
`ifndef GUARD_SVT_AHB_COMMON_SV
`define GUARD_SVT_AHB_COMMON_SV

`include "svt_ahb_defines.svi"
typedef class svt_ahb_checker;
  
/** @cond PRIVATE */
// Note:
// This macro returns the width of data bus that needs to be driven.
`define SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width) \
  ((`SVT_AHB_MAX_DATA_WIDTH > width) ? width : `SVT_AHB_MAX_DATA_WIDTH)

class svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  // The Analysis port for VMM are declared in the ahb_master_common, ahb_slave_common
  // respectively, which needs to be parameterized to the Initiators ahb_master_monitor,
  // ahb_slave_monitor respectively.
`ifndef SVT_VMM_TECHNOLOGY
   /** Analysis port makes observed tranactions available to the user */
  `SVT_XVM(analysis_port)#(svt_ahb_transaction) item_observed_port;
  svt_event_pool event_pool;
`endif
  
  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
 svt_ahb_checker checks;

 /** Sticky flag that indicates whether the monitor has entered run phase */
 bit is_running = 0;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag updated by the active or passive common file which indicats that the
   * address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag updated by the active or passive common file which indicats that the
   * data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
   bit first_reset_observed = 0;

  /** Flags that is set when a 0->1 transition of reset is observed */
  bit reset_transition_observed = 0;

  /** Sampled value of reset */
  logic observed_reset = 0;
 
  /** Event that indicates that current_data_beat_num is updated. */
  protected event updated_current_data_beat_num;
  /**
    * The configuration that will be used for the current time interval
    */
  svt_ahb_configuration curr_perf_config;

  /*
   * These are objects of previous transactions for tracking the active time to calculate 
   * throughput when perf_exclude_inactive_periods_for_throughput is set, and perf_inactivity_algorithm_type=EXCLUDE_ALL
   */ 
  svt_ahb_transaction prev_write_max, prev_write_min, prev_read_max, prev_read_min; 

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_ahb_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;


  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;


 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (`SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Initializes signals to default values*/
  extern virtual task initialize_signals();
  
  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Returns the expected data value for a particular beat based upon address, 
   *  datawidth and endianess.
   *  This is invoked for Write transaction by Master agent and for Read transaction by Slave agent
   */
`ifdef SVT_AHB_SLAVE_DRIVE_X_IF_MEMDATA_X  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`else  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`endif
 
  /** Method that is called to get information regarding the data/bytes for a transfer.
   * Currently tested and applicable for AHB_v6 incase of unaligned transfer.
   */
  extern virtual function void bytes_information_for_a_burst(int beat_num, logic [(`SVT_AHB_MAX_ADDR_WIDTH-1):0] beat_addr, svt_ahb_transaction xact, output int num_bytes_to_be_transferred,output int bytes_already_transferred,  output int num_bytes_remaining, output int num_bytes_for_curr_beat); 
  
  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Returns the data value read from the port for a particular beat based upon address, 
   *  datawidth and endianess 
   *  This is invoked for Read transaction by Master agent and for Write transaction by Slave agent
   */
  extern virtual function bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] extract_beat_data(logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] data, int beat_num,svt_ahb_transaction xact, logic [`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] beat_bstrb);

`ifndef SVT_VMM_TECHNOLOGY  
  /** Returns a handle to the local event pool */
  extern function svt_event_pool get_event_pool();
`endif

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();


    //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_ahb_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_ahb_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_ahb_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

  /** Prints performance analysis summary report. */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Returns is_reset_active value. */
  extern function bit is_reset_active();

  /** Perform signal level checks during reste*/
  extern virtual function void perform_signal_level_checks_during_reset (
                                                                         bit                                         is_common_reset_mode,
                                                                         bit                                         is_ahb_lite,
                                                                         bit                                         is_master,
                                                                         bit                                         is_active,
                                                                         bit                                         checks_enable,
                                                                         logic [(`SVT_AHB_MAX_ADDR_WIDTH- 1):0]      observed_haddr,
                                                                         `ifdef SVT_AHB_V6_ENABLE
                                                                         logic[(`SVT_AHB_HBSTRB_PORT_WIDTH-1) :0]    observed_hbstrb,
                                                                         logic                                       observed_hunalign,
                                                                         `endif
                                                                         logic                                       observed_hwrite,
                                                                         logic [(`SVT_AHB_HTRANS_PORT_WIDTH- 1):0]   observed_htrans,
                                                                         logic [(`SVT_AHB_HSIZE_PORT_WIDTH- 1):0]    observed_hsize,
                                                                         logic [(`SVT_AHB_HBURST_PORT_WIDTH- 1):0]   observed_hburst,
                                                                         logic [(`SVT_AHB_HPROT_PORT_WIDTH- 1):0]    observed_hprot,
                                                                         logic                                       observed_hnonsec,
                                                                         logic                                       observed_hlock, //hmastlock for slave
                                                                         logic                                       observed_hbusreq,
                                                                         logic                                       observed_hgrant,
                                                                         logic [(`SVT_AHB_MAX_HSEL_WIDTH- 1):0]      observed_hsel,
                                                                         logic [(`SVT_AHB_HMASTER_PORT_WIDTH - 1):0] observed_hmaster,
                                                                         logic                                       observed_hready_in,
                                                                         logic                                       observed_hready
                                                                         );
  
endclass
/** @endcond */

//----------------------------------------------------------------------------

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
khdVSCPqK2EOeRvcN1IddFaNOz8ifOb4Q6mktktpqHfWlo7Pdo+wnz3G7Xtk/29+
JiR9nNxv2PC1P7crerF4IAcFQxCQxNUtArUCKCNlW9sUlh517zqBcE9Y0bRKgrlc
PcLcp90S0ZIgwJJECMzfG+N7ybfl+9sRNpwitJ7iylc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 336       )
dbZkyvKEuJLSauPyxsFY5zs1EKdOo++duzKmI/5ODWVmmKIBQpdfGNvQ4eUMUEO8
bzSpfJLwFsOmioWlQTNdC0e6uri32x89Q7G+4z0Ycf43KDAnMMm3j+a1ccl7Lc/8
25IhJSI0l2noOeaqGB1qP0xFJ1GHFlcFKUTnAQUQPyf22dDA+whKnDi3A6zhlAfd
Mx/3ffQkZn4AC+GFQTWzuSgDCWMk2oz+QZ8Mc/Ra+JRs+XWiSqEI+AiuMWWT5a25
7Vufy+eaN7zITRe4w7Dglrp/5nj2BwgJM3Tl/ZNxmpFo19isxHO/gnBztQy/CMFw
V2nOP2NNDknMDFkyHb8iwVvzYkCh+KKMgVif9sPHzOTdtNOExK5vBTyFRWTQwiRP
f9/cUUdyh2PamV919YRfOo3L6Vfvnfh8KpaWzXUX/7uDdi4tyaF/7wDuVwzkUN2t
R7C+HQhi/4hwY9dDkj265w==
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mGOEH1Qr+YBOazICHU5ixHlJnHpNOyboVAwFp4S/B4K7rxkCcJd+96quVFXYZR0D
hWepPpFN+te8QzTm0gHanylIZghtTNXoBLnv0Tk1tACG+oK5OoATbLm65ZbA48SP
EAHqZize46rQL/8sE5WEGE+ponLaJgHmkQyDXYuyL5Q=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 28420     )
VIJoP5UzLOeWa6bz59PHG5oJv5l9jkX6v+bwm+/CLenPWfUmJoPYZr4aKM+ZlYRE
QvJUAthwhLx5exa+/V0FsLiPFL73LOLdkd+//0amQ9L40AdlqcGcTmBG08/OjTgN
s/LpKta8u6D5zAIqPcPghA1p+fzSNcxPvzAxG3hvqAnUYRdMrvzOVBsikgSPLP9W
RQA0AlY8/7+KsyFKC3ncvHwzCCz84Q1h6997EPn8jhWB+jO292risvfbjQ7yHgOY
SCGiPBZymkUG/6823BMD/ET6Dob4olHoRJmPl/PjTvGbY4ohoED0g1iW+q7L86Vu
n/kcfbC0XYkZVtTY4dG6x8AGRxsh7ayhdMR1grzcS3sK/fw4+H9DZQ9hYRVsQbsG
sanAz3ftEbqbsVsx03TDQreqi9yvN2XgwXCcRMZ/ZUfeBU3f8eqPZnDavPxbZ+iX
PKCXHo+dndPphiXQmFfkaQNxnV8hvODs3Y3bHyMcQXggTwFgrWmVDKZaIXhglDJX
PDUjxiG3Ph6LLg6Z/JSIRDm9QMa1bp5+Mef5X0moshFJZrfT3flfoiHXPx8G3f3m
gUpi1yt7pDrfjukVlkH9fAiMlqIlsdqrkGCiyzBVcTDcNXedtF4uLdX1hmMqusgJ
tcyhp1LC9SgzvBc6Pcg7wbTUETpID3+piyi+V57BXnwgemn1gHCUchaXdOo4Iu1d
TgpIgv7/7u+y2Uu/YJPUtCVzfObUbNbuBDKQid7sNFD0ABhaBQepisaJLtqMJd6k
x6xOg+weDbR62lbR8S4M77aZrxwcXh4fnfo6qT/6R6OG1RBK/KlwZ5ANgca6ooBR
6JahZV+P/2XPCj94404oxCEc8rPywuDW6ls8ab/N4NOn4/U06GJOkUmbjb7nEHrG
Tc3Hm4ZElZoyET9RkkD+MnniQjAa7d4VB5ULLGIjJ1yZJCMm0kUe6fS7SRvRKj6h
ISP1D+aky2F4xvuRH3xhj7kQaQLloeAyRN/j0K9m94/2QFWqaaiNvMZsy9g62K9k
Iw29aNRHlZHAuO4zIHWLsP+bARk7HXAtUsyBOWJJa3Zts87ZteVGzZfwUqDDsDZl
kKBDeTWb52flfxG6EJ0KmF4dVLDdS/gXrOGnwZdmoxb0SEYIAihptW1ACrQFzXyj
EcBGEY2MAzUcsKNJPYcW7BrE5zBuAm9Byt8deq8AgUpW4V3AYGYOYf6MiXZrRrSM
q/dsx2/yU1ey0DVx+dEa7s8aVEn9QOw7dVQWgju9Hfp8PD1nS5fGnsjL5S391dDm
nevzaM9bqjn1gl+k3hupt9cSrZ8n+3TrhD7zmboDCDseoWfve/Rm0z/vrua17sc9
wXOv2kIwEc/Fhgxt83vQZEbGZMhagn2rCYLgShi1/cgw9f6K+d7aqabHgLHe+zU9
f+x6YQy2ror0t/MZfsixxGMwGXtijjEkn4do4MOshV9D9MNp9116T9xnFhbwm5y7
WEjCgNze6eYIwv0Rv8XbhWZa0P5a7a/8neSTO0c1Ds0d0jzgK341byNDDvAG31Fs
F0fHW+3UvPYAJffb+0FNIQSXJHWqqfDhjB9pRTmvyNQ5RFab/EbIlUblzn26Njlt
AhZCP74IjvrfrDcTlBtvqFeUxKdKRQvoLgvaw5maAjveiNMnE3+dwSlU9q7KNyLg
9/lhyZ8z94t2zsHdzZvQK3r0CBVhHdX41t9A/vVUFTu6m9U2QZuhjv5T5yL1Kgn4
GQvE/0yWXl0MIVa/nI24N0tSOE/A7dzmdrPUT/q4E3YAnwMfsMAfRGI/iQpVdJKr
lfVFbAsxEoeEdaIR3p0HO4kF2zYyl4VRk8f2BtqbTNBSyjxx6RVeyhtFcvPuMVZn
fyFLTSJV32E8X8ZdO4aiqOcrOoJWF/v0HK9Nkb1vQw0PFKwmhuLDtcU/fQFD6W2+
pUTvKotoQcwWAFaj+f4WdWE9uuFUdf5nC9kosQhbCtyLF27oRu+CE3zssGyXpIT3
8vJiw3bl4cQy/e2vlxmFoa28bK2i7S55c2iKJIEaIQj7A6AdWEJrP0i7wNayrTaf
+Y0KxFJXnM0zj0J/cM2ECWwN1y7BSfBYxrAvfGMHUaeBgcuOm9ivjbOwTjgfuhKr
qycK9MUnuqYcT+oDr3dRvM4J5Bz8krQiAVVpuBQal/Nch76WEdDWEJbAcMbM2Fg1
/ZIXkghXZmPiBMspIrK/3JiGLhW2ulUqI/CaPfTxfoQvtZ3YafaQNJyJehqxZj6F
e2r5u91a40HZWnmF7K7CAESyAuW7Ru2Uvmr0hIPydfUsaVlgqUYQFB1zgrESzqja
j8LpW/t0MxyVPTuelDoaDoJQWIbbkdTVBnEfKnye0OfE1Edp9j8dNJyzLqbgMfLS
5olQB806ZZhXsTe5g+3YgfiURui3ItIriq8YW3v/0JNmUnj/c8PJKCTbO92NcZpP
vYvGtffkOVLlRTgSzNGVFV/zkDTVvRK5Cts3sNsIK81JFPrzS7B5MOusyD37A8HK
Ch9V9CzxwzBfK+Iu7xyaNejcTRLTZtpnBB1Kl7bqwOCDkVp06IffXHNUqzDVpM1n
yBZHkdtMNJLWp6Eyzw/yobriK8xguLzG1gqjx90z0qeH8PMv1g+vme5gqxoTHSYj
r80ocGWMmmxMktxITb3ZjlDccvOP4FnxlHD62irf5VUYiqzuRhxXCR7+n0plnQZV
xn5FWmWTQXulovOfT15b8kFMjydYrdJFtu32oFlCWerpEIgEiob46OgaZlYVFHqi
rvsBNO8r4qBBJNYN7JT4ebXCL0wIzqVKp7/zuqR2no8IytQOTtn/SXIWiLt6al2j
3JpZ7D7e507a7vJOy2ePD8bckW+edbejrLtHE6++Qks+wuajjTiiuwhzh8y2VrPA
5AY4H0c1N4QpEZ+T+BK/l2coL4LDizS3GgyPxKYKXBuMEcFaAAJ3PS1N3SZqq50X
vG5Nal4r0XrzqGep77Nr6CaJyftjBye92OIW4MZafCce+vwhwLFS+BNOfZ51vOsx
a6za7jdujw9qH8fh8FpSBDeAV6437I9WO8biiClqKDLzJpROf6m7NWMiqFhoFZEN
s+L1d1KTPYRzQ5ZDBK5mWqYFg1RYbPiZiXMzrfDVDB/CAPS+hpjluJxt2qPkSjhU
42vYnjH2GHxsQFmU/kf6+TNjtoUjIm+opwv195OArLY6F7dX42yyDyiiCEC/hOz8
8+myCIOVyWUhoNEEuxI6UJP7Ud0E0fhAZwZiNyAe/zdKM73Wq7LQ/vbOBL7Iuili
6Hgjrxc1UyuAjuQTH787Jie6bb+/l4WzK3k8dcCzQKKY+cwukEoP0e95nEwQ38GE
Dri193xXgGC7OUtT4DtzsysevXpDvMbOxibR8GUqT0Q1gSs/S9M+W5VJggoqsNza
QaQ/dbrhAGLK4p0n+JaFx7e9zTEKDIp7HvlqKC8+gDjSwt82zGjRIxDevBEJKPsq
b2Ri1L8aKsqNmC1KB4cnpdjMDEpyZJ0duUrkftsYD8XJWv8mym3Nx1UsHN7OvXPQ
mdTk2rTth4UXWJKAIcuPX7gRFOKzVCjsZXWK/fxTlR7j65sgeJkeqXGEgYoySX+R
Idhrns0uOh33ok08nzZjzvluN5fUR/S/Ji5vUWgZW5qeGNIkT0jtz6D3FPjoQQra
x1SA8UDqNR5HvQ5fYXwb8rMKZhy2VSwhh/iEuEaJ3JS52q9njb4LOhmknhajS3Wa
3pA1LSwf2CJqERdNxt25dMLqi2R83FYeT6p/H0uCSRnwCm/X6e7kLmyAkaeG4HrR
WJTLOpLhDdNmeAebsxrsauXDfW1ST52alAmXNd3gByi6YEbd5JlEUchMzuS9R657
JBuDDf6ALyAfa8u1CfABFmz4zckjGlJKY+TFV2qbK0trK9lxv1DCD52m5yr/CSEh
nqx+ftDxS5bA+/X9ntDXdcNOQvR2S5lhQL4deC1UoQoRMouZsi/EcjY1yq0Z7Vnh
AZJSeigC9XCAQg2e3qRX1AN22SSNgaFpULxqq/So+iCtJ3sHcMRZG7L4rWHC07ew
AJPav+i1sLQnafyWe7Tn71gaRmakLz7h+qS9CxAcHg4ueSf+Q6yY0nh4nxmrl7Lu
WdTha/72rcyzcuUWXp82QcFqR0HUzPxKes0AlV4wvMOpn+lQt2UTltgycpZlCr78
SzxB4nEBxRYwNPE0g0jBQAsBF0rdlp+fnZOz1XoeJ8BpMXeki7mXN+qCm5o2Xuei
HoyjCeuRxr/HXAt6oJ+9wWsivZOY2Vws5PH/IczE9nhaZzlXSQZNAI66tdEyUhvk
82LgVWY0QIQJ/9B/Gdj5XXvF1FwhU1bQemFOThbZkXaMOIDtvCecvlsqyp4e0Z3m
dKLGdejPa8N9yUYZ39rcdz9lwH167DshQxQvILc7UMyMojdXT/3VLNGIqYS9CY7M
SnirBHZmoZNDlI+Kn9HTEyqCKZXbjw/LbetR6rmqb2L1cG5ig4Sn353D0XOj3IWw
aUazXHHQlVGoowKWiYxNsj4NF8yE0SvLUfmNbbl5Wl5zsQ9mG1Bb51Cri8pPjAfb
PyFp615XkixySfD2uNcUKxWGuGhg77IPkso1YSayq7ocGsyVBkPQfF/20F2WYBFW
cCO8k1FCcQq78irG0N9wqm2XVhAjCPud37djE5LQUTrX3IkrlvbYtSGnHyYYKdoi
bTLuP2Ug/J3Pgiz8K/oGBHR1SL5Fnfy+YFDYMF64ZtPImabq7Tk/ke+H0CyXJkcQ
Ug7eJa7qj3+jzKX7XAoW+qVel15mKS2R/68TiIqpZNPiHQuz5VgF91IVts2Pbarl
jB52T+IENibFtThCgavK6+AwTySgUSev6q9Z9QljxgbNZDuxvAswoetyVA6hwsTh
vNssNjpliPZUiUWP1jZMfcFlfZ3iSvhxV8qjlY2nqMSzz8mkGebjGXbw2QDeefdE
nYBr5eQDD1oYrmENQLWEcJSa1buFFjL1mLOK7k/Pq4KoSId+fOABzpv5koGPHYMK
t4mmNr9QHTfbxbBGyUX9JN4fmuNF/JMB1c7TV1qDy2Bh5m5V50jiTABqVgcxKrcd
rtKBsrv1gHeYJ9GLTwTFTGzOPjLqGK9PwVUIAwz/7784Qop1YEfqdVXqnBGGO80o
kwEDN13Z6JrV1PoERfW1H4mCnRJBjVRRoac0Ulo6QYyoCqQoAosUFONagXaH3UrE
HBCJBsdJXcZosMf2/TZQXSb5mTJ36JS7DgLRhVkYoVmbuer9kq3fAA8sT0tEVYnn
Q40ktTQLWVhX4n6fP5H07AZNq7yoX3XFGE9aIGIIRxhC5hmjT7kL3hD+9KV/9N0t
wZR9aifkz4/SCPjIOHWQEt+kDRPzVTDMoGElZigKAmkSKNN3uETTjfqvVcIQ29z3
ZR5quQysvPrxglsjS2Je49wvHAbef8qrGcKYSBWp6jtlq8u6lGFP3rX0yNfVNkKb
3ZyJt/j2P99oGPsJ2ofvB+OfkBKA07mKgqQ37dqZwoVfAQj0nt0zOmgN944A3jNs
7MX0wbRLccoOM+QmhPx1ifbU5RoWUv6wfQ/xA0hSvDzywu60DNaKJcrEHFenoBE9
LvbwnsaCaynDomtc/SwuLFHu/dfOWBd7xvJDVKUM9RNzedP4kkvz/cKvPWi2TrhD
/5xAd7/yFYsQi4jcD+ERn5FJZOVNqL/dZuN7er/h/FDjOfaQq0vauMk/qvFOUQAd
eieiUGYU7rmFlu3uDNo9a+9vVfuMZOEb7e+Nl2YR1KPXDCyskFnLLsZgw81K81dM
c4zxSDEIlepWIrPqihCVZjM12pOOdcKNjaP7/GewXcVcNOFwCBZAQNNShhi61j3d
ttQSlPBEVwLNPkqJAdg9ZF0VL9yoMUTM78DFRL0u8kuZW5lT24hSVQcExVnmDR3Q
BWxKq+OQYOhehD9ckDlWw2A3t65JouiovPJHpgIh6kZdShKgIGzuBoq/sTQiKDOM
dazxsQXJg9CTzVmZNLj/Lx+3J/uLpobwa32+wBPrbWLuNNFudGy3WJq2HLwVGPR4
Ca1XVvHtI2TEjNE4hIC4xejGx8P1ZwK1sVkzcuwBiHreoBZbu12LnPfjbWZ5vo0j
D4zg5w+0K9667Rbf4HnICM+S5MAZnCthFY1l3YK6w4x4JmXUo+z1m3u7u3WQYUKm
15ARQwQr7RGljVzqd1GEHLOg1eO3hWKZ1mOYg6DEPF6Tg1rm8L2RJETbLjaKmUry
08Com0UbwUGf9vYUTsCKWqV7xbWQ3218sBaU/YcUXLJWz06JW9tYfL0oeVmkYS/B
En1w4ZF2XBMlawLrVEOADG2TX4Gqa7MmW7OWyubAYWB8kYuNUvaAoRC0rzqOFtdO
2BuCmau3GyFuef2b+mRzzuBYWMMjb2PkAjorD6q9wfDOjp4ufc6Wx66iYwaBD46a
eJVvugfcu7Hiv8r/kx83zkmNLIuGyVimID+dnHDydL1cqociWszq+9Ro8YIwNnp5
n9KjoTFfWjE10OUTULgJsx2fK3zRNum8CsUWV9aMLnbcvWSSChLBkLLR6DNyGKEI
BoGFiJwznwycY9r14XlP7vawlxwcqhjLAPV+CV3ohqDwlJ2pO1Jnmm2rc+9dtZxh
HyotYYE1Qocz5+KuYFR+glKk20TPDQiHjbRIZcqIg/ME9HqZJ78tObeH6stw0UhW
aWIsE26m/bUwJcNagvfKeNUgbZ2NtRoPlrpUxRhM7NXgP/7tLf4BRAlIIe6ykU4h
87spqf+64/HuMxphLLPPkPUaB7rOWvmYYhxdF907K6AbTkofVwW61E0WTP0bLp4u
fDTaP2FtJhoAxHomK+vwv75zI4nUw3v+kTZ2Bwufk8jGwkW6vsIRctyvG5BwSx5P
MJglP1kMxE+WoroRFufuLUFXIgK1BAUI2d3YwbxwOB9oL1Rq13i+3ehQJ412+m4N
NgWEFX7kETo0uCBhQRpOLTtaO3csqlw+Gg/zIM6MwxgGQOU84OMk9i6ol+PRtFq6
53ePeVaBuI3izy8YHzxFbDLjTQ1/c0LviaI7TWUBAS7oV3ave7PiIM+m4UFpXtWh
+0xs2xg3Nx/h48DBH8hX6in2V9eXj5tXDoDY6B3YvCbLO+WGNd9EOq6ZPmlhK1cO
0s0CZQldu47CqTADNoOw7FLBKObPZU3oZ264Qpqfv+5Yn4ZTrpXg6m1d92BSFYV4
CcEUnb5ldVAMhkYexxtQ5d6Uf8TIPrlDZssw2iD7lV9O/eGglVzHgbXVaUcZ/M0F
oaZ6jsW75IW95hdAil+Yq25mzkp6n66LEIKVuuuJX2yUQkMlcMLvHfyywbzAUocG
kbFaeSebBlrfjL0+pESfOdPnz3OnLBms/jwZblPlaE9RokbjQFbTjw5xzjXQkvJl
ir7suDHngtbXUqEDHnb1yxBykNaVJ5NpKK17MP4wxbP5MwvSDPM/N6DVO1gdIytu
uL70AVlp5NKq0T4KWiDQQBGcyA0wr1hTCcCHKji/HjFtfdBGOeU+chNNh55f+Q2q
zhYSK5uZ+TWuyQcXKJnevA/HD+hJFBsMvhnRWjnLWUQqvgAMFyT5zEi0zKXBluT1
pAmEQgxDIedntm0uK4ZlBdXwfoEYGg7QeaLbJ2UoWQRB3ZYOskLEmvE6v+P7vknk
rVN3fncVvhYzDlaKbLPaqaHtUYZCLwfhuHlLV3VwAV8Ul6EayuL2nEw4IYztezrF
HtSRWQR1hCjNGgku7cZxxvVx4I+F7Hn5BPzpW+82na2Sv7ceAUZdVZ+6FI9w8oQQ
0CCPE7Bl+OrAwsmzv667Fqkt+9lSooN9gO9SGyYlHG4SieM6hvAi3yWu9WfKtt67
GMPHPsUxJ5TBsPKnE/UHRe9z1SVX1f7P5EiVu135Tf9UdCvny1ZSpDzoakwi4L+F
6rN5rc0t8E4y/dRmyhwoGWZLXP7qCVZb/H6sGSBgbcjw9KgK0EdLPQGF/caepZd3
Ux4QTsconHylnM9fCmeIWUmM0yj5P6PZyXRi7wA0w0C63yfTHkPUZ1LNnXcIZifC
bamkcrtspyJLbO/vqpumEEDADfzAA5uzUukBSEFV0cGQ2sQzEXcNnCB8aZXIynsj
7WuStOCXJCzr6YW5boIigo2M8d3/dElEBv9HUGzGTpmlVwFD77ouYLRjExBfK8OF
UPzqvp+SkDq2u/6eoipvnqGcqGxuvGz3TK0pA12E9X4QmyLM5ExerAa7V1lNWzcA
MO8Ra06O2YYtWwxde4PaheJNWtCIaXpxvsp/58Ty5P7NV2SM7fQBpmD3c6qjRVFk
/Gi8VX1UGSxTCFsnq7wrTZWkYvUSELv0wFx0C18RrXNYN+2jkEAAI/Jnz8+uf2Fu
YqPRTsxxotuTG0eyNtsgRtf9Kn+QJEr7+9SOTSS+sWJ9Sgfnl/RST/woAVVux2nk
xQYhSwEMip6kqb/vMPiy3xjn17D5Ji9G4RasNrioiggY4zuJIJoUUN51CENyuiN0
RGTMDQXMAxdVn4athzli016wzuImXJYh0L8sT1Zen0Bgz5jpngsIIJ3jwlYqBQA5
3hmUrKI7K40P877J7H64uouKwO0c4T0ZquGe/Dsar8EIrbZjcuEGuoJxTlT20/vL
rFABYCI1eUWYTBkKt1hzPsDpACyzNq+MZlt5pCWtGPOmGF8ZZxJG9Q/olnojHD51
u60RDamhJxSqqt8BZNe3hCo25PSuB4ct/usSglrC6yarLKOCZjJqa+gSuOygzIyv
2q7jmPdN82IAeHkZMDcr+nwy+k+A7bfouwCZw+YcBsUL3wMEc1diNoh1P9ux7VPi
lr7GrcrWY6fBfE2CcHMEL0mvJ24zo1P8o3Qago3kb8FxzzRdc6qi3m+2JSxK1tQe
xCLTGhW7uqEPuCzqnqZohafWxEnC/j0iH/b2WW0WpGrsvsKPxp6IexDz00LRrBK1
+FfejhQaXDPoiIz5E5Wmc95CSNTRK7CvWTMhJsd/UtHFniUfT11Y5PS6UMrBBBec
YZSMs+dvlr6pFgpN+MruRyk8MaCz8SndHkQFbTQtk69E18mRNtmd4ZmKXcC9oYBP
s7Zfa4+35Syul9EipEf+eq8MdXMirrZ+QGtDsl+p6k0vHXRHUSTczcwE7rg2e8BI
7ZpO1CdMmfilWwTid5mBKwWppo1T3zrFA2Wqsh3ITNpfvsGFnrkAi7lF7/kw7mkO
ErEZTT4NLP8zD7VpL+CplpYoW4KFGdBA4qRk9W7tf+rDMmcDXwu3Aqg1B/Gn8f3T
9ljzG0pSxeAk6EHF9KNSaD52oJp+blXIrRLGogRNONVl8vN2gAzQZWns4KpZQL6s
7bUnHM+GlZKgL/yLfbswZ8LhrPVHoWSLNZqBCtilXm662E787GUHyz0Wyqqua85B
FAcV/tJ9AnnOvU5uTwZipOk7PZmv78phVKJhjKKrj1fqBLffJ1gDSiL3VdBvexk0
6LKCgJ+wFx/6wbvQ8QRZ2XLse/FG0hXeSvZRvsmPxHGj4V/TR/ZOvzPTiTSJY6Lw
g5Ia/C1bQQlXCGaK7eovCD63kSCqVHc+rvbpuJwzltxwXZW8RuJB93ujj4KoS0yA
wigL34ZgH0Buz+md8TOwW97pvcvU4bDeqRTnosfbofbQFHAhDBwH9lG94i5kMS2i
9EHAv1PXt2xpx6RVrKH6ApUmb+bD4FTJqdAz//7yz+M2JJ3kzB6qo3gm4Auf+5UG
uMOG41le9E2wjbB1cElzkwFWMdgM8nQLr1z8ViYjY3v+5ufX8K+mZxtUZloIdM3A
UV+hSF2+HAFNPeKMjRVEsT+lghLfKAxb5HhVykWOUNRrFw+JOs0W8qD73Id4bPrI
oe7Om5+rhjgKBDE/YrcVuZGdeOWtkGe2ibK0CvoaSPTrwPCDADlVfXw78KJBKkzV
ppdGKtTKdZb/a5vLM5ePwPgSeMS1y+e9A8YMiV27wXNyEHaNTHTVTSknOSYeY43z
Nzxo+9XuecxS5m/OT8ZnMkc6cjDhc2kSmJObaWX5SULt03kHFY3QJnPyyy1mHiZU
DL85tDXYoF7Bs+9iinteT5wzC4HMB2GGtCeI7pSJoh2iKB+eAuc8RHiYx9mjNC+/
67o6z5ElfG4GRJ8DSxTWz1uWA7KziIW0LjplB82+wNkXBPdMDHVe7JEhB/W0eyr7
xUKO29dZRihk4Yx4dq9kNzG9cId757I3WaXCy3lGCT66cnKgMrVg7ixQ1LInV3qI
GiZ+9A0Y0wJWaq0i4u0jGBUK70MQJaoJnPDaudVhKwDHbyZwQBD9bVPN+Xb/5/7S
IIlmN14bvZy27An9gLNlUeDfRMffDnYf8W1cmpjk2ECSBIvnarXFL3Hj+ew97qzL
tzvEnNAFVJ/S1Vtl+XDihY76H2KNvw/B7FZ2BoOo5gvStQkllFySRfW9YdbvZiM0
fRw/uJ3qs27D86ZhS/CiyTtyaFxsX+X3ihDHYJFRV4jxIsSDnInZH9GPp9vxgLGw
qJNC3pba/FlJdGuvUmOeEevc3SAh0uO0P8KQch4mAKf+wYK2awrzSDJC5yAu1aeG
8Oe3ef6a64oXxEO3vpQMAt0pgwo/3Oju91wXikq7w3SI5Dh0Pg5sYyOTscfTELMb
ro8HM/ILIM0BkFNKr9icccnaJIzktusoxo42AHzLLGeThANKJGdTRU6a4XAcE318
2XHj7o8MEaXKto9rmDPd6ZVPwNLAGsV5129DLD0MKMzKjNvZh7U9cPVjOav4Uy12
5gUjXqh3bMYrTKcRAYqGpUWs+PiYCpf2dYYX46Kqy54Q+lskMaEBSQBlHPDrk/nP
EQ29swELd8VYO7INXALPSCv8nquaHfMhtx8ZMWjKDXLEkTb/5DQV3xVQKkQjIBRg
3cklsjM3A4zvk/anWTb/KVlxF9hKbDnnoOFFcaNTS/go8Uh9KYIrGbbbI1d/ELrq
U8qJZx6BqI+K2ND8n2IEvi3V+8Kl05FUHmLtX/mcDJnUJtwfwsSvc5/sj5RHXbOd
duhArwblbIsC8TkMu04Ay7kc71ImuI7+MlYHew2H4iFKQVz97n+j/mwWA0sQl1ym
a2Gm2Qh6/BAj8pPAMuILVuFpgln9wV5OirzPrm7x7i9WVOh0negVnUz41309qiVx
izA9qqvoKKQcI0XcTUx9pNth6qINt00mOufBoVkyMU/9jImursQimX8IEnxffiSB
5xoLHS2uc/gT4MzdIkTHvUIsChquBl8fbghuqSsFxp9gDrsbdQ4AIm4HgNSQUZeM
is+8/BRTAhEmmAZS0rwPa/7m+u2HEU5yGu5xb0NC3YmI8Ppf2Br2gicVdVzZIkrV
PeV456uXaYtL3n2NowkfnD3rOr/f8BtjFhSsGsbVeBnsQSJm3cPoGmd+/6apCJSE
U5BKvPaxWtdzThe7Covn/hns27a/8MmTRoxzE+tSoVriYnyLWd9lxBPoseOVOtpE
d2tJYm20LuO9via7Z9gNTHnfBHSdMeffta/8Zk0LYNAxsjVfRPS0zeDzNtFLROfn
yPXOqDwfe/NgKjI45SoCP2KwTakFCBsHumaFsmA3IdMF3EgDj+Aa+CMBKaSI5TNh
W/TYFu2Oz0ST5jPWfzFP05fGiOQYKDp0pvTLEtK0cZlDMViYoYQ126SdoRwPT/MR
Ee8yC1NkwutsARbgCxkQ9Cb4o2NIxnC90+5zNvaCaJ6zp5ZCVjjeX6wAiyml/Yf4
ci1Tv7ID54myKCTYbbM1tJbkvXpX+H9NvaddwQo85zShBuZ52ZJu4TtqZznWNmlb
O1vRf7AF/FqZmMaz2TtmKgmZuAaPsn7SSHz+dj38Yiz4+RaD3fg4ZMPA0j50PTIP
1lCSEWRfWM7TztzN76ZeP4/7+hADd01Si5CQQaZxD2UuIfD2roJ9U3fENPM+fwZI
Jqctqjj3DmYMtnotn11o4wWDgHIt8+bKTclrDZUf7a8sNdO5FMmQPK1Kng1JOG/5
jwdFBCqqiQ5P7O/LxTEUz3x8kDn5K+tezX8X4Gw2DlVLN2w4iZJ4jtc9+uZSJfXe
ReUdTDDGCVneb0lnSfsIkLA+b9fAva76PTC8mYcPKCMzxPXBS4KgjeZhzHTH7cnq
nDhLVTntj3oBBaPng07aLr/59l65UG4Nb+K239+LogHa3viMjF4SPCuLbBxpvEGq
vbJvUoS9IddMyONkdPey9WAHu0GOFHbENl63q+3Mxn8nbLM5J+RLtNpQf6wge0N7
S4Ml/HxCFlgBSssTF12WZltn9I383pIxMEs3hI7q9C94UuH0VKZxdnw8+dMPGfAy
Ejwxeqhk7CuT+yJCrT/q3rhoOn6dwfPBzTF/zWzJ55/CI8yQT2FeFGJWKas6i7xb
eOkR1HmA8CSEE2C5BZnRDmA1KuxY1r4K/kcSPfBsjkxdkRTKjZrzWHdb3xMc/lJt
ePPDnhPnC2W8dxkw3R9MuluHwdTM65NbM/e7fhcNw26ipHDThR9YmH+3lZRTkYZT
YNsLgul7jKdMitjpA486Dvh6/c1yTAgNg+T2v/sqQkkewzeuoKjetoku+r09XARI
FDq7Fw9KQbPRlPbCAJP/QLfto4MysIXX73FITQ2E/O0yjmZ0CkJKD+GyUXGhmNXC
XmZRgqjSK38QpX9HDTlhFM/LFurErT6WOqSyqQjyLKlLkVj13xuGHE8gxNht4q+H
GrN3WSAKfnXBC443j/HLIymKcepYrP18CeP51yidUneTcErLWYLmknyg4fDk7qMB
1YsSmTcuVfsy5InVNeQ4mTjqZkZiY4a70v9/uU9xuq290n4S8OS1vEEQ0SH7VO9O
9hxU4RKi94G9tlXtQWgTOS5matUnr4ggxa8qkzIT9lOpQBJzaltXX9n0sovlad8f
oYGRHTDVmRH3nWJOp+XW9luSUjBDTbUHMYJwSzkKAArR3PN7FbfmiCStEpbtnhPQ
YQ9/m7UsCHnE1dxOpvqzct621Uv+FwbAQOIsHo3TyRavii0i9/j/lLjpx1n667Vi
rqSV7kMfPRw8klh+OcDiujLyaXwqe9diqRCOglPMsqCpwb/pguVjvBGmZpaju9ZR
LcUcCgzJT23yL0ST/zaW0/YwHXuxQ6pNpwqvL/xJBX+wQpAw3cAIQmKRegoR6AKU
OxHD1sb+YnrfrbdaySmkgQtYSVCCnSHithrhTvuP1a0+xJUwIhJzTmmJAnJm0uTq
mecuHkv23WAqXui1ENAYtWt3+L737JCw6zX80ordX17xLe+oJS9xnUf0IWnzRn2T
J9EvyPYbjh52f9RDA8yNtb75VJrkhXw0EhU5IPMPuMstX+krQoPRxqKSR8zf9Nc/
U0gOqP6iC3kRad+yXkkmFTc4WtQT2RNl/3OxzSejjwG7ErVwfus4KjpZSrUpl9rP
dD9xF5LFxaW1LActeIQ3fUXw5GDQE/u0i5xZwrlj+qJgvfyRJ1naFj6uwk7QZI7j
3KGiRe8vUgyNzn6PjAy0MwSrg5yqLlS2I/IqBZaRYc8QE99LVJ3sJY51agG7f9b3
UeqXiI548akjoaA1Bm84vC8IoVVVWA3FBXSQ57W/dBhBQXM6dN8MLT/zXGKtxBqD
6ZU7536SB22tlEKXd7ouwKpRDvHEGvZsPqgGrL0MLV+G1UU+XqscRScI6ydpB0vd
MCopIliKlNR/RUNOk7Sgr5F/VcmgTcidOiiuqE/qjSZJ5aVGWa3YSanNV0V9yBaZ
MmTMTYdrEKUHrs4kIk8resp+8cIhrYfI1FqMNkowFfhKX4fyCbZO8XMIy4MeiGTA
MZDPjgmlxB836I2AGtvzdBuVhDvJOUuWpBMxjwu7vMFGn/cjNaonUns9P469JN6n
aS4xFEmBQtt/HzCtU5zJBT0FRHe+UlH3DXomqi+tVnloq5GDj3/kd+WJiW4EOBIA
7asKeaN7f67GcDF56QVCVsLMjkSbyRJd06c2CO6StoUisyaEdQDvy/u3M0KtQSlw
0qAWlMUJUN62ylLm6Ie8EMYBAcGmDfrHtE5oPl7eWdhF7y3xtA7HTISov3iZyVac
+5bfZiHwBjvnYrCvxLx1K6tksMW/YUwhQkk+pp9ajM+iTts8ea1qGarhWkZupH+3
L3Gz7X3Nxah+b/FsO+10mJYUmjl/ZX2W+tHUbh1CInp8fkYhlsJcAPWM6SX/nwvx
frcXfiGsidrHxaE91QYDW2TBtvI/GbQOOxri5WHulS3FO2Vjq0jzoym7mqsxmyxF
ha4ky8qmlsvB4Dz8USDmbxCNooScDZ4D31/M32bt4j1w2tFZC3Tv6keNa0vtEacW
59ANlUAipUuK8h/S6/jnxA775GNZqgbOoAPvZd9o4AIYzHRwLaAF5jbCS/Cp/USd
FBdzrDp6rwIFmQxrHNdbxFkaUKO+vroEikle5166beVwaedDp8Kw3zidvBznzh1v
J3t61k3Vr0UknuK3gCdaXrIDcH8g7pVnZZcJmJxsbGduc/27FH3WuZAV1WO06OcH
RB6kzp0hzhUH4GxTh0IqY+lVmVxC4YgfegkWqk9lLO5xwPb4bOpv28V5HYKo4pIn
Bc7QbpxaCunXb/BV7qm8UWJMBbvGbhq31vhPM6JQiw1485iCbMOlqy7YpcINud1+
1Lmre8QB7QqBlnAIUrVYU2iINmJE/jkVCT9ln0YPQ6iDBOmc1Zz1+GH3UgiXkshN
ZPG9Y+tYHq695KmwRtLsyuGP5tMJzDO4qEMQfAqNvpFdUgYVj6s4IpXGOYzh0zvw
E6ydXapiPl14OzAGjRCZDS+Byd4Z7dkojVXnlUKQJTu4CaW/jKTLWj3Hefy6ILPu
T81Gy8A+GJVOLD08meMao0HKBUea10rEgveJjlfdX0TuHg5vXqUjGYkCLLrvffT5
v6U/uVXu84icAVgT5sg4SU8nhATsUgcXoOlH2MCULOsC/YJrIvk8dQM4O6CCchMI
8RYZGhxDE+mmeu+ZFuyiNpAEpozFlyMa6e9AIn4HACUGnpYUWWzIjq+B6Q1vqjVN
sC98m8JVa2UkqyRvVRF7hX8ySt/avRcrtDGPaIy3dxe4sLBEgAVh8jB2NHIhsuKY
zrVS+p5GdHxF/SNN69VVDU31qreT4zTyUCmbUVwEyYa3+LHE4QKfsfqvVmJmuXpT
F+DJrGytZUwo4Dxsmbky/+CNVtMxdgbtBy3ifAbNymFU/V7QY0UYnmBedpfvIaiW
fj0roiUS/CObl7T4eMFHssjDBmgsPAMPrtrlvl0kxqTRFws2blrymZ3dGrbQTttl
CZveX48upzvUlw6y5z7zVbu1eSNUXENFBzmTV8cBrTzfCS6ZVvftdz3wioF/EQsI
pBT2u8/bajzX333T2GZCHUxs5hOva7Y6bYxp78eDmzJyPM1a6eqfll3ChlCGslrt
5Du0mt+qiBGL0XcUwjR+WrCOpw3opj0QYc7J9Zy9R/w9lb4i9Lri2qF5lB+CBQse
2newcf39F4EjERSD1UrZ03uc8IzaXWq7SLy9wP45wkN5+mUhQxT9rVkLVqI0BR5k
7OzBPc/zsPQ+hQDbw/bJrgSUqzV9HQpNNUs2Sxv9OD3Mfgmly+s2UiRqc+RkXnnd
foxDaJ3zhYfwCNAoixncGOjO9y8mJQ9pD7/VSJ30yvstY14a2NUVjKY8PHl15eF0
ToIXpzcOrc8dVCn4rjonuQnX/65rI9+XZlfCmSnC8AsH9kHcbBuj3CPGywV2Lmxa
5WwF82fP9JKhXQP9E0JyX1OH5/f1L9MDzb1be9zT9Ng4PNgT74NGgA3r3TY75mwR
vQRbo63oD1vJ0E7qMeRR2XNU8ZfUiSk1mN8u4mgwx7l0PaamQv/AJfOy7UrajKV+
IDvxyUuqXyiATDNTBvQOh/wLv6+bv7hnOtCeTSd4nZQjAENeGVnhWiL9BUJsI/mM
i2EG2GcCoqjNKCob39Pulx/UR62mGx8f4oGHtiTDoSPa+wsR5ZckFc1khE3d1wPB
1NW9i8Uq6QLfdCNwTqMh4kmvzVkiQ/RefN5xrYus9jU7VVbvFHHbRFqtdMC1oBGJ
/0PhTFEyHpptXpRLh8yOxt4SRpGZkWFCqNTYb4RwyUcBOFyZfiMLPHfoCjQSyTtD
qw59lxx7d/nuxwpcwFMBBQWS2XJkwnPozAxmzObQYw/cVR7kz3ZppNaGvY8nbMah
qNw1WcxsKTx8fkDiWaKdXiDCJFqC6XglL2QeikSMJSk2ylTWBYzYFPDb0qi6MCEh
Mfc05GUtLxXXuE1O6qLThuR9wBAQ46q8lKhBK2wroSBNZ2jtYTpoikhFl8epGJEc
2JMvCQi8MSpmdGaB01BHFSx23a11foOEQtIM1KUH2JFG75KsY9k0mZwtcw+UvXwq
Px6vZVPaUziUDd3Cy3Wwmhn4LagIIeP44UfULova8D2hB3n4msgW1PpK1O8P7AEf
IztLCr0qrttc5iZcfB5Tkxo3p6muL5vg6qQKwi4wjcszTCBTsaqftW3h/JfHSkiE
T1BMF8yhhxdwJct1/vYQhFWcDHQILmT6ln1veLar/74nrEP6PiA4uiRC5h6IxfyC
1NaokEH4ilAXgrb1x6HeGTqfutZOG1Ob8HBVHRpNcqoH130oogwxAVu+ASSWwW3F
BNsOgcxtjh8MiCiTTVSbBg4EQII5n8q61QjBHzAD2gHVRHhz8SIBIrnrfjZV+bKU
DiIYJ0i32x2MTT1Ai13HAT14B0Wf+NLfmN9ubPj8WMKUd79Jpr1+xTCXg5UlUnsw
4QS2EJa3bW43iYJEiqXwcm+uBw28z1bAWqJIYIr/oqPxcKgC8G7ecLNNgLX9hcCz
gJsGGrUrEXL7AOdMwupXVPEagGXeBiYsiFuzSitimP3z5SEJwI38jtP+r8ROKCA5
qvrJrTa3cAEd0MmoPk/k0sq4FvTJV+8zCgoKa7bNycKm9WPsIbtXz+GwkXR6+xUS
2EKdJMN52Tfl40e04fUPUGN92rN7CxRQqcFPlDCBnWhGCS4t6HX6FvPiqaYgz//j
paO+COzHRESOYEpB4h0hVTrDX5bH2SvfA7usqTWdbXO/TjIxctvUi9avoJsPNeOv
0RgkZTolpnuuNS4A4i+opuJoTZOx7xzbegl9hNrT7CCDoy3xln7Aaml9sWukz0aZ
qseEoORd7hC9A3VOSuyU52hvALTFOKFd/VLBqaOGpbFxYWT6q91PAlGmqEqxwIZo
2aOiF/JqnKRJULkLtckiEp5DnkSdvV0Pg896tVS9vP58xX5X82oOKgesQT3jIWKl
RDjJ9vJr6sl5OinulkKnzz8suKk8VrR03CsxaFLZAUSmRSw40tMghLDMivNR3U8r
lZphrCipc+VL8LTjtgYzQMDP3MM1b6wfyiATWo17ypoqUjYwliWenkBmf1dvFEPb
tVDrBCTfnypAW6XZQFD/LJnceplFao89xnPfGe5acY9TFXRDsa1hcq2uHLdel18B
vfnZchWmm06+zAcskVIwXD4ObctHXOB8QTTUBBd3GdMuDikhg5IoCLlbj529ND3F
ojMEMJTBsfHCr7IcsTOdrSVBw9PlhUaGg2nXkZYdU676LKvUFFxDng0kiB+3LIF3
lxVvYof6DcFbzQA/62zuaM8SEsiIUoVT5+PhnVON60z4StmIAV/4rLztzqndKRSI
JxSVZWL1kQ+uO3iVzi/wROsQnijZwyX624GtaK9bcDKCxbszKuw0Mf0fDs+v6aFh
NytDv9mC62+5f/hGdAYAHiU7MTR0N04XscpQlON69XxSIvkpca+xybrtDJ6Jipfh
R6McOa83GZ0Az5pEEd4QM2cO/2cJgad6SHooEcMVJwIs5pGyLZzclFnpFy4sSI7Q
NvFqLH25SS2AsGEKGg+8dJcuchwh0iD2Z9GdM4fX0onQbcmlVFhOj9k35FaaLDqz
WISFww4OhbvhsuvP5uNG49IAGRG+B1V6ctzSglKF7Y3hLIZYiJgix5/kW1wXKPv4
+jLUFhbqqFMNrVUad/Ml4B8da2K4BP8nMw+Q7znhnHs7nsxSuiXbqdYr3hcJ1Tx0
7Yi5eM1mBXcDWrsrLD70gML9ZuX9fU7Gvcy1zpsm69dH2GqK59Gg/Plk+98ukMt5
AN8F3MTHaXv3p+ZIkGfQQjFgJ6aEd0jLAq1flMjWGezhR2rH/5yf5w72OfDnQVs7
E2WHjzqv/qxmTgqRijywO0kCW8OfV85xe6v4fHafotyBLXi5qbkfbWLWemlnafHX
zadkoC700ii2tLSrpjqV4zoVerWvEhgliY+Q/1HANkrrcSYjDuTSto1cnZK2E9QE
mv92djmrZ3Ev7BgDgm5oW5q5EcNTtlvqsZiqG2Oae5EK6e3hQIFWJzMpuzWbM+N3
22aveB1AR7kcCwTsUys/6LZiJvEEzAPtZo3ju5KeQI+icZtB4g+YUcUlGSWZT/fM
SX86kLBwNIWCy4COzxa/lEPDFxx2SqvDD1YRnfTZvc1kuWa5Z+sapS1dHQD//1aa
FFUjAbSEKYE93LNSW3w+DVGVOYkNzFzahYYQwqD/v2o4nc+VItxNAqG8AnUPmCgO
7THd7QHhUfbCWiF1ZlTbTZ+mSCtzPega9j+dfT6DFiLNQZ8zuJoadlhdJzUgYsCy
TCEzP/tsSmrvxtaNpfXXmqAuTvzZm0JkRjy5cKQZi5sKxZiTEtvts4FeUbqS4UJX
CCivDttFOrYFjjkp/yB3vHcYlgBVWhAUE++aJKJ6OeVXeHsCfMLaxJOJzdX9iNUc
JQdO7lFbBwDKIPDqHFb9QTvj5Yj/KJFuTYZUptv/3xcA292geT5oTQkY1PWFkLGq
/Gnc9tviPvlDD+SZWRyKSUQCidABl3XsA04UItERvLr4GH1nXt3ur4h3q8OJoeeU
WvZU1F8Bv7bV/1eVa/0SL85CI78pr2LvalxMTQMTOTkZgsKq0ijqJGYD7ThUPX+D
6imLmN32JHj22kxMXzCtCWyqRjOq6MJrOA9ABOTOcIO/cTCo4vq3YDJDmLgK6Nma
KU/MHHW50jE4Y+cVMwrL9qvj6qECZoyU31BgeOjBVWkODBxCyUdkY7/mU1ijRrLt
ZsFjeLvE5RbqNuste5AnvMED9sjWI2joAocAU6HtMDodKRfrSIopB6A0mDo1ZfW/
qVc8UwIuuudQCby6S3qRQoeSX6pjaUJLrkZma/Qc1z6CCDVCQkgR7TQEsLeV8FAm
tY2rGekn6/OBxS45EQIN+QGxFVrm00GH8wt3Wl5PiHQPy+CwnyNvgEEhMtEeA9gU
apONUR0bzseZHzsm8JnrJXre6jdDpwl26slIZOSqXD/wbRI5kCNJtd3FnFYUD0q9
XGaQUnCfjJ2/0mGqPk4Yl/b0NSHpwFgfgwSGgs/ayDMeKV92IWLWcL5zASjAoDnO
sz1ICeuu4j6lIXOfobcPhj+mqZpYoEeJ/RlDs3kE5svoH4IJTjh7DueZpjdodNcH
9D5ZOeLvBw6EqG8YiNvMzvnVVttjZRN06QpwwQXHR3WXRr9sDuZCMphCXOcvoBX7
52R8RAdvjuacIXS5iY+x5sBeu+gJTJWTEHI/PhXiHuQcHCOaLlFgBC90WJ+xavX9
Ecx019Y52qAnBcaj0tJiWbZLFozU/TfL1UFMUst9YdxB2L64IeuTWMPY8pgU3BUI
LHwNzXLkvopo63EYPfs8+cIcV8upaVYnfecp173oHMEZRPa0wKys3k1qYy67euuQ
O8WmGCas6bsBwxND3bL0Wqg4agTrIXRs7QBtHLt+ii5EouTSew3ifwbBWZvZo5+C
eethybyd1e4LxWs9TPHNMu22M+o7qdCSVFi8WYLp2DRUHvKV7vGOIkdjs18uc12w
7nJd42f4s/x97/r2W6OxfoO122Mzv6oyTdwDcRQOcs53s2vi1Rqj0t0Y+S5771xT
H67zpxDKb3SA7XEU8DBY5XnULruqduda+iusHZUtQeffZWCNtet6YjGC1o9mPfzt
nK+JaxwNjchqEsdhdFabPJmgNaxv6R1d3xMoQ+r7IAp8rBIjLwXkk31LkAn/Hxfu
/EcaPi8epl9/RIVXpINd9H2BxRmCEVG/wNiuDyZDssqUE28FndQbOu/d8rGyh9ui
IUtAAlgwi8P0DoYJ1ukXUUIjnUe7x309NfsUiqQHVgjKvT47nOKgCAGe0jsNx5DA
YlbM7IxI96Z86lw92jHFqZj6K5XOGmvHzgBtmBMjtZ8NhSumiP/F75CmC8jxdNfS
8z3Z0eKH86CXa/iYDQYRYu7sQ/qPA26HWrlO5zTY1brP6bMEik1ZmB+45wsHl1aY
wGRyZ+x3M1tDskK9AB8t91Lv5RtQ8rHWErEn4/nTyq/VXWitNH35cIXQZWs608rY
TWM+sBTNbxp83pOgGUt8VFDc6SHIgs4+8O/7UMv7bp0GZLyohwFSeL05Aed6nKnr
2cHKACopWqYp6ugBuxfpYcilJe1PLyC+LtBB0mffHzLmWPPMV7MnMl11HWHVtV0M
J4S6SsAKqI4fpIMSajIpig0Gx9ilk+uxZboyw3WLLiDcVRddR/unQ2YBOboVQsn+
fPXVkQhQ+fSmK7UxdAiGe5A4sfd2PkOnibt1Cd9cKxKqQqHhD5ZoC+GgM5aBvy7G
VaKiyz4aSE6seugg2spGAWJcqvu35mkhrjr0ZzgIIq1l75yO/giKnpm6lg2K1WHZ
slzkGyfwFwKuFxkoFdrFfE8zk3HhKwW5drSBeTPhgm64BKkQfF8lWx+zVMqLXeGn
Nu1jjKj05RFnU3LB/aClsYPevDa7UsOkeuOv21H8x8W4quHrLGJk+OjjCMmBZcqa
POguvA3uqeeA28YRj/Dt7VpOg8LwfcgxM4H/nM459sWf8Dl3GrScUza5cu1A28cZ
siCQ93R6avP1GwQMlD8Fb+XzzSZlV0WX+7YNJIIw48uQ6vFGmRP9nS/q5IL0ts6J
tznzoy6WoB/9cZHrNUGpxQFm/DYU2JtSd0c9jzYLpp+QOkjKuE0BnVonCjuwWGB0
h9ILmO18AjXGQogSIWOs92Fca1jl6Sgzk2eQG4P4ZZVicG0zKYRsJbLKlqgYp1t4
mztDd+95TpAIeaQZVsk6yyk3PRKCdVklTJ/l2OC7hrqBTSAbDk5xGYK118DANWde
w4W6R90ps3nknW9M1REqM3mz3oPWBz9TC8vz+fc0ZvumdS15JlP+B8lWlCjcAmUu
1IRGvq/xX0T7C6yde4U7LNbkuTD9NplcjESgjI7wHLl+NNDDbuptVUvYwkk9XCMH
zgJpRZsPI6UQ8+S2iiwVPPi5QY0LrSkjVs0jDQF9VaSR0j7j2LZL88+yZe1yQF4t
E+FLB09ePgIFA1EiZKzrWkHLN6EFG3mdnENaoW6cs3l5JcuvkDmpqWErg8HoQBGv
dZjk2fPXSuixBWaYmMooVU3VmG57KM8Yw9tGQrpU72t2JBZhLz+9iAPn5HmsXvsL
zjD0rBWO5SUyynmwgi3k3N+43qgAivO24NQSk9T/SOQfee/kwiNBr2g6/XyNw6/4
ui/0QUvWZOjo7cz2iVu7Srsv0DxOPQWGwD32WIgR2diOg7X4dgVll9Q2lNWzjkjy
RU0SzUE2VRSJk7wRdZbqMY3xEuNhXmpVNx09PEqNYYpA7c+qUW6xK5TnYb3PIlY5
jTNrFaxOAszNQO60kYKFN7W3Tjv7fRFJ9IwMVzHM+c1xvxzIPDWwl0xAJ06Gxe4n
SbaKY1HeOToVY5YBZgGvy+qfunVprxb6seC5uiIqWfvsFgwybVN6lKBZCNqZ8uLP
MRT/KuRIko6wCUZa09m8e5bVRT4smZr+X/9Tb0Mr6IbxbkNnjFEqpv1ynBIIUHOz
vFJUJFYJP70LXnGnMHcBBTiu3JitcwLoj5iYmXlYKks9VIFS9x2jhJvyAhzptzMo
8AKcNLFLeBIHg9NFqxP890cdQtL5qePzo0twcpH+pH/5zhliq3aEP1YQXRMYCXGI
sLj+TVK5wMPpyhVlQYj1jto/AsDCsn1b56v+o0wsAakSdr8REHD0GjXTkonODF2X
h6LE2W+nl8hVdpYdRdZp0yliwH/xUiwFdYlytfZYHh5F45+VsdWBfgRAnUcU8hIm
MSUoh3eY20p/SHsivHJ+Q1m602YE7lsyM1XjEThYdshaeTU7U9sdVw7b2sWUnG6x
BTs95yUmd0/uK+ulqmYdVdPa1qCa/ZAImUae+3Sgpiodj9kwnQAeNqsaQBvNVGRX
gBEOQLLpcTHh9pwQqFOtJWGVZKINQx/tNGOZwi6XVr2FrUfO6iH2RSqJRrDrNjSO
JgtqFz5idlYaFlENybOEzn5lzsdmQHY7eqlIM/3aW5ZlLKE1s000mXNjHH+sjkbc
6bvGtYZUPViQdlPieMeTS/572yN9PpMhh28YWZ0WtBAFGuqjGPBXfvNDX/WzhG7I
vL1wOYO+T0z6KyHMsOl765my/9g3LR9jHtiOIhE5cOYJ2fHnykwpfpMAbpAki6Xj
yuzxN8SrcZC0xZ2nM+dXcWnDnV2EWwyxJ7vwE7ECcj8SjE5wjwDVq7JbfBVXnFWJ
k9wVIijaeei0VB6MW/CkRpqMkTZj7m7kO61hnQmE4v8BfcvuGlfQMN8PmnxvfXAT
+VzFijwau1gD9eFG1d5s/oODMVdHJHGC/56O/COOeMIdMvVJrshZZ4RM7RED5H5y
c1RplfKQ6XuGde2yh3e9qZ6VRn2WBYC3jnofyQwYiHXzqlxaHEQbXljVRDrEEtc/
lAO8trASKGeYsU3wAEgMkFJrFXzNzolnCCbnkz+zoY/WJRXmV6o4M2xJOpDPObuo
h8j0CX1e8CviO6/14Pf7m7k3uaN67U+WIbLuTrH5JZBixqSt7Bl4He5ox0/Zm1on
i01G9Lis3Ry7fLnz7BysjJlHCiB8UcBs63AyIG0fEii5DI5QiBS2kUAASxY1ProY
HGTf6uHYwWByyJ+3YGQMufbIVi4J0s/h9VfUQTqAvN/5gY8tKU4GqLVCvWWX74rj
ODcSeZW2Jw+5u9oqJtvrgfXz95Q2DQlPWlOiczPeczltstvRkeDoDZJVRAaNWEUw
qqsUgP24P8RD5IxMVc9Dzld9Wv+UDX6JAhvYIPg1KBHMGUHNCDdFNdrPquT4SeO9
wJF5O8s0ERgmZnSmkizxYBE2OkYoswlKIjGECguARU5BktfxhBauk7ls48qcfcQA
GaKCEd3T/F1CCxhq4AoI+Ix5DkefwDOXgDaShq8p6OuFg2WVhNDOVJUHrWU021ph
U8DEHcz6sW+9hw7RESeVY5FS+9YnDy3D3oFts967PkdIl7VC+ApLcOUrehlerXkj
C5ye3hUdNpx2W9FsQFWTLjy/05QE9JRNw61QAZMUza6hoNYd+LceR7Ml112Xhx2A
ShE3sIFl8L5wHRh1zyaBnE6UOdjEuwDJ0wwwCqDCpyEFOf9LeCxPJ9lXU0zWf2zB
KoRb6YaLc6xYlREtYQhOipOHYJDKP130meZe6GHLPtIAxHk3XMvd/xjOkr+fykMv
xegjb6FpeCuufnSSDHu/tFhxfePZ0vBvaj4u4dbdmC39r9Ev/i+pWFoCsCbVQYUY
rpgO5NHN/w94JKpR77fh898M23scDEhpRwxHlqBOW7z7IT/1pEqLTnwQCeaKOQ6k
HLBi1Mw1unARneDMXe0e+8QCentTvNWntl6LPyBHaWR40aZACQASenvCC1cDyMgu
zVyImsLcUTgcKm6ciTiKM6Yw5hr3y3I1nKU7839UHWvZLLz8YwANfFtIxJWibAih
k1xNRg8nHXZcIQQ3MX75Fn6w1RknPSE2Tb8Q4cELA0wRZL3f5hX6HYl1pfQsjecx
LkbkaLAB7mpnkPOI0BXuOEoIRCcomplhmKEC3r5f00vM6rhss5QNA3iTe6t94E5Z
fq5fwk53V2G+6fJYCXZlM7goW67lHn/FdBtOL/TNjGzhZcI5rajQ1WQR++LzSk+f
0UXcshsHOtWHv8mIkV+SmjaFlqMGbos1AVad0x4CTd3HEjtCDIpj7qQvCkLr6qR7
X5UHI6xMfEZflFZK8uFkXh6jS2F/JkTAX6ia6LvQIvXJcRlTfKtQ5AoFp9Qbv0fP
K4CDo9o1v93PmFLEJLYs+A5PHY2WfFuyNPK9kmynXUnsV8lC1PCN/8SxkCgve+CU
uo8GAV3pB2KZqwU8qsyaONz7VQd3JxOyIf/gqc8FgsDWJVvEgfEnDsv3Ed4fuCWL
K9ATWLXPzqKhe7JhTlstQVUrqQonE7V+soARw5qoTOzEeKjNAxT8J2KNPjdJv4RT
MZf2UNWXfBQ+owkNZt8LLHKSqr3oHen4WAIEvASMdl+BXswUhuaGCOnvzcP0uz/B
CtxWGfB5j9HTCpf80ZQfcUVFzbr0DUtguvUiKfAWhB+9vk1DHsnQygr5HireYL2i
FprmpWg2x98C0rbDyew/+66tM/2/vEUx7a0ReDf17qCKUXyU/8UOa/Qa6a2yg09s
64Ty+BNHNkzg1/+k+jRLKUVm5dXMNxetY2djcY26WmgFbHyTXNR1FSW20cN9dt2/
wkqMZetWfC5iqEmdYjTUKk+2JrSxmd5uNd3e5nxtLyJSkyOO9ScIst1FDeVmXQmJ
4zTblKGjzDMa+c3sAAG1BTD1JB0tr7v0H7A/LMPnMT1AI5ITBtNKs8+eDwf/9GiK
+Cj4KGtLRYJPNItZlqgEkzHgM+hvNMqSh/YDrm4uqiqqeQHNYxzcULDBsn/Hg78Q
b5UWYWtpUCz5qREurlOLgrcUtWJwshVdMLRI0D5K/4W5FUO+4eLP5egaVDOzWFab
moFB21IEVKt6ToYbSGNmFVse4KXw9EtIAplXdEzzM2i8y+pKRkw3rTj2+zUktJWQ
l6KcZ+uoTXls2ZOYZOj7A9BxE8AI1qTsOfjP+zEktYdxwjqwHXs4dc7Xw5KjpSOz
fsvAJNE/NxcfUIzuN9HZ1FySEuPFEUFWxlpZuJ66cGVtsNjb5ai759IODwSJRhdb
AvF45RTkQrzRWoO3gY/IbIzlDQfclYqWvjjCpLNuifbFrRPw9lX5d18454xdIaq5
Inc5KYHj5VG5GneqSW/XH/s6ZvInEIS6a6n4+nRogwN8+gcgb6nJ/9oPa3sqcQF5
PUHNIquNp9RLHcdUn2nviaBsaTcXc5a8m92s0JLw1ERweX8AIe1mdJczJR8GRLPs
WCVGabQQQXjpQ8aYmUn5LmlYJVrKRaJPaqVHy/E0N7ore1/MCrCJMqFqbRQRJvdP
o/e3t/jUe64lrR8DI2TNsxheaipJaRaGKomdQDzcW9YzXH5JT4tv9BRkUd5lUKdH
3wv8iYLPR0aA21muvIAvkAKFzqxqMno+cN57jopTyfZsRzTfTuYvAcZFpP+7gWgP
6Xq0Gr9RiX8PC7NxGC3NtOWdHvqZCwOiXMGRuKnWInqvmpUisUEz3ohkKT77L4Hk
74eicrE/oAaIJd2AdCn9GD2Wx8rXaTOSD+OViSUKMjmscRtfqtdHx9Ab2Vl6bzVD
clL53L8CDYk3pDA2JljSZYLnd3A1p92OhnF/xpcWnVmaHHvj5PKandFfztD+ynAj
HUainCEIxw+JAQHY16xpcJWBzfKe6BS43M8JGpJwP/MPso3NPEA9OqjEl0o9XvGQ
wcehwqNT5l8IF1JXIzaQQjnP5Xornu7ipLzi3L3NP2IcvI3sPTUhH7U6UCLXpTMC
C1lZQoMlHycZsDES0knKWzgNTnrGttxNkKbSlqAMmd1F1eYZE3uwlKNOi04wiJlx
j0ImmzJuu83GIgycCErWj66m4AdR0eIQ+bzoUhry63BzNPvtb/Q/miPIWBmZKkUn
jbn3k1jD+wYi0iMRgvk7zx+aiWVJrAbzVbVB7wMy1EkmDtydSCFbRe/rM68egpP/
F38vwXEabesF8iHixZXTZGwXbW7qRuBYfff1KYKpQTUpBjkY8uH9QJ5D1ppTIvon
tGSdKAz2TI39JwpwLmnVBAHr6Ep7696o/aCNDDT4mVyg12930LUjAvfYUgR+MEnd
E9tKopwCs7A/5ixnmtk3GPchm+0UGnEjA+6OLU/C/FfLvO1KKrOqOOPkdF72X382
aLlKoJzcHbPVlpqQEEPCZogWEczLPE08lvbPppSC9Yze0kjQMb//htxSBzdnu4E3
0JjHTdZ2Ntx3U3izp99vSrpXQL2SrEAanRAkX+4oZ+uvzFjjXAtSwnmDwq+Y2UmK
US72la5asCShG9RfxgEfMuuj/S7HXPgXWoBGtoARFrGx6TGlYEwzBBiHhEt3p9C9
nVeov2du+RasjqJ33KptbwpeqrCXfsqKXz5yT04zFVz9TfE1Iv+8oxyVeCdHaq5s
xpW6nzU0Gg2uZ5I/N3L2rmb3KwNstCv4pJRoBQuFZ9Q2Sy0Fpo7QmzWfRbUcfFV9
vHLu5dmOiWx/mRuE0UjgQE3kY7YIxq320RteSJHrgX++cOoNIaFAhnNKIutxDXSq
owKoTFuwZUdrkI8irYZ8ETxXJ+akd+Q6b4tB8fm93lEfK+VOcqF6ugB9A9WQWDk+
hm+kY62HstZXWPfFg/tJesI8+fxyYIHDi/Cbj/3Wxyyxl71GMt2At1YbhpDHeTun
knnnQ994GVfKCrqyUhCFRA2vke7cSHZwUxrDcrWqCM380PpIAC+klbwcp8lZ3yWN
G+cXWda22GQFvmue7auQSig/waDuKk5/YSqQgZevAmn4SJILgCvlYVfaMlZaJ/yF
+en9VGAvHCI9ihOUiL0Ch3DzvPHLKz7QBmyscGhCK2Gwp1ynVMyDGppq05r0KGii
yiXO9rggkSqoPZAcTMdgRSV6w14u3z35pYa32sCHMNq/rFEhJTZ+c28aUnS2fiHP
EoZQUOTTX+YIC41E2a2MjtUd/WspxhH/IkYaIs7YmsGz5APb8Wgo16Z8dxJLZeXJ
ffSWOR4ZZsJcCKJaaVwgdEQnZ7TdbPmByQ41teL6bQDy7QWIONWgbUqmMhvYFmnx
qsCk3lheR104eGa1Q5DaeG3sqCnpcrGgFOfRyi3obdU8elqXUwQq09xipRLcU7ev
0VCtApfvaC6bTpz17CYouNpbpJmlTJdAMh6X7F79ZM6Bmnk47WD6+XOpxbcJTz9z
52sPBf/F5EjyxNY2CZn6hjK6Z9jMkK7LOgcoyNbS6ME5k+hKdgsUXIQqL2VyzJvI
Pa9CQHOw+bmCqtrd2koFxlAKw/rhfWv3TEzbelu7Rj05eDGw/quKiO0I0cM8Ch5m
sG8ypg82YOykdalsEvoSXmoanmwBAnfZUSgmFAVKC5mP3LL8OuNTyfAScJjJahhT
nQG7lMTib6BvXERDokUoI5WfPih1JbV2m0jnpkNdFb4iCTvylp/9t49Cy3q44eCQ
MNtp87jUzjzvAv9QOR6KlhZrKGXHwmx5VGjQBbwrE2Ta6dLkF6+ZRgFMgilGWtKC
rdHvu3XQwyOdR3qEQEOYRBC77v2QfFZB7ga799ct8xhBLcbZwBfOxz1i0FidK6KS
0Mw5fC/LjYL9GB83avKLDOvIT+8AJiQ3YoNKu2BMRgcXCz5rHdpaXhBVTMQRbtzq
zZLaDw0zXPQAX3zWl+DKbDnNBMJIdA0OOF7gzr00KMElMh27b5DfETlSbRAWVlwQ
kEp3Thpr2IxUvAIg16CaimOvVjGL+FH6atX5MyQa+GfY1XtTgjvhR8QQq1CmyoUi
b14QawHVLEP9kONuKJg9irlPYvqEMVbPn3rVWRtneSsvsNO/QtnSoYoPHrwnySAy
tZYWL4zo1SdxBJX62gI6Dz9U2u0jGU8AR1uecA6UKHYopGJZ5pk2bjXh8HD2T/48
5DRBCs4oyD1yxhsEBwU8polc4Sh0Z7WhzsQqqc/SDIKAJzzCD+yQuvnIDacMcxSC
QC49aIttNWuZrF30j0brSBIEb6hXPp5wZLxu9X7DVxJBlv8ZzJg8adAsngCGV7AD
hsgj7Q56nxSck9sh6oxOdR5qBk0urUEXV1Lne/3eeYtoSjdBInXEkK/2UVxFSkVZ
rxXoTcM/Sh0khjzs7UNgGE1lhb12AvLwJkOhl1MvWMsqjB0CzTTMjjI0sL2I7np8
qJTRGfnNjWtlWmVbz9ouGHh5XoPqLDD+NBqbmUjNwxoKLAZfYcFw+II6I2iKCOqD
Z/T4jVGr+sWZpE1Oger8R6xCiCSasM0XYTpkq1bCBAewC8sUpsIWc1dkjJi/j+QU
FA10RwzjxYKpjS73q1JBsUfh69ky9aXGDWndYq81HykxkrsNr57/onKNthTGl54W
23Zg31XBKU+JdFhgBRyd40MTI8nsFlLLO3bbQwLbvxoTwEMjKAdvQE/QAb+mStow
EuM8QCTGZoNwWZKPBa3678Us3b7B006MrcKc1fG4cRiAyj6IRr8IRaZssQ24xudt
FkxKXB9o5d1xP71d5vpbnsQR6vezmRv/uReJ/9SPuV10TdxfMmqSYIWFTcg8KdsJ
32ql67ibwFte4pdiTpF51DE2KI4UGnhb7SkNNpG/ECamx/pAb+nStZj/a5HS4GEg
L2ZeWzhgJNwRYk6qGt02i7xc+hGSWt/GkFsJXJ+oEoY8kj7ypABRuJyC2oYGPjhF
4ZxqneTN/i6Mqn2xnjndLvqUyVcfQSswnRnj0A8/VjfkmWOBRWB8/EdSAWvKgabs
nIttJ1SOdfUrurhY67HkIs1V9KgcYxTgXeP49751zkQuRwET1lRNYHiStFPB0BID
El4vsFu91sFcc8KRmo6AfWkT+ZMEJy1W1o2FBmtyB00XmYn5yyiNA9ULQWKbyGzO
F9omqDV77QNbe8fNi9EyA0zs5GwIsaSQkPtgTrGWrItpp8kHB0p0a5WFAZJDLS04
V/wm+v5RMiWOdWjhzAsWBQrEIrY2gGJpI1/MyB44CugAm71IoytgLR+v6SSteoav
G+3oqarGkk4IvoeZjLxVi0F29MmVU/dePEGfP6t0yldj+83XX3ioTaYvpKdlop7U
QZk7iVh6PhPBscKV36JJHj52GOxjpXhWe4ULjyq2baFiiuZi9ChGUHg54XfAYl9N
ln4yokRK6haUtlivBd740wuCsIr8RuJZQJd+WTQSlam7HTOzdOxpP/xkCDJachJf
BJ4Y5sHXix1sPkRnFnAxX60iP0MHRsOgSFPU71FTFMC4RyDOrzdqVDgncEgZJesM
aCNtspPX2wOUD3tN8qLbd9T4hVwIBFTZJxdmjIlFpX5hNXbfnNwRGjwDRZhiQZjO
kG/MM4EfBlCqegB6bMRb5J9LNsI8j5MT4/iPCV7F+GcnB7r8U8eYgTBBTqQ1B7tO
TC93U02Xuw8yYqFb3NS0UZvGrDaZVsYu1uyDz4E8Lq7mUOuYeHMo4Fy3v8ayw+Tg
5be5p+rcKdCsXjF0bbfDkA0AqNP8VXf0FRyboipNcn3BMzaWyx0bsGnWclw7xNTC
FD7BonvnSw9bdj058sHrSElM9IiFS4SiQ3UkHSlDWqcHMaJyr57P8VxsZyNT6SxM
QfKsHUpyUKGt6vvcuGan6a3eNnwg+pGbhByV7rOd6PMvH9tdPBfgt0ZuSbki7Mw9
1Tz4dr50da1tEni/5Flj+Ujj5IO3H37e8yO5borLSs/Mllcf+o6CBCWfdn+ZNQE1
7TB+x6CPQlG2wU2VFDJCNEWE5CM4g5h26Z4tZAYy8pyeALvnDG5btMq6pw2nWhKR
J+IAyQ6q1UeCNyqILfC/v2hEI0bRpNP6uHYS/cxMS41l45k1G5s1haG+L+muze3O
0GTVTou7fGZLiOsJ0OTOMBLtntwxAlLrE8vrVXfQ7qoeaVs43J+2F0lskgXDRZjf
xiTIzdn7aLOBfYuvX0rJWw+aavqa5L1z7Ff9Jao9Abk7vY/y9q1vN37WRm+yQYOQ
1OxITN9omyXEdTo9RGpmcgsyQmA6MZYFbJzRNeXeWpW/nUPCewbimvHbqopKf+kx
wdZ55pJ9wVIHQjZJzAhBcow2mPpmfCd7WpTj1UWjG427D70QOpmaKq9RKu91svp4
ARHYLoc79FiwshS34/uOJSgLD4tqG3dQb2CVqyhP+mD1wt+HEXQMmwe9HYz/vxE2
+v2fpANVOpb1ECzxK2HNeTdvrosW3lJd1j0guwqT14eluxyu/DQ9xFaJUhXyeKJm
vfm672PBRz6lv8XGc6t3LOBInGzDTiHgQ65K5Jh35etfPpSIHJl8/VeJkBrG43io
kGrdtaFlt9JfhBZg7QkCe4SkYl8UJcIiDK7A+CVn4gZkiHwFzwc31TtZpzraGEqe
zigbVJ2eYe3LmdDtI7zGJVnRbJWOUWpcCNE6xSTGR4sI44QuQQsd66dVMwkq0Cg/
45lbXeu5vyEMhBoq9OLhQ52xL/UACy53XTFqOhqT7ASfSidbuGiV7a7N9bnf4hH9
XxtNMLVNT+Fc67O+QvI7zsVoOeYIVIe80vZaj+bRJCwaRbFuzebG0F00ajBvq+QQ
rWxkQg2NXkcbO+kgm6keeUrBhB3kx375rSn7R0bgK/XRqsbEM4JGtFqnJqSaCSFE
IiG6WAQoz75DDnVWGWuGHnVTa4t4ZgwnuGMaFGElzXnDt0G1q5/R7YIcUtIzh5f1
f3Ln7gYXy/oBjCPANG0jA36AVY9fcIi5sjBV5raWRQXVaoFvFbnAivwRA5iiAIwU
4WnD09s1qdcDvOFeK+2QV6z6kAAnnuTS91yVo3pKF5H3FoaeQAVFHnD7ZefVRp68
uN1SgSQKoU2P+c4+A8Hid/G/fzo/JeslWo4En01i7Nsazcs2vrOG4yY/pCyNhjre
w4yc9SO8wWjwfLQhAYFbpinsqIv+asWU/cj+FuoueIXVFw2EMzL0xS7aHUrGAd9n
CD9wq0B+2siqExSxPzIZMjGcFK8jB6HYVuit83w6TX1XpbyfkosNBWMOYpH6/+p+
q5qdfFDat18uhIIJcCWN/T2ESvXI70Viy1WxyTk1U8b0ZBlLoiQK/UTR76Gx9fkl
W5pIrO9k7NJ54nU9t7WqsoO4s8+TucL5NxM9ynBpIQhOXthzFfoiMSoygMJbmfAQ
seP49WyLNpVs6UArpPju51l6oWiPTxuqnjR+yXq6Egsbg4B2+zQCHKZXXZj7MteU
TIVyLDqDHH2kAefy2S+UrqKBSm+A0FcCrm/ar0lzGQe0TGkFD+NIGU91FX8oJefr
ipaZOoptzbdrBaptEqxypMWylE7oFYeMP4Aa1L3upP/CmxK+HDEkVGIBhdPWxxf/
Cipe+7/2SXnx0SIoEOeHsFpmsNsJW0TguvUHPjE5c9e1UVp9ahhIBnyoGzLjRY5r
icwowBU+Wr15ea3ZdrIvCIZgRHejhC7gPq1Sk4gjAGOxAtLIG4Zxr6vJMRKSftQ/
cy4Z3WRSHDZ+ZcABkT/Kjr7g0bGIDIb/yNmhHGdBTjfvA22CXoLnEnt03j/mCiX7
8rVaQsnWL+a79Y21GYCZ6YUQM3YNE6bk0v43SRMnofjQSKBCKwbjfT9xFrFlUdv2
0bujWmxyUa36xUbK0DcFuqh3FfP7aAGEnMMZa7D77IIajKUmw95vg4sc7l9ziuSU
RhhD26I+CNmQgDwtDf1/pkhGgpCWy551qhr4Ru8bHimgN03d/2wfEx9braD5hfgg
PDGP5CVbbjSlPhOU7sgNuidq18JM25R014T9gmVTE4zDEgrUn0iIVBf76KfcQ0do
pVaw9kRrcuOA85eXaw9DH+6XDNI2HwsJEeagWwWOnMxxvBCPrupW9M1/4tHmYnEC
II/uHXeb2YZyb2Pp8snaxS/j0ipJJdfQLuoyIdjQRc94nuRfaHmrF5Tk7bK842JA
2ZRVFCOLX9kYgUeU8y4gIGYBYaGUQC/SJtcd56VlXo0DdHqq+N+lIKmwDD5+QrWv
bbzQGnlbm43ZcFDbzkYb2rZnThj7drzcvzrJBCE3QzAFWIRyvtupXQheAB1UKZuK
yi5YbmGIC7Adv9S8+DmotJMe/fMkn8cwg/Zxhx7KTdgTkcn0JpcEJ5EV3sApEpqT
zTd4b61eb8jqq71qhiHiumIPnbFEL370vmN3gHMwa8rkCqu8VbUFzkrfm32d+YXR
pa6hyjZPhcdk6LqSfsXewsvx+KU/LfvucK/KIGp4Wt3eOictGEVZzylbUQfyDsQT
1RJaF7s9tufuYlYy0/Z1lixK80kl17Jf5ekx4By08Vw7ea7ngz+PxtkeqoLJksjJ
p9EralnptKmmknlpR5FWxtLXtpEPIA0WuSR63Ebb7bYvFTQCBF4+xj2Os/ZAinH2
8LGiDzkYNPHcG73XT6yNoFbpvEpBizhdTcwSazl+e861C+NuhJxBI8z64FYyEzjP
BImOnmZOVf2cBY3JhHSdzTsIoVs+W/jHkOP/tfB6GXn18KPW3XtFqNaHUoaeFCWq
I6djU/n5l51LTlnRdPDVlc9EgkX3LlOwi8MkeIdi+vHjxoI2nThhdt54rDn6uxkG
kaep+iDM/qqeRHXkBD2qc1QoKu+dnj7qcwakPvWrRyrumaM7oEF5hUlk5OiZgQLC
8qO/gwxZ16lk3eo4N4DY0KgmdI73g7kGQGFWCXi5A2AUyqHgX2eXZbMn+mXYLb2b
0yBi2dQ/Ef9nxgvv1xm75NxVEji+maHrafXV+V5z5PoRaBuOUsrokxzNsucIf/on
GlXHeh1BEx+LTmoKta9FVttcx6N6qUbIYp5MJw4TfQRNlYmJdZcvY8pjosIE50+p
OkgtUT3dZwijeoZrEHweqRuyQKrS6n4+3e0FPgIjyzL/57i4ha9co5HQzCoU1/ec
aBGagoqco9FG1SA83djEQd7Fdn0s9ywcyIJBWTS87QBSKyOaHjNRlfcLnfQtTS9Z
frp4AcYdJOn4BwDiWSoOFOjDsZGILpNGIQ3M/med1OEfVQDt+XCHwmwkRUyqYdp8
RXnvNaf0Z47G5eDdFccPLCaL06r5fUuRuapxy9Ailm88HmuC20m9vSw2q2uiKHmZ
x7ql4yeT4iXZUgMMaIpeE2v8gXCA3nP6Tm/0xoPLimwdXAbpLk0FYzQLFxKbsyiD
H/g2S7GqIr9aH0o+ewJ8i7D53WsoK62SkWCk+vwMG6vE3drsmd8eanRF86m+re1j
ZTvooYWRk+kXdhxMpSrLeXEk8XpB/uP4UtQv20OL1LJODUMAuiPFrOC4QwvmQsXi
2PDTgJQYs0msxUIOI8NY+FaNBXVqecK80xStvscbTXlA1gGsFj7VS+ZT5ZZAvgwx
9TIBewiCXDsSuA2FCi9cGJ5y8HwTHAIJeM+WZW53373mbrsV6qwH1LrkUY5RVK11
1AMrcKqkB0rCpcDGwLoMR21sqIjWcAuOSHpkh++yiz9rkSk4QjbMKbShNeYdwizs
KpGgfhrDc9lCyyHowPxxZsWABpsNPzKrY7yc9DUVSL0Dre14qofubnVttV/fLIuE
lfnMTyzZ49gWnwDeBjNF6seL76Wsv0Qtkp8nh4DWnufIHTaw8iDobz47v6FNobVt
v7xh3b/tG/vlrF7VS21vGRIKz2y4SPxwrbsF6wlpJZ4uky7sK4vM/gXfhw2pFiFU
B6jFmYKAAfpSWZ7ajZcbrCry5EhDDHeR4UX6dPEN0LwfKqm7xTHZg46r5Kc5QSGC
myWYv1mxElJ7MU7of9+/LImgeIiTCJezHzh5KSEF8SNX2ysHSn0ulL2bTQsfNpjv
Ih256qFdfsGKTDSNMjZ/7R3UUxjQLchB5YMkh6Q3Y53FPISqppODlYKnPGmi1JEh
OYRTi20Go/xgnc/Uf5F8zRGWTuzLkxJ/VAOhADIvBrYGiY0Izsv1IYnqv3vNlI0a
v3S/dXXsNFD9cK58qbUqknHAiJ1c02G1l9n8ToIDjD25ZjnxiMPPX2L2h1erGNzI
VyuIE/5bYC2LDyw9Yc7RTyhN/9CzbBCPMBau+2r5d3/5CEadqThU48VgJmGX9v1R
bM6re8eVPLGj1ydmV1cMIyHu55tk8QaDt2NBUDbumF91a8dz+DpuCTOM3RLmOBIL
9rEmr5sX02pmROqLAIZ3z+R2Y1p+OA3NMyGY7d2zg1En5GcxpAILHf7hnXxUUv2n
HoSdfwGH2pQ5acrQFXK1ZojPt11Gigpks4rfDLYoT9UkgKB1m4pXTDc2Y7cLDPq1
Q4uLydH6JVxOERWJH17GKbwgC/lVy3Z7l93BOyazb2CbvgPe/v93vW2KcSUvob1o
qtSDytdKba7Nc2sZrHCcoLiigrs5QzazUg010/lrUge3EnICqxiDdXu7MZj3MKaw
lt637sAVKfBuUUa7of+CYOluQRZLji+iRdnUu1wtUYnrE9ym6+YYilmUG2XFG4gM
LQ6pPhPGsx9mxf0xAdRxkxD6Yifq6iJ52CD4fE5gKxTVjcKLufKUv71zjpm1ZqCm
sOFT3F9mvZzKZfJChcDA6xWf9QQgnn/rpk2OsmFr55nDBYgTDUcQBzo7iv0+i5ik
0wHUxLXX8RlZ3Do81HTYxniebAu5mDHx1hAYh2aS1yBPKtzJySOZ1Pnw+5VDnwae
/ExP2pFUQ+YJ0eJZUA7M6rgHOkzR/bXZKAqtaJTOA3xU716sG5DHYihTqUVhBo30
Fw6L3TL3G5mGXRIQ4j31fxjgiXTvE7Qhe94zsR/iDmkobETgCuFJ4gOdMOHmFNE/
INFZFH8LKN7G3RC3//Fbs0g8BQq7vq1EohvZu0ARZLVmi2Agwr0NeJRbuES5vGq6
Xg5RGaG9lZIMw3uVnaagib6e02yD1GucdOA4NmfImz1BPteZZ9IPnXIvq/ku6x58
K1/VsV3jtONVuYsQ3Lf99AP1P08gMKXtAKSVg9X5HZzgA3Lp3OI6oLil8dEtxQQ1
N5lK4wN7gjXlkcBGaVCV6hxC0c/Sahlq5SnpJdpnmspfb3lotyYNQi2KG4/PA4u2
2dUj+49bVDDjBGZuVcOWEinCCCk/LWDc7KO4II0dHi94qvSQ1STUjnPISlh/baFG
nnqkR6ixHuVOHPf/JBQADla3nxN6ZTGXzsZK1nALQKMryXkw2k5O/rtdxJK8r2RC
1TLl9uKfpW1vkovzBfcqKi3YmCqJPztEWuwpKUWgzSRsa1No1ul2OwghF2GRxZV4
Rv4nCUwGS41cVkxkwSyLRPy5BsGIq1B7r0fAW+9wXYgSigXwu3or221hfHcX36PJ
q+bLdOJOCoVlCA8DwEROU6MabHDUpFh/P6Axfl1UyFyhjmQHo1hCq3h1fUczi3aA
Q+F820/hRjM0QmTks4kh2VrY7fTX+4XLfzOK6Ax0eRQBDoJSUMX8E6brrtDsdm0H
kU+ufxqkUXfRDkRKCSz3+O0kOQfdZkEd8VqI6RtBEgQpFW2WKb//qgAJJVjbGrAS
+kQSUb9fs9+eP/IDoDRCdCYT0NVRA/33816Lnvb/acuaTSzoGlgDuVnaE6Ru2cSG
X+3ghAKzlQFtVAZVOazaqzrdM5q/F1+4yHCSFkBgxWss7LKnqS5SjtnAUnbS1pQK
j9W4vBNuADXlR83hT5CwG1c1570t5JoucfFursxd5mogEVwJQpov/4lymcJPSWxk
WQthqKX7CcFZirQFDhfwpdORt8Qjs9Phttr6zl9l0nquJuLoPP4iIHxETwGZQV1S
AfwzSrgGLa2E/kIhcJY9XhwZCC95SeKHd1W2/TtfcocAvv9quKzjAMEMMRM84tQu
8F1snq4BnM3+psiYNJd/Dc8vXBuxz26/tLSkR/eKymXVFS9fVms3MmKqhKValawo
7OQVcZfsU1l/uO91W3UXQVStsvIHgQYvABVRkZw6PmGwEa5KstqEMMield2tJqiP
UXwEOqdefsgg2V58x2nEabaDuE7NvGiS2/QsBfdyr6sMfx+dP/zkjtYwT8fgju52
dhe41yMAm6diB6E1NyIKZ0eXMQfGOjKxN9SYibwkU0fW0VyM2SPSvKCy3eCxDVcW
ilHm2ZINwbI9REfBo9PU9Amk6zGHUiwLsjfiO2pMxIPig0C9qorGPeBwOPFfhaYh
DT83CapU6CRrRdzBxY5BVHdGbJWCAKrGfZY26ZT4fPAXadn38XwT/vZ1hhydaK+v
E5ON4aQ2gOVQzL3UI1HlHDzUVseuF3l5KSjGB44O2xDJsNRoWKX3Qx+gJqKNpe/5
odeZ9WJpYEayPwxhiWlWTa6Z9IaafusTEHXVDTup5OVsoAXoFl5JtcBCt5sm0hZ3
Haa0Wl6NpqKrq11v4fXNvZoSXzoqWaR8yyEFVgBLdpVEidVpPJQXOEwPDenlc3/e
RrGBsfxBfKbX9xNBQQh9H5NLWO5SdjehseDJw4RxDKOLvHHMPsBnm79jfFCXYnZF
twEvLkN1HkTiyC1618F7ojdiNBurHGVw/V94j/hGXerozn4M/cGUUwL/51nx4mLQ
LZPVcU0iVvPFyHgyOKYFtI423/flSl1M+QroMTIsPbLRKqNvcXgnHLfY3uzporY7
EXBmoklsNDEGPAVJMY+eXUJAjHuNyo1mqsWVvlNzWQLQswcc007I7H9xfrE2VTd2
szzFQua7IU7InY4q/Z0qVj9EVMuBBJHON0+83obZzjIkwSedmn4nX5dgkgZGfzHa
J0GP9rkeysT9ocfAkUFVIn1D7eegsIsVENh3Y2cYDvVKsd/waluu3vcNoBwDumUR
OFf+c814RXWomnd1vdytp3Bwtc9aqBlSB87WzKjw/t2m1G1JvhzFsvusPtRECwYE
W4MkCYuHm6kww/a789H38la8+cGnSjnabo+tCL4gwEE7/LoB3LbcTpaOTLNJWzw4
xYrqOhvNznnXxK7Q0QNwcU0KsEaLWCZGXyU0Y+mNlW8vd8cG/cp7vZX5PlP/+TNw
MG12KT9vJZcRITmaKlMv+r91LxjyXshv1UZrCjrOlzWIJB+YFrXqyyivUrgSxVIT
GdJojS+nDCSohXeN6bmzvL3tViBcUc8zh4wktWn+1ee2stxbO8T0ixBd93/d/zwg
UPFWmURwJ240O3HjiePiSOt7IkbQ3DfRpoCqxEmhhAxZGvKrokjzzbCdjBygWebq
715pWh3dRCd3YxrQ9MmqRyoWxgOPXuGrb2dLM9GcwEsSFqMI/c5+9Gs3Jb2IV9v4
4hDPfjMioVl8pLbLyG/PYR7YdDrTh8MrDaHT3jy1dsBoNgM7YLE1HLxms0FMuO4o
HL8kt+IUEf4RROJ//NdaHx2mYyz/S1O+WkuDKKKnw71vMQ0wwOdHnvY20a6vBjpc
qT/BzwICLSzrCog+uawpZ99DB7RZIABCjTUJM1XJtXVwh5lSP3dpBQjAwj/ZGtcn
zGNqxjm7pteMWsY1maUYWWvhd5SKg6geDb8tdJKYrlNPfD88kBXD4PglAeYCWoYA
+C2Zcj+Ntey5RG9W2idoO1ni4YqGMXwV5iS+0VMhn3x5gMIZImvhJl6U+8C8YUbT
/NNYWoyT0iZjOMRI5qENkUi43o5zK0vHEumrIqM0rNI9UCLAM8DiZC8QQBSW2mvq
c3SqkT6U3Kcwlf4CEm9s+xE/UIpNABqpZQh5iDPhLMa7PByWeygavagG0Gvt3crD
6bytDjss/I1hnMIpEuS/CXRiHn8WUloRIF5sFM9mVPYb+PX7bMy274TIvlggQMfN
tTgnt90QcBO+roS3XM7CkkEoG5iuKcnVGi9DnblCecLE6u3bvADxYM2/h8vA2A5j
CeUOQwUx2QezHl4zZK0pjw==
`pragma protect end_protected    
  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
V9PNqntu3j04gmTGkM4IZx5suMlb7+HywVdLe3u/F7Slici7oxoZbqS1OGRfMHWA
X5Xd+Xtyxkfo0m1/gXsyTgTKaaVIbxXeMPTPZPyaQx+DUwQYIeOUpLKOIrbnRRVO
2mCnU62ZNNuU9FHgvEPQS4bt4xBVDVeNH5vwbXiFUHM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 30051     )
iMERZQLgWu84bke7zqkcrMQ1CeF53Ar1ANaY01IUATyoVTYB4YjvgXPUMJLa06Tz
A2VaGOSwgUhHLdTw8n/9BC68hDM2W5S63JBelJJYw0RCrUo0jy+iAA4O86Q2iLuL
vaA6Bco1L6uFK2Kf/a8lj71fW3a3l5iXTlHEhn6EYGOEaSu5R+ZJC6RkIXpsfKrC
RBEPf1ecK5DzN+E1pJ4CJg67TW5kmbidQGGfl716htGtoCRT2opeqzIj/8cc3+RC
AXrQMte0hO6jGcTGFvr4kqowsxl192VTBj0q5ew/qj2NCKgNfO0k9bEHPXzfv1sj
agXiqr0G4j2yvERLd6nQKepH0sCJNiF3MVhMuWJ5z9OWmwZK26Kp9bIGFnun6Uhv
W5mnu93tMkvvhmZFbUNOKWeL8q09eU6O31/fUNkfGwHKlmcRdNnML4+sv+SviJ2j
nKvJg4O4ULz6rLU6Q3hDjokZtCP1WttsAoTb3gfZC/NdVZEohEzdbyriyhiuz4rN
rIg2Sd38l9OHCQWKg7Z4RyxsF/IzfXR4SvcGnjWpyS62/B1KseNV0+M9j0VzqXpr
Nc+ZXTcdwrC1uGHp9N2xWKLjrauSlBgQ2+lqZca94Wgx+T1u6NciZ9ed+iVqp/M2
NHbFuo1zIRMLe1O/syoNddb/ympLk9Q1GdXJ+IdIfEONuwEkw/fAVhvKuzSzVv55
SvaLzb0kWXX9OhZQcJXqHuU3TQIOGk/ENv+4LtaGOZanpk5C+oZi4bFmeobMBGcr
dJ4O7flNmfopY4uSOUtygzXTEOtRG+GkfSvyF5U8WK/PMMRL9EA5QJDQI7hYsHIu
XABsltpmqBUheXszEW4GrNlK62A8+XC4SjdhaAJs5WXWWNYkFEmrg1ZZQd269Ymc
LZ4zHcKvkQuEha+0gKQRMWGhykNt/SENB/xGDOkPNakNzJR3d7B1JZDz5VNqf+j+
MGELtRopuzj9Znc4enmjru/JhJoO+0HCCf9491JFv7r65R4bhVAa80mWygQM/ABl
T61I+r9gAxRPmdFPQX46ck7AJAFg7xn6bD08AIseQUgJ7gKy4WvLOMfmgeRwH5t6
ETyKUNSrNN+jNLmBtpBxwbHPtRUyFMMC+xPvLRY4v/cmFlmHhz3Do7FoUFmKTblU
rdxj5Ypta3AvNFGPcTwYJC6Tzy9k9s18zE5F7r+WOOcKE0wyzILnDltWVbwoGAim
3k4y0yDV6NC+7VqmEXPp0HHSROGcpkCnvBl9fHO2S479O2mmL+P/E9sEIrccDg0U
fY5Ust0k5OvIlyW2/DrK1N6gi/HYHi4adDfmxVBD3qRPmEhYRmKDaIeVmCbh/bxb
fV6mbSltJNpCrG9RpQG04vnGECfBXSBswCeYpVxNFl57nAnGB0n1wr2II3U+50cC
3dQ9kX9OrMuIha7e3u0J6Kr/v7ACcWPuRV1DPlFRhWNswEGhk3kpwc+pj3yS6XzV
5Q1PabN+RikJysZ1U5VCnqeBHi7vciKsZclH7VFkW3r6h7Vp3LSMUlWS/V++FqLR
ptn+AhuOAk3Sl35jKPSOYAHnzx/jdrv2ez43/hwqaTmUOmaOYx811REpZIclETip
l77WjVJHSLVs0GqxrHNjYVywO91QziOtvUq+1tyV0apuIOx1vGJltXpRWS0KXJMA
xx+WOnH3Jx7Ybq/oEMALIqtRJFDoPmLrNA2QycxbvEeTCpBGkAIOIl+TLe0UDKzf
KT3mh87I/wq7KkC9AfQYDVO9BtBZYk9YAAMR+ngpCB/Y9nOQ9c4O7a5/78RwiBnN
WD5rsjNLn2VG0yG+gkllpHIslq/4iL/iYB6u2BhbeSQb9zXEiAdQDyrH3xUPpYT7
kZ1uMMOslKOrR6ILt4nNmpmx9jWNSYhXZTKqlVYPnExElMq4d4aXZtERgZvYY7dd
P8bRFjFWF3Pw52s++GxTsNvjJpTevPeFRIl+LVqw7FYXiQzkOxzc2LEUN983EolQ
esro6a9ZXOZ4ObfMSc9B9vGWGJQMiWOSkG/lEOZXQKmcsRkJFgzjaxmBoCU9/LZw
o2EvkVG3xb3cJE1scATQkAbENyG1x2HqUDVdCY8c7hYdhP6FxrIZF2z4Gryt02Mv
DDOkmlRpxUBhMnI/x2ScLElPfdsxVlH14SzoK4A4fzDCHygfX3glVR42eznzolvW
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ovazDWHVWM5Gyn40yxsQDA+5DrAwg5eYxj7EURtqEhQm+pU5WjQ+ZlA/KLvbag2h
bLqVpP4xQaL6bF4IbvAGiS8i0DqrUrO3uDbebYvkQbp7/KQKFOFz6o0Wvf6rhPNQ
mmk3ebXQTtxiOlDHpJ9RCzMDVHjPGLVb1NF2WlosFpg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33313     )
usJWVSgNheqe1CsNzTl1DTtsRO7CQc7P4oKBVSiwgodvwF/0Yh0/bhLZhmp92czz
ySZcsq1rOKCjd9wbQ286GGskOiwkqnDNFTm+HeLdDYf9Jsnpq5HgHS1VsFdrkqB7
EYUy+Dq6mcEe6fWrY8vbS2n/ntAYeEAxCbwnxQYhtEgsUfA/iJsWfyivVq9pIhLC
9y2ic576U191qfrb6QkpYBQZMC7EGgr0PNiJni0f1Hu0a62KGGtyW0VmWHbpFC/+
gUc14cOZsiXaJlqXJOR5lgV4JxHbJXuioEwv6ESZZxzHZH4RKKgtUdBEhXigQMe2
66jQdluolnwQwtS2u4nvDWT/rt4Gf6FU8D2kp5ufsY2Liin67Cen3EndxNM4mXNs
2WaCD/aaxdi34j4UdfdFaBkAaajAUCs7pGV3epnBGqajr5SIyvuuG808hCTISWCY
R6+9w68xv1T4d8n7f3WotDCDFWYbit2ImbSVEjYLfMSjt6XxPOUOuSOZu/AyOsWM
A+mjDoYzA+HOU3vQ9j4QsvP+D707NJU3jTYT9aFjveSrxHopYbkgs+KOy9Ge9VK/
Sv6aV/+k+5alkpQUwQcnXh7BIFrd1+jeYB0Or+H/8i1UGK12bt9JcXoe42KH2FIs
gwk7FQAH96dapB4ATsjCiWx0bab/rLvAgBOTKKD0vOv6Ugdgh4jF4PGNZAnmI+6A
B40tGoJkELbdavTDAyt+5DEbeIgdd7r2PcjXJWqTcTWdInyLgFlrf/jEv0t5JuJE
ce2foQ8KaXu3v1xVKqq4AuUBF9m2kaAHCyxMlItL1jDapucIyAOHHGHlLHEvmCh6
gemqmY5rRuyOhKtMu7kbg4STTrvQNZ0LC1yNyG9nWS3pQj0z33caV+2e1+o7Z8T1
1FMSMmybC2eVLdzRYSvJpHmSDpnKIfsdVsQJ6Bkia2V4N0A0N8xi0TPoJBR+ixFs
BHDbMuvfVukA1ZH++2RWsfclRaIZNbsldzWwVYhAqkh6DNBKajKN5qHxOeV/WFpL
ScESgH9AyBwY5pPUkIu2JrtfqyLEgq9M78ycIL6u5tABpLx6toDDfwOG9A2CwDRr
4w69DYAIl0UhzrqQdgSYOfH0m+1uo9hIthpojrzcjp1LWLb42/UGdlVH4oNiFMEK
hGYoXqKaPQmqlQm6gBlxVplp9JPx3wNaKSbwT4xSqqqkOk+LVno9fxlbvtNWBRTz
6MjRcvIkldBkHuBKK1DGk3NT1DoHCGMWpPjOIa2U91EdMMF2yqxgg5Khh+KYoMx2
oAs0uvUj4rWujPsS7A36p/hRClMVdZSKXUUQ9TurA2hiDqq+CHrm7ZuXxWGdXAg+
hom7c/ydvyPXjo9mdx3AvPZ1+FINXY+X75jOV5S8SxjR2yngUG3Xzl15POGGJvrV
E1UKcjm6Y7UI4SQ4twtaPyECUOLMcU5BX8dJ8IY6jvOuSWnIaajE6mF+1Ws0NRHV
x7vMSFwzCmRHzabivNWIIhSljd4L0W3fdunnDN5yETYi94YRer+7wmEBaM/eaXf1
OqdghyowikbNB+pkHTaR+2GNpu3DshklpaPO2GJ9d1k12WEGOyPP0j5QtdnQQIF0
CBykg0tO2mdUhsfJY+jBEYBYckg5A1iMoDz5kxcQYa4Ja/4r5Q3DzqU33OsClKN7
uFPC0X+sYMX+0OasRh2SZdtnCVXMbJulr5s79xnBET5Th2oV0Lk4HdY4SxhOwCCX
tTJMkQJ+9qLcWn8tu6dUrHyWS6Pb4HbGwRdpHifA9K6DpNjlnN5WhuQ5NqsJmiNQ
IgxbdMBmbFlPk6hF4hO1NZmypo6g4+3qpqoyYstTmgZO5Dm7pAEzG17oOnR0ZmJO
kk8WpS9vl2akyeTb/AYz/YXV65Yv1Aq0sdbg5nQUS7o813/zqoauUlECVoDQjV3e
Pcyr5tFebFi6/Kx/mREK6Ul2yZTW1ydZnFCIIln4Cv2d8ztSIwGTLuXhU30jjNGX
RXLcGYPbfXx2CZvxNkikt2jApcTiSzgHP2/tNrcD1zicrwROWjA0Wz+p5bsrrFwr
ljYkQpufcAmEQrw+gbDqurWEBehtrJE4kIoNFFBFsbtntuRLOlkDgNXsUAtiVTZz
WDCu2xYbWrtHpFjAtSKFyhz+G5CgMOIQwv4FhXUg5NqE8FCL4Q17NZU8SXPX+pxq
zptc2NXC9sJgPqT8x+gicjsQ/hf27hmoSRJydABEAr0X/e4FpSFVTI7Fr5nGrtNd
YoSApWh2fXQYkzjH23FBWQvH1IgzEHz+zxjTlAvK4HRvgE0ypC+MbKsFobi0pGtE
SQkHn2V4e3GJZbZbyYv7/4/f3H+ot910EuKAxq3tSqV0+HdXF1ZdGWBK3ZaN31qL
o9YpMQ6f7Nn10cjhWY49hTfxcQwtApZqn8ce8Fd9QA5YcAi5SZhnZ/F+akEoUV2l
8CG6YWc2tQOCdwy4Y05WvENiUHzT71NRF9nLSrfnzW8UD/CZ4ffiTv+ENbAZutWi
XNFNGaXZoaMaaPfbFERj7kjT15KF92VUdkfOFEAfJUop21abr+ByUG3YAA4+m2Ir
CDgE2YTOPyrLqRFyrJAwdTQAIxUXXgqhiTNzlEWnR2DfvLn++pQBIIplLbe+RgS6
I6SMEClbRQUIH7luM8mgyBPoGnYQxq8Li0E3M9heqZ8YKF8bByaMlJ/f9tptmFXD
qgoZId/QIdfPUHSMKrguW9gTVsXfMiY/Zf79H+aiO73QaKpdfAKJYLjt1SbU05Qf
VhIbtSwRcqy9QqTn+xReJPggZI/EsQsn546G1+sWuFNjk/LEnu/R6rts7XnY0gTW
IoIF63l5qT0GwqTa3pov87L2ahWBesB0fbb5LK8WUyo3ubJaUyRp44PbrfapVaUG
CkJfnwfqUomPsvTA8Qv9TWY30/FgVeVjcjetjMd553tmyK4HXIqMwp1KdRaTFCqB
FIrVLCOiOnVz0j/oZFOp/5PH0RyBl79vyOI0bETsKoEzC6SjCOONBSoD9oqlnN52
zxuUfv9+si1H9/qPQp6ERIC+QetomBhtUjma3ReneEk9sqWCBqMv7Mz42AiEjoAb
SGM3Qa7aPfDyxsHaHcr+nfUHdn3WExDaqNsmqWeqIQ5iMWlkpGhnxTtp1SJWmW0H
hQ7Giakf0cLXhrSUGkltJUolxMENecdLxqVuHTeBZ3FZ5SFb81Korc76c0s4+DSv
gwGxID2JVnX9uB0TIzcOlbzrv43VCcqIzB7e9DYh/AMFgI/A+PW4iQ5FCD92h9iM
nQH+uq7DH7NVN6EKDMOJNjjOKmq2riDKuqw814hgJsraxMDAIV+Xpyklzlmhj15A
54Qo1G03OV5V0njHczOCMWPm/n7P4krZ4erxkXhP3HX695EQ1T090NAYM4Q5dgl0
0qshoXMlJCU7hsKKDxayfuqSy0f/+jRTi1PV+YJ1NspuLmJyFZyEQtKGh3aPcrFu
lSJyhmkGxt2kYKISW17corIKNfb6KNna5Mgdq8SfLVfNqA2gXwwnG+JM93NOuJBQ
7NwCr2zFOsecly621EBCENDtmcDi+kSKFduSw+Xv9D/Prs+jOqf4cEfNE5ioL228
RaoTfymNV5QhORi5LISnpAikgNs0shtl+ynNrAsyK/7vADV9baCdWh1SyrnV4qkf
tOG05IObI/s9JyWvoA3/Tf46RIexhq3IEIEwBg0ImWk1BPS3V1AIbkM2NrgpewCy
fXy2M4anUYS8Nj9p0LNdpyyls3SU6GUv7qE5U9wSv6s0iyr5MXD9AE5kk9YQhdZa
9r2BML8jeHhp91gRzq/xC+UJSyW0atUVdi03V5S8LO0Nz+7mkxHnHPNDxJ9cDtFw
SnuLf+P3R/V74GaXx3HiOBDBDK3xhUeabdypia7GXV658sKmGJFtF8iDABwh4/9g
jQxRh5ePAhELxKjyn140kfr1t03czKIxnVHr5MUKXw1W9CibnOyKoTXI6zGTYXyx
eazw49K1swL+HWU9Z+gMVRmiJcpy9DW6eJDLs9JOEv+h85p5PtoQKYzA6fzfhjsh
PAWIRyRh/eExJE6E5nnuZbw/X2H2g1UZm/hVsCDnrFRDI4wOvkcAfweK80j7NxOg
wIT9TsEKlmVauMFkmGVuXqFX3aD4sEMYaV/SElHZ92aXwwxmhmKR/XcmWCaxeQhD
dmRoTuzNQPW78l/A+t+JGutvIXa7LcfF+IJ6ocftv/NEx0ypjY8kLRM5dr7p7K3P
w24ttKySQMixjzYx5pHI1MEPNjWPb4kafxlJ0VnqahK37nxXSHgLnQdwK78UKZTz
JwB+Ru6ksHHQf2x77GYH7zk0tCvlAIM63u1hcGAuVAcDc+kfzEGvmWnBG1lZc/yp
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RYwoy9bVrrTA6eam1QvWvJA81MG/k4ubIyXlni/JuyNQ0Gzif5+RW6+lk+iO1Gx1
mr4rNqjbA0KDcjv9AcIfYLI9qiVc3LWDQvx7J8Ede4QwLj1Vngkne5E1594vJ8XW
uXmh11xc0AuaqkK+c4ODZGZVdqE5vdE1VbC24BqEaUs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 33472     )
3vE4bOF3sVxC+08oN2VVdtnvpexFkS8H5sL+vqBPmNr+btZMcN7+Hb3ryY3qiuEP
I7HWq8OvBukX8mff9mET8QvUnY1foicxye8ul77AvFYzRBQV35159kh0AUfKdfss
abL1z9zBUGO6gxS6fFK2HxfxD755ehx7ONDgjRnDSPI7aTq5la5m1GFFmS7oKw9g
vOT0CBMUZrVzB8C9BOMEiA==
`pragma protect end_protected        
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
QAnu6wd/KFj0stZm0apBJjljNX6c/iupBbAmp5NtStxaitAaDxbuuiXozE2EveSN
YaolF2kEt1+P9PNeK8ICQqr4jcdr88eS32V2b1nfVK4+q/82Nn5MHztSX51dsh4T
b5KN1lRHwA60ULVFamYgBs5wHYtgL+/wKX4UR8dlDRM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 95053     )
fkM3qLCq18ODEDozgRc5tatbO9snuhHbzpa0t+krjADBXn5B8Ins/IVo1AfFPmXK
1j7n/ASJdqw46ZkwG/tZgMSRxjY1D7H3dWUoZ33yzUF12Rw/NMfHcK87qac8s0k2
q9+Gdyl4KYIb0z1bDiwHCDxXTSL9oAN6V+GNqGG3/YXVWSmFEzSFawzc5vupRzp9
yqwCquOHouw6QMyvAYMXWGfbx/506YKoetvHYuxrA26zpGwL5zNUtItm17h1l0pl
hHFG/H5WwqonA8GlXWROeD3wlvTMDJKfWJGG83vietRpSi03OdzLcVeh3fhVFigA
4jZ6b9FGmzguwX5JOIhYStGAv9reXkmHU3akKNUGk6pziw3Y/L7Kg4K48nQ9hwrQ
92FQjH5QyKu/JKVEwkaaBq3VusqkWNgZTr8ExlA/gntjJNaxiS2rDiLpD3aZXvkr
eLqPG4QBFR1QrDRa0ZuOZcK7bmFTiBi/ssGfp3y7J/rNiy8LlGP1f/NkwzzshZq2
0pfpEVHARBUEeIsaj/hj1g1ldLCj+y4pf6obwMqj3/1+jXobH1Q2f4EIIrHfsXC0
Nr12pV+5vzAiB8xOYitsbQZDUQwF/v2Wb+7l84M4wYgVTAXxgAXefbZ908E1qpPk
5dIId+9invqWkwP6ffviI4yNa6DAIzUXZLxvxTA25jLAkms48cOSA0W28+k/GNhc
WP9i37jF7Fo0rXzalkpHNAcwy8KLYTRrG9S/MZ7oLusZy24zArHTARGKuNZlxP9e
cCXh9DOKJFcRAt13jFoYfNEjAEQgctP0c378UGw9n9fbHHEO3HUqeKHB9aNiwave
T1lvBMvNOBrUEGUAaUUZThATCetQz0ACDiQxvlfOnlmytjp1DAbHPIrKmC94KZgh
d0mhjoeT40Wj98/1u26vh8dheolXjpuDGJSnrCNO5cN5gpwg+wEPA/XenvUbI+lw
wx7IHv5ptT4UqrV/UYBgK3SietdHgmR+e8psvYy2+2YDM8f+ueD4N6jFv5d6c2Eg
WoCtJFGZ7unRKCuHIJojJnf77IZ+Ya8r/oH67nfZWjZmeUshkwyyLus9CNjT4GZC
ze6ME5/0t8b19OnxH9NJTDhdXzVDQDFpvx3+NTn774zQLM4L138LquqScNHndONS
XhnR174bqX8G89JJOGeGNouitShr4C3UZ+4FgxJ2ENumqucbFoNPMn3nv1T02ZMh
M5PzPLKuudaFdxOGxDlB0C8kYKmedbn2HF3OqYMN0BWviR3HpzxTQI/4Apqddz2u
4axzBPiOcX/In/HxCmRUas5/1kximM3op5IagS3m99jNHGnzo5yFAnBDKbQ5f307
Dq43EiPEk4XKNJow4pJWc6SNKHQdqsX1LQIXku7nswEUJDpmof5pdi2h2ttIX1k4
IvwiKITuMLaOaSiF/swgXqmm/ufDYv8Cgt4sh1tIO8IUTPNmuVTdqHAcIg9xq1eB
iQJHjBGlw0VnOGlWZeAXSp4E3QjSQpJl2iObHfDHw7ZX0UUsQF9JXUFzPLooozP9
sBo+OmCugyn74rc2sffJAQnuGgE4K4OEEXfJue9CnkvnqrEgDI/t9p73nrPzVyEl
GjXQj+kcRh8L0nUZxquxGAMXA05k3oMy4XQA4e0/FKfvcRDfP+ZhdUgTJZszJLhL
Z3pzpg8lui8AtWjvSZsmetmvCMgIg3OcHhCCcq6fcjdI7FQ5NvmscrujzlJzcf5P
tVcLbNXkNibmnTkwu4DQFjqwO4LUGAXxVZW0fM+S+lPkgw+WGSl506xMPKhaHc0p
bab3xVIPEFGWCwZN40MHjqMYQHaUVfai3YSaSXlHPNEpdQJptIIS5OzO08lFvrg9
cJ7A5/CXeQuYSRX8zWmNWCzN5+NB/i3DhVs+lbaQvVV31rHvD/rMwWWY6zqSv0Wg
2DgIpLFKvV4+LuzoyElrwwJo0Nduvf3Mf4BJeshYzPkTmG6m6LMWQGbUEXS4lUAE
SbujfjLzUxWZnA5mby6pJkUiX/aDuCLnzRrvLJQa7ZQE7VdmBC5ctA4MGUA5Weoo
sHW7AbVPiiuP4+qV7VBwucAVECgeOG2Sw5wDz3V4LdhFgCu/kWfEKubr4zBncn5A
REyJs6TBjVAjVlmxVEjPRK4RHuRQurJ3suuyZLsbVUeeL9P9kDt1B1y73hC59Kkd
WM/j3tc/cas39yXO2RF54azl5LzrQlB/c4Yam05ZW7fMEB/a2wNciLDGmC23h4xf
5G0h+isZKJ725lNtt9iVkLCWbne2yE23hQYnke6dkrV3OqHWeDTLoyitsJc+U6qG
j+KheOhTfJUYCXwpMNxO8FDjBoxqpiQWLyY6OnazYea4hIvtmKG73ZzShtaT1zr2
I3Jj1oBUQYsPco9v/NiVIwG3jGezM3/OshcSiatKfyubDLdGLh5ZvyD4iztf2ydF
sJUVLY3SzSWmM9DOF0I0SF6K05TcDwaqSWO48ALgX36mha6mSSmV31J9UrhiKsyX
yJDmwGKvgdiZ8Yy5gpHFijOm6aqYsS3sQ+pwIWeEyGsojK/XuimY8LVX54LCFso5
+QeNqE1BOCEEabNOZ16UUCQK0PeKgZU8xGPYUElk3ue65BrWJldLON0DdTgTkzFo
ZRRKblPW8ModFww7u4zLxC3FWXnPqu90iFY36rFI2Ux2H0MgFNCqKwHbOUVngVUr
ofvzvPPGAOtEwBE+YAwXyIlxXIgk8rRt9CkUnegQLXd7KYZeQ6lKO5MBweH+gL+A
TzgYs4/iXiKviFvdYd/3SioNnQUgRwm4slX8E9XE5digc46ZFRac/bxckA5UshRU
iYU7CsgmvHTO7/sIPLz/xWTjnSsG/B6YLeTvB6ZihvIycsFtTrrWaWKdbZB1l4JE
yuWc8enPradCHlSGfvKoMTuGS0reLrM+qN0ARo4VsWqFFe62Rx59sVbeB1LKV/kB
gFbZfkhT6duw21LjalVWhpBjnonzsFK3+HrL5iBitabAn4IVaX2lX5JmKlMEZsdu
p0Rmdo2EpJF4t/rdre7zQGa/YczjOJ/ut1iP0ByxIQdoGZz1qHb11xa7ETr/Aths
Cr7pn/21wYfoE0Id18dABvyvg+JqUpUDL47GJMWDPNK8gE7teHObbZfSfC8ziJna
S+5NGfJ7yUiviIHZ+SHsuxQmQVUDzh6E6tRyVhi66q43j6HUbAr4QITFCrFoBIJ4
SFf57g8tNGaMPGgm1REvRYvXlK2N44wClyS1BLfRSXSeEJhWJ50yYxYxSSzkEaED
e5zY2r5NAymT3JYljVTULexbN4pQn6aYBt4HMxqSDy7gmSpZHpjxSEyz5TZ1L3NC
YDvIQyECV2fbww10adXEe/+eKb/ONyCSjE38dcLJqM4FHpldu6GUAwvMMrLzquAv
eNJuGCpLF/jynfaP3MyQcMIhLQitbrz7tbk6gRJx7+ubbQjdhYTKvAlA/otBm8Nu
yZtl2XOaE4IWBYtAlAoy0635CKjLKbPJapLMLBSGHqX+t2iG7U7AKb5Ulv7UNfSi
rNAY/6+zGeKpBPD/xtIi/6J0PpnxcRQyRE2uZXVkpetVqevOPWdbo+Pgz8sE7pKq
i1qF9gTePPyG6lpewZEL71bQvOIuckZzGsW2Mu9GeLJsa3+lPzzpK3HU8BQKN56v
xV9qSqrShkgGNCSxGtPTVD3wXAoCY8rVl0UV7lXHulkrEl1LOYAnD1/uLpA/a3tr
S3/mBdjnhSlIyKMLAS+ViYilN11spSHLouxrMamtvFz5n/c2qM04hChOsftAJld3
72NOgTXBY2agbOp02ZfqF6vDVg1ZneU+B89BCNZK3LAxLfnN49xYgykk2tUaRcr8
bSX657VJQ3JgN3ttiiiK1vE5cy3ql490DUbsX9IUMGLQ4Xc7NwIwGEKhCqIqYNyA
yTQI1I7DVlFcKYD3TNJVGBeCu9kAY7pfA2KI4a6HQvmw2+LHmQV1IzAPxb3w9kes
vFOYWo64qEHTA6SThoy0oIeG6bxp+VgudxeAxbn6mf7u1RrJJQK/PBV48jC1PLBq
ZHQiRvDWkNCHIAD1Mq8ksxA7hpZ6GNY4/1eP8zV4xkIKEuUdoy45vbS2YB+jBTVu
wReSnOB6fis90zHpn9GUBSJcJd2DFzcLVEA3cAilb4RQYec0ze1yar+0zekcZfka
Pq9K1TdcFxFy8VSxwVSwnsmbKihGaFhO+SS962Z5QBHo0MQl4NtHI4fWISI+rPE7
oiZFZyz5unQFYvzajam+0Hris+8qrRzxJUorZ6DLIFOAABzlqrSNrM55XHlaN22o
PYnrH2vj7DOwo7WmtJn9rRh/MRKynj03MTzBnA3HA2VRaQQhJPeckFg64KbUtFdp
CRBA/opo4Uwsv6aB/KCuMTBAQbmcmZKu4AlZtzgM/pl3ADb9WhNwCXOC1N2Doa9D
fpOe2heG4Nril+c/9IlS6RBBSRYqSRy8H+UURFya/CcqHXuTmA+ruTKeL+E/1TQA
UrErjZLciOBQ2xYNoCxEhynqcJSzS2xbXBpcFgyxybp1LKxDNCvubiay+Q1Kr4iP
OCT27KDynisIK6nC8Ijwi9U+HfauYGEUuL1nWcQjRUzvOJ7GpikSGyHlCmpzmUi3
SnkRHqOKZro6V1fhm16TBS/QK6Jn9oMw8m7O/3XlW6nASdIg9yVxNZ2ZjfEfMzf/
qfkGxulT35vgYtVq8XgyCzspF4IGlLuN1LVW0A/Qnp7TGP/4PDVsCuE5Ymnsga7y
cinaTyNmYgrFCmhX95FZr40i6z9rCKD7SKEJ7SPxUNHNl0h9dYDLQvgEBUDGOFEl
R5m3vQO47esHo5KQmBz23Z0j+xHWDM9KjHj+RuOylhDjEczKdcgHilEUJLdW4qyM
97PC44Gl2pKGM6yVV4+XKxhvfTXtIQZa5Hh1P2R21r4IRecTKvMub9g66vw43QDF
w/uKpALXKkDYcEzR7ihetI5oh74yi63/my3JDg94VKwDkL3FgvV/A23YZqaUKdbZ
JcLEdRWJ8O0Z0GhcvJjfia252e2ueKirqXLtakUrlq/Ae/Y31KtRTfRDMv3tAHEC
ioQDZLfJNK6/Qy7QFB96TZ+GSwwekNc828RRUewEt6TAVyfKn8dp9kz0hAKTIAX+
cpmPZYh1VDsGbXI25//udI7AU6PmnY/57Z19OKzjwTboxeD36zaUcoi/614ipgcG
GmYzhwWHOd6ghmKPXdfJAGB6dZniCq9lPP60TevgXXhVXMJ29bJw8gKs+Cnmxtzx
Vzkl9iBS98R1jEsOrrMG6kK+otYc3BXSDO2O20uPUXkpAvMyXBCwCftG/Jz9ID/Y
sDYjsBvvNdqZI8P7uNbp7Oke3YFaFM28PIW30h9WTBgBL3Sblg7o4wen2WaGZjzI
l4cUkG7xCtmePDNBkf0vxFkwa0PIgobn33ePBwJtdzRANeh54gmLTuHeQ/g9Qulh
yuQFTSLS5bQRXUp3bGfaoUrN1Ciuaz7uckQEKJfKsCta9UN8rEyo4r/C5uC9dDmc
Qr8BMFvluOuQzloTo4KCXimogOit/qM8cjXr4arL+pshmQlthEIODqYPCz41odpk
JV95UgxiqfUCvfRAAzB3HsKd6lNraBv7cF+HQT1iyFVf4z8AS0b4O1GxkAX91qX7
dwpLdUxwulrJwXpyx3V79aiwRtGxPIg0v7qTKT5Av5LQXn55miVAEd6HQcl+CepD
oBO/20qPcvF9w+6DW/4MY2ciV0miK9o5leGNuVKPSN2e3gmja4dFRm3HHVKFPypl
PDQwV+7fJM2+M4utoujJUqDgvg4gqrZvDN8FYzOO4FY8ZWeZwSDMD6XkPkRaRd3m
t3qiV2dXD/ZB5dJGDYjZ+Sp61H6RSjzDgsrFpxPuUYh7JWlh+Qn1/vMO6E36oSRZ
M8FEg7g0FBYpmSBabUmMnVf9e3Wkzxnk6bSvHeizTWq3zDZ+fvgblUrIFTcx7U2Q
zeio2VpCY87ZZuJOOEs6UbQjc2dNr/bxdbTpSYv0EzYVF8HixXP+O+8Tyf3O5GNQ
sTsCZNmOXvNnmzgmxNOVA9eN62Phce6PcZVmRv3E9lM6kgHFT0+v3IFeO+oOF+7A
uo0rICiHz1BxAD7I15Gd/1P+CN9OEu0zyhw8gOJix8rIQI7U0Gc59NJGBMYOy+iX
WN1mIOv/4qAfMVD7vT/LP1cdP65za/VU8hTgLTsY66OFCxNl7lA0w5Dg5HTm5/Rb
udCAGO4hqHGGIj++JdFxSVH2LNQZ6r0wJpdoNzOo7iPMN4tEt/hXXdp+r/6ogcJX
PdI3Ho+9wGUjav4qtFHdkq3lK/diwIA9g/3Tvw8FRH09w3DZXEgvaOp44j+TVmcC
olSP8Cwma8jerXFw3/ANufotZPfMwD8i5hbfiuFqEuuoQ3IBhnO7+WRiG5ZnaHUY
4ohdYMxhaKMfq8KLGhx7qu2nWSrGQ4kGrKdeLVbDtI+/eJ88GkcqdlLoXgUbXlnj
zsGz76ylm8TsqUADmUP/bTEMREdOjZ1eR9S2DvXn4t4G0KChuU7ERnLh0LPuGusm
V/5S1Z/OLfd39Q7ZfEVMpEYhBKmBPtzF4Qfz7DJvzDh9Co9SarDCoEP/BxJfOKnh
szdpaBS1kjS6DsRVlgoP3KG7yEq5xjN8eDNimbkdbBye0MWtMQXOBcPrb1RCntUX
rkIAJcgol2JdK/9rXFgkEadpYoY7XAm8kVAoc5gHKSnXRhu9/17oMZQTJlbg0Uac
VVnLRSC2Sf8IFS/qIJA1fE4IqiNfEEICBYrDWjqMTlRu/mKL+6WmVC2fCLCMZlCj
sD+sK3+dK/CeaIhNZER+i9U3QlATwN/nadwwUDEAe9D+WbgE3gNTGNmgcm/UXp+e
rgG0tMTAKkgPnTDdliVg3QIFhhPZZHBwaFPOEmJ/OD6OrZyqfe7vMePfqn2CyyGL
ENAg4V5ccDriL2sWg46TXiqZcJhTYAKPEtw1KsGDN70RWy/Vpp6Ms19UNTRNQ9PT
UXFVUTIF36YAn3lME9hH3t3r/yBhIx87Q4dZAM/6NJPvS2pREzWdeRvlSPjx8qI1
AJm2T27srPpb3y+XWk5rYqlnTqW6bSOAbLdCMFkti9DnEY3htEWw77w9KW96+fzq
G8o/k9poAOon1xffZESRpbr6VTlkLfuN81Nr6SwyME5WI0Oog6YXzdOb8lbgWltI
uYNcvPpsPhyt0Q3dZKDQpwoEW7wNmVJT1mNN/GF+Yle8D19c8RsJf8YvP5VFfZzX
mNWxTh6b2zwlLRghhFev0a4asYQlw2uI4r+e+D+hiTGrIVtP9mE/6aLahEbMRPAl
w85sNI+9n3XVTgu0kSNQjdp/syPQWut1OrPoXPE0UShnLitQraQmhtU8djs1l8fZ
Kv7+i7Mp8C69//vG/k7Nun8bCon/XWOJ5vpW2dGuVYR2hVGdlaLBcVuq647o849n
LaA1lolZHirZbKTYL/4tboJPFpQl4XGhtZDdZfwNpfa+MvfSy2ncUa8EsKlDKJ0N
ncv1+vclzjXFNmx+WG8PdCaDzyxYFzSiNq3uBODw8mCqyuP6BOCKTyEYn7Ht5pp3
1GNhZVRmZnmkdXlOzY1ZmvD1lTrlmsm27GGM8waGBIG0qK0GGwis3p/mMYtwZTRS
bKu6jXcsDsvD4521ePJXxJ7FV5AyfEnrKZtFkVAdG3IPiR6tDCnON+n4YBqv9jR6
o3SFUo7GAKBcefSHAL+Up+g47MHSenhPurg4q5vAHzOduKrJ5ETC//c8tSiZMfmG
arNI7FRtvQR2LJHKo40rWNCdcG2XfGXKiVvsPsgDel6ssNStAO5lXGbJf98pBjPT
cREACUtURACm9RN6Hgw0995h+HwdzCbQwQUyIhvOdAXWDkvAaKG2BmvxkAmUqPwq
9Y29BSRPkbWc0wdDi4N9YunlgUlVSWEEt4tKee0HmO50GdR4vpLvEQZ+iQZwzjc0
Vr+0VvEDqC5sSs9gjgMCngQRsFnXuI8/ItjPUCOBPCbfIwCPOcUjp21G0pvttwNv
ZY3abhPnWiPDMm7lguvZqZRv4t2UkEj2HyVfqgm8m2OkFkOZjYucKihEGCnVjrbH
HWa8SxBqI++U7Ti8skqbHHkQvFc2VuhSuGsPvwKXW78zcfZg70qSQExWGtSaamir
AYNf/m32xYYqzfZuR/r7eE3/B07lrUJUvuCoQHdKWnNncL428NvV1vt3GeDST5x7
4yBjy0jSR3VFDyPjmHIeGDWU9wQHzS8OyVNsHtwDh5/uSXSokhQIz4X+YcX12a18
+xd7ImgK+LLteip0I62CrHkjvBs7kpRSmOUTtDr/1hI6u9LBNxSBIGt05IQ7LOjH
4ettV1WCECSIRJLkNzd+rjyxMPF0vmRhNXE9Qiyk1eSzCfQHWbLaLkUncziQYVtf
HfXrGbdoCyIf0YInYjQoD1nUZTDCnbcjU+KSwusjkaybFUrOnrf1pNXRsZ+nikWq
onIoXqWTd0n1S1kQedK6q9DFLWTxWYj8XEfpVRvJoGJ1n/RawpSbicqumS543Iji
AJcJFD/7sGt9kMUGlYblITXxWJ5P5ucj5M0bll492G/f2h1xiBpbPTbHwiQrh6AR
radLP8b+LVg8+RlNvcmrlDzDOO9rdYkm79gKQ+Xe5ClkW8dBzDDEbygbFJ56Jw5u
5gwWGa7ayJ4C2dpQUzTiYF2OYNZpDXVBLr+SvP6vO5aTfu3RMs19dMZ58kWnuC5X
NCJh/YtY8bmEyop+xO/9KpDGCGWu6jjrQAz/V4mS3iaS1sWJcD93/SLpMBYqncZp
gCglP2QnLbU5sSGVDyYw/JooUJ11BoRDludDUlLYzt+ve03rsmV8TR1RS59WYb2R
kxswY0Z5SFDgB7jpS6Sb9JA8gVBcjfGSXJdzGrWGDuhhlsdtYNBPVVu6GmpgItPO
ZRuS6RW6teT2Tc3hlQPyQB8tx1F0gRq9NktxpdMB3BtO1lifaHCzGp4LUngrkUIg
ahiYWqiAMJK98iriZ46brsCIbmVndhUEguUxOCYqPOrgA8ZX0upnr617qDAiPx1L
Naqv1NHGxeKppcd/3VsWGoCRCxn8Y1AJGraPZX0GID3rwwVF0Szb34/UQGE9eeJS
xVTPUAaqs1dC6SBHvPNhuTxevH3BwviC6bj8Fu3fiK2Eaqa0Gw6eB5qASPxDzIsg
3Fi/0vfehISlwlX4I0JB+HnBDT1JAazbhIY8egktS9G0zGYgFlrAUYUYCTcGvDc6
Ueaea/+R4s5lhnf+2a7ArMDwKHLXbk5B/B9TkAnEreuUXT5Nf2QRXaZcxAgbnemO
Cqiti7dVLmi/y60JHtALcfsq4Wrl6moUMJOAhKFpZE2KvRlv+g8vfwB4o61veysT
jJKsfgzo9poAdM6YpmAtXt+gCLeVsqUoRkNEUgJNOztiC66SK+InsalyPBG24qPQ
iO6rKhR+9maxUP1NVdCpRbzsiLU0HGKOWd1ydkciz22Plg4k17N9wyk0Nt3O8FX3
DiUqsGkVWaxl0eS1x6aUx0Hgy2PsOinbsS2RyP0WQcp2TLGTL6KCWb4LeZGhRN6K
tDK8LdP5NopTEIsD/H1KePylaaEPYvBHQ49eAZMGTwLT+S66GL2j8uqhd4jldlZ1
JN3aSnLZ9vnrCQK9qF5vawM/MzdFN2yY8zLy0ha1kCl/9pjzeMiiLNTlVWKHlayI
6w5JVIxnd+4vOOCEWQ85XWVT99PT+3Kqxs9bNwxP5f0Ov72ZTY5T06M3mEIyM1rV
A0GUraPqy/UBPzoE6x/ZAOmyFibNGzuOT1fqBJhgWf9x7+LulWvETij0+aNxEsLs
SbxJp591qyRLLzfQLQvsNVUWEBYVAQtsZZVb+fTQGARxvvMDN6SexI5b19PnnAPI
PEDgzhd/bsJgARh9pRBYNDhkjEOKKWefD5fQIfZxq73D790LPXQC2IyogdXGU4Zg
HS8cvWmz6f1j7zS/o8bqZFPDr4yjZ2JTvL7u8n05S/hM3lRPRvrccnTu72swyn1V
BjFyRg6s1Sad1aeoWMiXDs/d97Ax1YVDmb5WiUutXrvtwclDQl1W1IO0MWjhAnAS
iZMT6jLMGWOToEF1Sa8Pwjt0swWtfmOmf2SWbXHmR9fPJ3EwLxFCLa58gixjkpkP
UYHFT14cICons7YnZhVlk67mW/EcBIcIPkaWu0n81PwFe5qWRnhYIkJZbjK1FIrS
osePvTOkA0rYoZyEhnU5jtKAODUgSf4FgvdG8KDox+LXApqFaoiW5h7WLoVpQ9Yt
wSPwoDxPSCsSd6FUzaYDcvuwKEC0XiVgGjIUtGiEbCtXodTrJCUIjtqIDZBbLznP
BWkH7g8EsyiP4sHj+dkTBj8K9i5a1NTQmKHJkNuUTDhrEno33pYR4++yO/1Reu4c
jC0/MG8wy6rt4lThupoy5NNMpA0peCIP8ok5tqtLM5ZohHDVugPeeS5/p9DfX1/N
5Q/GsO5yLzSt0aLmDZBF36yUUrXnUkIHCBBzU1dNon+X18weGqwt/VDw7NJcbyFu
fNTkNX476XVJW9tI90hubNiFaOIMHAVMF2YzHDtMZlX0D3YV76/3ZHXVdKDV+uEP
eBtPNYV1B6q4/Pz2IGdouBmAjLU1nnirsqB1zHNiJHOh+FYXyjEFyX+clg5Pa+8N
cmK0ncoL0s0qEY44SBRmJvy0ODLhjm3rklOhlSXe8LkXtDqiQPobB0tVLJ5qWodO
1v4ShRAnRE4UVwiyawhJJVgf+DOUxk0ofNczx0+iDUX00nJEos7Ay2ACvmlNELyI
tbu1GDlBVQA6Yb3PRe66puxYDt8Nra8yuLkiyflabRjntqByvp+jinb3AIqgtlsV
rOiNL9XaXMiJ6mhrhiBBuraOmJo6j2jPeLIah9vz3Qp4/Hb0nECIO0jds2uLd0wX
KJoTGHTtHoWh6iiZkK2EmJJSGeyaGil+NTMyAqDPt5E++TYVk/t4ahcENb42rPi2
2szOJYAYHPNx/kY5FwLyuaQZ9X1rxb0csUvmnJe8icdLg57pZ3zTEfSic57s7HDs
xsraCHr0l1FwPBsw+QcpbtYCMS6irHbP5raHBQlgDbc+sctntQQC6so93YVu7KrH
2mYS2DwtwJFDxNd+IZcr1xAZ5hqTBUQlDqKHNe6WWLL6AR0vax+XOBQTZvoFG3R5
Ebsef9umK4u3SXfKwy5mGTV6el/3LQ6remTnU4NpVgn3GVnS250rZzpxhj3O6lwn
sdWUATv1huIAhbGcwtciiaBBWgoMDfT181TI0IlsCVkgNoRu6SkDYYzm7xZ54DHw
qZCkzCMQxe7npFX7njEE//kmNnUdKpiArTY5J1FpdWVam95nxsqltAb0i4TJU1EI
b8vBwY18NB25C1MJReuIEQVjqlZLQq4wKs3Muki9KELNf12khVQ5a31g6Qs9+N+6
o0n/JokEeJvn39szzgr7rwqlUhJM4J/n41C2eX+TEy5DZlxFFRwrVzCuJYdxZXvD
FrUN/ho9gV+98kWJlQPClAVjqxrzq/DKmW8MPglKTf4kHwSCKfS0xIJTcyhb4I0L
lR9grBcV1V1L8R92YOUcW2aFWBjWVBhFjxTK2iCQkO1pJyziwU/Uhrf+q6TPkaTZ
UT5gZ2UKpH/4U7F2SfeC+hG8mxOnt25hLxnyi4Ln+SxWkm1wYv+rReWktN2imTIf
3BmvW5hfIdhwGWCZ4ggfqt6zXBxHpLO8tVd0PMz7R1OvSpwqXGprd5wJZRRwLebD
rPgHbnJ3k4YxhuuoroBzRuJnp2NaGuTS3FIhLDVOGrcuScnDvy9cgNh8kTxuxPxS
Xii0V33U17kns8M43fYAIRNvyhlA1BxtGzUcTkh6nbzhKhTULg6ehG4MTDUc/yvp
Fm9d5ieIs118WRq6e5H5347C/7rQJs1K3X8BCYYG79PAw6tZWGy2Qto0rQpx/6bH
z+Xnu1k/GqBQCQHy9H3CztZ0PHHqVHccq2QYuC/oGcAZGwXhxCq75m8/18VWgd9g
lRF/dmVBVmM458RM5xwEcHVFVo5Px3jqbzlK+HfTXrMKZ9tWOeIezRsDMQbUiT+v
E354cdz1ETJp0SqlycHmObUhraTxHoCb+Rft3mxt+DMNWlxbb2HK73bZ0GUKH4ej
tnRg4VmUuNwKVws2Yb+joSEcHpPwm6jZm7x8LJ0laKbyjhe1aw7KeDGYb8JAVTkj
guwhNB8Vq8jbT8zIzLNciNg1ckZ2rXIrvLaR1IseVc+uLhEhJPFWi2/iWwyLHHQL
nITHQ9y4suk8AXW8Eswk1hzkUTnXleVw80ek5o0qbrnRDChZ7ufSgPv0zWjqDYFY
t8umOR9GIWSvignrkhU1484CF3XbM+zylAJ3JmSq+KhQ0kGhbwRnu1mHVNqXBJw9
ApInSrCNbtHaMvq8gWntHNk0bdPFdjMc4VejEgwLFLqJ+iqXf0PpUVXD6wSdiveD
vfu5X+3xStHukeXxwrMsO15CJmj/ogdtsIKmuHHQxJ59TLSsGfpNI49Zj+wDoisA
EMTMM9NfAS0X+OXK/DF44J5cveb8qtJlsVH5Oequwh498p2vIqhNouzQjhFUl+1N
Gg85jwSob1cA0QxyZtrvxhy4aLo+4ral8mc5UTAiCblSEnZeNjf5KkduauH7IeUD
d1VwmtdEq6VehpEgAfwvUKh6mEQN5LJbYW7BXmeh9+wCogFDbqNsV5fIYPP3X8lq
V95Zq7pD+69Qq7UBwc05CpWUIuU1az/Nv5azXHiGs8F2q8q5XguXY2CUMuXSJnfm
86tiy4kQnFalFCvdY5qAmfDK2E0hxPSLEkpKSL/cI/Jfk4DVhc/1pPbdTUb7pvcy
OFkkq6P5XPnM4nON+287ZO/ct6ZDpTTAgrVOCDNNkN2m1xkIdOGA6LY/sg5bKk65
d8nKethMK0XsWFr8DjiZfvkHhmNrQkBJu2YARizoL17i8lNFTzBrNzxuImnDitL9
kuR5AT/UX5pTQG1oVbqah+D/EqCuljrN7rQqDfNyXDoiCaYj5hX/gZRICLEC0siU
hLyK1rfJPRd1Z8NBYqXVfpo4tCqo+EZLi5Afu6K1V7DJyvp1OgnJGXrZ4a1KeZ+N
x8YILK2TBT3fd1R70gQvFtYNdGd5lX7oJTReu/ACH83eJox5lbN0T+hwfNnN+e63
goRebC1bRRhAsproqdsl7uoq2T4yIASE6h/5GW2eZTJQoXyb95x25KGX+mkaHokW
S/WgyFR86GYnFbJSIW3hjkmwKCbdsGMB0XuS/AePR5WVRYlaIXJIWaDvXe9cd1rb
DuM9sg3wsHoRlsjUXJ0MIYs44+sbPOw2T6NlUgP/nYjs2ZQz88VqLyYq+kh004if
L1tiKK3xJErwtKTvdvIajFRp0ifIcyr2uNvwk/IFh19W6buUKZYpCfI/wLyauNWK
jsiroY7uY4pErsJbJsLjwkCO4L6u07sEPnOvoLRvlHtOhTwNGxMxixVjI6zX0kqR
U6JkRc8dXkzd0Dt56Z63R2h3sueJrtMbpuGw/5auyLyBPWYTtAqlk1R4GgQxPTBZ
DjSZ8aSgLAeWA4kFzrlqf3dlPAUZS5vuxFbRddIgSyLXa+DY0tCSwxzbyaE+fLrT
dHRf1bQyTA1pkwRQqiSY4/U4plcW3j3ck5MnzQfIo0+ZyRk+HScDauim9ktogxwa
FFPzvv8D/27QRV+Bp4pSo8romIY6g1h+lhGlQ63q4E9vPBn7lTA4RVALySGPPDMU
pxAPu+muVkO+RkOYYH+8PL/ZfE9377C5gvcvQXMu6LGDdoC0MKOBIRyqfzWhblKh
EMfhPnQLuD8FbHh8j2gzccvRlYauyEDVW0XPbncBDl7uiF1xTWhjHn4BFKGkUqvj
ft86aNgC5Lh23w3Ja60lNn2aCJbI8eM/61GAQJKjvj71E51CBcJn8G01lb0M/PUZ
hcjDtikBzO1Yk81/FUQpEPBFg6qXTOYb32J8+9ZioXmkGtXiKGrDRxAG0SfIaARI
9eHfHmWLRpW/4Aodiu/rJhcVc5BPQxJrp92dWl0+rcUOuyJJ1f0pBNaIXi8HFnO2
npepWzlTek5hS0OuFxLE2nzbNsICanycY9lKYOVK1GQDKGBOr2j5DAK1g1VX6na/
1XMaPSIC8E/5ZayuRtaIQRH0ePLR1eUUChDuzG7OjmDx3VXKYQK9c9TtqCPiRsuw
eh/fGYqdZ9eiewPiMESO9D6ja65AleJCZhLz0BlZ1T3ylRjTRqbl8VKXFTxTPMsr
d8Xwi/1ckBeghpfeVQsXfS3p3Ul/UnUJtT9Dtmp5oIsXnB1T3Oot7ZXa8Mja1CSQ
nL1Mq/Cy5uea2+b39VCA51VvuEb+DlfDxHB8uxF+kJfn6qBy+E5PxjP6P5EfFjE9
uYmrdI6E0HG2S54fg40sKfqVvTasamBrkaDQH8r7gy2YT/Wa7ZB27OISobrpmSCr
cwAoR3Rd8Ce7TEj/ptmElZaK+qEhH7rDuQs8hWGpbdyib+bFitPCGuTa7L8FKQFz
pMAlkMhrPV6AmKBeK2MspfLstG6UBH1035TLIX/sOxrmDXfniPQRLeazBWl/6I3A
fAnnhViwvDTdQ1TTvxCN9nr0wO17q066CX8z64CuF9515bsatycxElJL4O7cdScm
2K0Itaw/yyHs81+hN3VqtO8ZZaWJAQ2dI/2+9Hxfy3YFzagpSQj2h2eVw/x87skl
tZ5S4kn/tW5qv5MHWfXi8kCcPQ5dJt+XKUCurJE/Y8bz/uXj1zfW/QSbyQEQlL41
ok0iugB1jX/n4pVuakbk3bgZKaHXY7bTFlowxUHAEspBHIZnk+4JBhQYNILcPFC/
IROaoR7KYjWZbzFTON8MPqGJO42ycQB3deUwRwom4/pZYIuj3kyQwwI/VGfnrKFf
iAySAw4De4HCd+z4xJaFDufXV0sEXYXYMXpT+LRVxOPLT3BMqBP07vrXj/dieqiM
6fIcu5wVsfEsxpTUSQFA37JnzuonHSK/e8KhT0uMlsnlnQ4VoWQMl6HgbSIO+i07
fn3LQJDxQOFxO9NyUeUtR94w6zkT4np/DsgadKNE+3Nmc6PyOYrXoUOlOFLr0Kvg
PIDiULJhP3WEde8TtfjVqj4nJIZqlDMIs/YPu1mJ86qBQwhhybmmkiCOzKi00oe9
11Oxj1ANSVXHv1UCMywoeCOYckI/psPb0xFsbZc7c74bgXf1NzWlcljVzucoeFE0
j/ZXh5q08Rj8IosmFqouDPsiiUB3xgbRmyAVHSpUht2i4C+Y3VlM3uOHQVlYxwFo
u7sQFm0Ol8x2MQUj9Z4v8N92LC5sXLs51lcuyup9+mGn7LpuCBb/OUTE70dkKHll
nbMia4EX+nZOc1UxuBMAM9Yy8niLljO6okc/l0NOoxKJVJsVCvo24JN+aMBqzjYY
dIw5sTQ2k1VC5LmDzCF9J/YmuMgiwuWhzARvpzx/RQfE2iK17MlTIcIIM+PVJiei
Dg4UyCqB96sgAuyC47/u+q0L/+SSRqEuNLQ4yJIfuTAwb7p/KTcSWbMr0W30BJgy
u8xPw8sr+kCxAgmGEg9zHdKR0+ZKhmS/dWRq52l9ZaHwiqrfW6F2UmhudW61zYO7
7kaPxY9huhIn8Kfu0CmARkzwVF6DfabT7yR4d13tdG6eXkGOlrOy8fGH4C/aJ87O
ctVzZ6s35VVDTz4RNXGktJ2F7jqB33A+CgqRj6HGFA1oNNEoGtN8xQd5lgwX8jKI
XIpvRgykbftAZxedsuXIrALwqwFGuCvZHTtv55ZNb/ZbjM7RBebJ2xgXRFmvZVal
TL3+sObgBh5pZ+wJM4j5BjXyeU4fPoyqN1IwtSDqY4CxCc0YJ3grnMKCWP9Nt5F+
RR1060JfPyFREajlIMS6Oa8Vi8MM0pVTEq7q4m5rFab6D2Qc/7LfDv4WkHzYIxA1
32E26rzzf/V0ioqa38G+YImXSmH6SNObGJlco9Oynvj21jMExyv7OAAgc1/JVu2e
5UvCfMmbZUDjdDkaHdONuNB+91ZGD257mIbwecepk2WqaOtz3tTTyOW88mLP0csr
Xw5mlV79OSghQ2CvPamCpZZBsatz9vb3bO3vYguJCiSXZFC2GmkfFSPmXKfsSbXq
pffsqdvPiqJEZMGDmpondwmb3uiVlwHP8iQ5w14km9JvAHwPFUYPEY2mYIuRmpO1
9HiwY9+9qxc0KAntqaNZ+XIpYFmwTPuxrSw5oPJxfxSDxkm0/W84xJllsfevS+ba
Pv/8jbNIEc6GO1M8+GePWLrbSbi/MXv7Yn1u+hQ4Pvq1WWFjnRw4dYuJM5UgKtPZ
zxBuVyG1myWLnqv/YUfxijecG5/szMMeIjfuzaGfOCBlLJ+hZ4pD9/ZSR5tT3wGk
4msuP4wEPTRYp7n7RMCj0qwnNEYd1ElXV8gF5N0/gbj7HyfuK33mcZ2XtOPqtBos
dKXBc2GFm0JO2MmP5c3qOC1f20svnMld4Myj0YnnK3js2XpiDssxpKmj2aDHLeSK
t1ISuQ3sPJCwQQmx3FFSjymX4iQ9hbemBIvi60P7NPffLszMLCetUgPSuzO4In13
3RDU8Y4z7QkM6ka9/3tFrhOlNuE918qEo+YHVZAaiNy+kpobyAcLQbLQf1pBqm60
iXahV0C8FRUz30GGO9hzL/oFcevTFVjhnOl4B0ANZF8cWSUAnBzc5jO/zSv7RnSa
LK4ei8Rw/TQYYSZPaQShkFMASqzJlQT2lQlOi1hxla1eW8buSNyASlEwkpWE619M
otXqNixoxtRiPvD3Px6OFloAuY8PvTVNSYQvCMX9T5A+rSEIvn9jGtU5L8Eicmie
7evueKQzW3itp7LTmIbkVwBQGBfJ6Mi05c4qDmY87L8MvqY4aF06iXKEPON3I7ky
jJDNPjV//IoaSg1pIOg6/rQH0X8NIsTsY/rCa0i5N5szCiGWiftNTOVh0d1PSm9r
0lhaXvVBvf6Whek8U4JRERS7Fq9o9FTWboTFhtosCiMA3DMWYDELcRpM48KfpToH
2sh3TEZGNDUP9lFYOFZkdEYPdDkhr5S2a3/3Wm50tADMpkEWvMQRxYawGWVwRMz6
X5RVe9dhrMm4or0TLevfPkTv6DlFDVCDpbDExpLhmEkTwafZs1irL6LvEFQkEDOU
GY7zQcdVleHcFeHJBm1iXfK13wZccvkNkkhXOf6paqTLrCp8O6Hqc8aZJrGbqweY
GgoORZKhS3laAu4ng1FVR4TtrCtAuEQ5pM4HFlpRwUOZw4mgXxbCg8fEsL8oD4Vl
gw01tFRgQ23vxYCbKJLP0bAH0ChlJW34i8RriLtjzh0qwY0z+Y7bo4hCNeVndXQJ
jxr/F8K7rOKadm2+nQ+h4tmtYsxzHZCLKH7vfHib6ob10bBJcp15PTVj4uJiIr+i
Y+GiO22foKUfUDbqRfklM1Ta+AKnPNc9wjuHaL8zLq20Bwl31Qse4DPbplah2MNo
JAJjhTKFvlLhgzAAJ3JMdy3VdzK30LbbtddMY78GiRMmj/PaviCISoavvqaTHFRi
dgwOn1JPnAxPIaW/VrM2cKDaW9buJRG0OCcT+B2HQlrsaQSFE207PdqoATiEEM8L
zgSpaXvg3fbqn56M/Su390vXB5AUN56OMVv5a9I0qltcn7koz0TQQ3oaEDe9RfDB
w2mt6RCadpSxCfabuKvaadyDJoT+7+ATFtPbtNjN0Q8AnlSr17LuSLjaEwM8mnnw
cwrceo1NW1Nkyww+1f+FPRz4dse1GrRaw2TKBOrA391YX5yVkwCgIfMY4YtiD4pd
J9fcUq1Duyw+ioS0URQOfC11cZcqO1w10j1S9Sk+RNUS8w/vsEyLjrMj98FCAJ0G
8ZIpQ/WWCGGIz5UmJXDyxVkXBSRMj1XUwmDGwUb/Fxm7s9mo7lAlTmua8Dub9TYF
+Dx2oXyMV7jnkbLWHMGoGaVWODaO+yoChs4TGTfKHs8KDPGWgWtL/v1XNCUBIvWf
/zxLYOFxfhjDbDSnG4HAyvdNxI+d48hCwdr5O5UfpvGMGO/kDHS1gQW/CuPxVIP4
t3sxfdF8pA15PHvxwxMxgv8hp3gMAPXFh2Roq6o+Eek87/XpYeM7Lr3ssKPNz6qB
nC0IBfvyY7JkmHgzp2+nsGvE0qI5LJYEpXRsB77nikvc7CtA09uQnb+XP+x8BhFt
CDxPxt5OJqLGcjCgYvZC+0ano7aXxWNMgz/PzWGWuUaDAzdLr2YpAfsOWGQ5l5/g
8K80OK5H5lDodn1R9pO4Dk2CpYjsvz0B/8NYvFt3v5LoeM4D3NXTuEDtk5fNJp9F
hwC4sZvTX9KwlHsh7UySLHfVWlhnuJQXQRs1bTvpuczQ2Gh77JCPgyJQL/MDC8IV
ZyqtvdPjDZkDpiKZN80Hy8LlU3ek8QsuU5aHy2CqGCgcM7c2bOg/uvNXuPCA8jyO
F172Pneo9AgETXG9QTSwwel00T2e1LAKw1mfbPNGQMDhHVb9Zb1nRxryDhXm5sVI
yiL23h42u/yC/Qk88P9EAPErijhxFCwvZ2nfZfO3cvrHoKZY8ZqxBSscPn7Dligo
pZkdlKk63eQ2FnlidDh3B0mBH3iKPwGGiK4ZT3nHQc2jifn0KNZPYrjKP7S/tHmU
drhTl+LuWrOwVbVgsvsJh6FWoNzcWpD0SNZ6Xb0v5DAKggFl3pvMSwgrEoTrBrl4
1FHhU5JXfi71W2iBBEtbPrcsdNBszg/dmM23GU36HvjIPrgQkXP2IkqC3WLiuIhK
kX0XHYg6L2is9rkhfMHEb9lX8pqLnT3SzrflS0Bbrv2xHlIvBg5eH4Gl3Y4ouO4H
/DW8aFeMFB6XuGKJDU+pKEWSX7wZgBmM5ABWGzjfVIYCnZfX6lS0UfdPOX1Xex+Z
plccP0ayhmhpA/VT8gforsdSJZT/6hluokLIzn+aOq4Fasy5vxw0Zc/ZqhsXIIP0
+FRVjaBkQPfdswpJyKOY6LHfGlHVk98ymeU9y5Ab4EvCNQ3ExpoU9IcPq83/biU1
A3s0UrGzCkpOJm4LnMGVfaONTDZa5JsNNpszFjKo1SrZabCMl19rPviRQ31EfUxm
xosTxMme27+w26BIxIrA4oHVgroFN6GJXswwTrfwkXwl98OmTp5ysw05qc/p+7ib
Q8UgGDW9EKifE9ogOvGMw8oHPSo19gGRKL6WOIxvEwWAYbZ8lyV7hABFZBAc9QIs
qL1AuOeWbTmBFfnnZUUnhdSwOdy/XnU1VC/4wuBKQWQssxCCv5ZvcoKMclft40CF
0owaSjOYgUXLTQLzKi7il1uVjofnttOZ1HEy1sVUxFB63ynxxXEoombFWcu8WbAr
Wxf8h4R/JSTOXr9Y4aQn6WL891oS2P4GwT7ZDSgKE606Z6NGk3lD9WJvn1uQR7GP
74mSmuHnms3aQaRT+rA44CEDN6O3FSz2CXs4sQpGZR7C4Azav/mDBDNyrpYaxZc2
XW77gWzCfIP6r3qxURVuBiM8m3M+lR824/qpd0Khdx7Qo7B359P/kKO+6XJLrUfg
IAW8KvXIBddpZRGOOSrz8tZY1Zy93luM3f45nLXiWGJmKMfweOEBOZEVxcMrOv7r
qY7FiKVc1g93aVnxZIiOEbjvjYc0fudSLjhehou6oT2KDQKRzKFkdxapIWxHoVQU
mm60Vo1A7rNz6b3lkBISYIYcJeXXUO6JBqPvGAnyAnEbvQvXJs0/zndzyiGhrJ1S
FtaFTaArThUAegW2epy17be0WVfz/4dJ2ODY/r3gPDk4WqZFhA4eQ7E4AbAg9k7d
HdPfBVP+Ga9vgKHqKv2QBG3XIGqiCN/OZC+APT01y6y0ngkOSsKdH9hAl3084tTq
R6jRcBm68lDLjc7ZGTXBaMxY5Yb7tV6Yf4GAuIIIdj9UbJpMrQzK5PvBE4Y4BFfH
cYw6GZ/CPFTTHZs2HOUeQWkB071nv5JlIGr0vWJLCe81ME+5KsXvqqQ+mvrmWdCh
WUvpzFXGMFMwBtgrjl/XeQq04sqxfaML1PMJIxKQjKjhpRripp9pN71MEXe+DbFM
sggYgl4zgknU3QLM4lx8CXdMYMcSxVYqhQDg64Q7TkMUBZRn3mNwih7mxfPedPKe
guuB5hERmX/hz0+zODZ53GbtEVO3b6YPVcCsS8JE6DVGO9XhdR4xEjhrXiU1cY6F
yX28sjb0qq1l+fecv0t06oUXDT6c9UJD23EVOUdvycB+sEYt9SC9RcHxRZ62fc9y
3c8uJy8W+/kmHG513a7er/NyhyYF1QtU/pUbF6Ee445usxhTdy0Vfb8+VegdOcIa
3UNjMImh2qmP2NoldK8vgOejXjDP2xGOkyhjw9QUccvpixUcZva0DpkE/ObXM6gw
Nq8d+h4FNqUSTRvtlwagFX/sfUkMasXxSY1WmY93mx1yERDUkd4dwW+BWssmxm2K
4SvCL1Y9Cur4yzrJXE8XBgP0oWN/AdnbIhRdd5aTcwlyrHSNLZln96bu+UI86f4D
Spq0mpEFpTCzSBAPXELS0fN4LBzFMCW1JHJONuLqe/1lCPDYaCNB98Oz7DOLzR5k
37I7pdaFeHB9a8SG8/bRLDiQE3d89TdNs+1f9O2ySasrkRJ3/3UWiLxqturyJCBu
Ik7XPCya6xfo0w8nNzE37LcgqU2yHQqrxH7C6aSM7CYmTwT4lyEKjYY5IvJKq4sk
gCmC2Aeufq4RIbxStYSUtTIDSGPj22FsTwJANOaUQePlGmInyDPR2+jv3AZDwq8R
8jfSnK3Q2thZtLTkdWqWLnR0YF7P6qgisRSqWpo8U6GR9rv7+IEE5CgHVEmWsGOP
JldU34NBQhN8O7IrDQdhDsECgrJO94ICeJ6xQJa2Vu5pIwK5OT5SBm5Vv5VOuS8O
1zV/qcf/Y8oVlPpbtvV/mFOWl8/cIAtvuJisqR+ku7DjmjsUI/YozRaEAwUhjcrp
A60xbKZkS/1LpMQVwUkQOh+Io6nlqKUdVO2QyNM1J+k0rzp/FQIrUd0oUGbQtYse
h+2NRLL8C5aCLhXn23/4q/uHiNDHrvzJmD4GP4NfSq8zNYLCfw3M0YHn0zGx4KGS
fEatHUFPTUDUdtJPsyUPpSeJGPaP7zZhMCK5w+WwGGncEJWI2xL84D48i+TjPHcy
M4rjq/uQ0RFtNJ2mgD/+B5m24azSQAcIvgUggVfwoyEpmYt/47U2/82V3S1VJnxG
OHX8QUQoRA2lFha4sBY8KDjqcH4m1rYCCEF/yfgy7Xmn9Fd9YAX8ZrnMJFVMy73R
McYX3PHcZV2+LwmdQf9/jLvW0m7Lxw70XCODTX++5g17A+4fLkmltU/uzs1/d7mb
aki21fTLLdVSD17DmGJr0g2EavgWw0SHfQfkyds6GrRsndM2PBV715ef0Y5WaZHm
3PhX11t9BPAMFZ4CfHB30DNe+7D60Dq6U26PLwuoKXz68T1hNNIhfs4sOq13MT67
A8pCjcbcMGWZNV/ZjJznPbfo6gqK9vzZgPsOd5RG+cQs26nJ6vrafHSeFhlwCu5s
GxmRFX06u6to4Ygd3fmB8hU20s/nV0Sfxs501qzNCBe9AeeDClvcrFEJiy/f3dXr
D1n2IZI27fE3caPSk+3dn8R0xmwcNa7PSyy9XMaR4MEeANWF8tQgV7dJjjj5ACIb
ZNfeBsoqni8so9Rq4jrkxzeAJ94yvL8oF+Iwv14bl2YDjq11zQNhHxYBdfsgBljX
FD8qHtBaHWixyUFVaaqZukw91eExLopJLACDh8gqH1pM613s0W5qmgtX/VhI6mBz
1t+P6CRoYUVJjOnzIKtOtId5stDid3El7mWpCA9iPfaFyY269dvlzE20WqNFhloD
6xZ8GBN/K7r2gP/TUnaJiiE9BuXDWdpvqpycUDsxcEZ0X34dPsi4w+NuxNW2goiY
Ej/nqs9mwiEuZnkW7LGw8t01HgB+24zdj4JZ2Uj72u3vALfVIjPKse+1axjlyW4N
M+4vXm1ls4XPNh2Uu79mHAzLSgIuGFiGlxd2r03/hgHKPIBKmlBGwt2p0mvgiLew
jKGxocTx6KCSD+svqv3UoB20sAGmEs+99pr/m5n6j3AbEXWnEA93UYCuHMWu0wDl
LBx2qndj0xgkWW6au/ODYgjkb8MuJG9r2G+UD3EqtBWSdiDtK32FU4v2eN1ecA6c
ymSgYtT61yDPCEOyqI8qt2lQA6XZUbGa6m/6QvxMSrxHnGcAvw9sUTsxVMQme1H0
Ej4I1DcNmgfG66w/9jyWTyc1OW0yC+PImoOX9rygrSfvPRt3ZFnVfZSW0eyT+dx6
nrkAF8PaHS/4L1VzB/tJvoPtxgDzBDkW7cakQ9pZknYJ4svNGEuinO/NBYnhdB+l
YUQDFGTizfkG5E2SnNQNfzV9ROJlgp1ylx9vWtWVPfuqwSAC6hMxZoPNpr4Emm3X
NLoqHNh0NHsYRh49NjXOFkZcR17EkOiTRPLt6zsfXtIDKHF7HP2X+s8O8OhfPrto
B7nphoZR6EhzDyOhCeXM6OKho/I4eHSrxyWXkVbKi/0N0CTufZ1LMWypLEbmXBuj
IeIxJHIO4RmHtBrl3vWGeGK2bGJ9P98HktJkcL0qLoB6+cL0i/38oYhgtZq1iJ8G
5L0FRPwJPE1WB9Q5cXgqobtdAakJmrh/d7+ueesn+4oAFucLHfpWW0GI1qZDpsOp
6r9dFGO300h+TeDWlv533bnqWhszRW2cxbG7ahdQXUywOAc0W8PvOSSEiMDA0Xky
WCkOFyCTsGIhF3M0SsQXqQt16sZZY70hYFWMQ5xSuLmhFdbZQgLjaqhL+XQixIcC
ARgPor2ygk0hYPbisz/D1VIQgVgkAJGtzUsiD0WYQ+m5MYFEi+i3ttCfZ/HUZ4Uq
QUaVFQDVAEhqg7YeV0JB7thm4m43O93VE4EcRh6e9RO4GY112xO7zZ02SYepCr1P
K0ky79NPuYL/T+B7clHI36NNP5rHwqXWvl/vcSO+2qVhJL6cR/I6TLBOEpCLENgj
RxEDbVWLkq8OyI9MtqD2lh4MujOBXPtMvBJL70jMNVzPQmlSkyp0vwwotQP4RYrQ
rFV/jOJilHbf9y3Jc0xBv2KArd7eJijc/O/mzMl/DE0p4KCZbSJGZKmRAVDxvcVn
Ek/14xtS6LCm5JdfMo5bakrBhON6IbgdvNAg2CYPIvWp6pg9+CHgVxvgYlNJfjwl
SmhD8NFEUncOHW++vZsIipO+bW524OoXP9MpAtKp4xqu9OvswOyheGHW7nJGL1Ky
g6Z/xmMDc2aXbAXI8qVkfjXG0opb9o5HlSIERsfFaB7iwoqaMDGBzdwcMB+Ma4bp
GzTSunqvnZRm0Lwb4tMFEF+wYXT9/opJDEzMeqzuvIpd9qDdp1p8bnX/AHnMKfic
XZbgDkKqqO6cxZ2UCtStJChuwrR8BkmRq8reS+6kcbQ0NqR81f/UnKVwoGk6srZe
N3/0tY/oF//E13C3IuwXDwPLX9IctMlThOpsgCZRFv6CPeg0cUvqFdyA1JpP3Yz3
RN4SCzcpaY0hu3XnohKj97WlpSOhi0RcXVKDe7aAbvgY4JbRTuYA4Z7/bKd5BPsZ
fmbx8+/16qmuArXbsEGi+en2cp6iQ8AOFtPzQGOnxMQLYybETdmTAbn+3zdmyADX
o3Hi6dY1BSm65k+5+AcK+ptDXE9xLsa2Vi5JR+wRqj24D3ThgQtY4vyOqNd/Js0+
yR3XDJ/SswrmnI+ntvvtFMwlPXnwNr2qUEFhCzdhm874c7ie33H6915YGjLKtZf0
9KaDkK19HWWH9/2mPrToIrbpYUoF5XrQi+mKhXN2vAFoEDAzMJY3ssCVIJoV1UJH
bA0xiJivgJHlM7rrqeyS3OfROTDX+OJ5yA4RJwU9cTFPScJOfWTnoELcQ8+Unf11
CVElisGFgO1lDLtbqP0ApkuGFerJT8OxQZ8ncupPvX0oxeykUjI6cGSYMI9AYiis
5RrqvwUyOn4uD72yb1XuANxta8z+DYlQAtB2NlQnVfWps8zYW2bxz1eC/w5JvQ3i
/fWlUg1zpG6qVDJZHNSVejHNvjn4qBCaBdrrka2A5ttKqRg6s7NsSCqcGH9fUXtA
Dmm7tMNffh1x+ZS15mh9JMBXpF4svyfjf4kR9gX1LmHwUWkEbs2SMDLA2BOl45c8
f3UXNTIYSRIWuOAsHuokaeE4fBO4DDU/6VzUrv6X1Flzl5I//BTB7B1CUfgBSUEr
Vm7pYYC1thVcupbtHTAHPGx5vX1u8c2+cJvbn+t3/ihfGqjXj6dagUECdjjeJfWg
e8fpQtjjR4p2hPFgY7qx+OWxAaO8kDYPplWzcjw1LLTIqNiGOm1T4b9ndLT5YTyz
O7uOKLqtT7CtDTYZnQjrQzaWzJbjBD6Jg9UhKmlkikaRvGiRt4s0PenF4MM9xkjC
rXgH9MzHXwqqvbTcyXBFznyUEj0Qh/miEl4WQfn714B4oii9QaIAXhKNQ3fugUBX
9vLg5RQ3rxrZbKkDtygyKlT9fJN5g/LzJ+7wcXpHkfk7+ptQw68KxNMEZQPpTL+j
0ajO+vERhGvdyyKKyt5j2aC3arD4uytL5qQptTRpNWKVZi68SxIKqp7dkEvu4YCH
XSXzkygzImx+HvQ9NRqySFe/+sn02qKBms+/EWH2sUnMUzboYkmH2Pw768sbmd6I
eEkDHlL1R0En9DD/hsAQMGvkyAi+xbFkOfvNoEoNfu9+6vzdF37LQN3XmZ8EoR5k
B9AAOB7XD0eb0+T3QUZD+IrQ0NcgIiZYFu8MW+0ddWrL4w2FMXVgnzegcEusWj6m
0F3R1yBqtN0AE5+tMVaa5qCeREB22ah4oMsi4BpyiCiHCI+jJ15GZD+fArAefhr3
6/MXwQsXy8KkbMhsQbnLiT1u3N3/ZaRgQg4zzzpvJzwqD/tk1bdeZf6+u1+gb26M
Fs6QCYTSmtplM+r/EIzq45iwr21cPjApuTeUJGHk51yK72xiw4KVTjyKtIeJP34c
fJHCX7r0kq6Ys82+vVa8yPQC6m+2E0RYSDIISeLNLuH8xn5Fq1jaMst48gb8QlqP
0rtJtNHnrSyqSiu0aQz/kCJ9DBywqf6cT4iQkqW7Vya1URm9MMdE78qEn2GI3Pvb
mz5zW8Bj4v6fS1jQ8i+0SRuNFzv1Hzkweo4P+sTvVBgkw+eImf3S0TGl6xGpK5UL
x3h3aT6eT8FG0FYgR2buExdubRuhWfCA59hvNQSDVHPGvx4Kv6H0ogB8XGq8oc9f
IYnMIey9QhJW73mG1/7qF+zCNQZxfzCcATgp1Sv5oS+/NWxbR++gdwONHQ3sb7K2
eK15lHSIC9bUIAKIjhtWrtMKkbyFV6day/liH7i0MHEZVmguTV2W9CToxgYJeI+n
4/l9KYxI7WxUfK+uQZEqOqIP1czDJ5KpFwOPZImHGogxbq1lphO5hTJQwEgI8Uvx
+AAaxZE9hA7VA7ildhv6QAhcgpuJYWqFTyK2+2EHTwULAOnJSOqE06CXYUY+eF/5
oN3iHbzRAky0WAXjqTuQSoddv5EhUzg/3FayOmsNaGMxEACEsk2gOMndDE+Y2FRk
FczBiO6sUzxoPdk0ZMfjLvPpWfw0tWu8ddyeFivatOOGTCe/WS5Ikr/iFiw6IxmV
NICCJnzyin52llIm8/CMU3e3gHQwB300GNbwHiZ0CXWg+nfrrBV/Mij61JyAGgxw
gbyiKkqlR813g3JgudY1URjzIeVyVRWoLH/DO15ocWmw326Hb+rIskB+erOwHBka
2hA/BrxmDRV2PXnL+ffv7K6Dc2ZhSvnminxG4asYyo7+lmIqcYki37si6yFz/KBQ
yKXhZrG/Ro5IaFyBaeWVP7YMcglC5iNmrX/P+w9i/pUDFGVLgTIKFmZ+QyYb7sQE
VeM1pXV1QXR00qUCJUMCAnZvU3pll+mbSqV0RAsVbWaGY2Hg7ig+pmppXtnq8JiS
eTn7MdEOnQQIZP5yMq61MZNabkol0EQIQw2qSu5ojiF7WFl/0cr4QXFNxSzV1R+8
C1ywAgLQ/lITzBVABTOwYV2BPas6T7pikzme560Qrgmi3FgvSZ1y0PITrDEv//Qm
0Ghva6G/YwPihhtuEhbugoF3L/Td9MkTkI4QANWYZIE8I/t6Vv86xyLSy5M+w481
jA5wZK2zUjhTBizTNPGmI9Cn9O2gLEXC/1vcwNbF/D1eCdtksdCAbu+2AAEG30lP
Jo0rvwOvnSqmsVLHnFYlFohAm4gV65KUQth+RTFG8urPSYWh+0JJx37RYJHxd2+J
tKsiREVmFv0ZBjLtg5NLAZ2ogZvpGK24uO8UsT3Rhds+5gXmkYAkk+Vq/SH75fkh
SLTceuXawZHKTrB6kw6Bg0arwHqyAdxlFJpBoOh0o2Pm1eeI1qEMhxeKgaFxT1PL
LbOJhXMVqDuVWVyr8Jl5ppNfDQ5JR1ajF/UHKQzuYQFcs5KuSmHx3v8u+7bKkJWi
ce/SCPAMCUdUJQeXLfsFEiueSaY+ayWYp35ubQl2oEvi3TcLKKzAS13UFnrOixEh
/fC8G/njN7iCnPMjlSKSAkJy6SpvClSRgMn0p8jztcNW3yEegrLsZV7Fi0fPyYaF
JHpqtujdjzEhLBynrkjLJofHNsv5WWLPIz8J9FcFtk14AmlVFPi/fb9jTRdHSTkL
KuhCvyu4P9GeuzLHz5zSDYvVq7XvFYfR2n48iDIy85Av3LdmPNarlfEMurIKsHsQ
T8g0f52/OaLlG5snkad1/KcmWUwh6eAEEiqq36yQ/c6wWfIvgqHlxjlUf51sDHUO
yTotEhbLzKxTNtAythrY8+hk2svjEB0Zhs+4s07/txVDx0vgRHtBN7YmyU7TdGMp
tirmrQM4VvXeiK9gJjS52lYFPqpj2JnR4n9kjVFIwDU1c3Sgn7uSKM8QwNybZNYm
gEh6SvjdpukVRlf1+IUdRcaGms2vYneX5RmvDF/L9lnbsGpAjNTuRNi8DV/JMol2
wl+V2q6wEi7HYN0pfa5QUeA73OjB+RwBhT4rXNkKpUmHA25P6Y9j2PCOXWI6rAYc
PuLVq2IHTDuF9Ie6RVzVl6TIHsmwBMfR+mu/s7xkTNxenxRBtRCJKGo0qfCL7V2Z
0h3m00WQ4ftYOjBq93lZsno+Nj/Zsgc7E9AwUM2eVaah+cyERiPc0yxJJSnGC2+v
e5w1PndaY8yw14YT5qk4BBw7+IYiUCDA4zYLcnKgJ8Hu0JlmDdTbvR+S6jnclpJ8
BkoWp/SkVjTY0/6KCo67J+F22/1itcPCMQ0LIDTkyvqd+QzlcaKcoqD9iHJguW0N
j5mMCKbdpw2yAKiHB/Jq+MIzNXMAtId5juqy63AfvO+YJJZIy/e9MhA7GmZv29Wd
uyCcinbt6IJcFGmgKuoD/3/z2yWBzsoMpywrOzZMRU9HOdxh/Z1NV0gNl91AUnck
EcPxMH0116d5XcNu5NTKwf7lqbUlyQQgAGJnPcs1pZ34Zel0kXC9aDoPlLBgyRYq
6nDWivh4ScB2q2KkB7m+mERqtfPcO2IDnP69sDKuxvETTiJajSQHS8BzXJ2ZCBdb
YKOIT/puFdZCKkpR1sUMnMLC0Ozv+JLvHLqY5pfnTaBfRp5Sss7QrNLo9gNot9fQ
FF4lCVmx70WSc3RGfu1VpZ5S/ZyFrvN4FKGBrrknBQso2HnQ81Wy8KOtFlikhEyd
1OqzjdY0Y6jww6IK8lBixvuGwuKOu3WJmgo7p12V32JQk0HC6GcqsPvYnS4xMmiJ
WXIKEt17+dcrpFagt+pn3+59vjRdl9rkBnmdaNAw0730OHxnHzdqIOMzdQyvV5l4
nb1kvxp1UqqsLrJ0d/KKo+3tdCkPxi0ryLUqz/X7bAkxn/E0OBm4oJ1/jMx89uW3
SboB6VuAD28z2KsCz+z94VuS3nfYyzf7NtFxUxyaJknqvV6WKPeIXKc5M5BuSeSo
re5MiTgKoNrxw0Y5eEZtWaIQ9R0y9yRgmnp8wclCHCp57SYoCLzFwz85SAMg55i9
5NKzJEKbGbZpTCLhsP9zklo4Pr+/F9apQLxMTD/r9dHeU0wj0q6KJ1xAgv0wai5j
PPwXnnc5VFTs2hp19+hDjIVujBAKtWG+61VQZTya9ZMvadhoc4YTPoRXKY2LRhVx
P8mOhsSRy5f061aH1dOZpfAdu5ai7QYctHXjy1NZXqBR/473YWzOhBFfDcrIE/M8
4ru3elHUH4ku2rEWIo6Q7xo7B/77YSA0qYeaDFQzxTG+MFeyVQI6bW842FPh9zGL
9ATXwR+YJBkHLuyvgnopk9Ip0o8TtJXKmsUyZZ3EFQs5GBds84QKcx4uIctk/EEL
gJo2cVjg6gySM6mgqNul0w/yZa0L8CSjXlduS536u60eixvQXeJEuB8ydtIWW6Mj
3aLqSlg0GA4vPSjC5c0gOcapiK7Zayot6RjYEMCvEYrQu24VvgL3baw8rdXD/N79
RUzYN3fl8JKeByNUsT+W6xtJe8OK9mTji5gLcYLr5hy7DzKpSJtgVWnoEv4aUi6G
2fxUvVLVaR0Q/6yoaDDhBZfhlx3UJgpCktyeGOgksprsLmv6TvAhEqVHq77IBY9q
L2v4N4CrDbfbsapBuP8xHtET2zcWgSXWZ4dFqa2E9WPP7A3P4IvVomjTcoHwYO9q
esX5/ypM6V1LUxC4QKRKX3e98B9kNmyRnCTnN1GV0mfDUINafCjPKj3BntODqm5A
2gT7Yqg1C7fRidUqG+fXAVKJeLZyNGFEfnqCIeJ2zVzLWw26awVQT/6kGLyR1CsH
nlTUJyBVGzqPV1RQJPyiKY13bb8BMlL5DxccJGOhOywuvK34gLtaWhQIT6/0VYV8
SNZyZfWKz209eEEWBM+iwUxB6zHEjVTeV3KJW657dhHPDuwdbtRjhZjdgaGHXmJf
h3cUrYqFBUqR6XI+bQAK044JuN9/pl1RE7EU16BccRrymKDbsk6A0IHb8Wmy7MxN
YimDPjI+497UXNSdAwYJXJE5xc24OEu74K+GD4RP/OUT9gxRe6oHoeOPFIDHIh11
dgoq7JySJVpT9HWwK4IakyRXf4Xtc/EKARb8S5ut/TREIe2R9M8sEBuGIybtteba
s7eKTuAbrn2Kj5WK65uFskiL1bhkyQxq9zMXvGuTGHR0L18mgzirDZndjSLHmPD+
6dRi/zZHE0u40NcDMYAbtGk+DujeBLQhFH1Hp/rQd8h4WGwKUOUOelWaZqDdubDZ
MDmmdbFE+XLOE12d0q+qnc2OIRJRafYS93XXgq+p3IKjdVG0xsd4MhUWPdnYNqsN
iA50ChIWLTW2F03hwvcpFnvwhRYvSFEUt9hcCYaJNan0wQwhyD2OM/u/MBBc01Wd
3KM6+qjxbkHobQxWN/nOlZYOblBWGAUIubA+1bSwqesiEgfv+vV7IbBawqPggOXV
jZYqtmc+2YkRlrM036veKOsW0BYcQ8qKpSIdDocvut4rjxcP0WSAkYVLc1Qf8KVt
GWYZ6hpIR3UX5TyGakpSb4MrXiIb1IiisSc0GaTwToQx7lJki9EwY58TpIghWB6e
tM8pNUlT0L+r3N5bBZw6ErPrkFfhIV5bzo06Rca8eAVj4Af9FGLvJOUFvjhsHILF
JFJN0CpA1Bc9s7+PCPPnKb43zJCQ8PCurUv7DNZDs0g571/gYXVAYpYHnMTaRtU1
jwMaz4yt7RaGX8FPps+DoWKTglYIhJpJ4A8s1YSvoDw62l5+m+PzruzdVq5N6DQf
iRV/955vPBmXCSHY9Z5fqFMMtIJVeBDqOz530iXDt3J8e+s0sydZwDcsrtLqUySl
KShk//MPCBPS9tD2XfqYFfAV1Tn5Y1oH92ZLbx34RJAoeJPeBm8o2IxuiTFzpeX8
xrLgk6Rs6SGYTNyhFrsxTyjQ1JMvzyIthAVPGD/i/tsLQ+hRKrfnixm1qlCeOSRB
0uvzSdvYRZRqTQ+6TmYaDxMDxBBP5DtCZxz6Hiv4Jk4GUlK4PNb28d7SZlNVqQau
GCJ79yCuysSYA5vn6hPFnDfOcDvdkJQi/HstUxZPiTYSmknAzBP1FoV7H+8ouiKr
IEoLEQJmwZovtJnKlaLOy0TmQxaReoDySwKisgmk/XwF/MHVQNCyrfqWHTuWCMd8
0hccquyqsxsCvEQohfGzTden4+xhc8bnwhIaq1GgEWLMBaiYFex89NPTD/CKsJej
2CREU4DDvix2ZDo/9nKFygVQQtWcjPm/RHVtOWvpk6tOwfnZS1D/qDLadIvko9aj
T4bik9gRHQ2KD+e7XmMHaqXuX/d2VIpIEkQCAy3wfnFMgfCdwFo9viKAKUZ3kMNg
KaDoZMHT/HfiZr9NYn/uKHhNsfEqs/Jma9scN2XdkdpUPXdhjF1nxPbv+7gjKvR1
X9Pe+TCiObl/UrjBoyC1jUDLrqK6sABuAVQW1y+3i/M8vfeyrFGusKLSdHplgKH2
hCdTLwRizHk5tCok5mgyTAXwXPebnYJam0KPd38Gngj7v7zlPHMUOefbe+mGVIrw
HSvR152aGZJ/Buo4xMWjMhHIgM7t2uD1ddOKEAOXbYVERrQdpB1lF56dkJY7G7Am
aRf4QZHHWbwJVhcmQxNr/wPB4yteasd6EZKla9425XLkrzPduArVJoi/Lw+FyjgZ
OcdXhZBSzloCg78hMoW4tyHL8QVZgU6Ps+Tpy0Bzs5VfyJy0C7QlpV2rrO2Hk+8G
tBx1GtQPngQ5D0mFLNVDDWIem9tj55NE4rw9Utyr9czkEPGMvfZ99mTDnBGfNT/a
OXZOvmEFQWv4lkASlSwpeIpa4lhlkW9Bn+Xl7ILfrlFWxw34HV/LA6qs5bBlOY36
ubolzJ/xGRsUYmOX2Ufx337GZwtmqveZbXeQ0GULAgD9YYQuiGAtY6voAMJAlDbZ
MbM8UNcZWtTNHBNcglIRRj/38N+uu7zAcdQFIxuBQoWrcdBiqQxee2lfpyLwd0vM
KeexVkIRjkanqn+9nDZReOaw4Tz69vJVNtgUTimT1aDGAPaqzAzs8k7peEt+2JlH
x8E/RLqgvL23K9UhX8rRV0cUymsbODVtK3TPwSuiYze0PT+34JwazorW02VT5yRE
JIyMDxPjYAYy8yCf8TMVJ3qJvsyX6rVDynhweDS6L72VlaD18Og31gZO9KPxVW1q
3DqXcvWtmjKlvPd0Sf+zfrJWiPTEK+cxXhGrYGXA5QwPVGXfQYUjkBbhBuH8pKr7
9BkswGgjzJqEzUW2hfQK31VnIv9eulwmvhzRxVi8AGfszz7fNZ8ZEwr86j4wYQK+
CW3r9ejflNun0AAfQBkPzaec3ziSCgSFQXNEik7hckWCWNnyOX+nQHseEI8QchBu
CXcusjVmqEkqt6QFbdqJEZEGAq1tU8pg6Mz0kOAkA23cJqCdJbRA24OG+KHeDYT6
hNiZ9KxJDhgqmBDe+J0gNHjliEpS/Sfo3mp3mVqcFDkP3/GpdXmR39q5ItCTWpJv
e8d/2thKZBvRSd19dWFxFlaRvwFLDeDeOJLBvtLYc1UptdkoXSxzU8NOASJ+q1ce
9hfBGiL7KupEusDoWU7LIhYn8V3ye/YQVT/Jou+oV1JyCn29gSrdlBbGCkxHoIm5
KbuyWOL7TmFI2AW01VY1arKEdlxkTl2qlxILxlBZ1azW016JeTFSJ8JLe+gV7R3M
YP1KOpoeP6LxWULsNqwQR039TszR0f4DgeHb9fXG/40BJiHc78+P9yztP4G2AKpc
6WZRzpcR38zmH4LhDbcg94uK7EfBrrV26ODHSyCozEo5BRsYoU21r0/5JRP54ExX
wBDoeD3ylaQ1SuNCO30Aku3EwpAe6uV/ld2QxnxbsytW7uIowXiO20XWpXDm7FZE
6TGwJ1Rnelz1tGkd3cR0Q62rG8mYZpNl1K5apAc0WI5uofVPvYfoBE1EgLknG9CA
dzDB2uVzaYnDTcyWouhX3mm8jm/efLWuHvFN1PFIdFtOuKvZbjJzhzIodqNjOB/O
MBmbYh3R57fKzp0W6bNGeyKse9gPge0nw9+nuZjzHfXkiuwxGyvxtsIMBMKtV64P
+e1qihRIRNC+DILUvr+0Iwe3sCQJOWxgoEnGx5U1iwlosSr2dPvhSw60b5t4D014
a8wTMDLxIWwkgTXP4fScggeDPJV5fRh/IpXS2++wwdea0gHLOX5pAy3yIQMECp6B
n9TnA6Y5Xr238uh51n5nngx4k+aQ/Ie8wX8xpm4muD98Ck8yn/nqNfED6wfPxb8e
WBUu9XoAanu0ca9Hovo12eCPgXE18iXSKwY+N9/rqTwWP7FvXosnbrvHgGbPQIsJ
rioKAw2ZzpYZEzbrjK7N4kv9orftwspk6Kh1Z2ZAbZlUwxhQNJWxJUD/CdGwBGwG
AiCsE1nBRUeG7YGuVeWTppp5ubX3OMiFFa1P/ErGopSzXeo+Q2sXdP8mebieZP21
cRvv+FFb6iDLZwyEVT7sMjhwlTkM4ybcpCB/fs8QvjVZ3SsqPWm/asTD3HjKnBxo
UiNnb9w60jnLz7bJjmzDlccnqD2W3CmfhYZEQIv1AXP8lQa5Dt80qZchm9r75dvk
3J6jCeMzPNlEih8OoVju8bebPSMgzPLg4YfIvA5KxASqNMi3eIuSA/GSGbGRH/y7
pCUqVV+5zl5L9Gcn6F+GU5zNmtwUdj3YeqNqEpvN9ycACQy2cHDjbFVxsfzVaWZq
AlnCM7RdofdqxTvNyS3WJLCHCORUKx3F4h2lb3qr4BUowxNDg77hI8DtcuNelWY3
2npDr8Z9Gy/i+Vn2SPU6+nozVhXTE1SqTmssZy/AhM+cKHzkkg8zYhqaURofHpdE
1fN40FKKT3nWNE/ec/fMyYhHygLzonXNUAadbby/Sybd/ikRw0kMkIQxenRnc1BJ
96qLsymPHTnqIa68CjRor/1g4fOEBo/l9POo/FXf8M6NZenoeLE11x0L/uxP5jE4
VPYuXxYcwoC7AIcdXO9DSCOO7elne8Ti3/8LUp7cAq+T2V267dTfmDDC1cX5r8K9
4wTpd+Vy9kOsMnU2+dga7RzYZRyYGoAbz2w4UfmKlAZceAeRU5ZIqm8gUzwyOIB8
94o5EcGq7y218lUCF0XzwXlhUddVgORXKTKgtfv0pRSv1GxB+Dd/XmvvUkS1Xie4
t2qMyH4OZzGHgUcowgRfJbIkId1krB028+QielwvJ7wSHLfnY9cD0Z1nFTw1CmYx
VnT/Puqo6yo7zf5NYMwV8Np3PeGyltrvhnaofjdBBlO+w6h7MUxEJVzcAIWR0CMg
F7Hu1DkC8rCBYKxoG/H4J3FJQt6ud/Qh5gLrTOUtnQxK5+aU71sOsfj2+NEUwnYW
H7ecOd+E0V5ei74BnTT7s2PGc/rYEvG6eF3EO3iB5vwnOjFK8ybmksqzeosLq8VS
ON3ojkbcVgDcHM8FA2OH5tm105tOBAWUnMMCp5o9SnYX2RGCztz90zYqc0AUyHZy
f4v8tC231cbSjRLepM/aURlKj5zGL1mdfWzYZgvShcEgqbp2uvx4gzjH18TtPfqa
bbhABc6+UUmYEBJ3Ja9gM+q9RPaWwW2mS4sC8Sus8oOOM2quLj04rJkPj0qHhgmC
YJHYq0ROZfR/zMDYXbQ2bEBw65M5wZ/PROSZm5BxizZF9X8mebyp+KQjgudMfQbP
H+N3uTNrH5zCwbT4osow1EkX7hOMebRKzrUJn3Jnp2sqPiA07yubPmg2CW4KpquQ
PK6e5mpNb2s+94nWnRAwp3NVW6YAJGK6owZ7pYKkxknIpOve6DIze4dIUZQOxMAd
Bce4wzveeOZ/r4cHumJ71Z3bf/22zAZwAIZSlYjWmXDhYowayj7rdJMkIleKAOFx
jbwCT9+6DuTrA5/ODj8fvXmvben8Ee9zdS/qQGFXORW9iyAQjV5E+hap2RWwkvKG
ei/4CO8Og6uIRTPWcEDKVq2y1l1HKqBT9QquTMVfU6A/nLOsy64zhY+imxCI9zBh
1fCiYNv4T2ET6IeVY4u/yABycR/+fXNwR3TivOy3IhDp1VnNjpQrPbKRih4FvBhk
Ixc01BygO7C3lRleWNknn0XKDZfUA1dzsYA552MVz4XgSS/JsLQW10SCA1xSGaS+
RCryhIz0LfiN0LfGxudM87Qq+cCWZw/x8VX8kMxhzv/PtgO6/uz8gEznm8NyuMnt
aSQZDB8cDiRuKQZbMqhYgKdNApbAZER6c/EGrpWNcY7/FaA5bMfX2v+26NbwhUFz
gHpCjK3cnJ7nXtCvNzfWjOxs1gtXjgFF2l38T/zroB+LkanFfO0YatM7TnGZzPa4
ceJBXWTXi6I8eflSULulcXdkF/ZSq9I5BhuX+2/JMMwqUY8c+JFJpBefCHfnf4I1
2W0v8a6njkHnqbYpo3AJGFV+ICsQd0YO0bY+Q4TwwWNKIzPELAeq9HJ662f8kSKA
kwIvrxVPt1S35mC4OTw3ChrtdJLHwLI3aDQo1EO4E88wHNvcun7x2X0tRxsxUa/h
UQpuAQ++TLwKScCzNwL+E+sduHeqq7QPVz2llE/ImZvDmZdCUr1rMzzZ1wliEPqG
SWu8Q2aCmX3EtsvhUlMnVh8fNgJPUyydJMRytKFDLYRPSAVpNBMqP2H5uTOSPIUK
HfAHsMd2T0dizXJfBlzajKUdJgeSGe2XrN+1Ih06eKaWvf4QtM8OvhHuwHO62/wR
BtuIBQaZ6dKztHkdIqw4oh8NotnFC8GHSCPFJpX5y0SBWNiPtF14NY+tbGrn1xNm
fpzvBhKXnDRk5xM71wbSeQXYJmpP8bjJs8GjHecMYrUVCRM6TLuzAWscGUwdEq5f
4QnReOfjYGehsTacObag/sLPt1bDovq55rUqseyH1+yR+/oPuMlrPR89YCo8v8ld
sEGQ/O8ndztOGlCbGMhSUEYe9pD58YQNlFi85lR4RU17SG5l3avK4FsF+pTo7PoK
UjTwg4BYpJz7ZC4pL8bOEw3p+T+rSIcUgzQXeDC8vjVfy0UUupl4aFN2Yz3H8JGU
55RIMDa12+63lhWX2CST0mH/ObPEfTUAsl5aZGED213Zm8p19firjAZ2Y4aXYTBX
qtgS5tDlPea49yFElDoufg3MNIbWxlOkycDGDZZYOU22gAKxpXiRZmTY2xCywY6x
94wqOYAPQ1RGiEvCDJWGn2c4uuYUFzHH2Ak4RLfHBODI7xN9ipKBdp1b2swKWIKG
djDMj59Kj0itjYEPU4kC69gHrBZLEMbptuvvxDtTEIGqw4xnVuw2F26petDf1NAD
7Ypblavi6uO31Kjmfq21vOIP7pNKxS6R6AhWbMxzVZL3Mn6C3Tc3zK2WNJQ9Mys5
ijz2QzJexcvl0N/ea3yj9VgKrUkqpR5UfxNpr64cz5F7KwcvOLI+QuhWR8Db3Obs
5gPJXi5lv2I30gfBbsDZhDvwAq2IkTMECcyqT5lUGgJkn/rgZsqJ6pV27Z4CL0Ks
jErs8k/n+fIuIynU8IlQdFlzrW6ad8EY0H8o0gxZo2DYjKVsu+T6Is3VX8tSCeeR
l8nYuAVKGULzMYyhDsI/mfalclS2WO+/8Jf/9mMRKr8gweuJKVQoEH1BXtAegl2y
5NIldF6WFCUBhYGO3FCm0oBGMiESyaYPy3qVTY9udlIK0huoTQ2l/+s5alO/4vql
JXzo2C6IWhBLQFkY1wjoSkrkzaZybnxCZv4CBN+Srx5ahRIVhsdPEh98oXgmfD6f
xZkzIUNGkMGqfZ4UJckoOWlHPlrYJhQtJHPsDjSCY57vQlPjq+DHT56+LCxSV1+S
whCz6utMqMX7pvA0Dpc8j2wE39qI2U9Pa0PnsixZwHKXrZUXyiJyCfLNN1a4kqjs
XMbLwZETKAlC24ARx8TVom+uFAUuOii/K6u+kaibPGj5c67iUkLuMKAGz1HvqG5s
2vVcH+beek5Vh433ff1gbaG8GcLJt/VbWm4BmOcFOl7bWMwicu4SqK9HTEqXpQ2T
dcUSIqsyZYTFjENeYoPUJCblBhD/cpHG3kXgqFQ/vPKgvq0wfddysVkBv5YmoT/+
/6M3M9lDu5f9nAjC1HgkO03yQDOOpN5cIbqQ1pwMBPb7Hl1Il4xwsdYNglM1lUw0
DAsMoDAuGTtmMKckLvcCsZIZ+ru2WyIn0J+HZpdcd397AN3ESBsxr5bitR/0AltY
mTnEUjc2ED4K8UVo5qHkz12BteprOez9SoY7+1giAwLYwV8tjrH2o2+qniBeyXm3
W5yrq9pDiHVM8QZQXGyB7Fi56Kn3wy/NGMZv0v7owbUD0xm5c4wBvWUMSfSqgwvH
uNGkOgwEwkW1sdrX9aFUhBgB3iQ9mqVh2NyxNaxyiEPsrelrQtgYpbMAWr1VyWB7
mgEOgwJH80GPRNYPpkjdwdhijQFUYakShgY4j+FOMPOyeRBi5r/brnt265fCSamn
q8WVztWhDSJ8ZjE0xKisytCCvrid5c2IJcuBAUXOkDKE5TgX6RJIXeyr7cMcXH3T
XTT5XNTiTg8weEHckUshncpCZD6xDnoVJy5d8GimfUa18IwoM8bUKwEOLDxb1yUm
zZZjEAyRgr5VGDS5/YC3r5k1U0WsEwRzGodaFQt7tMj8E6QzTpB2Mbb6hjykl0gk
zE/ea4Uwu7Bul6PjTrgLeRr4j2IIZ6XoWSFlUQwzUP8V2T5DgqQcQYxRdglC3qJY
UL0ONQaDcddV45hD4gHhb1Yos341iJhEVrlN6hP3OCsL8cQhguOZ1i8oDK+9Sgd2
2xnB9o48oC1VV9cZqe2bnhhrmmOctIePJ5Q/qZy/m2ZaWqoGdaeOyhfZMrttpY8P
yxbrIBHZbOk+d0EsA9A1qw8MEuiDFE8qObO7JDFsRZMa2YkHfYHHDl59l1IYg7qn
/E1/uqTWm1V0gR8pXwxBnbgNBmNKkR9sTyrr2dsvath64zM46npD3+mCdsIuPwJ3
M2PJHAPUN5EDHc9iGS3dK00zlutbpbAOLLL8xbxOyQtgy+4H/z8EZHPZB38T+1Ns
f4WIh2BsOmKGauu2hwAt0OD2+Lm13UAL5MeBhgP3FKBFOW9Iv2lxoEk9NAsltv+D
mnx+GnZxWaetXOsYzW6eROxKhiC23dBPYmFyzslkKGmYGfAANowMVIGmkPbzJXhi
tOA9CSc5U/gpjbZKTA2fFsbaY0uIbZ1FJQfxxpXd8AiEKMc2mnpkk48edYnCMclG
3IK4Su9xlLKwMHQ9XTXgaHZYQppUdDdfVA2YC/3ltii/g3BhM77U3w55CvPbWzIA
GvvM5AxnF4N9XiG9krHvxrIUkx7KO5AK5RI6z8ILOShdVJkA7N/hqv9olD8BK4xo
5i3K2oOS4O3dErJkIWRRGqMGlgNfuDo8LSYBLrNmuUgvQJF7WhVoDAfuj+VEux7n
UX4Tqcss42YKV8ZsPXUQtnbV6SZNAzoRAOyKlvwC3RWj2q+8+AnP1tZgEKtunGp0
Cdz20TGubGBXtkCOGkrm0xpOPoqVB/yLf0HwiN0u+1gAG+DRg0Gd8nc5y05sY8Ay
lCLauvtL2Z6y+dthvcabZH6A3JX+Yu71OAL5usb/+HwAPWgHb2SHBLCRPUyIZ0J2
joesgmpmNRpguyJzIl0LEOVPUk+J7DodaAY7CNd3R4Moisdk8DY8dEv9TRy8rnBe
NNg6gaD+jA3Ld8nT2m0zGRpFi2EKePyH86BY0qk9LzN5x7m7Cqp6DA0xsphMPcM6
7AZXW25XdSdFs/sMNzey7NthXBVdfQvxHHq2X4nq6WO+wFC4AN2+BSa6kzmlQrHZ
7ZH33utu+6eEYyZBEEqGNeFy7COIB0+g+KSS2rbGozkPN4D8yPPx5Bjk7YBuhaQg
q8WcxkyBW//h2ah1xOD5oxZmTKiRE9d7Bj9dh403c5mlPDi0e4TZyt55DMJNkc2y
IUPWG8ZaCMrrbU2u09r5g07ioy4mrtUczkEJ+xbNlHQ6O6cuslD7fLVsF/PEw6hE
EIgw5RAqq4CJ92k3y335oyDg2WUwlH0pvXKL5X5rO8QDlyz+CYpua2/XCWtJovmb
lqqxObcwcYUPTBOBASKYKGItCfHkfM/dgalFV8hChgcbI6Cg9Irf3hS5qbGqh7xV
nD/kfpy4P7LN6I18M0DI12YGOz7be+jgNOZiHxcwoiKOWLJxokdVmMKDJvERGZjH
tBUWtihgGYeLbfvMQlnQFuJ8ytli7eKQcHr0UpN2/ubqigpEwwNlOsLX2e4glLcI
6MtpCPUXZ1OYG7Ac8THTI4qXIwMzXzKVZL4CJ45iL0jMUpMUHt0Q7DpNWbLRTQXa
QtSNO2vLbDV2QPUxw0fBa2e6GtkLtBi5tgkceHqgdSDIGhqHebXRHjtp4TWRxr6d
m65I/Yu7USw4QUml3iYTOM+r39zuySGtOtNNHA73lVHSMhPtPP+Kx6Xk3BM9zFYU
oOgCeWDqG5m8wcJbDyCiY5zSy/BFbyAYb4b8iMiH6Kd2T7T05Z2GXFMzh7Tb/Mz6
V+omXKnRDYYLMH16hUasfb38tdHXHlJwI4AqCMbspK0R0RGApiTvYwzn4YEcyZJK
9fbylpU0sMtdVfM/9oERHGNmRE4My0DNf/0srBlrPpMWrX5bVw9jraSO6p2Lr3f0
LeT9KWU48OO36VNvp5Wn1cz/x47sj+tWZueJ/tx5R6giHwwPPvUl1Nk4nyqUzggi
FbkGdtcJ7g11Qdect++lFBMyiiB4hkX08x2l5sNIVjYO75DPt458dzm+Bvy5Obi7
OSZ6oMZuCma/yFJeHOMHiXO4kwCIzfT5ad0NhjOezBT2iNiiRd0lydfiGqlaoQZr
o3WJoYPQ7ufEf4tn6fiHq8ll/NHlwPO6i10eYJ0wDs9KKouGrpDOaF2+dl2yv+sM
TcoALhx05nuWhRRBxuKAuT8N5x8xAp/0IJuSHhaPwK1/alKPjfcg8NwKiimNcjCx
FiE63S32P0mZoPw6x+/p6V0funKCZw9EbhkjJ9IxbRBrTH29INvMjl60FwMYvbAy
jva1WD/nHW27JnGGSgSDEjeR3kbJEajT2hz6nlgf1sSR9UpJm/GPYheAYSy6MTFh
kKwjCSzR2wWoNdkFo5qiOfOYs/U7CQycveCzDEbBDeGVS43OOxTmaLGZ0/xsmFe9
gCRP/9Oj3u0L6IiT9Z8hVcL28iMBJ7i9Zy+HxNeHN6lv4MMRY/fvVaaIkKwp8gj4
Nbg1pxSJGswv8HsIZ2I2jIAU7kN5C0j37C+lLHPLcusIdXdfjTAoM+8QrDkJEnPB
BhenS1PbBAfDLznD4uNPKKm071tzirblF/7q9YHR990rweTz8Ytd0BPe2meokrC7
u3uUiLBXj9C+4HJzaQB+7GW0L+vocue0DWlbXeAAadBrkUf6MdDanZDgZqEXxAXZ
cjVHCn5lQyX/0lON5XliIOtcorRkOR5l3MErHhkEgG4q9DQ3SzmAqBQCBbeF8x/x
rj27kTwnI5E2wa94eA8lrWo9HuofoD4XQPFbZmAqa9kSbxEOiEg21/jjmmxLaoUa
V0IyekgxiyuFMHrLWUcKLi0API2wdC4lKwqQpnMeKNVSbCuhiTtjvjaDgUCveqm5
NlNRPCXWTxY3hrJDOxmLtbKb/DxgnrDV4oKzjVNiS1kryVYvwgN1L5nhvzhIlnpL
++4LKEkTHaQEFk+pRxSkn+nLOOn4l3qiwVcD9onNj1HsGf3j+N6K979+ijfaWfYa
9IMOElcAX2naoJLy3IgxmXX0cOOnnHTIzOmiCNE/m5BqJehmnn25hVzGbjxQiF0L
pCPdJ/yy6GNrZLn3kFopwRHtaPPkI+w3b4b6y6ksWVAfBTadvzif1IqN1B7IFHKd
WBCU+a5zgmx89e5TwyjXKnzTrOQk1WM1sFUOiSsoS0aYM5O/G6MLPp+P6ib+gl0W
/G0DFTlUbeYRKTZOFiiE+cUNjRq0ZCdxF1VOjJsfqJPn8XbHRKu5d4iDo6+PJvfA
ThfVEf1foshLodGscye0MZAZ0hiaryxMMkqc0WM0lDOIR5I4K34FKfnUwz5izBFs
+OVn9D0sys9abdie28eHTZtamsVjlMl4Nn6qUSa1Wi0KCW2dSLjIWMIEu12cfuhv
nZ2UV9AW+32nCEzDa4zP2URt5mq2LNRUPz7hzViwmEjHFdSpRrU0YyUgEFP+q/Bl
fnhZ8zLXHWG8Z40h784eVLmZaCJ/7fVc2xJaTSrOySDXpDgzufmVzCHsyGarNUgh
9Po2ty3HWzTyCHjYCPx2rD1cNA/S4Ip0PL1OQ3+8DetRea3vXfHm+K2usAMrbn6q
dH3rauJdQ8olsga5AK+BrH/dzgpHpZ+wNOGkk8GiIX+nGXCd0Q9nQJvLjRMN3KE2
bPFUd4MgLDWjMSKUaWFgPPiH9eofqf2dWg9xoqMDO/x9Y3izjjT6u+xK3tqYRBvl
HD3+gQ+yZe8tuDlN5zl/QAAFvdAljEysAmzMW2gdxuq+EyY+du5ws+DzjKCIeNcQ
7pvTsYOb9tOLQdNp9MWORO65tcAmpRd5Vftadqlk3wSEa/JEskN6f3rolTHj75re
Is3Mi4idk85/pb1iINN4v79Gt6ReBkCvbuGcoUDzmH8g8QINxeikxCmLjmPiF+IW
6OOLgbaUDnsfIRRMD+D57FbaxeenRLBhk/3x4+uZDRmGBqhXvdfli02Yg439vZgY
A+1tZWyixq3t7p4/haEKN4Ek7Kym+/ZshH8mysVWEYm6Js1SwhVBkTyJBfzju9hh
uvL6TZkzGIw3QbtB8Rv+gjqozPE1cZMcAL7Ui8FqjI7qedhwKHQIi+KOOGv/mYt9
lKo+QhM6jjzm2PY6iZbzuGwMz5UFk1gKL72dVRwliEPIrto6FaDozhWSSIsa+JN+
AgbDqo7HDWfeaCOOnqRrvK8BPZqlKuAmnnj8hNv1iaPJ31Qpd7fRSqIo9q029oFd
geIGLIaIgPAz8oWk3rKbn86kVh55pGNeCaGuAN0eMQfuRK8IiJz78ejhIrvkzYDA
oijkzqTZgqOKRS4uL2MCfWL7CTy09fRo0AB20J8bbzk7cw1ZRQcB5a4tn9C+hQ0p
WR1IkeWcs+6JvessbhmeAlWDR3TQGfhe/nIJy180Vk6oN4u22rNzmqgpwEozc417
18E1M+MqdUR2J28YrzjSsLhiOxhhMYJPEAYfDqdLFSN2VLKc9ztg4EWhyECglgOy
HaXFBX9fqebq41j0OOW8vZoq2VCH5uAsWAQck1i5lWlhd8LaCnBc1OYmVY3C4adV
25K1VkvUwKOonV+0+N31iDGOhcjdOVM+d9wmKDvmKIHZz2mWjfUWk572s5jtUtLL
5F/tdHVdpVVjTap/ZcuGtE34xLQNlxQnJ+TJv97UFQopVcBGrQw/0NXyqMN/+jTt
UMyjR2WIFJAX3L36WIsxBlNWcwBIVT7tVy054oCb7eXqi2PWSOe4HXPrPWewz+Le
8eJq2HI0fWydn2DZ0/iyAWSVVtBmHZP/0Vd4y3VWYWyu4AG87z9JE8O+mjiWv05f
rEyVlTShVMtWEwEPryymMCJRc/gti0Z7l/Wv7uILG+beS0eU+hw6VhaPGgM59NLH
vByBK2zpi0uD/PRxer8YJc8zja/KXuurtQc2YXHuivdyZEVgbioaSSFkUO06x6xJ
On7DbZAOkFSr60fJcoVV2AK3Ol1vyBmRqODFfGT/bDqvCH3lEGpJysduEjTt71Qr
Hih8l8pBWrsCHTAxJu/gXJo6lvOHOirWiHYDmOx+bWPr30CpAoWEtaBFgjZdpBbX
ysIteSO/smxIwuFajgD35Za3kmDGL6YRHHK/tHbL42GVmz03GSzxvcCEzB+Aoaxf
ULJt8dqZOe8PT1ZVcHtim+1AQDj4r8YJaKFg+aR5c1NLf9dLMbw6lzKnVmn9zUgb
d4KfNHeeczXrZ7CHs1ObqQqjNVBhnRGgnKoANWlMJOuKP3sNxdoe4G41IxiQH5k+
qL7XrKVGiWca2BvpAB6JZmOVujvp+4sIiS9W8NW0Fospz8BpVAIkQ/AanbF0oO06
JTwAAGtx8uOdIynIYECXF5xegU46PWrciMb8XAEwgXaTfZ61j1SeHy3/OeNgNaar
0S3s6Niv4J8RxpJuqsfQY9NCBZCUwGfYbgBxPq2PANFH9Rb9tUANvmeM2t5bnovN
ba+1JNTo9BddiDOErR+gNIC52r7Z5vszYUxxsTxiTQXGj0ICOdDAPuVFXqrEhdvK
I/Y+1SDkIyIN09QeYRKmVGLp91WGf78zY/m9Vr4joEvFhPssYvupcXfqd4JcMgG/
PDQk7sw86ShZjLydv0sC1BUoEJMIUrrittaXE+7Y5bQedPBmM0Oh8uF/P+jq4IlA
H2xJx+AjxOb0iWCBFR6fzwMEXIy10IrgXdCFWWODCfgICzGtQuvpfxz5x7YVfXQt
ZQevjZlraSq1PrbPNehgqf+TnMepTJyxncImvCjTgY6rZ7v0Rkm1a075ix1fd0R5
eKFqhkxDo8Xh44ef2ilURsB8hjIMMEtpOsvz5IxBfssLoKSTlxqAwy5o3aGmOH34
MpxbLGWnW/nGnronzomxqJIDAiTH1yOmaYkUJQUgjUTDgfRNf+r4vaM4c/VtJt4g
K3VfyRhrsjlYBPavpcIIraNTomHY49smq2UbHS/wyP7q81neh9HGLq0sq0nKGuAK
WwiJcUVZYHkF9ERCVTq4KL/Et8T7XQ4ss6HDL6gNMiAUiwgGXA0amDy5QZ1r1doP
0ZHugicDXsvFGGudIA2xZZ+ylZVa4H+pv9jjATV0BE2eppMhT8JMLfUiBK/d2TvI
61eb7iyjBlU+ufyjV+UCYu4eNqjmPvBux5i1wWj0NNNTEzt2VNFb5z6od0SI2WoM
bjnFrEWGtZps/yaIf016gCNqKtrcFNyNJc6OwgrCt9tqi0BHYbrLtbdth6oi3EOG
uRepKEUfSdPi9056taYVS1zHOYmjezFvrcC595+EzakCm4Abxo3Dw1Yse2mZFLYO
D8iQ/5XBxcyb6wV74DbKSY7nP4vnaXSsyXeyecRDiyqHdy3k186Is/DMEz2USUva
vRzLyU5JdJeOuLSKJ1Z5XR6MoNKYwbRMUNxgXhfwRh+DMr98tEsne/iH/Fa7i9+Y
LRwV7xC/iJ4UKmKRxOEdIIzQK3xj9YmUuVZzIREo6HU1zfpeFu0kXLCm3WqpBYxi
cfiw6BL5ZlBJEKPF0u2MUXcXB0l9cSzRf0zE4rFy+7enVuq8jypmqlJ/tAWs8AmD
2JX4GxUh0zUQEw+QBCQDY/oMQrX47BGGQboLjRztzPU3JWyW//jdjQwJ+lQNKtgU
DmlwJLxWJ691m1tV0cRJg2xXyF8anYKHRDWWQZ7g6X/H7pC066TZiWJYH5d6xlHs
GyAlCnALMvi5wuXZA+sVO3TjAvseLT8Epk2eHEbWaMC7GJrDV3DgDcc/oZA/5LX1
zVdFna4LakgpQXTNXfT4+F0a5wOSQjoaCk3fbUNJSUB8WVu4IsPVpXWeTIBzb6EF
fEPFnmDmSJ/OCL4U1vpFwLcs2WxCRqxuDkVcFBKyW3ms/TlUwgL7szCQs7cfb7X0
jnLy2Ylm5ib8Ra0HdlV3ZGRckoDdl0PFpcHi7R2mg7zKO8P6kY2EvpjxAMlzseBq
udytFzns8yYMgfyMUYgzckvjnaVLo8tBHeKt71k353UG5/0Z7RPFnf2wwzGIAgjD
iyW+SaYz3A39kXrw49RVzOEDKsBMs7b9Xo6EK438UvACMrBx46QmutyhESEuERFq
XeEqubaOFCUVK9xa8VDzVOVbC2PmL0cKWLeKrIi75tJ6XvnqvyCSnlxCmyErd+cJ
ibSWxX1RbOe1Te7OHYN0q9sYbSIBzJia1tFjNOAmvqIWId2KJxPZgXcwloZXcskK
DX+Mkw2+ZIsJhkorgBxThJBN7OMqN9OIv/5hYietlT7D+bYFUuUPQir5Hy6M38Uc
foWxS/G7sIHl10e8DyA5IWiZAELfNk2Zr68yJlsgfN3uvCd8syKVCNwaHSP3ma8z
eTIijNPYofBDKzNDP34RQN7ZyYtl06GBxBIVRPGCBQjcZULctCO/IPVDaKgsM7+n
OZfUDI28OEYZIVu0QwmQOTIwnVTwYHELV5Om017Q6zoUAPYrp7aTcI3MyKfFo/IU
53cH2PkG4f77jPcPYUH8+g4np6h6QixcSG2eSxcNVklRFrC5jmMvqmOi8B24HapI
MGV3E1G0rlXSCofsHo5Ju2g13VgMXOWgoMracTJN68PnEo+U1agZnJZwAeh46US4
Kxu8u0Q7LCQp7jggRvA1lDaTUstfa99aMqa4nKmEb+wIvhMl/ktC62+Tx6cBNLwv
sMhodBKnn702IfdDiT6cMvL/bTWx9WsXFQKCLoPq28wtEdRfbka1dCOf4H1j//ZD
VnbzfSe0pBRI8I/nTHFORzJBuHa0ISNpo/5CbyaxQJAwqVFDHopV0awHu5LfB6ob
f1ALOAKngUiEYBEyuKaGAZGjG3eWA52PS78+0o2GHb3C3lxubB0L8JJ3RO3Z7BUn
gxNM66FqGzy2dbmCirkJgL0d6nMV+W2qgMtyqEDJBle6Q/4PMBAxHrf67OC7cv8M
9brp1XRQvH7Qs0QY55wK39FNOq/9YBOz3oAvN2GZDpExFsrIdNg775VbkUoTsOSN
xp4isEv3CQNdLwjSKHgDEec4QuwlF98FMDjScaJvXVEEtUb4VAmhaihLI0Nnx2Fk
hQt2j0ufyDfLeUC3YawHwEttsrNnIgt3iS+oDkjj9g5iwm9OrCxpY0D4MEGQO40x
2yHVwo7EPgVWmBJq1Wd1sYX2VG3k6YLuFsWBp4VkJlpIluhpVWkVag6W2R4WvxJg
Wbcqmdg2vY/P2pvOMQ2bncWWw4mR9SUm6cczPSAcPxpD81eqlP87I4HyLpPyzXUx
/TpjzDQ0dIIIFmVetzrdcadjzgKhJzObhAoVT8MbpKgNWtjR7jvN57WgPj5E2c3Q
bvXNizMQCxBgwH7m9usIlM67OaKd4c5OvlFWuq5klb/bRldvtCvczSCCBvhzkMNL
drr0+5OTl+q8OWTlhoe4NqmnudZry8WvCGijrlkG1BD2B5QRPiwmcbaULPddjvmp
QtsHaTKxjcx6PUmh0nii3YCDwhT9qZ2ekzmsGkK2j3ijxpA5zl54u7jAsrj2a2KT
Bnr6MM7F5GpGrTxtsxk0tJTg7x2d3SiuVCIL7a7m1dCXo2NslPA+0lZT9mruEBAL
RKW2hO4BmMmshMgQ1FJlffjZALudzdFbZBFkaReQUoqAkTwNJjr5DVayX/0T0Y+S
eaifADnxvlskPp80wvHgAhAzQPxS1opfTyFSISrMCKgtr42JC5UR92bCvSK7gZy5
1cEsYLBFevQWvD/+cQTp7DDIblT1OAhGpsrGtmIZ5kLwE9JY6LfXiofWDOXflTDy
kYijIlK5tUwwaq+RgZd7nRR/gAadO/6qbrVelRMGACuVD+WEAdzKNdC3ZUQ/m5LO
TFWbnaMskLNluDhZ80GsEm0FIUt0XDJCdj2YSDaVIf+0n51iRakXPd3Xed3bmJFJ
G2mCgtwD6Yrz1fwQfcNUDypdz2RmYB063ojPfw5SNxXLmOqXgcPfcKfOXLbGVmP+
bBY+9+0sUS41XXflmFF0rCQFoGALbPGLNQriWbJ5VkJnC2hPhstHvKNedtCJS0qq
Ylzrg1X4lUeRN2tnr4KaQ+Jr4qHqUev/QgHfdZabYiCOVZx7jZ8KCt2Sy0kWTmYC
OkJ+H2LZjhZIbeHTnRxXqfsZBEAjmSNX/yRPMD18u2GC9TzdgNIiOYNKjn6M+p0M
QvsHhijeNglxzLfrToNhUh/LA6uwQQ4K5V9yWBAG+UbC02dyDG6Cxy6yeWj6QvIU
1nZzEZol9fE3WZX3/Ukvtme4k603fCGzy1GYv9xzw0YyGQXU6d0pOqErnc0XKjqs
T1m4ORU8qfF4VIIvQiXdEHrfISfLNWovhY/G2SFYFenENbG+/VZ/9FY+4EGG+XgD
CJ/KJDLlwPUi3UeB0uyXrFGLqyZ/i7DsuGzXTy45Bm5+uEqMLKDJDCrsz+Zyco3X
Yx18BMAJemnQZnTnhI+ODBa5LloTaVd7oI3wLrRufNm2tFK/B6BcJBE/fyyRBgpn
4XkcH3EY+uKnFbbsCrCBApV+Zl8ANOupW15ZQh4Nf8/yd6MzdX+jZblJoxBv2f3P
q/kCusD9sAQOopT8RiP/1x/3S2N7C09CfqUscEQJABrAfcTulHVEHaLEioFXVFop
lPZfENx1sLeABSEJwP711yqgpSwGP5p9muNw39WECzu2mdcghH5zDq+UZs8B9d+P
uIfx+9aWCjOrUNX/HRteEOijAbsfO9Er86PDKPkYMoRHsN0T+Kwv9+ceQwvtZbah
6f75RfGTpOaNzV3ynv+nYKqATIqIEIjeDSQyYdBbv8QvgU1IoiJYp+pyNgtItbKx
z6EXdg3GEm0l2kfSTa/DbIkjBJ/j2sdstUq1F0FG+RHZPaMGiR+By5fsV7tjKFKf
EzwzXsq+3NKI9mzxNJokKTqq28Y6qCLHKPzISo5G0vzXN69+06pJgFJg+iUu47oa
9lDNZOxXDJwrTpAZwUwOyJSQhCzmIjb5phdTk4zr3UcI3TmJQHpGwNVNxTZuojTp
CuL8mchaAnd2p5/nwIblugGyaYHwqSM3S5foYe1JT6/e3/7a58Ps37x8b2Jp7bAH
L0hP69Rdmh/p64TSulgiFMxGBmjWxaKwb/q24HloU8wCrm2G9sa3SE6Glgn1YL6y
sAgFFvMMAa1JicC3Xrx7c0CNzB3SvRAKTskpPPiqNaB+jqjK9Ry3XgRf3InnBuCy
W6lQcwnnfUMw7x+ugzmWkD4S1ghYjUCcdtFM7MhjGoNwZ2XQeE3PSIu7lDdOlR89
ADhxf/HbALfdv9ZgdXPjST6Y5AkqfxNSNkS+lM2HbLLVCC0Wf853KOpnpUr7n3nF
4ISUQq2oFQ4zvLRYGMn42/eVAwbHWgRrNSV/YpQJE2rzRH+nz8BY9pv4p38DrPEr
U3+rDXlK6Fg1C3ZJKbpqZJe0CGKFbJi4aTP9QHzgySijkmvrb8ZN2yT8Ac9q/5ej
P7B1L9T2kFSFaZUvTrJZddM8+TANizW5x/adc5D/7dXrjlBI1/ZRBTHk3l105bFT
aw1bv/pStJUrOI28YUFlaP72+skm3J8soLDtkYoqwrQ6Oi/5Uu365ACkPAJx2K53
zS22XVenULuDpXRyXXgYyEW5p3rvuTF5CqYNwOhjX8PkerpLREefQ1FqhRTp1aKO
G0LbNuYq/Yejq1DuVSmcaKKbi2hv3AVHMd+l4n+FfNtFlt1MGzFGkYx8MZv20oqj
5Kfahq23RkunBA/dK46A2y1M4CX+RvY4XFfAw51iIb1fBx3sDGHfEI+jLu7ph2ul
DlkXzC8En2dUHUCQ76AH47BGQXD40ZanChuAHRuNPcUAxYUnu9yWBFw5J0zOqKMo
SB3DBDFm0SdkDPIvxikCX7qzZQ/SvygYYWyIGBtvPBvBm7Xep5huCnXytoqcvP7z
KWPXruKIQpgDFXRdHTi4ONuLRVsuYhoK/yf0g+89niduvsukv7sIoaAOtX52lRcb
WNw1LQbVpfBwDhECbFR12sIyPicw/zeoxWh5b0sA1DHx6l3ADmtCkxiqcghYjF2K
H//K1Pl57HkoDn5v+v0YAQyn8wfk0zDgOAeKn/3p7gP+Dej4t32R3U41ktUAxmF6
GC1YpHEy/6x9xAOhLJPSnsoIYuygPo8hR00RSvcf3FS2UtRJJjiGPxA6FT/AsWKI
ljOhGuQFR6bHw6W14KmPYmXWswcM2M6pmrUdSVMJemvaxnzOl4CK62opScOrTmyS
IDcevnzX4c+w67BuyrcWtcRlKGN606qFdQzY1dZxuk9kteMzQEtM8ii60d7LJZj2
c0P00s0kAnuwt23O+jSztnopVt4nKlqI9mbcyYZTzpQtnk/XnAW0PCw+utR0bZyA
9mNTQInI8rY1JT1HgY5I6poQrpEOQbk8lfKSpDITY9c3wBlYIZiNfO4wv3orq4SU
WRIDuU+w4WVFuft3Hi2fbwv/4DDyEWX+8kssYL9NAGs4iUMzQxjBlQ2Iuug4dSzU
yjGEb2SqjTY9LXMgiCz4jKyFkp9ARvCzAY7RmJWKe5LhbXhuTXuv9e/QrLITe88e
B3XwpixJqSDgjOEATdsjJ+dWGaF5Xu7na8Kp4BgvQoktPBl3TcS3bCWbcfNFUi4d
YnCOK2PcnjZr+XQte0KV7BELYtVZ8SfEyfgORpEK5opCu66CKOU43KwtTMJpOLIO
8sYOEBezZFrCCO50fsoFOMRUaarGAz4uj/KmLc+OqiL/HoRpMgZaeAT47vTd/50D
5+h5ya4vM+skBRSLWBP6MxFe6BE1n9moZJRqIPw9TME2/a3tPN1vlqOfhIgr1NHe
+OwDF7V8E+MqjTNZYv25w51C/HL7jXVVEWHcQkbE+0h2qe+7cDqGE+MyhiUBws6s
eIHt6/wQq9806nFE6eczgmmuDIei7tObGgp1e6BrHObZBys569+vLt5ERetdU6/J
JNZvwWLXucXb76QY+Mxvuk+h6IzAe2H286yT7zt7VuNxB+JHCYKRmNfThDTOPYUa
fXNpuQROf7JwU5yOTN/k7m8t4NGiWIMHjNjzqpN5ThNJLoZXbQ/neW991fsB03TD
QxtP22X3lctN8GfkrOdG/+hR45n0qnquDEbNiV1VphAzCJ2pueyDI+q4m0swp3hT
xGvWQbyhpW9dLt/eC31a4HKoJ2qwy7bac8zh/pHZewOLeZqy6Eqh+ZwyukmbfEKI
KbS5vKpv6x80kxlg8J71cx/zgyJQiEPlWtn6qygUeA6ZWuzkHyJQYz+qoaemSehC
chB44pCI5miP1lURFeYaqERggkpKcTg3xah+7MaA2IpYE1gwX5TftnH8dAx/T0VF
ixz/ciqGBzl7If7R1oaLmw+9iM+5CO7HILaiBYvfmbNTI15yCz767j5PqGW5YM2v
njNjpoaeEJuuMcvibtxXwnKw8ozVB+kwU3ArdSj0VUCKP6aVDurNxzdBtTtdsTPS
Pv8n6qL+s9Uv+xKWdUaEFKpI3jam60sfhB+kZ7kmxLs5XYTC8X2d7W9HOieeEg9x
1GwvMhE3Lfj6dPgAIOR7iNZ6l6wel8hU6jp4F6eguAYZ3jWCJPgZFbdHwxb7Bl8p
k/kuYIsnx0eFIxGY06Y2Q4OpH6zLwD9l0mOOk0+9gD+LLYcM6aJuz5jlFbtYoiM5
UHBODTuKpgyGK8YfmfSXON/eHga+kInsrC8JCt26V3yKvsdS8OnThqYpXqLgvmW7
qqhweX7vTvWn6oK1mKr2IxKEMffUtGuZEp6M/X+BVD3eHgZz/2QRvjbmGAlZuZmS
XaXGl2LCmg3OLjJB05lihGh4lfjLHS9c/XrwS32ahyWqRP+PfPq5IH1HcARTQ42z
GdYt4XWA9dDTLSXFoq5amIlQDgSbZc2xY7RxZLlBmXjTzq853uSg4i7atPLTkqUl
pdHhAFdlYPjVMh8CWcDYRh1A+0TmRlECjOVErkuBCW1MXtnxqUWSn7MvtEya+G3p
39edSQ7AYyjsZPWehRZqATGAA7Q/oy0bqKIQ4LUcc9bvN8HQ7/jnOrYfogG0YQQb
YnY9VkUmHh5KjcHs/Q8PuRkbs8NOb8a1CuDmNVCmYXdmoYHzeT8O5wXGfeeKSu6P
2nvCY7Yutu2jJz9+TCZt7abIcUIcRB5G0eDBx3+cN/NYL76BVRmc0ozBBmSam361
vzlAQxmLtAiBTKnTw5EyPWC0F7wm+dAgXkTDNe/ONRa5E0hoeD/vy4IpfM5vuysI
xBGWGPQjkQM8TGHFZf7E/W/TYplVjWEwAItt1JZPl9ci5e0+hmCXTfe33rbSusN1
xmXlmSGZTUXt5Baul97/p9dG4i0/QoYuNbJkpPaVNHXm/39PcVqBsafqUvgKeKeo
Bfl7OdHAFQr3AyOzyJN6UHV6h8GOw8/yIkB3tp/lWE2DtdHgfz4uRfV2z8DGqYo+
g58xRPiXbla5RzKi0vZreBpLp6n5glnCfLVLLs62F3NYufit/THBcD77TNob7rvN
8zSigia2TUHLQE3lKBQPH5ChnlAYJlby2slqDK7FEZfYj4sjzZ24MicawcK9jREA
L5pfBPOSpoHSAtZrrWOvcXgHzM8tQJk8ktiis4D3HW/vP+IYNsyVGVi8KafS5RV8
AvVZU/48XaNJTdIUnO+c7O2vn8rM6sSZh1E24a9SvK8Z4tEPmY5d1q3rMFcQE9LT
QGxdQnXL8yxUL8KtP1gcFy9OkuLZUQMyho5PSF4jH7OfrCAn2YZ+QgmGC2cJ+d0z
4psfqAfRnXoJjWAmK2fMFS1YVKahfNovGgYo9JFB4vSzeD0thFO4WFOQW3Jd+8ID
8sk37naByN1Rt8cN2xQzWlg+VTjC9HyFDDRzH5KqG+Pg4l34r4DlVu6deJPRnfSd
yfWEizPLjS/ZhQul+aDHL0qTLof0iSQvjc+pOvji6b/Gio3UGhMLzfBSzePrg7XN
XjLH6PuVHglaRzpy/qKRAm6tSq6+qVh8oK2jSGxVpZJQ7DSVPvihQ1Oj+FBKERyF
HQkWLxfHs36FhMr/Lr4iRWb6wp2+/KXRWj1kY6saw8kbDNSiMpRwipYuy+BcEYb6
KkFey4FOzRzd3nLDh/DdUaoHEUSYQMmQxgpFrX2v9roYOSanHjkLcSvmaZscRUEw
XJ8ttflGIn9Cyy1xqXM610QyoipxVuNDqyxW11ww+2qfAcH9pjXI66oa/YC3zb1n
l0BIm9sOV8Wh0wyxlFu4kULV2Bv3OprtHTMG03jNmzSsBrlKxJSHEKmMj+qtNPFU
hBa/UI/oTofpXSarT8VEvIOGGwdTqlZLHEgz7WRCCH5sMhk9XATkfzInftiqAEXO
C7ekH9ZixrU1wJS/TlUj3tta/v2ufzauiIsCg6jzlSd/0h949Q5vmWpE6N2Kev3X
Sf6+mGUiJ60DbmJmzuomdTpZJ7rCVrJi4uWK24LhpIOeOh33gsWNdCaMs13H5b6R
CiLsB4+eqiE0gSGR106xQPaMyitAx2jiqHfrscuMHpXogatzfmeKLg3J19PFiBXy
0HAHfsbNHIDXnoDWmIj9SwuvhJ7YWEkFg1ZT3XIHIhx6KTV+kD2+mQ4eSLBJSDI6
Y1UsATCCTU8sLk0T8puMy2yhRTzoKZfmwYwq6Qmz7A/p2LAlyjkVX2U3WSLfxyN/
VbKR1TZL6QVzeyfcl8BVdl87hCnUnHCttwCwKazvxvbLyFtameQkFXBHnA2/qeYS
JZ+Cat/xYpCNepWHam+GdQuS/jlyXC5rTvZt4MfVvub6PL94YdbKP/H/WB1fHQL4
xQYWdP/ei0eJFUBQhheXmE96laz8DJXKPOVlfRqpKiaf/h1D+WjbKP6Jg+qR2D19
WGndOyrFMzxBiOXpv+PiQtebs3sE6qUudKW0cKGDKbMccDkWTr1329+DsnaZPjrP
1AlybW0wUxZ2amSnb/a7WyLSTzkznNB5o2w5iLfWflBgdmRzD6x54JyhOgj4cUpV
QLXDzkeXVkxaMAkk2mLMdMURxOaaqzLZFefUeA167uq0Qz+tEalbAK+fY+fF/Ryu
2Cm1sUlFXzh95gCJDQIe9+0kfBzPLYr2i0Af76n3TQ1LVV2P0aH5hyy5Mm3qm4w5
GwggfGcIrTTxB4Sc+sDJNy9SAz98ftlGqxMRnSE8L495JVvEzww34/v7RT91qyUA
O9yE/KZU7gC1tuaSPJCQTSsu1SvG44YFRNEaaXmFLtH5aUBllIVKDqHGzgoAatmH
UYmb2EOqd0R1Y7DjpaYdjr7tbFFgmHQyTyfQSivvYgvQ4Owt4IdBw27hF2Hmd9Pm
eBhESjdRm8ewEi3wTctRIVXErm5dosOnLQiXg6givGu3u+d6kKcwKpXOAWvQcYqc
6dTYBinjS6O5PtXwF+IKKBMwFusClaf+/yMPRq4RafggtP+oKWZra+LXxunkffpA
i2JRqmXc6QrSjHZu3MRf1X8PN9KLqmPHRuoXwlM36a4tnlPnkmG2YLP9Z7nHU5zk
fv4Yv6mnnr1K2fqEn9Gwpt/RoweokDvqTEcj+BNf4CbSppzuHwptQ9YR7+FEtsAI
m6VBt4FYxbyBd3vbXY4m3fzZnVLTtLSQZCQ1I1pB2Ht42dTEGzuoYb+yclB1P9yl
i+4Ld8/mbCkelMs9dUXQlaV52MFKURH4jB0XusV8cir055y+K/iQmag7Cl4hO1nR
8GXKtfT7FG8GKeeSUKqnEI8v6jCUMmBRVfybHByy3q0LQiwibu42Hv9a0gDG8HtZ
tYyZm1iKrsfXA5dMB+VJpkHnQFjrD1H8SvEidVKZWnsg20/eV/63M47iZiOWoWjt
IDH2OjSasu/0x+69VJH/snr79Nkh1bM7DrxGWcoekNetSb0L0iKKF9ZgoVheN3Jo
0q3bJGRQzay0MWjqE2NrMuom5n/cMGUIjOkJmAQQqC9+biwZUn5ACxfeALvNQBST
iDebNx6O+Qw4aM+3oeN4Zt4z1JH3JwrCzvaikYlb+UpDjaY72FeOkvE6LwrI1iOv
uARUuLDMciL7jmxfe+dvBWpaXbYKXLt4mg0uwqDU/awsWVXt8CsSfLIC38xjjFjo
zHEK7pxU10snngrMl305YSGS0fNQKdv7vF+7sPuGGQ36qY5bpfKLe85R7mrnKGFa
hbMGiiaFIbUM2WJkNP+g3WecjR/4tJqdhhFDZ/K5Xj1veLLE3tfsPKKpX3p/d3QI
6Qu0Po8TglBn9ClLJpWf/cdsv1R6BbIqaFa9LSoSNhCGUrkXsWvjI7xEwsNeVdmv
5rrBCIkGAp80m4HUrSgjZFr0aTEU1QsCEjnFgco1BBD2d1EZDatg2djYgB4uQIW4
wpS3QN6Bat+3cD70q27yZcS4+/LXSbyRNl4gPGDoWg6cuq3fioKxi/+KxkArI415
Ya8VJ/8BFP+pG+wI5VIKnR5Egfro2T2bMavSuzKIfROb3gnPxP88tTIiyE2/on10
+SA5r762iNaX/Nghkv+ydsrwuAkNFJgel7S+aiyMBO7TFTZXlwlxZh5xhGBEt0tJ
WFAH7PypD7HKdrM3uxKAVu/F5m120pTzFJWqBTSccO93oBysDV0kMKSECLnzSzF6
U8wN2itWW/xiolJXh53H82oc9BE2uRlzIu5UxpdIGK9ZVGJRx770SpXwSfvXdw5J
T1llL3dXNP/O/t53IxvypqmlcNOCSjkP9VgW6L+0xhF7VAgR0k5DqaRxhUkSX5i/
5oxMvlTZRE+96O+ncnRUxUKcsPNnd6CiDskaIumtsUylSDm8VfCEWG9qE/8AFNsw
Ad1mWWC+uuUBHfUE0RtCy5ZevVx7LDrIglnZBAOSDCTF92ks1iSyx4hU5xuX0gJG
8L8abMJaAAfAz81ogF9N7RmCNJ3qLeJGIYNvU7iB+DotC6LkQ7irD2qOXsitIvLY
yyCX8x1G1mEati7f+EEb3A3P9hFvcvj+1s8OTxmgsnPAqy6TTWQnPJTUMGMVsKql
4mj0dQjKne8jTTL/Ns9Ln0tH4HO56XAvwwsAqiI0nP3XPXC7SkBMB8vcJnOpWARQ
mtlzdhc5pOkDKwBwtxW+DJY4uYew789+C7grKDhQpEp70CWUG+Kg4alJUYAv49EC
PrULaVSi/NbLC+wn0yrfi82B9cYBwI7YHhOXJgzD5Lz0aDg8uzOS4zCYphnNoct6
pQTEP/citgiBwhmexFpAMInSEFN2lnrIFR6vzSi/Qj2+L8pxTJJEn1Fy4y+kboGs
448dLBHohBuXyiqVM3NF4l7Nw5yobdfGkJ5n0vNt8M8DVXx+uGiqicVsE3T8qWO0
38O7EoOBofpw9mH0iLfoh9JjscewHkgJQyKT/egbAzxdd2FcJRxBrikPmJrHAfPR
v9SK7W82hBJMRZdMN+i/xIR5wF8HkdMSmk10H3wRJKjJaom9MneMZCLFFOW4cHxu
k174QJHpXYvFBrVOkfXHd+LxjBqJXjrEwnqtd8MRIzSiBFCFIwUncHsafYct+5Bz
QFpPxg+nSyekHXX0oUNX5uvvZGIdBkaf+tfWbTVdG99xAsPvquyc4gJUtBLbpmJj
Qb9WZ/o12WHX851xJqkej5BFXK4eotyTKQEqRVpEoyxJSj6uL+LWxGyeg+tpwEIv
shkRf/mJVPFegDav4JkfgzWaQrs8RFIxzWy/6MKJi4RDlxW3lnBamQCPkIRU8juo
dSd7NmEouzxxWsWiT0EPhaduBmU5ySvN+1L3yxBM6oNmzYZDu+DbtNKW4TOh55MK
tVPBbk4x2aHBM8Xt2B1/1ZNcZjJppr+kW/lwRk7K0e65C46a6ZhF9FTz+ycZ+7Nw
QdYfBCuOn3cQVf30BMpUjnIvAemmzErqfPIWqOuF74O5TOfyvKRS4hIfiC5QG4LD
4Q3ogv0/bSYJKU7j61N+kS/3O2QSLWW0rWouxjRVZX3gEPG+PZnsfXXQhZ1c5nWW
Dm4D4eXotH/18x+NpDa5T5vrAB4pHFyR7HAsldRtMu/XbT/4bA0q0O9GMyZ/eKwx
EO95TEdlDBuPazbGaOL8fJf6Exbbdxu8C0V47YClROhWjEOuwP/BfWC9GvJdxM0f
Fr1/zoh3O/zJ/NZm7/KJjxsO3tHWLd3I0ph/nv+8PFFFPZLMYXTsByneOACYNtHV
SJ2zLq0T61IrHj/h/TYHhxIweBc+Pj09jHgFvbqv3YGkAmfajP3KSMxs4TyzziW8
V4E/Ghqq1WqAwf7VyZOCgBMNzg4O8ct/77v5Or4XZdtJYskTaja680f+g7hVzaws
epm1qeWFXHaXDBkk74GZkVNwJnZ85hcvNE9LRNxZW2gAi1lzrzzS4jkK0kmCeLZk
if0cxyMNre5PC313NFevkCIAehwQa/ljYT+QyTd38JJilZ6QlliWi6Cu7Z/l6lMC
oYuSk6MvasrJ/Pv8dxWKlPVRok/TzJrrVC3iIns1zGfmJjHEnpvxjhN5HEzpLsz2
0IH1InM8vgvgTRcNjwtEzSHzMEcZFa+W1Yj8wK6zRnaxd4PU9JXFNj4sueenegRF
QXIED1L/8aee6hSUTayjLq7LrDPBKGmH98Y84KNBXEGxhjZo+C9t/yldm/cgMFAz
/MixZARVE8Rhdt0mLoxssux3H0696aDLTPdOfsVO2ABuNlar4gyHG33LvBVGpxsP
l5YfYKl0Pd1HCqsTWJLFHcQpu/+VAYDxcMFh3pZJ3nV8zUtViWeol7dYSGxY8K6c
EYICM+Zfi1lS0cXphcMA70qa2hfioyU3NI8hFM0Y3ZkG0NUrFi3wFV6juLwsKDtO
0zStjJNH63MTGVK3dPsa33Quu3xdQNyL2Czqnfyi5LA5N5jfn2hnvz3/jEhYwHoO
pRDGKQRte8EHxQpoLGAoMW3OtZjMcDtH3/4qDWyJ4MzBHVY3zVjZCRW0Da7KW8tg
8pGrfpMbngZOohtSWK29k+jjzmR2BJVQFRx9j+lLMclxnQzUM7P8OAJWpCKne15p
kKvcahyCNMqNu3T+3kALSAzkDbKirh51uHdlG2Je5gndJp8m99M+tJWxpxdw8RBt
YGIVIJwEND3EiSFODGOqsRQ3jxJLV5Oad5pvEpXeP0Tha6qgfFgT2eRcNLU2T/nU
0+cV+OkFstaNGaoZef3xjMNenQDWIL3lIXEVrVOwXLerdemUTu0FUn2j0rmNIkRE
8i/c8BF1LE55zp6j2v01e9zdBHlY6xTzLHPD/X9rnG/X4RKIt3eA9b12vTo7QlGM
qxRUhuq4gGc0XuYGeASqH1yBl0Yx7d4RT0hfoMk0d6613jdBfoJoVPiQKUEMjtqH
17CBQuoFwOsid+MLx4VrwfOnpy0a+pAjkoWYn2Y7rVOkYuZN/12qpgJtCi7KVGn3
ysxJgONrU69zrbbAAPf4FayLdyYC7sQNFH1tOE6XpliYfhCFAXY+5bQCFZec1y9u
fP6tXHgiFsx1L+MWm+OGhDpGyrbgwaDBXm2flrLUoli8F4jEPLtJdVUd3828tIQS
xKWwuOqXYM4HrAVs1+X4xwIrkytCCumUqjaoNFHyuLRXmzDD6DnFnnpfzffZXUcT
L3nWqqwbGayinD2SbnwC/UOeXCzcPVxirD+7DrpEiBj1F8GyGSPjmxvTKY4UjjgP
PAn8N+ylsMYLzwWOllUYBRRW3N0AwMjGIzXI+qwJzFO5YRSd2G53yS4A/em6xbEV
FWMoaGTzJnIeK1F+7AL4ewAihSHjNk9ENzUzue3X2Rqu4oljYHBPoXgfUji14Izm
S2ks4oLgmOX/pd//LTHcDM6Su+JjlK5pOPV2FXsOMNogg7SZHwD6w6jxy+70AzW3
6wsn48EJtM5l5Kb69I+/b5R/W2unZ9LBd1wUBaYJ1LZi1E/aY1CEjTu89mjvM5nP
26GKh966nkcL/zlNM3CGi+BtcwJHLJJ6TyO56Ua/ntFvYoAcv8STnfnd1WU2cEYA
rnk7bEgPr+FpUZ+8FpEsCISVFrXzLjwC56TIyu8kD0HBXR3JCJ21POXIAbbaWnCG
Z98Umu5KOw0ZqchE5tThvMp9sICeU4P4vmThkJ6G1dt5X2AUj1Zg3WIA4a+SIF7d
2UFkdrhNhjHjqeq3ySvNTXmvCivQOfgd5cE0suzzmfdSAjZHx/91qTTaFtm7YTaa
MUwKWu44DbVhNIUNVWW8u5Vs8yOVAAIDab70ax0m22h2V1a5BTyJm21TxoKfdLO+
WP1vMr/ayKHck7OFp3WEegclkFogZLFaQi4fC+tdndxr6BjA6zeJXRvl0elaWQzy
QpA8sNvs5zS8+0Q+TyqxD8A129LHT1xVuBcUOzV8rj05qWYwSiJOQY64+MtP9HqX
GPomHhXR3CM9EQ3eLQg/TMvjVYIm2Hxfp0Ais3dxKxM9l3azxjybmGOgyZK8L4lH
QeodQ1G1+/R/tqih8sepu13u0SxSVKQal2nZAtsM5oSiqAuMzVKK8qHlqMhq11UT
AfjaXCJwvDCsB15TMleKgd3Md1qyQRTDP/cXeybjLQmiTfyyBTUUxh4zPBPbdzen
8M5AEUykryX7FFyUWMKTINZfG+3ZH2+KJwplO/phGVzVj6cFJ5KI1GOhlvESNMNT
2uaFAZY1MBzJFeoa9dQE2B2U9eQ1CpvF31xlJQtz4KuJIe4eXuy6e4ZvXMP3clLy
go2iOuOsez6o+d+nRSsLl/1nPVQxc8SUFR+g7vY2FhQAvvQ7WgwA1nWtTh2o987n
iXFDLu9hufdNFZAGFi0yXdS35+POdNggDwb7IGRGYtOd9qu6uTiG5asXNnjLsxZi
Fn7x75vkIv5Yutqc5VYbtaXtgcj8W6ylg2Y3F1raAw2JGdkJLeEZWZkrO1rS+2FM
M6sr4D+tSy80Md2pAqM2XrVJD9MCsUn77eE3tukajRwtBhCHsZJK+lrXkBgQyooS
tBNMK5rnqiB1OzzQE2HQb1lx9ZMZYEs8bmSowgCraFy0KoeZmlb9bp5YM2PQVrWp
GFjnDmfG4b0GD7iAIXbs+ZT/VmHhUwZh/ZPKxNgolMB2TjqVM0qqJlLhabEUViOG
0H2xOyF3V+Hv3Za7DfY/Sr/7X4w2MBi4GkOuMoDcChSMfrGHXgJCGOFBfxY6dAbp
FoKB00iChm7/oDalihUA5Nyj6ubii2s0/yIUXHlt5etgwK8LjlgCyCNQCpGp4wZc
n8/Qh6XH9fAfoHSmCuE71bb9j2SY8phyE/GUSc1brmu/o4rXOwPAfsICjYIdg+hc
nrSUUKc8sBN+N/otpidVtqH3JLNnOsMZI2ancYgqURnMrRYdlTE04SA1iJ7j1FQ7
9A6hXn10sXFZ66Ih8bGPCsT19pyn4HI2W5mn01lHTOf72+8GnqNwP1g9MDAAax2S
l7VTLzd2qqhvNZIheYJD2wVNCEGZ59fEUuV8+t58981UrNABXsmlmCZEWvMLhFU2
ijXLOu3UerynDW9BEmsCanM9CVwIrfkvCRpYd7ys8END5GY/+saTtPnmlEKctkfJ
+VegOIwjfXennz+50qUgNVkxHRjr2njqbi26NDFiqLwSTRYjToV0b6hx5s9w+4cB
lxuHzm/NKtx41GemQrJboshS7qFL8rCfi23s2VhE6q6600RQuRuhmCw2CZhyYDGb
XLhdSlpXQ4xUM3gsRcCg9Up9tLUunkv1njRyheunm5x6ztlwBC4K1mXKSi2BjMqC
pnacDu7ABpclFpt5WdWk0lKsfBXutbk2pCHcqHCX+2uCpvxY7IL3ydAwuc2s7Dpa
gP0BiepsHD9lTkM2LYgYXU3BNz/IsknY4AGyUbJ1iyJeICUXEvQM6J1XYkbF9ERS
sgk6NLxXpAYLi9BNWfDKurh30ZVbZSY8C8fucGwNJCoB1aGEQoObWTfkpKU2Wveu
CDpBnVHASd9tFZz6KhnuWE39NLQaow3gXcBXCNEJJ4yGoTb4/+YOOwMqYMDl/YBx
Yt9r7sIXKlRQoUflD+za7cimY413ROudkZ3EDcl85zBHCG/PrwoskfVYsCQ4wUor
eVO4qvoCtblw9+6EJ/fHjyu+A0wxo7Br3gXnu4tZFfXOHW1kc450qL0RIanuGhvO
3r2G0qkXajqJ03Yc4pvJelrdXKRXHfmgO81I3mZ0RyTEcaoJDqBBQThuDBjj37oR
9dENkq/6AP23Lx2DeGPxPqMdP3o+apR0/L7IcY7+cSOQFF3KAb9YMmXhPZNnb2gK
wt6F4fRgAm5BNCm6vRjGuIeiQHdvrfiMtLqdgy4CDaSkikPvw4SFh7E37qdq17Wy
E2TBssV9BcoSAZUdGkOTtVkhiVxjss5evDLvOu+9JLpeAVDVlSwXiS/apl5wpcLO
ivTIdSJxJO/AIZwObllAw0SWxNECMbyd1zGZ5NR4hILQBoJZwo5dwSVXPIiSoDnC
UTJHhg93sQZH0GBtrvzoLo0wLMhZF6spZQ+6Q9Pq6gh+Sdy7d/+ConfDCIRizn71
uDltCGOUosjaEVtvPUayLzCEIAPvWF/8Ze0k8Oqkyfshue8PqOhClH7BbDuN+b0/
3YImq/FF8t4fU+OVuRFv6lo5KI3kscsU24fGh6x3fgd0JQNxPezFEQ7mmPgrITRp
THds9UZg1mOkjYFYHY4AFHJ5PC5WwFxGOJECN/1ROeWAmBpHEdeEs1ZMfyJFwlx9
kZdk9YQ9do5XasiGAX8mmfRHMcbGJDv/rhdlcue7Gygc9QoFUyjUkdVrXg13x0QK
Rll0N2pmUFm6Znj4xmVCzS5uDIeU8plFTQDTQjITTFX8ogKydsu4Y356Bda9Sjr2
XiXFSOXN36DmZcpd/du39+Hs0L9hfKSS84XgUJujZkMFcSFwXPoIK34Wdnig/ZMn
YSSszVOxvAvLH9gKTNNJGv3O8KBbzpoPccTM9YVQSAesXBmpoB49982WfN1bC0dH
kpN4wPv0HkpeEm4+ciHCrQzIBZBdikjbCDq7WSo7vXhKrZq8Sfh14e9I9oo6Gw7R
+zIfJfByn9tLSGDmcjay2IWIBXnnp0h7rxUrHBQs2B5MAgi/yh7CQkVJSTQm78pV
uJO2F+r6DLpEhUkYfmcH1XGkGpd663l/9fDPhhnWkiapIxKbp78AeXINkppq30X3
APeV8M+HNied8Ydh8EqHMeIa31nOXqpzfg+nJSIK1+rul8+fLZEAHHgv291ISivU
+H30ZxNjY7z3RYOACWHv/wvfhnAoLSaVAyfGy/UOd86EIX+7gL4hlHt48ErpMbpR
9hm9C3iP3GNp2uY4edVag4LFjrRinct8FKgrRLkZgHJ0YnO+jzztwnWrqeAhKM8p
0uZ+RGFgmdLPRTH5aJexsp44C78r5KmBQGivKzjoT6vFVvQe3qrR6oTDyM9y+u9/
kk3iAuD/HZj1DmQ46kJABJZDkMrAPuUu98Mmo78tR9UzXd+cWv3Ssd88kDtMiWK4
aTEs/xjnf42gsxJV2mol+RAnlFk3xBolwTZEoyCwTg13vuyAMZb6WO6FY8nbprrv
7BHIg1ktowBBwm+QAZYUlOQGyqF/S/g2TOt0biqcIWlustqbTelS2dlsXzjuth+W
2DZgmfupxPNEfVVBctTB+MglgwZ2+6eRpKgUob9SAOqgjYRyFsxgEXDkgFOamwyO
pOAw4ATAiaaN9TgdOFmldC6bNy/TSnGoH3RqHVDi8lLWRHml0E6fMhEQgANMg9rt
jugWQHU0AmzA2QxsL7gZWLyM7wTVz7ehfj+3EtCdm2n0k2CFqXT6ocVQx+HnImE0
f2hH6xbujS9gBrEmsWsTEmUPnUn25TkazsShIKaK+TSHhSCDE93Z9R3LBPU0tAFV
o/sp15egSPLgqzpe4bF4/TUZL2rd1qRzCssu2oHh6WX+puFWqiqhQ7sTqMiNVjFz
hqMN0WiI7hsVEwSxdJETOmWHFF+H/F8KbjmU3Tlce3osXBY6/1AP8wNUsPX4s/Qe
KipMLphFniS5W2epjg5YrfcFEfzko7muv1CFJSR/489LSZs1+9RuUYJGisOs/X2L
1l1xhHQVhEX1/HBrWnu1jwKss1WJj/nYNSFeijtKhTekz28uf86ROTok8rwk/CkM
6MA3iw8HcILyk8lhcnelQZaBamlTYuS03BIj5fmHwT0zMc+yoX4By1WOdWlAgpad
+P4CM4nuvbRnxqRSQj6/vRiukDXUIESqZRYl+CX8BgujNI+0p00Jib7VU6iN14Uc
stzQQxCy2WowWunS1ofzF844zvVmwygNdQHgDssjUptzf92DSTPGdAKrO10NtqVL
L5pval3FcnQ/g2QkqGVI/NYQ8cvXHXVThRkOKfLhypf66UJIrELMzpinwtAhZmHk
i6NNj4ftsejeey6jtzcJuY1bdSR6RexP4WByo+MBhywCeL0hmxxRxFE/mSSxpP2Q
ctmqeL149DcHW2/BxOH1DohcHpPm+67PkkrvWKJCWyjrklztZgan9GKE+bTvzn20
Q1DtqTWleMCwEWupaL86+mIQDNo3UTiDuIfyqGYiOeG8lCKGDXb4fu7hrqB7hbdg
eLD2PuJ58ycqFZe6K4edkT6XWnMMrQTYsznQp1wLnOw6Qp59t0gVbLQQHYXTzv/U
HO5TtyR3oZIErfvdxUvOCqAO4Ko8KIDJMs8Mf66WhLFDA3fiMGTqvvarrJTJk/vq
ul0cWjjrFJ0yK5GLVu3owyFYV82yFG0B2aPBpw+VU83YILy2ppOxJeixBbeEcoie
Z2vT+LyCEMuGSlPuCCqXyPazj+V55TFwG4cn8dmzuk5rFZ9uO1lrTKVqfyrenIs4
CLZw9HCHvyApyXaENL0rS14AGnVpDZ9330bWUrbZV2wAmbMB8gUO3Rz9CSmAzCJm
t2C9eCPYaa1vH13s/IS8WmKABipcRXZDCDjnlxB+l1+NQ4KfgdtrA3kJasidpf9u
OKSfwE4jzWTaUtuOEKRTig0bfntvi7JGcSnwEdc2qRvTyKHZ5Rvn8hC1dgsYE9dl
lPpnACNWYea/kmAFdOjnYcjNEQkOMiW2VBf4etMuvhimpOe4p7nnkE0DrbL4nIlk
KKWTBWv5MmwPXwHcuiESH/zOW1k3yNb21m84h0HUEym/gvY+nN4HI73+gdo8Fvr4
Ni5QwQPN+kwbHCq4vvuAAtWHsVLD0ALx+mKcShJpBYW5F17RXXDhhkJ/BfpPI7KB
ukIzNwwSr5eqZ1FJAUi80IUbmyRbhIhpkMcps7I7FKGElfjX7a6i1ASzlfR/A+6o
6BXlGuvG1xPT8LafqDtftk+g6CeH6FWXwG/3qMBhm3NkUnMtBhtekEX1bgeLKc/T
r8bNseV3cthusLH15Pb9XDQms3H3Cn9IJjiMyJUUwK3/aTmn0Gn9mCCNGpxncCbY
OSfzzlMS50rX7bSbzgn7oyPY25m4qyqeLXoAAofxgEoiVWj2eweItw+FWvz82wlo
nq/Rg4xI5ucfMx1X/YIv7DRKWv70TJesdepHFVjig5P5Y6DiBOSYZziESRdmM4lC
J8pdmphjRrP+XmPlB8UKPB/au8DMquXh4hEPP/tUaBgo97xTPhlVtT+ztl/BUYYt
kbwluOZnv9+CAIRAYYl/vdHQK/pFgWuwLGddAn91qAdU+jTfOL3xcwt91CHKnHWs
ljYgoTr3JJoh8ithbAf4u66d3LmtTWcriPb2FsmWSMYLcXU5XU8ouw73T4wxd+AK
6tMvNVuAoURKHzWL0A4qg0lx1CprJ1OxUrF9lrKR5eJNVyz+uBjSU0I5TOawbsaB
L0UOAnxxTNTuzM2B+CbrpTUJsO4T/hjK1JaCM4MyAgkRidduPDrUo725Zb122jzR
OuARyhRHSGXifzdGE/i9Rceno/ElvWQWj70M/z5rU8tzcuF9Tk2TOTB1k09wtifP
iqgMwA/aqnIvq1AStqRxIrC1p9xHa5B/plqWhIaK/Ql47qHO7DXO1cO7r9D64kpw
U2I12o1FEvd9HAkPB9OS8V6es3+r4VFLSBgT81eIkexBAA9tgd4i5euBkg7BsB5o
f8caHNji089OS7M+tzv2gqKp36qzQ+NYYA+u/rjI5ex6NCbUMlVw1ncgO76hM2xT
MWYHfyDEJP3v9MT3vFWPP9CwXxK4KhhMWINnLRPGs/XrNTfSlSuPPyI2/+A+qcJc
AtvuIXACgcWCkNUrFAPBP/sLJ/Dnwazp87Yd8eJFGBJ+mnJPdWdV7PcbittVM+nt
Ar8erOfny0fhiDX1zn8C8Bdl/OsKHCSi9jyobstbpGra1pVZsFr0WZJxdwG30yrI
+GFzF7sz/30PEpQ7qy4CSKPgkEpbyj/drEy26vdrsDonOEZGZI9WOWuX7saNoMmY
OQbigrFn1r+tv2JKw+/8vniHZUjskTTVDEpKXFO4sJrkFg5XYm4uPTwDb/pMwuIj
6TBcQxZRzLB25EFn4pccKit8o7lFAlfpnvrsiUD4ckGSigzA7sOUUTNqYP+XKbdu
aIfysljgbUs69UfmShXypJa+8S9Hiw3AQDMY+yEri/u+dIah6H1OS9q8wWZluPKW
dX17/CeUf3jtxo++5JAKz3MnizhBONZmATcDzIIYrf0DMww/HWmCyN+RAcF3RiUe
k9i0Zf9uAQ3oI7fVKGUKe+vR6J04p7AxRnr2zV1EG6wIf1uxq2uFCkwmrF5C94Mj
S/aDiX3scnsjQVmP2vN7goNhZ3DgCRjVwxj3MeYazgTPrfR916cskIiSIyWCBO9+
hU/nN59NElA4ajoFCt/Ny4XsJasjw/Xb6UhpYzGs+f8LBXJ4paH8fgthbl1oEfG7
1X4moRKfc7mV3wLwVkmT/4TgtdaUlw3a9Q0VPxRp5VXusSQSY2dI/9l9JcjF0w5L
tin/07lpGUzlbdmTy56OdY0ImwI6VT6ELkLO9hG5kYGPcMFDNOyeuzpKImw/MxP3
N12ZsslKdXsTyJm6SqVotrXOk+ogwf7SV0YOD90UekBWH82qNg3fAEjfw0UYeUfr
oCJEYRIn0OBttRLWMFSc0pTAjE88zmXafj6PfYq/0KAqcFPrZPjmYu7jtKPOl9ws
4C5/RYlUtQKsWJBKpJueHC0f2PGaTM9TBq7UVjPXdqk0Dnav0CTIunSVAtKaLFOV
yVVZbWET1Weu3wH6qRTO6PnjbEbhmw61fhzBuRpYnzxZx+eLEoP/edKJVDju6kCF
f9Svq0eIviAIzuLhJwdRJZO7gBcsll8J753TCnsXSgKbGcoqTj5tZmvLWDA807/i
JEv5RPpeLk4OxIMXkOZ9DH87Z5pRxq0AJtsTGDEAVODBw5XVUNy1mVUoZkErvgum
RCbtNFVWriVtIKU1K8nnrzoT1Dki4hqy59s82u4xg9QWiFzATDNccvxY7eMx6ayQ
B1+t1Wpmo7831iMKTU4e5PCH+IKz1V4G80LtgBDCaCWrB4rzvv6FDWMI6i8z7Ddb
pNGcLUTJE3eiqMvFX9WBGvGl8VoarYpjkbjXIDT/Rm5zwCXII0Css14gorl5qlTS
wfBQFMisCvZpCVRnhPpiOyJi+iqoyYmlVjgTGfj/fMJ55wYzhnhl8Ygk28hA+p9y
vAGF5smpnGENLc5Y1HaeXtqFQdzk6eVb4tsdMCxkHAW7jeOMJCbbQ19FLgxnrISm
PIVOxK7IUg1JtoUTBFa97ZsKBQxe+sh2z6WTJ6ZLaxtg+r2GQJ5OJyf7Xq1wds2y
C4lLJkjyfnNemxepNhjicLr9Xq2jlC1GOoWauHo0gj/asHbBCkChLd22udKmDZXT
xN/zKyclVgRq8HJEZ3fW7mQveSsM+3J3wGCdPn2XFXV6EiyE+dKKONcM9hPLNGL+
3y8KM+iay7sXmxZtKWmwDSsqhljGNCtzvl2Zo9qW1kZnOQY4zeJcldZ2hh8e2N7M
ZGaGsuFsxOpzHk+0zi+lZCC94+lIa4615wup3F8LDwMad1NXEezACLDsRMZU/1Zx
HZwqw10vxVyKC0rwHOLruEi6akLetk4F2O6Y1QtIT0eu65tF70GitHnV0KdKGQsr
f47I+aFMNoJFHKq+yhTKtWAQaQUobnRRK+5aXAsWdbEC3sILJr0xS4G1iJunNUrZ
tzDPid6IIe/fbJSCL7mgE1Q8Re6V6QREj3iWMXgdKON1QY4cXboKBZjGzMzyR6Bt
FFzthh0kddlhRpHb5a4yJnhxZdflBfX6dBQd4e/aMgXPi9Ea22ENCHh8JT2sDtXS
5z9+bwNesi6VDcM4apWcsSE+b80qBnaHT73ol8+kjeLg4Mh6xRCboFE1ooOQcBBZ
xpo5B1ogRh0+DhGrrxYV6iPNrB3OGJqxfy2Wd1ZBo3Xq07D/yXQaAz12E8WYfnqv
xKnHoaaA/Z/PsUoBdlsLkkU+YVbQF6aKYcNFzVNwEla1UW+2tjwSFtXyQA8gT+AQ
H1UKjC1G1T/ZdQs49s1WCWZr77XTtw1vs+RsDKxMEJFOIwIrQJ0jkbeVb/Gc43Dj
sxlSGPKmhwpwvLolDu2foNgxiOLjkcdBb27pi0I27xFbC+lDBO/Zy0JU3HGJ3loF
nl6tYqpye4e7OctotPVl7h95lc1NIG6FxkUS97pPK0rh6UgKfcSebltPItMtwzFp
xodhXIp+AvvFnpvE5oHiTCFZDm2+Sdrigph0Cbn24XoABeE1O9PBfrBXr/dGK7VV
Kx8kIK0Utmef939fmLivUXMKf636uO13gH2mQiE7/qcusETL67BCbUF27dN23XZm
XaFN5IGlB/b3+SpodFSn9AQG9A+N/GkCxf4e75XxDEe9lZBZQsTHTlYWODfq/ATK
47fW/HG6rZjvCi6Sr4v0PsNUdpU59S1wfazWV3j+WoApP24LGPdXSyoAbz4Bh01h
rlAodFqQYvINjrMbeYEHxTbdbwMbj7K5OnrQGgO5WaqsAz7rhlMeRD29x6FSEhOk
Pc9mV7C3EqsAbizwU169akHTFYtVsZaaCKoVGjsQOQetJPEkxlk+tkzuaRLMBR5c
h2Xn89hq9OmdcP3o4OXLwD80BFKKN4VybE1lUBSk8ySVZJumWOIWp99qeRJRnPIK
G9c2/tXjzLk9TLORWWq9DLVawWofhh9/pFvJuHxDwQ0RoOoGS7b9j+LEh1vDCRVA
17nLIxQrL6lGK2TIlKdOJ3X6xzM0cG8AL22i71lPCclSs7IrCwgpVAT6b9ozbAlJ
m1AiF/dyY7bJL2zNZdlVHrnCnViORvRT3WqtkQaT7/gO9w2WyHRRKcoeuFnQKBkb
b8zQ6FBtRdunr2GatCUafIDLrCssNRrEOo1lGTpiX/YNLL7/nIV49Qt6MiwltGFZ
E8piCxr68+eUtfNU2X9W/qXzXTVqoq7hClzjxZMxqkamv5qwlBZ60ALN2PNUUDS7
vluqsz218V03VWW0A8G4TRwElG/s1qiSpULQuuWrgBUuX3OkEj9ecgvGbDMfjuwE
b68x3OcaHTWRoQfG3JbHEm03XLCP3HjVAceKl146sOgt/g6HcspzvtuC+j4aGBTY
1+EWfI8mepEyNbgFjawh7zaORlsg7Q4mKcV/KB5OEacOv6T/b+5m6TfXm++L5Df7
787ZHcv78cWCVaXTdsyI7cvzFAltJZMCRUBfFW/MxOCmKBF8/aOZ2tjd79DD9JUu
rhPoIUTwpoa/WoBAUbEMFzQ3mCEr3YRXTXuBl5aXJ2urzDtJtW/AJ2TPOPJGVQ+N
O4Ym0obwT3oF3jwF3LULC4apYK3DioTb5tBkaI7kw48ovsGxTrOK4Jib8tHIUpFn
uB5+TppYsL7zQXQLiQctFrtxr324isbNw1hgSq6E+L/PPOG56wOuWnw3LC9t9XZ5
Rl7MXIXI5RWpzI5U4S6IkhEFtSKUsSWZIb3V4itBHTcX8kr78IwQy7gzZ9mam+CL
o1aQ6hwEfG1T3JCq3YEe1Swe2r4nQ7Be//bpbUbqJocyZnuWccqVCxE2uiRsMIdl
eweZ0tbBeoSnsoVY7WP0x4BBnnT7THBfayemFLokkhuUayySAXHZ/6Sc2q0A0CrT
MBpY83TrqUyCFaWhv0/Tm+7x2YeOVvBRtz84n13A2I2KjJXeIPw79RkfAD64AP1M
V+4L3TPRSvn7fWQNutbEHUN/dbaINof8W1aVbdaVfCio9pvaKoXV6j2232jRfY9g
/hslmoDqp35z3cg28hHC1ImeWMMRgW0VRTaQ/xT8HJA5o+Dy+Ab7wAS4iV41Ho/J
zGVEcrPGpLAxJPitwvkYXywtYUd6HoGHP/vpP+8TlPZiIUbaU8WYPTi77Btp71pl
ec8Ggm3FbmlPyow09pXqmcM3ZRhi4DRujNI2bgbTcw8bmBd9uDYQ1Z58b74MIMWz
NU6D0OojcaTCb1J2hXKIq+0peF6ziQIVvOU5Bi8oIiF9Dva/AVZh6Ofi0BGq3dnH
cJQH8k5sNJz03SYo1Keo/+CegGeCQtvQddJhVpAl9JDkIxc5shzaDfCbOaDdOcok
dO15RvYLpOSa4pp3njPLhB3n4s6gX2o40SfTvWPySw56B78jdak40IQ3eckPeEc2
IJ4tGUhWohbeqr5R7WathDcqkRJZteWl9h2Ke3ARrDL8C5ZWXy3aq9mD3VmuV4uZ
QifThhuprG7eede5NyEw0oqBHToN8VnaFJDvBGpKxpvwZXmTEc5h95SnVXwsZs02
C5pdlyIx2tqGMhoeqkwiBEHk5OoHmsQlWs1IjnF7faeed+EmKpKgkUrRuGx77Eyp
zhpWHIXZsaFGeSjn+O0Rxovbj2U44zTIxzX6/e15tXF2jfPneudpGGDIjjtNc4uu
MKyMULfPvqaCMc8XVb234xoRsFSPzy01xDAkDcCMWFPzw/khfxXD4n1KrzScmEGS
fTXWqg68tflCSPdzwDeM30VpEU7ffrnLWeSkQPq2XWxuFI5aYv/bfBtf1peDwyQq
16rHp9Agw/Q8vaF01VbPYs20zRXN5PC7USut1pCXZv2yKPLAcOF4rzy+zX9oyl++
gXSdl2qS0AHn82L3h8AdJ0jQjmofo3JoP4EgKpp9cOy3XDwEKjVYpv1vncqykvqf
7iUbatpeonB+6II6itXquDnxppVUk19nGAL3LHRVI/O0qUjTm5O+55DSh4vyTb1w
xz4DsXxhO9mVDstZxDtL+xByzqKmdv/qW91cx1clW4tJUN7MGMyIGQ+NFUq7v6Vs
BSbc8PurVlIvHNgxoyGlSi9CGWuBDnhAX3KkCL49BxTWpUWRwwDyEMb/HqD9W7B/
va1jXAUDuEEP2vtsDIv99mUMW1DRfDOluSjBU8NFPZqpZBTCS1HsMv67XPRMOKtI
Y7HH7kRqS4kcUeX2xbDFTBJ/TL+RrsGvo/PtvoBM29bYWwQmrKix6/1O2MNBdELF
CBE6uG68xefadkRUjS8x+4kr8IHaaev/kHdMjN8gGPgTkbxHfSU3OlpPQiM3ef/o
7qq59xq6pAYjuIBS+5Y62T1jgf2w+eKK9PJERUM9mk/w9ED8x/RfxZBDD+ojAP5W
fUByQmud+2dOfSUSHfX/fcgrQ8ya9U8rUdUoVN8EdU+SjVKVToohj5mEFXray9TP
fEQMQRVW50XYgkNnTOfCF5zrp1698KmHq0gbHAKP7FrqQKBmHBi5Qe+9KM/4Wdvh
hKwAFVTCRIX93ZYE5tEVGtBR2oSW1xD9dgtniTLgXMjJHcDHQjB5lkcI/q+CnVxl
C5TcW7i2tikIv2Ag2lpTux/Vey8tZftpIfFBRM8GgTol9x1NhzfmWBxBT8cF7agq
ztzWATigsz2lKM/2cSXD41pHp3LWgTUQlelCu1iPS2+SDTTzVuFESCXvCuKClRbB
hfLdm2zqZRl61Fq03FPkNExxTLpSugzPeD6C6mCDobaarj9i622yJl8thXOFAUTs
m0rvOvnZXtvf/vmmKs37t9Y+1ZDVEQJg3LA+EDZ/a4RdWv3I84f2D5tvwC9hwp8P
ftVDGjwCrS6uwgITPnaxYVaZCvwCYgdbnjA7/lb5OdOSh3et6nPPNWbFDCkXtPLU
InvLdQYku134RFCgcUj2fRfsoJzdKyRn+aty70c37mcVq9NxYGb+R7ZhPBEv+nJI
FVfWL6DpAWNVyfrEqnBOGj4oagSQWD3yRxeWR8XzVPmudUtkZ2MIZpcY6DH5U4VZ
GFstU7keNh7vyw9HUGkayMWHIFaUP5yg7t1d44u7Z37tDVycwlnZCAT2yFvr5VW1
GC9IfAXyEl9t7VnqFh5HnsXbm+37CbAts4WZ4lxQGQ5FimwevOFM2tEH0e9pjKWH
mvBfYLnNKB3LiotgjN0iL5XPfa0xoqoWjXt0Gz7FynSjCeWwJVVeosUMY4Op9r/3
BatmfKBtE8BRQOPlMLL3BLHH89J17DadKm/R8iwDp1A6rZx5I/gaezdwZupFaR1M
oTeMbZnWv1iey+FfuR57o/rjRrwhK7+EOroyQEB+f3nS/y9BwzcLBn8diUprEt/6
3e4wKXQGmcli+yQDFu/ezI+mShDqNwH8ybYGqfLPIn7ZDV2eONAbkN+r2C8uZ5O/
RkoO/Ko+60ZV+dEoQHJe4AUEGv72NvxXej8WSyAZdZk2dcWF1AGpz3aKkrUkgLNT
avAFcrlKypeC4qSLTgg0ZpuUPBZyK0hsNQsXipAzr8g1+SjGN9SnGj+hW/7xjfMD
dDDEumfov6xSOMFVZ9i5fQUnyS/PArlMbXibCelLXJl76q1b4HOLrnGdlwQCZkpg
ZvxLqEvTgm3th6oEeH9bRoz/q9k1p0nzwHMoUYkBVl76Q5IOz/gbKFHwdU5fCW99
H7MaVYtvg1fq+iIWZiWAgh/pqm2IQk60Tr5vW8HMV0Fu31ZXterA8IwzHM0bowTd
ByYD9uDQubnaAyoyqj8PBDM41TWjVFLdE4WGXPq+VYFnEVYVN6aNpY+XBwFS+636
Hc1vl8X6wbrOsR6mGwoPpPzHF/yXU9/OJ/xszJL/aXCKYpQNqYqzMhzSoglWRGhW
PsmRz8+dAQ88ru2QUELqKo+zDFztNu6Gl0cadrM2hJT+F7mQn6MqcCdJsAjDkyZc
ZIBqqA3+qE2YfXURhXAla2TXye1gbAlLqxmEd4Xgg5ckBn1V5HCFoSicgk8+bP1a
neT/B+5yYhXhxMfY8Bc21djFQikS6bmXxuH0bO57lXQnsO3wIfdo3COWkox65kDj
kuB2IGlXb0H8sW/7oK9rXMAIN0xgJb6oTZwkmT06ivCPED3iuKKUvoRfCprJ5vf2
IGRClrIblC/UH7cwqs0kOGsIaANcVxU4zUvJNxwnq6OO0GNlcUV82vslzK7ap4L1
lguXBFJWKp1Ry9edgD0l8WRYfWpRSMBTPY8kjDITdVLnezo8hitq9JkuEfwGtJ8z
iMv1+ViCG4Rn0qOV+FYIeWdtw+OdN1qiKcCMgLFYfBdJod8gBXUzhpmN3prOxgQZ
J6jCkirYZ9IimC5E/LlMrcujeBdZI6HmQsMWIRpHjpInst8Cmg/jZDCxKnMq7InC
5aBK4RahPfu421pfsiQkwdmIagHNL+ySf+T1U9F2axCRjfYsH/nNfxvdh4cmu78b
fgZ1yhrrADVPCXG5rxboLUE9X5NGDJO60GuuBXDQFj1Rv74ds0X13mdXGi68Ukj5
nc5jNHu1HTHgnaqkP2bdxV9S0ZYDre1fWZPqZD1GLg52VKeMbfG4nrE2DsKqcoTo
8xdbJxvXHgRrh7jk0tZzZCD/CRrIoufGE//oRfwGo28u7nfI+oq8YVEL2mGATV76
lwVRwp2lK+MoS1WpWG7/RGKXBi61KX+F9Gf5HoKnszKMH9tB3nnmNZnhmjVD8g7r
l5QuUkEWVAv6vBw97qmPf0plEuUA3bek8x8gIcrVdgwjFaVa//8911wFMJ9/mGG1
zSZif7QFj2NlIjR93b75ZyYbU/qpXNheivgpE3RBd1PmRPgvotFYiCDDiAkUX5qU
gEHiQcUmVUHRjjHpaMiprgg+csp75arVKCTCq/b80RX6d5HndWUdW1o0l4LZ1jUU
0uEHHEnQUXs4GL94Gm/jVTjpUsrJs/C5ILni0LPx6QUEo8+ytvFPquYzifRdsW6u
TT7lWem1LBWuCf3PL1Jcij5wspkAd6FnzuzPk9pTKynCJoaIMVNX+9+6WFfNGvNh
A0KqJAnLx+ii1tJIfhQcJZVoCGwugxWa7iu7d13pTfbeHWNKMi3kbFijj11hM1aQ
Uw0Ymee1Xk6JAiznlLfF3WtJLdTUdeT8Bf52A+8DVEu/xVf/o574/9Km4doTqyew
bpi0I5BAUTxNJfLB/EkQtmk8ZRLocJlNZPlVCu1b8GPLXwaRY4Y8B5wp7jpk7BWV
dRdRX1HF6D4p7MhcwsVCZQAsgyYIYKM1WkFB4Uxvo8SXRShDBgna9Wg4W+MKxnE3
QbV1XWmSxsdBn6Tn5QVcMo7gsia+TgNP70cVS8B0N2+O6yKk6Hnbn/JHyESMK6bt
oPkLTbR0pJEKjqGkfNJfmBRBqxFIlEzErm8IbqPEbKEh9Mwd7O89tWb67LHFpNlK
6J6yWYUhzzQx20dlmwshM/bOzmC3K42apb7dui2TYS/D3QTjpN20XeY7Y87sZwEF
7ArPBVb9wAu6BMrNc2le66ly4u+861wExyq7HG5xO+z+gYp4MOEJzTmWNO36pCBY
dI45+M7zL9q6q4sX2NMiA9XRJI+NjYvLPeMY7fT28sLrafHn/g0WglKfjTq7YYwc
f5eO9khz29jEa2RA6YGi6kyWFL+6vuQc/xOhBwLdusRTqaczZbd0OTuFtCtGEdvH
erRQbSoaMbh5OiGQ1BRW2Qq/Rtkv8xpO7ehT909m9f6d9AXIXzqv4hC5tbDtZzW9
rIjPcd9RpWyNcXATTkjknYQFkrRASg5jR8emZcCSMmsTmXjufteyGKpdg0Vc7jHP
22PPJ7xjH16xU+xHxRQs74dLIG39ALeBECEKjK78IUaiT1Q4ESeFojefORRrCAsM
jTogWjJBn3ZhabZGKQhsI0uN+/Z+QSSPGzsU2lfwriAwbnhuOdkMojvUOX6L07XH
D3nLI80drqnFIp3LrQykkZRkUVSafSWftMTYbsCkVoruKbFJhK3pRh1CZ74tEEJ8
QBB1fDU5NaiCSxhoATuSQVUoYA57GKd4WYj1ix+mBaa6KsskGYj2NaAszf9ThAPE
WEugT2sM6oYZTgbeldbG8iys0xFiP4eZT/Src1HW6qNdr5PEMBjdYAWj9Kz0jKUB
Rz9tNKkGgFzJG3zBkX3K+JeipJ3x77632Rlx1E35A+SWe3jlQC3ktrx6ltrtInCE
A3+Sd3WSx1HbnQq91oua+Hdk8avq5Qxbf1r3zFxFnLQ1rCn9LhN8nvKyygJ1MZPk
q663Kpwx44RBsLUR7uLrvDZRKDlECv31cmkrhMdUkH9AJCZucGCURDTik3jP11gF
Sh3dPRJH3hUWSBwH8DlmWf2kUNK7w0Z+g1LOvk9vyXQgRxTKhyh2wn1buaaYFQ6m
wjcwRlfzpKD4wjdZqO6fVxaZUPp6qBD9PjtwUaty4PKSaUIRCTzgj3IMRxFhEES6
42PIOwH50vYtzRYor6277R/wKFnMq2QfLwldSG9Tkkq97sn+gOZOQb+CuQ1OixuJ
8DXxaEb3h86yZoK9LtrzKZOVFfB2H4FYUJT0GAScZS1D96D5EGwIKOXg3c1doUGi
qrgO2psQJ8r6KSVRnRC4/8SiyY7TanmXxicHQdmK4wtNLx2kOwD/gwc+yZKsj+Tc
5PgOEyjamofe9lUsJnVffilNuL8XNjGKKvnfFx39V0sF/YQdad5wH5xK8zNoQdft
ll70GghA0v0sNZdqFu4lnYbPRexmMWCPeGh1iF1Sdl4MSi/OKi0LrAOXU847zRvR
Z5amGdI02WllL9eIGzfZs/i+DmFgWCdaAujzYPi+lMoi4qD1037jfkJpYXVbhKf/
drlnQldRBuUPL4JAt6/avpxXgoPG7wIaY0oMFZXOzjBNHI8kxyBF4b3issf+BMz2
BWycj9bl3EoWcnxe2APaF/+deHN2P32qAh7kW83ODJ8oLxeNeBSzdwThNE/q3b/o
gyMpsAbdDryVu0C/rohcVTRZfrA7iYhNjBhf/WRJfOxXi0Cx/I7GJQTL63Apy1nv
D3bKzzzf+abDqJyPk0Win3eBUU258q8/9BfeKRQ1lDtHtYH6/9+8Ie+KqNkhnXeF
+4YIGU4rIRPoo30ygYN3LWlZVnnTbrtGo5abRQMfwuNQKG20k9FvYXtQXntN4Ei3
sh2SSYJXn26ysPB8n1cCE8OcLPPxDIMeESYxHg6ibqCUMMLJOSVuWhSiPx79FK+6
I8JDKoCnyOIhvDhzhL1zr51Se5H1CK8RL0tjaR9JrlpO8X6t8oQrwyzExn7kJIbs
B1TtivEGJ9tgpNccZHMouiFiE5XCZrw3QEBhgIhi4QLJd7oxvWnini0nnpusUH7B
LZ931RgPnR44a7OUb0frjb812iJoburxqhALU93SfuKUITIYGijApp5cjLKB09nV
7mp21d3fP+FM/Y8M/PuB/2Lub+4dkD8z7d6IXD0hpncbXFZBbEpsbNPOOy60pG0k
dTQiESjTD8KXWxkomSuYRRQ4NYTfFW/wIEC8Yl+h0Mq09VDFYSM3++tNgfnCYTvL
UGNs/Czf90rVNrbO5hCBH7bp25IwWoQl9EmG89/KQoLGqGlX4ReuAGlChIq44HYw
JAbU+/Qx8QJSS99TcOZ4juelojy6EK3v8XU+afS9QGjVeVZMhFCxA3qBhzDTWKpW
1AAUwtOPOcKvWc3zq4FSRG8w3ihpgzVBzu/N9EqcEeRHtvbzagrEiwi6gE2Wmxgj
i7aQSKzpIGCo4Lo17N3w/F9v+Xy9+Vo8OXYzuJMGBemXFGbhDLrcNAxv6/at+kPM
EQk4A0QXwAyXEHxOKjBQFXjgwmVlb0486lXXlmNUoV6ISD2KAsK8MDn4hCgoKyu7
OX+vpc4S+aBwl+epv3fsLHm9C8l2O32wsODvVGzLyo/5EoL3dguIFTFkPaHhVC1R
BKtDRDi43pv4fL3Tz10AecsfebD0OLb+USVirlKLHHqwuSRZsIg43ioza9UZy7r7
1Y0gAMx4cWlpReGmaOAUpsaa/L70yCs+KO3z2WXcKiNEOEb/AZmyMHaWZ32k7aQf
5sXmfUsyFJgR+vzz/Ho+Yj+TW/dqqDXdqwsEnj29Y5yNoBi+Z2U1GDz3kApHG0Oz
Hk2jL3TAvSZlPJl1CChIHy2RWNaDcft2zUUSoQEyYNa1pI1tQxFtuHy3FzlOkgLI
ZR6j3A3/+2KUlWmMGE57Ua47iu+k8ktEbIM0l+aQRlgmhHrNkInQil8DShioK0Zi
nOpynevBAMjaugduPk7DmL7yYwozQ9UOi3ScH0yq52w7u91TgqSaZwt39fpBKLKi
J5B5bAewi3kyw+C1Th1cbsakTD5QAA8HnJCruth2yMPNKfl042BsVXw388SsAb3w
8AqHKs8P9ykgiT6e9DORA7/M+4R2Q1Il2RjUbCr7mlZXgtoUc9k61bVuKwJ/Y8Hc
2UWpYZMBErTLSHAGrMpet4LUyQV1aLMJI+Q9IJfZ35b68+DTgtli2AkkASSLH0dR
u4EqndcTF1AmGPcsDeIFxsvhQJFhA7OIblVNe52QD5u+iTkzhyIAbkVuRJSF2l5k
nWBc30z8/ebcv64VEPsr0MdkicELSpGtOB8sS6nZfl28hh1J1D0bX7Q1t2ZLacyE
Ta8OWn0XhAxe9DgeovPJBWKfFvNz8UPG0mhaRPZM4Do3fiaa99r380s6Jsm1Bcqt
bu3REoVSXklybnXKPk3Rnxzhd3ccXWHEW0JkldMu43a85rlB/UpuHsrnxY0Zkyla
r8VZj+uI7IobFiEnVwYkqK0eHofG70unCe5XCsmJQeynoh5C66rdAV9UE/qYQzvN
OFWcviNfYpN+oi0SPQRt4UN5HC6RD3i4yFYsTDNf7x0HrWb+lStd9w0Fu7QiNiXp
TaBFDX4VgGKmbUWCMm5KAeQbGBo2obG8ndNyIjU3HcbWZigPZLoDqa2AWSdrWF/U
+dZklYNaw3BPsFTZ3k9b+n0JO2ndVyZ7yj1JtWmJeoKwKAzVYqVfQHkAbhxemLKH
6D4AAKVDy0vnzA2kMauT1byPT89sBLs9PatHPLAAn0uqnj9zBW6NxDgIT6x8u40X
JgrWE20Qm8UUjCGRkzQ1AxFY4ivTWMnZqPpOcydGtsoZmQ/psekM1mTNqkWSDt7c
93bQGu3oHPlC+9PeY1Cey2LKRB9VndhyAjykJFG/zq3aNyZC7qBeKRXWjedShjUj
NSyHOyeS4HiOcgI5YmBidfNvBm2BqpAqrcgObe5hVg7cQjEmxELluTNp8hFpJclt
KpAWDqYPa8WP7xX6fGmmF38DrrZsINsIKpcw+Qjg7v8quxsUSoqwwBsVvWCEXYNK
JZrZem5hmKVUXwrcLDnYBjsZNHqQDB4fZjIZr800vEhT261PnxJhXZPAsYlV+wJq
a/zJJi+qW3CUjOQUKTpNeu+5pEwVzCmGG0FT3nlKt5v6u5v3oj0nhwurRG5VYPka
KNKV2Jsm6nNXvzpv8eYwtfjprVlVi037KgNY6HLRBQjXfSGwG03OqUp4RgPqvrZu
eobetMR9zq0PCav9194JrTBXN8Uuxh2Byn9gai3bJbjMfVmkZIJuCanS0OWnsWot
oXZTMPNGEFqetP0xzpLsOeMK99Df9hHiU2jfSbSQ0JEGj8KGLbYAKixn6LbcpcEU
kgmmAaQgC+M3Wh9hCaHQMo2sdcuJOMtyLEuogMtIh/H208FIhdo+foL9W+nB/YN9
cAXKkdw1Uy0+FbD3EEl0KrbKScv+Mu2G36R3kGpR2XHL5B/q2MF801LLj3rCBoft
NbVXiZKvm3tgxKD+pAz43wEjwaaDBjXpRZ5hyq53y8Ca3jaCBGwrtIWkSgx+fbyL
QGalQ7nP4zpyvgNZNtJ2Qn9K6hGlgewNowdNkxSfdbcSSQRIMSIqYV2giIQ4MqwL
DO+mcj36Qk/kGZR97mhFmYowShlpvHNORMoyb+o6+r8y4J6r+bW4vz4Nug873K41
jG8+u+pkfAZG6Oy2u9RLULKZaLH7XsjIqIbJ4tLOPztEOEZP11pLuZS3f3H7POJC
SowcBiSxxMuxwQt3J0nUeW0A0cY5Am1udiwEPFUiAmmbsmVeJBRG3nFNJWf/gIXX
NyaUAShEod8sk+gW00t7w+ct2RN8AkCSaQykIN/fab9m+tzi5dNMplX4roGv4+dL
W+NsTmU/Zo2LUzvi0SATPOXFRNskEZqYusIFfITFA73LFNPbR7UDBGAyh91i4Six
Gz23NIN6SEns/w9wJez+yKWQOBpvXdOC/MKiWjaFWAFDvFq8jU0TMycJmAbHt5Ht
ZKprWfcsiFGCyf2v9iZKrqlg6Zih9PsFnwNYr5ePqnoYQ9sfesMdZEC1B13wZi8i
tcpZ0QIWTzly93fNNZGFioh1I2knxxQEHUw8DLLB3fDd06qTjzSR3Ir+h7l8BoIP
lno5WO+sbLbQR+VM9ZopIo0iBYn9Aq0qxmqDvDkQBWdATi6slDVoZDNNn08VDFix
LnKIxD2ccuIjBoG11MYNPxtwZ2921qO5W8RFinQR+l+hIBzV3mmgayaOhPBMFM72
snbJQhkHa5JQpKHu4p0sPK4gfAAd0ptq4Om78s7AE4TTEYK6fQibBCm5+yuq87Ue
gPlABLHrIbzkyzqF6N8NDP6vc3q4fkM7XLSITSUwmPlxshDLXjCD5FLuWSYFrJxw
K/lzJVOhvYo5PfWgHySUgJPUgOcms3KSNWdP1OY3t9zx19Ion49lnYr1BaeXJ5dY
+ejWLv9d5QBIqlWiZwnR9X7Go4nqDfH3G9DES5+ouTJN/wzeABBJ0StQY6U1rYKo
9PQmL5eqSTcQoraBzAE00X3Usd3JDbVBSByCvBrZT0eTgbglPmugp/2XVK1xQLsU
peu3Icbq5da+H3ri2Qc0Lv7yJdcVszcuZ8nOEVKLGi57DW5WY6K6L38EAsAvz5YM
Ix4XmQyMqkqT8Dsf/hCc+bjv2y32SLdGhpwiRsZvkfY1IsP20kB8x0x+S9X/J7tx
DI0qJ5lVIUGZnjCSkkuMqY2XDPKlu3g4rSzlcYxYhX3xGBEouwdEmWf1FlxfhTUC
UX4gbyPULzI1NPCKt1QsHHw90hWQrfXj0NiGHuBXDz0hu7QY9JtpOA9eO1wnmbod
ZLkf9ooUQljv+hRp2QnpniZNmgNtWTihSiRZQ3ToFChGC7cDX3DL2ftOf3XOR/+d
i0VvM7mLvjxgKqRDLq0sITsGY61fiLYgXsab/ROCVl/0Z7ACzGoYPetK6qcjQWFB
hzV/Ob8TUAtqwOmVXCCuT1kUNlPsqWWZAUBQdU96Qusdj9mN95V4kQlKxs86m4qO
Fuw+TwLNDlXIbnBYySKRmq166NiIGWg+o14Nj5leCBiRRJf4RTk/ysQ6uyzqz0FT
kYIa2Q788sta15t1AKlXPX85FtHX1qeofx8oFH49HyxCjQVyDKbRP10Izo2Fx+TI
MeZ9NtMc1clUN8g2eGDcGwPMS1Q8pjLJ/sr6Gfca6opvTpy6/fbD+3lr6qjF7pgF
Ws68fhnfWa6rp6c5Pm512hbHyfM9xGr82M+ykVpaNTFa7D5YNY36S/AJ6D5dzmfb
GWEKTyIOwtPHqWtt2Gvti/WGmXWZODKfBD1jD6J+vxb3lyDPaSUK72ssBp0HFlDw
/oPSIJu8AgORJkiMuBbpoN648uTEIvsC64SSbqMcP9CmDZ4lbRX+DFjhjdOFUrit
JTMeqVZ++Czd2bjr9mvTAz3i0rU7LJ5dwlvXjX93hCamdnM907feXCofPQ0q5fYW
9DxapYD1F/MP+NXzbvUxU+4x/T0Dh4G1oMmu5DzNmK9ubz23YnhG3As6wC4bcfFg
svOKnF+64l1UN73vJ5SeGYyGKUbMzG8tcLRsYmlahiAirEg+rbXhy1nPIT67n/Up
1lP8vpgGwnTo/seGbCkM/Y0+rVSNDmQU9BRphqt1qUkgoSKw0B81UyM+o6DkCJOQ
gSn2HeYacY8awajzlM2E38KGdYqb6Ptl5IS7QKj4s5BQUB3X9aWZuy15dJN9ARAt
BGMFU03xFtxrXjZQaL9pSRvWxeNAvq8mI4ctaV8B2duhh9Hi2Q8igTZXEuKnCYQn
6oa5VdJP/OxTRl493YuyzEJBl7VSzeJYb5pK1bVaCKSQNJ7THCQaoVqGHjYV7ETL
UQhpNNTlqroRTWCfrLQ33nPCTe5vokRHnh0yWfjcwrQbR5jwDbDXFxb4acSrHKPR
20BzrpEi/ut5/22Kb9LPbnnGd9WomEkK6iaCbjOM8002FUcwh2iJJY+Af86cmcKg
UyZmF31Fy0Y49XIZM3wlbRcVfQa6ea0yvJ4PWjYaD7zkr+g9H2UHkxAUZoLRT/lB
bm1KPdgY/Az5s+tTNRV2ZVJRefEx3VPA0vqmcXCIIo5DB1sHbOEx3nCTxQXNlWF2
P9NKp0JuBc0SmJqwVjKpUIDpSDAK9eSYCS8omO3qSdoqFy2IffXzNWe8nsBngPrh
fww3iT791IlORIxn7q3vX4u9rthD8fsTd4+7ZXebJ9YddzucfK+ev9axCGTkiakO
haDJD/17/CnnYWDj+ErckYC6T729G1BpRFseeZLzsQUu2M/EUrvd0mK8CVT7JraF
JIjD6dCSqo8kHH3F98jPxqbOgiJJQ0F5ZFqaFfFr6IgvlsRCpv2KRoxEb2cYvGad
WUNMNHJCxPNSOCmjQ9kFIiB2Ssa5pi5dxnpJljp4+mjISegW27l4LH2+hzgSXlgo
/QREXQWHpLMG/L3sId6QTyXUVObEPIB6148C4D2KNmahBYOX9go6cgE7GKMc7ZfE
nZQLZ3Vcb4BEREPU9OlBoV/Jj5W3WAhF5pE7OD3bu+BgZX29vybzw+eW1/3/kOIG
iAavx2eeOeTE44dWZkfuyclHB5w77YI6uY3cA8Gsqh66fnsxYx06J4IOaEF7SdJj
Ld2CDzVCEaSe6YHN6SXtJL5GGfa1Ih4fNcetC5SZoJdUHSuI2KwO9As7yXUi5npH
lJVimofinHCqyyVpJ7iY+7KoWUgfGJ/GWcPq+W9eAfH8+wzZ64SIdFzfQJtBQZ0Y
ZG+R6ezaGeQzinrgUhlbws5svfuUaLGYkz6IK/sqbk36hDz+a0t4L4WTB/uI08GU
aKLNw8iM4Cbr2LLMHxNK2OfZPAwtXE1cX9ADain4oTDPNOkYn/R1zG32pBwZfXws
Cv2Jq32YKJHMyEGE7tCEahfdQtN8COCXO0pYyvYvVwCrbNpJVQoQsHVGEaAyQzSr
k/Ypbn8g4Txd6jW1h9LBmzteLmPbZDH/P6qy6Llpq79ruVTXtmM/qU9vV560aKHc
jyqcN8uvvEnG4//KEw+MWNZdzL5P3wkzpB/xMEejo5dpKe4cgI9/haBDg4fUisBu
s82eK5itaE0GepK8SbipasKV2PbCqY/X+QHB0pjiFAePZBMqliQtGFfFkNsbFhDj
1MF4oakujE02v6vumWRwIvV2jKtrBaphTJW+LxFuJGV827QLZozn1URP2+uqYJzZ
um2jBngpf+s3YXmksIXdrs6DuyAJwurZrGQfIzJlUyCYMLKG+7MFLxaimvFM7y7m
j3Wzya6yFJvTHGgwaSEY/Ogmgj7dCJBJD4+37dxZhtioS85dtW4PdUThD368JWbp
hDvP3IqKvv0eyFIFZgeMl9Orf+F1ueqAfctr8o9O1vz39BFLwfKokMisYI3tgmkg
hpa6nOIznA+zlyEyOmcrgyHA3bwez191OTOy69wRaCC0lEkB8BSPjnZYe+sbWIOj
qLPKexxGu3pTwSZdMIBP2nns0Nlqco2cmtRjHAKR0tRSvrEAhOpGwpamgTUtLrg3
ud+Ohe7R0EK3soXjUxIJTOfpQj7Vo88YG2F6SHSw9MaR6d3faCzWm+7sPhs5s9el
Cifpwby0PNst4qruaC0ogR8Yoz9KJOpzpH6MpbatW93ta5+uEtg+8llMIcOG1Xp5
dPyVKrrIb44MfRPKOs85DlTL3P7FVrB9ZbRS2Xo+lcAnLx98Lhj/mRrv9cxciZFl
9DJ9bWGh/Szk+w1ZiuWnO5mCAiQohDiUFXFLinEwrX/85Q/HqcfF6EOdtY9g5HDl
pCbk0BrRkMP01+5YOEAiFqRa0s9/nLC8SFOFtmQqzEfENUXiI7HGul3E542Za36A
kGqby8A7sBHknThvgopIKtx5jMTGTbD+JxV55ZKsO8Mw79VuL5AUaJDwnM3/fj7b
hkqsd7LPzqRzH3QZo6n6R5ZMciVNm5fbQVobwEc25iGyyogPkPz70ECqXRdo+hmy
HaPOtAJzoFESRbLJCeD+LXXZNCtaXNquk9EOX/pipQ2ZqsEsfeCO5FkwJrPQ0sBr
zzWonbLTaUDsxdZxwpeod+18xVl9oEZ/bRMEvIgHJlTJ3SczkXh/7RG1Ew2LtO8h
GtKTmYHLzt9R4uHGxOAkrVeavkA83VoTKN4KBb8VACnAqo6HNgho3MxozG9cTz+V
sdjyD/V6PiKRQZD6Il618dHYJDmGfjNzpMf+jZLLdC/wsOVw3xQxmra0YiCwntFc
+jtcJjc71qip97zQhQOoQ/lR4n3eY3MljG/61LoY2VKuin5TAdXtT25k6T3cEQjD
V/WP9btNV6lhaaeGPkT+wCXwCvBlOqE9xdmXRJicdWjxeC6NBBIFmNIX4+IpdRKw
l/7b6ONkWZDJg+y73lW7m3hZFwi+jaF0ihBYIWSlyaNUB8DrhDOwyuX2thzwSZ7Y
aQ7KFhAjVBpboRJHTGbnB/s2x4JUsNSeae6EuX0Jcq4A0NcUTQ2nYqEiHvQcwXhN
89DEYbL14oqhkI0nOe9LfxUOpuzThXkrtKW2vPY6u2L7RLLMsL49xJHt+81T4cxx
eF4QeYz3RDf5hEvPoUGaFbfTeqngXFsI8E65qb8yZmozA/x2ECdbudpiCukOOglD
cHO06QHWoEsWh4tVAbo20GQIzD5w17rgIUvtCtVQ3CaZo6usN6jTCtS+hqSTeSkt
9X9JTLijT4k+/BT6cBVMtl18ZZP6yGFngmSKLM8C9YPPBv7jC91veqkGRA+ovz6J
fQe+PbmSGrQQ4AyBAarq/Rs/6YADGR7uZa1IcHo9oJHM7pH/dhRk4oosdMzyOBU+
EDxh+3AdgrkKF6dZTAsKvBkvI1btqRu1w8efGCqf8qJbdsXJ/tr/oep48eyDZSxc
34ZbmnWAooHXs1E7iUws+KwnfAUuw8IdUamhLDW4QCdypqnfH62outBK8zLxf0Lv
izF6aI1QTUvYr/byiOqNVG17uhR5CyR9gtyeCpbkT6Tnk/hm1zrnV798FgTvO1NR
4DJSPB1vx7V4xuk5T4C9WtSZZFnosUWZbW7xAj6I9NxwXRuhslsqrbACJhzn0Ymm
Y4KOlcxoHAHEuVpUQY0rA49/iG9w0ffp4Z5LPZFczF38GmBG088F1QWgaalhl753
RWlDNW2xroUZZsRE2PurPwkBkJfVu9S0OJjcXWjm+IoNolmyRl/HQvC9erNn7XnL
XMUAeP0AunNE7HEWYdYH5YzBiOIrUkuPHpjpSHRP8YyZgPVwWkcMEhjcJqa77l8W
BASabf3TK8GZoPKa4Xv3XDBpDYUK2qWrOU3nFQQZenaHbTRM8RUTh5FwTmtyVGLZ
hhG7k5YJrmQVC6EJ0kJZR5/1wTaS4sPOEexKbW1GStDPXbG7IcbhE1Qb4HUb14mb
8d+wWHlQW6RXjGFpKqWOjGR/r9XmeprT3Gv6F0OTsR8VmUd9vJLwGyYLCJlNexbE
5YfHjUpCUWv8HojPXhtkUqDAuM88Gb7zHuQOiKe7VZwn0hrGtFXHap6BMhX/JQy2
CEmoyE1/0MyAxHrIWE6wMLson/tsW4R+BWOJC9dZyPXGB3kjHNajJW9yqb+scT2m
8Wuv8h74l6lWXjobe2xDDU++PLoLWkn9749y/+Q1izFDbiTHUqom9ofmDqVdfAxJ
CeEVFZOdQtDJL8MKd4GQLVGR3/sWb+Mo0Ffpcq4Pe/6K/tfqVHlmBRguyVm2eIF+
DGsdD7qFSoaQGjcEKZHbt5M4RyMj8ceJAE2Mwly0p93k9ddtUKaG3yc0e/3nCvCS
87P7fhJCVA2MBuD/uEZHIf8eHMlpR8MYw3chfcfwhflK195EQerjguPG8H3Ae+l0
gotgUgFfk5zqERSJUEx4QI29cOBUs70uKS75lv9VlbKPIFYKdRPH1U8V3Ryu/5qG
YlVjSOSfW+INJ9HvqTWC+fXkDYDW8ICprIw3G7hZQ9qkTjbDMRNu3Mm4YsuGKxHO
9r78imQmEnAIaHRYWFYDoXZfg55tUzLoli6FYYZofB1mU69vXAPgj2ulbZlahRIP
YLqAViu5YRpgRj/OgpwwRr7ygPt2CQnRGFgDM2TlY2pfsAfenXTMuwnutIBiK5hk
fqwBGY7CRvGlHxIwDhVqbvSOOPZnlEfUfnUPwn87at7PJvVEhnxKCszmJFiYG6+I
OOFYy9iqTPZXqamOioWZEGlOqISTXgYfYiiCHuloCo4bLHq4Nzoma2jHNKAnH5D7
6KG5Uv8oFpHmNxGLMIcEJMA9Iaw+X0ZBRMLDo3Z1B5xq+tqJa5sAC33JkXjGp7HL
11AEAHJPCQT4VYG+eEBqJODfghB5f1U2XK7bei4+/0buaEdRYIAlmlF6CoY1ZWxw
XDxl3st17+PzNq5+BLt+LxFSzCjLt58OA+puFpewGppevFIfSKwaLvUzFf8R1Sc6
haZyvdKt1m8xChWL98IOMaYu/1KU+o3Ec09vU0vj+7MynP/viCmIPBKeeZZea9Rx
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
h0h2SKtO7uq1whcsFy6mJfoMH5kXK2PHyYL1jvEbLov2qJ7Rl1n3Ifwa3a1rDOb2
rqLYhY5ycbs1fV08WEq495jCBiS9s8heDCFDxm8WvEb4pNGiPTvGgrADWcX749EP
8cOppxE4FTouafHwYN+0R4iPaM4T9YkoOm0sq9W6khM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 95136     )
8OlG2n5hoSKfpsjfN74CSVuq8I6SRydnym/Xm3trzDHLGBVFzpaxSoyccWH42mdE
vazlzj3Id/TIt0rSCQjjotSdD+8mrXh6Rv73+FXC2z2k/50JNTr1bHhmQqLPZnl3
`pragma protect end_protected
