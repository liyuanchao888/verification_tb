`ifndef GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_BASE_SV
`define GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_BASE_SV

// typedefs

typedef class svt_axi_ace_master_base_sequence;
typedef class svt_axi_ace_master_base_virtual_sequence;
typedef class svt_axi_system_base_sequence;
typedef class svt_axi_system_sequencer; 
typedef class svt_axi_basic_writeback_full_cacheline;
typedef class svt_axi_basic_writeclean_full_cacheline;
typedef class svt_axi_cacheline_initialization;
typedef class svt_axi_cacheline_invalidation;

// ================================================================================
//************************ START OF ACE NON-VIRTUAL SEQUENCES **********************          

// =============================================================================
// =============================================================================
/**
  * Generic sequence that can be used to generate transactions of all types on
  * a master sequencer.  All controls are provided in the base class
  * svt_axi_ace_master_base_sequence. Please refer documentation of
  * svt_axi_ace_master_base_sequence for controls provided.  This class only
  * adds constraints to make sure that it can be directly used in a testcase
  * outside of a virtual sequence.
  */
class svt_axi_ace_master_generic_sequence extends svt_axi_ace_master_base_sequence;

  constraint reasonable_use_directed_addr {
    use_directed_addr == 0;
  }

  `svt_xvm_declare_p_sequencer(svt_axi_master_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_generic_sequence)

  virtual task pre_body();
    super.pre_body();
  endtask

  function new(string name="svt_axi_ace_master_generic_sequence");
    super.new(name);
    bypass_parent_virtual_seq_check = 1;
    wait_for_all_xacts_completion = 1;
  endfunction

endclass
//---------------------------------------------------------------------------------
/**
 * Base class from which all the ACE non-virtual sequences are extended. This
 * class is the base class for sequences that run on multiple master
 * sequencers. In addition to being extended to create new sequences, this
 * sequence is also called within some virtual sequences like
 * svt_axi_cacheline_initialization and svt_axi_cacheline_invalidation. This
 * sequence cannot be used as is, but must be called from within a virtual
 * sequence that is extended from svt_axi_ace_master_base_virtual_sequence.
 */ 
class svt_axi_ace_master_base_sequence extends svt_axi_master_base_sequence;

  /**
    * Enum to represent the relationship between addresses
    * of two consecutive transactions in this sequence
    */
  typedef enum {
    SEQUENTIAL_ADDR_MODE = 0,
    RANDOM_ADDR_MODE = 1
  } addr_mode_enum;

  typedef bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;

  
  /** variable for selecting domain */
  bit generate_only_shareable_domain;

  /** Sequence length in used to constrain the sequence length in sub-sequences */
  rand int unsigned sequence_length;

  /** Configuration of sequencer attached to this sequence */ 
  svt_axi_port_configuration port_cfg; 

  /** 
    * Indicates that the addresses provided in directed_addr_mailbox should be used
    * for the transactions generated by this sequence
    */
  rand bit use_directed_addr = 1;

  /**
    * Indicates the relationship of the address of one transaction to another
    * - SEQUENTIAL_ADDR_MODE: Address for the next transaction is incremeted such
    * that the next cache line is targetted. All transactions generated will be
    * one cacheline size transaction. The address of the first transaction is
    * defined by start_addr. end_addr does not have any implication in this addr_mode
    * - RANDOM_ADDR_MODE: Address for the next transaction has no relationship to
    * that of previous transaction. All transcations will have addresses within
    * start_addr and end_addr.
    * .
    */
  addr_mode_enum addr_mode = RANDOM_ADDR_MODE;

  /**
    * The start address for the address range for transactions generated by this
    * sequence. Applicable when use_directed_addr is set to 0.
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr = 0;

  /**
    * The end address for the address range for transactions generated by this
    * sequence. Applicable only when addr_mode is set to RANDOM_ADDR_MODE and
    * use_directed_addr is set to 0.
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr = (1 << `SVT_AXI_MAX_ADDR_WIDTH)-1;

  /**
    * If set, waits until all transactions complete before exiting body of sequence
    */
  bit wait_for_all_xacts_completion = 0; 

  /**
    * Indicates if a transaction which is not constrained by protocol to be of cache
    * line size (READONCE and WRITEUNIQUE) should be constrained to be of cache line
    * size
    */
  bit force_to_cache_line_size = 0;

  /**
    * Applicable if use_directed_addr is set.
    * A mailbox into which a user can put addresses to which transactions have to be
    * generated. The sequence times out after the delay sepcified by #direct_addr_timeout 
    * if no addresses are available in the mailbox for generating the required number of
    * transactions
    */
  mailbox #(addr_t) directed_addr_mailbox;
  
  /**
    * Applicable if use_directed_addr is set.  A timeout based on which the
    * sequence that waits for a directed address in directed_addr_mailbox times
    * out
    */
  real direct_addr_timeout =1000;

  /**
    * A mailbox into which a reference of transactions generated by this sequence are put.
    * This can potentially be used by another process to take these transactions out
    * and use its parameters (such as address) for controlling another sequence or
    * populating another sequence's #directed_addr_mailbox
    */
  mailbox #(svt_axi_master_transaction) output_xact_mailbox;

  /**
    * If set, initializes cachelines of caches of peer master for the address
    * of the transaction generated This is done before the transaction is sent
    * out. For a description of how cache initialization is done refer
    * documentation of svt_axi_cacheline_initialization
    */
  bit initialize_cachelines = 0;

  /**
    * Indicates if the value set in directed_barrier_type is to be used for all the 
    * transactions generated by this sequence
    */
  bit use_directed_barrier_type = 0;

 /**
   * The barrier type of normal transactions for all transactions of
   * this sequence if #use_directed_barrier_type is set. 
   * The specification recommends that by default all transactions are affected by barriers
   */
  svt_axi_transaction::barrier_type_enum directed_barrier_type = svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER;

  /**
    * Indicates if the value set in directed_domain_type is to be used for all the 
    * transactions generated by this sequence
    */
  bit use_directed_domain_type = 0;

  /**
    * Indicates if transactions should be sent in blocking mode. Only
    * one transaction will be sent at a time. Next transaction will be
    * sent only after previous transaction ends. If cacheline initialisation
    * is performed, this parameter is not applicable for transactions generated
    * as part of cacheline initialisation
    */
  bit use_blocking_mode = 0;

  /**
    * Enables atomic_type=EXCLUSIVE generation.
    * If unset, atomic_type of all transactions are NORMAL
    * If set, atomic_type of transactions could be NORMAL or EXCLUSIVE
    */
  bit exclusive_access_enable = 0;

  /** An event which is triggered when cacheline initialization is complete for
   * all the addresses of the transactions that will be sent from this sequence 
    */
  event cacheline_init_done;
 
  /**
    * The domain type used for all transactions in this sequence if
    * #use_directed_domain_type is set
    */
  svt_axi_transaction::xact_shareability_domain_enum directed_domain_type = svt_axi_transaction::INNERSHAREABLE;

  /** 
    * If this bit is set, the sequence will initialiaze all cachelines and will wait
    * for resume_xact_transmission to be set to 1 before sending the transactions for
    * which cachelines were initialized
    */
  bit suspend_xact_transmission_post_initialization = 0;

  /**
    * If suspend_xact_transmission_post_initialization is set, the sequence will initialize
    * all cachelines and wait for this bit to be set before sending the transactions for
    * which cachelines were initialized.
    */
  bit resume_xact_transmission = 0;

  /** When set, a check that ensures that this sequence is called from
    * a parent sequence of type svt_axi_ace_master_base_virtual_sequence
    * is bypassed. The check is required when cache initialisation is required
    * since cache initialisation requires acces to a parent sequence of type
    * svt_axi_ace_master_base_virtual_sequence. 
    * This should be set only when cache initialisation is not required.
    */
  bit bypass_parent_virtual_seq_check = 0;

  /** Distribution weight for generation of READNOSNOOP transactions */
  int readnosnoop_wt = 0;

  /** Distribution weight for generation of READONCE transactions */
  int readonce_wt = 0;

  /** Distribution weight for generation of READCLEAN transactions */
  int readclean_wt = 0;

  /** Distribution weight for generation of READNOTSHAREDDIRTY transactions */
  int readnotshareddirty_wt = 0;

  /** Distribution weight for generation of READSHARED transactions */
  int readshared_wt = 0;

  /** Distribution weight for generation of READUNIQUE transactions */
  int readunique_wt = 0;

  /** Distribution weight for generation of CLEANUNIQUE transactions */
  int cleanunique_wt = 0;

  /** Distribution weight for generation of CLEANSHARED transactions */
  int cleanshared_wt = 0;
  
  /** Distribution weight for generation of CLEANSHAREDPERSIST transactions */
  int cleansharedpersist_wt = 0;

  /** Distribution weight for generation of CLEANINVALID transactions */
  int cleaninvalid_wt = 0;

  /** Distribution weight for generation of MAKEUNIQUE transactions */
  int makeunique_wt = 0;

  /** Distribution weight for generation of MAKEINVALID transactions */
  int makeinvalid_wt = 0;

  /** Distribution weight for generation of WRITENOSNOOP transactions */
  int writenosnoop_wt = 0;

  /** Distribution weight for generation of WRITEUNIQUE transactions */
  int writeunique_wt = 0;

  /** Distribution weight for generation of WRITELINEUNIQUE transactions */
  int writelineunique_wt = 0;

`ifdef SVT_ACE5_ENABLE
   /** Distribution weight for generation of WRITEUNIQUEPTLSTASH transactions */
  int writeuniqueptlstash_wt = 0;

 /** Distribution weight for generation of WRITEUNIQUEFULLSTASH transactions */
  int writeuniquefullstash_wt = 0;

 /** Distribution weight for generation of stashonceunique transactions */
  int stashonceunique_wt = 0;

 /** Distribution weight for generation of stashonceshared transactions */
  int stashonceshared_wt = 0;
`endif

 /** Distribution weight for generation of WRITEBACK transactions */
  int writeback_wt = 0;

  /** Distribution weight for generation of WRITECLEAN transactions */
  int writeclean_wt = 0;

  /** Distribution weight for generation of EVICT transactions */
  int evict_wt = 0;

  /** Distribution weight for generation of WRITEEVICT transactions */
  int writeevict_wt = 0;

  /** Distribution weight for generation of READONCECLEANINVALID transactions */
  int readoncecleaninvalid_wt = 0;
  
  /** Distribution weight for generation of READONCEMAKEINVALID transactions */
  int readoncemakeinvalid_wt = 0;  

  /** Distribution weight for generation of WRITE transactions */
  int write_wt = 0;

  /** Distribution weight for generation of READ transactions */
  int read_wt = 0;
  
  /** Parent sequence of this sequence */
  svt_axi_ace_master_base_virtual_sequence parent_sequence;

  /** Active transaction queue */
  local svt_axi_master_transaction active_xacts[$];

  local int log_base_2_cache_line_size;

  local int log_base_2_data_width_in_bytes;
  local bit seq_initiallization_done = 0;

  /** Indicates if start_addr has been passed through uvm_config_db, or is directly set */
  bit status_start_addr = 0;

  
  `svt_xvm_declare_p_sequencer(svt_axi_master_sequencer)
  
  `svt_xvm_object_utils(svt_axi_ace_master_base_sequence)

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length <= 10000;
  }

  extern function new(string name="svt_axi_ace_master_base_sequence");

  extern virtual task pre_body();

  extern virtual task body();

  /** updates parameters needed for sequence. This includes port configuration
    * handle updates etc.
    */
  extern virtual task initiallize();

  /** Generates transactions based on sequence_length: 
   * If use_directed_addr is set, the directed address is fetched from the
   * direct_addr_mailbox. 
   * A callback, pre_master_base_seq_item_randomize is issued where a user can
   * potentially provide a transaction. If the callback returns with a valid
   * transaction, it is sent out. Otherwise a transaction is randomized and sent
   * out.
   * If the initialize_cachelines property is set, an event is triggered in the parent
   * sequence so that the cachelines get initialized. Note that this needs to be
   * done in a parent (virtual) sequence because initialization of cachelines
   * involve multiple master sequencers. Once initialization is done the
   * transaction is sent out 
   */
  extern virtual task generate_transactions();

  /** Randomizes a single transaction based on the weights assigned.  If
   * randomized_with_directed_addr is set, the transaction is randomized with
   * the address specified in directed_addr
   */
  extern task randomize_xact(svt_axi_master_transaction master_xact,
                      bit randomize_with_directed_addr, 
                      bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] directed_addr,
                      output bit req_success);

  /**
    * Gets addresses from directed_addr_mailbox. If an address is not already
    * available, this task waits for direct_addr_timeout before timing out.
    * Once the address is received, we check if it is feasible to send out a
    * transaction with that address based on the weights of transaction types
    * and the corresponding domain type for that address mentioned in the system
    * configuration
    */
  extern task get_directed_addr(
                         int xact_num,
                         output bit is_error,
                         output bit randomize_with_directed_addr, 
                         output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] directed_addr 
                         );

  /** Returns 1 if any non-cacheline size transaction is enabled, else returns 0*/
  extern function bit non_cacheline_size_xact_enabled();

  /** Checks if there is atleast one transaction that can be generated with the
   * given domain_type based on the weights that are assigned.
   */
  extern function bit check_xact_weights_for_domain_type(int domain_type);

  /** Sets the weights of all transaction types to 0 */ 
  extern function void disable_all_weights();

  /** Checks if the weight of atleast one transaction type is set */
  extern function bit is_any_xact_type_enabled();
  
  /** Checks if any non shreable transaction type is enabled based on weights */
  extern function bit is_non_shareable_xact_type_enabled();
  
  /** Checks if any shareable transaction type is enabled based on weights */
  extern function bit is_shareable_xact_type_enabled();

  /** Waits until all transactions in active_xacts queue have ended */
  extern virtual task wait_for_active_xacts_to_end();

  // Task that derived classes can override. Called just before an
  // item is sent. If derived class implementation passes master_xact as non-null,
  // that item is sent.
  extern virtual task pre_master_base_seq_item_randomize(bit is_valid_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] my_addr, output svt_axi_master_transaction master_xact);

  /** Assigns a weight of 1 for the transaction type given in master_xact_type */
  extern function void assign_xact_weights (svt_axi_transaction::coherent_xact_type_enum master_xact_type);
  
  /** Gets handle of the cache in the corresponding agent */
  extern function svt_axi_cache get_cache();

  /** 
    * Initializes cacheline via backdoor access 
    * @param addr The address that needs to be initialized via backdoor
    * @param is_unique The shared status to be stored in the cache line. If the
    * value passed is -1, the status of the line is not changed/updated.
    * @param is_clean  The clean status to be stored in the cache line. If the
    * value passed is -1, the status of the line is not changed/updated.
    */
  extern function void initialize_cache_via_backdoor(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, int is_unique, int is_clean);

endclass: svt_axi_ace_master_base_sequence 

/**
 * This is a virtual sequence and is the base class for other virtual sequences
 * in the sequence library.  The sequence spawns off a thread that waits on an
 * event before it starts a sequence to initialize cachelines of peer masters. 
 */

class svt_axi_ace_master_base_virtual_sequence extends svt_axi_system_base_sequence;

  /** The parent of this class, if it is of a type derived from svt_axi_ace_master_base_virtual_sequence */
  svt_axi_ace_master_base_virtual_sequence  my_parent;

  /** Cacheline initialization sequence */
  svt_axi_cacheline_initialization cacheline_init_seq; 
  
  /* System configuration obtained from the sequencer */
  svt_axi_system_configuration cfg;
  
  /* An event which when triggered starts the cacheline initialization sequence */
  `protected
7?Z1JHW>e16W8OJ\C5/]1=PP>J0M0f&::6aJ:E/I>A8^Z-T,>\B04),-0Q84JEM[
3(V0_#@Z5GQN49]H4JcH#9)g.4cNd5[LZBQVB,gBQUOdf<[L4(]&7-IZ_1IG8NRgW$
`endprotected



  /* A semaphore to control access to the cacheline initialization sequence */
  static semaphore cacheline_init_sema = new(1);
  
  /* An event which is triggered when the cacheline initialization sequence is done */
  event ev_cacheline_init_done;

  /** An array of ACE ports in the system */
  int ace_ports[$];
  
  /** An array of ACE-lite ports in the system */
  int ace_lite_ports[$];
    
  /** 
    * Indicates if cache invalidation during cache initialisation should be bypassed 
    * The initialisation sequence sends MAKEUNIQUE transactions followed by READSHARED
    * transactions from peer ports. It then invalidates some random cachelines. This
    * invalidation can be bypassed, if this bit is set 
    */
  int bypass_invalidation = 0;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_base_virtual_sequence)

  extern function new(string name="svt_axi_ace_master_base_virtual_sequence");

  /** 
    * Gets system configuration from sequencer.
    */
  extern virtual task pre_body();

  extern virtual task body();

  /** Utility to print caches of all masters */
  extern function void print_caches();
    
  /** Populates ace_ports and ace_lite_ports arrays using system configuration */
  extern function void pre_randomize();
     
  /** Utility to find all ACE and ACE-lite ports in the system */
  extern function void find_ace_ports(svt_axi_system_configuration cfg);

  /** 
    * Gets random ports in the given domain. If a value of 0 is passed for
    * num_ports, all the ports in the given domain are returned. If
    * port1_in_domain is set to a value other than than -1, then the domain
    * chosen will be such that port1_in_domain is part of that domain.
    */
  extern function bit get_random_ports_in_domain(svt_axi_transaction::xact_shareability_domain_enum domain,
                                          int num_ports, 
                                          int is_dvm_enabled,
                                          bit is_only_ace,
                                          output int ports_in_domain[$],
                                          input int port1_in_domain = -1);

  /** Gets cache status of the given address in the master specified by port_id */
  extern function bit get_cache_status(int port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, output bit is_unique, output bit is_clean);

  /** Function that puts back semaphores. Typically called during reset */
  extern function void clear_semaphores();

endclass: svt_axi_ace_master_base_virtual_sequence 

/**
Utility methods definition of svt_axi_ace_master_sequence_collection class
*/

//vcs_vip_protect


`protected
NS]eK6R2JJ9\\EVc]e.R:@JW0&P5YLE8=Q-HF\J,5OaD)ZbY<U7<1(P5P3N:<]f\
g4./TOd/A^0Ce?[gG&?a=1gCFS670U#SWDH9)4/Oc47K,bf#DF2>Bcg@]^6XX=08
VLYAM9LVFP1]BB]?V[cA9[G3GB-XZR^@<(4SSc_QT#0eY]b2<RN0)/N&)+^PX=gF
,:Ka6gSCL28QKRR_R[+&g(d,#6:PMN/fD.^99A=0<bc[0^;\W?@Eef#R3c67Y^[D
^69Xa2UR_ZZGT?11c@J<H-KV;2c9E&CMVD)HI1=9W/6C.9=Ub^Y]3MR:0Y/OU12#
6Ja+32LYW2g0=;+89U9e;baa:W[eP?\,G3Y,>>_)B2<D=WY&/N?4)OeY-U;Jfb/E
b0BX[0AO5RDc+d/C;A+N3/#PAd>SX2]P_54[;V_YI[fP2H5/KICe6a\[&4d9>M^<
WHV5F5JAOO1\VPd<-60@1M:QIGX&\,CNYPR:LZ<-W&B\B]&=))S&=X0//1,DH&PR
f:#</D^X\@_\SME.d#&/]JM>a[1_V_D5#N[O4\J;X3ReO7fE6WNb4+C9T)3,Uf4E
/d2b[8=&#\AAASc>_BVM(#<Le_YOUa^P-[R4&(dI,Ebf@e)PD7E.=6>J2H7FA9dR
IY@,3]K]S>52Ad6IPX9fa9/7&JJ8LB,;1#^?bZ::Ud3)Y:G14@N\Q)=QPUQcX;71
G>RPJS<C]LC(gc:2f,8YKG[J<c9]7?+OZUWV5.AZL4S?I&=(U/?,CN:G<^<f)724
g_=>Xfff4;g(QRFN_IQgcFC4>9-[dIX?[73OVEBV&H\7;3Bc.3<4,9gP35^b&f;Y
J-U(VN\A)M_#5fEDAKCST#I)Q<DbF^Z58FROW3#:ZZ;#C0+\dV5/BIaX0#(.EX45
Pf=Xb=#0-C0J,>Dd/U3TR9)9MHBD+DTAW>RH>a0Y]A4eV+VaD+Y3JTe+8LZTW(eI
KYMYIbLMB&B=/SOH@YEF^<TV@LRc]4dBU9DC5I_J\\+@f0TTUGWMS]F:QZN.7Q^V
3U^<Uc7g\+@Of?8KMWP1:L[=A+cF6JUc9dD+]c=C]-XO8X_=6?\HDZ=R90+1a1d^
a0>/M=U;JS&XC1@1ZKK(=c#_ZbN+R4Y9>MLGFS/dLEDg<Z92<HdAD^WBZP@C/Ae5
#=EYG(N>J>@B2NU2EF8PDND09[1Vg4VGEICb&PEJNYMe[6e0RGL>Ke0E:,7Xb.JJ
W?,(a+/1USeQc=D>3#b.eOE[)A3gBU=MJZ1V>daKNY2FBE3e8eIdJ-0;9>4:Rb#>
.6H6Dc(XY+PIBM^Q1DX#O>6QL+-)YY)=RLbK+T@CJAC<4DWCcUS-8S5Y/Y(b9_<1
M(R3DL(@@&?PY<&^L@P[R+(3TLPZA0_6E>fM@ee1UHA.TUUI0RH[F?@@6SKAg)dX
V?=f&/7agK46,9PfZN9W_#SD-fBQS6-FAC.P;eAKNP^X_1IV40(8[B>Yega98fPI
GfME6b\+_?U7]CZb)/N61[<-f\IFB3<]YTN-Xa(\[Y^-6Q^J,YdSVS6((g+3UI6[
d@F8AL[E7I7:3(>?Md_YfEAKRBYON]LGO4H0\4gM)\^^#,\FT0Ee<)W7N9e<JK,W
+H.ZAS2c5D:B#AA>:EX].B#eJbWeBVSA5EWGZP4[FG)2->g>AY8<8T&A+?/H/+=U
A@?g]WH;fdJ.A5VXVeCfZ,LD,H#;SYB=]XL9DF1-O4ANeVfY9;cdc<0X<@O8da\a
I]DI_9N0YLM,Qc2\9gfJG<[XLgXRg[Q[L>JAO_K4a[/3@c2f-QSdcW3-DX>E0J<B
-NL1;-&^fM&E&WQ?&T[OYV;TXWMWLI;(DWe/+#K<AUS\WJN0V0;?@V&Z\DS2e.(#
dFDWHU1fI>E<4OH:09A:QF0Qb<EQ1.9?C#]0M9@@beUEBB9Yc70S;FLV/<K01,@=
VBPF<XG&GZ_L_Gc5g_Q=[IW]338.@E/^[OfS49(]<Y4U+)SR>c0)[5[#EVJFd8-5
=&@MK3T[+=K</cH9VdQEDG;_K6RWNP65Z;;6#KX34&J-K]1JC.[]QYeT&@27]W#I
+;-BOFgUHKQLT[>URT5]8-TEZd6e.212#0Z?9M]L-\?_FIJ9aN<#&L(;,/@e&H\7
?WQNU^Z@84,+0<dD+?KV_Nc^,?&a7c>5Tf2>44]);YPb[?(I-GKD6gDaQS]33&@C
P&YaUPZ82:6@R-1+)\EQCaTJ]JQ:<?V9Qc1cCG6Fc.]L.Y[1M.WLgZ+S4Zc3,6+[
A8-\4UJ]QJARLg.52@,a^=1U<+/:JI5TA:a<TQR,_XfHOF>cT88RZSR=bR^\<+AM
;e[7H645Z5K#>W58.JD7VGc-JEL?[7Ue<gc(E^-.H:Fe8_15X>C0K(5OF#O,7TXL
:A525#X.SCMA01(V<2LD<E.X+^I7f([F@;f>[G(VZ\E)QbSM/(ZFfF8HceXEdCd1
dA]T@]UR.IW\cQRB3C=\XV0C4^,ZbH@6_#TPZAGK<G9K3gYA9K7[<8V28a?J7O2K
ZY06;P/;@C;LL(M)G.06GH/G&K<M5<.ZEP;?79>WU)H+-3?Y&H,d9/XaL.7@6eRU
<D[:NcSOVMCa@&.-,JX143;P_E@-]b34;=YYYe6L\5Qb0ICEU?<YE0JYZQZW05N-
D8K^UcCY/;)#47f4-U/@YS801&Q924O)6-?5WXTfM85@>.&(0]&11K6ODFD2XQE_
-]0I/?NcKAc,JE]BOXXQ3Ke6bPQ.@II4#J6Hf+5V:<>[XW;,9+g-d)?O98NEdf)&
[9-;<H9P];MdE/8a/E(H)I(12:HCgDUHZ9f3<_\9X_?.OO1+Sa5U:0[(80.D,b&N
#I1BC^,_A#U6T#GD@XVbaI>^LT>5C9B)H-\<-,dK@_2(Ye8]Xd2#11A^RdHXP2A=
G1e6?<\O/G,,;Bf;T:I00<6c5OBf7D7Og.>_d\\)0^-AH^X]#gR&7V)7ac-R6C4Q
Le#M_KYX[d;HAA-\dR7I7TfM+ZEU+1bDW@BS6bXLTR>5MDGM/9E4AcRFe#CB(&6+
5I).JYf.eR\CC9F1\)4OLd66WXT;L6_,g?/43fa)f/&1M13.=Y3?&Uce^S5_HJQH
HL.Q]QaKIE?B,;bYZK,#5TfMJaOV=NcF7FAN:cX]a&;9X;(HIc,IcF][,/>fR8@,
OLeTHH:UE>BX38UDgWC,K;MJ1XUY9:T1--H/>2M5c-[4<Jc?3S7RR:3D&4XE2bKY
NR8/GZ5agf5]=2><>DI=VgbW48]OVE\@=D)d9MIU@1;)6W+[@HaV5;/:A8-MY7WW
e5QHcRd]5Z5\W&&1+gUT5T3_d(+&?(E?0UE]JFMSSSYV;JNK-L6(GA?eTX,fR_fe
3K9.K6D5C-S3A@W(5YV)<ANJTf\=0AKX\,H+a1CV7NNgNd@73WBT8,:-6HM1K\VW
6\1gb/[U,L-?3AZYJ(We/T+Baf6-cM3SEC+1-.JI5:FR.Nf9eZ_XJCPI0[RYV9\P
4<8E?G?>(H=,@9BeP05b+:6?Q)Y1M6Z=-ZBD_=De<46gg]fa-_P4@.=]LEFAZc^:
+fU_V9>/IV]JA]>NU8/74,Y.fQ<U##K68PEA+W[50cTM=XeC7,gLT::2K),a1e]U
P_-(1@Yc,#eC]eCK4<U?UBdZ6M9JVKb7<M6b9bB87#0Q3Z-OgH)JV4D:XMQO^5:#
;R-I)5;QLY.0@6M\eYNNe9((7@86TUI/4=/d4:,+\=?PU803P_8(N^7[<^Q?C)4J
1GMU-VS)0)PT#N&=CEZ?#+#&8=Rd20CQ]N)H:<I;S=;4#-0.RW<;a9&7QO7#46/4
1JQMYDV[D:VC4.>Z-7EAXWZ#K;74cZCZ+B6&aF4<L=dT,@5eA(G)9Qgg3DM:R(3E
(:[QGLL2#[?B76:a18_EHPAF(:[/X,:P),b;EN_HacC#]PD8cQI25fTSBYOY0]bf
O[6VE&B-\3Z60CE@D-S;>]_gZPH;gLg]PY6a60T]-N]4D7-:3&d<<MZNRGI9LM#,
:7AEA_VCaBggUeB:0EW;.c0&D:a-V(X<AIZ&-gTbR6^&9IYQ1M0,XRSaQOYJ&.?T
K0[Fe7JF]?J))Of<G9Qd&Y2S=J)X7&KfW;XV6];YcCOW_dYQMG?dbG.GLdC<MIJ<
C,NUGXaG.N0O(1/NV^3dFc4LZNAFM(:gMMA@&O-M1VY._0H:1>I\U#5ddbG<:C6S
0E^CR^D^-G(CY9bI#;Z&A,>(0e>+?4&J2=]-7U<E2ZO;C@TQPf6V-.JZfXP;70cI
&EY]I9##B#]/b2S;^T1UT8(4M7U_59^M?<Ed[45@_QNC?fCQ.[DG.\WQ:D[NE#(0
)#IA:HXc--@>C;=G=Pg<7/XSDaU[BbB)Rb1_6O@gWXH>d0XB5,3<f]c<]-[0c6?+
^<?PJg3Of64.)<ZfB>8.))-N5dC]RCH_XDM<G(RN32E/ZGe#0gO7cDUGd/4>VY-\
D\\;2CN]M=b1EKWLXU,1>@07>X4&0NI<bLc)[D1I\M3CV<BDUK4NL^fZULU+DH9:
)IMD>AAKO14T)]1-A[O5Uec_Ub[LV&0a7OdD_H85?b:M4XR]H/T6@#NG#<0LX?Qd
Z+GSDJYLJ52c5D5>V,31HB6W7JU2UK1LdG(XB)1.81M6IT@UK,ZJLTgUWE]:WF<V
5a<d887Rb=YG^&G+H0AWE\?[7Uf(ND4F89RS+NYUBaQTLIDQTRc5:9]>&Za&Pg(P
f@Ad,KC(WZ&?._8(6Q2M_VZc+F<]ZYKXLQ->A?SYVHH/2>Ug2.3f:6X04TZ;J+I<
<98B4NS#c13Gc_#7[:8=AF2C,7<6;/,P;GbR))L/RFad5f.2XQ7@:W+/J7G8=F>B
I0WVGFF21aLKH0aAX(TaGM/KM+dY88>UYGJ-aOQ@c0_Oc,LAUG96RfM9LTBA&2R;
a3J^PG6gH;MS@68dW?&>d7)Y4&Y@8_5=6WAcC]Bc\cX3U.)_+Re+LL_?YfH8,gH]
29]0OON]^)ZV<(=_Sgc99FQ3P>[K,WDc.2T.#-[BM_@32Z?QPTec#,?g68V^4.Vd
,BPI\Z[\JL#@/YH8/1+2c>GF3fZ18;\eR+PNe7cBc:cT7157N@e6Z+[>6^=a+BF.
;eYY7K4dDf&Y2M<6L<O+<.(L..AOLC4EVdA(cN-4_:GA3EK[?Cf^#IgcGIW\,,Rc
A:HK=TD&?7;1CI/;JFR5+[E<0dT-9[CYR6P_3VfZPD##A/(Z59b5?:0EGPgIL)-e
U5^LX])f++[Ad](ZXdRD9&^cWHR^YN6.(/S)QS7\d/B__8CPWA/VC8SE-W_.f(6S
8a_\Z.gT>&Q10J#U55SB3/VVbCDU](^RVZOJ3W&_11TX2EZc#OfOO\W3.a1QV9GB
O1J9IO:>2cbT7YbE1^_,?gdVe3:>_BJS=]DXXT#V:f:ad#0VUc#)O42A1(dNJ/J@
@GZGbg9f]Ua_17IRCbbG:e;MbC(</YVJdedZFf.:(63G/DaC&A2<#;-V?3c0<5cR
JQ&bOD<T]R<c7;J\561]ID9UBU/IdeBTS[<eDW3>=Y,GMCN+J.Kd[_+MC;NQ(#+N
N>G.NWg4Zac5Ee_f/I,]+Mg7O;VdM-L1:M>c8?RN__.#E3V6./AFE2RJ0,Y,LP;a
Ag,?_BY(ZGe;NeO>[5[g6e0eC=)D^VPcF78D_+AcOO/?a@TgE]@JKG24W@V-1]N)
&(QVCdWB1/)9.YaI_SKJ84<Q\Ad>Db.JX-.QDLZRO>)IHUS5E4eX97I4W)-13N43
N)NJK?)>Y2bP_\f+D2G9YGa(2NdN,Y=RF\?>^M=>=/Adgf_O3e3+CKHa;3<&JT,R
:==U/9(J5d9)9SPQZBJ1QWd.)GU)+PI>AbM3_8>?5X?[[<5D?/0>5a;.V3Z(FO_4
\X-8D323RQ)V,]_2]AFNO&ES/)a=##9(\BVD.W[P#4Ga8P2SMCH/M328P=\C3_4I
2e7a-,G/_B567PT[8d7]CMI:S2&P;,TR-&#1L;_R?1^F56>D3@]H.<a5cRgD^PG>
7G?B+,8(9(XF\;,+@4UM&NY]5f<NdI)Z/+BJJ4IJ\ROdQdF]DQQ+fH4DG?[Z0P#A
&Q+G(-/CIUR#SW(8+Z_1-HB+?BVI)G^?MBcgW&H\6OZ_Nb,).5TfL+Yg34XV,=L>
OHDZP6NK?J&OE]E[H(JX0,6JPG<-M[4<b3XMBe-V^#g&#I#[fc2T763fZ[?H:9&P
V,124);gUJdT24Y^>3ca\SWeg1_YAX(AXO+)3H5P)?04]\W:->64@?1TJ#gOB]JQ
@AQHYV&YH>+b7\T(H6;3FcQ/,HgN.;J7.D8#DB81BB:;,7(KN36B,P+77_T;=C,1
)9?g+eV>LEJf0Ye-29T+4N0NEW]+)J=2[@>-55,cJYWT/fc&()TQA_26Tf[f>=>-
HZSM475JP5+V(>K&W].aW^G4S4<a+fGGY;feYN1.Q7QYO6f(,bJ9G\3cZ=^,ASKX
UYd=aV,SR:1f=U8/.W\6U4gc_&&c8-2=>?3abd:c9REWaF1ZN+Q&DN14c::,]/NY
14EOd4SE[IDWK)HQ20GPL;=,<M<aOH96[98#1g]6P@I6U-8f=@cYUKc\/Mf54HeN
;@H#9d+PI?A/d==8UKg\dfgfSH?8f5M7=B1CRGHbJBUQ3gGVNF#9U#@Q?U/N<bJb
U^6D]]<H1UP?3-CJKOBP(X1g-DEEEJSeSL7-<W@b?H\G8T?DT;(ZR^<<NZ-L6J3F
<B4ZCH3(4H1RW)ZS@VAUOJ7F^7ee;T=#_C2Y[QHGg7XECC(ebM@Ug)A,01#E^>O@
@b\OVIX>6Z68W3)KPAAS,4cd5cSY:dXJfORZLX=O0SG2NN?3bQ;?\6edHK#BWdD]
A^46a_WfaMZ_B8<5J4RAW2X5?=<F.KOU1a2S@WL13J9Y_LXfR[QM[W7>5gWNN;CO
4g\;,CKTfXVbGE:7K<aNCd&GPY[M.45>8Q@;L;6P>\4V7V:DJI&>B4aXJ66&5[4O
LQKUT<:.eM;1,2fA36F]OO8fd832\EY_eK;_dT]H[WH=+cW7SbQK]NfVY]FOb,gK
<g:14>6b8R6YU(>K,G/EG@.2bPIV/)(R\J40@.^;U<>g<f/;b,0LWccI3JPJ(][?
_0T\EeTYACZ1>I^F=E/<=C6<5(&(RA?\f:FZ91-RL9=I@J9A]OG_ELGCbc_,,VDL
4f53gYe).T4L8P??0P>\39]LIH>]31egcR?)66U:U<V4_&9-\VD3La&V17\P5;a-
.;G=U.&0MA42V9=Q[II1JC@9L)<UJ-KKK2&^VV6C42,LV8?O:&1eD=0=E@FZU7VJ
Cd9[IBeRV;(SVg#Xfg9J@aCTG#T:.ggaeQ6>I8_B@Y:+1HC(7E?63F9e;^K:79,[
+6JaV;<)>ZRF#0ZJP-_EKNEJ6G5)>9#]@&RXM_Y54eK8OYA3B^gd_;RHb/3XNe4f
/egTF+P1>_,>V<?M>gH5P,+HDfXVKS/:JbM^\D^FZf2.H2]IU5>#_B8@.HgRSP@M
KOK1T9fdc,RDTUZ1c1=a&3@N?Y^=&>#dV+#0K#0A+3I>N2BIFMVf)TXLD4Z,8]Y8
ePe(@CeLbQ_dAI,JLCC/X(_:3(R@abUNb[<EgT\C)&M+U_/;XBWE+X>P[JQHdM)_
G,?50/\VZ,0V;XJ>:BL1_YR&?Z<Ed+7BF5#BfS36Y7L1E:_,(VCA))d/1Q=_Q];P
&+(^d>HC-T>H@W7f.EK-#O6TFcY)65_(5MF&\:NI2&Id&PAX9>N+8?dJ5MH0SH(+
:[)KO5#g0eC<ASW;I]+LHIY4?V3e]H)fKBW3G@6b.;S9.ZFD+D(/4E7\WLOL/YTb
3Z=aH2eEbAX9]>I]b]XZ,PR3:29]IYSX@8V7=D3OHU?7,0BL3<<91>M8Y&UZ3&Uf
.EB+NO[YX]/Jd)^L&GPeVbM9de/34]W-Y;eAd[1T@/:,@BP\TTOCEY+Q,0g/[]S@
b<=/cJJHb4S3RZd=R0;XeR/:YeUWCN;1,g4SQW>dARNY:c&Z5cFeDGTeL2CX^@(g
#,<PM&C<56e7+++JXN-[>7\A,f+:=.&)]YM4K@^?4cHceRG)4EaJZU.G<CV^a6KO
fCZHAI@Ya\G.)5;9Sc]M(_C5-(IHFb+O7A,IZ@7/ROG.S21-BeRL0Mc/,;_RG83P
A>+3c:Y3IRcgO+f01)QJb(,QKVa=bRHHXHTPD#+<W3(9/?4I33[8;(e<Zf8YIL/F
A;KeOMe4SM2,V?UJ)/ANa0CYUV8VdP5+T1-ISBeA=&#T97B4:4]X.Ee(V2JSSQ3C
VF7GB3-3H9L6DL?C06&[I3M\VFV[W:-0CX1.8SWQ_f[1>X_ARTJc>V0O&5>Y;KQI
R1ba5#]\J7[+AVG7@T\I8Z\EDVC6^]g3/\LT@PL2VF)OVM+U6e7DcJMR)D3\2\dW
O6YXc/47b(LN9\,KZgVD#@+PA]W]KC(6_B-J6,)G?_Y+H80L,ITc5&<3VJ9Q#PG7
QL0.be[]g\D<,W]NaJ8ESN_\.A9VSOeVK?@<cNfFMRKBQcW-3OIV39Yf?7R+1T@(
+N^1^@<??B#DOVa+A)(]fFO=Eb()8WL)H3?4[?=[_&L_((/430-V:Lg[[N1F=7H0
Y6(1dY@_4JQMCF(2@4OII>=^TV>-+9@aZZMb.1VCReR,Q-4bFY_KHRGS_T,O&cB4
;e2RNe0D[.5>ZfP[>B^HbU7W)_C&N::=fHE:V[>UXXA&fV^RP<D6Uc/3D9cAb9Z?
;M\4.9D,(<?F9beUe;?5PKHYX#OX<V20HS(Hc]DYU;HT\:IHD(a5CGe81_UBS@QL
CVC\2WS5V+FeK0_-9Y>GZDcB8BVJSNJNI7HE]8c^b)@-M+63&#R6dN5JceC@6/Z0
Hc3<IWcBF=TKCfPLRKE(@5Bd:KdK8<O_76<\JdS;.]NC^Y9a)U;X/?OUNWJ29BcJ
QSCMgMN&E):?_0I?49KPWgEf-RHed@(Q0GLBaD1[#U;04b)O9T:^Ob3:b]b5G9AK
gRDB>9OS_DL=]8L;-=+&;UTWJ&+?F?[5D.05-L4T?b_NPIFb:@Y-SIV&)Y<:/Q_5
e)g)WXC_\M,A4:>4QS&_37S^c^UYRZH-58/Y2PHSU<CeFXfdAS3\_a/2+1GRYFg=
3X?-f.Kb5S_B/<Se:N#C6.aUd#e2(K<+8[0PUgKa&5bFU8ZPAA7;@:?@.H/^,Y?,
#2f,9eSLGe[P=QQ8a_Y/M^1Ace,Nf56DCB+A:DbLEaAGP]F3a0aT+KPL,#66B1:f
#SV)>/8OP<AM2g\C6([+4I(+:aY]LM@\SJ8a;gf4+QHNI&cI8KT9[gWR4U]C4I<f
22^6/JFKFc(Q=2DN7f>e]:4W-=^W];0=@Rf>,Xg>&D2\1CF[-[EbA&1=Y477X1NE
99D0<.K9J\)MCA8C_L657ZgU<@gC&/gabZOHT>G_^^OWZM2M/3P.f1=--2A2]7Q+
;F3g>9P6@R(3bST:=RS,<:3G0f&(7\2+07[Q0T(Gf.P@)PID=GS[Lc7JL/VDPc_=
K&W:F2>GV^?>X:V#VAFSW-LfJPDfJF.a6>4FeLKWS9eb30DBH;/#G&[FQ[cW)H](
-.ZAB,659N[]Q3>S[@\KWN7?Kf]01d6gEQcO4>@.?5cB?TcDB?<4,&:F@&=ILF_Z
[#[JM9e,1b0B0HJ.VVfV,-cNV1W?D;XB-)&I&-@<S+gEM&6Q)9-Ze<T3G2Y<[8G:
SC=1^>_;H;aJ7MJWEH=VUOZ-LEd&Y[>Hc&D<09\ba+I#\)GS7WKgFY[>\=VA[\@6
d\=BD?1(TFL;2JFeUFbI/ZR<IGX7-&4[F]aHe?XDBBB9T(J6B>?GQWH5:8?G#A-S
=g>d83H(f^BI/c:f2\NX5/:]6ALV]5-K_V,Uf>,<[gV>TGFUI0E)a5SQI>36N7L[
H[MbP8CAK+.^#4_;HF1RUI&5\NUdeB@RXO/)@f)P6bf3L:d>U3fFN;-I-5-?YWca
bE)F=G0SKEJI^P)#=V>W+)1TcdV7U<Q4fSIQGD_-^CJ+9YQO22Me\=/][VVeV)9B
2?9@68a_S-?/N4^gD(+8=&A[g<-^K[40=#:3YH&S6_@XV#QIaJ:Oe@g^eQUHTKFX
ZK@#P\5\9_N73IEM\ST2LU5-TWJ3:dQ+9V0G3aFf<,A2X,Z4E9=JVb>Cd=M\gd;-
^d(b,.]a2(5+8651dQG\@7OFe_4g:,eCCO<:7e1ACRc/IX#(@:ee.Z1#,]=de^#S
G9Be6g\cIe4b?/[95XcR&RPUZ9c^5(e4.S)R687eEMGB4#e=PQUZV1U60&H#LB[K
cZd_2E)C2TC9ecL\G#0RX/81fK>3IPFe]W,N#GNMN?4YJ=(&cFM&&&D,N=?,e^=7
#:<5W:3WB]0/FY>:3VE:>+a:BZ?.UaM1g?D86;E+e^BQOPWB@fN:^PZcLXgNcW6^
SC@:5)S1_[DQ1Wd)RLB6;DA^3?<g>VdP+=aBe12P,)>>)_1dAPE:dF_,NO(-EGa)
8^FS?O;6P@0Z:MPE,;QZ_^/d:eVRMYHWRgNRH0M28dcbQ#eB;K3K9<Bd-D\A5O=J
MX7HcK-?C&VB/\4C0?TWS\A&(Fb#[P/_M\BUV>ZU1FU[D8E3Z?E<O_=40FR&Z=4b
L05#5.BS#\XE?CX7Kd+&(<UNHDcT#:_3(C8MMVS5:#]K368X5(2L[5E?FKFE,eJX
[(W+N0Y9_bYRcOS?1:15,MK5,X/[)X3G1LI6/Z9]FfVIdE2fa2U9\36I,#^G5TVB
;Z79\[^^A>)0,FCMXR=KE59/;[3(&;gPe9K-_5b;gDL&RK+-S;-Mc_RTA(f?7<a1
ZSAJE=T+6&Ib0B^LTBM.8a^C7N8U/BU.].eCI?(IAc2G\gH+]F3/;3FMC,+C.Q/&
71Pg=(VH]5a9MB91[2U1J#&)?;#JD;e+Uegg5(:3A0S,5#E:b.Z70>+(db\Y>VW/
F7;FITC_8HgP8-HS-AZGL).1TAS>N4[C8[<ScE.WdTX9PL/&Mb3(bVE(9YQa&.TE
DV.==@E:@=C,E-.d.(E=Q8g[@74WU[WRBL@J\9Q^fPB&:,(7a14RI@]W^HH4LEVX
EfX/O1#9\[FO4MM:b3f^bH)E@D8KDD(.SWQYL<W=e?YHW[QH>4Q/FJ;1)deKW)_/
+b[T8d]Wf=)c>#MZ&Z-@GDNF5P:FGD/YB[Y,WAR?U>:B+9>P.YI2bU\P&>=OM4YH
XPg;Y50eV&\c2>T8;8EM6.<S:CfU2/4OD5e6=,QbYdgaA5F#7O-9e<AJGU<^WKS[
MdZf??UBN-\\I5fM8:7.EgP6fAF,=SRWe--.4]eda7KH5G4OOAB#^7?_63#PL5D,
A0b\4_)UVD>SN3gM4M&X2ZE0._;W#1&>T3D-2\LGYgcfMZg[/dHFQed_??a9U4D3
D[Z;B3CX<+.Y)M[Ab2_^dfg;Tc6a)c85A6c]I3EeeCVB4XQO:g=T\P:Y\HQK[,ZA
+51IO=7L8[Y1TD0]+J?fYOL.N36W](b>;_^3=EI-D)YL-SM/-AJO15T>3T/=],;H
YfcU8gL\Q<,.0\>\+0Fa@@E,Se(@8E:UWN?.GaYc0cb(VgQU)T7K0?VNW+--_:;.
Sc7H4O)I-<ELILRa9.C@FOO=^KCWK]C?E\:AEgL#Lf;KK2bQ=(ff-f^(25=^SKF0
SCS6UX:/<)[9;bK69Ic601I5H@#-dcN3Z#eDHFW8-T@:>D5fAI:0UM85JcDb-9(B
,15;)(D8HCgH2&;>(^3HI=gKC[)bV9ELX;<Ha)b)gJ[TO274\a-YRF<,cA?BNKB5
=0a-@#\g^#>3+9HV9?M]S=._1F=+55e]A.Sbd3X,?4VD]H2L,K@>M7>;ca?#F;<R
[;0COUJQ##:RE0d/_BP-K0/[G&-fOUMd51#E[S-73Ld6VdV8a2]AbQ]:R_FVgf7=
[^&Y:;(&SR]P\]O:8NR@QYUgXB&HYHN[g0f6OO9H,>G3g;0G:Te/:?<4eP9W7/Bd
-.\d.CT-1P3gH;Z]1a^e==1b)_MA&##P:Ca+eK28NZP39T:?Sf]&[)eMB8\.Y[20
6U6VHJ9U:ME]/8&Qbeb&dd[\RaA<=3:)3L>43@>>?&_.2U.8<([Q:FQ^eBHMa,6D
PDc30V-D8+\S/cV@JL>\W<\20_b+aN20(\a)[7;]?\NPLRQ?6@S,FMe6M##HYUf0
EK-093E/X]g@\\Y[O/@R,3H=:F8JPg)L+dSbAH>N/<d<K84-Fc?END4d:eNOXEZb
K?H;[cCYS([.@b1faBe;fO3,WJeDJT5gY<,@1L6]YV^[BG#8O>:O(NPOWf,_X-fe
7YDBAF1D-TTcWBY+&TZ5#ODS67\-HXGS4G:94?CA2DbdD>7,B@e_=D0IGH_U0U4D
3WIE+)+&_?81WZCK;Z7+e=;Zd_(eMPJ7#[/@?0a>D\E3TGc0\I\T1WGI#Uf1P=N#
&Ae8&(f9G;dSZ1aWE/+_CAN4QBb>E.RD;#;_@DZ#7V:.e?YIY)6[I]@;:3W;aN\-
CN]+5X72RAW]8R[XWg&&]PE5,28TS+Qc:5L+.U#D8-[G.D:X]^PN](8eBGU=V0)1
/6I)O:=SQGHN.4/2=87(C_=^S9Q&C_7K9GM5I[6A?OJPd6NeO]^AX9a>N)+5:eSe
3U4@9Y^++N\/[JDNg@<]>bf/Y_CdO6R-b142-G,4&I21\g-GO(I4T+[M<-C>.6_O
/N>MB)].b=A[@OGOV_/ZXbf0&dQL6_(NIMKOc1fD0;7V;ed/+C/5B&.^T#(319D)
Z2\20OJR43BZPSLdMgS-?Bf^&<((LDdS5f?.?6EOVfUO98^fC@YYU5OWJb:Yd23:
.B]Y+dIW&.SY0BHMLCYf#gTK84;eY(Kg[TPTEbIS##-.LY_K@+0X;bd9WKRaB4G\
HDS0NHafdAQ[ccH87A.>R5E0a^SQ@OYL<P7g3HL1TR9#.=MaE3RF2AZ[75MUU>D#
bYWS+d)/[Sb7?D7Ob^c<.JMbWLUaC6(?C4D/Fg+Y4:QJac;fE(7&=g8;=dR+?3+-
IE>@DdYeDSCHNfK8]Q-TE@TI44HScaSX+g+ME#Fb(egDMBbWW/[CIf[8V;H&HR.\
-9V>@N4U::D@V<1bG?IJTO9.>HR:faSA&fVEJb,ZfRg]HVb[=,WPa9L;69dQ?C=Q
XA^d.#7dJVQ#^gL8M:J:0B&8Q;Z1&ETc^^W5-C/:,6+#TbY;?eD)A:SK)@3WB4Y-
b+JbY(ZT_aAcWg/=K9\F9@\,bLaA:6Y<fMLb-_d//[<MA,_:Ud#&2T-^3F2=,d?G
)X27DDOY37^-EZS,0ADPAK&)X_8.5)(a95]PQJD.9Q(Z2g=XVS[N0dYNQ\A51O9=
-0KdQ&afR_8NR]L_5^DSXQ0YEQYF6-/TA:).)#cZ]UC]Q<gY^IR_&UaOWdO:Y.>:
J3\O:CG9UWL)+^I./[VEBVVW#<bbbJ4)b>JDP4?DFd^&S4cb\C\Z>EXYQF,_ZY_S
;a.XQBG#P/Z_].>a9@]Q]e8,G>.fbVfX.QP]#^ZN^PdQKR[:Sf4,#4O+@U,,CP-e
6.ON,W@A4cSG=T9T@Z@>@2(:2f2,8(b;B0V5]AG\U(@#\ER&WQ:N)b7?LA;BII&#
L(JPS<6&/HgGeWfSZ)b7DA;\>L_c80@SKO)9f3X]F3e&R&0B#aOKb,H:+.W35^EZ
JB49IPcf,-T^[2)fN\F&8JgFPB4MFG1LHW#DSNge3D(?QP8M)eeJbO-SZY6?dY04
VF7LbQ.C,0V#,\B,V=WaL8)<_UM>b&X_\&SJUIWSIY]J[][;246;>HG2K3F/5+RY
I+:0^5EJ+Q1VNMY-d4LA^8[B<)K4#9gS#MI2RK?a6;T6?<eaF7S3QOW-c8SQAG2.
N,2_a;/8@+SbODV]cfa@C^@R>3WI&24)?R?I76]:YK>P-E_B?&??Jf95+2>S4N.3
CASVKe(T5[4:bWSIY:[Na_4a__#P+,7=SYa&VGZ^M?O7<J^U[gO6&\HE:c<B6DKN
R/#7]7G(?CK9fd<.W)R3Pcf8Fc>\0,HYe=:S;Q>f9,J8Z)]RG0@\O\ab74[S=9.1
<JDf.?63T1=BNR>JIKDaLW0XE5aZ^JK[8?=P#MY-H@FB1c,/1<)5F<+KDa6(0B^O
0X]U[T-1(>/Y5.N#.T#AaB?[(&Eb:W)@]EVedg:_8(F&T+X_Z)CHDXfRJG<B>TfD
Y:[CY^BaJU4C<Y1DHC_)cMV5-,60+S)JFL4IB(PNY&gVec[;7W7G=^8/7,8/)NZ\
F8<(DV]/.L#gf6gW)b[)>>7K95+a,-3UAI5;7-QW:(G9B4W6R3FR-fPPD14Q9E)/
8a/I,DObV>E;<?#GL[4TT.1,Qc<cJIT8)\Q-<,dLDf.d_4O>7ASfa0^W#IAU?O;Q
=[?PIS7+7NEA,4EW;HM&\MNQd[E4.H3B.Ac3F?;8VWegW46gVgPPbAda;OZ9Z.7;
X?VAEAOb>V^.7DA4X[)/C)QP9ULZR1#N+1:F.)<[FTL#5-DMCS0I]H-D5G]De=.U
P<D8]&HY@4QP?EA7,_D]=TA<]75=9\]d&^54JX=1NO(1)Z3gCU?4)9&_ZU0A>4H,
e1WEZ;bS._G2&]>DNC\:1-PRg^EDe\Wd)8afZabSNWB=7=b=6X[P[QTR>O39(8.f
-YbGTFMBaZ)4Q[E@f&&7?M8ZPK2b=+-J4C<cME/O2L:A<-RT?PB<5WV2,G@/MPB<
9?[K^ZW0dLK5gJ(@J:R/+MJ(KIT\JLGAQT)78,P2D??6Tc=QQ-Tf<0S2b-S?_M(,
7DdeJ@6HB4I,+7=K@((5/;&F]OgUb3RAQ(O\\c)cMSCU>DS#ZZY/47NQO&F?X3T@
:aGYV]4R(D1bg7,(VfHNOLTa).]]/ENIf1JedC2T+@;R-Y_X?#DPXccTA&cCY\C:
ZJ;X#_]BKJ/L1;^=U\8b(9;FR:aRa=)3TDc]?PFB2T@Y0](./8Y01AdYA8eV_#,_
,c@UFOe^;PUg?T\@3#Q+PHB?14a--eU\WAUa?X/<5Z4HO>:(0Bge\5REK^Z_;\7M
C3\+?SKb-]Z33G@^#dS@<F=GQV)VRRFT(S/X58.\0V=-M8XVc1Xgc1:a?0Wf/E3/
Q2(MZ+b01VRQBFaO_DT[AL@,SN\TPMJAe.@K@WH4XM8KJQg#2+6Ib6_J37W.KGbU
JXOKWQ91,:Vg8Y?KE7&<+Mge<S3B(COLX8fd_@8R,bf>#83_2?RNA>)G_2gXE+Q@
a95[&P+<)Y99^TTb76.U4?e\VDc>/[229PP3N^@(_W67>;;5bUeO70_V+DTEOBHB
dCb2/_DaK8[PY,<]8[DID[6baC1<]_YFe,:E7d)A8ZPS0TY>>:OE7<0G[6=H^&+Z
L(UB=<26V5L)KLJ(W:9FXY7&E[^?[)I?;4eR:=(I(ZeDgM:_6,6/aId<dH.YV()2
MaMA+HDKR)+K.4(&D,OXAY6=3HL1-.4CV6,3dCFF>cI-3ZddME2M[C3,II8XBYaS
;56V]aFc<NdcM;H#5NY1:FHG]E#MB9[C7e51&b=B]KK10GgAfgc\+#716F0]#R^)
QT:@c#/IQTR4>/U>:W7Q.Y5FC2QK(0@AUE)E#2&Zf(AdFW:,7/MC2BG:.(?1=/O\
R#6\W@;_5LH&H.:4M\9eVB2Eb5,YRZ3Y;e,bVaZ1g9J=1+@&D#005eg.N57+1BdY
cNcH);>@WWERA9dS9ac@7aO\=IY=<c00X2\2XA)9Tae+23BP&E;+b2HA<fS]b,ZA
3:BF1(MQST&.,BZ_H,(Q[Y0E847;d<dNOccd6((W@E7^=V93USH;@2gK9D]2d<;I
QN\\T/I]-VVZ914.>/c^e(6MINEU(S_41^Z.TLeAQ&9]FJ;b/M\.P3#4K5NL(=+1
LaCXg@O8RU>Q9AB\a&WTb(VB+DTbQ5L45+c?>7#Z5(.WNS-AJHP;0L/.K_g.fKGf
>eP5;DO+YgR0JDGNbe-EDH<dPQGRRY])/aU;;e1D]:d^]S+SAJaK.:0gUI?[8LN.
E&AHdX]PNQPQ/b&@]QFU?J[eU[D33&QVT8,>=#f7;N:U(0[]1NHDW(RIM&FK[K2e
G^Z2[H]:#YPG2XYV8)8&N5#5K<]2VE8>K#V1Q<+(IOI#2P^],D<#Oa<6R16&O#F)
Q]Yc91PN_E7D<aIDeS@4[)-RQB,PP=)RD?_:M@/EP0132KE@Xg(d4+T;L<._K(BT
NDUL_&N7UHL6;T;+J0OQIDPY_2+OOdI0HBbUg.9KcENJeSQC<#;B6[ZNH\K>_Z#3
fD5D8\-O33:ZQ2g67F3VE&GS>F&V<Q^-a3.O0N&42L+\^-RQ:5ZLM;;0->KV<M[)
PIV(7EdQ&abd3b>D,FQ35?c@K<F(GJ^;1.7ZO6S,H\_MA;;;11NY^X7PD^?#;O6M
g34[]2(D@D-+_/e2OW>\bSS@#HM\g+P?S6\N8d(N89J0CPSd;EV^42E]abBNQD/@
?J1VN3G@>KEQA]K/c3dBV>[7XA>@U#;=&/7Z1?5_fA8RKH=K:eG<KQW=VQ#Z/[5X
5PcPDg]42K.TgP6S(NEBJ26WO[J42HQRZ]g.a,\a_d>2/Qg4]86^I.Pba1-45;3<
>\4Y8@6ZagBaQ:L&-FR[W@>E[Nb7?M__26;Pa@J[200aW.eN/ba8(+=g+19M(:\0
0B\@ZXU;a7=,POD6F@AgRR;DK(f@0HP8O:B.2RU\@e,:aZ^TCGBBJF9_VMc2)GA<
-M+f#]eWZb:[QR-YRO3DfBCWZgKB2H[0W^VG)NZ?.#FPQ;64.ITVA@I4dXMQf;D@
U0L;5V/bV1c7,.5b(P9<6)e,GC].eQ;](B/G4;A1_^3c=&-^Gaf)])^CNK==PZTa
-+TZEVS5:.d^?89c(,)#0,GI9PRARUYY_@L6;?dZC7547ab6O:3G#O&A/^5b0JUe
fQAUK3^VJ2N\?SH<Q&@@X31D;S(b;L8-8Va6OEO)1\?LLO5GJ9_UR(b#,IQ&R?K,
.N,H<68FR.aOD@cUMW=4KI(g_AI+,8gY+)]Yb6J^&KS&XJ)=2(I/YSAg)B?5&+?D
b#<>1811U_8b@^G@1/ZcKW;V8<<J@1)?<L-0,I[+B@F7D?4R+[@9;7KY)G,XH]d_
LUgMg4=(]UY,H#/2aN1.8GHCTN0J-cOW5O37O:=GObP9cEB:7gT&(VT9-X0TWC4d
SSG/>M?9eA834ZD/+_eM;d1@R=H.[+Hd>eAW[R^JBV&(_Rd;GY/6W^Cf>bPc1?aU
a:-_(GgDX2)ae+4a4/#)88BP0KM[FN&S:/AW./3/G?YU44c?dHJWHEN;H=g@^#b(
[6&>[b3=>Q)NBE.87>=DEeb]Ob4^E?6DMDb=DBURB^-eSDC)0IJC,M#YE:aSS<,_
MfdJ=OT78^V,Z,gbJP3PUYR&M.4JPeH&VJdX\fJaC9CHRGZI7ZXa\\?SQZ1f<4gL
Q,X?W-aOcR[dTXZ-S[Rb^J,_H(K;1C>eBP4RIDJQ(cNf=224ZZE)<)\AS2>;;]:6
0Oe8CaI+B\=R>Y7(;#8.&b.NEQA(g,;,3gMQ=UNO^?Q;DFJ8M-T8=#UHdPPVG17W
6JMK03cTQ4M;/\#agNH-;+ZTfW6/N8TfF:Xc,_E]D^IAe?\g^U\S1>Q<C,SWX5^f
^8L,D>5SR<@>[)Q,ZR_LQ/>L>Hb9+Re@?RB#-e\.K,-f9)EXe,>?GNVdK:F&TM&O
FOWKAXFeL)SPUV2<[_+I_Z9[aR?-:[Q37:DBTP?F^HdZ1CES/@/c)<De^OQY]0dH
aK,]Q>O,3[f^-K_7+.A]CUL.U&:39\3GGdTM7bWLd#MU-2OQ819g#7;M(3H,>WZB
fJQ6Z.UO9JM,(+JGdgE,fa&)C<1R,]cATa5?/2;WBW3WY1ET3O;TF5E?<cX;B(SH
X2,KP-VMb_DZI4#1F<H51,#?+9VG<gbf2Q:F99DJAQ9O_Pd62X5fMCUTR=@EQYRQ
1=8C-_Nc+Y51LMCdgbS+2MX&Y/QRcWI&BgEA0gV/J[F7LQ9LAeNJ24;GE>FI_E5[
WRH-9J1/Mg-H^YFM2d\8NG<DbNICAG9#_Ma>4DPI0+EQ_)Y,,Y]DeI4_FH>9fT:?
:N_V))92<<QJEaTR\FJIT?D2fE&cH[7MQ0?YPe^:.@45fL(9bOdGg^F(WAXH,0GH
TQ=:01DXCg?76Zb65Fb6:IfXU0eb5I>IN^E2L(O1,\Od]1XH1F)AVPD[c\1/H=T@
Bf1/7UW;[^5^Kg^VETKIFG-EBD24b/cgeBe#2HN.Y5&-UR#<Q_.GW\cZ+I<RQ^S1
G)V(ZaQ@Z3WP=CS5E.bD3(fH/@YQW>&>c2_0\].RP,G&V)ELC;e,E/,FT#_O:,e&
[ZE3I;DM+BWf\_OQB9<5D/bMFWG0c@@80f&3N&.#ABW9(\5&U=N0G^XTb>g+.G2B
/_g6DdVdKCL1AALgA4]d?PM]#S=O4FU.QQ7=K_0D5=f3[/2XSdUMLUSGGaCNcRJ>
e-Z=>2M(77(H+[c]1Ue8?U[Hd2ObKCVB[gB#7.LSg6;V9&?7):\e,08-G2)M-X0T
OMeF35+T05R3,9OZ[7\,VacID(Mg8K2D_E:<34cQ;].1D/;c,g=]X-EgQ;&>3&&;
ZC6X;2Fa-[)2GTU>X3>/XPV5KG4P(EZ,@/?/8_#F;-.6H5DDNQ]1JOB67&C,P8=6
,g5VCQW\FJW_<P>I8)d,@<N?(/J5)]J+8-a7B7RgcNQ@2dS=fM^M+g0?99H^.-Q<
MYEBdYI/4,QHASagDW)7@@Y.-RS&;eB\>bf@:]KXH+VZ3ULGg.&KPG>.g;P[]D2.
Fc)gFW4NLK?+<>>#C07>&R_gff-(.=N:a<8]^G:@<R6]e9dFCGW+cO^_UV@QRGOB
4>dC9;.Ef=AEBHKSd(8d6X_0U-eMa@.,\<-D,EG>M46]&eD23YF_<Eg^d-AJ\CBb
Xgg3P&JJI8TN)3+Ke,K?f=_05$
`endprotected
        

`protected
?IVFbOWZHGCdZGfE\KM,BU-<)cJG4AY/dLdUf^XRVR<K;2#5R^Q,()K<;=._?@[d
&B38LeO,CPaga8ScdCUGH<-G[R^+;LB8;$
`endprotected
        
//vcs_vip_protect
`protected
UP.VL&Za\3V2ceHb.O37G77;^@4>2V+#d(@f2#XX)\GW++0JgERT)(\UdIA#8XP/
=>312SL_9I4SJ-Y[1><(:<c-=33RWdY^Bb;=4ZBY+BcO14^f_Y+<#=2EL<+HEU.5
E@GU2]5Cg2K4AJ&c:.?f3\XZU+D(=;0JL3B1_BK0<P&2^K(6/#41Y#MD4)S/<_U/
UG)+C1KL2XC&dI;RJ\4FI:NeBbe_R#OYT/,(&bJP[-@L@B[1VFa4=-Y1J3-9/LFX
97&A8VS@5GC<P-FF;\=]#cO?),B_5[+Bg,,<1_?BYc?VL/7adRA#BZ?N5[aa;583
(D,+IBRDU7UD)\ZbdF5QLcW=5(eR,Z>>-#FW18KHD(J6WF2LEDG;2<-8)5.c?G,5
NS8T3>H;<6CHCG>.EGM/aU\EY#-O1S]H^](3>2[2E]MaG^eZ+/3WaW-8K_E7HE8&
aK.]Xc&=f[g&D.fJ&9+KY#QLCSg5D177II_O=_^9VWMNZA/?6JK9Gg9?]LTGVecG
:KLcQK#e8^<>S-f]P-&-_LD)Fb6LVH4>0]/8eVL=B;0\7Y^_<]OP7O[]/FL;/4cd
N)/.<@e[4M#gKQe,F0820^c?JO3FCP0Te/^T+LR=4fga<1e[=<3-b=?a93RH82RN
aKa^KRYB:WR5.R[);1K5&,7TW.&R[+O]/-MGP:_Z:G011W+=:>\GbNP_UgbLdIgS
1&bYYc=.:5I<\MW3OgD7=.9#=&E/ZC0:61\Aa+4GK[<,bTF\Vc>,]@Z1V+DJA[NF
^AU?G42V\?ZaNgVCWQCT/OF^\=#[/?6(_U(dZX4fQ0X((Y/b#[=Ng??HRUTEGQ27
HZ&)7@1PPA2PP84AKQF<@@cJ]#IK,:#b#_dVTKd0bQ_1XM_c_F=VN]#89EAcgK?Q
Z5gRR_eU7U(FdCOI2.fO.ZSB&?a(K<XcXMB/=^T:9I=C@(9#=3Se3I2_WM11/:Y]
#7bYE/[WgOI#d\g09BY,,ZEZ[YKK=1,[;E6<8c2Zb3B9)43Vb#+Xc2^W<>a,@6AS
QN@M2LBf^Z)g6g?7TC>XFb5M6;E&U6<A]J+1ZDgT[\,f_e?B6LdV+;&)#IMG/<N?
5FPBT]N^H2_9K3=+(?9O#KH207)6XX-JYaH(Y-4(U)F4S8#@+MWT/IO>.#<(]Q4d
5a_4.gGY5f7D;RRD]0Jc_fOVcY&:_E_<f@^28D3819aeF,1]L4b\eBVc4<]#DU)H
bW9?J]b5BDEVY[3]KJ=BX2,6:]>U3)3Y,X0[.]>NQ:G)?PI0?74V4@&?5UY>OaAg
]+P-LE.P>301>G8[/[H@3I-IOd::D324MAM6;D+[DHPA,#O5]^E/90<9Y;W;c(W6
cGVb4J9-:/XIcBYec<+7c;0<NPQ-We7#ScUa\_dNE?;Db)adJAH,NJUP:JI<,.6H
\bA#JVaE6OXP8.J&@;T&HDR:NQ.5UaQWJGS@K4ML\4^H67NZ9,Dc./:=/eE2#CW]
?A@STQG>dK@/Jb.>fH(JKg^;2dY0NFT&U,3;V)<M2E&E(^)H<#f6<fX(RKb=,6Og
.B(=U#-N^R&cdFcB;@T3/4I;^NIaMR0NOICTTL7R2QTZ4f0a_@#eL&X(81[=>)LQ
T0T@MR>9PZadOW@fKU3BXSUF]F.f61);UV<]C,^Xd)9&b]W4(#Z43UXg/Zd50gV,
,]U04K3VdK8J@B7=[f5]).]@A_61\_[Q@\>54Q(C<LdXTaI;S^V7VF5gdE,V8?I9
TR1CZQg]W3JIS8S5LL@#TKBOIMHI7C^SJfg-QDQ+A@9P^;PKaKeDXAfP?-<cZ?V&
4-[@P,O1X]<FC(;VJ+3IBB4.fE/0e/>WG1.L:[>3Gf@LgFY5FGKd1C;3.^165E\_
,@QUAH7VHS<&Q]dQc#>;&67->T48/E^#W67aZMU&4LJ6,6#GJ+US:cW,DWP+,@NL
Q_V;JQ:3&KM?.L:HRdY6IO@6^W=\.]&ZYY\<f1B8=f&)8N[R0SSEZVf3:N,N..@f
O++SgeA1-[FI_2a1VMJ8/.9C4SOgCST,RD.Q##R5g+L]EQ?;#AT]N+B\M92I7SeF
LRaKSASZ9Vc.c-CUXBc93?_PcJ)95:KKdeC&,gXKUM=CG__CaHN_e_(a^\?B[8QM
?@]Y\<ae/YAQDQ&MPb:?Pa6A4?#EYg:7^X.JOTYP0d0EccJRFaT22XM>AQ]Gcc@?
;:g_)O-cF0K9WG)N\a:(VL+.?HT5QWeDEWc&PHRQR@WKBSOD8QLU796@^L?WYA2;
EGSP[2gL3)<bV>,^SR5&\XB(BR<GC&0#41f+]P^&LgE70bcJ0I57PNd^2fZ>9KQG
]X)>PceWSTFWd0;fV\,+L9825OG+B1UUTb8Kb\:_fgY6HGfHIe],a).0235J;Adf
/05eTdGE@.4D/R,M/J=AJ.1f#,SUW7+<CX(/A_HWH+^9Q,<MNTdObYJTfGPOCfSg
TX1FSUXJ.fdGAG_M_(U;XOZcaV3O,][?-FCKYK5OSZZDD)g#0dMXR@&bE\16aJ^V
>-\]M0/JMc<Oe_I879Fg6R3W(aFGFY[;_Aa/1Q3CT[_18G74(GcaTb;BA]+B[;fQ
=fGBYM]CFc1S?&?a+g69+Yc[3SeU)G9OD1\K7<<FIO^8/Y-#@2KP47&)+@,([e4#
GHKCH)18^;JBbE/_YedW?eLQTW>;>3MVZRULO\HdfE&HMXR[:+A)aE#RFX)CB(3f
dL]HIHaReY_<9B9^<@U5b<NOT.e+:X0)J>MY4HV4eV6\bXB0bG#Ob#1L[\eCc&e]
eg?(R2ISY=QZA>XFCSd)FJZc&?2#H(Y0_X1\SPd/6DL4&>VQF,2=I+f@N/c[XQV1
KBX[]SZR#B>]YE=<[fDa9Sd:>26FTG^PQd9ZPg:VUg<&L:MaaDV]+=T1YCAN3;)M
/@RH#4]9)=EB->bFJ5H,TdXV\E:EX7N)@M]fCR/.NSfRGHGL,M\OaOOB6g#0^2^[
,2Bc,_Z[O>K1MCP[.IKb_/AK,++a_<O.aNHOaF/,Kf7_Wb)5)Ybf(0g(I+O2g]I:
17RVDAAY0/1N(1>W?8Zb0+LT:8\/\=Y.3\5[#]B111)<\UV4H)X=3->YYSf:R@1&
(N2;1[SFJ6XFG,LB@K1H3TUL&4E.<MNK_56=d=<7:dO[LbQ?Y:)/6S+C-NHZ/R,d
5ZF1DD6_b6+]#[b<1423PABZ?=b6VS54G0F7EE]8[1Ib2A]fYbC;1Rg68Ff=^<1R
MU<2.K=&:OXXQ279B<B_RN&Ad;aF&2.aLS@5[)S5aAOcf#gJgB[&=C0GSIH+SV\Y
fRA?;#]PR4);)WV<E3#Y_G.1,8G1)<[PcRPZP,N&PG@_;2-DN-:]f)K[@P.Y(cfd
ZUYSeaBc68O\VDO0?c)4EY3/J+da(]EVN=c=)8/FY1-5baJHDN\b<GOV:A8ICIDC
@+]a;J?@T5C4JH\97Q9J&X1g&#\[D8[)>b>P1>SF(.6DR=YLKAJ3b.b>X?AL&3N.
50]C7T2VCI+WEXgD67=BHVN(13IYM^B\ZQ\T=3@&@L7>bGS_IE,_CaM^+RM5G_dF
AcW=V0(JIV\OY672LRSHU2PbO9eV#4-1,]A.-E=aYcALJFCTRCAW?>eIgaVEXM=(
9:G>JA0edHM(_d]1,):X]:9CAH7OKJ+=48]_C63K,[1cPc7R2]RH4S@0+&)8ZA)B
1B&=SE8(U3AQ,<b7fPPLe?RS2-48f45;8EgQ.>-6?gB&=_aN\U=KafV#e0_K>8Tg
eV2EO)8X9BY/>.bU?Id?0IGccIKRH\ACQHD2PH__V9AMLQT1R\LBRZ\WBQPNabN+
(,6X;CQ7Z:1KB]XHgXN3?A]cCLJXGVIQH1B(6(].IWS^41><?3JT/)T4ZaacW5(g
55.MQ]UI]SAbWbA[9X[eG.W#E:DYI5D)GJ+]06WOe/2dJA:/GSWT5@-86OB+8/TO
H\\]b?Pdc;+V3+b&_JbTSEZITWM>QVZ\F+8:W);aBD=aM/W>UC^fN41b9c7_USNc
ISd#ZegNQG2K()>dXD8#KC[>QV1\c.U(RaT84IY/,;fL7-K<g+b-56Te\-(^ERBK
T8HEB<d01955DUOeR827[fZ39S>2,=af@CQ@=bgSI4OF0B)<-BR6G\@YFM?<-TE\
]A)7KD?N#gf0=B_P5+D.0aO&U4Eb-7:K\<?^2F)K>M]bCN^c0NMQIG26D^[#UDTR
K6;]I9P8\V7,S4L1cP>#6Y/b2^D+#HG0SQ<8LZ[&\P)?Dgd^0WY)96L5d?S-U-b1
N+)=;g#Sb)92DN83TEC]dZ\ASU6LG6TDd]Y4P,]4UJP6e+EE&b/Y#H;Xc(E;T(XG
:M53&KIfJ,8g:2(Td1\WS@W?R:#T+F>C=c3Q,Aa0H@^\(UBI]]a>\9Se^Q#J]508
\/IE3J#0dVJ)gW\&TPT@eEb][W6FQ<;@]<Y5KN1eON/(GRa&g8@5\aeAR+Q(OcV<
]\U4cd(2&eGQ-V224ffI=DU9QRM#YC:+1V28e9?G3-L.8FK4VR<8&\^5DK4:=,;M
US+d-)/8/52F],:7HB?0F:JR)TeHK,\S6&S2DOXZ)gYE;d-,:JG.-)LW1:_TN>:Q
^B:OJ82KD5F^DEW4FHL\SIQ[@C9,,Y]WZ-FQ4L#gc&]X/-Oc\<</<SKa,VRWV@BX
/@g\?1DCEIDEV8a.<(/,B))aA@)\97.VE]++OX^&<<B;,NW>cH^G1&O=H+T[7@W;
:1LDe\R1PB.F)aLf4;A/8ENK?/c(Zd9?+ZKbG]=-1Ag^DULS/E-1]PZ^ffIf:<O5
7MZC\:c9[>0MYFUP5IcDUCPK&O4d1b49)6/bTV[#]QI;N-WbgLSLR-(-H]S-NKPB
/^?d?ObLNUcdB/K8A(7@#J,ZL=X<1D4gbX+Sf#7/c_g-WT+0:A1f@1=#:3_E3Y_Y
BP&LbA#X#BP_?^7^PZ&NYPMa6.cgPGb(:69ge1^fdISd5fWEG(>CM_fQ9:@A8a5I
+HMOg)c7D0<H6Od@7(f(4;gB;7]NK-((A^NB?PV>CGFd.?I:Q;0RI#b7gbH+-YT+
+32IR,&[N7WCXT4a91P]D:dZ60Le8_\?>8]cBY0#9,<6G#f05_FWD#IN/^gO1N:N
afCB2XD.GC-&7c35\FH5]/IZ,XAf.ZD>9+Ia;?5B4^<af[NAU[?]W,FZN(GG9b,J
/Hgb>g\[X/#MM]egX]0BA^79]fZ4<G1?<b),PQ5&>T8]cN8#fO7SBSg._/ZKF5/[
WH?\UYX,KL/cTQT;MI,LAVKf/_JV0cL=LEA_b0CcVK/3&a=.@F1V-Q+@/;VaL[5\
+ab=@]3;LD^:eIOZ//L>K9J-W0-3Pd+c=cfdYTF,24\9Y1=P:8#W42E6A[Z_R#8^
;Z^O?83@@JK+RfZ9bX/\Yd>J[/-79-B/RKMII>/R4,G#WQS=g)gc)5ZZ5Eg3Me;a
AP]TZ&>\)gc>+BbHe)[(+S-MaN7<\=8:JTCC[IV)P3DK/I.SRMK)K@.QPU9-[?HK
ffM5FXP4YW2Ge&XN)2N8)4,X8.=(393_?cYcZ+/RKV8D@SWV3,AIcOQfW]b\B7VY
15]>YbUgO_H4OI9RCeZ]WK>?V:QO/Q0&<VJU\&e>a@EL9ZURK10BLOF_7YDM3:b?
0-R[]_W^(9cL9N#fGB#,S(TXTJb1R2eFO^_:F?:@55IJ1fFK;(TIN,6M,+0b)>b/
97fIVUXIIT&adaUeB.WS4XS>6>PMYY-(aIU))&Rb[I=-4,>U&4-fUEQWX/HMDXeC
_)3=C6cC7^\5ca=@:FQG6#4S4,++c[dRAJ)P92:WFLega.g=\1eg9\2?;AJ[^(Cb
Tg\^C_ZWP0MP.RF5:=8=FI3RCI(;C[M4DV<Q8S7C2,3]5T^\DC[N9RKS1Bb/#Qd?
fd/7G8WQ-00JUS1H))<T>fTPEZ2?4)G\E4+9A4cTBF^Z-1a3Y&U3EOESDSN,5D/D
)#_?0/M9+gH^EX^=7<VT#-@A\\VIb_VV.BYSI&.CEW&W;61_0)U>OW0C@d5dMK+N
6RO#;UF;<N:GW-0\GQWbFRaI:T?L0:cV>\MF441CE8&UKM621C,I&,E13]0R@Y4g
4SF<6b0GGV0DS-9dCg9R+;\H/7PY+EG]-)W24V/<TQDU=XFPdRcACN(;8fcMF/S+
.I;Z,B.Kg(V6:T1#@;?96:L)73b)Xf\TJeO::6;;0X&]bY6K@B4a5I:SeGF&M8d;
Td6WgG58(/8XW,BgPZVLM;4W.FCHBLA/#,[6VY<LR)3NV<WN=QUGPeJ3[.ZE]5YG
+AHRA)E6-37>E5^+b5K.MM65UOP^+1[daYceUVLY_fF=,^U<;D&E_&;MR:.L.+Pb
8>f=dU6=H/#(K5I?K&76^V[L:9RG@2_YQSR4:K@8PX?;X]5@^g\6NQJTVUWM,Q\M
@/74Y-VI/:WJ(VFeWQ@=-N/_VIUP[TIC4LGegYKEe2Xb_M&B?cVYDLKKe388c[-_
YH177Ve\Og[_1GI^T_07[P44ELV2RE+G9.YQ#g9KA+CIKFGSO1=0CO]\JX0<C8H0
Oc.>W=Y>:ZSV[,YM9Qa,911/6U2>3G->=JL[D)W^-[(Zc.LO_72fHOW.C/GU+6M6
+c7=-4dX0\/,.=]7JcF@B199WaXfPgR/.]_3F1JE/eC-OI6@-OM8^bOII=&PddKg
TSBO(H/c6HQ:/L:aDCLP)PE-)^.,L^PL3,G?OSSdI+B[[^Zg/27XH>3Rdd+e_HaR
eMJ&J)7Ae9J0/P>)33([-3[g<d4G6-Q7fE6>dMf&3=)+^5_?4/3\9BS,]-N)gHDG
abcULJZL;H-;TAC<Ab3c9P[./D/g<)F??FRXII4dJN#)LdA?:0+1ZO9[2?TIA#b4
YX/V29ZRLQ,6(@4@ZW;/+\#Z32DeY81_F]I_@L-(A@RNO(7cg&MUUIMLA&E/W^N4
E;=gg\/QAKL\)L#AN;aATW?#R(S4FNSL1[WcQ(9:LQ9;T[X4d>60:;Fc4McMW_Ud
aCZEA/VT1&N,Y+aCWQ4a9[:1RE,a-L@ab1A(c:JU=YB@fJMM70BfeF?X[dEdb>.H
JDD6WE&^C<>XA]UL\1+f_c.dUF3Z<#EIL+Zc(.&A#bC]J8EN6@b2(MNV3O4Tbb^]
<#.5eR<-fHCc:3U<G,L9V3WT3GdWHb4Qf8)XR..XE083>dOL7Me,2:@__=2I/M_.
:1-L@8^IWJOOX(33J^J>A.8-Gb>J)3AfSFV@[9J[2H;>6XdM-dcO+Wf7#L,aaR<b
=O;g9fWSbNTg7g_c[YEg1,<S0FbFe66N-)X:9(@NSN9HIc0#MPU3PWZ@c>9B[12+
f/L,BLPN,(Ff0O/P+?1EY3<f0DUI^Ia1:0(gL9UM+4\H:6&P9,Y(#-27#aXA+B@<
dUdQT4AT]@2LOFNG;<]OH88Z\BFP@T+^E]8;a,;AV.LZVbJ,4JFOGU8556^E+&+M
,AZ]^f>SO,Y/5_15DP)C(fG53LeP=@/RJ(SW<1)UTC<+.3@&<2,b>8GVFaKT[ZUe
+-W3gg6TQVYXc#R#b1_(QJ0cb2YFGO:Ze[5?;<IN;Z?VO-&>X,<d&JZFPbZUb-C<
bH;e&Tb]O1#2^SGYQ^XeRLPHSJFI3;8Y,E[WK7cT>)::B0Za;2FEef--)5D6:+MO
YS)(/U),N;^:_7[WGa7bY?a=cOe9IGWbc945X&\RHa,]<Db80K5]]Z:;4YMY_>7a
./5b6N]\a<(>1[K,,PVcG37XZBB?+\D4_8[::<Ce/CU]Sa;@U)4<Z6R1]5>867RH
@/A2W?9B0-==F-&3F(d-.;33b2+I/Q?>7Q9,KLUePW8IZ<5UMPFU(^9(-I.d/QYV
f,ag&O:?D[>>HT2P,S5F.F-KP-FL6+gZL0BI5N0M><XR4gTJc6X8Q2&XOXF76,#X
R4gBJR1=J)#3DO4#4LR=-2b2H31,JTeL(NJOE/<H/8<=(eLU,,YZU[F4(QR4?#QB
6G&U;QKcd@W\0-@aYD.NO7b.I3OAe[(aWMF?,5U[3b&c#_0aS3-_TYcg(S+0ITB5
:gVJ/-;P3D\M7152T65:Q0GV>,5+C<d]6G>>&@<2JId6BSG=fSJf:1+#N116/0/,
8CbTL@eAK38OdMR@R[fKQEIX9Z##M453^(;/H/SUKV[+IZN)>dIG761HfG7COf[6
<-d4\V]-T+/6JO<6&6/TNC\C)E:29I#8EGa[TYYD[C]bSM&@UW6=a6#OOLVCQ?f1
L:MXKAFD[H_a0PVNe)caK1gd=BfIU/,#Vd.0G6XZdNY&C(HF4I^?8I#fPeAe]>C\
ROJ<eKU,(ISMCG6d4<FKR#C;bMR6Y#=eTZ,G-d.3gR+QVDC-=(N9O+(b^H;&A/A>
8JX?<34GQW&Z)LSdFXA)\L]df]2O[+/.^.>S;g5H^XH>_(BR2fGAWQ.F/2BM[G#L
[JgNL/Sg;+I5N;<>TY.VU:XZU6.7\QTcQ;#f>bUDSG,WGS7-()J:Td.N/Z9E&PB4
)E4_0;TC].CI2ICF[Z>dT77PI;\MOSGPb=0GQ4PY?6PLd@KJ>M4&P#=+:0SK?JM^
L_W\K+@L_?PAW\^E#c55EQ=C20e7KXF8(IDGR/SO+YU^FabcV<ZA,UH^geNYR#)]
\+E@QM6dB>@QSL\01W0ZT?2@FW;.0@,P3c)(NaG2ZJ74H\5W)#JU0ZV7=TJF=9CU
Z@[M#0S6;7KS#9OFWQO8cE5#;4_GS+R2P4FOH#4]@.W1b\\EGKbAFP8I<WS:ALK9
9=?S=+3Pa2#c&4NcW1dIPJ4_9F.g>?_fO7&gNPQ<:bL3;9P;GBa.HUZ^@N#[PA_/
>QA?5?P<T0a._SaMECTf>:62@;JbR1C6LHS3dH>TOJ>9C@bW0[+@55&c/G>?],bc
Hf,+-.#QN9-b[7V+,QPX^QOJH?6[W_(3EaUZ98F[OVe?gXV48^f9&T@aQ-CB-^I)
3[K;Q49Bc;I_CSe[W(8E^b=PYZ<)E4B[1EL;Z#XgVR62YX@7[9^.ZJI+QG60@E(B
ZXHK>d_eN;Ic)WGS#JcV#4M:T_S@.JP;:8GL6705\0&;CdIA;,4#XaKX6K#dIDA3
aS=NR_<_dP&(\/eMVIB&B4K+NRFB?U1gG8Pb1Y+[,0=OQ[&g4(/Rb:.5\MMAA6<?
8E^G(@L\?.XM_J71U&IaA[5BH:Y5&@)XZYL@)A>3K]O@ZD::;<2@8P-[U^?N#/9[
&^E.?P9f(a>][JI/c0D0UEUI[Yb]WN5D8Hd[)_,MVA>X3QSU08I^a1DV<2^dD^[3
F\FA(^X4,XH7HF7eO0A[6;^?L3Ed2bG-/TMA.#Q0Qa&bdb@L+E<SY1Rb+><..@:Q
_eV7:,),/S8#G75:N0JO?\+^<0FeYDcPY_Wc>&&:PQ6_^_+=:V9?_?UI>T60Td-I
XY+41WR?^bM7U4N4FQS_C>S1&+0[R@aJ=CD4/JaBV+a,/a,G]P&XUMgO@U:38.]9
&=-TYeb2b+32,(8fCSSC\,5g[G]8ecX;5gK?3:bC/E-7cP^,GWFSfS+g,-A?8V?+
,6X;;>.<0Ad#(U0f@<+@2-Vc4;b,a_/e6(+;)c#/\A5aN8ZS5#/UdM194H,OUJaM
Y,S:LI]:5e45:=09YFL4ST+3V?PBO38?)&_VH#.JObU92M,T?e3Q3e++R_Ng@c9+
,^U<KZY<,S1gA9J#KeX33EFAUN?1HMe#EN&cOfVO?cKD<-ZTeDJDNYUHNdAW];g)
0aWV6HJT-1^b<P\O,fb^aH5(a(8A+MV_[ODM?RBbN@&VRV/_fO[bHI57N&(]2I0Y
?[P-#UQC:8,_[#VRL(fV7EL9>D8SFS-TLaU=c:E7/MNZC0_-RY.,2MJN2V.,7bCD
aCB.b5FBX3>ce4GT-J\;R5C@=\+&MF#Hc-7F<V6K<D/TS2HTLfQBe@G,d2G2c?.,
?9c&8(WA,B#.QV&IE2PW?[E1:#c5C36KBd=dSAI5O]4H<ef/Y72=e=Y/5a)(<AMT
]BA555;b-YQQ;g[G/[b)c1718c+c?:=HK?U16XGZWY\fBf.ISId+4LZ<-P,Jg/7\
Y/RKA^2/.4<e_/bB.Ra7ec2c9L2Rf6,Ma_VP@F8#V0bC7SLfF?&D^Q^MCeAT,(Dg
[fUOYE^]00JTW9c]3VAZ-BbW\,3;dc;+>W&?Zg?C9Y2[-5+8_#HV5URbE^8-W@=a
7eA+[JE2SgL8VaJ/1g4T[e?6>eIdKLV6a@-7,N_T-N]V9Ie[F6J[,C.95.=F&/W<
IJE+7R9(NS[HQ+WO4M</@]+Tb2B,NZWR/(b)S79P@J>@gZ^1L-YRDX_^>R1PN/5d
b.]28S/EJd@0-I&COL&1f,[GL:Z0KXR:Q90TXY+<C<;WY=7d;)Bcf3SMadId#X)@
]#cX+\BSI@g3K+T?#((I62bFF1OeN\A\7d)eKH9^G]QVX/T\UM]FRR?@^C@U7-d\
dO-MBS1GW+3/-,4HF5gfLO?]F6XKK^b\CWPbbNTI@>?bK<#1D+2BdR)?NUCALVWU
[JSV#]FN3V-OOZ(Y1AV)bHZg&4/6gZ.QSSg(PYF-<fg[5>F51GUd15[QQOYP0E9O
E3\<V1F;:4FN^PLdUZ_(BU(1VAa?:#cEE>3e(N#:ZVF.9D#c1?F_)UYA+d@<aK8K
9^eM,g<19D_Sce9aT@:90#GZ#S?S6(?Z1O1(Z6K:Qab7#D2KeO2;[>7=@f<A9-&=
>Z-PT(G=NC+E#VHN./_BTFZY6DS>Bf4Y.M:9RE#LGS5;JO+ZeU[MFBeC@K5#?@H2
b(V<3R>g2W#CC&N4U=WX/FPLD=]+M9:&[:YN?:B@]FT[&15&[F@;6N@3N[E>_-IL
XJX90<dVaBf]B=/JYA2;]K/Qg8LA>e>V<8^DSV4_F63Y<:8^@@WJB&C,M_X]E,?+
R&-<.7L/)g5HJ5-D;<]E&;(:\W,f)0<U;g9UO;S>>^13]^ffE-^F5/Meg1bA),2Q
JX/&UY.9YEFBH]U]@Feb7#SDdJ2VZa;H)5cJL>Kf0>+BCX])-KX-4W3M^]aZS<@7
FSbE[-A-LWSRVX5C@;a3\RCFRCLA)K@=S)DJ#&QaAE#LN9\Cc6UX)B]&@[WR7F;2
U?fSUfXZ#aO]c?aLHPDe(S@]>UUCO^?51f[3]\#@e)D:[Ca2MXJ^QeW-ED9?[D,)
=7X<)Z70^Se4ag_G/AIG,+d,0D>I<,=7P.V[.6-\0:P.M^dO@\2O67OaJ_>.N?28
(Q94QIV<g#LS5f/-6=>-:FNW(=5SJ9K@5F94&JX[W0c(Q>0)-;L9gdRBFD<&G+Pf
g2d3dK?:8<BO;YOPW.SN(5Uc4-M(7?[#WbPgB>3H:P<[[=HYXHcJWMY?[5TNMPB4
AXF/?Ka?@69(5\W2)9JH=EN#DWf@H1R-/PIIU>>g71XLEF<NJ5M/#?ZAXF<9E)?@
PI2,,P@11,6GFg&:5E2((-MDI,[/M7;\9B/<+M9DT.E,AJ(LEYRA[+K0GdP-JWKN
1deA_8-<XW=0@dK6(R,RW/@8Rc9X6F5^CVaQ8+^=[a;3f8DI/_H(F>)+bTHT:66M
D/HH1Q[H6;,#GOZeb;bN)-H_B;=UG_;5X8(BTNUOK(e;L#SQ:3(Y#M#Kfad;DGB>
V+JP6(?4\W3,.bb[A+BPZ(#Ya(,06)I)<PgB0/]()a3I:dfQ4[#R66+302][DRGU
eDDD2Y#U+]<:&,YPa[d)#V],CfJD&1,2Q.#=NgB5]<aQfO9=Y<J6H&3[eE/IVfM.
LXFIS(4:e=T.KQ&gQU;IA\d_5[]P&M.<Z,@#LFO4V5KP)N9b#71,[EUPG+((^]=X
J^,7L.H=e;4^feB3-dF9A7G_2?//fAFX_>,Q#eZ<-H5+[J^K=.A:5ZEQH>;=?cgJ
D\VKeB[G3MZBeVM8<^bT-D1+YAM<1e+ADMdcM:=:Sc30N3N)/ZO[BV_0[><a\+Z?
(>1eU1)^VTKSX/#BI#bI8.aA>-8/JL7K7;9_A/WPQ]01[K/C33&Pd:QH<A2:3W,e
U\>L1+f>W6)3\?/1,3@PJg/d;GY7##PcOM3f[5PPg[IPDd=?CV?Ka.f)d+F?90cA
I0fYP^E]F=M(A9e_<,g:4<^FB7+++480WOJ099;<9BP26g3;SQ)\OT4Z@D/df3>4
R[bKd,2,4HBC@O1S^cfg>Gec8RL_88)Z^JaZ90Z5)V)-N:TC5dT;8OLQF6LDC4@,
d+Z2_.X8FCTX8\JZc\=]7L<>1CAU9;Z/2g6=f917>J+_@(7U3[/c<._(Ea1]aKPR
&A6,3fA82faS-F0UYZ8_:=GMWbedQ5eIXTDG64bOSQ-8M(?Cb&>V^Ja31.J[KQZS
/X.a5NOD-FI,V1YfTROB1aK?:&DV;_3KJ3LVQVPI7J<ML/7^]-\AW\JY[3eSY7FM
a0Z>P/9M4>VXS(09J,bEFI=J+^>@O+XD;\50D?O.UL21BKf)P>EC&F4UMHg=FLTV
N/ZeHM04@K-<)e[4K#OL#-D\LU>GA5Hg.CE7c.Ng?KW7#D?U0=R?S8;)UKKPf),@
gLd==(.Q]A)d0KHdefBEXJ:.0C:&TH24VEd8dd@I9V,BFA.3<V3<08dL2cV_:^Vd
d1XM_,CUF]?AU5QYOG2:>dc(0)WJCD>/24QHa/9R,9+^de5HUTBTQ+?_E\\Z+8:_
HRC?]/D9;IOB>#;>gN;AB25\G/Nc[(dL90RcX2f^\-fea]DEKCYJA@]f)IB-;?)(
#eY2N6^R9<TPC2bHVLOM]1FA5G:I)N)=,6#SY@VR_ba[Jd#8S7L-g_BHM/9.+M,I
6DNR)N/=&1,6#0Y^V.dMGV4VV:K?&[5[Xgg(+@b9XQ7P#8+6U.GRc=1E6_;W4.EJ
THb\<?P4d[8YR6@RT/a6.\\-6QdN&>WFT<^=#>e^R@\)M#ba0BdC;f9d:CYb,KY,
aSCSVTg@?+T4K0D:M=H9V-d/_E6)F/6e+_,]@GUU8U_-D5E;.Ta=gWe7[f=Ic6=;
^I6Q0EFE36K],WP,LcB4&:.ZTXJF)TFWK,a0gHV+bZ#2_PF<[:VO>1=K[.:-3FC4
#.;CO=3+6YWJPN4>^[:,S8V6EH(>=VF?R?8d4LCcO]4fEDU9TaS#6]08Z(C;Y[<8
_P_aK\B>R3@UNB54=Rc.G40:]SfBP9edH1+67A#6OKb7KdXI@(FZC,fE1A1V2]D)
bT9(OK)ZB[V1LOBRM-@f><ZMXU38]2:_PFCQY;NbGR6HF0T+M4S?6E6V-=]A>^<b
:IUJcC]955CKDL:;6\Tg=,XZWK2C8D&T@4[^64TVOcPPf-6HE(P:,^.T#A>]Q]6Q
6Yc/Vg=^:R,BfY\8,XY?)15K\cS\G+7X-R<.GY[G\UX9fY:@9WJ95PZ^>.g5g5XT
dI<fNPQ?P?ZC;ZLT;A[,I;FQ+F-6^4=e;]U^W.a\;/#>CQ@FPc@F2E?GeWK&3L>&
CV.?ZDDE\cRC<O^FB<RUI()ZG7B8U_=W[E3BJ4I1Y2LJ\GNI2Mg([0B9]T<L6BM<
U&=:FB;5?@:bHA/&+6MbF[O;6I:MLBf:GNb<DT+?)10+Q(QNd@7<62N&TOCIMZS]
^#aEZ5PQZ0==7Q-A</QeQ=dR<Q#,GYZ=@#O;g/gB5M^UYVOW#4F_S;@62^=G[1Xa
g8:_^EQ<FIH?8MI7e(fbReOJSO4YYVY@N;A-L#TCV;)PEGO.bRJXb1DVIZ&BXbQJ
ZZ([<(^LM1\I_ZT-PL\)YdV[a?&E1C?^J@aF(2DgDgEUX;F+b5Ka@;23CT2Z@&a8
9E.g9>_c/bfBB,K?;Hb:].KaQ;=3HI7O,S:X)Eg\B\,#b>#4F=]<dX;F^OU2;=VE
C^C+@JRKU5EP6GX7L6O>V]#aSgRJ[XN_CgIE,F]1eD:d#C#):<e+4CZU/H[;XT6<
@MSW[5F+BW/F[>/3>L5T;&dd?Y#R2BO=eLM:MK8_0aCZ(<UI)(&UBbCWZS0c]X]@
a)A]3B,Bb5)26@FFF(6C\F+8NA(G?^<:FA),OK,AfAX6L(:#/II@]cgWgYcDTB;K
E(7@J;T&>;=F\]@[YTQ/_2I2N@2HI1CA]P7BWDBC7C/.Va_;]LVLgd?+]F04YbM^
[S(S;2EbgMB^,+5bQTRWKBN@RAA^+/7U(OYI1U0B?S0a2K>c8I\UaL[:)fA.]2LO
e5&Cf4G7.-+=/a/3(/R@KALcYK[3=.gc?B0g.EH6E[CW1<3?&a>0.E(?:AgTO^.(
\e.8c+L)VB<f5C(P8WRd.&W.9(9_>BI&6[;5J9AV-dY:\fbK.dG#O\P(O[:-8YgA
H/,Ff)+2P>:XB<J6W9/RgZHY&?FAEWQGG\+Jfe[T;UM(+GO<eCCUSU3G;^Z)#Y#R
42X^ZdI1Y8b:F1FK82(QR^/_R?]GH//?IX<Q=^2]Y6>;WOYeZ[[T9CVGHg0A(@(_
gHf[1dKQg3A=VR]L>K_8)cJO&AdBOa?J]5YL<G978OY1<1cZ4]J,:T@,;g_Z:fTH
Xa35ASQb:L3/4;MBMGYR(LEQc+XV,bLeETdHRZ9-W4DM609cIUL:CUYXCb4T()@M
9=0PL@-,;F=/1&BJe6Bf-D;8QCIFVfSF@7-fLg7/3U;\@MXeb&YNS:/E-IP>GBRB
LMN6BAf/OPU_>58cfg]dNc<?9SEU3:,I_b[OeFMQW,52K:0SV]B\2)(Z@NG&+MY#
#-S\TL=.4;[Q#9C<CXQaRFZKDQ7:W;Z#)PA8@K2-J2;33RRZ^0M@K0D7.dQ,.J:?
g=)e<&(d>5ND67M+PI-f9EY;cY(M/b7P5VLSC9U:#eK^8d\?2]P#eDR//TZ)KZ=9
/?X1UG,UDcNf6Ya7-(]8e3Yb<TOOHO,2_VCNa-;HQ-/X8]?3CLF(JH8)6_D1[UE(
XF)gK^B=a;)D(?OcWOW7Ve?Wd,KAQfTf)>.4GdR/C<L>8)HAOC3YNaQI4?\G2fWS
6IHZ?#AeQN0S@LV9^2VRV3N@E2)b;JDe&C4:A_R[=d+/3dDZ=V]:bF++gH^M)CSR
)5=fVME_.SPJJe-=P80g<_AT\L&BZR?/&Q.b-)O+fe)U92JgB/e\d&LOJNa[CBeG
Z3L?2[^^Z(A;.W2&1&+aE:@=+ON-(5,#DPD:=5f9SIZaE37P+e7HUYf1NXf1N(EY
A(>bE8@SOA/J^[+I.:RKd\,1_-X5fMMb-Q&?WaMJ0#O/7^J/>MRKP2G5aL2,21<e
/+CaY?ReTcB4_LfNU[MDD>&#F\e><KV1c8>B\4fd[FCB:>ZYM]BJ[G@TV(299UPR
,R2dITQAX3];B.BTeLbWR46@JD6EO>2ga1[M:eXcN<<)]Eea1Q(=543^(5=/X_?,
)+P\VbA+0GKM6>W8.+[Y+9<G;>V]T^/[cFbJ[>[D2YSa-@[.DT,F]f[3P:SYHF4Q
.-9(Hd7[46X;K#3#@F,@9L&(cEYHLOE?)[QAN+dSA\@c9b>ENe^EH\gJ@T^ZN1+[
NbZ^),-C?:(+EHT8EgY98(,5:Jf48S7M:6f98+VCNI\QET<H1K0]BdEIf_<2=a95
_\@,a+^(UNZ#&DJYT,<OZ+c[,FV:dg:E31b56-1/eI-aE)dPcb&[>I;,EW#,;HO&
X=FgP>^R,f+6&3Yc+F,R52MFAa.NF<,8N0(,I&FSdGGT>Fg?PcfGZAGe3X6CG1UA
9ANVd=8X<I==:6R@G@\DZEX;X=>b(QP0gPb[(WQ[.K/_4QIJP;9WJ18gNN,Y@LbJ
):D47LJ<Z#9c\-^e,ZK(L>.^ZK^:85.=<?da5dA-D15EX6F9N<U6#e4#QOZgNI@4
D3KR=_g@2JG#-N-N_(a:]7^f2aR6dCT;Z&[6\UJD[fcLg+]MKDcWO7^(#NJ382SV
ObYC.<:XNV16E:c(DEJ,_6I+NeP:fM=g]^KJ1cX=b,ZPLJ)5.(g+2_4UW(^74.>O
8P@0Oe)0-8C-CXN-;<RMe_<;Q.<MVPP&(eUe.JEI4e-I_+^PVU;R1RONbP;,,OG>
E]4YIAb(W(NE/\,YM0c4B\TM/daAFB51)UIO9+:cKD=2;,\2D0Pd[K+YGL9V]Xbd
0MW7I7)bZOd-dJHB&M]),A[7;)^RXc<KRZQAd7A9()Bc742G3>H7O-bJ@Z7a<#^4
d;+&4LS?-E894Y([/4W<MY_&^;/#dF#K)]TMZ+1>N21^X]6QX0c?+C2H1FZXfe@:
bE/\>I9BaG;P=?Ief:EG7@d4)AgX=/b8WE>[X;&&2aLFCab6:/_P[-XeM:23(3ZM
ea;L5,JK.CCDZ#9IO.3)7:&Ma:NHKHCgNUTOO:E\Vg?e7)A^9VDJ7_32(4\TV>f3
S\)92XVb)2JWB>=61M1^E_R1J)]2XTBD\,E_.GNfaC#.@YYH,a_=+B<02gdCERF5
&)M4fc,Od[V1F1G(BKd<N7<?La+eL4Fd^DXH29^NJgK<9WNA^B\.R_fB]H.E>ZHI
O;,T-(Jc\@QY:6=A&S8Y3)2Q4=@HR<B=8T]1@@G4VW>]=XSX037VGB3-_EeQH9XU
#-e41c[\4];_ac,?VO3f._>UTRa?RSgD_-=L-8_GMb3\;<=^1N[\1eL+^8<OJg1E
gS)-d\)H,5TALUeMWR+I.f<C9XV)BHd++c)g#(M&C_bS9KM?OJDKJ;/X,8S>S6;)
@I)#5S##29OP)=L_26ROGJ6;/@Y/6N9H)WYN4BJAG7TPY,J<QG>?F:fY0.U).ga-
3XJJPB_8CJ9O>RB^=[;gDC1Q-Lb@5QG5+d9=fcgQ538J_J;)#cT3/N/eT/:6JSJ(
V_PNUSM0JCd9NCPLaUN50aCTA\\+_NUL\^OFJ)<1S3&3(S3IBE[S4TIbY?bV.S+J
bMb@bUN=X36RJEX&RaaW(JCd[[1&#.JT\L9V69>W8T_.:g7RFf&f=fU;&@63UY6R
ROdT/TU71^f1;0]B#OSL8VZ5HQHFK2@bUMQ&<gB3U#@,?0HPM<4GZHTHSf#NE3T\
8R2-KE[B7C,+7P^)3T&_Uc62RUQJ5cP2Qa#cIfT?L>UZ2.\I?@NQB#ZE1^/3H@#B
B=Qf?AFadR9UdVN,dZR0[HL]:E14(/@-E^?4eO;:KEU4e:E9I]G_>XCPAK:+?&Se
T2:f71U\+HVf#J#_?^,?1_1]W??6R-#JfMDNf<IWZ73gA,+EAD<2B8:<HC.DR,aV
-+4])\e#EB1;:K[YXF]>1[K+-AR[^NA=7F_12eV9EQ7RIUBZb.OJ)XMPRTf3U>VO
]K],M[?PeIDg\OZF+[3H:]7JcN\4^^aH7c(S,=ag]V=cL@FUKbT^H\Xf&=\(C<E\
e2Y@M#YN-=df<+5FT(M?N^\2N9Q<KK?dW/#U<S5eK]KY+#RG:PQ;A[L[8J8W;EL)
A?(P8J:dI9]YJ+\1=J0d+5EaAIQ^a:bM/fc(,db0.[9DVDEFEFe+Za-97V?T(eE]
.a@/.d.c==F@g>&9X]K)OI#5@JN56<+PbD]_Ag1&1,I6]TGO(J)VgMbDd,NdMC/Q
7\-G\Kg\^g9W1AaAE=_T6\DTSCOK@_c:DE;C)D5#K<0P=XK2J(Q]>V8EQ:6Z[8^&
L:d0c_\^&)=X?]H3[RN(daF=]WY7(Z?KE5WcN2@F]_Q/O[HeL>SPg#OG[\ZWW)[C
Ba?P;PcW33<cc_=YD3[cVg)df79e=^fD<ER3A99,8@BH5G=)GZNBR8)#f4#_^UeL
cf^^GdXEGP+T&T:N3H70O0[[SC=Q[2@bXdgYYbL7]FR,d6WM8g^NSI@?J=P^1JS>
AWMgaSQ=#&eaJD#VU#T6?Y7d55URO>V2U&K5Faaf;.6Z?S?,5END8>fN/ILZV1],
2QbFAY9FdS#QgHJ#QS@_3d2^^ANfP+GbURV7aRYR2-D&\@XM3TA\\X3);2&C2@</
1@(>&?L)S1;WIT=LJ9C78_7J<dUKYCV\ULO[-\O11_e)S^&7]-=5ZZT9?Z\e4^JF
+[\C88+41?]M;&7g7c=YCSL\I-S6dVEX3/K/>XeT(T:UGaI&?dAa]a:)6HU&\/Vg
G8;4b,+67?T,L^@(cB-7Q04f0,UN9GW-Z,d]_f<afOe#Ig+AA(7UHK&?D8EFZO:E
1;daC;HUaTRd_?e?Q/L)@IC<b,2(A9VcQ-Leb##7A/Q&+R2LUM.cYIUR-BaR?O(]
3W2&KJE;8Z)TCcYMQA@1DJYVfR/1W7b9Ee46fHd00aF4XD^Tec-Z[V5-Y-FL?@]Q
H+KKYU5^9FI7cJ@ZR#T\6;X95G,I2#1GeTM0X_[@ETLfR)e?f(<)BH.L;]TeF#1<
T;+f=:AI.ZCDO-@)(]^PSKCT]@R2;+#XO==<2bZ1SBBV^-T9g-WQ>0_?dR2SPJ(;
,:MCg<+=2UVSWDBT2Ja-,\Cbb&g:I8/[,8_K]=Lg-OKT[PE_44-f@EWe,86J@T\O
+g&/+=43R:2<8\F-PI3=U6TEgT)_CF4e8=FB0LP,5I)@d07J0Y;K&6=1UCX(0]_?
IXRH?RF.0W<B.dX>F=XQ9?ULA.=3@34EL+G+4O\PJ/A</)[3I/D.8-VZc:=?5]@1
];?WX==f\YJ,9QN[Rf2>8?BS29+cM.N1XU^<9V8;X7B+V.HUg?],=[cBLBP@CY<f
WUS;ZC4)?d\:0LJAN_f,(U1KS+0QK,F=DYZd.1J>]\3UE+FDLR.b\M)2Y_1c#5EG
QF:^TcC+T4a7BDI7afc53\=[X85O7PXT9Z>E^<[C;=I64-e]R5YIWTEDbKWDYFaC
)NV\UfQSTARIeDDJSBGRR#+4a]\^@@(gGfJ>7]bWD:FH=d>I0C.2343@I]I[EL_9
+J^NH6RZ6I,XQGT57=KI:d+[TfZ/O\b&P7+_0+79(Z.MFNX3f>P@&0-:+d;U_TH7
G4g-B(4V<PS51K9WA]0ABB1PMO++]^[bOV]#gOU]HbeE]0(O1ZL78PYQGKNgQN7I
;XI+TF/F+/\405Ydf[eLV1b04ZdGX&2,O)8Ja8b@H<^dRcfD6,GC].N8B-Aa0S[J
#:DaC=I]59/HE7T_[9TY_8,MCIIF+-</+-=(;1]S7_/H(?GU4_ET&3g]bc7bcP7g
fOW#caLeXCaR6]9F,,3G(VXQ#-,ML^JNVe-aW@T8Nc49Y9LY&PXebCTC::E[\#(4
)OcB?fMG1?1VP+_a8/Uc8P^Cd,f^P.Xd)Z4A)6LCM9ZM_Xa3215EGfT+b\-G>ea;
UG.e4IHWX5Y&GI^<VW(<GNW>CMSBAX/J:D?-H#E4#&,6H)A-I2@Q).S1Qec#W)0?
>]?GY[YSR>YZ2@OQ3BH1MN5H]MgH4E4/M@(Z[/&Oa>?PK55ef(AQ1^]HHb=ACN>T
X5@O>]&0;MbG,E#Vf,gXd=g\>KKOM5IP;&ZG)e9JNV#SPQ=QBPLU7H[/#2YF(/#b
-\Q>+\3Nbgg?D)O;+cOLRHd,5(0OUJ8,e)=6B]XSdTS&J3,PbN[bN-&?=U(Ld^GQ
-A)/U6g)_D.=#7]bgaEZ@aU#=V/gJT<OW]((4)GSb0U]D[H(K,R3<3,4(e]g\f:g
DOK,:LU;WF1Y_(c=^J^\A]ZZW<4\(WL/I:+,1eL0WX/.63=U1ED6AJ;7+7#ga,cZ
_cX(Xd&U.3VHL\&>0/;aY>MA@\EP++MV9U0KC+<@LAD\V27BW8ZLM^#H_.3OC,E9
O.LKVJ;R-;@]7>X1:OeAJF<0@7,9E6[J#&ODcH:M1N/#W\Xd5F3&;c?QEJ6.3_NX
I.;31BdC1\PM&6.W8=bDX<c)B+B+RHXT#9OGY]4LG/QH.5]26/9NHDSZNX&KMS7)
6EHJ\A&@Oe.E^43.6c-0@4B;7Xb<E.\1,;BDC;)[0eW<<:^QCTFC4>-IDaV/;D\Z
a,+1L6F,5aaXf_BVW2]IFAVLV7:+Y@,6D8EOGBS)_Pg3\>&(aC11>XIX8K3fA6U#
4S^W[?Ta-Ncc@LY33(C3DVB>IM.6b53cOBZc]fO\aLbPZ\5?O,H+CQ<)^7?KS@CC
\e,ZHGPbLI@.ZO.\\SGO5^X)/458aWF#L.^.D_PV27@8YXaAU?b0@=SO55IU:E]a
<7:XU8X86]AMW-J:-_bg:8I>7Zg]?_I9,cHDW@b#JfO21#8bWZLLRPB.?GA.ZaY,
c4RCe2?0U15R+RXcVeKfN1L6DF1GU95O1X^,YZQV/#<>G=#7^1>V9;TaKR:@fWK7
XT>&?6B0Mf[9T#_DfCC[6V-7]&P\U\9R@QG(BU@:1dKUW-=KH+0XF1>=f@<aH,\B
B>a&8QFMYe9/N,MW11Z&]00/@Q&B/QPO9KeT5eDJS&15<.4#3(b-0S5)4\5,6Y1G
[SCd9eU)>^E2=/^Q2K\TIT#5W+eNe+[?cSW5f.EbFM4.=.&JU>6KY6:SLU_4:#\(
c=D?-bNO_<3N^SJd?RZ9=.,RIO<XN=XF@(df,c;EZTaN?4Kf1>YTG_b76#7<)KCN
]AJW/UUL5U]\)c>JcZdf3/+YC]JRQO01[LZc)J<Q=2bWT?CRF=3<b?&:?A]aHbZY
-_EWV]5Ke-+cI.HGX0+7,6G[7?J+(N+7\g6C3+I/,]/GU-<\8S;Pd+W/fP=?fGfF
Q\9=KQaBZ?MV^ZA.[IE:J86M(.gASeZEQCVgd#dIg+-\[Y+WE^dI7gQN+1H31:_9
YAbfRggca4J]0)(T\OER6eU?S/TVKQ_Z[+3\;\JXWG3XfJ5PHJD<DZF27&a([@.5
:Y8S,-ES@NGaL>e&[(/0<5C?6J6;W,1@VC2[Jb\XM<[EAb50W51T,cHK95JMeF&g
IN3L<1?GIAd+F-3L_H3O=Hc2eCLcXd>(Yg-gK-@YWeYEPO-/X/\EE\A&3d+aWKFY
6fa6Ab<@<V7&Z10.a@UP(eO#>^FPH5KCRQ><VGQ6JcP1cKX]TYT.G,4PSdE,>9P5
@2e)-KC^04f><T810/EONbOHL)2]f^6I3B?O-BC3+HZI_EFX^:DKBa)]8GP(g\15
;(e3cEB[YK\L.gg894LRf<XUKd9-T]VgJK-_.QV<8bO5/c]deb,;_4B7>dRgG6VL
31D<9VFb&1?-ZABg.NC/g3#@ee)U:_S#<4)F<0Tf/Qc@I?T+YYDDbT;0[GG\/cX0
CL.GNfAcNcXf9.901g&>MO2>R=F;PKaa\BDaS708./&.eD-BZAg))1S68I(&#^GJ
:TP]D=>[/d=Y?&+H,.JTc9-QK^/MR(;2:aILCI:0SI1,geDgS0[+,L+6OeM+8X9G
MU=RMAESBQfe15cNQ_/]DP?Aa5AJf6M^;@cDc6H@_0D]6<eXA5/7NY-OPYcb&bJR
<GNC8<?A6Y&8J?(5D-?DE-M>?1Gb9?8=;C-1&[D\b:GAeYdA,)8^&F,<^+Ue8.Kf
H>2BPHM^:aF+(B>c,+81aL2:Pdee9V1]/3Rg4>ND<H;X9-G5,VH(&d7N,^aNG#SC
JR;W9V^W-?,d&Z\FNP:d#<AUK\PBa_[(29/U>Uf0G=/D.?R(9W(9E^RT#I(+Y;BM
g_H;Rg2/+cM,BZ7R6./9cD5^5;39e70a;J2Xd9)&LOHO?N76N[E<T4ENRIVF)3O(
:cCCA/&ZB8)&OAggU1)HQE-?)9PS.;MCIZf>)U[b8IgC/XBXQeX+>/,5d()6A1,S
aJV^KA:P6U=LY2?R&D8VR8Ge\_2GKP2gUNb&fAAL4R@g7c30GK=KK>5#^.2Z5UWc
7#C\;1Mbce0I8I2=B#P>AS^[-X;-_=_IU\cXTUJ(<S]]6Z>)^&?4BUDK\.a1S2CN
91PO02MQ#.FbF#^@B/D.1_08-3EQ<R=@YJ9:G7.Q\VZ=NX&CW;96L^;<008C#:fO
X>44VB9B3c(e1^a\\[HegN@.Vb3c[VY@0(/1DV0C?HHH9f[,I,cMB6&cf?]J6G;V
/#HEf90[S=#g5Rd?]A<QQYF9UG7]4bK<C6-82GR4+62L1Ka9)2OVJgd9E75T-Va3
a:)YH\VEYK923=XEbJ/G9X)(Y(J]21)1@eYQK=UcX)W.(YCQU(U#:4YS;JSUgD>d
S&+RR)O@<&8e]PWF9M:Abae<-F@N/e:A,].?&XL6bBAU7X+)S9O/e\-GcKA9/]4@
Fc]/YO3c+:M8ZO]:3#b;273BT>bCE:FBZOAKT_DY=4GR74(I;:+e-KB?#5R1I<Y7
<Fe>,C103S14_F&L7::CY>WU^\^W^G(7PLX([F(L&eNTX94SHLSd?QR2W#gEBcRc
#Lgg[@T5U^H/NId^2dPK2HE3>+G4:@==8:OZV:+-Kg)1AcXX:O,32P8,IKS1P:bA
5B.&)2CVe?25RS];:Y>06P(QX]5XX\]d\:YBGZW)\P-.(d9f2e]>gF/;5SC:3S0b
91>^^TS(XJ<3XHeZ,/-dL&I:T5<&bK&5P/_e0S7)0FDV6K3TMge#F2[/>(,N&S@M
8.e#9;g/:G6X:0Z..[ON28\C6PIZIURJcE]3a^.M:A82E94<<0C14;RXF&UTV_(O
:IAD1#_Ag4T)XA&B\V.9#gKH8:7?<c=,e]f;P8WY^g.U1.>GZF@0QHQTH<+:KZ)2
W(&bc,BC:ZDWFX<]Cd6D6DY,X8(@?,&4Z]\Y)@PL9P.\P+XPI0CHFCFf/-1=>B\I
GF4#S7WG,VZP6G)@DZ=aF12B??_(0),JMcV?9F6>/:QV=LT1P1+A6(eEP@EC5.:;
KS9@+eL,?[6LRH<1(b&W.b1Q<UWcV&.=cLZ4DPB&4-.eYN__AQ[4O<2,.CZRN>@=
7#23T-;M(Q?A=F)g-D)82G;V6Pd)L@Re7U^L(X)AfLebZ]EZ\TfAL=SX.\HDgWKL
2Dg(7-:_4Ge5UM@&LTUCP2b#>,B:FP(\Ke&f[86@5CD?V&C;(\Q4gSTMS\NRY4O9
+H,R&3J/XJc2#QG5I.]GeM3+T>D1?WA^X2=WJQKG7CeLPc>]IJ-WC[C;7G8g[[V:
T1I2R.@EPQQ?9C-1<9A76>CP6g&(L;R6egZ4c=J20aS;HA8a.\44b9<QI[C40\7;
Ee\:YLIQL[#b[N?:7[@O3eI2.<M@T7LCcNJ)B@b@]MYC2e,;K7R3d_K?7.G,?]Tg
J)=H)2AfN,Og,3UDG61:5UPBLL@26<fb=+LU2I:3YEZ]DceQZD2RJ[0dA8LB3@(+
8.;EeZ56#7a#6d>dSO16[.S4SB?I)/\SC\L^;?2LZf)aND(/_B7/N3Le>#<aK)W-
\Yd8A0e9,5>WX,Z73:@F4>HJ#7)YFfR&_2^+,fD7dOM\YG9OI;Ae]-\^WK;2f5eg
N,?BWBOdLM.GYeFP5KCLG8S1CWa)NXZB\e\K<+g0MR6<35fKO[69-12RGb/&QVNe
e\+FZL4&=YV+AQ>84_,-VgC_PG.2fMTf<-Vf7-R(=1WXMeeNcE;^6d_D9cG6&-U0
JZ#A&AH<(Y?-NV>6F.YB500M<[7POZ26O_Y9JZN&Md6eUG(Z/aAc5-,Ze\e/2c)a
A\&-ZWX#,#P]5Qd10CJ+I@UfD=4?G@T.A/)g,^U5Gc4b=8.DX(86.5c;H7OP:Z6e
?AIUc3JOD.>S..XUWB3T0JJX&de)>>+F?9/\gP2dD542R-0ba9LdcK;],N+ORI8)
Yb4OIXAX5NF<@fWBIC;#Fb5XN^.<=U6\XVI7Q>,A/ZFU/H..g#VIc+bZ2]74HgYT
0W=R=3K6]-gV-=:/3BON3O#.PAEc^]2M_-_&/BZ[.8)&M5g/68eeM>c)TI+a8L.,
I;++MGB_-dJC&SHeW5,4X7S\L9a:UAfeT4]Y#+EAK5,>__L5WXZ/T#afII3_ZXP1
>0C0d?VP/G9;@^BSBQOS/?BT0=-g<;+43Zf=+JFGdf/d,c8gXHO8D[b7a.VV53;1
:=-X<79(366A7.)DZP\99b7;Hbb/^5e8LBSR3bfN;AM61C+YOA&D(S(DS7L48V4)
5S7fFO<c?0^e4f<UCM;_NXW>_Rd?_DQPM>Ef6JM8a1N+eAN-#TgA3;=W&L7N:KPY
>QbM>E^()g+?5UbH8R@BE:cbIa)\,9UKffQTUN?]XG8gNHT+^R0JeP4=_/SFO8YJ
b-D&AQ+@0c#M0G]U.^bEK;A_#N,X+R>-HWOK-/XIL:_D=gbNO:];FT6^^L//XCXS
,CS<0=2,7N++=#YXg0\F+@.4=8[0MOJ<RSIg5P;M.34:EL,+U==DX^MO++Pc3USd
)=FK:ATOJVd1g4D+TYFCHL4RdUegQS5&UH]bUU]\ef,#9DWRM,43B]Q0Ld8CF@]S
d^_F\Sc>>ODN+C=(&>.YX#63Q@)Rd\eDH=R9UYG/d#0I7dg&<@4N5OQ<S7YBD]f+
58R82KJTXSY;2BR;#_7,NYLNWH^R^@VI(eN\517^1C)XW;;([]UcaTL^1]OA7Xc[
QX&PPg#,>6Q5gKIYP1V62+XaHeHc[&U)7US2HY(@=DO5aFIa8WC-0ZQF1e1O1Nd)
[]&D7R+<=e1OW&F#4d5VE7T^H<L_+>d#7K2Q;^07D)BU@Q83H2DKE4@=ab/eU44L
?7W3[N&(G\]VbHdaXc>^+=V_3J&.@?2:V,dTK=S2]<edY]]WEBN58W?S4V6K;W]?
D&aDSUeT,_c<G&[45^\IER3R^cGH^RSAY-.S8O>eCBM;V2E@[HX#e9\)6W/eTS\,
KJ31aA@7SIN#@+F@=cY_Z20NYc4Ff_J@8QO_WE)D:H/Q_.aS?-=^3a3.?5.+OP-0
4^(=LKb0/-f1ATb((.3YOI5H0<<g[AK,W(O:5CV9;D?G_)[GZV85B7;-^V3JW04c
NYe:#/EN_&^.3NZf+TD_.BI<&#XW0\V?-T[#:0BEP/P\32>FAAdB?FNW>g]g#K-\
]0LY@(WeQ88\cGQ;U^F2;L94ZCNe&OR,Y@4F@NaU,GVG#Xe1(F^(X_2bD56#447C
AN@H4.@9X>X^#c,-U?D@g6eCLF5)GHaW8JXE9YTD]?fPIAd#5C=HZK0/OP^Y:X(_
G@[>LQA\9#<eMgL4XB.@&A-XRF[1f,<=GR\GgVMPb6Sf2E?e[9EC7V]J,)ZE;VQE
E=U9;1O+g@,SU6Ubc-Df=ZMVA5YBQZg8ED,\DHaZc7M]_]VM>PaBFZF)80UHW]HR
<O[.[0PK)ENX.^U[S:)_.?.?R]9I./6X>W:7_03MLOgNS>[-fX;>90.\a>U(1:,C
#I7WE>0CWB1]FHJTXF;Qe#a>XTIH[#/.e81NMO:Y\6U^H44HD2_cDDC0bg0:-SR\
LNP=b_DXW_968/,Tb&4I7A<+b.5fYNP8Ic?CV.#6YZ:--IPQX8/YSE<+\T>)&.bD
/aEaIH.]2+cG?G>79]+IKL[Q(TeWE=Y<=eYA2,A<5<,MG5779;Z(g-&CY#.#7T[M
8\B?-9(7C/[_Ha1LM&].UD0Y:cD_;JR@TINbNMD=7Q78B&\g9?D)Cg>&Z_G&M5YD
7^]J1QOe#Ld:O;.3.]RAY^;^V9_e>Mbb/8d<7\(Q+e3G:5:^a^2/-Ig@gGA-DQdF
ZcRe:3>#ZWE7Gf_[87NaVaJ;=8_+BM#]1.g0H<;1a>.G](C3?FH2bQ]E((;P(fc\
_T0Z3KG#7GTZUKT.W<7bJaZZJ8/BLV3/5H6HYC9g5=OVQ8SQJN3D2N:&Q>Ve_J=I
5&AQ\A@E,Te4;E]/P8GP2XL__8>.OS;,(IQ7QVX,KM1#?I8YA_1dK<5&NBUe:X^L
d&S/07?cZMS_#gBF_d=Z^b#+OP6E8EObU[=:[eU[DB5QM/@G5/[/cD7^/0f9=ZP\
E7^\3&/+a\fbe^6NL3@WY^.]C;^EM[MB8X<e6(S\[5PK^H2-JWRd5b.UURU<bY_Y
],245B6Z0-)YfO..bL@619e77(F7CW-<B3M5>EH4Ka.<)TRWRDN+53-,JI03BR28
)<E>&aBJdI5.RY9KB#Lg6U,3(SZ_2)I>NDgL/+J0;C+SO<1Se7[A+@:=Z;8\<^.(
[1fR,?@3)1O[AA/NZ<>^QWCI=(5Q2@9.0.HZ39VgH54/)f;/XM;G7JdP]SPRe_[-
XSC;,d-B4]1?@\&S_1g/8(ZQXV,S#+c,>b#^7U97fQ]Z[?-(1)I@NJ2\+V9?&+DN
9]C]&OJT(e\Db:J/fR3CBR>?;H_\T76XW^Z]Qa,D()N4R-Mc2\\b509Q#>;afaPG
#89A-[;<]@@C[NBRLH?V0Ef2T3V#)S+Z;P(F39-9a>_.9NUF=P+04&8PH27#DZ:V
D-G-?d7Y0Rg8P6U]cPH8J;gD;14)79E[F9@g=b>J^-R^PG[GJ,#;6&ce&b,^]U4U
7S?C,)HbaDGef08<XIO>E:GOB([#N6VLB.&<6-4c([c5A(>,^Q.g<F-#-UTI;0H6
3Y5;7?#D)9[MP/._62?>;/P0?e(D?(K0;I.8./I]?>eMG)&A-X-D#]G,U-.e9D>^
XYOB:L4]#WSE@+,O_>dSI-7&8ADVPI(@JQ^YcM7LD8ga@+:B10?Ta+7cOU4a8).W
J\#:3E>SC9,\MGe2@3HNbZ3SVCFY=A/[cD?Z[4T&&_ccCKMP,V]A2G>>2D&Q=J(]
IG4R#29T3ZMY6IGNOgfD2cQYBW:RaMU@U5LZIBDK/NVdGE3E<aAcW+X[9Db8SUE&
5=P]6CFDYN[F0IfVbZ;[^(O#K@I9;E646,?)QU:5gf6-A3U+P?A<gP45P(2&^,Me
Lbg=#aLXg?d<&I07&A-bRP@:[Ob?FES2HC0cTg-^7HZZ>N9B&DCeG^5YJ8M:6-cC
=Yg87aPFOV1&U+NYcaRfP5)_0AYcV]f=\KeBXW2:L7:E]Qg<2/#c>W>>_d\S+1@>
M5(^/(\MABBQd5+:/Q#@.8@5T9#^V&.S:T9dbDBR[MF_d(O>Eg1JY?B,68&fXc2a
TP+4FU,,SD^J].L,GT/3O?.3WD8)4>(Z+gb++aCR9BDU+[33,4b1-aB.;?C#@G:5
TgELcNSHXS&[/7FF,3VA\L)<1OXZ(W+L1FG=?=0=Z]J;Z?L>3?=J5[_Ag[HQFWFN
3#0Y]@dfa[D(F2,(0TEd&Of3<7EdbC4VI/O6<g:Vg9B3:PJ)6L78+;IAV]-0dNFO
Kc4^L+P+)UDT0&@fg/]?S46&dV]1MPG1G3P#X<C.fZ<bQ6304f^]?KPSgHS3&:gU
#2VMcU7+O2/7CLd[-#fGggGX8J@H7f3?ARfd//D<Ta7HK@[adf;N54.<Y^bT5f96
Hd#@_R,a2CG,a#NeV++1Fb97c>XM7Wf@X1>W#e@^6c27-_U1+XCM\&2C^e4PMMI/
IHJbT=\Q4#/)g]O^A)8J;MR?S+9_<X()/PR7IXGKJZfTaCS0?>G7YTDTRK@RW)]O
D-QaO.BIJc)N?KW;-)e1:8f)85QFS_D_OV/SUcM(1)ecOP[P<3R2JHfT---YK#Y_
YUY;>DbfQ:.R6NSSG<ZRWYSJ;cIL9XG\-Ycf9PbU5<f1?9YBgNBH+0F@f),#()4f
80[@ISMeTO@+?BWfc_N/9gJ@WN4U7C4W&3XQ.3H(KTga\C=I=)&S4NL\N&F@6G<@
4_Nb7^8Gf3]JY280L@IZ1CQ-GTOSXFbee)bY^0<6;/A^PUA_1@@5OWQ6M=[B:ZWO
>.NP_&#Z3f=/<4,=T1Y309A?_A=Ic2X^49U5C\Eg4?=,2)Q_QA<HgYR\.5HLQDEW
&JN[g_Pb#REC0MDL]E8)ZfR]&eS^>Ib+ZPY5R)XUI39@DCG/6AbU_a5900Q3/9.N
XG2I0:AL2(.513bNDYF+,<Y4I)UG#JE.<H-M0c20Q#E86D#T=F/]L2g2=9cTA:R6
V:EVBR]d4a<:I,[U51b^JMXP+g3:\35aKHB;I;:3,?fRM&3V#.W:NYG56D[VMJ7.
+_3f-DVIf1/@=69YgA]c.__6T6)/+^b4_JKF8.,8ca^=BLF6RI>53@3@8#]^?M6c
:7IG7N=VUMa=K3ZH=dFK9TX4TdB5bOZ).c,9.cZS<8_Ka39AD(\Z7=KV8(U^RNHL
I_]e2-G#F8[[T@?E&9224IU4c@&J=&0WI9g&NLcSZ&R^?:QP,a-,_9+cE:Y3D1(Y
Qf7XC9>Ncg8K=SU4&]a@4BBC/N=a6S)/O]]O>?V+6)TF5f[#ccU32Q/2+>TVR,_e
6A@YF6ZNJ(VHGD-S+gY640R\[g/04K&V1-Yc45bZ.V9+OSg,>6/[;XM6e.N+3aUe
P6TVc5&IRHTc02,2M@?LYUS4:?g^-LG1>.g#XZO2[G+O93#0Y+E[Z;^,J?4]_^Z<
.aa9VFOI3K[SCNO=DMOPG_A?9eVaZ[6]UNSag]5>.\4Rf]+_NRE&W2Y50JW-F[=<
+52#NG0?4TXTZPX-,Q@(]7>()9eL=#9P7#cf1_LO9Yf]Z\>>b8X0OH@Q5I8;(BT?
c_gB.=]S[#V?O+10#@=Q<UF,ZELg\O&IHIGc\)Q152&eL.8P>+-=C@:2DQ/:D5Z[
.N8QfcQMT)HB=/OT@W;K0AeC-#T;1IcGXdQM3495&Bbd^Ldg(LZU1Z#Pf_fXPe22
48<<9e@gC6#[&-50SOH,D9BS0=Id:(OQ(YTH\)?Z=VfOaP477:#Z-[=>1c&OR(B6
,/2a3XVT>VSbbXA;O(/,\E[H_=298JJ[3-1LFT-R_UdIKDREOF-.L/OC>3WX01-S
M:SXVXZW,N^7?JG-(A,aGWf++MGBVE(6_8aR.I(M@GN7Z]BI&e2GV=.GO3(5#c@O
U/YD?QT;Le,[Q-PFNYQY9Oc,E0)4AIS#:@M,4YNMEC)+SLKQ]P0>Nc;9>5bL+^fc
L)^=QCJ#RGCHJXLSRCf+@>2Ae3;<e,1=;D2?X8?49VB=XgH-BSR_9D_-.XF5)\9_
<ES3I&HHV\GP7PNI4c7Pe\EF;B:=NJ9WOH651XNdbB1UA5DAXc+5R9Q,e[f0YK&a
Y2NG^?(:5]_Gb[:BOcb#K9&9O8)fP^H\(EcQ;HK1cXRb>A+TYHObRMX8RQ^bH,d4
+3?#VQ:2#^\WP3bREH/Y#]dY.CTR?0A.+(@9]CcPMWaOfB])/AQ=8VJX6_,RZRBX
S#VeMXf?K,:5JTV>(6,S.e0XOUb6@:8<:;B1)[<&B#RZc:0Uecf[2WWE_9,O9?@;
Z+V@fcg-K[K#6;J\;bG-?.Rbf[4)DaG4L1J6K9c+;9-5+&F;Z8B;^&GV#XJF#6^?
Q.N/2Q_d=U?(V,N^MEReJ?/\]:gNSfWVYcfcZQdVZb#U&U-BIg/=],^LYX#C@GL6
#Z>Y7VMd_^PXB-#748C-4GLc<g;@#K@.B<HMf<TQIM]edbPU=/\WK752X;,[6Y;f
5/3)>(;_VJ#13<W[Y,>Od)d@F(?c2]eB1GV[C;8BXa-H5,GYXJ/M.&@];1.&5S,@
49Z.AY1e#CJg8NOZ5PU#;OBRY3]FNN3/)2]@.YC<ODS3,/G\,fGGd.T(NCI>I0I8
QXF_^Q3\g0&J47..J;WT0UaZ1O.@O_ffR5&c<c=(F]cC.;A\(dTC=;R/HcgX(]Y@
L#:N2F)VeOP/O-LKC;)SPL2[6K.EZFUO,,1b+e/U3gdVaJG-\^,91eU492A;:-,-
F9F7LRA;XcBD&@KWCMdW>W@RY<9UQ:3N7cOe/b.YJZaO)U6g[84A]=^A=+F-6&:X
Cc<MNQR+TT#8.;3D-_W,V&2D5=BH;b^/D^PM]/M0D>KX?8>(:Laaa6Pdc5daQHXd
-\K<^3TZI=,_9_MgeF8L-Y_HP^..VQ3;Bcgd&4?&829#Db[N8],(/MFQ-SA3.3c@
I(9AVX]JIB8FQH8G4f8W/7QIQ.^9f#fWAPcM-a94OXb94?R0O&CCX750Y7:f;J]R
c[A.4g5H4CZIC3SLg&7SDBUH[R]<J#^)I^R3e\,&,QFD9.b8R7SLJ_A6ZgJg88^]
98bPL=4)612^X+.&b7FQ3d0dZ6LKd^C<CS\LJUM@XMQ16+bCa:AL<)OO7&eeVRMa
W\@]W7WfeR;2(ZGKI@N9?P7e)&Ef0BO;>7_TdJJ^H-6V8fX4-Q/Cb)K.gJOGU)D;
4L:/2Q\F=@7^<F^/MHXEU+1J)M/[QY=0H?dYJSB3JFSX;H_?IR<-:ZJ4e;SQ37cX
<Q)5Zf<>Db#e5TQg4;C#.C]Z9EU;A+-+D6T:U]badb^ZRD2G>^Z,3)/-eL0bFC/4
5=:?d5(-V+FBGfSPMNI7/.T.UL[)3@=NPE.49LRP8)-g536CS?9TQ:gQLU#WB.>\
E;dfa8NRJMF:&dd:M?XO5TC/)9&;g1/a.@D&Mb3gYCS\(TV5WS<VRKXD0F)VBC,g
YW373+A8;J4=_VLdN&U7[H4,0e#PIL<bA:_0aW?]/_ZfQ?+<#Lc?AegYa]7<H:28
V0U&Tae#d]VfMOQBDb\P-C]8=4?P<A,+BI[HScKgU3#.YUBLO?O6P.12MCSAG-d,
B;B_61&+6Ba-?W?4-TaI5:&X6W0G=/e09e+T?R@T8-J><,Z2:6AL9>I5EW,3RN43
7AAJRY@2LW0],e/7J32faA6HVU&1@591<cPA?1+V6+U(LXL]EW115+#FH4b;;)M>
I4]9a7O=I\G:NB@>W;d(,2d)W.EdWHL?O;QY])(:K=-+:gCe./63D9;+:UC<2(c8
dRGA?R;C1?>)Wg)^-9/#BVIL=1\9EKg87.8WfcdO\GB;/U>\8&MFe]_ZKRe^MRH[
UE3?[0<CYQF,b+9b5X]6e>J@X9<;#e&^,WR?Rgg+4Gd9g)dOU87:e0=/Ie@=V]/(
A\B8fJJA8+,87^<12g.5A1R[]61\D@:)Ede)5eBWQ(A\LZC3R27=M\;8e]gOQUPV
2=M@B?6g@.bM,)ba)8?EFV9/+;S4]1(G&3G^&-<9aC-J@X=b@>TK@#>5I,R+=>,7
c:IbZDeda/Jab\C/]8TGC:--Sf>LN(_7HF-IJR^5P=3-]cYO974H&YAP?DFQ@O2>
O::D4WT,4a9//JH9=LVfdLa=2&>BF88+e9,87Je\2.YRBd^8bV4^<R9ZHK[+VI)8
&G/V8,?)2b?METa\-&bUJ\VZ9M,:[bN;[5+E3H4/ML6TA;(-68Y9e-Va+@A)-YJ2
d,TK7a]?eU-A@069D-0@RZ#UI\QM5O?=&+OC7]XXDY:Ifg[;7[7GZ28DI?5OLM+B
a&H,]e0CLeYa5Q@g9S=b@JFM9Y/6SH&DB+KO:IIO.4/0XO7QVLSS@O0W92^RX[=D
V/ERUJ6D,[T0J@IN.X<=F])SeZ;N6XgAEI-10::3Q4I9ESG+IHT9Idc^,,N93T&H
g.E-HSW<L;<Bd2#LF=_Q>TAY3S<_:X5E[UdRdERQ^\PPbE+@H)[<Y-eR=eb(J1=W
F78;XZ?MSf<)3U1Z:+]ZH]SU-#Y:T5<./HG](fY-V52B98&\?1O,SI>Odb6)@JV+
G1M^U#\Me<+CFTJ/#1&-F+=(),L+AL+E0A^,FYd(7M6_LF^Z:bX.bG(7IabF92A9
Y)d(OEc;1+8Z](BR>>2fBI2.3a^d^>KRNXSH[Bf5</5V0Za(N,<7eP_EGcIQ7O<A
/+BQS:8Y[HWPb[9ecG.(1WZ;R#T(YFW+^Q<#dEAM:=O(KPcJ[T&TZ18NGPGN(b@X
dSRQZ?a@O:CO:W7T[V,V-&[@cSL,NA?,a<NWTBUA9N]07R&5CU^^D:#E_CJT.W]<
:19KWfHCE#6N_1)^9Q@GfZN&YZP#,X.8;W71-Y)3gMXGcN=B:gYAMN#0TLd=+;T@
?>>:_7_,F8=DVFBW19GK#88]SH)IMGSc^=b>Of@@D^0I6]0>O:TY#YeJ[?bO38#=
#9]a?NY8(H1a_Y]&aE0><BE9S(9,)JPU:R4Z+QE0Ic5c&K9M>V<\/EG9E(JQQT#/
5&Va\:^a5,GCSf@&WNWKfR@g-F1?<CY].>B=932/)T.-&L)H\dV(Y16XB6:B,dE9
[c@:FB)5JTM1b@@NS0R&_A-8KC[W-fE9=1;W+5@P9I:O:R8H(0c^ffQ(Z77/HI?G
;\^])H.CKf]Tf=gF_6XKXMF#2YNJ+DIR6\(=26CT7B3]#7d5OR>5cX[U-2J5Q1K7
+G^,BF19d^ZRUB0&@??7T+=;?AgM<&(/^&0G.@4S:B9V9M<g@5[VZaM@(TP8=#BN
+Ta3.SB/LTL\fa=RKFHISc-L5>[g(3EVVceOKLMPO3,.>Z>)H[#W)J^#XM;[J/gF
0PCgZ&^A,[TBL4[-(-4-<GW?6T&_FcG#??ID&_.^/Y_1D&8PEJP,=,BbIC&O[>EZ
><=7M&MC>#0#8WN=e3Rb1X8=A:\HT8VRXU7I01]7d[,X^:KBE?U&@PK)bffc?LJ9
4+S0XDA,J8c5F6&4E^aB7&..-5M(e(\79@CQ8c8a_7[ZD+@gLeK4fU?64R0NP#BH
cIQ;(IJ,LH6<[8+HH<VKG_0^C5KBIBRFQVbE?0V,YgaP_MDC+=Sa,b]bE,F_A@#F
Y?ALd-6S(2OV5K>:0(1T9=T]c3@HA@_U6UN8)IH4RY&/TT2f;?6_XRPXdM?G?FHf
NUKS8_aW8;9.3_>g8V.C.WN2B>Z=K:X_VdEXD8A\7MZ8c+[M.SIR_2gUA@D^HeSV
WI=L>-X1dbBDedaYD9]8,E;-;/;Y_[9<Y72ZT&:_\I+eJSZ?T,[/+ZF3Jd)X-KKb
<.Q#@IXR<FR5U^H155UHgIA3=1d&f@45T@5;J^LL+)QG^261G-AeIHVHFON.XNS.
X#Td.aF03a^<^61QL[UI\7@NS=a7Z7Z>I7U(MKEJV\3GM+AAGUP5VFPFB.=#@A+F
bN\0S,6dGN.\IQ8,RGa&YQBVSC)9GLDa8gO\/dGe&c#;CG6#Q/X#EbbR9f<PO.:+
W)Kg<BHg]QN0+Pcf.cP>Sb4@&(YU\KC&Z@,GcSW=2(g<-.[,c&6G7-E13[=.Vb#?
S(HK1_PT]M3L20]?Y,g]S7-4&1ZVPK=N.G)NaNQLCL_@]2e2Q.>#B+EaeN#]@]cO
GL/I?Z7a>30,F(e7?\+1gDKQ-9P6V5T4L&XSca\g@/OS6?10>+Y#2T]Mb^95E&bg
?3S#7efeNcVLNN,G[a/9_6WcbWY[.;R@g;>c1A30g4c86bVN<KOVCA5VDR3C,&_L
&&04:>>[d,eSC[1c0WIW+B+1bU/c5c(cN&X[c:E4APA4<@\P(.9=K&<VWS2+9BPF
EdGKFNYLXZ57T\9bLZCWg#XHKQb:W)(9N<KS=?dDCS[V<9]Z#=>^QD.OO_];,#,-
Gac5G)Ub,0\M6CP3YaZ9N/gS-[d1?FPXWa#GbIO&^R.8Y56/LU2VQ0(X/C&EAcLG
aX:,BZ6eVB;]2H\>SW44Z@?,D_P)fTRK_JX@KNW?&7a=(>W7a=eb@Z1cO]a-2cC/
VHLY\[12N):=QB(#a;&GDY[0-1.&SA_^c,1I;?7,&LUJf0OA6BHd>O+=f#JL/D(<
I-II^aVa20bJ#K^)Q.GgfD?JJ6@K_GW\W@#WO@+3#0?Gf:<QL0L@#=&T7(#UYIg3
ZBP+G0H,HABKU\8+&RMJM6NHC@48[0ZL/aBPIFDM0+98d1EeQ=>,J142;+V7D&bg
&J[>;:QJ?<FMGcD_+8JW,WISOTJcfe&ZIF.;f61_S5)Ec:c:1<NcNDM:O?1V.1S,
^EeBAc8aCe=)<C>,9Qb-I.\]QGIY4b(@c4T]ddVXTc2RB1.S=E3[D0#I9<=]W4Af
LH#.M<[cY6&YY#/UYHK3O.EACGZ@YWe)c.BGK@M5W-8=/eXE1NBa3Ag,)0e<MAM.
Jd.2#=YIP.bKN<PO72E9B]-fPEZ2YUXY?=0>[R2b2dY;PA,eDc?-eOgQ=8;[O^[>
I^V)/>9E+3c(X.4L/aAJE<@7PgKC6_5\b6I2Ff)N:>?I16?Y\O>9VK54F:cASCPG
+Ld8>8:IbK8G>QEU0V29<^Z3DZ_K4ZW.E:0C/d]5S_3;QSRIEIDT-V&)9)W9&N@d
b(XHEdT0[OgS]L+Ie=NRaO\?Bec2:#5S]U>U+8e-,f::V.X,=6dYbEPN=^-3dEc+
CKPgb?f[/?g9Q28MS5V9UXTTS@M&eJReFK^eaPKfZLHKSZXO9ebbOJdd=c>?+Qf-
Q/7?<EWSB@IK598Z7?gbSC&TULFBH@d3?Rc57&]7Q<\H[0[9C0\Od8A?QI)M7NBJ
RM=8g[gca2;##9^gc6PgPDa44FdQIY516g4Y+,.DefFU4N@MJ2/5U=DESB/(GLXQ
D\QHg)U:-,e--(5e7dWSU(/1#P0[4-@P(?cP&]=RLM93eZL(BO9KM1^]?BV6&Q4#
0N4e6/aN-fXL/Z\0MMa>=2dNgYH)LMUX1P83+L<QCO,@2QV=EEOeZR(3Va_g-=45
MZHQF3RbZceE4Pf..e)6PaUGL89ae@#^YJC\U&=,6W8&4[U/AGdb2+P+R-g4-);\
[HMGW]44YY)VH[b>W=O6XcIf7TT?)><&a/KMZ>?B>Ye3?d=&e\0[8E3g\>MZ)a?Y
M]W;c&5KA+8>(Jc)Ka<<aCeQ1)D#bK#0?W&K?)^S+@FN#fINL_X,]f2f^L+&TC\e
f#&MU=6B<+8fb0@HL+)LM(7I8):Uf_816[LGY(VAU2&2J+Y/.cIT7,=XWKeCagD0
>FPFL/B0f\#;bD=[B_gG&M,E.M&F;b)[bY#O,HACGc3]V0_=MV9X)K_@6f3TT;\;
][)6S<2PA-H?\J2JM<XY68+N^]Y-.NI>ffT[/Q5FG5R.:B]M8^?^,>P.Z06))\]b
=#)f:dP0d6\0,Ue04LE7)FH][0+=T<EEYT&:;)/=cf0?UJAT&-f3Q_]T7^ZI,3&O
_Hb5]Bf+FT8/DSAd/V^OA6+Z)O\1cdK(R1WAYXAc):XIO.9<Z8HIB/F0/NYW6d]c
Y#U0/\g_@7S]P;Hb32=>g93_)bKg)EJ+U66#V;(U^B.R[Y-aBUffFC8,g:I<c<)B
\L+6X_:bOQ:^@LI9]_^OL;4=^a,;e(ec+0ADK#3_EU:PO-2_aJP.-5;?A&90DRVf
]T-T3J9QUZ>28ZI7f<=8F\4.[Wbac#a[+[H9^C&R-eVa&;1VB(BE#<UV\N/D4G;Q
.MZ@<)aXO5_P0_cXZ8f1-N^?+/,b7>^<767::T.80#@;Q3/b,<^6WEVYMde#OQ@\
f?G\SG[2P0P?7?>F?>4B^]#[XXEVDfPd^?[\d,Hg23A+^29RBIGOB+<fV[R?KbU/
g7&0GAV;@NPb318f:\^C6aW@)3G9MCH7)L?TM&B,aLL[U)A,Ce)NME6)1d&@]-b1
,^U05U1.4)DaZ14a>259Te^P>?d13-EY,-A:I6-Sfe4Q5R.J_>2R^8_.CVJNRJEd
MJDOK80J)WH1B/=Xb_/Y]-=<>bW(5d0W[V),cOBIIPb8L[[eE932JZd)T:b#9d3g
D7_GK\[MF.(b?LH[-R)?_-O-N^d+4Nag.A^Of.#[>&WK1F-b5_QZ_)MKg6a7g]NF
+L&6J<W\;J(Xb>J^-A\&1O2-2d<d7PX9&1Vb\+=1,/NEX=>-,Zg#Dgb\]@WeM/>X
)V)(TR(_<0<D(=HT57\WOT?T7O=fHI[Y_A:[.P^1C33RKR?+,IZ4T&=a-E^Q.H\d
09#6WQ1<M50^dM9;@d0T(<&RE4U@Id[1FCB:_#YPYPTQSB1N5S:V\KTN2;4PgCg^
JWBT0X10.?Q;#Q\A,aF,FCLMRW0U6Q;66B?TLR8:93G\KBc1>-Jg#]>E:Q#WKRb+
W0Xgf\_W?=(:W&3IFYG/:d6+]&)gTd[1N_.eWb2Je[1[g5gU6EgE4=R3<B7OBN2>
S2L,><bA@g=bMaCYJ-4S;VYbG?8I<K6H^>]/WX8aB^^L9g+&AQPZ/]6^JeR3P&b7
2CZX@<I\_f4C-)S-M.AUTS6N>AS5):gB13QIMN9SC-Z<JL4?J=9\98ECM&SPeIEL
9)A>YJ;@e^+#38-U;-_#&:UTTFS3ZLe4UX)7\3]A\)41c549:aOPI;.E]BF.<#_(
\e=_6ZU/CC<f<e2;OGQX-X66U;6B6a[;)ES_#Lf<3b:7e==1;IL@b+2KQaFA:LG;
/aEfUJ9TDa4LeD,9MfcGZJYIe(W>K+(a/6BAZdRF0@D+Z6T3>[f>EUd.<FZXbaa(
2QYG6_UYV@,Hd:6]:;#b9eIU?DMS+23SP:&+A5FVPDJTVQ>[a@Z:3_REW#Kf24E.
CX89CO0RM534IFdB>FHJ0LXECIf2V&N1E81#+5#aRZT2,T>1<,11G\-\QV[ZGU/X
4DSETJRKQ8/OF,8d9L53AV/cKBd6/>RbHA--e^\g=2^G1947LD8MD(?#70+1AIF]
>#W=a<][T.[UgY#(C;YX7RHd94EQM/J(3&KD4OO&1+JU6:B9,Y>gJU_S0ZX96Y/f
.=6V_F6<<AScVJNZ[<T2aTgKAgR:L>;#2^>RaU2=H=:0P@D[6HMQ+-ZTW1B7Z50?
a3&L07^d[LM:<L)F=L1Z;JJ46DOQ/VM?+L]f]#QK?TSRJaZc,4MAB+_>03,1;BO6
MI7EN]We/fA(?)0f3e?+[MX[F#HCCMG-9ZO/##d5?Q?Q+>c,VXeFYIc-4BZG6X:V
PDBEYg^+YY[-GL[VA^8JNMf_I4HOF@#8H\QSIBLR7dX7]X(>e=FdLEF5:H_1Zd5e
4?F+@?JgLg17X?AP^OB.fE/G6Xg\.1_?-YTE7/Q[:Q#,_(O>11[6A3Ve>#+ZOe)P
D<:2dcd0PDI,;/W_QX3_4K#02DEPY?DB6]=Y]6>e:UK+[HMfTSfg(9A1K<)\>DdY
de9PMf3b6g._\>1e31::^RL.D17](M6cT/g:2=74/S7+P0YbYSI)5b9O3\,5US4K
;<OLJ#KLK_72E[(E).Zf1P_85MD1\X#d<,eUKR7FI[7JP&ZHOYH,HQfR5NDIR4#5
LT[P^5G.aJIF3).B],4U6=aLH27TD.c&YcQ:_/3)=Y+JfHK3K^?X3S:-:+A2b_.(
:O>I?A3fU.?QXeZMC..E7F8g1\=:g+2XaNCRG,EV,X.+EZI6_4[BfWI4=,(3J0F.
(a(ZI+/X02[M5]WLILARYO6^16X8TF&,XDcH4M?A]MHWdW?V4]/GUC<KX0C;)S>/
2NB=V^[G.4;L\4:^fUV-ZD[A=CVM,-aT\M;e1;>fU;f#>bf2G_1CNFDFb+[])5P>
bAJE,()H3J.V>),01NdI>P>LOdbeHXMUeEYT4dA4cR.[M_a(OG4=b/HMSfcOFD<e
\[EVcFHK^\Z=_)3^K_E#;\fZc[9RJ5.;)^]1BEDQMc[>QCBQ7a;NAH89_?.HG/U8
D9e,4FX&NQQ^.U)XAAM4bbQV]C7_;ZdG;)G8KgWCCNBfIR>DP?HANPCbXS]0[4XT
+6cV#e1-5?Vg)N8]e)W7E?Xe2XJ>@8VLN^XMU_e\T4g:?;Vd1CeQ(2\PeCbYO(/)
/Sb8BfJ_<SYbc+f?IbfCA6<e,LbX;FG6]QA?gOCeM:L5GIQ.gg]R7@8[U#AT&NNT
5/7;P&S/>:I)18gO,-/?Mc730f4A;fA@[7a7@)d<5F&&X##2S+Q^5OER@Tf1;UA(
?-LZ>.(7RZ\]bUD-8A:=?;4O:SMR&,-ZTS-MFQ5[46.(?#c\6:,d+RR9HP<0-.XV
aE^b^fTW&SNgU3:L/fKLL,d@Cb9Y(TJX[JHAcK1MdTb#,BRcaT7BH[a,M<1KCc7C
ZAIN6-T?B,S+LXA=J-+3-R#K5JNf]?eFCO;&bA4NBZ@PS<Q+?G2<dKWC=+[T_-F.
VK.e+LRa?IQTF4LKbW/g&QH</BAOGIX[)OYO3]EGXU.9:=:Cg7S/T]3VGZ?&Q7^H
d:Q2Y])db-]Q2[(TQ@+Zb7&?LTWH?OMe^.;PW&4Z1676.GLN;0RJ5XEJZE5gTV;\
3R(e3?Z#/Z.Q9J7Z4e@;?;H_^d3XEOCXC9MUAF]@^bT(Q@M/c:JJ>R9[]>2&6VTY
bOG<P[91<,e5#=_1JWQ#b&LM<YeJW<O8[,0MNf-#Y7ea/+;Y730+&e5b3(P9&cKF
-XU\&=+3HH)HZ]>caY.U753K37bKP0A,G/P5;N&97_S/\B&D_OZ:YD/+0Q,^^I=Z
(UcIQR4Ef.#+/-,KHXNP.F4;S3ZEP[(PRKJ03@aBbS3ReY)YC^UG^g98OF?9X:f@
^b&BT@V)FZJ=VJYM8fH;bL?-J,5Vge+E)BUQa:UM7&</(01BO2^@((@NBc__?&-d
92c5F8cIP-CQEG.4#NGb#8Q\eMXN2fB,BC:MPfV>0]bYDNX1I+/G)XZgH:.Y<D?P
f,)RJ>Pe6[255WGY2CFJ[R_H&\c-/O:ATa<IcYI:(JY420Xc)Y>eg?EAZ@/<gIe/
=I1GAF@#TZ1fIf_:]]<K4c>0O>eM)VS5<E9(bO<AYA@C4?QI4c&P]_IAYTI308;d
_+@SCYd@NB9&A^MDN8bV\5fBL7C-<KGC_\H7^?FDBRC<(JOUL?L:>H;<NPYE&/;;
T8/[+O4cDA.gY7BfT(LRHMEM?9bIX-IJ=G#g=YES[U1H:Q^-14??5^P/0f3S10^F
0P49I9+TDL)?b;Q9^&#1R)HLZ#c>3VQWO/?e6,P9bN_Z]00616Q,<S+\>_-^VfEd
7:U;=C20O#e>ETA/EKK5S\,fbG/(2bNTXJVA)^+C<<7g5&g1Y_ERWa/12H1T&[S0
NY)TUFLHAMD\^F@LDD9?g&?ZU_OZU#[_a,;2)Ie\TeD>.Fa,K6P#;2cDB.?3QOZ=
&g0H,L>dN;6KHUaW++G?X^)01Od[)LR97L(gAe::bK1c@Yf0N]#Q26UD2C[=T\OL
2W[+6E7b0f+4(A10084D7OJZ82b^]b/C4VI_bU[B9X+2]ZB_//0\;CCaZDJGXK\N
bO95M[7C>&5:8G5A;:ZDOT=NWaN51&>^T+9O:L@OgQ^_Ab;JbXgNA?9JM3DHQAef
V;?54#<D-Nb?6F_EOf;eUG1gJ[XH[I6]P/LW+7Y?<4\S1UN:/:I[#DS7=[.Gf<T8
@POC4@7EO-DY6KYKd=4;^]f<;d.D3].[(3H;]3]e&@,V].NSRQ63N-H63Z8=O8b6
?(X>GgW(2-^/:0BQ7L4a(Q^bbSJ:/89GF-R-C97Sb\5FP?PH7.Ue5[F/2M3b/<fK
4@GBbG[OE/?gU@\IJTA5:4L7J>E25/CJ,EZZ+,4;YcAeV^W6Z]#&6D,df@(gLQaY
eHKJV[P5faM.7G+\&]39I369Ne(+1^IVH-T\.;Fg@XgJ)@(20=Wd=+PcLLTY9KI:
aZ32NKNN2PaLE6AJ:WN7T9Z;d#RGL,0>bF3.6YAK7(J@gMe(.aG844c.DIJa1TbW
;,KVg1dYHS:HD+_&G5^0[g:da4fTSUFX9dEW//g5;O,-T5:gK[ZeBFF6adB6d,#;
UFDP5Y9(U8?V]XVf(V_=HYIJL,>YJfC+Dbf9IA)B=.eH5eYNS64TTa/ES?P1egFV
-Ag1]D(7]7WN=,gA_K<V])KG]2H/E.[2@E-0H;Ga(3/fa2gEf/72XKQfJJ_OAD8b
Qg/8e8Q63<;\c]\^a3IdbYF8;OdB13(K#FBP(HaY7g:5(3.HGg2V6&a8\H1#IIYM
E3+Q8@R7YBYH6IbLOLgQ3+RVbCf60O8f.2@.)GRBf]=-#J0DRdFZ0W_)8RWHNO(N
ZYFJ[49A^PT?=MCB(D\YE3_Zd\CBAY<f4BEF.L8aLKTd^8M^5@B_A0Ve?GVTOOM9
bDYG_([@MBVQXd+)BKJU;)B[@DSG=1aDK&XCU<TJ=Z+CeW,:&:61]>AZ3PZCddEV
CgI;Fdb89B-G;B0T8#I3(0a(SKSdaWG7;G.\5ODf5T[Z8]FCY;c;6]O><R:EcXc^
Gc-f=(\#:,+06>e;9&bgeEM^O->VE31^dX;TH4WD01X_Q8XEZFf^+Wa:Q3X:Va35
6>#;C+/,6MeECJ:,;O6g0-IP1-/&<&/(8CAF+4U)F,I9NQ/3D&C)Vc<<M0UUW])a
/W:3R:U5KeYVU<d4HY=VU#Y@T2IP>FP+R?/OK(O,gMGV/U6SY>WNS-I<TU>eYT.-
AH4eHS0G9B2<c+A;QaH#^;]ba#g;I8#=B?IJ=W/-1b[9.GTLPK4HB=MMLQ@cBJE9
C[)N[(UU:Z9+)C7MM5Q5=YA.TKIc1aWX_]YH^BMR6Ud-bOUBOcL]Z15L):IZW(//
Y5UQAL57L\1&f5f^S+N;SPcE4I2)S7#OHDcVUWQVL2]?19&985Qb0B8=^7-6C5>F
4e04ca#67UKRWK[GD/g9>NI&c:I=F/b8/LLFJW:AFcQR(T2BYBPK_)=ec/:G(BWZ
KCB7B8Ib6V2=LK88+dG7g=\^:>.EV/a99\c6QP60Y0]RWHI@8;41<EX=2R1WgS:-
gMcB.-NO+I><>RI2L.6WX27Gb-_I&5Y^_e7&;\Ra8F]VA8+XMT7\T,)K_eNL3+3?
X1A/V^D+?&K=&+KQ(-/<[]//HGfdVGSZa@cb40_a;e8RL9&C@.KfBPUV6)PbEWZY
MTdLA(6\Ga(O;G1gP&#1[K^c&\3YO/\4bG4:Df@>#[\XV+I)Ub,GG)P_H>Y)CfVcU$
`endprotected

`protected
@V=aJ5c>^=@UY6ME]eA#ACQF#d.<g1U.V^6HaUf08\0;94KaQAO62)_/IK]H2D70
E-c/,B.^Jg+OI=0W2JXQ1)QF1$
`endprotected
        
//vcs_vip_protect
`protected
Y0F7XXA)Agf1^Z#.4bT0K)ZH_^51BA;)ZH_]G(9,X/\4fSH?U;N;((APTE:<7L;-
b?TT<[62Z0a\DfD5]G_>=^XB=,>MeZ&B2\\_6PfZ.BJK5Zeg>?dOXJE3OE#)eTGV
@aZZ+^\348C2?J4TZ+9]D4VKZNS]C9+.J]&;7)79DGeUS4=2G86\Y.MT-_/74NM=
a5(GBVS>4KHI5AD?V_X#,DS<K--_CRGVL7J&B/0;Y&/&U)61cSdM\YK9Ic5V5YDa
VBRa&)X-CTX:(V\_>DJ,aI44Z9\Y3/ZL;I7\4+g;QL2f(deU36=d3EJ<NRWK-ECH
RH(K]E:2R,a&A-AV1PCN2SD^I3:aJWB\^dV/.VCfPc:A2&Q0D+&)Q9K5_TabVa<U
6<^ScK7Wf\D2Ya;#.BfAad=<H;PR7/OZI_DOKO(93O,Q4M.ZLc,63P3Tb[b3^^bF
^DcgI7@_PEWD55B(gJR,3;71_/\.)Z92/QY:87Q8+.)Z0+9K.^0BC?AeQ-YH]<?V
ed[J6HC7(LOeCBEPTL(3bEb>@B.<\9;(]6^W,8\SFYD/5c^L>W/,;4.-aL^)W5K6
-QJaH5.ad4#KM?;NbbT1/6PK^O5I+Y9-PK/<8Z+_7A+CMA#c9K<d@YH(WD9[X\TF
f))EB,TE4:bX=JO4>@N\&06QXb)fR35T5.D/&K=89Gb7Y2;.#W0#J0Xb?<MMI09I
_\O3cZZWI#dX-VQT^BJ5LJ/.[g1VAYbU&QG-2U;d#ZEI].,Z.E^,GA>98#:GUTIS
->f_NEDY81HFD(?<cFW/S_4a#e:K]4).WJRfW;0A7MHEG\>.8gIL(gd=9[-C9#;@
DO/(?(Q#(83#Y0/ML&(EU1)G]-D#d\X>\BcA[ZbJ<[^L42S&U+63D&((4&ZZZ1Hg
01aJcN[d\JT12,,Y84KB?d;<X&2@=)@]>7TDRT:=L/e#f_M-_\[L0dPM>2N[ZS)a
:cO61)ab=/Q(aEU9[WDEP+=eBMfG?5f1339=&;(CY3\HZH]D@-NQ=,&Gcc,X+++_
69O>+F5e_V.Tg:<YJYZJ<?YDTfN#TDDXQ9)@VH[=GF-ES4d&e:MX&NR)B-91+PYg
W8Q8fL+4#H^50b<=;DGC-VOLa&C-V@8.Z/1D0;VR,DDL6Y)XOJ[HY6/O416:[-,_
?(4JOPSOCEK2#]Ld]5]aGWS+b0YBVTbfd8][M]S[E.dN/I#4A(/=:QN>4(2UGG0c
OHY\N)b;B3c;>[?Oad/G,XA)/70;3E9//XHFD)SI9DB21D4S45eV&a=3fKg4[_JQ
dYK7a8E_;SN@RX>-2>SU\4A)5$
`endprotected

  
  /** Populates ace_ports and ace_lite_ports arrays using system configuration */
  function void svt_axi_ace_master_base_virtual_sequence::pre_randomize();
`protected
O6BG>f-])D&CT+(TY/0\O?D01dSW>S&/7:FA(M+TGRJBO2GEGNW23)J>/KQFJ?)a
\.:(7;1CQ>0\TS?957YI0GP/[J@gaZ4&dC\7Y[H^RF=XN3b=>fB4>c]S?72:XI/K
^bbYN6B:fbSXY-O.Ac]Y)?,O?8^)17HaYcRU^H]A?WOQOc7)QT]-OY^#_6&?BfD?
ZKfMWcFeA_,)PW3.b3E9L3:5?X1]T:+eCVJ4,.)T\C#]:PIA2CS6gH8YcO3#]04G
Z@b65f7J,JN9=.0>AaYT?_+P,ES47ebfR--5.V[+XRS]()G3^0]G,4,SFR1P<3>C
&7Z;[5Vf/(04^_26[:M4/Z_ZFOA3dcbO^P.[V7->g\5NF-/VLBcWB@Y_&PP5<bPB
;M2a=D.VLQ:Q,Gc2AG3#?Y_Z1$
`endprotected
    
  endfunction

`protected
4RC?Sef^#\Q,VUC-d@,3[4fE?JDdF#<Fd6_0&T6/fM,L[-8W59XC1)caX]<eGgHb
;<_B@N=[6U>+A];KbNUJ7ZO/KRE_J^<EdZRd^Ef--2EcQOU=3#Y-<PJI4RDFF.60
N:fJ6;R^B:f3PeL)IZ23=gEb=aQdJ+[):U_/c>aR_cK(H)5B6f\0M_KdGf6YE),)
ZPPF981.#NDPgg3Se]]MU^2Xaa0R-QQ=gX&g<I38FN:2[>c(6E:/[>^)3?Xf)U&V
f;,=WBJCJFA#KT)A:;1FH02K0,=MQZF(Q)Ce8@HXRadda<SYC:0c22/bd#5VTIPT
>]-0KTIEAX<)B[#7^-0QA)CJ6>-faE:ERI:_UW16UB2RP&HQL?O]5AU@:UNC<c?V
\0Og)_#.;0a8cR>NDfcMBZN-4#gDAMP#JfgK>McJTSO&Je-S)5TJcM+G-.2YBbg0
Q]LHL@;V#E6/gcEU6EJcP4A[XbKJH^M5c2=ZL\\C-_&6KCXUW#Y+Rg;6/YXF955F
B)/?R0/NECRS-S8FRU7f;;X_7IL2AdfGF#RGR<7N<))OO/g8<cX(99)CA(=>:E2N
7Za[5>7WL:IA8IFE[14ZGYRK1D<Dge;Rf+L26>EH1-_:JI^[JQ+[UH0[_9RMQJ[2
A1)Q1P25RE8F1/)0ObQP^BPVNF/Y<Q0S&K<1UA8YJ:HAIbC_6]5EUfHVMdA>fQ[D
;Z3[edC;.gdRdgI]RRME;QJ2[FMBR_//]V_a3\,>ZV<^RAW&AWFK0.fe>[V]WVcG
0>4d>#(gOQ=&Z86?EK\\7OHIc>/BKM6W\P.@<Jb;Nb=OYK+IQG.<IfMV(e#6B,\A
:LJeOW<e5bW#4#.Kc?P4902NgYc1]Ee;#[VA=&K5=ZM)Q.\^_\O8+0aB<4(WDga2
Q3EIO_@U0997(Q7PPGJ\U<dY\3;KLU@TZDNaI>]UC>KP];8U8=^A=E:@c>d.?P_[
NJ:a+0@5B/H\OK;57fM-:/JCD0P&OMWD^NCY=8HT88-D&?[7V-NBFUe[f2gg#NMN
[2W;@:];.)LA8_BfR]IWH/0JA1L?G7HDKVW9)_ES<.C]Z/a6LN0-F>RDQ9#[X7LE
UAI?)[NFQ4Y54Z#a:0^9EKGV0;JUN>/RMSP288=D&614Y[SE=CY5g]#RAJ)>G/4-
.ZSXB(4B(:aY,#H/@D_)B#cD.(QfYU6JePOUFOgf-Ib6CMX?-c7DI92UG_7#3-NV
_Uc4Z_E4TKERXdWeP--d.4U=[fP,[K[4_76F78\(\\VUYT[DV^3&=P:MZc,CCf\Q
+<0Ia&d+@)NQ7C4AbdgRf?(-3FWHT4]2(JRf_D@>+#9_;BN8DLR,g[VJO+I&<F4U
5&/?PO^_E:@+XU1#IFCD3&U1TN)HP/abJ+M=#.@Oc\NLP\gOD?[,6aFI5Z(,U9g_
>4ad@)UBLdE+=RI4g0\IZ\2Y+\78@\R=7I=IcMUQAW^6RNcg_7ee<V3C:U:1Z56C
NQ7)V70FUKeAD,Y&TVf+4<J_B](442/ND,S<Uc=K<Z?dOTXJb8^VCD=A<,A2(g)B
^7.GWMCON\?1[d@J#F,^#@3S1.)5,/HM&.2XZ<SQXSb,9@L9?0VT/5V\P132&7(0
]T_Q3-;f/^=25C,=W.22&/Zg;<fCD@B&d_]-N12Q<,)S@@RDYJC1;Z81,[gAF^V5
_Z+.:9&HgQ]S<OV8dCWI-^T;B02ZRAgK6>]O8K)c_c;dT;&LR&L#R1g[>a0\]>_O
X:_WON86SSO/FH+\)&4?Yb@(3K(RX+CB,;BMe8T[C.U5)(Y91+;))Q]VdEg0UOG(
I>38@RG\OM[g&Q69Dc_++X_]2\YXQGT-6KK-7-#>\@=WI9LE@&P+E;ISG+=DO)A9
63<,YaC@8(bJE=M/ZKV9Z(C=96TGXU1BQ?f7V2b3acYWQ>:7#Q+<8@[V#Fd;E6YA
E&I[:G<LBaN)>SQb8JG/c#Vg&e@MJ\N-SHcVg)ZCKC[f.H=)=;_BU(#A-D;K&2FO
WQ3J7S0OJe>>Z)8J5F(KOc3EEG\-_(L@?Y5Ya[UI4&_<T46IL[R<]a/(NbX&Ea8S
C0]@RUO.8,6/Z_=(T7Y5\bPA.#@/0IXN&e.Dc1&-9=c:(::fA7QK..YI>LE-d/>P
=c]3@6;_?D^DL2KaDZB.X[FaG00;PIP;I]STPRW9.?acCAHU_^Z1?QP6@N](P;,+
Q/gDHXP2/UYF>^B6#J1R90B)aeG_9IVV.PHA8I-D@+WR>cYF22?@HQ>[e,.8)>D-
_H0^-GEGJeF6FL<e@.JQRH6N?#@3Q]1O)D_WJVF/;K<fK]ZLg?BZ_XZ>6M,)e[,D
7VTULO<MH>7L9c(0a(>@5Kg&]=f]c[(T_6NJ[5Wb.B5=4CI+7R+4A1]_a?eaJc/+
WQBP2^62XeCeafGdG93<_M?BfZ](.ZDIZ:3Ba5f;7Hc-4fDS^^Z0Q_F8=e5Q+.(\
PQF_))I>R(VLN4&f4g1-.GD4]c:MW,-:<T\EB6#W8/T2^76TK8XLM;LV.BQ,c.Ze
\?NO+KfUOfIZK1:/=3S<T(8\9=>F+X1^3BR2DI2Z&gH?TY#g;XUM829:aB<3]S.^
&X06=(b12(gG15Lc)\@AV8@S&8SR6NeCPKR.Hb^5-6YY:J2C_/K6/3LI<)Tbf.c+
[d5d1@?M^_<;U-EV13f00O9K1B1K+0;_f\A.c>d9?fC^gbc?>+A#PE<_DZ^DTR<&
XcB]LcTT.+b=7G,HW-ODF-0V[aABgB^ac3[;LF//LfA94;7;]KI9Ng=^]1?g+H1O
[c5+ePgJK)8;[ScI9a1ad+;MB4G--fPJ3.Ff\A?3R2HcO>?C=2d#3.GMc6E+J;0e
YLHNS]77O0]C:99cF/SM@UV)f:(-6GQ0<,KHRdVL;BIDa?)U.OYI.3,H(<)#9YPf
C_<CA./QQgMH<@>M\.N?KH(5J-Q[6.QMNeGe0UH=g^65TZH&CfUFc^\1T:Z_,,RZ
-@^#YgS3gQS;OG3#D#ZBFT&5YZO-(GZ@T-Je1M1bC48dW9[fb:YA>4.abSLg+:5;
:ETUPMH/F)ARUZ61cLY#J0#-=7R3>X,WQ+CW>WPM>ROR2C,UcT,4]1^T@2-GTVJE
_&]>dUHO,@0S3Q(_Q<R9A?f/7N)b-H@N\A[abeb=gcg.18V6F2FIS5?O3?g/,UUc
EB#Vc38.?V6]=F=af534P;^]4ED/YVJaff;N/2Sb=IZO=UKaR_H(;4:4<d/_Mg6A
a<A2()>-c<<ZJ//JH9c]7Ca0]=VPKfLfOBNY]0@VCMT0_4N@H7g[->fQ,XO-4/Y-
9_#^)0Ba/Edc5)52MS)\C\6LR/7aaG+CegIT1HHZ_XP.=0Q^dXf3,2J+A/XdW5U-
a](8-<g@-=,Z+61BfJ#^EM#1_3@NJ]RADXb84R_,C-UTHTRWPXJb;0IK<?KBVMa,
0UIE6)4THIBXM[aSNgd6>@IG)bf@a?/XD..RC953K@<?dT--DXX:QO7<VO(K+IVb
@J(@bUG5dQ59K+9B-UR16,FSGJ/#O@^0;^-4:YJ/L#=&<4N_9P<b0K-J#GY)\R;[
+a<7B)RgP7JZGOg0^Pd7YKTWPaWY(OARc\HM8)Y7F^g&&J;K7:H8EU<T-TM];CDR
YKZJSYTI3gCCFR0-8FY==V^9c0;<Y36\\YJG:XMN[3_;:HUK=#0)?+:G^QLSS,:Q
^A/Qe?Rb@OU/4U<S4##6[fTK^XRc3f:6=;U2+e4/@g:HTgN?VV_g1\/:EU\,6>3d
b7<HA(UgMDT])g<S:FB\IS2+Wg&QTdB(V/5RaW?SW4Ua:1E?,=DAd_\,#3[OEJVW
L(b[Y:[PVQ;4WS/RA]+O/cG9;3</W1VGY,-K[=UCYdNW?W67CIG<]<L[QRe+Z^g[
<2YJ2aKG=W?SEIG#[b#3,\YFbECfUP212b<:58a6A,?)I5)4-5+R;97CAJ4>D\.O
@c01:Z3D@H&][g)e#7R_f5b_d_Hb6gX&8R@e+Y\A>a^UXf0P6IKg_,(We?25.I+G
W&[)<,W0&.VW#M8=@53)9&<?+eNd1I_bWc--8f4,=R0Wf]@64_RI3-f]L,KBO6Cg
EYPgbAK7X4=R-2.[;L^3+M9fa@b/WaB[#]MV#A>Lg6NEEFX-JC[V[NXZ9d<I[;-N
)7>;c5<L]aKVU(-^[C:_P8T;1/2<MY3=g<D85&[R&2ETW^_X4\)X^=5d,-.SMF#F
0.)EHN+?64a\;bU,cdEP,W,C353b[RN=[G7Z=K==Q>XC2b@Jb,,0^5LES@-G+QPQ
bS21GP\49C>-QN^GFO?6,7C0(&3T@^Md@E,Y]OY:gf-UFV7T4]+H#ZD8-)eabV2>
J)X>86<2Ka/C5>-HGJaJJTb&H.a0a-fP>2@[B=K>&_@?PED2&:Q3DGT(F[_E=VRd
@ESeLe_IAQ[Vb]UWf4B5FH]2B1=/6c_0e,<AIFeFe]aX-ATG=IAZcD5>c7WgLRE1
&.:M9N0d_O\F#4ZD_DF<#eV&/T-a=:_F@Y6,R[dYdWdD]MeO997JG/(M,HZg5Y91
RMY;63P8U]cJOB<)-eeK-1K[>4U=VdG\A-S@a<B(\@-1VTKX1#W#5+#]4U_(Zed9
(,a19c@-2&gTfL]H<-G5abSZYVg[\Y_NCBYOD3Q<++XF3E6OgXJa&^[_/@Y,]AcS
GG=;Dd0A)Q-e0518X[V[_LW86=(DH(OIOZ:W>FQI\fGAM7?ARB#9XgT)+0f_fNM-
P1T5#6/f\5FND1U1a:abHNDZA+efF#KXXbS\.OHfBLXH2QaTKMJ9#cOJMCNf]LQ7
J8gB1dNK836/>3:IEWNFXE0^+39-fe^/7K3_JH>\V#I10e)[GZ,b#I8T3LYgb\=L
11H<7[\VTf^EP_cX-\U8aV1ZS7Md3VOgZ1I/9=F#@QY0ID9;@Q.ZB7AF\ZHB5bb0
[Ce:DR9g+7VQf_3V/C6c::;Y])bVYCY[ZT..7&6^=:ZFUBIIQF_a04;OG44QfaKg
4AZ>^C48T#/AW=CX)FK85R[ILOE_42P)08I>Z&01L)@K+ggK<V(fDS>Z@-1)8<9d
]+4gGQ2F1SR67.Q(T7?-.eBa6JI9+V&Rc@K?_F?cS-T:9K];2KP:V:=6g0N97bd3
R(e]<K1N-((7]144Q-7&D<>efKaVNe+@CD?:2(OCgJ1ECL);&4J_HYA3VMLA?beY
H8Wag5c&X_7I1cPd:^3/]L/+09TgK\6a:D):YCZ0SG(-,PO>;5[H#2V51dd;dT<(
P6T2=<Gf5E\2,ZXQBNb)_,=XDEWB:B;9095e84dSF?05bZIW,f)X.^)+(A,fF+6=
=VG?N8^]8\:G=-50cHTQK@f@;#)AeF1E74N=VU7N,e.c^R3:f,BXWSA^#Ze1Z_Z]
7&GL1A143_A60EN;E:]D?Je-57UTRCC..==D<MT:<Q#RRVR,13)JNS4Z#L0#[6VL
aW4fN@cW#B@/ZD1\_9VZdSfWALdA3Ob2;P_8.3]E[+KF3UWe&DMCfXJgTF8-c8A>
]a4-3e2X&2=:]7^+&9S:HR>#QF2&E5#fH@Jc78A89)K^UH9?bU/TNf=Y,2LZF+GC
O3[@+V=:<>-7+9#-ED@O8fBY]]\LO8Ie23M@N[a?P[N?KWea5[-+WWNV1Z&5FDb(
(FSBK-:Y&bY]-d968:)?FVJD5H(<8>C)MC+@7N?FPY@Q.O2UPHf:9;31N?V108MK
d,2@YV:ZV#4F#/8KKT.CI-e\MCKP@A^CK&d[fX2Y;-K=8=(I.G=5AOE-)I7N:8K+
QVMO;.H->e;:G+GJVN/DZ_f^)Ke<(,f[K]YX+?fNT>Jf^Eg8ML-OHH:[]KJ<Db.-
VA,X9L.9==@J=FEL^eGD]R84ZY3NN(1eZE_SK>4)4\Nf#bC)d?bO(Z0LJbb4Va.#
J.X>S<M/MI54CH&KJT@LLP:5MNZB395:6C=_>9f\BS0J;Eg@.Bd_)37)0O8_Z>)1
XH+Ib^K19M2aJ(]#f&ECXK#O23VM&<.cVB/efL8G=-08MQ7I.AMG.0A.eUQgG6<8
cU6VD?P)E9f#d(HYD+53)^[K^G[\b5V0CI1]\(OY#DSRdA(S,@#A1gMU8d]9WUVZ
_=@(Z/.YbHb:1N_>.d6SBY>A,C26ZB<0MP\&X;>CP1;D[YTgK1CMa)>bDRE_DgA>
Z:FKCIa,[U6cVB(]_;E2Y,4gM.^Y(.E0>NA<Nc]\J\)3aZd[4I&1/Wb3gC?2K2C:
UQOA(eRQ/,;]&=Wd]B3C>?7C3f-LBL,?=Ab&=&8OPXgQe5ZO3gVUM1VXBE<DM1#H
5B#(B1K(K6R;a\4/)6C03-4C;91J:(KUfRaZXJ1IP9e2GGMg1P>3)c6S,2R-9f1\
U,5C8V^6?FUD9[fbT#4Ee3&>DRR?@,R/VQBb8I;c7<I77,>K9S:?B^X4MC+E<A+6
dSg2K][:>:T&XMR:RN)IKBU\H(gPg-5YMad\geY>KR3>g8/N7PR-e3,A,KWKFRbX
X2f@7aDbaRBL&P\_g:-<1aKc)cZU6?=-@0(@MKgD^4UdU6C3=3.dQ1,71;MM_AR>
5c[_-199D>I#>V0BFSKXV#O3OD)8f+DB9,ed?STUQN9#:U98P:EeIEMRHFIZU[T&
V:fLCE/@0;)DIP5C0=Y-AG:IaQb=eb04bMaM;gG#ag_#fIJOEd4^+C_2\P_W@RbB
VH(JF8b(TJL^ZH@6FZ/,H]K/5c/,b88\129#VLBg:D)fX;[e3@EJL(;D0BY&S>I9
Q#PN01A]01<Z;XL6-0U>2ZdfC:JW__<NQdbT@]\N;DHKZaW#9,3GUIEX:NJdE>3N
&>/209.R+LUHI][I#cYDG=7RE24UCgfRQS3V=2.PPK-_4Y<;,YXY,<9?WEGRFL-g
IK#BC+E=D+9F0BJ6)Ref?=&UG__DP3.B[/)3L&cI01c82Ha),.@37=Y057F<N]c]
HN.U[G6O>,e\9^+SGfXR:8_>V\gFW?60VX9W0]4&9:dc)/YS-DT^I8.Kb(-5Z#G7
;=<?)@=/f6&WO/-XPO?M_P:+@[?dK#A.cCgPM6+b/Xg84#P7NO85@Na05/C<Y_?9
E3\4>d[EA&eT+J\^[7_9;.L+c<8\;67Dd=A:D(3(.-/gHS=.[2P/^cGZ@N3ZG8?U
(G88RcWAS3:+1&U5aY^^>W7dSTY3eZ2I(8I9/R81aN/W8?RE##DFfGVP9;#;A3>e
S6AGH>U^3?:Q-CWSeS_2KC>D6[b-\B9\[FYR,Pa4I<3,EFKJKW).7BOBRX-RO_3/
f5XD2Q@E/>(Lf@45)_34>.f;@1Q.1QQDV>0?@LaJ[R9=7K>cG+.Cc[b5KV8#GC5_
-TfcY7,gA.D-HF#J;e1UT&<S=c&g4]A7:cU:HOQ_1S>Re#Z:b)K[bAW<NCWLMY^.
;abdRUH9O1e<E:K#gW);8RK@@,H/0M(E7\DB,d_fZI>F339C/]YgB)S2DB+-VR&=
8PK/C_F9HJY/GZ-LR;KC1fYD+L_RDN?UM<e>dLE0Z(\#>JY2Q,WN;UeXbaW:?J+4
9T9G]Lc+Q-O:+Gf9T(5W3(J6U_:0<&=T(X-/g#8c3HA.Q:Q7M4HOV0/_-7<U#0e0
G#2?L@PQ@;5MZR\X=MXR:3O35>8W)K\<B3cY32;WV<2P6#e3@&=9;+TgFI_?--OO
-J4A#Yad3A6_ZKODCaKf.\?5W3e@9:YY?1Z[[e.gg3U>)2108cbQNWT12N<,U1;N
TY7\+GE_3.ANV>(PH6_[g7BTE^,\G2/,\.)0H),/2G#BXgZf0<HYXTB:6F2-#)1F
XN-?3BG/3TU6G:QM30CD/.:L.-SO66LH0]G8\c8U4(.U8PMa_E2QVbWbOW&X3Aa2
D(?AJB;<Je3&)+c-B)VYOL=>]4]WcHGP/4fc^e568.&NWIVU7:]4LKG@.0V.GS7A
(bQgNWd?dC(KFJS,?@-R#K:L1YWXeRCL_?Y:a@N1U8@gL3D5P@?IdR1XH5P#L9Q1
YM)1@E;/?/(,ZC8#P9VBL.1B4:?D[)ZRFF<Hc)2H=LY&EeGSX?6D&/gccac]LdTd
/6.W1VD7^<^H/aEID;7J[AXQ]dSO(?()+XHQJ)SYCJP<@&UE3Tf10g&11RHNbZD\
e#X-]Ib]dK8T7>ICS@/=+BATgTc=^Vd+#OJIGM:IMI-:4>5CU[WAYB=-4KFTB>dY
Z0+(WUXB=T^_MK]2MQ6LB]G.N6WI0Rb;QM+I9]27D8NKKZJ.])aT3KEREX9)L7\&
)S[SP#.&1Y=eaLLVES-g9U1(#-H1(Q4JgPT1OK9Le+TG?0aOTf8;^GDK:[(KADY+
D/\A>5e71)e+X/@6g=MIgXTBB:FUFA^IRBg&EI,RgfO5),8IVCN<QDOAIU^V4NKC
GIa4a0/(;AZF?3YSKUJP;EgMJZ5ZK=R.[47Y)L[M.0P^._@X4I;]L)f(\[Q6gEHb
($
`endprotected
  
// =============================================================================
/** 
 * This sequence initializes the cache line of all masters.
 * This is done by:
 * Initiating MakeUnique from 'initiating masters sequencer'
 * Initiating Writeclean for some cachelines of masters.
 * Initiating ReadShared from rest of ports that are ACE. 
 * If use_parent_sequence_params is set, this sequence initializes all
 * the addresses of transactions in the parent sequence. If not set,
 * it initializes the address given in init_addr
 */

class svt_axi_cacheline_initialization extends svt_axi_ace_master_base_virtual_sequence; 

  /** The transaction corresponding to which cache line initialization needs to be done */
  svt_axi_master_transaction master_xact;


  /** port_id of master_xact */
  local int port_id;

  /** Base sequence used internaly to initialize cache */
  svt_axi_ace_master_base_sequence  basic_makeunique,basic_readshared;

  /** A sequence that generates WRITEBACK for a full cacheline */
  svt_axi_basic_writeclean_full_cacheline basic_writeclean;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_cacheline_initialization)

  function new(string name = "svt_axi_cacheline_initialization");
    super.new(name);
  endfunction

  /**
   * Initiates MakeUnique from 'initiating masters sequencer'
   * May initiates writeclean based on random properties
   * Initiates ReadShared from rest subsequencers
   * May invalidate cacheline across masters based on random properties
   */
  virtual task body();
    `SVT_XVM(object) base_obj;
    /** The address which needs to be initialized. */
    bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] init_addresses[$];
    bit status = 0;
    int target_port_id = -1;
    int last_readshared_port = 0;
    // Populates master_xacts from parent
    super.body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "bypass_invalidation", bypass_invalidation);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".bypass_invalidation"}, bypass_invalidation);
`endif
    if (bypass_invalidation)
      `svt_xvm_debug("cacheline_initialization","bypass_invalidation is passed from test");

    if (master_xact == null) begin
      `svt_xvm_fatal("cacheline_initialization","master_xact is null. Cannot proceed. Please provide a valid master transaction to the master_xact property of this sequence");
    end
    else if (
              (master_xact.coherent_xact_type == svt_axi_transaction::WRITENOSNOOP) ||
              (master_xact.coherent_xact_type == svt_axi_transaction::READNOSNOOP) 
            ) begin
      `svt_xvm_debug("cacheline_initialization",{`SVT_AXI_PRINT_PREFIX1(master_xact),$sformatf("Cacheline initialization for non-coherent transactions will not be done")});
    end
    else begin
      port_id = master_xact.port_cfg.port_id;
      if (
            (master_xact.coherent_xact_type == svt_axi_transaction::READONCE) ||
            (master_xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUE) 
         )
        void'(master_xact.get_expected_snoop_addr(init_addresses));
      else
        init_addresses.push_back(master_xact.addr);
    end
    if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      target_port_id = port_id;
    else 
    begin
      for (int i = 0; i < cfg.num_masters; i++) begin
        if ((cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
            cfg.master_cfg[i].is_active &&
            (cfg.is_participating(i))) begin
          target_port_id = i;
          break;
        end
      end
    end
    foreach (init_addresses[i]) begin : tag_foreach_addr
      if (target_port_id != -1) begin
        bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] init_addr = init_addresses[i];
        // Get cachelines on target_port_id to UD
        send_makeunique_xact(target_port_id,init_addr);
        // All cachelines must be UC
        if ((master_xact.coherent_xact_type == svt_axi_transaction::WRITEEVICT) ||
            (master_xact.coherent_xact_type == svt_axi_transaction::EVICT)) begin
          bit makeclean = 1; // Indicates we always want to make the line clean
          send_writeclean_on_rand_cachelines(target_port_id,init_addr,makeclean);
        end
        // For WRITEBACK, WRITECLEAN transactions, cachelines must be in dirty state.
        // So don't change the cache line state from UD to other states. 
        else if (
             !(
          (master_xact.coherent_xact_type == svt_axi_transaction::WRITEBACK) ||
          (master_xact.coherent_xact_type == svt_axi_transaction::WRITECLEAN) ||
          (master_xact.coherent_xact_type == svt_axi_transaction::WRITEEVICT) 
        )
      ) begin
          // We may have situations where there are no other AXI_ACE ports in the
          // system other than target_port_id (from which we can initiate readshared transactions). 
          // Initiating WRITECLEAN for some cachelines from target_port_id 
          // will help in moving some of the cachelines to a clean state (which after the makeunique is in UD state).
          //send_writeclean_on_rand_cachelines(target_port_id,init_addr);
          // Invoke ReadShared sequence in other subsequencers
          // Cachelines of all masters will be UD,SD,SD or SC states.
          send_readshared_xact(target_port_id,init_addr,last_readshared_port);
          // Invalidate some random cachelines in all masters.
          if (!bypass_invalidation)
            invalidate_rand_cachelines(init_addr,last_readshared_port);
          if ((master_xact.coherent_xact_type == svt_axi_transaction::WRITEUNIQUE) ||
              (master_xact.coherent_xact_type == svt_axi_transaction::WRITELINEUNIQUE)) begin
            // If the cacheline is in a dirty state, make it clean by sending a writeclean
            // This is because for WRITEUNIQUE and WRITELINEUNIQUE, the start states are I,SC or UC
            if(cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
              bit is_unique,is_clean,makeclean;
              if(get_cache_status(port_id,init_addr,is_unique,is_clean) && !is_clean) begin
                makeclean = 1; //WRITECLEAN is always sent (not rand)
                send_writeclean_on_rand_cachelines(port_id,init_addr,makeclean);
              end
            end
          end
          // If speculative read is not set, invalidate cache lines from the target port,
          // if the port_id is AXI_ACE
          else if (!cfg.master_cfg[port_id].speculative_read_enable && 
                   cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
            // For these transactions, either a non-invalid state is allowed or
            // the VIP initiates transactions to bring it to invalid state
            if (
                 (master_xact.coherent_xact_type != svt_axi_transaction::CLEANINVALID) &&
                 (master_xact.coherent_xact_type != svt_axi_transaction::CLEANSHARED) &&
                 (master_xact.coherent_xact_type != svt_axi_transaction::CLEANUNIQUE) &&
                 (master_xact.coherent_xact_type != svt_axi_transaction::MAKEINVALID) 
               )
              send_invalidate_xact(target_port_id,init_addr);
          end
        end
      end
      else begin
        `svt_xvm_debug("cacheline_initialization", "There are no AXI_ACE ports in the system. Not executing sequence");
      end
    end : tag_foreach_addr
  endtask: body

  /** Sends makeunique transaction on the specified port for the specified address */
  task send_makeunique_xact(int target_port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    `svt_xvm_create_on(basic_makeunique, p_sequencer.master_sequencer[target_port_id])
    basic_makeunique.makeunique_wt = 1;
    basic_makeunique.directed_addr_mailbox.put(addr);
    void'(basic_makeunique.randomize with {use_directed_addr == 1;sequence_length==1;});
    basic_makeunique.start(p_sequencer.master_sequencer[target_port_id]);
    // Wait for MakeUnique transactions to finish
    basic_makeunique.wait_for_active_xacts_to_end();
  endtask

  /** Sends writeclean transaction on the specified port for the specified
   * address if do_writeclean is randomized to 1. There is 33% probability that
   * this will occur
   */
  task send_writeclean_on_rand_cachelines(int target_port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,bit makeclean = 0);
    bit do_writeclean = 0;
    if (makeclean) // Always send a WRITECLEAN
      do_writeclean = 1;
    else
      do_writeclean = $urandom_range(0,2);
    if (do_writeclean == 1) begin
      send_writeclean_xact(target_port_id,addr);
    end
  endtask

  /** sends a writeclean transaction on the specified port with the specified address */
  task send_writeclean_xact(int target_port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    `svt_xvm_create_on(basic_writeclean, p_sequencer.master_sequencer[target_port_id])
    basic_writeclean.writeclean_wt = 1;
    basic_writeclean.directed_addr_mailbox.put(addr);
    void'(basic_writeclean.randomize with {use_directed_addr == 1;sequence_length==1;});
    basic_writeclean.start(p_sequencer.master_sequencer[target_port_id]);
    basic_writeclean.wait_for_active_xacts_to_end();
  endtask

  /** Sends READSHARED transaction from all ACE ports in the system other than target_port_id */
  task send_readshared_xact(int target_port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, output int last_readshared_port);
    foreach(p_sequencer.master_sequencer[i]) begin
      if (
           (i != target_port_id) && 
           (cfg.master_cfg[i].is_active) && 
           cfg.is_participating(i) &&
           (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
         ) begin
        bit is_device_dvm_ok_for_interleaving;
        if (cfg.is_address_in_range_for_port_interleaving(addr,cfg.master_cfg[i],0,0,0,is_device_dvm_ok_for_interleaving) == 1)begin
          last_readshared_port = i;
          begin
            `svt_xvm_create_on(basic_readshared, p_sequencer.master_sequencer[i])
             basic_readshared.readshared_wt = 1;
             basic_readshared.directed_addr_mailbox.put(addr);
             void'(basic_readshared.randomize with {use_directed_addr == 1;sequence_length==1;});
             basic_readshared.start(p_sequencer.master_sequencer[i]);
          end 
          // Wait for ReadShared transactions to finish
          basic_readshared.wait_for_active_xacts_to_end();
        end
      end
    end
  endtask

  // Invalidate some random cachelines on last_readshared_port.
  // The last master that issued READSHARED has more number of cachelines
  // allocated, so invalidate more lines from that master. This is becuase when
  // a master is snooped as a result of a READSHARED its cacheline may get invalidated
  // (because it is legal to invalidate one's cacheline when snooped by a REAADSHARED).
  // The randomization of "do_invalidate" takes this into account.
  task invalidate_rand_cachelines(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,int last_readshared_port);
    bit do_invalidate = 0;
    do_invalidate = $urandom_range(0,2);
    if (do_invalidate == 1) begin
      send_invalidate_xact(last_readshared_port,addr);
    end
  endtask

  /** Sends a sequence that invalidates a cache line on the specified port for the specified address */
  task send_invalidate_xact(int target_port_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    svt_axi_cacheline_invalidation   cacheline_invalidation;
    `svt_xvm_create(cacheline_invalidation)
    cacheline_invalidation.invalidate_port = target_port_id;
    cacheline_invalidation.invalidate_addr = addr;
    cacheline_invalidation.start(p_sequencer);
  endtask

endclass: svt_axi_cacheline_initialization 

// =============================================================================
/** 
 * This sequence invalidates the cache line of a master.
 * It checks the state of the cache line and initiaties the appropriate transaction
 * If the cacheline state is dirty, a WRITEBACK is initiated.
 * If the cacheline state is clean, an EVICT is initiated.
 */
class svt_axi_cacheline_invalidation extends svt_axi_ace_master_base_virtual_sequence;

  /**  If use_directed_addr is set, this variable decides the addr to be invalidated */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0]  invalidate_addr;

  /*
   * The port on which invalidate operation needs to be done.
   */
  int invalidate_port = 0;

  svt_axi_basic_writeback_full_cacheline           basic_writeback;
  svt_axi_ace_master_base_sequence                 basic_evict;

  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] aligned_addr;
  bit curr_status = 0;
  bit temp_is_unique, temp_is_clean;


  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_cacheline_invalidation)

  function new(string name = "svt_axi_cacheline_invalidation");
    super.new(name);
  endfunction


  virtual task body();
    svt_axi_master_agent              my_agent;
    `SVT_XVM(component)                     my_component;
    svt_axi_cache                     my_cache;
    int                               target_port;
    // Populates master_xacts from parent
    super.body();
    target_port = invalidate_port;
    my_component = p_sequencer.master_sequencer[target_port].get_parent();      
    $cast(my_agent,my_component);
    my_cache = my_agent.get_cache();

    if (my_cache != null) begin
      bit is_unique, is_clean, cache_status;
      cache_status = my_cache.get_status(get_tagged_addr(invalidate_addr, target_port),is_unique,is_clean);
      if (cache_status && is_clean)
        begin
        initiate_basic_evict(target_port,invalidate_addr);
        end
      else if(cache_status && !is_clean) 
        begin
        initiate_basic_writeback(target_port,invalidate_addr);
        end

    end
    if (basic_evict != null)
      basic_evict.wait_for_active_xacts_to_end();
    if (basic_writeback != null)
      basic_writeback.wait_for_active_xacts_to_end();
  endtask: body

  /** Initiates an evict transaction for the specified port and address */
  task initiate_basic_evict(int target_port, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    `svt_xvm_create_on(basic_evict, p_sequencer.master_sequencer[target_port])
    basic_evict.evict_wt = 1;
    basic_evict.directed_addr_mailbox.put(addr);
    void'(basic_evict.randomize with {use_directed_addr == 1;sequence_length==1;});
    basic_evict.start(p_sequencer.master_sequencer[target_port]);
  endtask

  /** Initiates a writeback transaction for the specified port and address */
  task initiate_basic_writeback(int target_port, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
    `svt_xvm_create_on(basic_writeback, p_sequencer.master_sequencer[target_port])
    basic_writeback.directed_addr_mailbox.put(addr);
    void'(basic_writeback.randomize with {use_directed_addr == 1;sequence_length==1;});
    basic_writeback.start(p_sequencer.master_sequencer[target_port]);
  endtask

endclass: svt_axi_cacheline_invalidation
// =============================================================================

// =============================================================================
/**
 * This sequence generates a writeback transaction for a full cacheline.
 */
class svt_axi_basic_writeback_full_cacheline extends svt_axi_ace_master_base_sequence;
  
  `svt_xvm_declare_p_sequencer(svt_axi_master_sequencer)

  `svt_xvm_object_utils(svt_axi_basic_writeback_full_cacheline)

  function new(string name="svt_axi_basic_writeback_full_cacheline");
    super.new(name);
    writeback_wt = 1;
  endfunction

  virtual task pre_master_base_seq_item_randomize(bit is_valid_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] my_addr, output svt_axi_master_transaction master_xact);
    svt_axi_port_configuration port_cfg;
    svt_configuration get_cfg;
    int this_burst_size, this_burst_length;
    int log_base_2_data_width_in_bytes;
    int log_base_2_cache_line_size;
    p_sequencer.get_cfg(get_cfg);
    if (!$cast(port_cfg, get_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_port_configuration class");
    end
    `protected
WM9WCQ2_H[cI#e\WJ-ACe/I>/W7KZ4fG8.[Z(&Z:dcBPfNYZMe#9/)B/G4FHaNN&
[.f_YFBH<HX7>+Aab\ecXaS>6R<UQ,D8:M=bP4+:IHE@16L>-68E#6eET2c<Kbe7
G&TV.b&W<P=?bKS>0A80(>BJU]VILeKb?D4;1a35I.QVH5CLJ;E/c99JL1AJ&44F
3(;9Faa?/:B@E//5\1Nd]+Ye5_-FUZ5+7?53^FYEb9\F_2X^O+Q_H5I2]K9Q9[\X
4Ua2HY4QQ?,>SQ+d-e5=.<c[;ELcMG=W@K^WfI2CE96cI6VD87)e-W-7)0HWWB,.
e/ZFV5WF=U4ef6Z.WKRBVU>8DI[_UX?d_V)UN_E0W#](;D9b,V(>TUd99DK^TaIEQ$
`endprotected

    this_burst_length = port_cfg.cache_line_size/(port_cfg.data_width/8);
    `svt_xvm_create(master_xact)
    master_xact.port_cfg = port_cfg;
    if (is_valid_addr)
      my_addr = (my_addr >> log_base_2_data_width_in_bytes) << log_base_2_data_width_in_bytes;
    void'(master_xact.randomize() with { 
      xact_type == svt_axi_transaction::COHERENT;
      coherent_xact_type == svt_axi_transaction::WRITEBACK;
      if (!exclusive_access_enable)
        atomic_type == NORMAL;
      else
        atomic_type inside {NORMAL,EXCLUSIVE};
      if (is_valid_addr){
        if (burst_type == svt_axi_transaction::INCR)
          addr == ((my_addr >> local::log_base_2_cache_line_size) << local::log_base_2_cache_line_size);
        else
          addr == my_addr;
      }
      burst_length == this_burst_length;
      // burst_type == svt_axi_transaction::WRAP;
      burst_type inside {svt_axi_transaction::INCR,svt_axi_transaction::WRAP};
      burst_size == this_burst_size; 
      foreach (wstrb[i])
        wstrb[i] == (1<<(1<<this_burst_size)) - 1;
    });
    `svt_xvm_debug("pre_master_base_seq_item_randomize",$psprintf("is_valid_addr = 'b%0b. addr = 'h%0x. generated xact %0s",is_valid_addr,my_addr,`SVT_AXI_PRINT_PREFIX1(master_xact))) ;
  endtask
endclass: svt_axi_basic_writeback_full_cacheline 

// =============================================================================
/**
 * This sequence generates a writeclean transaction for a full cacheline.
 */
class svt_axi_basic_writeclean_full_cacheline extends svt_axi_ace_master_base_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_master_sequencer)

  `svt_xvm_object_utils(svt_axi_basic_writeclean_full_cacheline)

  function new(string name="svt_axi_basic_writeclean_full_cacheline");
    super.new(name);
    writeclean_wt = 1;
  endfunction

  virtual task pre_master_base_seq_item_randomize(bit is_valid_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] my_addr, output svt_axi_master_transaction master_xact);
    svt_axi_port_configuration port_cfg;
    svt_configuration get_cfg;
    int this_burst_size, this_burst_length;
    int log_base_2_data_width_in_bytes;
    int log_base_2_cache_line_size;
    p_sequencer.get_cfg(get_cfg);
    if (!$cast(port_cfg, get_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_port_configuration class");
    end
    this_burst_length = port_cfg.cache_line_size/(port_cfg.data_width/8);
    `protected
G<4[)QUGJ6C)<WQZ5)K(@;]NbEY)]Y6CP#Ba5AgG=B3JI6J2E2?e2)/L#P00.PBd
Wbe1@0VC-+HQ2(;JfF/c.BH6#[(3VaDd(5;=J6aR=6YJ6ba7,O#2_NEU#=BfN--;
QJA_XbfTPP,JG9<APG(A78GcfDXd#_1D)65_7AA0W#0-eZRM4W?EFGEXK8b26S[1
Hg=INM\,REZA5f^DNda9)#\C]RIFAHJMLQIF&;@PM>.;L1PC:.(BOQQ<GKXJ88Nc
VH=)<4#\JNIL#?C,EOSC(OP?&NOF>[A-T)D6IfQ]4VRE,[\+^4(+b5>6M-?=MRUV
Cc]=K8XKP5@HNCVYN/]81/F2S&EE4gFbTB1cOU644.]+I;BWP(OXRI>6P$
`endprotected

    `svt_xvm_create(master_xact)
    master_xact.port_cfg = port_cfg;
    if (is_valid_addr)
      my_addr = (my_addr >> log_base_2_data_width_in_bytes) << log_base_2_data_width_in_bytes;
    void'(master_xact.randomize() with { 
      xact_type == svt_axi_transaction::COHERENT;
      coherent_xact_type == svt_axi_transaction::WRITECLEAN;
      if (is_valid_addr){
        if (burst_type == svt_axi_transaction::INCR)
          addr == ((my_addr >> local::log_base_2_cache_line_size) << local::log_base_2_cache_line_size);
        else
          addr == my_addr;
      }      
      burst_length == this_burst_length;
      // burst_type == svt_axi_transaction::WRAP;
      burst_type inside {svt_axi_transaction::INCR,svt_axi_transaction::WRAP};
      if (!exclusive_access_enable)
        atomic_type == NORMAL;
      else
        atomic_type inside {NORMAL,EXCLUSIVE};
      burst_size == this_burst_size; 
      foreach (wstrb[i])
        wstrb[i] == (1<<(1<<this_burst_size)) - 1;
    });
  endtask
endclass: svt_axi_basic_writeclean_full_cacheline 
// ================================================================================

// ----------------------------------------------------------------------------
// BASE CLASSES USED FOR DVM SEQUENCES
/** This sequence generates dvm transactions with all possible dvm message types
 * from ACE or ACE-Lite+DVM master ports. This sequence is used as a base
 * sequence for higher level sequences, with proper constraints for sequence
 * members dvm_message_type and seq_xact_type */
class svt_axi_ace_master_dvm_base_sequence extends svt_axi_master_base_sequence;

   //* local field used to set relevant transaction item fields */
   rand svt_axi_transaction::coherent_xact_type_enum seq_xact_type;  
   rand bit [2:0] dvm_message_type = 3'b000;
   

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_object_utils_begin(svt_axi_ace_master_dvm_base_sequence)
    `uvm_field_int      (dvm_message_type,UVM_ALL_ON)
    `uvm_field_enum     (svt_axi_transaction::coherent_xact_type_enum,   seq_xact_type, UVM_ALL_ON)
  `uvm_object_utils_end
`elsif SVT_OVM_TECHNOLOGY
  `ovm_object_utils_begin(svt_axi_ace_master_dvm_base_sequence)
    `ovm_field_int      (dvm_message_type,OVM_ALL_ON)
    `ovm_field_enum     (svt_axi_transaction::coherent_xact_type_enum,   seq_xact_type, OVM_ALL_ON)
  `ovm_object_utils_end
`endif

`ifdef SVT_MULTI_SIM_ENUM_SCOPE
  // Property needed because MTI 10.0a can't seem to find enums defined in a class
  // scope unless that class is declared somewhere in that file or an included file.
  svt_axi_transaction base_xact;
`endif

  function new(string name="svt_axi_ace_master_dvm_base_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    super.pre_body();
  endtask: pre_body

  virtual task body();
    int unsigned sequence_length = 1;

    super.body();


    /* randomize the item and 
       set the addr and coherent_xact_type from local fields */
    
    `svt_xvm_do_with(req, 
      { 
        req.addr[14:12] == dvm_message_type;
        req.data_before_addr == 0;
        req.xact_type == svt_axi_transaction::COHERENT;
        req.burst_type != svt_axi_transaction::FIXED;
        req.coherent_xact_type == seq_xact_type;
      })
    `svt_xvm_debug("body",$psprintf("Sending DVM transaction %0s on port 'd%0d. dvm_message_type = 'h%0x",`SVT_AXI_PRINT_PREFIX1(req),req.port_cfg.port_id,dvm_message_type));
      /* 
      Please refer class reference manual on details of following fields
      svt_axi_transaction::is_coherent_xact_dropped
      svt_axi_transaction::is_cached_data
      */
      if(!req.is_coherent_xact_dropped && !req.is_cached_data) begin
         //get_response(rsp);
         wait (`SVT_AXI_XACT_STATUS_ENDED(req));
      end
    `svt_xvm_debug("body",$psprintf("Got response for DVM transaction %0s",`SVT_AXI_PRINT_PREFIX1(req)));

  endtask: body
endclass: svt_axi_ace_master_dvm_base_sequence
          

/** This sequence sends DVM Complete transactions from ACE or ACE-Lite+DVM Master
 * ports. It takes care of the ACE protocol requirement that DVM Sync handshake
 * on the snoop address channel be observed before issuing DVM Complete transaction. */
class svt_axi_ace_master_dvm_complete_sequence extends svt_axi_master_base_sequence;

  /** 
    * The snoop response sequence running on this port. Must be assigned by 
    * the sequence calling this sequence
    */
  svt_axi_ace_master_snoop_response_sequence snoop_resp_seq;

`ifdef SVT_UVM_TECHNOLOGY
  uvm_phase parent_starting_phase;
`elsif SVT_OVM_TECHNOLOGY
  ovm_phase parent_starting_phase;
`endif

  /** UVM Object Utility macro */
`ifdef SVT_UVM_TECHNOLOGY
  `uvm_object_utils(svt_axi_ace_master_dvm_complete_sequence)
`elsif SVT_OVM_TECHNOLOGY
  `ovm_object_utils(svt_axi_ace_master_dvm_complete_sequence)
`endif

  /** Class Constructor */
  function new (string name = "svt_axi_ace_master_dvm_complete_sequence");
    super.new(name);
  endfunction : new

  /** Raise an objection if this is the parent sequence */
  virtual task pre_body();
    super.pre_body();
  endtask: pre_body

  /** Drop an objection if this is the parent sequence */
  virtual task post_body();
    super.post_body();
  endtask: post_body
  
  virtual task body();
    bit status;
`ifdef SVT_UVM_TECHNOLOGY
    uvm_component my_component;
`elsif SVT_OVM_TECHNOLOGY
    ovm_component my_component;
`endif
    svt_configuration base_cfg;
    svt_axi_port_configuration port_cfg;

    `svt_xvm_debug("body", "Entered...");
    p_sequencer.get_cfg(base_cfg);
    if (!$cast(port_cfg, base_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_system_configuration class");
    end
    my_component = p_sequencer.get_parent();
    if (snoop_resp_seq == null) begin
     `svt_xvm_fatal("body","The snoop_resp_seq member of this class must be set by the sequence calling this sequence")
    end

    fork
    // Wait on DVM Sync and send DVM Complete
    begin
      `SVT_DATA_BASE_OBJECT_TYPE ev_xact;
      svt_axi_snoop_transaction snoop_xact;
      svt_axi_ace_master_dvm_base_sequence dvm_complete_seq= new("dvm_complete_seq");
      while (1) begin
        `svt_xvm_debug("body",$psprintf("Waiting for DVM SYNC on master 'd%0d with snoop_resp_Seq='d%0d",port_cfg.port_id, snoop_resp_seq));
        `protected
/bQAL?PW=/@=GI#<^(:8a[cS<0Y,J+P3JO8:SV_SbR5977&G@d:M,)CLSbB]@35X
N]#7;D8D?_J2[d^K9>acY,[I-VHCc>LdG7:PS+V5PZF.<8B+<Y-FVQ.8/?9=V@;.
4]B\W;./?gDN@c1K/Yb#,K@C:[YM],=?)IJQ.0Z-dY[.H$
`endprotected

        if (!$cast(snoop_xact,ev_xact)) begin
          `svt_xvm_fatal("body","Transaction obtained through EVENT_DVM_SYNC_XACT is not of type svt_axi_snoop_transaction");
        end
        `svt_xvm_debug("body",$psprintf("DVM SYNC received on master 'd%0d",snoop_xact.port_cfg.port_id));
        if (snoop_xact.port_cfg.port_id == port_cfg.port_id) begin
          fork
          begin
`ifdef SVT_UVM_TECHNOLOGY
            raise_phase_objection();
`endif
            `svt_xvm_debug("body",$psprintf("Received DVM SYNC on port 'd%0d, waiting for transaction to end",port_cfg.port_id));
            wait(snoop_xact.snoop_resp_status == svt_axi_snoop_transaction::ACCEPT);
            `svt_xvm_debug("body",$psprintf("DVM SYNC on port 'd%0d completed, initiating DVM complete",port_cfg.port_id));
            `svt_xvm_do_with(dvm_complete_seq,
                         {seq_xact_type==svt_axi_transaction::DVMCOMPLETE;
                          dvm_message_type == 3'b000;}
                    ) 
            `svt_xvm_debug("body",$psprintf("DVM COMPLETE on port 'd%0d completed",port_cfg.port_id));
`ifdef SVT_UVM_TECHNOLOGY
            drop_phase_objection();
`endif
          end
          join_none
        end
      end
    end
    join_none
    `svt_xvm_debug("body", "Exiting...");
  endtask: body
endclass: svt_axi_ace_master_dvm_complete_sequence

// END OF BASE CLASSES USED FOR DVM SEQUENCES
// ----------------------------------------------------------------------------

//------------------------------------------------------------------------------------
// BASE CLASSES USED FOR BARRIER SEQUENCES
/**
  * Sends a single WRITEUNIQUE transaction that writes into a location within the
  * given domain type. The transaction addresses a single byte and is meant as a flag
  * which can later be read by other transactions. Typically this is used as a post barrier
  * transaction to signal availability/observability of a number of pre barrier transactions
  */
class svt_axi_ace_barrier_flag_write_xact_sequence extends svt_axi_ace_master_base_sequence;

  rand svt_axi_transaction::xact_shareability_domain_enum flag_domain_type;

  /** Indicates if this transaction is to write into a single byte (meant as a flag) */
  bit is_single_byte_flag_xact = 1;

  /** The write barrier transaction to which this post-barrier transaction is to be associated */
  svt_axi_master_transaction assoc_write_barrier_xact;

  /** The read barrier transaction to which this post-barrier transaction is to be associated */
  svt_axi_master_transaction assoc_read_barrier_xact;

  svt_axi_master_transaction output_xact;

  `svt_xvm_object_utils(svt_axi_ace_barrier_flag_write_xact_sequence)

  function new(string name = "svt_axi_ace_barrier_flag_write_xact_sequence");
    super.new(name);
    // Dummy setting so that base class does not complain. Not used.
    writeunique_wt = 1;
  endfunction  

  virtual task body();
    bit rand_success = 0;
    int my_log_base_2_data_width_in_bytes;
    svt_axi_master_transaction flag_xact;
    // Before we start, create the transaction which will write into a flag location, because the second
    // master needs to continuosly read from that location
    flag_xact = svt_axi_master_transaction::type_id::create("flag write xact"); 
    `svt_xvm_create(flag_xact);
    flag_xact.port_cfg = port_cfg;
    `protected
g>9HPf(R=.7?#<S7B(>:EJTL5UfFf?MaCcG:EXQH(GH>Z4JX)BaT6)V_CTV4@e7#
/f=U2c2C1A^>X-1_U?dU>KIUV?U\<\(D;08#8d+40+Xf^#]^+E5O4Xef7D>-(?=.
4AXP?c&.DZ&Ye;PDNd@G#DJ/MZM_/ZYK:IJP\B,X.G:V+MW<)YR]fFUe_&Xd;5ZeQ$
`endprotected

    if (is_single_byte_flag_xact) begin
      rand_success = flag_xact.randomize() with {
                       // Align to data_width
                       addr == (addr >> my_log_base_2_data_width_in_bytes) << my_log_base_2_data_width_in_bytes;
                       domain_type == flag_domain_type;
                       xact_type == svt_axi_transaction::COHERENT;
                       coherent_xact_type == svt_axi_transaction::WRITEUNIQUE;
                       burst_length == 1;
                       atomic_type == svt_axi_transaction::NORMAL;
                       foreach (wstrb[i])
                         wstrb[i] == 1'b1;
                       burst_size == svt_axi_transaction::BURST_SIZE_8BIT;
                       associate_barrier == 1;
                     }; 
    end
    else begin
      rand_success = flag_xact.randomize() with {
                       domain_type == flag_domain_type;
                       xact_type == svt_axi_transaction::COHERENT;
                       atomic_type == svt_axi_transaction::NORMAL;
                       coherent_xact_type inside {svt_axi_transaction::WRITEUNIQUE,svt_axi_transaction::READONCE,
                                                  svt_axi_transaction::WRITENOSNOOP,svt_axi_transaction::READNOSNOOP};
                       associate_barrier == 1;
                     }; 
    end
    if (!rand_success) begin
      // Error
    end
    else begin
      flag_xact.associated_barrier_xact = svt_axi_barrier_pair_transaction::type_id::create("flag_xact.associate_barrier_xact"); 
      flag_xact.associated_barrier_xact.is_paired = 1;
      flag_xact.associated_barrier_xact.write_barrier = assoc_write_barrier_xact;
      flag_xact.associated_barrier_xact.read_barrier = assoc_read_barrier_xact;
      `svt_xvm_send(flag_xact);
      output_xact = flag_xact;
    end
  endtask
endclass

/**
  * Sends a single READONCE transaction that writes into a location within the
  * given domain type and address. The transaction addresses a single byte and is meant as one 
  * which reads a flag set by another transaction. Typically this is used to read a flag 
  * set through a post barrier transaction sent from another port.
  */
class svt_axi_ace_barrier_flag_read_xact_sequence extends svt_axi_ace_master_base_sequence;

  rand svt_axi_transaction::xact_shareability_domain_enum flag_domain_type;

  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] flag_addr;

  svt_axi_master_transaction output_read_xact;

  `svt_xvm_object_utils(svt_axi_ace_barrier_flag_read_xact_sequence)

  function new(string name = "svt_axi_ace_barrier_flag_read_xact_sequence");
    super.new(name);
    // Dummy setting so that base class does not complain. Not used.
    readonce_wt = 1;
  endfunction  

  virtual task body();
    bit rand_success = 0;
    svt_axi_master_transaction flag_read_xact;
    // Before we start, create the transaction which will write into a flag location, because the second
    // master needs to continuosly read from that location
    flag_read_xact = svt_axi_master_transaction::type_id::create("flag read xact"); 
    `svt_xvm_create(flag_read_xact);
    flag_read_xact.port_cfg = port_cfg;
    rand_success = flag_read_xact.randomize() with {
                     domain_type == flag_domain_type;
                     xact_type == svt_axi_transaction::COHERENT;
                     coherent_xact_type == svt_axi_transaction::READONCE;
                     burst_length == 1;
                     atomic_type == svt_axi_transaction::NORMAL;
                     burst_size == svt_axi_transaction::BURST_SIZE_8BIT;
                     addr == flag_addr;
                   }; 
    if (!rand_success) begin
      // Error
    end
    else begin
      `svt_xvm_send(flag_read_xact);
      output_read_xact = flag_read_xact;
    end
  endtask
endclass

//#######################################################################
//BARRIER_MEM PAIR 
//#######################################################################
/**
  * Sends a barrier pair
  */
class svt_axi_ace_barrier_pair_sequence extends svt_axi_ace_master_base_sequence;


  // Barrier ID as randomized by this sequence
  // This is an output after randomization of barrier transaction. 
  int  barrier_id;
 
  svt_axi_master_transaction            write_barrier_xact;
  svt_axi_master_transaction            read_barrier_xact;

  rand svt_axi_transaction::xact_shareability_domain_enum
            myDomain =svt_axi_transaction::INNERSHAREABLE;

  `svt_xvm_object_utils(svt_axi_ace_barrier_pair_sequence)

  //*************************************************************************
  /** Class Constructor */
  //*************************************************************************
  function new(string name="svt_axi_ace_barrier_pair_sequence");
    super.new(name);
    // Dummy setting so that base class does not complain. Not used.
    makeunique_wt = 1;
  endfunction
  
  //*************************************************************************
  // Body
  //*************************************************************************
  virtual task body();

    //=====================================================
    /** Set up the transaction */
    //=====================================================

    `svt_xvm_create(write_barrier_xact)
    void'(write_barrier_xact.randomize() with {
          xact_type == svt_axi_transaction::COHERENT;
          coherent_xact_type == svt_axi_transaction::WRITEBARRIER;
          barrier_type ==svt_axi_transaction::MEMORY_BARRIER;
          addr == 'h0;
          domain_type == myDomain;
          burst_length == 1;
          associate_barrier==0;
          prot_type == svt_axi_transaction::DATA_SECURE_NORMAL;
          data_before_addr == 0;    
          atomic_type == svt_axi_transaction::NORMAL;
          foreach(data[i]) data[i]==0;
          foreach(cache_write_data[i]) cache_write_data[i]==0;
  });
    //=====================================================
    //send to VIP
    //=====================================================
    //send trans to VIP
    `svt_xvm_send(write_barrier_xact)
    `svt_xvm_create(read_barrier_xact)
    void'(read_barrier_xact.randomize() with {
          xact_type == svt_axi_transaction::COHERENT;
          coherent_xact_type == svt_axi_transaction::READBARRIER;
          barrier_type ==svt_axi_transaction::MEMORY_BARRIER;
          addr == 'h0;
          domain_type == myDomain;
          burst_length == 1;
          id == write_barrier_xact.id;
          associate_barrier==0;
          prot_type == svt_axi_transaction::DATA_SECURE_NORMAL;
          data_before_addr == 0;
          atomic_type == svt_axi_transaction::NORMAL;
          foreach(data[i]) data[i]==0;
          foreach(cache_write_data[i]) cache_write_data[i]==0;
  });
    //=====================================================
    //send to VIP
    //=====================================================
    //send trans to VIP
    `svt_xvm_send(read_barrier_xact)
  endtask: body

endclass: svt_axi_ace_barrier_pair_sequence

/**
  * Sends a single READNOSNOOP transaction that reads from the same location 
  * as write_xact. Associates the READ to a barrier based on associate_barrier
  */
class svt_axi_ace_barrier_readnosnoop_sequence extends svt_axi_ace_master_base_sequence;

  /** Indicates if this transaction must be associated with a barrier */
  bit my_associate_barrier = 0;

  /** The write transaction to which address this read must be sent */
  svt_axi_master_transaction write_xact;

  /** The read barrier transaction to which this post-barrier transaction is to be associated */
  svt_axi_master_transaction assoc_read_barrier_xact;

  /** The write barrier transaction to which this post-barrier transaction is to be associated */
  svt_axi_master_transaction assoc_write_barrier_xact;

  svt_axi_master_transaction output_read_xact;

  `svt_xvm_object_utils(svt_axi_ace_barrier_readnosnoop_sequence)

  function new(string name = "svt_axi_ace_barrier_readnosnoop_sequence");
    super.new(name);
    // Dummy setting so that base class does not complain. Not used.
    readnosnoop_wt = 1;
  endfunction  

  virtual task body();
    bit rand_success = 0;
    int my_log_base_2_data_width_in_bytes;
    svt_axi_master_transaction readnosnoop_xact;
    // Before we start, create the transaction which will write into a flag location, because the second
    // master needs to continuosly read from that location
    readnosnoop_xact = svt_axi_master_transaction::type_id::create("flag write xact"); 
    `svt_xvm_create(readnosnoop_xact);
    readnosnoop_xact.port_cfg = port_cfg;
    rand_success = readnosnoop_xact.randomize() with {
          xact_type == svt_axi_transaction::COHERENT;
          coherent_xact_type == svt_axi_transaction::READNOSNOOP;
          addr == write_xact.addr;
          burst_size == write_xact.burst_size;
          burst_type == write_xact.burst_type;
          burst_length == write_xact.burst_length;
          associate_barrier == my_associate_barrier;
          atomic_type == svt_axi_transaction::NORMAL;
        };
    if (my_associate_barrier) begin
      readnosnoop_xact.associated_barrier_xact = svt_axi_barrier_pair_transaction::type_id::create("readnosnoop_xact.associate_barrier_xact"); 
      readnosnoop_xact.associated_barrier_xact.is_paired = 1;
      readnosnoop_xact.associated_barrier_xact.write_barrier = assoc_write_barrier_xact;
      readnosnoop_xact.associated_barrier_xact.read_barrier = assoc_read_barrier_xact;
    end
    `svt_xvm_debug("body",$sformatf("Sending post barrier read transaction %0s",`SVT_AXI_PRINT_PREFIX1(readnosnoop_xact)));
    `svt_xvm_send(readnosnoop_xact);
    output_read_xact = readnosnoop_xact;
  endtask

endclass
// END OF BASE CLASSES USED FOR BARRIER SEQUENCES
//--------------------------------------------------------------------


//####################################################################
// ACE Exclusive sequence
//####################################################################

 /**     
   * This sequence is used to create Exclusive Access Transactions at Master port level<br>
   *<br>
   * Transaction Sequences Used: Exclusive Load followed by Exclusive store 
   * - Initialize cache lines if initialize_cachelines bit is set 
   * - Issue READCLEAN or READSHARED to load location and wait for the transaction to end
   * - Check the cache line state
   *   - if in Shared state issue CLEANUNIQUE 
   *   - if in Invalid state then restart Exclusive Access
   *   - else do nothing as Master can store directly to the cacheline no need to inform Interconnect
   *   .
   * - Stored data is updated to memory through WRITEBACK transaction
   * .
   * <br>
   * Please note, for generation of exclusive access transactions, svt_axi_port_configuration :: exclusive_access_enable 
   * should be set for the targeted master. <br>
   * <br> 
   */
 class svt_axi_ace_exclusive_access_sequence extends svt_axi_ace_master_base_sequence;
 
    rand bit [`SVT_AXI_MAX_BURST_LENGTH_WIDTH - 1 : 0]      exc_burst_length = 1;
    rand svt_axi_transaction::burst_size_enum               exc_burst_size   = svt_axi_transaction::BURST_SIZE_8BIT;
    rand svt_axi_transaction::burst_type_enum               exc_burst_type   = svt_axi_transaction::INCR;
    
    rand svt_axi_transaction::xact_shareability_domain_enum exc_domain = svt_axi_transaction::INNERSHAREABLE;
 
    svt_axi_master_transaction                              exclusive_load_xact;
    svt_axi_master_transaction                              exclusive_clean_xact;
    svt_axi_master_transaction                              write_xact;
    bit [1:0]                                               cache_line_state=0;
    bit                                                     exclusive_accesses_seq_successful = 0;
    rand int                                                exclusive_axi4_slave = 0;
    
    // Nummber of time time exlusive sequence will be restared if master exclusive monitor has been reset
    //or Store opreation recives OKAY response in stead of EXOKAY
    rand int                                                num_of_exclusive_seq_restart = 2;
    /** represents percentage value of sending random non-exclusive store overlapping with exclusive store.
      * Must set values between 0 to 100 
      */
    rand int                                                random_nonexclusive_store_overlap_with_exclusive_store_wt = 20;

    constraint random_nonexclusive_store_overlap_with_exclusive_store_wt_con {
        random_nonexclusive_store_overlap_with_exclusive_store_wt dist {0:=20, [1:50]:/50, [51:100]:/30};
    }
 
 `ifdef SVT_UVM_TECHNOLOGY
    `uvm_object_utils_begin(svt_axi_ace_exclusive_access_sequence)
       `uvm_field_int     (exc_burst_length, UVM_ALL_ON)
       `uvm_field_enum    (svt_axi_transaction::burst_size_enum, exc_burst_size, UVM_ALL_ON)
       `uvm_field_enum    (svt_axi_transaction::burst_type_enum, exc_burst_type, UVM_ALL_ON)
       `uvm_field_enum    (svt_axi_transaction::xact_shareability_domain_enum, exc_domain, UVM_ALL_ON)
       `uvm_field_int     (num_of_exclusive_seq_restart, UVM_ALL_ON)
    `uvm_object_utils_end
 `elsif SVT_OVM_TECHNOLOGY
    `ovm_object_utils_begin(svt_axi_ace_exclusive_access_sequence)
       `ovm_field_int     (exc_burst_length, OVM_ALL_ON)
       `ovm_field_enum    (svt_axi_transaction::burst_size_enum, exc_burst_size, OVM_ALL_ON)
       `ovm_field_enum    (svt_axi_transaction::burst_type_enum, exc_burst_type, OVM_ALL_ON)
       `ovm_field_enum    (svt_axi_transaction::xact_shareability_domain_enum, exc_domain, OVM_ALL_ON)
       `ovm_field_int     (num_of_exclusive_seq_restart, OVM_ALL_ON)
    `ovm_object_utils_end
 `endif

    constraint valid_burst_type { exc_burst_type !=  svt_axi_transaction::FIXED;}
 
    function new(string name="svt_axi_ace_exclusive_access_sequence");
       super.new(name);
       // Dummy setting so that base class does not complain. Not used.
       readclean_wt = 1;
       random_nonexclusive_store_overlap_with_exclusive_store_wt = 20;
    endfunction // new
 
    virtual task body();
      bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0]  directed_addr;
      bit sts, is_error,randomize_with_directed_addr;
      bit exc_load_rand_success,clean_unique_rand_success,write_back_rand_success;
      svt_axi_master_transaction tr;
      bit random_nonexclusive_store_overlap_with_exclusive_store;
      bit repeat_exclusive_store = 0;

      `ifdef SVT_UVM_TECHNOLOGY
          sts = uvm_config_db#(int)::get(null, get_full_name(), "random_nonexclusive_store_overlap_with_exclusive_store_wt", random_nonexclusive_store_overlap_with_exclusive_store_wt);
      `else
          sts = m_sequencer.get_config_int({get_type_name(), ".random_nonexclusive_store_overlap_with_exclusive_store_wt"}, random_nonexclusive_store_overlap_with_exclusive_store_wt);
      `endif
      if(random_nonexclusive_store_overlap_with_exclusive_store_wt > 100)
        `svt_xvm_fatal("body",$psprintf("random_nonexclusive_store_overlap_with_exclusive_store_wt must have value between 0 to 100, its current value is 'd%0d", random_nonexclusive_store_overlap_with_exclusive_store_wt));

      //port_cfg.exclusive_access_enable
      if((port_cfg.axi_interface_type == svt_axi_port_configuration::AXI_ACE) && 
         (port_cfg.exclusive_access_enable == 1) && (port_cfg.is_active == 1)  ) begin
      
        `svt_xvm_debug("body",$psprintf("svt_axi_ace_exclusive_access_sequence - sequence_length - 'd%d",sequence_length));
      
        for(int i =0; i < sequence_length; i++) begin
          exclusive_accesses_seq_successful = 0;
          `svt_xvm_debug("body",$psprintf("svt_axi_ace_exclusive_access_sequence Next iteration  - 'd%d",i));
          //get_cache_line_state(cache_line_state);
         
          //if(!repeat_exclusive_store || cache_line_state==2'b00) begin
             //Get directed address if set 
             if (use_directed_addr) begin : tag_use_directed_addr
               `svt_xvm_debug("generate_transactions",$psprintf("Getting directed address for sequence %0s",this.get_full_name()));
               get_directed_addr((i+1),is_error,randomize_with_directed_addr,directed_addr);
               if (is_error) break;
             end : tag_use_directed_addr

             `svt_xvm_create(exclusive_load_xact);
             randomize_xact_for_exclusive_load(exclusive_load_xact,
                   randomize_with_directed_addr,
                   directed_addr,
                   exc_load_rand_success);
          //end

          if(!exc_load_rand_success) begin
            `svt_xvm_fatal("generate_transactions","Randomization failure!!");
          end
          else begin
            `svt_xvm_debug("body",$psprintf("Exclusive load transaction %0s",`SVT_AXI_PRINT_PREFIX1(exclusive_load_xact)));
      
            // If initializing, first initialize and then send transactions
            if (initialize_cachelines && !repeat_exclusive_store) begin
               parent_sequence.cacheline_init_sema.get();
               `protected
bb1_@^3J6-Abd1eLIQE&dFCAdRI[^^(H)US6;#OEWX3#6Re.;+g]0)/^AFX:&H6U
@8ddSML1ZC5U4Q]#O8\g0CAeESdOeg9Pf+_cGYB>W9\&Z+)NH_eKa^_:)QB7.3a)
YB[B/J8Q)Jb[;2MO_@,@Ye@A9715)=(Ya1E:RE@fV^AKdfU2\BK\Ab_Re1CN+2b3
JZ@\#ZD?Ne>Z1OCdYT6<Y?@A4$
`endprotected

               @parent_sequence.ev_cacheline_init_done;
               parent_sequence.cacheline_init_sema.put();
               `svt_xvm_debug("body","Cache Line Initialization done");
            end
             
            //Try to finish exclusive access sequence for num_of_exclusive_seq_restart times
            //if the exclusive store fails
            for(int j=0; j < num_of_exclusive_seq_restart; j++) begin
               //Check the cache line status, to check if the cache line is in SHARED state
               get_cache_line_state(cache_line_state);
             
               if(!repeat_exclusive_store || cache_line_state==2'b00) begin
                 `svt_xvm_debug("body",$psprintf("Initiating Exclusive Access Sequence: Attempt 'd%d",(j+1)));
                 //Initiate exlusive load transaction
                 `svt_xvm_send(exclusive_load_xact);
                 //Wait for exclusive load to finish
                 `svt_xvm_debug("body","Waiting for Exclusive Access load");
                 wait (`SVT_AXI_XACT_STATUS_ENDED(exclusive_load_xact));
                 if(exclusive_load_xact.is_coherent_xact_dropped || exclusive_load_xact.is_cached_data) begin
                    `svt_xvm_error("body",$psprintf("%s Droped - due to is_coherent_xact_dropped - 'b%b or is_cached_data - 'b%b",
                    exclusive_load_xact.coherent_xact_type.name(),exclusive_load_xact.is_coherent_xact_dropped,
                    exclusive_load_xact.is_cached_data));
                 end
                 
                 `svt_xvm_debug("body",$psprintf("Exclusive load transaction over %0s",`SVT_AXI_PRINT_PREFIX1(exclusive_load_xact)));
                 //If exclusive load recives OKAY response abort the exclusive access sequence, as 
                 //slave does not support Exclusive accesses
                 if (exclusive_load_xact.rresp[0] == svt_axi_transaction::OKAY && exclusive_load_xact.port_cfg.exclusive_monitor_enable) begin
                   `svt_xvm_warning("body",$psprintf("Exclusive Accesses not suppote by slave correspond to address - 'h%h. Aborting svt_axi_ace_exclusive_access_sequence", exclusive_load_xact.addr));
                   break;
                 end
               end
          
               //Add login for programmable wait
          
               //Check the cache line status, to check if the cache line is in SHARED state
               get_cache_line_state(cache_line_state);
             
               //If the cache line is in SHARED state, make it unique 
               if(cache_line_state == 2'b01) begin
                 // Initiate CLEANUNIQUE
                 `svt_xvm_create(exclusive_clean_xact);
                 randomize_xact_for_clean_unique(exclusive_clean_xact, clean_unique_rand_success);
                 if(!clean_unique_rand_success) begin
                   `svt_xvm_fatal("body","Randomization failure!!");
                 end
                 else begin
                   //Initiate CLEANUNIQUE
                   `svt_xvm_send(exclusive_clean_xact);
                   `svt_amba_debug("body",$sformatf("sent exclusive store from shared state - %s",`SVT_AXI_PRINT_PREFIX1(exclusive_clean_xact)));
                   randcase
                     (    random_nonexclusive_store_overlap_with_exclusive_store_wt) : random_nonexclusive_store_overlap_with_exclusive_store = 1;
                     (100-random_nonexclusive_store_overlap_with_exclusive_store_wt) : random_nonexclusive_store_overlap_with_exclusive_store = 0;
                   endcase
    
                   fork
                     //Wait for CLEANUNIQUE to finish on bus
                     wait (`SVT_AXI_XACT_STATUS_ENDED(exclusive_clean_xact));
                     if(random_nonexclusive_store_overlap_with_exclusive_store) begin
                       `svt_xvm_create(tr);
                       //tr.disable_all_weights();
                       void'(tr.randomize() with {
                               addr == exclusive_clean_xact.addr;
                               xact_type == svt_axi_transaction::COHERENT;
                               coherent_xact_type == svt_axi_transaction::CLEANUNIQUE;
                               atomic_type == svt_axi_transaction::NORMAL;
                             });
                       wait(exclusive_clean_xact.addr_status != svt_axi_transaction::INITIAL);
                       `svt_xvm_send(tr);
                       wait (`SVT_AXI_XACT_STATUS_ENDED(tr));
                     end
                   join
                   if(!exclusive_clean_xact.is_coherent_xact_dropped ) begin
                 
                      if(exclusive_clean_xact.rresp[0] == svt_axi_transaction::OKAY) begin
                        `svt_xvm_warning("body",$psprintf("Exclusive Accesses sequeance failed, CleanUnique correspond to address - 'h%h, got OKAY response instead of EXOKAY. Restarting exclusive access sequence", exclusive_clean_xact.addr));
                        repeat_exclusive_store = 0;
                        break;
                      end else begin
                        randcase
                          30: repeat_exclusive_store = 1;
                          70: repeat_exclusive_store = 0;
                        endcase
                        `svt_amba_debug("body",$sformatf("completed exclusive store - %s  repeat_store='d%0d",`SVT_AXI_PRINT_PREFIX1(exclusive_clean_xact), repeat_exclusive_store));
                      end
                   end // is_coherent_dropped
                   else repeat_exclusive_store = 0;
                   `svt_xvm_debug("body",$psprintf("CLEANUNIQUE part of Exclusive Accesses sequence is over %0s",`SVT_AXI_PRINT_PREFIX1(exclusive_clean_xact)));
                 end // else: !if(!clean_unique_rand_success)
             
                 if(!exclusive_clean_xact.is_coherent_xact_dropped && repeat_exclusive_store == 0) begin
                   //At this point Status is UNIQUE or CleanUnique transaction is over, store the date to memory
                   `svt_xvm_debug ("body","Send WRITEBACK");
                   `svt_xvm_create(write_xact);
                   randomize_xact_write_back(write_xact,write_back_rand_success);
              
                   if(!write_back_rand_success) begin
                   `svt_xvm_fatal("body","Randomization failure!!");
                   end
                   else begin
                     //Initiate write back transaction
                     `svt_xvm_send(write_xact);
                
                     //Wait for WriteBack to finish
                     wait (`SVT_AXI_XACT_STATUS_ENDED(write_xact));
                     if(write_xact.is_coherent_xact_dropped || write_xact.is_cached_data) begin
                       `svt_xvm_debug("body",$psprintf("WRITEBACK dropped - due to is_coherent_xact_dropped - 'b%b or is_cached_data - 'b%b", write_xact.is_coherent_xact_dropped, write_xact.is_cached_data));
                     end
                   
                     `svt_xvm_debug("body",$psprintf("WRITEBACK part of Exclusive Accesses sequence is over %0s",`SVT_AXI_PRINT_PREFIX1(write_xact)));
                   
                     //Exclusive Access Sequence successful, bresk num_of_exclusive_seq_restart loop
                     exclusive_accesses_seq_successful = 1;
                     break;
                   end // else: !if(!write_back_rand_success)
                 end // if(!exclusive.... && repeat_exclu...)
               end // if (cache_line_state == 2'b01)
               //Cache line in INVALID state
               else if (cache_line_state == 2'b00) begin 
                 `svt_xvm_debug ("body","Cacheline status - INVALID, restart exclusive access sequence");
                 //Line has been invalidated, retry exclusive accesses sequence
                 repeat_exclusive_store = 0;
                 continue;
               end
               else break;
            end // for (int j=0; j < num_of_exclusive_seq_restart; j++)
          
            if(exclusive_accesses_seq_successful) begin 
              `svt_xvm_debug("body",$psprintf("svt_axi_ace_exclusive_access_sequence was successful for iteration number - 'd%d",i)); 
            end else begin
              `svt_xvm_debug("body",$psprintf("svt_axi_ace_exclusive_access_sequence was unsuccessful for iteration number - 'd%d",i)); 
            end 
          end // else: !if(!exc_load_rand_success)
        end // for (int i =0; i < sequence_length; i++)
      end else begin
        `svt_xvm_warning("body","Port is not of ACE type, or exclusive_access_enable is not set, or agent is not active is not set in port configuration");
      end // else: !if(port_cfg.axi_interface_type == svt_axi_port_configuration::AXI_ACE)
   endtask // body
   
   // Randomize load transaction for exclusive accesses sequence
   virtual task randomize_xact_for_exclusive_load(svt_axi_master_transaction master_xact,
                bit randomize_with_directed_addr, 
                bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] directed_addr,
                output bit req_success);
      int log_base_2_cache_line_size;
      // Get config from corresponding sequencer and assign it here.
      master_xact.port_cfg = port_cfg;
      master_xact.port_id  = port_cfg.port_id;
      `protected
AT?MLD&C;LU_@@:GV\&NA4PT@#QR4YKY?O&H/aIVdMNdG;Q#Na,96)L)Y>@,]dLT
><<;M5G6#M1L][^]5QL@Vf?H;:K22^O]XQJ;8RMEV-B/S\GC3M1=6YBeMQWS609X
Ca+8YeeM>I401e\C;S2NM2K;]-)NYgU-.eBMKfHE@NF3f)GHXN84f[66f<3W3K&WQ$
`endprotected

      if (exc_burst_type == svt_axi_transaction::INCR) begin
        directed_addr = ((directed_addr >> log_base_2_cache_line_size) << log_base_2_cache_line_size);
      end
      req_success = master_xact.randomize() with { 
                   atomic_type  == svt_axi_transaction::EXCLUSIVE;
                   burst_size   == exc_burst_size;
                   burst_type   == exc_burst_type;
                   burst_length == exc_burst_length;     
                   if(exclusive_axi4_slave)
                     cache_type == 2;

                   if(port_cfg.max_num_exclusive_access > 0)
                      id < port_cfg.max_num_exclusive_access ;
                   if (port_cfg.use_separate_rd_wr_chan_id_width){
                     if (port_cfg.read_chan_id_width < port_cfg.write_chan_id_width){
                       id <= ((1 << port_cfg.read_chan_id_width) - 1);
                     }else if (port_cfg.write_chan_id_width < port_cfg.read_chan_id_width) {
                       id <= ((1 << port_cfg.write_chan_id_width) - 1);
                     }
                   }
                   if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
                       xact_type == svt_axi_transaction::COHERENT;
                       coherent_xact_type inside {svt_axi_transaction::READCLEAN,svt_axi_transaction::READSHARED };     
                   }
    
                   if (randomize_with_directed_addr)
                     addr == directed_addr;
                   // Fixed is currently not supported by interconnect
                   burst_type != svt_axi_transaction::FIXED;
                   force_xact_to_cache_line_size == force_to_cache_line_size;
                };
   endtask // randomize_xact_for_exclusive_load

   // Randomize for CLEANUNIQUE
   virtual task randomize_xact_for_clean_unique (svt_axi_master_transaction master_xact,
           output bit req_success);
      master_xact.port_cfg = port_cfg;
      master_xact.port_id  = port_cfg.port_id;

      req_success = master_xact.randomize() with {
              atomic_type  == svt_axi_transaction::EXCLUSIVE;
              burst_size   == exclusive_load_xact.burst_size;
              burst_type   == exclusive_load_xact.burst_type;
              burst_length == exclusive_load_xact.burst_length;            
              addr         == exclusive_load_xact.addr;
              domain_type  == exclusive_load_xact.domain_type;
              prot_type    == exclusive_load_xact.prot_type;
              cache_type   == exclusive_load_xact.cache_type;
              id           == exclusive_load_xact.id; 

              if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
                                                      xact_type          == svt_axi_transaction::COHERENT;
                                                      coherent_xact_type == svt_axi_transaction::CLEANUNIQUE;}
                                                  force_xact_to_cache_line_size == force_to_cache_line_size;};
      
   endtask // randomize_xact_for_exclusive_load

   // Randomize for WRITEBACK
   virtual task randomize_xact_write_back(svt_axi_master_transaction master_xact,
           output bit req_success);
      master_xact.port_cfg = port_cfg;
      master_xact.port_id  = port_cfg.port_id;

      req_success = master_xact.randomize() with {
              atomic_type  == svt_axi_transaction::NORMAL;
              burst_size   == exclusive_load_xact.burst_size;
              burst_type   == exclusive_load_xact.burst_type;
              burst_length == exclusive_load_xact.burst_length;            
              addr         == exclusive_load_xact.addr;
              domain_type  == exclusive_load_xact.domain_type;
              prot_type    == exclusive_load_xact.prot_type;
              cache_type   == exclusive_load_xact.cache_type;
              id           == exclusive_load_xact.id;
              data.size()  == exclusive_load_xact.burst_length;
              foreach (data[i]) data[i] == i;

              foreach (wstrb[i]) wstrb[i] == (1<<(1<<exclusive_load_xact.burst_size)) - 1;
                if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
                                                      xact_type          == svt_axi_transaction::COHERENT;
                                                      coherent_xact_type == svt_axi_transaction::WRITEBACK;}
                                                  force_xact_to_cache_line_size == force_to_cache_line_size;};
   endtask // randomize_xact_write_back

   // Get the cache line state for the address
   // 00 - INVALID
   // 01 - SHARED
   // 10 - UNIQUE
   virtual task get_cache_line_state(output bit [1:0] line_state);
     svt_axi_master_agent              my_agent;
     `SVT_XVM(component)               my_component;
     svt_axi_cache                     my_cache;
     bit                               is_unique,is_clean;
     my_component = p_sequencer.get_parent();      
     if(!$cast(my_agent,my_component)) begin
       `svt_xvm_fatal("get_cache_line_state", "Unable to Cast my_component tp my_agent");
     end
     if (my_agent != null) begin
       my_cache = my_agent.get_cache();
   
       if(my_cache != null) begin
         if(my_cache.get_status(exclusive_load_xact.get_tagged_addr(),is_unique, is_clean)) begin
       
         if(is_unique) line_state = 2'b10; //CacheLine is in UNIQUE state
         else          line_state = 2'b01; //CacheLine is in SHARED state
         end
         else begin
           line_state = 2'b00;
         end
         `svt_xvm_debug("get_cache_line_state", $psprintf("line_state - 'b%b", line_state));
       end // if (my_cache != null)
       else begin `svt_xvm_fatal("get_cache_line_state", "my_cache is null"); end
     end // if (my_agent != null)
     else begin
       `svt_xvm_fatal("get_cache_line_state", "my_agent is null");
     end // else: !if(my_agent != null)
   endtask // get_cache_line_stats
 endclass // svt_axi_ace_exclusive_access_sequence
`endif // GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_BASE_SV
