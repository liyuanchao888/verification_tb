
`ifndef GUARD_SVT_AHB_SYSTEM_ENV_SV
`define GUARD_SVT_AHB_SYSTEM_ENV_SV

// =============================================================================
/** This class is the System ENV class which contains all of the elements of an
 * AHB System. The AHB System ENV encapsulates master agents, slave agents,
 * system sequencer, system monitor and the system configuration.
 * 
 * The number of master and slave agents is configured based on the system
 * configuration provided by the user. In the build phase, the System ENV
 * builds the master and slave agents. After the master & slave agents are
 * built, the System ENV configures them using the configuration information
 * available in the system configuration.
 */
class svt_ahb_system_env extends svt_env;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_if svt_ahb_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB System virtual interface */
  svt_ahb_vif vif;

  /* AHB Master components */
  svt_ahb_master_agent master[$];

  /* AHB Slave components */
  svt_ahb_slave_agent slave[$];

  /* AHB System sequencer is a virtual sequencer with references to each master
   * and slave sequencers in the system.
   */
  svt_ahb_system_sequencer sequencer;

  /** AHB System Level Monitor */
  svt_ahb_system_monitor system_monitor;
  
  /** AHB System Level Checker whose checks are called from system_monitor */
  svt_ahb_system_checker system_checker;

  /** AHB System Level Transaction Coverage Callback */
  svt_ahb_system_monitor_def_cov_callback sys_mon_trans_cov_cb;

  /** The AHB Bus component. 
   */
  svt_ahb_bus_env bus;

  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_system_configuration cfg_snapshot;

`ifdef SVT_UVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  uvm_tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor */ 
  uvm_tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`elsif SVT_OVM_TECHNOLOGY
  /** Fifo into which transactions from master to BUS are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_master_transaction)  ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled */ 
  tlm_fifo#(svt_ahb_transaction)  ahb_bus_to_slv_transaction_fifo;

  /** Fifo into which transactions from master to BUS are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_master_transaction)  amba_ahb_mstr_to_bus_transaction_fifo;

  /** Fifo into which transactions from BUS to slave are put when system checker is enabled 
    * Used by AMBA System Monitor 
    */ 
  tlm_fifo#(svt_ahb_transaction)  amba_ahb_bus_to_slv_transaction_fifo;
`endif


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
 /* External AHB Master components */
  local svt_ahb_master_agent external_ahb_master_agent[int];

  /* External AHB Slave components */
  local svt_ahb_slave_agent external_ahb_slave_agent[int];

  /* External AHB Master component Port Configuraiton */
  local svt_ahb_master_configuration external_master_agent_cfg[int];

  /* External AHB Slave component Port Configuraiton */
  local svt_ahb_slave_configuration external_slave_agent_cfg[int];

  /** Configuration object for this ENV. */
  local svt_ahb_system_configuration cfg;

  /** Address mapper for the AHB system */
  local svt_mem_address_mapper mem_addr_mapper;

  /** MEM System Backdoor class which provides a system level view of the memory map */
  local svt_ahb_mem_system_backdoor mem_system_backdoor;

  /** MEM System Backdoor class which provides the global view of the memory map */
  local svt_ahb_mem_system_backdoor global_mem_system_backdoor;

/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_ahb_system_env)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new ENV instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name = "svt_ahb_system_env", `SVT_XVM(component) parent = null);

  /** Obtains the System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_mem_system_backdoor();

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the sub-agent components.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  /**
  * Report Phase
  * Reports performance statistics
  */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void report_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void report();
`endif


  // ---------------------------------------------------------------------------
  /**
   * Connect Phase:
   * Connects the virtual sequencer to the sub-sequencers
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * End of elaboration Phase
   * Displays the environment configuration.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void end_of_elaboration();
`endif  
  
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the ENV configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

/** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /**
   * Obtain the address mapper for the AHB System
   */
  extern function svt_mem_address_mapper get_mem_address_mapper();

  /** Obtains the Global System Memory Manager system backdoor class for this AHB system */
  extern function svt_ahb_mem_system_backdoor get_global_mem_system_backdoor();
/** @endcond */

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external master
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external master agent handle and its corresponding master index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * master agent.
    * 
    * If system env doesn't find any external master agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of master agents considering external
    * master agents and set specific master index for which external agent needs
    * to be used. It is allowed to instantiate some master agents within the
    * svt_ahb_system_env, and some master agents externally. User needs to take
    * care of correctly specifying the indices of external master agents to this
    * method.
    *
    * @param index Index of the master agent which is external to the AHB System Env
    *
    * @param mstr Handle of the master agent which is external to the AHB System Env
    *
    * @param mstr_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_master_agent(i,ahb_master_agent[i]);
    *
    */
  extern function void set_external_master_agent(int index, svt_ahb_master_agent mstr, svt_ahb_master_configuration mstr_cfg=null);

  /**
    * Enables AHB System Env class svt_ahb_system_env to use external slave
    * agent which is already created outside svt_ahb_system_env.  User needs to
    * provide external slave agent handle and its corresponding slave index
    * number. It is important that user creates System Configuration including
    * the port configuration which is supposed to be used by the external
    * slave agent.
    * 
    * If system env doesn't find any external slave agent for a specific index
    * then it creates one on its own. So, it is important for user to set system
    * configuration with correct number of slave agents considering external
    * slave agents and set specific slave index for which external agent needs
    * to be used. It is allowed to instantiate some slave agents within the
    * svt_ahb_system_env, and some slave agents externally. User needs to take
    * care of correctly specifying the indices of external slave agents to this
    * method.
    *
    * @param index Index of the slave agent which is external to the AHB System Env
    *
    * @param slv Handle of the slave agent which is external to the AHB System Env
    *
    * @param slv_cfg This parameter is not yet supported.
    *
    * Example:  for(int i=0; i<5; i++) ahb_system_env.set_external_slave_agent(i,ahb_slave_agent[i]);
    */
  extern function void set_external_slave_agent(int index, svt_ahb_slave_agent slv, svt_ahb_slave_configuration slv_cfg=null);

  /** @cond PRIVATE */
  extern function void set_external_master_agent_array(svt_ahb_master_agent mstr[int], svt_ahb_master_configuration mstr_cfg[int]);
  extern function void set_external_slave_agent_array(svt_ahb_slave_agent slv[int], svt_ahb_slave_configuration slv_cfg[int]);
  /** @endcond */

endclass

`protected
5DR2Eeg.=Wb]RBL1f7G2@f1H9;&WW57ULGA66&32195YE/\[UZ\..)(FA[7e#d4.
f8P(GL_R4ESYb6&&@,;B42?7.H(Hg_(e]CMfVb?_?5:4=+VGKF:BC]7\\M=8?U7g
[W6]Zd3e.()^O-^@/HaPfKTX@(IRD&.,XMQ-eX#H//0Vddg3:N\[C,PRN[SG=&bF
WDgcC4#LCGbRb:[>dT1)KCc[/_LLN[LNP^)EX_eN4[C5;<;g--BI?^(G?SeD7-6N
U8bX0g<[_\:^GS10ggJ&ZC30:BA?++V=.3&Tg,<GEaNS)(/1YOb26U6-D6OQf]7I
U8?(@Ke?+0d^/$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
g@acM8VS.aHV+-4aI6D5a]\#0YRFSS=E;10SA.+#;4bTK/_1NXgY1(J@C8X[HDNP
VBOPG7NTVG)Y?IJ6+LRG0_9g>/eT&O;VOV,UW@)c25FU31&\=/WcV3OC5]49-d#<
;1ed7,OZ:OE+Ng-=;W)6TS>A1M2]P8KXbK:dRN]eO:2/7>;B]7RdgUY1Z@-^,X(\
cS#(G;N/D#]I,,WJDGKWA)FS.-^I()1GPOc:<O]RfI?fX1Y.BSbY+Z4QC#VDSD5E
1[4Y:+SL5?;(NgPda\WJ_YFRRE<E3[UgR5FG(WEXMQc^T^aVF\JFWJF48[_/ZK#b
\6bfV@a4O1_1P6_/@(?Y#(_\]KgQK.+c/Ma]7HeM\\N(Y&EDD>&U6W)CK(/JGc+N
Y@K)Z/[>\bGN._A>H+TaR2L,>Q;161V)<W+Ne=TE0U#/S-5eKH3#-]3_^^L^+(13
?CTIH+Z5/GA9TX)JbSQCVPg;0JY4T#6/KYV_;ZNf[bTCQ>SS\1T:S&EJRM@KA2>)
2R]2AK)O>D?&E3/M\[\gBGAcOYWbZa^1;e[f[)XS)&;1(B=5fE,<db5D65cA#M[g
@ZKdRc>,D7\Nb>NV4X9)W?e6Y[C;YZ[\AVA<,eB@#OF^POX?&SOM?4YgT507GQ;g
c817fHWTGA)5PdFP4&+N&VFCZ^T-0UHZ0HfdU1X2Df57K/N6)N)2:,,#c#a7X1a[
B2?bNPd.WQd.5/=/:XgAc.7V2#U7AC]cF4X(^TA,ZVcEAZAO3<T:4@aFb]=CfW5S
SRE;.f>\[\c9?DH<-cSRe+#LV;A4VV<6>_3d72eOC::IZcIHM3L54_Y8080GC6U?
>&LUdZVSY]YX.37Rf/5QA5GKXC5+,M.INNU8IEQ332/.9;;;TDDLC3H;,6\85\GB
93:daC6A2fZa_=Jb.Kf2WQf6[;fZ;3I2>MX@@OO,Cbda[V]MbeFT)4F:_QS?W+-I
L.#DJRVe1fJd.[S@a#aKRA[)+]WGW(D4&MMdU4Kd.OAT?&6+ab4UVLc\Y+K#a@^-
KEgSQe77Sg)EP)\0435/>I^<gdQO=H-W6Q1>aD^+>R-AP-,&+M?K:JfBdU_Z5LC1
DHJ1=^HeSXX7f7FS_cYPDaG)WW1W3;KA3>DR4V,VN7JZCBQMe4BTBg^GPFVQ.KVG
MXAAf?@^\H+T#.6<3F+f82]#a.KG;[^U>dX/SG.>4?f4c:f8[^J[gTSPJD7Sg4&_
Y)_YWK7ZX]#VCJM&VdZX\A.d\afAW,#COPE>aK_BZN4WFE?3DTXFbYbINE?IA_KP
:;R,f@^R@X,,>UIc>ZF+M2@FFb#XK3R]PIKMP2gSUYS+00KfX?-=/cH]=M3[R).]
VX#K03Od]8;?QLefPCLUA70D#XO]^HUIYVFA^b7DVgWcaH^\<L:dg91Uc^&H/;,3
.P#+-UDW&63W_gJ<NDLN/E\-Hg3XG0S-cacAUc_S_:;D#W5#D?a1.3PS7gM[CJ:;
f7H9Bce^3d8N)3).QU1L8AVaQG>.?aUF^FX0UO&5J@eEGQA0JJgZLIY)VTO]E<)?
38FX:Xe<-UeR:E0DXFN15D5(PF#feC9^DeH/#A(]D46(QY(5b:CK)-CCVe_[+[QS
.2&c9@Ae_1b27J8,I;42b:5-fPZU#RO3W?(7NUG)A(HNP7,4MV7SRE)KRD#VZ)dW
+ZKN0\:)F.c:/LB#/43O=9#BI5C1)a)<6,QTMYVC/#CgA[VL3VZbL7e&\7DCV#Ee
dYHdX@bT+_.^b<@[BJ[UR0>S^BMGC37H^:.>FdLHTL[[4&/3[PSW^C>[;W(44cXE
aNY/P;(f>=?Eb#A8?S=UAE9a<+D=O#J4O+X-IaQbXNL-aXR^1\5HN1e>aMWHV/>g
LZ[gN6DQ?>g2G+Uc:4BF&.^/:F-\Y@d6UJNe\A^=2WYEN<8VY]E\YFD<WEOC:Ief
87KMB#dH6f@K\/EJN?eU@5=MO+Z+W)\WG;5:d(,>R[9.DPG+ULcfA2e3\d)@;EJ1
baMJW0E:Y=\g.d(GHe]A?KLX1,NBd<Z.c15H.-59U(=9&VF)DXNMFDL#4&/;0Nf&
?9K@C4\L@/1KH1=+6Aba[>O6Q_E_&KXQ8eFGYF7GL1+.11\ZCGbA@\0MZ4[,F1b8
A;NaAHW2B:A,:APeTda?6672\fbG9?&FYf60b.3eU.;.HXP/F9V[X@OWJSN=K_Ff
W/B>8.eTA5>O0--&+;fXY8;g0;JEaEA(HfIFg5QdT:5/GX62]DS))R05.>8eC^:/
Y:Q])=QJ<IK_SKP<d;#Me@SRPOW=YG3;9E3U=eXOKVa9&f9HYfITMfJBTDRMbS;3
4+@\J4.:C^4L\PUeU+@&YG-]VI6NM)Z&K<JSK#ME;c\57AKCgJG&D.T6L_N49K/e
]7A@dOP\U,g>[UTW?g?,.d/[BJU;_D7,+DR9#Y/LbTb?C(UG0ZA,377ARcW0[P6.
R<I09PLG70g:JUNb^F>>EN0DZ]QINF9-1F68>e0G<97c>HWdC64R,LXZU-f^0;H_
:7_DS[KGbgC<I(X#^MCAY&27YcY\6S0#a0/(?gBF2<<EaY..]N7-#&8,H:(QZPM;
;-(_[:a<b^9+04CU\,6@S>##:c]La7G3ZT1+K8bJ8JIf@GT\UQ]W9IQcB@;(f)WP
2<Pgg+)F>&:>g(P9b<G/gbX56#2:T1d=JL8Mb0BcSN&dXD#D;LM8G.cFI4U?]fUd
W)TW1;5QCTQ:D\A.7H(M/<g7FKU]>?9YTZd<0fc4b,]<(W4>JLZga>a)4YH2eCBP
3PB5-4DM#:JC+EEg_V,^7PL)\IF)CgCBXa1GN0^IBEQWMQ]>8]=@03@XG)C^2_<#
GW/RR^JTEEG\APK;E-8RbAA(H-89)c?,S8W0b?[6X42O:dNTee:(F),g:+5-F)9;
\PY&#K#1.-f1WFfJUVc\:+=LPEW,\]C5=:-3;S1[aPaPaF9Q,[aSC)M8FDX)O_HC
/C?+M>@74CcdgW6(fDQOG<2#+4f0JGH=FXL/(]^N]5@EV=J>>__gLf;P:69ZIC[7
3SH,URg0@9OQ2^O:\8C^I\[.>Y\4bgE3V^#?+4_BU8cc7-M;=[7;0Q<Ue6060?>g
#@;Pf2EQ?TM\@7c3]8;CV.VO<NAKbP,F.&gVT&SSW?@V8/2NGdQZScY&>W@GI=2)
0#e/@<75>WUY&LYXMY8JSZ12LC^(@T,Na>[J(,-@96a;Q#cR2V/0DXCfR.]),GF3
e(QLgBLOcD:-#gE>L7??A@IAH>SCS^9fW\Q\)YY:f<:;Q#eO@Fee@[JLBTG^-f@)
&d>O>dDL_E[H/WeJC>U])IYOaPQ\QD:=PA,EJ5d=04ebWVX)W@NC\K+ZQa5OKcM7
;eZ6FF./MFWagS.4<CEZM.gCBXcb(QP25Q9d+B8Xa-P;_.WS8U@W:Q:)=/Oe.eDa
4M;SQ704cSW4J4H#73#VJ\a]X7,bfQ.(9cF/\d=GJ<Y-D/GM[5ZaN4)OM0TbJV:,
e,,F:RABTMK71VNM+>ZI68KdJK1B>UB3aC>,If-(P@A78/G#8EcGadJGgON;\;G0
>#bLRKg+^+;W7<_]B9LLVNX4IC.KX^2/0/@#LE9BD.UBH--C+HBE)2@SC)ggbD(N
Q8=&RYUc=#aV_<^-2.>MCN\bHZZ>1B.Z/F7P;.\+-f1NT;\.7#>AL^N-O6g?0-SY
UM5Fb1,;92US=NWZS>G+UX/GX60G8VXOI&46daO_+AG2ZW4gQ^BGS5JXU&a>00=7
.G)=A96J;bPRM8(\\XV,A^UW];/I5;Qe=6C22GHA<Y,)Q=caB04UE.GGg2FH9OHf
[a4V=VPR8aOYB-O1LZZcS3KV3L8LMBIN8+B:#EJ,b/,c+.(?Y+].+fJH1G?[;UH0
BfZDJS0,CB([+;G94[)J[F3QWZW>[AQI,KL+U-g?Q1/LI9E(0T7W?D7g]FSedG@#
cb5P)[YP[f@A2^L5D#=^)<Q3(g.7V7N13KNKc1QMQCDBc+551:Y7N3YPe]K/LQ^Z
U@\&UW1[HPfTAU(OPcU<=1UANG.a64FOGI&,c5FS6.BfMD.,LJNE;,LPVX>5V=NW
4\L9K/1&b]B8:&OH7.YCN>(:++a2-),ge1&?27?Zaab;0f2JcaW#a_KD.0@b32-5
KAbeE@)P):PKNYT;>aNdgG5g3K+@ZR)c-KZ>0R@]3\c@2/G26(eK<a5Z#9HYO7,8
)Z?EBNa.Y;ATUVE;0UC->\:)845ASOg.VU;W>V(QLa?CbL)M(d>O@6PG-IR7A2af
>cTQ0W\ZFBFcC(:ZF281I,Xe=LK--J><5<9H&>+&\e/5<;QV.8&aYHc68?,d<:a#
U;O>(R=g0X7FH+#(XG^W<VXD(A@gJ6[eB)18&c<M4Pd^UCQ3+H\Q4.\>-M&g-M/=
SX_GEB_d98=/Lc4b78L?\Z7+[QQ@O:BVBJf)&TTd[g4gF1D-1>H>=P:&1F,ZBP(_
2e4_]9e5gW^3dea869#PX4FVNCDY_M&7T/P6<1DdTVG-1^V4gc.OgX5Nd],L_6T5
D0a1G2.+@7J+f7VeVI/0RL_C[eLbEYX:[Ne9R&OH//EW)ASc?,)Z/Qd;X1LMd7?0
XR,AGaU9^a4O9F>XL+IMXXV.-.TOS)?8:_)aLJ5@V/SdO/KJfCAIC<KKIM)(UIeG
6G&Y&1<dbA[1CW<;G4B@ZOW;.CfX[.3[,\QG0<Q43&U_P2Se?/1X)L[\UN07eGWe
N+YbCXGV#\2)Nd:]L>76&/b(F&U&-dTBM?[9+[#L)7[2dSKDP7#DK-a](6g42-EB
K:(N>JP545)MTP>U.Y>L-&[_LZTR:I56X5EAcJ0,+&5(X^_EMAXMP:Y,YEc-D?VO
b(@cJP3SP+1Q@e3c+JZRYK0<&1FYA[JMaB@F1DH/C&;^<<Y2AE^?/P@&S^&&SL63
8D7Q55S610aKJCC9@7SBV-HM^^R5JFV_3HQ[Dg\>cHd#J.2)Y7,Q/d#BcU7P[+JE
7=-LMT+_X:7K1T^N>:^GE+\]gX2PdQ^=_5a.,Ne[4XS[X/S8T.YWL&Ia9:[SB_R@
fQ(HQgB1N9f,H.8,E)1UG5?)9TRP:RdI+.FDebE@/K[^&=[ME0,QWa5cIS<;5&K9
=a7H+]29:NT4?TO]R8Xf1+_;GYD<&28J=IgKHJD@D^QS+c9ZE@VK+#8)Z?UY00;7
cI>L#M5X05>[I(PVZ=26aa:)I&[Q>/f7];->+4/7W[>=AZ70C#fUZP_(#9HU7;;I
@-9_W=LJ4Q\=@0?T\Z&dc[JB[5Cb0#RUXI?06X9L:ZEgA5.a^Y]Da:GKG6:&Ydd0
&1:SQa\GWaXFWQ-\e0CN>?-d6C:MW#a120ZE(I+?DEI&d=LW36+)aKaDSF&6E@c/
g@2>RQPI[9:D:cd?D(Za1C0@8eJHY^=>Y/4?WB2S#N6P0&D0P9(MM].3T[KOgT[Y
0>ECecgQ5-3A2c?gUZ^9,_K&4H)^#)09Z;S]bPUbELNT-FZI7-H3>]1,XD&A8JRW
>@I@1K8+ZO/D#93;ED.c1/0U[,b718G.6#fL\<@<-50MCQQD0MQRLZ^Zd^7#15AJ
Z;P5F)V671D=Tb)7I>P[RS(\Te:(_6QN>9D^O1.QUB(G\/^PVHLR1a<C-86=dgEd
c990>\.Z4DV5WN:fHBdM>3dgFf+V<HK>G9L>Ef;X;2HdC:@@#O^+gM3UEcZDe(cc
_VK5ID8N<^C,^;,/Q(1A[9(C_bRe05TdNHJ@H\K,XM;AXNMIWfCYT(M=9dC#U,e[
MYY=C;U2&HBLc5-A.F=(T1(.T(CB=.YA)P9E@E21^O^Kc+8_b?e(JIQaE/cBEP&2
2\7V-gR56ZSS2(#MO04XUV[a5(5R-a>b<PcHD3)P=(^8d]P>G,9b=_6V+6+>782-
.gZD5(1S\W.QZd200;]VXSMHH/D,JQ8Jg659U7_aD>LH0\VO:e8Cec=Md+Vd;+25
b2)7<KDZQ-^:)2-.1M60S9-eHUWV<X5-S,XM-g1Ae<+2B1,=Z2X=9#/Q,BAc\aY)
#e^BG?Z:4g=X&;4FA<VEZ<He:2fTMBX,,e/J3(ZR1XeU8\IbGWF41@(I<UFXg,d(
@5TYQ,/)1a^UOc:7+(=<3,I_b\PXQDC;/E,H#?(V8e(8e,V=#IQQ,H&;F>Y5[_XT
68HNaD]-R9T^5(>cL/6HMf<]:fe3I\R&@fSU]U8J/GVW>SUG5KCKU\OSYNUCDSD[
c.T4@9Y)8<)Dg98[)P0?(a1NIQ7&-<c@LOcdF8KY^IPc)][R4XC^d7NE2:AEV/SS
1F9],\W2YYZ.N+]#D24#HRCW8T3cDe39BJgU&SJ3OOC:WBUYFD5,JH?[B]P:_\(Q
Id7HS3P@68KC=D76>O58X^A53Se0DPbQP08c>b<c?AW8L(_^ZH.I[D_>OGI(&#+K
W4[)K/f03gGK:C_5O\be^FSN(,.=U&6SSZaa0OC_@+F5.L^1YQ7=34G4R2G6.MJP
9ZOHb>W:WgDYPO;FT&[U)3#1&fD>,Ja3JAQe_DfR7PGW[R+T>-UOKd5CG?<\Og\T
[\Q@VgK(dd=OT@+#-C9J7JU?X,a2SKR(,.IaW5geR]U>+U&\PXUOY3<T^E2NIL46
=2UM[9Nc_(MXGHdC\C\HLV638.c0Ub6,LdS-4.+U0B/NQ1a=Fd59cUFe97X<+9LA
0M_SF^6B\cD1UdHg<FQYGW)QMGCK5MP96TgQdJUT9,Y>(3agNQ+ZB7K_VWUdX)#,
6fU6<2.NQD)fC3U.52M(&UZ&PaPCJ[_CO9eEF;N>1;+Je[gWb7Y?^:@fBDb02fON
FG=8:U85c_^#J756&]5gCM<U2+^)_1eg:GfXRe0Y2G4[>FfVAHJbF@aCV)1TbTMf
[1UU[BA0HfC#PNZKAT[+T7+JBJS?.#f[:2&Oe+4XO[C^_^&7aaE\7QEUX1gFgGRE
M?S)?5e+fK-eA/g+(=D:2E+GQ_7G=4QJBe_3-8:_cMW3.G4aLM2OJKG-1D0:.T<a
?c,;<5d(3J4?(7Sb=L=,:<e#3R(g56R05:^?b)^7LRWGMDVAda_V3?85&>^&K;LH
H<G3APZaD1fL&-B2IN39S4;C&E2:aQ5HO?E9>6L,TWFGOOT77bC.G6[AbGFf8(C>
7RL6?H)fLNG@U3,P5T.),]ZRMf684g3NB/CV7aI&5M2<fTf0EZ9b>3#FWf6UEUX+
aV4?DAW=68PFfB9.[YYe0VYN>0_+0A_2#&O42BVN0VA9d#_60.WGIcMXC<0,#=#=
U^e&)ATO\8gg8<S,8WWEZ.?&23eG0R6<8.3Vc0J3_ga@E\O>/D-9?:)GZ8\T58)W
^UKP^Z;)JQ]eO3/O.PB3ZKL4;Q]:LLe3K@HS]22A_&dUH]L@8N0R@Z.IK&S&5&gX
TZ0F3VU8;<R+-M/_b866HO@6_@N[c46K1OCIb17;,V_@7JH#:@e_AVH:>e->P-<0
P@_e6V.-V4I0),WBVKgaF6@^a/VG,Ec4dg(6I0+OgXcXg0\b_SfgF+BK6I.XKVVG
F)_=PcQY/UV8_fa:N3<C9JGEUE^I\<Z3??89W,dKPa@TY-N-(Ibc&1fI/)gVF]><
CM)g>/>+e/L(Bd9aA[R4OfC9.4.^SX\6@H7&T:f5OBB\KGE1;#eE<c#_O:>Ag6(/
=P\_E6\J,ZF32\g;CHB.XOAOXU55\;C_00QZ=QE<GD=JXfRO)1Y)f\B)9&cc6)>N
-<Q<36?_?XVX/fb^HNDSW26b[^4D+IB1UPb.6RBcPbHEV5T@>CA6aH4]49;[<7CG
1<+W-JKc+Dca62U:9ObQUTVM\&f\>9EPHQc(Yg_<,.(UAI2EbMeK6_#PN/HOINS]
>#eaRV8^DN@Q)[KPEdMHNa+7Vea@[A)YL<KY2]1?;gPS_ZV)-&Y>7U[(AN=F07>#
Tc<A(;DD-&O>,NYHaU0QbP:RV7?3>I7^RLBNd@GdDFY&1A>_eUB1&eSI)LU9RL<:
5A[U[b4^bGB=(6VYF+46beZ_R[IgcGgG3Rf#Y2<?[^Db/Wd/_0VM+_^I>)@@^G,O
KEYU:1&8K:GVQdf1@UP1(5R8S6XBYU@3?_UD_-9#?3:^0)4:C43UI3Vf:d<a40d&
#X,\9OS]Q#X?1\KU0+9C2^:66\;W[(U7-</NfYEHIEfBLL;ZbA;OJ?^OaIZMd,([
UDGYR5cEN<##>D_eYJ1UL,Kd<4]D[L.f:P796DI;YE_@OFUA>4R=ca+,.ZIU0>/L
AR2cS._FE<g=fH#W61/<g=113R1\8-&@5^3^[)XE#BR7??W>?-17VK@9[ZHZFUcN
e9g)Nc:JX:,=ZDUFHMDAd@XVK7>FQ/8-S@@\MB-6+BUc<((e3/MO#]Eg]-=]b^)1
-0X&g=42Z8]PD2,[I[GMP+4b;LH/3\aE:a\gXAYP\)L=D@Na9#^T^H[1,FU]5e_L
S/2VO+HZ,3a+F33K#;[<>#PV\)DG_9X[@A&,)PQC]ca=M7&B:6Q@?gLR(daQ9UdD
O@5K.>UDcRPHd&X9]cOMR\H&4D7>e>\YfJ(RL<:#?3aIM)UF,aT><;e40S4ZZ3f_
L5B<MO]OU&d4.de?Q31cFIJDfg@,U?+bMBW#IWD-Tb53G<LM)1S(Y=8(gHL#6FZV
A.2WO?I\gMZY7IOP7P1^.LUNA<Y.FU\&WJBHa9Zd>eB\A=D\=[4L,1@JG[B]_V3^
)@W)DWRc<Z8Z/SX4S\L96a:R6S(U.HF,efL\W])88/(Xdd2CE[93E09AT.VDedH-
Ye?cF=gC^8WWC&M2UaK;25DUc#<8dK?NVLKeM#^I7b7f#Xg55?KX9Jc;7?@EC+-0
2=#B4Y:OH@+F3V^M<^b-@Sf#e)8NT0.[Zb;1@ZG]673<2W29(2Z30Qed2SJW-;H7
W[Q7[c,L>4#c#a61#S=08-_8)V3_OZV0&<Xd]V,d(5LWAGP3aH88.UF2-fNT;Q&;
\+H5M4Y2-b:BR/5+Z@fT#R,>+eAc?7LJQNGM5YXa]aa3(,_XHS2\gS?7/O@-(4LZ
cF+cddG-+fDJT+2I3A7BB:&Q[_g?>fP>7+UgY6Bd.K1A(?L^g4Q^]b_cEE2Je(WK
FX0S]1=gD5[+e.D1bF&c#P-OV+W.?7e31@7)cWZZcbSK\6d>7GHG+?_.411NCL(Q
6@JGdSRG._1GN99WMJ,>gH;P9JN-?eLC2Xd@6)1BZ^J/BGKV4=BSAWE7&#,AbH&R
BGFP-ORb8S^8Bb.8B6-R9K=(c7aID9@B;f<aKK_[+>#JI-W=9MUP(a/+2O64KTM0
EKK8eS9<bEe7#TMLT=RPGb,E9(ECE)fUB\F;2]O5>IYUF9/TOaSB#LfF<A5Ee2HU
e231J)D7YI9YHS3TFB.V.AQW^PDUI1MR(&#1;FC;727S2TS1gTB#H.\CZ0VS;b:D
S6B>G.^d[H9cKXKefPAR][9UM22e4L82O3KHY+SOZ#eT1Y[_e;2=)1:Ld59RVI4)
_5VB@He]WAKf[[SaXK\>;THQR4Q+,2XY\@[N-#1.-2OE]I7TacRH=\CfDaNT0BU1
->U@a177P9GI11bR(.)S[d\EfFO7UdG9A2QBeXg\^X<7F^^UX;0]-);/+O@:1IWM
SDB>aI?B^NbOVF:/^c(?_R[)a&.=S)(SZ^@VUZ]\CGAIX@bSdbZb7[WIUC#\A7B6
H<Laf^>]G49BE&7S3Q.d1)=9U[IOL?76[TUN[+e&:AXA3T7_@=^VB(9OO0X24:M7
]C^b&S\.#[(:aN\\4R=/Sd3H(4P/A?2O2JaP-GLJT3L[1[#/V@-P5P0Xb-3#^O<f
JB?6^C4<FAd.(74b807__(R?dEQRM+=e+=U>X(]X1\c<c;NH<]6L>;V-1[VF>aY,
2.LMAN7]1QHaSI5,0<R,8,BN3KcKS/Z,W.Q(9P=8M.T/6]Z@;G4F/M5<CA\2^fVK
.TB,+N]I/M,gM;K-1c\=5,a-A;F@TM(KJ3-U;DX]<d]O_=V5eQR/VdV<_KQ6[OGF
WI:6L,T0W.3C@?+cZK)DV9D)6#F@9CdPIA,L0U@a<@W120#+YG.Ga+J5S^KZCAL=
E+T&+11b\<-?2(AWGY9]\gA=EO9a&Cb=M+Zb3Z[ZK+G/HY;FJGGQeU]C=M/:_4M-
dQ?YE-b(GJgD\R@O<g.&(=U1\.^\aM>::6Gb^:ZTNC2=BDcA5CLD+0\2=ZA&U3BA
3?FF\T89LBf^f)55c/g:@@Z\MDd1<O?W\1<(Yb=2/_g69:#CI1CK2LQ_R+BbK>2D
EFFZO_PMB\ND/[AZ6B2V=F1B>F:95We2OIg)CUIBA163F[PGS4UfC>7;_;N>D8F9
X&B=GMF1R6G1+N9E@.5<EKVQIgdO[Eed<R68O\X9[dBd(IC<8bBH7^8X_SOVDO0)
W&_6G1J[_2@N;cI38+)8^4B956dR<?.)Pfc:=#VT1,GUSGK[U-[\DO#G9e2WK9C;
cDZW;Wc2VWWU<M;6(C8Yg?LNF(<=[bOAJ;L+;d.X[D;8U,X#f3WO]]LLb#bB,V6]
bb#Z3]A\9f@^=.aB)_d2d[d0Q28JBP?/UQeP,M6Hf@W_HL.0W.(V1fFc-N[+&=^\
PbT&=ST/H[B+88bBKaN^J/ME7Y,2.d:0^:gN0LI8/+\8^YgL2L8:>VNUR5J[_&IF
:Ha>;We4@J3ZJc=F=-9OPb-MJR-><R[Y=1]+UE,O,AQP87A[KJPJ2Z=AZb[MW/]A
/I(#9U_cCa48Ud=Q]\.g<fOe)L&g[O?>J=ZF]J:&g&LEa__(c4>^&KCF\K/beG7]
ALD?FM1]=]:5A6L+(g1O@>=K[aF^BAQ/ea8]AZ<5)-+S_f5?^2b>/SX8^(U]YGP9
0Bg=M:NE.d?/&B=[,>75\Na^NNAN@)^VEQK5S4,c=8)Q>.N@-Je;\Ze-ORJI2O]I
aG3TJ1K=TL<:?IYbF,.9I>>JC^^.+IWa:=F1-70OWdZZWG]>5U0=Q75W0]M-ZDOM
HK3BFCC@L,,5=;WZMCR<Ndd>OTF0EfLJ<\.@U(>?LYQe1B8\,W0TOTI<9E9Y\e<f
Yf/SI2fKGUOaZ_Q:)B)B_Y,R1dOBge8E=&S[R=DcdXQ^_b/-D4MCI<f0XCb:NGXL
eTOOI6H3c2.RJA<5N6GS0dYa8AK\4S,)KUf<AS866F4A8KZF+KB]6XUfe=c(Q-0#
N(O5eH;ecYPXJ#&;ZaEWG/S&NK\\[1R;YCSU:+G6&b34JMJSR[C1()L5POeb&4+A
+WM(\51O[\H+QVY6UH<L3QaGK(A;a.#;DdJVR.V#L)O+bF5_^dIb^3d>TK8\AID@
eK)PAf&U#fA3/U_KR-A>Y6:6YC8;:H+bP>A8+eeb7c\f@P?Zf8?IQ67LOG8cR&TL
/C+6:E2b+#QMcfR@(PTKg)NJUg^T&976+<eL?LW@OZ6=?G#Y>7YC9If15<@--eWG
R.FRZP/2G^KQ]@.[?AZ#NY=#T8-F\C6GI/PI?S6J<FJS:VJJ7aLCQ]gBHb=B;F#c
cC+@R)FRK<W1eWBZ1g[H3/K7A\UX(QAa9f[ZH_gCObdV]I:#5ZI+fBXR44C^P,C5
@=&\FW2R62A;A@BI7L/[ba5=&]0a1TbQCQ#R\1ZYT:NU[T-\_/VG.H#T-A3YcE_\
Z,(f?HV02>.,30T,?/gT3A5H,)2=U[CF0.+IID<RMR\_:E;NSISV7_IXf=0KLKe6
eLZ>\MY8?(W4,D^b1;D7P)283;\E9FN=^e<aX.QTIe@&D86/-;&^+I^=>&3gKKaF
B5.LIY_Ue.=,EgD],7-cdK]HKB?&JK--gN_?0[=SRC?Jg4<3ESSY?JX@S\DN:CO+
2I6cFPK=c=7VH>L?1_^&d\BMe1/V#TdgH^>fg^XI8Cd6aVVfJFUcJ2gfM@Cd9b_2
gZIT_D=L/dRAI4(Ne786Ag7)VE<YDcb<LLa384Z_Zf0fZ.GDYE)U2QU_b)JO-2Z/
E-.aYJ=6f4bV)+HWd_>d@G&6ULReFWBI(G]+,CEYfDfLTB1Q)>^Q]C^V1A/H9-(U
,K3dG@0.fUQUFK,7f4fN#1]f)TY59BEI=AbOL5._d2SE)V<_bXdb^G&O)AQQLVY^
F7XZ@U,W@+FVAH[;V+Fe:G)1\8M+Z:H-T##\dU,]AP-#W>2(_CG5(C+BA20N)42G
\M2[[c:dg-VFL1^3d=gCb>GfJ-KSS0UW;CI?E:d0+]Kd1.T@J)+5e5/W0&_FZH/O
=UPHf8],#L[#0N)8[QDNG+DT,N,EGQNJJ^.1)NdOa6,N1XbD)-4@fSJPB9/d<Kd+
FPUG>-CYBN\?+e.B,e2JHEP-L.]Ub@B>,H-a,ER3\59Nf@62+Tgf/c)XLBQ=<YGA
cJ[6,HH)ZYNMgE@1RDRN:BgZ-e@8UXV\4?-2fHeT\;;FS_?2Q2B<_<YH<(B^B+aP
_;64f1a>NPb1M/5JWK)IO]P2K^)U_\b75<M=e&5L5,FP68b+AX,VI,UWV-OA7:A\
PH2f/+J4^8]ICF:d[>YgM;fWK0T:/6-Ug_39.,:;H+1>[f<>J7+D\f^Z^IY^c3Vb
XYa539[cKc,/Yb6OC[MVK>L/W(AeCF_D3:9f88d#RHCQLJ<4cbM@J.;F\4B0HCI9
?3CdT[GU\21ICZ,df/C)a8NEF9:A>J63RdIF/MGE\X&HaI(SBJ<.0L]RYK^64?c7
/D^5_RTf&E29,./5J:;Yda>0327_Y,XC59_2[KV6:CP:URgMRcYQF=<7:HNRO.c5
[2Z=C/BWSWE=\YdY6-8Fa8/C&6<A>#.a[Y5S1feMObM/Ff8IJ\_T[JOPW8V@3([6
-AETT&d5G;K)?bX:]84HKJ4M_X58)WY<0J1/:S^bX8J8/YTVB3UYDV(LUY1L9O)I
.UW8KH<_A;ZHK5g4F,>6>@e1K_DYW)[2(/L2M&9FW:<0T+V:XeMWZbaI<08)65)2
>Sg<@0R,E,=.P&Z4>@YNa=Z4N[(U&VUH591Y7R=M-MOK\Y^WI^?73eH8]LD[>P7C
FR4E]K4e.:9):f^e0dc6b+_S>RGZ,gP1)a6[UR1VJ+QZVS;2C4[fO=@X<>3<Oa)T
[L]DYfEN[2;R<2e]<AVHaE]V3Z4_QX)QV5_/e/IMP4,e>f&XM@;c@E9(a>S\;O:O
_Z[(f;>B\\D1f9BAH0Mc.7f?1JY&[Y>Xg2gMS/O.Iae([T>C/OSA;M@+E7@_VcH&
B].J[VSXZ:2:5V&<MZ-8__;Y[#40.A;^>[P1#?(NH(W/NUOCCC#-,:W&YG.]0U3P
CB07O1BeA(47Hf[UDA7KG>P:PZ==00?_E^/AI^892XVL6J#_[X<P)7MRS8PMfSY=
U\BOI7?<O=.bAZ4B>\[=6@^6XCbW12D[\U(HUV22I<;6]eT4@eI7eUQS5;H_?O<0
d[Z3L@@)VK>H?,WI\5=dPN[@=<P]&eGCa]48_J:+S^7XOIaW7&-NWF&6SGa05B&N
F21[64[6\(O>cVeNKO]JcYH:TY?QY20?XMT0TI2c^DOLUYOD(5CK(Q7AJ-BTc=B)
TQ\6M=VS#976(7>2aD&K,]e,#IHDa,+4Sg)Q^fIG[GTI\:YZ\UA,ON_]M5cR2f)6
1^D3#(c6=9)J:I,1\c?5gM/&^;,gM&DN&8J=]Q.>XS-&C0KfX31ILXf#TR7=aEGK
U2J_[=^.M@D@a3(2VG9YHM#\gH99&[?G)cJY@?/61DXA9[+AL:Y8&gII-eS,AFN#
/(7.]\Y(eI=T)<.2e_gc+&)T6V9>TM]:8QLQ++.<J;?/IKHQ#gU=UI(WE7WY9JS8
;e<Bf8./OH_>[J2TVNICJ685-<S,TQ20TL/3PdG?aAgS5bL^7S^#B9;9X92_PG??
=K8fSD^.IXVg3C/4]GNA8@ee9dB<Wf8CNd#Qe<A=28\A8_YKNJWXd&88?O3FSCHM
A8+b;US>X;V?YYWDCWQQW5J8F)aJZ/DW8e,+\L@1GbSg310RJAe^3fJ&0\dGNN]2
,e>Pab=_AgEJdL@G?73Z@V.LB7AU+<2IB9TX&USR=NO^f&56\PeTZ^B__<IOaP72
S12,5QM9CWGfad?\QaPa@+)7VJe(GBA0CYO#G@1_3D8GC1])Ac&-b/4<QfDP2ZS#
\/47T7cc9(WEWM)c85#9aJ2]1.M:8E;X.b+JRe2J,4;7=f&[aeX8@R:(YPdVU91S
,JXN1@H+X&ISJP88R1,d6J^:@>A^RT42(LE5V#8Y1P+-+AYBI+_(^3Ug\8\U]3I,
U2#@4,-X2RENc?=B.-8&b4;gIYH:KP&Eb?SR)F#,8OgSPXY3[VOTB;CT/F,-O,_<
9-6g7\6UJE:TS>6^]-XX^N37CF0OT3PG+#5[7YJPg69aba9f)^FFZ[fQOFdP]L1K
KVY+T[#1VPZ0TPW0:A11Jg,/0IKNV7\4X\#951Bd([VfPF@94aNT@J.M0fea,[c<
VaMEX)YF<e>OFKg[/TV7K(b,e75ZMgc67I;K8+JK]V/b;3[7f?\CC_=ADDF-&4R\
0)C1Md@0[Sg.;7&ANRRT3e1+098D(-=\#/[a-<E:fWB[[.ML_,ZFPHQ_e-@g+O_f
DJGaKIV.gH(A_0C3[,PJ@P-OETWTb>?C--#/CVVg82;]E(5><M@4_@d8UCA<aS?;
,BG04_=Og+@SV8>C-=G(Pc/^)^9H9M?=cN96OOb?R3A2[fX-cM(WEMRd>7B8PVVd
@B&.OLbE-Ae<<QL]<1]XQc,g>R;,K>8KF]3:WUWSL0Dad)ddC0-/BA\2PF7,3AX&
A+?TDD2=J[Y(ZJ11HbQ<9K&(U0Q5[TFKZX=e8TPRJPVU-4&MKMS5@8Pe4O],;(\M
dK_&,83VdF[0cdKf&Md0H\J^M7Z>,?f2B3caQ]F0GW?g1^=8C@C8927:_\-O1LT_
Eed?4308aB\QE[HCXT-LI;L=^a=Z6Iac>=S1a<C=dX,>E[L:&7gg0><dATN1IC:@
:Qb/]RZAA-9#6I(LGZB?VZ+F6d]WbXCC]e-;aIc(>^]&K-<@/B@(TR6^:5\K(1Ec
1,eP??f(MEW]WCU:LR?NN4@<fQbRQ=G_&N9,[GH:09U6FBYOP<U&8<9f.Z^-[=Y)
\cYUCJ1>@AY:O(8[Q-T4&AYG1TB79f=)Y:/X_g6[=^WdSYYHU12c3,P0&L7XaaaM
1\2.d0/:A\YOfKGS<WD_gF-bZGMF0O_cX&:XY()TK#GcBC>6VC&H9S;=bX#e,;cV
cV;SQ&ZcG6WKLb[Ma3N0G1@,4&0:T?+09N>M):E7K^U.-DZR1^&6K3+F<:,g=g3H
&)UbC\)V<=f[)^1SB[@gNIYU1+3&SFGYRI<IIAPUV3N91XWB\]4<)S1]_6#N?K[[
&?;V.JAC#6.D3RLUQ<^G=I)8^<P_ZPTEf;RWB#gKVUDX4D-\-d/&#)&[BV2:&)>9
)&V)9Pe;AVa=3_;U?UW1:_dJ<FMD_1.;gPDPB(TV,a0A0K#:a#W9_MVQHeV4AT[Y
XQDb&@\]\9?J&IW^_aI_faSXCI[CL5]\-Tb6H@4]V)8?Y.&YHR.9U(SV?C.W+I^I
f+g]4GJOK<WE/?T.c@X0Q+QA6DYYgf65>K4WV82]^OMK8#<,LRdgA\VbB9K)XE[Y
T\6PLC=&Rc+@Td5H1.+;;AS_--ZN#I9IM9VO01(E)53<I(39VD>S?)adWN23/a^^
K/DeHJ<<G>+>_@,3c\QE#[L]dg78VTYRNFeESS/0.0;)YZTS6e<JPOP,H1-HRK]#
N@[RaGYbH@;[S(5;0>FVbRSJfF2PP[J0b]9aDE:MO\?,TRZ?R.>aL@.gC;FUf+Tg
JD9caZ<M7(-\7Z^/EZ#eaB,I3LBM^a2;FP=0-29#@bL-:A]U#+gE+WLM7c?4&[(3
_Cb2G\^V8T3Kce\)UbNeeN5N)V8N=2<XJZ]B.J<+LF^M.75QRTRVJ\0gABG8fcYa
8ZT3Dd^Sd>I>?6U,H1WFdM-?fg;-5^)D-7J]BPGe/UgN9_PD8-7@fH=KI,Pd3[E6
EfHYH+1aP8^a+?LMLTPI:a>]KH[&]JgCR(UbeJ]^#56<FN\B-_]ZPX&aVSg&6d9Y
1)IG5?S\=T9:cH7KEL/-a?I@W>&T4O6PJUXg@Y>33FfG/#.]:ZU7J4Qf#<Cc417^
E6cA>GVSPZMX,>42+=SMZ.,)Y?/9&>G7b;Q8@HT<.S.K<:)GZ2Fe8SbM])=F>=GM
Z:SPMWW8.<BXXE1g<_-&V@XAND;Z.(X[Y/E^Y>GXdK\EC=(,][]\;CY7>F?M@--S
Q1TQ68&[D9\e+6\S7)e,0dg^BO+ZB>dHa3LOVFbQD?(/Z1<7YUI.3KA.#B(7<&BK
2TFP6a21A_H_8e@3a(7O3U>>JH2H&#+W;fc8=]4:]8QfZ^<I[AC9]O+L??C7Q(Ub
=BAUaHHME)IVJQ3@d(WYDXB(E0?&J^^eZ3X^bI?&N07R>M)&.N@_>dA9JTR(06L9
3L)+E>R?&3RO;^?_F+,b8:L8G#Nd,3B)X_EZ&D(eGHG6W4+FD>VgNS.N(QE<3?&9
/&P-SE,X<,2@D1P3;FH6R90R+/bcN1<P+VJ^\OIPLKH#9;?\BC)2QVOeb?(4N#;A
b-O]EDZX6A&)Sb1MG,OPC5&8aB@gTb[T4-CF]W[+.GI]AL-cU_ODIXf51O6Lf/V?
ZFVP\H]-TQaJW0\DOYC][HJHXgfA-bgIWEgWSJ@S7XWd(PGV+@<G6&OU<>6WYM28
c3e)YHJ5e5dM&S9HU1gJVf]S+X#)@PJ?]._YUJg\Bf;;HbH1;R>(71FZR0]BW4_3
0X3N()3ME<HL8.fc9,&BR.Q,g\;A3X#J@gW]2S:8C/UW+LVa)eCFT5+-S,R/14@F
&gKaF)B)(3:/?]-H7X;J?>:/c#f/JG>.8E4-QGLH0OVXU7.,Oa<QeM5J1+.S-^Y9
)MX,^>33]/S(f>K<M(125:\c.J,@#N6TNHC]&Y-&dUSQ?Rge^?,OfW;J>34X)_5Q
M]#8ONQ=#]YIMI:T]R73G.TEI:EA6Xd;/X9\4ZBK7F5.deeMLS+2YI/BM-e5T28.
BY:;bDH31.MX/#0c:UA8.OPe\W?IN(ZQKL7\aOCG2FCW\Uf1YSYGgY7RL)Y9)VSF
SW1g:^^L]LTd\5debK\0f,c;\f2]-T@f1B[.9YIG/^f,Fb[0+HLIb0aDfIJ=S6eM
7df5/XMOV6/8_[O?ZNP/b@U;IL_OTaZOAYYSXf<V;?5ec1L#PPDJ\g)DfAfNX9SA
0&CXc\BeFg&aeQK<;MZfSb87HS1808NEe:F(BT/9Xf;H:N;EbX?/T^.1JW.+S=(<
DOfd6_CLW_T3COD<::B1SB+_RMVD6g(HYM(?OX)KTU-_[\NK4<LH,K4aUTBSC/P<
(f.DV&e&Q<VNBU6+#1B_,6,^LW=6cCI6YSG;R;-G7FGI8VT[.V,PgL^4G7:^:OS:
9dK#AcI3UFAT[LUB3[=E)[3e(\T\JMMLMX)7(>:MY^6;Z1)RM6KO@b09TUHYDBF;
]EO>Yda6LA,fDG#G:#[;YfL;S<Pe&c#>RP3MUZ9QKVWNWZ.CP;]PA+AL^(TSJ,CE
XW-=]4AcbD66KN\TK7A\>cd&a/\OA+RS0Ac-SL4G.1c,IcI0,5de@E7KX?fF.^VF
bELP9,#-M^XMXG?Zfd\UGADd;=Qd\1aM8gMP+/9M:T@G&;#7NaNV#87]2F0&JE7M
62R[?eQU2;;@5bS3=I.g;JS5KI&f/NQGc^SGJRLAbe_Q8+CM+L5INFb21@A]-S@;
5R/d6<Z&gfQ\Z9&8/_(0C2VBV>bcD&S,g<Y5X[Ue8=0a_PJbBL@Zg;IU<^1W3G\+
C3/4_G)HV2@?]/&C?da;=M>EQM56\41Tfc0M]3=6d-fV)5,(6JY8^>?OF;a)e&2O
DcL4[2P(L[e0ML7DU:b2>(eP8I>+</Z0L<3YIC5I\b?AW;f8gC?L:=L&UD,YGL]_
-dIe3Ya37D7L7NHBLb&L]#CgDC]8B^XS7@@#9RMgHWE?&]^A3ONE=)J+2X7a#1,/
])bDI>A6KPC\34D^Jfc>LFUd8R48)S_O-<Y95g_1YXQb]_YJYbN/f5?.-J&^=U>L
4O1@C32U3R32PEcbeJB^0F@+&/QI/6N0L#PUCP6,WL+N,,[P-=]WbTEG34A(^@a3
:O)^U-\_b0A2@Q+M&XC5Y0U.Z)ZZ&[R(WU6&,Y3X>/G_df1^c/:W@KN^J8,O]#?U
MCWf/N,O/:&)QF&4ERP2W[d6NE8L4>)+)YG1a@0PNG@B.@5ZOSb4)ZO7JX_S@/;)
A2JJH3R4V.,G4,dXG&TWOTYBa7Q40DHMfZ;6&D.RLASZVX2_#([)<E#6SZ1WM@\3
:0N^0XU5+QNDNHXXeBEbWb&5Jc-CB.2?D)aA_L=;R,7)([EL0@D4J8UY_4T-4=d&
2)e7:98STXBUDX5[.#S9=C]ad6^2dQ](f\8VgX772a-Qf]G_3eS<E7?VB.?cD)X\
NYXV+7Wa]5^4XdOMQA3X;9gS?Ke-IK)41=5F;f6:f>?Qg11EV.<GS\_Q?6-LCB[;
M4YU#e30Oc#(5P>B^R+P^E4ME))?2?CRH-VNW:Q+#YR8b]9Z:2aKUA/B+Kb,E,KP
[/@7G:#3fJA.YN;2KeT_aKd>)7G9:F921G;:B<&F5PBF#5^^S9aSG]6Q@;GL>8&[
SLV+HH6YR9XAf)Ibg[GCVd/RO]CTYfc5/;dJVJG1Sc)^eE0SNKAI@?IG];N^U02L
MD((7\(X[ZR93;GJJE,=SJN4;aF>:5/A,a(cbF.)@BBQHcQ02\R@O4gJ8O:a[ce&
FM]dNJ\BWef4U/6f@.03@5(=g=H;@^/XUKTS3UH[C0,ScWX1&TN0T)6Q_3((73<N
@]8GTCZ=Kde\9DF@97Q,LK6K:G;/gU;R5df26^<SF@]J:4F,<L(B<EC@(CU#00-/
=?9SBA\?c1,AL<ab-3]TPFCC#00]TPPHO2#e0g(@T?5[/Y19]PRR?:dc1ZdOO4Lf
X5\bF[)N\^;AMc2_,I-TT91]-g]-OH-3a3cPS@2-dNNS4G,MA^\\6_XI=1_.QFJ)
5_b^SFXVANReRC(=).JRI6GZX#8LA-;N9P_58Tf.;H<^0.7HGL(.IQ.K[HU^-=8B
LCP3dT0GgX>S))W[54D1,/E:Nf&d77)I^)^TO3,Sd<[5^.gU?B0D<GM6^FR1HfaW
(XVHHTT8@e4JaAGAGYVWW\3.A(GR.H#?0f65-ZX-;CW?CX86KRUKB<gR3fRA<6<4
)1?_W/[1ZXWIXBa\&47&eOb&\b#8MOFAOZND7<NZ>:(W(FCe4[5?3G-8-aU7e2&J
CY2=9>U&MeaW),:V</N#AP#CW+IU8O#COAe&:-dY-TcJ8b+X8CKTDYDJJ6:H8&23
:<06PT5Id4LJ(6JaJD#f3)55]CH]R8A6&MP)X\-8O)1[)T/L>_B2K#5USFCP.<OJ
KE9H7>e4(>B#4[6gE:eWfYEgCf?g:L.22V43=VLD33Fa14ca^-+@5JNBDbXS:R7:
0)U=#+P083:]TV=bS8C#KMgBNE69ed&#_S&Oc&XE#>/^XP5DK:[Z7d<,^QZ]?5[\
OW-/;;]aR+5P^)(^2,a8VG-1e7/6U83(C?<gOCb2P7X?#-G]Ba/(:C4Rg=:Hg+7^
(R9#G-(#Uc71;&,[a<W4]8dW\(]<Z)+B,81f+#(5fdJQ5g6B0[LORKe?8D8VN,+E
8DH/@)IU4K+4b/;:Y-J+94X:IB;+J:VLc::7^;]gS.9>.P4Y#^b7NJ3H[2-2&K[V
,BI(EBH0B1F(7,dMI[Q^7,/N+,eKK]P1:K7Y#)LD;V<6]70C0?e#SP4K1bS0YKf\
/K<9[dG@RAEK;9SbYBC/;7[AdZReR5MLMIJ/:@G4g\2UPZ2;@;X8c4]AA#BP&QO\
=d3:BHG[TePBAJP43ZA=(cZ9#_=^8.>LAUA1PeZ1VD\-39^8<)1^a\Hf6E\^\VNQ
:a:NfQ=/4>d4ebcFA^_?<Oa3OPeYc.YH+LUQDKC0@[#\D.U?:MBb^d^&K82I^(M]
+1C>>\3.3g8d<)C,:;JRI6b+E1cP;E]4ATCd>;9M:g0R,,EaP6^FKK9;MN,SX4=S
#4H28Z4PMA96.:>J8AgR6F]FNXO7<IWIOB0&TN?S@GKY?8JJL\-eYV]&?93QF\M?
YgRG(RC(7U2+c+EcGE5dM=4\OGZ)YE^UR-)6+.ID&<a<;=F<HMfM;R/\TW#]0,&#
aE4TX(J=P?bYJV;)PYS=R3DUPCK<)6[)4bR2:8+]RCNGR(;&>gMe:?dgdG4CR,@0
8,(F+TA]5R0_KW)^6\LJ06(R++aff@gZ;&V.&/=7]/SH#D/;M@#:D55,^KcL8.BI
##<#+5VOgdRKLC9Ub:UZ^^-BU4aRA^]-79_6,#]GGN9PXI)4#F3[Fga_L)8dcMHO
94fET,U:F?Z0E3\J08.\f#]Xb27a+bOQ@J<3CdPbML84OQ1E;:37@fRAb8H2Y7=K
>A1FPeY2-=;W>0R0C9_3&Y0Y?@CU8:Y(WaaW4N[K-=V8E=Yd=<[WeUM?[-+TTAK3
gV=_WAB1#^6Q&IY4N&\5;L/8,38EF3-dS:6cgEHWGSW=+SM+G#KF#J0>cVJF3P>Z
fN7#aQWg1DZT_=()[L4KN_e.83UfUM/&]TY7PQ>#3PD796_CR\=CY<<DKVBZef8B
B9.OVHD2]LUQe._,,8KB<,HAQC?c0-ZPN;WV0:GCQPQb??5#(BC[IOC4eCcG1W+Z
@,IY>82SMIGSSHA,Q.0QY;6C/FR.((D90H;?\3E>:Ta)[<>2[NJ1<44W[F^fBUFU
S1@gIA5b+Q024QHJf[N[M=#^.B3)#WUcLJcJe1[7Y+eY1a1WVbPaX9ROXCK57Z78
:^[+gMW^[VUd(EDJ22>;Z,EI5Se:&J/@G(+aE]_YJ&+8+Sf/(W5@&3(H3&,UddYY
IY8+)[e_NcLE_C4W,J93F<P<:f\bR6YP:eee:]ME+5BI1?<L8\32BOTcOOEBT)[;
FFYFg0MI,+=)JEO8L]+]L+]GK?c/08M5RL3Y0gae\:YHX&_)aVaLUZG&+AC#K7ML
CTIJ-P5=\IGK:#_-Z0.[L[[1CI(GFZTHWKT+c2#RI3==@_>c&6Y3&R;e]OUT]INM
03=?ON7HYMG8-PG^Va:cb=\DE+=gVXF6f)B)O^X95EW[]A.=_WV_-a;f5U>)@(/_
?9@;F>d)=dJ@JK6UJ;bHW]/IR)Eb7Sg#\^[^1\HW?=[HF#\LYFCVL0JH\EO>W1\S
P+_5bZX05=N<^RKK-W=6LJg#@bbF\SNQ;S>GH5V&#)T(.GQF[V1X04PRb83\2JMF
V2c1E>GbZPFF(=(SdgBFLe/MFD@?(5^R(0,M^egM=_EAT60]cXH=X[V4>aDF<XB0
+#Q4_7P[gc^<^&3bQ,?ZP:]JFZX(bAP8B3G].E_-/<2WI^+>&CFZ:d,]=&?Q-R1b
)ZSbSc&daM62DJTd\S9SAK8_PN]e#-Ra<\g\^X[T5g0SN4M20^N7/RC\eD>:+bFH
^G6Y/HC79-f,#4:#PT[M,B_9/38R>_EV+B+].Q=8:b#SeNES:9&;+Xa_,7Qe+cD/
aKV(RU]2;E10U&J9f-W0HKc(J@d=+J+I.aFD0G&LC.edQc,7(ON@fdcZZE/O6HG5
]?&6BD&Ba9If.d=_;Ka>.bE_#L-Kg#aOOP9[(F&C[/T_;N&B74O:@SVE#ID3VWe+
,gOVGKBMOG;SGAG3;W1;,3819b5]a+,/YMa6Y::JD&B\LQJ/GU,PX5D?<C.8g6QP
_E[g8F\OgZPT./W,][)@92dPdA))4N&f#.<\aUKUeUAe3R6Z2M9_]_Mge(O@6UDK
geC?2V5_W?K>^TS;G3:JK+b1eN8cV\FEZ[D3f^M&IK3IA2)&WL\A4:>U?P\a)R/>
8Q4=(Hd+QBR5_#Vd+,/BJ.;@@D5RTWg7YXO+e:]\Fef;5e3JI,,[E--RHIXKd<dc
H;>R(EU/MNDKT(51181+=2MO9PFS&g//Ld<4TG&.B?#IY)b>VD([\.IfGF2=.[5K
e#GLXeP2T_/a29EC\73+IEJgO<]YO]/ef75O=)Z@@RVbZ:a37QZDc=2V42-7FRUF
R-C7Jf9440P)cI,EXc,B@9G>GHE4>G,cZCAITdK3-^=-H.8eON+4AR;.+F)M9d_F
[72+NVY4S^W278[W\fbN.VDW,C3+2G:Q=XGQP3>:&,cNRQ^EIWAF&(6:O5Se?TI^
958FOJAG;RbeWV1-X(2fH7Y/)bRDPaR,QM>IfP;T=ZHb_5]eP+9C5>._=Cd-<@;:
L^B]eY^]-FL@1SI.D>Kb;A@GYY.B\<6&4ZIF6N5FB[X_QSE0MLYBA@_<91J_<TQR
d4W61]2MT+S&)NVUC0:)Ba1:#RaNR\WW(2T=7F;T>PPJgNCb<[UTc.0L+=6S^RR&
<MH.BfdNcL?X#IZ?&15>J[_^]S2Z)\&UAE\CJS7<g/[RcdEQ]Cb-U=5-L^0DNPY)
D+(3H8#RXMP1IaV4983)T805BdY9=\VI(0N.CaC7.;73\2?HOMD_@cU5CgQ9PUcC
PKa)H)HfPM4XZ[ZH):UKYF(eN;.,bVZXULO&)g=.,^^L>E+,9LTY22&HC5;JD=bM
dUbI>G.7O+JG.Nd[(QH3-[@)JZT2O&.#=#]U]7:XR+S8Ic(.VGI.L9WV>8N.4,2Y
P\IBFUfe9^M]YH0SK1&IYTBN2]RCZ>]JN[5R,[6QVCP\N:FN<60@+_c:>B)0P5FK
6K<ec5]5U>8J\a[[?:^Ab;D2/Y_1E;-b2+B;76:2]Y[T2I>OB+,1g=DQ2+W)6^TP
V1f+I&1O<&YWOZ,VWG,()A1;,b#S-BL15CT/&MSJKM_8P0_(LN5f)RQQY?N\A/<<
Wd2T4=:2M?XcXDe+,(;),OI>\f+RYV[O^06Z,[c]7dH5Ua_?JRUL8Xb2@EgdVg=:
e>I-8bKZZdWTe+NV>S(aJ,<8NCDYGDL;Y)g54\0EH7W9R1&/6]V-.)_5Ld8_7G9F
;G_LM_2QOI9W[I>V,.CC+H(RC\.CDH8Jd3T1>Za(,C)PLgLD)Gb4MMA,8b/4c<J(
Wg&bcI)8\]e/L-(BS=8,_d9dL)ZVPN<\Y.^eU_AgC>)D@IIYQ@YP.O3^^<&[R<),
_;^N/B)3>3^#T+U6:9_Pg4V52WF45GHDB?IC&0V\6=<(EUPE)A#EMd>1f=Q7X&BN
.<P,(]#\@4H>XKYRfS\Za-?R5I:3\N8RKC@-E&.H:3GD8[X;fLJ)QbI<[KZNTg<g
fD]::9Td\d)5gNR0GX-Z-dK@f>N4^N;[fE0X(OQ-beHV@8#76cW\.IL:^J>H(IPZ
VPGCe=:;Cf^LA/HY;Z7=e>^)3=4S[1TB:^YY-eJV(/LB;L@8?LBa:[A7DDZO-GI=
@AI/V_NaB:U?cEZK2\A3NOT/f_>>IRIW:[c:1Z&Tb^QM0LA_H#S?)?7A&ET33A<_
bfS-WI)1LSf[LWd=S9[SR,SYYZ[<6T/J86&DO(c8A07:>)&B))a+.Q?D7H^+F?Le
.UA]H;BB;B>R\-DU@I14c:F\NVc2YR0QFU6f)C3O(gDcK)db+-XD1gJSW(Z<Ye3L
a_[#ZODd.@f<fUf/Q)-Ba)U]UKf03Hb4c/TN#/_MB#DN[bY5P0.;d[:@E1B,e^&(
<AOc)VIK3#@gF@TIQB/8D//)<):C,G:@+KQ<M6H5(2aZCE0O&BDV45@XEbP_/.b3
Q=BR14eg\L5K#N@95NXU<McI]QDLVN/HVJJg91a?-CH68)cM8Cg._QVY.9IEe5G#
80\efP#YCF\?M3ZI;ATg8bUI5G388SLRG]),.Qf0eD1)J378&IP]f7\@03Vg8B-a
fGNL^6]:BZ.IO#,>O^;YW;XC6NLY#\KOG,T.UX&LDc1Efa5Hg<.Z\BX5&JdF9)/S
35>5J]/W(/RK0TLBOIg;NHN+;4CHf4a@MP_[\7bB,MgC>=.YQ&@R+Odf,Gb&Z37f
eH.909A87Z@aV]=\GbFcFN:7>;W]YU>Y:A_3VBd.0G0J=^;-Ye<41XV#_6Q/[A.D
KYUaL0<TN=d3WW3#8-/BU>>Y&dC_1AX>5gF_U8?HNO4M^P.JZ\)DV2Z]_2W#Y/dR
H@M[GS&.fOHfC7X7Y+D,KGgULU\f8a-&;gACO3.H)dT]/aK]R[=A3bY5e@T8K1F9
3AVKW/=T[O28[Q:E6\_3,D0B\K-))11GFd?UP>CM.@2:0Mb&ZMKfVO?1dH,e2dSB
NX[U>1H_<gB<(L:4V^b[4\LL<K04:4EgTeP<_E]&&8@Ae@P4WZ.57G?C(_JgdB5B
T#fAP3#EH.c_1PN45&PFNOX;YdD#FA<U0)S0F0Ae2Ogf[Kg54d&#W/a3^]?/0LUg
PKYU>=BW>O)egZH849A)aa;0&:HL]HVBXL8b&M>Md^?;(edFS:I10JZf#W,_N0HG
4\5(\<-C<DDgKB>#gXNT@++N/D9_7RY7+^SddC-]IU?_:U>-+N#:gNb\?g8#LRS&
BK]5F;eH_b^Y6&2UaCc#DAOD#_W?T^Ya@=8N30U\LEM1U0E/<DF>(@5BW,1<F4Wb
A7Z3f,8?,:N>_<GYKd5F7;.^gbfa:X7O&a8R]I#cbQ?L),T,56J<&:BO:Oe.?6-9
dA64VH0AM(ZG3,+eSUP<UQP14.H4:ZJT0-:/G->^HcdVc<4O5R6:8HYfcE:9+#dY
0(L<BR4gT&IH0=<J[U[Z&9/4XI>5QREJ<?L.U<ZOU/04RS)>X.0&[YfaB/a:WI+V
(Bg75F+2.__>P&bLXde8M?/9f#19+K2YB9FB.O:=+d_RG.(0[Z0ga+-d-.JeE.QY
)&[I[\Ie+^76JeWSL5.5PY-,6?8#K,[3bU<gOH^6F^YecfBGFZ3DGg&812U@I)(.
-Vf:b8@.ZYH^3+2VY.eG,Og(:R_(f+6fF.cI:/DS5OdLP6>EdZ4BO586A\8,X9g@
4;N5Y7=cO/YX@LPB[JTdU:#)A-g5LXSLR2V:Pa6gMA?:gI:W=,^V/J:Z]:^-5?O+
&.5Ia=ZH5Q>:_+<5N\G,ISKBbC##K92_BG+f,<>,@&T3R?dZ,F83:]d=U\3VTa07
J+^.gI^]7CR>ELg6O((EPMS(4;.(cL_,5L][D&U;Y^M9;^H@Ag\RD4X.<LADYQFe
/+ZANQGHZ9^dD-66)+BQ](#H[?&<55<4L-G\DP#8c+,8[MU)1#C:bfIbBb.8^8M7
U,]I&Q/5BH=JRUT<]fR5IKK&fD9)(=9=WNK(0[ZD28W&S:,T8cA^H7B6<?M3],Qe
;[LG<.C7^M+^]451F<8GC@SGDG_e>7P-UQTS5RU57T)LCLfbaH4[RN.JgNc(02[5
:/HABG0f)K>XDU:;>f9Ha52(I?_TLQ7-Q4<JZ?P+?fM8XN6eGO3\QI,<O0=]=::J
1NcOf.,_8SJG4<^6UVA^CK?:M.^CT0;T3U=,cB;W??2SH(/WMgI/(F?;ZT#T.#AE
Z38(;dPbI1[N#bD>2ecPE997-.T9XY^V.&5,>1?@SN9bXA/O4D@4IE#8_]b/BJKb
EcL9/d3Ad(a)_LAYX?84GR18?PMPT6B=3:eO-9UJVfS-V./J=VK?AVDP&(#7\<FE
37-g/C&5]4)C24?@2#.G.--=Y(1[&<H[#-O;OS5R3<XM&/,(JS5)DVSde]DH7aZ^
TRX6f.J\d^4XJ+RQ8QIDA=8FQY3CROJB\ga@g((\@OWPY:/]]_F)Bc^2eHKPe8#6
LW[\A3PH#0K&=@f]?6JCHM=_+D\H:Rg2Q<A4;U?Bde2O4C<76?,XESC_)ZCEMY\Q
ZGE/KX@2,PBY;=IRYbIKPI+bL_K:?4)3c^EMMO+,.SEHWV<b_I[bPC/Sg,FI(2aX
X<M2)MAXIT7:6\>V:ST#B:4b/W2N\?Q[DD6=OG<Q4e=+JDC.&P7S)ZF=.5##83-8
O5QQK6gHGR=g1@2UY-e7gLC\F,4X1H+c>_BPd89GOPVF;(bd-H\gV?B.Ad/M(_5b
128\b:.g6=CN</QOYdb3<L#Z,X9^)^V7W8OJ,O;#H([&\1QT995-?/5g,,Y?_B<c
FF>aVS&P5@UB(\^TTA@2TB2+@7+Yc3aS:A0Uf+VF<S..7I8gL@Wgb&Ud=BMUQ,0M
6SF[B]SR>;XcT+W5:XWMWg[-Z.2J?Z5IcGJQSe3ZOZC23a36X?K)N?T5E\GDL5@\
-M)1I9NVcgCON1gNBJK[0M/Td:Ee.6.bJ6AG_#P:GEJf4.)-ET1-BB_/,>1(5/OA
=#\WOeMT6WFN#YJRcgP,6=2Kc&bIc&3-7#A;+(0G/bbdUT7()7,/0=/;\Gg7+be0
N92<9O87_6Cf=-E(<S)Da]ca59(M+(dU^##;dG&-+#fTB:6_AJZ+@R24IaF;&QK7
?^5I[H@AW;EDWTOB6X5E4J[1&\7A3Yc9J#MC[\+R=T9U[6ZB)?ZRXB/dCD;<-A\S
P//a_KP^Q[-1_:F:MT?@KbC0PGRe/UC1CZS^U<88/YG4_g_Z#_Vg&^5&Q2P7SL2T
0?YEefAg>Z8<FUSC12b>dWF.>EF0G<(FAG5)URXO2^6;Z>RS5]e]3Q>Pf>C,1##:
/0ZX(0MS1QF(OBP]Mc&IG/RH88Q7.R2B8@W>[C(:YE,Hg-C9H3gMEXP.C2HFdF-MS$
`endprotected
  
  
`protected
bH6)>2XS_Z&UYa7Y\YB7@/T_O1<<C=R^NTaO3G=4E.fD#K]T1G9[5)H#EB9:cP@e
#4E8?=O(W<[\=0[5<78D/\cW#Z/E,?&&XdZ_R9+FHGC?Y_M@UN4J-7DRSW7U\LB8
C?I:EU.Bc)>\/$
`endprotected

//vcs_lic_vip_protect
  `protected
--<J-A5==LQ[(9g0:D,W@eC2QF?X31)74)BHF:+_b7@RSX;TIbKT,(5R&;QTa&M0
P=7,Fa]\7+W0aT.[MT6L55GF)c=ML9IW<XJQ7M]5=2I=&cd2MFZGc#)0CA1g_I@f
bX?a3/S>E(U@3O1A5AQ,1Gg4Y[,UMM>gOTf:MTZF7Y#]V?65dYCdKB&/U+GUc1^T
^gWe,0cX33?FW:ZcH<:ZHVb[@-EB?;W-[I>6IfRS[_CB;ZBP/C,-@]1AYAb?.HcJ
QCIE22MRd+:PWW7?PMZdgNIA:/SLB]L:X/_?V)Qg@<40gKJ.QB5RM8Y7/QHga=_L
VI5<,3X0g[AX)4?OB^054:.5d9)D.b+gcDWGSV65e,]C=[/I#G1>2S)VPWZJ#G/e
bd06;LTT)MZ#Zgd\M>&eJ0\?56.#[NLMTT/+&ONa/T>^RfU,A2W=>48U0a8OZG_-
FDDH#TS<b4Rcd2bYW:<D8V-OSJ=7)X<]<U+=.WfT.^:^M7B&V_]IHV2J+/I2aJbS
2AY07W?&<=370a3fRXUe(H/UV;cG96->C0Vca>0c,gCZdTU(,.]d?AK:]:VgeH:_
O&;3Q[YI#/2gD/:T(4NKF2Mb\,67\Y0&e;a<A5#EF)fST-5/7>)-BcH3<82fb&F5
M30<SeQ.N4?)#/CAU2S&b<c&J8CSJQIM[7J3U>ABDJ5b@/3bScZeI>ba(?068+_Q
MO+9E,HgcZKQUAc9JOWe>S;aR.f>6-E_FIWgA\YYSTgOMATL?JO^7][.VT\L=RG;
KHD94M1MfY2cECT(RRFa<HIf9aD+,GH?.@GPOcX4If0B200^IGa&fO3V]f=a+OD0
LV\3ZYaLHP?O.^^F]+MC<#JBV^UD60\/S8TP[+=K3deB2??/bK@_)8g9-D=MXXTU
^b@-ER:EfY\I\0N=;71LbD+[BN,E.(;G#^Ub96LN6,O3VaJVe(>P4S>Z705b4#:-
J0HQF6=XVH7(ac92b06McG;=MO_W3#MO?79B;\]8c8[D(dZ>K.)<4cd=\S=,U=A5
@E/USPSBO,R7GSbF+9D64E\g=>IPBB,?]-:KAN?/QQ)_)ZA(f[4^TWCR6Ud04eYg
#(/WW9)eVK+3#(?8dgGL#Bb_>&K?=+CdQg:A.>=A1c4-D=T38M:OMO^C,K)1BFbK
].&?TZ(TMQJ3a#>)&D8N&O_8^L.f>;D.NQ59^B+X/(#]dg6<-Ydg]Lg1gPR#,-?8
ffM2_2f;d_N=R[8LdZ;9Y&K>9C]60]8QOOQ)-+>/3Sf+A-<D9Mb[=gJIdL&MJ]O/
A5A_&H&3@8dcCU?@SXC?(MOeb\@b.)<PFL3]W^_5;]a6YR8&+-@DQ2;JF.J,HS3d
Wd,=_[a8d])?TE>.T)WSc?N4P&)H\caWMR[A)3d&b#3]a+=@;)^bNV2+S&J7OHfI
]OXX2cda<XZ1A[bJ3;7-dGFVOI\AC/[M)Eaf)WM-B/QJc<gb5JBC?e?N8/dY@T>_
.bIa&c/(3?NEPSU1Ed:84CDZ?NE[D:(SZ\Lc=bc<.K+8-?56dGEM1)b6gP^a8VZ]
/e?1cKe)ERM#gf?g,HJ.gC)E&LbD[Cd:BYDc(NU2e+_=e;M[2>/+D\\EV^[0VTM&
999:Se(?.LQ?9?Ba#,1YLY9(<V[>fS(/15.>/[45:=R5<_[2eY9=LZ[E<88&(+>H
fQ.+gRGg#HbI8^HY=cS[4?X>V[4a\>b>I.QQ6A<O4=45ARa<#d.D&GD&8fcO@8Ef
NGI^P9g^@a5eAPW_0T&8_S-W1T)KgBE1+9F[/_99XFR@G@S<P+0\2IB1Wd]_L9E[
2H5<6@K[9X]-W&<T4WI=aS+J3T&G[_CE04\BKKSB5\]<GRV4EWKB5N64PdDR8XJ\
f,V<NFS-TF:NP4Nac:^cE@NEX#.(8\f^B>G5MMNgKd7OUNE[LL:F0:[GK5L;TNYe
\;#1IM0,J+(HXW6dM=A&^J:EbPGd\NdcLF(g4S&<aOFeNE6E8XSTD/]<Q@9028b.
VS4bD&VYOBKU#AYL\cb4/SKZeT)BCNI>/05?)\_MeLKcU>7AUWB^gPGg4MY4IRfd
_4^ed;QLG:EF00cPE=L0HUAO\_E3K96\L[X:5A3f?TKgYSVE:P,ZQ[bc@7ACgc8&
>#J.\L;846Z+<]B181XPTd]+4VS7/.36-[RO@\6f?3SY>;;Fa=PbE@/4;<VS</&c
fW\FS99M4;572=eXG&<D26e:-ZCgJYLH61g63RI&8:IE7<)eb^>d-AYNZ@JO8-S&
EH9,.3@EDR<BN#fS?6aK>S=N_bR6IAD=3@NG_^RKGaa<8=N/_N3f\X=FMfVF0_69
A-bV.Z9@QH)O<PR<X)RP/.BN(XF?G<X<LSWV,PY[TACa&_1P;SA,C#J#ZG?FXeRC
0PFCZJV+\YNGgZU3W#XK>MD\U0fCa#?MeT7N\+Z<\N6@AOOW9D>^ddQQP9cI)[@#
-eb/b_C/8Z_\NC=\c18:P/4T<_867MSeaY@P74S/2C5D(/3CR5IWVFSS[5_?CI<E
7a:#3PZ2Y#P(Fa^8+DL([0K)]a#_E[c<?&9V<QHT2M<TN_Y5e15HP6;2_TZW/4IA
[;.;3/QJRML8/=OFVN9)N,0)D=K;bC2]Y7I?NL6NSY+(U)TH37ZI66B>QNB^9f,]
g5DZ6\JeWA_&6fbbI<C0/;fB\[45\FMg23S6d-,g6^]3W9V^0PV=9Pf@fW[@T2I#
8<1@-We/a3(.L;N@K;4>8PXC&^+<:82HZ;PYc)UX/K?LU\f;Ab?I.K7W:4JV+#EP
6);.E8/+JbVaBK8P-HWH@94_:N7_f1L:I:NHDDSSK]5EI/Vf)d:QMN@a/VS8UTMT
9OZ&Efda<QK7ca7(UaP(LV^3)Jcd&RH9NUdNY\FbJ,gX(LT[T&Kg]C5OJHP;fD^4
B+4aY<M\K(@;.JKO&bCB2ef4=?<G6AUZ\2J10+bEU5HKB.LM_6YPf?=P)D1XKO>Q
HE-:>YR12cV)/I&2Uea&b:<7M.F-#b(DfWd?E55&_\0Z)=.0@9MgbSSU.R__^3C[
/L2BMgJBTL4TaR^8J_P+-LU-Bad5U+JAfS@/[3Da6ZS?Q.VV4^;6/2TSSYL[[RJB
DPE+[(&9g47GXF&Adefc0>9[.UM)fd[#BET;W,^/JS1OJKTD>PHY?02ffSfK(<9f
Q5cUPB_ZP.<dFTBVZ>RX+NFOV^)e-L)5O2#MO&8BePC&b_CG]BDI+53IEW3@#Q<@
YTC)#DZIQ0@dPHJH;M=3S5O79ZO(C&;/QX/Z4,:B,PZ.Zd^/dGXXa7R<RKKWF2FB
IDfE&fRD.I&R6IHEc=YIVFKV^\S:O?>:TSfD;2G?,QZ<]_H47(MKO5NQc=>^GO#R
?QI63e&R^01<a_Z4W#FZc-&2G/UeR<NX59I=<>MMQBAD210H#H_D2RBC,=VD=)O0
aQ[735#A2CE86+28;<Q,RI>Nc3;Wf4E)fK9UgF2:?QD:W\YAED@1QdZZ?,L4MGgF
AC,c>-CScI#]d+g0>e_[2.U6LDI(0A,+a1Q=3QW5daVI,]NSN<3Z[Y#P/FMQb+[:
?+Q=<b1/X+42+6+>L::O@ZS0#O.#:3]AORg(U1a695N:Y:f>2(3NLJ<O6A.2WJ[3
@ZYNHY;(TEd<J\e>?D\;G\Q04<(\9e6FZKV\[9CTO9,&?OXc+<.4F=^@7]aV)cH/
9#Ja0F^H5,_2;EJCDeOPT9Xg]:a_R&Kg1:+#A6TKa9JaCLY2JcJHLK5JWd.8a5S\
ZFLT3+54)1E,B=O:CT68AP;9Q[g:OV^bIO>65\SM=A8I4I?^A6,NWQ80M68MJ8)R
:V,=<G\19E_@aB6K<cK28EOCTC+dc8U??0d67c(g,9YHI6DSc)/80P0fA+6g&QMV
#5O>UdK07-e5GFL.P:Y82O+&NQWP(>#J9-JM#_M;ZVS&^/Y/SB2eR:a2d/T/2E90
<a8?Vg3b_R1W-S?QgVa&CY.LfdROR,(d^V^(]GCUc4=(ZSJE(,Z3bD.]]()CKRGZ
6Y&>FU9AdE=05V>#Q&5MU6DS3:;6WaB76EP4C(.NXV_=@6SR0?ZX@dZ,+<<6D@YB
;3@>Re?KH08?O>PI2GU,7P5/]F&:#HY0NXSO6b:2)\fdE[4P,P=/f&gbHZXGCY9W
53eXG]L36^[2EZ-S9^+>-ag4^K5T;U[6NV](H4ZG,T+D1U?aRN7A:gE#Z(N9cB3F
0,,/aRCX.(NB),Kd@6fP&^BX/&/R4Qa1^c./cJ;X^WP<8?C4fH;[(94aSP,P>[E5
Q^JeJ7<)FLTTcEOd,YfZ117_O;>f94WH^.07/U)5TYS@;ZAE8OE25=:;G@+8K7-8
-TKRL?>eZ_UM\I&&BXP@BR9CX@6P27)MKdAT;dTa68P6e->0+TCVJe)R]7VM4N,0
RX@\=-BF[FV2X9L+57>@4e;5=e\F.:X(J?S&=[(=3R9Zf.K?EB4M+b_L\5>3?c)J
1O5M3AHYgP;,?S<NKQ2CR+9-F\bC31H#6f;2eQ2IAG78OH1EP#B&AM7e],D:bFJO
KS8cB6N\.SKMW\H6M2dbRR2Cd^-?N-Y<KY<O]&1a2C2E-V\9XX]8P/bS^_0X9DQd
SC<Y)&[Q;.=@bc:,74/V8Gg4185Rb4TK:8C[JQZT3\H+K2(.P0/gW4AY1LgZG,,\
Z6]CBK\J_\9C.Wg#NBS-/(Sf,[1?,+a;@D(GCBcT7bAUC-22I4I@ZM^G944;Q2UN
[Caf0;SfT#CSH4<_-E)Ya?^8+_)F-ZU\G@(eV/I+g7;K_GF&5dH.a:,JcM[=&c]7
P8Y-XK\b>L[0/_e-]Y7#3)Y_S\/62WULd\c_UQ7,CNOCeUQaP@6+.W5g#L:J@OS2
LV7Za8.M=/K@DG-6XG6RW(17M@U\&424A6=50[@-+I#?\VEY#?PC\Mb25OB?TS99
caIKeCCV(>#+=,e#J-7PVRd3J2QB+LU+]QeHK)?Z11-a<e0NJI3[bS1OC2aea^@I
edQNYcAd>5M9[N\(,[5D=BMV3[Z:&NeIHG.fW+\N;0AJ.V&D43d2dD)::VQ9Wd.;
A(6dNKQbP6@[5RgZC#Nc)eE3BUeZ;.9NB01c?,=Z@,/BUNfL1:?bc=CFWeQQO8VP
J<1DdTS^LT,)c1/c?3aI#aD139H7(KA;3e44[MRbK1?8CN);\dL);7+:\>/:LKMS
@aS6&_WTR3].a\5B06XLE18(YdDHFJVe#24_Y7DH_PHV)P5@f_#I+UKR1VF?2X<G
4;5J/=Rg380^L]597,8f^-Yf&W]8P_Yb^K84,(#K,Jfe+O6P#L?-[>)6XF/<1R:4
I=HLU]L&S.Y,I6+M2XB\Dbb<6A>dQ#dIA7TE_cE&bHE]A]R/MNa<ES8P(/13LMMd
LcDRXX&[(W(7I&9QGCI#BF8HdAL7X@8O);3?U<K)6XB5]K&M>S(I,8-AI#>BB]^C
>P4X)0c/7Z?N(>8_:6<VLFX)Da]/9BAaT&bO2@bgcJ7(R,K?F4>Z2G#a#&UL?Se1
OK#,+2_:]^3WNa<@YJ\dHJMHGJ.I]XVCWbRF,\99?XTXF8HRQ2J_N,4eHN#g4bKH
JYbVX5aXU_R2SX.3-8MRUKTc/QN4^IPT^b_eg#Q_M1^T0N6Y/gZ4,>A/KK2LRX:K
g[HGCV&#X:?-IN^O:RET6:2WJAH/D/=(KOcE-D@WMNHdg)7f0gA:&5Q39e/cWQJR
JJ1U#I]JKUF>GLdAQ6A#866/U-U(-?0IB-IG:Q#M;gJ:#3[Kgg(3\:CYIV7NaVUC
Ld;<7D>\FPGdOPd8(R:B_#.<YZB^=55[<<CEC/6U)JU9b9(/B)\&B29\dFW9NYD,
D;@ZF@>+\?&OFQ26Y3.I7gNf.6E<+.9=Z0@YcQAcM4Z((_c.BVJ#aJ<QcF]#/&LX
3,JQ4]_c8@Q6UdOWV4BP5ZM-ER?1GP\.RKJ+>bPK^2)Ye4UJ#fc-UUH()&T^S^N0
a_>)58.>6/d0^.-JZC)GK.)a_9]&Q1ga,HQ+_c_]6caFZ>KBKc0CH:?A/_LJ04?<
f#U]G6:T,e,W/Vf57&7;E&g176cETRJB]4)=cDSU-LeQF1a0I(4O?Rg5:dg67NT;
E<Q&6EF7@bOP:bVaRX7fg=PeSN6BY6g?be:(LNQ?X[[K7VfAGL3O+<,^=/LZ(0\C
aZce(ZTcDC7/b]RN,S1&P:cgC.0@VQ+a\[-HDZgD06_;:[YC#UA09gM^0V6c6AI8
U,3Ec^1RI,D6dDcXF:@aN#]5AeMO^/3IZX(FJ/NTe^XBW+MG4RY_ddHI4QbeX8JD
).>Ic0:K>La.F7defS-)+Z7,e7a<D+deA,VgJZQYCJ]1Td(?>1B1O&EM0<NTa4D+
cAFR.YFd^(LQF@U.YBYU.#MC-#+IK>9/0QH_2f.TL&E@@1eU)[a?+_b\[;#124.D
cL.#E?/T;#8YX-[1)9D.E[P]E.XGAJIE]^/5>1P[Z@WWVBHbb66TKR8AfY/R7?B7
K[CB4R\;VD#MeCT+RgAIC(T0EY+DW1NEFgMYZ0EfTY1^e<&-8NNDE/]6_K[X-#7C
8#.==O4Tc9cF3PGW:-FR2VW:1Z56K=,,_FR7/RdXW^T,C6=.TZ<^EP@-bJYWgQ65
OG/C1^N4dW&<,/Z\()5J@b\7/)]K\MKT;XL&)QB,fcAP44AF.(ME_-SVL4SM:b8a
BA>8E4P7=dCDMUHR.a8We:,:SdGP]XNDMSHW-FcA0WW4/UI4EcfV=3#Rc(;<]?DJ
:#fZMQY;H8<2RH2WY+B_KgBA;WfV9ZFPJeP>9+B;FVAU/V>Y]7YX<AAKUEHg?RE@
><^M47T]MU[CCKCC1?f/U?[?HMDb]5.IA)>\b)@AAEG?#OeacXZH&^P8EXVRH[Ka
/]^>7aJK^39<c8.dT,gTeQTb-1TPYI?J7^b]T9TgcGc-&+BH8a-)6>.A&[He@:A=
UECd[;P_8L(7<]>(gR@&eAVFU6&.eJM:@5:9BR4W#b/1RgNHJZ1TIW^V>I2A+cVg
3X^^>Z-[/#,&C&#>H,+gUffd7]Q]3f^f-\@2c@JQFH-V?X7T.N<49#\,YD;FQW]a
<cTd?M=76bE@C^XR:[/gCd8f<&\#R]7g<&LI^D=G=W5f4M:?)[J2B1d/GL3bRR:Z
-?-;G,[1Z5gAEI6@.d4<G6B):JZ-+.fM#<QX,MAOEU(9Q#JE=\LVVe31:._BMYb_
WQX<H7YV7Ocf^W)>R0eK8B_V585I:>?IYCQ=5bMHE#UMaXX9(&YHPE2D6G255U;T
]5YHS52#\K,CNbI+5eH5<P?e;-CQ4L&5.IN(D>_9:/b;^38Y:Ba8O3Ud]b78PTFG
_Ge/E0+@LML982BR8)W/ZXKZP26@=59>VO#ADOIRcT_A<O9?f_TggE>\\XCPT_<H
=IPQ_\bW]#&\2EZNPK.<G\<TI[cH0g<\^QEQG4d>GM^eA0f=J>_bC@UDGH+.CZI,
)44>/JS\Cg,,EUHO9?^6]SRS40PV(H2&\>GSX-LGf6C];8Z8?JWdLcXD?;,&PD#a
7bR;S_g]-#b+/>ITF>/0EPYcR3CYU_b[+cNNP64aG>Bf2NX^6F)<g^X<:+J^+-/.
c^M4FL<2TC2+H5QOTBPZELO8=[Ed6e6K.+Y0L],._f8CFd4+@^e>1OB+/8YZ?I@-
3Z#3&5P&<4Za:)5>U?D6g5gVZ,?gVaUeN60SU1_#M73(+ff<^cV[#[E5;Q5?8&)U
P(>.[X(6&#SD7?EH;<E[TZ9YMd2FB#^)fgI2P/K:NN[[,(RG=OSRVP#5#=[<d/Z.
d;Y5-#:8N8TH0g.g47=<9&]B>@=J_58N+PDNV?6QP7[PGbEF6Y2+UL-:((I@KR5:
eBO:>e(SddO^aR(f7-;YBC5cdQ^Q]de+VG)D<.TRDGN1H?M1Z4([0:4341Wc+HL-
<45d#807Ibb:V:6N,b-:F_&I8Y+cf48#.E<3OD1>bOJ,(XOAN8gZ+L>_da]<TL-C
,)<^T5N>,?#CI;,\cEK][P^ZK287GKPGH?@A@O;P-=+XWI>.B@>2R/\TNL?_2>&[
\NKB^=<CK)9OKJ=EDe^#T_A_#3(P6[5#UZ]V4]R](0>.]F1OWQU.K2=<R(<f67O+
+K=BQOO&c>6T5ZEDX,A^RPUFM_^O#ZgZFR\#cF22W8#Z8:8bG#D3C:<@O(P,=[7?
(G2Y<_Q^/?:(+2G+2/K(F^6I90EEL^SMPJD>,cYP23A&S3Qf6JG1IEb[=E;_,NJ0
aS)6#7=,RZG:S&9fAO4H6ZO/-<UacMJS7DIM(B:HA_f?dNe+=FJUP_.YTc910<KK
V0VH_^/3ZI4c\\.O;7dI7/f8Yg<-0(H:1^Qe&622/AO/1[a;K[U5>V;2fCM4[<&G
^PE=[(aT;+d2@ZL(\EV9+@,UGQBZG&Gc^0<CFb>D&U,dS;>M>O:IdL&5gQKd3-@?
IFAOMdS8?TH0c;U/[7Ob>>W;=#?GP=FIgb9MSC]NL8/#[Q,dS,P=ANTZ\aQ]KKFc
)F=WTce0ATWJ\dRP+a/IaSZ7dF99UM,0_80KOAZR\WV#;YT:e75I8K;/QM_N.FbM
H_e-cdQ4B=YF@615JF1;AMOJ,+PY(5_X>DRM)De-Ve9FX_:)/0XLSB&??A?\37UM
YGZ^>GbDKOTR:QZ@?J=&S]]Sf)Y/DM]6Xd;TGGEJ8)-e7X7MO_SDORN#U8G,F/T[
94OQQEYU.dNDFZB8WXNAN;A.dWQX<\e:ZQFY>]_cAJ\P80?Tf9f.Ec7\-A>QcSFY
D5GUUA=D5;S[5XDQd_WZf8C\TWX3SfA/NIQ_]P-c,<cZ,?E(G:AOfHeJa0=&].IJ
H)CA,FJEa[HR?WD7.IdOO4c_OELR>Yf(?_b@MAEQD&C99\NX>BP#7D9VP4IR>5JY
?))LOQ;YB.3]T,_F&CG,ZU[2G=-=+XcG2ID?LgHf;J@)D<>71]G_9NVgT&7^(1O@
Z?Q4ME)F[<Ea^^0O/8&.fZI+,UHA.4:EM//UEYD5D=AL-5f&Z0/Ze=4Y8)dJCQ4;
(J?:G[dC2[Pg^cKC&OL/CX-07@Cg:S:>P]IS@M<P7SX:3CU>IRC\eFWL68:4KS@.
FPYK+AFU:]D+ZVNZ2:D\0g2_ee[IL+f]OB_5P&D271U(C(<7YaDY?^XL<-96&OWU
.XVg#NeN?[4]O_bT@^a?1P,E5e\@\._ISdRY0(P2S;=Q+-aX8@O]NF/P6WI3.UKE
?7DPac(#^.^K)gc2RA<gP5M2F8UGRJ^]MHY3LA9NM3?J,6>)8=_=RC_[64KHP(^P
3N1+?:0gJ.>E>L&J2;PPI1]\?R+W+EXE5Q/Me6(,c.9ZS8J7cMg<<CD4_\-HDJ+=
GHKeQ-f:X_fX>UEV.73IU18_]0EQ5TO@9+[L=DcKLEQE4#cJL6HU](1VdM#JYN5B
LO\AB9ZM._;Z)U&CR)S@8Eb#/=H8O+BgXFYZ7JA8?I)ZFZ<2K=bLCS0OOUCX1bX9
X&Q8J:.3VLR6eK)&>A:E=?N^(O=8],a[0801:[RO031ebKA02+N4WFX9bAc\@N[?
Y56I@U,-Z-U70QPf;J58-\H;8HO.M?-YSgB8I5TDCP6&GgK.+5CIBK7&.9R32c9L
&b;8P?&BMNR2:D4eFT(8>1&.dcgREAT.H\EYa.]B4BPZJ@KLHcZgc/T67R8@^/]1
cH-3SX@ggY&J3;dbV8I>F_Y,/-eeJdFeN7U:/P4AR5SW9717WL\O6MfFYHLZ99(H
KE?E#bZNE\LgMR#CF7S#:bC1U291-[RUF?dL2;,M<-)U4V>K<N98^RUYXO<b&GOE
ESWY.dNB.5:\O9EccIX9-dQWX[_ZY(RSSYffQ^+AE7B<Q,F+eA00YT(UKXTgGe0:
DH]NHSEBG)eXOD];0J]g#):W+0P.#<L[ARNO8Y.^]I2Y^/<F#DH8#.aUBTgTSP=6
)_;B9#[+#.3\?MU/XD15_Rg\,ZWO[+H)KIN0A?\XfF>:AP1CQB)#[4aR,)3L\VD8
TDaY>;3LUe>c07a5Q>,K28dU8RBd#ZADN=7=M1VU#\0X-2AgAK_FPQ@^]FSA#SMX
Ug8(QYQ(+>[XV04X=PO=-CS9=[GYRI]Y7M4J?g?LUS<XP6O>?@0^QfB_X\D@W_JH
VT,Q?O/AKPf1?A<Z7S.VSK(>C,QG,B9a+SY@]-KWABYXUT87CECPF.e<]R-]#0I6
A>J,dHS_<JgZ6PXIR4-J&M737O<^fa6-:gJ(9:d#7C9-;917AgTYPU<ZGFDE>J:b
GH7^WGf:@B(99M2A(^[2T(BYegK5#BEY.GVH:WI4I;&Zgc7G@-NE6)#59fKJ;1dA
gEJTYR<8=>05>?D]Y2^Z^N46aYNE-F7/<VgITW[Zb/]fc5UILWZ_XfEN47J0(ADV
A@gO4]2,ANAVcCOBKd^RN;N/2<NFgE0@8HQI2T52cS..#02EW-[eAe87f_L#3..)
4baeX4Z6Ma+Z0e2Q,LP\;UMZOE<J4GK9=Rf8]cQPDV=RAfTE\0;P8G<fYdT?ZLTI
fMfXR9XK5WJ4f2S33TB]3SOM@DeK\[95G/I7+146bS:ZcFBM+RCU]ZJZ)6Dc7082
NOBaHN:W=P[ce,6_Lb7E1PgT6SRRW5;T=P[;@:WD6[Q+&dJ1aJ/Oa<KO@L3P[<)G
;4TJW)[ENBK:LT])F8SQ[OcF-:,(X(&E=90DY3T@U>DO[JR\1(g=XBZBeI8e\U7?
4f<eF.;^&g)<@(Y,+)Dd+]7bQJP]S0eHU1NEeb><;=bYGEB=3^AF3M,4AMaOZdP]
U,[[Ec5<Cc40g7>B2.:R+)CK/e3XEAQ/RCb_3H7WS(adU?8Y2UAF-5OCP(T60e2[
_FBPP1C3[_N)L?^#PQQeZ0T1LQB60+1\SLfYHd^C3GB<X/[#D.8bC9UTEZTA@@;F
4<&LGW6g1&6-]CK3ba:+^J>7WDV/.#(5Je&5Se7@3?e4RX3SXX-+BC+Z[b&N3>;8
c4>C_a6IOR.?^3LQ0bH(GYXa6K+&&5>N-U3]J4Je^K;0(;(T@FP8MJ#Q&][\0&IQ
2FK.M_J8/AQbN[;bQ3gHXCAc4<SEKV1c3S61AEB4<)N\QHT3GY-+.KgfecW#?eJc
T;+V49AbM[4b_[e@53K3CDXAM)K]AR^H)REAV5J&E0NRf3_GIRW=/YF;/E^N31Ic
1bB@4:E9>dA[-c9078aCLD]2.&,RB.e:Zdb5>e<[V2>U98Z^J^Y;;[U>>G1dC#C^
U([3E:29E]3a-dL1M9B&Q),_]U)fg=1SQ2fN<K8[=US&HBJ9=>-9Z+&9gU(K5[B7
.MK+?4.-+<+.eHQ^T5.eP]Z_\O4J.]V7(S-GT9NX)0[ZWPRRb79U-CO8X(a0?O9Z
5dfTAYRTY3>S^WQYdI6V/T9+Ba\a0C.e;P:3b:f7F<7-.DJbbU4#<J&BU+M4dXH@
5_c;>_da=,0BG-EGV)Z6II#e52/f.KTfOFdCO3d#/Y),F+EB+6A-<f]#V@XA>6=/
G+&SGg^,^)(dE]@]FF(O.K[3Tb^NAG0C@:M3A&VfF&SB].-&JE:8f+AEIXe96dP-
?e)J)?Yf#a<WSHY5:W=[g_Q32D8BZPAA&SWW]3?,\P9(U=S=N44gbNf\C1D83e7M
.MeS^Y-17F+bc+[2^7/JF7>^7T.dO(F5)aYS-&cgK;(DdZY_&<f/C#U^/S]3RXL<
)B?fB8HKcMI8ZYYB#FZg@Dc0D@@d0]B3\3cQ3>\PX;K@^c47\67LEC<>]g<deU<L
[WFgc@cHa7gY7-;4HEDE8F#HLK0g1=,,3gDbR<1>RBI]G&(D^8F2YT2RbVMWcP6E
(gR>>Q=.&O7e9.2\1).2+.-[/Qf5U)I=F<MIS+>GNP)c1AF-28_5\Y,6K&X+LIPJ
(eT&VP+:@bD5><&A=@CAc1U(?]e+eX\38V#8O]A]3TABT5#B/KHgQ<cad<][438?
b-\\QKb460(aWcA[B)g7DJ1_Jf\@5eG>05H(0P,Mb+9B&RgMHPD;eU3RGc<;eXOM
A-7ULaAP,K1H3N,RLEU[LAM<AQB53dAg@XeZMg^Fg8VEY5GOW3;-A:CRNW#\I@U.
<<Y<ZD#c-[M,_d]\+8=JR(f&g5A6;4Z+afDJEMedHZEfL-Sg0:&2[64HP_DM,a7F
_gT/<N@?,O)H.0PaD-&XRRXR.+GNXZ&+eABW=LL(^&OfZ6:,+(9BX:\]MOJ#91VE
2gZa3eQe&Z772_7d,&>-^]<G1J#J/NDN/DJC9)#X#G7-BG#fA&0R.e+QVX/QH+OP
)KS</aE/AGZeN.<=beeb>N?KSO)==[#LO9E<GUFVEYO,)=8d4?EW0:(_FS34+^C#
?S6<I[g99Ed25YBMBUOc?=?ME?7bBg:=FS#aK>64KH2W?MS44D;UcH11ZF.OA;K4
fYMeF_?G90521JGEMUZ44VG.>5.K[>V_85e=OR]C9&QFU81Oc/bf+8I+WLTY>W,[
dAM.YQ&RASSb+WdF/:V0)^&979-MXOc8,&7R9/34PO@5DVXAI(-RgFY]1M0.b9g&
6YZcJFRPg&d2O-c01H(G8e7GaSYL=8[/F(QVDIODLd@F9.],>X[+W00WeaC+]&FV
b]SWP^SAa<gUY(#85dc6#P_K\14-Gb.]/c_cH[(L/d]>0A7FNN^U0[#FP1&J&+K(
dI7WQCEYC#>B>BURYa3SW#_&X1;;SgS[0OR8H/-1X(4)V-6JWTC[KfJ,OO>XE=H.
F=/cZ&6UgJ[KYZTTVD>-K1PUWP02aYJ?IY^H.PJ?8DgX5g)/d&b<:VANb_]d1fE\
L(gB<WFJCYS>WPSAUZR>eTcLbPdB0>E)=Q1JEF&XDG1TA@2?SVJ(/J)fN8[+NPZK
/2Z?:#H2O#A\^K7RUe/Z&J2N^R\.ba8Z<@[4e#Q(D(aI0fNLLBW+2LGOAO>Z)E<C
@_g/H8WJ2.=WdA[:H\;XY_V^TfGAT&&_.2Z40CX@EJZO>?TXW8C^,YLc@@?cP9,?
,&1_BSLA0E;C7D[-:R,O=,RXHS1#N@\=UaXHKf),:YW.R+=f#(;DU:Y,(Y-f)98V
_Uba>ILOMgA(Z.bL2fTI3H-a_+Ga)3dET<>a?,Dd7BQ;8W\+d:,\[6WM@8B@>a:O
.)B/K7^(eDN]H5T\U1FM4Va?=J#R(<2NETZ(J77/#D<4d9^a@?<>DCMdES5^M^SH
:LO.5FDT-,F<8Z\BXLH8eKbMLVfJ>0<2;F9K9LA6\U@6R#0Z3/HS^9=P468[<#f@
&Xe[bAG^ZG(//U=U?WF:TZG4K;K2G8c;JPb>;e;/<GL6F$
`endprotected


`endif // GUARD_SVT_AHB_SYSTEM_ENV_SV
