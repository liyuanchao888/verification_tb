//===============================================================
//Copyright (c): ALL rights reserved. 
//                                                                 
//  Create by:
//      Email:
//       Date:
//   Filename:
//Description:
//    Version:
//Last Change:
//                                                                 
//===============================================================
                                                                 
`ifndef CR_DEMO_BUILD__SV
`define CR_DEMO_BUILD__SV


//m_pcie_subenv = cr_pcie_subenv::type_id::create("m_pcie_subenv",this);

//this.m_ctrl_regmodel0=ral_lpddr_ctl_top::type_id::create("ctl_regmodel0",,get_full_name());
//this.m_ctrl_regmodel0.configure(this,"");
//this.m_ctrl_regmodel0.build();
//this.cpuss_map.add_submap(this.m_ctl_regmodel0.default_map,`DDRCTRL0_APB3_BASE_ADDR);

`endif
