
`ifndef GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV

typedef class svt_amba_system_configuration;  

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
udx2srhaA1qZzSKsDk2yWFm2fxtypXMrPt8SAK9H34HoYniBGg/OWuEB3Zgsp2uE
CuzsD+M6zEKMFG3diNZRj46uIAwMTg8sOAPsFaspY34dEEB4ZnnpwqEssUwFlAtx
lcACH1SHr/cMOa/eDy5HDGGg3kBdVT9VA7At6mnPaBWm52SO+sMffg==
//pragma protect end_key_block
//pragma protect digest_block
ca214nbto/x5mlexKouJGljJjDo=
//pragma protect end_digest_block
//pragma protect data_block
QOA3NkRIefEh/ZIgPIR8eVFMWt38E1dZpXhjM47NZhRSV+sAkKvzerRm8e/bobVH
Gd649cU//qw/OjQfjIewJEpcz+s2pbm4jUxq8a3bZACKbZbGlNv/9DLKD35415eU
VBQBoDnrStnMaS2b43JDRmn56pitsNAXoZBEBdctAiel0ZCZHyepusdbwbOChzkQ
715M6Xq6wP8E8368o7hiFv4FLPmDdwtxhLdbDDDrl62FYKvoqmz9gWx5XZi6D+F/
Xoeo4kTGY6tCLB/IL5fjBsCuaHZm2dUUfQwbN5FpgXe7DEa09ngzxDTJt/tZJvkG
2WS0Pv0bUYfbpVZn8KAcSyAXRoUyiu7nFvTYxkR3eLy7veNRgk7rIBt0n7sC5P6x
liCTe6FjFMdsfxm6v70nYbGNCo3L3nV/CBkeQsG1RZ9odkKnFo6+9MEKksutv40N
Q3/wtiOzf5I7yGhKNskt8dAoP8lyYAlVscllF9RQsM++8nFQTvF0itIibhnAXaxQ
2yttXfJNavzrGn2AO2MFVl5DpfwW4Y0D4tJi9xTiZuXnUltzd406oMBYJ+JZdoH3
2DJBDgzTtN/Pir5TmAx+MVIN03xlNGzPw70dPyWbl7sqhETZnvt9CsGkSA2EkXFD
d3+6CgMxhCIjQizAh7pfxjctNhcLDzIJ3XIi3PEFJCLS7rlc9Et75X9JQ9V36rex
TqIPKiC5G83A91DSo1kjom08QvbphrsXDf3i99NcT80qPpPVDlaCqAF4tFk8hq6D
rwHROBx+QjsvQGKoe4cbsFz4fAEVF3DuY+0z/B2ZpbJ+/0O2KWkZcz2SPYE5Ebge
BcvM+qnjanphY6KENdMpqahd+3UrEz6hOq92vic86hq3CFpM5iiqqz9GjWahr0MX
/cYHgVH6q5fPvzA2jUp4xvtj8SsOk4SzyLtBUgVeYe1cpgYDhs1UCMpPAy7/K90O
0/T/gJYn1OEZwrBez0MbmrE0lWwjBt3Q/UToAMoeoCKrQkQ9u19s98GjbL3a2nN5
8kpU9OsNPYMRessxvlNCKh8Ht8rMasn+rPavOiFamR+kHaxbyhdzuY931lajEMjB
bQMp1DxXQtResdBYk7YnjV6Vn0Ox2noR0+U5PLqb9XaZIcucLSOBF2iQ7KsSZQ9+
4xYV+acSTFKsQoc6s8QtAS5voiDMisEK4VuqUX1KNtrtYmoaFxPtw9hRsMIlFa3n
nlPu2Kj4BRrXH3dsjoDKm3ysmN6SKXADi+fhkNQh2k4tGrf3vZH+l2y+ixVJa+C4
xBvK0M194Tn7vqtHPFj09t83m3uwtaGcYljKPsacn2t8WRGpRM+aSKDqnbUayaue
au7JDDsbZQqGVnU2ER4zaRGnytCZ3yF1nFREnWRiA1HK8wRfnIuuoK6NyiN3R70w
1byq3EKRetNgu4R+5ABijvjynEVsdBIw6s3/9/q1feANk2vBzXFN82NUXFbeLRDc
UXh3g8s8M7SV6Nj4UMzkaDkJZ+W2zJCnHB3aJqCMu4H/Rd7OX7h1l2x6rWvAYfEU
D8oPnQd0hDIrWucn7uohmF6NnjYZPfdr3OGWvpF7netas0YXVAv1D9126pXNbHhG
LFPIFbYCm/KR9Rr5cqz4JXEdKRCBqaCm3h671q2xAf2WSfm9dd27jINHktSlxebF
q7PKqiayKb+MwI4DLkzoyGPoZTJCs9+elm5E/aL2fsPY5LnsbmaNOMVa1QvbLhCV
efvefE16UVvYESi4rKEP9gDb8RxY9dIYh8b56a3ijyWUs1ueQqt5i4eJYDtJqpfb
GXnJmIt3BSORdYi0BdDv+zkPCIKyf3twkQ6BS2ixnKJv4kklvozvJIWyxzw/CTzN
4y0Hsc91qdUrfiYnJeP9n7a2+K9eSw+xfyzSbgfapOpAfVuFN+0ESS60jPyOiTU/
YoJKfoYSFjogqGwLW6I5hcl0k9Hj0N4db1yVZVuWT3YKnMmOuhnENX12HLE1FRTz
EPhpRd3PiaNo6FBZM83Fb+8XEtEzOqXOYzOzz2Fn8OrygmSnodVDDV48WC1tLiak
CZrdHvw0em8Y3cqumst/O7h338pQwDvDMss+9zyWhj2gJHKDJQ3TfYMN0Or1byMG
ansZ/p7N7oyFQX0Iq+dIWd5bptR6SD/BBxclcUl+/mBWBD1PXtM6uw87jUFoNjlz
LEORVQaFaVgwIuzF2xtERLBMfxb3FZinFU+V/KUvg9OECJdInGgoe3ZZeh46f2Ry
iFNK/q9U528XuulzLlt5aEr7ixyKGp5zyXb+wob+Qi6d+pcR+X1K6TJuI2Ng19SJ
EZiS6cX1bKvrSAHCOl/1SDef3RF9XgjAr+1bwMsKIdkfQnLpd3UWzjAFqMV2UhA8
4XFtPOslO3UJFjF44iOuDIFuM77ZBcAC1Nn2x0qEv/An8ANa4bvOz0UERV69shhQ
5BjVSSHlBtKNBCC34aMOBpLAePu2VuvFd12UT2jsaZgeZF38Nz47hIkvNhKASNkN
ja+uISs8PcPeu7A6Uf1o8WvEJicfYMxLrY8aaMwSeqKoTlFmBGz9eUt8WXfg/OA/
oQQJqDNiSYT1JmxnCA7OeQRU0YRw/gvOr/mUvY+3EQDRzfCrq7wcvuZUQha1HdTl
Myx8/oVTrXFkmj2njN6/Bb16NbZDbdjgf1v4btkOJYfgywdWLfsfWKrAudzcu1jn
zFQMD2WmJ1qYD33FBQLbBj0JqPKzgI/Q9/c57FDF1d6gsm5PFWV3aOuLMRVHxpKx
A6NLzshEgjJE0SC87rkmWOmXMS5/Ay8ifEFvuWn4bl8nXRDtmF9zf8dpRdMgQREl
/mRtSmXngHvRZ0ESIcDp6l4B5OcqLbjB9UUVYeAO/xixS159lUfy8W+vMRjs6g8W
Wylvizmaf0N9SsZWU/vcSu076adP2dayszCOOFrDE20P/P1INUKNvG14QU1xxcL0
3V55DXI1Ewiml/ReEWOzyfxyB7SR0ISFJFOpejnUxj0puaumFbj7Bg0gAtpisLN5
L0B4R7v+ZwoHMgwMOUIN4wjoAImI3OWTLduu2KA4Y33DL9JbVlWvQrIFRuSxC095

//pragma protect end_data_block
//pragma protect digest_block
O/uADRnZCSbrjnlSAzgI7VP5ziU=
//pragma protect end_digest_block
//pragma protect end_protected

`include "svt_amba_defines.svi"

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tf8oBAskK11ubefR5vzOIFBc6NROMjwyU2UY4MzZ+hA1FSSdb0DBoBpBVmgCRR0E
Q/P9y2Sa/VU0q1dw6s8HF0x6qJxxZP2jUA7Y6m/0kdgJ+18mxK3AGAt9MahGghES
ricDkZUTCtdt+aQOPigZbNmrJGBeV9TlVwoi3fiNUOP3cI6p+k878Q==
//pragma protect end_key_block
//pragma protect digest_block
0UemS03OEffggZVCWHbZScSuA0M=
//pragma protect end_digest_block
//pragma protect data_block
oySt1vUsi6ylLr7lD6dpSomcBzMLEu5prLnL3zPnN031cJJEy04/WwTqlQzwdbDq
NaWc+cnzzB8f4+kifuKmAk5wUYqSJJl67OPR0Hqj3NSnMMxtro1Fv436khpZVsAz
5wa+ILqQjvjyewIuBHwghbBBu9ln/uJuZercAT9lCJ24oeHu9pQlAb4l6QZf/JFj
6v4DWC9Y9CrnsPykfs1A3SjKgSOayccBMdSJaN4M4OJudmly3/Sx0B4keBiblBZQ
sbcmofC6pJpMB2yCacbFp2ipLVanB4THAbzrav57zZIwaGqcr2/tuwn3gUeU37Bk
MOU2LDoRxYzYwnrdm0sAOZl/6YFuI7kGzP8hE986tuTglOBaAL6jpXhLiJFrH5tC
hmT4Bt5aUSqdJnV8qvcC9I8ws5Y2mjB+sH1tXlJj+XicVAumplJPd17tDqnGnLRU
f4TcJvzqayqtdX6L4NohyLb/0ovGpjJwdqdRTRrKTo02QfUNWFAUC+XHzyBpazCW
XlxIWoTPU1EjfHoO6yFIz8WN0E2voEFJApbyt2CPqOq6lPuPWpJEPtnGxOwTT7iz
oPaHvLh/OkiA1s7AzwCk+p5dEmTb64HiYf0gl84vUS3GB12PbXeW3KeDn2KxTRke
RP1ZqyE7Y8TRU/pLRZ0nzsBJxBVhIj4pp20/xO6jcyE3I0Hkb/YDyhBN4A5vXn6o
n+zKWShgB3LrpjXu56JC02n1Td6JUlUmQU9QOljwSk8wOqJjroZWskC39JUvR9Xn
/mmSpw9g77VxcCOS2HpNUg/hftkySZEKfPUU+wwAiEAob88zylwYBicA2OYj9VeG
fvWkemYOPlqdRCQZk6umBT3rvPLvh8BABa/k6BEDH6O7LjeeH43Rjb7w7opsjmdJ
Z0xNSIW+vD84y836L382ZaiUuCVhtZ0C6K7b1QMSwBuPREQ0qDW4IK6XzgkxCHJv
m4sYR3BzVzaXfDJvyg3blPyPJTdDg4Oo4Lo1wJ8pmDzdFWgVVrKtaJ2PCykBqTXg
C881FKWxP+XZalFRVImSGqbEzQpq26Km8XJB6F2Tp/WdQcsSdgmI5dGTvreCRovJ
OEY6fhxgi+fwF9zHKaiGXMeq0Lzvk0a5js0ZsThRwqtyE7kqCYmWiBF3p5m2K+jC
uiZ52UqcGAjZBdNaodDBidGRNSVya2fKWzSru2UBnYrKxM1cAhFrU090/Lm5XD+D
Y9jYAooIoWBl+0pM5GXERTKM0cnSLxJOEhReDPbezB/KHQE8meaOB0TKwDJsH/BG
ci4wMf81AnyvnkIRVqK7Jn/kMl+PiSp65+xB0ZCWjNC/7i+mLYyZFVR90FYf2G3O
3GE4XiOixmRVXFwlmGggD16dPm1zJNyczzDelsPCwfEqyOsrFlbNSNVd14vyaZXb
nwreBCmcZF101CZLlKtDuoTrThcPy21oMjLTAF+KmjMMBDKq0GzzSx2fOf9CnYRk
jg4ylaC4XLX0VUA+q3psRhky0XH1REGOVsslO4ap2Do15CCImgZQBpasXStqS2Sk
PnUnJP2Yb8/0UTBWFOp3S+IeYhnwU0Onkma/T/fb/lk=
//pragma protect end_data_block
//pragma protect digest_block
xDOX4Y+vYldXcJHkz4ClHJsf7Gs=
//pragma protect end_digest_block
//pragma protect end_protected

  
class svt_amba_system_monitor_configuration extends svt_configuration;

  /** 
    * If set to 1, the system monitor issues an error under the following 
    * conditions:
    * 
    * -# If the AXI/AHB/APB port to which the transaction is to be routed
    * to based on the address map is not specified in the downstream ports
    * connected to the system monitor.
    *
    * -# If for any transaction received on the upstream port the transaction
    *  address does not lie in the specified address range configured for the
    *  AXI/AHB/APB slaves which are configured as downstream ports connected
    *  to the system monitor.
    * . 
    * Default value is set to 0.
    */
  bit flag_err_if_addr_not_in_range_specified_for_downstream_ports = 1'b0;

/** @cond PRIVATE */
  /**
    * Applicable only if the system does not have any master where
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    * Enables the AMBA system monitor to handle posted write
    * transactions. A posted write transaction is one where the interconnect
    * responds to a write transaction without waiting for a response from the
    * slave to which the transaction is finally destined. When this parameter is enabled,
    * the system monitor disables data_integrity_check. This is required
    * because a transaction may not have reached its final destination (slave)
    * when it completes at the master that initiated it. To enable data
    * integrity checking for such transactions, the VIP correlates transactions
    * received at the slaves to transactions initiated by masters based on
    * address and data.  If the VIP is unable to correlate a received slave
    * transaction to a master transaction, VIP will fire
    * master_slave_xact_data_integrity_check. Note that it is legal (though not
    * mandatory) to enable this parameter even if a system does not support
    * posted writes because setting this simply enables the system monitor to
    * correlate downstream transactions to upstream transactions which may be a
    * requirement even in a system with no posted writes. If a system supports
    * posted writes, it is mandatory to set this parameter to 1. Reporting of
    * orphaned transactions is not currently supported. Orphaned transactions
    * are those at the end of the simulation which could not be correlated to
    * any slave transaction, which indicates that some transactions did not
    * make it to final slave destination. 
    */ 
  bit posted_write_xacts_enable = 0;

/** @endcond */

  /** 
    * A back reference to the svt_amba_system_configuration object in which
    * this class is instantiated.
    */
  svt_amba_system_configuration amba_sys_cfg;

  /** 
    * The upstream (source) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB master/slave configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int upstream_system_port_id[];

  /** 
    * The upstream (source) port configurations of the ports connnected to this
    * system monitor. These can be CHI/AXI/AHB RN/master/slave configurations
    */
  rand svt_configuration upstream_port_cfg[];

  /** 
    * The downstream(destination) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB/APB port configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int downstream_system_port_id[];

  /** 
    * The downstream (destination) port configurations of the ports connnected to this
    * system monitor. These are CHI/AXI/AHB SN/slave configurations
    */
  rand svt_configuration downstream_port_cfg[];

  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_monitor_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_monitor_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_monitor_configuration)
    `svt_field_object(                      amba_sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(upstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(upstream_system_port_id, `SVT_NOCOPY)
    `svt_field_array_object(downstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(downstream_system_port_id, `SVT_NOCOPY)
    `svt_field_int(flag_err_if_addr_not_in_range_specified_for_downstream_ports ,   `SVT_DEC | `SVT_ALL_ON)
    `svt_field_int(posted_write_xacts_enable,   `SVT_DEC | `SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_monitor_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_monitor_configuration)
  `vmm_class_factory(svt_amba_system_monitor_configuration)
`endif   
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ygxDR8hoXflvnL+vwlY4iFbxn75ddJYbT+PaMlZG0tmFcPdLjtryNVeY/s0KNeiP
kA7rM4Zep7SDmrdAVTBoVXZRAhHEYwbVvcg25IbQ3Bf2eW8QX4f5fSEgw/q0P1Ik
mEuaJqlpmu0PqBy01dyeRAL9tYQnW8G8Lvkl0g3tr3OeajAOML+ZIw==
//pragma protect end_key_block
//pragma protect digest_block
nQN8r/g2wdFMVNbIGlp1pR4zlO8=
//pragma protect end_digest_block
//pragma protect data_block
wmaYnff6g3hGf1jRe1rLk4wjH0ipdcJiY0xdLk0aP5vSjy1q3cyjo+tJdH1Uya07
s6VvswtDGvTNB1mtXzQFSx+wZIGHK0NaBKg1aC4zITDowqijLNUpGYNZO3cVXmBI
cMCUzRQmlaSqRJnpWHMgnpp03UO+7t9p8X5Q9rduOldWFE2ccRnVz3ggQ5Qm3YIU
Z7YEBBBs0M6lCimTQ3AllPBfZCk+Ri6b7xHP+YJK4bRDDr8u2gwUVv08m3RY+6J0
k7ShhJK9PMtZJgoC63S8Q+xGf6V1uF/3S+0KFRateRjD1zAuykXhR244u78aLzIh
ITZzDtT9EWqi68ov1wcAyO9N6uYS8tigrC+nkT8cy7WHX/7TxMszM+8hPWZ+u+vL
dNG1k3uIMRMlnFlhCfPlpmxV51L3U/dc2ySa0mn9gTM5f2+fOMng1pM3l30LBDFJ
g9qLr59+GyH0rQIppqYNJif6n4/wjEmFNc+UPzR7B7hZnh+JV5XQhJMp+89tGmjp
MYH1ofDFh1QwCwImMbLaqywHpyFHii3vF6FB4DlZAi77oaIjUKYE88GgAkfFAAZg
qAZo00iGA/h5ZxeM39fNoR9bcIQdl63TRSWRbou4iSdHTa93Km1lFe2iqg461cNH
6EH4GVXr02AVKdS2SZm66u01S8Le0FrpeIFTuLX1/BCbZt9hYvnB14n7aW8D9QNM
KPlVm0mE43ZwUZBgHUOk0YdILAnZt13XYZh11jH/78sUMGtLe8wXilQ0Zy+CITTU
oAh7zx3B4MjI8O3TY4x8fSrYD91vQIH7WKMabmmdDkJl8ELE0Ibb5195mzoKdM2i
SQTXSZwd3+Vrwp5N4HfkD5EzcmmKXQP/LOliU1KQArIPdaAJeaW8zruJFX2vnbCt
94rRDlv/FVibb2XJrFVBsBQL7Lw4AgWTiQApZ4kFNSn5XKeIfJn4OVjWJUqf1RF9
UJmHsOJTFWFmZ4UOmHiFdNdhziYV9P2vH5IB2KeIqJdm+FVxtZfHOa9KvKGcBhRY
l7ch6BeGAJFXh4DW1XVnEwNe89n+XFeONIrgN2nhDY0WJ9L98AiiVTu/31vxyCJ5

//pragma protect end_data_block
//pragma protect digest_block
PiYySH9OWhH9E2794UldKIXEQbg=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XSOUqZREiV6qsNv9lt8Q0dwBAgADYJF/Ceihk1kIe8BPEyK6DNdfEgdhfC7WCUJC
BZoph37OgFBnDfGRvLzpO+STYp8czhYKNp8OxI7ONWe7x1vVTKI4f38fWxArwGfH
lqDfJyUyhrxcACXaX1ezd+E8YDV1jj893Oah6JeZ18sWkC/UkZoktQ==
//pragma protect end_key_block
//pragma protect digest_block
9JjECOgwkTL7PQD8064gsp/v9AA=
//pragma protect end_digest_block
//pragma protect data_block
wgygD/iO0D3p5Q9pxefPP9bGATI++2CAVU8CCN2C4kzTsLpmakZX5RuD8uTVUHls
e2eiGZmb3IsdCj3aE6LQ+E132s77zHwVhG6y0mJx6vqhxrUmkRiM9fO4if+FJGg5
BB6AsOYh/PbvxReiqXhg6lDEhmVtBrLIsDWJQpbNkGG4wBe4DGWO+R/1ZNkP3Ova
xrcEB3ty63AJTtGG0TaUVRwdXkxi7q2oma1xiYYsdc8xgnWmklK75joF0Q4V8O2n
clTHU1owQZXmTcDeaFK76FwwCZ7dJ7N6ECHQAb5SI6yrbMfN6M5JCiU9m9RsbObl
ev53CZ3/UyMPkOsXJ1Owi17PZhJlt1pgRpL+LNwKr3rYtU2t1V3vwagIGvPPr39l
Ks4HZ5uAiixUO0KYvxak11Nb4bgqOsxJfAd8WKUpwa2P4sDfC6zKW/35HyIoUAyy
P8+A3mRi2t1/858F0USwOZqqGO0IaZHITRfzgvJjGMtj9nI437CIOBebIHak5m1J
K6vae5NbfaT6m4eHnpR5tIWBeT/sepAxTbHE14/HTaHDiQxHlfUgSvYFh6avO7pW
65jex8nNi6sSd2miLzOXpGUODm92A3Z7IeE4/qAiIG6eVxagmc/kKqHNuvTb1VzX
e+9l0j5RSc8fJJccwEKZEhNs0+gW0x6n0rPB4twLsthgUbhwaj/IW0ozbMV/KFxh
y3rIskcbeeaPAdtyADk/wjpyPMdsZS4pBvY0zun0bBW4ZBZf/y3mMhc1eNGTtdi7
TQqN4FgLcza6QhD+cUXESfGGyfZLxGHXZgadhop2xuEjXlQk9NCvuysxIBRGzx7p
+2oLfRx5x29hqcKu/5/zDOTdgV0EnCjyb24kTS2AieXnrE3PxaKx7iefmFvc6OaO
z6huhGgfjkY5jeHStOqnD5jv1SbGMwHNBR1VrKBYZtsrrWM5E7IkfiNh1Ykh+HOo
CnFDmVj6m3eLA/wMg2v5mYd9ns5VQxeONaVjUzCtWbwDqSTSooHWx9GjLmXzEUXY
rtgl70s3j2pohj6zP4QibJA0xQVjJY7ihp/FwW2W+IT/2eyROR2mnS5HCjDtSnut
eVwklGuRIw30+eJ9gOEgZVtlnW1VzPs+i41V/XHBe2xMBxQZ4rQ/u5wENCLd9MzX
e2580qsxJQpnVsRXyItxsp1gQeshZMBlqgHF6CFs4NSt1+PDXyCACcLiuaodmMDo
Ox2plaRap8ACfyZgfMkDFTLDQoT84VzSO8q07CLKOUsagLM/uOWGHNED8Aqd7vbC
2im3aH9AhQ336aBOFJeyTYH7lH2Je/jNvXQyh/EUm73KIuiWkh4At3+jwI7DSqk6
7y3QRCoMk3Y5zGrYS5Y3SbDbkiQie9PnIbPc2wrYtOCJFGSF2b1+tq5pHUgEmuDE
5J3O9CS2Dc9KadeSyf6kOxDHQYmgsQkfi0s7WgNTdwiw3sJEnNjILYHQ8CZ5H/fD
0Xe5EbQ6jlrYPhKhkFkddB+UNq8SgHmb5ZU+Xs0dfJ6KofC6bWw+NCn5Qd06mzWq
gS+rn9HI55uRfLMyzPc6kf57jNNV1d0nSGRxsLMQfv+CP2FbtkkH2UtjzU151C6a
4xCycbiudi5/TH7rzGClITVBOgzTBypc1b+AUZxJ7MdMuJxV4+2dpO9xAHcwKgIo
/ufJEtDInIIfjFDe+GU7WspS4Dkv7IZvv7ua34rG21vGWr1qrTCWStNCJquq/xFM
ObdHXYEpfhMnMtkUirnBpqMiUocYmPAwuOqZmGQ0+HgslAV0a1n8dkOj0VucmCYY
x3gFXq+UgaZjlRq2nswI+fnodJyNZYPSq8kamg8SgLO8Sz7Ch0okFlvN60Q+IAEY
LfshuU9weEhKIvI2pGJjAKkD+KHmaGpHLoIvKt2mRExVTdZVaNsxXUEq3dScHtLx
CKJXKa2XYewm8T8gT3EQcSZZkHyq2aOvWjKJdmsEaikikuckFob57D0PZ/tZQ7Qy
dvPLwFhFl+100jl3TXuE6ef8XSGVyHjxeuz18ByWpyAqr+gKNznwAGUz+R8usQtd
f58x22ut8dkSdT34F6MyoCg1JPtRaWD28G5vBnrVks6wP5I/OTbGVAEuSjxsPHex
WAlkQ3HQwjoT5lpx13eKR2dchJUCfEEXWOHk9t80qIU3ypF4kK36BCoKERU6Vg7B
83eVBRUKae2qgThmfryJ82u7D0twZ70cqECRiImJbaD+bV3Uo7zCmw2QoP0d6Cpv
7khtCMuu8pGODoqwaTNKSisNf4DhgDSBSl2idRxJXi1KpnHlBT0rNJpitoF67uh3
wmX19I2KO4V2mF3hfpELtNvFWAwVkt2e024hNwOiBHO81SwTcU97yccfBYXwV0zU
EZm6O0FqqlFPBndwtRzAC6CaFoepoH11FLBCXjFAABGO6q1YNVRM+Ox3Vf84hOkS
fU3EgLiDjWSZfuYGCLigNmPCnDncP9h3Mn9tgIQ5hYmiBnH2wSrUKyfdszGXgcy1
+XoPnfxWRYIaYIEkY9GFG7VFbDQxhOYHae+ffqd+NrQghz2BaznFM2KuOUNI9pmi
Osu/4pMwWDjNGuDDgquyjblJENoEmz/Cb2nt/6sinUvWfB5Qzj/fWSF1CVtPvRaL
JqJZYcAlP1SoH0k3AVW0MXZmjB+nUDlcEHUe1Bf57aEZHQGF/WbRnNHafnNPKtMs
goB+adkDWEAv9kWFd9G+9qQAjrYFytbWydfUSTzOr3ueGJmRXjSA98PTOAkOeUkU
0ja10VukhM4vf8N/hij5SQaAcBmQG39hA8drqPhJG3w2yGDlPJXlMzC2ZfB5jiL3
1UMaauWujtwYLhimTlOXLkzKiDWXLUIAduwhCm0PE9oTonCutx23owHBqUNffFNw
JqKOlrbNWIaWSNXobm53douFHZp7eDiL/VWmfyLiWtQeFbPi33sTUm3W1JTWludg
gWAa5M7825uXLR2AfIcGxi1sWErwhdNr4G+FXrYsT/+S+SIzW9q51hUGT8VNafZS
NQH0qt5G0/KB88Lqjiat0YmckkvpEuWE9AnMpcA+eanx2Xuxr14WPN5AHNGvknkh
Dg0TYLtCPR3OE5rim6oRxeH0j3XgtXuCeeBxPSzJ4iRjSImDI3b1YqULzr1I7vwH
3iawIn7/Bl9bd96QNm7c139+9CCneCSLF5e2uCwqiNb2BJGisuwCsEMoGuSbsEf9
Hu/2HCK002Sk9+i6IYWebQ2DGy/lSINVotrg4zjzt7Qox0aJxgofWKaSYCO4UEfO
dVfAuFMpY7cZ9ea7ODMq/XJlk5IC5FPtWgY6/81EjBe++PVD27BOryPunhF8oWoI
eDqYjobdcXbiySNU45+IK804Nc64TPMeG5Xdwp63GzzDJZl8K5tbGVWIZ01h8RU9
HCVQz94pSKQxjtbi8Ux6S1leqc7BdsFWk6UBgz7QLU1U52VSMZzNYGYBFZ4dpIcF
V59FONVXGx4RPjhRzaekFuApWgyHTq6ib3i1fFKNHdi3696hoxrMweiFK49Rb6wH
C0qxU1t5/g21fx83Zdf8jsL3Hdy6g35lgg36rWT6CuYeh5iz6YMCqv4ehLxRDTCk
txoVL1a3X0P3Ov8Z5WVYKBRHYDoZBv0a/ea7rSHN0GGD+aH87MhftoemL7YJAijs
qW5Lb4bL2mhfGbZX7mJY8axn+7nXmhMC1g6BaHN4fyXg8SzLz0tMvfIxYkfqIO12
ebVi2qq3KV6UkjypvjyphuvqQy5iUlvCtwHutFy7rOUcpgW+PWG9c0myCvr+Ik7z
Za9MM2PB6lzEbg0Jf5pGVbQpQMLBiFjjTsFQPd8sx6vIy+OrIHjzW5gINsfh1Bko
dhzlYMMmwgextV/2c+xFpWuCqf6lwLNQ/qFx3qTaBxrTlu+5vYQ4EBM3iLdhVcnK
8uOjgWX3obJs2DCZmaEVAVK9IycZRdK7M534pbdlL507Y1FLbmkk6X8hXa24Z2V5
uDWjfLrCig2ZDYTkYEs9hD4VlSH8MwRvpM6+1LDgOQoHHBOIiSwcHRc+F/M5+eH8
wBEwPoqc0It6zOSidYkwo+9hGmzUdtSyZBgObAOyCxFu06/gx/rFOtgafPVkUE9W
9DBnAgkFQPcDTAc+AHy6861EEtluFlsSIs8IbU/4BPDzkIr5/oPEh6H/i1E1bprE
EOtKVBVjnRTOHl7chvYPNuB5Q2aO+szghqM2LmN7uRu4+lApkTcRXYuDH8FSsdGF
sf/U0/qwCCm+voUiee81gkTQSzxiRsibKw+pBUYIoTW7ZCzIwxrGNeeM/4aCkr4s
IkSSroVDCwLshlvbCU2f7UhWKfcGpDkgP0/418oZw+xyHIt3rauO9Eq7tMaXsxYK
AixV0uEWOYR6I4irV72M1byEk4ehyUlGiB8itPbJbU84X6uC2/ko5DJNodvOe+me
LJLFtGyLrBc9laC0oi4akM70ZVMdVsOrjUqX5PXtCfgv33FoQERngGmeiIWYsiBY
70IC8Rv3mxZsUUDPj9MnEaW4McpPYp1codd6ZUDRL+u5ag7UfOWMAN6stL5vZXZ0
rQX6NBdZL6X11gYXIy4Yg4i0gnEFpDbDu0oUXhRE9SjJhrpxP4iTkR5+Ku39SnfE
GuaHyzIYFU3fm6EulQfS6/cxZ0e2yC0TaQ5n2Jxs2fp7WmQHSV6qRsNEBRwjnENm
uRFoyej+aXgF3IHeflROLPN3+S9cM4NQJZbRN6jF6daNCCQ5eHZAjS8/8g0sbdBL
86qQQTtPl/JKwyBBbCFhrHkZp4kSxhsxTazX3evWuJwq2OuVhjU7H7pyrPUf4+k4
dj+KnHpAWSQq3ehE2OkAKUalbL49tZQEphAIA5B0sVm1m3MOi4hVRGq/yLlLCzbc
tJppdqhSBO6F2at4ouO+8KBGS0AaPpwW+OH/XB3+fY7Cvs/p1gK/wF/XeBXydrBj
XbPlRCm/YeljOxHU1ar9lFxS1eWhqFys/JzeijLcQcXtCfnZR0TrvySSMFLUuzlc
jt2wLv3NHATqePNkMbco4CeSlaOJWCE/ruxI0MOJgGgugrWaRJpzNVNlD3LvI6B4
p7N7hVBPa3zat97TxOzT2O8u25PJ1leVL/DpHx0E6FEXKHq7jqdkjGDgmil19WZv
iWU7hUrVN+U/pPV7/qXnAKaTeYunHW6+BLjeOsTEIhu6b6uOq1WrxIdAsk/KwOMj
rjVmHzE2ppSn7gpfA4dHp/DQr/sdyQAGQoR+ZvWrbyFGcLStIWToWqnABseAlRvc
eMQTX+/gFkYJsBdRklmp//mHFB5pk9ZZ9t7jR6ez29QbmbafeAkIFENlxsm+DfCf
/uY5nM+xmsQtLnsVIutD6B0Gl0YuS3VynfCBbfLK8HjqNvZ6v8H/92Lr9iK2smsV
ssfAouokpgReKo9NDUSt1YZlSAiIaeZMtHzN7PGS3dwh4/D5V8uZlhKi1pSy21kf
wRosOQXO+HL/iQ8WUU0LY8dtQyFgGzlM3Mq6LlJLWsBGMGv45BimIydMgCQepoqk
1kV5HYljRC6R1FkwhCHt+Ia6R4iLdlfjBSNgB19rfSI/QXfj0Ob+2FpMHbH9CM8j
JsLVmXsoLfHiAc1qlx/sLymuLIotDD/vQTaLTCWu4fnvZ0cTs4tSfgIH+L+g/Sj4
jMrDWlGpXBlOIKT7scdTkBIrX4pk68W/bO3uxxhvSK8O30CXY1S5zxY5fIxny6PY
e9F7WNDARn83KepFIqgEqga7E4+vOEYYnLYUGoZpcZrgTCIR7I5md7h2OvanpSIA
dWD5vYjTJ8UEc3PWqHAdCLtZXPN+/2nc8oKfRV2rzVPHzRUj8VFnMJcCxIo5EdYK
vKDBQfrypkoXdB30hxjYEZYKrEf6DzUeWLPIhVMddJzxIE1oF+1rVa5OSTohAutr
d/qR4vMlXYXwTqfpFfYBtY/M84gYXj9RocKsksfL9IIIFnYnptdjlWf2riFYpXSe
xv93zwfI9gqd9ZMj67II0XWHNZ49CtAjLVgRrgMU75owyalVyLPIZaRpCyvkW0Eg
/PES9g/Tez1pq/IOimy52TeyOG7AFCFWYGPF3CD5nAciuy4QpO6IY3c28DOse+ec
ZXFHmxILK+Djqw8xHYvojAqOcXjmSO0mRG0K/Vrr50/ExFdxf9wQRn0LeAwnAyid
R6JW0xYnNQyLReX62FGJ2Qq9FRxTEkVKsavxm/wfbm8UqutC5wspBbXUfq+GaEoh
wHXorWYsTcrd5TOhQTVPJEe7+CyzdQ+0dzjzhk8CDsKUszzU8BfHFA830xWJJdQH
B6oyuZoep44Ok7NiZ2LWbX1SWNJ75zDxBhvwpbpL6tH7eQlImS3fKL1H9DpSXwmR
xaBZVVebTc2bjTh88P006n8CHq+Jw/NG051KDlwsr4pcwwbVoUv52mg5GNBGqaHB
b5QP7UsCRMakCgWUMqsWsK1+4IZjSHcO6jSLvuKmc1SdcAaK3YbgFNeK14TDxadr
iFhqTeAF12fWKpE9/dDkh71Q6ISi4loe5WfxVPDf/zmzQwMfDAjHPYAaZMhCdJ9I
735aRddcsWtJkme/L4vduBBid5cXykzg72DjSG8xclPA1LFc0ItPTOLfVefP+x5M
At2Rkz6ELmoEZs4GL+ZIyW0UQSP1pC9G4S2K5kJsbWVyikdpIEjIg+fGM81TJEul
7vdcqJVIdaHM6HS3lDFHTgElT++EXEOaKHNoKaLfl5afSO0+DpC8J2UXEkZ+OWuA
bjmFgzWG7Yr6lzQ0mM76A9f31so+BljhwnmiE85lgqHJxflDqFIWqld00yMSwmhS
cp3GSB96hvd93RBN2jQq/TxhY36ygZQjvuDGrXPPiyx6/Mcv/dsQJzZDMtFodsLn
FUt8FrAtU5ZPVi57Km1e57iBM/W9xqn8W3jQxBo7EEmFvw05/EfLbQeyLs5w/Oqq
fbWlQUU4UBO2K8+8zadvhcNk5rvPBU6LlHSu+DoAUFfvjp6HtgaghgNisb/nCFq5
uBuJQnVgTa9aDSBpoXjdN3IF+N+Djaq0BY6JrSxGRdFavfXj3Oe+lXkdPW+orFON
2z51Lr9BEy8N12sOh38e/LIxar+2ZOrT2s1p94Lhc/TazWjgGjfuq92v7wH2L0xV
uHHJTdtFaUNZJnavGdo7oX8zbVnNelbTqQhZABZsU3kfagnM5GmeM1KfeZdtCEKL
p/OmyaNirbQFoUR+fX+IbSwl0VCiCIBnelQOq/IkJLPU2i+YiuJuOIhu+EvnFBqt
97rO7e6K1/tD2sxcoQ5pgc5wc70upipkKbgnfmAicS242ka4Nbati0ny8IWSZEmv
b8to8rv4Wl5MqU0YAgC6x1QXGOu/NC2xK/l9LjFKBC0V8uNd0RGGIzx4BewsaTwE
0mPG/PvEB9rUSlG+FSnLm/ed1xP2NrK9Gx3fOSOn1tuulrRz0hGFEDUhSOzbii7F
tqZxgP6xwBmSomAVRvTkwNCcYJtgQZcASAvhvdupErMqG0G0yrvdhvn2yzrgyR/v
PjO4R/Q8cUzWkMhk5NKmmjkBQInUwqTCTmP0Jjcfy7zOcTFldzFbIGPx9MeIHJeJ
ZMefQt6PKRoiIMitCStudTz+D4df//BrsPgnHBcYL47LmZt8xMI3nRKuFZY7geWR
2PZOHDzC0rqMGpb9ibj+XmCC149G+3Zl6IGpOEz/7hPjnAwtCGfYowJCLZ6B2KDp
ewsj3B7FFpj4MuGzxBioHu2QmZgqP8cNg7MBs+bHH/LEilpuSx1T/JeUe2pABRSR
20yAzv0Mi0Y5tBRmEfrrQh7x7PEYd95nHZyQpmRXPc/nbHIKyOqPgHpZEMIopxE9
GIG4hWId68LtvMTDCy99Vt5/xYklnCzHfcOX/KDU3ip3n3gfdm8nGLQPG3WqDPDE
q3wF4STDmsQBYfCaybfc+AzheLNigCpVMkCEClkCOPaR/xwJIr/d+m8pUnOMrf9P
PrMmdVWqWx8TZ5UxB0AVpRkHK+OUtbQRpw+RWeknmHUBXgn9SmMtbbNUwTUowiGe
eUAAZa7vVFZA8EIn8OxRcJnUbxCoRshpOxETiaqEnkIu0YqfygMWDWNA2tXwViC/
Id6M8fs6FyHVAgsWMA3N25AgAZPAo6vCuls+VR2ZGxF0a132SG5GKE6/Z5uBZUqp
vNeM6rMN8zft8wCvZWAhszzDfyqSgWUmDMw0j8j1L8eumNIc+uKmMXRkrmP5yyBn
xl3KNixjzHcP1Pp4VulfkUQyUvu3wLdHamgb6bPctMGIjCV0Ez0kXqatzwlOgX1Q
a1MuSN71/X6jmRfcmjQ6ztMaLI1BrpNB739ZZmz0qL5WWQE7DuXEpOulrxR9VhNF
E3ctbDsFOnjezUaHrPS4t8+hZGJMJmxzGaC5myHYHRNwQ98a4x0N7Qp0enmwgv/B
fCiJjhoEde5cG6J7UcLsMy4NHTMNa149wiJUK1XK0MTPGwPLyw0mCbfwyKbZbSIZ
G9I0bJl3wHgrMEiN3AzTNwQ3978kdhD+weuKkhqT6KHuQ6ZNvDHjSDSM+79KMC6F
fjNCxu+S8laWLCaaQvlGkWuit4tLsqEBmEyA+24l3BrvBCDpeIxg70zoTeyNJ4AA
ddL5mkRZtzwwqV6KexGqpnh8I93nt98ZlNVIDDC1PpK1/XH99LcFuC0IXfVJGo91
gbKodEY1WkztZYoDiLdPD+qoBL8iAcFx5P/t6YcW1U4QzQhdjzPSBsICYEccgQUA
rHgi/IkGXtF4iFI67ya1+9pPoKmX9pDX3g78jYxj7KsEqeuZP2aTqKZeWmI0jsx8
2g5bNpjEtYczWKGFlAPS1CT8EwZBN8kOucEk7RzBpuVTKVD23FljqFt6illD6zqO
YrmwrWTPst5mjSFCCC4HNcMhGhMxfz9E3b08w6cebBuB2Yn2+vWGX7bdS93lAzSk
ijgsA7Bl1ImJlxAW57O4Dsg1Bh00G1DgyYnv0jbjGCON1vpUCJjl85qqnX49Z37a
2FigQJKI4KM4bf38Jas2jqZEghXX9E42/UFs6Hdwdox1eNmA5IJ5AWAQVTrUy6cd
IaGx04mluKkt3feX5/dHV3NrV0h4zCv/m3wVpuu8aYA5M1/+oFklzsvIanbCWoUC
RXWZK2n7+tShIqFBvQABZBYYEufwpTBTSrQMZ6C6IuHqBlsfHrgY9/BinJqtYWvO
WlifHimowGLdF9vvN92a8hvvqAUA3oS5gXppSboQGpmCtUvtY3XIj3f6oXiYqIBm
0NuDTATb0lhe2Fb135dwmstryKPyUh4Cr8iMunoEjihZmpB2A9suLZmXtXunPptT
OetWeMXTqNeNcOVxgPfSQT8edyiJZXTiBBMHWJ3fEkYA7x87H+7N9xSNIlqIlofZ
2pypIUEwIdvNWwxuOfSpo5l4HQfflfp7NF7PGp0ak+e1PlQQ+iuoAuq4wAeC/xEN
G+4t4YP+M1zRZDjRGl4O3jU2nbDFZRvT9NyViUy7harqnhSaMPzq/mjcdPY7UIO9
F6indh1UAULFRJ+Bx9i0Qc7C7k8h1wGaMVT4hIcC8Y3wEk5D8jiPP4O3pMzZ4K+d
9bELwzYPlhMg8Tb7hciZfdjJG9FoUyx33u1rkNy+jwao8Pj0t2cJo9YOoR+9bfqO
bR45fTuk4GO1SPyyWfIfF/TSa3Sd5X6GqcmuwJtoBRwXC78Dtad5sEC6CXl7gz5p
i7jDNssxRpIFocfesq/U1FmJui/EaLJt28+PXRQK0/hanf6UJXqfrgdW5me9Mx2X
xfYcCtbfOuAy2ZV9LEA8yGmIPF1NHJm/83x1+iyE9HWdYpn5xGoqga5ksnP64Y2J
wAX53f9zUKrMwjW2Xu0qE4IfThNH7JdiQUmdnSHg8leaUxDb4eR1CRCToXAtk2RG
hLiHG/LSnvj2sVLuvC53OEOd4yDEqwQrmCKkdTZdHYjpPt9O5Or9HpQfj0gIrEt/
QHy2KYR+7MFFrqAKyyu6m6QcI4UJcL52va/9ntTxBB5EHzYJXRpYE+sAFqEoVNvo
GFjVK+/sQLsUulvOeaMbE2KZ29IRgDAd6E6ofv4U3mxvWJQwEKs8mlcivT9TeM55
G318wtt7QbphZkvtmpJIqL7jFbuRiEcEz4N2ZMrWzQ5O7yhi4blRlR1JhdIUv+5l
pmpZGvgN+GWwW8ZOTt9odS8NyqYpwwrogbtykjCFOf7YyfxLl2c3GrjOyoF3LGiH
aV/xTD7RolWM7wUG2Iw7VaizO1AOkAvowcjKoV90TqdkvLhpgwdiWTrUwlxq/yAh
BDhuc3RmGAcQA0jo3IacLiARwzrvFWvJ0Q4DARRfVlSppx35+TFUOniRVW5E5Hyo
MF1Ib0Z3NSTII8dsBRfoOlq1Q43pbHTCryx6l4vGd3b+JpZBpVA2w1OcVWD95PH/
5aGpq/jsT0DpkmhbbIgVrfef6dmMxRONTrX/Mz6JDBCiIfwNMraPGbnr/nG4HEO5
ZBBb2tekgranhMYvZ0saE49pUzVaBiNRV+sgX1TV8Lav/PDXt82yu2KerbKYy1DG
OQNac462azUP+4D6+WhvRgm98CPTunKTjLzGZPCRYDhRe6B4UHXwP2N8H9DNNgPR
IqU6ecfUIuFu0wmXHiQzVOd7IRZvWTyo8esAqP0bRO1rlLyF6qoxHjvJ4hAFEGbV
vDIx/qS/JsoP5Vm3oiNfUK6+LZmQJPhaXfW4KF43lXb+1DapG0JBRsiF+Ttl1Mwq
ycP8hY+1kpXvHQusMfNtqDQxaT0jDMMMfQSoHwksiuXKh2aZ2njIreLKmLk5nDRf
P3CBJsvU++OhtfShytIJGUwXSQK2x8XQgNoQ4ol9u7Xd+55D+40lJhOrKx2enKmb
qMEZW8+OHwzNZ82IDcmFT5Z9kzgzhedXRVT+S0eDleCAtlgsBSLCxK5mUvzjc6TJ
pIyb0WZ/lxh23dS5Gg4iS+Evdd9Py9BOyNgFLCNWdnscfhECAgyvPfhOsfnp/oW+
Ss+KmceScBmyRIAHOamwOyUxA66UrelDeORFEu5+8Ea9q6K5WeX91hF6bGhKVf2i
sIJZyonzUlpwS4z23pnht/1JgZybrnnaeCdwKvCmHRvz/W0C07kE1L9Tt3z4AdE1
7tIqU9baWiZgcMLUPoulgfmOrRIJMvRKiKqY8CFy4wBp767vhPgOeHwIvc6lpTyK
D8oxHDKzzEqxzH+YDwF7E2ilra867DY7SVPCwcrbuAo097/NlpMQPg4z1++JVasH
LQ1J9hwOor0sRIIDobUv2LsiRJIWvFbQDBfyzfCzNikdLchL/gwhEKvqx8WTttbm
kWPOwlUsO+jhQRkwDs75qIYL3pR43+ncEQihpE4WsxQWMmX9LA8NB/508PndUhe/
hjeH0I9N3uAIqrfnBI9b87WuddZfdOO++2CCjwstUOZPiyQbSbSvjrQFZZOEvD8s
Y0fS6D154fmuzR0EF5/Fs/jgm7KAeLHqCODqwuJQl8cTU5f3pwQP+iErPEbu0kB5
9xU8XO+lh3sWUn0z0L8CJnlwo85wTAuOUFqguRxOg/2YjGaznG79hJ4h1J56bqtr
JKQEiWiiDnk+f6RM5Ak4qxXrOTaNYjx1koX9rR1KCneyfdJfTQ3fcbuJnA2By2Kx
3sSQ7WmkvqSYwKfA4MEwRNkhk5JTU75eDrIQtcUA22msg/5mj5O0XZlEVUCZrGP1
KuEmLpwUOOgiLd/j4UfZ/i3VguIoV3NulnmtRtJqRWzaZaMtVLahyocIC8+pIeeT
WKjgEGXNpSthdJ6He7wR1XImgfwN0lHVzImxoMvH2gJq7Mi9RGHq0Ov5Dfmtgs02
ba8rgSUgB4ewbWY+2xzpDJH/GWhw+UGuOuI8FOyWb0tJR1He+TJLHEhCBdC2XS3C
cMsmEIUu6T2wTzdInmSGwVyW/ec9avos/Wiv54RFjfzoXrO8urjg0jVvaaHifCpE
pY7ZVat471T0AWx47yi+gez2cpt4nxFZiIlnN0pLf8dIqV2awHyNOu8fg5/rkYQy
2rWldN+hmEHQNu4yBxyWdRqRapeOtf2d7L4W3MWqXg1qjV4eFWN5g3CQgAknAUaM
/FCwrvUycC/NtQ/mG68jtFkg1Cv7FXba2hVW2GCS65QIBi+8A2i3RXPrsmCKzPTg
HPyET25nkDaKw7veLLftVCb1YwGP1MoYWJph37fRhnaxgWINTuBF50jl0wbsQUUN
h5trmBdmFzFusGGb25qGiXHSGdc5fsUFXwCebR53WeHwc99Shm2rxnc4AQ02jm6X
5n+6YRNbhle4R6AmB2sDGnmiR0mO0QU70GUdfM+ID9VqZ2lrBsdNr9MKDC+t0EOk
gL8qpjXCt9E0IbxmbGo4ayA0JovLO1MvvYtmtf3b+P8Z9ofWS0qJQNOW3wGk6u5I
K6OclLK9rK4g0uNUWUuukY+7n4+pGBQ+/U97G/LqpVoeYT+q29G9vAAGTSDzPC6Z
Fv7tKQqjhTZpOif7FhzSAoDHp6mb/kmh6ieLqLAwIZ+Zg3F0z7mRlkz0O9Cyfy0D
ngPBjBR2lSgNPTS1+BER/f0F+AcfbIzRWxebNcFX2Lycjfv5lbZ/mreLjbgIEU3w
eaM1eucz7M1lPGf3J02vkGXxyntF0yOfImm6kkg9+C5QlpkYD+zPykYsYlBwjC0K
phZrASftApQglsJesavhBC3H4J56+zAl4kq0OlTGhuctExda6kUQgPeRao3ChIrE
Z+ga6smt/WwIhl/u9F3aCJLrxUQARV7vJfvRDQ1us72tbsFyBprhpp8k8u6UX/3U
GRHynpln6pVjSG5C5ZOYS4wsvbQ/lL7yHp47pAZdMUJzNaLRVih3jCf8rUOq2xJn
ZdlL/cY7tmfLCXzP6FtJKi7FYzH2YbQNVh7AIC5L/Bj7c57TJzQL2a/GF7S993ni
D0RgUGnmkpCk9gSZTMLTUPi9eBQmwtU57uZv8n3kFv0oj0XOAiwQXow6El+KlhOh
+YGcIEwtv8orrW0tOGWBYRA1V82lZ/jls024xNFBi+G3jpaP3/F6PdRt/SGCdZMj
cgL/5Xrh+DvZIIB3/RahhymJQ4emSBua8CRNFWBWfOXPsa7ycCbsvQtJTOugUbYs
7R0i95TRAJtVwS1ObIAvl4q+zuO1itZpelMHOW+ScZZf4SgXqyn+K0IaGF3oxV4P
/0+zLiHnJJx+lj7njJ2bo8W10UbL82U52PdjISykIR3D2JkSamozNYRu5L5k1S8h
Ro+3t2XBEq7gj9pK9sjz3VdVRyqpTb1m7wRA4KbG+GCJfhr93Lu5o9c5XXiqWxbG
8MTYFDVecJHO3oaEPhD0RFXvaS/oMmDUS557UEDDhalNkGVr5ylVcyxxPA5qir2x
6on0p0/MjllriznfAyXsz9a2oogTXZHcNd8Vuu0JdUdj7F2T8ccDirlDqQEWT++8
qNbYubUcertrwKjCexsLo0GxMs+uCPMO+zipxT8+aZXzXo80rzpxiyd1+NbHRpbe
Cx1TVp0pSv/56+t3i46Be5JKyRswTcY9DUQdqsdz8zftpizon+SMIZ4m/WvRf+E5
pNIAfq7LO8d8vK/P+xuAJnTvDfMp9wEiZPAZc4OHvvW3AT6fyLX7FZD26fl0Bd0K
zIn7o03A8+FD/cqO1dZz2PHpT/nrc457PY1AevoXqiVtBSU2ejFqdGU5CiGcoZe+
mNOFI/JZ11/2oMHU1Ji8T9TNgH5TBxwKfOwOlfa8qVw9zcJVRia5iqWghxvGymLU
HMSx1fm9GePQQPsnxjWQDH9IeZeiXl9V2tRqhReWZDMhyPetjbgKMeh6TQUuUoCH
L5gZR9IwgCAbEABBseHQ5x+Sdi7qucMEr77tkyB2fT2jlMmQYA3sC5nEWNJY8JGm
LtoTKYIpNkuXDFfknLfBSdkBhogAj++E+ERAs5aWsrApwHTq4OnfI7MoiYb8BlpS
ZMCcanN0DjMiu/DHwt3PjUgKMApoBS+KT+GWKwm5sLaTXF1b6dJdEIzas6pXrsJz
5qcrzbJPLbimLof8Ve+ITwW5fI6FYbMIyM+KL0IPOIfj9JoMQAmCgR80OPqkfYc8
ZOpAkI79GnDytt8e0IQm5WtS8tTZb70bXct+3dUEEmqYjmh4TkwclJuzj/rEeO5u
jId/6HSm64q8+QlUZz0ZgE61axuwRVyyKGHr3Vh1btVEYIN8pk/SLZczcmG1F3X1
ZYYIxtnljwgbxKZznPsI6abVyCJ6JCZQTF9Qt8rNmr7ueUQvPLXRNnebRgIekdT7
hqRY78ugK9rnZl+X/nU1N2spTReuTrCCrUFnvQj3L54WufHkIsLg/5/4+mAx61IZ
IqqwW4esHleoJ8qPLdcC/Q+N+uZncTg3KJPmkjNrSgw1C8oKyTr74+sYDfblq6xi
Lbx8YJLlkyW2QaRd5w1/RaQj6lxqv4r+l+NVcOwnhzmNrPni6JG3j5kJNKcMdnpP
p+xrqTTotLbTU8QoyWR/XyT6usWvEMDzev8wsk71Hc8wzUrggVIIF+PMzVlA2Gfc
kmjTJBLM8ZO2EMBWRbHRWtvgQGSUtWhjCnOXCQQ8RluWNQtabXdMF4mwlrC5DvVX
E86UqwHZqbKKh3wiXdbdrmyy1dCi+3dO15/KTyySCopEEK//i5oArg2SpUgqu/MA
WbI4pqY3Yxn2DTXylmUJ7VUSrt5DuiNarbRYdNQMWfIVHZZ0Xi03PtlQrFBpk3qE
seIkHbcREtzNyxVf2GsUA63jmdKI79dcdk2tOB869AH6xE3LONpoh2Vlnu+hhMtn
M/WE4dBsY+Y4O74AfNPpGoUxzyJbB6NoOcbkunDtcEbBehgOnuGsRHX7guynDWDZ
hzGPnSkVDcIpOS5S7/fkIb6m8rOUejUmZfMNfr5pFbOeIp+NjF+GTLMDJLC330cR
7GeyiO3X4l9tFte37TgYDTdbqNLsiB9LILfySuP2IWTLDq2mZ+m1DzAwpGeCsfjw
jUYikqxEEQiU4SkYATTm6brXYejk1h+GsUJRFFpLhuwuOSQHHQiMFeirwstRV7B2
RSEuEsj13hnsBh3zpnDNgf4WR7aUEHcc+NY74gUnbKBAK4PSJ2Ji2nyvE2YAraFP
5QhbIa6NP7kCbAIU7J27ClghU3sUZlZls1Ba6DF3R2naJx594eoS0EQ0Rk5Q3+mZ
W1UFLrlG3XozDaG338LUAUBW4jl96TwT4RSu9Ax2+2wfvq3JdxHynp36Cs4c7nbR
VuNutWx1eAY5yXk3ufSKkubTWRWySnVQ1XyAg291xKEbYpzqUGZ/+hpl5p1X6fYD
DciXEO/rso1zndZA/8ZjOCVy+BmIK67QqK+9yiuS2CmXG3MB8a645PV4XdBmaV+o
fwdHTxCRfwPR2YdhQUcL0VJ8yurh+vuum2qd1qzqRWDBM8EVqA0epeYpohkElE74
8AEQwa4XQTdCuACgGIMJ6TLUKOL6KqzA52sRyZvFwEK8JvjLJNIYE7P+0DqkptGW
p1qk7mW0clvaEVK9pPVxNwnb6K8z4yvExNd29xtgFkqqT5di3Mc4WxrQC46VYuhB
GWjwj7x60JLAnkkei2OUXsQB3hfIuTPxZ0gByFu0rLBVATpcYauEEeAwDABQ6z59
Mgua/lGe/MB0Ps6J95XrujN3pah4fDfx4Tv8758JH1Q8Kc3YJMJ+ruNx2kPwSVCK
phcjjG699+aVGbdUgA0pX+8smGGOCIXHT80w4SttaLLMyDbRm9aM5CGHbYmfxnUk
BYMVfEnCr6Cz6mhZ76qj6QPgswOCJx05Ps68b1ZG5LhbYvez5O0Gxfw04xNb43CB
BLrI6v+fyy9rvkXT/lZwaDf7JhryGvmIYS02K8syIuIB6zG3jNRzBcwxmg0H5+Bs
xlbXCCR9vm5MdeZEIQHn25o/QHTTXsdmWEOmXFKosd87iQjwzvXIxGHsOXFiObHd
Sz14qEujfchMwAT7O4ulSkwU0Ddt7DqnMPqTE/n9AJ3G6XGyrfXVVXbzvDAog9PN
IyK9D0/H7V9pOcl787E7VYJJrKXMWhxG+Gt+qeg66Gaoc+4k57SqAsfXfWG9MbLz
a5oao9RaVWwDtYUDu/5soeSnzzOKFf/Ozb1iMa3F0+cX57PF0T6rihCcjoqsZkG2
uxBqJ1yRJwIgN2PnVRzGAfHbNI1AwrH/u5cCggph2SfVRPXCzkMEw3t64wCKo9/U
KnrhGzDmwsUJ9SnjwHrovPRJuOS/4W3lZEdPcMfVXwKDrpcWBy1OEtbteloOW6NP
W/SMbXSxtUzX4o4oy3qJQ5qybfVcWS55aiKeBgslbkKeZX1eHsSP8Viw7rro0SH5
Q/Pgo0uWGF6NjBFShItgdO+NTQU066EnAhsGGkToCJVtOV0IR24AEjmQRDfRWgF7
k9Zx5wed6nzazjyhl5sMO2nqcElxzQFcAd09ZuiQv0I7DYgyEeAvo5d//IBryabR
VCaVo3QdnsU63drazg5DCT0dIKpj2Jami5/1ZT7tUu0Frfow/mqYmZ8j+tQafSNL
4I98fXnWqs7zZvMt5oMl1YpXVsjqcsbPAkPkPsA91OVtWwzdjoSthucl4n4XHS0m
N2vBbCjajJeMaacjtmCyREI13z8SqquolefUwtxrIktCXYGUl747e072XtZCn7+g
ECdtuq8UdEv38fNG9J4IHNtwWT57JTr7DS+YPWDvNGfGFhue4DQaTiQMmHNc7rWA
M++73HsYAz9pMmCvKCSE5pwLjpHzUAkImoTjjhxbAdwzyu/Lo9GkphU9YT7c1WVE
fMT69ncyIxz8O3vQSjpbOr+qpP+kJauZBHkpT7BgmFCs4BcHzNFvPO1zRVhs6zL5
BO2B/8q0avNpPSf0Uwamc1Bsaqn3KmwMjQAb/l9dMllvrt5gannhGYsZ14qchi2C
3PMRHdoB+45zthHAgi0Jo0s6Rz8SNsmo821FRH5PP9l3AAACcjl1byrc0+aJBh+K
r4b48mTp7W3SJWRHPSoqz38vZhihO70BeTL7urQdQzaDVwVut4JY3JgXYOfD2Gsw
dDIBb2Y08E0TYe+EZwOQq1mLrlkU5M3pxdKOqv/3Tr1RQ4MGrvBypNs6HtdGVjVs
Ol0eLI17waBMITWlM8feNG/7rbQmvfBSOwYRE2I5VxN1LyvO50MXnWyQm1M/t4jp
Yw3biFklqbg18465u0wXWLqQ8GVHAB/vJnA8pl7sEScVW6ri4DH7ZxHx4MXkExQr
TYwVm3aE86lwD+1I3OOkWIvQbIQ0OO7w3o4nB4z0mrnmPqVHpBD8i8+BtuSpVgGS
EHFS5cu1+LQm7cu+ezURmDHNtkVWl+csgR1l7cEV+HGyH4dQIqiJJ6+yOSXa/PlJ
0t1BWPnJheLdJH240IJ/sEzCO/SAKdrUqbBORJVp5Ja4zKgpb5opHUW+kD14PzPu
UEn5ZFU299N9ooPrjgQOV8zmgErHNqEZEV6myvo/sITvcNpVagPwdxskJ+ZEgF0t
MpchyF8OI1IcwHV7ygNtB0qCjbKJM+gE5qP6rtwkG301SrkJwYOXJrxoWM+erTTc
qe74WHs5hXMXFJs3mN+etYruNIU3s0ECTTg72M3jhqimvTVl3DDkdRWizvZ5D/u8
e2SDH8TWE4h/QOG5F3Rzd9KTVjXC+JZpJX9VGDGVUxzV0OambV82/GpMOVdzK5t9
+tJjzoZ2kyBCbA4rV/M6bILpOTHX804WrAcFmIbOE5QHDCQrxlsTWAshhqx3moWl
vhppA5aEj0umdVfWKDf0jQM7KmDA0VXzyoB+P1R6SP6Vcx/OdwvqStkXVLic+QLB
tpTjQTKjYrY15Ds91SKot8rabMIW6UdoUVJfMu+b/FeCX6fjEB4P0r3xfiJ5o2Ol
hQZfkPjFedZkLmVphePJSFVJ2brT8G2D8UBNiSsMb8jEiXPtkfpzcLY4T+V87h30
P/7vWUPLnISLgZQ9V4/WfprrYZmWjb2IJShG6y9QxwdU60kv477N/LhFKnZCRsaC
kICGeHWdWie2z5pr0iOw40UB4cz1P1wQ2ONik53QOSXHhxZVWBYIUz1sQ0cRXYYz
xlcz49xvPN0+/zs0qXH/QkTEGcsoLrT9P/lJXEsTqFSrx0HWeMgGcdJqbd2suqL3
/RW4TyvDVvFt/OIwxpxM3ezTq5+CySKTbky0umSvDQt/QZ2/UxYtOYoo6MNUMD+A
TuAlDtaAfP71g6ODFaWudsOF9cxjcY7UFAdtcWBkNE1L9vENp/HIbhaMNwoL2iKf
OHa8BI4i9lz55nsNP0B1S6EKR+cNL6JY7DpCNFdT2ZG6BrLQhuIpAtqROXSohioQ
TktX345pszSWiMDkddfVG6HUrG2ajFVoFddUmQX5JdL13+RT9GRThwGy6nJTSWyk
Y7mo7EQrMiQcKsYbrM6ccmKye+Kya5xvLDlDCD20AgLUy4sklsY6yolRklZZzF4j
yXYinQ4achVzQfXlxGpR3v4+zcIGghz65JUqZDu+WM0WGvap/s4tG0roC8hFzIEu
Q5FPE4ObLH1CFlLqPdX0iHpg3yWchE6lfSIrXu55Dwo6NhS7ZN+YPUSWhqI4Lt2m
5HnT/vsm//fAfaY9ZwO/LnTCVKr3CWmwQcbqAKQdfWdVlWusCK/udbhOQedLP5Cr
WBVJYSk0cs9aFhE+7nFBJWV46cxvi43Nzml5uS0wcluQVB3B3YLdo6988D618CWC
BYtZ6dJAfM4tAf8060s6Uk9vfmkejrJNfXRSZZxFVPO+dtVmBfRLrp2+UpaDcNz6
OHf+tyC2x2q5Q9tz+yGfwNA/UsyQwOuSUoCE6mXWxWPNrWNyyMARF5VMDV5/k5KQ
+HHKXpQ2GVAEdWnBk4NbfPg2Rp12ISRnjMEfhbNifp+ZY4BCrcat4U9NEb6/Y94V
s5zoRs7lGHhz+quENIQ/a8BkHUpV4bHjrl4SSj8+9W9j3rJi2xQQiIp6dYKWavOp
dp99GD0srAAIECZ5gaNEgwyxwVfK96fmrXGVlbGu2UzLAodRbTI7lkkLy/42SiCH
BGQf7PfZaySPqOp4Omuvti06qexYMPC3WjJISLObyIDumItVw8Gh/xk1wqupYJ/+
R7VnFdkwrKkcSGfugYIs3kdwUol0WdSs41+MBddRIQRVDwP0v2enKG/sOjLkm6XT
ufH0SZt9ur8ZXIeTPvWMRQP+b2U7RpIBSjEvZnb0LDkloQxD2DTRiv4fm/fWtGlt
udOytc7/nN49qzT8VOPYIAJrGOA2IxJRk9/DgIO2PsSusNCpN10dLUoJ+wWuM4es
nY/5Z6osJ2XUtl82YJsPg+EvEK1TYhQjLz2HDZHtK1gHHnuhReb3Sg4bhYvXTOYj
DobUqSn3jQ8jlB5boTgBdVJj7IOwso3Wmj1t6C9aJj0Ha4F1Z9/Bdp1oNE7JIs06
inX3TPVDrnl9wy//nC4dgiv52jOus6E8ncirf+5PJP8Oky+475q+you3upbZtWlt
DQGcfUlbuITdcdjWxHkHof21oJQzyA0F1Zec59zJCd3UW0eMBHSf8OLlwlYGZsRu
sycuaz+TaxiqkCWFKBzhA2+yVMkPEJ8/LJ11QkBtXCxKCjDRSdKT0KoBaC1MS9Dj
c66wKdlUtiq1ASojUUGMERLw2ZkOcGm/zbiXE6CNVf6YPHg9DqjjPs+YOLmwJpY+
Epl+l26vguqsE8wO32p/q1Rnk7p6pTirFKK30yvHsclnYHZtEKytgPfxWlzrf5PH
AHi+P+u5xPJTPzVAWKAfR6EOLxmx8KptXB7SrYD8Zj+xQbaKxUkaXQ2ZjyEFhZbK
vn54pxQPgovoSTpco6PNUlkgjWWOw40BCT3N+nPWOI7vCtU6HZjp2nfzXwa+6S3X
UcQd4Y4oe9LUkDlmZRRa//JPXj+7hYjXPx14r8wATaDRi/gxsIe6LQxyCAjRj0D/
O9A7kJ1u2p+8I4AXcIvijKizGbIzkKqRkc3y3Ev6Wp6IfXJ8jnpVUjFEGfYjE9Oc
stngav5ayaax+uRtZLsRrsX9SK9dYflfb9uhx3L06iMtF+jbk99T9SsZOBOWOhdP
CP6BYJLFRYa6jYiNdcbOKINYI/tyMWwmwdcWEcalWsQqLZpzN60hJEnNdUAz9lJR
4hH8iRE1gZsnK+gdrQcYFNTRunqHiiCk3K4IM/4tiEkXdu94jlY96hK9dqeD9zcJ
VRvK4CCS/hHFaFmhppebQO86V4uq2av8k6dMCAj8UCQVGhwBVDENgncbJ0IBA5as
1MhOfbQiPejZyHNZWQFN5miTChBZ/7mmvzSw8ArifQrNJcCC6n76yE3taSyb689n
Az+R4REftx02Let5TFvc86FD25U43GqWVF3NTlgox2TV1b8pSZyEKku6Ql/22A3/
Uz/fvoVb6+ijnHmrVQg273Q3beu6H49YoIbu6W32bEqtnIttG9LpTIG0HahQ4plo
MDKor5jOX+tbykFKH83r94CMJUSjvUHMucFpPvtN7YaJWdXAiPXB/4zitghtdiBU
WkhcBJiY02kUQy34mqxycKnSDhayiU2wDpIys9nI//vljY0oT4q8sixTzsQFg5IS
wJhKD0RpsZlilLCVtbbWB6Qu9WYTXPMXMV9HG3hfst+1th4WmTtGRXdzbVjrAtre
s5Dp60rqWwccdQNYHQ53QIwkAR3T256r2IM1P4ptacbROnX+jatkMK1nEz6XmWAk
QPMP2U7wOiKwjZLyk27XuHl9IO3nFEMb3DtcfTEs95Pk2yM7GD4jFfcarGV6emjl
qZEdUkdusxM+OxUKZkRJ+BBxov1JGIf3Uf7jVtUuWS610fvgXP7G2smOmRTQG644
SvTIyq8PxPk9uJ8gf64rnFOAT3uwyufdQCqCmwzVA1COkIxIjzp0v5avugtyp5Mg
FB9S9+WBKqTsjX+coLPkuFfn7HL5VcEUBCiRSwWD+KH55h38G7alZQGHqqVOrt5A
MwPZ5HZddRSw2RIrDCq4G8wB6puPDHPrSz+ERHeRHaa8AmKmuFb33Zo6hnIUBOrS
fh9TQfViG8NKH6jzrrd3hoTWCIPqldj2AcEfQ6NBnIg6YK87BS5UATUx9GR7o0bt
S2ZYMVoI3Tzsml8woBDdsEjx43vAmIs6pxUKiOFVgP51qs4uHxe0SppeT/BHkpG0
KFrMuw7btJqxqmqxY8qs7DyqbVr+MOfW4zCMuYoDc0Fq0Pi8uFhkUBZ88hApzVG4
WUoIxFPzyZJwsOs7f5RONAOg+5wQT9REqvZayZyfux4OYxYjKqoAOjEess37SdwZ
XkvJtsA69TMJQ6j+iZcERsWs1ssJLmCvt2dci8xkva+OKYGTHyfgOp0MU1e+A2Zv
Dk3LBBcBAuTKxdAyZauPy2yJWkyNHbwuDa6SaGGl/mVYbAdCKMeZO3en32AxKnmK
cFIR3kQrWQePks50M5XYvgEZlYX133ejS96xQ5U/P8JMF8fM1Ac5wHuNHGMbIl88
IHl7UsMe8tSshb6emTfeSzYNWGDfwvvaj7sNKRWGJcb386T+oG7Picr4sRShWnA9
l7Nnjz/53N/3q1vkmLfN2Xo0jNN/EaSlXksVKhUx+TlQbRWIrLLjuIfUc/ddu0/4
0+eopnwERYDd5Ow/HQ4sLrtOyvo3wtDras6ma+oUGK0e/gmkwIFt4IN8wTNdtigj
AD95N6s3OhdLFLgbGFIFqWlxtUtSq0UYa3apYch9QJwAGKf/tQMFbLAmwiXmtcj0
c7zdnIDKtjaxx7mcrjGIBezb90TbQOemDcDAu6HywNrf/ShkBpNXWBQxcUMsFFAV
8WeUm1aFktnB+MUCTUCRkUUeDlDQQ5QIyYfBxIu4ei/YUa/F0Dkmt55B1Jz5pA6g
1rG1aKZLDU5zn/UYMHVWQ5Lf7+o0lJBmw3K9GvwH8dpRRQeKmCrkpSP+2E+vfw0M
+Dx0s5g8Bbm5BQxiFhT/Bg2GbP7zX4jSNK50xP0BEUl4CXXmkKzt27d7MFsnIvqT
MQKEH0PcvCNBLo91dZdZz3uFEhRrcB5jBgkIUxlXGYSYzB6IjVtWXvlAWqw0vy9I
kUt0Qb+wXcZdnn4NJvAuJt+/bN8qEjQQrwv8qW/umaTBvNXAVVkcW0HuQHEA4j5l
d25mu6nZ8OaxC3dt43ZsfIJ+MB6yExgLgtcdxbKpbrCBucS82t2N91Gb1ie8QOkO
xtkdMzfyDvc2TQJqraJ+rMPssuWs9nB59z+AT2J4g7PnrJoiArgKswOHJpY89rck
22rAEd7L8CLIffE/CzL98BJJ+JpBmAcFQMzgw/irZWGIjsy9Fy2dXKzpWmAb0uza
kmm2348tFWghgTnozTjJDTtLu8nNPOssQAh5y6v9BhOEFPhH7k4veuR/pTF6J3gW
Pxt05B6yt+gKyWYuoAVpsfWDKZnLWZPofqA6oWTIHQyRQAUWqkpKF2ImPKzrOY37
tO8IfN7vkJHRFcedZcBngEuYqp437c/51wRt9p0M2QZOUJzk9+Y82yae7+dljTsC
rnwNq6pgtZmGeyE+URV6J2BJLjSgbiezGCKLADu5yCw5KwJhwlVNz2VjFiNgQ0vR
OWvkWDn2VdyQpAE53FAx905OMJmYtqIWBb6kzV8KWKYKQaE4TaY+306etrcgP1Wl
UHU4aj8seAlsxJZXdgoDYwFB0I8VVJlodOIDhccyBqtRdcR7NJVnINoayu7QSuJi
BKkccR8pd/FA0o/GkYuiYoleCtba9kabWFibH6z1OEv+dENiYV/aYeJUi0VgFyeh
FrCMRfDPgw4qdUv0KcTGgzwbJoEG2bB3K9Uvhp6xPYP4bQKY1oG5SCZXCZU1wsSG
h9lNVRVWphT5ecaGwrWKr0h0COvDh2b5Wn4WOZ1uuV2tkEHxUdTa2wMcrXxxFijk
sVLdro8CNPWxlOfaOtvqaLHF8HJg74Le3jRz6FxWekZ08r9tybbTXdvddwO9G3Ng
s9/ItxI6rK4RCqQvLAPzH3ZVgG3jJTD3M2Cl6Zclm97NFiJbCAm2s3JUQVErquNy
xkgfY7Lk8AxVDGi+Dl4tMj2IMGIllTAHxgy7SzZoI2ApJEc0o3E4Tm3lZwqPOc07
0aRlsl0Y47jJDYDsRcbsLvu8s4H64aLynw6aIzNItMh7JKu4W+LhgJ6F2uI4v8SS
YeRRo44eqwitQ26t89aOtk9I3EknSbimhk6mVZQPuvM4Cq6V0tfqEOneDn6TzYsR
wXWz/k4dyKIjsZX8TcffInhPdlvHhS1NDcRVbkG9sDYcVCSxBw6ccMHXIRkI0Je4
UM63G0ZMQFYGuZkp21TpWdoFUOGO4Zw4Gano/jLvVkc7VpYmPMqnOgQnsFBteHZx
dp2EqjKdx+Jcnwk8Pbd6DflCDLiMNLBq562DnjcRSTfixHF2Gil3BOxewuZeoNbn
Ha84wd3cqIHumXB8rtCySUz53dKcmagka5/9eyds9apwLOroyQqyXlkDBJxh/zbc
CWW8f9/T0sPdCDzRFgtOa3mjc7k7Sg0wlUZx0AFPlYgzlNqzl85WeD/kSfydhD5x
v8W5y13yZse9bUZ9d/+0Ap7Z8OUiXoHALOrM3Z4VuUZrhNi7+asdTSX3MjmUnJnB
uZ7WvwXaL5wgJw+obMjJ51OZAJXIn1S2GbVCQS3o1Og/UJYgNIShfLxAZ6sdaIL/
Ob3CZJc3NArnp+0jqUXlpr00TGlND58U8fcEzqpKZpffL7gvJ7Dy/vqXXCNbsNdM
OB26ccgznGDMLoRig5spSC5zg1tncL+c1eZstKBp+NVYi8wvvmcc0MjmdHav6hQz
3fKCiu0Ry7W1UgE1snlc6xoBBKFCHbWyiJnj54vZKpyfvoT7yPL45AJfQiuStNlN
bw8cb/6gqQQFCPqWbeqsGnu81KryYEloLCD3XzIRgAXpL/pYoU69uIkWpvEVeP0N
j0GF72w4y0pKJr7g4insPT1LG3bE+M12ReZUCGXbwlWwTIrvraLX/JO4tigNly5v
TVKSBvDNEAM2YTSjgtAFEyckh4gQH5/CDPqcSAiH9ckJ13VZwQXlHCcDV0ltwk5/
LmCu5NJEEv8X5RGzJ0QT3DG0hFuROlni3YQcBQm5BUvbTgL1r0J7uZeS1wu+/Tah
lswVtLQYS6bddcAzEmLBnB6piuQzn3c/B/llu3uWLJoOGMJ2JtiTsMtMlQE2dxf9
1NgXfGwCsJrp7IXeGgelgidsuGa3ETdrkB8Fat8BCmsSooKVpqx2645CoL4w1C6P
yrgTDWUq1EFMlK48j2JjDSU9PNj/an1f7UPlYO7BS26rMGLbHZYDIVG/0emZBtQ6
IitP/lusylinYqdDqYabaAKVElwPzbulRmY0q1/DKYUhI9Qikhit4vQH24BdVNUk
P+FOjuBpeItmVHu6wVNHQHtqsPbYEeL7kFVRGCG04/HX9x56Gu7wtdTEuKNUHJhA
NSM+WeqmQgGy/bq7Okfkf8A8iyVoFkvc0TxnZWLaW/uc/wvIgivs0SFoyPw6I6f0
hiewnOPLsVWzH9hkfWbwtu1TqJl1+3uLx+/3Gq81DFPoDB21KCr0dgOG717/g+lR
/JBuINaXvpEMPTuSNGHyQtKjJMUbvmzTBcZQp43+ivIsVL++upgH+TlivmMh10ib
SDlxxuBfEwVlx9jX5aj+0S5GSj8kTKL6Myo8VhnfSqFi4P9aqWtOF6eMMG9BNlkK
U8Ukkm4hPn8GH4UpV0cHohC271Ox1hB68rZ9sONKKAYqd7XDIDj+lcCcG0Rr5Rmf
kH6sS8cUsnrFG10ZsXaNgf4i/xmJdAYXdqy/y6JzugpARqc4/cBcYjYQlTHd4uYn
17LCLGRf+/+ONFeMhjDsOZkWZcY1ruicyrVXn1ETVYy2m85aNaIbTsg28JoGYc6O
Opy3CxWQBm7GATpBOBL4/umLQZTHQ6gvRkZXuCMRn1MMU/42vfOdBhsECBr86uyU
ga6LYa7K3CrsiPSTpogdhvvuMSFHrQKC0HwQww5/tcH0mUipIaF7EIAulyeeJQW5
x9r4NzyGYIFzpBiaRJKQlkm582FsJ68TdWIEodKu6BQOp8jGj07EKRFMaLrZTH91
+2p4ouvyzm1E80k9HQyJnjJOoeCrHVLpR9KIwC0iJzXCqRWhyVv9dEElCuY7mJXc
j6/lATcIms4ocXI10KztaUk0N/b1GUoJuvw+1ZGYe2YmDGpwkisromG0Ofn5URuc
ZcN7Ap21LwXoDCovgTOA7MnZuH+6EfomStRjv205DEpyq/eT1uVzvT21Q9gUrqpY
CB5QNKRNBm1oIA4rqolmvZjvLlVIrazw144jCKaW6v0DLVZmm/uXQZV1HsjlfibV
PXGzhXsbPs/su/f1uUyz9f7Qkpx+AVj4MByBaManC8+gOvI+YPD8Uuz42ZePne1d
mtwxOe5Z7kBsvTXfC+/LQ/dRdJ7KyPL8dVzWYYa4dPPpPbGk/DsKoL+dVJN+0sFK
z2dlDODWpzl8IZlElISUcSe1CJi2y+xuPsLAfsSZOxv9ebDaLcwFUANLXW8ZT92U
ZIIdnWfrSerlaT8bzXZbIh9YJl8M02YJE9nlkwlddCRUWTjiFDOIBmsnT8MdGNz5
IOquJGzjrO4PjJvepZuw7LQUQd+Z4gbQHMcvRtKXhsaABpWfTIxDfMmsSIlZlTT5
uRL2vCBzLg6f11iA2j2GgURma27Ip+WyW/zcxDa+xwlqedrmza5fUBoc42wS2U8X
m22EfKwQ1CqfV+HJ/ufH76jmypEsmpICByAXRNPPyNLplg1TfTCXLQ3EPtW2bacq
w3Njwi/7XLwjvsyUf3XR65M9VRkwwXFZMItziYBeYmXsoFEgXF+bNacZ3x7agrSl
nrB8vATS2YxZnBRyG0pF5Gt7vlWScnFTh8TfBG3qsRw0i/e0o8R/qMA9tHxHV88K
RLD3mIUX78/z58cQv75hRU3RYNLhE3mjUwzolWQYR9Z0vT8jqb0cSw4q747yrxqt
m2v2QtgukCEHvsQ2RRXAYHcSG0sHrP1j1Um3A8432fdw9k50z4zZrBRjQaYVenLQ
aIhYCwyCFJvf2efITCgTDJyx51dxYLJP4vcqOcQoxyzXJvQcLmKHBXSaW19jKGHV
EOAWvGPu4jTakm9MriDMgcQRzPBQyq9wNFugHnthtjyiuUEU83izM1SvJrCFqAsU
u0VRQT9wfcsbserHfkDJH0KOd2kbQpAYuYyPfyUWX3/PlKSLxDYzLGyyLhORUq83
TZJdWHTL6hWhTSCOo8xe9QPCYBiS94ip2/zrtuPN3ArWWdAj+o1ksqSUU0rJlNrH
O4lGCyCY4oNBeHHJduqxa9TiRs4bmi5xHtcnJeF2sl9nDEd+HtPmuAohMQ3sCwxr
abZqR1m9RT8ltIS/7vN3nEqxh63Z2a+8odW8uaKdFZ5KyhggRUMEQXcOWW21ZZiK
mMpCWUgoJG8vzcT5+Rkg4LIl0jwKU95uVlq5xfq/b2hUr2oEq4KAKrASFXkg9Q6G
Sg8T6jhDee/jJOgaTRR3Hg4IwP2s7AXUFQqykKc+XCguSbn4j8dgp5OKtrbhSAbH
B9p95hR/T/n9k5dljmBrwHgV5qzFGK8/TEBh1Jb039xCZlnXTIU2EBepUkDV/6bw
NlaKOWqCYEJUD4C7w/KrIeI5GU9nZgXGeoSf+cKG3JnqOoEADrP2nRjImlXDGBRT
5ER+YwqFz9rtsD/gtl86RDz/omQRHMXo+Yt0EI1roKBTfQP6MEcm21ihUXnd4xS2
+1QqLLNgGDR/xjDoIQd4+sWeYc6Nudot9ov08cKHq8Yxt1krTKOzIB7v2PSAzs5M
o1vZCC1qxlDPLBD5T8b+n2uOYuijSlK1glATAUkzHFyRNA6yv6ttFhXWj3H+E+n7
pJJ1yxVtiziojIEv33b2VLRloXLp6Kpmaj3S7jKdlHv3EP2YIxFawKuudgllzzPt
x1hioLuVvgS2k2CaT0Maf5JqfpHuPuwPy3FhsFzDvywN6HEVw2//UKArXainua3q
ck2RGHRFM5keovHzyI8V+A5zO4+KkHyyesfLdwUIFsRoDZdI5zHByb+duNA0x2Jk
7JPyN7ESGebOUCanBRYROgTRp7wCEN5jQNjcItKES6/2L2746PR170FOsQoQuHYY
CUJMcIGRiJUlCmCZk978JHUv0ww3zngnVJmeaMj+mB/oPbAZ2vCOnKdVhGLPM0So
ZriYq6V7U8otVNZwWNbI0kGruP8CvKcWGkjcKbNCExrUIkQOQ/tQQnbaOApWiu0A
08MHuhRt17dIf7jkINTlEx8jHVJRLo7NiGA5+CvD9PsF2Ftu+Xnt9lKZH+9Q73Lw
UVCH3S4Rz2eGIKY55i2B1qamwDNY2as0tfpKL0O1FQm2xbj0huWkdEHcipSbqPSX
z5biV7uuPAsSctQQyugDdm3WFC0HQ3MCSNUrHHroJWs7fa4aWfgZ7T/wC2aB+LAq
DbRI4VfmJeFsDweCyxYRHDgnftHzLNgk9Iax/0Yc52MAzz10Rel7OMGkdljPwVJA
LZC8zD6JLE45xrpWinhJx5deAInKvw+GzczIf7scFRfAKTGf9XAynetibVDNTonQ
J8BEBqKHce0dFDl2B4QSELQFD0B8KdWN1ZezBMIpnbuv9YLbLV7svAD6GjJKgXes
ErW90/uxczyG8aADYAKC8Q5hxPnP1QHKIOmbdjmHaQO1U63mPrz+ZT4x4KprkM7m
hJK4ZZ263MzF808zZRtyNmKjXCMw7jBB9Uo9A7+JBOVVi0BYpSXYu0i1K+3xdWFF
poC5yk8oZyO/tLwBCqmJehvEprA5Gwq82lhD4yyh99QPYpvOtdsp9uYzWo5UlLMZ
NSpTYn3t2c8T/Mx29WpX1gwFORhbO6sMC1BzU8v7ackBamD9j6nc8ZiCP+8e1oYI
nShAXJlZ3v31VP/sVSte286lII4SXy8T7LolwblfA23TFClHb6G8mXD2b1PCkzch
PdHP7GXGTcCaNVSULPbYeG4uOGGqqbUMdSkrNIFQs+Eb/vuRJWY2z+4o/bHT6LQ5
g1Ru0SmNDLRKo304zA+o0p6mFOik6PrfXgb0CYZRiUpY+WV/rRjaQ7L400lO0c6x
Z5tKifirxz2akkKjFAz4G8nbrfvVpeq22T37eLnvJgpAFtpnolIetZEyPK2eCdDn
vQ9Y/CIcMGWGvyTJKiV5J/8pEGbV4cnzMlxJmQoOaF4x2/t+oayZsldx+td7bXg8
hQebG5n2Hc+V10kWGx4zqflUKTpjgpwqjPFKhWfo/qBosVm6J6v0G7DC5fnIep3V
TZPGllNeLABOdxwZmo60xtRfIHxYEfadU1AuysoyD8PxafpiP7dwqbcGUlI+bz/Q
qfr+/tEqw06WRhRlyabGcBI2pWpmWz4QgaPlnIk9ptKllSA858ezIKnlvxwYcCI8
0iCKwREOMkQtO17txCxIgkXnuI3KZacA9MSrlYSLeXie1Xdj+s501zfqKcl7uyB3
wk1LRxXbKtWkFkX9/rgLMcoS5nPiiYC+UXIFjqR3/UjJqNQAJUkC4B4/FeMpyEY3
UvLMx5ZV6AgtR7CGSIrKHAA+262lhejMT7hbcsCiz1ZYrhdQ2g7z1sznCTXiintb
f8VCyjxJXKn9bboEechv5dogiUWFcXsv64p3ix4Mit1D6gK/Rzt4JAhFHWf/40fn
CYOWqiFDw6MngtMOb4iRqzCwbY/ugQTLPwyrd4CbPIsvwVjdng9QvH3dnLfkJbho
k8KWmbj+AXkYKzR82LsFo+IouF8K3/Gyh+LQobPbc+JO9B/UPDlkoKnxbH7+RpZa
TAEf/dg2e55EZg3WCeb+rXzoT3WsvsG7zj8r+FoLLz6ghjiKfT0X0vRp5q4fKSkJ
ewn+bxnZl6/BuIuE1PCnHu21W1NwqvkN9v5sf9iwyH0suR+a7yjzBg9antwEZ1bd
eQEG9uMZei/uZ9zGvCxvopL9jrHvG/IL1hBVl2OmvWkQx7I6XQdcADdUwwfyRooe
evDLZ6au8KUl1Hm4g9/uqmXCDi97HdWvE/q42EN0OewotMSbxhMnJNUloPUiLTat
Ux/NSP9k4nLX5ti1nK7crlkFmNg5sFrVpEvaPw0c+1Ky2dL943Jt6WkCjJGACt4z
Ft2lcD4Jn+uxLeToISPZQ11lE7sy6slBb9xTlA0qGHMQ7NE47y8JNr51cDKtTxjn
4I1CUiTjHBjluUiP25vZsgWbQnBAF/EXk5rrzjV6RIOGbZ9jJYaYlVG4QqWOYMct
OSyrPUKivAmw5c2dNo9Clx7wfOYuGUcDDIpG5DYGnnhLvlVWgfA8m/VZl4brQCkv
UPv2Xmgwp6EOvwUfo1K2OeZ6Ulb9cVxP+tVCAy5boM/61sFwQVnFyeNm4U5MBFWi
VChCxaJhmUmBt2zhYw0qshwl7MsyWsF4lZjkOzOnVSZo3BP6kWKpRRMJSrxbSio6
DvVpWAhh9uZgiugYA/mJvCZ6IanAdPXJxM/U3yd02GqlHMEHps4fMj6Ijz7E4z4O
MljDnmHkqE1Rwf5QrrXIH6A4cqHQYOvyuqazXq7TPrBHNqKLvKb342sd11gJWo5n
M5YetBQOJyxrbfcpsxsLPG3jmgeFsbTffaTv12NxdWUk3XqPG/6nhKIaYDL2QWUi
M9bhbolyQQwr8nP5NdyyMsm6hUg1zA7plwk7fYNWiYbjegu0kphviaGrj6hfeb7/
q340Pq50uN15JLv4jlR2iqVQfl7gyC1OpluLaXY7tAKou8p458EZ7/ikwq87iDvv
ew3mtQFste1hzbpy/U6aXe9ayAL7rK9IX60YoA9aGs2B32FBcdR8oepCScd4QtWJ
HSG1EztzVpRGoOI5L3Ql9a2JuOWSRlLIOyI/2/IGajfyyu14jLRB/k2MaG58xRUr
V3deeY02dv82FQnWfg0p/l0jaYBzrT8sIMBPx35FT5I9RW8yYWjgEvqYExodEIBK
TtfrtX1dwXwZUgyPv9RNmGiXuTI2XORc2mxsQPP2UJUa+QDIql8NW0t6VEQGjPCh
lthZrq3AWzIUn4uRHOyOTk0PLeyKQ1QJZcoqq6F1/yR6dqlxhaSddoqpR2OKuvSK
meS8hPyZESD+C9l8TWqd753zp6YsqSEOEGTH/4gruRRVBtj3xQidE3Y7W2llT5D3
PjaJVx7nfv1qWy9OzAOWOowfoZ1mT3zBvUM8+gjZGHBQwYc5tlbLu1cWP9LmGxc3
0+iiGMDbWG//rFSRxW4lUPnB5qdsBHV3DhyLvOiRs5WFzYpKutfiZwSnaXckGepc
+U8xtVFejaWdID/epFZNWqccEs2XMsLOYQGJuP1C5fP2RWcmjuxjQjqrHZ+YW4/j
+vPseIOSHqy6J8lA5o9wrOuDr8oGVl/g911ys9Mhq44vHOx7zMI6YKanktbRMVAW
vfl3bYOKjdhwEerQYif+ig==
//pragma protect end_data_block
//pragma protect digest_block
E47s8SpiKZbpqerh7AjmxucbJ5k=
//pragma protect end_digest_block
//pragma protect end_protected
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
/**
 * AMBA System configuration class contains handles of AXI, AHB and APB system configuration 
 * handles.
*/
class svt_amba_system_configuration extends svt_configuration;

  typedef enum {
    CHI_INTERFACE = `SVT_AMBA_CHI_INTERFACE,
    AXI_INTERFACE = `SVT_AMBA_AXI_INTERFACE,
    AHB_INTERFACE = `SVT_AMBA_AHB_INTERFACE,
    APB_INTERFACE = `SVT_AMBA_APB_INTERFACE
  } amba_interface_type_enum; 

   /**
    @grouphdr amba_generic_sys_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr amba_axi_chi_sys_config Combined AXI + CHI system related configuration parameters and APIs
    This group contains attributes, APIs which are used together for AXI and CHI systems
    */

  /**
    @grouphdr amba_multi_chip_system_monitor_sys_config AMBA Multi-chip system monitor related configuration parameters and APIs
    This group contains attributes, APIs which are used to configure the AMBA Multi-chip system monitor.
    */
  
  /**
    @grouphdr amba_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************
  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  /**
   * @groupname amba_coverage_protocol_checks
   * Specifies number of AMBA System Monitors in the system. Enabling AMBA
   * System Monitors in the system also means enabling AMBA System checks.
   */
  rand int num_amba_system_monitors = 0;
  
  
  /**
   * @groupname amba_generic_sys_config
   * Enables CHI system inside the AMBA env by  constructing the  CHI  system env
   * in the AMBA env.
   */
  rand int num_chi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AXI system inside the AMBA env by  constructing the  AXI  system env
   * in the AMBA env.
   */
  rand int num_axi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AHB system inside the AMBA env by  constructing the  AHB system env
   * in the AMBA env.
   */
  rand int num_ahb_systems = 0; 

  /**
   * @groupname amba_generic_sys_config
   * Enables APB system inside the AMBA env by  constructing the  APB system env
   * in the AMBA env.
   */
  rand int num_apb_systems = 0;

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_generic_sys_config
   * Handle to the CHI system configuration object
   */
  rand svt_chi_system_configuration chi_sys_cfg[];
`endif // `ifdef SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * Handle to the AXI system configuration object
    */
  rand svt_axi_system_configuration axi_sys_cfg[];

`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the AHB system configuration object
    */
  rand svt_ahb_system_configuration ahb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  

`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the APB system configuration object
    */
  rand svt_apb_system_configuration apb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * System Monitor Configuration
    */
  rand svt_amba_system_monitor_configuration amba_sys_mon_cfg[];

  /**
   * @groupname amba_multi_chip_system_monitor_sys_config
   * - Indicates if AMBA Multi-chip system monitor must be enabled in the AMBA system env when there
   *   are multiple CHI sub-systems that must be monitored.
   * - Can only be set to 1 when the compile time macros SVT_AMBA_MULTI_CHIP_SYSTEM_MONITOR_ENABLE and 
   *   SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV are defined, and there are more than 1 CHI sub-systems to be monitored.
   * - If set to 1:
   *   - system_monitor_enable in each of the connected CHI sub-system configurations must be set to 0.
   *   - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations must be set to 1.
   *     - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations will be set to the same value as
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable in the svt_amba_system_configuration::create_sub_cfgs method. 
   *     - In case svt_amba_system_configuration::create_sub_cfgs is not called for the AMBA system configuration or if 
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable is
   *       programmed only after calling create_sub_cfgs, user must explicitly program multi_chip_system_monitor_enable in each 
   *       of the connected CHI sub-system configurations to 1.
   *     .
   *   .
   * - Default value: 0
   * - Configuration type: Static
   * .
   */
  bit multi_chip_system_monitor_enable = 0;

  /** @cond PRIVATE */
  /** Internal queue where unique master_id are stored */
  bit[15:0] unique_master_id_queue[$];

  /** Internal queue where unique slave_id are stored */
  bit[15:0] unique_slave_id_queue[$];
  
  /** Internal queue to store unique id for each valid accessible master slave pair in a specific amba system */
  bit[31:0] master_slave_pair_id_queue[$];
  /** @endcond */

  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level coverage 
    * <b>type:</b> Dynamic
    */
  bit amba_system_coverage_enable = 0;

  /** @cond PRIVATE */
  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level cover group for master to slave access. Note
    * that you also need to enable AMBA System level coverage using
    * configuration member #amba_system_coverage_enable.
    * <b>type:</b> Dynamic
    */
  bit system_amba_master_to_slave_access_enable = 1;
  /** @endcond */

  /**
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_global_addr_from_master_addr()
   * method must be used to define the memory map for this AMBA system.
   * 
   * When this feature is disabled then the legacy methods must be used to define the 
   * memory map for this AMBA system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  
  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the AXI system of the AXI slave ports
    * specified in axi_slave_port_id queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_axi_slave_ports = -1;

  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the CHI system of the SN nodes 
    * specified in chi_sn_node_idx queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_chi_sn_nodes = -1;


  /**
    * @groupname amba_axi_chi_sys_config
    * port_ids corresponding to slave ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_sn_node_idx. This array should not be directly set. It
    * should be set using API set_axi_slave_to_chi_sn_map
    */
  int axi_slave_port_id[] ;

  /**
    * @groupname amba_axi_chi_sys_config
    * node indices corresponding to SN nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in axi_slave_port_id. This array should not be directly
    * set. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int chi_sn_node_idx[];

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the AXI system of the ACE-LITE ports
    * specified in ace_lite_master_port_id queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_ace_lite_master_ports = -1;

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the CHI system of the RN-I nodes 
    * specified in chi_rn_i_node_idx queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_rn_i_nodes = -1;


  /**
    * @groupname amba_generic_sys_config
    * port_ids corresponding to ACE-LITE ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_rn_i_node_idx. This array should not be directly set. It
    * should be set using API set_ace_lite_to_rn_i_map
    */
  int ace_lite_master_port_id[] ;

  /**
    * @groupname amba_generic_sys_config
    * node indices corresponding to RN-I nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in ace_lite_master_port_id. This array should not be directly
    * set. It should be set using API set_ace_lite_to_rn_i_map
    */
  int chi_rn_i_node_idx[];
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_configuration)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(amba_system_coverage_enable, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(num_amba_system_monitors, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_chi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_axi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_ahb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_array_object(ahb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_int(num_apb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV
    `svt_field_array_object(apb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
    `svt_field_array_object(chi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV

    `svt_field_array_object(axi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(amba_sys_mon_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_id_axi_slave_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_chi_sn_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(axi_slave_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_sn_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_int(system_id_ace_lite_master_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_rn_i_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(ace_lite_master_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_rn_i_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */

  // ---------------------------------------------------------------------------
  /**
   * @groupname addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param system_idx The index of the system that is requesting this function.
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int system_idx,
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

    /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing AMBA level system checks to a given
    * address. 
    *
    * Note that the system address map as defined in the individual
    * slave_addr_ranges of the axi and ahb system configurations based on the
    * actual physical address, that is, the address after translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] addr);

  /**
    * This method creates the sub configurations for CHI, AXI, AHB and APB
    * APB Systems are currently not supported through svt_amba_system_configuration
    * @param num_axi_systems The number of AXI Systems
    * @param num_ahb_systems The number of AHB Systems
    * @param num_apb_systems The number of APB Systems
    * @param num_apb_systems The number of CHI Systems
    */
  extern function void create_sub_cfgs(int num_axi_systems = 0, int num_ahb_systems = 0, int num_apb_systems = 0, int num_chi_systems = 0);

  // --------------------------------------------------------------------------- 
`ifndef SVT_EXCLUDE_VCAP
  /** 
   * This method indicates if any of the sub configurations uses traffic 
   * profiles for generation of transactions 
   */ 
  extern function bit uses_traffic_profile(); 
`endif
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_id. 
   */
  extern protected function void populate_unique_master_id_queue(ref string master_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique slave_id. 
   */
  extern protected function void populate_unique_slave_id_queue(ref string slave_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_slave_pair_id for 
   * each association of all legally possible master and slave pair. 
   */
  extern function void populate_valid_master_slave_association(); 

  // ---------------------------------------------------------------------------
  /**
    * Gets the handle of the SVT configuration corresponding to the 
    * amba_system_port_id given. The function matches the amba_system_port_id
    * value given in the arguement to the value of amba_system_port_id of 
    * AXI/AHB/APB configurations and returns the corresponding handle
    * @param amba_system_port_id The amba_system_port_id of the AXI, AHB or APB configuration
    */
  extern function svt_configuration get_port_cfg_of_amba_system_port_id(int amba_system_port_id);

  // ---------------------------------------------------------------------------
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the CHI SN configuration within the given CHI system, corresponding to the 
    * given AXI slave within the given AXI system. This
    * information is used by the CHI system monitor that receives transactions
    * from an AXI slave. When transactions from an AXI slave are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding SN node to facilitate
    * performing related checks by the CHI system monitor. <br>
    * Typically, CHI transactions are converted to AXI transactions using an internal bridge
    * in the interconnect DUT to which the AXI slave port connects. When
    * CHI transactions are sent out from a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. 
    * 1) Configure SN nodes in the CHI VIP's configuration in passive
    * mode and hook up the output SN signals of the bridge in the
    * interconnect to these nodes. 
    * 2) Configure SN nodes in theCHI  VIP's configuration in passive mode and use 
    * this function to map an AXI slave port to the CHI SN node. 
    * .
    * The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts CHI transactions to AXI 
    * transactions. In such situations, the VIP will use AXI
    * transactions and provide it to system monitor. It is
    * important that the SN node indices provided in array are not connected
    * physically to any SN port because this function will disable sampling
    * of any signals on the SN  node indices provided. The configuration
    * information is only to facilitate association of AXI transactions to
    * CHI transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the SN node.
    * @param axi_system_id The system id corresponding to the system in which
    * the AXI slave ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the SN nodes which are being mapped reside
    * @param axi_slave_port_id An array that consists of the port_ids of the AXI slave ports being mapped
    * @param chi_sn_node_idx An array that consists of the node indices of the
    * SN nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_slave_port_id and chi_sn_node_idx. For
    * example, element 0 of axi_slave_port_id maps to element 0 in
    * chi_sn_node_idx.
   */
 extern virtual function void set_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[]);

  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the RN_I configuration corresponding to a given ACE-Lite master. This
    * information is used by the CHI system monitor that receives transactions
    * from an ACE-Lite master. When transactions from an ACE-LITE master are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding RN-I node to faciliate
    * conversion of the AXI transaction to CHI transaction. Typically, ACE-Lite
    * transactions are converted to RN-I transactions using an internal bridge
    * in the interconnect DUT to which the ACE-Lite port connects. When
    * ACE-Lite transactions are sent to a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. The
    * first is to configure RN-I nodes in the VIP's configuration in passive
    * mode and hook up the output RN-I signals of the bridge in the
    * interconnect to these nodes. The second option is to configure RN-I nodes
    * in the VIP's configuration in passive mode and use this function to map
    * an ACE-Lite port to the RN-I node. The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts ACE-Lite transactions to
    * RN-I transactions. In such situations, the VIP will convert AXI
    * transactions to RN-I transactions and provide it to system monitor. It is
    * important that the RN-I node indices provided in array are not connected
    * physically to any RN-I port because this function will disable sampling
    * of any signals on the RN-I node indices provided. The configuration
    * information is only to facilitate conversion of ACE-Lite transactions to
    * RN-I transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the RN_I node.
    * @param axi_system_id The system id corresponding to the system in which
    * the ACE-LITE ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the RN-I nodes which are being mapped reside
    * @param ace_lite_master_port_id An array that consists of the port_ids of the ACE-LITE ports being mapped
    * @param chi_rn_i_node_idx An array that consists of the node indices of the
    * RN-I nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_master_port_id and chi_rn_i_node_idx. For
    * example, element 0 of axi_master_port_id maps to element 0 in
    * chi_rn_i_node_idx.
    */
 extern virtual function void set_ace_lite_to_rn_i_map(int axi_system_id, int chi_system_id, int ace_lite_master_port_id[], int chi_rn_i_node_idx[]);
`endif

  /** @cond PRIVATE */
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /** 
   * @groupname amba_axi_chi_sys_config
   * Returns if the mapping of AXI slave to CHI SN is valid
   * @param axi_system_id System ID of axi system mapped
   * @param chi_system_id System ID of chi system mapped
   * @param axi_slave_port_id Array of axi slave port IDs mapped
   * @param chi_sn_node_idx Array of chi sn node indices mapped
   * @param report_errors Issue errors incase of incompatible programming
   * @param perform_sn_cfg_checks Perform checks on sn node configuration
   * 
   * */
  extern function bit is_valid_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[], bit report_errors, bit perform_sn_cfg_checks);
`endif
  /** @endcond */

`ifdef SVT_AMBA_AXI_TO_CHI_MAP_ENABLE
  /**
   * - This method maps the AXI/Acelite transaction port_id and ID combination to CHI transaction LPID
   *   - LPID[2:1] indicates the ACE-Lite interface port ID mod 3.
   *   - LPID[0] is generated based on the OR of the AxID of the request AND'd with the programmable mask defined in por_rn[id]_s[012]_port_control register.
   *   - LPID mask in  por_rn[id]_s[012]_port_control is by default set to 11'b 0 and therefore LPID[0] will be 0 unless the registers are programmed to take value otherwise.
   *   .
   * - If the user wants to modify the mapping based on their requirement they can override the method defination. 
   * .
   * @param axi_xact AXI/Acelite transaction to be mapped to CHI transaction
   * @param chi_xact Mapped CHI transaction 
   */
  extern virtual function void map_axi_acelite_port_id_to_chi_lpid(svt_axi_transaction axi_xact, svt_chi_rn_transaction chi_xact);

`endif

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_configuration)
  `vmm_class_factory(svt_amba_system_configuration)
`endif   
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bys06tozaIpjWwUHvMSUGXEqo/SwKUWTXqSzpilBwW4EfrInJSR/0X33FVtOU2ke
FetWUhtjTS6RXvwlPZo/6zCLpLIcGPEbhvdYeSgXxO2P6h3jc//xQNeNY5uW3Axd
mnbJkBr0pqN7zTaGDl9q5MvWJbhf9DoHa5iKWIrk797VROiDOd/xhA==
//pragma protect end_key_block
//pragma protect digest_block
2iKkW9EmESMe3HzAT34OK7AQdqg=
//pragma protect end_digest_block
//pragma protect data_block
24+8+QFou3ILwhHnxCYlIuvTXiKDdUK9RGD7b1sFpj1C/ZiCzYpAR6qFcnuG1lGA
mhRsZEPrqcdbSF/9fwGmDUB6aSx3BJkyShU76KylSL2uwOu+KWc5RaCmhlJg0t4y
+XAgAnuZ/XpW57x8fVspm3bAZWZR7TmBjjs5LM8k+RVIKjMBRmRGOvsBuFBxVWw0
68EO8AU7iTfStWwACrFlOUnDGD2dMxx3H0dCm9dCc65+ZpEI3vdW+bp0/1b2xJKl
ELyEgpL48hPUpxWHxUYd3bDD/CXvCkbxNcv/L+WOCUkJ4HvBYBYRTlZ/tjx9IQD5
dD3qqwz43yt1DXO2jL1F25Z0RJWbuSSGnU92yZ3oD9qgC9locuN8qebuulET1Uko
gXxIiSM1OXFKzVl1/aVd2UUQFhVVAKXOyi5FUZteyQWOncXNFV4HhJCcWih2h8we
hvYGFH8As4dweK3UsL7nW5rQLE8zXhn5JPcRy1zuuJbKdez2CPJZSIyP+fBP+Xwa
ObyBjU/LRVPbz2kYEDz3EsrBypqUCBa9KJZPgfkrFftkri2mJCEP3SAyb9Co4hm0
f7D0N/hHhT/YqoSjxZvAioOip4KTdxMDOn/ISGJBgVDkbGylzkuz0DpZP+uPvsXR
et4YfDHziMVLHYpld8JF0bY/C3qxoceBELhPXsElMzJjSNCejOB+4bpdQtpj804l
Rg23eeQqnlXKUK6hrEFdRaqJN7iPnZDrHljBX17+sLw6kIKQ/tMIs+QNPATtLB/Q
pmocPxxwe6NTPz107jC6z8RQXkv4hWw1aLuvkhNrCK+uWqEyJnqMHhO193n9WiMh
hPjpIBfhlGPgnYrdgdXQIbRsBm0zk0DTFh700gX8yscFMo3GRjFuHswbqJyd4g8u
S7NxgD+bxGhbnt1tyriMhqXdNN4a3mRMXQKFxMqqQ1t4UlLIWLjG9e8ButMItUzx
ktHBz5VODRYl76SlNM5Jk6k2E931JORaqrfbtwDl1C/q8Db+m7BDoQFpq2mz8srW
Yi2p3csTCUecWafGMVOngw==
//pragma protect end_data_block
//pragma protect digest_block
GgUlCrd9sP5DfV2YN0kwgJeahYc=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2oKZcbvexZ+fTJSq3ZmvaXIu32hSRm2kN1+m3qo5s8wfnkPVw03TW8q5yEHq6x0L
lr5vBXcyyKtIuwdD+nsRdEgTOttM2syMYB3dIA1pYaJAII48V1vapbQg3EARyhRU
4+MMxG4I9zsDYRSKF3trDG4x8cxOOrIuKREgQKgWX1ttozkM0gR/bA==
//pragma protect end_key_block
//pragma protect digest_block
wUzizYzJi1q1TzSz4Q/c6uXx5I4=
//pragma protect end_digest_block
//pragma protect data_block
IH6S604dJvGZs9AWJkYsQZ7zeoYMpAgrrY1XY1/S+MokRBawneIyKodyodQNgDmD
bP4nXd3iicgFs0XxezkRyD08BQSKeFf4bLK7C67QO2AWTnSN3RikqTnALnMK00oY
ZLCnrrcIbFATACOJWXAJsXmPDvbrP6tafCPv6JCkzj1cKyg1TfcNwI3/BoOg90Tp
yXo8RXsinZKMtwi9T79dPPg08o8XAdgyg2FbCVUWgXgAaSPA0YievXH/JLET4slC
9AzbbJYAWCqLhrjI0npjtdC3H9i97SYHzP18N9l26SwdpBOrfUjw5Jm7fKNaf3+U
BVHJ6+Ni9Mjs4NctXoCLqBzDh69v6eFIIUNyxmyWcbOTcHIbWyQsQvq3//cT6D1o
ScbUyp1EGBcfpK/F5Sa82a7dUP84Ci60iZ7stU3ZKx7VKQXOVG59XVLXAN7Y5jEz
q8vaiAHAgUrm/2N5rKEzX0wYHBVOCgTTqBmvG/oM/0eHVmqo3M5S6neUCH8INZbD
Rf6t6Um866y0CQdEFWvfzn7BeYNMIR1PVfc9fgTeCEgrhVaCtCqs6OfpzcGijqBn
CkvikXY1oRPuishyUcLlYjX/lfYKnvENEVxUixEsPxKyQFZlNLEm0CJ51c1K1QkW
yhurNb1w+1qOAdyuvET/igcislAyFrO17HLlD5BhhlI5V/TBfPs2PWB2oGYX9QU8
VtKi6+J5+GXfabaOKwiZy2sM4dG+uyxlIWP5ZmwzfiYfxOc4QpVmBOmeNYhlW2hw
CkiVoVzOAMkdFB9INm36RYMsSkcSSmupPhflsDAJphYgc3ES3LHCymYcPp4tgfg1
/8gdZmV6o/VWBPZ1SLf0HMsPLHj6wO253XER4pEJXMYnOtkHdpv1cUFCm3zToUUD
em5WYVQUkw4nT4ISYndISrP3GDjG3LvVsrs/0ExIHU/d+SRNNgMC43u7ylqcQANo
UAZOUlIeyFVIUtDlRhjA69rA7lOEYFLlUSEdobibAZLX88EHkc1QWeJ0Jp00+2+O
QNQk1Bhr1HUVieVs7ZEhbkzfIBuOJI+QC7FttvXhmf9lYYRaySlpb4iHcsMJLhdh
GRrKKb/zRUY++xbR1VpBE0fTGzFGRQpsSmBdfn4v66vNZkgWVm4lMrrRnzegix88
3S4DEIP85N0Zt53sdBg5fJljyY35gMIsRJsXUJM99HjS4qs+ZG7x1qzpjQrMJjf+
PYdjuqGvzSMqMu9pJm2e+1Q2oEy2m5LUeVCb0s1uwWWXE85J8sKg5KY+nS4w682V
NdwTJ/FhkHM53M/V80HLSiSJX77QwZrMJw6eVmdKzlFCvmcvAVQALv/yEhjRSpgD
s5HPZ3QdEQa/jjLjlUOKYv4yWYp/zfwJLxekQVVTX+xjbAFz2aP43ZpNAU5em/IG
DNshkCQdrJdUYd64ly9ktN9XhXD7+kv783/puRTpcLglSjLBmMEfXsFRzp0/h5VF
VNZlCzmXXJHfNLN38gyYjjYFg0U+OjKcGp7g8VtxzzUJj5Sk0iCDCxD6W8HGT1wv
FAyZFpTCBS2zvRcVA8jekZC31rZf9RgdjauW2Iy8eBKAeNfUjKY1cqk2TuwROY8r
j87cjjm3cuEIR42qPwomUUQVLO6Tc/reB58MwBPsXFuNJMVWYaLkvDSYY3TYsipP
RH/rjvmD6doJ4nAJR6Q7Isj3fpsSiMxPWwzpn05VKQJ3KTA13UhesKPRUrrAWjcg
ZOuV2wRlMM+/1iNkz8D4MpdLeT18Vg0oqUSAjLRmTGicO82yKlglGiBLgociBKKx
DcGr/wt1VIOBu7hZ5BWuI/llBwh2Fo+IWLqATZKgnUY/eeF6+aLLvqafhIUAa8Tp
Ooi/WPVD02af8KHT2GPRvtHoN5KY8K2W1kz3v3ZFZM/rY9yx/dy7zg1ycLNxP5To
HbZwfLDmDlDK+hPE5jySJE3SEzhuBgY3ulBVpdKmrLzLByvlZOjFXfPWXy9no8Kv
wu4D0qJZKfmsL5lcrtG+NM/tAZe5r7u25nkyWuWjzvPqILgCyoGa5cWesSrmDFQC
0ySeeuDFrVTSYrx+UogWvfLUau1QzVv1Hduh/lN4jUlNevjHwL7ZS3zJeEVv0CU8
FFaFnh8p5Gj2C2yiOGeNsGBFk+en7HEKZ3iJd1Geab0cAntFmtnJSNRRbpmMJ9Jb
8Y4b5PkDqiNoZGzrL0PrH2LlkZqabdsQh1UUqzlaM44iSCwuECfvadInHCY7tTW4
c2GJbNUf8oZl/t5CtxYo9TKNhstDo6gHwiBwkzvsKWSCGqqLA8Wvyz21LPaq4Bru
yLrBpa8K+Yy1wzne4/7HzzjVgdCT3XKePYlffYPsbRM3DKGxSJYsqaJb0cfIIwlB
sKVptdYKz3nywpCk87bgk+qkP5MofpaVy4XvzVFzGsPM4FG0dL4Z6IdgnckEgvl8
fatO/cMAsmSglwPANo4Rox8DManyAcx8EoDzkDG1pRgZjeO4/TUKeV4mncMrGjHn
aTMDi1tqNkcX6B9CzIxMu10vRFs8SeIrmaTjQghAxEnml6oi/Um54AWw8P6x//5r
WPsZG25/f3YMx2Cg2tBaN+M2LWiyzQ7bCEOUFvnj0zWpmFjB73c6/8fSHahErN7W
0nBiHBoZf6O9pbheTylaBiUnEI4RVHUoPdMY5n8XQpbTI7dNesgmg3cUHWfq0BHO
BILT4PTKvbjp6DPU3Ndud7ezDjQ2Tm4/CubNqgO2y4iwMfC1nXSsnvn7id0Eb7oE
BtiJSy/ypPXDFRATF7TMQvxKU2rzOTeoSLR4/17ZqiufG3ZHJE6p2m+OOzMRWLur
XxEY5+u2Wj5SCL/t1N0s1Y8RM6L1pihtkEzXKdv+2rFgBtE9CdaTfcsddpPY0XHX
B6xOjVDqtFGuQMJMNNoxJ+c8aIENcdncsUTz8iB/b76wIwwhJY2jk/A28bMXdZz8
+M30jYB9KKxoTbizuTYEXcVAWeeLb14/Bqjz40lbe23nu3M9XXJ/zdlCKj5iKxwi
x9FqjGxXyJlGVIrPjKwQJfpzpX+GMBCiCYa7dXvrgR0I4vn2V7H6d7ObOiB6ewir
l7PBsgC3bxnwp7PlR4sj25SlSpewPYNFF1FkcB/6g8tos3KzX17KKTPzMD7mR+k5
4qH0eOkKtrGK3TN/q1pMV9jetzTygrE2KBYxaxLlztpt/azT3r5JmO4lmir7t+o9
xvOQBN5FrG9Z8sB/oxHJ3Tg7EVKHvTvGCgxvtUusS4XPfYCWdoFrX2GbKmxlIVaW
DWeoNBcL1AVzTNNOZ1MYV4SWFJhQlw9YczfY6aNmtyNyzGUZZcRtK5lPDx7y6B9A
mF2RemNvyReGvmxx4LfGGzBVXw7Ddj27Q1Wd7dc4475YGhMMfMmsJlMbID+8GIPN
i57uiuh28b9fHInb7lI5YESqkkZj9bD8Xq6M4pe4D0ayoBhz59XSKtQWo/ZF2oJK
DsMpP6qp3mVtN6SlacXVxIlXvaJltpzMywoIs6pwEqy3FoH66emP8psZXM5rhZx8
u7/18LptncmEe21lPFx2LFiGIX4tc5LqJlbAncpZalqr0ji2gAbpYz9ziKTWzeAe
QzsSDx0xxTNuKjmMZxKBrGi/IYwNyPX8wW3fk1bbBL+tvHcoEWFFqGmCcu4aaIjm
VBP5oEsZ8rFM581B5jC29b00thsgZPA/V7zXjPft8dPhhe2meo9IaM1mOK4SGhWq
CVqQgWi2ETrhpKZLJpeMCf8bwhEnEwu5IhwQdXtUWjb3dPvMK41oxAcf7gXrpuBO
zy0SmibBfMw82Tyr/ucDcfdzPnshd/KyHsUPLAypWFIkdNNWOyJ0U75GY51TpSop
UpyKdNLOfOZZ6OYEflZdYlwNqUlY5+KFANr1PJMN5lb+3c8NmCRFhiJbCxKk2Ekv
SyM+VPNlCzsFwO1lJ8PEd8hkQSCDrbUOd14fgF3uf3Pmu6TZBhnE/Kcb/IgpGNmJ
0Iq9ddFYQ1vhP90k3fMtA4Ar3j5K60DQs8/ftgZ0QXz5WtDgiMmItojq4ZnqQrLe
fe0iYNlpbt0fSGogAldp43tNBS4QJzKK14NbJmgt5yduffIUjqOw9RIjQgWs51yJ
4kNebFI7sQB/6kFL1xVdQqWvwC/s+x3gVpal0v7UAp78rXxnlWekSVdj/1Vi4kOl
guFyL04JV0ssWhrQeI9dDX921iVCmSYc2ds5BVlyRDPZjiwfafNXgl968KQOV0AK
iONo7/S3Lu1R78X5bFgnTZQw9Zupyjgk3zNSVz994Q2orX2ihAT8EqBWoTi16qmh
fCYFrEZ1M3BsW5FhrufWkLO80jqQz7FuQ5Sdg08cpcgCHuxngC0gBTd2znvlNwEN
143X/G3tMLUkyOf8mMXm31JE5LDzMmqKB8V9PLk2d56rttR7qLI6t+hMbCgqgeL+
ipdvm4d85TnQYW4cJXoodI6dvmFKiXiRzG0gBdp10Gh5dZYKYZsGBg/2/MpmFwWV
jblL0ZTX0K1EKdKpt1KpAdPuHJAzhVl72EypA0hwaa2PvL0QqqTUWkd3HGYgDSJk
gTcv9jovXVJOR3igDPq3fQYGUNRgIvHq291QxMDFbN/1GSq7UcQeeRMB7ySuOxbk
mO7PMLf7ZhVzvClsMbbhwjSYik30v76KZDn8GILBGibG3p4kS5C5ZeNc6p2W/LQT
NDKxziQBzAJvKo1ritvhu+eE2zqrKyXNeTauM56SlT3hLSSFZ1obhpgZt4oKXTE9
dnz4YNTPxDWhXLp4xLFq+3sPx5TQIk1WHq67xAsKf3NI1EA1Kb+UxRIqQ/1utg8b
0LbE1qVDf2ibgNXgEzEmeVutDNvNxX6I2HzE3HRuyNf1drGNXuhrkyOv9jaF/+cD
je1uuGe/awQnZBczcwyrLFjmzp5o4vjsYQitu4343Wb5HlSxm9yFPErzPo4XnUEw
S2VEa0YI3nDUaLSBBA9+6qZX0mWyvjo5egiPSTXb+QGyk5uKtogs4NHxnBDfHnTR
oTJsjbFX1f9eFF3ObLEpQyaiV/GP7k0wjYixKG7boYgwRLAf4thOK2F3B+NrpYkh
ErGgVpn8AsJANnDtDeppexS6VWMse9+GdKilgBBQzdT8kiHg13OTqhvxeBgb+Uo6
OxTaOuiNQH0qHk67MQAFW+c7JMmniynbnVsUH4DmNk8xVtOmNrljYM4xzmJzt7rA
Q7vrzjX8M3LNYlEwoxlGpf0crb9SIM+fYdv0u/W2nb4rywtuRw5/bEBMbMokupnk
O1Ps/75D4IvYNksggEI50kSbDFgeFMXIzFRPP4f5tYbDfS6VGRNnE9fYGz1bcuRa
qjxXUpyx2+5TxVk19fy2PTJJaUZvZmR7YztdHf/VlAD+knhIeqtXCakZ/reSf0FW
+52DtSoP3Zo+pNADLgjz9XjHVzEf7iOCYkRXkVV8iRhC05Qhta7PBaFsKNwraXVJ
GxRZM6FcfleYzpyFyaxcvCqSrkea8WPi4oBf+EMfhnCt2+hv0PyldESaeASkWiFK
Aux4HIiUbhv2ywXwkVNI4PEGhxn8pY65epIdGKHcE+n08IbtAw5TM0YA6fMhspyP
aQl+qwnjhcEE6Kkl0MP8NmVOmt+SG+K58sRTPD0/BckpPu4tFOq8kSKVLpv/1P4R
tLN5bqCmsNT1HiX+6K6yWD7KklBVD5B474DDS9prqvt9IyEUjOEOAbJuxjcI4IOk
FflhafYbTl4MXXh39KVf/TBXErQuyExni80zGnzq0gH/hFJa4QRUIhx7okVmWHis
U++6mt9MuoTkl1YKw7Sby2QYKoD63WYQl1vqquK/fwOGYtFIifAa05+036Jbui1b
WkhSINnLQGd7DIFL0+Hspm5/G2ITmFa2ix+JCa5TqvPmUosqUL19Cig/FHM3MlPx
DhcmAnN4QZ5EoOildfJIOECG7yFkr03ZORDRVbU/Pp1YvGIgMGGZRWNl14D02Nvn
7CVY37C41HT5ek4Sv3PiwgB4taqorWX0PR22iJ1Qhpb50lXwsc3iWcL7HlBkkstk
mBuM3wXMgxa/t8V8O1HW+5UEPlTJvY0droIpwVA2hjrfhNUMrAE4OxaTzRFSjang
GwYbpJw6/tT3W3ydO70Sy4HLwpGFjVlCccTzuYXKLJuOnikq9zBhMhSjxK0bB0kj
QVzZK9qoSoudAjwbIprH17fxF1RALvccl+tP9VvkkDiwAF0Ddj/hBFu95uhT+wpP
xFmOKbwEFE4VwcVGm9rriQjKAm24NpNA6yh4MegVmD1xn/IHua/SPM5eiqyPcE+t
4KBoi7sAHLByS53K7w+5r5TJv+tY/VFUC98pkK47zrwf8MOjz+BRTz3kgwEKnFs5
pyuv4AmDIWlwb7Ky0bv3PCUcMPvsmeVWHumxG2DR25sJubd2mbujMjAr3J3VkgS3
jY/H6ETc8W0Z6M0kKS358zuxhVakPhPknH9KxjOFZIHqVKm8fNr5smTsa6IscpZ/
DF8UCfM3FmdIwK2nJ8Rs/SJnTF+87vfcyG362nLP3PNGFlgRe5gHZPZMGu7NF7MQ
CYxekFyjzVQYkP6g1OINIz6M7soH69tkJHa/VgqaD2kZzPk06lzk5T/EgO3hLFf7
IsvKe75g1xZuUIctcLTLF1EIZrODGpk3//nIEFeJBS2f25xlK4DEx8txKuBNiS1P
NQ5OYR8gn2LAJQ+4KjZKjW3PN5JFd30URrguu6fuJDljg8uQNhnTqI2n+CwoOuce
pSesKEkirio9g1OcgtgNtm6sqjPs5caDaY6p8yvO61msDeqmBw4Mwj1b2XH/fWqJ
XzKzKZFklnz4WiPPzFTde9RqdBJkyNOj1qevj3voDrCFZ3s8z7VSplu6PHv6pCQe
9JbdXj76aXJKNdtFbE8/kGmnKZNtLvppLJr73wDZ+DwJ10FxPraHsQyMYJYBOlv7
vMsRa9WswCuoGx4qUBoHgyMzc+qS8gWgf0nERmgOHDbKDzUhRe13lNOdimVoHtDK
dK/sCTigMV2ydGZFsyQxDrLcEUNm7LqKvyXQ+p1YMUhGYS93IDfbYLSIjCvQKuT2
Unt7F6V0GYGx+MAwTRm80ZPOIlcc7Ry7+O8ETeApSWvQQHDc+DrDjBz4vLA3Is0s
yn2AknQBZpNUe0/86Oebc5AwxUpr+u7rXoR75S4eCvYUQEvknWHIM49yuD8tSq0t
jAi4s5bIlk1QqZ9axlzf+ASFV2t++KoKx4d29XPmY0vnuqmmpjvT/hB0gWi31kBZ
X3x9VZ3Y9O/0vg97zF9MAkFbBd2nztWgynS12EaCdiIiAHToHlbn2ulA6e9BxnS9
R0mADoWpRKDx0hoCCM53Ihb5i0uz0QRbWPWkXgMX3mA9esTmOwVvKxUlUIErdUul
jhgViK6zYYZYPA/7xAQD1cD/ncStMKRyIUwx2SgvY+Gv5t9G96Xs88VASPGId/R6
fHrxXbXyIAYJ+LsSqoh77+6VMA9t5XpbhL7iRBXB+5S9E5lK0Q59JW+7tT+zTBql
i8SnldjK9H87wJCXlejdIDCvy63PgUHJKbvHOyApmPEgF1WixVqKo1uw12UxjSl9
pIZt/wWtx5wqOIFJXYg82vbIvXAmLpWqyMQEJPgt6PwATK7KBR7KI3XqIGLUbs75
3M82nQyCfwB0WU5genca7X85nCESRqXP63k8BL6ZdwofWGxJvydgJ/0Mpgdn9IFw
jjZIM2WiZqvhn9I73Q9ece2U+0Abq8k34ZSzgXkMKa++09jFDbPpYkjLXnV+oUc9
g2pWhP6w18eBuDGG3A5+nRSmXGmN6NHZ5oVdPORmgHUg11lanJ28KxSf+yfooVh0
XKLGV3eIO73z3MEmX3SQuK8Fo6qAhZu5xbCcKtqIQGa4XnqWYKTEDsg7+HjX0Zxy
+RjZw/bwmv5+EZW0+NP82+AGNwqdkBkmViNbOW5r5aMNV+7D1F88mAb7Dw72mYqR
cllO8pQJFpCNGi6yKBbm/4mOdMMLLMGBd8TC5ZG2z0fpCu2RQ/jw75Zus1SNUXuU
HYp1RlVNnEZ1SUzg1a7WGqTxJEioTWxjjYIQT88yjLrOny572jfwHUP277Ic8Dd6
fF+21a5XVVBkAvvE0oZH0WiDbATTRkDLfedbnNt6TEBwU+Sq+jg60hO9lvFHEGX4
tv5qz5S7GNlSV21g2J6rqXxNy0wxgUSM2UKnX9Cj9i7kND7ss8fWOfDNGYkYYvRq
D3lbkrh8XCgRdBPHIcYTCNNqVhLlwTw6vJ6tm+Kd2dHkGPhOitT1K6iGR5ZOPKGx
l77EoovPJKuVlNp2xpagHpcrm/Zt1pp2VOl3OIPBLjHZ+gz5k9VYAK5VmWN0ApSr
eQhBjVuaAckZcuH1/bB4qC0j0kWV7t6szkeiy4xFDiDn4GSXDLPMvXqgmAvlBWKP
mmteiwbLkYQVV6gHjH4l1EWX8mU18bm/QfFacKnFeSBU0KAIxLT8W4JvMml03WF5
j4fExdZJUK+m1k85NSiHzMHGk3A+JuPx9TScQrGxs0es+y9SkZBf4W1GPhqjn6mU
soFjZ+EGm4AVAzczxAnSPNm0Mg/jAAYzySm/kYnlBm3sg9dDmu8NbpgOChFpN9wX
aSOJWVa+8Voq0IX08N1KLCN1Xdllw+w6iQILz9Lguruo28AnaCPUXeiXRpE8lWg2
5/TaUsHyJzYFtxqqueP4id6AXxCQQd6+f1yYV345GLZW73ypQeRFcs0PGaLGhjwM
7N7oh0JRxaMSaitbvqDrNVXkvkjGgmZtkX5kOTXlf8IQ/XgtrZbnj9UwqlBgC/3s
isHMxO6yIhUprmw2NYHB6cekCdYygJpD0KUnPTwoVSZnfea7mB1tp6X9fi5iwGjA
AISPYuvjh2PQ6JQrf8F+NsUvAm6tjHFAyf68By4kUOyKAwgNeR/ED77bjAYmlRuK
ulJQnCjvbnwmkqrTHjU/UcJEvpvB276mQZtONNppFmI1Op8a/qobhbJvI3cuGjZW
VWdBRfcFfGas0i21zYsf9MMCoND1V2/48MHAeGeIGucHVDeLXsEQLAamDGHXfJEy
KSJ8mgMZjMzG2il5kXPU/tWuBtRqYI/CsB31Jyv9oV9brV1wlNNrGA2K95x9MC8v
naoP1/z+X63U5u44mRtquTW0MBIEgFNbr95lKZUu6uchBinS6TFNVm+r+7ock+Sz
DXDh+Fkba3NJQzAllVpFzbFXz6vMM0E8+xiPLMvf+XWkb5iLn+9IZRWXgpn4rZFE
VXoBA2H5OX+vvC5eTyeo7k/wRSWlCDiEhwfd2xZu6QRBiUelh44zxsQ3Pb11X1BG
Cfh2x0rLWmGBWW+1qlPhPb2QJeWr4xpN8GCRPjSM37ajRN5DlNNI0i1WARELW590
Y2jKyRgSWmiW1MXC7NCsGbHSvY8Nc5kW8sWwPmoOP05M/Z7Z1woLxswIM7xhUTv5
Gl+wsQLFhpN8yHlRJBluwaf++4afwHkvXNuqN3cMYko/Edb80RX/nYaFPw0OoYef
fLycAQslsjegEFWZ3Twi4ryVEavkHGfsD/G1i6MjTkr611vWmTcp3kgc0VKhZizT
GLKCEE5fOkIv6BBm1U/t1TWTajFwp0MGm9PRbsGt7XTTaG2APpc4vs5UE82mB7ab
9m74snfrihOQULjT9ow2XQneJBcgx3fcsLuAjtDOSYd7WbwPJJtqb3XQlJKbzCuw
5AZPY/chxaEpQYSEGQ7MmA2FF3ApASGBhftUAmWzClwxLtrPb7rxXY0zA0TCAdZi
7VT5w07FGild/SFUV9dE0wj1xrzeERTiur/gY1Lc4ZNiP0VZ9PhfOsWI6l0wVNEH
Psy0iUld5Esm7OTntscymq5kHr2PeqL/ljAPaIJla4YffVurQUBs7E+K1zUc1wpI
Qu76UKU+BK1ECaAjXrqp05V/YcPly4l/oztd+ZNvumUJrTgnrKj0XpKFXVVLx0uP
mcKw7auIE2IchDydjdxpgNTn62XPU4wQ5rnHVev9iGiPdKna4ewkOpCjEDU8igd0
LYV8ZZB+a1JgREUpMRkICjSKrS2v6O1neTk+Hn+1jPXiwCgj2RVFdQyi8g4ojRxi
y+Gq4RhD/BfdeVvcqz+ao4fXjI0c9BgAb+KF7urDMg2OzUgU9EwWw3Z4TFfXsE1t
ucv7+Luvag7krQGFLb4ODD0cLYsr8xs3Mubxvn9Ugg97b4EIFWCW7ETm/bBIwGT0
vKIATfVkzzz7dftBziq0V3BR9QOM2XJc/cR+4239vPIsRTWnNzCsu0vqYk/qOdwj
mL6q3RMW5/cZ6wqNXAZapgFhqaCVVsrN5J/1FVgD/jRwWt4lcr+zkTtYfbr4DvYY
+qlWc7QFeWgT9PfdxYFIhzMO38EHWGmf9fDtycl8l/Fb5wH4kOqqdzHK1sEZsAQm
oyrTF3k9Ymo2rZX9qbth187c4G9Y6OVO8cf/WaoXGPID+5AbEZ+/B0O3pbeDtQTk
2RL3U0jKn+I8RRc0jfrq6XBvO60MtCWy8JXi8dBWF+g163D69cATFTGTV18GAgE2
m9vMRP4nf6MeAte/beQZPyy/OFsYb0hgQfy62q6iom8cR1nZx6bd4s5Duet74PNf
QNz1WvU1KRuprYZLox7EzkNsM9TFlJFBZu9gbxyIgWPoXEte0JU2WJYHaRX23baT
Qu2lhYRvQ51Gm1Pg1Qh7czdljNZleuz8ZgVoz+xHOY7tqGKSsi+NQw9IWRu1NyPp
WBZyrJu9h7qtQ75P+uCPkBIbiBN/+T8BkGekSegiiV0Zn/uBBvkLkI0/i5pSAosO
kVVuwP9m/tIuWCoHyBq79d4SDWPv07R7E51AbYtDbOz5m/w/lC+rRQucysg1JVp7
Ow4ipzn866NhTJmuc9WD4sEKkDQyj9v6uwOs9BRJRnQWrJggB6VxCMBP6bh0MgZm
0AikfJA7rlkqZbzoWlQj7e3Y1vzQdPyflLk4kCdtFAoi12SC9kkEyxaH3pnb9CFz
lNfHWvxmztch3HxrkJVhqHj3lfXBxHpofCQ5j5sDdsdkTG7y/OpaWwADVqW2S9XT
/23bILzqv328pY+R80O2U3UQCJOkWeb0V1IykSVg5BU9CbaUnt5GZ5rYPn1vGU+N
97K+pati4nekEniF8MgxvJDvItpBp7TaRAoxDyK8KJ2LAKwLHvMIYjQ0Vy6bVNwe
iYXQHbSLsAcpCIQ3BA5SE5qr+vRGNfYGTEKFT9afCHiTZneg7vjONIUl+x0kxZZi
EC00R5ieRNCafMy0H3yvkwnl6oQJoI+q1d9HPGrL1ofyczQtOHGV8oeUmOTMrtec
0k9DcSeitYtXtwAY1P6g+hG63Bds4POWsWydptcEK/sp6PIWK7zX3XhJDHNXyhs/
xNjuFsFqcKhiBYviAKQvhUT/mimi+9rV/A1ScGGNk3JCiixrPbfyVkRmB4gc+v9r
inLW/QhX/l3xLdSlvDgadmCv4Mct4bgn85tPRjvJX+I2gAHiEqa8i4zoH68qshmq
0jyTapNQQqowpMqayYgCjf7pQX44LFyUiencfXGJzgd1+ef87nuCSicDYBa8xhpC
0oun2m4f0zmy4XCrBsoQjq6EnUSwg+hfEoGzGEefOYGiyR45yGgNTmxQd2Soji1D
OK9eZmG+uO0aXjJLQaiWF3OIkkR4KWtkcGw38eXvPz01XDgGKsBaktAQrAfxkUu/
FHyMth7v2IVuywu7FDDfyGkzFlJX4uYmtnA8cjPWPlUirw5vJ3muDuVpWCtoLHC4
hmwHkKn2rQN2O2aR8XbnpDZ7TRXqOfhLp7GBo9kfiabq9f73UEer2u2xrsrokzSD
MmTNnzuNpqVYIWUJhh9yY5sTROoFifP/0+sam18oKKh/zlSQjdc3KJHKmEIH6Nnt
Nbc2dc5uxhlm2b6W7lAyjq1wYS6r+AqAsMaqbqsGRwyLU//JF3F3Ie4RLE0I/92R
axJ5CBg2YqkLRBW+aBe1ttcT/ASg9tTBsTkQw/ySSyY1HnZ6As9PuunNO8m0AT6S
ZA5BtBVTmjrWU33lc0dOTbnkNzeL0KgMZdPW9XvXC45iQOXBgMnXS6vSHoNES3eJ
HdQ60ySfmzewEzwusI5kFT4vHEszSw2gpJpJN4BISKkzPUlMEQ9Nvrt0+5PLbziI
NDkwlw4gQYpeDpKi/jksdcvO5qjNPF1JyHWcoAhCGngefV6XTcXh3KTxxKdib01T
kDHjvNwUCi3PVHu5DmmSxCvYrWNLxj+QiTPZUp5nXs60RYWyPQNhsJx2VHDBh17V
z2qeFqL9JjtXkXBPNwX2HGcUh6GQfNVkZjpX0TOMYYjMqQd9uLUBM6scayZ8yBjA
1LEFyWd14C1jbBzDRYYy0ZqxcOIv1WRzo1vfS9e2DI/v4rd+MX94+dj+G2jM7cK0
W4a9xzHKNVWqlzwEk0aNTtWcURGkwGKgsKnfYxXcLyHGOfiQ5dMRqSfYDZD0VDnp
7vAXOb5RuTvxk6On91bUxXDcDAS46CkLiXmqnCzYmrZLn4A8/R5HoZMG2jYk/IOj
EJCOpSxX9bNqUbO6Lxc3zcaW9u+pC3iOm+EmscMp6Pm0yZmlx0SlE6UFHT8rm69L
DVw5t9DU2FF8qGcyFzvbAROT8+CSjjBWZqwCvSFLZCTE4PF/S48nNpx4GpWlSYen
Wt5g3jctDKRFupyZjETYdAA43c6RacKgl6kiysW9DcJTO54m1nVYpkOKneePQ/Pt
fqWBC9BFnqOtUwrrwaJPsb1H6ByDirjiJmN+J72m2cf/vVHj8vQc/YbUQZcU0RcU
uN8MnVxdFMnh3nMmNaKYxOpws/l0QTr6Gm8gnSoHfS/3VzTGsIx3535ZL2dzJXx7
klX27tbDZBmVIo7Ah/T4xd7gcvQUaAyy5bVJGZlZDFm7gDksFlVDrjLRxqOmdvqs
aBFd8Den19XpZU7vk0D6FpWZ67S/jHugUf1EbaAyEM1FtMKEXWTKj28N6dmQlD91
x0ZInSy6rD5l/ftBKpEheH6ZuRnkDzk3cErsFAdwmW5RiO5+7SJeH6VPi47+cPcX
g7fgNZ8fWopmtZCdcsboto1YP5rpKTtGfw+tmNlpUdDTFFQhhGMqnbm4FSPaRBzj
rSTeyYyDtaqfCOnaraAYnE5lAHzGGG9ND2Oea2H1si52CsoT7zOAyNcOmEzFDD17
/jHu5o0bXi0AQHnU02EVgIAZY8pMDFSOPGSO89KxIbx36GCQ9KT1uxCgf6Cwy/ea
qtBfreStMmNFd7BDU6tEiBesu8uB9I/hXtUKRYXJmY9n+/BZQAs6P8tiqZIOO0FE
69TQMVQGpa328Xy8Ivq2g2iEUDK/xcyTk+DEV9aR4k1liiC64Aputc4DKtYuhALF
/aDepySzRFPohaazyuHBhJP8jShrqZAtBO0Ic8uNadBIh0J9PCgvScrOZk3A2mWg
bhU2HsiEvw9o5isewSKxbl/cXsjRNMuEwh38JBqPJyoFr1Iz0Q9Fsdp9ROZ2H2zX
68miyw0NuY9IPkw4rIa8GgU9nZVhY1TI0yakfkC2Im0wBVC7CFbfnW8CL7Ybsug2
FbBz9fqmcIisHiLsFLdfwWJVgw1jUzBU4TCdwHtlutBkvtlgJ3S9cIszJF/GjvWh
7GgSoNDtOTsRKIxNuT0z+MWaqZ6CxXTappIZyUOaNoYjeUYKfhhm3YFPMwyZh2y/
RZ0acAvjeC1FiU5OQ324jOc9aZduD/Y3jytVW1T3r5sfTNhI8sAMuPAIVCI+Y6OX
pnc4v/HSwJwgPoCnQaNY4eWM1LyyD6DikMx+1Zkfu2PCHVpq/B9pRRS1Sxu3+fMU
Mz+/IyiXrYYHZzDqp2SMUZCQBwFvy1e633uLluTGD3dyz8pufvy1jfX8J5tOMskX
h86hw6Udp6ZaS3/hlT9D6B1+0oGZEBQyU5l+guKK3zNE/JtTJ4Ms/q0rUlN/G/Fr
bUOoOB+aBN2jo35udxEBIOqyEYKQJgYJQt5rfN6HXFZQ7fAMV5ndVK5WMXR44aoM
/AgWV9nZYpGsxh6ZarXjJMHSexKl7MkweCml+Fmksg6lOCt+liUGE9PXwDqEpP1p
QYjfkMk+mgQKZbwwp+S3jJh9ezS+W8jzDF9WPDXqFJv9ydJoMN0TDUPzPSvosyfq
COsrqxtRfkzwGpThRswcqBmglFYFB2BtQFojcVfp2QasI0EJBp8MeNCBNN1R36SL
va/j2TIfmSyccgih5V9QY86JeEwOKtdT2wutqXcPYBLKAnMa4Zd2zhKkoHtvX2ht
+1hmiulvfUK0lwOQIVkp+jAvgtocC5p/QppHX7+VQ9BMjzObiFeuVsYOlgSgYRnE
2YKEOvdzM2BeG+d1HfiW+i+8AoUnitiPUOKqPUs3eAi7Y6A2Ib5QSrkYKoCaTLca
XoLdFcjqDU+HF/21LHf7awAlstA/ecFl7WBA89fxNxCCO1Z5d4kqP9RR729rUstJ
RqC4sKZQdUXh52K7hT5HqhnniQfRG9WeOhsjrhUFMIAAL/bt4brV70N6rKwrEZMn
WxxQ0guSlTKFSXqt/zK1niQ/ZT7zaCi4sKQENzEUX/dLynnAjV6Wxnw2mrh9WE3o
UKMY0WFI3e+NJm8a8m2T2qIwhoLlNovmBiifYfZnNprvgzyjBrNfJ+376kNTWpBX
rIRSAqrLJrhZtNZ4N4xyy0k4cAsFX70LkZY6wSHW58jB+OOy/kGE2zbgIO/Bq7mQ
DKVe+tvc0G5wba6b/F4hN4xmryE+C857sz3tpTlzz8zZyaQljcjw3M/mQ6ZumFAV
CYv7cqC3gvovcIFyUReOm+jRhXoDjJBAtpeHi107GXibWaOYpB8RmtBtWwh+OrDf
nAL68uEbc0fAE42ypAiHAFteCxUqrvnr5kKmKm3RbwvIWt+9sbl8kqgWjpekPepR
5aiGxsyoUXsfiWIjoSEXrPbb5rw/Mp8AviEB4qyAXRF8G/aQTdJqIwMOp8KlYwbY
EL70jAv6WdmV4M5kREvM/Ohs7Yypx4rsf+P6KqJwjo+5G/kJZnCTbzVxvnVGKkKB
Vy5xKJK4aLAGc2092B0uCjMZmEOgwRMBuNwLYtbTmied40A0GcC+kRWl/DtX+LNT
qyuMDRKSy5X3qp80c8E5bTkAgs6A13ap9mVWKnRyHZYCY3aLp+4Rw2YHoOiFXm2A
lJd8wtb22RjNSw3inyV7ES+UOmxSQlKy3lL4DDQjq38l/TOJYEsAM+n4fXNADjyH
J1Evo5LiNTF73OvFuFM5fKP8A2PIEekmo1MHsNT+JB1YVXuevQCMOMpKQxz4GadP
3w6nFPfclmM9/0jv5WYRpeOSRtN8QIPk+QH7Kpp9GUpPnW1mmSwJzDnSxWh5a4vf
LTSJjUpsKmY/0wdeWfv0oA+gEDoMZTKEje1cu3JbeMaNTM9NxKzVKPvRysZiDvdQ
LkbMCRavi1RvkN/xhk+N7U+pOj/T/mGbPC9nwlaDB1/B7icLDHvhNCAafSnC1N6o
ZXw2T9rGdbYyf/1GVywF2TlkjjzsbgUY3d0tCQssXpPbR5sgCkvqHV9bJWnVImle
XjzlUOwd7VWVwRT6AKnWKqwBAYQbgi4Mz2S/M59ZDBU8jIqiupa75TkUsFaaW941
8Q8WiD/Capgvqu5ughe1xklizJoORcugL0QRb6qejb0HiFlb++Q7yyWTFjKYqyhr
3rZhiqNES265F6QmlilBMKHgkJMEaCXChejbjKReOyMdCaLc8GbaSSW1/zsEMIv4
EJY9Vjv9t3ca0ov5zxPAokZE9xOgGH1+atYOzXlz/pJOxugjxGyMyUK7Z2Ndx96g
9QHTeGQAqzLwaUPmPOPMCqZ/WGKoXqPngw0g7yjr2Ieg1RBatrG2SVYyEor/br/x
eA3pjZNJ3TO467RH4zxDWa9PbK85otsFj35+HQfde6ca2+GeEyce9QTMzCq2wsO9
8L5RojsEitd96pRNc+X4iq7sjzXd2CXsTT2WoqjSWMlIAwv5T6yYyg8NPaua4CnK
jGT/Ts2A8W6EAHuZRPfE9uPOlNuyDsqOgAZ8/XYgFjlNLYcPtswn7kAiJAah9G+/
yA2/tWmdCbgK6tuRhIllSbJuKXDRYrx7jS19qhhLscPVdz5LJ5If5z2mj1R0GGRL
nj5Rd+2Z7GQtON79gB2ddnvdjQfLHqHX5zmMrOaya6aWvEr/osekzwPoMt2Wm4n7
LAvNJLcOt0ZSoI0CH3QIgn4h6lHO/oJRzOeL5K43xsWQZ/vd4hL3UqP3lqpNlRbI
0cflGGpsZemhgS3KRBlerBCsFZ3aIHuLYuYm+n2EOsng/PmwE+u/q+cFTKgLJ12W
5gk9uxCBpxlxjOBBaP4Er9sy42I3+THuxSrv5hkcjrSYw4Fozc4IxYdsJmy5Fv76
lgJ+26pt6LYouKF0Y0LkKwH1xdagzHXOw+e1pw0RlNuUv1ikcZ/PCx97CXv9lUG7
1wYn/bbMfDWGF0MpeDdbXLeTRfpJLLP/JrSBdToSpPVvvS1w7iZ0OSXAwbInuw5u
dASWBHJwP4IBFJegVesOokOjxC8xJWxVSIocX0CnQVtC8v48wnm2p8JOFb/JIWer
JXBoEFKBWrKE0rY9IhWMBwzOsXj2xQMXIB+MmD6/W+FYzjtt3tMSuBKafcbCWltT
POuiqCl+5F6CTwcr86oAPxlOHILdDV0O6Rab/s/slnG9HXH/WcMu8HUO10yopLMG
fAoKeXgUX1zuf5VblT+vT0lR/Ny1ZFifvsw5gV51RcRmLIVHwymFBfm/O/nbRPDn
ZEzBoy43ES4cDogfi4vwZaUGphatNT7kpp2ewS6yqsnVl7HeefWX/IwDXWOBg/hs
0tlVYeqMi9ouBkNBTKSju2m9odWJU+tlPRzfyvEBeuGi1IoHUsA+9POvf2cimPkV
0emSoF30GPZoNOLvd5oatwMwRtbvbIsCDgG/zO1JvOCp/9wYi+EWb7xD0TGYGOQe
oaceBu9gZMip/BQgBbtPUYCcQfxcDGcvOX1fmaYZYxg4iAqhr2QtgN+MdKjanpyc
B+Xp1RT75y3JCLBSe/wIxSQTPJPfAGGFwKrJqN/Cynb2rXnnjubWQ4oeNZPTsGZw
62A5/WEvgKhMeFi6JzQoNt7UZ5DVmwTSS5oO8TV/3f+iw3dTEQh4cbAtQhs4cnUX
TqmnC6N4IwuvwDF7LAYWA4kUCq7LNTxCpZL/BlbWFNJrYPYRUYm/oopnPKUQIX8l
xxxtnRGvfgsZfZWWl/h6n2vdHG+7hg3fLYfSsMA9HfE3eVIZbMtabOJW42EBP9s/
WVBYeGWyx2L/zEVojs2J7OSL58jhIwpgZpmCIHJAIulpCN9sUKxIMETlFhYr5VCL
hzpNvkIxFQJjY72LwfPAu5VAYWsgFaixq24DvUFnCOEM9QguqVewIoUSl1l2AQwD
yFqBKxRXOwh1c88jtbOPRE14E7ftDek4fbLrbTxJeqOyGA0kzzvVnAErtltJr8sH
5VnfnkCitY+KssylWfy81IPQRv5B2tNQlgfWhA5eYhTleVMEO60dEyyt3eN65FSm
R7f9ZNX5le60SHgS5LNDWoKI1Pb7Vdh9R1yME/aaFfgyr9iQV/izvaPxiCTyrmOR
5hrPqU0PEoUnuz2xXKWZan6g2G4E4PFNnOCVqUGSswMmCLeXA1LYKl/maOm1zGx4
K202nOlkIpzx2gOTPJNV8aZcXOTbuwCpeZulDEXwLZgagIIeOQGMpptc/m2u2IKp
Qta8tQyVoOYHqZ+4nc9PQEERZJMt2F+CKLx9e7yQdGR7hsA5glQnB8l+Upq7uU38
UAxpgcjx9qNzx3Xeyua15fnme6pAsCSKEHhpV1/4u2yY7ArB4TNZsZMSq2rcewpq
tL4G8J3rKdICSjqklwx+WPLBYEqjie+ZK+9q/MIljb52DgjdTpraOiCSa5BCw1lT
Frag30VZADyR62yIXJM0/cAkcdXVEM2n7+ZgtuKuzwARo2perB9kJ1/20j6Txpez
cQ1S/ivE6JSirdXJC+w1+xHbBoz4/0mliJHyTHO3f6TmrvQNjzUa5/ef8OSx7ugr
+IJM+n5LNNDi0BGJDoEP8uz5/jmtfJ25+nWwIM/rg2l/NtQgPzmC0RWb3pFVbSXM
hgjMesQFCnGWjv6Rer5xA9IgekU+mW4/s6J4Y5fce6VlAT04RVjuTFwGWIiJvSyX
waP+Gyqh1e4Yb7rRqA90rdLfJelGa5k9JgqBhSsSu9UFhgsr1qfMNRLaxHOkmBIX
23LIydA/fhuXhNervkvpwkDSMq9SmBZQ0ChyqGwc+u2kf2oobMF8ccsuTSBpVGIH
8nD193CHA42tK0Y7EufU8IXLKeZUDncJgXmf5KENZpIYeNLe+HBy4mQNPd/KPpXL
LvmSCnw1G7wQstawj7/lqQcXe+d2gLCj2kY6UNbZ/XojgH2KRBPQkyyQNR4z6dlk
uOpO5geyuAIZ9USPSm6V3L2EF8nhtN4oZeAzPElX9XCqX56Apyja3JAx3YCV1Xv/
9XCf92Lu3pFxWbb1jzVLiuAeMNwuIahKOB86/yZNurUaZ2iHkNE2Gd5rvyJum3bb
eAVD5Cz/oydV0rYLdnzORQqNLB4yah9dSqDjz04IVhy3X/uPqFlReYN4N6B2Cxet
E0apt1rjycCMrn7JDe5caVgWeiZuyalrEiB4R43a1iQrQrsONM/cKr9qTejgv37D
EviA4I0QQTjo+YQHvVL/sMTNY8Z4WK03+3UhnnPsC5hApANJBqkrBAfG5FmByQN3
qnd+RMuidrukfQrBtH1u1fEmrqNwf9QGUY9v13hJzjXK0yqmxdbdLNQo7b/vIRtk
c/CpZmJRTHCMNmfmw0O/37GnTbc4XmjbIvs5AigFqNeyCFVdqWiyPlZ+on5t7LfX
kPsJp8f1/vL/U9mYMssARH3FkN1Jz2HKo1Uzceo8706QmIsGhg7ZVn/HvENA339l
0woD14HevCpD4WyizVg3dBvERsWTHB/Ne9bv8Z5w3xCrV9y++BJH4NW4ghxzscWb
sh5/1iqSxd2MICt1tMPU/+BJJAs0nCIxciNBABNk4nfylzI2bBxkRlWyPLWdqcTW
AR/zzPuIW3R3H9Ni/yZurqvBg/lMa6Nq5YueE/yvfE5qaUMSyvkNEfKUyl1Hwjvz
Zb4RKIydYXtBlhwHu1p8WRIDZ4mgJKHHzA+uNlpPKiVZm9taV+gMOgr3Krcff6A5
KCu4Vn3dfNekSwM6eq/NbHdtrcA0yLDdIHoSvnjGE0a2IBj0//2KHwm5DhiFgjFH
5SHRmNe6Im2atdPQrYVaAgff8cUQekgJf8Q/mJRS7vyjH/8/cqo5iIWnuOS/cXxJ
QGC9z9+xvh1lTcirw9uRtVCAILUAQXPfP51o4aOKIHGSL7mrdN6/n1MXZ7K7ufzs
g/+ifOeHaCHRfCiJovCFDIyNeXmdhKd/sYnnCA5AiN29J6+iAUoZYrABlyqUqdk1
RKSJL/oKFiVFgg6CjDhWExzWqhG3egwCd64YUmjxfE8fWO/k33mwGqVGwpbK14Ex
6yHw6kFT1ZDZnnM2IXXvUHt7rZCTw9u7GBVp/BzhFnq8TOgcFgsagNZABweSU5CU
ejRoDfsu1FcLIXca3lyMcG5is4+C9yCJTWPxkQFb2FzCk3AIM9iC9UhNOeqX/Q2q
VU1upbrVJIGxGXCU22DE73tdROmtmnVPg541ip00zcLJbP11ip8XOKhHpK8XCm65
arEH0KCbzMR0Th73Z3tTD52XFIQq8A9s0NB7EQH0PjKAlh5mYUlbGCnRFK6ZmwqT
NmeDLBrg1MeUC4ji6TdvNBYhkomniL+MiQTa13ojJnXykDsRqIq7uc9Go2Ct5+Lk
7vFwbYTe7OYF0mtsuJ1TeiWa/A7zAMYTPhyLZZJKxNei4iy5/eIQRR+0PFNHvLZ3
mWA383qWrlJH1Z6r+ORt3hB1Iw285UqN2GirT6qpE9iIH+IzsxgDq4Anp/hPPzls
E9zJAwu1qDg6PCBYdHPwJN4aDteirDhRQKIht2MRBEcDmhwh4hXEtwATpGkgPOz5
RXQrum9nag4LmWZnX878Gf9m7EboJqD5Wcvvmwtpt7fCVxnoLZEg7VCP3HJUlbL+
m0+tTcSg+F3/mAMnIxn0Q/JAtOUgsjJ5TYCn0E4eOQOudDyH3eSwxxEuq7TTJW5L
3j0AM1YbPbWqrJHwlkLJVgIw2rwVAV1sWpPQsujn5Gr4oYWGI+yXMRkacx6Drsq1
R+KOZ+/HF8tsjPnJkBrirKvOpFp5/fCKmjBIW6boJ7PusP/t1iKzmOssaZGKFM0s
fs3W17eza6b9fEk9EdyMQjHc07xzEb9gCAqSTkzkxvEpQnkH5+HVJxRTlzdCmJho
RwVIoV/mS3SwiafmsU0xSO2NFG1VXBLz1uO3+hDIXfLz7pSfzzmySQIvUEjb/eBY
10WCgqI+HgVu2RV1JofivIlsPW4v5czU6Ukt0MDetTJfy9og1EZ3g7pvBrf6SBHn
Y67cq/tX5F0O2rhbFZAg/xay+FbWTANzHDfqNCApOIFupv0MMcy974r7Iq33L//x
5rB3SEyuFLg/9DBtKdXiX6gzJ21xgn3TtjUDMf6JIaQnUSh+HnRlGr8Lur/R8Jk2
M8o6Kzm+QTGZ7rGv5kBBI9t3Hdw98PxSGHpz7f3cL0EPAZIOOnhk2yJYumimUbRx
RkNV0WToJ1kWNwFEnAmw6KUvpb5rOzdoR9FwqkqoDmBBa2RIk5NKmQzFbc5mRF6L
qiwZU0ANeJgdbUCoj3gtFI5FBj++K8dCuPn+HtQwrtLqrydXw53HzRiCQUNG+AwL
AUHoHQKoT1bW8hGOJBQkCs5FgojtsryWVlt4JUbgTYSocEeL7n/Nplt7kU3RiBn+
FraXXoUFb+hn+/1bsXDgNtXdPdtrG+eKZGE8cFpYMXc2InMqQ4mWLDmNEceU0G4m
wBKd1kLdCBwW1Obo2ZZpMZgrbmEXBjhY1ztVjgmPdURNxoZ/4q3lq5wlHJ9pVk0h
f3mCMLi0Vqp4VX3KjM3K/aMDGPgORTxUEKZuSP3pU1XWU6tNUOHnWGdMeKCqxv9n
S5+uGJvIx4qDLjeCmAN/mFDARbEnuRk9Hkl0nz1mTqTtGrJuGzJHrppI/xrqzcfE
BRR4RAtdl9vtYwTd0T20nxb5kZDsm+eWTHdqhY1QNM7XlBOIlP3tC6gfV/x1c/Cb
tSEB+OGBzwt+VIiBTCjLv/u1yz7ICLrxEfEuaSERbXtmh9nD98OR6B2yk1XL0dLB
SwkFTTCvTVyhLexGmCOgtuG4AKDCTNpg2uPC7yLD45MNh5sQN9W7/pVHfzwvXPnX
opt59hSrrsSOpNc/Xng1oTg6rPYANLG5tb7TbBcGkYwWTByK0AzWSIX3gKyHMGik
vkGeyxpVWhJM57m7izrZF2ZIrfCF9uhm109590WxD/otj9oUfNWnjbNsAvXCIpra
ZVypIIn4gBeocHTfpgzVwr2IwtCDdmUnMkAzqYeXvauxJyDTjLVZnCZpPYu69i2Y
i5b079CX8tSiorrtvswXX+TVWCjPY7+De6QUereUAbEGyVjNAhKW/0KAr27VHi2S
CR9/R/yjElhOFSJYlw+fTIOIqLPBkh+28CxJZzFjhW8JL5NJUUkzugsE6WuM+hcp
PoezB+ChxA7zVDm+23LHbvYzDKEJCeOUICzRDX9RLQ4so+Y44n5yLQDjP8/bDT7C
5VXG+xxk+xhD/Xgmoo6goqL+NMEzuForfznI0DMxpNkynxLnUS1bVvVcdMFmZugy
SWK5f0BAiIDAVixE0BGyE9lmxwF4uW+AiJ9RIaXB1mgl/mMjKQF77davcyYn9GSy
Y7fMuexcZOZrk0aIQ1NQhitl2HdgveaTiM/IqxpNvEx+5ROND7j4tPJa6Ej0lLpP
NWZH5grurvEXEUWOlkg0UPsqBpiZN6lL2llk8tdwwXEzT0Rorm8bOSDtRGhRulnm
4Z3P5puW1WGQ1qrzb6/zpgLhGSwUbu9qbM+AvQdwjMw8ERTvdezZbyMnZWvkB2RI
bxef3PGKiS/IHZ8fO10g6CGsRdABxkTocF5qsgD8PkbGlVRl8LY1fIn1COgjiCdF
g2pcZwNzKkzTgLd349nCjLvSBRQcCrUIHNQ5dNO+sJTX023UvFm0GpuGg/YPuqo7
47PY9z/7i0hLVhXGLXLLi4refHPvoYWLjSaSgTk8tkEPvfUqxmyhx6TCTZFB6U5J
/oIEmB2TVtQO1sCUrg1Z2K0/SzQQ9j/Tibw4KY1wffUfIxX6EpibKn3ZRbrLxy/4
UKsokEWH99v1CsH8/X4EWViF9Lg91aufhbfqYrJmtVDo+8doDCiCeRfyL8NK+uVt
DofGh2F9p1xLRjsqEFSCUgcLFlLSQuMeag2ncf1lpKz8zVc/dMZd36Fw3sjpTpKf
hqrbFyUX+U7etYHOXFFFaQRysEpW8aMQ80fHqQ/4CDOXqVrRCwniPbWjrUNy1NQs
RoVjWEqyKypKYdBVpZUgKKGzeAd9MpW68EmrYTm35FH36ohWzFZyZheknTPS71Zb
TnWsh0Yrf74rpTuV5EGkg6PahJ7v3naHQxhIIEJLH9Mm9XWo6W48st4ViYasapPS
8Jj7VTdyaqLsgK9/UjxWghpytlWAHI/BHDyD5ZQYPDYo+fEltl6vxEV0Rqjpw4t2
JTf/q9b47aoDbbgDHItrjbaeSNOulSL8vricP/KL1o4UOHq3UqpjA5dwcYkoUmzA
GO4jlWICZEdKpTP5w4oRURS1kODApKcIyRjmXt2N2FiUWNXt653GVuHF02gOIBSf
QqnDxSxucLhZyQ2S223UtzXMa2LmUJrJGD5J0xIF/ELq3ST1tbHUkFV6nqY/ejD/
7ZwzBNPwML7mx/Xka0JZL+luxPHr9Z/YZ9QokmPLW8HCgXXXvuO+UHWr82EawVwO
wlWMMmeRC/tTFftlThTB/MDwuJoPkJfauvcg/zLqGmpvUGKfhixea4+3Tq8yjnLq
+bgVAaen5w8O3wRkQ79s4JwqnagPyBGd4K4JYSkTtHRrNi5IKflHXBIk+kOeA5e8
Br9O9lLGb7XuX541nB5/X5ldDyO6bOFTpo1lhHhiGAXYjIsF1TRm0n3N08FgI1nk
PT3FyhA/PA8MmxqD4WRW46CMk6p/wRjfob5eCPE/wrVel7Cp15M9TDdBTPP7lX1E
+8XMlKRLhCXbPtF+HCmE56O1D7/ACsNraDu4sYTtbN2ucdMgCL2L3g+RwPwVOszg
reezxU0K8yznygoVQQJW8x2OAE+NjUlB5o8BXa/1p7lSgRRY4l64NP+eeMdA5WOK
60RhJzJrNXhao9Bf0pco/8U7DNWe+P+SEz8AP/ekKdKONrqvK0X6231Y55Gza8gn
fZkWmHMIral+0peqTqR7dUpOFXC0cXuFB2V1zSPEEz0yTf8K/7bthO4n3MbW1BTh
PMMbI0sepZ9uiQ8MWo3h9ABRXtCRuFY1gIONbhD6vPubq3rNhCrYVN/dsO9g0KAl
6Px/lmRY+EsM8sFCwgc+SOfeb7pRwmgwD8iXfKXJsw+S9MNr+LQbOQAV3Rz359Fh
9ZjBtKJ66Knr1tIaDzLtXZmxk77zikOmi3ituVp+daCREA733vOKuOwAYJp+7NMi
eLSLBLxoJOCFpT970FrzEoAPG+z8goP7Wle1OfoEAvLggpgR7TiieWnFoHpGCnLv
B6fVcmjOKQ14daIi52aF09Higre8TcsMikDKO3cm9lrDCQG+urN439AZ0fBSrmps
cL7MxOOHRuhOMOCT9+dgLkI8Nslvh3cF57zIXjBbXkTktEDWYSi5FgCUzhKmopu3
FE5nIhw3vyjb/3HEpAd56Fu9akoKxvOk435icumdVLgVGTWYe8sVAcOsKgCc/pn+
K5cyO0PH8ZeCgSnu/rPnN5kRqiDaXNcEO9d2YuLhwv/eq4bjvZ53urg/0ov7Wd98
gXDz7+RGX/G5NEK9WjC9UhOwKn2kX/y5dozPfs4eaexSCPcauyAhV9pmwxsRt2/b
mkOyN9xgkn+X5+XeJKs10+OPuevW56p5h3z8zfK7m4GLS1LUMo+sIHsjmqmSUDO6
9t8armwQpbh8nK8TwTrby9mCip7zv7heKkbc7+IMn6yvv/kT82QjnDPkDvWopck2
kc4ptbYWpWaW4/qxjbAwAEhWXgg/YU3sjHKoB8CiP8lJFcKBgrbXr67EFxkjQLVG
VyOf2hjbQbnTAlBAEtvE5WTNYsGvCejgtcL4Hq2gknPE4AL6nIFYn5FcPY+Ytm6q
NXrnLJ+dP+VRvu6bdluI8a2TBZFyg4jgJmM8i7LIJ92RQ7r7lXuKbsbGvbS0KwWj
wrMtIZDd4CYjKBBizanxzsK6aNf7aFV7tlowGg2GUrXl4LUEsT2I8K6jw20Yklel
szJFouD7jrCfmjeSNqVIqEUfTW+dMirZLTRNMciWzs0DRj65lkAKRnQdpx0CYZZk
gLjTLV/EhDwnnCDoNPnkCvVRU+TJ03aITgLm0gTsTVLALvxnjloIvH3MFRPVe5bT
MlNNkoQ/jQH7gw5R+Db7Ape3Q0DX8K3960GzvvFKRNpuS/rDWMufF/61UGwhflF2
8J7/yegS4j0fQz7kayVdZKh0lgN5A6mU9W0ROsg3fK7Xaml0pNepYzMjwMXqUqkc
SaaB1U7MsyBIA+mb4B8oLdCXrMReEAxOTJjarI2ZeVx8hjEgGkAuuswccZE+OHAV
PbvwLKrzsMEavn/T1aT4+RQ4s11REmX/vrt+hI0XTNfcRvOdPBWzxJB6ij9X2P9i
wS3/hrfs67otyqJEmSsz05Zu+18vs+2ktmhAhRP0iapI+2/PSsaO6jv1dm0YMdOH
Dqb5aG5sMqFrBC3ir1JaCSHc9lXSCSCsCFa2vNCDzfPN0KdKhGMoD7XDPkP8oot8
/ez8wrsMmQdKfPlyO4J3E4vGr/ybBs7UmSnaSOELD9+nXs8dQYoBtivL7DDlgZsa
NbKVcpzi/BIgZ4dRd63RwSI7sUDK43kHqB9DoM9aYgN9nFxO4O+Jqwb2KiQFiAzw
+Y4+Az8eskYQEVTimpOmHpki9+OeJRINoeSu5aOxwu8ceHu5Wo4ld/qFmFTWUsyM
a0Mk3EdBg/23VhSfPxw5nUIcviOvCcD/dr6GBZ1+M3Y6khy7m6XrJZmxBtc3eVpF
kXS71/qpvKo1kwkZfY0km+tkhm+qCLTlEeaJid0+B8SXb52a6gTuXNvtojVFt5Xs
BB9WUqxSm3XM5fdED5EPFVs+XBdW99m1A8JBPBBA9JLd5Pm/AzUHNF2WXHRx11K3
2Zz1vBxjST2CkcCd/I8C0zzLDPm+L+wBmSun6MbGcvQbDDAD+tEllgLKRqK5FIUN
s8zAisgI4BNOC5duMr9DQH2r4Wfh6zF2NSRmmPFRXNFGJFkwgVr3wBE6WLzbWWge
a4BAfJ4aXzC1E9hjCLHvFJ73uMe05gkIiVBrkkVuipsRZPCPuro5FloNOa6anqK0
Tz3XYS5Vpm08c+vaq+ZXSV9E5dKwwLIjHmpWpKXsU0rjPgyxBZUPWe948bCNeCyn
4v3kkla/njjIt5jCgMTERGT1FpQ9mPU9dY8zYuV7Jk8Qhdc/iSJfMgTi9kEKzHiG
RDr6nFNZgQUFWmVonhlQQhI+9Oq1sggFkHm1F941NvTXdEAAblKKEwxcp+rgdNFL
GC5iK36iPntrv3QUG3+DijCcv92Ic0eyF6RHlxU3lKrN+w6GDI2Hk6Vo5eePUDNE
p9bqL2isUbhtJdU9xTT5EsE6xttZZaYRObhC6TQJ/nSHNtV9vjrJsFTKLAa2FPUO
J4GB4Y6C+JQqEQPFnDc4WZZhQSUF7cXqCiORaI3VdtkghlupyMT9NQA5+RLoxqdU
4KAZTIDOgitsNBbIf/Y4httZJF1/AFw6Oin2BhMLn9p3q+oCrzp39sJdckCuG0OG
n2nGHJVfVvjP8Bb42/h1ydSKMg48Nf30O2vwPmwjuKqEt9a+Iv/shw+BOCqXDjPb
ZQZVyw6h9vSOnpCORjzV0zU6y6RuUFglrYgnQrkMGN4hlXmYOzEXz10CRseoc55b
XazJCZmH801PTjcD1kyMTIyV53Aden5p+zkwnaQ7rteJIeNbXH/MWqRJ1GLSnnNU
+bfy9nK4ak+Rbs44NEQ2qmUO5+GCIdcOoGbnXWk2li+XpaPdWzzue7BYGTz3VJLN
lrxN63sxW6ldI9H0O5rzTAH8ENXj4FCBQzlXoVjdXIJHn8MONwZpMbrfJplhwV3g
dl5wQikDmJGBQkcWCuq/eTQcesenPgT0h6ce4uigkNxfF9N5Jqd4o9CWAluZlEhk
xqA1eNcQmwhq7SckyX1l27VRRI4s0eRgnjlZG3eDWEM3jp+ODdT3rY5kPfeeM302
FPQAznP6oFzRHOqAaWVFKiGWsM4HPNdsEvpFL9nNd1C11PY5CqHvzLuwQtXk056k
flR9+hwfu6vJK3JUrZ2uBNhqxg3Jp/0VEOdwM8WL7xfultpS9fhBES9BUppuW0mz
CwBtuSk17mKVI5xZL8FvStfUSDf7GEziq8vCQ3BOVHs0lSzanBRIr629KAQvfJjd
PQU1k5ImAdjsczNRO1hS8puyG2YNMnEGrVEIuQItdOerZOSvvdUCiJIltu3XUEdO
cy6qtc1VmwPiPdAEH+lxTrVypDKoGweU2i6T5XTpSCrLwCN5S5dL+TpUFmoeRANn
HsXLmWq98HlPX93427ay+BZYdqzOER6sGA4FNqHnVw39ZA+cGFYuwGz5j3bBzxX1
eIOsN0KbwM3+fgFnj0CeDEJHVq7AHv7rz6eQlq6oYnrn4S5kKXdSWSnT5ZO+Cf2Z
oDWwKJ9TsyLkn9gjjzyVIzu7o/RHRmZ1C5ZuSvGtpNBjmDi8APKwuqOZZzvEGPkW
o/6WfrkMnRkKjh2IedBDgNVI9HicBnHiC6ttsBCDPRXEmjXjub7baB900VG7COQI
QWpZNQUrKHrjZJBvieBr3peBCGd/tCPIcQUVyUY2s+fMte89vaxG4Y8AMGNfSi02
Dn7yNQ8K3p5d6qKLkNvmGtZ27MjI84M49V8uIo5NrBMjKQWhQnIbaKKrNGxi0RCq
69kxTwG/3LkRrlcRUIbHs8cVIUgktHjF3EUe4qxjPhIk1W9zZ3EJVnaNNc0OLuF0
G0MYXB42fGD7THKMHuZHAk8W08qCuGsCniMzYSysRnNxNmwCCzglkcaJOxui2i/H
ObYkjgvpSi62EkZ+n7i2xaLLDPLcvdyg6Wu274Y7qOG7vacUhugugmt/Spn/JVPZ
/jmXeE/HLk9DuHUg9rMtXPxbDN8jDHBWez3kro7C7cOIfrhq5ICm4mpe8uccE0MF
/939+soeW+qkcDiAtzaBs7tIIJpXAgXoqUKPdPOrqjvfKiw2/ump5OEIH3EL2wBL
mv/fMK7rlzK9n6I4Lz1OgN4JMEHqqoPxqGu1G/Y6q/7Yo1hxiSEohQ4ThsH3jMW3
S+SXXpY1FocwNaQh65bzUoWOJwSHvhwXSYzzEL7RsqYEv81vGpVyCPKEQ0fcam2C
UTp+BrSk3sYqv2f6Q61hZ0wXSsUHAcG8JODo1hvj+dnQmk+TXAq912OswGRNxpE9
hP/ReYuG3+KanTyQyhWoFsDgr4ECNhv0JfVkZvorYlw5TnQzPa97uj4Sheyjq+W+
J2kETHVAQBwFCRHr9A8uiS8fdMN1WGngvGJHUiA+TV6kGzZbiBezU7EeYRSLKIB4
xko4kfLHNmXIQxlmg5wZCTiOUyCS8+9MGnWh/nufCvgb22PXuNGzOLXHeR6Nd3oX
DAiKsvYQJJFtw33NLo3ySKmZBvN4rqOKC3aOjVHUowVpMYSK7kkawoe2EVeGIp2M
eFUEcxjEHbcTw4HVpoAOut0LLUTa4OmZpDuGHKjtArVNDz4DZSbkmNVxR5g6sr9M
6P9QLByJHdXCTDKJMrye29gjGt6+RgYGSTKLQADsClMELfKTJSjaMYLKTcJwdMaE
CKLnuDYdrboVufvp4ZDj2SGP1hcn0rpJs8C+3dR9G+0VlFYwiknv+D0ebIeaXCtO
6YSLF7jYNSCbbGlFSWku5H3tNVAUAWZjbSFD9EOQ2D2orV0Kk8okV5TS7U/4PoH8
AK/crxMPimOTOER5OYg3K01r3uxA4ZUvE0Rf5Z2wvHr36FOT2YiIaf8yhsk32cdd
3qRci3InENPbKE87VSJnNaPpXZXG4m3M4r1q+kZLx/IKSJne/OmDJ5SMhokzpAr9
XYDeEQuyPmVgTBpYRw3IURhrSpYYqKZSqBp82vFDDXekniUhKME2UHD7UA/zdYtI
NFd/wAG4jeoD4/PvbEqPJB0NMz8rA+E10pJ+oN20JPcvZV96n6FLzjAj1WtCbtFY
Mo3f2mn6N9OKULdCqOJNwWrP1gygRV2cE80MUKqEf0Am7237ecitFm4g0lJGL1kB
kTRZeVzbatQtX09IZ5ugkLQqhzr+0jxmdR74WruxbcxXlIa3qROJ2A99G3SgL1q7
HMJxAr4wOsrHaSQISqTM2vzgvE18Y7xB7H5+16bnKWqm7MJRLot0Y4NKR+PyGkaH
0ybZ86hksQERNXGCQ6PkSpmS/0hUC4hEy7RTfndsLCxEx3IArgl+e8YlZkJvOraq
aQjOI/Z4wYcQhmbU9T3ALRDAKQsnKIXMhQtJCh6szhmuKVQFaF2Tyd6dJnMuZJB1
5eZMQp+1wb4PAQQYDc+5XOlLj0a995O2UJJG80jQnUPDWCXfNvRZs/33AguBmkLQ
JbKSNhaX6P5qrpfF/ziIm1pA5TaI5tGje1m0Doi8IyWMS5Q4c0G5CUZXrQJ6OIkF
N4uoSyYhP0RZpIxyE6EWqDSQh/aJS2Gdtmcbzkc9ihKmTIaY03Humnm+e/oz7Kft
VX3HUCbCLKSeu179Da1dMZ4wd4tvGItgbRqS1qY6Wcb+VOCprW1lx0AuS5S33p03
SqStrFIy+vryicOHRGjBI2vqPFrDGWXZSKX1Gz380b1U7NzZj9tXS4CTcyShXfTO
aTkmRLaP1WjpbsHeVk8FL4z4eElxVg1oFUhMaLC9ieBIsrNyxAhZlUuwJV9h6OQD
3w4sk6zBIGwlUmL+Dpv1rOqFO6fFAcQ5NDXYxTajXPDItOp8tdiHimKGj1xxn/Zn
EfShTLaozaXEVMrdKHDWxr9B0H64TqOQmHzB/vCmWWBgQdoEyFAGI5y5ML1GJBgs
Yn7G8y81RFl6T9xNd7zU50kOGas1wIbTmbQuTRVqnc0m5aLPnvptWYRSpi9h0nb8
XrXJkoozNZjTkcMhYJTtrI/e2zSU0CG4psk8dSRTptPpAV2BNuBjcZ75LkWK9Ka5
SdVqxHBEx/gDj0xZ0Jt8kQkJl6RhQyTkeFsVtcD6M05JfTHviv65CgQ7Pol2ppEg
zt725tr54txbUSDFRXPmrYbiqx2r/eXtmlFxAn4VkTC85k88Ck7Pzo6VN3EZvHX1
4MoEHyT9NgMW6xZIySzO5uKDJBdf883I393w636nsQ62Xjycr7NtMiKweqInHq9J
HOIv1lCGaGA/MLZzkp49kl3NdGoxHGwzwa4XXOCuQ7X0btMuoFsfLcqvv6a7YOKZ
p9EVS9Higf3Ss3ugQX3Gleq7JTkX1/FZHMsgjQQF4S83tjl/XaRnu0pU1IdFW6zm
+2rCvP3QTG9lGjozE7OTlOGcBtV+9Zic1LoGUs5UqR7BGW/T87VZ0OJCfpL8mvrK
UiV4VWtESinsTjHIhVXEIWYmsgyOYCGNWHuetZhBYDUfMyYO2BY9gVyClYIUfjn4
fD4XkBO6vNpd1zgj384PYWdZzlpco7eQX6JxJbS88l7auLayOS/WxHAPke3hdvGo
QzScSxQAa001PgtoBO2DdzUO7vl8XFca/P6r2hI0Uhf9QyuXhA2EFyADGG7TfU3l
mRPB4YJDQ0aZJT0vyt4+PVYOUQK19tNSZck13lrPz+wIMPknyXaJN8LvlL1DvyW1
G/CxI6oXnbxv2nqINuWjxX7/DGGIIavbXJzO0n+uTELa7lDWhi1qYZcaVJKnEV9Z
tsPtcLpuR9hF9qA1ZaCO5kuKDO0P8LW3Jo5IsAr3r5sBJi2i9heWKHWtezJbUTmv
1T6A+Gn0X1M2/iiejvmCleTEuO8USVkpSW77bXMfFadVtnb0JzfdxVqCcWz6b2+t
Ck026eBZHj6dsRLZblof2Pune+f/O5PZfAdBHAcyfkDDgqQ4oRawWXzEt4fgpBur
waNcT/3lgMVre+qDF+q9AsKPpfH+PWl0h/RUFoVIFt9nr1vaRO6stSRFeNaIuTMN
xCGpNcX/f6ONfLgrdT1nG5wiW4o8oeane5GkKBRi3XtOj+6jwq2a34ayhd8VMV83
vKNidm/iPmF9funiWmO7ObqQ+M05220nIEWE+C6x1/S+cFLCnkGbMr95gNI9QXJP
d5KNPk7j50gLH7ufYreWEgw/143aBY6A/fJUAhMpQOcklt/3WA5wkT61imoMT6h1
+rFY5tJDb9y4BLVzLPDR+MBNQfmH/VZJz0cvlaYDEj/rzoTBkb2x5BGwRKkV1vwJ
3jsVkeD+nyJO7WohiBN2WmUg63can+KoAVLPPwgDoUWt+9xh6Bz/a3jwf1F4NLqG
PP56iUuQNtn6DpTGmAhVwQFIjB4A4CDb1uKhv7makIWOiqMNzbJPJg+Ig9Kf/7pb
XWKrcbBwferxOQW5ps0bqa9V5wOe2d/Elg7N47nTthSmTliY2E8VyIeYyRK1OEl3
sBUdULJKAGnWd+uYiGSwGe0ukjaGPREBcg5Fg+uiPPARoCk6jeYryv18v935VA/7
TFiYxSvIMogmkGNDrOw6KQgHxJcXUj9xToIiwV++gjUeXPiSXFZfWNXGQ0gHbpEX
lqcdrRuaWKdQmtTNAeJ8sCygy5rjv/vlW690PKjhXNn/2Zub06049zps0UlIyFWz
6pcFR4D99whm+DaUeCnsz18lhsAy/jQP5lrbZghjGRbMGlArl0BzgtWCG2d1EYYQ
bB6RqLume10ccMWHDLueV6viPcM+wYKfzt4aePz0fRhS6ePKpPPi4am0OoKsyq0c
2vGTzxhZvW+Znjah3ZXBnRWq1PneWFjbQg8Ly5VEN0NDPIP+Cpn8UEuIhTujfsTP
u0rT2Zftuc5ToTsR9ZxoDOLO7g4xb53iar8pitJOBB6CZJG/pKNMh5yjWME+Vwnd
7GWY8Ze/Ss1txluGVEa+HTjCty0VnSALGaRNSZZh62CB2llomc1ifiFIoeJqqp5l
mplUiN01kBbDWfyyNZB2vlEY+j5cADoHowUD8938RwLuJkeR3mx3xFvvq2Q79XXf
yXCnlmNbJT5S6z71iy61KYU6T2i/zuCpdSBHeo/HOkS2dxL+4jC2+WDdyyr/3oc5
mSJcuBa++X3iB6yMW4U0mntnEc0suuWyttqSO0U3MUfXx/6OqCXbTlVDHVj+8rBo
oChU5fnP4ya3asIsnT6AYaxsZppUUbVZC74ZEClGuVm0HR2dxtiB1vwwtRP5xbWm
SSf3WYPdpbzgPq3cqmbE3JS5knx1Ca7sJ3t1oSrcKZDnge9941LByEVshegiNLXi
/RSj2fszD3xktRVHi1EI/moSQ9wFzjjyauQDDuN8gwqHage7DvJzAj05XrfsQD6u
4Foow0vLAjC3TrAKi+lqHeAUyY7KmSppks3buWlw7AuyZ0bLVKiH0SkySqCYoge/
StSvwu5f/yIoCgCuSwuyATBibi4Om9jLQok3dENcFINgXG8VP38EaoKHLNlluN+t
2ZL55WrR7U/tFqcKbGOKN1MV3ouExxN3daRMYTnUsulxZjTAUgoLtrUjrv9r7bcw
KrTMBqtAYwwaBVFlBGHSsDvA47Q1+3vcpTNdeBu6BkRdj0fmzFh1mSytRep4K4Rh
KDwqspUQ4NYcy/UVRjbvG7Xh4+K7w/TSMxmLboU6+6XNbJriSlIn7710IgQZySAq
bs4in5al9qXNiF33Oslsj/iaVFudCPWFSi3Bf2eynPh5w64JQK6oEvsl3pX9V86w
Nl1G1UmOwk1iRyqwJfxDAqtNlpEty3QBIDY8WD4DQc9wb3wlsjBvaQvjFcDRvi5J
LG6Go4kQMhngbjEuX//vGezzVV4Guj3GJa8P+U6ybu1Iid2p8kf1RaqWuZS8e4OE
eEraFeMaw9/0zzdccknRkHz84faQIhiXLJSjaku33H5+wcYAevYbUR46XoProMyQ
cTOCJOpDd8vT0AhwJ1ziyxMfyVQMI8gDbo1+SP4UEyJQ65RPWsWoyYXMJPDs+7ln
Y6PDkw3wvo3cLL6sanQsvPkP8VBZsEYZpJAig3KLVTtIkr15BZmQmF5JFOknbzRz
j3sVCrErGYhdFOVGZQk3DLqUQJ7PO1VmNuQKS3wyeteld1yrDKjP+n6QwQI3BzQ+
WjyAAp1ad7Auk3l8qds3v9Q4/OwlRTP8LOv83DpkzKSdGTg0OG4M/+eFhun2rvXF
KQLYtmcEsYmCkkIrLQ/wSDGlnIwjQMHnzatGLqlkjXchMBcT0Bz29kxYFZXegmTG
hefZCioGz8fxoMMM48JiJiTwhEoFlc7fQJmMwlaaRuEiqRWFrXnoU7l/3fjZQsEA
iDuaWFR/fRLMJVxgyxr/1JwkfWEKiAUA//ElVp46GLQ5zlCbo2N3nvUAuQYdHmuu
0KMHUAnXEzsw9cBOuQ7VXCcMwr2KKhJcYw4kvs54uf6S7pdBG2/sb6GvRIftb9Fa
ZI9wUpgjnE1Dhd4cb0D0mfK1Jh2cASJp8P1jyOcHqeSWUDppJ5A7X9bAHrIUJIHJ
eomtiCRuaplkokjuBeFe6iSNDO2voxSKYVZsrggkhNLmiREpr9+m4VHy/AKQNVen
oil5PJI7vzfsovG7TepG0oEfEiARepIuF4J9xQdltKNhmd5Ps4oWh/i2ET0ITbfI
1DsNxdm0H1arfGQguNLpmM4LzkpAFjg5lg8VMMPY0X0tRvESuHxDkhLaD02+rJSI
La3BRred9BIcZqzcN3OSygnRPDqJzB7pNjYKcd5DTXiLdoFEoARx++5ZJS3edhlM
9tMz/G+0chajJaQkxa8dwUICCg6W22eEwwBROP1rN1gjjK6+g/Yaf9ZYnwFyj/lX
PCxAiHsIfygYju0ug3cCFVSVBnffk4WSiB60Lb9HIUjnidnqX5NJQSQkxfRXdjaC
ZqAbTMrEOHX/+EoHrMGNwfechFZhamWHkKASTHKIT4hC0/1aY/2zec6pYeUBYLcC
2oIb1vmudU8kjDVQ29sWFZlAOLRrp0Iq12Tzp3aImiZds2+E50O7MwVXyfBVfc0Y
8/YBp6xjdivR5sgh245PZCBSphYsdExwTOu2cbUFI+c+HMPvIWGfFdPc3SHD22u5
43pU7e+o4N7R4TXqnNE8YyE1IAlIuWOVZUJffgHf483IaKpcoynZoVHrWvKAAyEB
C76WKXVZqubwEPPpraEq/4dJuKiKrp7mvAWbeA036v3ToZtJU4Dzw32NSVSV63Hs
pohcjGT/I1Ghf5xhysaX/vnx+/gGkcgVbJBOvMEpah34JLG2QQFa5ODIurkk6bA1
JIHf7qWLkTBgY07FtVOsGidX1RM4xhUFL/MIzYxF0SKzLdZe10GOAwirGOmp9i2c
D2lMpQk3uKd46TZdLms4Z95rP2W91dUnRHSxPj/qPGA/QT0U3fvU0C3z41VXJzP7
f1AxXh2OM0g1qUG2K/T9yV3crXEqqsa2tf9n9e1P2VDUIdvX+DQjSLwNYuGOh6Z1
fk4KQx6Pmbc4FYhr/SKdfadWTAya83cAe2rLL8Tubba5/kCloGU5D2deKiiwQygs
tdA/fMhuczLKuqVxjBQEm70iITnJ4xv3aVmFe6b/ZLpIfGQ33LwumN+MJtSoSWta
IxQX2AHVvcDCrsoCzwVz4Wc4lDYsUSgdvxd0OoqP9M/274jAGrVMfvJYuU1i0i+I
TkoFV2FmDIEGEAGWueKx8TukCMXTiAnLPkrwSKdsi7qFO71X+4G/2Vi3+zbMX5jg
nAKcot2VrT2pRM7wzlsowZecyydA5UHXLPCu9179108hV5q9wpt3tUl7kOh97YD0
sv1d0D9gGqBsmpr2c1qxsIvfC+Cjefbk7ro1sSAMPyG7/Us8EwktvdvS4aeFvI26
6/ddXxvKxXpHDe8elQjqw3gXHpOGNvqAyiQahFAJwm0ZJM/hlc45SE0ayYvfCwbm
/33+DHFaRE4da9Pvxlv6bBllaZ5hH44YlvqWh7al08SEXInf6chCV7F0dDNJGCFa
6K00Oryywj6Kt2kJxSa+k+l7g4d+kNqZkHjfA8FD+R1km8z5vHITiSBDEgXsU/l7
VzBRoSkkRE1dyMMxgCKfZgP6OJ2yeWMlFwN1yPDy51whSGTtU8dC5lzPUVT8Qne+
/LGtDLnvxV5+AE47xFM/WzmX2TIWZL+REKZ4CL477iK2UQoe6U2Qsn9cWHBEC/Xf
zMKVV3ij6WEuGrmIRx6CGWm1ryW3Fv2GSJNod+BBhwbdhJy1yCa/nL3hBAmlcRQc
cpwELE5hn1Ndg6lLpqCLvga0bWdR9VO7jagwhFFTu5KNEpgvYQG70FnlxYfCQwZ/
Btqj/XCDCpYSs0JPmR1qNsZ7dgfEnh5B/23lvR9eUDX4MqKfPtCSc2kh8aNWxSsP
dqvIwo1k5tt2BJxs0qxANhOHQbEDKXBs8SovZvThiC/YJWLp8oWyUUzHiZrxyl6d
OGyPVPEInSfUdX1av/wdflo31GWpgDKI2K16xFAPAaX4cTFwxdUlJiCEoKetYRfq
BxCxADLcp+gHOsfd7MhQ+ayMNLE3A0bNwHQChbdA8GZnRJGnN25cHJd8klBE32pf
sh1kJ7Yway3bmUEUdGRYIxZDzkFZ9hoFw55u4uEix3Bt1BlCYQR0uSVDDDP9TbVa
UqqD7ylq8NhUUnSAM5lE63egXUAHduSNKzkdNkvzLdgpfGA6rln3Wvb3OeX2Gk3K
Y1f06zTfxro8Az/B9Sz4oppakif+AFXs1U8MMjiT3B2nXyOTZjn1rUBqJgLZiTcD
Jcl+1GYKcXI5Npoq04xrec3HpkkkmiflHmqPy9IC+3z+HITyJS2ZblwS7ZuzRczt
Ph7b1GBR/M1Nr1S8fp0mlde/uPRplOJSUEu/ON+gU+R3s28bLyLajE6O+DMg1Hn/
HW98iVwh0Pz9ATFl5780lMi8Uyd8M2UEHmjbqIG6kQ9m1dAhNV3YXQ34VHTo8NOn
he41zHp03DlwFokEW1N1plrYopjeG4tpkbF8Hv5N1RIycCeEdHFt07gxSuynBKez
tdznYf7oz5R6l71ti/Rp6RNHPdE2Jg3FJPZK3Ib20apSzQR82Dnt7fAbi+Le75BI
FC4HxCZqvy3bZwBfubThfoWIAAVmD87tWv17oDPhbI7LOdlvjcwtJ/p9FUDqAMje
TcYFWFw5YoRk2yrPNfZcztnoG6AZMRfa9kpNI6IhGLL325OF//eYUXH4rmdkh1dP
uclqfGVtSZw3uPQvQRmpJ8zylYFxmTvZWhsqFBB5ZW/SGrHg0rZLcRO4V1D4YhTo
0FHvrqtVRub+Mb+JazGbp+4hCZS7wAb8OW7/Ekm+afeoAUDY51z+V3an0Jz3LFcD
kQOg4lSGcMa4yLtJiLhnX1hiqJuKslJTIjqZNx/fWY+wpmGJxANDsYDCyD5Uuev+
DEauHDuKFmM9QJWSUjeKtCzetwBv9eUFh4Q7k0QPluFBrGZSjKycJfNZ1Fh9Sp1a
u238qShOTsXhT+/cxZ0SzEBco15k/G/ByLoQ2VHAesV2+3D06+mFfYLavsZ5wMwa
bFU9EW9UOR1XpxVm8D24sN017BrcGShi7/lfQOPZPnhnaj9uOHOb6pyowKd+Cm4+
1PnSTs9vvYmsdf7wBNZLxndL8fVJtroxd8oRUr9W/KUVHH2pUspFfEU1BW27B+d1
YlqLI8bIeo45CwEX/eo1/Kis5ACRVl+j0fTULT7O/U7i2rE6NuKmycR+3xM1XSll
CxAJsR30fS2atTnv3+oyroY+dDuB0gexOc0b8T96JQwz7bm/cwoUHA0UQ85ooKiW
RSH2ohI5Ol2IwdedWk1cTQ1JidU2vAW2RGlPrpxF0DE74Z7ULy+lJrqz63S8sJ4f
pGX/OQXa961L0ZUzIJDaJkEzt7cvblf/PggDZ2XKkwTpQQ5VS4cSR1mKzue0IB0u
+sK+TEurwSHA7jiku/W54floiUZg9/jPoIW9f/udGc/Ku3eTQ0NCHKSIc3GUFvfY
02j9Qz0j4nV6QBJiVqIu2SetHeoBMUJRjjwwb3sgpBHJEddOPRNradDNT+cTdYKT
1iUXCfpVe8HvDZnK2SmKTtorv/onccyYJpmRverIjWmp61ORcUrzecN1kWbbZ8aO
q6y0DvJcyRS448tuxlDI06DjRFNfVsdXTUPRZgRxpe7lTvdOaAZs5T9BQ7CBsnbK
4oZBEY3aUhuDYBoqZ0fma8sWXl68IC6VDZHYPQoznvBkpAIiTd7qSKtLZc6Rtl/k
rdxIhBwpnv08zSMOqTuGjuV04lJ2L207bYiOeQ9GrGqHSOfZiyuMlXpr92X9HC6w
dMUwpxRgy+opfUFR96wX3cdovYZoB55t8VPR4yjoPAAIHz8OFgHT0LWw9oljMLW9
Y3c29EWCpLYgl2bN6R1/3fqYceoJSETpa/WE8i3CweY/T57We+WCylNLlg6YrBDu
kZxy8U7WV0FSaOjmutYLZavxVndsUjFAD96Top2GbcEW73tr2RDb7ggO9E7Lc4sP
rtw1ntfVII/mwI1K2atGM8gyqRmKh+rCm1dySJQDKbiXhbxZH+EW+FvOxzgGhBgt
ye7Ul+pdTqA2vsQXRsKz6XRkpBKLb4KLaFre2xADslS8UpsjO/S1CiRLelPVfh9g
pTArMdioaTHktNsUWcxle1TIFAmJr5+5lm1peBR+QqdOUV7IOfzUfgyeiUsaS4rn
GVixi8MfHZK615KLEsiMDVou734+yhf78X2HmnBAOIImHBJvbIVCZQ33PyevTigQ
5MPkpdKosPO/q1t3+uBEwogiy8KJKcWj44gk20hp1WashGU893yMsRo9zcFf0/2I
Kme/2NIG9CbtEQeWiqj7Hdc3anjivrKwysSyys6rv/ecwmDGCBju6Rg9kmswCjEE
kGgnmhB1aPSsvTyZ+m4bt3Dx+fOpaw0uk+lLjojcBePJVcm3I6/0h1Ni0+wcoEVe
nrbMvtoiJJGFkgXKRwR2GVadktU0aJKQ4ANgRieYsPX4IMRWoTdj2BYPM6WfWNNL
bxQgvLZRmQJ96TSGAcVOeflO/p2OpM+Vfn5ALarZ0xS7TXbkSlkf1lxurzIMhvTj
N8JNp6sMY55JVlB2VCa7Xbtq+tBMidkycDKJqgyGTQ0vHOzQRMd73jZzeAaIkA6I
AyFUrP51+OBFq5FNbelt9YXqZB+rLujjwIp601K+a+L+fmrRtWuBkwBNmh1BN314
yxP/MHEDqgpLAtTiaxeb4FKMXuRnc6RT6OcMxjdwVJNlJN6NSn9Fkg98+lnoLhi7
pUvDCGM4kDDWPX5e0J+9Y9G7cl8hJdY9JSjGc0SPV60mpVe3HmKT9bYjanOtezH1
isZMpOADNzXVz2naSh4GXnuhBpO1kyHsG0zlB/2AguRiRvwy5CEwp2l3pnHx35K3
0W1BRIxJ+7OKpLErqn4NgeEYNNsUYQ7pR5xKixTbdoeCS5Sl3ftenHnsUNxw5kLP
7AYnnTcJBHQdZevXG7sn2hbvao/H57ftgHJefHdL1Oxzjo8hD5X54IZjs+IZSCry
d3lBWdoYHDWMsW/ufjP06t6KzUfYm3/dVy7W0ACZLkF7W2bQCpCE/796mAbkJUev
TP76RMVvEkYqOl4V3wA9Gh3Z2bxRZv3iRr6prJPYLcs77ZRrT7fLx/HmwNdYAC9h
xtI9oZvH/rZuV3sxwd2l+VjzLNHJ8e1cCygvdgwVi1UnQP6Btkcw7zt4WQ+HgKOI
IVs6dmZVcM6N/CQGpr9gwwh70RjvmKovzZRvXzoggPsoDR4poJ326Dw9FfKb71Yg
rCG3VmqV+rKwgu4UWQhNmcbg2zkG6hUajE7sBGGfuolpZr3VNtmy4StkHUKE4F69
Y9uARkkfybM5l8fNIcqtBsF0ajFiwDYvMciqo714l0FdukuGJYKqVYmZSP3hOcP5
hxWjHb6tF+BSI+7Pus9iYGG/HfQUf3a78Dx8ebcttdURFknI7cRl/FOiamiXxu96
G0+2Lo04ul4/+Ru6NCf0i7ICsgM5GwtZFR+CxadLrWQvVhoMjQduqcDh1wGpzdHs
1nd5FTx67rcukk9l7MnTD7aqd9H1bt521uI2sZu9yPRnNQ1b3wzc5OyUzSD/tt6y
R7yWOvA7KTbvBM34vlJcUFZA5pvOaAQ0P056+h3pam0xUgK6zbcMPeRbvp1RXnq0
UYl9QtyjFamIsGdbp+pDM+5X1xiWeni0vN8sACNmnLCyTv8EdeVi19TZMewEmrqB
bM5wMA3qZXTt1+rDbemjbvIX3MJap/u1WqJmkBTbN2dYujjaw1hNLZnE87yvaCUr
3wl1Y5kWqbJviaMHpA1oj2HoTCGYjijllA9eTiJKx8/dOxZtVhYULehYJOmjaXqM
bNKpdULgDK8+IVgfJzT5TB7TuZ6cAmwiWXgS3sTAFdYEkBw4kQq0tXkpaZOobBxh
26Mw4Q3mrsc8GWrB6eapNaOgvb2ogSJUx/CVgZJ2ZsTCBhlB13v9o/PslGIDhdhM
4hh+4lHOSidMyzxw1s0I3uADCUqmTUy4HMZKWEl33SRGnINuFOOAiVDtPTVxZqcY
afoyYhZtS58QywzmzMS4pf4daPbg+Xooc78GfrkvzHyW7JaXJKSXJ7Wbb+wz6Y++
awCQcADozi1CR+rsnbJX7RJ49IFfqH9ASM4dlKM5JndnUUH0c3l8K4dJNzrEm66b
F9r4JPX1yfmlAYvvBk3R9BQQe6cQ1qVlAnMvUXfSPvrWjMJw7xzNwSl7rUho9rWf
pS4hG/5xzo97IEg8eZ+qskhgdMEHm2/bBCm6p9nUL8iAh8ul+RG3hA5Tiysdo7zA
TbcBhjKVQxdGNKfKWW0Mm480s9DH/gAWArYCsp4HYhggHBJsui+9Ao7wFQvGTVDl
+Enm2kP6awq/kfLWqSieeHWmjabaEBY7jIcicTCchWjEm5n8B9FjgKrgCjob/JJM
ipzLIzxwJ4CWFrJBkkfTIdUN+oz0xrH6B4AQs6pVQM7j8RkQXpmdUhSz5HZPsKcF
0neDRMIr4zjJVEFShsz9TKG7ln76IOA19PL02KSkWlr9cAE7+8KCi1n0+SoYoaB0
z/gT77TPCaIs9cP8t8Nc6xrjBLO2qgN7tLTlxWZ4F8+2cRizlYdXhaq5svmkcBgq
T6iGQPDvhXEoQNZy+VYmWkKbmFQXfbijfGxaYi+cFryVdbPmLLEnbTSwtB5D1WOb
1lvNLl7R9XCfoFN+AwyqdgGcIlaaC5QZLNUHWS1wxSofyPIXOFeM5VORGdXBMsMa
K1CPXn5e3i9ZsEM1Z9cwUSlGKZl1/PwhOlqdngbTTAmjMvoP2V6S58RVknyzAPwy
Hxkw/5Miq7+I28R0fEsR0Ggf8Mu3vcd3El5YAWsNEeV+gbnBkhTVgvekfffNvJ+X
p0UHWzkdoFfoTK3pLrZps+JVBs/oMduOyJF3dckyOhv7F5DpJ2CS5Rh7cvdvxjEK
Ogu38Y3XIRlqxuIOf8Ns6dKQjajbQw3juGp3VRAOpv6RI0GLn/G4dt/RQA2RfNtE
ctDm5G/yhOrm9xMGehUcA+0Ot49psjLBuY6wZ9xpYOuJHGBWRxB0LW7IWvfRIPQv
5nqjqYXtOoBOcW+MYWLdIihTpm0Crouu1ZQFJ7qVzD95LjO7EGyEbVc7hN4E9ACx
sCADvkx87Q4efV4vxxsi8kxevdaQgDjFVp3XnjqpXAlva+6n88mwhYqrGhFhK7ee
JfZJixlqdQtDZKesmxVvBnS1ea/63FbNwDFo6yx2JRj+5Qq0tJLO3kp1AS57N3SG
ic8mdHcaCjh/iCI8KRURf4Bc0Oqq7DjHps6VCdXJ7jiEo3mVswRToJMn9z9k1KZy
NFhaIjKXhwM/DscU1TjcZgRlcJaXVIda49XBE7tPYq+UEc1p8c9qfUV96ggJbevM
uzvBpXA+BXlM/GASawX3xsXvjPP4knMtoX9WOLkYhkbOTEIjEX20gdfC///gEvCd
FMwDmefZRn6duMoNYH8SCiksMh73ioWLtAx6CFFtem3PFnl+ta4hknl0WCbmQSry
fvLIbAfMawkymIjl5ii8aTCYOKBUZkdGasTZzDc91ZGS1xbpqiq9dQ8aPPUDI4lg
VJZb5MeC7/nzgCM/IbMbyrYzNMKrsARsB7kYuKKRhd//KrPxO1+VytYpgjPSVS/U
CHNXPqn+myxQ8sUcJi/VzCGYfD7CI6HcOKm699/ey6dfyCA8ghTIeiKzZC0FVLLp
3FZ36j69NtSrqrR75f6id4CXBNHz0sEnyBmK/XdQIIFabqzFypo1Y/aO+533yvpV
brW0AuLDUjIUvY5LAbmVaABZy1HqXxFxQLQkyt3rSwozk3YB4dAzXWhWJLDqO8pJ
aYO5rQsb2DigSf+apDztgwGD7S13DGXL5MP2HmCKAw7g1T5eZSm7gszVYvrAOVgm
M1Z3GBdCDR3V5mX6u1OP7Rg9bvotpmFQjrOXNhfCmZY/MjigOS3ZQEjea5WslY20
P9i1MYRGWdJcEl8rwkbuBPYSi3DZqwGHWU/72PMyE6AiCjzqC+bJW0kWyRfty/5u
XrPXonwpm1HrwXFvOtp7WfXC9ex8vqN5mwx+iSIZXfitG+uHji6iQqekOpHfmIN/
bo0o9zHmjRp7gQWvHEk6NSc+gDun2i58IN/IOGMjJ9ykzQhU0bPtWchUOAYbmXz8
CK8yJgtoFVe28llrpqH+SrUUS22UsvWRPyQyqrsnzD7fWRmQOaVnF/8Mt3AttQlK
fIvNPRQkrTqUfOYA50f8xvYm9uCZrWQXgx87pSBaw5Jb4Dtx+GyotLGb3NVzNOaR
w0xv95kfBi9tQP/1wDINW9VGUg4wEVFWHLkWBzkR1eauRRGlr5qX6Jm2pJEr3Y2c
hYw4ftn85hhX12IJxKVLlIrDOlsBDncMU5HauvE3fJ3WCzRV98cnRY1HfG77+Rcs
mDqWLmzJ09G+GcfcvkfGN3/oQ4JfyGqAlPP2CvxnloBEQvQZNkxcsbIWJJFo0mnH
KRwy9ri+BRNtS1d8u1SQLyil4l+7m6nBiWkArgiwOlxsvr1iG8Nr2zkwxPp5VmfS
iF4sdZ8FjvRvhbqWz3hZof7DP4DWfzglHrNqqixgO8xnHF37Dt8mwTtYzOST9wUT
uNeV+L4TlqmoHcTTPUCbwuQPWz4SsznSiAmCJa9411NUmu5v8WfqP4DBwzZUDhRt
F1IEmJewrZBxHBKXImB7k9p85aULg87pTSMbQfyOqH5gxjNSmenMl+7mOqcO5bEc
WaEDzlprlkPAE2Bbdyy8CWuFn3vQDfKlYrBru01qUe2gv3daOFMpCptu0K7jmrdW
NM2foZKbwjOCQUOqenFPYXONbSwhSKKOJz5k2osClf3QjhtFcP4kh8y1RNYiYbiA
89iNhRBn0nDjnpk/7QIhNpnV4LTvjG+/oZkpis/4ukVxOaUvb1XorZ7TWj+8ydsg
IiACmFRN+exkVkx8PKKYYy4K0o5psfyvY/9Bu+dF+PLy6qbX3af6msTfZuJ11jAh
yAodI80ztiDt//AmsbVW7aeIDUY4qs9bdDJiKqxavCYseUc3VIJmHxwLBFl5wAkD
WP1Cm17RkiaLVUuKoPRqw2vvo6sbGBfW20CxXadqRqLpZyQC+NyUCSM7UPdEswqD
qgC62kw55LGHY5Nf9HCWAqL0bFwIdcQmL5YVkFnd4QyLy4DehOCZD1+Uik4rA3Wv
Lkld0Ki63B6ao4r00VTlxqhh9rmuyVfvHVd/UhERZA2FIaj2r9Z/K4AKEq+8l0oX
fQNLAyoCUkYUw1A9IHNXhbUcy0YAxerK/xG/aa9RXQbd57OSSXIuOhEE5pG0eLb2
p2QGn+Ooe2K10df1DgHWYOmT66vqYi85+fbYk89J3gvag58rDmRAcQkvKWk6Y11Z
c0ub4+hWz310AAb9AtKBKaMbPldOjPx/25KG21N/maKwUMaAGx4B05/5aUD7RoLY
nMxzLrkeJDPzTbMwK7rKZP68Kq8cuwwqBu+6v6FLB8xzTtPCLgP3paep56uqrbwH
7MvNeBkyXLKdtfRI//bNsRIGi3m515LKT4X1Fn4intTWtfDNooVIiYJvUqlWqVEw
U/PtCJF5KUQXGMzvvVuqWPRI/Xz8XaDNatOTFVuL6iHUd4g+E64Q/AxrxSmz9MC6
cwdlfZNpED2+TC+LxuugyfPUP5adeDyZdqSmSqOZcP8+jkxxBSXQpnrgGIHcJsnl
nrGMvSkTY0V1hdFj4nWGtqZphNatqh0ch8DWwbum6yKmxb7OLLoxzOI/9aOyjEe8
DCVHqgcILP42y1cSh327QQn6PhUTrL6MnUwB5sI9rxisn0B64oOhuMhem9OC1jZr
wcL8riLm8Wrcv+dvOvMERr+qxFsYdI+skkeOnaYMRAjpJR1gFj6C57KdxWW3QkzA
24AX+eFVHOcTZY6TY7AwQ1ob+UrC/3b19Z22l/7oViCWunlmtU+jYPnN2hhdtAkL
BXP1zBb6ZeQuEyB27AbBEjhvU7Vt+QSESgQXn7kQphinMkiHKxB5YUmydfGlzeXf
w2MnNMu/LjCl7TFIkUGKtnlGyJTLsMmimPZVa0jHUabPIPF6eAXa4xJGWcqWlSDI
XybUe5jx1130hhbwmTSBG+xo1Xh05I2V/LDUf+ktK2XfORXPORg47i62cWoItqeb
48qAH5bMrAF/3EX0V9zGKum1t5tmZatUp3sxebBORJOqgGA9gtZErkn+bKxQUIqP
g/CapJWGXbJSV7pnx0PJ1tFpccE1X8kLHP0s13Q95qYNVWLLiU6e4Qy6kRHON+xF
IHcK6ubjrkpBFTgbrHEVmcRsULCYYn0XQLA/ctV4P1SS4dl2RSDdIRUEt6QrfIn8
mbUPqBF0J+/gZChIz6036vHSs/rZHQPVFt0qO5pkCb4K9VTPOeyZYM4jHyfaVt62
+oV5TaSME5LDZ1Bv8HdhE3teBl1Lu85nYhypsALO9hk2IP9v0bu3aLbQ2cheJYb7
+A3z4PdT2y6vzsAUlzIqae7AXUVzEYR18NMpUVzHs9UFmqIKZ8bctk3dv/FAd0qR
R0Mn5uz1uqupwgHZwwzjP5NUV3Y6AvllPTC1Szu+/pB3lZdlIw7ZykdnfCVF5unX
wN3ElINJq59KzIHE0+C8wlq+NiD+WJO3URtzKSD/2NaT9XRdPR3uBXlyxCEewgFF
pKffLQ23xOq2bD95lShhiaF+wzyg/M3bzgnvi+ccUidAKXEjcrRSUswVASwUjgUE
4M7wdTPBm/7gXJtrPbsC8WHz/aOuc0vW0C5FEJJGezratJRvpXTnyhSL7JAuyinx
ulieRQBA+8ANmirSOMImq59IIdR0+Q4+2fq/c914Gy4RGpWRLHjtJfNabQA+kpBE
pDmte0cv+CF9FHDUgqqccLHfn4dxSOGMZmHNxSgOJQ7sHuCmSxHx60OTFTDfp7cB
tDiHEXl0AaNuzwJAXl0KWwqcF9ok3f5fIYBI+a+984SDwBYIviUqoWv2OmzfDCy8
kpqKTBx1bLAPOOew5OkfFy39An1MkAJASUtkcT11zOoyPGKlfKM7yVyW4T/JM/p9
lGktJbeVW6o1m9rfrfRDHgYQD2jm/gGRUySBmENd0LXqhMw698i7IqpGdT4xqtFq
700Xjeha+GZ6ig78gZiAuHhqnlVUrqtVCmwqNM7ZLiwMYhI3fS2e4tb3TVcRwsLH
okwiDQu5I5Z4FJOxAmfV0OH1ql4d9gg9gw7ShX5Sujax10vGZ7d4ixazVRrG3d3G
6O8cP9wqM9uRPp36iju9HD1CRbsvKC77ujoJhMNcd0CmIZMQ7w18flf/JTZoT3/c
jX3iM4hFA6SFBg0sDwJ5+ZaQYzDRwxVcJCu7tIBUs4V0f5zthj6eWhd30eFzFHXx
BE/rBop//E2OrEYmtHtQnaQ5C4CehpbDBpzCK9dlSyhVtvP3loQOD7ebfHgDzr2r
Xh7PWiB1kPoAnhxxb2mJCSUiI4nzUwH6eCzlSVnFe+1Dj8gE8rI4Em5IbqzAe0bi
nuS4d2xLbU1wtFwaoUXEiQq1NwsvWRGj/6McOKb0AJNOsNMTPSZay6OalVbdaSfO
+u4f7yQkw7eqAeI2zmhgXViK/8XiirhXfR04KrnbaWfTD1zgZC5MZQfbFpgh5htQ
9/seYyTggHUpn5mKWzky+a2U6FPu3QBiw41lQltncQaRMnvfqeMxp0rmTvxf/bIn
m7fGTUx4tTHkcjAgdio/88HkBDIniEJ995xJOhW+Bh1qHP4vmsLbdMrTNCBffnEg
NGfkuq/amW7PKQBPhV+iDupy5JKv2ohyeH1HXD+S13/c/4AGLrkw4h0dSEVLAWFa
d/96XQIPUEk5Ikh76JyqCbWfQSqQAU0yMAkcAxfusPkVrtnGerKg+ws5xHLB5190
nYuw1DSt9OhjxPxq1UpV4K1zEJvQM9/+jBn3cfHV3glXIBMZmtVH/CQjlGpu2PNP
TK6NyGidoT1MOuLfLccpFIStqVXVNqPKIMZ0SzWp8zrCqkRVV+uNmO8pxRn/fSMw
n8clVWb0w1gPI7pJ0O5SP6MSiTveEMGDQWJ0qg6Y9OjHHr97YOBTlwlUnbEooCCx
pIg2dvdwgjmoRn49WhHx0EFpwfQ5P5didW8Vszo7htya+PedkSMP9+t1Kxjikh/v
9I4hxtHUJz0HugyVtEMavSMBBZ/2PZLzzIoBTV/hbdkrN0HstkU1CGIJY3FfxEIb
EIQzrn2qoRlX50dK5JISFCMQzOzVbT9EUEQPtv1LRQAn2Awx9XaqJxols1Njnwoo
v8ZKXHY0R3IE5OHlVCmR5vSYZvcE99FBy8DNizKklpANcZzyRaxZp7gxHrrxe4a0
cDDyWuHxNmtNIxQcpl2M4Adfma2GA+qLYuz9TPJnvz28JXDcz/HIAh/MkfMiINsf
UmaS2BSKT6W6MKZxK8DdBGd1fr3Qw5GKHQrvIqsXiVpQGHeq9GDtqx0DU3ZzS0ta
zMCJ4UYr0pgULJ6kCy29FCqIN2FjT7Mg1KE2AaodZfsjOwSroENeizawseoX5Ew2
hQlH3Mlb16tTeFhF14p3XIoMIMhD2lIg9R80JKPsU1lPhtHZBrF2mp+fMK3J1uwY
ZL8TUUimMiiYcBHZi8nidKxsaxP7wv0MPjdad1tyXAJfy5ZxCiXW55rC/J/iJSoX
s8+xjrM/3gyjQCDkSfNdZc3q0hA3uWn2//u2XOwCC5OhkHqbEuuLZmmr6DhX33Rw
hLftwT4C7v6+C+V8EpJ0BpcMwQ9mxoCB7vOAKbSDEv7mHWT6MSUoKztUrIMuvBf0
PGVfOW6d+H7YkfQ5y/zwiASjRoV+vptsbCrg5CTWskVapfnp4K67OGN0+VTs3Kye
bZL/XXrz2FtZslyjV6Qpr9rWiPSS1/jIwY842OmwisaV3XyrskpJPY2VH1+zd4A9
p2YMAXkIOO57idvemLl3vEq7r8DFy/V1nLnEawmQlL6VkV5pfOH8/ZQ3q90guiUM
Hxy6gPdft7kvfoKAcaET58OXt5mY6h7ffLE1te63sA2NmdUmH3gK9Bg596Mcdefe
p1AsDFBkbivZa+qTBQUXT+zbDw+uKKMJIQ3tgQtW0QrBkRPsGlTCLvYz0rKbmKEd
UyUfPBUBz9Yk0163c35L73Z8aVnMz3b7j6yaYDVcPurs25ZEDhj67v/513zeFsqM
Qm2Klo0t7pKJ8lVnOouJYCfcuMe5cbRku2P0In0ntVr+fSzkxtuZ8kRIuBwknxqG
iCB2oWb3gHijf2/KfA5gCbE0GBZdxCQDTxPdyvKh+zXgN/qR6Y9QXWbo2IKSPArA
mdZbjReDhRdVymfyfOHm1dwupeTeOIkqg+tkglZ19ffUU+82aktWJLr0spIt0fDc
kBM7LNT1uLbgDYiBU257QGUDHf77CTCWciicnwHt5uiczM3jfTBDXwq/7Z+eWUd0
r3u85UA6EKeVaYuFSj3bj6lbUm4Li8u08ilCewQ2RbZ/6eevfVnRDEzuvkcCHgYd
jjx9Y695oJ7UjGLBEEnirdhJuxmUJunQrvXDvoBXWBkDFlkE+EZnbsoAfJeVuExG
P6h1/f20pToi/YllYNwL7nx37LXPYP0avi5CVcaiopROdGMJvCR6Xc7LBneQj0QV
VNEuEfmcS5ujVYIbjs3itvoDpAE1iEqZScOXid7fD4IOOCwnWB3hGqCPr/jznyzH
9/x8K6k2X924bCtDOnmBzVdzPHu9a4BpYAcQ24krkhvfnVWwoyotbUEOKkRhIAPk
5GMGVM3LN9Tr3DhwYd+3QZOrcKsW3f5b6WteJ7dR9XdpUHQGV1S659f62Lq8tWWq
xvp8zeKkA7UFGajq9N1Tb1j7WF941hXIl7XIFxp1Xr3UwivbfprCnTDwYkp8bPUh
DiLhX5E9PRCK9du/zNrkobfyid7/Q+aTyULoFXkOfWZ2xUXiwOiYwSINjd3Qzo3a
ztPnaNOsGZOC4XGy4VT7vfIe+3sQr2jDBtegIn/4g/gwgBAwTPTGMhhsLywPVrJE
rE8+YSdOi4QJFJRM0YqiH6Vwuhajxu4Z5b8Kvrfe0iOOmcW6AVy9LJWkmF8cpGkE
vrTuF2BUqWF7bQUzYrvjAuMJ3Vk3/w3YKvvJXRHuCKiVz+5NWrePbzcuc3g6+AVI
ZfHEtA5weCdxew/GuOCCKYJwKrtXB8sc15bDursTX+zDmDozxJvqtiahZnshcjj4
csVBLDBkjpwp4x1J/q3D7ncvXFbN12iTQ8OffVXicbaDpW+MVojxY+XY++yyi970
h7ZAjk5dKH3KEbvuNYLl9aH2ankEJjwLBmBz1UFJYQvGAYNMbr4pm6ASk1fK4vUv
dtJ7izJdGEfmmcvjrmbaLQL8Vut00cU+7nYsGixDii6oPoPrBllkjlb6ZJVgdlEb
1SgkY7nF+XhS3L02/lW55mQ0nCmOXKb+DQJuePynrcX8Yd/1/DyKF6FDFZEdBzST
L33qO2+7y6AQZrxwlQdTxgNwIOodRbR4WX5Hphz47yzzS6bcPkecVp2LILUGRMDe
KxSALwvUHbUNaIoEksaU1TkBIppQmEEcgA9k6EN7rRoQvfvEnwextH6AurfIYt+j
F9TG2laMv6nEG+HxhP7iJEg3bv4Se3UWOzEqOQYw34le86r6Gj5Rqd/x77r92Lc/
YvYNaTpjkj8WnX6obPTJKyh1QEsArkjNsQApaFQ2hVrRd2zx2k5xJvYHX3MLqkbX
QuQO4tEBYo4IjhKDVSF3ZtUspIMX8OamB8TSkF1A0InbZEfIhMtWRx+ft66GqjwR
yXJVOOcDjORro+UvlhZLwfSeEC/NCyQU+XiAhoB3XbaZyimfFXIu54zX/Ey9X+jz
TWJmDeNnYdekkKR6BURML75QTZeyM/vYzhtUDSbbKng0cS+GWl8xjaZdZV1esZ8S
Jx7Gg7adojJ0d54Xd40yAt45TV2E2YhHTW5iZOawW3mHxyHfRoB7ninbtR3RbXQu
zRrytGls1Whq1TKJaLULMbTwql6M7oRv1/mOIGqtkSHhtbcRIq6lSRAhjbGDBlmK
7vOJT6kVZSkgkIDk6ssa+CWujbSHOTn0FDbp05pMm3hH8OxHLaklWrYbRvWrw1cS
A8PmV0xSCqQw2yoveip20yn3IzO4iFc7CkLmyztCoPO7pRdPoiClJ3L93BRjiUnN
R8unC7O5Q4kmKvg1wRaR1NMeqYgbDAncOoBzbC302B+rXNZxwtfS14IaMKKThQuM
I5y3Ykl+NBjk1YjTATMQ+GQsnqCz70I6aYxT6IqWVZ3QOikAtOT8JiRUTz+r3S+2
UONycVeJieGOZaZQ+IvFBKXYqkshpCKp/4ITOU9V09iFvWcKwbzhE8UuBMBbtrDL
jjvLTyPok/qikMkOvIVjzOa5khWOXuj7Ul8P9W6n8Pf/cwDQ/CGtGK0W8FYZKdim
6ne7wNMHWdxW7KK1GJM7CO+M63KuVxrUV28649ND1Snx0NDOVN+gy7Slp68fknEW
ijcrGEm3aMXV7LMFfrmzNwsqQ0Yf3fXDv6Q1FdYYLiEKSXDP462kx4dnajy20zvQ
AMLPVy/MDw/oezoFYtIlnFD+JaK7lIX1zLJv1uq+C25PoHco1roTzMqajgMlPwbD
rhXtzEbHSc4QT3duQVUlltMFucgTHjDj29gOmEVSawlGfKYktNu6q+sRwqeCAjo4
+Kr3mIYMc4U099Yu4fgAqQudchf3NIlF0HeSkaaW1b0dFO94I0ZDF/AQ1VKoEiQ6
I/0KacCCAUaKFXigmsrBokn8Cyy3RECib/CRKHS9zkWLMmz1rp7ugURSF2ZMx+Ub
Id6qbKrr6AcPncmOhF4cniaSL+s0s3CpLBTjIF0sghfn9o3KfjMKYq7v1zbbY9+y
swBtWrE5EtSeaJCUeGDAZ22hcukTDql9F/gV+DeiJ1tMxMQu5lb7q9hdfpFAEC4L
FxNclAwr0jgfC0qP2WdPnIkKyoqXAq+kENo+YHO+ws+3yI5XWWtBP7VfkKVN/Y/W
l198w+DTvscRLpJFa9hXKwPe4syCvimfR+3OEygva60lXwLc1AXQWNwxMZUhoPhs
e+VgMhaNkI0Q4v7uvxgFEkhSjfCDs6QAe2zkO88kUuNSWIwFHHZ9nS1jQb0Z4Iji
vcQnueXd6kX+4Ix5J8xix5A8qT2houEOIoLYPQgByMuJZBz6AISr4cU0eO5pZVxV
lH6wM+I81QZAYmyDdZbPwepUzZ8hkNc3z2SWc0l7XF0xnpyc5aA5IQCiIx0CStbf
tV4bgZLT2Ep3YkniZB4ib5AJd0ODpkHvtySXPQo/+mKlrh7dUpkVaxzV4MXixEqx
vVDBuxSC0wnjACcpSwJzClTHNu/EQRFpFUcTon9M3nIWSCrCPGfG4eoBm3o3N3Zy
LU5e/XLJ8ZdmFPnXuwTEedCUavBD9udN6jmO+a/sxTTpv55P3H0yvwNMq4LAWGnm
tuzWYaRzH10mTcLKbRvLPGIJOWT1fLEL/ewztCZjVg1b9IYSJTqPs3r0SYYF10ZS
WG9EmlDX6ayZUa2DRqJl4uCp2kUh/oWdEYPsTaUApCLt/c0ap/s5Q4rD+FrY7sE0
It2yErhxv6/8QTkfAiaza2LLDCOJSnieiXGyGbiwrEWPxFHLIy+4WzX0cPIjwkCU
Y7AKzDB/U0hfiq6LKbvuocZVc23qaU+US57NTmU7U95sAFsClOGj2G5tNlVxKpU3
w7vUUAXba2cra+yK4lDGRcc6NvcjjCqTysei3nE9iqKKZ98MmJiL+jqIin2jam2A
/lWTlEBeBR8VvSfPeFYDjfECfK0kkwO6ySZeOcBPAWAHaQTudXnYjCF3RDQgXQbS
9xu8rLBNU9UZLvZ4Y2E3BmIGFbpZ2sSRxY9Ep6/K56fuqBxkRn3Y/GmZFBMLUX5g
oDHVRS0mCgwDrMv0tTGP1ljTKId89+knWR+SaMx3MGe+cEDBq28Vy2+fCiomQfN6
JobRO+y/RWSeCduuUzz13mC2WphSHkfA/7DCs6DgeXSXsmF/PtnNd1tNP6hmpq1L
LRar2blmkruT119MKTEpHcYijJo5dA0mFioNN51Wn8vhguVdIIMt4X9/2yBXo2js
/WANIe3zvCd+Hg5/lumoU6lJpvkl3bJ3VkXJGRPzjgwp8M9bMI0b6viGXL2YWdiD
vKOHGMCYEuuOQEsLr2pm6Kw3srtXS4wyfHfFpHnMGFLZM+uwp7eIhuImPkviKS+X
gzYkURKh8n0Uh9cTI1XiA9uKdvlzJCN166G1FldSsCBQcdLC6fwPxDeEEiqD4gBG
dHVtY+WRZD/jIEPydQWR7RdDj6l86y0rT07n/aUcQhmW/5V1IXjKFnGCt/gn/XIy
uINdNP2idIu0nbbaq1Fhh1EoauLD6Fl77iLD4gIaXDfHsNWxf7iAyJS5SvHzS+Dx
QXQpdmztlI5HXcy+wScIFj/hns9wydZ1pPzbvT1isjR7bHadsC9fjpjFXy/Ij3w7
4BnpdwELIBKX2agF68uCCVx1nPkjhhfy0dV1wkjYRlvJm3awk+qACFYVhA2zjwIH
4qWXMnwlyR7Aa5xVBaJWsKtOzkH81EYmITzomsrNSZSiPYdHhjIqohgKIaXuqrF3
gNjv/OYjKfO95Ej8ooGq9VmUqWEd9S42nc3WPIvVYxCdu49Vb4+hKf129f7333SQ
FqFRTy+pxCFMJCkMxLRfSAUuGbRcVamFMQbwoNvmy6TmHo5KDCD+hiEVkjt4d6IC
NhUIfftf6AYBXZ+fd9bSo4LE25EC8LCpXfbnfHWyhQt3Oo4mzl+6JwbxV+ZRlMwf
KMBwTKU4dAvHkUqqGphoc2WYjBJhUC+zNpAPEjSQIz/uUmWxMtot8hXHjkgOgH5U
YSrHR0Z3F7xGA+4kSXJPigS0Aul9KGePB6be6WDtulT1I+v46pvXYdM8YeHzzdYX
dk1Gy66eOrwyG40mxy/EiKBTYDuJ9kg3jtWJSDrwNMO3cq4gcOOFe/rIZIy7hxWz
IbYE6RsTfRv5x6jWjCQkcduciyjdVL8J5msCmkkh4vFPH6xVwYsJsAQ+NBhfJV1W
0WRO9yc+cEnyx7L81LtnG/YBHwMlc0PIf1SFS1gLR1P61MCNCoXp6h1DYojdx8ac
dmJYJPzfMnulIRfoJhdUNwPfmNEZUpwaCNbJin4Emw4/5ZUA4nN0tHdlggikFdBS
PboIFWRp4OqwOjcpZfIMfOQQtu7aqGUgq4r9mim7xNFKUW/syI+UKvfbLYWgDSJc
o3Pu1ScG3yBGHe4R64t3ijI9x0nJQEZ749hTwl2PT16apNxbDcHjli2d17E8UrTq
m6iWHGmpWkAaXabsZ5OBvcV1lTzuPqEesJnMgw4tLu7K8T5GVc5D96ocV7/vsNqn
USHLOFqqBUJhfV5eOi3hq2ZcZ05WtNZa0Ps8ENcw2dr7s/du5cCnTi7rDf7+0e7A
8HENoVW5haV9FQJpwHOxZfh6aksWgceoWG7GJ86GwnlGf5oP9vnyI+k0vtp3IY8t
si5PwiBp6ECt81fxBbJnanlTMNUit2wGF/O7/izG0cFHpcmAOvxHi6p9zLwCnXEs
QTLZ/B1wmb/gJIxLMHoDgyyqLGPSqEmp8yT0QzaLoaTI6x7bHlFbOy02H22WQCU/
eduDv67MP+assdiVxHOYZIZ2dKGKjEZmh5jhNEp1NVl9mRUqW19PYhaeJgcvciit
bfAWo6G5NhK+cb3DRQQ6dHJp3XQ02N6XUpJ0HRrqyZPJMi2MnWN6SHj6h/UnluIn
4woicFx3eTdsjLgvyapPWi+s3nj1/fR5D4mZpDol07vUzxyRk1U20DEW/R16TJdq
uuQEkCm4/gdSZclJ1VMx1dIqISXAWrIq8BN20vKO/7RYu5Oba4DoZvYRSHivMg29
jyRoWjS+nUemNbS/Mu1047eKGKAaPNvM41NFxdm0qldkZXmYaPpIdvK6pT/CqiQV
1yz1hliDNxmNSid0wBAL+ZE20lgyovvB81819QVlGf09FmtzJN6H/L/s1z/Hu2nu
8471GxGJ0wpVq00ryBxpQKFoe2VInIa5qRcoHiJparl0hwV5Gzaq74ugBfAjwuxh
Fo8urnBrl9+bFlO82qcvLanZ8LtLaf0IZ/EEScPANngp2zmSzil0Jnln5E2D/T7C
ubtIFfvR/i6j6lHRwU1zqrVmuMDhUZqcg1vgakM+1uUxJ8hcwzI8LPX6mD48wA8n
0kFiTyM63cr11Zl/2p9PI+83inV6w/18svSr7Du23ZUXDuXFGKMhHFw1e84AgzFv
0Ygu5p1n8ElF2mvQVmLbjnTdpNoXt2K+9svqICT6b+95FRQ2zorqFCM4N9AekCtx
RGfLCK40nO/EKpyAvei9iI9/+GWwpsPVpqE+ek4RbM6FezyG4v2frgIusRHV6ege
/IwhVq/Qpsoazw6Ksmt52T4o+ovQs+bJnfP5vDmTayVyau/n2uMUVJc7vlnePv2c
zc1cYxkXFWfDtS7OHvVldJe/GsbujhC/AIQi3SktBwXdQI8W9yBC/PPFCiE8Ah2/
Gs+3cM0NhCv5e+gCmdq39kKhr3u7LPpA+Xvw3HGN72hRf/wzI2tZSgNFz+ab/N5C
S5Snnihgm3gqpnPzEbqPpYsACOXRZ954ZIiY8rLCR4Dc3poJCKK7ehkEWw7D15S2
euyv7PNFBebyY0/QDMILgiShtfPnFPuRTWqf2jeGMe2HezlNcBYWfd6ughVEIYWn
lrnKgPzHNM4zf2tqu34E728DfhYVBcXRx1v7aYc+uMqRBtvK3FUdrc4lQLtq/Kzw
z/0rDd3iLtd/4FLtD42SHAg24WluObpLDWSTVsjbz7DrJ0dHSEeETAEG3iA0wj8A
UjIZPeo/VxLmmP6VXEuZLarjvahC+MU6VJLBkHuEhv0zct1EtZL3HdnbO2AYKree
jDdZ1xmq1mX9a5GK/XmK3Wv6OZQmz+pODgrQnOIdVUi0vjQzXrIW5WS7u5IallYa
KQAmAMBPbr93GyrJVXtzsmoLD3ArjAPLGqgRY0jQh1VVgnOghFwVaAq1XRl5FN5H
vzMSJ0MaJxKXaB88cc28xz+MQRsCXqZH5KLYWshlRRQ/txybwjR+2qklYfSFyDJh
mQGP7PQf4woPDCFocBmGL6E4hAMZPV4LFuH23/C5Lt3xKWbTBW2OZVMN5yfB/Ivo
i6KLQYP3vW++yzgazy5L1nK0WuUNwC70mb2LejQrPLsoJSRw6FwRRM5jSR9t70Ns
F16XtnDg9hnzQm3ubMDI+pFvev8rcV+TsoZjgn1vmXWknM/x9rbKnhf+79EyOHDn
g5XXsBTlAi3UpqFMNl7RtsWF8jpweok0WZy7P6LMc+EGgr/qJr001hlzTcKIZSmh
VlK7J0OhE05zcMkevkWbndrJJFSRFdA4/EsVjpyFbbVZ/A4bwe5JvyNp7H4Uy2Ks
0flx24HMJhryFIfmsm750T6vtxAeNWHTpWK1jsJWMLgXHbaBKrGnMKG1YN+ltfWX
zOKBMWOgEVIMElpCLCwlprodTgL2U0f2i98yR9OcndnJVsQy+1UMCZ9nxD/uCuaK
FQdO3vfWw8GzAG177aMBfR3LlvD6LaZ9lpofPwtIEirk7YpjC2RANqky4rsbXKnp
Fxhvk9UsbrjT1GIcM/0jWvDEkmPUcPJpSLMAwjikXTLyZZCVzvpflfIuVSgbg9Mu
olr3ektUDzKhS+PrqbUJIv86tM2bE9Kg6+/3yQBUdQIEpUgMm/LQ5dnvXClk7Eoo
2J6QsUuXBaPUyH4jLrN+rv+r8gM9vWWqaExciZo4Gz3Wzy5T+puYsY3BlD1JhfPy
RiQNAvzwLkPsog7YdvWtXL8WcMJYH/fdJx4csnTJgx4U5qkWJmw1z9HL9DRiHjxR
jL2T0n7eJ3EMuAyQS5NhAcwyTbUDucd50x+ynq2yekrQ6uOnsZjgzZi9Sx8PeRbN
669w8v5Ub7h6oxQD4vAElz3tuLZmE1XRoCMf3BP5Q73qeFZt/TNDRLHbs2WpxtV8
R+UGsmAJrDZTxuzp7WhYvKmKKx1jPPpqEOjoe4RiO+vCebBBGwwQsouvJLIY6CPO
UnqM/q53AAdExTg/r/1z+q9T3ZZT9wRXceeFv0OcXIiW6u679sRt3HNBMMhZjONf
EyPjOu85q8zBZJTx55OuXw==
//pragma protect end_data_block
//pragma protect digest_block
h0pqJSdxIV/JlGxvxInpyoMSN4M=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
c3yz1IpQDtIUw26kKMjMUTJdcDE3b9BlPip2ameeXDruCYPmAAh2RR3NKHTENZh3
49RHv6OZIQgL6c0F5qzZT0mHdo29s4XmVEIVrazXzPco1ziWeWpX9/XBC+fDds7B
PNJN59Hj/d59aGW1Z12Vdog7ncH4IwnlURCGq1PhvXfvFFzaSbGcyQ==
//pragma protect end_key_block
//pragma protect digest_block
PMdEAGU3nA2wEXHQDEUVq6HZ8ls=
//pragma protect end_digest_block
//pragma protect data_block
ivixLo8x7t1z35Pz7XiUA2ldSk2CSlU1+RwkAO17B4PgSjtyB5jx6RbHBssQ1rbO
mLwM//P5YuA+KF5yqD8ZRu61VnuoprevZOpRJbiYxcMWMc21i6V7XY+cNZqv8H62
m4z/zL9Uh+BeBZen6nwwl6zrBdIgXClCZ09TuSmAIm/jkntp7MB8rF9mg8ZEPnS7
KfwS2IPGyMWDizWbAOWqIYHPO19OGHq9WTVttLCj4jJ1Megv/uUKIJJCoQ+j1O/W
A9at11KwAMIz+O1jdaA+DQFH5QdSJPX1+OqgdyCJPM1It8SXENyz4B8Zm0XrfP2Q
rnABie43iN72EBaFYrSoKLqiqmltu/JVr4kZfnK9oHe213ExLIC4U1ptLDKNLnVN
gNfz+meHj6SKECXOB1N6blp6ZnMqZkGJ3AwmpzIMB+em0mEFAq6LPF86LdJ6XwCK
b2HPlsesyIfWct0JTJ7Cgg2HGtfayrYLBKUWh/yLhnSD1NdAZTYkYqAjHJ6iiCUW
JzVEFQe+pnHRQzxv7Accx4GuPslNaGKlUiq8S8LM4K0=
//pragma protect end_data_block
//pragma protect digest_block
ZxeE8zsbTEeApnloSJWjhsI/x8s=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+lHWJMmUywxO5ZOV4p95jjIthDOkdBGrto6z7tBh8fhFvNmXEWx+sZvjseNN/LBx
j7JWy5/x9e9xBohegcJ7zmqPV2srxR9lYDS0C9AzZTOOqJ8ORxe36TNSjNzU5LuY
DE1L3K8xNqkLPKl8YcMvwJRhltVYnpdJcCars5KRjWo4W11KRx8odA==
//pragma protect end_key_block
//pragma protect digest_block
lS+4HQQxL1TmY8E1s8nZuSiF6/c=
//pragma protect end_digest_block
//pragma protect data_block
S8EmO4kMJOUfO6VRobtRNKuYmTcQCAchQ4VprJQPZxo1OMvqArq+F+XHmUXOMRKn
xoCr5lFwyfJYN9gO5BuDXXrAlgbxtkDl70WEJceyWRA5c54uyK9VJhaabrnjOBPD
ouSf7eyIOnQYIqu20sHeDlVQS47tBuaaSwP/0a4nblQc/x4f9yCdN5uL1cLembOa
bjZ+k31Atr9U69E6FnUbZBg1/3vCMmp9pXLGiLwaF257OLFcPzzepf9mYRPtno+u
NHdvKiqLniIncsGs8bA8ESJBeX/wqoBSp1eHeA+auhxdE0LOR4u0e9tGXqH1gAw7
XiiyvIa6Ahbbmc2EsQufbHP98gRlDItIevkpFsEOJvWElIg8VA3hd8X6hNvmL3T9
lVy3NluqE6bXMJ48Q1NNweB/FMibs9Nfn6Fx77pTIKE/tTPnBaHiBnNPXZHiNzKY
J3aTXhuw9+SznfPitY5o896yEsRL+WEA8Mbc457nwGJibvyLp56+/Ol/podkucnp
e5ohOm3zIZ+GbY88NLbPeT51jMbhnfWwpcc7OykBy7kN+XCRu8uJGDBDmLVPXjMI
57pwjqGU6AP9Ic3jcInfZXSz/omSyLQewcBvCZHGixTA56lXe03A680chAFn4FeC
XV8u1t+/Q6Bl9tRS1hZVWiknTaxsMOdFwXA3jRl3u6OUAn5t0npYmM6TXQDgPW/0
Tin6Z4m1revmUI0joCMDhKBHaZVgq86aZwSddc01poRM+Q/q5PXAT9Z6M7sLaujM
W3yypoREiz3KsfKlM9TcPR74J5Sa22KzTlzTSLTag0tlZv5POoEyTmJQKW+iGhhA
pcEtHQZPXE8T4bSJgflah5yko0PIVTkHNKIagldMIg/XGCFc2RusgUgZ9DyIDWk4
b/hbEHsKz4uXv7n5jqqU59jqZNzmmF/toxX4dOyO6kTHv1L8hylmz9XZ8YBpDQkh
6Yp0XwoxFFv1P+XQkV3g+FH6wjrYQsAVEpMDeNyMaXNtQEsHHXRbM6tNdKrecwCg
9J2SwWexthy8GqjrqMwUob4YvMi77YgsTD0XCC+t03N20HBJypfNxHegyCcBOT++
7gRnNf9nkywiy8m1HE6+sqmbeIBpQyXfJUhDBqIn6QDaI9305iBiepJCbgnz9kS4
sAZ0hqP3JNXGMIcsUbc+wu5Q9frfO+KbcBqmFTqg64z/lTOPXm/D1Or0h3jj6RuS
Vow9vRmYs133dvccLdGRopdIBvmCZpe9sobOfLY37kuZGbeHK19OZK3ytUmbPAX3
y84Ow0BBsT6Z2BCRwF6A2aJ2v2jUTSd3hWE38iuLLmlY3an3eAfqip+gf5Spen+h
bgLk2GGlPWHITvtbNU26nh9CV6RNpcVIwDJNF9o3U9FVfytVhocabUGSgaVyq90T
j/TMi37NEmvp0Dv+O9+nzdwt7K2Z9Tku+K9drRNcn9+3aKgeZ96gwOuUguKFqj85
1eTriBIo+v7y8aVh8KNNrSxrjeM7HpN/g09zu5Aupf1vV8bwZMB70XI8zFpxcSC5
PnjavE4hddPo9nwqH6e6SHfyU1YLa7krYqBx0dP4+Z0vxEfe6ukb10N/bVn2NP7e
ROdLAErnijwem1K1v1pfs0/nKi+oi51sZuS9t4BHXw42I3dqOIVZALuZZ182vBbJ
EW0Ru1Pos7cOMa6ybKCYZYDTyBv/gsjtSvvTYS/SzN1JH66WMqzzCC9mw9TfevQn
3qhuvQKt3ys9UfzegWJJYvpeYY+3m0XpJifvIpu/BsMEDGwf55TtRNEbgeSgtpLr
9sWPo5rNrQm0ae98YNV3QPXvodg3mptip9FbKs9zGDRTv/SqND8KUwQyhBWF0f+5
1sY92i9uWe/WfAnvIblDhQMZi+ySDIBu/vxwwUqFqiqIfJyS4TVqHfzLBZMTb4YO
993NHfBD3DWbS0H4Pjle6UJKFHlP3mKam0G2v4ky9V/+UzIZ42i+4wl2CPPxw+Bj
O+CUDa2RajI0K5xxawA6817QHylCZhsUppLJ1Hx4Uo++aK5KCQMWOjfWB4GMFkD2
id1x7/aIYNMv6UejHCE894PBV08/Ml56nicQhoPjdTlHO/2l6QSntwAiGn/K+0Jl
BOKv01CBPIkq56l4JVpcLSS4UHaW8Fxlzicm6gZTvaaFxP1Zon7xrT+Ox7TZmj/7
UdUJ7bVIciVeA0rVC8LH/hmg1+gSgw174/nc9kzEP8WP0CqPhEO2OYe+f3gxAZoL
bu4qpUz1IbR/wMrhJw/TIMKUbVeG/hF8MeB8yQKgtiPyofvxmdDMM3Nx8yYNQFiu
ebkhqWj1obquzYEQlcpgTiy/8z6XTc2aMO++j1Dg4ZoMEa5E/jt+OR5OiWkwrgZm
L1ed1GAQ7TZBibrICXRaooNKDAF8Qt/k7NAVF16x2s0ICLk0lHbu4ZcudCBp356u
C82+utx9SA9dyhhn84VlJw3YCeY4fdlByDB74HkXPxvQRx9VqLb4ExyBxnh6mqs4
vjvQ8wFy4Pgij5nrjriCxPXBTq6w/1XjrDOIUs11Fe0bnDD0X+kYARdY4c/xDGw7
/WDhLcMmUvIRgIuV9CDwgLVOIReUjCgu1d3ZCd8QGmQHCn+UMuJd374XqmeRSwGV
WrUxlqBfHoAp5vdlLIzpL1raQGHarYfVcue43JlIBgs8g5attYwq6sdgANKllhJX
HyXgi23/fy5RUwBPmWgd++ps22dZ5pUcTcPZX0bBaiLcTR/3Yjbi8npKtasTVPjs
+Qew1vG6OtiKKY89cpCQ+DUMXgfluiFwx2wonHitSF6sLXAP396IPmnMeBYIOFmT
lvSgditkTtjJdmW1TzgIyX4a1Tau4sNTb1YKAZFVhIcf6dqt9Ko4FKsd2qx7mb7u
+FsjumIPIteAp+g+5JH9aWqjoLiicZ5aU2XNa2meTuYGtpcrgHGydc88WplIsJ7m
c0cJu9HX3KzAFJxV5wJcCS23DUAbi7DKZZAe06HTsSFVasecGCBrdsxIgmFK6Sa/
uk4awJTlpwzKKtgfhyrFrGu0VA7l5DAsZpqpxq9JY8ig7vluYwWHl5vOdSuA7AD1
dDG6Qr6kQjmY3pyYyjusjGqpiQSprXCuekDwzJb22w1y7rnhscnJ+RGDqfVL/4qr
XmHgXRscmfrVyJs/B+dy3Ech+8zHyKsQOZ1lBYXISy8BNziSZ7u2CNxSmdSuYO/6
q13I50jvOzMm9zw1XZxTY8A5FuKyqWsR9J61r4WMwKWZ5oiRoLguxwdmjJ1dZL1V
6tDrWMCzW1ZRubKSRYM7OmZN3u3kXgN8mpBr9XanRt0TNpN/dkE1EUxic5L1Sd8V
Rmq3RQwHjvunAXpR5ZphngJVDU4aHr0Fk2HaQdUWdwdX3fFf02IXi7pLxBtd3KQW
rNDg5ncU7sLRCliL/sO8m9MQeiC1MyjTIK31Ij9Mjqw8x1QYgLhRhlavaxJJV4yy
XK+NH/pu7eLKT8hT0m8sSqTxtR6Q8Sau+i4/cGRoRKJkq+QUCs+8JB4HJ4XomzzY
jB0ErUtY0J9OZ2LD8v783Y7T5sRzh1f2NZYyvVXyFjsQnavUcgCffK7dWoBcZA55
mlVxF5b2hy6r0xABdxsxwKtTOPtHon8864GFi/4Gd9XxOiMjSyiVlGlx+AuIqTVG
gQ5z1vLbLP/PVoRvBF0YexrvKtJIYIyhbqGmV0RxxkuPGtEmjS7BPZzV2xgXFLWj
iUsivObPh/wy4k/dPw3y0RDOLwUW3oyXHybKfuVguD717voupskId4UJmFWqqBH6
8wjaO0isVdWpEOAHkvRGcqJ9Tl1/n2McC231N6CSI7yAfTm+0dcPvbZuxXoBWOU4
8Y9suZmYoqvI0BLzD05qlft1fTpXj0gGSBmaqzpZKR3+9jOigP6EA21WUFDmxJ6S
Rdyd8zihMlCG/TjGX9x5yaUGUF0sgKeSORrhTifPYZR/FhzA9RuarhVzSoNHY37R
xDx9RBhoGOBVil+7GG3rT5+C5dLeDn0Y8i97klpaU+vkgPVcqgMyHdHGo2O7NohX
dXp1bI9coXho2zJoQHhQeExibXsfPmezziJkUcH4HHSRa5N+gXkPGxRSw5X5I5UM
tKuM6QI9j7otYD7BgTZjrbGS2u9CAs658wRcp307RM5Yjfk+c062jH4P1wPmqDLo
z7sXuFC/52wTUXusVQPKVEcgW/aezgpIjjJ4s1RA0h2pXr2bsiJahb9D/iesBHOz
YIH9/CioZBdUyYo2hREyrtfTeJYAzr9cZvm7JBOOsyylgERNLhKKBv34WS8snfg9
zrjrdaSlWxygRnfKf1bW4lVjWaUY4np9LDyif2rS2Ledjr63TP5MR7JqYczfE9rh
uDpDe0tmJC0jVm2mKNrRXyVTK6W/7LpNhDwsg6cTftJJJKzNw8EwYH2p06JrhL9v
pDY1o7IBzvE75pM+N/Ltfh1IhPizbS7D2ArxnabLWFG9hEU3sffRqp9aP7b4BhXq
/t7XeXILIwbxBCtu3x8o3lik3GGkd78ydPP6Oe3gvFP2CWS9Dkgyv2p6mn2PQQog
evwUiyjYkhY3WQLmKKeCsGYOMKTsK9bfwpHqO1vsXrOEUnwpD6IPQyLDDnbX/M67
teh2MRsJnYQ3pH/EIef6PaDSU4/AKlFmviKZ/WddB9AbFcM2/S8Zh2AEYVxgYWFD
HymZf70vO+80f+6ajOvbeRiBcGY0j6O03kCWE5qTySFeV36utW4NQqSaDecjBKty
sL0F8kGIoS7+fKSWKiSFUx7fHXT8rfdLPWsjKIXwbLYi5E02/lPaOePi0Hu6tYop
Yqp/aWDbaAwdXdd7IlK88PYdqfM2Oig4ES7I3M/T2Q8ipCPEyPzT9VAnyfgNLFmT
pwcVuSupmi6ERnO+1vY9nqR23A8CVOicATElmmTnGC2EiJBuaeIjyaF0qDmfI8F1
omr30vi5NVYNoj4d9U4LFg4YjOgpm/NrLQNDViro+tY1MdhDZWcUevh9ifFj9Lh8
qc776xj2qtS4GXyI+5t46fvoG/9lPB1JGWlITBJdpJWrDdSs9SbWUT5h9M4SW3y5
9Iw9IH0WGzp7xfOG0P0h1Q8L2HIZ0IjkC5bH5dmvllgDWHfttpee+TtE4DcVG/km
B+OzHFpgW8awkf8qckzQvYE1/U9AhOVGx4TaFV7lmE+vV0Eoegqq4wb5PwZYSV6x
tXBhV3AqqFYX/Seac50J1wFkxo7iXp8jHVCppKnHuXZ0KBjGWmOLP4FKG0Bsvxqc
KZe2h3xJQWWqcBh7uAHJ9eNlFHgTPzZn7NitqvoP9bBQAB2nU6kcIxy8KQ7cr3vc
nyLUua2CiuR8BiZydcabj+05wPU+HCz6vyc3tD40g2Rg5RiTcrIikH4lT8BCwwOA
hDiX4CYW6qlLNgf6YydcwcZfP9I5Zk050JAaX6QcwSgDt24nIO7h70y7bbhYptW9
vx3Xekt9S4ReOlY6HRFuy4FfLb7JcOt4d8buLYLZpap+UrJOhk4HDQEFLr7NT2H9
qrRjtMFg+28rM7/fvLr/BvnFPwvVRoagNuT9ot3qlBUlZaC+Bt/lPN4+3R9EeAYS
4+L385cGZNs6qwDe2z/dOi0AXe/8e595TNL0EjsAgbRI1ah2qQmXnxMrOKnQb3Tv
lUhwk/2+k+yP76s0kELW5KYRsjqeLA5TGNAbewKCHev0ry/C9ZxCciJkswMTJlOg
WTQ6LoOnn/8qItckWjykTamRouFu3BhjQyu2DKdVVWaOViqWwzU6bitQghrndzOZ
YE52F2GGlt3fY1g83JydtDCbAo/fjkQgtUBagCzpcGuR7zR3+l26gvrL/tcHpyJ8
DEdgZ2r/Z3moEqRloUNQS3WDATT36RQfU7maNeNykb2K864rImIn5Yjbf8TokQa+
iQVI9mXmKV22zi00L+gCLLA4i6kA41N+r9BC9aLxOJPaNGgQEaRMT2gyZQedUoyn
imWRw35oqxrjbObYPRbFiHCYCW3tVZyA9PJUopo3wlIID95SDEL1sHaeRegu8sv8
jjPhLElK9BgUHN8BjRw0SBYzIFOuPMIYKT1rgybvuZ7uqmqsInQ6UMo5E+cf8Hnv
S+mgdOMa1f7VZYjnEf1yTJ+VIqa9OSiAokA0Zc/hy7s80S1WhcIHxW/wPMicjA/I
GcFVr7vBhsX1dkUZFRt/h/uToyioGNvY+nzr9DBLnDyIGBvcXmzi0G9IoftFoT4/
IiMGvAdeyBRIdtMDztVzwVOc0N7IVrmicwbaLpHUKSqQQcx5xvythmJKcVpqfuFN
InC+CHCKbPH/uMq02mB6CT5B4Yp3S/gZQ2ZDo0jsfj3wGKkKyZigwNf9l5MLS6O3
8WHdEZ8v4wYmLfsi/WOTUo36ZiKAhJH190k2zMR7dyPaSuie31S7CRPmkRAeSUN9
OTt24jprk+/NNfri8b5nilpTcldibf+xPYVVLQ9CWRqlhzhaszToR+6htJ05hbMX
wyaYyxUaslyb8DKgLjH2dA0xmVorTRJi37UKoLo9+cwqA77GhNSmRCFkt9RYi6CY
cmLqlBgoFaKq8bXD3vxoS6qOu4Hqeo9BR9u+OLXY1Z1NLJeNV42z8yxcnUIgeQou
0YFUOuC+Xc6gIToH5hr8/ZwpKuYfXVs//OX+/hlUSuwG8J71rkgj/j1YqjK7vIah
QRR3FJG97smiuypNerNFNnyGQZxg0njAFOAtXVXIlmgRpJOpWoAWKdKwoC4Y12OG
ZVtRvtIz4bKF+marqacyWCzFlAZDoYh/uJ0KaVEJ/blCSPUIzp3AzoU/OZ8ACRUd
MEPtBXTV9IhkxRwcAH+WPd1TJ4saCUgFdTk36gm6tn7fTuP8zMlMTea9opV7ZLgH
puIh21bUUCiff577fNp3A27FuK7gfvjzgmEWCoFUzDzsbc2IlqHS9UzhvG87oqGO
AxG3V52I7gltlaEDD61+3Rlc7B9nmtOZevBMQTExlwnYenSDBmuboeTJnHa+y4EZ
G9JHbCZmgt0oOzg7ySOJm7P4PdrwNy34PgATiruMqoDIzIgSObQ1GZIu5ubBT6Uz
AvK9kEsgELbGIiLCUFp1BSe11ApFzac3mEAxv43aOrLrnM7nBwOPmF5P66duGopf
9B+3DkzQmFHlSzO55f8I0uBoy5ZjQCGpkYIokI1echfzkXmV+byA8AM1P5ZTD7jM
4D6+Mq7697elPpXnhP47TnUgfiD2mcOyeiCzyAw4/aZCtkMxmp7d9CJeZHzr/+Dr
sxGqYlI0tVfWq9+yQh4QvnlgCKvgzkDV9IihgkVUMVYEAJ8StkDhlGA+XgGwiXrF
anR06oka4TbHPWuWsqgbL1EfE7YsmvV9gartw3LwRwbSc+6v8ihzCnMo4ptVAVWy
t2MOC73DldoB+z/oCCURKOh3fA1XetCsYtOjKgbTkaTImzY6RhJ7yFeFGhljepHV
MGt40lkgO4sC4kfA1WuMgvyV/jWDQGG9viRKRqRX+kIiJAZBq42D7trMASuetrc+
hPkR/hiR767AfJxW2ErCDSaEnfYYnEonmRTVNkLF/ZyHdVDT94bmfGYMyc/52JJp
TWFxo+s5cHOSX54IzY6hRg+cpi1D/TJlIs3qllMFmYu2ZOcAqLGID+377jBJka+m
g/7tGIZkC4pVp+1hQ/9Afoy99BmPEhkhwvbmnLYwENOk6XqpCkuPVJXnTPDmF1Go
Or+INCWQd2av2Ft6+TkkrIDEWJSre0EkJI1GrfQUw7t6DAa4uTsqN418Q3g1ML6K
E21lsbB4bPxHWpbOodHpTq+1xiDEnQi/CHBXZhlhHBL422pdFrd7WSNc46pD+9l2
s+XxkLmNxjVcdqDVfrNRSjkVkJ87jTeeTq345XjCC4ykg1g4eX31yTG4mtvqnCOB
AMV0F2cx/TzWwzMqeIA7BSobcAwDnE3Mo/QLgOuVF31A1ebrVQ3Oibuga7uI8LY4
4LV9ENI0lQBt0X7s0bwLXrJzQdg8TmUq5P72gcHTR8wpsLMumem1EoMJowN+Z66g
/Qejt03PmTOdTfhUUEH+K8zl/KWA8Ox2BQj8szlTwOeGppP8JKngdEdvcph4uQ0f
PUbiUeHG+Hz9En21n8hDNYlmuKSDnB6LTruXwvilzioeB+Efu2PYJHkXmnNBr0Ix
jJxsLX88ESkQ6Bfmk8xoZb6VUm0kWSxUOcI3pjNFGJJ3AREF96k4WWfwrFw5Ql2n
RSTNaaVV3NWZMUs+fASha8rlQ+4jWxKHdx86WUe47IYVME9PEyaHFpLERu6Cvodd
gsaqta1PFFZC7AQECQ9831568zQ5ys6j809Yf3CFOUP0Xs2KDdZ1rhReEDzTm4TS
QCkXk42AKhGlzho489EFoGXwFfpCx6qXg2Jfk1VhYZhCuf96S5DMeRaVxf1+JFJA
JhEr4o1saaCYrqy1vMjlwKC2sjHfDKo93Ge4EJ+HUv078zSP0vU4dAFsI+3QxVjr
DNnGzOuPskUhtJS1yf9Yn95B24lHYZ0ODstkvX+Bm+IwKHbImflxuthsWfrF37uA
wUMf7HeLDTEwuewHDgEuTlK10VPIBaUYH+jg5q/J6wcepmGzsOaho1WOJqXCYAIo
rs1KUryqwEvljEKQoenbeH5fmzpDYLqyQCrIm3SqzwyIIQFR7Hhm7+TgLOhVvMHe
hNH70NmacwhGv4CDMJIU8B5LWVH9GG2wTahPKJdjWkDLqn/qJdi/643MRmdSu1fg
q1N1gECO/E/rAPwR///C2MqJVFf4hOX5mHCXA10bqKcYsiRUb7DbNo6qXPk5oczB
I/81V2UXf1OniZCYhpUdqwmtBVqCqrvwdjM3/QaFtHNhsOp5cAqufLq9GlLNdtwU
CRQr3cC5wx6oGZpYJoPZUFPrqbXx2N4o8HXzgFY2bUWRW4Z3Hi2+BD++64Tp06fO
BsUNBMj0zyIs4ew3MsCv6t9LmSF/mAeIoGNLmypAcFAKOjmBomiAMvD4jPhRaiiN
l46wJrOAW+qNjEC1bGIt0rYBp3cN3We90DLmCMQ0/q7AbTOv2HYjYIEokfILkwvV
bfaPAsp2IlSTSMCZgcqa9GmLOyy0s40izj2qkxCdSTYzLzTzN/13XImnseQh8nty
GTPkh+u6eMe6x2rNTblLa4hC5nsYHckxIzdk+EQinIJhdTNu/85IuH+DA3/DtI9k
ywEGfBcQTJUo+stJmpNLKweVMVViVO/F27XUDx9XHUcLFajkAlhKNbph3+0TpJPr
niXxwzvqbRQ2K2uOri9pBsIYdB9HKZxEckxKj8DhPG0ZECtRaTja8da7pChi7b/p
4fVSefEj21QEH0ENYh3DemC3m0FtOYvclUo0mkbgaYD2eFv6JrSjks3L8QlNt0qR
Kw4VvmS6CUy+9NDLI0uyWjyGQu7PTEqt7NLvsR6NStPj0CCVj+hM1ad2ANnmO5Uv
ukBqXCu/Ei5h2Mqb20ruP7zNuw01K/Qve5RIva56daItFXyYsDuWX7RaZoMT8fSm
VysMM5yTOaBT2IlX0066afWDX+9Q7R1FWwRgRHelF0nqfPTA93H0xKxXr8EglZHj
O5Axxf9Jm4/5Ssgd9yLzgWG38wVYpWTTHRptDupYjE+vQhuz1RTeaMnXYb15Jw4O
BHpoEGYafCirS1SZLcwhvkSWtTD2LkXraor6pswN6GGWkxFA/HOOzOSWyo+rOyXY
cDLZN1Utm+JSVjNR9kHpcZvr+nJLlvhYKkburDW5X4XujiCGOULYuv6ryKdnrJM+
CgKl6LSuJCiZ1B8x+d6DN1I6CHQtK8wNsem3SPi1xZuibbYulkjBIm9DvYNoTS1r
LxcDWPL9fgE1b52+RdvAV8IoBislHgUogAP8BeikC9UDTCZxjqjQaIV/TDGfIvrn
ArbRP78SB/dbQhjLmE3A704pGD79M4KWavM799NCuE8ZUwLTV6qSzSbjtRNcHpYh
hBb8zUJG1/DpvI1bmPD8rfvbC/EcwsJiG2n6DMf8oDIaJ2CaQrjfOReVzOSatgIm
919GUVUHQBAUbMKlAJCug5A6wHKFeBrfVw9osSOK0PhJKQ85Dfp7BUHCcVG+GFfr
QJJR92FB8ABnESbNWX1OWSKodHmaE15MuIJOqAP6X43K0AYjm1ZwReU4ievL2D9a
t4dEu5EYdej08g2JShgNbzfsAjOKohkpe3XAzFbs8ZfD2v9DGlodotkLQyJM1ZyU
spn3xeWeXjqmmgAraXYMVUcRwq627o306r3zzZUqDwO3xYb0m0wj01eBmmtvaIbo
5Oy3/7bcnuapoelj2egnu39vUaCVeh0GYnJusiXMeNKrwE3LBXQx7Rum1Y8fGxM4
CWXojzkl5oNlbAHX8wg6RqAHu4aWsPPRoKa36O5c6eTMSGRn8aN1fRsaGl4w8lEj
wHHGcSkf1ZgV5J2yFbxXDZF3Mns+mWlOL64+iJKmtQSXS+UsUxwInxSjV1o9N60F
uK+0Lo8CYC1GY8HRHMY6+pW45Bk/06mN4hR2RAtxR3PebVGm3ol6lXvO0vADjACu
rGmWM3RGTUdfDT5D5KadyRFAiWJ3rf27kBQ9jPYKuWaXntHMxm2RaANDgjWfefpL
FyvMC1OWrl39jor0Q7/039zCzzAqpytlW9QZm8N33AIL7ngcwnEn3x5W6ICzxD5v
TMq5QT5G2FUyg9Y8tqnMw1SM5fGSxOR+dh0takF3VgSOBS2DRThMKAPx1bg0floZ
nzFEJ+NjAjDaYOp+tfeqLLy0njRvwm6cmC1p3/5INURbfDpMTnCvJrLXMGB9xJAh
FHgSvR5embYbm0o3axzgJ8CDk2NHgZpd2KPJCh7oy8bzRlfog2zHWbr3qNmkBOrN
AKCDKItSa/QkxleHFVUYRYhfELzPWLYV2HHNrJ6itKGYpf/8Y9HOOnn7Vpy3MYcB
v8m6gpElvzGv2qKiduYaqEbc1gqDQF0nvivBe4mm8QP5jsNbc+zDrzX4VmRvkDcy
lmqXIIaPE3yIsimCCYadoiU3mWMbg4QXAoOVaPavhqPKrRYWHql34RfmEK7AZUuW
CItlkHQaIKuEj1tkzYHPrQIV5W5vAV1x1IXXsOCcdnswZVta9iIrWXmUD3JBwMg+
BkH+1u1sucg9NoWB3OtyKsVJtAA+A7pkOArOEYzBqcMF4golDot/jutSTT6C0yb3
nt0AeneMR2u2kGX6ix5eWSQiKm42x7MmL6G27QC/Ivcon4Q20bzNnru/1PSIJtSL
VzyUEpmOGUrqWwypgtGRsP0EEEbmBP6hLQ13pDbppOk7jIQs5rknU12pq1kQnSTM
nqLj24JWRj+uOVc9ZLwS42FqeNnSs61M9b3Al/+g2Hopdd5xd0vIHe4D64eVf2lD
XH/SIVS+ZXIB8NcpZNbruw//iBrhRc2bBxJUZ1XfJ7gyid0yW6qePdwtlWlBAjLI
k5pUrCe/InGmzGBSnGvUJ09T8YpJM7P2EpaNb6CU2gw4gcC7veMtm9+1NLD7SIRW
4iEJGjNdXn5SXoEpSc5qTSGcrjr606EadSztwdjtZWzUErJay4gCYtP9fSuxipVy
XPbLE5tOH1KykiGMppnWmWohnZmESS8fOZCGngdMaYLuF7RsZpyocnKs1HvrGiXY
3ntE+Ou7uNKq0MYE4AscdkpbXFEEsrer4sb/Tjv+BEYUawkovDgNxwDJzg1WZ9jK
Rf2kWP1xRBuPiGQa3RQl2MLxvimcd2Ps36kqM5rMWF7QhKvBlZsKun5tv3PB31lA
OM4q8xea2vxjNPL9YY8Gkb4x2VVOIv+EulptweFKdxs8yVCWUGpmaBSOpTb+xjBS
gIBPlKo24oVnTleOpNDSkpnLeHVbcB/ZIX6JYWYQEPH8er33YC08M8KzYPpLL6G7
QxGL9GhoEX+MeWEEFUx4n8XkMx1nRxCSM+fUirmcFwP63fTGjRe8RnXQPAV7icPR
MhzDw0COw6j9uxiWtmDX/4zoKuqNNuNn+lFg/2R4E7dvX9WxZgLTQZeE2h4Gwi+4
euaSElg8qKTtMn2CJGHnT5brzF8flwRERuFx8QjKsIkl7S27bMIJL+OngPD8gUgY
/NE+II+zUyFpa8YE7o7B+J6iaqNNB7nu7aAb7UotCm3PB5oBJes7/hduSYm6r7uA
AjQmyjCmVTnCpTNpfgk8LIjHwH1nitLxmcZ3BdpoaHI5iJIvA++5Of7JY+rlvE2K
1/ZopB8hY3taK5QGwQJFBkfI5sDgGEYOzBQOynZ2WsujHpfuWqz7vEDJKXBQ7cAa
vtgxLbtpBC3UcHsll5MDp/cUf/YM93GOiz2+25e5Wbx8oqP9eXa83utqtu7ZHS6j
iDDnANRkGr1D7UaW6W/cKstWJ98mHm3ftWPWUZRZhhNjVK4LAO3TYrFxw9fBTPI8
1XdLgD4wQXA5vbXkN/b1fAReuLhNbw3KRzVouQ9FGKHkS+kzt0vUIKkn0kzw6lHQ
79rz9H1MC4dHmVrNgfZNcFQzLspTtJib8i2I90hwhEIr01WZwCAIzImFNM5HmMMp
AdGCnbC2C3CBTw30epaXo4rvn6o3MJjWRRSJTUbCVqyONa4DGr+NfIlpSLBXLJQR
cmPglnC2b/3M+KLrBz1hK7YMetEJ5RMbFNFuarOAiqNj4sKjcUVdIKJ+g1cSxi8l
K2t58FbkxgUgwF53g2t7ZuIRbV2EaTpmSb8dzmDy9aGBJU0/yZYqvzCCh3u0XRQd
ktPh7WSv76ZzgxBZVwNuVVLcxR84zwAHNbaOswgVK/gQly+FusO+n6DKqD/vKSZ2
B7I5rzX1BKay+d29SjGN1QofVJo64+SJ9fCQvG3x9v8R2gICsOLFgb3Oo5O+kxk6
cszCWtFy3amQYkkBimzLWXKQeO3ND0WqDuwlSiWbsGrCyjTKBS9xdJr+XTiuFGBc
8Qd9ZoMMXvEU+tRL4000Lg5YnQ66IE1QnYslE2iq1p6rCQMZGbscwrUlAWg+O/ZO
XVDHPt+wcudBFOkU8cnerAfP3oc2UHyfRnBt86+gIQGIAjwy6gQvqDSvUfFdiERy
YbKTpF58xEG8A8sGlUdafJtmRXUzw3sDXucUVuEjilrx5WSH2LrGBusUKd/wUvrH
RMJLYrXnxFTeN20aU0fcRhVRbLwj6crYcDqACU7ewgFLl1y1dBTRvYDA/7DIYGyS
9mXqmTY/CFawSp/fKWcXXeOxxvnvBUYcw7WJ5i5XEP61B7AfWMEHjbWiw8fX2YEn
cGaalaSxnCD8zpL0Qj+l67NwcUHLSXpgP0DyuxpZeZIZf7+WaMbfrxU1IQ7lEEF6
RkZX6t6B1Mu/g+vvWmEjIUXzW4URfpYbrYQDbXP4Byk00RI0z3XyqaDEZ5R0wu03
h8b5mMkz8ZHuP34QSrM0+weeKu8k2DrdLzascWBwFfsukrpMWECEARpSw9KgaJ/C
FBsfg4FYlOefbhNNH0xXjGKrBqrl0UJoq9XoMUGr11BzbVKh6oRT2tDG3LYnuq/G
G4KD7fHi+Q9HHL9yVMNH6TOVEglTYR9ywyyrIT08lZy5aUBwiIGT5My32a/mCA/T
/PpU7OyGovMO1WadHCh06NhksglJoNHOKN+Q3Q3nwQM/g/R7A6B2Pgf/o8TSjIfE
0x0Joi/5RcEVOLlxd+e6Um/C2k/s5VToj7LpzNoKE087V20BIcKZD1awm1FNCExH
CDDQe+nA4N9pVHvh58zTuV1xm3Sl8ZrAg1lgdK70J/oIPP+BirAg1UwP6LaYsSWz
fO6du0nAXQXchAbNzskYnht5Z2KPvPupwW4+BEm0nkhhCcP92GYp2XJf0a7P0v6P
wLtZubLtDLffHYfkdHJTmUlsS+hAoWpKhhG8TQLq8pNm1QeoDbYKdiFQ1eF1IcRV
LOe6jrE1B+lyQhGScvDFrtEXZMsuMer1rNQjcIaXzkZqqEdAJ7eaa8NSDS1shitS
osdtRpiUU03YAHI/hNoA6Bf0M7c2Oi4zCXZv3tRXluoPRjPiPT2lEi6LZ+hEasQR
8qSoi4i15893OJNsCSR7UE9WQLwzDh4sEifbeH3ipZS6QV7umhf69f0rEA1OSLi0
G9ohDtBeYAEDdW4TCV3a4fwFKGw6G6/mcZD652A3W2XMFjfivdKH3qBgjUw7XHWW
GahKW+gl8zKO726l13Tivos4fDh8ca2Ym5tXseAda4HgWvwVoHkPINGuFWE36D0G
Vd+FkNFDu9yOX/+3+bELP8r0ux+e0arXurullTMfT7wpdr+Jxi/u7h/XGmRgLs5D
9e+x2ZiR/VPBgc/1dLtbC1Pa5f6jlertE4pcW5uWhmYKeb09wo5zEcMaxzyGrQhw
cQ/yilKfGtE6ObgLGjuLkHNDwFEewXBImZ1tS++XSLqiInp7MDwvexxH2PZD5T0v
WHu6AkB+IXj+IviPnPQBV5Gfact2ci+vwpW5TXlGxIOftYi/aHDr3UcwsRBMNSLQ
TXqVS494D0w5h/wkPXY8ZNtfJ4XeHBS/QX2gBxV0Vef1pkgsmHBiMM1/JsfEnO2h
k6z7ZHkQnXx1eGylWOF96VX6SXpJ65PghGIRDd0c2gbeA3UZZq64csLyPsH1EvfE
xo/2Y8cEJWwTGDIVxd7H0BKhMWoiDHJzqNHyuwe+HeUFA/Q91LAJuuiHZCVaXbVP
MtUIRfZ6Z2QhpOLaZ6ETP5/z94obq6kLvxeAVSKF/EAlMudQgi7ePCee12//DTbJ
3OR6cL2cwgKxLh8zTbe/eRnBfoSYOmfTVypd/6ETec+t7//Iwa1Uu6UbqWuDqvnk
LD/f1LVmIB4Vx5XhkGvcjkd279VOKUoNZPMHuf/2FAJTL6itunSn6i1e/N1c4Pc4
fT1qK64zmXNDzErFkZmbQsf4ywTH2nF74cz/SuEgwDR3UJEtsjUIrUcuzMb4HVfE
zg6cu4I1mBXvMH9o8dZJs3/3rnwrQPuLcM/sksIyKXZ9owAOMKjHEY/77PLkcX9R
SJnd8rim4aO2rD9L5GLcXjZaDlnfdbvaFUNTKvDfK7LXVhijEX3YdydDtp+yu0p5
QvbGLXZGsJwSPVJK1jsHkcrtfVXWcy5g0ZZRWnqPwwSzY7kFxF6HzWf7YEwv322C
k9Du4JBqycTKrrlaIK+svqtnh+wc81xkReA8cqgOFhvOmjQ/6HeIfL13h1Cv28hx
L1DA9sgiumirLN820bfwzk/sUBlOIhLmrcJJtlFd+Vt5Emv3AWNrcEj2geLQs2ct
bu90JnN7jbXc9U7UqHYd639ADUBAUfJ/mUzIYp73p+VVnFRHCFbuufPVCXkHsVwH
UXfv5Ef8l/O0tHEPm+EDkl4b021RqYTBEGcke/rOS+jeC5Tr4tPk9KVu0XlrBUue
yTDJQyn/nhIeLD2e7IDyHsi7o6wmsoke5ZLIp2B/SMXXw6wZ0RmShUDIwT+DOOBE
HLiqPaRxPaWlTijXDPfeCKidmHqfQC6vvYeRAPQx5EC776cmuEYsuChRuS1WjBnu
00DUZro5ctTJhfaaUsvwQ3b/jFp8aeubcuI3w9aADIoJn55FbuTI1AxluAiAjJEf
QvLFApwxezkUEYrFd24/1RauDUG4cJfvNNArB1ZJUOrDpHUFnItgHxeKlv+bnp5J
UXF4bkxWqyV2MvcZPS7rwTyZzBrkJCHAbqLtRY2yMCuPiFIRA9XO6mIprbj3BnCw
C1Byx+JmxIglC+ZuIF5GtLuHnV1E6a4Qptvfk2FUH7QsdFcC9X9a+nSu5Uufepkw
zGN0pREx47S8wnuCboWho8nkvuBV09NkwGPWP9VVZWaAADOxpPiYVVPi6CRxXG5U
aoa0npGaewMqN2lnQrEXZdW2p85kmZjWgaZt2w0eCsH8Yd2yET/AHxV98drgTKh/
fliCi2tyrQ7bAGlrxdBa9i7Ar3MR6EapNMj42KTh1FQeaVvsuOmF+vJAewHIezUc
IyBJYPz2HNG/HVjm9QkwQdPhzWMDlHicGYNleRaRpI5iT1X1yQqcUTEyZnB6u5mR
bMsKNC7rwpSp2A68hmDbU5H1KuzHyazJN6msjALMMolW88qoIkyIbJkbQ22VxMHJ
bSkNqv6ww/svUQivdLLpB1aTpIl5URpmGOasRZoZuCwfg1FdhtaRkQUUswhV3CvX
H/6+A0tJpLFwhVoI9ccMuxYbMCuh2MAigA3pGSbZE+Jc48iQ6lEMdQxhA36ajdhS
vO9iBFej4WxdFJWd0qsOORSqdsP5Q0GJBx1kLTlg7J3GWNEOPMJQre2F8Tuz2xec
NhS7NPowaYAPjV1fEhA4FgrRrgC5MuJQtzBTXuo+rMf7ldKAG08Uu2D05JBSjPHE
cb8QPLSkfCSpWH6QXhg//71gxsRwwm9K1SbWy1/vLmpbn9Y1MaVCLLzOdxejd4q2
HyX3q4uURC2qhAV6RrkJ/oFPS7f0RN/snV/nY6q0WsdH9yYQJd3+S9XZSCzdyAMR
SqPW+1MmQjSxNldSv4Z+DhirSiok7Sg6qGyal2n+tUamMc5yUmu47/iZR4ejV/un
hYeWkHJBGwKjY8YgFLhJ40jRHM9fgLrfnGuDj3uICgaoL+lQ5STjJ7ElYkoF3ouA
3d+3CCZE+mCZdwY7/+RAwE0+qRU3Z+BDn2W7Bmbt2JLiACtIWn9U+TTaTXd0mpFQ
/ayhfZ6GVfLD+cK85XYxCbkQQCqoPOpY58ppJ2oFiosh80lQFLgy/QOQnlYUbBrL
Ibsf1W7FQQvwqu/KE0VwIe4xedmQDns5YczDXSxYQWEHJH5WDNNO+mnc691wGTB9
f7taHjfda7+J68rXxYxd3Hb/ccft9uz6K5sJbtBdJrsK5xiD+henyoF3SDM6gMDz
AB0MOanSqkiB9t0PfUlDa+sXB9Y/428z+ljH2adoMWZ3CFpvr5ozenbd8Js2P6IO
vWClzybqiS2/T9o9MqzMu65KQuBRV/lgfH6cMof0UoULgjxuflkl+z1fajsuVbJ5
VRS7G3JFgQYtoDMvOOkif/I+Sr1lbN+6gpFLt3iRXCUmH8lVe1ylA0hQV/Blk0Ik
PTgrJ9Tgdmvtzouf/YcdGCjqI2BcxxiYJBhbjwxtowR14SyDBx+oHFihtvSV28Go
M+NlpQxoV3Ai7tPTzNZ+ofj18N6EGmZiMFJneVgPJ7Luf15aaF7TsK7YmNsz8YhS
ExvNQskp3LO73CiwB2q3i21DnFT6615QWoMhE7mgnzO41IzLkw7h/cRwSIfZj+S5
w+HdUU1vIay0lWWubsglqFoJakqhH2edCXPxGIhswZgXCvrTsIB+XA3HjJ3ToAHw
b+GEgQHXA4RHCVXcEH23uwY9XQ+A3ubUldD9aXtxfHkypTfAh12fmQ7pNsHqzEE1
AQugTIVuuzQlyPq7Z9tcT82Ilae/5u/h60f2uNzhXEeKwp0016ra+yTH8bQAlPdH
MxCHTPO5x6sh8scXET4tgUkDaz3L8oH0oroh9DceNk8czGU2WorJy+WbOVI7qRiU
7ENiJkzC4xyc7/DU9OLF/92PQXfZPwhJDUQ5xgo53YLyOUEVlr49Nb4Gpe+/wSMZ
gS3GCs1q9cxf+VYZKjZixXvk3Z6eoYeskHlVyPExmZmrYcZBRoWZR8ShVQOQoRIG
rJl6ibOYYSRMEZR0zJjqv6Sj1yy1vBdsHcY64P+N8l88BTSk42WHHjheSduQCHRu
0duu+kigzMbJ6jORE0xyhronCAM8Ns1Xmjz0NWbX+jwlf4r7rR6o5XbHnNqy9wW+
J67njxtQbjTYbrrxCsG7MSYeBqmhAKPNbtgFL6xoaAWkdkMZDh7A7GlsJtKKXR8b
jZEN+Nh+7jeDFCbYXRkWDYu2+F+ykC9kfSePw0VRStNkzfEtztP75e7NDVud5+KC
hj8le/vNi+0w83qmX9l/jxMjlDCmdBXQbxhM3tUHM2dNu9wo/ipiPJiNFE37wX4O
pojBqwQrqD8Z8wmdc5YjGoFbRq8ALDYE+oocyGmHUr1iTLrcfrWcgbIKWMuxkR4+
uMn4sg3cuxSV6+4X8PEJddjGMywo/7MCOUy5Z6vzrlb5KiNnCiDdoRrTEBAbmAsd
djt+0HDNruO6r+MoaM18hebw+gNmprgImyHSXJwYzmil4yCx17dgvrfE1kE8Dawf
uF+tWFC9hVb/1F7p1syPwq8e3/b2V/vY3ArA6haqQHO8dpU24h2Jw3g0Z1Qj/Gxt
nTMqnNv5TBAF3CdjJ5KU2//q69AjZ0nPS5C+QCrOSEVDg9tbGwEmcuXh2xDBvF8J
swuaiskT42tROarQzWINmY9T8yp254s25fxCcWiEspRbO2vO9sC2AQxqu6+pKW/z
L8Gy4mLOxIrYSmYvSsd4HecUwX2Dvn82FQ7N/e+e4zfVte7/wKQXrMU10aAsnu5R
mkdsZEA6sAU61fTPL3IA0BMca7swepd+db46eez2QgNMslUqrjOuaYMNz6n9HRM6
njoiPdF6PSqgFBUZjQFydb3aAkFi9XXy+FHLR89d3EVQoJRd0efbfyC43kkF1NFw
cPxPz97NktBOi2OvyB59hRLk9SFU5cyYKlO0EfDX8okSeX1vaL1SPBQ5WaBUcGNA
bst/XwyHxSOq8oNnDZTZyKp0x9JZ/uqDXqlnfQTq63yP5CP9qjRi/Q3j500+9HUz
qfoSNYyVjVEnZlvYRfvK1JjYjf2peZtsT4pdcohBMUBmPyb8tsLmDWLEI9H65Y+F
DBRtp15DAl4KBHNYNiDzNjy31sA160fkQsQgf7K3IzOsGzsp40Yd7XCXtj8pSqZK
h7zekoQQf6/NKy11sl8/55wi9QU2VjHVTkinNzvkoe+tNQVUlyMiX98WUXQZFN8o
0lhfMwKjI/qo6QpGh2K9/L9MPOQyj022qTTtWL1fEpnXViaD3HxtzADR3MbUPb/L
iilAgxg9olCq+P8zWr0DriTmCeq+ybhMVcfyRWUuTR8qb9AGQx+KDLTYBB+fhxKP
FMRxVdNoTnnPjoTeZNmJjwAMmyN8Rte8u0IBWLT8ejW5r3eMdnv1BFemEkRdYHg2
LRtkqcx9aZPL0Pv0BuMl98f5RfK60yJNjLL4DxyxF64zMsmzrLJXpk6X6vGHa6rP
ksN6z6bkP4H8HsCNtL6YkvJSuEdQnGlr/CCg7KaMWHUnBx5wxV8MTCi5wOy+M+hl
wPfNqs83PdK32+LjNBOxCsso7U4AI6wlaxNb8eiI4KRi1F8uQ+zG6dPupojd5gxV
I4LyHS4W9sYlA762ThoqorWTKl03Q/3CLH5UZBfwW/YXLVplGk/3ksjpcolY8zjI
MsBwl6p55kBxqDomGcNAH7ip4gG46VQoWGb7M21VPD6PpzXpkXQhGx2CcZteRphC
xPmfzGHWpMl2sVm5lP9Cq/bXjuAPQUUUJ859IbibLiDomAvDLpT+ZHz46w4E9Nmz
rpwjm1wLTL/N9R0jXe8p/xJaOAQGLclRyGKp266ogKN7TtO3or14IZi/VTj9s/k8
hj1IPcBiEnCT/Zqlo20EGXZnUA7yt/7JECZD2u2yFZc6kb3LyAfI7tjzYU0xGeZ9
gwo+sI7Ul6Vu792r7iFRpKwvPQVwV4wpmZ0/eC8ijBD03wTWP3+2FSuwCcKL4Zao
ijuSdX10e4vYLbJUFrpZdsiPGPNrRuyMlP7GuyUstKm+nogRwJTJlfWaEOl/8p3e
ZFZ5QKdwEn7L/CukD9cumE983F6GmLd6BKj4nykysnG/wBoWX0Y4VwmvshY6eTvc
0OTE8ZRJhYmn5pEN89DfQZ9VGm1Vjnvo9yt/MK+MWrYNYPW11pLjYocP9T/dFK19
1Fj4WYxpcrrSpm2OTVK2aFnTOfuWb7uXB7718HBl5j3V8BRhJwUPrquldzX5kVFG
dcve1UtxDogHtdBlHi4J/jQMvWBqrAdniFoWSa2nRhpgcb8laOmDflC3/YbU+6P6
kiVe+KyB/M/FBT9mSHdRSI8mGWgRZkhzYH6SCxctP9M+Stl0RWz5fEZ8qYrfQUkC
hZt23159f1U5uOf1ujTAEdEjAPwvT6EruaqR9vml9grcL1OBHFA6DAytkwd8Jm2U
8L9PVjDo2EgEDH9B4sMLzjqz8hDAvHw14JwvS7xu/vO1tTvsT5Zdq6OMxPkFqIGS
0LgwNVmc4yFhs+1KFHAjLNVRfA8cscpeGA7J/Ac7mIj5ZVtz6EEvoEiiPEhWMQcA
+lholhtaDXV2ImLYAzJsGnAvgRngobCMDPGAEJ0VvG5u/4iMvpdBMx12TeyGLRi8
Z2NtVX4zOJJRBkfe1VL8BgfzZQX5xKUTDMxshT1HfWzx+oudcu7LfatYsqAnGPCp
n7V/PCDE+QJNNXMGnBc01rDhzlVeUllAFg7qAySNn7GmR/W9SxvXc6yoJJeHKZfm
8h3/7K/Dn847a7sdWv0o6dJPU6xXHolzATXCMEVJTMw5KOkG/PUgmsvn+TeSaMbW
6ARNzLipeW9DoqomOLWSDUGqNCfuxkioSIQvjA6OyvqfrQnQAPKkEby2NbQi5gN0
LX150tNA+rlpme9r9JHARO7gz1IlUT8X9091D3V526VpgzVcBaCl31C3WUjaHfAW
C6CYqtds1a0SC221uffZpACdeqMxGYOqYUGfok8HX3X+Zp7axhfvg3z1pNV8qMUG
0GvA0dQHIDx9DoP3lRy81+AGCG+RYtyRXZWiDaLl+W2dJdFTd7dhorX/mBbymMue
jeW8CSVHDH1ZsEWljNCN+qCknznB9ZLuROH54Ncn+o2G5e0CajL1a49SeH15n6/G
OITG37aX5pD+ESGhSQvUl87QHywIYEIRku7jMZGeXKiOd/bBM1tAIz/h0pMfD3qo
hPsOEoJY93+oIkdKcdXW7hSIQeSH5fiBwv9gotQri50mAqQxZtMfGHm143rirtwV
gn14rtUSrg1fEOHjch1dCaOJbXs+wFZcr28RYfQrNez5UB5rCoRYXcgQUCHmMjgl
3GUhiwAtErcQGB7RQ4ittBBlFqK1xftbqpMZSLIeR8iBLNyvuA8xPeE3ygLljy6j
o0WkEFpAROcrLL8+roXRCDNd9TinqKGs3Mu2kHCqUjGqtOaGWbuMCf07ukQKFkYx
0vxv4b7KpWqRXF5jVzsXDAsRl5qxyvyGTS9L6BJM0GjOq1L0xMk0Bz1iGPTqg+z9
RcLEBXXgkUkpLPrFouC77t/5PaPSshFze0COemsbwyn59lmYoT0zJkH62DU+EzTv
eZydZodu5ogFZylbPmguw4SnL7aMgnJvuKcxyTnElgTcxazt0t6NlskMl5IeAyRn
t/ydvt9KHzVmmzkm/SV8p9Ty9aaQ72UgjtCbBK34wsnL1uQNHs92E9zl84TBKr/c
sgPMsHUMd3QzvXL6uFCmo/dH8UpUifEcDvubv4F8CXzEOFXjzQ68ikRTq0PoJmuS
WmelddmVzR0LxnVqeRLobAJv4/CKw3Q1n+4mdbvFe9haXHOmRK6dbTECFAnn7Jjp
9IT2I2gZzPe71ZVSaQFLk0I373iLzpEhfCT7mXzPaumGQ2iE0/Ne6san4dpBmvEB
e05WpBM+oM1UPEBtptkSsUO4wXckr8/zMveDlDBKPfpBiSF0pIbC9BnBKtAQi8fB
iDomlwyPJ9P6syGOptP+Ke1sB55D1tyluh4B14Ehls8qPK6tKN34LKRJ7OEyaRpq
OjCkisK0cedFPT/S98hoICXjQfKVjDCLsbgl0E+T1csdjtrmOfbTC9TdtrNgOQ9k
XpUYKxlGc01KvGoUoiz7hec+M2x59Ex1PUg8jG5tACzZiQRgXtT+JlY++JhQb3li
h5IOiTYGoAk2thfrXLt6kWSCsstt/DespDMAHclkgGp+/fME/cFqsl8PfaGnj/fx
iAht2MPuZz5srLqNNQCa67+v4SM7kjLU4xiM9dwaXIiJ3wXf7kdd2HRVGiM/zh4a
8Qba/zLcFeBAzQGESeJgLg7h5o5BO5rCFC/nNbWJmM4n64rd+ViNSWeAkGBB5EFR
O1pV3h8lDqxBE+LdrftwP8KJbeOjPT4/y/98hAvCvo2DqKJvWU53UZodJK1w2E/5
+eFpao1L/gzsGZ1tkqBVtdLoQjpiTM+GyU4XMVKbDgNvXS8tbEapEPXnrOByjx+M
nP9+3qd74jvjAhdLkMlGCzSZt9v+puHqb9rD5BKgI2xu9YsmcLWa7HAxkf/LBpkz
+j6qVTbfuuHU/eVomrRpKBeS9Dqvw1Fka+vcPmppVwaO9goyc2/Pnf/9RlipYSUB
d52Nqf1GBx5OWT6QpoeGMQnHBv/oFd12tjXi1tx7P5zaqSrBtn2v0o6XWXyfn0L4
sWb64b5FX73/+VE2EnbcpMA6buHFH0CHiV1UpSu6CPZahdfO9Wxpn6qJwueQOYGs
ty8LnxPC4jxKdXB+BKaF/bONGLq0qDuBVHt6db5Mx4Ce7gJXjcLUFM84Sa6cmK1e
pJmrERGpLRXzL7hDr6ndGRmHUFgJC8D1Cvm65ZeGxqVr3ZQYSN6LW3MUuxDkWGtB
kW27H21n3RZskQ7XIU0J+rGabdLAG0n2X6hbm4cnkl4tAMe80xnRuXARxLXgKcHg
xqRaGGUWOc/bDFbZ2xMwTu1jlemeN5UCLfjKkDxmes8LWkCYUxNsZq5Bl8YIuw8N
+soEJ87b68MaIyhLM7/RBfuPRBLGWwCPNlSjJQEoGjUSVQCUg2kbXnP1d4TXjFuT
Cr1QNbAsfzgd0mgsGGiOq4dlRJ5LN/YnUfYkDqaWl7kUSVTkugdBuEHFSoF2Y2lK
/FC/IBqGLT5eMcnxbASkbjj8+V0VRtZJHXCr+f7Xzd4zFafQndaoaulY6yB4CyCx
5ygTeGNO5UgmswnkzA89hHCRzxaWdbJOppcXwTaONuQzGVbqSkHQhYOn0Wq/+LsR
kyolEmVkSIjKaENgCEhrYhQRm3U+N3gqGlgw6BrEUdCA8EzKlMZNL5Xm9/Cko0GS
lhTL9ysBQCbwPL2lg8sO/DTGHVuqicTMu9WI9mzdeoWSBk2cT0XNGrRgmmYJR6Kw
TDzrNpjJbw5QU+pgu23GFbdJc2efu6RY/zujHYeLwq8skNye3nWYYwd0YGI/YEnr
XhmOVkVc3JlZi9IGgPx5E+ozb8/F01hQY8cyCP8qd6jUWpItEIagKSKB1f3G0U0C
VGOHKbsh8rB+d3AdcIN6tdapXtK4tIQgPbIEec/JTZn0JL4ji3pEaUy+sRRAiD7j
r1RY2n1euHJizmWSODESQ9rn9Xl4zj3FIe276jzyMLh10SXO/WzBvoU1GY8wx30U
WZjecdnuhWeXeSGxEGlTGwn4jGr4Hj0fA5Er1eKfVLoN9+0dXxmcyeKDi3Dk73GX
KDg2WoMdRrHWzIoUAQjh3qlLBmRm/UTnOdJbIf8Pe8pEp9edNmLopB44h7v8+RX1
/z2umip3YfVB9l6N7BCnbcgNjfwRGtnglPMJNz/BzZErQSWk24BQ2gu5iwKoUHFC
vIGWI2X8IPaRZUQ5O8hoRcCabsa8GRHVFQpCVuaBa0HpEjU2IJofZbC952fuvtgc
WiWEpE6mH4taJWuiCRjvC7BsdfSTZxSRRcMkeyHa89aTB+Rcg2B0KOXm5y7asb9v
o/Zdbu8IBakvlaJnHlkSWYLlb/ZdNdZXsWJ5s6jc5OmRcEKtCqSfAOUlxuSB2oFe
zkKNn9dX8p7sx0McrZnvu0x/F62aalRKICO9uc/OXMs2ZVio1vKiTzfLvZKXEO1b
+RCle9edUzz1G3o/UMuA//Y25HDo+304oPz8CoqEH2tTE2nS9IkVn3YYtfNDyWQ0
U9iHg/vzMq4ye4Rbv0trKdxjdpgbNRyg+NDFN1vfeebTqNufspjp8IZSvobO8rOi
lJssvOSB8qKZTNr/k0MM3YWW/b/J7YPWojr0eMi2hAjCCJebY4PeiKryIscmfu1+
y4xtYSqi8EZkTx6BoYMm+hO64TWTvhz4S8g9igDgiU1Y+/Hv7csYRBIVpLSaIiUz
UnORSmwN5JhxTAuK//T5v1HK4klM+D5Z8PurFhvnhOsAzZz7GBpl8SpRDvxnP/Rk
2YgU8dquNHm27AqMEwpDvqBmABxU9K3lR4q3yx3GA8yMiF5PS/ZxBDa4uohXh2YU
YABEZPD5AtjJd77dp1g20vZWRC6m5MIlp6sxjwBZg4+iGXsLTvv+sFWM5wEj3ghg
HMtHEsMBb/8XwysjNVquHZY6cK4+DnaSakRIe6vE27ThXddpweqpGUwCN4VC+PHW
P7SKngC9687TN/UHQfCQdQoegQJdRPQxVpuJejgtXv0rpd63QFYCDi58lulTKm8R
23QD/jdUU6e6NiEBgtSR+qMO5dFLyDIS7PhyCSiVAqF7+d3IpTiT0Ylt98SqbAZE
4EYW48YC0MYUQ/qoDo19vMpZkzRMr4rE8vR61aa0zFh8rEXOq7QePecAC/1R0MNX
Ct9dGhqlDrDfWuAQSceB7g+jR+fKwmDTzGsRaaS4xcp1RrI6N+HDHZJG8tKxfy9K
jMHPddL4UbTXc0tct2ayUQ6XNF+0XUyLLRMeiL3cPbcsPX57DEDQ4O24295u+wSZ
XHY0Am3hoT9ns3W0ydtHB1jVd2po/HVjjOYgaRIiihqZvvd+7wEodfs9DtZg7sjx
p+tGAEmHQTHtJEMZ/6syTsT4nA2UNFAYca8nVOouK09otxIYgcFsYB/j3PzMhTXk
JMDwYJz3B9sz0Vf60tbb2Qcm7adw1huuovf+sPpjF3jGtQ5/yu/5IHm1jLz/8HuZ
CdAGmf60dWJ8Zr0tcchr4l6VaYMbnDgUbEuumHGdY6xzojvBYCxfu7niKgmcrWC1
Kw4bmUmUgdzcOeKAxVEtbuIxvkxl7MdSPaYe+mGqu9pAmVeoGprD6uBgTW+P+JiW
wS2prUwJXSOiyxuzgzeW23AyEVT89tY0lBS+B9S2oYPXh2+57QdgLyby5ka98n/R
2quIwM6JZ4+0XEqi2G88BAC/9ELT1wBAEx1g4EoeB5aSSVdEMjZ3Xd0uq5NIoZhd
QPn3WeHk6cVpPcJbRXwLoB7KrOMhb8SyDRrQfiuqVQtY78wRtIPmV1MYCnUBuPAO
YEv4GSpZlljhf4bC/IwT05Eaom+cphdfERDVNQL4r2A9xvKPYmlol4tSku9VLxVK
IBy5UNzKR8brGHZeJFtKRQH147iilmEaHOimPNqZ1Zjmm7WIsdOLDg+Y/cl0WoZD
5YkcNCJaY1NZFK857hKb6vxY3/kTmHfMheDuVSPO8Lt1vWGS7PjxY7t8FVpjd9Je
uvT20gQMQRs60+v07dWrXWxZ16qLFktm/W/8yHsm4fKsnsBjv8jHM8xNLUQOkJIL
1/BVUKFjG2lvMJH2gzKK2QMpKP7LxpNIU/H34sRXA9BpoFe+0Snm/u1iPivB8ok2
KBAnB85E7hh+r7JE0qc2hoelhfFfPF7yFvsWmV+BtlnZ369fKKlF0fCKA4x4eamo
yEhbfaEa2yGUk8I91bzlbCgQe2vwjIQygo5439E/AptJSUmWrFK0bA6Gnsr/IOo4
78Yt04dObQ5rehj7BW4WB9ZLVneS+Q/vpTJcLpEy5PpDJrC7yA8osdlXXHPSS09a
mFdPPHsNJsGDQNAE1TBTohNC1uBpUAErinkGlo0ZOKZbkuw2YwlI8N4z/meD7jM5
L4zTOqeVyCwltqMdtJoLBNcntlsDuO4nZfCSib21KKmV0MCQ2wkmbM5uNlRH5cG6
TR5LUZnblTG+aSOMW9pvTaD4WkPhCgWl/BakbeU6LrG7vZb9qIBSG37vTUd1YrPS
JExag3QXjQPSVkFxmkb2H+nRk2vu0lDu3SF8Lapeb/JVSHv3Zikx1ohr3Gi5Kr6Y
W9koFBNeWJ5rDQpSR4nLb/+WAYVaO29+n7cX8v5w4WB6tzIUJDg93OXDxcYqIQSv
9MT7ZuITgHfn1CwhEDrjrXzmuntnOXbJHZK+mZ6OAbK/hRjxGspmhMSJlMfuHKC5
s4IAFZ3V3rBoqeLRZgZ/4UFuLu3B6TE8MLC8/GDs3w6L9f5duEwML9zaYSDT2MTv
ke/OOZkAy15WFfAua62tvZa+UKy02rO21RC+NSDZVQShmRjxSm5reEwaha+l3lB6
2Km09Ij0tYGVooAoUxchigGj0AAqqDQKYBDdsKLmUI8lre1kfsKhGbhF/yzoCrIE
vk3+R+Gi1FN7nY6g8hfqXoMxRJ7GEYO1yZYW/j+hczDxE7qa2aFcAAZ2iPHr5JVv
QFGjz4uZK535tVh78XNnmQQJOfU0+c/j64VisQgcUkE=
//pragma protect end_data_block
//pragma protect digest_block
uQ2LWSE4vnedaTbHZfPGFc6yykw=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
