

`ifndef GUARD_SVT_AXI_TRANSACTION_SV
`define GUARD_SVT_AXI_TRANSACTION_SV

`include "svt_axi_defines.svi"

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
`define SVT_AXI_INTERFACE_TYPE axi_interface_type
`else
`define SVT_AXI_INTERFACE_TYPE port_cfg.axi_interface_type
`endif

`ifndef __SVDOC__
typedef class svt_axi_transaction_exception_list;
typedef class svt_axi_transaction_exception;
`endif
typedef class svt_axi_barrier_pair_transaction;

/*
`define SVT_AXI_COHERENT_READ \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == READNOSNOOP) || \
  (coherent_xact_type == READONCE) || \
  (coherent_xact_type == READSHARED) || \
  (coherent_xact_type == READCLEAN) || \
  (coherent_xact_type == READNOTSHAREDDIRTY) || \
  (coherent_xact_type == READUNIQUE) || \
  (coherent_xact_type == CLEANUNIQUE) || 
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == MAKEINVALID) || \
  (coherent_xact_type == DVMCOMPLETE) || \
  (coherent_xact_type == DVMMESSAGE) || \
  (coherent_xact_type == READBARRIER) \
)

`define SVT_AXI_COHERENT_WRITE \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == WRITENOSNOOP) || \
  (coherent_xact_type == WRITEUNIQUE) || \
  (coherent_xact_type == WRITELINEUNIQUE) || \
  (coherent_xact_type == WRITEBACK) || \
  (coherent_xact_type == WRITECLEAN) || \
  (coherent_xact_type == WRITEBARRIER) || \
  (coherent_xact_type == EVICT) || \
  (coherent_xact_type == WRITEEVICT) \
)
*/

// Transactions which always have 1 beat even if
// burst_length indicates cache line size.
`define SVT_AXI_COHERENT_READ_1_BEAT \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == CLEANUNIQUE) || \
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == CLEANSHAREDPERSIST) || \
  (coherent_xact_type == MAKEINVALID) \
)

`ifdef SVT_UVM_ENABLE_FGP
class svt_axi_thread_specific_svt_pattern_data;
    svt_pattern_data pttrn_contents[$];
    svt_pattern_data port_cfg_exists_pd;
endclass
`endif

/**
    This is the base transaction type which contains all the physical
    attributes of the transaction like address, data, burst type, burst length,
    etc. It also provides the timing information of the transaction to the
    master & slave transactors, that is, delays for valid and ready signals
    with respect to some reference events. 
    
    The svt_axi_transaction also contains a handle to configuration object of
    type #svt_axi_port_configuration, which provides the configuration of the
    port on which this transaction would be applied. The port configuration is
    used during randomizing the transaction.
 */
class svt_axi_transaction extends `SVT_TRANSACTION_TYPE;

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_axi_transaction)
`endif

  /**
    @grouphdr axi3_protocol AXI3 protocol attributes
    This group contains attributes which are relevant to AXI3 protocol.
    */

  /**
    @grouphdr axi4_protocol AXI4 protocol attributes
    This group contains attributes specific to AXI4 protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr axi3_4_delays AXI3 and AXI4 delay attributes
    This group contains attributes which can be used to control delays in AXI3 and AXI4 signals.
    */

  /**
    @grouphdr axi3_4_status AXI3 and AXI4 transaction status attributes
    This group contains attributes which report the status of AXI3 and AXI4 transaction.
    */

  /**
    @grouphdr axi3_4_ace_timing Timing and cycle information
    This group contains attributes which report the Timing and
    cycle information for Valid and Ready signals. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
   * @groupname axi5_protocol protocol attributes
    This group contains attributes which are relevant to AXI5 protocol.
    As of now read data chunking and unique id identifier is added.
   */

  /**
    @grouphdr out_of_order Out Of Order transaction attributes
    This group contains attributes used to generate out of order transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr interleaving Interleaved transaction attributes
    This group contains attributes used to generate interleaved transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr ace_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr ace_delays ACE delay attributes
    This group contains members which can be used to control delays in ACE signals. Please also refer to group @groupref axi3_4_delays for AXI3 and AXI4 delay attributes.
    */

  /**
    @grouphdr ace_status ACE transaction status attributes
    This group contains attributes which report the status of ACE transaction. Please also refer to group @groupref axi3_4_status for AXI3 and AXI4 transaction status attributes.
    */

  /**
    @grouphdr ace_l3_cache ACE L3 Cache related attributes
    This group contains attributes which are relevant to L3 Cache usage under ACE protocol. This is applicable only when l3_cache_enable is set to '1' in system_configuration.
    */

  /**
    @grouphdr ace5_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE5 protocol.
    */

  /**
    @grouphdr axi4_stream_protocol AXI4 Stream protocol attributes
    This group contains attributes which represent AXI4 Stream protocol transaction fields.
    */

  /**
    @grouphdr axi4_stream_delays AXI4 Stream delay attributes
    This group contains attributes which can be used to control delays in AXI4 Stream signals.
    */

  /**
    @grouphdr axi_misc Miscellaneous attributes
    This group contains miscellaneous attributes which do not fall under any of the categories above.
    */
  // ****************************************************************************
  // Enumerated Types
  // ****************************************************************************

  /**
   * Enum to represent transfer sizes
   */
  typedef enum bit [3:0] {
    BURST_SIZE_8BIT    = `SVT_AXI_TRANSACTION_BURST_SIZE_8,
    BURST_SIZE_16BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_16,
    BURST_SIZE_32BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_32,
    BURST_SIZE_64BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_64,
    BURST_SIZE_128BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_128,
    BURST_SIZE_256BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_256,
    BURST_SIZE_512BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_512,
    BURST_SIZE_1024BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_1024,
    BURST_SIZE_2048BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_2048
  } burst_size_enum;

  /**
   * Enum to represent burst type in a transaction
   */
  typedef enum bit[1:0]{
    FIXED = `SVT_AXI_TRANSACTION_BURST_FIXED,
    INCR =  `SVT_AXI_TRANSACTION_BURST_INCR,
    WRAP =  `SVT_AXI_TRANSACTION_BURST_WRAP
  } burst_type_enum;

  /**
   *  Enum to represent transaction type
   *  NOTE: IDLE value is currently reserved. Currently not used.
   *  Note: ATOMIC value is used for atomic transactions.
   *  Note: READ_WRITE value is used to represent transmitted_channel for ATOMICLOAD, ATOMICSWAP and ATOMICCOMPARE transactions.
   */
  typedef enum bit [2:0]{
    READ      = `SVT_AXI_TRANSACTION_TYPE_READ,
    WRITE     = `SVT_AXI_TRANSACTION_TYPE_WRITE,
    IDLE      = `SVT_AXI_TRANSACTION_TYPE_IDLE,
    COHERENT  = `SVT_AXI_TRANSACTION_TYPE_COHERENT,
    DATA_STREAM  = `SVT_AXI_TRANSACTION_DATA_STREAM
`ifdef SVT_ACE5_ENABLE
    ,ATOMIC   = `SVT_AXI_TRANSACTION_TYPE_ATOMIC,  /**<: ATOMICSTORE, ATOMICLOAD, ATOMICSWAP, ATOMICCOMPARE */
    READ_WRITE = `SVT_AXI_TRANSACTION_TYPE_READ_WRITE  
`endif
  } xact_type_enum;

  /**
   * Enum to represent phase type in a transaction
   */
  typedef enum bit [2:0]{
    WR_ADDR  = `SVT_AXI_PHASE_TYPE_WR_ADDR,
    WR_DATA  = `SVT_AXI_PHASE_TYPE_WR_DATA,
    WR_RESP  = `SVT_AXI_PHASE_TYPE_WR_RESP,
    RD_ADDR  = `SVT_AXI_PHASE_TYPE_RD_ADDR,
    RD_DATA  = `SVT_AXI_PHASE_TYPE_RD_DATA
  } phase_type_enum;

  /**
   * Enum to represent the coherent transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    READNOSNOOP          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOSNOOP,
    READONCE             = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCE,
    READSHARED           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READSHARED,
    READCLEAN            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READCLEAN,
    READNOTSHAREDDIRTY   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOTSHAREDDIRTY,
    READUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READUNIQUE,
    CLEANUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANUNIQUE,
    MAKEUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEUNIQUE,
    CLEANSHARED          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHARED,
    CLEANINVALID         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANINVALID,
    MAKEINVALID          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEINVALID,
    DVMCOMPLETE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMCOMPLETE,
    DVMMESSAGE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMMESSAGE,
    READBARRIER          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READBARRIER,
    WRITENOSNOOP         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITENOSNOOP,
    WRITEUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUE,
    WRITELINEUNIQUE      = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITELINEUNIQUE,
    WRITECLEAN           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITECLEAN,
    WRITEBACK            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBACK,
    EVICT                = `SVT_AXI_COHERENT_TRANSACTION_TYPE_EVICT,
    WRITEBARRIER         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBARRIER,
    WRITEEVICT           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEEVICT,
    CLEANSHAREDPERSIST   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHAREDPERSIST,
    READONCECLEANINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCECLEANINVALID,
    READONCEMAKEINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCEMAKEINVALID
    `ifdef SVT_AXI_CUSTNV_ENV
    , CUSTNV_L3PREFETCH   = `SVT_AXI_CUSTNV_L3PREFETCH
    `endif
`ifdef SVT_ACE5_ENABLE   
    ,WRITEUNIQUEPTLSTASH    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEPTLSTASH, 
    WRITEUNIQUEFULLSTASH   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEFULLSTASH,
    STASHONCESHARED        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCESHARED,
    STASHONCEUNIQUE        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCEUNIQUE,
    STASHTRANSLATION       = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHTRANSLATION,
    CMO                    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CMO,
    WRITEPTLCMO            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEPTL_CMO,
    WRITEFULLCMO           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEFULL_CMO
`endif
  } coherent_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  typedef enum {
   CLEANINVALID_ON_WRITE = `SVT_AXI_CMO_CLEANINVALID_ON_WRITE,
   CLEANSHARED_ON_WRITE = `SVT_AXI_CMO_CLEANSHARED_ON_WRITE,
   CLEANSHAREDPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDPERSIST_ON_WRITE,
   CLEANSHAREDDEEPPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDDEEPPERSIST_ON_WRITE
  } cmo_on_write_xact_type_enum;

typedef enum {
  WRITENOSNPFULL_CLEANSHARED = `SVT_AXI_WRITENOSNPFULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANINVALID = `SVT_AXI_WRITENOSNPFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHARED= `SVT_AXI_WRITENOSNPPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANINVALID= `SVT_AXI_WRITENOSNPPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE
  } write_with_cmo_xact_type_enum;
`endif

  typedef enum bit[2:0] {
    BYTE_STREAM = `SVT_AXI_STREAM_TYPE_BYTE_STREAM,
    CONTINUOUS_ALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_ALIGNED_STREAM,
    CONTINUOUS_UNALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_UNALIGNED_STREAM,
    SPARSE_STREAM = `SVT_AXI_STREAM_TYPE_SPARSE_STREAM,
    USER_STREAM = `SVT_AXI_STREAM_TYPE_USER_STREAM
  } stream_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  /** Defines the atomic transaction type */
  typedef enum bit[2:0]
    {
     NON_ATOMIC = `SVT_AXI_ATOMIC_TYPE_NON_ATOMIC,   /**<: Value that corresponds to non-atomic transaction type */
     STORE      = `SVT_AXI_ATOMIC_TYPE_STORE,     /**<: xact_type corresponds to one of the Atomic load operations */
     LOAD       = `SVT_AXI_ATOMIC_TYPE_LOAD,    /**<: xact_type corresponds to one of the Atomic store operations */
     SWAP       = `SVT_AXI_ATOMIC_TYPE_SWAP,     /**<: xact_type corresponds to Atomic swap operation */
     COMPARE    = `SVT_AXI_ATOMIC_TYPE_COMPARE   /**<: xact_type corresponds to the Atomic compare operation */
  } atomic_transaction_type_enum;

 typedef enum bit[4:0]
  {
   ATOMICSTORE_ADD        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_ADD,     /**<Atomic transactions AtomicStore Add */
   ATOMICSTORE_CLR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_CLR,     /**<Atomic transactions AtomicStore Clr */
   ATOMICSTORE_EOR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_EOR,     /**<Atomic transactions AtomicStore Eor */
   ATOMICSTORE_SET        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SET,     /**<Atomic transactions AtomicStore Set */
   ATOMICSTORE_SMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMAX,    /**<Atomic transactions AtomicStore Smax */
   ATOMICSTORE_SMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMIN,    /**<Atomic transactions AtomicStore Smin */
   ATOMICSTORE_UMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMAX,    /**<Atomic transactions AtomicStore Umax */
   ATOMICSTORE_UMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMIN,    /**<Atomic transactions AtomicStore Umin */
   ATOMICLOAD_ADD         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_ADD,      /**<Atomic transactions AtomicLoad Add */
   ATOMICLOAD_CLR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_CLR,      /**<Atomic transactions AtomicLoad Clr */
   ATOMICLOAD_EOR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_EOR,      /**<Atomic transactions AtomicLoad Eor */
   ATOMICLOAD_SET         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SET,      /**<Atomic transactions AtomicLoad Set */
   ATOMICLOAD_SMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMAX,     /**<Atomic transactions AtomicLoad Smax */
   ATOMICLOAD_SMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMIN,     /**<Atomic transactions AtomicLoad Smin */
   ATOMICLOAD_UMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMAX,     /**<Atomic transactions AtomicLoad Umax */
   ATOMICLOAD_UMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMIN,     /**<Atomic transactions AtomicLoad Umin */
   ATOMICSWAP             = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSWAP,          /**<Atomic transactions AtomicSwap */
   ATOMICCOMPARE          = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICCOMPARE        /**<Atomic transactions AtomicCompare */ 

  } atomic_xact_op_type_enum;

  /** 
   * Enum to represent the Endianness of the outbound write data sent in Atomic transactions.
   * Following are the possible values:
   * - LITTLE_ENDIAN : Indicates that the outbound Atomic Write data is in the Little Endian format
   * - BIG_ENDIAN    : Indicates that the outbound Atomic Write data is in the Big Endian format
   * .
   */
  typedef enum {
    LITTLE_ENDIAN       =  0,
    BIG_ENDIAN          =  1
  } endian_enum;  

  /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DAT channel.
   * Following are the possible values:
   * - TAG_INVALID  : The tags are not valid.
   * - TAG_TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - TAG_UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - TAG_FETCH_MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory, in 
   * -                      reads the allocation tags will be fetched from memory for read transactions.
   * .
   */
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0]{
    TAG_INVALID  = 0,
    TAG_TRANSFER = 1,
    TAG_UPDATE   = 2,
    TAG_FETCH_MATCH = 3
  } tag_op_enum;


 
/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   *  This field will be populated by the VIP and must not be set by the users.
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
 
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0] {
     MATCH_NOT_PERFORMED = 0,
     NO_MATCH_RESULT  = 1,
     FAIL = 2,
     PASS = 3
  } tag_match_resp_enum;  

`endif
 /**
   * Enum to represent four levels of shareability domain for snoop
   * transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE. 
   */
  typedef enum bit [1:0] {
    NONSHAREABLE      = `SVT_AXI_DOMAIN_TYPE_NONSHAREABLE,
    INNERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_INNERSHAREABLE,
    OUTERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_OUTERSHAREABLE,
    SYSTEMSHAREABLE   = `SVT_AXI_DOMAIN_TYPE_SYSTEMSHAREABLE
  } xact_shareability_domain_enum;

  /**
   * Enum to represent barrier transaction type. Enum to represent four levels
   * of shareability domain for snoop transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum bit [1:0] {
    NORMAL_ACCESS_RESPECT_BARRIER = `SVT_AXI_NORMAL_ACCESS_RESPECT_BARRIER,
    MEMORY_BARRIER                = `SVT_AXI_MEMORY_BARRIER,
    NORMAL_ACCESS_IGNORE_BARRIER  = `SVT_AXI_NORMAL_ACCESS_IGNORE_BARRIER,
    SYNC_BARRIER                  = `SVT_AXI_SYNC_BARRIER
  } barrier_type_enum;

  /**
   * Enum to represent responses for a coherent transaction Additional read
   * response bits that provide information on the completion of a shareable
   * read transaction.  Enum to represent barrier transaction type. Enum to
   * represent four levels of shareability domain for snoop transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */
  typedef enum  bit [1:0] {
    UNIQUE_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_CLEAN, 
    UNIQUE_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_DIRTY,
    SHARED_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_CLEAN,
    SHARED_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_DIRTY
  } coherent_resp_type_enum;

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [1:0] {
    NORMAL     = `SVT_AXI_TRANSACTION_NORMAL,
    EXCLUSIVE  = `SVT_AXI_TRANSACTION_EXCLUSIVE,
    LOCKED     = `SVT_AXI_TRANSACTION_LOCKED
  } atomic_type_enum;

  /**
   * Enum to represent the status of coherent exclusive access
   */
  typedef enum {
    EXCL_ACCESS_INITIAL  = `SVT_AXI_COHERENT_EXCL_ACCESS_INITIAL,
    EXCL_ACCESS_PASS     = `SVT_AXI_COHERENT_EXCL_ACCESS_PASS,
    EXCL_ACCESS_FAIL     = `SVT_AXI_COHERENT_EXCL_ACCESS_FAIL 
  } excl_access_status_enum;

  /** 
   * Enum to represent the status of master exclusive monitor, which indicates the cause of failure for a coherent exclusive store
   */ 
  typedef enum {
    EXCL_MON_INVALID  = `SVT_AXI_EXCL_MON_INVALID,
    EXCL_MON_SET      = `SVT_AXI_EXCL_MON_SET,
    EXCL_MON_RESET    = `SVT_AXI_EXCL_MON_RESET
  } excl_mon_status_enum;  

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [2:0] {
    DATA_SECURE_NORMAL                = `SVT_AXI_DATA_SECURE_NORMAL,               
    DATA_SECURE_PRIVILEGED            = `SVT_AXI_DATA_SECURE_PRIVILEGED,               
    DATA_NON_SECURE_NORMAL            = `SVT_AXI_DATA_NON_SECURE_NORMAL,               
    DATA_NON_SECURE_PRIVILEGED        = `SVT_AXI_DATA_NON_SECURE_PRIVILEGED,           
    INSTRUCTION_SECURE_NORMAL         = `SVT_AXI_INSTRUCTION_SECURE_NORMAL,            
    INSTRUCTION_SECURE_PRIVILEGED     = `SVT_AXI_INSTRUCTION_SECURE_PRIVILEGED,         
    INSTRUCTION_NON_SECURE_NORMAL     = `SVT_AXI_INSTRUCTION_NON_SECURE_NORMAL,        
    INSTRUCTION_NON_SECURE_PRIVILEGED = `SVT_AXI_INSTRUCTION_NON_SECURE_PRIVILEGED    
  } prot_type_enum;

  /**
   * Enum to represent responses in a transaction
   */
  typedef enum bit [1:0] {
    OKAY    = `SVT_AXI_OKAY_RESPONSE,
    EXOKAY  = `SVT_AXI_EXOKAY_RESPONSE,
    SLVERR = `SVT_AXI_SLVERR_RESPONSE,
    DECERR  = `SVT_AXI_DECERR_RESPONSE
  } resp_type_enum;

  typedef enum bit [2:0] {
    INVALID = `SVT_AXI_CACHE_LINE_STATE_INVALID,
    UNIQUECLEAN = `SVT_AXI_CACHE_LINE_STATE_UNIQUECLEAN,
    SHAREDCLEAN = `SVT_AXI_CACHE_LINE_STATE_SHAREDCLEAN,
    UNIQUEDIRTY = `SVT_AXI_CACHE_LINE_STATE_UNIQUEDIRTY,
    SHAREDDIRTY = `SVT_AXI_CACHE_LINE_STATE_SHAREDDIRTY
  } cache_line_state_enum;
 
  /**
   * Enum to represent DVM Message type.
   *
   * The bit representation of this type matches the encoding of the DVM message type field
   * in the AxADDR AMBA4 signal.
   * 
   * Used in the svt_amba_pv_extension class.
   */
  typedef enum bit [2:0] {
    TLB_INVALIDATE                        = 'h0, /**< TLB invalidate */
    BRANCH_PREDICTOR_INVALIDATE           = 'h1, /**< Branch predictor invalidate */
    PHYSICAL_INSTRUCTION_CACHE_INVALIDATE = 'h2, /**< Physical instruction cache invalidate */
    VIRTUAL_INSTRUCTION_CACHE_INVALIDATE  = 'h3, /**< Virtual instruction cache invalidate */
    SYNC                                  = 'h4, /**< Synchronisation message */
    HINT                                  = 'h6  /**< Reserved message type for future Hint messages */
  } dvm_message_enum;

  /**
   * Enum to represent DVM message Guest OS or hypervisor type.
   *
   * The bit representation of this type matches the encoding of the DVM guest OS or 
   * hypervisor field in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    HYPERVISOR_OR_GUEST = 'h0, /**< Transaction applies to hypervisor and all Guest OS*/
    GUEST               = 'h2, /**< Transaction applies to Guest OS */
    HYPERVISOR          = 'h3  /**< Transaction applies to hypervisor */
  } dvm_os_enum;

  /**
   * Enum to represent DVM message security type.
   *
   * The bit representation of this type matches the encoding of the DVM security field
   * in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    AMBA_PV_SECURE_AND_NON_SECURE = 'h0, /**< Transaction applies to Secure and Non-secure */
    AMBA_PV_SECURE_ONLY           = 'h2, /**< Transaction applies to Secure only */
    AMBA_PV_NON_SECURE_ONLY       = 'h3  /**< Transaction applies to Non-secure only */
  } dvm_security_enum;


  /**
   *  Enum for interleave block pattern
   */

  typedef enum {
    EQUAL_BLOCK   = `SVT_AXI_TRANSACTION_INTERLEAVE_EQUAL_BLOCK,
    RANDOM_BLOCK  = `SVT_AXI_TRANASCTION_INTERLEAVE_RANDOM_BLOCK
  } interleave_pattern_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    PREV_ADDR_VALID      =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_VALID_REF,
    PREV_ADDR_HANDSHAKE  =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_HANDSHAKE_REF,
    FIRST_WVALID_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_WVALID_DATA_BEFORE_ADDR,
    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR,
    PREV_LAST_DATA_HANDSHAKE = `SVT_AXI_MASTER_TRANSACTION_PREV_LAST_DATA_HANDSHAKE
  } reference_event_for_addr_valid_delay_enum;

  /** 
   *  Enum to represent data delay reference event
   */
  typedef enum {
    WRITE_ADDR_VALID                           = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_VALID_REF,    
    //removed address handshake refrence because  of potential deadlock due to following reason::
    //the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    WRITE_ADDR_HANDSHAKE                       = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_HANDSHAKE_REF,
    PREV_WRITE_DATA_HANDSHAKE                  = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_DATA_HANDSHAKE_REF
  }  reference_event_for_first_wvalid_delay_enum;

  typedef enum {
    PREV_WVALID            = `SVT_AXI_MASTER_TRANSACTION_PREV_WVALID_REF,
    PREV_WRITE_HANDSHAKE   = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_HANDSHAKE_REF
  } reference_event_for_next_wvalid_delay_enum;
  
  /** 
   *  Enum to represent tvalid delay reference event
   */
  typedef enum {
    PREV_TVALID_TREADY_HANDSHAKE          = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_TREADY_HANDSHAKE_REF,
    PREV_TVALID                           = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_REF
  }  reference_event_for_tvalid_delay_enum;

  typedef enum {
    RVALID               = `SVT_AXI_MASTER_TRANSACTION_RVALID_REF,                                 
    MANUAL_RREADY        = `SVT_AXI_MASTER_TRANSACTION_MANUAL_RREADY_REF       
  } reference_event_for_rready_delay_enum;

  /** 
   *  Enum to represent response delay reference event
   */
  typedef enum {
    BVALID               =   `SVT_AXI_MASTER_TRANSACTION_BVALID_REF
  } reference_event_for_bready_delay_enum;
 
  /** 
   * Enum to represent read acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    LAST_READ_DATA_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_LAST_READ_DATA_HANDSHAKE_REF
  } reference_event_for_rack_delay_enum;
  
  /** 
   * Enum to represent write acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    WRITE_RESP_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_WRITE_RESP_HANDSHAKE_REF
  } reference_event_for_wack_delay_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_ADDR_VALID_REF,
    FIRST_WVALID            = `SVT_AXI_SLAVE_TRANSACTION_FIRST_WVALID_REF
  } reference_event_for_addr_ready_delay_enum;

  /** 
   *  Enum to represent reference event for delay for first rvalid
   */
  typedef enum {
    READ_ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_VALID_REF,    
    READ_ADDR_HANDSHAKE           = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_HANDSHAKE_REF
  }  reference_event_for_first_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for second rvalid onwards
   */
  typedef enum {
    PREV_RVALID          = `SVT_AXI_SLAVE_TRANSACTION_PREV_RVALID_REF,
    PREV_READ_HANDSHAKE  = `SVT_AXI_SLAVE_TRANSACTION_PREV_READ_HANDSHAKE_REF
  } reference_event_for_next_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for wready signal
   */
  typedef enum {
    WVALID               = `SVT_AXI_SLAVE_TRANSACTION_WVALID_REF,                                 
    MANUAL_WREADY        = `SVT_AXI_SLAVE_TRANSACTION_MANUAL_WREADY_REF       
  } reference_event_for_wready_delay_enum;

  /** 
   *  Enum to represent write response delay reference event
   */
  typedef enum {
    LAST_DATA_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_LAST_DATA_HANDSHAKE_REF,
    ADDR_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_ADDR_HANDSHAKE_REF
  } reference_event_for_bvalid_delay_enum;

 
    
   // ****************************************************************************
   // Public Data
   // ****************************************************************************
   /** @groupname axi_misc
     * Variable that holds the object_id of this transaction
     */
   int object_id = -1;
   /** @groupname axi_misc
    * Variables used in generating XML/FSDB for pa writer 
    */
   
   string pa_object_type = "";
   string pa_channel_name ="" ;
   string bus_parent_uid = "";
   string bus_activity_type_name;

   /** @groupname axi_misc
     * The port configuration corresponding to this transaction
     */
   svt_axi_port_configuration port_cfg;
   
   /** 
    * @groupname ace_protocol
    * This member points to a barrier pair transaction
    * associated to this current transaction.  When associated_barrier_xact is
    * null, it indicates that this current transaction is not a post-barrier
    * transaction.  When associated_barrier_xact is non-null, this current
    * transaction will wait for responses from the barrier transactions in
    * associated_barrier_xact, before it can be transmitted.
    *
    * associated_barrier_xact can be set in the callback
    * svt_axi_master_callback::associate_xact_to_barrier_pair. In this
    * callback, user can associate this transaction with a barrier transaction
    * pair.
    *
    * Please refer to User Guide for more details on usage of this member.
    */
   svt_axi_barrier_pair_transaction  associated_barrier_xact;

`ifdef SVT_UVM_TECHNOLOGY
   /**
     * @groupname axi_misc 
     * Applicable only for master in ACTIVE mode.
     * If this transaction was generated from a UVM TLM Generic Payload, this
     * member indicates the GP from which this AXI transaction was generated
     */
   uvm_tlm_generic_payload causal_gp_xact;
`endif

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
    * Object used to hold exceptions for a packet. 
    */
  `ifndef __SVDOC__
  svt_axi_transaction_exception_list exception_list = null; 
  `endif
 /** W riter used in callbacks to generate output for pa or verdi */ 
  protected svt_xml_writer xml_writer = null ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_mask ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_range;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  burst_addr_mask ;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */

  //protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /**
    * Used in system monitor to indicate if all bytes of a slave transaction
    * has been correlated to a corresponding master transaction
    */
  bit  is_slave_xact_correlated = 0;
  
  /**
    * Used in port monitor to indicate resize and aligned data status
    * in data_before_addr transaction.
    */
  bit  is_resize_and_align_data = 0;


  /** 
    * Indicates if data read from memory for a given beat contains X
    * The slave driver uses this information to decide whether to 
    * drive X on data.
    */
  bit read_data_contains_x[];

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  // protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /** @endcond */

  /**
   * @groupname axi3_protocol
   * The variable holds the value of  AWID/WID/BID/ARID/RID signals.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ID_WIDTH. Default value of this macro is 8. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ID_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::id_width.
   */
  rand bit [`SVT_AXI_MAX_ID_WIDTH - 1:0] id = 0;

  /**
   * @groupname axi3_protocol
   * The variable represents AWADDR when xact_type is WRITE and  ARADDR when
   * xact_type is READ.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ADDR_WIDTH. Default value of this macro is 64. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ADDR_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::addr_width.
   */
  rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] addr = 0;
  
  /**
   * @groupname axi3_protocol
   * Represents the minimum byte address of this transaction. 
   * If tagging is enabled, this will be the minimum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the maximum byte address of this transaction. 
   * If tagging is enabled, this will be the maximum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the total byte count of this transaction. 
   *  .
   */
  rand int total_byte_count = 0;
  
  /**
   *  @groupname axi3_protocol
   *  The variable represents the actual length of the burst. For eg.
   *  burst_length = 1 means a burst of length 1.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI3, burst length
   *  of 1 to 16 is supported.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI4, burst length
   *  of 1 to 256 is supported.
   */ 
  rand bit [`SVT_AXI_MAX_BURST_LENGTH_WIDTH: 0] burst_length = 1;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst size of a transaction . The variable holds the value
   *  for AWSIZE/ARSIZE. 
   */
  rand burst_size_enum burst_size = BURST_SIZE_8BIT;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst type of a transaction. The burst type holds the value
   *  for AWBURST/ARBURST. Following are the possible burst types: 
   *  - FIXED
   *  - INCR
   *  - WRAP
   *  .
   */
  rand burst_type_enum burst_type = INCR;

  /**
   * @groupname axi3_protocol
   * Represents the transaction type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * - COHERENT : Represents a COHERENT transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE and
   * COHERENT transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI_ACE.
   */
  rand xact_type_enum xact_type = WRITE;
  
  /**
   * @groupname axi3_protocol
   * Represents the phase type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE 
   */
  phase_type_enum phase_type = WR_ADDR;

  /**
   * @groupname axi3_protocol
   * Represents the atomic access of a transaction.  The variable holds the
   * value for AWLOCK/ARLOCK. Following are the possible atomic types:
   * - NORMAL     
   * - EXCLUSIVE  
   * - LOCKED
   * .
   * Please note that atomic type LOCKED is not yet supported.
   */
  rand atomic_type_enum atomic_type = NORMAL;

`ifdef SVT_ACE5_ENABLE
  /**
   * Indicates the endianness of the Outbound Write Data in an Atomic transaction.
   */
  rand endian_enum endian = LITTLE_ENDIAN;
`endif

`ifdef SVT_ACE5_ENABLE
  /**
   * @groupname axi5_protocol
   * Represents the Unique ID indicator Feature.
   * The variable holds the value of AWIDUNQ/BIDUNQ/ARIDUNQ/RIDUNQ signals.<br>
   * The Variable is used to indicate that there are
   * no outstanding transactions going on with the same AWID/BID/ARID/RID respectively
   * and it will remain unique till the transaction is completed.
   * In order to use this feature, user need to pass the user defined macro
   * at compile time +define+SVT_ACE5_ENABLE.
   * Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_ACE5_ENABLE macro is only used to enable this feature and signals.
   * The Signals can be configured and enabled by VIP configuration using
   * parameter svt_axi_port_configuration::unique_id_enable.
   *
   * This functionality is not supported yet.
   */
  rand bit unique_id = 0;
`endif

  /**
   *  @groupname axi3_protocol
   *  Represents the cache support of a transaction. The variable holds the
   *  value for AWCACHE/ARCACHE.
   *
   *  Following values are supported in AXI3 mode:
   *
   *  - SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE            
   *  - SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY           
   *  - SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC                  
   *  - SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_BOTH_RD_WR    
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_BOTH_RD_WR    
   *  .
   *  
   *  Following values for ARCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE      
   *  .
   *
   *  Following values for AWCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_AWCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_AWCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE    
   *  .
   */

  rand bit [`SVT_AXI_CACHE_WIDTH - 1:0] cache_type = 0;

  /**
   *  @groupname axi3_protocol
   *  Represents the protection support of a transaction. The variable holds the
   *  value for AWPROT/ARPROT. The conventions of the enumeration are:
   *
   *  - NORMAL/PRIVILEGED   : Normal/Priveleged access represented by AWPROT[0]/ARPROT[0]
   *  - SECURE / NON_SECURE : Secure/Non-Secure access represented by AWPROT[1]/ARPROT[1]
   *  - DATA / INSTRUCTION  : Data/Instruction access represented by AWPROT[2]/ARPROT[2]
   *  .
   *
   *  For the above conventions, following are the possible protection types:
   *  - DATA_SECURE_NORMAL                    
   *  - DATA_SECURE_PRIVILEGED                    
   *  - DATA_NON_SECURE_NORMAL                    
   *  - DATA_NON_SECURE_PRIVILEGED                
   *  - INSTRUCTION_SECURE_NORMAL                 
   *  - INSTRUCTION_SECURE_PRIVILEGED              
   *  - INSTRUCTION_NON_SECURE_NORMAL
   *  - INSTRUCTION_NON_SECURE_PRIVILEGED
   *  .
   */

  rand  prot_type_enum prot_type = DATA_SECURE_NORMAL;

  /**
   *  @groupname ace_protocol
   *  Applicable when
   *  svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.  
   *  Users  who need to bypass lookup of cache to determine valid 
   *  initial cache line states can set this property to 1.
   *  In order to randomize this property to 1, the user must switch off 
   *  svt_axi_master_transaction::reasonable_bypass_cache_lookup constraint.
   *  Setting this property will enable transactions to be sent out even
   *  if the initial cache state does not meet requirements set by ACE 
   *  protocol. Please note that coherency is not guaranteed when this 
   *  property is set
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand  bit bypass_cache_lookup = 1'b0;  


  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`endif

`ifdef SVT_ACE5_ENABLE

 /**
   * @groupname ace5_protocol
   * This variable represents the read data for the atomic load,swap and compare transactions.
   * This data will be driven by the slave on the read data channel.
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the Memory Tag value in the transaction driven on the data channel for transactions.
  * Every 4 bits of Tag correspond to one 16 byte chunk of data.
  * MASTER in active mode:
  *
  * For write transactions this variable specifies tags to be driven on the
  * WTAG bus. 
  * 
  * SLAVE in active mode:
  *
  * For read transactions this variable specifies tags to be driven on the
  * RTAG bus.
  *
  * PASSIVE MODE:
  * This variable stores the tags as seen on WTAG or RTAG bus.
  *
  *
  */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`else
  rand bit [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the WTAGUPDATE value in the transaction.
  * Only applicable when the Tag value is passed in the transaction and the tagop field in 
  * the transaction is set to Update.
  * Each WTAGUPDATE bit corresponds to 4 bits of WTAG
  */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`else
  rand bit [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`endif

/**
  * @groupname ace5_protocol
  * This field defines the BCOMP value in the transaction.
  * Indicates whether write transaction is observable at the completer endused for persistent CMOs on Write channel.
  * This is used to send the response to a tag Match operation.
  * This is also used for persistent CMOs on Write channel.
  */
 
 rand bit is_write_transaction_observable = 0;
//---------------------------------------------------------------------------------------------
 
 /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DATA channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
  rand tag_op_enum tag_op = TAG_INVALID ;

  /** 
   * Enum to represent the response sent by the completer on the corresponding Response channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
 rand tag_op_enum response_tag_op = TAG_INVALID;
 
//---------------------------------------------------------------------------------------------

/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
   rand tag_match_resp_enum tag_match_resp = MATCH_NOT_PERFORMED ;

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This field defines the partition ID value in MPAM. This corresponds to AxMPAM[9:1] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PARTID_WIDTH - 1:0] mpam_partid;

 /**
   * @groupname ace5_protocol
   * This field defines the Perfromance Monitor Group (PMG) value in MPAM. This corresponds to AxMPAM[10] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PERFMONGROUP_WIDTH - 1:0] mpam_perfmongroup;

 /**
   * @groupname ace5_protocol
   * This field defines the MPAM_NS value in MPAM. This corresponds to AxMPAM[0] attribute.
   */
  rand bit [`SVT_AXI_MPAM_NS_WIDTH - 1:0] mpam_ns;
//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the data that will be stored in the memory for atomic transactions 
   * after the atomic operation is performed.
   * APPLICABLE IN ALL MODES:
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`else
  bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`endif


//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the swap data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   * 
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`endif

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`endif

`endif

  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`endif

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable is only applicable for atomic transactions.
   * MASTER in active mode:
   * For Atomic LOAD , SWAP and COMPARE transactions specifies read data as seen on the RDATA bus. 
   * 
   * SLAVE in active mode:
   * This variable represents the read data for the atomic load,swap and compare transactions to be driven on the RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the read data as seen on RDATA bus.
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`endif

`endif

  /** @cond PRIVATE */
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string data_str = "";

`ifdef SVT_ACE5_ENABLE
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string atomic_read_data_str = "";
`endif

  /**
    * The wstrb array in string format. Used by psdisplay_short
    */
  local string wstrb_str = "";

  /**
    * The read response array in string format. Used by psdisplay_short
    */
  local string rresp_str = "";

  /**
    * The write response in string format. Used by psdisplay_short
    */
  local string bresp_str = "";

  /**
    * The valid_assertion_time in string format. Used by psdisplay_short
    */
  local string valid_assertion_time = "";
  
  /**
    * The ready_assertion_time in string format. Used by psdisplay_short
    */
  local string ready_assertion_time = "";
  
 /* holds transactions that attempt to access same cacheline at the same time current transaction

   * does and started before current transaction started */
  bit overlapped_xact_started_before[svt_axi_transaction];

  /* holds transactions that attempt to access same cacheline at the same time current transaction
   * does and started after current transaction started */
  bit overlapped_xact_started_after[svt_axi_transaction];
  
  /* Indicates xact complets with out_of_order*/
  bit is_xact_completed_out_of_order = 0;

  /* indicates how many transactions blocked progress of current transaction */
  int num_xacts_blocked_progress_of_curr_xact = 0;

  /* semaphore to access num_xacts_blocked_progress_of_curr_xact */
  semaphore sema_num_xacts_blocked_progress_of_curr_xact = new(1);
  /** @endcond */

  
  /**
   *  @groupname axi3_protocol
   *  Array of Write strobes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  wstrb must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the wstrb is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] wstrb[];

`ifdef SVT_ACE5_ENABLE
 
//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the swap write strobes  value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   * 
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_swap_wstrb[];

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare write strobes value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   */
   rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_compare_wstrb[];

`endif

  /**
   *  @groupname ace5_protocol
   *  Array of poison.It indicates the 
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] poison[];

`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname ace5_protocol
   *  Array of poisonal value driven by the active slave on the read data channel.
   *  This is onlyapplicable for Atomic LOad , Swap and compare transactions.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] atomic_read_poison[];

`endif


  /**
   *  @groupname axi3_protocol
   *  This variable specifies the response for write transaction. The variable holds the
   *  value for BRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the write response received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The write response programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the write response seen on the bus.
   */

  rand resp_type_enum bresp = OKAY;

  /**
   *  @groupname axi3_protocol
   *  This array variable specifies the response for read transaction. The array holds the
   *  value for RRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the read responses received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The read responses programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the read responses seen on the bus.
   */

  rand resp_type_enum rresp[];

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE 
  /** 
    * @groupname axi3_protocol
    * If set, the driver checks if this transaction accesses a location
    * addressed by a previous transaction from this port or from some other
    * master. If there are any such previous transactions, this transaction is
    * blocked until all those transactions complete.  Also, the driver does not
    * pull any more transactions until this transaction is unblocked.  If not set,
    * this transaction is not checked for access to a location which was
    * previously accessed by another transaction.  Applicable only when
    * svt_axi_system_configuration::overlap_addr_access_control_enable is set 
    *
    * Applicable for ACTIVE MASTER only
    */ 
  rand bit check_addr_overlap = 1'b0;

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * Suspends a master transaction until this bit is reset. This is checked
    * immediately after a transaction is pulled by the driver from the sequencer
    * after the post_input_port_get callback is issued by the driver. When set,
    * the driver does not pull any more transactions from the
    * sequencer/generator until the bit is reset
    *
    * Applicable for ACTIVE MASTER only
    */
  bit suspend_master_xact = 1'b0;
  /** @endcond */
   
`endif

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * This bit is set by master if a cache line is reserved for the transaction. 
    * Thie field is used by task which unreserves the cache line at the end of 
    * transaction to filtering. This is to ensure only command that reserved 
    * cache line should unreserve cache line.  
    *  
    * Applicable for ACTIVE MASTER only
    */
  bit is_cacheline_reserved = 1'b0;
  /** @endcond */

  /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend response/data
    * for a READ/WRITE/COHERENT transaction until this bit is reset. 
    * This bit is usually set by the testbench when it needs to provide
    * response information to the driver (the slave driver expects the response
    * information in 0 time), but the data to respond with is
    * not yet known.  The testbench can set this bit and put this transaction 
    * back into the input channel of the slave. 
    * The transaction's response/data will not be sent until this bit is reset. 
    * Once the data is available, the testbench can populate response fields 
    * and reset this bit, upon which the slave driver will send the 
    * response/data of this transaction.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_response = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend awready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_awready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_awready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend arready signal 
    * for a READ transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_arready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_arready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend wready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_wready is set to 0
    * svt_axi_transaction::wready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_wready = 0;

  /**
    * @groupname ace_protocol
    * Represents the value of AWUNIQUE signal driven/sampled on the interface.
    * Applicable when svt_axi_port_configuration::awunique_enable is set.
    * AWUNIQUE is asserted as per table C3-9 of section C3.1.4 on AWUNIQUE
    * signal. The value in the randomized transaction may be overridden by the
    * driver as per protocol requirements. For transactions where AWUNIQUE may
    * be asserted or deasserted, the randomized value is driven.  
    */
  rand bit is_unique = 0;

  /**
   *  @groupname axi3_4_status
   *  Represents the current status of the read or write address.  Following are the
   *  possible status types.

   * - INITIAL               : Address phase has not yet started on the channel
   * - ACTIVE                : Address valid is asserted but ready is not 
   * - ACCEPT                : Address phase is complete 
   * - ABORTED               : Current transaction is aborted
   * .
   */

  status_enum addr_status = INITIAL;

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum data_status = INITIAL;

`ifdef SVT_ACE5_ENABLE
/**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum atomic_read_data_status = INITIAL;
`endif

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the write response transfer.  Following are
   *  the possible status types.
   *  - INITIAL               : Response has not yet started on the channel
   *  - ACTIVE                : BVALID is asserted, but not BREADY
   *  - ACCEPT                : Write response is complete
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */


  status_enum write_resp_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of the read/write acknowledge sent via RACK/WACK for
   * ACE interface. RACK/WACK is asserted for a single cycle.
   * Following are  the possible status types:
   * - INITIAL               : RACK/WACK has not be asserted
   * - ACTIVE                : RACK/WACK is asserted
   * - ACCEPT                : RACK/WACK assertion is completed
   * - ABORTED               : Current transaction is aborted
   * .
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */

  status_enum ack_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of coherent exclusive access.
   * Following are  the possible status types: 
   * - EXCL_ACCESS_INITIAL   : Initial state of the transaction before it is processed by master 
   * - EXCL_ACCESS_PASS      : ACE exclusive access is successful
   * - EXCL_ACCESS_FAIL      : ACE exclusive access is failed
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description. 
   */
  excl_access_status_enum  excl_access_status = EXCL_ACCESS_INITIAL;
  

  /**
   * @groupname ace_status
   * Represents the status of master exclusive monitor, which indicates the
   * cause of failure for a coherent exclusive store.  It is valid only for
   * exclusive store transaction, that is, CleanUnique. For all other
   * transactions it is set to EXCL_MON_INVALID by default.
   * Following are  the possible status types:
   * - EXCL_MON_INVALID      : Master exclusive monitor does not monitor the exclusive access on the cache line associated with the transaction
   * - EXCL_MON_SET          : Master exclusive monitor is set for exclusive access on the cache line associated with the transaction
   * - EXCL_MON_RESET        : Master exclusive monitor is reset for exclusive access on the cache line associated with the transaction
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description.
   */ 
  excl_mon_status_enum   excl_mon_status = EXCL_MON_INVALID;


  /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  current_data_beat_num = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  atomic_read_current_data_beat_num = 0;
`endif
  /**
   *  @groupname interleaving
   *  Represents the various interleave pattern for a read and write transaction.
   *  The interleave_pattern gives flexibility to program interleave blocks with
   *  different patterns as mentioned below.
   *
   *  A Block is group of beats within a transaction.
   *
   *  EQUAL_BLOCK         : Drives equal distribution of blocks provided by
   *                        #equal_block_length variable. 
   *
   *  RANDOM_BLOCK        : Drives the blocks programmed in random_interleave_array
   *
   * Please note that currently interleaving based on EQUAL_BLOCK is not
   * supported.
   */
  rand interleave_pattern_enum interleave_pattern = RANDOM_BLOCK;

  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  If the interleave_pattern is set to EQUAL_BLOCK then this variable 
   *  is used to define the block length.
   *  Please note that currently interleaving based on EQUAL_BLOCK is not
   *  supported.
   */

  rand int equal_block_length = 0;

  /** @endcond */

  /**
   *  @groupname interleaving
   *  When the interleave_pattern is set to RANDOM_BLOCK, the user would
   *  program this array with blocks. There are default constraints, which the
   *  user can override and set their own block patterns.
   */
  rand int random_interleave_array[];


  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  This variable will start a new interleave from the current transaction and
   *  informs the model to complete all the transactions prior to this
   *  transaction.
   *
   *  Example 1:
   *  Interleave depth = 2
   * 
   *  Requirement : 
   *  1) Interleave transaction 1- 10 with each other
   *  2) Interleave transactions 11 - 20 with each other
   *
   *  Solution :
   *  1) Program start_new_interleave=0 for transactions 1 - 10 
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Example 2:
   *  Interleave depth = 2
   *
   *  Requirement :
   *  1) Do not Interleave transactions 1 - 10
   *  2) Start Interleaving from transactions 11 - 20
   *
   *  Solution :
   *  1) Program start_new_interleave=1 for transactions 1-10
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Please note that this parameter is not currently supported.
   */
  rand bit start_new_interleave = 0;
  /** @endcond */

  /**
   * @groupname interleaving , out_of_order
   * This variable controls enabling of interleaving for the current transaction.
   * 
   * Example:
   * svt_axi_port_configuration::read_data_reordering_depth = 2
   * 
   * Requirement:
   * Unless all beats of transaction 1 are sent out, the beats of 
   * 2nd transactions should not be sent.
   * 
   * Solution:
   * Program the enable_interleave = 0 for both the transaction 1.
   
   */
  rand bit enable_interleave = 0;
  
  /**
    * @groupname axi_protocol
    * When this bit is set , it indicates that this transaction has updated 
    * the AXI Slave memory with write data and other properties.
    */ 
  bit memory_update_complete_for_write =0;

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * when this bit is set, it indicates that this transaction 
   * performed atomic operation and the result is stored in atomic_resultant_data.
   */
  bit is_atomic_resultant_data_calculated =0;
`endif 

  /**
   * @groupname ace_protocol
   * When this bit is set by user, it indicates that this transaction is
   * a post-barrier transaction and that it needs to wait for responses
   * from the barrier transaction pair indicated in #associated_barrier_xact.
   * #associated_barrier_xact can be set in the callback
   * svt_axi_master_callback::associate_xact_to_barrier_pair. In this callback,
   * user can associate this transaction with a barrier transaction pair.
   *
   * Please refer to User Guide for more description.
   */
  rand bit associate_barrier = 0;

  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions.
   *  In data_before_addr scenario (i.e., when data_before_addr = '1'), addr and data channel related delay considerations are: 
   *  1) For programming address_channel related delay: awvalid_delay and reference_event_for_addr_valid_delay are used.
   *   (for more information, look for the description of these variables).
   *    reference_event_for_addr_valid_delay should be set FIRST_WVALID_DATA_BEFORE_ADDR. 
   *    In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
   *    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
   *    potential deadlock scenarios in SLAVE DUT where slave DUT waits for awvalid signal
   *    before driving wready signal.
   *  2) For programming data_channel related delay: wvalid_delay[] and reference_event_for_first_wvalid_delay & reference_event_for_next_wvalid_delay are used.
   *    (for more information, look for the description of these variables).
   *      For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
   *      For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
   *    In data_before_addr scenario, reference_event_for_first_wvalid_delay must be PREV_WRITE_DATA_HANDSHAKE, otherwise it will cause failure.
   *  .
   *    
   */
  rand bit data_before_addr = 0;
  
  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions,
   *  even though data_before_addr is set to 0. This is useful when
   *  awvalid is suspended for write transaction and respective transaction
   *  data is driven before resuming the suspended awvalid signal.
   */
  bit suspend_awvalid_to_data_before_addr = 0;

  /**
    * Indicates if the current data beat of a write transaction has wlast
    * asserted. This is useful when data is received before addr and it is
    * required to determine the last beat. This is a sticky bit  in that
    * it remains set to 1 after the last data beat.
    */ 
  bit is_last_write_data_beat = 0;

   // AXI 4 Variables

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWQOS/ARQOS 
   */
  rand bit[`SVT_AXI_QOS_WIDTH - 1:0] qos = 0;  
  

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWREGION/ARREGION
   */
  rand bit[`SVT_AXI_REGION_WIDTH - 1:0] region = 0;


  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals AWUSER/ARUSER.
   *  Applicable for all interface types. Enabled through port configuration
   *  parameters svt_axi_port_configuration::aruser_enable and
   *  svt_axi_port_configuration::awuser_enable.
   */
  rand bit[`SVT_AXI_MAX_ADDR_USER_WIDTH - 1:0] addr_user = 0;

  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER. Applicable for all
   *  interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] data_user[];

`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname ace5_protocol
   *  The variable holds the value for signals RUSER.
   *  Applicable only if svt_axi_port_configuration::atomic_transactions_enable is set to1.
   *  Enabled through port configuration parameters
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] atomic_read_data_user[];
`endif

   /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER as they are driven on the bus
   *  Applicable for all interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
   bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] physical_data_user[];
 /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signal BUSER. Applicable for all
   *  interface types. Enabled through port configuration parameter
   *  svt_axi_port_configuration::buser_enable.
   */
  rand bit[`SVT_AXI_MAX_BRESP_USER_WIDTH - 1:0] resp_user = 0;
  
  /** 
   * @groupname ace_protocol
   * This variable represents the shareability domain of coherent transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE or ACE_LITE.
   */
  rand xact_shareability_domain_enum domain_type = NONSHAREABLE;

  /**
   * @groupname ace_protocol
   * This variable represents barrier transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand barrier_type_enum barrier_type = NORMAL_ACCESS_RESPECT_BARRIER;

  /** 
   * @groupname ace_protocol
   * This variable represents the shareable coherent transaction types. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand coherent_xact_type_enum coherent_xact_type = READNOSNOOP;

`ifdef SVT_ACE5_ENABLE
 /**
  * @groupname ace5_protocol 
  * This variable represents the cmo on the write channel.
  * Applicable when svt_axi_port_configuration::axi_interface_type is set to ACE_LITE.
  */
  rand cmo_on_write_xact_type_enum cmo_on_write_xact_type = CLEANSHARED_ON_WRITE;
`endif

  /** 
   * @groupname ace_protocol
   * Array for the coherent read responses. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  rand coherent_resp_type_enum coh_rresp[];

  /**
    * @groupname ace_status
    * This variable represents the initial cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The initial cache line state of a transaction that is driven on
    * the READ channel is populated just after the reception of the first beat
    * of the response of a transaction.  The initial cache line state of a
    * transaction that is driven on the WRITE channel is populated just before
    * the transaction is started. This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum initial_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the prefinal cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The prefinal cache line state of a transaction is the state of the 
    * cache  just before cache is updated . This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum  prefinal_cache_line_state = INVALID;

   /*
    * @groupname ace_status
    * This variable represents the initial data in the cache. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE. For transactions driven on the READ channel, this field is 
    * populated just after the reception of the the first beat of the response
    * of the transaction.
    * For transactions driven on the WRITE channel, this is populated just
    * before the transaction is started.
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] initial_cache_line_data[];

  /**
    * @groupname ace_status
    * This variable represents the final cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The final cache line state of a transaction is the state of the
    * the line just before the transaction ended. This variable is updated by
    * the VIP, and is a read-only variable. User is not expected or supposed to
    * modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum final_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the final cache line data. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * The final cache line data of a transaction is the data of the
    * the line just before the transaction ended. 
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] final_cache_line_data[];

  /**
   * @groupname ace_protocol
   * Indicates that the data as given in #cache_write_data in this transaction 
   * needs to be allocated in the cache. Applicable only when transaction type
   * is READUNIQUE or CLEANUNIQUE.
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Applicable for ACTIVE MASTER only.
   */
  rand bit allocate_in_cache;

  /**
   * @groupname ace_protocol
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Represents data that needs to be stored to the cache if the 
   * #allocate_in_cache bit is set for a READUNIQUE/CLEANUNIQUE transaction 
   * or if the transaction is MAKEUNIQUE.
   * Applicable to masters in active mode.
   * Refer section 3.6 of ACE specification.
   * Writes in ACE are performed by removing all other copies
   * of the cache line so that the master that is performing the write has
   * a unique copy at the time of writing. Depending on whether a paritial
   * or full update of a cache line is required a transaction such as
   * READUNIQUE,MAKEUNIQUE or CLEANUNIQUE is sent. Some of these transactions
   * such as READUNIQUE will return data (either from memory or the cache of
   * some other master) and this will be available in the data[] field of this
   * class. Other transactions such as MAKEUNIQUE and CLEANUNIQUE will not
   * return any data. 
   * For a READUNIQUE transaction, if the #allocate_in_cache bit is not set, the
   * data available in data[] is written in cache. If the #allocate_in_cache bit
   * is set the data available in this variable is written to cache. Note however,
   * that this variable is overwritten by the data that is received in data[] prior
   * to writing in the cache. This is done because READUNIQUE is used for partial update 
   * of a cacheline when a master does not have a copy of the cacheline. So a user 
   * can actually populate this variable after a copy of this cacheline is received and 
   * not at the time of randomization.
   * For a CLEANUNIQUE transaction, if the #allocate_in_cache bit is set,
   * the data in this variable is written to cache. 
   * For a MAKEUNIQUE transaction, the data in this variable is always written into
   * the cache.
   * Updating this variable is normally done in the pre_cache_update callback issued 
   * by the master driver after all the responses are received but prior to the 
   * RACK signal being driven.
   * An important aspect of this variable is that this data is not driven
   * on the physical bus.
   * 
   * Applicable for ACTIVE MASTER only.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] cache_write_data[];

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if update of cache must be bypassed for this transaction. A
    * typical use model is to set this bit in pre_cache_update callback of the
    * driver based on response received in the transaction. For example, if the
    * response received is SLVERR, user may not want the driver to update the
    * cache.  When using this property, it is the user's responsibility that
    * system coherency is not lost, since cache will not be updated.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit bypass_cache_update = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction ended because the requested data was already
    * available in the cache. This bit is set by the master, no action is taken
    * if the user sets this bit. A transaction with this bit set was not sent out
    * on the bus and therefore other components in the testbench will not detect
    * this transaction. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_cached_data = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if a coherent transaction was dropped because the start state
    * of the corresponding cache line is not as expected before transmitting the
    * transaction. The expected start states for each of the transaction types
    * are given in section 5 of the ACE specification.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_coherent_xact_dropped = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is a result of a speculative read operation.
    * A speculative read is defined as a read of a cache line that a master already
    * holds in its cache.
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is a speculative read. Modifying the value of this member will
    * not have any effect.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_speculative_read = 0;

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates whether the memory update at slave end for overlapped write
    * transactions should happen in request order.
    *
    * This is a read-only member, which VIP uses to update slave memory for 
    * overlapped write transactions. It should not be modified by the user.
    * 
    * Applicable for ACTIVE SLAVE only.
    */
  bit update_mem_in_req_order = 0;  

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for WriteUnique and WriteLineUnique
    * not being in progress while a WRITEBACK/WRITECLEAN is in progress is done
    * Applicable when port_interleaving_enable is set in the configuration.
    */
  bit is_wu_wlu_restriction_check_done = 0;

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for memory update transaction 
    * relative to the cache states are performed just prior to start
    * of this transaction
    */
  bit is_mem_update_pre_xact_xmit_check_done = 0;
  /** @endcond */

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is auto generated by the VIP. Transactions
    * are auto-generated when:
    * 1. The cache is full and an entry needs to be evicted from the cache. 
    * 2. User supplies a cache maintenance transaction and the protocol requires
    * that the cache line is first written into memory before sending the cache
    * maintenance transaction. 
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is auto generated. It should not be modified by the user. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_auto_generated = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set
    * to AXI_ACE and svt_axi_port_configuration::snoop_response_data_transfer_mode 
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC.
    *
    * Indicates if this transaction is a WRITEBACK/WRITECLEAN auto-generated transaction
    * which was generated to transfer snoop data. When 
    * svt_axi_port_configuration::snoop_response_data_transfer_mode is set to 
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, snoop data from a dirty line is transferred
    * using a WRITEBACK/WRITECLEAN transaction instead of the snoop data channel. All
    * transactions which have this variable set will also have  is_auto_generated set.
    */
  bit is_xact_for_snoop_data_transfer = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to a shared state even
    * if the actual state of the line is unique, since it is permissible for
    * a cache line which is in the unique state to be held in the shared state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE or
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_shared_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to an invalid state even
    * if that is not the recommended state, since it is permissible for
    * a cache line which is in a clean state to be held in the invalid state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_invalid_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set to
    * AXI_ACE or ACE_LITE.  Forces transactions which are not constrained to be
    * of cacheline size by protocol to be of cacheline size. Currently
    * applicable only to READONCE, WRITEUNIQUE, WRITENOSNOOP and READNOSNOOP
    * transactions. Applicable to WRITENOSNOOP and READNOSNOOP only when
    * svt_axi_port_configuration::update_cache_for_non_coherent_xacts is set and
    * svt_axi_port_configuration::axi_interface_type is AXI_ACE.
    * If this bit is set, READONCE and WRITEUNIQUE transactions will be forced
    * to cache line size transactions.
    * This has a dependency on svt_axi_port_configuration::force_xact_to_cache_line_size_interface_type. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_xact_to_cache_line_size = 0;
  
  /**
   * @groupname ace_protocol
   * The variable represents ARVMIDEXT when svt_axi_port_configuration::axi_interface_type 
   * is set to AXI_ACE or ACE_LITE with svt_axi_system_configuration::DVMV8_1 or above.
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_VMIDEXT_WIDTH. Default value of this macro is 4 based on DVMv8.1 architecture recomendation.
   * 
   */

  rand bit [`SVT_AXI_MAX_VMIDEXT_WIDTH - 1:0] arvmid = 0;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit is_datachk_parity_error = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit atomic_read_is_datachk_parity_error = 0;

  /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_transaction_type_enum atomic_transaction_type = NON_ATOMIC;

 /**
  * - @groupname ace5_protocol
  * - Field that indicates type of write_with_cmo_xact_type.
  * .
  */

  rand write_with_cmo_xact_type_enum write_with_cmo_xact_type = WRITENOSNPFULL_CLEANSHARED; 

 /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_xact_op_type_enum atomic_xact_op_type = ATOMICSTORE_ADD;

`endif
 /**
   * @groupname ace5_protocol 
   *This field indicates the value of trace_tag
   */
  rand bit trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of data trace_tag on write data channel and read data channel
   */
  rand bit data_trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of btrace on write response channel
   */
  rand bit resp_trace_tag =0;

`ifdef SVT_ACE5_ENABLE 
  /** Internal field to store the atomic data trace_tag for inbound data */
  rand bit atomic_read_data_trace_tag;

 /** 
   * @groupname ace5_protocol
   * This field indicates the node ID of the stash target. 
   * Applicable only in stash type transactions.
   */
  rand bit[(`SVT_AXI_STASH_NID_WIDTH-1):0] stash_nid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates the stash_nid field has a valid Stash target value.
   * Applicable only in stash type transactions.
   */
  rand bit stash_nid_valid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  indicates the ID of the logical processor at the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit [(`SVT_AXI_STASH_LPID_WIDTH-1):0] stash_lpid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the Stash_lpid field value must be 
   * considered as the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit stash_lpid_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates the ID of the stream.This si used to identify the stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit [(`SVT_AXI_MAX_MMUSID_WIDTH-1):0] stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates wether the stream is secure or non-secure.
   * When set to 1, indicates a secure stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit secure_or_non_secure_stream = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  is only vaid if sub_stream_id_valid is set to 1.
   * This indicates the ID of the sub stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit[(`SVT_AXI_MAX_MMUSSID_WIDTH-1):0] sub_stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has an optional substream identifier.
   * When set to 1 , it means that transaction has a substream identifier.
   * This is used in untranslated transaction feature is enabled.
   */
  rand bit sub_stream_id_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has already undergone PCIE ATS 
   * translation.
   */
  rand bit addr_translated_from_pcie = 0;

`endif

  /**
   *  Represents port ID. Not currently supported.
   */
  int port_id;

  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the cycle information for address valid on read and
   *   write transactions. The simulation clock cycle number when the address
   *   valid is asserted, is captured in this member. This information can be
   *   used for doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */
  int addr_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_valid_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_valid_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response valid on a write
   *  transaction. The simulation clock cycle number when the write response
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */
  int write_resp_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation clock cycle number when the address valid
   *  and ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */
  int addr_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_ready_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_ready_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response ready on a write
   *  transaction. The simulation clock cycle number when the write response valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int write_resp_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *   The simulation time when the master or slave driver receives
   *   the transaction from the sequencer, is captured in this member.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  realtime xact_consumed_by_driver_time;
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for address wakeup of read or write 
   *  transaction. The simulation clock cycle number when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  int addr_wakeup_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address wakeup of read or write
   *  transaction. The simulation time when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real addr_wakeup_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real idle_chan_wakeup_toggle_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  deasserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
   real idle_chan_wakeup_toggle_deassertion_time;

 /**
   *   @groupname axi3_4_ace_timing
   *   This variable stores the transaction consumed at driver timing
   *   information. The transaction consumed at driver time to begin time
   *   delay is calculated as the difference between begin_time and
   *   xact_consumed_by_driver_time.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member variable,
   *   user does not need to program this variable.
   */

  real xact_consumed_time_to_begin_time_delay;
  
  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the timing information for address valid on read and
   *   write transactions. The simulation time when the address valid is
   *   asserted, is captured in this member. This information can be used for
   *   doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  real addr_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_valid_assertion_time[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_valid_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response valid on  write
   *  transactions. The simulation time when the response valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real write_resp_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation time number when the address valid and
   *  ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */

  realtime addr_ready_assertion_time;


  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_ready_assertion_time[];
`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_ready_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response ready on  write
   *  transactions. The simulation time when the response valid and ready both are
   *  asserted, is captured in this member. This information can be used for doing
   *  performance analysis. VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */

  real write_resp_ready_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for the data channnel blocking ratio.
   *  The blocking cycle for a beat is defined as the number of cycles that
   *  valid was asserted, but corresponding ready was not asserted.
   *  This ratio is derived from data_valid_assertion_cycle and
   *  data_ready_assertion_cycle, calculated as sum of data ready
   *  blocking cycles divided by sum of data valid assertion cycles.
   *  This information can be used for doing performance analysis.
   *  VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */
  real data_chan_blocking_ratio;

  // ****************************************************************************
  // Members relevant to Master Driver and Monitor  
  // ****************************************************************************

  /**
    * @groupname axi3_4_delays
    * This variable defines the number of cycles the AWVALID or ARVALID  signal is
    * delayed. The reference event for this delay is #reference_event_for_addr_valid_delay.
    * Applicable for ACTIVE MASTER only.
    */
  rand int addr_valid_delay = 0;
   
  /**
    * @groupname axi3_4_delays
    * Defines a reference event from which the AWVALID or ARVALID delay
    * should start.  Following are the different reference events:
    *
    * PREV_ADDR_VALID:  
    * Reference event is the previous AWVALID or ARVALID signal 
    *
    * PREV_ADDR_HANDSHAKE:  
    * Reference event is previous read or write Address handshake
    *
    * FIRST_WVALID_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first wvalid of the current transaction.
    *
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first data handshake of the current transaction.
    *
    * PREV_LAST_DATA_HANDSHAKE:
    * Reference event is previous read or write last data handshake
    * to Address valid assertion.
    *
    * Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios is added in svt_axi_transaction class 
    * to constraint the value of reference_event_for_addr_delay not to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * User may swicth off the constraint reasonable_reference_event_for_addr_delay by setting rand_mode to 0 
    * incase they want reasonable_reference_event_for_addr_delay to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
    * potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
    * before driving wready signal.
    *
    */
  rand reference_event_for_addr_valid_delay_enum  reference_event_for_addr_valid_delay = PREV_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal assertion
    * before or after ARVALID or AWVALID signal.
    */
  rand int awakeup_assert_delay = 0;
  
  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal deassertion
    * after ARVALID-ARREADY or AWVALID-AWREADY signal handshake.
    */
  rand int awakeup_deassert_delay = 0;

  /** if this bit is set to '0' then AWAKEUP signal will be asserted 
    * before ARVALID with respect to awakeup_assert_delay.
    * if this bit is set to '1' then AWAKEUP signal will be asserted
    * after ARVALID or AWVALID with respect to awakeup_assert_delay.
    */ 
  rand bit assert_awakeup_after_valid = 0;

  /** 
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for WVALID signal.
    * The reference event for this delay is:
    * - For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
    * - For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
    * .
    * Applicable for ACTIVE MASTER only.
    */
  rand int wvalid_delay[];
   
  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * FALSE, this member defines the RREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_rready_delay
    *
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * TRUE, this member defines the number of clock cycles for which RREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int rready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which RREADY should be high and low
    * when the read data channel is idle, that is, when RVALID is low. This
    * property helps to toggle the RREADY signal during the idle period between
    * the assertion of RVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all read data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the read_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transaction unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until RVALID is asserted. When RVALID is observed on the interface,
    * this delay is no longer applicable. The delay specified in
    * #rready_delay is applied before this property is used.  Note that toggling
    * RREADY during the idle period may lead to situations where the RREADY
    * signal is already asserted when the RVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_rready is low. Similarly,
    * RREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_rready is high. In both
    * these cases, #rready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_rready_delay[];

  /**
   * @groupname axi4_stream_delays
   * Defines the delay in number of clock cycles for TVALID signal.
   * The reference event for this delay is:  #reference_event_for_tvalid_delay
   * - PREV_TVALID_TREADY_HANDSHAKE : Previous tvalid-tready handshake as the reference event
   * - PREV_TVALID                  : Previous tvalid assertion as the reference event
   * .
   * Applicable for ACTIVE MASTER only.
   */
  rand int tvalid_delay[];

  /**
   * @groupname axi4_stream_delays
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * FALSE, this member defines the TREADY signal delay in number of clock
   * cycles.  The reference event for this delay is
   * #reference_event_for_tready_delay.
   *
   * Please note that #reference_event_for_tready_delay is not supported
   * currently. Absolute value of tready_delay is considered for delay
   * calculation with respect to tvalid signal.
   *
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * TRUE, this member defines the number of clock cycles for which TREADY
   * signal should be deasserted after each handshake, before pulling it up
   * again to its default value.
   *
   * Applicable for ACTIVE SLAVE only.
   */
  rand int tready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first wvalid signal. The delay
    * must be programmed in wvalid_delay[0]. Following are the different
    * events under this category:
    *
    * WRITE_ADDR_VALID:
    * Reference event for first WVALID is assertion of AWVALID signal
    * 
    * WRITE_ADDR_HANDSHAKE:
    * This event is applicable when write data is transmitted after write
    * address, that is, when #data_before_addr is set to 0. This reference event
    * specifies the write address handshake.
    * 
    * PREV_WRITE_DATA_HANDSHAKE:
    * This event is applicable when write data is transmitted before write
    * address, that is, when #data_before_addr is set to 1. This reference event
    * specifies the previous write data handshake.
    */
    // removed address handshake refrence because  of potential deadlock due to following reason::
    // the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    //
  rand reference_event_for_first_wvalid_delay_enum reference_event_for_first_wvalid_delay =  WRITE_ADDR_VALID;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_WVALID:
    * Reference event for WVALID delay is assertion of previous wvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts wvalid.
    * 
    * PREV_WRITE_HANDSHAKE:
    * Reference event for WVALID delay is completion of previous data handshake.
    */
  rand reference_event_for_next_wvalid_delay_enum reference_event_for_next_wvalid_delay = PREV_WRITE_HANDSHAKE;

  /**
    *    
    * @groupname axi3_4_delays
    * Defines the reference event for RREADY delay.
    *   
    * RVALID:
    * Reference event for RREADY is assertion of RVALID signal
    * 
    * MANUAL_RREADY: (Not supported currently)
    *
    * This event  allows the user to generate  RREADY patterns, in cycles, as
    * follows:
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The rready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default rready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default rready signal is
    *       driven after toggling
    * 3. The remaining rready_delay element represents no. of cycles to drive
    *    rready
    * 
    * Example 1:
    * For eg.   RREADY  pattern (cycles) =  1110011 and default_rready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_rready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous RREADY value)

    * For eg. cycle pattern  RREADY =  0001100 and default_rready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_rready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous RREADY value)
    */
  rand reference_event_for_rready_delay_enum reference_event_for_rready_delay = RVALID;

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * FALSE, this member defines the BREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_bready_delay.
    * 
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * TRUE, this member defines the number of clock cycles for which BREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int bready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which BREADY should be high and low
    * when the write response channel is idle, that is, when BVALID is low.
    * This property helps to toggle the BREADY signal during the idle period
    * between the assertion of BVALID signal.  The value for this property may
    * be set when the transaction is randomized at the master or in a callback
    * such as svt_axi_port_monitor_callback::write_resp_phase_started. Values
    * provided in even numbered indices indicate the number of clocks for which
    * the ready signal must be driven low and the values in odd numbered
    * indices indicate the number of clocks for which it must driven high.
    * Values in this variable are applicable only until BVALID is asserted.
    * When BVALID is observed on the interface, this delay is no longer
    * applicable. The delay specified in #bready_delay is applied before this
    * attribute is applied.  Note that toggling BREADY during the idle period
    * may lead to situations where the BREADY signal is already asserted when
    * BVALID is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is low. Similarly, BREADY may
    * be low when the corresponding valid is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is high. In both these cases,
    * #bready_delay is not applicable. The size of this array can be set to any
    * value greater than 0, based on the number of times the user would like
    * the signal to toggle during idle period.
    */
  rand int idle_bready_delay[];


  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BREADY delay.
    *
    * BVALID:
    * Reference event is assertion of BVALID signal
    */
  rand reference_event_for_bready_delay_enum reference_event_for_bready_delay = BVALID;

  /**
    * @groupname axi3_4_delays
    * This members applies to AWREADY signal delay for write transactions, and
    * ARREADY signal delay for read transactions.
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is FALSE, this member
    * defines the AWREADY or ARREADY signal delay in number of clock cycles.
    * The reference event used for this delay is
    * #reference_event_for_addr_ready_delay. 
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is TRUE, this member
    * defines the number of clock cycles for which AWREADY or ARREADY signal
    * should be deasserted after each handshake, before pulling it up again to
    * its default value.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  rand int addr_ready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which awready and arready should be
    * high and low when the corresponding address channel is idle, that is,
    * when AWVALID/ARVALID is low. This property helps to toggle the
    * AWREADY/ARREADY signal during the idle period between the assertion of
    * AWVALID/ARVALID signal of this transaction and the next transaction.
    * This value may be assigned during randomization of the transaction object
    * in the slave sequence. Values provided in even numbered indices indicate
    * the number of clocks for which the ready signal must be driven low and
    * the values in odd numbered indices indicate the number of clocks for
    * which it must driven high. Values in this variable are applicable only
    * until the corresponding valid is asserted. When AWVALID/ARVALID is
    * observed on the interface, this delay is no longer applicable and the
    * delay specified in #addr_ready_delay is applied before asserting
    * AWREADY/ARREADY.  Note that toggling AWREADY/ARREADY during the idle
    * period may lead to situations where the AWREADY/ARREADY signal is already
    * asserted when the corresponding valid is sampled, even though the value
    * of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is low. Similarly,
    * AWREADY/ARREADY may be low when the corresponding valid is sampled, even
    * though the value of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is high. In both these
    * cases, #addr_ready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_addr_ready_delay[];


  /** 
    * @groupname axi3_4_delays
    * Defines reference event for AWREADY or ARREADY delay.
    *
    * ADDR_VALID:
    * Reference event is  assertion of AWVALID or ARVALID signal. This event is
    * not applicable when default value of AWREADY = 1 or default value of
    * ARREADY = 1.
    * FIRST_WVALID:
    * Reference event is  assertion of WVALID signal. This event is
    * not applicable when default value of AWREADY = 1.
    * This event is only applicable for write address channel.
    */
  rand reference_event_for_addr_ready_delay_enum  reference_event_for_addr_ready_delay = ADDR_VALID;

  /** 
    * @groupname axi3_4_delays
    * Defines RVALID delay, in terms of number of clock cycles.
    * The reference event for this delay is:
    * - For rvalid_delay[0]        -  #reference_event_for_first_rvalid_delay
    * - For remaining indices of rvalid_delay -  #reference_event_for_next_rvalid_delay
    * .
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int rvalid_delay[];

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * FALSE, this member defines the WREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_wready_delay.
    *
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * TRUE, this member defines the number of clock cycles for which WREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value. 
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which wready should be high and low
    * when the write data channel is idle, that is, when WVALID is low. This
    * property helps to toggle the WREADY signal during the idle period between
    * the assertion of WVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all write data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the write_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transactions unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until WVALID is asserted. When WVALID is observed on the interface,
    * this delay is no longer applicable and the delay specified in
    * #wready_delay is applied before asserting WREADY.  Note that toggling
    * WREADY during the idle period may lead to situations where the WREADY
    * signal is already asserted when the WVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_wready is low. Similarly,
    * WREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_wready is high. In both
    * these cases, #wready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first rvalid signal. The delay
    * must be programmed in rvalid_delay[0]. Following are the different
    * events under this category:
    *
    * READ_ADDR_VALID:
    * Reference event for first RVALID is assertion of ARVALID signal
    *
    * READ_ADDR_HANDSHAKE:
    * Reference event for first RVALID is completion of read address handshake
    */
  rand reference_event_for_first_rvalid_delay_enum reference_event_for_first_rvalid_delay = READ_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the RVALID signals from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_RVALID :
    * Reference event to delay RVALID is assertion of previous rvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts rvalid.
    * 
    * PREV_READ_HANDSHAKE :
    * Reference event to delay RVALID is completion of previous read data
    * handshake.
    */

  rand reference_event_for_next_rvalid_delay_enum reference_event_for_next_rvalid_delay = PREV_READ_HANDSHAKE;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WREADY delay.
    *   
    * WVALID:
    * Reference event for WREADY is assertion of WVALID signal.
    * 
    * MANUAL_WREADY: (Not supported currently)
    * This event  allows the user to generate  WREADY patterns, in cycles, as
    * follows :
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The wready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default wready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default wready signal is
    *       driven after toggling
    * 3. The remaining wready_delay element represents no. of cycles to drive
    *    wready
    * 
    * Example 1:
    * For eg.   WREADY  pattern (cycles) =  1110011 and default_wready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_wready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous WREADY value)

    * For eg. cycle pattern  WREADY =  0001100 and default_wready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_wready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous WREADY value)
    */

  rand reference_event_for_wready_delay_enum  reference_event_for_wready_delay =  WVALID;

  /**
    * @groupname axi3_4_delays
    * Defines the BVALID delay in terms of number of clock cycles. The reference
    * event for this delay is #reference_event_for_bvalid_delay.
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int bvalid_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BVALID delay.
    *
    * LAST_DATA_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for last write
    * data.
    * 
    * ADDR_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for address phase.
    */  

  rand reference_event_for_bvalid_delay_enum reference_event_for_bvalid_delay = LAST_DATA_HANDSHAKE;

  /**
    * @groupname axi4_stream_delays
    * Defines the reference events for TVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_TVALID:
    * In this case, assertion of previous tvalid signal is considered  
    * as the reference event for TVALID delay. The delay timer
    * starts as soon as previous tvalid signal is asserted. If previous
    * tvalid-tready handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts tvalid.
    * 
    * PREV_TVALID_TREADY_HANDSHAKE:
    * Reference event for TVALID delay is completion of previous tvalid-tready handshake.
    */
  rand reference_event_for_tvalid_delay_enum reference_event_for_tvalid_delay = PREV_TVALID_TREADY_HANDSHAKE;

  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the RACK delay should start.
   * - LAST_READ_DATA_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_rack_delay_enum reference_event_for_rack_delay = LAST_READ_DATA_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the RACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_rack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int rack_delay = 0;
  
  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the WACK delay should start.
   * - WRITE_RESP_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_wack_delay_enum reference_event_for_wack_delay = WRITE_RESP_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the WACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_wack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int wack_delay = 0;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the delay between reception of DVM Sync and transmission of DVM Complete.
   * Delay for master component in terms of number of clock cycles for generating
   * DVM Complete transaction after receiving a DVM Sync transaction. 
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int dvm_complete_delay = 0;

  /**
   *  @groupname out_of_order
   *  Sets the reordering priority of the current transaction within the set
   *  of transactions that are allowed access to read data channel based on 
   *  svt_axi_port_configuration::read_data_reordering_depth.
   * 
   *  This member is applicable only when svt_axi_port_configuration::reordering_algorithm
   *  is svt_axi_port_configuration::PRIORITIZED.
   * 
   *  This value indicates the priority of sending the response to current 
   *  transaction compared to remaining transactions within the depth indicated
   *  by svt_axi_port_configuration::read_data_reordering_depth for read transactions or
   *  by svt_axi_port_configuration::write_resp_reordering_depth for write transactions.
   *
   *  Note that the value of this attribute should be within the following range:
   *  [1:svt_axi_port_configuration::read_data_reordering_depth] for read transactions and
   *  [1:svt_axi_port_configuration::write_resp_reordering_depth] for write transactions.
   * 
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘1’ then, the
   *  transactions with highest value for this attribute will get higher priority.
   *
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘0’ then, the
   *  transactions with least value for this attribute will get higher priority.
   *
   *  If there are more than one transactions with same priority, those transaction
   *  will be processed in the same order as they are received.
   * 
   * Applicable for ACTIVE SLAVE only.
   */

  rand int reordering_priority = 1;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of zero delay within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int ZERO_DELAY_wt = 100;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of short delays within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int SHORT_DELAY_wt = 500;

  /**
    * @groupname axi3_4_delays
    * Weight used to control distribution of long delays within transaction generation.
    *
    * This controls the distribution of delays for the 'delay' fields 
    * (e.g., delays for asserting the ready signals).
    */
  int LONG_DELAY_wt = 1;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of burst length to 1 within transaction
     * generation.
     *
     * This controls the distribution of the length of the bursts using
     * burst_length field 
     */
  int ZERO_BURST_wt = 100;

   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of short bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int SHORT_BURST_wt = 500;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of longer bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int LONG_BURST_wt = 400;


  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

   /**
    * @groupname axi4_stream_protocol
    * Used to drive TDATA signals. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
   rand bit [`SVT_AXI_MAX_TDATA_WIDTH - 1:0] tdata[];

  
  /**
   * @groupname axi4_stream_protocol
   * Used to drive TSTRB signal. The strobes are right aligned and the model
   * will drive strobes on appropriate lanes. The model also takes care of the
   * endianness while driving tstrb. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TSTRB_WIDTH - 1:0] tstrb[];

 
  /**
   * @groupname axi4_stream_protocol
   * TKEEP is the byte qualifier that indicates whether the content of the
   * associated byte of TDATA is processed as part of the data stream.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TKEEP_WIDTH - 1:0] tkeep[];


  /**
    * @groupname axi4_stream_protocol
    * The variable holds the value of  TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand bit [`SVT_AXI_MAX_TID_WIDTH - 1:0] tid = 0;
  
  /**
    * @groupname axi4_stream_protocol
    * TDEST provides routing information for the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TDEST_WIDTH - 1:0] tdest;
  
  /**
    * @groupname axi4_stream_protocol
    * TUSER is user defined sideband information that can be transmitted
    * alongside the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TUSER_WIDTH - 1:0] tuser[];

  /**
    * @groupname axi4_stream_protocol
    * Defines the burst length of a AXI4 Stream Packet. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand int stream_burst_length = 1;

  // ****************************************************************************
  // End of STREAM SIGNALS
  // ****************************************************************************
  /**
    * @groupname axi3_protocol
    * A bit that must be set by the user to indicate that this transaction will
    * be sent to the slave driver from the slave sequencer through the
    * delayed_response_request_port of the slave driver. If the transaction is
    * randomized before putting it into the delayed_response_request_port of the
    * slave driver, then this bit must be set by the user. This bit must not be
    * set for a transaction that is sent on the seq_item_port.
    */
  bit is_delayed_response_xact = 0;

  /**
   * @groupname axi_misc
   * Indicates the value of the source master which will be propogated in the ID field
   * of the master and the corresponding slave transaction.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::source_master_id_xmit_to_slaves_type is set to
   * DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES. This property must be set by the
   * user in a system monitor callback issued at the start of a transaction
   */
  bit[`SVT_AXI_DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES_WIDTH-1:0] dynamic_source_master_id_xmit_to_slaves = 0;

  /**
   * @groupname axi_misc
   * Indicates that this master transaction is a partial write transaction and this
   * transaction will be split by the interconnect into a full Read transaction
   * followed by partial Write transaction to the corresponding slave.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::partial_write_to_slave_read_and_write_association_enable is set to
   * This property must be set by the user in a system monitor callback issued at the start of a transaction
   */
  bit partial_master_write_split_into_read_modified_write_slave_xact = 0;

  /**
   * @groupname axi_misc
   * Multibit array for different usages.
   * 
	 * If cust_xact_flow[0] is set to '1', indicate that transaction should be drived immediately on the interface.
	 * This is aplicable only for AXI4 STREAM transactions.
	 *
	 * cust_xact_flow[31:1] bits are for future use.
   */
  rand bit[31:0] cust_xact_flow = 0;  

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * A bit that is set by the slave driver to indicate that the write response
    * of a transaction has been provided by the user through the
    * delayed_response_request_port of the slave driver.  
    * Applicable only when
    * svt_axi_port_configuration::enable_delayed_response_port is set.
    */
  bit is_delayed_write_response_set = 0;

  /** 
    * @groupname ace_l3_cache
    * Inidcates that current transaction will cause memory update transaction for the associated
    * cacheline if it is  hit in L3 and found to be in dirty state.
    */
  bit clean_l3_data = 0;

  /** 
    * @groupname ace_l3_cache
    * This attribute is supposed to be updated by VIP indicating to the user that memory has been
    * updated for the current transaction with associated cacheline data in L3 cache. This is primarily
    * used along with clean_l3_data i.e. if current transaction is expected to update memory then user
    * can wait for this attribute to be set by VIP if user needs to perform any tasks based on that condition.
    */
  bit mem_updated_with_l3_data = 0;
  /** @endcond */

  `ifdef SVT_ACE5_ENABLE  
  /**
    * @groupname axi5_protocol
    * Defines the chunk enable of a AXI5 to enable read_data_chunking. When enable, slave will send read data
    * in 128bits of chunk in random order. If disabled, slave will send read data without chunking as per AXI5 protocol. Applicable 
    * when svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit archunken = 0;

  /**
    * @groupname axi5_protocol
    * Array of read chunk strobe
    * Each bit of rchunkstrb represents 128bits of read data. Width of the rchunkstrb by default is 
    * `SVT_AXI_MAX_CHUNK_STROBE_WIDTH user can change width using svt_axi_port_configuration::rchunkstrb_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1 : 0] rchunkstrb[];

  /**
    * @groupname axi5_protocol
    * Array of read chunk number
    * Indicates that the data chunk number is being transferred. Width of the rchunknum by default is 
    * `SVT_AXI_MAX_CHUNK_NUM_WIDTH user can change width using svt_axi_port_configuration::rchunknum_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_NUM_WIDTH -1 : 0] rchunknum[];

  /**
    * @groupname axi5_protocol
    * Indicates that the data chunk length is being transferred. This signal is for interal use to calculate number  
    * of transafer for chunkinig Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable 
    * is set to 1.
    * Not yet implemented. 
    */
  rand int chunk_length;

  /**
   * @groupname axi5_protocol
   *    This is a counter which is incremented for every chunk of databeat. Useful when user
   *    would try to access the transaction class to know its current state during chunking.
   *    This represents the chunk databeat transfer number.
   */
  int  current_data_chunk_trf_num = 0;
  `endif  

  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

  `ifdef SVT_AXI_QVN_ENABLE
  /**
   * @groupname qvn_parameters
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to AXI3/AXI4/ACE/ACE_LITE
   * Specifies the Virtual Network ID to which token for this transaction will be requested.
   * Same Virtual Network will be used to send current transaction as well. 
   *
   * Active Master will use qvn_vnet_id to determine which VN*VALID* signal needs to be asserted
   * to request for token and all ARVNET_ID or AWVNET_ID and WVNET_ID value will be driven
   * same as qvn_vnet_id
   *
   * Port Monitor will use qvn_vnet_id to indicate from which Virtual Network this particular 
   * transaction has been received.
   *
   */
  rand int qvn_vnet_id = 0;
  `endif

  `ifdef SVT_AXI_CUSTNV_ENV
  /** 
    * configuration register used to provide custom L3 or interconncet based behaviour
    * [0] = '1' indicates writeEvict can start from shared state.
    * [1] = '1' indicates no data has been provided as part of the read response.
    * [2] = '1' indicates current transaction is a block linear request.
    * [3] = '1' indicates current transaction is auto-generated by VIP for an origninal block linear request.
    *           this bit is supposed to get set by VIP. User doesn't need to set this bit.
    *
    * default value of all fields are 0 and it is set by user except bit[3].
    */
  bit[31:0] custnv_reg = 0;
  `endif
  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  local static vmm_log shared_log = new("svt_axi_transaction", "class" );
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
  local svt_axi_port_configuration::axi_port_kind_enum axi_port_kind = svt_axi_port_configuration::AXI_MASTER;

  local svt_axi_port_configuration::axi_interface_type_enum axi_interface_type = svt_axi_port_configuration::AXI3; 
`endif

  /** @cond PRIVATE */
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_data_width_in_bytes = 0;
  
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int data_width_in_bytes = 0;
 
  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH/8 -1 :0] atomic_read_poison_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_comp_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_cache_line_size = 0;

  /** internal flag to track if transaction is part of a multi-part dvm sequence */

  bit is_part_of_multipart_dvm_sequence = 0;

  /** The channel (READ/WRITE) on which this transaction will be transmitted */
  xact_type_enum transmitted_channel = WRITE;

  /** The xact_type when port_cfg is_downstream_coherent = 1 */
  xact_type_enum converted_xact_type = WRITE; 
  /** @endcond */
 
  // ****************************************************************************
  // Local variables only for internal VIP usages
  // ****************************************************************************
  bit [(`CEIL(`SVT_AXI_MAX_ID_WIDTH,8))-1:0] axidchk_parity_value = 0;
  bit [(`CEIL(`SVT_AXI_MAX_ADDR_WIDTH,8))-1:0] axaddrchk_parity_value = 0;
  bit axlenchk_parity_value  = 0;
  bit axctlchk0_parity_value = 0;
  bit axctlchk1_parity_value = 0;
  bit axctlchk2_parity_value = 0;
  bit arctlchk3_parity_value = 0;
  bit [(`CEIL((`SVT_AXI_MAX_DATA_WIDTH/8),8))-1:0]       wstrbchk_parity_value;

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZRypSBVsMJ/hicVIQ44U92je/RbUHxjfvU8fW5zht/GTH0Z+Qsdjx/TVos0EUbrG
fcpgCkQOvjOuVuz093DSa/VIzgCS4fH9FKyjUc0wUSpA4O9Gt8qw6DdKxUqIOigZ
f7f0TL8JU25B8CGLxFAoIktPjK1bxQHnXVuVVa1gNAu8CBaBLhC7bQ==
//pragma protect end_key_block
//pragma protect digest_block
CiWQwzjjHvnFosF0i+JK7jH2mMM=
//pragma protect end_digest_block
//pragma protect data_block
+R79qwVWi4RPnkudTWz27ZYysX9neBDWBtPsrALVc1TZC4OsU4DEhtVEAPfcFy6F
9NYof5CaIYuyOQ0GG2o5o2iJTQ4mLziyCp1Voln9G14ez9w0DnGvDWK8QxwbHx17
URiUeWNnu6jdm2enSS/NvAB7GqddupNUXsm2qJJrHzodxju0gql7sm6Jq+OTe6yW
i3FC5VHb2tsglBmE83WpoNcq6XGLGvFcZKQiM5ePTWxeg4zWag6bTjx2yZPKNpe8
uVes+S6IcXj6UTKuav3HGH7UbBo9ZX/KhrGjwA0NU2Pghf7z6DPvJ3aCjwmydPFh
wJ4dc7tA7a1thjVSFcXjnsW2776KXEMm/Y0rHA6SfZyH7bOUMJkGwUWZb2Kl0dat
040/o9NIziTmSWPyncMsdGIV8kmg4NVBTJMiZkalvY7DAvnnGgrd9kx3TsQlO/Yb
3KMsAa8+UFtuhER+/YrkFQeIYtEr+EroqMyej/P1I6y7P9fksXziZ3+Zz7bIocic
ziiLcGSMrYvER04ElTPr7NGkzeDgMDr5u30LoYZvtrr4Wfqk5dnQ+jmUn33BaSh3
JOeBzSo4fuyi2tfmkfSBqvObapjvWlEQ+1SYtKVSdRj0GGYDQt24CPHWvOHspBWv
BDNFNZRoBy/gX+CqJnSZ1w==
//pragma protect end_data_block
//pragma protect digest_block
5r0S80I+ECpf91aaQhOTwMiBh9A=
//pragma protect end_digest_block
//pragma protect end_protected
  
  /** Re-organised constraint blocks based on interface type. This will make
   * it easy to turn-off the constraints based on interface type. It can
   * result in significant run-time improvement. */

  // QVN Constraints Block. These constraints are valid when QVN mode is
  // enabled. 
  constraint qvn_valid_ranges {
`ifdef SVT_AXI_QVN_ENABLE
    solve xact_type before qvn_vnet_id;
    solve coherent_xact_type before qvn_vnet_id;

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
    if(port_cfg.qvn_enable) {
        // -------------------------------------------------------------------------------
        // Each Transaction should pick Virtual Network only from the list of supported VN
        // -------------------------------------------------------------------------------
        qvn_vnet_id inside {[0:`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1]};

        if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) ) {
          foreach(port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) -> qvn_vnet_id != ix;
          }
        } else {
          foreach(port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) -> qvn_vnet_id != ix;
          }
        }
        // -------------------------------------------------------------------------------
    }
    else {
       qvn_vnet_id == 0;
    }
`endif // SVT_AXI_SVC_NO_CFG_IN_XACT
`endif // SVT_AXI_QVN_ENABLE
  } // qvn_valid_ranges

// These constraints are applicable for Memory tagging feature
 constraint memory_tagging_valid_ranges {
`ifdef SVT_ACE5_ENABLE
 if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER){
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(transmitted_channel == WRITE || transmitted_channel == READ_WRITE) {
     if(port_cfg.mte_support_type == svt_axi_port_configuration::BASIC){
       !tag_op inside {TAG_TRANSFER,TAG_FETCH_MATCH};
       if(xact_type == ATOMIC){
         tag_op == TAG_INVALID;}
    if(xact_type == COHERENT)  {
      if(coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE}){
       tag_op  inside {TAG_INVALID,TAG_UPDATE}; }
      else if (coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
      tag_op ==TAG_INVALID;}
     }
   if(xact_type == WRITE){
     tag_op  inside {TAG_INVALID,TAG_UPDATE};}
   }
   if(port_cfg.mte_support_type == svt_axi_port_configuration::STANDARD){
     tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
      if(xact_type == ATOMIC){
         tag_op inside {TAG_INVALID,TAG_FETCH_MATCH};}
      if(xact_type == COHERENT)  {
        if(coherent_xact_type == WRITENOSNOOP){
          tag_op  inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};}
        else if(coherent_xact_type inside {WRITEUNIQUE,WRITELINEUNIQUE}) {
          tag_op  inside {TAG_INVALID,TAG_UPDATE};}
        else if (coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO}){
          tag_op inside {TAG_INVALID,TAG_TRANSFER,TAG_UPDATE};}
        else if (coherent_xact_type inside{CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
          tag_op == TAG_INVALID;}
         }
       if(xact_type == WRITE){
         tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
        }
       }
     }
  if(transmitted_channel == READ) {
    tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH};
    if(xact_type == COHERENT)  {
      if(coherent_xact_type == READNOSNOOP){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
      else if (coherent_xact_type == READONCE){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER};}
      else if (coherent_xact_type inside {READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE}){
      tag_op ==TAG_INVALID;}
    }
   if(xact_type == READ){
      tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
  }
  if (tag_op != TAG_INVALID){
  // Transactions must be cacheline sized or smaller
  //For an INCR burst, the last byte in the burst, as determined from the burst length in bytes,
  //(AWSIZE x AWLEN), added to the AWSIZE aligned start address, must be within the same
  //cache line as the first byte in the burst
  //i.e addr_aligned_to_burst_size + bytes_in_transfer < addr_aligned_to_cache_line_size + cache_line_size
      (burst_type == INCR) -> (((addr >> burst_size) << burst_size) + (burst_length << burst_size) <= 
      ((addr >> log_base_2_cache_line_size) << log_base_2_cache_line_size) + port_cfg.cache_line_size);
   // For a WRAP burst, AWSIZE x AWLEN must not exceed the cache line size.
      (burst_type == WRAP) -> ((burst_length << burst_size) <= port_cfg.cache_line_size);

 // For INCR transactions address must be aligned to container size
    if(burst_type == INCR){
     addr == addr >> (burst_length << burst_size) << (burst_length << burst_size);
    }

  // For WRAP transactions address must be aligned to burst_size
    if(burst_type == WRAP){
      addr == addr >> burst_size << burst_size; }

    cache_type[3:2] != 2'b00;
    cache_type[1:0] == 2'b11; 
   }
  if(tag_op == TAG_INVALID){
    foreach(tag[i])
      tag[i] == 0;}

  // Transaction type inside READ,WRITE,COHERENT and ATOMIC  
  xact_type inside {READ,WRITE,COHERENT,ATOMIC};
  if(xact_type == COHERENT){
    coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE,CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION,WRITEPTLCMO,WRITEFULLCMO,
                                READNOSNOOP,READONCE,READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE};
  }
  }
}
// constraints on response_tag_op only applicable in external port monitor mode
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE){
     if(port_cfg.use_external_port_monitor == 1){
       if(transmitted_channel == READ){
         if(tag_op == TAG_INVALID){
          response_tag_op inside {TAG_INVALID,TAG_TRANSFER};}
         else if(tag_op == TAG_TRANSFER){
         response_tag_op == TAG_TRANSFER};
        }
       else if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
         response_tag_op == TAG_INVALID;
       }
     }
     else {
       response_tag_op == TAG_INVALID;
     }
     if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
      tag_match_resp inside{ MATCH_NOT_PERFORMED,NO_MATCH_RESULT,FAIL, PASS};
     }
     else if(transmitted_channel == READ){
      tag_match_resp == MATCH_NOT_PERFORMED;
     }
   }
 }
`endif
 }

// These constraints are applicable for MPAM feature
constraint mpam_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if (port_cfg.enable_mpam == svt_axi_port_configuration::MPAM_FALSE && port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER && port_cfg.is_active) {
    mpam_partid == 0;
    mpam_perfmongroup == 0;
    mpam_ns == prot_type[1];
  } 
`endif
}

// These constraints are applicable for Write with CMO transactions 
 constraint write_with_cmo_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if(xact_type == COHERENT && (coherent_xact_type == WRITEPTLCMO || coherent_xact_type == WRITEFULLCMO)){
    domain_type inside {INNERSHAREABLE,OUTERSHAREABLE,NONSHAREABLE};
    atomic_type == NORMAL;
    cache_type[1] == 1;
  }
 if(port_cfg.axi_interface_type != svt_axi_port_configuration::ACE_LITE){
   !(coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO});
  } 
 if(port_cfg.write_plus_cmo_enable != 1){
    !(coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO});
  }
 if(port_cfg.cmo_on_write_enable != 1){
   coherent_xact_type != CMO;
 }
`endif
 }
 //These constraints are valid for atomic transactions .
constraint atomic_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE 
   if(!port_cfg.axi_interface_type inside{svt_axi_port_configuration::AXI4,svt_axi_port_configuration::ACE_LITE})  {
      xact_type != ATOMIC;}
//   if(port_cfg.check_type != svt_axi_port_configuration::ODD_PARITY_BYTE_DATA){
//      atomic_read_is_datachk_parity_error == 0;}
   if(xact_type ==ATOMIC){
  //  data size should be equal to burst length
     if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
      
      if((barrier_type == NORMAL_ACCESS_RESPECT_BARRIER) || (barrier_type == NORMAL_ACCESS_IGNORE_BARRIER)){ 
          if ((domain_type == NONSHAREABLE) || (domain_type == SYSTEMSHAREABLE)){
             coherent_xact_type  == WRITENOSNOOP;}
          else{
             coherent_xact_type  == WRITEUNIQUE;}
        }
        else{
           coherent_xact_type == WRITEBARRIER;}
       if(burst_length > 1 && ! port_cfg.allow_multibeat_atomic_transactions_to_be_less_than_data_width){
         (1 << burst_size) == port_cfg.data_width/8;
       }
       data.size() == burst_length;
       wstrb.size() == burst_length;
       if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] == ((1 << (1 << burst_size)) - 1);
        }
      }
      awakeup_assert_delay ==0;
       if( atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN}){
          atomic_transaction_type == LOAD;
         }
       if(atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN}) {
          atomic_transaction_type == STORE;
        }
       if(atomic_xact_op_type == ATOMICSWAP){
          atomic_transaction_type == SWAP;
        }
       if(atomic_xact_op_type == ATOMICCOMPARE){
         atomic_transaction_type == COMPARE;
         burst_size inside{0,1,2,3,4,5};
         {((1 << burst_size)) * burst_length} inside {2,4,8,16,32};
         if(burst_length << burst_size == 2 && addr[0]==1'b0){ 
           burst_type == INCR;}
         else if(burst_length << burst_size == 4 && addr[1:0]==2'b0) {
            burst_type == INCR;}
         else if(burst_length << burst_size == 8 && addr[2:0]==3'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 16 && addr[3:0]==4'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 32 && addr[4:0]==5'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 2 && addr[0] !=1'b0){
           burst_type == WRAP;}
         else if(burst_length << burst_size == 4 && addr[1:0] !=2'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 8 && addr[2:0] !=3'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 16 && addr[3:0] !=4'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 32 && addr[4:0] !=5'b0) {
           burst_type == WRAP;}
          } 
        atomic_transaction_type != NON_ATOMIC;
        if(atomic_transaction_type == COMPARE ){
           atomic_swap_data.size() == burst_length;
           atomic_compare_data.size() == burst_length;
           atomic_compare_wstrb.size() == burst_length;
           atomic_swap_wstrb.size() == burst_length;
           foreach(atomic_swap_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_swap_data[index] == atomic_swap_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           foreach(atomic_compare_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_swap_data[index]) {
               atomic_swap_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_compare_data[index]) {
               atomic_compare_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
        }
        else {
           atomic_swap_data.size() == 0;
           atomic_compare_data.size() == 0;
           atomic_compare_wstrb.size() ==0;
           atomic_swap_wstrb.size() ==0;
         }
         if(atomic_transaction_type ==LOAD){
           atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN};}
         else if(atomic_transaction_type ==STORE){
           atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN};}
         else if(atomic_transaction_type ==SWAP){
           atomic_xact_op_type inside{ATOMICSWAP};}
         else if(atomic_transaction_type ==COMPARE){
           atomic_xact_op_type inside{ATOMICCOMPARE};}

//     Address for atomic transactions must be aligned to the data size
         if(atomic_transaction_type !=COMPARE){
           burst_size inside {0,1,2,3};
           {((1 << burst_size)) * burst_length} inside {1,2,4,8};
           burst_type==INCR;
           if (burst_length << burst_size == 2) {
              addr[0] == 1'b0;
            } 
            else if (burst_length << burst_size == 4) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 8) {
              addr[2:0] == 3'b0;
            } 
          }
//   For an Atomic compare transactions address must be aligned to half of the burst_size
         else if(atomic_transaction_type == COMPARE){
           burst_size inside {0,1,2,3,4,5};
            if(burst_length << burst_size == 4){
              addr[0] == 1'b0;}
            else if (burst_length << burst_size == 8) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 16) {
              addr[2:0] == 3'b0;
            } 
           else if(burst_length << burst_size == 32){
              addr[3:0] == 4'b0;
           }
         }

       if(atomic_transaction_type == COMPARE) {
         atomic_swap_wstrb.size() == burst_length;
         atomic_compare_wstrb.size() == burst_length;
         }
       else {
         atomic_swap_wstrb.size() == 0;
         atomic_compare_wstrb.size() == 0;
       }
     if(atomic_transaction_type != COMPARE){
         burst_type == INCR;
         burst_size inside {0,1,2,3};
        }
       else if(atomic_transaction_type == COMPARE){
         burst_type inside{INCR,WRAP};
         burst_size inside{0,1,2,3,4,5};
        }
         if(xact_type ==ATOMIC){
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
         }
    }

  /* 
   * 1) Constraint the atomic_read_data_trace_tag to 1 based on trace_tag value
   */
    if(port_cfg.axi_port_kind == svt_axi_port_configuration:: AXI_SLAVE){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
       if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        atomic_read_data.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
        atomic_read_poison.size() == burst_length;

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}

      }
      if(atomic_transaction_type == COMPARE && xact_type ==ATOMIC){
        if(burst_length > 1){
          atomic_read_data.size() == burst_length/2;
          atomic_read_data_user.size() == burst_length/2;
          atomic_read_poison.size() == burst_length/2;
        }
        else {
          atomic_read_data.size() == 1;
          atomic_read_data_user.size() == 1;
          atomic_read_poison.size() == 1;
        }

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_comp_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_comp_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}
        }

      if(trace_tag ==1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        atomic_read_data_trace_tag == 1;
       }
      if(atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        rvalid_delay.size() == burst_length;
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};
            }
       wready_delay.size()==burst_length;
    }

  }
    if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
     }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE} ){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
    
/*     if(xact_type == ATOMIC) {
       if(burst_length > 1){
          1 << burst_size == data_width_in_bytes;}
      }*/
  if(xact_type != ATOMIC)
    {
       atomic_read_data.size() ==0;
       atomic_read_poison.size() ==0;
       atomic_read_data_user.size() ==0;
       atomic_swap_data.size() ==0;
       atomic_compare_data.size() ==0;
       atomic_swap_wstrb.size()==0;
       atomic_compare_wstrb.size()==0;
       atomic_transaction_type == NON_ATOMIC;
    }
   if(xact_type ==ATOMIC){
     atomic_type == NORMAL;
     random_interleave_array.size() == burst_length;
     random_interleave_array[0] == 1;
    }
     xact_type != READ_WRITE;
     converted_xact_type != READ_WRITE;
     transmitted_channel != ATOMIC;
`endif
}

  // ACE/ACE-Lite Constraints Block. These constraints are valid if the
  // interface type is set to ACE or ACE-Lite.

  constraint ace_valid_ranges {

    foreach(data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
    }

`ifdef SVT_ACE5_ENABLE
   if(port_cfg.atomic_transactions_enable ==1'b1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC) {
      foreach(atomic_read_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data[index] == atomic_read_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

      foreach(atomic_read_data_user[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data_user[index] == atomic_read_data_user[index] & ((1<<(port_cfg.data_width))-1);}
    }

     foreach(atomic_swap_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_swap_data[index] == atomic_swap_data[index] & ((1<<((port_cfg.data_width)))-1);}
    }
      foreach(atomic_compare_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

   if(port_cfg.poison_enable ==1 && port_cfg.wysiwyg_enable ==1){
       foreach(atomic_read_poison[index]) {
         if(port_cfg.data_width%64 == 0) {
           atomic_read_poison[index] == atomic_read_poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
           atomic_read_poison[index] == atomic_read_poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
   }}
  }
`endif

 if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
         if(port_cfg.data_width%64 == 0) {
            poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
            poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
    }}
   }
   
`ifdef SVT_ACE5_ENABLE
// This transaction types are not yet supported  
   !(coherent_xact_type inside {STASHTRANSLATION});
`endif 

`ifdef SVT_AXI_SVC_USE_MODEL
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration :: AXI_ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
   }
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
`ifdef INCA
     if ((slave_xact_type == COHERENT) && (slave_xact_type != DATA_STREAM )) {
        if( 
            (slave_coherent_xact_type == CLEANUNIQUE) || 
            (slave_coherent_xact_type == MAKEUNIQUE) || 
            (slave_coherent_xact_type == CLEANSHARED) ||
            (slave_coherent_xact_type == CLEANSHAREDPERSIST) ||
            (slave_coherent_xact_type == CLEANINVALID) || 
            (slave_coherent_xact_type == MAKEINVALID) 
          ) {
          wready_delay.size() == 1;
          rvalid_delay.size() == 1;
        }
        else {
          wready_delay.size() == burst_length;
          rvalid_delay.size() == burst_length;
        }
     }
`else  
     if ((xact_type == COHERENT) && 
         (xact_type != DATA_STREAM)) {
       if( 
           (coherent_xact_type == CLEANUNIQUE) || 
           (coherent_xact_type == MAKEUNIQUE) || 
           (coherent_xact_type == CLEANSHARED) || 
           (coherent_xact_type == CLEANSHAREDPERSIST) ||
           (coherent_xact_type == CLEANINVALID) || 
           (coherent_xact_type == MAKEINVALID) 
         ) {
         wready_delay.size() == 1;
         rvalid_delay.size() == 1;
       } else {
         wready_delay.size() == burst_length;
         rvalid_delay.size() == burst_length;
       }
     }  
`endif // `ifdef INCA 
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
   } //       if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE)
`endif //SVT_AXI_SVC_USE_MODEL
 } // ace_valid_ranges

  // AXI4 STREAM Constraints Block. These constraints are valid if the
  // interface type is set to AXI4_STREAM.
  constraint axi4_stream_valid_ranges {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif   
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
        random_interleave_array.size() == stream_burst_length;
        foreach (random_interleave_array[index]) {
          random_interleave_array[index] inside {[1 : stream_burst_length]};
        }   
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM)
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tid_enable) {
`else
       if (!port_cfg.tid_enable) {
`endif
         tid == 0;
       }
       else {
         tid inside {[0 : ((1 << port_cfg.tid_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdest_enable) {
`else
       if (!port_cfg.tdest_enable) {
`endif
         tdest == 0;
       }
       else {
         tdest inside {[0 : ((1 << port_cfg.tdest_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdata_enable) {
`else
       if (!port_cfg.tdata_enable) {
`endif
         foreach (tdata[index])
           tdata[index] == 0;
       }
       else {
         foreach (tdata[index]) {
             tdata[index] inside {[0 : ((1 << port_cfg.tdata_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tstrb_enable) {
`else
       if (!port_cfg.tstrb_enable) {
`endif
         foreach(tstrb[index])
           tstrb[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tuser_enable) {
`else
       if (!port_cfg.tuser_enable) {
`endif
         foreach(tuser[index])
           tuser[index] == 0;
       }
       else {
         foreach (tuser[index]) {
            tuser[index] inside {[0 : ((1 << port_cfg.tuser_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tkeep_enable) {
`else
       if (!port_cfg.tkeep_enable) {
`endif
         foreach(tkeep[index])
           tkeep[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tlast_enable) {
`else
       if (!port_cfg.tlast_enable) {
`endif
         stream_burst_length == 1;
       }
     } //AXI4_STREAM
   } //AXI_MASTER    
  } // axi4_stream_valid_ranges  


  // AXI3/AXI4/AXI4 Lite Constraints Block. These constraints are valid if the
  // interface type is set to either AXI3/AXI4/AXI4_Lite. Since these are
  // basic AXI constraints they even hold true in case the interface_type is
  // set to ACE/ACE_Lite.

  constraint axi3_4_valid_ranges {
    /*solve burst_length before random_interleave_array;
    solve stream_burst_length before random_interleave_array;
    solve burst_length before addr;
    solve burst_length before wstrb;

    solve burst_size before wstrb;
    solve burst_length before rresp;
    solve burst_length before coh_rresp;
    solve burst_length before rvalid_delay;
    solve burst_length before wready_delay;
    solve xact_type before rvalid_delay;
    solve xact_type before wready_delay;
    solve coherent_xact_type before rvalid_delay;
    solve coherent_xact_type before wready_delay;
    solve xact_type before rresp;
    solve coherent_xact_type before rresp;
    solve xact_type before coh_rresp;
    solve coherent_xact_type before coh_rresp;
    */

  foreach(data[index]) {
     if(port_cfg.wysiwyg_enable ==1'b1){
       data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
   }

   if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
      }
    }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
    burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
`else
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI3)
      burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
    else
      burst_length <= `SVT_AXI4_MAX_BURST_LENGTH;
`endif //SVT_AXI_SVC_NO_CFG_IN_XACT
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_USE_MODEL

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
      // Constraining the Delay sizes
      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        wvalid_delay.size() == 1;
        rready_delay.size() == 1;
        data.size() == 1;
        if(port_cfg.poison_enable ==1){
        poison.size() == 1;}
      } else if (xact_type != DATA_STREAM) {
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
        data.size() == burst_length;
       if(port_cfg.poison_enable ==1){
       poison.size() == burst_length;
      }}

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (port_cfg.toggle_ready_signals_during_idle_period) {
        if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          idle_rready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY_ARR_SIZE]};
          idle_bready_delay.size() == 0;
        } else {
          idle_bready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY_ARR_SIZE]};
          idle_rready_delay.size() == 0; 
        }
      } else {
        idle_rready_delay.size() == 0;
        idle_bready_delay.size() == 0;
      }

     if (!port_cfg.wysiwyg_enable) {
        foreach (data[index]) {
          data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        } 
      }
     foreach(data[index]) {
       if(port_cfg.wysiwyg_enable ==1'b1){
         data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
      }

    if(port_cfg.poison_enable ==1 && !port_cfg.wysiwyg_enable){
        foreach (poison[index]) {
          if((1 << burst_size)%8 !=0){
            poison[index] <= ((1 << (((1 << burst_size) >> 3)+1)) - 1);}
          else {
             poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);}
        } 
      }

   if(port_cfg.poison_enable ==1  && port_cfg.wysiwyg_enable ==1){
      foreach(poison[index]) {
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
    }
`endif

      /*
       * 1) Constrain the array size to 0 if xact_type is not READ
       * 2) Constrain the array size to burst length if xact_type is READ
       */    
      if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
        if (`SVT_AXI_COHERENT_READ_1_BEAT) 
          rresp.size() == 1;
        else
          rresp.size() == burst_length; 
      }
`ifdef SVT_ACE5_ENABLE
     else if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
      }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE}){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
`endif      
      else {
        rresp.size() == 0;
      }

      /* 
       *  Constraints for wstrb 
       *  1) Constraint the length of the wstrb from 1 to burst_length for write
         transactions
       *  2) Constraining wstrb to enable all the valid bytelanes depending on transfer
      */
      if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) 
`ifdef SVT_ACE5_ENABLE
|| xact_type ==ATOMIC
`endif    
       ) {
        wstrb.size() == burst_length;
      }
      else
        wstrb.size() == 0;
      /*if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] inside {[0: ((1 << (1 << burst_size)) - 1)]};
        }
      }
      */
`ifdef SVT_ACE5_ENABLE
       if(xact_type == ATOMIC){
          data.size() == burst_length;
       }
`endif

      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        data_user.size() == 1;
      } else if (xact_type == DATA_STREAM) {
        data_user.size() == 0;
      } else {
        data_user.size() == burst_length;
      }
`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
`ifdef SVT_ACE5_ENABLE 
    xact_type inside {READ,WRITE,IDLE,COHERENT,ATOMIC};
`else
    xact_type inside {READ,WRITE,IDLE,COHERENT,DATA_STREAM};
`endif
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        xact_type != DATA_STREAM;

`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
        atomic_type inside {NORMAL,EXCLUSIVE,LOCKED};
        burst_type inside {FIXED,INCR,WRAP};
`endif

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
        /* 
         * The atomic type is not exclusive when exclusive_access_enable is
         * disabled
         */  
        if (port_cfg.exclusive_access_enable == 0) {
          atomic_type != EXCLUSIVE;    
        }
        if (port_cfg.locked_access_enable == 0) {
          atomic_type != LOCKED;    
        }
`endif
        
        
        /** Address is within limits specified by addr_width. */
        addr <= max_possible_addr;
        addr_user <= max_possible_user_addr;

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        id <= ((1 << `SVT_AXI_MAX_ID_WIDTH) - 1);
`else
        if (port_cfg.use_separate_rd_wr_chan_id_width == 0 
`ifdef SVT_ACE5_ENABLE
          || xact_type == ATOMIC
`endif
         ) 
          id <= ((1 << port_cfg.id_width) - 1);
        else if ((xact_type == WRITE) || `SVT_AXI_COHERENT_WRITE)
          id <= ((1 << port_cfg.write_chan_id_width) - 1);
        else 
          id <= ((1 << port_cfg.read_chan_id_width) - 1);
`endif

        /*
         *  When the burst type is not Fixed, it must be ensured that burst does not
         *  exceed 4k range
         */
   
        if(burst_type != FIXED) {
          addr_range == (burst_length * (1 << burst_size));
          `ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
          addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << burst_size);
          `else
          addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << burst_size);
          `endif  
          if (burst_type == WRAP) {
            // Make sure that the max address does not cross addr_width.
            // Need to calculate this from wrap boundary (lowest address)
            // Note that the max byte address is:
            // (burst_length-1)*bytes_in_each_transfer + (bytes_in_each_transfer-1)
            if (burst_length == 2)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+1));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+1));
`endif
            else if (burst_length == 4)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+2));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+2));
`endif
            else if (burst_length == 8)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+3));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+3));
`endif
            else if (burst_length == 16)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+4));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+4));
`endif

            addr == (addr & addr_mask);
            (addr & burst_addr_mask) + addr_range - 1 <= max_possible_addr; 
            (addr[11:0] & burst_addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
          } else {
            // INCR
            (addr[11:0] & addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
            // Make sure that the max address does not cross addr_width.
            // Use aligned address
            ((addr >> burst_size) << burst_size) + addr_range - 1 <= max_possible_addr;
          }
        } 


        
        // Resetting all the bits greater than data width to 0

        /*foreach (wstrb[index]) {
          if (index < burst_length) {
            wstrb[index] == wstrb[index] & ((1 << port_cfg.data_width/8)-1);
          } 
        }
        */


        addr_valid_delay inside {[0:`SVT_AXI_MAX_ADDR_VALID_DELAY]};
        

        foreach (wvalid_delay[index]) {
          wvalid_delay[index] inside {[0:`SVT_AXI_MAX_WVALID_DELAY]};
        }
        foreach (rready_delay[index]) {
          rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
        }
        foreach (idle_rready_delay[index]) {
          idle_rready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY]};
        }

        /*if (reference_event_for_rready_delay == MANUAL_RREADY) {
          foreach (rready_delay[index]) {
            (index == 0) -> rready_delay[index] inside {[-`SVT_AXI_MAX_RREADY_DELAY : `SVT_AXI_MAX_RREADY_DELAY]};
            (index > 0)  -> rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        } else {
          foreach (rready_delay[index]) {
            rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        }
        */

        bready_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        foreach (idle_bready_delay[index]) {
          idle_bready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY]};
        }


        // Data Before Addr Constraints
        if(data_before_addr) {
          reference_event_for_first_wvalid_delay == PREV_WRITE_DATA_HANDSHAKE;
          reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR,FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR};
        }

        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) {

          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) 

      // For EXCLUSIVE access, the address must be aligned to 
      // the total number of bytes transferred
      if (atomic_type == EXCLUSIVE) {
        (burst_length << burst_size) inside {1,2,4,8,16,32,64,128};

        if (burst_length << burst_size == 2) {
          addr[0] == 1'b0;
        } 
        else if (burst_length << burst_size == 4) {
          addr[1:0] == 2'b0;
        } 
        else if (burst_length << burst_size == 8) {
          addr[2:0] == 3'b0;
        } 
        else if (burst_length << burst_size == 16) {
          addr[3:0] == 4'b0;
        } 
        else if (burst_length << burst_size == 32) {
          addr[4:0] == 5'b0;
        } 
        else if (burst_length << burst_size == 64) {
          addr[5:0] == 6'b0;
        } 
        else if (burst_length << burst_size == 128) {
          addr[6:0] == 7'b0;
        } 
      }

      /* 
       * AXI3 :
       * 1) Burst Size must not exceed the data width
       * 2) Burst Length for WRAP is inside 2,4,8,16
       * 3) Total No. of bytes to be transferred in an exclusive access burst must be a
       *   power of 2.  Max is 128  - Section 6.2.4
       * 4) Burst Length For Idle transactions must be from 1 to Max Idles
       * 5)
      */   

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration :: AXI3) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration :: AXI3) {
`endif
 
        xact_type != COHERENT;
        burst_size <= log_base_2_data_width_in_bytes;

        if (xact_type == IDLE) {
          burst_length inside {[1:`SVT_AXI_MAX_TRANSACTION_IDLE_CYCLES]}; 
        } else {
          if (burst_type == WRAP) {
`ifdef SVT_ACE5_ENABLE
           if(xact_type == ATOMIC && atomic_transaction_type == COMPARE){
              burst_length inside {1,2,4,8,16,32};}
           else {
              burst_length inside {2,4,8,16};}
`else
             burst_length inside {2,4,8,16};
`endif
          } else {
            burst_length inside {[1:`SVT_AXI3_MAX_BURST_LENGTH]};
          }
        }

        // WA(bit 3) bit must not be high if C bit(bit 1) is low
        (cache_type[1] == 0) -> (cache_type[3] == 0);
        // Reserved values:
        cache_type != 4'b0100;
        cache_type != 4'b0101;
        cache_type != 4'b1000;
        cache_type != 4'b1001;
        cache_type != 4'b1100;
        cache_type != 4'b1101;
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      foreach(data_user[i])
       data_user[i] <= ((1 << `SVT_AXI_MAX_DATA_USER_WIDTH) - 1);
`else
      foreach(data_user[i])
       data_user[i] <= ((1 << port_cfg.data_user_width) - 1);
`endif
   }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT

`ifdef SVT_ACE5_ENABLE    
   if(port_cfg.atomic_transactions_enable ==1){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
      if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
         atomic_read_data.size() <= burst_length;
         atomic_read_poison.size() <= burst_length;
         atomic_read_data_user.size() <= burst_length;
       }
       if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
         if(burst_length > 1){
           atomic_read_data.size() == burst_length/2;
           atomic_read_poison.size() == burst_length/2;
           atomic_read_data_user.size() == burst_length/2;
         }
         else {
           atomic_read_data.size() == 1;
           atomic_read_poison.size() == 1;
           atomic_read_data_user.size() == 1;
         }
        }
      }
   else {
     atomic_read_data.size() ==0;
     atomic_read_data_user.size() ==0;
     atomic_read_poison.size() ==0;
//     atomic_resultant_data.size() ==0;
//     atomic_swap_data.size() ==0;
//     atomic_compare_data.size() ==0;
    }
`endif
      if (port_cfg.enable_delayed_response_port) {
        // Transaction supplied through delayed response port.
        // data.size() can be <= burst_length since data is provided
        // through multiple transactions.
        if (is_delayed_response_xact) {
          if (`SVT_AXI_COHERENT_READ_1_BEAT) {
           if(port_cfg.poison_enable ==1){
            poison.size() == 1;}
            data.size() == 1;
            rresp.size() == 1;
          } else if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
          if(port_cfg.poison_enable ==1){
            poison.size() <= burst_length;}
            data.size() <= burst_length;
            rresp.size() <= burst_length;
            data.size() == rresp.size();
          if(port_cfg.poison_enable ==1){
           poison.size() == rresp.size();}
          }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC ) {
        rresp.size() == burst_length;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;  }
      else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC ) {
        if(burst_length > 1){
        rresp.size() == burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length/2;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length/2;
        atomic_read_data_user.size() <= burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        }
        else {
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;}
       }
`endif  
       else {
            rresp.size() == 0;
          }  
        // Transaction supplied through seq_item_port but when
        // configured with enable_delayed_response_port. This corresponds
        // to the transaction handle that is returned in 0-time to the driver.
        } else {
          if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
             data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
             rresp.size() == 0;
          // WRITES
          }
       else {
            rresp.size() == 0;
          }
        }
      } else 
`endif
      {
        if (xact_type == DATA_STREAM) {
          data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
        } else if (`SVT_AXI_COHERENT_READ_1_BEAT) {
          data.size() == 1;
         if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
          rresp.size() == 1;
          data_user.size() == 1;
        } else if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          data.size() == burst_length;
          if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
          rresp.size() == burst_length;
          data_user.size() == burst_length;
        // WRITES. rresp_size should be 0.
        }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
        if(burst_length >1){
        rresp.size() == burst_length/2;
        atomic_read_data.size() == burst_length/2;
        atomic_read_poison.size() == burst_length/2;
        atomic_read_data_user.size() == burst_length/2;
        }
       else {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       }
       else if(xact_type == ATOMIC && !(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         rresp.size() ==0;
         atomic_read_data.size()==0;
         atomic_read_data_user.size()==0;
         atomic_read_poison.size()==0;
      }
`endif  
        else {
          data_user.size() == burst_length;
          data.size() == burst_length;
          rresp.size() == 0;
        }
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) { 
          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } 

      addr_ready_delay inside {[0:`SVT_AXI_MAX_ADDR_DELAY]};

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      resp_user <= ((1 << `SVT_AXI_MAX_BRESP_USER_WIDTH) - 1);
`else
      resp_user <= ((1 << port_cfg.resp_user_width) - 1);
`endif


    // wready_delay[0] can take positive and negative values.
`ifdef INCA
      if ((slave_xact_type != COHERENT) && (slave_xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`else
      if ((xact_type != COHERENT) && (xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`endif
      if (port_cfg.toggle_ready_signals_during_idle_period)
        idle_addr_ready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY_ARR_SIZE]}; 
      else
        idle_addr_ready_delay.size() == 0;
      if (xact_type == WRITE 
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif           
         || xact_type == COHERENT && 
          (coherent_xact_type == WRITENOSNOOP ||
           coherent_xact_type == WRITELINEUNIQUE ||
           coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
           coherent_xact_type == WRITEBACK   ||
           coherent_xact_type == WRITECLEAN  ||
           coherent_xact_type == WRITEEVICT
          )
         ) {
        if (port_cfg.toggle_ready_signals_during_idle_period)
          idle_wready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY_ARR_SIZE]}; 
        else
          idle_wready_delay.size() == 0;
      } else {
        idle_wready_delay.size() == 0;
      }
      if (xact_type != DATA_STREAM) {
       if(!port_cfg.axi_slv_channel_buffers_enable)
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};

        if (reference_event_for_wready_delay == MANUAL_WREADY) {
          foreach (wready_delay[idx]) {
            (idx == 0) -> wready_delay[idx] inside {[-`SVT_AXI_MAX_WREADY_DELAY:`SVT_AXI_MAX_WREADY_DELAY]};
            (idx > 0) -> wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          }
        } else {
          foreach (wready_delay[idx])
            wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          foreach (idle_wready_delay[idx])
            idle_wready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY]};
          foreach (idle_addr_ready_delay[idx])
            idle_addr_ready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY]};
        }
       if(!port_cfg.axi_slv_channel_buffers_enable)
        bvalid_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        if (xact_type == WRITE  
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif      
         ||   xact_type == COHERENT && 
             (coherent_xact_type == WRITENOSNOOP ||
             coherent_xact_type == WRITELINEUNIQUE ||
             coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
             coherent_xact_type == WRITEBACK   ||
             coherent_xact_type == WRITECLEAN  ||
             coherent_xact_type == WRITEEVICT  ||
             coherent_xact_type == EVICT
            )
           ) {
        // The reordering priority of write responses be within
        // 1 to port_cfg.write_resp_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.write_resp_reordering_depth]};
`endif
        }
        else { //if (xact_type == READ) 
        // The reordering priority of read transactions should be within
        // 1 to port_cfg.read_data_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.read_data_reordering_depth]};
`endif
        }

        // An EXOKAY response makes sense only for an EXLUSIVE type
        // atomic access.
        if (atomic_type != EXCLUSIVE) { 
          foreach (rresp[idx])
            (rresp[idx] != EXOKAY); 
          bresp != EXOKAY; 
        }

        if (
            (xact_type == COHERENT) && 
            ( 
              (coherent_xact_type == CLEANUNIQUE) || 
              (coherent_xact_type == MAKEUNIQUE) || 
              (coherent_xact_type == CLEANSHARED) || 
              (coherent_xact_type == CLEANSHAREDPERSIST) || 
              (coherent_xact_type == CLEANINVALID) || 
              (coherent_xact_type == MAKEINVALID) 
            ) 
           ) {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : 1]};
          }
        } else {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : burst_length]};
          }
        }
      }
    } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) 
`endif //SVT_AXI_SVC_USE_MODEL
  } // axi3_4_valid_ranges 

 
  constraint disable_constraint_first_wvalid_reference_event {
    reference_event_for_first_wvalid_delay dist { WRITE_ADDR_VALID:=50000, WRITE_ADDR_HANDSHAKE:=1, PREV_WRITE_DATA_HANDSHAKE:=50000 };
  }

 constraint valid_poison {
    if(port_cfg.poison_enable == 0){
       poison.size()==0;
    }
   }


`ifdef INCA 
   constraint validpoison {
     if(port_cfg.poison_enable==1 && port_cfg.ace_version==svt_axi_port_configuration::ACE_VERSION_2_0){
        poison.size()==1;
     }
     else {
       poison.size()==0;
     }
    }
`endif

`ifdef SVT_ACE5_ENABLE
    constraint valid_archunken{
	        if(port_cfg.rdata_chunking_enable == 1 && xact_type == READ){
		        if(burst_size >= BURST_SIZE_128BIT){
			        archunken inside {0,1};
                  }
		        else {
			        archunken == 0;
                }
            }
	        else {	
		        archunken == 0;
            }
        }

    constraint reasonable_ranges_while_chunking {
      solve chunk_length before rchunkstrb;
      solve chunk_length before rchunknum;
        if(archunken){
            rchunkstrb.size() == chunk_length;
            rchunknum.size() == chunk_length;
        }
        else {
            rchunkstrb.size() == 0;
            rchunknum.size() == 0;
        }
    }

    constraint reasonable_chunk_len{
      solve burst_length before chunk_length;
      solve burst_size before chunk_length;
      if(archunken){
        if(burst_size < BURST_SIZE_128BIT){
          chunk_length == 0;
        }
        else {
          chunk_length inside {[burst_length:(burst_length<<(burst_size - 4))]};
        }
      }
      else {
        chunk_length == 0;
      }
    }
`endif
 /*Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios
 reference_event_for_addr_delay must not be set to FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
 potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
 before driving wready signal.
 */
 constraint reasonable_reference_event_for_addr_delay {
   if(data_before_addr){
   reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR};}
 }
    
`ifdef SVT_AXI_SVC_USE_MODEL
  // **************************************************************************
  //       Reasonable  Constraints
  // **************************************************************************

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Dus5RvTty9UOpNvWOhl+zv9XsCWfifu70kpx1f2d8TJS+0uVcKyDUI+iju2Bz8Qp
7M+k1uSohMbpojCS99g4VDS6id2zh2c8VuPCtvmjhP+gc90MiF83FmiQ6tY39Chj
0djEq2fIdY4aevcEBeYe1IZ4vmnHGGvtk8AgfyvOfwfdP4JTe7NAzQ==
//pragma protect end_key_block
//pragma protect digest_block
p/WSIHQh1dyXU99rgv5GL+DAjAk=
//pragma protect end_digest_block
//pragma protect data_block
RBKNN9TLGXMagOLUelXY57skvGhrQzycmeYebLBYDS/LdSwy6vVYOqrevYN9RnCg
qyzopVD3CY0swApYrNizdBH5H22+ia6TcT9upOTz1RBh4/1TiQLjsL7eNQNdG8M1
n+x85OF4QcysKR3nYBSmRZE+q8Lq9laBKFgUhRGxzfY9vz/s4VFshoEIMGXVMDen
aUGgZxfJEgUycVdVgD5R6IrDC/XxNlEaS3bn6Kufqdv7U5aDb4IQ8igON9jbxE1O
nFmuhBABjOX1C/YVvLuw8Q5XODa6cIrG5rWk/pmKsJyisNhXdwDWRUAtztdOupA9
qKfymN5ZVzhR6Pgonty+K/Oc98QIcvjImxgF7noTReViGumP4W0ExgGfWdBwR9Nt
M49xQV91d42EsAurs45CVk4kaEK4fUQ3lwLRZjGj7U/7ebeyU87EvbnErmG6mNBe
RhdDanyW+2zslYx8PGMg8bjxuDuxa7qMqcPhBr+zjcEROMo6bbnafPkcaCYlWZIG
rVdHrHitPzufr1mmdyLhWvnMuZcv9X8Di7t47pjIasvWkJJi2g4xTmFSPBJR6puW
Cx8KVAYDD8iFDUk0voZQXg==
//pragma protect end_data_block
//pragma protect digest_block
CwYQdZDZsYNGxngSuFkxFOVdnIE=
//pragma protect end_digest_block
//pragma protect end_protected
  constraint reasonable_burst_length {
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI3_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI3_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI3_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4 ||
        `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI4_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI4_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI4_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI_ACE) {
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2:4] :/ SHORT_BURST_wt,
        [5:16] :/ LONG_BURST_wt
      };
    }
  }

  /*
    Reasonable constraint for cache type.
    For exclusive accesses transactions , transactions must not be cached
  */
  constraint reasonable_cache_type
  {
    solve atomic_type before cache_type;
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {   
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE,
                             `SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY,
                             `SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC,
                             `SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC};
        }
      } 
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4) {
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE};
        }
      } 
  }

  /* 
    Reasonable constraint for interleave_pattern
    1) Set the interleave pattern to RANDOM BLOCK for the user to set interleave
    patterns
  */  

  constraint reasonable_interleave_pattern {
    interleave_pattern == RANDOM_BLOCK;
  }

  /* 
    Reasonable constraint for equal block length
    1) Constrain the equal block length to range of 1 to burst_length/2
  */
  
  constraint reasonable_equal_block_length {
    solve interleave_pattern before equal_block_length;
    solve burst_length before equal_block_length;
    if (interleave_pattern ==  EQUAL_BLOCK) {
      if (burst_length > 1) {
        equal_block_length  inside {[1 : (burst_length >> 1)]};
      }
      else {
        equal_block_length == 1;
      }
    }
  }

  constraint reasonable_addr_valid_delay {
   addr_valid_delay dist {
     0 := ZERO_DELAY_wt, 
     [1:(`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
     [((`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_VALID_DELAY] :/ LONG_DELAY_wt
   };
  }


  constraint reasonable_wakeup_assert_deassert_delay {
    awakeup_assert_delay >= `SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY;
    awakeup_assert_delay <  `SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY;
    awakeup_deassert_delay >= `SVT_AXI_MIN_AWAKEUP_DEASSERT_DELAY;
    awakeup_deassert_delay <  `SVT_AXI_MAX_AWAKEUP_DEASSERT_DELAY;
  }

  constraint reasonable_rready_delay {
    /*foreach (rready_delay[idx]) {
      if (reference_event_for_rready_delay == MANUAL_RREADY && idx == 0) {
        rready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_RREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_RREADY_DELAY: -((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {
          rready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] := SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] := LONG_DELAY_wt >> 1
          };
      }
    }
    */
    foreach (rready_delay[idx]) {
      rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  constraint reasonable_idle_rready_delay {
    foreach (idle_rready_delay[idx]) {
      idle_rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  
  // Enforces a distribution based on the weights.
  constraint reasonable_wvalid_delay {
    foreach (wvalid_delay[idx]) {
      wvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_WVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WVALID_DELAY >> 2)+1):`SVT_AXI_MAX_WVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }


  // Enforces a distribution based on the weights.
  constraint reasonable_bready_delay {
    bready_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  constraint reasonable_idle_bready_delay {
    foreach (idle_bready_delay[i]) 
      idle_bready_delay[i] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)+1):`SVT_AXI_MAX_IDLE_BREADY_DELAY] :/ LONG_DELAY_wt
    };
  }


  constraint reasonable_tready_delay {
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
      tready_delay.size() == `SVT_AXI_MAX_STREAM_BURST_LENGTH;
      foreach (tready_delay[idx]) {
        tready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_TREADY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_TREADY_DELAY >> 2)+1):`SVT_AXI_MAX_TREADY_DELAY] :/ LONG_DELAY_wt
       };
      }
    } else {
      tready_delay.size() == 0;
    }
  }

  /** 
   * This constraint insures that unimplemented features are avoided during randomization.
   */
  constraint exclude_master_unimplemented_features
  {
    xact_type != IDLE;
    interleave_pattern != EQUAL_BLOCK;
    start_new_interleave == 0;
    reference_event_for_rready_delay != MANUAL_RREADY;
  }

  //--------------------------------------------------------------------------------------
  /**************************** SLAVE CONSTRAINTS ******************************** */
  constraint reasonable_data {
    if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
      if (
           (xact_type == READ) || 
           (
             (xact_type == COHERENT) &&
             (
               coherent_xact_type == READNOSNOOP                     ||
               coherent_xact_type == READONCE                        ||
               coherent_xact_type == READONCECLEANINVALID                        ||
               coherent_xact_type == READONCEMAKEINVALID                        ||
               coherent_xact_type == READSHARED                      ||
               coherent_xact_type == READCLEAN                       ||
               coherent_xact_type == READNOTSHAREDDIRTY              ||
               coherent_xact_type == READUNIQUE          
             )
           )
         ) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
         data.size() == burst_length;
         if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
`else
       if (!port_cfg.enable_delayed_response_port) {
           if(port_cfg.poison_enable ==1){
             poison.size() == burst_length;}
           data.size() == burst_length;
       }
`endif
       data_user.size() == burst_length;
        foreach (data[index]) {
             data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        }
      }
      // No data associated with these transactions 
      if(`SVT_AXI_COHERENT_READ_1_BEAT) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
        data.size() == 1;
`else
       if (!port_cfg.enable_delayed_response_port) {
          if(port_cfg.poison_enable ==1){
             poison.size() == 1;}
          data.size() == 1;
       }
`endif
       data_user.size() == 1;
        foreach (data[index]) {
             data[index] <= 0;
        }
      if(port_cfg.poison_enable ==1){
            foreach (poison[index]) {
             poison[index] <= 0;}
          }
      }
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_wready_delay {
    foreach (wready_delay[idx]) {
      // MANUAL_READY not supported.
      /*if (reference_event_for_wready_delay == MANUAL_WREADY && idx == 0) {
        wready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_WREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_WREADY_DELAY: -((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {*/ 
        wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt
          };
        //}
      }
    }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_wready_delay {
    foreach (idle_wready_delay[idx]) {
        idle_wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_WREADY_DELAY] :/ LONG_DELAY_wt
          };
    }
  }
 

  // Enforces a distribution based on the weights.
  constraint reasonable_rvalid_delay {
    foreach (rvalid_delay[idx]) {
      rvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_RVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_RVALID_DELAY >> 2)+1):`SVT_AXI_MAX_RVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_addr_ready_delay {
    addr_ready_delay dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_ADDR_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_ADDR_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_DELAY] :/ LONG_DELAY_wt
    };
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_addr_ready_delay {
    foreach (idle_addr_ready_delay[idx]) {
      idle_addr_ready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_bvalid_delay {
    bvalid_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  /**
   * Reasonable constraint for random_interleave_array
   * Constraint the random interleave array from 1 to burstlength
   * If the  array values exceed the burst length, those values will be ignored
   */

   constraint reasonable_random_interleave_array {
     if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
       if(`SVT_AXI_COHERENT_READ_1_BEAT) 
         random_interleave_array.size() == 1;
       else
         random_interleave_array.size() == burst_length;

       foreach (random_interleave_array[index]) {
         random_interleave_array[index] inside {[1 : burst_length]};
       }
     } else {
       random_interleave_array.size() == stream_burst_length;
     }
   }

    constraint exclude_slave_unimplemented_features
    {
      interleave_pattern != EQUAL_BLOCK;
      start_new_interleave == 0;
      reference_event_for_wready_delay != MANUAL_WREADY;
    }

`endif

`ifdef SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, "test_constraintsX" constraints are not enabled in svt_axi_transaction. A
   * test can enable them by defining the following macro during the compile:
   *   SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif

//reasonable  soft constraint for cust_xact_flow == 0. To support default behavior of cust_xact_flow disabled and overridden by user to enable it automatically whenever inline randomization constraint is added
constraint reasonable_cust_xact_flow {
  soft cust_xact_flow == 0;
} 

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`else
`svt_vmm_data_new(`SVT_TRANSACTION_TYPE)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /** returns 1 if status of all relevant phases of current transaction are assigned as ABORTED */
  extern virtual function bit is_aborted(int mode = 0);

  /** returns 1 if current transaction is configured as secure access */
  extern virtual function bit is_secure(bit allow_secure = 1);

  /** Returns 1 if current transaction is of device_type */
  extern virtual function bit is_device_type();

  /** Returns 1 if current transaction is DVM transaction */
  extern virtual function bit is_dvm_xact();

  /** Returns 1 if current transaction is cacheable transaction */
  extern virtual function bit is_cacheable_xact();

  /** Returns 1 if current transaction is allocate transaction */
  extern virtual function bit is_allocate_xact();

  /** Determines if this transaction is a CMO transaction */
  extern function bit is_cmo_xact();


//  /** Returns 1 if current transaction is of device_type or DVM transaction 
//   * Additinally this function will fire an error if device type or DVM transactions 
//   * are issued from not allowed ports 
//   */
//  extern virtual function bit skip_port_interleaving();

  /** waits for transaction to end */
  extern virtual task wait_for_transaction_end();


 /** waits for slave transaction to update the memory*/
  extern virtual task wait_for_write_transaction_to_update_memory();

  /** returns 1 if transaction status shows ended otherwise 0 */
  extern virtual function bit is_transaction_ended();

  /** waits for addr phase to end */
  extern virtual task wait_for_addr_phase_ended ();
  
  /** waits for data phase to end */
  extern virtual task wait_for_data_phase_ended();
  
  /** waits for write resp phase to end */
  extern virtual task wait_for_write_resp_phase_ended();

  /** mark end of transaction */
  extern virtual function void set_end_of_transaction(bit aborted=0);
  

   /**
  * Returns 1 if the specified error_kind is there in transaction, else returns 0 
  */
  extern virtual function bit has_axi_exception(int error_kind); 
  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************

  `svt_data_member_begin(svt_axi_transaction)
    `svt_field_object(port_cfg,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK| `SVT_REFERENCE, `SVT_HOW_REF)
    `ifndef INCA
    `svt_field_object      (exception_list,                             `SVT_ALL_ON|`SVT_DEEP|`SVT_NOCOMPARE|`SVT_UVM_NOPACK,  `SVT_HOW_DEEP)
    `endif
    `svt_field_object(associated_barrier_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`ifdef SVT_UVM_TECHNOLOGY
    `svt_field_object(causal_gp_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`endif

  // ****************************************************************************

  `svt_data_member_end(svt_axi_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
 //----------------------------------------------------------------------------
  /**
   * Calculates whether the transaction is partial or full cacheline access.
   * returns 1, if transaction is full cacheline access. returns 0, if it is a 
   * partial cacheline access.
   * 
   * @param cacheline_size indicates the value of the master cache line size
   */
  extern virtual function bit is_full_cacheline(int cacheline_size);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
  extern virtual function svt_pattern do_allocate_pattern ();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern allocate_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when a full tranaction is to be recorded.  Note that not all
   * properties are written.  Instead, only properties needed for debug are added.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_full_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is RADDR, RDATA, WADDR, WDATA, or WRESP.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_filtered_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is "STREAM DATA".
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_stream_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the pa_format_type is set to FSDB_PERF_ANALYSIS.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_perf_analysis_xml_pattern();

  // ----------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
   extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

//-----------------------------------------------------------------------------------
/**
  * This method is used to set object_type for bus_activity when
  * bus_activity is getting started on the bus .
  * This method is used by pa writer class in generating XML/FSDB 
  */
  extern function void  set_pa_data(string typ = "" ,string channel  ="");
 
//-----------------------------------------------------------------------------------
  /**
  * This method is used to  delate  object_type for bus_activity when bus _activity 
  * ends on the bus .
  * This methid is used by pa writer class  in generating XML/FSDB 
  */
  extern function void clear_pa_data();
  
//------------------------------------------------------------------------------------
  /** This method is used in setting the unique identification id for the
  * objects of bus activity
  * This method returns  a  string which holds uid of bus activity object
  * This is used by pa writer class in generating XML/FSDB
  */
  extern virtual function string get_uid();

//------------------------------------------------------------------------------------
  /** Sets the configuration property */ 
  extern function void set_cfg(svt_axi_port_configuration cfg);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

`ifdef SVT_ACE5_ENABLE  
  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_write_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_read_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);
`endif
  /** 
    * Populates the partial data and byteen provided into data and byteen
    * that is used to write into a full cacheline
    */
  extern function void populate_partial_data_and_byteen (
                                                         input bit[7:0] data[],
                                                         input bit byteen[],
                                                         output bit[7:0] cache_data[],
                                                         output bit cache_byteen[]
      );

  /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane_for_data_user(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`ifdef SVT_ACE5_ENABLE
 /** Returns the address and lanes corresponding to the beat number for atomic compare read data*/
  extern function void get_beat_addr_and_lane_atomic_read_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number for atomic compare write data*/
  extern function void get_beat_addr_and_lane_atomic_write_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`endif

  /** Gets the beat number corresponding to an address */
  extern function int get_beat_num_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr, 
                                                          bit use_tagged_addr = 0
                                          );

  /**
   * Returns a string (with no line feeds) that reports the essential contents
   * of the packet generally necessary to uniquely identify that packet.
   *
   * @param prefix (Optional: default = "") The string given in this argument
   * becomes the first item listed in the value returned. It is intended to be
   * used to identify the transactor (or other source) that requested this string.
   * This argument should be limited to 8 characters or less (to accommodate the
   * fixed column widths in the returned string). If more than 8 characters are
   * supplied, only the first 8 characters are used.
   * @param hdr_only (Optional: default = 0) If this argument is supplied, and
   * is '1', the function returns a 3-line table header string, which indicates
   * which packet data appears in the subsequent columns. If this argument is
   * '1', the <b>prefix</b> argument becomes the column label for the first header
   * column (still subject to the 8 character limit).
   */
`ifdef SVT_UVM_ENABLE_FGP
  (* uvm_fgp_lock = "psdisplay_short" *)
`endif
  extern virtual function string psdisplay_short( string prefix = "", bit hdr_only = 0);

  /** 
    * Limits the data to what can be transmitted if the address is
    * unaligned. If the address is unaligned, we need to take care 
    * that data[0] and wstrb[0] are consistent with what can actually 
    * be driven on the bus. 
    * For example, for a 64 bit bus, if the address is 0x7,
    * data can be sent only on 1 byte for the first beat.
    * For a FIXED burst the address is same for all beats, so this
    * operation needs to be done for all beats. For other bursts, only
    * the first address can be unaligned, other beats are aligned
    * addresses
    * @param data_only(Optional: default = 0) If this bit is set the 
    * operation is done only for data. 
    * @param beat_num(Optional: default = -1) Applicable for a FIXED burst.
    * When set to -1, masking is done for all beats, otherwise it is 
    * done only for the selected beat. 
    */
  extern function void mask_data_for_unaligned_addr(bit data_only = 0,int beat_num = -1);
  
  /**
    * Ensures that valid x,z,0,1 all four state datas are calculated with
    * respect to data_mask values. 
    * This function is called under SVT_MEM_LOGIC_DATA macro define only,
    * to make sure while masking valid x and z state data also considered
    * towards masked data.
    */ 
  extern function logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] mask_data_for_x_z_values (logic [`SVT_AXI_MAX_DATA_WIDTH -1:0] data, bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data_mask);
  
  /**
    * Ensures that only valid lanes have wstrb asserted. In wysisyg format
    * the constraints leave data[] and wstrb[] open. This function is called in
    * post_randomize to make sure that wstrb is asserted only for valid lanes
    */ 
  extern function void get_wstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

`ifdef SVT_ACE5_ENABLE
    /**
    * Ensures that only valid lanes have tag_update asserted. In wysisyg format
    * the constraints leave tag[] and tag_update[] open. This function is called in
    * post_randomize to make sure that tag_update is asserted only for valid lanes
    */ 
  extern function void get_tag_update_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Returns the tag_update in the tag_update_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the tag_update is returned such that packed_tag_update[0] 
    * corresponds to the tag_update for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in tag_update_to_pack[] is directly
    * packed to packed_tag_update[]. 
    * @param tag_update_to_pack tag_update to be packed
    * @param packed_tag_update[] Output byte stream with packed tag_update
    */
  extern function void pack_tag_update_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update_to_pack[],
                                          output bit packed_tag_update[]
                                        ); 

  /**
    * Returns the tag in the tag_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either tag[] or cache_write_tag[]
    * fields of this class have been passed as arguments to tag_to_pack[] field.
    * In the case of WRAP bursts the tag is returned such that packed_tag[0] 
    * corresponds to the tag for the wrap boundary. 
    * In the case of INCR bursts, the tag as passed in tag_to_pack[] is directly
    * packed to packed_tag[]. 
    * @param tag_to_pack tag to be packed
    * @param packed_tag[] Output byte stream with packed tag
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_tag_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output logic[3:0] packed_tag[]
                                        ); 
`else
  extern function void pack_tag_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output bit[3:0] packed_tag[]
                                        );
`endif 
 
 
  /** Converts tag from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_right_justified_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from wysiwyg format to right justified format */
  extern function void convert_tag_update_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);


  /** Converts tag from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from right justified format to wysiwyg format */
  extern function void convert_tag_update_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Ensures that only valid lanes have chunkstrb asserted. In wysisyg format
    * the constraints leave data[] and rchunkstrb[] open. This function is called in
    * post_randomize to make sure that chunkstrb is asserted only for valid lanes
    */ 
  extern function void get_chunkstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1:0] rchunkstrb[]);

`endif

 /**
    * Ensures that only valid lanes have poison asserted. In wysisyg format
    * the constraints leave data[] and poison[] open. This function is called in
    * post_randomize to make sure that poison[] is asserted only for valid lanes
    */ 
  extern function void get_poison_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

 /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);


  /**
    * Returns the encoding for AWSNOOP/ARSNOOP/ACSNOOP based on the 
    * transaction type
    * @return The encoded value of AWSNOOP/ARSNOOP/ACSNOOP
    */
  extern function bit[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] get_encoded_snoop_val();

`ifdef SVT_ACE5_ENABLE
 
  /**
    * Returns the encoding for AWCMO based on the 
    * cmo_on_write_xact_type type
    * @return The encoded value of AWCMO
    */
  extern function bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] get_encoded_awcmo_val();

   /**
    * Decodes the given AWCMO value and returns the transaction type.
    * @param awcmo_val The value on AWCMO
    */
  extern function cmo_on_write_xact_type_enum get_decoded_awcmo_val(bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] awcmo_val);

  /**
   * Sets Combined Write and CMO type
   */
  extern function void set_combined_writecmo_transaction_type();
  
  /**
   * Indicates whether the current transaction is write cmo or not
   */
  extern function bit is_combined_writecmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_pcmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_non_pcmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl or writeuniquefull cmo or not
   */
  extern function bit is_combined_writeunique_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnp* cmo or not
   */
  extern function bit is_combined_writenosnp_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniquefull cmo or not
   */
  extern function bit is_combined_writeuniquefull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpfull cmo or not
   */
  extern function bit is_combined_writenosnpfull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl cmo or not
   */
  extern function bit is_combined_writeuniqueptl_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpptl cmo or not
   */
  extern function bit is_combined_writenosnpptl_cmo_xact();  

`endif

  /**
    * Decodes the given snoop value(ARSNOOP/ACSNOOP) and returns the transaction type.
    * This function can be used for the read address channel and the
    * snoop address channel. 
    * @param snoop_val The value on ARSNOOP/ACSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_read_snoop_val(bit[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Decodes the given snoop value(AWSNOOP) and returns the transaction type.
    * This function can be used for the write address channel. 
    * @param snoop_val The value on AWSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_write_snoop_val(bit[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Returns the channel on which a transaction will be transmitted
    * @return The channel (READ/WRITE) on which this transaction will
    * be transmitted.
    */
  extern function xact_type_enum get_transmitted_channel();
  /**
    * Indicates if this transaction is applicable for updates in
    * the FIFO rate control model 
    * @return Returns 1 if applicable, else returns 0 
    */
  extern function bit is_appplicable_for_fifo_rate_control();

  /**
    * Checks if the coherent transaction is DVM Sync 
    */
  extern function bit is_coherent_dvm_sync();
 
  /**
    * Returns the index (of data or wstrb fields) corresponding 
    * to the wrap boundary
    */ 
  extern function int get_wrap_boundary_idx();

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the index (of atomic_read_data) corresponding 
    * to the wrap boundary for Atomic compare transaction
    */ 
  extern function int get_wrap_boundary_idx_for_atomic_compare_read_data();

`endif

  /** returns lowest address of the transaction. For WRAP type of transaction
    * it indicates starting address after transaction statisfies WRAP condition
    * and wraps over to include lower addresses
    */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_wrap_boundary();

  /** returns burst size aligned address */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_burst_boundary();

  /**
    * Returns the byte lanes on which data is driven for a given data width
    */
  extern function void get_byte_lanes_for_data_width(
                bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                int beat_num,
                int data_width_in_bytes,
                output int lower_byte_lane,
                output int upper_byte_lane
          );
  
  /**
    * Checks if the transaction crosses the 4kb boundary
    */
  extern function bit is_addr_4kb_boundary_cross();

  /**
    * Returns the data in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either data[] or cache_write_data[]
    * fields of this class have been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the data in the atomic_compare_read_data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that atomic_read_data[]
    * field of this class have been passed as arguments to atomic_compare_read_data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_atomic_compare_read_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in atomic_compare_read_data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param atomic_compare_read_data_to_pack Data to be packed
    * @param packed_atomic_compare_read_data[] Output byte stream with packed data
    */

`ifdef SVT_MEM_LOGIC_DATA
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output logic[7:0] packed_atomic_compare_read_data_data[]
                                                             ); 
`else  
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output bit[7:0] packed_atomic_compare_read_data[]
                                                             ); 
`endif 

`endif 
  /**
    * Returns the data_user in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that data_user[] 
    * has been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data_user is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data_user as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_user_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_user_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

  /**
    * Returns the wstrb in the wstrb_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the wstrb is returned such that packed_wstrb[0] 
    * corresponds to the wstrb for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in wstrb_to_pack[] is directly
    * packed to packed_wstrb[]. 
    * @param wstrb_to_pack wstrb to be packed
    * @param packed_wstrb[] Output byte stream with packed wstrb
    */
  extern function void pack_wstrb_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb_to_pack[],
                                          output bit packed_wstrb[]
                                        ); 
   /**
    * Returns the poison in the poison_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either poison[] or cache_write_poison[]
    * fields of this class have been passed as arguments to data_to_pack5[] field.
    * In the case of WRAP bursts the data is returned such that packed_poison[0] 
    * corresponds to the poison for the wrap boundary. 
    * In the case of INCR bursts, the poison as passed in poison_to_pack[] is directly
    * packed to packed_poison[]. 
    * @param poison_to_pack poison to be packed
    * @param packed_poison[] Output byte stream with packed poison
    */
  extern function void pack_poison_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison_to_pack[],
                                          output bit packed_poison[]
                                        ); 

  /**
    * Unpacks the data in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data is directly unpacked into unpacked_data
    * For a WRAP burst, the data is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif
  
  /**
    * Unpacks the data_user in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data_user is directly unpacked into unpacked_data
    * For a WRAP burst, the data_user is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data_user starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data_user( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data_user( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif

  /**
    * Unpacks the wstrb in wstrb_to_unpack[] into unpacked_wstrb.
    * For an INCR burst, the wstrb is directly unpacked into unpacked_wstrb
    * For a WRAP burst, the wstrb is unpacked such that unpacked_wstrb[0] corresponds
    * to the starting address. The assumption here is that wstrb_to_unpack[] has
    * a byte stream whose wstrb starts from the address corresponding to the wrap
    * boundary
    * @param wstrb_to_unpack The wstrb to unpack.
    * @param unpacked_wstrb The unpacked wstrb.
    */
  extern function void unpack_byte_stream_to_wstrb( 
                                            input bit wstrb_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] unpacked_wstrb[]
                                          ); 
   /**
    * Unpacks the poison in poison_to_unpack[] into unpacked_poison.
    * For an INCR burst, the poison is directly unpacked into unpacked_poison
    * For a WRAP burst, the poison is unpacked such that unpacked_poison[0] corresponds
    * to the starting address. The assumption here is that poison_to_unpack[] has
    * a byte stream whose poison starts from the address corresponding to the wrap
    * boundary
    * @param poison_to_unpack The poison to unpack.
    * @param unpacked_poison The unpacked poison.
    */
  extern function void unpack_byte_stream_to_poison( 
                                            input bit poison_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] unpacked_poison[]
                                          ); 
                     
  /**
   * Does a basic validation of this transaction object
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);

  /**
    * Sets the suspend_master_xact property
    */
  extern virtual function void suspend_xact();

  /**
    * Unsets the suspend_master_xact property
    */
  extern virtual function void resume_xact();

  /**
    * Gets the number of beats of data/resp to be sent.
    */
  extern function int get_burst_length(int ignore_exceptions = 0);

`ifdef SVT_ACE5_ENABLE
  /**
    * Gets the number of beats for atomic_read_data in Atomic compare transactions 
    */
   extern function int get_burst_length_for_atomic_compare_read_data(int ignore_exceptions =0);
`endif

  /**
    * Gets the burst_type of a transaction.
    */
  extern function burst_type_enum get_burst_type(int ignore_exceptions = 0);

  /**
    * Gets the burst_size of a transaction.
    */
  extern function burst_size_enum get_burst_size(int ignore_exceptions = 0); 

  /**
   * Gets the minimum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_min_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
   * Gets the maximum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Maximum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_max_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
  extern function bit is_address_overlap(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
    * Returns the total number of bytes transferred in this transaction or beat number
    * svt_axi_port_configuration::get_byte_count_from_wstrb_enable set to 0,
    * the byte count is calculated using burst_length and burst_size based on
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * If svt_axi_port_configuration::get_byte_count_from_wstrb_enable
    * is set to 1, the byte count is calculated using wstrb based on 
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * @return The total number of bytes transferred in this transaction or beat number
    */
  extern virtual function int get_byte_count(int beat_num = -1);

  /** @cond PRIVATE */
  /** Converts data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif
`ifdef SVT_ACE5_ENABLE
  /** Converts atomic_read_data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`else
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`endif
`endif
  /** Converts data_user from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstb from wysiwyg format to right justified format */
  extern function void convert_wstrb_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from wysiwyg format to right justified format */
  extern function void convert_poison_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstrb from right justified format to wysiwyg format */
  extern function void convert_wstrb_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from right justified format to wysiwyg format */
  extern function void convert_poison_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Turns-off randomization for all AXI3/AXI4 parameters */
  extern virtual function void set_axi3_4_randmode(bit on_off=0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    * @param disable_msg_info Disables information regarding message format
    * @return The data as a string. If corresponding wstrb is 0, data is marked as 'xx'
    */
  extern virtual function string get_write_data_string(bit[7:0] xact_data[],bit xact_wstrb[],bit disable_msg_info = 0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    */
  extern virtual function string get_read_data_string(bit[7:0] xact_data[]);

  /**
    * Returns the contents of wstrb as a string. 
    * @param  xact_wstrb A bit stream array of the data which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    */
  extern virtual function string get_wstrb_string(bit xact_wstrb[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function. If xact_wstrb is 0,
                   corresponding xact_data is not compared 
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_write_data(bit[7:0] xact_data[],bit xact_wstrb[], bit[7:0] ref_data[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_read_data(bit[7:0] xact_data[],bit[7:0] ref_data[]);

  /**
    * Gets a single response status based on rresp of each beat or bresp.
    * If it is an exclusive access, then this function returns an OKAY response
    * if all beats have a response of EXOKAY, otherwise it returns a SLVERR response
    * For normal transactions, this function returns OKAY only if all beats have
    * a response of OKAY
    * @return Returns the combined response status of all beats 
    */
  extern function resp_type_enum get_response_status();

  /** Returns first data_valid_assertion_time for read channel transaction or write
    * response assertion time for write channel transaction
    */
  extern function real get_response_assertion_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** Returns data_valid_assertion_time for the beat number of given address read channel transaction or write
    * response assertion time for write channel transaction.
    */
  extern function real get_response_assertion_time_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** returns id considering only the bits which are used by exclusive monitor */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1:0] excl_id(bit use_partial_id=1);

  /** returns address considering only the bits which are used by exclusive monitor.
    * However, if num_addr_bits_used_in_exclusive_monitor is set to -1 this indicates that, user wants
    * use specified start and end address ranges for each exclusive monitor. In this case,
    * this method will return exclusive monitor index with tagged address attribute i.e. secured/nonsecure
    * bit, as exclusive monitored address. This models the interconnect's behaviour of monitoring
    * different address chunks.
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] excl_addr(bit use_partial_addr=1, bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr=0);

  /** returns address aligned to cacheline size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline_addr(bit use_tagged_addr=0);

  /** returns address aligned to snoop data width size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_aligned_addr();

  /** returns the status corresponding to the status mode value passed */
  extern function status_enum get_status(int status_mode);

  /** Outputs the expected snoop addresses. 
    * If the transaction does not generate a snoop, the function returns 0, else it returns 1.
    * However, if include_non_snooped_xacts is set, the function includes WRITEBACK, WRITECLEAN,
    * EVICT, WRITEEVICT and cache maintenance transactions sent to NON-SHAREABLE region as well.
    */
  extern function bit get_expected_snoop_addr(output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] expected_snoop_addr[$], input bit use_tagged_addr=0, input bit include_non_snooped_xacts = 0, input int cache_line_size = -1);

  /** Returns 1 if this transaction type generates a snoop, else returns 0 */
  extern function bit has_snoop();

  /** Returns 1 if this transaction is a full cacheline access, else returns 0 */
  extern function bit is_cache_line_access();

  /** Sets the port kind to master or slave */
  extern function void set_port_kind(svt_axi_port_configuration::axi_port_kind_enum axi_port_kind);

  /** Returns address concatenated with tagged attributes which require indipendent address space.
    * for example, if secure access attribute is enabled bye setting num_enabled_tagged_addr_attributes[0] = 1
    * then this bit will be used to provide unique address spaces for secure and non-secure transactions.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Address that needs to be tagged when use_arg_addr is set to '1'
    * @param      use_cacheline_addr Indicates if returned address should be aligned to cache line size
    * @return              Returns address tagged with address attribute of corresponding port
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr = 0, bit use_cacheline_addr=0);

  /** @param  arg_addr Holds Address for which untagged part needs to be obtained
    * @return          Untagged part of Address "arg_addr" will be returned
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Sets transaction attributes from tagged address.
    * for example, if secure access attribute is enabled then security attribute of current transation can be set from the tagged address
    * passed through argument or current transaction address.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Tagged Address from which current transacion attributes need to be set.
    */
 extern task set_tag_from_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Function that sets xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set */
  extern function void set_xact_type();

  /** Function returns xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set xact_type will not be changed for the particular transaction.
    */
  extern function xact_type_enum get_xact_type();

`ifdef SVT_ACE5_ENABLE
  /** Sets the atomic transaction type */
  extern function void set_atomic_transaction_type();

 /**
    * Returns the encoding for AWATOP based on the 
    * transaction type
    * @return The encoded value of AWATOP
    */
  extern function bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] get_encoded_atomicop_val();

 /**
    * Returns the decoding  for AWATOP based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function atomic_xact_op_type_enum get_decoded_atomicop_val(bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] awatop_val);

 /**
    * Returns the decoding  for Endianness based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function endian_enum get_decoded_endianness_val(bit endian_val);

  /** Returns the inbound data size for atomic transaction */
  extern function int get_atomic_transaction_inbound_data_size_in_bytes();
  
  extern function bit is_addr_aligned_to_total_outbound_data();

 /** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] get_masked_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[], bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb[]);
  
/** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function void get_masked_atomic_read_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_read_data[],output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data);

  /** Returns the masked atomicop wstrb and  data based on current atomic xact data_size */
  extern function bit [(`SVT_AXI_WSTRB_WIDTH-1):0] get_masked_wstrb(bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb_);

  /** Performs atomic operation at beat level */
  extern function bit perform_atomic_operation(input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data, 
                                                input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],
                                                input bit [`SVT_AXI_WSTRB_WIDTH-1:0] wstrb[],
                                                output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_resultant_data_
                                                );

 
/** Unpacks data into atomic_swap_data and atomic_compare_data field. This is applicable for ATOMIC_COMPARE transactions only */
   extern function void unpack_data_into_atomic_swap_and_atomic_compare_data(input bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],int beat_num);


 /** Unpacks atomic_resultant_data into beat_format to do the beat formation */
  extern function void unpack_atomic_resultant_data_into_beat_format (input bit[(`SVT_AXI_MAX_DATA_WIDTH -1):0] atomic_resultant_data_);


/** Performs Atomic xact operation such as ADD etc. */
  extern function void perform_atomic_xact_operation(svt_axi_transaction xact);


 /** unpacks wstrb into atomic_swap_wstrb and atomic_compare_wstrb into field. This is applicable for ATOMIC_COMPARE transactions only */
  extern function void unpack_wstrb_into_atomic_swap_and_atomic_compare_wstrb(input bit [(`SVT_AXI_MAX_DATA_WIDTH/8-1):0] wstrb[],int beat_num);

`endif
  /**
    * Indicates if this transaction has poison for any 64-bit chunk 
    * @return Returns 1 if poison is present, else returns 0
    */
  extern function bit has_poison();

  /** Marks current transaction as part of multipart dvm sequence to avoid irrelevant
    * check being performed on this transaction.
    * Since only first transaction of multipart dvm transaction sequence has control information on LSB[15:0] bits,
    * it is important to set this bit to '1', before randomizing the second or later transaction object so that, 
    * second or later part of multipart dvm sequence can ignore dvm address constraints for control fields.
    */
  extern virtual task set_multipart_dvm_flag (string kind = "");

  /** returns first beat of coherent response of current transacton */
  extern virtual function coherent_resp_type_enum get_coh_resp();

  /** returns '1' if current transaction matches expected transaction type i.e. for coherent transaction
    * if it has matched coherent_xact_type and for non_coherent transaction if it matched xact_type, otherwise it returns '0'
    */
  extern virtual function bit is_type_matched(int rw_type = -1, string typ = "non_dvm_non_barrier");

  /** returns '1' if current transaction will allocate a cacheline but, there are at least one transaction currently active
    *             which will attempt to de-allocate the same cacheline.
    * returns '0' otherwise.
    */
  extern virtual function bit has_overlapped_dealloc_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns '1' if overlapped transaction between read and write channel found else '0' */
  extern virtual function bit has_overlapped_rd_wr_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns calculated parity value for 8bit of data */
  extern virtual function bit parity_bit_from_8bit_data(bit [7:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_16bit_data(bit [15:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_1bit_data(bit data, bit even_odd_parity = 1);
  extern virtual function void parity_for_xact_field(input string xact_signal_name = "", input bit even_odd_parity = 1);

  /** returns calculated data check parity value to data */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] calculate_parity(bit [`SVT_AXI_MAX_DATA_WIDTH-1:0] data);

 /** returns converted  data check to pison value */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/64)-1:0]convert_datacheck_to_poison(bit [`SVT_AXI_MAX_DATA_WIDTH/8-1:0] is_datachk_passed,bit [`SVT_AXI_MAX_DATA_WIDTH/64-1:0]data_chk_to_poison);

  /** returns '1' if transaction passed through argument i.e. overlapped_xact is found active while
    * current transaction is found active or in other words both are found active at the same time */
  extern virtual function bit is_overlapped_in_time(svt_axi_transaction overlapped_xact);

  /** returns '1' if current transaction will allocate a cacheline else returns '0' */
  extern virtual function bit is_alloc_xact();

  /** returns '1' if current transaction will de-allocate a cacheline else returns '0' */
  extern virtual function bit is_dealloc_xact();

  /** updates num_xacts_blocked_progress_of_curr_xact with number of xacts that blocked progress of current xact */
  extern virtual task update_num_xacts_blocked_progress_of_curr_xact(int num_blocked_xacts=1, int mode=0);

  /** returns '1' if current transaction is not supposed to return data as part of coherent read response */
  extern virtual function bit is_read_response_without_data(int mode=0);

  /** returns '1' if current transaction will allocate a cacheline in L3 else returns '0' */
  extern virtual function bit is_l3_allocate(bit is_exclusive=0, bit is_partial_data=1);

  /** returns '1' if current transaction will de-allocate a cacheline from L3 else returns '0' */
  extern virtual function bit is_l3_deallocate(bit is_partial_data=1);

  /** returns '1' if current transaction is supposed to update memory with L3 data */
  extern virtual function bit is_l3_update_to_mem(bit is_partial_data=1);

  /** returns '1' if current transaction doesn't cover full cacheline */
  extern virtual function bit is_partial_cacheline_data();

  /** Returns number of byte whose wstrb is '1' */
  extern virtual function int get_valid_byte_count();

  /** returns '1' if current transaction is determined to be valid exclusive type */
  extern virtual function bit is_exclusive_access(string mode="", bit shared=1);

  /** Sets the channel on which a transaction will be transmitted */
  extern function void set_transmitted_channel();

  /** Returns '1' if write strobes are driven correctly otherwise, returns '0' */
  extern virtual function bit check_wstrb(bit silent=0);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_transaction)
`endif
endclass
/**
Transaction Class Macros definition  and utility methods definition
*/

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
spgycq4Zisdzt/+kVzeHcmDaTm4kNmiyVSN0i5oI21Jv4BA3MyjezXs0mRX18CnT
JIdMMJy9UPv519m3NagPD6LTw+mPAg6VtaRUXPdoaW2ch4smIGAPr3CAeh7wGGGa
Lt4TS3M0zDVXPCcrIdxekkxDxSRpX4KvAMz0G0/Snm406zvpD5QSzw==
//pragma protect end_key_block
//pragma protect digest_block
PU8+hCH2odAxBUrhhHJDeLw7BCo=
//pragma protect end_digest_block
//pragma protect data_block
kXQDIvFH3qQty+Kq9Msb4QkAY1VgF/JLkn7/nmCbNZyG0W7HZmLH6mvnUQMWvNyu
hEh3KafMlBIxv/e6+AzSggnqfgn6cCxyet1ImZGeHqrSqW3PkIBgcXftEhQCqf7v
za6SaT63fMgjsauqgnCsa+GMuJhivPd4HJwWYrgZ7KGX9IghcGxTpNPSd9HPd8H6
QTDr5LUIPpENwlmkHXk1M3hEBBmaYS/8rUy48w4YVJKyFK+EiZSHLPC+auHMJp4N
GG5HIMUYSKarv/6Yc80NuhDAFv5m0/19aOj3lMERZ8b4Pvi2OxVvcZq5+7PWkKJC
93G0HrNdVtm0PcMy9e4CqF5kjWlm2Dc2ONPkHMGKWEDlESw0qkIcxfl0a2OFw2gx
ozE7XIUbZju2HymsEA7xZF4lyrLvIW84nGlHfCVHf4EbNIOqiuN2rEYU6KMQ62yu
LfKPTNfg40KAGHvhlxYDfhuKES1pNv3dvigv/Lrd2kjM2C/xTYm696qTDuc7owFu
3JEmOpSNdhk+gFNUj9gdkW61CHh51XpLerKdUdRZ4fqM8t0eOoA9klUlWn+9/YPX
YQH8kKXOaY/XBtFry0jsml36RvRsJ8x7U30UA9YwTkcAMtnO4twzI6H4a2udQNAJ
zmx+MR1o/KqpfeNRpTQYxOhz8/Oxs/1fbgQGhDZiHSAZmGMO27EiPyIwbx7kG97w
8dVtxNtiFo9VWq7xO76DUJZ9ANMLsyJZHI2Lq911LotB1BlezXsGlNNAnpsP/dX4
QNYt4l+E1Sm5WME4NorFNDa7xiomSu6SGIrPrs+lBaUCNGCJWBbpownz0RDCyLwf
8YkrWwq022jUjSadhb8cHR0y/jR6IUwwV63stTCXjC9rFn0PEF0kFfwgtp+WNft2
IeE2/wgv4ge+cqiWdlqiH2MJxnvQGbWHTrunkwx1YGt3k7DH52FoUGC8jG92Jb91
LCohm8nlM/bvlpSwhz5lMJ+huvovOmbdoBnWfQZoPCijOCLzowgiJ8inAZ2dhNdi
JFSRT12Sbnhr3dDycKW8ml8KHMOF9upk4gHcFRh3JEZ3yBUts5PM7t9lXMAyx3E5
P19nMJqTLGPWAqIhyVMcnRHs5qEmDv27BC57miti1iM+4215Dm6oEXBXkh3Alx9l
U5rxPXx/eUkAZxXYPU2SfJGFTHz3q9I3y1uKk5bGIaN1VuCghnltLZxFjhhFYq/J
3FAS4V/FQWBocEBc9roKDkT4nca0Py8IktD3A9MBZUKJOX1W8Kdz7G0EE2ueDW4m
vOdi5Eisl0YYk5Jv4vpb6QLoIZPJEz24WTS/ImQkoaCcTEN/27/gfIEeeFfi+rzO
DzJ1SIXaCK6edVOXh9gsXp4cA1vsmOZ0oF6i4/uCAzdNcenxVW+Jcy7NMAxQkyOi
1qGPsOW3RgUjPMDo72Id7g2Fv1wJ47vAcjwUYIWFFk90Np2+tJ5YiOi0KfAItc7+
HQA0WSU8DkaNNUG9u98VYJQMVmJSfrdC0+ICoReasCqMVW2FdMA+OnjP32Bgr6k4
vpWzQhh6nbOarw71JmWA098IJcb417aAQezpojtz2t46p0dTMP0bbt6qhZ0x7ELJ
wSqh6Z6lLc2EtxsFAXlzqZDAKm8G2KFnAGZZyAiU68pdOtjvyMDBEnQGJjHrBtXC
CKcA1hiAjs3k9LYfA6ZXlSWD5tS4vg7QhS+nbvGqZ45quqWlQhphl2+Uh2onjqzw
QS5oY8aC/u6tgOxeYicC2hFKgJtoZlnz7FhHvD8Mixsc8eFvhCNE4ndtnYEJ30wV
kQxAF9KzdE1UDiDfAaocOUR2sbTcJRuJ2l9oFcC6jMZ+/QXLooIaKTPkugoICFAB
zJrCeMKoTXrcqtVLX4TwFj9PS5akr/gqcqpdD5ZaMDnELQEZHB81jmWGGRD53lbu
1d+/V8/17Ez6GY1ZkV9CJhAU11Zj14AzCQpXHiwBbvHfA/MrMB6QXBzd+u3+Ng6p
uOAeq8DP27Xhx1qdRRaZV0xevdOeVIbqb5a0t3m4/SdYL5Uyxt1OKvSzgF9g5Fb7
6zYl3cGFGZi5EeOdjCJ/tNWpGWDwsuqtKwG9YyLltNlF2hfZXjQTcQ4vr1Tzbcx7
TXeyC/AGBSf4x32WC83YMBX1holDyksvEfZSvX6JuiHFHM9WYc68+449zCN04DrS
cZGYd8q1CFCdUNK9/is7dP4BmluCM2AfSM6GM+zYtWY5T4/tU3UN/r+0xTk312Vy
JgMby223xv9zXpHMpqy25EjrCzF2t/7hAAL2csKAYpQd5/wTBSSDxFVWbn07j0Rk
DFjnJbnZiJN0qkFmb3Cibom5y19xbLe3MgMOQeSM85AsrTSRyb5bWqc3SQp0MrtI
QrOeehWBoXyasjWny4Ndc6GV3ZgwAh79SdUwBGx9whZ40Jkl6azk4ozBeYdA1tQn
epC7M1A33/vgLi0DQTrstBggpmsKu8zbc7C445OKQGzA1gnWKgffJO8pXshJBz6F
uqKzjmSNQg7/a0dgMyeXV/MoX5frnkpSMqP21ZN7CnZrjiFNcPXOu5XLm7Nl46X5
tSy6z3YQGRT7/oggK2QFBEwkfhOWIb/Y8+7NS9LB2ErybDnSNZR5PB+vK21xkvIy
7rWmVEglcGq6oqKOXbrmga96Vn+LclRzcU9+dnu8P3wNicc46TCO32anBOtiYHro
RKzGu62YfFTdZdLM0iyF+BjbK5QnlwfKbTAbKfsoN0P4yiuWG3nLg7V5s/44IIvH
A1S6bmPVVrkLcg2pFqiflG5siwubdlDB8Lr0FBTiKhG6YinCmHAPMcckxHJJMJrW
ynS1Gai6h4H3/CQbRPP9Rmk/ZbiyECej+9GwjTsBvpOTPaLtV1lZREPlWU83dRhU
4FTPt1zhJCcR0tbKf5j0abLIkABlCCqWaobDcCmF5Jbo5NO1REviBdGjHCRXd7ZD
ETR3P1CRGu5DshyuBvOEu9/1crs5B+3c9TxQTjjPwndzXNQwbb2MB1hclHfdhAVv
V4UOIwgQR6jVobj8lad7+EVvdc93jjWww1+UIOKqWONQy8fucxal7fIlN4JbBupq
mOwe9NS93oOZVp51PnhrmFOk0TS9aa5xnKtKPL/eBHrURSvWYYAQ7shG/1jgm9Sl
/GTpKZcUMeqYzDYop1dLlzFk8XpL+EMKv8jRlAHv4E320wKjRL2aaNOfFVl7svQf
U27VWSZXKKWUw1BDKzYY+dRpD0Q6fUj5PQ39FwuJ2dSSx+ak+EVokG45Cad1X3BF
gcgwkEVvCoxzMeZaDuMVm9Ru3ZOnghgKNxOIV+zqVxyALU58tuodQTMLabYmKjyq
KV2Qwj8u4AwIOCkp4wqpWodSVlSVpjWQrXXmTsILDz5i5YzOiOqwv2li6a51yQp1
a/lTf84Sv5NehH6Y2gfrVsqeUwOewSYpmHT2XVxvUsFmqPdenkgHEO7gLe7ybLKd
ljavRdcc0IgUfRsY3dJxz/HGVT05+AZm14Ve9qGDJUj0HUfadCjvWT929wzontM7
e8g+ONxYK1w+c+eWmFBSgYGg+haOxkC1Y9taLsWqt4q7YrQF2b1gFfiYn6OIiMG6
VB2Ma9cXsNv2MmWMcsTVwcQvPcSkf9ISy4wUZmMjXZXz0bUUZ4n3H/qcqQOk0Q61
c++wkHB6FCm4Z1dUOo795IVQpHx4Xm36X1KWXVXp12itxCazIE89XFUhOuBatiN/
qEIWJIQK7JVrnM/3HwoyjeMsAqME0mb67s3HyXcTUwGTrTBckcGPINHrB8q+tNch
gpcsVdWYldEwtVzpeAz7YI8O25gr9iDDmvxGWBU9zsv+62jv29lCyzRKRFn8O2ra
7Ol77DyGsNZeQeZnK6pgHpTqgjORT6o+24+tOdGLMErOnyHGy4YKocpyUFs0c49c
WMjOBDj7uMTALm62XoSPrV84spydtwW3kHb2kx34iBd0O8kjWI1u3eRVpI2udRN8
WrBAT/URfEOO94dFPRfgtwTSSskLZlURR/15HKmgVPFtrCpz3iy+npVH1PW2i+AJ
+swbCkMryMo3lwVgjRoh3NE+St34mCM7y+ESn16woBj+qUtTPeXfSDiGRrKFjsvJ
zlHAhCt4Dqx+pAPDl7b5EROubhADxyoqHOrTarQXVWIvRrxANHTWSPJ0xnbQq4Jz
y8beo+O9GhwIyljH0tMXTU05ghGGVs0p/DyeBdZECqU8xdaC34OCLbA/KGFAvHAd
EVnpH9KCQeHLJQ9yy1OtkbE9rLxg/g1oQiQadE1FIi/b/ziamEQ6GEJG4ljC992M
NWuU/sdp6SYZFF0vJUhR6O308lSo3w8a4q4HgfdOOxFL6K4CqiQ0CgEsSyIJIWK5
r27yIaTnd6GY6G03ldihgzQRapr8CnzxsLy3CxBZStKkMCuPYoNw+kP4IpLhvc0h
bCaQ3dANmnbcp44k5Ydn5x81lOQmRKrpq4wwcZCefbVqUapxmwW7x11rGxSU6dVB
GxcUki8ES4MuQtxodEleJ1wzhC+eWzK6H47HUrYsRtHmwOLb+RtAghH2KWs+ssTZ
NqUwV2lIyVqFgRNcfik40w0dgZOdEcUS8nflyVofZQtGKsL+/097rCtWv1TKkb/l
c03v4OhzQMlodHF3UOyuhtH+GgltDN8pnt6L0nkH4SrG0LthnmJa7YOkmQSzVx+/
NqKGshMLqmcRfcJJD3u+0hBIzOt212lwdEUMTPJPFjCeI+6Nw7Mca/ajRidN7nR9
XSqK8IggY//0mps0SjdjU7VskpRfapQC0xXNTcSgIOdZ8kBzIB9aeFJBjrKF9XSv
R8238vJ+f/HJa4V2CQSWG7ErtF7I4t7ahEds3kr/oqQIVSisKnbMW0dybqbCRUW6
QErfS/k3D9AvvqDo9034L654+nSS4gyXIQFupqrOay8xo2P/hf/ZJNkj1RVTez76
FB90vDVfzTg2ROwpwWAPsOdvrTDKKtS/AtBOKQFl9EMsFOKwjAisXeOK/cfYEPyp
tWQbroX0INvaHiHVk36DU4/hMC5xdEFp1pYafLRF8OsYveAtbwJaQrZ8faSPL0gU
JDoks2AlTU909YCqREajmXjPLUUxq9pNNqid4Zu+jgVkpFYhfZotTqcmLajgT7FQ
9xagNe2P2iXcYDtzwWqvMfT1YAy4Gjst5us8wdzBQ07wCOPe6zcj6qKQKxAq46Gc

//pragma protect end_data_block
//pragma protect digest_block
bGwb1wLowd3+wmNdus8QimHuMo8=
//pragma protect end_digest_block
//pragma protect end_protected

function void svt_axi_transaction::pre_randomize ();
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dG0YhYheWcQHREKIbvk8NcqZG7nNML6vCQBOrnQ9b1Man/UK5OxXeabL1wEPWtz/
lc+sWpkhiFtpHCe9FFpQKlRAh7rTpxb/K59nW1Yz2QjE5LH+CP3Z0VXxpwN043Cq
9wLhhzSOKTEC91pYSW5Inn7s6AyviyIYpIHBl7ie3pTaHAtNxQjEkA==
//pragma protect end_key_block
//pragma protect digest_block
itXTKAgVs4mLTMKg4ESQ1p43FqI=
//pragma protect end_digest_block
//pragma protect data_block
Uj9wZ43tZ5GLmrtTie2Npybh4hh7KSVcNRtagAztxXay9WI9CuK+MfGrt9Hty5A4
nmaND1YAX6EpDcPWup40qfSIwQW4/ma+8YOKTCQ+zuWQZBtL2f0NnXz3H3XMfYMs
S5w6AflS0Fa1ahOtNCu0rzQr0qRgn+ir6smIH0+GwSOIh7a0HpaDlHjgXOT6/JFw
iI+MUckUSk6YG5RVX4t69WGUQy59M95/YjazjMoIxRxLVdZgxeDg7dW39aL2v4AE
218ce1fbTqq6RUOPBjtM+tBcBVe/G0KH76rehzTzjq0QIO3LVpIyPpRLUY6y1bd/
u5rBsuY7P8WfRi7YVfkbl4GEjPjEt1lYy2ffK6gSWcu2p6UyCtUuZF4hXmRp9yww
x1EbUX/XOdYoIEDWg1lCR+ZKVamhRFEhRKgzsNSiisKOMsyy+D/Glao+uv9NZV1j
5vh3axlUxjzMTjGh5ItjEdZZcngViwbkB9lUhNwHtzpmvPsMAAR/rJ5PEzYqWTAS
qPkBrXB7exa/qwu9JoLmzFEr5NPdwCONrGZ6uTHkyKrZ4LV6MwY+Wo8oogEvSKsN
XEjGiCoej6XbIjArn2FEokX3Jur2ikvH603PgQLYg/aYUf6GBORqfP8kRKrO039+
vX0QIcUK2P4tYTGcJGFtAe4a2ej2a7ncl+Bd3GlVZ/c8XiEs/dmUcS6mHPQRD0Y+
2CwaryKmkpmB73SI8OhaH0P7VijE95VaSEoE32ZONC2cm9CxiDKaVJB7qOEhiDCs
gFJQZZCOBY7KtmuLEFr1PTDT++yX3ZLlTwsXzX6thKaBNexObEFI7H0kRtFoVr0m
heRiPCJKk/0/SWMqXM7/Vql8SGzOS4v5xOtkMgOFk+bq1VA6mMJ9N0U6t5iN5uye
LN3yQ7ouvVCOQbvt2ycbojeewNjkCF5+AZAktZEzRtCb3YXofsqMVOfoVvzfSLR1
fIXk/ofXKYGieTN2DYtX/4sAUTaTbrCpEIAk9t7U819ucj3h+tGKLXpG6WPjmpr9
cT1JGL2VcZngWktD3Dbq8Fr8ZzpmmPZCZryByIk2bNXNlN37JRu7dFsRs8q4Qtnf
qvF7n+Os+288kjdpS8jpgzl6rGe8Mp7bu1CpZEEdkcu1+x5o/AkALaygLGkSgQsF
KGIuVPeDB4n96abhXIC86oJouAwYv7bH/VyMmRExOHIxkseFX6w3M2DsLCW2MBni
GWeloe656qSLd6ZRHQAIfFkpfvd6hki6lPpfm5KdkQNpkAyTIxC5HsFPD670gpfo
67F2vBjlXB4Ai+Kcc9qE/Q1rl4voL/0ZE7+OzqSd/vnNtyBxUIqOju/T3L0UisW0
xrnmbDhed1i+P1WM0e80JNVvtt/bBfosOD7MZl0uneTBREEqaiqwJm/QmcbKZaLP
wdrmTVc/gbbtQuyyt2Yx0/6c77GvQQmEmd5B8HDWl/5GRjKVxtaijXY6ofPHPb6b
/U1T6jEgWlVclMeWfCHD4KfICyCSX5lafPpjspvtIcAHVPHkZwuQW6U0KYiTucbM
Tr/SdogqmVMLTGExHsDqd5kAoKZFOUjNpG7+pbI//t9SonIzarZiMlJVQLLTIA4P
jdjh7AzDke7szOdTWUglt9HL7sR00vd/BAGFygkVZKPRsoSLW65fHHz+5fEn0XVL
XeSn4eF/vNICjOPH50ycXPZhWT02f+o/LMlijFEKz4h48Gw1PO9kY4fPNfkX+KCL
tzSXiKkZjHyk6sWtSSZFypT3QSCBxryuGnachF9fqNUwLHeTjzCTzoblK2GFFj9N
UWftvtGZGOmump3c2MKcuJfjfeo0dv5Wq4K3A9Bs4SOD2iSFMh6jenIQ8VW9raSx
HIBL5znWceGifC1b4+oKCvSd99ck5Qmq8/4JoUH3Nr5we2Gohd2qDNHVJIJ5t6Se
4bIBqoWCiJ6wxkMHDr3hbwXKzU8MHA5ivfQTQPTysqIJnDQRX9jX5ace4b2N74CH
xX9B948bbISIF64fLtgNoaycZguGuG5/Aainr0Q+JcS1TO2Ii9kEeG5neiwafy+B
6DPLmv/WB37M0O66YhzdSCZ0eLktuy5bQEZtc9CXwbg4MRQknML0M4qM4Qn1CCaN
zN9dJlkrH+fHkLQgAT06RdJa6lMyhWNvT6HqUuHzP9GyUcD8aLSBruB8YbMgMSK1
j7S0dDKjA7NBN4A2n8PZBZZ2RD/WTocH6e+jQvBGTDm/lGzSOxKgDPnw9IQFTUh3
BLXKwetrA5xFSam61EUexfXvF2vsH79719lFn0ToLQGqpWFlxZtxt76DKmsXVlwB
Pe2hisblA4xGBoUFpS1AF9g9H9sm7ZdJNbv4fS/MEcIrZf7ijYYBNiOxcHNVgf/i
dDE0Nuona5rCtR/K1GH1U7qeZZgfopNEaXG14N3h9PCo3LbO2LIwVOLtbeh5F4X+
X90rSRNvERLtqFL5xptZzChEgxXmOIvXJCGIDZj4zqRsZQEF1s8zqOlLMfB07Hz+
DP2HAVTpbnxUpwGVlWP0so+lGQUxvfNaOhx4prQ7879yNoFAh1lYJ+82G9PRIfeo
Ca4QZwZ7bTI0qTmvFhUfbNBXHcOQOsyIh44V6ZoS+VLoU4H9+W4C71A26xe3VXlJ
vf/K3uKIdN5gWgBD7x7/Oiuorjd/xO23SgNABoCLtRfHGznlyDLK5WCWiQDDRRl3
JhIBe4+9gk8x1mQA6mtOiLtE8I0QgXlArkOcN/Cat9b5akhNv7kJ7TTT4paEKzdD
q1tLYWt0ttVMDHcmCygUuJPFKSerdrAuLhTGddEchpV5xO2IjfP7daF7nHph5QL1
gAvcPko0045pisTXDQ+oakvRz7c1ABIIrQPTpzU6tebuaxf2JJWIymrkuMnPSHTr
O5d9amb01Fo8G03aT2m86CM2nnauZlWrigxirDXZpDyMWm40BOa1y94qjeMzmX4L
009IyjgYVJC44UZ4Qf5ysEKcI/PU1fo0Q7U5pQGcpcEVztsO3JKgPqJ+90XnwzOE
K/rgzz2qKmxNHjzhQWQw/zNTgRj6ARPqZB2lVWc6AhPiZ2MblGgEeAtlXgt4PMON
uBxmOGc66ShrQadNBMEb54H5vBcdOuObSXqU9hd4z5RjJ1z42JX0+eDZqiEQ0apD
ip8qVgqxa7WWVoQz2gYlRLC8F+PJx8YBbICi3HFq6D4ji6slOyUA1IyN3LX3U8qI
kGXPf7/0j1yZqxc5PaHtT5LFvT+MVhGrk6rcwHufO38CUUCBilYoWQwLE/KWvMSo
1yG3HzwjB4nDRG2NMpJtXrst73Ij2eMimLMSwiVVIwS9k2V2/WJLdYFbNV+GQBIi
8oyO8oGKUh/NQdFxRpDUSPLq4pq+Sza16zG4W+D3uos3swccDLrMAhXvyIwksAwZ
aCTYGGQWX+m5fXWOPE4AmhbPi1Vm2ys7q5whg3gmEVNSJSnNdY8urjutCmkMaV8+
yuuVScfHJ472YZp4+0s9JirtKiCS5lc7S4A1iM+Jar43bh+JSSgvR5zaUZ7Xuudh
O6sE7uCc2TvzuoMZArsJliXbdj396mRCVedBGVsuWQqeQRJXvkE/FqjzuLcnPJQp
SlR9D1yD3m32XFe+Wu8ByVtRHZmoKm5wNJlDJU5ZNWi1PX2uSre4B7eqK6gdnliU
7U73/U++PghnbAEhRKp18Rs5QXniNaztu+WX0iBmraKv4w75QLY0tA8/+i2HqKU1
oCkbFVagiPA8ywfbN7dtNqW60SEnTH0qBF60wXXLP4QuaT4TbbPhc52N8RK+rNig
cCtmIKbV1jn7qiCnNPUpt8ywApD+DXRcgRBT/QBpC0EMyJyHQpSF2REmRWpTvrp6
hoJEcATY2m91RI6QzM4e6OYuDOKchD9/gtctmseSlnWsLaoAI+HI64JGN5PvJ+dB
TTtP9zehwfVckYLC5Pwey/2hYsFCbupWIBf3D7iqFXfZHEGE0JB9r56N4eeP/sHs
PQfrpcWTB5hx5K4t0Px1tBlPQwCopYUJevcPpit5CuJRqXxWofDSQnfJ8pljyyXY
ivWvv+aavfX1cqC5e+VD0zZHoLLymJ610nbDbsOkAh/ZBeV6+mJLglAvAj4KpGPJ
/j3S0LVcDjbqZ5q7kME3smK4xYyJ0xaz0l5jAL2gNqTexUHieY3hEJdYutoBrQsI
Nz0aap90yhA2hreP/oRSa9JtZlB2/AtdRjgWZDOsqU3eRLtIPt6xnEZ984rtSs47
gAZWWybEN6SAJ6HpxqhOPzdEd2X63NMqjz6uB+d7/QVuxOHl/eTQ+R7141oS4Uvv
jEybQ9rAVeredjD0jKPrlPgS65G3XB9CCT2dWzwgVDlNnMKNlUgQqHp86K59bIS0
Cp7ouV0v1hzyKATAakyoNATriajn44fKoqKvexxxOrk8X9IcuwaSaHQsYwT6yfcB
IqJyJAtRbKMW5jEr2HunCcwx5fEH7CHob2I/q1LUzjTFgJpbcNJ/TQb68AU9XmIp
ju6hzosTOo5B8Z0SGneK+0WdGSLNfvqz3ubronjnu5uXok6hpwzBY8OogS/yMNS9
rlb8b5bYTkYXgR54AMmszFFInNVm/dH1E3+vXNW0AZgpxeMmJmJrAzwzlgpd76W0
Og6rv3BNxgg/iOW2p+3S4w8jT/+sdtYTJmLH2y0vBT2kucGH2TcbG8zrZvhyDXAp
owsUOfn9e6+jkwrrSZElgjcUYUiLeSV6K3i95PbaqU9FuiQD36D+HOVz2QvVmEN3
7D6OHv+8qDDUyMPpTOIg+NzDlSAJxYDGuPU239d7yaZNCiE7rmb4GlkL1u4R8d/0
z/T8lP4lPNkhCssZWvLNDJ6gxTFFVUmtPCSB7vO7ByzFzbc35UtVw70yaGpjrcpe
mHqyq9Yzd2Ep1X5zktnIpbPJZB8LikjZ9NcuyELIqJklKNBAUlTx/BpWWUAnzoct
ScBbKlBjISnDMEuD8E5nWge4pGP/OE5Y6FXYZJfY+qHFEtwTDD83XGB1nywT8VGD
C87Znk/AYfWrCrc4MTjrSlgcZdAsKqGflF6lEFshE4KIVA0NKdIEuPFmES5vpUgf
CM1Zna92skuEYg79+GCzVO0n25R5S06OApbI+RATZ6aQCclz6N5Q1Ba1asB+JptH
CkvSkdE9kZpPhPE7raqz7C9gE3t4eqpiGjjzjrbJUB97nCreLS43RPlrxtxHQIs3
Z8LgsCFE67AF/VFEZVpfHNI9uYWkDCVoB7o8D6DvuxJ4tUXTHCAh7dNBtXmdsqT+
KuB4cSyW45iPCnRw+PC1CeV0A6t5b7S4u5HG572he/947SXe6tGSQOu/jyKX9xpt
4jxaxXD0Qgdmzt8dGjUtKtELCUsHg1CTNgPyjOJ73oCIQUSzsHoXOXvKtP3zRt4W
89wsuXqTqWHRuNpd3m+MDdJwKKjnen7BSYICTaoMkVePULK/inelTx1Q9J+rBWcl
mR0vsUEdJrjoRa+ui3f1Pm+3GIf47QlZkFvjkz40OtbVRmbFVwSS4ApZHyC4KtSx
STkCpQTc4ni5+fckjrnfvn5Ze1uvtOa8SJlI2FWZVcg46ZAoG6qUcQRDbXO82s40
9To7HvypvXkMj4kNSlINurttVJ7zbAzxVJv3Ej53L90DkY7CnzN3wCfKOpSi6lDe
OwFVUFMZsgODIFtJx99e4yM6W9oXULL5fbOu/FDDIpKQTS+nvc7243DcNFwcolW8
FHWpb/b3iUd/c1qL0bwa/MiwtbPlHTtPiO9Han+ZYyvwHqCL/yotiF9DHMEFwDW9
pws6XvkcSvsUU3OedCNiIRe6p+/9YFZhic7FA3VSHPHiZbvmGX2k7sEJgYSvmQ5z
mW5ONQ9ehKrcUH96iRleR+xHrmqdoZtLgEGJmRSYAKZQM48F2PdlhKvqEjphA8XT
HmlL32CIm+f555C5ol7JQYZMVABRPLAU1AsuxtmSeRRpeWgy7NA61mJsDav2K7q6
SOViaLeqvU2he+N5UAsslS399QlYrdjzhvGCGEibPcA8UcU66hOphlRGCGRrxKgL
74DgUGXPZqwRKCu+yaR9WrPcwISU6YoybRLBu8bpcjFI5dZJBRZIz5wega+LLIx0
Eymlt9zYLUNa6z57KZ0lzo/4uIGmVO/8j9W0HJuaWBn8Q0bxEp64hFb187Mnyw/V
zLvDA51Dma16aIElbXTyawCpNAkvXVXbwcvcP0f7WEo1gUY3OcIgciInTwEy+bYn
z1BWOlvdY0O2VkFj0y4zQW2s/PLXvJQjPQSa3G9F9iUo2V8eb8cN2lh3SjOCjpB8
MwDdGQTT6qty2ekvf4Vli1SPwPD4PYLEsd6/evwrwZ9gbe9t8u+bhqtZII/NZpRQ
CoW4aAXdTH/MJn4I6R+mE3Z3IO/e3P4GLchMMs9ap8Ycd5ZGTBaynajGGHLB3Y9S
r7QG0jMJz0YnentjWChYHnWbPhjzjg52Nx23pmV8Z9SGzlAGezNhC5+BhKqB7mrn
1LQ+Jj/s1Cj0s9zlkhvUDErKjq+DLeZhWpm0rC8ruY0ixLuh0XjerIo78TdIX6Iu
jYgLD6QhEOQlgygY6L8r44XNdbnqflgSRQqYbNe+thRUJhUupefOPH9vQCI1wbZq
zR7ui7zKWdI4eBdEtaA8OkFzVRJugIs1FlL8QDCQHi0dpAwNUXQF7Zf8D/4OeWow
6FgMOfc3hjfdYunjIoSBVmTf1qFCBS7kLUmU5GCWuvvMOy9FZqEAx2RMBN73DrDU
OyTQFhnhpZOOwRySyDkyciyYe8imLzmDfd9C6HyhTOZmSLjgq9k8oGHd+cjYUIhK
bsXIZ4yZOi7TU6KGUzdsczizdgJm3S+CfvvilsZz+L+V2z/Nw3zlN5ClXh4f5/HM
dbLb/DyBlnnU8tdgzSioSgZY0mO0NwommcX4V7d/71OJ/CSazwihAwAQekh7mBkX
KZXtLnmmUINc7UNco3+PRbzbtLUPm1hk5lJOekKj3ge+RQ9PuamZVrtkex4vsQNu
BTFUC1glxnAzXHDjI3R1H9/IKi3tMqk3ELNmEvXcjNfnLoVJXfDNzytIHUfOoOAv
Zh+/KmjmmOgx5JeuERFohlvtMKx+dIn6cFlfM4aDI7zyPPSi2CMxqHsVwCWxVh93
M7uGOM/zy9r06s0Umq7h7H8x27XC70IT6CDoF91uxOPywk1+sS03qJtAKjig4OxR
+Qb6O1UAG/sbSLETNDsm/xhvdwpF29QANaTNAmz9lkBOdfU9n7jnKMWVGrGoM0d0
dCm/6zZnO2H/hJ30nF9hr9/mXRtz4+GoMZKjkr+iuP3xTQSfCzzRnFsGJPyGle2+
m30ZsH3NZ/E0xSs3biXR/JU4ByizGjI2V7QxPk4DUNVLf4F2NFrTVfVoR37/xbIT
fYkDeB7CpLafk/swXJk5pVqSOnXQ9uDm+2v3Tr4mvnh9BHnBwuFCblNl4k6q4kcV
3DtL/y/lf57ieMmF3E+c4Jt18ihfaUY4YTcssiUuI7ImPROl1goSHAEHaNYV13ES
9Y/VRB7Z7230h6MWwO+H1fdi79nMpmfmWzsWP6dEUoAwYjFYSZJHyKDWNuWLL6KO
w0epC6mvFT01zosdJ49yWrW7UOG68wsx4Q2g2PNXB85Je002z/9x0BoawlrGj4N1
7sW/n7ym2+OKWyK0cH9leh9f8hzJlSNy6erLB6QIv72g6b7mvPqxLVil0/o10evk
mNww5nIZ8lu8l8lafucN6OrsIm3Gy2J60c15WjqjnNWf9U2xAueHxxsEROCTcG+g
fYXTaeECOXGVa8LlMbBH86eseKPuBuOcZ0mT0XX37p9US5KJNTKCkltCddGj7SrP
zLrf2Fs/K1HYuMCiw6d4vN3qn9PZ8kyyyHh89jeuOFxVXZoWGeIXWtOruvF6Og7Q
6XMK9iDtNTdG3wu0GYVsojGRMfr1WUxIfrXos9uozgT1RauLLsdk+ZX3pH1G7fZC
emqHNSVqbuhkYwiCpuVmsAnpFU7JU0SehK6JEyvObU4QQJYaA90VMfhpSPa4pqxz
SpfB41WX0IbpOUGvW46BireWMz0XPy+6A9HYw0tiRVUmIlCxR4FyzPqX/xEgAM7r
O+gqaYvozrLdwN+BWg66bxHLkDu1jQZMnSS7XJJUb3nTy/PtfBBIeySgYiPvHJvN
6UN0s5hZcTQ//IW3jON/nheQiSltw4tnizNyrMRMPdlJ9tnNxB8ClEmtudjNSJ/y
LOuS9qEszrpoRSFxFLoA3T2KXl5qWBrfZmW33ANpo7B8FD9qZ8xiqjt0hkrIZU1h
hSZHU8XEn/Wyu0UlelEMHpBEFk9Hvjvl2rT25GJUcDlOhj/H5obDgSkTHUdHJVnT
e0B06mKFbRYfCIZUGLRUi5g6jJyvcVAy4Wxbx2BfSnqsrQfWHqfoLLfNMq3FKtjN
4TzpfLMus9V2jBnfYwI8N3tQVTqZl3fpHNk6jtMEa/zrTQSjpNwmtWSvHXaM9i7B
CDwW/C4yihk4b8rV4FhFFRJzcxeJH8REK9R/q8gBiurLgZ8mCqzYPH0/1yb+M/oh
xCFBM+O3UBL4OCe5TOp9sB/1yCBOWDTZvS5zHzk4OMLvz3FqRfkn1T4nhdL5Actz
Pt0cydDlYv3NPFGgzYtxeoBi1pEWB15WdlSoalgmtNZN+uFknejso5aMbBVs5wJb
CeQtWF4suZDA9Rs0HHuUqqcN6FaMkCTNneNVgCSinQ4HdFpOO419Fj9ny5VQq6B0
OP1qAGT3QfxYwCfXijDweaC6afLMZtQi709OX5Uoot7bdVUEpBGub+2ja+QChflz
fE3j/NPE3Z7CICrVqymdUH2+w6nswrhHU8SyXshl+chFTjXuZWG6Agh91etcfxwA
nTib2HUxyMcI2nTBmWvK0ZY6Ws5R5o2eslsTy80DRTYNSPrqpaTZwdFH4G5t15zZ
guauW2OCl39gxIH8QfS/pP7HpsTRL7OXgBLX1vPCgUbfZgb8mRaYsMqxqIpIaWha
gURkMn2qDIMNMnH9yqy4Us7WpWL8iqBV+mQM+bJR4EYOkDE9vBnv/kjxTKXeAFdr
qnpiiRNqoNKd6bMe5YuVeSG1a98t3uPS0LzFm2Pq7Bb3/Qz2l0xtQRqMM/lFN0+2
0fhHT4fTi/huka9E7BY07gbEXQG9L21osPrHwIv7xn37wEoto5oOcHTAsVEMvPrz
y/HbUvReMJcDH7iVPiTCnCnXLE+2bFGCTasxNwTtYEutSUSNgCquaRzL6U65f+Z/
bqJp+iui1DqdMLjn/+M/tgt9hNJI0ZfyuVqr6V3J7OSgWMwEPTBioYbouteQyQPJ
4fVl+sl9+/J95dD+FSZrD9O8JcDqcogIPSHEnX7LKsiDVmwK5lO7/vEDdlhxC1xg
9KQ2762vmsA7EDFJLV2AmuexQXHRggEPEisJq/JnWw2TGRBbLlMfru/YsAzdCRHK
ViBMn7Jd0GUxGnruj4DlGMDZ44ddXuzvPQ3euyvPIojzeObBcbCr/KKcPMIbSMJS
Z6tlIPRb70uTXryUd2cM/VUXmtHwfyZiC0YNSXd0AJa+7tW6VgFnnc+lbeOA8WZJ
yVoGydu2P2ZwKiwcJeO2gcXYz/Dp2NLyOiRfZgdXPZ5vL+0HM6lZVjXwr2qbDN9l
ZtJ88YEr+U7yJr6JXS9LuJa9roXziTrYHQ/lvj6vi5jmGpeIVBiru7wNDvoQ3an2
JQW/7oGpjXEawMqwaYxQDrNEBJAWH1jiXMKbMHxyrEh+EaKbcRqQJz56vLYQ4tO/
NvC6mCoVeS04l4yWOVxYi6GlpKzFyME/W0tBJ4/pJbgdolhQwq2Qv9Vc7V+bNxLV
ahnd0h+ynnrqHVnYaWFXslQXe75dXFLpEgsYGo5c0cbuBzpZyrOoWXZ4SggRtkes
hRPK4nbYXp6BfbamL5rmjH85Ms1FqVnBksGe6dJVzJgD/5XiO9AtNFh+FQiEvFm2
TLNIfpfOstH0dILYldiKMYPpoxRta7GwAORa2uIpLmzi5vBQkY2bKBWgoLfbGGrG
Yts97vrvFT52qaeXzF5Xm56aLtZo3eT8In9rJqhe+4AeQ94eYpYZApQdoN/9KTk8
ZH/xUsQMf6U3HNYf+AVSM3cxAp2CTTEYJjKZ2BFXORlUcMUcvtVkJM7wBj8EESHV
Z4tIUuOHWdyTAe2s8SFOp5tg/CTk8mMRrteUHkWNAsBID3yh3tfu2g6cnY5DhdUD
hxPanoDXTKVvrptwsHcvPvlATw6xHj78wTzQ9hEBzWApF1rIAOaE7umfvj3Vb4Qr
PSyGHWL/8x2cwI5bjC2tvZoqq7gAJ7TSK+Kx0FyZKc40o30ZiGlpwKOhskYEsztk
4Rlkz3y7zdJt3nfkkY34cCaQDz8va9DSTx+jr+bVBB1UVaasEKm5n5myfUjBDEei
MbX4cbY5k+JKswV68ONhfMdLoYSBHPvYfJ4bgNHOHaJHudN0wI1LwGN1lbHBA85E
KqotKyPLEkak8CrpshQeY4KnY6v2JXycRBsXPEcHBRQD3So8EZ10OHeiGiJrAYFG
+edj3jF4D5cZH4pcOBRee/bLnjnVpUG99XpM+dk6tbSpk9Ba99t1bR3JtdMWf9qb
ctYvoaHeyG0DaV7N5MSd7LWI3Zv9/OgrZWzCUl2UXxvv5TI6+BwzlkEwgi4i8Gtt
LKQxX66JbLQanqzvi71xlI9Ek9+Yb8rfP1z3QfuU1hiHm2j1zo6hZ3XAXkIXn1F+
Z+oPztjWqhPy7rSXdjYrQt5/iKCIUx221Bq3PxiEFHOnvyLe1ygonGzhmZFkP/M7
qKy5LlVdqHzNksW/hvgh5K3a8T5t2fhkyuZfBc3Ot8tYkqZda7xXNidDjp6U44kU
vNaSgwdC0aQXp7dvp7LHZDLcKMePvMo+OwXuwVhmi+5b4auocccv6M0DOjiGoFFv
t37H+hfLXC7709/zWFCO3s0NdwAUw32EssV8ULG2vPgZ42yvv1OrA/gCNKDemHyG
YAgWCxwkkBeZh92YCmsP205z4/CxtAh/ABKz+lWSkA7ipXZ15bzczS8xmWIzcGdE
GwKll3CiXHDgSi8NKu6T8f6Sz+Y0nbkPGreJzeFV1MHReSOhMhrPIY8cutykxwN7
Z3vnR98d7QOwglVnRS4camt8Vro2p1L4gD2gX6kDDByNq66ZJn92YQ2UbsMAXTyn
pPrdtyEwmdCkafmWO2mB+znCocwk4l07BZpgMujGrMTt9yZ9eyWE+8wAf9UHSqBy
EgWuaw00qLmR8eABF56sFrakw2bxZcXQKfDqjMgLbFvv1Qu3a2HovYoS/4impnSV
wZRrTADCutIF/7yhOaIT5oa9iiDJLgpIDm7A8tGfT5g7TCHU30Tcok6uBUux84MZ
iYoeoWI6UFa13698EOhpyV7SPCLzZKLXaFyxZ300yNw2cQRtIKsmmAoenTreijLR
fqOaFcdXPokYXRlxj17O6z4C+bl7mvTD5JJB1GlHModF+Nu5Xf9vtvzY6UloreI8
s1ki8XYq1Q8Z7VHG8w+dFa6J3svo+pXHzM8YDMVvNa19+b63Qd6w10wKE1A5Sfdr
8SIn8M1pIdDZ4aq+0okwyIJC7O5i8dlXa0iJOk0EI4QXQGX1v7uyIIlWo/t2J2/U
ahViEuaF73q3cObg8V/x4RJHm/O5I/c6Tw3b0IHuN+e/r43tSqB5/PTygWIh1LMr
y8MDkSDq8Ugoq5hhrYKAfK6x6hpFx45FOBl3PjJ7gIDUc/FrYfEZyvZAY+V/e5JN
SbFEWN7bGAXBcuIBH37LlxqLTpGSjB+5/s2LQGw+4RjiPxzDY9US+FrTTH+1FxS4
C7WLgxYDZcH6UXjTmBug0eMF+gmOi15iqPWFpVObpYhANyYKeYxnD+yY6NY4Z0FT
WJ1FbUk6UZ94Rha8BIEoBWIMJnnJK4IlHuOaJ1aYQKoeNzm40rqTwwpU4DFEgXeP
3+WQcfvSs+RK6gsIA9zu6SGPoitPbvyspUq7lZNH3o/i1qr7Bnruuvq2Ao3/ypC8
0cDPpA+vIFI6PrT3P7bEO9bMydFiZx3xQCfS0Sso0c9KNDwsCZkplkzF/8TYorHj
Qie7km5P0XvN+0Ej3i12OiPZSeMOA8wyTq9AVpZ/iwJKfuLZkX8yuqzAMKtTMjw0
y+mUQm64zualpqgDPc+UmRd0LaOHpbXxkBmJcwLCgp4L/tSY4h94C1wh+3T4HgTL
jQuvQIoEmo3zk1qvfG0fwGmgP+Sugw/o/8QH1MzxELeoBWZxyC/oZdeF46Rcn5Y2
rAQkB2HQA+gbY1twS3vPHMtvilP71h7T3UlHWyAWoIqh3zisvmQVaJX6uf7KhG44
c1k5Qr3r+PoBMP19YItFMhwntCfLa7P+mT+hu3oQ79VlpeCQRyXKHcVqJZnfxaKv
E3gVWIPD+RBV+Kxd/2BCwzXgspyeyx9km357pMuUCC7si3QrXwdTP1E5tdBKuWTW
zPJd92XQT7IwP79sC9XwJhiIz6hXvv61QODrybR5VT1QbG6Nzdt51GPCHfAMAAAA
caPG+qts6zcRNENsr9LVvspuogjgN3LdkyJAKp/FEX7SuhCCMRsS8qR08lY5Rmrf
xxZLAhFNvNrWELSQYccsgqd4fVISHBNvBMCoN30Et/Gup4FJgQESM7Kwr4dbCMOx
vh5zXss8hIYSaX2nQPXGRUlq50dbnx72eYwLGrdOqNNXxJCywNYKgk/w665smaYV
ZOfmmXw0LJGFKfhV0wW0bWCS2gzwj0BUeqwFIGD5nlOE3b55GOedl/tjGPqfVMUa
AVZj3xgJbYAeopJ7mkEWra0MFvOUZpwa7lRDdZt8m/0NJuKGEt7onTOXaVWMKHi+
yCN22Vx6kZyl6JrO6rU/3IppBFynt+NpJqfZPlWfunVLAIXz7O+H121pS7VD2hBj
pdi1Ww8uiG+q3+P343CI6feLM7i1g1AtHsqANrNX43n9sI44C2OsAC07MaKjG4j7
altJnndD71yXICnjsPs14DCFeNFN1KxGOaXSL2tHoWWwBSeF/obFuZsTLhnJ17gv
ybm2K4XDnqWBXSlUCNRUZUSr2DztIBOaWfq5wXxmxP3AXAAhp/rPisbv8OOmQyRR
+kYE1E+d1lKN4+8tTU0KQQH1qdK38GF3giWkcJfy6voyPknt3i9YlQJkwN7OFagZ
9ltm7/70WJu1RQFyTZvIhAZGzDCQFHYqh7hz08l6O8v9p+epkMeAjl9BiwD51WLo
IVnkG9WhZdhrf87ZPIuOWAbc1uCCum7lhayR9yiqNLkwHxw/gszQOScLO7+D6s55
FYh/6rSTLRqjEzyLrISuU2BBp81PHlhdz3qOxt611S8GkxZsZcazyf+c6XTuGFde
5zD/KWv1aQUrPuLk6sT6NHywhgQzzBBFXTxECDzE7EWC64fr8FCKorg653VZqHca
yc3dQV4KklEydE79nZCK21MDZicpkoCZmtHTF9hpx8Fzhl9fFHvFprRtle72N+D2
PVeZuPdNNJU2JZne0kujy74Ay31kLrLnPuwBTCl+uO5Uooie28J0rZ81+h044bTj
d8v9j99DoPphoXqlp2nZniNq9iXicnLAa3p0EdWn2PUdYkUiHaU9C/kwuWoGqlo6
3+JRJUzScDSculMvIwchMfXF2uD7Ftcy0HlyZIdAMbMUGYxEGzQNYoFcfLpWs0eW
rcSkSeyMaDXwldERBv64W38UtPTmBqpYeQpPf6W9DeZAXxJ1+cV94jsA9xNKGJIs
K9AquvfisRde3iyAvd6+TcNfhIKbbd1blGO50SBXTnYK7nYEOeZoM9z3PjVEiWFT
5OSHrheRx6KYkCFlafsoF5LGlXHrzvwNrIkN0xb34AQrb31gFvgrz0lshrlZXpAZ
DqYriyWbKKukhEd55CiC4rAzBZhYhVYciGXVScWuz2w9jTEuE7Ho071K22ZmPbgP
E/7CWnYNyDeBE2YmfKYq4ZRBSTRyma9/zjGYGeLfKczf0Huuxv0jKWlh2wBodnkP
9xwiTglx6x+6/3tdT1dJUFBADllHDtuS0Bpdvb9L5CsbbUtTlDT/C10c49LMjTuE
sdATcqvwZ9NgkHJwyWbDd5ZqZzRjvAhtSDnY0ZcyWQxHJctCAkZzxNIOiOtIcRNP
nA8diIF2BwWhcjkhdqvRNq2QTZqArpfyq/ahRDPUYuXQq0pkR2BMEt9s8XpqQvfZ
mjRd5K82VY3U6SATMrnwDNmY+hEHylSUjGA7p+QNj4Xm+I56sNBCetXDMJEbvKMH
3gBaRxgUXI4XZrqXUIdqOwgo8mhTShw2XhFxFj/1fRhyr4OXHOolLZtDAv0vXlo8
Ul9b1CFLI6Rtv970YlIBR/ihFL5qnMaNRIJE1LHQVLDAmGnLjxQ0h0NNuTCZjt82
zaA3apc4Jb+SbpdVrUE9ZFb/wfs4hCNoyDuNpr31rMAd3+OqfiCFY1Vmy56ChlGU
jeonYt2UpTSjVov1bfPs1jDg39+LbqpIL7jnsWUvS3/trKrADa/pMV+/iyT5dW6P
/3F1KsX/l39QucOiP1rLj8ECTQCRcKHEPVL2fmxiaegkIHtuMIFgPKJ0SWqJ4Pbj
A+1VbL1dyT8bKiTZtOc9t7Reoy1FuH87nR3SAneKTvoj/EZYsk1rYKKy4MW7EtJV
HUsUb+usbUHh+aVPOeeK36Nq3f1U7Re5J4xnL6sXhVFsTiNZ6apwQ3LA87tt3yDX
aJyssVn88vpPJi37JWrazT0gvAXF/GBQVHTu7JIU4W11j8LNAm6oSDQ+0ox2ydkv
6Y1sU7G/Ne4f0CDqv9g5TTMMMV/Y9zyHt4pWA+eM0gdMQEu3ftwqdxExoSoPuscB
LbwM7bcxce7O8FHT9/A2q/40BOWWCIBVdWY9ttjmiJIUoWthm7SW9De2JoWOpMhi
qTO/Lc+0J60OUiZYx8U8x82SUVAswLCm9mgNfLcbMTQAhns6Z2gHNdjRUHerfWoL
sHnMn3XqfxaDqMsvr4lVgeoyaBgAwwX0SDoy7LwPQfYz188aG4jxWsm4D2hEuOfl
GkRGtftjASMkmkc7YVxM0m1VqhOF0yJ2vK4JXrtQIhslwgCWMgz3gpZEepp2j4b0
q6SHadd0V9UZ/yr3+3jDx1aM90ccdgn/faqE4VwUAFsDrd7ht6IOYCi1At0u9mdQ
4eIvocJu77vUYzJys8c+X3m8g1Ee3wjDy28q140FruwmSKsFcmIkYyOERN9Q567r
VB2HIMWwOt9JTdbZuqVhwkVWT+o7q1NRaLp2QubshVUBYcY8J+4vLfeJMZEN3srg
TWcxyDUUDl76G3KUxOHs4PNB8YOM/TCv+d8SbDKt9xkI4h88u38c0jbcn148OJ3U
BfY0+jJRJ+9bL9qFoa7acCNqNO7YpuoetOUYtQzFGCacoAe+deNSbAD5PoIBd3HS
2JoGTGjXMsJaStt0uPFXV3co5ZB92RJq7wJhYFYKM9vHV7VHsGRjxWOYY2xnVSQI
T3qIPynCstfTHoWLHDbVVyenPWiF3zy+jIBA2yPw139kf/KOYh4CXU9dCcvZZLAE
7SshLCq8sXX541lpspXwLyLDzoWOvEr/P1v+iBxtmuB0ax53o0SOBWEn4BqaxuSS
dBxqPhejPnqjZ8vaxEAvEyq+HTVvkbQOhLQEx1Zjk5yzxa6TZ5yi1PVWHCRKoxIb
ZGTdRXXDKXAz3bkU0byNe6fIyRkGdNfANc1P7r187APOgJUQ53u+jZrRycTwbW7+
fvmD/ElIYq91AF6LVtTz/+AhdPnEMtCU0ajZrOJ3/4ftmNRomAk7zJ3L8R87SxcY
Lmf+Fw0t+FAFmMUua9GTvID/PsTsBC3LX6ej08YmQzRIFc3fs/+GxPB//KU1U3lx
Uc3DY2CBR+i16GwQ/IB/Q2MdENKI7imhy+2t8T3d/hNibpuiSLZB2fJJyg+sPLpT
/U9StgWe3ddRbSBsjOnSfbOnYlW9hLLDOn/KaPVUZ+GhrvNQDc9B6cI2HyQhWtYh
XeZw5LeE/737KNYTQoxeaXLtKU/coRqdJViN0W8SStOCS4ty1eRpXwBuRxyASyn/
1kgMNRs20osIaykTRgqAcRQMalTPfXp6DyX67DTPO/zekuY2sT1tTugemiSrZxlS
ar3JIJZ8ax2gSTD97GCF5lX0Z6VgToFphtIcKAFcwdVpc4snAsOv7iM/JHZ8kAPc
8z1jEejLakMZ9lyZSS/BOE/jvIVJuDck464wtzBRljCYocEInDRe0vD0ucQfYoBU
F/5I4SsiHy2fhhtGDUYYkVZL0dmTUdzQrkdfbdulqjbdxgScLoz9tVQQG3nj7s7k
ofzraGDb316MHwum9XcfcjXL8TuGdpFkulTY0ZQdfsW9TzcKlV+FVsqMMCsGgLBC
4FmW8m7eFL+HYP7yxR8rNFl//YXKKdxqXJyimV3zrtU/10gJXMqni+9F7rTXm01g
dQ0yLD2XY4vE1VgeFtlhnUgmQjCrWwYgG+0A/SoXA01tMCI1R071H1DHwXgNeTXW
c07Uw3xpkUZ0jvAnvywiD45yoy8vD07812/Ipp9BQzFFNrDVNuXL8GckGn7/An0J
I2lTPP3FxkrBGYF1ygR7KbQwSrhAAUeECvpoLmnYS0S1onqWTrsOytOjhsklc28x
EIZkqW0qaf45G9XWWwPMwqkOAkChLKfMysi64GCZRRzomHJPOhzhBuBYfzH+VID5
aFlGYAobJ2XCMkYYzb+aveA0hcjhUEEOquhgo/7GkvVQLEfb47I2W0Xztj/OTgEj
mRgWoqgFWqzCmKMZB1A0dxhYZRIShg+EmfpJ9ontHdE0/vym3rRTbyBT4k+Ugy92
nAgkVAB1tX4W3V8dP3oaE7f+pcgWh0pW+wmXbCBbziP2XhkU5+SmWr57Wz3dU3nQ
eDfASB6MyT3EZ2NKx2DvTKPoB1jIJ3K/LrwQOtSy3mrF5VgR6VHsHQHf9HdFH/vH
xnqWS2Rs06CjHWRPlSWYvVzgiyoGgfexcV4LzRAcc4SVIgwJKmAcwFuz4jcjlSEr
/IB7khBEpB/jxzEPHohbLuZR3ETaXlq5GfkD/kvyw+Dddxl0xZW0qnJQC/C6FFPH
Pv3vMfJTMZkh8+nw9O/LVn/Yft1lht3qeW9cGkUM2HR8NZtYEDWZZNWTHgjIatTN
cB3TOWalTsNG9R3Bf/qrHV70hWvNXmhHxUTS3TFSrw83RdiAyY8elR34LQzwXCaj
5xmEqCkFAPhdB9nILtYPEEkHkpCIRol9VOixtotZt90M9ngJmXS4+WwVAHM1zY2u
hQp5dw+rWNQbgpRSNlq9a8YplM2h/ypBk8PW9yuV7e1n0jXdCj4bmhtCScPE7RT7
A5yUCQ0uSfv/mw/lRgq9ANnx+jJlmjH0ud7GwgAsQHtjTYSwSAVeOKwB8ik302Dq
EEdymPjkwb62w871cRYBKR25OLA1hQT2LZjJU5L22QF+fu86VXwsEAV6NXFU9uJ4
H1ddtneWhuFyrH5ZBzAeHH5Dd0ffXj8D8sijbgaTb11s2nVt2hRp+Ry6vOfUMvDv
SNZIHQIGvu8+BVcMI01QUGfi1sUb3GnlwQc+LDSua5BmO7Uv+ssNwsrPX9SpbZ0v
Fk+b1JeyPrg0WwEjFzH5M15ERSCYUzaUEJ5Qu0xF2sVc3wkvqPlgI3V16Df4tTX8
lD/MpzC86p8XglnrnkvtOWR0rCZkhlmVYd5bFInq4uWpcA0SjCjz+NDijmpoQXnT
xBjeBQmzh4g6YaEV1KHlc4yCPl8ZEoTI4J5fKf2dc8G44ZTihU69+I4vojQE/JKo
UN9nhjfWkf/g57szKcec4i4+LMmLdVjGOTBgblZxKlk=
//pragma protect end_data_block
//pragma protect digest_block
wDD4Z8OYEOnKMpjRpEUoXHt543g=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_transaction::post_randomize ();
  int log_base_2_total_bytes;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KI5j7iiiJeHTWrxsJWAM3X1eitOWLQWAmtYroge+fNcMZVVFHGRyreKQTpT0ytpq
6QAzMnSZ7pLfnzVhbnJo/LEzkddj2wT9RsCbp51fqq56vb5D5q5SJDZqSU03mX7N
P1sACC8YXUtwrD40UM/2dp3TxJWU8XXBStMEJ9lG/j0ZtzmunNAcbw==
//pragma protect end_key_block
//pragma protect digest_block
XSGV704FF0VVjar+ucnLp4/5y7Y=
//pragma protect end_digest_block
//pragma protect data_block
I2fGKMmGvelHksAbiGrMI1GepUTkXR0Ak6lPtjfKagA0GEhFhSDSNxiWxPEGsKQn
pfRmPLKEw+WZO8nOajzNtZlvAsDIUnXOPdFAR8lhkjHIfVn/gZsuvKycAqHvGnaZ
5mE3y1J8WDF/+0Ml6uF/zF3Az2zfVaLoRyAfPBNj10qqubHo4mkT0ST20AZFdGi1
itSJvKBdsMMok8kB+iypXIhJRmJiQi+1fXyt3wE6yfEwtUiaFIHZca5lz3FVXoxZ
EzYJEmBPsPtb6QAeSwHFvBEy2nk7ElNdDYEjIlTkDoudYOjUvojkMZ/8CrsE3g27
mSXcSDhDnhS2CvJbb6KhXnThNVaptGEFafYwIYMvj2RjXX9gsX4kwAvHxPR+7c3n
74PVA04AGRw1PDqupoH9DjNxFiTkizWfMAVMJnNlRv1yt0/qV22qE/D8RVCWN1u/
NARfykKnCUcZCAmQZQZnpJxXUG0NWQdtfrdMCD7QJUoB9ekA5/hgtLsv7YBnzC5W
Ns+7pfnjYqKJQCxbYX/tmj44qLIUodYg6cccNkIzERXGepGiOdPOeubTAmfhFc4B
jOyPIIqmneNorHDeCel9GILStoK1zmRFF1EA99BI+DkCjwiAux1mxpsLowy1sMCi
5ofuGlQYO5LY71+GHN8Jr421Vd2TD6p3TXiM0FZ6nBjVqOEma+eZhCiQpBVm9A4e
dFT9eyvgR61wCyRq/brI3xwZB8izGjRNNJLfSAeX6B4HvcTjHG5rEQ37kvjb+2u1
RQTGfqiAoacLSJhuBp/N9DZKsqwWqh6/87FQ+6rB0HJbypVsSztuj/k7r3s4RdAt
J9IJ8itVuAjS1/qFUBcM/MGq+GIRqND28Zngg2hcPP81Cap0lnToA1VduSKZ86mj
uPFAXg8eX5XTQ9VluGJjDSnv/3QuL3awbSpW4JPMNR/hqxwqDcevsEV7nr9SN1ho
q29Q5AJh5z5kW5qKZBvwFW6krynovRfXB4Cg976nRgZNTgTUGDXdGGnIyFMuN2BN
ed/rxZoZwTuXjMPhFhquL/t4qWHdYwpaW07R3Zwgi67mvmZNoBWb2lq/Ewtfbj9H
PXSAvulYnv+XG2J0cRgr+lzum0GEw/kUekjaamMqN2Rhw1wXK3MZoKbgcns+h6+v
TxKqZ5CIUgwfaqwlZ3iFU1mYtm3k2fNz8HcR1QPdc1ppHzzE9RL2vffmbqyEFmL4
F7uA2BnK+wKIkyLOsko19aAb5lidiCtfBe00RoM9cGA+Q6go5Ys0SRRCIpYA6H/1
8h9fmVEISGR1BkY2wSernC2o+1eS4Iz2WUNB9Zst+8PjcMhUCVUoFoWRzVSx+CZU
45ARRN7ltDwX41etl/Rgw/ylI7MKd/7zI2DZC7jMvh1JmP+MvFUoCKvmx+IqUEvq
1dbi2tGHAu6HrjDoukotLaR8xPiu8JJsAV+hh2Si/GUB/U4Uh6sh1QfW0T7d9GNR
ZsWY4AYo+hG42NzplKmRvWTADHGgxgEQSYiePDneIKbnohVOIu+N2uAYjNvyse0D
2PRqRE3NmxDfUwW5TVpYPsm0EaVFerBlcL6whvh2wArnzurCzhBa8mlh0tlwiFKi
c/pQ2ibpwjx/aAnp07rQB6TDgHJgaHqiDkldGMJZ1vG072v289itPu9HGH7olg/G
zvkIimih8AyRcR+9T2+iEJEzlllqYyNx6cErE8WtgMPBaGKVGjPEQPV+rshWjRQj
vPj3Goj/Bd+k6Pp/CmGNLdiqyRE5Z0ovXSB8blPI93dWzCbVizlAnqlCWf1yDtK3
fTBKP9djRdChhk8aBtiehH7+XCr3Sz+Xq0zKYgB3fA0wpXuo5M58yIN+BZst/QLw
feF3z+25erQSjdLvSOvdQX4qkNnbVeoAxekLSl8Yvo/QME6XfM17yRfriqodyCq4
KdQKbQkrocp/OV9Z8TybQrqymv8/RnVgDh8WjtONHfdxA45v70omv3PeBbGXG6Hz
lEhWUJ+Mv285dNtuUqcA4kdRC1+sncKaUfsCny0rFxKZuzk1Ol953eT3tuWV5kkX
wih56385ghiCymU3GAG1+0o/I14SXgB+4I9MMnIcYlVGlQbAdzUzvh5BvwVjpIyB
hGttB9LCtXBCjknss6rAgEKTmRE9MIrcOI6kP8ns5/ED+1VrXOMbWuOrDbTo7SKp
AhJWRn4pFAv1SiBLoERCYlIJxPV9u7VIPQjhxvQrvzltEuqgx6OCnQTYGnbEqwNt
Wo2+CUb3E6QZ+WXbgeCXvHzPpIiLMkpZPhaNJvYResmdfleInyGCGBkIbMbpwh8U
0B36EDYs0jAk3unB62jahZDv2Vtd7con9iVuvWJ7pLlcRo4cHaAH81sMwhBkkgBm
sKRXeeJO9YGhkAkuArFPo+A2rLUd1HDf63sK59qNguzRrXmY8Tjv6INUpXqXjLAT
f9ZGr0uQt9pQD73ag9Stj4786Ry6WExefuUN6lRodVz77kJB8mHH4iJcxQa4rSu2
LJNgHIHVeLTjENV3ad33+P4EUxithyUdqCeR8ANOKitiy/MqXROgytkCad7fUmg3
iyikgbFTOtZ0GpMq1+MVbL5I2PkQsRlJFZvSFjukce/4yJCnuMmXo13Xa3dngTj4
2lc7cMVe9KBb7brnEClLaOQVa7driRTx2ZG+N73GRWV8fkpWt6LRnrlbYCd7cXGu
R8DqzAV6ecX3BCxyvX+ylzzZRwWAG0AqeFViRdW9YWcNKQq0QEr4RHAduNwsJVCj
WiC6dQgwm/aBZXrQ03b/4dRz4lEmSUDprZg+rKO9LxI56swCT5lxwmFu08q8Qs/j
vrEF6vnLKB2Tvz4a9/NB6FmYl6vSd3gCsbWshGzIctRK3Pgvk2Wyhko12jvmpYa0
dh1w58kikY6Vlk0YmZ3u05ecQOHe/dOdDdSLI0Vsen+MN7eXGSDaVwT8Gik2iGvX
8pHQE2JBUN88A/i95a/kT0YiyyGOCia+W7wGGnpHDkyYW7Qcc5qTLq/XTGPuYyWA
FkK2j1D/0YhksEUJTtWsd9dyMmoFMTYeTgqOY34c43Q1YSCFlXrZKnm83/+mIJVw
ohY053iz3cSEfybHkBngnraVTg7suMYcrwbsTC/nCJpPiJ1g91Wn5bd4HmEUbW+a
DsTi0rYelFElNOXUDex6SuJAMP2zHGYranQ0pJl82PGoRGqkvOoUXJ/zNwzbxw7A
04QDmVHrE+1KG061ZYGg3sDCilh9HiBO0FJGhwY38K528mOBsfc6uyTv3ahThX4I
JuL4+4WP1Nn+BfIaw7kMTDPk6xeAkxMbnRZv0vpGYOtwoPWiUMlfbKkEHn9AvX3i
xNB4spiKOq1KVlshN0Yn2fcJjg9uvLCJ7/LhMBYCLK2zMZFi0GZyG4r0HpF3zYjT
utHiTweKwvhXFP5dZltk7VIDFEkHs6fs402xUENZNAkzRdcVtflmgRmcYv7Zr/Y9
Np0X+qATYyxjkcEllRDnQgjoNkeXeaSPXBpoffQgwLYmCqO+lNzQMNiMONleOZkW
G5NHvRtp7SUswQfg6eLSwJLtApvdTZ3Zhic3KEPJ2ddX05gQu/0y0L9lGb5RzYuD
WbIaWar1PS59FTqrpJQOhNgMO3t947wmC/HluC+2f7E9btin+CbO5SzayAmX/OCU
JX+XxejXPc8zk4eYYIzld/94yYDpBALlIWH6nhhND7F7SALDuNs16g6IDoXUzt+a
tWQ1G7Xd1nKhQU03P065rL+KBIO33vNHbRUbIh4RoxE9JJ0GzF6DFrYDBVYqnT/b
11xXOSw/GU4mGpF9EnatvT2zAQmE8mjDEkUdmyhf18ZnUjClZ+7OGuhvGFwvgXBN
KqMWxUoOWTYknBnGmdngm/vgXYD9O3JLYPoyTKABVRpewnQ3sUouPNF5j5kqligQ
ZSkiKib5zOx/AJrxFbG0HKRc0AhWBuMiu/yA8dmyIEiWJrHLRmvD3eGbIaUJRrl/
gLi51wxjBI+bzIbnJ0gLTUCboykPEZ0ZJD8XPj8kqMA9NEINhULr7q6CB686EpFJ
x3K3VcnOoPjeY4z8i1c03jaF+Q/GTmQi1ZhlOARCyfMMbMvi3Hvj1U4SJ2mP+wLA
Lh+ORXAdAVmscf8jyALzG+sqGeNx+6fuMfcGmw0niAYHRiSlFo3Rl7UfkbRE/r+w
gdT7GJckNxOHA/H7P/EerQTtCR/uk7/HZS37R6jOcEAJW9a4wH3xEh1BcjSrlL3b
p29aBqecwkSk2Ktk15elWQ857HBTtxX9CmgA9jlWcZw/f68wZQJfe6jz98IFLf/2
VlcaM0IH+JSd8iGeLEDPQPYCJVMCsN/1NK5ifsFTwIojEOwtF5rQVBPXOK+nW7FH
c2i7RRC+SpNMSsjMch9xdLPL6dVWIwpaHpqgZQjkrK9EfMDPOt4HouszihJDX4hJ
p2UxTeqctF2O9At6DdTB3Hw3bnfRi9UTvJV/aOfS9E2wL7UmkouLzAyBARiXwJYa
pZMiOtMoJPBf8VBBm8Iduw6tsMvSCbax5Z52r09rEhP3eVYM9C/eADOzzwfsEDu+
elIvUI9sBHGmUlcO8VcuPGw+RgB2T4/nBj7XraLdgJPxh8zCymFb602aLfTU7pAe
RbS5esmqJ2+bN/zj3MPuATTxAz3v+8ocprkHYyjaBEH14HmR4xJ9QO5XFxBwq4jx
xTibzE8IFVhLF3PMwaHBunm2tXe7kTEZ9Nj4w58nhEApa2Hb7TnqbGeCIl+Rs5g/
hASmNqfYqRoe4AJ9XnFzRIjsGtkzPkP3Y9lPUxoGsiF0mmZiy8MstymUhsjibNlY
ewTb1sD2vxrHnG4saHv6heDuAzcV5USQClFzEy/Lxa9kmUJIivlQLt4IPOThYOjR
krW48nYWLWz0GvvssA5LneXfAaroqiP1FJeeZk/ZpEFOXVIpf7qt9/ll0oH/Cp0D
guOWKAFbwhPr9rNdTYS+m0TnVAm2lS+kJl2AvsLR7CeYkPK2QalQiuD+AIcOOMbx
8ukmZUc3F1lqhiChC0HWJ2ZWdUYioyxOZrkDWKLsC2CxK8K7Zow0YLyPMEdg3tbQ
Ajsiaa7ZyRf2F6j5fCWOmIczbasDEzPdza5lkPZ9XmaSOdChghIj+7GC2rHDSINr
AmIsr71QzVngi/Cdx8bdv8L3A3LSz/eE8lcExY481SjXxlkucQThPOzAeyG2z8eo
VZUVQLtaaRzurh88nh6o9YtNMD4tPItma5QMD+7+PQ2dOOeRJGc7NpkDNjlXg2lB
kDCtgHmvDSi0DYFJ9KbltuQtBeaYBYST56cL4Hr/ppUi5yRnhlCT6v+7Ly0Dml64
RdfQabDu/vKTICqE3drAMZHSaLMSBu3EZHE3IVX8H/fDvgj90qUDyXh+3x1nkzis
XyKHL209Q7KYikd+iT7mHCgDuC4B+08VZb6apbvx8MO+ho/ebW9diPGAg8eqrtgw
9MWGzXJDZdvlMOasJWi1vliXBM7DHGbmxba00Sv23GXloyalP63GSMq92lQPPmbo
Jy0M9aaZatXZQg4oJOMTI64NpZahY64XZ9Up6jj5zS4bkH8IHxbbltRkJn4IevmZ
7XV6neKwB8qefOIeB9WszW5HhaoQqutzp+uhwtZCtefzpYu8Ah/PzO/bWM2oMWRP
4zfo3w6OIuFze0DpzAJiininVJBVbfzJgvcVnga3m4JQ4671UXcI+8Rnohme2zdv
lllEywbrqZwFWaoe2hyyFE01Mx5QNByjYQMYrh6SopKxfs2MiPz1u5fqLzIma5wq
3inlN4ZG+p6+BSdJsDeu1etkzD1ugsqRkkNru44aINjEWZmOWzsbiZrvHR/K4dyH
bgNW8QskPMgRf8BWLxNOrJkC7AKTYF33AKa6GNOMGcv4URWgQDs2S8tEmKdRCHaf
NQSVW1B5VmXuvHlqj2J66q0Gc50xTvkaglH3O7wFBTF6/MarkPyr9j47UHoK7odC
gHw9h59IXBASuTrr5ihbef/3yTqKDfnMz/Rkb8V1laZqxVe6xyHerDI2yIT2r0yv
eKm/3FQvvLg0gOQ7EKd3DrVzI1n1LNGHjkev5MTOVtizlg2hdZe7tYELbnQjI0Vj
zF34+JnKF+4j5Jl4KBg7Dkf9Sk374Dpgma8R8YqJi6+BAPx5OsUcMVtPNiJmIuZg
x+YtwTRlhke7zWUkFMGEFsaqBdbG021AMx3auOPHyKvu3C3gV/RGTKQ09FGQ9ZnO
/HqOcZBw/9remf2XXDhOEGXmMstfkztnqs4N8quckoO3H5yGgRUJMDHRfPl/js5g
XeZMoDMB23YwudUf8V4JL7AMznVTPbo5cdnhX8VKjFedbd74zWaPwVsKI4gblr1b
LV9n/O4dseSw9PXThwVYOPbGtuz+Gyxv7qjNoobqXLtvPodJxxK3O6Ws2H38jgp3
8SjN1sDohX3sWlq7Ps8ttnjfVfLOQAAJaeMv18gb/jSGyZLwjyDPzRdJAlc3NHTM
ZFuR88+e6nD5pHqk//MAKLqcHPUiNqO4E2ql3TKE6RCfWxg0EBFITYx+w+TqJjV8
8+/9VtH/vtm671eONJNZ3BtlR0inyFQUXB0yTEWOdPxwGY+u5TW026roTZH8S/Sz
n6tau1C1kUsreoBCX3SPW0VkMav41/QHyht/0HQ41ec8MyuWoRegCvTMUkmQOpis
NmR2i1EnqTL5mEqPlaCTzEy0mWF1LoPJ6mk/LWS0UVFiYECECA5ad+HK8KicAMjo
RF7IOpDGFCi8EdpqzhBI9CIsc2TJihdav+7sRU71P+1jOA2imD4m+k4XTOR6zYC3
JrjsbeN9lCMjl/WEdrKk2MLCCRTFEA5D+M78KOim1dEYj3BqAsHGPrcNJJh/z2Z/
4uL82Me4gKtlgM+5LBswiUOaKWLDDq9PT2YdLOWEVUfT5ZvGoadTd6mKo6nidBp+
mpwgmM39Z54G1s23GADNRaZyqxJmZZVZ0fNzjcx36vPi7hSz8wp8az1Sn0lH8Sml
jtahf6R5h5Wuk0HepFJ8MLIkeGofKbCT2CSmrjJeRYeUXcikHcaEzcVRuvmPE8HJ
1urc5qYdafPQFUqhyVBPw+NQipLKtC1seBHCe5HlsPXYZ6UFCk3YDQfkSjOaQJW9
C2gIKPG3d7Vi7XhLmAzVEPRv49y6O/31Djpr0BT7jrZfteLzOjfqBsZ/q56kAZrd
yw5ArdAoIVkpDZvsk3Zsr0COgwtUmfNCLx+7LqmBOMVCm2JqpouAwDvwUU5Kre8P
XG+s+nulfz/SwUFsr7oi4pWfuCN4iyg/FmeHX/YKcoQ4tGTWq2MfAWdLDwkpBvU6
aCqDB+VwOx1VvjfnFYqlgiRkVIuTYV/34707lintpdGcQgWrqG9Anl3tWvX6QsVJ
+S+X5Io4IPfArDwV4gUtGb+AACwdLmIZ1NcB+HqkZ5jkZdTnLRO8BfJzpmkF7u2p
uUR/AVEG3caCSEPUQmPfe2YEb4XWOSW1ZomyzxUuYxdrx1V/iViCKwFOMqbKvftP
kEVZhiuJT9K9aK9ahmBe4qC26oCJfAd1CXPAWXlLXDEHD9w7D44iWTavBN0JtDoa
UehavO7vWl9M5kvKsTtK2RYSP6/vlOqnHDmIOJx7xpljKGdRfSKbxtz2wuN2fg2C
TR7uPQ/fERsbMEXxAq0oStC0GgzArjwzXKNRvrfh9LcQdKq/YMKNOX85CYAf1iDz
kunYM1UPCUA9VqjR1IAZreHB4rjQistr5DwRp5vRGC8wdO88dzmcMgZFFoFFBoGm
vOCdObzPF9UORtsOY3WWLuK5H2b3AucweNOPD31nwVUOdllvZ3wIvZq4RsEsvJWo
r+bVXLtaNs3yHciy6TVErbMgVNuntdH5J7GiGDRjGQLRA5i95MNgVNgIIeqv876d
O7EO9OfX/R5BVibyvcSsvPsbnD4Ndg0LcyktcMq0BNUfAu3H8+YyWw/Zhj6+M7SY
Y6zBeiNKHu+XvcVlUqtQbVmYzPfBMplvkuls6pevESFlFk4Zq/IVd2dOooh7jko/
cXjFQiNe+hTU8g9tJGEvaBS6p3ysAosgsFXBpE4mLWpVH/31cHIUohHXIhW1V6xw
hhzsoNIULRpbWwXRmwhXM2xsTNJXzDC1uzJb7hLdyeHLfZVB3oCr3BceOvEarcpM
pswmPn4TlWfwGWHCcH7Q4JjAnjFM2ctXkfYyrGUqwoKF+kbPzS0KosIYDtgk7Iqv
bZ5H7wyau/cLCCb0uFe9Ktrd7IzzQttNn1QX5uJg44Om5InyLtdXxH48jHoVCZyr
KRG0c+zjVs5RGGYaTgxovEDRajOPvMGXTLt3c6HCtVpmM4T1SQEYI2DDc5HjWbkx
dPdS0Q7MT7P78ye6L4nOstcgz7GWeT6PWHyBOURQs0BweJLbak2U6UwSLmoNbgjE
co3AzG2wfJxZQ39eDfY4wrs/ocknLsKc+vtT7JQ7EEx8K7XdoGOJmsD9M6eTTTYI
TQDwnTL+914TWxG5M22Mq3uvJ+71+yP7SH5C51A3xvaV8ED1SKcfDYBsdQId59rA
0iFGKXtrmkKnglbNSFsSKhBQElkhMnuWCfcvL1+4wQA+6nJk3LOuWHUojt67ioin
dAuOkmDt1Af+46Fv+DukkC3lr5A6/0BpudzMkiY+8u1/MnrgmyQdM+jKL542H7NS
Nu2aUgT4Mx5EQkUGSFGNZv0T/qBSdfSdf82ccvYsDDkr75xa7lqOqTBPOMZtlbm+
67ozU340JHUgsipvoFeTn1q59rw7UobHVorrOIt4+9eHiAZxb2ietNMSOmTuHqTa
Uiz9W0rwPFPvevQdXu0WNiwCxvQ7avZPEvgeRVOnBOgD5jxWUm40CXqcAvSJSrRz
to9l5G/ebvnNGNdjrAW61qxNRUfMIAaX4Uqfsy8p6twDZ6l18XESIYQubqvyNFJP
BK23FbsNG3urX5XgAmg1j6MVPBztFJtQkRrL6oPLpxsrxe/ye3vo67bOjI438S86
PdMEEUvWjRAp0YcF0anonkWoiwBA9MTi0SbqzBJNBrhNcRoPRPAy/EfLBUv0d7Qr
xeZsvHk38qNmX737yStpEKP+BQY6ByPalC3tDtuc92lFxFUM6VWjwILq2XcsiZLJ
CFFob83tL04uMVyRvkZEKR25fSpYaR6kx8t+r8SeTusChDnBHMjbwC4z1ZfXdLPT
Fu5qHc6+RjH1fuoqSq/F1jB0kClZvDeKwQSjJx0SoKgnQcwCcFjI8t1qzqkUqMNw
8GFnguqsvE2nlapoTPvejdzyfMKOftpo3oGlMXVaYYoZrbVQugScGDxfq7oMHhRZ
MUEAuMsyAfzfUhmN6bVwrjplt1ACBIN1Hg8a2mcBbfbCTvjFFfHiELrGopq3CR2+
/UOOV5/3HPFHzUyKNwM9HeiMA+My9JGYCDJ9ern2AjE7U2x0WG04YLm7B8bpDh1V
aXyQ1bYc2JE/UrohD8V0Me0aNDiCK5Dl/JbBYqWPWXeXXMh+ZR+KU2RBFymfnJNH
KK+llw7wCkwZMf89q8gDJLHXaS9yz6ICFdDJYIOhEx076EPQ5ee39ZFNSHGC16kk
0QE6Ioc7aoZiYfGsB8/gORoJzb6dyvUiHpergHRtHzBA0uU5OXXtL7LVN3CFOiuj
hhjUox5qf/9kX/FR+Welt0ECcXJXS2KqidVI+vp+VgLgo+FDRb6p+SlKNGhKYEzo
+cJqOe2xRkeLhAr/DODMl/90qZOTqfTPaz1pislE2XdL4zZs8jwlQBnq58QSrYRj
09eSoiKeU9FYd2VgrfEKJ1N6BcLYSXUmxs8IJiZ55ka2oBecvbAwielTCk9PjQt0
Ln5O2dJUW3gn/4z3Wmg2Xu+NR76So2JghaTnc3ze/n1PDxJgW6Kngk4yxpSK9oC6
z2OI290rkjPBE1CNEwjNL0JZTfXAR9nJ+jQZ1N0IQEoveynJMaKndU9lWrIYoFKq
Y2Wmq0T/1PrLp2UPjo0VpoAYWAr48bB1bHX0OPZTZWTbcyT6CGCP2FXVkj5DWCMQ
l72CGVnZcI3vndaEDun/nLGHzRtqDih0zpDtBSBIuzykLipUt+ZesVSmz+1G1+g/
x4hOqTHXD7y1RYritqZxWIMAP8sv+YTTKq+ubuEdlptV63DB8IGv23P1/a3sMksD
NhtHCdG+K4O4LRz4BNzL6nf+oDYe6o3qCByFtSGUVafBxAPyJdNA/SCI5+chWjUi
fH2iUyJL+Aj6y6reQIpq4SsiFYHR2qsPlQMKAnC3Er5nB33IgFCUNMWB3NdF84cM
MqmlqStTVw2MLXrEw1+d2nFPWyPVt2HWH821ohbvuqw1hrb648Myg78tAEfDCLeM
4RDO1cFKUXvbXnu95vflfr1dWaqx48B8dlaCJuR1n8OnPMgD9qg0EKZtBQDwPorR
3lSNiRJgwAlsFR7JUhHIf3SlKQ2gH4x+x2hOOMtZx9XJoRuinafMNUZI1neR/nFC
wadOS0JdjZrqSu06C5F2fQq5HQWpcQwF13Nh3i7qPSN8r04w2iO4zXbL5peJVoKL
CMgtI91Z/4mWoyfB6xrOq+OdmuYW9aKBqdC4xKJWT4bwmMtMgq2qrwrQiEJgP2Zi
6nZjgH2WTUUi5wMiw8FkqRZSXZT0ddWiRGm/MJ2G9NM49z5jknZtW0yW9MGoMHr2
cF553q6mK8S4rbZWvplVg+U3CSGAyaiPAs3TeQwTktslE2+T8Jw0J92m7s2o67lG
HWhAHKRG8lf9XujGiyhXCTZ6QOj94N9LQGOXj9Ivg0tcuyuKn+cthscslFOf+D13
0lmuh3DOJaFN6yhBGBzhc072IwAMBsdShYwU6yqFmpTQP9fNu+oILFGai4J98ajI
/jyFvH6mlhueGRmhaqEzxiClSZpHSIIvIebVy/faIDODAZWd9pkvAI2AQ68oGGet
o6vHiODMDSvJu+m6aTiq76PukkWdF/WJxBXKAxP1iokErmtuW8bIirbwPNpSpxD3
DaNUuU4I8D5PsmgGe8jnYWYQONIoWP+XddbGjeA4kTXV8nPAiTj6t4JFCNMMcGb/
LTR3bS3joDJEkaJm/ctMjTaO6jBP3W1/tQCdWprUSXGvQ1MEkawWCDXebXpHWVbH
u+495xATwUxZmljZM9AqitatNzZNa0WI+toiUqvHgsjJoOppP1+9dmKdDE9juphT
zhwXAmIybuqBfdwkxP428NfvmQ0TCaRDNQmxKpwC1JErg0TvhdXmfj4jdZ5KcZEq
SfIPya2xFx+Hcdc0beC9rawXrVkeLCvAkJRTVEdxqlGMInCV4KrdlwSZ+a1mGAkZ
RQnOIgfP6Re7MKuQDvLmqJQtqpjXMWaa05aq1VNXGm7UhQRYpvxQVcx3Jit2mXhC
YW/t0OLbr0iVedbn/v7wTv97Y3LdnBDBsQjsWdCiytENooMWcuv4woONR6EmhhML

//pragma protect end_data_block
//pragma protect digest_block
WbwxjgZS3UHHNDXdZL4WyzlL3Wk=
//pragma protect end_digest_block
//pragma protect end_protected
endfunction: post_randomize
  
  //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SWQf4rkLaFPinGmEufHy2V9GrxYaz8ajexvecQ0Zth7eVoAr/nHfrzInwD5hSMsr
9GbmzgWzvJIUCSbwDI0iEN0XHbhR+KB+K2R6shjTOwHZA7Ii1ely2L0ibCU0q/4+
TT+0kVrzuBz+dSj3KwKw8VSeFeOqNcmIfU4L7iYZNL+ci2Wo+c8gfA==
//pragma protect end_key_block
//pragma protect digest_block
gHgiZy10G4xfdN8jW8+YDa9zXDE=
//pragma protect end_digest_block
//pragma protect data_block
P5MuW9+8TqFPeGVppjYG6XhPTbyyowT3/mWSfAdpJlckm+aKX39O1hJvAZZ0cC3g
12oFUxRzt9Kc3shYTkBSz8BusXwkpHRPEz98VwxyNgGVA2PPmSZBBk4Cx6Kdik3s
gSqu+elvAE0LYUcL50hDt4+/HDfT9NsZW5N0HUUBycN2XgGEczBH5cGVsMO+VA3V
i9M+ApfcJHRQGO87Pbhf+Te8D2wGM1bSGCQfgWmuQH1LNhXVAnJHAlb6zJZpkkeV
ChlAgeE1vYCaIQyHfWDixPOBmMIUBQ9a3xcNS+BRzQROPoP/LOqdQBS3fbN7XeVF
/Dld4Ll8DFD+6hL/UmUx2dteFBlJEPyWX2eXkmcXArtCaBcAMPQSKUQpVYYKBCMy
0i9V5P1KAl65lgrC00JE/0dnbdzrSR+hPoAgp7bTq9vjXGHbaAmWfcLpFLr2HYni
h1NDZVsW0TzAmBOj303wPyxDk6EFD6EwMYZDokP5FCOHlwkeFPZF1Wh95B3+eZab
irSOVmAJ9qpFAtwjyEUeMG0wK0G46lo1DnDQbCiLnHdcaLqF+lIaCYRGBtMte48X
gX2+IvUkWEdA5VAEBSWWjVCDEeUgZgpOPoRrWYKJ0G2klrRIL977uf7Hu53eXWDi
pX+TZPhLsVBBV9RVB6q6L8V77D0IDdtaDHOjj5iJBWgAS9zFfFVXOss5ACvmLWhJ
eACtcSVzK1GZNaBNEy6d2l/lJazwm+ujTjn5D1vM2WU9M+q0ZIS9N8D93FCYgZvI
kJj1E2Wl8CZabc3MaChnkLlfVk2euBua7da2C5yAZQzsgV7RdSON+j4w0Gbga7K5
Hbq6fYYpFCmd0JIaL/1ZGaUPsQIbWXKv7YLL5YJk++KF3VcfLCNL1TPClwJIH4Lx
w0Lyx6vAkC7+0o0dFw0n19Qbowkh3Pww+1njQaK3NF8R2PlPI41vo5e1+ztxOeZp
fzRQ9unKlq6ggr14kNYY78lQE8B0cy12PhjXgg5+JK874oc4OJyb14zLmICiQ3yS

//pragma protect end_data_block
//pragma protect digest_block
ja3JmvWHqhq5inIdHye7TVi90KY=
//pragma protect end_digest_block
//pragma protect end_protected
  // -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dsbRxOYjihzXVU3aYGiR2w3GUUrBkfLxrmU4qQH62WP7PEUcJWwyiRrbJPtaozGR
AQFgXClNmubkhMkt95YnMzsKbpQ6P/lZnZcNwvWDtu5pgLSKuzRN1WCSa5adv/rK
X9r178jtHqZvyXzNtuifJY33MaxI6lJ0PnJ0b5CpAfh8CTRtwhm/Ew==
//pragma protect end_key_block
//pragma protect digest_block
vzI4o64gJgVzZ/ccfht8GuZn8BE=
//pragma protect end_digest_block
//pragma protect data_block
u7j21rnLFDZJWOcwzrBDJP9NemoLcg3Pil+RbcsM7D0dJlH1N7accldY9o0T1nlh
jGbi7GPzzNbZzZl5TNXa+2bURkPLkuL0mRfz70PZVFkt31+osuDhyhX0lltRgRI7
azqDAxSxJmPVn0dd72TNmSV7ulDz9NM4R15U4E2w8KnlYZoYfAqtM6UpIydup+0V
WSUsHXx3TjuCgu7zJWRtBu2ahYCRQlssqqFaQnx2vxmQKmcWeuDNcAz80HlvKvRm
VtZoXF2oNsa+dwuJav7GFTpBHAF94T+gZqWAyoIO99mii0eNkVfrY+teHOZQDXRf
yC6gtjoyR1edES6jJdTtz7TjtEsqYsYB3roNtL1wAe6DsilH5qZd45W8pbcHkdx8
zNZr/+r1wvaj7B7ef6q1Fz1YDdWDhRmoLF15L3TN+Tc1WgP5UTqifX+82ujKr4wk
qIiNuMpZXmgs39iK+iJwOdTHtfmPSFIte4RDIthUlys=
//pragma protect end_data_block
//pragma protect digest_block
7xYmPdTAWcGFvPV9l5A0Vm5yMdw=
//pragma protect end_digest_block
//pragma protect end_protected
  //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7+26S2wnogerN9kzCDjAsAWYRAysSA6NOIsAFwk/J/nKAW2vD9XYYcS73IdSunY6
ygFqAMc6MqJUJvOHgT7FE77CMe8voT00BuKITDznGULU5Rkl2Q8dJQNSduqgi1/b
+/iWCqSNg2CtJ+x9s9FXpSgHmA3jaFo0HrinGQWWw9L2Yy8FcxcVuw==
//pragma protect end_key_block
//pragma protect digest_block
aF6HljKqsAO+YjHovqPB5Sc1S3o=
//pragma protect end_digest_block
//pragma protect data_block
7LUV8ZcE1/6rjyXe43K/vxo3S/YkHjERxeGO1anNhy+U22QRWXsHvc5kPPYKvfwA
YToyOnU6UIhaaP9nVp7x0UNvOWhg5kfIVfo4sw+goADC5nwpkXt9r6RQy4qWrm/A
ofwpZosU176T5n5U43gLcdJyGVK8YlA3+J+vtYqrKWPDDXvQEWM4FvxJXi5p7fUh
Wb5ZYBzXwQ8SkCaFOmjs+lQO25LoownSSZtIXjwBAWNQSjUvVYwswoOMY0xEWdUd
pSgOsfUbnbTIK7aRDJPnIpPJs0oNjg4jbrpX4ZJlfOcGE7DazzxAL36U4lij0Vf+
QJ5HvQy22d1eBFV1NQQ06Yv8B1a/gn4kZFoMcLYZe8AyeF5a4w452iLFKpGQSkVT
KzuRjsrZ3i7NNX+KCQp3Uu+qDVn2RC+RMZ1BAeohdkUYwK4lvCgiI4K6D5A/8KCr
tup8JvjRt/IsiRD74EiO8WVjdPx2BJrtP3EmCUxHUGhvfR/ykO+XdzgjcHzIFbig
fZvWfgqlu57gOfmirHf5euTTwvwxnWSuyBBPpF0wgoCdzIiFtx7tO72IuOT223rM
90tEkEUNGsbEvKdjLi3QFhzT+6OwvZOZzlXmHLVh2cAfYIiPENObErtueTS52Il8
DLZQBdD5MGi8v567LJEDJKq3XbqwviSwCm09FYsa9raAp47U0oIWoSwwlQx+guur
cWvlqFGOrrM2kYtHqSpgCQWxu8V43q/hYySCgEyMGtItNDPivSDy1tCSIwR6hJrT
6rAMTwDROOEL9M2ba1SPI8X6VbOfOUEWmTszyJtOBtSh0FVLQIgEpJZTxBPVmoU4
+VrxeVUwlWG2GCdHscdkGH+mzejEDaH2+EoDNuXIiRlQzpQRXF80TIv5CTanZk9b
Jt82sBicNjcyBM0xCtQ939H+NUwPClfVNcmqhwzrY6EyobRagvATQP6vBFvxcPoN
MXU+4ih6XUdVTO8P2bjwxbUHCm7YA/NMSllOHbLppx8MfKPiQKEf+kH7VZZzG2bM
W22K9QA+mNuft4GMOQ82yDrg1V13zsAivCbDNq52uoq/vly3rhSeAgAiwcOx5dcg
Lcg/VZVWYhPUWFwtY28ce2O++WWfTBSLdBRkm3Y2On+NvJRPWvTIADAR8Iwv2OwB
7vER+zHQ0hRUbv3hierBpUj7BAjYAcMoFVC8Qyn8LbnQOGf4JDPDWiw2HmM0I4SZ
LszJ5Y32Vkhc0bnVYVZaHNsBq2ipsMaGkBbPxIzczP/wYRO+/lgPzCTWg1YZ+gME
0ju2e6AEBHy7IfV6j9DMyeSgMfZ8vFE+Yo2ThuFMvipPEFtoaogWveAGLNbqKG23
bKy+b0PezI6NBUH1WK41HukCduqW3fpbNlEQ1WCaDEd36yKumg00q9YEfMeQc//4
SX8DYWYrlSzg4BEzfiuUTgnGKqJXnT74Dt2SKSNb6ILP2QY1wO4R1KnJmdWKBbB2
SaHNb71CYuT+J3ijTezon1cL1MLTqTBG28kUp3aZ4Uc3MJvVq3wX6aGGI8/BF/sF
YQUJv83uYU0IDEjquBA0hGeTVe/GXohqj4FGf3l+diLTg92nCYxwsKy3f8puap81
Zk77/Q/gYI72CmQSi4nptOo94DMXxTHV5pQm9PtDuX3AU6eiCn391jVIGWOPzKLl
vY2N3EGCn5DQkUkUz04xg44J03ie5MkLBiQC9EZr+nghry8IVYueT/oPIO/GxS9G
P3K3/ed+R6/MMnxr+Zd4Hjb/NyxRrnzHTKw5indv66zRASpQrPLT8qGXM6a+cNjv
QhTRyJcFc2pFDu766Sk2f+jlSfC9qNu5MkhyuilwrJopzhzx0TysETEZHo+wIjtN
wJzT0Ur9fIYGlxgpuT/wjqa4Mwrm10MT0d6nBkbcCxEbX2mSWl6/Xta2uIeGPLYq
oLj9QeLyT4xsrHcHAtREcKggxKfA/a45Jvoye1vzQD4tsC0wM3BszMxJKOekEXjP
IrJa1cppTdltcQnCaD/4/GXCjFciiyE4jzG4JMUuyjb5KS6B9iUpkzzTjnPqa6lf
+tM0jP8gL84yYeLinSyR7TiUi6u83JRGGcffYLJI922FQ20GPaSyYntfPj1MHaev
pwPOIIm4HOGkdN4stMrgaVZokejqZJF2NhKadojK++AXzUBqCo1uwKCGf97KXZKF
hoaouKze1A09kQakuiPZB/jc5IS4yGfITci86QhzFsg2vY6RBDoLKb9rBk2TMI3N
FzxRAwpHYWeZ6bk3x9K1v5AdOiOwM/cdVfzHjHlC2wldvtkheDfP9ds1NIdP73lV
jldRjw2K1edBmNtZkMOiJ/XYkkEQXpODxGLFYVrmYtTn91LgDl368LC9yssyRwBI
GWc+H8zW9qO2tJB3HrVd3p0IRENInesMm+aBk7Y+aPG8yh83aiO4P2jMWNHWyL2c
+2N28+CaIXEboPhs+1mitjQDwHUE5xYv6odUxnPzbXiKo1ButaXQ7pT7CoZUGRLq
KxIHCgzpcHv11FShqx+o9A90BrRl+m2Saxu5zwQ8yIBqKoYo2YU3oDC4RD8SPYIW
fum/pWvH/tW8fV907v0V6GBIAYQFxXPhOnd3jSAQMo1xDRWAxoMao+4KB67fm6z7
2zgFkS0NpLITn3shwJQCRbpI2jt3PV3O4BBGKXtOhRJ0Z7FEWWOnwHGfjXi2nY0z
gqQ0T5q3XXr729QHo6CBZ+B2eHXXl2jPeEMcAazpILr5zI/mMSVvDwmkOkZ+PR3X
G78ynJkY4VtcmBeKNO/Q49Dl2surJxJQqbO/DCWEopYyGz6Hm+UqTKk2r3EJehgT
JyXBxSjM7Bxo2LkE6GxG3YX9CMq04lTDzdm5EwYaOJ8WzKfPTiq4P6RbJZTHPujp
WzGn8WLsCSsyzs4zuOGYfqHA4SvxBCjL922W1AlZ6eWqqM6tlde8PacJiiMujuld
51LtY93x4ko1JthdW5YsyiPnNTPKh+B9dKWWHdS20cSqu0phFworzlkSf2D25+xt
3hlq9maTzckPfXSYwLTgaWxV83buWQpI/OdAj/J4U/kRQ7+9DYLeN7505zZSZPkF
JGFlLBfRhqh/gQkRT0t/naWPCFRJhbiX7Zuzi6SDBXdZ7AJWrxoccWmY7YFRR0on
jwKbEbqNq0vM4tb01HpudM8emND67Ui7vdlmm5yIQSdN4phxB7yPzS5q2fC2+0Jn
G8ADjV3fn05nmZaywFee1NFgoTfXtYsNx9w03WUunVsAwy6fpIgW7nOdzQqdhx7D
moA1YsjdqGMQ9A60b3QUFcPT2izSeeCMT086jVvi/2F15MYBn2AIf2rx7uuvxYs5
ORw2Ys5QiwGKR90a1BxkrzwX3EgkjFsLXFsLZRcvbuSXSQdR2VWr1UwED67rsjzC
0hrsTkXYcR/eQmaLdoBoOxLKm3G44+Sw44G9VDxvlO8Cz9PMT+i87Fxiu/aB22de
cyllxgxVHMohVsyAa/JMCFzdELmr3fqEIzGcIe3Swq4gytQeK1j1Jeje0GmH93pP
Opw9GnxnPUJK1DNrw1ejHG5LzTTKV6sHJtpgOK9TKyBI+ZDBBSOtreefI1Y3JR6u
q3bWuY4yB/zZkzD3vNEP2dFGELkGU4Iq3RR7l2L0dlsuhTtX85zsEHxOCbcRA1OZ
LDnVL2ll+adjWtbaOYOsiEAgUKriqmHsfn5hoWygHLCTW1kXp15hATgUbfA4kKXS
9hsOtXb5+sn5mHqrZhsYymE0iRZiEOwccLoMKI6cJs79xEa98A41kzsFzqMkN4hj
yjaYO5/Jgq7SPmkhd4S5tJLTKNWtHP7OAoasRqDSKB6Wd54eoE6gBsnvZjNsfOmW
k28oEiNZiVpkS5Vt+t6isfEENjYBpGnmOcveCInzf3+5eBGZXXeUMHYqVwvaACQu
5NqCp09D0Z9Fv2PoKsLN0fkG1GvwQ7qlWDltUfIZqeTsai+t8x5uDdm1slSKgmV+
M5qBv2/rXL9LApxSW1PJR/geljg3buRJvGJOgDSpGuf5Uj/u3GHmwvrGLiBOHAgX
KYPniDtLtS+1FMkaLIrnvYjV2MXzxir10Kb4q0dMFvMaAaKLswf3fDFREdoHo4Y4
xQb0DABRUtfHA2BmAOGsnZ9bO77ObpWNAlwziwz1bSf54Qw6E2DSrm+5kjOznyPo
cUIPJKA3+IEg8lK+T5/4lqC9dHZoD5Z12fdCDggVrv6EW5OJDbkhncD98j54Ro+e
56t8LGiYCYfaLY8hgL9IO37aJfLT+PLVIt2nuCzrzknOpfR5NWT48WaCWo0kGm8R
UdzS03wsnZ/8sHu3ezhH91UpCTjUq898h3sz8Uc+ufIrSqoMZvQzFGI6VcRqDYht
fDG1vXE12mmHd795SKD3cSY+OaLP0+/xea/+XbUb0Lkz/0yL1GLQHeYTs/FcH62C
Vfs1E/xWxrRsRTrXymoeCHW0OFPQOvRPP0VH564Ca0Xmww/chIRGCmODLQQNZKoo
YjG1Xr334oRHvJ2n2GWdDIKugeNX52AuyXvOvjBiVL8E16EXtSPRyiL7VMdcbP0f
tVNwNwjb5oMfIJPP2rscyVsc0vRvzxnrjnqGVzLUIGly0m+mMdYD0WrEM2cM0ZYM
LRG/W9fVgYSufYQJPuaZ2tTkifqX5RR5/aVZSF0PToO+lUTDXpFma+4oEujymPTi
mPCRsiNE82klMvyO6zMDBOAV6N+ETVPcr9GdE3rWJG5JTOmE2pFGRlqa9Utxitwg
qiWB4VEZ83d3Q2Ghnejwt6Cv2CBCFJog4OVus1jYfJ5u04agsOnET2M9IAy0mkFp
2+oM4kBZX/fjc+0moL1efs7i7Etpcl3NoyaNZDOr7L2rfU7MjsTow07TZ6z/jV1d
Q/34lQaFrw84AJjcdHQ7alY5UYbvevgW2SPWvljwuLvU14c4IuD2nXPklG7C4YOV
ohycBUuj8OeNYXwaWTZUeYkVUK5GqbjLEiXMnBvcflUZOLeYsmBBxHUQJvP+HPjX
CzacSl7t1uw2jMuHNp0ujJAbrmghzyMij2wDoFbow5VyoBus1jmm+mWwUpfCO034
zWD2Re8kDy2Qnnh2MQ/oQ7G7rJcYTwbMhp/gSXbHpA96PxCdK6fcwkWQ6n064suP
sThYYlhERx75IcmWva8UhGZzLQCz8oRFbUArJPagwsuEC+Z+4lcWnjJS4G51AZus
8MoWNlicZBBb+nG0LzugiaObzxk03dJ5UTfQ/eR/zmBstqQdyEZk1SEbeASmWffx
jVZJm4ZUQicmgFjClHWZeIp8qBmJk5wef2WeFI0O2knzCpkx5iMKUFE9kjJd/a8z
50t+CEousA7CJSY2GAXO2SsEzW43TcxzzzWLZiZ2ihmLlz5pm4nb2pMpNNp+LdRP
hnTrpV3fX0m7G3JvEE2ABxk2QzKs1u5JDc7c5zr+f9zmJ5aFGjI8DRs2BXUXBwHZ
14vU6CBW2LWQykDipO1n2GNALB5eEVuIHp9wOeRt2z2z/wxpxpxv+SRPg4iWPqlc
C/YxS+3SySHPtKGWVEsFm+sYJXENdYTrq0GnnojoCuoDOf/j69J92vyGlYET13hh
sTH0QfZZ7H2Zb18Ql8Xwdv279gf8yaC9GOcisivWuhApq+BUm7rs73rUw9OIbN8X
GhznCvwt4AA8VriSlmOjyE8hcNfBV5tjtjwF/i8cjRv2ecmJsYGOcKafQGI/m2LJ
hbVUJej+G3JV99fhqh5VbwHxOKtr4uZytlbElx31ljyCC2xnSkz5CUW/x6Z8wVzU
mWhPukXoVF+s/dbNeNFVYl8OxSx4tZr1sbOGFcCjGDNFryrh5J1eT5FPNF7Vmmji
cF+KIWzhlkwT4Cma3UsGydqwg5MSPqlWEw9Ej6iDjJTlrQEnEJAg/h00ow60hbHt
x7NMWDHEuoNzsVWjpdb1RM0gxWEoQZ89TJT1ITq1XoA20AZWL5Ff2H7SNWktfJj8
LblF58AYSJLBtA2RjRPRJs3iC3zmYhbyB6jMecnkXOk+bKECxP8nyv5K7ze4LY5x
nNg4taUptKd9ldJd/798s8U1sOstYoFQ6iAzZuHCQ4FWscv36YIJp9VVU75mjtyH
5UlJP1Zo6pJ7ENZktUEF8UVvSsrvK9uf0dV85azkmWhHm1McmXZK+6+vMqOOswe5
C/mYENWaixMOWYanBFogSqu04N8Ty2uoCi4Rsp9EQUFqoKArQo9orumqCPmaOCaD
8eN4Q2t0HnJQDQspcHJ2s2WD4DpiekoIEeSoC4z4qNGOVOqxXHGKVYiBMn93r6ka
00qVxhSvkjkE6A4vO/ZaufHrt8ThOA+ZWnRtk2dM+l2DjbmTKlFGf03L/yT6H+M2
Krar08fX/smHCtUpERdadGNOfE5AEPJCzq0V/TpQVZ31w/M+yBFsgCpL2ds6JZ45
PuuKR8ioqGL3V3DjY6VpMKW1LMPOm4DWHgOY0XiEh9OOer9WuPsj1Jnl76APgJi9
Ryn1vVpTp4QG0Q/8yZQNyCfyV5Z6WyPGE0AISjLlgkP35B61KK/SPwj4AEVRZKi6
XokpoH12B0/JuxsN1BTt0n2pwnL8GpY18pTH38tsf+iDh0YdDldiJvQV5yj0S3+C
3BCiIb53Ry6b3VZ7UnxIhKK6eO+Zx2eiPUiLxYQZ4nywfKoWSX90WZ7AR9imA6WK
DsSA0eYDzQgxkxaelfA9JPWrGef1W+JLNeRMiiEPUMJDYIK/oCzcrFCH1GHy1voY
lZDSEgN9iD5J76daCSb5jzpTqedH/bXjwZ69iCl1pUPVFh8gxtcsxJUGJtuq2bEE
L2md45Ne77KgzUY+7mn1EUyy6ISH8oeXLkzcSJnhPSkrZULPVczae3HKbkhtwH6J
46wovOMea0JQZuLOuzaWRujBzyne0U3xmQiiIpP2aAAGFQAwcsIi5YrFm8QhlBMT
pVl8hGNr5m0Rkn8d4MTq+rcXTxVDauZsYTTuQrw9QCYYgexvL5Sllce44PvnQE0O
Uyq/ucftQ+rbbdk11/UNsiQhQTt/4bxLPQ/c6kdKzUGZdAfBT+eEgqOV6aC/RYcO
K3MtGNhiEdLSvzWRZ0tAOldXhQZHxiXlxZyYlJZAbpW2MLPzmDfxqHCs+1SOuIK7
3j6k/7gSWda+i3vVtmBgRYe0q5XYEEI1RMCIgphPhE8Pj4VnhqY6HPhZzLrol+r1
WpayEfPy/GLE6yannf/A1+kDqJ+ZCkxcn4M2rkbWUbukWcOFFjYuCvBq1Qld6enU
B83ja+L33breN6o5178jCt+ThO2ULDZbBorK3Qu6AuRv5GLVq8R16yvgyuGGJGsd
7JCGANVlEjihfaY0wi/VjSI+YyxbZe5mvX5nSH7GZ7QRjjxX+6/ZtZgmmfm5VkdR
oiMCNmt+LDqGigISczrx3Vp3wnNU494IXzv8kp4wZZ2l68gl82U0vSn3U80euRnC
SiP3X9pWuaVcY94Hj6Mir7qZLIZIDSbqmTQSoM2pGnxSPAUAaOtOT9eXgexMaDLw
kFXjVg2V+cPTVpaJRjC1eiT08UHf1Q8rN26w/b5BSNSmt+v392MiF4BooGZNeQkd
rIDTP2JK2LdaTnqXfOsGg8tUP2xy1zhEK+NOBY7GKdlD6RDKK4pVj1Abba527l6m
TewGsErAyULyiDuGMpIh7cIiY1HrmYQNLesgIqZDzGqlBhut0n1huSeCyYTfqhfm
iVeZwSAHNAspqkjHKqZhiylRBRaHuE8xRsS8mzpQE7XYhIhANv6mVZUWOuflEAlW
SQdOTf/agwpXoTDvz/0SCoR8rZFcZeehpDdks33Dl8PTq+4eyy06WoM7U69W7oVJ
qahSToJptTejqbPRK0vqlliDkAIWWXfap4OuI3I+Mcq3eTMCkc3XpYxN4CuAdbUY
UCBDHv6k3tF6wPPQYrxErftxG2YE6gqyPCXz90/3JmYw+wggb1iNr8l0TRBI6Pco
1XGWFfIgs7IXKob9ZigOVJhjxitExBx9ArqPGW6jpHS5AK8axWE9HKmGWeR8Tthg
LYxcZ+1BNEk74a9TatbU6RR4aheL281inFlyya27Q0LUbDdRPectTVnOJ6S0Qd+p
+RH4ssT3z6L54H5X0X4t4+v1VrIQ2zmLJS30566qthFS7nFOSBgm8lneeW+iqPfp
T1qQjdqtCA/o3GNsXV8AmQ+eMcK2xYgoYP5ozzaOAIHhY96wmFxj2ET9lmPr51Ia
JVkJbwrwfw6+6wlNvxyWKqwr/dKgUuGPKUvNUa2FyGjZGz00Is5KiU9MafpnUp/y
r+E3/ljROWEyeZypUJkPXyUuIBk/9+/X0phNCy3S9yPdGXCMymOKYY0ItTrhV5dW
UEaK8GX3DGyaBj33skQdX+ms12m52+b5SP9F/zoWXqgTvgKq28H48aYrS7B2s6/c
NWm/t+OMKQR5twnqT1v5w4yXtKPSxk7Bn44HaFbwnKo/Fda6Tohevq5RhCgPGqyi
+AjbGUnrRdFgmkcSFVkSz9PJABSxlpWCZni7NH234942DFcsn3XdjupVWC0Zqv8J
Oi4UUyYQ7qKYaIGSZio3ZVDCpCFEEfl6n2XquCVZmOyixLP4/kTkMw4HTlDxvRqf
BIuJWQ9TBwjUKS9zB3QYdjcuZzS/yEpPmaiLJcNC6vvDaLI8pUwABbZtU0EfIHEu
GaYidGt9RKJ+1bjFbgPuhW/kU0raniTC7xRjXBYGcyxEytEdw7+BtIKTZQZWJQL7
TO4hoToTrRQkDduW1EoSWtioNDfpFgQq/xliFkA9FJ455KZv/cJnGCl6DZepmse3
bzn8+IZe1BU4HkVNk/qT7jAGhm8/HpoNXPqOBm9Q3ZaAuVmhi9lgI1NiSrqon9R4
1SMBbuOV+QKWGoxIPF0KjW5Ogfzz0iAgc2+7DNiyce0WfQ0gmpxofYP1xTdCMf5e
79uICigqOD3XLyTAU0qjfJiEmNBHr0QimqAq3QYlP2996SmJd+FrUouaSNUwEznY
wMwvNf+KeFOHBna/oRaIloXt4ARm0rRvsFz3RFQfZAUVZWXCiEaFasdkYvwHJPvT
Jn6Pbc1FTaFfMGe3aKquFdVV0wuDQhP55GxzeGVpSdl2sIDGlDmzirpXWP8jaQRk
BlwQPNi84mOuFwqwyw53gEwzfVgcQmi+2flExTfA0jTcnXtUjkgsA3Wrqvhykkb6
mia5+rVz8LYjlAs1HYutFEGjpd7YFE+bmWHqzlOevxAQ2uGkOYNoeBD0yN0CZ7in
UPryU8u3qCCxS2Ii6uOCQB3CCKQfpXZ2sIO/wzAfwz+iQMh/3Tmm3+A9umgq8nsQ
sP37w/nSvmdFeRzFCkttX8/k2+qLeCI3EOm7iHhyFXPHkBFuxG9SAf+PRpa7rtAa
l0CKoNn1cCflRgysfmMQv8buHdaQUF0ZjdvgH+5OXuhlp5mWXG11fUTzLPqp6Atk
icnaWheWJn1mmIMhBjJ+qVQFuxb/12XIyD8Rp9mXFFnBGASSU9st050NmwlkV+DC
wsIv0EQ3wy7ESajfQyki95+/mAUPyVC7t0el1yogYOejkr6AmGG0q8WTyeAVOfUi
nu5dH71eTXW+XRQ9IN2imf9h2N6OY7xmCrTuooa9k4YZlU9rUDQ/3ju5ELy/DC+T
I7ka0jeG6olu1qnsbOmRd7fDCDpoHnTho2HCSN6o4trnC8M/OiCz5mbwrNPN8L8R
COo0t74LRMtbfxTJH3SPMLUnVD7ujObjLBpN/I+NW4VH/2eSbpFz7EXBMy403Q91
Q0Rlp8UqcGvG7oQR8o+xDYEUG1wzVkyNisa9UKnlSleRBAfiz8Du6zAzdOGkZWqr
Xh9f59lFnzB3tvgqn1V4y7XUg8HJdk4SfQY/A5YRk0p2bMjGKM9roxxnesnxvBw9
zimj28FUuHA+nbIbsA9QrRDDAL68TVIy04lpFtegKLZ8fr7urMZpgIIGzEK5kjh4
D+3KEb/tAaedFaE6faWCwAVq7FBVOWu7POCJDL0DTRuca+ihmw1krZRqkHJIDGoF
PWwYt1+WCJlJTdw7IQJdPaXObG1O8vj/dspAuTzm+aWyPAMqWaEtpt3Y+s9tZoHI
XZoLkUVhTbVZ3cpxTWUpE8kcTHs4cccMAPpvcRyVPGTWemwcOaEOo2TJyk/eLLQ/
dDNYwcQ5TJf5v3ijLJkYHe1i2YiJMUWoNwQGwJJ9TYmpQcLCewKRAyWNclwfrxv7
UJNlYQi+Qme0rrvldyWkSFJh1sS+oELbiPUpk2ZwWgIGuhtjfxmW3C/9S4PagdVl
YZAUZhBvFTqXleUFxVq9t+Rkaw/AaYFyeKipSRPYM+Gt74pVwI1jHkvRUjzIDrKS
hIay+bSF5qHbMk/GHAsF8y8L1HH6qDEpGMRxrRHI87ee7FzqaJMVRftmRQp+Dkg+
gOXUhegq3bUz/zfjXCLdXi0M2S5G4m67j6vjYIXPgMf++YNko1d8GX2N7E/ZrXTY
0VpvX7gPs+lIfDyR139o0arkXCWSdZWANB/8gW8bdnyqrovmmqrsBs7TtxIEjBCj
8b855u6a1RIfbblXyhpYn8Hgt8PP8sTffOWcEe5veeX5qqPGAOTUpH02u4qlsVY1
ukzg0PkvfQApVjqLBzBHolxCaDQ45y7uW322PIzlW4wyhP4G9VHDnF8uOl3HlnPW
3FGBgLcSXmnGz8m6hdDrpkbRm60wctb/3kslUh0H+Nnstq4l8nvH2HpkoLWkUbUJ
62LC8SigLJKv8AGvbxbRx5aAQhn1GrAmrWT8BUwTImGSgE/0R48JZaqb/7v2tttK
D9rEyIEpWAVlP83r/dCbxxuk8mK7e34AlXnsXaxkccyYWIours64wv30D/+yIpJk
aJzlw1dBBqC7ZsrjPuJOT9go9ntIaVZKLHFV6Qi2kkrPNwS89DXM7Dlf/W3Y0XAR
wwhwHrEEfZ7Q41OzlJCbpkDAbnIo0XhboRcVnf93SBPvDlMS+wxRulnBP0jTlou+
H14/4C9YdPde8q2PwTra8NtSQWa5ZXVvigs7SEHRvujayjkEK1bMpnfnhrVpOikD
Amh82624zhNauY7rfeL4/AkJlQG9B33+J7MyrzMkV/+czMZfEtsuVavmxNSPO/le
cMoA7pmxHzyxQ08zSMg/wIcBOwWcnJUGj2wr3Be9MXz8NJm/hFDzG9ivyXrvlwZw
6mRNHuOTquYhUqcWvusxhcTxxcsmmvQ508+BjK/wg3g0aDUNf1MGvE3C/SCxqdss
AS8PsEG9i9mgqx8NMOr/CaIdM89I9aRfLtD36iPsSJuiX0DQLKqq1wTKmbvpI+Cu
XJRzQdYZhF58ufaGVfOvsxebdmQ5pPPFAhXRYMitCl5ZU19VgSlkd2Bcb9onEcBH
KPZ6OdRiT/C+N1SQcRnkuDrNOEFnODHP8ZeMkclxGC65zIXDLP0P4KuAtLN+a+vk
coP8qHTdVI/eiGpBpqP4AdorWIRRsPaN+LBCiL8S9B1dRBbyZleYu+8A/+rZCVoX
1bi5xG2FlTk+pm7qTJ/F5NTEU1pLmX4Scyl3sTYyfSMETcBCY8KLhrCedaLABIkQ
FKH1ucXEKDh7092azLPzJm8tzDSH+VDmuzPtv2hb5Ct73G9hQC3Kj1DxEO18xClw
L7cBRUkpnyABzV5SF+icKD66acK9b3pCSAymapElE98+FpjMlpJ8Wi51DebW5pSx
u4asXZaDPrtJsYCCB6E9hrANeAy9c3bL5WIjS5CHjv2UEwtI3ucN5VaHWoGv+RoO
ic+ONL9eaol166KK9RBsuanzGy+ngLq2fZqGQQUbXfsdAAT2cMZ1XaXnlHl1LjeQ
FgwPV/wRIQAsAcyhIbjj5bGUzoLGH6JzDVzfrZC8nnliOJR9tAChPuifGVqyqD9D
Lj5nZsBbb8p3ny4HNii73xexA2qKaaXV5/bnca+4/NentKJHLPGuO2rPrvE5M/c9
X4nckM10jnnepG3upswYuNsCmylPVzIG+3BnsvX3hgo3Z9WtX1gLA7Dwf/z9EzqS
nau8kB/y1g0Fn3iPyP92RRDvJ4v73ERDO77ep6lTlBK1E/ragSPhsAj6hjR8FpCb
fpOZHp6RBPdawwyP9HobuBXC35sdwDzE8BPQtwnc/dLfOETnRD3ByX0gGSXLU72h
haRZoYEpt1320ZANdea3ls31QWrhc4UuCLHDNTQ42jkSRpj2+vEbmwqC+fZM1Clb
YKPITA7CAB0XhNckH2O3/QeJB95qhTVZGHJ5GLnF6Oy9ztfG/XnkEZ2t9GtNh4Ot
FGmQpO5yahw6S/YOlqpSMR8kE/LwA3H43cs+Iirgru24BYnZsUe/eIhb8Dfyb59b
4PNL2DHGfs9mDNj1rLwnRHB+IkW3dqojCQMRqaKuLBL8QFUhOde98KireNE9EJHJ
4LtHUUk3D5hzHk+OydqJaLZy+Pm05aGy8Sv+NswWKZUcC1oe6GDYx7Amvjq+pi+Z
38albmK4+aQ5+aN+ZW5+bBuxKLdOmFA9q3S7TsqcpaItmLL+XBNWpe/gkIjn5bJ/
lm9I9N5Fy7xU+LNyxHtBnzRyiZ+6lMKr8t5xakwz9iJXq9vCjQhiOANPRJuKJLvc
NVWdjg3Q1lXMLEzEMqjnM5PZUC0bO7P6sGvK0vS+51RhdsALlgV8WM4HdY4rqkbY
lpcZqsf1IGYpNYYE17cZpWY2xIAXjHUkXA5tNajx457ccUULghHX5ZtUqsh+vkPz
QLU6aGF9p6EfVO3BLPs6HodA1Z54LZ77AAQfB9D8U5pXnMwDwccLk/NouaRPvo4T
5tinPrPA3NhH+J+1DxHvY7Ala/5VmbKqHOBGWE3FP4kmX7HEyQxcwGrnsX1Nckz2
RiWqDuhdeVEnxGAtENKi+mH7plnlL7zuI35EosbOnHwx6AtqE8/voTM0hPeJKEoN
t5jXELlMc5OzN9oO/N9i/gWJSWxRFNwhGOVy1Gdzt1KLAxhFuykUnk3wWj38AxXF
QNSN3mK4/tvRLY72vfGWCmTJ2kPcnz1Juls08iJPyAX8WSSYER/XJ3cOi8VrwtIM
mZsS4XzdASJ7AYBVPQxzzlrfbeyI0j3ajRzFbeoSpOOUhDH5xN0hwaQ6GNFXbnu7
ErW95GuGmGFIthZrtxqPl4tqekDVp7Vq0fWNwM8tCEBN2Qp8jjKV6APCLWMXB8td
QhH+4zPsjn+FZLx5LRK0bji5VmqNPFj+El2DBzuiZft24szxmeXkM4a2u8rCuSe7
OWAjiQtspMUhvLvjiZHCcESz2DqPKCre9Vd5vvqebL2vF51myn1j+HJb70WBLY+I
1OwPdcN/0XkeUj6HXem3TjapUNYTL4AxTmQhAs26fYLjF+2c53iuGs/cs5TpAa4U
jjYhXrBjoHVIWfQgqNDnfsfZmSHCtUeHuledTn9Xz4sOY7YttkwoNEIJ5vLV73vf
to6ApDNd8GYNLqXvcQvN0LNtcUbeoNuaLgeLQckWECAgGe/7L/hUp1l67SbUQpGu
UmXJ155QWkUjOyZpm/UpPv1tga7NqEPqxkcnPLfH0dQKYTzuzbNfNb7wh5QG6USC
iKDUwVzMT/6ntk/2NO7Va6BPicgByTX3LMabc6r7yfWqp310yBLEP3WSm0T27M/y
5sjVzF+1HE3ufgl53IwBGQ1KXwNeO1Qr1a5RCtJ/tlPiw4cScXyEfsLoKCxFApDs
1qjZI11B1JimurMwJLLw6ERm0xPeVay5gj5hkBtNJjwd0jaEHIM0C2t7/uUQkxGo
Vh6au+8uWuZLbhtw6HoPc7dx90BHl9pG5OpFRDhdwnL6JL0b9Mbbjbtlra6VJj5c
I+VSxmZ+AlWWWQPskENWn/4byhM+WNentL6KRIjl8D2ZObB8vfzJx4few0/HioQY
IwBV0onXibB7udcGfTp7kgVPL00E5ys1UZopBaMQzMivLEAuboyKYd5NEt1lhna0
rnk4kZl2bmyNGuu6kiJBB5N3UfheQJbnnPiXPhTFTnHNpcZou5vmCKm9ZEPIPTsI
SUw4CYyxOem21EBMYSlJWh9lR6Re3pnk9nAp+2pRue8eo/fvhTR2ygc9j/xJs/08
k1bgQtyiu0+cMiTSxCS0ns2zETVLhEFitEN1kHcr6j/bSsE2c6thiFjrnTKgmUCs
q/auDq2cRaopwAodye8r/jiXVAOoVxcWIjU2UtC0DW2qzKHvE5xcYeAEXmLQs/fP
hozxz0z5NtYZTu7BKmcCx8ScZX8XuBFcRwjLxmAreRoe+yDCWmYcQPd15x2Zc1d9
atZ2fUUC3vz5fOJty3rTzCyVlPDOBKgXOr/4Tb5sxEtDsp2Q9BdEr9RyG6XKdcYn
d3TRHLl1pAAUStYj9LKn3tZDT5jKDWhPuPD7zVAkHvSc7I2eM6YWRSDa3da5qluf
u3T1ppxT5z0U8RhtfybaGxrhr8M+0B0f97lSyo7zyBM5EDY1snMYz87Zq5FfjTpm
iezXMG1rUACegZ5nvT8tfkKV+FgEFVqn15zvDi+6itEmxELr+K9NrJoOIvsy7OEQ
VcYEVP27z1kLll4eGinSqLH3imZYyoA9Z3/c02Jt4b0C0//daBYW0D1iBsOWFZ/z
wayK2O3RMY9/foAITe0uaqJE6xQ1PDSl/HQp8ScF1U74Ztyv9eUB38l9MMKLzip5
ds5vM65TzO7ZVcP65aHhu196NSJcl7MPhRzaDW3Vydt/nr0+JqB6+wScZDSZrkQH
unj+2OZ5dNV10hDeWyfO6oPPeZ4y57hqRi0VlwRMMxJYFvnSH/fuTb89F5Y09GIa
75hCgjv8hwIoKSSdSUPZWqw6NyiQpa7BzMUnWHgmAKtSYdLScrVavAinoeUKrMBl
mHedDNlJ2V7/ErTvP4fytugNpIYM10Lyc+ciUdFHdWp6jNAxCV7WWagBXAcpOl4I
xMD8fVYvo/tpCsSuvupOrmGlj2y+mGKXWMUexoc90HoS7lmgXlKE0ziKX4Mob3lq
rm/SQ+w/hoa2hPKKvozIQpSxalEZT7760gVpVUcC46NX0ySHe1mZiE1MkWYek94v
XCriONKnC3MYxndmqr3ToKe+YDVIrATSsWxLvwm2M2QgRKPNtcYWMqDH9sGOntna
rWSdjymaj+FoGLL85T/c/7XTF17CaDjaTibQaeMGX7h2qSULDu+MCSlb43iy/uKl
jsHDmETl+y8o9TcePPthEjv3OiyOpcA9vlZ9lwvG+5jWXIkNqoT3iFYmBxnIQ3Pt
KN9hYjj6jtSmGM2jCjCHXjvY5lQYiRO3UVjUDAMQl5PTWEp7eoMRXMFGdZLCdq3S
12DmxzjHLeRsF0sk0jN7sPsfeOxIcGM/CrmNSAVL+4BJIcIJyiIshEL9l9FB+U8w
+3iDyJ3rt88Ku3iDfh7pzsRVzXg3St+oRPJsHDXu3YVTKkN2XAdeETrNaktyBovb
ia6E9PGBjKOmZqhvHHeW+WDb3y8G95FCu48F52sFxlYtItdiak8r3H6y2myXR6tD
pkvuSwgRNC0cZUH9qhJ7lNEa6+GEW7EUvG2oTiHgV9mNfLK9xcH4pMPvHXseN8pl
v0OYGoaD7TGZd334X/Rk2vclD79gL9E9oQV3cRXcJZ8YjEynYWXNhuzsinYKoyCQ
Kgy+s6NiG+2WvjfeOwVtG3AuoNfX6S43gbGYBdvWq5vsrpyttJU5QokxVGxk+THz
Yk1XevgPwUPGSxs+Z4mJfRlrKaLu0zPzcoY/xgtqYiPUL1WB1HghtqEQYXlAQ3hz
bW1XpKHJ5IIiP35S63lCemfw/+htzeRRgZeB/EewUBRsGhNKJX5gDsZwTWMr+otY
mADw/VbLTrNNNgA8b/NpRWqWieF7pPonebZQCUqnOxZzw9BN+38lRz4aj9tQI4ij
UyxhUznQ2LLQzMUxLR01MUHo+9RVBEgW42mD+XRfI0PnusJHUgP6mrnALhcyj6p7
x0hVkHwIWN+vGjK3Vs0eHg6bsOPFazuk4p0kezYjT9/BSqiGAU7nlmVlGHSgm91g
/9nLhXrwm/KYfUqxW1CAZ15miTRJKUJo3KgUrfaOfVz1YuZxHV/V1gxeF7FvPR09
55i1Nmn+OIt8q2/HYLjvCPmB8ZgG9BhGphkt5wxhmN0fSwS+zRJIuNfE17FwN87K
enDwpwWZgv4HnF4t1zfosvHYILhFq6ByWu7t5gVs/MdReQaJmfQm7j9MDWjj+8z8
KKDyyvuNgJMTwMFntZjluVMdEzGwc+YwgUb0Jd7y3cOmJbFM+MzcoD7pozJl/ZFI
8a9XkiEBseI6TZlq3c7zeERdd6MRPLVfFqGlO0F4yXHjsxajwr0kr2/+TbUTFmgb
Oh7VQEZuD7nIc5nAZed/8cdRw9yOkuxERAxsxsKZ1L2gzozgE+N40Il9JlvvFsW0
X4VpWeHG1b8mvKLQyjKik8CwIo0J/5XK3/ziaWyKcUSkmhOgUz1/+dUWczyck838
YbHKKlf8x/8h/gLhrICAjc87gjodCL1V2vrLyXeYhRPk+/K54tXdjco1IBHD+AOX
UNAzpmXgu2+9AGUK/9uyH4RE9YTvewT3RvEo6z8Plp3kWHVPBh4RN1R0QEblJ+oh
GQH2MDnJNuH0jMk+r+jzfgNAWMeZ+2bQozD4zR1ssPHEw3kFU/g946SJvbY3jJ6s
i3KpF+vYSHrE4vWYVxh1g9rPwU/uirCeh5nK1Mptgw0wc093nvSG01fE8GIGSA2M
exAk8dA/ml2jD/o47q1T5M0Jd5GCvQ/udvsFJ6AW/zmGkjA8IsofH9y0yAKNowAP
bJge19LQ2u6HAalGZfi6ulLybFNTmKa7bRZEnSZ9Vs4LF0vgvUkL4Y0zUp3U0IIj
2oxaJ8dc5PNRuiKIeA2vGSS0n+eBK8bGRs2G/CX3Tuk8+5hcNDpDuypKAbkzk+2Q
2l4Nx9P0lWcnQh2Ke99GfiV3QVvrD+rHl24+7EsZwT8tlpNDRipLD6eR2R+j/zmm
g95IPFmJ8R3dxTfbz89so/ocLSQyNV07kZSAiPtF0HAJ7DpEpJAWVAd6uFrJ5JnJ
DuyFeUfPk/It1K3DPJjpGcq5GIVa69klqe5L7K+H4s+8mVr+RcaEWawJnn+r/CZc
9FUkS73WdB/EJ5JB9+tp096uILmcOUfb1hCp4Pkx9/YnY3oO22COI4U2I5xmzkPi
535c27fVxxlkFDihevY4z00a/9X9oE99mVd3HktVxy/P/htXAjyc2sxk48s/KxKJ
IbCO7Oub/b9e9HwGFdWryDzAd2ffpPZmKWF6Zp6RvfMgN7kVFSG7+v0r47KKqZvK
Gf9eOwoO23Aj0bZdxumkiF/VvMtBn1/2Nm9+29OcNHI2G53xL9BxKfzB5SF6JDAG
f0BxctAgORsXg0AIJE3NhVcc1wwP2otZw6pVkieU43/iOv6plCN55sR/vu7u43zy
2qCiNxkbTz41WiwualKxTu5oA8WgtErakbPdDLA2Nw9b+/NxWFNmcHutiQSixy7T
qFrrbH2tbD+mFjukvvBIf62bh5OEqtCnBisU1MhyUs9ty8mU3mrBywa80K6dOgXi
KvrcrGmowfNkGHSja9HXq6XYlcarfMkFIhuwudbF7Jewg5LJgTjktLoX6rqLgjdp
M2WN7DfUBTCwnO2BkFXo5uM6MnTDXcGlVksZ8kPpbwiILS7+qoz01VXlEysgRf2b
hNbcTrI68jwWOy4z/3169Rt/MjASqp7fHboGU1Fix7+66M4LrvUw1LMmRPn0DdPi
6BQcnwxAog3pn5PJnSn+ymrb2N4Sby5IN6tdXCd4zGrewzKewbGMMy4Tg/KIA5Yv
0/prXSgCV8rKymx2IYIppj5oWeg90UM/NwW6CVQ9/GxE3hofgvwfZZ5DdV+xoOf+
NZs8G7mSTnwUylynRS/fVN83ceYU0DocA5cOxrjOTz/OV9LG6NaVgiGjd6GGmJU0
cXyKQ4UHeawTIR4fLgWIuTLl8JCxukkKm5bfAeytYWWF6FmkbnQkH3M0eKJdeLda
hHvWweyWMQ6k29N7VpFxEzqOZELGmnT3DTMVK8ccBRWFYlFEQ91zNfQOx8KjsRNm
pdzgGRt6/YKm4TnO9U2CsJhFjNejBPDZyGcO5OLmlITjWcVsi4aR4nR+AaeEkiWI
K0wbZpsfKnCwGCSa8/PIkoupZhe+fzVsTWvUVR/hgqIawC2nDWdgm5DHET5dbHzf
sDR47whFAxcZ7ldVHNxSSvCGGGIhrGqlaeYdhOA/f9wwvN2t4L6pjcAEGwFAyWs6
Lzc5hsx22L/F+QaBOf+ZMOZtgWvLyTW7zU3kiyQAQdCHaH5JT9oE9w9aGmBKgtPO
Ah/uNOpgQ5+a0YoWapeotDVUcHaSf+C4CIAxtUZSUTGNRIo04TwJKj7HTTjqbRVD
IAa3IR5CgoDurIP1j2HT2O013cxKSjeChSGU+Ej0BWJoUW7WP3WyhDwuVeq8Q2fD
rSwhZw5itZ8YOHsRUG30ENYCXWOl1gCbWurRc9id5Qs3GRvRjZGhclhKW1841S43
AXKXr1R9+J3GwBur6/aWcq+n6KrM9VGSABnB7P1Q2mbOS/h8i4HUasR2NmGnHCsW
xHGtNvxQf8ahCTlkzyEr4MyGBuuUwaVtvAT8Ex8Im2pE3IgWrrmHYIqsoJkbF6nv
ymvPbxue7D6YPpJVzpNbRSig10Ozzulf0mPZWTYhgoahtw5f9/jsimGnN4FD/5Rw
DcYyTwZJep1xQgS+m+sTNe6nma2oMmZBkO0bzQs1A1IdfsDlaXT7YhWWcve1GcH7
iauezFr3XtLjYYVAHEBsK1eIzXVfM4btkAavaDI+6i79Vn0Oi5wPRySED16G0AsI
hu3FV8+GnSREbLDs+kYOF74OsfQ2TnyW6E1ueVdRcOsm0H8nkzjlYSd0+4mI387w
Ew5KBDneVTO6qkEpAC0wSt8EHEI9czSh6I4EUo3SAe2PO2Vk4fp6ARk8dHq5dCTO
KRwo/nDv/P9ZYJDjfSThKVNGVo4kM3JQ00rx4xlghpqQtRsZwuLOAaaCvOXpzjN/
fx7WHLntcUTGnC0QeX8jKwwK5SJ5cA91/mIqWSlfEvInPcLmPzu8vEYWc1V9qQq+
e/sQK7ZVKLavSn8PxAvjIpOdP850dg04AYptgZZrrSXnO9GWnG/okjRGNCgNfkJs
uojc4e05AiLxF90q6zqTDC+j7BDED+dlTZxBlh+KX0aXGu9JWfDeghAArIhkcU/T
pRrSjQQlzEppfjy5A1B8ZEAh2GDHoqCDSgRXCh6LRpaDpEhhLxet9fHVbAh5JiRI
311XXa0gjAMMfA4IMwMn46pyPUZ9W/8PBbjNOIW5wNQGUpVRCPcv+RwWJ/5iST93
wADr7e9bK0LSvZE15cBFkrcUftuWPsjtk0ISTnKM2Hx4FfREWvEIs8GD3AF+AElr
5QJJds86NjzMsqLP+de1iQNzXQ8cKkBy0c9bOxcbU/GYQELyjqUOqVawNb3kGoVU
hLKWbJg2aO8dtMLemJ6vbs1EJOVIkZfG9r+Jc7+YsxYl2f+Zb0mzHSnF+2KgQrZS
rUZlj99o6p5DcyecCwT5twzZGlsY2PzFxG+wouCNQ+RJIbWGoZh7UccshQ6dXvm/
jxlNqrbg/ukPGaNO2I03y5hxoLNd/LwmujnBP9F4loSq/f/3ndnOCOCadfJrAbNt
efTg1XxcDdbZY5MfT3mm8BzF9y00BGfEH+VltIrxVqciMj647VlF1TQdPJi41vri
OS4+62d8aRRRBr0Gpt71jHw3A9Vastn1Y8HppgE95Xz/Ua2VFswXoDc+isywYLNy
H+b2YXKmR0XdUcczTrF7nhHGMbk5GEYWjDPCbUkw/dIAV3Qe7jXTFRIyXYmd7CV+
rxBPV6uVUomM4tHzo0NDlAR9lfgrODg1I/20mfRwvJhTT79KQKZtfl3bDYHl0jUi
G7phvEYCfC13RHEIjtxxgrnai7HpnTfIgPgCWFjr3YtDa7Mxv9HS9Pg5pqP3zmVd
EZ+0K2ep2ohfRf4WYo7rmnHAOweyF+y278ia5BIEKXq8y0m8D1RQuSaRNleV5K4E
TmmxZOfzUXaxwlygXsSRD0gGzm6N03IIFNxwbBHOK6Rz+xetWZ8NovUiVrDpnNMf
+Lp5LP79r6VS2AzMssNTEwwVB3M6Fd0mWbWAR5if/lLga70KhN9VgturWMvIUgdr
0mBLsa/ctvKpU1LOO+T2nJLcqH/uDra4//5peQWxhxEmds0y6ZvPyd7nr7RDJQZP
bCtF5qmBQl4CgYB/T4EnD9cFI9wgK/gMPrBK1X8l7fF44CFfZbLUbj3RiltaI68q
G4Lm95ekxxKQihDnXHO4Ol9dxmDcG361Aiym4cx5+dusRkjCfN9kHfUbrXI5y7xq
C2ITaBdeRFjSWTghe9/mGl5XjHs1JSYDPhDdzfKu+0kpb8aLRIFw/I+aPLdAXovd
EcTcbHBIevcSJEXi+y2wbpYnO7Enz/oSUhZQSRSSK8nsG9Qs1aIvfLnLmShTjGEn
rDCzjNAU0R4fFkM1yaL/sx1zikzPdtYJwpjWFYtn9QnyspxcpokXEVJoP+1rfDE2
tQIvgYGMq1xgcv/B5NqqEKYWCyKX0irISN3dcaiwjzTtYTWVhLDQuxRjikNh2Imf
yeGbmi3cnN4/Kto9yy+MLorv9l0KE82qVteFzz8hpKnr32ph0w6ERf9Bm+3KSbMI
1A1kYmg9raiN9iy6YrFtzyJXC4OneGbY3o3dWKVYYRF9a2YGRnr/nE9QNQDLyp+i
1u14UMKfKaP8JQ1KBGNFwCEunfleOBFqKZmiA4OEuPAGqFhwEftGxSf3RWa7y2HR
+Q2uFyIFA1oazO3QInTWK7i4WqDOzKSNxpzbqTE8pst7zcdoiwYdsyjYAxm5uAO+
Jeb690wBKJ8Mish+SV8n2RyPM/cu2K8IlmqHoW/2zYGrd1Moy0CRSCP+F383d+gC
iDHL7b7ON/JieStSfpLheMe7RUeHtcWen6YN7LETV0A0JHDn9b9jaaxfp8OcGF2O
w34UHhTsx665r5bJUJEZPN/4ps5gS1qPdbWp49oXlpf756a8rGjQV1WaIiZRvQPl
VAsmF0tH1q5BinuCVcunqkVqXcvRa19da1cBRgJcWmn8C3rFBWTxz0dlsUpzEQ7N
xgtcheEycQNLGUGWTQn2Fi4hwZzqiS/tfzB9fBONpgNvc2S09ZamdewZ/jy+G6RA
7s9PdYgSwEVMu1zg4CcAVup9t9P9XfAk7Hz2V7OhcNJSIFKcAbSQp9uLEISHG2I3
3c9ccWnterevEEJFCz4ykFdRAYgSK1s992iV/QP0rAjZK6pwda9fDgVO31KkMAwu
KboPPA5mj3EBs1PVRSpixjSydMyW/zoAta5atvKWnEDjCQSleALVL7hrSGC06pt9
HMw455YohI4uBWb0uscc3E4MQcerpyz4LmZbDA3FNLx6rJL3NSR25lfJ49NhAl7z
q7OtrXfN9TBYwvPgoHVNeFSBtFwIIHLbpgwdy5SLf2d2IoYIg7ClfWIoDKtquAfH
uSXQJNcXOAH9JFO/ASvkXq5iA9VhO4TOiiR0JDIDOJbqqowQhjGHOEb+I+GkFEIU
y3E/Dx8aEalKGuQacZah4SONX52b99THWK5UwehKtqqBXK54pGuwldYQI0SdhNpq
QR/dZqZttOm8x4hLxLxl2OriHEm01jxjAKDpEmBFBbxwZcZB/NDUCxF9RfAPBfbJ
22eM2d2bfh7mSiywz9/hY9XXhxO77KkuYJXFoXdkRkkSWa7bmo2H7rRs+YxbNOel
nHz+2v3euqeTPSVmcOxnUitvzcOUTGnHyeCGdp/h5ub9Z56+eIZbhqhFhw/KJSAo
lLGzl09HeXQ1GEBTzhNa8BlhabqbsfhdI9r/RKfTch5yfnoEiDdsWTcf3u41JFks
NvMXLuHL/fWMCSPhc02xXTE00g9S1kahYqN6nKPp1TmYiIK3Ig2AqHy+uoVZLpxG
eh9qTnJRVPgWh9SkAd0/BIrFi0BurxNUyNB2HQor9BU7Gz1ha48Bfih86QFJoUUG
eFzjpByBLSsOw93nPa9IFa65l6huQT2zUVx5ajx+cykWlm6sQYndSECqnZkJRM9/
NiFS/iYZfZpm0Dqs7sIOTfh4N5mHg9CxZa8EKz5pSaD3G/2pSvlxdt6fUCrBaRLO
4UB0LiFhFHEmsYDE2xYF7ZgLBMnqH2hyecFR5m8pOUu8bk5vz0rXtoBq+F5YyUlE
Z540brDifQ1K0wrRddetILm13W9kxjk27M5/iwaMhfkAGn7b9DF/L/DOMxtSiodA
n9D2MbcNomp/CmUiuaopT9tu/BwYXZWr9tBHTiT8IucBo6zIWuNmKXf90Ps+CQkQ
tFwhVLECmE+8MFRR47pzw2PUw8zYgtPCAXSv96405TzW/BGbJoCIdCX++AHbktfY
yF/+/OF0aFyeXsjPCcN22j0xi2pr/PveKFV5s0TOrG2+4CFsCn6b04r6echYBucA
zKbudQt12ELMFKhmTzvw5hZMkcrvSha/ueA9B1k/C+/4/fvc90muNIkoLaMrlZj9
RzRarvDmTFAObHkz1QZdive43KyBaiqibRaoLgwQVUnS+vybXYSl0X/EpCaq3RLS
dCJyq85vM8qlKl/6fQJTAZFPlG8mOjqC6Vtc39yY7aSQq2AEmpZYInwPhJiIMix+
OF/aLasz6tAT0mB1PzPuA1l8JaDEzry6CBm2SntAyq3teSczVfoYGQp8dmC+0yJE
y50z1wqfjSS3irO7m//pgJmS6Jtjqul9hl1L92ZrKwBLXK4jx0i8e/ZFY5vkQbJM
YWeLH8hm28ECaZWwQBk/YyeOreIJ8XTYFWJUIcugCXtG7dDRWlIsR6V0XKpkGymv
F6cUnue17aJMuT9r8oZgjXyDxTGgh4ziOiropJIMF85vT2H6Tb21RLKO5klbajHU
xf6pAX1BKR60tsD5WMwaIcHbZrThXjvp0oJASXj0WeTqnGbBJrRChvV5l8AlJnVC
hhveAQj4BUbJ147Xx16wQC+u167w7085s9Z2ZhEmmrsrD+9jCopQWUaZ/jw1m4Um
d65RIzSdm8b+h2xJ7GZ79QUMke+x8N2SZJi/uWi1Tjn6mEXM2Cnza79cq/0Wxz8d
Q8WpLGtDMU5vK+bMUM9A4jJpXOhgGukH+QnrdnPeFNXwoBkgh848TKeOqUjaoiMO
qH4NmIamBm1hoXNnTs4sbr3sgiT20ZvBniy2qxazOIYojxHTrCnNJXyCjj7P3HTa
r7nPBQdsqTs5rVFK73GcGCK0QJkiCMNNA13C0CB296u8nf6qcUVjcVIAh1VWtm+b
1wPq2xl4D45PTmZAWQJBmtC8zWceMmFbtAUVFs16qr4Vls8ZctFMldJ4vJeviQmx
B2lC9OSbDUaBN4uO+iELvbZNQ8EpY5HtfmHqDRWMQdxFHZEHhghy1ArcjbPDOK4y
JPbX6uXdCVj0aiK7n3YqxHiwwGbKZbRCYPC4Gpc+XuN4GZCsMsDzW7AxGdtq7EoO
Bhn7/lVgwlVvqBj0y3OCZ/qxcKGEYVeUdDgRQR8Rf2NYAlFdcBUVERVgZe9cGPeK
sjB8DJ5KnY7DwdZUpuZ+Zsot5oxqFF743BFa2RHRnTjnCHlvaYogkN8WBOM0OZuC
7K9guIHMiz5cFMlVNxhkxpGIcGPy/7m9qxECVLdo6F9+rHNHjJvOArbpDo4dANod
V6z0ctYeeH+V38o7qsU7V5sqvjd305joWNZGVliGUR6H3Z0ewjnOB++pkQZCOnyn
vQNghF+IzKOHZtESDU26V0oGuRL8lVW14D9hEWsfwp941IgBKz9ecRmNwCGnJDGR
u8tXpFjscN3l2qrX6lIUTmMgu1gLdYW3dXar4MlajWSxvBdM9RM25xgmidzRwLkX
iUwcO/efJ5zzL2g0bM9EPaaKJUHWprfPR6JbCugLqULzdDZZkZ+19Hxc9UNfaC5T
pAiNY9k56/RzdS7J6zWwkMcMQbtr658jz8pUZl8cvs7bl7oLIHkTnrgPdUt0Rkw9
iBVQyu8PCHqK0rCIejW58U4MDZfUpQLmWej5XDDOX2cW84DTzKeWreV7S0qsv433
/gCRJtt2up6SpNT9NChFrV7uztMicdswG3wwOBtAvhgFmO8QpnWMVXOhyNPbwns1
1nh3qJIvUADA4YchemfOlaeaTfwo7w4RaSVaKFLmbJYjtzajlavyThYOfI/b7VnM
2NLiP8xKlRHSEjhRyqzkwbur4OgkR9Qy8jtW141M5/xSshN1TqNG+Yo7Nx7j14pr
yi5dzz0pdcnYndgL+7mHUTHtcClgR9TnP17JohpzS4N9n3RYj0JxJGrPcixePLw8
ox9ugvGdEhN/k0QqzwPydkWjjtyu7KQahhxqQKV2+qeQHrKJpm1rb0s1Kzc2joMy
B5t3I2T+lZMCSGLPK7lKeSCMIL57ztbAQ+HMFvPkDPqkQRjMfBRv0a/FkQXP3yG9
fBDsi5vx3P/IuMYftM6AMgbvhYkVGr45QUubbhRatvzwITBLL4V2y7sWC5Cpa/Iu
5T8QUChRrlkIyqD1nOqtI89K8N++7cVcMaa+QrwpzUH+/bQ11KyfrkM/CZEunuj6
BmADXutb01/hoI7ULQMVk2shAs6HkhR+LLrxiCuzPRSQC9Ym8sHAtMyVOtmtwIjH
gzNaiNK++IXMOcF8d0G7R3MJqg/hshkIlxyPf+gO92XIdtYIk+GNzX3sLVTgiYVj
ZDzrVNgk0Jgw8XTX7W6gyyFc+BcBVhEak7c/7Odpiwv6pibUp3pqK1w3CQY0BLdL
/v+v1ANOTOG9pLx3R2oArD8OnvckYlyiuQCOWd749b8DunHFFoeT65S4TJ3StbvE
DbiqTXgn0t/O5OZ9hTsdf55krFHQUZUbyckdaB1ciwe0z1ufupUzXF7zc7fvT8yf
AZV2aHTlXsbE4tBI3f9c/zcyS3KQT0h8/ED9SMzS+nGJaQBPCyhu8VYGmz8fgX7D
bmHxKLbecEom4mft+7y2LqQOnulvioCqwUizdkun35I/eCUKb6A2rQqGEygjk8tg
qx+LDIUtt4C+cO3jGM6rBEjDumO2tQnnuZsIdUekQiULwajjFFUTNVFz9FeQbsEQ
hU8s9VwRPKz8RlqDJPdjvPk6IcXAV+iQu5YnRyz5zrOnj7a3uqzKlz6qfVccbHkc
/v8gzvHWaKayrr9UZohtUry5RTpE2kmst8tBlzA7ItbD4jzR7sqqFCH8fK3ZPSzE
JQmgFotPbov4TikspS26KLWGnINWn3gWAor8jzZisMJyQvNBKFnv7bDDmRkvn+US
WhiboL6syyRo1dbzz8umhq8alOXXmw0r5C9OdVEkl5STNduPsWZ+/4V1d06azm72
qEUFtqDqtDrUWmT2bme9fbrEYRxNg2QQ05vzV++N5qZzDR5+3S0seBq5z4Zlu01b
YVjrcwi8dUa4AB89POK/1H6HmJS775sZCNF77Yy3p3HwQH1vr87ZiZzHRYphD59+
JmC2TPjrvukDjXNlC80kt06EWe9XYo9sRKaIYb9ihU+EcyZaAKhfRn6mjnwv7yoX
jLXjPc8hsfwf4kcMIrOJfrEVZ7FcnOPpQ4zaJMX1MjfjyeJKBdQEMCfOFv8SrzI4
J435vWQDwGGTz4wKFgI2aqRd4Br/o6pxOiBMkRLj5n/vJeh8f1Lwfk44D13gbA5i
yugzkFZUJmNQo7z0VWrugaJOs9CZ9VSEzLvo8yPQxWHoS5SB6iY2BkidnXCBcGhg
t7IsJ6DMxSkPliQvCbkSH7fLLEfoH9q5DD15EYP/jwj83LyV5S6XbzEQqGXw8nja
O6YmIvRKFe59CH+sPsxis5OkT+bsjtWx8JYrp629AeqrNsGwW6voLcu493nZuetX
oxoP1gcqwBaLIqtj7kjIAfNDIqtqtHBw7+ob+yz+uTnR7d3w3S+AIzlVRStnchC9
jnHw9D9wcCd9Q6bUa+BPwcJ8ivA2DQutFStWfFlQvSCJVEty92PazcWFy2EJCKop
mzaAdzwSDCr6tFvFlPTYvXfF+6zKU47J8Wc9tZH1+EaodeuDWlr65xFz1bXDzhBA
4qhmlc0I4OIKHdKwOxGivVeU/W63Dn8vS+FEqjGDDMJOfLiiKBmyq+TA4nFZ/EKN
ucC7H4D4FrRPEV7dx3O4eT0dBq+BdpEIKRvrxJLRlFRox47zgoRPgTBjEXRbZLjQ
6vIx+e9nVmE9L9rD4JYYWy+VihYzhfTX/wmjBXjLq5XtXz9ckxVLvuu4vnXyc8kR
y0Z5i5FEMEG9YIWscjTLmVwsmNqVdi6tMjwfPW1G2XWZwA4Nt+YRf7lSv8vN+HpV
n3UEPxkgyIi6V82HUCjX7vmd6BCkYJZANx9TGOx4mATPMLXQfcEEZdRbVKSMTtRj
n7dFJ3oTSpmpGLL6KJssXCYERiavkp6GY3UD0fB6tS1GtNu0AADdmU5/65Q8yJl5
VU4otnjjfkxAKkgCxu55PtsIBI+MPxAefV3vq8OMBKUjNgUmF8+Fgmj1WO87jwsq
XFTfWi0UFAeDMJBL2lyARIVwPrP4q9ZSH5seOPY0K0nQaWB1cYU0htmEcgNRlHd8
eJ+41VNWPX3XhWFGIvbO1X65f0UwxAD+8xd4/pAKXLavelnYGN+3fhXSqXaz3+i+
BoyDlG+LS6YO5+lIwNTc7A3NE9A9DhCaatZDtDra4YoJ/2b0NPOLmn5omv6ZOa8f
AZUH6QreCDJNJ5oFsQhjB98C7dPa8k5INHo2olS8Doh2WvScByyksaaIX+cYgClh
zjVphFAaIvN7znDXcJL7USbo02GzmtkxsgaBMWDU0wduQV8cppU2Zl6a8F8ibi1C
700L/MOZVXgmGCMUhI/z181mpfmwzL6FvdvrGnGUzzo/yll9JMT3X/vX/hoy44yL
sInV5DTXIOPMs/zT9sqrSDGFqLG8h1zxwZUG/n8OpwHHSDFk9bsmjfFZVwmEsOGZ
G4qFnOc5x3kJJS9KOee533XwqZug9gcIwcfWpvUv+QHVyYo+0o+bZzrtcnoa2fdh
K15dgbT4nnir4gLO1T2P+WcMogbh7JEnhw5Tz03rZplnkeE3HJ888TovQEeJ7azY
efujP6bWPlzB21aSpbxrSNvy9rp3vxrG9e8x2a9NY85WfnSfUbODgCnESdxOJ6Pq
Zx6OctljSMzQDCiIIz7498sTd/DRRGqWe7n+iw/8m50/0HIQPutpRtb1MkBuD/rf
Nmg8TY9YHnjY90IwGNtYPnh5LUOqBpNvxc1Sfu40E3elQ3+gXmEJwizW2y2nRM8F
ZxDvow9ul/gxKEiEMl/H1HiRakneyuy5m0GiaFv29RU22NFptGQKzzMeZnI1Xfi4
+mt9kTwVPzQJXJ+bSE570SdWdMkgm7vEwEHn3ydVSOxeyDblRXuecJqD2LXxVsxq
P5VbIGkCCHLYbe8hMnjY+4fgOllF4DqgaHaBakBIXPHuOJCqID7JWhp2zBskLEA/
kEqmDgzSdeWs/NW3V/lm6MQ5GC+Q6pt/HuoCiDYVj1IIjvofHI/nfXXbmMhB6mfU
0QZtU1QPTzhOhsIPfq1Y6gvVxy+LF+SYTybnX7r1c5b4gYrZTOe27MZQ+vWyCy3h
sm6OY1weMiUvFWSSPASCKSvvdWI2fBz8b7lL0AT7eAJNLHDPfsv/5wuHogoBtiu2
rNvjerETy+5Yb0J7U5aY5DbRPT2ryCmOZRZxB79ZeGZn4NJgfvGSNs4E9Qq+csTo
OW96mj6G+F3AOVkz69VN0n0ycdreezVdrP+fUzM/QQ1O1HLOdXfFqvg8fbXs1RrZ
WlzXkounAbhMf3xci6bK1wfV4+0LvD87PHrIZFUKVBsYH+DHGEjp2o7Wpg7d1gwh
KWaXy4EaW3eYMBab1c/pxMbdTNiU9yERtKx1S1lzb1VB4WUHGH5edKLD1QxUoyk8
YV0BC2bsx9y02z5Wo9HZB7uyhTqDz5//VZ1yCbFeQ3K2+XxbFXWdTlNcSi0m9ONX
2TzbP92QzpOwuTYx/oEe1TqN+5T3c6vBVvqzmMgONWgMjBUQzpRFaygl3pTa5Kf/
+kpWT/Jq+kzVOxIV0ubeElalQ/ZpoBeDIWyqgSd8FPCEvQGHwRJuwhacl7OM84Bj
/3mz4KcMN6QjanyaRS0hd5TfZZEtGyMNDKDA1uSxe5svRvuePErQSX6DmNq5LygM
WiAXqm6fxKx6tAjlQl+B+d4j+EBOsmPCmXYmXAlqIjxcm2peB4boZdq2ycd/c2L0
v41CNU4ercnwHzejCli+G2lqUsq8dVDtXT4GrYWYQPudRcOYo3XA4ufyCcmN6B7J
yCDPAoVHOpD0fQsx9070zY0iABWS72tC2RGrOYswO4zvDsVkHYalU9u+tRuKiRHB
oZdzxelhrszkiEfZZvv5bnfTxb06hCk/kNJbZWEHaNWfOVwGfweQh6vfQJMhqXRe
aAXSi35NegSNg2/VOUofIeWwg7eLmbNJQxyGrReeGueGEtKbDMG7Q8RofwbPdMSn
sinBNcx76gM1io1xnZ+Ak78EGpAFeJQV4Xc78XfDyvdCG1UXlhvGuDDuf6AD4XJU
F28632+DvJyA8hmbl4d+f5Q0O3QV5bTFZmxonEEq1a6zTQqC43HbakQunxsIOuiz
U7A/iXT1S4WUvF8PA8njSbmvR/TMPGo8yJwVmRK3oalIwkYRUrcal6P1kFF+qqug
8okLHgx6YHTaE5TjANBf067TrrVzY7mseeZQqK2lhQaiDUaTv+SDONxXyGpiAZBM
2sya23e0apTZOQAsnozvwMcZ3almPpx7L35TKJ63ZglNLOsJmxA9AUB5Q9CDJDmr
4VfGxyMhLePPq0cCxT4hxJK0vmhNBV2iDTLbMtCwun7IH/zA6Zpr2nh5ISxP4LaG
iA6kwPv39KbL9rLfGiA03ZZ2qrva6G5wsNzHH+rVSB8J8P3JudIK/BnZVnfJgMDJ
zaFBmEfPF0yGvnbUgcj+DfxLrh/GEqHpmNgM4WwGsVC/LwfYmjbxz+ixyJN7qmtp
hfblWDLTJOfmw+B8Qq5Ay3AKskvt/T7QXHfwQJ/x8tg/9ztBREpI0XVXZz7SviHx
9pEq3vR7G3KX3lTIh3ed8eRPyard6p7ps9Yov7yRhLtSnOmRAeIqaKhdCpByh+Nq
9ESLNQUPaPDD+jqc2GZZOG4NdBf5KsOndLXV86sSg3aDGCa9d25zuxLjpv113tSC
L2Uzdp7qDmi/7kAvhtbOHAYxdmr/ojrgp2xhiRm6aMgCShByeVkq8gDMUxS+5Tyi
7Q5csN32nqMH/Pd51UmmXAgoh4X5C+u89T+JvFH923hprASJmX5WBxsUuSGUJj/Z
gNNQMeN9bRlQI7X317kRYmGQey61STQfvQR3Nb6xsgvsKwA4lysfAuChIHF6e6MN
OzVDL+UUuvsKcrKvDsaNcCEES3eREI0DwA26Rle2TdKsOqHScyrHpmuLnb6R9yW/
pl83C+RrhMnuk38flTvqYgcDX0xCkzi7KZverSGST/kTMhwiyPzUIonXgzIZnmqk
uUXgRTMd5LZ6/9GhXs8rbJqL1zCd5Iavny27Db+7kjDdV0Tdr43Q72SqpMQ/1Dye
qMllEdoNm6qViGLcCtvxv/110R3THaY2KWpYYg7nRiOUbu3HCSA3fYj9+1wWDHax
2yXEJh5fRRzOsCV1Sze5BFc8D8CYjIrfoVp/3cPIFmKuxBoYbLFCXw6VXqT4sRoo
9NX8Hf+6DSN4i+2pOfTJb3xPxn9EVxFPScYIv04unpM5J7dY578D74cxKYy/UKbN
1vTRLrpCzMS1GZHO3+O6lwXMxv9pXAaApmTDdSC4N78YxizmVUMJHLG8jv9MYWdb
nIqiSwi8cQTd78wHNqnV9JGJJoSsUV3T+0Qj8T1OP5vhpVxOoHQHRXDltqz4XZrq
+zh63Xk1goxClsZUpsmtpdGAtJbvQ5GLyCMJJTRIj1/F1SnVhbMl6M8ue6Vzyc0i
nlNSJDQ/xzJnZ2RFruLSgt6zaq0HEUPlP8tNySw2zq1lPco5sQ0FIO7qGbuPru4n
y7G0wNzWaChy81k3bdHTuLa4SlWIb2nsot/aptYkRRHHhjGH5MZA4aQWaWmfeLyQ
s2/rXCFUP3Nhp/L/2BJLwlSVuNwPZDIJT9L+BSZDnePJ0OMH3vS+mb7uIk1cQm0u
EFAQQaq+6Arwm29KhLuNcoF0nGlBnsy6Tmli36Iigcsk/kiGYSWG6/akmsnl4qXk
D4kAtORpHD//683LhU7h4FawXf/75SDqIfvJT3pRslh/TKR8sL+74LdGrzcp3HWf
a/R1ijE7/QhK97PoID8gxPaeTQtM6pXz0nwNRN/h5D3kh5SmCCeFrnYjQ1i7E72V
5fLFWaJ0uLLwsv2CSrDtkDKsos7YUYUJ6n2nkeW990fniha5qgSPuM5qCQM40FbT
oJ72c+8LWgsVWSVCgDsRUJerME8U7InGwgA46oqrKSCwzPMWqHCbzOLaTlyjkibz
c2djnhR5FbO6njt6dTFB+03sgyFwS6XNtxnTLOdlgt1sU7FdHzPBzghJunucwNat
quDOh2fnN1zkB/93ionfdAQ2IEA3ciu0d5oZo/ZAB1+6CnkTPqSMKoSHXELfABEi
lgIwJc+f6ivt1JqW59ThRsTZHVkCRLZTS2c4DSeBH01iNK7gkWXAgMju1b4CH7mu
UTPDe65+7Slu1FkljbLuLzcmPiC/9KdUi8ii5Mwl+RVUw8wXpEflZKSLPfNxkbt3
hzi5A0UeWpSHYW4tvtogdVMtf0uROvg7FHTZ4IXb6tEbmZ7zI1XtrR6ilaJDjuf+
1OrnLdlH79xfTMKDhwqzWfRCsFPJ9Z3AlyxCNsiCNKGKTnam08XWehznSG+Hv8wd
H/bQIKIRPevmEFqf1fO1ULigwGPpYf51dyM6s1QlYpM4X1fyzbAONp6XwFfHKUPm
HxklEl2z3WbrtLVCaZG+FT1kbdHaLRdfmdYkb3oSin3dqY0n6cHWxldI8pCW4dm8
uduxG3bVXtDsYU5qCvp4BrZ0FRWbQKAkuZnlbcPFyKhvCdnspUKmw+XPbe7d3bqX
tt8RNCfU+PTuMEHvkUMmVzrPRH1+cS49ldCkIH7ngXfuYz1CV1aKPz3YO4FhWAYK
oeI8wuaLjemM6sXYsUW8jqCnu6hYbFSihiyCdWas27UHES5aDemfST/3zdTrvDUq
7xi300lAkOEI6SezubK8bOdk+gJpm3dqAeg8D0kH9cXp3iPx5y996mAp+/njuU3/
cZnO8Bp/r5Ds0EdUiLcsLHB7yANtd+iFFpK69brccprsOhkNQUxJ0DkEY7qLG7pM
6sgLdRzch2hB581w665oaDe9H63LmMfsVApNbkl7I4DQhGKdSSfi/+3XYuNUCV9Z
Y2czujjjeKDaNGrzOEI2LSmaILCvDMUk2q57IkTUl/TWVIIWh/urm1sY2b9BzJI1
nRF32o/l2KZ5ftfpQhUd22ih6O37JxjSIiAuWAhSN9ArVBUgDZyssbz8QB1p+jtp
HWgJENVrWqg6cTfPe2DlI6tWRCSoW0R+syhGt/2GpGg65SmyEZgzrMTTLP5E+JNx
s0eFkTA1S9FmEM8exrwRDB/pnL5HLkfqdnoydnihDxXIyaQMGWaWtUU6gmd9wu+f
AkM34gYbgOLNHJ7Yh98xpeQfVuENHyUtAK4+CNSsys2fwmZlqwAO586DpiRA0Qvo
A9fKh3HK7BeVhrEp1TN+qpa1Q1DAeZL7eg/azumZOLbEa211WTEzhNdTHSgIjLRU
0pMkMEMGQC93LGqE2Kq/BxUZrRZEl6iepcB7ejONo3b9V6UsQrBsUhCJlPxTrp8b
kCOLc7CQV7CQiYW3oyo83sfqC8GLmhyvavj4Hg4xYDjASxf+J9ADoxgimZJ2dSTy
ccfzEBwPnjldcnck4njoeujRuSCNj/yI8NtqNXMG+zVsQvr2QU3NeNchIslwYmOL
WOlgvgluVsfrQoHJwHfqbyBdhogyg3tkuqwd8sfYxUvrnqPiNoEaT6PUCODCMrtb
hIPh10YumWbnNpavpxW/55z7rXd9QB2ZMLaOWDLbYSbCSRG70G+ysiPI4Zc5z2yz
nGPWcTRf/5NRNSuAXR1e5HmpaeKN12uJr3Nw6lR7eIiTZTwdAgZuuXLV1MGP+OCk
to0RcaiTz1jkZKe8brPYDEwfkWAEFbRvbYR+fsv+j3LbBbAhN/0PEilSQA7HhWRY
DdFiuDIWPa3lnYSwN9Mb1tdWOi+z/AaoZ6KKNintPgXAoXxHVZQWrSFW1wSC1geD
npfb6aOXKzMnHBNb0CDbalVK86Ngimj7IYkJ0PFzzv0xBpvDr7SFbIThen26DhRa
Ljy1QS2NlOBApClAzIWt3JMZ+TXbDx91uW9rdd2fVr3Ho9D0P2L4hQR0+Iu/A76/
EeOBzV1i/vo5tw1qBtEcke/TURy9JuYzDQXGAn2SmwqG1g6oRzCDrgifvUYwq+8/
txencUDYOWJIU93MrG7XY63Gvg2okmYJkgr0+Aqq6CSqsSYorP7059XU4tkL6bw1
O5fUiGLBIw/OAsRmiSrva3REH7AKX/y7EXcjPNZvlh3PwwpX25MNMeUwGGeFVg/i
Z15cz1t4DXWVmmqpWqM3R7o8hq15u6ghPjypWsZkUQ8GU7QB+3PyNlXdmM83FyYo
ked0hp5A8MXiOMOseXBqc7rkBZda8fy2mN0bF3uS/2dSYsy/UVN+Zr5RhafTrnYU
2vn3ySovj4twMGyyS503e4ItTTtq2rnpKrSAB6Gy8DXEr3WNms9K7lghVt9CD7LM
DLkp670oY8fLghfP0Oa1CgwfU6DwKZQKrSwmjPtyyqt0VKzdPQoOE3roLoLkZqgB
AnOIuUGz52YiPwc8GdDbzII/SWXLORLavmS5AddJwY7SpW+RmFMbiXqubuu73ERl
YU/NGGa5fPFoCTwfSCXK5468lUAKJVUcYJ5bscWr7dLVWcQ+J9sBZgdPpxVgIoaX
Q99UN9jinIHrM9Og34Dnr1FHpQYFHNK3u+aAiFA5KQrIB638Y1Z+9s8vifumc1lt
ehMqc4ulK9ycG3KbOXHlQtDlSSiJxFfbVEEA2j5yLxU07Bv7XUs0VgmvH4u1OuDS
HmffKrP4neuJyZvsxyO1H4Yvxud3aethUEYOiQ5bmhj34sMCN/Q6mfUlsJfkjrOL
mG6ld5d6t/Eccnvz5cHK1MEk6SLM9unrnoWLoN2ZZuPzzZPZC8yu1cdRE2x0xiFC
GtxMoCERvyRMpUonJee89JA8R5DBEo08Rf2yKNddSe7DGcRXEpw/ws/GncEm47nQ
foiS8HvfYGVU/hXpDnLILuvDDwcTyvYaqvtO4cMwWKuYpnoGWJMkKyonncZY7lEC
36bsfauU/vyoYBFty8Cmmu9VrTHyXvtML5k6jqAx2iv4gnaAdUuPNYEURTjk5nob
ZVsmR9Xw1aFwyqH1fD3kA8kzviOt1/benacLtCDrQGZBfdjE9c8RavZ2o+eb5ygf
iAf7SYimyS9VJLgESb8NArbf6vDglfqAY+DcXGjLoV3CGA0EL3bs7SGKavTHWg5H
HgIgw5rNAR2LHJlMR/Tjup72eZvEM0v9yUTGyMko6o0A7KRqTZIKFNwYmenQMyfJ
yRIY7Lm/fzCQo2Dy/TLQ4IYGr4z7XVcrYJfTr9v5CgxkzHADDqOT8ZL+25EHbg1h
HPkI6AHwSXZ4Ctq/VXTBjKggq/bZVme6XznbQZOFO2vqdoEA2qPEBSjv7XGWtYRJ
eAAsEkVZ6ZlWhsHtxNQO6e+XfpDTimghpChM6uyJIuNCU1A+8rQToo0bnmqHmDU4
I/Cm0jdhKGv8e7s1bqQGYpKNzMeva3fL5T2J7BPjQx83ULY+b9WGmCNlLKPozVCm
hLPRbGIyzchNaVIef9zCifzxVjMmlI0Fx6uyNrS4wd08HJYYfLh8MPiIV2b2l/Et
1FpFefWhLZE00q/BdzSwDnkZHhQgeQ4A0N1rLUdm7DuA4Z1YE6EJ7AWTTWYmF/a4
qdV/PSGdbOl4kNJuAAeCMJ992spux8yecbHWlzfLNs+lpCEzZ62TCwaoZWgiYn/V
cGOQgml+S4po/umYLuXJSBH+9dtZJXAX9HPWcuseYdm6tI1qabpdsjEAs4FUguab
QUXZhHVrq4dNvaY6HhGmhj5fuUKHFw2UGJ0fWETrJ4G+Dc6MIyxZPc1F1erL5CTZ
5bTgbI9Xpvl56BCwnPQNYLGb/o++3o+agh7+GMzZcIUTcGhSovdt8RROH2dzM1Ny
dyFsSRshRPHacF2YtWUXHzhj6231YkT144aFC/FpTrDwiNIW06PHFt26OnseOq7X
gZTAcY8uGZpG9LMxy3DBsVJcrED9YNt3wU++tRHyJcd3vI1bIWJNG9JbASp8COk9
vtME4GDdpRPi+cHTYdPwnYCzFj0nXc534hbSjUMfQuFZHRCm3RXTKpZq4wLxCmI+
qwEr/95+kmmDOLUfmqj5nsOdDcnA20y63tXSuKsa+j7W/LY2ZvBSkpW/tr0M+PCA
DS4Nbvp7FKf0aoXew4TxQH/SfbrnU0QOTdLbMwjXkP5np5A1oDRyURhC+PLf2mbC
XfjFvL1oTCbcKSjAtvNVtLpNeGt1Z6Yyyx93LDK874tmn5+tmgFjlhjVXzt4g0Dr
t8NUbuvLrIZMxXAwRJkHBB1rNTizlXI9awMJz0uF+htTdqqQQIM4wkguJdhfV6cb
i30ZHkzJakJXNodv1lq/kslSv16p5+wk+8YBcNr1+IM0nX1WU8KhCQnTATKn8NpL
iAZXCzId7W8SsxPlnKd7cUxlDaSWkagsbJXBSUQQjluUEqpp93sIFAOQ+hFi0iEJ
5LMlyZKzYTNX0O9GsAXTHh9yim+fpXArys6/E3SZECmE9fgDCLJ0vX1IzJEou4oX
DrvUYyTz0toWJWBcBJ39Q2pZoj+rzCw6GR4hqSy/GhoFK0WPfkWl+AHcZnOATJGQ
2hj9akM/Rz6PmisAJ5LtRHNUL37G3ZLIVL64z097J71sr5p9A4T4iYfboCeKT+em
LX0V49awGEmuZ+oOaM+jTu5vwN7pH4e8ray8efmKcfRev+nNFy9LJLuZ8kieUUdJ
ISMqaPS4Id7IzeNhViTtgNCuFu2f37jsz0RQScEQcrn82IpTH9RlBG5CixhryB8g
jNEAty/AKDhJCn1KINNlBX/SFkvy+g5+GZgkQq3fsnCZnzIwv6acLX0l0P8Gb/WF
VVZWzjDRowN8dw6j+6gC+WtwjY2Fm8PgUeuftV/lHTpV13wChrbADQ6VclaYahG7
8NOKy9LtxdqkKlEeSTYtFJm16UMRIkKqOJ4lMhQV5en3sSXng4Z4AnkKevryHbRY
t4aKIp6iwKT0yfnNr1efSZijDXtvPDERkdIYGH7WxEBsX/V3zRbbsOh3NEWYdVaK
FZXg3ga4SljHRoH4c1GIaK+8MoUkSemy5Z2tYn4d/Ovu2K4/lIusVQndh2ibcpmv
oDcz7cvqMFtusU9IJf2G6aVFAgYO0Lzm4hCvmvVmqDDnCn+ftA5K3FTj4G4v/qbf
Eh2EUCQdyqhRS0RI8ksd03Iuo7aIPmSHvYDBWjqiscvs1nTzaDUEZ6HhQq+2xWKM
1YLVFCCEJ6OEdFL9jW6/kGfZR7dPwVZK4VT56tnbCVUNN4VwVQLn/fXsBzRvbiYd
0RNmYPCHAr+cgvMkPqMOoNnsPJvU5hh7KImvSOdTAdfXDe4d8y1bQuz6rp38j2cC
2Axf46hNExsuzZOSI2JjkCoqyP/3Qe8vlehuZNV3haiyuc/YUkmQtjl72n0XyuLC
crNBp/PkzpSv5lHEWMQ6lEQcJphzikf5jMpRnLcoTAPznhxKjYEY/AoJ5ZYZpZOU
heEBq4gVR2WgCY8qZzHZQ/Y4740DNnOZkurWVelUBzCWyxE26utz7PrKAsRLB0lO
YD2UJZszQaF5c5E7Nz+L4pm5xg9LYqsKdCDatGSt9mpqXul91fvIzEtDi6tz22VV
OK3wW3yhMrasWS7iMUjKsiIBTRdgUPjycMr3A3tV0pxaKGR35boQzuMOYZeYsSGF
RRmcQv5XjDz8Varu/Qt/C6cHvZe2IARTs0ggTrR/fvZKnr47RCgtkyMsp81vEy1p
K12plcJTr+vtlFpYlOjU8rtsIXLvdzO5eRzojXGTBdjixplPaTnrx/43V+xWjXp5
fLD4Wv1XTwm2RGhVf17KKs2BPX2MAhgt9UL3SgofyXt3Q+uVcofus+pkMyg4WR81
XpaIxwy2ZOlEJVcHe8ka7m/tqdiZZ9wQDObW1TKIrZRJ1KddX/Fh5IACjPnKGPZM
zsEbMJ+crDAkP25zmSVttf/VqOUY5TFpgZz5AsDBDY5YQXRKilvj2JBaIFtG5rkr
dzPDjmzXZ8l7EIILCnK2+3cP6+5RpigKNspNXW5sRKQ5b9ZiLNltaBdA+Agz/g04
GlfOD57IwpCYglWtc44FlHAMTmotNXHu5PU/DNwtj9Cj6zcHbh+oKr89EyWCGWB5
LPW/GTbAOuqw+bpe3W1eT/uw9nZsVTyI2kHlRQSV0/97TzcrZf/3qdwGVFG+/vRj
qrvGJfYeueUs1/HHwMAcZ7zffWd0dR1DLaY9RirSXVRsce4fmKPKGE9BkPSWBUKK
VpdkFVTf/r3iCLy9tAndPq6Lxp8lm3O/zHHrOPSR5ArSircDE0VXm50+lUt7ivcR
cZpQURczee4egyluTNjy4gBKf3L11HifgIFGajXVwh26vziUxTe659u8NdWTm80/
CPRtd9nF9rPXKgf3Ol7/sxssrCqRsM1qZRWlMX5Nij6Y/kRffy/29YuTdbrlxvKH
1Axtb2AsSdSiLh9rHxzTWuVzaAIprMg/pPlwSkYAnZdsBcXtm7vvYnJAvTNmpljI
B3KVq5xhKHba5N1gDZJM9t9+Dq57AZ4UI073fPuP+5NWEQG7w7jktPwCYPmfFmV5
q78aS5hwL3f37HIaJuT9T0wgUu3DlLvm6+sleIKs+9O0mWz3Gy0MNydMWBR3J7jS
5tQTvZyia5wEymCRfBbjD0cc0Q2KTpzJIcLAab4OFZ8dB7tK5TZhnRjiSqKC6FWm
ZvwApmEBbVG/0/nwjBZ+Ils0aH0ulkQTzeCc1S3mIxoLh3XrCQ4sOPyH91bsE/wT
92A8FrnLO2KLgFNsKdzYP9oviaPWnlwm9b5dZuMXQwD2tnVz2VWaqdklz4RkI+Yy
8NI6+AHBV6uhHVD0nitQ966MBqlZhbEbXUUJbInY0bgpR1uRLsBJzKkOMjwYv2jN
QEVjF0IfNl5UgfZ6DrFpudsrO5NE0QF8KyzmNBxZJQc60Ve38NNtxCAG5x5ELnmb
s5bgo2fLgIlj2ovW0ELe10rfsu42+5WC9rZ2XConAulliuLlyke4P3wAvZbf0IZg
uxI0vA/JG4naxBlCixk8w3Fh1x0vNDLhZLNN+1BK8UnCSzbhBWQ7IEf/Bv2r/0jA
2vaD2M9NiGOdnDyE9Z/nd822bcvFMFBVMJSl6i6bKJVu0zclqqHitcQPqAB/jazm
Lmi6Wzy0tRoLSPl3ETXFFYT+ahG1w9HTFM/piKG5QlZrCMVOh3SR98YlYHjOpnX1
45FYqISqQ1Ar5WD7lJ/ZkC4hUED/kGNAuKP1BXoq5qJDHaIHATnTXnGAfjaUq5yc
BQNnKlHw4FNFtsqDCZ569RFiNHXDVF28fngY+bFxg/j8qOv+fWlTpquaPxL4wR+j
XQjJFvnR5Fg3rKYXjkd3d76G2z2LDfOJkVvNZHOZAe2FFMVqXydr+fPungWBEE3v
591oyHD+WCZolyGKe6M4ginkSgKHHAQCCWz5V3yT1oBy27ZT7yIKCByyuew80r8Y
9i6w0reOvF54elidV4cr4DdXn80c1ZWAbYOg+NhMBkv/fZx49xyDVOrEg/2HO9Zp
XyFAL9eK6+ueX1BaIr6hg1MC9Y18GUi5sTZOLkgPfhW5UCwf4NJaWAXTo3LOf9dm
Vm5M2zfrDJ4Lp1ZhuAbBflr22iY6zRlxq4xSLzkAK2xeSH+y0vX1X6E8HjIT6QMu
GwoMmTrJOb2Ai76l8zuk0DwR7CHeUpYhgGRdPLDy1fII/engrN3aFWmqF0SkQKfL
4FpdUFpR2xgDUmP0AakWrY78uXwcmP4OoJS93+gUnnqYq2EXs+BrpU1h7498XMYt
oz5ICc3vsefnkcds/UyHD/Deyl0i8rhUkGIA4ge7LdsalpbjhFLEr3bxaGvlhT79
tgsqZJjN65xlKWOcKYZKLVJZ87lFoyqDVtP9JLrcOzkLKZbrz2CG+LrxDr00rj5I
wuBlrNrIkQPIfjMaj8hMIlTFem4TMWKrd7O95qrHdCCu0xyIoiJGz1l1ILYAkDpL
nysq+S3ocTRelgmodBJnOGiGoJu+LH9Un8jC22aoLwrWEydF3whM3MHeOyC0KVqb
j0LDpTlUwKCvdUDoGChMyxfDvHW7c6pWDfMrJjQmucUU18LgR9Vqm3dLq+Tqc6f+
P1/5Y/msCqNQcxbAsz9dn5g2BdXQvBZyjoEDMoG1XfnwS58zl2fX7SJhiVxom6ly
jwE6bqXc3uJzuTGqYoGuN0fBnjnNZ/f5yrauopgIqLmaF8ufDukCHRaI6nWzXJn6
VVaTXk2+gANcEFmmH9LiWZ5/TcC7PGLOLjQnnq3xC+d76oiryIN0Wv2633QzvDfD
TfElPR5uJIoSmqil3e3Jiig0Ebq4P5Cs06O09x3Ms4mVGSNBQbRDqr/bIndZkhcQ
YtWua5jJdFbWZwhqqJjUXqTzrVuNvCyCPn95SP72k1v75HRaQzG68aqus2DgtspV
VgoiXJTxWL4xoUTSGeZ/gc6q1I6HLKTh5Gh8hyG/6JZXBvZ/k2IuNRV3V6FAnmK3
o6IVE+IdqhZzKEj5lG/PZyLIAqmP2Xd3Snq91Qe6oWPLHc4EJDsrgY8N4E+/g2Zr
LP9unxf9hBs3MvTVG805HEcxJ34zZ8pd6vLL9vmJPnoEfrvqRGQSiDmC8qKj/goR
mem8szh9WbXVjw3OUWrNsUGbg1SvVemgq76e3ZvNoRUhuFxGqkWGE2xLeCp5ou8g
Hb7eBcWQ1NLSU8dRjpteePctNyu7P7QUxtMpyaGjtzpHmz1C35IQPGcrBrkyWdbe
qy/SbHV6/OV7YPeV+MDy5YQFKj99IYL6Ov+KFPTK4nO+go5OZRRDmPstIt/6IXd8
QHk7p1EWp45yvAxQMn6yyP6R1vO1AIxSMekY2uLLID0yIkaBS2bjZ6ujcTgRIGxw
pR8iIjUjcjP8aB4IfItiZZWOkuJ0GyHGXLtXKJYe/j/PjKMUGogd0ZJDpWEtw3xx
K4foVLqG8DXYXdSDzRyzZzqPrL7tUdoUrIof/4fg+EgGOfejZqgUPDL32NEwRz6D
nLxdADdWL6S1vRI8b+miMrgdYlCxh7yfTYtA0nSXC8AFNVm87iYcoPTEdQ+w5FmJ
b2atFsqhFlsiRcWte8qpiJQn32oov0TriDYb7HjcyWXnk/lV9HlClM0XNC8nV7C5
pppn8d9yI/kDvSL2GQ9OkD+26R2VEVsdPKbJJ/CS3T4kBMMkT2PaIVrkgaLSkaFY
wHH1vJpUAurnaKrCTHNJ/5Mbm+WOFK4emub129g6mItI54EERpMa1DtMdBh867FW
sh0R0aGNXpx3+DO1xvtmK6NuBvkTVNbSMmEd2Wv+3BbPVxMQVLAuZqpn1vGvUIoG
eH3Vkz0IekDAZzkatVmjf+vR1OL4+YDedIuKeG9aqw3ibY7dREJUSKAJEsZTtzpz
1QC05BfjKRe7YwhrwdV7/pVXpYDYeuG3O9OT7ejoRR71DUHcfhUSKKijXYmHTdw2
2cJziOAb1fHg23D6qUdiNsS+9+7ue4G7yvWlJBqdKuXcMZQtAdbZPsvxidlgw8ri
sPqb/bLu62sV8B686TxyQjx8T4W8fGq4Bbd8dNvM0neimwY52jrBqHXk9VwNMYf1
ruJ2OkUNv5PDV8wGH5xigOvc77FTG6C2OUMn29sPNnNcZ7m3Sr1iRPLMkBWAd7pw
VqEjHUkPmipz0HSv++cXJVhrlj+McLIky8MMQnPSY9yIMWn1Rd3RYtawHg7VjDk6
Emfg/VY2QUTZr/y3mz7xaUANHZR1h6a/JdLE+0sRimEBmeme9b8UixphLx1wHylI
H3hJU04VaIc58gH6rIw9qpZqdeO/KaPQMuDVVwExcKDlYza7ZAU3tIsK3ma9r1Jp
P59Hk00Ms3D4LUMohEA/z3hIE/yEFZoX8IK9y7B5uSXsRPBdXSqyaavpub4gJHLx
cSxs4hRqMOseM1nzl76ZjdbGvBw800sRs67eH7+g+IG2FzVshL79ZaZXCbuCK4bf
iHTWihVRQ+d2sHSdtVVcteYgkXhcmgJa/EHc01USQgyQfckxGJ60AB83XWivzfud
6vy0YB4O6N/3/Ur/qk3KyobA7YqYAaJWy9F9eOEr2OBlBlkCOTh5IUO8NI+VdkHz
/oRFJW1B/r6oURyHQovMhIKcGBGV5bEaWDsutoyX63eO5RIvbCzIGpfB01Ik8puh
3UDKgQkkAxg6cVxeXn31HSYsD/xX5z90efd04HIF1aHYY2AQThCbAy+9zGKQW1ii
XYK7Y5idRExwUtzp1Fsgw5yTYhozcOaeEbY4TrnXDWA1/CoojIUn8ocGA8c7FdJ+
LQUJY15BFAYGVYnGJ7ULYu4mEOKjLBhQVKYUQT+mM/ess5r1KD2a+uWoYF4v6kBK
okDuSjlgiB4d3sahps6EZdYItMOJhaNBvIwIQHA2MJ59zDUAf87WCrRKb2zm5kD4
/rYfPl9lJnz3prkQvmAic8Giu7sXJDCcexmam7St3D6TTzJgvWCWtiUFUxZ/tQNO
W67ktUSptEI8aAUg7oBQ9Vrja8Nhma15uqnUkZh+vkaPFKRq8jF3zb9r1iYq/BRG
447NdTQKZbF0de+Hj6SJ/8kiobXdAw7p0v+/wS35Pg4+OqB+CE0t7yWN+680dk4b
ybpWn+os5lJ3PMvTKV78siCtvKpYaP2EsAz+HNhxkk86zCj4qBSa1bxJM2RleHfF
XjqgM0xe6RBg+GB4n/eUkDFMTrgpaYK82s6m120ZJFCh6SEYmZjmaVyQQG7erz9h
DF4fYYBchZgy59MBaxSF4LZbFqA6By7AHPP0Fr8pDa5LaYtqmdDfsUSAUGTCw7mX
n/hGvVYl0LfbnLyAfiy6x+1soS6hYPs+qctWSUJDMnkaDzlt95cyQQNDlKYlVoFs
V9va+ttWSSPwd9QUpqXvZFeVTOiT4svVy68MyOhYceQlWTlS1rd/QdbtWUBZtApR
z9c7ntGY8oL/lMG0KKLK3ZNnCWycQKOxkoMwTWh5YWN0I5/JdnEwULGyxM07Xd0x
SKCEkLgdOZ0V0qD23a0/H9ctcneNM677ucKd8xQhq5RuM7V4bEm7LHyBpSfyXs+/
kcgNAbbaCmh8N+IL/8mWstz7Iu//te7d8sE0XwiH3NPCTbronaBW0R/NGeioN/LN
X7N2a+woSW+wMcBCbGcP3OZBjECvbK9e4z04kaedCHeoh578xe2sP1jZxpkIbRd6
JS9TlmZR59TNmS1SVzL+9/mHtksK7acU/JPVqxPBdfyYra92intD+qqzqeCO9hQN
EkRoxP8LYzQJJqmNgIb5/605D4l0oxUHLj0FUppzbMGkLnuhykWguwjsRgNclYUp
4R/wNc1iPPupgvq09GPl7gzVcaQYoG0DvArTNRR/8qJgXUpnZ+w3NQrwST5ZsitP
RDGp6/oRlfkYKG/2skCpnkxwuDeS1I6SWsrV5gvhXEiQ9yF/AzhAxSlDtRnoa6KN
No1jZnzLtMS320e8nOMkSpshI2rJdKg2u2hX+vD3ywPmFijIKHl3+T9wOCSJDDcH
OhEFAPFqdxFoXGZ8WkvG+Ur00UFNVViztRNXmhU7gNdtiIcqApRQP5+V6SPRhvQt
Bmiw9Ev36o/eq2Od+4gK3wHnuaHmNtps/Dxm8nqgV/YILKa2O9nOGmzwNrpQMCw0
z15oFgKubgpL0OnyGtXB9OMkM9bD4uxeRgjAKa+eRxpuPPSFt2aqiRXr3L2gN/JP
5TRNDFdCr+a/1YVcw/dycU9h3VQxpOB3RZB+mvqBSAufsqnfRRonCVG2fdn5SHGP
zh05xXjaeIhWM2BF6NXnYsAPDV7FyXKc62pQs8evwvgIz8vhz9bLvDNLibyO263B
9IhrimhJD1d4ieeypcPMbxLCEfitPZ6/+U9W5omxPtZb/w92hh58G3nYmLXEGzd9
qshN+J9puVIBpC5JJqv1FLnDXtuxeACR1b5+KoKAZOLYWRUpyZw4IG2kz5116BGA
OqZGayGhZg1NwC/05XmYRHhJ9KbDjjtzJ6zMDEXurpZ78Tik8XZM/GJedJb5uVos
XgnbnCQiw1IZgI2PY7Kpy/mqwU2lwiRhV3YGfGjSWKOzs/LheNn9KyufEhvzH62c
qpquV5zpdT4OCs0FNF2+GE9HE7B5UOMtBn0HFH0G6ng1QTuTdW8Lru8IHV0Tf0i2
RKCot+1A/qR6HeJfROEB64iyf8POjFvIuPG8WqUOgcxgeDpHBkB0HdEXosIZ9zG7
+coQl1rehJVxPoekIDHPFep/nPJ4wP6MJPrNBoGf7Rq2qQL8Ha8uG64zO0CIQCGB
eqw7uNngGE4j1b6c2/0HOOW8wZtEQG+Gh6czYGzq9cTGhAmWgxx/I5oOzHnXSpN/
xi0Lw149Ac3Sjwyzd5SOjRL9VGwCnFI6vza2Jr9YkWCS75UCv0qXeG3uwZ3ZbLI5
+brwlzj8dmhV56txH5BGHIzqIdUFgAzzfY+zp7Bb3hS1bQ68lqsiu0nM9VVSn51v
bcyICk4OQQSbmiDmNKxWoIPDUyuN2yL7I5K4kStpMIVO6sw7uCFVBtqeIKKvPk1r
41CjQadBFLSTIo+MTjudxyqh/MAZu65uS+tpBCUYZs0JSwOHddOAKlMhfx/Lpn/6
xNYlmOGqj7P3bOhWHyfXc7IcOe0p6wB2uU9BILCl7CD6Z92gh3dk8Byk2FC9xOQt
2V57KpDcdleJ66kPDP7WS6ORxJCfdTmY2ygvFd4mqKyaAahEaLX8SODMFMnwbUAG
zDEWYQ4akTddZ5q1QxCvCrgNGbzrkTOmgIggAyXhECs6sbeZn2OTPLFLlpue4T24
Nn1NakM2+6p57590d532Ym8O9CkojbKFlLQw1wU2nVtUzuBAay4O5K5d67URAfJ+
rOXOEqv6ycGIAEoVJB9fYCApOHIkUyuuMxCJDm8ntz5c2Ha/jK0WJcVKwO5X8wDR
wDonmQdf4MuHo7ZPK5ZZrK8BNgxBpz0xBYi/L5SOQRaV1a2LxUhTDSULOKhEGyjW
niSDEPFkl5Byw+JaHoMrR4uMH2mhktRX+6IJNK4/eyxa0PDNnYEclS6i24wApopF
qOLTT1+PKtrC1rB+2j1BhT7R1Xi2sqrE98WAdKyaR62Lcy/sMkSByLl0GS9rB6Ev
R5ml2D0Bcvz1FVzbgQdQ6YdGSibGCWrg/tvBoPLQMyUAMFOXF6PhD4hkSBNA+ZhO
Y1Z+k2LCAMQtA+a/EaF4R5UTgxX3FxZCLvBGNwIbk2/6W6CkGMpsAlFkhq7UTvSu
9suJ3CeIq3yHLg1P2ysW8E7oUVCwT97jHDgloAbarumZK8smPkuaDhgzOA9Fu+5J
zOE/8g5xcY3BkheF7AoNTyTekkgKubHYn6t9WsLMizkmbP7IY62/13r9KtYoDGXV
MJbf5hPxfbimsqYzHeHFp+q9fYqWVbxx2O63RFOMvJiMejJ8/ub0VTBQTnhDRX50
h68vzv6yfUWXOMoHzXCTZELJNg7tkLPKvY3E8JHjyyiI1QezWtZac9WSNS7MWtOD
NxaV9FHr+6yxLf3LqCl3fwP7Rme9WETDedJgqueTdXV1xkShwXHgUl4b24E0DZ3K
NBqdV89PhANIN7ekdH2ogNKi0U4O3XnZyF/DAJRv6af+9vaSQCXeh+ZvSb6jsTJ5
WJNRhoAabGz2PPhTmec0FOeTfjZNtyy5jzUAR7IYIhgf1oQ+3wsYCQEwfOPtGhOW
7ZxKJVIAuP8KNscS+VDhU064yxHYg/DmVsiGZ3L0fekx/jFAMwwuZKJE4mRhN9+6
kxTprX4ytPidyA4hdD6Frd2T5xEVCW6/QJnMJWBlqaCFlAPgnaaqm4Nfw2K3OVLb
uKX26NVfvoRjUu8e/oiNBUfKsB0SobV+rrVRx9U+EwdYw1laFrLxwp7ta7pvCHhT
MrFT0uZV6jQJCUOCKoi4J7jHC11OOsDEg/575lsdIuzifdROMf0tfH3FnfOWRPF/
a8isUSEiYqOgmnP/64C3ocEj8zkImoIe+PC6ZOC6wxBt6NhDEnD8ZnLkF7NFcRuL
KUy0pVeFMfiuUjgQvMWL9hN6k1ECVNCkTgg5CPqRcxOnRg/wJyCBoIUoT6vjvJyA
oVvHV5F/xsrdDE6U/wSDJmboGp9KDjFEWnYdunoyd6cwKJxZNk1ufEZllcwL9ZD0
S6c7MA0RpVfRStGJLWrUTkdRwrhorTaaMr1x8q303l21JFaJFpRvJ4DpCDlWIwxG
MU26AhkkvqBHNjr4k/Kt+K174eU2hUgXyOeOyYKkpBPPcHLF/9sjN0bxi6HVajp0
Df+HPEQBamnjQJnePvftA5WDqc1yTiQ/3fudQhgXvBuzOB2bhd4e7qDltIH8//2h
YWL00lJcUMA8FZ5RnaTsKLd07FyAQkYwATBdOKCn6j2z0/17ydLc2YwQU1hiVO21
uDX4SNmpE6MMk+9SNI4uzXjy9yxqWNOk6YfDSzZuCHaa4d1D1Km7rt5J5Ikt9Sqt
47yG0iQqW+E+c2Nt5yHy6s4gl36au1Y4r82M7MI+0nVfqlrXnD9lH/+ZxO2U6jIv
4+u5DRDnQJeB3bV1RWulOM66tDfIgvfHbd3vi2Mue/zPwbrGZt8ODr4PE+mgdCcf
+ngqldFLjflvOsJ7Ew1T+CuRNGE3YfElDN4/tSb1ck7EnImzphHdoQP3xE85w5qN
FHAozKvY0ceoEx6DVHBhKQjKI64T5GbmEJDRfYC1C9osWdjUVDJRhiU4VpKji9Fi
rC3WcnHfE+BWcfmev0Eplw9dyt4VoZrnso28++0MxU1rTVx4sNxcY4nAmmrcExp2
Xaj0jf3Wh+AssnszAizX9uVJt0J7LHCFGEcULPa5qGvUiHX6qXsHIVUrNke04TH7
jkrBoo78o8rsFTYsZtVB8XW1b70waDk7ocsRJiaHogfTqg2sDOF2QUsMU11uRJXa
lxAV8zl4lQNt3H1Lb33qr0sxeoCtrRsR8zcvBNe2FcGJOjUzo1YtYMlHICHFcWG+
5Y7F9qO4C2Kcs3hZhDxW2jEdDYvIVjpildNcRDbTvt3MR/YiNT5+aokaMQZjJL4c
Wtzt10O1l+OKXkp3ncrTjgOzy5yRhYzv28ZHNMJJczfUcLUVgiwqIxLVa28eQZFn
0TnrEOwzlhkxKZbmQoVjQfaz8olAlUB1S2fCPVUrfZQo1VNAOl1fffen+vDbwOvv
zZzPLx8f0GW3RKAlBeUbIDy0BDOCvozLclGLpQFWctGa5RAlF89QvBbRpXt6bgAE
Hq8RdiEoy7rmiQb55mByDnQTaGCgBGJe5Svz4DvjJhewiIXoTv1q1SbGG1YSwU+Y
LmxOdiCdcv0owIWMxHVAPzthV//+eZpK3yc2W3qL4kjK4dYaMlvN4iZ972eudIKM
yRVe1Rcln9vPWqNPKUn1XD28Jw7M8pASgcRWN6Crzk6oXRf1Ln0+sRJEIu1bikHl
80LyW/kFTXm1BGe1KGI4xi1dc7gMa+vg0wQOXsZi4KpdQIjZq+2xueFwvsjSKSC9
aG9+eZz3bR0ysnRo3LEuoZCuWZYyEkRjfVF197rqMynHWweYlcf837GncM7Dvc+a
6INAkW5lFf6wKos/d+puvPVuytyEo0+RR6LpNb/4po/VR67LQ/EtftFmm3zpAX0N
RpHzm0ZXbmHzrxnChS7zCVK2k/3uh+0Iwzwdl8yMttlcRPdJqkWxFiOXWPeVNcFJ
jeCFGd33/+Z+OqDEaVdQY9ufkMsSCMlzFtM2kdnaRfFFL1nVNFTrPgIUn7h8C5v4
C/lkBLpRspHrKpi0amnPl9q3m2FsCYHZs//7E42RqSINA3J4hV0niuCDGl0PAsEf
N7AVvp3qiYv4im3Sttr8iJO1OASpm3VrF1SpgmL0V8lID9dQl3W+a/5Q4FR+hf20
kzjnNv/TVAGNxEuV1RhNLkdBoMrj6xxLuaFqF6N5v2BdmlR1e4dXe/4UoKIfvTdG
1j1UAIdC+140s4Yl5Disaeor3rmt05MHpdT0tANnfvMpfseCj1HiSTD7xmTWySqN
noiwPG3q+5gH9D6/aVq3UYkORGBAa08M77G17fRYGNpGIRFUByo7MBI/y+1/M+dA
DPx71VVE+f0nlba9tAWxK6HIUG+CN82dVdZkDU91aeSTizIYWQplU6fT1pQ3K0Mk
RfT3klTInouZKOCrqnoqc2lzDywctWgCsfkBMQG//UdJAe5qKkzSXne4fcyXoBBP
xKqA2i/1e+A/GC3OQOizdwTicQUiDCw7pESKCjSiV4BUyc1lcCO++X0P93pEPQ2S
Q4wQu4/qrDzXHTmVACVvzbHtrHdHon3OiSHB94/Yvlt50dXQTmZwkV6/8eObKcSj
BfM8gHi2XXFYi13+qcvDniDEgTO2YYiyBuKXWtslNyhUuTsqYxBnJHjTgFv7wy25
edks4NNmzj6ly6xktgUhUKxJawYJwZFyeiVSs7WmWAuok6X0oSQvW81NFXmXyZxa
YdOFKhe3MPAf34SiREYZV8G7WKcouDoG4NxBr/2dtog/E8cx46VpbvJAq3Tyevwf
MsCAGlcPeN5IphQrPhPTQORzXQ2UZHJp+Mb6MM5jWA1nrSCK55fh28Mw5RZa5NS9
B7vC1NnCDR+xqDUyixaZ5yTsQtraz+NICIcLGh7KyjzjZiyA7OCHrKpn2VB3wkys
jAp3u8NVbfcCEH0u+A7Y2GeoXKT+Q41p5zYMikgPbUNlzSTi0rWmH48aEwWEVtys
d0wFU713vgPuUDK21wyxTGKtc+lLXPbW14OtTNqtXXwIQ8tUvJlKrC8hxu8wgw/2
G5h2p7rwMv8irtMUUYsqtkdj1PRMREiF4jogvqYbeJPCumGG890CiF98ulszS0fz
/TgrXLFSuY9LcX5g8ehzgUzZf34hSNtd16YrPecxe7Nr0h6QIiAJKqpPvvvDDN3w
d9CX2X70xJPLbp2t97ymVHjY0TIK6uo++K8NCK+k4AVcCVSxnopXFwM8LEjXjtx9
YZyumCkKlHf+LTjO+0YJxrmTLoHJzs/krKpaGpiJSl7TqKcb/mKdqfvndZXRUSa7
4W3p//V1pV/s3oukapOoOQFKF1iZ55qV7vxNyxdkk+F9MlFoDepz7RotfVL/JNFD
kuwAg7Bhh2f+NSLlolTDkDgnWgBnLG0/+fRw/cfKGSxRioHBMor0UnJcpD3Wo1v6
+h2+FQjZjAvY5H92MFwzBF4y3xbPX9QzV2rCUsQdDK/xh1TGHEGPp3NGFXzOwCOH
mqMabjSgitiYWv7/Rex5AWalbEncNbVEIhqCt3MxtbEkem+KJ7i30oejaTZG8Q3I
4waO6CXKBcu7ueyRC1S2etT11nW8pWfSVTCpkt3Rvv+iW530x3BhQOXFYXtN/nC8
qvtMn4I7IEqdesxztSjk3zXfH1QGGTXBIpc15Ijv6wP6om+Nm4tagbKnQacsEk57
C9aiAcN21tHX0+jby2pHYPeNzMu7dGgWTsEHTeYnAU9ATO47vjCDt8oF7YT+G9A1
6jV6crcQLsGmMmCpz+aSnF8uZWzYW1OD8p24mF3CvdN+g/t5G80n0t5tjdtDwZnr
WHs77dq3Ufw1a7BbA06Va/I/kmfu4gVrdq01Tu2l1qt1Eyb4PdwY87m8nKLb4z+M
nehmtKoLeP3Vk4RCQtPtKNnDUP0jasBZ3u1dy3JXdqagvdQWeA2DYTEB+NlqXREu
iwjTnm08quC2yOSE7+7j38T01hvcttWq0Uy8xjLmEqEFlDvI/2dV/ur+RRNRKHzK
ymTOWQ8JZHZZxCZYkT+2286XeRXNOLGlLYEosIeNJMdCtOq/1Z3paCyue+17kNEl
viu9LgZjIBkEpr64skeiuevJjaJaNObF8WOBwRgGOv9NVXHe67l5FId/mq55PVI5
91zyiNqdhNuORSbQ/jHBKsGQStkwikLmSZgvPwoMpXnjzdZbnROgdV7Lt3eoF0WJ
C5hD9e88LfkMLqRdu8noodtGJGwWhXoix9MH3by43iLmQW2c3QvUhge8Us+n63fA
iB1Asvk2EYmn9iRwpXs3VPo1i9NRfc0pZND8dsjLH1GCCX+cR8lRxhbqMJx0wY8V
0OdgUbBqZ+D/pL5HViny+vySV9uUT/z9IJI5wT448ZXOIHl7kPu6L1YNfhX5cSBB
GjQuVXpgjkcUEDsjSrX4o17oTgwP8lD1Pz+4fshkGFP+UU7LavrPC+buUrMvEFAl
23XdBt4xAjF/E4qPZSjcwWlg6g8Yk0lEdL0cIRSORqkNAsloIO6GqZx/mHksUn99
2WexagCbbBk9ZsZnPulcflXmx9XM+ApQp5DoI2A3/5+K2g/IQpPUZOdE7kkih61j
MLkSqzXq5cI8pAclMC1pKI/qAqGvwIdziIXCzjMjabONV47BM/GT4xpmh7J0Iz0d
vannip95ktZpNMsnM0GaKv+hSh9NkemJxEjyCjTQT641nOK6d7ejUtNKPB1nZCSg
qeCpgTwGIHAfExNdEiZabe8Mc++LAnN5QhGynfjrXVVTLLqHz3HScYWumOm58rjo
WX5WW0Lbn9Dcu60/SwGt/0RniWGgclODXeTwgNecXjyLIBSDAQ5sGTjWS9zmFimB
s5KrskNGIg1maYDKL8g+AJ67RmPq47nEq7MNI36wTbvpJDJ4fXNU20qJT1035VsZ
qFSOscoWMtS9nTcy8RoyB6VKZO7egBXh9EEwaEXCH5Vr3RAnCjodg9YnGrgT+H69
74CeKCB8dY3H0+IQMQshT/MTnOfE0z9DsxkTmd0vasfHarWGQ0OW2LLNTHsiqB5y
UjtAZOsix0WWnLlo3GPOUhV6OOd5sC6XbP/lRXP4Ltd6++om/cof84HulHHpWLRR
8H60PvmL1z7xparhRzXtMGct0S55h9hR6J9dAUKszs68Sxji4dheSQ8T9531YcTN
1XJ+c+S2McOqm9QVhi+Ce90LC4I+EBot2u1BtXI08fsnkbuVlOh/M5V53AMHDan/
2gs5q0t3q3r298D1TdTk/kPVOFePGAaSC+wZhS/Z5o8ZaC3XUSzQGNyG730Jg2mM
xdi5kEoMrqeMnoVgp3A4qhBicmIY0IEFse8TGBmgMn0xnyC/kIT6hAMBx40NcRAB
4U5KhOdCNH7tclnPFACmnDh4L+pk6fRd8rDkDF3jy20SUTab3JyNfdixywoZRYkJ
8flV6fHE8PpNhpCu/nz/Q2VBLmh5Xzz+thJojqt4ttn7gVjb+JgeAuyVNK3YcU1A
GgtOuRnUpjiz7SXF42DQrd06/PeNLnBLlzJwXfOAub70Q37lAa44JCBvV/557VaK
NX1uQIU1Jkw4GTFgeZ3zaKCoxsg7gWoEyLHx3W7QmbKOv8dog2M4m1/t/4Sfy33f
9CfwvfmLFF4e29HmnmVtS9Fy2e1cZY2LyTqnzjQgaxX39bJjy/Tg22th23vecYHL
7nPuiu/NUNqk5N4as4f6Hy5/JFGLRKowco5qeTqGVNnEFJlMA9chQW8BM7Pl/b9g
7MNOJbaxJDm6Pr/N8KfH385/3bdB8yI986pbwu+cVihLSxRGoaW3S0UP3EJGfOCk
ZD/tp6s4fiZR74drWevT39ov677T/WroObxGAB777/bJgLvASSqToxY7T2LWP42I
0wFkQF5WKc8KzZ6MXr9pBYIiw6R38G9ZWSxnKjk2WAGMNhw9F6A9TZDIPgTCDrnt
txTq3kT3Cgdg83n3CkI1tfzOsQqOb3TIalZnevWwWar8pMlhGNAdqs1b54bVZAPv
2RISBOVeZsHIulwuc0V6ws3EThBijsCiZaY1JWHzSGMwzTqpLpH2DfylLhqH53Z/
U9Pq2h3wzCpByjZp1fvIZ7KABtFxO8CgZmR913uroEavGPwbmSK0/hSkP4ELUQcR
LVGz+2w6bxD3NQyj3B/jYJ3nQof05q+G0rWNfPrxVZ/CFF7nFh6ZyBMrcS/HwV01
dyOEB50YiP4lovV4eDMSXzuOtjXhkJRogQEVc23OaAa3a5wvJZ+xVZJKpkfZq3Rw
ec+1on6J6gfPNdOlOnRM7jU+tVBppJZNQqn2+oQrP/8zL/O9lPw9928F4M32u6KL
E6pLku8x6bOSmaa7wpPo5A12q5j+tqoJLjh1b0cy2MNW/qf663UdDgpPXhEUv6n0
TTuV7n2l17B6wNEAP1YI4TAeJX876gKreKewErsPNwCdzgtW0mDaxNj6fZcB1ntV
uwE4S07h67JBVlKPu5JIiJOTd/AmkqCnXmI1lUr8uN9/weUb8VfqpBd6PgzGq65B
ubcG6jht2HT/lxfB6bkSPE9ICsg+jQmfJOUwTj1T55F85AwmlILknGvwpi68tWIk
HdGtPQBQnJEYHf3si7gv6Df1p1s4XBIG3fpO5IRsEcuUEM5gwHeQR2KbLu6Gls49
4odsKyrd6Z8FCEV/enj+80ty2xH/xQvjmiNknEt/u+IpIlS4bNBXcY6BbnKXGSLt
Vybx6YfLYU2xGsAe1Sn5jEdRQufqQJSu2MUNPai7ULWoYwvCeFE5/1UYtbQ+EgdK
kgFVn6S8lNaXgW/ZqOQvGstNO8W3D0jFXC6eGI7DB46UWIW3YV0YeMVpCdFnBmxe
Zk2QszEfjlkQrTrwzHC2JJMCDziBygePl4+TNSfVxRKHz/95dQ5/SQ9GZCGY9mtr
D0rXXlcZmrnZ6LuOIAH1uPM9WDlP6DMXSp8XYoUVOL1Vh2bPO94J3JiReJdQYx3g
terEqXnGphol06fL8iYOTpv9EcNCu457pHzrZAnVHSRaN1g8joHHwfr5ImVXda0N
stgY+aP4yMMinaifAHXT7/1DDFvuji2UbnLKA8kR4QHy+5RyHHuW1eiQOfKzVjRd
zKcOMd71rRh5UpZwVuA4h6F2huf07+TLjkiFZNWTKawFsQeg9A47eGWZ4KmEa20c
zigvAtcMpREQyoNLgiTska9fu9GoBkdFj7Ec/1b6YLphMNzL2ilNKh1HMiptLqKQ
8NkMX/G+lQXrDO9n0dW2vl6mGmtHGJDB8mDaWYJm5GQtdaTsOUkIOPTiMwnn+BNa
jugoeJYYDA1/Gb3W3r4AZqujjuTKzXGRTjbgquysz9qfyJmuD0rNB0TNgjbfQMz9
3QxvQ+tBnvdSxvZGO9GhlWVIxglbQU6XjEV2zpSsUfG1wmQZFk/tcoSbgZg3RWw0
CoJirkTPgcp1nG5tNgrb/HNtxmyn2cjxjD4EFds8EtJuYGcMeSuANwqspYndzm5b
e8Qlp8Qr4raySAAUfKrrDk5gPVRQinGwFhJtqybjDeTcbmB/grdyASDodyqWsX7G
ou/frrMG3P0/5xmhhg7yAVQrKcvUXrQzHvvZFrSdiL5P2CJUR2lFSD0r71UA10Fm
TG3YmN6vfaEgqoGtnZ/52cn9HQc67yHBUraoDhmxvFGBSYSbX6Ox7OlQdAfJpFob
nAL5JnSmFVmYmD6h20tbzJhWCZe0sejYrbJVHimpn+bdZ2Y7RTSROnBUXDAX5qB9
ZGJVQYfoKldSEiZWwZ9foZSVVCyFuF8KLRoodvYW7pSzhpeWnrLJnWhWxt89RdFO
ojn3IZ5MOOYVSXShk1FS3923kTpgfR1KS0noDoQ4qO0aHf7XAWa3zl3S/u5S7tI5
p3zJSxHf73c/k7amJe/Q55DqXYd+2j34aLrKhccluLzEuupumrT23bCsjEo7N7n3
RR0MRtewXe3qzkXxDF7UsObcIDMFCrnaIw515am/Z245iBRhO2mN0a3Fao1TUbVv
xNjvCu6c7ryun4BGuOQ7VLNH06CYffVIXmuiDoKWr2claHP1aFp8sq4FF8T5tQHg
wGyVIDXER+XOI7mTIcY40hLeIt71IUcqQBgr2+aMbOpMO6r9kY2qdXfKQkezQYb8
o/wlVGkYbAOlGra4z9+npkW/pBR3BmxoEZ8c2OS4ivT9Uy8Y5MMQ0D555lG55gfE
/0D7YJzE52gLVhmXIdicy+NbZrzFDZbtKPgMgiufIKjcdVYkyO4l7/AYlYSAlrub
3CXhhIlqpv7svOvkeTA3gGJGieHs5W4bvrRwQ6LbCJ3RHMiM9/6d1HEAOnwLWifu
8VcSUY2ce9hUkIT+LPO6OEL/QC+HZeMKhvphL0H7mpsG32InCjNa91aSJw6h7aBS
YO0RgZZqt3YPbSfPQabVh4e1CiCrs21jRr4I1agsZtPQepwCBxSW+iEx386EXcWe
OtQLwcGO+yDhDJ0Fd36Bw9wTuJzJLp97V0/0IyMw3GzHBmPJqKbBbay7iQKhT9ih
P2JskBzmz2HkoCJz1I6iOpLg5eejPXfeyUoxPIsQrlrDtTE5WYEzMcdGzfxnq3Uv
pdUfk5vpAw8/WBmnUvm8a3DXPcsJqKvgimPT7zAmC+UpBno7xTS5GerjwxWYDyB3
z87hzZweBHa7e/z3+buSCx/daCOPnjcsGfazmRHHnWy1PNyc6ssMLocd68NS1Wrr
1Y/j6lwC2FnDmZaiEc9kIwIagAV+++QL7Falq6vfxF3AQhYHs2HahEaNmzMSNexQ
S3zk4a6sZBGB6+zv/C7o14ubgiKryfu4A5nK45oTMsiPVvcvTem1XG7uh08gU/dZ
D3S3DeWn4o7Frf40mDwTrTV5QqIoebtgEvGxqb/RO9bWDKce2eX4xnu81njWTBOu
MjR9tDQsvk9hwxahXT/5XarkZpE09YRBnmh5bhrz2pADfkPGFUHZh/JxPeWheoxH
j2YdsYbV5+NZX72ZDshfZqznaIPxl1YIxasUAvuLfE2OU9aFBKeSc44nr6OZ9tEq
9Y5UnLYmRj62RGFto2Vy0aeh7/qZIMsFASrR6HVClFa2qhDmogHYj6TRsHpZ9d5n
l3Hflg4Em0Fmwm7kcGAETXfwkeftQHEZZZoWgGiYQgdMWCdl35KRt3g2G1sASpQL
2I6J926oN8sPH69lf2UoK5MQrPa83+ctHbhNDOM8TkJSo0eyaiLyBzaz3bn7Sbcb
JaAczdrdY0XV7w2JoPW9K/ue9MLjIBgnF3kQZ7R4EZmCG1Kjg6YZCSSwosiHOEV5
lX0PfExzICNdA8wwBNNK0HF2sZ+ZUS1x1Yj8J2X7EIFTStUabU8tQZjKGq2JcX0Z
wGakKdH7mDmZJYu4Uk51YwKF3RWCKcMhr/+NZ/e0pH1nDK5scT+u9WWWn9tIN7ow
B6+UYoECDQHFWi9+//zu/mL2wOG4RZ8F5+M5CkFsJfYl5MQ20V+vLhFEx7sL079L
Axrf4Olpjano9g3r84Q53t0qhQpMkI7yU0MErO0p5iK8z+qysx6zC6CZZM/RJRQ2
yIWxOzzMM6CNX6n35ZsGS+ybyVPBz1c1wOAXwWT0B03iIQESUZyiRpL9Vp8yZx3f
KDm5cmjPSnQQdHvu2DKrPd4Lqt9walp7iu4MrOwctplWI2aEuSsTK2F9pSiXFNl6
JO3GZ8ApByLT8zUsQWF/lLK+ziaVCGvrEosGFXEWNPrX/mq0g9bPNGBJKQp7AlQx
L55hgcGQeWCaa42kf96ypy7o13oxukjME2707U/ucu7YejSLaqlkd6EHqoUAHnm0
/iUnrTGP1XPHOEQeaR2x0cIMgSWPm6ZnscokezUm1L7zCizYVO33Twp74r0wH1lP
EEO8ZXRgi+Bv3AS0zmnJRIVLe5BmrnujOYuXB6sXcn1gZdXHeTNTs2pIlJICOtjm
DxcymR4iBNktSYUfqz1GnJ2WgXR6BaleeGyZEPix0RgDrWz/OatwHxekkKfG/Aea
JjbM7KuZMTXrfFSezjGhSkrzJeTIQk2/U8lH/Ji35iP4WhzOhQPY3w9e7nHPUKWN
oFtuRmcc7VFki0/3dAmm0ujr61nCNQQlGhflZPw0IEmusQilVEhhopT1xK9mVMCi
0mvInbryI4v2wSICPvumtbdWKwXqPbA0AFDtRIGtes4zTmHJQkTzI23MpmDRUPTw
ewXwRgHiBysrtBv4fL6JpGGJHVyoKpBBf9AmrwavzZOxEO2zQG9SdiddJGNXda3P
Vx9JJi7VqJ9dhIIPAizSZQ3MH47BJ9873iverpeEhWkPJxVBOzuYMruAZVdOCsTT
ClpJXpX636Aa8LeUYbuaUrgJjfBHB26rM8nIOjLnsf/TX3rnDObJRgqPUlPqDXXe
ZdchLspoJpEwXhMv9458a/r8G3ww6OI/04VhKOtj4ZjvLN997YIbb9JxZYGfzHDT
ebYbpTAwvl/BnElp6rZoqcjGQi/EvUVNMHUTwjV6pGnYB+1OjdQKVMDaDt3+AXMC
NMaoYNRxxgY08tu0L8cev0YgkqoJdVTciP6TJq01aNImy/lqlgS1ol8N0cReojrb
jURnlgVU1To2SWnphc03Kfv+xtsRnTvLobPiJDmvENKYowLsFgr1Fq3cqZ30IZbg
mzcQvYOoTt/0MbhjulQ+od7G/odHmcv5P87FkoXyp0EJpGZtlXt7/mJus61A+3zE
zjEhoQ8ZVT9kHarj6JxPug==
//pragma protect end_data_block
//pragma protect digest_block
heWzPl5Xk7BiGnulsYViiHLEPng=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8PFsDnrx2JSPs9xXsvXX20nYpvQj5CdGCmlWx7MgmkN7MqiW6Hwxpd982KQlLJ7p
536owxPEmnTahTp1k6YjMi1/975A7Mk/2IHdbmptRDd0UfcEhekIy9NIpHSX95NX
/ej7YuWA54dJVKSSHPmYPxXFBQyToZcMDAFRJYJGqshWSa9gy8zhWQ==
//pragma protect end_key_block
//pragma protect digest_block
MbCklVDqCfl8thwBWUB4GFcUsNk=
//pragma protect end_digest_block
//pragma protect data_block
LQKgJQ7iAA0ClII+GhiV6nOdhoXOg8755Z1gr0xsIOZXelIyeIbv2BbxgccfZWKL
uddxzX6VLDQ8srB2gz8I2h+1qRekIUVSx/tyge6oEbeNILqBLjt6jIxPHu1GtQ2X
Tj3ZlxIj2B5k7lzBP1oEBqzH+xPdz/9Sq2csS1UcKMrbj7bG32LA/9jfOW8IDcYZ
WkX5v6FSUyqpOdbtI22U5EXMomqRWx98Q7oED1/L9qRz36NA/yUZTfge9sA331aC
rBzLQPAPiE6n05fHfM2gt/D15HiL64Hmdls2MT37g6AwPWTS3i+PXtKQ32zwNWyE
zcgJDNPE6Aayjjn2W2ANFTssnbxk4Q+uBNFG22zvAYY2QIT6izaNUCG7FA7tB+Pe
kMoJEbdB9vuottfjfX7WUAdEYcFGC0ZKD3KKGv3/o2/n51JKUtpQ5pOvYE1cF9jw
LIiyCSQ9g/n9IJNP+aujfQ==
//pragma protect end_data_block
//pragma protect digest_block
ODXAvHoxdeK4SfpP2PYB5DtLJlA=
//pragma protect end_digest_block
//pragma protect end_protected
             //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
sfTJ+kHjKoPfhzaDklQBa38tpoWRiVO+DTH5hKBZ/Rmrjppq0kzXKfNnE/fqtzgX
5boOxy4GKN+BJSKEDKMPbPRzuvu3IlGqSn9qeLJ11HTVmV5ZR8OJ4vErwsaA6qW8
ItCtGvez87WU053p/083yxki4dD2SZJ2qwJ+Sir51YZ9L4ur0Bq2TQ==
//pragma protect end_key_block
//pragma protect digest_block
gCg70PdqUznXDyjOeLyS8rEqJA8=
//pragma protect end_digest_block
//pragma protect data_block
LK0yqTrL1qYLGSSKvxKoMHdN3zNWMZMQslRviPqptoyrAErKpuzSgwwBmo7c5z8g
ipIi5mwrqy6UoD/MZLgkyxe0zNKJMHtlI/59laYpPJXPey1E15a3Zc5rYYKwtgIt
q3nxyyxPi7m5X2X5gsTo6Hma69zZDyB3EX6lRS661sncDRY0xvxYpWaF9bIt50y4
gS4cmC96HBvQC5RVSK0ISPNYGnZlq4szq4JYH1zltz10uUSCKx/8vTpTOqC2k19n
GmhFZej5H5p+/Mum/y8JU3FoTyhSTIdDUYvCTyOQIF43kUqr/iHZNrnOVi8JKbl9
tsRDeaDUiNBzhlqq92XSm6xgsAFqBJRgoUCj80llGS1p2K/dPFdf9PXYFb5Y6erm
9ZgZXHOWGAl8U65yoRlHZxz2qU8Nnih2l2agJrNWq+2xUsqrrfHtpA96S2GJYQnk
zUOpjU8jZg+7080bqCR2qh2Es0kUCkmb1kNCw4+5l4Odw68d22xdRBIYtGeETjOO
G70aEAE2aDAiTklapI5C4poEbee7a9EHR0DFaaiAZADeJ4nEZNKKLQZVawLTWl6i
89k0+LM4crgwXe7ZEml5gh3HHEwPW84BFq00WqmbdDONYEiVhjA1WECyT+wp1+ha
p9mkLP/G6557ncptpiQT4a6tgY5KWq+ESEqSlUFyBzEFfYebER2SO4FXKsi0w/Nb
zeh4EwYtsJb7XszVq6wACzOIgPKPdE1PQRoB7VevX8Uzvd9W3BtiSy10MJ7AsbG3
5Ck1gNWft1/9SOdsZxBxaZuzDHY/PnELSlXMVxu9Zn8jC1gd27ew8ma/raZxJWQn
7/jNzFt6LIO5ds7O+QJJEYSL9J8xCYV3AnekrHlLGiHHs/hjGLKWzENuSjV22kAj
pUogRwZqL92eZo7q/qecoLRsDAl1gHt6SH/98auIBdeUmieKQoruDdaUzp1h4M7L
tGVCynHVHLiOk9qlJv16clsFr+q6KgnrBkXQRTgvyAqkwMdMlmgWMEYbzBv3Od4W
PxGr26et7KbfUPwa0AOSg6IR2HyD3v2lcapMadcxgt/CgUIsmMKpn6onxi5EKHZV
WS4+cvNUtTsn6HfdopDvs6pqqlRPgk7jRDhhOl55LhMstSbtyLjpWIpbePlz9xVZ
fhpExMJ03tjmfi5XWI7uM4mI9uySDanNFwZeAEpHdoengI6mKfXyWrfR2YQfEV5C
NLGWolDdNEa242HGScYs7BgpzuSJFbQQQEMp50sfuIrMBt3e9XLB/6PTbqwHENEW
+RmV45MZemGkdpfK4tGk50gVP2t00UXev1QV7QjtmQogr6vA2I/hlzSWJ15RYh/o
MQ4Dofb+bczYMb2AQgWuLYVvMxLjELLAJScMgeLJZg4Z3NpuJ5shvHtquv4nCnIw
nZD+UWg88senV8e8yHUxPC74kxMMC8EUSdVFLdcVdXAc7iz4MvvfHzdlGbEnhi9/
iTcbAr/+57Z5krUyYfrGee1Uwi3uKb/FVgo8qZhHf1QG6/cIc8LGIobIH2X6JPMY
akt0oXBPvwURk1E8RiiBVAVznjTIg8lP41lceAmKol5M9u9Dyif5fXO6goufnTbQ
O17PXA39tfaDyXG8iQ9aulLeDoguTXSboVojudDAKpaoA/0pVPHX8z2diPkEd9Mg
OWIqNofOS5YybiY3gPFXXawtuUnmLLphrRCHioeEEhQv3AW+pKO/jaJ0U4qSEGQc
Ju4Urw9icdVCv5te8TTQAEInKlQ6oEpiG1VoEtOwH3VF32TjoTVMHoWIEJTeQyds
HMQ0XpouREQI7eMB3VQFa84wC6jbM1DtMFgiK03fYGNrPIAS1n+SsbSlQhyy3YK6
Ezhjl9JxYkDmuVJuCQSNpSnK6z39NSSipGIcq9qduI+NaANZDKkl6ef7ZVpLiP7S
fmWQ0Be6Yb4Z7pplAUAk3W4A67nNCWUbwrFR6FOGUIpcMfri05S+fg3c6T5P4g24
P3ip8OTf1iSgCMnip07bgDN3zWGAimZ1SGh6s1MJokoTrdaCHqsJ4Jobp0ZG+V6M
2VO4FbB/VJM2ilm//e9bZELxPdnKu/f5wKBXHesFmWCRh/sBA1KYZkzY7H3HHeDA
34bFwynJJ/tZ166IKEqhZIqZ1+Lr9F4n7pVsV17sjA1iKoJug1BwOrivL2yt775s
BKqAROx1RPotd977gPpDFAFtuzS58AXqjK7IfhgAmit9Al+lxrfe9ypNCwQ2gMsY
mdUjXwZNf++BR+s6APxDWs0q8Rltu0T8+Xbgappxn+JyuBh5rkx2aa10z4j97lTQ
LX0/QvmrzYOQ8ZdrNkWb4CZDN5OUdL9fO+cd/sLPDTP3gTMQXFcYiNG/NjNPZVLK
UdH+Ey3gGR0n6CzqlQlS6D7+kPAgcZLYV7SD74ijivKD+QkCSFrQsMWbZ5rEL+gy
lQ61toPANZyzBPNt1GemvjotH3e9qC923KjIzUD5kNwHLlZWJy8NOesCe7b1gH+Z
vKp+zVOSA9X0xojiMKakm5KlmbXjhU/z5l4Qh8woV1rKh9JzxXQazRlbe48crFkB
C6ctOYRShsxXm9rpgynApK/PLMWyNgw3n5XY6CLzr3ePX+QhDSzS1zr9JHJ4N025
hTCf69YyZWwE/Kss7GrTxyiwxpZ58GxkBox7OHXCr/ULab0cGuN2KXhFU4ABvkv0
FJHoZml3DD3tt2hHpJdgldbeAgcr49pJFr7mwrPAKD6LubyoEVESgjjFysxS2AOV
3SSE5UE3PIU1rg4HMUE+4ADeoCr5VMsBOgp9Rbg5LH/2VzPcBYogApVOifIFhliA
I1tz//aRW2FgeO91yABWkYBFMkzoMwlRXcg6SaXAhpvd+X8laYntfHOWwPn8JwQh
xIV1QE6L0Skdr3vmiKzD+ftP0zJoDgIjWoIWYZemmxM4DeiOqzx7otziIDdQ0EIS
ABfFnx8C2Da+OVODY14A2cUXd7LwwZODSEuZ/hW/6XAcnW5lT4d8iHgSc2ivD78r
CnjKxGCfCbzxhu0/syGuJ607mWiZClbMbHKs2EbQCMaOm0ZLyFlkOgmBivlzQ466
bDS+QbUebvjoU5Z1w4epYLz2bZpaUdih5Riu6GaXfccyEO9/ye5iAxGz33HWm+za
UAOl6Q8wZ3sVfjuxdV3Iapv5oSCcFyT9w+h5NDSawHf03KrjRo2HAs50rS71i/wb
RXtR2nsDn/0oVyNO6Dvr+fa26RtvCfdN1qAGIEdrt+aHAivrFkOl3l7XoqqpOkB9
2wVittT5NfFstSc6Tyi9AEzUlTvSjx6LwKFmxHH0gCIBWLrr9j5kYPY21mumV95m
Ma/DPdTOTp7vnTh+jhh9KOpocxXPLy+7GdWdtk2joyM8YZZS4g/oceRpJWqDP1q9
vw949aafcTnmhX8YvWvg1tDPgatSqmGqUYlqjuP20WDwUM5HRxklotvsSFZrfRYC
5MKJ6zDfytvLsrgA3hfvTa2Sr78+fpX1Yd9U8TxEV8jA6UiukM+xlYSoXqpzZeUj
vxms1om8RoSzxoDAlabbX89tMGCd0866J4GWEgukD3u8Dyp1qgeqHenraxJwbtni
KRpYfvj1IIHu2DzCQa9kG6wi1gOwjsw3HJOVH8ygO4MDRE+zZYj9j3FKtK168x/g
wJgzSMISqdInrQlPDunFeMOP930tsLOoghA1ctYG+GibRH/ECraqhJSZpbqWZdjM
ce85+iFaEm5BO3JVz8XCCRPb33SoM0h2plWJ7sVpC5HxvUsyjL+yKDE8KqFoiTiz
PWfW1tKZ1m0cEzrIqhDu+/2uH9+gMJ55WPoy784jd9fHQ53hk/msCsxa4XJRwQu4
S/17eB7k9ZfI7IqFDXPn22lTswNuRyljwTyZyK3qkiKE2I7WgxmUvK1t5y0/PUU6
npKvQv48RphE+GsZ1xvxJe0++pBoi1riL81DULXWjyV48ifxBYYwp+02schkweTU
FWbGSwamVLRD5kHoPceQnOXLtaNHfjuu5zh/XOtpb/boVwV3Lic87JxkUNMLjrwy
yeGWhBs2vT4RgVfXveprqpXCOG5lB08iNUJhIjSJJzEnsno1HBVl2IrbScZjYgoo
9SIWU5q9+E7kdyxubeHXoCINn9IMYLgpucyhp3vyZRp6T2fcQFHGfO5h5GdTINaX
0qwo6eD/ydw8egDx/FNSQ7bDp4NDP3zC0BBjIdN8dg10zMgsSXw31SSNlrF0eSY6
0hlShxqodNBHq7ysBvoDW4/BuKqgYZhbGece4ldB/FN3nyJGnc0urMXOG4Vv9xoq
xmWxJUnhTSgDGXUuYalv8eo5VlkvJ1vdkbuIB+dBN24tq85xhN4hevnIQ3Q6QRpc
dzS5YwafdPNyUI6CptSUaMCjXeDk7vFl84EfKKZsOflIIiZdlnH/jhS0Pe44Xx77
Gcu6vK7oVPmZT41U046HLbzEInKzhqA9fshMsttbAfrkCvpcgGmLMO0yvSj7O+i2
XmBN19JaMFB7URy9BxM+TTeM4d0MCndrFi7lq/G2VB090oyAxqlPUjm9cnqkYO0X
rj+naJ5hj78qr/su/lJ0rJ1XJ8wznxDFz4kn/NeeI1nwEjeEEABbtawH4+G0joNJ
RqwO57jNUsPaXcbVHR9D5YvB9ClTR9L5d2M3dI7DdhTASL2eBvInfP7B1s8bP374
BSJ9HhTf0JBaByZRqlkh2UgL1q8GWXlqKrWfuytylma2Alj33Rc54A+XffUlLx0K
OTlDrXFzTGBMi+Tzja4u7QbfxFqa+Uw1wgjpo7eqV3RwfcZA1vvY9LoWt9zjmqEl
GNnXxfRh0c0QcB+iZp0Rwyx0FRVZCLfuZb5XyQd/ihNnUiAZwlBszamvJ/Td36Xg
iEjLxyudbW3df/PAwtq2TzD9/xV+sIsEZMiJj4AM1xQsGCrcdvPPkqXegXgX63t+
x7PTT7NeecOPCCcSGG/8XW9TJWMh0U/qUWeFF9FwlIwAn7kSdACVjMQI6AlSKlzq
BUtfsHYxEGN8br7wwuVmv+i4NxDufrnZ3aeAL5x7K7weFQRIVCm/cpWZgb3UpvNW
IqvaKqaa/K4ZhkVCR+xT5/CGBlDmXODL31P8uvwQvTdx7dh1hnkH9XLqpqQyuWzW
Ec9vT4ofwAgNb09736yBhbWVcXBQXKrvVlXVJKR2G/cCScVJa9bf/CMsC0nPEjYn
l6LvLnynI+EqNu75HltibTXbzD7nkQw7c0dZt8iJoVicqUoEVBj+SGedErpRr0EZ
vg+izugn7cngXcy1UAorEc/49/FohmWM+kgY5d7RrbyQb82Et87SnPeNcP4aG+aa
akBnto3efg5Pa0mmHS4hqzlVqtFe8MFDlD57ccaE83/bc12fHZuulcbwOYdZeilT
tWua5yOU5Wtm+uXuelGzsecuchemaRjEHyBmMTlMaDMItPxcYJYRcBcbQWOIR5Hk
rxnAkYJwVbIz5Xw+SfmJFhvQCQzTOzFxB/cUzNziVVWoc2Cb3xMNPc6pNTk55BSa
5TcVSJmxRMVYjmDPblpQJRs/3UT6BxGUt9zX5AnmI0SHatupqA40nVtwqLoxGRxv
PENHxuAVwEJon+fcaDWZQ9KLsnrF4UHHQ5IPkst+1uYi8RzeQ0mxk+44UPeWQMCU
Rdl7DlDVYVuK1UDk0ihT6o5lhMpypCGK5k0vlBvJDEpQ8kQUKyJ9dnInPYrsBuTX
DOc8XBrgtq6sNVrBHkrBzviAHhaXhlvTQ4RClRFXbVHbFc4H9Vs7WDE9bTDA+I5I
q/IYOtv8ILJBH5lotuUsUGlbMT83PBPkvaccaC5P/osDttBw+LSmQPf8J5X9yRcL
/ufGZ2SpDZ8VFJ1drkj1qmjyWC0+heHljHlc3sGn0Dw1DQr/QaLfDUZ4Wxbmx17t
xTMgj/hXjmIe/71S7YUeznVAWSGv/YWtpj2z0aAtMGQ5fvev3XpqZfmgf7w7e5Cf
saNStOBNSgpB9V6OD6OW5+PqT5TUSy0j0qY7ZlMgY3oPG5h0mSQ9krh6o/NL81Ll
gpV7hVw+XmE4hpcm06r5IjanoUmsG92OKxxrdX6YqwCWL+ccHTI6JuFMMzMHhAMP
OEr4buXljXCAdxDs49HDl7OZk9uDvlPA/MNimHsQ9+TsY0ix0pSB/o0MgG0pwauZ
mt9hhG99itBui7vvmU20B3tCcCKI3JmQPnZyW07NHi7INEH6n+o/7347DQO1Delq
pRXS8gAiUtfFMzQzek/qam3SMgdSnBP/KssYt+0BVhlzNpPzOp/AsGSX5cr53vPk
3j+xWcS8aMvlLQPtHayBsY23CVArR9LJZ4ZMunzTCy6Idg0c0N32+GY+S9MC/ihc
F6N797ZFKUwc69nZitnZxYKzhK6Z01AiR4Nvv4GlAi35csfO5MLQGOncrRsWtv/P
+XDFIoav3Std95q0nyZ3Qwx9Qt4L4Fi5EHaBD7LiR0T/Uu8tx+nuBPLGux+pna1e
Z59/ADgsL2xBs0E7u2QNe+hry+f1elB7c8YcX2/nKt2nwJaRS8E/yEL/khb+14C7
FjCjgIEjrBz91zyWl3O8B0+ajMNHmsySYcJULEZIN1HxtKdA2ALZKwfxpLOXOpFL
m74m1SQW/KfsP4MovHMf0revCUlM5GR8NP7zY1LErx9/SaqV22TEUXpSAqHsM/hB
SleNuLpojb17LEeN2vTYCMtN/lPNaNpysLaVThB1ViNJcfRDV2KtSrk/0B3WCWe3
UZ8mU9KugjA+fnoV7vHYO7w8HYu+oSfCY5UZtQTgQ0fPN28BEFR4rbMELOIErWsl
GOYY/YzkkWG4erCenKkBo+Yp3c9954+uho1oJv6BYWWfSi5fmpfTJV1IeIPvzvx3
b2kJc61ZyG89wRLM0hGiWrGYsjdtP1bhku8NGY67Pt6s9T1IHptB3excTM2zxPj7
+oXb/3rUfUIELks0QIHVIEtB5ZOgWrYiVjU5D6G/q3kXLWzY4w/00ac/b7aPlL8c
EZiET4NJKoohxoo1wY8Wrf2y0uX8bESnybuww3STlKF+q+QC5rq9QRATHEnVVFHe
sm8xtG79hTSy3CtmmflszfavrOv+iELWZOw8dua5paKPhDI1oC6HxVN8dhfURd0C
P1QrqOBwaz9TvHyTedeq7BSyAEwO/sLxnhzJuhkciZxjpOGbbqIII74OYIRsexup
Ivl1P2pqk0jB5w4GWm86Qa3UDU6RlQ16xW+XAQzRkyFFCkK4E0ZffPj8DYe0hdEr
LizQDnt3EDUtF1s7pHkYuYEconQ+kKnAxAF/TvYiGZgu3asTrxI/uMynuqZHoRgQ
FRpdwlf3YMHm15MHk3sA5eEWAMlfLJSJF7rTW7LFfHNCZYqc18xh58EAZIvSIqwc
cNprspUzmNlRrINXUknHxGXHlxDsC7qAwjJFce7Le69EsXIhmdwgF9s9c6yrepj1
VN/vDjOLPUBblAANJnE8pGNo5I1EY1Te96qrCYIq5a1GNH5JZMn3NB6mK+2LhsmM
6qyu6uW8vLvVMSCEuDEa8mo+R7CuVCjJ24wbTwC+NxYrTXeHkmSXdIHK5zu53gxu
4VSvjCylVvDhEVKfkxHNFAYk6J1zWFV+zcjLKD3DAVfSAJUvm/X9p/Lys/ajtlbe
BCwdpBLOcK3UcLrJc0aXqBuo07v1vOhL54hOPJd/VqVc/iWs9tYIQT09DeXpBX+y
okA6tb7AgRvSSqUIIEzaKu3L6rINbK31pP4lXLgm21FPzVywmk6s+GVLhndHNkJK
XteuT9872zY0rQp8YuUOIUsLDGRF/dkb74CWtIXYd/GdCNF4+vlRqF8H+kNLfnHS
tch3UxJh8kOCDTacyJCnlkvq5FibqtIZK9iOf0AJmPUJsXzfaiJ+6fCwUE+6C64q
//R3Dz2AVFMVYDzf3P9uzcXKYxMMxlADVh009RQ61+L6VZ4491eM0es7FE+K0nM+
wdSLR6QOE0b6QXhydh9BxE0CAxDg+cyHsNB7hkKjGvfiq4ClVTfHKYBoiO1bDcLl
n0SANckRc0CEBDBz0jWDMX6LwlITrRnUNYsRiWlHc/eikzCj072nAvKm4+vkNGM3
NaqFF+7Arte3nbyKSdHkgynYm+aRVnNwGeDNkWXz33vgOWDDXBU+cP4MX5oLYN8a
3V+S5n5Q+9Q6zCWzjo4lG+fTc0Z99XZnKo5jF/Mb7hbO3CHqxRLIlu7yNWe9oE2q
5cChShSe3r5xFDDUckPPWZtFVzbCyhn3zvwoVo/dxcJdAQt2lHppfQ3vVBIJB4k8
x5HNv9hfJLD/jo/9+Is0T2WKynsTGtw1yS3TH85PkEDHOzz30Qfvj+lJpW+fjhPK
R7gSKA+F4J04+UwR5WtVd3HaQ8IVwO07v296P7JO2Up13G3l60ubMjrmOpKZNveF
N+eCse6vP+0EBsV8hATvYv13TWZiaKEGMrYAisrDH7xTEhE9lCtbTWMg86R25d4N
5wL8q/vRYaCUCw6ehd8rEqxYITvyzfnF/18m9urLPADqDrRJoe2wx9sI5cCITkh3
oVLdHdATsli1DJpz5ty5LG1KyenUl6zCZyl7/okmTbWc5ilKyxag/fqjv7i02yGO
F9fmN8d0n56yrmonvLl7QwwutwwtFnmMo95nvurpdAOEL77Km7sIvaRW+CVtg4xw
nOYsYN++ZEAgavhrppbz5SFt5ppsrF1bDA5I0t78kdl5u/0eKLm2R4zWvUVagENO
ZY5wjerINKE7xwo8+jzY/aLfI4V997ZQVS5zDa3Kx3d16Zcc9oegGuZwAJZqylx5
p3zBSIXY90GgoKcQzSKlxyEkmYgnVLvTk/xlyvIBtizN1flZq+n+92bNRQfsSAbY
HrhzOh0v3N0QkH7EEpiIvI1/sErd1WhHKj/WilaoVXwV5U4U5p3GZuucI570V0pg
Stmiamtajhh/2ldkXtAleyNS8BZ2QgmH0q73/U8rqv60PZ+jpPyIfDBDcVLDnRWb
T/B0kzLAMunnvh4LAEO6SvHjxb3VbsfZYu7mo/FE86fbhfV+F/RV+ZhjXGLMjKzA
4yu/T9IubTzBdRxoBtHIILJnwMooS9NagoHiz08uwJ+aAnHaAqS2qsFOPvewojIL
ic9FSAcUTFpyxLp2hJ+oanE6HP2zvihewv7mgLFTi4INBkwOR/rGYBtu5LusYV12
KGMpBu9QAcnIxUyLmxCt9vOZ7d3mL4ppyS1w+dxgm9wSntElj/et0ubqnKIQbvuy
6rdYMP9n6LyZa0SxrwLv+zIupUv898TCaBxXolmzytjZ0b5+mN9miv+UZpEaaEb6
pjagXMOZH4lGLBNLClQ2kuO73sMwq4DW5/cq7/T64SPJzkYEeWzm6wMvX8pTf2UA
Rn6vN/JEvsZPulgbK7qcgNS6Fuz3Z6oOwnZhN+ToRGxBDvoE1wsNmSSsOYWcwe8C
HlyaHUrlPLfJOcNEH7RGTdGhqPdJ8jJ4MjeS5LnoaVvBPOIxLRiRaL3H7RBPInTK
xR6UMv/dkZ93Qp6QRL9Bhc5hqKzVc7YtQgawSgEgUCYiuzoYGsGl8ISQDIrjR3gv
HNgx0CrHwiY213xbHc2PzngJ5D8+gNd2f3Ue2KgshbTuJcc8mZU+7eQQMS00RG8q
HhqC/CHdMH1PsFSfgwh+XtLxKBAgZWsgF2zfDxpU2pEyg5g2WQA63yKMV11mbh/S
Siy99RgZNRb0bF5g8bPGOSIta46og0RTWq590zXTQpoKZVc6BlAmYSJkaCaXPLZx
Hp1iedg2R1Lc3EVrpFQXEDnH+TG9EC+iExAoZ73fCvonUZNZOHsuTuCUqtOmXsYS
dyoU8wI6uvzmP+VlTgxKpI7WrLUX8+dM2iB/asq3GAUlpfDvosA0jORDzmJpKvl2
Ts+pcpnLRFa5soz+yUqAZw9zcMg+7gpyrNpQPnn9SFyiWqckaFXZKc2UHRDwrsrG
BzmIsJWmUtYhv7F9z7pjpXzHG2iHudDSXlgtVPHuJdq6l9Qxjz0+DXYy9LxjhCBq
hJRE6Pfm3YT/+MMiHqCNNiKCPxstSeFC8pqaKJ3sGdHg4mNYjWdieAxJpzMpYXUP
T7PECWbLJhaDfIITmzk+gCozAoZCPqyZfdMInrs5Uyv2EATt0T6i0Mv/OKhKzArP
ngMf3CMNagnZLWxQpZb99nJ2AAUg3RVeGdJ/iZ0W4W+6QpJsIvQhdhFZVAUKMsGE
OISQOTsA/4Hz8Jb6SOFZiGjndEJ3quQ3CnmaTCVwAmoehR1lqghPo+XQp2dZirk9
AlFF6CRkhh8iyOwPqeNunxR1gggOxxlGGBrM1eyLRPHtvwElQXUyjIxyonU1oVX9
KP+Vp3CANhjOdBoEPuT5uGYVfy08JVOo5unMwdEyQ2UFrfA4pqHqenEPhJdgwRMT
y+tV8YKJh9BZgOrge232lBMfvOyb+Lql9Lj59FbZ9iCCqV9I7TzQ1JgXm+3P6qCr
KR1iFNcXA30arkdmG1XGbPg05ESNhGnRhhSiqFW217qmsh0Yvx3cf39kUE7tjtT+
cf2z+9hlPl75o1OigWOFAi09z1AgGgCCHkRBwKIZb3vLsl0WOPwzatTpATwNWENp
uqGIaCmidnVEbEMWwHd2OgA6enElPVMSNNRJDi1z6BssL47kQpN1vUfb1UXZ7fPB
1lZNcg734RQCEbjgx5+ODTwClfHyraORT15VvX89dFEwgQaiyvideVKvokhu06Qu
vNwqusDbeY34/8YS2cLg/71Ok/cCUa2ehfOZL5fPcnHtRRrnqjoD5vxdQq0FsGX/
CgaiYsnVxQJ1zl0yamEzDhD7kt7jy9k0ws8JCObMZm5Pqv7F/7BcqPqP4UXzMK8V
NUQM3Sl5JtMOOakj32I+4XeP6+e9y2VdMW1uV7aGeEv5DVIodcqaOYD1ncivitkp
+Quv/+NOYUOW7/si9ws2BObP69D+fCQRcnSiGvW9PsUO05sXqOXP6Yhwu1VeXk1L
u/XMdvCJOyKiBaENKuY8jXi+dSBIuNgujxDYWUKegeJM17bnyBrW1/UywH7W+dCD
S8R0sPLvTy56m674MNK3bVqDGJ8C8iCblwq3Nz6HwAuN1Jq+fHT/XBxcODP9rtJo
B/9ejKZR3hX+hCpiEoGExP7NOFrQOEk73gvJbJaL+C6eExflhAOh5OUA7GGauxBT
/ld4v1IuBDzG36wgFLxh4+x3zCwKTa5bme+oqQRVZzd5p/hooeWnOcIxznqo8sVY
RXJrt2UCuS40TqA9ysSVdk/NXJPoc/82VYgNO1lcGFjNxw2YpVvO9XECqlTsNulI
NmPIuOK+ljakuuqkfa7zJZ2btbEN4+MeU7IcZ3Dvlc0YroZ1Xxih0BKgBDj4Rs1o
jAdT5t89iSUwzi8JdgGlwfv/s2YyQ3ItiOO6xX0aWW/kiQaPiZ6CA0lxOMYVq3qD
7OUDi3xTLe2KBu2R25kWEKYmRRZdxkC/3of6YPP/iMkQDzEa0yjvbAd3rBP/NXeB
gVpNGfywE6dAaCPJbD5tRW9lL8jkVdRoZumOtWSTpZwSl+ZzSl6CxqTiZ1hgcFRq
ULQOBsWDNFJu+CRlrm1KiubmPj7iMVpGJNHxxbBzbOjOr6mYWBFCRSmk53WbZQ01
5F+75VNKRvQ6P84BXoN953czk6YB7XIzP3Z8yl4BboVJaIj/bwm+lfLiupv0bb6U
0Nj2wtwj+yYqdX78Kq1p8Ie3DnMTQoqgDHI55fv7zYHivEMBDSmZN6/DEjUETYqO
EkUTS6KnwbfFDht2997G2SjiHpVVrJnlv70nU+agO3+J4sD/ed16syzQj1sN19GG
QSyVaGfgbb6xmYc0MBXKj1Twhdw1x/QmHL+XcznvFBHFH3xp1eGDZQf+mKCmE1r1
ioncvK9zeukLXzKWPRULouiE5SpOD76zI6iX8vI/fVNHv1/gsSAsNoldAUyR0w84
DKPR9gE+Fn6KFyWruHJafLTZtZVP+JwIET+ZWrTihMo+ldVC0EyjFCQnB6/fJXV9
3Pq2KwfSLaNT+fZtkfK7SYh8rN2sX1pmb9umTpKb9UlyJpAZ/aLWfWHbhe7haU7z
aMFJJrW8JmLnheUo//PjLU9eUCh492FZMujN3KnyvBOXLCn30exRWPRLzOSygKM0
HWlVQogrBU2N/nv4RIcZ4s5rMlBEzoT+yK1Rfr34AifQ+Kx48ijq78U/lLsBekOO
+5wb2b+jKi3iar/faZTBfKz4bnivsDCf8PmJJJ5DmccvgRbKWL/R0htVJAyz0zbT
LB9rw9qX64KiH9e/KJJYlONE//Lw+I3aIWGpqFyRL27opV+lPsEtj3LwFkEaIVe6
f546ot+GIaDxBe5D2adqKKeQbkncuYcjr7tkQfBorBKeifY8jfkZu3oW5F8ubYgG
dbbQQ2aNXzCT+bvvcy6eFOfWW62k2RIh1Oi0EjyWnFdo/s0UC91+FBG8Zf0MHXR8
bpaVeDgoyiAXhmRqiDArHN+DICp6GhHWXOqqJqnMliPxyL4cV2TWklQRsDXc9zfe
udmgcKDuyTjZvBEAi0HgvUbiugjCQMv11LKyVVlzefMHrX9JLH1RKmI7wCghDtai
Js4y0nnJSpdFToArQ4Oqc/heoafzd/8B+21Wrf5vN795dDO4o95PhyosmaqxL41w
UkAzXdAwox5cs+txoiHLy63quhuA80g9QdYprbTCyehlR1dQ+8JKk5dRgp7chDqD
kF/9tocb+VyKvbdCRHbHXx0MAY4wC91TG+Or7fOSpaHRqZKOhD21MZcnPP5G9Vx6
AzBNkojnTacyRjLJFRRg5CbSgDXbjMOzHygEM8JErSZLjZ4dIWGNZdnBPrQ+76aW
/cwtkWECVLaNS+Wcr0MJ4VLKG+KHI0qrfnC4vIYUBjT58hMmvqn/ff5yS/Nt9mFj
cZvla/gGB+ZCfl5AmcHiTRDMbcCpAbqa/cnn+ezUUXjAsl/Q01E4FyhYEqo5nK3s
XHZ/gH4BaW/m4pZ1MPfWxxcGq9Orp64bFwB+fg+VlQk0U4VJmDTEDaR3qehF7hUK
TdCjUaciv3r+UwF7JPHFZijiTJxoRqcZtWBKYIWdZcvdxFL5qjnEMkHRxZ1AJ4As
m60MprqjPlusRw6AGJYZJJdRb7bAsPDkUvAMgTb5n0ZxP+L2x4mzQp2htOUuGLnM
X9OItEodANOJvsSVKAe+C1mu+p7fFx343ibSX9IpNoo8U9ULkPAMianMb7WdQPix
wq5AFzoxiEGSvXIM3z1JL/bJ/vO2pZSexfaqPY5D8Yxjz3E9Ae+U+zUlBWwv3KsR
EUR0LbzeHokYcKL/sRouT3Ng3zJyJbVl/VujnT5r+sw/+MXqrucqDzQqfaONIU53
6WB27rNvNQiWRDku7LB+YDZcKgHMqu2cgi+3rACbp+j5+pCRuG/QZRGkTJKC53dN
rehjJpwisrTigmvFxIhE+RtRWdEbNTid49nKZcg5q5LcKatuecZjeLOIMuaWjdla
SqzAVPLH7N8rP05a8suJu4kHjGf8CU65oNn1YYx1Tat48uYPW8ZhMXHJBo8/yDAE
OEMrwMdK2ue/V8QLp/TSBScYZQABGXtGRs60kp00oHxgt51PAMAZp5l3fbMPXawe
Plfnb/n5uthw0aXJel053znDfmQnNtm5Qz44O9A6SgwflQr4bHa+jcMvJ9PG9Tca
7Kqqe8bAHEsO8FOgiuBRd9Ovoqili5w3viKLL9buoyb/9jlCnbYYPYrFHXCIGqw+
hCgBAVuSoLiPFLF+9V4i8Amuj8nHZ9qBmjb/UaIL/I/kSaWL/lBTGDrMUxnCGJEh
euaL/BmcTYSMGUUuK1DHJqXUd6Wsze5SAUpXDwHT8P5EuUvdnHO4RLyw7Y4+K+9F
1vco9Ld4dNiu9wOMKmx1T6gKzha0S3EjTEwQ94y8ZvL424dXsrW5jA+uqPlDLdZZ
RuvwpQUbziTvp3Po0ZtAFf1KFL6yutD1BjjksllT3I84z+tQXn8zabyxDQfrhiMd
ZVKNW2CSP6Hmz67Oh7EbEFOvoPMirddqYWH+ZZA/7On3vbqKaOFJ1x6WYRldy1x6
2lJsBWvt7ItlRpzzU3/PFWvY5THyyuBfLLl87VnNwBTUr02t4rJTVorMPkpkORtu
xIJvDLziqiZxOljDd0ZIopd44c2Y8PESc7D2RH6+nIK8w3otHaRBlG8h5XyRxIMd
GT6EPnHX9yhBI1APORBbv6H4VZ8MJ8hMGprToQUSK2rqBKakSmhHk6hSFoZjQw+g
XKDCzdibIaCqzJpv93tKb+u6FnrhNP0hQqZ5oZvVoyWnD02lXFmcVQfSlESCruLB
AP8xdD+YZZMN4OAPXE99INVo45Z8cBbIosAQdpsTvZKHdGZBHH06Vy2gFVlYpk3z
JVjbyRPxYL0Xx2T6F9oBeNNyyCuUzjF4bO1D4glDQ7egx2oUT/h+jFoe78xu9Wx7
E6nrHuCoaE+FKBBYy9Zccv6PJcU+KVd5m0ybiX0FyeJ5noeMzVoUhfx/YgudhJDV
awjajX3amhkdDOiQt/YxpZn0PF8sajrHMbvYpDTxxDcnuD7lUcFh1GCjEA6BC2Nc
cJAO4X2g9RaSA+KbrMWxYria3lnkQgzpDIaNy/r3vWNF8RxgyYoRLhb0aZMigz12
UB5fmief9vVe1bussM0HwUcR0ekeKOQ8VvXtADcQbzN0F8V5/3OWhZ2P9ribjfHR
6z6MPAP47gPpZKDa+zgaVpOQbaCi6UwMlUOXMSvqTKYlTagO+poFRml9rqqVnnab
m0UPKDZv07c3vqudTKi64C1GPsYZYx1tK3qWgeEuRD8SasmlDZt6ef0m7xedzdv4
LrshT56yTXQCkWtNVo3e3Hqocq4Mei7MwI50k4b+p29RDuPkqHNAirnxFtiMQo3w
f/yt/CBIXHxEAma/hSj1txKh3fw0DYQkQOE3DjxpR5WH+0xDIaF027743YbHvmmE
RQD/M+Wf+bCloJZSH/Nol4oIaZ2HMvUDa7dL5iPUOD2Ssok5y2rYoaUZZ2y2JfiA
80wDN1mdvxksolihv1sKV3mGj4yy1uXtPMOhXnrXurDpYW0xK0i716WIAUk6cypu
xvmtLLyqH/Kh4T9oxvn586AKKNwj3HXdI9482iArRyVJo99/75znYLnl2FfFVdOR
mOQw91FXeFqL85lAFzZeO8MTUmSjXI1yAAlHGk7LN+9HHOolfoSkCByXBhuve+PV
Bau7EtDgluGH+jFjN/oo/se9j3uCpw+5P2LOhdFdu5j0Xku+gvZjDbG1Q88uU5zx
1mAhn2MRP8OdLIhuxb61TIEfmsVYRm28prcrilouSeCjksRgGezgjF8T7yqHuGL0
e10z6dH1yU0vuqmE/2bZuTz9hE5vPMXSu9PqpLw4tkOH3QjKtST/WoIPShYsVFLC
n/zakAXDLJ3PFwFQY0QkovuFNM9r2c2lMlPHHQrvSXPHF5F/uQ0Xv44rVsbKMYuQ
lxSYKLlUuMFx3fhh8wCcPoqdKN8RhroHG4wIOlayQF/bnkpOtVbMidlupkU3UGGP
eWvZbTLtxpXCcwDd+TDvLEz9s6pDp2arnFv2H3jc7ZBFDVTJKQOcQwmHimWYnsVe
JN9SZdVADDt5kFtJI2WmjP9vmQ8j+SHSKmutduh2zMJYNdsTVgU7Tyj0IIenRZIQ
Ny8QOqzm+IciB7E4ox4nrgQAvArbxh+JPPkkf3GOjkf0KZYnXmhVyvFZA7q+kb8d
nZqsyvnedKeqrlrHEgwF0DSj3DxN9a9b1MWzXhzNfG0CVyU+6CUVBuP2GXnnvh7Y
qxRF5E2hsP5XmhvGCvYudPdNpkZibb9uCIZBBCItPrQXPvXm4SS3I/3CFz4TkSG6
839JGvxP5CWufACO1C4Sge6n16kXg1564NGf+YMfka4xC6rAVc6+50ZGljLNJ9uV
UstKtZEf3h/1kMteKOQUebQzWH1DP+0nyGow3ORETD32ZUsxEEUld2eUNHg9Qz3Y
tY+fbaqfJluUr8znjDlEIZ3Os9MseiHJ74ReAJ3fZnpW7xtLRrOEeza3f3sVKe8J
iY5Z81jKiGuY8JoFdZS93If0LDgHwDK3NBZ2I+mHlNaiX9FPUfFLCSP7dBwMQ1lA
j/D0Vw/xsnFf63HULZAIR/HVPEtIVNAv/MZ+deUQHpwzMU519ZohfP4a+Tbwtm/W
LnFQ/Vqd2U5BPkXmI5y8g/ECxqw21szKiz+NyUuFunhEHUZ0Hq4Ay9Bt3+8D2e8v
RcqglJss0z5lgS2B/VgITPJ+GhwBmPLOzV3FcIr0lFXsh9tgTu15jXp5oYRlKex7
6dgsfYdfqV8wuZeoHLJRHgUE6RlCkmDzeTgDIRo6dkpHh/fy1p6XXGIUnZg7u20r
Ens3q0RtBm4HCBQZuKFZ9B9IN4EnjWJE6tGHcGz7pdXdBG6IhF80Fu3t3A3pIaSA
bIJHNFEJyklOp6KjxK96l44/da1Zv62/+hjs1ZOWnxhOYQ+NlMoYllzTZDexp1Od
yVzRMXKAxtGtkctTsMYBF0TGXxxAEmoqkuQ1vCaCLb2SiE0W7vdUtw/uYzR94TcW
vlJCyLULtFs/Je5QJwU1v6GKoXqCm4n8jrA23oxZXHThYpQ7kjmDjnAY7dfhGLit
cjcmshj7COztLS7+LI5Br+vBmYx60C6E1o94uh05sLkF1pLZk0I3myR9PsjneZIG
W6QfSidypHLYGMIW4DStgvXnyZI1LttS7VOXzpMZQpOybncUJ8sqGCGEXj4VDwyl
Mt/9qt0yWzaKf7wYkI3d58Hh3e9hgpvQmhukIJuMgnl+Z5o8hXgRlOTHT+UEZibQ
Sd0n33zDwy8G57S+ot8+ncj83/VlqaC7t55kTZRCLocSDtte9cBWNAQNxhWQo52I
X8/ZYAXYXsNlmOd7RKirhMZ/w2jhvEJsU+LrBJHtK4CmSbZ/NhaEN3NlpV47wKl4
Vtp8hfrbLfxzon9iopBMYSEvi/vka9D1Rm5OIR+kHmTi7UqBUThO3TczekjLNw0b
ooVOioR9VyZxOSj9XdAfuBHT7UB+AblfAA+Y7b5vMeNQo561pNyloW1eFZ6qJ0Cf
u81P2ll3pQxtfleEGKz4Sh0xxx6t+H7YM9pVnKlfIpUphRuAo9hElONHF1wMb7gL
KkSTjt1gjKfWBtZnzeoNVoN+bvrTVgRTTnNrEW3BqQHnWueqKxz4KRGNconXWKGI
pJmwIy3RsWYHyjEuPNvaPExFoy2/gLWUqgeU0tdXcrtLMfUiTQxYxCxaHHYmDmhJ
QKJ3vzZqsw4/7sdNrxAY3f3MVBz/hAQhL7iQPgcTIgBGr4ICIFipMvEejgR7+QQa
Us84cdIqpjkU+aFCy40oHX2gXbAulB7GDcQf2uoIdW8pmq85HBU80PonE2Kd9bxb
bo57jl0ZaOR3iaklN09Df72pY2HHJapZsqSDQDXy0377HQ0xXCI7iBEsnMTgGPJN
AoS8t9eoT8PuEGSa9CO7ghaRQZku/zglKAp6YlC20dYmueCoUdk+XbY6+veIujUh
5jGiaBLSAV+u0QGqAat4jKICIc4ecU9/KDMQpeITQKQiZ7+Ch7bqIULirHSQo3za
BOOtS+9Rm+OHaj9wSNPWm5uhJnQcj4ehznCU5Y4wTMbnvMThU7XBbtUcNcwOPYFl
ZLijStrrYrV2zzB3u/IqrkK8SvDN2DY0NXMqK5f73zfHz11/JfbKKgjZtmERtz0u
CcSg2tuEXYKWhAyXMG4UuPZDvOxEPbqRsnyOLHUIvxpQRUurW9xbuOWTWpmUtDoX
Tnrmq8FAowR8oQlVeiYTCTJhXjIxpZ++v8XQJNHI3xh+r5zyLtvYESxCeYcF9LmV
bo2UpDNDfNq6J95OtRIaxKROeAJcqs+S0/nTzQOtdgx3FKHOn94M0J66rvso4PAI
bEmnSCMho8O/NORr+pm21/4GrkOyX7pwKOzRqwOzt5xFDgiQI1LklLh7kw5PpSLv
90ohDRP/HJBsNpV6wQZHtqlMzjiCmoJtwkalxM/f0UsZXJ0PkmyOaOt2wV+Jpain
zoRryERJvZsCSjmn/hjnpttAx+99zzI3JmDpomzXYbDN2GsLvMxpkO1IiTiXXXqN
8BZ/U41WRyEXT3ipxK3CyUj9LfiFC7igl4QzSuzny/iUQDx5KpSeUKaoOya89dgk
AtKWfD7bMkIkT1NPiQGwPtY7BjdPVZbLva30m9SWDfRsKwmNlV13K4nU0XCwRM9m
wQsJPbIOUJ82rkC159NVyjvWDbEEvolOFr+hyHsSdFLP2Kjo/THeDeAPFNQdKsgx
HYMBRk044fIZAJ2PmS0IaXuWB+C+DwQDtQzfxPfKhLKbsEU4lQ0DhEB0IAaG2V2s
Oz6ruFai0HoxwjlpCjkpGePpVmQDzNHA+4zeiN8UO1pldoWiwn4RfaK6bJ6bXwm6
YfavcdvxUMP/NXgT4fHFm+/AYiPeH93Ym5EqBsIZvio0q4YV3oAxJZXUm8qOZ3zv
eah2cwWhmEuJKMuEDoRuZc0l/JPg3Z7LIq1gKS9aEtjQpqWItOYt4Q0aruGWFkXK
qPsO6uRIg8VL5LpU4pu6GWW83HCOw+rNXZagIT9ahHsTosVeAKqe/KlCB9woJPDE
rydzkDdzsL0+PytIpNQOw4j/sBgE8lbgYQQbQLTpV7V7hEt+BINy6+px+LwitbH0
s/ggTRxKxbLaXjSvbVlgMjmFL5aHB4p5/1u7iLH4ySKoXKkv7v8KcuX6Jbc7J4wV
yfkYuHIZwfxPLC1p7oxwcKRJZ73EQ5RgyslGAjwxey3nX90j6t32lqn56bEIxgGS
vk8SzOpm2QMJtn+yVcLV4mRyf8D0sh2k0MhOukjmcdk6yZSGDtueW+a3oXnInL81
JKpAn54ao8DC+ShTRfl0b0KYfx0l57+DCs3Z+V2fC8BHg3YnQ8ik+EWz6QVhuoBr
dLB8KEVdlEvew7fX8/y8ddCikeClqKmlD57choOUViqVuoT+p9dJ1ENtmUJDkFQZ
DSSdTVUm+FROMRXFCiBPaFtdGHlzsYw76lzAu3oPJtApdpSX2bmwdcGv39GoEV5P
C+mKGgJAMdDJHY2bfngAEbTWLj/PQ3k570IkTEYnUrd8o8MdCM9dN149IgarqEhD
zeTPxru4c90Ba+bVf8kDFOxc1ER5kDUkYyN54jiuRkaqPcMVYhQJzYPB+vYkXbXE
hHUrx0Wc0/CBinEUx9sXoZ5GsX5J2l2SGXCA6dphemvRYKfL8gInGDLJSN4FWUSI
h5ep5P6mDpbllQGnBfCMyIReIOSlZ1BShLIsWzhnFS5hRNp5Or6rhwA8doMY3yh+
GGaiV8NalfyGYcInb97q+058qQWb2FBcAYdu+kzCTzWxgiLRdG+6M6g6eF06Jscy
LDAwKOwpl+qt/3HNzmh0vlsvjNVjT5VKF9YSVx6/4HscfofGN2p2tAAi9VfHislH
FXQanGgzfRdVod2iZEoqqk3dydTNU4mwIZawxVwudJBkGBwDCysJoSv3u6gGac/A
1/jwD93lOSrcW0Vxrto/ymAvOXN20lUD2b3squ9QKwARNxRafhcC3VbUI9Gs5nqq
2GJwutfGliWweAS7phniwOwNCDRFqnYJS0ZKxKkDErTjzCmjTH9XSQV9rQ/IS4jX
MsdGhl1gWjfzGn3bnb4zEn6GiOfdf1WdkF6ZDrjZ76Mm+UlzITkW2hdT3RbUpehg
DUVRSO8Sthlw9NiBpoQXO7ADoJhJ8YJ6GeR9gBaMfPZ5jhh8EISq8cUWSBD3SVPP
QuPHpee2LcVuTESjiHSb1dtlxccjOtz7Xiyl9xsGPEsTRQtkLjblURQaH9IddrqP
ubDm4iB5/sKQgz6EomKtG53RyFu9eLdDmkZsI9r8rZeGR2NNIqM6UjuFZwtWVCsZ
fuZ/rgXmbaAhiLFHEiTtXkR+mVh6fku5PVGn2OgEVS1FTacQYW0zIjtOgtRxM5Pl
tWdi19o4rQT0j9Xa/I8lDZ/ghVCUcdlHTvAAUvuqv3I9+BaQKPCbf2FZ7rz0c9in
e3KmqK5ec9EaHw+QSlq9FWUSnJDRz2d8bGNHvV2ikmD/3BM3PK5RzqXSXA4agfpk
LQV/fgBpyJrglLZi4XrnFkSijHWicsmzHPJjk/qLT4wAgRAm1UmZcTfYgqAwcXae
npyf4FNBJmQoRGBXDuYWILHY8xzRMZMJQZglYyx9RoxrFmNXPaRk2IcF4AHz/xBL
ZMNwscFTTCfo6Eq/xlWhwDbyTEGUyXXdTVeo/zpaiLfdUqBirrT8GgLvOwEvGRsw
JsDzRevRu7jozIhlR36T2vSoHGWq067jHoEInVL/8Oiymr8lSaQSC6nUK6zf7Apa
eKlU8C/4ufPtU5RKrqWDdShTjwoLrCh9UMlcxqFqFqBEqpy7OYT7FzBmS0AnQDeE
DS9vipwLamQTfdTqb1JNyIHNBdNo/UWakNm2WQ5YhynvECEP0tymqYOoFCYhAUsN
Otj0f90mvnAwkpWS3gfdCyxcryzsJOxRQHbVmYuB32pFEYaVRyBmrbmd5ryFTESW
e1WR+qs7+9OMVtzq1Al7YZe0VDBxvnFW094MIq5tNFEBI1QPOsTvLQ/3Kl2PdSvY
Nfzm7/1o7x5GG+jb99wOCKpOqQ6YwEuB7RfdUJGxMeEtcGekVOMtio5q2kBH75oZ
B5uaViPKnrOPE4FTXadm/MyFlqoYQaWIG0XNu6/l8mafY+UAb/4YMRFQoSdENEI+
p47ao9u9mf/aDIKDNGEEtaua1Ips5XW/LO9qkAunlhOdRZKK2rrh5QOdYJrRSz5r
A3HGsRNwxSfJepzu+rolhNLbHmb73ht0kI41hhKZOSrf9HUyM/VDf8rh6PKioS6v
EoeNHiSwHFwYSd5oDhQF4C7+woxLr7DiApkuPuTF0CpNh1PdccZMR1v/tChiBBW2
GoHSTXrMklNaxNIurcLBmG8Xw0JH+T6dKFnNcR1FXvDYf63tIWwRmGDPklBf6uMN
whYPPOMVj6bUGi1Nd19boD/G9CECwAqKoVwi0efKFDplFqEfcnjT0K/PVNQQbizW
60Kl8AND+Mi2F3rdCYay5bSgZm780HI19Ok70FvUe34mr1z2dm8v/za0QYM4B1y7
G7y9AhWOf9YK0Yj86bj8r4grdMrSKStRFcZZS+Q0fP1ECSO6WGpIVBGRJkFW6kBz
u7uGn1jrtCysPQBOM2wLbJ/dTKXA9p2agRXUc4+rRbMn+Rvvt4MP/mpECd7CM7mY
Efqxs1AjJB+6GL9RWk2uQmcYYVkrQcY6EntQo/z6b05BUisrD8ByvEP6Tzk/7lfh
lMiw8riE4OYQ/1NuI9C732UmL1rAty7gOYT0LJzNccYQTEou2vVlkVuOajbW2Wtx
x0WDhfY9WfBq2M6NfdjwMhchW9+G6rNTPDV32b5plUTrskaw9dDSQrAsYTNqbg00
EXjkJRuEkwp4q4BGO8qA/EYIHJ36g/pZQa1srOW85Rz04dXiIUdcBzsqn60wEI6Q
VHCofzJL9eYglctTSn88RXDZTbSX2eb3jhidgXaYnVCHG1UXmjQzFk3jrhSGnE0B
DrsIX/bIcEFGAoAy+wUa3dCXRJXLt2I+r9tROYM91V3I7BjvvWas5UQZelWD89yB
XrToWr1fJGeq5+jRvBB3S+jKZJOlHszW3ghv1NLktGmrqU6vaRIilQiLd+iWL3z6
8wLDEc7dcmfW1H7BQzV0YNNpVSsBkqUua3fK6FNIdQ2TSesoCuxow7LJiIvNvIYJ
N9PW/Gxt8mhQ4m3d8VJCvIDFHAOXrearrN1I837hU1hLhbBlBq4nXDy/MPKZBaY0
Z9r56ga9XP2mgHGbYYAap2ShYVUvg5kjyXE/7z560x4aW5esfhmQEWYRLCTW9+gD
kxg+jYVcxteuMurfPaGaE/NBF/O1bbWJs16RWxbcJe6WrZR04+gyQCA1VGZJ2YFo
efD/klI+K3YV2qCB/pV7/FCe+9GA6L/7A0bZidRQsshat3WQzTf1e8t7F95DcYYn
7vfEOl8ojZQuRVaAapSJBf+BfGf6IhER+0ZI9AE6knrr8ZAzUM1xu8uCJWSZPf+G
d3UmEZ7ZE6v0diD5az+mKwyibJ1qspFDpmU3hRRPdzWom3dGBocC4cFHairpXXir
wb9iVWgzhbKKM+OhROjZBBaqEB44gkbJgpxnddHFTicfv1VffLQBSC7WxztykIpj
gLo1hyMcRzpFqE/eOlgcFIYzEBq5NnYMSitMxuYeXsxMcW4RX3r+ZJo2RyLH3gLv
gRufS75jGhWhuYd4gn1WvAt84jn311XiYq5FkAiGa+b2i+NuZ99C8Utd5c+jb27q
bAWKBllnH4uBkrCzOz7/H3BP3YE1f3+sji7CdTR40VeoxDb0pizd8ri9oc881cYt
mm5PqzkcPg4eH7Qdf03gfc5kIUaClMB8mBWjGPnsSwIB21HibpB0mTRwMzOYf3fV
pPAQhCWUasn1CMdd9lse96RpHHGrO3dgRXNZDGihz8wOQFhbwjQU/pcY8n0C0Nr/
9RlbTNnpvqI3dTPKTdCHAoiLKaWX1YTGP+9kkalcDbAbUTqWafDsbonJseb9/8os
kQ47ohdavPYwKGhXA4aU1NSJasPguMybZ0FMYG417nvuGMU1BVJzQZWInwSTU0vk
Raf/SC9OLW8yT7HZk4NyHp7TvmP/C2gHEOqANbuaymPsOGK8xIrC9UQBYlPQRPz2
uXWoAUOvG52ceX1lnhVOpJ22b47v3/hk1K+4aYq5CfUfHW9mIAdq2uOAit7WccQx
SJAeHSKI67WniFQP1wUQROiuO7RfzjyDwJcjQXhclOpE0hlNXpGU8EXcYw+LMroG
X1wHVg1X/f8wqqonuYqVtF5DbnI39yJzC4xNxZtxNgrq+JuTSjBaVqS2s8Hl4E3T
FnRkyCzith45+ICgDbqfIErdTipKEcn1el3l3TH8iqjBPdmZ1iYNwVjqX3taJCv9
EXbDGT6Ua60pLpicdN/VnEsPqporAK6XoQ6V2AwS+ipEykbOTy7ynADth8fhkvGV
9FnLGA56TK2IW3doqH0vwnoi2m60p6zXa+o+JpVmAyKG+u/BoH2GM1mWYm4uucvP
OSwCN63aW0m63BtswOHvHpuRNlUn4ES2hVlF66VcPkMsALDDPN1EcbLCVZZ9if+V
SKzH8tJykd4E6yB8/Qh/Y3X7XfLf+aH7i5MeHi+qtNyEfrTggbEoGFQfguLx57dv
nkolLdHTr00i6QjUMqie7EqMMx7hrJbyc0JsML4aIo0vQ2mDfdOyPZzdCceeK3pA
/16u6cqKK8NnA0HJvnfzO/0V93Kg0DUTRBhdouV0B2XSspLXselEHXgFztQmNARU
kXpvzfjvgx5L2+OvVklOAVts9WyHqUSno+nXjguoKR+Tap4XIFK0m7NVU4TieTMI
5SKsgweGnoxkpELeaeo8TReFVBOT/BgocUvy0bzUbmrQd9btNtPNaghNgOlpeKT1
/AP/cDB58zwB1EmO6sued5YVjMqWP6FNWV+hNahwrMlKH8yRbf/8j5nYQJOoN4Ka
Xt5rozVKhu1FNSzzNJZi8V+1i6q0MfRkS0MnR3zIbWNMEtelekPqPcCY2KbXKog4
z1a8G8GYOWgO+kfYqqPqMEzEu6QyyfCcemfijbygoqWs+Nhn2hk8wMXXhZ9GtxTr
u2Fqesqc1+YxigXbMDOObJdOhZ0XE445UF53OQeFaVkTg8JXBVFBu8xXHuLEXlRF
GzFQgmRkbt6zR+DOq+lC3tFuY5IW+8oT9NzJHfhdPvI/hw6Ou261ngWvjlW1kdBE
9rbvhLSsBZVVPobOplVFkGlfIrOw6Sb2pV81zCYpAuZRFi/Hc2tng65LaM8DJ6if
X7A0+dUf2N21Ei9oYKUTAGLCkFvCFDCAo4TMW7Laly+Eptc3+/hKiUQoNRQHmjXP
n/NleR7T7XEtjqCy/GiJsxvXA+Svr8tFw2W0hHCaUyI9CYvWrhok6GUF8IUWomqt
zEXN/R0d/NeTKP1iX5iqH0R/cRtvq6hGqal69Z7Kj+ocMmpE2KYc2kL2JLPocd0Q
RJj7oonsWFhKV7aR57NyE3gnWaOigoOM6lmm47vzQnbwmcWvTi7n99GXrWezGL1w
utqneZmV8LpdqF+/YvjLnHQ3Fs7cgzgWIgAkFGzPDZxuXhrYKrzHnG3jWlqLjj1W
O7QEsXVGyQlaqIVXEqsxe7Qm1dmLB3wCi/OZtTLgN+zJHOrn4Ywg3r6VhWqr1Vgl
iQ8DfndrEDcFU5GSVflXoje9p48iHCGTUTSIDH5dzfXKRwi8Ia12Y/8R2beSzOVh
yzd9VXDdoDi/3LSltUwiExIhlLZkKl2e74g0252fdMAWfu4Lt3LRZgbAcKnLOBsJ
LPnv43liJQT6lSwWe0nIwkpSGjtXfghrpCmfyN+azzT7CjJKvEpSzVxRyV3Xebh+
w/syIEDQtKOGTXcvjsxLfKwEqQ7PXEQEmXT+0a8wNfE6AguDm0ycCmPxxG1JRruW
nfkOMzbzogL3b0B9u2LqY1/iycFWFbyGD7d4XBcy6zhvMM7QikLXpr09RKBsbS/K
cttAbKOBXYBpNxb2WbegQkHWsEomlH7Z0yEt9LMDF5BUZnj0eOc0r2eEzVwO62rq
2Zr2eBmUiCUY/nZo9f7Kav9fkoR+0ZXI7IjdVZ6PbAxTM/n0Zz43USskIH3K3rup
Nf8vDbVBUBYRThXqQRjjBelbrPJkt2lJm0cx4BZaCBnwuUeh3g3/aXl/ySPKxavu
4JadfA1KhneIRoUXqbIuZQWk/PnzNMiUP2Bh1jiocc07Yap+4fDoUAfAA+Nwvb9t
BHTifouc8dYD3BYhZIqLR0DP4mDbiIFF1i2AJI1PNGDp+2bwBnKSoX2BNkQVpYts
2TkWp9dsmRJsvKzxO+khRC/3+ZL7bKWYPsB5muJvv6hVHQ3cWxcDLIsCppLOyAJ/
I+qooZjXaLi3zZ4Cl5RRfnQ0iQPUaO3jLwrt/ws+ZEPOWCLyEH0W146ByV9rXD2V
mwA0U5eIqQxgmre8vNNHJJM9f6agorqNOiaVsiVnee5vZosvsSaYmF2IY+/uXbqv
wW8LTtTxuJV+uXA3W5PtF6WaIhqincbwJyXxgRmjwkgsJ6WqPWYHmt7ZbY6qDssF
ZRH9TMxcJUxGuOxZRN1/2FVlpnxMFKZFn7d7oX7oqVIV6Y5W4EQswxHxuM3lHlTH
9n6j+oYY0OORPZ5gsNBn5QRkvSq7/eYIGAKHTgKJd0nlUCEj79H9Y4vaNT4IsbiJ
WyHi7f9Vv1WySaPai2S+rZVE8lBt9LGfGJ/LEwD5uyIgq12PNd+qZ0ajhSTXSznv
HxnpJc9VbSylw2FGmna010sfIbkkNKHEaMb8NjdYQ2YC+rvzOoi+l1aYZzhmMGVO
nT5gajvzmAVrcmVb42OOzM8khTbRZ7t733nZOuTLxyJE8jfmSvHSWM+/Cy8Ykze5
3wTf64QiMzWpjU0yJERNc7UT9sw7rFnO/XptdPZf1kucUPGaAJOrhw+VWK4P5mWX
dnVXL6zjOZisVq6ELegS7i1xlQ1M52W2g6HxwuyngxOsxPmtb7PLuAK2irDd2zUe
U5h4bfgn4lpxGvNIAliF25+YlRg06MpS3wpgQLU1wZzz/ep5GAwCsEiCfoU3FJdr
aXgfAQpYIM3Fa8abwi5SlmJ836bZ2Qgg92+x6rEqdi10oAbtsNAcvtgbfkfMiRxi
gm8mHb4foXL/lnqM8ysiNU0O+1nFeLNcjeDqJxjGG2RgDwvLd/sMVtT+uFCpmzLA
QqkOKzATlWoiCfM7aD5TqIoOTVSj5p0TXet2jT/MuUVRuHNqOkZkPVVgcgNkNESD
QD0T1sip5Nyf7IAnU6n3rpLv4KOJNO5Bn1oqMIXtqGM9cVcfZAltB77feWASc6Gj
pqoVz4NoVWCjc5Az1ZU5Up1fQxsXDVdk0zGaOpQOZ/tJ2HLy54FAiAsbyuCnVZRo
KfD7LrjGqB2Z9lUX6M8/YG5oADGZXgj4VuPWHwIeLoju3ZDwAzbL4S6tLyGcah18
jPknG/qSmplFlFhzXZNjG/dUziCgF6d8p0gnpmxevDnk3Wv1dzyAn8zMsLADKcEE
qMq6bFflTPO4Q693ext6hRu3gvEkYIqLpwXbKD8qkiREkpG8ghC9rooX6Hae48X5
6WplXTOCZRhdlW8GA1JQTXPfenfVNmNc9nfxrsJEVVT7756hegqlLHdbKV/H1+h7
9eIQ7OIHGMSl/nvX0C6FRB+QBShwO4iCPoBrPKs2dorelwvR6+iDW0ETk5112q5P
kzPRndtWbSVhvXYpH3PT8RCjnuTfm3M2b4Se+jiZ7SMRSG7AOiWFrOhH+mDJ8kqA
3WS0HAzpLWR+ACBcSeQlQPmZtyZTpqPIwtPsuWslNjAzr3kgZxQuNHKaXdChEFpF
g0ooRzVSfDrdWClx+gigVy6BGOBIrbGqh7ItzxjufEegYTk4Rfc6bEFKMdwSDk8V
JwoAc4ep5HkSnaTDM5GkABkcezIbFF/QZJ3424odv5S4QN7U67NnrdFEuKktZEOg
n09g/o2mHyVCxnVspx+dE0Xv1hrHEKuT2SzQJK1sJM7lS8XmdskLwnwZtQo2RDeH
XLwGemTHlxltoTehkODYrF7n8rLut3ACk4jXm4m7FcndtyloqxSFQmUqT168ClYr
BJZ+P1az1dJ+t7Ie/ncI2yZgMy2mAfw9NEOSHSshzlV8zrhH/yJeHR9yKkNDrJex
oYyKVRYH0BmmR1NyXvFQWkcMVpMt0o+oozzrtzT0n5rjVrWN08U2MZng3z2gw0Dp
WPXgsTugR6bgnSunA7gBG1ENayfh4jfsr3mokndyzKzRKysY6aSvaLCZtabnvUvx
3ozZM8sQrINFvJKoub8npk759RQ/Q2H+x70Rs8jvDkGLuAufkhpYMiJFqBLWaZ73
43WdFipK9ZyzpWudWDTEHMt8OWwEwtWYv1ZWy8Mj7Djk932uef6VGtZ9X8hc/FJR
jtjhjbcEQaJeWTzAgjO31va2QhIjhVyP82TKwzjXQUL6lwsMcDMZdYYbXrGYMks8
vgUSV+T7up4oKhbZlx8Aa5xIB5Ixvh1iCn7WqbwtFVanCsZizKAaE8HKZsxJANBi
UNb6iBvbwuWFU8S1Be/0hq+GfR0T/HKI/RJW1ClDa30aB5hNR6IG4GFeHkYtSpAv
I/4qX75/Z+OhRz/3UT+i1OYV2dwWenXlsHDmD6s66+lQGYqN4P/3PvwiDQVZeydu
QjbZ8jE+H+rcxQpJxT6oRzsz/OD2R9wV7df7dj4qL/f/owI+kto3YtZWEXYQoFvy
fmtue7IB2xJatiFfFM86nfPLciTxSABoy69hJqKOJp8iumsGYA8Jrvx/4zLduknL
tKrvDmjYDgRJFKHPBsLRwSY+nidnmoJrwK+/ZwHFlGvKDoMIOcnL+WlXBN+7h5UV
ReES74MMhkdjnZU9xmfn5HGBNK/5NQuseu+EDz43lVDqszFbKv3VTh0yuq7tNjrc
gt2ItO/DOVJaFtc2prK3hN5lGMm1JsiO8Cv161TtvPb3rarzvD4BlmRzdViMm6iB
FV8fnvdvrRg+lm/fMyqXq+DxmTlAzua+gnJCAAuyfz8+EHRb+VUYzZo9XXPvoEB7
yLM6wt268I2ABT9yiiMx9b968mROx/vMgrXlxdKcw01E5HmCsb7OLZUYooxKtWjG
aK54Cgu+/askYDfGko7AhvaTieuIG7e5loLk5UbX/SLLOLgWvt5+vBIKbFBVaDY8
AgNZefHeBBwUNGm+IX+7oNT6pGbSTsoymzSG1RA8viMjVVRwqVKSvI/OMJH1jrf+
Rhh8m3/1UJZlP+YdVoSwZiuGjUBz5uTmvv0XXBEYZ73KM0HPbNmzvjMI2dLmwlrK
MLgnHTJHFEw+38vgtHRNuCt9tiPjK4k7nhu4cVj+J02lqDy5IUD80MW6VRV3nbcA
RPHz9h3zAn/kBSi3+Oo/ia9iFqeyXmFNJ5anRVs1li+hbQfYaSxJApiUWATROhbg
mTLGBdnX0zU1LMeYiBsz0x9NgueUZmZ5vX7kqGkWY8heMSkwJ+xUohVpupwoa3Lb
MWA1AGhGopoMAujbiG0PmNz6j5pKrFXcqIw6GYgvTpKJ7TUNWLxBZKZzIoAV6qaq
pt7yTR7tnm7LIu1rRm+8BA10tXNM4gOz/EvCc27z4oI0SwcJEyhn8yQYhx5AYlx/
Dy1r3RgnlfRM5sxgy+9H8x7v9MqeXvMCQFWmZoh2Dhntx/U+Vk7WCpmfeQU5zvSU
SVtTla/1V9nQsdVOOvO9a+dGalCFXmwtbpX4ed3G2ubqqb4MJoWdCXjYpV3wh6qp
CLVri4BuRMpvnAxCo8EMXAhHHNbKyZcxNgJur5JVgFLIPL4YSK3ZsWiQB69rFaM0
5zx5ww0MON3UCIKbL56/1fZ16/YTPkT+VnGy1cul1F03qThb24l4hLCUaberpkSA
BPqRB8Zh+TxXCWoogCJw2c7WPHJh7hY8KQ1lhDNiioUdP91AM0prctsBXi3WShMb
P4A9TCNkGEzmmrluD/4EcmCZxftwzs15EPdEei9Uzs03sqlkFvLJSUhIc+la4SQ2
Fpmf455PbbxQnrfM/EkgqT+NudA0jP7iBg5RAoBzYDOKDi0cf2fLmcnKiAHiIsiL
b93Mi/kZkPzBFcSvsIKKaar5HqqjheADjbKyDJpqfPm7a1QN6A/lYtE1AecNWgAI
n6SWTwiNJJfxACiSwLlF2zDe8U6eC9skApOmItTPDdN/UcDjm7u2S6eWMMQ35tT+
bTXl3K+6AAbYImxoueJNvcEtt22jOqUrfn97/17SYw5pO3ZTR+rHjrVg1mytDY9V
qnt53hAGrcES2bqFWyqKP4+b6MHynzgn0PMm9O4pjOD+3Xr2bG71EqA5ga+t+2QR
yv6aVe9d501bzwKXpMfvsb1nmYk2dnJKuqfv+xIGzb2QlMqK3DoQMjlCMAniqyfa
gYujy41cDYwFgOrXovnPYaPmHZwQna2gHfS02fQUU5NmIxKQfp9Go05Bz5EQCx66
a2y27YwcY5KyE2QZUWUvupm2YSLcCQ7KPLftcHfFGij8p4KUZyBvXV4yEWmf60I/
7ENoZ84+/lz8OqWYVxc10uRLWFN7Njj4Ni4FD/K/GMQ4ZjySVmjrKtlk2RxNx4M3
0aYGbiL5CTqgQ30fNpkw8j/atb7wEjPhh0sllFg/5fDfy0acnxZQHqwnSIq6E57F
Q1ggx69WJjRnO715QEkl4PhdOrO8W2oGmhsHgF7YBZu5+DxaployJznPTGrV7mXK
Fp5Bj5LORrgj17enT3dHDfx6ne66yg0e4aHomwZ/Ewzh67l3tAnD5MKvsLTuAno7
1IoEEzZKU7z1JUPpLymws6QT2Z726+fI0ui46eb408OS3HDDeOd4ES7TJ/ws4eP+
xGq1T1n+jPNlNT4jF5wogxf5bjTyTuD4ZjbGckSHQURtSuJQ3spySuA5vEpLDbEp
cDRRmXYLZsjjl3v3Eu4SH09cSi8PR4XR/GtV8Wqi4at1t0ZIaO343i60QpsWC4Mn
zebttDBI85ZZMMs2E4Im2ESC9Iij0ZJUd0N2PV+dm9QGbcUzIgp/YGpXdwSY4DMb
ZfPQ3i/NRxilz3r5UQINyTzNY3ueAQk66zuoO4cJ3mmz2Uo2T+FublMJ9vrEYbhv
Wq4zDH3IJ6Yl08eXlJzDOrHY5iS3jGPJdM4YbZTY2xRRKt83RnQDlggto9vkAIeA
iNKRM2nR7Tb/tj6mJKQfJDyMEwvlFd1KxpASFj3mgA5pMl5Ttlk35kp89hTYdVaa
kdspO7TcJluO7gahuwak+pLEv8nhdwEQMMq5ltKMxFoEIIC+md5SPlPP3zZBkagn
qCbEe4gE0UgObzmuhOpA9MRctZXBtNYakA/f+0uOxXMkYAjHRGDnndcb3Q42EXib
FJoit0nf1yfitd4oUWig2GRm2mafXpr7FhrY3hEkHcUMROHwCu9rHLTuFI9BsfLy
xs8bbxZlHA8bLlIGFhExLp8Fk++3vUsWX+DEgJd4xZ2GszP8pSPESv6/m1YsaiW4
x7vhiu1CvGAqx8Gu4Wv7EBflvpaEQAiXkU+XAR6bv+zbgLLu2nonItL/7Wfqq2nN
UFPntGPN509mP9p67eUcfTAEhilEcUGS+z/JaxxTFgylD22E9BJ2df422SSzR7h3
4nBrE3To/mv2rKGKyFbMa36Vr65STObu4/8GAwupuiyJg+oEtFSLBcijR5OK/dZ6
uufZLt3voq1fL/GCiZtac9VLeEKJWxLGhCuSVzFwRQYbkoWFAfy47NEHMBFt/vje
fApZBwd32E+JWHCK164VYS2AaBAps6BSU1IBPaCBK7QJMJhkxT2a0XIivpqaHF49
hnyFFZXAgZQRZbnACDPSMdaypAhLVBRevkDmWS5vrVEkKTN8HXlNE1C0UVQQFm6B
B8qoDlcil/KK7+6WwE1dn3l4TejMIBzbdq+80Jfo7emXgTkiIlJc9+1y/LnxZJhS
oKxgi0BwrIGjAoGfAF8Vc71xk+BZ4zbSl8Z9XGSNRLkmZpIoIQ1pk66V0AoUTAOY
xyZch293vvID+yxn4GmPDgM9DlC/vwZxIYiouXuVbh4SuTiU9jJrZ9XKuDVjmNpa
nTjtgi9KzpMjLvm3VDh0NZeEV7rxBuA+Fn13xCr1ZUTc9V8MPZHjDI3foPqtVfch
8HX9gKQOSOqXXjQC2KSS+jCAKetaTmH3Vji8WI/2YmihnxtYCp6DcYXdWhJ+3g0O
8zpv1ZAAu9yJcmCFFlvANkmrqfPsQ7PgRGZCHKe2ULPKQOCpXI59XF8ITyYA2y/W
uKh4pVSm8F2P1eZCTghajv2AtEHOKwqzOp6RQzowYqCADS9Btpo4xyYQ2fgZ9C5n
60YCktpQfILAMDkOjCNIGuyQsKvm7Li1ate49EpEymW2UYB2qwab+RP3IuTjv+Gj
wyszyF2mYLlSv8TXJeFzKR3lolhL9mxLQ/xrUaF6BSpsz6RhaF1iTOScrkDGLhyc
AxSiEZe2QRe6VdCGeU0DmRzJvJWu2BlSxzAj6F4LyW0nXFHASly2X1dSIoDnhw5j
nKLYszp/UXc2f6hzdUINYGFLLNM8Vu9+GN7UlfDQx2gxW5dYFZzI5A/2OVsv3ia6
q/Mkic412ey+F6QJh3mOKYeAimHRkgmRkjmlofs2t2vwt3LGq25UtYAIhm42otti
Q0WK1VFlsqowTTl1E3HTLPi/TeJGpHRJ764yAAKqWBfeLQ2GxezFg5PsjXxlhvDm
M1MrKQd6o8kUUP99WYIZi9sym76dRu3grNV96m3M+aucw9b5R1xKCs5IOVwN+geu
neGnu8j+2Y+5+x1qQ3IlrHOYxB/+jt1R3M2p7iHJvKKkkZpz8Ewsc3raxAyo+crz
Wa8K16FHC4M+k9GlO1NU8PrZljSiUjra/Vmdh2TCOEyWWSmhKIxQBr3ju4TrB82U
uM3c2YtTiWggX3aRJVvCl+bLU46LbE6F3Ap31QpF1txMBb1BtLuAnd45DyUXEzqV
kEYahoJVmVRGX2aBRleoBNF1RW9UeY+D4nx6dQaJTRHyRX+pJK6wAE9lu1/KXDKp
Ry2EfmHEh8QYta88yIIxon5cnxtADNtZxIJov710prMgIci2IyznOeSIXEgeqgkl
F/ypqVDUK8aixeuvONkBjbb/MkYRYyFczan3BBeKv3gSSAat4rjaluKR63sxvdk9
8tPUryDMbidaiYqdWiepHWL9Bp6+onfy6KAQ724od2la/QW51BEyS8MRnN7chDBR
LmV0lfn0nmtflo3TyC0Y5+3ucdF7mcPjRzNuenKN579ypF0+nG3kFUxjOURLeib4
DRn473f/9ww1NngYlrD0zlQsNAwD5w0XReWZ+96p6f6bERBxQ3Dan+tfULSO/xGq
J6pUA1B9T7jgbEBSxHy+bKKFOyuxneJhbxbLfhGsIZ4oiag0y0T/xC2fw3cl7QU9
JG4xy678poxZVUbHTkf6Tsqap6eHizzL+PBpsurTD+yaKKPY+vsNcBdHVkfADCAH
79W7TcqhFQONw39vb5dluJwB9f3SkKWD5OWoTrwAaiLRI9VMVF9eJYEnU4/SWJdW
Hrwz4an8Gw1OSXOQYw8xnMDzEcmY1Fw8ukSjLZde/5H8AnDAGUB5npTcDBDtTLbG
o5u4lQRRuJXdaLe/RIWQiHzBCnpK4KzJxs4M4heOBTa5dxrgb9/fTrHsY6OYLArz
LDLVezFffws35NNbRy9U4XkpNaWfC9wTsXN1fm1UAwSpWi/04X+w40J8QUH171f7
FwhxqqgBp77FzC/a0Ij7L60cvV9WcM1zqpbVcWUUrOBj64KM6vL9j3MshWEPgosb
qmiy8Vh8zRAKq3neMNkCgP9iNx0r9jk7lfbdMrm01Lm0HlMjD2wCc0a8hdzblb7G
IBUa6OP5DP9jCtslikDH83rxohJsEGveqPjrrZ3txQKs25AhCUVCjspxGIf6ehdV
F2V2oVqw7RkZ3COCe+cBDC9JQFqSvF2HHcjNWv5z8eumNb6eEpCSucH2vIBZsrRa
I0KI2HWjRVzQcOUHps9HjfDNdY5Sji4CRX9SMA1CyTO08rtIsvjp+0vzY1As0rPi
Skmp7B/8kophky4WjvQNAeoP6x2GcrGYJLJJ6JvQOGAIcx+utROaajRBeIRpy/zb
//hbW4/8Cddb7uCWeV5RqnVVGVge1tSJjOHi1G8DzNtXU/RXv7O4RZsNkmq4G45I
c5nc8kNRWMS5XJM1xIjqTGo5biLOdhJn8pxUFsDpWP5Dvcb/hbE4OLV378Hp8VQp
lk30wKJ6fzYDmZJ5d/KYb1P9rR97jJx/ra2EMpg89eQY41J+ZkVQaiqDVZD7zB3Z
+nC/U2mA3BEpTxPN3SOX3smUY/B2EN5cWy3Nx55Rz7nuCSfMaTrJzvofo3pdInCU
NyAU0N7Q/tauiRkUOfZD6RDKuM8oKkez6vwnODAVaxdwGV/zRWkAly8Cd/iZBHt1
FGjyPRIFcOBJ2nzwkHXoGg2V1JYWdrpQKEMj4PisAQ59j2A5z2/y349IxuWPVyY0
RVl6w6nS3odEoERlkGPV9MrIdW3a7FZBymE6R7pCvEn98cIj8YYDlSLrbvIEubSo
UN9snM7LAsEz4n8HAx50bUDS6lyCD1BUxPWNAKrl/syGhz79+wQ7dhimTQ3RBN1i
oZrC1sZNPXaS8/9nQXjzhcisEBCu13DF7oHXtN1W1H51hyXsX1h/kgExJeINUIDL
iTCcyCtHDyeOCFEUEb5Gez9yN6JSwgpXQH86Erssl8LTAgL7gaKmajbOpBUD5NzJ
ilfjxo1d1pV48SLS9j6NGRp2oCPiGPH5E3PmUyQh2o56wzeQoJuy8VBf5NXHvGM6
qvjL/tSjyl//yGdTLJSJ2qt5eyUenzukNBLp2zaCL9wlY8YlADpjNw6f4c4BKMZ9
GdcotMh616OD8XOJP8P96TAPnozkie1KDhltpQU43EfZuk5RtJWX7KAKlyoWGb11
8yphVEqjQFgZv0705RIw+CsZWiplseaBCMLaUmNtMVZqo5z4NlbLPfV4CUbWfAZM
rcvqEKFYHZa/jd9GAIbMGCnlUBbp2XxoL7AMSxq07DFrUBatDcJjIAABQV+nOiL6
0GpJvVosXu1RIQKRtxBGDkRahQujdpNbEBJa+X5dJFq2LOBDLqhWEwhRG4c92N1A
bALyoz+H//d3SUhZuc267qv4oUvmK2e3Taf6+SpUEKmPI6qOW51Pt0PwmEPS7RQE
ABLlvy2u+RsAVsh4d8IZvErdBJdz1RQOwB0AgY7xegeMF2HQXZ5F0CM0EaSyOcVK
u/KxYKD5yD047Ikus/p3ouVz0xiSg3V7VDvwznX8TqKZ5N1jCxFq3JYInTCMHKuR
hqDDwfejfI9OqaDn6y0KXCfPktsZTMeg1OAwF/ckpLBlTvvNE2SY/w5GCzVwZdD4
N79raPL2Wm7Xn5mijluNg/LM9mckFOX+bevIdHdyWQ4o1cpwCKZwIKHrD9xEqtxA
vF2zocM+YJhkwQrwdumIkx9mjnBb0bXbGm6wkUy1TDqoWTg9vOOCgxWEZPBktEow
yHtc+b0Ul5qQriG2HYXkdhWyBUEN7kZTerZVx9sLS9LjZj1YBWCYycJhi6C0t/oT
F3PZv1QcmBbBUwi4ynrc+n5ZePyiZ9FoUbe/VGP5lT1tDLnnd2CyNPJipWDWfZLc
ie+/tzrhhhWfHBpyRPSEGmn9E3HJK04o+kHkZoEhQGzLme5vyqNb0R9s19tDvjrB
6nBaIgxCjT2Bc93wHY821OINJt4SxBsTqMSinYyv1GwlAEKFa7uYIQQi0gbq/UTU
yw4hLUdkAqEWCDnb2O4OiG/+j+Bik3McLU1gcMMsJ1xrlz2uVbgQVzmKO7HS/Ls/
DW8pMnPe6h+HFnqgX3NNzVG3FVSipZmIiW4Xxv02P78CyOE6iZ8702eO9cIgWyha
Y2oQ3lCy08M82ln/BYTpT1/s2HXuy6C2hZ6I8dXt6EW15tvgauSItRcLoNw+E4qI
NPogXcGv3WfgwgldKeLQVc+Oi3mwCivUMtNr3GSIFZgtqE5cOkfaWZXI/aj89sKV
vwsNoBBzLuQF3glX9gZrVCLsl0eMebAwUn/Ld9+zxEUBFA85/ZD3u7z6jPcCFVrW
onahrsxs1rMnCTxNkMxtIof7vV4siaDXXUrreKCwrjPmIV1LeRrYO7o6CLhD8fi+
66ouX35C077C8yuevTEWHzOmAr9SwQeEz0ocVIzJnrIyppqQWZbuySr0xvk73cjS
m+sHE9UviGna0WQdfMV8wLSomZKw+eXK6yl7N9BfsCHnda/XcMxOzhNdviKnJxZc
DLam4+u9Iq4lWhvk+NwYJqzNTqwgOYvwJV54T3RhZBrVKyGIVqmvakuUjS2p7hlL
7bUqz7Tt7W2p3EHgfQtPUFCPE9JBYZP58FPosaonBnKE+to4yKvlcJWeqZSEG6Gy
wNbLYYu3hYnSO8aPV17k9KaOHR6pMWM4A9UvSsXLeNpOnMgIpYUKG4/t7MXBXFz4
/CjYjjrhKEHtb18T58rqCukridM3DlYRqeVZIzOH0DZ6QC/rGu2PwUckiXm9R0BI
qeGjDSVzbaVV1gD8G15P6+vcIXf5e3ug+mxQIm9hjccs6n9S382LMlM/dRic4S3J
W/uhG2fRxVJm341s6eRLJp0ROe5/3VGE2T8vLJDF16m/4BV9BWTuO5dfE/MsG/m7
UM6TD3M4PQzuKguFF+jcp5ODw6xfgLMbmvDc4k+I6lL967HEPHrbo99/GZlZk2/j
6/Yi6HQHBYJpfSLxmJbsRbd2XBK8WLIiBYRom03Z1c3VJPAoU2/fXFdfonxo7Q1+
whzp1BhcVANNdT8XWCueTQEn2iXW+8kQxC2VOZM46cALhVefpNtdB9qiqsXskrpY
0bH2Fmep764Z5co10kO0QhZO8XEG53Y47cLrYDgaFpcg7HgN4Rh5IoSpEBLTHVuq
icljK8D/8JS9z7RTw0Ls0nnzNquIOaqvYb6iBYVr9p3W6JfS9F0iZGqgRdfOeLJo
YMhQ7SsFDyQf/Gow7uAvYH/yC8vsGyd7uS+dDf9O7m6SVKxnr/JK40hbZNcbH1Lm
Q1Xx/4GemKCuMZxgDtQIwCt28EEXIOwL7nXpyneny64g9dA9ZqOW5U6yNpUzTomY
Y3+Z7g5l3J5UJ/5+Na9tR/MWdHYj/cMxPIZXtH+EDcqRTit/pRgO7PCC1JTtyP3o
tvh4CdAZl7Qnf77/qW7jZyDTiv9ClkD0MUl9nsu0JeKd0zfDRvJAlqoBHiIl49Dy
0JZUHaCbUO0RovFsWs5yHQAL1FH2mufcTAe5oeErX9DOZ6jhtTd0PWlseVR2GORL
Vb7zDqWZoAQ9iirq2N0VFyrVZnZ0stXCgDWyMHPlwABjnnzsA1KvcnzZ9kGHw/6f
sCeayrJbDqPan1d6jwzpAg4TIkBJHnnYBXQKIhh1daaOXNjMJnekk6xCYk705eSn
g/YZHm1N0/lj90MD4nPEIJhMAv4gqCMGeAbum2udwzkvbPVjnBZS9V9eveH/R4yJ
U3zadc7GjSS+Bc5WqLg6oeNHNNjfJ/lyrx53r+79jtivIZOQt8jGa82+9+GqZI0v
k8vvI6qEOkIDsb63IAzlnN+EKlQ3AyeD+WFcKsrvErrXhH1KRpab5Bz8dMjG8fjx
m5fS0BUUp3JVma8rdljLX8B/W3V8icrYEFb5gE1bu9weas2m9xGqXKW5yKYHnOuf
nA+tE3w3jBDSnRqWzzelipY9fKXH+GPTir/TUwWPwm2iqHwnWMencuEfgriD7Ay7
2J1pM+Q7VBDUu/hXVmS7uBbfoOr3Huzyh1oXdHECzQnV3zriqJ2vHQ4R02+onfwD
GBLanLcyDDGjGLg345uwaiiKfOp/CsmJJzFgXYFC8LqnpP7CytqXygKA6ac6Jb9O
w4GSOTgEJXzwEZG9JEnRYEtnV1bAKNy0ty6RYXOFWM6dO6M+WujIvDH9wMUZiwlc
oIvIn00b1Ycz2gZ/sCqbnlcyannW/qjdHVDZCs5Gm2crp3aVPOp9b0uMJxfqT74/
9S6E/1AP7pb/C2yuFTo8mNGrNEpWZMXjb08u1p3tvL5ByXcQ76Q0Ued/c8uqZAMO
42sjImOLCbxeurdyFEi6Z89/RfWgXAwov2wjNgboa8ZQqqi3tRd6TAYLIQ15ijxD
itwGeHg+nZ8M5zAoRg1wC17wFq37lwSVqZvVX6Ep+3LetL1DOHF+yYehSJMNOiPu
4Yykl/DFpmoS5IrirAegyJCOLCTPHdY1yZYefxr7DQ2wNFkgz+GEhQRVKLsqc9rT
exPYcEtTcl1ClmalI55kRsqVMKPKAk6q9qts3Wq8Wu9vKWULGZ76jdwgiHbcRTeG
Ln5F4XQmsyiQEsagxKct1SGadvS/wbyUiqtXQBEOYe4PlgVDK/mK5bwmhPZE3Uiq
+DAPEJktwnSpzseWgniaUKr9GDdZjeF+5gjvrHagRsxRroD/GV62tVIedYfG/1rR
rpBjWqQBr3xhFIjX9nfpfakarstXGd4neMMuFEbhB8faONmAy3qxB1Ih3bP8IYtz
2XCPZhUvfLBakeLrXON42VCdPD7GkobZxlB3jIzuOZA52d7K3qwbjdhE/6hy3Vee
hjnLc61AG9HRGhwAPj/CldtsezRjG1f9pS0fRxZtQh5i9tdMaBCTHNz/Gm6RZfXt
tSIOxfD27bz9nCyZSHRKBcrPMIU6RXcmC81nUWRmBVlJtxFzRFMCX1TqARDvltn9
lKxnNbh2G42e27hUFXGFa1uMlPThZ/E95FMfVwZa+XmYNUeE0v5Jbj/JoTKRodkD
teVb6SsNe6ee7NJbAERPkGcm0b+o+HxK/jGvRssPF5pISAnfRQyGPfR8MItH9X57
RxygFAF8KQCMWWK/ZimUbNDcXNxJezHiFkokdvdF0kCeVjONU6AylR26MZTFeuHc
4pYXmJPrpDjLSzNW8c1otk264jNC0rrofUlvYKm4W0cnF7KFsZInAgt/Z2ptutcB
B8e0X1L+mnjDgmYH7bJvgu/bMHkyUpMMTnNSyysCBB6I/TA3pE8RZX7haoKK69nY
rUypFUoAaEjbRiAJ44t+RHBg+CavztewitiNKyrKQW1KgrJf13ycX7Ulkwzve/LJ
IOw8kV6X0x/5rNr+U8p7RL9S17RUYDs2msCCLfQsscUDCf9R7Y8T/pAXfV1pVTeW
H6ieFvj8T0/O8XutltPJfFgqTtpuWzPIsFzGEjSN2rtKDDIjnElQ7d/pT+tuAXuk
bII6G4WN/JgVe5nInSpZitUBbXDA4FgduB1qD4VNIhxJ2cbRkTGfqPAoiHtgNXZK
74neK6WB1ytVpI8FAkznA3Hw5qsnoGmk0lf0bqLTqLDJT5Hqr5Zv7vkorLOXWHmu
XMqDQutU5lQqakHWwitR57EItTa8ay6gJ5MsVYbyFM6AXe9UAgakymsKA9cBftrB
tPMi2JbIkR3lhCoz2+QjtffcoguT0lYMU/V6tn1FgrFG/7nMOzj1pexOIa2tgERN
aRPMbSeofkstFj6XDvcKc8x1BGNaP6kmYZHyAobDxZUCCEkDOm+W35CpbmYnFBcG
hcavM5oxaP7pg68sq/cjaChZkx5Hy03p431G/O2Vw3KqOA6XCa5yBtVP4J8K+TUi
tZ8Qmy78Z7AxjEZxZ5T7KzjjlYW2RRvpeKvPmf76iRJhkIja3MVHY6Cq1J/mhHs8
qdmAd8Ov8J0MKgQey+yz2llQApyGNpF/9WenkQEO9uG7uwN/xV52TboMnugUFWk4
Ii7buShWCoVxaBAMt2nj9SMGBZPVjsl2lglfPwkthhToV3zEPuQnvSDXu8nYLJlR
8IkYB57QmYEpm7t1GjkLwd71nZmYkicTWZmqARW7JfD64aRNzP5W04kTPiBVrqIQ
BkxARXoeAiZLH22PBC70R07sVJFATI/ybKLoaQV3Sz2X94EwjLJJdrePxX/VkeoB
+ccCi5xB3M3WTGnTrKazQqi/Q/xwyPVUs1I4YKGQpK6SJSNW6aD/dlJsKa2bUsUf
zOWEIurnjnm3u9VRCOg1Wvuc/3DWgvpmet5G12obeFMrBI23U9tAJl77QyliPZCs
k+i8XYl28rt9eXJSQGYgfCqS5G5goQ0jXoP2pvmly0P3A7eDsvsEZ54TZWgnd8Ed
81WSKNOwL0LKC3OE4PKmuTx+tx0D2u4kHxAmg5ShddASWZU1aQU9dKW989dh7sjE
ezORiWOKncpSUUjAnYTrQMtezjncjkERauVYveJThwE5VtiU13jqmbudnoFyYYAQ
gTH7x+JJbU0J7XTypBYzlQmmgKPm1ad6Y+TpfqjsAdmfcfXKQqBEoGC9fPXvH9DX
iy5w2D2qjSzteRY1l9Bw9HSlBT3J5qGJIbWP2QrsA936we8lq/aQNasjBD1pKV91
EIIXd4Aiie3EbwHngkHuH6hxLnFLGQFcqgR5M37GofIBCoWqZa4IzTJVfTf0jBcx
KBObmYId53q58gIk/5EqTuRL+BHXxFQt9I6yTy8wji+yXwAA6tMIXBwUTKCozsYo
1a/wOLK7PprXGLO8reyR4qsI8yPM+R35fp7jDhQls67XkdSdO+7kBj8YrQnCyivE
samoqin77F8Wu4v9rWnqmHp1UJO8piK/3vWV5+7Gydc3WLjhZ/xlpUJ3invMwFnp
fDl73mSGoYmMVgOZUDdzEnyxTk6qUwZo5JwGtvkuxZuWKZC4Dm5CkoL/8dx7Rems
38+9DuqZX+AMFFk1TcXQRF0k/d0IWDdwFZ5u6k6GFgCscqC23YjGPOM+G8Ya5z09
HVWmOKn44BdgzzTUMPSWZqs8P0Pa6UME1LuXhomL0xR+HSgAov9fnecxYNGAn9cB
n+bplbwTTvxngEECdJy6Sf+m5nmqpiVFg14RYEupM+6cYJvpu/PMQ8yrHU+Vfx53
ao8b5W0BHnQUiJli7Pc2/xy75ZKJsanKORtaOhYWvA4L3MNVvuB5HVCloapN7cS8
10sCOdpM2lIQsZQY1nRXNF9PqRh71BDsAGRleSk3+vj+AkGvcC/FeZvLakQlKnDD
DyLXtEa/2zusg/Lj1qTNJ9XIb7JvSCZBE/Wmv5oYZm+XZwjJisidcRmBv4YhS81x
bI2wQjanmHoHwAsfzsvrUKqOYTOQpnea6wfRDgmR7eo8S9B2QAOoqENwwo30XFid
DRgX/DZ3QoaMK3Y6pGZ4p2EGc8yoGKz+xKUmHIGzv1MABNWlQmtvjhYEN9msGiFS
WNGKhtafqzf9XuRK79kl2maoH6CWhXXlxNpY3JUqwz4mf4/hrIj8LwuPus/rMMq9
rlh91amNjtSME5e5CxpTqKt1tNJsnbSqrjxYzQHIgWSpz5qtPMWq6AFHdJjX0iNR
SR+wxYEHRrBUaGGqIvqaYqlYa6EQFxXjNNhyG5ENMDcWoms4Iw4jGBoiQBJ8VoHh
kH6OdVkbopbHDOFqEZDwCp8v5ch+uQxqXEKlFd+T7S7oL8rYQETE3f36NvqHB0kx
ktFS5tLCEixSoiikduCOUTb70IqfyrdAlS/8pN39R/tbX+jVcp5UJABM91Oo8wOM
rAKq+BpWrLX+Qx5vkx3mVZG/6EUDPZgpTBwR6W8qZcNRYiX2jZaXWBRP/LsgC0F0
F7Ms5bMr/DNAngF9j+CvJlh8eaEUC2R+3OFOylmNi4F1JQlwD20/2w+ClZoJgCtw
GdEfmPvwZPYhcl7LaSr2PA5TqF75nXlOPnoQ8i+cy3CVcRBEGnUanfoOAR9lwEvd
yu8lAlM6X20b/IWAvEdy4HXXuP3905LENE83e4DtZaGJR4jFqyaPox69DyUxEA99
O6CDGf5SrTc9b/8l0ukTCFT1fu+yaXDJLBAV4sbLIcEGjSQJR8x6dKswT9cB7xia
AwTo0lf09a5T13c0riqYAR3CS74iW7EZzY2NjOhNXMmwGHjqSS+/6V0M5e6H4NVb
2Wm8AvfcoDj85851XuMod1BDUiiJl/WNefxgkHTmBKOiriyseEzj8T9YxZTKQyPl
zJcag2NXMbu4OtQXzb9voPuOcjzuVGVQa3nAkC1We8vbR+dkqvknbYgrA1HgqpRz
kiz3hIHKxW02fFSOLVPVD01Nx9Cy91MfPSw9ioyfgk1HjPq0qyNrTjKBAgcRW8RZ
X2XsIhvFCXHu1HtYb4FWRlFSnQCPmgosty3gqKY+SHYE15e+clgcDQRTF7e9q1ZK
FydIkmRFrsS9kfy0ktv1UCH5L+pzVYHmmtScmvvYfDRzF9LumXOnKsFWn3aTrlpO
iEPXjQcXwKE0src1FmVgSI91WAX7oH07yTFV2+GG7wbPoG0Uyy4Ld/PBupakknWN
KiMs15P3xkpYqsDKwetagdcgrJ0D++2WDx62tpVJG4q9MAUaZmmlc55NqKF47Rcs
uvCRHwBUC9srQ3NKG2gHBSBBW1G+LSJvCsGi4e++rNEM6gKpwBuCbhLT6HOETI2G
m/sp61sV5SXyXLKpy2tgo7T0K2ELKnBUi8jMEymdamC9BdmCniXGIVq/7Ya1L5Ak
egCOmGYqk0/D26D+N5BmWaqx70a40ZJZ/6wUfh14C//Y0k5ziU9qvKFuFERjcQvX
07uLPWugyZKuLx88encg9fujg6I5XwnZvYgDqbiCOygBGfO2d7jSAEf78pWSPqDx
VlOZ8/aaTfPvwahOLuBVlWMvLD1xSHdc0aggSPv+WIXlFwMTm9FG5RbjnHFqnp5L
bnYt5awCNmB5bh2PCvcAg3FSe9SCIL5egDzUtr7LMgQbjCYDFWfXmxxjmQOoWMvR
WVFS0rwgmbeTcHIhqBaGLKvEkNfV7SwRP5xwWgQkst5TVvskmY+ikY7HKb9BQbHs
Cy+MridbO08ZJ1fz4u7DgTNikz+4Wt6nzdT196ulSKRSV01lOtT5rjwcXDPjSgIf
uzVDRkh2DpLS5ukwnkSHBeNsQ74PLB+CZA9qacMnwcOF1SsMoLsXKgEa8YTrO+pW
eCHMInZLHttoCLCiaE6dfyBsIw9izFctz4CPaoGpm/3jvOWgTaI9njqFq3eb+Uq8
xRHiKS2TL1Y9ehJpRp+V0u3CHPF0arR+ejugVwMLxIeMRlGHGI3QZCyph489FIqq
JtIfFRgEMf5TsT/mu+RDm43HZ4oKiCUkz/+QOcXCbZN3WoTuq2r9mg2dn6de3Adn
mdmFLciSIsdZ3MtFVFHBaibQ78l4nIqhryal98wGb1NtJ87TSmu/Fkrvv601xkO8
P0gSbVnRLXH7Bzj17PeqzR1pSS1AJrfiiTNNYiSk2E/9LKnelNJ9FFBKFR1Dr3Uh
N2xipY8BoooP/z9N7P3sXQwDjNW2oBgxDQmyH3J29uUkzfG9Q498pGiGSfjCz2+s
jaFOz9KIqDFB9Gr0JeW6fNK0yR9rD1ZhlWKrpquckX/mqePko04BAgTjRMMCzWYp
rbUiTLzBfvJUU0YWuXse3FJn51ljZpp0Ip9t9+ExXkPQ0m0mHE6qlNmizeXGM+Kq
1qj55RGZ+kyfO2H+7szx7INaLZJgyK+QWvy6fZaIwcBGOEd7xlYFJmNGWIQWM2/7
hltY/62F/5ia4usgmaAdVdX6jZpoRz0J2FvpUbWFcjajRKVFKGd+A04VzSTkka5V
dK0VmfXAkIbhmSviNuuIEUfijf56NB6TezmxXFVYMu77pNNSC5BgEwT4OwjI2ptJ
sMAn17GSgC8gAxKJZQtNHJuhNOhAlLvHuMrEUK77Y9ULDU5BaoZHZWmHLlUR1hT8
Z6PfGo2OaaXChnZ5i0mQlfmPOcDLddJdR4Lm9R5tYNQjmD8eFLvRDZhvz6SGWjUB
f1iV1pm26W4oQhIj49q3ZFSb2Mel9I6XvGWZsrI5bsRqMsaZWc6kmGKV8w+jtFfO
9EPoBEeuzINxto3CyIIQK6nZGWVMHeXjbeJ16L906i8gI8iIw6La3guojQ6TCdCG
SAGkXmW+3AgcsuBfnwLmI/SlP0CTomeENxZtu/WYGjKAlMazjydxMv9QNiWt76MP
N8ssNAvgh7khSTj9ymbNBssdLNEVjFz/xCpwhfIIV9HvS8Au1ihB44I0BoZ297a/
GTLIYSwFUb2Ihz1FwxBlhCxUIMcwzNX2rE0CsQKGVuFpg3rR1yHTn8aiMW/HWCiJ
RZNiDrzf5wZuKyQPywDlm/RpD3zP59Wk09GtudDWnBwnu1SF7OKL4lyVFlrkit1/
CyggGM9yVFGYWZsBXPirmO+dVfdUE6FERVFX0VsXxoO9fcCoyav8VkaWtL3gBPn8
b+arh5r1qTNNKd2A54tPwDvWwSRZ4oJ/tXP/cNqEQD2Cm9yZHhy1wF9shjZ/ErTK
tP3U6Ubs3spRZFv7r1vUYeTNocNX93CecCZveqs8337fgG/81Xv5rTw9q0WdSNVm
RdVOEfRKR6nveL5CQpMtaXNg4spvh4QrUtE4hhgTbH83cem14HJ8JQkQ4wttmOyX
w2rqRObBfh+MLnSQ/BYWrliSCGyg8gBs/hX65Bwj5WehATS7aMabb+vRcj5Kxgf2
zA41lydiQWHp92PpZH6EQXL/QXT6u+77628hqvyjQc42ZyCnpQnYDD9X8bYwanM1
bpHWO9OkvFPyUwVwfo+dcOvjHfunm9NNnda52ziZr7/O8M/gEX+qDOKI/+OAq5Pt
sAtoMh+Wj3Az44Pd6XuAkBzw7ZH5t4ChCqTIdaTw+SrclPbd1BslSPwLlLZvLIWZ
xPepaC0VIm3PLB4h7PKNYutxPOilPor3Q7tJbWK1oeflHLvKZWbU6oc6bAdHzgen
bMGmcoujER4BkNLeh4Vr8Y37F6X5O9DuYUW3zzkCzj/YbXYOEDtpB4jNHg6uweHy
0NYM5QQlkEZ+hvw9K6z+XKyWKQDyeASSk7qASrIEKaM7tHTnwQsuN3qf/rD3XEkJ
upwcGJzdKqs2knWVnItEYp8SLv3pTf6IBojgZ6noJmLC68w9MajcDIZ/4vECiSIM
froylW3gibW58m1ZqPtTxE7lFWrpQ/b6KM79yclM2YMunrRD5rbfIb8/vsJJNgBq
uKsezazW7XNz0i05Gf6GhOZJNwjbP8jigig79h8AGv2X2uyHyAkWCshnb/+UwpkU
igBpiqn1WwL9YQ4/aYD3nerNC9oku7u4HOh2kxbrBgMaWQR3aI6biaVe1+H+8SkR
QkrVDGflJTKnBErz+KtKNfhEsKKudQas8ez02BiRC8kkA5MerBjUMw45j29ZasHB
bgQFwD/fqF2WfWyHM4/xbJisSTi0uwD0iGShTmBPOWesFqCLc2pCnX3zRDZzsTAj
cd8+JwVcINRuYrpsK8DC9EXmyRTF+8VgQe78IOYSc2b7aAeF2/TDlKapEvuScHSu
neDikjdsH5smsW/ZCoALOxJa3WtE49MN2/W0IkwJtvU1r9pGzQ5zV1ZozKjP/eDM
+NNA+bMM6ttGcnaa/fRDdOSwV1BUPVIQCPJ+DOzjZfasca0jyUV2iAMjnDcoG2ZB
JxXsjEs3aWW2GDRK12gCuII/GusVevJrcriFJXL9cpu4gL+bykS+04ea2m+umUmZ
W1HLs/wnNsVuvhMzU7IOK2KFxmu6tuWoEgovQ/DKc2I63Mltsorx6XHt7X4YGSa6
fhM/M5NfvC1qT16kZajl47kAr18XGqS5m1xNuwmbpQm2pW6cx6dnPrb6cUyP1SAj
Uumv7L0247gNspPdC6WZDj3f2huILUk2PttKoW+pO4b+BypUF1CoYSmlbePuZi2N
f9lRMCu24LkUO+idShKZrIStODvHj5IF8H9rpiNuJ/rbhwmxp0iOTnaKmCFbBiFt
HkcUnh4PlzAwiVdPZDARXgWxtVOz5EWLFkJFiqGxTDH+2Oan0PjyqTyd5ltm+3uP
RBt2X/1ARfMo1fsVovjTqqgtN4smjIE/HMcKC0dTQrAkaZqu2iAP8JKfR1r8+1Dg
PcuKxCMY9q7IEEw1TagupRr+ZmfSUCmanM5qjfARE9GEkau5XB1bM9NNUc/hCu6b
vwKKdesdVTocdxSXYS23iUrSnfQXOis+VJItALmTF1fBL5+GRomCcQVRSmzoiefM
KbyEH0WMcd4uq4Dt8C2plq9iMlILaA44GWznNlWKEuKFQmKGhgURgHYi6ROs4W1g
A/mySL0BaQ/+r7X3umUlFS9xsUhTAD158yMIdTJQ1amUJcWPXcXfjTY5XPZY6pFF
JYJhIaZDa9eYMyg9Nca51PwvTN9NARbTmHSqJuk1/1cDJQT/hy6LTypV2HhL/ju/
jBcX4l6vcYGbU+bQ6VNz0rZrNsUqJn5lWIYO+MIWZUxwfRDY55O7y8sROU06q7Bw
rsjWCB3k7sV3Nm0FyDlLaCM4MvugPFdc8p5vkKFqKIwyZ6gqVWOWT+YWMolAswVo
juGkzj43ENLODiOupeDIcTFKLIqwtyJBPMnXCIOvT2O5FSn5Gw0Pg5IvOAFYoZ5i
5B9RALKoCFSZIs6GORGxWOooKJ9tH0qqklN7XUmCHpQWoYqG0ax++Z6s8jElRxeM
BSRjSDYjJudnxoUH8ByQd2poJmUWAYIfpAB8b7gbCbly3T/5Wpb6UsC4Ua+Ji5WK
KW8SnT0GHeLSb5MKm8KT6Sv5xQNTNmZDvvLOGj6lgjabjYxGNkRrNDM0QwMkgPlW
ZJAIKl2twAYTpgYzOlu8QSzeD0f5mSdjOqETJA7EqLIdQDOPUt9rSV0fOod3K3H1
JZVZd3IJSuEY1scf8JRRx4KzT22moeDDcGi+IYJnA1ybbR4vqr0X9HXgd5tuQGzP
ymsZLmoS7tOvYYuQmG0aBzT+vFvGlKndIV71vpaambJPHt+7riPRBmhHaR61cpB1
W99BX6mEdU87jSmXSiN2MaFFaOjTSqYaivglis/A46CE3qF4TCG+rNaviW94iYGx
1/0ucR7inzYuPQhumVuVYLI47zOLXps7OCKbymzaQNChdvXD+yyZZILZbgYyI/dY
+w0FpuwFGYUEdiaFyFFzWvxu/CgAO4Nh8hEoJqJg2gIbOA3RzekAu+dYbl2didZB
BCHKL4QRoZGP1vlP5r7fVV+sEl8CCIx7cm1dKZqOxIKlvnUmVdV1g8vGqiRNxP66
XnlEKHKsiDIrwMkTz1nzsRSND6qCE75MsM6TjHKoIwDtJ9V0RvZc5nlm3ybp+GBF
jOiRSKmZTIftaA6ad7sZfOVzrlnHr6un703LB0CfuyyyuBfxNSUhM9yd+UNk8AeJ
MIbfvy/wBGxqrv0MLDo0Pk+pg4pdRwCax/XP9u/xZzDiJiXME4hVttRpU2I8YR/9
ov75rw6h13742ltjRGxMBvxZWfq5V4WhcWR/CiXBxPlXyL4/kXP8/SNwG2dEv1tU
VI7CWiloV5jkl13aqPuduFiqY+KqJY3mNgnghwTF12QVoXnqHOHJsuCSQT2uWShk
OhD6jqZwzWw0wex0sKjLyyGOuIine4SL65gfwp/eMWWZnWHsK2Kko6hQEyOq8JhT
E+c/YIcUPiPrW63WmGiZPqiG0JOXY6lbBAY7ujH1w920NpD4DtUjvSE+ls/OP5+Q
SfxliTEJBLHN/JoEj8P3RK2zfRfyR776YjL9wlO6UNE06GYEh9U0Z49JjCShA1SC
1qNSBR8Dg02fklTbsAx3VMrluRNtXVc7aEC6wLIc57YVKeW2snyi84bNq1SdPdm4
ecutwdUnzmFxvAMxCXM7xznyMTzvuYjTXXO4hvp/W+UALDW6jhByHrHMITnf5NNN
BFwcc0zWIY0iTGX8tAH2Gj9RjtzRgWn6DKpp/QoQD2Yg0nKthu48ImkkB5s6yM1f
gBY+ct1pRXngWk0nmJPj5SWmcqjl+Z9ePPhVZxKney8NPDDnHM9X1VhQp6KxVV08
WJ6cW0KB0Iqm3EXXlq0LGThbtKq7c40HkN3bF6VgRENnfzNvC2nnp5jp8a3jMmWy
D38o0jHN71frg2ZKRKxDufNgfpizWTz9bjmy9JJ6SOY6XB/fOAwVAQgAT7tfxHUf
qg07wwb1aiHYdWgrcJZzsLtgkXCS8OC3AX5/IWaXmFs1X43t48GIctpsBKKFeIHr
evtagWDzC9FuXrAZFMhLYlnEwpUP4Hf9MXd0NQOR6Idjgz/K/Oe/+W5X4kVtvU3M
RG3TOqWhFApz9tJ2bYCgtWJG1XnA1wwiuk8kwxI9ygcppoeeDy7hSRBYTYhJEqg1
YTmVgh7s/l9dRSD8p2h9egFC2FH8ZHY3Zk64/z9Et2Gw9HYziuxj8jPDYrIVuyfw
CbBknIMD9U8kgGy/fwmMF5LF3I+mB+RNpCE8Y+b9kPQzYRks9584KFpXyvx+T1G5
VuocGzYG6UiomRcza6NZ3BpOleVzGy2NR3bRFYzbFWhWggWqVlZm7Mb49XnMckgs
gt9aJOw7kaBtWC1bAM6spTAirr0xET8651sK+z96ZiZ+enEuk9uPw0lrMEoAuKQi
f6z+IPbRUOKJABPVeStJ0hKhZetaaWpkM0KlqQGcP1vappMfd0opfvgP3oPgMZrS
pDoo9TJVsSFCG0CDJKxVYrsdfBzFSioYhcH9E6UPzcg4ggeC9L0oo8xt0GBfBdZR
l8NmDaY7S+aSla9qSAn/RYediMYXqPLUoL+w2NK3F16iTQyRVldn6Bd9X9/Rqk59
XaNNYFCjxBQ0wN7jVnmGf1gRHbOeVrCOUQO0cVCiSdxVRITSgoHyEfhb5OtiJpTB
5cvpxA+D3MXRSc2oVyuughQGVIuLuyld5lGVpokHL2kaVXgGx47eWt5cDr8hgBKv
axbY0U7gXR/3GeIo/ONwbS27lrgpLCLuB7TCG0fsBnpX7SMFo+5VGb5IWlnjFPfu
rp/MxYqpeTzE3pTrM+LlCQYfp/xJTUMK3ahczSNJHpuiIhVK6LP6j15lexfan0QY
xfjNWdHnvCUnf/qFq08drfi6CmNNyGaC44ppC5v6qXSRyCisgw8DXL96ULIrh4aP
zUPBAMW76sMzUSPqXFfspVmOJCMGOybi5grVyd68Of33lWwS8BiI9hP0laSGKSj+
iz/7uJJ/j5EU/VycRccikqDr7dxzZgikFgMyqfVygMozOq1t1x5f2YlN9slMhoea
QOFSCqD2YCnCJ8KOlvaVHfLJsjtjW9JQHAFe3DpdnSWXO2/feYvsgIUlfcfoxXXd
fACOqmEbYdB8vt9RXJQP4o1F+ZNyptQIe8eWWV1J24E0ol5voOrCOWQE4LuCCyU+
IlfxSkQhJS+53NbYoV1ae1Ig7C5arIJAVMZA5L3JdkMgpsWVAoihUNONuWjKvlbA
WuKFnGlGaWxLmL1VJtV36fMqr3f7mhcXvVBJ/uPIVcmAu+/KgIqPjU6cC1UkTWv6
7tSSy+ViJXIFDKHgrLnqddPPAfogO2dnpBHpURz1km94BegLL0+8n4jSX27AehvA
pQubcCtlhQtJ2WxYqoOlxMETrTGUxxjNgykL+K/a6JNSohUohz5N71iJ7r4F8/1C
z2bRENYmkwYArSa6k0nYOBe1STv/sjbbetTWcGBDpkNxxh7tk6TxNRZcQ1WIp28z
+i6AaK4fnpEnIgvYFondqjUzl0Rv9Zhz/AVWpZRkuI7wkWXFR3Z+tp+fyzABwrhh
lVRFMYM/bKfllruGbongfjdNLkSsMueHQuWlLjoalBmde8ovGfQVhfOlHjoWTNdg
fovAQWwavqIu6V9LV6qcNxYU4x4eyr2cgpjVLqbn0nVvrjDhZw8BaudKJOgiHuDn
Rbz7UmEL1b41u0BK3YRPak4mVFdeUvTaadecUqiAI5QcgfFhhudBjrexq50MJ3zQ
qylEtKAIkuIBg6MHDrZn4uxFnU0QBYY9YQIV3zetz/4SmqcmlE9yc9hjq5MtrXXr
x6HP4oQ7yoVLMMxgs0KRjBcn57hc+gdIdDbGqcoq6etGfXM0zAH0W40dpaUO8LAV
j5tBJspb8/kZjB2uWBxsIfgnvRg1HwAGMPkn4J3mkYXmGebkO26Uh9DCpSTPPxA6
FEPA4VPGuLyykDk3sneO9mgYXmF8Yg6rrjEqpH/NrNPOOszzWr+sTSqSNUo1sNpw
qnQfI35A/SAr9QSgLH6/TnnpJUqkJfFWO43PF+paHHDggqUIkVlZbuExmg1T6fUa
EF5f9bqgpRZWUgqxwabFi/+nxoDgdgRIN41/EXQ6lGAj6iQA/4PLs2t7O/OW4FuZ
bcX5mteZyII8bTVHJ868WZgS/Shxa4mFo7smp/dnydGuYv7hJSdt0bSjs615I893
k0SXHOmQGyX7YejFVt3J8+gPRtI6kdxg3fTmZ3HXKa7kt0b1nHUcRUzL5FX2Jbfa
Gks1x3cbfr5rWWcJ185w6qBWA2rfPkCPzPQOqEzn/nCsH3CVhfKyHeXHj2bO5k+6
Fzd8vzyIfo47+0HdH32ekQ7SxGIfSWQeUXkDs+mDBJv46KrUQFH43+NeMuNQGDkf
ZAlAEN9KQaH7js7SGwfp8WYMJ4llDby9qlhYFNdJRFWLjwZHEE5s3UoYYFrWgooS
+ZYgudI4OP6Ls3QCGxk9BEwuLNC9cUNw2qoz17YuU9eZKrP+46xFhw0SMR7ldxYe
oCzpsYkYBC6Sq6l99xszP7eJfEA7QIJ8AKe3DopOr8smuA7vtA1YhOTX9asTqKl9
5MO65rcnfx+5O+zU4+jn9i5O1K5JLeXme8P7AV4pH/gDHQxYkzOFtIfdSu3NN8M+
uhQqv64AXGFCkbcFYLo9TUSuvEj11tAtuMjY6PU5DfUDQKvlElMeNUBendOHUxxr
66Ic7rN1b9RYLZLeV0V4uwJqTylb7Am0MIchUQ9oOOOAt53mmDTK2UMfuQV4vnwq
1ZOMeQ9HUet7Uo1kGJQuFQ6B55RijlR7OvRAfPMfXKeC/FDvREr5xVO8Uhe4dONc
+O+1q14LR1Hd7fXZa9Co9zjuQcOnmu3QBA6LFvJq1ulLdTWRwrRHDx10aYHTaluj
wAoDXlDPYKdr2dHq5DiUo+J2UK1MquWw0aKE/xwZOCNx8pgNTqWYcYiU5EDbYEJy
ksMBsJNj7tZNxl9XYs+3j/oGx8Pd+TKxULP2BqguN5j06xFFNcOS8fwE7WunJ/Cp
86oZO7a6n7+BZ7icZDwN0tqJ0X+kaL/PqUdS7SzjkH8EvBWkjOdaDB+90sDLm1wI
A0ozSVVC/8My8Wfaeva+h5aKfnKb/h43njaF4Sx3xeJzylRgk1lipMOH1lXPNw0o
BWsSiv/zGAR0bJDTRNdasVK84nHk6Tl9f7xDSJ4zDanlAC7h/8V7N/ZYqdz/dYKJ
guKpvFK3U/mAbXC3PpT1PlrNR2RT+81UV+bC/4+d+sbQZDXvdUUpefu3NdG1OVN/
FM2RGbBSK+x/7P3WtiuY+5rRPQQJvkpyNd6cL+X62w1P2Mll6Q6ZhxLdSJRpjvcJ
Gcx9PL2+A682gONZujCxALYGpOJLoTb0y/AfJa7cC/z00947YSlBShqQEovIWdsQ
ahLyCf5SPVQ19mJJgelRWExJ/sl7SUfBoalWaIUVqU3i1cavnkwhC5ChURjmJK2c
Y7EkIVNSRPDl0DRRHFjxrZKnyPMrCuLWXyJ+XWo3KGd2dnRuQPyz3JZdrQH6SvtP
IBUY41JNu8URFxYJ4WIJ15pq/yuczRpKdMDPYAX9ouki9TvUXx+XXrdEik7nqDKg
+rHBgtLnHM3PqBheqS8ubVqgKwG0zoju6hVw8uqg5qFaCRcEmuuDQo1Noetl3YoJ
ymeX1tR/VvX1LLh4ZdAiDUp3RxxAUwLlyTHmQHnMrNDzh/i2eSejV3iFnQ1Wxxkt
Wa0+p7jMVnML5wzsic+cBv/lt+XZpoEvBbgGURMLc1TEUXf9YawhtGRpy5/9QVvX
s0BJc+sYEvjxaHkTzKVtuvoLbazgW+BcI3X8ecDbqqjmnCBlX9F6ROWY1EQB2GoA
bCbZyY+7V153sm7/bWcb6vPyipdt3lQxG2hkRsU68iLyh1NmKoGEOoPbtqfTCQv5
cZTKKunkoYA6fl12qEQZt5M8/rHGR7Fa4kXfPEz8DfguIl5qbJlbkRCkPWPEvsth
SE8Nkc5x1IsZ9BAojYp8Rlmp8ebQIzA35uAUxBuPNwRki+WwLavrNP3QrFNs6W+/
GusxQAJOWE5ooxvnxkZChmqtC93aaEecf++MlFUZgn/oCC4GYm8NX7Zrcf9M/s4a
eMyaV/x9ZJvwPAQirMQlgbKu+mA/l0ZvBypPDrwisPr94CTZH9/cnuPDgawTJ0PJ
sG343ai0hcxdCkVRKR3Z3m7K/WLAthnLDKd4nzoRGFb1CYfr8yJFROZ2U+nk2+Sx
NEVui+CPshcPumfNx0qiSxIiNsB44TMKaa/abbs1hTyu5ZF/ICEsqx8Zz6CyZnUh
GfaKMr2wQx3i/Ni0gdl1RVi//UZDHBr2nvNUo1UeuJt/mOCvcmIDiZmtNVQ3wcIg
WhPrg35Qn2FftRee9rXfEBN9oRm6ym4pqGoFrfrvNNa4B8Quz959lsSWCwDgYUWc
UQEicXo7Nem+2N0vCltr5KG2iB5DyRwumuKDoKpAB4rHXWqUZ8BvqiaLCR8SSYwL
5F3YCYr0/HkmFq5kbRJpo4vzeWgkrWn6Umh9gRGRbRU5HkOOEpTUCyHEWYMqNsMB
VcQbG+BiBx2tXPIZS5ovqKaHcpd6SpkG8mLxOMIu+Hk4w7ZjhM2BivrCJca+io0j
QAAuLulpIuw4Ad0laor52qOg4svQbGK2wetGA4C1hgq7u7ZTYLbMmI00y5MQsa8r
IbXs25zJY12iczV3CZd0qmdBH6I8tD9J1HVwxeJANPwF4GTzfaghHP58VDjjC+nb
Wa//Khr5rJLBKrjecpzM/CEXogDZiHmXiE0tdG9LFCR8YHmcosAfhHJ6QajJmQR1
pKgyD/Bl/cHy/1seenaYs/KSTYEfAHqaAUilksV8EyKfPVUBPKl1HLY7BjeKlSWa
6M5tF8YxJ5ptNF0Fgg8FWFOAgULuxCLO6JY5CYX6Aw2C635IkvYtB4ZZHugNvuud
E8p9wsXUXLgBCV6UZZDSdVd7hSqb8P78H9oa+ZwTMvl0rKQbKNNQp2zLaMEuGi9a
WsReGA1UTLEJr+dCo52j5sqlHEvIb+tAdaY7xCkqt22iNVNE1Gr6zRInLzKdEWZE
pXQ6cmTD1OXRTmmkWyBJaa0bdNDBCoM8n5TpdcnkxVvxJ7a1Ow51uoXMOYCAbCCg
InvcFTEDmER5DsGW73AYPXs6Xl4qx2bFRt5tZF8cyWK8f7Q32RnNMW8pUISmu1ph
safQVSKFdflvZFXaaota/1lOTL6vv+lOHeAjlfOrOehSeDG5rAyapXVTaFiLd2Xn
I9Bz6p+A/iyN7vOjELL7EPM+bWXFbaxs+AAX17pr9/NeeHxx5LvPbprZA/pkDXzm
numT1rE9AXtilfqfTMTJadYhW2L3opvDv2Hd7LkDOiwKvvBozxz1vCXa2rBQp8dB
tag2kEeHVOIpUFHa1BtTn3lJGL6kYxhfweWf60yIwcYnGGjSuqyOLXytSrijJlZk
Pt8/jZbiy/b8K8HN+GB0rJacYGI2jjCSi86Ie8oltwJsUfDFtoQYgQseIvC4heVg
V4n5AAMhnAUHc/TL0x2udHC5/UyFg6ztFYRoX9EiNW6L64QGQOADcP/KCbFDdQkT
g8oBZKbBiPfLNZiWpjveDfdY4zDBj8W8hnPMgev2GilwBU/9Y4Fy7K8mFlEgxU2y
he+7xZyxjJpZhtYDScRW576iI4plXs3Su6CC7jXA0C7mSCQmYCWQrcMsXoTeqBKA
3Viyf1ZszKShzkLtRFnBEVsEYpQ+I+2bejDHDZPzYbzHgJsURVpGRcdkvkkBIAxt
HJOGPsLcIjiYaBXqlJMdZrjPowSSfJkENzHdUhSjPb1fsYbthK/tU0iC596HIQPv
rDcbKi9sFhuRMbzhmMWmKTD2Av3D9VXDCnrTvdE1W7Lb/AmCTvvtKI4M++btDMF7
rS+qq71gNWhmpKz06jPgNNQ3eueL67YgP7VAGqw3R+RkSTuUXIAN2ZsxtTH5eMts
pGl0yKOToWD8zpmnwdkE9PsYANucNcRKUqgenL7cwNNR6zIx3UBNHycsNPkILQ75
K8e0/PnB/l8+mXGgibri96qd7DJmxp/DCaeKQxPSVXL6UI0k0qWJWZMkgajRr+46
ek1zTuRfIjRJySTWLPNtENDq3ulLNPgamp12mNwdCTHoMrTkhIl+0JDci32QJ669
cmN1fraYkK+ErDNAlsjuM+FiApCf0toZBlnt9Cqu4gblnzDmDFXdqFFe0kPm3Onk
CNbct+FYluSVRUMIDvuYJUg0Iw6eYnQT4p6LlDiavIoPg13rMyWQ8qrAFpBNiNYA
7X9YN+j47I2enZjuy398M5E84qUqB3Bf32r1WF9FgL95cDt4ewfLyIscAPQnFUnX
211llGLl0J++9iNH0Gwp1YG3tCDWurCDxwJUz16/lTKpLBQJrkjt8WDtGQbhF0LF
1etfu5EzQ0rhnYH7xpwLUC82lZxuZLbPlMeu9X8yyS/4PfkzO5s5WkdJZZfzfebI
5WUmcVGhoVgUjHlBhKocm+fVZw81408vzY1eax5s4ogVeouWVAo803ru9AnLBoqp
ZTgdzZ11bdoxpd6m7ezTbOBBBF/jb+U7CuWXPnpNafBneOb3Isn3zB6YKzPWcfko
zBIYklqVxrdgt4NWeoFG/O7A+TyIMXv7ugHluVYFOoMpQSfLLpwu0WhrB+o3EIfD
6H1In0yrIyNEIEnHvG4sATbabflc2u6pbbUa2GePUu1gHqp7zyOcK8HhWaPkNSvi
2dzevt4LqR2RPy4Jg0qFoMGEMDdWRjOsnJS8DJfHRwiKf1EcVdbuO5cx11uaMGDl
JihRfmVoQ/gEc0nbinqSKrTvQ+vwJfZ68/SC0HZjAMNz0xekGJBLMNvND5ytLglw
wHsUcV8OQjjKfauehKjjZ92+fWU1rgQe0G8M5TuGAq7NdloNdl8az/W/BpzH/aNI
yJdsGWH5/l5+3Ro5R3AO/EH3B0GhntFKEbSYBgOz9QhxyzrsriZWK2cG1OFXmoyA
kMH+9yJESrejsctm7h32SAKNtG3U28tlHn7iZoNQuPzaWir5m6iwAXkdyxSshjd7
OGQrkBCi3AvJ0kwrkvzwa3o1gN34g1lBblxKJvtW+rYXo3e5Q9J20oIEb9lxbEkB
fho33JfLRyvILdWoIRIM8JN3hE44gDKk6eEMcVVXMl3+qFMwiyH3LjpSOvlNNO1O
z4/9Rl5Kh1HmRRgoEudIh//NbPs0DnuTO/WSx5kXUI5RDoidsrsGR/R26FiUCSiD
hYmT+4EdLxBBLUgNO/xAe7Sj+6pXyd0LteMOnDYYwwvtRz1O9PAcvUB5s7BM0m+D
qiCqg9eWViryfSBvxi2Qx0vuEUKEM9IHtN12Dvp4sxZIuI1Li1k5xgDLzk2lHwar
KEk/Le9aPVgF/UzznTDUpjg8Fv2FZCInZK+FG6m8GMCEnw42N3TfXf0RhTzrLxmy
lB2UlMzmQpFnTXo90ueG9Ulq2ePORMklsWX7IN9+MPGeInI5v6jPaTTnktLIUeWv
ivSlbDf0o1Xl91Ml+a7IIZebU/bi1prbNwprcsbmuEjj42TlY6Pz6XVaDYCPgwyK
ywkDqSDKCMcCr8patZpTyJ4O/ethC/4iBQG0f1mdv88wGPa8XwDUoivLxSRcueL/
krf7wCSj6yosz6cPb/hanM2HaCgPb56gnLPAxVhJOv2LmeoQnej8Mfh3J8F5sIqR
Fn5+U1uCc7tQuOfRRr5YyQOa+b8KFgfVnVzwKOUXCFDdN2BL0eh1bzbNb0RiiRrQ
uvCCulfFEfXFzyGUU5xcZdfVWyct45f7xUgLQ/8z0iX1ybtsiLtzTfgREWEcaEnN
59EhAe9U/58uI1HXg1B0Niw9dYAMXw0MWBcWcaW/E+kWUAMg6nxsJps5rJYvS3Rh
J2iM5I7CsHN7BidwdTdlbpmijJpkQuJjfb/iEBNyHsT1FH8dSk80fpVhEUWTtzly
i14RVPO4Ul0AOTQTQf6eQMt6ll/r+lW9WXMUrr7rt6mP1EVjp0MxnMfBtY9ApiGv
q9BUfNfZShCkJeKQL6IxMlqZBpnlgxkpCNlYhTfRet/jMPYs2teffiL+WXAXYlQe
YclWFtNmGhRpQ7N1SHPpMjbYxrw3/kZVvClQLg+iTBfGAd0Bi9SWu6qW7TFPSc+q
8KYXJOm2nyX3FoApuUg+xK3o2fFIcvwtPmy4VgpsP7fe53zP2lU5mNkwi9kYlHWQ
/xboGPhILUFgofqLR7YU8F1UXrsMlHmOy7170zDtCBuHznMg49wspv7Mzdxdl65P
EA2bRW1kDP4ev6VY8vRDzqVYhXehe/MIC/kCpRgnpR9nnxYPIdY5yAqVk/1OTehR
xI9sjFStQmP08GTtwVbOFpltNM0kAice/8KH3O6ry6C4PQfUXOqxrzEo+Pfik4K4
NHPS+my6+7QzsAsaHwlEKzZh9ecS5ufX3MOCHrQw8ZNF+O3nwnHp3/9qytP59q1x
7bHcp+vFlCuyMVckHXQonq7c5wzHoXN/7TpyJdLbeXJhj2fWS3rOvG/QfX+svdH2
wJvxFpZd5aZfp2b3wLoPGedRYL1F1S5oxfV1Ygc4o1olMOMYzadYziyb8fEk7Awu
g3X1kk0mxhDyeyz7j714vtXtJTKqhlErrznbmuJpn5WwjsvlKYxji1kEX5P3hzbS
Jc97kftSX/BixaBVf8aTctCa7XGd3gNaRnXbMJVmciOsOnchI+qMogSNzaKHrENA
srr5JuyeAZAKIVRx62HDL6NXUNUzQpwY87Hzkfs22ZezLojd7wve8YhMmDOhOrUm
IugdKeQXpbRnAiuyiSEpIBz4PfRyW8jK+eMwpL4OXELzqmetJyBx8pdX2TBXXmRu
7K2SlirPj2mfOoFD2K2IZoShwANTptnse9o/0uSC/Gz5GhW9WVZF5AvkzNIJeczC
tLKzoUwTopabzj1+fK22IEG7kwxuPoVASAsGiOtsNlSJZiUI0OyipGNuyeqOj+96
lQc13PSx1uPGK0yJn7bzLO0szeVsiMk8Y2OOmkqdUp1YHaL6foC6R9XBL8/jyXrF
9irDPK9cTjFMnuUJ/86WBmsAHyB8edn3yrJ5hO7B3z0EMiGN+Pkju6adKl5TaSLB
O2Oo1jR+Ctc91CDUTyD6LCZli8Z9KZUXZQ8z/j03LygqSItsWyCrkJe57z6xufHh
fnJNHOOVXBW2+tcb+46IrxDfUIabrloKumsQ/YNABk60nlfCHMI2fP2kSULvhlil
4CrtY5YluHZvLHhztjMwHjuT3u8ZBp0Fg3yG1HTEamyUHuDAeAeDoIC66OcefU5n
INwYLLkk2fIhlIxskDOIApsMY3Mq28em2gh6iK0v04yN942kjn4F9BaCPwmS+weE
TBad5mBejWIxv+qdbczoKwBM+L1HkeUyFFJtDUNh33DMVI8c+8ekCy+FEhCsIvxD
wbuAVWyJrhAFEAf46RalBupApDWgsgVbfo5P48tt/GmLjSvaQeQagtsRRc4pIRKb
QBmqgRO6Msmx4ePsLXh7YvCgFAueItzf77x1f9VehTDHqoOOt0qnmBL6vhTPPFOm
ZU3HcX/wF3HqwYLLthORphL+UteRiN+9pX/cqNZnTseFHvmm0d6ZlX0CMB3Eolky
2+ZhASmkFmEYBC2sb8DNtouE1JTDMvfi1QAU2zSJQm5GuaMtB26oHzJOMyyvoIsv
4U/DYaGgNIFpmB3TUES9Kp20wuBPl+K+sIqMGFSs0u7K+yzG4tTjpVeRxWEOPK/+
cxVEyrTpzXnPONKRV95v/vsVUfU0aLOlXBh6oOIEfI7NuEXsKg6LXLNFjnj1mewl
KEGuamZVTZVZ1CVVJf+7xpdkCEZxFIf6bcHC8/LNzxl38cXJUVguxvi33iIoHcQa
QUrZG2RyNqTIzYGy+XQ+03p0nq6I++FB5E/ObOMC0bl1fx5Z/MQ09fkyJHeSCpQz
u65q9qgWQI25t7t9oNkTfhX/TwHCxfDDm7FvNe/KCTrywUHJXUwow/5SKiJ9GG8T
5i5hV4TW9ggVvHaK/f1+YPqNsj9uMb9EFqJGiTcWdlkdFeBK4glRlLiTteAcxrZM
5bg6RFPrznu9eY3UPBdr9a1ZUiAl2du9vKqd88hAlXnUSb+dSIJiwZiK+sGliPAe
RAGLl8xryPKI75SqmzPkxkVutYeX2Ktoo/JHN6J+ZIbRO7fqrZP3rjYQv0xqKh7n
8d5dvJXu7YDNMY273wVS+LwawfCtIPYHF1G96Z1WgPdaq8w+Y8zzcitFlakJ1lYD
fuCwf29lZxfwZtKvfCgp9tP1hrQCzxDyrY6Twd6vebfQF7R0Kb4iCLj+t9Egkx2/
9FZEAE/m+gBq/Ax+PqlSfFCUiz9xeu8/McTmEvWif2P0U6PbwNM6HgGd0CJhMESJ
wIH90UG0LJ8BwwAeG2++vj63rcLANtUFvS4OLIQ+g08yssadnInI42MSesCEyTBb
oTVMEY6a4HVf1O7OVd+KqQDUOf+u4q/eXQgxYEWE9j9QSO8uUBU+2beILT5BP4XF
sTxBjBFqaYTm4nAH1z9xhOJxTgOb+cJt7GLXmXwHiZcB2vCQRG5jP2TfwtVEhLp+
9X4MpiSil/rkF72KrcS8phTW2OYtzP6k2Ck/oy+rUYJs1a/S6+Mb+zNKAUnZDyGp
k+Sb2CRUTpl63iQI3hthlxY6d1zuJ/uKc0+wJZDl9KupodvChVZjYaoF91+BZitd
hIqO+CmKym6rc3s+IOM575PInHRdass747hrnuFfnMtp4Lq/+nVItaiFDvRaQ9sJ
aCD21vMwQGGb9oFlBjOTe2qH9K9Cc0VtD9qODxFfwbRMy3xHy3dL9d/xxV3IyEV4
bZhjtO1T45ilc5BW//iNRrtYCYO6AwvBSdemdGD+ZI6EK5kSxAunN+pLWn0GRRMd
gKzwMZkYoIMFsa39noSJz8kfHbbL8rQ7+jXAwCD0zxeCXrxBKb1egIYVQA6J5RRc
60ogGZfv48YQxDE1w4BRpMxC96ZI7VvlFujrqsfCvBiV+B9a7h+RIb/Ls00zdSNZ
CSFl99wM18GOY/VaybRf9CY8yLrCXZ7jgTtYKsRcvTy2IbiP4XFlLYSNgjCWF/Ec
WG98y+V1fN9ii2NHNhHhFDDfpFQlr+9bdUG04wi6USkxMQz50Snl87WaYMXx9wYq
z6uxOePDVjTjrsgbDi/VE68jygj1tPQLrCO0/elxVXgvBOIe3tI887WsJ0+7Vixl
+wUMDDKScfgCtmoPLTL9D0tCmcDp/UkzC+npsgL3oCUxSj6mI3ysF6jAIxYwvjsd
/VaP+0j7sojWixgxNvojj/leB6/4hQdlwpYrKASGLC00R24BmOg3gHCCx+B9erEG
5M4d7SWnkB24cnM/olMPtLetY7Rko1R2EB1OTiN9HUFpZ/qHZwys3nqZnHgh8tTh
8h2ASzygyz7DZ0VuHnCf8qS4Q5qh9U+iwM9Ad2EiOBoxpcr6ZOFKhm9Odk4g2TGF
yaFHC8sIpvyMp14p1vPL0sYcHAoWsBNeTPVjUfouwfF5yo9dsL3vbxTKdn8dHA3i
I5KQ5oM5K7+ioaTrQJizzuWDxWOGlUIFP9JrnRMRChIv1h9JpDdM6QkxUZSodeJ/
8Qa8Icjc/ROSLjh2aEdZDiPA/uiQXjKznURByp2VhgvEh/fOwRoa55CE618d3pET
/tX3ENjJRlyxJa+zVw0peuqARLaDaQADTtOGnQnmtHVo30XNp0VAuQdR+TI4g6+h
JRahfOUmpHhsq4WCC9ryKE0nedkcDAqdSKh4eI1AtAmxDWbAkv3lByKe8QIaZt9G
ahOtpaTQXyx9+1M4/NaVH/khEVzA6R3iNotShw+R89RgUmOBzEwbXet59bTEy5+D
hk/Cle4B+XX5cYPnF2QXKVwu3rfE4orK4BhQx+7SYns+55IhRobZdTi8qiFGuGHe
MzdjHA5dEBva1n8jQv5iwgsENHq8sKMI89Nehrym7L1m3F94jTC2EvlUfzycRhco
Vs/Qbwx1g6TOTl2OiCa3q9pQGub536gKuBDhqqRLo6ZHA8ApHnj8BxpMDWO2SumQ
5Fi27RAzCRDWFMNroBGz++8LX/2Uc+IvJOlAO4rfyru2k7NGImPv6I4Z63HnfE7c
MXX5oZ1vnCf1opcoWJV3xOB36il/Ex7fPcNzdZM3Po2YDLFdoCtPEStzHt4KK7Wg
iDQ9eLbE5rNIBEmY2Qh8yGVwfl5+LoM2jXNoNBbkW0VYtSede7cve+ynHNWdXrcx
4aJY2cuaRylOKRqq9AJKX4EJCIgeWj6doRY43brUdbyAyGkORI1ol6uBqaFQVFL8
8VY637gMqpgrPq9IFoM+GTiO4BtkLdj7HOdvVLbXeAOAV+M9/jlZioB0QI22guaS
146vH/fc9ZGeSev17/MYkkKJGqVZdvR6lCMRZPtA2EetYIoH+FTbHQPKBJIl6QWc
F31N725f7NJK/nwsAUz1PAKQR86qdMMlpMUX83U6y6f2o3LpO5nrk3sYXkoIkjl2
qpy1Bh5Kk4ufvDS+T9dPUJjopKzNYYYEkKTF0cEBgQBi/Hm4dBaNGoJFgCB4Kvow
qfUbO3by8Jwrq/mW6TTrskegb7PNZ/tSoaW9iBw4X4UDgxaXctG10kCzAovdormB
C8MLwtOkUo6xj6ilDTdl1EYixViUi+dPb0MDFiYSnKw7zTzZjKPZc7m8hsHW3eoH
jGKrN4kxW0wEK0JH0rq8NVr9wUXrPB1ipe8nngV3IO+OiEOoCB4HZ+YVQcW899Wo
KCFuP7JqyyF9Ixzg8EvkEl9hKgV9QJoL5XQAch1rCpmPG96hmukHM+GdCbuuL2eL
CA1HiH+9o+pgh2jpSs/Gjb6PnhXs9T/K6myOKm3wl89yv2Akcc6hmVvr2u82hCw8
G7+ojuqiQiPS4vfVL/31M8+NjMIM93HAtwBTAOwakXVhnxivrGGhiSjBZCULyNqU
rLs1XmWI/BaOMTk59kjmA94VM6nqyFE4fVb2CYfq7h2quDHvQ7c9oRAxR7N6glTc
HGwQVl9gyeVWrP9lGQXXGmfQYexs2ERMlg/PDlchDxp7QNVb0i1YLDt0Y4OsZdWp
cxGqA5htvcd2gMFnmyrWxs7DU5rA3tYy77+xq1hZdBUbjcdA7MMsVoysVY03MyQP
lRnSk9/U5EZtB14FbmnJPPpUgjN2qjcUebVb/ofd5SLPoYF5UFlKrHQeVG4Ronmt
3213Xo+krArQRURyStFmECf4E8Tp9pqIKa948+08x5SO80hG0GdXVNVdXlm7YUO+
inwDbRguRBvmdH3/esNUUSmxwAOv3e6rlUvoD1d9dX9fgNuhZc0S8HR9A0vqyRg/
AVYqgcEezR+gptitp1l9sNgPV7cKVb6gYY7k5QSNM7BROmQZNm0F4/TPQ1w1bSRX
6YMnbq6VCmiynhY37UbImIhXMQvJ9i2H04pQpN5s49iCf7qCKtB6f+mFhG9PXHUc
RozCPMCXPNolY5qN51EaFsbWvPyUlgP62oiPo0Hbw9NdvRQXjYPpmUM6amgtm2Lc
jjefTLR8QhTzKiVsX1FZl5/8iSv0i73KeKJUqO6HWuzCg6HX+I9+6aw1VNoi/Z4C
4bYeuRRH+NI/wXpHYiBC8tja+dJV479clD29FFIzr+lCtpL2Vpt4Hx0OTCrwAwRw
h0dhWvWjDanvVBxM7vzEucLIDg+0rGH1KvjqZc/nGOAA/PGFzGfmjPvAFY1h757S
Mqcdpxhm14o+bRhnEfUoLVwbpGfhclEbUFcuJb2DA48UAEHYzYlWFtFkoZa13l+g
TLT1cM23FLrrt468o7eNKHF4EGcTq5PDheyaJUSGpWAtemecsYZYnbtOevHEXXe8
/LTYzphdkLObl4r9zgX5K84AVoBMAUj+S/+G74nL51CyKE5spn4xOgOoSmwzF31R
E1svrO371Y16COOxI/qmbqmyXuQVnHS0RKzMF0FGr1Yt3B4NSSrRXddi9O0pxLpF
JPq+GNitGS6IaBpHp3WmDmp6XlTgEIjHr+9ZXUI/Lk8G7++wqA/tdDSm2vouzxfH
Yg5/Mw4qBMf2SRTHxEM23RGEtqfFvarfRfaU3AAW+Ts46YjW5GgBluWsFuFwYF3O
AcdvcF63nOoEpL4+WPwIoFuc2HK2khgkmNGqR+JwhwVpZefTKl0Z46nUMgj0halh
q8dGO+7y85YpwAOjgLQDgNvCuqnwuDeblQDziY4xn9eqMeIVOn/RFZvmT4YYcR1c
1p5SjNUaYHw3nFWfFGZKqh4Z4e/ToDGCBv7l2p5ODhwcUcJwod800yBQPd6+AQj1
4gdUreMF1cI/NZH61wavj5d1dkz7VZwaZTUaXxdhT2vrd5bUO+So1Wl0RJstZUA9
rjts9sbR2OnNHV1J242/NuNAFBTMEL6eDXjpJdpvlqRjQXX+cOLKFqNunGvxLDUZ
Zenx1Plorp7EZxsZDHTAXIK6Hs3+gl5Na996eT/211XuX2SoJ8oxi+FsbxXw10wf
JcUQVxVcNy3p5PpCwsLDUDFAUm05yl21/gm9z0wRhBv7TS6iB0sNT4K4J3Kr2/s6
6AvwaBLEBl/5DBLKqxDniNbi/9cMTmG6ngAILtCB4jteJQ69/urZZWBDeYuB8IJf
/Uk8lcH+kttV8uneRZflCF6ua2pgUxBXMihdyZwdMu71Uw0ElS8sTPaeX7aD7OxF
TyNBZAx8kVuxyee8KQUDcOUJBa1Ko34E/rzHg7gOnSmzDEohnYj7xLZNXWAxCyo/
cFJH0KsgYku1X+RlikknccKBYJHaH7JKQaunr9rdM87et9Pn3wp4n6m+OP9Vxfxq
ebHOEWVdgcEK8gH/xeUM+8VCiKWh5hCg0pB1nDESqqcJ1FKTg9P8Q55KVT89gezT
BOBaMaUuw2ew/A6xLo1PYJ4iECwTy7xb/QdqSEYK8Ow/mYrtK9R1eog2Wpc+OT3v
QI480eD06OB4uUEfRnbjqNYv13vdMpghUY3YTUbt6fjGmhmdUah+r9yzMkdbteT5
lx77X4cz6z0WC1Lmb3GzOR5UM9PHtRoufdZE+3bcy2NK7yvC/nzksq79SUjjUb0a
kxmJebmiV5WulJqubzT359n9dr8Hlm8L5sf7OtU9/fCavok3H/rUj46M15oUbpwS
OhNy+q58c59D+vy3xGe/FwgPPZAlBAm1RmVIU6EYWDHX22kEMrE6RNmG9dtyLmM7
E/RacLxtdMZFYlcBreJi9NWdbd4N8dqCQH7tlA8PZYhnBJl+MIbA7xU4QqF5wBzf
mC6vavZapIRyM+r7hxF+q42mzQk5hGOaosjeMBE6h71NUgmiQzkDxf+DJftXKV8h
jpjJJzAebQ7aJ7JH1lEv3hhudZS9WAcJWrrW4fvn5kWf49p2g3HQUq/Qi9hjr52O
OD8GROtsUcJ3+69cyEXS7mGgSOiP+bLR/8U90XyBVS7Y1hAzb0orGMaeZF6VOKWL
cfFnQtzTKO4eTJOd8EGhOw2Y9EWsnpWz2qcv6CuWs+ZfGN67Wpbyt5AMRtu2jOWQ
ccRnGitqK+yDp9vX13pqhETo+zfjFgbFidItRatXuU8MAm4W0d9/V5dQvYQ5I7Dm
0mDVmji/Lewkh87fN5WA2FAkAflz1TS0/4dJg+kKquoPXx0eoph+ujHPaQRpwQEo
EYbS+bPkJhD5sp1/l/mXATogbqNyQ9r0gh2rHSibBPQM+30DJCJNk71W0Jx2Wl4W
yqlUTs4yPm+1eGMonuCNox1MRYnusUQONqMDeoePKQJxIOJR9ogG8MxKQV0YTJuU
UoSGz01nQ79IgXbwfGfyDm6K82uSL3fNUV7QRG09vhictuJuvEnleOHeJ4P7c3/1
ytjWQgciqK4wNiMjDDuC+BmUnia62Lxvoymqnym06LqjrzhVeP0zocIE2IUD1jEM
Tt8s2N1krbHlvQdHrSwcREWitHdo52MXWL/w6gbvq9cWwvAbNykCca59fJT78zi7
AYKFAub+pPHz+0PD7YWVl5LJrCALPWwVqHJqYWei18kFt/9aDHnlWm5XcBLeoJgs
+QhCtjUTWDDiLCQCjSLZsMQ/SbRpwQMtgiBYnmsX6Hf1BBejBJg+QoO8dxLTDyfA
3SQg0SjwA5//zJClLtZEZQXiCtMbkAwbfln8W94gWVyFi3+0kod9ssGXA1Jmxib4
cVE9Iu/4dPUhBuUOr2ye9qWIIMAskclfMAGDsyXIXNK0nuDy4Y33Wpp9XWw9Kpu7
jquxxlcfaNuCr0tWNTI5Qis5g27ADnNHYrtHdIqQqjGO/tjRD2i72h6Up4cWaOdQ
kVcErhgweEuivuVp5PifUpNUNAiTMLdf7XujePN/ghednaYZhtOGPapLlY8TfnRJ
GhXtfvuq3usBLYjwSqQtCsEi4Iqn0TGP8SYkoJQ91PbcQjGXYV8/V7lzrmO1r+gj
JoN/s0NfR+AH4HifQQJCnWBbej3KgvH8lZlTtTg4t9AV3g47onJTs3l1XElC1usD
USeJm4lKKVqB41Pjt8JktH+XFgEgnyxihqQKgcER5CKWEK8rp4KTHRQxhfum/76C
UMIasHVXYI7diSryoySIPH2PB/CocrOMSz0HqFQPEYYeEGzQPl2rHl7hjp5VtgK7
zQacKWaYj2BSb0f/DDILVi2n9py9nGhI/ULwNd/sBx4wqPYAzEmj/dLE/1epuo4u
YkATRG0UHL1/5SFQQapSVO5YWHm4WKbyAoOkNkD8PxTxbIrKayISXm534arauFIx
UCG6WjQfl4PkPR1PaCCrjeHwUl5GffCnbX7cZTanXGjDxadK84ZwD13ylEX2piQp
Ux9yJEbI8GfIMm7xIJIOHl/AGjVnqr49lTLtjJdltEjPsEwSOLRf/k5tyANNsQZz
AWd0E3w9JDa0kF2MNzmeUuRsESS2XVcmQlkieoFETRSdPKuRBjFz5Rt95GYqI1SV
rsRMNlhhumoQ9T28SnfhHaADxY4b3CBs9G/sbkAI1PtGxlnEXur0xjF4k+VRY9mb
zmMpXDbPSpeja6O4B0uoqMNpCUdQleBLAhL4s2x2aSQjcQd/FN4T4KIaeyUTrjSL
SG91WSz1d1KY3/Nl/VhBEFHyBs2pzBug66aq1/62ypMmQPvt8OtNdIs/V03NYhVo
ui3U2a/SPPhsujBinNhPZLKvuzi1Aul/8BGwI6yOwY1/N8QFtnt21wRmoI2Q+k/b
xxKqEuRvnF+8/8cd6yem9foel1S2a9/y6c7HEXf5UwE6xJ5nqmk+gKwb0pvSgK1V
h8qjifn+9Rtu6mdNdkflHueZTRLZ389uDXbXGZRCDQihDY40LI6/75XZ86JTDG91
BBfwN03hRlgRMOFVHr6xQpGrUz3uVsAeSKjY+9XsO4ppu4xJgbfbwVp4Qouo3qsb
z7fVF+HCyRTFD7gEtqIkUNm90Dc8HjV3bRgMTKnV8ZmsYe3v0EgPjIEx9fveY26N
3hf5lPWJlDn7whtryE6DaN1TQhTmaDsT80VbaOjRd1l5F+/UCHD5GVb1zupK8hzk
JJ+WZCAMi1S+qsm+ed9gdepJW/UZiGrUBMATF6i7kQCybSIT2aaNvseVS+2APHpJ
F96h1WEJfdSaBf+eZvt/XkvfcelgHNSYCdjC1NhK2jyWBKZWeFX5x3VjI3wdh/9b
t1aeXGzDtMBtT9VMCYa2r1dGGLg3nLWZPUrir6PUJ3d3qjVk6KmmXfNuHpf73nKh
bQaQ5vr9sTNRxSzUk01oanMCDpcmVlB2oId+h5EQPJXATopPLF0mM/f7ev1nSg3b
57wfLFzs6JALFcLE8fMfIYZlNSb4Bm9wDEGKQ0lHS9/2lPEVZajaTQLqTtzN3MQQ
bA3zPvKFpgPT/DWNypDRjfAl2pVNowM+HFgRooCoZBp0c2AbH3eFshn8wBl/PJFf
dJ7/R/0FCrz24SzgVr8vJvOs/lTScM3BsWEoTUL93L8/c5EeJpsZfJoVzV6Rm0Gn
yesmq/VqTqVFNEf9quG2Qh1bMoGpxfRAPS+x8LsLqV0tH4PwY2dvx95OJE6+LzfL
GoPK/Eti/b7dtdYJyNVsdGC+m0PuFtE9FYmCOK3ONLrEkenxKQ/OrCnAQWYNmRlt
zmfa1Oeitf3CzljglWScRpspDEa4AY+Tge7t1yNlHsSg9wH6eU3urY6SVfyeMP28
i407UVZ/bpimluaVCqIdNAKw5ExT8ZZaEN5sbw9k0Rtb/fHaHGlIBCjjtWorHzxR
SKcMCMvQFUnG8Jm7HDTB+JGHRfIZCFqHkzT0cH9ZnUoI5Xghmaa4kgvz0lnFExb9
KvQp3iU4bHryb4x1zpDVU8sTBmMEOeNII+DK476zRgdppP1aGKpc8DgAlUM1JwdF
tr+Mfh7Y08c/nn3o/jQI0TtnttYrC6cQFqJlgUeK+QbLI+5X7O3zuAiwVORgKvzP
LOKkgvu2RAc9kFRgVELLmPHsUyuBadsasEYOrCbR6p3VTsk3OoLoRtwDoVMkKtiU
DEJYnAnUXXqz/J+rhkag8bKG2pmrkqJCk2qGoIB1pXRjLx7NbsEu3fydF/HrWwlA
O0mGrzRYIo883+By8yGvMu+7KJBcAGGxW1V1pvGu5JBmB0S81ZmYQXCIkmRnshEG
yE9bm3Vb9dOJBDUkSeWyabUGs23FlW0dyOVyVbIIz4AvtdhmziM90Vk80yFLYciN
gs7abapK7tRvIAylYBvOr7+fZ7UQC4wpWdzfp8YObk6PvGIN0jgnMfdx+ct8qCp9
0bQKtQGe3KXCa9CCc4ijhVfNkfwPUb6YtB1XXVTuUrGKQ9Jx8F2IRLw03i8UO32B
o2rdt85cVugXoWjkaJj7Nirb67SqbNlBsIplCcc+ZGGbGjQYuDrN2bpu30ZR/xsr
2859WZn3OvnKZPMarmWRLw400Q4ZTgWBweoK9InYSbV6VVbcs0SnK6gYHEpKw0ev
oJ9mCZ6M8dDrlkWapxuLeKWwNMXNnFbQyOIGgh6xTTl2XBCkIHCTwzob2ecaj7XZ
2SSCGMx7VfDRBImzc0V1rDWNlIQafTDOq4+CxCr9Z804c1k0oKNzuTwMnJ+QxEEf
2ucd0K6xZdmzJeERDFn0zyfG3NuzrBY0z/p0U8F5tiMstPhvl1RJNrj3e5F6FF8d
/WKZT91eIfZaT/qT2CeidD6MuYp6vjcHa+LoxdvI2/iSZlLxJ53/b62LWBzy1KIN
s/nheeWSekBiqnF6wLkUkJA2hwJQqG/iZlzUXBUadbWH2GvxaM0euaVNk0zliG7d
fUZOef8AfiWr7+P0UjO3T2egNWmYM0278N9lf6Sp9OFwHKFASw8TBVvMFr8Evg2I
f6jJHCn1lcpJWIlej2ybF7Bmlga8GPeuyhFhFwzeQDvyO0rgrk0U2v0HNfcNYv95
Vd8gmpMOGpvV0rQDNpBz+5eufKPv2VuaB18audgXRz3m5TKYSbxunYpukBbM7+j6
RNXC3v/ClgUMu08mQu725UM38kxI4wCOfK13oRI7XrWiQk6uB6KGi3SFgrcejGk8
A7IIhGZmVqkyS7VWv5JLLcqJjfJU2q6SabO9XTpSKat+FV/9v4rlOBg1qmAYhBNu
xb1val8nO9qW6CKZ6tj+Tb3XXZrZ/y8DXVP6m1ejHMnNc/V8yUHUM6rb3rUOu3HZ
42NTbE+ZnDzMX7yp4POm3+fcR3AZ9qmJDnojWnxolDBXKD46rer0iYjAa2wS42Px
TpD+TgBwP9WzCu6jyQCbTtrZMp4U7lCTPDUobTwy1PLsqCn3xH9de9ol7njj9X7b
7SY9nMFXUrldVtu2GgmuMXEdJtZmE2CB+k0gTrW+3h7+03rl/k7oiQmWUDmF3KMi
2FyF47K8x653QfEAC4cuvqFV7LwjrFlZBZiD+RjU/pmJ/DER2mFQGU1oMsBdLjOE
73o0xOF3U+0kxIanHJkHl/aGcLdyY6WS0DsrhVWr9gUJWdm9yiRZq+xNoJkBdITl
TyNjJ5TwzrSfdBOopSe7wz9kkAgTgFv4V8ZJP+Iqv8DB19fptl4gK1g8tVFFVJ1I
K391VtpXXzwCH298CLAM94eI3GhFpNwyzv9b5sTwuYuLljzl8UraIXIG89yCkXdD
sXMcvIvQJv1PkZRc3r/P8QYVPbNxSv//ectAZ4cA7flKANIGXml8L8dZCgjiWk5Q
zC8svzoU/ft1K8BeKeLvwd5OzPFvo1QkaHk0mRxk0CKmofm/Qfu8mDpnobTXHnU8
T5E497MOBGRN9aOMuOHQu1vlweuBGCdyUS2bArcvDIaM5hum+/czZXT4fM2ZXydw
LYhq3EQV8/QQvEmUWf/h/Oli/CsnuGyxMHX0fOb+Z+ALv7b0rDGilsdYJi6Mkkyl
e8tcJE+qq4dhPEXHhs/mZYRr0ozJL8yS+GlwVozqk9Y9v49Ypj876wZn+5c7E7BE
zSAW8b8TAwSB8GVqD7JH2eoTt7RTp2wtzBqIIxJmFHHEzdAqgygMWsqx5kyQVzzD
3hEMlfy7AdreMqR0RzBqYAG1U0kdKNYaEyQ8ttcPFyGfaSUPPwaMXE9kBYNz9dC3
3KWrYqFLkIHyMdzMcQCwxd8gY7D/BFGPIbxFFXoU9l7U2ulznXMszGZrgQ1vY1Xc
90x+gL+57Und1QtcexsLFio5BwNnixRJ3ixbIhOMLQXJpWkItZ9j6caWwWUK29Yv
8yeUH2itCz7wlZk+qmPIEBwuos6dP70aB1F396Jm2EY0fTlnRZr5fbXgMjD/Mak/
elhmallHdYhxPjuSeBuLystEraz4msSw7zAXUAXxBLb1RtmOYsYGEVkUBOKZdtqk
bAS38TBDV6EhmheEeLUhN3Ucs6bxuO70UI+/TNFVKLl45fEHENuy2qtgjIWQDMAO
OeDcZTv6dUhYUWg27Bptshos96b3VWm4t+ksHNOlWtpn9WLKblk85ZuvEGtK2b+U
4OkTlbNGPlNR81aEOtG4SbViq2u4Js949WhiN2lEtcYw6eyv9UPRKfAK9WQjWWq0
ied2iSpU4WwMFfxlPcoroRHJFe0VHC9GXG8IfdGbg8vhap2xcAyiyyin9DMA0WoT
EOetRxBfjJIu7OfK41UFws2kNg2c1NrLCWcdxYr1gn46evYqIuJk7UvraZqsh6Iq
IFux5SF9bjuAiLs+xOSNmDpR5RfgsKrGA8byMDOKdHVJbzKBMPp3s4ZKu52rTP6F
p7sIsigr7026FiPIAeHB2uxmDdVgqMBu+uz1FcNlRkwSwzp5fv/dXVwYCh6TxWUF
yN/VAkTeasmVY+VcaF3ZS9ktpOjMLz5BnD+Brlj1FubJ8zN3WP0dDj1/s69eMfxo
Xa9vP1Ioj9S4hOL6pDlKe/vSQA8QOHTXkoenuzuwKJKYqw8kv9uDxml+tjiCCjlk
uPeGtmgCwRkOnTpV0ZqpybfyBjVsOwg4wZYeeUkhJkWc8e27GjM/i4Ukf0Zt+HXj
XZJToSDLeIQvN6kYVw7oi23BlKQdrJMtxwEW1ZV5/l/IaLwPOQqe2xX9SRMwtT1o
E3BJi5KgAOmzdv7lgCOS7YECfWcV7t8NB69IAx/5kBCmz7VT/ajMXdJBs7Sb2Get
BZB28+myDvhlasT8hxMtyQcx//9NcVI2CU/fj9Mw/61jcrbSQTK59HDE8isH0rDI
PnY0t+GvBIRe7ynOhBk7lsQ2trcKwsk9IwZgrNi31ruesBAXDdgG6p56swqPh3Gq
O2WCWyaUKY134GS/Rl3MeTAt1A4mgTnuh1tHOMbjS375lM7IUe1sb0gtBNVM7p2u
2NY8bWrrAcuz2ApJlpD7BzjBGPWOsb/WdYrO/3wQM3H4rY0xg9mYhz199cGCFC3Y
y2EUhckDvwACuM+1om1NDy8UZMJifcmKWMw3i2VWPEScB0IVoSgZLMg2CByXp5+d
ZGm0WVmHErAPR1/BDJjdl3Kp54sTX4uidKMsGQwl+0iixfZ1BCAfLHU8ULCoEOEz
gHpTsq4RFinZk0QiBnzIBmo8GLi1oeBBcg+Oy4YCto5nZLv8ki2Yo3z8GZbC09Ui
W02jCScR1XswgrVzEvct5x3/k5zIVl5Ny3fneCn6Q7w6vuOJHtZc9su9zuJRmhCH
qI7QIRrfWeR386Le4HhwoatwvKYQdwDunx+CLIW4LpL7v5ogXAbOPZbHe2AW4d/h
dDldbewVuI2xtEy4wHsm7iSF/4XWgKOL0LS3HXFxyzwdby3ueLOEyrjv0ZDtd3rT
qLSP+5uy5N5dBdRnOci3Y7Jlbz45hhExd+U9RthpRRiv4Mq/S8NAEJ/jGcxPbbUz
2DR8f4Enxyf7TzazqNK6p1Xyem6A3vBJ1VpF5P+soXQJGkpIdSi/TSJ8XZ1o3253
R2T48OVlB8Xo0N0+orULTR/yDl+98SOIgtRwkGv2Ruf4dUUYOSOZ0H99SX5cW8Ul
4PscbdUvcZ1YKbHiEIvHDw9QAI9F/+GTqfBijZkR7Xu7wiPJD9HEhwwpGsZdLzTU
iYiSA52wxs1xDo6acuvCyqML8xOtcfbBxm/57HSeBN6v6/OznNA8R8NHSVj+S9lJ
jx0KiYY3RgTr/DbSDOz75GkkdAUNJTLmhfgqpuILxjM2ILiL7q4Wzp7XOIj+mz0m
7LjshU2Oo/n7WgYbUNlJM1Tc8pvI/mIrSdzE21CpPXH4K0cnM1oZW+PIKtM1MN6P
8BaDwe4kDKu4riufH80/RWiWXpoQCHJovV/Nrle28td5gUt/3kXQVh/xTd7gvyTC
1B6fKRc+dw2U/vJi5uKUIACoSy3JGbi1vuRsSS9aPQ/YLA4hXnblJeHYJgJH6kgv
i8sHKOYtNfMwnsALhAPQjDniTkvMwq2KW/zrE1UwM80YtD0r63PAe+SiVTmaEKzA
nV9rVPrADIDyqeLSxcrCx1/o2tNv0VGqSh+SMlZvPbyUv614PV5RkEIFHfXEoFh8
J09LtvwnyWWH9IzWEjtHEB9trAKIzpZ3YwJDFARwxsELVxaj0q7T6f5ffFn8cQ6O
++YM+kpywgR87NhXuSH+418f21lCa2H2aU286hUMDPCo+XgbExjEr5lY4S/JFhT/
zsl44NGQ+86VfdHCPAj8rOKnOblIm3741w7EcRBrU8Plz4p77MoF3Io9eAIKFD/N
XX85A7AhSUi2fz1aAyg3Wqrxwp9faIAZssGA23tHaMtZtlDSX9ZJ4r1FVlmYadvH
YanTlrqFHV3Xuuru22TOshcsQXxmsdkY9UI2IUqEXnlXPOpVaXrzK10RXNumzGh2
uVTYHEeBCoRGD7dFpaQGuKGdq9yLm9pJ8CG2AdqCnfWNsCDQ7lUQbD4iYbrUQZuI
oKzgTpjWqhpDbzws2DiDrwJsGp4XLgr8ZwenXkc4v9MeuZ2LSlkjpUnQ4+OHIuNv
MTcc/xqsoWdEBCxIxL+iM36MWMHRjGZuBitSSGvpM3NqATv/me0sY7snSAQdVMdZ
Wy5IqsAu/0djaMqRGIBf537RiHmt/7COgAHZOc2tV20k9eg789h3XwIcq+nFS6Pm
8SwypzjROj4DWV5R/Yqn00tp03SxE1RnlIClGTiN6eeJobiGSusq26nlbQMB8Pwp
sk8exWsQbxDoLkqg3bUQXwZthjXJ8DmB8DKde8I8JfwG5KolLKabV/y8yO66sD7h
L3PQT90QF7FS6KlrAw6GywC5A2zSVuxPh0Hau/Ideq9jG63CovkgIO+ktE7xlb4l
ncGqivlFw8v7ZaIkrMhffZiZKJ1KthfQwZ7mctMsY2wfSNzXsPvMFdnP8Ix50FMh
5tYH+pgLZ5RWsbwcAQcgfwC94rwCafg+GxXvuSPOntunexsTNUk61ellzhvpCfNo
Q+5QrrWFBCVWEAqrkCFhdNzPsP2sEwdw/bzXE0Uswndm07zztvdPFD7hFaTMp0Qi
ziJWIrFFox4sg8xOxF8AeV9rCS4P35W8nebI0uaQeRvfyjePLRcgfrCzlYLu3Wy0
ouJG3HBcB3bC1oEgAgtmL+Ff5PrwQLT87WfjwhUZe8LxXSJ2W2fXRMiVV7r6lqYw
U8hUY8AeDq0FOhYpbMl7VpD8ckPcN1/XKx7Fr+4N+4+NonrA4O09E3depaUMlRiT
k0uMDp2ngK8GQwHWzzMCMUEFQSXImJFzgbm/53N2cX94Cui9jn4mDPzLkn2uWTIZ
Uc0mNmiyg+IjykdOwMEvNWavuO5tNBy8lruD0V03kZpWJxCF7dShtGimA+DYpjcJ
9N1hJgSZb5Eb++/5r9uZ+AT67Z5k3Jl9xGGMDrJvQfJQDDkj07xtHbW6GHFnQ6Cl
vwyH28XGMN69XzEhl7Sy27lnyY1lvIqOX0eTiYlF+psfiN7eIWYbhc3qTbjFKQqK
DlROrMjIt5CV7TmH1S2l11ODuvHykAHsTc2UCEStYxnfEuhTt7swRtXQC/i+A3tJ
UMR2mpxcAuS/ypb+q/GMHG9AlatMx+kggvaljom4IRFo70EX2r8fV2cS4BFIUtSn
aPBwwXUvpk8YkNJQXHx5AsjjLN1TzlozK1IDRsVFpS+6fI5L7/v2ccsqI++cJW7/
AV1Ng8PavY1v+35avimEw6ewsi0D0P8cC4lrEauwSdXddds+jc9gAgRPjArsYZFo
XMuvX9ZG+Pp4xZOUOcFoJtnxW0NBrGy3o/5QDjl4MboQHU5q5UusKnzREGDypiW7
kQFl9kFRlMiKiUeQ7F8gYAUR4NQHyh91X9e0DVc+0mHNkeTJ+JeCKGp7jkZD4bHM
W8s8QXoskpuT5oCEs8GD0SrLOaj6cu4ZeHK13PhRwQ6uzoN/SnTJISz3UtTksLr/
ZtIuaICRiUXnDbtQbbZjc6NLj8wFleiDtIDlZ43Nirs76wYfsJm6CxjZvt4tk9w+
+7IcedQkhZa1JRgWw6Q08skG9GThwyihDXGDmW6CXxf8uFVnC8QQ0t2+J0fhlPcA
+7YeUvdkgDV9Qv9zMUA/rmwRvbj+nqfacmhRA1xkPHQFKWcljosJFzlfMTsIC+JO
X5sc+G7j5GXMrYQCPIkSwbbd6W+srrkGF5CCvA5wPynkE/prHev6Xp110AMEvn0s
7pQpEih2L+Nxym2h+L5wxahBKvSVtnKsACzt74McDIm6IDW2N21uEkdtNnI+1teP
YiFQMXzfKm9uxmx2/UGTRNrWwFX/qYpwy155ZodxkEBS2skbmgBPSm0JeqpMoJ2B
LQkuUPxr+1hIZyWp0hTibSA6qyrYgNp02dB1ciyt2xkd/6zxUyzeBV2pmd+H15mP
5TuUiteHSp8qFb5K/cONXHl1S14bsqzvyR9OUDAs9dbwuTl7ucA9XM8Opdd8w48R
lAWdm2yt+f+vjlFUb+Ww5hZsiMjo0Q9PbTTT7vP0WQPe8UpWWMlVsOZKnsRrwp8d
1GupBeABpoVbFQ4R7rSqG9N86L6dH5TwB4DcPu0gZ6EaFoHKcdGgich9MsFkrBdV
X+Xqj6DY5ye8zVo9nrvf0BSAgnOpfI9nLfwPnpMTP1gNnh63oDJQ4pBnJ2Xb2a9J
uF4PvZkubWbv6YSq+PuyhPibewekfohgLZ4bAUufGG5a269YYLNuFlLs/XgwH2Qe
RSoVL3RtcEzfmelc5Ktc8Yeg0G5Bz1jxu9Ym04bU/RMHofFGsdsnHZiYDZ4o7T/j
QW1rRuxEnIIw5GnpyVHm9KBJ8MU76+n1z+Wjp0uPnikTI72DMycTbAlTYIcxoCp4
82PgaoLp5FNhp/PhscBFHS0zpS/MMHivyTnJ+0C/ERT6h3nBNOzIKjRN5HsDBTPA
LdqBWPaSsVp7B2znp9rIRr1fyKJh1ece9HlGBb5kjuZRY4a8OZEziyZkfuTYPXDt
mummP9lI+t85xJMA4zcYsbZZNJQzPJEYLQqsEgmBaUD3a1Ri0jUP5FYJXd1Lh6e0
WioSIbmnRQY7+kdGDmpUfzkDCj53ZtwxZ3ntu26J/X3ZL9T4A7mIvOFvzN5qKFyj
wL8D0B1ytSujj1nGw1ps38x5MRd63a8CPf0pox5dbXyl1JqFcVH7l/DmZ43v7v7I
pfoOr4Q4nk5tGX/vK6/0BXgOuyI9O5BjgCSE8HUA4Tp/dPNNs1x/j0E24dFNPna7
XcXxJ+DyctuLsJyaedR9vm/yDJMeAoLNCLhAXP/46XPE4Rq3SJHnyn3JLTXL4bNK
+TCX80So3wwfIpeN2VykYPkWm79gVuXz/dUJu4JHRUDW/vUloShagt6OcfnOD4En
FHgfK0Kcc5IJQnZrG8rrIdiMO9HKosD/5Nvj/zIeB/cNo1eltdGCn6frL9qtpBhO
+8C/pAPr8d1qHSHYSYUku7odNqq7S4tagjCdHqE16JsZAXPp/8NILNhR1B2BDSt6
ESX2R14StmQxSSHRcocesHROj3amvCyolOuuWq/LF4s0jUgUnoEBijJcRqK9NXqj
WpZh/cDI5KN1QW0zJEGot/RGPo8Eh/zKpux00A8DUL2Dh7Vs6rtt6H0dklOvbRup
WINORY8K67iDuCeSyMA16oolZD7pXzfXSS/7l3SguG55zVfQSdXqlWAjRgSQsO4P
kzJP9fE65u8BD7bkDLH64NZaisYgA1qRGDSfqANdysEm1RcOmzIXIdqWo9cYgTar
AlvZ16Mvil7/4kNMwNJmMNkbftI2Oh0svViw3pceMvaXXs4Lct1OoBAmA0AGe7YT
JwKhRtEjQQqq5H2IZdeZRJR863NY4CsLA+lSlvVH994Ll9uS8aD2EclEaQ9P4c7j
quA4q95ukyBBGvN8XGwXabAq/FRgqFtbAaBxpi6UJmsiLTLldwRPABdef0jVfdEm
WAsBqXUT0iYb0HvpcQLl0rmYA0lzJQTIZ1dl559nAJHZYCjMGsk7LQjplWO0wu5R
TyntomQdK8MBPsjvWtZ8t7Q6BtXaGVJvvz2QPazorzm4BZ4gffMpbV2Jv15ahdHT
NwlDeNDYrVHVlQk02XwfvrqXrXZoJGZrn8SVhYIQKp/rl4IPeVu5BjgSSrfbvVT6
3TQ40Mqb1jMwSfZwYqfItiPcV1x/d66kcSvUfMUbCNocLhiKLzAVomypk503nWX9
fYJOY1sidqMAzNt2WfoIszwjZop1Tf6tiq1Nw+197RbxCJ6NH+tlmQTSglFJQHWO
sm7V69r4tLvZz9CVOuEJYscuOBj1SEvo5TqDab+By+zdgJMJu5KmxeWQy8Qlj56l
hqVDKApkECR8MC/rrBL49G/OZCtNWRBrqsvvergb217Z6SUk5wfcpjHVp+0Y/baj
as8Skm0qLtd7xSuUEZgc0L71UDfw8D15X0swhB2DKSfYfOacBIdz9KxvVbtHUTAP
euOc/V8P3YMQO11+A8ESHj9ZI9lBES7thwWVGJ/q+OpaU9bQd6lHUUkvQsUp6hW5
a/ralQ/ec2ueCRosQjOEINKogofA7nQd4jXF1jMpAp14eykiqR5avibhdu3w86PG
mfS989WcLT0cVENmumNIn+LHz8CPo3W6bnPWwZJxSk1WDepjYYpUhqUiFJKplnFf
cp00HArBKeqGK+0qoKs5jDZ4P+wF4IuTWYHBWEaJVH2iwjUnXsPdi0eogiiX+7e8
jyxUH735Kv8yYYsOBGzcQKrmhAA4vR7JU6/1bnVcCeVaubvMgD8XhDdOcOmv1Av3
77Xx0MB6VL1Ix8uGGKasm8q2xMPh0h11T/ogjeQRGqZyvQlN5CcnNReMJcRYpxmG
y99pMVbJmtCiEF6tsTK76X8fU8RnO8TqA2tPfsNtwcOAV/yuT+9X7v2bvKSDo8iy
vF3PzNTobbaui2vMEv38Sd62BHXgyNIHnEuam8nu83jfCXnCkNZ26PMAVNTR8+M0
FEezTXAwNrNGMqTsTM6lJI2eEqbx/bYDp1oxRTIS7PFHpI41q1G7adgFF9CGdTZY
bW1IIjCYvHCbVr+VRl9na0zVMlPbLzcsfg9xbGeJ97wj7Pb1IxMc3VL6+OqeE4Yf
0bjfqzrPURA7M/E51GCuaA1Vcfos5FNeW5O+h7mlk30rGzcmJqitxXj/IpYk9mdE
VAkZKXfncQ0BSH4ZlZQavYq42d+zv40qusq/Pbi0v6+Ayo5LbLfSUcW5xmgYC0vg
MZFOzGKOgIzLnEhExTe1qPfCfSWYB0fkLvF0fZhv4lW7/Fkn2ZaltOVHt3/Lq9xD
XukxwlxIfyNtO1PGHf2P1XJYM/6QXwguFUSTtS+g7O2GBWmlSKJiyZmFWvsrIipf
Xwr8gQJgHTGB7AIbQ6JAaayaPz4eW9xZV3H6ZEd74LrM+1irJr7X1gH48pThUbbB
42ceX75aAzm8PTRl39y1GCgq3F9lqVEzZuSs49noSJW3UCeXxf7Q2udvqKa3LDOn
8r9GzBY8tZ8TYuOpU7WixDydhP2k62dN24iKd5DCWk5PSQwS4BbVgt8rB4OpmWLe
qv7Tycb0Q11crOyZ4/R0ThUzN5bW82HneG3pOECKfbrNKZyKb6at8QoNXV7+skMj
wzkBeIomOcQ0GwxeiK60jZNcMrVQoIYyNBInSz6qzNZnM+s3HCktSQ5rlCrLBmUm
aaMxCH7i+Ay69snmLO1B1o/m32v/cSGN8qyjwyTQnQ/1/AEfUnZpRFcHJ2qHNq0p
ncx+krKMoAx+WMiVd8c6yDpfvKak/0QKQRYP/LhFAaH8KiUArvY7Wbh3tmqk2gaH
hmnjj1GtV/ULjB6W4GvQN0ne+d/9Z2rbjMCue5JIit7tlB8yEJ0qB562NnYlrrxD
Jq008hz/IOoINVrYTl6yI6qLn4Ul6t6x+lG+OTfX61BPdqNWBgdQ2mNj0eRRExkF
UidqXzhQMAPkkmGrnglCNQMfvSuavXf8pXUoJT3jOhJc+SegSqCJIT41BAl+UpP/
PWMYV8/MITwIyF1sbUnOzlf0jnz57PIyrdPuY+qColb4oH27vZ8panAtfDuexih5
F0oFe0LnAeqyJubIOtLNqOffeV7aEenVgSSuCQQdc2FNXqGFze5q2032i8Ivgjjb
wGjm5QPdp6voURShJXrDR7A02xcE3b9U+otpdj7+vFHoKuWSOfphxtXAx6+NkXoG
NgM4O7cpB1vUW0YkCf8wCZCHVPDJQaj1LYiBKGU5k8yQ3ItPwqeBMM5uOoP8pEpp
kuSQmZNrzotjUr6YTbSY7f8DmcEodXOj5wicMgfNfPmAvShg+fwNbimm0zuDiaSJ
EMH7r2DloJcubjFRYiBTQi1ZuXq+aQ/fY1l5X6+uunt3ULYieorqodfTcHMu2edE
Q9+v9yWTujdgz+MU2KEK1PsEqQ1runlCdgmBTftF1+4L0oDVD0yFFYLbeZkgIAmy
mec9inXFuJKgds86tArByyBx6MdndOOc+/jqigg51o4aHCwjQW1VHIxDzMhZoijX
cc/s7p/VDcCx3C6rlbxRNyS1iAetWYNj1skmr7Cn6CkcPOOG1I9Me95Lh/Vm2Hkw
7vO0UtlvQUlPid2F4DynPZwelGZVkPj6nyf3XcGEgUv07BmHE0XokPeWsTQLNEwF
+DdbAsl9558syVUHd42np4DbC3y8fkEY5rraHiUKOtMffiMo5zPKIOTQqJouiRW8
aqq9fNwDF/QKbuCZyZ79AcuSJHfXa3PBzlMyHQqvq7iX6znc2qutZ6O35QRyKjRH
sG5NCE5VzXrfjDMMnXT6kwPxpK5pwi9EVZUsQfDIy+JL/8TWr6XPhrO413spfNHB
xkti7krEUkxPR97y83I7QA/tuiN7m+5lrrOJMZr7X4k4ikcpFTCIHA67OnsIpDir
B2Va6Zvtobvgs4lVzoyZ6vpV7o40RPHEYO4DxqqIdOHQ0TC+T0YDBE7GF2jDuihI
sFKllJDy/xsx2ARRi7xiT78HoYtLqpvTMYxiMxHKGqmxhaBJRR05Gnc5NoOWdOHy
kMuayaSeWiG8BpvaTuZhcC5f1EvxgcDMS9+56izJttVIa8RaYinAJcRLuT9S1ZU5
SddsIykmCMCUXsWmKqmdi2ru2zHnZCGmo903SHtpuozRnlXuIjm9uQjrAU9XecII
G4QtPxKat0JEHIjlAez9Ftmw7w5YQMJa45CckxnSQztHhZlPf6iS6ourqJIJmqUF
cO4qUK+L8iuOmqd69oQhYHy/3+bnswJrFVRAtK236tu9Hwe0SOLHRb6mFasHaUl6
8yncin2EcQ7TMIMvGRD3L/PcHzMRwU557N75MqIXjPR623gjQNMSrWW+BICRW9hI
DbVG/bkQrpQ0GwdfKTaWH5rmizcrE7NPw5ohDyVQWlG1oBhF3rT2RVpdnJdUhbA7
fQKyRKgJkeTTao0t/de4/m7954PlM7SAuIMRc8SezZPosG8tP/EARg/yITP3YV4X
4/f7PwBh4NHc7YCHf5Ij76umAG2mGzE97uxrKUeTtuAi9pMQL8B+kpT5RqQntMtV
vt3+Y+3QtAvkaj+H2EpxLVSsUhNKOXceQpe3jJX7uYor2vl1Lu0W1meRDG+7rJg7
MLX0ZbU2DKr2WSmm24NmQ3sBdHVP15hd9JCNhKeENoTh55t2DbUA4Ju/61Bhj8Fj
Nph1XOe3idjQ0tNwt5twANPvtcOc02wm/psmHlug5Tjys2iKBv+tVeqrk2eOT6gn
ELTFoonEEJ7MMk4RLkPJnw64gh8SdmGUYeBF6qx0dZ4PlaXbHbRdvUqdXrMh0qHH
x4L+tBhcRq6UsrPBTlprZp8BglHaA/E19+2aJ3nvYsBMFWCh0HvDfjx0aDfLC+VH
ywPleJONdAS6TRhRHyr7jBsB/LWItuP4OFqafOxHdkhDqDZSZ2vaeaUUs4P6mINu
+cnfFn85bR3khqQmF2p+Yhw8L1c0kXjxHXhUjdJWD9w1dH90aEPCWiMDJLji845Z
2h/7VOeuRTn0TXRRlNIMgcckP9k36jg97AAaHu4EkDSUEWQFcgLsg+eLMJv8opWl
EeX7HjGEqxLB+Qz2H6MHI5a1t6MhZ3QtRfZlyhwD/ZjbUeuvHF5PG1AFKwInhkKU
dQCYKgeBRmPMwdgSrUyXIs4o41L+h1FeSVnFTcFq6qXqAoeJBU315gfGdJs+QbzP
k4A3wXtPQ5nzecdvNo1Uwu2oBOyc4/Y5fwqznhEVgI5ZwQnxWjpIrvZv7tU1HLuT
Xqy+SgaKaLAiJx4rr34IVK6sVPra3hWbFdmK0Wd2TjvqcyF7K0eTSDS+X1PHWDN7
QjQ7rB0AG8kdmoVu92nNTGZxuJjLI0orS2VAYLACKwlXZXLorhIr7r3+MKCXOm8y
Gna02FcPf0gEWy/gcxkM8QFmfsYEaiUmGrY+RCIOBSQuPeLYsoBmLoknrjBDv0j1
IRrSmIB2rxAIahMFfZzSGrqqzM7woIRaelUlCdcDkIDshPTlqdVvtnl3BxI0fwny
0Kwr2T8pP7H4C1b453Jm9Yl/ed7ACfitH/fx4FfHlwKZLH7qNZb8WJtHyjXlNM0Q
UwjTdAV/BTsXRGgDvISA8dRiE0h8aShybZ+nCj+8IXbnT0/lh2HUTU/2tTMoxpeL
eO9PySp3zNeX/a+QFOnN+1oGwiY3IgTZSGJzbqfNP62uvQJbsbpc3wSXDxV8xz/y
fDNLpaKUlegdajRh5fVitXpnXv8eqlyxRZrv9J8N26rqFqtvDwM9v9nnNI5sdLeg
agoLX9f1VDEGdmVVnwknOtVAusYcIBEbSVbQHkDqIUY+QfFP4EIWI2/xNXTIcXFn
ZUVaNjP0QtAcu8GpBYRU7zIzPmR0j/MwEOeYdXpzGdGuRtnnuXX8gD5luq+Nvy6D
3JqtpeZKlwZFF+1oKcgSZMfbQvFQk1k9kPfHjvfHOY5SAhofDXos24Nlpy/YDylP
afGYVM2WMUPU66Tpx947ueaP/1lOEmKi9UE+z0wlTAKnxXotEhB7bTqb08eBk3gW
Pf8H6OilVBapNxIS50Lwt0ftEf54PR4SKd9I1fV+fzLlgilnaXXxml3mnM2A2xpa
x0z5gEjst/kE3pUCAOevj5uXRpnI5IEq8Tdb1QYXhs4bnkyRaNP/cwzOTGQRLzHx
j7kErjLF+F59xoCs/Hc45oG+tcZAV8euA4GCiiJlPKwvRXhLIS4tRI9sLFX3FGHp
FZKfjGADV6LBGbQjpbExXJCOJCUshXWmYzUMmHKk6mo0ybnaoxZdl/63zynzuBp1
VspYM0Ttl2iSz/mD3FXoGvc9JILAPJyGxQS1APP17y4zTpNPCqva4erPbteMsDhS
oBmTGHTR/Am+UFv35//fpNCwgnA0K58DsmPSescEQnyWHhY4+yFjDlZeBTw/kJ23
iuoUzNU0CfOaSufQ8Fb6FGgQU/GFx4+7D1QiaTCwzTGKgpMLEhvgKMXeC1uHulhp
RDQoYt/JGgmCSmvQqAJnSLFNTT1bVhcwUe1q4W1gpvrDuZX7cfsyZi35GyLKTML/
Kq/1ENww0PB/rze4XJVQtiPKyZPBmQdm9PjltgSPe/V2jtqlPSJtLBWbuMw0FzGH
UAnZ9tuXYRGn3piMSq1td9wd8kDZi+hi9YeqJN4SJESYyHz5WiNR1qfQ9Hs9fbAU
We8wGo/7tVw4mKq/b3oKRr2XxnPTSRHuqFdRPFxSHxiLlinAPo9YJd/+0h4+Bj8I
4oSZMVQbfjC6DmMa6ASx7dWW+QuLyWZMcf/K16gt+86KjLcINikzTVgjowGFLftA
aGsA9Q87Uga2BFg3vXo+3lhFs6Q2Ocr05Ym1H9RDf3tDoSpAS5S8KkNr9vyvwBCJ
PBU25urI7+4As/yfyJTnB3qcKLItwRGu9k7H81uafIajUUZ97jvQysL1i+y1txKI
lnZwca6YcQhw7Tz7fXRCAITNmmF9WvapK7issBGzyh9iQuZoIAKyRjlCSuzUwpBX
zwX26sz1UQfe35IWEAfSyuNs1RpgdACUP2DNW54KBVXPMZeXPSb3q2XxWxiyR1tF
V1U6BgtVHfaXu64oK6PuAutuIngd+7Yot7pyOkL3PDyIfqjAPz1LE8tA6wRbjb4G
Ldj+8tgdvgbYNp8YK8TVGnTF0wTR14+Gx/fsBjNJhz7woQT8kqnEgr/h15lUDlSo
BjuLRIpzuFekdGY6wjZOa4tDgQz/Z5gHFXHUWdU85nUwQTcuTijADFwvNDPJQbhw
nKJxA1CWJ86Nk35m60QpATyrLaVWiEn/Z1ZINanrlC7occCbDmWfGuoVqpeI8AzW
9laiXLf90rIOwDlnmXWkJDFf/JAkVIzLfD2S0CyOXVmaZ4VrbaFePWdYo+576TFy
O40OmvtGWSUxn0HivVXGvXK37vVb/7TtVvsqDfBUJXjJ4QIIusfl27C8pjqOwQ5s
75R2LieOvY8iWVMyAGZEwi+sW1tzZLaPl5S2KgJ1Ted8wlgvMO6orbqItVr0o8HT
pTECJ1Wr/jwPweDmRGfI9xDv79rqjZyypLPVzHQtzia+IzzHBhOd2jwEyj8NDEBb
n3ToVStR01053Ilz8JvWZBn3fmsLsoCOz11t6S2WvpvzHJSUFLMQia0RMwRJvP9G
h4DwpYBHXDzE03HHqYYp5vhBMk/G7rlmb16Z4wIPdPOlUrhHPkTsBjBOC8OjhJPl
x+0LlqTI/fvCFZG7FEmFPVe+DE+iNGBmM/cWbKatnIyUuZA3wT6JtAzsURgzplWp
T9UJpQ4wKhdD1fFxGu0jEjL23Ia/VmnCTOIo8NSKfxnCplCAuEhm1cs2DC7xjAHQ
IBz8mZn8bo48PCsZAiZeVkd8CeTvvqmC6+AZac2JeN735vVkFxrFqLXUNBXS2xrI
VIGBm9GsXJfuxtqfo2magTG4mUlmoeKDWyyv647fT7h5iJUug0mEumxjXZe2zgo3
uC73iPbE3RkzT3vqfsSopbbOReVkEwxjRBJdL6YuozCpOwA7XNksxhdoCveu/Pco
VX3USWlkdzNluNUGjLzquYX+sl9LBrDiZ/kMObfazXyNL/9CqzfjZrTFoT/WdbCo
8NpRU7r3gMA1G8GXqrxj0POvAbj3rIbkExsgSHuU9tPT+CJx3hd20YwR0jMmNr73
laTu+7Gqco79bCy5WEASGW/NSUvinLcwFthJ5brB0IqN7c5UBOpSkstId1/SlOPD
GK5aEep5xUaIEmNxfQEhAX7FqlupgFNVnA2Ys4nn0iTy72MTlrMv31kcT5kUgDL/
HBeerPNFIBQDP9AjCf4kUJBsgOw8y8RSGi5KcJXkJLSWEtI5uAmRy7Cu063Y3EbH
JGO6+2xsrFtBwRhktnYJ0KSCvDQLwCbtKO32SahJLYz0z8na/lMys5KrYSxs/IpB
zPttceJgmZazLeKbCJxjwIzmRGH5lJiLSJh5DFXcihnu2vWvQKonDWPGWuQRDYsA
pmqUfNWpdY8w3PwXD5y4I8pt0rjjnYECfxnV3JvahRBbVXwC7Lr41unZu1xoKGP1
ebXW7AY/sdqt47m9g7N6L2Oy8JmY41/P6gaoPECwsy/KFitUj1G1k2yGxK2BXHw5
8uEo9m27ONloGfO/dn0f9sbORNrE3b4wP6s1S+zIXi4S2b7rS6Rlq0LgA6m1246m
byd6dv24e+2S9mTOPaoyS1dKT0q/L43E7ZJzophyXSiTt/hycfIxmY5aqa6+Lt6Y
BgYupVXNUaLuGYF00ONAn+gzKT/MUD65hCpfGWF7SsMvoWIJk9yHMwZ6a7J0j1J1
IBjZ33npO15wkvGXuh4RBgcM99N3UmGY7y6t7BziJejb/UiXuUJT0PQtUC84eqFS
Rk92KuniC0wlLcqAPVurkeRYtb7ES+IviTqNDqPGRdVPDBuWUvB3EEzGaUZHb4If
MZekQLmBc2Rjc2Yf9Ne5qRnkRDU7PtCLYrA3Blg1gN9VzOVBNfvah88pBLkBwt/5
9Oi0DHDmXIemdLB+W13sHRpk8QYSgpCa9Jeo/LY7gb5AM3eC5kePJH/nR5mUwHwX
Z0scDQ8LhTBjHwSZ5BLWv7pKLZshyoifvSSzeRX+b+LMpiZKd1DOzKUjcuLV75fq
EkrZQyavEndGxBhbCSMeCW/1ejRn2O0PZjw6KFRPbDoyqc+Joledt7SnACCDY24Y
Yk7S+9BD4akGk6X649RoP1vN39XpXzn/FAtMGFocgVwRrJEx3Vhl2b5wkvtZtnwu
9HouaxcQn9qSk7a+v/XmRnNbAvWXi/SRonRONP2Bt8mAQ8r8a8HN24ptVlGCTHHI
ZRBnKK2OsiP+EEoYUSvTTtIrTDrngmGU2dduPgwAH/Cx1dA2f+mkx0BTQaY9+NJY
xUtU5+wppCKrhWDGckTVnLGkeUXfB4mjsPzSJ0cvjpBERarSphPBtPWsiQyIMGHY
QX+w2UfuT/zQ0Pfw8UipHUtLVnrscWlXKaiLv7u/b2m6m2u6ZhgYLFwbSH5dvMut
CZ92NX5SIiq5jpZH6owbAixIitB3oMVbjfRTrK6/q3FyukollKwNzz7zVixUaCD8
mFV2hOZOKAThpTRoEMCi1ggb66lmW24fVZalMqmNsFBJa9Eq282OVW3PMQy2DD1h
Rw4S+CByI/20cHQmG+UE0H6Ew7EKjceEReCm2LPqrQjS+KWbabb1BvgYZCHG10Fz
yJkj1YTRgVU97PW6TRAFbEKYaS0EC30nryc4vR2/bgNy1dWFD/2H2goLL547TOfS
/s9+0kxf8sfI/g89pB1/7Wg+FUj/xo7y3oAiAJJdBtV6CzW8W0xS68kvjRj5VKeA
P4J06UsPexMN+kEMMykKvvg+XadPnM1DNZPPQYOXk5eBf/rRDsZUaai3sy6HMhQ0
07Tb4z5TFAkEnh9k+PygoT2Mm1hNR3fqSJAFm6YVVOVfBjdM1bv8KHCgjxCXhit/
kzYQYvZbamhVMnguuKnAwwVDdwoodx1p3iRGtXxfonjTUrS0tdpCngroqW96dWjT
eoTDzGy7EeffLate4uhmdVW6eJuMUj9RmKFAarGU5QIJVGuZ49aCIi9+HvvTFy2Q
9vlZOJaxHKxZKSZc6wv81ZI5DRQEatWNPtS0thve18ZIrZIswGUxetmgwVHFyX/Q
53+kR+MtSPtojgluNHGFwQq9YSIFOKHeKl81kPmqmMQChan4Fwl2ok5jZqJvEbSg
zfpZfze61d3V6hYmdPGGtaAgaSJWVQSfGNmt7FBE3ndR0JBhbATqsXNOZbxaqJzL
j5SkScg+Mywr5FCTc2lTQMIKOpFvWOiu67m2TgChTFgkuOI+P19XM+mN1AQQR5l0
Y3PNx6ledVARRRh8EWDmHf9lao5vt3CDIlFOZmTC57zb4liu7ipA9oa7fpv7KZf0
yakelKHvkWfZ9NcnQnW6io0gtInNQoamklJ6kC8YlN2EWeLNKyBucdnSeW9YrEze
5mco3zkf25wEt+2cz8EJ9ZRC+2CjGfMumh9ALWPQOj+FAqu/qeGopNNpdXO/3pVe
r+k75pd7TT5HDyNw17aGfN1AvLxSiLRZ3BW0CisKNHbgES6P3vFAWj5FBucr252X
I2v6WepGOF6o/pnm+VRneIklkWxLCr+/4rISFaFObSjhGnrjBqtXbary/TcwjnWm
F/eydJcxLQd3jVy8BMifo4/J2Sgf+lqrODQ+XdCNZQvdP4Bfh7J3UOy/ea1+KusV
E91OGv7zY8enKbIPMqki32znpU5ThzJx/HNk7vnDzPAl+RGLgK6vLSbztyKW0ytE
0O1rcOTF+2wYGNv8+ht/ULZDUGxf4KgHl83RnfSckJXn8U8HCPtZexzM3Cn4//i8
tBpKe/ba8MBhMan8cvQIAWoEGguoSPNwN3Jp31eDgPtUQZrYgwTio8nJEb4DTajn
l7IS6gugXhCeiF+Y/hKOECjVvV2BmiYFnpX//uJrUF62LGe4c3ZCTkSddz8Jj9bS
lumYpaTwjgODq2CdEw7qTnxT8CT3r3+PyiKXemS7PTgct6xnxrg5ZT/T3eEknymS
Vhc2xhmomQ9K/ZEBg7q5ctRR9zdqKDOdbzfcBt3AGss1eNnEie3psZNAqx63IyPf
MUaBw8gcua82FWuqCAVjLZ3mROlQKfjVfjf+OXlIs044AT7zJe2tskDjQPwFzH4I
aBO0Rn8PzZhU8qHSWGtu+25yy96l19XlV4rLfMR8hoX8hbNJqP4EqSoGIzU6stkG
JeO970tcfuvW31/68axXqAXuRomfS66QJl0bRoATQrd6xAbjBTl00eQSOs0jnMLX
sejsh48zeg+CFtRk6JE8sRWDK8zjd0XKBgFeFWQpDAFhmboTA4tmQ8JQL+M05Z40
Jkm8Z5O+V9El0z6fW63gd5l1I+1dC01ZHh9UpVmJVDa72i526DkfADxdp0rOMycm
lmYbg0Ww/Gh4QIEWStCt8J0A+lD6VplIz0PDS2tAlQ14SH/ZR165HOFdK2u8pXpn
kL6Cn/spBdeWMByImGEA/8sBEl5e6vGcWWiI56/KmAKLifT7ZetsHfHgYrT1keqD
PSPEJMRLQz7QNujCIJrk/DGNnNBElaPFCBv7XBlDZIpPC8A2YUR8LOwiVAnSCsP9
X6ip3wANHkwwvuV1NabtmCSZAzHGPv4vorOTrxdWdxaMBnlbHKW8Kmv63BAJS1WQ
84Yo2A63hRmmn9dc39MPRebE9J0pWJHi+zKfX58Gp+0MgWE2yHPi0vRRefZBrayu
k4KTD6AT7DdD01p7N8P7BHWIhmZztvnU824aNKnE8GSNGv/vxGGppuNndRtmNw2y
AWYk9jlhwuT0FJdasFYja4A5f7l7xcPpjVNiu7C4WhiaXD9Ab/eGwa7IHMNavsFh
ZKduTgDT7zjiBeDxXXlYoc7oNNUlb+NnY3LChXWgvE6GZP8uf+shzgqK14es0VPC
bdRYqPBWnStv/01I+NZpnsFP8Kb8ToDFeAlRPY630k7VMEaBlGn4kx9eF9eH6T5c
xGMK6T1tloFKIEin3FPDibzPAFt/EMVCRqK9CVK4k0cWmqeLYwLVFOm5DcVRQuq+
29FxMCu6UufrLTglXnk1ecVbfggHEBIX8ESPCs4tPZIA6yycg0YYt5SQ7e9bAFKo
RSH6cdGrUy5gn15aQPXER8FKD5Nu89DIt+2Sk6Tq5I+0z422rLDj0TJeaoiNieiy
nu7x6+y9f7XTCxD+2knUL5mYrl91xAWwhPsRxWaLmEtsIBHbMeUjAOXkPZt3/ZBl
QgTOO2PCHONYGmvPFkRvwkXM7WhxWwHNltU/xewbrpj4SrRefuOZMuq4OJn/JLUz
8OyCUZ8kyIjUfm1VZAKfVg8FfLU/3yki/Hj25VOwwHkDivmb7EGtQT8abWIK/6L0
Ll5yFAqqfqoEsZ/WFKGj8ANdh6YwMNh64hmYQalPDXoAj0y+LW+OVfAj1TOkzDeL
/0Fmmbi1YCBDRPgpRsRCJU4d5NRnhxg704iO0ZHqmcDzk0QHiDV85nW6i9eQPQWJ
IHyi2/QxpDuDlVNjy1cevPSTCaecpO7Zmpr8enm0DQ1/PYPxam/W2xA05wbBE98K
mWBV0MmxLg7P65E3oUdzdDFEJmgbZBQPcsTwop4AppH7zXPKaljqTu3FPGdYCl78
SGncesFNwXseijMUFP8qQM+67AyE3tkS4EzQrIMkMtINYOgmCzJehgsEEjYx7A56
CLVfaLHLH3EJU5jgqHE1UPu+ytECr7erl4vpkrIXrX8GInKL25w+gjWbu5aq3pE5
eUUliWJcIlKUAjoBUKhCF5AxfJWNEOPewvc58GloxjcSl6+QCZw6p8gTTDrHgsAy
0CYCNi1mOrs+y+mSXYyMwHeEjeuwgW+0RrOPcMofgTFn5ZMFxt7f/NGXRnyqDVwQ
HsDjws1haS8nzvoKO0I19WY/5yfzzT2kkb4XV94jBd4gW56YwgIhJOF3Vn/uMkqO
7Xt+0aAi+8vsdKa53VRs1cQUTQEQq00YdSsEI1GW/8VZeD57EpSdHUwYyThZUIZO
BLxB4RidpoiGFalAeksjWVNY7nQDTHCNSNvaoO//zgZN6CFT+pwjrXGDGu6vUs3b
p3uQ8iDAmGEkvHCX3+h+deLgroPlXzZgs8neub3+aixO+oqkfzhSNydh2xQhrZ7H
ZW2rRjT2C0EQyX8exjJZxsSzjJdWdnHK8SFDRj1GFmGLAYfSLPIsnv406D4/yuMb
UcxfwWcqCHa1s0m4/dPvrrUPn3gwInmHFmnbNG8Uibb1nZIzxOaMT0jrdsg5JzPA
usJxT5sincMOHkmuB44MCIfPaAN7K7N8hsAXp9remEFu/K9h1bes7TnpNK90y1pe
JbZJYl5F2gmsMZv1hgUx/zEPJuDUUgkOFSl11Hji/awOLQrPMSBvnSCUdY5Q43LX
WAgqeiqVzr3PP/PNSS/72LFx/5YC5qfzsvIDfi1Th/WLHgiW1Z9rbjtDcwOVo0ft
TAI2p9FbG7VHS3rTF35Oe7YxGvhvVV4XTMJWqF10Pkdpu+9s+/2+vEAU8893tRwo
ukd8SwsmTuS7C4CF1aChqZ/8XL2HEhO5q8JPKNDQlptxa7cs5o4EN/s9u2J1oHjg
wtgVCd317Za9z46U91P+9Qmqh5TjkQWYQe1BuYH7+fV16EPHgy1GW/XFdLv8KH3L
sZ3TQFdWq3DWZDLxl5H/P7APGye4kU7/gKY2PRXuhPlsfcS46YiEMkY8LhH9d9t/
1tttPoPHO3Gzk6mxYXhgYn3U7i5tFI5leOgX7KKDS1cqeoJ2XHKYDBPJmfR2Z9zg
KzBvSxX4MuIh4dRRoCiF1Jy7nUpVdsB0DpRzQ69qTyz2YjIUjE8S9Ji5X7zRgBss
vEaK4gON2ABsdMeT2zu3BSIOZCZIQbtcgPaotrCwGZV8P+j2xGK+Nx+D9gkhtspi
3Ogn1G2mbhfqqV4EqnL3eIAROzCH+6jlhL2yLkZXbykX9IqAUZ2E4dj0obBCmfiS
c0elGHU7vNuEmatSZV1DQmfnDeTXGPmTbcrBu56kIQjmeUp13mJkwqqemh5aCWN3
jDRocJZsou4biR3dX7Q9TwMdVmXuxJHJ5ZJTex+Yh/fF5eMmuZGzsA17rJBicUgz
IqxEBq/zCzSaU3mIQEz9oNAQbRJwtYmJR0jz7p5UFh/h+v3ZOZimhuUNt22BxeOO
ffy+haXJnImH2GuuOkJ3qORFh+o2+Nxu4wv4Vn2AtH1eEhPmE1GykRq6hWo4oKVy
30wdLBMKmEXTRsK+JdtXjm2xdnJfATnsf/8HQoxmjBPKoVp+iLG4Brm25wlIr7kU
W5el7Q1ABHf26xEB17uW+sNPmaD0+GyoZKryLdNnSOQ+ZpVpLJois8Z7xwUG2fYS
mXsbBMgDwgUHpwuugltUJyPcdMwhvjmMK7HX3Oz0ao32LJOqQquMFw2ChogXGqXl
ORmlyi6tjl94aAzAIozNBkGQ85kHZVolqHBOKEjm1GT1Z0En9+isq1GZdtVg+Tx8
mpeyVZ4IQzIpnmI2qeYdA4dUMZCkrK842w1aefVEiUAp6RguRtb9rhpt93o5IblC
9Gk2Y14jc3PjlgBvF8oKhA801vNjYnHGTDD+KJ0nHzdXv5KPsZoKnPl42Zpq8uFa
fMObiqMBbmtorRBsVQr1TkHn69R/CBH8tG9J/oyRfRFqKl2ZLnigT2daHPjrql8W
g9boVgJsMah4KnRzbe7G1S5iNfHDlLfcURXWMhNYTmKNtvFUqfEhtw2zUMgSATOz
smZd4oWekIEZMMI6CQqUuVHSYb9+0nRLteEnZLlWJCgUKrLObI2DSOweedmdgZhF
QetvmkgfB0eKnNkvlBFR5CusoiX1K2T+v7lDoVGmcYjK7/qimn/pjGMUi4cvKUnr
n4g0C62DPLtR8YOiSEgoxPyFiuoRn6yB6qZBu8KvaTU2D4mlqmP2gf3DcyJbqSYZ
5mB3d3MlpEzPUvNHCbNdI9R5694Tz8f5hcFa+YMDGPViCqRFRiXxbNks15szHiOU
zOCZpGtSe8OjzbQQneLkY+tODmsbyMqcvYEtsMkZ7GICxeziu2Yiz815WFURqbAO
ASZupsHsZ4tZnysvOk8YMhNweQfl4w9eeBQ/dmoyUlQqgv5VuHCgKWRuFP9JcGHk
VTcc26bxMyk54SVvf9Li6Zq1CmLAnG6U1cJaC5A1EjBnv4RikWUsa0x2gDki7lhg
gyjEeo5yaTvM9EpN05mMIuD3PJmtH/BxoM50XS7tzhouQ/q7eGuboEQjz7XVIQDo
uLg6E4VNfH6sHPzj61VW2E1JpZ0kFHln4i3OHoBxUs+52zizi75SPR5iWEK3F428
EjmtiE9LMgdjbJa2shOft3HsPJ7VcR/pyi6LaEiFsTTFr5g19/2GRa4gmRBV6wZM
fx792e8cWFeZATPJCawID7lG6pXH4AkinLt6IFhTJ6V2zTlHvSaRmRkE4WkF8Q03
KU2luTM2nyMqv+J4zO5S23CyN0l0rdFRhSGBy+8z2KWbkDAErZrgJjNi21euGHAC
xv3G8FVs2UHc/iaJaFalcwtneU3olvSmeD+JGnYnZ5g6Uc9Y+21+qpabzGK7p5lx
0rTFd1gmAWJWbVrAuAgZ+5RelufTqp7SDKOIkmu4Srjcq7Dmp71kg7gtOxT1EmoF
3SnaMVrXEmMIr4YuWUkdDQTmZVL8Np2hlLHfnbvAE22WE2SVfTho2CpJGEeP2qxE
4fhKIr2l36F4uZqn4m/Wkix8VW3CyE7Efg3opp2poLpPU9d7MqEb9XSeCyMg+qhM
64i8J2jhDeuMC4mYuwpXI5KR1D40afuM2Lm91szb/uhz5XHYfn+EujjhUVtGmJyC
LcoTByfGK3cb9fIxQ35eYVgbcXEG4+5L2qcLG0dMVkDuxibbKU4YSI56sNF5ZVSA
CuTOP0HUrh9eeKOy8KfSPsJY9l1xCxb+0pBJtCFwYEEYatLZKgHtsC7kksMsL+9k
E1KBVlsR3+Yr7JgIBOH08fgL/DJprFGCafoynrPDREmM/derYNtFN5/telSS7Xr4
ENmrImY2dO390usZ8mgy4+DprVpVHU6daQ6dn3RR1RueNAMHhyqcy5mG/uFdla/i
RV7zMRJi/IW4JPssLZEKh06tZXokDcoH6bB6HZlcbByCuZxrwGBIYkefctLdc2d+
R5DdzfD+RysmAIAu5cor7saDZuxGll06tZ3rUGBGYnosk74uKFulC1gUoWCI51Gc
r0vBONJerHUp5imW4sQdNS6Mj04iPj2FxoMdgczFsY1wOtyYv1Sp2DD/pZ+WgkPG
BOfZcyMhCHheIvO4tjsnsA5F5qZkeuN3S4HYoVLZpkCyxGHSXl+AwBA26hpmf87w
i4BBrpoLqy88bGBsOlHq5hk34qwD4l2ayNMSjsJ1ih+JgPr987k6it8vxpeC84i6
RAvqgzXS6X8itzGzkYqbmObx5zFOQGBL0YbsoRFmK9mkNSXHmXm7B7QXKI04KGVl
vsmHVtvqhR7C52EE4Xihf73+M3aKgdz4SP51h+IfdnhEeqdWpFzD8aF3h8+jxpsv
h//U2YUQaxAIfhqBr98FIk4wrUmeKA1L9MhBidL4XJqcy0s+wwbAqTArD/A8MU37
JvEOCrcIthb+kyqrxVMTfk4fZzuq6QxpR1hb7shu7Mct6jlkG0vCuiNuwqaFEgK7
6xmBUmvnSCfZ3ettoKtnZYOwTy9dCNhdyD9NNcrblwXuz23hM3OB71COmlpKuD+f
C4Hrbq6drD2ZozX/TU8DBW/MMaN1g5iCrN8c0QMDAX6ahniECkLx19OfdOOKfc0r
Vf7l+XHQr0j3dkLKRwhzgounPxQKlfYJDPTHBWIKppfN8gbo6ZyOSut2OrGprj6+
LNVSeGD/+fZfcXoU1LM28+oxXPCxEbFxqFdk1aIatBAXS8bpJC69xyyCg41Vb+LB
xA8P5iBnHe3tAE648meFvR3md6zkVdENOV2a+vtERrNOK3gjzqubSoaZi4artn4F
wh6nqCtoBEgv5wlNNDibnbrHcarV9XvXhRQdYGtp+m/xbDYR7IdS4cWgE/LIGCJO
RI+nQ9KU8aY2ypY/wfCW6h4AVNY4rxMMaHEMvC9FtamplcZbiEApFTit0iq2uF2x
tfeEqt8a+rvRAAGHjL6kC2oMoZl/3qazXm6lT1zITNjUXZO3Hy82RhX4gKe8IEiW
ALbZuEYiBxLZ0yhAqTc4oDMdPx+gU9ge4EekxvCzSYJh5o387N7He/56Lrl7MP6i
EIUhazDkfWyMOoa+Kh0lcOM7AOJNUdXk2FIzKUTpBqfP9V+B4epMUAycAfA8fSLp
AhVwj7aRT3wns85WpEHY0CSuGyt+tUBdGmY/m8WP17cg0WVVYLA/WM054aFtL0C9
tuxH/FRu6kV9lXeQuNI5UJKBfK27rHUH8JhmuRfqtGtFVNKcaglO9kP9SB3DwFho
2iyRsT5DOETkY+DttE69v3WarNCNBLctLjHwKjYnExC/rVD+JOqjjQ9JE6QOwB+m
brG89POf3wztPwvNC1AzPUhJOjTh9wWFiX/RyEOICgASCPrc9EIspLeHaT4Z0xJn
U8B5u0yDuhDwRyVRr56n8OAtvWuye2MS7sAD7lqPDs78PaSlPF/Un/C9KWrmnokd
sb87/tvevzyXdA08bvClAZxM6vmlzKhsim2V05ABAoci3etLyPLskMXnGYB9pmyv
qo8pISFKlmBi7UcAUbEnrMoMYiuGRFwPZCeOZsklfg7G9URCHhro5OSd3EA1MTE0
fi56/ccbHdorGhQ5XwNcjxsuwDUlmC0H4RtuYcO3yPLQncZWRi24jTUtXLlPT9eK
uuhAkxSkZwyoqdMg5v0wIdtkIJ0GuisqeY3Vc/p2MwifE3TiqihBamOJL4EXYFNJ
9gLzx3G+/QZaYRt+pzLiATATjAVvqNLs7UbIhdsMSaNic39IGcJiVeOufEkLtGGS
1fpO9fIs0n/9D9AAmKLvng85xwbL1hMA93J8f4n8/orVd8qxB29+DXzVbP6toP22
mZf1Sti63/cAIofUd1DH3TBK0Cn1Y6259cwR9//Rjpv46EUuDIijgYGX/lHNkjpx
wgRQbe+Yszh0eOWQ9NSwwI9dLBXEnR3iQiygCelVag8w3GXQRgjtT1+5Sd5Kqdc9
eTr3ivzDA52fULm/HU5j8/tqJ/31ymDFTOnR5C9OPIlV3Nxj74OqNOmh6n6Z7D6G
kVcFwbjI23ifFFMjbxAeV4nrb2idDevNjRNrHIVwpb8XStvqeGJ0t3/pTEJ5XtGR
P++PUMxnr6CFzeOVnp0iJrLNIus8nfZV5im3MS5ETSfCfbPaCwLaISwZSxTxDYQ2
oJnw0TQI45DBiKB52+Ms+AYBmXkbmhF8LOQZfI6WeRiIGgZxkYzH3XEKsc1Z2BKM
tOhr0Zi++xAEZAWv9Shq4IL+xMF1YqXwrX6bu+FTFKDcxbpYvol1jGip1vUy27dy
C0KfKMS199M3vbo4uiFgxFK1ON/6nxwL6K3NAAPZd9jMsSd7yDWV+56uzBRmXZJW
yet+qVuo4tGVwQlgkpsIwx6wCDlbqVaziXhC05ZrCz3p7ORgRXBpK24RdUsHZ0Td
9whsS4N6MN0HjDJ1TXV9oX6JMFwl5EJfqxWQecHdb3PCmpkb0ZRc9A9GMp7YhBia
KmxJ/9yFjL69SJaQ3hTkJpqh0B74hgrDTdnjwbu5GLtwAySjylRQeWaRhWSD8cT3
kkwP503ri+dkMPHlhLfms1BLmt9F0QJRhIEVlNLH2WJH4xBsZ8Iw2023/Hc+ezuQ
ZH+0HSFlCWusYjO+xnqlX/uM4XFsaz6O+IZv3jdKn6vIdFst7ePtGRkn8PwLmUNR
6LOpx2rT3yDOFoy5XFsM4poGJfQTurQtoLCMX4Tgo2CjrBPGpgj79Bb3BpMs2FMN
To0WKQkOgXwIwlQ6sDMeabHxUszLw0KrJPDCAn77CZHb0sYiiyobZSxwDdimkmbv
DZaw2sUMzpoMN8fwHqaEwogsQpJejaTPkKoztPtKosUtNYUJMSd/uIms6sxx7YTc
3xHmSiFcsQd7Gkv6SZcxFLEcogAsBhYkbzWb/F2Kl47q6G/K/o1iCxUZWzM89gkK
g1imGNObpZ5BZMM4r3Wi9jTZ5PVJyokwU7MnregfPlKj3FxE/vkL0diWo5Idm4Nf
hD15IK7hT0bkCUC/fR6L4iy8yFK33BeUuwMjBfTgOJ45ltEeaUyMcY3x3iKwmKJF
ETRk9lUEU/Xr5lSrWozaECHtmgUYPIm00qn+Ccj4KUM7EKoj8pqiRbGSlmXUVEgW
u5npEReNgTTLqPUwPMgqM8YVaYrKyeqKjL7FHxp8ah2bWA1K0nxHBDpV/gSwDHI0
qD20bGMtBRYUeLlMRkz8sct4mu2WRXEgrXrl1lIwPjGblOiMFymkEdlOHC5Sn/Sb
wyeBObMThadB3XoKKULsFlOwwAB1S5lIjrWaLotNmlQlamtSnE0YpqD9qVBTmdR0
GWxURBGMYmlvEcqFjbzyiMg/BoCiQcjbaS7xjS84K+AENWqVB/ZKOYSiklAnWZnS
1IyO57Quwv8HY2br0dc+Pz5fG4Z5QZeKWj3RdH7w86OrPCJhEal+vVNYYF2MIiqF
keJIvGp5fHBARJ9ldmIfbzaEGPB4noWDUi+pqe6GfsLqTM+JEfBNpQYEaXrr7cpj
mzuc+RT7chwfdnq3irhkxh8taqJcyn51kn0DdRfozH9Gm7ZXmJM5y2lOBbSTlORb
1lmJYabUpR3zwmXAYbgIhEKLV8aAY2qQsLifkZFxTNz0lOANZk4JdWWhZ3wjgAGG
lpiWtGqo7Y82lbAQNCmi+HW0UKepwOrJZQkxQaK/CxgccPyuBC7Zg6iUi7FegipD
c6tSNADEdaorbGaCJFLMSbcWQfaTJfaNIAa9fim33kJqHdz0TesTit0SbtevbW7w
ajyn4itJgo1Wu28CMZMB5XaAR7GUf/xLXp+EiLXOBYmW+YYhttsjRKlQBscQBK4u
dcN1IXYDttZBK2YoG8AZPp3GX9tBIdpfrXPJqGeZbllKVoxPDksUKEkjJPsMyTje
pVUZRZJxx0ZgXVB2WYSUusfI1T5ZOJL08SS7GKwF0QEBZgGeptHWnF9iIQFhndNl
bNXSgYP+Lg9B27uKOT+wcioBgvIJ0JC7KjQBdmUix9seDYPDZIU7pKN/Xk4j9QHU
5bvlnhaT2xibnD6QLZS3CQF1vNkO5RhBGhZvk9VKKbu5WA8o2C606jtT8qR3m8kU
8yuOEzK7fJsbf8W0kNZYkJk5ZYWfwRMcMG0gR1pP8lp80CMGoV8YTTBdafEGisBr
44dvV4ic0L2++JXWr5qd/uPGz0avR+3/mcAzzpLuSXPdS78TD0mva7eRZZ2dyBKu
xte/85fwia/2A5Jwr0Dh+g/x/YuWJc8VIBjitkXrNzWMD2K1oSX7rn06anmIwzkM
oqIV0ZE0QdZqDSsjqFXWvZbdUhU5YYP1Cy+oXfa0505jW4ZzA6TJfylqyBMrNLf0
IgmOry8MJ0g9As0vwnW6HkBEVa9p81u7M8gMR4Hb4TAqoemKkhCMwbtX5BUKMtCB
e0tPtAZYToPNySvQw4orGsbNWp4CI/NjOwbp1WHgxWAJNzZ7KnWGxkJnry5JpAGc
lnqc34ClKvHfQgbBD7d43KfT8dg8YqqdV+odKYUTD30i04/vWMog7qSR7obR3mN5
tto0QmUONWjPCjZK80F/JlbeF08GgJ0pxVbqkRlyQzrdAg0JhijU+NNfvRThef6l
V86lXVo4a0SAzv+BiTQzPi/T/AIHCr1N37prhlUEH5eAIOoYkRiF2YbuqCSbFRUS
GYrsxVbl4MmErFRcqaYQQJPpnbZmw/CndzKxuRoH5pnXrH1TzKU9agyBBIlpkRK0
K+4jgeMxRrXC0qjINXOS5eVlTNq6l56F9Au0RF9/ytcOV/3MEvetW6/NSKwYjG8t
Iisvw5uo/SP66tqfjp8yZFtAbtPEzpd0ZeDWxyhcrxUYUPhoow+iclyiTynZHVGt
Z/HzNqTC6ehJ5Grqw0Aw9WuQYatGHKrd5+MlIpzXcjyulPmMHyaK7SLMBkAvGqXg
HK8Wk5zVmSufmiZUMzq4VZ8tg/PYwgrhf8h6ij7ntP3228CbDFDVfw9lhLnAweyF
bNHdP5X/XEaLgyPLQs7p7+bcbVyyTCzhfAmWP3AIdQV7aKvp5vTlAxJlANkOg3IZ
x4OPNWgo4MaDBy1Njl4e5RJeGlwV37CrUQGk0jJgdP5yv+H6niXkQJGbWaa+yu83
oyu/Ryr2oNNZ8pitaLYOQgbwBIfW1kYG2LuoIb6s9nwJULOoXQQNNeCHTTc9JXme
ynI2Fw2L/CtqmxOjIgr84Q1ypUCsMpd2Gi38zeJaLEwmBQHnLYpwXJ2NP50kNfE4
2TVvo7sRMpJ7BefQGpWqCBy5GUZZhkKCi2aAKgWLKT953r08x02l4Qayq4007nC4
1KqLsNDSZPf71tf6VByaLK3q5RXqTdXmTigGtvuGWdfXDCm4xG5oM/QBvloTCQWp
/AulDxEkLfvw2sld8gclx+AmjlsvxAWgq9BHT5LUWxgSpxSGi2uTAgfj7PY1dU+a
+eLTPHXrPBqG1TtHKDLfqGzRn7jo2qC0CZdLpYjap8Zhnf4/xET0Sdsw3yvBsiWq
UCVsAeBB/OsydcxkW4RAlJHXWbJt+mf5xidTA70YwilF1A3tTKB8HfHon++V++9l
GjkT1rCEkbAXZOsGo+TDxv3wMVQCMpo5JW2toPopw4LjpsGzDnqcuww158pV25ib
HOhRtSg0QIZY1zHl+GWJQ8mM/cU3k/d/sOUpd4Fkp8aiHK4q2wi41SpEjqMcEjkL
/oXuIsn0OP4aqtJu2qtgmaE9cOcIzEvs3RpIzujVAN8llCK9+a8AB+khAatpDtCi
loWR8bJ3oa0ujFtgBpHRyF+tup/Idm+4InY/uR39k0YjnO4SqDXKrClkWXvC7mRV
Gl+zhRaA+l/CpdKQdOmZO4hAvqGorFJj+fld9vdKo2GSSQ6FuODkrJ45YvIzSVv/
XNGg0DFsTC+nVjJ2E5TW7lzZv/TUwE1W4pSAvxOlhxuVmB74d2VnLDyW2AXz7hIF
OyV9ojtuODVR7uPteYYhpJo1rOKHDgjTTv8lhKz/YAg3Uf0NweY/N+ssBg02I2C9
cNoFddmn3Igudv7Z8suKer2z+DqDg2wvkmgc+cIkEoRcGOzKBE00/6omDIIXmivD
oGw7wmap0ZbP05iuXSldCAWgFOvMDHWYImlfkt7rzi13WhpPtJ+cvnGLwYyEIn1z
b+cz6YOF8K60Xmvb88wN703bCFobGwfoA7Y5I8CalMB2JPO6RIyZh1rgqX8xf+H4
Xy/U8x0ncBHt5bSVGAKx0LhE+eNcCcr7EUw+yaEiofRs1vMNMCoybAtBCXfwxcSh
n5wAh4rFDlDWWgHg9XYThZ3LAPOFW0X4+OFcsxDvlmfkwDhOLrW5N07tMw7lahaC
G6HjCSIqQXaGezUvZTmuZ0hVKPJDMErHcnxmq+DlTsccVbwCvgbfdYrW8CJX02zA
/bQuYyYpVYQ/6tav3j29kKj3nW9mWOaXC5nbKB5/j2mqm9he/QWcLoYNWHR/bpD3
RWiPk+5dmsubqXUwsCY7m+r1Lf3WBOxjLOlsq65BGpmMWylv4ozmw4cAYnPaArRQ
bcE9W1MUbQ8GpfCq6KZbxC5Z7qksZyydwNyVT2UmAD+IDBL0BR2d627AnTnowm4Q
ZPkjS8/Z7rL6Fsm309kOEmuW0+q7tScIVQpYrxuPn4Pm2j3lRhOnw2qCP3bOg4YN
ZOL8KSUaUnu9T0u7C/qcpasp1J5MuupaYwaSd4nQ34f5Mtm9fqrThfiTnkjjrHuO
/T1oqkHOqfMHAFstBh0rkGd7QZ0CdOyIGJUMYtztBps1vjgIm8bbGcsxWR/Rtyr6
+AS0y97qQNjJdU6OmR0pKA8bnpKW74nCldrHoWkhdPU5R/x7bNY8BLninYURDLLK
2R2k1ppaLwJq3vz6Gnu6maasGWeaopDbh42qT7z6W1ccXAx27q6diCQQMR3K2GZR
B37phSvhpr2IswwAMfx8zhpCFdp0qxfjA9E7oRJ1WR+gwSdXnvJHx3yCaP2+Y/Ai
K9ovyGW2Z6vM4xeJF67ZyahIFFGt5UQSvl6ptE50dvFUWRwLVV+WS9n9AZ7MMTET
7I2w2m8JfKnL3h3xSIh8IvMJdKTYDTkAB/07w9GdNMVU/Sl8RVNV6lk/C6ZFUI9F
Bw8SgrSttoJDUvFQENm0pMC7GZXus4lFS3+TRaeAHPCluH7LYmgDRXkOeqpU7dsO
smB8I1huqm50Z0u9Wmn+06myIuXUQE7+L4TXKfJdjI6zMgOR0AbNBZcVxi5N36Ok
gkhInyI2RO7zYrIBIRAA1von8h8CW5ljVyF5eJH22gs//4V/MGqXNrYxGwjhhwSk
lvrKRRBgYxx8MsDtwJWk/5WHeH0kW8zZkXtMH3nhYwqdHszbsfdkllDkzfTKLvFg
KAfVCp5NAJo9Vuu+QpUUB7bxn6DEaGn1sUZSNetI12nINcfAh1TqEBddEkPIxVbR
FQ2Tx8NNM28FguEBpWQe2/PDE7jb9ABoUiybhwlQGvsEiWwdLh3342XSI2z+/9+x
rExW6jtVQeC38hB24y9Sq4XUFvyZjBZouoNJyo/8fsYzdXbD6ipibRfJNcVIxqwu
mPiFGT4x8tamNfV2XjW18R1IF/LadbSA2ikQ5f5mwUt70uSAYw5abonaBaHc8SyQ
cz+Pflwi7EKbOdhWPsSRsQewIPUbOX3Gu3oI8+lOcvq7G/CILyM27tX5omgfNMXU
ey86hfggM6XMBrrhublY9cp9sZbSZesUdorml+gRAqkZ4z4zs7Koi50BTWvMsQ+1
kGJItTPLldD2fHsNBUeDfN/vaUO+HyzolI5ckST7T61CWI5HVlf7OkiG65RvW9fH
GD5TATzu9JNvfpep/+I4xwfWSNR8tnqQ2XNjN5qEyWTwzCTmERYVMxBjN3nzwue8
epL3M3lLoPo57aMl/WJ3j2Vvde1J1DJw5sIMeh0kkAR5c23QcQdGS+HYXZocdIF6
x4opM2S0I4tk91xipV9TCZBbgI2dYk8d1BRZmO9Xp05+LEvI094Magti0CqhMj7e
jotMzBKHqrhVSQlqwCH3csHYASn/s4+gD2IFqQqvCf4VFfbgKzh2TKgvUZyNOoST
GNq9zTPfyX4mGvM/rOt7waZvA+y5Bc9/mxLEFqtb13eyejr6k0jAamGxD6vdwJyD
AY237sHKuoicynQ/I/qaF+djXIx9ORtoXICCvwrplWHQTe7Zf7+dT2beQ+E/4jQm
JrFOheDuDXcP/afwHoGExVFVXCLau0mqPRrT8vq8nC3eSDtiKBVFcHsRzQhzobAH
h7TMjzTAZ4irSVRzuNqjT3oGJw+wN+jV1Opcw9TaaUXE39ui96NlOMd/rraopH6O
plEoSlmeDrFx9odUEu0hIDn1MGK7+8f1Phan+Nk1DOyAnGyBKNqIawkS3ceInkVz
TgNAB7Kcje9uOg54D6HuEObZgRsJWWLKK2PItXybVvG41Xj5QtY1QgPyUwF01gol
XUcK4Ie3jHvMzjeSe8OY9QFDVXmM7FCYJTq+g1gHMi5yGRFsmllZYXUmn0NrhSkz
cB0HxKDm40qyk1oySR9P1amvdG/sv43Lhbyimjou/4WkMnNstSfBjh76DwT3BIi5
Yx5hb3A14Edyn+6WCHMJCO1BNMW5XYdNDfOyQQiZ6NO+jZ9N6qAX6f9sMo3bR/LK
jjjDf/XXuUlmyQJa25UL0XzcmZ/Z076KzdzVp9PCkFi98h/Uc/f6H3DyYiejLep5
qHGUTInAGlxUWUrAbgu9DQQlyjAm/o3wI8cez905XRCx5Kfo+OtLKR9o6q648bOD
0xnDk6o0KxIAjmacIMFytqE9fS+egxVr5xNWf6wTAzqlqlz0v7kQ1b331HnNRnGr
yEqrXiXwP0pW8XzRhGNrHdEVwkrBfIweF3NSvGtcQgikVdA8jVOSeL/z2073Kni/
I+akE0mP2yV1oXBUonaeafer5s5LlHG30W70gVvE4X4yjcpUZWje6SOuPObDrNL9
8iyl6zYN9Pv2MXbf4KOJU8BLRCoiBPJpOEqppLqEqU9uNP5AN2K5sojOa9XTCO/4
r1+sQwjj6Et9HEbzDtprwLtdU9ADRF2zOK6qQB3C+fqQPjhZRtr+CerCc8ckiC6p
wsuC0G727s5m8rdTETBKqA9SVpFpjnIyQTVGojtiU8YJNAKqtQvcLKyASqiwF2WP
HyAjwAbY0cHsJoU4+RdBxn9nkIHFVra7JXlBLzX53Bza7MUeKkmnbHIVqBgDmCox
e/MHT4HI6QkMwI2BST72DLoiH1oyIJXrq06jD5Br6Vgzxv4/lFj9shRyviUZBIrE
YAL5Yy7mlbWP53PeSUU92ho+Pfg3QTR3MZtxUg6GsBqeekMPRoMVtMj9FOof2Wl6
8f/On1xHNbsaRT2OVTuPOOeEl3xSo8pQxytmkYok/FgkD60Dj3olpH7cUs9p7mod
RbTiiiS2OFL1MHCDPscC2AOMVYcbVP6mrXQW6ulfwKQhUhuoqViZkV7GaooP7b+1
xILwMSkxQesRYUJszHj7kqcn9uszpS6ZVtpVzmdHr5pAh0VQM6vAKbF1BwvOlRH3
aNjGqK4upFnrSG8J/LDV7yCpMf8vMUasmtmbulxJMbCLW03yKn35hemhISrrzrHu
5a4LUSkEFq9D7VNXeqt6slvlHTgTke8Velh7VaFBLIzn9awE/kR0+VBAPYSL7gZx
NbtOmkXoXh6LYvAQ5b+BNByfgD2IkqxSXYiBTjFftPoUquJ+kbc12p3c1LtQYIu4
tF1KHTyySsN9EwS9DtU8rVKjeoUctO6FDVIiYYGGmW5Gi6sIJnPN7qPSBp4j8la5
iNnL0Z4DsajBZq1zRChFA4HZkhH0qRYCgi9uKx2jlaemDgA8Lmsy1vr2un9ukH86
1XrIVCtHOcFExLxrNb3ilq/V0/xHTU+Y6Ljq1li9QXchl+PRN5q2WXyRlviZ7VS/
ZpegqHZiV6qi4gzx4PrZCd7JR5h0xGOGK13lKEuJkTBPZdxy2h2AmvGScgsOkN08
5MwMQvkybkh6IvnYPM3MJB17g/cyjzgI5N1eoN7xsNIdey4chB2h+7WzjyRi/5mA
XEa+/kbFlAmKEJaDqYySs6gqDjZdiOkkqKgW13xfYMuX88FLvu08m8f+js66WyTk
KgierwzDndUpV2SN4vTXr7BeBhE4YOPYEGf74PNNh1q3hl4wK66EfI8dKfOtY1Ci
/ZsWv3T5/WnE6C4ju9W5rpdmg9lKD0+GkBvNdXuCJh4kzjDhVZS53XNSD7w4UME5
ESlKFTr0qva565EHakXjGd5S+LTAZgry3XVLqX5G9+GHBk21Ys51VTS2Sk5wG9Ap
IvaRAyLX2NGHbeGzHkPK9lw4T6F2EcuGSszFmwnmNfJUt2Sa+Di/hejYSo1Qd5uG
4rCVNgRbm1/cu7FEgrjalMEYqLzoATU/xnEcsFZci09Hrin0H7+GPOarvSPP+ujH
aSauCdq6vHZmYe285NB200E/FExbGw8/XlV8nNjxdU3iNLPEqoIOe098IaqWPCP1
hSqmjhzhUKU0cd3165bbty3IY4J3ntNrkA2Q8Wl8uyp51hxxsiTRVLL5xgeQm2N/
bI2+PXeUhhAdf/3gPnngGNDoVb8xja4zg5zMLgJlRP8n8O0vUucqo1VHGiWwD54J
TWoC2mlFN8yUJZ6FpM+/9QwIH43mVfQCWba14EO2oBF99CTZBRka7BQaI3tMjgkg
X1rNnbyuvJk+MloN+zzJ9a92k8g3ay7uAvn9X9i4P6KQKuFU2kWoQK/mDfys22fg
HtRdtd0CkAzzcmXlm7ANC5saePP7PXHiJzCdDsPmzYzioV6ggxdez47cD5xMnQMJ
4EFjqx853yWcnTLgE7VHFm5XBzyvRVnXSSiv77SYjtcrJZ/QY8rTJYjXSQLXIe+L
uft1aVZmmkP9sBhEvyQYwuoLrjSYiX7R1NCUDz5XdLwrwmSToBKhGcZDBEMbpiXW
8OhClMQ+EBmY4CckRJy555FvMKDGhoTrGkxi8n2hta2IrDtDdohuvaVRFucHWMYR
tG0C6a+oogqZEJgxaiBOUpLe0ZQQJeaJk86pfQV2N93kCua4/pjGjexrKpgR+Huz
3z9eM2j6evjjPez6GbZs/4KLlaQ2STO+5QCu+S4+Re/zRP+ZUDg2b7YeZpgTWUQo
sWwA8XDSfd21EcaDtZHyadCLnoBqApnzQX+v1T2wdp7rXybPvnR3ZpbWpRIOo5Tb
YkQNKDiebWtr5zvHYmjyfJ2WBS4tNFPNx9M/LMy6FW2YCsVbJiHcErMpo60cmXxW
lD26FxrTe18DvmL+DBE72xAY3vwZt4ynvpU7WwiJAqtoQOVreGp+N1pNZjqNk4Je
+zcQ1spUY+pBkgM5lzTfm2OaRobR2eK+N98ejlYJl9wUy20KJpr1m6pDUoO/3zOP
OyRUdgasiMqYw61+lt9JfQyOFmhT1XBBgQzICkcnW39w7Ujdb6qTjjHaLHj5qw32
f1HYQKVxbjrU8oWfm+T3XO5u7RtwxrEIsPwgDi8BF3CYWgunjeg/v8zg0IXo356w
oTr8GQGw2LSc6pAVqS4ljTlivymAi8G4iFPfAtT68OWjOBpa1wTERB6MXSxViy6h
HIici5t2iZSn23s3nfAR2ifSeT+Dvh9wkExaspyMcwySH01u72FHeHF4ID12WNPR
9gwaX+qm9uPULj/QsvCJ7mGT/Xg2vWL+FsBYMEaZaUX1BNEKK9c5PEzag5LwS9Ee
RPZRjrzGmdhU4wqS6EQjxY3LDHJXywzIFapqgrWuu48mdP6iP1LR41oRxWCmm8nS
UVCLloIXV+kxD7TPbSuRuvwJixHjpu3IVg0g+lgfGBGNyndzjOQQfclSXF1Hmrv/
i3LrIG1G+zOaN/Efvcy+cyOAe/OQmxDf6iYyFFmS+jw7F/DBzv5xbVyp7S3H8AR0
xoO0SKEMiKt0Tc1HmAwz0AJHcdu4v2mVk/uIwg4mKjTnaMpoF0wzTxPzsz4wf2zs
wMJhhu8ZsQa6cUtJv7G2BtNQN/FveSYhw8rAszNBrxX9A0yYGxnkJFcOTVO77bpx
KJOntSACTw8mU6bcsS/WAe8K+AfR8diasokalmw9UbsN8AtNNjRwOx99lsiJ81GX
4O4vs0JwkxnpSBOksdFGzS3UV/GbjvXvWWk2bWDtem9Jq3RlVseTQ0A5ozqmO+4Y
JELIURvxS2eDaJv9i4WV6T/SQNSN7ksdBhF7pPEZe/IwcjZoHssvCdnJJpYAQOv4
T3a0obUjGOKn+K7ht4BH/MIxSyMeGlLhzPw5SgGRdRgsFmfVoeQ4EOZUSKhev5DZ
uqH4ertsQCElWycIYk4YzBxEkp/tYZuuJEWjx8eH9rV1atYrYpGSViQr5NOQ5hh7
pJUI1qpgDR9fHi3r21zrxFGfP4SfKJb5NdU1yeWz0+ziVXSvG2vWYESvTapDs4wS
b2vKit5iPNqBcvaGwbFelVZlA8T6ikJ6j0+ALixzCJRoQqUGgJrwVF3kVmc77jWE
UyG2tm09Lz/K0o0c3iQiwTosbDRRiJhDasYnb5WgwugCJrbuRnaqPWwCPzr+mHT6
YwuoAHVVsVdA/h71XWVXZowItM23wrKGcwZkr5lN/YeENNluFD30ODGMXXWT6Tsu
Be3Gtu89bvFN9QL6QHSCvTXmf3yGz3WGeP4NRfzlgbgfgGW75ZJi7EYVet0iyKc8
5t2m026IHWsYHuyfAVnEaxPRz5u+zNIIqcASSbZxspjqD8kugv3is8Ztvp+dKYDu
rv/7FVVLdk1qALiygTF8HIKt+tKw4XYeJfsOzhOaLPRE6ftf+/ZV9Hiu9gLr1l0y
R9qDZfVtz8FqaQbge3hJFPUt3NwP/yF8F0pIhCyyBWdOWbVPl2oqVuQzi8ssNcol
X+5qmv6oHeFJXZEgtIJ47q1GgMhvcx6bxYilvAf6ZszYG+MTlP7Uh4iJMgrkBGmU
DC66SDMfapA7KM3KMW5CoHqngX3sfh5A4PTWJqeFl+d7JNHrp6gqa00p3ncwGcN3
v/HnPAn0U9pB0526s1T0j2n3VCQBiZ9FQmYrqNhGfykoG7Gx+y0KsMJeO57sS4ZS
uHIwwIUuWZloghwKjHYHI0jLQ6zfmGkHA+qzmM+ePMV/9YINDJkxfXC41dJea+r4
9Od2UrjY4GdEw6j4ymLGjQBTa7Ut81ra3CnMNSbhQedNQw0KaHEuezE5tamC6T/m
SI6Mv8vEhPirGnMDQZ2ErEOOpSqfA3CvS6g+zZJXeHjClHeBnr11eHsru3KTclfV
wv7Tqkvpx+yPKgHTUGRBK02wFZAptnVyinFIVSIow6G38hlOyCcdTtRrO1LNided
fqzMwSc6xotu+7oEz5oekhtmjrcxBDUTy9tdpJnVKmbeytbkNjGs85iuEL80IRbA
igxfgObLM4s0HyZnFAbGNIotzUWVJ4o2UuC1iDcsJ7Xbuw+cAu4C9tKXifz+eUqu
QLC8PWGn79O/SjC1D4OFUVfMaks9p5on4eOGhY0xQhvt7qNRUAxA/k0joOq/y6yb
UsvfeODsHwhRM1Sq97sKhz0ou2k7lL0S1g7n7qfd7KmePtR/QGdVSkYvUJv72Dsp
5uJJvhxmA2OWvFoeynCP5nZd+PAxEM8U7KxDqHKTkbIxy1N1sqGNLG9tSgCpttsL
yGRWODZW+kFsWmPin3d2WaA0PxBdKx5MUYbmxfXJy9wXYycWPzKKfjGW1OpThVSQ
WjrfBGMN1c+rfV59yZBm+gFOy6j+SHlqtsX1pTXe/PqUeyg+HIzxSAUAeiZM+g+L
v/iu2rtVSCxH4HF9fpoUWnon5dH5gXdKvEIIoKyd4qdU7kxjH4OPbf1rS2pbIjZX
Tr3b05kis2PNJc6336HTjJssHOQpBqis/sJX/TC6QdPAkAMbU1gu2Y3moyvQgqlj
3/c7HUVWbN1+MzAs+X+SC0IgAleqYwSP86bSxSQU+OQXkta3sef9VrG5lAFKu374
Oq+fn185DvRDrqh1Obdt2TLZTdXBwJQf45iwTf2GpE9JQadx37NaGO49gM7WPnAw
yDJSzR46Hd5tMj8o39pxqP8h8ft9HgWieEBhdy7dippFLpqMoZWmCgAcwRegRzp5
+U0n4W1/UpRntuRzwz2r9I71o6+sOfz+UJX6w7napHwNJbsjIzUbJfiY9et+mMRl
r0Rfwh9yiMSCvA16RFxHJ1VJ/zx5wgGoQZBavEKshbv1u1mw3sqnFeH7Kof/3V0n
FwccU/z0NN+GeJeKtwAz5Mvjqe5WFRY1pHmlvz9DZEm6ueS4bNgo7zYQswWdQbim
SbxHKNPiAhtD1AAPbcXlGGhfgQC0MTDNabpDWR1RxjmqI5TaswsMG7DosIsO+4nH
7GfOO1x+MGJKWEUqE58hQMujw34bH4pObh1IfpDmjSQbXmKcM5Q4Z96NrSohe7mo
EDb9DAuzNteT018YrFl/2hwtJ9SwotBfBJjH/UP68i3ILq55tdf3jfrSQQTNpVL+
f6LTuKelrO6Jgt0X1vdRycWt3yFfGd3jS12fuLv+Y//CVpiq5eU0sL/vcLQNZsXh
2vHJi9eMF1UvKEEajZi/mjgqxHw0YOvzOxGz9oB4Qm2TxQrdFFvbObZFBnYiQRNw
myEQ+EM6YquD88WxDQsu5eHE8cBvZRnSa6xwp2tyms0L2cWWlBgyZcuRjFsSwxJ0
4huCxiQbnjydoDIMPDurUFdyFcaRyPlI2XjwMp+ZFHZzeHBvij/Y3H+Dc+CfsWAU
g0jgpHkaf1Kn8Scvov9O1BbJY04049hBPYxptdmaKGCVLDOYvrmsGJS6TFWU5ZlM
2XPS1rJTEyjjYmQCc8hOPW0bYnz/SMOG1mle+UZ7scVUbE2PQBUDHG3X11sFdmmQ
pIYK6GQhzHbaS3yfiflmpZpsSx8OVOQFDyZB8uxKAx0cPFMYUfWK6F8sTsyfATwU
lGdT5jgasOf7CY3CL8Lo6R2FNxGLht0AKknuVWadEYJtlRMYza6rNgSRYi84ITfo
MBFGrg8ua0/7SHY+BKypuGlIlpw+67OxJQCUyCBNrolwVIkRJz2lOov1M7b0mW3i
6r0omd0fwSoobTyTw0tF+5mDjCEaVtPWl0kGtkzjkzYwd4PMzs2gajNaLlaRgcze
gDZiNqMLQVxblPK+kZS3gUyFpvN+Ed0uqWdbn5jB7biGvWFE0Js5/2700gJFFqgT
cU/HiTKCK3pTZM7GL3zPJBxPTaafkaxXydVirF5tyNprICiY3NUMaoupGpkXysf2
6g7xEBPiPCquhdKYbI2uSdqQl8LcOvoBKo73IMznfZ2WXdNwBSURF27H2zCbZNjr
L866Jyd6hWHU5E6/WSLX5zVX9LmkEkG8icJ1H4eCm2YXG8dr9h8NZIIcjlHLqWqT
C6Y68P+nr+aSI5jHDeZwFNxdv4VrtuXP2LqfuiGOBtw4fYQvXnF+UuxOK82kB1w7
jH1F601W6LIHkUi2Vc5FmUzNvSdDRmaRn4VOAn3CI4hrp9ChICT7qH18nopY6IVq
pYJNgnhVAo3x0rko/TDHTkWa7zzIboqk1wPlWeaAgEhWHhrSWVOft2fHnWoSBAlE
avYP/rhyMp+yfVT6H6tZaQMnS9yHQnQLquqMP7lZWBINWVVaErCWO+PHpOqqJvow
Q9x0aC37rQBqICY8wTgJr8jn4daI8nklVtm/NAUjGIokDANgyYvv4z12UbXSJkZb
ssWE6nwyccOR/i+9Vn3kSUoBqr/q2LeCf/wQRRh6y6buVtx4R95SzKP1hqoBrqRx
FFMhyW1yDVeX2jnVcWHeb6d/aRITkrc4mdbtnqeU29WToalZJ4Yj4+TOnegCE/Jp
8xKCmwswHtqIqG+CMGQuAyee4lyxrfnrbIAd6Vc5hrHir77Tc6+10cuOZq+5ORrA
Lj/TlcCJ8q9JPGvorW5Ait7lYnS56guPbthwaRxmI7DkOTCucj2c8Z/teObOcU2z
6Hij2hPz2x6TawI+bQL0oCEfcZ23HU6Qg/3WnxkXG5nOT3B/+OCF3RC5KNNev+V+
YX8aLS5OwgtiPJikmyAE+WOHcSURCAy7q7Cw2bHqcH8iAKbbvoWBA/mzvmyYIBMs
EoK9dzV7FZ0PbtzMZjA8UY86IM8sTSq48dmOy0Y3FGGVM9xipeplzb4TshEQu/M+
T8S8lo/pusABUIou5tSeyr/aFHzob6aBfQgZa7gKqj+E+ucHf+lW9eP9WbF/BcJ8
Gph63lk+X/UNx17GqmmPNeQ0tCJZSQO64iiR5pb8DDgH0/fvLu980LFKD7hA3UQp
BbJNhu7n03sBKJH2yLr/h6Ev2QlfMDdGoFwd4RpRSbQTugAkTnDUd0enbQMnm11M
Uh/myTirbmsNdBTiqdNCVTRUxlRdZgd8JP7wnuq+Qj6Ho6CqcNoZ3S0wiDNTuD7i
WUuYQyYpHqUFDk5ocDSNMm8PX7EJa0L7ENLq60w6lgo4W2bnNA7TX67PC+joUuAW
Bl03V6n0tSPSPnbYBDXgW9t3faX8Cv/hTu8xPzKurh8/b0NmXqprDhwidHQCo28q
C0q8DoFjlnPnoUlAUZeTuCTkVPEIrG9udqxW1Ggi2G/n2nkJc/EzCKu7JlWpEHH9
JYQRQrsd+72tFRjXXsa6KdJ6lDOjgAfpHgAnRbu+GYTmWldVEEyDcUM7XTvIfGg2
OBLgZTZei+pIy6BGmS+BlpbC5bo+i5pxe+UH2S+08sXsGyogxtUbq9KfBkFzzOdD
SBC4ADC2PwBhoSfdIYGmIolrO84yGtS7xsHxo6EOUIQ0+NtHT998HwicY+DpkIxr
tfujy4Rcvk1d4kqIBIHd44utBioEjFa877BG3w+91WZxOEmJuGsWNT5cOfRxKBgZ
+JWy3rx+yv80lwxONU/D5Apxc9WrUNOdKKGoEud/KyitHE3q06i6Adz1GZ6fhIOt
SM8sOQ7McOUTQJyHD7fvGccxLcgQIyj7BcZrrLj4NIGA9wz110KJPt+rrkOCI2Ks
nQeeVM5GbdBeJwQR0So4dM2oIJ2j/Cc1NEJYwFwMrfruZlYPQgTiN3CWBy5sWBJp
ZPpduYo5TSCYdYzr4gEQ1s3jGT5BBIq6TKbpNqCrKXyHk4i3lNZPGjLGSrQRHeKs
ZOE4hrMwjU7uAGLuAoKDERWsNscETZgB5qfONksnhePt+6C5Al2d5uC8R04J8SZa
ZtuPVa5WQDs2NrNYYcl+4+mGJ2PpeRO8WqB9jcBXMw5i61UNLSrukZbu8x3UXHXk
6TGBesIDhMffXjVMZTufh29Bo+LcJr4QIAhx9qaBV8q85QQRYbP3O/1ScQMDUnNb
PeatK898HHjDiWe1PbzAmHea6C2B0YkGU1ZSVueignvTvvPOavD2gpSbLQuasuu+
RfxrEWFrCv+OoFBkdk9W7nyT5vn3OCyabLM5ZzayJn7JkrwJPDuv3Za7798oT6/S
/j6j09BVHbVSuGcSt+6yvd6ha6PTlXrLiz5lGB0z2wEjUkuCZPKdY2wglg8/KmJe
4bvP+maBNo8vsfkD9oqIHiGRlCVFfojpEvLcTlfb3fXTA3UonlSYHE0gvLkEnIcb
kqF8kD7QXxhQewLm1NIfD8scYhepEVB9z4o5E9HWKS23CS45EWNK9Fv3SElz91dT
stl/ntpIPd/W218YQb9W39dkMp8EUMhpImxxli27DFKN4Cs9tmqszDXdxQXSssAN
I9pwoRshK2uLOG65OBga0ST/meD7EZ4tq3y9P3zIlQSjKmTRUeht2czTKloBETz2
lG/pkPLxmfcWe3qBwMDdq/lxRLI1d3jotb8C2al4Sdg6mA1T4dJ4XEvBho/s9d5Z
0B7azco0YXZirq+15oEXXVoAj+bpWJhULVw0uj1lC9/vD+NToC+bsq7BH4VqUvLA
NRp6mkyQ1/igvJlBLgtzXRQkxo3+8OA7HpmkLNBJ/kkSAmIk55KZkXN2ssqllnou
sxsZEaEyY3U0wPZ6t1JVYMXveob6ebVroNjJVRx2vV/dgAkWI2T6eLku6Jp9iyrU
nBpL6pM5a1FSjCPDhfYE4iErI4NRP0cDfCfBpdfbI7Ny0/XhlPLGEDFWWtPkBcTL
JmEDqheVAFn9TKdUTow+CaNTeNUiVCwD32qyySN3xqfuJaEmlQVdiZ7nsnM89cdl
aH+fmjnUDQLCU4GJ/Cehau2XYGxE1eZZz0XP89IJ05zVpmmC8StqKCZPzm4s3uKK
DFOVucQ0U7W9CdEQciDKWhEqNp3od5RNlg2I6HvEngJMbeUdywiHcthrcFYglDXt
n8YaqVqPk9aSiV1T+EbdTQze5uMyiMTq64tsZswGLPrgH5efMze1aTteAUJq1hEI
SqgtCKUrwHtpK4B1YhKhkMeSWNTcPZXuC0GYdC87i2Za2lZUhU1Tu+NszCBxfdM6
G4Nu6f3c8DULWNQuSJLcXgG4gypQOJzbg2MgIPgjNzp9nk2LBPy+4+dlkx5qbCi1
Vb3yB8ZozTKTrBTFhHVXF3eMP4Y/yEUPs3HKDAs1IxAYmWEpd1D3jLOHlLMgtGOq
p/KQomUhTzO7zFzZSCdIz1P/IRUMQCtHUw3qLPrNoJOWTszEM0uSz0efClMFV1nb
ALvzu1a9TGokDL2VNV+17tdukyinw4k6vfsrTliSu0ElkrxNWsqWSHoKVGif50MF
ECtY0HpwHyMs7+pfuElvdhB3WTRLs71nh7NCiE8KeGSzP5ihkd5mC9yl3qAuW/vf
bouxBomeAR8p7ZhRJse/MCnq6eJu5ujLR+zIiUomAMkbNTxSGizbdFc4GYAQ7x0a
U8lDXGMEKL/m4nGNOYUcdWdxnmx/ISv9UBHVsgTjCJJmNogAyIPZ7TsgA+5oHLzU
QFqELWhAufSjn1zW5P1O0zxhItnRE/VoRMK9BEHabeVtcbtnlN4880s1/Ab/8zsU
LXINh0C1eYT3fj0xZwLzG0c5cOXtV15mJOU0JnxT4sWvMFEQWQL2/7Wv5+usIAXT
uwEck8R6v6SbubE3nYBiJ6vO5SIrDE0XBMyYASSAaUPqNiKXonawBrMb+/XCXfko
P0gtsHif1bNeoiCw2XLxCHroblXTuoTpLHW1cCZpxiXqkMS/de3XRSyn2LzPchDp
T5QQoIPCGpj23hlhYiTB9ww1VMwQ5ds9VkDO8IjUZGy6tE0OIIUzKm05fjgF/oYx
Ry93IWpdKFo0X7C57/y5BLq/uuxN1Jrm7gSKWWNlyoaQUSMwc88Id2NSEao2Qrsu
tG0eHhMxO+hda1al701QvDCXQ8sbdipLxQgytGld5ioJFdSRfEN2AUQDkvgrtwCe
KDKyJAdbYJq5Bp9V0P++sjt7lAHFgvTSkjeepY2Km8GY7/Rio7R198DaHMBP5o5v
UAolmj9QDyhZlsu4huHCbqTXceCVZMyNw8etT2+eR1UHFRbXh2wY8ekxvJ4lLwxe
TXPnJKv0JgI/c1PnDbo9/oJaHVzIxySgQMmZEzrN3dt87txH1CskO0+BneRsA4dj
uO1ZXADkCbvAU5K2OfMg65Ju+bsOTTt8fgXp2N69zZCWOOR6vy2mCONOzjPOry4A
0wLU7A/h33YAc3OpD3R34NippXHmflZacPqjEI3GjgEEdCm42VvEm+5C1KmViipr
MKsGavImisHGiIAgXWXU/tkKRV4FgIzlbm184xyUZk0iufasCJh7E1cuNovl5hWh
gmtBAjM1i8Y6SBMzKZgGeM+l+68G25ujHt2SP/3etLo0nYW4v4oTCowKbtsMntxy
480VWA/yKagd3uv2TjppA9/Um46NRGhsNdFJd0dFc+Ko4yvjRR4PL6ZYRqHY/HJK
RTkgbNsWKDxQabGxcNlA7wX9U+xqbNAMlkoccH/Up+z4unGu5h2XQQ1kktX/aH1a
1h1ahhj8KWLclZfp7yHZ9zRQMCGOvuIwV0IGynXgiLrwox5EFgOvvEGyN/GRPXww
fkW8wiCs29w6yFtjXL1rz/i2LPmCXiMSM8Ur8X9KXcaQAbDxUGun131w8++s6Cws
swyizS5xhyMf/4fDd/AIBNqubR4rU2o0YWzqJ7b3s0e3E/QXFXpuYkxAFwolpOLQ
0MupgM4nSVU+Tg4ZX6ujD3dDSFDvlUn8IZYkYDtyvRAxBPe3o2WwJy9345WNMZmb
+E1Q4RxAjpR33kOhP+8iS1G9KGbdNDsyoPY4LbFrQeo8oF1O8izC/+BgIkefkfoO
g+Cv7kArlWuzL5WKKjztuRojQwRKwJK577AuudctL2oOHUsgDEP2bqfW55t55vEv
dZp5z1dFyXB+0/Sd1bs6oRJmf/n2vIYFNwP+u+FGt/6o7k1AjG0dUbVwlwjJ5T7w
SCAq5q+E7kocNX1H5Xg2FMlG/fiwIrd7O42vievLMO2gAB44Yp7Wrrky4zlCZQuG
gr1NphFfBbjtQrrBDQVtnR6yagkWfVG39UVaD8EITSBSmPVw9GK8hiCVG4qEAW8V
fmz2LHTCQvPEuR+bgyXGBIGuOxpnrPGlRTV5lWlSmo6wPcecLUk/HTZtPb9E4rJC
R+ZjpU/RNkjuFYZg1wwe35dR40/66Az8J0WGSZcCXWKr14bKQumiAc7bGKsICniD
Bbnw74D/ISzvBmp1vSV50wfgU6ACjFDrr9sR7nZyeMya/s8RY5sH8iTb1mLvSA4Q
ExBetIw0uOpczARHBKEKuarIJG4KiBCk3R++53jXQhW7Lxm4O16ZoPXbp9GQHdAZ
UFjxWFSNGIGFq1YvzCKUO3HVJ6lNQEkwXdOWGpAy+TRuYmZEQlwGT3HPKnbAv4u5
DeK2VTvHKjkgqsucfl9HyYGUYjl0HcrMrb9MrnjFWRLcNbIQ5UqlX/vFLqVXNsSF
dCSUZXVM0nGu1+TGcGk2NLhZeXDHFtCXS0d8r1dTH2OkRjmEg9x3HHuyhM20WmZ0
8zYskSDp1c4XINQ60VBJJRSVOHwmmX57bzsfKkynaMCF/bTJNzc3nl0hKB8pT+fZ
CdqPgrEqxln9ZaAvtiyszvne6UPodP0miJaOCYviEWQpb8UhSwlI6VEBGvok4VNZ
vjRxsCK/qoPmGg/ye+rk2B5FrNJGLZ9fR+VbtwS8yHJ4uM1GjbOYwXHCDu9KI2Mn
F5R9tpylT8xN1ukmyjJtAcYxb3JbHqWorcms0gH676cZpBFyIWFpiEDIpZcAFFaJ
EyQ7bYIkUtf9EuYGN89UkTjdptICx/9Kc/KVKx+kjM57Ab46cWUWIaCaG22AGhae
6EANgadGtuBKzhD+lN+84BfiSqLafVnu2jiEGUbUXx7CFHIKNEU7BVmXae5aGXgt
tkUNFjFwrh2JXnNgzjlTsukfA4tfbZx3AHbSUyDufT7o4nyhaT/yeQig4+5LN3ud
yUiDiuTxLlikOx8fJVu6wFt+a109v5DjDBqyRAyi9Hp0sf5waj0NxMukuRgnRmHG
vdPhUJTNOT+5nCNSp5eZTnMmZHu+No/ycOT5Rttk1eTiucyO5DbuUlSHrF5Vgn61
rmExyJHAtoRve8W3YjrDFYpzo4HuMLapNu6QLjPOeekoqnpgv/+X/B/ra4U8wuFn
zFkSfpdSNSP0jAodMg7W9EBJK0Stkw0wwlcJEOSiOiokKVjPB0rXTsVLreQzdpn6
tgOPILmmEY0rMKZIHE5kZ8zB9r5QqHUQj1RGmpBBHYSJJc1aKJ2obL7hgHb0Gj3V
EHnPNwzed/N+RLcTI7FGTrC7Z98YYeHM8lkQCj0HUbSzaKWNe7gRvIf61YVsPf2w
oe6tl2Eaf6+flV2ElIHL4UjMqyekdxGiEFsJ3a6PJmPQgl5cidZiNLKXkMaSVdm0
uGjioFfII/Q4qrO4BHkKHyybCS1Pq5XlEjiqrX3qhV78yqUeRIrrxYNQFAGFbnce
ZChpnonqVvw0ET9ll6FrV0YO8x3f7rErBHbiNUbl2akONMQeXIgPrM38m6ZqAvqn
hl6HQwMBq3tVz2pQk+d9JuWYR96xs0gW85a3M47GVQlhRqawH2sicyEcSzX1pupT
fjTLQJWjwGLKi+7OGFm7V92C+mpih7oB5wrKruAG2FboWa9iP2hoKLlbRk19erbg
agVi8fvqKIBLivNfg5NFzr5DZc3wvsoQPrgV0GQ/wGLPYkIrbnFpmUUw4+G/sXgc
IrTs7FcC9xXNwuDuiv/YOw3qvKKutQYfZrX8TDhPDtnlN5ySzsuU+deB82Bi0moj
2B7lJYHsuzr7kzfS8Ubxz4oauzptjIdVYVSdg7uxkAUu9VnXSbh4LaS88SLaGJYL
VS8E7zZAJuhdc+YjgP8Q015Snzud71JMpcGVOX3Na/hX68ct05nYvFTt+oRjfn6O
X87FWZA2bLYV9YiSM8hDp3C+d6VC1vW8WTfEk7WZBWP8TvdV7YuJ9UAy92Xxqx/3
Z6iVdEx7+sCjOcxM68wfbj6GPb3SGofdCD7Hmn8DoIlrcySnprhD334qB0rgcdIN
LWZAEqcNmCPHO0R8dPHGnNw+0DwXOVP6smXc0nKgrnHmgbYsz11tRqcg6ZxtX4XA
8JHWt7HdD84xJW/tkydpk86xTqFZEYv60/R9667femZPAvqo5CicRyyjEd7Su1Jr
NnIOYU98OeOgzFpltUduZGzbsZfsTlUeUI37FClY55zpLcb0cEn3gOlJvADSxX4r
JoOBQgwMBTqmgOHQYGiFoQigVB6vUPHV4kmkgOiYswjP2LAzgQhfHbE/8mjtCb4x
saJ9rm81F8em3z8MsmcrMFmkYxMm5ynpd4WTpVx+Jf0zjyulaojzmfOlThGtU18g
oqm+yptDjhwBsP6vx5VCB52ZrPaj5snulLOKKUmdDjQX73qlGI2G16LMf/sdW3KT
6bfLWxQcHiOD9yhERUy43rTxmN0VqaLEwW3H0T9Dvpmqa8o7MCSkS14ppjAzB1NB
XuYzfJfXYvbeAURWE/98v4++gvlb4OChFBhilg9Jwjp8Lrj6ucekrc73MTCfHKZH
4HJWOZ5+5Yb5/w4GPegu8N+VgxOFk/Hc4UmrRjl3GOa6fYzLpQZbjzEcVQ6O9CKK
RMtEnc6WQIVg+Zfw4xLdC0QLSw3mRhPFEC8oAESu8EyUArNO76vt9UlOt/GSLqHC
Go2pWzfmDo86A88fRkkySLGz60AOBIhbxAh1EuEHp93wpgWLDiAwkqhgiXLOMGhG
uClNourXg4rMOsLp11fpcEoybS5/3N/EnDVZH2Fd2+vMRBnqSfgKFKjdj5LJL5mk
vvyKcfOuZ6a5UBwgOUCvEXaINJohoQnpBka4OlE7Vc9h4GibFWpGdLQv82dZwVQf
aoOguGo/kuN0VwGS86A76+uMhwsnYhIWRYu5X86QimeCxLd0ZHDvwpBLavAp0xMe
0X4QGgEobiE5OnrqDr3TMFkJ6WLp7c0DCCCR2kuOsvu5NJKh5vCvCJ+vNQA9B/sR
MsZEfAL7A9SWQFAbHjPh+7lrKngf3wkl8KAKYV/h54DaXBYSTFarjzZezWpQnwC0
KG0MnbJmFZYHw87J7GVQ6LyyIf9gXRYeNgrrQVtregr98KhBxQsWSgDNXlSS8gIm
ykZTCefd+jLki2GU7sNG4qm0LZWyT7bU/i8j90pbIJHLBkZSWfzHDTZ6dLwh0MTA
+MjYHpyQoh0ToQCB1WAEeIzq50jBCT9T4cvrdm3bdgIlDV+oDH1dDKAbDBcLuirD
yTDedQ4KaRHpNsxvkk5enP6VXWor+n2wPMFxHJ1X2eEG8P/K8+KaN0VfNvcf5JH8
lMnn0SlJzJZv6gfdXJsyK9GqlfA3p6Im6sKul6OVcOwIKUMDYmT2kM7Uo8nut8op
7spJw+oolXUJOKHz/gzsjvLgNJPP1UVQPiJvWKVJVSJooV6PJItR/rLWCvYaZfaQ
ohcEy/d/IFDFf2RMydbEYpyDO6DRF7XC2qojZ0JkJQW4TiGx1cpUKsDhHe/Sui5z
v8Et0GZRSQPFqhyg6NwhMZTYY0u0ZRPIJTm5ASCuOg87gHBy+7fbevY8I6cb2ob8
cFBtYB5zBeiqYXqEB6dr2cWJ3NuAFl0VM7b3JQYgz7sdHN9Wpm1ypN1gPbJnr9k3
QzFsBIDq/IBNoFAABJ+GfLtV9sb2BmYvNTS9T6M2N9xlqMsE3dFN+9oWK8hoqGLT
zrKQVeO1dp6O9P03qq+D9bxJ6z2tCfqeF6vUyuimJBvucbUbjxXyy4U4CinPYt9j
rg4fyizIPtP3BBcQOVLPyWUZgnm8g72e7P0hrs+WMmIwPcvEOH6oqXVzf51oZ28g
gEm/t22do/TVBAri7U4iV5wKUkLmQYA//fwjR47dOoq9+zn5i1M/CUo791anRQkI
6lzI83rNFj4OCHJbF+D20lQK0EfHVApS58H/yIXaOCQjvnPuUwDBHT5ShPBjSq9j
Fel8Ehs8eclvLeBuN0M7SLQAVpZV5B7vADlLGnRerVBbHq1HZEXfdkFPzR9SmwtW
Q23VAZq2/3MwF9XR0rErf4J+E4a7ecHWytdijyYihEf5AsFBuh9Hykv+OatMDfc2
LUTPI3ErTculLLNa+ZdZerkLLyotE45kkHhCiIm8Ogi3Zh49l2IVi9i8l0lWK+QI
adqn32Jabv6fIS//yFZupNKvqdMGWNzgmSZeiRgPcXVJ/cDlKrKdKdQi/iWNx3hv
WES2pdP4j2QhmOfbn+2MGFW0apw98q38VStEqzmRpW02aWwTtv1khyfNGlr1QYt9
bhyX5RoYBS56r1uZp3mLx9215sR0T2wPRot+eXfpZsD+l9Eh6Naq17vN3+ejbaL8
DV8/jAx0i1cJS31Ri+VrYq6rPmId864672U9IpF/hIJvV0URrSRkW8uDSmAYOhXu
WW1YNowYS2XAQkncJ992E1HwknwEetDMWqZSGg1FJLt2yw/C2KHhFvaoR3J9kP8e
2rHUg3KvpEdMomljd4aubf1tYJItxbWxBIuVfRKx+5xLtc5w2cLgLiKJcteUSNIU
7luHdP2lSXskFECkrV5/n2CB+7+Ni3mzkkztQYQ+p6e3t6sPEu8tIbdlUk2UARtF
pWPH/P5jAc1J/CLpScwsGL9OocgWpDxcFcm0JK6YaPLGKZCim7IenpURxYQoY4TI
3yxfzy1Zbc6VKevfyuYOsGxFY4vXi8GEmJWNsG3vIno79mAJlLiYCB0Sv59uqYlf
x4yALxiIR6sIf94N1PxGzZyx1kPBPbEwS1aQF3sLvfUtH4QRoqFKRhan8EK0rwkK
ef0EjAIUxkgDQ8JMqy9yfoQHfvQ41OG37GgcVoSBhaPed35a/Okx/zSyOOUIu9sA
W0OZ2t3JWSbTOu/WmFXwNl9cGHqJQ8/dxmGnyOTR1FjQZuTM4VtM9PKHNwAFfXo8
oxGFWRvgJzqpKk35uJeN0/spW+TUU5l1sRRcvIpc2meVxFd8prgv8//yPLp6K9In
XNJ19YlvE1PKJaewtIIZuyTH501PJA842v8S9sATwo7R7n+JYx663LVXuyblvDQ1
yBYa75tcOrjQemJVRksJB43c7X0xUE2PWjx+2lOhjkIF96UIFzYc5888z6USFcPN
pF7Sl8y3JXj/VU9vm9kYnCt/HIwc/at4Wu4l23gAAI9uFUxlf+rKu5aBktKTl4u+
S0YiUczpb1Gjl3mFr7eR1y3Pw1l2eV2yj9x8kYUhXod0buTvPJ7OosrRNEpBZ7vG
YAUdeKuqXGLITrYeogdYWJBg3n33ciSBI4B6Me7+0QXMwMQBFk3daMW7am4A0Js/
phyHCQkgxciHCF7fOg0hvgJqMkCyxXPoMtRO5gxjPvVKB2j0pfnAKXr3EnGoDi0j
CKzxMV1nZN0mHHHC5Zi88UIRVQQFXvYzuXsZfw4o2n2cfAGhUlncCJ9rtxhVVcoM
J9At7whNeMupUOvrNyyTmIVvB45Lfd15sF6l0pMOZ8SRchUE/ipf2jA+X4H8K5Z3
ii67xBMc3h6u9ugfPDts2JbtMsZPBSw3tGqBL9al4nvz2WPMN2HgKObWY1Rb43kM
HUWp6QUrM9wEOOzEUM9Zb/f70mXdBo/U16PBF3radnuG+E671+6W7SrJYZUOgpLJ
EU7nWlRn3Xr+CsAv4BtceHPdtiutFsKkfCDT86oBDI6mgKgLoewlvu00pfyaCWce
iiagNWrYT1elVTcy68DiDnAfgoNBJ1JuodZHmsud7K5fIc5pCmt9h9XTGtrgsRyL
kIirOuaAxOzVytQi9D5+vmsBn2K8oMlgphsjA7+EX+f92Zcx632/TY7fDctXg4KG
ntgXyd9k+5vSfZTUqgturQbecRg9/yXnLft1A2gb9HHHF3dHlniGiGsejkdsnKwn
aacbbuK8ig0SB6b5gDlijffl6OxlO5Np0nb69HYyrQWk9tR3kl4GpKPYUPKQFHsy
AsdH9FZrYv2c15A4eUqtnf/UFY+QBEOvx2CpTlBcQWfWfpAsmQUXoh2uIPzq7Nks
8KM592dDL+Sp/eA4o6L+Nhm9wR1AAjkdFwCnO0lT+AjAOYwijH/xn8gN4jX601zv
7ktzMLqi1Vl6RX6evUxoTodpvgnoU0UYtatXxT0vAE2HkKKL/FEEay/FMAK/ZZqT
szUxEv8ozo/lYM6oLZUE7l9bdh5t6AmDcV5d8qrjJYR92QzIyhL/ZUYfSyQ+e0U/
/UuFgZiQUOXTdQXATxq0CamwXxD6ZwZt/ztuTw87MqgbDXxzaB0tN0GWB10cXNRa
BpR5jBJ8jBAeGrEikAoEg98b0yTZ4eGLnBLUx2vBPb7zjwOC3ceGrB6hxHx6ETFB
8v0Mwb6fEoCTLl7oxo6EeRAaSAE835Sv2h+/67Oc9MFKofqX0LDoFq0YyvOWMDFZ
Qdvaf/BGTpk86UykNTLc2cP33SSC/ddH1cc84WKptC6WdLUn+Yf6SiaN2Oqi5WAW
m1vGawx5MTzX7zWNJMB0ouuPoxV5bv01LZy72mxQNrG5qglsqHUW8fuPOnOujdgi
8z7EW3zVbCZQY5UYSDhsCJ2PyuZatVroZ0VSMUGLh00G2OghzEiC0g+lfVh384rM
neIAtLA5tlTvffAKwdPpAeAlrjaAWS/SVgQldyGXn0+OLxCV4tnF2hvs0scNoaVA
07HRtyU6wlRNGqtXYhWgDo4n5MJ40PgbNmsfqM6LofZSAkfoy2ubcVLrwfgBY35D
ogjwS+VJR/6bkIpMbphRaxv/trd507DEOYvQH2iinWxORUg0681zFTTxcZR2IYh7
MzLddOqY6WPYWiAcS6cg351k8mW//HWwAlKsVNU2Gdi5E5gXq/dm/VGUXNl/C8Me
35XD2fyXRPXNv1hEwfDcNdO6hFnnd5u9qIa+lzeJHnpxcuH0nAo4E4ovBeKBpN+/
TG+/+BsUaaz1iFzfiu1w37IyS3YcORGHxs9vAEUP8NFoujh4AKznnXlYGxyz0MNg
rW8NQCaIXTpOGRqrVM7RJrQXTJjH/mxObXyHjbbkUqg/Eox8r8d0CExrNRhsAY0E
Cvj+X8gMkSd5OkgQTDGQ95RXDBTFEmQP6SzqwDa8wxYneRc8XvvuooQz8JmamTyQ
YZ4v/wue9K2lFXt9nT1FZKVFgl+wTrE/lBrPzEfGyXmxE+zRSv48ShLPXkQ8u7T1
8WYOQo0rb4vYVKHq84nerc+rFdTd+vPyw+UDPKQhaTMTY8aDceFRyQjqrXqNFNVR
OxA87Zcdav3Sus0VzmyqmRxh84tJYnyC2/sdESlAprMsgCtU4XaDLmI7WcjHNZrz
SZCsb2Rdzvxi8joEACFED+692JGkzcOEgDqO1eNrFDV/CtlY488ioA4JrDandZqm
1OmCiq4z5nfLBg1/x8opDTN5WJaLNYNKapWVF2pPmOVaRitQN8C1F2Oirwvp2n72
LGEU4rTZUFcBmpi5Ycn/vRtbwmqAI6ONttsgLXqAk2d3p7mvwihFEdtndsCgeABS
wK2JwnWg7BysLgzFRTc8vqNv+mKgBvNy4djsZ4mfu5OucwHM3zdV/1kiWMgmP4lU
2mcRueGbJaTV0zy6VM/c1f1TWTfq/lw6w13PT2ikosIHfjZfjcuBBTn5tDhfh7jq
71MCeUhCCdJ+KK3RCMXKADncY0gIB2kydsd4LzG+DVk8v51cV6uh7mMFAsp0lNeJ
czjZiRQSUgsp7ILmhP0gbD3af+rmdTLvU6ZIgKsTzy9bjMoJTlWdGZC/GKCIT72y
CR1VRdBQ0R3gZQiE7IXklsZ5LVGF1ofjOYCFNbn4CdnyabbJx/A2yH56Clz1RhoV
LMpjN5XXRhmxuCETsGlv1If1V3Z/7oAjonEybhATZmSSVlIXmzCNO5xxghdMZ6QU
dh+29UEDDTjVT01UuNfbJ5f/7fqNSTtKU/qQVZJzTTwxOYiV+DFBlldj3joARGTw
QvTrNWTqzaCtEJQ5CeOXArYdDTr8wIecowJgI02D6K3aMkhYNGRj9EtvEklTWa48
D9sHGzTVzTPUx9Wb74E/pj71QGcFd1NDPCjzF6yoHVnqL964sagzIHv2ZwScdXMo
A4PieZn7dblWJHOeowdmcINe2rI3ztJOMJ/+9iOWmpS375ThuhlWAw+/wDxTmZv7
CyKD6QY3Dc4lwxO8vNG8ZFwKWXj9SEPHGg9Tyf4Aex+yghwkA8GSzvFzHtWGt4m0
KtQ36vU62vM5nGteB0veeHwHXJOpoWfh7N/xDX1mUhOd4wOcRlykhuTjGNnRjUAr
jCoNbGanf30Y282MxehWipQoU/cM3vK5PndUiqAMSu4wIYm2KX8YYXSmZ2bLwjwo
oGG3qJTr1Cwd4E3ejZ2fb5f5FbxJuQhiDXERkjnJrc767gNbppfpR5PLh80u8/cl
GyJQsXs0vYz1aP4b8TgSqmkb+3yH4DGIvjtKG7mmJ1s5bP9uVPW2FUwhHIvLnHAJ
3zrW+X8UFR6WJoFR7LWDhKMxfGVYMWAeny8ALqA2DPrLQCIh7HQ1PbyyH6icpyMy
ot9AV6rhnX+tayGq1V8kMBoIaufBU2TG1lnYiIfhqdGQ7t9k/uteAIWVbkWsZXMz
zAAbNL8EyLV27NtuwJPbIv5bOBr1OSbRVXH1hEYSLcPQGiyOHF0un2w68Vl6CrWd
6LdvtB/X1/P2FEFdw2WryY0muk4Hc4TizQG2q+o8l/uFnk+zMWYOuUyC7Vk623TH
CGxRSkXKvpEdcimAy+P1kZSxK/JWXA7dG+E0v9HHcC/Lw3huMZiO7E4ws8mEa4T8
8q3BxRBE5EgPN3nb2c6sSQGsS/lOggToQUDzZsRTfyml8TqQ/yk3IepJK0NJsaip
l2foTeZsTu1i+xcbYmIiHt+aJR4N/nOOiVuky6jrv2B2yji5iVxXZpJrCxJb7BR2
Jnrf4+TfYMIDxKtDbc++Gmwyyc3CUJMywHbss+2+GbYNNoHG54bl85gkENZq0rRZ
v8G9FFg/BAw2W8CusD6YltX2LKgW+95rlOewIaB0/fgBrgFdjyTqX3rccsiX2Tq8
dI8Gt2WK+K2a/hOStIRBQS6/QldhzFLwzuFR22CObH41VYSAFWoh13jyKeZmeMKf
YKUFSZMaQkWDYoeRuwe9dcG413UwEdyr+cGlaQRqmnxDJnEWm1lKKA32axyKtNuX
mxxsIMgh7Fz9cjRNbwHeQyXUlTZ4ZOZ1oDiZvel3Api7CImrymu+0PM1hMQHpWFn
vxnfP1epeDHUT7RilcU4fuyADIodElZ1D5kUPentKnszWravRfBRGxx6uDlI6Neo
Zj7S4dg+EV3PbUKPTVafZbCTe/dFi7+ojuEP7dNhUdhDBfvG/HNxir/2wi3j8CU0
j+XMUMJE20Pan1aaNH+hLGsVwlxspyJamoBsipXKmlfd4dZVlp7pn/ZiMxMb59Gu
Y7MYATX8OeDWirl57sbFMzqQXEK48iytCgBWj1FD49r4I6W0NEIy7Zvj/JrGQK9I
foi0a/qvb8ssU2+t6AxdyGazSNsHhMF8V3mbHHS4Epd/QMdyGzRyUmJ2w3fmqULn
QT+30CEJWaB1sfe/YRTu1m7D920nz1kbmk4jICGMimU2dSN5N6fMvBBiCRWQNSaB
wJxr7QYFLEEvgHeFGDBfJ6g/jebJSBfC6PrJL60kxhBJ9UKOlFUOJfh/1fqFpU5t
a1+/3KNUpnFTT8g+JuGqWVUtGOBqphYbR76ZHFEv64sVJS9eaTb/3GOkogxLkQpp
96Um9SI0AFKIGeMswJrVgZF6mNDWfDHB0SCldQZFY7FCKBLcyQLYQaeU1U47Je2n
ZdVyyRGyu77bOdX4pr5xXw6PzVQy9ERn0pfPZelypPA1Q1EkGJaua1MAWrFJqvVT
ScVfxh/nEoidn3ru+Kh0P7F/efKVUqNSgjaQui6M/RcEUe9dhYEv8n04ajudaigv
F+BPmjJohOKROZ41/kxqFFLTWuJqkRl5CoCGMRDSqtN5UqfcvtTnuNKLBKmBKwIZ
E8QEcErSXT4x1329nGpBTSbrw95wbO3jCEiPrLBlj+TH89rnORNn4UkGCHEceX97
jQQ+UX0TXdmK7vp4n7GuWlkjjNbYXvZj6xzsCvYsfF5oVcleuYtGGMSNYiFUYaJJ
6QbgR2FU0BBP/Esd2ipMA8NqDkr3vuFo/FLaWY25s4aGUVWvkIiP69AyXLPjDmjl
BBhcguDRsgJKjCQ7NkpvK1C6IIRj/tuDVXC4S/4iyMzIzDuYaaQVRWjV85QYKhUf
FuFSFfy72/Msfq7/IaBKwaPG61WwOElp7HXC/5WPjoSCj6p6YukRFiu3lSR42iDv
ZC2Zkz3MYeplU0uITaquy1Yh6p2yrkeTEAUsB2OOYEchQrxpCb/5QxGfZBkRudGS
WWJWYR815d8vB8Jqljk8OC/xPayLT5cJEUdKFQNU5aQLyyvVweqLfnU69hLBssZM
EqcvebE6krWaPg5EiAGgrn6U9Ahv60CuzVrr6vByfMPKXly070i1C8W5jYsl5kDP
U6iy1vBcsNtKMuvghNNd+8OU/HLvRcyKIBXY528QXuQVtRucRRwtBXRkOs/lKUWY
SoyQoV2ATwej1/B5tMEnlyVJw7PkDplyEadj3zIsK6Ya06tSjHSoXmJShVJewS2h
CXNynDnPcixQuPnFiTCFaG0qcdFubrvdk5WNs4oaFzdJKDvl1utiqDDlzcg1m8Y2
wsEZP6ZisNoiSnkrdHSBz94ZeHqYi/gDjWjOYw+XhXHNRvFhgp6PaM+aRN/0Br4j
jCZ3qwgbkUvaAPdYZ9fmWF+q2CrDPVHd0SzpX1WdMNAMjEAe9a+UzOcBk7PvrOfQ
VXKZhcg5/rh/vmuF2Fz8rW6kzTbD+RvrIgVt/qciAJc6ibSNXZGtS0KS20S1jfK/
1o12yG3PxHJ8RQBEpweH3VDI8F+1RoYwTypo+6Gw441oWqg5tN/SK2hINPVfN4M1
TBO1PNEhY6j1Pbkp4KxS2DniOOWosjFmWo9HWS6HfhkzbjplanEpVAKePd3vNlHe
H1sMbN2eqhQ8A8B05MBCQbU8gSJe4ZM4CvqGcm8vtHGzJ4z+RmdrXGRCYxH1TBwG
tVWUV9EPjnhf7lfvVmtAMFteJt1K5XyWtfB6pxlbYoFdmEjWzdr1e5qGungaawY9
X+3O/bPIFWJ1rdcDtuPD6+Wz+gKhcTuRcPYQheSY1MzLNI3sXUWYtH+BN0JZXCib
9MITBIbJVNAV6uWOjgXhYPkRoCKEYPyQe1U/WdglvzwapnCpdlK/IwSFLSdj4eHz
ENESji1v5kgiZ0ApGNiwLWxcYXB9Qiep4ETGo+hLPRN2th6Qf5tJhqO87W/yGFl5
tiRQtNTLn4ziZvU9p/SFJcO+TjqZawScS5FdeFx4OLlhc4GrzWcba5M8OSKw32Cs
6+k3uuEmsrA+SZnQ6Dfj9Vs/h8jey1EKBIjedXA29qWk9nLFsd2UTHqwZ6seZQcd
JFTIVIgJWyT81JCodM7d1fiPMY5Caxmsw84plvdCYV5Zz0KrGpnFHTWIN/nzTDRl
wXhoTZDwviupLxXMsQsnzSNlhnVjwPhd5Vz23UH0vuxNMkccwSY+ObxnTVtT/v1V
2Tr7GO2lJi2cly3Htq3m+cJWy6J6ZqH/1cEkANVfhAVVrif/dAcnwRYVDsplbhpP
520XMLD0APqdUvDtafzehELLvX5VCYjHnpZWzwy0wLYtq1EAS6o+2fzrCi8NgnrC
Gfqg6jWnNZP3SIHwt9fuDtslVjB/pm4eFG2ebIX8pO9Y5sLL8/A7jlM/T+4Dy5Cv
pf/NvCb4bqBN85pUfbal16VDhnFA0u7NVQFo38XPdJNE9l6V+Ts2Dhfp7OvWgyK/
Zy0GjH4++gcZVOWagWeu9OidicFXg4E/NV5WMT3hRSn4hZBKHEKpUcihLgr4z5jH
H4Kk7VVPi9Ss2yPt/NHdogVyHbiFdP/tqSmg0szWdmL3qaWg+Eth7wjJwrJO/C3M
npgVb+yMUcyvqnO90T0HJ+aKhpKpnbeV32v1qDem8CC6WDiLX45IAZWZRi6AFepw
mbAK7eyv3+I6U2qPaRZuEdRYOAJesZhKzK2DMD9IRobM7Vi734XMj6eO/BapSFWW
Yfqivm2pWaOZVxmr6xImFn1nKntqdx0Z62cjY0FVMkDyGjd8IXBzfsEbEn//v5pB
OOBUTseKUg94XWDaSJZpEGWCgC2LTzeFz1uaLQ3j+42wKYAVx/yHzgPdVoLoBB+Q
GD7uDF/GnYCjxO4a5Zbn4TTBWGr6mk83QShh2rWTHKSRWYeEpwqVYHoZ07wuhnBL
I8ek44bVgmHcYMpOICgSOGhypOZn6VPA9AXIeAIHUpBEONAYb6PnQsUUaed2ZWrG
ef6crqtGyBIFMY3lIhwhy2fFi9M+0rzUnMwZhcN0saHL9kze6r1ott61yRBacBBp
uDqmQeGJOJN8RA50MSCl3ti8uUw/xDGBmzFtw37gwlCh0E9d0Pz4jkPc0lXUbDAM
0V7EA4+1fkSICmnsJh0YintbwSOLExrorIxZ2QoX8cKZiaPSlu4KCnuY6PD/TNW9
f9kCI5yEB76+bas27kC5DNzC0n92KROvwuNutNyNNmoOeyvPa+kZKk5hupVp1Jfu
qJrdWLkIIHKOoFNryJok6MmCHAMcl4xTFaK0v/MXiDfwKlc3LVsv5YoMsZpyl1c1
g1DHfMCCVU6dj3aeQGEw38t5NFJczcO8rGjUmGj9STC5JVpy6uJTObqRldsxf/Md
ncSxJA67dItlSmABKxbJJlBcMdUNtr05/z06MNhS7ZJohNhuRT5BbAqvg8p+J/Q9
ZnKGhSPhpJrg4420ObWA8TgBovSKHl3nMmaVv3/qUqWte6LF0N0vB6VRnd6dwrtn
vLZC9SlCUQDPuDzgBM97NpM/DiiGH4153G03S+equhlW3Kva7lvJc0rldBIgKU9o
45RrjC7tRHh0jTwoI5vDDEwsagCy+WvKXefVv6Nv0VSioP0RnMd9PtTo3jTQTdOU
VDfD5qMEISY9pVhInJUrIBixRxFIulNu2j+LcFp8F1XCSwfRb0GXPEkojqRQ8Bbd
8I4phD41zW3TLVx9vFHOhKI6W6amHomJJZu9WDPiHKt4ejgE+djdgvxi7pLYBR3W
5wX+NR0R1MjUJpbQDwPHUAcsUHFaA9ARv7jV7G91i7SVr+AGeaGRm/S3ZbdnbI/b
dabzon4g0hEgwPiYQQIvKaG9xnIBYAFBSq51mbeH8RaaevQcQvO9A4/uCUVZ4LsX
T3HKyUoYRIluOnNfGKdaBNWqYkG4BRnZKw0yctgwH1OiIfdwAMUWIc0Sgdzn7VPE
Xb8u67GI82iSCAFrvVCQ2q4pA7O7s4sNJtwANp1T08WrcfQbwpMCio5eW1gpsYw8
jZJ/osXe2dx/0J31Jd+20VBdR1zDsQ5IdJtEEHNKXIbTHT9Z5HvdIPJWsda4ySOT
egStmGfse1zWbm0BNikYCOAjwWfIiliLfO7zbGvvk8F0WkWQfGipcvsUxOWNPft4
j6XjQaXs+ffgmS/dmSjflJ96KCzYdiD4mFnIyTUskaJgPdlDTLdMcsNP3l1kyqKz
UroQ1cV+gcN7vN1njfEZ31WQRJ8pIrf4Zycf+gIdvimIawPlYJupIiBo7JAh3s7O
u5xJ1mxVmZOAu5f6Raa7P8jHgfjcSdk+qelIRIUY5upfFbbKHxMelWYgpEaHMEtd
pjJiq0Aj6OPwuz+yfi1DNQ5xEJ6N5uDbQEx/CXnkTdRAn8D2tshTtTZwJULb4Ggt
ZJ8aJ//0S5kcmjS+OWmYh83T1uMqjbJrclNIp3Z5FVmoDQbKKmfxxFeBhGcNcsV6
IJznqvBmMtgbW19SVMZSx3R3QfIbqOAKR4neStd/fF2VwdScRFSe5sDxLiDCt/dP
T4xsB/rn7oorqYjwF9JvzIcIsoFzoPS+uIXbWclItQ7naQcOyZ2VrYMOFW7ZI2an
m7vQzoQGflLMKAykIzetRx9Qu/Q4XqpSqyMDdTV3RZh2iaBCBqvg5Mjq/XIqeHCy
4nyUi2rVekYWilRTGf5YjT60ZX0kqfRB2KSXy6t6/w2gkrloxzzhjLfiMRvdBABh
Lvw6mAwvHHiey4F0MY7rYo32DmeeyI7PawzVEuNCnTcoKBXfhtnsbr+JVBtQK31k
z99K6k2wJLNgRew+Q+130An9SnaAUMKoQaa37A5NfRphSTFBPrSqU4gYNyt2L/tK
EjWMynGADJdw5U9SPVa1wtvSuVSHsygMm96GifrJI+aGf/Wt8JSldaYzgm4XSiwC
aZGKAtGUz/ZPrtT1zGhBxusVIf0L1yB46UxyONDIa/jGVy6BqgbwqPKUtlCiu1Oy
apmozbhc81TbPrLCxP5CCh7sv0/dN2+OuuiSph7MDpLv4TbIW2otCO1l8IJ8SOZa
R+JZtqyPYBqbO7g9/iOQtuHTVKTAorbM98ERO4GlnNuuIhbJHH9DTSNy21FBiw29
21UQqJOH4Z017vJ7KOablagDaF5eZxmotu2aodnr1tsmcyjYliqThEoulxhHFTbU
NuH8rYr5dw0sgbrHwqQeih2FXiWVoq/BRId8M6kmMXnrxOKTpa57Re0QsBvy+dhy
xCVsFGqfqEyaQns//Zk0gK4mcCx3DUOP0Lv6FcEFtNIw1zHwVHokDNa2omcS5Xn6
P2fF6lLPacJza+ra53kBJPYWoa3VNxnaq16MYIRy0TYKlxksDnBe5u82/29Fch7d
YI1C5kv5Y/H6vFWm90iTH4OF7nZ49JbbjGzWNTUO6KhpGhe4hYDE0CKdPLuJLuUf
BnTnLWGMJ/73F7a88ri12gKaylIheUOF9Drul8GUgWuOr6I1/nbj4/GCpHHyoB7F
e2hPdWgOQLQI8E1RvMrnmb6FZhhbQMu/eG8CPA2ZaBgMbzFpvMySbZTTWvio2e/g
rVu0gRJpfSXbNuzcTl0wvLTCc62F1ymEGkaIhxMIIOR8Pc3TyJ9kv4m4P92jBtYL
72astSO1e4jJyXXm7E+VS2mjmS28IqYJdimQCs+jSvJ477AiFNKoQ6Dtf+pE4IFR
FRcbmkMd5HSHyO/RZsKdt2qGIGRwicWdiUuXxLww/Bte8P6MF45K5k9ox51uiNHy
fZVur77olPHtuUTEv9c65vVGpm4PT+EKy9VeQ2/U1Sv9/bdCCNozgVWUoCDfqTLb
o3pEyTGQUTFyNrl9Uv46RSw2b6oHHtF5Yd1+hlAfDf/p59yomkW3jXwtgVm3anQu
kl2KcnBMaIwXelwQaVCTv5hvDQFzGv/IAJZnGsiwfGrXn3M3M4QHHR575R04v+PQ
eWpTRTc4S1+ClhAkd2Jl8+zQZnfoY/zm8QuzsV9REOzM+izQz6tL62Kpa5bEhnFA
MEL1yVaPB8MxK5KJ6U89wsGt+/ZJQ+XS1v4DEcA3x1L6hIaOe1BVHX5TKqIFdp5j
6fUSLbhwkOQdfrNu8cC+gzSIItNzCpEx+1USN24juskPoZSk5SFkTPl0EOywGo+V
2/28zrGHWVtRdFoGkMdqQywHLRwtt6T437MQV+s0+ubjLHmPp3dmWfHOjcc6ylQG
tf0FzCT+dMzZo1dF/bagX8GaKy7JOdFPvL/RWdFhe95OyUqE2YYk4vNWwbSdlMG+
2dKrolNzpngzEcp+SBviQCDHFXT8XuYDSoFb4A8F3g3mk9Kl688d4mxX6rm1Jmaj
u95ZLIS6PwsoBMJ8cBaqgxU7lagm6sVnUb6mgj4n2kQBLIPEenYCBuV/wW1Bb6uk
ayI//40xoyXkFN+sy5no4FDgnJEn3uD4hYxZwWzMttUBuuEJTEZmZPFgMPPyiGu5
m7+5hdHlJJUljCp3iLMl3SLwX0dq1rNF68g+amJC4e4M3ET7dKm/Fi8pfzKh6rLC
tdstwetg+gjb+TInEpDbW/3WsyS7T9ihZFLf6SIKNP3AVz6lqf++qjEXR2oeP6nh
+qH7PwcfHRU91ymQpm9uSZ088G8X1geJOuFjG1XdeiXUlFcTTO+nBGndS/f+K1sz
f4Hurl2pT6cI8VDOyIFy3En86xTWv2k1byFstYXQN1K1frEEsYyL6LyL2p1WKxjc
CjT3CD2Z0Q9HfzkaVuA/ZDqiFASRi4o28C+jTNUsxFMpSr1wiOyaDYmzpBxo2WAd
MJ/Z2Ovo6a44h5OU+If9lhQ6kS2w+2uc4lOkeYE75bCJP3xtZ/Vl2roCNOaaqHrZ
FuQ1jlVovId5yCaWNeaqxGmv/fasKA0MmRAcqXHRTrd/m1paY6GcyS2EANxhBdzU
yC5MknS/8x0Ih/n7P9+w+uyQ5XmD7ch3Fcxs6telYBD1W6iFJzPWbfTX5sHsfrOl
orSMHQiioLDg15LA/nfmJJIJCzUV3nMll3qaZujMnxSGDmScGqBz0VAyGtiWb2KT
Rz46xpRKYAe0E59MOiIayzwQLSvOcX4gt44uG9NGpetpQdoWzkWRjXqc7NFlsGk1
IX+fB5cKfkakrB1gSh9Ha5q7t1POE4mo4WQadDTB4AMi7OMteD9qbiCAD2XHR1KZ
S+Od3BDHLdgE9bnYMMILveWm7PRPPl7tYHpSR2FkMm+EwpuTSluFHTP7fe9bZyNH
w16L+rJ6UqC+1J/T1ASNVjtM6WfAAVa+b1FfoqS70kzOokx8DGGnmyhXATKCRBQx
13/hiKY3htSIyurfwBl5uSUP9EIAvqDZtTitWLEQBFh5u2MFcywBXO8ITJM+WnK2
b930fpxxlC03WCifl6y3FGgrUoM7qC0wcCYKyaZfHNtsk3F/GhxBRXFwxrIWBP5w
EpbtUljA4njjTv5LMUCthhCXv0csvfFRL8G/SSmYBT1KaA5KSedK7Yaae0lWxpf0
5QCZLpJRBOKWY2x5NZApDYpfvNqjxA1s8d19DG2pSrIjFlE8LVRvxyqDiV0lKD17
26tsVhjtEeCiLPyWJnvjafqD34BC7/AYeEgXKl6rAGvA+ZS4vb3hetVLZxDDjZ6w
jaijWQnJY1lXR9XpXOoQ3GUGZpSq3GEQd8+G33yTm1TrD/jAKVQeLjkydwXiZhuw
/XFZAnySwbtzbdQW7X6D9BsaX2RDwFHRa46QiW5h72tL47YGMNLzmJpIMHpsH0R4
FkSKVjPeH577UKylEqWrY9CRHOypEOK0DEZuHHc3BHeB6S2lpPjZtzNdQBd8bs8m
+tv65XS/JTJHvJt6mzhvZ1b/r8TPyS2JF5xYK/BTYs99wwWRdUN14pLB8C4G3+7k
ABKjvGxIDpvnlNzOnN3uP552npBiI2HHenVkPuCoj2qur17pDSMBsKVhPn+l6nvN
e5nPxdUyOO6DPUAWlo8n5mOBBbuI1UNJcfcwzAEoH5H1PyyGNyQCKC9xZALcx+D+
OhPh3UUMdaKl5BWY80fqJeS3iMMRe3P6QjOqy6QhvImZaPufX7x5xRkyf1B2bmS5
PPnwnq0J0/6xp1pYUfRNPhIV1+XKETPrd69H4A5krKIiAe/ux2i03XgUWJ0BSKgR
yhEr29kvQ+ESwqv496dtxLWzmvAtU6RPEEuROtHby51ui6/DcsF2kknP586QF7Fz
PhJSunGpeo1nSjoM3IbNpYegJVorj5oPu376cgJ9tcuwke78ZLNjRZhLNDocESM+
DT150yvNR6/HRlFWCkZzHrvkmZGj5uEPF7XKab4nnHTJ+zB0SUf1a3myTiULtGOx
Wr0L5WAEfjGFVPpijW9ZI4WH9HiWcmXsvFLoryfEzO8cQFxgBDzAhoRQCaRUcCRz
i83TDCA4TklZELwvt+tN8ZXUumdb/Sc1zf/2RMo1m/yKuObgO+6TpfGvwg7QB+ay
Kled9eHLiMsEOMjoGQlrJ9BnCk5X+AloBUtsTmtAjY1rP5K+Oj0v7ZdOvZ1KPq4X
BGFcaSnQLMyBuyFOtIU/3jjSrb2Pf4XmcclMeepJkfZsXNL+RjGocDkUr5tAytKe
ebi7JbI8cYGFAywJ9isY+0X1MB/Kfyseyc1Nf+j3dqGnvXclheRZzQZOemmDyjXA
2SgFLpxJGBzssmMaPr5pNKnd45++KtIc7M55oT1BdDJqK6mMABU2NLcu106xx0pJ
AUPd4c+EtqCd8ZELwjZLQ6N8Hf5oJHXTurP1QeNiyW8DQF9+qYtNKTXje1bAarzK
WsIJPZji4uAVpfwQYd0G1XXCstnicgsNWnqd8ASAjgydsgboGfYNdDrhHJjDTE3s
FJ6+LRUqZlbc53CGEAZX5F9bi0hCdbUJlEyBwooocy3xi1toePF3TxV4EWyMNwm4
SxH2DDhe6awfOIAdUSz0P406RFyn+AO+tLHy5q7YQAe3ooL1/W8VEjVE/peSh0xY
w2Hi2rEtiyYw2W/IuDt7niKnnygRCdYWnZnuxP2jV/X8tT7yYlTORKKpjzyfnLs8
g/F8zjKScKH6EUvixPFBWBPer2TahdICaIvd9BqTI6m/IWWThVhb90jlw1mhpwYF
rI6508ED1OSSh/2HTpwUe0cML9ZyE0pIYJFTJ5p9Gw4YdWYpN2DK/26ozyv8ZqQ5
7O7Ul9kDIeXbPUTLmiSO0k955DzUMyDhBiwLz6nZ6EXJ4v56ix4kkYnfNzAhnZcW
vPwYubKRej9Pz0zacS+vM4HC1hyZigz5qKPF/3N+Ibo4+TzSOzSZGR3KedQYm+ZR
EckTml0XzFP/QKotmAyfn4v5zaw7t4ML5TMevBE/iz6FHx5EBx6aPBuJe6grtMjC
1AJqr3L7WoNIjLVydfLk068RrGtkATJbZZqbAGOYiHDj5+GjNNuDFF8uQvbe1DfY
6Rl75VbvWMqbT4Fm/phtMG7vbpyOUmEvf/vCbc1Oxe7p5dx9PW3gjC/PDko6Rium
Olyo8v8EkEa5Ni7D9CR8yxC/NdsqWeCBEv7/Sy+3EbVJMymWJfvprPl9b3Cjv5PB
DySolCi7PJgw/BuvfehwKAwiomK6mLZJHqjEKffOxK0+vp1P//R5KQAoq69WgCQT
CYSNQwZeG08NRHJoDZrfM+uUEnuCXmAV513n/6KMiRjYfzQyrZCSFs6EZ1UMDmrC
QjdG1tJ7Dg0Z2h3EHIbHIOEKxNwNM9JwS0o/ushOoqwubMN05FMy3C5oAsCjoJwU
3YJjkY/udKVjcwXN3v3i6/BwlVGikYnovkAvQImRADz5xX6tA8PWsTREFT5RKF4Y
bQTXkQMVTqCGXC+9rfoUTfn19LleCagdVPa3LjQlF1vvdmKz/jaRcxE5koh4OoEm
0gl5X/lTtEIItkcVWMlRoc5W3so3WGhZDxk88eetkQtddw8VcX0Y44Qm6Ipiiavs
sj+mtbdO323BAbaUjywvd2sOEKVQw60CXJ1HPfOyi87F8d7LA2Y8/9prqjOUVWEE
9COOV/qNRKJwAiAVJZWtiCedb1WUIS9XLTJqwc112pPNuCGlxGYFPFy0oM7Q12gO
35S3pSjRcgkPRRL5CMK44eKbS2dMRm6cuVU40i+OAbgqLUtk+1I2YMU7v+fo1Ybk
1O457G4vq9N+wz4fMyZkCGK7B+NIk8sFy+6xIyZ9mBRA5MfkdoDQNL3cl7FSAFE2
t3sim7hrkpyiT0SBi2jpIHpmv8oC7U7x7MqYXdZXNb2RmFGr1cX27rifj3pBKeSa
iHSk/UgLWnrD4kIBKo8ookjQm3ILUtJyUs5OoF/wikVDpzgbNs6TSdfRGwSOB9TV
xsD+RB5v/O0NWMmM3kH1PlmyMtoZW5uZADmgvf4Ry9eaqQ13qnSSRY10nhZTtbI+
l72uCmSE6qx5PtD3hZc/fI5IdWKWr+F8BDcCa6WGW1s58JTaokPj3LmyTgl8wUs6
Fvoak3K9LkPcSMJ4hW8yE5NbRe1MWbSev29jCOZK6T3LJyHBO2LWq6xHJ00Jiwo1
FC1CP4hXlZBfY+7NObPi4Vkyg2fw3TUmv8sb9Bofwa3+AtAV4OO1OIUroeW6C5/B
cfH5hcey8qWzVqlJYXzRh5AShT4nxP5ryI4X0qq9Rx5EoyqVa89A6eGyWb1wnaib
xUGbcoPPv1C2k38KV4V2qmrnZyHwxHMNY088Ad6BldJT5tEWRRsPBYk7Q5fbg3Tj
nq33zHCmkWik7TkX6yS0HzVgDY0NwTIxYz6X86iGlzS6bvc3sUb+nJaGa7vvR2TW
OH+lcTuPHrkOEsWf3rE8U+KhUA+3zBvTyOkoNkVBZ7Tp+zOHLnZjJUYd2R3fL+K/
NveN/CWnTtxmsFrczUAT70n9JMemUD8NH5fbdxQka2QOyXXYDZPmPaccLmoWaS3T
XF7kBf2gOyIjMIDB/Xc3djplYR0Zpr7EP49tzezUkqSUWLr4sOv9b+QnhTCeKjHY
lWkRzBVNEyzhjebbnrZMLFvOPjbRC4pkO+QA2vWP5LMGL9c5b4UrwP4QZ2z0ftEL
kuWbR9gUEJoNAiqFGbq7KepNNXsWT2q+gPyUF7LJgKktBgkeIEYKkQbwYl6uAsLv
xPuvSVE+g3tTXJ4M3ggT/tu24CtzqdFve3+NpFDzpCWRqIRxIlFT93nzFcfn9Pj6
+rV6RLoeyRtHY74YgkHS+emfWfYhrDKFn2xNlNlR2l1NC2AMG86uEoq3ChRIonEE
c5qRDc7JeneyiIvPdf4I4+QSHOzyRQB0pV/o9wjSmOdx4d6fnfHMH2B+RTJDG2lJ
OeWcitRlP+Z6bv77xJEfN1OHsUMaK/KnvBPHrNRym62aXQrav+7pkUDNOT+FDit7
alhm+nnu3rUqw3PY8ln1LHbbqHV5sjIdaLATce7nwp64rqp2vSafmYCYXMKOwFjj
wnzpjnbyA6rT2EwDid6uz65o9JDpVr6Eg7BMmaHuqAlUz2kZz33ZT2IGiOgF7jJp
rszoEdi0DCwjPfsIaCKUJRhwm9t6S2ScF0QhxbVd07U/br/D1/gBn8hZ1l3rMOPs
FJv3rDdmCxoJPXDHtQtqTmGEMY5KYi0SeqYneiSluI+jICPZlUmF4HUvBL7PIFzE
d7q1xXS4hHHFEUnwKuw6BbtE0Y5fT5uHJzxRy6+B8pR1h0BC27OdMJ6vn/weT51s
7tNIKbGeKWxLHk+X3gbn+v3JbSr0nSzG/p2Nn+erQT+L8kSHglMGKEINaBcmFzcX
85Esy5sR4G6/KKCUPcpvY/f3xGZN10AfN+TEyPrzfZE2YoC7ookZsm3AjjvvJwHR
qv0pFE6BLZwo45WDKy16p5i7fW/B/4ft7V3v7sDGZRS6EF/OcNLhxd6AddesvHs1
1hAayUwAMxWLhk+vXQwHJt1xTO0Ps172G4qZ3ezyeTDna91tdrP3FeFUUz98C4sN
zFSfh5Pnw6aLE/vS3HPKEmAm3Dpt0BhTMI7ukXOnGQcT7wkmqocUJxyPt7xs14WJ
3a7sEW+J1iof2EZrxEagc8n+mx5ssK7hpqgbQF5Bw2G+4CYWgRwhXKRnJ15PLp1c
Qe/qBnFQvRYrMF3/WF8eFXH+/DUfWsC1Krb6bcSd1S2O61nhzL+0PqOp9E16avUo
YMNyiNu3PiDxknBpfqQEfCLMzisn/fpaueG1Zil9aKAcZZuwSO4878Oj8zwpUWrx
k7IbmV3OzpKCU9JY/OUg3bxKK2UtG5dTogyWYARy5OiSkcDmdrmYKzoXe35Ji/wo
fCtegRLr1qoeVB02k31ik3PUdvh0ddzhdqOzossy0W85LRvJ906Y2bv9H1D/yYhN
j1VoCJVKi+nSmZLNhcNqjxLQVatzGRcTEBTCEcFwLYB5wQnatcN/FPpphvkR2Iw7
eLTf+CZ/k0oUTvtoUgGuFo08hb4qH5Xo4oAQ+rcV1R7z5OE9V/Z81Ys4WPlnxCq0
8EwHqe18yeKjyc642nWXDWG40LZBYSiB9wN6A8/RregiLX5JeO7ai964VH4Ntd6p
Ob4HLOBujTS1ijAACN1W3DxB7hi7V2qS+bv6i3mhWhG8SztJEI4SVlQ6S5WeRoIk
Shg0QSCGaX2tKVVeEdwVeijnaLyi69zXAS+xHueR8a69SXtQAvJ9RqXfDZKXRmsV
9XCuXwpY+vWkGBoYFc88Og2dbdN6/avoDTO9eNOz+bKgTG5ploQ0rOMTnRXqhNSA
8Yy8hTkdnLLDueq+FQqVqIcfBfZ2I6oMNY+Z0Olil0L5G23ATlFTZgQ4wAAYH7CG
J7hqNZZlhGs4DF7wtVKe/VECjthWgOSOBfWi/SzE0ljl39vQRM6kZNiD9FpJbiW2
bynbFR1j3cVEmgTlnr3a7xK1jKgkoNXPPkqw/7Iuf7IjD+tAXjUOFSOd1jms//fn
l722yxhhFCmSBXD/ku1qCCaWCoQDGQwP1c+3Mp5BV7mNMlR6cQDZHy+xlVYCMfOK
g5pc4MRYrviIIgGjS7tXmJlHyU41U7zkmO6aLe95YZWYJkz1J3X449OV34SbyX06
WZ0ZfdORbHdps8+zZeIBrHGuLdXh9F6Mk5ogsLqs/6m3Y1aIdBKR1dk2hQfqlZ+n
1Ut48QG3Q2sAKGP23WePhhz0uJtTpGab/sg5/NIokJxvwMOZxX5vTU2aoeZ0jmNw
nRkmppWQ80BF9WLY1otThKq6yvZ6B8xuLM5C7aKyRsiSewO5HU7KYsyaeFFIktRt
8liVvtIbXbgqsxLlzFh4XGxKfuiD5tERNSTAGClEv2BXNBsmCEZGVDul8klevwXa
X4wTCO0Z+Pt7l4wPyVrLfpEaCRPt5y0940J4Kx2NQlU2vUqMvvCguECmIJO7ijS+
aFAks/jIuPPww/ZZehKmtFPWIQ42CY0px4D1FvK8ORCQzaR+VFk+iLEKO/+NwSzS
339DTuRtJOL+9X7FXBlSdaw/RS32+5235bLvFTnMDMIMQbRb7ZxlTd7hkwdlQJJG
FEdoV2S2X31FB+PEZtyXIrgJfpx0n5xtHjYlmpoH+ieEew48EY3DMHrR3NRw4/Ea
D8BGY1My9esdFJhVDPYOF+HTiIL0/7Oj0wUVgx8pPl1A68xxC9ItA4A/JCtk+TTM
s6QIDYyZyXROXxEH0C1JePmpAyD5tChnZHB2Ns8miuPwWzTM4VJJNdOrvcGJGl6Z
mxeyLelaB1UePNROB9TNRitlGQZDcUHFicyVEEDyjjSNlBtpvjQg5qDw7gGnhwiO
e8O5JCJ4egU8+M6vmrPTy/wM9xd0sovLcsC8KjELThsTZHxiMWFFNp9mZcbUaP/o
oIXQBqBe+J5jnaQ/lW08Xl8j1EIDBVO6KecqmdKJOTmBzJEnX64EOXpIx4IwlM3f
ya0uJGN2XnRgPeEgyOUQPfCOlfWwU0bRCOsIZcTzudD/1lO7+LWduM67e1lxQ+LW
jS1ogEsnRtM1rJByB8/07wkIbVsQ/GCQf2Omsf+QqTxyQbPL/T3H/mD/RoRAfgGw
n6LfP+6wXHlMhea44RHBQ5C6Sv4kyDkmNa+ytQdeK+BxsKsb7cHouVbmceZYDdtl
PYDletH/dc2u3x9Db9QcD2CSjFwGR/7UM9FacA5ZbBApNkXiHcsEFkxsqmHYcvS6
VtSnljKp0pHN1swETTAjjGDO68CofblNz7t5lwHz9SGht9foz++0eTPde7D1tGzr
+k383RJOvpEtEtbVWy93HJy3NKJgpDP/D29D+3O17EanJodACYzwVUERaivYykWE
cNmwqRMy/0fnK1yBFsXpM0CN8Q6AJ1xbsiXqLbXloIOmst9JjThHbJsJc4HvQKmb
CgPgNwbBZCg+Gjghk1aarmHgzK+aZ45iYhGnNeNKsF88ZuZhyfTiu1vQTNTuzM2t
lXqXQB8u5SHeLYbJkQm5KQGc89Js1DYLFB3j4rpcybcStXdp49cw8NogczW4SRvV
sgy15ye+YS5A8G6Rhf8oXWeWYWik2OoRCtEuI34t7vYXkeoY71stbSbok8yy8NmI
1USkO4ZSGvOUBbsfLmAVYEqExzII1C+poR01z9I6ImIEctYqSaQ95BjH4XXJ0lLz
a/lXYc9U7nuPh34cMXui4qr9g1tQyzfCadxijUURTfdcJpY7uh0zktyKp39OdgkJ
ykfYC7QU37ZnUaMyBo+UXH6GIV2NbyJfWpnYa5supvrsWv+OedTk+yfwjMXqiG5b
s2ivxh96DyxT1oAb0vCxIOIBgSML/nfUMOWZdm1/xzin9avOuTdGUcM7QoB4fsbA
oD1n8vf6Gb0OVHFq4gNvXQH/e53k0CQ9gt3UY8qEq5+7r/h3KO8jwMiv8otC1lm1
I9ZLCS7uG5GgFGjui3Jw8vxDDF2PYvj1OY74X6CtrgwDdtGLlsCgI+N1DTnc9mU7
/eHB009tsDgW+aMyknYL7yqBQO9HUWIsXI9IGhnIKESz/T1oOW3Ky3XXLsfXQYVi
E8aUGAAottC6TGkkOMOb9Ikv/GbQE5AEwaGi9GZsboav+1mQb20XK3NJbgEjLEuY
BDqQIKKVPlD4n41ZxNVQU1UXHKm8XZkCuaA3sdIyrg4nC8OOvo1yLAEsd7tltt+O
OZ+SoqK1kYDsipINlFpZEO5OB4hQmYUQ/ez7nvJrlp5YWwch7rclA/5DRnRC89De
/xI3Ie6+LAz1Bph5wGSRhL8sIf/rCWktz4N25w1UX1xF1tNsmEJYyx+PGmEdqDTH
Kg5ZUq4xqYt4UbEmfX2ts/35g3kt8/8lTTq9z9fT/PZDCwk2E+DlrTXnB9TK9a9J
VIelb2sFMQhwCL1wb9I9pv8+W4ucuMufURMieF/TBv9w1kkjDuBH4umMHKW7syyf
xcPABKoonJ/PBVET7ze3AccCfh4jPHigy2D7ZRymUsTbRVQov8HrA5R01ub+c5bV
76Wx4s59M0pBNetyGEkYlBxX2y92UUcbpR8wnM9cCAdckV77M4DEjClnWhTHKxje
t8n0v/qkbJ2NXAUMfevY1FR2QetEsI4fnHAckNk/809VrfMDn8pYaHH7uOL1KIWh
mNAAwenZ5lR4mCP9dpGxLm3pLh7CnTmO0QrGGmFEaUqBP0gAbGregYfn3qxUd645
UxEPqH/xuhTxuQhs19BSNkj5D/dXy3GU6ywnHVAKD2betZEg7zL3IYEIVmd0fTx2
lQ+Jcox3a590/hvtJbA/lRHcsQILjLxlwGPYUZz9Jky95hwLjwUTtNloOSbNuS0K
AszUiXyYfI+9GSby28KpGuAX4XDb3wkGKvcFVKJB8Ph060mmu1+LngfY8D8fDiE8
Mp0s6Q8EzZmKwMH9rF+m7FjgVRtYOi0wzgW9kasXKk4AiNiYGNc/eoIlnjoxGvFy
3nVSHruh4E6UnK0UghMGgnhVkVnZ1FkRFkOOxro4Ao6/KMfbfRENRz7wD6xJ2t4E
iRw24P7kImN7FVdHJs/cqF3yB2xuPcpceZdfaALmKTWaite35LPitm0M3DCJKHRo
FHpXx1LLEheeqpa5OcZdP8kVa4Q6EUDHDURcQFc+t+KOVnKY/jadVJltDgkvbbcN
0hd7mfmLuYl8tBKzTlr9VOZIYg1QX1QQDQXkPR/J2c/Yrm+knkjnsmoBiAshhgbY
qE6uyi+EwoaL1a5ABl2TVC5ljgPZeuyumt1yYRBUOhv1rC78Gicxv4CupdMD83kU
OO1uG2nxv2/AR4Tho9aSC1qvBbqiKdFWigcri77OrV8gebwqM25dj0cMAlSphsxP
Kky8xULjib08utnWI/JmKtni6RkVkIYRAJ556jVSdTIfsx7iod1YJiJzHTAVUci8
e5KDOKQDpWFU7nel9bqHhbUM6y6wU6a+oyrogZaR+XX7xnWMjgqB/2yj9oRhZqzV
HoJrvUWJrAVa2kVdJxgbS4RKqJCIkTg2+r1L+dAH8w2kb2FaH0GArTTJgsURmP8R
dUfQqYaaGZn0IMwTUKdTR9qICEDFk5Aiae5Y8mnsl/uepmb+AAqLR60BNHQ2zQ9w
wBankeq1/x2EoaduvHWun+S6lB8OglKtrN988BYHPlNG2LwXptEfYxXWUjQVnZ5/
R6khR9f8/TJwexB0CgY6Nz87Kwq0uztukB3th/htqewq8MhGjhg+wlrmhGHjCkv+
ck2gikx0t2bYwUO5bcNABf1SO2WMxqHqOyL89Qi0SUi/hC5Bi/bBQlSPf0fSHEfb
RJQcu2uB84bV3RYECtYRmW3XgWHDCAmFAZtsMgEZybig2zo5CUnCUHuZZAzf0adX
l21FeR5qFJ2n9Bnuu99VMkCM2xsuqcgP6TEyMifsnJEiC6fIKxnczb1rX+4Bm8fX
ACvSIP2X7EsBxYeDALhF62M00XctLlr5HzUc/hOSg1mPS+TKhS2GDCsc6WEdLVBD
IVkTP8bh5JT5K6ZlCyJrpAnN6LBCkn7Q+5q0+wvLGuG17n5ulfTZ7XdptDMUYwQt
6/zBO+cNatdfZ2pz93Bi6fTRfG7CSwurIiPO9VjAbCRXA2Fmk2K2bWCI9jG9+0E0
xGxasDzl9Hyd6ykoEJQkJoMaBlF4tUf7W4IdtBby5H+oLS9K0zTFKniDtD0mcsRQ
ML9NzmrgOmvheZgqvv/9q/nTh98vMsWRIKVJxF0pVV23zgAeRUIt/0EHk0QuvbA3
nxT8fch92XB5+dmAaIiZ209pdj7Hak72Gq9kMfkRoTnbrICnWc1aJ4haHs0/8yER
0meIKUC2PpSHtcKe2GfgJbDmOJ5lJaiIFB2Sbc3HS3imBsUyzx6oE6X3BwvUN78o
7p7UB/K0jq5Z/EYQA3ot2x1vfY/xmIaEwmjkKg5cVyDFV1QpECUrMfeNLsXF+oT+
Fzf7d9atnUm10rmkuW911PUp4fUML7IoeYBEJm8abRpbVZvJynJaxMyzuAXZqL9n
LD55NZLuoIOaH3RJMowCB9JRqQnSFu7P0e1mSJ/9Yuk3wrAeCpS65Q/rTnALzKVI
DLQMZSfn2QAfFuw8rnX4kMfKmHcMsZm4QSpylgCGI1sPKeeA4vj4mP+vqVBGJhDr
qwtEBb786koioeYG4fS90e5BfksNXjbfwOt+6e2pCv9twgJysQIgAJQG3f34kPxg
QekUPCIVEiuZpt7RgFx3ilTVYjK3exEpAEiGKMCd427vXvAuZziDdeR0napK+dC8
+DBZcRCGj6BU6xPbRDl72WMrakC3ITdo3lkC9dEjceqSNnEPVF3CdjZH1eHSH7eT
ph13sM/gLHX9U/ZBKOz923x8/xFGXz/7bNMspRWUfL4aAbygtARPQwa4VY2IRscm
3YXInotyt3v4bEMuXCTDpNr9arnnPX0mevXy08mv1mhjQ7Rc67vaEDb1A6kzQvDl
pS3xeHzqF1lsrj2KKpYgvrqSQN1AOV0CeCJxFdIm1GvU62luDePuBtL9ui7QaFjs
Sokc2YjY3jBgWeAFcOinkEYXDGwDNxU/Plfql8fNW72AS0FdeYsrgGF0yfCZQGv6
rXI6KaA3+E3Wq7TxQZaxMR6NrGtfGS+Ua3gB7qeH6Tq4MtcE+gLMMWDUCtxGH93U
rZTxFPJTTac1zrzsaBVEJKBFGL8hKWhsSqnPjveh8xN3hyOQTA/haWIGxwcRYBF8
/3uvIlTXJH3/Nni06LR49oBFhnQe7AosIruB/TsbNbEnx8PXaXUqf/k2NjAhnCTF
FW2dTI97KZHISe1abNrjkYRGhNO0r+X9kVdr7WADWSlwD17cKemvcio+idZpl7Df
9R6VWQDmXAEmS3VhaP5+gp8tgXDBFfEp0T/7Nnwhkzi7Y8ovEPLAxVxTLBOQPbga
na+m1PQpHLhBsY/V7NnmEof2L7dPigKwhFvQC+2kcgvDoCQP3PsK5JX44OM8MtWi
lflwWL9T7xuOcEl3ZvFKkp6AMwkY5Atz2JD5Xqh60cmRtdCMRLVSi+aLxeporBgM
J5OYqQiLmzNcFUK8G1AUcRllLfkoR7HUjo81fYzCqwMgbe5c5Cwx8P5RXrtfDBtE
i/3JPpxezZSWkqFUEfbLsP0hbjR0c2mNafsDsrSgaIs95C9DaSSSBkHq6L+Wuqao
OI67ITmvv7+mLXRvev9rAMmLz5PV8IhhWtSENSo3WT8bGZGJantyYg1tYraLPR0r
4NAWmO/2TLW33R9LWMaBwZAV+dkCaXkZicFFaL5JcxXCuiE4kyWTCsp8G0lFrHTF
9lc0RT1KHCU55Rb+P0NaD2zNDia0f+l+WYO26aFdjlR4VvSNp6GwGlP41C9Nr9Jc
ryeGtnN9muVAgjq4M8urmxap2CzPkxommJj5eJeSSJienhfxsbtP98q7dDmh8RU0
T5TpvK2pxs96qQwXFOOAygZ5/r7CHheTs0KnKJ5WsLZ5QEBnMyly5LWEnr9PwBV3
Ijef0wH7HXg+hsQjxHd8XIsZxhdJHrT8HuCstZVKAwrfZII1pdNfKK7TTEYPA5af
Rqr03cnqCqo+GW9+ky2BoIHMhRrSKWIIN2YTMmFZFHJfOzpNMUYCzj679fQbuUqC
SADPOGH9ZVOUBxQ+ihu1QqYkaSgYsXT0Jk4BsoMb17S3tcDoR2K+6LfRqtBUC/HZ
jlfxvw2pQy5rY0wyEJ/9riI7rhEsmGX7gegq2CmHEAQMwPBw7UCKa3ssb51l8680
NQOYzA75W4tzVqKc2MyqT9ECuytmzvT0q3Omx9QFUDU65hhkuMIuC2c2dBSBlBLI
vGlsb2nV4SW/OcSZMe00eadm400pDQtgtcN4hdO7BAA8D1ilUPn5W2YzB5VJ9fLV
csN5WZJ+kLG57MA356ROR2u7yQvo3HXfT7SXk4qT1AppF7FT3FLqzVGrFv2s2vlj
K810x8QDOSSbKeX38T0cGfwLweZBluoM8JaINlCM5grijSNZ9d1YanWalKCV455y
nWPzQl02Rj+U/hvhWmpkexMtc4KXoKc+DutQeePai+odxiQ932YYM5zyDvGrCMU/
v3G+d1IoSREpfCMBiKFIyO2b2AuQI3kyQUxaO5zzlPOWT9UE3YP6TzyHwcBk1Haj
lxc5QvDyBJfTCOVFmwfNm3vUFbIrB0q8Bevr+g0sfkWwMU9gVoiSDcfAcgnuIXn/
ypOuq/lLxij2ksHdgpg9WldWsTeiIkImWiz3bSy6WTbzSEOUSdid3IX+a3/IG/0A
4HuV+E79Yj+WzgcGbCuF3WlMpnnlcY+GmEwNwFrp6LnpMnACW0ctebwOrTQXsddt
aZOyLr4FOKwThDiIK8eYe7IZ+Ynp0nO+OPR4wmIPMnWQ65KbBmH/3UqML9qym2vF
Qx0LTcCFdbs4iz3GUzTUqpSfyqnY5F+UPEeajqRkcN4kj+BCceUMeNwvWdaJb+O6
9qAfN3QwiPFENvgwIpQKgNbJYUbi6DFQSdeXjTFA4M9iDZ/0dhrmKsDOFS3O1m2Z
+RzEr3E16FqvLyuWUG2ibBccCM+G8/rh0r/wcUYqqK9nOl/4nh2HZpRFoPqUSikV
GeiXbmiVByFk4ZUokmqHeWKTX4aumQZ0Z2shIpGSQXe5h9rCPD/hC0TuaqNJBdrz
zcnletKDfCS8ecVcraRyPkYfeTDc1UpYbF2InkHlPmoFhCXC6XrVNz8x/GfAjp4h
1xLDOypQYqc1iZe8bK9FlaRZbDwltn5bAzyGRBb7C/O2jMbhoYd9qS+/iGnH0tn3
efWtDoVvhBMRCKhT0HI17xzE4Oc504jtaw94jFGPT15bAGJ7YAdIFrienzn/Iygn
U/cE7hyRXFiMfd6DRPQZO3yxshWLFaQ6z26TpZEaKud6qw73T9Wh4waghe7lj1tN
d4nOC7ROrtMx9Z5W8E83s1mVP3Eu+Xyv6tKqpJy2xu9cfgo3AuZa2iKrqE+B78bQ
UrKeDXdeJZwSNbycpmoECQOp6nc+5IwZfx2WbtvAeij7HSGFpPIN18bGHQfw6/qR
KEtNZSU1OOBt6gsCZ53BK1MNdWxx+IzxSNPfXmH6DVGGA3VA8botfaZk18YAgfyP
dFXxORjpWBUff/6YNicETAbzyUO9c1fQSMBaJg+wHTsUHiyLGsDGRWUXWU09/SsN
KRyYytp3NMABbfpPEdpX2lGGgGiB61pCav03URLAFMmKTsCS0g3nDaqf1IgCrH1R
VvIEY1zKfqGmkdL0o8LJxGDBiydW7btUl0qsjcPVtHS09KqNBEj6g5ajFzQXsqZT
g3VC6RieM+j1ETI38k8uk8vKqf5Z08T+/MsJyYZNHfv9VBbmiZTMBpfNRqosyD0G
36jpFenX4aLWQUA+ovYmxsqsodLveLxGUMeqtFv/BcA/UYJktLiw37/iSmQaOrjx
EAVHnzKhEp3Fk2P19MjrWYJPZOAqd15K0wArnVbtMw1Du+IqXjuoQi9FdIofYp7m
dUHp8Ofw5Gh6oFMTuDWOIC5c4GjUU0Iv1iJZ+t7rwRh4ugDv/UFDsmTJ8Aj2E/OE
yx+OmiTqReVfW8aRG989kgyOfA8G5uxVU1iTKu37pE+Jv+inTBODX/zL/Bv9B4tN
EkXD8fRG4Cnx1e+O2BiTcami48aVqUVY9pWFps9ajTv/RkzADqAK/of/JoHQS/1g
jBxZgc4LM4mSJzhCqP/Fp+mhBV8ekJ5hOsjKu8b/zvC2/7mmSJBx3PQBhqnXNr2+
ssZ6ID6VMjedcSlSnShinHiMxHr5SXE8eKM31+zb5pLLB0raxo4WFssdooAucOsS
8uFgz+v+Xu3O4tqZEC/xVHXyoBgePArdvBVxkRCSTcwbK7o63wruZdzfefuOXSPg
/l0iX2pFvjG6mqDLTaEPMXx925iCPr5PKykaFtmrLYQYIcSi8jI273+uHr/oUjWD
zkw5WtzlQb0brvDE4667iLO7jKZ11e8irPG7o4GuXzOZUBP//PqvNQ3iOhdSrfpq
cmmnFQmZLshByaI6I393DQdLHjo0vQKo2jlOsat7Ov5iZD9nsu8lBsCR5RtSzx+h
k+GXvUB/N/jgzFb8bD9hvzpZmoS3XmcLCk/dSnQLgSiwld/6bbePK1DmMZmlOTbB
BGm9J7zLV8jW3yFlTiqUSpeOHL78LclkjY2lCaTT99YYnjRd5m2M1beQm4s7J0+Q
ZZ3xsaRRqj0kYMZvA7FPefxyx2ZGBFhAzTuiZd3/KzBsh6AxdDQrthxFfkScMCHH
gLoPVReTUwgce/dpyRqf0ua/vSybqrR3ste3pMq6i4U6x4l2irTxMf9xNGqLLXhR
pIa3/ppR+en1iT//bLw/avG+Ne7oVT7GB24A1m6k4Z4kyDxnP76gZ/RxKz+F8CTz
HpqHY7naS9wz/giNIk2y4mAjFo3+1Cb3TBtGcbD7S/IE6p6HCEIXlKspP4aWN3Jk
szAq1WNGqVY/25mO2tu7MGnoAEAZti5jCff0m7Nxyb23chsuUASHNsS6TAXb4YJp
fe2Lny/l00//3Fp+SlXDyIjJ9IPzhxjoMd4o/vl8biYxJpsE2FDqQ9LUKkEvJnG0
EVOY74OE2cn5WQSxAYQ4rsu+DQbiFRP3MQqqUI7pWWDEtymf82E9KucRR9fdimKi
HEdEZYSpYPyFYwmKtgRiMgPYSSzkG/zi2sK/x5oyI0wXBdJA18ud6Wuqbb2/oQck
mVahqqiHTG2iwCRovjfCzyjOM5ZvvDShl/qY8t7MitnOa0OlxM11Fzwcr+qSew9y
oQH4p/Ho16uHO3p1UHFlNZ6wOmekGWpZ60vVg9KH1jyT4MTMkbFGi57gs4W1oTST
ky4cNqPDoVSc9nSQWwrKMdsdoMxdOO/Ztz24Rp3EfIOm4KKjd/K0E5wFULQwlxuT
s+BvYk3vLbLo3rhayUIviscpPv/8zGaNGPiOKXGYNb44/qx5X8PU5mNpg0HAIfmY
3WUVF86phFDi7dw9WA7nSAr6IcTwVaQKeGfllRLgONS+inqPLlJhsyiLuWROIflk
3n78c1b3Bt/Umfs9FMYJSPavZL5hxw6Nui7ugjYsmooi+ghiScufe6Z7Ue3LA925
x0mz2Pxyh8ljShnPEXKemRpzOMMlPOe2KcWeI4R9s7xzcf2tIo8sK90O/h74z2un
gbWVBztQYATZsR72iKQlB6bqWpebnHD1BphkKwW2gckH/feTvYJNhO1phahkTW4I
Eqz4vNdkcZuSP3gl5w2HKajUMHNQbArMxqY/vZyShtixzsREoiH310XwSE7V78NL
z/K59JQIq4rT8AB9yONTm0QWR7ysFReRE/j5i1zhGQwGcf8ZDM2z5fCBJLLZVxPG
zdH0wUCiySrHJ6Cdo+bjQ6th6RSCtmZB9tVnHeTTaoEkacDw8ukQSDf5DQ2Lqu18
F8Ny8lBvhWnpIHYlFEWzFb4KUpPlRTUasDpt2PPdyhMmfFyBzOtWqbm/aI4lEFr7
k/9fpT7qgiqZPWuGrodPjf5yC8n1LhdonQHU31Iuz+IpNZPiS2HntTHQc3JkN6Q+
uaIdMfcFtGT+cE2cB86aDAJQwQMSX/T4Yzn8msmrSyagULGz2pyZs52g80t9tdIR
gfClAxqgkzrSAhDWQhFbfsGN7IRTxx7sESip89PTvWsjBwwAwBDPlWF88ZJtbhpm
ouSQBQ1s43rm6FwN2K3S6GlysvyWTSqHEFx+G0zZi89QXQYVhY5CM83eFQ2xqCp9
Hn5yz1e7rgjjMH9zp09Wruq6ivDs0Rwqfa3X9IEYUwmeOmSTPvEejGy9ioi3Ca0l
b+LOMy3XCcJh+7r+wlwwaPzN25KtXvI4RNtcur4FeyD2Rbw6VL/vwB4StEln9bSe
WA/eaajH/lL+G7K1wHc8CB3VC5E8OGTh3cARPnkVXZcvMp5P56PyVakNKUtoDkvC
6FD2/2ok/nNdxfOsVcc6B1Z3nLnKAOQpwJ2zcizT8aWRCWCJFvC/RLFfNuF2AK+O
62FNrwjYuTqx27LXATTGaM/pmSGd26m1UujPObFEChii/018bRLLUGITdKrrljtf
59tNxXwNEolMBjJ5RLM0XHqsIj7HdVb1tTPdNkJnM81N4FuFAE9fMfmQ+EGoDCkK
A1t90TTlm5Fp+Rlpi70E9VhDgXIAwGJuiQfyzCOZbapKRVDiOCigrHp03Rn2IHlr
6JdLILweWXfNN/Du3JC9C6TDRT7TY+etEz3YZ7ShzCwS9Ffuatcnqc9yf6yo0k7+
qjgiJHUu4azZHPe8+FBmVup6x94yR464iUls6IeLZBKedpwcssDJO0T7v2U+vbcD
4aY8Flh/udDxeq5ry7o80yPDU3dvDbeKhwH17bQpefVzHwjobJRYx/kqlCWaDABh
jyGBiBVuPwIu4tJdUHNVrNBiULjgUNUxIB7iZL1YPzGogU685QRTfeHfQBd7BH6v
BN5uig8EzBxVwTSOrCize87DTyxSxkP5vmxeBR3Ca1JHIA36GWOA6W0hVsR4TgZ8
K/jWLRSoj2sl5zvGycIx+IOYFGplNvSv9e/p3W5cqok410kWrWQwKJgYsv1BhkjO
J7783V4f2ylhkLfQ4lAkiR9PFmkjbYt6OJ1J56MOHF6Q20t/tX+tVfgL4GFjUvZ4
cq3aQQnJysTN0S2A0IwuoLrdFojDhFVdK7Lrv3nPhjceEz3LYRMJe7Xkw8uAFfgY
M6KJdpX/OmVo+ukyNB26q3kSB3DZpan0q+ndyjSF/87Ee2GakkAZ419/aswMTf1Y
MYw0udPdUjiQY8hKQQctBRsBrP/zDiIDRF+fpJI8Y0lbC79m0qYZcpI4vw8bYwVK
JteA1ak14WoSCXVyWgEZKn5CEJVU12Ns/mnCBzF+sJKhPwmLUv7TxSlsPv5Wlgs8
lvkIPQ/1L+1S97akqFfT2BCzlzVW7kmMWNKcIyRk+osAFQk519gChrdU0X/KVf6j
+S7nJVRoxlqJnEr2msdy6h0xIg5ummoy1ZoTsBf9a9hDPWyC/eOc6au52sqvLr4T
Hogua+F5L1P96+NzBuJ20Yvw2TsmCGmfAwxEf2iA2VL43iC2s0/xn5vXu5G042bx
YUEKidANMdsERRZUNM5jtjnypZPAmGYNSJelgl1TqSE0MWgey/a4yRLWhleJOjcx
Ioe/A38CNfCq4Ku8vJAB1kgxb8THZdkeMjDWF41n7nDBagx2KrliPBIVTFlqlhjy
MNywcy0GWgBBF07USanvnd6FZfYygvg6kpxNQPS0NiVV39kxCqQhCP1zxyPs4S16
PTdWFBH2dCj+sVgahrbgXPrz84kw0qQQzKnsbg7YHqlaEwWzQDG6dogQQwCP/N2N
JebgFpO79tg238Xny+f8GYLIBKcbL+toJym8w/hU/cva6UNf6v+DI/xk20F0yz8k
8ogqRSvzY8mszjoTTHPXyLemcgpJlpwP8R1iJxifQ/xxtpy3wcpTHCUYrGV6I+cU
xfppr/Zwhb8by0eW+t3MSOClZos0WUQt/L8kHCGs9pgfeRvrKC9kG5lFNyoG4RF6
XQl7YQOsnaZ+/ozKW10/AUEDu23utbQkEb2P20t81KEZiKc+xMNX+gfpIQ9JTYf8
EOgZd+0+MPxaTBjnetwa83p0aERqrE3yHQUsA0taVQaHL4PZh+YLXxb1DDhcCBjt
/EdsgS99f4YwWYqT8yV8/TNOMt1PLpHUPYB6g1o2V5Vi2USUSZgW2SRXfsBr8mFe
u6eUjKp8Mh0o6MX3VP1R0HUHxr+B2ZygxS3ErFX8OaC9E+GS4Y6+8ri6NSK+jK8W
eFpgHwoBp0Nciga9bRUkY1YXpqw1gz/1hfWELs6ne7wxbbELzKCU1LMsBflCCdNz
Ml04VJEi8H9VTSBZlTpatkEhzFLA5ydmCCHgbdVAc3JKj1NdFxVllE+rPhr6HQkY
mvxGsP1edj2OITV5ocGeYmVI6AinKWWTdjGLI+5uvT+Jszd+NYyzopH4erCwMPc+
6f4r6d0eT4/D51RlrSyWrQCt2xNfQKBaLsE7KA7f1KTuY/J9EtjOBHZxI3oyyKSX
ddYArPUwGQHIS+S7FxqzP2RQEvLB+o2KQ/SxeMaT7hIzYE1/rh2iqmOTWL0FxTuO
Uq27ltS4PFBgDGDopWQQNKDvs2Ym8i0RVkbcLVlVX8nahf5l77e2YSf2FW37hYwj
8pEcTc0D+qTUPF4xcOBpRu6tML/q01ZqxFtb7lki2VzF73ySfRkocMkH2WCoPmWj
It4E7hQhqakj0MyDCjBaPdwtVB6qQxcRZLc6fOtuhV28khOT8AG8TRzNfq2tvCrX
rRsx6AYDmPoIUyoPmW2Y7Os0CT0zAlV75ll6eHcYIvXk4Or2L8ptYv42HLbNtsEm
U23fQGeKzdsgnlsDtiv9L5LJjjaAg6JAvXU9EjxnYZRGt4rMop/GJ/p36ivuaJAA
33JfLw9u0U7N0wZne5FILCyMHgBJ3iVIT7JHVCGJbJD0AVQA/fpkic+a1Ow1O7dp
FO1TEsvBhk1EOKQbVrI092q1G4nYaqAxpGwYum6x/pG2ovLLTyY1Rnskf/2rQADw
p5QLqyx7SBAKDjfMNmLAueFWlOpImOCnclLMy4sK0l+x2KVxrAlY9JIz0patyOmt
uIFsdfF/c+dVtAkgRYf5dV3qUJHV424TMXmGswturvWRIZfnvL9Ok+bw0/XfK8TB
pp2WeiW1ixf7O8uZS9My5dtSdunII4dwhilHzqoK4Cc+ZJOnQTWHK0Ud8Wuug1JN
O94fB8Lo80c1S0oJQftYetcUxxz8IzJEysFP+GnCNY7nAYMy6Ibf9MDtvHo35xGA
QBpJlhbhm+ppDdHAfNfKoxJBEbqBPHf091eTZxN4rHYf7By6THU9ZYiR+KRMU7CR
jwbqbLJE/I0A1fnPGYfRTMqQXZ2pNsFysgmTUOeI65Grgr5fW5CuSkgOd1GBTiog
CAYhAJSJSr5OAM6KMIJqYWVaOngC26qgrJoIa7gZyPl1Tf4KkTCLgpg0jl+En85r
nUJ+QXBUCq2+fXnxvcdfd/LWmSpV/hufzUAq7+7dTV8J+FVBv1PvScEM+JI4IX/1
sVicGbO86YKxX2H83ObPduqKLkFiiCE2MR4/JEmSWhPWU8UJ/AM3hP0O2/cpMx5r
dZn0c0lHV2/+IfF/p3Ddsn7Ax3yoiAj9dnX1N6DHVfm5tSVQEuwn63XgEQYb91A1
Ht0K7gs3nUsiIbKe6khDqfQO8sbMGwvKbl6zpxYSSq9w7EXbj2KF9nh5xszGCeQx
lTv4rJ6zOYSpHuWlYfTQnrQIIRpB81Kuv0ScQrolbva90p7iXdU97RhO3WZxQj1y
tJ3259uB7hvIxakNlhvTVGX9JTWFsLnNiS6OWYM13P65IqWcT1/4TvJHMjuA9nuS
emdC78CeBeGnd+xvtfJIiW9MthYZpdT0E/tX/nidtHKjGZoRILb/kY8Qqy70RW9Z
8bIrY0C5uEpF3TLiv6MGdR8wAyR/qhES5XN3ivlbiWr16gYkwo1AwGIeRe4YtyCk
WaTCHYV+qwQ+/Q6qfyA1Kfs0umwgy+1xAAtiZ7L28f0e5FD2LJzu0ZuX0D1LyoTL
Ol29hPqLWKblLkKHPvRBExQSCYf9qqBlfXy4k8TI3MJQdaI+3dBOaKro4bY0FaWM
9HlF9TiTFf5czNPKmNa3gfFOQ6kw0H6hnsoT55POXMAB+PPwDp9VTuhpUFvMzVsW
hJ7OmzC70JSNnMRDt0/uBOeLElu8coTog2JlK1UjA+fIRJw/fFbGIqcc4CwM5IcS
cI0H003e8NGcwT+a2gjJNS3DyyUtXKeCxeagEvojSCDjD3R4cgSv3041ZTEuCrBb
UXJXHHrYRWHVnRWB6ATwot24VkJc0Gzpq2B9VyANX+oIHZ8hbLJV/VfqBp3lPm6g
zwVJlcwCyuPXtQUa2X5/2o35qs/CTi59mQWozgEv11PWbxpj7qIvoLG83UCAR4Ac
tpX1JrU0GjScP7Gm+myzpbcLAtKVtadaFSn7A3XvuGyGDOJzk08AxzJor5+bjeoA
aDDWeOSvj/SsVHLwx2Yn11JJV0zi8v0tr/OYp7wvT6pC/bIxHb86Mm7ACKaoKi7q
bOHOTrl7p3WUmpWfLbnouoHxR29qkda4zaWJgBSUJizPzGuCHwgSOz3zeSqloSZQ
b9uv0Pq3zESH/w7rFECzjh0CmDsxwa0Vv3iDMwOjQcWRHZaqzIRPJIuF7+BiEY2W
myglGlPX8p/NsOfati6dIXquvz7Fb1ByFIVKMerEQuIh+V5JiTnxCRAvjV02KGLp
TgSsMwxMyId411zhfHgPDW+TvyYiqLgJc416123LxWsZUmoY+akspr2LHRFFTgMB
v6AeWrc961Esm/LUfT4vMbBN52Z0rc1PQPqSDbTdZT4WEL628jFYYMyfuQfU629Q
CAJaAqPUiTCYYUlUQPTpPWNROUgXnBUbra4SKom8Qrv3F00Ud81EruCHHs6CaIa4
8UUBHxz9K3w/ACew4KiMg7p0mnt9Y7BXM+6zBcs3JL2zG4mKhq2X6JSazDULkuLp
6WpsoLNUmFVXHlzOATwTakGa5i3VEM37oroBf5fPOzLT4BonWmbAF2LJXZmuqOJn
6B4ex0Yq2LoR1ClaqnfLSZBJlRihtuWB4T+yOMLAMj4NXO29lvrmgYQU01S/hbyq
Xv9JMSSAj3AeQLmZ8CyPKqf/tALxgGWk4yRlup0swI1A50zwIn8vP8woiKDAdtI9
0BHDdgcios+4EkqCOJipocl19X9+ImoSO9NYrQkipwzoup3K3CqDryvTbEPoiFVA
hGvMNJ3G0opCQG0Tz3wrfjP2GTkmhgoJQS4UG24ts0sKWcA+nNOxI8uLSjQKmWW+
VkfssIA5rmUBPSIZnQXy7ep5CGl85K26ww+W3kOQOy+2+sTyduAIGLht4bRcgeIq
K5ag7Kl17RDoR9tnb8wBmQwf7B/OLUfl2cBIG+d6L+/Nrvj6OVgQVTSrZQNZ2DfD
obeZJPyEo632vdS1sIZ4rh1VjymouOa4JoSWLoOF7VRJKKEKw/j7g43mfNK1U/tp
57a4uyf0HYo5taYgAMTRFApwQX2BHO24JWnzvvNVhHvG8ju3/QOaG5VaLcZybrAL
tz9kN6PndyQ2/OA5c9RjaMO32MUCtXKB72vTZ/mw/OeCcSfzWkQ94sFtQIKlrwET
xhVHCCg0LgXZb7+Plf+PAaReY2f6kxX57sTBaSjbZzqI1Fs7v0hnBAhhLPuA8nRl
kAesJvgWtjdW9oI3kUSYmrL/RK5y296iww40iG9BlOXtBx9NMD5x1keV/SxGJg8S
3gsNnv4G6vCOkiqKjABm9aRm7D6XvvaWiEwP8RVNwL/ndlI7pjcU47zM3fbLS1fL
YBWX6w7aFwEJ7JhXXuHhHjFyhqOA5wEhL11V4wX7F+dGPSJ9dVNuEIVQWwk5eCmQ
6XuH66MI9iKbQZFEWTAg3Ve3UrZWIgzQaMOF1V/ytCT+TMMvSOlbK6s727c5MYCS
EEsrno+GlHJq4jTJy6gGdH3XHpsHkFsBhDsHSb1hwz+Rg8C0bkdjQ50Zo4Xls+YN
FhATQcg/3f3/NzieHPNkoCX+72o8CUuQoVaihb77Tbgx3hQ6QbVrcDiYDRurmNr/
Kfk0mcTIhSJfhN4vpZ7XyS3jY2wi/Z4vBZaumh0EWJTXgi6fffk6/6pqvOuIU5c6
/bWWyZypegmMnTWVbmNGGkWvAiNByndwpk0Z5z1vVADVIJ8HQn0WomL+1tUbLn6q
Cyvi2JPJeeM1MV1X5EkygT9hjqK4J5ZvQjxBf2RxlpmLxKn8Mt8X0vyk1LRfgUcb
uYFPYBHiAkXgv4mK+1xh11qmRqyfjm+Cm/ydgZpshrBIG/O/d3vMTqNyA+SUzN0u
qwaRpPafEN7kfVBjxjletV7aDIS0feqMVrsWbwTNHp3DdnCLJ7yeaGFK95oiBnSO
16ENO1Z4PElQxJBwzOEgKdOBFzwCmbtWY4vPmdpwyvTgjhtFEmiv63ygMNswtGWS
sijtswZKVWj49y443G/AGawi1DNcldXV3Li16kkZbEfcOfl9jy3QJYAFgb2L8p6Q
KBieGmiAXVxlk/RTPNxUoAv3bHfslaUAdin8R9HYT/WVc0G0J0PJeG4Gqm/gqNnn
wjqf+QHXQGZf2DHfbP2H3Mxx9wo9365I79YfskrZl/dQGqpLab1exMbIrtAjWaEN
6rh41ofA+Ll7ZjvAYdKXfj/QIzW6iK3qVMC/E3aYYyPzhn0rJwAgtoQyh7PrCtxs
d1PoWv07UfuJyvX83g1kfBRnEwxRY4quW0BD+CFdxbUuZDHow9Jtm1xzTFIFJldA
cKqxmqTvaWSgUaXgVEytaI0g7HuE7tuUPrbBpqICV6k2AeKoDyZss1hGCAlRK6Dh
nDJmnZR9/5IxdOjOxAuue3jPQ6FrXcZAkRnnqJTi9R7Glf9AtBwjUsb7Y13XxIQY
+w1Q5rWtNwo1ACUHfMEXl6WWCJTcLHhiX3Az0U+294jnwjOBXEuRavESW3BqulQy
zeXoU16odERI+judTOwoUQJQ7yROhIuAZWof/fUSLZFCqznvXwDokr23gFPJECNF
nVqqxDKQB4JXesVkjVzNzH6wMc7EVJEAM/MIsF1iniqLJt/ucHVz/g50lwPxid7z
pMdQ+tDGOkICVkPbNMmsafyIyz0iu0LrO6QIvzFxELoI+BHdCnHLGwVyXUvdza4b
jJUkVBb6k5sIE1r+6q0P1merboakgO4L5FyxDp0uWlSJUz9mwfQl29fF9VvdiwU0
zoZttigUJehz/QbL4P4PPea+76JYyYwFVn08V+q9trgSKsh81gwrJGZUwCycUM7c
lMIiIMowqHxjxM7Jj3Q2T1IoFfo2sKPH0mb7lBlPKOJZ6aIdwowJteA14OH9k2se
VSoMy7du8ER0Gmo+HrpiDUIHoTq/2yF7lIPD2NECoF9Jd6lKe3Mk9d8HHk7gZTDF
IrzfwqgCSsLZfXBohUmJcHcMHDcR3rczoXMrYn1QxOW1vKS4IcanMERXQdh/bxEt
jOtNMVyTvgXdEiHOM22a5hlsavWY/K96AG/8Ts/g3njGqGfkitB/SM3VW8OnpV+h
ZsSxszzkgGzd1WfoyE26iQif4GSYYF3Ip2FXjIUlJK6WMyaSB4gatECGcOG2TItQ
oEz7Rkmo1DSTTYKqneVTBttXLc0i1+ux++LZhhJFdCeCuTu8JD59R1Q11RytJvXj
H0+It8KrzaKfpvVcy+iEXARWa6AVJ+UjZRAUTm1c5tJbYVMVij1PNl7B6QGauwPN
ysWA113nzRRzM95j/07A+N649zmeTvoCTRW0m0R8EQsKrsB7Kjp1a2/sNHod6CLl
v7eUazSxSX1x7HiUVq5zqypOJhEJ9gZisiN0VVPboD5b3lO05D5USEk48CTlSidS
cSHI8r3ZapJpOBRh/uJY6GsX+2m5UH17cbW1f/8zBvtFYCWSXb6ORTKYId6qmMb3
1rRDfqBqAWc+uuiVF+wIePdyhMPAWHtoKGzkEZn+IQFycWB3rK01Wo8XByEBq6qb
arQeI+BhZYaHr/0cx9EofH+PxLo5hReRlILFi3TW3Z1jt0xnEujYNwpYgYs/okfJ
E8wKMVUZYo9eadWD7BzqAidsBxwN5ka2L0qX8JKV12+mWjPMLF6LX1mH6O98ItD2
K2mx5T9OA5qoK/MUeS032V0ZrI0O7XssR+N1nD4WTSj19J7ugCxEogWBxqQypp77
Az7u1oJEgXZYPNdNUGRmAp+J642bs5Q3bXKbAK4OlDVvU0DiIirj5a4Abx01Ks7q
1MRp3KmWa0Y80lW6L7wts6YiS+Y0bcK6eC9+sAMAS6g2kz/6ofG8MjQN9tmXmcfD
DFo0oqOil1c3o9T/yTaTwNGxjuOZVu1yne7Cc7wPKmQjyTmo8xG2jNULAujLMp7t
9jxHiw/oeBXl+eeFGGQcbfuexIK4etKsM5cKRK737ocqajw6fq+3J8W5m5HZ5HlG
4C7mUq9/zZwVkYh4rg9Bc/pT9L8tn2FOfNCvLecMV/AJYfpc1TFScd/o4OjpU2xM
iA0nGybePbAEDk2eczPAixo/Crtfk5IYl4eMh8MDKGQVrmlF3Krfs0gIl6ZZ60Fy
tEuOT2n5exvqFpu3kVSJauurxfLJO/pGVSf1FpXv+q2ixSk74rcBUSKkr3YIxzn6
YuQuBNrs3T5W/yGNS4qNF01qGpDcTft/ATYuxZE/DO3K2T8xr6DzdLFSjxJ/5pKA
gdxQp/1de6UlZME/NIOPxZcX3ue5mHtOIISFoMTFS3OMtUKF/awqqQhsKIPUtv9D
TAH/BoFyeyOSdu8FHqqYy/f+TkSZQcqTgkoEWh7vhlHYJzyHXL8hs4UCpQE52eZy
rgHxwAYhEufv80h5Vz6MQyTNBhZS/e1qFHPRnv+G+97F08V4gEwF7I/29eE5NDMg
X+V5KPE/lxOpinJFD0okX5DpfoucEBfI8a53NhklpV47dk1FmIsopnZN4FJMO8KN
fuc1sUPZPrzy/e6h6sbGJzz8HVN+oqbtVQPLuA6xd6gMlZHyQqcygiTW/+fkBcjJ
Rbq+8yRn8JpkAo1HyOzLIRK3DrKbYqwhnt8pMQCuWGxPiq+CktGYMvFX9pLI3KhD
J2JSSafIIHcs4jg5GDpyZ2c1i7m1vMjzeQrcBkpuZ/6YuW+NiJaxzQ+KKlGfAOzG
7THEsgq1GInHZhOc2uyTZi4CIduJYQOUnDumummgfzGpi68rpoXujxMjMrVQ6eW/
eh55U0YR8/uTQVpUSRUOQRL1YeHgyIoqN/uqQotWWTg3cJ60Q5FC8IcOzB0E5cyq
lOsICB3ulBX+h3dMKjUeh/AJGx57c7TE+Oj/OxeA3+6VQfjjhBvY4icYSlrFkONr
8khS8psf4f3zPOa0DpgMcHR7NfeVJ7xTAucBWRQ8xTYVg98WGfg4hTLXC7BxuaaY
Pqa8l8hCjVlcyVOZXCLRkp1GoOZucPS5NOgEJ7OXC4tPJc7MeMRx/CjJSTAeSFPQ
C1I8Y3hzHnP954tRafneii1SucC5BKHEbHqpGEvS5GUWv59e8VkgTCioiNvhdVTi
Sgd3UjstDOVsJKIj8qBmAeLd5wjCD+JnlNp7i36ChBWaATgn4A6XAfVtxdcdH0fX
6nsHvdX38TZ5/+m+4I0R5f4GwZ0mnVcp8h5/gGvy1UxB59y6BX1AvvKicttQuiTw
pOJ4oVDrtGaasqXiaO2IfNSzkfJuu1AXf3IvgJb9B7KHx7Wvg2VITFwK2GjGe21s
BF0A62vTyo1/gORKgpOWWm16ojUK32DBq4Lo7PzAu+jvC7B6BWlWEwob97AdXooW
mvEZ9X8aPYIojMgJiUe6ZQVN+JPpBNjpk3cO6GbcUhQA2pa6ntBrKKXeRRolyXpb
cIwHztCR22S6eDHQfJnzpVO+k6S5vCWHDHWMqNKXGkIbjyZR1ZkTC02rEDaA8dMZ
NV6HLVU/LCo1MhcFg46fggGPQBkILSB7wTa/dL5aIqQ+IYvSs2tcBieD0m1jakux
fizvs7w8q3Fy9WS2a1oSnxJRPyhzBDrhb76YTUSdb+5HL9yvhIDFV6gADsgyZiOj
Q5eW/CymOf8QCI+5DKvRxlph5p2IFNlMhE+9ya4GGv8iwTUQHtcH/2p7qMO5sSDl
VG1hsEXVCKd4abyE/MtZiLHy8pgQL5H3RrNrYtY2aJ5W3aVABNBtZ/6yWZzKsUxa
lQm+6vBTDARKo88KxyuBoW+pWIPmkCa3duTLMFOAQgWaaMh0l1F+rBTWKhrRZhWN
sbtizmk8sIdY8hXSWH0TL3FQu7Hb4ZqUg7gts7tArgd97rHcOZL7G09cZ22Hl7SX
9TsseSvWpN3gV9wTjPbk+LKZmhHkiwy1Xp47OyOek+gxfurN9I+Z5oA07m0BcWJg
ey0M9LqaDq8sLwhwUbW16jbYH38zv76opf3Is8IGeHuI+lbYzwSpdttc7qvKQ2XZ
zhmiZoHX0rmxTafpmSLT9npHxyn9rD2jscxYHNEkt+zCWBgXooz0tlCRFi+LbDcN
rAt5DM84MQwBPiJPeIJP91LXaR/PGnSAP0p9qYEZRIHO7HgMdinx9pxB25hihlxH
3eVulpQ9Z+5MHuRili3cT0kax4WDoDVv5Jj+l9GpX6VlrqmOgQts5zo+bg+gxlVT
9D7ZzKLwiNM0TyYeWutKdya7ULoa8r3CoDLRtoqHgTZ8e3ihMFr9jdpaVqorp7ut
zRoBhEJ/x8fj9jOtdjKO5psL7HlB0CIwF503XjiUavb7kAFVVm2xzJeNI1w0DYWV
mBXPaVtdY1uhN1odSXMtOb2GPfF7n+nvj+xD1JbveEtEmDAa4f/QTv8fyl5Md4yJ
bGS2oR8Uz9FRqfXNh3bd8lhoTnXqE6fc8s/a67SKt+92IRSNb5cRswKx04FDTSqs
1OXLyJk5+VGMhpCz6mgtVXU80NBzfgAgOcu5BKYNYnOI1fPBOJ3cwCOywOji29N0
3Z7YQGCZyXM72xvKpONwBU9aYlV3RIXya/ZvwvCfmZZ+wGXWQjrJQC12rDIdfXqz
d49n/88yY5qcCHfVbyiHC+K/tGusPvWGT3HcutRPxLI05DctW7+QSLywzNBZI0Oa
pw0tRUqP70z83Fl5p53jGuT5eKuKyVEazEALC6G3JMg/QO5EOj6lIEHR1ksFSXel
JafS801DkMGhDoSr/MO63nKIvwebG0s8ibCY5MfsoAY0X+78+Fx3aOcW0EwngLBD
HTRwUlc2cEyerPU+668wihqPTysR0G+bBf8gKCBmsjlL2PqwY53RzxxsxxK2F+ss
GxSqqN4qiUXIAVnB33tjOejt5aW5R9exmfyD7715bPnV8Fh6I2DbsVOAMOQQcm/H
uHBT3sB12+Z7RvI3UztsMo2WkMP49LdgSsKPOrK3xPoHUWkab8iMaJvitujrjgkP
NJLgLLpxz055ulON8pv6m41P7lhLKjEfMvvXbSQvUHE8PDi3zEBW4IKOMwBbEbKW
j6FiqC5hGkoN5Y5LzvqPQlLgY/vLkex71tM7fh/5Noy8VNm+18ld0R4NLK6vl4YL
+HfHD1DE4ORZIQg3LKVsPi7bIvx28zaL2E62MrCii+74IgRLZv4Si0qv8sWlQ4tx
YRCb4ustzRrertBOKTXmwQcHL1E+LpcWpXiwGl6Wsq5XxK5jfHArKy3SUVNYHunt
1BQrjXV6L6yAyTZ2zH+YQ8kDOojdxDHyyGwcpEaRxSXRdOhXz3xAfzSwqtUZYiIH
6jo0L+3Td1PcDMtzmfME0tXBhhvywujRRbY9Qp7vWG0XcgWC2ZTPDaUa5lxtxBhq
9mJyoyKZN2QQvPbkBXdZefLxDoH0R3Z+2HbdWA/fxCzF668OvuhFRq+so2HY5uTw
FtcQ9iMx8Rb4WJFsuHo68GZ0pEKhjoinKI63NEbO3uUS/dxl9j+JF0jF7kUo0Vio
HNoOZd9eYs2rdhGCeJVSP7JKRVzyhuIayqdihbRfJwMNfDX2THI0+oSPR+x5BOas
LhCw6kzJmlP0S0wApAW5eo2SDKYPlG9tspHqGmcI2todd6I8YqL5/6ShBUxdKsIs
PDyS+lnrVJnUvU8fHnl7AHC2IFHXGZd2f273Fvmfyn4VRcXztYGpsWPW7nnn4Fcg
cRGSmoNCL6KNXpSECHsHlRPANiLMr0EbpU4ZLXkNDsjoBYvfJHs4znaSaXwUuIn5
hfH98Kqc/y9DiFEHOrgBVIHyoxlTeMJ9hQRxPmlonLWKm1QLYjEmq1h6pnx2g/bX
zVTRHSHe8OZBlk2KcDP3EBqaNI2NexrTZkyjH9iirWSxHcqnEsnhltMLsKA4dZai
s5NvCZPseUpK1m8/FywrK36fTcAOgT8WTWhWPBWXbOulJ8mzIrVA3zBI78vivNQX
puwwWdDQXyBysQWcOLHnoenqIt/TEMJN0dx59Oc6v+HhOAxzpVrY9GnK/9aV+0Ph
EcNa5yjxDnlzZCbXLnz8aZnzETjlAfuLIhq6bvuulBcfsJ+4pY6KgztUaSn6AkzS
av7JlwteJQiOKKD+Svmm/sgDZF+lUOEBL1+G3TRpQol9O0I8Cqrqnl4iLHrPgX33
c5YIOXYNWQMd8lx2BjyuFS4jDBLFTDy+LT8dsG6zcTyJabnTNGgEHAn/e7Uuw7oR
FiTWIr8+21nECKN53QWC+e8fy25opjNhYzHoIi8KZafDzTH4XQ3uETrIHkwzSNLf
gliA1aNq2gjrlPYAl/ibJwW5ksP5mz0LlEK3q3tU2TwWbqmw/8K2usHxVBP25aCB
VPVT0NFDSJxrXViiBPQoBSoCRA9eNwNf2eK1kgbgc99FiISZm9+D9i16Ra1IZfWF
qSFXh66e17JiYrk9/VtYj3pBcNf434HMEYlw2M0kY/wtx4d/p9zrx1Na7df9t9qD
OXAnqClsEW4oMH7BZHxLucvskMMW7r8VBRQrBt1Dxf78QGxoCUMu3zKV6uu00GYF
isGmKiO0G7Tu4UuevB/cMG9rnpG0rHsfQpRondQHEtJJdoXsIYyEpGHbki0/7CwI
6iVEysdrk8O/L4ml103gV1dQzfIin7tezFzxyjb50reuuExG5GVs16TrT7GTRig8
nsuDKQ1MOkwlAWmQtLU8r4sFQ8XQJUwBkql4rcBfWz0NpouwRu9bDXtcpAg4Kyjf
k/v6mh0q6QVY5SrqMAKztw9n1QtIyo/Ma/2UV3HIEnH8c4Bzj/9Ehtg0lPQnwlTt
+11uRGC3TrNNeuzxBtouuCOT5VCtwslfCTsaI9muPwyVAm2dlui+2cVC6Kdg53sL
p4YcIEEYobazTvb9NupPvbWoEs1aQjJTJ6EFUE3oRVszatRBSoeH/PGXMNuBOg8b
IYgCux3qWW3jnkUPOiQCW93lWOBPSa+ajVZRdiw+dHBuyp47yQ/xoc5j4LWOYA9t
MJ31WehpmnzTvtJTuh6DN8S9QMo69fCHtigWXQBBUymdykWLKKnFyWHt/NPH594g
87YqW2heDuHPgkwzIBMx7xzaMSxQcxVPb3zzr4u2ZI5SN9Efz+E/KADR/ScipS0I
sWSTWmuSnnfyc0fMnW1dUhFusToWEqWvhu//o36S6tPFc+7vgZtKyYegTn39L+Tv
SVCG1S2X97IENB2KQrBW3cr6r2oj9wO1EOlFVQMyTLmS61IVpDwIWzvd96sJGY8j
Gij0FPqZoQ858brOF+vbNEuos1Jyji+VZ4X28tBnUoaiaNcFIYA0k6Vy+J06MFNW
VklSlSF5LpjAXZ8tZ+Y+sPJx7xSdGL8eY2gTDwGBnZj96S2GL2NhKf65hvIoSL2K
sgtoM/R14YYtiAkLYt3ibLsPxcUdJam0Uk7NlNztUdjhQhOJIIv3wnd3NGgrgroL
WqgJewboMCF3Q9JDDzcYSj6N28r/jv/1S5dnoUPMXCbhez8B6VQHfAJyPcPXCnNV
qXcl3dqcW3XRejgLecXwW3XgvhtdbQA+39W8vvLavf4hh97bEpegUXOOrD6hfAxv
nF/YvuglUKF6HyArFy6ci4L37ZSFC7VXViviGXvoaKugB6OJObaprLIpJQjPx5y0
lsL5QVyS1Pwx/5mZKTCN6NyGI5+lZnzRe1oDq/nY4oIuMl2cFqbG90Adrb3bySC0
z/NiinD3yOO5tJKvgIaXcWj1gebbw63SYr6Bqkn0wWkogK1p0jJJGMJafn58cXVk
nr1aR6qG31YRNkqHyVxQ4wvcorzic2913cMI0Q3avhVBxgpK76qznPodiEla76N+
CjWLV1AZfd70AhWkYJap8wpQFYAQ+BynI/SMm0S0Tsg4b7r5sMyIHESj699sybQw
Lex3OKq3lZ9UgFL/yJ11Wo6DcI5Fsiy6fF3vAy0noNdIHO/Yi0VAIjYt+5jT1XI8
6Vui88wTTPvosL37nzfq++oUlPNMhWeRifwmQPKz4Sc9CrLwwVnmCgpJNzZplGOi
kCSxrc2ljQ65GBEqq0XTfl/6KK5uZS2gFZ8FXvZuni6vSa5fx0Q3m3+MTTjfrgrV
Lwk5mdv5GhxM2emXWquRDMSjT0Vabx7WBRLY9pYzrXH945wlBjscXhoJuIo6KKn8
EMAdgXXvTeFiE4oGuZ/qh1GAZqB1A87aJTYG+pIa4oLzxgpZvtLevNuHNlC5RnAR
iwzT3g/aPrH6bopFOlGwkHsfxEp1WGbPP+F5x02FbFu1K72rg6bLAWms21NcbuGp
TdmChqv91n3ykgsjqGeNanXxFVSf7rIKYxRGKoUcWvtuijstu2nr5eAB7k3fTXRO
v6pBm/x6YdW7l1WzJnVPXSkQRGzCebRGKhJmBT9r7NjwOppCvlB1f9qu31Y4wqip
dfiY0nRUhZ33bHJxnzq3Yqh6+3q2N3THeJSYVwM2uayEv2qcacO6Bi5j8/9ZHrgd
5TL0M9OhgR/mmv9f55La4FdHzwRwO7FdwjVDJ4x7BChlZlMVrUx66iFm1tpyEZO0
WW0XeU6ym0zVJ4UPJv6Iwr37CK9QenmhBEnCASR8s32idyaufBDUAkbXx5q5g+tn
OOayqWP1ZXDNxUau7He9NiDLNjCun8zsQVXI28wwEmYI7y5zmHPeI6EUsSu/ldig
W9+p4lKkKG89XIL4WUOizNlqzoWL+fSd3xSmDsyK0B0fpVAoKDFWHifVdeZ853iG
x9aQrpO63i38JxQ2Zv6/5d/uUxga2H7ZA7jkb9SJnPXTNDVcCU332JsIuKriG1FH
CXPOKQyMVr6qhhaLObmrivfo9dgFWsRLPnSJUHuFuAdPHciDoRASjz7CGVXaAJbk
11qLu8qO4OvDkp7nPg5MGrCyVStT4XVNVM74Ed/PZ+HBd2JUDhBWMhVetUhAZDEm
x4XX90jsIMQbnNcrf3rdhaqp1QYbIGgAVEM9ojlQ2LqVLZ/q9XQX/cBAcZ0hWkd5
ch7iiazk6aPOXk8N5wcgFzVjVWxYTVyupeSHcT4MnImHybwa5agCUuwQEt9wuFmv
uiUr0wo+C7QaOBRTrgQ5cBJTVhzMAUmeSwh4lL0/r5Z/yJO1ckKmUxGhZpZmqfKA
kbwkja52S8o9BZnNOHEwnkiz6sxVIjGPLtiEsBZzWX39a+TOlVlWms7VMzBIkMwT
K0edXGYoUAxraGhfdLwYt2jJfbpYRt/SoS+YKlXYpJb3cnO4HCHcDDVfv0T3/Uvw
GEv2z3v9iIdZPmd503GSiiFBx+sKsYuNVB6T3B/dvehh4tiBomIGeL7nQne2RHe/
QBrqjS29tHDR0/EF07RHRd3GcMtDVOtX2FJPT1f/4HkoSmHGznQsT+p35GxEWLii
vUWglaBiWEgLAN/LGsBGp9yIo815CbgijszSuhSGyTcMn0rXrkZhVOdl0v144O4v
8baIk34DlhfSpqR8uGti2P3ujcAlg+HuonKk0ZlF73EwRFqBul7s8zf+K2mNHE+v
PY/ygZgUVqBvTAPmlu9AUM+923Ys6/VCFUGSa2FKk/dZea8baEELid5HxxXdjECx
YGyaGpHBdmFGPMcvwrl2suOIY0yBiB/NxTm5F2zqjDWFaD+Xu4bl9JCgMjNCJm75
JHNGEk3iPDmdQAL8VBke2sD9sOm8/wyrZdU9LOiNuml/Aus+AFMEHR0FMAKJ9J/w
cPkW+g8eJoWwon0B41/CkUqT/IP4nKWo4/j0h2oBxk56+Xt4XOfygRN2vDFmw+Wp
6WrID5jNXJ8pYRy9/QU3Nns4rBFRl8AZv9oCP3ix99lrrkdZZxInwGoMduNIm8Vn
uVKAI8rmGlylLzN/OYJHlRjLFIkMG0O75EWELmlFik5cz1hZX2UfEoKkXvJGPSuV
jEIKPskLq8rih20oSrEUGUZI3/aN9YgiRiPnLuNvYXFAWSNVNEvaZ6fbIjWT+9cn
MKMVPUP3q66zSqZRkA40yHUPZeO4WMaEcso/BTtJ5eEPLNZ2PG4WzwfVvXsG3fkh
glo0xUav7FPKn2p9thB4s3GDTd0lLp43eUzmmVPpsy25wYw+xC/XO+XP4f4FnP67
XDT1NHxTCUmMJiULOTGz9xTW38BsKY8ICffhkUzO/M86MhdNrS6EHa8lR70+sL4X
XbmVijBVXTeNbaCWW9jtD54xwnNsc42Hzq91JJji2kE54A4n3IOxSrfGUuaqQmv6
hquXlzBLzDF2Q6LD7GQjMJm99sUlHoCTVNIT5D0nQGdP+FhbLrkCNh3C6Uj8ZTm9
GjbSQ525iwbpsR++j39n1daEq51SHtsbO4r2MHjKXBoy2kqjLeTD8LLlu7vebxCQ
BrYfi44EW70JaZd2VUnKqeBPBzo2SQLw8XXOVJ4yE3S0HilFj9MFMK0Nh24Ruvt4
zBQxLSOZCiy0kCP0HHCpX9kte56MB8EVpe9HyV+umdgi7BnrOqy8CGZADoOXONiL
Gt7G97fTmrMjLkv0ajNSzAnoFoKHn2soG4PddaSjJtIzXmYs7B6gazGU2WtQOv34
Vl0c33edcYNdp9CgWEbl4bmLyoILblWw5kTkUcNhA4+VHTjrMDwhQPXzEwM2wRnK
S0JG/Z+mN2Vos11PNaK3OIq0NqQKU0Vzuq9R2F1DlhEzv18/yFi0F8VH79FErw0E
vhwnK4RQWrFysszPtyfAUJ3dUvV7ZMpDhhJQMpax63xJ0NxIlEyor7Yr10hVmtPE
9TLdNsDjVfLI3t67WgUTyb9hhIwfMfV8+bnJ0KIUN51PtnDGlLA8JfffUbU8uVIR
FvCds1ANgWpSpDm6XTq9Bk372g5Ra8Bs8HJDGus5jFVHe7W9sijejdims1dyyGq1
PXhridzhetiBlhCgNIpuVVjk7QKpsQExHE+u6RV0GnNCS4Q/uhuA3WujHZkLOYAy
RBoi9uFZ6Z6MmqgsVlpfwCaApv8Ie1WUynLd4W0bYzEd0pdLTsgcxpL/M3mGGAnb
uDHurSpgY//YZni25V8S6EIdftL7z16qJW1tQowzLn1bGq7YuiutjeV64zb+kqc6
KnaL7LyZJPOS1Ej8mAg0MNwX6UCKFgrh8H2hj75vlrjgYZe6XxINBZwFVgc3IQhl
Z/gYPrERhow83h5ZZGi7WZO/+86tonPHvhHppEJCoRu16jXetMKWVmI1zieHDte4
clj210kIYd6R+J/es9YVQUy7Ks7QPvmERFHzrjbJvRzlphxSwvmYsZdnlFi+DF7F
qOzqq4U2s3geCjzEXhgBwqp88dsR8v0nYpvIprhetzYITN8v7IZQfkeEKNA1GBx+
t0fn9YnGlbBIESe7py0aeThVTTSQ+kF6CpDVkHDigb1co/iVIyID1CRlRRc7iR/W
e9y7pshbcYwQO8OAHx6YF4AVt4Yp66MOiKApPdRHnxsMaadFHrVChRQp2mymGZ+y
IXWiZv99uibbplv5sYayOlcKDC+ZZXAvDmCIyUWmxydo9h3toUNpe3XSrFEYNam8
4JVgc8X/i2Yb/qHaQL9LWRJhVmQW4Xl1mwes3FwsImSHL2NXo8gcszuleogE0FL5
qUckv+QL+pu3aSCikdDOlAruXVcIyx0vPeKAmhXVSMBgHOcPZ2hlqDSGMezkSHX6
qL6rkf9itzBUXKvVAy6xK6aAvzlN//IJ0nz581GawoFPUe0Wmw/HS1WXJ3+QkIqo
dq6bbGak8iWrfNM+wFaUTd3TRXLQBjRYuxqkhZopqjBW8sAdcN9mH91LiVowUPTF
zLpt0fvqoLC/qlxhSjz8D7DWrnFqbed5gdYxPVanPrP2CHzndIILJR14Mob1PgBh
k35P7osktDprBtX8nAt01nReiAQLF+uH4idvz+j5SqqZON++TItbjzcHkLfvE5Hw
/dnqNYoRC6VHHGXsaFsszWRa6Ja7ZjQLAo72Me9SdJxLgAgcflNFshzA1ZkcWM7c
j5pgDoQhNFc8EFla9LjN4Jt/r/5JeIzIAVF8KNi0BAW1EhUvBGsMfmCvM0kHc2B6
NblESMR5537clEzd6Lb5pxqBuud4qIvJa4D+sktbxSstaHrn8nEBVlRJfMqrQwRB
LNA74NqtzncOzZWmbwAwfy5HLjyrR12cJWtSQZcvYObfVVLeneE0wgDVBjJ6ZmHi
D1LKCMHcu6QAqpjFJeAlu/fr1GAHAhhMY+kvKpdsfKxpX94mfJBeZXClh7TU7uJl
QjVtn5xAGfCrKoGhlldwyDXk1zht/j7QrKU1EDsa3W7MWxnNGcQg1e9sTaQP8mik
hWxk/egwv+9+BsFDAZ9wC9n0lSzX9CJ0FtkLWoDNgh3Qy1uqtPB5lk022E604bvW
KUdJNLaHV1z7fq8ArVdtNIL393KVEGrXESKFeV88raV6SwXlOV9ZGmCQFXAi5Xdi
r+9IOV3e0hppFO6bAjs5OfgALR5NLHBalpwum0zlEDrH5N/qa3SoZYOqX4t5+KX0
maB0maaZfRnsn1hAEBdsrFYWoP88/tnOkhM5R4SDSvTfDtvY468TvKxf4v+CU0/X
S8SVYNZVBDuzSOZCRP9I5EhxMRUvF1sDndLolFfOaanNouyYUTFxjs2dSSe6Il3J
sRPaaY+qnhVBrlxCFzuJ/lvZTbiu6pY6mScbpJEfsl7LuMSOHWL14TpZc5NeH8Ek
HAbIsdrBhF1vjcYe05EZxBvIp6bo4kDDo6YBN8XtFAoiDCQJsGxtPfGFQ4P+1CnL
10zKBopO5zRQUnpSYs15Cr99P+U1I1q1IYuK/G3yEWWK4G0NH7g1QwWcHPb7Blo8
Pc9jvGvYpMejGGx/PW0S44D+KEyp+KcwGrnmWNfjin4kUA05t2/rRmaGryyYyg7R
LtyhfFnjU/HCP8kxrTBlz3qn/5PSa+BqCRAoCl5yQl8qODuR3ykPFhgIPtgPLLFK
j4OZ1UKoLy71umM4VNmezhnmlST+jMKcMwFIaBtW9/bkWPch2MM9jDSlfYJJ4lAP
TAg69FfsSXF23Uz9thiL3Sb18GF48jJPhO7DOZO0cBuU9MK4c9E9mBnX5M/ir/tT
XrPJU/syGJiCTYzF27HjkfvGEhTnH6nj4WGeZLMg403BEc2kYo5wXsOS/gRH3cyB
InDfdvXfevxC50buxDHgzlXLLEdPoN122B3njPWZISwdXzVWdb+DJZmMBIG7msdD
Ua6kj7C48YhMiqUoC2GedknOF6vGfJaylBGctGd4ZQpYD2uR4Izlgs1VP/Qm+shZ
O1Yv2nNP8qOEfSoJILMmCotbFodxy8CYu7i3/pZmaX54BBMZsqB+qLXNLgyaEcnc
SiOgZ35UJltBqRY/tRdit6UL8G6Cbg0PVYDElc7JYxWgiUsHliaHQDsXw3xMuTA5
Cl7Z2LKt5gZx9MAgbsB5BcVphqFaN3OeiOC7+CzU14EwibS8SMwYAiN0L8B+jbDn
yaxfaYyDBYiZ9Gm4LxeKvRjNX9Cim4dclSjoaIcLxq/uaqiZQjEeGlrMl0i473W/
RO1Lk/J5XTVC8bY5FddlaY+u5n5NmKLGIMcAVZQQui+BWWmxNi1586RTex+j2RQV
XWMXzNxf+lmRokG1Fh7iInX6wEVfuFzwi9eLpQLKzKgkHaG7tjHzkkg7MLLkH+mL
OR3fNKYmsLXdNiqqm40qIk3aRdQ6PY0G/pVzaamuxoYQmxs6FIjSML6cFsHz/1EJ
wU9c3ekPlxdUCcgeDYieaWZDD7rmcjtCB2NNwKluZX0qvGZv6Ax26Q9vQBhoIAFe
b+YIm+yHwGOhtGUYWLLTpVQOqJziu9LcxK/grzr4Lcq9rereXSwiPUC1JewfpyZ6
MyK6l6ZyXKxJaAs3rwN5NgYKj6n/7HYiRtM3ajM0fh4KtCut/lGYQ22na0qtwQ2f
WveR3a/xvZpyITvh+5lqL5eKhMwS3t4KtappcfqozqjLaPxBlj8RBKYMFGjCFu/R
VIL3Ln897/j13PA2lahNBAALoxNUMBva/t/9LbipLee2YYgeF0kf7LecayDgJMoh
WRg2PkuFwBzENCqjycuMdEY3UFDU5EUqUBdIxMXWk5yo1PVvRSuHJ+ch5VaHgp6X
WQBWE+NimTcvlheodqQRSH1TtB30eThhATmTzYW79QVNpIlnCt+Vag46gIZn8zz2
jM9l9q0Aw2XGLB5ej0qSN77G01gN1puEqPAk+2yD9TIbDLrR/cLWrN0/+CIlwZDb
aRDMeuYrGGRpcfMB6dMTmQ0S5qMEJGlqqKRHCXvK2IbeMr/GjaDYJUgOd9U7OLg3
Ml6KFYE3aVuoXhrYghmlcIF8Fa8qaT/2APYrI9hEi2t/+Qb0NVwKuLokQYsNdgxz
Pblt6PlUr93nT8NpuMwJIx4R2pV1cTnSHXrozieTC7BPPP/GZbtmwodUzZeM1Gnw
mj6Jd8Vp0WFVrQp8rOHvfqOeBb+j0v47Q/cy1c4BD81G/tRcoQDhb/ZMdVEdkkZV
qlIvf9+3kKu3fAm5bcw+t7qo8IjApHdPP2FnwECO8Nspw8fB7y8rNFO+i4ZRHERV
bwSH/MXHYXDEAs669jAxK5+a+aYnAbrQovnlC9cBvOrEPzTIycwdrdR+MvLn2Gn2
TQsPBmBjCvqFSnTLTKCWX06pU5V3EnH3+v5oXRkW8Ud+WgnnsQG53YBPOLGRMAYZ
YjKRIDvtPv9r5xiyQFG5emqQROaCrXJ8Xwei5MkFCjY206Uk2nS9/wDBYE3bPMqh
TeNTyEum70TMnKo8bIjPXCEib+QwADaWmFsDdE73ZCKjs8NoYFsc/gbzOebjkGD7
pUaM6w/R9RGMEC/gh79hOk7kK4ZJNZVdXyMUyG6Xxsj1N51+U6FqVwNNUzonJAyx
JMy/IFuD+VWPAfy7LsJukHOVFuDa1cCJxt1QEDDtVFAF9YcF8peXEGRZo90xgQNh
Gmzx5C+pKzlxTo7s/Ns/tysPQltRlirbMAuGLuPczzbykktxzEPZeSX+iSX6AcWN
vbXT8O131VVSZKM2X7t0qn132uSOAfN4hDViGUGLTH4oMykbpCWeAVC1R8RbDoTb
ID5fSTofMuymCrSAGZeqZytbGc27Genl/33Pz6HU4ieee3e6TmD1fRCYsdb/SiDe
YWMZ2H1aR17Hgp1ri2qC44p7HT6Z/6AtSzsxJYDt7ycz5HiDDCXBNtJOsnFZ0Si9
HZwvWoPkRLY6GAFFW1PErDKiEmJ88a46roz6CPwDkrz8+jKyoprzzMonF4NgG0VU
cVOohKlRyWaay2jWBeTkzrqQiwjENzBxCAoCt1dSI123z8SAAvjsmrw37cdGYxzF
ByCdH6DsIO+QMZU6Ez8TXBqGfpiad7FnPqLGQ/ciQh6D/tQ7v0f2GE+7AEa+Wu5x
bs08C8AgSI+ec6xlNtenACAWlHmKSB70tuOJHl6M+2KbvyBa7dl5njZQG2HB7HvT
mcVV2B+yfjFXbYnCM3rXOu+d1mpdvvO4G80UGZUwnonYwvcO8YQ61lcC1BpIEHGj
KE8TICYJZuGZcQAJMm/uuyLEfjBO3N9joqPdZXzzWQGWstmzKJigRPgeyO49sL3w
SJ5mD0kn2oVMj0aDatP2WR0jpBf3VFNnaIay6EN0Ax7YIA5PzbB9I7jo9SM1qJMZ
0t9tVsm1RWpOI8Kte4l3O4EWlkDP9l5DY9wMwx7+Bt7SNnbCu9ctpTUn4t1Oql29
vQixFhXrctRJqVe1qwDaK4Bkc/bWUz1w5EoQIL/gxizgmmENV1OUml1aaYUIlN+V
SpSTRxTkDH2a9Z3Q83H+d/NS9XJN/JByhBBXtPLJZoG2VBVi/trZgFLV9qOgYdA4
l0jJ2K7dovEtWCM9Tg5/cY1BYlxm1RViO0WjIWFgbtxQJczQRPcMh+qmhAuj36vs
VSf+pInySktVoug1rU9hFekZGTPM+KHYbrODi1sVnOQHXg9hpKD8eb84Vh2MPH41
umV/OX57Tn9iYR3/JzJIBVB4XupM0RXh0OCQPG3hV4qXNlQl9UmhYy7OEsvhJyZk
dvUgRbSxgwXgcf5nrBLKWk9D4ZoVYThJxtHlK4g2K9ZjRX5q7bTLA+y0iYc698Vw
+L36WCY2mk2cbRG92h3+70/SAr0bDBxiIWQqMqxbmcOrgzgLqXO11Xh9ijSGWnGV
1YN8EPvfuqZDJu/KI/rKg43aYG0/cQpP9hCvBQ4A8ufL1pbeILTaHss3oCga0ZiE
fHtA67wMFpBQTj/4DGI2Q/g0s6H62WY50uaYbIz05zx+mYHDtWzQimBj8kUeqrpZ
0kApz8J51+ShPuuj3JOev+xFfnsdVKzwFAIoYkHXAs34qgi0peh+rTz63JV6pn1u
p/8xrhJ1ijRjVi0XV8Nm+He40hgMkoJpHZjaxoEibh3h7NwVLoJErqzivzUBP4uf
nCrNxUUh98GCofOexpaiJk8fWhrMzB7mjn2OJjN4mta0ImAQ6YAuEQ7gHI0jq+6P
5/dqIcmK22r5ogVDtcaI7cDiFGBdMV1HPyhLglxHWi00B9jzgdHp1VkEb3xzSW6S
EweVBu2Xq7oHhl+HImitClplqqVBsyhEHs11pR+9URr6nqKQ8QcqS7S01D9crfTt
8hBpHfn0j07J0G2JmvXzk7+pJk+kDF2bsdlS87AzuSq9dooGtTKWGtchlJ0v74Q+
M7JMvQ0NvPdvtxNmsJOJcdHWVQ7ZCFf91kLkBC/9vPwZrm7cOAV4nDiIjAYS+MWO
gdGLK1G6iWb4+PScnJIlYBWE6U/VLzcUs/k8KtiWwvVsgEVYN3VQZ3SvW6Crxx76
AiwWJNCua76eotTTChKA/1andQObFrLzBMZ7v2zsC7Fj/yhaa5kFqnndyxBR5X8M
km/9B11mu7A/Cy6LL6Zm7qP7g7qVkEG3Mvme1+woqS1CnnQrstAZ3caBCNkbGFfS
BQkoCHtxOi1WyScNUvvmwyOi/Sy5cfwp7JvWizwLBuR29oIs9H3CErIf/7IqR8v1
QO//pH8Wi8y1WyHAaGY/5p/Fp2IjRJjZz79knq0tuosjYHScvN3SRJYnOUmOCJD1
jnDMfvCvvlaxLpnBY2owOvFJpQ/Ve6bETdqcfxLBxJbkAyeyDW6cGJqLL9PD0xcH
x3jBz4kTbfNu5vn2/ts5ac1LoKUB0xaNhlHBINFdTLgoZY8XuxeLfv/DC7UbWldL
3BeAaBDO8zEAe3anytRISqfUEklhkTgITL+BfIZtiLpz+mQK5rsbdcCXSql8sXNc
hZph8y6QoFmsj0TfOTjZ0wqQ/xqQLsOIAvLLsL5STfDm2VFgvjlAANYT2tra4TAF
DxkvNJnXRzChZ0VTU9EafpdjvMQpih4wS4M8Xoc7hCP0pcz4DZenJTq5hb7b01AP
Qgpip6bqwayCb/EU01qLURHfyI4Kg9dA9RUpOue17mDUZCVzTBchas/5Xad6WE7C
WY4f7fR4kNnwfAGGAEXnBFFl7x7qn4ZEpz18gS3OyQmpXNGiK1nfe7O3VuhB34Pn
no0SR8LkC2+LAFn90Hp4liEakSSvnqOcIiMzPmxcFupTr53AFoZpTSNhB+SdAkWm
nyiSQqT8AaNV+N0YTv1i/t1vBFkPdJftRefzRAhiH0zMggLR8Y4F2EFQ73S5uFN2
ZPWAjOe9pOBUqJz9nndr/PDLyA8E3XFfS3mpN8MB3zUoJw7T/J8hqI+ZHSe7q1aV
6ldYVW4mz7N8Naz7Ji1OuWW0MoDLAUVE0SC/dwIG50zQOvKl+Sq7G9cqEH+J6SMN
ZwFVaO6PdSAZRkk++RmcyVV+h/OBX38SVpNFYaEiKWiGHg1PV4Zr8SN1KOt9Dw+w
yzE1IbZRUkgCKzt6VCOS0My5DZxAxCJHseMZ5IaFGpgFMf+6fPx5inVCPJDs5+1D
zwomDKlRB8nWDgYcEn019tqDmWfynO1X08dwO2sahPQaTsbVJzt+64RmQQ+W5J0g
rKmaDVZ6BDz9StHmPAPdP4r7sccMvMxaYRz8M8w27wgrGYJzFT21MoiqeHYorNy+
xejBj/FmXYZ/d2P8xx6DMOiz7SqwvodOC0Fj80Jw8kCuJfQ1Br2B8P1X/kCKCTQk
IF3i63+v3TyFEB8EEmGmTGONX++kjFiwFfK8e5OmNUlbq78OqCDBZxg7infG5UQT
pn3XAJN6AFigux0xmxIlTgbpEI4/Pjhs2htiUk5ooEMLmwmIZ9fWwrge3m53RVCS
HMnD9lto56Fo+LIvw0aEii2nchZOK3TeQ2/dNLauordX3n6T96E5ZrhBDstD0st4
MH7nuFMWV3Mnq5FTLww/ymp8eAPNNun2645n7riBXaCjcgBWZZMb1r7LMqiYWe2c
Xa0tijLKDB8S2lNAknWI1nraKR72TZmR9fHOuU083/joQdDzGYtFt4AxoKJQTq0A
ji5UefZwwa7cHs66HpfhvAxsn7uMQimjU7Qmfm9CDHsvt3DdRoTAHaYkurXuX7k1
Ku/DXTWmCWYpa05RtOZVIdaNCLgpAQH48eDZyk+Yuz+xNUj2dsiz0LdcSXSWB+39
0xDlS6TyJgZTL0C7Thwptlcbz5TVBgjnpYzguYcJB+oAdxum5/q+fnu9Bd8rtxO4
SL3kFwp2RlIeYJ2ElhvfJ6H+V+7A3gWHQ9WrJ9uLtE9a6IFcbQ2H3YPxDUdZUWb0
YAF6IXr3hJmMdKPTaFgyJ4Zzvi+R8doGJbekhWUXQqGC6LIatH5P5Fe8k7KNC4Km
Eg8t/DGpEHimFM/wGhAjWuALIqZzAR8oRoDrhZwPFcs5PQsX2ritgp1MhCeWpP2K
phrUsDdLG/EsWIrmu5tD7JfCYNCG+pO8LIrdQckPtvSfSP6TtLKnrqpceoi0Maqm
+ypB+ayq06A8DlgKyzw/11bck74ljl3tKi02ombMlK3vWUEyGkS1OyTN6tNgzg/3
noX0oxno8awAUaqP/vb77qkf9Ek/tSukr8VRLWWXpa+zrk2F7mKb1xtLWeZGJGyt
3rsD1bSHKFfuOemK3fiZdzDPUV4CQDIh8FwCNd8Cb93C/kaWpKvr4cVv41bo8t/n
/xYtTO9p5OJ6+NbopCOPLWeMldz4uXxbHSKiQwj7C2LhW71ifSURs+nKslKLkZMy
ivCe5hbGg2TFdSvarSTHujA7uZU+2N3LCAFZAleoEfkllU7zVpSdHFbmBCgdKZck
kAoh71YKFUZJAB9u92x+h6KLYVCJY28KAZodmNzsPkH1eAC9HWVoi8RdGIhsiKMW
3oM8uYv8ya1rw2JI1LjElXFd/kO+sBzqscSh5prsgdnSirkZkXC7eq8x8KEfwHBb
gqcCIrR/H5yflE2cNe2PCVt4vhP9BfEOd0IKQiHMFwkZW+c3tSwGz2iZ2hO3W+FZ
qKaNqEHG0UGT+FMhaGvQNlUMAwL27qJtacNJaRKkcJEN/ANVtpyM8r2LIApFbBDr
V03vC0i2Vg9vJ8Ze8SN3ZpI0ymrH4anofrO/4FTxm1360ZVVXCkw9MgIoD4cy0r4
/uawNqaQJyIBAjiDVearenBnxQq4ys7KbNH/6GwYLPuLA0xRASfTBWA+Cz1PP/6L
5IzbCs8duZrIz5qM0fscQL3e9wOJfl9o8W98/vIYbeaiT9rbCo0xZtsdIQ9SpRT1
t0nnYH1oYIdU67u8lFYKUNLXlPfSKu8+3q216XStsZMpAcbzukKKGYECGq0I3jRa
qP1FzAvzsJlLSy9B7IEa5Avhgwb439omcg9GiXXgqDne62vz3XO350zha9cwKtfm
hxOogU/5ibo1RhK28DNqh9GH8takRKwAne5RFjc/Sm0AufC7YhJtV6Gm/X7PgjTj
UMgLPknOs/oWc8tCito4RWfBHxGel/ogC+sPFn28RSEw8c2VmdjTRrM1TBpQItRF
j3/LP8aNPQCxNzZiN9aWO0iZfNwHzdern8sPbfgygvTIdpYvIXvXJItodP9igMve
I4a6OMyIXYVDC1trNEtw6du25WkZCzIwpz8kVjnFhKoLAk33aJ28uZStR+5e3zJk
3445DZCeldUBWXNHOtgGGRm/bYn3XaF1n2aHeayelauUL6/qNQ2zeIYrxwU2gBPn
sUxiBbLaDqEOgXZng39sexMKJsizODkqvKUcoaGshZl8mtl18m4FAfbHu/a1hGxV
SiYPuvlnaO5XhAFpdH/gzggORozVZ4kNF98eWAy78GTjBNGTM8wvZridDTAQuF3J
lnRBVFK3BBD1qPm0NOwY04FPcrDg0KyUyKzPVP/tW5oouJK0T3fiV6x7CycJSr13
shAM5dFjquB+ab/eakZS9GNASaaHbn6rSYtLRL9pP/x0qBmU8fMrdBi85xXRiKb6
THWRr6h0L9WfwJvT54YiLEqb3odmBbTmE4yU7Hg9zfH9KwE8D9hCU+bmk374LadR
zNE7vlxpxNnZYzNVE3XieSH+rW2Wx2j1g7k8oSFsvBW4C6HxCZxyMiuihHuhZjd/
2A7x+qLld6XFZ6jMF2Pm5HKJUx8PYXtO+sHcVUV6wwCt0FniT+4HmQ+4sY/OyYR0
bLi0yTg+d+6t2xYF5kzsDDTu/7aLpPX3Qq6Lm47HslnlP+jfv2R6kTF4IcqCvZLb
Qzu1dvYK2n30nDoxVSyOHfPxnF0bJwCPeQxtkFU8AQDIvGO5e5KWfOf4rCDixhoh
xV0tTa0NX9XzfmMb6DVEWRdVaI2vAueXy1OgEcb0dw7Efj+Wg9p8MH825Vc8u65I
88capbB6Lj59YY/oigPvsLFO9DqmsYHN/eBR43jZnbgOm9fRTOoUwEtkRC9b0pDZ
dyBhBKuToSKjHS0AgeawkXkitFF95d/HJH9Ixxytzw8Unr24/7BbTcP+f1OxYPpa
T9b9uOVnZYz0M1I5p64+9ncqZOa+QsnVM9fGIdVyGDgGqAVk03pf700FYwsui6i7
EiVa92IVf0q6WSHeN1p6p/gOJ3y/VRoJnostjeVZKQpbfs48p/Kk+faj6EBD/vW2
vkgSr85PRyNAXTAa52O3wx56CiXriczOGJcu/FXUKLwezMgkNx4NUqjz1CdWnx6Q
KwFG+X7opEG+mpi6yAll9ZYMbvyzhsHNIXcvTj3DVilmI5o7for6QZio3ro3i42T
71oVDodHvjTUltjA8HzdN5NV4yUZy6anxkzgS/xNe6uT4CPRwvGpn0hL1U5/p7cF
3ZU3W+liTM74f9Knu0vkTqQtujvr+ZgQ7mcWB/tzLvIW02zpm/qoSP9MnXh85Peh
WJV/HKMD8/rnfsAwOGI6P+ASduldaE6LNPW70MMzMF+ZLvWThKgeBfs7QKYZ+uR+
DJm5dBPZ6AaoJs9knaJBCqXH/ihnjSMr3Egv8a3NCsAD/svrPY+mzKJ6kUtssRKZ
1e0ZjPIPwpUv3uMCsqBz+VCPc//g5qMN2d3d8KJ1GiRvcsA+RXfRYs4htWGW4o1j
UL05SSYQyTt7+n682rr0FDi9jtTtu+FpwEiAZNeOY2tvhy1dEwWxeOssa52sizzE
i9MH4ZmSSPCwujNoI/mV6nHxnQwtuy6HKq6bRqYZ9AHbzD3o0GDwaxaZMCqRYY9m
MsuZYDJtiDl/W5AjdRxofwIqWHFzCmIKjNrMDTfVr/bOjJ0KoKYQva3CwSfGS1wC
Z3siHfPBVCUMtq1mD1jXZvqsp411DCF+vskgMAn8tlYCbK0a61ofqxNo276Ew3af
8/9WQFW9SiDullPKPrZgWC2TRft5hK0vc8HEhvvGZo9VijvphVzR4lxrBs+Z6t5z
ImUQHUoaayarhPKQRlmA7sxhfb0uRu3QtGaUo4uDpLaBp9JB+3cMqwkif4Son6GX
CylUaciV9OAuxeSWCiZW2muHrJtF/5JfJbQZZKoH2q6SmH4xQPWSdTV7k1QPXxK3
iXNTyxd/idvVH4cgNnpbFPUc603U7Ortt8ufKRE1JP1Hlvjt2LnAYnuuBnow7Erb
4ImtliLQo19Nb4mRwhcqOSRHzau+8nETsosSbziOYVa30mWB7nPCmAH/97wZmVXF
/Fxtl7QsBHZKEN+UDAFbIgJ+poqqWR7wmyVz/E+a0nJRmRbFvCEc7WIQ3mQhtil2
xZTtvOaz9g7RXrawoXlICT4FoAcFiho/wiV9Foa/ptmnSe92l6SxJJCshsYuASVr
i8uwHKTmoYc4JPnekPBsZjvLB7DYunhbAn7mHB1WWC8rMVlvFhcnRVTt8otedUdA
OLV8fdN2qOGIPagwAeZD5mB7gW1zJMNFpLIHRVfw52e4Rp0/3U6RQMakUTH2ewYF
kpe6atBXL3oDoqoGyASos8CPf1N3vpt27Gxuzl2cfPrWL3mU2vuovU60qSKTo+wb
a/J/4wmuMM9aLzX6hvd7oT3kdwfjnRtWGl+YMsUvqJJR2xzLnDex5g7lg3aeqJ4d
WyZOCeahJVe0PxgDBgwqS+ZiXHPKjX44yzRcb1qaOwLsGZCkhsKHHG6nuDF7Ta+y
YWZEHc/jqZdhyemDRVD1alDcGHy8fUELnl+4xYL6iQVvDCTWs5g1xlH8V0PtzP4u
eMChHni/INGcWcZeKpV5JVOWzcHagZws2Z5Fctz8Xe2ysG6hYtrbFfnKgl38+T/X
xUBSi6FW2LOLkcoj/ZW23hvQGBgcI5bp6gIIsPjm0+/E1+xUtJyU9NjvAGetOJ0l
+wvUqIBrm9320KFHIiOjFsDe5SjNBwcxqkqcd37D6zGaWqrb8GeTlTlLg/M6DTib
HJykgQXTgANWQ6dXporcYWbKexby9+Raei1K29E1OopKrl6xuS7uapBx6TbiNmwk
btfrmL1JQRwYbnzZ02N5+dCBzuSRtwHWYfae0CmhFuiYTHOpqnUmQP2GBLuQUDOz
cApG/JcXRWSsGJBR0nsUOM3fBCqccanlK0B4P0KnC0BfCZc6W6BuAQAAwViqlqKK
McDFRIyW5tqk8rgN4v8aF/nDpqsh9uve8GxdVN2rFwUeoYjc2gzxrxReIHCB0Xmg
QSpm8fqPLM18eLQPXv7g9x9jXH7bCGVcr/j/gF+UP+dyABxuvMsxh6EBxQBOQKGw
+fmOQI5zZmp0ab4hOeJjVgwN3yl2dEpKM0rEjDUv8I97ofPC3cubb2xJQs90rfVc
6s+UFAgCMsi/zG+yhqH2p1X2QvpLLXPrQX0sz8Arx0E8akSbp9qS0w1RPsEIMrHO
pxwM6kXyR++E1vlrCh5cs9lWBj/IqVKckQzIuRDhA+x+7NEIfydzcBEZKDSwojpj
smLCW/UMoaZAy0zBoFoQ0QhkKgLT53sPCnjM64qGZtZjF6ju09ktBhWWNSJ7iuFc
/b/OwJz1J/Qv2DuXNIebUgPoTqyGSErzi+pvkiHgs+OwhvzQYMI1A5SaRIiZt9Az
p/91fP5USEWsnkbGhNiTktWnfTNa6OTW7xByd6335/DBdsUch+nwjrx8Wwbh8rPU
pfJSgvasaiWgE9cYA1L2Iey1CgiVyDio2m/KF7B0OxktKk526cTAaMFPQ1HW+Whd
TPD602MA0ZXZOe/2wuSaqKPp2nSv2qYJ7mv5wMGzdD0MYi1Q7+s3EmtCk42pSWFj
q7pfXQlMnYZC9hyFu7eBpBD7WQnVVr7+xMhGckRTPNXMj3Gc/Y+sI28oorhTMjeN
hT73c8mr1sY5e8J3TbEp8/PsElKPgMU3LzdnZIKti21z/TP3t/S+t1LMxlVcJU8D
STFwv3q4rjqxHLB+HHkKgZBKxZ499FzV9Oc7jF0IFx6FeVAk6KS5Dq/lRQR1RZuM
5lwxamBOoXJOHekqgIqhtE0mrHQlgmOPhvkQQN4gk7jbghoOFpLUuf7NAlGEooO8
Eshg2mDs8tHX9eDNJaU3xgbjZxI7BNmHTRuPmj7yBlFPV8Vr6MSdFYzjVDOpnki8
JsbPAB3dvqBitllpQdbHEpfyHe3dkL7ipcUK0B/TC/46v9FUriUjpve1hc4hsSEE
F9KKtnEB64SP15K82Swx9ihQ/Y2RdXyiq2j+ors8lhSwlSHXrOZq4jWYo+0k2zXV
w5jfJeLy4XGGQzDOPSVkAMVXJRkBouleovbCp2mX+xALnMkwJhzDZDLYmhlAF2A/
jrf+sGOdwtCPPhAxW4xjOsB+0XyWVdOHfL4a1GHfcB7Y6wn7LhHrZ7PNHkM154aV
vK322LJ4zLjs5gOWH2bqOOAEKqUK0ABL9FGKuMhga/mny8l2a4y7Xq8di3CE7Ouf
tsUfMqhPq08r5v0z4l8JRS52mZsoawGr5HlrMBmZTleEI8zRrRA48zgO46cVqQ+W
rd1FD6H71jyQJTQSUMAjabkPnNiXrpxziO6EFM9VK4sbLhViV329MQQUaTJSbPgP
IRSlELkrkUpfdASTEGQVVFwv/1fFwjRo3kXvS7q6v+JulhM8X/JISMcdZgNMAedg
cxQlUbZILB/rYQmNCsAbGH4tbkRMvN1sl9qNYLlnY6DCv5No5LptOiIeF1I2jFm1
BbicBGfmnBGUP8/Rf9pEgNLtEsH/ENbHbXTiStG3mT+5JPDhqG0DlIZBY0WCQHQS
ZItIegV8tQOQc0ntsb+7Y6EKppSRrwE7P26RqKtrANqaTTPxfheusxYOcC3Dh8v3
L8v/I+rlCN6adSbGt8UAysbfgh2BqM24ZmRLowo+tZASKLHiKL0zTPDV5U+Q4WD4
6EsAGcah5qWlqAijtezdtTXbCQFDfRmaZV5hYETEq8b6vAGO4P3JvxTB54e+SbIH
66NqCL0zUkJpRCHwGMiRYmnc8c+5RLgnwGzQzpMB1HddVBOzPB9oAdx0H5qtDnBN
YZdIngDH7kj+rPGyIEcOM1v2Ibom5qyfZjBzdycZPT28dC8EyKDY8+qYY2NqYhBt
RsMIK4CY43JIFrw0Ky/Zl6oFqEXH87U4Btpn6PTpkAd/dP+lDCUclWELmc0RIUAH
/fJBxx7aNlQW2Ayo8fyMWVk62m1z2fZ3HJiQ1NWHscFmFEDJSPb8IrMCo4AL/QZJ
vrs0Xbx032eZKa83tHiatwI7DqxxDb5uKjQRfD76MziLj6cxn/5ASeeJWyA5IHda
VFbMJrSKV613PpTFiLuh+u1qFS24doINJ0LxgvNAeh8zEZqAn8QqNfGaY0Po96L7
kWYs97xDDutvip5Y+v3JjDZyuP8cIVNHMS/a/eZYAW3PlYqgkx7up73R86Jm3SZ3
8YC3SCwXlaynYei6UxAVHCbw/8XF2SWH89NMemn4lGRb0XtPyBIQeFjOMdAVAnet
29XfrjPzPoCw+PZNO4yFdxh18wXcV/zklL9SyZNrfy+mwYDKbC3YEefpOOZ0Dcgy
O1b+NLDqONyUqyI2DTaXZPBsNRgJ01MRFoc/BlGoBTIKSVwWCrO36vdNVE2mA4+t
BtL6mvbOkZOxhmuBA0G7bDGiy677VpI3grcWTOsx7RLS4Mid9Bytn84d4JdTy7M2
JRzI8KLzxIG3Y3Jub1jKW1KLUiGpjEa9ANrzfRgGAAUNRFwzUp91xa4lVPjm65JY
19nPpejh3qaXBNeXkDv4EuU9wan7I+En0pW1PXuEf6bdZNRibQte4AhczQdRt4Zc
jurqFZ3+l7Ch3k2qE3oifT9RDNALdP2CDiN8bwljur73mJCygOA/yGyTe1fr5tgm
Nw6z936uD+P+g4tFlDoFe0wQB0TLm2JYpLr64sWubvMnXujAbOE9VkGg8MGqIndL
K5GBmiCJOFjc3gLcaFZo+NXy7ClxV4FESpdU5bxVHpLGCfrO35qL0x9zoTy9ANAI
ns4r2ZNifLP0saic9CEJg8jrsB/dEV8F2ocCitBag//2S/6VXWNHhc3ztdrGCfDD
xPt+8SW9K/A28Lcb9lHzM+GqC/+dDP2Y+PBF/TcVVuyw8E3feI3YZppqTnAevsom
Q4DoxyStxV5K4Y5dg2jSXFWkTW77WLSZ2yg7owqbo4iFRaLv5g6mli1xeyTmr1Ih
19W2C3bW3b8pfBvwTETWCJEQRi0RzLB+eCL4zLSrokKOAqCfY9dIZ6xYmpkIzagR
nbbZVedVbZmIuireFR5JEzeQrP66GDuEGBHvtb5w6qaJ+6qRB26qvg1kjowNqltV
g+gPdIKy39suuwBz4j28WdndI7O1uxtTnDbhePSShKEa0W1hUi7hsMg8WB3Xkakb
0H6qWa+YikKzQE8d4H11LyjPkJYIAYF+DzLWUJUxcsGz7SVxiAYOHVq/bX4Yx+Sh
FXou8T3TjV36gGCnJZUqO1W71LylR0odf/iD/ZbfSBl/Hbem+sJO3soG0ap/QyzS
weXA78DVP4NoO3eEjpzsmyGWn6ej4kxSbRpLQdKCHEJC1HXNMkEZ/Gz3rXZ1dexL
vMjluR03ljfqHaih2UDsfO87eM0JWSwSlaJ/1553AuBac9zfFRBrU01WFUkdOH2O
ekuR32R1XPXi2xE1TDgXqQW0+QGTzFXTXGqs45VVW8LcTEVrKs/Ly9VcF87Sx2Jh
FcEoR7KOat5w47W7POr7R5g4GNNITVgp2oyeM6mrBnfoQYxj+l/8OSCHHdJlX78l
8uv6Ag/xaPASWMJnb2FUUejtNmlVeu6zwzjLGW3R4VMnxKw3LeDn7ywJ/42pvHIz
7g9cn4AaTMI5Y+6On2Hru2p/GylHou2Qdkmd1BYX3L2wRwBuBXgQpj3T7I+nioit
XFmA6fVdypP5p8v/MgEex0P71py49a6iVUCefpWefNF5K5wVel2f6K9Ket4QB/AN
af/lbzT1cu/graFAIvOo1+SHGX8NqWuB/EdrwufeaQQb5N/YpKid4PgqdMxkKsrS
Bw5sjXU3q1fXp2MlTrMzj1Sg2lwiXyYAoCuRFnLAd1tnIFg+1LFQ2Pc5dfCUkoLV
I36iPjxEX/At9AhU5pUOgI2kqh/TjssNYbMcFzyDWipAbJJxsui5NyMDIUiUTp8L
hxlSH+5nsICwXyPpziB1S/QkT6nKpo9N81XmphhI725RN/qpZad+gzBEsDsG4hkX
IyDJfVmyQ5+nvyviDxSuhGhpSt6ig8EGXOI+3v/wYI8nsD4N7J5CTzDmQY5fp7GO
IiQj3LePQTts3DEPyLFp8AzQdv8xyvR9ipoaCSR+eKZJLAnE3olkFrWxGzGpEZOA
u6xUiY0mzxKEkMbri+lsPmNCfpzqScJoaDf0KiGtj25zYsl28Eo70bffaYYVrvpw
EuZV79vQp7pScYFC36zZ11+5dqwcyt031mW5h3GkI/wwgvLQJEhtlkpGdGAqSASE
EewzkeeAgd1RM+Xrg2Dpa8Tjr+zCVYwiUsTKsKLTJ/NYOiAsnDB5jHfKQyqEct5n
Llxu9hPJrTRdrCTfpU/KA98y/fqA+lUrRDtwFQl7BNPXxQs5yXjIFpFAZeRULWzQ
VMjC4iQIi1bEA/GcYenTI1y+mYmOVrlj/3gKlyacu8jRVy4UGCDxze17KSQdPtXI
JTcHC1PB+GADQk2fHZwKYjENgyBeBlU1yLwI2fpvfKVwt0UFPZxDpAoIjQZu23fP
IU5wf84ttr7uv7xwQb3WQrSJ9mCFVlZqNbSAQFk/Xvtb8rye9qac7mA0TAgdfM56
JKgrZe9cgj8fqIIdXFdaYl0/sUuoXzB0m/GiKp59kjz8jeJHmTVEn+HscSfkNUDI
6Ljg70ebaHIV8x2cDJkX+H1HDWJOwqFtDNQN81ED8gey7kxC6V5spr4CqxYp3lEm
VlHanVeDXfjrIDa3D6BcvWrg3N9cn6btbUzmBlGte2zUlOoljTcVB10omrSjRikh
QG+TtOHxAzdak2smT65+5MyWsz9SmIildbU75fpBAkRP3h8xC2+1zUxvfLJYWYUU
6BUTB0umyS27iNdyNgjSOeDiFagDLtg1eTRGqTjmpLmWzIBnN6qRyyHXk9mfetEF
QHKq91UAAyiEpGpqs+rvZ/BL9v7CiY6GfJ96dwhtS9m0r7dasP/QdeETSTBrBcP/
WTREi4x+K0/P7XFkiBdd/koKqGhSuy2NTJ4papk+mwzh0Kn+pXc2mY12v7I37AfW
ySEqrjv8c9k2jYn/zXVXnNIP5E3aVxKwOEtD459nbFQ8g126bikyvpciPhsaENP3
R29neB9QdxWprm4nlBgv4n0AvEXV5qz/FtIhWjGxyjDZINxkFrnftK6hyVcp+kqr
d3RfYauXrJmfZCjqx2mio5icE+rEX31rx5gAHBKCw4Cl2dhk88LXVIAIkr6bk3pM
NNbfrWtSH2L9UsmTP83cU64roGxtdYjZyq2r6w2K2h6lt176j9OdPrcikYbA9ijJ
XSezFTx8djQsRwg4eb7GeFxzHDgQfjP8g9MUmdj/fvLfMuw2PZsw26wYzJvTVaZi
k+b22NuuYXU++hIMGVzFpjobxsRVEQOBvCF7/1MD4Wuu1eOiIdwEb3r0xUSeoGCU
KmnIVGGPyffQBNg/IOtHLAiTc/bV2P3w/bdYKifhoST3S3TAPAPLWUJnTZ/CMwnH
XC4/Gb2ESLplbgXwiY0QI0BgiinL+I5AokNCpi7/jwISs3Lpq4af5u2rND2miElD
OawQOlsqIElvN/2JNvlueQL3D9Y3ZdEKg19vMJZhodN2/soeAbY4PHTRocrmBazA
XPYFAC8ipKnQvpOdFQhyk9HffioKhcXBcpy/SCJ+McsEbb6ePintA94PGUT13LBx
B6VJZ3RbhzM8D/c8qGx87K745jO6jYMQQTqcIKwhk/9r17baZRqkQhFPif2RMDJo
PYLD5owORlWT+/Pq/8HNJv/R9B3zQjw6ZNWY0kdQz86PY/qLTt9NOkaNwiRjDo/j
pU6/++tF1FXTco05CoZwGY/06ouKKq4e6n9uhsSpFISWmwGjeIx6oNoAOa0LTen7
QQ+ezPEpwOtJmSFT6PyF7CASx2fepuNybmo89u1C6cRibjDDyeeuEoDolcMswy1s
2+Hq9437iUvsp3ogib4+nLnEEuMF10cjJsu57ceQHCyMzRrFo6MiV45Chm1Tq3EO
z1Gb/z2tZWUeg9pS8qW8xmyX0yjKOR3fdmhafNFzQxUyWym2plxnezxdMUzAIQjx
vmW07yDIWCQsastOYnMhIo3MbHuZVM1Dhqqmn8zyjk3BbItJbU/qgTJcwbHPIbhO
sWwR8cUwGBfb+I5Cuj99FmlQDMOO0hHhY3bSPeECXYI+i/IidoGrbEWMQC0Cxxqi
P9cGMzF4WmKVg0/tsN99+4vaKmno1R/WVUfrhi3PZG23qRRlgr570cPoW46DzR68
apsgE72fpDdur8z6ZvkQrMmfFqPqmajCUPqXRYOkjh8ULkHC0qsK1V1rLmvJyd1r
gC71EYsbplQYEERVk92uVcrVSlAy9qrBjfisNeJvpXQLihdJfytBgiTuTREe2p82
QhtNTb011FJyWsqblM2HpAr9kUGtp4DbHTG5Df0bGALdT4yIem0F++6RyW7HudVZ
k3466LfsGqJKK1xjAbFrpSGGvC4c+X2OFowloIwBjLeW8UnRyMlvXYQbh+WBbX7A
btyBsNGdESQ5inW5rvfaA4LYnjfN8hng/6Cy1MTYZxyl5GbLA+3u7qrFoLFVkixo
JVPReIvqjTuEZpHBldTk5PMpXI/q4fK6wTl9lbCJH7LHewHR/jxF7Q4sNz9oLnYF
SbYHE3scUbgqKn0CuJm5sauL46VKY2pdFJ3MZgKdBksOPjCJZNd4IB9izNBUhAXf
mW+Hm1Ur9O4qxgu3pvD9ZwrvgxHtIk3iLufBT/drXg0nKOXUHn11WjY3xunxblFX
jFkbgmMU24dKfRWqV2Axj/TTrAYuv5N79dw5ZZzPNfUGZklvz6wHxY0A/erA1fo+
TQlZi128rSSoaXm8QsUNUpbtNK7KmXp5tiMBd5janaMDFBIbG3u0LDnaEYB9ms1o
3ur2WQvN01mwGgAbqiIotKYzE72xkvC6cUj4/tBU76cC0jXygruy2zfrxKVAv53Z
s6xnZ/G6WFvEfZWaPzGFP/2UEjFEPTQtnj7K2NrEtWQ2NFJyypC4RPJ/TKH0xMt2
mFeaZEMbdPw9nHg8EO7r95JmbwlR4jDmWXWWWgbGC4dEIAwN8LMGknyjjGvGKKVD
Qms4sNSvAduAJmvW7Q4LcncKcCYWjjC721YAYQ9iJtf8Up1GMNsdJ8xYN8pMAyBu
rbd0twKbX2wqFucNfGcUmpU1R2yDDY/AkLh6wKEBZkmJ2jjtUARqNsApUyN7Ym9U
7M0Zi3kf/dlOkEz08RTJA43knNiACiANp2w1toRnhn2EXEnyjsHoQDPC+drLfHjo
hBVggNZ3ZWxqmHoxfulLtVkurXtiPmzE4MDcHoM5P4F6zgJ3wTyj/Rlh9L0Od8xN
oS+FtQ5jexCB4YdI6FJKcri5CRjSAhBGS/UcV6nZ2NO0cu/61sUZae7qdFnoYejY
Xr0ro/3P6WlCmxchi9X7JpKOjigN8YPlmjGGMVEg/+T6w6ezFTQzKnCumPtAGbkv
ilo3g/3lbDAtC6fKCr09pJc7fNlAA5iiXSQMy3h0a2NZSP80FqQ601fl3+qUmLmR
IQIM+scdxdrKy0BV4Kg0yt/Vqco7FooBhDoANGhtfcSma1Bsv4ZGMVVAEaSBTRuF
+Bl8lMhjvmyW52zk2iNiMmEBHFntnDtHl/H2ygJUEg6LuDe5MDr0xy67RgMKDQsG
oyCOwkoJaEfnXMaZtdJTGaPLy/hgHWgodejqBmjuNKUdCShtqAkA4DKNYAj8NV76
eTAUL/puK8n9Lrs93Wq8eMU7jWJQCvUWtkRZVypIqk9+Lsevi0tdO+M1GlmwUgCx
JbAYrP7fig5klUeIXtAaWw90Df/G+2pgM9423k7IRt+sJmsQ//0Sr/hvfbbhnaFy
UlE3oo20a8wtjfO9gFcIdf0EzAOWZ1ic7tMVrzokYXyLhuOLdS0xC11sAP6Z7bEX
ishpKhvCGjFxeXefH5muIIHdXiGvirMKgNoy5d0BJTdHTMpWkyH//9ecrq5Yw5hL
Ri0jQ0+j2zKfTyK+J68QWZlLkgdjETXaszu3HZttdgrBVlMaaxyo+Tr2f/6c8ggi
A9QPx5VSu6VqUNgk5gJvIi9T09HuxoN6AE1ZiQifSw6nNTIzOvLHT8DQTVl3oT6Q
q6FVr3eTGEzSsVoy6pcKpC89QFHN2DITTG7FmhEysg1PzLApx+PVQeTYFsEyuxqH
2rq8aetboDTyhftr335NGJSLUc2NjlMaQX+s6l+j2JnzABrZbFOwSWlT1HEo3jBl
cb6SSxFgsA5kjZzovXIOdZ7TbU/qrtY0BKYgZz79R/zFt/a6/3wtYpC9zx3I5Csu
FUapLCVciMe8zGfj2EpFtYmV2cceCX6VhrkcnLbaOEih1Fv4Bq1TiAVwEy1ywspA
LAVcttFbUcx+RzpFve6GrzZTpsR0/JgJPHxyOw4xNX5j+hE/CNJTkDyMEMkOTmBg
O7XMgENEs6otURZCY64uWMMY9UTBEGqNHOFhTknQiJ9RFPOwE25eZj+17oOyyR8w
/0coZ8p5vqV10N2P86RtOtk4A2XxbTbubigGZhQtxZ+CFPnhOxkOg5NVvS4AxczI
4v9snpCMEcXcUjXCiFFBJXz52jAa04JfsHraZ+HhT0NUwacdOY9nHW1cG+jnbEHf
3tUIPF2Lfsl/YTtx9vIs7wwTQ1ZYyWs6Rxbsw+hh60ZL9RkNAtt9GGnCKOKRSMoD
q/Bm+GmIYr15kDg1/ZMLd59UJBy4fvvYaXUSuD8z7sBanPN25gNyIt0HPYvhJZ3m
F+K3VvNIZ1Wit2LviS0EhXF95Ix3L4F2iNKO3jr3GwpVDICvAWKn1yV80vlrTIo3
voD+ps2dwbLF3cNkoHGAzDZ14RUC+mecteme3YFUXHM7KFLH3g7NjZyTI1NQe3Uk
DkoZF2Jb93wVnQFuZHrxyWDAJbonSTwVM/ZqJ3ZCf9hffNGV294iL315d7n1iiLG
rxM5bSznNMJEtw/sTAMVWI8lvZqhJVuhI5LrgHohU+p1btlFyjZLtqRMErGdMGka
5aH8zGmnxX1ve74l6+asTYKk3m4W/TmAtrVq4Xybk1bnxEVLEFGSmZ3gL4Fk6mcr
tB+WDiSknt1SZ+lF+Z1MRNZ0PlY4hhoyYeSJrqxxVi9tmFHyNsKGVjDT8FHj4LXe
OeDK8cSWbxRaubnTlLyPnam1Kq+di3g2rzxqVe0Z/XlTX7JZ3f+GOa9rbP5qtSmA
jH02Qr77nQq/Y4JWnFLnZ/M2UTS+0DCo2Mf/eHmJLgo+YA5sIxflTLY7wubwgKtD
+FC9psoFzKJ4llgGa1h7ZFEgTgYbFbZ78mN8t7jLl3SC3YiEFheAePtHwotZ/lN3
OJa8hVGKYSAjGWyzmQDf6RA4HI4VHvl0P6ROQn02qypP1GmAmyh+7iI+ofWYbP5N
1i9/OLFcHGSKcaw/p/PlZfPH2Lxo2LF9JnoJsctI/A6jfiaFI+bZ8/0zTdn0tFdt
SZJGNz5POwMC7Ep63UlIOUxNXACvBQz81K/0pxDvIOyceSyUAf8oJ6j4C5J02lPX
6oIszlHh5Cam0jwLSeTfGx75ofP6Lx6vhSr718a97gXj8ElNhs3IUIJvPMK+2qPf
yLhj30zKiscr+LTDeVHuTvZJCePDKH3IaXRjL4dUlZRXytC93PaxRBvSTbPZlPMU
/YvuPrHZApzuKUVxlKxJ+C9gtTBaITRFLhX/gXfSphzAA2f8PfrnbkjPw5KMpWF/
QTsnA+JmAnyBN7NfymFojraROBdhNkOXeUvsD1EgbHy6IfTGIeT+n8d/vL+mnQ6n
O8d837aEVxlI02+lqV9uRzuSWJFkewyMucOCGO9A0SoZB+WQcIZyPbr4jvNYdOJ8
+T/4DB19pUXvqpH68FIqARaWI3SsgM2kNKizADDCw3gpg2bpHmS85bI9m/XUiOok
MI93EE9RaaUVQtDGEfPN+LjzQ88lJ5M4qQbACR0MwDzm7RAUc7SrLtq9XGtgGOZB
gd5hYXwa2xTkB5fFrRFR/oWrByCfN8yq0LO2Qk20z6Ga1SKdY1rwA2M6HFPeFHwl
j7j31JnvEsYxTP6dEilC7xlAGr13CfpHVOR4rVp/dfdlAV8g5lJFfBJZ7e8O0Do0
eeXIHWKyu8itsabM8IuFb48YvzSylFcf3aCAvQzfqFJi2s+26CL/yR5cKze9qCHG
jF62FJ1+VUtBIKTM/oR29Al8LPCqeL6x5Oe3ajy/u3wtjL0KetMn2gDgrDMYrUJG
vZoHBNGJccXmgtttwu3ejp7Je7eZBlZQdgnQC9/ug/JWWjlOFqL1G14gNCELsrF+
CqdWRM41T9Yh6Kll5yyR0Q8ru/4vajrCiSmwiBo7McxppTZkKVW4CzOtHJIo7/sD
OixHXXsvm6ar9+gOO4bopiEE1ybhqZjCwfXz9kFbixErBkeo3nAyoUZ+5H+OS2F2
ziha8enqC6ho/5fas5GNd8FVp1KKDKPReSA0lP/QRuehNUzxIF/7Ceh9I050AN/4
BS1Ruex5r3TihV4XQ0Zrq2bhDdnYNh0x9PhyF0TmUdXI4UcOqd/Jbeh/XpmZvw2c
RsUJ2nSWOv70iEyMjdi5IWH0RinonAKbLXuI49YlfZYdEO0ZBtArqdwWVOD+x+ys
UF5CnAP4wU6ODW9LKc7sfQgm38lXzgclQNWWQc8QDcQCzpM2peCPeZy83XV0dxmk
f7N7Hb/e+wo23Nvf2bm9+KtowQ7GAgNTRl5UaJijT7gOWZCSiJG2poi7Nj0uR7bL
y6R7EBWVEKG5C4gpHAEY8DOG2x1SipFl6tch00xFWfepkCdaN5R3He4LKV1MWio6
4UMYzCGR4y1zkl/jMIke2O20QQYvQiI4fhFQi8+gArGXuJqpZZvoOlvFzKGtWASF
uwsjotNAm5boAdVXFZ9jKXDBfy9cQcVaj6idlKGY+kz9vIpOUiReddEK0VGV5dlh
ovFN5cc2LfTfQClfn/jLti9IkiGzvJEJ2P021sjVaRLod7tVGW0fUcXhh6sR0F9R
WbttInlbCESUHOS993Sb2vlhfSdVvhxDOzpGLSAs7JnCfUFIRjM0wLhBTeCxoxds
l7+SghXrFdTz8e4nJsabuEGtLvT34pnZoOGJ2U7Eidrj5DYXw4MfULJTyrmccQcJ
3t1y4PRdVbpezWrme+LCy9bZomFw0UhReqEucjFdjtwyQAnX20Xc6T5RNvtpGqbX
0tvAUKWmdnz1Tcnm6kghy4tDp+b4wI6lBoX10HhzQfdr2dzKTVzr9svI2+7zdfGo
VklbuwwI3BCBJ+XJqmH+JifosTv29hvNtod25u+HTuQbTN2+qYjzDZE0lLhflHaa
SbkKTKK8AyCFral73QpELW5Dzg9EUbZStoEMXF1cYyMemPZTuUWBwnL6vU3fxqOJ
UavXdwyFHqvPwP9C5qsNV8JOiHvi0bd7vEh3eCaXhJlVxBrIIAXN/4o1sZ+crns1
fuIvHezhhXN4iLPAoddPM4PDuUgqhMACy0m164OYyNSakLdLo7dg8ViLJCO0++NR
CuUsUc6RpahZhvAgl2k2KB/F0nxkSpbKMPFzRZPn+RNiqNoNrez+ffb9g0oAUcqe
ujmGAR3QTbHA4RREcLimmos1jImiZToCbSz+e/HjLc4VQaQbOHMPmYuQeDQPebbQ
dWjL23wzDjIqPBH09Fn2R3zAUygu/nkgOPPm2omHC7aQqbLbp16/Ws/oWxoYGz8i
tJ0PHS8i3u2Cg/Zsfhl/jM/dg8Ejzm5u1QyJ7y3xyHcQ2b9/LgYx6JC/fPn1Od+f
lfiNHmBeLY8G6WHRpQzVlAAVj2f1Qzo6PrD6Ywjsive7ut5FjhPkEKS9/RvN5RHS
c1WSC+7Du8ifU6lQ/YQz60bjygB3wLfibO+jqRtasbEdz4j4+VGcL0G0cd6ctlMD
bjaktDzg5ypJFKr9A3dgTlcBEbEFCVQjLXDDheOdKBm4IhYVs7uYJ4C7zCRN9trv
L7cKovKi7OzyTsiki+ivMjzgeMjy/xtHNGBgkk+ivGGqvAPsAfaZvTdBtKGnV/Jt
IsTBsarlpbN6xUV5elrlF184KDKphNGI+i1jEvUIvMEEeLSMuzMV08glecjyFSQF
vjz4UzAaXM8/xqV1mATy+gywA6auh6XtjJ7y/y1bw/3/9l771VxiT/IyvFYzqWZc
uaSV9SZM6QLRneliQafk/4gPfDkPpMSQPHdFbgYTmxZwHvWBlOKTSe6/lk/g1JBD
+yoon8s8hvVWNYGaiJDgqdWGFZHe3QU50a4sfOss8+wDuMtiWj/Uo5lzoHyyOmZY
oLYnV69uqK65QxC224m+7fpC7QVS7Q5hnBWcmXHf0neaIVI+azt9aYv8uKlPz+dh
ktsIUBUcKVV2iv1vtMTsUauCAMQdF9iZtKKodQrXGVkDaqz0mCWMewc4xm+HljnM
n0aUJTaNxIMbFdxrLLS0hPUbqlE5Qjxdo0JuAG9loZ3flmn6ltzwl32nuSTS5a4/
vqXnrURoQbU4s3ElprhVcBNBp7DI6gp4ZkUKmVKRtsgiYnffZRJH1llCi5fnsFEf
J5hyGGjNFem3W8i69yk8CQ2dQXLwgBELHzTHrBYbVPskCl9HSUTWMxJ88M7GVgxg
L/SWJPUOhriygwjJbWbTrTStFmXlBXJ5Wc9+ivSdIvkPugth4fMLlgS8Bufbb8C8
Cnal2hpK2peuEsAR3MqC3qb3Xtmb1wDzui802Ov1dSoN3jEsHHATTT5DZBLNqyTv
Mlm121mr31b89CdT2VuQ5xLxO9tHpKhbFurwM52tb7hD3/wgT2AskeWMUmp9yNQY
vGzITtEYY5jdFnPeHWXNAZWN8ctx3jqBPcmbhkKPjOfVTlu0xf/Bls//K+lB9qLf
zqjhYF5Jg+/ks1b+AzUglGHPQDzu53He+OpTTz5aeg6XBZegKgDNufnnRvh5oQsd
QAzhSDMmH0vJS6O9jBCu9nGOVps+ORlkbhVlpfe4gOR/4IjXRupt8VWo0uQGvanU
AJdsDnFPvSGoDt/POdN9JqfcmBUEmMd62gy1sufLD2753OuEpE84TehcSO4FstJr
oJasQpagEWSgV821Td3on4izVOijeRas/H+3C/ed8yvSYAxV6bhuqRLxkuLqW5WP
+RAd4Nb0hZEGgxhoKvX4lXPa2YtO8RWHqO5Jr5Mjptwjk6pvqQTczoE50Pe7jEhm
vuzmdf5XWnQEKWPEeJRIN+Cj/4HCs7D4FNw/jqYx2Ui3p++RASIQFXk1rmQdzcgL
hXzYCIB5DTeIdRRna+BfVA/RzmCJq5QAxTMJWqWnSR98nUCWpUzmf4Q7RmN822T+
/G/edx/Gp2Qo+EJwRuJHZ4hNxz+qA1DlWE6oQbm94yEK2bEt3xtCpzNe66A7/Xdi
bURWa6FL1Txhf0R74kECts9qGoEKJ4X7j5qTnav0UFkOslGanRoReEdrw0DZR9T+
qOvBp9GqeHb3bgtPLdpSsNd+2/vOJGGRJwVe+OCXrpofOerXoZZ5dcGzYbVBEL3p
b9A7dDH/5vNR9iFw5MDueTHtu3MhOPSomxh/rVf/hM/hGtdKtRC40tWEUjZaHi4u
X+FQtD0CLGdDLJw/KQ2rBNJpK3DDb0ebG5KFks7HV0KEQZQ4aaI/1oNP17aPM6A3
WZ978aULif3WR/2Tcxz/b2GvXJnuXdNSJymhnST3VqPCgVVZUn9+poUuJRN0ThWw
rzn5GZXxVm0MUjB9a5IHZuTfJALCCD26E1QwyecHMMYdUde1nOhg2tL6T0a2YEjW
IG/RI/M2ROqy00zMBljTaZjQl+bPAxXLVc96bhEQYq6xqUulUgvGrlzakaf6lnAo
Zw5qaOTrc3LUqv8EMnq8WtK4cRsufNIzOSoQbi6NLSKy3bvQEOL0GrMluDZ1H2um
6EcsnNaeLthIR9UPx8m8QM2RWt+g1WUm1CYGfk/7thrEBvV68buTQB+qEZQdtiU5
z8kGhKVU+evBGL5b/3WPb2QfbvSaVAZw8awP2w7vW6jhLGW4SBKCRRQtJ7CW4CFB
FD8zRPyp1iFLIS7rKDbAyCZ2nn480pCpF/FVNqjmvVa8+Csg+l7A5kS7g7E7NdeE
XuRRI3T/xDeBb4o9ePKLZnnzxmPRSBAWimTgVJt2dM4mEVPVVaZkzOk/3/2QGsF6
GnFmdUN3v9DALWA8mg5jzk/mhNG5xpZcpGvKIdfPJMMNn74E5yuTvPS7l+lZtlQT
KuOVtu4Ku0RFz0jYWenMpitT4VCOLD1JEpcn+W18PjnJw88jcCkTMMMOWObdxoqZ
Eh5p2zNbIP8X3NmXWyHPp26Nrw8rdHxxtBFXC/wj25FBxdoEACpQM7PG45bU8H5k
h4w+UXaMEma8hwNmmkRII+v03v6YV859ejIMBLN6UMbpr+Ui7ta42AfNn08IcevA
ALRGacgnkwI3+udIyrHC0HV/Y934U40858rsKzbRCa5bLw2N+sxhtrrJdxIoVAXb
rDQ0gWw8qx1zariuc/QTIs0xkuUpda5IDUdt9XstJ+W1b07q82PWydd261zEu+OG
n6ogacRZKEK60mPlnf3ANneZVmx2p6MQ20NdyIZJPzpscfs3hSNb8TcrEFctp42D
vnRtLsJ2pE8Mpjabmejd1ZYFoGddoSdTDwynDA90f08qIiGYceKnH5+2RN6G+BsF
0a9d9oGXsTYzfaHhp3JIb6REF22N5lKmSLXhXpo6qICJQ+mDFuwekT0t31XfASDj
ac6cckKRg7TwzwcD9vjfPprt6CVrSLmeNIvea2O3u+xoM8OdJ+TGbjJv8tJiygQj
tPdiZFe8tIt+8RhsJOyE81P8qnQaFe/g2ihuhjR84Lz1gqqcLj74VvVdmrQZTQwh
QH8pAey8VtFHOmt7ysLxLKzRHjza9hxz+/Ap1GzORlKJy4FRLmg6Nv0uuQFoL7/8
/wNfaW0KivgnFUJcdjbxEnxxmAUJMJRmRe0eYbdPKVmN29W5Zy++x/RriCLqER+V
5JueCJBd3naUAsekUQXstlYpfVlNyQChlJQVbAtcSJbau/SS8Q31/0MePJYWrsjF
FsFZFoUI2JYgkwFCxdI5CGhd1BI6efLxpC6VTB1jw8KNBpqm1zGR+PF2Je6O/J9n
RuIaFQuwa6xvfOZTmyPTZarl5bwjF37yqmAsuFUY6bV6PWy6ZgEH4ki0pMu29nm3
9Bx/dLzwcNdo6q8+BW02NOifSQUeqtNRaA1w9rORa+eP2jiVywNfOlDMHCzVYx00
xwEbAI2zGc741J3jbk5EUh78F984ZDYQ7AD7kzANzT3+PLeeL6y3yD+xY4LTUxnO
psij8rC5t2S6WI9pa9j/y94595Fp0jVGz+G5gMzQHwaRggjKFTLe8Hz0N7JOZCYi
ezheakoPFZlmvD9jpv90Dl7lT487ZfxzbKIklGAK7NLHBW3iwadD+BkBFb8OPjo6
G5r08mcZ+f6jInm+TyCILg+lUGb3di9LrDDBGC2tFRmAgUyU8G+sI9b6g8mSKDfK
RONhat/XlNsXeMfHTDVwsc53hLKFbsuiaVK0JBhK+g74wsYNesai2r1Zveg0M89Z
Q1ggEkMMyGHAgUIFlSpRgDSyfTWKohj4kOZMJZFG1XeiSMkZCrihwwR3U+8oa2jm
TlW/PsKsUZ/ZxbviflrMZ32G7dZoNnTn0hmtGjMFtxOrwKtbVnTb/BcYEIRQNhVK
Qh0TJyOKwyLYR8oLbIxLD5abntaHwhV76m3N1R2XVt9xhoRqBgxBIMqQLt+BCJX0
V0J3tAo0XMtI0yr17Ccj02WdmfJMDaA/BQ/UPSH1h92uDpGd4WY1RRpv8Lc0mueM
Y8BZKOEPeWHHD353nYG3HsK7PR7V3N/biKQwgoSniDK7V4zqYpTGpY5JYHChpaHb
CWC9nkzt8y05IbP/x4tFTucMGBcb7eyw92c8moFnz9TJeHSod3AjysY1kcayvgh4
l0EITe+fQdrcayS/7QGw+Ld1lLqLfd4kqfKQ6+yrioUiA7zb+5X9V144ou4OMtwK
SxbOmAKxLmEr+yw2ddD+r2j+rtFR1Nhn8ZInqrlkmbHn7PVqH23fZdXIsLYpIlsp
5wA5Kt7fD7d0ef0XIfykA2x1W3wwkwvgm1EX+v2VnMd7vMMi73ge1acS1NuRQVbx
704FvX7qmHQQPkjEXPNeB4gHxPaUBiIqpFHl1sdCtpm4yVBZ98l6Hq31Ssl37E5c
5xbYpcWGFOIORbujc9xr//05S4a0eDW99Ob4BByB6/Q6APIIcFt34XAFelR7s6u8
7AzwfPQx+rGgdH+yxPGNSQH7xkd5JRDm1CGRuiCpdBKre0CtptRKhsv63qGnuaYy
Spkuuo/y20izGCWNbOLOqfp0JYoz/NtkjjsGJA+3eWkEKYcvg/B6WTDKBPCNnhMp
IUqkEEZoCblcobYs4yGvX3bn0Z/3QQnwLtgcdXyKPuW7XJh7Q/sSSnZCJTZ7c3gv
p+DHYswcmr0GLQmolf04QwkEPu/Gtgui6yXwTMEjhuBU8po/67HOxFG0tv3G1F3w
M+VHXH/7ZWtMd3VEK63eVAUwQ9r/z+lZvj1I7mKa2jZle4dwf5v26OxE18cgHYvU
hGs7v9Gprza0OFwm9lIyHbiFYpG5I5cjSaUfWsgP3bcMh4JtkTZIXk8yHg6UhucH
dU1i2Dbm2TNqihT+whQTddrBHiY0vYCFkEaRg36ThFV6Rxx/LerLMkl8Rgb1efMy
BiZj+FMA9geUN8LpGs/N4ES5WiNwTdbArcij9DQ1kQ7P4v9UJmafTO5FCMRnVi33
umXxqqVERCQ3Iv5JZNlFWxQa4XBNa00W1pTjv/nUykmffuNxa5H+Ex+VxSi7PYdR
0b2Dt/JawCBiQTEs4PeTKkg6yi0xldxVKJz0Ays+OKaT1a9ARz4AOAD7T6+2uns2
GkLzm6sQsQvzto5WurhR4wexhtHH/96WXylyEWg8HAQ5rZLY5lrmU/a/Dz4Vac8D
3tz85mFAWCPyqENN9OetbZ6ab2GW6pZAWT/23cFCfEi+bwhggNBmrS6myJ2dsE8Y
CL+OUnBJ2aLY2q3vRKB0SjN0m9OjMraOngKILlcjR7ktB/VmsQvvRtuVOYrhzpGJ
I9eL16fug5l/Ju70/jbHuREuv4m69u65kxLjNK3/sQCQaQtoRK/d4dvT9wO0ZQ8E
6H5fypD4qmCsU+7llzMLGVEjwtyioDbGg7Y5QWYeQqNk0wSzYpPljWigTAo6IVtu
5p9zhKo4vw4f6fPbYyLABontM4lUrqGo+EzuYixHRgZXdLrAegA+U9u3rsOBljzf
FUnaSLD4b4AaUCSHRv26GIfzG6L9qw3mr9uSPwbpPM0KLneqG2kVo/lODjQq0vd1
ZL4yfo2Rp1VaQqFCYivgY7k3jEGOeVxee82OfgYEVPjKo88KiFVMP1LZVcNL5gMY
43mSn98SzJihOkV6XfHfZY5458dkxa5uhJRiOR3VryOU9XGHtP74HHqd4zZs2cMX
vp4E3KDna7rS+K6CzjoMzNDw5SclO0bZ9o1LYrWc9NvtUoNA17xP3F5JR3fJ8nwt
+j+3c4sqmoRLCGKgpcQHGvhlEf72EZiVnqLBvv3vzFfV0L1Mk1XspOb0plwL5vcC
1hRARvFpESH5sOQFkRRE/L4PynHoGu3Zv1J3EAA7aHPCJnpQRa6cGaHljoV6mqQW
h6DTV5vbbpob2mjCY9k9RhEUqUhmgJhl3i5guLcgN++hYAO8EPuyAJz5/tzSJ1nS
u32C2kBEOdbiL+taMQUuSAqBt8Hb3H80n/Hz1Eus7y5eYvC3RIDAT5M5Hh/cbUI8
bE0eewtlO8XXuv7cqEsBZ4yN+57VcFsPD7E69FBoN4O39BvWU3S4k+NSYhnX8+t9
+pM4x3wzRfJPnvDZZSK5THvhpzJ0z9Om3wSt2+P8jkB+BKHuRrYoEbP7FnX9XGX3
7q6uo+PykY4txpf7GzWHDG8egqgyWe/MYfxBxVibQSkkiqm1+sHM5xXBE9RHuuKh
jPREluS4mCPat6Bzy6nBRuUCBEK5nsGIYgfzucHikcguuY2kLL6OXvM8Ndr9iVpV
+fCCgCtTcqDNpztpZNQ6hAsBYKkPvRL1UxpynlUHqRkYi4DgpBL0rGdopa/s1Yoh
KmneTxIckcrPn/4gNxUPQxa1f7bJHNtJOUOLy7sOe8BcRwsXX9CY18QxLFWSqSuU
fr8afm3NvLq+SUCUmlTAPgZnRsE+W0OUZqVQKhHKY35ORTs32KYybRErO7m8ZK4Q
QjJHtjGnM3GgzmzoCXyRmYhxDWNyuXTmGKs6AhoIj0jbeEK6/VaciK03Hw2LRFAu
t/cnu81WVnY+WqyZ/7rjn0h+ab8YeY8CLWzf6u/NfMDPlRbsrhVkpa0AxfgCZhO8
bsDPQow+FHM2wqsauEj3dSudSnCHNvXLZojXQIrrkHDPf8WrTF6EAgPmdiEzqIou
8LM5CVu7B2I8mCC+mQ88p6xgeuxLAQtNxC1Stej8T0KejIrOW8woz+PC2PtVAYF7
HqztmYIZE4GWS2IW0+28D2fj/KZYyNHjWgm0JTdhqkCD5XZgxGCjX69cxf2DIQFv
oKstSPqydJ3fcotXzYSBJgSPfGWfljCkEdAbs8ZyxrfbQHdG909iY0wRR8kyyDGd
1harTShK991e55Su4vcbP7KSKFcVPtaxI7a/XzkWpqOdsuHRPpMlSgiym5sGxKTx
8XNmXRwogaPThIdT4Tp4lBgqFnMJZrQpCZCkH8wPQJ5OggTB8KsVZFrv+rrCtRBg
N8C022hYvbcoqddJ5NIYNRWwjF8KqUwRBGpvt/ZcJOAV9dhQC62K9mAnNVniY3VF
WVEI5vknaRHItePIL6WzfJG33gigA8mNxDgmFTcuWeXTBMIuTMo1ywGmNMAoOSZl
gP15ZJ6xr1GUA4xMWGpo+J6ktfsvDqlQuLNQKXi+tCZOMNI8R4oHpP2adKlQhvqg
F4ic1ZmOsCG9ZkQWKeNd9zOkm9vomqBj53FOegf2CeHsAkGXV7GCwpGMNsxDnMHd
G9GKy/79z+rdnyEq/6SQcHz3FUvJXSkyqGc3appQukmYKK1+oCYTPNoeSpKG7tSh
9FZPVDQ67xJvk2k5d+Auxj48u5f2BN8zAEIv+yWCbbCLwfzvBqjqWmHN6igyvwBj
g6wHkKUHxSkFxgkQkAIQFShrMYoVWfXqP5HbPxEl92L/oFA4s0jGSrLbuoA6+EJ9
FzuXHm4nQ4NKU2ufTYyeC8FZPNcJWzOJ5dDPv9wQcPQErEYbNR00QSQwvV7jIjCM
JinNdODMOLX4ChgH+SlWJVtR16JM7PLMYMPOgQVs5sqgG+MVoSUxF5gFgWXUqHYL
LTIujT7qP7ny3bSEOMcM+Ta/DxjQX/zoWctoHdO0hbeC9+aUsUxVT1joJCdGsuVL
3PzVqvqFULk7SXZ3juUS1nhEPQj9HK2KHwGUcnRffBeowbNFEPsN9D8HjBx3I9C9
R0XyxZkFDuUnCDf/06qXOZ5vwbNPTuYrjhNA8cOydC7WfIcxndjlHdxgP271dUDj
0lO8haTG4BSOsoKLrZsghpKGMLy/kAPtYtewrWN6gv8h6pkLqy+UVShVKhZNdQKn
ahy+tqzk/ienhZxsHj5zdOPWwP44QaR2H0xJCnKiniNO9PsCUzSxQE9o3qslj31r
9kQaH2L0UMsLB+GZftfb5Kjh7lgVc/OzvzOe2ZjVEod7Zyfmzp4RyB/c+9ONAin5
2UXff2i+gWUBaeSf6uXTxW91TamRdInkheG2dmgdq98QE+WlDoTC44sRTwzWBhEy
MvqcAvsqami+4tp/dxGe7MdqYVRIn8JAfwp247vSuEzu87zvh3s/Bwn5LJdckavv
3KMxmqgdR69I+8oTTfE2wKj/yl2ExNajVYaxi+eErfeCjmVvbLqIZVYKzZ4mdI+H
kGPKCVixRteJ0p7j0lw7OuMirToy1TozjkUBRbYZ7mY1twJ0dTOyDpbNaoCTyn+0
zUqU1wZGdSFCJmVoQxe7lF20T4Rs43M20XzoxuoaaBx2oCe17gjqrJdfhkXMdneP
JsjVEVWuYnqD9Beg+frfym0iPc9GmBkPmkrtD16ohE0plQtcLS7IjlNMk0aXl42K
mg1a+0OTtx4zAM/RnC4twj9QUN5m1Tj/Pgg/JAYD/dj29o4WXrxbF9Ku9AbkTK4B
uOZ7asr/iRCy3JcJ3xd48j0imFBuwcKY0VPgvixqwe9I4VBpeJuDFFQRcDH63GRe
Jx4GR3+yqPuKOJKA3qb9jocMO4lq8W/O/kUkJxqQ3+8vxFqnMwg8UQz+BnYLDerr
jqRhYXzU6EJIx4jvSx80EkB2Xav6jk+4FKkR8/uxwn1jNnQL44vfZhxF2OVsgxTb
6JKvCWXEfiBNhCeW1LBZQ3NQ33zsEQDaggX+e6WQ58yGEz9kAC5gFX1vYFy64qbL
qj757DE5y6pxhsWhabiCPzCgHiWXUvLcDElzQgSAkLRwDoQYc3eT6weJZEQ42PVe
IwNL3R0c3omXltako5y5yJKWE8z6VKIxj9sl/dXGWY1Zhy5tXJKZ4+M3HtqljESR
vmoq8sUr6AUNbHm4e0l4IU5mCRguIt4FaWJp+RMDOT3qNahtfkAX9veEaY0uGUzx
6016NS4/N9eaXTRil/9hU8CLMDzizq8uvuiV5OZU32TTqDKd5XL97jSPSdgPeweP
l1JmpWPt+KloMl9NbSALi2uGPc+4zOw2NFC8t3uhMOrSgV1/wlyFASleQWxsJB+B
Ov/Rp8CAtF98MDPUXKcgZ3R4ghQTdNJeSDdxJIhL1w+AoFpq3pulsDsEXqk5qrrr
ksIm59J0Pza1mhmeg7ox98H0avt6yiCVUpfdgOlR/0OgAUkiFXtsdxzH3r6gDby0
ZUDizHJ8NMg3jNy9ownTzAHi0L0ebl1Sh5mTdNKYwnlja0Rbo0NC73zeGn9x8tqg
eQg4N3ZBXokL9sm1Kx7BN4LqiZlftFUjOe4h4Oizg8yWf0da9P5cbRTHlERGfYUx
1zSb/sKT0glV4gfV8HFIzTHlMnEvDB9Y7UqS/7uEVXISjSfKy3BqDCoeHYMU/BZp
rEjUrr+aIv808825fEL0y5AeoFzivzydBo/2pitcrQAK2xmOsYEcidQZgDKSVfSv
FRdB5L5z4O+1td0MCtO9tDWTiaAiMdXcXKAOPiFH6fFtyjIUivlByD90IHGvbctt
lbXP0Sq8wCnp0I2vBU7ZTdwYC9MR+3e1iA0FXqpOEULxcSF1oEjSjHLazgvFq44f
itVT+f4k8rcw8Z6v5vz/E9uF/v3+ju+uXPN3QjqEgKZtRsFz+pJEppsdyQR7iEAA
1DkC3p/BPAqG3D6KjsOYzuw2I0CeUvXLENAuijqTlXp+cFoJ/rsbpvK7WapeJKkD
/bBHoddUSP985rsaFQUgCxgiDqQ3MbBdIDLLZuug3LmUqNKl5X9iomcoFNoetCNw
YhG08VXkofChQRn5YaaiNA7e2k7Qc7cZKOHo/q3UItzpR6IAdYXF16JO+LY4yiCT
T3/rK49u4zG1FylrxBSPqp5PMH7h8oIpKPnPY7Dfyi2j7jTEOR1pA7A+wbNHdxfU
ST8l4xnvpN/3Nm2Huq8NE1rAQIRgjRs1ZvCMJgNwKvMhGczoNnn2p4552fbK1TIL
FedD1aZVhVJqnwYwGowpmi7mKxkYMu1cYiNhOh+VnMTwXHOJXtDDnJ70YLjGynUn
ozZgIDzNlW7KR4IXdHK6oFPQT2ZmfVePLYaZ9LA7vgp8izbF1YbZOZQqC2qadGWK
uTmAWGQG408XSSSgvXuSzXzZN6JcnQ29SgVKr7i4YuY8f2AzQYCko/xhE2ezqAST
20UfkIjJfuG0QptbPyo7dODHR2M6vxcUqhBANlitOyBMnXvGrRUQ3fMzW33WG5Hg
utSl/fxf1+szaSDETAf8sbhQfJ+kGz6MTyNbV/z2pDqblAoSNcMgmS2Cfj6CKNFV
fumiXovuxRgF4eL+FHZeLzRWkecftYoqwDNmnJVKKh2TTZeom3UY4kJSRlXE37MD
TPT/1HHJbcED7U9kFV0mgtdznk1B3A9Wdv0Iiry8JHYzIksNJ/De2X07Wp9F+UyC
0HAu08mXxRH2nghA3pPYv7FGBuwpme0vXkpJ/GaLChNnsA2+dYjovyz3IiWqs1tb
y9bNdIKlWFulFYYeGTNjQ6NyFJgdi7cLvtbvRwHBqaDlgH0MDedkAtaus1bTSUPk
EczFWJgVq8KkdP5EqsR78TJRehgQbhVPpu8G93mVgGV1mD0VrnDg53XeCxontFlR
vckrAsV39nn/fP39zFC5j6wrsF++Lt5cGPDgIOOAslIxFUv2AL5HFx6IielSOrt+
ooubS9Ze/Tv9gQI9WEps4jNfjMVaOnbK1kwMidUUAeyexH3vt0nwGlyVyGi6Zw13
7xVQrQg7awJP4R7dD/kqVcx469ftPB+uxb80BnG2lniSDlHwoc9ItBYAm8D67Kzb
5k2XNoGEw37EyPRXj1h17SAlafpa3SKcsTnW7R/15oukr3meyP3QW3iUKJc0PN82
bGrtQXsVufBIXwr2d2ANrASUlnhM5lcibmXqzae1+ptGztDroYyjW+M1SjZnu6WZ
/801OEadzrV5hEXBV+OcOkyh2uxkCj1rKksX7Wv0tdg50IJ2F/kFtZ5sVyGcUcnS
H0m4sPYEJbcLOWByRQnFRy6W69EQQo9q7IrcOs7Qh/aS+DBiZyRwX2vJYORW5GvW
ZzYsbdTXP9NeiOvCKkaFmg21fwskUYXR1fslMpfwd4gtYkcXZS7ZXFv6CC8H+gvu
WT1ORNqv2GKuxDWGIOWmk9eogF4FP+0WUhmKqzoPkybeqbXt2hX9NLCyvnJ+dGiK
zbYVdMo3gMBkUkoa8fdG1hdrWm6+K/urNhppB7TY9FmFxEtCEOu2Pk/s68ujHY0W
El4daLCDf4nhf87ejTAptjBum33M3J4nlvooL5fGq6XHe+SbXaNSLn0QZwRGynB5
4FvVjNWcSbtAeYvaFapJ1uZn6O+jxtbwAsKbnoDUM/sMl2fPtUqqhbaUgr+8haYy
ZB1cF4j+9dj+nQ/1r2lu43KfOo0bDLx3k6gpWTOHxaa5X3Jtmpg5iN2Cqe+U2SnG
cnscW6FsMWlGmv6HUHuOey7u/5byrE+2M2qPSpaaaMVsqbGLGtVX/etaqFgA/suP
mNZVzA1AUXKFVCEv5tZSMePaeXcf/K2efyTavvn+cFn01TYwNBjkqNnwJk3QvRSh
r2DJ6iZOswOn8S/BrWAB6wmVERAXBADptHEyYR692TB7njMhsAMLYE3KcLpihYEb
vXwMf2/agjqoMf+pXM1AZVLeCfHs3PYrmVgrqIj95OTZOXoJ9kgu6SY6vpRzJotk
gscY/dFeWWzETq+Y6vaQ+g+hFEoM1WlggQR76gbIfuTcAS01er4Ck2MsaCTl06xV
qJBjzo9LhgSclCuJCA9tujxc/lyvK5yCj5liKU+jhJzSueQovwfvlFDnP30eIcQQ
hCVaaj5g7BIx/XvqMg9xaEpbpnCd3RgPD49hhVm6mWL46iQmoiQ5e8r9rfnYU/lo
Rbr4z1IsKf+6WWyk15dRy5d1wC5erMzIygG7Or9utQVqX2/5adZExOaRrphL6Fd7
NyqEcujCuZqNu/w41WvfjGig34fh3G+0W7vuFUfDdSySZKJA0L5gVNzxQ2KES9x+
K1YumLGM6iynvqaw1HFXRYYLJeCGeqX4zC3NF6jvkbMW2sBFsTfahjE69a/uSc12
7lm5ABPeFD6cDhjf9jgzOBIMsc5gtAwEGiPb4HzRs60fYV6hxFnKlhkDdcE2dRBz
FB5JmKJvVqoinlxPwZ0+XwyoBlJ9IrOleDedYWMhLCSIx5RHqVYXW9YcKTxZN8we
SIm9UHfCS9xIV2gtgRRlgRbrwJqO2qHwjsuQo8TOT1BMD9fg5VHxqvw8Nrcz2Vha
vej5caxlariAGRUvuW729KyhAIqQ8rwlVjkILZmVgp2kvZJRXIrWxdtiOTOSjEsC
BUIGR6glohHiG4GIb5ykcEy2/OY7FuNOg/DxlHchqwWxih/z0r052vzolnsBlnMa
F3nxmPqx7i/3TfhOybQTpQ8NbtSGmboBcu2Jzp6gXFrkZSyGaDlh219hC3ReDIuB
EWus3g+3Vho0TJfwz+8DaFBGNEdrU9s8IJO9HvPSgW8ZIAPtlbO1FDwdQUQ33/aG
+1iEwuAHO+22es++E/zuQD3YpxOn8DS3LFcMT8Kg6cmAZX2QM53g9e6bRRI/nn0u
uAxTX7Y2dXEYLYo9GPjfgdZiPHJXpdL4mDLiGHKQIjGozaST/+dURjZ6XQuXxzzX
fcAtp5Ryhx6KlcfFqQ4z0tWOzC2sc6nxRQI0qkaw9XA2RHu4piHP9UMcS+6gLBzM
KH2LB7m2G/hEQAIowWNNuoXMFTlWOfKGtrZh+3jNTM0Fb8IXL6T2LH/RYgsHsFef
0be6N2KQLm72+8y0HBdPM3ANVX9t/Yre2id147/xeMWsP8SeNg3yWpjO4VStlfch
DtHL4IsiCbeT0b0hoa6rWoy+FOIpRKNrRp3s/cHDaZ5KpsR7Zj4TDYCL49dAWqpV
ovMEcxCoG7KgtCstrzW2OAWtDbhA/naY791D1bbt9DYk0MsMV3J9O+3fBHLXVvWM
mYtxFlj75DWJDyqA+mlp1qP4f0U3zNrsvhqAVPnVvPH341B1eEIT61o6UUhOjFQ9
MbPuRUUHjgEB99IwNfNgITBQ1EJESjX1j0YegyZw+5bJWumAMkbnzF3B6MqA0VHW
AhUyqK+klo2/4tMTQwDxXkV7TlBWBsAVNoAemTZ3KyypmMgqUQ4KitrkVwv4ti/h
aa1OCfp6bfqYnjQUxMZrUgLgzYEo3I+474zD51SONirYDahnZN8mkA9A3VL8NHGD
NIfM5/FwBuYo8ly27e7P9EavlVQtIpYn63AP/9vo8HX4N/U68FiIn7ocpcZPbtmV
InczxVToWMTCLcvJ6+/+7rJEVoK+38OfLGP8qmn8rK4gOcq9udySH3LxcEzoPrMt
xISR051PbnEa/aGWgjdHuy9I2XDcw7fWz13Y5V78S+HhKBpJoGCnJnlc3YjAfiGP
mQ3RJ9f0R37Jlz5K7574ROay5m5uphFF0ILtzV+C/OxLPnfgm8rGAgstvwqeNwBy
I+jFRlQ1B/m9chLHYXKADgt8QhG0vaiaU52PDrdhgEasHOv94d/KR4Wse7aK/B8u
2n4NlQOE7wiW53XhVZ4Omzh3IS53AsZWC07wior+nb52TKungovLWk1JfsSGDCPg
iMgbWVaA/c0ahJeeAY/bvu3FCWp29a2Cis019vkdNwO9fhK0dTnPgBFYHciFyOjP
VTS1ftHwDAzEL2DylGGWJS/1p587mMlRljS9W7wf0CcyLEvKrV3fbuOEWO7aL7UG
s721HVldJ/qDr8L7H0gJALgS1Y/Qz2KJufHJikvRuTwNNaKBXhPGy4NUPeYw7pV4
9itJqRILdFwyQGBVnoRddqGBaz8oNHjh7XVhq2fIQIIhOQq0uySleo3lK7Sd7gSe
eChOZtEGE746lGMooH5TssBg70pFF1jGu3ZYZuP27uaWIJg4vMSzfyqMsUNECWdf
w4x67WGprq/vHYN/dws1ch06e7iD0P+s+8iFGy7VFxfmfGFdFPPwbTOmMuYVVEWI
BmCOsYyFxnkkWRvmMx2LJj+uIkktCXlkpAfxyB66VjWyIe6k6FinUb2SpCvEBo9N
Hh/Fp0wJUc1Zj2jfOKVpOIzHpncUfC/tSpFNMFCLqFetKZp883j9OTl0002WecMh
J78TMWisRrBaA2cQE9LOzExJvCg5ccVviJIj+l0x0ORvAAKu/MAitN1ljidfbEIf
vomeRsPtjpDEy06DyMqCQ7fHDeYajNrpwiHO7xmcr8gfA9+AgdAS31Qm1DniS/44
GGM3JobgkGpCydGH0w/jJJVuqHxkdCY3qfFK1PzwAYynRiIoe4DIV7Y2ED6KtSUg
Mk0gGP943LScTIB0Utu4YgUAxuglmyn0I3y+EGi+TsruJ/Tf7jhWUmUIgt9LzdSg
iPNi02PpdVxeTS94rcah6t150ATI029c3BEUtMvL+A2hO1JMUT183tkUALJc18GY
/KuOC5k8BITxilFe2BMFPyvTuRSsH2rKNpLrElpkntyyilMoRWdbnV8jnnVtfNe4
Jmgyezl2/XqSA9zBzairBV99cDfvGpTPgB0Ur/P3R1jE7SyqoAd1NqeyJKPeHTp/
3v6YeWpjDKeiXcaTZfOc6dqQU1iZTwvdQmaw8qynhfhRAp7ZNPlNh6Z5+GyWzj95
V184HSe51iYyLIA/q0VBGeRaoX7oLXl7hGcYQFGJfrZhB3NSWUBgXjIvhyz9GfRu
HMDR4Pl9aIIijslCzufEUaao4ODyNoAz6MEXN+C+QcBiBMzWwUk6tx7yjVgWy/lS
Gt+48TU3cT9QnJk2Uks4qijilruwBuPtsWUtGVkNKeobgwVKHHY8ppEkOEeNlnMj
mA4QltWNkcxJqGJDWR1tLkvXeqVfQxK/rQrcHVDzwSwkklwRh5XOVHbV0+7zSPrE
z4cpfU5i5FfYXZxZgGqz0snkhIwnd35dvSYYI6MfZ0EfVzXXC82Weg+wTmuMnB80
zUKrMq9luVMlsCm8JHXd5cVpX3hW3Y0yO7b8CzIX2y/V3XfLThhS+G5cCDs/8KbF
rbYoYvSPlfqWwbXwBalFKaVP2AXW0UQ7TvhMu1c4euisTs7j9LM1PYR5Adq6eCWV
AnYCh+w0YWVIMoGh+dpu+brUNgsSug65ZDMTnC4M+KE0xSNIoOFC9RLz2Z6YnIGH
UfCYXNlOur3D7EtPRaXioP/7JrhviBamv0Yu6pB3r9E0EGlOmvlWOeygngUicydx
xT9I5ckFyoMt4O6ot60xxGiAiSARB4qjXfFRP7pyhM+7QP3r2eOAXYhn15miN0Kn
HNCFJlaBJo7HD0Jjeys+6JalvIuGW7Th+HxpJV+eueBLikv/A5Ylj98Twq5Mxijp
QpabO/Hg6gT+5cKfSJCIoj5/Qe1iTeZKEVcQ1rYIP5fY+uUIg9zzlOL64qwNCTEu
62E6yDM5QM3rLt/5a1I7YqVkjtfesJ9/NFAC0kXkyfmCokrMlAdRj06cuJRxt+7U
EqZXnnLLC2gExaX35LqRqKwlT6EJcue0ecSBKkQ/TYqcorMKdX7PAiHdm2q86l/l
L9T22O5keRZNihQ211HBA8uednmvJwJB+sKP00/nwYEjj9PAK6HPpt5UBXVxtWHu
K6BRPkkHKfZ9DAD9lAHz0Bm6b0r4EcaH7y7wV3G7mTW0GBjRMaLj/lWProi7Qu71
/qVOCvVRtMLTB39kWHnXUdlubbsr41NAILNBvSZI5uE4B0q/Pw6Ww5a74DMJ12s0
Kw6TIEwk9nnF/3FWg5wri5kCCXF5p/n36atIQ36BCLoBkN8Ia//XDujDZH7/jJdj
qt9ZdZmHUlqH1ENunQNm530aMVTiuY3OwZQt8kfeYI3/QQVpF84BuALPMc5A9bWJ
AjtCIlnTJ1P78abAKkgMbvuOTZPcL+kTuq6i0+yJviEWPq2G534Mnz4VS9//Q+91
CgKQ71aAtcDu6/lXBJZR6nZIer4AZOQO/uc8Dl9puJRh4R6TAAN5nD2THIwAKXSm
joxWWS4ucWFLlYvGa6u0lDIu5U9fh9UJv3t46Aom8S/GOYl1E3T9UM2FaH6xKIe+
mP4MqLNDR/xPDviiBQsbj6eb2I/R9/7OxTQKrUeFuQg7jUrDU38cPe/Qhxn+7KJs
MJBCLpT6FIAE3f2Ji2wKCEeojM9KFTtI7hAJVjlc8iUmhv8OknBfFJfYtOKegHc3
pweT/l++htAfEPA6oAC+y8EM+NIZrndtufMDN93wIjgCgPawHMKHu9I3/GC1q8yd
yPEWt1ezb7TNj63BU1V63Zk8pm2QFyqxpdBrgVOq8AMDT/b/9yy401fnaL3EgxBl
Ei1LL7dxOc+PA56d8+5/0KNmaLNEZ1ZNTp00mzdJrVdEf5oRLLnn/XlJbCtFdUgf
j3YxniwqfYPK9BTVmAk96SHNWhq8BypIoCmCAV3B0seQeDn9AA3x7l3sRB6mRN0V
IIXQcyrffqTqtKIHJXNHGSsCO/SytK3Co57l/Cin41zfW5Lmpehzvnx9/SayFu5z
Tgg4JMfJv6GZKZGKZ/TQc7lx8FLEBy7bUIg/vnMFtNzfy7l1jeZ8ev+cf1fJwA9O
bTpZ793+Z5TUww6cVDA8nYtVZFM0cCY3vVNBQxH3aNEUMzvrEhesFem84pi/uazo
HAKaFra41WGnNy5c3Ajt8qDaYeDwjvjLZz820/HD7qMeuaUjgELU2KlTp3PSjND6
whkSjA/iMdaU0uFwqjW9Pf+EamPLmDWZgHPkVjAWqj9G3NNjbnMTJyu5o13Hn/v3
cmC3akPsJRvxfH7EkTkVkD+EcyiCrFm0RXBMb/ukVIujPoFSiQtOu9PqRciAqyO/
P1kBUU9+t0iAznfqT48Icvb/Jdrho3JDCf/YG/BODShRgdm2dWt1opdMkZ6j9ulU
O14RFKyMC5yXzGQ92zHZ600+xcdReEXkorEeP/GZfd1B9+tHBRk24pJPagbn27PR
z5UfNaY/lXlDX1g7So96fqqeZGa1mXb2jc1XqP9JAbcHNTdxj5JbxipKDgQ1DVLE
lAK53NMd82369Tro6k7PGNP6y+h+sHP6Yr8LbuhwGoBYMgc9cMAj8Kjky8MvPgkI
02UJe/gFUbu1hNjl8VidxgezzYGbp9JfGNmpoyC1jWsroerFkbFMeKCoAuZ4TtMJ
OjZB9NUSXMD59UdAVZBzdZuCa2ZRKzEWFjQpp5UBhiKNAm6jgKO0kHtaKAZr3yAC
+4l57QKtRt6lVW5wJrcWr+uOZp6fN9q6LrTu4KWviGIB+S5WjwRL7sx3m+qXYFQc
qei79fSHZjQR9uEUKz6dn4u0MkjBRYa8JhBshINWf+G/6CGUrPSbEephFFIm6n+r
cT9aByijiF7l4VzpQJ5bn+OvYskVa8EBZ1Qk+GqsaWHxuaHMhPuBoh4FNsWzv/ZN
zneGDzGM/dTyYzwoxm+N6Iby2b5FY1oqBXBxeRCUgMpeKQeh9s+niBHBXFsab8XN
HE6sC/iWnC5/1jWIBnfAy4roiiqcrRfXZ34QusV/aB1h+hRRuuC1mmcLqfwH5vHf
COM1Rdiq8BOfFvSMaVYs6N5r64Wg2fjC56wuAQJgtpH9d0jw75qVkKnjnuZ7ZZNQ
0lhA5cCehy891UKDdZqhfGVx1xOuo/sZIYSbJdornV86v3NrlNt2fIVv04DifjZ9
2WCIQ4DviL1UHl0SYK/WMHAS9lc6yUKVsGYhGWM2ADmay2mKqUx/Cgax8gEPNa/i
D2PVH8r/HOH9S93haHoW1rkJEHRlDUAt9muK25rxprikW3WPp5E0c88zdLt5PF/8
DfgFJKXaAvMWOeWl4NEwb4oPbH2xCsNrQyTukbdsF4apCkoo2NkuxHMBeBwDiPXE
i9m2z4r7bC3OdlS/sJmV/WDmWu4T2naDQfX/zwrNEypocOeK1q8olJv/7vZ2rzGJ
lljL+fpL/bOhHKSR01fr/cOF3rEkssYudumONBsX8QWq/rYThpPHT1orZaVAUnzr
QYdNHcYQFgZShpv0gSUZJalLmRTNbJqoivhxc8c0CnHEx+7harBn2t9bVZfoaSX6
ueL2S/zaiiGfDbIBFz2QxEpvoxGE9zGQzOytbwPGgUwX8dm7m3poLxDN9FjKiHAL
ZrwtQBwKQda28EYOPTr+tri9lPXF2KkxDBAx1CT2zfFjYvsnjra1/EwGDJScOPrs
xIBxkOGccoJvH8sd9TOt5IzcX1QcQF6JTKCJu+EmXAeskhV+9HTzuRm6c8565noI
8+wajLAfdWx0rgwmquKQAUZr+Bl4GwOiasiCmz+XZRHL9ysvQhLBLhhHicKL0HXY
3jE42XFsU1Hv0xMGgbhFZmvzZenGYWund9wlKLlMaHEzH4etS5j1enimgVKjfID/
+REhd/B/KZeK8Stmis5DGc0UBDf2kOyU6IgVsod1andKMv6MpSOTR/pI7ZsBXOG7
cUp3buQyc0mXe9N7cEUFd4LLa/LIPftFAich9BmHfvxKhQCGauKAC2mCNsIMk5FX
nl2BGOL/YMMvUQFQ6i3nWpCD2XFC9GBOiEoJ4AKCpGVvBsTl2NSCVsNUgw2xw7YB
OwUuy8H4y+es/edYXzOoSDTME7pI4SU3O6mm2HnqW7cE2wmtUK+vjAkYFA167oc5
iloXWIjXQuz5U6wWw7Qzcp6QTbfkZvMdNFz1zunRsGX95Eo0tYfB7nux1g03Svxs
E5jujMx7TNJeG1riwjxj5HA+ZIu35fYl8mtleDRI1aCFbnDcpJiKRCy5seDgcUIE
YF22finhe9NqE5T0hWTlmHiuEofH0o8dxgwEClHh9oYBup9ZNn8qcyYXNIRd8G1p
MRo/WmmWwWskJcxDQwANXUMxHFAgffqigWFWFDkCHJZ8f73YgMFuSC0Y8fcVpIrN
1+Ot7NaQavdOhzUd0prZPTH5Eer/4P6BpJUqTO31t2Z8VDsIeoYBXqCdf82aVX1F
5tz2na1bt/DCiGh94vqwisWbkQqK+AyX+4yV7e5fsdnNUgfdKhZ+5tpZdptVXEmM
FBJVz7gbr24H+fn33heirFjjkmuFJO0IPQXavbCWivUw6mJn19PbhO10tDbcecYA
7l0h1BFHf9n4kez+jGWQKVYKzWzJ5woYz4vQQRm6QkNFugLLi6rM/NpaIxylBEsM
LNHssmNDCyNUoPlt08xg+4uCSwUEkZZG8kcuxXqBN5jVjK/oovo6FwdU5RTYd+/v
IJqFeg+L3am2YT/SyiG9NWPELeyZWivMLiyFHcgA/10OTGBuWnjEcmUlESflIMHE
zxBu6FvrkDKofpK/Ok94LOKZJeECRAfqS5Q1WChIzrTyOSKIY9FyAwLcjXlw2TRn
pFCi9rkp3aO3RWsVRvU5RoyC3Z4sH2KMoxONG8zWH+TmoKP9dkMZ/9m2uM7kpVxV
yrsvB2ii7im+y+/yNxq0w5rgoMHTHrEOWCLqcYfps5oF99neGntfWjzBLbxfAKCb
tZIiEdTn0EmO/iyRGGeCGZnOCGmBhSyee8bUmAYO8UTUoZz7COUrSQ8qhxyJ9d/z
N6DoiLXkqSBQy7UIGQ3dzIJRUePn3ef/GLLIFOWIbrKiVbzfpr5bwzJARq+toNGI
DSef2KpNS1a23sVYl68JVILlujO8f47mvz6f+OAYJ/Y1YRTsV/7DSVtMqkoQtS9f
22Z6iGqXRMgPc3pkaTYGquPCr4f6n1mAOOcvdZcku18C0De8jhHLcoFPpX/Wbm3n
Pdbov0Kb48PZdSP0glGFbmfFfBzlgNY/zD3gTSkHuj2Mbq+gDX3HE9FVFr0qZm0q
LZwJ9IOMJ2nPMLyzphM0vluYgs1sQHf6ApRy6xlxIetPwQrfPvoBbgTldzTB/4TN
Z9gstC8K93UqCNliynjXj05HV7B4DG+nFxyD9VAWW5VFmj15NH7xnbbCri5idNV/
5D6yBUHLFyAUfmkEwXdIs12wDR0Rq32m4rP53c0G70+7wI5UuT2RRPh9l763qLyp
95Wu61UKs3Ut4tx77fhU3lQ54gSEsz01CP3BCRoXqkQdn/hpqxL0kcLhAx51eTXF
dO5ZQHC0DRn/p2Z1LvRrZL+JF6akxljehIIWprNMr4w4mUg5faSDCBxAdUga5F3a
4AttAkwQOH9djPcruQFaNFzppCFz/3doJmlZBNsLO97+6JRZB6kIoRjNmccFJ6hQ
B/38SIWfk/zRfNLStRNiJ13XgDqOIfpmRHOgcwuqy73Oo4WRxdCJDBQPzxSJgw1o
R7Hn/Qm4YH9YYXtnWjc9BnZlRgzx0/5O4ZTwz8gDTUckNRrXH4fuHrAy74VjhhsA
srO31g1jMiqJVdMyB3MD153rmF9T2mNizdSWO6400mEO93FWd+jcjsUaKZ/8LjhB
bSBHbrVS4OJ3QyVWCMVp8rCYUOqh7xopv8FbidM0FB1dBpyRHpo3kyujYchrB6Ac
Rgp73MMsX2EE1czABhL6qBqlcpTgEVCsQSdkkEbbVZWL5C0TleV+jXmkFwE/nRx5
3Uj/S7ir4pRmFnV7CqUEwOlV62O6lArt9Yjb+QqUeLAUepLWCvoITS24Il+rZL0I
WqMS/pjw8fXOtwPMbZTcK426K5KONDLnqzzjBnWjDxgBzVjSMRfWQPG8d/cCMYkd
cusqE7R2pg4ZoGhjfdU/5OSW5y0qg9nozQUlYT4YM7hU+ELPkb0nfIUwgaHsZl8B
L/Q6kZ3NNlsYT+ROgIyrW3wBvtr4XdzhW7FMBzJFIoq9LT/B9IJT/Yb/No7xN6y/
lfjjU+j8Ah/8NLwsWCX7nLEP1NDy53BdpjYnXtA5g5KHFTWNiIRYgy+1+YV9X603
nxeRBegOTfvikP8w28k9QW6fDhPD/591WFCkbqPzcXZoP3w8iXNxPO+MI5tPCU97
1Iq859mS8wq/rwkfGSahQ8zE84acoaFUJ6fuZeRTaKUItf9X8OQGmn0B6xAgvzij
gdzXiFmkJXCOfhCyBDZc2Xr0yIvF4TTfrgunNMw2/f+I7x15cyNGlafJ3EGc+rFQ
xGw7A7sI//bBrv5w9up+TuO9dzGxP5aj1k+YicIm6q0OCdDsS/7/InJKdk+BKXoj
/XSR+4+CtrWfH52Ba4lDlV9vC9uw7RW7Stovrha4L7UkS4AcSRc5X5tAt9V2bxSk
tzPyfyaVgB3RY9kO8MVrEkkb6+ZAlaEII/uJuZDVKZN+3iRZ5BcQT9lROzFvNb6t
xfUJy1HYLQOmIWpWoJx1EHtNGqm8QiP4CguPOpgOQbH/91TVOzBaTTk9uXIudRcU
R8hhkCdQaoCKnV5w9vSxKyhfpPzmClAnKa9M7n9OxpbBvzd4xLKv4GEGT5qkE3Sb
Loo9sfzWFvvfppmJNCagMD7fobgNQs7gfT5IHFWlVO09Oz3wTgsprHO1SafAcnMv
oYkXw40ddZvC028d54W6GU061mhlr0EHsgfbWBJ8Jc39dW2Vc/UkvPhZIIGJcD0y
tFl6NKAVJ0JU/a6AzkNUelenfuw4lOLkMZznwPVGcRUSuDuERFT/w7mwUs9Bkl3u
bmttv2xc3W/hc3AkYfQFxeSIF27KbX6tlGBpEtLVuF1sDi0vdyntgNJ7Oap4zB+q
ePc/0zChhCo3kv21p1SAKd/kUV0R3XPp4tktHsuFoks/baeCzzdDGXiStZ34FJTe
3VYriAFYZ9RsagRcrBq0XIiE+i0SNB070inpPU7JzkmfGJwvsTZLF/lPHe3CSNmC
TUR4ndnrh9hZcrjF0Tj5sU6W3vE5ddIFZKaNp/nNZ5/3lJJpUKHIMUsH9fgzqOIG
SIMHnfCNOs6AAq3pFBo0Q/WhA3VBS/nHPRlzDWBOxRQ+7AS1ygK6fbv1RO+1u7v8
LFgIqm+8//Q4/ZoV6+6X7aMyEdKje0djj6QBuqmJt0rU7V91dk3tU9OCZaXhJmpV
P9kW7j5b9c4itUZLbvkNPzVVw21acOK5Tvnbct5gAa6W9x+WsH9t8CV7h2iiGqIJ
wMAF9/JP6Lc1qAla/QGKMISMsvLLgj0nz8k73Nk2Bf31ZHq6NgVrDExT3GeTRsbp
gtae8nmmrlzQcehmEisQrl3IN1xzpllnHpguWplWYKLM1awUMHBjwEgFlh5Xp1MA
diuAS/zMBocrHjIj9fmklWOzxKfzFFlrPVjnsVkaaOVmz6OLDiUD714ehdEfTNqg
acB+3gyTWypLB8Z90uegz0Mbbom7182hCssrz36t5MszNoTl1HTiNfRrDlUl2ReW
1/sw9jTP6M4P5Oc6X3+DPNXfvdbCcGYsCQ6nKWAx3RVdtyt20XWQof2zctVwlXy9
picOs+FTTLdfYI2WUa2859AR7T6fKa/rmHvyLfWFXYGujDf8lxahwTkeRz9DGCIh
FQIQM0Le6HksagaqiiMpsUL88+mLc411SealYwfFZ5T9GeDDKg2GHqEq1Yct2WMD
VveFipz7IR1OSdKG7QrkN/r/53vcbjiFg3kFOTI2d0D/99RnIG88UHLNLSgJaypI
2z6xsKZUmHd+vAeAkHbzlOkhCif+hfRfxsBa/EykBXNgtR4yjI+dAafJAFx/B4Bx
dcGv19HptKFTTxJMTRSh1Un93oxItHUz6G5AQCtnG35A6EATQ4IUpTKseksA/VTA
I2P2rgcxtqP7gnNj2RFiyQ7e9fJ/nTgMqt6r5KGGSGeU9iQ1OIHI0Py6m2SSPi2N
YUWLbeNoCyZtwHwXmXHA/0EbVJXMKydzzW+KAh0jdn+ZkIr9C1U8pCQHvtYoEi/p
JQ3FkU24sxJHh95K5tSdE/ZBEbLWeYxcR6paXnlASa0LG7+t/OFnPQU9xsMt7By7
GBHE/SfoyxCvb/1Yvo64ct635ZJN+VlcD3DtMreRzosbeIaYinlX6zHJYDM60gq2
daCMVYQWKO5Bx58s8WEWh+hFJxMR6D88ykO3ru26pQQ4a9MK70jzlOWjp4wyoHWv
y459EaWnVoVamNBJ9WjmY+Ko9W4Lnz79//DAOG5zn87/IIOmg4kAwCz7JTXLHoQP
+DkwXi4BWYtFejGb7lxpJvyJQgryeMwLF8axCIeu3DFo3eo9vx6DP9UsUaQfH0C9
KzLswIvJfDHXjNF7BeY+BmP04bz+JKAPg3cLCHUWR30yO6g3X81IOK9qC9I8BgV6
MpUjihW/Urn0PELjBVN5dWs1ue04izGAzIDI3TPeKtjRWTG/fWije6wpZwwtqtEA
mE98O3pXcadet31AJOBZUZbbQ3kMrBCLHoD6qq5pVV12ucXk/xatbXzJWBrKOr2X
vVTXal9U7fUEf7IwY6BIRIg/l2xrhQCec9aHY82W3XfqT/lt11RyNmm1we6l0PMT
wmx/pedDPUigwtUOAW3FVfQ2+jvAXShua03pJJNScW/kaMcpj69ImZ3vC3JtPhKT
PB1s5yeHY1Vt4TiPmLdob4tfeLoDm+YzrGfdJSfC+VSfhbHbJ7/loA7fyB5FRx7+
4z6Gwj/F1lIEtGDpRV0pYCVY+kLNa0kAc/leYAInMP5VEYBBm4nhzGPFegfLdrhS
Tf+mdcedz6uOaK2gW91el0ImPXS0hrxH7wrR7Gp6XXrFv5Pbxqcw7qUQT7DNjtrL
38j24ewBdmcuvN97oPAVS3Fzbwpedt6MizCtj/1IthSPAxsl0tv+NiNm6ZBR805s
kEVAXZ8+SU/PekIJ923Lo3uFmG2TxkO2kj7pC4VmByjj3QEe5Vbn91wdKCet1428
7Kl0//J7p9+Sd+I4lJ4j56SM/HkT6GsNjSJ+icd5zppiYIx4kwt3lwcIw3sGAILr
MRiY1Fs97qMLz8bdp7K5WkJSCqx9D0Y8M9aWry5F2aJBE0ObViTHgT1uPOxMy8Zh
FWm+BF8VTEblf2WQUlwRO+Rn+wChCnDS1LP7Otr3VL9UtxxNQKqvTcxBaBy3MifH
Yu5Gyo8v7iE/zEQnsdPdXAkSTBmL/O5rQUI8s6hg13lLo3cXT46TNwBg1NSx4ArM
BGvue9i5/1djiryIoC1Uh3labtE9U8l0hAx8UTL5F1/zeK4MRzdwR1GSZwHBg/qE
wMElegflRYyP4eJdxQ6WVMdc+8T9MTjJW80pWy7jInE668e4x5BsOerw5eHpJNYS
J6Jfgm4lhOPIBfA2u8ZTjbX4fIq185HvZRsx1hLBuM/lAwRNyaQOmvEAsaJ0X6OL
efinKVqhBsNMTMaetkJVh83Em7WV8V0XEJUkHG189alR/mOL8wun5meRQWi182LI
ZpJZJU8XwmQbsNeczJQyERZTticbZfJkMHpMOALFa4pTDi2K2fgCP6rZFbrrxRJA
9QQIp80mUHNXguyg9WdiK962LRT2kUDxOWL7pDJ+hanyEPKQH+nMa4UEEcPGu8Tc
LCeHp3uppLYxI4zBr1xpt8jtTG4vnrxKnO5FiiheIdZ0p4e6lN+GytbU2ynmKoAj
YgqSW92xRMfgZmZKK4xWGfutN+MhMT6//7WKRKq2I5mTI2HC9ucUTaw9qKKG45nD
JlRARN6FbaNDbSpbETqxA3mxLIVr6g9pTuz07Fv6T7CIn+QlXrJK+2g2axEoiV3M
b/CyENPk56NofGIBAEU3Ib/xhYYcm6NLYL55y8ayXoskyzGka4b+YtB4pHVRwnUb
9pdec/Zn0MXGMPb3+6A2U4hs2CXShwX3uonDRfM7DoYZb2ikesrJAJvvB+0uS6f6
T26gu0A5Z/JShtu+GnZeq43mi1R9TanO4pHG2uaXTSqPN9jV/uZRupam3nowa56m
up/zHe5HwRIwHjhBFWh48EzO2iVNsteP40XiZBrhyR4DICnHIH0w2S2rF82ErE82
5ywb62GN3WQQUKerhS5Gg6ageNL2EPKy7rK7KaAmAeZ8sp3NPx0TurE6x0mp1h1s
DvhyqrcbYewgJQzzl2mSTg1LhxZU7Bh6/lsABSmZnMq2PSYhpGU2fyoeEiBaBIYy
VFfhbqE56hz+RSKlqpKG7zfKp191kWjl9hjsGGnDp4Ey2GgwzqK+4VlaCa7Y/aYX
WU+211Bo6Kv87CXn7bC3TsXHiPk3Q+fjknL5lNRur6stcLMVMNDjoNR/F1ihSpb5
z+oLhI4kd4YM9I89X01uNjv7gOeBQqm4hTnNX/BuCI8750KHJdYXHD4Qg8ybk4EV
pA4LUIFfa+en96TsxrNIMw1kOvi6P2SEmAuJpo45+mbIqJudEmlVh5F5+v7Q9Hcw
pywvqKEktwucdCFj0ez3bwbqs4GBYAoTgrdlCQsCkXb0Tv3vPnruKL2I0JxorQTH
xOrYO4Fdggrcn7ucOI3xNd1oIDwmunr9zEgV22/ORWPq2QNhLTV2MPUacds32Lg4
YhqAhV24o1E+BlzufSKHwg9APqIRCZtbHFpCDog/A4T+aOBkFdEme0Cp8KhRT1sF
9ER7b5m9TpXTTY9P6o9+M4OYeH4anARVSGKWZS9lq0FShdF6euUEn9hsWwt2aVHw
ecOIN6f8/QxWD3nljkg8i9YjO3/1SP2BfAZHs7RYNhWHoNU+F6ATvqVOd67cnFyX
QkT+cIsDbMmNZ/M0mafu0QXM9YUhZnNwknQYzMs1gJHkwLxjica3zJT9i8dc2mV2
ee3aP2eJvXmB8YTIGcaa+LwBT98RA57nKImLO3AkcKdKqOG7/zH+SOBC2gSp2wgf
gp0ogecdIrfjqYwExAtBCEN8f9s7lU+fwmhU9KWS31l12SXD9G6XROX8qLQV84w/
gpDcG0v9jO7Xrzm9Gw85kEpF087l5VdIcn4vQfQFbQfpfSXsxxuGHxLiMkKQo8Cb
kFPRN/Vv1wn574MKX79d7fkIhHEF7tLL95dZx91msXySTfJHCKV95BahYVvPljN/
vVziK2N4zZRbo2KI0IMQLx1wFGyn2gy5ksnab456ZYSo8ELQSggVu34frrFu0Plk
jYy345OjvwvtNYnS6yWzq4J5rXZekF4qwxRr+iUIpuq7ZvvTjq/yTRuQl/l37g+u
/zMthunOHGbO36/Fcoi2w4+aLCr0otfkxhP/n6TwJwMr1S4TJ51syGLCb2YcqX9D
7d3Fkg/7mXzZM0NeKu3ukw/WWr93MJCV90ssKzqCgNUz012iT+3bBIY6LTQhBu5M
manAvyolEOsIsLHayZ/V2xXsieYiUDgqggv3UZbLu01nZFGZhGCezO9AvrPK544u
X/VZlAFyM+JZNy1mdhDoRPYVk/7hEpkbMRiNr99bpC9Vxu4qOrbNJNcVhQwyJsqd
Z19ymfBMUgX8jsSIBfhuBx7FgDUNsh3SrPIPWuNFsIALaknpdBA9Q9VLK7mxZeuH
rkXoNBgpdQln1z2v15YhS6voYuCfp8y2gBP/tuBk8HrQzjrWrpkgm21FzxfNgtZI
4wBRxY8nd+F6nCMnFR1UPGwkSwmmN6As3+RTbNMdFsfrXlt3zjnUPzZQtJ9TQwmI
lspau6SQFBLeFM95Ai2m0RbKoQST2iZz5VKvoEEdMnJmlwRY5zJwKFQPrXmRguQt
eEsgyR1jC4YliMJnZpacHxvUOTzZUjOaTb/j6/HxKBn8HC8njjvNRCF21EEHExER
yx6ZLw554/UGmcq8SmY3MqoAJexn0grYDbG+QvqDfZa44sl/HMYC5jvQJT2TQ3Zw
svuhE9AZ2n+x3ZOb21PJdzCCJN1JtuGWUHFHdTwOhCwk7NL0HC+NNMbsUIxzQh5P
sVo2tfzwj7uNdO/sIRgYvbcGQu+nDfx45c6aemYNt6lFCkGW2IG0DWeLqWXQmphx
l2ux0WQuslxvLmQPZMxsZ8LgESoXmpXoaFo3fhJ8nfhEACHFW3KYB6kafolLj9ER
vtoaEY+0jsXLKd6bgtokPw45eetwccms3dFtXDfgGTqAvHHKZKyxFOvIzDQQkdvV
vSaRLNav5150Y4mM7HR1/9+7u+LRzkAYUImAmJ/rWfUmoGZPPOW7FloqytSlU6bz
h+EpgqsvIAAZ3w/zmsHaDBcelSqwGR+a7jdQ0ia2IEnsK9p8UvC7f3g52BOfEzv/
ajePkqf1rgypxTEcHW9lEhsHoIeXi0xEbAeXdzbeFdoV4YWdpMLKrLKh71lS/YPq
Ybr4BsD+Bv7aQiHJURM7l/DdiEEjO7feSoQ8lJP97pbp2NcPFSCYfTyO9PAWr2Y4
JDmwyx0Hs2tOCl+EXGTO653FbckchJ8mI1iD8wBebzupaQfDJEr9yNNrXQMKRN+C
9Qs5+FlfgpAg43EkBFk8MEZfmPi4DQmMEr9okW5kmtvVx351PuzCa+y2WvSR/2bD
YpkBol/zUBzDsGiVhpkYV/KRmviChujWuH93irxffANZvcOGgkM5RSS+OL857eum
1DEZxIr7CQgiYiU1juOY2ztlBO14ZFuvNhbZ9vxk3WYPv/Mxovaan6fP3cUqyHO/
Wq1MGzk/jp3tkQzkDMru4ztKYqcHaritmtvsc0EXXao3QhfWcDRJMuQa6Z1nIaZP
3aM+ay7gEKTfsIoLQY2JqK7M9G1YIMgabr897y1RXyiFOZrEt1s0D8H3s4Uk+olm
NX9FaFsNxo4NJkXwF37L1atMPJWBPUiUeDzvR5SM8Gf9FIMiE1n24RfeEReihWd9
oumzjhaTItib6/pUE15zhf0lk7gucA/PeAZm/OwJh0mAiHkzpxPGXpT3mmkX0mwI
dIeo2nbDD3/C0grcYPJUJSDyfeUslQ5oMlNFH8HFGRDbb7inBYfuiRwmXKPt7IqX
ZClrUS+c01r9nMD+hVyGb9Y5qMNVrdTCEkTRE/EkwHpj81jehbzPUTvpzpV+npXM
IMk7lu7/e/SoqmQBNRc1SU+pgYdOuD9uNhgRpn5vYrrtRNZ1QQgjioO4Sa8AbCjc
iPjtU8rCvyWJV4jakelWKqlCSaRyeCzuJvZaNqN2tSlW5/8Z5FATIPXUBcUBoYAJ
meE283y24d0gHmWn2MWi9scc3ToQuFCfE5Q0LJ+Ln2LXGLAMpte1bcrLri0qWq42
6iTDD6i48zxEH4LN8Cskna2jembGw0AyTdajHoIXEF/evT8zxqNtSZYiyvCVI4UO
PRqcYUaFLVkoRc20cJM/70rlK1eOuxq6poxaFPNdu74kQFwtQlco1plhadd0/I1f
T7rmDkDDwRAtdnXyc3uiW/mpJBcQI2+n4efpC+tKDVnqLou+feFCodnaHFGyiSYt
SLxj4kiw2xRsDQ3NNjnhCaakkn8pqim5MMOKiVhGuBsMHiaWTfZVUCPz2LlFrSk1
UoiAcyefmZ7frqyCiDLE5NZA3w7Uv34mhPSydF7LBGGK1nNxW8a6ChjURUWvlG0S
qqLkPlt/bAymSxXJyWfEWkGUNnioioFoD0/djx4xC7YuEiAiokwaGAv/mR1Unqbp
BQemk1hMOapF2Pgy5Vj/VqqLGGkYr9iJ4yia+VbJdxssJgR/C670kK+n8HLMW2r1
HbOWWiWCW/dsptJId+IKfX+WUtp0PxHV02FhG+5o5cIidTRVoU+Myot40cIna/OD
AvKPY2LKkSCN4Izss+tKvp9S8SoLhLHNIf7OGPHFAJYdcxs87Svv2mIYrXiBOVOQ
XFiE92R4KdyiX4r/FqaaHJxNa5gHFDZ0mWJIz5kK+Uy/wpeclPBtua4i0lyOP/VE
RJlniO0CUpTE3FVPr6S2jPpkZwWoay8by434FGB7IFuBgnLkrLnVG3qmgzKfUXU3
xH+1WyvEFSlY2TAM+Naf3NQ3WUth00TwPP/Qy9K2O5NuQ+E9aitHZIQcpTARz/N5
rZavqyQsNkHl2LQDuT83PULjiKHVBRXUeQxrBYZUI8DiN2B0p0CfW+yj+7bB78sP
ambTKBFv1DatwZfJ6s+zAm7ojCt3hpiBXGbkPpioCefSoEwlLdL1WybwOKaHLFUc
fU9KWPxIcU7MuA6czDrZn3Mgx9NCNhIiuK+cAhEtS7I3nsI8Ni2ucHfgjQ5KTkAg
p5j7LQ5IN3rSaaIuBLfC5vsLrS1f8KmsKTiOwYXgYdBOJW3JAlAa+Tox1VhQjLkX
GEgc8mvhMSSSrSxPguX9fO9+9XTnfTge9861pi1/a2u/y6XoFPYJPyKRACXszAJQ
09S32Gwr7z7t1fyOTDFvscGXDlRVLU7Y9UDq9qB3Fc6mKwFec2FCoB8tBypyiwo4
lGnHZM+XTEwgZFSf1R68h11MEI10oT/dcpPcrAvirF9WayLkZY2k8xeOqGUOAh+j
ZdPetyICSKdNSa2BjOto/1BlPLNZvJ8A3vb7y3q+WN2ZFmpecycsUrZnlrYUPNRc
76LQaFsrH/idlvvktu3TpKLlGLoUp41VPc6AWbW0vRqADcu9SB03NuUOkZdJ9bNd
tzdDLvD/uHRN5gKhzX2K8bi86L+BUrju2sAJsIeMNISsdGBMY2OGlfWXyfter9A+
D3CzvdtpUJy0M0Ze/fseBhp/BW9hkKUMWMNeHZLIvC/XsQCuPHNWVMJVcMhI//cQ
+gzDWVl+k9Tmajv8ZERvx+NbBYk6bFZuJrWoXyWQpv5I1ur2wINY7xvWTg9Q5J+T
OE7qLf8ucDBB0qCXkCNZmKcGlf0NFFt39Mp3XfmMkYDaYQ8GRKPye2L1ZHzzD6kI
4oXPofAtCKYuqGQDTSh81pDOTSzed4kg0vx+NW2jhl+V3iZ8YeuLHDF6s6mzE0zg
8qydoTvxBc6zAubZPcBFYM9FBO3E8d8oTp2j05Ugcmed2TZnBjVcZoEqazNkrSfw
bcyzHe+Z31ADMgnWtvIouYeBFv1WC3opHNSXlQnKLZjFxTQSmdMjpGapz1Ibmc8u
SXdjzIZrhiFY0XWXUlucVsU0led9usFcC+5PYcH0yK0izWNenwyA4u4Rzo0Iu8Q0
lQq9AR/SWLmyOrbYCgpsObn4B9cAZqnuwBVAhTIBSvUEL/fdOZXwjvrZf5+kn7dx
8MdwgtFD2rmQbs1KyzTnqJIQiqfUlCoJF/r4mA408vxKjP73dB4jb3u8DEA5FPoV
pkl6b/1JliKZ0cdT6FP9dpRiqdQPNpx3/41Q/oJdJ64QUHUZo2QIYQk6bnVGXkjb
Ocp2mysPslkPwbuufOY9kK5qBmqm+hwYE1046hn9KZHG+AHiA3AqcXghZzHnpLsF
GzvhdU1l+Ju3RjOKKDXWOf+0G44hikMbsYc7TqO0a/pltYm2GThwHLiMBw4IaLcH
orVLVIMYsU6V2L1e92oex0I7gguiSDQKFGxAdhUy2OBTOmT04FfPpo5y6xamtiVu
w4mPmuAFD2acIIPCnprNexk5UmNGb3nt3mHef9oYCRDOIDNNPGUe/SmU5v/QEzPs
f/tqivBgWK3D2ARpo4/IfOotYVDmRDCY1WFvCWCsayRSL+u/pkJBxT+J5I1mdRoY
90hA1F8GO1RW/eQgNy42+hSfZgRi8xXPm0rDHGPuop/DJAEcwgIUSkZ8KkjWbgdf
UuEVx4vlUQ9nqYOOEQzIrLw0erJmFuMmw8SOAqPCo7gmV/Z80sKexvu83FGzPKK8
oglD5whFS2FM7aiXWL0HgthtH8yQvNqdVCyumHUyc2aducLXR4Z1VMDuLAJGTMOG
rDOXUfXnJoZ4yDHy9Vacm4AYmgeqbgsnmc01HGyEW5jcLmdEnJilXAB5riEtsA7f
9k8NAuZ6Vg+lwqkW7bRTcnasZ/Rn7T7uOnrzsqvAIWTrY8Kx74g47AESssZpvliw
G1ysuNq3tuSakk1iRZ+dqaA9JZBJv4Urm2PYsHPsdTDoV8Ho7oFXwjWu2C+HEewJ
KGp95zG+pphs0CJ7qo6uZCtDSRuzU0Ir7yA/6aNFhtvz2OxSIQwEeOdTkK6ZJeqh
Z2ZOAERuCIDHdaDdhMZIdhjwkPjkbb2BRRgKytffsCNyRbgxLWlPmOmerP/RNuQX
iizRy/EIfrOmWCysspqWHn5rEPLJ1zkc+BPfuBT4RGveT4m/vf7dZyDM1CJiqUM9
TIgnFPrVtnnBce3vnxUESPVxqSKrDecEAoArYhlU/6s9P48TWOPgcR6XLhUMB156
aspfphQzI0seuBNe5hzFDHN4i5iQihddZZPL4RiK0oQ8k1PjeMTS9LTMwlL232LB
X6Nqui22GL37tO+oj46slJwjZmOFmXym02lTN7i2+3jJ74gWihTGB+iWmIuSgh2A
daX2NIaA+Bt1K094oUy83KYNJqOq/GokV/kBhBgEirQOoWotKJCW817IR7yw2CgL
j7SBEWUsBQ+69q6WvmXb0dRWd3UlkEsaty9Hs+OqmlIlDd8y2c2XGnt/KR1yvfJu
rmQXuJ9yKo1sWWESnWj+knW59L4JKhUfcWv6692oeAei3Yz3GvjU83FaaM90aSSo
LshigLVuKDuvmGbAthZsWl98dfWudZmkg4s5ysoqQUm92UZtG7CUk5Im+82N5lJs
w8mkzOM3WYl/306d1sdAsW1RiYWtx6HletdzYDqz3Y693T/W3rCHcvTLZIqpaf8Y
pvnE/beSg2YsZYzMREjh1ItS6rdImt19/210TQJAcTiv/UizWlhuHR69K7d82Ixj
IkNf7J38vrGx0V3Q+x79YXrIMi9vMEsxkmfzXgwf5dyZu9bduBqSl5qtbrNy2KqO
HrQWpDgZU+MdbUSvDuaXVEu5yvB486sp00RGTua6sKa/gfzTwu0glUX+Oz32Zsq4
+QAsKB/mi9crUj9aeJ3eZ07f4dNJ49e96MYhYT87IJ7pv+vSta6XtiNo094fcpAN
b5d8IDLBsDC6ZgNZvy2s8kuJFYun2DnzuvRCNU9a3bFJV9d4sbQSiR/tRi6Q1NcH
bdFFfp99X2fCmTxToGod2Mhvw1gJdlMz2SZot2q6oF8mGkdva2ZqzXj/nBNZZjMC
Qvx0OP8L+kifil5IlkMkVATXWBZPAZbmBIYC7kyx67LEoNpEcnpbOi1EZ0TRGl+p
sjO/YlRAWx1pkpW152ZO6fp6JU1qWf0IcF1zRRcd+AGhVAVVEtkn3v1VFBl/bZRb
z4JpBnG7E/weRSEJk+sPWvmMcRlyNjnjF7SiK4cCuP/oVloY/WVNNoAVi4x568ei
pcIQr8w0vOgw/1n3Qqub/nNQvARQP6aDkFyPR2Pl9CURQm9n80wwMiWZ9zUyoC0v
/InFNC7nCefjuuTUJY8jip5WeKfC041BZYvcWwUaNopftiQ8FFRuf9hO9/TU4ydk
l568NywLN6fgdmEBIxx7t93B3y0sMjkhPN8lhIHZHq4iuZTKlNwHAAWgE/3ZZozb
f6KIQVx+c5oW5mSJSo77pz+T34wa0hzVt0V4RQl1aE2K/v/Sj6UHA855oDPjIDqW
v1jbeP6QcuseYUq67wmNUnBwVDklYUkBmFOYJp1Oly7Cgtr0o58shkVe4kGj2kZO
DmZ/HEkJS1OIXZ87V5LidNBjfDZ+A/jhl5H+i8bRiuIseeJhCxGai2fgi79971y2
mxkY/BF9WUahAW4dtMBVbyxEGBrnuCVwMm8CWm8pYNoz+zkde3a5u8o0TqJyu+SQ
ScbW1U5KR1hJga+ioESgHbYfYPwMwxxw4mg2EKOngUmuwYSZlpm/TxxdoluptzJ4
YZn2fv5LnuZkZvuQ4lh7gDzY1sF8tjcs94I3XfD1P/GTUwFd91fqNR1uJlcWZ0l+
DSGlaVZOnLHr1GMwRb7cXzF1M41JuFSdr0BYXhcsG4EnriSZB01Il3lTGk1mZxDu
uVKQjGYBGTuKFbC4OjGfOYIGl9AMP2y446Sbu05NAYpzs0kxRlz+1Yx+hgh1s/KV
poiPfxbztJoRrDAI409f+5H1NCSTbyFZWaVGITGRmp3NTb1x1apf8OvR8IewjAVf
PE1hBbB2mveBPtDFJDoRopM6zt5R+TFYWpCgOYF6Chu74kleCe/+SAD+jbrXlKcA
8IvXetwDFGdF4CFC+rlKEaDQWlm+QrgmHrUqgmfF7K6i/ylCTNqovgbtwLU9wQY7
v7dMOD/yFLMv5WFGuIVHOnNQWJb/QgL5mYGgcH1LrswYrMONirJtqvGhmiXVo1E0
raZ3F5/IeGNCQ3QqMsqmGKo8QejwqfeQi2jYdq6S2kQYjKqhBZ6aqHnmTD7zTYtl
d60d1gu/+xn3rDt562EGqo0WRuKbrbJBQUaQcDbDGY5+cYKX3oXBtHWVOJKAp8wf
frUV5FJinnB1JQqwu/kt0u9SEPWydTFJFv9NdSj1lOfczRK1Rm0y2eA6+zY7guuV
55ENU03+i9e++zDklNVUfP+nLGty1/2kwD7rbdqmQgYyc6dfwGZtSC1oMQF5yCn4
TGqRtcbg7N8vM7iP+EVfxa/glcDNisOVf4tUi+MEPINZTn/4QdipfH/UkZEfo3ui
RgjMgsbmHu1fd96dwSIUReyniVI2WE0E16xuVxgr+Co48wbM3asUcqyuz8brgsVv
2FkauoFb1g3+zl8zn1SgBz4YaqXetBdZUEQC/m5+orfl44acARUU+VIM+7K+fMrq
T4a2u/Lk/Ga21K2LqSRFpDtJVMC7lUGopFnBI9Fmlu3SlyIuK1fBfiT6oaUshKsY
ibEocQBRpla39hAtFsUyUOK0CwJBRLpl1/LTf953Otn1WTLbEIKnpHyc4gSJl3ja
w09k7N/IxD0nkFqN3+491oNGB3FFvdjWlhQZ3+CD6SGoilqH4JUh6uMITowIJDvr
pXtwr94+yAyWtQNK0UN3d47x7x5DleB1/8lzWo0kjvGLNfYQqSe8RfaLj5COHDCQ
WNFS7M/R8ACec2QIIchoCpzqHN6qmay+/ppCiKRPo8bB8+MvZCrWSD32omqeC9Ew
QRIRdbtQ6Iox6IvlELJ8K/Tl9dQnvuyN4cxrehScCoirYD8+5cZjuiQzpBIGKrJg
4CGD+XiUe5a6lNrhnxQJNrPrU/6MkIgqx7RBBL/d/G/fS0ghDaiRGm9RZJEISM4v
AtV7sCBsRkAMoeFB4YOCZooadQCnLAoh5dyc/uBP39HW9Y4nrTBLg6DeDusLdH8x
bdUf+EPg/5b7TpPHquxhDz2aSHUDDk8zWlR9oeN2QbGyoyV9yelnM+7f2LqzvW65
+rTInTZW4+azRowq9PjWlCEPNQAqPkq3oSQIj5g+l2urpEGeLYeuQB7QQwgHhUYy
+J6tbOgp3OeS/JUP0QsgR+1Dn9BOfRxTbMnBO9Ah0NPqowG1y4OWC4acw8gINKn9
xTCDt9ik0jQe3E473D8bYaQ48xd8DRVpoHAbUiYTYW1MqG5UZuWt1/TaI3ThZPYq
NUkjNNrQEQ2wE0+dRMZHPUjBmWL2g55pHneX9z8RV9pxzqSAYDQ5u6Uo6J4V+oAt
/6Tw7M9SlQ6haDTdygGAXGB8jinJQ5Mv7R8zl+ZLK/CgK+XrhrS64vqpDE0hy9hQ
Nas50Rwu4bpX+Rotkox1aUnPvGwBKEs35vv45VI+ij2x2BajaXL6HQwJh71sP/TD
yjyLDQ7cTdmEkDBuc98Y/rFChl97oP87G+SqYhLFa5r/zDxVg7/xJCUTdGa2lBFf
+WlaayV4x0m8UWnSDy2bY0G7vrahuyVpy7pjQ4/XyRQ7+2Ig7l96yHoVA3K2LUJn
2FxFZGj5F6d3fQUro1iH2+cMEYIZ6FxhxR94fIEuytklZC5NKULi/PPFx8mYHdUV
pN6yJgaM4u4CDAKLaevA317hMsWL24PW01VX4sx6J8TM3EMKDX0O97aExv4WAyoM
h8Hh0Tpf3T46GEJn/OWTJWADf86vPbkGETG500NLQBcDl+6Kons29N2V1mV5N0np
Jl62ti7kkzk0+6LGQzbb0nANIbjp/ZNURUqBqk/OvzAL70AhFHYz/p1KSEnt90Om
v5DJHsaMqD0JVJj3pKTG7x1pCKfcJGcuDMf+ETcXIDrdP0Z1uWwhPXobz5y24XIe
rrOoaFyoROg5t+Kr2ynEBjjeH9JqmfHJ2iz4clBGdb7Pan5IgZdeS6mb4Obhcygd
4hFRxHMTxtYKhuK9zsjgL6Z6ednBbKxFpVO6HLwJzCPhXO4UQagOd6QPVCIOnMGb
8zoOGU0+Q8U9zHHk7T/QFPf3oToaEzKU94JiLPO6+JJSl4c7Kkxk+LknPA5zLWwl
HOvJh8+JDjyp7GKKwVmtBC+i81XRvL5sKIKL67RJLOw+OZ00zETH6lnoRe0qgnbS
TJ3HcO5SQ6DV+Reowwcn8byMUnreOM6fS+6eGhLjMIQrlQ9C+jYXJ4RFCzUuZGUm
vjC5b9hlk1Ru33MQYpQkDz/9QhI8xYVxR4AvSgz9Uv9yGKOtQke2Wtbwoxx/czS+
NBVgUf29MhRAVLB0EBd7g+uWw4DE02rRV/3oBijsqcj/CiVMqVzElhb4LacE+CIa
JDYPwqEwqDUwovTOkZ3gC+H3YAYOZg2P1Ml1LoXVqAiNvO6iErRZvMwZrnD2s5kw
o9il8w8kjoAiv52ePl4Uf7uC0sezMQ4nsYF0Uzsm0ZxDrYAbSQTQxyT41ONEqWIL
tNKRaz71f3QflurBECwvNAfJzYFPVxYTZ3CBTV1w10/QmTXPognRX0t6KLT/BkxL
oh331PW9lcKL8r4kNpYZlHxa1RsCe+hWF9wZJqHYxxjKtl0eWiFE9q3U5Ze/JNMK
l19StpQs1LR5bPVxplIKXnVSXseR/iR2FwTC1xSqpupPtEbSFqqBtSy6KS5yC1wA
1SJ/PUfpyC2SMgg4tGf++6xwrYamaNnHwR5NRVo7Sb/bMWE/XLCfvCJLcSrgjsdW
Qk0hhVRTZF6E+9LMEAWNHvkeLSBCfNUBeuA8rozrIBBkHVuSPbmLEbKw2h6iA+VM
2wG5WxJhbcyTWuvIiyouhAM6fYYXYPvrCsa4GmLp4jd1pVmEsTLSoKXxUfehCu9J
ymSuJlQ3B4qW0WIPOM/a6isV8cKfzheVrZ7wWQuXg2C3Bx4V4A/0RiDFD+qwhYpa
xxbKj9Pk4E0KpmHKvhRMjyo3ayfU/diAZoctH3Rl3jzg80K6zsFW2HFxaNtfR9kY
4UXjJfe9yhb3ki/fzPllEn+ZLNCEZ9uqqXwD+0JfuKZA5wtMRoSWEJZWa4hBSjrB
6sEp2GkRJ3E/S7USPohvhofzV3ptMYx5KffbgoypNM/16i8LKi0UmdGaH17EmGYQ
2f8hUjdPj3uYry1j0QuQvQXr1ijuqlcN0ccrdiZnQVTPsAuByMV85Q6HlsZAg9ch
ov2HdkHRZ4pvHO3Q6mOXIvL7BituH0IwuSgvKWaCT2RQaJF6w/QiGV/Bc4tF9bgq
749WI9QnsmFyD1p7QKtW3itNpBb29qFYbP2mwZsVyrYkuUG4lGu1c0CcdjlIKhPl
WWxB0XUonLIaLQ183TyJu6poKygc0WHTMX/KdBa2/5r6vSmWn0o7BYa9Mtkpcp6g
Orb4t9h1fIkAOxu9HU0rZPxDLTIw4iSGXuHmHcWxBuE+2/zeo39iSiovpKcvbKwy
sJ9OVLgFmwW+Dd5FoW6c9BahbksWxs/OZoRy7ziUhrIxIKyeHTK3YkTFuaqj4/0i
BQimI58EB9RfJZOf4dbXbrtR2wus7wVNE33kbod589qGLlD7dDGWjgZTUZzqfO0g
Q+G8r6uv6BkZ8WN2sBlzpl6Kgh0ClEoaMGN5H25WQNml+CR9SkkBEykIAS2BeZPi
YIC3/15P72I/DJCJi/sx0+KJIBPfToQZjFQm+9G1y8ljRauoruUfPOLTl6d+RVPx
JbY9VMr39h59Gn8adm1bwUiJ3IDfWLjUtYOcqg5EcwJ9C2tZ+WUiEcWG3RRZ+LFA
y84MHFxk6dRTgmiz2aDpApxgiFfspDSWB3F0xCVqu1LUstk7v9KpZrvOYNaND+yd
mcjIkmdD/pO5At108UKB/nRKlrlKhws7D+/k9xjNm0ig4DPvnyEO4M3QMhLXdEsY
2M416uXGWni1FVVZp5z1gwrZttgMJuGSKyMk3XIZKXzbIWRbVpG2cFKWRH2AaSxf
4QnrWvytlmDHsOap8Vxl/KHjDpZqJ48bGKyzAH6SO3MFWMphinW1/bYzhAj6gj8M
eg90aAKRNyxAguc/voIoAzjQz9bCtHOG474EzBatYJGQXkMX28Q3eg9EozfZzqLM
Sl9DJaPjOxEHJQ+OwqaEeVS09Cln6t6sa43XxlghiWyH4q/Tch9S2ELv+COVerq3
WnBddk5eu64F6n/EKE9+ZRKOikr/RFFpuopvK6eLSpBsD3IU9Yy4GkDaGK/zVScu
QVVuT7A31C8q9GAMnzYNh+NlEeE0BBmcnVDk8dqZP2OgLgNrsPa2Fo4Ia434expr
YpDnGCy//VrhP4SnZmhkFTLQBLdVBJGFrsJsAbMfs+VT6MFFsBlBp7+HYy7LF+PY
7B8aPP9/NQ2MIzM5dshXuQKsXKaBv0fgIEUa/nxrFwWkNMh9+N2MQ7/1+R/4+JAO
+cJF74elEyaqVFftWbNzXXlM3laoDfA+pPEkPnzhESi4p77C09+CXxyeGeI54nZE
N6SdIfooc9nEEqSwfbqTATkU3UiTRaNKRvz1qkNtq1XzDovM98GBvaJi2sBr2pDN
uKQcV/bsI+YSAA6T6D3ARntDVKroYt2kD+sAGiIjsxfFz8+7OTuQE0eqwm+/hKAl
O1KrEjlAbodPxy1/Bjfi4e+rxwkT3fE7NmMQdUyKohhtL+9lKq0YNiQmkW0aj0bx
cjJiTCBbpkA9I9OHNnsstXJeNmvqRF38H8S2qYKUIxg1zwEnXdnSG1mxye/BVv3s
Kf99UASEPDERD/kx7y6bwxR9FSLzuuJBgj3HIB9RZiF6Sd1eubl1gWnFRVFK9ZwU
rZzayFlQeU/Lu2fC8J8KTEZnl/g/Ey4jIy41ZUWavTUTIRR9BW5BJIfl63hIi2+N
V4JEEppa03PPJbkg83ihGYzcGVltfhIuIV0TpiqSZ3r2Sr6UefoCM8rjeRzMisIr
bhFDOfdNLyQPQdPfjyfLKxxll4gCj61PxPqziVZH2bvjOhIa/E3XSxXqP68LDJdq
UvGV9U0eFv2pkRDoMMD7NUQQGg7sXVMf6kA5WUvs5NMUV9ynUo1bT3dbdoZENdr8
PyfYypawtTsQ5TX22Rj5FSxfj9hWkZsxDnlZvlgAzOJygSKHs9QdUlKhinAcxVaH
dmUUvrMV9A7lPhV534LcyrVpG7wJ/IwlYCEOI+gA0I1QBeQOwflBRM5a+w3FyNfD
KLmgBEqA+iqlnY6A+PxkbbUsQAEdiT/fE2XVsu1NIlVkE0j3rv7gGdEymK70FBcI
g0wa2PZ/6KCBUWKXf1eR+55//A+UEyn7IbrQZi106pklRHnd0QAlWhJt+RMDF1IJ
TFji6wmeqt/29D7nT/biMAIi1MGZaPa5XwaVt/iyIc0TRGGJxuX07kvAne0Jzrwk
YX72lByTQB/JuSq1urJvwFNysrxXnFzJYyV1HAnGpx8URRE0sD1BO24py7+MVEI0
gCOOYLzlHYqagA1/dVj8iKLufIA2eCpr6EbZnf1S12KXu5b1DanfyfQn986vWrIs
FubRTqcHL2dwXGdTZGnL/Xm6etqPRFok01Jau9lUS9DTmt4jqepUAt5zaszmkkM7
cjfRp7If1i4VgKAJOcTR+YSfr/z7iYvxWQrVge4wZDjEqUMjEqiSWlvibF6AiPro
hRSoVnkPFZg6IIB6x5nsoCrkvQ0IEz1TckoRfhOPWLyRdjvDju6TCaNVYAdt2LCj
KI94KMb1/Y2uFUXVhUVbk/xatfoJewDpVuh7S994r9HhnpPUY/VMGw2YDc5ypRmI
D/SvE/XtIfpJt0lH7bSMVzu49eAbO8JsV2WC/oP5QkNDY2L16IPC4mvTClWY4UPC
5LdkzS+05/sZfvgPhwm9pLi7gYNtCd/mdm+AOGvDJH6/tDDjo62TxCzgeFs+cphe
HPwxeBXAABKmfWgdfGygweOZfyWh/KAX8qfvErDE7YGvrN0bvhakU6u9Zv8V1oIz
1vvaoHskaI745hnY+y9AGW2BwbEs24sbfzLs8jm3F0vYiw08Z7VCBzMMnZaas003
E2LOFioSc9z/4C7cJyBoCUaHeMdhlWMiOooREfWggYe8MqepF1kL7pqKJXmWkpTh
TT4D6M6qWfpzH4RFFWfltdzTXgthpPNWtqmpv0H0xuWg9hmjdn9o6UO8iV70tO4B
XruU9Sq+IR7cbriU0MzTGuO+gzUoG67sStZmbvq6RadupUkRA1HUCcvE4ynq86FZ
bU3OJl5Dw6jJGHpg7L1JE310LWwnHzQC7byQJG9r8+FZq1WOwTxFKLdp6Q5km3j8
tyLqqEWeNhojP+40tCgoq14WzVF8sTlqwn4uUH5dRyQFqydbIVEaFeHS5xJqhqcu
cyVcLBjuveC964EBpGIG6JYLAfI3ry6GZbIB0/yWqtDN+jmKotLqrSNMCjSdR7cX
j3EEm56wnJ8J1LujmLOc7IWwQaT/Hd00MwoyJVci0tnKUHXuZuoqxFJBPOqEdFys
nu/fLLCNrNo9LxQAgzQTJZfmdWiUZ3gvtajocYBocm5/RJ1hXMZvPiXYBfmpaz21
GFT05/G5KIyH5unsmgWxIzyaLgNHsSfsicIx3e1ahv7nBjaNWvFpCEms49c/I0KX
BwQ3tIczZtdE/mu0r9xriSIIbIxkxZ+uHYCAiT1dtYxIy7KjJ8sencttjHMq1EOj
jDXyCuXMfKrwFlqJdDMJ/jTsHtCXWlgIJcv84/OLZQDyBOlIRSvzB65hEVsv0LBH
tCXK8QUnOf6AnIKc2LRjXZdJjq79UPLaz1z8vF+eW9nphGCWfgwaZ/uqZD/h4i7z
nsGD7f+3ZzkwvQMq0Ih4lRo7Zph7ZHKyFGrxfkbcbTqsy84tuIIKzSCycD2D1P6B
JU8j/VMmOcpCqcH8XzHeBOvk8H3lgs1FyNpNJnOOMR+6vTRr6ak9qxlfEeWtvYwE
itjp0wvkYkFXKlE+COOB7j0WyPGpz3jPlruWWw6l8PdOBkrXHgGI5pOlaLSrk+0W
cNrr9eHsj+Ve0dOvhL6PRBCFzmfBwKXO42Olco7ZU4Pvw+xiTfnQtS9jZ0mn/3O3
QNAZzHrtjNzJoBxve2cSIhN09YoK8Q5NpH4AuCFa+9SrqCMBPzPSM45jo40JHSje
39VhT7hwGn//f/TugXV55fKtHaQ/Ud6CjcRSVj4GD129FzZf9+ngrkyjNcA3+sNv
LxPayA/GdOIrWzDG17nKVjzjraGOfti8nT9OMSUCipmuQDCiV6eFpWZAPxsdr87S
/8zwsGcsrl/Fl6L1lR9FDFVOTpkzvv3pnmHbUIThFo8pg8hGdCmXIvXKWGGgTZ3L
VuTyboRoLhG5B+fbM2Z+shNNdlzA/W/88JZzEn5mvibzjabwU5I4DKOexjiApVIz
v8VWpp4K6Jpx61j3WLj9SAFDn65NF93o4bbcnatzjokoVe5O96g0XVD+JpclfYax
QX1XLlqVr2b+DuRnu0e3JwNhb4A+QqnKXum5Yjtj4Gy8Hx/TV+pOha2kYrL9QM3k
zfrIOKDIS3/dg1lnYMXkVbnoW63v/SULLNTHrvirZkAUCfxJGGkLGJgPzCzLAbma
e+mYGGenf2txG+tJbD/3/96nn3FrndPY7EdMxe8cNPZBDnAGBlpmpGpOvAK5JRjk
kRBpYpuXL9Ql6NssTJFKY94Xy8hC0AIMLDR2fg1R0Tbuw6fjL2fIZB0F/ZBseYjR
eW/g+J+qi2XEOHyTuD4dMEyHZFA7cT7nPrjJ+SNs0tzTMnHcik+LlX0gn1X/aKwr
03X7bI1hhTT7oKiUVKvxpeN7CkcEdLwP6KgOl0Cwnp/n9/C5KNQ5uoQ8NxnKpro/
J0bYJdLBb/aT3UkfW8CxvvgWAQMMShym4hFXGgdAFnhgA7oXLi/9dQ6JuNcwsBOV
jjfAiO0CvO3H2V7SV2GgEKljWWYv2B4oe+NxuxVUGlqdq/2tl8x24ugSW7Zji4Gt
BhW7vfkuea4U+343euov8yrgZYraglCQ6rX96G/R4yGH/T73cM8kvafwj4RUVzCs
j3tvW9FJdJelI6H2GGD21pyQTiiBZJDaZSM3klkPK6EGzd/XcghlS1wk8hxptYLH
oDzSOzETkxn/9qKEM+qNa8v+AwGX4v+BcmrS0gbwBV2qVqCgnrzrB9fmOBybGMDW
pnmXlaAlgasTHL0jtaO0Tu1LuC0GcwlWYvikliDixsvxY0cyuSqhwOlO9convvIc
3ykKA0XDPeG26i9bpjrywqH9OZmTiZBU0MaG6bqu4yN2irqz/v5K25eMC5dRDmKK
RFYOWh4M39tkhVlTsLmUajKUErjUJG3SW/9nuVR4C+advXIkmkxuIKHGbT6tfZn0
slq1ctJjq4jiDYkTTmtgYWIFO4luZbtLK1TYu1CEQzFI3dAHwermId+Ky8HSy9zN
uyEJXrD6oi/kvOiZ050ettWvZeGGU6oGuobF4jKotQ8CH3tytyHeE9w1VHw9NB3n
3ORnqhGuAVtQwbLAo35PzbtVWIvFRKH5lVxUaiYTMTn4J0wY37yDAjvmZHPHDoPP
cxWMRA8ukMrr44TmHb3er8ZTVnyGKo4+SWVSgz4iLBMRBwJTkefTkMMjIokaXcLm
R6zaP8xJ/rB6bAG03y85zqI8AsYL+7bJVy+3+WkW/LTVGWQLYNaUf3WFxDR/Cv9K
y5ZXQuU1q3hvViSir46i/r2x/7bfxBwSI9uEAWm+k+/fWlq9Cdjq8D6crGlzdc1i
uFq7JkUf/cpFTgU/gFwZ+5tThF3a4txQ/J2bKf8i8Vu/lXWFgyn6iodrW8XUKmC3
ykBiqCQMs2osniCkT1ygiqX92ZIvQSXSY2I4M51GsnrpwbGqlqt9D9HRSxZdMzeX
ZgjfElmrWrj4ta7AhwIQkuPMyqbo8o1XmUFRLOuiQSryFbEgCY7eRoExUmykX/Yb
wDeYcJyOdAbmU3mruQjNHP6uRyKC1sHrZVr3YMOJKuRXLYbaPtVWPrZidCDV8ArC
XWkQ8TW9XealKyM6RypwF4CBhBJy6amNC5QjYQ+2U4xz2S5La/eLuGq/IjB+X5o6
eGLsouYXnUcxPJgCjDDathGzNSQDs/0d/Ch6NEZkQvh88fQ30Ya9yNDyuRFxAKcI
MtcyelP3HyE1VUG+YbmtkjXKZr4KScwMeuuUrJu0jQIS8bNDAC4dBaHls3BqxCZa
UBZZ5JcZnbXPHF/Z3cx5v4MtUSz51gSytRL2bodPwh1kqsOUa2DWBAfzukVjBtUl
wn3YuA9NAeZOYT0wtLBpRtrhIU+z9Gge6Dd6oyoTUU3sMyNAkdtQ7PIRd0rp48Rl
OGrhBfhWPaOxgbLsdJikRgwCLnAM9g4EeOveE3OVeRZ8MXRkp4pNhtRkmlG0gjUC
ULtJDpsgEGDc48Cxw1XLjA9yMIbfMZMcOM4bEiXfDXTqajYsgNutdV2ZVIDovH9o
Q5MXovuZ58irFJGTpHBbYubKsaGXIiRdzwhaK/GvlZzVZKVgiGvwJ0GEWhb5+V9h
OZ/VvhALs6G5g2aEH2wr+n3KSYgUwFOd2A9EZm0l7iq8CI93Llp9HsLiPG9L2Z4z
3jxO9Eg2lY5qG71ghDLgQPHuZVQaw7ipqA3k9za+Nt/RxyJg1UZHWywoRG6v4W3e
TdIgGJC0RhkZONa7w9IqbmGINCXzVQiJP0VMe5mTkUMdWBU53dqTS3PI8gjjhP3/
6r6uwej5AgHtsVqNrnKgHCYw3SBfkSuGFLPgte+CoS78iVgl/WpCGQ6zAoc43ooJ
czt4DyUC+VWMn/7IDx6xU0LB/lDXJmB64Yb5pB3b8hGTwW5LvJZpDnshXP+/glD1
E0Tb1FIHNHzLr/mjSrbGScYcb8ECKWmJxnhTULeZ9onDLuRHcKszC0asUYcTyvPv
3PGxHzCHKuFZxD7bSqGLqyIdp2C+JCjokRgiXknkDk3w9qr3apAu7hMqI4J7a+L7
IKHHHRXVYxrK2Rzs9N2IMSUS1fiLisVNeVDL7cytVhqoVrGRue6D8dZjAytyFjUk
00P4eEXYTOpsJ65ahAY0r9LB8Flu7mCoUWubvMVrDnv8mNeF/3JVLSzZyJtIsCKE
Ij8AfJSOiTSGyQ0EenStCgsi2Pa7737a9Csntq44PfQsGAC6Bxnf7qLadE1Cyy9E
z7ftsm71YELzZDSDQ7dFCfeg6lpltLxxl52acFvA4hsLrsYinOW6XBHwQAZHl5AT
EXCGc9Deal3iNgmpLT9hW2XI+y60yUUbwJ4fWiUjhs5OxTJLOxKN1yj7DgywWx/4
nnVYjAF/cXJHei1fDkMfRojIEO9pPOJGfrBIbmlhYUdYO4tSvumj4DvOUNIzuMCP
sSJvtKJ3EIOk87Yq0cWIUPef7HaC5sH+pt8Qvgd0UjBwzfifmQ9RAchJ5T9xub8Y
e73S4WvCzqAu9S9i1bzTUUnXMC+I7UNO2q79rjqhJGT0djsodrjH0ko1ega/sec1
PLJvUe+68PJfrCk+76lGIHMrgej5ikqIWbN6fu8AkQeo4aJyOFD9gtAAJ5XgZ04Z
fNssTggFiSL2DTqXbDnosuUsR4kd7E+QErsUj3TJXeDR7np0QzXYj7a/VonVBczW
LJFOk1zRuD1/DILU7rxm9JSNlW1xyi+7b0rWT4SrxWcKB+T4t2IZdHOs9HjjqRIS
O90FHKknVuwBXrDnALJs1+WiZAxcsdawjx73TY+Va3WcvLT1OlXpd4r2qb8DQpXH
69PCxNV+SKqE4qjlaLWi2M3ncr5bbSBXqn4ZngllxaS0tZ5juM0wDP7efwdOqjKU
tx27uDt+Xkn/XWmlmTg/Rekm5q3BIqhh2jI5/szek/W0hqF745w29jXtw7+p01FP
E0BNFKFu5OCgj2WOB9WiKQy5h7KmBJAHXuEy+Z+SAYiY+RtUgzZBETlwOYebwd9/
E5zWZRyMelukcLb0a6y+1lECwO5CAdWa0ctKEfksuIv7PsGSaiUJUCZXgT0pyKCK
juGvwXJYZIKM6M878tOdcUJa57q6kPXeOpbNMCMus5YY+ln/Gbd3ARpwsHlmQpyD
3JaB7RBNc43XW2hs7//C92KJ2D62i87ACOh+7ia/NdXfFmJ/wW2frGSNTfGUiLHo
yhiyl3DFpbEtCzJ4D1vCOWa/pwp5AC5h/QK8I0+KXLSnQm3Vim5jpUCV44MMu8ls
cGbvP/geHKrVPtdNu9T269zngczDOX406sf1ziIEHcO8uzwpTZCVJft6uL5DbwVC
+Sunl2WHgtPoybyT2+qZJRktDa4Qpp/xkVlydfijdYijvh/rczotfx6sU7gf7nlg
ruO91muiiotnacfNQTECQyp5w7PYKOrP3H3/9Wmmlg3VO0IUZW2h8+cZoRVx19rp
r9YoA0TsNzw/a1+pJmFi4/cSPYt6jFUUkuaIOF8f7u70ovrnbyPn30NGbtHjzJeq
WuM+Ux7WE4GxDJQ1IBzwjI5Twv67g3T34PkrlZvMgEhczkjxNdgPccw47w4azfjd
U33ykOloNe7hRfIFQimLAeijd0GyZe1j8YMBEcve+gUpQLWRLfvXNuXBkKQAxo2p
6XuIr+NwZURpcC/XEEdZitPdFiVz2k52orsCLd34h7iuYhJYDxogBKBQOOSEBDTv
Hs1mm8I80qBlFY78ngGjZEYwH8m+S8L+yuqbClk14fnEzGB/35MY3OOyav7GHwgo
svJ6+LcxuX2dmbAjYPR98ZqiCAWLfp2naHFHx1fAlwEfzjlPdDk0Z87+bJzkwOhP
8aE1kVov9Ku52/omhor2HCLpvZESB/ljujFDhYoE9r5fMJBicjPzV/1sWcO6IUUf
OeIdBpT8nxfydcKsdlCPhwJkkQo1ZcmclVBkF4uecQWoa4mxkAGNPLaZGDildtR0
30bU5eDnWnpkLweZolQNrnzFKtLTmfpaATtx7M2A4RdVRKjc5x3rIspO+Ab79qs6
VNMsz9i1mXCnBavh0+d+LVoD22Wj3lgml2slczamYZGte+omrkZbMZEdlCH7SLHR
UuyEEd0bFTcIBd6nGpUwrmkTCtEuK05QaxjlWZujwnQALpzhqF35niJRREaMxB95
6ATD04pIRWwPwbRIjnfSq8RAwqjlP+8cmk8M+oOn4JijL1SwSfl33KdFTMtCepPJ
3ZSPolo11Z8X5jcEu5AWSE3JLBj9Oza77T3X9nmH+0qJL87PsHkE/2T7jDq69J6R
llHziZbKwuHooxiohRV0/PKbCAWACHT9Nxht04eY4yzDCjV4ouMe3PNFo2RTKevs
uLkSUSj7/zwk1+LYzgCGhNVR/8HrdTwgHiiU0pZsdvXD/zIXhUKcGA+NxwPZj1Qm
S1olwFo5HIVH4N5u8ISXXVQSZQVV5Isja+5KJzc5TQXCCvh1wX/QduTaGDXmUrDc
rQFGBZZ1uGHO8DeNkthuRaFydv8vIJjmT736Fm+GsaRpcWc+CWWuJMQ5MKIAAptX
tJ5XmAFsNsL8ghPeapTvBlVba4KFUrWJE3hwugLEW5j1EXQbxHf9dk4Q/rxl++Fo
MQX+AnSckMvMNr8oIVLlqoTEv1b7k9iMmzcElSqi5veKDba3kiDNqwtCHhsSOfjh
dR40OBlTNA0Wl2EihxNbWVqgRIbT2qBsowsW96o2ILrfP4e7Re3/8EMOgofCDokn
SXbBbjpwseKl9ktvAbUDk1DUImhkiJckYncnI6GE1hruvNXyVLIWgKGHmIPQhGHz
EFeUZ8iPqYnl8qiF2pLdvGA84jAU8dO5QvDwErcRxLO/qf0MCQN6XSihJ1qpxizD
oEMlEATB8/wCGcvO+bpb+OQ0Gkbp002X7dZ2jblaOu8dfLNNMpcBOHfgi7vqubji
W+kVKhgzzSlN73dqwstho8qbOog6AXkoJL0bo7s/ayl+VQCXSGda0G2XGnOUWcAq
Myrul/en5/3kWBTnUR6hmZIlPLpFtYgGGBSXMz/x8L+C6axP9UULzq/q3c/e2Y80
M/pFxdgPXwZqn2bW9ef4Ntd6LQ4ebdv6j793gMhQAd4q18gxrdfi6EKw+J0g1m+X
AQrMWbkCUqKGin1Y5ny8U86C6ZMT444aH+EZcI5wG4o83Kc+ciLnmSWZfJDcK85o
4NYbhF/BZ63/LIKnBg8J4Fo4diiDn2fliKxIFA/aDDghIoykcayiDCaAgZ085UXw
iap6mhPIyPdHX0kFhED6AwY5xrZo9QdhCuQME3qRyazGgGSeiR64Ap+aONjqxiNY
S9GkHDWesik5TxSpbhMtDGCQnLduGTIyR8+knXqy8NQ+pD9X5GuGVodBiyTxfgGG
cxFs6WyYN7eS5PycFcbSPxO0hpHVxy9U4yvdoK3yYZgRae400qIfuqAIis//5XTG
xONQ7qjvygl49Ar2GA3f3BirP9JGvpiARkHyvwAAILGocKN3zNNz5EAIodP80ZpQ
caoWb/XqwUSdMUMFRGZUtd7WECvs9M350VS+tt5bhqd+sjPpCDdVDZSIMBZ3UdbW
fY8q6X0ygNMiX9e8nnuN6+BsVtWIJGIspOaLFZIkBFSm3fZsZ+AV8yNXaUpYcx5W
bNAKArdLSwMoMjEC1dg50BoAEB0Y1czdPM7zc8RfEPDDD/uffR3TGKi+SKDs+ZEA
hU0QWG6z5Ojs4a57gUBVNQ1VrhAl7OL2tTzt1+bso9xIE45XQH22TTM2ynOuDOTs
mHq9IVQixyipPBAe1cnoASyHn5u+/fic0nAeBD5MB1mRdaKMW/t2PMmPHmZIk6bx
k9yC6qh105yeCMOS2iNbHTkg/YzL6/kryHjW3e8MEA4Lv0hO7Nj0vPqFVMXqQjjt
tbugIY0dYgmvzGT83Avo9dvtAlQg0gRVj84nT53OKISfpP1jjv5DUbSrLeDXVJ+J
TVaw9d32tuteJNMPO5ob5ytjtcBS7a2Jg0MnvlcdswjPdyxqyvkaQH+miShRwbYe
bT99ewT1bxOzwCRPYYz505JFMMxU47Gq+APc6DmHFv/CM8xpkXIXw1g2kKTE/mqU
6iYhqZjzmJji8Z6A5RsFcCXW86wb4en8lWg2KIPy5A48VZAHAp0IKGC7f74b5Tjz
H06QZMEnHMdjQUeL/YJip7zZnP7qs5KsO3E/hNUsuNZ+IwNoklhHwiGQk5hI0M7z
3B2467uN+K7f3mgPAYaEsFVEIDmF4CJ8037UGKS4peT+NcXCI+ADWgYnkUg6IJTw
kQ/LVMowwvtycpErGyBwKocRWNOrEogNYqkFIm2B9t7lIpNVYPfXYRn4vTRgi06g
SYcl4GERydX6umNPfWGJ3w9xmCx+s7BSYnB0ofjBghczQEmOCyb6oQk4Es8SX4EJ
ItkDb9UZUcBvT1VGcBfjkVZpGkZR/fY4KhTWE5eD2DFmZmEb/v10jUrGFHwrenhF
wDwDdsut7VLY4wWvsfvEMgoUKQFVGnUa9DdDq7oQJlbiV+Xvwlof/EqTBaSv/nXH
8jjQBtzgjDuHVUELY9We0/S5hedDJgmO1oNdwFcSmVwc104enEe0wLJ3VU72lu5d
mjKJU6gGhjkjQfDk9jvZjQ4or+gEelTD7jyOt/xLaH7/hNb323X7OwF1yQ6QrjJn
DWtqe9GSrXAc7N8ZaPdfz+o1jXnD5fcGyqOiescgf43a4VBA/3zoUWc+xJTTRMAh
PBWX0kseQEs/BbGIGYwTNZ0Ayhh6uSpaDi8IWJuC3N4NxuyQK60J7ViTIDrcEVqV
f8qzPzKV5txzyRCsgaI94JPlZ9ckf8LRnGCuRnaWfyZmFtjuWmSoCbkBZBgv1mcS
zrf5SgQPdNWwIgQLqt5V5TGDD2/Q0R22KMTbBoRP1vf+Ol+Bes3Ybngbz584+g6h
lNJPlsqMOnHJ1mYaiyhiExSfHpg2jXI3r0Kiuq6EfLID3jGXi1c4WdQb6/542w/w
9GSp8ewPKBI4MlhYVOm86LNuBjYo2sZca2ETdYfcB1IWnTGM2WfINceHZu3jfwbe
wpwF1klfrBVZVaBESaHzQD1Tc1KGKVwXn8sCKU8L8i929T7Q8+WGsc+qt2U7RZ3C
Sf//G7gTP36doQRDAyo2+OK+Z3Rfmtu7D+pXbdl+lEHvcV8AbNl7XhiSjfiM5V8c
U8gQHl/6w8mOMYVJkki3aBWA+Ymupx5+gHdyUpDUNYMoOTNmRwSW5wwAsxRitdPW
21sbPhELdisg3YvhG2/J4G6gZr5pwg+Qtqllv7ZWRBz2XvbIbGQhkdN8zEPD0+rH
enFiU4vHb7k4uVi6GDD4IDNJ/Z3udv4L9F7NdKo2YQeg8MLfLa4SbTvHIA+bmpEn
5DVYr9QDg7FybIgp6ojQX89tcyI3xxCNMwaSyxwbqt9zceKaPSjrwAQ/X78xjfTR
g06OA9s3nUODRCQOzQFexMWTUgDnE29uIyXwuHrV6+qvQxT2VmTGlFq9wjvbjPWM
NMAvqrM9Jicc4nmsHJqSmeHXSG8X0l4DRgPbn9rIkwr6qJbgAjvXtF/qvNzm/VF9
Oe5bXccmWgfzEt+OF5ZMhELW3F7xqbZ2kWySH/jBovZLAnz7p3QXg/b9eXYG3gAw
4TnJF7QWRjyHRLC6oYWbWaklW39ZS/0Sc9x06dXhDLPDMiVR5CUR9Vq7CXMdm5tO
5xAmfhkO3XKJW67nghRpckTdGaA81kwqWFvEa0DMSdUhUcWeQLgLKbg/gch8PfJx
3Zwbr4ktqCEAQzvTBi8B35aY6El87m/j9p1R1TojVmWeboeHI9ASL4ef9QPL0PQe
6Yorf98FEuNG2oFTMloRVaQwxg6KCdp5zwg5yD0AKNVHkjpArf/Q/8qdZHClETdT
1pM3jn8SUfM7f9ZqqGoNJIWbEKk/ZMbWkR+I29XtmEsa5L80GPV4QPrUA+t6839k
xOKL2V2sFsgcW6+bea14TWbS+UsiCMH2PG3w5sJymUeKl2eNHYTGxqM1Qz8tRkiH
g1k1T2G7Gcaz1b7sP8ks089kvzzVDc9MxiW1EZ2m9mdiSEqotKDMraztn7yHYDQV
uevisp/r9d0fl9VEDiAtBO3bzAiBVmMsyRJ0YAl+Bck3wEm1pG9vSJM4qxf41uSM
U2TV8bPr2N+7GLURjs9Y1RmXMmaV0+EkrsZWhmrX2cqlUI1pg1MexITla97Qaupr
SEYQ11JP6hfC4yxmlVXmN30LWxFSAJpAHl7MRtnaG62Yrni2EACai4FCMkZGFsek
YprRWFlEZBgSehpw8rl+KZnwXUb9k5ZaoSzvZgcxPjYiaCoZ17STAPbLou2tRI0r
tfh8u6V6CwHgma1NhLCud/aIyX2ErVrqMWDkN+7q/oalg4w8YulUXhgazRb9o0mq
iaguyttcAI7EPLaJM1V1Z4GgC/7tNR1IhWJdiH8BQ1JLACW+Ll+QKoaqOQRG+9Wb
JKvbijaMCAdoIjdakFHS5CtFgvEDhuHjkyGtQ4KL/tX82xEJ9o98P1lMRRbayKc2
8lFg5KVrOFtF9GsGzW1FhgLZnfdFa2gD3rq6EFYOjhl4xIvdqnsaOAtqHRx/1ASK
kY/dJtv+9l9WEclft09pA4sqcqreiszvcqu9/olrakLFdn5+ONJFQgEwf10L6Fmt
BVBDpLEM1qcCpg2ZDQTss0WXEMEwQY/3gIvP9JfhPPAXapQ5xmGnLbPbHxtngJ9d
+98yNqH8uNSRcR5Ky0VGFNHMqbQe/K4rsU4UMr/CzUT83gbUg9Wj3Y4WIdXU3YA+
S/ziNMpkUiR9duI9VOCspocmxZYLzNS30Uu4l4W5wKLw4/LkTcPsxHwWJ76Mthan
iNzwYnTgcYjXQnzmk8GwiUdVymb4Fn/Dg3aRNtFpnsCLv4RQAV35WR6F6JAeKdiM
7QaYiL+HtQauqR4XvPjtObRK+QLASK58HTLYzqDizdDAfQNUrOzt+dpxYSeAWF4k
y8gvDQMt016wxESWSb1sqsvk4hlB7KHbaFlnS3silbIuR5JxZn3R1YB/seV4CXet
nwzetAklezs1o5rDRj/I32WmPcZLIW2SMJkbStVSKt3aeHHD3o1SYbVCVJr7aVyF
DgCLXRuQrY4/efHtuVe8M8H/qyed84cSZIJhIaiE8Z9kMbeNcWgFz9YsWNWT3Hn9
fuRHgTl6FghphUtfBpXBsRk3tQYx6ra4lWsWNhzohcyqrll/KST7St0DMoWP+Q+V
JsHvzDT/CsJMa3iVVe4lyyPbqW0rESmFN1TgBv48LuIAknYmjAFamV5i9LPGiMvX
Sm6zGdLzvogtLhbxNN0QgGZIA+sBWK79zo5g4YssEtBvP/w6kS0i+w1O+acGeSN/
lXrn5g0u6P/eh+FoWEqX51NsCsWGvV2Wo1eH+MPfO4/SXu3/LaLlIHo3BqrLOhd8
xqwIMn8la7Y0pzT4saWMxDRdofzdy16owsLS91oxKcosmD2k3eZferHdOjTRd15f
ZbZ5Su5Puv3pjmKTvib3qndKpy+xDAaIwKjrabMzRJCfqZc/G48KJ//RTn1g9ase
THiR1L+N812u6jfHgAiBi2VOlLkvLKha+HkkshYeWHD/Tqq0h2yDd+HQ0C9ioKWP
mxXfIITatu+IddO4uVO0TLidGD8wBwikRBAhKOgWICaN4pC9sfk5MguZWv4KbhSv
0L2ElugiT65GXCIjCftTFprkA2dIu7iKasngMfVcpXItywMhyuSw3t+wj8tbvf1H
kRE848wwxfSRXob2N+xWSEMFm/R7wTnRO6B3+Mc0CmdRJnwFkmXViqROSTqaGIFo
iQHJxJahg1PITjz0gGATIthQ9sLQtjOf/IGqbvwUD6JPz4s1rptduA403ce2c1xD
DmtWqigpbu6/qc2S/t4PtX88FWwfSbEb9HmeyGPWGkUKQ1b6jScPn3Zb+/upEfpy
pXJpMTzQCTqnAJQrWHXza47GL0SL0arjN8QiPPXNeAhKdnIVcZZFT0FtpTkyNaru
MYXpIPb75UCjbHK9mF63jZEDTPQ6drlqyoF8QIDV2xsHfG6O5CsrrO6yEfczqySi
JKN/EsgisU2azhJ7Lw0EtbGZ1m/EH6uyNCSiG7hh9omG/KvAHDqOoeIsG0GFcI29
XnoFMlFbT6BYjF2/CUaP7En6DbtrKj4q6xrlDndXeloaw30K7rLwBWCnE2cJ6HtX
Of/gpyjzYfV8rSDPWNaTupkmGxud/M+KQCHOaRD3iosmWzrTU2PdvMDh+3bjyvYv
6XfPIxFch4BAtVfIZj6WMzMURyPFGtJWPROZ9Xpq1oF6PElqQvy9A6whAPefNyF3
zPfdfd+h62jSajYEG1AKc0ya39F76bYduaJJOXMBWxMYeaV4pG/G6NS6IozgYcYO
jBEgSATTjfVGVom5kyaysfVarInfywHi9w+xhW7ydC9ocUmueaR0b8LOwJWfYJYR
WS9AUXGaOhwJLFCtLxLnJDk9sM5Bx6L0hGqmARGP+KuHpY4qX8iaWwmIVEzg5w+X
Uzhdq1Kk5TL3PJuvYRhsR5Ma6ygggG7rQpOkMQP4bevNzC7vApWFOSJ0h2ooWRBU
0cwhKM0Yxi0EiU1wIoWq6E8cFnBBgjSaQjlVT6k6R2o34JiXJAy2z5ujJeruYMYp
8Iu/qZeryKffOsXurQ8ElzQ2AgehbSZe4TGcwN1yxfmOkO+tF2NaSqx9So+fTZ7/
Ks8HghzKAjL1Snhn5c4no5aAGHwXLG5PyDbR0DY/8fiE1r0fOZY/6/AwJoR2dKyf
H3z/QvGQynYj46M511w7nBbwM23wOnG/QCqOU3JU1IWbDXSDsxoL3eF9aGVFLiCd
z5+jzzAj58UnchQFUbjwHRfl4T8FQpmBjAN2/DlB+EjsGy4s7Tt9haEIqnF44uYy
JiXLnX4zf7nHCPvZqgQ5myTHTmD64rWNUjW4phd/1aWfZVS0BD8hy8mnsVAkl5LH
miiI60a58hrN6hjwCwM+TU+A9KuC74RRuuKcbDcsKX0cinZwnuspKnK/1+crOOSY
O3bkxo4r13DIZBIAOWBvhU+sijp75VkUbZK81NImDyajqQW3DkuwbjyakaouX07p
qMpEdszpH7FkQQTAs9RIs9bUaIaxeR0YhQW2pixaG1WLQ49o4YooyhPQYRRnT1uK
2M+15/1/oxGhQmIVviBYmJS3+4jzbj3HMATaJUveHGO9k3ViUmY39JxKs19idRWM
WmSvGd3DKrR/eFl1hxl7sLoYeg0EbJi/JdX3HWL0rbm5+DWo2BsqStfGozbExOjJ
BMn5hkpGlzGgPY/S2jwcLnw63gzvcauvSlU45r4Up0fmvWRCWcSL43U41zEXc9g9
BvW44qqldgAY7kKN6z/LcQ9PiZ+uaVaSqDpScrlnPXODNKf/7/deSErUNt1X4DOP
YUqEZ+W+VCYRvBLK2NALJaKD81B6pFgXGdZy/7o3QPPlFHmiliOZF+qcV509eu1C
Gkz8vVWdxTCEXKi39NNQ7IZnD5Vv+40lTsupDPPS0qNSX2WpcYlmhXLmfDFCvvd7
qY7FojYECELTCFQ/N/E+wkRSklwz3WSL2UjoM4g4VWLYwKWxQehfho6Hjj2v2W48
N0a4RtQ+NQkj1QwUmwH0NBCRRPdCeTa2JHgukOy3rFzTnewEdaK5xkK+ZfUYgUsW
MwlH7a2Bkc5Ah+BgoHRUsgp5oC/0l3E5PAEu5REfRXn9THRD6u+zTzDb46Ib8gRY
gepqC3hEMZtlsao/6H8bL9bQYTtwlhc+WKILDPPbIHB8nVYxiUQ1BoSVXd3uDjyk
Irvs7UWApGGc8u8RBX5H0suzdo/8GPK90GMZU+hnjgYSCsGR7356P3mam1AUM0eE
GSxlZVeCJdW/PycHtNn2pBaIAfU4V7+OVozPdL0RGdeqNRfWWQngx4tn4FfijECr
4xY4ybyWh406avH7ZIVl+hI/UeRLgV3ISgdJ6iCWV87o7fZ70e3PNaZchOdyPTJ3
0AaAVupc3hgyz4RkghTh2kXgBSn/1mdsQf0LJtxEjGXuJudB5sPOEeoLbKWybw6k
YKc4ibRVp08+SMQAl2n2JVWv6xi8izgFGP/k6XAuS+wA11nYkK/7dMfh+dwHfwkR
qYuO3C9f2ZpHlIcVvk7hhhZDm19XpR2nFGlJZmkfs/AmYY0XRhlUfMyg/q82DF+J
SCQXKx7/7pIxliRdjtQ1EjV1/mDarWSh5ikRH/mCkOjnn1Xt+975OeLqvBaVBLOt
o0jWbjte9Amr6mArlsgBlIg/806Hmmr7Tnniki4VLoU5qMC0iiWiyYfSsfB7uYcz
Ja+fdAOyqayKpnIbkqgRJ71tDBNRTocPzYZBeM/ouSen1/iiufOv20QP8+fPKc5s
Vxv1/H4Z+Q4AAeu2mF3yl6iy/lrETvItc7iqMyXyUQWljzRccvA3PWRscchrW8P1
n3cMXoI/WkgL6N25zpg29n+wLLbP36hDNCUbtt/6td4zf5v1Rfv3UmGwdboL7fPj
I9U0vImYvpac/9QJPrprXipwRUh0fPuny9Aw61PRBItR6cgSiA1He72dCdgcGEUd
yiB9zhV2CtCgXdKYZeDmX9siYXKwHOYQ02JpBke9pU7qupMxOd13FUvwKRD/TRWh
9xLF7eAqPgF0whNNU9ajPO/60TttvtS/aM5Mq0VjpVAA63wUqeKv+W+upgoIlhVf
ZrQIWmh2tpNhxVeFEasy7LbU1R3nu+zCZI9MP09z5pknDS7MyIpAPLzjWW9HBrad
OXweirlunjAOHX7F9K51aN6qlvTxV43JgoUoJR7gDgsq43EdFppeaKp6/dykylFo
JvKhZ7oOeJyhDorpaVgzH8TLNX/0wYuAKiBAmsot+gcIR+AJYt8ebJWWwKhEv89k
OhVnQTWFa8FE0yGFIPNML5bNNta4jtkX7Jgpfy3kvzCdm5qP20BIst0TJVcly9/H
cZ46MHpTB5rSaJFWknll2oDuYwSwCT4KuNmXvKGqsjxM6cIbLkoRvtmoIjVOgCWA
y7qNbodWLFGo62D96nmDvEOu05LxialCHumboFEk46oLvo/SWEiSHqeo+uiMkIzK
ekm92k3/FW30c+nzX66qk3b2MzFRPAaFZQFW3pJd77jvTWUgLPef3Oz2yGWJtxpS
VBIeM3KJyd2Q4sQwqB5z0iuA5OO0O58YqWwkmHfeV0LnyoHktejbIf2X5exVUsSX
Gaww0iSj5nYOfon/BKD+6ZnKkY1WrsSIQDfZ8oQPVCtDpD6aX1QPqJ5sNNXvT2Xd
G+iSOcIuXtXeLO/rXlSf/J5VJZlHLy4WWz/0VHsuIFuGnCbKyOBssnXe6/b2z/yD
hYjwAZkQMNlQ/9OjekOXeXauD4ECpKIG4S4R3V+ldhMQ43tVQDt8u6sbK4nQQ7gu
sZatipIOHra8KJpkcGS7zDqucxI4k3LU++bB0Ek0wuXQVW32PcP2xvpdUde3KWrP
QDiKsJ/kBUUYGxgOEslVqTK6yU5BOrficomSHyeaCM/te2fEgk3wVM7SmPfPLVwP
LsXq5s2vU9+v9eWoaMuaI8wiwJRvNtKSh2xp/FEjulPHSHWPTC2Axi/xdZAIbgm5
670AoyIkpyqoEJb73hjJJOvYPVexef+m0OYlX8Fg5hVx/FaZzuTTlNtQfGnRkPzu
eWqA/qLdc3l1wWEr1nrM7Z0I0vhlGy2Lpn+UpQTEE4NyDYLT+JIkZvhpXf2aEfxz
d6fS7iv4KFl8e9cda0mndksh8YVClqGUWWe+jqE93MfLHg2uNdaYZPZbW3DGcSj2
GdiLDnWPytG9UXRDqpQqMj5LjJgdZ3h2IQPwV3XzTzG9lE0jVfnENVa/Nj+EZzc9
WP/LNutTNkLy6i0An1zw4ngKFRrBSqiwp1mqX4MYqx81aO9DJXWUjFYGBbCk6HQk
0MuSeFuwegkSgr9AGYr3CGuqj1gmChGv4Frp0i9F79CsrfcYZ+cHPmfu2stcZR+5
T2genZ4UmEr4bLRDOxt9eGXnlF5h0nALFAYKX9+nKK39IbWMcoJRC0I5Jnk+RKl7
5rVbTkMKbimilnilxcR/OnnFxWGwwRwTXDyxqYGGcSv+h+7BpEuzdDlgNqzmMrqD
QMwqb2qmS5/D2/OHX+x49GkUnrvi3jZakw1YVJUK0KyC9QrUjhIwYf6ZYFF003ck
yMXd79ZoBtg3XzALmiwexwNBKAz6OaromXNURtOljurRT+ZASfuICYRVyY51hpb4
hY12P2ukP7N3x4DV7oWXur9WlQdPFDWd5GI0joOd2LRxv3OAg0m/S+2kpo6RNkEg
ZPg2qZeEAC2IkNGLFhBxS3M2DsyZLFYATaksEdJWjrHJD+iSAAtiV+Cig3t7uBpP
KvH+R4LkyTxlhWD7zDrS8tiowjx8ZfdqdnbsiibRMmoplcRtfMGr4a1HPhNkQXHF
3ksM7PIbn5SquoMLOEkqCtqoOgdxZG/n8XYbX488qqMafL5QhfHn87hbNFQbFiJB
mSFE4iBRvfPZ7tuUYLxjNlzkq2W/Y7ahXoLB/B8Q9zdnhjfpHZQje+ejevAOTSlF
HTq+ajASfgjLhcZAp+6iAHTWrwcw+iK2LJmJwAlsuf8JArWJyQYSZlAIWkY7ntv0
RXzv3x+Qib5rb0h3497k7oCGGJzd9UG0ZfmHUuXv6/SPgfDptU18WCzfb9C5IuTU
z4FZNtFHQH4HxsNVtdrKDgfI16VOnYwvLHMtce2QPojgLWyjrcCbPn1su/zLlN1b
tkg2lg1L2nXVQXoNSmrNqy2m75FK2du57nmJ7ZmnOuWRuYOyVUX3fLYfkxUJYisD
IwJMA8BKM36oiK1bJ2swiy/UidtHtStHK7SgQIjbNlgdbLHQ95m8AUNA6217dLSP
IiQ18CtBZsAOP5+btCw3z1q+w8Bd4Gxdmd5xl+ZcThznWmFFXihPFCrxGKWSJdmL
WZPRYWbgun0JAcEiU6AExn6V71DiONLVAolDs9Ovt1fGQ5cVTv8eOgNiAnOHJqo6
uzGA8c7ABsXo5SelA75Y1F497ZHwv0mkFoy4GRGVp+woKXgHUElxovJtnJhnmzlC
OCgVcQ0ZiKJ5wg6jVJjWXVyFNJwAuDFeEh7fozfGCCcWHHSVPGCzKwSENeFd9qhD
DcDwpiDoByO+Akr1k1K/iG1B6LXa9Lzb5uGP3kL70KvwvgpAYpTxvOKxANHLemgw
HF2rK9zqcAqGt919jtE/i2KKfo8plss7ffD2gRHC2x54TTk1GQRcFi0EXxWWTuJZ
pJjFJ6T/6hDyAw4526aT+loDM4igiBjKfagA4OOFKTYARc8HghH+jIefKR9WJiNC
rkgcmqyuyIniscO5OxC0sRVdJw/jbeAdJYtRVM9I0JU7T2SS0GTIiESe7UGMdktR
rcosNb7xzfxhKazJFCNf9IorEtAQiKHG7EGftCWJ+er5iJWIJmrdwuyXz9ob2DpZ
hCScCFblgpEO96HWXDTFNPT5CbTN915NwQoLtRuR7Rj6KY23yq1aw5tJSnIFYZlS
P3FoLEwaMT6AfzniQW0em0vwQZ+LEcHNGFUTavAaCvLm4YrY+Oqb5AYp//KTxhmq
tFv9gWt3fwm+rD+QRDEktainVlS5trXlYNoDuFixBD4+q7aa0Kaw2hUTChS8qjP/
yzYxqDT5JB+SGc6XLW0QDSAdjIGd6mHOODfYCyqjzJ/hm8eiGrqF30qYWEeBKaid
PmxlBuVfAdILK5OEZ3ymOJwcI4Gs/rXOzQQu5twLxXuZc+KgYAZGI7WfMOiTalm5
7uayFCfEBCgT2UG+yiB+tKB2DhvnUMSyojKKzq+KcCzDszm0n7VUmN9rwCXtZBc5
Nabw7kbysF2hRgEOO9Ip2A9d8iYGesivz9G8fG2Boxmu5wWeRNRwOiIGZHzVhhFE
+rzzfrugdZQh2Huuqc9AGg3p5SaDOCyy4PaugczKIuKeMlyxokLRcaJgY+NWhl6t
0gAtvUF7LKuUvMi1hA8sjNhe6XKhyq4nV9itLLr3WISO1moC4Hl+aOeLZ7/hQO6W
Gi+wYZq3/tUVKXmdtpiVPzxbRz0KLolU0CQuKniD68sOyS5+JRg01pvleUabYBy5
Qi0bWSzIjThz5RbSstcZPNSHVCgoMuweLyZK+hMPpOAUcnICnE8S+cDmuLWMsESN
LgVPe4meyI4nnEkLTyo6RbC8gdjb9mttE946WqvS4l+rGJO0BhrUcH+8fanW8koN
nIMkxibBLzR1quonsdku9zicAJk9xcK7krAjKoHO9gRMcow5P9aOctKy3P/ACPcG
YL2wNd9NPwmBZmf3HzMdZP8Ofk69+5Hd37qtGded2pykJgBU9R3EBNogIaBoLLIs
NTahLegn65UVyPPrC8WOYMQvsBz+vrMqiL1ERpPVsXJbTnKsHV35/zIsTnqHJ7lj
YU1WHe0J8tlTY/X+3ijD2CTfwjx3So5ZLbL2KtBGcH1UZpak8zjtfA9LCvkSAhL4
2MCDNutPF7mtCzomPjeCs1f4BrKNIcqspd+aVEajyPBkzZRudYVI3ZC7O/4zh9xn
jqZxP6mWRVyhHq/SXsL4KGw8RIUwtL3WBNpGCxMU2yXmnpYPjaMt2naoe2QMiDQo
CCjA6GIEEIgobB3VqoFBc0FYKy3jkgw0jy8ipY2RP0ERyT3iExDWI5kgbiHi3WjS
4BEx7iCFDFAqZfqeyGlGTfcFzPsEJkLCsRtQrbfCNLf3MAtIhmBa3fVkeX4CiSKl
vGGCJk3+XsHLq21bHUcoqO4H6wKeUFQHvDYuH3M/AM5IolbEsdgQVpHis7SOzSDT
nzTzFbN6NyKuPMkdXbem4m9e9g2eIoe63FmLMqGp0bIVJlnliaLV/KS3xNIr/Nwe
Up+kqc473Th7SP7sBpDtUcvDJLOfvFtilDYOHttGVJiOGS4vCwdJfTHYFh02pNb1
rhExUGk3S9Xo3pWW+GDrrLA666SMUvda2pISFGdq7/nteggp+H9yoBlrOAze22LJ
LO0kMF+hkQ3Bguqorczqdpw1lsAMdINyYmNusaE2M1Kto8bW57CARgOv3jptrMk8
c4VWdYq9+d/X8Xj69cYuJelAG2teVkSdSdNd9JaMGW/0Az8V0NjkPTVYWLT1vIOr
wvnWkFTL+dbS5T8CfDQicanRdxJets21etZgh6/KmdU0CvGgfNUHPrF6Y0kLSx3y
7W/Mtp0SGiWhxizY2zMOQu3cOZuHea6dE8CUxdvprNV2yKEiF19xvFsV5Ajcgs5j
xe1i2OCDm1iGRbJTbq6ptrGWV/AAwAWcuBdTMLoTDE+epmhjBBqHZeAQwnxbgiSW
uuwBQVgKHzTA3ioKIebztQLqF5K/pzgavTvw99LOf9DD9Rd1Wsos67BoABt0axGJ
yl9ZL+/C6w76B5Gjn9yJf5UUwHd5PDZK/tOW8qsQtMLKvZvf3CH+OXt8EDAv/KMj
/aEpDeSmLLaBHGRVDEqvXsaJcuhgsLOc0N5Db2qWJ7ietBwyI0QtusqvaiLwaU8i
XW9kzdvy1rMIlVYzk3BAmydrh/Ytk6+JpbCdrxrb6Wmkx/S9xPyBX/R01ujJYGCo
IEoSmrzKFhIwy6eHiNocM76qba/OX62ZCBei18GipO4OKBTOAm81yvPY1vWlDrnY
5XdHXjHN+zPsJsgB4TyjJBUYDfHh4ayekK8CIMxY1om+a1Kg5a6+3seEEvRTr3BY
0MoYbPR0qKLp7jgyVajhXuXmZoVkMlXYzMn8UMIj9RwmNjAdzm12oowDG9cDTG/q
w81YlHYuE7ZftCXxI/i6uNP7ULlteL9ieNwTAMsOuN8DBX1DNLlK2TFYtJPAwmex
eP6swe+Tqx6zzLL/Yo7wu/2rzoWBx5kKqMkZo0CQvsHrq4RbODTAGk+kJ+hIF+h0
9B98t5WvyLtwWTsjIYuaw53v9WjIhlNa7q/Lkh/VWFt6JDV4/f0zL3IFfJD3RxQI
tYdPvAGEZ/1svpAA8KgAI1pSJQ/38aoc0o0Zocoj9WxPyo+t9iq5Le4CWePdxSOr
d0WEGQbGUjahUOnuM4lRScd3RC5PfL9U4PUhYJ67x0tE0yMlgUrJIC2KgPsgPj+I
dHh63N9rCltdgBvhqKF3zDdwskVySKCX0OrbC5tdS67gn4n3zWvopDBnII+b5qSq
Mv3Q/QeR1i2uqE2GuByptRceq3adsHx8wi+O0WeBZyWiaBx/fQgJqCC88WmgeAZl
U7m+I+5QR/3hKVYidT+xg/Kaj1uHCW3/rjWBoRX9NuhrLXD/CMnq1pnIKlJWwKOg
sFOedfByMfski/EVZX9fkLF2rL0pdhD4Wsk97QmbewAcYqHKx44UBedAWj7WJ2W/
RcNvHRT/kBev8vBAB+yRx3xjgDJsYeIH6K3lt+kkq4qWoGlwb3zoa5dfmVLfrNk9
WJXqsf8TcOCJhwdSZ7cx+iQy8eU5EYfKsZwALVLXLcS04wrTlEUKNyuiZRBP9ypF
t24szwi1igcyIr+yL1d9vN/UVVr1fo68JzIRHJDiOGNHjkU99vtmnDpuvzvTZ5V9
6X0YY5ccWnZdGXdH3ylLUhOWYediMdSUCPs/6vBedmzV5JxfUH2e4JTURJFgBZm9
IL+vBx7vKjYKD8tG8Fe+ABfTXG5GSP2yJy8va6mhexYeuRnJtnCMNqRO5wyq17oS
XMBMJFWmPe1oFyFp374nDLYDSkShR8i+09bYv29evh3tn7m0P92Q3WsqSpCHkuIC
bo2T/OiN2BTO31z1dxddRBU8fjiZS4r1qXq1sGoB3ITYRC7+b1Me8VW5n27CdNpZ
RD0sCVh3U/LbKINSBV52oAs2ke+76VwWN5vFgcYbaftXmGo39su3LYNBV3IPe4Z0
+Kbc8GCSUkElR+B9oztk447hzoJPLIZT97dCWxNw7x0W6oY6wS/83hHw0/GMOPLq
D4Emg0CTDCmzoiLcXn/fmbbovYMtVgq6f8Ugdo68ARVs8nt26nYhpReLJ9QN5qag
ETQRr9YK/wguLa4OPXAyy70fXxCwcOfyNnywE5pzzGAv/WKVN+jjxYzTilT1ILD1
S+AN0y3e4mmERUKIB5+5b5hE9vRGHDR8Dfd4VwUfuQMvfGpfYOix28Fvl4VgOq7T
gdke6VJtaRgLYjCKDPhu8zJ+CHBJd49kZrxmedmeh/k/4/kls4CcYksItq4FKjbz
7dLssDRewlcvhTiQnWbRJnUIrqGvTU9+MLxJdJ6Y5CEqRIRTkgTJlUsL6LpEwtCO
LansgTIsYichG7kRFfNsxdPXaaYkn3Nt6kwqKd/xG+1woYdeFApFudOV0WRv/mjK
yI/Zq+8AETMKZ+XXHpII+FD+GA0DX3l4gAkAfDqkF6zH9Zf8qY5mTPiyiTPjlY17
t/Oxj/CX1nTKG4yHi7CYVuKIVV3leCNeNV2loUXIvX9fMOkP0CASgihV0lbjXNG+
H48nQK4qSSvP4kGhmEYhzql5G9DNdECltR/fk5uslx9dEeUicbb2+j2sJKE9cVL+
YXOhydXeaa6V910hLkOHWuK48hmqYMQXOzMxYwz4RlSGJGCWMrZmj1qQOWyTxfj9
F7rwJFgJnByAOegSqinpSquMD9TChlcxEOS+uOljVw/XM09aDQpchrGnWly0nQ6b
nACq5zT6JT/+2JCTFpRkK8kqZoxGDTB6Qm4oqVbGzKVj2o7Tieq5yqD+IKw8nrig
QiSGiqz97+hPIp2cAzVWEmkJPbJZUFaQ4mtG+WqgJx0xSILMp7SKMZjYnW5anM1T
qY28phqQ/qm5KJJ0Emup50MhJJyUHCGhoL+EvwAGyx0Dq33yz3kmS8aJ6Cvp5Flg
HKXE4N8SNbrNTYJ1wmDmnMVRB2XZkah0k9OOwSHJU0v64emSLCxrfKP/6hXFACzu
p7d+ibviLII/38wcPO3LYfJ96ilMpyxl6gX+aRUTnvvVeV0aLF1fSuZlFBMNwAL3
Q6/jaD3gjzHsaiK+qhJCkcjf3vhCCz20cM5AmEqvdvr6bDssUqxtuiU5aKHE6zXL
fTIGUbzCFfTgNHQ8fvoWOsVqmWmQZq9dgKtek69uNME7VdOs/i1bTBIxCI34oQwZ
TWJh1sBExSx8KmE+8n56gPRL5KMKRpKILgFIy6AdE8RcbQHHPRZEuP29iDfBPtTE
mnXIQxIujnjrNobcmTGTVQ1YwpXKpS9/ROUncJ7tJgc/BQY8rq2BXrgNgsN2/qu9
RCAhrqPLCso2qAWTjFwMrTHTNQxynbNXAUUOmCHcd9/ry6pDTkaYwjoA3ekpQEgb
z77yFuC+F6PimQznqAWhXzWB4WRzaa//rE8dHS3PyphL0a7fu01Y9/iY/5psVCP0
bR/CLRT2+ARZ6jXtmfeforKpubYQS90vwFDT88gq6/1b59Usa3CPuXy92kAA4pNZ
E42+o/TtUB7QBfqKPhE/vNa7LLKyikjGEWdh5ziE6JouztiPB4fjiWYxJbb4UQyU
LwATCwckrzu8S3tEw1+f99bKMBDd4wBMeYkAZjLw4LHQ26kj50dcMdJzQrjR01vL
fwAjVDuYiADWnEVa4OH/3i0+Y+KsnI3+zRNvmrHgKXZVdOTz3e4IQ8JFZIuQ0bLW
wX6RBKCv1hXjeTC87hVH4zvO7uP/OLmMXkfJy6FxIYbp077HuMs9muUhrhTQLlrJ
9DFaKsk2JFQLgaqySp/tBzSfEy9zx6SYwp6aHn9TQaBtWIQlvf0KPhNYvYAhwhjr
wBEgEKRBrGqg0htjHYzkmj5PhrF62V/4/A9+1QUSd4ZyqJ6pBpuld4moXtJ1KRsb
WSBORGVxvvyYD/1Xb6zLT7DvBLZNR41WyLQSgO+fDba8jhOQas2eG878N6Xd3qws
iuE9bj78ZxHweUW7+vsodiNIWHckYXF/JiqEd5gLkuSJgTsGpCqRLiI8FhjnT4c2
YQIN8ZilfLHa3PLrOjS1VQdDx3HhsW11muAIMsOIV/UgUnF4YEpJiPpuN8RlJ9hE
9Bej9s9LskIDQaYTfUu75BWiTxJ6t/DRXVZb7WBYZOUOoKjXvvlf+8Qid1d46nza
+nf33IBlIKWsy9IakPC1ugXYPEVmcx0hi5ossRTCtWM1r4EuLH/WdVSFe+x2dL8I
md9K1oHml+H094tTy5Uj8SPYvTPNHn1b7wOB+TztHtQZAVBmSP/ohb2eNXONQ1L5
lXc3HZiG5VZptvO1O2ERXuQ1rNRZfcPfEJzui8W6K1smVeV5fa7NB6pRDUxNDmmy
kIvnlBBKVPuQ3HY1Lou4P/GbaqyZFRdoE8E0rCEONj/iKjzFNSRHSSr7H42YCeCP
bj73gfj/6A3fYl3nyH00vMMDn5DOhVfyzW2kyAiD0u84RToxfknR0fEAInFbWxOs
5WcBNvBsztfPrdLWiBuae7Q0+OD4IFjHg8/XBBw3QDuhSSO8htuY1o1ffBfF8sw1
W2m7Q8kOpejlxztC0TQj2xmjzXDBnKYKAHpIULdTab4wnDUN89zcuwmibHWSDGsi
qDAHe8g2H0SorAmpPNnoPsV15ix5ZVST3H/Yv6tFzbbJSXo03YUznKh4JEphIUxS
h0Y8UsJKgVnBx8Fvti1QQR9O6He8amp50V7vtlIPEF37wgmX/Wjgk8DKUaXsO2Ke
XKbN3PiMYnmBWmhm6x7xRryIEyQkxYI7zApLSIZG+9klHfQjWCXCkEJu6N8E5d0k
4+c685lx9UPvdYCVyv/Rkmi4snesFJQKrAfY9ItyM2PeeLSzG6g8lpFvw7uocDiz
8Y/UGrgfamQrDLOFGfAM8EWpurv35VcLSkJcsSsYU8iE0Yp7ZOKoEurfEZHCTnHC
KYREnY/v0KpXHgsa65oUOOb/jKNJvnTQ23XdFJdvZCmj4SrAYlEOl/2Flt1PmAcB
ljAGavZjpVvFWOIyxXUWqWKXuEWC+lTcIh0tdDd54DvsdgSfng0R+ZZE0jytIj6K
hOz/eaTKXsBs1oeJ/s3Dw2Axg4XYrzBT2lbZAgPboMJ2//xtn13M8VFJRz7Mljvw
YEZg47o0iTWJmutq2UUMplIl+57B/o1LQlzTRuTaC3AOCyBXcjxaLwZMo5AQA4Op
jYNaiqMTQ/yl2WnQDiDKaa3YU5mfxdpDVAcNbb9fi7uxU4/4suX+GXTC4u0oaAvA
R7VXWBmEATegRxcqvu+2e2Bt5M7UDSVMG6ilgb42nz3Cd50n2Aj92+J4t76XOmSt
MxkvxnScDiiO4MFx0+bfg7Y+SvA4EnPwB5IcWnvCWYimfel0kaYAnDec+MXEtq80
gv9xrYNw8fpQfscM4/gyM9XCI0Awz4fagi+bTvEjiP4rRzWr9Af6M/lTZW0uTZY6
NbokDjt0NJ+8+NX8izEod/bawkHcYfegeOZH7eMvpknoa21eGe5+ysAfvqyHUjFu
W2mX9QQhNrdAIGnIjgcRxgDq45/RYF8gpFTNoZYJFzlm9fOBnhSGr+5uS/3Yc10O
L6Bhx59OR1H/fDYN5wLuvvh356bsFRXRiq9ItnFJrqnoZFuL/TSK0YF8vDm7Tw50
DUKgpZNREqlGSJkzKyiqVGRs9oajTxQySKNznF3TlDGaFtQpTneQf33poN/C4kjW
6qVeLab72vpieS+GEfdQOJMQjj+ml2XHNMBwTBcMRJ/1mfOM+YRDB8VuJHL7Ec84
KwUyMlKnJqTDoi64uVr3VW8GzxW/76gfcXB3SDsrNkiQjZqesAjkw+5QfcscH4bB
/ZdwMrbnCAT3uX/30L6DPxGv26rZZloouut1UJyyPEZ2T7JhIy/LS9ar5KytqRzx
5O7xMuPAjccA+W2B1vF9Gj/W/r0YKVNbM2ObqE93n2ZPymZGqa8OYJ5qVBf6+Wnj
xKttW/43fSb2/BZfkP6//hRNYkQb/OWrc7gH5x1BafhV0LhnOU2HZQtI6gA368Zs
kqR/B0Y33PJxV1BJsYtXUU00yK4YUbs6WmQ+Z/QBz7uUMvZ55i02/zbXVC4PNlqT
INEoj0Ba3HPmC8lW27GZqlwe/vmLfiabtFbrPMgxEnN9ju6fBSdVrC3f70wbWe6A
Zma94/Ts2ue4NvD+/39DsgTTlWL5xZbjBN6fALZUMZXwIw1ge+FArJc6W7kpV/br
ll2rn4Kwb2V6JO4R2ZA6mTB1wBhvLUpuWmVX4epXcQS6HEvqCq7xGknET66Rftf3
skvNJ2Rp63sHuHJ172+EVjzAbDpSU12tFvzliji2nmP8DIMa2AyZeexWdlrkOkmD
3VccQfLp5f3EdkzQC0SHUNX0O1EnWhtTme6vjhd9h/fVslWfZ9Zr2EEdPcvPczgc
+XEw9YmYzduupjEa4winbYlGMdUleX757kAgIvnLR6o1N1t5ko3rrccGMugEO0od
MZAuk577EqXTKLsSDnk12reqx8u9f/VHQORvcgLa/SACvzcTKcE/DUSUlg6F7ABo
YVv4cj8XDoJzCMYFeUK7S62dAh9SORXPVA5+P7wPCSeBegWmRlkWBG9Nr0VIc/LW
WxlvPYSNnSGMMKPlCVtem3cRCmx8IFdh+3DnivZ0gowCie7Q1VAA+o53oL1Kulil
0gf1dy0zkfOE9Ik8eXqojkKL3UB5Z8c/jPNRSJjr5rUcZT6iShkubt57s8r0iO/s
j04UX3nPKUqVN/P0CMtA5FQ1vrL+iSaQ38GnX0qNM5HabTG4Az5bSqcFRsoIEPkE
TSOU6arzrpI4jcAUnFx4MATaSnD4wewt49MmGeAKvs4pegG8/a3loUJYLhje3/xC
HvpLrtJon9Fzwjks+9JYdI/IT8pVjJ2cPg83EgnxRxvGDeSzBTKcm3g/v+H+22pR
iFlHdeuJbIpYME0C9pawhORoFtXNhb8xysMR6hx9iW2i+Wobg2hY86VBOz1c5ceN
XE1hwzg4TQTLaMolf+UBxAtoVDZuxK9ZYveWEsOrCSPlI7kxduNq9zIYfq8jEnh5
cZLlFbRcI2OimQUfs1dGEduPSgDB2HVYULXB+WpDdvfNCSNBwMI055rK3L2mkPtr
kaYIIH1CDS4/2RPzStzmJhagLhJGtOJd7JzcxXgtF6BQKIpPJ7TPxOHwLZFV9FGl
vlArdBsE9fiPxo99XOu6oFinrDsZEKa8XafFMZ+vpwgiOoKpFqs5cdNE11hb8cUv
Uy6hYd2hB93LLU1CFfdjK88HOj96zRNliHUf/SNuo/HtfKqepaXf3pjU3HOVa001
CRD/6OM4n3lcWJedQHQJgQjMNjLbaozwvZaEXCL4C4y3m1wR66PiiFul0w7lmOMc
OIWNvFVxEagv/eywRWqc/Yo5kQqgd4TCWXhOyomLl8+A+8yhww/j1adHLccI9WK6
hu1l9Ez4M0U3xNEzwpqGYiHt0TAljYcTFHP7fwEpFzwkxeFCV67SdUbnQKuO7ViW
3jEuwwfNjqvCdVPCSO/xelt2H0BM2WFh8FfnoAOAC/C85MwpX6jv6G1UHcPz0lal
XnWECWYrpm6jUpxU9kAsLVMJ4VVhvWY76rAjzSGu6lYRUFcxusnLul0KrZd74PPx
SpBpPH8bz8UcvXOyWxD/RPmhmCeiG8qutsyjn0q06iJ4bESV1GycApieeVM9JOo0
1QfMUWQr+CCrwfggf6GkTAW263hIRitZ0osQnv4pRqEYx46xH7tZcx0tk0ftz5y4
lIjZJivaOX9FoBghV0OFJhzfrWvWfroi0+mcq6Indr3Kmj1hSA5PMPyNxh3SI2rh
WAMLaEoicBHVylTUk5bk4keZjAQzt+Mzh+k2pTLXIjbpPhurKuBBM4wM9ifaS2aO
Khg/TesQiYUquYHyd+R80dGyP/KwqDpcXJzjzAi7HA59Kbj7FljDdC+7c/j/U1/J
5rF6STlcwZgr2Tx/+L+4R749NNbfDdo7cNXT1Q3N4rjfq05tz3aGoFm8sb0RSTKx
mI0mfkeEJsf5AO3Ty26wQJQH0j7zKjfMvhvkB+QMrm6+t/D5rH2GlZScyrkQvTYo
Q0Z+l0cp01nJJnEXOHuIbbqR+XwtDVgz6a5Kwfa861bHqDWLry4NvkrXuW9gG73N
QzDw+GIbVbBbimHU1wueWjpupsbCO+slXAk9V6FVkD3x4q3xrptkNjXhY6Xo/6Zs
jIo2QekqsgVX8vN/IVhP6lgP/oP8hxQfWqUsTs8nhFq/B1gFFNpO4qIKKizYIGWO
r8J4ysNUjAquaCBlGGcTlnHUXrGDBS0t49hFT0sCp4WuiUNm7fSlScIgyjb7v+7o
q1N5+1Gr9cyZzbSLuDSUZm9Jlj1gFPq4+XpF+QFpFd6fXyTTdlHz8+abCk/I2+C3
VUU1ablXBbFDeDxdv41pMIFZU05mo3vYIl6MBDLUAAl1jsaN5oYAxKkA4QiRcAWQ
UqlsYtw4ZRISVm3H2h05pU3OhH0fUH4r6cbqMa3LyCB4cUhZPK5PveiXPPSbvTOF
Men1QG3LeTSsUIAtg9eGT7ry6AOjColJfQgxx3wB3S13541wB+642LOqJY/2MzlP
fdCznbQ4LB4bvFtb8buqgD1r43Kw6xLZ0i1W78cmmfr/+vlInc7PHdFF7rHOdJn7
1RtYqnbf8t03++QTlwGv7lYlWZUGdS88oTqu44IJXtKFEd/N7u9OlRYrxHXsMsVu
4S58noxl5aPfYh/P+9q81dMu1kAMQTqCDZi0rG4ynAyS00UAznq6KCoaLrLTk0FK
84Jvfu+JRm5aupdiNVn7CK+NTk4EwlG7llsCnRClfFf1jIcSFtiC7CPmI5x35taD
y6nRh3nFU3YJSrPFmUmaDJt3IA2UqWVIelU2NYUnh8hwnnzPjD0ijJzIT9AP/WnX
v8IFjncH8n2VbTkDan56yLfZIoFLTBDtUOAEV2VD+BFidbxOiOioynTb2wnH+rjJ
NmO5Q2GsEB4/BVQjURANmscHW02XqPkQevff/Um8xmDUff4N2obaeVvNq2Z62d6L
tklRP6J9u3mUfivp9k7XM44PbzQZbgAHo0GzD+cCP07oyzNrfqhQADM/lelw9IDo
9Od4v+zzkjztiPdvz8VzqPAi9rG51XGjjpar/4vlSNkgCW/j9ILoTWOONam/4B1D
aindgeuS124HYeWeJZh1tncilrx5z9mg5a+dHO1nZ/ZE1D5lOswP4QmAzhGZ8tdP
wo0OuipQye+IUKdXhyxCEdAzz2SZCe2XSNi6r+Sqjyx1lxJR3zXqE2KV36ivpGf9
gp+FR9tWmDGYTP7Ocs91TjbEuCGKQR/Vwb1dxTaDxALJRVhHSR/q04IOvofPktgl
9ZN2MamGIFFeCzzSWBrR17UP8YAwLSKfqc0aZhTQ59bEAcFAKyepbkFj4m+VvmgE
6bzvaSQYlnuWQNJT9tduseqL4pj5xHNU/gb9VRn/dv5hsjJj5dDKRzND0vIGj0dF
3/drkOADodgo8QavlrI9nLahf/6Kf6pPKZ+qH/+fpaiQK0jsHtbum+4fOf8GW/KD
6nC4Udg0I4A+S9dLfrYjf+BOt9Z20HeRZIRLRodUdF+i3M1lK4Mo565wMP9dIUNo
rFRTX3VHziCN0pn1WB2JlB0sc5jSFMiko6hzfw1UzCd7wHQLci5PpeRUhR3zC63L
Ct5nxfuXWCR4Fm359rfGKH28C0PNK2nbF6NylRe3wEu1fcjEACk4EqNw74wWZ/ck
+ieXB4zPh63/Um68s0ugh5zql5NIWCLBfTLVAyT86qzQV2z9QmZ/S1q/B8tLOs+Y
rrIZ/LJPvqg9ovcU5va2Wi2tVZhYyk1fRuKxzcnUmDZOVSei8LQJFXVJX5tugq5E
WO+re69NKtlXA/31nZYWi4FYYPJYt/PWV06Zu4bfyJxZqkxCiV/rfco28vIhwASI
iuylRiP4r9P26TC78H2UavAMcyn13kLiHPYAXgs6LsMmp9r/ihh2/5aeVXHAAXpw
EhYBUnbdemzXTXEZIPSWR0jEciPZSsquzeH+TiqbZMgLuWgvGSGd/cSSAXSz3CZ1
A2ZL+UjLJcmXWoBQmqIN2MR0HxXYF3XboLNP3KXuYH/FxNg86tJU/wNlvioNBkax
HdJyVAM+MRUmyYz1P74mAfiQA4J4swpzbLqWvmeUh+Qz+NPyDlKGSAdRg9m6XWJS
VPAumiyU+CC8P+ZDR1o91YLM1MyjjPCYa8HL6vgEnnLtgzbZeT9dsg2R+1pD/mx1
/yPbtk0OHLF1Qs6Q3GBUWhuBwMFfKBBQtIfUyo8EACnNcujlrqk0jHM+2U5j05LS
aG1C0/IEEOhMw/7YhG18F5UdQIH9T4Iy6isr+Hsoma0YWtDDWPNFZ0lvn9goSNu0
IFAdmnDF6LPCGah7lzsT6kPadkz1FnIrk8GcgP/9j8UOfOYII8a2v9b8yJOEgUlT
68yYI9XsWiPM7uMrNj+uJeNlfEO1G3fnGydbdufS2ngtZ6Ce6cwtwuh476W6Aljc
NnwIJ9P7vcIDUPQtRc62rV6f2imIJDQs/4BrCDw/QY8RqethZYMXeJo/3Dg7dBqd
i0+RR2x66QJy4kOmnd9l7mDkbBF3mYJazWo4OJzUZD9ClOrV2DKowvkuND9OqA+B
5RXBfQdjK9OqatUfHPasMAMgsYr70P8HrODmXWi0TSuWlzM5IIkc+DTjqbNVodDS
mGrDFZcfRsBh6ZkD/t5F2yg7og3qbKv+u8gAwHmvW3ANQglI34/HuK5yWSDTaTHH
mQzEmtAY8omtdNPQvM/wnJQqqLdkp+6FecBbrs+YkGZ4a+ULU0kCyqHTigJLzit3
VldUVOWZ0KEC/gbRpLH6xX79WefMhQgO+slwpFNpwdYNxDwhVsBFbAGYXUg0dZsF
oquIUHxEsDQ1zdm30NyhdtCF3x3thZ+7PsNEyF7DRjMwZbd7dQkNfrZMnDMdTNJQ
Ry/FHHhZB0CToA1BAPFS0mafCOVTKDnaHyOW3aTslyWT483HYXq5GihPR+JvWb5n
xaGdUG08tXPGcRv9PH1v2GEMuAlYqRx2xR+HWEYtBG4NoBQBCkceSoq5aMX6j6AO
w+wTbZzfba+Utf5sRT2U+aPsFB38pRGGpHPh1erhiEeQjVR7B6Scxi9fZ2xYeIdd
vs4Ltz3Smpib9pMCNj4vIFlNC0H9PthVmtSJjNHbTx4pU33m39NgcrNjwx9jYrC4
waDgYl05ZWJg/SC+qdW7SVN2LBU+Y8Qr37IJDy90mob3xtU4VS/eafZioXcVs0mB
ICB97g2f2x9C5AYtKWtDgzUgrGoPc+peVl2PMrRJVyLsdmOUItID1bdXJ3jKFJz7
hLZMsq8oMF5YznBxIBg4e50XrjjBjpBteFOQCeoe5WyA6TR1cRRLnvRvVcRGnDBe
ZmVU8aEZYoBu+vTznOYYP6pREBMI9dcYviUWWMUq8pvPV4aR+n4kVmn16aWXngYi
G4B9L3uqHxUSuvA3Eq5PWCGw2gkjsvEwPsqrMmMpyoujFMvjSAKfLGr3XKrwQNyk
Z5WUEonYBRi/XLfQ22/JDp6BnHDVnLC3ahPDIreOa/GQZqZAf8WSLGvxF4e8P1ns
NB3nfYrDOGpm62fLP2nWI0LxwrF5mi01aLhxnP7NcVIj6rZf+ziqmHUxiFvOPYtN
Yurx1SH1XtsGA46MpXzGXj8X/TpSClk5WO0xtGp24eqYDW5UHWTEZJT/fhzKKrof
u/M5BFgGSqOF/fuOgTjKOHiEtUtfrg6ftHiqPDM9V6mP8LWOMtFIuds6DYaBou86
WBoOHUc5JH7BiNJ+vanC2KL39G9LSr7A6wgdPvn2g2xXY7O4MIbz4lKnjKjTwZzv
28BLi+9+gxhFmaHvTkBP3s5sEiwIjjjbLpne3c+cKY6jRgbFGzTMZpTRbyIMRG4y
D/cYlm7ld9kRd//65XC2JfowGlGfBS281EzHr3JVjiXmpk7uQwkbU7FPf6ZaC5tx
zuWrJmRkj62FfExuqkn7QnbtixY2XIAQDek5Mzl4bkPzGTR50b0QBJA9lfo1D7Bo
pQWKmmTjROLUh9PtZ8I+NHu0B7zHalUt5zVzp8CE8z3IULwyBB6JFWCAgiwQEsXj
c1td/lRrOH1YtE/dZ3J3QkFnK/P8LxarX58qhD5oQEVH3JD8EYzwFtqOd38XdjhC
e4LNFk02JVvxtWwY6FwTzkwhp621zU7UgacHm7NYmzyoPu4H/10jN5eU3WeRpEkH
fPUVe1C0NUYULrmcBp3fYfoj4lB86RQj66Bw0NazLX0eL7cD/6TXeeN0R5HliwCu
F1jee/ZpdS0MzRe7IIZsTJJxj6OyTrXbszoadRmBjkH6ITjbngOEipNUVWyc6LoV
Ghhe7tGcRg1n+3a1OK86c7QPQvBXkiLl/WkVa6Qi6/2W9ysDNSq8iAqy30ziSWwJ
Mk/QwF84VrKcBN8zSMqxfPySc8T9bn9xw/XeA9Od0RAqV6mrnK8OdT3t5xec41Sv
AK9ZzCF5I9GnuvV+9pQ6dEhQxVLInMaMf8GxOGmnox5+vwYD4VrtutGzFTHSsyPv
rM+Vzx5fex2sDmOgc8p7fIPz4ser2cMzS7E8SfHtXGR7IZzew+DUEcC6V/dVJ/mV
xgckt3LxZGCIf4kSI9WOZiZP+fR4Amx/sZI1uuUANhcNuorLHP2xaeHRqtDRhciX
gJqIHBvzUEzWfVo/UXJmm3h4NcCHAli6V6hO5rMuyyfT3wk/BZtuWen57XGkOmPu
C0Op8L4spbKOzx+6LA7VUSUOfLVByGRnrxVccd8qfzjjgZyzylFBwf7XYqZFFqqq
WizCsYkK+474urbSZBsQLv5ElH29GGrG7jbVG/e+OuACv6QedvNlQcdhl28MgeVc
1MllZi1QgRn8KuZ3S3pZRabJV41iCoE0ztM2R4XUVmiqXKQGbWQcnuLeFwV5pCmC
XRNGusU3rShI8DDvAP4Qhk0bTw884UUR07tp/NSiZGJzBi0lnYhDXqAl1cb7pYU+
2KfyX3ZejVhK8cZ0Yl8cRRQvoLksZjeqdsG6MXBDbKMWJ0OekeT8p26fWbqTiLAc
7xzUooLSgbsRk7b7oDZx9nbMapJ9YIzs8dPxr0WSt277e6YeSb/NGZJwtbaJYJ2X
l12eUwyLUWWZ/o46Oh/HmtDW6KCbuLvGQ+jVdwpSethjpfAbrZG4LEhuv9pgAJyf
tDnizqJKrQOaGm1wLbER3zAUxgKXWOt4NVkr9Lmx1XEwqJyMRmQ7JYNgKuuyilZv
aQR3vlLQK1lXRbH6qBFmNvUlgVPZMS8LiDGMeL1V/KELD303YBSHim5H2k7aa3iW
5UMJu+e3w6zoIkABt70LwSONs6kThxWBgj3O3qL/TsONE7UKSDyKvXPPQXzjgPG4
jJ4r58ijDJh4Up3GXsgJXXfeWqGAstBFy5IZEaYcbCY8gzse3QAjIYAQUGy3Sfhk
FJYc7uSDWfaDkpH+ZANzrBDWmRPgFOpQkytsPaEnXf6qjp4nk975jSDhFmJteTl/
BJ7z1WNlsJF/XSfgGu6eKSaq6GZ0YyK6VihWAHwAC0PNEK2VhynVvF3x29h+M4bz
78HGc6bocFYPZb0D1lAsjFj5gEz/mw7RL/XFLSkfcMtLri5NdOMOFbL5GaFQHt3X
W1b+m/s8q3z347IhD+LSUddQ/ishXEskq5S5W8YIUBHEYyw0qp1Z6sTbg+bCXxmq
o9tDrEoX42inUEuBQ8il8ykALO2XThq7/mLVH7lJ+XWg6s35YzO3KIdRZXzeT1cy
lUKcBmyaH/OFzNsC7+ZJ8Kii01pLJMHPlsBwq/FWTFLIZg3Xag31p3AiKHvOncet
p/ReF7ZqHXcuWV+75hQWaV9k4Vl2Emr9GC/B03qHR6s0j1xtxnkE7mWXR3SMHtgw
ThZ4Z58RTgXVMoT8v8/7xsnZX8ezmFo9Sd1ItmhkSHRwMm3UiGf69ClNGpryCnRS
uttD5GQjdiR8ovC2bYrd3Q/07lhH+4lFO9ca6DO6m+Pyny5oXd36LL3LYhSqimQo
uvTvrN3UhkPpUbmCp4NcoBG9XEVzHJvjApoXlAqCotcCY+hwUYYJOa+2VH5hLEg1
iiRCF3UQjtB6irG8xf/gDQ4fer3xbHFPOPXtXRnRIjb1GYaCF1M47W0bc5NpmNhk
r/qKioEZT6vyJsGx086IoWdvvP55eMXIPMUsX/dT71jZ2wZYXd27ZAhcQCWUbALV
xTu6WoRS3ou2o3CQEBnLuIOjMaHgabmXKTAYlwT1+FueZ91thDMZtD3dISJdtKEA
OTYfW6h5yrbk6ONhfg0fXsjAzY8IPrVK6/Jxd2CqEDhCglh2vOfg/LduwiaPR/6F
bKxAPNYfxcBr3MyPOHSZLil2ZOKTu5Z3INUFE3IIgHez6R2vK3A3rFfIVKpm6DDT
Vq7noSiA7lvzvoSLIkjKWjWvtP1mY7HrsYcXaP//MIz+PIQVBz+PLst1DTMSKRon
MrsK6XGCik9VcdzeHbVclQ0TZ70C3Z83NMHyKYh30OlVFZgBCjNUiv2s0qa/uotV
p+WvdD+1jjDY7LJ9i64hP3PyfELt3hSUERcjOTz9zdlKgejMD17TD+1Q5KJ/FiWC
i7xVxA9zaKFqIqb1lnfRMhRf7iKAcU8wA+UC6Xn5GwLsMmOrhZvHd6GIUptKgy3n
q5MoIMCjPHEXIrhxMLpGPeoa4XDUT0rIfu6sVnYpK9yOIRudA8WovPOJQwSY7ZLw
kMnBplvfAoLGTEphCU67DXvxDwzIumNtnbCLCf7w92IJWrKzhUjINK+JySrZAzMl
mqkMVL/H1G6pevz5zG65BjvhBrju1eyS2VhD5lgcOE/OJeAdqEkW/xr/EEKW+vJt
ELk5Xo6b2Pv8XgSGE6KQL+RD2I9PHh7HKT3rncDppAH+3BDtWccp0tqrJVDQWe0p
keZY0Tr0fKKPUqsVagMGp28MC/juag62nsGL04IHSkXqMd1Y6DuNFfu3T4kabb5l
zXJNcq7tyAM2T6hbVR/2Vzw4uAmu2UuFbe7/RM5bllzZik1tb+6+qsxzzMjSGiyZ
4ooYGmsKuJUlQm16B2AkrfAiVvHH2ol8e5QWUpgTq3YsS6N++oPaXLQWvgd6rZEN
mgOkTjLr6brK8KVCJ5/EuL6FGzEiOzDiHycbcbo6qL/dIMpqTn4r6MhJ53e5s1y+
alDjsk8b5Aq4hyihh0aHU5hiE5lcydQDFPV6pK9zhWUSlpEErAOE3ANDisDfSRNS
o+2f/Kf5QbOH/JvKzEZ6PF666cPbLpnk8c1oij0Ok0aPYgobCflZe4riwRfQ3znt
252WCthF2h8jnlgdS2ACuOHbuqDN6DYyZsOlvt7dCdd2W04qeNoMtfivpVpdVhj2
zUlKPB11fx1txwssNXOGi4gUHMj4wzJ16dCU1/thLX+T7R47RT0GR4ic4Oj7vetd
acf1BNG8gYZ2PE4rgIxkgLWcBAem5hx3XYqVr5OLBN44iRS13ckhGalO0qOPrO2i
QCzVPUmgdYYaknKLOwRov+BKSnCcyb3TUq2alKhSdSGDciP2cLWeDFuPbNSZzz4j
/ChHZFUhOtnIwWigsvoZRvnDkn0rqf+PJ1qTaVkU5qjpLdqYtlKSuQMAaRbQ4ysx
NMWrIkRCECE3GRV3zSd83wH7QZMd6pCFBsQbM0l4KUWHxqDd9jfEXhODuhAd8wOc
fOJkSVGRdnhiFjNVyYVrZz5VErFBa/aMAruDLhiaojNg6jpcupROz9aNeDI3hzbV
e6uluTbKobdxeEAcfJdZ7WQtBqUIKCUWIhXLKY7Zg7dOXoTu1T0kfdko7IZZtxhU
Q2e+icNWRgl9yXkfStJ5lRjZGL7ZJWQJSQqoM2twfFBYR1VuS8YujETBqxxQz+mP
SMHbLoZy7aAdh7gahRs71FF+ueG9UPKkKM1xK044IgVheJ5YyH9pHpUDZ66JFR+F
4koFdN1YWfdxPrTptf7XYp3VV6AttPz9RD2+YU0HtX6xV8YUbZCn41qIa2RvlNyN
GEEKW5vdvpKhjf3ubKj11V14o4SzZMoOuFifrsYzlZ6Rv/lU5fv57n0mDkgAsHmw
1DtQPooXSYwvKXIT2t4+X8Goxjo2MSojSc52rlLMdYUkSUP82OpCpDxW/YVCqS2T
F+CP/noZ8l8mYBBdma1kbU3zugKObw9doBFT/lIWnG0+tWi9awIPauf1TFB6aoy7
i8yze6xFm8G6Rcl2TVG16lvI+RAGokObqjvrJxdxynjJE0shiNhNmT2hBNddX92r
T5mGO/eOeMglkfu3Rg4BYk+bCAPaa9uD4/uY8KdxDRoPqTdD7QRXsrwteVCjzTzB
hZqlqLVUQJSfgRSo6yv/hT/OaDrD1qpkCqHyiBffeKgwsOkRIDe5I3WRlN/MSo9c
J0UFtNhNHlH/8ceuXgCavTQvM4L37tofZ66NRncJExj399no3FPqK6ybFsfUYOt+
+KjVJvOvkmCbsiq6Y1gwcnqIxef8F15DaH1D10I85dIapICbvVKIDdBInBLYRFi9
HUoLS88hZahO55H9sHVbVeW1upGVtxFkJMmKy8OraqT9xlbIXk5E0+zF3aOIGDkP
TPwlEZqFsst+AYCEGIal7/PW3BbE4drNzb4PqWNO+kq192hmAhx6MozU1J2v7M4J
8siHvJ3phB/SqIbbQGE8X08Q6CgoY8JAs+w6SwF69njb+jt7y37YRfVLI9GrN6ao
fJ4xkrkHxgTjlaVRAO7qBN69NOTQb2awxp6bA5E4DEFDRbEuuoyjb8oXDz1v7EWK
07CTy16p0U+SYM7qqZQMLb1cYPVi1uG5yutsSd2QDfX0UhbnGjHXUQt9RZJDoMyd
w+Dy+7iQHUMMFuSLNhu4tu5vPAsQWy7nY78cttaszDLUMKt7D16ebu7cKsO4LYW0
/kSqDlqEFyoLgnU+Fmwg9sH7ST6/PwIGrfIzu/X03iAH+D+XEBAFxTAIXa6NM4+v
pO4atYUVzbyWGIIOIrl1TQjXhUbOeGXYw6SLA+HoHDGY9VxIUHSM84Kl5qgvv3u6
7gj6Ovad3NPyqhU8eVVSMQzcwk8qeCrZn9Re1GkyES6nmJ2aNFh58lkibEhuro+Q
cTs2UC4EVmar/S5Pr03h0v5Fta7sHdfLQ+p8c553TkYvNkDVElg9WLSNeGWrvyYz
yVub+0UXO+uma1Q2lpkBvMADMY2e9psYsPxDJoR2w5HPZH3zhlr2/WDMsPTolhUs
/V2s8naN0HSjn8CiAwlp/b8SGanS0C37wqtJmybkfsipEg2bvUiJd1MlEyyOSip9
/B+E4G/1wzc/sspcQqDjHb3QrTe41/+qPfzAm0M3JjWELOh3pRdgjTDqqrjlfi8n
kdMAnxjfeZCYHYHuNcd9cJcv20z04ICaREto7iuT7f7oFQHvYnp7d8Z76tX9HVtl
xDRFrEzRTnGPU/YZfM9paWixq8A904C1DQVrRc5GZk3GSzkPfw8zeuLKNzW6FlQg
OFgnNEqbn2OXVKj8Cjzu+BG9wrMtudLCkWln0ye4q9wqO+gTVpbUQpblA6zcbOrq
RMouSc2SS/lUM3T16oftKiKnDEfKUoSsHljGjWZxmFq0zWXbBIVWV8/xBbigpGf5
4fx9X7M+0UFNln+873b/GniNkGWUGH3zFkdATdccXJBXifyRmSsdVc3rW9Pib9hx
h2OMvhOcdP/pWafrBJMx9l6pT82f+3YoxnY7PP8ZWaus2byAqNKu86Z3PCC/roxG
EmZGYUWS9+hWYaC9GwUKe42Zpetdk2SwVjrUImTigvbXukyddrwpYLL9yuLlufs5
ZRMBfDmgojLDJzxzhDvTSc0XoMySVVNOjMEJ2S0zfCuE5NDRWpR4l58tYmxuvAxv
S5ncRNL65QlZN1xVtkX1J+TpTHJkYAdHsCagtOkDyX4gn2PEK5XNqMBDzG+H0JbF
KAMZN+8iKjn5FBZtJ9m8HCc5GYVYNmE+UM8i+GaSt+puksiGWMQsvJHwHH1m0Fe4
vBnJFVSxL7r/XKprXvMXL+7ROBC50R7NtBiFM4SdDPStKk0tTvPDTdlszXKg8E72
T8Ane/wwZH2zkY9QOr2Rd4JDh/yDbeUbNA6CXPcbbEYWR6EppVwSZSmdI7L0jqV5
SdKZRMlN8O1TYitMSyndEQkJs6ec2beugGz5o739riBKVLpdNYf0Gb2QDMJ2+E1i
v/aEl9KurubaPJ6MS/RUxhhwtteM9Tsp9LTCyycTcRkQlMQyFlJKrv5r3K591LvB
Vv0/y04zk/53/vtTVe8GiyVtwyZzMqsEMf2jpHL95B2ENQ1Tad39Xc29xepUvn+3
TJLrcDxXE1lK884bnrKNm2gnY2YmIe8EAZ+B6FAOHFEr+16AxkIxi0MEjfD4pobi
9bW4XggkaVtG+7Irxp12tEelKjRZbVzWXktU4SfF6PKfB8ocdRdIyN27twlbpL9S
//0TDmBN4wy4TAPFVebGIZMMlDRwLRw8OduDwR30I5ohvMQEErB73OcBEqr6hWuY
a2zYUgajfyBDUPMJVaioD5EEJGdByrwYTenU8GBT3i2FN30sBLIuBVcTm3/2i4Wf
G3kEgAmbbvJN2FRiFmE4XDjpIpBjbZsIJtgRr7pbGWbBRyy06aNCFiNy3iz3RAAj
fFqs6sZZGJfThC62tRSJt6oFfhBlTuhVpt7XyMA5iyrffB6BC4ZI8Yq8kICyr8T0
3RAtk9SdN/dMNTxNURF4YADXJjYKk9RiPINmoDGi5/uLjtAVBOQennZKgqrHkckW
iH/80OsnR+f/osd7w+YrBzS5KJUGHMDygSeNOGNrIVWQReIM4qWpPM0UWsRp16Gl
gP5zPrl944Mp/hqEys0XZjdQ2mGvuqen+5bmwx1bKcEu/auSOiqiXuh781lY+7+O
7VTtmPvz+goH1ZCKSxnQMff3ENgKjhx2J/yYVoKqVZ8R5TtS2/o5Wl1AbD0bUc9T
oeKn7ndIBE7COlGy4pWgQQXxVf7Rl5sYE/N6h0D8YmeLLYkZbF4DRggaNQhh/Rox
txweOKZvMV+PCfCICsHAQJZbs0CHrUrsDGUURVZDtJ5f0D2CzQrzkPGOR1RTYx9v
IqC49QkvCNXZ4Vbk0Vf1IObtU/0BHRr98er+M8ZXoH0+QYiN+q6h0eqeDYvcXEXK
LZkoN1f0QHEfd7wqxlMY2bEuJzA3x5bYietjqxjcUdT1PKns7pYnLR0xpFPAxetu
KsINyx+Ms7mn5LZK/v5RvV2xYScqDt04cbfW+zSKdfw1HYC8PT4Cvd+XjqpJP3gu
SeyiUy5SOAD44+DP7u+j0/PoWQRV31PBzLK9Gb0mkDUJwGwrgunqE6G1KpEL1vd1
tWAggC3+dpD9oy5UJNfcyFl3vbGypByHXKk7pipII4+eliwvS4I4jCHQ7F0AaHK7
X3qC6jTd5Ew01ddH/OvDc9ReuQIFlmbGrGThl6SdnZByJEt1Ig+rUtkOpaWF4BeB
mgso+zEGkJdH0pazDePDphyeTFrzDTwEC2N/zhjl0Ey9TLpRxo8Yhm/ULZfZnUMe
XuXz/wiOBcsLbWVqMGiOG0SwC8c0og5EsmIWO1cNEwnLPFO1ccB9NMXVk8lrsOxa
dn6F9eUVFFpsQjqgv1bPzilJAW2HzAPnTUvqubZKi0bYpkPvoY9mEYzhFbuK+I1K
uV8gF4fgHw4skrTerxz6V8YyWB1oA+TLy4ZV6xKhqhq7XzTjB285o6d0RckSyThF
D6VvbDARxU5cyYun4qFRJKmj1Ff+CJszzF2ZPYsIuuLaDHIyHnMrYnILtYPUx2KN
p+5O0fZZSXLe430OpJZKYujH9l3qIfEg1Hw3uQNCItkB2CK1xjez+xhx7vNp56GA
W0TzBsVmW/wn4BwjLCxEzjnGY+gZ/4YVrO3L5NQxOGTukqO4N+n9fZOZsfdabWJg
SzYJIxVuYVr7mScNk9X50WRvhcMsLo5o3fBY5h5pC8tbfwpmGZsN6EDEtgRZ2cNr
uTw/aD1xZrg5rSqPP85LSVHqkaHJ7d7lmKaj6z2cPptMCfhbCkRh2YlL+9WYdSvy
IpgpO0/p2HaByEjWrVkZtMoe7WmKpF4QnFlM5qvPw6Kjvws+am+VhwKj/nsb3BGd
fRilGJ3Xcvfn9ND0YIUTOHUocbW8rA9EiZ66pcE66uYOk6kMGjdnEH8J2l9d7FDQ
gYJXACfuKCPgBTZ6TnqPmXEo3oG9dE6mn03uMGLrdfHxJoCAJtdmFK9Hxr+qB1D7
nL1UC1MRCoXgEwjg23sWpUJGfH5JGQVE7dOJkkEwqfNMjW4tpifajfIBkpRZAM2C
vnJUX/6+0ZG2F/8LwtSbJ9gvUM9TXzYYwYI1vqQggvNZi2OmoWU8TPPE4+oV+hVL
S0niPcT8NiHbuipQqFZqddAseYw9CuYecoUuuYWVaf6xgewbJ3EJoYIVth1fgu1G
v+tURTZjUK7fM0OA/uHa8102EDTVz44/rlz4n6gABH1mOwJYO6Ux43HaL8cTRWiB
hD9EW2tWK4i2qb8bpOdzSpAfvZZtHehMF4aVE4HscxzjalyK36f4jJPGk1uzCFT2
HnNYIw/LlZ1q8qyTS6Fizwi594v39n8EH3V6JLfbfUl7l9LzULwpgLIKidArwfIr
G+li/PDyPCoZ72AJkEcTJoyovJhmwEoe4HR0kGEZ+ZICVoG9TCw43ktCkLdVf/5C
3+vM7wtYWRd0uXMmck/7/TkiPkmn0fq7UuXJdLE15hq/DU4GIsq7Bg5xiZfpGvn4
4gLOY2ZZexJCLr4aEoGpH3+YeqisB1d8yIMrg+PlR2iJ1FwfVV4uxk4qfASm9isK
7T6T4xBTGP1nnkgtmyL5ruxQ1uXNFlVX1rvVJwA7fQRZAmh9HE2epxSCiOHOLdPp
D8JDUNY+ezR18v7Lkga1DrGAIL8EwUrY5jv1P0q+tYL8XT8C9qFto1Q5HQj/3nZR
0FBJ25VFSUSRpLeAG4cWd8B1qboiwdMIb6k9tWf+O8YqVu5Ay/Yj9HAnJlJfVc/7
9qvdEU/n0YLGRhFqjHXWNFZ5YsbHvS56wvk3Qki4bOdYynNBmkoQVQ5+ovWtFP9H
PXyUYNFz8wS4eRat4iu5omqoe/C544gV/Po8+q3OKrgMfIjpiFj7OzK5cPn76AMj
Ql1PrbTN05XATZ3u/1dN+RzOT6WFuc07BT/dj1KgA/zZ1pdeT/Cj3mmsR5SE7OEV
cxtHZZsyXzN2Dwq8aPNkyHyiIS8eQmOa1Mk+q7weG190ZHnGEFYBMLU/gVhP1uCq
kSqwCk77I6JJJtunNEVp5EINkSXrS8cavBsXPCsMqtDppk8arKo6CK/LnplWWULV
LDKUz+A30PHNvpJOp+PhlXsLjbYuy7wy26MH+IvN/G0rSUqoWF5fa+7QLl58VnhO
xV/lKJcnM/H+uMUa8Gkl/8nIAs4OS1yroEJIPR0p8btUU1GpfUdMl9mXSFp3V54w
tJP9FPLHZjwVbEtbTU9ePSu8fkoBYC9vUO7ck5npJuTo5Dw6NEN4+JqpXq3eWWVF
RXUrEllRpVmC33rsInu6fyY7+ccL8DRZBmnNJ2wYJERE01HsGJ5Sw9ve+f0puPEW
p0NTVOhlNWnvSeo95dbJm0dqtfq1zrMK0i6bhsMTEWxBNRM+mMKhsXX8xvoHIBPS
mkMr7DpLEd/gQVM2XECreQGFcaaCmqY3KJZfSWB1DpI0t6f1mVHqJBv8UhginziH
qyhquWiv6sn98WFYIfzfblZ6bhjnsZygOD3EGPxIb+1w/vQpEjOfW6BNvIuStUW8
ajNIB73i802sJP500cpYLE4CafwPZlTtKmQeJjldwPVUJGtbsR7rHGMYc1FQu7yO
DUbb12peY21Gd0nvT8SYcrcxawE/p7sWuzdk8D8tWSqblVHk6GGSlm+NNjMhd6kH
lzHmfDkuJv9Pz1GB5vcI5jeY1S5/bCkKgOHmXPXrbTc1WA+VRb4TJdJicvWG7nH8
S/3Xmxx5zyacvNb3bx8+7Y9/vQce7pwZUnepWVMQ3o8j/YOuyhFqX7mAnMTYSgFy
3bYlfFPc2oW/BZ6jOKk5Qs0BW/ZdQuOLlqCq5t+neo6G+/Z8ISkVqFREQfFiYW2I
8w5oWaHeRIuWebneSNqYpVmhJWbk9zh02HrtZ1k84zT2ZOGgFuTKGIQ46kBXEYKe
kiAvlfB1SSlC5gpgsKd/ITqTdZitHtpE44UsqzTWrQ7dS0WCtrHJ83yrd/SjuQZm
beXX9PN7zWI+YsnaEVyqn96esA5EO6iljj7zEGivE//kdKc3SQLNATcxi5rxlKrz
ubdh8zhNZ9iRXHfJdempvcJb6N2LTLFpjOLgCDIx3iW465d9UQSPOxgDxMaixs1N
XfO7ZbZE25fNmY6S8dCIrCV4V1WGv2v3v9W9OPobBWWZyO5t8gXndPkDb1sG3mpu
REgI5b/+MPrNdxM/B1cXEWZEXNCcGHPKP49k4zjd4ATW1YiLgXZtUb3c5hQ4A3Q1
7x4s/WlFupxfGeKURPc7fVJdE0716A7gDM31CdEeD8J6rUEqT5NrBdq1y8Nziqof
9rAMxft8jB0MCCH88bg8iuTO2X6E0k+bB68MCnYzv7u0kN1uBtSmJrh1f7oIBULY
MqMyOaCKTf0RnuiqfyvyBu1UvNanCw4jI2Sw7Kghn2aPggrWOaS8dducP4S6tjZ8
Dz5ovSSbXtNvSY9PNWiYnOZ8NmQ6YGLLU+I5NlFhPJY3HXKIypme1TvI/h8LoC1d
nLmhGXl/vQzjGQu9/f1ed4hbMlt0JuPOA5kc031ahttdub6AK2fy5a776eal3Suc
p6qHrzxXrWaLLRQfAtCQ3X8xZ5hzWDtT0C7I72R1cAyVV+jRACVJ2MfCbGvdV1lL
F4kCv0sHDmySRMo3217K3SvZlmbu7pjvp3m9AKLWRR/dNu9AW4gYD2eqnCr97EQZ
h2+bwTqyAuHQ0afydeao3YPLYoxrMyBI5q1663/H0utyp0jQxBpq7y33P5OqvqxM
FLMXi4Utz1Fh9PZxY53FbI5JfUqDAsyd4EFWwxf3JiAApzBKtGNR6x2PQQk0hfDI
lbvVl5+9+0AZ7ouqvJAuEYYT/hymFQyuCTlKiHmUYFG0kRlgeXaweuhDwXSdgBeM
liy7pAkwJEHKArjUEZCvAPqCX/KqFxI6F6p5tATPdyPEC1Ml1+94baf1OC/uBC1Y
XLWsxlGJ7h64fP9lBEgrIXRulNsySfJ0KpIMMbjHys0lZMn6/AiGQikNIsjZHpm7
xAlb/ULrr9hClCSC6wGtg1wY/JB5ae0MJC1aMZdFrDpDVGSTCh1uC9hezhWsIkGX
P+/Y9EcfNlkvAkOvd3kNN8Bq13kIgfTXQB+hnQaY+rXYc1gZQdNnk7d8vtLZDZfl
qM8YbLC1EWND9gmzYFDxtwZDwwhbyfIRulcr8pzwwXjxwcvou89Enlip1XBau8gN
q8EWuB4S+6anGQRHehD3VyeTfvPk+3AsdPrUrlJ3XFxz2J1YsNAWtWnacmj2UIZR
JA4jhFF6NfgXo+6m5KDjVjgrOL5xwg22dAWjWMo6h3mQqzf3QFGd1Jdv8HaXl5de
gL2ZiV52WDDtIXirDIAQA1ZKDu24okR1bYF+f2H99SyZT9tQxWxX0dQdkdOAAVfn
vpLx8qUsFsu1tKI4nDPIg/Gojh3iXnmivuLK+j9z3G1Zyi+vu5wCRqhX+gF4umTL
21Yb9ir6NeIEEZSn13zqjUEk92NPUFG9NFAI5EWa+4pUbLZ2ChxcsNmmG0j0pdwr
vbP+lXpGIqgc2pu9nv/N7FnRoNbJOdNWgm85DWT18JkHZjfFCYBCtLmQEc4iTO7r
Em74yO44XVvlDINb2nYqLoqwKSbFdeVLRhtKWBUYzkPXpEo7a5vaziauNJh6awYA
akrOwuGSgCr2yuB+XNdtbl6QRnk1Ie3NRPWnGaZC1fmkt6WscXWCfym/EaAoaYGZ
/gFbLIafxK6gxGctS2Nny18YmX1KRwA03ZffRHtf4+1v3kCuEM8fI5cdMPk6x/C0
3j1U2HmWG3GrEZeBA2RV0jvTKgo6kYOLmObZ7hlcbPiI2uGp4T+fIfbmRqZQR4cO
fyCnRut6ff8zBy7azGC2rqVj+EkRfBgKmQ5GcyMWxOJ9qr0zZkCI8wecfo4QIwVP
HxzDVk9mnTVDDaoQL0tNyiRVms0xxO+noR6ZTxC7nYBaG2nEo49ck1RAB+1EFrGB
v0VOpHh32mbZZMzv6yYOp1a5FnJjBjznI+DZmOswlwnDnQ5fPe9PBC4ImcnXFEuu
kW97VAtld9nayLJWPxi3PjrkuwCMpjmIPoG1k648zMxSqX7EjH/8fFI35ewe0ykI
WN8787szkTimoji7OAER/IjZkAWkRV4yTq934+HZt45lauyhW46aotFGJyGiebqO
XGJUTF3q7NzuRwCGrQuWulaUNGm381ccAN2cAYRQRCIWdtobh5UlBpSvr0xXGjXr
twvhXPdPh4Dy0QxDztCCb3+zfvw42N8auvVgmt2SF3xut3cXATW3pzBBI0/VKtp4
fiqQPdcAtKQogf16CgfNpvo2bB1q8W7a7nY8PiDJo4DfuK94E4dDLJGj0di4oy5k
QaqxzesQlfXxiRQZaCxDrMe4qKtFG+Q6pATShpjIb39uB85HBEJXVYbIo7buTnXv
+6wjmq94zsYdVn6hCzM3v76w7BBHQxx162JXiY9LMx10WynDKmqkzg2O1tW6Eeo7
HypNFCnHEly5lzn4Ao47Q0nr9v5qj5rX3x2E7pC6I0X62cY0+ZPnmFXj2FxOMMnf
OTXLyaxUDybj6k80/RpB5UAFg0xy4F0b1h5+Ixpk0gqzTJLcbzOsBVvR7Vkno/c9
lqe0PMxaqLAXSn9CEll5PXyXISfistB+wIm4EbTRi/cOnlQbKndzs2n+zEc0DE/E
7jPaiOG3b7WRFmC6KMv+5yfWBml0Aq5lHsxqw0mgF9eac6bLvX+L5ic8Z/Okrdj7
N7SmWJ8ctx/9MdEEmN1Ud8U9sRzo6NlF6QeeNEOkAoA/psopMWBLvAg7tsvcQSTW
7iqQVOpFEhvrChUVsATHbR+t624Q2rwyCXMx1VYqXm8Boyq/HfMCgwjrgFdlHg/k
atMIlWLmbHb99J1YOz0sCLgLZqf1j3wTSFpRFvWwYJZqErbeq5lrEMeu+PEItZ4b
rsmEo17l+01RAkJWSBBkbAaY81JVTCmET7pruO6FbLM+CR4kTMa8gcFDgSXC7fXf
fndHykfn4HVjJJ1qfq90hp7t6FC9WjeaQDlmiyjGcsOWihGkWeUYIznSE/ct0iBW
wYWzdErlKdSrbDB73k31bE2nlIYxqWLCSF5Vs9/LxVtwfoA4aCy7t6SfPk2xxg95
pwNyI7AMsGAiYSIQa6oSvjrIGEyJSad4BbMwE2HoF31BDKFRBWGFIr5OY4xxoQ6H
jpWNTJeCAnsqUeLXPVRkN9T5+BQlygVVaw3lAed8ZRT5nVwVofjRMGvf6pBVst3n
IpEJSqJUKbgbmyXQfFJi/5OAGJY20IAXenhfK+bnopdjeM/dogFx3+XHFQUl6kZQ
KegskhcOi2mfpSKRDMi2Hcz/lFVNA5OYbj/JYsWEevaNJdBUMS6H86hM802s5NeO
dwDJph//hhno4Neh9NLGYLrTavVHLp5aDKU50GH9SvIHIEuF/9f9XG9QxrKCrg3s
gT0KUcUxf32YQp73rd5s+U2cTMb+3+JHY7lJuYH1VxFoDddNe1AjNYPmvSBhgbVD
gk3flU3ZOoS8b4CXUKtNRDdGK6GWCkBhWmvYnoFFj30PJeC4fX33xUDteCmKUDAp
Y6dBW6S/yycBYawMS7jLo9jIiGsZE28k0KsrSCX4VO+zH4fjYKPKxmeo1mK/DIFD
0iY4SCvLcAobR9+1rGN1zPGUkBep211egXRSQXYRYPwbC7/28SgI0Cuw4/CjGRiX
dYifCGZP+f1kcCzG+4nFTEhUeULzViSbYoDzZvqofYtxSW+Q8JyO7H6ibDzsJt15
rspPVl0tAVrEtxAHpS3k7W0w+nojFJ4NW1gJoF1zVzr32D4DBpBHfhxAffH56zF3
kHsH+rYNy8SQFKRXp2rPXDZu8sjZLm6pb/mtAAJ4agLemnNxbZ06c3GIAscNPqs2
CRJdVsR+dv54zogZMHZUrSpaUxgueMGaXla4oTOTon+OJD0e8BajKL1DB5URaX9O
A3yuPiCrugQbZYcJFLO/X3ejTptG/Jxp8Va7vuZHEnGZxzHppGmYqGnXlP2JLz1b
zkkoGBq85h2HjJOK+pJgSc0QQdvM7ua9PuNQ3BM320irqBvu8kHlvr6Qh3ksyEV3
LAkdj1SwkrKoOyauSSdwBXONXOqGrbKxFKAeUV9a8I18sSiRhEJ6RGt6UvhCDWaC
MNpyrPGPecEFLtK8ReOs+B+Tbwvfo5eWI0NvQew7lAaRQdDIK7c5aeyW6RaPGt0H
S5wk728tYUjnWj09+/KwruElR/+bNOvJ8zdKdGVTn0jGDOIPDx0OlI9gTQCYA7IY
JFW15er2n9fjvSIhT62HJ+gp2rpDDbIOu9QaOHm2uuQ44I/PTuZCpPvDVu8XqTlF
PuUjIhWnIXu6fIAbfGRvnWpF2KsRbWQAd3NNwKKstTs+AX2to8tE9TA57uSu5OzJ
uy3xwOdGJO1nMOcCQ6y+95yb0VHSwIRUVXdiOerEBBqC/Cdjih+cAZGsoGWT+9gL
txJNXqykCeA/VIxY6De7ltm5GitMoDT0l28EXPvKa2HCpm61G+FwtrhVf0ku0cSY
FhRg5WUXbJwr6PCjZsMC07udI5EawtH+CZZqDywg+zVtPMq9lEEzJOn8InOZ8FAJ
OAk4sL6EMQ1rTqtn8BBGiOO5TseDxFHPlOjFbLruEn4mEsyoH11oxFDnkHjT7atq
+lXqfEfX+6z5r+WUZgopEkIquQYcF8Emj3t82lgnTF0GcvNbAt712a8lW1X1+Wtl
GcOGC/+AbvGwGymSrh9tseXt7Wuvi2+s9l7V64obpuerE5ktZgHFSjTf75CBdrv/
Zlwk+dNc9BJCyRbuJVfeIwAVdLH+EsYP/IIseILwletciNj8eTsbXHMWKl55t4Pc
8J339dZmwNlq8ro05zTbJVujJ2Fq0S1AwfLHw7HJ0/HSYhP7k+emrg5QJbfpCjmV
GDk/k21Tg6o41uWNVolXUfzptIBX5ZkIXjFtuLSCyQqt/dxDP56WGn38ALgimRdz
5shi6z+FkX0kZPyiUnVoV//VgbENDha4bvS5WkZlE/cDYMcMillqTV+a9uHv9lUv
Wxx8JkW3GGIhLyPLbgfcOuOgCKWwpUV3xEcDp8XYF9iY3W8EDeFFPWWswJMyVqjd
SMKAkcR8mi8d6ToW3EHHmH2bHrMJIOcBrM2D0oollpWHeOjWCCGDmriONAoeWs1e
xLKe6S4OFCBzT7XdKbEAEwlvJ+ES+8frRWV78Ax3eZSstvQ5G/olVnf+6lLcNsv3
Gpf4NfcXsqDYcPCspYBjzlJG1xXgw8Qx57VEqR23MPjv0sWaKS7BR2cbkFerrgiv
MhtWPfCowgJ9KdEPj/pGhP4DZ4gTzHTaIJ9zEHztiq2RmXg7odgt0DbuzWVLScLO
TYNYymAXCh4oYbVLLa1vIA4uhsZUSQ+ScPcENpaJr6lQ6BJW36WFLyjmt1Iz8RNX
kIIfjxeWu9OejUSOpVfIjtQjeMJ9nPCxDZ2IZTbUpBmX/p+JwITtG322VhF7b1sB
zbO4M2vgObSes68OtXJik2x1uHPG0vLQgYiXPEA+DiGRm7nnR+1zCkgujyq6EIC5
JckxalzDuUx+xAjbrd/eLZbHeNsHPcpo7ztGmIkJN4YcNb6p425PSkOW3bqPloWM
P77dBGFkNh25aVx6DwFQoVBlQGl8v44KAHbaO8yukMpTLUQOrNq447pRmeUr1pB0
TSi6k2Wx/Wfbpt3Anf+uFvIyRFw2ayN22dXRA+fGoTLL9YXMMQlkPvUSYZNafxA3
MOWZ1XHV3fuJQ3EsI0fBH2KsTTt7twWsC0hCIcPumMwqBKXYsdGqfxrosPFcBYf5
5wE0eQ6VXJEHH/ZBfWOcu5G0WWRGrE7xuNtYbbtEJIti6cTKtg8dpHKLpSGwN34G
pEqfpEJxT+hLEos/5cU/CQOxFwU22JuoAhRM+K44KutYAm5GysnyScnekxrw6pJk
zw7G4Ewmc4c0ga4gPxgQncpEC4hjfKLI2Il8M6Fcp6zPG/LVKn9sPxv8+izplXIX
nz99mW6z/DUOooQQyBbQxJWcQpgSlsTUf4wBiM26MGsaEKuSwXpZV0RaKDz445SA
QapsAnm/Jih4XZxscyNVk7LYJfYKM04LBcm4o9D2nslvu7BoGxJ0bbQ9KTpOQYiR
WD4YhDGyQI6ksY9vd3rM7z2NgKFOPhzDI35Lf/+QqfHAv3E+xwwAFt8e1ATXwTBD
pYZJ8eyYkCsukEKHF2SI7H1i4Hr75ryRgrnZssCSg/DOeynTpGM/XOmUdk3HSWwo
DsYJGekMsuCjcThcAtxiUOajAeY4MutlvL2UIGWHQA7IvwJGaXLvIPm14QYqkc47
CbRV3qpsB+Hcln1JCuV1eGHnB3rNLTsHWFo9SWWXU9i5BO3wb0gl0BFjhkyEpGmM
utdTzfc5EyoxEK3NRjHOroy2p1UBfOu0AxGBELQlhRNbam6YAhV4SOoBJfkoA4YD
/EPU0mVxZU0fxxOZF7f/V2qEPtoLfpZ8PivH+P9TpNNIMRwjLP4DoCeYrG6X5eee
eNSspJSMNJrCVTcoFtwJrb0VOr8ROHGhEjbBAO92WdeDU9/Izbq57NfDjSYUhNUZ
56HkyT+K+XhzSCbD9tsb2PuxBg6xBWo7LComQVkR1NJG3GCyauSOwDOTgQcx8IfT
g8kqSX93yvehoGtF019vRSv5ea2TOP3egsv9gLXWypmOSa2oG//rYFOZZ9XyTYOp
es57RqIl3zu2m5r1YjtXNihfBu2iYBBwAo5uzZ413d9Z3ew9lJTiLnQ0EZheXQh0
amIVktH2937ZpLdhNV34UhoD8lvhQMTQelbzA3akpEWEQDeWyuU3mUyavlaUtpZt
q8yJCkOUuTS3hahl2wSyMap2zZ85rrtB8/zd/i1I+AdNHnw49YMnLXraAEstPgFA
IJM3SwrSjoHAWxYEiKVTK2PZqz3q4Bm2OKxvE+Jb5UIKyNFbpGuC7w+up3QM45Nr
xwwLEiWs0jlcDUWWx47r/poqCxfRWJLRyVBHXq1Y9X4pcL3P4qFOiaeZfEm/IrAW
CFFsqoyuFpvsowwDZTcb6c0/lstK3kPyPmTdMCDBi1YhO8I7YNb22fioPmp9tXjQ
1IlN2S0UGJLWzW4H7yom1ZUaxIJibrDeqzjGLrpYHT76sLxCED56tgQBHXljRL+b
Zw/7yCK/wLxWu3LWC/YZcxUfeGD/6zXZ/VZT6l+F/EOHEFxouBfKuuPo9hBusBV7
+XXmT5u2Xq4jrMSOrWjDdt6xZzEWpiTYi7FVmrb+EBfD/h0ekoKo/U20S2pznDQ0
bGj5xuCupsx/GS9xzc8gpHuLM8LTBUbP7nQfcw88Ehpkp6IMP77WW1Y5zRwQO/HV
XKtjmMXYMnxLqCB1wWBD7VO/PWUm3W07EFvS/dZ++ckGUpt99xMLFsO4k4NTYu+6
BdrbBqlf6RFC1fqqXUx4DeM6q+XJzRWxSnoqnZ+MXiAf/dxZSoQX/h8i6P8Umptd
nwqz1c6HNDMF7DoiMO1osjdDtF53kvFLBvUMjW26pupC5vJ04rEbpbfjSJYkq3Tc
VS55ebYhbkhyMKcI4oLbmBZb9KwArNfBjsA/Yv9Qmor2O8xJFaa9ksu6tg21+di7
i9lpD1KggZ3UnVrnJtiUjAZl3uAV3GnC+XZ9MrDwvrqdPLVb6GORyink6w5UPzl1
lGvJiClxfaC9HTxSSd/1wde22Ib3w+X0DozQawPEfZJ3pDSi5of+X/6f6oLS0ITq
6t07qG5ObgF/KMAAOEttOsEOQozQFsTILU+YgOChcRDdXttmelzE2WgszxJnePGz
M3uCiQi49zJ+O160/oYt092dTe8AX+njiog3n5gJDkIDSIAHBpBKhwwgGmN0rVm6
vbWvAL6DKN+xRhSA+bE1SvKzNmeOi+EqHtXbf0p4eio/sEr4cI0zPSuVDz2PabrS
lF2EXgIzURPSCm3D6APSRh2wFfEDvQYuJ7gpZpyFjvunWcNuUbBMECQtADiubfTW
X8P2tkgBS2wWrMpAYadOwhRxkBpdofA6OAi/+F6E+FN1PUb4lr1+aoSbs7T3Bl3t
5Px2GE+8qze1TeaXld+rb2/0/cIt02UTRsqVRrw+oVpmeu8SiAbnzUIIwexwNKqQ
FBfFSujNUHcD8MN7uMAkSJEVcCKRJoXlpLiFzdtHq9QGFJVLi7YCkyOkpilAym0k
B3qFPeBwkFaKy0inLAyWbrDq6Ybwk+zdc2HC0VvU7u90YmTOP2hQkKEqjqNRlkrj
8old+TbhuRnA4TZz86+3ciVM1KneZLZ0qB8s4rzJTsi0f4JvrSz0urAxJaot0RTE
sgOKYmaz4tX1CLAmy8ezJ0DdnpB75dXAAwPbP5PbLo7C5KsWY6w32nJi3LHB48yL
ZKviWXzA45eBQZP44NH1gB5hva9Zz1MIOBy93PjoN4aOxl2LXJ5CS4Cbonj19VPu
dyQtlxXPX/HChZx6mS+IJLPcOJnTx/DLSeqVQ9t6tb1KalgE2UzB3+sQzgqy10jr
SIw2L9NJO1QI7HM9/xwHZoSuiHfpe88GM46JE5oOY1mCDuVvZb8aInBEDIW0UW0e
Av4W94qQTmhAr/LwUCazvli9Ug+4Bi41+Q5yytEm8Z/wUq2hpqyep4F1ZaIZ343Y
9tUwiJ9lRjarnuPhyvspzjCs+gmvIBB2CR1rvsBenosXUjU1prYtEd0igvkrZPww
J6eDlsC+WIEqBvT6m1rMZz3h6qg6hRPFyGm3Wm0mYtW0ZCIvuvdhc7VoOapTfSlz
AYo8MyjaUZcpkSh+2OpVP+HvKnTH4hNAHxhbXzAawAK/aA7pojA8Fw0g9oHsuPFx
hkqYmffaPHshQ/Co6/rjznVpXAl2JQ/fX3K5S1HQ7pVrf9WFzFfdF7giGgCv/iXD
ycFLNUnz+Bv4WKofNNuyJxFi38AYncKkYhMUUFffR1B2glV4ZFI4YVp2oX24wdIp
QbuIeVtISAFYXvv6T11IWSHvmiDmMlt4rSdvTc90oGydr3wgpW2LjWveB+cYdHDk
szZfx99lxQqmaLjhwOBVGrSgFmTif+2q9tCrOj2vKmebul50qE9FcL+udH+63OJJ
EnqFnzbGeaxRsGzXhbP9IyUmh5SdxBeZTz7hUEaqptXVbY/WErbf4Y/cr2mPPlDt
/73HQhCBPOpzdX89sEIYBX6/88CDZx3xRpFndnSAgjbYWhlWhznQJio2xDjJrUCV
9QFlxZiN56b3dmis6wFFGu1Up7Zrk1SY9Nts7kdZh98SdzLQvGWoe1zrg42k1zPm
PHs/HoT/Weua5kGItSDbxhi/Dtr6gzQ7QNnucy83fJW6xcZ5ksXanBhpudyTyDUb
FKWSysV90MN7+h3i926e8/jnLCLRZk9YJPCg0nnpPP81breUzZcLQQOhxQqV7Zih
2xoHWYPoLfWQVEKY8aYKtuC2dXMMf8rqb0SDzZE10fDu3o31lRrblT3RcOkkvXT6
+7qbzIgbyYW7Zb4XWjtFheiWKF4RyHtCy2g5WdDzV1alFbaQgdvDxHjubx1KqdkM
p/k0GHO03Qfa8v2k3QcOfKcw3NAboDB3JbbfJ/BbjBKJx5TcgNKdAGbHUMLftPlh
2GxFQ5t/ADoKXQx5iGk/cxSgj1KD1ppGJN1TTEQEvOpM2H856scFj2c1/AWYIelQ
DhDHRjSdmfdNYrsj8KoEk6p+7z+Mo2452cpT8u/D0hMeliuLmCF+648fYINoc5PO
rhZOgebrj+GLrOLAe9N27Dv/tHHPt5gfuPV+71slxHgEwYKb0Qlcwc+58m1FSPBS
6LDag4q/wJVPHVJ0auVZyzlmxVBD4B9t2FvwK93ESNFv64Vkz2y1K2u/k/Ev0kY8
LfqnexKovu19ifR1n//Im3Mzg+KJ42m38fDpifMwyVCwdOtjFvjjRG9xuIGw8DY9
0puf1WHCgqSe+MzJ20dEhVel6b/7eUkGKuk/u1AkENPW5kQTv7EpwEh0SdKikIZr
thcsWqRWHD267zP8dWdyuUMUpInmULoQXNO5aw/xkhO78AZvboCYzkS2KEz492R4
KoyP2R1/rO6HWoXrRZ+CL2kpb3W8zqOUJGN5s0+wbfm7r0JkGNwRTQyWi3oLKPRS
z6BeP0dEmq3gfJxoKsKpkaZ5+aWWvGAmaRUi2BnoMZsNTEUKr06wpLlDFyTL544g
ZaPW7JLebTjQjiPe4d8YfxnyT9lVRYMRaKroLgsHl+g4Dl9vyZuYelnPx2AeCxED
sSgLAAozqlyltnG8vysoZKIPWpelsPygoSYMgUwKUk9hZMxwGKzI3iWVn1LLgfVd
gukSjUFfBCBseLQLD8i2j4K772Zk9YR24O2eCfeTMtDWk6ytFd8P58N9F84SZ8W1
xKfCEUXKsSZfjOaXg+ffNvJetulmPbanSGvT8FXE3OeJ+rhD9sMr8mxsXesG8h0j
wNey+WxTAK7bVyr2/nDlvKBmp+jUn7m3Pcrj1tqnDs8WC/cDiI8Liyr7B1NDAYF1
pUR1x6psZeNaWNzReKW7XsyTeL0HR8sI5Mb2nSMLNoacO0BDr37+L02NiIzZLwgv
nTXlnO1Xpd+U7HuV6vo0P9NAokil42pWxd7SEQMKqlZJqFgatJPe/1pGB3yZf4+a
q23NU/S+l8/XNxjk1/Ysy2qc5xhcOY1WBtpt4pQ1W68p79107HIeAl5JXMD8vYwO
tBuE/YWqko7fuccJYwKq/75f0v0/Tu/mLxSVzA2mQbsDlhnje8e/KkgJaLW+SMO+
BgrHQH0x5E9KMptHRegthNysjEsZzIjmwLm1MIzpnw8pJy6HgD9ouFWVoYBcNBEK
YLoOo/nDEm6jj79KGL+KTgi0BLTGwhkWbkWrNXlodoBeluMj5M1JgTzraqw2Cr+F
ywEmnaL5Q5RzJaaajh3udgdBw/Kb9hyhnZ79WLawEXPvhD66+QZt8cynPQICysuQ
XNJWOlwsiB+FIk9XY5T/KINRT+jIeIjzVO3xkM9aOVT7EupKgfeI2pNRB91hpNEo
AvdgkkRlgE6DIWJCgZWOrvm6vwWOgLrtVfNHWFAU34Y0I9XVPygJumeJh/cJBLTQ
+xt+iwqJ27Ux7jghUcX77WFSYK1VIhnWWLkP+sbkLHuv+Y19ZKd3ZUG3ILhBFFo0
aqdiCAPsMQaV8e9z5pR95UwnKON7RvMDcVhH4tXvcPY/yiUnmt94bS4MIGC/UFPn
B0uQBuIjkkVk0/0mIZnWTzJ1FKbNRtuld9eTeE1HPKU60YWcgAk3RdQ10T48Jj5d
cfDg5ypYgWGIGyAyjKdZfgyTpD7SLp0TM/kwz/IoWZfn90hVxelhp+esT/4TC1qv
1zBZWXz+yBvJ+Z7JFi8gP6y7M9soECWpjr6gCog2BgdZ9XY1YQXXzXc0bJntX49t
Gxl4ITowLGXfxt2J+lV8qonZXNnqVS+xxs+wdhy87Jgr5WXT4ro1j5fbtz9hn1/Q
YZebx/4RSuaOqZthpfro+LD6zb3nTcyaNP8Alo7kVS3mtOXQOCDre313bVoX48ju
yXh16bmxSwugV5DK8gMLssbhSZc9OOjB3Mrij85Z1jmeQeuQXdwNa8/+6RtF0hj4
kIi037ydOC0YlM04I8ja9NRqRaeXVM0sDXDTu1CY+MTf6as1f6HZo3dncWozqvo5
nnn5vzNfrqv5/1J3aeru1vOW3RWCVyVHDxQuE2fTGEEC5snOk/zpDlRenTfSXwCF
cBINhkYmRbqGhyTAMejtTm9Pu8io/ziBAH/vCbcVFH7VrDMNfUyKMh+ASRGVdtXi
2/oKbCQyfelhVTAlNywegeRYc3Nx7YzJFDEcioA+FhvmdB87ODqjRJCILqO1Hl4I
2gHU8q9usftggRqTlgxonB/fuCx8W2/Qy4I4PvkNdV0cu29p4WYpD+CXjM/fRN15
UMOjX24287v9DL54np+elRvU5zJQWWljmHiORh+CpImZpi7L++W6JstzBTD8uRMV
IGq3+NrgmnQ+BXTYdPW17n+gTvlxuxWnd7kTB2Uy1wR5giH9+vvFifmx+Mjszxw4
fvrU0WmUMc0p5jnyFEizOf7saem4XuwPxiP74HennCKshOfRCvFU6Mw3WcTkGmMS
NcPyL5yOc16xeLW6KcHN8YW8USm5SzonbOVNcOK9OAGFlQrTY5W4rIsb6laesRq7
lxnSKvDmtYOJ4iEy7hB9UXfBhYm5l7MG+Dk2vpqQmXwM0rZCjXUABbsFy9I2cLyL
CCWmu9CP7BACSbvz7iC+iId5hAxMfEqjcS6EvyBfv95XCq7NS92MEPRWmARtiCsQ
NpkOKaP1WkVsqgysMgzik+LuGC2S+2ZzwRWPJ3TRzpEnTPWsYv+IdFJdI6wRhTO9
0rhFq0oRbkxtxEpINzf7nLXjt/zFVbix/AQ6IgUYWCasDthjLh4WDXbZho9k0AaR
MCc8yOaN2BjNrjBYjwcC/y2pSUgGDNZu4vIWXknNiF1kEU04MjLtvzuceMTDGujS
YKwE6B+tt3KJSPxkDrYnB24A1Zz7h6xUJYGvnH3N54Aag58huXM4PoqPDarUshjp
G3D3lWM3QSik02QcOKk/tOw2FG1LhPyS5VwoIjW5/+hrODzKJz18HMWh06rvKPvX
dYaq2r3MUy7g1Lcc6u8I5tNMKrkKJk4aRgnqYbIKPDrDBA2APDOyreDOPzppl1qS
YoqcuXGML9Z5WGDhTU/zi8z2niAzxv7tpA66FTing2FMTNYG+I84wq5T77Q496TR
LWGSdOG8hK9j/yn9pyVI8FeOY+V7Wk/G0eqe/Kap8su+UV/V9/JEAwxCBVgMi8fx
mWtIngp4pC3nRS5YWL9vykHG+iPbyI7NKdqQxJm5KzJtjUvjyUjcmIaLozjTmT+T
KOYSWZoVyNJVfqHowoIMahP+W8fCftEfrj13x+OEB5t+bUkG5gh3C+8ahhVoA6jl
O/Xt9DKaaQmCJkhE5Tg4Ad660UkGmNO6BOwtbW4DOVfqVRWz1hkOvDbI6/BB/Cks
vKwOAILx6xrwI461bRycWqWvI2VZyUAGbaJeSOVHUUP3+PbGc78ua4Num0V9QMzZ
+6rPsksQYEC1GELzBlHWWOp6otYlHoLEPsk9ni0OVNFZa35yLcze+HfKEXRTCCIY
EZs57u3wkRA3Ro0JrB1bR5paxB4zINh+ZDCCM8dTMrfMmD1Euq+OZWDOvl/f7cbp
VzKR6r83PdLyQp304jW5AU1+YW0fKcmVLQGKv8u1/hxKrYpLPEaSPaXXThes5Kmg
XEhbUYUG374Yo1NT0BeeVUgOFs8rrVzzEWkLyUph5snx8TEdMUapbr+uU2gesJBp
YNJ7cFWmT45gcg+7rRFJvc/TQ+MmBv+drMuDNFRxKoFrVwNE1RsO/h259V8WebGb
mU5V4JvDD/HxRalMo7A4rP2kAWw+otd18WJY9Gqv+f41Xh78QoaFMfgRhw8P32wU
ettNtcYry97sRaHAj5vRy01/izvqJAdK0+nymfqHr3Z4VMilwYbtgcW7vHhT5NjI
HWty1lkaTzZI909rcBbX+FXFnuX4gjvoGUyqatze2KqarDZJZj68RW7qAdCPTxXx
qXxcW0vPeak93TpbBOESaRxB1OEd99D1JQrsKfmbift+an8e245nmD1po9AP8LVk
dpGcg3ZguR56U/xFZIEs7gXnvElU99coYdM0x9lDjR9Uf+4n2BXvTI+Q1mrppgb/
AOGT8t29aMtPaw/7n+9EBAr3EXzFn+7qRqGgvzjEV1lBp75DRUobh47DvZ+rVHlY
2fzY/4W0Xoh2AHKZ8JAPgnh2WRNlZNUvdUpqmvvVzLxeKNQM1PrG6vgzY6MAftvz
P2M45wtoy8rPh9SFqi0DfqozMrZiJgwIiy4FewjQIXRCEbvlvOLGzxJU3oZDU2aY
22BO1izqzS5f7pAL7vuodoJtJNcxhHY0NicL2TUv+b+bnnTesbBqaWn2aoovKGrg
VfQgFVRCPN4QqrnyjpF6bW42Tqpu321821oBdI+jTFZxD/fghmGKRBLuzJC1N5Hv
/U5XMit3d1kqA21ebTKqb5bv+B17rxxCeG5bozAwar5feI/LfoV+muLyDNQquoqs
LJWHSNHmGfUbJ7WQOb8/xMy45YAINZY6bC6Uq9B2Dz7oSXZiZ8ULFLgpRusi8r7O
IrjHr1YjwyLC6UC3ibsmnXaLXIAktYQvIbTLqjggrvDLdeqW3H7fqd6FnjjIQXHV
2mdB/kUrReW10YR7aFGdX3NHcr2SXqE6FMiJCnlY6Gc0wtJgP+pqoEVyTswQHRVT
p0Gi+k1J96Rx8D1mZ65s8178v9MKBXfFnX3yGiuznpyC97n23708+TPx5yP9Y9DS
kNFQTDw+TKP5X4ZcmtJe50+YM8crWRLfVoqyEH20s++2GA9Dz+jhSvTDRvTYMgPZ
nrHzzM6uTdW90Pzc2syT3QQF+SD/xYRZyK6mE472ZT9UfQezIsLWNl7/sA0XBgJZ
I9Rde2HdsnPnVqYPocJ0bQjfn10UwLBuZzEHr3VFmDwGFNBSZt0flCVqXW+kthxK
WIVk3o3WrMaMkoBgc886g8cQTZtRAL+UCw6RyDKbbxdslDll9x0sK8wo3s5GMdXJ
MdWkB7SKWAUCmuQLFa2oA8XbRcOTW4HNJKtZyclXftEUCK+KVJTS9dcl0uAgQFbl
mFjjotIM4zB/YcUVrUcMYZ3nVQOBWujOASemh5UULb9/c6N3xR2BTaFKMwDProDt
In7u148kiMEKy/nb47zRdf/0U7wBJ/CDfxlhXG9TAgsxg3KaZEt0KukkBkq01H3B
X7c9UcW6LVJ/xkF3otedF3boDYuQEm+htrxK69XxEZdSQqtoueytSf5en9EYcbOw
fKi4cRNXaZpcjJPmU67P7BHYVLe8m1nj+z7erI+ahqEe3uaxEaYoUsj0DVWdbS0Y
FJOQhddKkIqjgX2ju0MREYwV4jqPtuXwhAa1KJ9hWootIEYjNxQA6xsssrAL8osR
PGEDa4dI4VXjkT/6X6RRMmseXpw2xqoMMFVCsgizrtZBAR7LKpfqUcakvGymNu8J
7najqz7PNu1r15VlL9mn5uUzMBqqBZEfqIufsdzADL3gRha4bsUw0QgjncMOUISd
fffUuswrOot7LSLtCVhpDihztO9Qs21ndwddPErguEVsP6NGhRWQdgQqiw9riT7b
NH4o7L95ONqyy2kJk2uHGvgrubd7SsbO25pvCvC9CTd9pgCbX+FAxDGrDavuFl2p
AahUsDBSt87qDAYKGMyhRhuBKxCjvBOLQ1FxYlvEPcohWggjPUvd/Z5flTT+PNy+
n13JW4/TLArGXMb1a+nU9E79bE+XMo9oG/XUxXBi2GFt6wD4+yIXlHKBVBfmB34i
FK2jkRHZ4qVgPlAUFQeYAnm/XEO8NWbsVmFk6hf/SBlgStJbWPRpXtfwCAts6LG9
DPsvH9tDvfH6gZo8CMmHPqgtWpxRNiE6ia7dLbjiuNwXyjhoFqE6Z+0gf28z9YnV
kQ7/MOQHrF2h39BohWJKtV0PgLckcH27Slpo8bxZUA5whjqacg7xOkg66q/O9wnL
DFvsK+NVPiU4ZLsNIS3Y0zmgFvewgXg0xVBWBSg+xY8m/K0RhyJFh7UKVWBD2iwO
7CyHgaIvAZUIB3YxlZ0GyPoW6mucNdwvNyc1aSy09dyVTLyv049NO9igDuMWJRX+
RdsdV8mDffkUXajY+/TVs0l9ydgIpFkXROrHQlBscFwQbgogy1DiterFo9l3+9v8
HoXi31smW9Xr1eRsbDAK5Y+9aJrs72rPff1WZuZlgkTLSl5U7V/GIkAVr+8tLAcE
ZgS0Hb7qiSZWzDJ26OSBvNZkOodujBxlUt5hYaACJsfXDcUKaaVcsZDIMVAzAooq
ezWjR8G0oCad9zpOXWv7cAa5jc55QisREB6yx2KZTWkPmy3krfv+O9jq2DMwNa18
iBpkiH2HjrPS6JfKV0/mkkbkF1RQsCKPYo0pc5oy5XURcNZqpempyawkh6f6s2i/
Xj56DycZu3ySR2WFeY9wgj9cIbgcDuK+W1cV0mlvNPnxsAYdDQAZy/XgyeaNYpcg
LKlt2tGyw3MGTa9nJDuYgkO2Ng0yl3nQpA1QFTvm4Gm6Lv1viVV0EnoNQTCCfw/h
9s9dhHBNqRJ9onsgEAxBwakx6qAzgaauhOGvaahN8l2x8sbKllVI5UXKICJcCxEf
DclD+pqTBBKC5LixuI0XehXeg2PH9uz26zNsYiaOGSQ0it1pc75ey86J9KpWFKT1
qJbCjjEVDiPXGYUNB6ZqC7IdHGvpGfMQ08zDj/bXEDgsgykUpehWQdP9k7K19LP6
Ijeshms6LsB63QK4y4Swzwmi1XeIV3jLKwsc4kefrchF+mr8j2C08rdhVX6qvAyc
54VlX7l0vPxEETZrD6Br1uwkvZsnww3SjkEDgXDrgd7b2/Sw/rIZZi/axCrledQD
ScVQacsRQ69Oy8HlLcZ0EZaCJ2mNU4YpNXxs6CWXWoAeGXQm7WXZiyZz6QheGSGx
FLYb+9GDrP99rOgWhbL9uwdjF8oHHEGAB9ZMBUV1kluQrYbOZuF1HpvH48TcICeg
qQn0VTm1cd+ROkYmziBmVVZDgpRz31ctrgV6jZaKNmzfijPmh/NF/lNnnNeQfMSV
m/fvEs/h8SurmZzQFbeijUvRzfbxB8PQUn+Yt+iZPYQsn7j/Mxe+tG+qCgfoLd3v
8rFkSyYipeMtT4IRuLJV9oNukrVQGOp6Bm7mvRd1ikaypWAZPAjOdzVhm/73rGHi
OaOkKToDplMuXvMjpOC2lqXyMkfRir29VZM+YgmdgvbtGtnp3h4KEfp0wwa/dWo2
uyLmHp7GIZkMhPn8cimdACngcO9gRgtXaZMMQCYxgpTxCIlTwAR/dwCnYe1Y+JfO
XLFP/8uMLLStQe4swg/Cv2Uxq7Fv+qz82X0Bnbp5XdoQTJixY1g7fSE4SBReeLxo
HMD6YjojMiXnLWK6IELwHKTESaj+C0F/qovpYOxbb0aQaZUdP6gXKqBADNmPDNKP
Q9eE+QZoaAarDS0+s3q4/8SP6JrNgcg0wyQVCivDlAKNhFi1H7TNHzpBNowTsZhN
drGr6TpdjSqCjcfl3vYNYyP5tKZGY1KY4hQfxuCB63VeCkUBB97ZADuv6a3rgqTm
LkZ1KBzwycDQd5a/YyfaXDXuFmTalxthScY5bAZ0fJuVueOJv1vMNkq0qjjyXD2j
MWt85nrq85Cq71A7+WmizVVgIaJmwHn8ZRci9Jftj+vR/dB9RckE+PiOGc3RCgx6
2d6aLsH52AUMQ0wbRZhN/YtPetG+0HBDWQuJcGPGUdrdbQcsIdaAIVIRqPzySmmt
743/aIzm3/c+IGv5ua9hcr6xOgQQUXArTmjd61whTulajaLh3jF4pvGIAUPMTTol
ycDyJbBaa+TBpXHY6ytExhiZKPABTWTgpsS0fI6bwxsEcFu78NDkNRnrPo9itS0p
WwJtQHbYAyjjaPYpUgZKaFzYzsdYMlZ2T9nNNNWa9QFkQdvNTKS4BVdY5c4qWjqz
39ElOX3TFlaweYlIG1JRcHRzqccszuSUieSsBDVuf26cR2WmQPBdb/0ThKGcAYa5
F7Z/c62qO4pDg8AopHuCsRLs+hfS3RmmDh4MvcvdD+fOGT9d4spZo583Ot86s49h
Yb68y09Sp32HRNfGXspLeZ508vAJkzAN3OtGd3RAegFaicvsMEDO1gTA3SLeD3Pu
fQkYEtPtvAniOPN1rN0l5xaoQk+pp8wqUQc6wqtjx0oiXbA49Dm3dTvORdJQbFNQ
jZps+vJML5HdoMqiOhmUHs9JLdETkkRi+tAg/bQG/yEZJt/bTPiMxffDErFHtDWB
cGxqt5eCS1gDFqJKU+7FxhByT/642kPAC5XXgf2Di1TyWNcxZChNztCk2mUhSUvJ
frn9iCR49tA7fzOtSOm9IY04Ec3ACMm2lAkN5tkhV/c2icmPRHOvfcaZ0SyXIvHb
DLAiChA83Bz+/Yi6KQkFn2Py7qafc4rapD+mYsvjIgWvgIlKRn+C4RQ3KkY9EmKK
mDXkbqv4SfWWfrNYVjcTrbaDePbq1p+XcCap+ZqZo0iZISKBMt+vd0bPMG5hLs70
IRgvXqgBktHjRS13SJB5QKYuMxmuCykPqV7KwvP0wwSkf38e7ROJBUh0GyNleEJt
MNNfxioSLzb/E0WDmjhh2UAIwEz3zvOiLbqmBVlItXlZXoOaqNX0OFhK55VHUxh+
WM7vuHqGeTbgAYlkaqjkJ2Qf67gtJCrhEx6ml3YBrqvI5GnYnHm9QkBFkJ3n+TYp
Y4xDUw5EvpVEbk46tAENayMKQk/j2p86gtkT1VBl+gTuuTYAu6JfxfgtKPgT+aMx
Fb/bR726bsqTgfWcyYXY/luFyd63o+QCX5AeU/YP6ANJ5IxI/xgV3vzoY4SqWfg7
2+KFVj4T7VrKsq1AEM1yLizcaQ8PfTjFPYRtbVRFMZccywiWlkJKlQYaj/mVNQwX
22T1aux1jrNhKGy/mUqkeJ3zrLra66lVEtzw876kRT7hqPLfTX1gKnqrIykLQrs9
3EPNINxJgH4oJI1GhLH5QXdsZ0oTjm1ChbUkcs0XCtx+QB+YHyUDYkNVwfZFv78V
Ybn9P/gomew5gv1Em4CMrUYeeJBk3VeTl7tuhtG2wbcLAdup7rC41PiFdMtx+aW5
k4fLHhhgVA9rIamGBHvXnqmcTn7Zj0/m6ImP4H94X70Ox2mvz+hsBdCsNSOHbOur
NH0Ep9nnH6p3JJ4rDkc8iWANyU6fgfDp8EGQ7qOxZSfFRIhCp5ygiCH2olGQ49qc
oAjfY5p0MPfDEtAzfbi8/CPIKoc3q1Q+lXbciD/PBncT/nfF6WxVWzhsRy3cYBW8
GGcAziPUK0Gc6epafNrbjzBEiGeFIOveTrZle43pDg+WUVgZlcD+zHISvh7C2vHR
Ekb8ZbsEID64wKZbt9Jz9ctp6VgXHmMyXc9TdrFFIz8aR7jy2g/VeATzDZxMULHV
jPZFE6FYdduSp9EWgfp7txg+G8xBBEcKJZEYuBlkV4Dp7mbm1oV+xMJrfhXgbxcj
Qhzel3IxFdBdK2iGk9Nk64DioWMJpmUXEIxIo5eAdp6aey38kkT0q5VKBB8QvHJH
2NphPl4QMUMGRr1db6trNCjf2CDKH4AThzeiuiNHzFIawNV9IDy1C+Kq9q/uPgmz
Y50NYEEt/hU6Xxc+D1AGJ9d85fMNOcZYDHRLOyG84yngnGlpOJ/2kg17mNOTlq9V
0x7RpTpUE/pkMFYPIB7BpppDpOBW4mCObWSmYd0AaiXUqdctHaEYSGZTZJT8ikJ4
MIlO7rye/nswKdS+UiUwY3Ku2TWWiippKjSKflrVsN3Rtp2UPmqMHbuPzQ7L2YGd
7sbdyuXulLjvcTEHYWsXTtBMD2Z496X+vPLkHje7NUbE7slJ5NuIaYZDc1GmIrn0
CIOQh3iTqPSfgx0jlqU9XQ2KPfq+CygcZlQR9uZ9Fq1Lo8TZOduY9F+wiPL+ZGB8
In5+K3IBdT1etcb0jm+MNrxyEJ2uIRtUXrfh/Ihgakn5iFKUuU7kt+hgZPt58VmH
xV5MaVSZ6wRdy1ENelbOsFj/JGZHB4OQpyBkerxUD1KhoScgdtzv0rO+LKWVMXcq
DGXVOCU0zwlWbTwcCdsUsyzsYl7q793IlCXIIKBz2AoHhuwN1+y72EMPvqozMKdN
gWmaMmnTcxuuss18551ppD806FQ8+f5l4E/Tr4cjrNMi7o+tQSx7euxxcJQGhu9m
Ry2O7DP2b5VBMDq5h0PQXcvEsIKk7TgsE0caWsJSmfkbgx2xOr0SKYzpbvuSP0Ua
QBqQKBqmZyFlweJ3KGo5pyW42a7tNlbUUGBOuooy0sDewuIi8+mt4jUMqgRZJvCq
4u8LswK0Fy0lB+cfCGP/OiFf0q/LQyINKWarLL7aBgRswtcvzwnXBmzG+FRsUyHm
4cfkuJP3LAsTZORZF9SwaZvtvr0ra6K/5dPHABgOVD8oVGjUQjV9h412CUdQSybj
+0gppcOmSZ/pznWgVn9QUX6dCxtXZwQTMRXSMjwEiUbfDXBgAd5vYPkPBWpkd3kX
9dPSU3jcrEu7peKm5/M+iftnkhEq0jp6J/4t7Qs7MlPW8QB70qH579jXjAbhv5zB
tF3ASDsiuhv804Pp5Yg2/cWJzw2dtGdpZnMf0bQ9gjCdDE08BQ6fp+ypif0J4plz
kj1YztsFk93BloJOUxuGNy/CZ7hyXTDZc8jpTjmbq5ZDCiahLYinMZT9NqpJb/gu
9d58rdJMNl+bwl2jZE44bGinaA4jE/id8PUe3LhgtGsqNMCTk8eR6Pja70PAA27U
4ERsjPB1eg7pRhUsq3tn44EhW2K14ajBp9YYU9wKQZErffCz94EJRFsseoI2bLnV
u5c+YyiEL4q35jRpQtWufqSyx4QMM6TZLKjPr+quzvddZrn9HmLybTFL0Q+e+N4F
xuL/RJGSQ0/wH/ryLkQO9HWUdP+N5yf7exGKGghelUYKFd52w1TvGw4NWTVr4trc
viWqwvAj3o4i2aXmJRHRkGEVSBLuPVn1poWUMtMccyYFLlqBX7vfAs6Vy1cgo5n8
PHQHQKFz5DrIwCXBgG6Ez5WjqxnUWZIcfakeI4ImBRFbPAjoQN27abw1VdyJ4GYy
lmHvyJwEM/4E5CBX4Bz6kOrN4SOLwSltkrbF8rJuIydDoGAsI5dKfCYErMBrp2BI
Gl7E/UeZLGF2KgQ3lenGMMFeedSY8/aZMElAGCJ9ZX1sh6ju2lW9a6ZI6EQ3cooN
E6924UMcqPRqpXbk6wl2VLXDwUtFrZD0IUn6//4993aTgvC0df4IeLuUCnSOKUwq
dv3TeocYbFXzKtJWg4Q6zEBKUkwFX/CjpYGBwIf2149MfFNDqJc7dT9inQP5UpoI
t8s7ln9yDrEQmC6CUKTTfHi+6Ec17IAp6lA+bqj6oCUYKlN22gqx5FhRSt13LY6V
ZUHRrfiLEZlrhVivivQWM6+AXQTMpbA/zp7z94g+lJCLVItOjo4UmqF7w6Uxnalz
BbNRgYdCy/x+2049bnGAuP3pGmN3lg1xn7YslzmjpbfnLIAFJDKGGcbuL1OytZGS
yte0Q/AHo+ozfLI3O+4Vqz9R5i+afK8aAngwxLOr+xUD9l1VbAhj26shBiQdivzT
3Xwn5pWPdI7Btk+fe2Ef4VR+0xewM5mfPGzwVmYzg36MbC128jx64nTJGORH2VXH
m2eWOkIQscfYBA6RJi91wvizNKWZcDc+kX+dSxk7xry/IQxEN0YiaVydgEpb1ioi
RwHo9ANMg8nUeWT7f77UHMspT7gKiGEGLR+CTHe8m1pZn55Xp5bb16wr+LXj7F6K
oR3vNlcHJapp/su+lyp1ZX/XT35gs2UNVFG3/KPeDUSAhQHBEz8bt19JdllQKgC3
hZjrfG/1k6qv5Qj23WYtiv8ZfTc/xYFAjTWXayNkKr4+GXvGFmC/1CFquKfQS4wE
0saHlDgohmAejHauB61A2glG36bQ7BLORwXevKHwB1vK3YjOdGypD65odq5ua0xK
qoNZzlKmFqoqsY3Uy3/vYB6KOnFhDKkVAe7BdNFM3PWIZAn65lJx0dAWZoidFp7l
FZDizWoS2O52cqc3FjtjuFl4Eg1fTgBMW90HxO92VB5PH+SOtK8AMTMCybaY644+
vDFQdaj05iZwxcVgcEhtgkuzgVbF2JL6t56G9xZrzExCjhRZlyQgWvw118YD+gmk
wJGV7CCd1zJUP8H07LvQ9POCVoN+enZrvjDFUHE/UhZa8Gonf5IK0BQEIcTQMns3
/9xQkt0QbOEsLal+0+xJFQYrvQ/wq92q9Lvfwah1BMhCkG+gLPV4tqsz+GSlhiP6
q/Uq4xgSTWLMJaRSDpm5+FudztYGOQKVCN9B2M4tjRO8d2KjYe3AvMbubf31M9in
QHT5Ae8IRFnu/KlCw3oYT+QYN8GCLwy42XBh1t+8am8yRvsX8dHeJ6EILMmWT0ok
FOz4apNOD59EF/fxkGE0I3awsJ5mkhd1WmfakKYZbCmW/oqMgZOS7hxu65klMToj
ZFJ7KEkInSbLAcoLMunP2euYk0voxqndoo3O6EmLgYrgCQjrkNl1kSrYYSH/dn5g
AQqwfuNwubB9BjsQGrcn1taS2D4stPvXWqbNEVz/8KQ5riQmHf10jHXsyGJtMBM2
w33vXoEATorvR6gX0WifNAlTstkWA/MjpYUR11kd3D75jhhFlk0hThaDVY0ybdlo
s6Sw6cTopBvj7YrJpDE0CHiHfcbs3e5qfDVZVXiFOFng+wo5BstUk3Ruu4BLhuHI
SzUst8kHG3aeLXQgRxaNgxsNEaduyMQpGsRFHBOHrxVIUjn97VtChs9UI7C2qTKr
96DWjXdOOlMEUULIeLXIXcWXurxeMQFn/7v8tUPLTCaM4izzLL4/hcDGL4WtXDuW
Cb6ObCR50U/f2m59CiO0AqQvv1VaHFWZoU+K4Dc8a1i99gTEzzpGiG4raB7B3eLu
U7YCi0t7NXBM0KK8BXAQyvEMwdYZK0pI2vFqYYwr4e54LCGVMCxB2clt0LQhoKHE
UvFL3rDXWnFf6VAuwVSp5UU7zfJjT3VhEvEOrnjnh3kjoVC85l4mD39rDTtfa3Ou
jmvCINsJiL9U23eOwc5gKExe9tXYzmiBEFObry7wib5oHES6xxYT6dXK7FiquFCb
sIFa4GVq1ELDQxcDfEHV7SX29ouRqRX/cr/UyXFe3SjZh3Q0qq+msMMli+f0qCim
GD0zwugpTYpSYsQoj3gvc9asZloTaPieMd2lOnG+KLY0EWJk6d8qFjlCDadodUOq
S1wkbO6hgNXsMraUWtWKpy4Yx/HuU5S7evPllaJlAMK4aa0hDXnvEUbXsMNdENJM
du0iw647jfjtkhNcOVb5tjNut35xrs8QQV51iR0mb6qDAaJm85N709BedS1ux3Lv
OqabrE7xCFzSxXO7jVg5ODez8nKir3jhTy4y8cszGpTLdSy/0cAyMQRKG5uYwq44
q7sInHGC6vNwmbYeRryGK1iuzYQHPoBGCy5XbiEhiqcm5cFJyXQGc6TBTrbB8jLX
H5ZzFPcr1E4nrWia/hoaP6c8YMzKNk30Cu9lyWrBM/qORK0au7fMF/CgX3ruRQ7W
OBQ9G8Jlbvot5HufW+6h7OaadMqR0kQEwZaexHm0j07HDgXWD+SIs+JZbGXqPSLy
4m2tdBFZmMJ9qAStqwzUWbRXBuXImv+9wuSuiPe8EHU5+f8cQ3vU+Nw1dbCJ+xpz
/PSCIXbTtvgKgQmFNtm7VJhIdgMnFoOPP0qGpr0nsi5mq3kn/dDe+wfAq30Cw8jE
DpimNGx0HOsdX8SWi2grLUmpST2UZlzVn1+WvKBXnSmDkEFwVL/g3welZ8HkIWzd
JApfja86gC47ODgsMuiq+250YN0TPgGlV90jKstOoluDa1pF804TN7hewSRAT0eh
eBzPx46vlQIf9ltGnBFEXMHiu207bVw/hSh5goPwj0p0pEu8boDsUgvtrqiqkhSc
uQn+okQu4cvjyoTbDN38vJ2cXshKN4axnukFp5IB6uM+L0MPYFUFaB7jITGaipHs
3RfGwo55qS3Cf4zaBK2prOJlrrk+SXmML9fA+k8x7Fyd5mnteVFlEMDJORZ/lNwh
FrA9Cijw6wYP/4z7rGJ5WW7SYJFcKQHeNMI5MkgMTCxIza3rCE4DBsKq6GZGVEQC
9rgybeJj4CfU0BOsY1J9kfmNBRvhTFhyUpDiCbny1oPsoID0PxK+EeI81RX6bTyg
KlpVocW+BqBlYLT5x8aUGZm81xfbiq/XJIYKvBGm3MHqWDt7CoiE4ZZN5bpmud3h
hqhhv7COMu+qltuFqmlvY2mgwudRQsb3GCHzd0WeHYNcnr65jNFqOEHxlyyEnGXt
yYIUbA5TOa32I0BQL/9Nss2VIdW8K+ttYinZCi6W6s0K1rSWqIBjEHyL9ewz5gm+
jAF8qQIVmhHIsssE1/uI+/NvLyJrBUTDg8gAURhukEYR4DM1tNBHDSbKEfqe7g98
B2Gk95GcC7HfbY2/Ylk79NNWGTcmr0HoZCgumIgvIMnXB4ts1WPhqUgnRMNUj6MW
b4+EGj9YWdh3EUUzpi9G5RcELCzh30A1wgiBYRRhvbrGqYdAtOm/7ale0AMrhkLJ
QZi4QINu5sYOhwRECYVz57nW/4b72IuyDR8MDCQfdef+y3ByDHeBM1daInQKOdkp
WMZsvi/XRSnndcNDAkaSPlbZjoJCYainOK2qDHvLw5ZKOfl/+Mj6MCne3SwjCqo1
ab0Fnu7P74Cp1ztWYaj+xp6OcaLNuuj/92MFX95wwkZxIZsP8gNcfkCZvZ5y2lCZ
ubJGPxbtvhi7urZ/o5DnojjVckypb746GWboSUlbnlBNMPjBItKsUu/QzE8ObAkX
u5p8aGcPW1eoGIedU+L9QtWSbO8qSbrfjbA3/hwMHjhTaE1NMNrojrlL1YREs/0j
vFmp9uQApJCYoPyqdGQ3u/OXKuhNAM+0oVKit2pAKVNqRnJTVtcsO4kbzoD6W99O
K6lhY0lZaHAMQ+ABBqf7yIwRY5OtwTuc8NZS9wVoq5z1B71XdBYvKdLXjZ2+8Taq
2G35tWB02hF/pV+PeFJPa2JsP9StA0veiI3jjncUPcYD7NC94IoIzQbx0OVBZF17
GY1zJQXzIhsJPrhTFEXN/ABXlg6A/J98zC3rlqT2V1vIb88piVARxyrjK+R0LTpn
w2AnttP27iC/ThADr8D1lPhzS8ZugLsDuWJefZh/FzDiKPYXeI4caEmPOYa2rN2P
o+XF9J4JbSy4p4tjKEg0rtCeJwd0uOjNXcrpyrLXTMPiyjRZe4FVwOS5BVb+rexB
h/bhv6FiPtsHSqRnjcXqFVfTmxRecLJhiojXsNvc5OSIdJHnuEh5f2qhslw2PmOH
7mcB9nF1fOsZ+p6l9QHEKGzFbENPIGz8r4nlvAi50TzyL3ER7h0Na9B86lbtgJu6
I6Fo5+7eKaqwpO/TEdRCYMJFanz/jHS3A4P5a0FzJroj75VDr8cPtkRHYDDXzIoT
UAWMBrBJpXZaoa8LV06vivH3SWC5gmyNDvGCTj/NdiiS+XoocSet72b6nc02TL2O
ht5PKoyMAb69qHQb4IQ8Xd1jyTy4mbIiN1mOjZ3DJsHgks4dHML6FOh+X0azKQE5
XPRlhCTjP+/QtMjx62wVJiw3fRl4X6LS1BcVw9mfRGMXwVr4W3y9Is4LlCzT+Ry7
MPC7JaFVbk58+WtvUJ6DZfWCMlV42uMSYlRdNXaEVh6avxPAsTM1Af/Bz2d8sC+J
Pt4A9eSLIMOFgTEb/PMFIgplaLBkBK6d4OIHJit3vrEaU9an9TDI+ffw9DW5vHo7
LSoIHm8znurLmQcuUgB9SKqOYncBkrvGgGf9Fq0SmFS/blQkFrk8RvX2CeTzl/zM
lEJzIVe8E8bgHr66MzmMklqtw74QPuLq1jwXhKeEV6TX81Nvb03C4pWVs+J/MgRH
P2VR/xljy6XPTwXKU+DJXqrU+SLEv7IKuUHvZQONw8sVGsVtlEfZTdXrUEyBepf0
JFtmU/IKrBrmn4Unoe55+CGOZuxeckHMYIrfUsMm4NfN5CqxBLSdLQbWZUNnQ8Qm
4MDpPyb6aQOIlm3M6MILvrmvgrb3Ek3oQLvMs8BMAbhFLayJN7xF1+b2CF8ZzawD
AxfhIAt7eBKN0HLW/hB8FqoNIqIH8+GKL8h7S4MbRLxgXpTMrsQ1h4brXM2BtGQL
KE7p4ON7Pfqr3+3xcCydExaNbzR5RJxfBzTNo45EqPK8NOK3rtTjGwEhN+FjeyrP
rpQzBVMNoByKj5fOfCSwuOpzcvx6ut1qcpNwV/8zefUw1oT+Ju2SsubDgFfuB+KY
D3YG8BXq06pnvI9t2FAFahZWV4Hz5RMwHazfxngOeLK7/rOGg1Eno20g7i5EiuSA
YGN5Ff8+Cw2QQDBDUznZQHO6E7s0UOo/Dyrw3p0t+fG8rKs7izmNxLuvh1FnK0b3
P3O1rbyZaCaMi5STgtUM0juxP5WIcuCOcV2XRL32J/rkfZpcYZpAGsmfPeWE+QcH
xvPRixjikTWgIQWdeUeywyznOpWvae1ifjpkgRnoFR2LEmj2eZfiJAD797MfnRCJ
KN8tktDl6oBkvULl7QMkW1jNRMKnw9XYjDdJDJAVlvbe1LE0t5cZJUZxRwscPqaF
MO14l8x1ixeIuTv7Q7AC9U6Qa6Xm4T0Il4FgP1mOFfr/8jCIo+Q76LNvRWJlPMvb
45gnr5fihvBPOi8ojyCob6Vq2pXq2q+1GubZd10Vpk5qKbXFrVe8HCexErNSkTht
o7Ycn6tORNy7ccKQlw8EYe/rQlb0pGuH3Ik7OlI6mhVzN1tW12dL1GMzDCvup2yM
na86NU2KVh3tnrXiDg9nnAIYYsgmPyeXdRPWOZSmbBftZ597bqFoq7dICga08h8g
+W5FgN7V7TJm7PrPBT2drF3fnnfqUsQQaNcysFPrHoKeH5kapH1GsleyaKQ/p5XH
anEE7CCLzwYdpzGb9iEU/Behsd7ZwzFxsyYvAZJw6++7aveDo9uGPTyhtuPZJy46
F07EmW42Kx65Zc62e4tFUWlI4+nCTq8bL2oG3p9AxSOpvadHqMxeVExMYKjYB0mO
b98RXTKhSJiS2yVRSbGPc4Uqab3kdMsx+DJwVj2k2B/8SMdD4p7p7AmXboN1e/zq
5fgvqCOh4ep0VCjjrXL3gMjEbrt8lKPs2J7nDRUMGnsitaaz90QpdfmmuMPo+TeY
DlNQkmmkDRX3D8khDSmQO6vktwTVIBYoyKHgqQko6ltPmR941Y0xMKKgDl5NqMO6
VIOxb6OeKQiOJNwJJpZxVjCtP+ab497RLBMhVKwbCOE8227TMegCSll2tQ5tHCh+
3+0gqM30Vi8K5ASjHHtW7YgwC3yWZZjuwaYgD5KX2Ul/u6xhrHbnC9GM79vf70YQ
RoWnTA+3HTblv6KH+gpXtr3X8nOPV2Me1srH5sIM+emmHjhxlmc+hrdARQ6c4KMc
LaEF2XilmBUAmgUvI+taI05aQWnXzgE2dFaM2mdYxM1v2A0Upvdta55KOQEVNe0w
13jBhOdNGSkpkRwhPS5r+w1szxVD79sAO5TbiClmej5PBKZx+9hQGHH5F66go++p
VuMK9acQEXU9eEqM0GDbJmKd+7ln6WuVvB1kfL0THtGviPzlf+6kJSblaS6g5uhg
VYJNdCczpV+UQD+Xeh7qONzAWoTh4vlgKc/Qbgke8UryVfwbR6FBo4JgExMcHF4B
u5hdeqGgV+F+zwcbRymBWNZczDYPCFwEUKcWLZxC4qmSJxM0hCbciseEdcft9iSz
NZ1v88mC5sb2BjgVbK3YKEg9aaaBsOOFl3GqHLaEcb+XGiUByb7UDuGDj36/iEWe
yUK30pzMXTzjvAlJmOe14EyBokhq7R2Ye1VVKH/zJZybLHfyp/VTZ3g5XT37FQif
/0VsaqVF2a1Tns6A9IBP+fMWpMJ2OvjRJLrk1GyLtU2hdrOkun7R5tqd12fXEaW/
zsXWiVkrE8VVAZzBXVkWGz7Yztqx/PTV7ZV+ZAwdzy4Qz0ktea0RIO2CjtZ7MBS9
1pJaDK6KHVrAYFMo88fn8eRRpaLj6nwEnvxPLDF6fpfADByRFSM+BJVtr5bFcN0k
WkYVd1wMSZK2kqh/eHfaWuV71CfocE6V4ffNUPKu2Y2xS8FekKEFufISARXny8Lx
K+htmamAFThpnOTEJS7ioIDxY9oFCGiGXeKemWINGEWcFhNy98/PfjH3jWJwDdAs
NWjWw4rBVlhSM9mZbKdtQA0y28XOgFQLoqOcsTBJJ62dhEySztVa8hjT9dSm1zpF
wKq2XcLxE9XPbyoz1SHdzCVd8t/TNHKmYs+tjV3kt7Hg0KRj4EX4WPN4W51KZb+U
Kc1caAZJmY5THEQu+zfNd0NbUTBU6XKeDqPlCu8ZuYVDyxVIIgD8H3kmy4k6Tsq0
OA6eBzFPeiHV5gDYP6Xs7FCFJNv0b0n9eOYEI1hv/tzqIxyZ6nFJJoNgGGUjS823
U/AB3tuOjHC2iFGfftBz5Wg3l57x4fkHsCjpFLh5Kne3j55Suf8//gJc+1gidZHv
n0W5kiulYgKUTxmbt1y3Ufa28RuXjezzi3Qh1UZlN1odlvWNciAz7Ic5vquc0zop
cfgn37lgvB0ryyVST3DVphOa0KG+PlHi+ouTZGodrzMRtdLbH5XOngViopfCpynC
lV6yVRdIJDGjJByOZWhS6tUeU/8LWeOgoCBH/vUZpcmKX0/WE3LktDWZdtDseoB7
dLdcvrCcVRumbAf7We6GNgpAlWir47FuLaxYTSNUNoW6AABZF0WN5Sr8kG+fqGKd
Hrly983XZfD0AL+u3LnS5BzFphV/upa2Do892GF/E1q/TSTV+OEYN34geQmRftfg
7H3AVXtMtQQQKpWJObP5RQvP590QlJXIr/jwNWIFbaik2i3bTap4LKVZv7OJo/7G
Z0F/LSRAHy/5Tp/i5FlPk9+soTN6qlSmzSyYYVqRJIwwSeqb3R7OqLmPSaOJxYRQ
8Orr7T4coqRq9m/YtKo/pliI4WZzrzNwB8oD0StMB2WGsD/1k5/h8SSPQYRERN4Y
rag5pAeTokDv+XDUDZagIc1SpsbwhnE1e4VQA2+POLyDBYIQ9QN4TpU7ICiGrVBE
uqa/OPOvVOA8ykMCse8xAqqTCuQ3mktCsNKsGKq8SFqPrvzOa+gwJJ7yssi+A6fa
Gdqgcnn6tccy6C9G+njdFE+EpHCIWRKfkzsX9YeEccReUmdsKjXR534x0eOJl9PP
HZc5un+0b/RwXrjZCev00vhZG/yQ2hpi4KrbwuflEcppGA6qwDehe5MYsDA4GFzg
l3NmAFPl1iPBCa8anWVv+dK1lKS1hGvxXmsPCk6Btrxx4c/fXN6Ot7TzVHW4Axo4
GaSV4rVz5M71DLrbLJW69vnsI2Za11sagY9lVZow5JG2WW2BnEVnFZNXio9OchZe
qczr3BCPmdvHJrGx9CO9AJoH/zVr8yGf5g9n53R/SGHH4oOLmR8GS8kSuVzE6+Eh
kye69Zy0gjuCRqmw9XEj4hkNX4ODkwZ3ADQO2H3ELDRVmR0ychaaA3MKc98zblUs
ld2HSm6scmdmbdybrzHg+SljJgNu44CA3aaqtgZB/MSnwXDzIk8g6BX3Y4zF3QLV
H0DcaRsy7VyN/Wi1MVUdNl/eaFixSj04Nz6/JVVdbtiQmbemf+SB8Bw7dB4D10rW
3eOIFq6fg4OtIomcE6+A0cBizEGbYnXvamqRVyzy/tFOQwew3qVqmj5kF/YmV/ap
ouxMKF0PKxQp1ggKZPhyvaXoFu0ByHIb764iclIN4cdWIWG2JsYJwBkSo0ec9vvV
nku/oQ+NFTdCbbZBN+X6CdbjplB1EmjnsnXkRHiz2gr6SGQ2Z7OcLgDvwP7o6atD
15xZeDMNe33+2156RY3uDpkP6wsyCuLDR3+J5vQfmxyh+DjqGWNC3p9yP4cfp6WB
o24H1k9UuBDdowhFU7KACCxoQA88tm3WVL6szXJwMBFwGb9e9Y6rRCErymCj6nLr
eicA2foMPUb2ohv/ULZrOjtYuaGfs2f+It9yzBD7hfwpIXHYIG8y7MOKc6OgDoOV
gGq7V7GW+//ct9uwFXcLnjB4BcbXZqcbzwwuOgykLwRNsLjy/nQXfGk3CXY/4tnv
Afxtwjx2usyiMfI44sSww+dcVu23Cx7dEPfPr2qDX4hrLIMhMbiA49o+QtNRfA/r
Cw9MZbWPN4dPLCwxJ5k2b9iTjrDdcB4KSYlbUp3UeA8iVZE+6Ta1sI32uVANZBjZ
Xo9e1dUw5xFk+ZSKtVV+tZxAk173nB5sPMwe+ib0Wde4h91d3xPmS4MNAXxMXEx/
BC+808AVKUiegQ8YUaBfv9nfy/wqR8yk2CJuShFCthi3C3+8jwyDopMD9m92xc1s
dUcYDRADG+rnpnnf4FPpzlb/H1cq2a0RJSSCuQJjqz1qZ/BHSivKs+R3kuplubKW
fYhL0c6qkRLjHfT8AoMCzhfCaMAdbdT/bILEgihBC8LR3ADBpvh6qx6QnS9R1MG8
KaI4k1/16QcH7WTuGNWB5ljbx8BPa9tzdBUdQcrAaGmMU7FyZ+TIhRM05CVZub6O
Aui0tUN5xV+vyIWSEgY7NykiAdhhX9NwVKiI47I0DbpkbY6fhty91VhN0zKYm+4q
J7ng6/ybin8IoFGR9j7L8AHTi7CFCInbdQzMNu3/4upHgigrAP8Du+/hUndeGCSX
vekzYNHgg7B5IA9ItoZwhCEl6hNTE2m4SMHt+h/mQOgA76yJ5RTOYE+gHJoFdbpO
/Tkuv6uwhlG54SKQTtL/finoMXeU1rnz4u4+t7GxMadp9GITQiHq4fLW4M1lLCA+
ZBK3HKu7415M3hoc+5T1Jp/7SoFv1PwP8/dJmhiZTQyJXKM1d1qMdTl6cZ6uErU9
vvEfoZPw3Nw33GqY8prWP2/OWXIFKRq5VbbM3N3CB0+ODHXXhqUf8jL+ifQhyX6J
R7qnDBsn/F91qmOo6XWtRPojDSJESFyPfxlhQaxyRvH+f4BY4K9G5ZNS1BmRXys4
4AMXWh3VIJv7cvS/KBsklJcCXPHLZE6jeJj+929SPhOZQdPjwdTkR4x6rVxko/gp
v+hPeERTOfp0vbWxpqwuW/N3Ju1gUoWWCyH7gONxbedSYf1Rt9jjRi8tViwMLeCS
53tcd0WxrzS9Z7slt5ED6M0VRNiyLvZzMMOT6dwfcptUBED4nQO59S+pyMZG3H0w
21JqRFqhjn5iaQNkaGMVzC+YOZgRov3mQLKxbZLe6jc2DPExrTGexQj9ClUyU5Ui
e2Xp/VNtSD3xJbaeXGYBoNBKBOWmbFNSIkuaiBSUalK3C4mFjtXnO14LzhTClQi1
gBKyJmX+cVTIcSzNNBaqFc6c3SNhH3h+GPIU73dS0ehwpw5WbsaWerWwGgDiBYnb
DZsNaMNwqYJf064IN44GCS7GhbOGPkOP6SjX2mPCAQY8BuwH3Ha1/uSj1IG309/q
9XQSOLo/bUXXA+ot4FRSCZLOp7wldPaE+N+d3FWmf3a3atw4JBlqgsQhzEEqdvLn
dUG17BWCU6PmBoUvUY6HDXcV5jJFY4zDGjNIvp8QAOh2+BUVYlhp5r9YY/8GjeWu
SFt4z3SgG5RpN4jdBX97k4CtWX8Xqy43SwBxsbkPvWQNH2rp1+3ymbWm1zCykwm5
jcsi9BQDaz+2DcOPjYJSFajvXuxbBmwnkt4wiX8a1Jsm2UwAgptfzCC8UcHDGtk0
3BIqxrVxRVOIUqZ3WFp0eKLJ5LDMcN4k7YvTXYXG3pyd9/kHeUJBIWUK0LxUcDBY
2KNaIFBNY6LASH/wCEt6C06UUb2fiBODoxRtyrRYhd2YiLlM8GVxbu00r07gIXUN
d9Jm+7LBsYf7iGveaEcy5kPr8Ag2mdFrQJLlj7xgAJiPEWJzQDPUagHOd3y8Hjxl
R/x5cdB27jj2btGX4BmWnvMu+eevohx3bcaz8EdukFz7iJCl7RL/LgMPB+8dJtXo
uLeb5Pj/M3KpDg/hr1N+/Satm3aiVAS41y6AKkZyjtEU6JJm63VML1rj9uW9WZ2Z
AjZ/CBTUKAlIanLswYaU/873lxnjMjLm3qTA43JlHqEVnzOcXffqjufQ6idjH4DN
r2BuP4DnYvwn8M7MoW/dC2gkTmBErlhSvot1ANv5nTPD+zUv+hW8z/oknASwuh1h
ySLVdjhjTIjq30rpfP8uIECjDHm/inqB/GSjD5TbKvFRhRAgfOXR3OuSrkzmLQ/w
MtlCE4B+j71bSN5P9Y33FPcsDHRmUUQlzIDA8yWQgmxeUhFHXJ+7zQHWEOIuKCMc
cmjo4a1DftHKt3OaSP2dSPBbuYbjJsaFKlJF07l1+Ht0tI5XwY952w5kwMzMJ8wa
T+/BBZsbRWrklK/8F5pTJ7cK0VuK0Ri/X1EVmN5gzrF3duBHL9of6B3LnMaVM4nf
ooSYqxuYE1GO8tKkb3qTwdi8ECtDHmKT5Q8h+pBNGjXjEW/TI0+7pcofXQ9s70L/
SytqAdRuam+9hPxmiv6pEWCSZI6tkvnpmnMlacAB2IErvLMqkJgkXT+LM+gw716Y
TBUpELxSRJJcurua98X+orHj+518PEG9ycGRim9eKpIzZM38zDzXJn+Su+bPnxIy
vDzQoseGk6wubMjvyxBOGrnTJv0uThTwmU+kA7+UY/BserBM0QyD4lcxlFBU7Tc0
7OCYIIRjBNxuY/52W3zf2n+9dFlsT+fWH4VfRz23XqFBq6BCxdQIkpD5jCOH5cCM
Ucgvp+Hm4nJny/GTZx7kn2DlDxQ4aQ8FWwYFxzoFCMEyMR+y6MGkFbqdjsedSgaP
ls3wqUHyL2I+BEkRtwsVVZQLTKWAcWlI5pR+iU5GYqyFIojfCgHvNFqLmOvb4hfn
C0dcPTFZ7xKqHatv70wmvOoftYdGWsdR23+hyv4AN47xkBnytRycrCb6hOyS7LJi
bDIxMs9PqYoVU9c3IuRNBzMVqWzk41dbKWbYVDK4EVRMpg8RFgAr07Mbrox/uVzj
pIYHhqNKm9Leu2IClYTIGaZ2LS2Fwgw7MuhrFcq043MGR8e2jIC0A599iGyGJoie
r1hgsCmu5aFHy6WZjMckAMReduqIxbdnkvdvqp1/LNuDMnnGjBg5fd3GEH0/hO+t
862fBNFHWslLihqRefCD1tT/MWft2m9MQqfaMwVXF/Ot0mOUhcG+ezvEAkG9wHMl
cIMs3LS87NewBsta5wAP2dk3VLGGaZgSuqU6TsVBMoemJ2xyPtVhIxVhmDuLmWaH
nCDjZauUGE0Ng/7dhmSwGlChhKKi8a3c5td5EllG5TkmWhKNYsb1IBMlGxbpbC7x
ZdoiUo3tnFN7Y2t7JKa3nJFTKUnvcrgcWcYLFdcb+viql69CYk8ltXmV+Hm3Jrk3
UXlYh84sggA/rfPt7hHvOSyqnaF6Qpf0DUrsjQFBrN2cKeZhrWroQis2pbX55/9a
i7lqZT+5Hv9ZUyWZvwjXRzyVkfLOQ/mkI7SYsVqoOp7dlIj4IWA2VFOjjZU9ss5z
kqom8a5cDYZpeM8lW6ERNPO3g23p7qE2KF0GwgVM/JZOjabYxF2CX12BZauHHzdg
3sQNxW5pfE/Am3QwCSQwihsbfGG15ynfb6wR55JN/99YTKhZPqfArhQBhbviowdN
iAbYOrWuxw9nvkNb/eRhWiHsuXTKZRKg5p5kUik38sw2kx3+w4s55LEd/4HESKvH
UpGP4ZV3+TVyAihxTRU8k/kycroHDAZrZh5GxVbUphyouJ6A6BkZaaMjo56/r0bt
a7Mpj7jaPNygsug9ipsmmPe2FYuc6f19m0hDQ3wgAYbcp/Ea3eHtiZiUv5PrcjzQ
KgpZclSQlHzv+fVpFbt5HBD0JV4OANlv1iJghklcd4+1PI/6QbYpx+AZeX9rpRaa
aRxkLb7/AD9UNDwXbjBZf/7jhTinj5Z4ROWhFnZ9dCbsBk1F2n77xg4zKum5Ny4D
oITx2VCyqnW27pHUhETEUYN2xNTJiaYTCHoz4QUktSLIHaAr6bxX5qSFxdaMaOgh
Jn1F0EgsElYWsxI1OevUBUen2IfGuF6pBfF5xCiefGfvWyRKmGceNtxFhP8l5ZXE
gQLOQZfLl1xcBYMQs6YIP/F5Sy3iT/GxqaQWmZxdVqxGfuWmVqUmFwCC2a5u1Pm/
3YqdESGUmGl4+nMorIT2GZLWe2f8EQ465kDogWUk1liYmygNcgOUYjVMSGc/eLMh
8aK8PZN3mx8C7HHRUAplokkvfxICRWVa8dmXLs46BeXmDzPdi+//+XRM3TqJokyP
18ONhSj8s/PTSwmRGoun9PydEUniQg93RVqWc3pWcU2uzd/XiCzpC+QsOTiKfDOm
KeN9KVg0q5boK6HkbAXazTdrlirnoNGplSkq4FGejbc75mGb8mgeRmYTLMnLerWl
ZVf/vHDyPmPwv/AyUt+gEEbw8yn8xLXkCT8TohFCQJm9OENCxyu4Zp8GKaPIIJXA
A3W83tqS4/hA7E4Z0mb5BGCTUNZNESLWbxTQT3yf1UYV5k/s4fBelD13M3PMBb9O
k2WPJJPpxSZDXt8F6MZvlFrC+AyzixZDY9R8O7keG+LvQaV5l/Lr+/VN3a447BPU
lMi8mIeo7Q/aJQhgX/3TKVPAwe82Xy0yERMCPKhMI++ELNek9SB/kmVH+xO+bZmf
Tstz0YzT4fKg3m8frFZUPZm4ff+CZgTUNZvFBFx+04ca49nU48f0CqkM2fForPWt
ZpBbakJGFF/XmSwOXuZwMNpCCGAMf/96M/w1tr6+aPmkB2L9a4wZprgBY92K+Qkk
60c3SiNiBPBHYQ5L5mCf631cgtfBvfMX249vDtAHjfy0m3vaavZwJe6wx+fyDDNc
VfOhHw1/1R62YcEmzil7IkX0bmwEFKo74fclKkebNuopA099fu08bUyymDvHRUKm
qf4Whw46fDPORyvw/B7g0Txx8CpZNmuSHXd9ycjlWDobZ7O9nu6ISb/zvkIN3ZgE
G27UNQHnCITxl0UkX5IouiWNnZb1KaawzYwYPEgXSeNQJrr9EFI6+Vnjqigql4PS
gNTlC+vlbrkj5duP0/mpxTDOJSNRE0pUMV5TVG6met32vvjh2ALlI5WGyBaDEtQK
Sr0HQY0a9cnsqoQRIv21L3YFYRaNvqFz5cTj5U8XunytTkD4qBFjhifkI+ZNlyU8
A4A08oP+Lu/Bfk9S68xxqudUdiPfN/+a6043ucX2bmulr9A03dve4nTAZBSsoRY+
OarqymP3HVPfRe5M7S9c0pQjYRLH8H8HfyCMO5q0Imk4dlFWGpGuC6XPW/tSl54Q
w0kX5UDcVJBSKYRAUljdJcYJCBQ4mVhGpYVBTyPbtGNLCP2yYHDYqmlUya/l10bo
0i7aVtOpRLP28rJEMD+WdZXf+rR9JLBB62/GfmVYxJLvbKZBScx6jur3r8Ndf1Gl
C+FwLwMVAdJzVfG2hCxBT4f1+64PiwWvpY27T4P8LN6E1+xKCVzqteB0RlC5YjGx
l0mpqKwhJJ3TAqcWcyEGEK/5W9XGJGHTf0jk9m3XVtgH7hC5o2kUWAaKbK+17Wq2
uiVZaP095hgOxKQL7yqy5PBDBBumgxskP0a7ykVA0StA4OxjJ1meR4vSYfVL+qiK
U4isixyhzqCZlDwqfEviU68fwD/JkzDOpb4B0M9RgUY+TV9QSG0P6jBcoRPTptX0
zLnesp5SD0UyorOcxmBnKwdJ5IkDj6a64Ijf2sWyKmh0fia9qQNlqLEudztZJfR2
t79WlSeQKBuskhYDym+/wTUnNHexllLdcjibqlaFGej4EFvYUt4XeN/4XdmZnVPQ
g4qLUoUicf8a18I+MaxFvjA+bU+0SnhevGGusT83K38blmMzWoeUffYlpUaQGWnI
Xu5udsNj1vt8PkLZ/vAxVZJRZgDB2k5yFnXJe1VDZdK0Tp7laXr6u4gT9u//RV6O
PVnkKDf/r+9cL/CJetUYfchGIL2y5cVlBAdwa+rfihMUq3xe+4YdZgNPo17UDIUD
ug7ozG04KEEbTPs/x/WDJZEOs0oC3rH4udexXax8jpeMBvQmJwmqg12C7Cp+N30w
cNagsUTR95WnKjzRkQzEa8XrkpNuEUC9Q+ipAHzvKzwgPCCbnqRmS7WhMtXXPeG2
qSkonbwly/Zp3FL9+ZxHcWxSJqpn9LrGboJvaWTpi0QQ93p7qD5p79hVSbSd5J26
ex5bv1OXE2MGsh9iJzPPVNWwYSvcA1aCkbiWSuiOJIFnzXbAds37J9IAIsCFTbcU
r4XTHovqLhSHN4RHdXxbqOkKN1Fv8gj/MFwNC8k9IjbQvNGG9vsPGYPzD6Adlno4
Yj5njSRD3SuxVT3j/cGbJOogoEJXpJqShnte5zVSbWKM+hB+/5ronHbE4/TxTnIC
OZL+SQHez2kI+jD2yvxMs0tSD/qvlyz0DjAmZp8uSKNsYM5muvwxtF+ijqAB5NoU
yRX5RTdW0rg0ZYn+zbkywINGrkS6HeRSyn6fTogYFizRFdLpGRZcJSF5NHvYRL2B
ZfYsaYW+xlJlwzVjYn/kFerA8LQMrkn4oCdKEraAy3YZx2J1capsYpPAnwJ8Ppb1
Jt78bPoJb+SdpeBydxDd/5ZdpcfDUQ7tXqFCI4Qd9DOvLgK01DyhSREqqcysmua6
cFYZXPf8lIkPUrLptT4l/4lX0YpisXE5H4ZO8+N0HykkCazwMRsoJm12MyiMyMsa
T3zjIENIpab8++mAJnqk1fMnIfCrC4Y75ilWAMKmbpPLM7aEHmDWTAQMugApd+1i
qXMbdCpDHDWcFDeLt+eV6ig7WAo+l/VlpGPkhZcXxCanie66xeuBZLwPtBop73Y8
DuasHK1vWLOWrhPYc7lMO9I/UX8lh+pBQ9johCymsiLEJ0amXWIw0pZeG0wstjFa
mT7hVTACHiL9mGCtlkNQc/REhbVRTOWdNZg3IIUK5z46U7Reqs5IcIxDcdztjldH
xoMJZzuMKSD/KrL0+O8FrO+3OWqjA8gIwpFvfSmU4dwlb2Mz8+Okmj4S8vBKuQWS
9tnEGE2Rwhqkokgv4B/4LiLedYRSx4FzAZrVKw9r5uddDvOsUuCU6wFy0RUDwP4C
IgNu55AEmGRQW8AgWFDGxtKm/k0h1KrJ9o5ZLyjruERid4swgIT/Xtrj/sq88NDX
YshD7Jm1hFGqQ6keNRag/aAiG24IX7ZlGkF18hdtAGzMQ6rDD3aK8Jyw7fc0JZhs
q5zI3KfHVmfXzS7cD6m/QON4d7cFMQgd2/9NaZQbovJwslKX560oUgsLqAB7/P89
CV52v35+8NSKj9tkkKuWFqfK80XcPJJs6YUbOSoL5Kdk+58LffFPYYI9RmI67cBZ
h0XYx9fgQn75WssC3bTlGPKfYV9WjtFmLewMmjINPVspnD+qpzTDDVOGjMPgFtJr
IvICeZTXhzv6FnQcKrG8C5IyxwRHsvqGF/kTR9ogZU2dBEqRja6HxTOEv3ADj3fP
E3TbyhZqmfasP7WMoYhJRiaqoRId+6yuDcICaKx2wL5EPt2A8CuaNApcsLQVGxXv
H0YC07th+p2TkrEZXf7afhXpjEIWdhr2Frb1mKPVrMgyp620aurpQhzrfJspyq6A
UcQufE8/y3CqeAHsmKjYRZLCaoT39NsFzNt7M6ctdjWHbAJg+xZm904yOYeV4uRJ
xuQVJ3pEhxO9Wm/1XzzdGmYJVtJH980/CKgEBjnPF+68mGCAZ86Yj3nPi6qP/shC
i2MeDbsOQlvMJ9SXRTm8QfD+X51+pJy6uCWD9sY8peyx31bTuR2CsN/kIcwwi2aI
DaBSj/CR950dVI+HBvGdd9lHPzLXGpx89tDdOLy4sazpx3FPhY6zFRQEGqCizyW3
gPFnUc9CAihw9SFZK5nqZl+3d7gSmIXhqcnSGFT0b1Ae8pm2WvHAQBBcXC2rnQpj
zDgbiP9hNqH253lonJhqiTnFzIBneJ8qvN35hKmZ2DF7DB9lraYpiSyu0qh577X2
Pm60hci0xeD3g0tJqy9NRtKkEHwavuOC4YKvswdhFYTOqDhRnXt0MgWybv5I3rch
T+etH7+CwXdcDc/9rI2zSmQI5eKXXIPNglYIIzCDuxA6oE638VwJZIbV7UEVOZyK
ygj6hklWUTOkiHKZ2c213pmWxUdoz57IVYN8lwZ8sUDMveVldH3OXeFK/fgTQ2MC
mDJnaBT37iw0WcKVugqj9u/btHZBZb7exQQysWbNEmMnvkRwoUBWP4FkgyhbIn7U
Zy3nKAanvr31Hof/ArSIfUKr9qbosoD41Kv2ZwZpR47cagPL7BL0yuaUUbPxN6fa
kw4/64XIQ5xtTJn7yp1zQa+q+U9Jr8Cagpin4VmmBKm5be4oWQbmf+5JikL95F35
v67AycE64Ck37mJtq9Do/85UIBFHyhGEzTwLWyoPyh9seEK/zEYxoYTrGsBxuYF2
4wgQT+J0+1d3sJJE1T6bw6CTrtFdHhk0nle0Usbz7BlmmRkqJd3QjU5omrSauhbL
pnlp/pjd2rA4HBDPiNabiNVGYICAmlIBYGExmHI9Udi5HnXZcNNcjnUDHYp3Kh+J
P00CrJYN7pG7cycgjcrZqYg1Ww9nl8bPAYMUnPcKa/XAydVVn5dMWmWjsJIfNUEe
Mt/I6w2TLG/Vk8Bgx8pwk/J1PovL7K10hfg5YriJZmVHxmu1o73fqTMOy25Yb4LX
Pbo9r3MGN4W+DXpOnlY7BuZFJZxdFadvI/B96GkEnwdI+7fg+R7rmZc573sP8awc
WBlxsuD+/qtbPJNh+QPwa5l6ZwrgHkePXY3tgbERLDEBrd82DYhFoO1RHHr3Volg
x2uzRlA6colA/nuUrdnWWwAeOKw+g69plrjOwe6oiOj+h4c7dvJT9LK8VKKrtrtB
bejVL93ZXosiAMA3foQ8Gy7xsE2QIGHIbw/yj4FibEnZZi5FDgakCyVk+QbHiSsh
lI36RQtyP2ffzl7SKplJMhPstzaGYwzFYqOi1dYTYh0xJbV27lHNnGTH3A0oOH3X
suDmlL061e1e0mo2/GwDEX9tozMQK+9Jjr47aUUXIxXAxlmkmUn6n3Y4LsPkiqoA
15U1QM0MDzd9TLLt7DEc2KatMq9oFnSlodtgepH1yMXEF+BRofHy0k6xAIyQI1vI
g6aaLbpz0FMKAQlMM0719YE55b7DfpfHbhxXIsbca//UQYDUtyR6l6HpQ9nOCAvH
ZgQGRitLuOQ7AjIp2PRpCyml5JcbdDhV2ztMovUqzhDRMOWf+lGmIFd4hb1dprA5
93HtzBHji/k3922wDOeXeuRRE3ZposCbn3apuJ1U6BwXgI73KK0ymKeo3f7wEry3
sXqMPQlDWVXCnpVYaLSJ+E9y4YDMSX0L8Pfi3Ui52ZSbW/a+w+qNcKX7hxEVedR0
pU7T8FwaV1T48s44n1aCl1Ou8BerFl1mlksuszbZ8tRJRm1CNefYkq4xCBTYdpRp
LX1ltZtkzxQTn0coGWhyHONYhEjNakTWLnp5PGelJJe4uk0kGb/H2ZWOV78iu+9D
8LlZlIFTwR8k9RuynZRiDZA9gDldzRNZhi065AOBpGSz8N9DSYMlMYge0+rH1mP+
UNNO3NES7BKCKfKsSYd9vm5dJO9WKIdNE3f3ICk5MxL/dmwRi8nxZLluasvZ8OpB
HBWA7yyRTRSMS3Ee/DGfpXx3QUQ1JX4gBTfBcfgPcQJw16LMomZ+hkVB0g+NI4JH
XoMOJzPopnMMXziuXTdm/Ze04LIZ1knUCoKSsWv4NAt2Wm/I77lgsmt31lHmG1Se
fhnn5Cr31m1yYj7vbGHzKSxhAB3YXB+u4u9IRkKH9qsRQbGoAcalhc/xSxhdzcds
ugqGTvxf9FO1Pa7iuuGiarGE38P/O2cl3kack3ei1JDsJ5Q0SyqwAS35R7QSDlPf
0CGrEZcxxAhc6G3m+3yzv8pmx/XXIrCuXjzbMO4JeIYNe7qzZatkICL56/WJ1XrI
WuGomSVkns7c0hQVcN+i29k7wBTXzYQcNqCH/C7roiZ2QUVHUz6iAzLMccGiZ+YZ
WlUwnsoUnM0llmQ16nNrzMi4iW+1rHcbc1Btm9bUHPjFXGuVL2CaVJiKNU5twhWy
WYbi76NIyI7mlXsi9u44TWlVnjcynPkPl5nG5n4/1SeT4ni+CSdY9xJUhm+Sj+9j
atc80yTZC9Vxty40x0+oV7F8I2jQabuPpa9O8glN6XeTqonz0tnVhm3Squnix8Ws
KEfooQMWrK0luoBlcDIb8TZdODT8YRv9AT2hpZNL1f35h0lRRS9vg2ePdImwp+wQ
ff/bz9mRFHTti1JP/YIgiu1vkecQNddiBeFKXAd4KiZQ+ArXmKQYn3Am0nJWHyHb
T/KRIR+vpHrMnPSSHDMzW0vqcGfSVDKcbh0X7SqWF8og5YlXBFT5QDMOBs56zfGn
IICkVBqWS9u3ms+FhaWXqzf14Tzb+TAoJptxypPGymOXHODJwdDzKlP5y1uoyac9
xwCEq6/D3Tvjc4F97WuhJ84l287Wb2nkgX9UItoonwL+5EGgYu56oZcXkvn5zurg
i4gefpH3Tors7dBrKdp0QMX0SkyjnA0cmTkOKYn9kZDSALe7AfV/aEU3fhIJUMjV
/qataoPqTtO1n/pircLLLen7CwVHSh8+9+FDJrF6i2joE+aTYr3pXt/3//zPuLBL
5UJYqhpwjlEzvTOiNXVcbIxBOZJVuN8NDgV0DKLXna0WGZcqteuGwjz6m6nLB5iZ
aggOpnLQD/6fmL8h/oMADUs1mRgV7a8EedtCQkrbcJolHtqkrWThvmB6UgCFTp5X
Faj1bLDBGpHL2g52URZtJSvSn4sz+bsD7c6xf+g4U+4uT0r21Nm9SjdVYzM9de5c
uxyBICqIKn43x76b/+Qw9OEDACicd8Hvn/sngpY+zW8EeChGMEyXQ5vWM25KfKnw
piJa1invizGzYtXvWaaLrdpsM9Nz7Y/EqxszeMOzkrTvDsEh2ww9SgNS0d0hBrj4
CSIyM0nQCYta0dlASgdNkY/OdpJr8qENxPYmAdGtYZxLxHahN+nizJGgPZCdh3lc
q9CXGNindcJIO1ZHqXgUefW7kxTAg+TPU+/IH6Hj25gMqwa7bZ6vyHLZhMYxp1fh
XUOFCUfQ/9JIhJWbovba9VoqMlnt78/2vr9luvB8UVMyVPsOResyCAZlwDicarcj
eqa+AUJe/fYgdt02OioKqOub38NdsKz3quzdc3//gMznJTiK72XSkaHN8+3x6oMc
h0CXedhqWixu9XSp4xzm0Ik2Asz8PV1MS0Be1Wg8DgXvuIdj1aAC84jHV/PnzT2A
QuxBenYOeKsBOKuvc0WI6LvmUTLWOzqlubJ1MDBHhNpHj56HiwKmISBimIYIP6l9
M5AIAhkoZgxMhr7x5XHVv8FJkxhXZtlbctquFdkh91wmqG/ikSdAPRx8/24k6aJ+
odD4VefWqKqfK7oiCyvYHKG0yIXwaBoGDMTTt7R6nGRglhbFKD8fRzNGTX/dKvWA
ft4RYKdI/hZbZFxlAdGEG6x11lKOfNKY19wjk5WKQOVpHrgxwdiUnEAYHl8uR1Is
H/PDzO8HPcQwpSQZu+ZBpLiaC+Xwyjalp3+mx8DnARzNqc7tV3/Ptv/KsJn9pZEe
bqDA0r5f3ADHVSjwBMNcNmesS3WWVGvuGL/F2ztM5yk885VZxY/Y2jkDzOsamBYz
yKNomW6pV4Ui9aZ1/Fxu8/j44lpKQHsFQOT5uMu9F9HoGvH21a+MPsLs43HZp2ek
AyPg7e3Vt1PgBZBQ56vfv+7YQlBq6xoeZmicbeODvjCSN8AFEuCWpKBmSsm4b60n
2ivSIyNf9VTa0QVk2iOE0/sP3ljftV+E/9upZrnVO2F1BLcx3Md9wPM0NoJKeeka
opL1DD1fexk1TR2JZe4chofBmpHquXof0EdqyprZVqrL/cwYc5u/IhzacKxFa7El
r6zVv8LICfl5OfyLJlF23BpTaMF0Yub5TUWtEXEWFKI5Xu84iv2Xv51IdTrczLN1
Cc2twc7vC+fkLVA1meULM0HTh7+RcI56EhAVzNjkFfbKFzgCUdIxzGtKz3RWamlV
LEXg1Z9Tl9XiWa5aXqBYWr+ijDK+ffexDdXkfBsRDJQyXGIIVWxJKEir+bMvG5f8
3GI9F9dfcWjGol6IydGdm3nEUzB2cpcJ24AW3HlgZnZiz/LVSTI9MCJ8uSy1oN5S
6bee9GhNDDBeXRWTpLz5r+3Qrq+Tix8/Nb2h3+E2N1UWfXMtQ1kNfvqQMfqt5FX2
ryNx3g3eb3SPOkc0F+hr0wIvbfVMopXWT/Y/cWNXNaZXm6FxMry83abPZTnX0KMu
RixHqmUH4yLK6GP00OWWZcuXD8d60oTnOaysanDed5bB6AXu+Q6C0Zm2hy5Y/LAp
cCX+tnSZMoLOkxpPPzvtk/rksiYmOmlKHlIxYYR7k5iLDMioYHccedv+91Da0Sd6
Lc3ZlHYNoYD6epEOBiQVZ9tclDVCH2fDSzPwsxAq6ThWavpUa9piXSstTSR2ZFHY
x90eptWrPlvnxZGZDbLOimk1tIT27m1kfm14ST1rYYXVcrWMgRIOW5ad1oGuRR4W
jmx4nvUOU8SygICPJNR3RB/PMi8PVvnY+B2WdwREKIwauHmSMG6+8ydtXJlqf2J3
RdyWVs4AHgS2qLOQ9fJ7pViXqvVdAMUfaVhap822aOwyEHYONBapyRE8sUdNup5k
+b25uGAUhkDyxWVLqV1I+3hArTaX4iE0HFd2HNqd8x6oq4Wx1OqtbrtVwntCALri
ecNVOOlmD33JldHZBHCQr7Yr1aaVr4rueviflVL5EaPZSy0dWsPmar7JMkaYu9vF
uC64rGzvWEtK9FEXZ6+Dr3QBcdOnlXvsDpz7p/lDGbumcu/s7ppVolQZ0HIc75Rq
MxHeOzxyGvhQG5cxJ2NHcWAqbMDTij5IWEmsMq9qO4BD3HKIu7Yd280j7pf2vDqi
an91y/nbhHMg3pdt3ZYAm60LgAk/xcfDe0z+XR/IkVPM5NADnHzb/IJQYqKGNIWH
xlJqcsnslPdJfgeP49Sdgocsvq/dDxw8GGf1jUm/IoDDL1yoq3Whnf2Lrqn2xbiD
i0Ko7AuTkxfDHQlgaUoepi+HcVBCRQutNeJkRYNlSa47zT9H7rkGK5xsgp6IX3pY
VCkgGlwL6YUwCcyBK8uQHE268s6MPix+WifJDk3/D92TOMnPWfDLXbpkCWIEHrdX
FsdXvbalBHvgOc9dzccemBqgA14tralwDTsawUsWDVYddkgz4oG3KvohZmjjrNvH
2zEQ8l18GMzcSBkwYtNkeVLIYyDF4sBE7k0oQLw9bU95DscfXJyKVMq03PtfDvCD
9kpmqEvs7oA1w5lXT03GvNPIbGJJshBp+LM8xv2V7nlWYWz7VP5Gtj5EUuIUD8xp
biSQJctP+bieP+Zvun+Eo99CT9xmIanHopJ4hsJsn1WIZGLD5ZdNQccA9gRMoUD7
7wvYp1dFFdmfQuPNTKpY+m+KM4VPfWkmp+wXQ27bX+INyr6njdb4+K6NNffPsrD5
nm9gtIn6EauJ7/wEg+qTgMe85RnsVvOSY03qF9cltyMvZvK7VANSUSNW/Juifwz4
QyDdk4Mf2dPNSq9l7Y608wdYCG1r80hs9jiXtpQIolrocifqXVzPDwSXo5MP0yAC
w3oa3VSlJc0ELCzrdubgLIw7HbL++iYBcQJ/uPR/mO1QLquga9ZcKAjuH6pCtfXS
aWdv7tMv8iSQ3LV/j53YnIURT0h1knSxGZqS9UP5oWZ0B9x0R7ZrLmkPcC7AV3Br
zvdKTXqOTrGX0cRlRs61naJqWWOPck2CAAN9teQhJXg/hGtIyvnAYSYQ0UvFPVl1
Ucrg+QH/6tvpOUGd6W4Di5u6O9mNZOTXWpC8/F7gxT+SBzBr3mGcy7yunQKgr13h
tMeYVVoVstzPlHFScJBr95sqrZiRyIIQaqX6HSQ7mTml1blEJvLF4tB9d2Tf7+kt
cNB3TppewzAxO9FrfWJTYI8AQ8c/VwOdXHmztWxFH0tGCjV+was2GDr+UPWQx33r
EHoo2fs45hYlsf5P0pS7IxbDLbjxs90gGwCZRrlHz+ZIe2c2BIgs1nNQ2tSHKtrs
48P/3PY4zS8MytsESPNKXeO2Up1V+99XKALt65d9bTxTHffBltkwqXE4LQpeULkt
VZV41GKBx8W+9uVPssN7UMadfRwmZpfdszT6yBCjiBUCsIlZ4NI9mRHmZJTqqsPY
ArVIduINpF1ymxA164ICbPQ0VyE6AjpXOerD3QRuJpkM+gwWXq4OhIE+i36VhYsm
o490t0I3eytcDr6kFI94Y7ymGhqT1o5Ke4Nue0Jozk8X47T0F4uk0v2kfTyxW8bI
cOQJL882oINWSKOFRjUTZrQHtllad5V+kTn23nHgoo/T8aU47Us85+zV8pmJ3sYl
TKsqUZHsO0oYznRO56rmWWOcPSRaBVYLjCy2snvKCnIQ6xgMjUB/DZVQjl4befoT
glQH/+nFmS+YVYAVBO3vjmKaYkuCA94DmGakZVHYcXfj4F6VTWZe/IRXXEvclnyp
O8vd2MB4qNvuemZ72PXAHUrevgPbfzjX9S7YcU8ihtnqZ9Pv+jYDRLAdKH7sd7eX
I4/p/YkZ6yOpoDLQpHKvggK4n9x7DOXmKMSCqSMKc7FTVDVssQ25SkNu3iARd99O
2WWpjW/69Cf3G67MucCk7ey+0HR7mrgz+oZpjTrCWhkD/Y6SCGeicXi3lYycXOV9
f78wmEEBVjv/v0r60hjsjIBtg+BfrURdTZXCane6vKn1SaegIfk8xGUHHOT7ZJj4
0tBhlPClRaDv9GlkOyg6rdrK09eHyqLsevfupQcueK3CmmHj7F5x0pf549ap/1Y9
eoT5JY0ZYKuH0lh1jM9fE9Lp4bFg3SXJBWAiYXrfEuhtOm5S+zrHGYjtlqIdocQU
U7ivRJlOEFeKG0kY5cs+2TbCvm+hHBMfGzygUJSKW+1EtALtwhzAiPvD8Nk50rzu
VzCpb3Eo5g2QAC3nhNa5gN5P0M0+ulfVtuTGuoxr2os9aMZPte5zMwoFLsAk+7FD
HlsTMsMCy2Ti5tyIkVgCYhqLVpqqfjGeynGPrK4AfS7hc3sMu02NNEQlnB8+c2tZ
Rml9ewi6ujvfmbOHzGQoX9J4cOU+BMSU/fd5APQBF47LPkB40nfsgV4BCzToY2c9
v5fG4b0tFh9USeR12LZWZzKpaCv14gqEQtLSQoEUOxhYw5QVYrrSXzphwRrMEUTU
Zc7VDYpdePZhSl5vQQFyhRPNDFZWFpWxgqoqQx3V/kdcikzFo4sFGEtCCglMuVhk
lowiHuNBklqbN/FeK+pFbiaAMfmAI8EcDyRzCiSC315SAbdWlgifW0T2sSHuDRIp
QXAI2ymLpTylGYWHZlZhDi8zQ0CKQZ6SxpIn0kQ8npSXYrBm4uo1EplceXEpvoi/
9h21llB9bIWbUtvLnKOuAs2VWHK0ywTjZG+qYFk4t9rG6ufQP4iOQjzqiLNnQk8g
0wH5Ng4M0FHh2XpyHc37VGIVgUZ91H6chiKgPRImQzOS/9S3zQ1D9xyQTI3bmrB1
is/e+fmK95uM0XgnzxWZP7U6hhpq1fz3NqWJc2b6pUNq1TiGILgxYB8AbNl1Ju/3
eD7lOyUdEqATMqMM7qtr4Q2KKPaQULmaoHY8MWslaP3D/4lNFmwddTdjV53S/gjw
hpAiT38EuFohKqluHMzUZDZVf4vR9TFciqrDd7R60jwdwnrSWlnrZn8Diw2jaTgi
QlEzzfFibluXV+E3qcoLazuaf9YKxOmy9b2AM+FFx3CkV3rRzExmDJJKpCMh/gME
vkZeaMeQThHiRFIucj36478za818yh0IKxhuOSp1rphZ0ocgLuAuBcALQQpagWz8
DpF/0gcg5GM1jOrX6JSP4yo/AKOrkocVnSTQ2gQ3N5QkhCjgZMnW6HlHuahBKY8R
VhJsUbTQy5au0/Ul4jJ6Ef8vutqCTyfxhwU2PXb0CyHHqtI8/A7978c8qzHiUeLt
p8fcjcOI++xPeI0YB73xOVuyzNPR9BfplRKRZgS5Qli+pGZeW3hXB6/V4c3It8Wv
KfJtCAl9SEals8WinEDndfMXhtwIaK6KolqL8PjAZFYq105die7abjP9eGtfWITb
12tHvDeN6rkbyg9ehvthT63ZqGgGdjmdztvRFnRUR3vODbWvji4VwY/CKJbvQuBb
2R7sidQBUXVjUXAXyZbH1KfNM4k6zWUQxu3dmpMnELS47fbwZAHEgJHZPaN/d4DF
ZuxfCPoZaWBf4b+JuJAK8Me297uqmUubVCn/6w4K8XMcfE22EOR00MsYQmjhEM8+
F34MDVLdW+NoUxPbwWsxxJjqv9XAgsIKXlRZz7N+nCkNpFqJrlaZqRa2LuA5JfGl
vQsf3CuURu5RqgOaAYanPRXLq79Az+kJLyOMP3KtFFBxTK3dyoAO7WhmPV2nlTrR
rbxBon3F5JrUGZcSxbmILafPMEec89ET2piQptrBFhQJszY725siYwIDUuTaVS2z
KKKKE4+Ge48WYX4UipHK0T/QrawTr+XzHm4h77Cehgf0Du3aliIpm0MqSMTgOkFh
NxDOB6hQPFkmUxHah7dem0turZIN8nwGWcasxHIt9lOvF6qhwlH1Qd9TSD1zkvfA
BXr0wLoFYF9/oViAd/qQU3vKe2z6C9cTosEJhyGgtDsSKl2yWSrVCv3gfup45Qm0
gr9NJuE1N3qkpjcI+g1ljJQMIIDSjvD+QyWPsTgN4xvkjhyolc2O4r8X7AY51HbM
2gDR6+UNqs99yMQaKAx+vg/BwjyPXq8qEc9GdAeijXbytHn23abn5Cb3n4S00xaI
Ea4Q098Sop3lB/1NlIVJTSqsS78vzBAkHM6rA5zGVHNJHKnmLmmpGVPO7R9WjVnB
wdpL4WpSFStB3blPXRxJg5ZyOcGn/Z8YhDFmigYOhWQgoE6Ljh6BKU/7KAAuDe15
RPX4asxGoXJecdaetlD07C8C5ldCohOpkJ7iLxzYVU8Zz2fFpCHmhwsLd11yxP5u
GyG9oF74jd02osMAXO2ChhXuLd53U3quvAvkwu0ilseCrFfF+qHK+0zf76AOo8IH
gSqMklJAo1gUAXdRimxwObOoCD+dGH+xVzAo0h/WYjKtO10Y4nfCGFFjPC0zvV4L
SQZFbaGh9XaXRECVuYJQ09U/uFoYIDOz/7PLUM5w/5caUlU/twZ+OgmlZh17RxbV
2GIIyU3f5JUvjG+0hgwR/nsxcgTUuk24g4tKCFL+NVGmjJ8o738vDQUL6AmUU59w
UNBvevFc6FdDRHgOxZQhZ/BXUDbbGwLp3zfUTfm+MMBGRbbyoeqCwtbiQHzVf1vH
8V3tZqdixT6Gvdu6caihQzrGeaaMPLHhiN3M3nHPLZ2rjpLLBWJWwIUoIg6watq/
SawPSUE8vBrErLrJvbz51Y+Vyixykds466OaesebC2tbXdHYfgVH+L4QFbcsRaJB
xtEZYPe9NN/Dkf6mtDUvMVfkyPLv5Exi8CK//8U6s8rpC8i8fz3N0Co+8zKVxLek
gru2OtzoO8yxc/F+D+Y/U38u+WBFvqhGu7N5Ly74BUDPlT/aruFwee1emurj7OJv
Fu8z2Imx31aR7I5vWMwK24g+v66ad99pGzsJDUu9DAYnAbsvjIcY8cv53imf8l8E
nukBsABC6W4zPiwRBN5t52lmWBIgCcdKtK5pLoy3/MrLcCROyQiqIb0mD5XcUxFk
MFp3yrNOQGcqsCfvBJ8jqFgX9xMYxjZXXZurSkKiiYK4cmnqfuSgtWM1WQ84z+Vq
1k/T+MMfK2dRxVYn2s0enIqs9/umnS1hRqJC0Z78GFsUB7gZVaxYeX3VwSBgE6DL
VPaMUP/10otuGFgnoSPrvAH7GwYDb9lYb/oqyL3KLBASdCj88PQMMQG037GEqeE4
ZI9sJjQGl3/P5CWVxKkBTG7ifGaDUyEIhgj1D5InJ4o+iBBWo+iLEAxRlGP6Ep+X
jj10CWV7TFzXZRTeyuF0CMHRnpE8VMnZl+T2RfRv0LA7Mw7UyxZUkaeU4lxIrBbb
TPW2XjwObkjakLucmolzPSUtV534Cz6gNqpczb6MIkKZa0G09ubG/yNTzl/r6jiq
dhaQpG4EyXLZ6DnJKFO3BjrEcityEpstbZ4LhQvG3i6XwfNSZuiL3OfCLOOc8GIB
cVI7F3TbvZh9PDWPDs4etJwOjDrbMaJ5kIH5tjBXvif+VuW6YLiw2k0YIQhgeyLH
YwLl9SRkN1VIirsND6zex7mAtWw8PzYPGlByzuUYIpjLaCUMaH0F8JtpV0+WxYt5
n9cGXHoxgU1fSotdnDSs2BFBnWObPh58bc5VERIwKuM8qCm2tBB9TU1vBA+VqILE
7W5nnmpiw2on3C494kTQKmHdSZRdtK7UjCT+pUxuhnctogh6eA3PXVST/uC61hml
0oynRM052kDWuVjQ4sQFDb6WeJFlF3xyuqsoJMQfK/j426SwF5lvfwetZM3wWP4J
QUojlOL2G/Sk65+UyN9KVRw9a5gxb/di8w0XE9SYeSWYEpcNDCgowJXAJ34eTEKE
WbHC07npe+YuZkDqLY34tD0lema1T4oDFVBl7MAHlDtB7E1hZVP3PamT84tDCIQV
xqOgYfMwyGNdkJOlFhmQ7XWOw+xnj5mLzznQaL0jDgWwIFaC0pHJoDrtBQkrohwe
Et8I/KxrtqOnwYQXH999asuTLmFnzsBdQd4ZqHKX3zNeMBldLNnWBfR1+gTHnLsM
R4eYnsUpN5n+RH+ECDq3ZgkG+UhzFKh9+qx7fOMeoAeYvWIAaHFJkqsoZl5ePc2a
Ujez0NPu5cU6iCGvYpJAwTEfTVIAvSE7mCKoZXa9KYnvC53q5nPc+Uw1m1WmOljr
SpQPnUVudTagqqIJiwvQBYu5Bn9pXGV6IMgTPaPmvkCdJHXPf6bz7hhvE/0DsAyL
Li0FG98cCB84EVznW8/q1nqLURcTkDFuA9xH1fdRmptUN+x9kAzLARPHV9CzLYvh
ym2B1mlzGsvhCMDyq8Sp+2OjfasTTQepO2EGjWrpKS9VRKjH4+VOMMlO0YY1a68I
oFC9kAWuEKIJjzC/qklcIg+OkOEF1EFOedG+aYSjwvxIx0FdkgM/2wLp8s07GOKO
Og49DLaGi4iZiNcywfW2hSdjbA30LY/m3t13RyeCEIopsugQmZhEghEvMPYIF/qh
1wJKgwaIOvEHjFZxxJCmnxeZ2+IAfMcbCKA52ZNmBWmrUcjo1Juf/jdblS8WtysT
OAJVYmhJ+xBHuXlX2MlCAY09t+5bMazJxB7l11WJLdV9O2rW/ow9IDX4t+kszNgi
TsaM3+bRcrniqbZZ035C620Mu0vt313jebFW4folNnmWrK1JNaCZSMvplggxMzz0
R7CODRiTZvg6l6GAtrrupQMXNlTr9FsPWXjuqmPbrJAVAQn1aHVwU92bQ7QDC+cZ
M6pD4SI5VjyywA9MSpxJYpqt7qTu7VqHg4u7cM/V5sMRZyTYAX3ZUeZmN+yQJFFB
ONd9+bWYo6q5jqGSP7tkCpYncpEC+E+5iLv5jyOV0i+UZx7wvRR5sTjjT6snP02M
uW+oqpQIhCj0KaXUrWGuRkq3JkfKxoO+eJmwQxON2WXq9oWRntQKf1x+g6HJW1in
eX6RpLtVknM/DJJ/vstIN6NuVsp9LXxAaXac/qE7UhKJXKGAEF2KHNmLpHbqVnjK
F5iOd8ylszW6UJvsqbGdwljQSIWQzhjn2bEQlYIc4ew7BMv7M9nB3R0DA4iP5I1k
2qFdlWqyrLc7Az1kYP7oEF+h9fiqlcFl01UByVOLhQP62I+PwD2d8eKgKwsYrp9D
FfS9XC8ErtuAXG0TpdX53X/3pPseDstzOywKaYDVJql7pwxCfUB5NCugm+277Hn8
FZb7EyWCV5/2WUOn8Hh9hYQZ27Pxqdu8su8AvgoNtOm951O4s/ARF19iODbFzmYT
tg31F5P9RhRS9BS5VFrWxGEkFPXmQKamOM1Ys+GsIuiHYs1qId8EEe0vnxZM/qlX
K16LjaZIZuaaDjlNOp2WuLs4YKVTnRP+F+qwCSeDGgPi1H4hE6w2LlcSkH+saveI
pWxjfiuzCtEz1/GKNcTfABwEihwifUbmN1vp6Be9T/BmL9CTDQhSJvgkmJA1AEKI
hqDUdtRAoWNnM5rNRmYBUPZEPN0SObxjrgd7WbGq0RqCZZD6SzVI5/2rLHripacz
ciIbgB3hUq0BLaP4n8t5yFUoyZXisHfc10jGSG1l0CyqKPd4PKLw/ZuKDL+390LY
2EiwJDNZpXUrwXq67rf+SUh+WbZ5WGTQui+FH3Nxc2HOtyDfCRsHNswdg8AOfvCH
M9VRlxYiobjFOzf6+lpRDLrF3BVueu2BPDjVZ5yXcPo5L54+J6BqVUXb6CwBBsEc
AiIDorgI4FMC+Kvl28JcU9eanEjdGh0vBvZktVByCew+w9q34tR+adTV5lkG3Tv8
y26BoztPh730Dv63oVFz5Z0VNL4TVP768fzTpHLamrAg+4iKsCX5p0TMwPnaqxZB
gCICHxFwkXUfS0yOBFySyAZvyE5LVN3YIaJdwURzUuQ5ugoyTXLi2a5hYoVbb7/v
yk7WSVXbK7RsLHTjbVyI225aGf0HXGJfUV7n8ThFRe3VCD64x8V+yrY/gdMUriBJ
MbUZbY0FO86KKipd3HkLYqRzvCgDgLI+fFd29uMRYdAcwAZkEO0m14bNeRN3kwqi
4m5gT6dzsTElMc/RwhW16BE/P9IvkV+sqDoOh/mKMjnRkjuwLrMXdJFRLO6nWQ2b
1msGt9Vl8z6nrV+ljcLnnOMfjN4fjM0s0pSEM+JTIYZVr6wzSFsFcAAw9FDL/k/i
HF5/8l896xBJxkKn3v94qrpty02NUEG49nxH8aSQ3+DIo6XtJMYdQYA0+UBxsS1I
VyCvK8p2EITuIgF1I24v1BN8lg7slIJeWRJutruJo4iYfbHylyJaFqGoVFJ+M8R/
Kn23i4VPv6DCNU3cmIfBrYZAyX2ujHmCUTp90Clz8pESX9MhdGRMnObCOISeZBmd
UNrEtfrgUQ/74MjyYgFgGwuG6YqJq4dStip3jGwQxXxnqbxuGjLHz8QoDjYY0Huo
s73UHtLQxqk5dU8T+5znSZ3n9jIz3J03GkUfYb5mDkeIZHSSVJkD4rQFqW0B0kLL
mVuwOywhvid0O/Jb0zu7y1V4KdwPFJbY36d28TAP6NunIS588VP6Lc0XEh0URY9F
1BnwrM63PFVEQ3IxM6PxI8iHhUqU7mFD2Hnj0Bu0Alh0QWSQNf/WsrUbdRhoK0/B
BM0f7UekFaMpRFEIDVA3Wjkd09tYYgyHZRzXuAwyU8P83UJoyc7PAz76TstYQ9ml
rsmlk4svmPRTN1eL1BB7Y/A3w9cwdLmeCcRdVFAWa8VRin+1ffqLrx4cX3B67FZ7
kNvCd9xr6Vm99WX/5v/UpMzAIPoYfwz+bsfbUCGw2zKvzO9WkkyJSpr3molSzvqt
P+vW/NwSq+QxYbZJA0mJTItL5Am40+L1udGFL+h4/DqYC9KY3FnUopDlc02SiW2c
v/cjt59pMyhYUMNn8CVPOFEqsC6IAd70g/LAoMcnQnDprfFSOccn93xLtjKumuPU
pILAOrBYE2aJlullkKwZK7jKVOIuYUNmL0oeF6D+0jUNcDd4otgQR8mnDywoBU/D
UqeWLw6YXPWfD6e5WxWFpcjTTZWlqIsVpmsNkSeWfTh0hBMlvIkFIcXKX2/vTy2V
q+FfEHURK1s0IJjF+jkcu0sL7YvxxBySEuvzecd9ray8S0xsjFT0hmRfyCvmTnbO
RvxHctgX3dR4Jj8Ry3THg8WYrMy8+BjxceLI3OVUbLdJMPhGJ6tqF5B9nbpnuHPr
Db6R0kXcce3fquk8Wo2e4lTxgcXyoatA0DH/I5bqM6W6/RI3aU4j7QbbSnBuXqgx
LMfy9uC6EbV61aT5+z2PL9XdkZSc3rhrwQmw7s0zjnQm1TUWJq0dtRO07aUfMlzF
HrktlqhWgCp96Wzn/45E/8G1sZqlwZL0tcBZbC3JxUy3Np0/WB5l6OmL7UyHYzfJ
1zNwFrPgwFWEn/VZ1C6vNljkByC9EplJTG/Y/Q7GidV/copZ4YkWgBM6Qs1A15W2
hIVSIqGBPrHGh6v26iigHJ1HVEu9A/p++3O9VVCz85MeQzitEcI8ClBGHMRpBC+O
zipZ5zLx9Bh0Jq0tL3x344ys+z4Gyu5m+wKlHc3X+CttpCCxA7gYIiJqJJHyuU2Z
XIb5B3OPSIS8jGr6z2eLpVpOdaoBNgxt7gv7aG+7AiN3gLnKNEOky9qI3CbZ5Zz3
k7hwWuvl8DUuYKuMF7rWaNx1QW99v28OSJmZsek/UhCYCVcd1y6BMejQxau/nAsw
lVzf2Kf4h3Xi/eu5fdlKKOBBw65ruP3dSBt9BkwO642n0CCE/UT+3KfGxcO/TZRn
t+WnuFX+vKsHLKEKaxiHTX/WDHJ3NstV5b4vSH17gV/ELYunFlIhZA84ko1zgx68
85tCW/ijjAikLrsKgY6QM5QpHKFmAK+h+Ky/9sNuFhWWUSnHY0QbxBx56OJ+llZx
hTWwQ4csNMMhAzH+NMkFsbyYl4O688QLk5+PHf3+xVgMuWIslaEttTzo0j/9zg2+
jKbK5edKCKvyy7uZSviyk/Noi5SFWkMiOZ6zkSDrcTV5MgwvORnS6KjgMyp+QIAG
NqK4e57/6vJ39a2yTcPMDf6xqNhIXYHVMsFdDV2AgLuSfulYy8nd+VExOu6AI/Fi
Bavjcq7BkyoYRrE0etCg2Q5dW0qRiuc6cGj+ZlOO4U56a4ztdWxpvsHz7QSWwAAk
zQswPsqjMJyf8UTSpATuzJ9Ch2wePGXgifPtNuNaidWMhhNC+eMyADQ1wDezGt/R
DR5sg9acTX1gph8syw+tqzt/Os7d/uut0jLAqDDyyF888mOwXNQWogHEsbVdPpxl
/bYHDRGJcgg/DTbZ6Hkmjte22Y3c/0KKTXjxBp/ze1P2pwDTAAYf8gtRid0e3Amz
+ex5Hi1MAItuoDZrFQGfCuR3chNcly6X3ytjlLbjXKbnWz7ncgcQ+RyATjUidwCo
A4YccdK25RghLPN6fe/L7UnroSUywofvpnBNK5VoeO9IPVVQWYtiO/NWvMrpmYym
Ito4tOB8C4JVsfxOPQH6P78qr9xRL4EzjDCK62aszC/C3DwBIk4JKbXA4eo2pWEE
5b/LSmDH3x/2jPm4SuDiiftDBIUiwAjsn9jnZ8frAJLJYE5Fm2cjqP/Oh7fmMLHH
E0Zh5HYcPBPJEqj+sn481eArangIiWL60dt5QTp0e2M71N5tVOhXhjyWnpWSfPUn
eljYHxGLXsGxLiai+kBrReWfG+7GbEJGOVzYr2j6n5rXkc4R5eiwr/hJYez655gq
x77KYAcZ10ByQL54i67j8fJXCsw40iHgjNfkn14vivu8xplPcE+pTblxqC44MMS0
lNJDtTnucsofuqyrm/tvU5Hsu2VSXfGbmLH6VrXxciYOMPW0Q9fFInW82pc9zt/X
3MPIfZtZxXA72XmeSgtk/k43y35sr3ulBPS3e3PNsGfgIGqT4IpCbRoyArxG2qKP
09byGnM+/aYWgXURLNaTqo/asLDD8f2yZqLiefJalOCpAFW23JyY18G4jXrlA/GR
AbFOvLoAcfgUaiCii83Fq9yaVg97MKvvyQWNB1FdjALjKztpbd71GaTbPkRczb//
x9AW1JcAhoOyzMIGmN2ZxQ66R4FhVf7YNVh94QoZtVGSUvCN+6kTo1sqlOMuK4Ys
wzNvFTuFPRKRN9qKiV0T/32k3laSlhCy29QI0amt1Rfo+0N0Ap6abBKpFx2Yr2Vw
efbAqZHp1RVMD/SlfdEwsegT5VbV902/qWCpGEg7tneYW20MGe0MgWlXxgdM2UG9
kJPlfQMMkMYqOPX8GvYm+8kNL0MuRLG1MNqx4PfLNmPWR+hBhqao/3D0NW3nD6Jq
gO8+Q7cYnnKnjSMwmaMTLTBi1jILwIzdKwBzil13J0SO2/DkhWHNR6h+hpWlwZoC
c1NeZgYpkZtUY52QjHEu9L+aTK+ddbon+wysYqvjndpCQghZBtLxBNq0YdrnDCSP
jm/JVLiHjMfHPvm51tt2+hR3N3teQ468hYtRyr3rVrqDZvYCiblidLJbLaXRtZPs
/inOzSZasrYHJ2aQE4coh/xKvANTUzYEJhNupjJUpf9LTYhokB3Nu0Tft/YmYnsv
xn4PUzYH/jSkQOHzPzdQ3pH6FjCmqcvnOZex/kHASrtOu+p3XJ7AQJoD2JTByiFq
/hNdCASrIIk/9Kb+CByjrI8oCfw9hP5vymOVLEpmSMkmAIEj6HcM6aHQn9zIMiY4
DXURYT5eQ10LsLx6Hkq1EUGwIfX9v+eibXZWBJHq3A6IKSt3VTkYFgfmnu+oW3Lu
+oDrtnAuxBVZ2/swiMWyqy5izxT9BYhmi52V+cjR82QDQupsRfJFXBIwow6BE/sv
wO0HaqnhtrtT0adlMjtkmVHKkXhdZrblzS8sMlJBs9xVy+MdpxG1e2uWDXeB2zi3
a3AKiuD01KdyMyCRuUzJXC34Rgik9pj0iLWQvYyptTgFJX1tFuz3WYPw7Cp1tqp/
vlPjqBIs5PqKQBNXNOJTyT6U8jh4KqH7zKDdgU2CeNswZ+SMzSxmtzdq4Z9bi0w0
fMMMBgENwmittKFc1A2LdCXsflCZdXbGO/DX5HxDcVPt3jmfza5wLnKhkIxUonqz
MlNuNwbTSQvusz83cdmrD2u1yJYhHuhMsG7HztCVPAU+50kMcKlXf8AN7P3SX5dE
Zgvv1zN1EvE4IHJHX/PCcHywAX6ehDXnp9snaavJyvqfq9gHXPULiU/TsId7B+zH
TPMOn55LZW4fIRinZfJI2+S3e+qbrStsXaJXjF93yww41ki1roB9efHO3XHyuYEo
w+ZKMacBmlv7fuHf/kubQqiyHDdWw99q8kzW8JWXERnHFI/EAF1JwJ2Z6URwlsWM
0zcPPUFGOVTvKvhkmJSFXHpMHcRSlL2inSnlMGtfk17dP/1PZYrCEZ5rX0+z/S3M
AlufwVws6Eylat3CKnBSRvv8/2V7uK4JbSWypWz1DoSZ67mr8mI0k4nLZR2pNszq
VjWdfygN5uJxgjTFPwrEMwlOblmeEJJIo5UzCF7opbK18Alzg4vs0tuCtp9JZgxA
fkusXBN3ffrVE+vcn8gKgtlJyDJEwvJf/w1OTFEaDVAYgiCXPpuwUfn4sfBc5Ycy
bEJ+AdvWEBynG027c/0CIByN26UmO3pVZC+sF8qgt63cKghcgUu6ZNjZJzQXlDbi
5lnaO1ABpto++PbERI7UUqau+ILQcr7taWxmgqiQ+HTqdgJFzbGf3YLU6ifcuzqL
E0whR8XDN1oLCIqZuJH738SsTbU8q7lbGKZi9JHRcgZVH/gmeckn369sycaCLueZ
aDezVwCHj7nZjBobkcTN4FqF3NEL+PlZs6LufE015jK8UW3kJec0njKhpuBIYLrc
vBHUGzvFwpIdfZdUZP4rBZKgO2TXaDhfW/18ry9fVeNR1BzLXD2mtaLI2Qv5zzA6
I1Kp69HCo7ilEgeaIN13kF0pA5wofGtidQ5zv0kY1BXW6vs+WM8DXjdD4oap2ngA
1goCHqNy4cXPbPILweNsa42cLg2kVhApBTQuyV+KNJjcukhMbvVY5UqPmkFFdgFG
FBygCCiLJzmn7Df+O9PTHRkVAYcd53bVtjgotVqnSlywpDSpnXPWQPGm1fkD3wV5
POQUJCn5Yh/n6jmdM1NCIU6GQ870C/OdVKWWkNxQFoqsXR9Vbx6nCo/42PPXkDee
TLwY5OzVPkDTJmvke3ICmjlCYs3Gwti2Rykx5PLwyMZ6wLm/m7NE6Hux7P4RFZQO
TdkAhld/SGRfFwyKZBCu6iHGqEBjbtJAbMO+6XO5pdq9amaWeQ/OCFfXu+QnAXXS
10cC32Sk9JqA1IWFssddonq13Qdm0NpdVo6mLK0Ay0AuJ7uzMi/u8eUpNEZw0vJr
DaXCq6RZ5vFGM0Spt91grXnOAWc0d4u9kwFM03whr6oYamvr2zTd/Cm9PD/az6UK
MMBu8BrDokxHpuRWv8Aejx01+xRydwCUEKA8Tptb5DluBs9F7FIznbq1iQcUJEKO
MV9aNBPqItYpwR7eLKf5+ZBgmTbvIcV4KQnYqBKJ3hwmPw0PMFsLkwcm5IHpJdVj
rbi8WYWihZMaebinjH9J3GjbMtfqAEFGCB4Soy9YdhPhpQlHKvzN+VxHkoyPqTP0
GYpJts0p4yVxTgERgMa2kmebJ2aztm57pwPWy93IwiLjDr/h0PQ6KLgA6/y+Bb5v
yqVkeuyThLcXGxIfehyJ9WLIHW7iQ2C+fJMnjD31uV5pw45d1EZhRDyugTyB5spx
JEkydAI1Y/0UveNvkbKs8Sol2X+8AJF9I9C3a9/KfUUThM6tXlQeEaDrrXyeV5XR
MaTEuATU1crBfJFiUzEDUqkvfpqNMz+3TBa56uadjPHXYek8tnKQstyYhw2ZjODa
1EHYmPpBzyD05okvTPqcQ/syq94OTMEWJ/KQOyfhD2f9JrChwntMDKEQDiuyn5Tj
uW08jmmZymoB4Jv8shJpK74oAIJeg5XD6UKQ6SGf2GozqK0L1SY9yLTwk/ZgoXJg
+irQFdLwdN+aY5LOFv/qvjLM62fglQ0dKPgeFq4cSCbYwAOHDeu7nl6IyTYMEZWy
OX62tKFoHE8zkmr9bdgnSIyk4bexpjodqz3y1VXhwRJiDtF+HMuhqku7wWBkdq0C
IJ7hIUeYHd88Pxy6Ove+8rWm6sFjiprhPCAjBvV1MUdfzzElReNiQmVku9ekcr25
aXA/Eciz6hu3swBoAjziFY2PbJVdFqIN46d+QU8BpV6Ym3zZAAyzFFxvD46bPej1
jpYtGr6wME2WwKVPZoc6Vt8PdFKYIv/iOBBxOTZRnDH0iekJztLOuDYWXFfBMkpx
AhK8PF4v4hytKeiiAMVaQXvDa6xTfrVPvffuLiNa4FaXpiVbFr+Hn7Nd6EznKWwS
xu5sHMw0duwVDnFPCAxBdsuvDnpCRq2COETenUmQFU91v9V+16veClM1skodCYlP
mbmXz5Cr7nPSqTkT/GBCUzgggVmEPPwdf/sEE9P4KubNrqiwe21I6IzAvXuIDxnZ
DYNBmV5A7XUq3HjMnkco+bySWOYek+Mel+2/SDhibkMNUbSPGb8ZS0yJyR0wejGe
OSFb9GnNymX6ReI6JNPIStjtvi78pCvRd5rY3z+0zjT5xTY1Hwr/TFHmiMk+YW8q
62SzDh7/Mbdg/Nt3J17UO3rdZvvh4GX8rRpQiSrMXsFM2lA/LhCWi0lsyYX+vFqF
772gH7HLeaRRZn22kydW89ck5MgliO2JQxq+Anr6f6pS4X2e12SUevTxJLlBVjj6
SHuPLK5XMOPx92zbjlQmh9ONOvgR1gTLCkIsuFk1qecGoO7rSRrlfco6NAxaCosT
pznJH41/TIUuNvCmxBSXuX/2lSFfWLYnulgIxjC+Hb+2ChcHAlnNXMqrkSdYA8YC
aW5lZX8unZ5O33reJNT4ste+5JHqE7B3UqTwm86+rG224XKyuZByjKyD0/Xr4itw
+XFDbttoQtrAkHwJP1IeRJCKuw67I7nvo5zfOgvidt7RhxkPCVxTVGwyluuCccRV
DTvPleijxnwIPOcqVmAgQOxclxJJLTbzpvIP4Afag5l/z59/AQCzCfipkc27uEan
PJVz/iXq1EdAqdo8qbNc7Bok8Sn2Ua/sBE5R0rRoBi/AqOwW0kpxiqinzXti0glB
MNoDj/Qy/2RO3caDvnyLvw1st+JozRUaNopVQ3xXoI83abrTbcvAAu4xc34EMMGM
jTm+AEagtgGsQImsxf8+sERwxQfdcD9fMZOaZeggRv0IEekcq9gxs/Ehhz2YnS8e
8efSHfJkmJdKR3j3hNrrw8U/a3mGptoJiS9jT6P79898l+f5kv4MUMWZvXHgJ7Zl
RoAlEexyzTb7TRjRKfd1gXA58quqTMcuGCgeb7G3dPgXNqc4PGGgkgKG28W0stt+
m9XyhWETz/LiJD9rVyFzCdohJZvgDhT6uT83p9ZEEbCmimwgM52ExgOx2CxQTQv5
Bz2G+EzO/wxUGdcd0fW1mEf3T+rBjpvfKTcd179TU3UmVxIBJnYwXEpfsUwej7jv
+0R6v0uWpC9AF9lGNdVDTe/kXIJbnHkt2X1W9/AZ1kIpE3rVWdqL96cS3FbSffy0
jXRpgSKiOhYee3Ya67MvJearK3f9TAunBUB9lkHlfvMPXIXzUmQLfXUF4t5uipgR
97SLkYxrizbPoPoNx2/wgmIR52KPBJePVFdJj+Zw3xs2HY0cueRtrptBapl697jK
C1u+h1eBKqTsS85kxvllm9SKxnyZP+SX4cmVzMJY+5UPo/lLAbBpnZbx+9ZON/jp
pbW2Yxdx3cz1b1HtqlGfK/L5jYIE+2oZCnh8JzWOXvRlU+4VkHnvOClvqDmv3csP
NgUDjUX7s6TT/gbw1jcJr6PqRCWkPBfIzhsOZalVPuBdS4zuz3KIs3XaCvI7BTOy
ysRGXD13r2m9rxKPdLbVWjaZbVOqtk5tem3yPSr85KnWoZI9WJQR0pU2TFEMBhQ1
uQSnf5kb9Azkl6+0ssAnvn72Ju6FolhtR/FCvkMYufVTUkq5GsRou9gn6ZNZDez+
crujfLVDo47KwKAKI7GkLf91RaXxX4jxLcsVaXRdySARO4xVTVERXR+MGaXO09SP
twP1OJLXakXdvDsbhtDcRfthk69/EmdnXiNUfPLOKECoBM7d+dhTyPSpgATFhL8Z
pQuu8La67vDEJIGg0dtybApqegXaYOtMogP3PEqqhvnmN+6rnIC2nYMdtlGY+l2a
lE0W7XQ03NVgd9d95qG7YduaGsQm+uq//QLcNzyDUsp8coY9ElLmcS537o2m6kyl
LMi2L7HmHl5/nRHlmcBG+KpLhWyd+Cx2qonlfTJX28WZ3F/Qgijh+rnFzkf0pCrl
wJIfczjCoqodPj0emJQ0NGDTqjbt/9unNvKcyU8hiL1IvlANUWZAkJvNEKXnPSru
dv7keUukxLBb8Aa36dE/OydBx04BVlP+0GWrjR2CWfNF7X+/LZ3pe5kPy9TxXWsN
9YvxBveuczQVKB0pCWStY83B4vDQaWPG9XaZddYa9XxP0RtEV8ofVDxOOuGQXMBQ
VZJ44HnBBbL23u5BdVgY+kGcpQ392r9GYwftZDeWn6x2hIz16HmRntRRfZPpaZJ4
2be3eI0czhyAASt14I/sbjbjIopsvqBqIyyeBdO89hYwK0M3OenMpWkJ7N4TINUW
Kwr7Q9XC1H+L8U//y/lpBfFrjTTDngNeI+p/sk9UYGpob63eaBmXlx4PcDRcVdET
CpUXmSxoaAXEmE2crSd3h5xV8OMLQ5q4X+v6UJ/mUwMQroLvLIPyR39k+P51sPZj
1U5XutVWospnbRkpaFlV3GhwIAmloY9HMNZQV5OXxQfl+D0f284maXprq1ShUXxP
1KIJgtiuSS2RUVD05Q/uc8ZRdM21tVYMa/bnhnl/DWWL8v/bBAQXuUUgvnAFi72A
OnGIQl/kImmw6yA0dnOVRpRfjyQUJWDJGY2NjAEcGkfXJ8EnSPDpFQaACAkrqAmn
dhpw36qo3thriC4mJmHz0v3VTIDc+iRJqjV8mnwwdxWT/17EFOLPeKS/b10G4bQp
+xduFSskjXf1Rz8ab64GBWyMWPYFw3lqP4aekZXCotsbr+2EDGckEQ8cTT1o2f+r
gb2dqsdne/L3/4io8t0TBeNeJ9j/8mqLR/TjR/imvcwvat3yAMamFdxGsScjJdXt
lEuZDflfNV3LJg2OHzyIybd4t3ZQkOObG9usr9R6Oig0mmWks6/0ojbzHr9pWzQU
uh/G2mh8pgpSGhK4146LgIcVKJUM4PgfuM23L41TZCD2VJZxFOAMq0q+2Bjbl/og
YuyBOwKIFqfPgTs1JsdkaNoebDHZhhZayHPS4njNc4ZDIncazgeh6NTDE0ihvJ4a
hyue4nCA51HER/+bAnlrS/GnMqiqfqhJBEC0hlkDNz79Kx4A/kBatoKkxCVTvy8z
QSZcbwWdt44N3dL9ahhPkzg5X4mzU13SAdgLvmhvZjm/4it0K0bmho+xw1El8Dgq
FZyAykCQYvQbmd29qLafFH81t/VeMnxIZ/+vS1WQP49x43g9vLmz5bsfSADufWul
g0scIza+Eg+4R906TEPFW2UpDMJ+GgbexocE7RDDM/Uy5g8lyvy4w13AyNsVPK7M
e95a1Na2zASkzsaydgZoaaiK4FjtP4a1BuRAxgyYczBsZSM9sUCuipDZibSSY1e1
g7Pzc3Jhtr4mpb+p+fZ2Qb9pyGC4mwhS53z7IPN+R/oq0kUNPovCM5RtPIQ7M9RE
9qwopNaps4J4Yr2g1PPGtuov1+vkT/qcKssnqCjJcLr02bHeuN1GqVrnEWMqUEUL
4S3o8NxCP77r1j/bpSeJSkRiG9sTG/EKsddIy0xTtbdXyrKZ8tOC5k5yVQfuwQ5C
i3KD+oxrgXQtOUeiz6xcYGRJFo3pdVnmCZ76ikjEeurpowdx+RBMMcxVorBa+Wp4
VeffkG1p0QtWOQy1AGK8ihXyA6XAB8IbO2qxwVlMi3hqKCX8fC9PZJiDEuK0tqS6
trnSqUXgiZPcUJMyO8P6y77Dzv7zZQGJJanCtZQA6MpXmUS5EceWsDDGPMMRBqgi
GSWa2sR8c3LrxXyvu0Zlzttz6Hi2/7LpgSHHlbPnpQXnTET0uP3KlYXjEfDTGTta
Rrm5hM8RmrDTrykdJwnZtGz3kOJn2ZUgRcSo1l4QUy+7pEMEp567gL6YGTwDAmfE
UQbySkOXN5bQUHZAeRxiPSEWl1zEeVoJU7j0SQH5dKxf7a4fI9U/xH3dO9nwVBiC
2UN0JnpSFlBZqcukvy+W5AMEeEtWi3Zi6vg+yaT+k20b9ii6a3pEQwkkNNAUjmYN
6YRfC5w5s1KjZpUqj/CS89lJc1ZkjIfw7wFYyh2Rz258jey8+yKnuo5KG5z2jrWm
xBbcB35IZjT2QQcmZSzq7gCFoMlvj9wmVjPEFr21KtX8G3gcrWcZSawOInMcE9M+
uIoJ70VCDjdepcLZvwq8q+i5JDFvS3jjbohIt7Fkkk8lTLasdhd89Gidgdm/9SEX
mmwnSPndlkO6ujufnF/uksMrDHChSrYHI3bJ1NwLbZTuzJz3mXCsPkDN7zFeitgY
K0IdnbvkCw7WRjVDJGa83Hsud/vb50azRsyfrEOGj4hikBMdGJHdn7Ak2JS6Qg9q
Zhl2PAcB/DopqLpwqfXsP0h7j6zPlgCDWQItPpKdvcTkcIG1a9QMbFZ9/QF8UslY
beC6bLu+iQ4l9/DvKdefvXDBDJGJdtyZWFudc4qYoHgvm/nUkdi3mN8IHK+UOtZr
XuNmpwK+QZX+J6VBvpdeJRd2PJXErwc/pliWpHXOXXLaoPJZX3OSVoNIoVKWA1FD
QLETRrd4EG8BREYu/8Q4xS/dHPMoYdpZWLWF52VRPOjSUen6SZLxgdwr+2HtCR+z
8PF3P4dZ5FzZs3cfNojcRa9N72Lzf/Savlo7nZ1GdRJ7pPOPnTP5mi0idHgPXdCZ
p8jvq31p1LBbONFjm3ILOU8yXsYM6aT6JfUzopFsxQUon4yQDKyoPRx5J0VZKSVM
ha1cHy27KxHdvJ7QPcfjbx5aTy5+9wS3h0ctchZNK6Jx6YqwHpgy4ufyLYvptlyv
3RJChJNvkJ5R/5Iv5GIdiBydv8jTOjX2mZUcbq32cXzoPqNFUE2bNo31SkGtCVDf
MUUlqjL08LieuIeWLZbi0quV/uKDPduZ75aOBZprscT144IpyA6KcXNoyxYJ/Snb
3TsNVWIO+sgR1LKcG44X3l+y9Ti4HnDhuW94ZVXSkM4v5cgoN1/rZz32e6X0UxLl
tSnXQGUAlJTezsddl2p41aRla3qV3byvlRRtdG2CKASMfNu8NsJFkIyOO+DO0tvI
vj/4C1+PtNXGITKGs+V5SA6mdGBW+ZpNCxMSk1kozOOJe2mx2SBE9GawsywdKyZu
aMepvJNzV470pMxCBw9SgUIiHXzIKHZQHq+k0JNwZ/C3nrJb/dXmMC8AV+a9RS3M
//RNVglRly33zaxFmOAMLKmHpCFjnAf20pveOl73k+aZsQQQu4Lv3bMODl4Tmk69
0o2J70eufqhW87nGHm2B7cCcNPddx8BweymAlNUDnVVQsKYpTJbr3ht5tghdvRi0
2X+1X+Kf18/CTgzhwIZJkyC7Bem5bKKXPuZdtH/ndaHgeF8466U3/eDVVYJQd5XE
f3qE/MNLK8lU8G2RZPhG9H2Nv12jL/Wq13kb+gc+lFhqJvje9fZWl7woiqrPfy6U
sCgFlNGk3x4k98NJdQI367yJk/v5cLpMmWmYewXTNT2oU6cKppl485nMdCL4ETfe
wcDKk1JzrNH0pcHl76fnvZp8EgmzjVBLELNya9CJ0YkGWylwgkwxefZ5GIpaO+ru
y+8OPnxjqtyccjd0UZ3zIMFcELIeOaH9HksoZnFRI0F1f+goY1/R0iFvL6GY9qhY
MBRnlXk2I0JU6xULCkP0hXoMnB/XUXW8UAI6Pt0K5zmKp0tL1xZH+lxcYAIhYTMo
5wgWOCqt1CCvNYF455wstphlbGG4bgqedD1iPr5jbxpag8GooNuWAmZKntasUtcx
04aRJkqO84eZ3yvQoZ4OO6TnKhuO/jX6OiBqecwN+SJfFjwupY9Heye553XOt3Rf
VfgFJsulN+/CUk5WxWbPtTUfDO+o3/Gc7R2iFMI1J33ggWL4Hq0MBbqsC3ojZFoi
jnB0gTKfszHRGbkDxJE2pdSLLhsfqFksHsehVmcRqhfFP9x6FvF8APumPeXE49tE
pAbZuCyG1bWXZG0bf9957EQioRiCQqVfg0RKKldf3EgtJ4EGAkSxukwwABKqpQPx
/NzPpI8of+43YoXsDKSHqRQmh+68mwVsRfVtF7HJLWdeKqtbrxuLceUheixup2gr
92yAGUO824mxGM0umJQ2NF/7PKpPUhbyAjjjWfS5Yr035OZezIiO+nF+XJU+3HsG
90KYkdJXWtdlZIeSJ8WPeTYrrwdD7ZWgxLfEYRAs/jDzDSEJyKRnQqa8V78YdH36
x2dkjKuD7w3Mbg/unueGhf7LwXWKyaO3H0p71+RUj3dJfYk6rDZGkM1Lx5eU7fwn
QdioGgPUI59/hPRDz3tPiUARSD/bNxiPcJ0SJuyUIpMR07r/0r7WYgnmSXOEJ84i
YzwMohkOT+lQYCkrEf+ZSxJdVYpLQaZrkmgBKPINEiCCz6/4Lxwh28ZEig2azeB8
8Rl/23XM0zP6dE8TlPrdAVErN2xKfnOp7+sWQmxL/xaBcpo70yWZhQ/2Ea6htbGK
6QrhkrrEiFxhhwofdakNol4G1uX3gyLxt4Ay61fPKaw+1MDKJ8FnG96+envK9faJ
GVXgWs4TDuf2rESQM/1KIOWpBIn+iQeAKMwI/qJ6SREDwjn+yW8a7qCHtywI5ASz
y29vbba3lHbr7mooMNdd4VlWKJlwUFiVOnNMQMmXrkBsG0/98U+B37T6dUNucQ0r
B033mH6MyoPPj4vYrJjHjlKH/5acrkhWxHBSfPX65X2P3oL3fLLesEKUtNpvjmuo
imNxWsMLouLXOyUe4AJjsk4JhlqeikLOGRq0z7MJEscCZ4ed5n3MPf/YiajR+xvs
opIWO5pl/uLE/V5iFLbwdNMVTyu5qymlCRIoCqRgrnwpFYPw9sGaI+XpFSsSNtDn
CuaT9oLL9PGISVfEn3bS0TMYfaxhedJWhZbXSKMHcJIY8fKl00EuhCP64OnlZ9LM
v43lzQXCVQPUVVC6N/d9hEzcEb9ZccMkLF6G107euCiVQK62+IrtKicmbY6cLqFo
QbPz33JTMPb0AO7QUa7vvvWfyEUdVNRZF/MG7r/yEUal5xXu9PFnH+dUyJB8xUo/
HvSrOEcJ5E/bpfKii+sRHACFxSiNtLoImPfZb6B5+eLbrlKLvRP8QyM+dckMpiEx
Inmw9u0Q8/uLK4rSxl9TLxw7L2nDRxrkhdqZjb3+X/Y6FgZ6KsH/bV7Jelmkdz1C
4DhBU+pAeF6FC8qZFxzS3FSK0hip++SC6av3CQoVlZzO+K947fL+OJBhogvj798s
y/KPqf3nOd2J41Q22MtynoDM8pu/WfUqibsIqHG+Pf0BqmUn4Z7mUjfBXy7g9ad5
nB7UCksdmWX+8w9Ev6ZAXODL/Bbw9xx7rKCSFHtA+uOFioo87rn6f4r3Y2aLz4XO
Zw66KwkIDt1yARg1/ehPZo9NUP0wIpeRCAtqdqXTlS/2xU7/uFdo4fuoGEMTXGKx
UcDKbKYPjB/D+sUig8KQ17ZEXds4BIzryvxHrm7e7sMSNaCTsQAbYcw3dBxtJGp7
UxAnQxkqvKI9UsVXzzfKTl8XlXHN6WcFo2GFL4X/WygvIW3U0rbYIPT3tHKCju8P
zpdJlu0+whsrGlZaFAvdH5tn6AiRMnsA6w996bQ1f5RVmgCyyW10jtXWjAJUxrjF
RO0R46K+O+PHSBPIgGGxIOobY5jPdxwHfL6ezF0lVC0Xa+zoP8EdmhHictEfCvpu
BH+a2xVLruJ2XQ7YIOk3CvwGvfjqqIu/3EZvJrCpqCAEEvo0B5TSJ/u7q4Xutv9L
TIYZ6mtApYDrJ533OhUDLPLiVV6bexiaLK/J2Ae2sIq9TfOcV3WJn62dYukVktpL
CWuWOS1h+NQ9/8eIe/TqMunhwTqSym8YmzFLnkvCznK7UEodgrk1+VjGEiuuNbxI
Qys834CgL8TtAI0a6g1N3oUtvoc5+kcqU3D3U6k87WJ4Pz0pl03+Y6SFdfRLdiBe
nCg5W3TfKfSvD2hQXXFTaoXpDVWnLVLdqwH1lgKfOrjIQPmonuJwmbL+jlpw19YE
+iKhI7BsE+A7yDMo092XUNz89xOxENWktlOvY5kABXXs234MsqiUm/lZNq2ui0y1
Ug+6gsGEaCt6hSo14dXqDMSDZv2UzfJR1ZWhCeUoRPmGyziFxQsXgbd5yYB8/AMs
Ul4EUCFMW7YkHKA+ABPx7NDwcY7zR4VqX4MxbEs5hU7JViKpphO0VuAd83p6E95K
L5eaptbitV3p8blb+cJHLCWRrjdlI/N4jAZtuFRJvnmEG2gvuEyk2wTyz7Dk9/Ld
Yt+duqKmZBwqD0j8paVq3VUPV5vMmwBnn3In9az4TD1vc7OLjkZiNeLhMVMDtWKd
42L5jazItnDU/w6WkKbEi+innTCIuC7mNN1Z1hJ3+6Mxo8ql451XGkvqmi+R6Enu
e/zyBwsVmxvjWVWWBCPfWdoMb8WIEL3ZpvjD2rRffQNEwLt4Uo3doUiYfM3Y5ESF
H1ih/m0CoFeUI5Shmh139bGw4kGvAZPO/nc+uKybaUiDXrL4cJ72xrNw8ZKs3fH0
b2DrwCFvuY14bk6isyHflUI1Sj4rIw9qdp3u7qdqFEuSPLb4IF0Xrh6ydojQbvVK
yxEWSZV87Vj1JFtB/gds94KSTaTfzyKuHCtM2ShfYAnhsE5Et780ITIaDKKwxlJH
rDs51SiObyH3FcCEQar1nx5L4ltAWB2/Tk1yqb0JrJofYKHY1iVR+bEew5FC90Do
3OkO8rpsaDOi2QxIB9MrMDQ0335yxdWa7BSzAVJ0FyL7YvYwlRsHSfk392GxWVRR
z8zluuVXm3NXCcmCXy4DgRrTcDt2wiy4hRTy95AQgsZYjwZIJYHMLQRTWNwtPiUM
Q0ORO02/s2TiP4ZToPy2w37cpp0cThKau8DKq0p9vVXGewrFh3PTkInB6Ya8pxdl
kvSL33wagy5kCY1itHN2CkGVojBqIsCgXdwYLvQq5AlrybCuXFhwrL8PWxIOQDfV
PzLYoEhqTjJTfAI2xdq6Di23oDDthcMRp/32aCPSLDn3ioEUOT+/rwy2cTu2SboD
3UmtduKISAF/cKvy7YZ9PuVWKrVq2hJ8QLO/IigfaCWXdRn3jDKt0KabVk/B8iPO
8kqSkv8c2dVdPXsN8v4Q3RqgaTqvkNNN/WB+1ni/Q3uKHxfSO1wt5ygNbmmONlQq
3Q1rzlgE/OQUhNICO3UA9E7usWsBvkFLxW8AYPPceDkPOoVajT3vybz8KjUVT5PE
3tOb5A4Yvc6Cb0YeO9GyCv8UMer7oH0233eJ4gXdK9roXYN3oSrSCupsZvdkc/4A
1hIxfOoirw33R2GpErpqSH3FShapayKlHpYuSynLv8uTJo57l4a1m7BULMbflI5e
6RJ/wOxeIQYNIMO0QlqgmyNdtqJFyMKK3NeBuoefBW+T3pG6BV9SbxYiOWF2Yvv0
hT+QSddGvoszEO4qdHpX8udyz+a3KK5juF16qrbWzz9B2Wr71M3pVNwp641kSB6q
KrsxH+tGio3LXrTjlLhhz+R6eWpuCeVkHuA7Jy0pisz4UNmzKdK2FZhidoJf2R3H
X6E05esuM0jB/AEIBr4711F5JBn7fP4CkLLncmstTNkOXAUGMEjFwdyRfHG7zXLy
ieTjFsO3sLPZQJuAFR53P+8t8JNy/PHgOFfI3mo57GfI8N1CRnWaJAN0jZFYVCZn
LrrsTZB1LivvXGl5hpiVIaZc0FMFoF2pPgCCZZpcAsk8ggjhz7OxH0d6DSEwUNce
bN7XUUwFNy24EnNFOOAIgsvvpz+9bZ2rAyO29a6aTOpk5HuiJr/4cNa63np3U6WE
Zz+MeJVNAAyZIP62J0cOCX8BOAIAPQDUcmUdSVz/hdGrb4bdVvNb3aWUQuwUhhNu
In0Qm5u2xrl2kbBCH0GrKsZtSbdQ7WruQROnI90PpH/6T5qmxFXUoQrAeYHsWJWQ
y2B0d6+pp7vbwtiHwPUl4JtibbWn3nvX4ZoibAWszWHF9SFDrobXUubRUOmLDKWQ
rfzmlKJisDNK+3LgwcKNi/3xbhPsJjdvCdtjBpoUYOyTZm3Uc2ouMhmjFTY7jBCu
ZCIkZz5UY0AXBotM2HxO46XS1LG3W5RIHR+iELf0qYfc6FCEiIWUxjcQXqWUI8dH
Ll7pLKGga2zs3fZSQJMBKbgvxiXNnTgGSHruPJgEUDvkyCz66VOXINc5lF9q4dD1
IS8ilH9yfiKynWqHdaMloM40iwlkAr+9lUBB2EJ0+liUDxNO7l1gydh4LLN4yqfA
Ee1tIvXKu7X7O8LPFRATBkFhJoyL56yI29FOR27iXgomQm97FMe0D+mSW55s9aJL
ThjyZj4ex1k/tnIC70ClpdeIRqMnJLqv39Wo53JpFUg2J9qtMyhvoa5u891fwZDM
Qyo0DRM40kVzIPsAyvNwjc1ktZny4Xtlix0s/wmsy/oCMb59O+TD54THiuXTuILn
Q4pOS/ovbU8uY8ODCKdY2W8QgMPJmh68VXykmhiAkntXlqpx7TJYKadYsfCcagbS
r/O0DQdexRHVRsEHoOvMi043jybvZel1Va/TFBp0U+dRNJxSKMI8U971Vm2B5xr7
qmxzE8vJTKx5bG7LQ5/HWsYH2dnY4WyVFnGl7a6XvnMaZywPupgHV6Ic9vgAFygQ
yw4mqa3sxQlNvUTP/9AVStMP//G4eJP8bSrubZyy8X+F3qX+oBM1u5ppgsEXWKbp
dDbt/x7ExN/CvHkBghYDgwn1L9JuJ9b3YWpQ1gLnk54vkJsYVB+2ax+jU5x3+e2q
9rfmH9LHgbRV2UvbEwKst4LMevS7vxH7bwyKLGC/3PNHkRoHDNZEFdRg3sZw9s7s
eDOMh0wIiwMQdCuQBt8t8wjEAFaLL+06fNG9VPRYOxj/UHhxlzKBW2zY81l6oyA7
NOvdk++3lfuGhVH9lZXQnqxw0JZgqy14ULTg6P7nckQjGDi6Uwu+TnOrVJB1HNh2
QrelFcpcS6D8ljIiBKHcvY40t0G1hCiZEkQ2NKDL0MNONPyXeMJAS8OowRHRg9r7
hPG35fCEkwJlJKBGce0bh5XEfk5NPjrfZCCbgmI60X1rwpscq5XZK3bf5f06tzBa
bT4ub8ASOouctkAy9h2azq4lcHeREHqgSzH80lKLrgJUdf7qxyVgxcMLgrIrzbE6
y/0YEAahWmSeNWIxySUlyKudVz1e7pJ+TARNf9oXq01AbTqIUA1Z/PmL4cGjy6kG
GnsDxSznpdAcxG8eN7wvC6n1otX3bI2B+w6K53nVZU4E3ho8ckqEKH63qvzmUwt2
wtt5zQBcgXFUHxTacRE+j0G3gjdZo2wvXyaNpqdHZaK5WwKRtMz55dC7rvNOvjTe
6kKJbXGWzPw6x99l2eNaSzaOM5S3d4QirlBSzDPzIpuHTeBJwzLQlZqcXuPD4zXy
RCGk9boe7PRkiT+X1iKPgychYRotgJV8Zv9Oq/9BtqqlmhLcSdeQWCjWppDiR+IA
cynmt6JktCSWKHVvXma3jxvDrCpHS5t6kxY+J4hUypfFN+mplElxfZa9nybK20EY
62LyvH6MXxBZJrjw/lAW46MbiKe6GozcnblQipNwt7DiJCBs9YawM06VRjskDY9L
b4QEQ7Vcq7uLWkJAudqI3BqMJIdHRtm/H68kn9bb1z50u8Fm6UkJke3LxKqH+gU3
8CDWtyU0L8jnHpXp1/IF+zCYJOisrLBzrT4gkosn2j0G36mB8P7Y4JKyO6GavnyB
HZA5CoL082ol0h2XUL7XAh9RQth9F3MhNX+zaYV0eqFljD1YWo9dOaeXk1Fe7lR5
zrremeo5iB/2JkuYcbf6H51gwEUYppjyaAziFgqQZz8eLUOzQm0YJkxKPwUc6SLa
YMBqNjYVQEl8RIzPauTqyYrUGQAU+iu+96lXLsTC7RMhT5VD+lzA028eTxLsT3iZ
+DTrTse95Mc3RC2CU4V+r344nPOocSivmzzhYIYAzdG73Q29V0PRNFKbPDZJQVpd
cxOnberTifiztbrX3xL8SfARs0QOT19WTF2yVH+ETU+Mg1z3DPS9BodxCW7ch0tB
BrZNuo5cTE8TOTRLq8//52OLC79O+QpzI9lgRY0hnaGBRmRiypFxGohLV8ggSWbJ
gRWyRwBPZEco41MXZdr9dTv1J1rAZSt7PBbGBkk7bAOhEWwLvzBedTfUIN84qyCT
+B1crwOEcjNagXCcooyJjySSWVcUqZZPNcEJ7/JIAfpRobo0h/5NIN1lK+WCEsqV
NWDc+melAsxIwsguxLiv7pH1MNXkz1mLmj637Ia2ld7ZJwGQ7jpcyQ5Rwrholf+z
6BoY6zNJVlPPwY/Tq+EJw3d91fFfVoQGeAikoOo4WCJ6g1SolEew4YAa8GQE9vNi
0mWzH3z+Y+z0rmWcrEPw1eJX02Z2bqjPYQ14OXY/t0b+lBfh22KsOvb2gla/ZqEa
RutJEWIhdWq1rGTjsEHRgOXUxXLmhsZGcaEOWQKP9br4p3JtFgWi4foJMDnG+BNH
SSEx7Dlo3H/0AYRDTJUyKqkkKR8jLW/Isfr57v+bMXmUm4Y8Y/pI2Z5nFiUhBDsE
spBcAa3qj7RLhQAqQ5YuPNi/CEw2OFdNOqQjHkWxmb3qPGWE68v0jAxR8PM6rrYw
SaL86Jkgeanu4xF1PzAVzes+enx6L0cVHam88bhlVo9OIOn4y3zE04Ag26mz8AVL
cw6BKKKhRcJmX9AVFmnh9CwAXkbG1odREEt/h3SP3RH1HQoaMzIdYNI8qU/6dLVK
DEHwl9Jf637PKhKYve4wbg1gJSKKxvPHah/9dA4d65KNtYU1xYhUdXQAeP7mWWVN
vf7wtExNxo/HdA79E0MfHFSLxvL6DRkVvUnlfj3VoBa8IjDVaLo7woNKUWEFFCDq
CLLNlW3rbwgBwE8NqlGtB4rmz6yIvcy/+dP/fzljJyHDf10Xo1Ho9sP0LSLjrgRN
BZ4HHKCK4uEHgRt3PYa2ReCfKrwhECbT1dsbYzq4hiucNztRVT6OJxa8kOr88kqr
WW9B8BuNbUc9WBqnxSQZsrMSlkMdGRoG2ddskgGZ+zYpxoXeN1D+ESEYCEQLoh+D
sFvOm5r9B6QRS0ik6u7HLOxk5wu/iEzELOcetDIC7ZFXCjbcfETGwU0mrrYHyuWT
ch73IBET9hgrhK8vy6ZB8oi4zScxbj1gZ8zAytGwkgA5ibNlkT12eIbRGQMAqtZG
PVdj4IpviXN12FG68pDn3OyPZRjmlaNTztXTdv4/KylqGoK6B84Z4A0nE2Eafh69
jBYPtTf0SXn5LrVMFFu2GHTlrX/NAjDGqTr1ZJ4XEj2oJkKYiCL6IHwQ3PIq1RiL
ih5tW7NhUHuYBaax9jYui6SoC0uXpeuRmbX6KFbCT8nMT2LA8TnOsHCQO9CNN/Yr
AnX7g5TM+xTrh4et8AZkmCVpHd+izCCfoSJaZ0m+DMTl095qE6d8nKFNbQv0+msJ
+eJCBrZNlmpg4pZFu/o6bp2/mqiHQNVAxptDnB+tuKPlcJNvNal6eK2hzs1z2TO3
3K7S2vXfgQha5R8DExmlAuxkbgUNZPqirDkLgYTaVJYbDGncbtLM4EEWbXVOW8Ly
PFD6h8I8T1FfEvDSb+CzqrxodtO6haVHntGYNhtzeVz56oEGFhqGDJHrNtiQk7WA
+Isk6QZIdwGLYAeCc2/y0tfGLt7zgkVUHd3qt9j6uECJ7nOLqepL5TTQdh0v3vJc
UIuKKBVxKFn7VEpvRdUQFMGwgPb5HZR+Z6bgif42JuRbXQQF6Z84y8d71lQE1g8n
TKj2t0N3JFS3tdd4DVizwbzPAXUEMr6Z9VQ/fDMec4u00+rEL4s0itGozmRoch61
1+P8WlrgWFf6yd9oGc4YkPHmwA9h0fu8yjJ7BKeVPciMDaR31Yz9viddVcyrlop/
OKK41eA4o64KOo+Mxf9AU77f8G5Lg0Oprv2lv+kOMqSRrvk29LZsfvq2XtAmJ6Do
ELIpXvQHSc1HN7ciWj+OhhOUH8t/ydSk6SBsrTWctBqMqNGFCSPRC6bI0wgaDYvE
6rHynnl2qk4tWIrnLunS/izN7vCV/EO7hjvVkUK3zOCCs5rcfsq8uePBMg4j47jt
4XPGUtdqtJx9GrQ0VGx1V6V0X3bJ07Hiu4JcysLV5d2mvj8teM00ujeJK1qd52k/
0Z8abnDAODtDfh+zO14TfxCTm9PloG5yQaArKD+5kwWqPBLwZjHr6n42+Zt1NTJ9
vwQ1rJUyePr+FpsWJV+D9uj+Qub3QzkKFBeIfdfKWJMVJ8kRXkhpfggP4530Eolh
y7xW/WB/xc8L3Hm+y6KK/WVxasyf5zQCd6YNgKS3OlwGhGmhy46Ko16uITsa0Abg
ZunfbHt1XFQZMs0wuTGt9JdROiYvpq9UiuwL9iDIQmOpfxOybPolFE3X2yxVaAKs
9oPr/FgVBVwRypF/nfO1ntjGRnUWw6rSseh9ODVRO4kxczXKTbRQwDOO3C31adLc
TAKX/2ufdPmSuIWdkZeUf/wGO32bcqSH/5TkKZTQHLCYr5GLhWX3yobPml3DQlPv
HybQ5CiRMYqi7MJnVVNb82UExgrGO3tC3ihRD8mLicy2ttctiWufUCP5MQKclX07
tU1usVzHrDdCz6moRcEzVX1wVtQZDYywKuECMfSiagIxOeZie7ZmVMWX5khaXtSU
h0mmzM/W2Cs1/CJSjBEMvT7Px4Apr+L7ZVkb05VBF8NnHi+ZyP9m4OUBXywfKdnO
YYor3WmV+DA9qFpNw9NHQ+27l9G0HHCqZKxys8jOxpFpJ9F7NXW9P7+h3m1GRmqb
SwRfFBdto/+QZP3/PKlawuJBJqy6m1LzqdxV/uJFlMlDXxjIeZrKqqSO3kAOeKZZ
NsfVFOMebecdexWJ3Ftx2qYA6nqA2Z/E65O9WRdgCRT5hstqUCGdP3jzo8ize0tp
ift+AaDJ0DpLqglx8ih6CAa2dIznllP0PVbbUWEQxMDfG0wZyTWV23zzza1sGMvM
ZgQ2QULu5AwZFKPujX/C1PHx7Gd/71t+XFa0e80V9gSn3ZoXIn/hktvgG0aSevCZ
Q4oUK0t7l2hTk2Nmdr/uydb0rbYKQ3mGganCpNHeYlChej+1SUvcSkfo9frvYs1T
qaXT0HiYv0PxJHxZh0TKDdUVS9XIfKxRX4viC+7eMljbaSR9ejNUuUDrkFVZw2qR
/0JyUAvNHe4OUgw8cJx9OuWL840OUr97IWcdZovrmlvpavMVbRM79P8b+jldhC8v
Sre/TmZjlZJd7CjUmRjkqGbTf4ugwttugpl/3nj1Z2p2XRvQuWQpuvPkngyxxJwv
SDGUxsiVlYupH04Fzd5VGTXQ/JYsvjd/zmzRVo+8o7EyGsVAS/5ku+ohKP1sR1Hx
yMNy/n7MXhimeyXn0gkA7epinW52gxhTVq8CRV4+gB52K2ZrKeeoGO6KIrPgv3Qq
Vl1s9hdNDRp7UDQy2ca0qW2bz4aXBDQ5k3XRrc+WeimZH18bK4/CY/jqz5YOI6O1
Sv5LxfUV5fThuD4TOMD2HESYkaGuvqDXmzu2b0C1NLB4RSTJtPdASlojbP6k7sl8
+Eb+EggUNE7llJ1YCE2QA+edNLBtdO4a1VQcY3wVou+++4+OfUA0m+zHD6geVYDG
httdT59r3ilCIwrLszdsnRzEHOjUH85yf4owgq0xlSYEULS3bIqNo6Hg9w0l29Yg
486OBwJKt3FF2HJNiCuynUws5mjNsSMYAY0qfNq2R1EsTjKkNvhocV7ya1T+cMhB
s9xx/0kz2vhAm29i5Ed2FuedcpM3J63ETVKsotN+W9PoaGv40WM378x8bGBBEICu
hXxAdDz/+XGuB9MdZPyGA4UmVaDkUV9IWf3DJwqkjk9PIzbp8uzrg15CDR09We5q
guRC9b79hgH92XwfKDz2wvkZr+OC/gWI2xz73CIgPndisGjwGgQPgmaCnH8w61rH
ddv7o4JKKu6i3lgwD6RJqEP8FQOF1v80xk9T1G+ifzvSFYuCxvPWZT9M6MAE5/+h
YEyoAVWM01koahIRDNoThmLn+heuzRyEAUxwFF8NRYdFgoHvQGhHscxH8xRRsPE5
ABD4LJaf6VZASX2V/m9i7jnMniwit68JIfzHAM0ZjL8MyfLQMDe/RLNhYp7bysOe
kficdwq5X/zlDgqS6hZsUgR48OgiJgm9ofkvMLd+UGVSTyDvhI/wtGtI1q09agPB
/pqOS3sfDs/5J8+6eAo/M19/21wrO2ZHzSmgQLOnvsjOXrDDuO9sGM8jtTg32WVg
9GmjJGSx6cTw9v3bF3MLRMaBLj5rWM3Xq+Cr0rYYFMBerdJtZ8xrvuUkdQPXDek2
yv+P5j06Wo8Hn5BJ3ZwfK/f0vDVbjiIITHpEOJ5n6JJKJDpUn4GIzC21gn8v6FL+
hljZMK2nfJysE4zG0vDn5bwP76E49CqL6BKRZj/+ol5mC3ugM+AqRUBLPP8dDT3X
tJnJpXN69ToGl+WUBPwV7jm5wODOMQ9rYbS6+4TUI/jWzj2bSpJ+jRGhpqwVOliY
HhHQovg4bcnh10nugzVWXatx7xoX4lN5K7mzD3IDZHuC4/GSPiJHmToJeV4MPi7U
gewnDQsJhAgICvRnMS+R9MH21x8QBdU210GpIFAKfWA6ERcxS0sTFppB65cXku9n
swVVbtN8UYZzr6HqLCqSxlK2vfBijf6Lk972YyF/xKxmg4NJkw94ZQOm0s852j5O
x5t62DK6kotRIvgQE07Eu6jre01P2vs/9nsN21Gpte1p0S4EUiPjenF6fKD5TJcL
JmJSzTw2hXVOvbKDJKnH0ZNOijYSbQLLILqrTlZXVHe6qjgeaeBiwOS4slebZppc
BVU2IG7ckSwsOjw17AUiZX6QYZLXphYIZVt+igcCU7EWBzcJgTNCn1QoYU5RD/rw
Tl2tQdDaVaeRju33h4HVI7Cm/Ty+yTIV59JjM1xjdrfWW+660Q5CRVAGAIT95wKK
Z5orhbxJ5KaS1DWkOjQdzcoYSNUVzA2eTPUB0lzueDUg+sip0Rm3DbUkufwiH/fr
k6Kkfl6rC1Ew9zE/fcVsc5ZbzP1kAAkLBE3m3SigYiDAC9D+fAgEXbgOSxFsV4DX
/NzemnVhYbkX/qYkUdj9mjQz3TMFNFCUvn/icoxUf3cn792/iNQQUJmjnMV1XRI7
PNULMlx87ehMtgpF7XIFSF3XUzyJ46pw69sHi3wEJq04EuY+ay/aKNv2XgE213Nq
yIXl5hbGI8ifDCEsVnyNL/T9us7geMUsW2yj3H6G1DUI/IckeCVYonI210SaJ+LO
99a7E4bdCZiT/ZOyNT1BzIquBQwPnNOCwTZr4l2W9IiOZEDpOafoQUhDkz3tUYG6
2EXmastEhbYAmmzEp57Ojde4g6HkUL6u8ZdySQtW+HlDMvIwuwnAiKDOIAMkGyQA
3/rTD6JQKYsSJj/XyDT6tNbO//Rah6s+WeTCJXKyID2Xqps13/xRwIve+YQezlSQ
lX9pHOnL2gKnfJ1I4aS7FhRKRXzaN6hOtlwAOfZUNL4as1/OH8mz5BJUG6e3MK4N
F1ZFIm9WLHeyv8Ovz7iAduIV85Xu2ln8P9cMcRO1SkUWI8kl1ORo9DMdYsUIlB+h
nWXw89f9SdFtkJwWhgCdsnqlBwnwS7pNwsBvS4HXjnCKHt31GzAMqo7i1p5Gn0rO
7PH7I8uMevVDYpRfQsQw1sbMw0kkTB/pPOEJq4tO0uISomxk535qbyc/qSYWUfZu
3r4NqYvsE03rYtYLaKkFgtCkebC+nOhHKhVAdWY15pNKC/BJ/ss/koXWNM3/JHK8
DfrEckT0LGFnoJyKZ1RMnYyTQZMBuGv1SCGHVYbuWKwYkTqNmaznvxD8fGjCAyUI
zLolso1t0XKjIUU1eIXcKXSSpyOeCikzxR9dgYhz5Z6HsAX/zMZXRiqVL8ZB4XfN
n0izybdjD7CHP/PczxtYJYanRATwU0D5h1k3FbLJB3d0cpnnQmLMfTo1ILkEj3cH
ZaMCDCLCl4LoBNweCaiXPGthMzhGFQ1YuYN653Zmg/9AC4Zyned4Tg8ecX5ojJqO
ckMk29vVdzjIN5gncukj+ubR8/tH1aFH76IXKzVgN16RZkZj8oAbS0IPViVtG1Sf
T1wDHUnpHKW7oTHUB0YQoyYMmyKzbnieq/xKG67nRvHNoatJ/Kh3ekg2F0G0qVWU
FuQ2SA9rdRo6G1ru2hMqXLEjjEnsVffOXGTNjAsNmU25jOp48YCHy2ACJS++cbmr
ZF3h/bPKqg7jKI8nOwVbawIuOCERkXcaWmaxQ9y+DLFMlpDhgNM6AUVk3/GDZPNt
XTNP+OGixac54O5JEEm7ked8uKJIl9kndiMStfJQGjzdCaZUp6YwctrhqKTfb5dt
dNeGK/xN4nUXHIomxwcubbP8zhuNZZ/U7g5B6cbCQBuP0o8AUZZwdNzdTvUojS5g
41h+YpodTe/tLuG07IYs1YynDvnuJEHcPONdr4AFIpuDVlHRszWeZDsdBFWGKBKu
foBBLShzDd0yuGbNrcrZXSJPVXAJGcg9l2sDnCniVbwBhK/bw9HubOqkdOOLMVEh
XDzAxQgllnOzB8x6e1INXXeHwWOqN3zv+KXWwQWLTJkhxY0m0fxS7z0BpMq3+NG5
6KhZihQKhg3HTRAwzFo/i/eUxzs0d5JeKQ6gTnx4Ts6zAwNH84z60igSrobkenrd
Zs5iJpwrJEpPE52yYRRJmclTHEoFjdCxGmTSXFj10/UjtP2hfOn1OCQGrgRKfV6Q
FabTm4QECQqHStiR301S9sA7XuhtM3ahFDtthK+NW61rFZdA8zgYDUiZQg3kb7j+
kzAQAS3LVMeXAGJhU8R95CBHyJ72HqwByzmGlpD19OC1tAV+ZSIbQ6pu+GzckomG
leZ2OToQhA6nuoAZKBy/aIwrratxwksSFNRZGo1uYdy5am8+z2Z9yjNX9V39SiAe
DNym6Dm+SLljdUXObIk4qmFNdVcABq2alqyJXPW4QWadbCpxkvXPNjSUN1TrMLAl
2ceFuBxKqYa0STufvdr8RqK9mrSrq8Fch6s11ulUPcMMoiJWCopisafmTBIwEX+L
Pr5UtIE1ET5h6JfpXGMB0pO3SE9GLbT7xwmQL9qadJrVc2D3ufovqfuDWBj7bNyO
TJ3elChiT2NXpuo/zQU4Fnn471Y2fnOuPnS2U+id5788xpm0ynZzBaCpo0h0H2fA
zSaixlGQmDNGvJ6IxQbC5LGMQ/TIzxqjJ/P2jnMJy29YFE+IVNiiu6hs8vYg1F7K
7O3SMN9RX4WVeeUWXKq00QNozj75xHhuzDSrOPg0z9EpjQmPhrGdwfS/GkrP+ATz
vkbUY+SpqMuMkjDgAAc7eFhQqkydR84qfuWcuukJGYN98/SOkClfJGRVQGBF9gwt
JuB6zkgz0vqjvUF1BqNrya6l1PysE8HqgoDsYEZfUpzpyvHkMKfYLF+L9y1pNbp6
EdedIF1Lb1a7Jr+TWmiqpLwntN3ach51F8ENW31J7HUNgBso2xGCiEowgUFcsZ/0
M454QfqIpZLpnvj3DaIDrxqqY6Ml6VsB9gdsd2Egy07gs+xJioAQ6P/W4xBSG35B
ICfHyc8RHBhQjl7JZWfLukGmdb/zDpzH43YSdSJistuxAxA/dFqIXJR/AcWHCSV7
tYxsm60N4lY649Md0rNTN2tQE0oJLCVXWCP0EzDcIcEbH+dVY6nCgLUxWMFTEiMP
RHMHW8IaIpbvXCzGrRnRmdqXqwZlOlLOppC07mCgMPA91uuGB5Nj92/2TkvnfYO2
3gkc536Xb8+74r7dFdgPllLM4BSkDIPiUaZ+zEbjhz/cSZLf5dUQ8cJSiNE2UqrU
MFH6BEWkVrvMOeh+8G14wTUMsDPHvuGnNp9i4lpggdeibxPMHtwXitwvMDwdSxM+
TAOjzAsIEowqtvYr+nvGx2mZLu/tJgSqw/ywQ2Wf+Q9HUqqQ9LBQxO6/3G0xHWKc
PTykEelfYGX20wTDKw0oZz7+m63Og+bq/y0CBm5+Z7jA0wL1a1AiTRKw2FU6E6Kp
iI9I0ZVU+9HnvjbBgPgYRrRnq/xG94goSY+OkERuGobQ7y+kAwHQdR4x63SO+zF0
BvPehyo09kUoug+ZVnJzZkWUOhCWuzQZro1zWt0Q6oXX9Tl0R9XtL7R8FqSextw1
QKcChxrl3eqyUJBpYBoXmRBC3imHFQyYh1T+VHxlEvThNZfUkhhHRJWj+2XvXmC0
oYmoXz+vNbwfr7yB720koxMm/LifW1gffrIpNjJg/2WjAkkf9ATyyEebiVDfho2I
Q3yUimmdWdZXa5TJSy5pLgxCfH8wyc61A9ia3CRVhdEJgIrHNbTksJM6+1dHTber
Y1xvkQs3ozUmAQfbTEU0iRiIX/7wn08xVcnVZYYF70BUn92SXDDrpQeuu/+4qe03
e0BNFxeToRysTS8fjE/raUgaGOcDeeeYR9VRXlc/UVPWNx7Josf9r7pDsn/zy5o/
yDJmD87PlfaWDiI39C6HZx4zbcFFxrUQ0PqiJAE00+0CVPjVPP3tojWi6++G4Ocx
XXuA26WY+huV2up6Ux6bhWYXx4dI569pXia+zsD1nDwgq7GcelSMGKJl+zXJU51h
SB7bBa0OwqITjth3ZpwziXIdOVUD1pT3et/tJHphsUk2kVxrtpkNa3PrllKotkFd
4NsrFrGJLAhuewxGdLkhKf8YdXDmAADGwWr5Gh41IlRjhOo1j6gxakYhWU+RIn2j
hauGihwjFCrpVXg/eK6YswKsQ519V7/JqSMUJQ+BIuuRMxBMiKxhxrv9kfOzq7L1
1oD53FE58lBEBHYOaB6WUYnPpWWBL9UDujpNLujoj3l5BA2hQRo7/aYMtx92DTQg
/t1Tp6ITVsebbn65OmHToyR+YhqVpsMx91I4N0dw7SwFgePKsOiP4NNliEKNBAFo
Xq16ZRxK8LNAI2tyL35nsSh2tNqe5aGp2NfBtJRjjCm1yQBu4UzaukMkJO7vk5uR
CHjGnp794iFVf4HSETwLdc71+jqSTi/DUSqB4l7wq3grYUwn0HMVQnvj6/XSE49p
5470DCnOOueDsEM0W3RLdSVkzI8+Moh2stZKRycWOfXHt8bDV5EG7jZsZEd+wK8r
wufWEhgTyZnOnJfcExKjcgSHQYjuNYzcZOvKSouYO3Qa6gQqu5idPMq8LjjnlDcX
sYHR1W+AEoU1zQbn3wDhRB5XXt1owEKYLnI6I2wutE3T3VhtTOYyQ+2s4CaGegHU
BCIsn1QpI1Q9YHLsBc0eNE2MIqK+cCiVNCq6KGtA5za/p9oCd9XTLWSiQv+0zjr+
WURS7W1dvQGUL4+BnAln5fSww8H2PxNQVRg6hpuKP+Sw99MgU+70mGQcKePv1+z6
skp5OoUrVICbPKNZxyZP7ef6OCauJ+yePLv82GTP7XiUz9KvEH8FdA1v3uDWEUw9
AwR2DnrvE/vBt4ZPGhG1HTsBXOq+fhOybG+lbjeehGPB0zGl9gHd1CW7UP+qeWs0
E5JsMLMmcafgmgfIA9giN0ptgqO0z8+XCNqlPM9pBANzQUj5gFSpu+Duy3MF4eJk
zR987hTnju2xH0naYPAMc3sO0lxBQed4kqYGDQiYVOPxT2nJH2d741nMcp/Kqohz
nAxZNoaJ4/oFBlKukoEwzyQB1hyNhsAzrXcL3aziJLSf3vaqLq9RtbEKtkcJrLF+
SPr9f+VbaBov3COX6tzZ5i4+D4iB7uYtgRhn1R3XsFy7CFl/g3r+cPrqxEPuwXNy
Vi7Bg/bD/EEHsl++gnMHwOEFDfd7nsn5tbb3OSKaMt0Uwa738p41xlCRp0xHXXJw
hQfQDRb+FkhC6wZaHh4g3y6d8h6NXCWRy4Zaja0jKlm3SpBwA+trziPHnwIIlRqf
PBpUs7bOPKyNMogAjgc5lhQdfJ7E3qVCt81+2q0XgrCSSUYAUht9mbjBCEqoMkKB
DvhAZMvQMYMRlKTtFldxSz/2IqlORY0P6xuN30Hxs/UvRKg9esM46ADIPwlAfqGj
FrurSFHv7PeJhJafqZNLUc2KKXxz6dq+JRJVAVBPkxQZru1Oqgv16zkCwL1ctwt/
MVOgt3n5gJdDRTyWtk+enmdjbEcLS3ZqNvu7UinhMBr9DpYQFDC/KHESPtXaeyv9
9m5+06qXkrUTkgcOxPxXJeWOeTdFLyZCN1u6byi+TNCNodbp+myDIG1znUxk4enM
HdjCgFxnNxn0eBt+rHUeABLN8VNlm+5PD3YEPWs5Pvyxp8sH9E/hibDyCEjvmbPH
TGzKpzmY4jj4xvWvAVPMkt0Q+aRVrW10/Hu2Fw8pU9q25rl7m/4PkoSA1kzLE+NI
q5nrWflErsg+Vb2BIMAfAqOriqRCcKKg2MA5iLYmADBC0EDVndY2E+SCoOKempTV
6IsUmJRQphedJav09Oq8rKlTBYFc4EhCEAbLx3ctAoIwm4KuqznhocgthbSi4EMc
gpf/UwgmgifCTmJeXmGmeTlt24QXQw6UVaWEqrznlRHE/JzyhGEmLBX94k7FZ009
cHKmtrjCbn+iwCjnwm9YzRp9ldL3n0QXdUwyBZUAvkECS3B1gA6UaZRAzUBIrh4P
YufnrrAXLSzYu+gN4BaU/9tC0ESt/8EzMkXkhNdUbUAAFWwFa2NGpXq34c5s1EhQ
nwZnU71sPrd3S3YSaR4fwMTJF1+UmBzXayqSk8kk23MoVV+vytxE2zKXc4aSuSx4
lzPlffbyTkaHTi9J3YwF0VpvDOXvyrD+zTAs/+vEE0iYgBgwzGdJiXX/qFuugwLA
ymIQ/CEb6MEvfH+8Mqel4P7YUPWcJYKl8U8wNHz067xKPqO+ZsqtElsbMOphTQtd
8WDIapcwjOpIWniXDglDuOKIuIAT+mPFFYyDipfjgQtJf9ugS7+7v4R12KsIvnOg
dxokS9Gwpvuxyo0Gr5IvGY2mG9mmRFowzN+Gf3+l01pdAZ60MHEqsOdAvEm1Asqg
Q1pcDyaEPnHwCd2IZ4MFtKecx4HAT0zzorz9Q7JAUJlvEbfvUScHsQh5AoFvgmKH
l646rn+2LoTtddZ0fQBMeoMqrFJizE15/qTZvltpvoHnHba6slr8SxCejKzZI4s0
AqWHK0YrCVxCioahfaccO50OtfKQhimFiBwEHoUq7pUkoowxC5vjhA/1o3cC4rg4
3ercTZKiu+0t3xEOjnhGqU4PJ38X6QFsklVu8rv2j06iEFrApkoGCPVdx2//81O3
myLBOc9sGpNY1m7Wm0MEhwzOp0Q0KmSm8fD6mDZU7ZwcALiGl8NTUnnWYOPRSEzG
LuNoTnxU0MZ8NSX4hhp6K6vfuSc7Kl4F71WLANOtuQdtUMn627W2M3hXps3ozp4Y
bTyAntBVRuo6Z/QcJZGGwY7PfqDtFyhsU9HEdaVvBZM5+EkfZ9TeFZQnEd4Pvsso
iThB5T/T90dBkuZ2dnaldJdOSZHyt5S1lgaB8Yily1Z2A/+AGBw4jQgckpjrDqEG
5P/sVmzh9Vez99DChrkpYNkNlPHbMobYJMbDhBrQVi62ECZan3Z6JRQszGkxaxYy
k8/Ra6KOiJRpxrfVBo530dfcVNacoWCX1NTaecJm7EiJ8f74lVyNqKhAgY+NcojA
+YqPl0jcfYfbs1sIn8UkMoO2RBV/gIZ6zjBQrFfRjApzBAGQM72U3uwXxoJnF/1/
4YVLz4BLmT1f5y7ZC9BmEvHoAKz0QnQWvRK1JrYu/sw8jZX1kEbUR4ux3a7OPwLb
5dZNJvmeBKGEgz+EBMMEzujs4+fV8833mnDmS2cznUtaEy6bQe51uoy7DfHO6VGj
XhibP4ibEa6JF7ZP6+JRGQKe0ex2wq+moMhH6+SD9/8dHPjGIjWzdXFUh20n15Jw
9KbFDxnMb0xFlPJGFu8oYZrzBZQfjDG3k6z7gUODiurd2UPn/rirIF6qPzGW+8tF
WMGPKB/dCN2g31Qgzvv9ypEUunuyT58fv/VPqsKHIOZ1quKZ2zOSLpIKjBNuga1t
oO8ayULb6ZJ1bj9WdcfNzPRW2lcMdYeWcUjdRzgw9cLXRg8mnukZGSxE+Xc/Pp3w
hJXzAKBwC3zjHnqaXRPav+3nXFvyVfw0+EdJZBhm+wF064qeB3WTofQtYegHHmsV
Ur/m2qu9KDRd6QO/YTHOE1kX4eu1m9ihVmgQt9Evb/8hvPF2pE+E4Mi/Ot5aitnr
2V063FAW/eG3bPtzBGZzAj8lz4vUPPtkONU1hCFVYMSpxtydIIm2Mz2qPxXtAp+1
d9SNplsYhVEUTP3KyDVXq9kD8NWfY9OJXYr1DlpLX9ZxM7L4Uj/meoKwiBxPhUvt
wMpI52hSl++mYgJ/7+BHRkdKgGYbJnSHW2t5j7QgrRIb4RTv1iMAd9PlaY+15E/S
rSQvfy/q6lCkkenwoSDTuP0/JIt5wbBoA6c2nieJ0d8u02l7xK7gdTXAwdkuNFil
t7Ef4GWaGEQ4GJGaZrlava89OOqkARj5R2tH+Z5kJqg2y3NPVK2Q/9yUWCBuchgA
5iWpUDEU7wBF071gTjTqFi/Z9mxmfL4n/boRpGhZfTqwuwnM3Rmma30ygbmyI8oa
F8s0tNe59TnH+uKQZsGfKPIbRxd+zhrUVMfsxgdYSnp92a+bngDk48Gq0S6SKddS
1Tdv9ujRhXfM0Ai/tyaju5yCtTCdjb9RjjwEvOmMo3Mw+l25Bboh2ARwvoNi6Lya
QSinz1jYMzALW5TNpr1nvnXZXElk3o+16hpYw+BbteLvGrIBp0g+NEKMgLj+9Tob
0Bi3Y8Kj5X+wbsTKfk6ynnDufGz4ejpmWGoFLUQ5uQy/6poj0Zqy1NImdUKV16tV
oNOB9TsbIVeoWVPNMqIh7rjHEz+dmoJ86WJf/Qg8dzS4JYm0HuCt/JK13jZcJOcj
aEcinwjoNohSbMZtt/U4deVMPLlteobcJVgd27gT6pOqYyTayS2KE/qcZPV2WDkp
Xk2hjJ1lZVkcI0mjWiP0oy2Igitxbc3of2XS0td5cNhzU73DQJ0I5dJGyiozvrYj
pr2SzWllpGnZunsMBldUVjyfmNKb/cAGhFa//dojFa5ZUQ6hWwp54InbhF+BXK+p
mQJ4tHr1kH4ZYcy2ykYxLLfvDxGl8lEfHZuI2UqdtCVJJDtTwrsjOzL/dCAbfIkK
2TNBVPC0pJ2ZhtFGwEMo7PfqI3fRn0j9JXLQdayIwg84+h8CL/rcE7W53710oIEt
q1ydhY0giKa4FijpJUCj83lmR/kPXNvFfUHSX/AfWt/AUAMj2AfgRL5tR3Z1mkPv
mQqR8IOFrpe1VKuQEHh4S/+3XClA0f1zQo2m6EWm7bFIc622tXV2yrePsdnOh8Bs
NK/Fce/EWpRCIL9rKduBBgLWscvC4JndVwPjS9tdYW+auG4WCkdyYpbn8PMXMjOB
cu+cjUW4cRZbOKTYzgHSISg5lS3uZzU2Tv21e6Tt7cIK1Zq4qpM+d4QYInSnT6ul
Qe5KCXnuslS9Lrf1GKBK8tHU1HUuOqPeVh/YxLvlfZTDAy0PI4Pu6dzFYBXCBFst
z0xO/sE4kDt4C24lTSwGYX6T8ATzIwozjo3d4ZBmdiPoF2c8wll0ARgP/4ZDUCd2
ANv1Ax8/5RpSfv1XJhpwcTFt73Sbw3XQn02hwBMLu6KYlun40z5T/FJRvcWcqeZR
v4dP2LR4Yr5O6F0DTo3AWup0kVKbmRhxhD04W7sy0LfBrPjdVGhGfBc//5FbWz5n
FM1rhGvu6ymn9sC+SoGsah5BWfyBBAMkZx93WDqtlmi3Kt9TVIcyM8bXHcTMDRfY
OOh4IMjIs42xuledmx1q4/8hTKVTwwe3ZXosB6/RrhkDz2ve4dwtwyYqcWqOzO1O
3UPoJBsmCwMwnoDwXaNiBeYy+tnKl2sXGds2n2bs+LBBwxToAcBMvC8A2LrnFqmo
3R7LhL8ZJ0hg0cyqeeIGNoLh/o7hLjaEQ3rkA8cVt2wyHQaxPTuSq0iL5dbz0hym
ZbYe9FurSHc4kRbYAQxy6sr0z7n1qckpxO+KGhmGltkG+fpBIT8iooPBZAumyC82
qsWO0cGNEb+vlnyfEDpCChAb+AJnNWQ8M+XBdeqgPQfi6wQF0dN7DKJjqCk/zGQ3
0MvAeLx8IT6eGK1yyHp5k+Kj+fBPGJr41UON2a4LQwPe1LHiUvbBCETjS93WY1Sk
+uahbFwSpoaHJb72PQx+CBSqSCOC+HzaId20PdJLH3/Dbd7JVwXm9OGZGqtiJY4g
BVReKnnkjgw72NlQUeI5I8MVySJfWXLETR/QpsjpFPIy+ys/JV2tWLt1VhcEi/Kr
FfEICin0VzrzoG4SQaadQ2GgIm2AF/y0aIttZkN8bIq6Qos3jAaoz0ua57Be08RP
1r/9OWC+SvYCwhG5N15JNZtySGsjHJAogZ4Y+lqhYI262x0WZeoJg/wL1URMDST8
pRKJ168vuUk1wLpwQwJG/zsFDMk/rJ/uLya6WIhTzMsuyIONJhttjSeuW6TM9xeG
3Se5iWCNdoAfiE3WTfcK0VUXf309WMdWM+S0LXZkMzNkdtDscihUrXy/EdEQQaXW
2cWpusaFF3J9c63FdxqXJXIIHGfdEveWO/w3NdAKxnZapLzrwWJreQk8ffDlFhOL
WhQcWofHT+Oy1cHaNxxCOUrOEmUe5oK7mGsVjO04D9aUgXLerPYdV+Uur/j9OPo6
MlswbrxnOYxAfL1tWS3LlMyJasvLgWzfu8b/BV41h3vnaYuzzjtdgn1Ax5S5IzG2
R7R2GpUoCJZGm012uSMot1BHMi4YAopEJd8ONZET+8GPJQFurh79Ch/HNhWhNrwG
08/hCIS9OS74U2F642Sm+eAJci4Ec4bAZe6Ze6RxBa2Wpj+S2qBUR6DdXy/LWrLR
posBXWGA+u59y2fRyhx16QIz1xzQoX9yqaHmmm5DtLQpV8/sRO8czl7W6jW7WF7d
pIpkkeE9PbHTKfssRroNmU5i+l+P98yyimy/etYbbbJeU9X7uIozyWQPQNS1U7Zx
XYZUtrGQby1sRkwFOc4euWg8bGllvg/Qpo7rKTE6QuJhUr9Rpo5QcwfBzoqEgFle
grhm/jSqKoOTZ1lNUoEMIJp0Mo19kTaKo0R5T8L9WNjt7YEmZHCP8nERt8m4BDTV
f8/gKAvvpISBEickA4n1vdPlnhGZL5ePG4SyjLDonlrwck01LurM4846BJKWNlwu
znrwWTOSsH4knbtwn5yn4GLC5yxvrz+EXdusIztmmuPWa5ARg0VZSMnso9sxBptv
+oPFK9RhNfdAEOfHFrJUR2787n2zulV9l/yT9LZDbXeM4yMqYwgOP+3dqT4Lx+ky
tYKZSsS9IFEhxMEVcmwx0Jq7Ex0PudWatiybMepnpFOrGPCfH59wCLM9pTx0ewq2
PcH/rqJsehOrylN7LphXsu18pM49G5zg7Lg01ARUa+jg3z6WzdI0koChdB35brZz
M/MPEm7ZmyKvcWB+SdL5/KKd0GpTSq3DsPeZtwNBh+uAra3HHW8BYyByyFUebuWi
FUQGIbpsauAJyZSilpbF7qwZtluEtm5HUrLLmVcdfSpLyLGXgL29xo2WheJbk/wz
dhY66N7/bC8nGimkhK/ziYH1Nr0qM7QhTAYNETV7BvO77fHfXaRerhrDSSuwem19
jmuq6pzIRjjA+ogix45TEbDD2S39S6ElckT7s01658LOecr+z+QjjL8mX5TpNEDA
ig03noFAgUrDILGJIGTa96Q+py1vJ5CjphizluXx9qU9XwlR5k4I8k1H8eO412pg
FHY8Ye/IwFP1YcRxl5gFnSmjWT1c7WmWgepmeq4D44Ec2xkYsAAzS6M25mA6smF9
pM5IP3VKQiQ+KDTOZ2HTBi0ZJ3jPVdW+yoybs8ivjOV/GnGAicf0e8cGEtU1XkO1
028a8iwKtTVJfgFcvkbkAWpAXxxvyvVvEBfyB4Zioxv7j2zllDozogShg+zq5hBq
vvlr7Hvair4dOR8iT3L09+5+mhAMV548oRM1pog77iyApRK9SXco9fFdn8vtAYfu
T0lIwyEJp3rK/6ltQy/Mw6yYUdBN3pY0/s++Z8U7fndbEgOpDuWB05OEbCneihd/
3dIMPhu962XJrwJ1zjS32XJjMffEutmHbmLiyd6K8oi55zWm/w46SVWH3ewpD03S
iEAbZXFe/bJb/jFz4yagIeGPdzTf+nnwUcsU3QgbEUE3+6I1cZNPdcAEVBlYGAdb
q/h5bNrb+YBDsOY9hxMjvQte8Z15vhtXc7Tz90CgT23ZGCWZx9SGlno4w2NDEiHg
4tI7e1YTaozL3PJy0skTPPjNSO2IeJNt80O03S23a0BRlymUmwF3qlI8c1ahJV9l
TdF+GYGhFNW3Vq+jPTStn/mMp3Pwqu4m3libB7g+sb+kxtTs8I95hZ/kKmZ+vPWi
sLiuABloa5QQDxt/fbw4lwcjY1CpWBqu/OpBKfkZ67IiJQQsvrWa3JdmjctLEVZe
Q7bHm0f1uoAk166QI7Io2+3dTi1/9jdyL14NP6AKlwDNzmgcoiurKW5i/OI87EAz
90d7rDtAiN7OdYip5c4nF3RCy2CMSX1G6GQUUnXDV3YCvc6GJxe0yDbJO3NwabNk
tjpdokaokXzM0fAWVMgINe2FvwgXnqPTqf91C+Ca/OHVQEG1R2fh9/II1XZwXzw/
8q10Hb1X+vml1SCJN18N3Kj2iyszPrNLduiCD/FVqChkW+7v6LDcSGDhjqY/bOh7
9bayQBDOgkn/pyKiEpgrrkIwlNdLpSvAuqKDxytix/Tk7xThpeCl2U3xweQ2RN0J
CsPCphcCrRUWwAvvxyoyKzPlgOWB0UsMsflcaHdtAFiNG9zzmmvFvWjHblgJR6TP
2p18XbxgVZPW8RmUfPv8I/pWV+tr9mL4iqCaYODucA9MgTnG03EAJ5/jxwM0Pbqc
GjxUlPbrFb92NGMGMptPR1xdKCYAK6xtr2duq4lOKQNy6XMfRtXj9fUwDPQpWef1
XDxnjKjl3oSvrny3W01TI0nkxETVhQOF18el2kA8Ka94UJ0Tq4xLaTLo3vbBkyTu
99VbITRFNQJveF2PPfuVnD2XYFK4QSQZe0VF96z5LIMmm1PgG6qYL2vqPeBFZRO5
5JXN3bjUrbcqTLrG4fU07Uyp8kOc1oHobA4QoOlkQhdLwmX7I2FzcDb5sc/rQoFi
2+9IcZktDt3R1zoRzfOJpJ2yE7mmF6bJvTKXaZizpjVputQN9NpJyP8YOLDZGwzb
5Bn1f3bfoYWhz6RzxXvTxo76X0h/GraWjmba9CULCA0mcokVpJy8WO6MZbA5utSd
JPiE86HfhKAP0dkInoUnF0cG/7yJr6HgLS+vrp6VxpsCT8FAYFhfH+zhjwYjaiBB
QkKZoWeV+GscorOUPU3824HIVD9fuHMVy99JyHRHMxn3dRjZBXLRKvpCR9D39/O4
Q2QJQkg7fMYb4lPshAphsQiiFJFXzaApyybD75SjGovKL3LhUAmy584/0RdGeKZQ
uPM5OqfCcUJmbW0NnP+s+vODglRA/WjiXBQeDAv4igEyU1jKyUnNNOjh+0B8djEt
So8fDui3dTJhQbvvge51LAeXFU84+fB6cNVhFebNExo667Xy7Z0Hj/slWQ1Jghb/
btlekkva26V6CGcT+q1H38nU/CKGWPzMGhceYAV9eVADJDjf7+SyWdz5J8eetqAg
987AnT740ryQ300HZ4nqxlzW/63wqR2C8YxT/BKhENYzgBEUKjXUeU1TfETJWiOq
FnSLFvh3Y/s+wxpcYVDQZ2T21BmDzPfc6lWDvzZc3l3+pHIZbSwLfq8bm3+qTA5Y
jcvu8u6zM7k690BLtqiLcI30ZvwKEpve5HCFGT/LHVjHCPdvfes/mVaC6sfkHC3C
yVN1mt4TUS90Ex2Yp0aO+bqhvoToTlGBkWZ9UIZd+kauxT9NaEmyZGtKoialRnXm
9vunZlvz3iOqDunQik84Jhuv7zeZPate4z/F2fuOavqK0LucU1Gm9iNpiIWdOE6c
cuJU2jhcfNluiQj57sJVJ/iIiIqp6v8yEZ2XrPxPVxc4xqQlMQ6qpPtgMjD1IDtW
hbn8uOZ0M+jFh4FuLZcGzsBSqcXOD+glAC8Te9WNs0yYdBOTGTcq2UM8jQSVIDs9
X5tQPV+BCdY8Zotubxa1W0InMHf3mSAEdrzD1l7gKwVN4cyLEZGXen8CakRT+f6o
VAgG1XkJjCq2nuI2bXKKc6efD1eQSg+dN6V66YgKnVklW4HWjyUeuNMaDKO3XOTr
DxMt8M7BMSUrKslXxfpUKdPJSrsRjfq4Bor6lX5tDsUsLvQPAh4dkRnYCS+fGWfV
8kP+7dEB8Y2wYOGcoWucMzkvKMw88ZNHS2TasOqdNABVlr6L+dIy2ZdXhDPGmfBz
sBgF3+SG5liK9ChBEnyExa2RtQlCqbnB5lDpx7TbfNU6mq9p1/ycbymi4HKv5bEU
psBEvGiyMGYTknrYyW2R91ytVWOSpvM6g3St/qVtKd3n+TiT5E5OjE5zEbonYo6r
z/S8vUvH6obc+lwcC8+EwyS820ZbGhetcsADxBdqFIMndBDSwKpbBRPM+qvmjvmS
PuzIzA39ViqTYBORhDXYL/kKLxjtnfr8VZIZVrk0fE0OCn+b81whDFl/atVksjig
QHTdcP6Rc0punKPItKMwxV8CvEpDq0EU4Byfjjwjy2IESNBmYTBpQM+F3TFn7HeC
Ax8++jt0YsaNwYSS3afe5uccm0f+g5UxHlSrHKFpvAPBx7iM/gC1E81Z9AgIcTYp
EYi1JRHXiZElywXdavsQ+ayHxlUVMJD8HHUbh3El6wckSDlXv9Sh7UhNyYVC9B/o
885rQAq8fgd1okmNnb5HVGTqTA5MgLsaZ/3WkfCB4BOkSK6lizvLHmaDggwmzOiG
dTF1YPaAm7D8BLIorwVpwUYtiWODGvncUdNa0YtDsLXszlco/c1LJ7yFLZqfTitN
R80cIYe9nGqWZgOdbxFryVdUB6wAkR/re9l0BW3Ldk4EzHScn6SbSfx1CCAFVntb
eCKKroQaquoSchic0IP004zDYsYhwm8IeZNQACdkhU8diX1uGf/vEYWOOMnV218F
4l97T9o64jNO7yieEnHsa2JgVp9e5ZuT+1rvF3aomg5o57M479Gf7j3xQplUlTks
wQi0PkuKqgTxyb+OzXMc10Lv6NWKV+JBomxFNDTI5l2Y2aShrSI1n6QpBGQl+CAX
Nm95OnfNeTGHnpb6Rdk/dISBgpMB+jOqf1thSqSX4zxYyuL15CI2/W06vMnV28Hs
uHMfmJOVMpYj3/ftVldMRUDCfznUdNyh7HT51qMq8morNUV9K1wmnRroXOHucUCg
mkqBz7HrG8J1L/b+bfTWMJMSht6hCUzVxtpWp78zl30ohD5uql0UGQQpKhPXpCUa
4npq5kQt9azIO3lkwFZXNSwOQs29s+zSRCcUK710cQYyGaMIQQz1VNsSQnAR+P/k
0k+3OIieECormI8fXu9m9M11Q3WafvhrDaEqgMVcSCXG6ep1sIJGDCGWpIXqXjso
hAbkg8ErBuzXX+cK5ryMHZvxnHMmd4QE8bh9CpUdubYNrxh3xfNDseCHtknHcCCT
fNdsTKa0v18bLyyx3Ndd4XUTJXV7oWBD9tKHinWqU5Yhc/RCoBtDMrI+5zjvGqXY
rLGFUkH1E8vbYLzT5iutL/sVMlhxfAydQL0NhrKAKAZopmmvrC9jk7CRNZxSnsVp
95jHOvhOFwJACUxBouG8eYMwwA24rdH6SnGxh1sc1sKyoHsn2crL8KxQ57hJVL+c
CPUUL3HsCpXZW1HS/mGAIc8xXRehw/iYrX2wyNB+d5mKIJmdm2a0wnSl7G1L0CUv
VD+KGDacK4UySWXZUr1xIw3k+RwFf/pBWJRY/bQeBk8s9LhdbRZk3VXT9sYhgw2b
uhS6ydYXI0RUP3cfAFjCyXLGzm54Is4npg+Ka9nTQgim798qlAB1pg+50KMICMkT
JcoLrgsaA7S48HilmASdBdkL3mp0s0velUl1JUddu/Fxn7Cn7xhKzAXbZXb1ldAB
s5poiRYXmvkEF8yQBIxHkxbzgTjHEMMHY8qbC5fYwtpKu3o9U7YjTZ051jM/a8/8
6voPSET6E35LRWurqdvntApj5yvbG62usjkTzwWlxaDKZ4xybZgq1BYUxPTxq6GZ
SwkxSn73PNNCUHYgg01qIReSi6PmE5viyFH2PkLJg3sk/jgFrU3BQNqG8zmfNrl+
D9ATT58IaIeS8Rhg2+ntu5dstKNyxQnaiBcyfg9KxfAL70tsNoA3YacXFFFauuYT
5eLvpLkK2kpluqKOaqH1UFe9L8PKCVzg3bAhQ9a0e3sybj+MjTJQ7FEoJjEJrAXL
fBDsaPEhVsOeLaXjP4urzExu1qnTZWDdhWvbt2Fad5gVJvmpkPmFzgn+WkGE0XLV
zHXQYpcr3tJGbDSayJzeMrXMyL9lqPufYsryzZwB8jMt+RDIrLPJZr2UcRCA5SF5
GqhQTc2rnT7Lf3Apmj5tRJVQ7kTLtasXHabN9vu1TDV5jvpz9yZjl9tNLiJm/7fX
X9w4Ks7TqxAODp7fjCgaFejJsHrketk6qT6jEIObY7YNDjkDOQQZ2LpnsS/upBOu
8wo8EySG6iQo82zp/7EbRV2GWwDcAjwxCXxSwLsKLXvEb30VlZ5S3kyQ+XH04SC8
FbWA+1hWLr6QPX251EGfstZbZFVTEtKe4pSNw+/PQDRhdM/XklhZXd6VNIKezMHl
NL0pohmPL4wirpBbHs1V3ziKgjOeBdYpg8n6J8dUY6Tcg78OLD79Gs66Nx95qhZj
wP9eGdH/vFKDilKWoyArV8rmBB07y51qkC6FDtIW8+m0PTwJXXTB9GJvI6lGdyJ4
WzA+F+HxlEwjlqnsAhhXgOFynrbsLdRmG4nSdyGu6NKZwo/U3HuwoWFV+z1eONwb
bDFl7L2m9JNzaN7F9UrjCjBViMyk7dMX86jdYliX9jLljKP2PpWF7X+gecnKIsXb
YZf5UdWlYHfdz9v8yFOPe9FQpAiAY+jGQomfwDJ0NF6vy/bCqZmNmhLLR3spV5Lj
/jsS/Rs3J6eBR3Kq2SXKzIE/7bX7OUXyqtNdA5kGlaoYpSwPw1EUqG8jf6SGFeUR
woS0SEspcPj28gXgJDIZFL8AvLKGEUfvVRtX0dt43wfMr1Za6CfFXwgG7vwZ1nQ8
87xRRfryPCJfHyAoETX/Gn+RqQlsshTiPmnhd8DPWEdovNcTSRDxAVuqbfeZD78F
HIHg6cxMymTQ4Qzxah6fldZbRCs5nC9ZXS4i4ck8BweV4LCBszecG7LwnbZPcrJZ
l7DvfIgy++Oke5LeKWCdxye5ZPUx4aLGfplgqSxpPBSqqUv9RMxLJRALhXM6vz49
4Zb20F+ICK3QAzZbecgU5hACViBdjE4L7UwWTH1QhUqLLUSD2rGoTzcuS+HFXkiC
YExr4rq/UNtH0SC9JfiDHan9ACTi/BAJtEwUTPHL/FD/RY1R9K8bHNyiT/BTswPW
HJrFtJxzB7rg0Htus5/HqN45vkUUBpEVhqEDwyLZamshlPs009Ob1LEnb4V7f/rN
zjqzpteiqoSL31yC9krofkaEulCB1Tmjo2vJ4FWdS8crkCaqziVaAa0UGXXAD2Yj
7RuwFLnCfxi6iLeG7NYcwfpT17whS60DK/FpbOilF7FkiG51s29SUk3kiONNERtw
31OyRJvoT5johnQ33OwWiQMXfJcioNEhgjCKUGWVrGiEZTqs/QeGfFToVmg3OHEz
o2K7uv7GACADKPlvNOAX5AgVddfjzXDe7TES7YUEnH7J/HzW1NpV4gH6+fR+XCD+
eIsQxsy1VhyFMKGPMMuDqH5XGIv5pyYcEfkRLfdtfqsmiqIf7IMY+Q2xX/Zhhixe
kiPMqH9+8WcihJ1CBwTdlmXrx2CzZ6XXbUCyZkiufMuFKiDB2+BHnA2Yvi+JZKjY
Brm3mZPNHz2gndgKfOhpfAw+QgVapwBOJN15OdSeNIfNk+for+NPQNTkTAwkBjID
/N/PeNiH8zryzsaco3u39rkunIaS9FQMFRV0UD0shCp/XYUWCTMRUSdsBiPepSE2
ZaNzt1AyemP0AX5gvpUl6HLB8D2v9O9Q90AVyNr78nBmI8w+/EUIQ2yL8p9LB+7y
NZJvNk9Vc/4Nj+oEnaqmHnvpSH3F2QSts4tUgw9dFArG+x8Ycu2sXRkI8/fiwDoy
q+BQmVynghl5rhimIEHeghpyCBXuFc4808Qq3d9gzYUUZi3CKJrRihG1bNxNSpr7
c0O3DLpB2X38vDzZ9Dt1gp/j01bwV3idhFPjZ640c94hiTa7zuAB63QIp6gWtVi5
Nj8crqb4FVqg5uKOqhOODtqvMT1KJtOdna5dV7CNAyz1ASzwnnvHC1gHVf7S6OoJ
hIei8F0/z0voeY1VLqaK0koojoA6saH5OdnnX3WJ/UBYcPowndV0sHJ/BeNgCkcT
E3Ays0TGC0cX4Ld28K1FjiQDco/bzU6nMQl/nHkB6YLXcp9AgTOWFCgRKAYxUiOT
hX+LVk00+TV4j4huAv2PLbpbWYCSn0pbaiiqp9Jl3e/JXJZJ957pWFBp4zrB+p7w
JCRojbllX/SwPGUYwtGnLNEmMyrGQlB91iWIBkFuyDRDF8vUA9dFc7JIhCbPSni8
/9elrPpYmtOOi9ko/nz4iW7ocRRv+HmGcJg0vac6VdUNF4RHN3ybe84fn0ZPjHuK
KWyXxAdcREI69nmcdcnlVuoYJqlsHsBtO51HOn13jwVNn1DTeUEdV2O8XJFKP2ze
5WI7jB8Lht7p99GP+XJoUnzuUGlRodpWf4okdGedrJtWoSL8mrDNe8BWB4K8VwHP
0uhtO5h8jvJg30VTpZpaLNX3V0Jx8EMBV7d7Jnu8Nif3FZnjD3XqZ/l2La3g3qTU
rh0XAU/sPS037A/PnaUrZ94c82ZQ9h2xvxVCgJpCPteeHHj/VwETy1t5z3hQTKUU
pGGIcf3nxPm31Vyxy7LsIHHkgt0bnTz85ki3ofXfYOKOGfTiKXhsQJ09gDVlOdzS
3V4i8n+7/6qtZNI98DpVp9AltRI3HXygVb1oCTPRr8ZYckycGNofuUOeySlw02N0
zqW/26hjNkjqwQ4syVUfVHGUE7ZAesTahDnvrsTAWDG6QKIrJUKOsFxSOdorMsgX
IDZVO8kkSbQHkTr8ySyfEk0FwGmXt4LaIIo/BfJ8ERIRbmxhQgA1iX+I4fB3E78Q
VUJEiE7vv7ZhXlY3qdbNplLplVhf9/aCWwMbxl5DMSZTLo9yTi/WjWs6P541yNm+
qkaf5CAu/jxjotWfDT4CBf53om7psMxGkSUHLIUKVoB0zwklYhB/dMJbUM8rcvLj
mmn85sxv6O7FA37JWKov3gPv5sVFiOD3XtIHUMnye5mtG2df/Kvn+krfDz5pmgZX
9xQXwReZXKx7qDruoLkiVRt+E1uIo0Rftk+sZRY41Zp9AkA9aG/POKwOPh84PwlG
/dXNDRCT380/wTWSbXZNXseoDz4KfaRzF3NK/L7HkdWfWnyONq46ZlpCUT5foLWv
gpgbMSKjdxSFCuXgKOmY85hMw0BXcKjUvpZ2bneVs6XYxX2SeAebn9LL1Ji0xH4s
zeJQq6mscROszE/fav/4Dqd6+07HJBWsQWN9EkdvaQsPLSPWpvN3z6dI0ICLfxF+
iWJLPP5s8MsnSraLkA8ZSpqW7ChetDqNkSDDlwjakm7d0LCByQOKcm91YyV/w3wX
gfln+FRQB8DKUT+VszyT9739yAZU1sP3BLGC40gaYtV4PwPpeHnIkOvn7aHIg98e
xb4O8rUqEYufXgh/sfU0rj9NDnRdob0vDKPNTU/OBquEjWVrI/thmqmdMGjrP1jx
2I4KcfvfpMKm8e+D/ohs1oPaE+8DaN0jS4l2kv+Ur3a93tSe4PhmvBoJ9Ub+ZeWv
j9hHnBmXl2kkoYcfE0ffuWxNtFFdmVzII8nEj/7p1srvmtLfRb9+VG6np5YrS6Mb
Iy++NEu0ISfhrpzVxNsRDEbO8/3wiXr9zm50R/9MSwrRjF/ijhnL6pL3OqG1bwqH
RnkwcVhSYHUFM2S1GZDdKz79hgMciCzQHactNBjSM8oQwWnoLBm5oZW/6ucbJ/eH
iDGxi7f3NzmNeYe7kbHQv1TOSZl+rPbSYHtJO4ubNI7iK8xGMJ3NmGpg3MBxOiBp
C69BMaCSuZxINK0MruG5k+N4fKXLLKQPQUWXkttoR9pQi4wRdfTagj8a27Q3w1Wj
N4rqykxbCJ7haMDtXbOmnxXshqyL9nA6uvmQJ618689w+X+ky2dxty+WK/iKeHqt
5iwCMEyeJ0eomkLl5pp9zMUhMbzYEFTagnRNjeycf0tCe6L1CA8nQN7OK+qd53Mq
e0D/6F0jGxPN7twL2gpWrGELainnto1FMXAxfRV14/LtfuAmdoqVh21YB6+ngTM0
afj9py/dsi8vvXKF1/JxSSWFT8PJ7hwd2cexANutKYz0LaSkCN35M8GOD2Mz2HVv
7e4eUGKgltFIgQHkr1aHB9r3ju+66ebm+GHe5uJw6nfjIjRAhXvnjw5X6xc7y2QJ
zgJ4vmr4ArTINMsFp9WVwlmK0466tKsxgALaPlv7O41+6D/M51tIdlK5VqTa2ehi
R84dBz33xbQvs9LTn3C8r1QggshfvjK+hMiKP3tX7+4YT0V4BmgJ1lUrN8msnIuj
S+h49lOcLV/iGH/mX3EM8dQYVlDbvY0HNLunLsldTWBm62badA+NFZb4JfUwgV40
BDjkpB3h06BVvsPF+3PAsBKiVmHMeCsqw02WXVVTv8+j1qSYwE/KBzcmgXoCZB+4
W2BQkPfd2iv8mX9YGZfGI57P8HASvelLvGdq4YH/eFlSFJXO6IODsM0SLP8NMjnb
kcXzeatRwVJOKOJt50Vpf4g3i3L+UougX2QgMsoq7a9TibQtWAU+aLDKq8ofM3sU
tx0lcy50JKmgdBvYpQorQFCMZozYyH//jxAQEfVLXBPFll6qKbxI4CXw+tGdB5sY
pCwN3CRNWs+3MPugaJ0Dms6LAG6tHQ40sf0N0Ko0q4OWT1sv86FWt4REYkg4akrG
qg6vTbUrbsYQwBvBQKrU4vlKfxiVU2aJXsGGZdHn1B1fndxSAsO6sY+F0GOqTQOs
ZW2YeqhqhEowWzWX7uawkEL8Dm6PeKD/1tnQOvGnkowvMvayuWOf3IWGMkqjPNZm
4axlXDZXuMgLM6GDRvMvi6DPkzInh13JUwhxCOPNUnsmI8Rneca23VGip+jmlVqS
SdiSGNJ8XfBsHUHyxyfn0ILldCufqhs4yUZffBue4iVWcs6uUmXHcMwdEh4pA6UW
aTiukNJhobthPWe1cKGpkYFmTjL6Jsf4DXw1SzOZj4JWEMoxZC8Mm7wuShKPN/tX
OVEhlLF65Vj/3dvjjHkKbqzvRINpGz3t/B19TjClhehuceV8oQYEz9ZCU5aNgMWT
kvZm4PsJn7x7WLy2dxICmDY8zvIYQxMINM96Gt8kLv08AF6F0pEFZZUm8F385wzr
XLNtf71duMS+pGJvek5zBptim5i0gLwxN0iBpS5sgVVC4iuzdJpMcRRIOzDS7P7C
MaNxx+Eh6VJ1sX1SMsJ4GKx/o4My5jkzpaxUXDUr0U5YAJisALpI0n9rRe6PxyQZ
r4YTDgWcUVNMY7LYzOCiHwIJcr6riQE+cuF4blNq0ARq7Yx4DextHJFucep9sM5Q
P18PmxhuXWipvTNnSSukwd57Zrzll9ZryeLsUrokXIuRtjYJXW+cMNpDO21ElvEL
azOlFD727VVAJAuliAxAL5DRodJjhb+xp/I1acsKtiKUAWF6XQq5g9uWtJqcVGpz
XXf/BWfupYFNFOhTnZRh5Pf29Rzjg3x/M4+rtPSnvIeWvk5gjjWb1to2J1yL4cU2
VYiX0L6P55akPU58bSudTAFsY7MEkiePMpX6nRnJmpn7Ydue/dMHe5aKP+NXqZNF
9O6ydJPvNfbvfYsqtyHCYPDuTvnYv0JnXhhXFIwmjd7dYcOhOq3XDzwHb/v1W95A
EWq4/8kunxa0SriifJ9uUTgsdbeuhMDGM1+ZcqCkDCA6IjKGGQcWvJ/Kae1BHTM1
Y93OOKOjlT6d2zoehHkOdGyldmBZvRvJyIgUY4ScDLKjwdk5Meld/QnOurBzfVyC
ZduHbw2nbfwoU4t3nVNzmYWkZEgVhQ8CT8yj6qKpok6c3dXXp/1qYYCQuAqU51Gp
n0SPtu0kJJ8925ZTGMYJy5Bc5YJcTRERTsKL+G2yg7n9ZSXRcFvnipPEiDvSlxsr
TMINgBTSa9T2D8fIinDKorC8bGmGYAhItnRKX1155fN1gaQ2nGE79UCh0btIaLMc
NyGT5bMlMaNdlA+6XoXvMIz3z4ODMtOyFTJJ3MIJ9ZfSmKZHO8rrS2gW+kGf4d7n
Xpy4y0yYT2k/wa1k5DtTI+il+E3fMhjFswkhqVBskon3h6fCtB5lKNpEQNO2a6u9
oOsgxfdHixufM66YzyRD+tZRqEuUmZprsjf8rxqCkoDna5jkbzLRGCr36ia1NkyS
QLTCNRS/RSfvgZiGSy66GAV4qPkYBmnTkINmSxo/4/YX9mtpdQzQRBSnQUVtIoaN
vCDh8sUCgI/xUfMOtsirFVFZP9Bm3ApiPuW28TLViXphxQX+ZtPlHOnnhLODXTfb
OQogHEQQMxuGemHNkprAakdP0uBK2P45mZKyj58cUF4BYI1AYVlHDpi2vuEGtsQM
RK3Hj45u5jNcTzBs4qqxMCI00ljy1VOnytCocTheNDOz/e2n+OF0e2hYSUyZwJ5x
haGNQMo0AhOPeutWpiC3aF1HwVr+pDry3ooiLK/MIuIIgB1PUqb35xx48F7Ul0Yc
oLgMZqHfEwdWGBafPoFZYaa77sIA48SSrOm4tu+SSuuOBEOwa97n04qzGb8XAGzt
uiVeJg2BdX9aHdkmn6wy/UQdKzrGl8n0mQwNgHF+NRNOTeeK0O9q3PwBnrJjcIGL
jel7JWXcXS9FLZbObTwyfxsXIFfl+tzI+rWrpEC4NeEfynbtYF1fuTDosHI+TmFL
CI/tyrta3OWxffxEAVkvQxpeX2uocAp9gZUTp03v46iv2BoB1pEmJHOLLUCFTESN
ikE6CzmfDdFS8c6cgXyZjY+mOxpSIe9F+XqeHXcgD5HIUs/z9hb8z5MejSE/kYhr
ChQToK94KEq1xyJQoWRCQWfN/HbAUoWU7yTcTPAxsrj3SnIqAyrx3+mC4ejkGOnp
BWu1NyiUTygK5LODjTvwEV7slDw2TRU1BwhB+rjUkfUzCF+A3NcJk5N1fUdtMAh9
zaeOZIAAH9k1tD7g/q133zX22HUfrUNFhU3S/nHQ0fZf+Dlb8PX6pkSG/zYuqovU
xecVlAiG7GGYHs88nYJp4QfpDoa7x3sAWO34YbKxJpZvqB/tzHTTM21GUUZncgVo
g/6JAgmuD1GJzJW0idSEu2Z8HZA30VGUdeX7PHX64ZJzHatfFzPef8fl3Mlx8hWU
dSsA+8TQMjL6aNbH7+ztKzJzdK/RYqx96/pEb18++AVm/iyQn/RHpZ6Rs3A76KyV
quCtY20elpdgxhY3ra8tWYXU4IK/43JSgEl4jL6av8Xdb8TfxlD4QNdgC+LzSM6+
1tUags9kE2aMx3sv792ZUKsSgkfQdkMkoTEWNheoWH89GSjgIFBpElxtr5PMAcIq
5JmzuKWI9YXGWEDtJVQqWxB1d9TZAJFntj0W1PxidjD/JNc3hKpwEjaJ9DrZfDkI
gnpJPkwbJOIerFr7rqgz0Zp6vlSMf7yZW/P6u+uHL5IACeI65JqIPKU5rUyL3je0
H18faRwj16vLZNRolj1hVwPyYT3PAesfPI9ICNLm6in0NyDwHBzfcnk1MeRPJcIH
6mRzVGQOqD5aokFe6a8HikG4ryLppawKRI16X8rn/7HtiZuyhfQJH4AXa94wdGdh
4tcAq7jfGZEAhKzcYbtgRM4TIpCW6KNRmM05x9I8kLA1E74EtzigAtQKnViPHFHz
VG/ED6Y1U+xwKBW6xsY/8T6DBt/jQg9us30uzHkql3NtUYa0VNykxWAg3WFlCTqN
HHacWBuoyWn4BrYg/7KbDXCJuLJ6avVohh0292VQRJtA6COHvD3hfAlctFjSnjp3
7bfs7C8iXfPZDkxm/WJRjey5PeCKcHMzyqddVYCpBL+64NecH8Un3jaLmSSZTH7U
X5yfohfAs24Wi7X7jRkcxoWnWIl4vxwE2jwqFlIhxbo6p1Ff3ifLftrq2wrWxygo
Jt/UZCf2GSv1Qn212vT3FlI4ZO+sx34uAMjFnKzHNpoM8p1Q4z7h34poU0OEB5o6
R6b5D8SIEVfjHh+HwV1IkaFLaF5V6mCL7b35HpiV1jBCX2bEAdGA0tORhmykZm7I
ErMJvZMdrgubpiMPrbQNZEqykS2Hx8neL2u3Xyy3N+KQgp5CnfHDb98gb9Zbd4+7
49fwRZEylSPsG3jlZ4BCz40VX4LK7LFwxZmJSXVY17ofZ/twQVFCL6ZPMSFrjHZ7
ow3VMsmwHiBIZ+PNTGyITxvncLPWYv6EMfAVI+MPMDtcIJmRZmZ9PNpahCQL+EbP
O9TpeYFTSRrPP5q23KvQxLVNtwI3pGc3st6qx0V7w7ew64hQdL6vITG/OstSFjEY
e+e6ZopaaekvtB0pg06ASo8Fe9riNINMuy7+8+zSNBUTHAPMcpDL4VAHTzSr4CRS
6AMCVdcWarDJp89aEdi3Varl0gkoDHxRw/uy2iOu7hWBy1CM2rCsvTKO69BFuPHN
FWPNGb+wsvBiJMEN7yzLBjLgY/gY+Vbod+nQCbQsQgKiKygS2+afxD/h5SL5L2CX
VXJnkppTX4HA2Duz+Sd+mqbU2xMWcAe5fWS1TAKYNNT9M+thKi7VqCaELx1lUFpu
FWbj/9+TglNH7qE+Dkhvjyp8h6bNP3zxfzNRP7pOPxpa+LTRNo4qPaaQZVi1AT99
h2iuUanUvqUV1RNZpgtieM+a5sZUWrNXxNjRzLrOKNFWcVO8H2+7dIA9h5weMjXp
SKw4WExMS5f4SsuV9Q9DmZlG8korc0iP002cB1ozxvJ/tgTXzTyzaWls+/OjJpl1
YJ5AyBM9bRdwmNtnS5p00hdiZ3lCalPKu5ZlKSVVsbP/rX3756toEJOxmhxhQOIM
f237LAEvFy0yGNz77vVcmPDRltqMCVyQOTzfILABZuaQENSzk8n1WTqEh+hGfvAj
WwyLVLuRokysNAUZaS/R2516gpfE4+HQxYw3S8AB0EeSuPfNO9Aiqd4CA6SaaSUG
Xt80v3xj5BjJVbKw2zeTuj7Ia3IwrFYmMuwBBcq6GxH4+Dt5+1EIlX2OVdcchts3
rfr4RWg0aqhBkMzc2GFYdOF9yipBpuFLup5x5WILTlBYqaYuq9lJFOh1JCjGXHpy
nBY9FZ0KyY93gIa4EJ34+Yg9bMWVEMfdls8QtuoCYR3+NA0Bxuh3442SCs1we24K
Y1O/7hX1JIf/Qwxt6ImUaFBksiJhK6Z1ThoozQU8dO84GtqiiX4jML+0QN+LyLhE
w/cta2H8kNfBVP7HUl4FqCa7zt33NJeo+UUmrD/ldp7B4xVi+lpZxa68k1nzb3Um
wyl4Wyejf5SS7ExQpfQVNC7jhCKOl73W+7FxPz993WlkvAm5P9WhHPGEhvwcRTgQ
edgi2PuDINZF8njmCJESHSc41R9LvmJqeyY1nGf+n4O6SlkH/xn9iUHqwSbcSx5/
xS1TiasOeyLGtWtE/pvLFo6GvPtx9Pflmu4uxOj3CRECk/Fl87ZBM6FMlplUz/BO
r8JW4yxyL8HYWswOyHosu7ohBB8rIU9Y4PttXh+dP6beA/guC2oP9SVr12M7O6AA
JFXaDNFnSv+rciaBmepiohb+ewEejSQGaEHEPf4vosXhZydGB9jQBOPv+V3gBcMi
qr/PVXaucJzit6/LD4FPLwYYsM0ph7lMg4P+GhhxiIHW0auxcz4baaDMCaTbAJ7B
tX0ErG5jXxwlRVLCathBbQwLZG2QNFBboPMOUl1kzUEkfwkgE8tPn0WmQVjSzKVu
9AVCVXLDuDJa9ke0Hm+C3K9YvqEXOsNIsJOPLpPO4s69+mzk/OtfitUW/I+1m/zT
fnu6J1cVlEhYSWDHQV07UntjQncsWmAP5e4pOksjbytbm3nlS9CGzmVhV+aO9XYo
7chBm8KGGq7sr2+PCsWyAPdTunaPQ9vxYNks4GFYuS3wJcMZQ/wBLh20DX6cntjw
ud/AL1Jvdhiedyd5ZAiq/cXIJx/ApxhQTE57iDeDhtHVK9+bJTcDoi6JuC3k0eOk
yIFj4IH6B+v+OoPMQUwlaq9UxTqPAeO+8ZeL57Khhh5y2bsEBDQJ08Rc/lHr3R1M
kQdFQekR5HmdedM5vGNChUyvJDlCsXuM78cmpu5aOdN1OP3UMeDXjW1F0sml8Sjo
gLNKtaLEWbs4IFlf25AVIHiyNr+SX88+53X3eyf/NN2HRYjD5+Ufae3mmlXsggxS
gSMYcyAoldZbFEaacmKJMk4NJsmani/cHQb4mRKXS2h1qiOPW+DiszeiEEEjK8LH
EyE9VWrIY5gy3fs7+xBdJ1FVJZ5/WhcZONaVVQk6Hqgzcg1ki/3OZmokDhPozAoG
6ppo+2APSmYB377zezDPhTLGib197NaLn5BcQ0Pm8YrWYKExx+rcYkrs3SJ20xq6
u1YDD6OQIdlPpdLa+VuIpYGH7dXv5Nu00Ya9ySxw1n37mOj1xa/paBYRI3rMGiB3
ekMQqqP+qv0Cs8ebr0zt6voQEC7lyrdcZp8UMl+8Mb8ra4ZTjPep7C2DUcSPRuD2
qBQwtJkPJhtVM2aVfP41WyXNHpNz2bXwtLlYVdNW5kQvFaKyhkLr4OfYjIWLLtT4
Ku3PmveTpW53wy/fyswU7lSVgt7raPSXRehp90H57j8cCdazQzK5beEp49tZrDvK
ec5goLcyswl67bJ5l5PqjYawhsGgjVF3e9dNnCUhLTMFNipaSPB6Gs2i5SAshRlV
7FIdxos7FVRMBxifwqWIG2MvZAADd8/IDl7kBDlcLobTw8KcEDApdW0pnDRHjAPY
s5hnwXr2rMUQjxMpRAE5T5Odau9/tGnPhwm2cxoH6nyIALCG+nDJyG7lRzqhVcGM
8sd4rz3m6OzH0Hq0hk3B9SFOXXUHGEwsCK9CNTOxU7+ECFP3xt3KzhHmIIWl6NLb
rrl0iCC9tLZ4O/35QQouYqJz8cOP5dS/CknBLZsr9n5BYVcgp+s7TGQTcO4x9sf9
1Fgi0hCiHN/uqKHLJ7YgZ4HrqJrPaNfAfpatTwe30LKkcbo2G2v+vclWXhnXOakc
bIuG/TsZQZMrSQCCgv3eRsoL/PqjBnAuqF5/xuFWo96hntkVyqq9T0PuHdexQBde
Cbq1C/sCqdAkr0AtsT3SZ2bfJ5llAqWrJOKsJQt8vzjHbQX1zFdiG2uYixJEldse
ph6jT34LjsUSWCsJkzZQtQOsLI2FRtdhAcwW3F5aeifs6g5SZvAM8S1Zfzd2bISy
/EM+MjlCKMxK1YAvK7Xu+ZYjOIx2XnAGjVubs6f6rnYHRMKLi8AUCBTXtFomwdIv
1C5Sswm3TtqVno/jbjow95/hvRPDnY5I4rY51dYkZ5v1qJOxOou+niqy1CkK320U
6HyFgUslpoh/0OT1BDG2yF3IxnQslN3SIJ7eRWuXXCLX6pcMbb9sPsQD0r7aDj2R
WWa/D04KV+xdJpvviwcuSz4daHIaoSZkzdu5dRWJxzeExTkGA3PivY0lMDN0Y0IW
QpGNVv+qykTx3cuxWuwcsNM2YnHlRkYdXQTGrj3nGVTk44ReBRD9pdFMCFYZjQv7
9TsHCOh4kDeh+LY5MxBuh9r0CO53AgxD3G6FUfdDtyMCwcIEc/FPzIqgBAeCEI5O
FTExv8uvlHE83OhI/RH/E/UK7cDOFvWhW4S1I5IB0PY7XZB2NZ354ujk8q1S84Gr
yszHYxtF25aaVMTv8d95LWXZzLqeNK/LAoZwUN1yi3vlW+rEIDHyLbmWjrnZ9BVo
Yo/1Az2bk5g5ClGPQbm6N1TT1OewsIOzKWs71PzvF32retGA2ll4lci1I4Z1rJ+2
QuYtlGEvdXqZp3LLk60YIZfnHraa0/4VSWeK2jFZmi4Gg2gA0KgOAxAqvGF4L3a3
xN/xoOAB+tIXCkkIH7xyBS7Z4fhrytANi6NALpjgBb4pa4IAoCtfnnjncHNOYDva
0D/4FCXot/hzFX7naCKAIXQ/0DZt+XuW+V3jTVY8aRfoHN5MGE20VihhvDHIL5gO
bW+IsB2M0M+tux4D/dGDlPXGizmk2qPh1jhG9u7wpHnJ1jxlg+MZ9oNNkywoLuiD
jfj6y7DyYUHF3drJiabzwI1kfyspbx+eMjn8aE0MdN2t5+eR4/oQ0AJzeWvrQVnh
dt9SYxooNhCmKTZIA80LSn/I7dyNc1cWTltFhh06jknrbnBuovp+MY8rH02YEtWZ
2IqTRuO/kTISzeRKExYT+ZcATHzQSPLX+Z7JeQMgI5Ctx2q875g9JIjzwUz5p9a3
z1yPXiuCaLdkh43xELQVnsHszWPk+ZGMyH9zVObLlt9h9ftrhoxY3eLthxNTq0G2
owGmhiIjk5h3m9zdJJ9L5LbtUdWuewF7huePcuY4MdsuKw9fHZfgZUHjIxzoc6n1
iWrgwSBKxxkjq0DoVz4VJmOTIMvc1tbV6mNEp7n19cAzUqFshB5n2XWb6UthAh3p
TbESaGmP/bsAJBGtSzk6rCkZPv5Rh4C9JJkbCDeprzopokhgMfO7P1Je75Av85G4
+etHgUbi4lkMhRaseRBGWIqtj1/iibmJNgplTGqm4iPNZpcc+OuuVbptvl4asir1
DwaUmnbgnNSCWTP0mfbo8Zbp0OHOJe9bK548mAoMLbQLqdWoIOEm2ZTLvNjdhNRb
nAciEHAtgX67GWFYG/e3NvC2j8V5HF93E2k2lmA9vdsV9UPl80DLFA2y8e2FlCOE
TDWJJhhdux4vAKipJkQTzoHQwxHzQlkXOF4xx6kidXXceBuzoxZ9sdfZm7b0NG9I
BxVsVngG/qdtEFWF+Y59iLvpyCoVKkVrh8p0cNSx+9jO/jjF0eIKGBv4Hw5q1JrS
QuywfZE1QGTxWvTf9K9mxQLG2zzaaH1h7Cnnhc7MdoeVSVn+5YLXEvaSrxVKp5w8
lRgv7mvA9KAy0sMb0MWII6209uxGO0all5/De4Zd4Tv2hVttgwk5FqA5kVOa154k
yhwl0pLklNY9c4eKP4V/tCmlY/MdYZw5U40m46x7jqLnmBIhfSXMp6AO1vZjikET
rMvQ/RfNwl5/r58m/DjfeWdq/DFF8qb2uMPLKGSEuPWcpuL8W8NhS1Qgoa571tPN
Xg81MFkTruZva1xAgqAj03TQ1xWUF0V99yTPil6y+2ojB++f44bA3gLXT6GqMO30
Ulnpf2AFbSdhDehWWWhYPyC9ylD/KoKM+/DZP4H1VNf9POBzj/GtXu1wCn/XD+J9
9e+/Ub49udhPSpcPNP5otnbDPNkwMqVSuShrXShfr4uYX+E9Utism4NuHBLi3xn7
UxPLzryIlGmQ4zyLLBrgN0lFRJfWEbXvy047L+URZc8srKQcoSiCWwT5PnuiE8o/
5cIJXDc8YZbfi5o4gOMhIIpQNw6ThVljP4gMfYPFz4YiT78DtdD8AUOl+vZc7LyV
UDsMVM2k2NSY+Jc3nME7e+ax4IG5G3DuMDmPe78kaV3Z6FEBqczQOJkGUXy5aT+u
b5qgDlsMraFmje73sioG3YEpzsBpFB/Snj3797sKrWoqLlirlnjOxqysjrOF+EpB
tA8Ejyw8v/f/iYN7Cue878WG9O6KKUPLSND7EmSUF/DAwGlaCEpDPCm6ldY/bFWL
6kuJXtdXJn1PiR3NfkRsV9R/NxT7Tdlmvrkpii5mAH/o9iXp3/tTfur2cnenA4fp
uluIzfJmyS3wKHZFO0Uk0GFmqwcSxqgKtGMaXNH87jtKY7kRIQLYRosJUJSSYN1P
OezVRX6ZULj4DbVY1Q+/7A3OszPW6R/aTIHQFzmeHsDto8LLi/1deYfosE0k+Glm
NI6veVxuPeLxbUbN5pr+58b8pCu0EVGQeA5+cfLCfzbS3TZ7S3cxjPWdINDuyOnb
+YjuOoAVvM2+YCkHu4gl1t2r54UXNTmJxb4eA7Ht8GkGDfdlP5lwkGnUHlfJqgLs
nSzMFmublHYcycURl2b7QPsrWr9+fq/sP8L1Lovq1pEHe8JWqe1iRgzE1HYJg2Zl
oImYJ4A7AWu/oMm0e/kgVzDEiGza1dEhLPdyXzpaNQeYPgS5n1LsIKRnU8wjS6dH
1wv4g+kHM5q4rV/iUX0GKkmqtfsBTJ5b/E3hlLndJdq+aeWp/dtaa9cYYhlZK6hr
i9hpzrMNWxpgIotM1w9ghy1YwIcrJ0wPOGbjALDBJnxXMrY2y/NOWqO4Db46pO6z
9KbJQeO1Oydowi5/N98Ycf7Z3I6emmGBfFQEhYw2JIsdVcje36N6SHTYokisNtO3
9XfEH2/hKR2WM/WbTxIzCTAMP17s+Lwcw6M0hFk0SUS0mn8hmetANCB/HUvt3+3x
kZrPR6WB8CgSGo0kL0utlrcuOmXkjr3JriULhVpnyHc3A99Ku7fbt34qvmzirMYD
I1ogjDqmjXOOXNlIQ/RY23WkAGargMKJC0wMjmY2f/ltnbVDsChOBe8cueU289GP
Ea9hAxotxm8Mpz3M1r1fXc74IBbQyI15hMpMR9LBwHL+t6CT+LyglAoSsp3SYWWa
p33Dfv28LKhdZW4QmVtP7XNr8TmN8upYCZlpAFc30HxuGiR8EGVQQPaeubOqCy7J
SrH6g+MobfprYZqgMOE8yY0Ulxp0ZlThDzdmaw1pJFz778Jq6x6Z6F5I9H8vzKQf
Z0BAdknEfbfaOjUet2goYnGuDGc1Dgj1pqEvIot6QK81AJ/GE7ESffpU4x7yzSfw
8INue9F8tuKLM3VIKtvFx+hXcWf02KbqW6h2Uk+YctCP0yIjH89mKUYQczVHArpI
vqFgmoBJ/Rny/shSFMRBYb08W8heWYpC/GoQbkBgwT3BdB7EyKGhJNOdBuczKFAF
7EKBcoB2cF406691XY+0rqmiglVZPIYeeC7kzn5aOJyD3u5EC9/APl29GHOdTX4I
TtcRjyjk7KMVCoOy2yQ5OL7i54rQWA2iBrT+Du2Rkebe7P2Wb2KOUcj26BDHR15g
o2fPRxD8DqO2ueN02i9rJc86XhFVsC+WEARsPt+lcuD+S4Kz8gK2h0tth/zQIsE+
QJ4ZtszRQpmjypfqct1jRPZItLKTLQrlutJd0gNH7234Dz+HM7UDwnbQ/tsL1Z44
tG1HQxr656niwsr6jznOLzX+Ce7Tjm4rh5WjCMBLoppmMtydDoCDExFZUuKsDJvX
cNbW7xox0bBU3hwkO55oyi1CUKrH33NCEgW9DQ2J/OVA5GDVGka4ruiRqPdxxLO9
WS/x3cmZjjIYkf3XIstgnAuUadM/aHOtIlH9hSigWX1xhylV6QNkZv5AAvEhU/nD
huuCx6o74YrN2IeNc1kIpOjtNG/fkE/kBWuavQ0foVHVNEN3Wau8KD6qCG7N28+L
SHAMTd9ISe00hsvvIAaOq1eYWJwNKcIZsxjZ+Kye4ay1SG5m1FwGVO97mbdPU0qb
Jo4wsdMUpemkGjtpXiXkHisjxm79yh131jzrN7chH+gBG+HyIOv2IsT3eKORyY8I
iuGqjGi1ivaRDNmoWceRSncMLjtE6X/8SVc6Qqi2q/6Tup5u/Xbe5ACPn/Oh1kVL
WRVdGZ5hy0CpiS/mMdLARsNyjWMcVVpcsEFaXeZz+xrX2vM7qxXfdPln4aExzaQy
8voY2rzwssC6DE1oETjMCiZ0oe1+JUnD/VPBWkDCValZ9E+c4RN1UookFTS+h9Qz
DzexMDVEGRXUuUfh0/AuYVdVDHhaKT1F7iLI1xixF5FEyjGiseptDlg9suRkN5L0
t3C3zpXFcyJzuqaD5K48cX0vQ+9Tzb23IEigpliYxsenbC8jcrTKCzbEJBQtdk74
d/PXDkUtMgrMRy0z4NlmAEn4nsce1KZjisMiNogOpu444EGZlXk0HI8oHFH1s6Jo
Qk1pfIDMFaQPacjJ+UUrZ2E9rl1EnsonU0F6zWSZ1utBbzWgIMF+XZsE4qA3GhsB
lKbFqkWjkSEKRC5M7Psj8Fg+USKS0LO6fZISKoggjQu5U3NQO9bjpJ5zO/ThRtd4
QRp/1PImLl1lp3oh0XpHqqtgPVgGIRcSzutw99f+6R/pjGRmLqWqfOrDGk2f+5+R
YJyUL55n4xiGEycmgxvOPAhEkK0iq1c/xX5nuWodOO+xdVSdxGvbj6qgiAbe/AZ2
+Ds1Q8EQGcmhH20vP2IwXt99CfNIDeRuUKg2htcnU/bJgxk0VJr9y12Pq4xWJpeP
L63JKTms/PXcKtM5InJ4ViEgsAkeDR0Q7hjMWE8I8iXAF+7wUZ9cDA81QCEu44/V
hftLUfzqIEafOt2985Oe6Tov9rCeCQjqacRrXyW8p05/hJFk/keqwPETap9/pExJ
RNWA+9QVVnm6rx5lX9A7ZHCK8yWbEFkFJzGpZXpMXFUY2KJQomnjZTW8GCdYj8wF
XZBsa5AZgu32pK4V5Rk768DjUSPClRuUYM0DuyqU9HOZaLJD4OzjQhqgWTPVxkH/
9R1t8xJCgo74OovDRzFzRI23q73yKhgIdb4Rutlbiaj+I0+l6WHyj+nSi8YXYDXE
ligZiDwU7IVH/uNURaS5N9cUOCtMf+Gu60fHyS9/1gRJNLBRjwziR3Ct3QXXcPH0
lTS37PdcUDo2+XjZl0Ua0kpQaCcGVaaoyuO1iEReccRqedtfdEyBrEnG61PrDcH7
Z5jWRGqQJfsuJwwxUEInLizc+0XkW1ALlN9kW3TNx59eRBZCArrEgxQbYq6229x6
40hopYeRy+leqUuI4jTBJQAyH+AX62gseHVZ/2/PfaDuEQcopgPNhREjivot4fsN
qmdYSUeX29I1lWVgfTXO2+2O+/l1VU6sRKVNbGyO6tTHVudQ073ZSOy2PYHa8LFr
KrLRQ2iSnUOpTtNUvgPxwaegQfTrkVW0+rqQbb87hUWBSrF8YY/pzd1bznDrhoRY
63DpCreTJUvT48VPcMJvAFE5LCsPbhnqteaj7sdCN6+h13Uf0jLmYUQJZwYzbfg6
VxluZPQcQzvglx1OHePAjE7eRYC0UwxWiSjoE+QvP6mgPv9OsHUu/7GRM24jb1oW
nc4WhwNoBZS3yHMBS1GfA5gWEYFUPc2luMORR6aMFmifA1iWzBzVsTeBS/p2k+e7
3hIy+sSAHpGXXxIdurg/qrCtH1TS+O78ApxfL18lQAwFExnBbb7LdeOeE/I12Vei
AslsfsQVtgDxjgUM8k27mUHqiAK5Q2NHfg3ehqZHxWGLkmBiSJLJ3Sl2OoKsofWV
AeOmOcdwRGoEs+VTRFupJmqZOwUbYoTA6XpG2Rxs0GMuo5SZARjo426WaS0UfOlR
xpMRiSH/VHVkzrMrOOck6QMhvnAdlix+G9PkBa46fHsIfUNX/CxzzPy27Mr2JU2P
n13Ff6K1Uo3GZCLyu12+/XcWNqs3rH5vr7mWoPBQkBTyYpSCL/+EZBRgqLD7G30Q
tB9Gcgjjgbt6i2s/zw2lRBRrInPSBpXWIggQ1bja7UYKlSduTS7E4ym21y+K5/us
Nsul8UU/ZIx/hvLqAHwFjfBDYN4Y7VeIqU+WwocwhCcVTpXpH9fvBjieDnIWfHkI
A+vRsgRooJQO6fwjtmT0P0KymvAPxMnYhqOg/tmgFic8YA9W0XE5Qu1aiKlUvYZN
rM9W9onipbeYdLBAdymCgnmY8rqVEqjznprHkLU64GZF1EumeDKiM2Y1m+QbdrXh
dHRBN/TPX9tRUg8km7Bzb1xeQxDFTTiS6e6FUonZUISPIOSYYSHRL86D4Abry/Mh
x5tZJpTNA8/mo4KE5AszDfGlXqA1PrNmnXHO+kskrzR9bFVs77koO1WLmN4XZ9tB
qwbqt98lJZhqgU0yq6tJy1gLcGFPwcOHrynbTf/poOnrw+2lFdij7IB1BhwTrwKT
4soZbHn9rX0ba9oH9qMCNbFivTCkv5xY0yfmVmG86d7dLOfFARqsY00p/BGLWlYx
W+bqJT3eyjY5DAr8j0EbfcMs4CcbzZZEygcUhvSGmsnTqADW7uFwT4cA3I8POeEq
dndANiEQtnn1do0euhYPQgV8semdyZWIy5pDsqCxEBbBBtNURrr01BJsdBYrlALb
x76u7Nqk3rVGLegK/LinRJP/35ISGJfteKre+iGjdU/1QktB0BrnfoKi88J9kZhe
wrNvhOMoF6uJfbtJKDi4Lg9WCF/lVg9j3OeKFQ2Hp7ZKQxjR5r30MzGP+29o9r27
J7TXDsm8bP7lvAVHZEJn6EBY0vo8K9c44G8gSAyQF9/JYrv/+E0IpTkrgmBr5Bva
sho4K7tPQFRUrfHE6x9ViYvEHWKp6w2NrMdPcmBxduTWRTn4FBALEyOdIfRe2Inw
ZMtajBB8VdwXbW4Dptdc2/qszLPBP3b/Q/8Se8JLc8Tv8CcykEpj8aaOHT/r5u0l
Jdh5ctivjySQNvtkig4Nk7o5qgerI/qtKHk7ndbI/wrySyopB3DEePKUklwcw9si
Ux8yOOBXthCirpFhQpFvMnhuQXD6X4EBrL6xxATFDitVwBmhjFLhUniORav4Uyr+
z33pMVyO2MFyQvkLQQQEET3M8Xd36Gxh64rMooV+4nUZGhEGBwxSykHli8Emfrxo
USD+uqk8AAUmBiUnYT2LsIupX40qtvVUhGO6yZp2vWQQkROGylkvO4ySdnztqtJ7
1liFT4oDQDa9/GjMxqx6kA847q+UCkqeEHMPKsMF3xjxRd3UORcW30iAyHYVAJ1z
y5oZT/wGgZxn7edwJUp3EccYEUowdBjico38mX7FW+IeosGKHYc1ipYBNzgWU+2E
M85RfhAVpMNK03ecgD7tCIt34kA0P8h2LDOiFKJL4GIgBdCvXjSDvZZ/kPArVvr1
2WDBuwnyl41fR83vL4s/JkASsjaMOscz9tFN1j6bJz/DBnCnRG4py3NnU4ynjIA2
L3Sp/4yFyQuSrBYphvwRFZXQd4+MgtfKMVjiw19La0zN6+a7v/zYvgM9nE488QTf
dbAiI07MTo1MptysJcM3B1u0RIgYg3mlTXOKwDa5awmdBGykCBMNYtasuGriFoSa
XOU7nYAESQl5lUAzDkVAPwogHsb6s/NZrBRpFCf/u1wG2o6KiWYolbIF6xlad6Z7
aR0XKRmmNtMZ+Pf7qE/UoJOZn2JbRqSnMIgfRH5DwK4UH4FUSZuYd4z46L7nILmu
tZTiGe/tKR2/iDTjsBvAki5k1p8Loc8iS9ND+W0A49KnawyJKyrXdlVYMYOp4Wkg
TqwqPGUCMntVy092kC/ieHzjWvY7HfTXn16my6EGRqN4nkfoxtYdZ4KQoMlGe1HF
r46da6TL8Pv69lSn/mW37Gt1qIOzW928x4V5mgEZS9zjNm0+mtRIxp53li74iqwe
1tmeazxirSoBRVi0PsxJR07QzNGtfoPntzkgpaKMuK3Gkj6kPjHcJ3Ct00jnqHv1
2CA41qi4rs+8Y3uzkB3ZgNEAnXyBX9rYM2PtgSZY9y6IE/2BTElmvv6X6khQziXv
JSUUt/LLKKrfq5Nw20NPlSVVGCiUst3R9DphouKKwhWzBElJKaPpMwiCLssYrOyq
qjm32PpQjkFW+1OjPYjsFRfUGbUswpqvMSQk6F4+DCCNQnHzaI1Vaj1bklSh1p/h
xPIZpDTEGY70HK/fTYNt/1CSLvLy7O1dHb1/6VFiZGxuuyI7fqr230ibg4YHwhWB
uQmty+UH5i3yVKMx/XejF4AFxSm+BqHeFmdMw6H1ytll3q0EcXShkiU+KdkYyUPL
knJWnJ7Q4K3EUYTB2qtA/fpqe5OHD34rY3tJQxzmYqhIQh9ooPZ+6ojWgl9YLzSj
sbWL20RHhFgYX2tVNdZJXGOBZ1fHjk5JYp+zEkpAKHPIrl85VspkbzF3F+Xjt4BA
pvbrg6xdFzlwLrrDw4L14fUQr/OE3mrmNuRnvKAjTNjQ8MS39rq8c+ia8HYe4DK+
Peezi8KB7cOdoYfbgqz+NYoFk7gUMaOeAo6+1y4DshPj97Gp7NscpOixCi2ZH7c5
LXrFMB4Ii7ybJsc1NaCJDfe0olCB+ZgAWL1+wqfQIai27EmP0wgHO1KWPBVHlGVf
mGceVfU3cBaNda56wvvSsyPe6tj/37oX/pfxLSx/9c/TGMaWD/1QMZXQBxGtEPDY
efSTQMtN36ieG/XHyX/sraVIzDPYPXytMtLJa8STbQUO2JnmzDLIHQw/D6BO3mH0
BdSjVduNG+x7ZWo+TDey0fpzRSTd/FKozvFL7YDprS+Y7OquzRAFKNIYDSLGF32W
E9py04+5Us68vq7xi9TnlCtMBRx3gDCbKSY7ADRdMZo+XVqB2mdrM1frKxKqMdYd
hzKPjWp3BwbTTxYNnR/R72aWyiBBVJjG8nKFS7p+HnYUVVgRfy8/jGubZNkuurHX
hunY66cBMMoJSdrfDSN3i4xzcImjq1QCmNxTMEeGK7EOpTCSjGG/DU605aL03ylj
c07/PSOlCrcTZAoMPWYLOxgZrl4VW3kCxP1AFZsB9AhTBDYmzJtyqVpysBFHuzo1
iCGyGYOIYJFGjlBY/rXGgo78pmu+PiuyXxd2MNK+f0hmecKCxld738GIZxbv9NqA
C5y47Eb8lzwrvbbCi7Q18BJedXDwUBXblKsLTxMTB6j9h8dD7RRpbqH6yc/uTrI5
Us+jO7AYbSbtYulZnExsqSk7xwwYlS/5rSjRmx/6bK6ZDuMZbvb7bwdbjHujCvWF
Q+0TaEw/MKb38AAImc86hPBwtWFw6RdHbNoSLp5hKg9kcX63/sJ0qUdEy3KzSegv
FhMK+ARXLG2uyRcI2KX4aRHRPQZvn0McDSjm384tyTd33gL5PlUbP7Yl34fUZFxM
EiJS7qsQW/P/BtXymOuwYDb8JdQs6+FCGJ8lK45hdO+Qy2sFHE3J/BbeWBaDfA5m
QYdY+YZZDHsWL91xq7LLzvV3GptcIO2ZfV8436X+414ZI+WfEsH3wmMyQ2yV+nyk
4zhJhLMrd6Bv8+dGbXR/6XS9miOz3Ac9OXtEbhpOPRdQGBgXTwuAWu+sCSPDNRFI
CA91mVx+YotXIQWUwAlpZgMdzu4AFHqx1AqYWKHUyCIAqcH47oKx30EWwxgBAfzp
vl7IwiFNZzA+eQZ2Fn0+ALYGFlvZJ4IqB6s/9KoEa7NBvh3gCeqjwzp7Ik1xVse4
H6R7hHY/syG9dEmTehKATQ1ZHdb3Jsre6EXYWPwRwf3cq4wPuQQdEF5ADYK9yxUW
QtDX1CI+q9gsOm7wO8yzQImSNvyN1eHZHPZtfJLJqocM/DFDvUUbQ5sNFabPc83u
1DHwAwKapebE77zRv5SIU/RLIFa+FCCvUfAnwMkGQfxie5s2gs8Rr832vC8ZLWiq
IYMs64BGtWzBbFDdTg+Gj8ThJTGf7dS/hDQhxaneHS0OUuSMSaJlVV7gpbwNSnQP
DGI8uNogifxDuYyyC7+Bbhhr6EAGOTE4Z+SjEKhK3bxSiXwXgzXCzYg6cH/heaWu
rnWhDsul5CimUDPIbjXkTmvBTEUwRvjgKlaNNbTcQ+DFN/QDsxgadbWLKTfSLpCv
r4XBI90ljUdvU2WqKCD1baWwfq6BOLAELcWCeNEz6eSPVkPAd5AZsyNNJqa5UHEa
3EvPv3awIETwCtfYBjH6R2t48ZySNO/myBDbGk9GZX/xcApq84teXgz+9+RssFMU
9WiFQmoR3r9MRNKTLyko/8gLS4qQ8ER37louyV0DP5XJjnsV4rObvzM9UUU6CjJK
QFc2TXGUQz3RiWgd0347BTv2Wl7DFf6f4186YZ3uudjrMpgZLSRNxcqqSHnT2U7m
7gkKTTVGEQ3NEjp1xL5mYjkwcisHJ7IFs+qbNhYPBXqRtKmiUP0IezCOkfGI7qbr
A1lfjN3AvBFuSnYWfbCF+cUh+m2fkMJwwzFO5GlfK27uKHEo1Hhtn2vW10DXoBJ+
EZ0TbVz/7Nrjk+L1Be5L9UezhxdBsLmyCNAc99IQOZIVhFKITXL9DXIwomFh9o26
pO2GyonR3t8JgpvXcXxrTOpbCe9GYpF25YoSBm6BofZrlQz+yEUb33MqMCGz84nu
APyeYsuQSdOTM/vy1o+HDfRiqwtyGL/r6Sg1UeVcgVOarWYJXBnnJQg2To0t1iyB
x9Rkc0GAPjufSwB7VGY0GtfIKxURwOiaMxvdEOlYpigr17bg6sEP5fSYYUnCUyjZ
vN1QpxEqmu27hRZ/l89CZ8S8gWo+mUXz4djtlihLeXti8QrL5HzhzV0HbXsapB0C
6wLnxuFRulgWeRjTDu7Scxu3/1zMABGZTa9lPLNWj+N1pT9+ip1CDvoIuNAtQDCD
ipLuAsj7c59Xk/rqZBqBaegr8ZM0DW3wt0toKTgQV5kES8maPOI74iG2AX8+qQv8
lYXYbx8Ejuxs31xG5P6I8O6hglsxv6n0XnraH4AcynGgwNgoYILEF8wyTUirVkPz
XNVAFHWAk9kOms5TJXJNtH2hhJFM/iXrm0zieFKywC9oZXSnk9FTp6onFoUKjyaA
bNL6YrbL/+x5y8EcwYAsmGn3nkdH3Jf7pwLSyD5dAQ7RNJPgYFbVn2j2RDxQJQkZ
OLYR9vq2KG+xBYHv3WnK2RLBNZj4SLWMFnnqaFeO1hIwyf1D9cHbtGnTT5RJPKmL
fC70JAkqQ9Uz90dI0LH28egIc8dwtMWEF8hVDDb1tD6bFV8D7eoldVbQdPA221cb
124ItosXh7h7R+oaYSX0OqIMBEGS7LcRzSHfZ7rYgujJ8cYWtIWyYJBPY9DKRD1l
eQJle6B4hMnaNv6Asn2lKot5QEWo+xgoIT9vR8yKKVXr2u0k4MhN84naMggT4K70
jRMrRh2UswM0h10lW/Yf8/tPSQNpqMYndQfzcU9FWE/DoMGMXyKINIHnwZr5sgQ+
OgGBLB44etyKZS58pwqMmu9YbmNzXyFA0uGnjLV0fHUSPsmkTfx5JiGByn8MvgN5
Nx4HxdVMAHuVeGqQ2Sdotj/CAI95JrSF71ifW07Z5tKNbIKzAK7C/kdvHmOUin7q
vDGgFbs54mm/4T/vMoqyVJl/8mbxyB8eKDd01pCGn+HmCL8GhVgh88E+8JEmkY3C
jW9pIVl7uKGolThTQbnbjou6h5T9pLcXrV2XDQXMLY80Wq4KaSn/7noIAZxtni8e
v7WDnMolE4XheJ0+ITjOBGaz+g1a4BXDugS9hyRSDBAZjEHk0qesQiVbi0yd04Pn
Hfyln6Sizd7g/BBk9KmKJiNZ49brdIlZO4xFPUasKr5hI4oe1u7VknMBJRCQCKom
NvTVdCvNvfX+0w3umz/3FHOJGAJze2u2kFMq5rSUHUxKCJoXxYzfYQOoXHa9KmhT
byhtasSyBsAnp5moERC2M3a7AvXHp2A7k9tZnMPTXdaj6Rskm0HdcvIJ2FJPcEyS
qtXZGNL9r7nz0GPEgiavKExFNpJtx+t6HdY1iPwIXk8+7odKNQEA/nMkiQjMhNTM
k56OrtwCQLry4n2R8/plbrBaPo60s/OsuGUfXUYz0bMLDgCmOgu/44eVw74i9U5+
VG+L+zyEK1AxbSbWAFHfUvef3ew/OUpqj3Gb0un4Dc7ba/MmMbb+9TAc5y4Zt+rX
1xxQmi4To6fnbQk0of4s3IM3sErCAEUy/DmNdHWwos31b2hzEPuSZF8bIn6mLcF3
m6E+I3wBhXEmaMZbduTulkJHm+RMqTMAtaPdKGft8FVwAv5OkiFIaE848TnAriXt
nkecUI3jjHvAUJhgehQwZTd6XeAXHlG6Cs14/AlPduYOrxNL71RvsHizwEJGvgPv
KPBoysVp8eh818/EuDDa2eOs8AL91DsHlZxP6iLWsx/uCKdaWsJeuU70E7xNF3Ub
QxiRQ+bhrwtCzoYra68a4f1hjEdGfwFLmiY1XxtoattZI+RkHR4idLDnkYglGwFU
LavW7y/4vGDEampl9Id9xHymWM8hQLkE/H2SYeAWWp29mjat0+8dhTDd4MKTqxTt
bK+P+GzR/h5Y8s6TDl6Q4993ntHcI7ND6Juk7C3oQ25QBZVxY0ln8TUmWV+bQePM
+x0v26fgGgtMDCOgRe4vChBKoApgv7wWWsePqIAdAJVEPTYtYW06X2t07PcZICgM
wW4AIv8ij4vP0nETp+zVjYr9rglXcan4e0WLg3oGFM34dAM3EE2tAcfuDMe08KaU
/B2XBcIJxr/mvYWZivUwvdL9N4p+G47bomtYkR0EYlUnGeXmSXJ96usFHU1NYaEy
f7QL9JAbQMlqEolYv5GHt4K4j/gP5q07h9UXH3+wDaUoEfcHAqaniZ9ifoHd7PP/
WeFay8pNRA9g1eAIB1tGeztrkqGguYvzD5AS0yj3iN0JrJbsj2cIv3+h4vOziQRs
5F96hpHFJyCaV42xiKO08PSlx7yiHemzFv7iD0PlhOw/Y6sqjKAMRtNwLOaFc3wT
yYH8uUMq+74uW5MJBPCyXwnvl4982X9zIIgi9x12JVxRxCm5LMxgFUFmt3FZX7YL
0NBO0UySnVASHFPYEZBmjVCNPfA348MX0GZWQJZbfLp03LdTuv8tSpO4rPA6KqyV
kIEOvnWiTFN/bmodR9vS4rnxXz54iUcfd4JQLDiTo94q/RX62WXzrNf6fwLF5ozI
bsCCzfuBerFGI1uIwDkRiumNBAjvnVpfkG843PGgwnnl52v752rAoBJiN6+pNGQS
NlUInOJ26kf3Jk36mzvz8f6oVq1eIT/VI7a4lodxcOPCBvUZXr5HIn7vW2BLxt3n
Wvxmtcwmvhfm8WLK6gAjouSf2iSr2F1EQSNBTxQWleRFST3LwYKZ992FT92QUdrp
5uyROXamSq40uMIts7NEoAb4x98vHVQyf35VV8pXNz7IzCPKVmkD5+OXbr5QmS4u
Q5hrGLLC6CJsLuns4aWQHwxrwgoYlz6H7wHvYL/q1uK6ZS/DLFH9wTyImdRn/JXU
0JLK0oaalUn8tZU/xdkDg1hWJU2+pk9uRMiRWhi9XQroMibWAhC9HPpPN7I5eA/x
AMmFIJFjFJG3rYOL+PnYuh2BD3jvdgx57c93HtaGU0skIodesUmwoF5V0rNvQTcj
nBHpn12EtBEtQY2t7EJaQfSIBG2SLEp4Nf3UJXXiDD4lq81fuwKA5yccg06up/rW
HU8OFUslbt3CHLmquGTz4Dqb9v7TDpWUImhd1F10VGUI8EeQD6mr8l0VWm6iQqIP
p989wqWGNIR+dBqJi/7Q38jIpOY5NNXEvRSPz77IFazc9J7GdIsSP/oVtS/sqpp+
zT+rjPGGWDtWuuPMXLY91XU9eNfrqFnmQWXQu31YHXnGsn06Y0lDNRrJOqeHOTlJ
a3cykY1aYyXZ/GTc7NxIM+KEjRN/e4X3ugkDm6ER4FjcK27t0no3IjoWtXkmNyp0
YkkTviqRL875mGSDqVasD7bZ8T4pHf3Wr2s4bi5deXVGwhyA44OB5o2KBm5N7Qli
Zn7YMQMyG8qhrR8Bq7leiTYbLF0UIagJ/SClK2F4zzCitXKVYAOa0PBiahR6Q0Rd
6Q1yI/d/h/aeL+BKduO8/uxgfqyBLzahZTFiOCt1qhuBpZtLl/zPyOLuDrozm2/y
CqZPMHw4pyaHLIgIaT53SNvPEjeVcbreM7bMPjQiHXTxZIaNY5xIooODya8GHJ2s
wuyoAjBF4dVP1EtAf7iCk294zeyweqs8HY7UmrZxd7jWRtzz3ByAILT/wwwZ1Tvb
JUXaKyqn2sulbZtiVHGTiMnGI1mdgNYlzm4K/JUoS5wDLapIGCxB8YriLYf15/Ui
JnRHhde3UrA5rPsghoLdxaKUd6DB+vS8sXPWjoLeSBiU/Zy6TYbzegkEb3SDAA8l
brquSop+reRDWU+B4ujuU4CIxrWYcOwEvYKAd96O9URd0lmbdPPPaYuJyFpKgr9l
A1DCFAGcgW0gd9ER5d+xST6dhYNgH25GdL8UyxdnJSIqM2cR93yNY+Clx09tQVb+
fUPhN5JQQQ/aWHAl+tlF9gn4n2l2KGl10Cft7uqnhhJ6WnjT6xgS50A6Lr4164Gk
dx+CvNb4Zx2Vpm6swOmjrlHCTi2WsO032gLEx2QFXwgNwm8RJ8ErxMmlzzBqbI4/
0CcYJeWHuBu7xFJuULTaU+Mnk5gLN4GdeWmGgkHoa6rOeNrX+O100zF5JCQftm6j
qn4CgDJ2FTeth3ATxeiBsrp9UBghzJnpUEr07I8cDiEKbBybjt1C8/5RNMdoYZ+H
l2Om/K4z07yiVWeSIYsrr5v5vvR7aLq/VIRhhN94dl1fPMl4TXyC8eMMbQ4Pouzd
VLGcZA9VOLlxbM5utS53Fo5lD2PxnSL0Fai//xF3YmSVSwNcf51B5Qj/Eir9D+ke
UPpfCtsqHq2811KcNdBHtjst/HoG3v23zklKRP1Np7q7XnML5Kigjk+AD7AW++q5
P3B2YOuorxwD+eabye9SySkQBb23EcvC4XFpYhxZxutmpt8ncSmSHfZXVdgLHjHd
/mnai1x8XourfIPeT/F5N1KvR2X7saNk+a3W6EDNCF+eKWsRcPuFsqk/bQGCd3As
XVqxiNDaqCnAYVpdYhbTUFIsC9ynU4OKzahOabOlLgtvLHW5OCyBWJhg4nehetg2
JoGqO3w9NZsCFI5sI4g+c5ToMoYZdnVTf4GaZf/079PFuqUiYoCHsqhGcjb2GcNJ
OLbmABCYWFl4SbafXYA8QpOjoY3W9YsSaCqwZPX7O+40LQapjT9D7bt1SP/WfWR7
fLf0OuoJ8idXyEZSLlGiTXnjNZ528zregk3Cip6SimXUrDVUuwrb4Ojl8l5kcB7y
D/zjwpdTJAKnwnVxYuVDuDlwAgyp9LUsA0k9EG38YZq6YRA0BEudS7xId+GBbA+S
lCIf2FSLli6gqgB6N8Nu1iJMqjZg0EJmyt1kj73aKl2tU+jU/VIy8L+1YJZln8kg
ypBYWZrImQQcgDjz6yx4OdIeFmJYPKPh2vdLe2ux7s35pOhfliZOiFRkWuFbJnaQ
LgjanQj+9cKIeTqrzUTdGzsVVk/Yi3KTWrg/vwIubkgi2WG9D6Vjly3gvbcrrFlk
d5evhvTmZ/eiL46yPe1+nU2yICDS9vpDQnYui4xh35LI+wBkDZZoo3p/ezfdCdP9
pRyi+tBIUJ5axX2YVjnAf6wYcZeKHineZgbXEEpEJL+AkwzVgo+ElRJyvWe3V5xY
uhvgm4MA+JsPhlLo/bvdRw5WyHJ2GBjIKu6tggA9WzuR5oNmZmrV08+BTrdtz6Nl
5qWKTswWNUVB9qigSLCyL2m4KBA9vFLq/lLmpS5eBiMgiAk6WecV0RhPUlRc4TtW
GbiBIkTK17HfJIkYrEuReQ16p6t2/EJREe/pMiJEvPIxb18CUi1rtlx7h9Ci8wW7
C+ZcWp6aTNtp6QAitQiW1h+cooQm6MG6bPHfyy6XHjBDQvfXLAcCV5wYDEuF4Qko
mM/5wkoVdxt+mLN5W/nrhGeqSAPPkMzU0lMnWp1sNCm6KI+fK6DjlIJu1InkhC4q
sNcutNSt8lt963U092rDK48+3N4r8+f1zOCSBz6kDfX3H4WVtayH1pbgeir5mYtc
gQdsrO69s22dMDlydDlIlolM5zQO7tVN3EPGdhsQ3zzZmwKQaBFg9FbPVz1c2E+X
wHSsKL4W9uda8GtWurEXRDDCU/I6v39FToF9uVMucIP0RmDYV0bSK8fo24YzKbwV
vlvFl0cCZDY4WnRILN/ILn7ZyIEZTKWD2FcumwzqcFq7bnRWz8CYK3Vgt2TwZZ1D
MqRJGvDTSFatHfLiBnzgLsj3hX3PkGyn89p4auMbnG3siyvRrppi6DdN9+cdiVxw
txMrYDmEUqxvdhQXeADwA5oNPamHy7YCrCCvft0zsHyYSLqUeB4Wca/v36pyBSPy
ug17CvrY581zfZgOQx9FNe456OO6loUmNgZ0TCV2g4bDjA+BQv55MfvLhGjEq7oR
75pkHWpvfYhTZ+CagNjeFCyioysuBGr5AUd8mtxWE+BTWafix9keNUpsBklJS/xR
jdYXA02Gh2yhmE6ZeZk+g5OwHdbrpViD/4mfqum/wTWj5XedOuKIF+wGf+A3Jpo7
LGCUISpSODSM7oWiW7CSWB/fm5Bq07nbYlKibTr55NSQKX2/DGrsS124TWjtjtHx
6+6WJ1Nnf40VFpTF+yBcxHDb4fIunf8bde7WLbjmHVwpEhcigXiGLMAAheYTWzcY
KcP2VKVN2qhZor4b8XwGjoHhDD6JXnAdhBJj5ZoSnxirPlE2tXi9haVp9s2Wyqx2
NMtjkT0UGcYk08/8U7mJeo3CoLYf1LM1x9Zepqn1nLFq9qQVA2KvbSaUoRaDmddK
q/PrFSxt1jlqvL+kPVj0+g00vhF66nb4bNG0iLwDAMyDlZAVllYuREsca6GSqgDZ
5Fg77aFBFmDK/ugWd0s+TzmhaupUxeLEIXzlcAQd5HAO6aqq6OX6fKkDgGcvR9/S
jWDLgYoG5fhcoav7rHZBFw0dqBcuT4BERNTFBGjMU8wt3K4HttwMgg/wMJrebHaR
Q9pIfuNjIAwHXnUikISegxGI2YKAhC92qmCdJj7/HvNB5imW628K0lHVRkUvOV9+
7q4CgvvStP44+W9ZWsnTB4SoE377hbSlV/+bF+7I3k1F9TJwfXn8DDbJcmUUC6jy
LeB5LkmX7bsoAoiWOSXLuINupvt6CTLbqfhdrEdgINGZN8fzuwccPLh+kqUowQ1G
WlFkii6BmbjqmLBnUQwhigJhtyGp8CK1GIw53ah6Nv11wLASEw8mJZv1WgDBMaOO
RlV8wLnQ9seozuPSBgSqeU2HdoRcDVNLTFGumRR5epP9NX0A7+1gjHvwJjpSl089
8H6L5DZ7fk1R98R/TasF+Q/J/FyPNrdd78nDNYY1XXHR3m4V64d5c3Ox6onKz0hn
TdS8kofxTXZxlfD7/pvpXnykC0Hfeko3WIkQkQTSiA3LSeh/+tXxdlvvlqJXNWkb
ojzrptkDoiU1eYYE8qVeHCIi8LABcth/sb2FGkn5ufhhrvaL+UHS4zc8u9GviWYp
NLz9CkIJCosAGLsYB9e9NZNinj8HgZPXdv8+Is+2uHb/44/t4uLcE0rZnt4VwtwU
9Beb4PyqXaDNrJrKEpgXCRDVHaihyozueT8ikQotNdkfthCdUnxC/tTXth2E0ejs
DKorpuz1HPwHZZNIePUc49GJksXAmCPGrI+4uXgGcugJMa1iIz4aymrGPrRi+63g
93gO1Nr46sy6zMTSeQ+UFB5QtflEuUgR7fFp2csOTeZPIJ9lD4eiwfE2qkqUq9UM
0gIcpf5AF6RvcPl+AuWDCOnbA+/qbQU5Mtt26zXjRM5ZbV458rGy6pB/OUQvyAwc
emiVFNZQdS7OiTBZKW3AN6cF6GevVyDd5UltMkxHPJwtxOJfrqm8ZXTaNErSp4kC
+ybcxa92ZgldzOgYxZ/wUzemQ6YXTmnA8E+5+ygJ+cmLeqSOkkK3N/QuwFaeTQW4
Made5BecDuyaY3zwfOTKqzsNoq5ctOBLswYxzREbmyAwRqv9jEAvsezOv+h13zR8
vncHKa6sM79MU1mfHPchh2tl4MQXa8nrzxhjmIh/JZuayLGx9tiLsUHkMMjNITt4
y0oX+ndbKHo2FEOVpVlU7G+7DYPpdEHhb+LwO4YQAGcR9rFcD9EBoBi1vHIpWKpT
vNBcrYFEQ8RLMrraYk4uvpfYcAxmEQhQ6YbcQ4L1IebNYdxjLvUrHIoYrgFz7HXX
rVFtGgbOZ1q3Q4SImIFjZP7IFLqeAmaKzD5PR5OhEHEdcPpfirUgvUuTO6PPuV7u
T0fA7Vu4zhIMuo98og7QiOsruZo7HJ0ZAO0ZIWz9Im9LMLSk+m+DPrfmue93Kjbz
OIRs0t5FK40ouAg1mx3lYL/LR2Eu8PpOog9zJvl9QyqWC8wlNj/pf8Zran3VTV4q
ACOqMxx2Rhj5cZ8bLn8C6pFXPkvNvWqd0WPrqfua6lmc+LY0XadNanSsZRG5oYl/
AOMzdIDxY4b2CQ03vDW/8JwWQFY9SiJ4zGfYQAzGv13IRvhBljcnlgLih3hgGToi
iR0tk1ZCAUpT9+25MCPVYltD5m2+5xRDT2MapnJsI3Vq609IIe1+X3Av6rOK2/m2
pW387brjLQTddvZh1PKF3enTLQ2j74zsbzFbyXS92txNdPnJGX5HgOFCdxnjQdvG
xGcj6uTcWAMMpV3/Lp+oj9s3gtlJp1vRJBncmEH4JU1kQrWpRwMEaTXZepR+Xg/X
ojm4QuFZyr/z8GXTAUYSJc5Isd1SPhkMSQHaoXuQtabHcIxCp05rNebuhfsM8I6T
H23URhS6sTLkYYmPsIuq2pIevNPHcdpXadiOlS0i1HAeVMGfdlk6H6QWF1yG7OUb
f1/brnO6KgFGHNBKGU/CMDFZV7hrXHyzpVpjTq4UlmDcGHR+kut+d0p4ByG1IUUK
cwfzpCOakKrySRvB/WvhPn3Bkx3Nt7saoGm8pjkiImSJo+2feJZRNBa5NbL6hpcX
YfWDUgMshm5ixXsKRIN8ZDKVtujKVDGB2y0SZQcbhMgvJH45i18KLOBW72jYVeAs
df7nYtVodH+cZPeLtdRzbHBeB0dFqW9aHRlGmyfn0i3WrzGvPbGEADuQ+K5El6k+
JV16JhiQYVDsbuXr8GW69SmIWijyCDxFV3JxpNfV52mZd535bF63j0C5Ov/mLgAX
SvLoLL7lr8PtnqwDsig+xJwxeF2xwj4d8IT2SNhOKFVvLMBlEW1fc8uzVQS3dBWr
D6hKB103ZjZUjepE2X6NKdklN6eoQtyFWyQvHYs3D3Ih2cNY3a9upioLWetu3R0R
/4DEEjUkabGa1EUc5uRB3kNhCpsckSAbn6K9bmOKlWbW5e3DbBLiU2hpDSPi8d8o
/AGGYxbjf2FEio3G7lcXwjxQllZrS4mRUW2kn0BEiBFU3Q8YBnGf6Ee1YViS3Vlb
D1wEuPMmIJCX5zC6hJOJuJNMOsL5uaq/LX8P1GiS7VyaL+2yy7rCyALBqTcRWiqg
8LH01qxQcy6aiutViWnmkaaMu0OO2sE3u82IPvmJPH+Cb7eIOr5N40l4KcR511Zo
Or8dLaD8S5v/0T5OhuEItddz8psoxQORO98W1iX7T40bbfj6YfOkPOvlhaHKaODa
nk86Fci95jpAZm8+jDIuuGDDR5GsPIetQj5GSvTI2vcMTZM9ZmJK/TGoGIO4HmAz
BYzVGTPDG/0mJ7ZUrjRi6BvOeM3Xmkji/EOxF4Dy/QHLdPv9O9Lw9ycRogc429FM
LkO+RDi876iceeX8vAf1snhOvinHwDrb+zmXxhU9q0Kiw5ukQqZkLcBxbHEILdT9
QtjjwRRjkEtzjAzpHtsoUBhgzW9rueiBLIyqKzXuV8DpTZsZcHYR2X8n1Z5flVAa
SU6zsAbzrIBwgvLTSFflCZJyJ+itPCd9CK66Uqm/KA7Sj2CdgOm06+1dvarkaJM6
r8vRk5Y1CRm1BLubIdqo9PlfSUOxFTpa5/f4V3SzKCaVFAb7ZBRpYvW48SKdVPvj
0lLTolHp1oBa71XyUIjvfb6hnIZdxQyPuPsHVgYp8E5U8Zkbu30xxnvGe2V7z81D
LbZV4+LQMByBHa9YR6mDEOVPvO7+bP4UyPwGmlKpK0kQCFwqCx2L4cxHP0jnn0lS
pTmxondzHDJNVVPLP3X+5511sz2LmBo4OssK9Iz27VHIr9cM671MhANLzMTc6ExT
SGvid+AOJIaVlcT1zwUiV0ef6f/nvXDJiu5IOWidwF7utDKSH1UGo68TzMnv+Klt
Ac4MoRSKWxLwwH9sszgyA0AL1f/eF4PDkd63IUJJ0Z3R6Ih20mowQ+jxtaHqNsQD
5XuqEjrdP49/0T6k86etiX/JrnVhAYHMh3jzIBQCkgmCXvb01sQI1zNO200tjAqh
iING9DquSCv1MLHqzc0eXhdLhB9pEV7O+Vph1C+sN5T29tNdLvDOi/n3G4QczRDL
h8dAgZkKdR5gXLaEbYRdB5WipGXvZl2rXHuShBbMjjdnExQlgN8xoexQB5tK3mtQ
NEWzPBACeA6eArTlHZstsjCGhu0JwMREMon+T0MHZ3T/FIzH0ZZlNrdlGm1P8uLh
PVK3FCPbXfemByTggsQq0IFNPhaXIFdjMtkDrGYVKBRKo4q7wPEsv9+3QyE5N9y5
wzy5sg1ATZ5/0ygHjqlqBGxe1psc+QrA2/DOmt2LAQK1ynOlBSUpLFprMDC8F4ra
DGkO+wqm4oam4cCHl+gg1h/hDFFdsPwINWlk8JQNsTPp7J2jwD6n5hCj/8xuFcul
Dp7i2jLycRpnXanX5tam8pjUoCKdADGqalakxM54mshIg9RMfOoAlavIJtvv0hZy
dfluuVHUa30pmposEzdNfb14e/aARSG/qFaNF1En84Cqaek+MYhJzuO83uKrfFNn
52pDm7xESHgiCKfu4FJvgmX9VfHSZ0NrQsVJEFNm+pGWw2oVKXIKDibm69vzHLLr
HqxCdQJ+ZmrFOxb1sMKoRRBZnZvOT/ACqbbBhUEn6nM8R+Eg0i/DKYjOkjJgvlus
Bffysjj4Mi7UuC5icEGFQL34hvX21Lq70G6Dreadh6syYRCKht6+YAY/mzyV5hFV
Ym7sMx2bKNdEjyB+9nLda8g9DqyvSjj6Nld+nam9PwviatcrEpzEATMIDThGL2G2
4KLFQnmBZ6CE7lTHIscY9ZDYPV5Z+WY+IxtujO8jyHcKw4+xw8xnQIiKRuMhW8/A
6v/52iSU2ATXi97eUK0/Tgeput2sjH4Si24UwHfBnKc0DCCCQEYyi1s2UQe6WCG2
SwphbED6cjRfMp+nIabJcRw7dZ4JphHVN1uaCbIDl9Bci+tFreh4LDBl8CbgLfi9
eaWfy7+N0ndWZyd7GHv19ACs+gzo5JC1Kh9VDlKInsKVJEakMUPHRsczGyWp0BMa
KmIhaOiQAGLA28MA0rJddY12gB8brJF7iCpv71Yah/eQvstxGQ+gueT+XFB0DMhh
xp4OQF2X5Tz7KbtLNFx0FJnNWqggMgu61Bgi4Nr6RNLmEwR/S6DiRpVa6Rc5qMjS
5t8kp3nRJcbBxZPyQQUsISxdm3AHRuVdM6bxCRABGNsXKmPHUDIuN9nNEYVEW6ud
v3kjEmQTBDAS7e2/c/tnl5KgSlSTYX67J5op75o+0PyK5eJ5zmWuhOno1vEbBqtg
F4stD4H1+Ml7XDyak860GhYjp3VaYCx1EAyWIYmIRafZvrsVZ12Iqa3G9YGRjheY
bwmwDdVbmYvKCuCuFDdhB+OxW1qaa7LrLvXItPtr2LhZkSZIaGQzcUBJm3hrtqJf
7J+uNQgwAN5UJA0enXlDZe3e9T82khpa2KVNcoZZNqF8PEHcmbIGi+WfPOaRDNiA
KWY6WwA3N0IpMtq0fROxFG+wEa+dHP9C4MSRdk8VHzxov4b3scle91eK4HhKaKRV
gY7cohwHWSTYPwzoK2/kLQ1/E7qa+XpAV6eAZAe8fVjT3beiacaYrvpEscFGCbDN
oyIb3pVNg+D2ckKPnOCwUnFkOwxPFx6FqHttaXYMmajsezbGtoy3lSueHu0sHn4g
vqGi50cJ5FNiZV2WG+t9gjWuzB8zHNT8tStWJG4tqGpZgzbjeU7CkFkQoi2Pbp7M
sAWa541+ng4P9s4grcjIU6aUJ7xEyhq0fFx/U5U2Z1RkSEAb5UPSrBHEbpw/J47P
DgOG545Be5IjtX9nGIYt2/a9gOuTYezCvtNOwbuJ2qE4A5dUVuf5PPlEZym9SS75
+JMtTSy6Y66DwRf/yk8T6xhjoVKgJAvRUIvjqX8m/+v6EWUhPXkwQaojwYW3PVuV
KAnOVNElHOVmdYfJmnWTixVEFDMfSpJsbhxpL1zcae9M4xqtYqpH0grxtvGWB3V+
1GEpL8XzNGGzDZ16bNyFN5XO9jXVGeQ9mcY4quWnad3SSw/BXw0n4nhu75kOeSNw
8fQFmh2/JtDIMI771YX1T3YKgTun6BtdvsZelgWY5nTrE855s4ZFXCo+ccvvCP4P
H5/GbONsL5VTcXsQCVJy0VksOMLpleDXExpW/XVjN/nqjBg+C+H969LvxemM9PIX
SnsrDSzm8b+OlJMQYHFB5tGnDHjfKJsVuykQS826YQSrXSP2Y7YSEOJDflP25fKp
kgN3f4RkPD+bbvs2KMbxojE2jvuVuZYZop6m0XBCovjZMzrTud/L/mZjG7OcZGD+
sOQG0bdCiymC1jGcKZYpLW4a+wJTWMzMj/g1+ng7trn/pAYx1/5cuFYG4XrjVbtG
P8sNaH8wBj8n+cnb0iX0kti/6uPu741dRSWtV+fTVJmbbidKaovQUxxFwEbFA2iZ
rboVbvabvjfRTg+Hmgi6t48T+FwLp55OIugXo0lk3722Ogy7AQyAupom/Y/Sq9Sj
1AUvScXtTvVsk1TulmXYfXeuxo6dgRx+/lPxQ/PPD+WTBbyDmB3MN7RmyLS8CGqL
0RdqNxBxiwDelTn/wJuDy4ACN8zOH3dzTjYyl588+Gy57ymsQGYFvLTPfdU9sUiX
KHMsRpIrzyxr0x8/bQgp8zZfDJM0JqmBc9bbjqkq8c67tNpaI7z+2IVLQ8lV5b9P
4EKoetvCD5GJDgCBS1/cQxolih+Gj43whzms0G9Afl8WRSK++SpOCdp+YCjNCu9+
EvN9ZS7X32oVc4nP4katALG6kiEEDxQtQfZrr3ecd4/ZnzELuYLpam4Cbi2dS51U
jCNkKZwUa7te+w3ED2Ct4BKliLiprbvlq1ozPsg66809FuNVUOBrIe8i4srlItLw
av7nA2ac/kYSXGJklbJYOxpgl9UoODKx0NkZAm2/qNmiG/oR7m5yFqy1B9jz29K5
lUIBnFzgnYJrW60PdTD3LBruUa68i5dqUJGIGF1SOP2hiCej2HW5EhkWVnXnkKnm
4cWXCqbNBNeTto0mkjYcq0TZTIL1Doi/HKtxLw4BgfjiMJsgodEL9oXJStBH4dpX
swClySIcK01J83J7PIvHpP47b77Z9/O0HLKp5H5N00NZosP46b2Kmyf5/LlGIP0s
7s8WzpY/kBfUv14xmUOgcgIzUhCIkmuYSu4mfFhpUnCotCjNMUozRT5uGIVQ11xI
qK0TvLFCZGDiI0cmH6f+qbuLK1g39T4JpzVH3+GrJiattusAJb4gUkNb3U/4/cgX
r8QkGzIQPwktpEH/qavMOeGNQwz4To1lg46tLP09qmv3Yx1myZxCvYQTnjU12gnd
tcv8/zfZ7TOHYF78kM3tzoMyZ7ZJBcLCV5f2vpgw75QT+Zm6ZW7f45v9e0nawfHV
BUU99iV3uIzO042Vu3GvbcO7TpweAVOWWElVlFh3mahj02UsVvbxzd3tz+223v3O
dw4ViF/Pf3GnDvU/TKd+ItOtCbV0kcYF/lO7Ky3KDGCUZ/ykGDivCvxFcmrCiGom
3BlGIwnWmzwmAn67nYMpZKJUsWdt/5ShKv/EZwbIVPfoNGyng3Vx0ZXAUCby/TEO
EHyqAcxr9sd+RfkhQxL91JjIv6o3W2b8bPeWZX4b/s1etW5lWWAPGt4dd+p51V+n
SgcwZmphLrRALvWC24dlB+m4JoYEBkoOQNYGjEMxSjwL7GOiU8dc4tXim42rzwoY
rYpwQTo97QWSzMVe+dkcsfO+XU8UgAYU/CNjddsXoDs7skl3g5nxtjzYyjcw/x9j
ESZGmZtMmiLv0H06Ie9qHELZj3GWXv+ZQXWwG8Pd+Q/CCesvGwbTPc35X/CZcEjr
dTzdCtFOrfEbQjBgsVOZiJB+ymYAqPp8VHH11Rgc41mRTsmNJtxDCoJ1jbr0LcOu
7G1damLK4pFoGchbs32oQXQYkqSFZ3oySlV1iJlw10FI+IU3znjsKT7Hd6hGvvvK
vgKiHirgZonMNA1iHsJ55xJzZWWXf8eWwm2rxpNITPn0QHzYTzTurHhmf2yPsHt/
BbIGvc7ECRd0bBwFqoQB7fNIWmaQfqdP0WUMgr+u/vQXKxadf7BwjdrmisYFaeRR
XaJvfrTS0YGXCU0Q7O7RD9tnqw9t57X+kBsy4tUx5aFB2dQCcjoSsle7OxDVhfDM
8GFszU3xDWpyaOkjY2/mtOAv/zBgP9gnlsax7mHLAOdfmcfQ4tdlN7x8UoS3J276
NW5xuxfjpYcAm2AjkVHplWh8Wy6phQpQCRAoB2qGuxxGiIX2qlmcV1qITDUx1Ico
koS4ZT9/N4FwmH5of0GZHOchLLZwwcNa9SOMumdkXjh0iVZfxtRHThjSLUsbzpTS
VEsa8N/meucr/YXxoKm8JP+kuQGbApkFTda8GGGuj/XjmGVY/+CouWZRoh6rdJ0J
LF6mgPOmC8N0M7wMEDCKt8S1omN+D+1K3LBf8931w2xa04quiHUq7ZPuP5bkjeq3
Dsfige47Q2tPdYLjakIs4DhVNoVYKKTv94opdEBnYbmsdWteyHSyz+0xMqaqYS8j
reYaerMbiQ2FPqeQhp2QWHH3G1o5qTjfinYHHqsIytUUJYTWBgtLAH4xSyXI+rXE
kmJF7SRceyCPHgBRlbb/hGWPPOY5MGy1BpwnO3EwRC64UiOOOx450yXBSn5cxRRb
PYWSALpwBnTly7YjX1918eGNYBKrzeHcObRte8I/1FB6HVwwiPerKuTvQIWD4EvY
J01haND1l4FiSrCsw/6/yY9+OzaTfjI8Ko/G4rKjVm5Qc78hfErlRn4lX/HQfNct
MccIy9slHi2MtmDyYgzXCcNABZnxiF6+OhCaJHnC1ZTO+rbP63eZdtgutCkVhi3d
8GhtNgSZJyEuGEIoWKq65fPFjRzYUFAAVxknwu5NtAoKhCR0dckFKP1hCtSYrNLx
cSiCB6zOCn5bctt6hvtdZMCGxnmd/Bp0DXYy0+X8MOPfUIQw6+JqEHib0lRx4jBn
XBIJXby0oLQ+ljZA/GS2c7hvWP1Jjb5iYfHNkVxwaEQ0gxmlDd/niKL0bDk+LYV+
rBcn8YnqJ1SuMlqSJ8q/IN/u33J9Oux1LHuPzeeYMHG49a4Snt0/7vVo+3UsDScG
g+cUvFQqU1yVEpEayPDMNPtYB5vKFoVZRF6mpX/ggaYz9LN3okO2iFxqRL4I3CNo
WsWNiWNKHWqiuMjymCWz7W1WiM9lVs4iNLQ2VtDa8OflGGKgPokskXvuWElWhvMp
kRFtTBZoJircUcLVjzhwBR6fIcsTThNwRQ6nUJ7UATDiQYskrXPlkqOR7NyfqQUk
SLF8rAlEBxX0Te0nzEdyHR0KVc4hOiub8nYtzjr5XNkWzLGAX9kYE7DAmQQQ3BsF
zk798aGoytEzh0fWpfn9+j9/2wddlieP1E+gfLmtHRBlxRXaYJaSVJf507uxaJW7
61daoCVrQPFr2sSiiZe/NLWDbHu3833SzwA24HZpz15/thXcSqfVaP/SZmW46YUi
VjlriBQwdywUYgL49MNhAl4RCcI3gGI+IUdobqmDlKk5kOMDWkhuW0IxB9l6KrRe
gTu3XdZyQPGllEA6zOyyfUc4vmvXQIouXyRfXk4UY+MrfUVYVxcv7z1q1fZPixF5
AbQNun58GfC1RxBKoK6dsiWJHad6lkZ/jE26anlJyBVNd3nVyn1Xz0H1z7t/cpQg
ybhchpC2mibCyj41sCf12fPQ7ckPoTxJQRAMQXzLpxxdJWvsLLQVhCjEdXDDs+Ld
dTDPYVsC2tMoBUsB4SqLdRGSivu0TxZ1xtJdCBmbkSfVhR253P7sgyZrBSuQXnE3
ZMxtJNzFgHJ3awE9GOfK44YC3bEhJ/R97Qq9rxswlW2ERsaPsRrGdoN57gk5zSzR
BAX7LG7xogSReTxMkvMCFCPqzIFiA9+khykpiKPyDwVTsc3F3vpUJYjNvCWv28TK
sn14mNSUjJjs9a3uflsp9gnuKNsiZ401mvjC59SobK43U+/iwNGHh1z3sANs7eql
ZR3kmIgNkxqULk1Sn3Ly5cTK/ZiX1/rFfPepK7SNv9iIjmWj1Zhc1lTPTCVLNczk
ePjQXV2W50Q6KOKrMeIFxcJK+NCORBCl8Suwv9tr+VOxENI1RXFlN3/b6He5rQ5l
g5E5EDZG37sZzL4rrVseOEbtXlWJ2+/DFu/StJp5/Dx6ZXLvmzC5GFqXQpML/zUh
mnnsAKEC0Iy99uiuHtWt0Fqe59ZUmgq98IC1kmEtJ69O0e3m+XYF3KBsGbaIfn7w
morvCY2RI9qXO+m9suwZEwTW6eOz0HbQQ5zowxh95CYHSPQ9ySK0CjVQojaoty3E
SFLPJkhIP0+3GNo5CNIu2e7bSu452413WLQOenfVYpD74eBIipTpvdWHwhE6lSmk
5ZuRBsZs3VkXtxcGRDNAg10Ngtjt2AUfQSFusaTdkm22Uv9FZPQQm/jI+4IFLu6T
XKE08cf/XMoHkU0RbopKiZLtb94QdL28/D2rwtibxQaINVqLr0MN3qiTRAP+s9U0
TdNIMVNArOzUaOoxpoALj2bG9BuE4B1C1XPKtT22JMx/Je8DX1NQPXogvJ2dTbf9
GJKFOJ4jdB8cE/oeQjObFmtPW+Bd/+7eIW5NSagMIlNsvM6PF7rhrOhje6gFMDqA
by6R3M3GZzLeuo3bVrnV2472pSo2ld59Oug2E3xYp/wn/YeA3ucmyqfuFfHANSq7
vNh+oopDrQw+xGh78sfrMBbWGwLWY0n5IS8m4CxZEDSXkgJA9cLEthzi+DIpeQ++
JgsU99+UKETnELYGhOyJtxlv6KBitLJIm6zSNRhcKuwzDt51+lugRliSTBxkaXxb
BsihA0JtJTpX29pdROJLQqhJ5fx1sejqtAj74gDpsxl4MxH6mQlE9WscVnlyqBPs
g6Ys/hPkmd4R53Wjj4eMr0RjbnVqbVY7AKdlZ61mLPH+D2kba4cgrDqR6Bx40xpl
15LhVAupIODh6RLkNFJ5B6zasDYJlYVN1Bamb/VPiejUOj4W0BU7GOtk5wEw69Am
uowXahU/mci50btzozC0bIaj2jkRILv/f2iauoFlgGtswzrjCqH29/m5+WQaGcNu
u4Fv1tfR0gxvEk/nG4tlb0JMum6atWyWdkSksKOh8tGytadE+0n6Uej0HibJg5Pa
TaY8Fdb2E4rQuqC5uU2suWZX74Kxpm8s4DjsrKdwQHSKBEn00PeaznoDQXLNjKEb
cTRk8pl2DvBHg4SOH0Gldo8LYuFURet7Fdw6DA38ox8nM1MvRcWwcP0wQ2ZX6DRR
0KP7UNnyN6YQnPSelTJQ7xqAJ3F8cm5b4A1tHnE1Gn/dNbA4aOcTpXeU+E/cgVPJ
ENecRFjpzzlvBZdbfwbQvTq/ULQtqhQ+9dj3xV6RNefKlecq0Yl6Fr5Yp5xucz42
OVbD11SONIaCeGr1bFRnh2ugb0fDmOk0TzxvnotqMq+t2eB440OZDJKUdTqsNSsy
RwVwXEh0qUDYZhmtfkOI37pkNYDGOwndRzfm2/2W0ExoZu3g2+vc+6DAqxTxs/lc
AxuYVEDPukQdQr8a/6jqg+Xv9eQufaRlsz4Plw+4ofX8k3Bf5AQoyELCEIPKpDYK
ToB5VjrttqPQNRc3+V94ksc2nReTUbKKyhgufhZVIxro60UNthnnliQXk42eHkVz
FLqjUaSbW6MF7iwnKqMNBPpHICVJGJZZMuTErb3qZ4twIHZNd6KNr/Xp/EKc4p2X
aY6uGp5SQY/iPaAWRidwkB67pqH81oC+OTDYoiPrs2u3jE7fGDEFpuisb6TY+d9l
bz5veBV2XRpgpuNXFEJTUxAbQQfO+N6HLizp7Y72ex+THQyJ7AzyUepOHOfFxyek
GGRl381uqIgf3qrw7g90VP+bbTcO8aFakoBh+CW7qvfKb4JvHh0NCFDxg0CCp6od
S7IpXvlgvKXrQGhELC3S+82L7SYWBausS5AKPUGTwSCxdbC19cztAtvFUXrooRzj
Ka0W5qw6HnZimnrDGJrzJH9llnPl85CN9ZNjCyWyRjpktxV+bZ2hXp11c5AB3wdR
PzjBxzCUp9l30RHO9UwG5LUtTg+d2a6MzLWXO/fGWxDrtEf0AFCVwLBjGy6wztKX
RejZ0nCsY0WqyeMhSUGruLdCLRWQjOW7FZ+lxqwZQsJqtCuj4ZGAJohiKfFnQe05
KwXJhgdXX7b1YYlctSIrq829AnsRLcV4Uy6tYUyKo187QANtmXQrVn4upobdzYhw
UMarG5tzoI57hmcHeLF+Gd/IpQEDxcHXBu90YCUseCyk4I9rZKRIVoWWLwTk5PrR
+LBFVeWpBnFHrGMIWfLADUj0Tpyt1PgV/Mwtbpf3sbcHZpGpkn480C+atIG8Eec3
gHP2MOE6YNRlVGNs/csDtRy4KPJ+N9fAROegGHy4skzqN5/8K2PVcIo7Mi+MfuVW
2LiEvMqkJdZc6FSjk9cqDIPIcJv0wVs2HVBGEFbIhEwW9wcl3N2fJWAMaKNa3kEm
qPpmd9P1v6wv65ZiK3tnVlIkXu2tjf9Sy2mNDBBCL5Rr0ZAe5i6NkFdk954ewZ8x
EvUX08FM1FiDpqAvvNeov1+e13R84aGK3k86k82pkGRouR4a3EbL6kXLtsscEdxs
mpztMz6Pun0u+HkvhxUdILc8YpSDP1eTg/cdCW8+5kfQXCxn4Eds9EPKcmrmc9xI
gddhvgkYCmDKBxXQMlcHTSZFH59kAMEv8fQWRAxq0HSsfFwggSKl6W8uZBOqtmaf
zsgjPDJEj6NdiO++k8qL8YsiG47QjLhfAogCbMa8eg5Jj/v56NNbwDyKojAGW9i1
nn2nB5Ryo79APpSHsCMI3hNVruKHeDodfgJ5xxnmQTJdGyZivyoPVz7FzsYWLYSG
s/oHbpD1+yo3AVBSnG6FGUAohZRJsTDl+j9Lp5HYlGTkxLglaQ6R4BVe6FSJIENn
A6oJaMh6ipk36E7h6hdbWoc3vWvdHzX7K6lrABrQKXlY53AvcC9TX/xCvQmpMe6p
6QzPtnVEwngLASfJg6+QVSep8WM05iZJYlYvX/C/C+Hp14liSQ5Xq1cq1ja96IIZ
dG9rFencssHyeDU6f01gK7gTPmAJfjdk7T+bdcrqpK2Jw+W2fCGu2M8LGmcsXfiY
tbHsAfgObKh1d8PSlG+A72SEG9CM38Yk4teIR8eu04d844LwhnjHusB3U8jKCjbD
Omo6yFAG5e8qLLVduQZVmYi+M0V6PwQqUHox2Y4T/Ua6/tUqR84M5Dc7cotAbez0
1XX8jXG/qpTwd9/OyDWKPOLQVCY0AClmoC0qAXJiDOBPGpxxG+Qg8mAtAv8ktGLT
3Mzu9vz8N4MnXsV0+dL5qb2V7PV2EIH+86OI9UB0tKZdocWrn3uWBQTVq7xxN/2b
x5PVESdSAyLLvKtyfGPM+Gat9d5pjPW+U2et8lgd/xFyWcJKNBZPZ10K3NqVklNf
znk6rPHoCPT90Uyl2RfgzV7aaLMseFyMcuKmQAzvQD1MyTEeTRXV8LHUk3IRcSVZ
E8cDmdWEb7QtC+VzlE7vRdeROGBbVmSxlwPLwG00lRKlK52/rrhZjQtboz2aDirN
IGCLG/ceS0Zcrxg1yvsNeCveALjamkOMNm+XcZxp7kK4mG6HKCX70F6+D20HoUQy
/AAJqgMsz4IRluHTiTw1xwRklZjyBYlMl0QT/g28JbS7WU9kedgpQ4aYySkLX6zI
KJzAGVY2crgzCCY9W5vQFS1vR1iCjWLFcLRYbeLHuLucHG+xiwjBRh4OESEnBoSu
+WC7cO5g7LeNKjNJcFD8rmn5Hb+2svL2MRdjicqGkHaSgxBwSd3CS1Q8HIkanqN7
CthsCJ3zUkIGVe/tqrRfHoxYE8dBWhMtzD0jlIkcIO2mRzPJ777QxYNIJwOvgfmw
r0J1Ocjfsny3BcOOdrCViYwbtLnLLn508TtyP80xWmSkl+tnS1Geuqo/9bHjxID2
g9wl9O6QezUeebOhIAW2doQhCabJ/NNR9chVWR4DCyX26bt+WC52M7yLWj6pMUZU
JENkzZTyNcFMN2t/impr1DDaCQGNXgMR93piZje0CTuUTJKRzC4OZKdXm+WF7hl2
lkVeFIJXD6UxQ0PZWXzGDPOy2GoW7420noVJcAoOH2pv5IOz743rchyFc4uO8V1+
0XHMvstPHNO/CDKmreGBr68CCnO9veBizAFD50RG0iVseTGBXsBuxgI8M4ppYQb7
glcYgRy5dxWAO9MjiMQ2rkg65ruegdXun+DaYAkwtrH32PsWO19c/R7YH6NXzAzn
k7WHcxpZ2m8arTzAO4mKlT+Al8SwW5MBNxzmuFZ6j6HcRlg/mvCVDrmrU6CwGcEZ
6uxqVCqoIU+ITcJC/9Sb1KimtahOIHMAYl/ru3gy/p2Pbdv2aYzi55Jw5MbT3eKI
oZoSwPvxLcPlavVeeUfI7roMQRkCjoJMcw/2bb5ocUm806NzMmVXNrwTnk+d+Nda
etd1nWinn0pHP/Fr63mJL/7u1NiSDK7L5rNv1JpNFKpOiF+B9Q53sr2m0zF7XCnu
n4nhvCqkzhg0DE30Zr1SjBeYeku1lUeztAHgr7ob6UFCK2ytH954LYZSvRv84HQJ
uUc8rwJQyf7KrFAtWXLJp6rRTt1UQ1YX6Tkr8Y61GJ32Y0qGvRIiMLcYSTBgnwR1
VSzQnlsX6iLAz8u5S3vOmgTCKs9J82pNxK25IDwnbqGep0uc7y6bz4TVlHHgDQFv
cidYQZvy0SWXvq0ER/GJHNacKo2D0y779YH3TlLSm4I6S4m1NvcvPdCk3LuNKfIJ
CdiB9iGgpMb8/OBGlQjx+cKjlGbZffxPqw3hS8l+HVOgghqVNC0IMrj62rbfwYjJ
bzuQgprJAFm3bCRObiD8WvVzE+Xhdef+0Snos4WGFYfuKTebmjUjEy5kEhtf4TED
z1CWedg4If1jxYIuk8btBhAv1oIpDsbZzg8n05Qk4T0g1TVM+USmikH22aIFAvrA
ELBIC4ZL0MfYe5c+2zzNgIDqLNbpZycfci1422JRotjERG3FDwpzGLkisV2Hx4JV
zGN3ubTBv+aZyYlY51Pv+9e6xIDIUkI3KOrhtXtfjy32+TMriBTQPBvdTIeBh/uz
5cSmwAlFQwPYdzMxxpiDwDaSLepnS926uxQf6OmMqGkKv27e8mKxdM57lCPyhMz/
9MhNkT4D/nde1/h5fqm5Kd9fFyPruhmrfyZCvDrS+Cu1QnPwG/PlZKv+MFZ7UXNW
2bjsG9FTp1K8GDTo07o5Tn3ieXpwHl+XlHyni+Ao8BACcClcxHdlRn1j0aEp0NVs
EpKJ2HF31IFxpgzqhAiwdi9iLVNTgL6jws8KvaLyZQ6Rvg92Vr9rbof8AtujVAdH
QSoY9O102KVnWQW9kqcNUheE/Xx8QLkOYT2ViLpCHFx8rM6pLYzADrEkUfCmVQ4f
qedIMciVwH9RSIvgcWgAg9TlWLw5eYskKfFDz0jS4x7MIVckl6yok41aDVBogaGm
Q4NgYDMg02c17box1CYGKgyUf7UtBKofkBlvteFWOsiAwsnGHXwFEpvVovXjSO/5
+cPfaqgh1JSUoYOqMRalUAJ0yo3FD/b7tKF+sTGH3h4eY0WH6yANYnctyc/r7/oU
6i2r+nJLomINNRDjRn5E9ihSTchOSiNE73EmEcBYa+s/IxdGkMJwtKEvvvSFOLG5
nl06iDAhNPwhdHC2K4TE54D/DogSIiio5PSdAsKvNmfV1zxtmsX0BdXkJe/N4Ad9
NSIuHhRu74RFtrC+8yKRH+52eB3+iIyBUBH4i+oRgFaWLUg74ChNY8w9laB/AQ+M
pgNZ8IUIvmLPnsQvsUPsAsA2fihZnVKSrTZFZwhYefHVZxHlkA4Zdiwvj2vXin/D
tDGi9VFCFuM5k6QcvSofv1w3uMjXV0JtqWmXzrt9VM/7VXM86V/mn8rnGKVOIHt8
W9Rl0uIMILAOVFPkT+b7OGbX3vsNp6W73FfqdKE25HwWcmlxiZW7dr+EFYkweZLY
DDBF8RZ33bzR6eaUZzwEctR1jf12mtTsb3BbTmVK5s39lkm+loxCYy1jC3vNP/y4
wwZ018xMqaIvAvuHACvFDTpxj2hf9xWKBXIaYc9NaOtCi8SaR0OpJp9CteUiAKnm
Vbstfq/49evNH6utOKsxWN7X7tcnuN9q3HbGjUJSjrXBWEDHK3ZMWnST3z3GrjX5
LGNRAtmOO6C9nLxsYEb1uYW71KeoF0VfjFf0uVHUjRRe1d84yEwui2V/j/+gX3AJ
+onbPLBQBmWzS5ov+DPgz0ne60fsOvlGnI9Q32afTdRxudaqvFKX/Y7ehRjapttD
+J0PAmJktbI0c3kN8lPoWZcq0Ryj13Tp5xS23XVI4XpHlovs6PBoq2Z6acNynKOt
t01Rud0WV2/mRE+Is6em/CsWpjaZdX8SvESHiEHSRhWGq4vdzRdU28QbRCjiG4tm
3vipdSHVIIvu6SauKBN6ps9Pye15ItxqWt6svsBIVTGVb/bHaZOubGoXqonwZA1p
CqZeaUfPKn5dHYb6Mp7aBRS5pLp0A6c9Za8WNuWZWzPsBJwItmKIomFYGspjIc0r
uKSkDzYbdvP8hLxlY3uf+1JR3Ap2CFzqf2jubZvedjxBgV7fRMZiIenwkL0F+oXN
u05HAqIjBTHXVUKiOK/YV81pffrmT3pHHDlC29lSUwC2hE9lieHnOl0U2xyve9u8
W3ocnLw7Rar6n5z39xPkg519Krhcntz3aQl2ITpCtz7sgUQf0uEoOjbv+uvV3PjR
vYmXLhEUuDI/wSBV0nTmqrOeyOtMWxNVSMHMLZwfEEWNFCXpxvgmJK+YqnmMN7vS
giJF4Vbt5Cx0gYLIjmP/ZfNz5qXrJDx5uSwIUJM/rnV1p661HEXDo3TFYmP1JsM2
vM9DdWwr1NvLM5FpEVNCuvX0MnJc0wfUNQ2uVJejRP6aV7l7t0ojTPOWulnkD/av
W7DGufA82TfYCBMzh+hOMr+cE/aae8Gm3lpqBG3OK26T8weeBxXqAnSI+fELJyN6
mWujml1lQpu0Rz2pL5vFJIPCD8BRItztqIhpQ3vKl3v0n//+J/hxBISnalb3/Ppc
tCaIzEVkc/WV10id0sf66wYNoO7LILK4HMtqmC+8jYyApI9sIc3TIKvHrDkjk0eX
AoynqBEwZpCZErKlUdSHUpV/AwPqHucuuCwgblCdjr1BIKWaLSk76VAA0f+UH+Ot
plP1yLaIySjWGZxu7/EABRu9QWMgmbvWID7BRQm9EsdBZQOcdL4rRKcBagIzQElI
iLDUAvaIuKgxngYnSMBD5btxvahMBxUwE6GPQR0jB4qB3R2x2GctCAC1cupYJtf/
V9clQI5jpZhpC79WjuH+8vfaeqPnwxZNDnFiLzf+JDuNFjjlkpE0FEtKz7lkBQQY
GnzZjR7N4Ddr3oYIs+v5y5cibfasiIV5Vz/LdS5NkwpEVD6ZxsSPkFxdUlZfkvm4
6ZmQpASCQotrIFChOqpHxgrEgvCgFrTjwngK6egnXwOVB+7tUX7jUt6Ia0vshO0d
+BQYsIgUKQw6dz6ZDReo+6pxZSb41kluW1eFE3NRBBxhiMEBwMo33WvWh05NI9xk
C/I6v5Z+HBQ5G+HKl32Ylj2pWkjM7fFzo3DuZw7CKF5OpolIAY+dirCSP8zgXRlW
RSErRK29JrEUVEe66+raZPyMoBj245rKdeD85IL/NVRHcZKTh7CrBIwe+yH2L5t7
Q6MET0TRsePntYespqvmjItdIW68g+Q/WFOg065fvI7PDTqYMvnNY4EIR2JGzhXG
OFsHvLei5IkT89Ntum30U5kkQdZ0P/eznXJUe/ThlPgSjL0mA4rJWlgqOOefAz/a
nxuie2kc3f1DTLWVJG1xUi7ZRx1BrvSwnMhiidZM8J2We0UjjSwVtVYpplmYz42r
pu8WkEe2mCyr3lSBc7VRwGinYfVI6n38UlEmOTonWgnmH2I+tV6S1xQ18Vf1dbak
6AxGCcVZdNmMppWm6tLTOTq/BKEWapvRL5t+EsLFpnGWroEsiZDwSg0k/C8DHny0
EyDcODdYVjmxxb7p2GEdFdGaj7OtXjp8LshiTr1n7oxx424QqY8+9KFtxP53b++w
U+derSqpFJPG87qrDFhmItVODAGaV1Wc5Xak4+BM29wg0r7mJpl/7PAGWjMFGHMq
uwkiFEkdySbjwWxKwtt6TaFtky7iaVvYQCiSkkpqnAozwnMTgymNCDewc7uxdiaP
wqTTBxC1treEznrqMbLaTFyrsp15GWEHMyM9p8Q4IE+pBGvOw1d+VqXqDyi8aYt4
+S78IEOy5v60hB2rvk+EHMnRrEAKXHCgRa8rpKNcp3ZoIdkx/eoI1n+ErD3ZOIeQ
obJ/oZmsOtN0jquboxy+PRepcHJmLOuYTRp844/a+CByrGI0gjFBnq8bI9S897/4
SbAcb/UpmQong+5eaPGlwkrHzuaE3nb8liEKckcXkWpg88VqwoKQvY0ehxwihV3C
ZkhnUitP8lHSYVXGUgQ/ZygQ0vDTGEBXXcY5oMbLiZ07wUQsKaBfs+VieDSEjRb9
w0OMWasetMvyBNB71qiTb5U5mpoQxnMo6CosLR3RzpEFGmtd3YNlQMrIr3APYUss
tPOGoDl06WgXEM0NO6I6BAOGD46TP9TNTExuN/PGQ1U6NHMaYWwSG4Ayg8/rseQr
hnxp9rVGb6AFmXyCojOsluF3ZlBlYh5M5suxwB6AiqqrCynXzl7mMYTKQeFPi1hB
6RyNlHwbkDpVOTFTc/slcT5/dL9uRQEmYav1kUU+4NXhnW5bhlsYh/cvtXiPla8E
tkfBFZTT81mE7eoTtMl31mATP5ag78ENkzmiORc+Cy8ycBv32d83p7XrwSYLKIhB
6tJYLyt8O1WUKTK+4SuIcNsuEndyB8c7htsoKU6fqvqi3Yx/ti3njT87rIQNOLEr
0Hhm7MESp2nwoiPf6XfMuIdONzQAMrgXqKTVNKZyapIlice/8fFVoDmqv6W+LOPI
UfkLIioacIi9vxOpCiWEXXwH2XTGO9HBoWoo9oTBhK8BmCtPByq0Sb1DvndvPQsI
2SpqUfXRjeF1zhr6vkWisf0rw9pN78+1d72pgYoiV4O1Z6jUygh16zuf6tMSpl/z
V2WfHKgbFh/eWF7kLE1U5ceCR0hcUtS3sukp078QFsst17Qf6WFLpmNH87KpH2Bz
wIZsuOkMvqPayvVssfdzE/xrGeshVDYp6W7qO+pQ4U6eDrB29hVoqkpt8llwFsnJ
v6k0v6MWIl/eCpwSVYr9qnSWu4qkLGzNy6ff95MT8zSdyiGMvq2BcrPhNXoAKUyj
hAEW/DqeRVRmclYFwaXBImuTgkV/NMhZ/A5LAfFGbgkJ+q1qTkzPNW1hIYYQjqgd
YWwZrn04uY9mLM+UNjAWkdNGRFvidjYxKUgDo0omKI+BShtmRAGt9QA5GYyNBYim
4yrgig2Ma8s/RJuSPgBVjYNsN8h6z3uSYmhCmmtENxVXhzMxJkO4qJs/IyLKOyp4
DdVT68DkUqewxO6d0T5CIuSfnDRbH5o1JApVwwh8VpoMtCGrw1sPIFV2JrQrRHE7
uBRkRka71TmKIx4fQN/6rZWM0gBkMlbnFj1nxa+yyw6SUWW6wyDKFqUTpmYTwuQ7
cmZ/ookz6nhlLljYLUJ4YPAxLLDc8lybygYhwbcvT83MnANo+UqPBMifgP7Qt95I
eSp1K/9yjCzP+JyTHsqmgI4doER3CC3paIVoIerweGra2bmQXdFHlhAfPJ9QIuSP
fqPL0QlsD2Hs5G1eAQ8VQuy9NK2+h6CUUAC6GNrFLByhs1TvGGPX1CbvvCFNo0KU
a8s4LT6soqbittAAzTXRPkesmZfPiGmZwHo0eaxOv4EoC32wNOtt4fQjqBqY3MF/
0+Por1OSca5ggjOV7/itRQ31xl3qJBpFiRAgYLKbZrjS5h8nscixxDoPU9zrnizP
VzPQ8CvYzq5RNWJBKfCNcc/uIZYNdm3PSX8reRLn8vz2+2Ulf9YIGxksr1EVIYjo
TTGkaRbmrSp1QtK1P3MYranc1Et/OO/ekE8MiKVPcmgO0C9q1HH0GVmRiQyUhnrz
FCfQQZHU/q+izWszy7ytbMt70VINZZ3QDhWXZGOFVuYAgp+kKRvIJGbD4qpns7/G
SnJufRhW/xqGUemLZPdTn9JxxqArkvq/W0rBBKd2RiEVelAHE75Q3Pcv80pvDd08
sl7i25ZhI+oxkkcOQYrc0T3WH5Mw/5fJBEecdGC2k1+hCwb8xhwaUDpuySc+eZg4
m9hHg/raZQQ6Y/Lomecauo8MLEHE3ysaktynMJjwtDhWsDmfizGWIeXAJKHAbYi1
ZmLArknIxMvwr0O4yqqDQgHwCuY+MQPlCsZaa7Zu2OKzMAwt0M8xReF1soE3H8L0
JNQiSjuyeX5sphaLhl2BnddtE0kQlvRgynXVNSToV4CE2dYmDKbzRxIh1NSO3Hzl
XjrLTlgfpPs3yo96qNFK1jr8ckLbUCulcaU+FtpWnQtRlxOCD1Zj1w+dTB3PNtt1
u3ZAxgg5MtQc8S/7quoUemyNXaqfFr2l09seFFXcQYvBMwFYEkRT4JvUaNj6vGmE
XLrtOqQtwe3YExpidcxPyu8Mp875zKY3/IAKHQ63bzOuuDR1+6jpPtIlcuC4s94L
NxPN1S4Hyd3CSQgh4KCTuZDXJfy5/2HsxoKx+vKwiUu5OL4yt595ftKsnOhMdVbC
P5wmOqIu/fj5x5uV0Qxw6VPyaNFJQ2YzUHaX7vcKCSkAvQ5tushqByQ/RNUo3/n2
yQa15a9aV8YkHoAyDpHBGyTUv7EFpY1Yaed9j9YjXEqP2cdtcrzhxF5JpGM/oePI
0j8zpNe+5JVjZe3CfRsMQT+Ywb42Zumrcbpwi99avWIs+AmOQ3kJbcKzLVsbefGL
ynMI+ISNDD46eXn2l1CRykrT0I1rB+3xlsT61Q+JTNB/R3bylefDL5HFn/Q3h+Xr
EVSi75l2n8c5hZ8Z1sg10WwZGZU59zA5FIqGez/Xsh4AUkweOqkYp5MfvZQUxnEW
VlLfyXZp7NyHUnM6NglGc8adtp+BkDB/QlOcZGOcAdvyTu3gRzHXC2h4+8ZNtqMH
FQCALS9+O16EY40SV0/FDUG/WyU5x2hfzbWmpF6ahgyqAZ52GGK9iO7ZVMHxHe8B
bOqK/brT2O+QnaKbF0Rwzs/sYYnI/x4vw7yop55zvqKzlaGJHj959kcjH5gwcaVB
0ob8H22o+ci/eYXdsajH+lVj4XH05r6NcxAyS45HhNPaNm1rKfLY6mBDW8c2BqG+
eIC0fAq/gAG0akzbABU3OENgAaTsoCu2noWI2cdmd3Rc+lm56Wdz0m8rPPy1J29a
y3qyHsGDKMFVv4bCYv2bHmmE0e2ozSAjn7TaqGl8KAhH7O1g8jaRX/LI82cc1tXL
40fOHfgT8hwJcAuM6wJ/nUIZ4X9ohTWa/S1o5NtjmhuRUOK8i7Bv6YRwq9PnPLf5
p8xj+LaXdbRQPuNv3a8WBuebIqykjlcz6SjzVdAkyyxvtPps6hxIjT93sJPUAtsl
06Qv7qwerf2/fx+tfX97Ko+nDWRUirMg3kd5zhl/w3A4u3mVu7nbCu8Ta2GyDKU+
MZCIsZzuV9PcCXk5dNoN5Easz2cN/0Ie9kQzdg85so54tWP7Vt8Lda4t2dvGGJSb
RoZ0xnNgpkpeQL82w6kwWhKC+GjUNFgZiFIMO8RvJGYGEmRZXaS5zKFw0QNK7qAe
KvvdAnIRK1FTXNUzPMEe2bsBuoxrRNSCEsgK+U/SuFRxM884WIEAd4WxfB76bIRW
TAXIiVNvizFBzvwoov1Fk7myAIOCjjSkhaQjtt6Fx1UKxvdSUocz74yN6HsgDb5D
tmYU+dpK4SYMAcX+NzDY0oHpcV5tUKoTHtnfUo9qEoJ0f3JSXUcziAPnVtlpuaim
pMd9ztGam9soKwypyCdqj1Xx/i/O2+kK471IpQ716uizi54efPLHLUGIRPLEU8Uv
QKy1shfaCyCSAG4qT148qByq7OJH9Zc8TOhx7dvxh9FZab0VlERK382IytxGY2Z0
E0MgBq5G7eSnP/dlphv7EVxvrlIVcwACs8hXnRwoEOxcIY9KWdvDMwaSE4uPmBj6
BCqkd/BzPhdSr6V20QhMr18r3YinuC2WaaDjLuN7TujHSd3po0A9Q5S6Z2pSkyvx
iVCo8VU2yhFmN29F2EYESFUBLWJNVYBU0qR3NoBBgN9637zD5NEZRu+xpVAP/ipN
jEBry8gGPxatgRxEDuOkjxtbCsJDZJT2LfjaIv1iBlzaGgLKjroT14v0jh9+af5n
JWHiHlLCoSY9S4VkSxHaHNsSrizCMMRMucCdo3Xh2pJ4mkTkXEkRByf4iNiIMcLc
JWSnq7uVQUaZJNV4ZoteWNn8Bkg8C0j2LeikNlBmTlUedExF0z537ljmMg4hokK0
7bPhoOSrAOmttO0WbrdwIjNTdDuSZq2zL3yiRf0s7QKWnzslVoHxCXPNXxZWjsh1
IWfZuJ0d9DpcQGHaZnPIXDMkffDyPepl64wNjXqpEiK6lN5lapBjHAiTe9uyotDw
G6g7gmpV+zDHCJmc1qj6anQ7LvBrhFLyV0l+tWaXDAgrHo5E93uVPeZmhidI1CRD
jEsnwzhQjsjw0VoyvN1agpFY8WSODFWQbeMowMxnxjYS4pX2MxbC2KIzX0e7IQk5
8dGfOWbi+ccDFPZOfc+NGkgpvPxiBTFpfUvjS7kaSWpHKu5Bzmta3MTBVsN7bdtu
HF+tJWiABV4t126r1SppQoDIl0dDktYiXpDWqTaIbBFt/fKHl/VX6FCq8OuqAmF9
3ElSjZkCaNzNhoGJNRElAsZdSj1d0y7REu2aFjQrwnuC0RcGilq1YJwoGJZQeExE
liAiCYIjgJA9VbPlAkU6husYjd6Wufqbs0daYN+rQRBXoAxq44Vxf6NjZC2hn/QE
U6fdmnhkNZywr/YWHGuryFlaN5+WyVYyn5yI/tcHw6MToFlx2jUq9pW4uNLPSXlw
Yj/0E38CnVbFot86swb9H4hcRwiDmcU0hZXYsbc53vtScdWkfmuc0U9EgvWFVupu
ickTQbiR1xu5xziFcpHFSELbBAiAd56hb0R4gAkDSGxIy8DTohxXAKsLdVrDkiBy
tlkZlhzIJ1XryU4ufbRoiF9pxKM7VoULPD5gxb2wm6V/Jlnzr7ebzO5IuwbwyWU8
HB3OROzc5QtjglwYgaD3h8e/xCiTLmeGjvXomfPyk/6Bwbl++XgOUte9JxOvtRex
nW+Pfw+cuJHHWh1xDZghiEvkWgJw0sOU2Qa53MzS0C1xXyWpvzujgaZoevKZShdz
dTSpqOEKOin9SD9hjEz2/C7t1pU9lwvwzw4rl/CcKvwUfwBenQOhfrVJPMyeDyYQ
70AWbM605xqf8nDkgYi7UYo0fpPhWXTRh6RfVRG3iQzUNCPpiAGmn9kmsASIVRAV
R8FxUDYhaQ0Wb2v8+WATpXFycfxc8hEPZltmByFDCTPL9Rb9JPL0WONn0E05XmE8
wCi1ANDApYaRCqWoZi6kn+KT0kNPyAGexgSHP7/SIRURRW+304+SYfPtuqoUUnJG
T/wdyPAymxzx2d3BE7JVuYriCj52O6Bm5o+89TtTLoNOL93zTXYvUx+xd+weZBHo
hw+yH43JOpFp4Rx+A7yJe1lXOyNkC3rAnM/ld6s5hxPjuuOVMjm48nFewbM9ssVS
ns1wyfIGSIEjq66Sd5JSOXGisKLESZiFcQ8Xu9zh5GNgG249KL9Iuv5TsLwJyZfJ
OvAQzNb5Dl4n7EpKMrH+Q6pdk4HjE/+QTg+ADKU9vV63tk0y8exWkl37Q7UU8UAf
cB6fGUK1/Syhs6ea1ESVshp6Af2PjaU7yzuPo0nH6yq+O2PVdPWAay0tBqts4664
8HtNd/zR5mtztO0vuyTIW96Afj9PqV9qWRJyyAareEe5THhVMFigY7MIHMLKO4Pl
V5dMq3mbnsu1cmAwMOCstq9dcNCCcIGIUPPMN4mJOKVkMf5n6V1uqfytihpaxUj6
qzY1d6z31CigZjPD29jFeeinleAEEG11el8z23wK5VMUQhhIjauiIw95XICifzqB
0vKgpPFIresWfKru7iUBzwQxPplav5HM/7JIdTLELBfPxxephEST/tWPGXuXkl2Y
Go7R1LSJ/t4qUIKBVLVYDwjRXtxSxpMnXQ0J1by1G94bOPb4j2mCfVDs+6OZ5FSi
/+rs+vxO/87GxvTBk1mmuO1L9kA0eissK6fS7j/Ynh29s20/c26/xFvDNEfh5g/c
h4sOt5u650kw3MbxwFFjOW3tb3eayEr3CZCnc6cm75pPczVxwjapISbBBKj6eWIi
NUs4jgPNl7KKtfymk0Cj/aCW2J58MeSJH4KF0E2c3zNZtHyNf3jpLePbJI934iLH
Zck+CFqRg/szbG2v7ucfqclJ6RTaeYee1eP6cVG1QGKci6X33axfSKI/0Y56dwjy
CvIw5xwc1lrSM6kS8p6h3fstnEXmqR/Gwbn/KP5GsoP2kqf8qRE3S4X/iAqySdNS
/BgGe46tpLA5SAWnkewcYiEbsej+sC7BjzQ/cl0AVe0gV+Dv0O8FjQbTd3uTt/ma
23qRHxWQxIEohzAIQyp2BrotFqRcCKkOntDmwFoyMMQ6pWGQTIE1UF/mRf/Rxy2G
r0C3TBY4ugFRO93lo7B97A4u41+lLl85lFT8AkKfozqPikxJvZ3kthH17dDYEQNx
3364ZkMu5t8Irh2/eYZ7PUG2CkN7B4ivsy7ePiZtigUke3o7t5t6v7LBzpMNeUQz
25blJvN8UnIisIU9w5CZut8F8b0R/sIGazebKXol9TTY7o6BcQaTluBiVBxV5qn0
qZWuz3qLPpmUP+XLsRSXB/1QrtX8VZQ9rGFDalyqqx5c1unD2MpNde1oxNhcKI8T
cQIsC5WpSTgpSD37n542VFIjlCDogvxVo8Y/Yz1LHI9zEiHTCBg9PNOYsFo6b5/W
CHry8FuFEJ9L8xjU+g1lfmuXzN6r5QiKzzYQTXbgT1d2FAq7ktNh244gRNkc/cLL
HWUsIZngk3Q/qNn1KnU8TrccgAoEYRjhFWn8jG/7GHuPbMurUSqxUKmIvnlI2bZP
QmzC/TQLvONUcC8tou8sylxGPT6ZT8tJW/aZzE/VGaHqYjTRxcfUk4voyapq+Zhv
lJg8s4XktALsDpVxAaINGCWFnSEa54SQztLP/RFLlmk5eA/6ZF8dmNRia8nsemqM
H9YrK/OTsjjN67b/PLnFhDk/1szLL4CVh7x7feclXhRXVbMTxD4RbQMKavRHenhy
j6dzK62bIGHMq4Fq3B/9pBOyRJFAU0FykjBLqDTDckfIy63ufXlEsQtuPSv6yYd5
1xacxGTDXTCmYs1OyEItdIdAts+hWIWTpEkUL+WRHmtigjdUDpKknRzkzCoHimvp
xHQDtT2DK0zye/mppohWoQdDq/cUMbgKdAdkFLOfxcojrh1CzEudduAolNOY4HaD
hisIHvYp70czEOV/ulqNtjCMjpWiQefq3fYvCy/WLDF3EuEPPW1C95CDA9PC31aw
wXvZiw/wfg6tB1mjyXTKOXh2VUrD4fmTYAVJcwDc3k0/sfH2X5hZB6SddyRmZaV5
MLV3q2NfGE5GwttAAqqonx+8EAFsqVEbceEme6fd8C90ucDEcB/OolqHbMioZ0Io
anZoYGA1Ycn8xFukbqE/xv5QxiKEejcGFKxAGOqY+V/EtzYFiXKocmqldvr1fbHH
TBVJpxldM3WUXfMzPIGrQsIIL0wo+Jq9JdrevLjkA+f7ZwcxaKdICnBFNOGqGn1F
F2VhhhaWoQdLsc0buxCKJWxueAIyyJ2ozHFs/0Jl++rub9CaXIKYmK9GCe/xOs88
FOWrXSfeor04PbzioNulIT06wzFCQQG3zRkmvkzVfWGTn+EHivJO+hofNsT8jo7N
6Yuq06/vezSEJNIoQSA9UcLcAeZ3C4iN7l0EdvATvdUOuw78tRG70F33lVjo6rnZ
yV1O+LhXfNQ8Bjiz9qg8+NSdZctKkb45SU/43D6X1Jnrq4vhg2dh4I08uNfN1KMH
+a3kz7k657roREL7uzDyFU1kRaghV3RgegF/bhyvZmP/OZ7oMcPz54lbiVkADarB
B9XK3oRXDRZPlbMyB4Bhto1M+/NyTszx/0pjf1yTrAT9wBFE+NUseYVEt3vWh5z2
KzDyktgtaXSowD5QTS/X3ZH8ItyXkgwiI1rl8HVdm9vfAcwyMJilPJiPALSmDu9G
NS3CzLe5ZDk3ypgWFZzwSUJWCUf3zDjojBl/0z6BAlTnnZ9lgyfMmPXWrjaqbWq0
3NehLsZYIXDRNVkGoVtQqfd/sm+Idww/9QdKjG9Xbc8Dc4Kd+Q0Q2OgbXWzVft1m
Ic2s1r8vjxRbnUVFb1WTNfISDRkD+A4kbzBTPPTuOtkJQFmappf9FlhuYsUgugfX
W9SS5r6X+ATgczA+CAf4Ukoi8fwRpbjpQPqUehMKnXW74XZFqqF0QB0X4/ldqjSk
pcwU4p72GEVVaOcZiDzh9Lb1GScbA//fDTpL4JDhzGvxiImiWF8R24f+AXqeAwME
dAkJdwEe7pXrRqycEDAEfXH9Danm/45lsuXclzGaKJ35G2cJtA+zocX292POUiNu
K+Rsf1r1Sx9gZmeYmJQGDY8ShvgpRm607p9lRri3l9uEd4vyC9/M00VlBq52BuA9
xseAmArBKwktsrg5zePciTFkeq8PCym+xrwyRg0fjdCE4ISXhmKB0kA9FcIPc+Dr
heAq9sbUsqCNKfuD+oDwpef8wIdASkki54GUaM1MAZA4k7tVLocOwU0FTIgpg7tW
/tsES5YjRgKC4ukpr/HmwdCM9x61Ht7tq8fmTwjjOtay/M2eqrNqZyQvmBPga8iF
JZ+Y7PPq1vrnc9smeb8jyEXqjwpQqRlSfVcdp4A0h7TPhlZd+ghyg7u4ExtwG75X
IGAUJIGliKAugbjNN8ngM4dYcb7Rp/vgYFEVitZQhqYCP9czZJjGTS6y4PLClC/n
wG22kzZ5VSk9pie0pxpbyN1T/C3G6d+Q6A6KPpY+CaRU0zIma7P6NYCE0OpDN7pS
mgwcyiS5AbppSNyQ1DntLcuaFyMvz0O45UTGnmhuvMWI+gJMh42yJXbiyxPJn2pe
kayJn6aCG/en6ZiKLgYhXx/SL+kj6rqN/UGpLXple6Z1jsbe6n2dsnYYqMkXwAHd
quQXH8LsOP2EKEBniUl3krLlSBx4KtSAxOwd3FcYtxBVgzYWToBq5tZRA50lJOUF
AQ0/4jRSUS48lNgUrCXYprYtjY9ZUDjCvq1VYD+9r0BRpWEZvGiUqqswQDA+yxpK
JORmfvJGnbKyP+LU0472jd0dEr9IpMZlc0dTjI33s6epo7ydT9IS2toQsrpkKTxR
Zp3JW49qkabl04WVsaBjlayAQZSohhkzkuL1FdtGK/RQ/bic547+TwJ0iOkMhzwR
zQzKdSRC1mJRptajLragvxYlHr7uByIQ63tHWP8Y7wXehkfHP2MLSvyoDd1k/EBK
r7OeFst6NipsVgUTBVJbpvziaqRqa4iBFVV8W4n9TNf1S/rbD9cp2UfwkMq+YsMq
b+gR6bh+DLooUmOJJMlxSQyXmir3YAsHTZL8e8OeqdQk3JpbiD/nF3gPvrqyOrIj
v9jPlFCHUXzVMkhdLsZobV6zUg+MbV2a8cQnVMEQpxHjihIlHSQu54xU9CVSCVkm
XUbrXLChdpwmMdfB0AV7j9pWRNo/lCvVxddPmVpjAguMteJQDjmb8L0tr1SUd+tg
xZPuGh2kJpYh6uaLl0bCUis4t6QDJfOTcFe7vlX8dp3vbN12vHNOGCdRaQZPdAZf
1FXLq9R4PckHQzoxXoypRhByb2ktI68XdL5cJxuTerhZj7R95winzMUzIVSfqDlO
O0rbJtUAwIYI56J7xMa0fhWRBoOEhDN55/ZRbvttXrbRv/TSmhBqOrDCjEXDks/u
ZZIQkAvW0I+ZCxWhcUqF7U84F+Hom5q2j8+xQtN89gRGupVllcXenhUhcfmoOWCP
n4CkNiX+2I1OdHh3C6FcZF5C+ZbVDUVLD8dXJ0yB321shGhjsg1orOH/R/GrTSL2
QNPFyMCoF3acUs01tpWvgyicwOVW007024yOzjTeilroct7q3LZJxrFyFE+14Asd
IAohX99RQrpzR4/uvpDoGY/rePHTwFdZFc28attEHHsE+snsOtOPkR5fF+MPOcKQ
ZWoemb0obNkfFqvTimunPafnKTRA+GRrQQEM6/Td/CRm+1gP2brzwfB4fyCrLXIQ
uO9dBP0iIvzqA1h0CVi1EWHuN9GZKdWFYEeK7mMV5Uav54+X3QKWFO2O5rv59RsS
M2vjW/Zw49T2kqy7jjcqWoI2OLKkcrqMWdHvthX7ezjTzW6UBNf1KJrUqZPZJ/iP
TAw/F0IOTCsyIyMrecOhB4gmaWiP9pD1YjNPRHsIlv7ieTFgm4qtIQU6+nqcWcXc
d/jbrb4kRzHijaa0YXv4HIOD8TCW5zesjzyO8Av1+XeB2ACUjGjz9UK7HORNaJam
0MD+2ddzHozECjPb/DhbIRBSE8OrKwI+jWE8fBxAn7wzQsfMtUz9TKQwSAOtw4Qx
ZG45iLr9Fe5Qgs+v2aKsi4Z+koDHNcx51Xn9Ol9KPKPC8e+DJzigGf5XJysRfojB
oJSt54or5+yxYAh4dF21XK+NCa9NUqKVWGLVfLqmpuE6+Px0XoBuY/CzXy9J9Rew
rXQRg/suUvvnuQQ3FTAPpxCjzGDCcClYkJwTaO3p1D7L+K0SHWMCLcZgCF3V1iE1
Ozud1LXy7vn6bTXajd7ZAOMQvmjEfFUMATzDd6/WhTPgj/dl8226z4nKESGdCTjG
PyVdqo7h/CucKw8N1+r5BSIo6jU0Qf8QeWcHTkr6Ea84WDeALoGC9kwT7anJ8R79
9/bKkiUClzk2Czst5r90pX85Xu6oFp7grvJFV4dgT0c3bq1TPalyHJYoo4YdLs41
qudHs+VfQUGqK2cbAfPq8RuomtSdyHB7MZ5cJ0wTzi128hccsKPsOFLtVRjuKO9j
nxWjH27AnGXuA+RjUalSL7kXK4B7zb9r3JobRNbfPgyv8Ms0SVpVowr48m/Inl73
jYolw68SzjfGRYb/DMQnoVurEo02Z5Em8+oHwgW8vEwAXGkxKlEvw+rFkqLL1Jzr
C180a/2YaC09+QJpB/IepVXBxw0ExsE0RJPJ0Mdi5UiVDypS+jtTsEMJn3rZwJ5P
phWXvqQ6M6HO76mOKFCXXW343YMMT3QADbz0HPnN3g3VjNn2WbNsIyDctuqlHtAW
5qdtjhbwjqkYukUCh+OLlI+2bPtkL5FkwA4VCDGoj4mTiEMSqj6pQ8plm51S5g4q
P24xj7U91mmme7RF67OyK0xp0gyojT0Pp1NuntDuoxcno2Y1K8qJSxgK8hu5ArLp
F9tPZjKVXhxlMMlCI6IJsNLyR4qxuXmVHqRWxwBUacKlAQGnX98hgnrNX2iynVYw
nlfcjPSIqIrfL05D+4R3Hl0v72NlxD8Aa2In3gQwYztZdLihA94rwAapE1xHfsY5
WYjqgSUltDGP8gDQyEcedjbk8TA02sejVHbGCdw7N6wbxWw+GEUtMUPef648qrno
kO81vc5pUEAHqZCqEDSbDtGxXLG1gq32S15qw1EqNZUdept3a4LaHuAFCzdRREMp
lMHBJVULUnOcqYT1+ckcYcmMom6x094IvWO2ApsrxadegmLh4/IBGV7fAcr+Un2W
os/BKDqmcRnsVwXFn4SMSt1kkq4UvhqT0P3+kDGOE/byy0+EGj2jYX7gC1qWnkRz
PL8Mn9Bt2w+fnpJosoJ/tbWWtD366i+aQwrEnCvgi4gQQpYXMMx1/DxGEWIfatRu
WiwjMeCbIliimqYVedmn6eOw719qNVPhgLa20yZWV5IR3lnRk7t/9a6kHMF0IX8c
8cgY/n/+/mb+IY+xU06s/D0pjDIKBAubxdTnklj4BRyc2OQOueB6qwXyfKcXaBOh
g2Xa02AvtEX0Ky54CznJ+13w0yR7HaOGcic2BQV/4tm1hRv0AXgV3mWMyOv4YEio
pI19bJkmXIBhiJPRydxuSUCezmC0zXn80+mgfnbX1xseweJ4hMiV2rHN6Kwf1GBT
0W0BRUA7mhOkxv18JIcIPgGvlg9JHCLvd0TaP7T2J70SAEtxO/IpOgk56fD2LjN/
WaPWC72vCqqonkQ4R1ewsha32PkqKVfW7WzRz6pAF87X9VplxJleePtv5H9wvWrR
+L8ehyrQVKYlri5vuwYM6FriEn050ZxfIvmR435gr6gz7KYi5TXwf/KVpv+9rfxw
k1XvGt2NzAMUxj3gw7D6bmC6CIK+of33teb/6IRsQrxzSFr9rXebyUa13eog4WUE
7W4U9LeuivL2iybQezuxBhrHZMdXeImVIHa/TVxjzaYpzvOYSNY4eO1rCDkb1/iT
3JYdxxygQZdeEQdNwVcFSLqpBoQHhf/3MWV7Udq1LyUDWsMWlNfTO4GWkj/nXSeY
sxER68/2MYyOyPsrvbvxpdc3n1Kf+BSwfaW8PSIFa1g/T1ZbKfDJvGS2Z2n1OI/o
dvhwHteWjJt3dpX3uiyaKdpGxa6pllI6mF8lwr9g9kUX98qbl01g0OsreWBRvlhu
ItmtVkARDsjEvBWu/OjpGZ1EbYH4cVjc0vCpP8NUQAs+5UzBJtP8gs9XUKV5ohkC
wOgjFek2pqqeMSaQS/aQtwHDHrQAAz6LWS0+PjblbXZ2SCk0/yDsebeGPTNs6M9z
Z6oKue2I+OvdF2gd4w7odZkVn13/dLh3kdq4egjUYG586AK6GwXIoPTfHgu4NuOS
Qdu1bRqqqIgEbJcfs7e98vlFAA32NHTBhtn6woEGP9BR3XHxZOJbk8Ss3/B//79r
mR5DKm41ih64fCIoOq1ocxGOlHbOYx23E+V5BdCiudyhezwMvSfhHbYvZpJv2NKM
Oz5aztAwOKWgpRghwxUOZzrWa+I39a03FkwIPV/bbVIGPCZ1IqLlnQSpKKtksZxy
WkhCBri+zQ4/WFpvPgvACaJGXUPZa1zt6Zux42NFjs/TkQG9PUvRpDLnP0CW9FpK
H0oieL3EKDTEcPHMJB/2+0v+s5rfnt9zOhGPtGFxPQwycxsqLTJOFEKswp/+HLdt
8bh+g1sb2EigbJAp/7eUfTMzez9D39oppYt4UfTCXmz0N5m9Zze+R3RJQz3V8c4Y
ZVYuIkRkaEY+SCJjEVpoODl2ZywedJNC9YwBRPbHGoTwraNWq1J75/bVBWWR87LC
fnhXZ+eWjatZCPgeHRjU6FWSwHHlbxCYDHhqhp7pndzTuwFV/rpVHeH1+pEe5rCv
afW3Fcbw3EfmLs4RSRnuYabzpV8gIjUmwPzURCF8mTyw3Ltzsy3Q9jPTwlloYPmN
TiS9X50OgEJyr5nhpMcYi0j+lXf66Y75DCbJmokClVyUVuHAWdNNxz/aeWksiUXa
pL6O7M7XjITOH24YPq5m/NaxbWutYjpxV0CPxiYE02i+h+tQfQ5cIRbRYZxvAcR7
2x87UVFLOjUFWUo0shQ/yePgc2Ya/q+i7ptliweCqIja/88Isqqnz6L0NCYMu9Zq
ITsMK11NlIJWf4z/I5Hcn1vV38naJhZn58SiC7q4pf3/PbPezE1nTF13pVbVZpqL
k6UZJcBMg1JXvySciQWWIkbO4p/waaIONNfGLTrWLv5ENIgkpOkl064ssoxcBb8+
RgwVtvGLWvz7N39zrEyDWDaFm3tbjym21U+hpOKZghk9J62pnEDUrbNIsxTAlZD5
gDzLrcEP/wZN372X3JDdu2mFM0htQ7nRn0XD6JpsisAR+SrQTsbXuo0+0lMsc0Cj
38SzQjtwUhpeoWw0CGQj4TzVtiC2nGSx7CcaM7n1BLdC/E3UfXg1hqOuv/dpTgC7
Dt4BSr5Et8PaVttS1b3GG2en5k4Xc1MsWKF5JFBtT6XtWGhKhd2Wza7ectGIWB9l
tcofVKt0gTfr8ABm9/XH+s7CzRVYzM/2m1SG2JUV1xc56hjzNqbhow7X6mcAq9Ik
uwwBIh6ipuM1m6xAU4X/VCOQYQlnN8ue0W3UrcITFLhWL28HW1VMKEG/D5qAmCVZ
eJCqfNuwK8uNSQGJUr5h05BWyifLZWhy4YRFMOfvHsQ/WCo3iYAwD4q3Xm+qlP4/
Zz4Mr4SKJY28qbWm+N3sexOeCxEC9ditiaDn2BT498fW5kQxnRAOqhchCYyDkzyS
e0GkfO9ZKKoljzUrg/MUvlQtET9lHpEBd7mgaU9wLd5DHJfABXjK1jacqXzXAKlb
PKtTNzAogKT4xCSKiqbppucQkhNoVZir27kRwRo04dBJSdhTaWLJRumaJVdFvjJK
Kq9aOUhywFJAmprKLXoPDwz94rPH+u8gAMIq7effCnrNYLICRLYTECD1LpU5Ndvy
GZzJdhXX5yh6x1cHjp+hhJIONlgw0Zi2BkZqCMULYr1Tda7OZvIsbvcm3BPafAAO
G/2f2agpcx3iQitZIi3obWMIe1sN8TD/u1H9WQw/SPF6ixhiSR6Xfegl+rchtCQh
o3uSMbcx6yAqgPBA6wBYrNqIbCoorIF8BL83C5FpBExD0Gu6Pb7mP2AfDkRcn9PB
I9LqTgxWe7nyLW1LMzWlV1ZhH5zZRoiGC266nF53KEEGuxt5lU951RC7e71l4wv7
fq5elUfZDUsTaa1Ng/x14OZjsQsnc5vO85gwPGnrig06FP9gY7BKCQBYvhccrbnr
Y+0Ni3X92Yq5Hxu0y7wrG6cizjpjHEkYbF3e9CIXCo2MWf9BtCCOE9TalmYMB71E
uBjnrnDrz3zQZOLM0hftupuhMbdOtTNsoevwoAV+8fkUrD+QgQ1MG9XpWpi5bgeN
SgMTvTG8LoVj4CewtXVN1r+UsfFg2OFcV/E+b/MJo6xWItgGKyXWZXNsJ7dTDV/I
Pv2zlkZZr7VXfX2Oe0JkP7d+W6E1SJqz/j0xjr/e1PC7gL6HXDg5fKZlNqjncGFe
ePmJyXkhzqg9zB1ennhl4qGNcCp/6CQcOFr/2K5VPDISVW6b9tfvEzfxYkCoggEJ
6HVTvs7cL8ykCqGzSWDoFJ1yKZhqObNf3LjNipsdJLy3UwZN37VfXtYHUigV7eOL
rJLzVnWRaEYRdFyFUWQ/ElXZPOQ+Koi1QJBBE93j9YQkLQ+5E3pQ/MiBt3WHdAeE
NwDHYnwkKUr3+5OLT9M7eWLdWFor1XhYxkbAUt1YyqMQEuV/OM/hg6FCrGRytp+k
uh9WgZuxB+A53zjvwtYmikZRyZQG9ahTT3MldVf3JAcu2f9wUctX8XTEzuD9W5aB
UBEzuf36MUJB9WaB1zvfWqMyJ0lmdUSGsn66+pgfbzeehuE1tCR7Rsq1e+F6gvYk
IWPNl27ngmW19v1GSPCRmje4AeTKBvncKZUbJoReHZ1yiSOMpVRgfRywmy+24OAV
cRo2+9K1g37PBfIf4k4Rgzw6Qch7pYy3mT3M+EpfGdNCcE57mtEoQySh706xFfIm
TfHmFqa1ucfQNBymsNKcXVQ+8M1BSbNZxrNNfoZnpLeSkC/3JbxpFu3qnS1lq8E8
Bb+WEoEwK8IccxLt6D3GQVyNLm3RyTgNN+Wgjmlhu+XtDwktAZ1JZkOVtIwrmzV3
/JVoABGvt3P/sNdi5ubuq1J7+U0rAZWwxAHaoHWxxd/l3Jto48Sdc/F9b5L+GapJ
zyNdWmRCiwIlrLUPODUADcM6yv/0Hr//cjGj5HIvoEveU1C1a0eotmVomOzguZDG
tVywI8P23xXnc6pAfs01kHLa0+Ayzq21f0KkFd33FwHyED2Cy84w1lAdHpLGvQag
3A466pyNdAQmpLJMNFc/+BpuASrcDbxVwG43Zmrqy08LY0k/MOZnKVTYqNtVub8s
qdYpRdMisDEMwKbHvSW5op7awR+FcHmjQ0EFnkgPkB6ghLkkogaru1rH5B6VOkF/
IlH+pBmFW2JOfLtRGybnWWrNyLma8SsZReKh5IiSsGrKuR9zI+X+K7RMgFIJRuL6
3JZTpT7RVtMGWfuSLgGWSMpIlWsrZkTu+DVnw4B2UmxEBkxHqGRTpQRNW97g6Jdn
ijCMXWTxeb06WDJutocTVVUK21y8AaUnBF+44Mao7UJYKy5E2nkC8qhBMkSbLg7H
E6RNNqO9qRA/4y9wCx7lMMPrKeW5drPdcsseZ+5cFeo01gzmsp0bsrctzjZhIXbK
L54hb1NC6iATMPzQTURsVhCMjRvoE6dabVg0f6G5vaQoC0DVpCEhx8xIqBO+1fEa
0UJCBnEnOpz9TEbX+CWojxEI+Mq5a5kLGtduaZ5WKNgy9OmveG6CHpMJh+3ks4Xw
pWdSi5LZf4GOdPHnJE43zSYroIFHEVY9/i9SKcv7SGF5ONU90ThgSnL7EGNixatX
6Vq9QbNYyTetfyATk6fZRCakf4pb1MMttzi3zqtgK4eRLKVOnLbtLLeofzW0LTyF
So9meLnlGkk5E6v1gMDru6wkuwkbR6NmZ3DmE+KtNtPDuapGUrX7zVkvuFxnLVnN
+qUh/RXmOGnIFV4+HXqKbBPfyNErXdRNjoNjb+T2yLdNpCDFBLn2M/MEi9bYbIjt
6DUiO806K6DG/clAHG3KOc2nQ008WtXU6UH3HjNKpSNMAsqifTIVG4tr7oBHNkwC
AoNzwLKC0ATsAn+ChlwRnlE12EIiHBEZ5AZsA9s8G/ONN+P37Z2KR68g1hRFstqx
VhL8GgeMAZSsNnXNXOn/svehHiZbusD1xljZHqKndWqCVeJPYmWSawrecOnmKIw/
4tOmVlGtNtzsxEoBXjeNPoyZY7NnIrgVp0OEOYsu7fm4Zwh9ti8CtKd+XQZ6AQHK
thY1o2wDy1WTdL+bYVEW64y3Jd32zvzXQDQsWUZpohaf5OrtMY3NHhzvdu+c+t5v
cLHsT8Y2YNgwkVLQsiEdsnoGkMJhWylIiNgdiSaArcYzCNg9A1I1nviPKr+UlKvW
QUIOO6Ywm+nVodhRUEPNgauyyt0n+cia42+hc11qTFAZ0ZgkIcbmgEp5yIJ0b6eq
8z0g7IvOJRr/ITGGJueQ+/1oQ3yrBWR5KEH7Hh+HU+z/tBOUwKPjggmHU2FsuIjA
JfayGyrhmmUl3KtM0ZfTVzzOvxCB0+rmlUgsLFi64TeJSu6jtMM5Kt/dTWC8wfFx
RO5/u7BHsHtnNhrd0cWQ3z0YB3bA3/bjm/Reb3tude7aHsSB7yRaz/GTBqRO8ovf
6iGZ/KQaIcqisW3ucHTLzTmk1tg3+I0GywlE9sywRznX3C63yOxEV2zAa+ZT1tf6
qcV+Xr8ln1EdB6N6i0rR4B2nu53OmAog96LN3cYDoeUiDjBpvZ5B5YfxyMFmMhog
q4eFZgcpEPf3/yNr1rXj3oDJu4FT4jjKiE8a2lo/B3ShEhIMQ58QzS+eqHQyL9es
EyXURlnCsz+jcx5tDlTBn9t9Twhr/3V6rIpLXnzxAICHAGwb8q5O5UaJ2UAv8auA
/iGNOF4/fl1n9yiGwE9T/ZZnY+uyOotTVMIMQA44l798lJB8bSKRQSq06i1EB+oz
N68P5bsFsLY1TWH2oEOg2U/FWzQYhuDDnBX91ZeFLc48ySv3Ny9WnbOthXUSuPOm
9RWTeyUUDcWIvZ4XAdYb0karW3GS1Aa8hF1xWbuhPFtnUmIyD7FBbE0kMVBQ+td1
RaVqzuNEzuOwESJWfG0yqmrgcfOcIvsChDSSXt4uhqudhkD6zbi5yWY7/FnSqlEa
s/WFWhAKmwy3BA1xRVikyuRZrykhh+cKVkjss9Gre1/TFI3uwXEDGFLQ0qi4ChVL
7H0pp/gxPEfRllJddyzTUl39tET2qdOVu8T7p9SMa7Lrh+6wgIpEi83PovWt1tpU
r4n2XDn4N6uYiLrNWZ5crdqlDWUy4Veb5SxXh2907Nv6t3JaL7nt9irjiPneeGE7
fq14p3rm8XIr2YMJbkSjWbSqNReQiTeLmgba6aNtq7EET0R/gRvMKJfOeYKHcupZ
N37MvQ1dKdphXSGb1P6vXpPhw2A+8qSBx4C1+a89Wp2bSy1miGVQvFHVy0ZJNaWa
Eiys0IC5zYBcNHHgw7+3g1NEUINJPMAwHGYtv/iFUcqYzDs3SZAbU7L4u1831hvU
TO5zZr4DEXhqKdi9JtbJ5yD6f7jalPpLuBoDRzss/9BFkfn5psGwAEGipLuu1QbK
mjHP+nhD9vPOYMetHZijbq3SQOtqerVfkbkTCwnj7VlVc6sjJmn4YzP3IQQLZ+XC
XMr8FDnB8t8bgZqco/iTpS0ZdmljZVCVmCb06boXSvMb+BQGPWNtz8rOwP/kcTOG
GJVeYfac9bjorZLyOgrP/KWxLW+dPUpeX6iXX9hwjMvEpbg6R8BYsvBvTjHMmxqR
mXlj3TBKybzwOU/aR34u0QHqll6QJlq5qVDd4wGRbrlsssGa8UzXIvrBcYpvlSIM
BZOReXf/OJbJul5iXfgTCrjU2ui5AqQNrk6F8TJmCIvDPWZ6S0+cWhE8lJKVQFKs
j1BvZEXWMknjtOOCAq2mc8vR5d+TE4GMDOKMMSFvSzXkxxEejS8wHzr484fUkYAr
Y1FbCpvDl0YcV9i2Ab6IFClK5GbMeGc63WWidnwMj4Wld7eBnK+kstRCntleGQMl
P/mP1RUa0VuoQQNWzI9UbXItyo0q99A/koLQb6fXbRFGpoPJu6/SHkpwpOJFZIk5
24tQlgX52fDUx0cp3K/4q9DBTsxbWqK6HDz5UmNHlUcHJ9h8lTkMSvdeUFP7xnuF
fWslzH5C3D92L6VAGzfB7zvAgxp71hMhoW5uJXmDSj5kNRyZOJ24xjK4ZwmyeJlM
HmfcMhW938l9VvI+mk/6DtVgigH/kOI5XZ7Cl1+RZaCEaNwwvBmxqYhzqmi/quiO
KzML7ZDyFigSmqQLwrrT6TLoMHOh+uOzOMyVcltcPFWJfQgDuw3CtvyLqiEgXCdK
VXcHu1L/NnkHH4qi/ApK0vrYbzOuW0BqaqNhqCxWLwHskYqAIarjMb1QcsDVMGuR
FvgMi0NSplYyMrElob108JXjA7k6p8N8r+rojn079FI0yr9o2bYP0SHg4KPAc2Dv
lv4y4an2YLqMWSOFvW4Xu9u3+s0QGXNPLEISum5goEYs1RbATNKvOkfx88nkNMIU
yspwBNnhHXGETq7laDaNT40wiLCgY6NDi8gs3aFwry0txK83lWguHiTO9BUOGmsh
Ed7uYngkV2kk6m2huKYUZn5py/kl+pHEnnOS/B+Sn2SkZlrU1yMcY7b0o4aBjlMd
EHOcCtEUFcXlRW0cHbe/TY26xAvnHHDGXcKMW9tvpQKFnS0su6TYagV3DuysFZ0V
e/pG+hk0fPUW/lnmV8xsnJEOIESRVRAapEBfZX6x1mR/20/HhhkJpP2sCqBIMcly
tKCdwiI4sSpkVf0bmYjRdaT9SsnMHwrIJqBWMVtBoAavNqFir/6v76oU2RogWDiL
is7Wo3IRb11nJkBl7J9VqUPE6UOSsIrs5SoNbSGUUj8rTYPbMmvaffhEOGVbruiS
9IVdT02uYY3H84CKVVr8MhIS0byTvRyoylB5nTvABFA0BWeORy045zmFrh9ut6om
SN7NUviADtS15N3ZtKBuxPbAr2Wxx22Q5PsOPsexbJ+nZQxImDwGUzSyZcvpT1Qv
hHT4JF2A9JokiCdDFkcYY21piEl+DWHP9sDA12EPabzwzXCV7mc3FokWNuXWurvY
4xH3/xG8jmqUoJrJVYjYmqzcmcS9uQx1WUPhQZ2Y9mILe+AHviNMI1uTCGPvn8T0
jDoGd2BQvcnuso24ue7kpxsDT5izXQeC+X1fZyKQ2qvN2UMrj9Pj2KpytvNvzfMF
DgOEj374ugDCiWIvnRiK/r1psQUrOGc7aYBwdLOHoWwLrA4zWimwqaqayHKsB370
HHYROe/DAPakZmMKtHL5hlNhJkaN7B0iELNTQqv/dcamid5TIwyBnCeWTBdSUuvM
K5dYBPBeHVJGoSK2wjqlGzYn8kTfBBqlzU8Aj0dy3LwI/kuQBPnedNEI4CiR3a1Z
fqqtjQ98Zx7o64cu5gcD3HAq7vFJ+4HOPYaDGC62tbZZy8EkXRU359AoXFuRO1Yb
xaSOFeh9IJ2ddB6FBeVxvRuotjEB8lBVZj+d0zSnU8CxhyXRDd2UEvoheZWaQ93H
TPtG3beavHGMmsWae9RKPzTKjeV1KhyWtarCNnOZaYvvSMNgdaiXqs11SMYm/R5G
3vKfES0LdrmCsGmJMiVT13jjtVEGk1m2wm7fQU4tCQ8cjMt5BRjY9qkOaAb7oZUl
fOlE+ELd8saHWqpl8EOcyA==
//pragma protect end_data_block
//pragma protect digest_block
AAsNobfEWUV+8a3nmTOWNNUSNjE=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
f7nTk4rMeFhrD7JtKzMe4KupEDutjRGeYt9iWHNX5lYb0ElOMdCsUQg4ounFK5UO
vXBVjorxhKkq+C51ULFtEfUV35ltZbKIiJIQ+E8LTxRP/bMsMYvIR17SSMXV5jUO
UhoL29YEqcIi4oC0+jqgk5pml9GGi9OD8f/zpplru/ADkfrn49YRRQ==
//pragma protect end_key_block
//pragma protect digest_block
YC/dI5i5NWxwrfSs/gw0AqAOK+U=
//pragma protect end_digest_block
//pragma protect data_block
TRquY+goJJa9pTpRoefFM6ZO3vlp41AbYh5Fs5M9UeqPfsRFyDSlerednLRHGuCt
ESVR230B0I4t1Cu9iufeQSxAMkfFY5+Er2qExBGy5ii9TD2U8z0MdJbvXGJcwpH9
7ofezJGXn3A8D5Bzpfeeg/WKOhFM+WUSz9EtGvfxHp8yUJklken41RdO0euqDWDK
N9LSrgwH3iIqv7qLSV8y4q+DL3IDWkurUybGadsU/MsA9cMf2aZmKRVpbAmQBND/
uiQesVNKLvNu6UcUz/n/jrpHwOhFU6bFb7OVg6PwukthJ0tCmu/gGIhITYVH1tBh
Mri1Q1Z0XRmDqFV1ghhcofdcW0ZSdhFAdrr8urFOYplAMefF2dOKwiaNuMr0pZ9O
NC5nCRPDJdMEpPHBifio1gwaW93SBFzY+5pS9KiLsI0=
//pragma protect end_data_block
//pragma protect digest_block
wnzhr4HL9fNAvEjD6zG0bIJVjUM=
//pragma protect end_digest_block
//pragma protect end_protected
      //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
j4VJkDfbAO4xgO3N8JxuKsxSqQFsIWAo7g2woSHeGivA0y94k8S8oqcF8WuS+Bde
kEnTe+HwNMGIuFYuDihqMWY+8LINbG/ZIyDcx3Tp6hxiuA93RVDmICpDjiUEAAU2
nlFMq2jG1wIVXwpRBFgnd5MUXZRdqF3iiqXHTuqCPr9k6LRIOtD5Dw==
//pragma protect end_key_block
//pragma protect digest_block
KaVKdCyXUOtziX84ai/otKGyZTc=
//pragma protect end_digest_block
//pragma protect data_block
vLYH5ISJV7av6dZ3dj9SU3AlTFQ/n+gbV82hNwyEJTEqpYHfcpV8YZIjd3aV9Ebe
zv61bOPRNyaHtpMGFwx048UguuXGLq1fMUGY+VC3yAt+LnvsmAVN8eNkKGC21WhY
SywfJ5QrqqBwH2Klzc+k1aU4adImX7C2u6Od7yEdzZqVtuknHD+YRffO4WiLnpje
jSFBQ6JFjec3tenqUWqL4IKCI5jzJFu+PU4FbESHcl+bW7KuWXgdsDro2dacwh+w
TDQVTLB2QRlNkrotIw8/6ySVUeCId8tk7mJ8tNJ89E2VqiTwBPqDocTqQswvT7gx
cHZ1+W0iBj5XVpj85h1ftbA4LLeyKQ60kknf3XywSXsYowdCut6TRzudASpdQnml
kyTsUdpl72kvfTpQ2Ifpb73R3Mt/lkqo3ZLNwlotCu0S1KVJfWxSrF80ZLYG7D/C
AEPmES2lFo1gyIdJzDhuuxJeKecix20WUoOyq6F4htCOMpYFmgSOunhT+RSJKem8
XP7yYYQ6HVCzcYqRQ0rm612YuBYdH0PuchJCfWgWy6NEPjg/ko1aNuetmqULhXc6
IKql8KfA4F8/bunotwhSJ6Jtmtkuucgl5O4ZX+z0sK84jH/R8CcgH+kv6XRwnHyL
x6nAFpPJKsOFEYon3Q5zyUC907tI25n+9aHvi9s0pPrtGcIeyqYuUBaYRESTez5h
5dhIb7ZEzFHFSaWWY+HZPySRvTEHTu/OuJEVTFaXqgtnB9xGsB3IaEmXFCK3tvuF
ZLVP1ia+PDcTbm6I+u3KHoOwtrsnxsTNFLkNm0KZRRpoIQCtwh749APbTun28x0/
VskeW2ibP+DzkJcV6Pdof425Crb/4cqMbHiJ38bIpFxGn0XbLXM62dWeP1wSj7rK
jQF8TxDRwcRbnMUTWtfF6sX35MenEWfpweU3kBGWvzsXdvYKtk0ZGrtLt6LUDWG1
N43HPeSF5v/yj7WLDobDAiZWesHB5P2V1/PvXJrF5gr8JQ+E5uiWkRCDSP6pgeuo
zSQVxRRdGh+RVdxJe5fbJ9s2cdx7QL2IMaOX30pQx7Q06eDobI1s5Ekg4bn9bLG0
Q/PApmUMU0jYYtga7/Ov61mBuafciYGqBrgJsHrDZXXreFdx7F4B0/+xXj6WqjGk
cmUeIMLWap0U3fv198unw68pOeSHdrSV3/vsRytNrctqhMroxZ2b8/wSuNfxKFbR
0/T3TVmmbDAZwGD3aZYWIcMU8TYoQQCn+TKkhDuDeEMxqMv6NwVVFGJI1xDybja0
s/ft8o1QShkBcUUCY7sZBz6ZpR4kxyHPlL6GX7O/GKfAMyKa+rLxtQ5HhfD/Jsom
EIQ+Nf1HtuE8MoIQ5nQGLaQPM1NCdp2eM4ZAMDdgKEF8Mgxd+WUcFfez6JpoDls9
BFUw+NI97CNgGvNRIwpFbRrsZ52wL9Tmb+O/X61+duWGX2H63JqCjnDg2Rfda9RE
YGsXDD+Q2DuElAj7a4c438d4RJbAFgBu79TXK9/6V5McjZhNt9SSq3/XBfPCEUOl
X+9ejgtbK0IPKbfjfmFy1dapTxhu61CuKae6gUora5UbCQyAh+9kdgPSYvQaNiJC
dPAPacvddh9YgjDfNkSW29uU6kks1Ht6QxUiE94lMTw/RPwtf5Ec0nEeIl0RG3Bq
ZwzUNyezblSKaB9Vqc5K+dCg12AytWI/EZOLdIdUQJ4vEdo4Xx6VfTTBVJMyN/Hj
c6iUHHRsIH88FoAxA0O+UFJy5AtFmBOryzAIpISAru9GloL20jvZiaMUJMX8e8Zz
hv/YgevRfx3U0KPgauHpJ0GUxRY+8TQdNskl9tB0foelyf+Nni6motCaPkpgiiHd
bIURp2jntxDFnRi8JozsRwJS2+aG6Q1Iium5LcTfavXrFq7vgYfEC6vu9jiVy9PG
CH8L2RhibXiP7EkCTsTcsxARargMIIAZFMcXEkNpGQjVpb+5CgiF+qM49wT0wZWv
5dsZu23pDPBNLokOhcIvB8nliiOelnNXnywD1CxE1E8sNrr/h0c95hYjMKLlFN5S
CXYM9S/2Tia6a2E0pVjLpSQA2vK/kxAeZXG5RuZ+r/Dx8177FHSmMPuqn3tomKmy
5xrvBKJe7+YOGDdbk1PcS4S6qnKvzt8lE/y8B6/omz7KTzViYzQZ8n7ufyY+Chtm
UaTfuSGnocIWLdlgOBKYouvQo77u/JeHZWBBKb4Bg9xOulfzG9YEyhufoJPjs9K2
hiH81Uis58Nz7sIFWKYXlFNz4wg5VmfddNJTRo1YqPAyRxHElG4/O9d8Fj9+FHeH
6v+fB+vA2WPwr5WMh89CLRVt9eH4IfObKYThNfJcMcW4AL+EvkHO7hFAopFMYEvj
gkHFDgg0IRR5Sg7ckv+KdJcQTEo1tRgCASa72nDzw2aHDoT/rS06DpSnqRXtepcA
r1/6gmMo4bMR7La6EsVu4zGDBY3+MnHPDbemTyYHHWJ83Lcm6XPf6+SxgpV2X9oF
DtV29dvj1MziGtjT+o1eHVj8PVTH+Wy0IeeafL4QV0EQsvRV9XeLzXuPcSpuG1PT
5TMSQPmgbQA3b6rZwqp9Mx7MWpBvFfnuns5XRc9GDI2iY5QqohkeYtEbFP1an5Nl
vl+Aj+BuCCxQujzVdtoC5ViyI1F9tAumFZepe8F83s89c/b786Wq4hqecF302b8J
TjEmIcWFdj+MnFYaRb+KwFhYUlq3fFaRVgoE95+i2vKp9DRRUKvV1VwCkjEM+Wud
1/2ACDMcNIjnEhH/BfPF6WfVjjrFY4JG9jNiOFXjhUYyj//0ljSSBcCaJ4nRpdnE
rBQWBdErgyT/foYlRALzN9xshvukqqmDb6Jb/Zp/ulKJqACdBoKGpgezbgF0M4rZ
nJRNM6k8cSRn8N3Ja1Ih3lRLvnQeNOwxyR8RXTyctQPOcIHxE77n5OqmAf8h7cGW
MK/Dfz2uoBe3uPRNFMFGchIYuIuLbaVuJeba18TL0UIzONFK0hPpBAiBxqJxJIvh
WFaWFrTKfDjlDQScG/xbU7JJ81OSXNGDs6zF1fv5UEZtXBNZunP3T0vXu0Dj+KBC
03ScYuJbc+/LLRc6CimcYyMI1c2ymEKm7vshHH5Yqdc8LY5ejnvY6TBtRbsnGAO+
VNUigZaZMoyVFsnH4ixz4JO3LgdLs1n4XVP3bgM4GZIpDiMB8a2hdRndOoG/VENz
sc4WEnLRkG8Z4+5c8mPHlQE73t1fuOLVaD9e5qTw+MuDK2vmDuBYhPjlxGu+wgEE
SIWAHx2usVWBqwbnNsourtHwfXxYeUcd3zz/a+U7XIaiHKWdHMSSzgfTEpvFL27U
hpFZteU/2ULkzgYjC1PmEGe3ryDVdirkP1/rC45CfA+z2p4khTsf/7pvnetjoeFu
O7XUUzv7yaEIOXxiYg7avZJTbom6mIK4i1QKWpeh3yZHPtLmCof1OixIQ+GXE/Pe
xHxxoKhpYOqHuPkhkTMhe6WyCrQG6bGm6pOtRcrFljmJB7ma5X3hkk2VLCiNVpD4
J+2u13VctoutVviKarVPh5VzvRFtZbg9AsTzjnIIJt+XLjU2oMkl6wcew95NwTiT
MFavute3sxajZoJ1ernbUmyux2VbiMQVH5b66AcKp3C22bEmb5Co/HsO5hSVubj6
94uU6knJhFvJ3yi1cC6skDsyGlBZ3c/cZ+z3q3lwM4H1IcaZ70BtspeKeHirI5Q4
CFw4lzXNFWRj3ODZYdid6955LzIIl/2uJk0T7tZAW2ztY1vfd6Q0TPBUykJyX48+
3qVnvC8tUk9abwrsp2A45CwK7pN7kAixq4wjfTJDPCbxkAF3PZKEQakW+5y46iPT
Yea0Kh9fBS2gNV62liSXcCObO2Qd/CFqzBF4CI89oXoQkkPcmj1EnKDZNx7XkHOd
js3qdFspINZJrpiGbYZsDc9I6U7FgQYHqEh9vMx0OWNR5R/GRcqmppvonve/Qxa0
snLjQtqiABWnKFHxg+Slg0/cowY5oaeMD1+/IxPvzdPnPqMXnCntb41AOYnJE1VR
Rnbqipf32yKcwyzmgmjz6Nn4rPvhpiwuYLNG07XPt3cmCNQO+SzARRFdJEQAiiD3
zY1TVwwIDzXIoMj4yUSLrnFCHDhxoMpTtK0BAlMAlxziRlzyC8hKkkXiRr+tMMiH
2CTxpgpw+5U5x1jP/N/gjmdgkX4ZJOdztyReNxvj+g6r+68pS3KebOhz2Z9nHUZo
HnjXwe9nFsptSUwvvPTLnuGb3XnSy5SmyUBwi908eQsItl8caUXfMgWmkhpdVSBh
rCmQ4jGbqXETiJPJVPCvDkDK0bC7rIJmYj21d/mizDgYJ+E8KY3MO0M5BH/fvtuG
4NKja9+1G5DWRgTaJ7ZWdwgTtxh+5S1bMKSmuvDeP3sOSUxnkUsqa9jwU5ZeXM2B
Bl5Rl6ncCqoqP8NdraPF3cq5bysmewoBJHgpr4a63tmRLFSLCFXk+aOLma+cbAfN
mYjf1NZwtiGLdgkx05CSaDz4J306sQeOqjyPIUFFVIjh/XMmEHb8EZpVikxA9cT2
hMKtzxdBVZTm4nP1ccE4U7gs+B0pHrR5QPgSxD9TzMUSawohQeHLXB0ZE8aGNuEp
kVVWX7peNp/o9awIla/jU56geFLS9s6CHNZ4KHm66FM5Oo37AtZuUci0qExgJMr0
80nLISQeCLeBDBl0vEoJZPCLfPJcJ4doKLg/c+2/+3zGGAyQxq07qEF2zsgPtmcl
aKIj1J7NLUFzYSahGgeJ79oib8gj4++RMcd7F3cXtssV66z4//cLPiTR/TINBkOe
34/I51251pqh6vzcA2KLdvyYAS2IKEUEyOyCZvqOM5gtKegDv/5+UDr71gmKcpa5
DzrGRyLRmSawZfjRB2XvHWr7Z9ONTmSHchFHpkYeOl3QdUEQ11SVRwBqdAlp19kW
VDB3V5sSyS12FgmAGyVARVIV47N1Xa1XbP5WUlIB/xfL32kABhDveWSlRH9kH/R4
C7MYHXOdxACe8Owq0C4ztp34aeaf8Hjoq8v+ZcSAamxbYc0z3eFoKx1T/fqXGRjn
vQ3crylqrecgnjBLyg4/aKOJmcghbFDRqHD448mbrTGoc1UanH2bEM5fx25du1H7
nhZSVuAwPnFph2at5XdT8tHlB3PRSWUXe6Ryuiamno0DIPbX7FjJuXLVMH1gzuQI
fQLgLa2CUmMdHuQxsbJmj5CtzApmnmIQerMZKx86o+0JYzWzWmEEiIaTiO6BZUh+
zfhuQaJWxuYLJlPlYpGusJ9MW36quVX651jgsu4tB/uRgpXiDhYtoVo1juqAYQVI
y/YLPLOHMwLIvM1etbKSMP41lfi+hwctejVmz+Snh4qFzbPIc4ijb2eOVJaoKx+H
JaIzj2mHfE14VCVfyjOtWnnIMTP+CMLcBdHiQgJr9c2WZ2FZnvtfiybIDr3i/Gs2
6oKdRlJn9ZaTqHFLqpF95mQyEGTYEfAhFOiPXagvhLl96/4sfIY/NUs9ZlQyWM6+
ZIIIm1sJqY8bw3gsukU5n8aHeu+AhQ6CqwI+qSP6ECLjaVxm7i21HlQKylc7WC6X
ONu2rzvZrVC6W/N4iKYeIX7aVuG/UyUmvMAGPzDtIeQlwxLkSXTH+fN54Tg2Gqqq
LG9PetnvSWw3c/EyZZe8TNfiB7CrIoqVM/+VpFLdBoc0gxjKCxvrXPqu9yKm46nP
926b/ojV4UytVN66DG8lAgJw6xKGE09IV/faAh6JYk7FzBMhFyulJixbY0Ev9dLT
D5dKgx5pjUjRzm3jW2DA0f9KiMkgi7iJtpOOqzj6zc3WSFJDWcUDkSE9YHDYJ0+o
hLPNvvSIqxKEtLt1gJNruYMTtY7vw7HEhPr1pFIFRmshehFAfUJP/CwjVtXKyv1p
1m7K+gq4KWMk20J+iPkgEPUFQYnaOmS35Rjyeuy5x/N60A9TVMEK+/ykxqFIU2Pn
2zuOaHpi9kCfYWRRgslOsWJp4aH6/bMF2ZhG3kUR1vRFSIQ7as0EQ0OGFoduogab
LVTZlivZC1QYSZFNFN/kSulda26g+zUa0nhlFMb35WgHCZr26DW2oQtEcUrCKLj+
kw7aS36vcJm+WHi1QxAi7G74byU6TYqqWT2T//oZeNoBhqGr2WnEN3YQJb5fvhkI
ytPvi4cMIlaSo12YT1ggjXV3c78SyXAxt+Rd/j0ZXAAU5GhUTwuuJZRPZMiAdAuo
JOAahpzxcNZDBp0xjfGLs11MfBKnfJCQZ0XwAa4McRyH8ZNmKxIokXxaaVo4UFe3
9id4XM63OBbLvoXRZKivom/31eI1sWvQSJoFFKWENIbfJRuNBx3jE2DSQGWDwN8D
AuV2YfCnF7vRRCbyyRaebwkIHm+4teM9TZXejA+i7j7i9oVX5khlRepmsatO6WHM
Mn6lVk2a5lLZrjg7ricRxkjCqoRuz9P+pLgLy8jyIZphzHYDBR8tUMYRCbdDpiOS
2MrBgR73XrwJRTtEwGKQ3XvgxEi8noPuLCW0uBRchmaJqrrQQtkzbxORN8HEe+LI
3xLaSUAPBUspmTHm5qDkumJbiH/0zyQvsZijHLk/cOpSp3eoha1QEqATyhnU83TQ
A16yLajntj/RM3ryPf0ENT+kNF3+wFlHQUe5KWqzPOXHHwSiHv8kJKHb7+j88mvo
UHb99hRpWbJZa/A7KdcqtzzgzJnvV5S/dFG7NVQNV44RJkLdXnIK6s0T0MH0jY4m
ApcytEJlcvZUmczYwDdBcpKQlXMtWJtOXBkLBP6gfp+1Np2cSo34D/ue0AQAT8PT
QNbNt9e0SjnkVmrhI4ziwVPGV8lCNxMkM3DPTcAG8U6+ti8AbHe49YkIrgV1k776
T17O+Qk/fbzu47yxerNhE7po+K1O5+l9EOagYFFtau7F2xdXerM41wFy7Bk1Fep3
U3f4veDooGTfI+2+2T0uWrlEn3U6Lq35RUirBroGKhEwBoRqkCrflSaENkyCb8W7
TWMx3JuFT8UzP3nvvtcIftuhCJPx20JjGBp5UjWxssEif8O3+fI8LNYFTqgybDy0
dCqfCcTpD6pubRdW9kd5daVhwJEaR2B0GVCw7wZy3k63HaqoiGG4946RWhPYB3i7
fthWNd8BtN8SSHPSok/NFoCfquSReQNJnUZGFGLlAhibspn3nMJ7JBo9NR1CmqyR
EaRnb/OUoz2nbcmrHZbeh0uUmCDnIRB3xyJLUXrIfd4vrnaSHmDr+Ahyfb96QZBX
sQCeH8DiVJ6swKRsb9+CnqPd0lsaFG+pbCA8n2SgfKxF1KtuMYX+VA0qh3OJ93Em
TcmkhMpIt7YnnF3SaEFCvx1CzigFx+Yuh5uu7WQkT8Mi3SWf4+7btuIy9b+cJDlb
QKL6bs8fc81F29XHgYUib/EH2UDpeLhLSf4nBu8W4AkeXJa+7m+5h/cp0c2v43Jk
sa23p484+JU+aEs1W2Z1qwXfCcKV2CLUOqascUZG0hehrfyy0scB3NMEoj2Xr6yw
x47P820A3ZlUCfk2xO5m668Q9pX9Wz1x4Rj6j6eodoF0pecRuKmvNdywZLzdQLD6
Rk9on4K25Kd0wEPJG/5kMOyEcWzvtDSTJ+yQ8B16i9usnv9z9Fppz4iYfG2b5okm
gtCnNBh7yimX90hTk4EY4E/btCDmwYFdrZqSpHV0s8bnTKdZoQDQdKLoSspiLTbZ
cQzyM7nEuzJrePhNPaHWN76ZT+fW9VcLlBYZ3PD96MBMqPZ3rCVYP1+d9m6OnlVu
97yaX/IXEl/c/VtZ/u+dHidaCfhPYqOkqMCv9Pn47c+QuMn1D+h4baPB9j9Mag+E
trp4At9XekIR6qETpBzEPIgKrSOY07oji06PkMEYZKv/C996ZvGb0iZrrWIWxmcw
PGo+0ewf8WX2D0L969WP2R6+q8ZuG1mSnAUACXrmlv0nwV+SGv2qVbec8mHpO9gv
GgpKlZ31RwMGAheyfTe3EcpH1JLqDzVS6Y5eeNteSK3sv7Z3ANBlHDJ9IwT3rMKz
oBY3Kp9XlDggvAjypR+wMRUEW2AOYquOoExOc+0uIDgvcIcw8/3k+5VPqpIdr5iz
KnAw+4jbh2tbkaiDzDX7edYA4YdL57BHFqOX5WO+3Qt9DDGpH4viwfjDvnbUn+lH
UsBnKSSs3+O18AuLhWAvce0liNiO3YFVuYgypiGaW5mWs1nC0zAFzuhTwgxkdUqn
npz7X7y9kyf96jD1uReun6r/tC451YORMpyczE+1zrv8NW4pjBp50XPa/4KaY5pP
UQDu/q4axx27mZ2kNm+TRjMxzGalqAKOxnFlor7YTp62Z6AdGqd1U9gCjb1okmQR
5f2MfvrXiz2UOGWcW+6Vwk9N49skAxg9XzwixbSEkh+iKN0dKuhiEq0gOvzUw7jM
4EGidAwOck5Yq+dntHa/4+r0nvZoJqz1v2SEZvuVfAioSNWo8rABVVIDmS72ZDze
nCBSOcsfv1B8g1dy+YSrsbdCkabuPcYSCDZcsWTu6ixbUDaym0D+cRQnKwQBSLXO
30I2d4I/Zv/RqwpchcMr06n2kUc0E5r9mOGUkmESlCN9VA91V20/2dHWxPl8fUH2
aTo3zVKkehxWh6aFoxowO/u9W4cQrSBw69SaxA+8tM/SQq98XvXqlDmiglprzhFQ
BzBs3TNKHZjVQGnQkwugRd7utcCzq9Ce82gKABo/QVVYTPX6sGo+fMxWQMR5MuL1
0DKl/pNeR6P9wR4LLSwKKcQGoEQtnFRtSqNhjt6AxjeJt7BupYnVGJ1cT8Ytg7PT
2PFOUFmy5Z/AGTZX0oh77FHF07TyMpVvISImFglhsVHrR8yYZM/1Q/XnAiyg5L5l
fqqh8Dk+r9gtAQ3FBVfoDqmzDJ7kZPbS7FTVtCfeYvu0PHx9JxiaxbYnCI9BKRi8
eYXLF5YpiJcbfzY6iJfcQ8Wyxn16EnEYeiyd1H6Jxf90FeEhQzDa7/Kz2yJufpSZ
SsgmKAfNCFxO6hcYsLdgTVis1x+KeJyhWPoIjEO7KDEpdHVI32MQSGG/zyYVVhN9
EqlFKJQ1b+hXfcYov3ET9Vc7oW8lu+Qa9WUgMRmOOhYmqdL39uHs/CX10BHyHtNW
d/SktC1+rfXoKL6KJ4Hdm/cXIZKsW5QWY50K6eu79B6TiwbmUGuomX1I19CRavvf
qBuDA4dRMG0IlZL7lwj9EZaURNL5EHDtm1q/MSDZLsfs4AMimAeMmkoPLZjCXS4R
68/geUoeJG05y96HqVdBs89Ws/kEyJroDK3kf5E7PURguMawg57xjo8rzdui1rsC
OMnCNDErbuo/GXFjNstdR7OXeh9STtlT9TaqWkGCaaE3kWV+EDwpBr2gqBvfcq3v
J8NII51nvB2R3FoD7EmXBR4P4Q67NmE4F6UVVUp1fjgM/VJEo5pOVWZuYY7HPwC/
zTi6+zjPs4Jk9WJmLdeTRLub5C5HyJeMvGJzYeivWLIOMH93iXv2UMyRUrL/hgT7
tKNsSsFc1ejuWXC3WqwDeb1SKZ00sRFAqI21NHbBI1JNqxRMoZlbJxmSU7QffP5t
pjItKDjxS7Ad0g5ySpyndMZPPF1vlug77ftCeZzvgZK4uZtnc+NzuUEEXjt0dVDf
+yWv6sQqTZm+qe1C+Z57SLN0Q9AnSQa9/wTesjS3BRjLm4bmNaDhH4JdK21gYJAg
r9Ee8jaqyyPnaNZxN/BylqATQbKCpS4zwt17VvvJ0bovevN2b+LBHZSyr9uaKd5b
hw1je/Tyl5jJENaR32Q4ed8TFKctgF2fr3G6AmV+h7yFVa6fpD4ZH6a4yO6Ncscu
1MgbWJ2sDNgwxI1stli6BmjtemsI4Q9pJSJ87Ni0wzKOGkLsVPohPxK0DV+87KDg
u9b+5VRJjgasg9pJfKUT00HZV1kXldRojeU2/1E4+VZyaWzSz7D5HeqeR3KZzFLD
IQwVpL/2pzxWM9LiJQNp3DdB6ru2YuzZTgTFue1fY9fyc8cV1Ab9nWiP+gOr2CVZ
ycSBFY/hf9Q2Q5UvPix4SJ+v2/0rMul6oib5Spthl4i8ujsHaGr/tOv016jYcimV
9nz4VE/DvJ1l0vg3hZpl8FRLQ0G2z/MgEBqZGw2slvc9E2/AwxH0Amy9tCELupFd
bHs+/3BnWdwSVCnE/lU/IyXf7B+Xn9gbAGqHKa+TQSUinhRqbswVLfdUIYeNuSE6
TInm27Z2IZUMFPNmeF+O3V1Aw2FJXOpNqj7QDgO2D2pnLwkpoLLCq/Oz0TMsE9GT
olbJ2PAAb5ZSLOz8Twk7HAHvW8+rBqbtW+dHIfB7phei+ZVZAfouK3B2zHQYc8my
sBXGfcy+a4iKLR+X5nXsbklFbLPu27ExxVXcs14/3bYP5XlnDyCKbOcgToTka5iG
L0pOOLHAA9ZoWG+TolqbFWNS7bZmIFYTzBiuauP/pezlgcX5Mg3oga5E7p54QwZD
q4TN5cO4KPj/Tlg5yAOiol2L+BX///7L8xif6xbtHAsvKFSR3BVaxHtUrXoHegzU
bRxbBO3UefdqpAPzIRT8oeKw5U0pinVNHUwAlZqWjvOsFoT1DRs8Vg4k7GA3j9DK
P2t6QepGyFCF8X5fzHOv3cB3mQA5fuVwbne08MIQ0iPEL8FqPkpihG/Spu6zWPg6
jGjAaLM5IyCHum0PCLRTPiBa/OteeIFE9i/8O5D6hIaHmxfjoOUX0+dDW53kSrnH
YBUVFcgwPaj49+mGKMgBB7PmzkO3JCyFBAMbH3K1o9Sm29tCwU98IQZ/9yRK3jEe
av8iZVK0WJzAklY4KOu93TngHltvqRo+KWmbVZL7Ymc/EzQZVCqcPwQAQXrlBQYV
qpiIWReeGQtoP5oR9fNxOojRyxkf5LkoRcBDoXkVaDRm0sjq5Fz5tCO5qOe+TufX
Hkr9MsdgHWMX8JQiVjwEe7fkyM5zJvEb6Wy8oZAeOjIYNN4ndvgFrg4D1OBNd2mm
sgCVtv1aaZ8W5HYFEgXcZbX2We59BEPSOgeRDOL+g8mIbWBzWmdtC+M16vhAJdq/
1aK1baqGBkpbntF6PyBEk+rb7ekwTYQszsCChuR4QfecXnm4zZwIbuyLsw7PE0Gz
WL3/Jh3WZIwfMgMDuLW3dFkEY1jjYjUDV7XKh4fJ6oYWKSIXeXxAH8hC1n2fpfIh
w9UkSYeS7jF+7KceCoqjIBZ0SoomR7daf8cw3V4c8LuTKEdeC/+QBQdIYmBmhfHs
OUJZ5Z7L0rqeJMRdsKsBXcBm62uqZVTUTr2xxGuBN2Jsv2VDg5Hu3AjwoxLoP+qz
kLUBJjUFSTeX14T6ZkD6QYpvcdeoXAa29CzlreOBv/W9/RK61N8ZfVMm9HQISn+4
AQtQr/H0FXVvuRaPm5im07C6wm2y3WstsiKWd7cqlcp02u+cc4srwkQVLHg4wfQx
bnnG19m5m8LwlR2gBWUESz9oBHwS8dffjlQr4zoMQ0YiLtMGDNi5SDF4S+Qd2/2S
Og1PzZe2wV8rocT6hk601bgBqs3yQVGewhJp0zQB5Yo4Sjoh4T0v1D/z91ETG7Kh
UV1GQgSb09Tvq40t082dZqR3AGLxha99B/JHtm49UyrDJHyJ84qX83Qyz7KJy7g5
v4i6/2NLWpbNQzxmVEDtfhLuNr8B2nLxChDkH7DnNV8aWW7X26fXkKhUHhe1mB9Z
/d+nddNSoyt6n4uUd9z7JUCsRxjTA/y9smGCj/wwLQftdVtfcI0CH0NATtObl/oY
fgkAJD4YwctcMVEWnnZwOPA0Azfk2cawum5gQ0Z97049Mm6C031HUv9cSRjyjKGl
5MXanU8nuv457vBiLWND8d033I4Ba9CV0zIscZq6VToaGTPP/Rg73knknpv6VEAy
yVs7eCpQK91hGYXy1CXoEu7OEPwzISvWjDzRBWZn3KGtLpKobr5b0/WEdb1lVmVz
Ajq9to5LqnZXxHxtR/4isdH2NKGZ3diE2QxWIJcsPbpnd7a/dhJgiOI+PPcvoCqf
mzVLlylHS4pozZsepIAXOeB+nIYNB+wXdzsT6tULJTh4bTnxRmzJgAT9Yv+JOsJ4
giWd4r33zhNS3QlT6yWvHNIhVI2RjeHAD6QAO4o9Jh07x6pljxfG2frrqTFJ4GNJ
mWpdkklagIlTQHieFhvBTLm8+czAdaK8IydBPPQjjESvLmd9eVONV/cshLr/igoE
Vd3LRWtorIP7emiBp5SrRxkHNNLq6Hp6iFOESoVU1pE3a0OHRBoxPrIBEuQTgdMS
6yGdJZZUas9nynwrJeWjbzDw47liUzaPHg5nthZfXNsGGByF1kK+4VbZOIOhQ57A
2l0/BdidG+OUVD3zYOzMmT2klCk7S7q1RkW6cH7KSeOf1BZCW/7zUbz4j7V9DaAN
D0XmBIvVs69fVSZNBF9Ck7cztc/BguzwiXJtN5pqAhrsSSuU0qmanD0LY/qNdwKH
ow2M/wkkaLyApqhyFq9RuJoQ+EO2QzzEgiSQQ6+Nm5fs31QTCyfjRvKhHyy2g6Ql
I6aekwGBGber5f3YYcTH5HICYBcRJk4WK9cpFCbPiJFhVx1hlegBOWuusPsbSe9J
bJxm4ywnacq+cBPzcdMtHJB/ctODUQ9yJrDGCzhi50HEOPnb60cnFPYDYsQxMb0M
r1s/kcaxzvT9NRkWuOvd49/psxiQedpROgfpEoptZ+rTOs177z0nlpISW1vlAMCj
TM93mbpPjpC4Fnd5yvwg3+yF7rW3nkhw519TcDQRRsYyUFkMp6HxzAqoW7iPj470
IqAAX3QAZdt9cALkqmAuIsZ71tN4U3KqjSAJzm0OGhtI8t4GjFUtmCFIkEvEffUz
0/a79HgJv6tWUW2sXmA7fL5KlxZY9jC90z9MODcmHly/Y443wRo2p1krY8ABw1KO
3DoTwU/BwBbUJh/Wvs8WwYEZTYabkat81cbQ/nY2bV7WF6wHmu6rb+xA7iClVQPW
flFef4e7J61KvknRmWQMoEM6k6ocu6tF5HbbzQSs6j1aRY4mhHAzfR2+uJtOzvsG
8+tiHPV9hVj0JwGWZ1nLF3txn8s00Q1DTqZwZBeA13grcd+Z51ltDroBzakDMAAF
oOMR68hHfHBvKR8gTtoCdoTo6cNteubJzv4BEHLJWT/IPYy1yUNxTpqT8iGnNj0Z
6M5hmbHxPC65rlJTirwojM8IoG9/7UGkbdgZeXXelNvodcSE2Q4CUf6QNSh5jqNf
ij5mGSBesd55yhd4SHG2A5pLYW+fbu/iv47RtLeCNyEHB855CaFhFyRIEkfBetaw
Daiumaxy2jBnKRJSHb9sfMKyUAM44KKSg5IVwag8yKtOyK79Cc75fTI/661YQWl7
FIxGHrtWI49yGkVU1ZxH90qDaU3FnAo2nEui5mukAJovqw4MDCnUmgAfNeLuZ1mP
LyFtK755YUJV9+b8zJJ4Nj5+4yJySEF/U0F3WkthSrNMkBxEgdRi4H+qsHkPlulY
SCityGaymrDdpfNLCvjyXYIpV5+fRjxtVD/B3SA9Yii4TYrFA+UbIdiGm65olewV
POTyUj4mN71NLey3FG4eEKWKOFi6860oh45UpxG/pbAWH+3mcMJ20SQr9x3nKwuN
MtpI04n1rl+4D24F6hOJKutMm42O5bJrBOrmjRIK+HTiWkNIVfIdkom3Gy9+RC81
dvU70d8T9ZLgl8yEbqgRIQptNjUSkFNuLXF4waX7gyhoX3JNFwPCrY7+fZjzrUqS
w90Za1MiMCDhKPIw/I0n1YxNsPNPAV22J/sT/mLqNfFdhjBPaImA4D3LVfm6QnJf
Pv6eMFeDpdQOz9b4c60apbM1eX2rxm7yASvHlRq7nA/KXzuBJzsPnJUEAMaxjNgx
+cGt+ZFZTqfHMuPDn/QzO4vsDkRMr62I2VspXjLOf7t0dtm2davvvk4pv/CLLduI
cQKXcPlGoX2ulT/vxtt4FUwJYlPn50wnXkpywtxyZ3DbfHVPbyWeJB424cauKOYj
ui70uP4rg1r7Pje+O2fp+vI5t0ykHqbXcMYoN49c37EXo12/RCQvBfNzZ7JanDHh
n29cud0KYz7RDz1p9iBhv3DXD5PJXl5FJpVvaC27DiKXEzI3XpDc7w8Q5uqp1jG2
kYq4SNfb09kWfLNLSaReKMc+FAaNyNnAH9IoLFU4Q6d+4kisOrEVkBpRrv42sr7V
4X4BrQF9PntXvOGqpv/U1Wv5MA+wsvmUTcxMgD4xbsAje8C1hm2/Lb2K33yGoEqy
+aVFijkHwEBOq5Dv/3ZA1CFbthdpvu9QyLwNUKEKob1b/Rf3V5SK8OtMafQC2q5D
73+2SrjCZJI4ZnCaGf0o5miBVRHawXURcvsUgfQhn3ieLVKQK0AXjQbDIEGj5CXo
r6zdnV1gyddVnkUE2W6ngpw88NOYiV4LAwjtG5lE1B6nHCouiidaAKXdSfXeAv1J
5vMuyibVLAuqAuB+pZXTdPQLy+6mOGDM6iAMv7xFgt+iLEeP0mXg8N8L9HtDE+23
khh5IeFHb/Ardq6bThx1sLySNIfP9cwBWlvkjZGWMjTHMxO3xbIFDgi12Jmh+G2N
sX29VH+StQRqmSCYfG+1nA42gIZIRL9u9wj5Q9HdFu3aZMhPq/vNCu9TIn569kgO
saM2arDm0e3WheLksUjHxpwhaJAQmBgVQs12d0mWXk1WKQln3HcR8b2ZwdLlYcIh
B3LLCWQX0KftyYMoSz2BB0fpN3ISVokW2+GImEBibBPFJd1ihmd5D9Fx3m+SS+H1
zK7eW/q3WdnYT0ARQTF7YMXmXUgzu/fXxZ6PSFWSHwSGKiul5SoJiLMr4MZFiGG0
D0R5LnwxvxZ6dXYAtFD3aRJ7PMnTMmaKHvQn4xTaiPleNEVAn/LiCvHqy6TtBKug
U9OWsA2gdMrvPZh7CLJ0NHoZTyUbAa4TjkxsOQvTbWNzeacO4nAjJ0Zqs6RSrYgS
PzwaZvG82aN5ibmHGZrMVwjLuZXFhKMrFx46boLp6eVMzTeAgdUNOwRRSEt6zGPa
XtPYkIq3NuGuD+AyJaCX/1aDMhWNCaabXt8MXPH6YCdoIjV6u8Av58R+YEfpP0Hd
boEiQinODmxyfy8IyNdfBSez5J0tzI2DlMhpHvQIt417NkNTHtf0qaJ51ZpLfRoK
8QQaYZG6Dk/cSe5QJfpuAZJ2QtCDAt0Ksz8S6K2IqyRfPrg7RzfChcoRSzA8mWah
Sc14p8t/ewy41B5u6nppWcN+mYSWXXNlwg9Phtsuu5+nqtkJN9lGy846metaZiQo
Sri0W/gtu4C2hFdY3t5DGcc9H9AefT6soIJAI/hqvVEVruYcVRo8Egv0iDFnqRSa
2XMZysaVdwTvTK/jGx/gzfGDeGWQbHBf/hrCcuMJmlz6SR23+4nK6Gi/H3iBDKpi
yynTZJZf20tbXAb8a5Wr2baL8/x64ArA+WvRyh8+I0jer1ops1y7PKCwBDuk4NFR
3l9lp+GDLLzKogx3a4Oi6YURjfRwTLA/1NlYQCv9RiKRuorjdzFKhAR/kRTerdHn
ObdtVZTmKbaJO2fCMkmtjJMWtQjc0taFPHXOlNP4i7Qq5Ud+sRgupfRaLC+49s8Z
Jkf/c2x6axYTErwRD0g6l+r3iDirNr6rMzwjn1P0nvr5iHqWriFWmb33N8xCzVne
vf42ytXKRobqnWuynPnhz4VUB8Iqn+0TblZnmBMt/Do5HKHd0OvEgVphxAPHf0Jz
rzuthCLc1RA1gp0C+0RFrw5FSCJzkEIFIfubqH5HpsZ9GdxjBXzuMSFhJdxVvM2D
uWMZhDL/DJeie1YRsX1aXdwnel8aUNvqluEA5et2TlgVPBaC4+Hl4++nhRZfdRWe
uuw74rJIXWfS0PizMHWpVXRQ74EcqCq/qLk8EuW0NKyUkiylU9eLT4B+Frlnso2a
osc4by6aCd6mMpGrf99r0V4VOzw8P2TJ2Yr3bkKunxwibdX9pOpdjl2Lh6PtAEdG
XYjmv4mY/RIzN7gbTXo/3AYkYBFTdBwTvOvH2uQCZB6fUlNjwFV1XYeq8aIGSSdh
j4g1RAlUgbNecbEg9Rgfk8Of3Uqeen/+6VA9Bnk3jJFqOcX91fIdz84v+e3bOoRc
l5FQmpEG4wUAArHk2HkjAPG32qo00VrGeoPCuQ6KvGXk2OSnaz3Xowx/zxyMLO3G
n9zhquVuH+2pqv5fT3Yxy69dpNAkggFPFKLP0/xST1VeqgofVod4CeEBfFUWccsi
3ymoFhgqIEbpeoMgLnZWgTX1n28vBGWseT+TlBSuTg+dDmFz2kT5MCGxBZUDvBd5
FXHRREgrub7JbT+eKVeATljLOS6DJ0gYvzlNu0pzyRqdSoeo80HssoI4FCu2F2dY
UuhIOznTqOpog+jvTYA0lIwKxo7S/8MI8Cz23/Y/qWvERQYSvIb6658hImTxwv3K
XpYJLkHYSBDFkj1Bu4nBso3AIMAWuS3zV+Q6CaPJo5B0BRbc1wILgBrICJiqspa8
Giud9yXE+ktsYTrx/MLidQsF2i5QUQrKr+wJXlH5/PJO6j9Dvm4Me4taqVqX2gQM
w6yuP71QnL4DO03K2zzn6PQlgpFnp/r9GdIm3eGi01rU76rjHDr9iCuZNAA6haRs
vz8TQLwQ6YMrrasdLVO0p5YUppgDYuLdfeyUtvwmDRRX6z00xy3H+cJDV4mUv0eV
tR/C4OVQ9o0aDqWh6p7d5yic2HzQaKFOU2guUyABjpg5WMdK0k4ZinQBPSmnxs/M
Tr4cKh+W/ueDK0z08czezGJjyWzUTtA0gW80XUd8tRBQEXucozRxuRB4t9+N2+f8
8ly5reEOtSCNRocimijxP4bzx/2sS+q684pR9AOiiccZtNdnsFRRvPrzalVfbK9T
NBXBAKA1UAaHz1rqm7oa6ON061pDRjNJIoVJNgpPNRaBTCwXEa7ZzzayLqCweZGr
FsbX/wYy2mi4BQbWTXl8cRqmaXjJWDkXGWNPBMlzfS/YRJQJSGboclbm66+T+9Yz
5vFFjI4RLJSDkJdNhWACup2NeMejEAmvOL/pp2rqWPowTmPnAxBNYQIULxplQ6ce
PJ6XYq3Rh6RiTqxAM85OQIqWyxH945jJdGkVmFRaIZjputtPifpXYdJXTLgBFIr8
FlOL0KNUlIwJWgSyDO6jbdgf+XBsSavujxZ9oBZoP0kReezVt3jtW5KdeC6PTlRo
CnBoguyshi7H7KaFIxrK+DwHyrS0mzItxLPGshktC2BFT/TW1Evz/nbRTgL7IjMB
RU9cXCrKY2vw1TxJCj2inGnNPJqkVIQ/wDke5jGempEAEP0Hd+ZqqGq8tktJlp3+
ESZvo+B/qMMyVnoHKeEBSqNOIb4Wu5nwii7fQK/qRKIXr2/TJwvbJOvP1SrwORZq
Ny/x/kxyWCr8zAOc8cS2GSe/3B8F5xjf6H7Sn2q3G8zKK3z1SStp/nBAJjdGfcen
TR5sdaYy9O2U+1da6MbsTGHGvPzwZULSRJHSB0IcR7Y7Y2BvKzOnSvYYWcI8kUuS
pnrpOxzNO+9A7ZHLZA0xYnRGBVZDeMgKhXwm9Sp8ieGaH6ruJT7dZg6o87H8S+NF
4ERDoExCdgXIi749wyXFv7EMDYQwcqd/J5SGsEZKWpuoD+oDFlbqXX/LmXuTOhM3
ANYhwwzXezvOC+bS517Og8F9Fz21Eey3LFCSeQbBij5hHAsffnl7qAnotSW3des3
Ms2EcXDqWafSoFr18tYqP4SZ8jCUFLplli8iB0tWJeEwiVZEoEzdn2Z/p/BwdZQH
P8BjatZ9SiYgirY6qEHCgrd2sxkIUjFomlK/hHnvu0URYw5V4vhH6KNCwh/Zu5DD
0LxrLbPa+QWJ9hhAoGui2+JXZ3zhZ6GgtP919k3Y6I6svLPMPQ7rXRSUw0CTYNYa
HF3KILHWLueIwf1DZTYfKCoNp08NmI7H/BpaFWvQYOz298aYAL/ZporSbLPmWYXS
YvIyaO7qqplUgsoasWAFqUjpI8QzXGqtfN/pKjkfa7GGSWwXlNx/w8LXbsszhPof
RE+hGiZTUTq7Y7h9N0CuI4PBTgr/yeUEO7Rvcy7bwGqXFVgWOzvzAFazdf2GEwXG
rPWEZ7OklbXZ17q4sJnH6P2l+Lr/L4O9SkNjCy3ILSNEWgq0Hond9lCsnbPTpb4K
htFYzNqhzWgcbRXqMihM+fjdNqvLX2U6YxSWkNNec31RdTzt1PAHk+jIVWJmOFfe
NiaxYHu+R0PBo07NM2lCcYUmexnl0gC0qzKyPgs6cynGXY+OlKHuxmS75ufIPyq4
x15gDFtmBpP6WNMLqAasIodpJioKwZHVTTGtsH76XgbhIkZ94jEXMj9fVP1FnPfa
g2AxHRTTdFvF4Y1Dv9moaBmsvHJOPl9AiBvmCUWTEl2fMnTNmEv48RyOkuTdqZHV
7BBh085J9HL3esysIR6aBuMK4z9fZBsPnuyRD0XVza1+bAFEFz4LinOh974x08yq
YiImYsx2iWjjGM5Gtgn6UyV6creSQCw5YM+DMBIjQ84VXN3BV7IMfnv7EtJkoPbH
UbwFm7Gi3giGkl2wrZR12MSSPSjK525glFuOzjvdc5UTpY0Blj39O9UpfULXoSRN
46/i10US8KRoKsBkbzrTpGJmEyK1Jk3/3XV5OrAX8FrObbsHt+HxtvuWxn2YTlrS
VR5uU+q1/wsBGuciIO5Ttupd+n3IERXTqYdfzj8rj9JyngJbTI/Ws1xBlFGDlokr
T1HwRtjyE5EJRx+FANKm49O3WmrTcEC1eXUyzoaPYRZ58ettmUVT9LEUHQSncCID
tQvJ3UzhQOxoMyPAI2Z7gTEwyCk3CZiHsOTF+wNLB3d4ogzT+uqILtvRCXlctcoC
jsJZ8hxE52U3p3NWsuBl8Vb+A1AQq3LlwtA0cmPcHN4814PWapp8N+N7yAndMm+8
pBNgw1GTGS35WJdNpETMK4adKNNEo8izPo7nscFVywBQDuFpsYNE+2OM51b5YZOt
pimZbO/aXoIc4uY4KHp2dddL7Yg6rT4VMyKu3thO1t414UxcACOsSYlwc1Z74dGw
TcrwwYqDGXLoPpi2q8LEOCwkCsPF7jFefPg4ZHolY/+q6L9pcKzk0ICbZ5/BaJoF
jdpfCQKHbfPiWT5usnambWqAh/nK0jwAvN6CkPQ2mSA8oeth343Xoa4t9fvb+uJ1
i7o4jzflaBKK8IeR0+B0kIshPUpisdZxcOY1srDkZQFsAIreJ86hntk78GPhplEA
RwPhjDTfY+UUC8E3dtu459MEVi+by+tGdJPk+kuW58HnTpspKAePdAUAUVZ9lW6V
UiM1kzVpfhdFPyjDP+av9sWpqAFtoaxkF8EK+ud6sCqsolr+N3SK7wAu9SR0GvoV
/AOHt1h7glAgYvMoG0Wm/z+10hxuqFERq9gic8j3HdtTGo+94kOao88VWgibRytO
iXQD7RZwlA7FeWmRwa0BIPMk9TepfKaoO1e/DpkuqGeMedGVknGGbDIsQRIf11+b
ga2b+ZxLAKJxDTPtueqDaBdzlRfPQ+m/Uhvd6+tJaIBvdl8rjSmXdWkeEhKkY0Ks
m7gEjO2mc7uhm3+EaPwcEQ5tMABlvkzyrtFEFBFWojiN0sIWFSpHCtR6q3FTWr+z
vM1LlraHMMK+qmIbGC4j5Mu9rZushftKqEqmHEHsBAfx7ER3s9uO1AGPM1OdfcYN
wu9eUg82AHUN25FxPP3Mf2h5xlIoe2jbx9Df0ICIhgNwI0yW6O7gWXdxt+ksdw4A
E1aBTS5N30SVBQrEUvx5/1pYxaDO5mncpgjnldMe1IYKPPZHfoFRXzZITOcY2Xvw
FNvQ9yIURu54s2aJ+LacPtmSpqSQ7kLUkp6J6fYpcRKgT9g3JYhIPwGseoTVCELB
ScDHG5GaPAfL8TUfZ/DktdkA6PJlnzOZn8aWP9GJ5f+87XGFqRUGofP4BeHkKZsN
lNz81MudAf0mUwbxzXUejf8rnasXHBYL0oGVngUAi6zmgefTRF89NwhAFUcPf9hx
CeY2iTpdYfhcOt0JvQCr415al8bw9aCPxiX/YtkKiVUoAJBTn8U0YU4xEXjSoUnX
G7sdbQowgGo56tqPrCs60AKfV8OtDFz79kyUKpPxTxMZGD9k/O4fsntcrBc+RRL0
/xuvmLXnzLN9pGLSzS/zQtmNvDYx2VPTDOYFEwXAx/fVwy71GPELRgQCTyDxiOw1
ZDpxOjbI6AgkC9WG6GV6eGnJHV6ktR2CW1ahjTmfcIqDJYZQ0VxjhE9JZeCVC0Ev
SJbm5Tp0CvBjzYqUYzjhJPfZHp9Z5dGyiWChjRAN/1JNLdjgTE6CQ0JZSPFXtRqC
5faa4B/g7EYRffgnLNi8r/kNHM6WaAPEOzf5VVGlbEyZaUrMPyPnBjf6luWGaPAs
jX1M/cVIQh1Ec7wx8EDxS1IAsmjS9KYvQ28OPAl0T/acrr7yVjroM7VfBNlbbJjo
5bJWBSochGB63f/2BxPoAPU3IUGix1Drqt1kCTyToJqq96r+SMusjRc88cpAYcan
DhZFBFom6LFPF8werOWbbBz50zIAlW4Y2UcaRmA+PdeNWHDk/khvXFq7rimiwHTs
qKQJzg3l/BuwbJXUUaX+VB3yr9JjATncQ8YxnK+P3ZwynbByLZkR4YasST8vh4th
wDzxoHtK6Af9Q04azO9MLRUTrmXd9dU8ZlyyYWBydtpzzq6uRELSMdMAEXPbiTuD
sZphvPY4ZEtPAD37U/3HQKZKrec7Xq53qeRRc3VHHF/t5LLOHUEPMen5TiTZBKAM
44ujl0sTC79m/IzKMEQoxqdwEo6WtTxtJoXIPlrBuAjzTSSKBudWhPDfxvwak6Fb
2uslmQAk84mvj+Sr07cYtskP51e5jzhl/aCbRhW34sxFtPt+6ibQsKdyagOkgLCK
x+5hlP2VeHyckaYJZI0n9y6yRESB28YLNazNCeeyN87W/E/zTuyQZawM8sCwwtcr
TOhAk8cAjHbqhckWXjXaBpFt+46ZeaEcQyPGHKdfgV2qSrlfnXh66i5hhyjtHdWQ
ImOZRVYwjpol0nghNcxIaWU7YjSubG/2yMXS7PZaukw5gyVXFcwNAmggNugAQKvR
dibRgcvXX6kJ7rQdF5ZOkX1Vajj6AUe8qH1MFa1FsU91wNWyO23L41sa5rTibzA2
fdGBurTUaXCW8b7JBW7zK22rupPpWexKUbrfQ+BvTOR+l1+QaAQp4Wk4dTu0vl5K
PLCvDVsHNwZG1+TXvWyWipTZm9Ud78EFH/wB2CvmSewk7G9xYBA/90rRqSn4Xnut
ynQuqaWG44ZtxNEyvZoZvB9kmhuE/6XOeLN2UazkqzxDHt6pxMf9zoNE8xLIa8rJ
CyqcU4YmjFroHqBvedWBNcz9lKlgx2FIgcM4woNV8cgs0iogNbeu/MIAr1T/KZBm
PPqYWBqFx2EbIOIPAb5MnM7AIN6RTVWredF/J4OUN66Grh3hryCzYDZt14FyPOXt
kEa3oYzdeSzLpX4Pgief1TPBm9+a3/b3taPX5HHmPtJe2hwA0fZL4sQllmW2Wylw
7qYCkcjZhBoXtJH0N/fvwTq0+E65oAnIYKxbi4baf1DFGCWcdRlRDs+K8uhdbOBI
zEUiTnKI461Pu7RIwjvxlAQtnKujNW/HTQjfHSj0Z/eDCOEMU7uHnidvzgdWSo/J
TlBL8kLFPZYcmBgNVKBKa9/UIlO+S1oIbxntrHaB1EiJVt5vEz777F7DmaCAQec9
mftGFRG6GA6MjrHqDzC/XpfOhnq9ZQZ1bNg6Gou4dFIumAQ5c/vRSnxSwhrM34EF
ahyY2nFow53WBtSozEajeY0xQ6mS1i7gimV1YCkPYfH/8+zkMFOFvWWsqPSLBo4N
kGKRYFbMFv9MjfIgnU/jLJ3iP1grsiSt1OSEKXtuGfcRywu+CMeyUTGEdS1iZ/q0
Jw2l+RLsTiftMTcR5nwg2qPe9rLa6B13GaWKu2bmVNkEsOCpB+SO2eehNw2MBKq+
nVKEIAsOCKedsQDPMJ/Ey1cL3xilmC6T9qlQx0EceKO8Q/jvI/iUuspPU4JJCC/N
w/VIKtX61nWfr5tfONQNBkh6zIyldqiVQu57WeX5Gu7XN+S/P72l4RT6jzt0UWGY
uG7zHm4tsDfqhBSXPozOiMNNqveV88UZJMe17jy2o/fXGcGR7JJJ/9SNpVGpQkmc
pJGrrPlYgOZlbmtHPzVhSr2K8IRnGaZOR6T3uo/6PY1QzNRmE+1/LPEwdXgdHrx9
wIjDerMK1Kts2BLEGtNxybR/pm9M+lrGXJAcK4kxt9hKpC4/quuqGYCiXx2RziJO
T3ZTILTmVMu7RX/wdx9e2A0r3YWtv3GTrxwP+4UkR8kGF6VIwFldG1q6NcB7pPR/
xajL6x1g44Dbx4qyP5Jm6UvGMqkxJE8WPHy2IhNm7x9mT49eSZ8qBP/CBX3zG4rs
n9MTmT3Axhb4POS7F3xwDfSfzot+N/3Wz40kRHhMz0dTGMIAciFlZjh5e77qTUbV
vGcDA/kcgLvHJU9RgFCCUI769qhXwIzioOQajpnWd0Qj142HKzb/1S/srt3WnsQx
wA9p0djxyMERYktkUD7LrpQqa/D6+8Gt08rFBumL3V9tMEPdg1tv0Un8+FFDFa5Q
GhTYmC9vvVS+QnHBTBFYeHfgTWncJFYDnxkt8hePIFV+V45YcmU6HAWFbQOw9L+Z
iI2opOfEJeaUYPdtpPtBs8qZz9YPTH+DSnHl/tFyIr7tpY1G8Oix/cy67G1uwviG
rIWyiX0EpJM3UX/OnElwucBEJGQl+OCEx34n2BOL2F2j5DHyZbr5XNJLGaGomXVD
QK8Rs6bny+1UvqWIBQW7rFc43Fookft1o3Hb+ZvHNVR+BTwcZ2OnVtdDzGnMDUE6
hh22qRkyzu9z5cWMrKaQj3Fz5iSiKIK0u5fFfUYWo6Q5i7YlP48RWH2f3U7b8stG
wE3WdAJ02s0/ZJQJI0uXQhwt/ZmlIl3aBGZZsEucclrIwU2zwBkvF29mqwH9O78G
tUCrcqeYSwfj0TOzFJNg1D1j2zL1TUDKYn+mitvvWA/6NUtqY2dx2BLV9HfLG38i
Y+Q/K24+9/jKd6v+Sy353+xDFo7NMywGUHiDJJAgIdyTiV2v33W/oat1dMVqEU6H
O/js/gERtck6OYmY2Yz1UiOVPe7XMQNg15Vq1xn43pV9w2kgNRr+bB4Nv89FfJHh
k8mRFTr2Fb9H9eq3rPd7Wo4zRKqIwfEz9xdYgHvBNRMlLKe7+BxbU9U1g1lenRYa
NK+9MnPRebrj/URtu0h/7AiV3XrcTnCapXbeC/SqTZDvkpNYRJXAqyhDA02Nd/60
rG8Iz+byjaa9ufAMgUd+Z47IzXB8FtItB6TItUZiRpmLIHa4qziGvk49Oz74kgyT
Znc3laj24/YrWB8LRI4YE9xSWoqyMksaQrW7PHTEgv/pO94s7J6iiBSfEV6L9N9s
2/u4rssYC1bVCAcP4gptRLinAGb7jBJO45+SPdqvAffyyk1KrXCLlsdcJtKQoMwI
wPUzvuw08kkaTx/a8qodC1Ci4KHuZDwPGfTBUwBFXq5jPtDPIE10TSkG3wa+lJjU
TuHjILJ2mN7PbZfFLeSNXu5bjDhatJorXolifllUFzB3CfJTc0QY++BKd7Mz1KxD
g980b8aU28c2yxYwwqtO7eNXxasPPCvhIHBrtaNKfwspqYjprH+uRll9T4REF1RR
BhaHC2osXvxSrHhbPTX6qhgGXCvyoohXXAJTv1mDcDxmKnuWGz4Zcfbia7k5Atfq
zlvBa+2jnyX7f8YM3fo72AQd3aFVaBf7DQxUolm9qFTeGgcuHg/ReTxYiRmgLabt
1lPi3XfgjWjh5HcsbAIsJTsUd/prFXJo+6unz+3mWuaCyLBIJRF5wIGD89FGvg+o
fc2MGEqLSbpPCxfyANRjS2KHM9qN+MZqnsWTIp1Co1oJX8fV0vSxrBkrXG8QPKh0
En9EiaYkXL61jG1Mw83gNoDKaf8yoondCJk+cD1LlCwrG0gHuaWKvsga8MB+MiL8
rcbvIyuzS/DIV807rramOW27dGRg7oU2+gFZZucveImCW7QCJl/D2THj6ytdMB9s
Eu0uOufUxyZYtuS2NoofPsfEDDFK+C87dWu051Lpix1ZuG2n7Qg1vOVAEE8NOr4P
Q7/1ctUNXzaBBXzMapB9gHGxUZYuxRow2ogOIesZufka+TIYw+Sbls1hQXsKw+g1
TINQ0yEnTaMEjSTgZff5ts13qJ02Pa0sGxy6QfqDtWCrkp3Q0CIrZtWMxRNv0qxo
kSPNun4ZdxDr+xB1tgMN94oF4uzeWLlFs1lt10q7tL62xjDkbvMtdWwszAP5PiKl
QjaltMralNKDgd78akxRrDPCOrB+HbmyzcgZvZS7FqCU3iQrMi64dek3kDZh+3l7
RnVbIqPuMooai9ltTAki+4XF0fHlrEwHKDWtUvBIzEhV+UWkVOcrJJfR4a1+kRI2
eY90mZ33xfJHQC8lXvZFnHOu0VhyPCf8+qyCNjiicIa1R8JJ09xwPTL5CSV7flP9
KqMgMk5DkXogvBzBi67CmyhF5M59meTX6WuSwApHaMzBnC6Tti/Wap7R61Vb25ON
jw4x/QXPIcVUXybtxnosrHlY8t0hCFwVfEWUUpUP94lnt0HmHtrqSiytOEJb4Ujv
7TKGbxEdaqvsLKdOl/S3U+TVMDNI4YqETBuRlvLNQKBf4kd7ztwNnZlCTFUUpZIf
ZYShjudLKrXaBrWIEwHGX80r/3+uM7pgIa9Th1Pmy+Gue1artcH5IW9sHnffOoSy
ioe60UY9tK5/2+bUdYhicVOiFEnFRWTAEHxMg6lD7SirnT0Kj792fH5XCx4nC9QE
q6T/QFAJvqVgQcIvX2kBAAmDT0p/1zWKWKtMdh4RCOVnzr11GTV1js4AbUUpK9xn
2uRU/C3+BAHX3tkLb/TAPKj67nDCOl8swC6GTwBm5vG6PWjYonW9KAbclihQTJvO
bFarRJcPfmEf1lR8KLx9AjQlW72jHhtKeQr+WrcaLoB/KP3raoTOudZ1WP7Xvf/Y
zENSonydwBy15mNXwQjOEg83bqflRFQSLskz83Ea1TNUhqd4NZtmqVR4CGSmVwyG
jhgEbPDleinCVnvIBRguj5yzv554KGmS6qMJUlu4mvKonayUf3x7IL6rmmr6Oy4i
XGvo9QydAHuiEjeHeooU+78rmo6nXcYJ5Ra3kBG4qDTD7CVLuWf1qltp8PfnPBHu
eCZZx6BRyI6CMOdaOQe9DwBeR8nunalxaQu/3CAc9iYbTc2CRN2qR5OHUmKWo667
6ixlD6LWSul0+V8dM3Lyt5XQLFZuu6S31JHiesR45B+O51dtIED4b3KpRG820Uck
ue6jopBHGAft5xkrOzpvqLPACf2S3ccMgqvdWaOx2XRKasf1rm6PFoWwBvk3EVq4
rTU+a2eGe/ZiUFGzQhuKX07k1jb4d6xFdyHsm0n1sgPaGCYYCteIS5dQJ4Aq3ywZ
y/z+OG7RCga3XruIw+5Utd4oeKiDTYd/N9ADIMlhZ4uLN6yTpUDFAWJYRfH4y8Nr
Psi2gnl/ATFKeKiAlLL3rqH7+vAISJ0SHCTQKSBeCQNA9Yt5HFBsuHZ1uarbzdm+
sZhXfmFCWBkm9VoVJpbd1LdbM53js/WN5GWJN9VAcTm4jYse08k/GMAIuiwIorC3
GNXXvvx3ILuyvsr7OEAzhV8nkPiKna6ZXPY4bUczudaslwPmxZUYmNzwzoG/hIF7
aGAu2aWQfJPuYab+7W+I5rU2zqIzoEGpjXHvt9as/jmuRrnURMzxy2nV2Cwzgyxt
A//DrlhkalrSl1ON2cUjdczcUhMc7JnjUrgfyvXt5IITG+O07l0FYyO2kGUq/rxD
1DsCk3KQzYtQ/UyLqnGcuEZ2wah54BflBPyjTJ6NqcinWLJW2w6LWdq916QQnxGV
dnC2+UtGGML1FVLP/ipu6x7cXz5/GHClS4m6M9FJNeufD56oQemMZPiXP3o3h3Qh
wiuk9oo0EbwdrNHWvSgfJYlzYmCAOXsDJ3rNqsU1jYMFENPjX5ZILW846cnriHnM
XQ2vF/Fh9Z/mAGBUDMxU3IEuOS11eIHKHdq2mhmpXeqBHQDODDLuxrjQisgqFtmQ
x6C/pLIePRElDtYCW5AF2r9E5AtWRj1jxgIPG/5p+Bg4Edq1/dPEGFbKv0C686U0
S1P+w8+3gzbVwyu8R4pNFY4XSwMjnwsvJeN1Li5Em9zibKiWVQRThZUwGzv7EhWc
cNsWET8GOyaE4ngTIQR8+ijI4LFCMEmz+EM44RoLlAP2Z0pePeZEVipEZRvxazD1
R8F6xVy1SIFQ00LGMBPqsNJRhuA61E7revcJCdccjpNfvsJW3cj9+rdPt8W5U81i
eF+MEUayZDo7CAEBUcM16EGOMCMoBvjyyQDSWO81k/hoawSGIBg5k0S07qqRAXZ3
fLtEx/zwr2Pd3plr915DkMw+9pXIjwKyb4ax1AIF6hjDijbMvr7y0TnnQ7DbIhaH
GahMMdAI0KJcCMFo605bmi+zPfRM/beBvwbZCHlob4vlJBHPStj0zEQyc/EJnZ7l
Tpu8/4bsXhLoUQ/+y0iYiX+a3xzLHBQbqCKqxl1VU7lVWy+STk0ZLSvZ++f4bbMC
6NRq+1tKTg3tPCAObQqrWm0j9I38m3+nvQ0Agsg43UuR21/BoZ85jxvBbyhxjURA
ydQJTN/pt1cFvbd1ExPFVf1CbBRKTm3N7xDQjyIz9qKamI07ZR1/TeMsA3XUXdcx
Mt821lNcZRXcOofh379SDkGQhoy4MvuD4UZJYyQvGOjcGW2f6vzXcZHt9Tj00V7d
V2FKmZzxaWXG1/MgMxZtVIHrK8hFWC2N3WWNq1XXRCw3Sxd8/Fi/eRQodRmFTKMn
G7UHYmaAFamt1G5QlfJxOQbVpPcpDB80yDkSSuD0rvxVRi2knk8L+CksjmxiPWtx
CcFdgttOnoP3wfuw3g1YG+Os8nLoWKFnE3ESBXlg17/raJvDO7Gv3j/j7SDvzgh5
u+TMyD3fnu/MbXi/Rt0UEhmuD9Jj2LxU5VLoAGsOloggaggfkh5xpvh5kowSBQjK
dT5ko/w5TMOcP+shnPTEO1p/0UZrlSc1NqtdNXPeIz8i4w9TXcvuREWyZZGeukw/
8F6yz+/xZdhstTt2jdwPKHJJ8BGqKktcxJ0U1J8FjO6CnEGeYt69RtT9ygeS3wt0
qTiMyuZp6B0fBFDRAvEmb2gyrdwIjDzuKo0MSly7eDWCHlnymcoN/AC5gbTtx6a4
DDxJ/N5dw7YcMoG8yRsKBC1Xc/6706guZsJWzslTnr1xuEyMU2qf3UYGS0Qr2SRt
cLBc7uU0PTadjvfAxvRqoZep1UWBnuZLfYoUIg6L2braLxtl1HrpZ7pkQCcJHpSe
Nyghb2Ecdnhf90ZjWqdXwYElSXlLkcL07oo4YhvDN/uDp6b+VE/vrMwPiFRVdWtG
6Fzg/tGQy5B4ISb1DYtFxIcy9VBkyv0qbMPuED1UMBpDFm085JFYa0XD0bY/6Lp0
zQ48wyJZ+ARQjLH8E1RhvaaMTEUrjv2/Ihi3+I8zxq9XXNUaRoaj6KBXMVDj0D4w
prYJ5ala/tWSgF98F15qNiV1ZAwNL1GCtdTwQFlFukJxNkoOXladyqBEnsi/JwTe
gJXIeYBKCdffr9kL03BXAhunuE+qtxO5DB/tRbvLbO4phlpC1xDZVU5JxKpd77t9
vbcUp1xOQCsbgrK5j4wpizV7HMAKpE3fKHDxXH4GmNPIj8so1o/iWTE5Y4bjRlZ1
BzWgMHrajWm2bMYkHQjNq1IP+TVKf/ureelc75GQleZY45QmoSSBk/07DscJa3ta
NFDfzAkgv7R9/lPkHBaVJa0TbdYcyPFbNIe19XrkA6islP76SbaRnpVBY4lRBD7k
LDvtNBQbZEqzn+0tnCu/bLrd7ty5FZdgOj8N3p/+iXmmiSHVXOjbrI2HyNCNmgNJ
VgZ+hbsKX1LbRxXxeH1aJnrTb95Gri5xqodH8nXFBhntqwaByjhx8SvivqlOmg85
SgIviTGNy9e5Ba14XI5m/s0ma9wkyZl4iTGEY3cl2nf0HHuCMWH+tYPEaDdbx8VU
wgfDlgXHCKvrLNzaU2YBtThJk64lkoPDU8+I/AQb5VVemHCyMKooFdvdrZSIE31B
0OItFuqvkDjyccReBzbCAn4+IpZQ6IzRSyFaSnKFEaxA3XMky/IeeUjUIexQaQQQ
S3BKwd9HJKo9ofV5Zbtu81Xt2ZeLV2wApGKyoTUER22upMTrbBvNBbss2pPDrVhe
mKvs6qrfo1lQxRkNBZWxFUctHxjl3Pm8dxqLwSLl39pwyCz6llGW9MO6J8mDZlYc
hg+GXzTqK4sdJMeRHhje6itJHVzqSUEWacv1rk/AFPnTu9F7GwybjofDbXbzN5yQ
ll0E1fYgK072NHwEYnwHXXpXS/Du+ph3dZAmFKBi07ypNq4J02N25rET8+Vlupmj
s/JuGuUmPL9DIFRnV0b1nTZsxIUB8ncylj7NTvy2RZ0QhRiEEGtRAllIoxRvJxfx
2cZKFJ/P/BkQ+izXu0vf5m0BLvzcrr4Pq7wvEJu7fANdftDYQSeBGnKIlTGGtPrP
vJgQ7YJ+PsUv4jxKJEjAnpUjUbuR88QFJO6hxC5Xe7xT+6o6p6FAKVYX9C4j0/q3
htUtDkiVPJOHvzl7WA7rmDB7Lb6pHPSgJ6ODoOCLq63dksre7dAuuwEwuhZF5bTh
xpoNdC6eD72N4OjY8BdBZyGAGvrm3Q7+guvzyi5XqE1RG77pHRIqvYEQQzCmQHew
s3DUTCtwqeIiRpp4doQ6cEbY1n3fe3dj5nWPKkAj+0mgeMYBNB0n0CQzq/0JBi6I
dZYMWy5LWoUDHba805tTjmdaDCIbMAYYCyy7EmkUr7w69F62Cs6df1hx/hMJgHas
q31bPQrEDr3tDT73aCdu4JGBPNkkZ35LIT1ySykLIgduwMzQ59hAM/CWX2pgKTAf
AcipCj8PJJ8BZ1utXpkQGQV5HvvCNoSbu7+Ogkr7LRK+CjsjPfQnXgWmakqAIvVp
U9e0kSaMvcGpAY3nZ4OJqQ1U7YHwTLmoC2fZwWI1GNizatatyAByjuRWpZSBHiUq
rPrqAaz7ULv638vLsUuWJyesTm4RTtt1NvlD6ulwv9FOL+IRKaLlY4TThc7ipbT8
5NsmFVTl2LgJ6bUWg8EsJUD9Zj+lK82UBQvcXjW40aR1gAcEYSvniT2z9BpJ6qyE
uDzyUrQ14jERxu2XDSZPspvlrP4qaw97j38h4o9jmRqjmCX6dUMBKjhtZBlnVUSl
/PH+qfWarpdUsvF0E0ed9KW+Cfof0TuD6Z08Y++lDJ2II08yiSeZ1WOntQu2zEsv
NzVFbmFozhncPbvJoLC3Sxsd3dYUPfqsSKpRGQtRotT/fog9WRgIeYRPCeVHPcXu
wWLaJgOI0LO9eNwo25eUk8V6DjkoAY4G4eKL1HODAQQ38ws1Gn6sHi8qss/xNT5f
Ss4H8yIJzBZQiWYSUw83XMiVCpDq6NRJ7Bjw+ZuqTuDm5wMptbQuDXkIKi8+PaCw
lMqlg5+u43RwAzW9zCYkgnAAK4ILnhzCRTnXQ2urHU6F9N2sI8AIbBX/ihqUOpms
Rg/DUdHzWgH1Jdlc7jWCXTIdGwXPmAYYYo/Se32DNxyBCOFH6UJg+Che+LEXNc3e
Lwwcmpolfph0zR8I6LA4W1bpvLwLhpfB2A+j9LWVn5E8r4unk+rON3ifv5SkO6l+
BiQ5ghR583Mi48chIhh2FsE2oljxhv4zHREXe67ZizTeH7GmHfgoSkunT1pEhB6H
th2hK+2Fupr/wkrGsvJcVfuZ65Lx+KjjVzb/hPqVBLKlDfFJJOG2wA/+IxX3cx+W
UvAw4uwDKih//axu1Tz8cfw9CbUBDpkri2yYWfHxTB2ctWWZNyr5TIwKyy51eqLA
e/AkgN03OIbkPsMjfUFW/TSuoDnl9ZOJNaUzo+ynG33AdnHWxZ/NFgC+CdhW4Laz
mpwY1lCrHRKTh48EPvNPQljqzNCd1Y8fW6vETH2lo3LMEAUc1KieTZwKX8bt7vtR
O/CDyK3cRxqXYkQmEzqH2NarhUK41lzIxsBhPn49xVBAL9IbCA9lYumDk5PIKkVk
jDyLTUEKbBtHLVadjlHGs+UitAsTUS1x+59LFs0xRcTiLsqdTNVLYZod/QRhYIBT
eVdVGP59Pq5Tw79c23r5Oj2LYaJr+b4N2yY64xBOYVExvsebY1bbwns5Rio2S7xB
WY0/26baTWRl67yvLBZ5vtKMhNI0Z8ArWGihDYE1VToYkrAItnXFydMCf2jweG/r
gj1VRA1Q625wTi0JKMCsKRlwadxwqWPwoY4YhMeRy4ecV/jyIAbCoOtitRubU969
y+XISdvYEX359nW7OJ9pXUgrSJYpF4R25syowICZN/djw8C8WbnDLq+dZEZ63nf0
Wp5DGJiNG5LwNS2RZVK9kAAIKmfQaKYjwwDZ3kvHxpbmpU1S2Ry3dS4a69fCoAv7
7HQ4ioAbt86wu/mS2MAVrM2XjnKr8IAGbQHXzyNKe3APtgI23cxrT8Zxsma6KkUu
Z5fJpzz9fwpyZ8Xv3kL9eQz2xGRj+0RbPBCj1ElKNRZvt1CMZlshTLmix7okG23Z
NJSPraeYDm5/YQYr03AekB/ySZ0AgYwhnExqXZ++AbZgKMRfn6rDW8yK47uTJjsa
4ytW7i5hWDDDDSGm3Bf2z678UZDA/RH5CkU5mmGoUgAwBea6rcmX4wYABWNFwXTh
FCLIXHRvIDR6wh+sAyCx7VVgxd2NTpcxpcXugumPI1i84e3q2Clz5hwAM75WP6Ql
5dPKgP6KsXvcZZJsnWPZrVcahiSTcJwcju8YH9Nmvid2I43NPJzW76afFM1ua1FG
OIdmXdWwJWbUHs4+wPhdTDAqjB9bzPeKRUGqFwjW5adQaSe/mDjNzBxvmwl0v+hw
EVjr1YQ29xyQyxJbDmcswgUqW/0UgCr81wSEuxXV3Q2+zZtixMgmDpiHPcmgXSlC
QtN5OWbhtM1EeCokFH8eKigvOPlOhPYi2gWmF6/tfWqbo1h8ad3QyY45IGKr0I3E
f7Lq1fh0J8ahFcA7JUM12tmXDODOuIOxWeDpoRhlHnLu0s0JE+amA5Nq8k0jMU/d
pBmhtkBO09mJRgImZtxVly3z+0ipq9JZEmquOxML292S1cYQHxGhcgMJ1WetvwPL
l9qlPZn/IUpfBNJj9u57ujAV8ocv72SDFDCQoh9AM40raHRbWgLX1tAaUVUmTpU9
rvLnwFnl306RxGtlQzf9wrhYjNN/VTj/uGFla6Vnj3HDv5kbynzWF0qSneOS2jqy
qojoWDpK6YWhF/j7Gi3txA2V6z7Rsa4S+FIXJ/GrAgRfxskmvlBr+MCdBN0u+x7O
UnWSJUHNNQMPq6Lq0rVOoMIM8MZ3/CnHFuE4ZNctiOQwIEvncJ/cXXOW2jVRUkuF
LYnP6n+Xf0WXXK9pKe4sTlSlRZbq/W23nL6vnKSV+r9NtDdNtpWuisKgmWmM/tqF
6lenOGdnGLeA5fo/ZXrPWjYSufL9kW/8OZG7DjR9aPdNCP5hK2f32i34Ookq1py5
9sQ3qcBrAG8FcN31TJy6EBOwThul1qEZ/L88a4zo0BtDALkuHZGuVXBI9JPW7BRZ
KgDQkZ6WY0VCN6YruiM0SIGDEOJ/ijtqc+ULEyJSlZ87239dJc5veBSh2vBqgodi
30eQddWcqi8EhsdoBWY1MVeu5f4dAnr6/DoDloPaPOn4o3L0tNBhwgbIDE7iz2YC
pPF4hGfILyz4rXZR/YSVPn5spd9y1T8vqrnGsHqZNW7HPnpPSs246zoBgfVcEKuR
Ri/lbKTXrcYBmWY3QIq29KWnqhu80g4Kf0N8wglUzoIcAdDoLcUL43fswn4QeNj6
KlHzw72B1cBfsRFvdASmq190Zo6w2i9vkF7EZF0TKOpuY7rL+ltMVzpGJueJZjZ3
qCaAz9fn+3ii9L/WHoRXROefT79dhx8x/KNdUycEdGZ9pPjQIn4ifVsY8o+ExeHo
U/Gas3GrlNMW6D2Pn/aMN/jD5T8wA0SFQTwxYGDP3o+OZzJDaOsNEavYdl+EXCKg
hGd16hV4OcRoskrJDLnTBuVTW5Vxo6UZfMOs4bD7HQnY/7Wv9+yO7Na1+C6PXkPm
jEC2kYY/a5887COtShR6DOgE2yYw/qRwX2KRCezCYTRfv4fRn/E8SaHO3rQ5lg7c
FI7k0Fuhl+tgNrfg7ArV+oHCzL1TC7JtY6iwhfkOHsRWiQZZ4bZ68Dvaz+f1qGXS
z+Z2LX/i9mf3AdqV2lHmYIzlnATTsBPAXdEGv+2weoCcki9884YvvNp7LuDIONNg
cUpCVOLiS94ZepQymn8WY5AC9xJevutlFD6BszmYk7z9C9PjFvSSF1kKRy0gY4mH
AlyNefda3E7h5jYSLyLICKS6FbyIeBU9H41+qYopII08LrMYCDTNAB+1Tv1tobns
hotazb4Qsdc9OH7Nf9e2JXSi5dLiv7eUrczxE+9g2bWPRVFn34hfKHW+Rb/oAv2k
ZKtP9LeUIQMHSUutQVaGzjC1FDp/dGIj1NlqlVgDBmiyRq+Xi+01s3xXt1DKLa6m
/qhiHF7f38iUoxWPPuKMWjmFy5SroDEp5SvN8PE0fmJwzxJ0999cajf327VOj8yH
+k0fMd1FkWM0tk5nrWy0rdDHdQoYWjmzH1KYuybwFMi2/rna82CQQU5K0v64Mn8F
s34zAhdwXLI3r1UZeAfntFI4M+1LviA+1YiauosJ5iZyO/222jMuO+avKs4kIJNu
XhRngh3gafx4UAVsl256fH9A8Zo9+KVA/erhJsm8DbdqVjirBRbtAYba9KWX21GX
R44I+nM4VgDhNK2fBptCH1w9x7t0DqsbgSlruH5aWzjaNo5O4FHCn5nuSokmVVJO
VH5VDj+nyoqSKekfK20uo2Tomk71RqsZjwPsKZWprcNjM43u5LpzLZc+8NM+lL7p
kgSOqLbeQxoLwiQv51K8U1w8WPlETnJ4q3MHACeJlAR+eN4eU3Cls32KhOTWUA4y
gSLVFmtv8dgyVrFRSa8LpoZiY1JQM3Fey3gaTqZwNSvRlKi//4NCYenN8iIPOKuT
Lcy036st20DjSY4MXpG5WlEGYsHGHDB8nS28xqxaepp9HszE/a0bQjVtNL4mBylX
bda5BfQYSUkEv8qbvekpmbCBmDWpKD9J6hTL+o80BK2u8QSSy5uDcHZOtvWjqK/C
V9u/hYPCPZAJZ9yv9WsW6X8T0pIIw9NX4+z6wcsB5R6WP+5tEofEtso6tHD06TFV
fSOT2ElECyw2YfpssCuKZPibVa9YNmVRXo0vPNIMnoffc97FMFOQKDQpotGP0OoV
tSttkjWONLqkx97dHSfyREQwEkBhh3YBuEWYHx61LTTd6a3OAZuSFdODsa9tehVI
i48m7GKQQESZ5O4rXKLraJOGV8HFAT4Zo2Jd0fGWTGmYBgYNUQFwy+Ttgin2Mpuz
9Yp0VsBZ9Z+QzrwaVKhT16Zi8KHiTPFCQOEJCwaVy6J92cY53+XQI9CKF1sgfcgE
eOqNMgslRk7i8RIY462/biHdmgzB3HKU7T8UXjZ1BAgyAB3/46j7bRVe+JsYpZNC
qSWPbuezqaLyHL1zfHNZIw6saZcMxs3lwoWvyMa16b5y8brnPtynTEaI0E2Q6Qh7
8qjVlieZsqy7l3UWWA+UYyjOHmtWQ6FPz2WAhVH+wCFmkN6nef7rWFM5IINo39w2
VkLoTEEHctNJ4bYNwLRF3e7IdXNzEh7C6vqjZyyT0c/b3jJWfMkzs7+MR4FXZvi6
kkbyLEEBBe4Kdes0jGpOeN1bxTFCZ34IpvuTtRHtQcMMaLeHn+g9GUeCLNxIHvHA
tJxyQ5VqS6YO0YXcRdtD80MML7EzTynfZ1hxk3kAAlWkgJHtn4jSws1bR9qpKKC0
fKQKNXY2M3kNvGRu4Z5IoAbkdA4ha4pxNR+KvPulva7y7SRQsNvgbEi1Mo4Wduwe
YAdV0lbPAhhWXgB1u8Jwmp6S2+0HaaLNfWcojo9WyFUu+tKf3mrBBl557/coUVX9
y2/6KCD77W+en5dO4m6HK/yyO8m7v4HjuIKjwsTSlKehS7hUN1i9nELPdS3WG8/j
/P4giEFut37hfEewSyznJsvA7GSAydISESyZhdubrBvMpHVbtCnmPclS77jp3hes
o8MTO1d3U3+88rtjOgdLO1xijdwsNX9zMqf0YAQPLbQ9888nkOJfjs6uG00F18IT
P7COiNAizC081pBDS0lgu62XVsaNdDoXN/GBqjgwX+HKrmHi9yJobUkvgr0o90Yc
woHwXqj7H3jmapX/tOflY3bJZueaZm/Co7a6fpxyuLnVYqFHYJz8o3vikbrUl+kE
bzLlQ/rvezCj8KC8BiUqargOZCAnLkZEuBEYP0wLeeQUbbEYvecKjpwozMRcXA+Q
7s/fvL0z3hp2tYvB1xj/QNpU2C6Lh9uwpic5onnrA6RlCPsB0Eo+osGDApjekO8W
REjr2AUX/v5lfjskRquuL51I2LHyWBOT+NJcsTbkxa60oBUsnTwgJ0As9IQCepgZ
8NWljcW2/rwWPEsocIwi1QGthAJdMvlqf/zazuRmGEsOexoPeJ98qwe661G9SzC9
b7ByNAkNLhJnwhLqoP9F7eWVtQC9MirbE1Eh8JcCLxkL6BibHLWD5b6Y2exYnvFP
CdppTc8PX6dMHC9RmXRXHe++AhpBIwPiEQYhD6JREVwmu3OLCTcaJ/bOPmBrcCcH
SvxQbvLHDnqRjuL6AU+Y5DgqMS11z0RKlKMEClveryFWkCCPsOx7w7weSAOSvBck
8TbN0XV8mBGgykggI+cK4Q52FAD+wMwDATHosXs9nELNHnSBThdf3IQszC4inzIy
rjFOuSRPlKPN6PHnD2V+EG4+oMxK+OXUb9uNwHDy46zt1P1EtBhEuSPsIPVyuvvJ
pFx+54SEXm1fgty+gVYta3sTFhKVmNr5nmez/loWrLczZGG4x0Jjyhudpsedk/y9
iaTmQBW/F2F8nMku7s424+xloZWgceQpITL3XaTsaAnyvvhNxwSsLhLN5aH07w5E
kXTU3u+mJqExV0bAfYd7xX4fDl0cUZthbyemUM2rCfp9OfFhCiCIhjcENHJsTYLI
rZsDrdfNvB7lgo20s8xYI3x9bew8RBm34QUDiSVwIXBi4RGr6WK9K1aRs3+k29+/
0t2q9KPo+hKy+kOEn3JxO137xwdCqWilzNzMd7s0UQ2G5rR38cIyepDJJP0NubsO
aNjWR92DBlPH2FpZP5fvts0rRRyFQT1q5mZkAblPYHTvE57EuTpi/X4fa+ADjo+8
Hpai1Cu2dYTaZTHIoFkcz2pMR/jlQhWF/coTAlRw5unbKKU2FI7jx3uRebdmhG7E
UGMZWKLiOR/u6dg+hSU9GPo6Seg4+YW6HIMxMJxXk60w7dyax1Ehmqu7ktjT4Y4j
u20mQ3VaE9IEsBV5oenrnQH1sB3btnfnaM4C8zPUszWcHNBck2Y3V43A0UvO2wnh
q8XXVP9Th3CxDFDzxAg5OhMcaUIKBnfFh9fGHQuAD7sQ1VnuYEBVbLIIdMCcU534
wPrnV5p1RZQ2Tkd7Jpkw9ks2v8UiMGuBeNKQNGPWgaLH0jp7FqrXHhSYxeX+i2Lh
/HaDllktSN2stJ9S/8038AnY/YdAyU7LF9AP9zQg/PXpQPcXcLHQ6vVPOxVPfgH8
LsiE5hrsaPKs+tWHB/1i/PSO5+DFO473G0IDIS/1XrddfD1kEuKI1SYWCPdAm9FU
bj76RnWvrqseGSk4M13spaAfOva7NIsv2A9A/O0qxjvQjz6JzeL1i9LxDH3pPppL
/ddXo/qEdAQQBS+JHnCjY63/4Czk87cGNmAbqhjINPkmewTtehVSG1BwqXz0he0Y
kuWak1WBnRDCPNnC5aLcj5ho0ea9fG1QyRZxv4bbKE+yKxn1ezwOL2qdvQN1Q27y
REFNkDJSjghP61eTv/wI0Pc1RGTPMm/1AeNUM7PXsrBKsAsrKV+cdkgvLxLzoiYI
n2TllGakWvxxvzgpF0IMT1kXh+orxhAlb7MJ0jffXxUoxkW5ZSxcEYT18hPU+RPq
4ckW6joy6HH+n/RNeCB7yIU/Vnxd8PIxtHtvByZfdUACvI4sJDgU3CkRgLdNkBBS
d7EQkoK0NqYMZwTCchtW7+GWbrHeNZPz9hE7pkVnHJt+ol4YTKvptq1mgakSz26v
iWK4DK8w6S0SL1BMQGucGW/q0SqarRhzzfrgc2SusP5ItvUzTC+J6FoRNdlD3UPg
NxfCAmFh/1K5xoJYmwgMWGmw7J09JSGKaIHUJUlafh85kNb7fWn+vCl2hQSOjJEI
RRlgv4dE3kMMPeGBvwftIXwXHOWeiIVUa/ai6Mbhnz8CueTX59J3LN5DfNMpKHUy
Bd0KO0h4JlizGj6cErFtQci4QJUi/+TC8wr1bGJo7ivu3GM/022zhH4uVV3AyRFf
svYPjXmCScBjytew0IXU30oM2U22IYYGYFzw4/+IsPn3F1I7IUmEqJUO8tXYElTo
ntRjiR/7JLno0FGBTAxlj828+YsxAdhIwJJqnsSiQ46ZDBrehn13QQ9S02cQqtjZ
MFnjNriCJYplhSLsq8ljVtTZSriI6o15+1vW2eQ3aU3V6nFZbFgKiMBhgWhv2WCm
zF8Gk8ZcFtcLQUZmpepPUlVfw36CeOUVq0WyOlYygRFVwHJnbzIN7EvuHW7Y/LvD
R2qHUJwn1lCbKwtqxuq7r2eSoQaoWHJJHv5BjcAGu+NHsCDbOOzKr1H3WwGP0FIj
EqHgx5UyPSXGGMCVTpwuw9GEgbWu0dw/dqEKVBZhUAfU6r7eZbpjQ7joHZC8e0kz
QRXUIjkcE9DT9vl/LTX0wFs05YmkHXsKjAjR+THMM7y5LJWCUaurRD/a6iUKMxY+
Tpz/iy7AhorcfSg4s+FjknDOftHF2yoW2z1A6rkwmDVn2W50pNMe5NbSEtHB6jpR
qw5KDAoweMzEQvxdXfe3xtdwJzeE7uQxK6NpPn5ifRqYZTUU/ZPwqkymsNWPWTDK
osJyJoojCDk/YFgECmnkrF3U9tLYM0EPGzylDAFn9riOxDSOajlhJ34EWg6Unngn
DESRyA8yeltt6ckNP5yyfKncHuvZJqpJZHVClaBToqy9BnBxsRSGUPMsOYLUJzPh
sRI1UbvgmAka2zw0T+dydgdecLHEkaq3OG2063/CS9pkYG+/UYl0wwwFbiquE6j3
hAdfGEki7lDYr7M1d+tdzoHiA8H+PSaRMXtBKiGGSmp1C3loabiDjdTwSsMZKOMc
BmsQVU65mSFxUdy3xHwm+bkzHg8kwea4RKB3N+UjYEcDJO5uEkoX1TyD2PrH3zYp
r+9FGN+yESdKuEW06q4pFTI5ZAo4YieOIUxSu/nfQ1ARAOdQNpaHN52v6AlVS+0A
uKVFFGJz/mtSWcq3Lpsm7nrt9zZb9lEddV8yrWz2yx391TmwTNu8IA7b1GlWgntB
bNAJas4esKZHbNuSZ2Syik2WM2IxYgpvICiJGXHIdg5K5QFTFhZVjQx+yW6RRe01
wXhDCZO7s65HQBiM/x3a2B0ILWB4BYkF7tGOmMuqwirY4f7dWolZrE38votqsbkP
ezyZoOPjB0MaA9w+88JBMGrOSroAo8YhnyrqwPf8qnR0BESUjdksLTOUEkIT0HFL
ggRBL34naJN1eMJmpP/zkyXf7KkqAywp0SebEy3Okxk4BchRQWSvzAKUpuS1UZkl
38Pf+maE6D35p5c/JW+049+IxBFvhH2cKYXOFAPNlD7VfmFeaLqhIVvdVaarcqtF
WMc76dwuxI1gMF43fY+REH8HqyJ/UlKUoWd4yZlue8LkJdWmVy3Ppltb37PmBIpe
CfYcTRNrMwHshUZoSjqaBt1WgCFs0uYE5VqHwUgTRQfqsx4P0CM6Ep4RwP7H6iwB
/1Wjmjsco0o6lxMwWzM+BGEXG+8n3nCn1NBMju6CdZQXRdAPXJNFqjvrTGkBLhH7
5jzjQfoFwA57fP5lw1ixLsc7S0Or/x9o20p/2L92kDPrMa35UU6+1GxXgHi0dov9
NNKgWbP+Qv/zeZaoK6m/dmLZDtNpqHMFRZskoUADymSVW1ANBrqJMWP7JGIIe92q
6CeW0zY/gTI44zIvFPpBSiU8URjZv6sFBh7P2G0NIpNUDsRIY+i0B5/skqd/qiln
/KlxtTv4hWGb3kvXppmSeMMXE3xERxeU2mFB/C7vEs3N2cRkbvB3EXj2JSRaDsxo
6xQBiLb0ZaFr4CETfsLSJiIeBlLIMqWId44MrBs/yQW6VG9Mtm0BtvmkPmYox2B6
b9R8aV4sKQDc3pUgoVZNpn5n4Zr/7j8ufHbw+cUF+qlkH7IZ2+ioW3TtqFqGv+2w
R+BHuiqIRujslsbbx0Ig3NdjQwLqYd2dAJWTVsbPKBgvydTVU7Foyrzmcq14ohRJ
FtuXzv675skD8oxP6h+UMfUvqBFkURJd+icGmdtNuneILyLGOMCHbKKdkTQgVHyZ
mR4VVO8n15wj55wGaOptmyKFsTUZapOZRkltpRbeeL6v8U5XwtM5N3v0jm1sDUym
LVjGFwsZFQB7mKoW8zfKzxznoNulttbBt76WJvOYfrsL/3gIvTXVXvn/ZDUaSMHd
YhEm7+IMCHHtGxML+JaRmV3LE6C0OsAuSV4JNe1ZeWfTgbhi2GnMsFviGgTJvK9C
zmA7lpqkDlS5jMlAQWHfXnnbVMxrRseVW4oIBwnXkgb25GSdbeEJcyHjcleihHAl
LCh/lCEsFPP0pmX6MUnPPSeS7mnDltYD9UsTQSVxScT1PRLwY2FiYJ0X7JBJ5PHQ
pJaPJE5yJi31mQcaiJEGIkeas7bAF6cp+nqkKpOlNx8jCQv6KJd/NxrEhvWK4LQm
TPR3XdzP3YPfp7in7/UFWcmksbKcbo9kotcaqr4PnhCOOC8dkAwEpqbp6FxizACg
5xJOmDWVeJJF34ec5sdjDV1JiJKroT//LxoDR3SAXwRHwnwUqZmBdEk1MVrR7Twx
VV8HjtHWBmM/ksU7K+gPUyk0twZ7hMeW6sGqgi6TfWyEx9VL6/Hu+r/U5nCmyFB4
fu9e9QRLNbtLQwI89kmTbbCjI1uVlyUxTNP6NXzdpOJBxr3UvhpvRVk/SuRf4TEo
azqWaXh0MdY/YR1oWF+xnUU5Y/vglSOQymAKCj2uWhL4f1bP/Y27SsyNdrb8Uf2i
8T1msOYP0iDYhYvOl8/HVTk1DmYUXKiQYCKN0iD0ywvXxDYn4CMVLvj+BWYoNHNT
QrXbBUKeQBr5Ug3nK9GOGCDlmiJqVEPcj+k8EnDZpreu4r7/Zkr80MJvybPK7SGu
vcFKXeTganO5vbl02CYXiDVIdSJXgCWy7vYL76iRKjl61ThwBdxZYS+8TdSDiDAj
3su03I70uFyY7f0WN4TJz5fIm2MPmY9AazdP2Ivsq/mO2jmfXgm37skRqle51WNJ
1O3ZKkLsEnmWElGnPYMxJphGYRa0Am5c4w3VXWWQDk4BvY9hKBGZEzriPfmJ6cyN
S/qOK4/FRVRmRlaXaFjEhllBQDVkKBV8OBY6OSV9OMpmkdx+RpVG5wurcQKIl+Ar
JaTMe8itEt55tIxSMaYgPMb0+YOrXAxrxJs7YMhpfh6fL0qvSZm65NML2SBN/PZN
Ptw3gWg3DTtHaUeaX9bSqtYkrjuMVu7xNgoAdMWtMb7/7Z8pLQsgwNb032CbugeW
ajesSDC+8xWYrx/U6x9R36KmFrGf473/CaVrDfa7i88xGK8umQdNl/PDYONTLP4C
gjorOkBOVCL2ZiccJMKJZpDoKNDUvmbjJh+2VR1S/0pMMIL1mNXD9MdSV3o+KFlQ
3N9+7w40oeePa11L1GQT7dQ/UjbbbiRfOqw+sRkR7nkPB24h27k1LCgfjkxEaSFZ
htc/gph5ZOi00Rre0BRGh7ED3KlGxHFuxWYPb6osASKNlLyOoikivT5BH5mGpT9n
uMNF61pd6MjzbaOgPQ/8j12Yy1BDDNSk1zFZnys2HLpPDmk+eLrPeL24dM+CIRtt
i2OJolgLssqb+gD0Mo8dC/U4/zBUpro1FmKYgt+vV7SBeGqrp7/vKGmdvs++Pzpm
eeU/0Vy5nxaUBRAHLsP/yRbegcI/FoVtNSnqdQ1i626ZP73CAoTw3qvHFq5TXYHN
FeHeW3K1iR3TYyMeWMlnRqurFRN3kbqUpq+X5FAWL9V/920tUoR2Lh135oXC1D3z
gaqQj+r70xqF6pCTL2ySmm69gwS4ShR/+fXLhH+7VjjCEiZOEEB/i7nuIS7Q/GU/
twJGyhXaHX3tw/J9JKluhSxYmbE0o/0h/j+i8bx5htMjoEo+fLT7kWhofQir2x6P
6WaPO/yCTrRhQWe05GIuJ5386MRhg6pgM098LIJc44OiFWwuIU8F9MYOKh5Wm5AV
9qA65w40pox5n6UbqU4aWlgNxC22lX0+qcg2JIU5mAfsDrsvWn/H83vAqx8Yfza5
sN9sP+VwjECILTh83hJahBLODF64tbtQxa3brymq3kwW63VVgLQkccU/WgI1xXi2
8XOa5II0exNTms1OF6N/k+BWhDbuatZ7+i+GGZqVzZGlytULfBauG/bqQXPThcCI
pXcXfYB/JHtgmWrW0F4fOyR38h81Np+A1ms/e6L+2Frqq6+ktKd2ADA978v8j/Mx
vZDCyxbplon5tISRymiNVdnsKtmQNQRxm1Sj5PUPzSHR/9i06FrGvsgWKhLagF7Z
ppTBdZmwB7DqJwcw6oYKtSnTKjMKjAuUnF9hWlIWneywBQ8vYELdHhz0gRxLR6/Y
HYlI5raYHiFOx+Nx91fCK3mh1Vbi37P3tQpsaMwiixE8shwGhkfHlDT0+4t1o+Hn
+oDxy6x9FYRPHfLYjbYYT7s64l4juVVH4vAxx9qdWDGlQ8UpH+GRNLb9NjwbcCSc
EinAjfsO+MnTCYPfnvrJKvXglbNalZoTcwJdR4Fzu88ulOxt//oixUMTbx1Q5i8w
VfkaddfgLaovzYlAv+8FwgvFsZqOgAlwLbqL9tEGUBBWawRazwdRPcqanNqmD8OX
BGKoYV3w0++7ZBplrtFlP1EGOVUHEWjN3C+Awbh9CVe63KE+YPgNAVRvhk+qQlwZ
Ai9BI/K+UHrcqqJcmmnBIF3HygIXxkZ10ros2DfwfBZ3C1V+K/o/MWYIeyH1j91j
zqi72vxUS0pqL5ooYARNXQcA0O3L2JuHZBfmERArVAU/zL8MkiwSOaueKXdJlCmr
72zBeiO8+4Q7xwqH74chsuYT0QH+98qg8gNREQfuECze/bLvL6i+Y2X4l0V/rYtx
Vzj4SmWp1HMl/97JpbzVlQa62OsFHTV+zhyydh0+1ntbZ9xY8vXSYberS06k2L5J
1PLIv0Harlloz34B2jJsAQ5FBOzVQlPKn8PMxgHDKOyXDlaNp3EFtGHLmRkIiYwO
Dsqeg64nkm9Wrk/xANnUz4yDC/S3yH/vl+yJ++rh4QGGV18dC4GrXXsWlvpWgPbq
PTUmVqbZz0r7usJLv74l2kEQCtUMwukP1FPBBCAp/5loiZYn3mfvToYS6W8LkwoE
CtYPLiqyviXmhasgXLvB+1n1Mu4XvDeZKEi4TakYrpLdioZ+fYCshXFfkBH4mxfg
vKZU3eOzb02HZOOTUvGMjczGj6PkthqvJGElyBG4E65h2WafDrkZB8UMRuWfr5s3
DZIcQDBLZJ046CqMC7Fvag/QWs5Sx9nwPUjCZpv0hqFd71jKMWKaYVeskldMykEo
vzBc2aTBzt5HCPpmW3O7EQNRUTkFXypjpszeoE8Xo9FxQOIgy/MFshrZ3dUpSq2j
KvHKgSAv/1jtwAWlut4Mw8mC2frgdjZwglaJ/W42HDH1p7XlbGfLaTVlrhGDUdPG
67XzsVftU0Rr3oGA2GsLPVCLr469vfaVUlK/9S6spviLC+w8MXb8SLaBvudxnXgd
RKlLZh3jHQaNSSPKeo9efo89nLnt5T6S6fZCd76qqseBtZIUGHJJjcPO+HjnpbBI
DEpazGSTaTH3QGTjSGKvIyQf/AuAw9jeJ4DteNG2quZvEGhz9uvjv4lvE51/sBVD
0Yg/FQ5EJVFlNhebemWo6e1tRU5sdkzim7orTqu4Yc/7hUpaiakfRt0Ly3rPCYm7
xqyN0KztktQt1YNdMaAv+KU/CpZE0dOIiS4y5/DCRCHp0g9V2AEqQwcx5JGo5rad
agIkRL32k0G6mjg7h7K7UvDcLmrwkV8V0DXxMf0RwfKi8pJlkJiiCtikD8TgGhJ+
HvdE8oYNtTLgE6/NZWZAdcSTQpbzT+78jXRAkq0E9NKvDFuah4H5Bh29UvlfdH0C
gvF0osHwz0o1SW5P0IhBHHFUjk1SglMD+bPOHhloDOcXG9q6ZO3aB03ZGjohJO2n
k2y83dsGUN7kQWe/bgzK9vmu2odqS4AJh+X18/Yygz1KqbLcwDdWt3r+PPCxowU1
xFwZqSUOF5eTPfKhLiWGRbROccHBtb178vQBI6S4gx5tJ8t+dgtvgytEBhLGgw1M
ckB+FKcTkzxNbF67KN3g38LpRJc3pONSRznCM5/RGuwIJrq7RKWPvxM3wgMEFPtq
N8reEI2ENZUJ47jU/CeUBivpfz7Y8yhUV66QDPAJmhvF4p+qvKVjIUutLpDBRmvJ
tYBE2Gh5l5ShqZNCw3w4F0gKB2YCtWt3LkXgg96fdW/Jp/8YyuR6jzcptq8/yCat
s2OLo3PlOekvQwK7e7CoCbAZuNJEtKgSuVg+gdORIlzd5xcFIHYP1uWLaGBlKJBL
qI3YyOpPFFIihKt6PCtdAozSAYsqSuJAE9HlrFAao34PNDEN8X+Dn0mVgZcuEwsU
GcxR5eI+jxX6CpW/SpeNF+UWKkWMa8Z8cVtpe9l76mPrGTB9WjuBhQteRoIUprdQ
WVgm/bZfZKVO8AaqgnSHyL506Wjep/8/ZTc2CbHt2yCk0oJDX5y/gJJutV88P4KX
4Rl+PleFrYj8p9mUc9/56xuHGWL75fj3VxWuifE8wm4qvxQtc0tUieEVCFn/b5oV
SSFST5qtjeHMWCGevH0LO5PIm2di2A/J9iF6fQcX8qI6GlNTVZF6hbfORLvnZJXR
NOUNA1vt0mv1gBFmx00z6jAxl2ztpnkzbBX0FK+2mbTIVkwmsMS8Fepc3YQHhFWC
aXGO6GdzjZ4hU/wQ5Spb02O4Ejp3z0ah9p+wTEyUw+7rrfpyqjO64wVG2e5/7ez8
Bu+zoKmfm3wX//t3BAD76sMb6v6u9Xf+BLGzXMohN6gaiyeLOsYsjCZ1D5yGNyKo
FP0ar4wQ/ex83kMiImzFGr1EJNdHyC0szHV1iTbr8yWh4/9JVy3FjqZ7FUsAJFld
n/V0ljI9gbDCyPn+7NF8oxC0r+g6e5N/YZkVTyaZamkQesJQbG2hqF+QEdE1EUz3
1BAzm63mlFVfbQyHVGf3MiEKvi9hRPc9rz+H1/f0Rqzphs9usgAbP0GYbQMDymh0
C5NamHPhnaTCIxnl4s5ZORDSjmOZEWaq+s0xBSoAaTN3r6CDzDZe6fTpkQsBvFAS
VrLWigfqehC4HHQ0ys3BnCauXq1WNE2m6JZjKdJi6IuG71fkGoZsAL3aPJv46ljj
dPgorHLSfyBhKglVYuH/GaYPnH29CxulpYnvlplfWgH8zVfTX7wr9f7KGSlSuBne
28lgIRjti0GldfL2Gd199nrJA4nxk/vcr6ONJIyKABWgWz4XtBvGP9iVDlu749JA
sGCS3v0mjUFI1R+LcAw8oTDTEBD/2UNPesVqpU1GOJJWUhNjFzQ2TCFrET1k2BXc
26XvTuYdmcQS4x/RElpeB40QM68P4+exN1ugB+cLe0bbxbtlmaRdbasiuWOc6AWw
T/x+Iyw4yqtxl/Z7ZQgs1Wt7iICXlJFUBZM3jXwPpWo5XmGxRCQzV88P7WCBjnxG
/jtmRFRGcQkp6KOrpCjohVkhnbtrzt+Nl8fnfHo5f3DioyeMs0Q28lXOTtbf4qqV
GE+Yv7jTGkMOgOBp0eQLEUJaknDXOPtGgd0iCHTWN01RveUd8/x6bzWu8VF9hm9k
vaXU5RGIi4dbQ+iTxjbcrwfsd7g3qYWLESd9LMP3OsQ04fYH1q55DDAQHI69rrlq
smqeJ/2VU/EML0ijQO2LOzaaSinpdX2ZntqVKpIZUHhSfV8Dg7BqHzjlesicLD6F
mKZ3LrD754RzguNSkvpxxyF2kCUr4lFm15x4TfylTASaMr3Tiiv3uLApwqHizknW
6SbkK6PtFnlzN94Grue6kOMouW2iZeJjO+xT6bMspDUQg+qXqmnXSxIHvTn/x6zQ
jDvuwVhz5oZap1odcHFdjJKvJIL6SDGgHNrsRukCGsIfzYYuMyKvRzTSpPgQcMDF
Lw8nJ6Tv/eqeIRJmedLZVHGHcroQm0JSlI6J//WFSKOZ1RWLvn2WfHOevMpdUjaS
DjgII/Dt7cOsaQdDz0BY960+p6SdBKlW2TLznS8Cw+TUq0kvN2HV/saSOrPVawHB
HZg5yclwXSrTeSNl1Z22p+rWsscquEScvMDHvxpTsjiDOUyNgL6lG6CEFSqAcwMP
peGXpS5qcmePbXUCgmyuYRIOnZ07XenWTdq3OQcH0TwRxi50sF5zOxTtF5iBBRpT
eSJZp6WFIQdh7Vr/5szBiravezxAEvijOmMjfXHnQBerqVS4UFm5sxlIYLkoXptc
o5xSSwD7OxGE0VsaXElVmWu3Iyfj+dhl+O/WvKCJUJLbAcVS+JFS8HzCzneR/DRA
/ly+LccWglkycbmZCdeejGoUKcLsUzHebeayG6yldpKAKDuk7AFmVl1taAb6Hz6D
LuGFM/OcvbMELmfE+TH4sCWkYmZOZH0BUM6O64xjx5LxbMSSWNDAYiGA5uhbY1wF
qqaiB95O0HCRhbvn9XV5wUsxsR7JYrNAfJan+CRsGDPYK5rnHjIPXrdqJZQc//q0
dN9y0tNLyjKqGnqm/nuKqo18fi8ULXFxzxl77QBlJC+MRW/OAP/ZjavQdDpCwYIy
SyA3jnOTQZ3oxCNMH1pUbQplWeFoyRHn6c55pVTT+nq/3XSvbf92XNgpztdYYJ1Y
z4DCszJ4GvDX+0nS2D/Zg+EqxcqfNgh/ROTxfQ0c2wzfIqh09QH/x4+dNeSSq++l
JxclOQiL6he1z9P3D8DgMbDllTPQVyMMr2lhviFWx/pIlaSuiUlz6BwH63L18FLq
4ED3Qd5G6+4qIXYCQ9JHkk4sVLbkGwIpHU05MEGQtrvGYjTpHCKiaOZjzzv7uOUY
XBO/DX7A3l9g2fm/9whBS/UPlo+Sc7bPWxEZ8TC0y52jGqFH18n//l10mz4ZZ29q
TFek2Ex28jWRjkrnlCu+CKbPecC6dFNhiJL5x+H21VzPPdtIZ/XZG8ret+0cDxKI
wyN+HkEFcO0ORCntO5hned7tyhg6Qxtq4HaKXmX/c/+zMeHiPlcb0a7aloSZ0wIG
r5VQPQwwdaTmalEJmqTON+B0TKeo/YoWrGgTpTwI8yroLDXedQEmM3hYpleCAIWa
2nBZRkkpJjUS49zmIvqSyCowKm+WLMetd1gaVi65at4IP89cFzCakoo0PIQpeJLi
E1YGO3kyuBGb3VRae9aljo4QEEUi2We196DiEkGsTYMiy2g9mHusS+sOV3NWAbsd
of6LCPDa72dcPh/NR38ROH0hBFV3x/xH1EsK0jfHRHCkCXX/O06lUPeMQpthdvTu
SX4GzI0TviGqTyj5Jzt2sMifu6Mvmd6X5EKc9q5kOHBlE7otnZ75YdImC4fR76Iv
fqLeh5pxNVT12YxveObctC+sMojin/0ooQejicUUsY9okUzH0d+lx8dt84IqsXEH
K2LM2XGA1pYiZgLvTAy8s3ZECi3WQuzGquV+qFxNj6fJcovQHnaO7b7YEB+51zy+
Hj7y7Ige27+QjUF0PXZxXXWHV+xCj8a3S8HkMZDEXMIxvARngMxYFVIwOb+hT0Tv
eH11/Y3taQ2YMUwDMlYb+EZjsoeQ9OsJ246M0M8FtuFvLg5EdvesdHs9HXlS1v3x
u7UgeTJL1O4fdtz3paRH2R5PilXrw7f2qcnumPFUuLkPbQSOR2u8g5GxmuRTxe+7
uZ9MTTNzVkL8j5sjp3ki6y/XcJmm/7qIhsSuMVOEIwHHPQ3gUrh0IYX49HGkY1Vm
Mb7PMmPehEWmFnHoy2wxAHpRbnkPee38CZDvVfs/u9V1kF0E1FX7RQbkK18vqgyi
WNPWHYzeM/YRG4gxNif86yUPWGHpXOvoSIO+p9MjCxKwA4UbKfojzAMd2eNmscJW
+fQVH7/ElOdpBqCDrDNMLbslGHFq8DoyZHIr3RodvvM2iVaoxbj2CtHCnIFQYz0+
uof+MwtK4HO40EO5YnCwSOgyX1cwzGV/eClvTlGA5Hvs0v2foUrVFIkjkTnuWVE9
yVA7zd/qWnBMvspxzcgI6g6LZ1pNo46LjkxyGXKceSa2+zjydIkIveZoIKeIQcgq
FKDEZkKCEzzkydEiyXnlQCxxrp55svpasduNDhXa5ZYWm3q7aD4MFze7/bmbhqal
sAWP8gE2p2cwdCSDG4zbbeiOwNJ16FLA//WDGSHoFUnm+OTgJEDPYVs3QoIrVkzy
YVBZX/tVsRzTj/ynFjkyy2PIMI1WQsRrwWJmqkQBQHPAKVrG68/e3KJ5QhMCRNl7
piZJnmW9RAQORAYRzOu+zODbeV2sWJsHXNPZBnF5IxOa9jC0MEqLyqWSyQ954kFk
jYO1bwGmjvif8kcvZAl4ir5ec8q6zig9BvRZI1hpU0IXWjCPpu0kIIsGYq9FrDqg
C66ptHl1inzrMSt2WLN3vhUKZ+OYnaTFzImRZnfSGYVEwrwqtN/1mF+knqlo7AVM
N+NLt6WaeYB9rttfrwY5DdDkrXroEQRMeFysHckBegDCXHVdzknpnlPAle1ioamc
UeXGnk85Z39BfX/b3XvYvwjXiRfs6/+MGNLAt0/uPNlDrwCvxSInn0i74rU5v5hc
/Mq+XcySTuHO715G5kr9TMCnTboJwo4mukpgQEzWD+Le6AfprBUzayaYnPKT/pt3
kPVhV6VZoQm49xYcMEDGfnGMQygupetRMow5vdpxUZkhHNT8bvq0rAD75fvydjit
ZZ2FUOJYLlJhiMrKC0hDOBDyJqtmWtu4aTrGfpmTEN9Mui+1sGRlkyjAWEawqctf
P/yRIkA73MR2yrAdtqRfzjLuHeyge0JHNC6e7ZgDfLPvlKtfyKxblbbZtNnAzOvD
dVhOfEzyAfmxGdQ9YMKi+1aYT1wGEEBVWSXnPzBxhqBa5NgWoFWbFwA/f4QI/+o4
0q3WxOGvXbhV+sWf/mAkZSiEOFzDgWXf0z8gHoB0KVnD/3PGUf5nB3NwTgVDkZjn
pyR9y3mJj/4mi/1hYOkyI2L0O7RZXyxLFralJHIQ4l77T7E+9iImL0WidiE2SGsz
+Sqzs+zLMlD7LMURdJTndib9SDqGdr3VtXL1i/qdKA7fnwHqkVn4shaLJ1EIeG3V
whMwbY64IUQbjjLcLpBBCWgizclM2v5TW1PskJLlY5PF8rXpczVW8buA0+7BozKa
26Q10jRisKoV7tGc+pn8Lm80Y1h66Lvg+4GJAEi88nZcEB0kMndNjUDoGoobrQqX
gb/zd8p0wVKZXsLwB7PxaTyXTjs7ZOT7aYdlhYsU4Fk0H5gt4Ln2PojkMXT7JGZe
7xMm8PkPFQ9WA6jOaLZ1XoUv2PLnVLxgrP+deO9mkT5LbPh+234s/MevhPlt2ywh
PUqXu7UOyN342As6tysDExBq9iXAu/z0kWXrtH1EYFGvHncDotYhzl8q+0+zNwKK
/eXehPC1So8NuYYH6GaC1bEH6cNqIDg0KHx7dnXWaVVaS7scw+QMrzcAB4B1K2xl
HKr7pYSMLz2m4abG8u1S/MXKCtMA4SAjfvhr4sXuCS+CWLVfgWpSrsf1hl7+zJhh
KmSncFOLd4Mm1p3n0VloRYDC7m0iYZllJRQkBvOlQDnsz5719jJ68f3i4dzZze9p
OzhMmtX3FQtjRcQlOnDYiT7XoxS/SgtcPcSNgjdYQcui3Pjxj1nFUnY0UcJ7IRgH
TKZqPrQhgOBe9iPvGHxm9aL1QZjZGxw0Uq0MIfIAztyJDq32UywNYa5vZU9spSST
iIKEacjTI6lPTSztcghzbDm0r3YXu2hbofeWSAbYSApply+eQG6C/ZdnHJD23MZC
jF30qckhCO+mQ/0yNIfP1ieiFg5mnBEOvwgy24K/jIhL1ref5hwM7RiWzHbSjGxm
gnEHz5WxpvFEoAV0x6goXr1C2nlzvCaCi5jbOm0J2LojxV9/iqBxox2ps2brb8i2
yLv9f77QFXd3Lno7r9KQI/jHK8E6vJCvOYvNI2Gp0JtXNb7T33TZ3dYbui6iAnhv
q2ZZkkdVwpprKkoU2GNx2F/tkJAZsrNlIUsFbaenWeJ6V0NsLGpx5KHuaq5UNChb
qSy1LWnfWfddtc2LUwD2BYdpmkutJtUkwCJ6nAaXalP8YgiPfYYdAT4B42uwPPxd
cVOMkNhPh5n/GqJg6daFa7EeNUUu8R6yXJsdK8rJBO4l6qVkRuZWsrYj1Qcg7gc3
mhas75Eallwfy+t/K/PLXnDUxMPs/YWZ7ggx8VcNip6LkS1lz63RDrOx68ueBDSb
HutOAnnrnMdwWYCkFGE9nLmNuGjr2W4DH4E6phduueGSTdSlJv0ikLLLK6gZum3X
X63E2bLWoAnYUQdbVXu26aOlLRspthyeMvKxEBNvKLPOHYYITZw+o0qz2ObbnPNW
NL0yGuYRMGjMz0PxyJAeTLHkW06tQecGWFp1gBAKoBArBIHDE8vgPgBgI2Og0AX9
8vRXhf/9GjPooKreicuAF1gl4V4rLi5JTMk5hA2VCK+UmkWya+n/JfGlOfrNjkLv
Qi7lx0XIoKlh/3gbRMgVb7hy7tZGLURHq7V7alG1f1QyC0D0p9BwWUGekz+Z9T2C
zd08f9+KWiBx0Yc8Gd/Sj4UggkJi1ckXHkTHC5Su0Si22OkmpCsydy8It/QEa+Mk
qBjHGIQNfCMwNBo5kvzl9VzFZTlFUPn8LQCR1P4dJUzd1PC0lFx/uM3nk9byE01K
E2f54ZSwOkt7PvC5mMIqK/V7nKUUcVrOofBxDOvNCW9uZsp4QWwZYdTZkTO3u0E9
QZA1IOj0noMC0SrSqWoTR2RuS9d18Q3EgNvkAOJDyBs0jdC4vfTQtKUB4iAHGGHK
jIP1VF0GtGV+X+GVKnk5lrMYiwnpl04g57PbQluR2fgr/1ZN2Q0mZxW7B4lfoOkZ
/C6TRPYGY92ZB5TOUUw0n/kVCkcXUfnerFVpOnnH1LP26jaIuiNGm56Zd2O/7sCL
xdHkyuoa1nICnvqHbyBDuu1qUChYXkqtUeLKWAPLpSIO8OGi/uEUtn1zeY3NGevP
fgmtRHQm7YCE0zVGreP6stmkQ7SV4QMPA2Gos70gI4OyZgJPUaHie7qGZap6qksK
kA+5aAfl7Js5YB8HuUn+iyzpO39UgP8OQEG7C1t25ldE4pIRTS9fJv5DoES4Bch7
YKGQfp6evWpO5OBlBFSC0J7R1/RRJD9iI+GueGe4rmLCJz9pjbWijvVpoRg0G5H6
1BSmHLG4TKeVdOlmCAAj9EVwm/o86qRjh68WQ2OOE6cPpaMzozhtVoPhPtSNPEqv
8H1v6rDpQSKN319+62V6bTjO2XRAE1lt2JyrFf4+2k52hxP7Z2fiwiT4klK4OhuY
fBYnsA7Mgff6WqyIM8f1dRJwNQEYhrLhIgcYOu6KRDiUwEunphlq0c2AVNTxx0Ey
gkwN5HcGCVwF+iHZGdKYxooXN375Ahn77tWp3QkillecZXvO4IWxD0M/khQCwAIZ
HXDq3GQ1QpUWXMg8MHCajtvFPn61CgqLjKY7nDKOmoS323vNfi5WFNPBDlmxnQr9
6GQgE8G+RCIosXsSmDpN7rMOImi/78ZSZPAun0QjTxn5SQh9kIQWXSrrn4opKgmw
7o6/MDNBJVogdQwtaiyoEiaPFrLYPzdH23Xz27WeOo5Vh3RPbMcYjKdvCD92MIY6
JUkt+mr4pYRPS+JzZOUBblYoRy/xFkJWY5Nvr2gha3JPaLYPDiKJUW2I2sXnFTT1
7ikMCPf7+elz5UsmK5ZQdtXphtOrfHWYVw7tYc42If9iZD6v0BK3WRzbMcl+EA/U
KR4Lp6U+Tsd4hIQCIi627VLoE6GpC2Wo18kCCPZ9WiREw3DWH3wkgIiCu7uF5kSo
lZcdprsQ7bhTWvoiOtKTwqIhQL5fZ2FIqYBwzBytWIri5fnao/KC3UtlO2KyoOlW
K9sHvR+F17tZKby+T/if9y9xcd0eTdCX8QZDB/EfTWK9DXZZXXDQozyzLn24kRdX
PZfY0v0hMTaWfV5+5f9BWwSaEzAkhk47Z8wfwXtWbxz04MLIb+JVxAO4VVEFynp7
kextwcN0zxOotVYqygd6pnkQG0BgeNiHC+rzopbFAsWlZNH1jHEWSc3wJzZIAXIp
V57zPQEtHg4bbg8Fc/CrVoDSL4FGGKewo2IvCYhZVveQpGegIvmkCk2itXVaPb2d
5ddVllxRdyvijTckbKMvkjGavxrTBGswM7n6YiDOAIw+6Ctp3i4739Tnosx84rP0
T9n0q/M1wRLg6EQM67DHwc0EyYU4H7s57vrfB2BnpvnMgTPSuISgPHGLtU2eDgUN
dcCFWO6qCD9BvrMTj/e6ygaaYxhfZooqj8tD+wtOTkKlBRfP8JEm/FJ1IORz2NaA
9zI3wbH1JcH0PJy9cYFjdK4mXNMYkZhTcqNTMn/aGATAdCuhUnJ5VVwADAMMMgel
JctwUOgERCh6/Hp83JyN5jgd4uQmMQavU5E7oyY5DbdRWn9KnddiyC14KF34jRqt
ppiCSzqRnnEOvEOIHvuo6SjTpkiwFCl1AgJrZpCDNGveHTVtLOfEJ+N65oc7bdGy
72LmktOZSY6pv2yPLCoCPdXYfeY0Ht0oy97cQzr7UfMSGRrN3zyRs4anAhfmqbk6
sJxeWKlAv4oP5xtXOJRpH0eoxWkM25FcjKCZ4kZRP7VK/xFl4hK+n/JldvXWyRQS
6e6FC9sMQPDsvFCPiC8vhYC7Ysvj9+sx/efNsCthC/6qIADBsgdKLVoyXDmX+JXw
xW6C7nV1ufQ/lSbOQQ91vKhALoelAaaeujEiE3GwSVuEUBUP8vmngOh5wanZ/Puj
jx2PUnNCr3yxo+qddoOKCI2sk9W3bvR3fd0WzCGj3QZgFLJtDmKQi/f8FQlMfgM7
AYA1RZTC5lXnZDkKySwSJF2Ns+8TvPCC2V51IYqG+GI+Kob8qOochFG9/J9iU0is
hIJ39+/UuwwWsLbRxFJOviOJAdhrX6hpa1V8yxHKDI8hyJV8LeS0NBDf+9NrfhdB
6doc7wRljZ3j+zd3AlPv6g4OdTPu/WNE+hRSmHhz3IOj0ThnyHJARF45ut/K32Mt
vgi3HS2HOArQAs716Q5uO1Vb+qMfTNuoHcfv+pyYOR+uhvNcGxw6uX9c73mUe8q+
Uw/Fgkrw5UPgpasJVJj7e+cDkvDWq2S/9PlJhFgZXXJM60KaYAp0ESaefLbNa34l
klUjhqg/CXmjmbbea19MM4BkzQ7m0N/nKebWjHJhTW4Zoi+JMnIeN3h7pDWsFEHW
N1ei7Nk/lzSULaPx4d4HGkVEDwL6YKWCLIGyG4JtKdCqDRYU51Ogv1WLGTrEMobO
BeboBbVdOG7oje8Kqq15/9VKCxl/LnZnmjzdeFqUZ2RhxndvfuRqKkbMnlB8cZKo
kPOo19zbZn4Svr2cyOqIYD+3/5k5Z7GspE8a24NuYTeQ4wOs3kd+sfgiFasN3lds
NE4O/7zKmBmATJvE6vg81DBvGB1z+cMaodR0chVVTsEnzUixf6RdW7LuDkioJSF9
a741ugllG7BxiXyCDbo0z/+o/Oeo+W3bszCdqOcaP/+HoH0c+2wo4Iw5XWd0pGjz
HtQcHiUiBU16xP/3lztQbOTsxBR+T2n29wLAvPtYZA/XVF8RJsCp/4rnxJMNYapD
FRiTeBaczhZTj2njupKJlcp/RZ/vNYSDWtCT6iZFSIyRKu7rKpkFDK7nLhi2OGvV
GZY4lCyzw6cAbDhgvQtIXQDFVuL9Da7m0Ys3xCAl0lY72NwwmRzxVueS5PmRmT+d
r9Hv0VlBlVYZIOXzx8W5lZulMsbBjFTuXMpLHyWPFWAv5T+yb8mUaNDt03Z1XHYF
wiG8U/wjsPOXc/MWu0dGCRpGqgUpqR4nJzMDeXDsfMMOOwUvi54sa7MfG3s2OSwp
oMKVTd0MIU6JFK2q74BtU5nEb2amMewiAgNVQTt+tQvSgon1MNDToT/QNIbNHRix
/tfmqDQt7jz61LDeDCWPDxZMPTHD0PvugrJohj3d/EDY2jYCxvJu0PMAddANE8Tz
CFJHBuJAr61y5gwgUCe3p+hNw5sDqlakmdblGotpm9O4jBT/BdUF/Vs1i62CLsre
bCZC9lEXYWM+beBAifuqyQgLoM33gMrUO5zr9BNW+bEEULZkZqjiQa859MSkOhdB
p91EHCLIVH4PY36XGTJgCSGG8LD7oCqfylZN3o8WABshUdca5EIcE+HS+1w/8ypb
MOuNUz/ctBQ0irLdu3JyU3g1i1uuqt+0vNWCiBakyHhAxR3o2EvMpHEAVo4Hkwna
sZtLcNiGmbo+s/Ur8J+edsv68iYMTqH4WEAmIATEuIToVB20CzKUanQzrMUE4g99
lnSXnBC08XXrEK6nLlPRd5MxjsDBZLRZjI0p4opjMNjgQr0VU2mJAiqQsg0EQvzQ
yK1LZ5rpg0jb9wGyhosPXcyvS4f/LLu1O2mNWQonhSsqLV+u74J4GVi/1TE0a/9n
FPw7XmoatC5uI5wm8g4g9GKjzbowHQD9ML/F5UMMJ8r/AazOlmn4chrLLFLkJ3RU
f8LB9jeKk1YmbvZW93bQMy5Twc1Xmk5Ql4ugE6rrLPS7YfjwRRMEBfyEeHL1AkWw
/YtHHm3dx0Jnvrmnhn7HxvoxPiS76VtQEKY7v+5HgwzpysxJc2ZMUVwVOynN8FZe
lSmV0x872GoKCWQkI+ycvqLMVx43GJD92JQxCqk56QRpFc8CsaXmkBzpFaN4/9K3
OBbRoppXl1KGi7WkA7B6y0FTc100hrDwUstwKE90nyamJ4v2/IZDXxQaxvUxFest
zWLf67XH2T9XTsalflRIUnjAMxfnO1eMB8TIrYOw7aEGnYRyEsrjhd/r4J9arust
BZzheVbNA+xBaPp2WvAiEdNIzd5yo0CYVgn1thwiND6LSAbmdn3KEoPKlroeMnuQ
xk6joCyJku0nSWJ1AwEzDPWaOxHUZwDERZr85LKZP6bBjG2N5lmcEHsysuRttyG+
SfF1Sd7DxqXPkN05EmnXRVx12vt92tPx4afVH/n9OfAir3r0YuZtzmEdUrFwvRNP
0rakjfGC/fbz+8qDEalk++uT/rSzGW34EtmQdzZ+ku7qtFzSj0aRB3fQ9uGaSVf0
4ttgv/5hKsLRLLzPimeXmv8AUyOdi/qPibyG37k4+CaEdTLZO0ZXwq36v3xJJ/TO
CIT7QeXbxxX8wtq7QmpoVXWmAzvIF8Plo7/CN1OfPozvXdhLczjXih1b/hSr8dad
BVMJ1yv9ZfOoE1IgNFXTE2XnCXJCjnqrrghykXRWIyyne6uxq9O2nHhPWqbX7h6w
0JVFChguP7oiyeUe+HqoRRZpiLjBV/wKaHmB3GRJ0G+RUFlQHg9Uq3CVmS+bXNbP
GEcHQu1KCjeohVRLW4YaftNM9q9NSxA2VwKNN4NRn291el0/qn91M6j9xHfMEFdc
q4chp5EP8/Ifd1SAhsx02co/J0T0sTp+OULi9kuMdRxPTCno5BzO8nJHtxGrUBgc
mSFaanM508QF752RrAPfvsCVdZdg2sj9LKiamhCad95lrvnq7KMHh0NfDJ36da1Y
Aec5kFKNbTCbjelpfUvuiCn2RjkOVR4zALoUJ4Er2aCGftk16GYDqYkVzXTszsJ9
94Sveq4BZ5fALzdwaG4rTtjW1Jn5pfqJNHd3iCewATHwd9QztSuPQfQPk5WtAkXp
6S9a7M7n6mEd4veVC2F2td0I6IOzGOdOie3q0AIRywF49MOE9yUqT45pFAVgoScY
cDjSmL4r5rx9V+iFEx5bBGk3E2ZKU/5o2nhJQ3UWwMNkZWj7lB+gyL5w7tozyLLz
SpJj2vJ1dQ/hxwvvyTh2NKSuxa/vhCo5vMwwv19Ie1Xu+qiaWuKMJ7ZaBeUeQXie
fWPU0kZH+at1sCfqDq1pP6+cf7DFaFZI5MdXvWhkiWlkH35H4rHbtk3HwHlfjDlv
NL6LqOZiyGtznIUIXkp2Jh99lKSMxaVxotGHAPKfbDp8dX6n40a66SJG7uJW/fJ/
yi1MpZWohghkhVK6o1B3nnHtIxbJ+Q9+1udXs22vFLoYyL8yA9aHUMgHGjo4+5iI
2CMiEFlyeTMN23fc4A2hfZOFQT3GXo92zcAv5fCAip+RTxAmzXcKXvo0YceVcfjV
EFHdaGV6d3xZ3icuryrSnfw+osy8J6mK8z2j1rb+p93TYzwxXS4iOR0F2wsfOc2v
A/TMUZ2JWM1PoOcnI4A3zZipnMkWD8PzqoVPaDqUiEvcLR+hRySAVTpoLQkqw9Za
2J4Xp2UGzb68LgF50jP9FrbCxSQBqf36r16Bh9RENrcvm8vwAN8+0g5swuHoLMIO
lUmhoxfk2Sa24G1TDbKVZKumd8ssTz9O1eKy581Y2IW1WxXmavFgY78Y7qrVHXFd
Y7uqpFrx9MNg2f52LASSt4RhPbo1O9OGLhg9kA5lVQ417LJE63vYOg/lgW1i0gkP
0pgDlRyQBAMc0V8xMJ+9eYvpoFJkEk4hVXkGeN3U3+BeSVibzcksfLyE7lwpTKRs
nsM2kRjf2OV+/8i3NK7n/7j6xhk1xeFFKxAVD/tsEn0mWEVdtdmL8anFYolURFQy
FdgJQfGi4eG0qbG4tO36Avk3cxx7CtzltPVSh+a8W58C/ckLAs4b8/irgZ0CtnsA
lB9aMx8xmK3aDnyZWxmgzLETYrvkIFNf6InESjwnRI6TBrak8ppkQl7XVyJ2uJpP
Vpv6P+RGBfUCo1Xy3Tj7FoIYZRv5+WO8ei7ur5TsbuDbKO4j/rB0ZJq7tHoySH3/
1Q9XKwu0mixKlazmztlhlt3C3+rSe/zkrZNMyLXwlqYoI9tzDPjsBSMpo1Y9+n/D
/fVGeInbdqylv9ajwaLkmrGSKzhj7Q4fqB3BuBxcw+a9PqCzywne4JTPCdb1OwIF
5ChMwlPpbUJmMFosNq02SRyeQE2KM/DFzkOpAPcd8c3DFWe4oJZ2YlyuuCMpB+Cy
K4JlSahVYJbInZBqClT6IhKiaWrcGPScirM1G/JcoW9HO+odtH3gLFH1+iIO7o9C
Af7NJ/DfdvdZkMKKysQ6I4pich+no64I0UWv06uXzn2Wzw7lwMaB/duvk2EsklNX
MUa7eMEfDjYCcbuIbjsrXajc/N3vKTsFSqJ6azCBBOmO3mhP7xTavzZL0eEvt+Bt
fmecXG+sJtWr3vhIauAZ1yRN74MB6WchEPU1w9aT/Dy4aSo9cWcyfpRp3JsfLQZE
p4C2AGuZFDdOnNUVgKiAtSwMEQOLuG6arVxcs6q7JD1ucLxk0V5eX1WGU0ROhZTr
p1Wh1deD0t1pQ+I7MPJ8NlFHkZtuSFIx2nNKwBsPOnJSVrDNci3f2dZMp6ECq43i
7vtlTm+eJfxpzteIbVUFE3ETfW3aYZBTIA4rS9P+GtQ7lWz2BXAEm6fCooG1Hrj5
uRPzmL9+a0fM9DFk9GrRD2ysTKzBzqxDX9e6X2fKGYtQ/v0HodGFvaPzHRcGejhH
95bhZxt0q6hk5NFYCYFMhKomRdEu6W+6pRxLYgqVTyIDZ1rUKdSHOwfpqkGyw2/n
fk7tvZ2/9H4NmmvFHbt2+hDXa7k9rPOYV5WxtoABRagpKflxQu8PXXnfv1bklVEI
4R+l1HTI1wGavk9afqIi2qV6NRsFomyXDkdMwYNbOnt6OHSdHKrImWM19++oD+Fj
nBdDjOWwlrT8sVpJ61ay0+JdvcfcOLg4QASY5jdBimHYBCp24liBo9LA/4FLcJvz
q5IU2a3atkkGb1waqhjSgsoLAepaqy15KNVD3ktfVPE5Fpq72ksUO7X0qCsN3IiI
4D/AWVD6Hn59PWdBkwY2sCNZPwG/b3ROpR+INZ6eUwbOPY1Yasq+//cSS58FcAFE
OtW+vsepJ+MWbSZ0cdLKmygIvJ7jTimKgmA2bXxD9SbsugLGB99S6c6R/40hLKx2
hUYyiq302TvhCCGACl+2/pgzP1EcZzsUxNhwon7Zw1tw8QGr4OA+0K0fjFSNM9BI
6EXGU3UIXspgc1dPYVjwxXInMYQeTs4VLQZQpZWnoa4g+kme2c6eykn9SgIf5wjW
m121fqMkoTTGXHV4VV78MK6FUWuBEi9LzlALy4qDapS4ulj4ZjOjO+qNBI+zDpmk
Q2A0AeMogp1PaFE4B1E2oeILlWWnd4bBn99fDbzMNiY/7QTpE5rJ3huvzlWjRqjs
ebJ/34pysElyTkiyrcyD4syRXFUrdlhnFc/JAcIHt5GSpBYfhTdTDg8ZSAJF3+tz
9mkaEM3sauPYA6R/yD9AYlSpdO1RuLNoSxxfM/eXCK+kIEZ6yTfkLfYKrkTgMcpI
ZrbTZCzbvvusdt0bvxqZ2rT3Cs3N0RHbq7r42QrlqzPx4QyL1fHz1cWR/8WWXEb8
zCzk8E1g2o85Df761haznMWfbbrAbKVQ7SAZpLD0bRppg8j+3ec0kyX01Pj9B/Mn
SXg/twK8E/XTHoQg/EzQcSlPgttVETt8a5gK7bu8FaCAsfr2Y5r4OCOnDxBN2tkT
dgQh/s8ZDDdLhlD5nZNL91LLwdl2SclImwY7gDM012IO/X4E42xJbFnRYgDYdSe/
tkaGDKXSGbHnKZlM/hRE6s0Z9w9bxjY9bZBfmLPPke6aY+0oaa6pUZ1qt4Lp2Hwh
yozHTCcJt2KGA8gXqR08axCM8sm4u/PXKqy7r2WsAZzA5OYVY2Dggzl9hGD2CctV
G1rK1TGT5XNKpd8Bz+1Se4keuQNF28bg466Gyyokhc58zrzjOwWLctWjpaGx8KR5
naUrdi/otqeWn76UIYiMImCnII4Mq1oUj+VMVqbqI1ZBi/aX7/Y03dZahvtlGzX0
Jgc2OJcidmNj1qqqKurRuyZJOa38S9SqRgoUi21p1Hh1weO+QaxVvLJC6PUeMkDD
hu6doiqsKsM50jkjtFvTMdYBFdmpcEAup2vW8wAdmzkbRJQE7GGEzS1rVJlObsLx
VLiK2KD9NyYWXfFLW5WecIkwatAlDlLT6QktfmF7RwQDmJqMf3Pw+SReaJz+ODO9
kntNv9t4fkMHRlgGZMtL01jYe55S3xGJDBuh32kz8pQ8vHwP3/JWwun79mfbg1iR
l+RwEK8yVcchZXgKNAhWZQkAgj+99TJHasI8VLFnd7gTWGlNt2Xyi+UH182e6GT8
YH00tomJylQzhv1VLyXsrNHysPn0Yxl5Gf6e6v9bmugpQBanL+eVB/ubgk63UHUb
1SyhgiRHtmCVs/j66XzZpFfXW7JFJlawD/Bnv5RlQVcSP2gD4iUWE43dsNAY+syH
9a3/dLeGXWZAsFhbJBx5mwE4aqpWZ4yeWWiNxo4zAGWSdt3QA/ub4Zs1GPsQME2A
W/0ocsaa3/aarfnG06Niu0RdmzzyqutMs8oU+WkAiObTIqOSHV3K2xZihL+jdLvq
hcIlpZq1ACxbw07j9zC0+5Up0mesTOyVSkJh5/3sqMV42Y5V9NrpXGi5HPwISmbr
2TBXXDKT4RHngIwr6W0nbkXS3ufM558gosB01iVE+B5ZRUSmHsi3SFEYM+x+bFGE
RkwaDsZOk50pN+OHylvxx8vryfG0IFctJxJF/zFJTyp66r+4uf9MtCfzaDsRisAT
JSDraipKea1IFhWrMSXdyraQa9kvKQ9X2ZhKF5ZmFIbkKgnCblmCrSNw60Id8pCs
emK03x2OwDg4PnBME5BFVV7qrzjSm6dQvCUjupIZStvEFgqvS9B/dciFSvh9W+qQ
Q5JiiM5pCa6ZAJYPGjzu/2Ba+LZC9glthmZIFtfhk4+vk2daiEf8i4yHgRuuX/TQ
wHCiLlWs9FA7O+BLeSM8pBo/qaFSf4rzLFQEfFLY/blo2VarsBAR9GIFfWZcTuZf
UlYqe7dunuMRJEqjq4CYZNqQmRKpY2KqgKw9O3lasJgeURcnIZFRrMrXhAY9i7WT
ZWBW8MUz3cZMzoTmLJaqBY+Ka1J1vbOy/wrb9Ylb1OThNWvStPDOs4MOieDFOkpZ
dMmmXo4XvAn0C0SwOJnnioa/FBkUcs/Wq0zzhHn/cW7BhekQ5xdDYsMQXsTMo+4Z
HSFwICprPsVe/aCo6+EXWGOST0Dvk7DQlxIpRETGCyfGcJIg5mO2D5Co1/gRwC8X
kFXawlWJySIgecn6XrP885Ll8z+tFNWHZ/29qmx4BiqM/tYaFjOPUNxPX9To2uLv
o82aPlaL8tIVidgVp3BuowHflCW+9AzoF8jWtnQ3clLjYysFhu6nZhs4G3+jn3UW
/+xwqJWSIzDJrOWt5HXetu2vk/JI+b8ogzcolyG2aZBKJ7/fufXh0n4095ZehNXg
pZwSd5fTIRC3DCYS3ZAPtHdw+P7dXZKuY4oPTPATBq8RfrzHWZpajn+e9NDyJt9T
vLtPctv9L8sifNCr9uZ4sHtCz9IXm+i+XvBkvHWcdLDO5yJB9I+TTmZ4rJECLx03
r2DDR3gtkd/Yl5xELlX72xlNQgjwlP6FhPBYqNVJKsZCYzkv/NHivQHveKuo5yfx
02dQpElNsz8WhLn6d8xLQEzryTtMV/z/xog9BfbzrO5QrOtKF7paqByDfufFHa5P
rG910RDdymuXEVwPjZGgOzEiVedscD1CQw6jtpXumtvwS1PbVgIuWYNT8oaqtO0+
h6KU4PK9yEocYPbIkaEOEfI0/0j6EWcEQQOr9ANx1U9+Hb0cVFIuw7Ptw8n5BglL
q6rC9Ec9wAJKHTfu9VgzcPw+FpIm6AsGWbWIyJFJUbGei6PVE3cI3NzZMq1+0qqg
mEqJIVf3iDOxOCVp33yKqYWPhLbhKGY3x/VvPEx0wwtv2sJqUMHvNgNzukXtxxRX
+h/Rfo+JgpozLqAKMoo4PSQxPDZfun3Awlj2AyS6GzdrwrHMwtjo1TXBk+BkGpIR
pamrfWaA0lTvdh+KZawdiWRJU9gJvQ/hMl0GfRqbRdre9g5QsxLeJVhVZ8DZ/aP2
N/Ovedq6mKurZWSsbXRKWgATUCro8jAmefYoOEaj4pwhm5XgCM4qcVWqNu3ejKDF
c+xpLokMMdHlOYAwaRvPxOIn8IsRdVAy7cI7vs4cmS1yBmyXBpIPvwJlLbsKzVJk
OkyDmAsL667C0KLBr/yKEdC1iGAkSSyh5LLcuzTkcPB3RB/SQMd3fqIaVLTLz7Wl
sVb4aGEJF1Mfukghwp6JwyPcf68KK9j6wbRwWapOOrUXGWDzgz9mZ0kYTcYYhK5A
o4HQr2tB1DRQRxBXjtjEzsLZkkVrjnDhXZG6u5N3AjGFrmhXj5x1Msn7WlmXgGEy
c+kCe/xLYUzT+3rVePPxUlbSdhlxK76VmLhgRcjUZOHSjogS++dMxEQmjjTM1HuD
32GxLapbCwIUZ8YJ4/z0baqinhjJUy40+tsM+/uW0DQm+GCe6gUcnpIFDbNgRcdb
FNcL/xRHtSH6DG/CQL824GtOLNrQK5NdjZs3+MJ9zVJVSiSfiGgqdDAdRU0c2teV
FRbqcGzbY8Jt4Ot/P6fHojdButmtpzK1rkm7jkuPF6Xn7rcHwVzZFYAWJa6edCej
hR+M7QjlCoeIek0chj6Omm56aUeYkv3c+WNLToAS2y8bOaXCU46FjVzIhh/mxtcB
WKgXwGnnFMhm2YcNf3THgJSiXr7GqYhkK1x0oix6C87VWhyXcWKVNHB9icUiNIcV
RYQdsrC+m1in5oMF3FI300pZMxT+ETW23e0DgutBeAieXuZeYMgfAnAKxnEbVmON
e+BDOxiXOhyfmAJkgSIVLePouCr560fw+LWzPagSP6CPxwxoY34gySrltR+p6lFl
A/nt36Zxfzs4fx9VukI3SGoMiL5SW2QfT0LGqn+MnuB+Rylel3Mk06IP+NWwCPSG
13ZIPQs6prquQTCgcAZeciNGkpkOS010fQ8TIKwynTpckk3utzjIRRSk0GqLhRzo
vO7yf5Xc+ZBDc9Pe5gaCpgtIuCnXVPPfIdwHkEccO7wOt+Qpxb9wmVVk/5OUKGlE
f6cYuq4iipT1utWFKtERcwUILyAKcKzFlhhwKqRDIxBpXYkcsv4nS8Ok99jDofH0
BhI7FTpoEyIyhmlRah+IuSBCA+suF2bRMXtKYFEH5KT/oBn4zyXAL07Yt/iC0hxT
pBLpiYOQLEvgn22xVnc+lgc4nHZdVOxcAei2buaQEeF92O8igpt0x5miG9ynP28k
Yf2h9NyAVKcctNiVV/lvCzkuN8yTFRgqr5cCMJ00P3TWEjjUxOVyskii4f7LJCIg
tfJJylBGNh6RV+9txwnemmbzd/crcGoj4u6cPjfcuPO57UFmd1/XV9C8xCDOsIse
xPrjreM7ADrvJw2QYgIk8Dy3gVc8ZQ7GKGGTd8NQcDgdLRKZ56GgUbc78wIzRGFm
EbMoQXkeTQ+/CeBKVGhNS8hCtdDYySF/2Dk83xwQfjNu7jOugwmk6mYBHfkN1nDp
R0eqICEqCyh/bBNW4Gv6h83g8tjZqKSZicDFvB3qRMUc2NrrOiAV4i0Mu3wMQHym
ZPSQLuQ//DRa3dP7euH1ZVVXWZaPEPM+c+ozsrJU5bhmvPo2PvmcZcODgS/9JKDp
NiA3UhKAi4CMNdwuGrT+nmz0ZXZO6mRRs9mNAS/LbqRYdsUXM79SY8ucmJ+TcREh
dQkmoYFFLg3h3qYHkOhqIGbpDADW5XPtyDAsNSnFvRPDzGNYJxOSfeQrtf/V4buf
zcSJY5sPGmjawXjtyNWHzf2Ik6/Vw5V08K11KBThh6R7pnw3Xa/gTRVx6u1zI0JK
L7aCMM+AFzPMwP/84n6fsFofmrr/rHWAv5RntXv+jwPlJD3K3r7HBY3pWtQNtQjM
zfdTfbysrh+H4hbor26GGlU4WAsFf2vjtpKJ7tyM7aKLe09rXGe0OYnKXF4ZBoiq
RJzWXGoplcKUn7Z/hlyXncOZ2LwR2FPu9eFPgbVf2ZoMspy3i5aBQXTyPy5xYJRh
F3t9cqPyGc50TzWfdzzZropxyEy5KnBCgE6r6/B86KhgiGMkUOZie8k6wSHBFUJ2
3vz/iXWObZ4QeVx3nER24Hz/RJJ27YRRU4T/p5MNq9AHKesgfWOTBRSRsGxl65DJ
GnVAKlbsaGoUaU3oT98pNLqc3FKI4eb+UE3M9LoQ0qziMo8+SWtgeaCGvevip4wA
MKdzmpPldO/zvSLIak5rotnA6UizJ2d3Nqz3o+oYHct2zF8LwUku+t+hIFR5XyA7
0GSabcRg/TNewNTelFWLDyLfhYucwRLcgngjjj3VmeI94peaQB8xW+cxpGUh6+QZ
uNBc0o0O/ZHXsoxiY5XyscPONz6ey0OuacX7QBJPG7f66HLuh5PrKGLoOyBb8oLj
Cb9qoYufRNXAl8vbpuILF6et5IvaDN+w6/UGvvPnUU8d7WEeRXIVZq7lSvF06Cx4
dOl4kdL+m+we2uu23g+OM58WxbFaFPTVf7qjA9n2025p7qa6LmDU8j539s0+NJ1I
rT5C0CNmAEwcz5eG/qgas3VtcKQ0/z0yhxojU3SIRCGJdOQnlZ1AwmVJvIgnhnih
A6QFgy/xJVPpMNfdqt3NdG7yAHakWYnFTU41PSmRZJw/XwFqsgiKR1ljyhbDjRbR
FgBZ5tw4rOyijbhQHgUIR/Dhw+8No21BcKi82QgsJ8ek0CzDYg8stBgeMDjo2Q9H
Uyu5xwiiqZfQSVBruagyZMe+XRjiTLCbS/kWELTcKF70Ge72hxUOJ6eLRca5/B7x
/6CPPc06DE9PdUnvoYecoq3XRnfjOiv2Dul9Ldcnbp3CC62WE6ASDPVa62qUyGsP
QWMFy3W7ypttGd/UcJMPEGEAsA+M4sCmfANnRXd/hnblLZtqnCorwxpX9UupfdLs
N+hj7sjaOyQ4EuUReA47pN1QaCsUbjAyaUMXXoZslgxd3XuK/kx/Cd/PmMo1ZpaW
mMOhYQQ9Ssd7GiLDFQvnvd1ZsQAtssMolOBoSg6dPvxXJDjPVhxWgTuja63J/9Z/
pPI8ObWWJEJRfPDEoMiXb3DRgYee2vtbQ8JsTHNGQf2ZofizK1RFf4HUzCFHGIAf
oOKHQELYUXTkW9916AxUSe3jhu2injAj4SG9koCzSwsaf26Ff9ThyjhmtJk+VFz1
o8tOUYFEmwkRqF//WB4CBEE3a5DG0DYInZdf7329q60/YlURLTlcsjajJvOq+8xB
D5xiKzI/WU1Bnv8Fx0r4dQ4gpxqnIOryU+K+FLdn+MvyN/FTMfGJ6J9uIu/U6bfT
8w+8Mhl6Ju5u7649T0ct7tJAo9sY8LWQ35p2NjGrkpSGyREfgN5BY54Ofy7yxcUX
3WljBk/LvSKX4arLpFAM5KMnM1xPzIK+zwkmjBLU4Tb7J5Ey68WqRfjx6SLmfZAK
BlO93P8rfBFrnTAnR7vKYCspL/2Zt0tKW4eYipXAx+lC1qxIlgYmAJYH3W/maReh
FzrDcdq/DEZVRYkNXt7vEtKTDnQ9h0YI5sUesk3CTtPD0jlScQz8Vq2ivPVmcXQj
m4pbnwJgtnjjnpIoKyeJDzWrcjfBpjkNLqFMmUzeGXRxDvkm2SIbU3XtWhT2PtG0
tZ8zxPk4gyikOpSfjzOM3dU0LyOPTzwJE4WpBrqiMaXt0PxdZ1KhvWBMrdCuMveY
JArn5uHxwUExikHs3J4+ceP31AYscHSEeaPuf9JtO4bNW4ZLqxPr4VBgWTl/xXlJ
ztX1LAs4CNSb5SJ9EvVArrkxO/fmJVfhW24PNh1hXBGDHQae/uqqO2xIMOJbuXPw
hfxeCQ+bzZkVLZUTcvvk9KeZLAYkAF4dx9b/jMqVO2n/aBz2q5PzrCpbtZKBTVuv
A/qjyxfbRgDclcUoa9ukCSPRkgujSqv4VDzYlYkYoKJiEHF0nEaSnE6difAL1DSd
Ye6caEJsdJm1VUPr4pkfVIrNIapHv8BP5LDOw+JNjtKU2jIVhBhkBU7L2zgrQdMC
GEMYzUwHLXZA3JikUEydurCR2Lv8A1WlO5kN38kGctAtmJhiRFaOEBkHm9XuWcQt
A8dLk2kDfHK2VZ0RwI/W0LNyvz2K3q3+/DNK++Hjp4ARzq3IM/0YIrLNgnM459kG
Z2tuxY4UdNHqZcLnEWZjbIlsivaskxEvh500HiCYfCqfMD/toE0kA/D4ihWwjR1V
3uzdfMaUYGmEnIa+JV6LlwbPHrgKv4c29JlVMeyw7KRPDz+uEcZpVFoxRQrtmj5C
LzbSGIGhxP6nEBLTajeYikgCgOLzZ49Y8LO5lc3LRAm3CAQEp6lDTu7h73JlgpGS
cK4EMX0F6SqwClr2xqZaIAXtPWmtg4qYibAHiLYjiHu3FO3v+HfXTyghSYtIpzRF
gvB7LPG8Y9NOxZT4GxrOjHT/waFidQcQdGhkIvxtWg3/VLPHeKMyg9Kxc+nRxsw7
IktuuWLjypG95pwfJt2Ci59wLCquiW1G/0zyEKum2LlrubovLb5UQSZt5z0aILhq
pF5JAz7ZXBYnFoCfe8PQG4l5GJDY35jlrz3Ikc8RYz3W+ZSV5CTMQ1OfTEYjVC1H
fa17H6IcaC/v1vXznt6NDNefGIQ6GsUamD0AZmZ2Krkdn7FhxRZKm/0NQcErLqxd
fWmYsBZwrE5QgOBd3r6s1EM48IZis6tutYsNj7np7qyyziKKIA0gILi3zMehLA9K
hfVcFOS9IeojyLs3n1O7TYLU7RctaAkwk9OJTJuWWAjMd4Cg0He9nxoQc+1na14K
eggNZfVVapR8dGrVdOCh10sbGZcaWrhGMzDKOBWeLsG9Ypb0axsnY2EzOtR7CBEB
sSTmy48YdgQcJ7Q3KMD+vpUtuWBFVKwjF+2U64DHW6xy3P2ACmsmBmQgAhvXXrAy
VkPd2LeM161a7laZt5RaOyG6d9OiGQQuNDtLd/VR9jyQJxO0bCelmQvJMXchSNYG
hJ/jbPn+IcDK1pydlBVxftsIZ4KfK+E9j0JR7s449x2Yoq1MtdmMlUUkRkJUF20J
48VTFbzLxgwYYXj9OeBTQtxit3c+k0p+EOuzjHDPzU0qNZWZHmj53MnFof7Wfm7P
lN/hpV6UnL+mBZGJvBkTV5WjRx4IUo8mTHfpDBXSaSu6OPqzHCFlltDsSxGBnKxJ
BCJhv0bdnAf7jSXlcurZrNEUUeGS+1X9d7J9Rus0a4f9Ou66l/BmHx1pVpzjFFk7
J1RFgwLeI4aYY4ruPjbujBl6MfxV3+GuIurVXRvQSvAsdhBXZvLiaZAmdByeHMKl
ALuxaq7jOF3OsE6AUrIKa3/k44r84gA0Gp3Ucv1TobI/tcV8uXcQfMSuIYWXXwqT
cgKl+APS/jCMeIxJ9m9Tom0lJzVCl0k8/UDxTDqmE9k3X4KiNA1Tublyv5Yu7k9m
cIB3fW2mtQESFnE3EvVe8QaYAk22GyizSJ9jd9knSQRkYmjdso8zpDnS1Ym85Sw0
nGHkuTAU4ppjorwzD6II1Rc3MHC1lBBJqGWN0f4oy5zbdGHKg021qR64m6g1rmWc
VVO07GUWiAoOHRtVUiECxygvwNNudQlYruqVmpJ9xxICKziT6XEzFsZUIs+q97Oo
Zifkzx7aM2T3DwHjP5rfsgSpYR/mNVi3fy7mnWJYD9vTCtrKVONur6w/oEMAd6Bu
1H8yBt5dS1ibTIru1uVLrazX/ZDwKEYs1kj1F4UeoK51kD1Zve1t3N8C17yimIBb
iFOdDkzAh1yGCDFHNvKd0maAzazlbN0g1BSSK1w1G56CjoZ7if/eE4OByFGSSmdu
W8DuYfcx7BfvOJzD+v/Z1XD3TkabjkNrl8pxcmwDs7LANA+kJa0YDTN4ICvewhVy
OfJqb/SmGGgduHEs0CnHlKtAE/2pR7I4A3HVd+rRm2YlqEvkf2MkxYRW36mhNDto
ViPH8xHqEWWhW1YtTzvG8SafjolRRwQavN7N3kGOwsFORvIXyxnxI058od/ODp3Q
ZT9hRV5rS8KZstQPaouL8Cp068lLHTxeTbvngL6VEC1gS3bUAJkQVXMxcIN9fmHY
TUebguNezKx6R/S2B4DQQn4pvddFd3wOZSw+8xOSaFxgnehwku2bAbEFAFdMiG2B
EXuLEkCdicRbNoXRzPGaqArKet4H9bTlsOx9YvK+ittaN/DNU5uPUuuVp70w7nom
SfRKSgyvv+yTsELaqsPuayp2MdhMpxCB98Y/TVQqcoG+2elHtE8/i174ieE5NkJ8
ZCaKEIsrN6mLgANRvt3lzTU9N84OklGGNKraVw7ZyZsO5Ck9YULn2/vnvu28geyS
/Bw6Nga+JNxBDI/0d+lulD4XvSG0cO2Mm57CuJwBPncef9FoBInxpjLP9cGwTUXw
G2HO33vEgzRiY1ooMeptifpuCU88EUssc5HgTo2IC4b2tN5lZnSfcDZ33WJcnvJx
rW1LWi3pkZMqOf7RhXjaMQbmpscwPr8UQGNZkgtQpsRNiuYiGyBe5ntpTDRe+GZ3
/sWCc2R1BEyGFZso5PNKsp3nHDbWBQq1YHZWdrdi2Tq7hLNEjFw0gsA65zkHSk7d
Rl2DD7bvS1Wp1nWsWTIwaxLGqHF1DGu3fwMGYCT05msP+5Ii6tmzi4aeofa98IHb
fGdLXYLkZnlucdJd55isPQV52R+KjyGr2dv+/cWKBMF4geyrIu81YfsPZ8gJNbH+
x3F7hJrpCfnu83sM4kp0D+84Wyw6QNlYKHEw2SictxWhn/HKQs1dhOv/vUE4EOPy
zwYxdgE9CmGHJHObmrJcvQmu2mTmcIaos+FTQJ3dj3VUy4D1qgF6Tt4BingkNXnr
gHPom/BTXnj/yW2vN4JU0Z1H3U6L0DeYnNAd094g+/6QB9tMvx2O0CwajUZKhmtz
wYseFR8psx/7DMiB+CICLvg/wjHTZZsUHAtGAXYLvdV6b7NvfwGW8lT4t1637o4K
7RgFbzvgUbgbCosCifGWkavrhuTt7esGxltTJSL4by5gvZkUOz6MBHTQkp2+lJzj
iANTbcBYDEQ/sQNzMu7kOoKeea4EtLsq8Fp6blyhCMOI+ifrE18jL7ae09TjBEtC
NJsSkmb3nhR9hUSPH25CsUYPhBiUawkyKUWxOXq1DYH4FdKwlB3C6IjbIetjZv5u
eZHu2WiwdnNi2WJeNDgkJeLLsINuBe1Ka1ZOSuH0hNqH7Ky/QeITxFm/w9/q1dy/
xoX9eRfYnGNcL7ELjxe2Z9ie01t5NcIl14t64qGBxxA/ZV4S+MWlz2YRBBf2OEo+
sHnHB5IHcCMsS40OgV8eGDcltzJlH9X9yzFORwfr7Hyyp+DTZMD0kAxGd3+Zjf2Q
eKlRb82gwoKmixCOGtI4ZRdCXURz2Lyx1L4F5wIdG1ilGC6hx97oyocR/1N4LYY5
Y75TskTHaWGUDjxYnKZwBlMZ+Qx7BFY8Ig+b245uR3IPGtUEpyQybRlOkjSRy4yV
zMvCQ1H3XeMim454ubDfJEI4bXCu4zfoMcIYm5nZ2qN3fpDybci/MmbpvjrTokP9
ISeBFaKzJcAKwQh/Mkn2nTtxzK6MIfNynJzPFY57uOCnjEXl0MZsbijW29GhPVmn
1i9jC9O7qmYhYMo/1xQczeUQXGALRrklW2gVDz16/xef2JAA8We6vGmlzpRLN8lf
Wc+4svk63NDLzf3UDBuCmZL9fTAKDGUWPrEXJ1IcQmJdIlJGo3YWQ7efUvi4tBr8
mrndHO4BApeXLsmFlBQWXujbLDz+lY4iqzs/pYCcxLTiO7olLr7Wo91M3+40Nnmk
U0A+mEt2WHcdCm+jOxwk0cBKi3k2XL7ovxx9O8sPVXNGqSCbWpy50QHVvXz5s/4F
NyQ10OU6kTIu3Mroxjp5Yc7UuNNKVWqxHnokR+9NvLZ+4tTKwZGNwxOWHQIssTW0
31HEwimdpcw6iZdAoRAaT1GA2z9kk/qhuFNh0Uo378bPTxqOplC7aJUOVoLu+URm
vSt7l0jlZ4iduDdw1sgYKWP/NRBdC5r+KjKcKOCGpzAnY8FTAOFYzSK59xcr2z2N
U3u2meaTpLZLCMvJCoI3L7uNhK8wxrR5dZBaHGbGC8hCgbVLhtGYu/mcJY8g6r/v
CHBzzHxchrkWhekFBAkfIzvB7J0kYHYoziGg2tD1tpNH5i9mTxcvbtiClB0iW6nv
2DQQMZz7wRjX0xO1XeO39/yXaFRGZ02+98ZlaiRZDwRdMGzxipWENF0Yn/2kPXJT
8BrUAFtiJctUSEDLAVr98+I9jCGTHf4RDILTK1P0jCot5Qxk9Evy4rU/241U1WrB
ufTrH2s1bRYjlT0qfLnT7vmVJg0ONs9Y2+UJsj3XdqUkOSaHb+XuNha6mAkJX70z
2/y0PUL3+ZI0dAv8cO76HrAQP49Bodnu9jDcSinMi2zl9EVIdsmALtDiY7yeJovt
dTt44CVHtza60pm6k0EQZFbq7E1fx53ShhV0qAvxakwJNR/3I6M+B6ETU/P2zxh/
TpTvnidDqtKqBzT2LUA31sLtcYWPtK9t6W3xtQA9b/UsOZ6AzFvVIPGcY4NVvboU
c59/UhhjfNQA0yO62TAkIvWsOK08RpOase2zwX5OzJl6fiqY92aHtuVMPFFkyplS
o0u5F33Io+L+y6sR4Bnx6v48SYBRBVMBcA7XUcj2j/+I3g5r3ms7sdcLNBmbUo2s
7EXRp7jpc1mlJcZMuZJfuj3+07+nGrqqDwDRCoP6VufVF5CHnwr+DmiMS4WPVMug
umyFrFlDKQs62tsx4yKatzEqEwX1HBpxhr8LYIYypf0xYl2xZsFIvaZ14e+RIqKS
wAODfEp9DKgdt+q2zV2mCwX7FoKeadWewBfUGBc3C6t8dK0NHj6oNLhGEgL0Ad+u
1mFnVzKT0msIQHM5ouX8VBhjFjIH3v8LzvPV6DQwhNuCKB4QRVhf4TcpfXt3xRyO
rIG3q3b7geFRnjgYmhhBGZKBwbdjAu/OoBZHymLDzUI0sQtnWm7nmHAHTgu92g0h
q2Hohjsq1doIU4MdtCFlKsk0uUvhFeMuex6Y9czlIXinxb/KGKoJ2NyF3GP7S3mo
TZCFMpYhPcIMdQJ07M09kaKJidwlMPXQ8IshWDhlogfdcyWPhZdPsOH62T8FUNN3
dIlsOcZXibu1eSRGdPa4o1iSN5sLxk8k4FiGp03mlF17ro3H5w43JsGNbLMJS1aH
MNXIUEe5bX7snjZwSJ0ZcGpGB40/+02RC+gFjQNLsm4Rq99U6Mq8W7ukfgo71aS3
CfAOvwq6sIa8hqBg2FW4o9ozRnjQ+UihljNrR9IXdKhuM4KTeaajuVfgd6mYGXsc
gM7ZwtaVonZJKMncl9t+zxl0hK0jQ1oToUvkA5MsrxAaWhgtXX9cqJxEfvFZghAO
i+kGXtK8Gvd8BiRFtZbc39E/aFbS70JnwB7rVSRcApPMb9Yl18iprZQa0igBFLFL
KcaMBr7XcKJPyQ23JXGnHypQ/N39Dun6JKbQI9za0AqjCqLgMXFE1wmJVCphm7qW
EhQGY/6zlcUQxa6eQEiNNTDV3dENxcQD0X4miT5VtuYcl2Fd3YPpK1lhw7wyaS2v
tdxCLNC0zavdnb/oDLePtYo8x2DZUS8SDzKuXli5o8jzmHRN33esGlSP1cvNOmry
FXuIv3bNzmAqNvtFlxC/o3q9trXXa5mfcSAU2yoQehKNSY2vE3ISExQFTAatm2Ep
4OetKm/ZR2m1TanWkWDuBimN8pXv8tTmJ7Vww7OKCINzpDJ8RrPq7GtwPTmKmPr+
Ec1Q3xv13IMTxnU1kz2d/QNw1S/w5e1sa6jlg3CdJDumWJgklomPuUMdDh8M1NJy
jGIcmDHD/ZoL5SlQCCJSMRP+1dTkHPeUU3o0XyKhBVLEkE95NWkDsNni4xcyDsq0
rfUd0Civ1D2Y8e1ceeDhuPs19LIPk98vKkCmmzwMlrx08edChH67JE805Dqi1Qke
p5iXALfhlF4PB4BRfnfc0UvLM5h7iq5wYX43N7M9tTJ5BIW2FHIdFTq/etqNph69
PUWzRtiiqfakrONPX+Yp5CyaZCisdjvjRBqxVdesQOAIOsTCG4zJtT3UZOgmdwIt
1hSNzlw1XwuqoyzLJ2ERHFwIfZ6uLoNcdJ7uHBRsDk9brdNJZ6Pt+lTysfA3Fhpk
wB/AMJVga0kLG6W/szryiZHjprje1o/5dzs9HAQ3yG9hFWglXVxPiZ2klAbUajwG
th2fp0vE6rZaAKcHEOGK7nPwSA9UJdnIH/RuOpX9KTNi4SWnDechJvIANW52Wx8I
6d40qOFo6+po08vuczMezvivzaexUrLyComiQ5LZRvJaX7TCvv7PibUuh4cdGpeW
18iQi1y6mAbCFHaR0HOaHkMEa/3xutTJI4CncEKuEy0s7Ul6ambEyul/0FHAQUgk
TsL/DD0NFrdDjAqbTjdPWmpnkQUwrqWbqX1wzR7TKZJqU0TttbvaDaalSLh13DLS
63dngB/Jz+OYJ8hOzU0xBwKt0z5WI35KRVOD2Fc/gJt/1g5T0o1Hz/yq+ahugJFp
RLfrObi0023kLKa2ihkpokp+BuVsd7UftqpfdKls5b6n9n9U27pEDjm0Nc2kUcFE
fpzxFiA7IAd9cItZRnUlOlf5dBxLqzFX1yCfPGbMg47ihmwYsJpEW5IAqlBx8w9J
mFAvujOtHzy/E0iGJYev725WoIqVbu+g+BfQ8a1t/fG/xxh+pjyelLLxhybqX3nf
8KqfFyG9wFa+8N58AaBa5DmLeDzwt42NQzIyjLrnSV7L/KtWLgwuhHlAxbJqdThZ
UR6/tPBTTFbv0g61XK3Tu1Cdqua0g8FPBEsORjLVL+PMGkhZ8oYsbgdRAugEyW0a
TbIXB0tk6pkkR1peoN30KHpSW0LIwDbVQwZMVj8eWDN9/UMDcEECW9tOPJISsRsP
pKCGps7qz97qXd8SdIrf4DG0czRSSkHyb/oUcTDz4qpWu3cktiExsRHEUU33+b0n
Pmt2LSykCtqiO73OZ6f16oo5wRdP1vLvk5apnk0CerWmEpFiyGEVxsk+/KmEG1qB
CozqQCC7r9VnF4BGXq3lbmNKPRcRTdXHr0oREcO4kGsCiC49YFAXF9GiGs7j4g4m
YtppQerMnm748+qVYV/F+Eytlx5qfv3ObWHYmM5xYJTJuf3uPPL6+hJpu/H3P75m
8hrEMYPkvix7EuyzThXPkUhamEprS8eExHx6V2knazokrFHyUmZznFwyyXyc0lIe
1FCdPb6XmA0W0xnu7yEfg2LNsYJz4PJNrZdcfq47EZvUwOtxRe4Ulh//bJtSfSy4
vvCEQJvIryOUqcCL39SEoOtAUSQTSaO8gHV7cz/iS3PAve9+w2fbA4fFiZDvN05a
okt4PmvDDSDZPpR0Is5EfonG4pb6YaAUYTtKsRZmJncZm/+pKcNuSeq1Xbt410ws
cSN+30P0yPW9V9+GtR6d0LxXJiMN6Dfe0c6T9dhNjw8nguZCLJVkn4Lt9TPI/Bse
7hyOBxWJpFyA7nwGOG6Wws21svTNjppwwBRQ5Pff/KEkRhOtbuAgmqXmZIdIIxas
GXvmWWKSZGa/SLJgehiv6YKaEJjI1LpfClpxiASRnPin+TZSPThavA3BczY14Xp9
7dcj1YJ7Fd41Zvin5jB8hAN/lrREkKHL66bpEyYlOCz2dqL6bpJkxxcQNdezqNAa
j7gTloUQ58JHUbtZLvll9si54FIsO1zR8Sd8bp7AXQWBY/3Lw99R8axvUVm9JEFT
siNtIj0/73d4pgup/sqauPo+Elga1j/rVCgBeEp8MUz8ZhlTiUvsqHZZK0DrZjkH
L6voFGf7is6V9DleEG+Mo/EZqR1ocsqBY8E5dFeLLGG/dRbXy/L6Mp8kSEWFgSSI
44pVrFAHzNS9gFKOrQAaIO+3851Oyb0Crt7NsVAQ43uViPEXtQMt31EVyR5FggBi
H/SIDCmDX/B2jxYAsZL1ANF8/qMWzIS3XaDxyIJzcUPGS0aph+9N1dQubi5ee82g
7JfpCHkTuP3c0SI7BbKaF8SlqwHoNhZj69oU46wlKprMbV1i1YfGZ02VBQTKmc3A
uatsUi55e9/OJpcEyakUBCAXPhwuqWryYvdRDTLfyItbdYW1oO9VtXpT2FZszoEd
nLyMKhx+ueaUHGUOuE6I3/rp0BXLS+Y6/YOC4H+3kZGEXt+FjmRrH2yYqWaG3vww
ZuEoVdZQ3zhW2ghKfmBQartXCE5xxnpzuKClvdGAgQoZ8Aw2rLANEqv0Vlc9OgCf
g1DIpd56gV5Zwcsfpjn/KF63uOuDexEXiMyJr0DKJgHp3YRONZd2m/8Y/QHJknXQ
n54oz+dO8xiuywarAW74pgbkHq6XF8r7WpZiQsCUwgzMJYub+8eJCK+h/wLf2je5
4pFithZ57jyIY7uZCfG4T0fZS/YovHGtVl2JpzLTnOI1/BhJyDjAJuTV/mpO8adg
LAOyta8P9iVib9HMtUtVvhGZR6s5j89sX+R/Myfhhda6mJw3xD2oyui62e8xIhM7
4gSfYuArDweUarsfAkkOKp/ps0EARjak8vKV5RnicsaeeezyGq4FDxi4UV8RgMPz
t4CPpMierN2BJdpXfbzpTX71V1SBuRpXyL0dPBAgWH2g6n/nHkPz+NnE+JFi6Kjt
BvTLZyKf9CV7xrDJtsLCbsTfwbFjsDXpn3AGJZiobIg9NAenPuEAmtjbd2aM3yqg
mUhDWGhK1DvRzoa+70v6LB3DyXrQmvZfkTy0/k9CNG+6xv3qjPkQTC3mMhmasfcZ
9dnfYfb7Giv5sofC8DZFPykY8WQ+wj691Ei92d9t/hxm++7AE8IALsc9QvI2Tx83
6beBL2td/qPpakO9YoecS8RHcQH3sovZg30bcJAsNRCgwEpnDqtJozU3S7Hyzrq8
I5oftxbJJGMglQAYGVdjtbxG1MfU4y2vFx8PjWKXnNSok4E18SyxxfqUTBijMhXR
bp7RlVofdKtlRBbnpmTcGNjLfQPurgjYujtRJQXtPOhimTd882kwNKjY6YaJLwm3
VzB2qG9a3j3NeB/KsHCVy6lgEw0As6Y5itCFv1kTL1SorgqRlmXg8WtNxekOQ+Gm
MUtRWfQ3Rd80QzH+j8u1Ali20tsIWehhk0RrjwYA4zjjTR7wUokuAoNK71Mn5+s8
98rHNREN9vG3MnJl8BbvvklLFmYNyy1fOvMtdzb44FUkDU+azGeH90uf45hrXmu7
wkZGXFq96AkDxNG3YgO+01MWB1Kwk7mahnIeTy3kOP/HgDqHIdUQ2gCdCMr1Ij8M
xy2nAWcgXLVg/lZS6yF2kpBtE+U3zBTs+kv1ROO/ifVLmZEHuJgEEanPVcj2KzDG
sxXdOMumlmTcQPBxaoaYGYniEfvQi5lVQutw2v2bF08qdLMXn8UZp7sMXm63VQKA
mV884qSz1GP0tpaqsWFFQWwVYMsBtZTGV4TFlmEFleHN59ZWrV5xY783UqVSVbA5
chjZURgQuuvFnzorl0CiN5Z6xsPX0kdeWy54vFWTl4xF8qI8CMiDKTbQjHrRK6G2
OocrYAsKk+mFCalV2AKuPdlkSBuQn70MtNYboSwN5EpZTaVkgjhCISmEMVtSCtVl
x1JMVuyHFRqQ4x3ZrzSd+iqODZGvxSwbQzZ/WIGsbDt5zzqsZ2J3e/TnhLSVEVU+
JeVYXP1rumZWUDBFUskypvvb3FyRB/R7wOA8o/h3eBY4U7BbF30/0FQBi+kxBw07
uafB1NDEuTblA67roGPEfNZALZZhCBEspUII1JooRaC9rChVyRoxXO6qTSDdptf0
J2cmJZh7sP6+k/wh9DWc2B6ilQAkmx6PPyswEMbc0nDkQSxE2LHrLtyxbYOct2yA
Bi1c2Jmb+N4paBry1/BPjBUTkSpndby6RNcSBKW2VXUWiZUWX3lbIA7QxmcN3EM6
1YyKALtWO5szdBZuaWeLvzFalivICAisuwyjNweUFaYGCARCwxqWMvQIq7BIZjEN
6nQPms8ueAdRUiJMjQG5p9RyTIpb4x0m764oN6Yld89M4cUEeaymgVJZq5i5dA5e
B83xIwZg2Fl9z0dLL6opGOhwMIjr8iRB2QXHCc/JhMdbHVksF5kqljBeJmJfs1HE
z60xMcBDsIb4L8p6bSX0HS8FTnJB0i2HQZ5uOJ8XTD+7mYiYCZ/x4sNpMpKcOnpg
nq6sbfb76HtHQm8sA0Lo29GtXT20KHWDa/iH8f3e4qXR8h0Zso1Q0Syhby4kK77p
EYr2g4yDEimvFzh/b0c4V8qrqJQyfMINHkudL3oLZ7/W1ApSfxklHb8Gi7x89rkS
H+yzsIGBXnDONmISLctUlL3TANA322lQ8G9Ec6MDGbMj6SjjFkOVdSmKFBGb4LCa
FD9EDY/zoHzkHTlwp9dnf7ynZzSvfWjsm+i84m+Pdtd2eL2HK4r+s4F9kuYShuPv
HDJAQjrCFSa7zuA8EhGk6qOS0SqP4KEhZrifz/hjOJ1npyaPTl4GJpUfWb1vrYVk
wqlRyEAVHPc6Y3nBEGYWFiTJrDsJ0AntgcVCs72HZfbw+qT3YxSdQxUIDEBxHldf
bhGE+wp/ZG95Girr+c0O/IOIafZ9bo+z2WFC9uBonqvXnsmFhN5xcsostn4BJcn3
QposRpVZTr9Mf8SvnbzWI1sYDebG9q0QlwhPQxUnNbEnIpGWuQwtTGO9i1QcjiTr
7W6Hx1by7y0GOnYuhz2V/pfGztQZfSj4TIxlhCU6iudZ8XuIaEK0hd6nhIYarobG
gh4w4WtQwTwY6Q8bNbWkdhi/pUo6l04y87ZKIk2R4fBSJPsphPnDiqLm7eLAhqLa
R3gZyZY156mmcz9E4a4/wApICBOxISijOBFLqp8iuTQdqIrKyWUSHY+NbTlv+9a6
7XPZe+5fK8+4nBdRPtUVoBoOA5lQITKSVE+OSqqlLjuGgb8I7+lrm8t3A28fLL8r
C+mx1fpjF9iuoUM1TonqE2bfFY3M+eYT2dB67M3JSOiPb6tmj/zt8y2y29WmqyTV
ygXfo5E78WMFzRbwnaqIgDwhnXwGfXJO+CRs3dvuIxzHgRq25mwZkfqYFq2T6sr6
m/Rj7uZqbVp5rBV5dwY+aJFpP41gV3i1Hso9XJd++cwYXlqipE+newIuWQ3kv2fh
L3tazbJgeIDVREndp91mProQvGsgoBzhKAxzuR8tr6ANrjxsCO+vZtxxCdMzoh9G
SGSliNcnYMlGJQiLvWOl0F94FMUhKtm/yt5+j5qcCYfvXjch9x6vZ432pgK5ig9h
OxamA6GrA9Y5sHIpEfifnwTRHhTsVeMCLo3F3v94C2Ob52TJT20Ji6gMDhlhjw37
0x2hekuiASPDjroQb7LGusBcXyS/n9YFwdfJll45qd7DSTImNs+rwJUH4aJBi0I2
+vZxYAUvOKsGW4fYeS4kkwWzfr4WGv6E2TG1HMF8bPbZTnbi1+/LEpZHYvNyEmsR
HTOLnZso95lIfqZNCVX/KU5K9eEd7W/uIiXkGhAKcChi1+XVidE+CNXIEGNDGhEN
+fm958cTPT2uSrPnbsz5k80oU5l6v9xfe8t1NdTt4kOCRHJEUw8bGFXXKlHqlchE
R70jh7umkCGFoyJ3h1hojes1aOPuPwe8LjwcVLJ+1oaiYuso2DGgsq2UdOv28Oj+
46G3lR65PDbPSF3x/d6VPyPgwfR80s4ViScT8z67rqT0sSsMlotwW47ls2pxG2q0
n4UIgbPcmmipMI/78UUyl4/8opMBnVC6vPAyu96OBdcsRHtaEANQqbmX2XAhy/xm
ctlwomZ21Nz1fdUVX7OJDF/Q8yj8heT6N7UfosvOSpamZsf+Cw4iHu2r+XGWRxzB
UPDo/3KowKy2iUbFd2gaB/zP3xHhqCa0KTWjPVbZJy8tbdp7/4WvgAROorwiiJ2I
jYHoKv6Bk0jnaTl5JKS6JicW0+9cOnFx+JNdW8y/LdZ8atEtQwkTinxkwL0pJDT4
+e63Q/wFFS1xVkEtoLwoMXlsS+o5I6Mt0MPsR57H3LsnM1DMlQpTJMevaXj3aJkV
IauBHLVGLp/OGmzcivI1aa2rM7EF0WVxfQZbDqjljcttj3a32bmdkDq1BW809ksd
DZ1TzwlMHFLzLCggH1sK2EkQuV7K70Z3vFCdnJQFrqEvlrzSrGeKcIHZPCAduolQ
eJZSmSibk17LcHdlIKSnYb6/o4yBSl+2Z9+07jGSC52VV3dWfzIH3cVIkz5lUDxS
WX183eiW48XuMu4k1VF2XPjwQg+BATdKk5CadZyqhZPatVM2feU8xPqmm67mp1h1
0KW5U2o6OVdGZl3Xr2ppWzed90Cmf/b27+IoBw97fqmuqneCMpMJnigLGWdT/9o9
LUetNGXRDZ14n2eHYc3tvCQOjqlOcFM8293niVDGr/5hYFSVrPYOgQisAOcHI+Ow
YptVtj/FHxx7MffoEiMRKsWW8Xw5e9UCjHsrGdxIbpFRDmoge0G+LsQIumTTxJeI
8U/zL0SThmQrRaOdT4F754QerDn3WctJyuPbt3fqGzPqYI6tF85IMkrCzqYCrbh5
IbC/s7AggXar7KYIlDYK2srC7imhLYH6Jb09wWKSnH2lSeaBMU4SiWGVS6/8zgke
759j/WIGoA4DOmYJ/9h3tupFsbl6e6Nkwx0sEfJ3G8S7/Zt1m8y4I5uPufXS5lSs
+nt/Hzhtdw7wNCfWNKXo6qwVydwtYqJ2ajqHV7EuN4TYYFSEuiZi2GLhaHJ6DYNQ
afa0BY48uf0UKt5Xm8Dbo3XXc3J3Jur83wfBC6Fs79u+TZ5jsnmI2xyGKXJuGRbU
egkTZtP2G8ZltL0m4cVs5bLUx8BkcDXITv9N1e3/nz9KRUG/1bLxKOmNVH96P8Kr
NBD3MfwE7IN8SDXGQwyL8qTK3fASEb2VvH8TeS4NykFY3EloiQSvwPynoDmA+UYm
8xlHD8FysTkXa9h57aTI5FmJiZ+Kd0WJyxbqesMbaJzHNUpjd62rSd30gF2sCE1v
0R+8N4CcQ5jhQMfDMeBRwXmN/C2qqBB+5AVyyqzXAY/0yv7rEh1/dAk+f8/CSRk6
mbq2GXaCEhKuwvBa2pueEGB4czd7e6lrXecyEC0PzIqP0dzLq4Zgx2YQO60BiObb
8JX/6cHkMrC1DTAqW+IYf9ncbe75hO6PwiiVHIUFwUYqVT2kFka5ykxbRkQXbM0j
DuX2tANYjTFA1G/WcsRt27hYUf836eW9Uvop6DYdvCvyBEgjh9j50qsjaVxdlmmR
cDt5pAiu7RmBM5BBBPhUdl3jkk8NfKVrxPh+Mb6WfXjihrjCV7yWmHlfMVKv92nw
q1yyrvl22/2aCC44zRGlRQUUNuaeu5J2Z24R1PtakcZhFob43FCwtyt1VUHo6N/i
AfuJqaHpKuZ7It/EXldOKCIexo4k1/Mpv0MOwETzKqIKOUzlq4cbyw4QNPvq0ZQh
2boDPOtfnGkcZPH4Wy49qhD0rhA7E+/3etFBVkfWQrFvKmoMj76p7CJS/b60jxkv
DMPpY7ohxCB8bVu4HyKtSjzL3VdH0/dhqS7qnJsige9jg5ZGUoKzztZJZC7Zt6A9
Y1v+GDQDSm8kKbsh8uGwo9uoFBtxGOqErAJC8PYPvsAFI2EtpeYKk4O1S7Tfq5Gp
O2dhmUH/TvoLGPHyx/TIFVwvn+h4ijgg/3fyB9tfJS5fnc7S8uXTPunN9h8jRzoY
9imUCe6gSiWK4zGt61bH/Em2SgZ+8llJMIHYOiOltjVzbZfKMrFoKf2SARob7+fg
KT8Q90WDaREpLmkf6WYy608sNVODLf3JCxw7dmHRFLW2e9fhJDcybkam5uNsh4IL
JGAeWk4/IPd/CT+LZ5clD5SXaKSxhUH+zso3V2XjRxaM0jyV5ZAX0tctz4kqJR9D
V2U41xBDvV9O6bMcTjdYzxz5DY9pSVMIgI8qzRl6MNR+fIkzsb8hH3EJs11Csvml
uxSB4oNnaDS8qQwpp6vgH6EuKV09lVY5OAwRM4z5QjpAArAmbLWSKWNds7fBZELy
L4sBqtnuNfPHM25XbjYfduwn44X3xdoAEVGkivqFaLr/NvxCML6CF+PFv9XPfOeI
vEcA0LRva5Uh9+YAXMPvMKy13b/XHlP21YhbqhShOaFFKB3CTBZnlsXQ9JxpXAR/
KN1P4iL0kceGYQarNjZSR9KZtf4L+ha32p01ff3J/cdAJ5JbX0g+Bpjt1xP0n5+d
2G1dXIXl8rSWSRLQjlKuvZutEM5EzOTQjx2lTlUDG4YoyfV8BFHheI2uKh+dvdZJ
0zdSOXSmQUyuDEnAvMzPI9E57vr37xgj9s8WTY9Rg9pNwjchsZ4KqtJ/BHTM+E2Q
ColowNxh25S5brzs4i88UvFm9HDb2b0W1ShOqAVf3tOpRXEfH15IPPgtqsp8V0nr
ahaGz9IMpSbmIYKDLJj9OrwWvw8TUffm2mIiYemgrE9FEeFA/yZ97AcZip1outUo
LLfOZ3IiKX6vpZzEXHmCig78r0Y+ASUGa0p7zH0/MejpLcLzU55PPrgGS+PsO4UU
W3BLpiz48Mg+15YSnU8zZqaqzGk2bpdX5rFDfEI81BxcS5w+nk1YB4WA7hXi22RX
7kqMMnHTVl83yEHpuvNbog6gDtxiplAygkZjuqYb8VH0kkv2NC/WQ74i/0G54NUp
u+ZFRwkrgnHX2TMHPhMyA5mpEl74UqBL5UtRwfIOuUGxpYMs379qk6RvKYo7R95p
WbYGcEyJyJ271MJSi8irYMh4FDen6W2Qo/EWhexW4HwXMw6lWiBPUfcFSdEgounE
jVf4pKBIFjV+4Mwl3i+BdqCaGXkcDqr4dC2HKwQti76IVREnw5hqmYjSkVmj43/H
O+MRss6bM2XDR/e33wKS8tvSEhM7V3CDzd20WF9XoP+l9o0nZ4NWjh3dvgXL+Fnn
yCvvhYOo8l487SyVpz1SU2gmv3DLKYjivmKe9RP/6Ops7NEYRPZGbMSh95ohdatO
ZGDMz2knpOEZa6IC75Oa9Y0qwZ+Izf9FhxVDYDsRxC/T7CmEpu+lUiizilbpJhea
FtZCYjOK+wudTSuM69JkhpKQQguY0fqWvRShtd9anSzkFPPhLzG9JPHtLJ1CyzX3
0aH1X2rzTrpM4dc4tQTH8anc1mbuVaVK0F40Q2ogvTPob70Y05wlMLM3tv6lJokK
ppDQAeiqLstUZNsS8VJ/JX/aDC26Mz0nit95TSaX+gUrjATSG5EfAMEA5NYgUdOV
1f8JzgJdNXKsTlzRvTRpQQnGiQXTjNYIH5pdGoRh2bY/TE/v8jQ/j6GSNekSBc1j
y8/Bs4MRLav+NnMvUjO04roTnCl8R5DdjPKPcUS7wqvOFdHDLQoT4gYeC2pOdJdL
GFY6ultsQEB21salFqCLFTu+e3XDDcICuOPJ5mLX0uhrjirJYBeWuNg4tNP7L19e
BDa1+2CmFFu1QScdeMvQAKmBdLErpKB/dl66OODwaUAydyo6f4SgdzIwvLBaNeP5
HY9Ac15bnWNzqytHRMmtDr7rAcoAL89yr1QTQSr2BVE99jktLGyp9945YOmpUNV5
/QOmzj9URBwZD8I1ZEUXOuAtvMsfVCx2oK7Cpcu1b5TDLFf/TjQRf39wIeT4ft/a
0qd32fjzre2gWNMli8UihJnf4fFjnXtsOTH0ArBluJ4RBDuDIctRWXdzuBOsbV5F
1jPVUum0VdKTHs7N0oqah7CKfXUfTauE7ucyCYdkznPgor4lM5ha2ZCbc0VObaJr
2ZkRg9toPInmvxhVENoA5W1Dbsd3qBcWnNCqcwRarJkcpAE4HsPis7Qxc2SYxZ9E
JNGyUpL2shV+DNApYi8mq+OqEMEIcEqBCQnrF+CxKzodrWyTckRglCElr8UFJKxy
kLBwaBSbBFAy+D9b54NbB+wNiCv8Cja/EVAY4INt7/LmSmHdgHxntr/hUOQ+yN8a
zJ+9KECJAwRToUSZEgH3GzMhPIiRMuA33MMQtq5KeSSDGCr52vnzQej17yL1q+Sq
rzzhaxyFMZ4kyk7dgBjCgmmtjA3DzhlIuqty58sQF1sJmemYaG3BV+alPCcC61ma
76K72W31fIHREtx84GAdpNYBiJdPG6fnlMNEtkIOFe1/dUVdq7ppkWV48vALyPxA
1f+lPnP/vRKYJkDJkY4alg4Z+BWzqDzVfRKR91TLlpk1VnFhPOoUNy7koYQlJUnQ
TMqEVqZcBAQuZr8Hvk3/O9jNnI5mF0PPb8pf0rgiHkZgkN5EqOEhqOUGuycUCDSP
QnhUY0eb4z7W3DYIGL1+UZ7qzgpmlqBvIu8x5k2TkO8gua/+7BHC1NddWyi9FRSE
FQFwOx+/x4jTAzxRYGlkBIHio/w4eu/nWgT6kW16FmIe2k92OWMqpy+G74Rz1kxN
IE65arLpNj/kGhGB00W4F2NWC/gXnxhfUi57wPOVnlq+hjFZv6njFAnrHnGHZvv0
LwkwkHQR2ZmRVnlhbQzoaOs13J2VoCuk3I5KTDgk6teGpBuWOyHLbyFe2S8H4+4f
H6XwYVQurjlJsSqSG5z9B+b+dpswbLHCdIb0bbg87KOaihntkgxWysCqcw1J8g0A
zkXrdkGq3zSWo86+xoQluIIPoBaJnk4E4OTSIwOF4NPm9J1Fc8xqTEjycJ4ZFfYh
/9ILbHDnSggh7S8c3M1TX/L4G6eSPIUqavHI3hGfReNJ7rKJOnLYxN+Zp3tacn73
EBZEMdkdNBAY/HMz75noDepvObgOCeNnK/N9SoT0NyDgeIas5bqq0OaTW08LMacO
2Nn+WMRea6mwvqDQu5kurcshybcQR6SOcEyIMy/KX6QLn+aCAQvNXB4+H4cbUnCW
gRRdQfjdvjqhuk0dSGyDbNHHifpql5W89eoG5YhwX29nn81T5mApjAAezNC+q821
x0lqTU4o8CZ2mAx7BCpIhVBNr/wTbNY/IIxlAOdGkveUhmmIaAx8hi00JedC6zZl
eYYuLcNq+xDItbEzif7P1XoBA55+fgguD9D8JQipPzvto/5/NM4gznj5tgJYO1Xn
m7tPGWdn/qcG8B1smjeXRSm588+ZXYYlyZRQeZq9vox9qItNaIhK0BSFqB71x/WN
5qDGnoGQRPS75Ul1j6IhB/kTMB2KAuyKo22q1tShubkOgyA+nGIoH3SBwYMTHYnc
E+aNEsK90nbkwLtoprgoV7K/dV8wirOc1rh0kEHzREHlXnzpK1ffBoc0Ry/0fzne
qnz3mUML/GbK4jnayD+1e71aM8eP0RxrYlV53tBl4fMBqfxBrDnlzhYRJvX/58po
etj+TOkWARworM7b72z9uuMAuaptLJ0r6llZCyctMOjiNr7CdDFT8HGLFFkmXPJ9
/kqY1ESxWL7h5CZFw0nKpK38rrUZ7Y1dHLvJplsQJufMqd+oqQr3aJpuPIoh7J+h
DkyKkZOzZNmHFcvSZy4o5jgYh0rf0P6kTosAqoLIu7aT9NAPqjBkYxzqTwuxwZfV
lY2tm7pgWMsjMGV5vQxbKYotGBgoTuOBVGR8rl66fAaYNt7YAsnd1hT2zQl0j/5C
K2QKsEOJ6cidau94TQ2jVl5sE/b+9wr3m5Xk4LVgoc4/qUTWUa44ywCMdaLJAFuG
2se1gy5/YcFxK3oefAAM/FjtCa7xAraWy5gI3V8qiGZdr8SfqTDCkrQd3HHbTNMR
gO6u6tLj/vJC9FcEhEEkC/6BfU8zGsYplMvJI3HRAImerzVHaV6SfVLrOLXshWx/
sEg8H0bSV73or3tuDuuQiAps8ozWJRJ00l/P4Z6kTRObB7bKGnQsfuAhS4mNvoHv
WSHyYaPW7ty4c7VA/+klRdlN2jX+olnPgJJoJL5whA5P+WMupQgrheD/AX8MhZ8q
1ibyQ9WKWFoQ7yOmBWi+ItuA99HqnMognPyjTGJbfsc6TuYfH/pIIVMemIGxeoXj
EyJWjbMm7uVzneDSIhgj6Ihoot4jQM/bxClbrrqRcZvbcQHOj2iet1EgExYo3eBU
OyquxfktKWnW+tB80p/mVzAdkGjFvB+zPYo+CN+013+IOhn6aXEmjvLnEbHnk6Gp
SBrYSh+Sl9F6ZKiCmjgcb7sHkX0sn5kWcM0utG16QGFgqKGvwjwOHaa84y5+Z8DE
BD493xW4E7eYSFm2sn07aV7mVmKxSbh3MFL6eF+Kjvu78uQWrAnbuUuLa+c2Po9R
6jafy+dbXNMzUEyLf4JM3o+d9yt+Am/Qb55IYv8XTxtVkZwbhCdPA74WKxLPoUT6
GxkdPtMXSKGUx5mipDeTdyUTeKIlplWcf6Jy0d/AJyWYu7E0PMo7bPDDgGBFnHX2
wxUvvaniqNQqNJS43+c0QzhkaC840zxf1iNComy981rMy2nIKCGSq8IR8HgQipNU
TG5Nz4dRFxdvI21+if5PkBLvYe+VZ2CqLTv2PlpysAk4UHr4s2YKOssGpJbAND7f
4PRFz9p0NjC/7rlNmguy3cAd9fW5te1w90Ws9eCIO98I2uSeI750yD/LiCFJFhEw
gyRf3ddA55rB0Vxm9L3Uhxo/DrP3osJGx7XMW4u7XjM63QsBOr1Ns2gOdDxCsJMD
G0hXmwcEvU5ZlR5X9NoRwLHnE7eY7KeR2ApB0plEqXXa+m3zn2XIZ2P6mJ2v8Y1j
9ojvfHYTlDLTE1yF41pZIkYxFhLN9F+nkPG1BruzegA+3/Se9RRBMGmSFBYgpn8t
He7LwDVPFlZpWDqIzZdAQyQyVjKhWapm/Cc5Ks3s6I4e+kYwEkO0DuSVtkFzE2/V
5u23nC0y5x7SAtY1Y1DuN5LK0gWS2JS9rFJ5XiDNGDBut6Io+KTvr3jtyrttuOGY
JEQjTKv3ZQixiMLhvgSsNNd9HL2saLiRfwhKwxFHLonMdaoPSskq4MWf6gBgmFl4
8pPK8I4ne1y7ohKI4xAulD91/EBWuKSWkL9Ykw4Z4a3/+pYPB2SR3KTi0kR09mqT
v6Wj474MJBoXhKI0Jl+g8QuT8wzud+7g3i9/cGy4W5LuAkseJAvImoTllKlK/q7O
3WDwVQpc9wlOPGu9DHW8YXvKgCOK4p8Pu+Pnsuv3FljDSeIjuEHUCuyoCZP5lcXa
879+9CVWZTWrR7Nzysazb/B5/Nq8e0MBZ+zXlV7fEPb0+NOz3sE8jMQ7vey4Ey7P
IlmtmcaCQCQmg7w14IyW/XQ4/tqwDuWOvq1M5lI4k1Aw+T/hgR/ur54TqZZ5LtKv
dmz3YIwpzawBNfPfohkqnFLM+sB+fh/A1HGOwAc377/cVVrQuHfdavk7EmnZNejS
TEU3dQRSOSWYCkb6p35qIQ/kGwTrZQspbCl9nZLwJYSPoCKHQ5ha9LuxBFYLBjN/
R81W4161LdnlOKzkyMAnMFyk6UjdqAGI04xwhB07SRTkDQwUogg4k8+KsqCezLLA
LtKHz7c95MUCP2eI+o6NAuj1Ec3B6+P4RIXPTzqYmWZwAQrI4BRV6hCVPK1xpAFZ
jR9zrqn9aNWTIFLIsB6rOdkMoo1IAKWw8l99HdfE2/Xzh8SmEo5oQNVate5JdpBd
UrcmLUpSsZOFEPKN8HTxtWV8FZ3iO0oHexiqxy4wvu3ssEXhWMrRguqmxP8Yn5iK
WmCJTi/Kffu11XDAUVZwdtD6/2EQ9iQE6ADYmZN13y9frhXWhJTCE9jC3ZCyCQ4f
u/51vJ6Q5/vbsuGhNr5x9dmqbYFrCgZ0zTU16ebuqaI5abAQVQCqLN9oFCuTAf9S
k/YsTpmRc2Dag6F7baC0JjdTuugGzmszyqQrHAv7d0wMpx8d/ESuzK6WoHgCqSD5
osnmcUX9R2opGLPT2nopy24NZGxZoJaHU395Pg/JRaChXvxFVJu0AXMIYNZplXVy
EYuHVF4X/I0/tBAzaohDB4dY1P3vMpARwwA/lpVbmkXGzfcPaZVX9qFbt5gf6J1c
FOmPuYhTfXWA49kzTINJxEmkklmGMfYunKEeCJvGgpXlkeKDGTZo/jDUt/aoLp3D
R0BEbwsKxmxyQRVjbGscfqQkCsq5n9qy+LrOmQiNueMzztLiSmYAnRZupAEud2/0
wKcTDiuyFnukxzpdJjGdcXJb0xw8tYWlbH8eGUpbjqJ3TnbXfolTXe0nfhhmfdJo
1Uy2Z9U/qNcl1/pEM0tsQSDwR8+IMRM47w9kgZGSrlof5nAm3lbwopFCyZgzust/
mFb1Sxf2mQeawB6gqfrgrwCYExjW1xuMZ7d25Kg4eoAIbXKCrjoAuUL+c+Lqg6Cx
XMj/7qLm+RyzqOvppX0cv5pns7wpXM/IEoSb50AS1nByfM0PvCs9go97HDsoSY6l
uliSffpouDlifdjmkzWzTh+XrUnma1J58u1ApE7lAaOmQSwHlCaDRNfj0de0II1w
ibJ0SzCujYC6ez9zF9fTZos120dlAQeRmXthW1+5mMRAyWlA3XAj/ziXnL0tsOp1
yrSKVz4Csc81w9HBXx29nm2TSITdFcOSQhOTI0D2kW+LhMNBxbnukQ8svh6hW7YW
ZniHPAkHNe+jrUDFwNlLa4R+7wIItjhPcGrGX7E6wTUhJYrb4n4SxBI23T+JioOP
vPJPUxzuF649qEm6VWxZgTW6mGLLsPpTQEfDeYol8yqFUeALgqVJj7wgXluPY7U2
bF4XIDA2tX6s/j5h4xO6acEQWdIXjBqaWb1qvdZbPwBEIFW/0GG7n2hUdIommPff
eX1jopJRIRIuHK6eXInFEYaiy9ghqH1oS0xKHiaDeJ1zqAQTlAZbqOmd4KWcbVdh
38827I8P+SpEMInC6MsEMAI3pRk2n4sTKWigLoYOncMWDOtXDSaOw5Hpn/W7PA8Z
AIKS/h3DD3smgOF2yERKYDL52XO37QTsHsHJfSSMSx2Jd4FHgZs4HvdfSgJVBmL8
u1epoYvUizRAKsjOXuwn95+cj/EFLg3EQO3UW7N+1a4PkkswoAGGof5qA8/kbMnn
/+3xKrBTe/8Mxc76TtUYN6l78X0oNKqxpBzSCpIvlfXwdxVJmOiXNcpFDkq7fVRN
YNaJDE38nlvoN+mXphrzk4z6QE+IDY5HUXPckmoes58NxWv3iuw5Du16a6nDzZv6
Qm/L3CEIr+L9d0Qa9CGffoODe0/l6J7iFeWHxz9NFVNuGdwq8dS5fu/ULCq8UgKO
czmW5Y/xfNydyl+5tJCvD3/L7pVXckD6zLn9k0CP7FuJMDToNH+DWRRedNhiEp3P
ohXZGadc8n3M4rTFmk5HJzUYmmpvAy6h9WUqGKBA0XorUhL0SVDYLXIDNi1WCSfK
tW/fJRuG0LEGQeuQrkKR6mju1cwN5lC4BAyDRzG8K7ZZwJ/KwHETk/VFTJPECpQO
YIu7p9Oc3vhN52fgqNeCPklXv4ebBt2CHyjUgM7zRDNbXllQXR//ym7DqvdZ2r1F
KaA5FHwg/w0Kb8DInnTH8QT1a+/r/Wt1EN9UNj7c/L6WtFe0xduSaLvZpl2DE4Tr
C69aJYgjtPPvFDbEGKjbwIHGKstBcmPddGNuJAVD6bpuQ0MyDTLP+1ruljbbUwJo
QkOaJGwGYHhih8/eNjkwH6y7evuDTG1th+OyOYibQtWu9W+fjYBzBDNU7OtQeSoO
R1RVK8TLXBTBO0v2B+VoCxG/FP2FxR2TFXOpJVCcfYCgCYVxF3svNUcSb7ukb+9X
JDJWQAk3tq7n4zEyFJO4KBqI1ntamWPeHFS8VWNxrx0MXaMKLuPOkwZrxNh4r/Q8
B4rAVYh4sJGmBNs90wf6NY8Z95WDo5gI5/OOw9SdD+Ua8abwmeH51vMGNVBIP+aB
9Vd/DxaWTIEIKMs2vioSwuk6ejsYqnF9umWzer68v/IaUnx/pz1721GmJrPpjnKQ
JrDZ+yRr0UB4wAdIXSjPLz78EjudO0Z9+ZJ/gtOKttLl2EsrzoN5HdmVD8tyxHFg
rypJn4B9PDzz34oK5QVTb9BA1lLXi6XlkLje3/fRiPe6qs4u6M22sidDUpQtMJ6J
ejmj1zD+TUPq+U18XwHMcfQ1p8znMMV3o5j3qMK/baUEsm8A1dkOCxXn8HJa+cuI
ZeKejM/5k3Zw+tS0T0ZROYez38MXcil+aZ8KWI7+o0/7Sa07cqkzsmLxPs6P+3R+
mJyghcrMkKOSHuygQGsqIUugfnOghp8cKUfjoEBtImkPNmXH3Vb2/gUOVhrKwQ/b
vv+OJpQC+SA52Jamqv05PLBSXV4VtFocwN40THCBC4oHoR1NVL9JrWJAmLfahzhz
yZ9b1zrV/RzXEyqpsn05AVVwGe2+SQiahTMYZTz1vAdoo4sfhMpgQGvq/JDOfHVn
6QNnFgn616QeMDSa0MTiS60OWHi0ieHLKTeydBkCjy5yNG53Jew75v1C4UIB7ZfF
Pf0QDqXqDjFMKhA4syNHMQJnRPp8bXxK8JP4xKZp5YIvVrKku+ytbibn3bYxWCdn
Oan/spNZVAbkJi69RUCZayXAVm5BgVfohFTzR6Hcyz3pAHAy00CkH7YpuEVDOFhk
sz31FZl362B6/AcZbQumvi02M18qY/S4AC5BjcJuCb2dYLVb6jINuqYQcESgQNTd
meMEuID8+iUwX0NqIRDsBioe4rQWOW3i3kcLTfZ7S8HKqtNMHbJ/aQCyr2EgRWTF
0Zk27wsWLEDegmOEDxLXcQsWQo5LEbVEfr75NdLqpxQw4ZkcbcL70HSncCsKgEK7
nKvCCrP6KRrOrDmSB3zr565dSKjI4ZIDzBR15MlVX/swYSpGQRrSb2LDVR3Te4CT
FDAA9TjDPwJ7u0NjiTZWquep4+kE4WgG9vPEoGiHjBOus4MUyoqwOhyBuUUtivOk
w17dj6ija3UjgzJ0ZSqIOc653NSgy5FBQjC/BGKr/wOwVWsjiszLf8LQxtCbggwg
SImCva7/pNTOBA5hpLfj0ShJqX9dDiSpQJr2Fpq9fA+jE+IFrecMEvTHoHdzM3hk
J1QW00sCbpXj8mxF9yTsAqYlo4RhFkBvX0AKiRdFw74n1xs3DogQYdePvhDnP7vu
gQAzTsHf8/8WpRbwfudQLsbrjIX5J6+N31bN4UcDHkcPF72OP1qyWzSvNwoZDKl3
k9xcmJw+6kAi/EtF6t4Bv5SqjHJDJYBXFZgWF6viZ1VEbvLPDjQ0JSjJLEivZTtN
X85DBNjtWK5u+pAXcxawrPrbLiZzKBAGN7Vow89ZN9217fhIzrhcgnRHDDoeqCPa
ffbVU5cew07f7wU6UBKbq4LpQxNvdAGAY6iduIG4BHwn8DwIN6N5TDareJCjAZwI
5OPtf98Hniav+5Tz47Hfz5UhxK+s3XG3dxqk0b/vqbLQA+a5CzaUYscsj4t+V8Cm
Y4wOJIDxsuVOsT7NjShoZkxDc4a+3iT0fHgXkdkamqc4qeWJhvXjhLk18xZYp3+e
c2V8WFQZrzEJeV/zfhb7wLev5ZiYeUbTKyF8qcJjLN0G7J80sQOEjYoYCc78Rrk6
7J+Hd1uc0NYZRG15GlByCCKt1LMh0K+0opPd7bQN8vkBs5OcsxRX+4fbDZeJ/PUn
kcVNHikeKPfxG9prtdjRsqcmZ9kAYaxKs0KXJhSzzqeJrgnNoBl9eBZR1GP2rlZ1
91vlET+j6g1z0gL64ATVim1xw0Hqhfci1z3Krc7BkPaeTwqABoJnbYQ7a+dwWh6P
HHx46ugMDLLAmwFd1XqRtLXadSkjyYwaFuHkCBOZQvOcjLW+6RYfhlgzN95gIwGq
QZ18AZfjsJJT/pqDWU1yxmkcBRPzUfFOWh4LeasM/qoD7UwbdTIw+OznT3bJVx3e
Y2SwBAH0N5DQU4gCccbBJ9Ow/HL8Y9w+NyTkO3KHmZOpjYlQJ+xw32F8kFwFwrM8
HOhKeuqgBpdqgD5t9p+dkl5oHU8YGLni8YyGsZ9NRA0vV29Zoq3TvsN1HnbfKOXq
PQxeyQDg8G3O6aMC4QGoWwVXn2vlEzrFvo0+mfkn7rvnPWduLVbuaaCYtOy/y4Ny
zdLb0icLAG/CQzxGoHq/a6+aqJQqllxi63Sfbrrcc8g+XGvBoY/DYYwdXwaaBWeo
pn3jIuhofHtOHvPizkjmtzrt81RsYaENUTZmFrlBzDlt3+fQhY3vbpQeuKyZ13Hh
wMZ4r8ta/tET26MFIWcZOz7GIYwFSll7jFc+ObvzZfQxSD0wZmsF6SjmQbXYlzKM
vSoVDBUATMLvT2Fd5zsT0dlzyNy/RnU3hEyJw6Dq3+sUwnW9ZIr4tVGr/nVeAml6
/skeNncCG03qm/kySHAtIQkhKG1u6AmtISFl3DXxyU3a5ybgBe7qJC4ZRaVnrZgX
hTN/xFK7mhhw782DDWxEuozt7t+czAkMUEVTAMule7UmFcVbn/QDT8YgoDm5kW0+
dRr6khtgr09uNYRhfuLF2zStkXFF5VPt22Rca0m0hxTrhOfrJ4sdZSxcS+l810hY
S3FWQLu/CH5ZLIknLT5cjlgUw4eVYnqAJ7C/7Oh849oxP4juYnd96eeHEiJQJV69
ab5KXz4O9FtxMPGsrSk1qlHy/bgxDnxu0Ya94isfJGmO1R7kQtPXJosuVxLiu1/e
MIXr+3+dwcQkuqqmSeXsWoGLtc6vrBHmqfzBGdQVXekjhnMDkmQNl4kZszFk0pwt
R9EQw4qTDSccqFAPPZkesq5CiuholN3DVloPbbpD15nE+gV6MxemqhoXtVVPUt9c
vAnEbeqQAQuZ6Ojt17NKmMlIX2ZM9cxuN9mlqwrxCHL03ZkjgVsvjUxVSZzIT5NO
WU26fJljqCV3D4RYR3Yjqm7aLyM7Z1vrEbWCez5hm1yJVUysfFu1ETAsu1R/NoNR
U8S/NhpdIYEkfGNc0cBJo7GpUj383SEBjwlXfkPbiG1cpcVeeY4MJIw02ERDDzsD
xjQ3NY1qlaADLvXLH6JQtZqhUpz7ZeNnhnYIBW9KqU5UAwAlMF6mm17srSfzKuSB
KgZZ+g7TGDvs6oFOdj90l+EIEV5oVZlLnfmKUYnffM71BOR5e6E6vIHYPbRiUyQL
11pdCUGyawkPbFlZ8tDQaczT5QsCVXY99bkt8AwzRLxcBRd14b5lEZ47bg2TP511
IaDaqon9AesuZRfm0kImiGRqeRtQiBQh6eh+HuGIaQS/F6uNM8tLVG4lPYAgf9sE
qpM2ttEszkLmCgfmEuVkByxg4+AQZ2leuouSXZ1LR0sX0tMbVMZVhGwEgAIPHghD
iYKyg/olyjF7pc9WnZJ2Diaxs0ZlLWO01g8YyrLAl2r1x4NrcI+SGmLwWkqfUuFN
yEwQ7vpR7ihh7erNcRKSKMXkzVLQVik6q/WcYIjVsezRqu4xVlW/U7hEpQyPgYNe
cxZVL96g0SkFQnbRpehIa03Pie66p0KXUsf88ZNEzp3cQYpjbuwvLsJoGFxFRXSb
6sQv6j17J9mSfOD0xokXhKyxXbZEu73YTXk+RaqG6oQ0UIRew+5VRn6JGrTTENxR
aniN/QL/QtIqhSqE1BfksgwWaA4iHAt57J+EKFoWn2027ZwZSS3hv4f2GUkoy7or
n+njD02ypEJUj/+eZSypqq7RNLKiTrzhZsCI0kezn6pf0bcil03N7HmoJyW7TkQO
Cl8x+bsPymk6JoHmt4ti231bH8Ko+ES/9WTsJGWPkZkoLU5c8QNLnLO9UVbYvtXt
zbsRE+TXWR/486SevSKJSXejKRLZ2/1M4hNn3BwTtCKL/FzCOcJSo/SxOm45k5uN
dEnbtDYmUtB0qUuEgElvVw9WcjAPOBE1iGDk3yz7VO31FKbhCgvZo9R5t29/j5bb
z7eenioFUZClJ+QL0HVeegqAi2hDJOtuZNa7WahtSsR7llglJEovKk9dV6b3O5ty
BYyO8ijGFvGlKCcsqE9Qeh++CJYIUZgZ8WGICePA9wVKRm+1dfXLIIdWP0+Rf5oV
3jZerVuiGhOX1Cwf4txNn7FI0XfJmt+80mekAbtNWNufUpWv2FJ4Ch14uobIUhOb
O49RcYJ2fkKrOEcfNj4noxt1kRa0vhjiPC8gAqCsgg5ljlvIAtSKXw6CU5DBb6Vj
y0U1LXoAbbPS4K5SugrPdlbctso2V6ROG9Fg5kYK3IX+lT8rPmo+HSUDTtmy6EW4
ahyOQ59P8QZeEqol3vVspnkpjTHRNxwhfxw8H9QiXYRnp6Cf+FCyeOTEXYjDgNzj
pLUiyF0pav8qEIFlOZbdM7OtwPMT+wlxcSGZNpCkaf8Iz+VQUl1hxkDAuhPa1zn8
2VTPWi8IrXkPuHGw6yzqTJytuw5sXV1GmWxicEDL33zPCkOfnBRJ6lkTSdcVZ3Uo
VU9VIBFcXk3ysNbh1TrY//8lM3SpmW4GiyMjfFz4updDGpE4+3FSDNCWXFmOFBow
XFw0bxhFtro/36qWeGN2m6SbDrpokrwM2MWgoSdJXXostkpK0WG8gvwtNSYvxZHy
GQdZ9r0xMNr/WNAffu0+yv87zSiwNsbXVJ3YD9suOIT1rG7ZgVge1ud4x+pZ2pLW
RdbJlNb0FBz0UViIqNLYeuyAniubfQZOQcCZJqHghb4KWkWNI0aP4F3Np+60i2wS
d7+FR8s4/TUkrJGW5Pj0qihTOBakfaGTeeaeCxSzhw9xLiQrSeiUoaBUdJ4hZutQ
9ccFtsfrvbEaJAIARcQA/IA24l5sj4v/suNPHHRCIOqfYwFx5uZ1tIco8lHG7B3B
igf8UvIiVxvGHhKmLX7jPHehs63AzydP8z0n3vroONOWEVJ2I4VUt//YAedWfw3P
+QfsDyGqAtjqNHninKnpabNv+31t/flmAb9OGewUdqDI//GsTbgi54aXz1XuWMus
0qAmXlMK0Ot7Bs2W7rFiJHySNSh4ltkQPTTAJR0A9DvkdolQ0J+rwyGy9xi/Ha5r
LwREN5TpzPztEyz8+zuodO0EjLzRYAJAJ5xOBsxeDIQlu4ZQcr/3budTbtQYoLv8
O/yGXio/BOpxtG2wVQqR/xISMx9R5HlAKGalggF2vtv1U2YUsNV0h82UubGMWmz0
nZNmTyc6WyjICpIzwgShhgaHdjbW+1nMQdhO0btnRf2Nv8ma6jYxqNEkICr4AW2y
Jedyzkom+tPRZ0TMZ0D9mn5S09qoMtGwOF+HwPg7EiwkGmY5c3aLRQMe2t4+6t0I
KYjF2Xgj7bjulow4nqR9V9aG0ojKZtmZBtTtant8PG4Q50ITrDxXMU65Ti+4IKde
zrVUU+twJKmrqQ640HiM0F4CBgWR6EJZxGWYiNjDesA11yT9cmo9EA1Rf/6cNCU2
s72XSzDPVX+45xpV+pcrD8D30IYOdffy+zMefFlmrSAXiSQP6L+L9hlmQaujYjfK
NGZ40ekYP2QKKfE+kYj9rEtF54vGf+LI/2eAgWeMI9dvIO4ogn8VQHWRtfE8okiK
VkfFHoFnxv2ae+oTTefdJ3Tah5S9NZiySevgg+qeUv+A5LjnRFEg0RBaoQrhTSjZ
tgBpMWZzafmbP/B+GNLN7swmaa8xTJL2UFgyEgBb0j1WtvFZ1luVy5fFoZuXkpGp
JDwsiBrXp/93oUAcEvIugGjqvGWQkp5TU90kjBruiInEWagnbv6fUgbeEDf74XpF
MyfDXbwkzSexxyhy+D4p9zjORNgoDWMEhvkaEso+fjLBeS1ycV/pgYCOM53v6aB7
JPT+biLiIVQzIFZ0Tt7xJe7YBJ4Q/ntNkGIkPf2xYBVzgrFO45VZuWd7Im9bodq3
735fk6RSFlywucN4/glwxdLODCQ3z6+gwaJF1dYsZuoHvG5TOSOXomMXn+A399Nf
jjkG/j+MAG+Tzjh+MaHqv9F79pwFrhTbILbN1sTyGVXN0AyVnXJ9cEz1Tx/m1Eim
+9Ymmvqvw0bv8xwSUrjAaCruSCQOSXf2J3TSUFB4pmVBBGZVYQcdbiDS/sJKuItW
atCrALehzuvtRq1PU2dUthFXYjpFpb3YeNhg1J42IEwDjQrYZVqcaGZpGJ/qwKA8
B0Km8wAXLj1yM53a8/IpgwwCQW7o5z34d/mM3+39R7hrvkEWR2U9PwwwcLGS28WL
yLo5325PM6pBvzHX5z39w1Xxstf5EDFjHCLMl6qh8fU2ATTggKPgTxzHHJgmev3F
GEx67vaKXRey8aCNM8ch4cWU22Dey//EgryNG1+nupyaztAfMtsKzMVowDCBYR3h
Xz9CjfnIPavAEvCtPMWWjLSxrFotDCo/pvLBdu+riuwEbddfTLROyh9v50a3lTkD
qiOti22uAUiA/vuQGNpC31hOgdFTvrmU3uVwi8XXhtkoj4R9ghQMw9TrPPyXdxz8
BIHPSKjnUOCaQcYekA1Oqj7FIdXaLtSEQv0rmfvC29N6q5M2UcKWf8oS9fbxgwT+
/kQfUjivvL8+QAleKnnf/V+uK5cTjxVyIjiUFCNY+8KerqsMp7nJt75Zn+UmORpv
zmH7/s4D/VvhloVpybbph2aStA7J3gQ6N9fsXKvPZhJKEMGWIZSGxZXC4TlCwp3B
VIwew2c6soLmyeODgY80ohoNJarofKv7u3s/wyas0K2DumqBStd601wTKl+gpkV8
s7g9IdrqMRNvtJtMRmGC+LctLig4nGOvYfg/0F4tdQs/w3VYOLBT5FffXDHqSaXs
E61DXU7NnBYh17WR7a/q6icYGfIAlNIcgoAZkVu7yZ+Z0xiTIDQuJCgSYw1i03j1
iH4hWEvRkcV7Lq7+ODNGpXBU3YLWt0c1dQCsvwHpjc0jXYGbX45ytx+0mfkSSR6Z
GJC6xxas3a1ofb/48Bt6AdmyeK8y4jpzkDk7Ynt3Pd0rDDL9iuiQS0q4dARET0rC
EItU+t1zsUj3bJ+b33aAIiTDj9aLAy0xjzyho7KBh25Bf+084z0uXBaJIuvmpA3Z
mQRHfTubZJxhXPwA98HV0EhN+Dfrzi8Nvrqsn0EJM6vxvEpp+SFZFuTUngEIx16f
cnUbC+igJU5OF+KkWnzcM2sV/ijwOfKkqH1sHeDPKdgS7kZwDokiAW8YDgKFF/Sd
usRjafbP3s4wToj1t9Ck39tkDRP9QWuPoAnK73yFgzvBK1mb0TH9F557wN0zKhPw
Yeg0KlD0dncraG6lQDuq3B1gFHMTq2Rn2zCvVhksIfuBa98YS8PPYrHPiY0359mZ
biNEehLUU8QJzuQtXQTiisUcZbLZSBZsXbcaj38XGwGIF504BxtAcGsm32wTVh9i
rtvMBrHmwNtF8yBDjCngSuOCn/Q7cJ5qRg9dFvSKbM31ku8gNIY6MCMTzO9pU1E2
GC5jP3gwvqkTuMxPt3z4jVALA1aI6zGLuad/pnYWOc75lwUpPoT/0y1MsVdAgyoL
OMEQjWpxMcodSzBYME7Saqloq2ZY4+DwWoPpjgwPH1TYTl+yEGj5s8UHhbEiXFIR
CyIAGNaKr7tYzgusxWE3x79W42HeNZIPRqj2iNLcJS8+2UHdCKB0t1fX8+JXg8hI
0o8I1S7iujZumg9Ht3GbtrkY8OsH9mXBEJ99LIuL7VlwMiBCrwQJLLpYRbddqqTn
0u7ikEGnDWn/pvRmd/zxHJS3shENCrFHmJb8MIT8uO3QkRS7htm1gJhfbAUjijrp
c6jOpeWlIXv5Wweu0qnmT2Kor5IUKCyvlYDFIyO2kXjRo/Bm6LwhWPOKwXKCjuHM
6Z47knn5FNlZXFdfriXLEBKrMR3EXvgFtVlMQYAybgZK4fc4eHphhg3XPgAXCHDD
NMR/XinuCsoUkO2WntNwt973goTjU1O9Ikwiw7Q/yutRuQjg6zV7+pIrP6JQLhBt
yg0KIMELAG95ghk5R9NESxAGVdmN6AMJSFBuG6crnP8HJHzgHkUtFxizlDqSJ06L
A82l7/koXmUPKfPkrlVoLdikoXRVGRPoI+wJiBVb1NqLI3K5N1mH30X5akilGafJ
xcBcFNsZ8XohxWvw2CoX7zwt2CFabAo6bWhKJayaVBTEwrQ5NLJU7XDFrs7dszy4
/+soCATa/bDDBpFRUjdxWmX44goY+B1n0z/GXsX8Tb26T80Grx7Exns+1KSAs4Ba
DYTXe4u+8bt/gFoeUMSJEWgwbKVhlnYcTkSR9Wtb0e8ATON/9FFiUxhXwVthO0LE
wNmRQgcm/3uEzprhXILi1wNsgpXsael6SzDpYbhccYccHwlwM63ZFwAofeBUUkaF
g+dj8PFUjmvosAOnm1ZGv8rgt575ZgjejqtvH+lknOngyVqyAi1HB7PoEq1NnD9t
A4jQ7fB8ZMYxEQbpZhjWBWCYAzJBwrlE1XTPyuPwo0E+TpCxVnZynXVGeCDi220e
0/uxKcHv+z8i+IPd+tq9+O55pAyKpRrtQyW9XB58VNm9proKLy8YaOMZWrxuPAKz
S55njlpl7d9bBKIByHE1Q4SFTzwTPjkzvQrz74Uk8yTEvLWEvKhMS7Ebx2bYIw4f
cd652r7GPaf8mVT+R4NVEl4IydOB608/YPW9S+fSFOHkzT8KVmmMhx8wOvxBvpij
fhUOeOMYi+wBSqeijzugPO+SvlczTyt1/KYuGAk5nw1gCzDvLJqjOhiH/pEkeKC2
OP0CsJVFyBqjaoaG8Z2DWx4Xogc0tfiKdo18YE9+S08Mrf8almlwfNNuYJR2RQiy
7NPJ5onBRfvga3/VyOFuJApOSxUDetz2bSn/OYyQhM6mHo7aIXfOXbohVulmhMIS
+yFH/TGEKDaOeNuhceIg9psjDkDlRAAk4KTbHZyLoqmrfv/3VtmuTTqhnQZmD6eL
8fGgJMkeqz9FfYwvWq13VrrJJ/Bp9rtLUxpvtj9CY5xloCX/0RDvseMOt8m3QAkp
ohgVgOQ3vcyT2jMQ+LqWACvVYZReg5VhMhs1PiS6CBWKNrKiLCUgCeJzB/2laj63
+O1L1dv8OloW0bwPGGV0QxTO7lC5d1/iKLdLC87kKnZ0GA3vVYtoiN9LPCgfqqSC
macjknR+HsK5vqw41s5uTZOZ9UsSCmAggCbZ6ozI+exCbmUIDuBCEQbi3lOXgZNv
pS/7m9LhZ5D57eFXd+7dwtL6dWZLlUoii9Cb2oAE8dnJy8HyGDdDgCwVhd7iXtFX
2mwZyAdnf5rv0GZqD8Q4J9QSItQrW05rLITrTJrd5xfRB2dPJJURfjsa0NF0KuN0
y1xUbL7Ob6ATUMojLG3Y4jI0FG5QYFL1AT5LlSkCgjHInCI+XV/fd/h+lBz6t9rH
206s34CPyxnuK6CKnPy9O7+WLXKxOrhcbmCpXoHcHruedyp2+36eopKBbsHPUULi
VP1Qqk3mQy4Bs2BG7ICQBHaAVcLvWmYfI5thbikd6eNNa3PyYqX6Vcxe9kLffP7B
WLlNVeZVv4uGEFtUuuwr/KJLyGzW8DKAEdQRNHfBvlJD9nFlhvbLf7frjovaxnpF
MXDjZ/nKD9kJHbfr6rFdKUIXUjBUceqE81EI3hCzOyeWaDDY6706P9b+bkxnirwV
VKT5OJY96wrgv+ISo/bO8Ip7LUAd0ObwMtjVBdTuZjxnetoDYFXyd5p37WaESGWZ
7pUXWYpfo+W4M82vGTN/D9iOOqiVBbdx7e1qrMyhjFhuVNscAPDlzeGejISQbO+8
UuiANaEtgEGIxPVcI+vzrz640HZkzlCtmQOZiCbSIdqJo0OA4NaV38rsnAAAupr1
Cy8zow1aQV18ySY8y0STphDKDWy21VslsA5BS5Ep2/k76fyjxU88w+X4Szu8/AGl
Sc+RyngQcA3rKYeS5L5dgbHJ2HBAbGCCyNxaD5/pIerpcWPiXuLO636bOtujSSsN
dYBv6/SUyrsX5fAX+6MkWarTIUcK98po8edIloS6zpaNOWAmKy1vHt5Cfwqk1Mcs
yPij4dG3jg7AFqPI72x97kARiCQqNVYaDZpinNLLKdF84jPcVkvB3T8VC/X0Uruu
4V7dmG1LQz0ydVUSv+pTfl1M9dVM3QLHMQw7oEgo5NEprUaBh/waWawWKoQLjL9S
jmLc+8KBPGwArFmpL8hZO4Lf6ljRlNEeO9q16raU8YerkFiMspTitTEkNvharJ4t
DrcMPuM6dBkEVbm2ucYX8KzLirwICNVFDVO7fIjSuzuh7G5JIsANk+47yO3CSSJs
Aonh8KnBmk/qBqGolnc+KCCxSMJP1m6XQnLUW/OUSCDztEnkCXlifRv5CS7LEzJC
E/VUOJCnoEkIcd4YEtpQLvdcx8A2/um2q39JxYZOcz5thduAXNvJADT7SdHfIDSu
/tsKnGScPrsuKD6us2IYHTXJzAemUl7xYHa2DYtfNjwLodG2n9sGDRzQMr5n1/wA
FiL81f6hGjhif7VyrsSooLt55GxvKEkzMI+5se14upNVDKFMX3+0NgtZA/JHeRPd
0iufxqnV2CEtTf8BnGE+N7Im3o1Cc5AFaqLBU6G72ozZl1czRwUKM0hXSYiVzc7k
i6Db5R91FC2SmQngsxxfv3sf9PkWP7KFFKxB40O0qo9RLAytLuCyKXdhnUZ3JvW1
E4c2MMoNFQ3JIUj6BPIb+6GsLSyICVC3x35Om6sb8k17BGOI3wZJWHXedf3E/HF8
UmggWO671DaCxfg616NtowVeLDa3NwzyGiXdNpAUW/xP0wGTIAHVnkd6Ubf0zLHk
lGbq4ywNAmNu5p5KGJrZIokuJDDadVMfsuY2bhMhOf8FqHdwRFp+1Ab6dnJ9/PW+
ImKJSijrXSiL0fuSZHbAY0pmfPt6Nd8y0xzR/jpT8xD2WMFI7mClW3W2EdHswafh
Q9pylpbw7xTi0y3nwgEWA8ZuiFcZvCAJ/W/rXpQkKcz5Bqc0O1ZkDNwdS6PGT6TH
KGd8jSUVYuq91LWIvJuecR2IvVVHSKD1qdM9fO2p6oFIdomP3BR0Y5nKKh2oDVHq
TL+aFl29aSA5LSAKv36gHRE6+hAGS7Fn89hHrjILT3L8po0lJTTwVkvRMn8w3O/U
3/SzrEHWrgsgENkr1SEiL27fsralbkQWdzUZjeRvu5HPoYph41FPr5OwQ23bSTjf
7JwHIvzHHE3mYjfoi4zKB4OZwSjY+aNZfZnDA5Si30P5fkzj0HYRhuBuPIkEVANI
9c/VwlodQHGIr+gjq4f+V1HvAmNt+E96Acye2/VdVX8IOZyg/rtaP55F8Ojq1Lz8
3IedPwLoYIpGb+9TvmHgcs8Temu3yODbA5bba+F8NVyQlIFsob2QC1XX87yKP0jU
6sVhJVrfoXMUQf5PwDGocNJJbymLT2NXU70IK1mPpyUV2CwtOJ7NkawGpNisylSX
pz8zYw4wBHTOdnKSaHE5YRWPosHcm4Ta9IBBJyKzZY8XuIwyTvH7k5h/633XJGsJ
edDjuIJ+NN4kKmd7TIWqUzdK/FjkUYqcPbUTYjR+zlGF/sV564bv+/iS9JqQyH1T
1JaMteLJY4pr4V0zl52NocXSoUbWOTK0wLnqAjdDF/8PzF4Ti/njhxaoXTeoro3L
BoVB/ZTTFbuhNL+NvB1jdqe4fe4tD/5uXxRmrnO4f9xizh0vJ5uo/aUAZZ5O6esE
kQQiWZRGhDS3Ec2+EH7RAZ6TRx7REQl6Lf7y8pM3BQGth2A663bvaqeNTM/Sl0/C
zmWDVVIRdOVAGv/eg2UT4e1lAMTtJfWnI1CzojzHnQJ0wg6ljQ2hzlEP9UEGPLT2
yqRWhUbdUe43CniF3aUt01JzHGthUm0901vIXAJtZbZI5DxivSOCTng0bB64R1l8
5sPPt6Hcuba+/O9s9WldnTdDjsVmuzn7r0Cil/h4xJv+nkNNcapGlFSBDgzUm/MA
DHP6qEn27lejQnDbLZbEP8gux+ra+cfTqOyyttDkCsSqSPE1/Wk3DuJ/aCbVV/cf
zaqAKC7AKFmNPKuMFSPatVrvEWUrnQ3/GwhIdgjzzNSZVDc+cMob/ZAJjfXv97Xs
+nqzNPZBE+9wVob8uOEAtmvnWUWiaLSNfBDkYIrOkJQ0cdVLfzhIpMS006pctdXU
A08q/iH/VW6qcaXYUB0Yyd8w3y8mT0tbRO9FcHTAuzHlraAhAyjbEjj8kuYHbxxt
xuQW1FK/4ffpReObJfkKaR3Az3mKmewercd0BoxmQU3naudruOdhhS+0NNjLcWyA
sKjjzYeTg54Hc5FCWjDqQh7dI/vUZMxrZpd3XNvTcsTAsTOrPhQphzUYY1EDmjQ1
JJkvtWGul9Pp6jEjE4ZrPagu9I/LUiHARbsiFpjQRYaY1OOY3gbgxUxhGbgoZPpO
4wBonkacz6u2tjMH+2V53RJ3Ruz3K7zeduYI0eKGPCy0WR/RFvoII6VkPZS2NrDt
9uxqk2b9NR54lNsa96Lep5cWa7qW1ONdw4tWWbdCt7jUXYFsOq7AGOzx/YdJBnxi
U6UIA5YAlIChECvVC0Rsww7lozm0bfuIF4n5BlLHWYvhM2mHp7v5mQe0M2f2BueY
g7SI/5mQtRm4XqxgpFBlnUZgX0TyaBaKk1NfVL82ru+VSU/YxV5oLeSgwybaob7E
YsMahvY4E5lGKg6m3GtIVBjDVCeTcO/YF/oSMYiMXR4/KwwfXFlDROJfIPhWZBqx
doBWxART25HJnOJsmz4nTBdzHDhJHiFdteovwTeu4NkcmlISt7RJtmSm+m/d0f/c
Im0RxYJr/xA5U5V0l3YQnQcrGdec8KnGCZtV5qU2dY32qrYFlqhkxkJkOf5qvuP1
fkRuY4TNu7RhihzjJaw1w4SD6nSTdHYnoxsk82VNPufbejprIvsIEWq8Uq7VbQfP
ZNN9HRnH/HM9gKXmWBAP4v6SJf9nfH2Yl/osotKxQViANjsh1f/Fki3UdTMg0xqi
pGPooYXwMNGAKYGjYe56VwdCsuyaNDcZUQtUa6faLssDCBb+3/5T2O0ldVMb0RPt
vE8a+6ayZ6Z9JLUaUsJEUYSXZ9DiJuWcMAWqbyK74ajP+dTWPGZiA4LWn9dIFmXl
oGvfOWDxSQ/p/HfIx33CZlvUqP/oMThHtzOKGdIElKbhyViSWBPdtB/QwCpIwiGp
nX1B3+KOwViuaHwOLs8iTtI6HKNNrgHRg5OxqzHSPm/4rzJzccLgwfSXYh1aCXVM
9iTcPEPlBUGbuYhwzdGGVHn5ULruHL0Ek6qAhkHknDYekGU1FHGQiFmna2UqzEVy
ebOCrorS7OB/9W3xGJL99BRlIndWxpzIBnUSbbwInJR6aPhkI2WjcofokNC4CyrR
E9yUWwqAzAYO+fSyfPLJBQdNGQlxQolLM4o/T8T78Bx0+f8NQZmdSeAbmTs4Dk7t
46pi3rHOjydS+e7eDSPKBZkeVqbteeaeUgaS6QPXR9+d2c4qbzmHDwow8bX7RlrB
/nQ98m69jYNV/T/arOh3qkCvLGKJnEg/bFCrKHdxUpYY9+hoUbdZ/EvtxULIewqo
7MRqI5FQhpwZE4VXOBKQj9CwpAqvaMxVq939q8Norqs=
//pragma protect end_data_block
//pragma protect digest_block
TE3MkYBdp4jPkY3ifP28cSwL/KU=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Vv5xibKNMooP+JQmxRl3FMu+QkSVBwrEjMTiD2KbQc0d9TSwdZVuWAmETw83hJoQ
ILZP8ueDPlLY6B1mro0OSRIk79a1BzK97CweGvoCe0+/SIPf844GkEK7DaVCQd2U
eZ3T1/NfJn90HaeuJTJIJVB12Lf9GLKW02c2xyyh40HMaXnof+zd5A==
//pragma protect end_key_block
//pragma protect digest_block
hTuglAPBzXYUhQiNjkHbZvjY7kQ=
//pragma protect end_digest_block
//pragma protect data_block
RATBq+1Sf/TC0qHI8EMp0D8+P0SANdM0lOcGXMwcIAqxxmWt0BT6A1n3ugBUHUdJ
+fAGodis1kvaBD8AwDhoQHP7DllnV7TwjKc/4/p/sho7UXyyTJDw1EakqZxN4ofb
MPA+sfBv9bVqGWpAYDjsNXVQkdyH1+KIHEaV3un9D0ZSZm4EQEJjvwqjLFZFNn/5
SdwEJh+dFNo0Ae1rj1ow1/LKtm+LfNdGQhiAXTLO+CxqgXH3TZUJedpQJ9oddrLU
dT8Lql5ugdJPNmMoaq8PgQCaGkHSJ/+saAWlWgbjD4mdr86Kv6MGAZL6pVOncyiK
8VITWOrehS29NB6Pgwte/hm59e+Sunqp4XsDtEgra2yp9jLiYo7irUkhvhb/vVW9
k/lZXcxpf7SCJW+7TLtYCrlo7Grh/Ymx4f+ZhtwDOK+W9gBs67QslKTxXfBnwwl1
KbVGiWg74V1YBukjH8XQrw==
//pragma protect end_data_block
//pragma protect digest_block
1RpmPo2cBPLIUzDqY4lfpHyXFRM=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yfgD/njpVMUsFrS/De3LV1U0FP/jD5dWl3h+8XDADh2dHdu6X+4Rv2J2LxoUUnkH
vaZKdhMMydOp86LJUiMyJgFIValwfqxyOo3RofRotNWfE17WBnRWak2OAxmQj9ht
t/jGVEGU/gDyn85RyjQW2o42CJpgBPYeoEVSE7PySQHlxLUi9LxVCQ==
//pragma protect end_key_block
//pragma protect digest_block
9y8RfP1WlD466gO0XKrYSbbyTLs=
//pragma protect end_digest_block
//pragma protect data_block
DH14VlHw3D/1Iumcn/i2VT2nLSgCrQdrCe+UbSKO+fX6h1IEDMbbq3SinBx/tE3u
/HXxIdXKSFR/LrR34nbM7wrR9aCmHOcAKS7u4lxJSWt/6oGk6Xnf8gntcX+3kIyX
iGla4j+aTaYNocd+ztUu+ov3ISO8qb2lAQWYdzlibmi9rR6Z66++XCj27xXMrZzN
x6o82fDMlnb6ZseLOVR+6hX3/JJiw1Zql34YZ4yM+0fvuN0sB9AO7pgP9iGwNVbt
5rKb4hyHevpDR4mi8yco6NdFPQ0QpOthOQvdUBFSe5SVJe1HXpcXTMxoetkq/5hh
bG0QV4T5BXVkzN6wJREQqlbVSaaDO3tAXAZkbC9SK1tlwLVwWs9pDrfiqbxzl9LD
iRJeDg0CifyYG3Pwpu3PCpfHJ8n4x0LXflvNIcQbYXvn2oP4gixbTMaGmUERKLb7
w5DjqXlT8TReGq4DlR+W8l5+59/wiOzvmOZx9mrE5QDxEsQvuQeGNwTZcSlpKH2v
6+051y4/h3DOtJnAsstNA8fDbw3thUKw0UDr8oe6KW4eKNMpMZmBlJUi/ID7It6v
fRnjg59AuAdj2Wn9x6jauX0yJgDXZ2OuFbNSQHp0PyAUajcitaxnBTOE5ii/eEOa
MZxGCgf+RPlsPj/6ea2NNVNyC/qYlZGmLynUzumodxqzLxheZWWYSBEBQFf1ysJH
O2v78oOq2dDIR0pIBteE1wTd7za/W3Gns6MedzJMPT6427MgmeVchZ6budMB6idK
gK4dW37CBF7NGtjCH6jpG1a81532Kv3cT/X45H8GQisTIAL24RNVs39qPQp3tT3I
cNP4LCXbMpbevVyNxSU6jtVUdG9Mh2DAjnvywVD389/VYyn9XeMwu0wUprY06kji
RjzNtlyaKtc95wZjQaFF/CigBBSXQQ0eUixgqCQfmyEEtnnTXizFx9TzjYIEAuK1
x0o4SxgRCCX5XtlJ911mSu+O25mWOMtPz3EU6xmWkQIq4OD6l1J+GKUssm7wvnfB
ZSXIcJkkLC4hFVXiCtborx/NAvXcSkrxSc/1QNgeI915IQm1dISzhxSX7QmmTs20
nRurIIbrjTAIWLDWhtktWxCpbYjAP+WNyeeEJHqsG+a8DERNzLDcBaeKp3A3yvmi
Iso74Bh7k3MRyNXpyPE1oLn0F+rzBZvlvWu+Z17H/qCVY3DhYSxdPwBv2k6s0gY5
yvWqd9w5UGXi0rpexHRkDgUCNG23RcYfAnFCNLwa2uIZUaGaksM9pEtE+KhxOCPO
O3XMQeYn7ZewTGyLWZQw/RsW3C6reaP3TYzlenuZNRNA0/U/Ch6v4DqfHzaYMkKl
KJVdS9CbS2CEXHguKbRSot8DS15IWsvQ0845YpqP6cnM1VQfTDYcpUVNfepa2aa/
ELu1Vcqiqji9OEA0e5tvhCYiCjUXQqusP+wlIRf3b1T+NhRAdDDwLx5Kkgv+eOzM
Lut+YxIv50JU6fBUrrkg3hWty1sCO8oCNcIjoiDhHzpsAvPULK/J3kHj3ptKyVRh
VGZ5uAPITNSdkoNF+npvOUVQbg0q5zhyVkdgOYE26/2CQimPslb5xhNU7xWXxQJh
GYQ83x3ndjYiZV4jzN4vjDxcGoWh+/lN6bt8VLq+9XN3KxvR5f/4s1Zauf4D9UFT
YVOJz6nSsMWHi8+9N0uGGgXzy6khUc9zWRIOpYFRBvPQ0KReZ7vdpSfN96mkvo9K
UdCCfCYU/Q2kHGX3Mh2FV4dFo2BtdWikpAElYZyb/63DhNBBAZQit78Tz/RjYimE
Ay3cFcWHRVCs/KH6xSGTLUK7Gp72YrkWoLFj/d0p3c6zNgUs5SHFQIsopbeQvkzg
W4GiC0KCGejptSDB/t8cONJdylAyQ6tt0YH+juKYcJnGLGMZxUGi3CKjUgC3yXbk
RRnPhuNe0KUxqmsNm64xWD4CVPKESVIf4AzZaKRzCnaDWtacfUZkUuoBzWefEFHy
+lcCRWk+4oeeiIsLvQQfzA7wWeeCX1p9U2H9jTq/WrBog4lE0t//qmdBqN0wgdTM
uR82SeUBuFbG9PoprSSs5uaKQPMjQLffJPErnkIEyBmea0q05GlAmhx59WsLMRnO
NyMsC8DnkdmI60uvGo2Xof/VSoTUWR1uCH0atX4a6tQvgCXs2hTDJmR+WK45Cn6L
b3/2qY8q8Jt2YbDC9BRqc9ko/YbC7bAcgXoHjRzUXV77vqGHzBbkigdWjenMYAb0
7bIkacLEIU/dqndNbYJhT/8tRT/IBCrij1zq4+/0rj3hphnYDGSM2l2/JYCofkGw
sIYPm94uP1QwXhYsxDhS1+1PIwujtl4s7BGF+s3WHWWXZw9OltNBoHgTD/i4Dk5a
x408QkACFOz9z3B6bGOsIG7CGiIMc2Jf5oNnGY2Ez9oBNaom4RVZu/76iXERJRso
8P5nW13edjPDmQRf1ejFroNxEPekRK2yjV+GeB2lw6Cl5Mp0YOFwiBYvzfsf2ZyK
REEA4jIw1lF137fHkj0jWotdc2p+EuVXT4bHse/CJZT4YRYguSkCQDasM5U2NMWC
mPnZYIRUAsoK3xJ7rD3fUVoPNSoBuySNPYMmR5PQnuz83mpzn3eWZelW6zfBZ+Q6
O3nmZW6eUDi4pSxSrSsenCmluKK0h8eEbC+M3rulan889r4kUcV7IAgOb/Jf8i2E
lT4sjZvDiUrTl4al2SPK6VDx7Wdkw7D1AHsuWwM1Ezil6fPGV3ad06akYU+pavJA
HDQhQGrCfbO8MFzZ/6gkaRH+KvexjnqQjGgRU1xqEw2snwG6SDjEPIWltQ9CIq9w
pw/CkNjl/peAZsOVeBBSByoR+Cx+bYqMmlbOE0iRAFJWiVrdrx/IAwW+3TlcPJ5G
J6rwokypnvTKqyLF1hqYYS+VWEWZwGtBe+Oj27u0ZcVXmVPQ9l8Ra9odw7RTX7QZ
gM6WHOyc3mZe13jQu3Ij1hEgqJkO7GBhf+5RSrRdNeNe1Pp22OQ/Ljvd1NLN+o4K
HXIViMFAOaRDNZCVZD+dXImG2W48WkST9gNM9HiZAWzK3aTVsxV+hnfc/x5gSQVu
nSMi121+AstfyUwJVWiEVDUdNDwNVeVy/oLW95/4/SVgVGbOlm1Zh5S4HKOvz9bq
f/munRY/lN3vBt9j15CdbUmi1NhGROY6Xl6u2VR0tUyp1y7i6eSJZmAYWc62aXXW
4hTAILSE5+WA1Mri6wDSyhMmvTiVISEXguJsNTNuzKH1gEy8ormqKtHzQRw8qsp/
5UkjOPxRGtX5FGnYhY0/ejNZCN8TEXcWhJummlfR7ttdxMHErUuJwhFHtczuwhwm
GB4N5Jm5op+FYTWunhg8gCNmWTHbxUhoG3h+SRv9ryOyt6JJvKXNsoE1rCPLLS9o
VhJzQ+1rlEGQBg/z4Y+VMlo8aE51luc3j58jC4OfxpxWHJAMTkKP+TG0CLE2EM+B
0YqBKTjNnMw4uY7xlbX2fOJBNSzvmp/8sdRKthChLkE7Muha4/DZt/TZwo7s+RNH
mG3izXhLb6BMXqB/onQ14kFO6zP3w1IcAqzK9A6qHWtc/UHi65Xr1w1tqp7UwPWn
N64EOUHtamdjmM8CALyUdIWYeVJ3xO33xXdwHmhpq1ySaqg1icg9M86B+b+HdjBh
HHkf9PTbRgnbiOmm9bIbPn3yjNX/4vJp8doP+OxT9AEgXjYKt6JafRWmlOmrA7D2
m82D3/ujrgQO1iOhPV3bKOPk5Lr7foTpcyaQxYYhiR9dnEzjHwLCzBY34i7EMBVo
3fQuSJ95ub2LB4sv5od6mTB3U+g91UQtYwkGRi0QQYczqCXSDEz4qJ8CAg5yiLL0
YtVvdZqpjAC+2y5qz1fPMUte6b8hDjScAll5+mZ8vb08wUeomFC7z8P8e+Cx1xc9
q2K5y9ajs+36i9wDBcHWu1x3TY517rpvR0P+AXsDs4GWNf93br3/biV0F2/RnNqn
KT/Zvh/n83ifHhXWJzJxdduQh6y+T/96To80DJqTsTgrmuuZwqXNSNpKbkwzmF6M
/6d7teznjV20xwldGBZdYKx4QAZAtQDWMeSAiivzYMQK02+qTKZL19n9VjiZ2fxy
GU6UWDhfDl+1O1hnvtWp0yNWopWmibvVyFUQRS+dbuzxfNFAZelZZejCJIeS6oAg
p3kXuoGl9nxqYQW9demGIzLZViMQ0pMHPk1vRAnozv3teDMG2zwOQcQGNhN6iVWx
Sy4iIlTkDfIh8whyf44Usx0ToRLwOqoFbxOh69PKe7MBpdeWbJrPgW8xda9tbZJ8
wRkTBtXORUNprA3CFLr5R88AaG2/z6tBOlC8Aj6KHo9FkJIWc9BzYt58zD6+/v11
qgeu4CeqfPyTu8UvkW+HiibI5E5L/33cpJlesGZ/o5r6JAfxoIx9e1v8yUqJHSBz
QdLiKnZzWYvCUhNaVWtV6xlyHJqOkys1ZiSp+wA/ljjTN8drsP+jTKQbkPA25W29
76kdPVlEue/gRMNSJEzRiIZftYD4vpE5iTbGP6TGxynhSBDnZi4YT1nCSlQdpUwa
srTQUd84pVBES0aChdriGXuUcrOoX/CQE+ZOQMIJ6nWKF2nBhHzwQtoxZnmjiVnQ
9VZxjSzWFwDozLfpg5JYILJQyS0z8RvDX0rmo2czAj1VLOi8YuXeT38vSiUQyqMx
Es2iorvd59x7Hy20d9BvsTXmcREP4nuLs4ZV48HF2hZD/6Zq1K7VI6Dcc1mDpFWf
sOt1QsfyH7jsUYUDqIfDpntg9CN3CJpTJ/WvJfmVDWFCxxCqzAWAYYOw8Su0W5ut
vwBzz7BSF0HDTCX+wpmibCBTRdmeWcw+chWZVqVt6ksSbkOIrFXo5HgTH5kNmYVL
wC6/BC+RQxV/Uo0zBFGfKXeYGmIMZ0CkbStfbQqaWjO2qVLrAGPBzqA6QzntXuWO
mwc4FzrMeUb3SINUZWmxD5jp+qi4uMVxW2musD3ElZjvvywah3hoqSrtbVdBVW5w
WtIeM7us52Qfr5tUqZc2iyt3Yg8ZbjKKPy4+3Z0L9XHqWi/CV3lleDBuxZ5x7ckK
bxmL5pCQ/v3xiNGVOB51D8u+PMKPuLXy3j8Jn8Vn8cddzmd9Bvunr4VKE+mgY+Dc
dYMpA1WDYxQZ6iVafxUsmp/8thrZJeroKTUHv+xnPmghBzEsQ/952A6BapYvh4od
bVTnFw9A+vqn8nM4G9KjOIRstUoitmXUmLVYEdOKjyw0OTu3BTRMDKU7/RuEGCpC
4DspOv8pNyroFkfPiAeKkp31nUgYa4jhtMwOh4aZ9egeAGrsQiMqIwBqIIIf/KDa
3p273otv5j1nWs7k0ZFFpzsVaXDJ4jtSubsi8juDwvIVhTA+kSfciJUr9C2yqYtl
wvneihKzZeQFwALbisRE34hRPrOrM28ZrigQyli4zHQCa+FrZ1Qynt486v27HSlY
rJJ3qdkneHaL7qtjkPGYZ35vZCWZz9OfJAy4Oc5MaM8I2Y8gb0AxFJgftyheCV+R
qRQDnn19QuKH1qw0oWYLLLe0z/0Rjsup53cZLf5z7qqnwD+uYnotRkgEOiLYWBGe
7hRotUBzMYj0krX1yfoHN9CC4rN4CrATBh8F0+6/Qj2QqMBsfjbRc5BOcyAZ3M11
zii34p6SBDfKuYeVMNmK4zVjhoOo27t9MsedLfMh+wnLJ5hoOsW0tTwGEwdW5Tf+
vLICFyvFWEOPBUAe18AwU7DsPEpxWPgNCrZURvxBKHrKVlx96l7lY5aI486WjaRR
g0pIS+RjeANVPQKx/Uqq/HOObSpHrKdfs8fNpkKV3BsT8OEmdfgMa6ZD1U9LbIXA
HVByYsGQTBPKCN/BcJNrtrv0vemy1K5pFv/FijWAM4o6SGD6cEtFub/GbIG6Srkc
OgnecRVXLF4nfnlG6G+Qh5SRH5GMUQQ+TRhOWlSuybXiDWmGcl8J4/pHEM4UktfD
vrrInqYsKaRjp4qw/+yfieVkmbLVNmMMrxjSOTwWXQthWF/QUon99n5tl1WEV7Ch
6q0DLD+JGb7pQGbhGJtLiBQRrcc9hAsk7GCDYDXGiihsiXnzAZY462ywGgxAnkT0
r/TiabtKtYiuk52exxtI20JtqMYTT4BNVYi3V94VCd7rq5nita2fb4guJUcvsr37
1CTYRGJHOeXvUYiRBFlZMMxjPrlV3NlwBAyYKAsQRuKJujvp9rweKyav1yYaYVl+
5l9nVuHsrTP1RFiv2tlVeYJzdL6THEB3absoFY2G6ChRNqKbc/v28h0vaj9V4NUM
rRLCpEhbPXRfEY3PmrcKRNmxk+K6c7Y94ErRLydYsbALFV722RpypUTv3ImG2L3G
AR1MisGejc+lkV5vKENNyWTMXw+ryQKyLJpo6YDepN/YWpNXCUevCnyNtBnSK7kE
72JRbNe/HOrn2AKCJ/uzugXkgTY8n+/wtUMq6q7gLZbW+l4dgmZ0ZBN1NmUqLynR
ZAGPNV9G7dB3DYcgAVcYErVsT9tlgV2UpfDdyVYPavdVCavmmrA9Q+AfqOlVyboV
mf2vcxUGnpOQNsMKu+7pdIbHSXr48GUWWR4P/w/Rw0FcMJUdm/1asoH8nbeOuoqX
2t1j8rMcYNU+cYxx4oJLc+rGd1l3nDKPbdNYTWm7TTlxCjB5jWlwh+NFFZdVc/6q
fsgp2ebZ4zESxI5kxwVUeB60CkDwowalhoTkz6aWqAKYBy5xGZ9v/8z1Dyc3bJHG
FuEuWYRQ4L/A3xSNMfuH3NWj4A6xE2IurSb9oLDOqLeMY1XIFK3ENQYNhBign1TD
5wxbXqb2HpnhXhLRN2FytmReya+qQLdKyD4/u2CwntLtMrYNY+hMu9jGpplaXif4
uyaO2RTcSk9fo8fpslk4kkzdA7D+XagQydqo8AKT9ucm3Zc4m5n2tSMBHg8ytogZ
OMmz0zemm6UnhtuKE8bNsgPmNMd39aRFe9N7yhkDjKb3qoZIyg+GA5H8DG0v5/Sw
U6dIWXQNi+qUf+29tB2RGF7fktctoyStlFKlcGcZgQmZzjamVwvShy1VodAUPog/
okQRZDfayqq2Xaf2XGUuJX7ix0bVIczHtap5QGhpfOW3l08L6P+lVeVsWuFNKUXx
wsqmZ9KueinW4B7PaYGZjmmUmzStppEkc0Iu+NfXKCjqlP3q+rKfcsgj8nuyJ59A
vUhzPTTflZwyAQT0/570cxoBD7FMWJn9Pveg7so7GJCTF4R/NeERhfZLBby0sc13
fkkuCW5c1cDvau2j5v8Hq727SOwT5Mhnlzl7owzGBSNMYz5bu1LIfMcJ1JJhfrL4
HcofR3LvP/dV1Bg4yeXc8fqH2GT4XFgPrA9+hh2AYjDh/rc6rrXr2ldegd1Q+vvN
lMuoo20qjJrrdkdab0hFXCu4YeQJ/RbQo9m0tH3Cw0n6AK1yaJTIfiEnU8R4d3zS
4hDSN8skjAPeDeMC9MNVTzU7jlyP6p0nBH9atBfJTP/2wo9Am/Ea07vahUdgC54z
sBao0aMeYa4wpmKkGtETTbvvb1eGoVS8T7WjJHrf6zQWvBO/DEtUTb72tPBGOC5y
xd4pJYyD6UI1SA8442gVgZaUsrGJE15utRUoLLosmb0zQ+UzfJj79WOoIn3k1iG8
N2m8Osiqo5THZ9Tz1Igt6Gd4AXWFYDb7csJfqyv8yrzGWPlpYOCUPoXCRQPCqHUr
Y4pyMceDyE2GXn1Yk9qQKpT5rJoYTbXSjUP4dgwexY2E9KU/r0gpUSULrlSFllqq
mscTUJjff0kjfvciCoUSy7OuJ8RQ7PyNQsStZ1kG8z8cbwxTiWO9nfnCN8YzYmp0
GGHbyiJZ0Ww+jVa8LoEu2a3+Ja+Gf4/mwklV2Y85+KPYTrDuUycu6e6FlbBHFc7T
LOgjgd7I6YeXmBInlF9YvSTs6+pfG2W7OQfwTyzEWU9wQyTJlrpa0hvdlriHTnGL
UoaUvRIZIB2+1G+sB0lAME6nrf9i2sZOj9KnhQeF1UFuHQw9nf95Ju0LmRrq7S2P
ZhGT0BHVmBLzNnv+3hopO4/hfzUCVzI9fztUBPNO2hN+sM9GiP5qYjJNoO77AdCU
AFCIGRLrMJpoqDd52oRR2Nk+EbfrU/jyHeiK0WYEBHIwaUm/nUI7u6MZ3HdqoNfy
TIwRw2vtGZOn2I13YLUKNmxYeDKgvS/s8MMMV3nC2H+WMU/a3j7HwJ58ZBtSKjuy
ICwQHq9l91+nI2SVqzMxkWhgs9zf7VXpuEfry4nPR7WdwaqnMtKliCxLRN8tunUX
+sdck71hl7VriPHwqkpzT6PLuABhnBO7Xixe4XjGKHdIUT/eakRAVlgnVUIDUMJf
0qD+AifukK9JJd3Nxb6Unc1O6bzjlLVipSKbrXbdRZhXIQ2YBu2JjSDq5cLCvlg3
TorCzro666ZroQPJ8pEGga3kZMziBkWHzFCEHq07behiZorgRpsHriZRoYvOOuGj
vXQC2H5oDJaSgH+AA83UmL/LCe6wC4yzNlvNMTy7a2C6bGTmyJrvLLvOCeEh0DOP
67byhC5FvNGaXYdi/asm2ttPqsROOsuHNoVwehePoctE3Jfx1T8ayuPS6PbfGttE
vvvrg9R9kCYbqcBvgKxtMKCupIcI1OsTzIvbR2HkQR1sVgjw6HDCUV62PzA/ZrgQ
R87rFXk911SjIN87j099t3zo2kkelP6tVIpMuq5aMxZyqs5jqyTJK7uXKouiVCcF
Jwgo593crQRELU60Mv+uP3f8aa0HeM8htw0zjOKg5rhmB4wH3x+1OI4S45M90khK
PNMd7JYBkRiAfX4LAtadpxyvoeyoHYbmgDgyd6TC07u2mVHpNZjpU0XiE5Bray43
z8I3z56QReL10MA4U8fdM3nVw0gM2pmMBMABiFrlvZf22Op8/zpBJpUSxRUSqtir
oRrZMhBZB9HdfCYCrbx62YP9iUOzNohGVI3NbS8lNH/yD4RScWvy66POdooMT7Uw
lKaFjoDhm6mZ3FGUGq8zVDqdVNeJ0QHEyiud1Eb/amcveJvOZ4WSxJfcdFLVscdv
fSgY8YJ9T+ds7fOWN9Il4dUl/pHZJQcP/stzTR/LJzQQ3SgzYngFvk/cHySbeZ9k
tjBqyuNsb/XccCDVQkUZYPhgKMK4TE6zAU85MBAXvsJaYywe5wSNy6zYgWvd47CQ
dzwuR+N29e0NYCqZIk+BsNSC3RMRIvntf5HgBnKQxfNpjpyffa8g61lnByNSVIoJ
szmcINzTxE/WD5lBb4BDwAvUMUlekoKUo98p+MI/hJKjMwwtSeJpbjjXOZG8/gTS
vtDF9eSs5vN7S686hBmOa6KF2Q48G5/RuijwAvIjhL53akG7kxWX+MQZVHXz+3/s
FsfanJtLpX1sQeY0VJqbzgblFu4SwwiVOXiD+c/LsVS0CCDUO9kVOoiGr8TtgNgM
kZPMGi85vOa+ff9oKzLu6vulcBs9sI+FiVyy9mzJ3liyE6Srp9LmNrtyBFhifhAr
QrqipwraJj/6geY1C2eXTw+1BoOfvjRVGFGNoe1tszGT3RIJLmYwnPUahXNCxrt+
NKmvs0z9kVKFDy1aHURkK3scqAaRt1np+4cmjpNyumBILN8ZlbRVdwRbIdwzjcuA
Fd2xJjJAVlyWfjDSoYaD3k7skWeDWMEQNLs+qUvHtOnxFUotXVJ7fUvDTAKM22N3
5ILY7K6XD/HtHHHIlk3CRJRhgX6msDU0lHbqgvYcxu9B6i8HpVHeF1PWYv6G7mxq
X/XZEpR3ZQYbA5RsNKoufYN0eKuclDJ2r2O2rfmSWAd/xs6WF/YCynzXc6WNOlQQ
sPzxQrlgeYHNqiDVRJhkSIXHjXTqM5xtzP+5xx/z4VYXwq3NCmfR1CBXaH1lMp0h
JsoS6gwP0MrIJ5w8uUs5EplGDxe/+QzPWE0j3apd9K9Tr7E5Ly8ngZBPmrZMj4mT
r4V0u0lhe5zmgg+BhxQOBPkE1pDWhtI/GumM0SB93ho/mkZW7J46dsp8tXZ4FSQl
0Ew8wINDWyE39wIJb45ycW17Qwd2nwSQCEnwtCtWIKurihrbRf+TwprlR/rXh2Uw
bxIiOsdQiqJ72cEqNzsKvOFqviy8mVtMjKcN9JOEmMu5XusgoyhqskReWCzOge2K
wCEBkuPTac+KWfsuhFF2pn7ou64eeexgnOnPVBO3aEym2fFDg1LQ+NyHQXBUEOz/
GigL/GciVP+puskt43I9Q9IAH43LK1Y+/ypeJevNYvEElj7p3uBv/3a2iimoyud6
5LVh3eigsCc+4VyLye+SB4IS09PkpqCQm3Dqn9KhZH92w+ZpxhFNMBEStWypoeuq
BpK0ZxhNuXIL8pF5y8JVS+blixGhxR3Fw846Wsn9AkAw6IZbPtxYIoU52e+q4FWI
zEyAdhZHVkycaxlzGs0r6MoJ4naU8LC5yk6oBoSzSgOIOUwI5gn2Wg5BlcyUUKwm
szZEAyAKhYoONB4cxfSwAUEx99zrTXp0aQydJbBmGu5DxyrQVNgq6wNK84wtMpHQ
PRY0eKYmFzhoXtcFqZOhAAJER7wXV6eBIcJ5eFdWtpo0kkUzDf3tWqdjd6UGWaNG
s7g3UKmlwBQEyxjjB0ymtY8nenLkGLALSkZNThVFxa/hVxvig2Z7qhRjpnPyfuXn
TsLOHR3XSIwQ8MRverNmaZX42zxcG3deBgov+MU12AJx7OF8VIEEXRbw9/R9PJvo
1LKOIj1RRAhAtf1LudNN+5teRZojUMz7aOlAW/m/q3D4Pa08tRv9hy370YfDjT0B
TdapiqzGbqQNqGR5T+TAvgMAjwGhxg2YLi6ZspbU4YeF06LRJUClQ8PxGm9bOilk
L3ggR6XF1dpvBWKz+2g8jGf7aDIKdqSMVOI8oq296AfnuUOYPq7eQLSoNNksD6+q
KMpXGEmQQtKIxVLjv5B+ws1trPS56W0jq/fVEU+FI1eQZHFv9/vWhkOPp0pkL83f
c2DLKzeKUay517SLr/q08bWU6ZDK8hE1dQ8X1vQMhSTXpEG22V9fKTGz/tW9Obyk
nn1GUvXa6K8JP7RKcla2TA58m4l7vgV8e5pM3+XcAunnTnH1IpiR7WjjBKT+fgrq
5TGDfODgDGmnaFASVLFzxnFlhCF0Jck7xN9ntdtbN4Hz9x1Sbkjs1Js0baYfhA94
SSPlnCNQA/0dAEu/xRf/bOriaRH6XEy/dcT+wjFRFWz4GaKsViGoFcoRbiYwRBAP
CXziEDbPC+MNjuMES0fjM6poI/gs12ih8PmiWghD6lNQfLC0UPGlydfgveF+A9y0
8YlE4HBmqdoF/RoWAdI+DLDkNwZCd/AYMJtT5qRlJYgr0pRe8eiymZMv5oED2oAo
pP7tDGU9uNI3pPXiGuKZoaG4aKmVW3jmECfgJ+ER1kRjaRRVtWXTfbsvjNh16JhJ
EkuM5FPCUCgGrclCLQGSIrrr1pGIToAObzRtQqM187Eue0IZFRkRo3FoZTNxyGxT
CH6UlhsYyzGFL98mdiL3RTNOKkbwXLbYa4pGjwZat2iq1xz4dS/Gq81wVXhFGKhv
C9iC6zsKbQerheJNjPDyBZ/5ac2kgIoCqhI8SH3eL4iGIjEyzlLiQOeXQkgy7L0k
qhJCctMYplEYkgV0i97R+zsnlpmhMbVYT8D9x6nadC4kDBRWN2Uk5sPP/OkmxTf6
8HueeeSL4lqrTdQ3MyLCah6NljVMjZ2ibro63WcZW7dRq+rTbQzTexiId2Ilo3FA
cXnh2xZVxoK2BrkWf/UsAdUDfDFYiJUQAf+HNo2bT2E/6C84LSwbJqcIq+1Zkdxv
ju5ZX8LOUWnBwhWv+ye/IE4M8bE9N6pWGs+0L/sSmLyRfEP3qdrhGK9YEeTtAVds
Fe8HwpV0TZjrJ2BnD5Jv6tBz0jk3puyNUKZq3zbLcq6lxkLCpdEvHvu52uVwYofI
gA20KJyWngRMLFdbGa4+eKCXAZ08Aze9bZyGBlitnbVbrCQaa4Qx1CVTX0ufSdHW
sm2hyeSY56NSigHl64InNNP/AWMi3zMmXMuB6h6VVdqVgpad7740x7jB2Yau3eB7
QjY0ZegbJ7casgXvyeVr38g3eM+TXYLLbDhIE5DcEJOcdKh1LQPAB42kLM6bdgAh
mDMTqBkm+D1nnKZQiYEalngznw0jYCHfM5gmiOLC2AkVNTgrVjHNsj9+jxR0qSN/
GaZ7R0MjV+K0NboApLBaU6Es74sdceC0XEpHBACr++kRYdYdoBtkjR6bkAHbh+Lg
2XCmQSQTohgme+Y7lZB3h31tcggjX2VaGIVnP3qLEll2S52EEsoRFlPvh0qCPh2I
HnICS8tAOALI3cQ7louGqJEOvdoFBmzaH1MJOjx2of+RKCJRkLAyGMIjwB00IsXh
KaVh0waKGhGe3XF0gVB0G4SMCXabTXGGf2hK1T9J2/+z/7Bs3weo/hR/LF/iM2Ws
hcukTo7Tld9mHredJYw47Foon+5X49Gqv/Xebpz2pE5IUqNMa+aTA7F/CG7v3Jzj
KN3MOdcGl1hGpddIaGLLNKbza5xvYZ4T6EojsqImeeNSr6LJCRWWe5ObYa5lOkDk
8l/Oq+9BPrGMteOOonyuNMP0LDD6HHQkHWMSsl+uU6NVwIXJpujCUvk9WdewiG5v
3VDyYvuB98KMT2eF8070KPdMp2v0dms2A5ucSF0BKSFR8j2jDmj0n8YP+Pb6F98G
vgpsfai19yXaMqWGp/IgTnxU2JBvh3Qf7w8VaX5eQifHlp4qXwvhK39GwpfSpETT
4As8/8VFHTF/IjKah8QtB+jMY/noe0K4YoCLeQhavQ6z2I+xEKNxZFoo3SgV2NtC
dPxjRe4JTWEYat0brj3p+cTc0kqS9502mOXkjOhFqjg4EYDxoaOlIeLpB4DCYRyA
Ef/5oq8I7aaVlk+snbSx3AREI1+5F0WbDcXMOpFJ/C0yLdtNbNz3vsF4fKE5gF0c
Kb/wpw0bPJDboxwPQ7jIq/UteMkW0WrgGQ+PCzXVjigH9ELznYf9Y1fLqAISdEEP
x8t5/kYy7nc6t/CMpEbriwwezZ4oZ4SrSbANJJhOAvK5IdnzDZW2ExfQlSFRr6/j
T8xKpj1ZwdYGApftQjSuGrqiJloieynP9GTmgKbfY4EUj1AOMEe7HZMU2TvueKPj
ead5OPN1Za5zNG0ygJJ6oTFb9FfJrCA+GAZZQ32gTJjEBRkhe3ouyTaomR7zM7Uk
wr2FOeuwRdnv5Oti0bJMC+JZuVKp9JNRLDPuSfx2mJaRkNDf7+FlpohZUBH++A2R
8MzNTW3lSu5auuXaRjAmtOMYa/kzFpwXkmkHeZOcGE1aVFUfhsJwxAFXoOYQGWPS
V/bULSmVBZQDIlyWh5Kax0MroEBylGAIt+hteqZ+wdVyTbe+MEi0id8gOXYErlsG
D1hoddlXaqPyzDMvKpjHSURdGS6wYSEsFTrswVDTTCtyGiehocLwSlerznUjeVAV
GfMrdGwIPal3LkIV5HZeWC5OvgsEiKT9fC4OEeaXfKPk/BpdrsUNYWdVMQqZUCrZ
SKrbIwBX9ouLZuTkdbeivV0D3QUMkDYbZiAc4/YqvhbOASMK00nDDM6WM09tnds+
ko7Vgu2oERjIoEeREWjXBBKRgsGbArhbYTqCZPBmywxPTYf6wN0ncamG8g/F8pKU
8h3hKj5XC9+hyXQxEis68jz6KKZtJFBILJdeeIRbhDRpQlUkCox+IbMalRvz8I4p
XNeEErGsIENc8kGjKMorMniGORhquwqtWArwVR+r2Zzj2hWkPzawMl9oIcye/3jF
awSFaRwDxkpiLrCj5QfjtCvVp3rvzU0tlWiGL7WG1JYAZPoS2Wk9VkfBkNUl9bot
fG14RUiZMqnorof+on8a8PkU13SwMp5StyvAJVB3yZ6ymeW2QcJvueM3epf9d548
wr4JHNaRWyDPnSBtPOyvJ+cOyCUHu+BQomFov7kI/UYAjUOv/5MggIPDyNoHfyXS
/Ab8fc8gIYaeV+tsGRIY79WP6pQFlZ5mMWxDYUuP+k2eF2zrUmnulqaR3JW405NP
p3KDs1huct+1XwN6zLxuzrla+pwg60uoQcvjBDbv60lbEUQQAQxK/UWF4YvCMB5g
FMjNh/BycBr7bX6ZpP5URhhXlTHSPyNlm68F9bkvOhjkkNd4anj3vBVOO5dDnWJ7
j+NFGzsfNI+i01w4YOgL515JeSGtQ7S45V+FNn9NH4Qp/VxbGdL5SPiW58eWBsso
5dvqXcqI078K4MVLiRRkuZgo0nlkw9jCqt4FzOXrZODiFl6ljRgYjCHkydktbZRe
V6v7gv3F7nDVaoY8wKC+F9/tjLiTsGO8y2zXZo3hN1MYBdvblBo/KwgEPHeN2bf/
wF6KyHEaBDrwBsB1I7dvfzQ+llJvhg7k0EVavolxqHJeR8mgyjGTX9wFVbO4x/Yt
qi22198IpZP5HEISxS8sOBBaW32HEuQAYbDY8w8Gn/liO0w2pLMgaC55gz7faEO3
Yxb8sylWcvUD8akRnQq/buRO2gULc2umH2gCksFb11yCHlL6m7i5GyZBfkpBu1eS
lXK/9OyYUf+rjcHc1gt9YqoKruq5eqtiNgnGRMt1bOnYRozG5Ijs0X9aHH40aews
DWDHFIAoh8qPCdnWo4ZAOKNnBlDhAY38pO/INntG8nTs18haA2pjzh0eqdqNAGoT
CeolKUfnHiagKaYDAXSPzoYnaulZo3TLOMtkBqYQQ8zzATiarlWIZWyvvqUKG5uz
m1nVIPdKiQDAzpB4ZlWbyzQyFTke5hKhfUx7zwbRezeT566H9dPyr54UInfDeKlg
dMERPrtgzgXVCyENytySSAWSgOvulvZNKPCtkmtCOaiYQySR0p6q1r/VFL1K3ske
ZntW3WnYM9b6Xp0z1XGTAomiLNVv9aEjXb7w/TTL+GcInUknh3mIlkXiF3l8xGUY
arOj/CmE866wLSs63geRMoRLryO8sGrsbTayzArnW+NCmm/wmxakMu70Gj8QPhFX
XAJhHEFCn4atdG76fU/E5mVVQANr+7r2Dm8k7PYxDKwQ8wfssvXUUdmdoQlQNNqf
ut/bRd0RYXBxO9p1xYtcZVYuvGxruZRxtWP083QmS2Yylfw891kWh44NmFM329Zq
8RoAvcECb/Y23/hps0kNBIuBP8TwsUuKj7XwXq5zjqZJWNhCrP3/YYZ/Lcpqsy+i
3/vJrGqo0eeJvghEMHFU749iavMyUVnEI96FBpKM4nTex3WzeNf+AYv3v1GR7W2t
e9Tfw9ZLQc/7sfu69vopqvK78H5CmPvxRaeoNY+p0ZheJSeLaIEBtCeICV34c8E/
Ix4Ykd17eJY2iz/6HqYmwPpYpXYFcA+lEoH1anyqNDFnLrNBTH1NHE7v+aeplnt0
1zKLIJGHoDBixDY4W6AwI6cnR0IXejnujfk2WBLn7NHr3a4UO5HOzqSs4oNXz6Ol
ijeUS4fjORpW3xQX5CIPZ8kjx0ddUktj0tZEDbptlLLXnCdvk1igGyvSt1pY0RGC
+/3wwU3yPG06lj+ODyU10gTUJfUDT62ayhWeVP9z60XLLCzcQwz4F4VmkQtxvp0V
IRspcV0s2uo6QK9Y2FChW3mcfqmg3BSFdgKkoE1AGdOJleq+V5CnHw1gc1W0d0iX
5qKlBU3KgjVX2ItKCnL6uRAyuiTThl1u7R1lwSH1UgRNg07ZLvb2TcVD5VdClC4y
zcLBF2c1lxa4632jSO+DDvj9GQqYaVBNRnjOcHm48iITyudcXzwzWFm5oT2x4sLs
y8hAmn9K85uW7VDi45/c3vJaBfakp8X4KnBSEL0dahEnYVJvxWrKtUEBbHzV1zO0
RVget9GZyHfEWiRI3CVaGnLmUA7ZDBmAQqKbE2ubcuEDyEpmOAkNNNtdudKbKxvf
LBPUWKN0lOc0RnkDf0ez+xHQUhIBj1pxfVlzungak83Q6zftD7awxYvb8vcKoUPg
51TMSK72x1WUdin13Ve+Jgz4a3hrIryQEf0CbtiM6yejHLk551LBgm0SVIzqt3KB
yQ7GRkTkJTrBLaLx8JkEwH6BniLR1GLWR2PLP1XqleU6lXm0pDcONjrgfrSBTcDg
9ydgtzAto13oLvU2PdTc1fkVExQTXmbO4tm3H+xd/GAWtaTAEHWCA749hUPRS4fw
ICATVV/F3uTZ1ZMB6F8LIHtsjfXnREZ30vpoh54oWud7DFlMT1L5CIIxHtGImQDO
XG0r56m6iE55i3mmCYGgiA8SFWY1PmX/jKGZyk4/uktnPG6AC1Zl0SGis9ZECG8j
HkXDdfOiP05sOtZVKc1pgQ2I4f1dyDiSRHQ00ZbuNt2R0xZ4eYcxC0Ohv9Yhyy7f
MtQcedC/PLa/w0SGB7T7Bl2y4jmTZk2/SibLxcbl03Oempu/ZYbzwB6NgRfmIE42
sbbq83Y4b75DpUTvePBuYBabFyQtbN3aqXHo3hFxTjAGmo7dUMhhs64Rb46uWhAh
jhJSBBhQYHM0ITSGxd/KIieMrrnB/85jgXzwT+zo/OuTMM3c+S/g9N+kSvlg67MT
g3hBSf6NMWTYsteXu+3jeoGgA1mBfZq8HuuBcB4E/2Q5A/I33SdHU/Tq42Z3EDpb
ZShWSYFVSLsLfH9OUsoZLpb0i4e0PrvG4F5yApycHqOFBzKdZ7xv+Ahrkru/7TXk
i055jlVRQuWO9gTplahy6PhncWszsOivIGKN2vSsLbAcPLMXHjELiptmVG+mB7aZ
sjk8BqxiY4JFwSQCeMAzrm+6jcIHvkTy3d3zw1BwVe4EM6ZPMmzbuo8uoG5in/mH
w0N6Ml+xUct1zQAQig18HWmwYsJWd1uAlBZQ6+hioyxIp+nsjOwwUSzv11sZrSf3
7UYkHKUPAMrmbSx8Wiwa/J2cQSYvORuUH1vJ9A0rjL52jrSA0VhiA75vzgTNffM3
wLn4U1QogXL7pOtfTDKEOs47qM9KNdfpWfEDNi2U3yXoVSpN9hVy8o0WEc1toopC
xfyYrspqnev2BKFe+t05fJ3Cs2+VvdTbK5K/G7X1jAsNo52MMUliFtOiqZ6dmTJm
q5Wpi6BW5VVgNr1SN1TqxLBy32kZU9TUDCxXj5YwaFG9wyrJlI44YWnyHlhhkodI
x9L6GUiZgpcv2CMVU+el6yt19Xo5GuwYDwX5Hmk5KmzBnVOCwSn8ZDv2x/glWy9c
BJQaom8AMpntos54rE1m3oR4C9A8Fr4Jq78skIVb25zywIhlpp1vhQH40szlVpSx
87qGhF2mbyxrx6ifJKR7scmL1oDU77kBciHpUZj1m7quCByfa5gUd0HC90/uXlKM
0UCkO4dtYi4x7qLPNBgdyWrqg0sKRZTReWsBQUu3TPlN/+O+2IY1CncfHxYb351f
E5B1HKR1M9HuuXvEsxhe7NVZksh54O1ONF0apeq73///fTMpK2kdclihIhF0o0Rn
7q53R1k3bu6EHGH/B55eEWJI+5ReZTs7Sc+kFMOHBkBPXa5hHxeKZpgyjfxQrxkB
tlydZNP34TNFvHSBFnKnuWx/ie9OeXmpEPyBhb3DThjgA+0yjeF7QwXr1lvSSNx0
ZutPSksWnt+GRGxR98rqC89LrfDGCg+fpOvHFguNzPeA+a8+Cx6fRCTheF/F+dRw
nN3Euci4V0We3hmV4xK5Im0BGRX90oggYPjrKkVymSmXFZncJ/ZCpiQd/D20ZS8u
Z6dy4vHIbKdOj9TRiQd+XMr5FNY5tMPy7v5NK/eSjgBxIp4R0gUmq/0TjfBaMHxB
VBxWyzlLBf6F54lUXKM9Me0GMGYkkP7KPERbIkRZfxTJcpvsPJSJM5b1ZtTTOK1P
tBSwbRN1MqP8Hcr/xNczKGCvVs1MUfTtq4t2f7mEvpWqOLEfEvrz7eSYxtMSlGYJ
VIQICvC1vJYfq3ot2w7vo6tswlS5ULGUrJ6uAYSnFl55ljIuIUTnZynCB4QyrvO6
bg3t9sl+rkJaum2fTPx04bheVd73QPgXRJf8QN4cNjoe5ByXVJ18T2HK0lU57vHG
I/JyYMJJqUmS8CNwOmiRjMWO4fgP4+ZE7MyI4UeywC3eUYm19S2nMIeXaA+As0Jm
CwyT4ntcooCZNv9FviO36gQkeOkTsx5nj+BWg3LnQc16PXWpVUkFFsaxEVSgoaFX
DlGyylGT6irXjFgAkk3GZ/CidSVhecoSClGvRayn/ZpUoJ2mh4UubLTYbpLhuOdg
E5FEooQSbckMI5weneef/gBVQg5deRPxfby0t8jiLySMuBk34ORvah7fnB1jO9pG
sDSOdjG5TDFzmjBrAldLrhOcivCOtF8PhrmlCMZLDLHT8Qod/GZi7VpK3X35g+P5
BhSL0GNgNCeNOE7ozQLTmjHbQ9/AukUX0OJIg2ho623YN7t7FV2u2sWtQGJxAe7e
n8NW/LKnQcPY573pgNBl51cwcGisKpvbDlYbwskkHUytjbsRlHm2Sg7E/cWBXp3o
xqnemh6W5cXpiw+Aslze2Zaau+Nd4tT+OCXXRCKU25WWqR55V32g5CKP8ApcWgYT
un6kWL9R4GPi6JgNk/a3G9Yi/OM9YKrxBFuzFNtTq6JR5h2AJCsIumis4jATTDXS
O39r7qYsXjlYVKRDnE9ofSxbv53e9ysZX9/4frDofbgRqNvvKy5HaYtfo3ykDHup
i0PwAm5fm4yizoRgG4rvwLlrKkVU/7PBttnByHxLHGRVpiAeRj0Ppee2owhD1y8j
rwEM81rFnRr3MEOq5GZDe5COdjLfvwTp/uKwtvHPPtQPcb/nLiRCXQCkbOJts/6j
PuhD5UyDO+JgF5PMn8IgvZ1Bd+namIB4hun5sJaNywjrCuYAo2haIulA+/cmCUxx
4S6ejTp5C8KDEZL88owdhUXY5XKKJxtcgzf0fjdGjqX710FBdJ0czZujX+mzxDeP
ryoFcSo7TvJ0JVWGUBB1Ea9nxlYDczSPTHZrNFr2p1aOjZhbw4EQuMT6FNMewa8C
FiZ2E6RkurxToie4ZPho9AoF7IZC19c0Ush3Ghome8mdLnfRjshyb2vSuFKf3JVt
kE/1KfYFXtXsOOhRxqddZIl9bMFtp7zO9nOeWHSCRXXhN2WSzRAB/fZxsTQQppU8
SeA2mlfe5bRe5gAPnQ7roysYbkjwFpZLBlBx19HsVWXbaKopPVCMKGO7qxgvgHd3
0sfq6U/zkFtRbUwB3ySyTqCXKnqZY2/IWtGUrLwx1tEF3NdIG4czbouK8mUvYTU4
Cl6P6Zv+Xg+TRwPkKCf/UWjdhLPy8HllOxUPKoddC5wXgS4S23W70WM5FDMe5OK4
JYIKZaUGckrQAOYpr2NtWfmrHhHXUJ9mujCyDccJrIOLJ5a9kGDKq9np7FaEGan7
HgTWsAbn4/dEO5UQ188gIn070AeDcmnxhleWJUc3xKEfXmjQA4JSEBFkCaVd4Avc
4MBApF4zb7eCdpN90oerAa7gSHlLf3/JKtNLE81T9pVTpBmdInrseDt0PQnJRgqt
Y/Ul/LMQGGNaF9j1Dfj8SS/dIsbwnaAeWApr0nkaAIa2VTD+69p40mrT8u4Ygew8
g+9kxFiJvb8/mM7aDSOR2G9p7DJhyqZsFQvS4Qq2MztxVs+TtuXEXpSyHxP26eYv
7U6p1gxoxzWFN3UqZV35R+pzMOWs0tfTXFr7esARe/euxPxvqeQbkwfPQ0M0Q2lj
1slVPpuzLgxHTokS6CHGw9Iy6jB1wXoUnV0jbWb8h7dXnugYnxO87lIyRmisNJJC
N05gE4jauou3hfCwnsM1EGsBPsQtQf+AmWs736shBc4pEWaseCa+Z4Faui5s9CSL
hKcxl5jJfqBJuzyAGaRWjq49CYCEP1vp+QmGlga+XOPaLOFw1m9f5Eh44/qGKl1P
A3m7bGfnecaA0ViEYk/Bo1fFsX0xqIkoFOw3pawqiI8O34jFxCPGeTHSQfuSean7
G48Yf+IX3jzL/cXr8l+vtA+Jv3w7jjSJH0pF32I7DPAhPl4a2BKLToiHEpBp5GGv
CB+JfaIG7Lu3E1kk5T5oIzr/p5+VK+EILO9YYu8ScNEF2uhXy7h1pj4hVvlXy6ZA
1UBfENvs+JyZTGeIwNZTCK8yOCKOSvhqrxZfa9Veet+eEKSJkAMEE2KCGT9jrxub
l0TkwhbzzzigzAjG7WH+9j1oD9EeAGuGwW8aZhpvm0XPggwg+g8AhkWoClXVuQDW
a2prD0T+OVh38Co56t8q3tAObEnORCl9CrQsCjIhXEmvv/MbF81BpZlxYUIssM4M
tT7KYM7JwTbn7AGJgAJO6GX0gbnVF6N7waEtlJF/wy4vE0gMNAduYL596obWdQkE
ulZDvy1EQVhRIIlic9x6VGWEn8/9TiDXeupnKYln6T8Y4hejl/7EFPxStXHe6rCK
0MeX8uQGe5tBvguKZ389GQHxTKx9qi3dE+NXqmMhI7YVHwZe6uejqZgHWDe7AGpk
l5nDN634nqixxd73mLsAMJ/pWZPDwYq2kntHMxr2jlWXkTkidrjIUnHoGnDbzR8Q
UQVpCw8TZD2jWUwDHYMdeu6kQ5YI+lJqo04FR2oPo/M1B6XuIdw+OXQb1WiaTrAy
ariPUcpwmX6Vg0g40Zmr8yKXEWeAp4LhUMCmHImPz7rSds6J8oQoEpcuTanvHbMX
Ods0eqlIu9UIDKEdZvVUh0sqjUr+p3Z5REhTmIHyMRwWOrgMHYm/TDGp5kNM7i2L
i7EqY/zn2aJAXVO3RGc82AzXxdgkfbUd2VxbV2aPVvbtGXmy9aiKTGMgc2H+ZKK0
NcTQilDBfvLdE/IyRP5Nv4bbuaQRF8CA9iLrhJXjJ+YLsnjUAOr9GbeXi9D+8kiT
pmZsacINRS80TBinE23XAefTwmdYy/2GCEn1AR0TLj9F+bnmBKV1/gQ8ObZFW6We
vbZ4V5zlc7kSOFZiEd1P4eBddYt1BuIGQI0NBSRkgbKf50c8hcHdmX2aYuCmL1Ur
3UDUOKC6ZWyyNHGATfZvctNFOa05G3alJ//11i4Rp1Zfww8REl27G2yGzIBDeDdE
6E4bN2kGdZR38n1SPYWc/t8nLFP+/qXTCPdJ9KUOW3vNk0Sx9ZASoYhCDJPjNdBC
21Mm9V88Gc8lBUGf8dzgU4k1OMsgdQTNHT56wAc7EtGCZOilkLsYdYOONWE1H7TA
csFIA3147Ldtj5c2MVeye5lraWVObeiHXIbGLlXB6DLdWha0go2HEb4SMe7yRohm
ebrI7pExrykn3P8EjO/l5lk6CGE6O3DlFTpbytiSlqPrlKntVtRnJRhynM9hinzQ
cEaHaVQNrYN5P83n578ptSL/PDXWFeZbkzk0S1Sba2FAhWFUf37/Gbpab/PfnXrL
U39CfxQ5iW50KxB8mSATQ0yEoDgp6tjJDcHVRSL7ESPuz46UC+FZ4dETWN7mym7W
WSD4v2NkNDErbmC8xDidciGqJjixgw47xCZKdoB2Ht8AnM5q/1whWMI9orAPc9V1
w4XOp/0fYodO+7tHFNwfO476A2O/rgzK5Sk8pASXm8ub2/b7ttRQ2pKwMUC6bWCM
ES/K9CQ3Y8fYBMyjP7Pscq/o0UP8hiN6wgehU+Og49Gf+rta9dBPGZUf2HBX6la3
8i2JmEu77rS/AojLQdqnTxB9yD46XJkdCDKRamST3pBndgDpcTOS4f2HygR68BXY
CLJv66e0cqlORlEiDxTBmoyRQFnllsT/jXaVxWBy5grz6zf1wrMveztXSeP6/JZc
1fJJJ1EGQ/FYeJIKS6NmgSf6Yc4/puNNHjZ23tlc9g4eH6LfgACEphRTcAe9rC6o
G6C2j0KiNHhb6CnfEtR4ik94DZzBrDyyn46vnZWA6QbJwnmcdpdjr6XMTSF8NFO0
LHeV04X1P6nX6HrF4CgZ/ZsPaLqOVVFjf8VTuLsRG3OAt4xR7v7ben3rs3VhB9Tf
OrEGn6M0fZQyOkqtoaMeRUvH7M9ez1R4oBXKEDc2UX8Oo1DwaZZeR6MXO1sJAry3
+HUr+PVAG+DYUbO85+DyTo1ZAvv2RH43FJQi3HylsVZP1ndPDmWl83Ik1T5i8Z99
nho0v5XuzxOwt/H/lbxx6xMQAVEw0rlrKZQEzANpro3yC4gr4JQZFoPx8yfdYpfw
m9Lwmrniidus21qQSwKbPwwKTC5iN8KeFpalWOjSd1Nk4hFVwaTvhlDRfrebsZPu
ymO08XYaJ+MAYn5HCtdayFu94Oiy8LuQW4AZL474IMzUDbKrJqD1gmdc7Zy5XHE7
I+W2H9Y8b6TSCk669RZoxao9jpWZgrNG6vJjEYtuYKkd4ozy7cJp/bV7y8FqI6Rl
MuIEYV3m8pAPXh1BOaxF1EZEi49H4gDOWz+Cn3KUiuxDkEPrss0X3XLZXSmPO3ro
XzIPrvFZzH9rr6Hqw+u049sAGIKytkt4b++3yEvjUL+h5Q6BnIa2lqPdxja4QR7y
6cb2kc7bwoqqEFE/AXoC1HgC+/29hABTEThnXUfHX08DWqDHyoaM8/QzMvCo+AZA
zDyAks7KwR/MIjIjxapk1R33LuAuQDm5WFDYuqWQDuUmG/IxHxpVTqHh5t9nQZlE
LnKfViMFHHB4nb1t3ANNMi15ekr4M5HSXNBRlvorRuUftnBmUImDbP5+J36jdJFK
o2kQxL+fuQEmfKsfj9XhWkSQzggGiJl94F793t2taDcOv1+iH/lGphHJr/NUUxZr
aGUIrrHdwLHkTorMdD1xkz5AWDRZ9/s+L53ecrQ7S8Cok9naZ4BeFfe/xLk5MqgO
WfYD2LSdrvGCHiPpHVkZTKlyHy9nssGbG3cFmimchDX0qTvlQAOWXXt7AYt+EDSs
pAnlMmTkE6APz+peBUJQna3lv3mp7nRjzW0tHdRS/oiVYnO57cDSnMzbYqx3My+a
QFiqXEsiA6v95ivA68wEJff2URVIuuq5V3i/P9JRIsSIxSFA8J/BSuF/NxoUwYrz
8hl5Zl/rEwwvAFq/9Td5npV+3W7Urzn5nhXNd2uyxegAELxq7YBit6m9XO4s9Vpm
HcI6wyUPEX2lIw4Gzm5748Q6XOMIV4K6D01fnfA7NCbUgGaux0ddPYWaCiJJvrzo
I3I4yaLOzLFNrVvWlVtHK/L3vaAMmk/gfPxnw5HCn3Bseq7DvtKpuWTV0qG+RrO5
XD65uDTf8N/jUrzgqjmW+Ghr+BXeM2QkyMARz2ZXYjZrPqr9raLenkUMKPhx5PV+
T+s1PI71bg8m5XjhNztlPcdYzeYCAHVXqStCJZLVCxX5YmprDQ7WZrp9v9inUS3d
LsFiSuTElhZPOmbFJHQizwCxlb1eiFVQPsYoFVCUxT0hZ+f9uKoWvTdK2So8pXbx
Ee5INU/UsganNkWxbodXdrB+uT3ym8zT8IuQ0lnKuj1iFkuZRc0jOrUbY/CzQprS
Ytdzw5lZnxoRUOwfCyy9gJ8MVBdst/nFw3R6dR2nzgbVeCO5dhqHJEuFuqdw+xM0
N2iqEuQ9Vb6rIs+6fPuwkeyW7u5/XX7rKBmgc74/xPiC2n17qP3J2QSlBIurtSYT
dF5em2YNDZz8JBYYJqK7m7LKevETzYuhmAKwts7vWtZ5zPI3Bh9ra6sUhqkTW3BN
M+2abwrsIy/c58lvIN/TScONiyHxAv7L+pQhoCgwEmxXU33VUsb+oggJnqwXRsqH
1vD1DguYjCq9iWM096Nrt1Sw3466stq/ss9Gyx+B1Qb8KaR/d5UpQjbWdf5j7w5T
f0ma0S/9WZIuRN5ve0avHxBpgYFEOvhVNOeIwjquFeDVFw+arEIbGVKAAfbgcELg
ukQX2wCWxzR/8FftA6ySYueMygjRfAatr7YWMzQsFGlT4atsPwXnwNvfTqKDhYaX
ueBHegn0UL0vuOVUrmDAEVpAqIrWvzr0VzFP8uxXnRn0LR6XqI07rZbvxd0zFkxO
515SFeUa4m8bOvqxPzLu3osZZB4jrTl+EWQpdhgolMd4sTbBxGvxCL2ZjlQnw+u0
DXaAZGEOvIm5hCAApRM3vHOB3eKiBZAam7MmECzWUvOB0bU8POWgWvohahIp3dPK
u2nb8YdHzq05mtZjXA8Nt1t4Vt7X9N40+11UgNj/q60J4AnoBjy6zEy1hkPSvGJ0
hn+LmiEtotbfDCT6xbc+UJnBm8yTZ+VZ+BgNm3Q9n41rVgwZvkWEzahVxN9bLegD
KEpA7aB9KSGmbfJHaP3rk3QX6FMwYS97ZcGMNOaoLQKmJNayBtGthyutjLCEabzC
919oE9ri/cq/qHHT1DJcyGjFm3mQqkB1NA/zeZ/zDG7fJlzEKpaZxtIVZ82G2eH9
v1baFzr5c/oI0L9YoB4SgivszLHqd95XIvVKur8Qf+2J5+WO1vDcS6oF6UZBfcHH
8RGE8A/F2E+ZNTCJhuwox96fZttAkBXq2Ce+q5xdu3XWT24EV6bBrIgD8kgU6nUx
gOun2MInf1wlZC5iGtuXeTQXig+7JjtVgt2kQqRk5soto8i2+A+Pnr/sTWcc7ZOv
xCCp+RqrwE35czIXTqpV3Lb+pvlMJsq0WfEkHsJysowieK/XjMtQXXPchjNtQgsJ
3D/AQGfh42NH8WGlt5wjoczoBK7MiTSlvu6ATlDJ74JUo38fj88ZL0G13fHlJ63J
RihTtp6IaDdHB6LsN6mE7Os5NJshuB/5xuE4sj6b8oFZozLV9YQFjMas+Bu9nkof
p5bLAOULyjZ0gTxEGU2k41wZOtfvHdbpuyeGdt8+jMBAkRYlVBwOSyR/wFo1Gdlk
EFGlIkSyyGc4nPoga/7oHM2eZFD/PK9yM7daOreQarMqS+13dyNQI0K4+OUuoPs+
7yDQhpuEzyMEqMnY5OB90loW6yarTnZLfLbrweQe7x08YGCxeAk0N9VvH9GOQYQO
bOQfIrlKJ0/gdIeXGHkUL/THLhey5e4mF6rjegKKTM/e3TPKUqF08pwgN82HWC6q
jrrb8yl3aPL2dPJ+8v4Dpeat7DVPfvq0/4JMCJrKIUq8DHC85TP1afsEZuB38t+h
LX9BXxXAiNbFWE4aSA7ijTJFbTl+PXf9iTV4zoM9SPY1B9q2vKq34/IJLM4CyQnU
sasDMfBHoLNsf2fdS2yizsx/tSiso4wMOkm2Q26ljTBJ9j3pzS+gXiktYXt6gIJW
UxARwiehXYt7dMRnLBxfhkcuaHs2qWaIfDhSbgdyEbmcqHSXNsrhrDteyiXTqpkK
5X7mlOUGJRUJpg7HF1etROVIQ0qEqEny+pSeORG3GKEPsNvGeEvcLMRkX94+Ro0b
nvQR1CmQNmzqQeK6jSNxNVg4ZtBmGUFpkAdtn/fYCR7s2W+WAOzSqruTV4zFNq0r
AxJPLsy129oMsVJbS2ghSTpcbzAr0QM8ePM6SX6nkYuMma2caskdyLPLfHsoNnOr
WLBeFkrS589ze26GnLGh1gVSpxpD3GKLMq54c972zVHuy+PHoED13h80oU5/sMy3
ByAcb8X/Z6mgVIx1PE54vdRWwNzKvcK7x2CXrnlXhIZ8ApN8i7LDEvKXPQrsiI5V
iOj5nipMKXX4MRzyRctC0AfsQvfYYmZagYs6c+dPZlsOu/3jW7lq8OD9Te6UcMtW
p3YfqEwrwk52M0atDb2GtbGLcrx/SsKpyXhjIV4rwtsxDNOOAIBLM4/Fc1edairj
lP3LAwNDe4dtBBPZLUxRGKP23Z3EDJzoNLHjO9efD2wsS83BC0mcVZqkd+TyGD/E
CHr+mSSAknlj4WVy8o0xp/Ld9Q5qNwB0RvF7/qYz3aI5JjQu/EzFZbj6dZbSzo47
Opd3JdCgt2aaNMZK8zraBBaUWYG/0CSm2RCVot2YmesTHB/iXYBWwLvZd/qpUI/D
xjuK6/Nxw003TDpA7OzIkOpMCW6fPDlQAArur861utJUZqT14NcwMsWpnuaKloBe
vimIRSfXpYXUqTQlmjM9vNqGedkUNS9u+6VYgBsSs9/p/LS8KbOpx93Cb/pc7mgb
q6zjat9jbZpmm1r+TSVjV4cX4Aoa6KDGpnS7fQM4juYGVTJFAa6M38KMJAhdhbpo
1k9FMz0Zl7OWnmMOv+BY6Vsx4PUAvDwdpqh4Erjo8KtlX3kh7wNgkeEI2orWEP7e
tuDD/xca7blPFFwOsfu8olVjXhQ+iDxy0Iv7W/AvoRr3F9xPid7AWglazHsWQ2Hw
tdb0rihu3paM03VYYEgrMFmesW/Nwm0pqDDgbJA1gDn1ENrFMkzMOk4Vr/gfl4W/
26fvtfRsCMxiwJt33i045TlPLMbDiX7iWDELcTTU3JHamXqmrS6BLvgaUqcUVXpc
FvHitAoPdv0MRngw3mkhIXJoqwBmu+aOZIUTuXXiFgWiT9R5y3JHazIBjIC7G5Bo
RsaRsXTzVHmWIcHQuvNVu+cr8MgmaEYiQpyXUggoeBMvrcxy1S0KG1bEG1PFCxr4
9OOjE65nCHGo7gRzGMUnVAnKhhijzf0bfS4I7mGeMa9Vr+MmeBX3MiMMv6gWNj92
2iuDVE4k3wuOT+dS2Mu67x7Ted/6bzWTyAElvU4z6L7u7k7QXdIbFu6ls4h7tqV1
B4npOM7Jqqq7TXPRZ5cmnsgkM/md3Qr1cqMhUbnvbiUo3AK4c6Ki1Qz5IEkqzmC8
KlLFvKkKyTAArUCybXDwZAY5bzMSTSniZazMbwcEJui7Gy1/rAgvxuFptxrSCxbg
MS1xv1Oefko84G1AdgP7jzLcyyU23CwPiHqN8Skof2p0RX5KLONPWcXGvr4B35TV
V2ptwd8oV+kOG7gu/aglIC46Z8Dobl5xIxOZpwFu3KbuUbkPJzqz7vcCJT0hYx3w
Wliric6/UYN5EOBh3cYI1HpYlMVSarLrt4y1JtxMQ2kmmYKRO/QEHcSKrSO6uTvK
RZeu703x7IyeKZb2q78A5YlxjYjpcXcADmBig4Pk7oBUjACKn9Le++05koVU8Hpy
HkvF7MOQSHUOkORj1I5M/qebFGZddYF3Pl3rn6tye3V+ziYEjwa/qZAB6EI2/8ci
ALpGbPC+r1zCRqC3Y/YFKj7Vk9MprLXpf7bGj8lCQd4wGEiojJIEq40M0f6FdyhJ
l1gzwUbYUI46oHzFVt4KEPVlipLNYKsRV2YUmjVlhFDXfu6waq3PWm19Ei9ppoJP
Gn0Vs6ryYi3GslFw0YtSEQh7p6X+v/kMgDax7BR/vaCcfK8qe2cjdJfefTDps5Zy
VSfwtfbrldK+IUrM7Zzi9prSx1/rvCQ0+GB5WEhPHo7ultsmN6LSdiR8OMF5fA5V
EvxP+Kd/203dg5Fd8YKoJcFN5+DM0/gJAIxdKaMFPPfIs8p9qkMjJj0NJg8Zz5qJ
Y0NYQYZPLrtmOGMd0B1wPM95T4JyickDgpMxFxlDamkK5d8eFQv4haKbVCBUiOqJ
wmg3Ombd6KZFQh5NOU77Eh/mzTL1mF6NqU9x1mCgsS8jrPBYQrgWXhPbxLrBxAzJ
+kwGdts1BGcgWgtxBy4bBbiivfxLWHmUYg2uiaLCb+CLmkq6kEKjv3fYTTztiaSJ
CAvKY6Y6NC7mfjB+pmijTkJvPECEIwSd0C5ItPPPV4fxzKUNtztWgRGR6Za45dKq
sj4QFV3y024zEjTfl8WePI/JC2Ti+iVKuOou9jo5CP1ic37H7PTvnt/zSsquozQM
fLRRkt9khN+dwulZDAvHzysqDN5tfINfegIosHFiCvocyrOm0y/hYmFRPeIVqRM/
QNMOiEXi4Op7jNXZC9CX2rXv4mBCHrKKeMVqthn2xAaJzb8C7lF5YXKZH33o8or2
wmEV9x1Xbj3sLcCWcZ7Aqm1mk6/vnw4poA9nz97m1pdti6gKZZgQemRSeCNTbxZt
PjZlfiv5uRU0w9qG22b8FgGUv6M+DySfou/fgJ/i6/Aj74AC8Rp7+Wqxz8LvB+J/
e/aBPOl9oCbXOAMxJO7+WakJ3bBr9+5epdUcufvtZs4Vj9/j98wNzrDV/QhMiNX8
x7ejFBvFOcRNjgpkdsoRj+66uURad/os1DjPtpyi13e3Pr9ugBJKqD0SgQG+hktT
fGOw33bOFMoYD1xX6fjj3eWoiBNbOBJHwLUWy0rwz60do2FBof4ZE5A6737S68Ts
QWOfW9Jmpc73xNK2IiWREiwfK5ohCoT393P+uZ8EjJgfellYo+dAINOBgbUrEzTv
89N72uKs6GQe7rpGuN7PH8JEQ5sfu5o+qdytmlBCu36fiG/nPR50KUXccWIixXyX
I+R9tR84NIZK85riVldSUWghpzna+ogXNaV8HaHCa6SFdJtifXqrDRTPkLiMayfR
I0TLmqxSOZybqGgsWiwvyPI6zQSMin9Uzr9f8BoaQRFNlBnxNjeXK+2VzuTp+dfU
/7uNEww1hy0jP41Zi2s0jnQ3RlgWdURlp22gvaGMR/5TvWcoPXuzRW6GK6ZWSVSE
n3u/1HOw9D8UoxHa3u2dAQY/kvW5EapocGilloOz77kDSnnW4IPzGIaK8efxGM77
qRuZbRHX4qFu1XvoJpgVww6UtZ/OV6RUNM2Ntp5r9VEz5p57OPf9LbGRPiio0PPt
+1x1XofpmmbJv6fasgZCmHIRINk/er/9rpJD1dzXX2L/D0iicI8xcWiMGIvaUjJd
WYn72FrR4HN+IAQby/yODNoDY4vK2/YKo7fp5op91NS6hyVMwHkTYCSU29QO+dGK
56TUkp6IW1pj2vXpokJOn4dXRBdszxeQF5OePWduJ1TYa/BHe8gu5zilAv4rBZBQ
AWpb2k7PLXjyj+Kjlw6bWPAChBYO9x76oomtG7rrOKmCefrth8lAGTgODF6YixZR
ytkB9+IdRHorZLzjts9LjX8wEW8spZwPHI0rubErIMm7U0sbbPmqsk0jA4pxSVip
ND7GaepRKB1vXbcEpuPX/rQETJ/2ES5nSTuKqtl8V8h3yJu/TApTnPbLs88Xsy+5
LAVRo1KYctTueTpwuNzubBLTi2RehM89x1yUy7GELRFEKZmo7JrzPizXg6BD4y82
JvIr+XAeiKG1lOTPzNGi4l1bieNJd9kXsIsinpMSWZWYTFce2RWz3tbEVvYOlcuB
pKe0yB9jixue10UmBdKfOBS4GlMwUAgUix/vp6aKfeHen44ZAkyx+EdG7SdYbByl
RJQbRJ6vhQZyqhZIdCxys3G8COdmlNOdDAjCg9Llj8yVB6t17vWAMVuG/45NeM6v
XGpPQvl0VXi2qYJ7rAdcie/WSJEsMkc8YcB0pKxGbcxh/BFSuFXcTmi/GNuL+l6O
/GH7EgZn943n//gqXoE5MOMiAJzU+GpdhHlVo8yaBdRPfmjvfnfe5smyP7hRrhSm
wSE1LkeztvoXAW5D8s1iOHgIliBG8XvuVXh58RbnBpzNn+Gmmu9QMHxOlfmzwfF1
1+RQLkUNzFdYS0l9KFvUy39K2nTZwCJqkXJyrPHOfaRk0Ze/Z5kc0+x2Edq2TPjC
knt4JgXc6CjDoXe+v9ehb21cW18Sw7q2eWxC8Vrcxswj7bzzV0u3Kfi1Rk6PvwRF
n/WLRX3Q9rCKfYyVV633fqPPmUaQQIf849JLgyLUKxIMKUCv1Pl/6WLLmrM2cB81
Jn4oISlMj8nQzu3kXmrY8JLuAAb7OMWdWLcioqWT54/5/JaqIE5gtFfLeV5UGyGu
bw24gohv1/iEBRdqwe2cTyvxFKL2U6HM/Xp7i0QfNUWhbVyckPajFARq0sNHylEQ
3vrt0SiKCAWElAszwyM7s/3ePcZkh74CnG6Z2w+Tw+Bxj9efIfiCSdPJE+wLnDJM
h34XV4A0J91ppNzPjSTfHNfd2sZLyDkR8mti+VsN/VtUF4erqettouQj0UhcWkca
9+uJcHewSxxxQxDJPqTQJdQLmJoxXx98QfO0rEPCgglOfCqeh+854X0Fa9OTpGQN
51mE24bq/Pe+Kmv9niUXTatmuFMK1c8Lsu7/Ucm79iNPLhNsi7zjTyN12VUIP2/A
gONLSLIX2alE83eaUpoP5o3XvF7VZZuymrtMRweNh83VZfuoiQKJYmn3Ylh8NAsT
dhfZo+rWcnQOt+0tmQC6Dpfn5OFyiCAuZ2B6jdvVkF31Atsxotv/mMTxLl8imAUW
126x5hW/FlVzIiotHO+9AXdovyriBPykALEZ7wyhgNnYIz4GqdjdS1J6qiZhyDfh
ukeUjdaERRE8tqAVklxLkZ6GaSGD2U8yW+WRi6ImYWUQeEPm7Qq/bZmbfHG8EN7T
uKiT0qDQBajVX++VqSx01E+yTDlGwwoG/AAdkqVHtEGjR4CWo//sAc8YMQO6Iyqj
IX9Mhq4broOoxzS06Ezz0bswyGoMMlvZSOsroarl2nV3WEoFlkO4v8/QgheXlZ6V
hJtriNwbARV5Gzl5QTiRcFhl9vpdcqP95IJuKIqbgMvsqXLridyNphBN2AtYFWzR
9KOtZTu3dNRN489ozBXQKRYCgeR5npSEYrmqnYr5RqNyaLwZAsEft7uMYG0/lEKF
jtIFhkPIJbrtCMUMcJAZW1ycxPfAiTbGgM2ilNWU8ntBFDCmbylwLz3KuplWsUGO
qpmEt10WUu/RInUdLFPzsqFKG/CH0yMX/092Q/jXrB/1ZEyifuh4k6I27UufK5Kv
IZp7NmbmsTrW/Vajk7NB0Nu6O/lAoNDeB13KI+ei/l0Y/eR9ZgzMEBYEVaVAg0DS
s2Mr7Y5qb0YpEqV8yABQBU1vjdyJ5KI61Gl+SbG3+pSiG5r0SfBw4mZ/pOHZrQ0J
uYChLZiOUJWGsS6pXCzLS+bXeKrdZD9Bt1uqET/bCJvDXmdIVCpyehCgwRr/wZBH
ManQnnvMGMIao13zc3Tu22zJZa+4FNmi+fjb/RgcurLCn1aQ6J0Qky/pERBn8mk2
fwnQY6Rcb2fNwLZ7shKWoiPrgPsa6CUdKM2a1C+HfniyLol6xUzM10+6ciMSDjYF
fIFlCa03faK8X/3drFlbMGWTWQq8ciKtBfQCcvh0+3zPNo5/nsfITKcjNJxXyFfv
RzmxVOwH6OevlLwb+ZDkEyXluIM86GrHe1e6S+erSG9eAFIxQUP6ysS+ZW+nOV/b
9tsg6nLrHAy4+eqWT1bJ5+EguZes2mNfE3tGQLU9Z7JhH/uxgPeULT1xGReQw2g+
7FleFUa+Pk6UqeJK/LtMmz3qsajmp05bQ54SojvUbD4zNgzgm8JjRZ9FGVEYokA4
UG90PlwUQMtz9BZ434rL3EKvyOXnBpdQSR3An1U9HXrM0aJjf4P7D6+k98u77MYz
O/yhwxO2AwL0CPyOW0MlrRTF1a/FZhX6BXpb04xAFCftl2ad6hihwaC6UXN+QMsK
dr8h0zBb/mdHDOQVBcsKbGLJtwDnGRgmDZPQMYwjGqyEVtVZWgMP/NMuCjgCKoda
/VEtjCc6ujqDh1261Q0o+JKcGPiS4q9VWpSSWyzsUziPgJmHRJ+ureNlN2EDSfXJ
qaL8ZWRcmA36kmFBsLtqkUxSpG8j7PER/GpPnIemoQnYXKwmSgxZkGmZS1MO2w8r
8zLamPV/AUR7jNdWp5RsXrovfx6NOHc/KmziC/wo9wPYzwUG3dzDle2QvKie6Giz
uyVWz1L3rqSqtfCtkyzvJROx+t2quIV7lu4fEvSq2ZuMI0S+8IR/qFIY7D92OujF
eGTvQjf5bMEF8jio9RQIo9qN8HiE+mYt4fq7zgtwUkTjeo3QZI6TGFR7ba76FUt8
+4COiweL1m9cY9PE9IYuCUPL421/AgGSWfy/dwD4odtEqdfKh6P/nNIV+ohvPmS/
fHWh5NiLcEOiSyPqJMTJZPxal9OnW4kCzwBex5XPriveByGjSzp3sJP1s5gOV1O1
Yqc07nMSfIjqST/MFaRFVCEBq0niwH34fWopKTE6CbN0c8zOFv6Gu8f9joKbwai8
A77QzzTwvgbfEO9gTgKMVexuodXacpI8j+ryuZ51PS7Ru3Ej/5j3AVaQquNX49Sv
Mzpg0PZgsCAsm5V4BooOtV2AxLbn//b+RdZ/urDtNZuNnUCw/DHiqiXv7er7wRSr
TWKTHK2msSYqwWcKPg8MycL3vyoSVJA4CGONduW86MuUTCmDtGcxDHHp3JakFNnX
9gKD3vlpr1g4tvwwg7iafR18ESMdXIQ64xXOj7+QokSpHDIOJyBx1bSeyh8KOaQa
1d0exIx2UKSM8TigN08/LXIY2OEqCx7O4x7yo1rv0JMb0FGs5fryyJipoalwuATj
0ChhDhhF3TR32vEsDH5Urw3a0sz3dZHh4M9SOggefb3gbWNH/TFCF88RM2P3ocWx
/hmw/UVBFUDzBLlYgwkCen+37wLyVzJzE3vQ3hO82RE/F1KFZ5AXlaGQCKIZjuWf
RBiOuZz6ntR6+33uhlAg52l57K0xqgEn9hdBUGDd+wZj4AaF69SIh+nt3IH+wXYP
TGoaoETBGjrnIMPh5HsnJiKCMAlizMhZ8mrefhYHWR6ZaZ2VkvdjvR9DnyoTPVa0
nHtoSYO/c4FowVM5xdmz1tJ115U5aQdEtndzRofozdNyEGgkNWJ/7JNz/mU/qOJO
UCCEVrqCvzA5Q77tPOu0z6fT/+/NTIA/2WZFtLATsb8DKQoofYJKXGwDWJmijryz
KIbEfMhI13LA/YfdY9h9oBoIvX2THPn+vwE86NMhbRYgxnM6J7rK6zz8IHixlLL2
KKmmS48hO0DuMroxBOxXuDtZ5foGNCkU2StkfWs6VDGT2S0bgqv7N2jm5L2dbTQ3
QixdGK/d1P5ZOD1cITagOY4NhLF0O3ilkN0mOUm78VTYXeXCsvtwulQvyOLYOnCq
tMIhPaZ3q+STc2YUGOnp78YP1IdWNe1+FXxNxUKg7dKbOyDUlbDOvXMWtNvJFhK/
JeKxLwajBkIMjYqPFGs1gJ1uWmliMKQVVWX5DttolYbVHLJxlq51qr+tdg1cV/sv
HyZIdYQ4Ku4ExNjf9+kLU3CeiBUSmxTJ9KEV+L04wt3do2AQc3lT/lVhPYSNwAWE
KwTn4IoDIKQgD1+YRTjKusRRTIJuO3jQMn4pbe2TuyjRpTLGFBPZU4thSFcvttE9
CeRSh7eGOiKkM+sxEvmqJ/lJm7D1WRkrLSU7rVRn25TUWy7TZkfychhDynrv3cdJ
s4BszZMeN2NR9pRMjn8MF7eEcxszxiWzTe9RY9wA0al6aVshBUB4GV+5cL6AI79C
wE8UEk35UdqnGfZ9CBwLOpUd+bcWvaNZBrCrqDnDcfDNKWfBV2sC1Z2sO8rYE7wI
reQAXUf0C+ghDFEei4W7YApBwdO7wLFHvCDhrQ8WFRR9TsB5bLgVv3V8Vh6Z+awu
e+HTh2Iz4rWkbdh/xOjfTHUbjN3R+PzEUwdlIzmmzYON7fw085MV1u7SMEi5Rzft
bLGH4GgwZVpTsuFsiI2SU7WFeGj/snOljs8ewMuLmVg91PvxPStv8XeSt3uVevfQ
0O0k3MqpqpOW+kQs2yTDSLeK9BRRul9Ve4SIKKj0SxVle6nJUxPWoiY5odrhq1UE
1HAKnY1HKx/iEldmaYj9zM52kvKmNmbygGVHuTyQnKtb0bnr8L1YQKc7ivcsL0J+
21d2w8eVT4P+nHJKbGhPvMzw3x7VxkZ1nMWQwhAtXVcR3DWedaP8Epc3pyrkHgFR
uBr7siozA4YL/GmOvvn/fiAyoBg+VwI0Oi/ACWDUf1azQxAeeLejhxniHL71o2Nu
zkNkFAHQLfEVuFiY9+2wYZ5oKtltbbezobZ/T37Mi7bYwOuglU1LWGvldTkUJdns
LVBRtVmXB41P7QeaNsBJEjji/Qs+2LogNxphWFKnmvIWSehvm4PVjOzHURpQaZhW
7NxQmmm7/jf84DR7IJoPUzVNhWIosDmpUN/JL2UCScmrYnibbaou7ZScEaLQrLXq
3Am97NFQ3XxdF0eDHKkcmuI1keYtPXaA4ZfSRZIGrKAqXS2Def8wBqplEniIGVCl
++mMi/kHGMsSckFPkPsclYS0TgblWxYVWtL1HlZO8ELponCksSdbO3iOwwfbQbHq
4X1j/Yn7JWRbslhIGFjgAGnoAApVrs3bEcmQBz667caNeaIxjcfKDcdMfjbpd5ia
mo9toKgwUOJty9bkuI3TMVWuqVkbQkhH9EHW0vqYn3baAM3IsGOcJO7T5pi0DH5I
DqsJsm2o6axHRBlgk6j0Jy4UMdXqR5e3O5l2A8w7+XmLaiyP0+GOnZpxlNkc23bo
P63E+GRrfpB2GA2PmdtEZIh1vrAT2nHBziVDP3QxCvFr6V+ARD4xMHl3vg201iu3
T/05GXppuvN0julvl+V9ZfSruVa9W6nufHUtOcrNRp2nlx6cPKKe7Lf7vDRWMqxz
Q/2nFtSWzTjOhckaoqeBom+GQuwuzPRZauXItByXvXNeKZOR9fOFZJpN9SVhBxYQ
gJuQVGzCr0LmJELCAM0nN5nHCWT3rZwslXHfkyKWl80Jm5DDPlXWoymet8mNysAa
Z5+Y2a2apnHuVgUr/x4cSbqECRlaDKf2utRRUAFy8OPKbHSlb/btDj9Q2D5IxFPD
7hZIHK3Z14CwvKhxuWvNmoGn2n4l8XKgfTxhVFRQCY2XXY3F0RykD6+nlqB2JLQ/
+nJMKaouHQFeWXlXRzyliY0UYMSyYBaEkgx6cmz5nzW3ZRL2R4fGmtCcDwYVRKVP
9ThdQzAgtTZ7A4APR1K/2KuEr8fURDa3ehH1LJSOpkARgAck9DEK0RKJP4B4DNRz
nyZ7GQBL0KW+bbGucUcZ+N4/PUW+nu6amATQT4CngmDwWPqjlXn5zgJiSIYkQT/g
rIiE8Y664KLuUbOH9SuZ/PwgPi0ShKt7+IZxGUGo4L322IxuZtqcugORh/ZBCUFd
fonENroyX3xtmga7VPvpx2a4hjEF/MFRJwvNIQc+e2YmRLOftmjEbUQ1CVikSjji
j6Y7+7WWH93oyDftVWIX43FoUQvFcqaI19nU+uO7CTy3dEapqneq7Zwh/pqT4aLy
0C6E38rtjzfqrpGdeMXhBGFTe7PoScguUeh0vX78J2YxcHPpkZqEecq9CtDOKm2Y
DXWV0RU4VKf9k1NRRwU6nEyA+Yks/L30UqUJ6aK+hb3tX1Mi3+uPZaQnjGz3PRWj
z0nygOPesh/979NLyfmkOt6/g73IQn7dCuxiDHFATsIMkEf0we8mw7xpX4hSnxpE
9jmKCjcXavjBTY6jYGB4qs3BDIPruMEKG19Ez+nKxY5HoQ9pb2p+utqukgJKPiF0
XmoqG1G7ruZNdNSpIjBwRF+Xpv0EEmKRAsfkJWjIxHwAMEvPWyK/uG9vETEzucSr
a90Ev8vDLrwipGodqpTf8B4gzncT+1SJy04jhdHEqP7MiRH39iKoN0ho0uUerOR+
5i5pygTdX2ibOOEFVJ+zkbOT9wq789oWjh7kiWvL4SBEmBod4h4F7DkF5PjUZmIB
OsQNrYznozJVfu6ORW4K5EMZiFUHX7rP9dAsxj1ww0M1D0DM9r1VvvXlCMPDAVew
gXR6FlnUTus+GAQTSftFHvyoifCMwgoUIVjea2EsyMb3gM/006TRrNNglJG8N98R
QpW95ki8BjrK7hqLO/2mFz2KmMqSEibdZuWK7UlgusCXNHmR9Q/QUi2xYf6B6ApA
AlynlTx4xwSDuL0Nqg2+Uwmj8WnvqnS5mrf9w8Dg9itmjSIhgDq4HB6XlZ1ZZKaq
alPdBkp/fFpAkygSI5Muu/uKRdAfftOezk+UWEf94ou2bb+Im/qHX70udkcAZADQ
R9lHLWxEkQDEHu3Sc3uA6JqgpJxflRVc6IJxFmU6/x9GvY7tBFLyDBdkNvGiYhF/
JmwqANn3W+sutKQ2qVSHqtqf4NJVdth8zxIEfNj7kcaDwbvpwsuMc/cVGsOn8tLU
j4pq2M66gHcnZ4MOKuDSjz1pWuzG8A+6vSgE4GWR6Z4IdigNCileXO8Z6phSfDx0
Xf2AiyUZ+ot3Jv4AbTFujTDMGijbc0RGTUFxwAoQpthiVit1cUlxgoVoDwL228ti
N9KrJXe4HVdd/l+qpSR8cd3bjhkG56yjU/s24Rb68yS6IibfQ9CTFS/xYKGLjnV4
M638WfpOg1MDIEQ9ozBO8pnO5cvH61CwRRX6eLjLS9lTzg2VUkRWVnnbMOTkDPWJ
9fHzypA987cPQUQXhySK/ZNhhh7u3O1rJcPON9bC9Qrum5XpwfnITGF971rrrYGH
mkaEUD9Rij2J/dXeJu1E57JmclvDNUaF0+gKHZ2VQjGdQ1+eCp7bLsF6qs/+1E9+
02IJFvl9rE2tVxgeWFNImqObVuvTbJ7MCA13IK43ENxJOn+zOPN9qD3XL+p1jlTm
eRsf/+hjacHqvCCy+AkFD96WH0pDxM7GX/fNlJauqY5bAszgo2k7j6PVEjH7j3Zr
c1w9y7nLSBNdl3dvlNQdAoISajHf0OuVgSfENdXDfVMhIGQ+JusF97Vz4UvDbGEP
nIpCR1nfiR/cmHwhRJXc0FL5AYhYRG/prv6yJ/idwJJxS473Kv1bZlZAwV2Z+OoD
N4t24MhVaJsgCbJJWxZyDWQ79mD4ur37A8GBF8uTbHy5ceA2vvrkhCiFUzdIL3/n
HkeD2fpwtBRsL4x1+euLtzlZ006p5q93fwnCBawsUI/tm259JV2ZTAOEoFEPchak
ZVObHQe9dYtn4F5DsIKgDvO3vX6lnU8tM5ejRuNue3Xt/M2GFmBnNZ+iBFmUw/XY
9Xej0sxBNwTXb9gOybAZ0hFlmnYNF8BFP3NWYUJlWG88tvaEbVjkAECi4GfiSGy/
6dB9T2k0OSyJG6kySAPWEypb7Mv0nx8VdcroKpjnVIFE2SDGAiu83Gt87lqoBthV
bJ0y9xs6Ycu9fiDDM9OQ67x6KvZEQ92pX0x2kFszdzWnLnKZ+uFe9vbOYYx4ecMC
7Ys4dcC8oE2b+ep+mxmVCo/r7NtyHQY0Mi21cvB4wNdlsDLz9q85zMNqYz0rdd8j
+8SqigMoZnWa8sBmCkmKzcEpACLPq5209occ/TO44vHk3yQBjT+8G4cfsgOkA8XB
eJ6/DYUUs2R13olN8jTS7BrLhkpmX1VIMFbd0Qh3eIWyAF5M4cohFpsQVz7BkdGm
bT2dY0M9jC5lLK7VBpKmmKSedFozF2p9JXBZqsFlDnwmI5w0Kb7n6wTovfWm6FQH
zlvI8zAMuJ3GzWOxGO8IgnOmGqF/WQJyl8r9P4p0phS5HWDC0pQ8u7qJ/2x5C0R2
vdQzSoJworRFtX6dbhp7eW1QMW4nQH4XkpZSglB//tETbweKXYX8muTeIypHxpwa
G4sy+sTVCPn2NtGuyTIv9XnR6NDJ84YHBgwLy24Aa/TKArwYB2dhH3eXM/wLx3C3
QjDV243ThmGfWLdo+wFFH2S1yp08HS24HdFgWamjNDhkKtZHPK4Nkmqx6/bQ09gD
p0YU7elP4XEzzmHP0ONMFY+PIbdX2N0YLqidVjhTc1piUXG6Rzpmy3tuW+t2hFQt
4SZW4ItVwGHtVIWrDBkiRWL+twkHwx16I41ODUZ2BlsT0pWdc7Uykdk52QV0YyYo
DdEd6tdqwKW8XY28BPfNMDFvhFPPXiqKJTVGDOvnrEZWLNTbcn2U2YRYF3fTpMjW
9p7KbnkPMijFpLA5TlEkNYZiVkWdNpkE5u6FExbX4jmGDzWnopDq540Ldtq7L6Hp
KnJXANOs8kopzSNTyj6OG448kbhY3CHJcsD3ZhT+XVtbQIpjUzctDy8QzNmPPNTo
dYjJvU47IAOtbh8dhMtiG5d7EwhMDaJioZJijCueEjceFkNDdNvp+eX43AkNswDu
Z4t+YyFLveyhA+rhSEL3gK1jPtA1+4WzGF4pVTmMA840PmRV3yJ+CIuJC6BSEttd
NVJa5YmdrUCPdR9uoHxg+PS8bvqsJHf6ALKdzMARGM9/kAXaIonwMWiEkOstJ4qa
Srsih7efEuxACBMD6vzwwKEtkdDy44lC4FPbNjwV8w4K5tz6V8ZP4KUWlCBEdPvo
o661XRqK4m+LTDeRwCX3Y7CIhYUQ/Cht5ZxI+KirLxvwIsBy+4wgZCfVLnZPumXu
OWQkghCrDvxytnLQeDSfZ5673cUpmrvclQ3PPJGVp+eTgYiBHQej0Qm/93lO1dZK
mIcahskyBezu7aF4jbYXZEeokfQlc29igZkJEVrrv0rjs+Hb7X8mSVOSJANkdSLJ
FAdeHeYA4XfqEXjr3luO2BQNGXsoCN4BDiY2qt6mdRnWfN9bPIMY4zsqIdaolsxn
RccOInFUNQEE3XdfSG0kKFRL1XYg3N3Mg1CRuSBaQtebj7K+Zt0biT5MCavP+Lxo
Md+J2lHor4kyeSxncSdmC1KF7lWV+SZjxcRJjaxzfJFO0AbQqY36D/dl5vlePRMv
EgrCXgMfokFkojFoOS8oliKa4n3k6yFkQxbTmdKZhtK90IaiEKPw7sK7WuCitjL4
QrAV6Pua7kis2qzKgfIIHZNs1iNjDejmkKnsEcm0rE57NNdMUZLD2MpfF/noqmcx
QnxWg4+QWSV7bwdR8M2oFFQ+pmNSqdUv93ahzlP7lajwTe19hgFdPhpnhz0kL8VV
myM0pmIwghMfRQK6OUx6SIno4s2cPFCxSWZ7aTjXCEdBeKr4QpTWpGPO9SqYGzkQ
1ZhLRc55cvOYYr8ZCfE+RhHLkjyVZLNGNqh9OpagupzQUWn8qGcjYIhyPoS3vc+m
SGMQSOdrKfCpLq1FqAPjtas9tt+hs77852k5rO+LtKs1AiWEfMdJvorbU87hySXa
LHr/90Ujd7lHqmZEB5oWawyd1z4NS8DLW2QNnwOednv+87SqvB3darwbsN0H4As5
2gCsIHNgCcEQbOkfLWLDfUXXdNZW7Glp0DW8W66/d/M6ZQvWqTu0Fan8MohMhg0e
SM8il2x11HLU6GeMEybCcBybNM5fd23QG4t1P8uUi6SDd0ELUff/xeusnaXssixc
kiil/sxbvNiPQ+h3VQ2aBnGIFUdiVxXDEyG1qUTxoDRkwPB9NbvEpLiuK+0mat7L
ZFVvjmv8BR34RlUXR0Tt3lCC2ZRgNQ0Ekpbcx4to+qooMIqBcscTF6o3oUw3e6SK
bgDE+ICXB7Ar/Ojj3CZS8oL+pTSG++eT5g9ymb9t01Yx03PplJf458r/VPZCmDTE
o6sC63yByzu63gIx7kIi210EvHDh1ae5Wm/vilA6tYv5xaSUH3mU7OPI9GLyvBt0
4TosvNBqSddPo3w/IkEWR1Kea+A+rheLRbIxA4BLX20msuMH+RiDvVGeFVGTzNX4
26t9HNn79+BWBk2+TGbIWzZK3tEP3yAxEcdD0T0JyUyrgRo7NlFIaR4v2Vvnh90d
4PkLWm0t1v64XJVHuPedoQ4ajBBAM9V0WI54UxO4wRYLxhKFcUzIDZXF6G9xwbSo
XqspPtUy2J7tU/oXLG4eqvfAZ4tv0Bbar3zyAGmUvGI3H1WccDX7GX//CP+yGcor
KZrU3z1DBvJOSG9QWGzi+3Y4R7FKBJGERlabZrFMDxkmQgVRF0+hk5/te6f1sTMD
1gDICRXkuqu3tqwOE0tM7oBwxcrJ/yNS2UngjAhzt0Q6BQvH3Z0DHcpkLBzU2xVN
UWtV/jdCFykf1by7GH6iGg8CnI8oQoTVKQiDgm/nxu5E3QpN0Z4ZaT723ZDubyrT
BkViDM+LhCp/gA+FcUVu1+vnYlLghMIR2aj538SNIq4ku/6xn9JSC4pcqu3F0gvt
FUaxuG/MU7eBh9p7jmK4G7weTxouw61S2F1Efo6/QND2r0R5FF79DgWDk61HqeZm
RcE6Is2Q/gYULeHyTUE+sWzJNHY7lidGOWCBX5KOqfyOzDjQbU3+zGYLzgeN4Ixa
4Sj+lhzyfFXwZoYfrHIYsXlrLqiPmljwNDW2+3Vk2SsQXKPW4nti9RhbzvukmLdp
z85jNFPffmWPy6p3spDmOEzaHWBwMJlHaEjdlIBxNS/lwnvGEL72gqBV6sqml3WD
1dZaszNnReWinzT36WFRsydFRECpmpcESr6j31NC7s6iVzHZdnLh5H0+TSe5WWdM
pGogcVgnFNH3NnXcoN5SYdpZXLxm4pGNpun3ApjsZoDHhmiGrCR1gdiFQr/0baD/
TJOGllCfPgRK51jxeWQ/Rq689WFP0pj/2BRfpn+1q89JDHPVH5Bp4A5ZgQGHWFmW
7JzCSCODPEjJghsVe2KYL50mvZk+tfUroUhy3nlK3ahXPY6FU73Mjp0joxUf4Wlo
ROPIoJ2waWSx037830IcCKgGY/+mgmV/Xv4cV1fLSk/tHSg76CyT5PG27ymmE9az
NjwPWq+YE3MVLAwtLCyPObm1QDIDHW8lyPc7a3A9h3vpDEPBHvQvgfewy4IcwxS/
M3PlzlbKaE0SllLtytEjpTyXZnr6LkGh/xZQR+aWWo/q9Tapvx9zlO9x/VF0Z5CB
29b+gZrFZWXIxKUaBd1cQiGOOl+S5wjzeIQH+gUOqVw9dJtOIuoURa73Y1W9Dx+7
xHyFpP3xANajBMc8O859yIG+3T1gMj1P/fl5YuzWgFVOolPBHnLFzgG8HhXhRVe/
eN/AIRlQynhDKGJApqhK1YzrCAQ39LjVucMXN4sg0DatgyWvawjOKMhKRRonuam6
lPWs8AEp0D1Zqi8uWg2xLX7J7YkLtR+FMx4blY4nb1mZVNV+ftQwa7eP+G/InKh2
8XWZMfjdicaz6KIF+x/VZUJi9sD8GHqa65RlDkQ6+2DFKKg3mWTjPZySVtVHFEeJ
zEKizlO7sETMoNFPBbjPQ88dPcB2pAIkbNOCAa7kqZXoFbvI+aS8kD3T1JG7X8qL
Efm7BofzfUaFF+BcgLrt7c/SBl+d1YbZf2vAY8AgRItt1y/PokKoDd1N2rTQYwJK
gdi5NXdtnvyXxnW6V6eSS8DuhjAG0wm/5I5UjebvjYeaL+FWMOt9KFnV4W/iUym7
WbDOr5f1A3wLF3CoBMOxfyDYx435Q+VL1ubg5s2mp08xu7bjEU4+rLNPLJPR88Jb
6r9VqzXbt6Z/n2Zl67UWoefKD1xC1HnnLEyJsCcXmYWaWC/Okwt4YFPoCvIy9rYL
eykDmtfB3uM5z+QmX+G6DLHmdVXR2m0JwIJdSGU49op0iW6o6QrHapkTjVc7S3U+
HBS+iZ/VJihED/l9+mlmAtmYedHVKPnc8SmvKvU1+9Vsf6Kz2ZhccGOEJdC6tzBG
ZcV0cdmFXE6aU1wQJ1YZiFiVuwVatwquGTW0Ac5fWfDcRi6Z6zpHmXOE5kzhL/Oo
ekR1qxgnulMkmRaGkIrjaI3o3XKpCd8MEcPe8xSASjSa329ATXoKrV3zXqG9W6/J
ALWi9p8r7htP6rVhjIL3A+C6R35TvIsQ7YAXVmWEnac65qRfWXa5gMxMMjJyVh2C
q/N0RHkYmTcFU5nBQGeeqeMpscpBYpEcgIXwei5ai9hTqet0kNT951inflXhkJuH
Uhs4Ac4/jJgbXXr+0+OIpa/d2jrm1TO4KA8auVhZYuPUeZ6yoa26CYH6zagFGoKn
AJ46BhOLx83dgZXBPtIZTHcRH0iXofPjPPLhQ+ZoMJdQPNClo5WH8WLc3rdDLZ9t
YlcqB325DPkk0eNiz/zdJx7BxajbOcoHTCxKL/j4Mj1BlP++Pm3ECbrmPrHlTb2A
mlm/TG5E9MgCh5vXo8Ki3q3uJvP4oj4DygNuoDPB5Afr+aJ4yfjMMhXIAnL0r+FQ
4FANo9vgkLk6cQdLWalTZAMevDHSPDM+GfPNgjLqdeYBibBmAXWC6TgvyMTdjfsz
978GH6aIJCuKfBN7ytd2pCEDfcNtQ7xgJtWHdVJy+PsPV65HSdAYfUDvKSZFddHZ
niVzKaeO0UQvD87cdP3R8bHEsthrP8qzMZ26YTD4C8TnCl2aeY5Hz1ylklx4xShS
hFSTRvSKtvMTzMRn2DaDR6T5kKiueq94z3wlXwkldF9m241mQ4mBOPLMgt8I9K4+
XwQawd40iU+mBOkNTxTnTzO2yeGQ9P2Ufi27u+xmC5F/rRfqDYv+hwyWp2iPMRos
8EIkL+yHWS5cALyFFWJpDcyC7ah2OKGw328R7OAavFjaXGEAtU+xh5zHVu6OIlOU
BPt3eFSkc+VwSx3wRIzMBWIS2oq5h+bmS7yMBmg0EZjJ6XLxxA3bJ8DFVHFbI6MM
YFvOAaZ58LN9l9cZGitAowrO35za+XSKTEwhIldqHYYdLJIzdmpTYoivk8xLh7ft
SbeCC+/AO8D4MiF6zW2NOxsbvQ2+2Z/sa6WZpGxGGZliU//0y6YLogxy1ODnyxnr
bUdquKYupwLT4HUTXEguThOdBLudFHpwf0ANO4aDqqNT75e3UHpT06266gTdeT5b
qCI+VHodlKwgGK8Ek19DLxAfiZLnItozuY7E9MeS8IONS6LyXTGDx0OJ8GZzvyqD
+DsZKT0YRo09PepKYiho6FcWSTaCcL4Ys8+18mTOxv2hL2WCG5w3O3wNwBsXR4Su
/2Xk1dFlKFS9SFD+EB2hJm14Ql+WlhN+IoyvE7T/C+6zZ9KX8B8npzXHDKDAYz8g
1Uw4waF3P/ePTppQQWDAuuTyMgWbalWlZj/cM+r8d7G/oQHWNv7/VY2RFwj8+Jph
Y4N2VFJusPYnDtil3e2fLFV0dlnixJdrGUf0NFLe3XWraEeyrxewNYkjPRnoF3Oi
jgcqiTPikWMzFsoELiEKfEJDx2ww1abRHRfPyWyEOPehZmTCLnvDRjnuHCcHVORt
0VRmM+yCZs8vt1wZ6+tyOgimZCozgL+mUoJ/4CzkzUurAmGBipcJrTmJgjiuAcxd
4+gMxDRLYc1+ZYsoPs9ZkHWKzjpDdTJxrdxXgHi5uE4uIaolgrCHtixr3GySuEm2
6+HDrIB0D2eO0/AZ1GXjtyK6AOtCHHrQ0Bn/j0+rkl6Sy+KtgXzb5qCehUMmfuY5
IGcku7k2zlgXPVwdllGlozWxOhjzw/xKUnRGBNjxISkCaYNrhpNdspwB+qWMbkDG
NLFE5rgBnIj5dBDfo1rcb1VEkOXz4LRL7EZwGA7irgET0sOHcLFm1pVRCRxDkEM4
M7w7IzsIiZrsALSLPtNUNxchj9ENCo1NWKgactUL2WbsbBKr63EyPC53T1zL3mnb
/IxN8rNQpI9cLl6fAjOQk0+bayCxOOuaWNzT2fGbj23R0s9h/a/f5DJ43FU5Tahb
ZbM50gdv9kIc9QDiP/e93mjQxR7mDCEK7qpJYgTEUo/n+hw2fYDG28uu2aT1ANfO
dBEUiEm+R2XbYt063d2O7mSWw1+1yAGgX9tq7RtNJ29eNpYyWS03MG9qcYX2bS8d
a1gW+rysDpDaRKAimlRvAN2hdg43HpChqTWPJ7AJNUUW7tesIPvElG/86DDgU5cg
r7OLlIkbK4GGlrmnrqo3AWpT0oUpSdpVQvIN+uy2hKh9BCDH/6kO+B5pX/Kx3bnI
lKaM+EjkAuMS+xVU9D1vw1BjFhOS8XQsdjGVR4luGRgRI0nymtlRYZsJPT4lCskN
0A3eXacrxBUp9Al395/+1K5SmLo/60CXWavIUkmbkpqD0VONVcQ5u14/ruOzc3HU
3tzYkHSuxIwBlL92XVzT0TRwXPEzzi45z4Iz3vBBo9lBrA7cAnkFhScRSrdf7ZFl
uwpo9tf9F8/8gq8trLi33FUKujRRiVHF64Rjt40/LZeZjPmDseLhe808Wcf6LsVD
OGBLHOivxqo9sjTiVSvOZ775LOPASYc1vxVPDXFNEjmEp4ECgJQpTfuciCpW39uU
/hZONU5rk58IAnFSI4RvPGLL9mfl8hnr34oSLLRcx3YeAfXjnvN3faY6PLetixzc
kZG9A5iFbDuDQpvrt2jOE8ljn2iP9AGjNUw8MlNm1BYBGoYZQS4/oYKiG2nBxCw5
M+6BzBuxAWo1z03qE895P39pBnY2CrLwJV8A6xsPIuyUMGNW8EtbUagrOldndsU4
14TwoG83XUjsuKoiy9rYp8hcewZS9xzW3/Aq3Yed1NdQZtvGzGnefaocF7d9ECrY
rkGxbfwB2eglj9EsccmwuCZ6UPrPwn48b5mCy9k8Ze4HxlSZsQQhxVPxX/29ciJO
BZARN/Ay2OVY3I27col8UBzqgJGyWYLWQm9vBmSMat5q2T0jIbPA16++6lDxOEKD
hN+HebpkVCsj6hHpWBz7zaYyTicK55w2DZ+YBRkzl7aiQwa0Vd/gxcVaj67ij0Wg
/0FreUaFzG29FO6ClDFgNz++7WeyMsOZ/84Esw4NKymsvvB5XmyENhwyEfYscXWF
yKGtMPp6Cz9ADTx++ja6gQy3E2gHh7uxqs8u0xwou/VV6ri7wInDI94gA2PYqTym
SgipqO6rfn16LjUwn25LdDDMdg1hb7IbieSGLxGqeNFNzey+NYES1gJFhdIYeVmi
C+2ZhGL4yHp+7fyGKQBZK27YxgshDnYsEJUYTtmnT8HYVxeKNMKIOO1FIuc80YOr
vOaENBA2jS1xW5YSirl2Vcb+Q544QA9j4Zy/IH8f6MlJ2RjpYqrFk0qwpsSobJOV
yMsHKPQHUsFxzZ7X4xmm3FR/RUxxzrf9J2ZYMD7sa4Jb63AhmQRlxFnr3L9apF0s
YGorgMgpK4sUZJTZGC+1JtyPQDKZhnTlbX1D7kLSHcNsjitAYaih4boZ6q1OG6V6
BmPuTom28EX0t15aQlAp6YY4renJ/O84k2lZejW7I39WxMoT2stvECS8Rd5nJwoM
vZe+kO1qqf5MAgHAClLGY/VYUNBK2GmE0fgyMOOOtU281GDUXjIlz6twiXonBTFy
hRH/zurT7Oi46Lpo5K/rbH2gcuE+Sn5yxiguEHL0vNgk9u5DHc7sNrkdS/GqFEuJ
nkIoXklJTIe7O0tKnsByvg8GkpSktbhuKKGwKOzDiRNSwIav9MTUkOiW/LnI/7kw
7+I2zlH5xRJtIUenUufaYMwVqYL/KXvuCFIU3mAIdC9Ad/ad8Rfp+zjs/oeqlikE
sTuwMdmvJwLh1znw+MZfaIwNKQDP9cZMi0DxMxV6LWaBKjNJ3btU8lfY59OoJ9rb
X8B+YYr+Nmt/79JuMeR4Fl9Xa8HV55hiTxGFheuor+oE+Dt7gq4aonaln+f7RElC
iuKF8fmdR31Djhf1O/7Tv2+C9z7QaH5aAuiwrAvWJAHMar+WbBvtlzneWW8AHXOH
UmCf2jGHyp87zLH7nq9w2ImFKKTT4LsEEXD1w5dlQ+9RiOsw4aO9tFhm5a1HQNDd
nmO+vbn+aIgE2ID+ir5ac0Br+LKL84qql/SURtvbjs8DSLOg9fN04SA6IsnjR3cr
L5s0Sz+R98ysVgSWWVMTvM8A8YekVZZmLDddIducLiPIeNHjryLcFVK8HctO4i4B
ywkPReKSGqH2GlzE84FIyjQicu7WEgM/tyPtSWtbaBJ8038qjliMy3ZIozlFlH1b
ClX4CugM7oyl6rac7lE5DjsV466nwWuBDDiySA5ReYsw/GCHh4wn50XfyyGzwYW6
DHUncRcDThx5yNt3qHvLxicVpjuLpJdl1+LKBz8/oaMCdyt4ugSJg9Lvop3Wqvjf
kIOEc2XFY5kcu1Myp2d/qU1ymGL3usxLox4QgY+A1lmqLSLoSyd9k+hpc3v34KP5
YUIpTBruE1LZlYR7zB6tJB9PVqHsgeX1kirc9oQZwTE/fUoM6L+40jlLpF1+spjM
E3E6swwJs5mb4I/X56b9X7QrhsfmO11s54ozCK2+RWrF3htk533jbEXDFNzXkaR8
7UAlF/xe0baon051VLAplEPSPLr0fa4h2X4j5rqfRLuZzksxOSzj+XjEXfXdWXxr
fsG0Im3GWXPEOrXH2s36Mf/SVjRkMQ/6lu7iPQOOP9DOibpy7PS94LottkLrIN9R
paScVp2qkxpDUEtC3HVcv13VNgh1SuaRTNGRIgO6NWpie/mIM5GOalQgnM3k+4c4
P7wJ5q0xgyljT7VQawoxDdomx7jLVJuUFrjnnwMG7h9VVAeO24XfY/5spqeMsW1b
ZFesh0kittnqLCasQCVM6JdvkkWE9DeJZUMTDv9hr4ca6YQMQQCBhzmjaLfDHM/s
pTuZjCIc5D9mAXTJ4bFe0/FFNFukvrS26JANb2f9QJPc4dqlNiIRp5gtYz3L9H8w
rhsUvOgsc7myfc4rCBhhibB2xKfRgTLkov5Okdxq69XX+6y2vlYnaIySJr4I5IS7
/mizSHPy4jckv57E0pAMf5OuE1/Ty5s0DunDRB/ZdjWZ6XNGfWQBx08AP7Ssky35
cVSzK7eRYEAAXgZ0ySFEH0GF+50Hm6tDyAPQiMr7qe6iYteigl0nDHQvFq1/uK3H
v+HillfJi5orqxQYrbuL7znmZOGy4LBpxfbonWyDRC5XjdMLj2yyq9GEjY5PpvLY
lrHPFgP7xecTnH+EE0sjX9v2EA4cgLJl/amZV7LD+dq5UfVFvuKAC7/ybnOGv1V3
LmvNTTFZAt44xHB9eQkjzi67Kh2Cq2+uTHlNdPHX6sazaQ6U6D0WZfvggi5wudSu
ERDjdkB7LXk0pHCCBoAZBpy3o+71HvDqOq/tg3HXz/DtOvbw4ZSNT2onCnSIOvMB
hr025wq4B16Gd07FJ27arBYcGZvwJeBDlZLgJnGs+/yx/fQkpRxl03iBGh+ApIZm
FD1mYm3OF7MipViw1XFYSaY4JkEH/OzZ0he8EFs+x0SSShqHUBw1RAcFRPz7EErS
/T79klx5A/YN91i+iuWWDn3PyFUnP8hZEfi4VtyswbOvLTZ8ImnLhYEkvPgRCD/R
EYpCZLKi/yQu0JSxCa+IXIaNw+2sjtn07+fNwg9zLpdThrHRvg4/X4SvHgwcgXEQ
4g8PMUvvRXfw/rafdIrjtEhRCbC6JAMef66qYOChf0PP20ePTek6EgGrIu7K4x+W
JLXzs4xZYNSoVV280jRCnVLvpn8VF/HCq5zzXS+7MAdWtyKSkpebkea9HUTUMJgT
519zigijyz1yaSH+Dj5O/d8ofjxxOrFe9klEpW9HqLMFe5be7TqDETwQrAH4pvz3
KcV4KRwVsqx5Mz/dRwcK/lBppXYLvBK2mXRjKSeyjUwgjTFl6LSKkM1Mpav4xdwS
AhxmRjCT98P/N9aT1bUEdKcESsQo0J8HdVs/iA7hvn9FBLVjCCN7QbzjR6bxRtQ5
V8cozoMAF2HS6KJNewHv0G+3wWj0o+MB7Y/FKo6jCaFeLVkS5cIJSq6O7L6ZSYVV
zQ+DKpwBJSMXOVVl7p2Js4YGcPNWwxxjxczz7wIDTHQ/Bt6UFiVNKkuKb0OTHD4k
qwCjRwN76O14WqI9+Y3Yn1XAiConl3PbJ0P7bFcDxplfGLZuSsMCWP4nk/g4xBzj
o5AOGUm7+moZ7KQd0cVxrU1TDOm3owMrDHia4XXKTOZ+3VEeYmoyKMNnQ7fBcFAH
tVRHXmMtbxcL7RYXEspRrIr5fsplYlnmbc9RziaUlbjCCf6jC/TgWvbUa58RoojQ
Oz5GtTuTxgjGrlmOKEAnMYJ0v16oegQxpv+6m6mkUa/Q80hzjUshU51J7yzi2UU6
YMy+gWHlIoBzspI9kAhNd5px6f6Tr5vhM6/OibCR3IDdVKojd7Ls3TN9wGozkxDO
TkwYjlL3hqwc8vJgGGACx16GOKy4q/2UfiwqWZ18upUji7DVVsiuSwgwgYb32jlz
gcxxl9R+ygXjQK3zpsgVN4MMc5/sDrBgNJJ3Sn1WJHayXm6Kr8Q4i3Lf4pdoVUq2
3N4pZfoWNzV7DIKS1NeGuhTNaKEn+UCD+3LXA8cmCu1N+kX3P0vk7g4CAVUA+mLY
nKQycIrDxFzaf9UniSn/HZdOPio2z54yq/jgE4SxNPkD3lQkdo6Rf2OATp20apYl
qr8rAgry+7NbnKd7LSgFyvY6+0F2ssZCYZesaa6QYGhd25iGWj67DVhpVeETUXMX
gvTRbwDeZvDQdkL3EOb1Hr5Jx3lHxL7ugVepPAR6OSUUi2CXZSVc3ZjyXMSZMcEL
msG/NyxLE2UdoLnWjbMPisi8O3YeuSlrxcp2YFR4RekLb+/krZevCP1YUsND6MTj
0efm6npsxFg58StGIJniL62/Xeg9sX4rqoiibbik9M8K7Oyn/3XhLpU9RKprwATT
m32mZq7oB5KK5zIFltVObIz3GyAmk9aM0ncfcs5c4Do2A36RHJVorIuGJPmhO4ma
t1ECFa2IPTjRtZgKv2y1lYnDs8Do+4WBL8/kJGL7Q3ot76TPY9bfsChmCOefOGnf
9htQNMuLQquzbW9UvcBZLSXLnOfjK3wzUS04N0e/NAEbMPYtIg5yqd1126DUfS+/
DxlAuoghCpSg4rnOtt4dpK2N8d730FMkzOiY+GWERom5h5wObjRBd9LcdNTDf+T4
LsKgfJRmE3ZcCDQ38zZNUcKTNO+vj8jpW4K/soSlchmSYzVO+g17SjAP+FxY3pJ0
JcLSHWWfi7wpDFCWrBzwlI8ZbZ/C1aj6H8A1PGfSTXndQf5X3dsRsnTs+lVdb4sK
mGAMdkUbugWxbAOfjEC95F3/JTHTXWpkon3703yZ+hWis74lntXd+eieQMFURMFf
oXSV+tc0209R4n8NpoLvJdTAcg0rkHNP/UV6sVqZ1VeGZkt2uzZCPCO/2TRb9Pj9
kjuSncLztI5v0gxHuJiLp7GGMNlhGWgYh2jNf8QTUFUS1yzZH3+eGPwpCMLR6Mjt
EMmf9Y9/Ihw+1fazJrZyYO0XB0w9b0zGttO2GFZ4vTnvynNChWD1kt6HCz6h37+d
KzD7qd/FoV/JnoFyzSCXxhdBH7jodS3Uy1KSDF+0mEO77Tx0SSRrh6YTspTw0rR6
bNyro7QbYM9IuBN6mQyKHqPi98GM/jVp8/OFH9Bnwwx//0TbxvDoVGe6JhS1nqhH
GOuT8Te0pbv3DYXwU3J0Ug5VXMevod/nAoE15tdYQCG8J1E3GPIypIOSuCjXcKvV
kD1KgnP6Z1XDOlfDPcG7nmr/onVHtFzKToCKsW6dxuMBVgc+F50Uwa2UCrLtACrt
Bc2uZPASG0zQBcyFH6/YQDi+80FiuGjB+Q6+zyrVJ3hffsYX2HaXmFjcsc2Mkxud
qs+heLlFhisS6Io61A9Xg4LLTzqCAG5SslIplhDCFettDy0gf+CCGeQjn8hUVZJp
G7AwKJxGmv1i2ZxYtKBzwhI3lVgIuQrXiQZH+GCXeJsFfPJlTxOLAW7YtVLU9//G
sqK8yzQLF4k9TN6U3PTvdOsK4L9wv1kSWF+DGfst1h8KQskFf90rkXZoaac1jGYy
RQRnfA8wTuB5W/PXduVF7ekntRtoOSENMyl8CCFQ3hBdGTgx0/4UuJyiIUdNLTKO
Rg3uZqMDmEwng3nXBMQ8muH/dH21aNPZDNM4v5JckzbDbzGKsMO22nmw3HPZLJj6
g3JjHU2V2ZEt9rUnO3nY99JNcMznA+54CUalFtif3BkBjKwPqCAwECzrjj9AsFmJ
kCPOTNqWZcy8i+0C7jWDPvn0B9gOXMsnX4eNIy4HPBRshB4f20KK2+J1QaXSzHRR
QPjKk3A0R4UOkEdpH0J6coVbJ/U1cbzWMJVSTvoQSc8Ox4t01sFc7ybKGQX7pXFu
bfzi/B4YxjZamNipV20MwktjEGtvsu4aU6Jqiyguumkm0gLm3ftpjx+2eBU3cMee
ZJO210apk/I8tp2mHPvwkp/5VF6LXDLvG6YtMWAP3ek4H6VVRH2azoKbelN2BW0+
K1G2bw8YfFM8hzppkOYdqxDvxSprVeqmUKMGJJTrk1RpGKYUOH/j0WDV39BfQHGK
D/BhEoCLI+l2Nd5adbKifli7Hbg04aK/6ZGQfbIz0aEggSn8NYUvMclHK1M7WSuI
eQFnOKKdRzxEugJFbnS1NqNoNDpRZoES/BIdBPNcIH07BeKjdrXI9ZwXBew7Mh4M
ppJ/ucqraEcLsSIjB62mozjc4aKM95pcrHbuinVgvQgfhg3S4iADgTMMVJ4jB/HI
zTic0zccr4vicEKTFUVFu2Ft4cdxx+wK8sOP7CW/jxv0oB5Bq7j005BOy5WYjAw4
opZAwXGtjktXD5PY6jjxqOMkMe4s66y21HhibC2gUvnXk/Z5q9JopXxhOYi1LVv3
WjCdLIwYyRsbOZlywPnvpQICgHRHXjplpGcGyo+9PmSnIhqtlxLlD4kFW3ge2IJa
a61mT/fOBezv1aDV9MwCuMMRiPfZx7uoehBPTqRCPkNToeeGQAcunrjyTwTrrFJG
QtGJ408vnSAYr+7lYYUqL7TagxlXbH3ztsDNLJXxtkgEJFLInCE0lSrCvHwgtdtZ
Em/gEPqOCC2pXSt0yan9KqDBNBEWIYJ7sBgSgYtqlctvbL7uiacVAxpFHD1qLrg/
abQqJpd2RjYCrliz0C8BCRhD45aqV+J8VFpH8sJ5NUgCzOw7pEu+UhEuHxnpUSYf
5lsTGQO3CmIhKWCdY3+38slaCpZO41xYefG0gyeZxGYoNCgXnyyIL+qH2mywhZRC
wvRtVoIigEc2085Nf4XUZtdAv0UCqnlLD1/ICBMn22AWgYf+2b6uDlozkDM7NZ/9
mEqqV5MWI3fQGczc5sJ2oTrhEtyBN6wm0xYqfthQH/OCyfY/Ds2KCKkTVyjWOBgo
OoMPfxxMIxewpNY7N5V1nsMk/lwEoMHNaJe7dorujIMUHm1DJOxrVDZz3jhvqtqy
P3m20V8SHdHSyCOZwy4oAi10xASL3YmrHODdZjuHuM8znsvBiTKB8RvQ83Iao+XX
8//QTy0Mhd5vF58u3l06DXhMfGIT4VtfNERi9j64zKI+ekMCFCc1EPOyBmfKdRXk
MTibDpKu92r0H2MIa3jR5CMSkiwGsBQPb9ouwQzdOE1Sez/HWk2VPLGEHV8h76uX
8vjm7IQzBv4Ctlqqb4CqJdBChNsoKkiDqe7k8vHinEgVZsx2644GhPHzhRbIs9g1
6OfJ+v0s9rAVmROcTQto+UxeMjvrmCLbnULAo5ApB3cKefpqn4tFPJCnCQddLkeY
dBulwD2rsufna16gUk8vh1/ZM7QI5g4eH1KNbeHABtYvteR3EC2a3szCCRmI1auf
U4E6InfudbCH0rOlZCDQOlcw9v3CFVJyFjByWWUwERtH629se60pWfn6Y4g4jP8e
guj9QsP0lLZbwJTpB+S4GiGWYkw5grusDN8Zy/bjuo5NsqlLYl+ek1rSRNX5X9Gb
+RgEqo7gIFGvX2AgsK85KZIEZo4TgqvDaF4/s8tkbPHwb5HEGa3F+cinoYWAKjAu
5UG/TDykdDAdjIQYdVZevM02W5FEDyBAGru5QjHctKti7bsGQezCWks8Sk/Dgzp0
dP6JFueJHNfhJ0EQ2G56Jr9GjiQMF2ldo3O7GJDZbj7nhGo2cPshZfWQt78e3m7+
6REz+aGBFu4U7LRV747gPBNxlskCiIexc624S+LCQneNGhyTp53/iKeKr62X8vgf
vkwmwKU2j0d7chcfYHd+vfiZVwsdZesOr8/Xsqt1MPM5TeNi2o/e+fzA7jdpnlXY
o4Z1WryPVUhHaUHNeulVh6T5FkRAwWr5gkJhZarpfLx0TJXKruWi/uL8rSLtui85
lYMJpkewdIXqXW0ivP4dZuXnAjAKNMTeXLvDsCeTg2RthFNFxsf91fODw9knKFGr
yWkd/NTMi+rlJyUmKVfBwq5UluQaVW6gpSZQSWul5ijdsvYrryWDuPv4e3iI9/IX
yd8lCT7B0szXVuqOY12Hrqk4zdfYZmzTqx17hepmYW5oDsdYTTu5Gb9Em43YtxIK
k/0//5sBERy3TxfbURApNv1H7wVPK3pzDwMdoEkXmZe9W7AbnhUO4psVp1wndbUM
g6XbZgoiNIenuzdp9JUA4BWXoXlJJ1M9TQbO+kt+t5knyAnZsnySIMw2tHB5xYjV
e9WLi1/0eqqOALXWb9AxvzJHqOFyT+DcDt+CcMwh321V+bZvOSJRiP8BRzxt4iNq
vSyV7uU7wsMVX3pq4iR51kgvzCuwnU6KvHUGzPJisFuqCmwEI7DkXmagHpVtATsj
f+Zni7gggnQLBl6bnLJQd63qmBBdU6bu5maeI2OQTIzdbj3CeP0jElHkM9t/izh/
Cyffh8KAgCBEosAGlWvOxZ+dSnMl8Jj02WHfYIUCqFVyu/nQHtIbJxHG/L9HmSEF
GVhORJbVOsLAloaOHkow/5ni6o27lEigY0JaG6uivmWeMQyXq4thcWP2xsoifKDK
boLIGtbbzPIVtlyfJjyb2yCGUt1ZSBM8ZgQ7AvbdHVKOQ5RAPs3CRSGWqLvBPQtq
CxICM//RfG8wGenB7RaTt36hsx8XHpWJ5NQfYZbgo7lITKzmyN5PLripqm6RCBQx
BDBEmYslRDKngTEHTbEwhT6zLpa/ecZ0jatLSixIDuRfcSh9pGc202n9cCygdfuk
3F8zO7gZSTBLJJ03jLbstU+hUjyO7xyorrl10C3m2vbCedNTcLO5WeYKcC1T9cB+
wTeWmGMFQHORGPoluvsjHyR4wtGQVvqA0vpnovqEhLGELnWudrA+N0CkSGhU8jOw
4HkEY0zxcfEp5/ZUx7vTXeketJJokg/XRieK7eTQj4CPdW37sa6WbblMs4eJnZGh
urU0kLWVsvHgGxtIRiG+KZIRKPOhy+v1piVJFlAHqyeihOJkTIHwEBfz9EQvMjaM
3nhFETvZdUd0W9aZKsxkAPWid0QLmXQq3UE8q0yUy6kJTwVPrzAWbk/hQ7r3ukPS
7pg+vS/dt136wyuQFsjKa4lITBxkuuCpZyxfCw2LUEythKGb0i4Twc9L0N0bNXW2
WA0ayoQsn5nUbLRWbP2RqpyrvAeX9rX5xpIsJA6Ah2beGaTQ2vXpByK3KvwT//yo
iX6kKvCUkr3e+kBMRNKDLIOgcfo+gXoOtk4T45QCZ4WPBrEVnfN3RiJ4TQ0pqhzo
L0qvfpLNlWzTTDpuLjVWQTHx2K5ddcH/ZP1niMrotvGXUOvWSvGbV6HNSyGHlGuK
qLWk8a/zfGJOQ8om042ZwmZYkE0O8PacPOMbVjVzLfVchXnc2feSgRPmx8o43jKQ
kbP2XBAv+VL8HzJ/UlySBtf5Oa8aycvHx1t4OOWQ2JMNg0Y2uzBaKl61vbMsSZPy
0FGP2mmK84isljmCqJpCp+cZh+sDk5CHB2nYyhMsSHYrJU37eFmPABrR9qJ07Yku
NlsuFAwGe7f/YpY/IOsnZVhaU8cRngcmlnPRQZECEafR1bjMEb9goU80QZT8vuaX
SilYcBO72Qd3CpquVJZ04Su3tulDgm6uQKTVCaHuX4XdHB90KTsZNKg8b7ZRU6Ja
SNyVfdZRNY86WInQbZFP/VBYsnwTuSINDKSTf6UAbvxxLFCtNCM3HSIImF4HDGqo
IjF0NDsr0OPhZYSBVO1hwGyZDs53Ou1T9RGih5lVQBDvWXvQ/oWzVyUheXHeuI7k
Zz3k9BdRGjuDNd1aRrE9OXKcFXt3BSsaUPZs7Cxx6s97BijPgwlKVKzSBLMzTqTr
PIIoU5vrjLHqxt8etXM7YopufOPB4G0def8TuTURnSTASL0c08PLLFNkXwoPlz06
ybQGsUw4Abg6WlVQjb+5hexc0r8XaDf8nGmAq192nmRraLuzyQansjtqwy7Qf/5a
7pwIDSWjRJ3A4KMVo2R33ttRkfyyOhoZ1nuGnO9H48ANl39YbIP8I6m3lJHkfPcq
oWVs379maAfdGbGEn6Aodwk5l0sR6Cv23bGh6poL8GxJa2xfw0kIlIFL+A/NCqFf
rl34QcH/ZboYLXQdypjcUvvZWDXQDiuMCRIpR1/uL9xt3EfcGMZ5OKlKlUmv9pSj
gdBYNhLPAuyJcPO5fFr9SIvxLR4EmQBJAbhdO22wqcOPp1SO1VevijV4hcvua6vZ
Y9gmvttgLVV8xMviXpuonErOWMWL/AtgHvVNCGsqCSQhBw28BlFfyd2RkUkutO6C
fUXBVkgRy2/p+lVGbUjRuyyuK4ERe6vrp3am1priJFA3Oote2OFDLZecNL2sg/7n
iVKv4Zu6lN7+AsKtD7UhgBuZojx4WTFumpM7nsHxzcv8klvbfbjXthMVdFYHEX4k
asbIfGYvyxqx7ixIBBo08f84Ft88Qq/QgN1pDH9zDsx0L1+NRrbdRDKburG9sbs/
K7y+io3V7jcmgolFhSZYi+SUQPCURCVNM3sVLnzo3MsStG8KcB5QwzqgPkqzp/RQ
mE8fJF0uePlyxHcpwefNrvT3I307cG3o5L8XOpPruhVU2frBHTIQ6v35q2Ca38bV
riNBfuK3cccC9orNdZumnAjyxKTwfloUv6oMz8KSf87WIbEdapOKP7gmgmeFZlWu
D8m4dyDec5JrsckFQtSzfDFpr8MZdM3T8/+uRmZCDFafpfytHZtG0dZrwLvcImQe
QnTIUCxLUWaXAvQIjm4nbGaSRq7O7Y8fulYJL4RaL0Ct36AtdW+c5vJW6d1hJ+IX
s2T5y6ZaX8x7B9f2/tL/xzJR5+nBMOYnQnNC4HdwGzt/kCBl0txTmuGLdJ1vSCaa
IFOfiweuxMyBJoTHceIwLpgA0Ca1SJgjsQ1N2FzCC2ZYw/fjo0Ehc4D55wifxR6m
2jMQuJ0nLFPYCzpIDZgKNrUQPdhrNenyOKF4VNstj7jSbBtT6i/3I+GBrGu33lLh
VFzDzUtT8VOig2vvW49Lp0gP9TWEkGClMlcUGBKNUihtPD+ZdELC6NW4hOhzudND
tDKNcgjboxpIfFl3xrqDTu/qr2uQNkLP0bwQ3pdZ7832klz6SOaVoM1gj8shvv/Q
1K0eBDRhXK5NyRKmHMIBSCCN2Pa7H+HOPajPfE44gw4liKGCBReQOn5PbTsN1+jV
ejbcuLFg3WfnIuQznXAvk7eMU3E0Cy6ttYKAoF/QOpj9IX2m0IrHDgXtvD7f1HVu
/EzvgmkN1RhCFlbzR2jxqZmO+VaRXgTd4dWTAuWjz0KvozjLviE5+lZoF8IbmGN6
H3RhctuWc2/jEMcBEsM/+r8C1Nko0PkMVfS4Ez/3paObuIebAPI6S2zAYyZq61Ug
CwXjSG8gzQuNawZ5rds3o6yBjFz98yW7lKwNaxtSLCxtJ/KspbWKDuFepMamgI17
JFPcz6r6sRbr+P5eDD/YqUfnKnXNNNtfB75s2q3/KhaSWG2qnxIiGxMePlfcaAHH
MCAzOZHqDp8pdHnXKA+AVEquaf9AGcITF1etvl+HBU17cQaTTRn9PVO4BEGunNhc
Nps3VFnvAJdbbOxCNBkUILyAaVvXUhbjSt69gquATGcS0wZsOhXfMGmVGZ8FQUDF
cZtQnkDLl738rwzEYDOeeucrKQXzWoRyw80HyZahrYVeszFlxPAhPCbbIhAQ65nS
m1MOvoeKInwefsA8vcQNzudZIQZCEYaEVaVtkbw0G4jpdPXQeMqI9QxxLPaYmvXu
tCrMZ81WYgEfR8x+HJgeNTPasOnrSXljk5AMqz1QsCbBWfcE4LkbWbWMhzQknz5/
s5Z8pVwHdaeD8UJIA34BtvzN0ydQahPpyO4fdEQYIrF/sjTFCUgDZTDOmazwtRvH
1+y4x8ak+8YTop7vrtoHq19ihJuQoS/4MVBXZEBxafXzUvWzA0StZBSopYJVqQAL
neojp4ojU9zAtzo0GDzIEBrUcaHKOL3OZAr4XRmH5rp5nTupdlitu6LX38dibYgM
FQJSbbxFinMQjpxUG4N/MD+8yNUPqhiAYJaAL0PUQ4+SM+w2j6xwqncmW02/cAZf
5Ef6cSPqHxxtsZ8lduwnTSQWzGIGCW719rBDmg5VlbNe3D9E39vkc4xHaJwS/sxl
EemZjWWeftfNBlosuIBr6gAK5Uf7og9fJ3Ul+CmsMuXqKDTpSBDm6vEBWpDkRudA
SRWyY+i7e11fVjXyh3vKTVJMuFcqPysjZxDiIngtIKZl1Abq+Nl9dwj/0sQLUEiM
kBfGrCCELixr1jE/NqSA0lixKq3RIrlHXptUmMR2pddH7m9Y/1bRd1zBXa2sVyeQ
McRqTg0Azyo/UpJyhCWH/5yAGYN6cj2zKVlSnovvqngKyWjDjQeyclpdKjg6N5dx
KF4HBqclEjaK9YqqHllt8xTuYW7aIo8gxFcLjUNoiulS/qVPFtlwtaLSaMhaonnH
CLqIgwcKW2jjPaO4CIBJGCGoYGjvpECcOCjezhpKhvtOcd5IKAKh9cEedNVED9QU
Ihzz1NqF/YTmnG8q7XXyBxOEsyIXO1oqHlK1UP1+F9ZyJb6NJLCKRCD3Z3nfvrd7
uMhW+Oc7xt64YN/9dLTtQ2dKL27/BiIPtMnzdrVwiRW0GdG9qvhAuTBa757fX8IY
ulIjTAbxma/6G4gByEQiBoXTPFloKbyGzBZA7FAjm0xX4Ez9Y4iD2ieY72gwORTs
W7TSnYnzaC4yFsFHXGvsJYgG66jU4f/g3eH1daeKku0bawS8+Owdr5E9t+tnOJc1
sr7xRx8yqnAoTJPkKFYTXLxV8t0nDSwhQkTnsU7eoy79qLs/ATiGmSwb2AXYSCbZ
T2yYATkgNeWPbl9wSwQHpJK8pL3zXLmHm12HwX5WsArjqIaGVCH76fEI23SiPNfP
ItcT7XITHtfuOB/xou63rjKXlAFHrs28rMSNpsp3RnCqfW+7tV6XwWrlgoe+4pzu
HELkDqYVXIFFdvYXSTofT1T0d8sXhIk6hiTKw+qqoj60vRMH7rx9xwBFfluBJjZu
PdWoOT+4w/G72aSvK6n+hjo6Fq2+HjEXuSZZGCQd6cJamtvJ1Pt10wKfhvWsBPpH
lMaNzEpVpvYrhAfLitvr4b3FHsUS+wHi1byT90xZd58BOx3HY9jaIw+ab+GjQVjr
V1TozGr9Jz5JqmkL1hUUaNlJxlFzM9eZ84wEYw7TpBY9M7++dOCUktP0y2MeGyzv
gB+eBtmfkB5mCIX6aO7xWtfNQ9ZGWe/yaBxeFgOSuB6NwM8VGld/lawV2PKf3ink
f25ra3errBRbSieWDM8Ad6rCMbsLg+tNcbt5WXnC1gGI/oomQbPNNaubcNOw6LuA
zPSzdMVyovIc6dYpw181rFaMJxsC2K5Zk8P1ms6uBa0fHZbMCcCO61kJdBGpWQge
i82lJiB1t7OPvm1jQFNoio0dHH8mCJN0Fe1SKb00rjFSnoPku4IyArTwk9stiqWp
tyK8+h8D9GwT3pdfCSy6iobQqDVEV58tNbPkUcGyKR3uGVu/t6MTMJz2Z8R3SBl/
sv419uJYPRmoY6m2Xt2LZukN1F2bu4ZmsiLnVIF9TQgkP3xUeO8Zx0F1pK/Tr9FH
iPvueO3OjnioWw6P9767qHFpD6pbyb0cVwDEMqOwC/sx0gjtvB+qzPbfwOtBMbZY
XTtZ1iCK1qsjRxx6zB9UdqsSH0Ixgm9rQD9oYcWDg1la5MMux4+Zf1co42UmOADC
VkTmQFJvl2HXpzxBr3vF9yxsFIh4qqw3OZ2wjVfvzH3ZJnesirjWWuxdK9uvxuaD
t9qPjYjQ52IUxRRgcZ9hqElLoPO5Z1RhpVGvasrNQFie2BbbA6fPJYi3HNjCSZPK
Jor/447OVc6iR/LHRw0dKCEmHAUUefTqwUt3QTcNjMhMFDiv+vikWclsTr8CeACt
TyZBowaDJjuFd5/XRnwIfXY0B6icRR5AwxbZhFQTwSsCPKMTKi1GUEhQA6wYHVna
HXT0cXrDXkHvhAmMOdha4PTrJeV0zZac9g/DFDmre4NlPW6quJZ69af+ub8uUnGC
B6eSm4WuM6dWC5kE+9ARaC2pgOMm6scxtadY4QVNXYRG0yj50R2UezkdQpfARI6N
ZyVcuRKycwpNe7f1Y++qdWG1jBsh7mzglHtGQ3BIf1M1ODgdX8etKz54MfnanYvz
OpoeIGaCG2+v6YS8/vJNcVnFaoMO5bwj7+n8ofxv4DjIuagcoG7aA2gbkkB1MGBh
DjuHlZkZZ5TbynHnuTCJCwS25dMi7EurHx1erd9yGoR610cFLBfxd5VGHC7tkzrU
0pRiVeGaeUB94ETm7Z5eE2nDOrj2zpBUfRc1yVvqs/4yDeMCww5NAqLxpIodHVJQ
Uc8EwtmCuzKJkxM9W0KablOrvL+VxoGe4gYZaW2jzpeY0E68nXZ7bpDOMZGHYztO
P8Dt+cFYmNqwEJ9gJNvnrIbKRO6mh+WHEBkGdYFCUD/vUCuI3YlS3ovZGoOMr76o
4L/et0gk/rgznfo/6Ep8dn/dsIqJq4gPxwBRS2SA2yVbSkGy2uMr47GPHPO28bPU
RyapirYPhKqHhP7Vez5fVUHBLEx/NGBpBUB5tumD8cMAqy3JHaxYYVBt8qqlCHMJ
UlIsJQQD8Iw/Mfxz++DntwmSOJQ/pLhIkYaOSeqaL1hlvphZ699BEYv04luK5lxP
EhPxROgn/alZI8CgPvo1AXnRgyjM/IfRpr3yP4w3B7w63j/Jc9OGsXl6hbxdAiVP
NzkFCNF02kZyQoXwo3zseZ6U0sQ/Y1XxeEomb84s/fABSabsG5IVRVshbiW83fYZ
P1x7dl+ap1IP/DIXwrgBmQipWX4G60LomYeLJVxhBgnAgKpFDAA3G7SJbkIWvsWy
V4zN9M5cnZm3WuMlBc4MwHPw31FpbeP/7cqAqvRk3dXhFineokDJcA1BhCrgDINH
pB0bJzp8V7KHmeZMjXhrX6WZ3u3GMwmPcS3LRtXNTxmBfDRYSxNXeuuUa8Pss4Ji
gBtMHiF/U6pevsUoVrbaM8S854nlr896vr5x9KQW2tRKkXX+mDAlKCPvmHFbEQmm
OS1bc/bE/KEIUdrIgVud7/7A4Tf8EycjLXeqHDgiftjy9NbNVHnWxdVn8zuFShOb
U52LP5LpLtpfB7qliUt3U4QNjJiCk0JQqzIhCDgvrf7NDKFgbCWxDieiK82KCtQ9
XkoxbusraBEbk6SdrIxgPJQ2QyXMr6sQzg4xPh6YvPYb7QzWGeKJGDUEx0OXcFu+
jx8oG2U/uO+SzchHrvb2R2YLlOhbXFIa/R0pIS31nD+hmvf/zkP4L6haDMCL+gmC
h0YvB6OFbXJ+dKqCkm9vUiEkW8MSnX1hEpmKL1QbCVUHBamdm5XFvQYllW36smfV
MRHeXaL7qqzO7aNJ+Fdup77bo5G4FGyyzgTkMRLk/IbobZ04Q8nNfmr6yMDj57cS
Z4VZMMBs4/UhDWPQs01pw3+aRy8bLOFaT3Gv8gqQm1LF+FdiBy9iOlW0TVTppag0
bkemqJBBE4/JeQj7pp2dsGnlvGUWMVmZrs4TojFCICdo2qsHXtg3jIne5RHApxr5
+7mGlLxQGJOVosWG5byVtnw2l4XVLVzH6FE0qRUI+KgipE1A62+nARv3BZ5o7T5o
QexuDstg6qqu35fRaj3nmZglyW1ZfsGwdAio76oUT2eZnv8+OYONO2CwoB18NDwI
b9j3dcotjKnlLX4BP+hUzIv0umZjfyonR6f9UoMpll6y7YFZ61STl3G1+DyUvtyO
K/XOsisd6LoaKlBcXkjYU9X9mDj89IkT179v78PXT3iFbcilTB2lSSsCmP5e9qXv
tVgcsAJQMqg5SJmB4O1jZah4lXZLY1duEtgI9EMlVhPXgYcW3M74WS+ijbZh/7Kb
W+DPR6416GOK8rTpsDAhST4pc+uTskyz3pk+J8Cb8/WoUoeTyedByR0X3TLq2y/H
TWlydUSkiSNoGDI8FEGVQArn8XzuTQvim6L4VNA7fXy3HiCk0aMZXvv2C/ngMRG7
5NK6SGAJQRB4sD539qOl5kQ5qs35XzBL6zj/xlmD9goowVoxJjiERiFdjDbUCfc7
3Plia2JPW1Ya+u+P3hi7+2foJs673V5/gFR0kk8Ayzney/24TlB/Wts1BnmrwsWy
iwbi0I9uRXgxaQaIRU/RiW2jbVmzMUIlZCG0fNKDxNNTydo7aee4OfNPhuLFWLbZ
Juk1KlAUKPrqSXGRIl7JdF/ddRdqDFuGAGEwskOocKwqENc3qYSkK54v5iugoWFI
EQbJ7o9ltpL6+NmhEXLY62HnCKRRFUAbyKmVxhJmzp+OQuMaAAbSGL+o+yiZOh8J
81dMYxaXDvOSown16Ob+1ZE/7I9GsofEsrZEUAh3//7PFyax7IqOvr0SEx694GMD
nw6vMw18VX569lyX5Mzqt5+I36Yu6PeRJ53MIY2F2K/k7Nn8u0kfd2dktH41UdMD
qe5sxBpKc+rPT43vgrHpZnABBMMhebK1o9IC5vJZofWveNWva6g87PJxbiFPTfJ3
iJ+BaFouFq3HJBNMmxBJ4J8InE3hPWowIXzqZWIRKrjvFg7wVjjSjq+t8Tcvfq66
KfshBcrlAWbOf6bKm5VZ2j5JF0z0VjIaZ8wvV/9k+2oHj6Pm+qYJIdfFZepv0+Iu
QtC7pMz8HeXYywUvAei4Epa3pqaNsDMOuzuzBIrDp1zN3LJadKwHheDpdTRb4Ppp
/9YhvL2QqtDnbXKjXYdlOmwIUZI7YkvLQcb1Ra8hTF650x/atoXEQYrwOD1pp4Nw
xxNdp2uPMsUJl+rLV6jviNam9fmiV9ojUbDGpoYqoSX7cgNaeQMiHa8qmmK2UMPW
VjBEu68tI6szmYi4ynWwMU6khTVVEXvbPFfIlylbxLneKOmNcYXlWk9PQJUP01rg
Gfrq4Ovm5Pdfq7Q4xePRWlA1H0/2RL4glhg955Ecoe8dFxZ8ZWNS5m7LrF5tfDb9
k36xcgR32EfyJShw7iVkk9IYLOA4Mtg3LJFqwlEiygDQcL1uTM+3yDUmdJl2BO9J
+3y/GblthfwJ+DqLwbq2vd305Xv5fTh2duk+fHOMgrhgSC25kl5d9MBtZ2hr+cKa
5jtSq8vHHdvWYucCmZfMrKr7IvEBS99C5I0Kf1a2U0TOKfZ76TJVvo+uXta+MF5v
FMRov5vTy8STVEsQNorH/499pSdyC3JWe56fpCgh0JzyHAlfds47wIBXuN/ikjf8
SE2V+Rx/IcVZaGYM0bbWrq6AnXy8Ive/Kp5IS7fNcjADKNShS/69uCi6B0XULHK9
xc9VwpMtZ/iPyxmfSiZxH5qPSbGeGAId/HNLCaHrK9VZMmoAe/VkfjXUgaK5o0hJ
d9g5Kl8+QErYdqbqEWGd05dsWxZbIBRsCMNGn+U2ZymMVn0Vgu2g04JFoVyLuC+R
Xjhc3nMpXSFCxzhPt11bp5G1+E2IWsYZkhRtmGzzkhBrEg9PD/eb7t0F+zUxj+wt
ibVl8EowiwMudNFneKnKmS9DQMQWphXrFd1zdrBlVaHJR9m771++GcEu9zUXmgF8
S8uVXzC4w+bNFerul3/Fg2aUUah7tsjSG2uVIx6uCOHJs5pGIZUgZqwNaVSExsWt
ho6NkwPIV2GkjaZwsafLrjeJ7gxh7KWyu3TYnYIAKY2LzMynni4kTnKR4yxx0yhf
eGMnAfa1ZKMLzZ7kQI+uxGdTI0ik88OKCHmfE+jQXgYeWfCK1antV88N3ZN+PcK8
H3cqlvqCoKZTjqxOxSQM5QnO0uJgBYLURN9mHV8hIljIOLLAYpVFjtQRwFOgHr+1
ZTe644bGyxL/Pf68qLFZaFWKQxD4f0Hgyulu4SZn299rmInGCEYxFhWBt2euhj7t
OZAwp1dLifhfjnA5OjKZhE/9apZol/qyFg9jUDoSVHc2BTN8PfF5BmYcPvxhNBUa
5O9/oa/dVE+R4P2MQmdYpmsHP2SECJ3BYnXpFJknYdiX1vx06377GIfUzr83MgE+
2fbvimH9RuUGXGTQW39xvMDHfQi0vbK4qqUB99GHu9LbeAtXJXG+0vDqyKFtl+Jm
Asa9WR1Z6OcK1QQN3Mm8/j8jlcIgzDNj2z96OERkBcMyzDy99E/5NhyOQGC5mb6K
04xJVWPQ1yHR95us4orB18txq4vsr+2T+/LltsZ4KvgTSZaBQ0UPptwoSsMvobVm
VsOxqP5eZDOV7ozLz7860iWd/GANR7G8/PqqKOzMrsdUe3PJVyfmLAy38zxDj/tD
ThMkx0SOzp8Sp0hlNuPlYJdLXA4rPmX9ZCZMJlJj4rwoA/WjUcYh7La7j1B9xh+8
gEYVmz1vvj7Lw+OagreeQwkNR0h8cTlGTmXlrXvePo8BCpgbuCyv6CrAvZAXVVz9
z7NanCV4sJdOCM+Av37AGZD0Tofjocu1+kAYwvdATk8cIJPSU3yTjPnHbfDhl9ce
0ZdaDZum5ZJck99PmTKl3k3o3Yxc54jwD7gOarmq4/RUIkxKNAuQ2otyG2TrtCdE
CB4mDJq1YQzksbeSx6sKCJRdhh8ZiQftJIvj87sfXdOjHvG5jCkcpbhqStnwVZsV
4QniMdmbELkPNbrk8IR3hEBRN3ILUOErhb1sMsVUeVfve7mm+dyAULtXaLFJVEQV
1Oq5SKLjqI0MUyU4DfBpQueU/23z3TyX1NUmdR+g8tHWQniDwoHGFTGBCTYKXS60
T1/WrMQaz6cFLRumwMYY0P5UzqidkCZ3j0/cUOzJqB/9NKGFEUhJrzJf1TIA/V1F
Ug4/+CDBpfDfuoPz9MsIHy0GDveTPlcZqmcGrkcXW3aWfOrOJBD5hJMuB/TwR26A
BIyGxQNYTM/346JVsG5Oiam+yoIiYqALlv9V3hUkNZnGjrAHbV0lQKy0+og33G9m
sYXzD3QrbXkoB4U1KKdQt15cXE70sv0mdPv0zihM74FkCaQxoAiqjpUHWNTFgPYb
Y+8aczAXn5DJ6EoMLKxdLgxn1jwrD1S6Lkz8840GhTp43yKGgJgHtNkjRixbTIK4
dUu7Ho2q3q6fuZiqSYr2xzWHos6HGpf8MP1vVKCH0kyKR4D1e9pZsRrvSTUuMmtY
tlhUvhvDmfaSsDbbvBGBO1/laZZlm7BIhXnk6pH5IEX2nMdllmhVS70xTJcbydEK
TG/8rFqXW2foNJ1hPjZXKooBdBjHv982/EPqjyO9CRzni9ZxSmJziIjenfNxUTNZ
+kYc+FPFeMTw4FHfCxIJ6836n1OAgQCTU9AxPohotuzGlzKMXmGQQkQq4wSe1e4+
U6ujhyDvBIFA0SSvRDOfsqzP2TIU0Mq3Xh2Oj+krcEndfWYRSOKF3e+44P7K8Nh6
47ODgll69NnaP7+SDey8dJDho2rI7pIM4QtLpT50LtM3j4/1JVkRPnfqGnAhtUbj
icyz/jFlq7qQuPUxiLT3n6uZc68a4efwdQO0DOXSQmikNbR9GJUwa13paRvaakN/
VxI/99FNH17hVTwb6AJQw0DPw13NOVp6aSvz89pqOA5Fhc6eUVr5Or6qIf1C/oFm
EoZtS2TGTRJ54YANq2x6b4kZhIQwpl7izYOF1HLMX5Afq1pfBtRyAdlybhi5A2DQ
+Iqw/hKrsFFhljfOXbsCzJO+EvpKTsU4ezCza2NftVv0SSK43Yi/KFrj81Qe02ZX
eryxHaQ/AfnpqDPPYRj9NfBnFhAddJV5LlDcxKg9m1NV0SuX+/86uWxIJ/QDiu1r
V6pZbQsAtdTXoNdcYVItkidkd9mFTEKXPh6OAfeEbLo4kDVCejGEU+7TSxH2d+lc
nSyB7cOPdUZxh05jXjd/m+W4Z9oYkHHHhK/7/NwVIlMMxiKclE2dNw6KrHi5IzzT
dgczvD/Vo9ViMn+NXsPhBHNuJucwN2kZbKyJ5r8gN/9k2lzmz1cQk8tVCLAzdiUu
z6jRLIQ6goftvXXdAHJujCxmkq/w7bchVzrq/U33xeznVcI/QmIsDRgoaqZPNe38
YCRuMqtV1b6qwe1ZvAY79ol87ZzJMZlclCLIAy/qgMEYPJIDvVVV728BKgePNK5v
cmctdgfpjVEXgKFacc9aYgM9XWVj2UE4Wye7K9/NxJdDlpwBTjZ98CQU654aDj44
ioUeoTeEEbN1rtPGOkCub0xdCoegR5fk2VaLReZL+ecqCvqXF0ZW7F2PBwJRXPls
rcTUQXvq96VDzQ3AIqrPBFr3iModkn79dpgP9p2PbZZ4+GkUTjdhsdq0f8zhqbqW
LcUZIQKQO1F+0bFhnFjlWcZDvckTybm8TcNABItM9PXT1Gy+WL2/SDpD/idPw7PE
d+2tNms0dNlLqoqpPP66L1VLcOhyGgBJj8oMbyOvqaxSF9P3r/7G8JBLIUQHJJsK
UUKGkGLGTEZ3KP2FlU99ZP36Cn10PGwMDPT78AtPz3Ixy1Mni+qZnQ6RxhXn1ccQ
SOBc0QHkVzfIlxF54bN5LZ76OpAfWwWq3PFY5iMF2YiLKQWFZVfzqKR/9KsLaOR5
Qo4iIAIOsPCy8kuH6reOrG5aK7/9+m2eNr+nu/T6TlNqYfSnnigrkWa8zY1+fCxG
sjWDbGkChq5PEGg9dZcAUn5AG9ZtKRY0QFtqrlEpOlYT6m1zngAFUcWAo+33u5da
QMORga8swqskjyjarLwx+KAjKIacQDDGqZ+1AbYczNAs6WEAXKkU8K8nSBhxoZCX
Y46/MiyFcYJ2wJ/hyVpj/DjDAzeqDo1mVOVcnfDXsfgFFVmhL0TdOChPKt0hjHjs
lLh0ZkS+2KmJluzcjQ5vO396Ou6BliSaibnmq3auDwttfDPCSiCOHlhhcT7s5mb5
5uS3gTImTgYGj8oCJfhuU7+uByZHL0VY4B7yXzU++jE2zQJgw+hs8gggOo+U5hVm
+ZcFlm6YQ723gQSeU7hZ3m9PoSL1qqRCgnlExOyenyRbdNFRcMD5zrf8vQmYl/95
4lPduP2Acc6J+xLIKKbsQoNDDlzuhmJDI1wAuBnc5JS9PvoZ63e7m/Jv9numdlSW
lgMRQYqNlk/zbpddGepfxSx/TDLA6jTqutYaH879w3grzBz4gSwEcFb+GrR5bA38
NOP255aDfoaOGRS3rkNyDofOu0Rc/o5WGKTmDgP6BY0z4reygiG24NzBSUJ3FkRT
609+Y0rqLVuVY0WYx5uAfJNtjAKwLlVfmDV6csh4OpUcOpqgWD3FuYxd84WXiUbY
pkEBEINzxecgA8pODal+saKNt2x3QLqpWHXZ6zMVt+tAMwDNFTK/F/VemPYG/V3z
mg+eA4m4/QO7r4t5ePJx17LJ3Nv0iibPJIovidNvebFKls53xMXXtgl1+X9Q48nK
Xw/BAQiFzwC33PB5drLBJWtrzj76pEb5GTdbY+a9b2QBzXVcUjp4z+hwLpCYGJgN
uJSkOt6IeRMm50lFO3fkZbJ7t8xyModvSL+J+e9nNmJKshW3/7tPocJQDwB0V7P6
ya20TgpA3FZTwqDN+34QIUwQLTgn+3DsCoGqGqMcU1/MhEQo51gN095IT9DxGEOK
cecvVDdrQieRLZR2VO+UETekEU1fNsoagnsZN0MMPHee8hRYBzFeZXoEzdrFxjHO
dNrTDBTBAbWiAyyO2jvj/S02peIhp5vUDbvDG9nafp5pZGf9pxQe6BaJfDJYMpHt
qu+DpPrb5xljGhxWV/QHSVdflH1UZrd2KZ9d/1onHkdVAPTEPfepLUd97e5WzfU8
tOPLmdTiB9coOu4mHZpHYZL8asr3KVHI+QduSibGq+5EhgdMjAJsW6sSYVWyJHIp
AxPLRjz7AZYdn/y4sxEwQXj6AZpepWoaF3b8+912rJjjbZnSe3JyaXO9Jlyq9jEZ
TNijcZMdlmeMkPaAN4mK2SCHY0FnnF4pZ1BW7jNWSypfAs+d14l5ll6IMTDjVsWR
ihlXveRoHuk2z6dh+NqLQ88FUi9IFcsTpNNH1fKY68YsW41D8pIzgQIwJQbe5j5P
yXonFStCm7TNTlk5HLm/6lLxzH4iEjNRNS9SuW7CyZPb2M5bOYK/Z/RiS5R391ZI
IQUaZDTDhLJX0NurD0pm84TeRIrU1jVgnfl2pKxIDH+UmOXmKGLd7qXaVsMX8l6I
ldeC3/a8qkU+RxHkTyDxYmN4p4z1/JpjXN2pS4DOSQGGxDDCpt56aWem+7C3ZLxx
BjzJWM6f9T8w41UB9i6EkdGgDpDCe2iBFvRzFaUrSucIJ2WpqUdUaR6Zf1f6LZ+A
/D348unxPc3T9hGAzmtvpJGuWtJL4kpeBfTHBE02K8/i5grXx4aAwM0D5wCeF3X/
NOPMCWiDrEImSzgYRpvRGc0VxEAifjfoDW+FuDGbCGMHo8IrdQO6xaMKc8h1Yd3g
vjvZldeGY/DQUqvj9p1yg3qRID8VRdWYxXvUMch5FzupvHfZE/ynC+wivju3B+0h
834LofIQVfU+YGm08Cix+PmorcF5eAGPVOhn2PtwWP5js3IooMjgPLXUzmEQ4QTk
BW1GXR2TtcAR/qXE18H/TU6Kqxcn919I30egh5Wu0wEb9hnRrmEVSHqpLd+ARBLJ
FlGehqkCdhIrycDvzic5icOZ8vp8X6sD/ZiQD0ona1bsI3uH0LVIHLqMAhxuuag+
1lCmhRvGNC1rwQbiXCmOSptShMFAwBmwH4Y4vljvUOiSSpffSPWVqxUouZ5IaU1Q
bBVS72rjuv3Nb2100WzyMm+y1IzmBa+ckh0DuGbTGiURTNaLJS/HW8tGWVSqf2xr
XdeIHiCoev4ePaBIld5wgFMaZtsmmZhz5wXFd3z2SWsmllHowxeiKegktNubnI4p
wbdWEYzhZ5NIVZwcmd00lEBhz/vd6r15Z7wMMnqRpqiArtb00o4RojCZtFD42BkU
gAmo2sh57j1R55GEdxKWNfHgFpN56QJn2mmaa1ayxHl0aHrA2JYU4Sxwi6SvFh+X
89s11lm8sKogFegr8mXU7eKqNuXpoeFP5TUPIq38fBSjMSxL5zL0bUxAldTjxCfL
V/BYjLUveIvtTBL+by/MqFBisBtBIiR3EvclZ/2tiP3gSNnbgvrHQAePCHBPGey0
U+p9COnAHv0LIPOg5z2rtGcyGxQSxyUE4mkDUsYujBUnz609XIldG3QWtByQzhQ3
supsrMQ5cbSEcdQR+kzGLzloG8CqycIWbLhjcxqo1iaeRTKtu62bIu9MA61p/j5D
AYtz+fa+RjNfjyjo5nuqDJQYoYcm5boCtLH1sBnD57rkCgtxuvv75jKmNLD+MCWr
NRgjWUHAenzGc4NXiIMwADb57O92NA+H2tVUHfKySbe2JpVB99tGdFqAEQOCNVSh
CfZ5XW+igIHeO1d6g39iTLKU0kZtv3mw8nYS1ezV8ZrGBoVDAX0KDQGybQbXvVqD
fTwSf5YQIw3CAT3msO8ZZK+3CG1kV8bTrdxYjfIs0x86L4bOyPfhlass1W2ZSAH+
MBaxyDIumllh0JsoqmRRvcBDOMx3lWBaqf76lrlLsbj0SUiLCAioRPprWXJLcklI
UmTbudeDfITDcJRcGTbNJL/bUae1aWJLFnCtG+R7K9UjLWeSWzmGKEX34s/HBpvK
C1U40SQSduwM0fCuGDUpSipFzS3RXcxQ+KXw6S4xjnplhXHxBV/WSW49ubuowRlc
mCHdgZflPXaeNSXowm42LV7DsrtuqPdwNGAo+5MeWspiaqMj9y0O3eSq4pp8ngn/
8CUWs0mL/C7r9CrB5fdMaUydKIiqsCVv+MCQeIcEf2XaNkHUaJ2K0Vmdj6HdUXgA
OCQYRDe0cvTWve74uIMPoJtIDCL8KPuvpUOHN3hMp726oO/4Kodena62R/mb6FE7
COaJgU6YU0dlmsgl2uYYZWy2wN4uy4TtrFsDvGDZX32cuQRr0sOC+SzhS5+eUwfv
QXMOkEDyCXtetUhEAUmObywQqsQKWweAOzop18IJb7yIKxqU/0KHyj6LRFvdVTMR
YqyRgJUawR9cVevfUDWCcRjucMq9khuMeYvIoBu2ZHagCnD8/Wd0qd0B0A9g94wE
aqjifo6t/6n48ksBTWuVyNBbDyJKdafUGNT+KZ40tAxrvyKB2FWctmleavLSD039
IOhAkbUVJ/U3B6vmpK5Z99L1fGkt5Go9NVCQOIrOmlNcNTBMLqNupf0U80ReEOXl
wXdJOadM1qCPAcgjdR9JJo+PbpimWIhYz2bxMoC3ILwzG13POwohZySrRMRiBrqc
XSpPkjEaAS87u5YKZFsnOEkNMs7b01GLj+GODftoQZUbhsIIqNYbpAwjLa0zDxid
fmDAC/EYI6m0iu6C76QlhjxPU4ZhFoEKkngc2bc0XZ3WmS4MVOjCFrKSXqok6iHq
VtiNZc8yj8REZP4evbJ93afARUkdmNnluE+PiSYjHmdOBCi1x8E5m9AKTElLREzP
4ZPLg/eb5cNc3iK0o0/MrHqwftKmBgb617T7LWtKI102dUfQ5NHStFlGLYRVx//l
CloR8sSp105crKEl0TZI04KZ2rSvSLf8psWX0tOo2YZioxz3FPeHDhg4RgSpcasX
s3+gn424TgfTkkKhQ3ihVeToiZL86cSL0zHtnDJE/TOgm6nEHb3spcExoaBFCwAI
T0bJWcNrWOmA7kRISdw+PmvzAlhiX1Ox30EZqzF5ptcJjLCE5a9h+5dqJPcbwd8p
LRog9aZ67mErNkcojiJKy1DyGKCAww2WmUnVBz/19bn7LlPPYLjMyX8WPeiqwiBC
4dNymH1nME3Q3CGbgEvn0veuZeZijdQx6gIaGDAZunYohRlR5LksOrKoZ6UZL/en
1i04j0Ap3xHogh1UaUmEimGHeDKqrY0OqTaAj7C9JlV1drUgVJLyDW+AbGybB6Jx
d0xlNdO+uFU4lxrRyuM5XdtJw2oHA0dln8AyIJsiQWUXGNyTCcnruxVhEiDjwtZ3
YMfgXxkKOMitujBW+9mey5DkKcYtrm7B0iynNDZqrA0bRhfu/yzdWpumKQqU0C0z
6yHnmbSj9fYz0Pbe1VplUa5fUCUjGvzJe3DgJjU6Glv5mRfsmZ3cvt7cz0Jlansx
HqdD5EvFOMKME0jD3wu8wcoWUGHNj8gx6rqEEUmLYDZCqGGOdgvzJgKntFc+s1xA
Tular7+a3PKxWyv3VTffW0EnEVrNo4zh4Xvxiw+jCryvriL2RKC8Q7SrJ8ynLS8Q
IUQTaZIAcx6FeHoEioaP3VkuIXs8Xo5xlfMS0h748qjq1fJmDYaIawd5pRbEyY0T
Fdnj2In9TZ5g+q7d0KtxcBuLiJWGkFtesVq+vN9+xG6429LQAEqUA8KZXzAlrMla
RGsPodn6ikewU9clF3jJbMUwFCwzwat6FqQTtKQrWBoiNEd896d5xXLxkluDGTRT
MkWWzaKl5W7sEMlTNofZJNP5k2DXqkFO0V2t6VG1OUnuaDivulKS7GGi6c2+7skW
pWTlav5qyUcDcA8UJ1OZn8KEvtmFGCXl+tDL3Vh/A3tw7OMzNGP2eq7gBqVxha5H
hl17raZbuoEp2hXGx2sf4p2sc9BOjmbP0fS5XMFklCvYJ2Mw7CoYvYK+dAAioPFM
5TxPvuLMJEwOMrbFCHwMm3PdaeIMIl89wEQbUwQyUXAvB5X7ij04QbAHVt+8oosT
KZndW85D/Atrd8Ekm3I/Px6TAHn4Qk6VyrW2FTF/hO22jq7FYNKHS8jpHLFDPqWh
OAbVfNmXotRh46xuUDbFs7XiJa1Sbg2Aee8P3aPDCBiyLsmLzP1AHLekVeXPW5Zx
6L1jGfPe02v5Zh1TRFJsQxdg3nMrtl1Vdk6KXPt5+KmJDMYba5b/1Pz2t6pIFBew
W/vVkaBKKL5lE+KZ/f+PHGA1uAj7/dHrIg0APbCzSuNzFCHKLF7s9TVD6OONAHUb
5PTbwQhbcJUYDUbmpt6zDD3VWWquOVxhNfPiIdsMprvxsVgOPizQrZ0ciqKxpOEs
7mX0GwBPye+GsILcCPI07TKv8v8zgDqb/rQmawC5awCejNjhmff6JrUecckBz+09
Z6GR6zgCmwmObLoxyPtr0hCFaDImdLUIRQU+iQ/slMXlfL1g2HoBhU2OttjU49eX
7bwStziheIhD6+wo/X/sfWKbyIQL/IIWyJRYtAZKhaCfpVAO2v92GFuTBsBOlIZ8
0mTg+mvpCFrzaq+DeuhLo2IszEoqDDKx3D6KVBgyRM19h0uYySCVYl9VgHeRjdBi
ItT+mYWFlxvn/7+uTzqYo1mTk4+MCCdey1wSmDtG3D5D0wbdcX6Zb/unNgEnEg7J
75yzhlc/cUMRa/T1YF5pQqDC3XCVhPr9A/aFJiuqDlcG1RTxF5B8QOf5nPF1GbNU
BTGV80CJQpS/psTQ9xdEnCZhgnpRzFugWjjNMGV+j1SaEjs5k8XgBaDpkZ6yG3tF
Jm09zfONQ3dZXsiqTPE1ZxZr0VsgK5OR/mZi1/rBAxTcOe7SmZc76gsa966vVSm8
WgPSr/0bK9IpE0tDMD1rO9ijXr8AIWCGCfZOmr3RBZ/N0vV9AAy5kgxZTqHqaVbq
LDmKIV55CROHEPBT8iI2LrwFyBaPHrz4QohwPyaqKPGYZcEds82kssVroT03mg4E
Vws2yXcTnYGjvhiEa3ohUVVDJBa7udlAdB0OWHh6Nur6+gzvgVqPKaUHUX2iXKf2
Jg77lk9Cqz09GLNNqcAWYc56qyy4GUOToClxBC6jeeC1PA5fRUocCd+Ax2itYLDG
WDg/++nUqNi4TbvmIbSgoo6ibgYjF0jwx6pnzh61w4szkYBYxemA/AWJNVy8Y7qr
6ZtyLnR8MVO9K+aDIgdF1UJhjynrbar2CurYQ7ZyvwF0sGNqQKKSfL69Ju/VkZwJ
Ea04R2OX+GFvHIYyxfVQ3lrjIuLOC35IYmVufyC7z0vTmZ8LkPAQ176HBEzXCzP+
7jI9Uj7exKENwP/GFale7pYZ4rIBrAUsTMq19CSxUpLF7OkwPq76HQ3DkTztvwd2
3Eso57r8B1YFCpC6vcqMK/TIXt9FN7qQYyaYWnhtwGN7pT3GnPJ6nLzU+knSg+Z2
tpNTOisj9+eo+QRw+KPBCnmylZ4jpPLjbIUCwpQkr7ENosrExsU9JRXZWci1v3eY
r9riuIqfcjIodO8Ddh+6hjY8rzyBwobMbP18ey/DlFGNIVknPPNOVL8JHZgd6zbY
i/ivhNI2VHdgxjXGifMd7Dur0hRg9/FMlyRWYI3e6Db1Zu7BD4NDSEHACia2rFkm
FLu5Fjbl1Fty0o+hnUk63r4ALslUitj/dA5Tnf6sNIhuVOVZXuVTaUyVaTuTHEee
5N5Z18Yi2ruZ7rYCaHvcQLInAi11sH7pyiE091AHfLMZA6PCr5SuGE42xdyNAOM8
q9KkLdMNjO8c3J59no5DX7nDlR+9pImA90pkVfIukiUMYJF+fIj8RHGwlVs8jJwB
ZYgC5+KssiEsvJWB5GQYQ6QgYcNCo4wutFcflsh3+EF3Rp1xODwxFhvN6HnNrENd
Jk2og+bcwHmofk68X0Ncwm/RQlsywMnFSaMTF/KaIMMe6nMakS2J+NYV0iHNa7ce
U6ZByZKiO4qA6xadQftUq+vd6QVi/xLfV+FtWHT6Futbx3ucbgCyXENm+JJi3/xm
aT/YGHoA5+pVXP32NF6W8aNT5cDFbk3nEZd7gjbhgM5/YuF7h8ZDhLmhlcpYAoKK
ZXXP8odLPhXiieyb7EjPqBAxfZO0f4oikWIzaRMwWX1jbyrpluEJ+eIx0GcVrhkQ
q0RsebWLekJISkSuZH5BwK3+gsenwFzm5m5tXT7doaWG9E7eMPq+0ajJ5BKy0bnI
jncJHlmMDeZUSkrjkndxO3C10Rzz3pTSWU09w3O0CURG+mWi4Jy6mqTZvacKbddW
jQ4ZGdLbzuiiMVuTOWiCI9ohzTXf/9/YFovAQN+A0v7IcEyx8LmIk2TDVMD43QL3
sosodeV0fInFfKIt47YkzX7hIw4fJGhPl1G8ZHlDES+9HEkUkyJtF03An6J9BE0Q
yT9A59W2v3y+zFWu61GGl9GK5A788Tbi37iL8epxjsyB1ay9Uehb8IVPaVbxOwZu
Lrw9JoILmLwqAqsFYE240LNYnwyytfedtQDLexvVydvSxFhXFgfAr2OQ9VSYLvCz
zWAje7l3wlcenyZshs+EOvwuTm7LIojEPVMIDPJTdh99685aroEXmNB5hMsdqfpL
G07O/L+duyQARuwexk6S838AyhpA8yFY9uBgq+9XjK37te5MsrF5hjQSj6CfzAYP
aIo4zFCCgFsDh5cbZ9mXuyoBdYVOzzHqWB9x2XKp9aDieLilGovnZ1Ja/C/oKMEB
RCNfU6/VkIQPldYesN2H/8rSvGoA/fYngylb14AvwYnSPpK2iwb2YMGrHkLz/SQC
vtYi0jXOgXQBMFmobiP+/3rVV8Xigi+HkzU/E1GTxAk5UhnnHu9csVvWAB4iYSde
S8nsleWU6IhK4p8DkNRSYbMgWwqGO4+lQnttUbKKTdAwjrlUTEvoWx71PNkB44pI
F1x38gofuhxg0ECZMm7tFdzd4/zZ8hDmdt/mTYum0ja8MLeDkQtEcIAritJrYQbY
Mu5TyodZHg13OcX2nVbvq3oPelOUcmet1pwq+E5hOrUeFGForNUqrSDbnhawTUpz
8L+X5PwEbuc6hM0PR8n/uTz15FIYUAcf2u5pF1Bw5VJ3gpHIOVeprR0xzvbJd/kC
Cn75sl8CxXVtmPHPDRMiDMROsHE/nNYLJ/QXuAPpii6l4TwwxpaRtKrbGAiIupLh
QjB2r6SniqJbuAjtohwcsMcPpBCtXjQOSp8qCI3hrFx4XjVq71hZJ0ium+s1mPHL
WRfnyHerPNK899iBxiLKxzwbqYjaaRQVqaM6YKFtWVMqPbpJrVx7F9PggA9sXzhs
BoSmh3abW+3DtsRdgL6t+Jte917X08c7yFVvsvmU+pIJnLkVElm0kcpbBdOCnoJt
apgxkGwXmW/V4hhpHMqY6WNsWLyu8MktpJfXHY6W0DNr5m+h8yNNc8gabIXAsiMS
FL9yX7Kk85KquC4sm3/C6t3GEGXLcGu7vWr/IdeDI87m2YhAJ2MXii9DsF4YIPtk
U8DMgyqc8PjGffCWAK3WtVh4rdhM0PVYQrFTXFITr1bkbwIRZ0NZDSgy5MnXPtFN
bL8+mOVo9meU2J/sBcKsqjwXduc8Y2xC0j/8hCCJTgnYal7AAPpwZrfudJFZTU4b
vjdUe6zc4s+gwu6rO7apLp/lP/LzhVKqRHfbd9jPuWrrhNiUsCcwgR1B5Vo+ARiG
TRiT9g85Q4qAp+WbB5hP1RObpzyZO/SOkgpn13qxbo3xBVAexFKEfg80DwOy1oX2
OgSEcpqsdBFo2zv/Tyn5HHpn51JwnMr5pUSamankhHlQbv1tsXJKn84x6hbhOUqs
+I0CNL/cqmyWYVcP84ks+Yhn2Jqyxh5i2HMsdsg8Vv8c7Zfoq4V4XWy3BO/iLv8J
w8VF3jwdfiAgr11zRS3pS7ijgrM5Q6OApZ/IHNlFZppwWofEMRqMDtf5c9Fc6Bzf
Qs7ZPeLiBSrMFLteCNyfoBCwO5GKCPQXWY8Fp/w2Qtzy0aGapqEYEid895MbwkWK
yp8VeU0GUN8+zPcZgJSWz6X9vDs8iSEJFL4heciNUDYOeb7KQldK9HXq+UkIv9RQ
FDmXcuJHEvFf9Ap725BPiR3YCljWoZvvxjqwArG0lgqzmNL22pQ3WlR11iab4aC0
p3y6+ZZA7jNry23MZKCn1hpe6ZpFvy/w6ycRNJHFNUvpUGhmfs+XlH39DIm6V0W6
frvrPIBf4ALFK4KxTur+OknWwMJrNBluFSXdp6XRZL47GK4fkaCqlyAWMhHZUaH3
awD4yyZzV2zxHtKCiQjwL//Pr7XGGGTamLcEfUt6MpCqicOL/VRmszb7qgfCGHgT
qgmO1dFgf8PramiUttkudX52ARF4eoxekvXOAzIdxXpJkmljUoWnQbMnBjrrN77N
qDwU14UePJ6LdNq8db0juXJL/O53p6iaH7aHnId+3FdjQ0EbkM6F7qHvSy8EzATm
iAPRcfZACF6IW1PgKnY0/A4X6X5HIXWI5BTS3mTQ4CCtVqkFUmKfxws2hu8tBvDE
+KO+KIO+9aeNXwAoAs8t6cbLtMxge9p60JqOlnBrOQNqC3zDMyWLt9JW0VkfGrMM
onRJ+tu2EE+ABFE3rKonev9z8N/RZGxsnV2OgE255YrT6alFbvy14rTvtOoKrUG9
N5bNxmzIzbiMJLveR/vNFsVDa5XLG+O73Je6Rtfw4MrmB4qa0UBcRE80hle7nM/L
jSqkt6eKzH4Ke38uZfZs7SJN6x1VMk3a44htvWeYk90oYJsUM3ad8ZykrH8mHGjo
gyc1VfnC1UPMnnLCG408TOjBXfyj6ZftcqKcIXWgmE2rkrcUULSaaXJWbCAjCbla
VuMLtmVTj4pNIwkxTTr4WKBgsdQwnugGYkJ20HNNDYzWPcP3IzOANlqqJ8jFhLK2
cRuylR3F2wVlBYptLe49oXVrrGFthXPW+3ZH3i6NXvC6/PMv9mSb+mzyEu9ak/s9
GjfLLLg/iW1T38bR5dMKfW0tU9k0LaT9EZ2GCrUYN3lE4ENNJWNnZXHmsygzTI/X
zCnXhDukTehUU7XXhqVBiG+SDhDRBZMQQcd+6ssL00moqpDUOHtKpc7mW65ywOsH
hT94CeTXxYuiHean9LK2TeKv+rnGY1VRgpsQOBLUih24K9EZIn0gNHyw2+Vn1KQT
pRPzh3BvYc2AtyfksUMgHII94uGrr+VDFp5EE/HErsU12Nl4a3x9XzZjlzkC46vh
GgLOpRBomHWHKnkKsjbCk+jh0g/oU0o50VlsLQA6VuTveccMwmWlovCLdSUzsSYu
VjreCLhKrA6Izb+ev6819Ugyu1iKKqMumod18MsF/r3f5HgFwqCQ4gzaQ5iN+wr/
bsot9P5E3ypo3gcRCnAw1MIGsH90WnyxEOAM2zPiUdcZFuT2F7oKJAXuvNGixrjG
BSzvFhZXppdQL2o61rVJyYnGcy4b6uVXTOCtkhtcMOEBVAMxzafoAoNofWJnYbOQ
U4cFEn/SyoWZA2KaZEWiFEI7b5L9xb/mydwww5gV6gvpNvErFzcSdtNNwdBnHh5C
6P/LzJEGssq4NCnOW5iJzRyOZr8UyQHLozZY0QNOB5jqzr7/6BGlp3VPnFaKAfTD
gr67gyo11J5DvSkR8XmFJ9PEJyuoAdDRybK6cP2LxZqoUSSaruyMg9Byyi99b1gy
ID8ItK2NzIMjsurFwo6Gsf3XwqsLl/y2wfVNyfbOtNUK2o64AYL+WTy1TILEgDP7
XufuEatqJWq8AO1e3aquqar74pzRYNSD5pR/TOLq1gT8KTRGS5gHcucyTGL5KzcM
eYgn/pK5wmesLBwrsCVYPorz6fjHOuwl5aSXvuNIt5zh6d9JG3QImLV7VyohDFy5
Cg3WZk3RQHjAmPM3nSEvifRkp074hl1m61AV5l2WdIgL1wRV1NI46lBaoJhRtGVn
1DRmhdKEgY7n+7cHMI5HE1zsVPR8lM27gQLsTe6axQbjLY/4msgbSXjfscNTnagh
QWjjfAisksqnEXDSUXVHfdsibPbSHTUuxEVKp+pyMwsr4TGoBKDJUpx8kLv3nbUv
Y+JKQeM+r9pfx8gI2x7/clpMSxSA0o1eHfu2OFq6i8jXqnLAzXHpwH28b2StXt2e
Gl+UKJLJ0e0dQbqVDvUdQtx/cAYhN3CEdQPgD+ehpaLTIC6nNJoOp41no6Vxzm01
cCb4IFMyb1MaQ4F238zurqhfXCsYSKRYcTtSnKE1SNFZJUweshsmRj+Krq1sropU
Ngz52TeH25IfB7JVRIjL/hvjam1yZxy4xJtCkveK7q7D76kNJ0rW4wLhtPC8irrD
LAlgrtQNwlZ3JoguzThS9ALWMLrqrP5Uc2m6uVmA4u4oZVAiTa6M6XJ0u2ec/rzj
GQT8NnB8ZOyxWufgTGZ3mZnO88ayZmihHZGTOWQza51it2LPbcXC5fPn0Ia8/HP7
TP3jFqM4cYMHyDcveDD+Rje4hb16HDxH9QjijA40CNVHgVa4Jg+3BR5C+E2yR6DW
iCLRz7QToR3spLm7Xj2V8PiOHjmyltAQzFnNlWII+8l+voA+rw3K2PqbJq9a5a3f
bkvA9OrlbRODf6xGxZ+9ZMVhk4eaFH9cfoxY4HMRiAfdw0R5LjEOFMH8IEhzqKHU
jcDCmJbnhRSXWhFNfwJDOBygiyXgcn3LUX2yNNDhpe6/Lb2vQEk60qZpRlVesZZZ
ms3WMdSlUG1zYh1erE2Y1frgPzydPNrRE2ZOx6aDuDl1cQVAzJ3yW9bYdpjRn+m6
0DPcgV/Mv/HAmRkEjOO/Dqww+KrlV1B6taR4vJ2/bPF+7SziMUIrSlg+eggNCDFR
SS7UC2pJ0YgLkk8keYeF0u8QcGm8K1bpWBJpllaoOb007oMg8FCRvmLUaP+cKU2a
3/MSbiXBF5edgEJB9P8VFHq5ik76i+eZgamg5vi+IhkLfFHiqGbOsO30wuZEYait
vbgKjVhn7m4fdfB4wkaoNCUtWeV6VWVa2NOMZ0MFJNPXdpgasbIqf9KlC71E+EZl
6NRm6D1DZMX3q/ddfPmk89ZHQ8HmH1vY3/RrTS+THH4HzjM1ohYlj15DCx67x6IO
ZrP9hDXIrZN1UiUja84d+8RYFUjOaAGJbAwHGhLEkoNBsL3BZfLTUbpNN6rmJvop
zuZVKOu7Sz7wYFvdVKHqzKdI5KSBmeDACyz4VHQmQLkYaDsT3OFt79vszgR1UtQ+
2arxjvdoPNVyQGsBKvp2v6Lyxgp4/FwQWI2XnRmfv+F0bfXDe61okMXXwQAUXciv
Pa9gZBDr/j9uBOfaW4k57XMQHGuWeGO8xuMzYlmeJyDi8rPgotPpNCv7+KpZ89gi
6xIPQ8CPNNk8E6Da6eGJs7s8RbxO6J39UzRnw9D0vyomuPkKi5fjpLlMoXcqZg67
58t8a8+6Cc9cnJjO6T+IND3NP1gTQ05zyLddLK1PVUtMEIOKF7AOnsMQ7TCeLCJB
iJojn6D11ticKgMIAAGaVbsSUwKpeSNIsqSpmXQW3eWj6ONvkZ9d/IVxvmMc83xN
k7ePydEdemIMhqADo9dl5VhYf0SjPxq2IzAaCV747gt2sJ/U/5bSttPXAerb48E/
EBT2+7p4tuAe4Zufbsbn/lvDM2S3scjc+OcOVW/IpqQCHTLEzhNw2ujFdLmDyeIt
HYY3M9IZ1WajACNxoG0KEIEUowBaXohMdkJTn5DbgE+L31Civ93qhUTnJY253vF4
ClY9K3Nd8xTa6KbZEUkJtXWsRq4g9XCBBB57ywJKSU2snwC73MjS/V2jcLpqU9ED
5vvSS1++JLmMGPqs1KBNgjkokRzxknSjYqPrxwm9+/Fss5xzmCcXIERjsbALm/mw
WB/hpYynKWvWeG9KI0C7bQvQ6J90JzQEVIIqWp7evWOOx5+ZL5f4wQJ9L9kJuWSZ
scX/G4BVNIjnExVIfX32gJugQpHNInSjhvGjea8uQBtRUPKVJxxURpn1CjADAAp0
yuzqANGXWGo5eMDQMqvr0W1uJ1d7pVAnFFz6NjjTRiD6sh9dAB0kMprCuiBaGnSk
bhP3wZhvgBt/HAMoLfotmwe5Qs8zWRggwOlH699VJuRHWOcNiT0fEAlOp89xOWhY
uJXID+Lf6E62oN84ZLyNvfERnaK+JPrq2Y8ceLsWtUiaQ6xed4Z42PnxPD+MRdYV
KyIWmcvzNKirAkDbhK5pz8nWqe4i9Z5Uc/T9cGGlXRwMfK1roFyBEgQVgFxk4HBn
2JFnjNpW16RHFqy7iGChR1jTnJ5BQ7xWo5j90oIqMXGqrbNBlhzCLEjjmqWMKPA5
tPRWw5xSy32BtOivLy9/+AZEQqakA5a2/33QYN6dHswbRvnbbWWOROJejeGOW4ql
EeLuWc1HAR5PbyHd7T/RqxUNDNTxA69uWkmGtHI+42BSavixrMIVeGK0CQH1leBL
u7KXHXQr3D/ntVFIwnIvexCQZ6GEuZRgPUzeHbvrLCkLVpWehUhoB8L/cqLKYe4q
ajtb+ah/4txuuQALzK5OEs8Jh8xEVQB0uR1hHpgTYwLrU5gWM4tsjMNUU1sd1gFp
8rvgbfkjF/szBFBAnIQ4ROzIk4q3OA9oX7353+njQHFDOtR+7zAokTIIUHquGyYL
GS9OpsgCV9oK42Ngnew2a58N3xUPWztk28wSt5zYeleFxRn0YyrFlAIkwNiTcLU5
9960hmx1gp5KbMuaPHKkQ7QDJk3Je59bbKOQdWdRcOBjqCCe5QTC8alP/uoYCIYp
TIP2vm1chG+XinyvU1iK4TfTMB+y8CxdcNxfow8C1hFn+5b3fQ15kb6Qgof9b4vu
YzK4gaAJilSd741oJdOFDZxePyA7ZyRdLNC8T7EmBy3aA7dnprX/GTiOMpRnDY0r
xxJk89sD2eKYQYepp8WYIa1zTN6vKASEywRnv1VaseeNc6KyrK1InOkoSlnyhlhf
csNxHEM2BmP159nlvrycTGhK4V8Tdz0NQiMqQWh9aaEwpo8M/bjyzBjM4O0GwyNh
IZaNjuRrPuOpyEBTlGn+5Pfx4VuWM/Uc71JHr6spWmOoy/3Mg+fWawIvT3C91+oP
RVKYNT97va3ZlCBytsp/4YaEIOOPkGhmdZalA7Toen/5mpc78r5psDlA6r38emHA
B864RGqaR1f1QTF5VS2idn/h7alj3LnmLl4LM+VGSQjaQftGPEpmaNaBrBoa91Uc
nVMnRlH3LLybAXoYvds/Neb/R31SHVvnTPvh2hwiIAFNeksula4oESprCk9nWhpo
77BPo0EeTKHdW5GmQwOLVoPyfNKJe3w9FJ1vfqX7ZgJQB00tMyW0bjwhxjm/F3+P
Qsz5eIj+HY/PJ0DI4P8L00Rth59He3/g+kMHiGUrupzgZV74tkQe3l/Q7POyHs7K
qYr4/oalYuhNAyK99JMUq6V8+K/xjsd1MaeQjglnr8bDzP5xLph/46wl9R84+h5V
FZINBpnktrwDpLXI/UB1W5IqhucAOKIK+OmC922+tT7X0H/xGigqeiUBz0wBJaY0
Ctf8xOBXFVsXF8WG4FT12zLsAtBI4gqSJwC+V13CU/kYokwsnrFMjVfrJWV8sbG9
Y4rW3e66UoJ13EpEZqZaiE+36Ancb03FEirJ3IgL3ZtUKQOAGkIU4KKKXRkE0DPu
PzYqP8FQ1Ib6/2e/DoPsp9Vg25Wnc8h75XhV4jmFOIx8wPhr6FmKJzt0DefEAxR2
lC15nzV1bVkwpgRdeODxMcRC2wSD+Qg85DA/CJmKD5C5stzB1yhzBIYJeowBGs1f
+oKmneOXC0msuQG3H4PNDgNd1GPKie8gnLsGSjg3i8p8TMRAh+Os8pSN7YxWxgZg
bxR0VQPep6Sgg/YsP0ilej5vQfS2KefmMX50jvJUuoXxpsmQmPu8Ore6zMIQROeY
8aIUlfki38y6XKV/ItGEtqJg42HLUEuUvjBcf/HSfMzuXE8yscM3DlG0kKJX+xNg
um/myzGZp27huBJsacRm772dOKB6ci98FdV0rAybMYcB2jUua/JW2njCmap5cPS7
DDB1zPpuJdOPMLLIIiBhrZSAWGy1zkVfyuU01v5TTZdUZ4TATwysqxhSstEyySHZ
WyBa5POYdQTG00Rq1GZc8j0eSAe04nn/1Ab1/dUdd5qhRry8p2yym3FIZ/jJS0E1
GgIZ+ZNaPyq+ff+T2OkWg3ZC+ey2a25P/hph/UG9VEZhRG2M1hEDukZUqKrf7kHw
UbRn+53hS515KOcJWMj5rquoRnOG4sdD4m+axDT/iC5ikT0qpmDmGYt6Kd8SkGl9
azBJzCRMKAi9bayrhs31TCD80A8N9DrxJkbbtt3as8CpL6wQtPKT3bC4U0kiPlNT
gJPcAMMP0C4HkWkWew0QD0qvU5yX5c0xATXuZEoDp540N5i3n3kjIlkonWu2F/Al
FLoCCC8PATEhKQCLI784acGcaUXawEz2WtkcELy19BjOV8H1Lxyha7EOjjx8ga/5
ZUKmQS7zr7c21V8GmcEdO6acn5JHFn3pc7a+srTG4CVmUHPXz5OLkV9hg0kkUwm1
0N9+C4Uo2mCJx+fe3+hx+ITKMs+OnJWifgTy2XO35uYI82gVcxevub9B/upP7fmv
ZOT2R3fZ8MV3Yro06lHLJZRBCPjPtfUimqaP/PvxqUdkENqScCaQcII7tuNlZBtp
2GXb2/qgrjBJ5819pbdK/T7EWcnyZTUe5jRPr3nIo1rJB+mr6Inon9aXwsgbF6Nv
B+366g8Mp6tUBqRr5jEAIG9D1afisyq4Od/rP5I60Rje6tArE9lI16CAleO2Zd04
2ulKewHojycNrBnyRURQDLceUhlL+ASiCKvd0nudnwQJu/X3ihQ4lNn8FsFaHCbp
jlK97Mj3valR6BR6Mb5CRLsmwP8hP5Pjw6XAOs9NDCQNpLfV9WNig02BG4dfvP62
AIHyzGC3YJwrr16H+wXcN5HH8XFEd526BitWAqgl2xMfmETUbFqjJTyUa6JPnf5o
Rzl8GxR7hnorqnv+YWka39j4pxiWRJZ2BJ3L598HYCp8WFue78uRgYcZwoxmOzww
r/6apLlecfoXtmz3FBoVqlj2B1H8aAEm4gLIC55fiX/9gDnSIr3L3d+WgadQcCSr
p28d7CsduNtos0eHB46RMoGomv+btptNIoS8jpK9F96a+0V07G7q7hlgs6VeC8rX
tz7zD4iC11RFmyL7qZw0YVKGNlahoSyQykVoET3FdBg2p8lofxoShvZ8xcjdt95n
nQxRhnEo7IJDvqeZAvS27QMCFa6bJYVnKUBDzZRnotYL+s5JBkehKnJJfVnPjQw8
N6+XqibAukBwvU8csj5Tl/3tLRVvFQeSRDGsUQR7qcGvb2WKIZd10WK1l10TuufH
PHEw6I1XmaxKByvlcG4Q+7muI3qNgJ3C9HgVJlHe2/220N+S/0sy2aRNjL2ENk9U
ClfFxsewFcaMNmT8JIoYdQn8IOrO94q46UIQYIqoHIb15y3RyJMxatFwkm4CpgkO
0lOyCDWe/kNZgQ+x5dcofMV4UnxWeuZbe+F8W3kZ2OPM4NOpY3Hg1FrTLCNlBUPm
BR1o03uzkmCzraNwbWf6Mh1szyvLblKKWLCw394c5dyRM8tnLLi3BdF90UGPwKym
8B5duev3Vx1VGV5XtOxCPM8W2ETzx9vQTAEuByPt5x09A+b9lJGbo8JJPSF7PBoa
hdu8m0j2qLOoH0pbVBBNaT1blCTm4NyuXCuHbpYA1I5kckBejhT5cZA2PslOEHRE
1ZI5CZ3Wxz3BVG0Z9UVzzbs51tlyVCTeLAYDXzvNtLz7+QbcfP+rAtbt+exJzXqs
QMtaExotXRRkk7g/8SpVaQNvsu4910a42ftEKn7vviMFgYAB0RYMMTht1FCxo7I0
dJw8GWd2e2IG0vGctdo8A99ksvT1QC7OtGvH7De260skwMHjHg87IwBEodwan7CF
MBwQU03Aw1Qkm/RvaPEGv44J+dhsCz7YUQU3Qh5CHcG9ZP5NbGQVUZpL4HGgutFc
YWqusGQ5GaGaj4JfSy+udF7bXt8Uqo95QABXFNn/CEDZq3/cesQH/WhS4ZhghNtR
tUYnag2V4yaXEaJfoSK3XZjZfYyGXL0VH7cW0zRVoJrIaxc3/KkYa+soRnVmrtjJ
XcqnG4T8s9n1noY18YFPNpyWe3b4KmZaxWge2Hqi8PJS0aXNTHofXtMfuVvzeXH4
/d9ObHyr0elTxIM7xkq+gpRFMlU7qPFx8E/cs2N/WkczUXULFgAsDrKZD7jM2wni
RhBuiK7AQl2YNoEFYFo6SaBzYxRF6KamPbp3G3bHGNLLKZpimbRsVm2oGFz+pYLd
YVbdn0Vw7O/TCcKlR6h0JWByfDwc+78XqYVgocuR5RJKR/sqcDTHVaaEBCzmKR2s
0zDtYB+TaFBsLuRsfQYlPiCRwH1BRF5i/jI8TJuq+rvOM9R2MTUQ8HhgZO1wKB2v
Evl4kjQl+9b1Pu5tWCGouWz4i8vIkAxZqAmDE9uVD3/1a/TNKQnDfsRE48+9G6l0
aJNQALlz9K7HMfGuXChnmYh5llrbrg8eePr6/9Hz0Icjvc7hh1aXx20WvzuqOts4
2lLX0ttcy9na72FN8OYX9N9z4wzuHKibvQBazUxyjNQzYa1gDSpMFkjE2f4JDOmd
20+M6pX0sDeCzUjZrvA9gXy1UxrgPlVGUDRfhmT1z9A2nIGt/4opcM7v3ACVxh1v
IrT77Whugry/ghdHppTkh54AJoIbXOKcpOpGnPx8tR5P+bJRsXll/LL7muk4N9Hx
ZqjOhc7aC1pd4xpQiCuyQo26By4MNGjgI/HSPseeL+6LKVOUZ3Wp5pSerNIbVuiO
FrSFqO63o+mLmvMmgGeduolFocVChcCJd7eZTa2z9Qn3QuGklAh+w+vIrutW/dLA
mzdenp6Htm8KOdtn1AR0GlqPEyPI1PTmy/UdmYb5adTlc6S7YNpWWJU2JKqefBPN
9CW3nIqmR7bxNDQT+oWF3PQrSnhLFNUEOksnTJQRR4sIWH+7gNgcYZG5mPQSvdD3
nTgf3XSHNw/ko6JO9BEiE2aVVFZX0R/SgmWM8WpZT4mnzwYy1+bNLbAQkUIe2hLE
t+T42+0svdKfeW3hlFubxiDZnalynwQBQhGha/t7e+2CTA6m3zJArmNWXqh3tPD6
14Hsgu2X/D1mBHrRvJhALcK0NlzfeqzZoIk+V55TEl3PS6T33C4f2v7HZjym1S/e
tD7SWPQWPgrfT/CDIR57/wVmcxZI0tH6VYzAStYg4IHRCCey3iqR9e+MkgYcIby0
w4UftUFhVQU3him0WSVlSZh6Ap30PhTsGvSq0aai+qQgdzIMAkShHu6r7KvgVXi5
Z32Ryx0PZPMN60Gl4TgKMdJ297bziu+vpXWQjLgh1OyXNsfJA2WT/mVo5xM+5xuG
tNUAuNOru5cEpVOxVPNB8LF3QqrSJfdCvFfZtMsqyPjFshSmad5Z2QdNYM/ij6D9
V+0Arug/zFERFaZ1nQQiYuXV/QEHsM+ac5L9GXdajhPyLgXxx7lMSL/GNd71mOWX
mqo6o0dUxd73h77TTPaLdNvnrai3tb4x5jlOXsAoiEUW0e6AqFLz7B1XVdp05HjZ
kq9on+jE4FQW9tsvJUSDvkNqTEJxBomjXdG6weIXhwW+5V3DctI/rgiKzlCA1f0Q
0Ur94ogfLD9yatJCa32dDhtX8O41fSmq6iG6/GknJ0m5frEJwsJsS4S1BJtuWssw
kRBuFoHitEopSPzsS2HhwgsSdFAmPtF4AKM47ywa6V3ndNto9BQxZ7/EZhcusZ1t
kMsla7U0GoUQbv6fSEXJCye+TMDshyDb0p1z/jVAzeQxpNoRn51zlsNNaKSqtPm5
0Kw2wibyhF2dmpKdGFBiZieogF8qg9gLBTuQE6lRKQof1gQXND28eKEzOtIy6YTO
0NS4t6ZRij9PJcVeyqtxog5mK0NrZMCQCiiqwhgwWBJylTVQtsWHYgS6ZaPRR32U
UP/xdj0deBAHwK+weteZxq0BUy/+bT4EksZp7/qE1KFBNQrydXQL6M5zemxD5C7s
2ZlHLkfa9NXnidoBkJ85fo8VJa3I+d3CeLtRVb3MP69fSxp+thaOYuIWDLl2OYJw
rWlYTSnM2+jlU5iImuZmwNt7RjMcLHp20GYXZC471n80nV7W5J/4X3LOe8F0p4RS
Yexr6XIiFR+hHhCXmwXvTG4TdclSCk7n6uaBgK0gYDgTrgK9UVPQXF6p0R1iDC1/
MWXyjPrzPIQQ+RtTFe9hX/EYX3MJhhTP8wXcRt7iNhV3Mc7+I+AkNzGauf3Um4k4
sDpf42Cf74lwfnugri0qDWj7D/ijN72+EHxAar42XhC1nMI90g5GpkExrNIuRg+E
ATo2rgGngXYQ3Jxcp+Xo7mvLnXnXlH0uQf3Inzy7uhb1JEaqrYovOaJ0Hy9aHW/s
ET7dW/4IyYUWuK0GXgcfAa/F/u69McIf2CGxT1vKpsezWi016aj2kWwMyiPPV+/p
2MMHHAhIu+qNPkHNertK72a/aZAmoOn6DDQZXE5wNHlbVbONsNXNsmX8WHLsOqNt
pPvpaRNNNo5uUPU9YqiQyc5mk5HMgCwrgXQAzrf70nx4P1Zkxv82bghIi2yuRbFj
sVDgn/vFYi1zQbP0ybhv4lWzdnmh5X39UJFjSnBFKDCqryz8SQbYVILUNydebC0g
nQz2rrOjFpOfhQsX9w41ZM5PGEYIfe0yS2MPGUl1nODQ6h0XZ3BYHq/0fyRZhu/u
U48SdaM5mg3eBethGUPlMRTwF3JENcQ00Dv1ZiY1GS6g/rvnfv8qa6i0dSo+7jRy
H7j77PQYmtNdm9uI+Jl1RMsP0Dyn3z/oqNqcWRaanwVScjoKT1dj6fVrfX4wJTw5
riOT5j6flt1DKct5N/A8yObGjWHTXCI9Uyo3wrhCD4LixEu9WxUTYS/NV6rtyHME
qj9z6cUS1uAyvcPyCJHupW8m64KhmsK6vKkfuW5v+3hG18TbDj1Gpo/6PtOoJnMf
RM417if9KX7U5L/ZlLRWU7YAhiQjqWEan0Xpf0Jj+ueZEcK4t0GN3sYQ9eyjclP1
GK3mNWQMtz4zMw8mEuQjATECXSvOsXB91ON367VAPWnqIdHSqJG7/ZeC5tli2w7N
OyIy/wfADeZljV/nxuB6o30hFTnSb3NO0LqCgWZuD4YysdFMbz631znQGY6CDUfT
TNYtHVpJKwBaDBg8vmjE7sbyVBHtkgf2w5ipP3B9vDArJ5qaOC9PSAQt6uLjzGDT
iwUXp6BDTsjZGYG1L/xpiTmMZYKr7PRJoV2DJ6zqyroKf0DSRt2sFLbenlBOMOZb
lvaj7JFil5ZAVgiD7TTahJQWcdG01pPIMh614vn3yilqCDYMVJ+/HBQIz0qe57w+
aGlaW8ptt0A8fgonkyupMtmkRjsI2Pyh3JE1nZe8nibsrqpgJcnAKcUCXEuA5sO8
u5EmiI9stnNUw7LUdghksxdn5ZB+sDDG4TbJAE9F3ctALLWmzwaMm7HrB/+u4X4t
S1ik81zGhU5KLmOkA3mxNjPxaK8QU24ly2BsHgWFXdNPUiucxkuoIJ9SiI7uVgFj
cS38L6w3AX7tvX3Lpy3t8iG8a5fD+OOUpzs/10khDUoQY5q6InWDwpQIJH3ZAfav
bm0dM51TCc7MO7HU5kpn9AOlBGdKNu8OwallNbxVDKpSBz2IIdN/GqHi+bjOzfnA
gHqjl++mAJX9rK4L/cxw3YBdhACS88qJZrFQlKOHJxpMukargq9jyZ3JONEo10Mj
NtwTWGi14nZs21ijP6VQsYrcwbtmAxArK0NNQYgIMLbuXsFpe2Nk+8P8ROMzIQv4
8FBl+xQXdwOsGTvbUnmhU3a6eWKB8OYw+i3rroIAk7u0NFHcdzbKhpW3pI5o1Tfo
A2HJYMP3UyyYw96OA3Ya8wqlq7xMf3PwWa0Y4Qe91wVCFFxFCmNaBGA3uPOeJDP1
uvZkJxCryjHkCcogXd1CL9heYVr3TlD30i2d0uyqSYRUzf7rCOGhOXHj6PsaCCKl
ezz5TP/oKe+QM1oFRgDCdS9bnhXguw7SabSZUO9zCq1XKQTDY3S+U8voB+gweLlG
J5BFJYW1HwMPdbsYeb2jvAxafjwimnAE+wdW+DkdjME9IEzoOah6a0WEHmSylDMu
q8vopTumIBocn2DoFpRgFEs3KY29gjoEhQpqoIGyhLBxr8sZKioPPZRjR4xbH4tO
5V5JsOe/QUWB7S/0jCaPevgP4KadDrxUKu3PbqMECQuY4rny/N+a3/vM17+uVKOm
LJFUcybcw3HLtcjDOJZ6Fv5Xpgz+X71jOhQaP0EZZzob9pMq3wjPAmkZ+ZleB3Us
s9C3/Fiyls4yWT0oH5vY6YXmMqes25hmqawieY6zD3lvsrKjlFGwiNAp3/QRL2og
9jv8MkFQvZHBGXiMGvpJW06qBUA3SSulPc5l2rNttEHZtG3Tym8rqIxB7hb+lLvm
fwof1iDVmGl8Z54TFtaKOL40yqflZVe2wOMKGcj9q7xAgfBA3h+m5PAjoXDhCwYk
YuoQFLIjCUEm5GgiqbcNBWJrWfQcCyNqz7Okj59f6XShiLwjPOpVmk8l6rHeyWDp
SXuS0JML1+TMpCD2UFO+/SzTxRgMdFdX9YauGyM/rai044BEgGFtXW6UaSKMOJJs
0qZCqEQae/a0QNGmvQaXUliCzbXwlhgAjz8uXIHtxIInJ4bkgW8wMLlGtQPxsAjv
RS1sCG93LRZama3bWHCfAOAcgniNJ2+9qZtKR8dgT8lU0+SzkgLXp3B8cFvHs+Ny
fzoCVPWRU94bsq+jlhh8I4Md9+6mPWN/TaFEAN8yci0m/HB0BMlre3cfE32tLaps
Ah0K3/XJ5aLIOYiyFIY/5Agl5SsME7btAOQXCNcy0lOKiuZuXEfl3J6dgKRI1DcO
HndS8EYKIv1mppVu415wfHFI1ZWgqk7Lfj9rVdzlcoderG/9oDrHsad37r/fMR7i
dMxmJeBONDMKdNwjhTqRmrfwjppKPWmar1oFpDhVh39XFUqwy5DFfm9ohLW/Cv1t
6VwiEA3oRqVZGavftY1WWlg6B+70EbuGFsS0OCcGVDFkfxY+AX1OmDvOXTjgkqQw
YZBXNRS7665s3yXgReVHL8zNmxWXgW9qPXo7xoHDcDhKqGQxGg2Aoe1xHsZdJA6m
B/as2FzbjwBf2XFgI+5KzSQBluATF4JFQbCWBc7UiO+zyiJc/6hWUpzRYPjARsOp
DL5O19HiAPp7xax0gZ6dBal5UxFSeGaI9jiRGRsd+hVCDxWxX3d8y8hcxu0S81EO
6G1hoh6y5dkDOQL61GPsW8AV3DpyrGzLnicyVBYxM/Zgwt+Thn6lf2ocbMAXhKzu
dz3xcr+hh1BPRVhxYSTmzjUvs/Kn9a3LztlG2Aw+/j37mFsQOCPa2O3vrP6lL6GE
QiPJHaM11B1ymDzo5mMaotonfsMhaKt4O7v7kpEdExZQ3kT3KQ1LKx/gTMacMN8Z
h/f+MYvXrmc2bWkzrnp7FcjlN/noFfcY7kwTM7el9AecMNiebU8AtEspSLXDSrm0
OQLvtl3QWclFIrY/NSynDnnkhQWQiOOlgMLKqy+LUU1dLCwarZ/xsaSY0JL0NwOu
GBNYzSTGqDIT1BC2vnx5Xh6lR0635Hqf/kPUHdfkuFXOQ0AauJazuxEYBylEcwNY
QtNjmKnxISGLwmownpafRcHOW+pnG/rkg73iX8YYh1qi8Mq1H3wyNATPsLYPQ3S5
U8IJHeU3ERnDbuMq6/WLY0DrXiCH9NjkdJ7YcFgJUl3uUZyIOdKnedbXIn0BDA3c
6B0Ve9cn9jPRZAx1ZY2uDH1TT0VZ26Dm9h6mCblJ3GJ+VOHkVVjo6j34vEoCWalV
JoTI/cKXmbtNC71oT0+3JWtgA0kvYDHs8gdXqo99+BPNIPJlXvxb+EpJTsAEF0tL
GQZ3YTPTfzFu6Wlw3ru5KG1lS1O+2ROKx39kwdRjQTEwTxh2XCMYawXexqMwSy3a
MaU0r7ZVKL6NUc06+ocSEnkUVk8WdouxSfofTiRgJoqH5D3QNXV8wbrlOKYjcBY8
yERTXqTtrlJpLgxUsb3b7OHMTU7+9LE/l+h6hsjKzMmHskdrZQcESlnz80RHleWZ
BtTylq9xsrgHTKR9shLNHPzkcxD5E1KvzgXFPrMTSACsKTeFZAyR6R1o4N7Us8Ng
P+eEtUxKHERYA7/gJ8CDHcuyKwa1icFAIWg/maXPq0JCv0yTZnK70yZ9xWUXEBq5
aF4K9sHU2TCatsrssjfNmXVwxTAX9NJ659ZulDLLxgHrpQRJSzUpJ+mlQtFHi/00
st5iWHtPPQTbpptBFTEecvJNquta9XFjrt9zdJIpomqSihbdvL8bP17gvP5WwvqE
0ljrFsHxTXJIgpNlAfhmvFg2qhza6c5tnO0MJ6PtkZ4DaRc+3OL9KHb7N3q2nNwG
GATkX7HO5HVNSf9XohdqCfiODEex0DzsYc9oeCilai2Z3X5J9jbeinhxkYiXcM5f
r2654g1wzb83bmC/P347o+hdHihk4xei1WwSbfQI7N5kIMGuqBAKLYljTJCoZOb+
mF2C97aZfCxX6yiLK4gUQg2IZNe7mrANlnQIK8MM+pshlSWtGuWr8eNpM1rCGYwj
TL8yQ2ZtvJoxFTZ9Cxlz6yWoyVUYcR94zxRsGRREBotMmHfuSWGjqmVtN25+BwF6
ex4VG3SErqeQzEcsAVu9rwSgEQ3RljQU6DwkBIpUnfVB6i3MRw3vVaJjObdI+YEP
6sWGRL01pwsBquANR6aYjidV0TQ30duFJrt49GbW1zuC16Mm2isabfQ+Z90tC3bt
cyFf9FuRGedDYM4/5sOg3Ylp5PS17cRVC94ZSq9/nP4KWmXmCMnz+NN21RvyVNGh
7OvnTlWOP8C5jegaIo2qlSK4fbO/pKEKijzMstigebzvRz52UFXgcU562CCiostF
yonMzHOkf4umOZ0kV+KF3APnlpvXKxAWBoeQSJWMtrUDfL8k6hAs/QLUXk/n5asK
Lxk1OnGFCWE5KgQxI6sSkj2/pjljV6vptfM2MjSAWVqfbDSh/bWBUu++1jqXcKBh
DznUComGZLowWq12tN/oBnYhc+127tzTOwZPOxekf+UubMw/lifMRYsktd8vv1Rn
ZktZPijl57vodt33hqKUJsretmh9CeCtkVN99hZP5iGqoeAMGb+zfrC+cXrF/ldu
yptFFweNnaqrk7oN0EZ9Awq4Zj0zkR+nBhAVEG9YEtH21mGQtj9aGjzNwrn3ltg2
i9rFrG1ezaB0UNoYSWcFPzubUEFbj+hVMH2c5gIauhZ1VLTJoL1rSmE05Lbhuhsc
2D8NZ8UpK4CxpV7lFkjCAJP/4xDRDARVmMqWUpjcCnKTqyJ4uIagn/hUG9gSz0UX
2b+M4Nhfi6COGKxwH55qkTQ7N0E6wAqUwVvSdAEuJzf1jWSUCLsCVWd7WmzLUfcz
LaIDwgvZLMY3nKgOdRv2/1wSfUUepSJzSpQp5ENjRSQLuYJTMDDAJ6eybh8dAnX/
O+WaD914S8A0lmAgDZ6ZFqAGNAEq+9vjK8MVs8RjhecV6x+WoAmuEv3SQmH7zk7F
gt9Pkx7N9nZMu/HIlO7L9IKvRQ4tQAVtXw4kUADDpC14bMO+/hkjWLCIYnJoxl8/
Is95J0AuXrc1yeOiNXASfxUAwPwwTz8gq9rXGomR2LrLxF/o1fHtXZoZW2r5Q3pt
hcX+nNcCXk2+v0RLSA/3dA==
//pragma protect end_data_block
//pragma protect digest_block
2iq65udwsDHJ6AvKDpd9g5yQAHM=
//pragma protect end_digest_block
//pragma protect end_protected
  `endif // GUARD_SVT_AXI_TRANSACTION_SV
