
`ifndef GUARD_SVT_AHB_MASTER_COMMON_SV
`define GUARD_SVT_AHB_MASTER_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_master_monitor;
typedef class svt_ahb_master;  

`define SVT_AHB_MASTER_COMMON_SETUP_REBUILD_XACT(curr_xact,resp_type) \
if ((rebuild_tracking_xact == null) && \
    (monitor_mp.ahb_monitor_cb.hresp == resp_type)) begin \
  svt_ahb_master_transaction new_xact = new(); \
  rebuild_tracking_xact = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact.is_trace_enabled = 1; \
  curr_xact = new_xact; \
end

class svt_ahb_master_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                             type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_master_monitor master_monitor;
  
  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to master common parameterized with master monitor, master transaction.
  // For UVM, it is available in the base class ahb_common.
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_master_monitor, svt_ahb_master_transaction) item_observed_port;
`endif

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Monitor VIP modport */
  protected MONITOR_MP monitor_mp;

  /** Debug VIP modport */
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_master_configuration cfg;

  /** Reference to the address phase active transaction */
  protected svt_ahb_master_transaction active_addr_phase_xact;

  /** Reference to the data phase active transaction */
  protected svt_ahb_master_transaction active_data_phase_xact;

  /** Reference to the current active split/retry/rebuild on error/ebt due to loss of grant transaction */
  protected svt_ahb_master_transaction rebuild_tracking_xact;

  /** Drive data process used for handshaking between phases  */
  protected process sample_common_proc;

  /**
   * Flag that is set during the first cycle of an error response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_error_resp;

   /**
   * Flag that is set during the first cycle of a RETRY response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_retry_resp;

  /**
   * Flag that is set during the first cycle of a SPLIT response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_split_resp;

  /**
   * Flag that is set during the first cycle of a XFAIL response.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit first_cycle_xfail_resp;

  /**
   * Used as a flag to initiate the zero cycle OKAY response.  The value of the string
   * represents the cause for the zero cycle OKAY check to be initiated.
   */
  protected string check_zero_cycle_okay = "";
  
  /**
   * Flag indicating if a rebuild using SINGLE is pending.
   */
   bit has_rebuild_single = 0;

  /**
   * Flag indicating not to call the transaction ended callback.
   */
   bit drop_xact;
 
  /**
   * Enum which indicates the location of beat address with respect to WRAP
   * boundary.
   */
  protected svt_ahb_transaction::beat_addr_wrt_wrap_boundary_enum beat_addr_wrt_wrap_boundary = svt_ahb_transaction::ADDRESS_STATUS_INITIAL;

  /**
   * This flag is used to indicate that rebuild is required using wrap boundary
   * as the starting address.
   */
  protected bit rebuild_using_wrap_boundary_as_start_addr = 0;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;
  
  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** Indicates if the HREADY got determined HIGH during BUSY. Means that beat_ended
   *  callback corresponding to previous address beat has been called. So using this we
   *  can aviod the beat_ended callback getting called again for the same beat during 
   *  the BUSY or even during the SEQ trans type of next beat
   */
  protected bit first_busy_cycle; 

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;

  /** Event triggered when a transaction that needs to be rebuilt starts the last beat. */
  event rebuilt_last_beat;
  
  /** Event triggered when read data is successfully sampled. */
  event sampled_read_data;

  /** Event triggered when response is successfully sampled. */
  event sampled_response;

  /** This variable is used to store the beat data value once it is sampled */
  logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]      sampled_beat_data;

  /** This variable is used to store beat number once it is sampled */
  int sampled_beat_num;

  /** This variable is used to store address value during write once it is
   * sampled */
   logic [(`SVT_AHB_MAX_ADDR_WIDTH - 1):0]    sampled_haddr;


  /** Event indicating that bus ownership flags are updated */
  //event updated_bus_ownership_flags;

  /** Indicates if I am the current hmaster */
  //bit   curr_hmaster_is_me = 0;
  
  /** Indicates if I am the previous hmaster */
  //bit   prev_hmaster_is_me = 0;
  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GNuSa84w/Uby1gj1QsY84H3foeHvlePoyk9XDJCy5N1JJhzTf4fjinN4mRgkl9Ap
j5XI842GGMizuZ/hF+6X1b7BvZSZP1a9+KNjB0UKZd1FTaARl92Gg4aaLjy4E6fX
blXfeQgt70m8/G2jy1zQ2e8nfsBnd1j1glMunXXIlH1Tpp7Nrd1QNA==
//pragma protect end_key_block
//pragma protect digest_block
0q9Q3wAlQ9y4Vgu6ADWQcWviD14=
//pragma protect end_digest_block
//pragma protect data_block
lhWQA8R9BPIgFGo59eTUqaacT17kWU5hwIuU3THP7aCIV+liv+gSxRmmIPYydktB
mmzk/aFF9/HBloqUbdYJXJRZo9k1TAG7f99tyKxeR0xNPt6gf9GW2zIbIng8qDVP
qz1S6E9PF3CwWPhD90X4JYXH2cbeD1Wnndrc/14wDqcwCFGg0amnBFQ+hoLzM6j8
TGYuQqxgayUGJlKex8BXFWqALIQst6dzZWUc058mprOg3z3pV6aH776fnzyJtrH+
e6Fyr25gSGgHxmjijABPFOnXCHO9AI2qBCtVPVFyZSSp0QJdSyhqbYan3WDQgmI1
jLTr/HFW3p2aHgwCUTENik2EPt7VZecNlLOZcxrz+Fa3diWJq5OH3b6zHCIiBqY4
5NOTQE39+79tfrTlFTelnh52NQ0hcIyOS6HmLaiqCBW2VO4VcwE657D4qGUvcnVS
ESG/Rb+ELbA2eBnQuZUwgZwAWs6wK11JhLyGNVyptkfFAUVhTMkY7blVa0bEcNyO
ps2n1i03DU5lYYEAmo69Es/ZwFlsM8zV80vyQFVmkXOLl2D3yvyE7en0FMdOHXCK
kfbiftIeXettVtgbyGwnz/xG5yy7EILQvoewhcXCFXNVCVJRBjqiRAOapGp8DGCt
SeaEckua4KSDGHeW0xRWLMEWkGFoeAPxraoJdUQ79MOoEJpKsb3ilDK6PBVoKOwl
CnFBEnoBp+ktrPfqQq+9eIguPxxGaJM0plopPT/qrcKTJjaEUJ7QoFecBGn2ddpe
+kNpZd1SIIz2npMKzLIXJZAqqDi1ciWFF7w21lmkBG3BQT/TP5WjLjVvc9JpXnFb
oUofb7wEVn/nLrDfPl6hxQ==
//pragma protect end_data_block
//pragma protect digest_block
d2/7NzB/qkmN2f6E5goFpV2TwKc=
//pragma protect end_digest_block
//pragma protect end_protected
  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Issues beat ended callback for active and passive master */
  extern virtual task issue_beat_ended_callback(svt_ahb_master_transaction xact);  

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Update flags when reset is detected */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Monitor the data phase signals
   *
   * This method only monitors the data phase signals that are common between the driver
   * and the monitor (only the read data bus).  The driver (svt_ahb_master_active_common)
   * maintains the write data if the VIP is in active mode, and the monitor
   * (svt_ahb_master_passive_common) maintains the write data if in passive mode.
   */
  extern virtual task sample_common();

  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_master_transaction xact, int completed_beats);

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * Transmit response to transaction.
   */
  extern virtual task send_response(svt_ahb_master_transaction xact);
`endif

  /**
   * Executes the steps necessary to complete the transaction:
   *   - Triggers the TX_ENDED event
   *   - Updates the data phase status property
   *   - Calls method svt_end_tr to update the transaction events
   *   - Executes callbacks associated with a transaction ending
   *   - Places the transaction in the item_observed analysis port
   *   .
   * 
   * @param xact Transaction which is ended
   * @param xact_rebuild_in_progress Indicates if this method is called during rebuild process
   */
  extern virtual task complete_transaction(svt_ahb_master_transaction xact, bit xact_rebuild_in_progress = 0);

  /** Creates the transaction timer */
  extern virtual function svt_timer create_xact_timer();

  /** Tracks transaction end */
  extern virtual task track_transaction_timeout(svt_ahb_transaction xact);

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** Indicates if it is required to abort without rebuilding on retry response 
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function bit is_rebuild_on_retry(svt_ahb_master_transaction curr_xact);

  /** 
   *  Returns number of retry responses received for the given transaction
   *  @param curr_xact current transaction handle under context
   */
  extern virtual function int num_retry_responses_received(svt_ahb_master_transaction curr_xact);
  
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * Map a single AHB transaction to a corresponding PV-annotated TLM GP transaction
   */
  extern virtual function uvm_tlm_generic_payload map_ahb_to_tlm_gp(svt_ahb_master_transaction ahb);
`endif

//***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
rb8dqYyExqpOv1G7EjvBTDjSruYsdPJ+A7X8ukAS2tAoT049xWNaNjZQFaT872Gz
eFGmKMT0Ec9ZFrUUrI+xwG7HTCfZodftUsYDsABRtw7TA+9T3RokJuMxl5NXn0eu
VeXyrvAbRxBxBw/XxpIemnB0fxnV/fbMqUqYsMAe6GU8EFN0Cj0qhQ==
//pragma protect end_key_block
//pragma protect digest_block
mOVWbaaaWzcVshR40Kf08q1YHxg=
//pragma protect end_digest_block
//pragma protect data_block
UwipQONrwfYWQX2346hs8Ojj8pvVYcQmTtxS5TKfgpJGLNNvtssrPoH8IG+Hts/A
QIVjxmWrnRwbXpK5nZYmMyBLEZzca+oEKn9hxTVfpJEovSA9B7tIvROpHTuNlL8b
CpsuyD9CJjpan3fQlu5qrxJ3ejal/DujLuXMNHaxCKm03xYjyi0uKgBGegMUeUgw
Y/os0cKaCuQ74+mGn49MkIHOGTwCNkiFR1svnh4Git5hCQt5PrcWwK93VpKH2VZP
VHtgKQzSX/EYuXZT+GB9Kt9wNkn/W/uUmdfWfIBK26qtNzFTEGM0JAMHwBFTMpu+
85bqulOgRJikpcUPc9PSAv6m/ZiUzo2LkHmQm74pNGZRIbnqBoPHGpU9MKHzq50v
I1D5wjWtX1pXQ7+MqPwe7UkPMsOffXPGzrFuzGEqY0azGBDHFiMUpJS3e0uVjhFB
B7BjRVmuvg0r8KKmaflZlDRaGZgDjPO2Vj4F/lYutTgsr7s4EeiZWInB1mLIqd/A
uI37lni3hnsBNp/+CHYDcK396hA5zjDb9LCrfmla64GuO/gAjQe+Ky4uzDDy3kK4
ucLGyjeBHAojoTishL5OgRUrrNKTxOtHLyPqWkY0fpgQ7DFd9XhghSdcm0/vWykr
hRynXAw6YLle8IfeS0cR8gsY2I9sicsIOgfcvqkzpbDUuf+Xe5mi7RiDu5s1fYLM
lv6mVsVYtQz9LiwYyMP795tgkhuK8i3B+WCAL3VERS11ihBgWQJkjz6gM6snRHf1
xvBS7H3rgOKzhsKM6mOanDIKCMgn01T+jpv2PALLWNVLN4rK0Guib/1vC6PWITHQ
fWNxVURRG1PAJGW03F8cTaW0qEvpdUjSfFMA53qys7TOUfTFstx3DHRq0l7pG0EV
mI2x5f9Ck/l5UnOaJA0krs3ImK8j6h2ozuhDySLlT6QjlQRZW0VCjSPay05zxWuX
qHhuVBLK4K5/ngvzS48W1/EGDVGMPrp9PDhSJBjuo9OUKp7GJQMWDvFBjYlCqY25
JU7A9XTxPKiGLyvATNCQMxqNGmGctLmG/x8n5OyRqAXL1iPEwVQH/ymp3sSOH3OF
MyC3OpsKnoc5byYfjHV1KU6P246SXg8cgZ3kXhBX2/GtlbQi8rVTD/fSI362Lp3Q
zNPnNDLD7/hVJo/qa1l/F3SYtOxFI8HhuttvYypWrXWEQO/F74/bEAqkOM+U+ch2
uUwqqhgRmJZP3cKdZFOGUmmAuixyHluwpIim+NgUtWTajGx91dEQ1gyB1O4HQ06t
D8kLYG7I8dUGCpbel2y6fXhoBzf6AlU4fboBXIglycyTlnUWRM0quptiO/UTDAAx
0wC5z47dNay+jquUl4m5FtbvvE2NW/zawDQGpxOtWCzJWbL5utPHBJpM7UNS5faN
wri7D5B06wPaQzziAOYUHatXH68RXRbvM6DXNUqd79rNkklYaXriDMlus2AdpSte
ZMRc4772gfDpCzX9oD9Q2TfFzSVNbmtUapCJoavprMCVNE/Xn30Yb9p4xTH/7H/x
Z/oTBsTW6O2H/Ij00WOBbczx644HDPaDe2vGT4/uXP7QHKV5+9V9hHKDdPE0iRt0
P/yxBOLqORKFhZORnECRK/UuZQxu9sGqwt7AJWI1bt5Ah0BEW8YgXjBqIIj7O4WU
Wof5iNxmzdiPK9IcbD7DRJY5QzqDa5+0FUIrdhsP+KEjqrLnPhWVbERvvtZYDZHa
ADDIWNrc1rKXle2CcqOCUlf0MOZzrFEkshd8cks03vtPmACDweBf8cthJS6Lt7oU
2XsX2Ed3s9EsyJmRx61ThYeKIrqQlwuCzvwM0bGwn9IorQdSx396sTLRferueQdz
mbJt07/OKj0j0N15KVX1rh/v6mhBs4QtPnpcTrCu1aYX+frLXfh+DGO29IDJ0Nt+
LjFmixEcDHN89e/EibIfW1ELzLQIogHS21FZW0zZ4r5ZElPL9+jxxNLdu4nO8Inx
aYKUhP4fmOmt4QjMiU6RiUaVUYGATM2iHrc46pAbrrVxsuvvWBL3CRTySzpQAINr
ZzCv7tL1M9zrVLs0jjjmdtqZUYgZ2Z5F0R30/4o0tArGTdpTRP3WHwJcJUz8Gf/0
c0ObBIzYZqxJTYkt19K58wtNOPRH+1RRsjX36vShJeJWZ4eyLSqUEsR9Nc4nkwht

//pragma protect end_data_block
//pragma protect digest_block
I9dFl77XCyj+MSvBc45+zTpZTCs=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ot2HjQRzC3E8UW9uV9QiELgBn1NzWOPQ5U7CMJo1ozfo6oS7+LqfaS+WV/zw8k3t
G8U3Ilmm29cM88TvIS0KmsnxV8OK6h3/vk2Nx4Oqfa5NZrqLr6uh1HMj8WEklpnr
WIyBW1Lw/m5+SY5i/cta4ONY2WuU5itc6a7J6SknftXFTz47H2FNWQ==
//pragma protect end_key_block
//pragma protect digest_block
Ghcy+g/UYrSSfnW9AcArcAEZPWM=
//pragma protect end_digest_block
//pragma protect data_block
BAJdrBBsJG+cj84OXPcNy/fv5TgXMo2lGquISDCVb4Q1gRs4EVXo9D2wwKnA8qap
GoEGxf8CDLOhN5tYYxKzoSm5Q02IinaJhZ892bAX22SvDH9pajUwNQR1kPtWJ5lJ
TpWfFgJzzoEm7WTtAz3igW/pZtubSP9tQ0+0hyUWGEZI3dmM5BLk/epL0RJsrFvU
RXTqAewoGlQ01qspCWwSheRcm5EGmh43IbYXx64pMluvabd41ovWqayJevijlhwz
qr/r/20Xd/V4xYPQ+b9bl3mNu3QB4hKACXw8bemB4ikK+AWypE1NTRXgInGz3FnZ
NAvnwle2zFn1FYOxXTCErpK3CiXOG+H9rXjtHbEmDd83+TIawSW1KYWzlsQEz0sj
eiHodL7YDjl22W/QZfopsptH5JPcHVxRui7pCKISGHgnwu4w6OerEMVyqt7pgsiP
lgsXzSI70UcqETvznin+u3of+0mjvWXXFVhx6qcrtKBq65BViXtsK4gT58C+ewHl
n599a83DpLqyLYguXga319EWmBTt/hT527xey3bHGzb22wdJKDJN7281uzBxa/ZB
QVlVuiawk//EPAjOF/509ROiXKSpkXDdyFNF2S/5MfWiIjBKgI9yMehbvBFx3sFv
1TZENy0XhAhhKkQmLoOuTLxtUYj3zJdFHYAhEqRmcIXEw5DdMLJ//rrrYX/kmiPo
UxMB5ILcGzQq0d4l4z7TTSz5rDrvB95QCpYqOpGZGOZxPMYqoN/C415fxvG+QeNa
QeuyPr1xheueevwbWLbxXPOYiyb5KxZyygeip06GxzUQeyCQW8tD+u/pHSofWD5N
Wr4hhihfok2cZkoL/d4Q0OXlaxdDJDC6aK1361cQQIPKVd5bunI96B1Lgg1SsREJ
/dN/8KREdId4n3kqhK8sXiRHJauIPs7gd72UoCT/CIVitrjWjbYFh4E5fF31yJ8B
MXZer9/oG4iAm/dnyuQGfSKGEwke4n/BPON/Z9GtBEV0U53nbWvT7QR6LNR6nZwK
MtRczR6YHmAN5T5gQO9xgPvIZuR7uAsFs/bCY1E3X1TjpCQWuR6SYRZpfao6KVxt
AjPtOm279rlzfy2IdgPhTu22ADSxyfnIBzcyCAYBYJ7cY9mK4LcNnVepedxEfJMJ
ap2RMrx2JDKW7Gc/+azxa5//GMS+Jb5vCw+rp+bvmQu2urz1W872Sf4GHrBeYtQp
i/3zAqY6epzQ5eLUeJXmeTzmgx0jfeuKi7fvKs24ivdTOZorvQMXucBRE2jBZdpq
mufvceDPT43Pt0DUr9/FgOSVdApnYLaF1qInDb/tLadi2UWT45S4dnC/YSV9Rf7j
O7n7HRNzfEgi2cSLtACCKlDgWQ5PoWqKUdDz/KLtUayqSJmNVqwA6JREBQJgk/42
BUtuIw9FJR6CePmcHLS/F9Xnc2IKSQRcGCaRJMr+ysYAqE3hh/WKCRNgdrZVEL50
VZZzPnd56c+DvRg5g+Vpq7I0WZacnuOuI76jNx6AyvCDD2vYi8zaIuXpyXVTNxw2
XOqSD9/vuJGDW46ji23oOLhgU+chdzGGyQXkeWk5QopQ/HD2GzcTKVS1gmyK2WcJ
NGdXZEoElH9idhWjvjrO8QDr/v35Kwa1Pxs76BcmGmZBNB3XNp3POBnqbBeevoz/
WcGBuMhG00fp7LsxKAEY1+Csa3eg4ucDC7YSxVEAwkLkl2Ilxrnu7UX5fQhcde19
m5ejnGZZah9/Th0oIxGIk7OktgnM1GEsXb2rZez753xIyREGGlRkogR2fcwS8439
p6urk4C7PJUnR0/ilQXGLnKK+5VNhC0IfYUT04HJYNaA99RkhKt+gCqYwj9IZ6Kl
jYHx3PMO2zBBIkJwnGAqI2BLKjv1aXbCUGe+v/GCvRYSOVZ9YeLkeCnH3K63dT0x
BxRxXhdOGOYIUSGHkgUq9rEt9wXW1oYrYZ1t/1s/Gn76RyotcvlRNPQ6hagQVA7y
+SwmmuXRNJD+y0ziesGA013QgAtwkYvk7E9UPO8E7LBytuci6ZMHuo6G8JnTQ0fb
i/DOXzLs69LcowV1jNSzr7vOmWlNyl9XBMhCnpbFhgIon8KQZrigPMF3Q5lqMnGT
G0K7WW+T8wfRbc87KUnXUskh7oWujZoehb6DYSnNouv5gW5wFZtGzaPbBt8oFC6Y
eXqHiTsv+VaFExR57hENf2Ll2eBKDVQ7RKhIS3FPhyRq/hjskd7b6nE67cyNfQPI
dIeJOg3h9r3kMZV51Cj7vOv0KGHWez/ll4ywXGKlRs2crzsheID9Gh3qNadOE6Ec
mKKzpPgN+WS4ab7QrnHQ+/jsDhRLDMjFwuASSnaC3LX1AvbDX8F6rul9CXISTu8T
DtC2AU5zMOcGfS2a438WVwhbS7Bc6c3LWYbve4uOv/3VcsiI25HLsRfKtU53L6O2
4hd08cXhoA0f7cv2NNre749YExpC6qsYEYKa7J1tlDJbSsErN7qxbGDK9VDx0qoK
q/swfxO4l+SB8+wif/gPOU6tDSAuX+JkIQg9dR+9Btj4dDsG0yXPgqdX4mcQqW8D
hgcLAtDia9eS6Uk8MmacPHIiE33wlI1/GEPtzcFx7iS9Es+LiXXMkzII1BrE0F4u
NRoano1I57xWYqmgY8nFVxM+SKVZYw9EnDbl0qqiI8LGviF9TThCndLzpfBR0uSA
xh8WjsUfWgtT7KVDxSmAEMSk3+G6GsD3AmLJxrGVOY1tPXwqkxTEB2I7kDnQFvGV
mI9xGRCuGrVOQ9J7YFiGs6r+ZdX7sPk9nuIdW/xjOe9CQHkfkkUkq23mFshUwNvJ
nVh6/R6DYe8c6sgs6Z0haQ2JNg15MpmxMKhLQwYcvnZg30xJCxFR3aAJOkYMBLpR
xL/B9tj1OWRsBdoucyVAJTjdlaMx1WuAXTvAptzEI6gqJw/LNp5fHD3EHWmzf5RL
hDqBzta+dHb48CDyyP/+TJJADEhYAl8mPr/25zghdqDhCkxX2+wvG2sb9PQWofAN
Gd5JmKwQBNpnv1/A5RXCKAReZze7X4YiYRb0GPSvOe//GimnrojSe5i2nPnUUG9J
CBegKM02GWCqrf+Iz4WI5ikk3ojt5X0YN6cSOkwkggt/YmcgHiBI7I70h/5fR3Z3
SaOASbs2TPOkHsNOxuOj8FmoViUH2Gqq9iBCN7xWvxtEmKtpAopDYXwL+5QWE2PH
TN4nB2zO82Nh7MRLFceeGd5gLumK26sUhVD2KvOgovU4b8h0geFOpXVBMHzxkp2w
y4WCAXe5lBfZ5KoQAEEKTP8IFj2fMJp/gDnoXgezPUXOCoKH4ioealWcqt3r0Hlw
JpfEh8EXj8OKc14Hdzm7nt+WrcOXlfttJU2xL6Wt4lar+Md+gqoQoqyb4138SNyD
SK26xc+6JWUPk/aY3JKAi/VQln6csIzt0jogQ8j3InUeV+8k2ivyDgRoGsfXnymt
JtgcuzByDzT2SkQs3wtkCgmSOeqAInqgkTGX3jGKuPH3dvUQB2o83f4ZGh0+5u6M
4D8xtq3HE1FzFsZWwiJRV7hmGZQtH8XoNpNiqzIi/KzPE8jDE2l1oklsNc9GDbo9
NmGHBaSs+fOx06g0X6MMzOOvy1f7N80YJsdtnPvDprsSzKIIoIlVwiEn0t5bKTGg
dyWzkdui4MsNsxYKE7hH5MCJA+qYj7LrtQENPalTQpig+0JP9/CfdWJM3byvZ2E2
7HPSSojtySEKnNqwlOoLmFl19ZJj4sbBRPICq6aJi6q1CvAZnbTYGdgrW+j3NpaE
x2dhdiGoPQhJTbMQ+I1J1m6mQJ08gdq1NJK2LVkqomx7QhHrBenmVtwgjxmUCKrs
dzAz8YB+o7xscSKVkUGyGSgXRPeuKOuMBcIuOyIVXCbvwK+yRY+snvYS5QRaJplu
xbpHHT2aPHXP6q4kknO0w0KUDC4r63hgBFDF2tb3j8V7riC0ON1QgVBYjevTdy67
6QhGeFKYArw2g1f37S0EezT0QKURnVpySXVc4Qa02U564u7QPuyuM4YQ12uq2TCU
BM8dm4N4WRgl1EsV7mSzIJhMy9Iyd/7ecHseJGveGEe6oE5PS01qBCcZnbpHH/JX
+ZhSYEOJvCnXmZgVbm7zoqSVE6HsSj+3YhV5pIqL6W3C1jrSYN+YDdzhvBgxiq2U
/kjcXmoifZjPG0wHdGBoTfpFThkJKM4/ThimPVO/vUEQCv6tqrtSXVIcskqu0PY1
spjJKRAVEYNWDKLII8n2KaR8b097Bz6Oma30ZQxbB9Ck6AGjSwm/EeoZC0yPRXA6
FAH3+u2AGSK7ebq3PS/GRjU4Fo00hQRvmNUNETFfdqVgN/qCxAuYgbE5QrFQpu1A
0RWDzIU8MEdOkAda/topJzpyNqietgZ8PffWayS7TJ0JKiXukeHWDsDVXK5xqAcE
tKVUx2JoO14vvGo4jEK8JJkQu3Ut/dkcY+ish0o0vsnS8wdf1v7YDNN6VfIGAaAu
j0nLh4tmWeUC+zq2Es8jS7LOqUyecafadgLzOAikAorO1+/MHEs6zOx1wEFNBK6s
PUZv00tNtcygJXsvqCwVF11O9GYLlmWAmr7OJU+lymUhaWqh4YdUxOMw8zFx96D+
jVNNj73mR3QjprO3c9X4hmxcc2+bdKgcHkKGiA+j6ZzVEusc++wGjp5SAE9wCY60
vUZngt9Ehpt/bL/fAZnaa/P7rn7mKoWAZhXfSLw7XaV7e8deLYN2LhmR9lHAuyrh
cK3ZSGJXaqPZJ6MS+THvlCGdCcDINQvgq9+qzAzGVbts0xUZWTDPsYM32rE2MGO7
2HcHNH48Kth7oE3SOziy9phAvngoJ2iaDbIEKUURmPcTru88+CWX4TKPY5uD+ltw
GhbAjNAp/rdFJs7sNNKt9MbGqKCXhirppLH0YK4za+jO7uDYXhF2Uc0ssk6vRRIH
TEO5xkCc4iQeVb/TVTHcNqjGCLP6uo6Ub+wPRFdYtCU1E5vlfYlkvao6RvP1/NB/
kFqtso28FpJl4Thxqt7+/QUgcTjuYrO+Gb+JGchS3Z6l4Mybf+LxXPNltZJd3SnF
R+wKSrBz9cv9dEuSNyl5OwDbRAAD6IQ0A9yMujZuQkmv23TZfhpPSf8LVnHcFcAP
3TKcvNnrDfmyyoWUhl41fp6TuVuoKLGlU9j7fQkdO/qVc1UcMRQXeEnDEANCO8qt
y9KcIrUeT43UB5fbWs3WaYlt2dGy2Fo8XbaoYq1gtZ68RlphuNPXlj7NO1M36+vg
WQ9LNtEMQ/BkDhEbn2efU9vTJvHWKyVc9sIl6asnAWEMGKjhGzHUuM1en6S4cJTx
E8KddHVzGTgXez3AvJhj0TnFyJY7OOvjZiuYcqyMuR3fthBbZI2ccYltVphDgN+9
b1khEQszqeJ8DGuDA0EKC+ZvBtgaEfMkeE5cYamgFKKhG56VDQmeaQn7yz577XQy
3o1qR4yVwiXXdwPFkKJYAQH98MVqZxH6ZvExZdgXo+G2YZB7r3T3YYGwNCTZNyZN
J4LnC8cFbbqJNNM1ZjGZRJ+vdyNvfPx2WNd04BCyylwHnn/27mlrbTn4GM36HxEm
SMLbMrBkRYfe0zaq/3fDhTrYATLxoLwFThdJ3YjFSVF8IxBr0FD0kTaj34y9NSaQ
hmBqsHyZ4wzLWepQ8qiA2btNZReqzi8Pozx87/w12KUaxbU8C0WzJZyBB+LwlATE
q5X7zDytneCx2KHFT17RX2y9g72c6/afdoRawf7T4y7lyzTbfljVr5FqkA6e9T77
cq+UF/+85gvD1APgviV3m4pCVurRcezjNohp0Zm81IL2bSt9ZvKvR3XerhkxjAPB
TM8jPvoS2s7JUFdVH0GQp67RkzQ7Vm9cQTb+VP8xX+0dc+39ht7/jJgRtyGX8keU
tG9h6BAwFbj1sbw3hbnS65lvV0VPsb1AB2URGKgLU5Q0gIvLi92Ocd0LiJACQ16x
WlIE9ket5eKdQ36N6mlnKao8kf0x5Fot1hqLBwU91LCaFL+UTQ/OoxKG4ml5JzqF
DR/EawV+KGhGC5m5pgnBMpjgm9HmyUvOGjTr6f/1zrnVNAkQ6WoNw1NdhJ/wUtjY
gtzZZe6XPdPqto3hdbSgD7yMe2mdiiQ7/7SNnPznX65qQ85KavTDIzHMFlova/sK
UNjXbYJG+i3OILbi1oI8PJFm8plvy1OTQ5zhEUTQu46369pqJf/gt2k8p3TAh0iv
oNcxaoIyJ01YSvIzxbV70YVKh0UCKefGbFR8tXlubljNpHs56l3xH6GsEDkcd6bD
B6M0NnmBI0cq+dsTkaZFb/b0XWGgVGaRgv7VYHDOr8J7S0D/zZPffFmPT88UYmcB
XaBjAMopN/OjspUeQPcJMKgJloyRRI92a+6+lONdenrgw7RGTeUyr6c01Isa+ED8
MGdCPdUF8IsF6Q9zF245ZAIb3zmOdnPA1FELnNWRK3PmMHumqUNtQfash8ds70ac
At4InEcbrqsnB4ULtX9t/XkCX4dKlCmypZmJ+VWyL28WY/N74hqHGAicdF0IHGIf
GBjK7Hp8qLBJ15fIZvAe69O1n0mre8DSrlyKmRVn7+Z5F5Gapnsxdq4aBkxhxS0y
TUqpZzhDkb3BwrxxKuOP+MCQ9L3QuyWoOk/hcJboK3TXCMA7si+Velny5KdCIfmL
126p6nB4vF3muQoIcYAHQSdnnBg+TnM8oIQ5gqgYCrLSMEVzNRqn25kwp5E8CEEX
e9LQcM7hBhuwpB7G00mOqpjzN/0Ga3xeyl1Cg7HQ8bYvC2dqV88aPj1T9mYChYET
jACy0nO/1bMjmQ0saAq4yHf+r5M9pbP+1INhDmrmU6HGWv01ZCGR95W20H7YHw5a
vjmElDVYsVII+tRDgv0e0075sBJKm16FzwiD9O0ONavUpQ7ZEKGFdesM8NuszHmQ
ZSiqU64GI/zA/6CnRnnphDl0SvCxqNwEYTIXNHjwYPZA2fYnNfvRbBB9KFdUAELo
9Jtu/XMZtnS4D1yuEwKxKJbO8Zhq/woOv7jKTvhmh+WUkLEhPaLwt+oLarwwrrLx
EosW5wykxKrmOZvvy/LHbBVa0E/F+2wfWhWXntVJ2+XG5Gvcvp+k3NnWcQznVcJA
BJCMN6igQG0aXgbRN0Bievgq1cl7xNcyG7/saCxXapZLidjKT04lgrjTmDi+/aAV
oxY/jrQOLYi4W47NirMeispZyu/EtfB3JwsQ8TwjpAyFumv95VOFgRp20saaXlSL
oWmeRbXIEXUpYxBZXz/14h9rHB5byQnLp4dRnN4bHJM8pchsMBb25WKjL4coXn/n
p4otoeu6FtSR39KuNrK4URbt1fy9FZ7641GPTTMRBny4UBwk/MtozmE+UqSQ4Hx8
5O8P2YUG2UVdNpLV4Ij8WIinHSae94dgdmM1/8XeewXjVKW8cImnUrt2Ok3sArFj
aN3OFpr/drTqdnCyuhNiY5h818cqLHfSFV08fZt7h+ZJUHWkUL5ItPOr3jrGz+in
xGSBcDw9X6BgR1TkiXZD0T2xrNsead4fXE4Jr/R/xzsNWwWb1gwB4Yr/5It0GMt0
lDHbnEDgoI6SBAAdW5lP86CGfrykWDb6F9npHDsR6SHfY7Ou3fZrK83jyFZVF4cL
UHidHgHAsDYxAZcquiojIGorCoFx+C1b489wF/b3KpMSZR0GyacSdObMxMqUXW4/
VyKljOKQe1lF2zaN3NqhaMOK9h+CG6wInGiGBCcnrWQDdkMqmP1JXsm1x7Px3ZgU
/uZ2K5tFpNwpiWs7mAzqeIvULUQWZ3p//hana2F2yqb9/8mjxBP10k/OgFBxYk72
d5TMLCg9jfitkeCcWe5BtQAmTDkiYr6tyTkNFV7XfqmIujBN7k9IbUGvVU2s69vU
5AZLcfIy3Zn3ROtbYObud5crKP5a7TB1aW5toXnlTiHLwK/W4mlK/aIHPxclOoOR
S0wNNx5yVrEpg4qRcowdRv8bW3XqfTDeCsFie1zuzCgQhC2fWMyYPnYW9/Xh9WBZ
u4s1ZUAnOWkf0Xf1B8ISYfM4Bv5SmG0bqfFCUow636g=
//pragma protect end_data_block
//pragma protect digest_block
xRrS6bVzl/3yxPgVVsbfzBbQtsA=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Ak3It3hS6LnmV6ameGROQ2eYCPCMf9FGasBeUVyrQwWfSp3IMj3II+s0DjDx90Aq
JGw5xaQQvhzsboC01/ntU5E1RqpmxoN+yTwlNZT8TouhMv5TaIVQZyTVRGK5uQv9
6PpWvYwu1mti7T8ip8Sp6rBKVY4mpT5xpgmhSIGGO7S5bRM0gSBHiQ==
//pragma protect end_key_block
//pragma protect digest_block
C0nhojjhe8zVXzfMZsLd5kaeQ6Y=
//pragma protect end_digest_block
//pragma protect data_block
v6vX9oLo20t9/1/UC1XJPVGh/i+SSYUjaZi8/796XRCb/vpSXWof2M+4V3xgBRRC
Z3MZLV4DQSHiSVoZvGqmPdiM2ow4+/FYLvFghLMraS4nXgT77YHEuEopQAwNLfek
OrzwM89hgfQsMFNxqSe11Sx/QMjjYsX64KBjum+alzrwtfAP96KswMu4N+fkVrKL
O7lr33DqQbU8FZJYgghDAu6vaFRB3Q6Wtf/5SLi4JSqIlc707CH3TF6uKnBKZo2+
g4Eb/z2m7qpFSYqGJEbclL1Qf0J6YpHV/cnYDiRwjALps3gDhqfL+K343rcSHogp
dEE0MVsJ+6dGrWVvgd2IdpMl4EQXopjVPgni8zPERqTumEOGTdUBR8ZMr9rF+e78
ZHt6a3jt5adV6FkLPtC+GQDRuiQHoafg4j4otfO+9zAdsfL/rpRhe7ub3E4EfzFA
+kFtWPKwjhIEMNOSwXq9kHz2xhd+oSkzBivZ9MHY/ZKNoWpfGAd7HlysVp5EmDGX
e6UAgrhyNkJZqq1dxHLcBVbZBV/PU/+i0md0yLLq/tEZmHXtrNaIJF1c1hL4N8rF
iRWEgQrKIvPWtjvTPqrgFSihshZniJKep0sYX4y57DuK/lEcQoI00m37OKk0B/G3
u9GHfUC0vUa1Sxvvm81bqPcXthve2c90jHiUiefTBGE2c46NG6GUKBRkTFyFTGzb
ZV8j0XZJzW6d62tSTBntoky89q9if/fZ02nGj0Uc0BP3/XU1DRUMd9WrA7h40Umx
chIrgAkBNDzL1yt9nM+jUvPwfnUB5Ej+oHwBai4BK83oLB/vCiOaUET45h8JeIQ+
6yUKAdRtri0WOZ46bTGXaoCAwuPiWCdYsGTDmPSWR8PfAzFEQ7+SJ9or6utDWOYG
va+rgj3nnC0XlnXJyGpmCxnJ1zaW+5PgDdmhqlPbSKTQafTgQTPEZqPCsmqCtnRu
GOhK0N3HgIUIhjg53TmTMpvjYIKj3gd/lKi56+fp9dNdicqNF3xBj8Bex2QSQzp9
u9O+2S0SIzvIyKIkD3lh8AMXYRSS56hUY6VCO/mSzdGthEKRSxymwIJ+Wt2wwXqH
2pGHiUQ9Soeat7M1bv7+t82Qy2lYOzH1Fwxi2PLsaQBaSG8n/eXH4+9tRpyyEu//
UgVT4PvuQ4hi0B0E2uTSwPVLeGPOrhL5Ud+6lH9+o3q87yLB8mcBk9KYosr5Y+75

//pragma protect end_data_block
//pragma protect digest_block
uUyKH1LEfTjc8QstNM87/KBbmo0=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+VISJOYqH34f80rVglhgFuozj1mf0zKo9rcGN3jASdMptWdLyU/71UCrkzi1YPrf
yVGYCv46BM4nKGQpmWrELjFOPw1TqlLnvbPlYKspa4iLwkVEx+hY/ABtnnQJUM5t
ze1btm86O77LzhM/ZnKvpkU9ecqVoHwjj0RYSPC9pF2Q7iCKTiOhOA==
//pragma protect end_key_block
//pragma protect digest_block
Q3/AGvn69RHWOBVzeNwzrN2Ud/w=
//pragma protect end_digest_block
//pragma protect data_block
OCxoX+AoPfqcolC4rsBQI7bcapR6aYUOujuZ4L3gukeHrQaMTJieYjR5WxMRrxn1
PBtwqD/KClZMYYrDxv2N6Tvxd3+xSnbJZ1IHCcniDzDT+JzsoYLpomRZZPCmiqjY
aatVwt65x0VJyD+H/n0V04vqo5AgUKm8Xwk60OXhTxef+tpk+XuBhOY86Y4qHL1c
njv1ywAE3y35/iNyQnF0QDHONSpfWpu69uyl+Jp/MPvgTzgnzv4UHcxZ2kCwZS4h
e/bzina2qKBY/W94Icob3b/bS8LL39a2T+nNMFKJYFbURGxtxPvqjGjXcZZ9byzd
2SavpUA9qiaVHCchni6+JY46mV6cIwjgujhLha6cR57Or3Ol7ZLphvVtZeigAlEk
x/a2dtPBxZt3/HRSJPDBZFlQyxxu8WSX7n7ba5yNdFvQVnPKLIKRhnUkkjDPcwup
JQ6NSeraPezqk6VdWQYggwkfeiNchxCiRCtt2uvYudVyC/WWX3BqrgKIlDCYjngq
NmdV3fv5l39gGZNKp90ixlSYfmWjw2lcKqdx69cNw3OBXx6+tHUEsCB4rKquuId3
Hmj04VRxrtps8WbQ3otyVOhIlBCXj8y66oOCpFYrBsDvDk12f8e3PFUqdyk3Popz
fKm0FZcges1a1Jy8seKxMI7snGEbar9hhYPkxYuA602ig1PjVu+42U+HjUMKtEoO
mRo9/buISsi/fGK92X6vizigdjHNFKubiXGEno4y1ZBR9uMq8ednZTRZjK5oMGQf
Q1f7dbRkvNqKOCjdnQvzJgSqTWm+d47xOMSkzSahGMa5CJGSUExhSAEykE4FqwSH
cvvsEQR4VnHQFJQ+raAcIeH4iK8ldGVpDoRQ5asFIwDk4K2nVneIKjBEWnJtsZmu
9AGNx1hOy3qzCMW1GIqpN1pMk7gNGvf4Akg0TmpbG2QTD8WMoKGjKxA4zctQtHp2
UjYO0CopGeh0Hg2qYEHDrTzdX8TuBc6+hbrT/gbaB8MvxFzm4VdhcJTWQYygvz18
LpD20vry8bfA6eDHqAUayV7T+Nt8y5DZ0NH8OymD2lJ8FzVT3Q8vVX936w2htq/7
WMO/WxgCQhqdbBh6AWtJwLQzGhK0i6G5E7lxfczenhS+Ai5N3vqwF39fiV3GjZ6s
UtDzHk6I8XA0jg7fsQ9vRFE3c8ngt1tmIRDpRlsDRGpJzO5qmRZVv5GveiSrjVdL
URou++0KhKrNArBocOcxhO6lCJ12AmAyUzE/Tcmx138rgFeX49JHRIP/d4jEfMqU
tax2o+wN163CRMQFnZUQGl0Wjv4HT5nTVH/BTfE86pIuti6fj5gqSzvubszRzVIr
iNCBB8G/1TybQ6NhLSrKer7avF6Zp+QF7ZI8kvTqEKPQqzKe9rsz4NSy4PP36s0V
3D1Tvs55xukEdXqKIEg9gy2c7g/iIAbIIOH0tFsOGHkJchmlKUCKe62JwMZqOWLO
NzKT3kDtT+Z1lHwrw4kDGMFLGzhs/lQq9KVtH2iWbj6Lx6e+Qc4TF/IGSX0VZIMO
LGr9+5ITN6Qc3KStMRMPPRGBMVhknyMEhluOMpSOQ1oZyLTNeom7NibIt6i8XsrF
ZvR4FZ7zG9JvLMIE5k6zw+50SRUq8hSwn0IxjGCLU9/abrXax/wDrI2MjyLspxwU
0CUYksnsza2JFilVAkq60dxtKaakGCLXI3mRw7iA3zvPJYtHy9mc5DDDnsrqZydz
+7cZ7y3jZkQCKjrjLuzQbEBaTIXsS/kqAXGDm8NIJ64KrWW2bpkniNqKL4hkuepZ
KK2G51n6qt81GFudP3GsFTbsdTmFJgoK7L7ntnyzBXsAKyH/f148SHnPEKYl/W/v
WqR9MntrvNIUmJ1UlddxHPvw9UAT9H8kk6Ze78TNZl3IQoTi25ANlqmEn9lNVvLX
y45NbJHRKeIk+Kgm3NeGyQb2wUiVrzOmKDSezYFfrVpCwrZ1rzAcaZ4IklUk82NK
PfmvUT7AISfs0RQTkOc8CZeLfaLszBBZ5GHj2EY6kRNYxam5IVvrc/w1b6HvYi0K
GF1PBhMhwu/OOsqwSdc9EM7zw2CHznO5OrXSrWPezxw0dHUmaCt9oxdVYlxR0FvA
9FcXXClflmAIkouIi72gfEJTzoiV3m1cadr9G9SUPcFeE5tpSRLGiwU7CjluH65X
PM/9zsqwOpKbNYnv+IrpYd2enYuOs/7mRIM5uTuEAOBFLfaknamoIsr+zPcbiQ1j
j0qK7EmADUg6b+My4UEgIcUYl4cWxB9FXJ4Qfe67R0i7vep/kU09+nxmlgYNoIce
MNlWsZF+xwcOjljzrL/GaKb/Bo+awJeuco/PX4c3c5v//4EluJlH6VDsUooai6YX
RI59Cg92APSiITGTF+69jbVAOalmzdts/WQgvq5ySmo/mY/TulEI+ALILUMFlxYq
rwZKuZpSTuSdqIJF2WkxP0qFAvxY3bqbPPdl5vmIz58f+RAUsWDSAu9th2phnRY1
SODA86onF+dxKyXn7XLm8Fs0G7FaWFTZqEwcgERnDL8TODacfqAZSGLL5EA14jyN
t3AjVQNJYniOR8WC8kWt6OA5RjoYgzEcb983lDp4lAanvBZtCBBRm925FyP+1jcO
/sR7JIZj624VoiI/Lji60yV04tSY2Mw0QSmFBbH23q/g+dtMV/eiLuB8x61nGOJq
8rQrKadaLu4dbCOxDJz6cJd5+EheAntgZ6meXiVJFEKmHovwlckPNfN8lx0NBuhp
TeVFbjUDjpdKubRmSpsM92Ol0VYe/6QlzT2ndNEuWnIxhcP1u6WQnOgLLt9u3m2w
rONj/V6SSxQzwcZTwmAEJJJmE2AX8TwLxlvU3cdmERCp0+nmcxMRur/yrb7y+8ay
kFe8eJcl8JfaHY0p0yOjf2WsoLYsn0QXECYPIIf9y9YRtfQeA+pzUpo/DGH1FUtZ
p8bkQXuTJUsa7oRafIOlzGJ/d2poT+kd2UrMlrCDZMRB0duMW+BRbgg4SpHMr79Y
MR7Y54bTBp2QHNqmmAF35cWpvtavtUvu47wLVL0RRtkff5koFjmY0V++xyf6fMTG
fbZvsWtHnPY+7uGaxq+uyOZcbKClAT+cEDfyPPCK01PYNygvIlhh5m1Tc+sP2yxg
tbnGjAosGADkliLhrlDW8wXGATs8PPlbsm+vSQP2r2E3HlILhk8OXlXZIGJEpjkp
MIX1Z9NWllNSenMOqbRFbjNJwPRvck1weyI8o/w7wILygK7McHq0eMRNDD/ryaG1
/pPOhgMdgNP7BMwbNXH9s+yfLRta5I3BP/luZCT33Rw9sBHIAUElPdwrutgQtAWh
hkrWr86WlLY9YKaIlgwl+ifw0pAa0+UP6c8NFmcHSxiAwVjQxmFa31TjvGL2HQ9T
86qg21WdkC7gVZLkh/v9E68tc8I0g8UcZV9Rd3MlqaiWoZ3A5Qk9NxmE9j2a3mRd
LIgBWeyTUnNwqTxfWhDEG2bZ6SIhOEQrdTsGz3azuuf1xU3kpoZZZRUKPlhnzlhb
IX7uELBsBxgetpnKjxY5i2fCIXWAyeiYT8IqG9bofs1lSsG1oYQB7X7XBQblWg+3
IkXnJXLyNPspyeAyM60yXczPEZu4L4JxOPlISh9RUzmX82XAh5O/bkYLfLV6PyQs
MwDyvZqhkHzyl2sehpz2mvPagklSVigNKTERayUX1xuao4PVxBUjYlxKShC9Yxz5
DGfZNHK1hctMCS2K00jbu4TbgtJVj6VQEufumUuCojD/LK7SxnfALZuvFBImF1Kz
JulLR0aSq5mKruVQIg1zVRkThl8q+JmjgQGHfPIFEs+cqKINIVhkVyqPPYzxABb+
qcKF9SV5uzs7eoaqjz1Mk4p4YgRbQ60rdR40TNnMCWttEgVbVp6+k0delHcJD4Ar
Ex276+Qn20TsVFzBRaBPuVfidofOCydodx7TGtUihegPw/m6raydpg/L0aIa/PyM
H5gjYRSNHAYYjFdMAGFBWGfwyJyw28nqmyZiNwEtdzJM7pcgOjpOMneQBeM0z76D
MI/4pLPJcCHB/OBTETwiVFKQafzK2Rjputj/x64BiTmdHdYYZ02s05hMeic1ddzi
kWL0+IQtrWALvuUCpOfR6s0/lH9eASlfzIxObkFkaZgcmokaVTUhfqaW30Hy1Enr
R2sUjdqyQOQvK3LLYu/nlxC4BkEzK5VfXDfS1KDus83ZWSY4BehH2XlSxeqwCSnz
8WUTVqYjNZBU7Au/83AKexoWIA8pHmEwPzACj8gN3IgUIroecCUfPrLxExDcCI2P
8MjLA5uUV9kq31veDOK6WZGQ0U+3RL3aafMFaXbaJCnCR7r60crXdNXZt7M03yNp
L9RZUaXq5HdbWxxRy5DxWX0MbBBVImnuocQ2HBnF6dsd2kJ0e6vP4kRXSGEgqNx6
iJIOvksTldk72AjlDKICILbQ6t5p0XVZnE58+dQf+o/nUqGQR6+iMGA8+ehL/ZrP
fHenRD8Pxzbrc9AZyXr0knZQ/q40OOj21BF7UvKvROwMzc7SlUl9rbfnFONgnSt/
WgAw7q6JkEfklJPLgiHuavtRKgZqFjMeHbbV+svXI4khmpETLfK4GNtEhGH9PWLt
tPB4bGrWvEuT7Vy0Rz1feubjIMOsVCTtCmb5L2E5yqD8erWpk4yFW/SyLnHspKLF
FPSYr4uZ0IlqGSlbeZGRi3SZv0Fe2f6IHZd5eAkMiKh/9wwY8rbIUQUFvgLN2vkY
Z2T5glnR4szZz1wR7vmRZgDxs5yBrNBg+pPf6MkfAkQxd7WDNFY3ACgqQCqCE3Fl
lom4MXpwMVZHguotpUM1ubu58v50o9Hq2nqrZBtszWZUW9oSRD/T1gTxj7jWIS02
10bW56Twg2lTMQ1xtCrZBIso1bZ+r6DKP2rQVPaXOX6iz2sm6OUb9ln9uLVFIfBN
wxdro12unklU3no7tKIurcA/4f5NgGwQhgrXKzcphLoJGkuR83S/N/fH2yW/eBNR
xE4dFtRH4qp1U+WQJejHUXTHp+7Rva113nfV9A1AMk6u7+KOxs86rEMTJbhGvjKQ
jXdtRRBuMjS4lx2ElsBRrmnhX1eRDkZY3fOWWWahCYGO1ex4FfvX5H3ZAZ9z+WZs
qXK5eAjdK02yuT7jNtxXdu9sGPn5kkgjMcI/My63EfwnDkcYWOYtTBjF66lJ6v0g
7TuTSKKZDJKu5X1bXfhlOiI/VCo2HZlq1iMDAL/92sRcoA3rnYMevI2J+STqH/k3
ul/Y4rwc4iZw8uQQ/hl+WoZOoQaiXtBMhLMHjpQUGlQDAJyTx2dzmg00xvnGkIID
4vgPVdoCT1Ia32Zd5lB6d28zPdB2Vua0VJSeck5Bak1Qb+L/r9RCgYraTIRyiCPq
4BDnNtz5G15KfbMQqsklixkS5H45qxSyWmGjTTJP5tPuvSp68PNtTrLhjHKwXr/S
DrxAbAef6TsL8se8R/cjlYQJ4z1sXryk/mzwDErCpCTtzEx7O18AGXJtyR/9LREB
p/B93266cRh3f/D9+4Hn27nonit4xwmOlDQsmEdig4X69d7NZ9ukXX6fh8hJ0TM5
AWY+7+jDs5c1C0sIlwPcgdbC2/JfozkYqJ3/sJJ8Mkpdde65DrXgixDutvYk76hY
91g0zXiv6N9dXn2+6RDEHWrR8YQ/gitMvfBau1hcVJdTEG2VNfxdd+7jjOJcQk3E
k7c+lVBJG8C/ndeu3+No9xxmr9e+ZmV7AxqdcU8Shf2raQHl8+KmLHmWzPXpRHTy
5xOj44l1jFDHBAz2DMPZc/N1SZu3c7BGYhvzgBtsEVgqe6OuXs3caSRqZVnRWhEf
Wdlh2BgnJXkvmfxQGc2xGGfAWDyKGx59SkkAES0MyDSNNpVHN/uJoDrr15SF3QNk
wlYbE7vPjpVSdGRNzxQWbx0y6n2IHi71MBjfNrKbn9esusctY8j35/waOYKHkVp9
+Rk5JUMB0gUfFADQbFxk7FdldFJwbfx3bU8xs5hVHvysLA3xke+QaIh4fKwNe7To
SgdCV3zx3LWhkGNU7Nzy4UQC9oqq0gSdLO68DT9mWdXGMtvTMB7Wk7qm067zkbVC
fidFtnZKy4WISg0fSg7WEoQRkJruE0uCrVsWKjWDKbAlA+KlDwX8YFotZ2FEzoBA
CXybkpXHCDhJndPF7F1RjjHzpFaGkuR4CMjwHuMRzzSm3b+Ee+SUgAlcJg+x0X6x
mAwHdptRSLytSOyAFqZlvfe9PQZavioBIXSVH/uvmTtkOm+q+4z9xVs89TIKIp7d
I6TzsYsshm/oCqWTxjvHWGES87Ydisqr7JafwYw3mS/LGhMGW+QS3uneefEu9UfK
js8vt1N7ogySxy/3DqFezTf/Az7FmOCjALqs+das5UHl6ndNpTvZvUe1deqXRje0
BWQylT9uyk2FoIFp+S8q0di60NMkDUpyNNBdRkE6+xEP9c23riNaCKhpQNIV/a17
RzHHUZ5FyvcOtcJJi67JPpTFQkkXCvKZtvGfHOtbKEAxISndLB9cqXlx8HWguBFl
flovYD3BKDVranBUYFYRSBdmGR6UQR4R5BG68Y2tIUCdwefYO7XGgRpKSKTJvLIP
dWzO9/0WfKCczgI3vDaQBXEEORJtoHbrZQ82uQf+tav+2jwvPx3X9DRk2xydn9L/
tHVYwdKFXybqZP2aY+veMnsY9LPYPMjjKbYkF+v4K2hCX40wXmonO+d3qAaFdo6s
FaIykiT64mVtnF7tQTzLw4VDOy6/394ifwsP/We+pstKqpEQ0Gh2W6Z5tfgwUaY3
JTHK57uy+BFsw8wLsBN+HBpBbZlHsg57S+74e6/2GUtlhaXZpP1uDZ/j6PQsVBvZ
DkA7Uo+N6tenpid7Fy9ZQCCehZ4p4ZiTdDfFuwGddiGGwQ6vYF6gb5yZ1SODKZ/u
gEmEnqCymmB2s4PTuracLS/KOCq8kfmAAOU3yc89W83+jIvzZw6nnMgKoj8bYhiB
RXoQyAQl1Geslv98T+bp32xTPYMVDOqDisvUfPAAZDSjj4SbZPuOj1IBPmWCyw+e
wXOH/+ie6QJdkRKE1xcMPzkg6q2ayU85dMvaxXiQfaoDt8LfNrpmJTPECBd5f6X4
30b03+xJzlRGEAl/FBTOG+O9tca75OOUeNLogUFuap7OZcx68c3Ln0w2fJCgIytb
xkMbIYcquIkHxg4QR5fZ5XNJRUOnb2xnNIbFkBCPw8u1yJYXH07xNQucpND60Lhn
5IRkmWpl/Pylb9ejPp+FEaMyGphA3H785dhriSXJUhYulw6MKK5NJXbgCMfJri8r
SKDjL4XPQbTTGmskZaUwjc7ATWjn1OoWEpveFeJU8Ftzjs3KK+mxJfbUOJXuTXcQ
p8eFbwRInNTPK0wtZIXMnCUlDoD+/Ab6VKkRdpFS0rD/JTXjkYGHW5ocUFyW/9gw
vRLN0J/WC7tbqQynRdM3fTuCyPIJ40jYSjbNPmS3IwG8vyHc8dzEQIBU9RnC4rmb
Q+TgvIPbBWYka1cg3rXkp9/INK9xvJSclGQ1w7mAcZ1NMxaR5tyUodoXlKVZZeq3
GHRsxbEruSNXRyYfNudxSr2qrkFmsqcO5S6Wu59RTQ8BndS/2/WGEIaL769luLy2
c6CLz4wHuGxwcwqjIToK1RmgJkmLJGxSx9Wgu6jc+Y765LlVQ6S0K2QY8wCVQQ+i
oqtLHok89SyEgLC/sFsUd72SisuGhcRuK3C9XTEOmHZ2e7wIMaisMkQ7a7GE5OR7
Xl2NPT0hHndYRkGrNMfNUukEbE+k8dFrO0O0HTRlwV1lpudG0ZsPZ4WtYDHYb8VY
70mPnjwr7WpbCc4ztDzH/W2GMJ72kC1fglFs4Yly1Tye85YR19/p6GtPZ77rv7O7
/1AuVXj+gQ3mbWouF9c9qIwsAp8qRgR4OX/rplPkNXqcjEwjtCs+FE1mLsT+ZxNv
/midLJPr3gwQwQt2gv5O3rgY5waTPtQWBBoorB+tzcH4HBdTcDm2OIae6+pq2vCh
VyjcArNDi/GQ6JwByOT94bO1TdKKfQfMhh/7yTllCj/rQMlSufAa0U+rT1QYOxFB
o98UHgAp8GPpbnHHyY8YbK0BevtFPM7iXZpEt6Pm7/sqG4QqmMynQRGFrFMN6bdd
lA7aMC0s8g5E0iJTBT26gkSNZI6IPb66T0lsrhXAzjfhmTqJ8yueAQF3grauaP1V
c/+bk2KhkMjweUD6HVqmmiMdgRT5AYK3Jj01WB4mPL3d9PxclMbohCJ0XGgIg4P2
RbFTrDAOCscF+a8l93fBBUtQHH1+DIZ0EpgSknrqf0Wo7wCxEtvEiNS8AYS93QVA
FHPxlNU62Y38enMmjd8QJ7VIPUfd6p8dkuH+dur0tlKFx2u/0DlIGQZvotTpPIjq
ZPELJ8f6ohRW4b3PATmcwvBxwmAsrCq9hu7Meka2Q9ko8d8Rv+jCHWeaRN3302hM
XV9TgFYzfzUMyb3T2ShYZySXa4gH/I89YSrt4fzDUdiG+uziy6cHEbduG/vn4Xss
BjsGTf8QMn0lTH9v/Nw5etC5wkjCjmz88QcbN2yJWg5Rwk3atUxPOgcA+TOTDZZ5
j8uUjAcdvrUpBfbDCTREd6PBQCzO4WTM+ryqv5KC9+XOAhrXDmtpetZerzfG0bhh
+sWjao1vQTBx5UhG89lvmb2W85HsvkwhbDzXaj807Z3N11x3G2i/r06mRH33wv7Q
NhbMNXrk1TNC0ustoMXFdKbeESaLjzeXn+zNsuK31OgZiCbX+nlUtfBIIqfaTONX
SC6OPFUDeQLPErhenZiT1InMA6a/GQIneSkqHlpFasFxRvExVnGw/3qMbfVZKMKN
Y4VngjT2+NFX9qd9jIhVK6/yyaLD7z39uyft2uWPsi8a1BW96/sGKYUZ6scypYrI
LpZWKdeWZ5jkSXR2sOpfzzG5YNnOr42rrq24JpL7R9xT3aGYbPemzJ/wRpTAkPo1
drAE95Kz130HF1K595pGS2cyZn9kQwrYNnMniMQ+Fv+Q7YkDzTcga1HaQZdQFIC3
pjOzjJyj5CCbPXcvFQ30QHU+6MCzqHAzLG6/0byk8M3509hQqB/ua4VDKpRd12AG
cPZXlHmBhY9sCnJbD4AdYzyY8IAPYuU2hPbaehyBVjR0u5TcaIFc8abHuzj8EjZF
3CmuoCduHcnmJvYs53+6JsXeaPKLBMvU2/5J9FSlzsv9laR8Cl5Eriks1JB48h6L
B3AD/0XKEK7yMR8lHXR2XqfQEhG1SJ0TEGOcQHwPIaIpIT9poDSbJtiTADCwoKYF
ojhjM7Co+OT3P1rFPGZWFjep/9JUbgsNulVnH+nOAxyFfbaHvPoQSiV7IiKHyrh6
B/XRIdugXjqzi+CQtRaJLaXlxI6wcMdbVsiYM31AFDHtmqzbITks9h3lULdE+vQ/
4b/kx1uX0Qh7h9GCVedYXjHyqNliaAlz8NGpneYXQbGrTOoyi7UMb08mwFoHTDtk
2GQpA7uxW8meWz1cd8AQLQP4Vf0bgyhSJPqjl19IPmef9Jclh17E+xefG69BaNcq
eGCC5eVOPcUzUl1PJu+qD9wwsAo4RGh5BLiB4jt/zoHPyH06bn4x2YOS80SbCjMJ
xlDUdCa9cwJuZnwMCRP+v6KXWNbIA4tX/Pq49hQUUTjUcXe0RNolHGdDRrlzL2hy
kJHMWOKMx60cukLp7a0Sc2UxvQr+E7jhUE1JG5ss4kjU39lNP4/7bmLK061c7EdH
Y8eAMxtz8A8sKXvFpYQ8wz6cxrFxwAvaueZ8zkC1yi8FEztLPS77tA5JFmg4U3F+
zYJshIH0x0odft43gap3YDOlcCe7IwvkbCH8FSh/917P2c1U9vGnSpZupZLCKmfQ
Ts3ogs8UWDN94LTmMtzIajrxhkDvml1+PaJhFqGXTcMokNf+KKcGg1M+DdxZVmJn
yqVL6nodrDdsIDkpOnC1LGzxsgsygWxkF52UVmilLpGSJMjLeAW5WSGTSO1gX8Od
43Pm9UI0+Ot3HmQZlagYTuV2wSNdj6Gq5nhjbjRl15qFGw+4xGQOHyMFfAtiAzZR
+jSPcaE48bsjWfwov74oIdrmOqTo9Uzc1I4FsjK4yDe2rFH6QSsnxIaIIWJgQW6L
bM+b1jzq0prvjY/D/HXLQT/lcSIrg/jRUGVTGT4UXmBxxPZthkmwXYzoKwvrHHBu
aexK0x7Hw6Y1RFBtbD8ZKHW6Rw8rqJEwlJwTQa6jqdEXuIgnaEZKpB9ZBPmdnROk
RZfSEQQXkBCLYAI+lqlK7YBCleCAF8/MDPpbsmbQE7MjfcU7DmksAQb1TccngRQ2
98BDzCxvIUS0WOIzzOTxsC+4pLEYgZKITUCrJwUEYEahQHrIwmst0Lw0vORDuN/z
uCpslDQ4UpDFHCNo5C8EuuOAfHCFrbZVhSJOx8e0pi/SC1IIiW8IU574Oroo0kBA
4ZJEZlq0rRXfQReSyr+nle1wofvdf2LuZwZyUhjq9S+5TiTq7BUcoBCr2XaJ8UuA
mltvw1E1Fj/M2P1CIalNgDuOgQxV+oA+p9tDyDdjibYRUr9m2C2njS3VO1pxMcbY
G9Vgd15+knbABRhrwhMoT8dj8f0YetAyT+iodwQKDv3PMSr069hCQ7wOAbkSx94v
OYTDacUPAwOpKFs5BDy480tiOhKkyK/LjTikfuALho6ZRU59Uw6raIO20IpeALW1
nn8Ri/7Dx8Et45ey6I5QOU+Bu80Kemzl1jFkEWYv98P2QmO7v/dh/PItU62GdbHY
Q8HGiGZh2Rv3vbIem4A5VKJUZXUTqarS/qbUc0LAWSDZzBd+jXSQ01Wruewhv5vb
oqvSN+juykxYc4TYKr4K1YTn9SyELrajIylBprhh+58b0bW2JtorW3l+qsPhQ52k
TvFQDK/heo5Nvfjus52ctNxYY0fpwlVWexSL5LD8XyCoXmsRJ5D3g1tGK7kCyMTI
Ek94K1z7hyQWZQRqH40pKzOt0adwW4C+Tr2Xk6W401lscVBfX/KxXf/r8IvV/rLD
8Iv+QruqU0/g9dh+ADrjcSDRGuFRxRHOfzdzihtCiNJWgx8j+vo3DOaa3Mtrxbt8
5X10tDw9rWkZN65S0wglGhqdWI2lJEcdpBHjn6rUspf1yxzZvmwl4zx8QFLFP5MK
b/ETViB8WeUh/jk9iPh+mWh+ORCz/EqVplwtaM9B7qu+l+wPmko6zVvyqfU34na4
3JZy1yUjtdJEyEyl7V2kwyqtL0OKinK+IVITWNep7MVcTcgWnz7g7Ws0WDcwtbmY
4ZTKfp9JwJ1NS9q57KuR1erZIRXDJwweVWBXjK/FMkUcoNQIHmAfWQKrtyvEWDJ6
4qPShSYe6b/THDCkV6j7bSvbF9OHrdCmFRW8b3A7u89L4zEou9ZcbusyIIAOh1oM
G+RO4vSVqxI8wDj3mg4akmoG2TAp8w0XYsBlluoMhUVva2aE2KYg46YNX82qMuRo
t9hBjPo7J+/TVvdIlZnv79lFs3ofE2+Pv0d0Bgw94HOwiWh+stJD5jU6m5tCHN1Z
+XjwKPsnSYcofd4Q3rwxWLy0qDysCIdKnm32t5Gdi8QSWu5WpSdkASNHPlXU1LRu
XkrFokBRByipWK6eyhta7o4fLiffVJpUyHdOfybdDhuY9FVHMYVAeFri8543cDLE
jJRcmOhfSM7z5KSgnZTZTWyhemAhjqY08KBI/5nbFz/s7qa7WZOcB05J4PkXMZrb
lMlmQvwoNQh0IWxkZi3jO62I9aSvEVCSqXObxiG91xURtKd6R4wYXvkWPdw7HgV3
nkrz3+xDT05S2U0QE58SgKEebbzpBUNm3yI+hJLQHxw/Lf83ABdC7vHOVYsHoNr7
HJygC0JZKhGVmJPhs18uYvEkHSzvpg8Hf+gMhsgjVPzIAXMtMKF99hU2zVL4Uwye
bveIATYjv4UnpsqosS4uwXaFlPotOQ1XKSQPR6tgaRmNw7hcB9DRew7XW5wVIRa3
VKGI66tUiJDe8Sn1zaMPnKGgGOY6RWO8YHu4uO/g7mstdYbWM+MsEbSbBRoE5rOa
1CCfyF9XWhBcTKxAWi2JhiZPfKi7klQ3fyvIIH5UEy2hQDSl9KK26T7tI9fU1hCw
Qo2NyYBGHR/mKahDRBMynyA2tin1DFvKCp6SyNZQlEM9KonxwCUJT6LqM+1SM8kx
/MGmeQE45pxeSFWfTEjIn+g9SVInEfmZ3GnZ/KaDjSuOUpv0Eyzrf6K09DbxVova
jwO6vuSg9UosuMlimlR2XSQscic2uFAhOJqz/y7nJ7ZG8RWnkh+frDIleckzJ1Sb
3ZveshQmxGUdl/gtkhG/bP9t86k1MYvH/mkW9K7ywFNi7TvVtnJ3MjCy/blPP5H4
fX0Vl7Is/jjDcv+af8topEPb8EKjQHWTkrKm6ICMzWQrqoHlPAlNWt9wzHdn4ert
T7CXDTt/bBec3O2LTTvzleA9u5q7wFBZj/wKV94fVOy+vQNKbBoICIBfgfOXFwde
Qi07ELQRdaCdOAZcS3+LR/dBQC3X7FQxdp32gIj5Olp4njkXmy4PPPdEM4Vv+Wp7
2n/cIsSs+Wp3BgpSCJW1HlCWRZhzqoa+fTYLFqJBo0wCy2WoZ5uV0cOGHUQiI730
gXVrNJanMj4Ifq1wFCQiaKj2LbJeB1TYeIu6USEiQG8aw32kUf820vBVKrJV5BBm
79rMA7auGrID+5HfLf1jPVgWhXcckc/FgAZteqM81snMBFSovVXG9if6yxk3uRN6
EK36w1GfzkdY6nEwBJ4e2gXcy13HmabOOU3EKF3TK6wCfTvrVZS2FPoy26+gioMs
caThdG2FH+7nr/v3e1GJZMd0XyZwBscwbs1UGkxMrinLJK94bWN/o+nQdWAsIPQZ
dF6x6dm+9m18y4GfUhTe+LpOfBw992Arq4qmfakI2/3EJzwt0KSeOav4ca/UfajI
ceb9/BVIoZ5ckip60xOfN4mYxQUtv0yius9cEtiehKGiVvljMp1HzTBXlHiM0kEN
gV/k/NUO6R/iEhf6d/LKeDaAVxbpHrgMwetH7CDoGsRrVZJuPJRW0/Om4WovkcSp
6uB9gK/oFy9Olwj8zYJF/9GCW6k8YOGb+hCL56c1n9OFm4o2xG22O4SOCXhShhyx
aHUHl3KYnHxFa08PHLT6yJMzjpUaiDcGlTp1TP626TCoFBZJBsE5ubiXZ7jUAhOU
s1GNZpifQXnni756Uy3MOYbHbRrrtkQlJ6XxLM3udrcCc6F7O9dOxsOYb4t1Y/IP
w9o5vLhgVNXed0iCt7EaANB1rAvx3HFLuxY3Y6DkKsTEOn0J+y2zKRa1zvmaDYYM
ANHQK5O4iOb+Zo0DrcJFzREki2XHzkDfezpKBMIrSG6N0gqOdIREOCSVVhkd/TlS
XuTFa0S/UgNQMgF7i0GQKIvFsKOOTJN51GcHPuYz87gNzMtvefn5aJ2QHhUzdx3k
4ShwRQjsOl/GKZ9gGnwqs4l5Uwzdflt/weZEAm91/0RZIK8Z9m27D/dO9gloqetk
zHuyXONqVOIKzF9Ro6IiEXRX/6eLWggy2q0Dux7jvD17xdLjYQcY0zD7+rW1L1sp
ptEAZXkazN9HsPSUwkegVx3S6khsqxiQcGHSv43EzXJ4S2zXa2oP0OqohE0aGAMb
bG4c8afpUp+hT86oGNnxB7eDBKpKqgLal/bklCNp81vueYH6EHtoUaO61sVpAGhb
JhAjlebLt0yIr5pmEjMaEl2dsf+ZnC9Z6uQPLOSIQ859acNp9BYbzYDTiGtkjRbV
JJj0xYYD3DWk+8gTdso1ILSKk+A8YGeue5vnx9COc6G6T6ccAEZrMIM6+++hXvaV
MqiNd9FUu2deHlgnqOdDz6sdOHfm9Y2r7f5YdSb4sXfw4Tp0pdKA5rYPHdfMqrM0
1hVcYEp/YpJTxlAJjJ8vyGifl8zzn5NaW6tqnxs9IFxBKeS4fu8bZMFVqeMFsTSt
lqVYdq6yIs6/XBDoGoPDfEtUGGV+ctwluPYfadGO/PRjUP2o8q/DIiXrzorSC2Uz
nlPmG9Xcj84rMzeDeBI1hrlmOOT1omk0rXx9MEczfTunzhkZ2CvCZHThe6HFgLTR
tvw3fgJYQS3yCTU+3wipahLN2QkrtXVayONoZGMostfuay6ZSkFPV/AVhJwnMEag
EA8cxyMM4/Ewvf0eGXc7WxeXr252LJhYx5TKCc+9f5q8CKZXKBXCoCcTVYxoFqJg
O2jS7oLYSFh4x6d2fljmNkufv3mDZap393baSPTPEjk+vSF4yDaRrhvq1kQQC5Ow
8bdS7O1BB49jxH8fhSYcctY67W9jN8z+9MIWDhcO31givHMnx9JYmojbnzMbZCVj
Md0iDXTDFmrPCT3SOtS2EQhRh8dPqkf8JmrxFuaVeE/thVfOI7Ak3L0LzVr0rNCG
WyYR6cAAJKTK8ShEGPYw45tMi7QgXTkqO9feVF26kyfI4iZK7yzJVHq+y8lkWUW0
Am6rLAKc99KPw1ZQJ7g/FryM35uyIGpPohYLYm55CbSRhLbyb+ZSdVDsIfZGXu7W
ApNnn017xRzu6QkqwzQWyqUjx6zvsym/Fj0srwSitYA8Tyz+3Tu7bw5E47f9QvNh
bBErJablcpVza2j+YTHqAHcqmi2UJUXnfEfJkXfd0K3Ct7lzsOxz2UMQ6dPnx7nk
E+8jbHA+shpxKZhAtUZqB4zIs3hq9fJqwbIAQ/z9UULW7Q5x4uG4rSByYEfhElNI
VmYXrdrtrCnGSn8RYZTzJrOSLUzA3FLqbb45ccKQkqWXlKH8DIw4gxjW9Dc/bZa6
iJwQjfDrOGddmyPQVRbezt5OpFtIIPp1FK8cWrOUmy6Z+Vd+eI7dV1lUdYeEziTp
6xsLsS4TFKNwQjDjO2wk7W1LkEC/s0CPYsueLbfJM0u/VYBQU8Nbte41PI0nmWG3
gsL8w2pdGFd2zL9bLUVfuLg44DJuvQQlYUP9myM7fcs5hZGolets8wNOP/10wtx3
UUUvcF/BA8nn0h6MfXR78fSwy4Omndio4wWpMZruBMxHX+s6Uyr949XkVGQjpDJE
lsq6an/s28C80jVnm3e9k5Bbp6N4CGgAIOK61f898wvlqdiStA3fgeqHfWq/5Z79
Y610od5oR0dsMgYC4tm3i9Jc2sP1R3ckba+vMvNjeDMfrf2UGuGKEJCx2wXD5SSQ
Hl9/XWcGqajvdDlqY29PR5QjcslPd/sg1aMRJrHcNr3HCtnQwkJUk5PpQXFIkNCe
NRm1z+zUPSIVKaDG/u8JJTgyH55uFcvIsptST3AnDHAoVbz9LYyHVS0gHQ8Pf6v2
mcNnj0nguS9zsdSugIUo5budDm6KM6ihPwAZBUwJesGtdNTK4RoifdvMPVzEEWfY
1G/UkuBa5ZtQMEW30xz5WDMUJdbdqoA4SFyYg4uQuLRCywzdgmAcJMhcvSwgdiCD
LSTwGb3gBEDrQOq+NqVTRpCBmDhKBFKUSbiif0g96ib+68Q5zPBbC3ExcHHy1fmB
JZDDOTP0jHeQ9cTDzYiGJhhaFnsXu5QkUFsPEolL0V8m/ABnRON6kntxXPE0KGZk
Yja3iDywqu6f4wWBYAUytsArd8f/FEQWlF81AkU9fXR+a9tTOdOcPjIvtnN7mzdA
zk51lvcZMhJalaFXG2rhRCoGNHCmKf9za06DjkCyKvTHrKRD7nrob/uGX6dYteSX
SdgvbWrM/dWGVSvcEOlm94ryLY81gXzApZhdk6CMG/srrD6YKRTlm1/65eLkV4Kc
IKFGy+/SWeOFmlgZBmU1Jpwnn0exq9nEjYjqdo1dzY5BBb59PtY8EFNVScru83QO
tbNZrBso616Svz4R9RK6KcH884CHbDJYolpLt83AJvn7uhPSjTT8+NFSCSatfQ66
fznolxfVZyJHfVnkxxzCd1QIXfrwz+sGr83Yz6uf15UMAl6avqMZ4Iwg/zFZvkq/
8wLeTmvWd0FBG/J401lEe61lAG9WGsuIwzWpyKzsw/tQqFA1HL/0I1JMGS1ABv97
oJB1DihBSW7QBT+PRRZXHp9+b2LUQbg+/lnKHnmr28ocS4kY0+6WPZqmjc14YRkI
JIa/An3IE5qNA/GglmFN2kdZPVA+kMr55qWEU70WgLB4IuYHKVOBWw7VB9AMLx+8
05sN6b+t2PdI/wGe5OsbB5IWvzuh5kK+7muTTGf3buXiatXkuVgTcrwuURtSH5ws
A8a6be8gLCFI86gyG8hpm8bfRGO+H9EsBxSSyyyqJD+ngFnCe78LH5+EakvhU7gt
NUCnll8tMNKUP6I3G38M2hUauFCdPrGm7GrmwJZTW+FL+9qNZnyJ6TMp/j4fPkPb
xWbs9yvRi70rRXPaQnzD2Qt8YV+Y9/JGONLkUQF0W/Xnl65AuOEpB7HLlSI/9PVN
DxXuLju8D0OwYUmLoxLeHtqDbRGBaxah/Zxrdy7DHqUAK8VFWUD4pOQsFzLV/eGr
sQ0NhkCuvcLVGbKjdsQUm03msymX86B3zrrwFWQ7NjIlj6UPd5SEyjO3zsDBbObd
VKJ8/O3G95JVfmJaEqpDTeujXgwNUbjw85otEYfdaYi3Roh3vxjl2ugMIvjPlEMK
bHhQPGgDd13RF6aFNODYKCjZI+3YDBjxmPQzZWRijhEffJmwtti+7VhFs+T/859S
+9GPVli6W0nl5KBv4SkV0qaAU4qUMDrfWwyib6+TY74/MkVlirjWAh6SKMcFVy88
pvQmBwnFF14vFFz1ZKLRyJLV6PcvX7ux24wcpUU3txFd7v3yGy9K07Msu8+wHmQv
2IZ+bHrbPziXiLZ22JVjvOPHgxFdPkkTLFyHy5ZwhFFMTG5G7AkPbY9G/2ruNmmm
rtrOrUJ/PirZul31YVB0pf09vjqz3Jb6UhxiRXINTP3s12z9xEZTs7dbaKD40TKx
3lUNMLu3Dgjvkz39hb36xhxy5gZ7ogBtLfCU+zS8cT9/XmlDsNGI+ldCOwpImZdI
a5XWi0bYK0BnTmnWyVxNjSORJ3cb17Fq7+lpXf2AFFZIIsMAbzPJpP5HZXRMbIN4
tlHwfsGiX/a0HcadXBjZH5R5RBdFZ62C6ml0ujQz5c5SbaQ6QmirWFMyIEOlahb4
a7e2JGQVNKYolDI6Fv3G72MMVUQbPOVs/1CMSENaMG2ggpEqNQfHtuk4bKNba+98
sLg7rJIbPvyLSCigbLYvZDLO7obFb+fwuiWvoGfQ0cswV8nPlo7vv+Dw6yZUdBkU
vgWZgOYtHDuX3xa2ITfs/tJqWvnpdW3zqraw+JQWi7OxvUyuVt6FAEaBJ0GJnWHk
zlUoVCqW3zxLsEdy8ux3Fb/EMmKkIwtZdZsbN65lTf0f4inP8Ryph2IGoix5I8hO
/cbMgPjL7fjP0VmKlVUQJ4tLEWGMDWn9g8Ib0Wuy8MucM5rFIG2Jqp3zcicwIvBP
j0G75SDkqQvanv/6/RsJ/CE+hyAp9rOaZ2LBBLltExHi4PYOcioqbI+In4xv3AGg
R1Vf5KgVcccK64GyPQFaEIn7t7En7GrmcJLcyKDaEeQ/hiXNuvWNUknFW9CQ+3f4
OGCnNpyiTk2AQ7u7dlBtnOTaOje8TV8fn3j26Dzl8y4aTnEua5+UED+pHxQraKdt
U9TxIRZGgG3AbH0Ef/hqMFGAkm/O8rFldjCtye97uCpK+fwvUnVsIKOlnHnZJsLf
J59FYYTLoMAws/D2QGnlYOUhL0Qj64y6tE/jAKlZwPw5g/swsc37LBYvWvf+nXQn
RW4o90KV5nwXJQU6JJMvOSRC+pJXzZyoylYkMMrgyRlOk9CP49cwVneWSX/CdyRL
tKXofyv1bCP2xMtZuKp5dcbXg/ka5lD1rV4BEk9uvbDYmudwV0kt5QLUPze6Iby8
eTd9npTln9MXh9vqzLDsNd/LjfNYCEtYyrE4im/YnETqbWA7y0xOEnf0Py32vx2r
823zrlyWKXA8uNBE1nHjf8CVCUhk4IJbZHP3gYwH4d5zibRYSlyygQej1WjcmujI
yvEN2SyV/V53Kfh3ftqxYDIJyV03XRVt2AImzH79+REef4egBOw30G24np8DJINS
x8vKrBtPvLxH6lBLKt4DobiShtp9mt4oGthU1NdeJZX24yAyTaZ3tMspqatBUmMR
PAZvsY68wZ1DB6AAkKRGef/0E/EZIiYXNGKx4PkGx7a3tvDjh3JwQYcrM0BmFfSx
iMlj6lnGx7fLCcdIkwCzgPPIhsclb8+8VNUgatvBFqBsY8Eur+5SB94ws4rCp0Kn
YhoTSuNdEFY+O26yP8EaGuBocNR9EV86AQE04qOtMGI2xYhrXda7IKuZwS22Jr8K
UITkVsK8QpNMx2wlRrI5DmTGHzFwi7Xuwc9JiJR4Pj/hhspv/cBEM5Fv0O1oj0Ap
abOCxlKg+coiH0abP8lLpiSipcGp5Q3vLfC5RSUoHDb33HqGH0GyfcL8s0ZF3sPe
TMO3pGNsumbeyO6TW+tMVTrS73SW+ET3Ge8hlcYNyAO1uPh7bjlJxZNkgns/szlk
SyuCEAzYaj7fiHzlQTD7bho65HVVv3Dwr4jHab1JVlT2hhRJC969vDqd0P63uHY7
VG19UsZk4PpPrFtsPFz3L9f+BfjxKI0HoQUzlZzlqBKyCHUddzwmcBiy6Cypc4EX
NTsTFE1dCOVuhkjqBWRRmVSDhXBlZh1cMtxLZQZK3QBsFGuoO/c1US6VQnGSVO4p
2KVPBL7N6uSM1JFf/9upJiZ1DAGSBhTdoNUx12uG0LFeYP01WYgsmXEcg8gwg6uZ
cvyy0E3cYzcz+tXkczxU+39sEqgKlwSXsf4GWiJ9+tmzz/9n0VjvqWpaXw5Ne78o
kyf/g1FY7ffhewOMRtBMVA1QMXobnGhfwJ8pXqa21y7gCirHsriDsioxvm1mQKxo
54Wj4eH2SqiQ+lDlmnLGYX9TRJlZzHLEau+XprkwxM3e6RbocW1h0CxuVQIPE+ih
7DRbk9fFX8/57NYtQIyTAllCRvbhnvi4VskAL00YCo5yV2P8sJHUDTfGeu6zNx4w
iYafns/0DUjPQZ9GEsb7LeYMKmjHSXBYj2rBXJ5X+K+Kee3GHO3J71Dv08blkYJU
+WN9kjNjSrwmnikO61fF1HrMDytecSICJc/lOsB96MTI6THOugtFC4GAg6vnvaVI
QDNLtU12Be2ZH7Ko0K2sk5qMKQa8p0WxxOBLFBSF9LFMsa39QLI0Mdj5p60GAP5s
KacHrkghfOV5X9snKExtutzGXlHhRTZW8Arrc8rcziofDsTBWl++amH3I+oXutH2
mEX3Zls4iFVY0s1fqncbzfV6BQ7aZ0qdK+ubo5717/pB9jIu/hkjUELRh9kflRYF
J4z8ngponNCh6oj60Poo3AtCoD6/dexj+jzRGCrD4TPOhRWuuGMHCJbIHXDQIApH
QMzJbv7OyYesYkEYYMHiHDpj+DFch7ui7In2qC0Fj4MIvRwFgADQzBTnmuehRgWH
NvyKONs979A4hTCU1A5+eNKYawmnsD1gP36WSSJ7z2zSLBlQmcLrzvUOKQC1dvor
3iNSqzMcI/mlLpk6ey18U+mqur4/ie0tFZg7rBdlInoN5sXgvIux5b01ire8o0BN
KJzWDpMIkANPlR7UueBGqELGrGkmnHt6pqw4d00gGnye0GfftPNqOCZ3jv078JLR
N4JL+87S4NXhxTdz7io9V4eXsYIctWWLlTziJsKf4dIkqv5QKE82QoAEPGQF3QUQ
4FnHT+UR3NKWmySI6gJFUP7EDhTYL+Kl9j4my0FqXwfw5IT5gCVl6hfeBtBnazXf
dsiROU/raJJZtNa/Updxf91QoV6sF8kw+I6swMkzM41DT8aNGy8i3IBWRT7tEAxy
8dm72YvGf47OvMLSARhU6Ma7CjWAB5L198WZ4CIZL8IpGAbu9W+lOy92DjqMQeHx
ijNOeuupxCkIJamxA+Az7pjlRJqmWcuFmxpqZtFvu23O2OyYSyvZLcJmiRQs+3Xh
YTDMpmrwaOjwtzGinjNnbGYqQY0AZ3MyQ8ox1gUnEexntFw01EMf7kMRK01Q20fp
qDQ/x5mDw9Pw7hKRq8c0g11jn46D51DJJ5FPjwgkjIWFkpCVajTPQ6QcX2MoDojn
5WapcMv9lPL0/+/jLm93Qu2W0aKm7U1L576JArlWsPjS2mP9KeCL3YViz7Egqz5g
W4IrDFh9xhP7u+JqUfBMF5nnucJk1WRZ8rc1FEtvUqZIBGtP6vTzz96xsLyFOaPq
/5h/QeZgCfQJbKJZ9mfRb3W1SI3Gvrzk9thmp/u61lOK4eGMyf417nwJvZj1fujQ
QD8Cov6NQFd0ZnECYtYP4jGR9Kd+U7f/8bybR+xEYmh84ZUi9srTd3T2qZknE1YS
ZMdJoKBVb7pi11IfNeDu5nzZewOV8sNqAdGUYGuveFOMziY+vjzoPAo/Iba1Oy29
b9mtJmK6czL8Bw/bENARZEKeF413CJVtkPrjmkfIB6XucxNSBAzc1Lj9S1dDAcNr
jJ9yBNISVcTOTt/8GLfntbNgA0OJveNZn376MHWR64KdXLGSgh6rCtSV5t3Tn88N
K+jsLNX1wm44GXQscJcvDuKxmjAohjav+/ELFJc6pUzB0XOeQ70Ge+MMSGk/Efxn
Jrs41u9nYmzT4C2uf/pegQyzf8zm+JsWTR0UhQys98uGeV3x3HnBracsOnlzz81V
65eiyQJAGMp1zrKff+x2gpwIpPTXJVE88YeJLS76/UBneJKOYbC9mTz1E2FQFyw5
MkojWgwB4eIE2x0M4/6MbQZx87aABRAib4AQMugrDdfJyQs23hhqD9H6DFojoCy8
DXOCnr6Y3+mULxte+81sd1qwTava4AgrS7DNvGcd1Nhbkztya9SCSPd9MrSJATDC
6Dqi3G12GxoXE6USUlD3quhwBq5+Uz4AS0cmywl0QZHUecBbbThwcaxZ+LJGba1q
QaT7vx8Hv3+IPVb1wzfL6sActQcmKkuDF82lcr9U3Irjp4npdsDwhj5bAjmhHGf9
hjs4LZRGvkMqGp6AAH2FgyAC9MEx2sWoOBGa05ObxfdPmHcsFwhUjYw3TVtJU+LZ
e/La8Bzs3Nh63UXB8OqlGpdPDfho+SG3ZOsdEbmYGZEqTTRqmvAmCHA/szEOqNdp
M0oZaVkbxUO8staJcZcSiCy6lAdVl/6WveA1OIEmOpfMXLiHgtG9ykQywSdR65az
qeb5aHRfZRii/O3cyZd0C1+N4/G8gmAdtVc5gvheXHhgPDBVraHjzURW/lr1dxrA
tClEJoSVSoX3TNTauGa1xvwSuCiYBHo0kBhNV9UvNOSgbSU83W4CfYYS6hU3jcCf
pObddcXEvN7royGW6+iRIABw9kDnA49XyO+rPpfUYg8YGSj6Ob0UH8bL9YUtSE7m
tRKBXe4/PZS0CXYgGqOQDvR/+LDs/0xUfMk65Dc1K/ddbIWRPOiOd1UwbbkmTPu1
d219aY1WA/oDAnqv6MNptuGeIGc2wVxHkc1u+ICiWq46NOqneCi/oEgFhQ4JZ9/t
HJW8VgEgarry5wJCzYwGUz3VfXYlTfZ3hBKcd1vwVV+AsW+7pS+V47IfFReWZmBs
kGR/aoSm/p4Q/t1hYkcyzmml2Vr1U7QENlaD2n1V4uKEfQ53UdzTptIzS1JpYYyA
eVVNgIVTOcFdvS9R1ZE9Qj4amIxnZGdkFSTphWctTaUxr20qf+nusKEwFV8jkXMg
roYVCy71Y7uNGNehNAFEfSnZa2egxOEz6HFf+4ctcFEPZBjP6BX9KLLQt0aw6RWy
tD0ZI4R/fE520QCaOR9BdMaz8JuhHXM4JnkAECLsWGgplHl6AgA/NzTUKNH0tHuf
xreuFvYzb+ZzmK+xjRnYTo2XLwGvsOK5/V76AVYXPw5glao3KYzvQsb0mnsSy57F
u6utdyp68BokySc3yP8qGl7oRzvX6MQCm/cjCcl2GndmaTyf8PCPu8TIWPPQcR4j
CNOjUL9GrIVqZN3pfKkKrSTKrD1hxkWWzj7a5sjnx5jUka9Mwpjxnlq3XvmbGGrQ
ejGGWhkJhrJCr/g7I23BgnNZ5gPg8+ykrUesicIaucRvlPjMtiGmZbvaLw94HZ9A
wnChtlz3y2pBFtBjqqf6QbkcKOafX5ekKOZZ8Jm8HuZkbZlEVaLZs3fW/SakYvt9
lcvFYOkw0VVHTDl9cKvQPouWEzZb6hPCaKolXl2hblvgIAzhLHbw8JcgDxmUjgv7
x3NbvgHjyEY1sAjXeZhQw0MyZ3g+PxmYbcmjYlpVMsUVaOD9rFzWYvGZBuH0VrVL
1fS7YTL3d3v3hNTwJ47EfEJx1UTaBly/ph0sVaAbgzQt4shSqJmRUtHpsDGF7sfM
siYSLVfxiU2q0A9NVJXGLNXqI4WLRoZ8JyN/pxCTlN89+dXvV/niWR6rzuedMLVu
Pl90F0MZ37a09jpgcjMiW1ibheK7FjOQGiBqDwgARHKMMLqKC7bQ7R7MAYQ3uSEM
2OnGWdw+yIwhsv/Fzaa9suhRsvNaEvRfMP852fp3PO+WsiTNwVGEpEW7kAcJ32B5
WpOTqJ8cwQLziHwDE98yOrudFHtKQodJwJEMmoYZib+Iqr4RSz/cpVSplnRR6RHT
IFkuRKhKhD0wat2HB+Jxq7/XvEPdzbLCRtKM586Or48vzHskVZSHrqCdAfI5rhqz
Wt3lUYWpRqyJABDyReaQ32EcpG6MPttbROxc46foZK83ygk55k2/ir8A16MR/vwW
VnadXUw3f54QgOZ0keAcW4FZ8PogO6LMqTh5dh2DaTCjamN/titZUlr3xl4lSyDU
NmEZNsqQzBUPN5ouCHmTM7NFR6rNMnpSXMmsWm2BW7p6Bw94pHWX9DPUg61Sgt5I
F8z6fvhL06n+i8V9pwR6cIPIc8YUihvNRtga1EgM+J+MSrTeu0sYiFBmERzwk0Sm
tRYBljq4qxh3N9XTaDk+SWJPud0DWBrGHhl/ELGFwIroNTu7kaV/mNICSsU/x/FT
Z7LI5nxxR67cVRBdJWi4n/yF4gih+ztyE4Zf8MCf9NrxN1T+iJaXrDN7/0MgJKhK
g7mhBHxQrZiomNZziClUTOrAwYTZ/g8SBKFbjIXCkYfmWPmx/9emwGs+ugb6dnau
D3tKvFnAFXRUykC4D61nhIP/OCiMv1+INYyQ1oZbZ7XdhNNNd9T3wjoc+LPu9LHI
QMKhEyn5jITZ2X7ey85IWMUyLlmpZHeyUc+4m/H+QNIolOfdIodilkQU0XdC0gdJ
ktzHX1KD0Hvt8c1WMeYIiIyQfhFD1UmpngrsjueZpbV9+hT0hQJzHBoY6STwhUY1
aUHCnk5cWqM6Uy3s9aNEg7ItQHVCiac3eckC9XXdMtTJDbLtANtp5ZKW6495rx7D
S8VX19RPhVYT0iltTfIn6Rn3nugzeU6tq3IX3ekE3fJrYLaGsayevefl12OrQ3nN
6qOXRSmxoBT95MylGXTDgHt8ZAJB5b01UGXOEQ8dAAtPIOrvZRizn2y//2epunzr
U0mvPK9MrOFhknLRo3Sf6y6hXZnDX7k5qlleZsXZFwVULHEmRmvSdsVAAKndONft
I+e5WJYVrRN+MGSngdnhY24Kl57FNrX/xhNDUR34ceVX6uBBOdQXSqQ2pEe3c58c
oFWFwnvTznrZqG0xwtZySBlxpiSwPpxTef90ngwifRZ72bkfLIYGnOD1K7XmBYyp
6qMof/37e5BeyF6B6U4eMBKpV5vK6TXgwcR8H+5Qa3qr6kMJApmBuBXvrA77zUP1
5NJHig5866b0cwJEitaRcYLLQk5BLuYDMELdOufqVJhASm2sFMcK4Fr1C2hBcWd4
JyJX3k0xFaPru4Bb7qU6QbB1Cl6gxx2iugqWIrY++2XR+0UhWhQ055QvHifjPUyU
6TKSGuAaQnM3vSdjNpPapfXyCsCNs4bketAw/nYGORvZloBWJ4l+Y48rL+ViZ0Wj
rRlcy+zlIpY6kJXB1di99xbY2/T6gxWsdPgd1Um6Y3Ud8EXOrQqUrsPLBbkCJDOL
UcZ7jOIq1vU+g3huYQh+30ZsUrccnwnVEn3T1lApboHLEI41A0oT6LHRTEcFNCwJ
RE+FrdS4xE8vqLVEJFegiMgspz3BEXQjifjD9QNRPHTeSgqnBnz3Fwel0My7FYNq
XBZS9fTOESDcMLEqtxyd7ovyNyWMJTIIviad7XoyfSMYluAdFDVgLH8Gq+Nn9KbC
f1KrL/rFWsZ733McN/vPyYvKEF7LdxXQ4nv/GI115OHWhKjRGtjtxpnhs5dc/boC
oO3KtqTCxXyW0o6vDttYtKpNvDxbt4C4swWOio3AvwiRtZUceumid4RcYFRpLlh7
YVaJWGBgBZ9qjD8JVEGIPIB73et+jVeROMG4Yw10ORaVYMxtu1taIuuJJyXfF0iA
0FPVJNJNSLVPmQvdKJUeJk88d6FXRF6j/U2JC9MP/2N0aFOit369UqUYcXsvNk8d
YuQlJaAd71y0zcyHw7AmNGVYCw6WU5O+UkA1cJNVny3hdY/mackDu1iDdWMkKw93
zxkuxH0zza3DGzvyuoIP9KU7wmNhQT7nUOcsSzOM/WSNNwfs2YPX8gq3UzUcqlJr
T1/hISKow/t3n0iePovmck+5Bopf4pNJyuJ7DPUdSkK8csU/pU37Y4EJro17xEXP
Vyc51a153j8dBWGiiQ18xB0O72Z86U26UYkctJw3R4BFeMFX3ygm6HXU4/f9OT/z
YWco37a5xt4Uolt9Mz5lcP3A1ueNcmMCrfEKyFChOHLUPaNty5jZEBAUMwDgXoBd
QNE97QXPrKvWO2aPRKnnU6b82T5EJuA1lXPd3s1vkQT0hdyFEfZl12rlGdmd/v4E
IdXOLZStQ+Nk2xxafDKQQIOqwcuyb4TZjtRsahR7xRekiQFt/1Ph2M2L3HP1eH49
Bm+lMUzviuA3HdnF6ljD7pcTqgSQcaMpCMzPhzmf3q3dqy+jo+D1QcPnShx+oChJ
J1y8mJsS1W2LEpvzmlC3UsYn+VQvGXsJM7Z3umFYmW7Srh5T5wQrtH733dfhIcQy
MrvWyUntUW90o0xdDGEWAmJRKQx19afMpr0pAoLDEuctjrFgFvvQDA3zvZbdMOw+
a4Ru5tLrHEN3l2tpWUp8m/VJhIFKY3dpxBD3CetGrmQAlHDfppx3mbg7YcyyCTJb
jpJ1vpNz/roDAsQ+c8ek/b3LgSvt62/wiRSIDJTLQO8sF5oOgYRMwxc8sBlp1nZs
CriGCS9y8zg4nTYAtcjTTFeGDTVQX5E51oxM4MM3Sons7PMXYWa1SUmvEDyUCPY4
wvb9wDUCUPVpXOhn/BK7V6nvC+7SDo23oGIryLLf67jpmvnlhpVLFfY7z8uqKHPV
3n6zTyXt/sfsOnhTFnKPxcK3vtKcqLosII7B/sWROGRWWzl1eb6ipQBNc3Vn17un
+ItdMYQuuAv2wkRvGMG84QcPhYbOMB2rlZrRQTlzKPE7o0XEcveBt+f168vwvjzP
ahvlTswdr/jOCIaKspcf8zB4lpCl4hY2zWkjUtBHIP0MOKJvdgu/ClEaBcWiklLf
nT6Je8u9M4yP1bnA9hS7PSjYFwiXZlExwal8pPIHfFpDpw1tLf89pFkbrznYir/L
je5RNzeozZf1wDUxMr7cWyxJiDN6ao/VOxmDwc6AmtR+Bq6KBZwl0nCm3O9M+ZQH
8BzR9OWpxsuXOZYTGC7iwFUTMUoB7NT3dJxLwAGNx+dVjsTHKjJp1vIfLjOTBDdu
yVHsNr8ARYIrldVwnVtV7RBS8hBHbfUWmXtQwzpIS1Bp5fSWNKS/QRGzeSyy2tN7
LMRJqFBkDwtO6X0QSkEQwRsfvZKnMk2s3df9zfIwKy0/ZU3ewU97pqHdPS/9yaec
1tGaTETOMDQehOrjoDh627AlAgvzVw/G3eA0+OGJqG4e1BMJF6d9ziqUg3XW5voV
Fo09c8QppahDvmu7h1BFFrKU4jToFDG6BpgSc9GNqXlHHFB9VF7YfXUSnjKRBTUd
Rc4cwl58aQ0O+bAklQl8YF+Wqvic6sUTCKZ7MUL2sOFCIE2V5Ng/vKfjxxaGnsBj
9dV8AKUbLBcCusrHtPFTz1zx6jWky8sf6mNRTSP/+amqVQMSZFUaluNGMQVFO9W9
YyZOYdUTsE5oSi2YZUHTJDQ8pm6Ot33u8nR3t/AHRLwrdEam6xm8ndC43YfZF4is
EAxsbAJ7NBqgKERQBUQU5ZWoB51+WgCJzpA3TfWVJhgzWn1fNxKsco8xWxk7bRab
NNgDIpPZ0ylsQ/+gXxKKlg04BJDS7vnyUh5p8eW9eFbolm+UJp29GV+2Ixba6Wds
Lki3w4DB4FcM6cyyRC42RIyV4Gdv15KTXgVM1ZxDHpcWxsxrlGCwb1+YoeO0xbfr
xaypuR9l6DOkz94Z9dbeU/cotscrL39Or/QpzSz8tV/wGbl6gRC9Kg3wslym2uK1
UysmoIPiyqNwt2CeX69TPmLN6kmHk5waijaYE9XQrIvn6MYbxxxLq2ETFlfB6ztJ
rH+Ts5aOOI2rN3VFD81n4KBuPndjglUjfB8Sbtsu7lnn6f+4RosppHdKtWhSqbvA
jWNzmx9Li4pdL5B1GqJytHhl7AlsskzVTtS+e2I0NBDADdGfD7RJNh5+N+8Q4osa
E0kTtkhYHDY6aHjgNb2mSz1oJDC1SZqGobZYF/BA7udcGEo0I0JbNl+8csdCA1Iv
b92/SaD69oOcu5jIM+UAaWQsY8oN/VoZYuoL6RxWvSArPS0exuivVPt2ncC5pzSq
GN0q2lQmwhN8Y3tuQA6zMMGd1HwslPWzqjQr1qrrU4Pkcc9X+LEoSc5PEBgOl2z2
lB0YWpT5aHIAsDgRw1MktF4mANtLZB6kAEebIinpHv/q62nuLs5BK7OMgEViAe+7
0Xm27sGjoZp6JRAFC6D5PHD08soMKmZRZkpzqdLZ/bBiIB3G+M1e8Ai8YX7C2F/a
HrSvmcbPuVMg3qSnoqCvJB/iOXG2kh+09LMs96CHk+Mf3rp/7kNcExqMwCmrXezr
c/095eiVGz7Ih+S02ukAXfWgIPQcp84KwS7J2DSmdOrq8iquj2FzD6VFwmxwgd+Y
Cs3/2u008Zwwiz/TWnwq9gxsonUyUdlsGNVYtkI/qpY2SbJPg19HmzlNSpvKDZyn
E8Kouxn7zOL4MpYayFBOoJbq//m1A+50e0AKR4gE1dFTx0NutBMhvXz2OD3rU8gv
IwRANGLiMML4gkqSpwMGyQvcb2QjjNqEak6BD0tqT0xc9lVRgVsmeRC0Oo3Xrpym
N7q3Bl/koQwRt+sVWvf27O2hyxUKj/a62HZox7rdQSBz7quRFiH6uJK1uy7Ki3D3
/toEJCFdM8FwMnB0jD/Z34XGOsHh1Sz29c3z/MA83/FtmbNEHg8BEzGNVG9G9s0g
6OWQzgwKm02CNbK5Bl6mGhP0WBHgDYQmlpf4RSkxLqGJPt4ZKAdsXqZvAgXvcjaq
BvOAfOo9YopWJNUcj3XxqRebnbw/m0BqJdtEY0D2ro6jUGd2pKvfKg3Ut60moVoE
vyXw+lqeHoVbLmAKB/pKZc23Vm5lpz42XmURsFaZdqxbyZOHsfMgOaN3kKomhW2e
frx6xgEv28/VmB/MNSRXiNNv5mLDhJ/MS26k3raGgpCH5eqVlextav2IjKGJrJqI
22AQsQpE2b9BcXJpA568VVOOuhKTRtRVSZQ0REo4yCNHjCTyjd+9KwkTVa2aIh62
5/k0YRWqTiJTRt1c5mPR2LetELsijotnaiWEQBd5G/p3dgvBnZNgm5NJZqe6Dcea
fuAYTwEUMMdD75WT1PZcVA0xxhj7BSIbonBczDmEj8yNSyzd4Npa/BT+uQriu3Q4
WHeMt+FAtpkGw1EVwWAD6GxQMrqWk+SUDJ4ry/UVDdo8gg+zi4I9f83hJEaFb2GF
HI2qbxxaBWWw6MJgmaDyDE669aLw4cPtXWcIp7hJJdNReBSKPtwEfS6YfSwh+ZZG
+QOiWBwzog9m/fJ/lpU2++z0eevjZms0Nqnqifj3lG9F1cP+2pKZFjmgS5FcAS6S
oMKPzA6nNeFoLtH8pULscOq/Py6IgKp+0ZPBtmCF/U6Kdw/QPtgqT1uozvtzLxQC
aajjZ/n65YOHqPg2FxtlWyW33qe9PQj+P11sqqqnfuPEK3xJc/V8nwu6JJLA/DKl
K/8n3i1FfDr6QCSXr2Gj7YCaw0K5ObQJVWKbH415Cv6S4sEvXysM4QoxvDfyRWKE
54Szsl4SCcsWZCySfAinp4R7ddK6VpV++ScZ49i7x3ufPZiNBHnoBfBzIrgsK40+
IEBptz//5hnrxrUxO6c1U34AouQOT2lAN0cpHS7tCpE6VisNiGhRysDPx53uD0VV
LVcTQUWjHDaKyyPxzunhEmT4ZcOohJfKhiWkQdneY9jZpwtERgnByBBTMS2gtCoD
57wEkyrNy1y6/Efdkrmbyp9HFblRr8eeXI3Uqkslen1WhHw2HHAARqvOQ7WLMlk8
L5F+r0Zr1Zg1MQ5TPwYjgDPYB7W/RmGk4QNSwm3swmHwV85wT+yuONDGx5Yffl6b
7sYZFbnAg8U+B+DuYZsvNbhqeEi95Dm1uMMMRj0EKGNu/qnrQ7pxXXQWr1NkMjnx
XQs3l1aVhQzI+Z8cCQFIOcGzPlYg6Gm6nqK8l6pLMMdvAibMEuiFobr+HkfYVkto
xAZE5GkTpWtJyRXmylQuXWjJCVNsks+x2vPswZrm80jXRuzgnwKtWQMnXZtRzSIr
U+OoDoxQyUkwty+B5y49cL+uYik+qVewS9KmYEkZrhvaJPwIAaSU1o+7VHTSX64r
kaU1oniMHtGsiX6HdXIHU1tHMFsyYqf05Acs0zLFKtsPq4I0VEy30mEcACzTdXEd
rj1OJuGTTTEgY1F/+PS/U/zP5yWm+8+bT9Ihy2ZWqj46kLyZxYTObqnWriN4VUc9
swNTyTRBVjEa4NwOiuNUmcSqt2Sb16qI+W//u78PrfZNknd6EQuseQPYmyzE9f/1
kE2z8bFA2DfpKUnjjhz85bSwpAJaaj3VmeJbNyr3mG0t2RFlnhdYr8vqDB/kz2CF
taC3drG554pjuSiIw+RARqHcIey09PFCBNvsbvl8wm6Y3DUToGjlcFF4MsR/KkVv
NOmb/JKW+ajY9/jVPPnAMjH6hlXRKGWmKDGhFyp4LqalC7Hwl3ZLD2cI1S64EctO
ZWJLrNOdtDsg36EgMV4x6kJnJ43kgwFeUJ6a/REDhl6SefzuncTU8VqW41eGz9zq
7Dfa+1JrrR7Ec17leK5+gJHWN1eFRoRiDhyTjGNqV+hMEJqszp5AWKEOGt0QOnb5
wovJZBJNTim+hQ2Rk5/GisDi6ALy7CmmxAjMAO/O7tEUZ92fynATh3lRP2AU9olN
I6vi7ITag1+bfAZgI8s5NKywcK+GgXzn938UcXYozNJNG9kb2Jhu53ffPaqRVWXu
98jY4cUbGNjN9DCvXKWvzO6sLmaKZcQVPnsTtoas1bn0FlbDhhjSk3eRTiLE2oUe
9ZGKPuaw6b4Ljdi3wjpoapH6Allmi2P3JKEhL7u6ywyjVJ8xO6d+AQinhwAP9/g2
9gG1E9XWJeTL8ndxN8Lor2r6xmwSsfk2PH6cPmUl1+L4SAyPpQh+FIKk08sWroJg
aErJqmobf6y6oQdWs8dNogqBO3VW9qii8V/b4SZOtPdjJjwJHjrslh6LgmPginF1
qfu6+85fZuEwb0DYRapWDvelWo60uhTjr2fKhDnntuQm9beJmD4ql9hQDr/H/mr7
XI49Z8GPPYlqxUYP0swGYH+0xSUorsxEwvb5uixkdNCMEQiF78WMSC/dsCn/KSSg
KgJ6y9LZVvzyWKX8Dd9Xb5F9wmhnKzPjdDbTwT4Vc/l/nyKmVnTulP5f1qtbHUnm
DU+PURkp2wAzedYbVGBEyYRpQSUQwHuPMlXAVAQ9powNiCSi8a7GtKAITcpRjXDG
wLG0XSJrZ98NkaE3utilE1WOoiqPcGMRhs++PMwGp5Sn77XlhePyB89qfc9snRiJ
8y7sShDSbUzM/uF5WX/ZqxhQDStqcyLhsVQ0GWWGSk2IaXkso+mY9naKB1cuPAwR
Q8VZGi0+M487QlxVygREw9t+2PvSLCS0R7ixNEEuJCZvEre+kOZbrEn5xjTiSngG
QMkaELU1GRD/FB9JjHZCXx92LgX+hsy2WSnPowT4wmNqkOQu+wGgBZNJOWFYr3a1
IEhKoDEvHbjJmq5pporeA0eVeGPGQxtO43TT478TGk6V4uu3pYDMvhfi7i6DWjn5
pePP7wY3/J5EG0ugPim2XEvwPI7TAyqtvkwHa8A18sRmopa56KhrKeHLZoG3QuZJ
m1khSkXKsvkEpIta0BML3OyBEMqc2Xy9yKV0bPkGegWhiHr9ABV/+peltlmfQJuj
ZVMs8y0rsdgMCiQi4d7dmV07/v0pz1KxoOaeYHeXGyxuoiCZeNi8bL/3aphJTG0A
piJXqA69VlBhr5yvgo8W6Fgdqi1LL7uDIDQy8zZTiEf6OkZRZJs1qODc9G3+4PNS
Vq9IEB42jv3P9v09Kcyr1b7mrwyHg/Aq3uZ6AQ0ezplc04hWCdLawjIGTQBZgPWR
XbJQybMsyMN79dntPuDxSpJ+WzL/1EYdaRUKYZ8EbMEm3X6iNh05QvIpKJ+1jIbF
QY9k3cS+n0oYRvVXXhHyfWe/vf+L7hmNXUbd66LG3cTV6+P/Ji/pRF81kyYRMKfd
oiPwrRXMMS+3B5AQ+g/sz/D6XOaotF5MtGggZNsiOK7wzxuHz0i4m/kpTbvQUtZt
p5e33Cru5Lo50lsMGleDaGt5DX+0J5aqNeMWu282eQXWppibTaulJcENztNFmXml
9smJwbxHsyUBxGmGim026Momxlnx5GAPw0PljS7Yk82VQi8CBU7zLSBrO9TBGaCA
eT98j/21iIr4JuYB5y0vcatu0EWynKZWLhbcHWlgJ5vbq6Olj1FTOZA6Sk2i4DXx
1JNLffSfwNbQGcDVbhfoMfJzw3ZHMihZO7xpKVSl8ejaOWvkTriup93J3YHZDbzm
Lsip9Zzd5bSlQ1O+RiYlreCsTlrvm8riMTJqBP+CW3NDimwiYcoEGfLyhuHx4zQY
14Qv8pdiMIDjvLpxsD3dDIPX0HS7qXK9Aor9nQKmRGIsImQDUBDm3oWVNk0GbPx9
/8XdNYG/+6/bwZARQpGJ6gdwag+LfxLiCvib3J+Njp+05qClZpqmGKmfcmvLBiHG
0GLspDT8QnAIpkJVQ1Cx3nYTqgtegSsPk3ZxohTfpo0o4aYHZ+/GUcTpa++6faN5
bsOP/yml8py+wDPit8J66DmbvpeNsBWshSfDw7U9Uin2gIQv+VVesrJ4mLgIdMOS
2Lpn2g0zAau6P6nca7VZp+WyGlh+HC5+/bAK79s6bW21cj52o7vdE88DJ1ooQj3X
MGTBWE2sBQxka6zcjLDgqIrO9Vi0hMnCToh3ZwqI8ib3au8UletCRd48kmlihbHC
+Ser7ReKJJyAQQlV0oJxv5ydil+ONh63FJ1lEoc2KIyP8CC3GOpKXu8AkukuLu2t
/6zplGIFF+XtxOAMdaQ/3QUfJLgaNoYIEn8c3gZVrDQ5wRT9kvrCAj4KSsWfBj96
1gNpchMrVOnKsRvCVurY4ydLIYbGmripEgESh/ffAJQbfpKa6Z7BbOCU5+tFqYn6
0bYUK2Uptzy1KLEAFzFJlTxGoolCXShPvQizjDahK8FDbduhHpRJdTC/ObUIhpzS
2B/G4YN4MWSKYjAerGiKcJs61I+NPi/vxt1lEeaeX96jh3ruwgPY/z9SutmNevDQ
uc8pvosNW69HQt1/hqzz3HMJsLO1ixN+Zhd/pgvH99x4kJls9JsjUHZ1RLwN0rV8
yRlY1BMNvqfUbT1WO9cnxTenqAqsXL7V4CYn6+Lu7/mSFMRjQLn1h30yEVDIwgoS
rtXtbN1vPf0HDErarlQGO/P8HtPqPB1aIRzDGL20FYUFk3IyovUVuC3qCBGRZwDG
wRuYm1YnGZ3N8G0eEx+oPehwMF2MuVYzNVtPSb32UOjvh4MDo+ZBwbLh6bfwGKMj
HLqfCtC7TkOf96AfV2y4pkk0ZJ3PGBBA3wYp96Ta7Q4Ynll0YUhWerj0NgCLlecF
xzV7xcOckOFjyjU1ouxuMlOogZI06l8FhUYSzgo4+vC44QOO9a2PxlFNvUHOjDcm
5pTcMSUfsoJoLD4HRufSUIR1GR9fp6TRdV1P9J+UbuInHTn5TbCOsyluMj8KcQsk
/WAugZitfvLQBRXxGvMjDl2D7bXu6D7ukik1TFEAYSpOzEJFrmA9eJeLxqdnzcDb
iO+ZirhZNDZn0JtnWf/qks1IHAkn1Bjk2pC+4B+HgLX5oPWlRhnzDP/BzhTrlXFv
uvrXwsSu2SCT5BtxgbvzZ5rH9fVUhGLM+rQJ2sMYPelZhaxqXBaNtYnmqyDvoA6d
X10VWwXXvOLzxvK6qw/kB5t95flhaPw+hUk4dJtqQkoO4XZ1wZIrEXntRSjEmiWu
SakBjEG8SKqZQZ2avtHVNe45ANjTvnNuBTEjFlqNqYavPZdk7HCS8vR/qLPR5RhN
KMq2Svw7AB1HgWUXQ3Ok1SYZF/JBd07/6LIoAQS99lzf5VAqzvk6D/HN3UDL71g0
FMjg+eR0vv/5DO7/9ATe2artkamTylmOsDbAvzFPMWnZbMnLn06vUNNKWPXvedve
V9xHqgZk2sw6OUu6hpeMbPJzQYipN0rR7XDTRXv/aNGEpHdt7pezEujbQDGUHOY3
dPkgOERCOvwmoAjPr6ZQYcq8nJeU76JllaWf5ayh9MuSIK/mk+8ZmG7ghxrkgzPp
tkKtsRKLWU4jFkKWRvwFI/qmGaDnLHRmRoC8YJHc2qDwyRPuNGVx2kEnMaXUwAkT
eMgp1Tacv6M/Dl+MBvYn7ts8iHS+Zu6r1IAaizEeh4ZNrxm+RSO1oogvDUy7gY9K
wi5gsG30+vL+ke4Rt4kPduAJxIFJARJLqhORkzszmtzrwd0hD5BTCoKE3gw+WgCp
UgphB6YwHDwcIclkRzT3xz/Y6OQnbKVT3JruyOi2wHnM8lvWg9clAdSdK0WhdHEc
RZxlioGRf/RRTVTIsZpsfudhoIcKsfnhMKvRsIFoYjfRSG9wTx8r9G+q5BBWOnWf
I8Z0C5gCyOgAiN432s1zzWUjDV8uvVYKVWALT/YefWpmI2ndL6Q/QSJ/lgpppmao
yxSNAQUUao5zV7GuwI/324W/Mc7CPkJX4q1Fr6TEwXssNusIX+bWvXOK+uhXt9oB
sBPSzrgd5Wo2zZMaagKOEP1ZCHoQCIfzK0MVGMxJkHUTDlptjxaOZ59mUH7PTcxQ
xCmX6edv36IcrnbCa2EVMuSsYxOCO0iOnIgeylsKU8KxDWfSoGexDrVSvj+yjQMp
D1bjqMsYRWQehNoSMbUfjTlwVixGp8tRkUFBVgfL6bZqoiqd6nZAHLm/F9abnjff
DBUkeZKjpLoTKuoScmpMqNapBBfppsJbuGO4Nfkz5AkmsuPn78z2hZ6DyJjjG/XB
yak4U4Qya9HsJTLFI1a5W8FGpydoR/lPeumErPDp6mv+MQZEgfrthkaWG4KEEWhx
JMNqD1xVlrYq20Hor0piy9Nsd+MXVtTijNC3Cdi7cNs5CsTfGHhDaGkyS/lro20m
KObSBIx/eFw+HzEy14mPwoiQEX3tbuVwEI/h0KXP8cfnix7iGRcVEwXQFIcDsEa2
GrLea+9pMywBk+cN/YvPrHESFv143P+qP0dX5yDDnT5LQacao7eOGZ0JHPKlc+cE
shpEAUSP3OwG8UxiwDVCSXuith5Lb8UPe92RTyYHpw4P3miMw5z5UgUsErGF4AkS
lqxvUtU1P1NnYjCJXYL3ZrC1XGZ6PysN2ix6NzqysW75jmCGY0z+NJPrwWhidjkN
xIMiWgaF6d16IcHHGAexzJjoxAZInqduaNLxpcqotPBryac/aRwdp1ByppBX21wn
kRiHhBvoYS75nf8tSytgewRr9zT0Ma4Ms44Hm7fJhZ2IwlC12g1cO/GfT6PIXUNl
tFBAqR6DJjzcdeudtbuZgwIgoearnkp9UlaYOnRgPraxd3OZQ3dcNP18ClvXR2ju
jvAhNB9YIsyNMHNwrID8YDliQw+VwN2bSdNzihWNqbm9XZbMrEGAeXZ196uBLL4C
5TsemHM1dydxiXhF2KxE2G1sVZNYWFKSo5UmKF3mvdJ5qFpgDg08xfA7unYASegf
GWgKnkMC68sjMG3PtmccoR/94ljVZQe7udr9ZNUCrs+8x0GC7FjlQzl2qziAqeKw
quYutli8E3f0/y+tdrtvvJCa8dEVpk/FsYIgqa0MY1wP4PmNe4QOCwHDIsyXxT5k
4o/KSNSNZt4GowpNBGK8/Z0y3kdTjRSoOK3MeGdA7Y4/QeXnGbHrV5iCalpLn5D5
TV5Kq3VL3HbkVggvVwLwfPrG4DLLqym3sjUUW2Wn9Ka0CGzSJJX2Q3gJjwEt0m18
nsRtwctDel6bYuMj2gwzZp1cibRfl4z2OkYSezvazvdtiVReHO40v0Qy8VZfuB8j
rhluQT6Z5iK0yKdDytYPUv1Z2i7hY1jBkGBsYQbTaHY1rmMRhDqQFlIPTVW0WxhI
jZ0seF8Apejrf3PDTV3JOoS8D6PgNQZkM01306W60ATHoRedsH8Y3u7Arb3XfxhI
tVLnPO3lT0b473tuFHCZahkp0aGG3wAV7o/4VoZfY/zlNkwDYhpxdRJy3VwDuAMm
vDR4axF0tq0UH89Jg9ddwzPTTLU6ehUEtZAZVNiD83MpG7isx9eIQTXyFz8pI8Dl
WzY+m36xsg2sT0FAk/Zno2/F7ZLK0JcEJRRWWE1WCZWHVBvQgDSrIcojadQfECgu
0ShUODeOChPU4gqQeriO8HI0K6xFgeoUPXkb0WIqrbkTF4fdtWzySbnwmgqpu5gy
52z+c4Sfk/y2l5esoQ8YYf296O+3jOeCM9EItrH54WYeWmzlyO4qaYqwP3zKlWtZ
TaK2zAQgNthVyVDzvQC9SRI4ckZNcivHFg5rg+GQY/qza4XUptLgFxPjQ3s7wdae
7yMHuE9iumfVpy4Vrcrs8A6TCimIueLg20amiCYEU/iUD/WUqTfaoVY0i0LhQ3tT
1gpmpbC90AR7DTYbuXYf+t5sj94gq5r8MZ6WgEyKRrgaA6XYQwEfm/6ICs0A4eux
cQVv2mK+ITrm7LB1VudDW2Oe/+/wkEo5Uo1DEHdr1w0cww3clyyNVbS53ny0oppt
unePE4FBpVws153Ud08CilbxPIr5+a0c1TKsLuSUEZjQIU1sZBjF+chVi0cm4Y5L
vqmbn7pedZjkPfwnt2VWqwxNWqYM+/tRVcEhuN+rH0vM4gFF0zCcKUMqjiVGPdW7
iazOO7pr6k969h7ZHUZx756C3HRIXScMiI/x2ldCHoM1y2igFMcqFWBk5GbOadFH
pu5b0NhUgCg7AY47jSy0uFiMGIcrsm/Y7CTxHEyh2HnAOk6jvahPFhxSXhQdFApB
Y1CMyO8AuS+inySVbq+gylZR6e+WZ5ju7cxyHrpG0yXFmuJ107oVSFNkx0UnHiVV
AIBcixjfRJQWAgOE7PBX9N+SaP/2Laa5YvEkoVxjRCHNxdRxcUcHYrIJ+X2AX0sS
5TmzJ7Z/y+0usqXIBdRBxA+nVWRYmkB+x52iVUBlWity7dcc0ZQhBpCs4R6Dtkw8
xWVPtUGhj/aEPhraC7tRDB3bFBqoPRcTCHZdNJ+22hQZD1WjSzmTSdfq4B+eOJ3o
8mVZaS1kKW0P6uU4Aj3OgLy6/ZlDPgvTi7ER2J4Vav+EjfBRQCPD/JclYJKR6Yhz
DizudXuUndxAvdfcxj1A9/1YqrHgquAPaYxNfL8QtbUvBLjjdkiUIUVZTRvIdksZ
loa2u90bfZFsOx4MCIuKMciA9QsPc15B8WOTxw1dS7H48OGth1O2HQiEl2Siwk4D
bfBi07cByJ26XgAStXoe9+JyoOSoHutdQiipVsZ0aNxId8ojXvLQt2NH8VbWS6De
Wq4PTPDW+oopIZ56Bj7ufsQ/8b5i+VD1CTZNFEGd+VRar+U9+8R+8DhfG8BFv/h0
qoeBzA+3o1Xvna7ZXUdCCoySOAI5n8skZ4fgy4McOAgngHyZJLjnx2CMhHmKr93I
WXAfTAb0le/9Vnslwxwo89zQrg1A4o7vOfDkzd8oiik/BcW3Dp3xTyH7ztuqYpuK
9Xjk73qVnLonLoR2PKlJyMtHJ/msMlMAXwwIh3wOh7cTGM6ud6wfmFcIvm3a3W/q
jbEfionim5Y0QdpEnZDD+ypWUeAmwGdD8bz6bqAwzLo/R0vpaTJB9skqJ+qh9znT
a3LRFi18f1Lf9sXkahvJNAexn+ow/Lowy0wlurWfvRNN/MrMqGuInmCKZwYD4jMz
No1dk8m810iYXITrAUbx+fkYfa9aL33+i/LUFCrpK0GhgYoIiF3HDaaVyKQo8hT0
dtOcEEY6QVucoX1UbbMFYdSJhYadSwejCCd2WhAHmh3hw1F6mvPoPevZWgQB0q44
6A+KsfA/FbvEe+I3Mo/JFGICty2jZWgwnZQciMpwKoxmSjLk3Jo0J3L1qZsrqJ8Q
Z7z1UKEiChgy4ZKICBKH7+XQz2BPVNBhyGiyrUycUbCWH8y/xSV+mQ3B406Qzb6C
1HqzLdn9YT+FV63RkuBcr8XlqyNhjYiEXQSQbkZv0JldrCYvGPvj+6p9R18DKccb
fKo+UPc5I/Xh2+WzHgUCSDvV5TqQNevA4JOQTWkAtxY8PpQRh3x4C676swnR1aJW
tdbe+hMvlZFwBaAJ85yr/jaciyi9CIyE/fykpgw/EOdCKta3giPc61HvOnjjw/HE
r/wB2rzXI0YSBq+xE71xPgz3c3NU0JRgTh3dcPSbytw9anP1aN1pbXS3GI3E6PXZ
5Ek1AXyRiZyVbm0BQ+eZYz3b4g/XDVupiSly7bbyW94UL3wVpAl81g/VLr6sdoBO
ZHWgRBoWxQ3lsVJDGJrm1cVtXEDkWOsZlJktdZsjOFmtldnskHvWVlBgFnZckZq/
UyMlw99jJF3mbnq1uLXUoSUIYmCTuKrm9SNUjlzMfrOkFWQNQmAr6Ph8YMxdg6cv
GbbaNaq2kUQcCv1IYTVuB9kCor6FBQUI47UOHUwng8ITmjrITE19TfSazVT1WeDV
UU4ID2Nk7HKn2bfVzqWuXuxNaLgw29IInzjf5ysa9KLBcW2QFNgKJ7M0PI+aaijX
p4RIEWr6d5P7ZzNW2P/ncbzRUPpTGUS+oHkzf24oSd+0Bx9BWHuyuuINjB96+vec
FeTQbWtSHJyCGtisNT/pRcH10+X7iqTXeZhkUdR0IgoWzyb6TFxb6iZR6tlxbzB+
mzk41nUEEcQYxqSlrkK+fvGfgduEfponJSvsl9qZkarFDOpxpZoRlDWz0gTz6ftK
RngEMtbT74l+RhdL4or6GlsjAyjj5g4sicQ19Qs9XalGdNZ47RFcXKHAmbrZZgI7
LeFneB/9Fx4aFoaeDknhDjfMdLEq1ZrS12HgX0t73I84J2MX3jWOjwWNzCUfWL1+
Fx2fHwUhtaUDUkov6XgKw9bI7n3rpApEBPpmBU97DD+m1t1Ci9JdmpR2Y16RoqQj
HumtMvlEWMHhMaqN7ppXBh+yda66VhcfdSosrIH26ua/xcQyUSDrwTZGBQx2RopY
V9FaS2DneVQLMAMSAGovOncWRklDnLbJ80sdIn7OGlrNs9iN1p3hhF+F+CENNrWW
jkfxTavzGxEsrNVzw8niRgh0IaD5i+iF3jmZac4qrYO41UaqA8mROgjMIdpTBI5X
70OmZ8KEMVckLNbaEfKuQBEvO2px6Nie5H66J8lelxAlnWAKZOyFHOw570APWpwf
JJESIAOtnhRhPJpFO4qkbdCoD+xUaIBJByjGPVp3ZJO4urSHlpLzlsSnn8Yu0R9P
WdNUHQzmnn5FbyN44ZXwotZEr29QaBVhUuw2pRAUYVuPep/lOKITTdB/1gAAIP10
n2phz6iK/GMkrR4/nDrfGmFhHa5H/gXg+XDq6ECgz6FAZ/+30/tPHGAuW+Ia1B38
cbu4M7GHtRG9Dsd2lzuzhstRzXDHcSBjP9bRE/JtjtLvkmybZgzMxeyGcyB4SN3e
b0CvmPMnCgfv0sw6Mo5C6Z9167XeVLEYVHcKXlVg7hlxnJUGm52lnBDEKqaVjDyj
zNKRT6dfbE6UBp/wCyDLl8i9CnrVbabZHqH2JbWrZ913ydD7PzAif4OUgPXiRB9Z
y875SeHUSONEAKVJ2O31pxZurr4gxDENuZwrrHpLAcAHAXrKtFgNHWy8d4wT5yWw
LG59rA/MvzN3Qhmw4eDJePNG3Z/V8/MVMn1LqipkysAVk8vHh0uVv8OvDBcVlMEA
mFM6eJaXoYYMBCSDsq7fdBJ5WXJtYeURLxFKMt9PwxMRqrIay7xnZjEyOUWSkzmB
cn1x0IR7cEcVxreg9vTNHKpvx4eQnFQqTjsdhH4wBxXfxrKEUgiQ4gDsh+QYOfeU
qbQjof1qAbOr0Pbf1njaHxxANPUTgd1fAy6YUmKV+M9bqo6CZ+oBIqR0FSGjfZTw
356xURIeYeVn+X5Ixa+pQ2uoIXqSWACSmd+tBec9pTrQ8SfG4Ee5y5tKskG4kiNG
6wQ/KyNn/2MAHMwaICfioBV7ccPINV9gRAi0G1n/hvRyuDjxtyr9YcleFeXyxfVe
PhOBTqego/57lFTHKWkWiVWQH2FXRflEg7r8dfthkl99QLT7S7AJznyTw/KN7bU4
OI2apDnwtemq+1GjK60R82v6lLdFtyBhGAwSImZMreQJ3ZXKqshJQyHe/KxYIonj
CyqhQA0vW4jcbCS9C7lCPXN2PGDZLaPEILQ030O+Zlz/2E4Vp78fGSSDKzTuRh7t
r6sJ/6yR0B0ZezE8wUZ53fe9gnxrookyNP4KhDF9s9m0azNF+jCGnKG+zAvY3EK6
T3ygjLQh8UHIS2BIV0fhONfci9swc6xWgxR9RfoY4fRwkh60CDSbgRws5Ll1lahw
UMLjyAxNjAaCYrETcAQnztqqnJ93IZXCihRiAI9EulO6Z4pc8XIoSp/sIR1eqQ3W
nc93V/ivhgfxRoUCS6eRjfgquo8LgK9CMQ/Glh3QXTElchmPodJBezaWLqAqP5Hc
oul2auhNZ3tCgnAmIY0PpQ0XtOBX7KQlJd1KiUdueHVvbMsq33IYOCh3yxtw/fte
eMH0CllE+tlPMqIY4thheiDVOT+FplIm1Jaq6G4SG4aATSsnA05w3UsLb63Xd2qx
6ny94wRdlFo5WlCJPN6A5fgdWjQ49U8sIrJtptq07Wf5ns3fsrt0UzVz/+jUAAqw
ZIk2DYmd4tXEtlAGKjo/QjYYtS3/GNZdjef8OdEU1/qWp47oe+N2doDERH4MWWpr
OYrPQmM2POH84HtZkUwoKeto/01pd7tiMGfaKm2UF+r/7DKej9NkvjJa/rCr0fvL
Osh7eDd0V4NGYHEBPKvj9Rci67G+dAm0QAzgcdDl1Y8OfUke/PmJEfG3Eu6eZxg7
QKVh0AhffGRy5fm651b6fTjdFH98nO+fesE9JSyHLpb855FyiJVJL4Hew4BCl87Y
fAElMvwLik40C8O6woLLljxS8gN9K6IiZWODePs9T2tPWXuKaQW5bBKRsNJ7oNlW
anjIxoCN2BAz6wTS1iaXVOQiAjsGtDL/DLeN3mt/y++VJ2umVnO7H/ijvNmRnyiX
lvFd9Payumq175zEzuAZ2VLlDIAvUhFKG5YHsz4Y0MTn5k0MKQEy9p168Ba55qs+
XZ+RsTRBRViTolQRyQ+St2H+c6MlGruh1TuyF5HpIv+75eDo7gPedAbLL0Un4Oq5
51iN3B+/gpEr/ZDL2vA2u0lmT15v18cVw0DWGrJc5tIb1oVH2COJOcw5cz9dZ2ht
JBiHykxsPYfMDDFiDH9ri/YF0mCKzR03ex9BY0nm6sV7Hqfgv9r7KREuG8LNt5CB
+WQ1fvTaNwYj+amYDH92Kr8w8KXm6JXg1kjt+REhjr+ubQLcJPi/Yhb5hf5oboYt
DaN3T4780Gz6vs39AbPtRbkUkVSqZ2BY6tiN2PpaXtIP0S9j0oJG9YiHPdLwA22w
PD+3voPi/imkelOsoDcevypuvMExIFetdV82rf3ca/ldjZ1Di/f2LlASFArAzuQR
9idCypD6a1mYqLCoziePMMaftUCjJW/G3gEW9mHFal4YVQjtEnY+7SgEx3/fx6/S
HBqSM5Dknu+bg1eL+sWS8HxJeRV7652XBceYW7GhD3u1H5wNs8q+3jALMEoeywHT
oGJiyq+h8EwaCbDBkzNuofakzuImU+bwwYLiovRYRRcDURjRIqUcy/e4J3cRSioj
2IZgEbvJLgBru5ayrKlrbX4+TSOh4DeJX2qvfEyT0PDMfaPcnPqkXxpbKYBRy7Fe
qJEaYhvStX3jiAwpT/X9ADo2q9ydZNZpPFvLysLSDLgwrONr0RDLt0TOO50FLQig
OPSpL0afkZQqp3LAxOdUbS58wyoU8GizhMJtpfmHjCTl06HmDLPQQT+BZU894ct2
U2yl2Ty7dPEOexSQSfq2gcSmW3UBdVlxYJDZ+LIEO8tvP5TzlciH3Z5+t0yrSMrl
F0/Z/OMn0KtJl0mu6Nr45dCBzSMK0wYBu91zmyECw9E5ktk91VTJsdEkBTVbr9jb
3Xw+OEcm1ikkN1OfbudA3U0FuuPiPAUZVL0g2DWV0MTuWUPGSt8ZzzVDVTaQskr4
O/aWAUpi7gnNwCEezGL9RoAeS9ZPOO/SXDbqFLa/0F0r69i6m/8CYSUqqgjNqN9+
LktTYGRNg56w/AT89cvMRQgzKPjIqFwzQqTElf1jk+aSDJXx0dPJ47jqA/kBjuxF
f4iA/Iq9RS5VSBcxW2m7eWzx2j2UcRIzFW7l3+bPTcczPIjWy7sH8qLd+ihjjcHl
+3dSgmGDWS1Q8Mwj7eJ7vkY/uAwY3XoXXfsAqSgXVR8BDUvGJ19uek8plXnRlgJs
WjHjF9s3a2h/ORCrTYFCoilfifdKGeX4B+GhapF+f6l6tbIlzI5R/wzzsXro2FOJ
blAnaTj/OpMrlO8d76I7ZtKlCo0+7yKtYyhJ2CwpKO4e6K6MGtyhqeyFvbluALhF
Xygw9tz3o81bEAaWz3KQWKATLeWp/K7uymvrFt/PsU2yNCvBn5aSSZY8R5djBeFo
PtELEw28O6lL4FBCDXVqxHIWwOVdKJLWkk/bkKMsR0hbMubKJfX6JqOzzLmDA3R9
vNpUEQ6icGcoTqm1PhixDvAZUctVMqa2Rd3ptTE9sWBLamg8baleaKfBbLSqys4J
A/CSw3I9t0nXUGkv+GCBqcxOmvVo+1KNgAjUXwrXr1DqttIoSVC9we9nFrYuchSY
fpakx/8Wpndt6bO/Q5c5CIKG+Nlwno2glfXtJVJKBSwcnP3DJIVU8kFJZ56tUzxP
oyYx7ot7uz6mzfMA6sIa0nWytAXH5Wi0T1hQHPTceZHFwadcPnQeqF2XljirUIDb
F4kg+CTyLl82fzez0jN9j/n+BNwYdvKacKwg7OLP3PEMD0gzG1noGhLpGmEucVDm
PAR5Uy8JHRFXHqrfxH28My4l2J0WOwSJ5FT/Dp+poiQi36kx3B3QuTKL3J6CqaCz
YP8P7Wi0hyhttYdj8ZBKlXNvGPR4e+ygOvffYtT7WaI6cU7svuJygUmkvKwAJrCj
3ZsNT6fx3V+xpN7Rp6pPnfRORFMcuc8em7NSiMZttfQrzaJGnkvfCM9iUzaQ3nbS
8Sac/CSUShET6OHMarPd7ajeqE0I8JOklcLxZ3rjBRxZvMHJOqyT/ZMgng9pFjFT
qq7IkqvRYoJkPH5+BWVZ5yK0PCmRLiQ/TvePE9qN31ttrFZ1sRkGY2napOsRF1+v
zSw2CEIrjRaHegEVnVxjqMsZ8ttVrUlDrqWxUddRWVylEA5VfkVdZamEUOQZh0fO
fVklvfri0vjQhdJuTEVjlFtnSiSYag0mugFkc4PeJ31VLkNY237q+1QAiIKTstjh
iYT3qo2Ig06s62I7bsntP8Kg7JOQoTY6lXl3SVFiKdIZDDPV76Sk1VadwgX2ZrH7
Bvz0LUuBr+HLMvbGoFJWOL3l4eFltJk2SwstQaVeyV4AsdWOrzO0vKtLedFn04ki
/ybyZMAoap8T5MFxeKtpLx/xr2Q2UMuZL4P0Mpn9v4h/4qR1eB8KXiY/bE13Yd0F
xrreZ/PijmETQ9s8Py5xYL5q620gygnEJoaLjoh9SktEw+yPJVrr9rpYThgHSgma
ocWDphU/sLqEPaxgvDREo3nMSIrmVYq7172/utD+VwXLUPAqZDkT2r3yEImm1+vL
rtJZeIpvKpagHXmFRkBoMJWdEuB0vtRMDmR9Nl1b7i4qeqgDXjQcK/UE7gmwvq+U
IFcNeeoemhh2Y0hu1aTxTTE1xOc/j+Q2nCDdjltzX+G/2dTSJlGMBJcnULRnqBIX
EbGUsDFOrEe5tPzh5b29ZFPwdcgNt5XTQFNV0UcPzsIEcE0lSWhNRu3HWZPeRwOG
+s1rJV51x/mzY18yV56TOAhA4+kGJP7ztfOnMQgnZectfmVQAjtXRqQo7KIZNhFc
Utl94JAMAcmfwvT+eiyGVIshA8n8gDS4+jBfXUR7Z+/IS8gEeF4cQQefF+qptu6s
gFjWSzWbp7YZmDFqorWNfpDDMNPkl63XTF1GxOkkwyHcYChGejZP/z1iyAVSggyL
3PxEh6PYeBbiafH2TehE5kJeZYdw9HgkRT9JFYQQeRv5Beyh4f2zFhFA9/2cJvdr
Gm9Za5UihjGdtBjxrmd7q+C3ioWSIGgTQnqEKBY7QhM67pWbFulvjT7s4n3HBI01
sl53WzUslO8GxAp+tPcs7BdCimdyF6KDRUQEU1hWMbB7ZsJNGBuYk2aHOZcn3Ihw
JPl8UpHmgDrIbuFdO43CuOOE+v+8slxWP5HChxTnSAcdquGQYn1h4JS1yfvBwwyo
721kdoOJ8Pn8f6JhahImV2TlToy5La5J1qRQMIXCwf4fQGxBvH8Yh8p1EyPIyICP
Q3/MoYAxQaQB/4BdNm8YToc8MWDPnrq0v8rnVpYbQyOzhHoAPe+iMFpHjXpfOWQw
r6V2JPyxSVxaMF8j3ko8IH5xK8oeLiHh2ATrPmQrJdImsjajdmimhPyZ/Qjtvcxa
X74jGATIO10JpvOjRbtkdFC+qLcJEfztofq+5f+/NMM1fBPue+eyX7hFP0UE0/sU
D4ruEAj2OS795vz9rZ/KO2zeoAl+/N3A98nDbZMZDdARDj+mvinAMoqr34ud/lzX
Hv3xzm4Zfo9MuoYSc/88lZipFrt1+3Hy2xeXUJhVnNnwLIjl5IfuNa/LM3AsSlKZ
T6aNAt9oP4Mtav43m7U2cB4PaTVHhAdPhDIDx76FM/2TP6VDEcG32+CnhWDgEt4/
AqJ7FDigzOX9S4cVM0yOWr625HXRDR/6XewVZnNcwZ5/yBlxht86kq2SKb0qaLgN
SRn4rr03H8k6kbKXhN8TAbGvtR1/KLBCx19873PTVvFSu6zaZu9yF3hq2jN4jIwK
f8ZZOIbqKl92ZcAHNyTDcZRwoikFW8nO95T/J97JxVjVpOJbrZ9f8sD+f6mMDlOV
0bao8cyDyOiF/kco4dfP1jap2Jf7+AufOVu+dHlAtmx6DWpWiCP0WmfkvQ/KlQ0x
rY44PtNiyqq64LyFhyVdliUcMhBVYVtZAtxAKJzyCt68eHXs7FqGdFzaX52HPCaR
DfIQ4Dlp6LaMiOLHMq57K14CTadJjhuWm1g3rvym1/pJWlYaqo9o+d+dVibqsDH3
7NTshrpA7Sh7btwOnPOc4c3xLcVI0tF9fbU9yDXVDuZGrdxHjVRxJs4wRDMQ4WfU
nJHN/+1R46VNd69jheTG+mZiN3BIa/t/uxfNCWyCtcme6KKR23JmoAfk5ra9gMhL
oQtrJNk7IVAonNzxMVqZT7rwl3GTeONIIv02ijrKEVc38/H1z9xuijAra8xqnPQF
FcPbWE1FVpu+Tv23CwUeEPBDEHxK2FQX7I2eIPLEP9UXfxIuxDERVfxoQR/DJlv4
sAXtUGae5lO/koBMGNrRf0RLuho3a5/RS1lkjNYu5Y/pf6HeM8dBJ5JNPcS+sK2w
Dv1r4smHVjBbi+HhF4RQk4In844IKWI84g1ThGjpps0uC+bPtLPv9DO463HXNAp2
i2twtYXcryKMN/d5l3UhAcmueIza/EEptMFbs5de/NxJzhJscpqUEyco8oP3JJW3
LFY8MT72WII2A/15MvSW+J67p6fFj1b+OadkMJV54e9YBlbk8SheSaOiGms1CjlA
aVfyFXjBT64Sg7YiYvtH77n+bpXky/I/Orwd7xhFimo4A9Vr3gLMNK4TB/BSM8zs
+yk/RobcS8d5qLD5cFMP19A+qf7yDeKv0lxX//L3ThS2NRTQvXmENfDoWZjt/VX5
ZeIad1s+9VAd4ZS4Mu8VSy09cMUVyti0m0KLnBiIddmEYp7zGqlO/e1aHHEKjn7T
mmW7OKkEFB+bZI6WqmkjuYGGbmyqWospG/JDYlxn6k5mXZvB1cjpoPTFEKov+pRK
77XvTglxZTkQQ1gcoOyqdEq/R6hMQyDRvNykV1lQZu6dOIrIprDtMTX8VzbB0d/1
vjoRKzN9JGA6pc2m+EjxfDopkDP5xiZ6GDQQOkl1vvECKQLbRPKfgi3V60JfELxc
k0JlrB2zjQ2PXHsNsXx9a2dI9QYK6T7Oey1Lzi7jRlQfJe8C4ANWXZ2bnuS0g+09
p15rs26APvteU+L37zb+RvLb3SnnqbjflOQ8TcuIrxem7aHSrg57WYcQZn4Dx1sG
d4mDH2vHxlqY1UXy5tLaR2PMYbCmyb66nFJGNN74khviHHS2mvSUmjhZT9J3GcgS
/kSyQOv/RhmcG5oOd637pkcaUYFFPJ8jyXyr59Q2dzzuKeyKIV2t3WPBqoyMH4Xp
bQgYJlNiA4oZ8RTaKeRwzPylzUXd0CSmYB6rIH0Y3dEmB/hJRPRJs2idC5Y94IY/
xUAmySVGCLr7ojTBtXEdLqQCs0T/IrdXq95tVxC44QF0Bujo7F+YBjVv0qSE9me8
TKQRDpEXwDB9OYKACGsM9xi3u4fCOPymnpndUsH3epm+lgmhVu7FfU6WzrtFqPD4
KaSmIZxjh0ppMHmDn8vbCK9hrkU4LTmFpqQNJhyVxtTD5mCf1qrHTcGXTbvMbeqD
PnjJ8Jf6gW7OFVh6YL97roN6w1e/UwuZ+EYKK9sv9DeFR1+g4KONgeyPHftOcZDf
DO6n4sUgKf8XrCQSYZRiKFMeMbSQ3xUmSoX6CwqnyXQNxaYR7ImOk+t7X4CfHamG
Izquc8CEegopGCr2lral56oDOFIdqM1ouHVM2Ml28g8YZLkqgl711xIxbYKrK5PG
d9ZysoTWmMB5SDKmIijrefgbODI2vHsFEPOLciQzbJYwHtnw/IBcUgPO+Sl2hcWp
rEJ2OUIifxsUWskwrmcjuoHcW4exy8rZtH/Klxr0lVT2UVd2PwXkYOJx10AM0HKA
OkQCgSwdJjD+NpmgE2oP2MiLywgahCJ0C6eMM564IEXUZkxm9TcuFG8EnPS5W/bf
7Wmcd8Ec5Z6+HTsVJHMcr9/COmTDM5CFivaZsuVQkkE2bVnPppuNUwJePT2uolzv
HJ5JkFJmfG/idGD5yG9pT6eNrvNLoLhiD7qcenrsrE264cHNfdM9sXJN05Q96evE
XPaLXizg+KwUK/jqXOG6VmthEz5AE2skTXW1972q53JlfmSWVoQC2miRlwo3Evvl
vA5pdUrAV5DrHvFd38IyhFJX+eOUpx+3lNnj3QcdbdqE8Pr8Z6tXUyE9El0YfoZ7
dW1pSmBovejHPVFpz3+3qpWqVqhCBj8tiQzbYAbVL3l9y7QTPP9NZyFBInj7h6Au
dwqVwRv4NFBWh+8Q3vWZ7mYbpipsynOhoqcWoNVd6NCGDCy/98ea3HEsloEXvc0F
ToieR3/Xm4yYGpdAn7YiKoEJBKdgcz/+ll9e/BwMUt/65LwYlom1JpOoC0UXYjQ+
TTD5UAq7Z30N7yADjOMZGvvq31wDZUQ3qpNrECBFhpWt4uiiAFnd8toxS10pcLmP
wJVYS1x17i8tzpaeagrbj0S05rBx2L+V9tvtra8/Ro3rPr+Bp0lDWGcOh4iawb4/
eWeu1WorIEnBwIuT9cZ7uMHoXQ4FQPa3T+g4H/Ye/UjKJO1Vh+g2fKAZNbbQpJFm
Th0+61xboZ0P7x53uBM/+IqWt/p7d9G0iccD/h/A9lBSvHeoPv2CmSGZ0Y+Hirc4
Xp2lQTuBTBgOSDGH7RKi5ARJueAhQlazhBVE/gOJ9hh4JPd0cjCUKN9KvoyCgMA4
HAlvYY2IMX9PvuvEZ3s9iFnJGfJdfkF10pkNbDp+Ia7CyYeKQEtaXgRy6ykT7A63
RgwEyKUTu+oOSjk607bNF9qlmv+UYZOWsE2YyVasI+ZAssO+bsOvu4QnPYxs9eWM
ZGKJK4I0SNrwz14/uiQFFjXUdf96kmSjQ/qEAl96krnPQ3xdIepVTG5rLOaWkhGm
xDamZW7D3lz9YrqdhLfniyOHnSZOzrkq0S1zANfTlfGbQJ7oupX9LQRNy0tnBUhE
WMhckdCSCyinM+VMIINB7EGiYbXO7/WU7t7AgiBOSQh4v9ZeF6bS4H2E6TIIcs7p
zbU74QgJSN4+CEosumtZ2yk2Itry1+ei33w3ouLHzyBNMX180V7pDHLsXCT68Uu1
MS+eeWaLaoimLkbVrOWqpZO3G6MRxPTnCrAn+Ngw2Qx5eqkXeswVm4HZNgxzueZp
GBO6emHYd7uAsxAplfiUyURLxhO9T+vzARZ+B1LjP5CPMHbHRfvNQDV7HvH6V9rN
YdTH1/8h4m8b7RuSF8z3AWCYtnltrr2obyQs5WAoJF2xlzKp2cedAVq0yfre+I24
ErFV7UbWQtOsff3ZbmZdWvA73Yps7bk6NwTtVEsyGFzimrE6dsWUQ7bDN5GoI7nU
vMh7/lcR0C8ief4/qjmeD9BmCFCdPxP0aaajAHtqnWZIv9/pj4RIoR9j/at2kG5C
ms9wFczWCTRbS6vF/qblh7hvH2JmxTgi0z5jmHdAvIPt+LDWzdc/2tjjYCNCeIBs
co7HvaQqP2fGNFYG1Px4tRJNT3GzerWlnlCSVhtaTt2HdV6AR5c7CpQzlzWzJ4SA
B2Om+mkDQUoGQVSQQ969CfkLou3yjnai6RC+AMnfhncxxGkYr7Jkov3/Ijcv4Ny0
OMbtf1d5DGWd37IXqrvghlW9kEGFVOOeVZ4M4yXYSulqwSwUab1CHHUwPSd9lOy3
vQ5Sg0bjq/gjfsNRMXy6fPwv3wWHFfVeCAmDAMtrTlAM7btU8lfAPaC9R1uCJI0O
IRRk7z5isSk7XKnMdc+hlJvZaUCCmIAvVM3vJxtvbsOcnbdgfWkl1y8rafFTnGZL
sveOq/S05lUqQ7WJw6IRuaa4MVf7NWdYp0wZtsKgzQ3OjVJDhBnSKQEFFddPV04X
vps1D04sCFh344BHAmeBS3jW/21ZV2kQi45v6j3KMD2EaTnGRX/FS8U49vONSz86
BRP8ln6oOWd+9nv6PInf1w2J7nWtQZmfHndGFJm/1NZ2ntgN1Vs7Oi2x+PGI49XX
T1hwjB1LEx7CKJHSAkmCPSpeAgh3MqbkKDn/xdPeRPy8rREr/4jGtoK5fz+lQm2r
FkzW/ejOYSbuOp6Ga6pESfXPstvFk4TwuaCsjcfQBdk4a9nJrd93bSebpZjrxqam
ceTqXwWvd2sqToooCqfS6siW1zf2rl5vopLQ0ZS2Wmigze3UIJ3QjRQeA3XT4d6o
XadzJGUGb7jJLc7MmkLZYhYKb5oHNO+3D9/OJnW8bO4N8HYFXqNGlKNTcTYppLyr
Jb9k5cpd6qj0/M4/DVeF5E0gainXNcze1bOPzfJoxINuO8Z2yDAl79JJmT6EvlFV
N8cpDC2CE4TMY/Eqi0G15tAGR7Tic2vfvBAQB+YdpukLYwjTmIwLhGz/jFrhWafq
mx81VsTewJ7qEREUoKRMr2fmTkx6wtLIV3EH2wgK5cjkk24BkXQLryFpAYFbj2aN
wQto8BCl7xLdyth37WTaXqFocU9Dt3UWSix/FUGSJKqzy+voJqGKed+6RlP2Qy7W
xxNgyyfykGKb0fQvbabmnijghEvD+ATkYJtGIk5VDbnj82s/bB8NUzRgWjIz/PVX
dzvFbYALA23hvTGmxc2g/pcl1YXfJ9wWOb8VTf8zd23vBmr6bZMon4KV6fTkjUPX
tQI2UMEMIQ89vg96tZdncZXNMgBaRS5URC3aRd+me6VHd3xxtMNYJWeLZtw6EfF0
royB6Qc3xrnXs8K9yE0xDVIPJLQsFiokOaB8TAwvtJXNoApZH/D2YPXz0rhXbVvV
D5rItLjwfQ7Rxo9emT+zHodjLYCAN8gljbf0qm5VymLPeFAs9mBrSb8Ns1/K89RJ
8mKxMKuJM+BbsoCqgAqr2dv7mkp7ELZAC3iaSQZRWT7otvQ5+Lc7t6uaMnbGsrS1
6CQy1St7rG8RXgWUM9HF0qW4UqEGbfNgqxXdOAjFb+dEe7dL9XKmHJBbZtPmIh+1
piedNowPGIFlpJiFjAaVMcOf8cfKoW5W3Odp6n8dmgVHQ1pd3VL484qmxds8Kod1
wvAJOs1myLSpwpNzjTC1WQJ6fJKuFdSb0ef4dGSFj8PntHh6k1Mxig54Y9uLTi58
bq/5w85znajpT8Uxae++PZeFqs5RpzbIuP191iSw+daCO7ARFNxg8iLJVC531ApJ
TvhtTaEDIVbquIttUrr7+dl7qGvWO29GifVOKFmGzvBGc8hlTm8EpJAhEF0iVyR/
O9YCLvWOuzIyFxW8cV75A4y3WFR6Ay8ukxN6MdwDF5oSl8HIuy8JSSiDm4lmhlqP
DBM0/Kqky00s8UmQtBhXzNDsvMuO6tPJv/SOodQtJuxEPrhcA5FVMG/r6moasvAd
hcH46qs4+2rmHfh0beVfJ1QZsYGowxIPAeDIFOeohCHSN+B+dIm3E8It/TIdK13z
JifiEBRyU3pBnp1v0GMWmVVmmLcYt6dvV6JBi1v8QuiqjcWFLP7fNXe6k5Jcu/q8
20oKB+JCvEEZBbp7+c4XK+3Ljlioemk2FmFkc2nO9dLvdC506uODk96NmHtT6KVk
qQotKIFbR3gR4yLKCeGTZTXDL2WiPL27/cUV8/y6iPHBOy26whQW47tL8jtr5pWb
53GO2LnxGbgYEsZsGgTIeDvflTqyx3mhO07lDiJ5NtrKGsRHnPWrNpCDC1vfwKOe
mqUAMUnniSwBwKWavLJuVo/P38qL/4RM/3B/u1nVvppXfkKKFPLLdDVwD8McHSnb
o3Nuyp9yh0gTxVvy3oOOLrDicHXSx1AOMw42MpFwARTit/kdKnchY122FjpZzAvu
xYvUoQIZm7GZEqUb2PNPpSk/ZNuhhjsS3YTP+APNaGgdHkv7I8bojNnEZHXDLnfn
hb96I/KtAZLOEu36WuBHPXzKoYDXleNbLF884EfszybRyEpwFSL9yUL+63rxNK7h
vrv7a1tjJshT5uSBzb0Aq659jC06ls8cQe8v0re6CBUUkqnQOaFtnCVD1axJ+min
NovhDrvqnZ1/TbzLuCirYhMTMxLdf9Nwe8P+oGXtVCrOMGHseQczJ0s4S1/Ficd0
9IB5UWf9Oiz/sKQQwjuviIdqtzLgfEvQjkMPz4nggLGCtIFMuupWOKOBxJOzmywv
BMkRNkKsN0ACgNHv6tz6BJH3yUluyaElcAfJ3GxD98FBTCKY4ZyI/H+9hXvygYmn
v60T7DuJ+dbkldHoNpmw29pV/ktHjzBTgjr6VbI5s8Pycn5uSm+3BjocHg8nCkPg
EfrFWD2kdO/ad00bE7/q6HdfK+wKkn9N9rynBGV4KJDy5a1uGPZY+MlUedlf2sAU
/sk650079VamLObMKOeh/C2yCqWeIlypSdaT7JzAoSp2PwDD3Y9bwAJhAnThoMQk
M3yAngSdu1t7Uk+dOzwL11XocgUxX9HO8Ub+wzb9IpK14aDRzMIGG45iXgwIEaVs
7hg7fYCS2tFzfHyPcj8u7hECVO+FUOt41cNPEJcYtmQBkZlD9a2u1pMQrs5czD62
ny3/M/gdW+1LGAbTd6JmJSZkusWqcegPXZxE3OJGHBe703Z9Ndby944AbnSmmyJh
FqVbU8ov4loVREBKdgproFUdfkVKbCIoavxy75Ow4XNWAfiyqSDX5VpjXbAKd9ML
fu1j0S1jgohS+nmk/OmseRPbkqbr42ojv8jvH8JdZiiC6qO6O0PBNpm4rwB+lM1O
Z5lcRMdG1psyXJyEVOQcscwZ754+OdE8cPCVe0mBSIAdZ6Be6REvtCIm/XHIaL0b
scKNw/3k/dPCdQYf4ctEEml4d7KPivpsTbuDe9wrWh5eZApGIi5iIB6L+a0KzGSw
NnPvhsioTlNpGlKo4v9CSZxJa+E9sQNMIlLcyP5yTYQ7iFabAsRarzjNwujvkGxh
8vkLmOPi86vJh/FKh3yTgHK4+wxQ+E7EW+FIBMnt/1AJH/Xv3swJN119suBupw1P
TkK7gwzoIsAfeCj1s1PuCwHKFhJwMzZl3DT5WevY6X6c+9TBt9YSDHtUnrnQHPXz
XxAgaUpmFLor8HTyKx96eCDv98vLO5PEbJRuK7Xv8SwTS/Laz5wUTSVPwBERXG+q
n7AM1gTGRByk4FZ+R4d1f1jMPDmx1kpFDL9N/TfqJYDFIZ3LnUiEVmY2BJ7PaW33
vV+3tJAnhHi54/ZVZSbOkKLzAThe7ZeKsivrxXXjdjW1TodYEfgV1+Ibx1loKgiB
DtkLTizPNp4R5vaZEwGRNQQUE9EQeRSyHYMMfn0FqiJMS7lRxFrL+s2Ac/Y3kc7S
1XRY7TFnHsi6TWvVM7g9qrCzpRHG6tFsHokxa+9+ffKaaG/yHOYZqe62hto+ZF+I
Fj9ghR0u2RGNVO5B7TzvPohcop8H7jvQtzLPDn4m9Al2/QPhiFgMdF1utcDpo4jp
7yuDGhSiYB+9AA0aa+P/EbIGjyQvhrRSrA/iTPM8aTvyyNMRPF7gsaOrPSGDMH25
l4LpEeJqieOFMdHFWpFmESfAc+0mNYx9Nnh2wB2YN1zLwD+ojxPkA0G8/dwR/m26
Um1G0Q3jQGJvT3YISZ4v/oS23m/3/tEta+xXlos/vgT0Xtx9WpxCS0RCM9SctCIl
SG58W4SuB/eQ82hpi0cfGWCUCcqz+ha221TELyKJHLZQPOSTNpX7qw4weSwj6wLj
+AvLZTFDA3+UKdGaZUsM+UNxSksPqtaHG8UGXyMSoP5bc6ATDi0FYIE5svWn1Qwm
YHg8I1/gKVXUL9vnfoj48W00OCkAgwUo1j57JRgNTB8+8uEVw6HTOZBC0sca9BkZ
cvlEfjBf+Fnz9QrceXilCCVxABQnlLXMCY1SWQ3VvRJU/YUr1i/oBXNdUhkP6ZGp
QUk92bsCHkrEg7VJeWvPkROHDjdmPxh+EGeaR53ckgi5Qsqd6HS3COs/CD8kC5HB
ZRiXY6SWjLnfTrgnioaYasn2UhaWAIhk2th+YIkq0m0gNkH785YYqqviGcHo2/h7
9+Y0/doR1mnsnjSQMxaIQ6BQjG3gAryJnI4OyvWTqy5EROaasU+L9jLDU4JIcsir
ITCMR2qpd6XHY84Jr4jmmlXP+qUQMl8UTH5A5xUuyIng0EtKTlMg2VkeVF1vsAz1
h4iS3MqaVgNut1CVsoDrB6Rhg/mmIkF2j4gZ9uL8y51zJQzTCCas2SXZs+gemWUu
nangiKWfAHuLwRbS+0wuDyv0y+IOynJKd8XyZUwlZNSoeLVN9FqJEDusuFpeDVCJ
u6SlI9yiCXnKrt92B/mLNlcBb8I7Ll+marBgoaB410i1D18Scp8DXb3vbqvii39g
36cO7QbmUK9ZfFqLihWAXywnPMxkPEfkHzUH1IHvVm+yQo/Ml9ET2dgr70i0+15y
hmUH+1QckdBPUlmUxk5J5aUu0VuRfr8h2cP0tHqQaKuxJ/FMYiPFXOab0YL8XuVI
Gy9o6M30X9IhjlLor94ZhdO+1yGU/3A0Rfe0iyC3j7UjI3Hqhr54BfmAor6U7vLo
qXf3GT4jHeoYxUSuNBMG86+we7labnsRf9IuYFwGKeaLmmwkm/kvx5dVndHLRVGK
8jjoxwSjHlmQihEYlXKp4yhicO3HCWw6PFRia1Lv+1WqGdzMgsYAFlAbvFoVy5YJ
HEdzXe3y4SgGGkivRlBA9mlwXxB/knZrbTDg4BRJBY9BmRT65iw+4ZBtzTMlyvfO
9sZAJ5D8ivsDZccKX1oWt7SMFlftg11y07eV3m05hHfsGCkb09FuFV+MU5NBWsQY
mSIZxNVN9X78/ZH0S+hFE8FOccZgjKgGVibLrlRLp6l+l+DLbA/khhWw/m82IHoh
EAvxnznSoli4qE579t2YEX3tzvWRRTh4iU+0Gr6PVoE7XwbVCWzP+IJRhj6vtN2g
VHzUgX0JqtGo87IHKnnSy+/BcUY6Jny7X0gq4bXgMAOr3OoJfrhoFEbyxTCHjFiF
ASOIRRGYetQ5L8DRbry0Pz61aS9uQsRaPv/DhYbMwur6LFRiIOKhAszO/FjuFavb
kzDhMBOpGlj2D8rjPD6PI72gh35YHoVsBjt/8JLa5hsG5eq75hjPXP2pLgIb8xrx
UaZwjC2Xsfav1/+c4kPcykU1YKpSTzOAmwuxMpyP0YO7ROsNzkWN4gEHVcyf7GdF
ANytO/q4Lut3m12Q9Dnbez5vr2QLyBRHkuraxjwG7UjK1YPqL2kvXV9i0CHgsi4e
Pk1fzY1tToOioz+4Nq5cg+BBsHfBlQMMVO7f6plQmScApuCffaip+iTADF79rxRB
XFisixKPjsUjKp7migipoUSVht5bhiZzcuwPAnjGqCKaq10sGZJAySdkn9n7MNdS
yiECUYNSEqvGQtvGcJvxd8eeXYD1vP/2Hqmn9HD5LxEDzDym6zQVHpN2KB88ESYL
czfGxa519Vel/fdu/43XMQJaK5Pxxtfdu0CNb/090WdzG/+smRb721Ww0ZTdMHtb
HRoaIlXvFem6gj5U3a4Or7BUSxqMqR+ba6MuMwgZvfiM6X8YZrsY8cKkNdcZe0TB
DCV0kr+JIMTG0o8o7hehEP+/cDUSJm1+YtrZygj+tyG4wXictYLCAxBBxLE+uV3O
UeUN+l015GabqkyiLKIOHaeYfxh2Vz3wRe4XJ2YoYQM=
//pragma protect end_data_block
//pragma protect digest_block
Bqgqk0MLUFvQvdP+Pxm18AVlgLU=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Caug/q7GvQiWGFHZH4e5i4nXidUskr3J7r0c7T6pNhlpvZcgvyt9LUF026iDcH6Y
nWNDHtxdZaVJ5U7S3HkTdmegDMzwdCeKcFfVgZmqMG2pjebJbKrKjMTUwSdtNRLQ
uG7j3Q0PYJGBPMv0VWOMwXxsQ7Eq5OVIX45Rgr03KDeQdblabGp/Og==
//pragma protect end_key_block
//pragma protect digest_block
zyrcYbMyBUmnewwoUeykySG6DTo=
//pragma protect end_digest_block
//pragma protect data_block
FW58cL2MQWcMOoZRhrWod9wsEI90KQzTjO4nFvHkR2+XDnVbT9NwfLX60GLLvsWa
HUmEuvwi58fQEgzNSpj+Au1tz3oU84xxSKj7U3+lKAHBD64ycAOiSLvz0Lkq1uhD
VIEDsDjo1E2p2HzVgpvqLFT0r2LMhU0P33HXGI7aQlXj6cfjlObjfQ1sQhTZX1fO
wYoZXIr5QHd59QgCVghCphPGydshbyI8DsNJ3Gywlb4MZXqiaJaYRQJBqZWmQP9L
H+Dk1w7A2VquxKSCDBtUUXh6FuIruJ9PE/hgFIHSNRfjGKx8ggHAgBihkFa+K2tL
DXu/Ck9upquzG7cqmx1RrGLkjnXLse3BRX8+oEsYNmARxBy1w66vWa/vJ1i1ZLq3
7PrFEkh59eofTOtiEHhzgcNJvAbalyJ4+vAFiCQtR5IPuYivAvq6JdSOoeET4Sdo
SzOKinFhILfTInqp7bAYtVMl1bM/Y93L9mjHHCCM7dE6VLyJK7AeB1UupSfPjiWd
49Eld2zhk3+Zf1yr7Ve0KwPsu5ZHSkAm/nMdJXYRxwKQY9/9IAiogIWyv1jU/+bR
5UwAEIoHQRYETRjkUt3IxRFmIjTFnDeObZuR7N7vcvDYO24SJqobUCvDY1i1thwO
sh2AttfLE18yXZORMkFiBij+eHcmLwnzR34PKfDWgLz/a45c/uVHSUpQmMnty23K
U8akxcRqGCUm6Kls19lcLuSq+hnLYvG/mZFi2o27Y9XLGplL586uqLxxeKPyRI2M
4aQUnhrmtjJ7PKwH0bxN8+aLvUlM0dCGCYZWM9sQC/hmRg2Hxcbs7KBNqxM0zika
UkcDwtOaYltY4/6XVS4/HOj3HruOGpW/oGxQlzYFEm3EaErOt+fMne0FsUS2wds+
XZBEy+T7m6itV/dyc9yufJq8dJtG4NDYvQuyJiHo5sTak/omD3Pl9wJc+CJ/QoA1
ZOOd4++pnr5G/W0+wUQYg7OSNrOL3e0c3YLUe8eGM/MOTf1rUaIRqjGAwSa6pAdS
K8Nxr6xV3MlDNcAxk85uZmQg27xSUUPLIwds+pQozpoFd0gB0ObdFepXt4fIqjU2
m3MLGIX2SMwQzEb2rSBnC1TLS7Y3rAUZ6Mn7FwWR5rnksbZ9lKFsRYbXNn3B5eMb
vfD8NRIKF9nReYTrAAEBzwdnnhm6KZqCIg2cJPFOG9zGmgjvvOQJCRbqzoedsRqs
dBQfUgOAVbdjLYxS7dyLhXdziR2WjfeFsIcgseZJCG1MLVFazIEhoifeLxO4db7r
zR58G+wy14hTIOq0zoGzFP1zjNTk2yJWIUSMLW0ZZfK2Cm2ijaZ+yZg/WSSPkkOz
KyHZtIEY+n1PHYrCwcrRqOG6Rfiv54yEpCFPQvJBDq74iQDm5BzG5CJq2NgtVFk2
mlBO5MWym5LsmwVhk/rEgbZoGQRDJmNFqhYZRwEfvKYUAJs9zntefptRwe+TL4M3
uuBsm2TOjrFJJcZUj0zyPApid+fGab6NekulLL5W+UIp+yHmDj/UZo2gwIn1fPpF
orHsb3pOwOjYYG2hNuqDlIqgtrl1p4e4A4Q6v+Wbfs5biLqrCzpCA+6sqqzRUfpi
v4Eh23kL26M18XD4K6Oz4S3kvbZ2UHigz0zrLimoSa86f+wpDX1DwBmnKlFFRMv4
SQrcNifAqUw1BKqSzWvYG7IK6l+D2RkYDt+MxEr7zvClsHFJgNS8EAb68QbJRhnZ
QqZmZ6/6fhW2CvygmYcQdPbae5Eh3O1fQJNeN/08dg4iwz+L/UZ2BllY4S9CCXDI
WDOudgeE/rV2tZaqUhIJ8WDRSk1UBjqnB0+1z4vBVAzhbtC/0JL647MMwsvPGsxN
KGaJi/3Zrc5yaxao5XEW8i37vZGMLTyvwuw2zbPbF/ENFWqsYKCT9hHDX/N83ZB/
VM3raVYLbVTkgXZiUWKo3KQ9sCOduCTSwAs5CbNeIsabu03xebYGrpnYLIghelKx
rqfcbse4GnfhutPoR1i3qVjL5+4tL+gG8zq6mdjxiKehp7XA38hjjHxOVGrDZOvn
l/r3OHicYUNJPZI8IYbZR6RPIbj9qiIpQ+H7YUH6KT0Cr6zOyPr92WuWZaKoHnzf
TV2gDsTJQFrViVARyh80XkzOo+db1Y2GnUiGb80HYiuyu6Mzj44zoz3YUHL7TlKz
U6nDFZOUXiScdm0fgqKWPCpz/3avQJ/NzgQ/cQ36WsJcrvNK+9ias1Tc0DSJ7umZ
A6nTQyx0o+IE8f0xoRcr1GA1UelXGawm4ltgBEPQySHjkkxwGpt7lc5YT+w8uge+
XIyG3BZ8IzKXPWlFYMqWSWQapnUVsQSz2G5l2BZbDSk8XvrTHeVzSj6VKbtA2Dd/
DfnRUsGnDalnhxfKJ0pZadDjZhQqZlhzMKfyPoPZKT+PL9U+/X+awdBFlyLTBfgx
BYqssxF0eKjuztbabOE9XXdpL3z+r1aSLobmpGt6oQpaH3U5NWro8UkHeYpo6/m2
Tvm7ChTPL2Ismg0n5fRK8zBlOui3fa/gZ7vUne6lxQqB/3iNfapY4NAG1qSwagGw
0XRfY1m0dvwU7zN8i5bpOzQ2VN1x3MH9LJysQ1+8bPCTTLaHNHo2IHQ1XuQarBLV
Coee4T8cuu+oemVSSOUrtzdzgDtburywZfA+f2y29oYeX4v20/hJ//cTCbUfMVwb
LxUQx5qRLIDMqTylwakhSzinPFr23laxJTOcZ8zYBDbodiWz+G9L8omhLvPa5SjB
uUrIvP5naya/q2f7zmvZr0RJBXkUWP9/Ook3GEwcZ68=
//pragma protect end_data_block
//pragma protect digest_block
gVqX8bxPTBb5ChtfbAQxa0UqftM=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3NRXrZOwQem5ExdfI9QY2O7R8sNnnIBprUpYaM4wdqmGLQoev1OiurO7yKzJtyhI
MoWpWlQXrXO7r/7KRA+hbvT3KGH20jP3bYco0W6hHDGO4hX/aOlFGb5cStGDQkee
x0MBG/yCdx37D5frnj1HjF3F8et83y5K9yyC+P6DmqcKy8DiwjW9iQ==
//pragma protect end_key_block
//pragma protect digest_block
tfK8qBBcgA0M+4B/55MriwwRWo0=
//pragma protect end_digest_block
//pragma protect data_block
leWycT2aM62irUzSjBIAAg2xxhEyuUagja8paR4qcr8l/izwhEd3FlcZ5vYJdTXL
zso6F8y2GA58fSlnW/m1EPwhL3rwpxA8neI7kDtE7OQ58jZtHD09J2uEDRHcviFM
BpRqQYcBoNxAHWIWrS3A9kzugiJ3NIn0gHyMvOnKah6xCtDN3z9Oh9NySxIvHX7r
8KbUyrQBWywNack858k2IILm4NOUqoSm7GoVyet4tP7N8WEhdOXtMTr9X5LbAPSC
cumG46xQpi7AXikqRkTi4hTGbeO4+ZuXU9XxX5Bcbhoc2fjzXri5Gfaoset0Z51d
FIu69WlWahi4388y/z5jNw8+ShSTIlEfKd3sG2Bz6yNG/3d9wpBztoqwqciJ9idz
xK7q4gTuuQSSwjA7CDh0CxOaW3MBL0qkW0BZhURTrC60tymnUcdTWE2nD1buqtVp
MUfBgDtNQlrs1/iLfm5K/PDB5FDKD03KixJWrd+GPRuRnVV9+99nKUTCM0uQ3tia
nmmegcV6Y8+pVV3RPw68xLN1cMl8nIUuImlBzuaYQjlyQCMcudMm1Oj220tEm4qP
QvYrch6adn8X40LYFGz1FjRCkK0VZOPlI6D6UByQMDv55Ilh6Xuadhva1V0IAbKg
TduQnGN1se3SEtNgMORnkgYkt/YtjVRZD3p9M6RTsxuU7zG2LcOaoeoe0cwix4Cf
fy7OS5DlvDoI1yYOJjDciy7u6/AyEqLxpS79H2W29rO54XpBx8+BpvHNQWNMrtvC
F34ur4EaPwdXxgj+TGgTIkGDmGCW/591qYHGTxxfX04Avv85XJmvhwX+5vEBBuDC
KkIHzQVMEx6H6AvLttjKfI/UVhNOTxqW/zxbCAwaOQXkx14ZUEHj4C4cZWPnDggD
exw7rhITbor4hQkM4P5UllpACsaL/2SIYuU5xhjPijDPmZAbSZcOAuGqLWFOsVNK
rqHqLdhxQU1pNyqhkcvRV50kYLy1AJVbujOdSESFkDXLIIACw3BVA6+sK4vj7HuT
zkSDUjNDW1vl8fPtzDjirwBpnJswD7jQmrj8fB1g1ISt2WqZBu8tQ0bhMNG5d/Yu
82Jcxv2HSlFVVMmjQ+oZow8N7Mgw320Mf9IWX/3OuV4dS2sumlzQV+V4gSavEErt
Lc1yn3umufCTFjQIC3NkcIrTJEU99cC6uLi51HV6S9YndjtGchdPudBsYAdl9BLy
7SLAX2Qk/3U78FE5gyqoaH4demWgBWAIDoI0NeTmsBai23t5lzXa8RejP7LBvRCW
BuoTF7izYHOhVBoQhnqPInS6u586rGtILJBYCT2LilmgGshG0BesfqsasRg3yop6
eTkjyc7CC1vMiw3UXGelNpWnEbo54PtvSFtYxSrCONnNVKdP/3bAZifykSFWo8Ov
+qLHruDMvtW5Qfe5qGmf8mNxlva2QNQGSPdCsmmQo2L418IWwOUfJQ42BdOEpTka
TTNTbV/z1a3IkmHvaqjQLibeeaqiqBDShgPGBcYg+b6rgKBlo2x4qO9LRbNOzCud
HNcFv1fPOmztjvSrHeHtNRdjwGS7sBFoaycoYmR94hEpKdmeI4OIFZ0MmN4wfRBe
HCZN2Q5QbWYB5nbyq2yUGb2FbOdXIzaqMBQ7DQYFxHNL1YptAEg6fLLioCNfCfTl
0JG5FQDAzfAdWi2+ND7hZfgCcjcMU1akYaHVMvNmV2ZcXoKV7EmopMsJIGNgxVp/
WeVqzdniPPRducVGtplyxCntIpGMf32iY/9UhINDtuEvRh/O1cCzPRzOVfyzuIhP
T9seB8Tw0DgQ80yMYGdjxffSUiIIkipUwU75M7ECBci6SWU6kIzrslrxqNiSovbs
HKLEFuOhS7VFmvgivKRuLpz5mkPFQc1vWKYtY4xqDADN3lioUfHxSVxQ6QPTZkDD
upxls1fj0fkcVRYEi/T+owRref+hhPQucki+P62NZwnnonjCLs3sKJDH5PHFLuJP
xhaOcOg6KFTOan3UA7vjDjP9xj1aPBDAPCCQOvO3OdK0WyU/9CCb3St2GRj/woxz
UWvr/YMoyaApDR2EUUIQ+WMs2Fp5VthbRAyqO9HRdcsteWaApZ2hP+KYLt+YxFpC
BZFMvjzB5kYg6Qs9JbqL95GERQMCRCwD28KyDkb9cgBQBxYo6RBKaC5NRt0NV/Q0
d5mWZhsPKyhj3DGbb2XJt97znP9Syz4iXNfyU79sPBbDZ7f+oopLwZ2i+7rA8W7J
fXCnt4uQ2jaYByr/7twBIySlLfYSQNYjrjfuksXXF2UO1ZPnByDxsL7oXqzduzKE
dFfjJAg0b8ZTS39TZbnOKC/rSNtR/5LrcDAOCz5DlBmRLIdiN6aRxlEyKumIk6mm
ZNd0ALVPfsikrlRUtTbc94qxgcSimZmVBFH73r7HY1+wmlOpeKR40btOLOOzmDKm
bzd1BDwgSxXCKaJ5NFi3NHNa/0kH49vuikGbreR9qt7G4lCZPuVvzTMZQh/SYFYT
8ThBquM7BzUwywUlSpFekV6tkjUb/gET153dOmEYflvh2tRWLhGEkg8edG68euZI
ZkxdJqo3Rb/oGyUQnXsOYSJ2jyBGUUdc9zepz7U7HbgpUqAIBbeYsCpcFFRg4NuF
KqajWEhgeW0BHzNQFd7coZVVar0ztZSUxlQfTduS7ygxN3JXpRXkdevoXwstZliX
TSIA29ALLrWd7dUClsOhDDxGNQPSoZ3mCz0vTHBzA1JGK/eT72e1/RyKDQhB9u3A
3M8/0cdmkph6O6uIRObnC31zktvsXIwTARXyd9cYJp36En/YqAZ/zCFRmk40BDug
WoqbClvd6LJeGNNkR3ACsOoYjm/x/CF874wqAAswHcwLNDtiOMYUcggI9BSobsqQ
mmqXyB3Ls+58TUCYqcn0Djs4k4k/d92c1m3YFUkg5UaHFGcD8eO9Nu9DovdZlGVo
L2cviHFciQG4E3Gwy289Gac7LlP1uembyTKf0FJY7x7Jgg4af0CGO7ZIiK6Xt1jU
YdLIVsZUD0agvPI+T2oN0lnADGAYC0h/b6Msi0fFl8UzpLBR5ft58HB7HnWEw+++
aCTQsj7WJbHTP4dwPN+hIvT51DMV0N44PbzDfo8yi7FBMLy4JRnDSjkgX+9ZmokM
HtIkvgz8v+LZEBlCVIBfuqZKjOKJHuTVf+vpi9fJP3UC1txXnIj3RaV/8abA+3Rc
HW3Th8r166zNISIuqhBudjFm3kJ+aif2/OkOBkbjyrnGYL535WLamMMrukJMi1Fn
O4J8QI/fb9t5tV70pisvDN4x+VrDPS766HEGdtX/phxih6QDsOk5P6XpIAXQWTUK
v7tp+2tbmfnhXALo5X9bj1WmoI51hJpq9v5vQwHV4jcJaLvcdQNNKdrbjvO1GOQg
xIRlNvPLfkh96cC4nq9dQfQOXHFJ1nPZ3wNfkKhwEhxBesJJ9gvC3qnUMNBBqsEQ
QmA9SaTM8BeYd74e/Bt9tVZIEtCs6r0hZgxBf7oXZyXWK8tg+cWhNdEUDTO1q0xf
n4f/PDiK3VzaNtWAaChNqTal6A4qobqGrzefpw3FhBCDIdc5PpV7G8eBYl/gBgRP
K6uWvhxkQAtpCzFKYbwDrHJ/VY936G6MAPDB7MYWq5cRDFA7u2IuRMCnM4uytHO3
xBwFDK7vGj5pgfOO9n2LbGVB6OiwWV0x093tlKi0K79jTgJbWBZnGENe4SKCnBgA
DN5M0aKJ7TOyVG0c/He/ik/eUSDjeOyCMBG/Ywounoz7/CRisr1l6nRErkdIUQjp
BiAs/+qkyJo95liyFX+abmfoB8zkToiS8pOnLUByHwfqLXLhunCI+J+X6jdYnwOu
wfunoJZHP2v9PrqmbcyDDfV9wisf4exajyekqh/75HPoxzkn9Y/8zczkRbIwNF5/
kxrY3CGE93K/Kd5S0toHzhY7IyBMTI1OfY0otybNv8ek5FKrfffepzsNdVGJjo8u
+JzN5EuWLPoL1chcuVmGKF49oYu/BRMgCQT3XiyCYSfPj3gEA0oQ3gEw1pIJ1hW6
2LTeulrXiQzX47NJ9N4buXhYh8Ooqxa6tCggDZQkhDoYR98YuYMV/kY3pYhm1Qdf
1nc3Z3RcBkHpR7QeIooF4KYcLeLhw2yj89/cG7csKp0wWsfef0ovuFS+kwf8KKWD
3FhUIdneY78Gom1CxsjNBQ01E3NZ86lSkwex1lo1ZfvVvMU4ktC99EFT5Vmjhox8
T3RuK+KXdIuMdvXnVe1FUWpru4VPQMjJAlw23FBajfNhQJe4xdCm4RzcHT+Xc/fz
a1ElUObC3wz2J8MBfyXAQJgQ66up1vDdqzOQWS+62OPT6z8a32ERTaEGSclVzS8X
ULOQI0fAm9Hg12c5cGRvUxKl72icDDJPXcdsd/sjIFJIPBS6mmFAItj2QfJsMRCw
SWrtaA6la/MVMJLZp7DzQ+tSBE4FloPXUTEB7A5A7LEbNKMoaf/OMZps+ManvF2f
+saU3qT4DJvzK0e5ZbqOJ6301ssDq/wA5oeSm0baFitsK8Uojzj2BGnafYsVrPpC
jqE19IgNB7Tio//8epoFWMhFIkLnm6D2x4Wp8ctBqCyfvkj6vxEHWD4qroROObnJ
lqW1YRy5mGmT0sDJKOfRSZi42zYCz7OkE5jvAEu5GGMqjNSkASwVVIyD5QCwlTFd
H+VbsA/jjpSw3E80ZOAo+XOq3jn14OnFv1UHXFjEiwvsNjeDxrtZBtleA3Gp7HlA
qERQ4T9XDmqaUwUybyzuH/cxa17I4F4fkew9czAg+CVsgpsfrJMjcz6TKXNDN1vL
iDWt6mtErRA3zXMGUr1yHWrx1IMQeeGJvCDA77oJumicHwflAUFzUwervfsp+QsV
k4JMYrFJCPRj9NuNKtwfrMMCgacY2Qz8UF6UAaOUK4McYe7Z7G5SHNeGv3QTtGmv
t1PXvE4mcc6Epzkuj6MYGKvXM3XAAMZ+YYdSf7w+aJuZ6RMg3Bzq4/Q3d6+g0oLe
JGuphWp+T16cqaJiWq3mRG/q4OLE2Qa4EOQxH2o2jgJ4G15Cl74zUTeV/THjWcEt
UQiG1LzoIqul9yE184zbKx/0ngYN/v5j6DlNa4V0cuj7/h5zWsdmMLKn0qPonAy3
cPCelJrhJZpT8Q+qKOgAlz5y9czS5VJtoj+NReQLHiKxXpBtWyB8zb9kPBGbPsKv
RUhCCzaqc5nH0BOUPNsZS/qK6zV2hvtHJpmrtWln2j/fz+ZhHLd9pvURbkVDoN2Z
yQYUXImt6K1X4g/95pYwzqSHbA+mJBLrJUkiA1zZGrjlrVZQGrvL9QBRomT/PeGi
OMTMKYEUggzMj8HCvtbEffeuJuiyQR1p7OyXWkCaTp00p9Nw6qfNmicgB+Bo8X+U
1Ngsl7qAnAx3N9cV5bVYfZf+Uq4vA8l+9384T0K60NmEjSCS7QCDDjNqnw0Vivgg
AGar6tfxx0mQHxT3+87PByF/lTVH2f1rTVKkE85GHuO8XRJNXDOfcbBdvjjoQAl1
qllWYbD2IsOqWMXCah5cHPY4ZCxUtYjuK0QAq96Lcse3gU5BXGr8y0P6Ks3MYtou
y4Mlp+Yhh0IE55VL/134+U65Ie0F+Dg6qn9NSTygHuX7f0EPLQoklb9kYwAIPd0L
v8WwTtTGku8cspL3wtCdEyw2YhCMgcvOLi+FVIZnL6qxVzd1uvAdtwd/rjhTEQuX
iar7YL0y0ebcRq38+2172bk3oxQR/NlGvFwov1e6YiBbiCq7ptLI7y3AjFFXfafx
xIcPajYUPLiL/+mtPziiQFEKi/3GdLZJ8joTXAjl7wSTmISa4EXD2w7UmuAQ2HV0
WslPEu+p1zftE41rmiU+2iQ43aUdvHMT8WfJlSf09dgn+9KlOQC4+odlev6zdQPt
RJugdvkHJCLzTvqFjRWI69MdiNYiOhsHg11Q9cU5nmF/Dk3Tovct3FkzS6VObw5d
+JRnoFUuB5H+72OtOcs3DkZmHu8tJBq9b09Xbo4xXuOmlGrRS5Lz0dxOTsYb1rmX
WjT9coFAO+/yGTtgzPlgcyCQieMr+segmq4/NQOtwDlKrcC1MuyLc2mX5MddY0e3
2brkPBIgX5i/k7n4/Ll9AP6lFKtnUEFut0mfrwtQd6aMhSuAtjJtgqGWMbEWHuNE
sYbLeRYjb6MaMhfCvyrbP7H4mMrs2zRZBYAC95qndX2abaVhuNp3Bv/FM09A7Zgh
7U7L2OMKWxWI+bXDZU5M40Gg0uGtafC1CbQYeP9bLIliXHoMt8pkpvOgAjoA2MNb
tsPEWKIvYxEoA+i8bDHi4GwkqWuIt2e7g8SWnqrZ0lESkhESsg5IQ5c/o9pfnkWB
yc+cMlQtMpD4waEXsCA8hMQM2K9esk+kRdcwSzd353EHApME8JZecRSc6tG3oVag
FeTjRLfuAImwNKIKFd3rGwvrSOqjvREc6YGCkuz0XvyXdThma+pSobPO+5hDRwpD
QRdCD6Rc/zB/Vhc/PnRfoZIR7jNYNIaT5IYW5Ji707SLGmszt5nouIvXiXKaeeGv
uUzdKDkRd+NCRgnwuXTjorVQ7cHi3LKTvBjiP6Gc/k6PaRnbi3HzLrCStSnHKtHv
fF6g747dl9hyG0nmqm7b817E7r3QZms2vKSe9QkdshsojRAlLEC0PhVDj0CCClVc
qdTzRLWOSU5ZSlxLKBT7+KpF1cyvNcPhfi7MKZnAe7HcKPEiH1VfNqPXUZT9e8gG
9T2ng10eKotczX1cY8D4mdo8Lr7MT+WFwsaEKPaEdW9+s0mGNYGy5EqlMDkwlqjZ
HRb8hHpCJULI74WYhFsrgt4L9KKf6Oy0DiJ9X0Ohhtf35GQmbWCOeWt3fDseQbhk
oSLR40GZEzLeKLOmpTda/T3XWaI3aeg6I2+U9XTMfDxF/UIPXrdh92dLAbYGU9u5
yUvRgbsBDSFZ5XfrCzBtwybqahqP+WlQPikUQzDmXNcBqYVHjIEs0eKdCQ0yjwbU
DeVV7f7t2PKfG+OoJhLWKMHidyxOkuSD7BQNvkhi8Y40g0A4oEL037N7hZ4IR68w
sYX7MWUtb9iAfUlvvd22sLrGy3BVtJH5qi6WOnvPCMNv+lQ18Ilc4/Lc7SRJtf73
qDcmmlWiRCQ3N3l7pKVOd7GjsffNoteWbrM5CEnmHLiXC4iBzsZoA882C7ZjP3KR
q8+LCYavY7+CY+eZUPxH4vv9ZtZihdN9NLHAhnjWaj1tyVyiWH9UIiszWvr7sXpk
RbeAHmbow8Y2jm9K6X0E3gsOwqOolQ/Zje7mHxVq0ip6HWnOWaO7MeBnmVpaodp6
6cm7x/ukSuydfPVaMHT3kxvFSAqfarnDw4f2o2Tic9jh5hfM4zKUawsWLQ8s2lLl
SK4VU54o7nDsYY5fPP2EGX181qJJFCKZKkjInbDpCDzUcBM0ihspDwAhhHRkXyNJ
p8KMP5hk976976FV6kXt4CU1wME1s9v+amrxRTyluOGgUSynr2N0kC0b9iRwN75o
23kTu02K2FlEKMnKZMjTYh0UTk6+5t1bWQfZL3nX8ikVePND86iYHLTo5YA1ngpi
pJKwFHdqJHWsrQVMjFlIzGOZ16gRrUmNCTbi52yR6NS6JqpGZBheSF9ft7E/xPLg
5M2DHwfAsMKVGRhAhwaM4QGpn2MWm94Mw0dVLAvxh5lOmD4CSMWsL7i/VnkFz9fI
SMTAlhlLPdwzK5ZDlAlctoneHRteALIwMQtpxr44DEFvZmRcG8AQEQqoVVvmttEJ
XuImEfEOON+NAyvUJGJFE7ux0ZQIiHwKQ3pRkHsTc0e/1mz2dJRQcc5WgBESjRaD
7DNjuijJBtF0/HTkgw9o7AxZeQLngHquFBF6lTTqfgiQ2NXeWxwzaKmgSbCOs/Ev
MFzx0xV29jWd0IGYQPwd8kr5PW8iI72An0haa3dzoCETQNq8kZLvj19cDycf/WMM
V4VzMCE4YRvjYiBDmaxLPwE3qeI59arFjvhI06pNMLCGuZgVv4M5Xr0Baemih7/M
Fknaqg3JsvbkXdXyaWAqe/m+vFwsP+DlDV3EGt/Zc393v4qZFVSuVGz3dvZ8UbhN
Mo8zJ0b1buJzMPT8xkYM5Y50QCZylNN1LsAQgyRq4sDX8tbOFBUeocFoyQnRX2pp
/1XguTowoHMA3pRtJF8LqVWLGXjKLYEvE/N+O7ZzjoWIpmoBeASYf957KqalyKCa
he7asL4X0rnvwtWreqmOXDNC0tl/7UZDF56guRHR2flP9NETD0OjUeMyVB17V8Z1
fa4tx5rQjevN8NxqCs0WmZ4L27EsatGzKPVQ64RdZHKN+7OgkNHm/O7cS27bEs6V
8H7pbzqFKmsqBx4NVFs9rcqK1aZ1wMLbrMK+pAVRCdlIGeAAiMh5Zu5fwxTVWUnb
Hyp8gtfIGJXAAuahzhO0VReFJtZY8N1BEhMQR/LkT8Tb5Wb8EJCzEPsCrauFEwYN
IOO/gaEo24385B902YgjSkLjO+mDNG8e4T4MgktoRh4n1rVpaUd1u//PlzgvlCs+
SuiD7enWIunSE4LdC+mhDH8Pmy20urQZIO8H18iFKj+g9SvbTtx++AMbnMqoRl83
BbErVV2KzVUBQsTFc6y1X1kRdMjMWxXF2eS53WdHEneBpJs89+laV0dJrNBQS9h/
90p740CM+X9kpvdw2ssPIETlCYNiGym9J9JAMLY3WbL/VgkRHHlqDthUwxYUveHC
8RZOvzLH1cGiWO48D7cuDn6L58/GecpXvZq8s6IHdj27Shy0VGJPek5GlKxSKchW
JMNM5INucq5jqQhx1pMfD95HyoSlxDjEwlHb/rx3UqXR6dJoZT8EuQbE+M+F/zjI
0Q02dFcHP1lMrwr/jZuPKHW3vFl7D+P61+n2jENv9fU4XAZxBKYfI7pTpV0w4Rd4
SlbDXOx3Y7CHl6zzAfYT9mv1lhHThsK553hevV0zwKvFXL9Yeg0WQ6ku1DFkIoM0
otvywY2v+uFbjYosHPiweKTO9Vyxnq7+p7WO+5Yec9NBwJA57XYOTQjh615smRQp
SG6DQk4MdUJNxu7DUfEM4K6TIoikOBlr6t7Zww2+CJ1GSaqi0aMlxnj/wOtCjSiC
HAXPcRGPSqJOQN6avf2RLs51+ryCgjllvWwiiG69bC3ITh75S3TNV/fCCGWk4g6k
0eJ77Fof62quJo6uOZ1AjBpmLWVJXLNDjb3JrXbkMy7gBHeGBy3RbIeh1ZAYZA+h
ig2REzOwa6gppq4jBfhtVBWKN6b2Gq8hgk57bKmjl3Nkh1Z7sDPvSWg/OTIN2hGy
pDz1qnHYU2CyAkDG2xAym1BWAuNAJu2h9zLKX/AF/w+r4rhaPPTLqAqKtnUy9/dG
wWo/NAJcAnnjRIH6dLvDduQFZ+P92LYUDeA92AwBykvEAB/WpyscdYnWsWmUXOTG
HFRWq4gs2eV/BNdDRUZTnHPEwHrrok3MF4OsT2esMswNXhSn8kDlniEYyVfuQOrc
iiLImPRVqPPbQWmiisVS0shQUS+zqiiZBsqzpjBzMKg1o3eUGRh0n/KfZcIPfpoL
lQUh7ySDKHujyRG+imzDqHe3NEy3wa610kVzAxHzKLMr6sVL1W1Y6GQ+WWJa+FGY
WT/6GzBpI1d+sVxVNbw/oIM1krGOI+q4UX3Koj3xkKx11stDUvLQ+uKECfWuoSsE
FxpGifrFA4I0TTPmEj1h31mDRg7RIpYc1eo8IdVsN8crgv5FckAfv2Bp+0lPVUNy
rbbVFepR6jPXtEZ3oDDOAW6jObuN67i1BiYR8WABDq5CpKoLzSJ17vkkKfjURzmS
NSdXJabuJ7blWv61n3ul7RiyYF3UVI2v24d7MviWHboRa6ogbG7XE4dkqfoNX3P1
JJlsQCEJUSD3a3QJYTK19qXVmXPvqYf2QCQj7k9sBVpluL+7msv0LFGXVtySG3Xo
oPgzXD5jQR5U8ka9b53nbVVB3440mlPkht7x3JNV2hKMHCg8mIYXXIY7GBCzVvSU
hy/Ew+mWFXp5Q9mQYqHm9XGX9SNKkGt5pPuBSxbBnMqkRr/5W/8Z4bWLcAG/nTgg
ij1uqRKEEAnK9YLo3pmlRqp1pcOAGI0Qpn22cFAgiz3KAhhc6hLPqEKZ88884gLk
PnzOFholNqFfQAaZvG/bVmGxR46wMApzTyXSE4Aj3pceC1oW51DIuvj6uobpekHz
haEhL4rrCZbkWgn4cPCqhfwuIdgt114FL7EPl1KStEWTpFEZdQPG3EXZsK4Lh08l
IzXZ0iiIJz5DW1CfuDDLFt0KLUTGrw/RJhWBvvZpSGjmY+wNYfI6+crHGrBxYb7O
O67jmJPErdNIt4CAdqpfSAZXYTxslTvZUzYHyQzsNDzgAmZJFoit2ei1Wj5Vs8To
ISyn3kF5zrREgc/lZqJl/A0hryzWVniaN0KR5XW1UtzWAVIkls4IJ2KliE2LHSuf
TLTK1bIXQMuBMsI1LUHInvtjf4BL3AINRZK8KcMMFgOofpFSfRxsMuXHmiI2rATc
aRzpdZswGa+P1pG4JskyFFh7jzLAjFPklAeHwZa1Ln+LYoGYogEb3+eC5MkueKFs
6XUQ8vMENEhmls8D7QQN8xiISUwNdOjfABAswMO0DpzVsIuHCCUZlxIkhU7ZI7kx
mRFQhuJmr688K7e88x6M0+03zapYeqzN+ceZJZaVtgdVfQ2C1fgFckII/XeUQDG/
jFOdoDV8AIiwWjU/2q0WR36tfe8v9UBdphdMLPkfSDq1FJyzEypA9m/3ByfIjl1m
jlXKnDWWdBo46tchoVBbFVOwScheB1cA0Sl6v/K376SN785c6ZoUi78JDBY3vN9q
z7+N7Ap2ABWXZsjUodfeQBBTC3NZokIkxa+w76zhHWM7DCaBeJNIreL9rHDG0RT6
XZJwzFabWqeVtOMkFYvsn/skupsiKmdh2xFMGQrTAN2bI8NH7YijIAqR3B6xGcV2
HMw2GZhZCVoyoUhxpR1OjQGQoBJvREISoImr4tDnWgoEc7xZ+DJlUXTXbUB6Uouz
9/bjmCunCrWt2vMB7X8tdwRIBiY7pGVyJrkvv37UKjeTPFEHBYxUsBQkcxHB+Elo
AV0qYSNm1ufoOi3lVNwdVBJ+kKGIdm1Yt5K7+qYhEbT7KgCFYENeq7rFls4jpxKs
L1OxnVPtmRRqmZVmu+kUm4A9PFYry0P/4yoOAAJnSha6Dggr8JmC0hFORshr1xE8
TNVcl6jUt6Wh+N9mNJLLD7hB28K/SnG6iC8LZBqEmwpV2R1L+U6brTnXDjBTdYEf
FlrP2T4L1FVY82I2ldMFmMg8StHLRaqu0cNvG+LA0FmkG9/zRfjzFTXmTBzUxgaR
9zK8WF44RJTNE4mPCM5Y4zRgfzlkXgFqNjL5NWv/+tYEpvrr0h4JL9wt2oy3dgu0
JuVUsTkI91Uur6cmwBQlvIc3rt500WGS3y2Z5Mc9ntp7RvDctmwi9FTdkAkRg8QZ
P4CzjyH8qIM0K9dfSE7xbnRKz7yXRoMOGoMCa1TIXnNzuGeQ1oBGtxAU6zJgXaS1
qWU1Co69LzpJuvJE7dgY9WgIkzg5nEKr2EuolQIhPgjeMGzlxlnY/rShTM9QtQp/
nftcss2fTJgMBh6ej1uglgzyGUXGv0PWiaxykJXDQZLsqCeQQPhvzQnpc0QWJpgz
sBwlFf8OmhnUDaQcaRyklm/YrbbjRPxyvzYa91BXXKsJ+4N9ATzGqm8QP2qv/1WD
JcU96UKASCy0XHyfBbEdfdLvdJdYrXj2N9ssSkrXNFtGVFer2GkGxQwZEJsaqpU9
6geFtQFTpkQEE053VQpTnBHtr4jH3D3VECBWuT/mRzjQDD2tzyJ+8bgmYpRxeepV
texU7lmon5T7+S+PxMuX6NmRP2nGKmk5UNwnOZegGI+1AYo7Xu8AhavNq5z8OHMw
ELtOLj+6kQ9HedRAw9nAiSD+GrMBP0pOiwP8dFRcwrFcjGUd8d/kKfbMEzh8ngWq
KjjAt2IFIs+tqO/ndqYzZbyAEMq7H6d2GDoS+Nnv4NtctvEzZcLTl+sP2bcApGM7
iRPuStEseBOjvGHyuiGoxzOD2OFHLqptRHAcvonlUZ0vHKYns3VLIgJC96eE2w0Z
swkcYLXPYk0Q9vOsR5q2xEaF49llMWPbaB3KB62vRJ0kMmnAvmM6U4kYOJOjcpVY
WggJ68BtvDKi1Ae3Y7d2Dse61z8T8ImqGwm/9ZgU+7opy8BP1vNg3L1Lw5bFUtOc
Bwf3P2aK9uk3ktdAi0IXJbocs09k2wxF6UQZnKp4r2Sy4KqhydddpI84zHRyQN2m
UKiBgq8epPGqeL1rN3cm9y6nfW722SQtbJ3YWffWgm1ga2qiEd6LU20NI46NmiA0
cBTyf5bJula9JIwCUL27W0S2BErOp6LBFe4D6ym/yHX8Jhw7waokdIFz2kfTbGH1
bdwjCMRg48gCCIzi1EjbtkIewtLttaRLTZhV/tK1AHU019jrLDCg1SMMyDM31rkA
9y9Bi1OaPVkiAblLaC1gI6GfE9dI6dWGuGASGMlgajy+lg0ZfqToxhgueNzxtZUn
VSqvBNcr54VRBI92tB8ezdwIfBEBzP6mqoXvklsslS9hsKwl6fNjxTFUzIL5bgyR
AZSKkrAVt3izKz+zTxAIjIzocZsWVk7VEIN3YKqzEv7KEhEXdXTeprC5ORb7hXHc
oBz32GLED+yyxviRZI42zhzs4t+jpt+7S4hhiGBhbT/oD5DttZoospkL2/jvW3pJ
rXXaaEk6c2FxGietQoRUbwbdvmzTtfgMiRANkW6kN3JCsNoxeFtVv0GfADCwJLCX
AYdZU8uidKXN0nGsiOomb1m/GhNGipjf9H4/s+AjLcBAkLQUlh/jasQ9YkOto6EQ
afmzu0ayt4bXSD6Hkb0avh4jZfpEwXzwldi04F5D55DR4fNdf1gHxqVbjExZ4hqQ
wPbuViTWSDJ/IZWeaIBMSmvWMLJyfDtZOKQij3vhHDO/K2uxZ/F1FbGgMoVImcv2
iNhHVYq1nlnvvU3SnjYQ8dFkLcWRdw5XEfQogO0PWpXzSKd0L5ePV4ncAkpub9Bu
7/AOs5ruDH0IYeEEiSldTIpJ9tp63eJYCp21oHO8XNFCmCJb3sPQ1sOY5Tyx+uJs
YF34Kk5h/cEuHoglIUeeXIsDvcRnYVGQM1/sDk75WcvwHyNXKbI8/PjaZvILQHMx
Xy4gU9f8ov430rcOsQNOTBg9BS8kGLbIXvBJQOLVJFZnrEJpqqpg5vn2k1LiCH7e
Ik9zUCGOi3a+9ZqW6h6eDy6LJ9PpxkI0JjCMjhtBj+bOwDVVQxXbKZJONJIvP1+x
NYidrTqrsMXroUZuhOrGT++cRjs/9SzDCqmhVdEJbHw/trNu+1FkiIRk69t0ih+U
0qHVrvDSc/Imw6R8dGIYF95IQhUu1Iv739cw3haO0/fFyYAA+ea7b6gQO/I/VTg4
UXPAenqx7ODtboX9Op6ztPEvhWfdZobflIoc81gfqHJL4P2SyVkLz26gjv0dzTLY
Gd0tAbm5e/cMVmBo14RFJzZLSfMnolE/wwagXzc/Qm/lZOqd8E9ilVyeu3vJ9MFc
YCIfQ+yvvZ8g/CNix82obqiiYsrtMRD2gXS2cEUVICuPA/byPc2M0ozVZEQ0Q/Zk
Zgp4PxBsM+6cKgDa045df3Xrj7pStoKb5V1r9lF0YGJ+itLJDM63/60Fwz+f1B52
ir1rAXLYrB8ZNTa1xICCVVNUcdxNV/nuMu3zBte8cvjHZBVSfWLcmQpGuBCdbMBL
BVoS1Tzu6Jm0jEMPA3mAhP/PC81QVSUNsiYEAh3L0Zme16Tl/1PSxQ0euxYuBZGv
EcmXz9dYhAvMX0M4vYaTUykEhR+SHEVXVD47vIqcG/UYn2c+SQAxxR5ckBbXxZhP
gZZjzE1unAdB2fBfwGJnDpJd4j+HyQS2+BC+XRZKyJvoNoKNyW204Sqhv741bhwL
RNQNPAq8vqlUnktp2tBFD60h5w0FFSi20QQDhUZbOjNtQ3o+4LpztU04gpBxqTxl
En3w2klLLoHsOV8Y3gYDdicP4fRXkXVfhh5pw6O6kbDBA1Z7ZLRGbEGnqbFhlNH4
uAdHDE0H+7A+2kh99SEdJ1OGnMHL7YUEbfQ2wIevj+zePxmq2w4K7xwUJRjuRmOr
eeehAa5LB1W8+USKo7Gp2Go5PTrzz5Pr3plk23omdc7RATtjGrkLGSZTzY/eorFl
Pw90tm/V88B4y5OwltbQmvIhCUoth+K0aBAecpbaqm2MMa5abSV0dpdUVcPE5se2
t/dRAh9P2r1y3B2cptwJF6SOmgomoC3hYNsu1rcRq9uhW2U9vbzelJxBKdXRWgic
g8LQIwy6KMB55jzsbJtwj1cmhOGr+rFw6AgWUUgbptFfmHR1nE12ADXdrZ2Lwc0n
5eZ4vaw/Xdr0HOYWWnbBovydG/TkigVtgzpei2yd3NZn1nWqeqPLuUWelsGf9DxH
HWxfOEmyeuhN0iKWCxQDA0WCxXJWJD8w6FDx4/9vEYH+DqmIfdmuv5qt5pfZu7cw
J5K1JKNp1Pt4JHiG9C4Bbgro2ffTQEQkUqj4aJx5UKSO955++SqxNU78A2nrZyzD
96Pcjm9mrmx16Dcnii6LK58p/Ba2OF3PPLDF8vAC1Rj0+0OlFhA/rYk3z4KXXV73
Dv89wEPYFwisSvWuw5cJ0YDuFgOV/oWGHVT1yYVBr1jry9ubOYu91x+1pYoMP1W+
Lj8l+h/YtYHe66BUwwV4cp1mt9QlgRBr1Lc2Q5YabE9qQYrBPi+IPeqaRCBggckr
TMfAcrSAphlOIgi9oNHzvyDptMTIsPHodOr67uKl7/1JmfmvPAszOL6tKqLeJ4dX
S5t3q44Jw6WM/dqRg1nrwnfiafZtvuq4rZYkVOKRN7uuVMf++8IyOq/XpeWaw/ro
qh7ztsAGjkbmWaGtkvnOwjrMtUV6ixj8j24tnhEWlaqv+Emyjsce85qLpVGAJOF+
hknvTOiJFecEpXLFPY6jqECOwH8wFvtDD852LDLM4C9TM2FjC1KY/uHi4/eN15A5
WfyawFjCZwFNRZxbEOkZcKB8nIn616k+nSaoDsAE22IewE6PbhzMRWRPOTIBdjxZ
6pywb9jaq1FBlpwfBqS4hKUo331Ni6PNIF4kPlAS01eM/l73JOWfWWzitFaqBQwP
je+eWZTsibCfO29H2YmeDHNs3cqzERLQj8qyNcImUW/hceHiYg+GWVzhlUyiSGFy
im189vqQr/9DCiKdUEd7fl2K6f/FddC70YW3HfRmVegHePMXzMwZZt4w4QYVhoee
DGBKStnYsfOvPmvhQKWEfFnytN0hnzNeQitv18CvYK45/f8xCkDxm79yS7sRW8gK
+7nwF+aYoBxCL3cUNrk3laAPanjkhVwOHY1BigcqmRFpOBcLroawjlHYn3OU7t4K
VCpzVD5kSK5YZ/n8n7SjMfHVpupT+Vf2xZdDZid5xA9T7aw+0wu6p9YcQxQWycO7
7CFH5hj9VhAFNFdvm3KfFBHnqgAc17NH2Y93GdGofnoh8yFWeB9a0KgssY8KZrRi
rcFQHrmxQRw719ace6yOvg/B01MyBrwMj15dt3oOoW86KnOk9Cv1d6NgpfUW65RL
9V/6thX+G7v2+X0Fvg5qRw6yCAbGraFbuWPAQCHT5Z0hEAjUsGRW5TqKe2f8R5y3
ju/1/nnjY6jMq4zbkS6V7WdZn7IEbEoBSicztx+exM0ed7a4NVbNjbjmq4syPn4s
VJe/UCzPbDtosWYsTvVYlN3NYuzzII/M7EDctVYX//5rjqBQOfLxqq0ukUc2H5/N
RvB0SfEaHYpT+HOAW9DjSF/WNs/0luH+k5UNzUmMnmKQqEvpox1/uvnmhRt4lMdF
Zh08SkSxZVaByE/SOvrwNBPMo2Q5BYTxa2sfP/1bI3VkVEmCcMDSacUj3YQV/75B
alhYgqYGUGXd0tjDgrbiODkd/YghUafjvoQ8y9Cry0K9UEv4zhSc29WT1EnUdUEd
34vM/ersCm8/ZBTPBIa/iWN2joiW7k0iIeup/rIhSa5VuwMjZfOo1B9qd6Aq2vyN
d4aOn3PiehGyx+xyuXloX1DZyzc4RiJIl5GT4OFdTJrBoiNPujCzfEawz0sG2b2L
pQey65rXEBjcpV+L26pVCViCiIIagfFlOtwyS5wNoMZQgjIhiyQzUGmfBIN0XFiH
tu9QnWK8D6D36fp5nOlCGQk0keJKIWM05J5CGqb5qkzp4OqPzDG5z3X2u7jXBp+8
Df9QmP8KHI7fp3xnuDHvTnCr8jowNKHRWwR9v5wYy0DbDnCZzYSWUrb9HPRs9IlM
WOcnbpVATbaJCcWphFoOc8wrvqmMBZN1ESp7rDiJNDl3VjARknUllgBWMklB7JSj
CCAyBlGekn2fdMNki925FORXLGB6UyaT+Nk56A6IVh2aRgn8OiZ1cyP2OwcVlQbr
qcuUp1orTbjrdQBhfiJwSi+S/NQHnCPguPFAD/RO5G8cpapPKYe1bo9TmWayR+dk
gXBdzCa73YTw/EcMHjEDnX7CWnVlSMjgDJUHAMyVfroQy+cJiHBkch/qJVLTnX0h
96PUKtn/OPl0ovpataEV+cZ2bITni6lCBnairR0Mnhzb136jbNiR8AqYCcVsLE0x
6ysH0ibEuAueUFlE4XUV3qkvww0ZsaT6CR1r48qkPv0ZK9PDuZz6NOZkazfHbBNy
dSLtTS3YrgxQf9zeA/HTnBj6Zbd1fGp81IDzWrD5kVc3sQTDxDNpeLbfrEfio6uR
L0wrAe59IrB55KSYmAwQZbjK8lbgsnylxuW3UaSMxvWOIo+np09JVOUnx47fI3F1
odn+NdAkvL6CgLIPUAMMmGSTBmyy+gnjwpcT65S/BhIS/Zfd5oGQnN3mvv4V8dNp
MeK9VAmRyXWTyRicx3qD+Qu/2ahZIPW8085KL+J1R/t6jLz33ssw9jd8TxCISOQJ
BIiq/u0J2zN9SQiZryWGcVlE919nRSUn0dFHO3a3qJG/D/i+Q1SqnVOWvo79lb1r
9ymMWdyOomYygslhTDBhpdXlS+QF4EgS00kn4igLRP+G+jV0R175sT9FqzqGVVnQ
+LFOqhl31s0xfVnsK/h1bBfZm9CZ2KfpsnR2H4k4R3sizkr0Z9nOc7lWAdZiE6i6
NXj2/mPZm/CMNonjhP+aetMbTcLepodUqajc5cVMqW7wcEkKx56U64JZU78fJBvl
EOywRze1aBQ7tvu84lURORQeXsd585M/SvTDksHUGWptiUlqXOHfNjVJ8uXcWJCK
kjdxPa+v7V/f1bnzvFbqL/PDhSDb7Rdft0LekqM//Bmh5D5/i9o/VbW0z//xt2lk
q+qndnkdpvmNswhNvPmoCu7sA9Nn/tK2n47KNZCiwvLB3+e8P4A5Zi3Y4cwqEYXy
ThnFdTnlbfqGoMwqKf+EyQ6m8mUYX3goPHdwTX4lVOc4AQh9qLg1ovDyYITCTYtU
XmnVrUJzBe6XmgdpSMRTUISzzXo6uoi2866uF9Rz29Is5XIozauMM2TkGdlCyVMw
6+K90ClAkTF8cug8itiTOVj127oFQhmIOPfnoth9NQ8klk43Yumf8dXek2c7vtXe
3zwFmZaxpTxfvY0SBYl3FgLC+7jL2EXr99IM8P5tdxCG66kkGV2ACQ3XY0jqERL4
mJHPOizyJydDc62gmdmNAa/FkL/Uq5j4rU6NHZ96lCE07bCyCBExwqF95Hj1HG41
llcZosoSHhD/Y3FCY7YZ/JERI8IY95I5nNw8kb2IUTCN4V6wDsQ8kRmNc2QhB43p
h2Z498qffncd0fWa4XJEg7k4rZgh4zS6DErcKyrSwh86XWqI1b4ZemyG6NQbDWpq
isGV/xWimiXsKUE/vjwkuVZx9yRHSpSrNzWCuR3Wbxx8MXQYyNCrGMEODf6Vyz7p
LqBF8kvSq5JJ81XjGxu3uiX9PH/e8Ovbfup1VAFV0SuJNASMR4bxadqSSyFnFfDb
FQuGVZ5/jdmw5fhrzPwy1HusbTnCS3t5Gy5INPC3lVICHQl7ROdMBSLr9glaXb1p
zhiQQ8mzJf6zXHJHZOWqXD4MHSxX6PnpeeiehdIz4KQRuufAYYHGIVnk2h9xRsXE
v6jWKSGQDSUO7ZjqrDm7zMzNsPJhTJQc0rjsa1XOwPVuoFTJiNComYj5tL8Pdpe4
RNXn8woXbSuxg6aaDfy9tXJ9HDU+hwj2OHhyyrqP5Ai6WjP3XgOGFDcWRKR86sLT
pQFwtOb3FTW2DRZpj+gH3TNew1bNPc7Z3s9uc4/nyZai1XWH7NJm4/EdEasxEClz
+85kbGiJqNFOUZNE+/rs2j+fj5y7WarVON96qEUrVpigjkvSwcbiiRz2363r/KhN
qFH2sdEIYDU1W9eLPjOnL/UDBuBkHGG1U25RFh7kqMWJbpOx3vbtpJrw+XYSndBQ
3zrktIzMXPgxg760/0qoihmGPxloBYXjh2NYbAQloFDFjD2uHt6TlxadnqutIJ9t
/plW90x3BVEO59hXQQm1I6mHjG/UQwPijlbORNG7r5iZwpPPqOSlPAit7tA421AT
/aYj0HP1pNrv25aSOxXhZ3RE7dsP79yTbEKxGChytaIruDiqT3RxIT9dXqsyfbPA
zj2i+zywoKTV+0jt0vRRfNAa0xDztDI8zKh+MMqDkSaf5MgN0R0EAL5CEmxOa4/v
rftJIwfUwnx3T3xg9w5fqS/cabhshhw1A4OuT28YQkZcXUz5+MvFeo4I1YZORt0D
DrzAs8jTtJ5wVJM3TB4dYvFYLqWB6YezJTJaJMQsQkhSp5FE3n57DfQd3/D1WQd0
yH/9UirI5fa1nw5/lXWjWhW48DwJjNS7kcMdtm+ak6yH+bLqhrLl8joaVAXL25Vh
MQabfMPD4bCQ11L66rnjOwo7FW+uudawvTeGeYH40f7/xU04lyQz7DgbEeQKhNoF
ALRse/4rv5qLrt0yziBzpmGqURgi7xKnoMNg6VknmnlRyDpBgXRpZntrBoWa/sk8
eaLAJY9te8JX2qpH6c0sfPvAOW1SOL+62NPiPfaTaHGEpaBbhw4GVCdhjhxx55Xc
YtgnXdCg0HwPzQq5f/6J/D/w4KZd4EyUfd607nzS6xG9DuxwEXaRynfl6C/4MkHU
SuBmk0TIfSDg4CVUfUZzYLxwMJ0igEQRReRsQdUplt/wAC5DB5fB8pzb/qT53e9V
0YbqMCC/m+CjR71FpE0kDEZ4NK/v+1o6nujQP3HdvQVOkZ9KmUD1b6cfuLk2EAWd
PTa5cQkNqaSecPQo6FfuExYywilX9YF9msufC+3yAeSQ+qkG2D/l5rijepeRHns1
+oF1zWFM2CmGm1b2XemtGpDPrhN4j1lcncZnLtEqIKLwxF/y+iJcBJgAl2a7L31I
NJ+SDzRSYt6Pu89K8Yh03lQm3AMzvNpVrMCZP+dkibS1Hi+Ul1bTwTPYjn1V1bJ4
FqSdSQ6HZ1pbWobJPjI6s2pHidhO93GAf9Af9HxC1jOEoc4MKqcOgEXMGYzHO79G
JRwmUd3r/tG6OaM7fFkjAsapFSmqB+ljLKAxWncZcWDzQf8Sn1ZqOlpWmrZlyW7J
eRzvEPZ2KWJ31m0rqBfCh0EtFk/9rslQIg87l4dIqDPYnF5aazPMZofOtV+0PquR
of9wRfMzUt2TMOMZ4qWOddfQquIby0XJdLYxgkwRIlNiJEXlTaKPS2ESQzqIRUDP
JN/C+FztZGR7VNbSiCkk6C0DsAge9zB0bQ9oNW2s8j2vBAQAbclRJxj/UPoiUwaP
RbikhAmnLbMkJBPp1Lu88uhIXUd7LainJybDX4S7P0ey5pgPLpvhHGSJtu5vTkBh
pvNvtb5a7Sso9++dt6Sgjf9XlbPqWRtKwveP23aeCn1vjJTLZJqfsxfI8O8LJ3R5
V3zI10wa51PWkrspQIEdavmDSQNP6qIgiPzWD70e+s6bEy6kEqqV231KeJmeP7Nu
aOqODcHrEwGk59WGMRorjHLEuXarYNUWUuSkOGPM0JUpjHfZaxrDZGxRzOgpcUPA
2EdzSuQT3dM7LKzQFQYUOvJvS0ytk4zALrvcaTgbMexR4EIR1yR7Q36yjx9AgZb+
ltEtNCH/0+G6QMgpFNaT9QLa8fszMe12rYHarQWdZMV+t14FZDUSNwdbHRSEgZmB
sVQRfKdpvb9bEdOmB/aTbbYHqtezvHLjJQ9JLifIxGT1XrKPusMj1ypidLXtjcas
J2+21PnmDU9V8Kk+fFR2YQpIk9qfIysip5u4NymoZxvBgk5FkNNGjV5pSouKOfM5
7oCkiDh5HBUiGDxumGCfMsy9Uqfsh94hNwuqVl42CBFnGnspNixTFnqxJXlGWSaU
dupVHuP6VKOSzjvajg/Zi5/LKspiXaIHQye/mkwWGsRtvlKce2n3wY8PVR6MV3rl
VoChVk++LGI+n+C8R6EKyS+jZq/EaHrU6FhrKXT1pqjTSx311Bm5tWzNxjgafnxi
Cx7D1a2LpBrmHdxB9BlLbfyZozAqL8oMVm8e+MD78+6A0OVer7GSeet6PPG1+qdU
zKoxT0g5olpgccD6NSDRnPXmCVw8ddSDIwGtsZALZ8vhGgtD/2YpZF9iF75ZhADt
IzFX32Ms7WCoUT2nfuceWB8TgfLAzjXltMgedmyngv6S81O/VydTHrwObVyn9NKF
oe5wKrdQwdwyjXC+mW3T0mYVUqmESJf9rVyyNP6QTAAVBe9R5UYDGchQHc4MEIF0
nX7KN/RaGNRrgAOHP9+eDFLCKGIPxw34DLA0QmBqHPLiFokmAwTxo1I25yl1CRd1
NKB+gRO5g5mAf5w+KNJFcloB4wexMIGkLtlGJ/gHmGcTFxv4TQ3mgchspXmztH7U
tXH6Z08DvHoAfjaEpg/f4Tr4a0OJ8anQBr4pzCLVJ4WqBKPjGmGKr8avuFVadSMb
NQOD0wWw35Bay2JU2XMn3NXtN50NQrdXfl5Esq15+j/9l7OX2eQp0W7aTXjhYcLz
w+qL9dX70lp9kD764OWkdXCI7oKTlAOMnSg0xsVAVNPQbLlYht5LRDMNI8cuua7c
s3Fcufn0x/Ukp2sUj8AD7nxl09nqWsefDVRX47Kow3pTA0US+PaFgUwI5AD0qETn
/1qJfxV2fWoYSAB8E1kaIEcoQoCkvyjP0WdSkrxV+Azfwe1WKm8+jGHkspRKZakq
FV3R/PcmmNOcqgwqXWKFqCSLWj2Pbi/AWrRbU3akczdKjjrD4ikojZOVZYkDN5u1
tzdnYXlEaw1AJnLBOGqSvJ7LeeiNX6ic5ht2ysKP2uduZvZIRMIgsO9VPRMURbgw
/3uWy6TWaQuhB5scoqA2ds9aWbg715NO9MaO7x0LFshHfspYWeSENWNXYPB8eHlS
1c5PkIU529DiunUFlyiZaiv8KFz5q2SY3D1KAhfvKK1ra0OAyyXm6tnifGHte5la
Unw/mOBZGQpmTocVNPJdBXxxti9JCioqXo6eJ3ZSRNZazepQgfH+y2MpZo9zRx3G
O7X7q2YOs3DBX5cHr8kHtVyJ4zXYO5/k0ODR58QzOGf/zUzbOVqpWXaHh3f2xmb3
eCq189XHIxivk0JQg2tpTxcAgBIpVHnXhIdk+pxIidDi6xi0xTWIi/+d/rlBSpVI
y4R3rTpC2ZX23UI9J6VP8cj8DHy0IwaFEah9SpyTgWisgpbIjuqPxxU1ZUYcqbUj
bU+2Tp3o/AhjPk8QBGNzEwTSLrPAdNLPOycnJ2VVK/n9kaAdj5YpPMz4NwSe21AT
9Mn2WJWG6SsFkRHfOjO7Q4Mxkcd671l/SYIJibpCsbGH8443gtxa44DkdYrmS9Na
g8o+sl5/BWVhcvWh/nI74gsi545SkuOPThqpsqXo1jksZttcQB8ScOq39z0E7daJ
bSbSZnS1P8SElAYQ7DuNGMti8rdHrIVGIJ+LHdbWRwPDmVV2qBBB4ucDRoi+JFHp
F6mve/T1SbI6Girtz6ovx5g1nEBNMtraD/WStYznLq8dRoZYq/GTmPG8ISB6IYGV
AmTd1fbqL6v+l0hCaILmrJryM64oKgyUkg9xkyZZpS6Mkbu8f//9wKs28tBWytu0
JhbGjJyGenPrbk7zyV5Rc2TYUHqRmhGdmEuO9gkzgnWS6masHrBawXVb9tu9EpRu
wz/OA1tyCsHYO1+Gkmv9zB/YJEvAZA7lIBqm8LEgvuMqpyrHPznsy7vbQxeaouum
x6zDXxFlj1HHNaaoVhe3GtVnPWXT0lU0rig1v7HFAJBpyCyhugW1asoWU5AM9AIi
ilHPTGWgo/3widxpoHECqRiO1ZQvOTX+EUU/SAhaNQXMoM6fCjhPCRvzOtqQ13tT
IyCV8vvdUAyxqK0gt4RTVJ4w0pJqo7X/VTq33TEEgXWloyjfXotEdiytCZNvxzHd
KRUS8dWNvz0ecbYVMa5/THsQeovfom5ZHGEeK6peAPatAgX2GA08rk212Gutsjsd
kJE+fXJ72wc2E/+w7Hyi6GDMVicpyOCRTCMGPlbWeNJ/wzY5CHGz6Pv6F22Xf8bb
1xP73IRzFPb+3Ry5upqOiZvE8nZoZBhXuVhIgAhJGGFReCGYn5G3TEWfm9rtvqux
BEf6qElANffNhLhym0dF/GnjAuWhzXrmMDo4e1/wJ70QxxTVwKmxVpQDz17L5SEN
0QjxwQNZ6hZNBLM0s5qV8c443fRMc6BZd1DTeyEd9yb5ND0LJc0nNnCkdN1Tfr+O
btLKcuKZUIoTUM6cD2wdAuF8TakYdLK+yhfhwsqBVdBL4JeHYcE02TGn9hiwtEPH
2ly0JDKluW+lWhRqSRIUYlAYnMchY7sX6YYzh9+p4Z7GzuWZ8cx/NIPu8w75q/gM
5Um893T/KM1kUX6XwWzZ2Kzr9X1ngKyLrCuioHDsyZKV37CQqZ3BZcVHshrmXY7u
STk47NVYEYIgVS9qkpTxvh9pjPVsEfOcextbdNmTu3126ScgL7GRZA3L/Vu8Yb/x
roO+c2WeMmcM4cjrmVnWhypC1+7nQsRw6GEQ4fiA88KjCPI5EIrRXJzoz3VLO7e2
WsQY8Ivd8J1uvP8Qn5Wi5XAHbRSDyM3zJ5c1O6y2i5SFO2/ALEJI8NxvNW4ufXtF
aef5abe6dE3YXlgpzI62GRv/5+Kt9WsoN/NWm4Eg5aeDPKd6cXEMR3RdkF3taFUr
qL98Ohel0o5CH6uDfJ9K788Ao8MYTN9e3nzeh/XkHOYqdovRq/wsq4bU2FN/dktG
TSDeFMREeTmhLq2jwRwxsRbfzoV1rp5Zku04dmGHRs92f5smf+BXTidi1ZOKl5/b
wgjqazkho7rIztm6ImCO6VsOJRhDEQ7fYemZrZfov7uqvPdzFkR5GUCrYQAPABtS
dzv0uZmHVjJLbTwXCjuzQ48+R4DtyeyDr61fD/e4MVrrXw7lsUznVsDrIP4HJUXT
jAhdcP/TFMiqvTCYsFzTQfG3JbeB7yjMihCbck9kCO0PZUgZGmgwtl0nr4FgPUDb
GaSTGl7GodDLee/v2zMoeL8XSdYG0jKEk8G7wepKH+dwJRymH/ipp7paCFRVJtNX
Zps0F5Hc/7rRZ6Eq4HVn9rFCSPcM88VvZrpaZRxt4fZVeNxyhwWFJ6u0deIY2MiF
51cxLSsyxwnyZFYM2ur3VeE+zN3MnCf+vaGK1b7u/YFrBT8xfpuWRzMuFWCKR/zp
NNTw3emhLzpYVN5rxdL1cVSUB+6/6kk4QblpC+mRzWDOzPDtBeTBcciH0Cf/MBVE
vjtvElyNKFwoUkY4Zg+U/UzwpOp93b+qxlDv9eFoIufMJpzU4kd79BIzsbIrUmON
Razo8RPuvNtYbORMJcorNgo/Hwd5Ihg7SGAcgujGtDeV9885iw8k4U6GA8Zn8XaV
FPt2WPjKPMigaw9HQP0kX0sme+c6pePvUx5Oc6+MojhyK6IVoLdxi/dSQnrc9Qzy
O0oDmMSEqJcilHrif5jiAnAyKy4z4d7Qja6UeVfpmJuSq49DfFnHrrc6NBb2vWGz
YcHxkbH28iI8BIsZRMyBKDau/FaQVULaMKM84ErxTOcv7613KCn2NlCWdXFwcK/u
2Ag2OtIeoUlf4nOct8V5u5dm3v00745e9hQx7sNRgYoG8f2Sg1Z3UVM52r6IPZHS
Zb2e6Gs37ORrjbfqYWS6H5463FJQV/PkTRI8wcCQ1aRwTpKcNuN3OuVshh+AX4ij
4WOSz0flXG4tEW+YzDVf/8mZB0jTtlFJI6ktVb01xc6sx7ED2AVe11G0DpK7mXJ/
fxZ/IneDjRzOFpBaZR/01bS0JMZZMZKwKy2MDSrdO0H9wnrgxwVhK2zW85QUFSbu
n3zDLjXqx4P9Sqh/CArTo47ZZghJ4dN1ZS3mG8ajRR4ZmvZ4pimbLHF3Ozrnxxrs
NA4L9cpJ34qWzJu8SUa7GXugW4J9J1tkYDKP8+wF3F7ad1KSpp3Zi7csy17jC7iD
Dj8U5OUc9IYS54pULbxl8xryFq3WdR24DzQMhhOfgJGEwGHHRkFJw0iNrb/RNTMT
Vzhpb2e4QAMKG7z1Hj+IA1yyAyI8OnTbEBTI08TwQLSBFfTEBvqE5gqjNbPyCQB8
+Y6gBjsjhFE6il/rTZYnOC8rjGYtNIBxudV9IU5fKRlUuDetPzwmhmd82YupScl1
K24nlpvmzzUn4wM5WCsdfs6xFoyH7s8MkjrUb5A4DyfyqzRpnPFnskQoASQIWmPv
o/v7Aw8yz0p4VCMU3pLnLB6t7Zjy5mxUkj0GZSWwOB50cBzwfYlya6xEIu01i4HX
/KWLtXqWFeMUG1j56SfIFA4n9IylvDn/VXfItEUJNlUAcdLurTnCySDFRaBOJi1h
+qZtNEjZ1AwSKLbEUJ+5hSzowo+LAsAv4b17Aaw8s92JeT4L+qU5bYsf69JHpgTs
KhhpfAQl1skKDgUuSZaMmA8CICU9K8QGNlibP+r1B7gDmsbzfIpPa8Dd9Z1OS93a
g69ZTpeeZAnpvTXfcSIqWPmWCiMDbr3zHQ4RTXk88/oF3UDi8drq3K2UqAn1QIGn
R4j/Ixz8Vl6OiWwqACONpyOldh5rcdGZRxXgS8vfeQkKEyN7+pKEl3r9fsbQlszv
+8ow8MDIZ12SvgZo5kW+9pqC+SD+lj8CEDG4dL+1aP/0xfzC2EzHpcAgRqcH2hmu
DQ6jyVoitwZypyIvT9t9Yau2tggoFh1RN0D6s5A9obvSN7015YHy8Rgc58nuZ2SP
vI3zScuGmYV4eOa+/g5woIoF49dp7zhnHqso3heaV2NFInkRFxB6nNJ5Lq/mRf75
6A2ZK+BHRsW+EMEvu4K3Za9xHCROM4b8PMiI4kFDsGk1IdnuuJaL/MMgijfhyLAx
xvNA50xNs7yjW7li2Yxn0cx9Iczeo6aONkA8iUFwfdMJ+EWjnEet+Wf7euXA05rb
HYz6HZUk/K0lZzskYMpos4BAF9BLhFVJXVaSPdwn9706cofpUflIfi3auEeUO9bg
f3hhvFRsOSs7sPYLd1YI1y2UtcqyorNivunTtSV1TzY7/XYf6w64LptGVYkiZqa0
7NjjkDWrwo9poRG93yWP1kENIFYYFwA7JIk+NV4M8PU1OdFJMd4JF0TboxgEK/nY
QnQmTwfUISo1RNbZSxklTdRvOwjTXuXdK9dpgK9RfH1nLy1fTD9gjCA6/6Hyz0J6
pouYV7KKjcMgQhBf0+GXb5Ae8GdR2rqCsSnGbdbXeLPDKzQoqq/ErnYme7FflK3/
QTEf6LKR3urdhXohlNYYG9Whot8o0jwTWLSl6fsS3eS6EhzAAQnOS2mLNAQsDivw
Na1KBke7W8iF3CAJpcmv3UES8+GGht9wdOqXh7venwjYN8BX/uEnb1Uasqig4W4p
xlfdBLYngKIf9afVCF9TyqePr59a8Gat90l9Rd1zXUdx6PuIphR0mGwvZYgo5EvU
s+8/dszixEFTJIxBXOWocVFNZZ/2WRrToI1yygvZ02ymoJ4n3M/tQeRhivWoBXTM
clXE4479nX3v3K4aV0aeW3KCFRfOELohUh+wnPKu52P+QBi35yTekC55DJIw1hn3
MSAt7d/z7GJRJL1exlQ9OEaSxpRzUvtmmhEBz6mjka6xIvrk3dyNtc4SBMCNFtOa
6GFKVEddbZbxB0yV2lSTl+oG+9Fpqwxz5H1mFo7JyIklTKIroCLMJupgTzOcu/LW
ECw54x3tX98dy1zmX4MoRrmWi5TQgU/y/VJYOColL9kxPNozh7UmwVzurzntk1MR
2VVAMCArOWZhqz1TtNR1222Y9xqG638Y22cWitLbbVM+5MvtbMfHqRSDCi7WoEB7
9AgGYK/GR01yCFaVxp/9mD/Irg/VJU/q3thSdzG9xVm6+6dS3ZRRW1QvSwPZCLyc
U0P8Yty0o9sRCtGFH0GktkTbiYhIiln0ELYFrX+32HpYu7rBPTUh9KQFxM4+NwKo
E/+RzXbyYq0kBqYbZWvZPyNMLPI0l8pBP7B19NPat0SHaJlKZnYMYY/YxLZxfjYl
qCJazK5+snO4cuBoe3XpmMOqXBDk2qDmCeuJCFQK6Y81RJGbVMATN5Zr3CoerxiL
7/SD4f8AOVR+TZ/IB2Jxadd0ooIiAhdGCL5UnNxcEm3NkJZdqA4P47P2EWm2hlaX
tW81A7t0gCc9ObZKn0vWRE4XRbbI+YW8zfPgR6hhgCelwv3L0yAwokd2iTCdu/wY
asnmWxAO6ByXvawosGJrgKuDHBQH5mBa7C1m1h9gRbjt4lK1dM24soCWXnIRCDYn
vl86XOH1fdu53F8Y40WtsLqSFy7cu2ArmEZTWv8TBkF3SV0DP4Lw2Blq/Zsji6zd
OM/S/gomd/lmvig3SbPx+hHx9QFMny3r53/kdeu54+XIt8ypTSnFY5bsy0ZJ3HeZ
Pi7tNgUeowxlnL50qtfw3Oipn+IOspT8PV9ss82+JMka5b6NRUF2QsI3XSz5wQTl
MkDJ7Mi3xDJUBpvTj8oJSLTjh+lj0x2vI5wGrdYvTLupZ/bWXSIQtf7pTGTOnLoX
Roq54+WlHPasNDMM47UR8vvOLmM8OqSqOEh8OOVUCvipEbeo9fxS7VeitSWxnR7Y
D/45JWfbCVdV7ym1r8v6UfYDhxPmLEsCecTGmLSXcZp2cuqdhyeWiZYbtLFKmFcu
CygTZzbU0QSI+XJVQzPmcGxcgOu5BvlBTFXI0AdaVHF4AlQZfoqOEKpmoTqFkIQl
nuEICD6KZGEBxDsFWnO73Dl+SxUVFsAG7sNhfFOoXxrXq82031ivvf8ybpX0C3Or
GH4qekEsoEVwEbHyzFRAh0k0yVQ18ZPCWASbaERQiECztsBhzwNQKL4rjTAzpUCi
MTPYSqEqDkYlJWgzbqSm/v5hW6apk/a3plkcrNs33cb3RxTU2nTL8lkJv/Ow2gyc
0Vgemrb36U5a44zm/PU8dCFrm6Tnzc/Lk6IcLnWf7I+ngqGHO8zKXf4ckFTiI6Rp
4+mN/CrWjAIK14khAM8TT3b8NL3KMuNJi2LBZzE0iwE6Ywi/YgUNX2+p9ZXxjG+N
Qu+bNSAnsvqJq33GIsAYkeBV9zT8fNPGwcc0lmPg65AzSI8sXAvk0zL4rCUlPQs5
Hnl8dUdOgNZgF2RcXjpjTll9m2zBfSy1HaRFArD0FcfI02rYNhVVtlSIz/7ZJC3d
YzG3SMYt9UwiB9ZcIfuSDJscZv7USssIeHYkdAc9eu8U0m0rHWQ6XsNj+eL5qyZ2
YnOdmpjs5FsRq5WSxWIGmYNjxFlhHnXEg5zt0RiNTNdUIV/aFXfZPvEhI5bilkUU
mUft3QB087F94O+tDIAmKRWzApdXXgDtrfo+L+SlQuZLobThbeW85kFK4jSstK0G
I8EqZxF3pKQGhitltqYw1IajywQCIK38ItpaDlLPov/S5jW2irp1+h2UO7L4WGvd
QuGT6N8MxdYCc02YWJY/e8jYvpsZte7J5wHvVNOhuW9uzjZZh/lCrqJQB7GCD6f+
EH0WmHkCWp+2hTmS4e/QDFjrkHl7PXSONF6SNyhAqrKH7gIUHBxvQJpY3I2SrM8J
Xx2J4NOfZDyER7AzAelWRc+A5HLHwZAPlAdFd0yl0PjKh0RCVxrpkjPTqKvKADfN
cy4nIoEGjKElaLoE4tEGr+K3daL9tgZ4qz2y67HinwY5i9hGsDK6wszuHeY3RfC8
xGJb0Dz2GXMEpaKIO9HOsFM3VK1Til7NuchIRRAZzs/wV+tFu78voTHWRUC2cB5S
cFqBGqL/Y5kcdOcdDSc8GalRuAyQohYY/KqrkkuLBin8F5mGyXYwkw8jKdWPZz2a
73om1snBp42w5GJLJRqK9Gn+v77JZam8wdX7iKWB9+fx9hN7Fis7zUU/zd2Yja5g
cggVCGPboqKe0fLpNBud1iXZzOFKRh5tkeBiQdMm3XutsG7xGqluEpxerxFWcF+d
pMYbAuVWClDFCLWXUhUB0GCjTVzpUR+PvxdeEudMb4+sodc/kUYXN22I+VRXC11M
G93ctXl/59iwuFJKDoYCu0yGcvitQWopd5EY5FEYJCM06fAFtRCJBearySQ0hgrE
2i1Fb4sRAR5k4jdxRuaeW4hphTgOyJfuEmyUe3F8T7pk0nJun/iuya+1S8M2VWFU
YLflhVuth/I8FMJRTAeZcfs1H+3Xz3UrzmWkShNGQQC0K94OEDYvLXB/ehSu1ma7
EoYMVtkzwN1J/o2SYMhLL2hejP3CoV5VNxf6+lN27DcZNy6HiHRrTZqoL14hd363
Mio1cdbGdKFvOLi6fjQaDO+ipdR/GnbCuyDA8Cy/jlVJuAr4rQup45MPf2GSvbOu
wy93ym+hNmWkaiPkW6o1s/LUevbAM7Px+idsBpFzRq3Kuynnha+Oyk6pIIYwgfjI
YfPOQDOeBpffJFQUR/zJPUFlA5roJd5yjzt8vUl3CHCWMmeDOPzH+KQW8QEpcz0H
tRMrDprC9dxS+O8RAT/QB4HAdgOUsGiY/h9BvHayEfnzR1y4DcyqAAd1z1lGTiTw
rw/zP8W+cJdQZ8PyrqCkUn6t8tc/SwjPPdnrUoUNGCWH8Bcn43JB72ta2rD+VADV
a6Ej42eMOsV1bK2LsCbA7AcRnC0JqeHaAJHzLg+qSPUduNQZiwF6wktVydzrh2oF
Hs7VSBHP+JE4iszsHiKSbR0del3QmRBkLi5BZv3mS8EXtm77o/yk9pVRbDG83FRK
FJYiLgL117FReXe/PEEuBW06jLeMaZTCwW4WAAAsoE+B/Npic5yzMbocMFnmLtNj
4VlUh5Askb8TYKGHXLECX5uKpECON9XnYyQTvJj5zQDrSLRhB1NA3FDwL6Dqe/QE
lg1vg8eKgNJb6Wzf6gNghfzS9LLdywMTqBgEydAI13NYKjN/8/5uj2Em0gIPPXeX
k7b++alT7wYjw3Tbc0wIeTk+kIdlTCw4qVyA3+IuS9prjiPTY7wF6TXg5vx/LpEF
Aoy+MYcjMrTCa1gdAjC/mou/b6uBBkDieSCYCWizjzQi6MacVaV4cys8YLHrJfPG
As0R4BIIIW6f5JjNvCrmdftQyitdGGUaNEke56z8ZkcIMX4vrHM6M4jtMOZYHD1N
BmGefb1FhU7+sA9p0pSozUAM8Rs0X242qCfZROFCfgjShwzec1tHLhAaFCRp/do3
xIvmrYwlBzC9ZuvHLqTtWGAakJY364UyKd0PNQ2brsK+jo+roazqUnlrWw/wisw5
z2yglUSzpj2+kmIE3SdY3aD0s5Gbq2ZLURuptmyZxF5fADb2JMwRmFFohiTZjg/Q
GrGjLf7utewSZbRbZaIFuEJiJJl5R3gVqW+g4o+XqHO3iTNKQ33PJvNJAXkwACEQ
S+mOydbTmwJLebvuqhKUKUn2v46Jt4f+nnG6b9tGMj4qZjPOsLSxuGsEFFOHoRJJ
ewNn4H9akxyjELzTwk2HoGKMA3KFgZnTP8EMMObPSdhFOtXW+X4f1PjIdgObKTbk
X6NjOclvxYDWzeNVOzOZSZdr9f4CBD5LyaeRl5XuXC2UxOv64NtcfYxKz46ZLaQa
Bch7gKuDG2hYv0n+rZEtewRtLtSkP639tYJiEJkA7l7zEvWlrbE4P2kdHJmq51Xm
R7Xp8WjUTidQ50V9VXGr18EWrZaLq95nHFO96ceFj9KZuvKDIz59h8qI1/+z/FSi
Z+s/yNlCcg0tOcq6iooPiKaol3R1+82u3dOODpc2nZr09HHDDq1QeeqCs/vpm+Pr
77j29ZIuqDHzrnKINcOv44PO4TbRkUfzIO0ZTk7MS5I+7vzJCzL6qBeWRl3XPDvx
rJyhdnN67OFPpKYYigOfP1+KAvYIrtqHWYEnhaWcnqumhgEyy71Ruw2O2IikCjTN
NokqiRjaVX69ba33BczzcDYNkwDOR0Eab4GfiuqlkMlkNgGJ3C/A8ML+cWt8OKkH
7l8xJeFrgE481KNKj2njIjrg96aEro1rdpoffWw0M3ZzGtsVs/yMCbd5zWoxBAvs
kQLxPuSu3YAmIwt66b+F/3t9EqOgj/yXuWisS5c+dUOG2QrVzWUXysRqprtdG+9z
Gk1tju5G4e/1sU03X+qLEsFzyKjwGQt8HxGHD5HX93JG89yHHvWM0cMiSN4lt8Tf
ySPOBlHlKbNO5jOKZQyJsi1XJGQYyM59ueLRQ1TgP+gCLrApQjkfru0K1A4ejjjs
awghyRpXE8KpCtO2dlugLgRZF2RkfBWaSvpOJDHT1YALskPU03hI+GOEa3Zvq9x3
HpGC0DioJQ/PpT2QI0C133bY47itykX2mUG+JxR8PQveAchNi/bJoKVTFSNj8ReG
KJlGk+fYcuhMeh0hRIHAHO91BT50bGVZ4Mw55lLDIfdHVZi5HIJT/ffIgBE5ppsx
2E6iISnuQExKxSpuSPt8oMMn8KiplaDm5m+fcvRap+TdQdmeMQf8KLyF1DlhHFls
41UjDbo017rsSJhD0TnLEybGvZ0y7PlHO5rYZGAzgHcAerwKfCN8x39EYg8I7Kr5
GIlasGlmmQZQI2sjaWftFrLa75PeQkmtdxPeIp4oEXeaMdi3qIJ5GWXPL3Ldnth2
dXzVct0Fpd8A770c0W0NXNe2NnFJsdfEo7FkVspAQFUyQ0dCqw5vcLi+0mIx4Q64
HU0yAlkvC3aRtmtSu+G6P3Wm/7rUqQRjkYenScCmiQRWKHEZKAQnCiuCGix+dXcm
35pvnovxKfm5tKowxPsn+e4zb1qrZ+EMhxyWkShRTMnL82VHyzkNwqz5F8N/hKd6
xAcwpHXqcHgX4DW1hKlkCCibttoquT+ZT7Y/+eZHMcjm2j9gL20ZUkPqgLI5Fb56
jiUvrnumubuocnQ5RfpGu2zbleEbXXMvYEYUW4b3TJKEL26ErMD27jR+7YoNZRNy
ytnihG+SIpXeAsZ8Dl0D7POzyjHg38YzZogvF5zSHHiqjOwRzkCy0naTqoQqGWhg
zMMVd6C+6J8Kg5lvbkMU/siAwjhFf19XsoWix/9LkDfaawjxM2J4N+Y5TEw2Vjtl
dVfvIGKfKJ7XE85ASDJ5LUa2sCSCU6qbxxST/Jf1Nrt67ONrx5gSrqV+EWrhcnoI
ly0NkHll+G7PlkHKvURPot8FO83pKCI8NtZ7dcu6mw5fPJlY4a9p/OcIxZaLYk3f
NufTgOsG6kWuQ8BqZGVUhAPHChNc+sjwUZW2EjrOxTgXzWpXrE4Fg2FCQimZe+RJ
S/OSRtqPAFI3uUFB34p+vw9J3eyD8WC6nX3DryGzCuGBjvHU4p4HlmY/xMn54j/c
+q1LScDsfWDw8t7s2fxprFwXqUODbcWtgHEjIK3Jshv6+r/o/ZcanhrycxI2n6II
WwpecMpRgepU/3ZqKRQ1kG4vG8dfzl1TxTO/iM0HDC9gA/Rl6FKwkAd2hNJM7b/2
fCbphbFzXyegMyGr8HcS2+WhhSMk+7ZwsxlcHyEUiJrYvr0HLP3erMSyQL2s0zsB
G+leSMG4dWzt00MNNKakfldIpHtYhSLI0N0fnNMpmdKHF6UDD+aerhL8DkulIKE/
Z8sQW9WHd9Fernt30oHnJjNBhbeHf5q+T5DNfo6V362hIl6bia/1Z1YgAlj2qa6k
p7R4l2iGlzhXf8ulji0nqCWXKUcDEDZ0KrvSan6udbttTvfom85uYgmNFLYhrdzo
xeUuYoBLqvSYQxedzMPdYJxvAbFvS5hWXgfXFwoC7AKaYn/jLV8GsTeKnOS52vxW
FdQJG2hJOSYTarUK/SyBR9kLljc6khMF1F2/Idpx3kfeMHblkjGqkH4hH8QkOw/e
zvFrADpimm0maG2rsLzWzRsSc/IRiojMhj0qm0DjzxqjPTvaO/pw0Lk/vIdNzqUD
2+8CVInd/pRzOyK0j1AW0YONR96Jwucb51rbovBiBFANpD5cAyzU2jRibRXgBV2g
+1ilgfA0YMq6cemNkn8nHH6n5/33C4fqLvXHYbXLOq5z36EzTB5/WXDbm9h7OXl8
RbQ6phxeCvaC4Md8UoJ17EybdZmdbgbdhYc/pCml4wN8isC+djMuIoc7cYOQ/LTd
9MatbKwmVHV8Q681atUOJGkw45tIX9wVzSyWAjgUu9G1i51ca/TU4ZEamRTVtT3h
eLnN3q6SEzx6h78Wu1N6e1PxB4GkxxYZHIHYyHQDTreN1Q6pVmgzdMFAbHVgLMSM
mzTY/txIOngnwcFgruyfBW8sulQQiriP0rYnpLBzK+5P5kKK3ZDR6of3UeNRmp1G
nK0zefo/KVOivgYHsOmgfAX9glSZF+l8ix3eBSi+FnzKDtLSx5dG79Nc/uWTQFMU
bowLalhxpqKmn2oAQv4kPbw/8nie8nfXn1NLmzYLq+IsxISK3ZRM9eRgBwzYglBQ
n1oG4ZmQI+T80md39xtKI2WNHgzOnV8dGidMfGSEerqPNyCQXLfQFxeO3UmecPl1
9sQOCSLQNdIh6rjv2l1mWp+pN8i14Rfo0Ux+3FNZOl6g0tDf2QBmuWxJ9TNRoSIA
I8B5ykfA7BsXWJQuF9y2+ssgtwzJhC9ErbNQlvEUwEkeBg7idGTj3oV59qhOZcOq
TUK9Oz/FuQaD+4yRXgzz0jlRZ8Swqb4tUIjdjLeXDgFIB+gaYbE87LF5qOvh85g7
41NhwRjA9gqNwox/OLp50VcR8gJjT0dvvRJnnEZ82qInh3aehE+ADyeaDH7/91kd
/Eey9FGgGUXLji/AVRZyoY7U7VeCoc/E4x4iTk+La9IJu8QtIobCu7MO4Zeg09WN
MFllEwadNIsYVC27/pCW56npKrYg+7UDzhmHCTPA1IWFmWFkMcrS3mVbmx3IWOHY
tg0mH4EJm2tzUZnmQnQOpnvqLTovCFoibpNotYvSxGEeDPjJwnp2cOIHfaL+6qGW
gWl27foLNDVrGPoppg2etR9fFPqpBHCJaqCAzo1FZqPFw9/ZuPd5qOtwsnxjAifc
4r0N2MuanZhuGKtXRCyoUdcfMd2DeyWGUbW7Qw4R0kMLU9TNkX5/UVoHd5Pe7eep
5dOc5VUro4FX5BMtdnL1umQb5Ep6g491XFygcvHsx05h62d/BAAOxKDYLIE/wWia
lmDXo/TD6IiugWsaIgsn4OPucr15rxaoCnWDLY6XRq8l01bpexkmpjrhClgeeH1x
M1PiFfi0WwvV7MfhmoYrvniV2q7RdNlPGwqjOvABxfEFsiDJBeNDsgbdPbxVhfg+
W1w7ciOJrcIFllPjuib4/3PABDqnfWbaESpINwErli/bwf8AU5/X2UH0ZC7NxJJK
Ujr3UHxxuy+PzHk/pZ3Wz0C5jsdtYXcmpgeUKhnOnInLq3umgCl/lb3JUdUW8/Yq
vGLhy8Vk6sDE8K0U/ZQahJvePe2ygkYh50h0slgsyL1OCTeIu9wBiTablw7vE60O
HxKw8/z1u59jB0G7RZCkt+tRSz/x7YCCLoo8ZWfUvohHGpPkEjy3L+HXJ91rThN0
p8Ofi7kW4uXlSF/iYa/HwI+mwKjTClJT1Xs3oiaYTkXviOQ0+wkmA5LuQCCpLubD
tL6ofRQSn83tn/X6QIosiQoKqStz83p50r3OOrxxOHdFgDqnNcMH9eybrujujltv
LEV5+boOlIhZaYtxBaNBiemZscdBbuoYenkJtXEbFsrUgcLuwOukN1/q/YWu8m/u
WJEhD3KxFXKxHRblPLw6Z+xvTPp4TY8kuYzNL7P1LnSlzNA3mWxpikGzIentBrF1
lEWb+COmfzwzoWRBzVNiKfpEsbAxMvQKaUUjIhBDaOBO1ZYWyopDmw84ADKu5vJ7
KGOaPKCsCgpdHIIqpoXtoprmycD7i4/1v/pMXfrTjmJMXdNhAtob7BBrCFPIAEsU
x3Ce7/uyYLKlQTUzZHFGSwrzeROKPdb+GlGdIFb5+qj+EPMyY+/QxSUA1xFOsKG0
zvWW9Ey1OkITkr1/aFibcVz5M7Sp6RibZ71ViZQhpUQm+fyCXvRdDDm9WOsFQ9qt
YjpqPtXGBlN5xFzBiLnOhmmmlHV2NbYWB12Hh9vgBplVNac7A1NbIOnRdk24KiYR
qjEWCssR1sQczRUp1S8Z7jximfeHt8B1MD9J/y6B4m0jHES2/cknY45K/N6xkA1x
2ZOX+i4jQy9F6aqttV4CzI1uEoZwS/sKs3Wez+zchRlscGnzEny6A3kw6zSi05Kc
hbL1Bvkk6J/eN8v7lAm05e4xN0dIp43ghHiLRwvM2N4Fv745ENwB/hJbgf6PuJLR
YnjvGZmLQR4MPBo8jgI8ajg4rsmRT2o50hZRR7y0Aaa3pbViFVehtyS8nAeoc17w
eLdrG8q8lZQ3WQIXGzy5zpa6lkayUPY9aF16U6dV+QamyfLZTHD8o9ApcAo9JfVh
7un58meuBetgEyEjUQhx6RMuRC8OafMtsGjOsFN/z083ZEcEn3T3STBSffCRUZQa
9+Sd41vpta/cZ5gEAJUPPqjTmZX/xqrmcUpeNysFex51BYcIIUseTf9lDiM1gr10
/quUnN2KVRoptH8SrDZfvZHJEarkX4TlS9grd3AlKh7IUn5dYZgM37Y9OLRdpvnz
0KVaYhBLcrLa1cNnw4A0BuZUl4E2FFOTvLgT+AGRF+aGrrnTCdV7aP9Lqw9T4chP
f8k7p9Uii0VgwvfDc+omLvHBGrhplSbgrCNYSK0E3pHepEZKAthWex8DrRwpjfL9
mnMBQj7YsH+ZHZqxvTkPRwPyctyw3mwqmYQxoFWKJG58NQnUnYpxVfZ9BCWwksGP
d7837NYn0IGH3mCNKDdwzj3WWzAZST3FOzPhH29LbpuZS8n0tOkfW/yhECo4cmlB
F7gmHZ/19jDQB7F7sk49Trno6kZei/fLwMqmtdxlUQm587eP5eYnk5H8GaaTgxth
/mYtIchQ0ZafWFvutIL9C/JfDGGKiYIkQnMTUhH69N7qYDMGAKLomiMNuO1bhame
qC6XIaGTExHc5p87n4NevBn+HDQrItbJZJhTyNcuTk9rf9jKv92VDnox8ObP44Hm
MDxwBkJxSaL+U+H9d+KV0R0CeVj1lrxGH80hftjySAv1uIlvG1Xyufti5INeGy3l
Y2g7+YJSNd2vIfte6/fFY4HHzAzBLr83zk9xZs6AkZrrRkl0MUcOUDcO8XidUpv6
O1OI+EOIarK7jeBNLS6GcQ+KOBcBENNrnObGcxjtwCUks6LJ0LsImGAAToOEXmqe
fPY4ofN4efxkgUdAMWqkPRzW5er36+YoGvGde35EJBM5yOfntSHiMoiDXoaPOWxr
xe1mUAcH8P2gOCkAbhl40hOQcVcH/XKtQKcurHfmEPxdvLpQQXn5lfq5Js2O8dg3
dBK8bfvkKF+7BFRwb82l4EORu/JOnlL2m5R+JjV8WkbN11h2LCXSuF7rUAFeX7hu
36KPDmOiC9I2DaJWbE8+BOXslxIKUagDl8OK7k8OIjf8b0ThTEf5Nb5qioQ+OG9P
d4ox207n6P3sgv6Nk5Nbrse9e0ExzhYsUriEIY9ocVMuLSj0X3YS02ntjg55AXyE
KS0PZXwpI3rqUjtZmThBfO39EhHP3C7jCgW/arPnHOjwT6zXup4b2yMzJFQEiqYN
q0DVG6EcMSdvsXC9C1bHLM7DbSfGjO+Qf7N/2HlnUylbEAmY6Oz/G6RLQRC6RcAH
ajhhmu3zkHkWK3KLWglEMms1ozAsPNMit8vwsXkbSD3pEcIwsb/Hu0os9OFqTHjY
9ET0uVkFcJ7BhiV7ZKG+n69yZJeqXpZqywZk6n+0xYtQ+hdb4+T/l9heEwi6zsVm
z+0DZwZME/7uscT+zlo8RmaxvNAVxqyPyQF8Dwb6BpS89DyyGWo5vsyRLFPbZFlY
hGmwf9uLBFQy7ya19J2kkEeT5YJMqL3nO7eos7i8AItuHf+G7g9mtaT5uAxHzmx7
Pn3h+U5vEWR5ENNITojkBANyJCM2AOphA5n4xrEfJfZAYc2f7NFN2jn+DJuflZhy
FqS7VOXAkAa6uRL3z2Y+LpMDNwKhZXqWritlwvkDb7iMwr2WIcRpOwygdzv7Y3On
1I+w0SBNnuUk3uEC6FnCuF9ewTkqJUJe+NnjwwBxyJAWqphO0UsJiYFvbHPFRKCM
LMIrTaff4UGMXhOOhBA4XlieHjlW9faiOP1ztFYZH4eyZuNrk0RUslVq4jBkSbS/
UDNkHERaigaNtT441Y5y9vnXN9NBN4uQJLcX106tXpQmiL4p2YvDU51WbrFdvnkz
QliDQZh0YIGpYPZWU3nulTTZPADI/2K7GdBHPzitc3Mj1z9Tu3Xn640QJOiHRJei
vTaEELPsIzijLo1WZqT3pa6VHA1VzYdBE0dsgydRfLKtTjOMIdGAOM6GxFmq7rBS
6uz8eZN/MZ07DP5jXfkijjp/XFnGMIBf6codnJpmycCvu0BVNjpEqM+pWLO51g+4
lbIkudI/Cu5cP5EM3mwBeOYPscit20mqZPQIKbYQYZANB3/R534y9X37ED/rrank
nnptbuFjM3vnZ0YCbcEsprfcucNDJkPgMTBudT8keyrYmiNqBkPlDqnCzF8Zthm7
Z5SI6+nt7I6WcAl6aiA2LqZ238pjlv77fWexmChQg6lJ8djT7YGJrexT+/3jlZLV
S1jEPkOpCdAowaErJve2YhSviYUu0tknFvF60mRBlhuN6/j1C/MU3MUeNmjCIkiw
NU6jX6E2us/UjipmWDQv4YvZ7ivF6/nngIyPx9yWASj30eEpyfM1f2fX2Dhpunsq
35ih6zlOTBRVFt/fbW3XK3tojvnNr77o61Zb1IEuF7Fy9ROzifHVXmotY7VUjMU+
F0zK4/8K1G/DfOYquvxzKsirIjX0OW/dGdaOYG1hONwglrCO5sa+Jyj1e058yE+a
RTZvruQy/d3yZArUWgXvXYg0EPVDbrp02ZvXjfow7rHlYe/AYZ1MAYGiiXRLC238
lqPrhtm/T3dq02VuZ99V1paQmrq3w4/b53tR3MK2W/XQ7yjuc4WRR+27sGyTJSML
PdgCkcc+zxbSvXNtrjb9SU2Z3APDkVEmxPkm9yu+hG9THFzFYkw0RBYSK4Fo8YhV
TsPSshei8Ym9zc58ZWyhhlMYxhKyNKPtE1OTLm3t/UJPrfRUFOswA3fKmfqJkZlp
fXdmWUdYi4EgClOw5MpvJIE+V5JfWw4Bv0x9oaoo5cFbGfMn25s95j7i+vzjBGnT
eN5gfhct7sfHkctAgf0lSOUslS1Lo2VK/OzUqGWCjqaPJM/lpPd1RJ2kSGB/CWS6
QYCdCyN+xRkWMEDnDxZIdL+XVkfalPaU26wt2PZsxqK/jGuAvauJEcrcQXufRPem
KHXr4kpVhcXeYWEWEyCxJ2stR31M46XXnprsZ5T3pnHEUHw3Mq3oJyaWBH2jEkne
Ki/OEzj2jzKtOfcsFXD8byqBSp0lqfsRJ1BsKpidUlrtinKDeP8EoJZZeR3RzPy2
/bPyn2ix93jXKDCCKBK0eG00P3f9dc90LEmsbM3grs2Tf5T4WmLLwX+hYT5nLTKI
+rvEQlgAptvTUeArtfyin/azZ6GcNqald8hBMrG+pfWoxo7YqhqFbv2egKjj7Cb0
XC9/BfiWTGnLEouyWFKolTXa3PiMa3xWNufRMSA820StbSbZq2WMRtQHKRjLMADT
i98k4UFJ5TrjivHLanGkrgpIacNK0ZgS149Dg6OpBr7xH8d2MW/29lle/052QhwY
WGHq5pYGjHTsdJQVDpu03tlmSKnNHGZXtvW/QJI/gM3A7KRevV5GVQ91lpmgg3fB
YY3w5uHiV4xYOr+RPYDxRF81315D2MxggvOoHjYd6MLaehgQEOgCd1jnFmYvOxol
NGfGoR+VfwpMmIAXO55xiVbNkTA8msa1/6+f5JphymgPZqBqJtwvf4SYf1eSV54y
nx8tQtjz6HibcTnCh6yzupgDTlok+twbfcpgweqnGYZ+R6HlqrpYWRx6rTSyGhQE
CdDkDcy7Vs4swXaf9njvHGZSTXxsS8TE6YDooIDudXLVfJCBf9rycPpMIbc1f+00
s0XqgrDD5iB6zqEMnjiw1Hm3Hl0p3pLIqAsct1s7XW7rANO+jCs8G1cnzO8/0Cbt
41MjBaeb4PLgq7TvhfWtvBDXdQLys7D52AWNL7RUpQQwzUXfmMkKY0hQgs18sjJd
/IkMInBcXFrISln4QPMAhc4Aqp1D7xUu2/MvOZ1uLG8WNBuMrA5ZVpXC6lDP4aZ/
1vo21sZ8Y72xPvMb/FpOE3d9zEmA8ieeFKuw20Tou/CfvnDzxG0INIMjWwyTbwIt
BciAGjTljFo9E+WCNZOyCH5S1yan/0n3UXNvMk3TLWKkTwZYyOei1HNftGCJvhdh
jxT/D+pl7N981AC164yzHOHdZM6KpUgehW0muS/8CgB6TziStKwhWyqLdinaqiMb
bf5LQL7NJ+Gj3PLLtkxnlwqeuRs5eDT7v6gjY0Jy5Kfg8vfjdy9gS7PY6UuB3CTD
WGIh2VYDFRYqSeS5E+Hj9R9RXJH7PYSJ+Jb42DG/OY/+bH8p7GcL88tStWZPFvMF
LJqnJkqRRo/0dca5m6PGyVgTKJkQvb2r4uY5rS945nngJ4A77RbVRjnxV57MYOOg
Iy97jqKqnF63uJRJwQfMmtZdQSeNxSeNDG5CAZF/zJTkWC+L8zlcch1gkAG16JTg
DaWrm07sXGxT55gt3qBrb1/yVu+IW6QX51U9BQY15Cknalc9ydE/lkYYLmYbfysj
l61Zyxjxj1U6/ZXuG8RYEN8qc4IC4yGOaRElT45g1F1UPzbg2TtXEah1hu/f+H0A
E2Nz8o0Rw/hstWsa27Ow+Z0LuLic6+QDAu0AGzGMJyq/o6Olvxre647aMYE4EmkR
yikXcWcLK6m7/S0HOJqxh0ShEJOB9CgcJHGSQRuYPCOOODFSrpMFNo2vvFBmnSlf
zhByvD29Jwlb+P5ssp0sn9WP372pzbD6pAgo2bBF1+c7nuNRqaeyMNMzPDxjrUWQ
Oj+2Ou06QYbdtTjVhPuS/kYQjgAj7/9NHlY0+JpFsOJDkQjlSLXJ6Pkpu+dlwyOW
d8sw3oOjR5+0I9FzgLkr6uM3dY3VGJ55KjzXzWkMec6jepWzcEMoMZcOzokkzAbR
1UV84KRxZGhDJeVOayJwqjrbUB0jGcjULFxS4yRuQKNI6SJAtRJT5/5gO4w6o/g8
5F1ddHXr2Rqmv2rrLX3eWtKIvLQJPo/5/mr8kqI5B7upSHXbfPGcAp9Ddj1UW87c
SfirH4vdVkyfrpDzTZRNnbDviedAc3rYeJkrNp38dUE/pTqUKTV6xYn9hpY28a4u
sUnzV0CR9fTXf8Vag6QVvjOzs9OWfAHeNsbv+Q91X45M5kuzURtDMi1Ln+weR78A
3+7YJQDNhPbTR6FgFmgx6bZRld9WZV/6xsZ4Ce5G/5ZFZj4OcBKWDSMqLkc9K9mi
cbeSQfNBBGnaIyW1OQLvGJ21Nlk3OyJrpcVpHLBQKZK/xbX1fHPIShVUihGyIDfk
n0hYtK85asCiYD5d07wFGq15qQcuWJq3rhNlQgRYkaTOZSgU2yQnXsUnBwCJRXLL
smSAQWYi6rtd9ZBPcBg7VHDanmH1L52ms4KQha4+71fyxehNamWyfC0qNPkbXlIZ
cwfZtOerdEbIJ5OAyPXnhqzHe2b9K8QTWsrG4pjmh7ukIq+vUPvEhDKMzwKGoeSu
6yoPB5jXzLjgIVYpQxzosj0M/9huhP0IiBa+1EYnvtiULE7aovLDtOeFgdReaVby
RLm5Bf9tvCBZDh1K/iPaUIQ5ash7YHFEW++UJAkEBeA+YJ4ardobTa61tq2YAUAm
zOd+G4mFKDfRRvcREcxT5E/Jx4S4bBPDmWMBZJ7nVVGCeuaTklTbZTgO+My9p3Wn
l/zduuaqlgU/DQMn+Wk6CEJS4DCtCOF7D18bok1av/JlAmUKAMfog4MW6n/L0I0d
l9dghi/Sz7wVA7EqScTWAogE8YlVrKNKaL8FhvH94JJMWA4SS6d5KcnY4PIeoXwc
gp/68Y5YLcGHpCCSwL6Bd8g+bGgTsCYPNk6jHhDmyRL1OBdWq3Y5ZYBBOCU7UTZw
tKih5TbC4svkIgRWAj3ULbkl9ZVLl0HjUPxe48sYQ0WeeLAHbuSfu1/Kl+9bwqGC
UY501E3OsjK5Rgjcd/8mdrOiGq2Q5mQdy+p6+xI/ssfh3BogMZ+6kKjUjI7boWr2
TlNgRb+J79UfCz701lwJfIe91KCiyXkDLWhzGlYZEDvopk53SFe59waC3FP0Komo
fDg0mB+dAdmWr0O++etG6SQfiwrHGUjcZUEnXSHkzJiYqEi2EJu3Oom8kTYj7SuB
wKTRRclTk3c3TUDqF+jtpPaNXg4Os1wMCrFR/s91lQyE8UsHogp4nnmr7rPNJkX3
EcZ6aYjCfO3Q4ixowbjRy7nmOCCHq1+p69VmOCei5UEa24Tj3yB0LJyagkOg8D8T
1I8xfq2Ctk3PRrTvncLU4rKDnmpZvl89L1eO4fhHuLSM8MtbEtiDaKM3kbNkkcDu
GEui0GfnkoFHYLz86cwVSjNH7ZUynYsgWKOVhYEbU5TTULPRVH7Y9sbQqIMqZpXH
QccsXRLSo+2f06uCbW1DNE/vtGqYe1SxPGhr2yE3s+DcoZfuC2pm/5cC8myLcdtE
FbEZ8jzG2cc0Zk7Ocx3tieYitGhthFrxIQABIWfgeEoHrtU7HXxdp3rbN01fMI3x
qoxPPnVwdsUAbZPOrIqkXnWrNcmemnCHAezqri9sVBRx/F/zRQaLrVLdKOrKG2hY
YIRBttb7t1BoCGnWOQ7Rk3O3HTbg3arQ0af96ucmaaQ7mzcIbx28YQHWW6qkpo80
oA0vsQ/4Pxlu1RiyvJ8BUzV6zRT8R7jWJ51IS+wNzo/im95EFWqbAb54oWvLaGQ0
BcN3hIft4bXjUgHDIAhlrLJBTybg6JCsc0NzxSiSR4QPZDWXdzLIP7JgWS2FcmOW
uXHJnEZVOEAoEl3iNXptmSuXspGiwr6Af4yE12QOuxnKie59G4MZHIARTTwvCSkW
EJpRQaf6khTeHwJrqXhAmWpOJNyJZFtTt56ogr878wdZ7eSt1FI2Sa1Lsc8gqoha
5YWD66YGbBBvgtWuT5KDg+TSN7Jl7IvPWu4pESexNvZ3CeLrhuAgijmiBs8KxWd9
6P2vE9JG9Lcoj7Sm9P41lr3G+3Z+l2YRyuFbW/ip2EYTSKOziDRFqXNPK9cE0zau
a0OST0CJoD/ubdg9uq3C3fzdlH0pOyFfdHqW8YLPXl5jk9p4fY/W5JQH5qg8y8vk
NRyNw0/74582zNiEMdMppuYCXsoKtfQ899LOpAgfQchnN1ZR4lBf3Lo8Iswxnc6W
ulBF/C+Ay53YlBXzx++VbePSswIwKtKaN9S93YagSgH6IzoyK9AnYNagniuGjR+z
B/K5+BvWedGeOVR+JwUCFx0sSY3VSOp8+H8q5M8krACMsDUaJM4S0Kc30ZIKTG2O
fSpWKJIfWCc86IknJjHZmVDXkFG7TSw81oeRsIlFf1358uTiznYwOgTdL/IiiyHh
6puAQh9T2v5q7S5NwITV4VgcfyNkoEe4ga2d4eh9IlyXD+iLOJybOChITjCycShp
/MBtPjj45Hrp9kETGnmcotjOoi+X1YhN8H5GwwpOvV2smTetzDshVMPiV9xD8NDV
xXBUHqKK2sV29nrtAHS9p5FyZbT7gealtmGY7Qc4HX3kzQGMM+OL+fUqyQPnzScJ
8rw4NPWpT7yRr9aqXWnz+ByFTPMyRIgGx/aVTZFdmv465/Qma0JsavLEQNWVVQUx
xk05pqn420J0f0borhJiUfv89fXiYYbVS1ScsnWzh+5nDHfJZX/Uk/XxdgXP81Ob
EtpIwLT3xDIFLlIXF0sZ1R+vCAcuAbmfvqsArni4qXJsT4ltZLtsmLaCHmrwoiJ7
Pfe6kZQv4q4cKLN1l6g39V309hHJ+3/DWyhSGYzWeFyaFRQ6qNQA8n4ySZU5Utoc
zBKfqL3og3rlYs4KYlPiNwXKNACnR31L7tyz1XinMn7OucZFtt/xRGEYKJI2U/2H
fkLr74m69SYaU+H1uxY9sgERPP6oHhZ+fkbuM1wNjx5YpXOXtxYonKYsyDng6GEM
k+sVS01Pd76ixBrHqCaP+PSwBerv1WwvPwAfqUXNJYXjPH1VoguS8QXYVRkbnhnD
qT4lizdW/65Wfnu1YyAMfkmk9nGqNYJCi5ujUaUxnWhsoHR0k69dNwbDAALEuZME
Wy9VRnYfvC78s0fvIu1O4N27ZSljuH+gpyHwg3539WLwIAuoovpbKYYDcyGcVQW9
qMDpTSqhej9mvz+xzSMBBGePtrph1M/MrAqDnl/Mwxr9c1B+uBuKtZSKD2CfPSZS
zsNQtUZ1pwS3U8InHCjWRSKKJBw4w6/V9PrhwTnWJbPpHP52oKpeadaSjEcabVBS
RRqRFgHHGN6yZd2Iaa7JqWyTmCsyRkNXVE9uXPyI0CApO9+Rro5jbKrjDCOnD3qt
gAKQX5w2AlAmCu+sAJmXisndpvmz7IcKDJoZmYm3MiQjDv6muByTgdbVOJBQ5Kia
no/bZnqW66hQQTKECOSxMp616NBytzWfvVTG2u43Bp9qbFCgPpXwaSlWweVIfVWs
GxsCtO+acP3GoyQFJdl4Y6k8gWM0pw6T/S5P+scUNULLcMV9jj/3hYWEeTtwuzgf
aCGknf8WZdXCNJ6Mr94lM1dUKlv5EL+xXuKugKWZDIUuHfGzFOsU0+qSQU3YUtNZ
J/E7nkg1pT/ziJOBv26sIeypU4vtFjTlu5+ZvtauX0+4sV1BGiEzcU1L1Dmt2Jvq
/7xZBbK82qOi+ZK+lStrWnWe9B1v2MbeW1yb7l5D9wtgZpXuA9qevJtT0DaFROIp
00wtcB8AFITUEo4pncnqu0d+DmBoXMhvTeSXKlOLf8bQuRuSOaIJiEieMBcL0qYZ
nxdk/VZ8PEvxOny5sDTzgqbW3/nq+kCv1qYiW+rDleUjaJEfA/K1Vq7snnth1svu
xgN2gohO9CmJyU9y//Hn2jaWq5Sn/fqHKOPA5a495JzLDW0+ySeJIH5MKSwvrU2D
ytXCPwQigcCR56CIR/1bKlEAu9pZqzD4zhLy3uYeIRW7oT53xhN69PHy5W989ps4
+QRZzlynS2zZ7owm1RybLWqWwO97O54AOP76aSeJDzpvT+49h1oZkxyd1aq1bumR
9LKndBeUdTNB2mKXNEfLIJD4RiOUCQYJhHsOz+FdVmSxKO00kgH4Nv4UWTz/EeZS
S3taqaUPYdShZP5dSYiCkIQAHU7cf9E465dw6sI+M+940mrv6MfRuON9kpveW70/
blXGg1wgvN/LhAIWsxrokT0KK5rsYLiQNyxhggz8yi6uNlUFmNEAu3zNWUP+633E
yq3OGAToMTzg8jpYHYZ1JX34kEl3ZmM75lPPXp1dfEa9mg6exZZ9x+fg9RVxFYDb
x4lP0QFyo1F0q7su/cHqU91uvfwcRQVT2N1bIGVUViWPMGDXy51mtkbGDS51qMfI
Sa+FCanc06uiIgxtbT2N94eytLMpn81k8hDTyzavWbP+Y0kTzyAAXO52DywyNdBS
xuznZxAOfZa57I9DoibTph8M2DJHvnwMZiY8+WCiQiLUspHcGk/30ObfwU2T0izO
wXi3JdFdkYNfU0I1camFG2CSDXuZjoOWjkzsotBRczLPgJiJVnSMhpsP/oaDPwsO
q5cDC7gciUk5GdcGA0+edvm0GXJuD/oz8aqfBO42BhxFX6H0df1P/BYRx+T3Oi+8
k+1sgntcJASqGqAcbX8zi2hWzXZOVRx8dHxWO0RyfvvlcKtZ9yjQ7NmE1+QoenBJ
ULU23UKFjIlk1/668rWqvse3PZuzF21Xwb4q2+xywF8P78pCv02wIOBdUxvAi2h+
/N2VMuJKk7UH4xhSpMZzBpGor/RSrYA10D7h6UyQyu3jlpY7ChHu1NEXv5edmvEN
3NW0qW3nf2MyuMDI/LEaoU6RMezIOyhRAicjTTU5IIgkwginF4odtVHe+G5UApRW
j8Un4Nf7+5+j/jdoCDWoLfWFK6QrNmSv6nwr1AWPb0q9yO9VoUOtmRkddVJ/N7Ay
3MRmqHff5HTky1+cOyj9ReEfd6QN9wlG0VEDOmcukVL9QxxlpGKB70Gac3JKJI0z
9f5xeP8ZMLUfN+ChRAnPxdroVD1Pa0LWyV0pLheJWV+Ulonnf3374pLSvHJWNM61
GFhKU76CQX5ng8Mf9oePfkhiFsvvbMRBuwSAoQSwhYeCW2FmJ2JF6r+5aWvKFZty
yiEEGXa9ORzigZV/S85HH2yBYHeMUsjptLtgWwizk/ZmNbAg7K8dDQGP2tleRPQi
vc8FhJNW5RcUlb+yUs7zkhYMqWC0p0HcBtYr50GiXv906B1VFHLQD4nHYwxg3O2p
yALJJpVgxv6m9xe8hrzU/TZhAZgWsG2Bn+P9N5eYYZlfXUYEbR2jPjXZIQwsgccF
W6Euy/t4uN9tklnZiR5al1DYff6HHym207eLu8dM6LeeDtI7B2/mBCFlfX1ek5zk
bbmYDZKn4vij98EFrZaTq4VDYkJSzQMm+AvcXEIv5baxz5Vce+361tm2+Qnm1bME
roup0arhJ93ubVN5sIkrO8ts5Km0c3g470Sdkpb7GDjASgEIG0u4tTLuMG+rUKBl
v0uKP5rSgJOwagwmfmWmZ84ckQRB2ZOMIrUyyNuY9zSgrk48HVglIeSC9gyTWKqv
s8VYhq99+XwMhcI1PdhSB7etXGnWq8JpYklX2wrBtJNrc7YV7G/EVH0uz7BZ5lBM
wTB6Fa+24pjRlfhAUxOurEz0hxVtqGU32zi4w0lgzgMfYJmzeg4423Mtowyp8l8E
Kl1+LpBw+deVZ0+V2iGdsavmlyzdr6S2z/B5+/b/iOji9vKQO62NaLhTlG6nEYTb
6ov3kbmvaJk6MwZEdrT1izMop1CcTJB/oFhCvmfVT/Pt/8D0Lw+9SvEaFD72DMPf
TktWYFcbehsMKNe2i+HxmwI5pnbOTc/Fs5wYu4y4LmmDJl19lSRIuSEPBkpZ/vvC
kkLMWnqQ0Rn1FqX52yD44dTExYuiLHuFu7EGixM/QDNdjbU9ms1ZB+FkpLc4OtY4
6xwcIzPXJCiruVrCMq5tp4ZVWuPEA+CIzNKm2QW2Y+Tue3AQ1hGAYyvPfa5YCzNr
+QVZEo5SmU20gJBntz5pQ3kXTUQpUdhimPsddD2lhKP50Vhbbj4jM9tM2BgrABcj
k4GirmvYDcAauDcbj8dnjaqW2SQi5GfAr9PTdVQScZnn+KI28juwqgApf9KjrRYI
8Y+mKFiz6A8UxKZ8LPoytgXn5eXk3rSgCOOZL99gpt9Um20frPD+vmaeSpWAWdfS
AXE5ny/InTykS0Hxg/u8CW27pRkgCTpFlVRmo4QzXlBrF5/9SQhFqLJzBzwux+X9
I+SrXLlFifjFqanxQZXrn21Nb06Vad+dpG8V21TRyCbcnHPKEzNuiU3iKgCh1FzL
1+n5pJ2Tt0j6U8EY2f52VyFPj3+BMokVUhFPhnkAPZmHzEIZMZcc8HOEZysPR2c+
Hw2g/JB3/w9b50hIdRI0aAyg7AC3rwuHSQzHPBZKYibTESiqIlJ6nHep6c7067hd
V7EEx7NpQUcZSTfozXFKQPDCBQz3YJxPqejTxQjwzULAaQ6B32MzazAUFSAYqZSI
1/OKLlbhCEjgR/LQLcr0ACbKcyqfADqnxqy4z8BdmyNTLy09A6slw/jEPQ2MOBIf
6gJ/ID/XefyXnJj4+rAkIGhPMTXKhKhbsP5fEuC6b2DUH4FmFJi/9dd/mWZB61FA
Lsp5A0eYuD23lE3PiawuSwuRUjtEwyDRWxg8leUE/XR25zWl54Mx9ayBWwuj67Uk
x8Qs45Y0dH8trOzNHycgylehk1Txw84FuDHWgN2RZkchtcQQ8HZ1T3wPrEuDyfWo
FBu0LEoCSmPSZgPFGfCNYxd+Lh5dk6wuiWN1Jk8jyZo2CsfDtGHxrVxALAVnz4Jf
Nnn2Rwd474XXBXUuAF1Lvgvrbk9UHnTXHDiKtu8TLY0kdIeImFF96ktLIRIH2ZXX
TE51x1urlLKjy3+Jg1Fiqu4v2L4fvPxZS0gqJM5KaCBhuwNqX5gp9ZU5Y56RjUWB
GDUocPMd4FBE0gyi0nXBdIMd6A2aufCjafzBuLncUCrewjtr26+oivG/KLuYt8jj
UvA6PAB8E6sM3MinH2gR73EZ7mCV7UR48meNHu3Rl1ia/eoOPOJPwQ/dS7EGmKTh
yRFzWvA1AFY0GN94epoNAUqDzYszAwiMQfpG2UaSt8fU/F0ZLDZINm8/ehZE/eS+
9av/CVkWgHjH2+GGR5EC8l2H71IGoRtj5fvzIWg1Bg3dmdliWRc05OTmJb1lGIao
O8ndp/0ZbvzWrhHSJb3Vbff6TpyHF37GUdTKROsz11uwdaVqJSea6BuXhA5oQ6pu
g37hx/vrhpQx6lU36jlfVQIWMXidToz1Of91uQ1+S9V3I6NDgAKGT4XZAGKMwLeT
cArZ4tSWr/3roPtULqqnRUf7HW1pRF4cSRlanfXly8nvNDfYtR8b6/cSl4+RJ+ym
pOVEWW87PBAj9o07MraHqtdMdLhuWUnCEKNLWx/193zMBLWBYM5n1/8dLuPgfFYH
voSc0PYNzFt8UI2mgzpsPk42x+HXOj48ixKeLpaW9VB67vzVHmegXYlJr745yUvw
0NNDK3x9hLzrfIb39l3fkWTE/KOVyP6zBArOyXescxl8w+W6L6GfgoZ73d0k62A+
lNprrsRVSXUXEFUINn6HgU1YDP3LJJ3Y+S6cImj5WFqKWQfGeVulalUg++Fe+yZV
pwi+1/vGKK9gTUgt7UAp/xHeci4ekyRObqab/qSlHdCplLu0D7khTDMQkTwFHqf1
mGRl92LPqpNQFzbO/S6/lQ8oIrjkat1z86abyAe94DT98wdOs8+at67baFHJqflD
JzngrIYbRaetRO2TQAph6YJv07+FZH+UXmD/qY5YzrBpByZXVPCE2cW8SqIG1vem
j0k5xLrF9KlabkHetDDtxAucCmX7Xu/bm3Xcz9V+Pe9unxdPbMSPHOjruhOIQItv
LhUMZ3E3m/8PzhMfA1ZjiJsiAZjQWmatK27ttcg+qQ2kWq+YErqqm7DOcG/a/Cik
FiJY0o7FFt0A2uLPr7WfveLxRUuyyGfsHsjQd+WeiA1rWRMB8+ohK5hbVIMgCSPz
CiJ9pkSuwDLj3WAHc7447YDVopd+L0C4cIm9kRY7bblZlW9p+W6G5nFIrGYjWArv
UMY69WokkLb1O2cwzCYGiiBCfBy1JrOQLdRMQ8/Ww0iVHikGiMXu2Lq3qxmZUYcI
/5dJ863t4+l6XGDCQyA1jxiEHJ7reKqDG+sKWsi/2MnHC+zp7mPKZgyySo/eSBVD
3tpKiiCaB1YvvP/1o6rsqa4hq1Nb6bE4zk3rgwMXbbOFIFpLCHVCb31AKJ2FNPWu
a71djgNubxksugqdNDdGIo0S0qsroDuDWnUVCE70I+K5GsHbKiJ9zWA/2Sm8CRBR
hab3y1obZc6kk1NVr1gtQQ8SLF2a379VljG+O+1C83Oj3QwbTt2sj/K2G8qne2Q7
CaHAL8+aJXh69UTieRSln2TZAgiDtFVNXy74ims6OoTWaZgZxoRofYZ2YYDPm6AB
111pBFo26TXbsWAPnM1taTB/WjIiDvBp6/0QNnClxb6X6cg3W+AV/xp6LiUB3Z57
7ahdVlVwxaeO1UVZI01oFW1Fj5hHCxKiwb22mAe0HjINRKC1JO1ZiklrVgom0lZo
a8SOvjMcgKerHBlZIfYkVGs/UfYUHDaMRDTsJDeBBBdFtz1p8ygQnX1J0uUXggSu
9rBQhNgbJK5UskOkq7lC9kraAhTgTk13XKHn+4JC2HOW1H19lKd4NSj1/g50OM5z
/o+THopN/x0+vgOWv/DJySMdemLxH0bt/bVQxy+DlHMG9YqY7802txsYFJMaqniR
Av78NTBzaLLVWRNO1Yv7WLWSdAGodd7L+QXUrdjJl/ouGX7jNadKc9CxYeVuXO4b
DA/dxs4MOUEG70fnYPqfqCOSCIeJWXjNCofSNgMnhf8Om8VQ2N1X4OR1ktV2E3K1
ZZb8Y7dtay+VMZv5xX5/0obGJ+52CNm2S6yoKsbUQcftvSnFnYDwfBobkZhzie0Y
z20+JH+IgsQ64xiGBXN/H1NrwXNckeWy1D7amhBZvI/M43h/qfb9L0inhGPdok8C
iTPcToLhNhcLeYxWeBpMgyLL2i78PPzQ7/cQyf6Uuti3BlJUrXelN+abcicveoV9
fHEQV2hNfX+J8nVdRsYOBG3OlDFC/xZoLcYnk/w1SYt8nZ89CQt2dqCuQSNOrJHE
H5STr9rBGW5dkh+AGEcrgi+CQPG/v0Vebb+c6CoexF2sYxumG5L/CsG6m6Vgnshs
G4zm5cVuZ195MquwXhFZTjhRk7mQFpbeddPg0Keq/gp4FN5HWIVsL551Kypm9NH5
RZoKqnkiyWjLeeIPglJ0C7MDz3x3ADR+ACSjRV8ZclTTnw5cZvICWqR71/aR+goJ
k1GkD8U/gdR8sYB/KdsSxxSmgt9Fu+TXoMkOgkkK+VbKCbIGVCbyDqxqvg4CeVqE
PWF/kI6+AywamND0zK8Ri8xWG05xpviw1A0hhTrHu5oasN0xuFDJhXtYoQvoe3YA
PTYN3Kp1xpT/RzULY3STyqgRuZrErRe66JD4qHLeH6q0Ez0E89A95wf2K9azNiFV
4NvkeeFEmxqNYITxiCwrp3zZlPfsIHSTbdt0+SgG7jlklxFbw+8ajaOJSGZshUDO
qoVGJYRbi1qbmEICMPL1h8ZkueqWyL1819hab/0cpAWpeFlPFYIlgNgu3EhnBYzP
tb8JavCTcZiU3W1WijYM7rjiwGLdtLqp2KfDqEZdtNT2aOCJyb9u1Z0/yiQmp6Rp
6L380082sIL2vAtT4wxk5Lpz9V3Ix93MC+J0Plq/l+RoJTUITbpgEqxXFZvIDN37
R2kYnkIdWqDj/0YM+h+JXeG8UoFaG8yRG0MDBpk+fDCBZnCN3n9h2LmWlryb1ZAJ
g3NNWuwf69GH/VPveL86rO/o4VSnIKT1mMDXk5y0HBZDukQPIMR88B+8eU2HxwYO
+jlM+VKV9Z9DBzupMG4hLiDXh0vguSmuPKkO1Q1h4UKjVZFEywzDM7xB/P6A4Qra
6IS4i6SJTMuxTgRw054w8PAECw983BS4mJVCEWC4+FYQjkpYDC1XUFtVtjjCtdJe
198O1xBbcx8grbsHexSUCnCCWYKRTl2lh9qnj6pbSApBPmPkGix66SbODP6iZgn9
Go1w+GH5FQLvvR4Alm2ncOg/AB4yb8A8C7g2GweGoIrSfXzZZ9uDfW4pnM/mgzcQ
I3zX9a/npISdfiWhWT73wB1T3bsi9tGrBOwB6+XkrP2d/LXWdDW/AJjcC8YpiIU2
c7kbks01HNxLmR9q2uUTJxmJgfzCDMFv14Y0i00dipaEo6cqKjMng+kt/zqoqj5F
GTdD9IVxLZ0OcVlJ+Mym95e40qzr7TW7Ve6OaolRlHVP4V3XHV/nNx0TtEG0V98r
aWJNJr63P1Ezqo9aS+qgU3/GCJGT3oTc7dHBF5+G8nrBejsW9GSu8yCY8KmaC4Y0
J2S0D3rkogfvExUPTKtAg3q1ud4SvozbSvrjlOmuZeJcAqZivmJmqJj3IDsExEy+
He9+1jUU1NN7w19v2EpyaSwH5n56Qq8wmuRb84WJFf8Pg5Of406NHkv2l+kImhZG
pC8YUzGD+P0mkI4NhLpV5qEmrT3huLPs8uOB2SQMMef71IYqdi9fakJ92ke3vkOr
kZfvPxmPZr7hdexCj6Rg13IjCBHAF17OBryWHir6T2oH0g8hlP/iUW2Xh7pFQgfR
zG9R6pt3ieVaZp3alHkC5LJCNnNxAaaR+OmiwfCJWWpstMQJjlFwVuupghd7oKwa
LK7WxdVFFJcQANnhouFI7ldKFD4hLRxcGSulHI8wZvo/uW5gsdW9S9OuyOI5p7ZI
8weY6fFeLiuaTh7IrQqgh5pTiz189E/OXVRx13B0Kbcrd+KM4V8v/zZrxnpBfGLn
Ldwi9/ozqk5bBnX++tA6gRXBr29jsxnA1MsZJYJ9gfcwYa5tmQ7CeRcBYAHjTMaQ
YjIpV8V+m/hDNcCFPwN46Q9mfBQ/+JIJGXqQkFCMP48l1GlWTnVKCb6zgWIsWP82
z4yxHp5p9x+uEmXgstisRM0hjQGasTl6gyqlTCtSCDYNQv1XSTTLKZVY3BxTTO32
45EKqX1zozMSISMig1GAaEaf3U085LvZQ9BX88bCPnxKmDp6LiVP5mhd34lHEt1H
hqJsurUgcJoNIrWfU3vM23KCjIMwbQOo9MChh7XQ80adi9ebfSzd34UpvSrtG9nq
Q7sQXNwVCVC7MVzlcAwcklhiFyvHv7JSrDriXkr6wGbkYugsb3p7sPb7LsXuQVvc
Hx34+LydG4SMl1KFzFaa3dgPuMla2EQjwWTV/z/0WRQCbgX+tNiAK1zEMOR0lZOm
PCbBnxYqnDhqgbau5K28wFpaPT+f1GvhlYYXUNcyZ1mb3NWtPTU2ulHAZpS+8hme
K5zyW6AIbD5Kot0S3rBBsnXLHHx/E9QVMbI21oHLKLmpjShjLBcxMNe04s8VEZFD
DszjJUdN9Rt9pEa2ttj1c+lmvitcD1zlsvcqLQN45InlaVVqaIXaQW3PAN231Ye8
USfuBdA9slGRR/VRBRB/lCVnIrX1Z7VQSB9ClWAksbeRgr83y+uITu3COzc3v+g2
mhI9oSEURFJoHjHBj6QOXD6twoM6b0uuYqECu6FTmKrwlzFZ2evMVdwKJ4CcpuEO
XFPVZ9dvG4WPE1rGJksdlbMY20+81XijuR+azbR/PeVNXrULYzLhoXz0SncFMk3Y
JWB5wGOLzujnN8MfCk+m7l8cW9wpGKuesyrMLqujMTFrs60g0mO7xJ3dmHvdB/QZ
lgT23tQ1iDvVZl/NxxtsGjD8OvE5cM7xgpmoXMQHOhQTrQsHQxirC0ZyXfHwWg+0
C465LJ9qJ7EnoMw50EW6wsR3uCS0W7+5bBT9t60tht0Lva8F8zdsZJ7OIRBzpdQI
eKCXsMCoHck3DW8eo1vEithyMGUIzW1/bPVyQsNvHTJs63m//gu1UIOVFn67O0Vu
U6vEvVmQ58uCvjpdY1LL+KlK35o8XkYeUZ2ONQoU/S7k1cUgOowxStzGjXGOov7H
wv9mdQ9YOfIVbvDWYqKovWBlXOMfcuOQ9SMtillk4Zr4tl/o3XE6edub1bmsoxW3
ncjl4x3ruNisVVRgH94ecU0CFk/bDlT96FBWl2jHns0Nsbp/ETh1F5Le0AEHXpBN
U3VBH6oPqsOeRe5l8EWyMcV4j8ILgAezCWaOK028HJOGer/aUAANBY5H+GCGYQMT
+HVk7YSrvDU1SoV+MhfLjPXfdBezM4WTwSR90QegUAw6qyVGi26I7Q16oSfVfW/9
sWjgwAUh9iTkQCX4fGcMMtNvHAQ1puUVnoLLq4496igcGip9+RbPGTFsXIPtFHVQ
tiuWN/2M6xFM7gdfez7Qr1kzG6ZbFazy9ZHHVoA4/JgieR+BNyrXM9+JFwzimso+
yV8s5l7wsMYRDYeJYlJKojMCm9DGp51CZiBgbkS0AFGtRFXysWGrXloY++6hy6Jo
/clAQAVn/IFMXsg480va4nmjJtADDFJDkwb7JE4t5O7a2MNVGHjp8w1Q2s1KmaKr
ENn0FVcBD3JpRGan9zIAwD2G6YsMNdave3K2A6BxXfq4TRzDv7/tQpef4WgPLuxe
XSsusgVKIcBhwzceW/4qjMb0GAHkzzfRrRLavoLbsfOfKvcj7Vk3CheeaM0jcRzz
5Dr+bOpz22OxG/e1nWXR/FchET9Cy8HfGPMEtWHOdl4I0e1QCR22F42gTqawZMUD
TWDlnbGxA4BFiSbxlK0a+/wEg9+0NBmtyk+5p/Noz8lswzDEdc1gjKaHu42Dj2kK
u4HcFWbZrAHSxGM6AJ6976USUng3SAKnJUtDlkh4105wWFDiV9+WUvWDT8BF1cNX
08lXjbLhsbdqFuFl+mHEYnBajbL+TJTMiOAsNBkvVZ/nZqUYmh2GSYd232IvXF+9
6iPBxtqm2ayZWyFctmbgPD3vgYKvdE8G7ueSfrS4fcTIhZ477cRYzPZ2pdGgNbRU
6qg4T5WBvSN5eXxyD85US0YYaCewupDLZsKSKVwYkZp+D4QqWZ/8T2HAUMuXuAy4
VOYaObOQ3u710FiBBsWZXnU/2gaYoxwBpeIU2C2clT8/ejcwvl8gTmOux4sPziZE
IeAFpGWo4brmA/subYiJ7FvwyKEIjI8rvubPd2bdg1sV0qS++F5IbaEuwNvMNdTF
pYfovylQ/ktlds7sD2d9PgGCbCeBKa0lF2NlGc0mFC9gLv64rcyhjM2oGafnBJaL
TAmmaPsoEv0CshNR7PV8ukX02VGfl4IpoqES70Fb326YxLAfFcoPo7G8DxWVO1x9
8QqmcgwSVDDw3PePM7memIMqNQz7xZx6oYEY6ZMj/mnBZ326yDAeGbmy9puEE/by
cF8Q8zvFmqDV1mbCCEDM6PeJvWrhdn+JSOYGynZ3mXYlkY+NJDrFZzVVL/QzaTZo
+3VIPHGtUi0kW2oXx5Vx4Bb5oh+hjlwT695fRmcw1Pw2GiM6A0H8+t7GILTor07n
J18ns/OZ+v75mNCjKPveQUBDRypl36t7QO0hxspxPmsR9k83nPyqdeYcx6Y5z7bj
Xg9Bk4OU/WBi+GjrSEmvMbHR8wBxD93AblvytMXTZB/KOYXiYNeeBYlHg8+cIbzk
e68LdGoJnE1AiPM5/V/lDxe4sAtYOFXz6g7LXX1lMyj2E2nnTxlSiJoWvN0L+Yt1
sIrjS3jxTrDXmAzJtV4YPBBmUArn+HVwkkugZ0TGId3R9fRNdD3znA32KpKH3xci
csFVnn+Lk7ZYz58zTsx49ZYP7m0b1YLdH+QzKJ2AZDjFkpTvepAKc4nGK1GA+kts
CNlam8io4b6ZHKN/WL53RUsnR45LlwMiD5uE5dYlad2cyh7EuC4mYvlMC5IJH4Q1
wjBOfp0hN/8XBGp3SE6QfrrZaXIFrr4mmhpadg02dT51ssKulZj3t6dIqIjq/YS1
APnHYyYfxUUVH6+PgxYpRBCMC8mq/J24O4aB4wlD3IlwYk/DjFGrU3857Rigmp3m
yVMps2dHmbGS8Y9fyF2u2LdmwlcOZtSRcJ9RhvK4W88F3XRIzjRr3dMnj7n0q6c+
iuv1MoEccOpi+tVgR47aRg0xcoN8NDBcpIkhdp/39hPcQACmYGoF6WefsvISwQpa
St5qmb+2t35bFzUs9pIdvBJZLiqXMmtP3tSsWf6P57ibenfgaywusEtFB+ou5lUF
1JU8L+AVrC2v0Sb/hhYpqpfe5KfMJDW/N3P8cL4o55LnOJ0KEKXNU8sQPGkz8zA5
bbBNUixVGBkBZVV0wVaA95KcZH/+2IDTZ2xUzx5WenbV4ozeU/x21T3hUuwCOuEC
iEaPUgXIkQ96H8fCYnGTVAOEX6IDrcjSZxO2dBnzu2XG6uVZh5WkisUKQIih7wCR
ALqI/FEMtkzun1bG60GZWgNGDEf8dVQuqqMdxXw5xF0YtwG7YO4exnczUzKUe9r3
iRq8N2TU+yTNX0nXfDNiAlqBXGWMfjHoRvq9UuPtcfATS7n2FXdKfIh5UxzP4biY
uivrIsoZsIZ/QnKtOhjusksZtdUdR2ZV7yHa5fD1tDkHBD4n4y+wnEZFmKojCDq1
q3ZpmWZIQoKHqNh2ifzW9VigaQddyFfdxdJ0yHAUZ51NnH/jQqBQ79W6tYyGlqnI
Ov7nr8zWIvr3oFynZaJ/7Fk4IUmQfYwlhCncH4VShxHAkQrJTctEO9p/ypgC464w
5nO0Me3zbnySMEALjN1bOnpr+1tcKgh4EDtl09W4D940PCys42/hkpRlGFFfXA2f
jFNK9DK0fmXhTt9CkIhtZ3uh4BQdQtXuup50BdbTTo21kusIWgjoVgu7ggJMLqEs
afxmXtdwTdTvY5kzMf0xBSuhHHxcsoBqYYSvKhagHxJntg3oQDNBdeAR1jaiWybw
7uqypIIA+1alcNEkEkVW0hBoB+GrMNna2iUzpr95svdfhiQgIRXNYRWJxy8Gagl6
HeaNQJx1wMrGNltQ+XQtfq2K4IPuK2QDeF6qX5iegB1ZTJF2DpAQWVbCw8OOk5IK
vTYGCQ71Wb4oqJy7FJt6Qgg73beLEfd+Ugh3BP7U9J6v2FfCdsikN9BQAwFCwLJp
/KzXhlTtLkKE/EM6rF8BwO7zx9w/JOJcenPZER7Hdq1a0DLQRV6mYd8IzNV5WlO/
Se4wyZxTwK04JbFtCvMGM/FIdSHc1qZAWt9vDmK7NuEqOEDILbIPxqVLlNwPiPHh
HmKyT/Kwqy3rFLHfBDxXl+EKa53l9uPqUB3/TK9p9iMyEptQIFK+tG2m9ZbD47Jp
tcshNVEDioJQFnSw4LMjQbpwRlnvA1Ui9MpTLMw689QLO/WQJGLIW3arjuuatuZa
EVINwCJ09EoQMcjth48M7WRVpAIjwpO8xnoDooHyCFE7BqJwfjG/m4ML2AiJ6DJU
+9i5825Nhk9T7uQCRoTMYB0be6JTv6FqTbTB8jrWVApDuG6cz1fUlA7IK84BZJda
5kp/7hyafxVG0e0hOUKDur7Hn1wIXg3v5mq2uQEr/VMdJbAtaDijtB10xwqRpzpK
xznWf4FNIgb/3aKHreMpxNmFo5DycPPHHmTNX2GfmF67EXBMqmXtH6MdSARfmhHb
QSS4nzUTT9CQ8ftfbsDuHZ6KS8r8PCTbsJIzYNzaJrvmT3Ejz2wL+40ue9vOdGhY
SirA3S66jndZZR5htokae4g9D3Wa7dg/Bf0g8yFQe7dt+bUgSPxVqUxZuUEJ50em
H2tTgvEAr+UOESBsJ3cj5W7twLXQPKiHyeX/Zjj707ZzaM/K9CENg07tNE6A+sCG
6kWKpEBr2K1C6koElJ9bQZwcb5RGMXyUY7wmr9B92iDa2svQ1/b18im/SU/hanN7
ZdgTKtEQpKCOYyDZQm7HEA+cckVKPyZn4ngpFX03HCcLmG5XL2Fr0TexZ4wU7oac
P9UgDw3+FECE1rpGrULsXJqOam64YSYYs76EiO2FyIhR05r8SAEh9JUF1nYmpv98
F8FbFvy1q+vTg8U+xyCabBpsLcMgnz69q8hgnYhuv/DeqyJW5Pgij9KhQ+Q6YSBL
6TJXlygfGxfcm75A3E3vht/vXqV4l7mhcVMWECHRpmBCl9j3mEr/l6Gn/m/zKACT
Dzpg1k4aW+8+Am7NC0Hz2xTKFYiq9ZBwaMp7ziBhjT5u/4LibwEQqq5KsxIuW68b
eulY4yhcEzu/zXMhk5/+OhcZWLi14+/mO0VJ31aFi2yrkiqMsiZhKh0aRUZtQhUe
wJqxiD4lFRa/dOQMQ6nj49+VKSOZjFykiq/yFhg5NnhrYT4sPiNQ4vXgC4sn8+q8
bTY5blezAf+Cta+dHMhxhWHDarPHg4z4iB6qmY/wcshFgkOCnRB9bSmgkfeLFJux
pJFDTjgU65n59vG5BioD9IvjDm5VACRNusaDzqs9eADSJWVLhuLdXhOehWuHNEbA
I2Sg8FxVrd/uPVbtuIWjQQv+H5KWujMG+5s50feyvR/Vh6Gme6WcxtgYV7GGKT8e
Vrx4oW185TF4ZiiiPIHEbsUl09lopYcP4hMssgzjQa5aLQ6MCzWR63axfm4UkzxD
7FYTbZR2KzZ6Hx0cen91mxMAfeK1zId06jZIsX8Up2wX+oaCTmWH4ffkJQtmAFm3
9Vw5x9AS/LCcanSZRGNK+YPaaStJGuZw1V/gsGqBM1IEKufGRWJe4xRmyIH/AuAf
ABdKXAXUlweB1i6vYtn+1DHN5/8LV+E5GDGJ5JziCikKJRbabu/3pptfe2MRWOMu
LKDZJMhBDQwFRckP0pEdsCNrqJCEffgg0dPcwbE/MamEQ7l0ZD6Usrk8RJ1F1CJ9
Lsg3Uce9SdAh6cfyrgnR816k1Ir+pYQifvUaiR3PGcuNwTqV8noqUgySYwwGwJ0b
QpIkqPjWY1qcOSsdCrZeOPhZKiodrp/bCgEVW9D6euV9BFFBaNE2vFUPj/xuQ0a/
UTA6Yc/SAjWjIMGKf3rfHZgPrMRCKvIIGkaR22XVQ/oiZRIE8dgkVWoNNzs6UW0K
VVBot+6vAdh2KfHqRDV8HwrlMoWZHGtg/RZy+TJIUV6gZFaXrHXSWy04sEV32DSx
T8llf2CmXZG6eBGNYhb7o2LRaj0gnzio2PKD7xwVsr/uSsOmwJgmEBLEZhSSDWyj
oGrFkT9hCMN9niNh/fu2Eb96zIbrlKZgcQja3SHxrwQegwlAmNZP+blLDf0cdASj
LSNpzcEwvyMi5Vp8eCTNU77GQ0itLBJ4FWF+vBX2OOp5YI8x7LEeN7EgxpgTpBk7
T782kcChP7HMN4Cku0jV7vN0YjDwc+x8AefuKMpIo3Iu2snSukZS6Te1Q+cT1qZk
INR5puUsSE+LN2LxwvVWFBmmL+f3Wo4qFqkfjpD/aiXTo84R11+1k6flTzW1AuuO
DOP3T75ZnBkrwp3s5b5TBRMZbnwNbZpYPd3XoQbiyNQcV2EQrX8jF0ObKEcpaSya
iHHu3fAh/NrDB5ENazybc+Wx2Bq6OM1Tg1MptBf8sK8RN3yuctY2lwEEjPpl50hp
qhQrENlo+4+5+akt1j1pCuByVCOfoQclYRWUL9SsOYhKB/WguzEmUFk3PEGOUsLr
raW3cgbhOxcOrV6bsboeNsNtHcA3QgFc03jG8LYyCWKyXHXzAy8ytSv5ToLnzNdy
XpXU2a6AGnbe8TFTt8mU6HnPXNoXP+ZVTML9OmU5y4nQ1q3MmWe+B8+pAsd7IU7j
t15onDu9OHEF2bF0ynJMz6FucV6G1w4wYixTlOGmACJfWnm4QyV1wiDtV963RU3+
SVnlvBASnPkschjaKnzBSwS+8tS/3fl6FLbn1cikVJBPYcNE8zVzPBGf07QVyEqy
ZyHen4t3j+1LNIXvMl209uGW3ExEcBzOwY8U7E6KT7mb6hcEog2MDx/fxucPke+8
mppkAwNEqFHTztQTeZ1416Q1UpKYFCI8QSNE8jXy9hZy4Ve2KfxcGdGmvdlzFUVQ
3EZX8vJuFwu1Pk5PJEkp7i7HwlBHIpq3aaJB5OkpeWAVNnpM68bImogc3ki0NW9s
NZfnK/ibpHr7wte6bWbPaPPa17ATGjd5z0pwi/qDexrFlbDpDtXLbeJ02Us9UdNk
s5rmYENC62vmHP8JKx9XS0ydBk0vx4KRyFDXPqyFHD6l2pzUP5BQFbkpHElD0Y2t
gDnbhSMmdPiREszL2LA7UBWktwWaPWvgZfYuH8xiCTm3od40DTx2TPNi7m0XbskH
ply+j8nWGPNwkUHLBDYeus1vuUkumsiUEvNg8DHyQWJpfagxmwt7ck6APNFaqBzU
lm+ZbqdTHLJ9idtDnplqEgsorFmM6H4u216A737hIUOhWxnbjDPNR5pwSudFtoRP
sb+zezat+3bI9GgmZmMhLEH4wMgvAsTbRyyficDT7rkUhY32Wub3/yRGSaS/rlLi
4yz+zWniJhEULVpLlSQJjMco4dA3oo5BtME3kE9U2HvBVuFj6DqrAPXSop+bZ+Xy
GKMw4nvkROCRrRur4MFxoQPjVYrWBDsdspTobSYHaMTkw8GdzDp6A/DUAbygZtRL
3To+k14xvqBCkczxp7dRmxqlX2UM6PrJ9m8ADf+8rJ6P/+NY8z4DfGDQz2hXShr5
+JkoUrRVFsNe96cl9WzlcVy9wGC53FJFGRh9fg9CWyqgHdkxIlJi+oP3ZNzAAlQr
4YZ3ws+m60cKGir5t8BoeNRTp4QdjfAziV2o4zd9XKyJ9R/LsTGmhSCmTxxqefRd
XheL2q8R6Ub58DEJkCPH8zGLhEkVJh7LgKPeoufnuMcchz/6FOrPAVDc0q0NMoEo
0Bv5+Cm0Q6bDZIYZX2PJ8fL04LxDOw3GoomC5GPqjBTTKzIw69ByoRmsByuwyrLl
Hhy8zVdDd9EbWl+n5SktVcLUH7u1AD8Wo0EKtMcsWa8t7uBNt59OwAR0lgOy9V1M
EUHFLtpaMR3Bson+tHkMQQl59eDsbGU69QKnzVh99E+SN/hM2hSrs60MiIZI25y5
4QtOpN3xo1cLl7zqAL13XWajOxomXMBZGRR1+BCmRUy22faGcLGFV8bxSs6xXgwm
TbHrhCLru22B3UguSlvhrxUvjY5uhjCWv6N08BLFxj7OuRXUN6ua5sjJ6vKq1p9R
oo96JWJOutGeZ474ozhQvUlbD2pmV+LzF06PgwNHiqxMQ+oWlwB1nwGkkMmQaXwl
ySbZuAfbPyiJY4DiYXtNorkbtSbYZavgjO4xJBpT4Q3TtTIicfKxo+BA42Im/pji
C3u8hqLweYK93QPI3MMI4Wd4iaN8KfvmzLtndAQoSQKZw9beWnzef/diJT0KdS8Z
qYtX/kobKS3VKKxxe0l+LzflesRmYj820ht6c0h0h+F6lDJ7E/rAvN0Zz0eRsCMH
UAhgyUwwhb192zS5BwwYOr/fC4ZabVxi9yzxgI1Qz3QXXU7HTeW5fLJtXtzm4k/M
1K/T/859u5temUgjZa97YNHfD/zz1Dtyvy3Um3OObLReDA4eSOgYAA/KQ0VZZzxk
LKyLEbqS5MUuR/D3Fe3Xed2AveCFYBuhor2VkcsfVjFVne1xP8ilcDqIJ/mCpeGI
mD74P+WZw7WlQgCuR64Tjv1FkSG6gF+yBWHUHzdgcsaRYIofYv4V/BYWADsK2uTY
4hsu7E1y5btKyu5nGbiVOmd5A8joUByCyPWbzSdWWOdMCsLpOGrl4J5QyFuDJuLi
gxnbJPAUQskSB3erx+ZGUyBVjy/H0gUaiIvZTW4yqQe0oXzF/1ARqSGERfmC8cNF
4GLJbvvPmy1leRvOTqGlCn1c5pemDfF9L9JfUpsdxKaQzuzJKvU4/qAtiwLdpJtk
mbzUziV9uo9CjlI7Q+Lkr3y5dblnqAUwaajTaxmtqMGtSINP99VM8wSygpKp6uT6
twxp0p/Rjd829ikPd7gkioAdabVa/tbfYzhKTMtNr4lIi1/hbGY7NejMVhy6r99N
ODLTSpndX9HznfQaAuokTVtBuT7Y6zBR8vUNKVVXvukK6ab0UmNubn1CI01VjIn6
nPmnA5Cs2E9LPZcyhf4wnPBOsCXq5My9MJ5MnGfiT7nrHRSy+z/UAjyW5zOOp7Go
6jIM1g1ak5hd+/3LTASvZn+oUmfPyOOD8XpxoJxMfkvdgGG+Pl2aKTwuaipPDUTg
29CFURv+CdtvZ8LcHZeKnRNg6l7iOo3z2qa8UjW4kzJft1BYXMgMSzOlZBf89OQT
v+3wh++5StTlIhecC8885pWIM1J2p9ffOmQXHDcSM7GclL12olWBnWry4kW72av+
3blciw2XZIgIsgE73imNZyWa8n9JSbzjx0RPRP8WmZEluIGViDQZq7a46N/GqMcn
QbZlRZ7U0KhCE0xC376yF4yMPsoTCLBpM/RCvvGI/xkExCl8zfKFCACrsrgV6JS9
h2GtJ14YsCh5ezlXfEtCxx9gcnO+R/w4YdYYZoJIII2JHQBoJ+Jn9lw0SD+kHBXz
XuL3/LVZ1uzJPtqle0LttmAfh7CFqZY77u7bRD04RYpqxWDUHwrT4ylFXOtKXi+f
cxUZlrbBjUIojGz841x8DdxSNO33QDYR1VN1lNny9OKKgqSpzb1onmAWb5LHAtW9
/TRcR8qn9N0KQ1fgwnRnbPQdLFUxx+16FtFL5ifbu9IK6ss7Fy2jg39GzbKRKMHn
q43gog6LiEgY+9Q8hcbrxAWMZhjj96cWGBoqGUHz6xfdQ5qtvGtn7gEpkesJ7NTz
kwBzH++BbfAOuBgG2roycWTXZz8R6FCkiI9NglPNYAetP882XmXMEfchaC71DX0t
ZZzz4kPTKzPjtYlA9huKnJ0COOzKTOeH0/Y/23ED8uSugN2L+DBwLgpSTbTILpyJ
hmd/QGSVC1WoE0Sl4/c1bwLEZrrXJdi54Z+UQM9RXblZ8u/M1hJgoICiAoOh5TX0
so3re8SSUQM97qMpp/+RvTDc0ezaS1u+5pSgxYm3HdL0JBMI9Zx46nlu+J5eeZN3
JVu5FoqfBX6oGexXF9BlNnedwIxl/GRWke9R6g9QcrxGIMaoBguJfyujQNpVd6o4
Os1gLQt5bkJkn4Rfi7MmV7qK1ekgT8tOZZBTJkOdbQeoa2W3UULQxXpgGjOejB+7
qVT8R8qP9I04FH/58uB2SpPc+I/J5gGqbwXqc1p0lXagwuFR0FjCRxu+8PtIQAos
vLxWUvrnI/STTiKvSD9MhdxBwYLoTnYhU8OvXjBE3YEvlVfinoWBozWNeH87sUFb
/YvCIpAf5KwDVkMSGLUIn4I9byjpJSMxJ7DceKciX9TmfU3+oL+DBy9fNskl0bOy
6a08ceDIqHnfQ6y8TyUwoLALvxZ8MBXTxGa574QSQaHhq/CAWgTejoDNnskxN7tn
QTt4dRq5iMkuhTPynbVhEfWxav2GWp8EK7OC8o+JA7PeVU8HYuccE1FN8B6PJAZh
fRfa6gY1HSnUTqTJc0/jflAiXWArl6hhMZQTX2XUA/gHOeDYOAJ6tuFYN+FHfIYC
ERvL0/nWqhRWnA6tCPtzCi6sYkT8Ou7XXebyr/0CQGu7Ca1rpj4Yeqe0L6vlfy2Q
7V6KCUpiY9clNod9h7rlPszxduaVS9PMi2aw3nDbeeHUWEkl21rhcMayFm68q3eD
vTunc+/az1YvgsAeoYiCmoEi4LvU5GoqOVm1tCdCZeNN8L4zMtsYFFUYwxSI1GcT
G0SysyC9DfYo8v7ecKCubHeij6KQfsTTFZPJQWNHGg/twelap4dlospCU7Ena5Rq
04OiOYczujzFZQ+VfFRxlmaxKA2jHApUIU020y4TVrRuCkA6+eZyUPIuW2pWJUH+
JvHZrLOjqEbiRMmwvsPtulHe9JExSwMbri6T0S/QIyd+0+NjLwAro2qGQvazTLZN
IPiTP3o7owKgl40pWYFsPb/11TT49qxLQ7C5lDX1uVvtUGGFs4UgS0w0dVd5ZASJ
NspenJ4ouU/pkb680Gq3mX3meoZZjBpTfo1nUlBj9EUqI5ZYvSeAeQfQ/AK9pfuy
WQkIQ/mJeNWsI+0KO6l0xSzg8LFRTRHsVxvKuUX262MD1jb/6yQSZfBVlUy+fxx+
hgGzhYLOiZhNS/klTgVi9pStcsJ/vQvRxurldPi2gASACCVfS1WLZlyAUacGyLdq
dTYc9Oq9DIuAA1IfQUS7KClRnwsspuv+hkX/yUHFxE2y2Uq3/XIPYRhwO7Zt7dkr
AtqIuVFKFTVAzCRei9zhAeH8blPofllyw/p3UR9slwtn9Iw1gJFFJQqgaTK8Xhvx
0cbJFnRR3QgKT+oDincR+n959G8kvj+yUiKV0naiQybr/lpGY3bqCn8U2PG9g3Mb
qg9iAHBeJIo3ZGCFgVX9WyLmI9DAUfB5AzpweDuzt/Y=
//pragma protect end_data_block
//pragma protect digest_block
GqNF0vA9Mb29er5nmBooVkGtEDI=
//pragma protect end_digest_block
//pragma protect end_protected
  
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PmeOa37QnasRpxodM2apqU4MtuOx3rq2bv1UUBMAcM+g3lB/ZqwKbYlTfmF4H81e
TFGfDtWZRLYgvTRx1MGVeN46pPl8UBxLr+kKwEjOBGi0I8EF06Xde5eITgnHzWDg
MrbZMI7OdT83KepgVdnHQXRRz1u+SfcQoCe2puIPTJ+G+zIDANqn0Q==
//pragma protect end_key_block
//pragma protect digest_block
7TrnDllYq7EAv/0TPqsTzhWrrIg=
//pragma protect end_digest_block
//pragma protect data_block
8nV4fSulnDvolkvQjVPzufIJazTttM48+8v8azABnFoFRBFiWY4VkuAdqX4LDiG/
4W6oxwQhwfYSjKEPRDJZwNMV34XWj2b70XT+IY8kFSf0/Qb1tDEkNJGjh4FIFPYe
2xTJkl266pHTTEBj3LmbsBzEdECQitG1Nxfhpue39E0Vs6x0Lx7BWUBtiYR1CRk2
1Z8i24X7m3VVFU/1JZc7KQwqY58wcfM3i0eDglUv36tsjy9pj0G1+SoCnM83tdVa
zxagRSEm2SlQ1edmmU6Jhg9LEkweQJFD/VMk7/o7YXVRqUM3hPYPdZ8qZqsl6Dm5
aditk9nvwniMHnIyEZ2OJvO1AkcjbsmikXvF+ztK/MLA+hvr+jT0tBR4xxm8q7ZA
HlocKZ+zvj1RplQSbCj2iovv1Ij7vazNit3paYOaqcs=
//pragma protect end_data_block
//pragma protect digest_block
57+lSwIdllYY++9uYZCo24ua4CY=
//pragma protect end_digest_block
//pragma protect end_protected
// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
mRvKHuFlJdrK3+O2Ud+eqks+Opkk5OaJbUahycVLW7TGeVSB7SsZKsmbSz8Ihxud
N7kf0i55EowcmFJIoYHZl6cb9m5EHQ7xaEJkezkeoT0xoGHWCNRN5maj753NJsKL
WLO8I9N1IKHXbyfaDIqQbW1y7rrpE5NA5FpO8n7PeVz5izNG1d6f0A==
//pragma protect end_key_block
//pragma protect digest_block
JD1k7dpf0ZDR474HvIIhTEh10J4=
//pragma protect end_digest_block
//pragma protect data_block
knPxZPacDwmaBAXlI4Hn/F8p2bUZj9S23M9zFwcWyrIhB+dWfev4FcgWrHJihiWY
0Pz5f1agYNAjel7onPpAL03g6vBPN37tFrKC9TJwdEqFmgX98RBmgwUPMlhO7iWL
3mM++dJPEDP73WIFeSdG4uEnbYgmLd5by10bnw9Sz1RHtoPfHh0HqEfhKSQ5eJRM
ZsNf2+3Ob7PI9l3azKFtf818Kbbxc+QTF4O+/1UGax/UW1meyXGzzrj6qA6eL2Rg
F/BZxA4w5ki1aOyPoCLtTCetuSQK1ERNZgNXOeFDiFSOpAxF9c0KhYXR3Mnn/Uqx
mVvC7a0Ix38Gh2iQekbNKQru+pSvkd+Kx2zm0AyZMr2WIMLxYLs7bjiKiexDW9Tx
c63l1k4POYJy1HRky1phZSDJ++jemgVfqqCCOnrE3EOB8Yl0KLWJRWKS3Jp8jPJk
i9447yla/mveiLlsVbuhvCjwjhY1N73N7HUfVOYrcyv33JeoVUPEAe3hTSkXoMA0
8kdfKmcODoKmTcXGXBg90E5RO5yGXLcIeB++YVWUJLU=
//pragma protect end_data_block
//pragma protect digest_block
j68UyzLvy9FBSJYKcZOO/sdsLVk=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
le25w6SgZ+HDEaum5o7/GWSRS+7AYIrCRVI/Tn0adzWnfpgEZRvZD36vw9vNp/jl
GeCNCNzOnpgYidf9FnIRsPxRBL+z8lwGUIAjjZbam6XesD/DO5SliAPdLDRYKsHD
1tK0joTQV/o7rT3cRzOpSrI1bCzS+eX0k8jWGw88LpvSagkgEvsLDw==
//pragma protect end_key_block
//pragma protect digest_block
wG7ww9n5TevyBP+5Fv1PhqHcTYc=
//pragma protect end_digest_block
//pragma protect data_block
gH1ntNC1voEFa565EPwXna5JKYBrrOMmcJ1C8qSM8WHsZdpCOlgDa5vGt7KLL0nD
yxcJbJnlSJcZZB6luyrSEH1Fs18cQXOGCP0yr+Y2yAIIb5GP0LcC3h8QLXiaqH02
OpuJHwsHnpqiMnRR3JP8paSf73KVp4oBkWwL7je9KVWj2lwe6YGAX2Y2xOuPkAxD
AAylJeKXLPTKthybczMiBQzvaFc0waP8aMW1mmI7nPwx0OIKOE23i8rLSAE3m02r
OK7fKT/yU63CZhqHL/BPr/Ur4z7+34sR3ZpRo1U/IBpTwIM7xGAnMnhHkr1IE4ke
0ObkisHKI6UqmW9TdxUD+KRqF+yV7AGloGSzDQhDdrJlgXNBH5RbzWBgxGhf0X2t
PSjUOVBbZqAlkVca1dAM3HTiyTrNFvt+lFRfyl7K1lcvrqXlu2B8OxfR/BfumaQN
3wnYPk089xswkrFciPKxTmuQWFBDKaPF2ChvaL1GDRH4w/JbJO3hqHOll1+Joop/

//pragma protect end_data_block
//pragma protect digest_block
46Oi1I2L6UhvRUfHVWQGgwYYbCg=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
VfPewn62JyDPKES1BjusJTReZe8oN/4F2im2EIhwvy4FN1AhPj8crSfNeW3+ynDc
+uQf0t3RfDS+/4i5LVi1DbY1LbhvABLE5Wpp6eHvyxkxjjPFqdupzE2jbQvJaR8w
uST3AgoZIzDCQLSTOqHd3lmPxOV/H1BCBGVpn/lwo9vIdhX9q4V+Sg==
//pragma protect end_key_block
//pragma protect digest_block
eQxFOy53aVFGZ+hxNsaolRcxYz0=
//pragma protect end_digest_block
//pragma protect data_block
dbjGr/wZhapnmW0EVwTRXCfz+F/qkZv/Eps0zkDTga97N5jbXUr+6+W7qVyTNa4f
2QrzYEujUmEhuhoNijSw37FUGUKY3T7oKa2B2uc08Gzzsw/vcCTMpoXDgJ1h+cco
FSi0Ng22yKpbVbncJk54vEAEESkaFkpLqB6RCh2ArEAnBmEoRNj2x3wKX43qw9ZU
T+FsW1E6EI4NmYzc/78X2lQ8e6IeelCkuKB67xEuX3D92cgGE2MbS0fwdOzFSbE5
dK5hhjvrCyLDbCueQkFTIdMj8v2h1g2F5OZxeQPKq5a8vEyN5JyjChfL6FHGy3Md
4S9i+6VY7jhvGZJoMP8UH/cgTiUgRoI5CHzp5wAT9SHc9W0n1j7I0O9POIJbDyW3
rKR9aooXvJ04KkibVUt5euzcnpT3hqqP7xdJjRIEiEkdRIbD3rs6v7hJFj2B3afN
P7fmbpyozW9GdMJ36MZNpV5ZQ3Lt99a5TSxSgxp1CzV/ytw4gsB651O4XvxAXVxj
Xgx6m0SsL6nd4UUCSAIBzA0rMMGEV4fK5AdzgO1irrTgPFTaG1Bbf4Wv40zUV6hf
2FuBKKji7O2hKcYvaJgmoZXYkY81FXup8E6msQoaubmRkPLIsd7itIKFd7NpKyMy
tVsURx0LTuyBmoV6ybkua9NUdmLxS5vqBuhaFWU+WTZlL7Rfu7WTNm4B/20RsDJI
b0p5IAPOkRvVbjlN7EkshMUE22BVxxUJqIYvGcjFXT4AiMPHOWYi00JAy1Ihjgk7
RhgdFd69ae1mBNvA65SRwJAyWwjfG8B0l0t5vV2YinHQZwBf7qtp5lybTp05GTYp
xCXiYiPs3CAJqh8UO233HjeTJ0dylZBIwmBNCKMf6/g+JEl+jVH+si9scnEbQo5f
8DtgCO6DPiaO324nnu/lbRYHWVQNHfNZxrkOXQJRkN+j/lXm/5vuMim40msZfFPR
nELj/7fpXZqKNsN6unF/pmFiGvM6KRcEAMTN/hJqDQg5UKtiNAobXQumv1RT9J/i
RkU/v6dyPahFJhdhgIt/IIcXVeWyenjm/ZjrRvYixZgmGc5I2lXQPRf4Nu51y+EW
QhVoULnO7fimhXcAX+hyGH1P2LFt7tMVwZjHhU6zPaU9My2FtgLVYT6IarQhl2eP
1EyBeMZl8Mm+S3Lr8hQmhXXLTGhRwByK8T32nsoL/Do9jDoeaohsWgyTgxovedmc
ycR2nFdUvpXpJd4MVe2CXSD6HqSTdq/r/OwvVySKLyTUNpiata0bJkYY3b12nj4z
5E86qO9VrQI9VVn7o2BMPSWlMI2otxH9H8HVxEALppq0v33vT3ufiKvguIxG1OX7
xVUm7yxJ5jSYVscf02kx1NCPOl4JX+LSaFgJAxrRiI7Jm4ubupf9PTBplUSWjsga
iDO3BK4Zeniq8EsFV/uly3gJzzeRcb0a7afYcDv3txljvq5CUurvzheqyVyBWbHX
mZSwnVHs3jmbbBSoamTLcVBTE2fio0+zYap3J30SozS4GzqOkDNtDT2KwBytBJU8
4piuGAxOODVq3NCgHrDURY1ajHx4snJRxm5vdaZNFct7buLZQopTIRIfROBxvmdn
p6j1YaOdGzd4jDdMKFUSso8iGNoLa0wOCdtSnL7x+QQIQxSzSyxvowypt5pARypp
Z674BF+kn6Mk35BRb15GoLWD4WKuf8KJ6ZDi2x3CqFVoWReQcznnEG6Y4Ixatt1u
XMvMk56vbU2wHPfkK0R1/xw0CmCdB+nw6IpocZJYOc+oleSh0NEzaUl2FSfCLIha
jftY4HOmQB+U3Q2fXlY4FRvCL8I7+Mi6ljn9a1FbmeOEg+xyR7cugyoodUrSkwOh
G5m3cuCZNt3NBTuwVb+JqeyiIzmkeyWFZx4e5+etoaaIvJV/6CkeDbznpqpUcdMW
lCPpZtsX3Vi+iREADJcY9Qr1XIcTiQvEqXzO59If+ArMkk07PuV/SeBNFFustOTN
prIwJgmmlOm536ydj242ysL6Uv9FZ9PypG8jTVxQii8Wv/cDroKn/PzxVxwtzBao
WP8d//P2SkLxqEamP+x/WAlCsM+kaxBYqDvB+0ONA6bJl6X6DJ9JkBarcNpXdLfu
56CwY0+aNB8Ttlgzl4hUr7v0S05rGK4w+YF7ic1mOdmWJcCrFhG53veBph06R9vj
7byRVKi0H00L/UN4+upmSI3HAFsjddWrW3yj9XpCGYmnKt/wURGq9EfIBfXPoE12
SQBA2WGwKb/RauuK2qWzPepb5GAsSEmKxN35ZjX/f4p9Ns1iQGCzHnyFPNVEMGE/
Vo3J9pAYnxGVcxxinY58LCl3AbpOFxuX0Fsuctk+Al3Q0hEnNZ5NYF+FgHbmRkNA
X4yAuyiQP4s8FhRNL63Ae0NiDWbZdK2fs4UnSKDc4TqIMmfhB26hh9H5CY2Df/iF
PTFZYJEAMlOoDccoWzz9XM5UOiNXN+rUh38Tgx1Xo+n5W6/LFvLEZ2cb4rvmd11O
2TnPX8XXGo1adQwrtmGXTrq3bPCwdLqShWDb8X/T2h0e8YOeNtLufO3RwWiT2H+t
he1cI7ND55nrDED4ytlDuiefRTh1bK7U7gCgVRl49qJAJ2ywbObRt8m5tpSrMxSQ
plLeNFQo3iJQHXZm9OULP6ene71/o377qnhKz1ooq1yc2JdI+up2dGi/kI9ZKCZ7
mrQrfMNlfr5yR7bvYTxC0Kc1i8cupH3A04/WPfxlexWGKRxu+4rlEisFZxMNgYcc
kuTpxVXkLyfzwE1IGyYPgaAEIhW7pbuBS+zRDds7Gl0H4Ea1C4bt9g4xV4JB9bdn
5Tf4WmUmdAQZzoovB7bUmQ6tUhQ05Ml/nDqnDmlS/3R8yxSJ/yruzlI0DiDqdnHX
bbDr0rxNI1GxrRybAyW8mz0AXObOFZpvLPLjqB23i71dZesGvSjUBUSVDrW86E+w
+3qM3a7cMbGE1EGjAonfCbeGSCbJ9yRoMJX2VXB+a1iZxRK82S9qXvoADm73VOZR
QkbKtakvHhQOX64tuDuC+tvv1IxxJVonJVkxtJkfPdXCCItsIWxOctlyGfEElVxb
yRvDjclf6DJkGug2v894P3b9Dk/P+EzODzFcAfy7sW7ws6pAOOiV1tp0qOOkBUeV
VS1uxSBlXC3YunDg7x6DtEycOvbOvapstAH/vmqC4MKtDulb2OBpvjw9YPGWNGPO
WEVdXKDWz3yByWLc6egFqNFl00fcSSzNwFOCM35NR+0xDKGM6DgojSn/ndk8H2VH
QKweaxKqIWSJFvY8jliI5FcLDA8qxKfb1B5CzqzKrbEy5w3Z9zdPa+yfRgMccBV3
33/s+tw8yz9Rvh+kTqCPcmEskQahq2BI6C84KWjdDfZKMU0BFTvBbjO26euuouXt
pgYx7MSTGcD4pT0BxeJf0f829C4zBT67a4tYcD/HO6fJyHIzFyICBEmOsRVyZ21S
nsrdRBRXs04JNsOlaRZ0Tfz+I7AJrwivz9Wx7+ZlKkOOeM7XeAEbhsiObERuDqfl
kjtRT9iwPwq3AXknIuRdXqrvlTUVRPGc2u68l7oxE5szVV5U5F6B6AbouLAofkQ+
KqfFgP/Ot2GGNSbO4zXI5STJiQkOLp0StHfc931UWyVtP0w7yZW3SUmKgKmYfgOF
4tvhcVQ18ZVsGwn92XIyB4QJlSfinOl/6kus2wrYeYtEwf1GU0bQtc40gTFIXCKa
8LY8utFcWsf+nZe6evurvpQvUcD66ErQ8SKjLxKQk0nniGTlWRYkJk1z6xOcKKn5
Ouh7dtqJpFg32MXzuP7lQGss6qLrrrfjT0lsj86MoSNGhxtA/kOAF4Js9o0KQAOp
ZqKY1N8kp6Hm1bJ8frMyc9SRtTvLRxCBrlHwioImZW62Ewrj62B8fyApCwhUsjsX
XrJH2wQ4CmCd9dh8qUnyRkF1ZTFDBO5A1e/eFb0zqifmE5Kt3NMTxrhaQ/FtSWbC
ZdXlTK3gXGxavkR4Mcpj9ZcZjdqSKA3jf959Vvh4aAxCMUQjn+W5VVCkt0BW92TC
aOTtUzJH845iluVNZi5ACf/sUFq/EvDUGVU1F699yRgb4+R61MFyT4DGCDCiBCUg
/2IO2nlT/Rgc6TfSMzYRqllrVQdW2WjjEq4Y/8exk4JT9p/OG+3fwX1QU0K2kMcK
0SwlUHcNa784CSPCpQ80kGfXfGl8nmFZWf7r5R2NXDBZMyZQdlzOqJ/cI2rRHTbn
+fuRiY9oinqkmPqCUU1e72vFIxX790tgSGw5583vToI95CXkuZ6sRyVg+Jq4icPz
FtZc1jUri5qRa+fU0fmRtwHxPGbmURm/FXS61vMmPStE8MxGttfreMs/TuQQaTOa
UCtWlacWJQrWrpcws6uF0JuK5epVOtuCQkX0PuYUuAIfx0fTFwkmW6Ot/rSl/kul
3aDAlWRwKVazUVGHJipo8b8JWNs8axOUr9cBu+sgT2SumtB6A/AHWV2Dae9hlaWb
KiGRazf+GGIuuE6Li7plBy05dOkC6Rv6/882cXPhBD3yxTnDitZIMeVVCF+B1cpR
IJQbimufRoPyT9Bu3FgJMxaxKGlZMx8XUqkhTDdNLtzg0+4yo+CqJNdd8KgluY7O
JDZUQ/G5WJEO+0loKNjlQslaZwEtGeOKQmSTJX/NP8ogBGPPn58+axDE2AWAG4ZQ
LQpkXs5KkicGBE04pSsnaWGw/Ao0E3xuQxWx5WqhUKBLrmcfD5mpnM7mc+ucKk9H
sVR52p4pPR4kS1ZNd/j6BdpM/Ya80a/pYC50bweCmCV/bf6R5P8ghy2NOqena2gz
ghAjkCn47oXcSl0MchTx1CcJZIfXjHmhDNaxvKRfwX2wTkxtra8rjYXJPdEBJitY
Btg86kTFom4yLk40RI/gLIyVawBOVGD/VWqu74KKVZxkXtkPQsjgj4Vah+krZCKJ
QNl+owGZrEFVrdMAM6pkS9cCvFkHXJCgMV0qhdg6AaQJjiyhuuIvJ8Ib1Fwrq5xq
bQYxIG5281RUnIYZ0Pu78m83TPbdkRolRcNoWQDHUKKER9zuzxEDkQ22U1ywk281
lQ7BFHGd3+gvIkr4nMGLZJf08SE4yqVzLAqGEQoM4BcXvl/Wct1BcDIAuTw1xsQp
3Kkd/8QzqUnC5L+hypfBOVODOi6AmXHcAKNw3MkQGp5x/y2u3vkyhLNQYjMo/TAA
ppdmRrFeGYkrdWjgQISsNdyG7h86BvHsGck8f1UvDPqDnwUYE5XN+Ez6LwmaeO1A
OlXOFI6Wi2TBmxGFRP9Z4aIt36oakzJ3yGGpbymAMuI+flLylqwafE6MJGpxcSnK
+w6KYt4vFzje+utdV3992PU/NeRf54ojr+F7rTtLOddAD5lCzwS51fsdoa64uWdj
k7VorMqgBKRWs+Hu60ZNCQoHXpaERtE9BTXitZGvH3PXvA0O1HPEAAw4Kz8BH2v0
lBmFtXEqNFPc6DanxJWLJfEd4aEq7GTfr3CqHaru8UmqjlH54cu1ABJovYbci+RO
WQ9Ra5UqRTCBCAV0+yBo7zijar3JeaWnt27hnnFY67qvoMnMyr6F6wqORjF8uAOL
fIemdaLqA/SY9lyHENc8/gqSz6xJPY9QqlIs9JBg7cKfAItw7GE6+3RDcEG90jYA

//pragma protect end_data_block
//pragma protect digest_block
Pe+HrOwoq2EsqeRi8fDmrvMbo7s=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
