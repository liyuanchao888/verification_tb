
`ifndef GUARD_SVT_AXI_LP_CHECKER_SV
`define GUARD_SVT_AXI_LP_CHECKER_SV
/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */

`ifndef SVT_VMM_TECHNOLOGY
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Dzo58XvL3H2Wvu74p+MNzZwmKM4/AfvjRKO6wUvGME0h1huzqM9S7DwkMx0LOquw
oeLoiVakbfbuNDyST0ub6M6ILs6oqbzm+myc/QfL8iciX7IBxSTaxQPkjHhUsCDw
RLiAU64qmGCPj15v6Rje6wZZFzC60YauFM4VOEgikZU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2377      )
w+9pYWdt8Td+FNQzSk3CedVpAsceiI+OhQdMxYhhKFTofCX5cYCqiA6qCMcEAL6X
vSqnEJLO6NQ2jkATNpKcUQX4fg/Fpg+jv9YgUOJSo6IHt82eEjOA0D5rR4Ii4fhF
Iv7T2zwV27MX/ctlouCkqw47YNoTEqfs1CGOkV9aHaqc1a1wYu0u/96W4obO9ze7
Ll/qHXu4PRSfiA8UuiIQxncSBguICQmMynvRC1HsCyvFqTYZzwnOSzBk8Q76Kn7M
S9PvYbk+VtDWpxqql20IzVeICxGjmrX2k2IU8sC0pHaKLsltcot1nBrcluqJRRLJ
TEdHPNCCf1BlTje5SsB9cfNC1MNz4+J3vxDUkoRhiHv2fmF2w+XGwhrMA8XskPPL
97/zecD4GbAG6iYqgPddMwcMz1txfolNfAXiyUcuMyWt4PctIUJfpg7Gm3aDeAdc
oH4GO4Wiq4TpeyNh/Ex+AInibeMz8ijjbZmy0wL0WEhYGDPNQbaMyOhZtDAMHMQt
6C9qAD7I+X9K4n9JGHNxLDIyEKyc/ZoLtAGO3D8ik1TyzRJPXmPY49O+xBW7KAwq
sXhkxGEwRMsIYipRgXvULO3uUcyE4csVHxcAQoiF/aozkDQhnu5imii3/lhKR6n5
rlU2DZF6No4XwI61rQEYWFGvUK6TKqzvH9sYEu0Qojtw9MQRQw0YohGrX5/zdjfI
h+jxcCoJ869Yv4zdekJ7JF0GTw/5ZsBKjmZEsI4Lb0X2Tuvjf2GTfNggb4ZsQS3u
1kMBVLhYgq7JN3LWxYkXCecIaAPPL1wAA0QKQobmxEgh70i1gEcO00eX/4fLNZ8M
HEjl0VmDLuLtIZNo1sZF+XJHe2Xmt29dhakCTSVG7VtPusrO9gyne6pk23ll/XoZ
DsSdOgZlk4KlpEd+FYieQKkmVXHv67HhezV7j4Yd9cfaXB30dwdz+q804GBRPvCg
7/IOg2uzPyjl+qe6ppEBGIzok6FOGegjEFiyIhSycGH6W16Xbfr+ATBDb5ITjjAh
kci9lluEJGOdkmvH8sUeiNfNuS8n8ALtgFQk8XDBGmq0IiSeicggzKC/cb++zd7D
saugDV78jI4zibMimqPgXMdKoNa0gKFyWPUJjZAWwRGSXcFbKzGLx8xTLICxLeyw
TbYEOkcyRiMy8L/gl/Ve9zzcAHwbPKlPsWjwbF9QMxaMmT+ixV9u/8B2GU14TFyS
HN5fN+AdnBFp7MdTGU2ZaDQOZt3N6jWCYjzPc86sQbzkizePBUb/i5ngSDnDW8DB
NshxgcBlbhUUY75ZlGsU8GNHUPXWr/Kj+QD56SsvhJfvRB4sEIvGanWad59/xwFi
K6JCQhWIl1H/PltI/zRPq8Q8SbbwXE8tHCTkDFfKlGOXappbr/ecV2Z9VIRGyVfM
+QVE1oq+zezoujIioEmkFMfzjXAkP3PG1X4MevIcavh1R2xd91YJzSmb0QK77/0s
xJ3i3b4vgHo2TZEu0GDHaqLmUmXCseY7PoEuYUDhIBkdJ7chXvRyx2fAKYYxAP47
b3jmizUg7jYJUI4gspJ2lJPYUzcgThtyo9LycCQqBEH7v0v8xdpCN9PnARa1paSd
3QRE7JRvA3X61LS96PlE+Ig8pxInsee78c1ZJLbwZxBTcpNOIYajA8iKHB4fXcZa
YpGYe8HQUgQ9PrY/jCnZSwb79dxursooIfNg5FdZGnXV9Ui74MxmS/0ZNy37fA7m
JW+i6Y6xo8gTG/1tv+RfSBpLSKW4rdncLIXAMFKmnZ20okSbuiHxQwg5EAfl/3wV
4q24A6rkgCt6O19mgxwi3GSM5QGX9jkdzw2Kgkzf9zsPnxDN4uiRq5Pqok7YP/v3
7QJx6iOoeckymZycreu1Dp6sL2pz8GSAf/oPgg9GT5fufjdNy36IXFzl0Kzoncod
rw8n5DdFH3Qih9RLXGe6IxPdo83SqzFlM92m2hp48WPt6azMIHZqb/oGUMeJ9SiZ
uqB/J3oDEKNNWeuXrwluoxjLuzhRawN+Z4M6lXPBC/7KFekgVKBTagLRZzdK6Vpn
XBtfRM1mFJjsVe0aU0diSAi3PPDVWx8yRW75rMGNoFxxSVv7Qg+tUlWAjeB91991
DFtWl36CaG6uKnFcP2iSeYSaiEuQIXAfaVI9ESve+x8ZPjNg0i2ypK1PPMCJtkHY
jbUB4JGs6yM/pNMUkN+ReSBauu26k/WTuYHdPjx0VMFNbfRt4jSYno/cmQfWx7We
caUMDFCFnwC2NHHM+okbM+bKnI0c/pHtXYg8MnVjLQSxwYAYTXKsogAaZ/1ZGx8x
9KhsclQoKB2ozgccY5WA2P0F/DuCZv1u0OdMD/6sX3GsFBcp1+8Sh5zYZVygbUF0
652cM6YhNuYsZ0EXOcSPl9b06XS2XPuiPzw0zbVskB5CTsJbUNL9rxy1ow49PuzE
80X0WIo9wtNwZCmi59YTxtC7dbc6MkyM0FrdvAfpJaMoH8cWhybiyTeeD8j54oae
8GN1aJO8yg6x4GRK35iY/AQ72Q7l/+MUkzqmLE08HKA9CoD2TcGP2r2gkjqziywy
huavAcpnCuoCHnAYKOJ/0Zvq5bpbFeV9yNlSVF6dfcaEkxyi/yp8xD9Y9LicyPta
J6+iFlF36FDd70ChZkLof0JMk/HVm7FDRGc00vfrqh4Qssi/OT40bUGvu8nuqgTG
MsfQRv7kxQ4h4LAA0XUMc8q4uHmYX1RTCrJZLZqtmvXI/uU1ZnJAZ3j5Onw+wT40
wMEaeCMnlKC+h3p//AecM5cdj2f7EZfOPyAVUZJh3mPszaRWsCt0t8URbLK5Q6yC
K1zhDLtrnHC/nSGTap9PYcjIDowfxqtlm+L/K6bA7IAG6Ly0OUNQMEQMussShqqf
xktp94DhfewPsrReS/ZIQybF5QvC6203/Wh8jOTZV86uw76TaPfk4MgoXpK10OUD
2+JESNjWl34zRzkRRt8GjKbql/2WK7NSvTMHfrjlOvf/jYdFGYLNv/auIfTVkhbQ
IJb8d3DwPL1whYW8k+vhtCO0YxdMEnLn+aK3trF7OaYJ3aVrPtyGYMiMIE444ZaQ
b8OAzexEHR00VcBr/8Na0HwHFHOyeb+V+VsJ/FPPvw9waYFlalBYryTXXgNKqX+L
aS2IiJptGVEpUw63PPWSUftsDO61RF/hSOFuVYmYQ08=
`pragma protect end_protected
`endif

class svt_axi_lp_checker extends svt_err_check;
  local svt_axi_lp_port_configuration cfg;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AFa86nx4Aprn2KZK3lnOvc0YQOSFYJPffc/kb2pOeY/0+Deh+HQMnpJkwrz5XX4L
F4hy02pSfFgaERioCgbRHfnXtq/cZ6McOErJc7uv2sP76LxzvClPMMZcJhVXa6M1
jqQIrFDKeNN29qROLDsQVkVeVUlsGuxfe+HwTVTJ9nk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2500      )
+kVzFdUl4FKlg9S8FH4y0LGgieCgPVbGbpm6qjf9BSZxPqTzCdU5fjovlC16MWi/
NdJpvo55rp9b+xMGwoWXUvIC1r8rg8lQvSesRaaXJw3kRYn2culLQ7sZ18S5dvsT
GPfisfFBjjm1Bh0dhZcwUJBsP7n/cKoHWaXuLxI9FWc=
`pragma protect end_protected
  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";

  //--------------------------------------------------------------
  /** X/Z on the cactive signal */ 
  svt_err_check_stats signal_valid_cactive_check; 

  
  /** X/Z on the csysreq signal */ 
  svt_err_check_stats signal_valid_csysreq_check; 

  
  /** X/Z on the csysack signal */ 
  svt_err_check_stats signal_valid_csysack_check; 

  
  /** while entering into low power state, csysreq has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysreq_before_cactive_check; 

  
  /** while entering into low power state, csysack has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_cactive_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone low, timedout waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_timeout_after_cactive_check; 

  
  /** after cactive has gone low, csysack has gone low before csysreq going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_csysreq_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq and csysack to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after csysreq has gone low, timedout waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysack_timeout_after_csysreq_check; 

  
  /** csysreq has gone high without waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysack has gone high before cactive/csysreq going high */ 
  svt_err_check_stats exit_from_lp_csysack_before_cactive_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone high, timedout waiting for csysreq to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysack has gone high before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_before_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysreq has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_cactive_check; 

  
  /** after csysreq has gone high, timedout waiting for cactive to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysack has gone high before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_before_cactive_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_csysack_check; 

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, uvm_report_object reporter, bit register_enable=1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, ovm_report_object reporter, bit register_enable=1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, vmm_log log = null, bit register_enable=1);
`endif

  /** @cond PRIVATE */
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  /** @endcond */
endclass

//----------------------------------------------------------------
/**
AXI low power port monitor check description
*/

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RXQ2nwzD5OP2FxaVA/JcUmlkBP7NnZxtelk51nLihW55KNeqIK3jIne6MmkFuXvc
IN/SozlxID7Rav4xB2Oo+QUt0TdeMI3U1CUIq0/4m8YUjfA2O1ZR6U7+bVywUipg
XloAXtWV6HgL9YD3UTxToc7EprjPElP0OFYs/3924a4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4040      )
strPOJDguqSwwrUAvElmW/Jb1wXpjDtRGaGtDuzYTilYblwPYAUEnilKJ4VJ4cmr
OBF44tNIY/hCqLgd3PQWJG+AewehavErf6HNfEg+boNIzymgMgw8c2zooVYReekc
C5yqHagdJyponTKxsOEmSJ1qoFM455Zgw5y4MsfyekVX5kWu/ftf4XZ80nlgr9eP
2m8Bk4m/mK5sLfnnvojWrwXZdTzu2Qsn/S7fN85jmIsjvM0qCcwvjk/7L/xy3XWn
xz6KwsXk/cRwGjh6jwt6I6cKiHY6/pPpyM6bqB0/a3VWZbvsHMaZHz3VdloYNkPH
Za8dbT0+AAQGvguBwvAzlZluZfnandJThln3xd+2PJEiQvOEbYaR8BAKsBDIEbZ5
3ia1U3LgMlws0RdJpGmzsXdgmvTZ0lfuOieN9/juaDFy2YKKKyKSCBFGqaNSMc3v
D/XOQdM8bknxmHGqGh4v7WT0AGjOgZ+K63w+Jx2JOskuE0i5J/YJ0jdrccVUUMCH
KjgZd5lP2ShVp9c+ATcM38DZhjW5VngiDKgYrB+5mkgpZ0Toiv+f9roYJ0+axZ7E
R1UBFl15vqdu3lVGfkivy8RpdR6pSgIDYztsysXQuG62MV515KscVc79m8BGBmEL
ZN8ERMrgPbXfw0nyykDRQ7M0KHfQePTJOas+RzM3rF2ANNrzVatEbsx4W9jbmPpf
4Qt7RUahd4QxwrQIUmhpr/zrD8jNDhJpEng9ZhGy/pr8BrBDffy7nyQQRq0fBmVo
Hlgtjrx4ce2j8qJw6fj5imUXrs/WE1f2NjRZew3kyc8RlnZXpP0sU5LLpw2lnOp1
kwcujLi6d1S3vji0VYX+ZF+Wbq/LH1Uw+Qnp5HsXD7HkpdfYaZ02lhUfdDHT8M1L
hSWM+nYXDyH3lF/62OfTPP4byhVNuKtVjFmr29HsNPjlkTLD7I/fjrTsyb6YywdA
rLOO9V3g8XHAf/7nne7JkSGtTTEvsWbpm9ZHDG2WaNU3SACYRnTPclPhUaTI6a/1
dyChi0Yvf5uts2v3kdWuhnWWD9rPCWlwBYidsAmbyCyyGvEWts6e+TTfgXg5JTUa
m8NMRexe6VrkNEDBqqF/yIaLxpq2xZCkAKRqx6sxfBBbQUZ4QeYT0Up9sDfMkxPo
5dA//vkaZRpEdaXVTfSTxKkP4FhbkdXx+pzTb5O+jSGElWcK8FX7mLXhM7fKxEjJ
kwICZ8hTqKH2d5XMjl4ds0P9AIuHP0dk++gJPtxZggSNf4LRKVbb2VRO7xRLxxdu
0qK7w0ns7SRmn6xEwookPl5NIRHsnByE46qlsJoleVBP9IuLRxJFKsMdUfvDFJFe
3UsqMIK6Rl3E6Chk5xkYawSGtKX6xnCvNth8VGaJk1J4wUJLJWA7Q23r0kDxXqeb
Jqg7U0hAYrF+Q8rzw7xWrktNDNG33OOieock+r4hUvVawlduPlO4JAJHRsnnMCcJ
YRkam1ivK9Xrb0k9GvXa1JnXPb4XfzEBSnMQOmWMcFub+ipnP2AWrKDUf5xoENN9
Z86VBukktgLOmc15xL2Y6/15XJZqOywuFWHL+5Rk7BdD7lDugzATSRG80ElehO89
7+ukLrLiYtG8NMVaGbLv8gGjE7GtUS8G4d6LunPxt58xwvbCcp54jUdT4PwZkXk7
Vw1zJlOLOGOMLRS0gEXNWKcePEu9PBnM2XQj+X1Me+hFUl/Zhll6wl0se+LypxLu
rGoPgniSHSta8ATzPfZRGhxs16tCOS5vkX8Vlc1OLTbJvkTGVr3qYZTdE4nVoYFT
0OTKrRqQnZxpCnoGhdUyNzJrh8KytrCKO+t3SuZvswxBqkQIPQ4gIXBRoHBsWAUn
EcXSPvMnIGVx+ukGi6e1VDPqWO2KxI442JkPiiz3ndROZ03MROlijxfEB9bTL3OQ
PpjI+jbfplnqU8IFoKR0dfjLVBq2duBGMGI8FE0SaP0a2JVNqhHYhK7A5bxBSRuC
Et+e5H+GKdhhAQVJPLq0FrCLf3X+hsokAL/8s7pf+u9HCdRl+LSfxz1+ytMSVoyl
9VbL5KdJby90rTCkWP+ETg==
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SWGOj8oqWfwmgTR4QVT8wsTaSQobUqpd7T93BaLH72ID1qah6ngoWOvSDO5a0bf9
1B41Jp4GrIvG/vMfdxlZhpx48OBKvQomDeOj56h4gjrGQJo+VsuNmAWE1uEYlgeo
fypMmJpjZxs1u/3YkwIzIbja6wxNO600uLnBqMnn5HI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9883      )
V5z2giQF9bLyVeSv+CAENncxXVBXlS68+ke3aB669hmFUJ0h5+nptbreyNsEuBga
70szijl15nw+rG//Hq3df/rDldAFYGqbTxVgcWfXPIyrNbu5yIrx9rHxR4spV4my
PYDIFXFwvUCPxeR5uk+W42f37lDWend/+cYm5OLUzZ+6iWZTKOni1JzgkYTpQVcF
YxPtMF5+/2xXl454cZQNTZI4jkNYKpLYMm6otdGWmiOGtiBNigJ1KSDownUqvVTJ
j22dX3NJrRKAXzsG3FltliJWg2wvJz/hGVrUUM2Jfsc36OIxVGphlCq4wWT2VdZa
B2DfnGWXQJT1ywnw1NS2gej9lsVucXKjLCpnOcfy7FYVdRJZxbdFtgiCrTnk4krG
uYrgFtsf/Wy3uWh85ZGGNCCfT9hU6WnESn/yj0Z/feUAu90mQR40P/pn0EHz53JF
RdPnXphVhEAILhvgfEPZhsoUu3JejhYkGKrAg5QWPGr/+8f6OeIglb7ehm6ZTqL8
r1VwpUbM1bSlaVs/ZxqeqS8kLkjjMeshnrqCimeaSM9sbEAz80HM2ObgDtDLVQBB
PxduHCr7H7hOmFgrF3+bwUZXF9CXjRFarXezrq23DgZaHd8odZtUJtq9QNngKyrZ
CFCuakd1JI5p61oKuHBO0SYd4OLQGVRru3jg7FNoeuAs17qQ/2Ld2vbMai03RhLC
Yiko951RPgA03s8gIASJzGPVe2sKue+gtboW3UyX8UYEHpIJ6/VJkB98YFIWOAr4
8aB4UkythjEVYxOvZ17BBX+P2Ha64Mc3ItgHKx7oqKg5MhMvKRVc7X422IsXb9Op
id4yc0K7ttffTU9uCxAzy+UWvU8bT8lJvYdUWT4pNI/3WLqVcHetfR8Xw2zWDZAT
KpZGE37sqjRkURtWNeZH2GiXWRpMXPPTzSiWO1H3Tiqp4chiRcPn1qJcPUXk2wB6
6ascjGfDyc/WXnwCY4jsGnWYLkoJ6cGsl064MABwai2rOospvYUCbyFSuFoaM8oP
SRk5ksHe4PaiQ0fovvNqseVJQUTlmTL1yhYQWq4dvyhosT1byNohSY/8hrjqdKfp
FXtYjRGyo1Xmr3gzrwKXeVhyl1hduheNbPLcUL+TEV7wNCa2Z++0fthCJVaIVpGT
beXVDJW/M7G848NAFWKUW00JVEAiPvIiwTrK4aXnviee4GIz5qBiKFf+3Ww7XjRj
jlAKJAIWH7gwebvg76bi/i+4fTMzqJ1wChZofOcy6kq4rrI7df4+aQyuSWK6dqUv
P/LYLmGAKbvjtim8ogdM42oPdDTlTjRTlJRFph2P85JNUkR4MkAuGxQHFcaOt/8E
2zslGpo2Lt8FoRroziWIHJLJvPCGgPLan6vsKfoIgiQwXnoCgIPi6Uzs1vhvnnCc
U44T2dqxrSLHRQ6Nd74+K0nOyPe4rmpBpoHZe3EdikkjWyear5VDfSEdJ/6Bl9j8
O5WGRsAdsGKFnxcYSCS4Z/jb3Ps0SMT14cc2gbbO5/wXduuChJy0n0sXmyWdnIoi
b2C7pDcKzjjLvpWXWNnyyLVMszVCHh3AjSmFuV2lqnxcGiVoNHA0Xt3jA4EegLAw
n6aOX+sROUXuJzuvAyVqRFfbqVi0xp0NB5/GDQkFi3ahG83eou+dTZFSnrLhynnh
7Zgl4P9I7P6BIXE/3QMI3cS6sLew+qlNUZ1DPIYY7MvHM21+z6KjkDmA653qqtDv
T2w9kIIsHW3J/0JgGEiv5SP8Q0KKYeqPzVAQ0yfGOHEEG8tCFC+Q3uolnCyha6zN
oF1rG/RH1wuQmsSz3jAFCk1gzinCahuURKcZ2Xw2nW/BaChd6APTTrXE3xYl8T7D
4WDFsxuhZTWyJMgHUmY+3vjqMnGiKo9DgbjAcHBsF/Vowu96vyKczTtHolXN6DZu
9OjNOPfoT2rkr7xR0g67GnncL41pIVN3uA6pKWBxSHofnlFjLIBL0IyvUdw8h+xQ
QeefPiVR3iAmHZvTTF848QmtkGqfd/O6uPn7qyUJJptY/VeAhNszADRf8A55hjlX
90kcEILzSoADDakSrNMRA6KhJ15W+/4xj5EHIKBUtZJxyfwcAWOF9DJPRXni7tnJ
JrpeiTLUVk7RyR1rfzwA5BZGLfNZyJGDZe48x3U74LxWGMibhqJ9VAHtYBumYJUX
a0yrqqZ9KSWCKMSZdFL+oIgWNbjSY3VOPr2X0F4/6I4VcALRylOvaJtzTHrDJto6
BMrVcbrIMNNCKnp/agHH28WPNbdBUs3K5940b8mVtzRF8EPLTwT515SDh8QK9dBD
tUg4NDEuylBbhMPSILvkhIhwPc552Rnen/ov82e1t6u9iHQC2zSaFDR2QwAOlnMw
3225ufdMmf8VDpB+b74XbfYjY+WMkkiXfQbIuBKTdCrbHCX10f7/+Z5+ncvbaCAE
UGGk1Lfw1SMfbTNysycv/tvMv9jWeBmIjdb7/mOTk1LGTLzoQHuc3vqe0STVwgRK
OWs637xZAcP+EBlnlRdVJuKdjnkDgf2JQBwQ34f1S8eQ3c7JNyE75eqE4n4bK2Zo
d2tcotl9C3Cz+kCFyZADSqoYqz4i/Dmc50HSrDcxiIO5vGtARtce1oPTiLURiaH/
Tyst0nZ07BVAFoEasXnJzxegsJcPhDB0Jubl0FckHZP+SbpD39JPNwPL6PzqUcoI
sak6bgNeyzsgx+v+Q4WDXw3vcmEPyr2Wikr+X4emwlpPlzuz1wlLBOui3F0JSNDE
eszouYoxCVEoU53PHCDPYM2uPS+i5l754rQB6FLk0U9ZqM70Inx6u6p1DJ0D9vCo
xqz5SvKzGpJrZD4QNhVVu5pBWYDqkHW3m/elAqmF1LfMtHUVoMbDXU8YEOACDq3v
IHry6mGY7OA4A02NN6jsZOIMyE9nzxuBvut6Z4FL4CqdvMQVnKd+JTD/Id64/ClV
VVQ2Tp2/gbwWYy9ALSXHpC286YAlrLQI39nUkPuue5E0KBY4Cva3BBSb6/eiHoja
F7K+a4BZxmCjlh5ZzoJNCAO6tld4c738QP1Vk7tPQmieYFNmoD7Wc68LSEHLm+Hd
IhdRRcNAhr/pzmDooLyqc0BCbMToNIPyG++mFWMkUsEI25dNwueuhHeFkHBNuOWn
kD+0qnlHr1HY9j/dVgs61cCoI1JDsCPKt3Rg2SMFhxAjkkE6/lL1NF0CrVrzC0W/
AM4fqUqRpRI0gJHhCyYOgBI4aMldLgmwIMFM3c2MY5BflUhg1d3s558JqxPajMZ5
XF+BdiM1K5FyNepOShmMtpQUXSmAetd8oYPjl9/nocYJqv7gveOwRB0YvlfDMuCm
gs4y+TBGEvVZYRbpMB4ZLs1z0zBULVjGnlxLEX6KaLTDtCf+13EdbAtGBmNEaOMT
8wdrxWipknpe5FWELCuD/j47pUqwMB1y82ssDdmYhFakAUnOVR4KldzVG/nANM2x
AKukdL7ybUc8EV7SiibUe8mt15LQJd9IU1A6X0MOYTGutoGewGUPtjqHePBOf3cu
EH28e1rFjMB1KsFWWTwr9UW98XMxqvage0gblZP3rhNwtHe23vlkwlIXdbSG/J4/
cWl3e/k6IiNEcReFi92bli5DuAlbMAGLb5dpo2q5vVfIZX1sKA3YpjWWE+uUZh6C
nuuNBUm0Py38tH97eLmJn3d4Gvo9onbo3GUkKywu/2zN8zuBiOlIB03k229viADc
F67zp7wifxXXVGdAOnrxe24XAsirtYz+9uiKSEam6Q65DXpxscyM8J6eY67O+VWU
0jMbzfE8eZ2oL/XrpOE8WSWRV09HHA+eM3Wqs0DLjFy/JehGb7efNjv+V7AlnO8z
/ehdsfq9Smi4tj8CvUlHo+g++ahEiK4rKzFh9wPp3pD8lC1PKq9MwUGCyiQm5zaa
NzY206jogqbE0mZHDZdO6wJzPe2157LcMsjJTNEkhV6habgHcD9Z0TQwSTD3JXo3
471WP2aUdyO7wY9H4Jd/b8mZU5jEVEdzPZhkGf5RO+Vw+dhgoidWuBe47dtPdqYS
pNU67P1Js0krcFqxg9Jj+yAHKw1SqHC13Xs6JiAazb9ZwKBlTFY/yxf3Rzpbkw59
X5Zjf2XBrQuup4hrTioIJsVtttbTRcdMXnJiIqAd17w+opZVAN04sSTNBX2UpFD6
JtuUoEU4S64D2AyrLQl6bzUe703u4VHtq6YRSnOeG1iDcYoHlipK5noMjVNJ1RAH
8Jekm7SF0wScuEQucM1FQJfO8c6SML+vyk+VOh8tqHo2bvKk/VKB9AdQwCRAvduO
UJSpwVYsCgbxjYAx6hH4UUqZauSeWsfC4cNUVP8Lw/XRjhBK050d6mymvAb0pV5n
fEy/xtUhP6p4Lg5qkPQSMNSICY6FcO4qUwaausVUH+hAK5YhrH2HRxyud3ApVmxI
xdM2zm3EPJ4KXInWHxkDD+Ej4XPA7vMpytLEHgEHUovqfZy/dYU/Nt5mXJQuiQfb
LDMR3JNFOKhgZn0ZRVQ4MdweKbv6zMJY81Fy9xvUsSx3zf3bCQoCwzEBtPJXtL30
6K4CPef7d4MOk2IArHShSPI0yAiRKrCtmyZo3Bx3qo/dGQYKclqKd5MLU9C2f5tH
VsKsGZdS4wr7wJuk2MAPS19R0bDfH4BVZDZzct1KotTnA2JNhCm6CKqkmpqPkuTU
sZCmz1JuidgmW9zKs9zUxOzm0F1sTOA1yX+u+cWN89pUWbRInl4hDv4oNzrHOP6n
pyZSGMu1Gp0OaaN1FNfnnvoq62vLkfqLcDLUIUtgWEb0gN1++WPImNAoWZGxPa2H
/fwdO0DlBpR6kGlSUHN0f0+2fPCvRbh8o++mqz0gDypU/dFE6Gq8gv663cxecIWB
Bt3Ns4YU0kluPaFdGGP1hiqs5UPy00GHkLnvQKL9u+M2+hVYpDepHv8vedOpnlHf
d3li6Q5ZtlRBYlIa87z5zCX9Yly3aKzyzYL24QsfPJIthL8hEZaKW/4fYvWR3KY1
OWwCWO5Z304MuoabTEcThmm5+ZfPMg9dOWfYwaexlkAoJb0f80aCFm9lFtU2xTQX
8+WCEivpqS9HVu7Xlgmnl6I42YV5pWzfzNIzH7/HxjC25pJR0kboy3UOpc/hyRej
4vezODVMDTMHtanGRCJ+iUKm0vARI6NJK87jQ/YFmwqlUd6YN3nsG8IrUoylygRq
iW1E8z7boO7V6zoZnO7SfidCsT+BWOLqgFM7+tzO7wylR5drihId0MXHjR39X+aF
Tdy8hUNMPa7VD03/7bdz2rfqbxPRdAyFev4Mebi2Z5HA5ssPIL5aj7d8Fv1sPU0q
Y4bI64O6RfxBjUngPtLE26UVKau2gWPy82FkDUyEshgi0iMTVZvRlSRJv+950VO9
vD/LXZyCx5w5Kq3QWWwaGQa1d6ZYGTjanvfbGNn4e/5/rmyZd16JlC11nitaFyTS
dKH5IPMbg5M2wopnlHHJ8VmsbN8a+jLcmAHjr7RzWbjWVrHZ3KfBN9kQZDiwRuaT
5zjjnQ3+L77ql5LWykeZ8o4CDqM/MtZc8z7gLoTHO0YS257IVW1/zmiPqlLpBlRJ
iHeWq4YyuiF6nZygQyifz1tMB8g5uGAHyEzK9I5DlDXXagQ6WwCw0QF1Qww7AUFH
flkMVtHWlswLa5wWa/298p75K2PM36xGmdefz3kM3Ov2+cv82m38N/02UuMFYd5J
xwHOq8cFgKOLv+iQRCmuwqTAA88NL3TMVWvYYysuZxEu3evUqjrTS0GhZXSjEHIT
NqscCxwtAkM1fdPViENO6vfouzk7DVf+6bqT9pzya/80i7ZiiMt1LSfkLfUch7am
TavNxvSosGsmPqWWr+7Mc/QvbwQxSGM4qnZ2geT57jMRBeq+ezmi8t1Uw8bZj2VG
PX/iEqodlLGr4ljWK4NP0Y4obzC8DF6l7wuimpdC55UQc+a+JWYPenqFRGGvH8Zn
QULhaIf3nkFme2m51y85KmRL81l03qnTM0Uws34Iv1xBKgQvKxc1V4cs6SEFrSWJ
zsVZ2E9EyHy9qLWzCoH1MUuHk1RQUpWYGcNlxewWXMOJc3gusq/xj9Wg+otRr2KM
J4hC9B1DyiFNcbgjduywQg6mwJguftMr1vHoiEP7ZMZ76VZ78psMiwygKz0UVnKY
j+EO5CKqLeS6pl0T+b48IJ5/OWgZ2k+HjpTE9jqdsvSCNxTpLgI7sFnGIte6ypDc
6pTE/L2ddWWdY877zVUnm2EdNqZfAI/JWQ3NWB0aj+4hOpORXW3O/GndrB4Uengg
bH7K0u+fQYHOOuZe7jfTInNIIciW9igYvOfF481sOqyoAnS3enYlZp6JN8DZfXZh
K8n6OSzt7SxgijVXcEg4Ukalb/QbJkJIJ9azkwFZ+hdrlLg2in6T1ZXFSGK3aUEI
M+2P4nqLNBsyDWP1ULPNUmwOyV50WUdriiDCzedtP+zY6v1phd9RYn109rN4POBj
qPwsNQ/VHxEy5AUvG/MyjtvQKzYDdfez3npq8ohIQW3Cat0KsyJd7ZPdKyO6l7pu
ktDQzRs6xgtmPFdjZXq0dstazZhZeLZ3DxgBFpSLk4XSf4gWvZlC7kohnFmqhSLq
TUa7ZV/TulUbx1Btqvbv9VtjF/LVBFLTh7da2HGvkQC6zs20RiELEVRiJNxlJ7Nn
3qHJgGjk4d6ayLQsHUJmnYGYDB6/fAP/sqFtdxb0sd+rbbXmiQVKF63ewmDKVMyi
X4R81w2GjAadztccSfGfvGuB8v0MiLy2RWCMZq+OEX4EywXvgUMYkeR5WixrhuGY
Vrqi8CKf3rVx/jS/osi+34mnwnx0bVmeMMtJuEpdQFM2Sf92vkAet/9BVjyW9Q4f
oeqLv0J07xBgUiF+RGBJCZ3N7NZ7YjRQfP7GVKA7VXNMlyz8Fnca9sx8tvUruW7a
qS8K7CEeVSciuvGLiXIfmICfd4RPNzDw1Bck2ywC1ml7aetZPIYdQXwUrUBta7Uq
RiY253zWbUnFrLDvXIrDVy0NuGNsWaUcfaMED+xAIONavFksmxmKnoiiVID9yTZP
69WsVdcHaiQTPf/+y0b2RDaXQgtxDTlIJCUhRcM9X5xnQGi02egj3tE2Hr+2aNap
ha0UWSsvUcAzOLc0zxMGU6YUEr65MTjAu0eRCRdujJjLUXWiS+HS7h7WpIF0j7OM
D4NDSQG8GLm3EP1Kr65eEPbrz/HR3/zvBBmBd+MBXEvLyjQU6PAx5BTZGV2jXBOh
n5XAVBI5cdbXB8Kl7QIHojaXaK5QonWbq6A6Ml/YmIGrPVeAAzTDXYgjxeXlXLeJ
HIO4u+hpWffb3I+6lMBp7shIMCUOf/VJxcwna2nZTma5uhbjka1u0mr1VNO68587
tfEgHvAFrTDyeGJynsCFIASDTz7a03D5kVrTp0YdpLLGFwiiE4CHGydaF+E8tDve
7oDy9B4OaZGE9FpcbAnnvd6k5xmWrYV4XZPbEZl2Kz+E9SzsnKJiqoZ39NUw8k5i
V3g5tsiBZn7hVfw3S2YkoUpzXO2ArgH29WPGC5pL8zT9vHwUfiV5aYiuQx8LE8le
k0apAU8pERj9w7Yc1drTNAC2VJIkKhHrmj0/EGEj74HI2l77GxlKjk0lkjcPECw6
AXiTOlScQ8V5eA+WxfacuagQZBFQdOszY6q9HtRM97pgUl49bgSTjNPoFmWMii0w
9L9xTHRvrLcXYEmxO9EaoEKfYYF2PpdwP/Lw2jCODWVjES3tQMsPRo2uFhOPFzwM
+ZhjbXX5zK19YV0poSbpk43B3DTeFv+7BmJb1ZymH2iZP3q6kUmJW9ZvtvXByzoy
`pragma protect end_protected

`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
a2rqOFSmnLzZ1Jvo+VkdGNDvTbIJPs/fgRc6VLTIsMQBsZ2N5rxkgzE21A1tWthh
DgCbIILBeE5kuws0V88r3NHSLeuA67gQ7jq1uTT61HJUP6e4z4AJAed7foT8hkwz
tVcj5kdAZrKv1w/g7rT34A80j5ntJ4fUnU1oMm4tta0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9966      )
JzuuLlcIw5ajESjYjYFyIAjUQNxGWxEoxiGwf6i2nQ8QGy8NAQAa2bfJ964tHW+a
M8S+uadWIY3JUBHm6IGzsPfO5YDAkmO01rKpMwl0jRYE7j2Ogua9pG9j/1uhAyJ5
`pragma protect end_protected
