
`ifndef GUARD_SVT_AXI_MASTER_AGENT_SV
`define GUARD_SVT_AXI_MASTER_AGENT_SV

// =============================================================================
/** The master agent encapsulates master sequencer, master driver, and port
 * monitor. The master agent can be configured to operate in active mode and
 * passive mode. The user can provide AXI sequences to the master sequencer.
 * The master agent is configured using port configuration
 * #svt_axi_port_configuration, which is available in the system configuration
 * #svt_axi_system_configuration. The port configuration should be provided to
 * the master agent in the build phase of the test.  Within the master agent,
 * the master driver gets sequences from the master sequencer. The master
 * driver then drives the AXI transactions on the AXI port. The master driver
 * and port monitor components within master agent call callback methods at
 * various phases of execution of the AXI transaction. After the AXI
 * transaction on the bus is complete, the completed sequence item is provided
 * to the analysis port of port monitor, which can be used by the testbench.
 */
class svt_axi_master_agent extends svt_agent;
  
  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual `SVT_AXI_MASTER_IF svt_axi_master_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AXI Master virtual interface */
  svt_axi_master_vif vif;

  /** AXI Master Driver */
  svt_axi_master driver;

  /** AXI Monitor */
  svt_axi_port_monitor monitor; 

  /** AXI monitor performance status */
  svt_axi_port_perf_status perf_status; 

  /** Pointer to common class */
  local svt_axi_master_common master_common;

  /** AXI Master Sequencer */
  svt_axi_master_sequencer sequencer;

`ifdef SVT_UVM_TECHNOLOGY
  /** TLM Generic Payload Sequencer */
  svt_axi_tlm_generic_payload_sequencer tlm_generic_payload_sequencer;

`ifndef SVT_EXCLUDE_VCAP
  /** Traffic profile sequencer */
  svt_axi_master_traffic_profile_sequencer traffic_profile_sequencer;
`endif

  /** AMBA-PV blocking AXI transaction socket interface */
  uvm_tlm_b_target_socket#(svt_axi_master_agent, uvm_tlm_generic_payload) b_fwd;

  /** AMBA-PV blocking AXI snoop transaction socket interface */
  uvm_tlm_b_initiator_socket#(uvm_tlm_generic_payload) b_snoop;


 /** Handle for uvm_reg_block, which will created and passed by the user from the env or test during the build_phase, when the uvm_reg_enable is set to 1.
 */

  uvm_reg_block    axi_regmodel;

 /** Handle for svt_axi_reg_adapter, which will get created if the uvm_reg_enable is set to 1 during the build_phase */
  svt_axi_reg_adapter reg2axi_adapter ;

`endif

  /** AXI Master Snoop Sequencer */
  svt_axi_master_snoop_sequencer snoop_sequencer;

  /** ACE Cache of this master */ 
  svt_axi_cache axi_cache;

  /** ACE Cache Monitor of this master */ 
  svt_axi_cache_monitor_common axi_cache_monitor;
 
  /** AXI External Master Index */ 
  int axi_external_port_id = -1;
 
/** AXI External Master Agent Configuration */  
 svt_axi_port_configuration axi_external_port_cfg; 

`ifndef SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
/** @cond PRIVATE */
  /** AXI master transaction coverage callback handle*/
  svt_axi_port_monitor_def_cov_callback master_trans_cov_cb;
`endif // SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE

  /** AXI Signal coverage callbacks */
  svt_axi_port_monitor_def_toggle_cov_callback #(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport) master_toggle_cov_cb;
  svt_axi_port_monitor_def_state_cov_callback #(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport)  master_state_cov_cb;

  /** AXI XML Writer for the Protocol Analyzer */
  svt_axi_port_monitor_pa_writer_callbacks master_xml_writer_cb;

  /** Writer used in callbacks to generate XML/FSDB for pa   */
   protected svt_xml_writer xml_writer = null ;

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE
  /** AXI Callback to restrict accesses to overlapping addresses */
  svt_axi_master_overlapping_addr_check_callback overlap_addr_access_control_cb;
`endif

  /** AXI Port Monitor Callback Instance for System Checker */
  svt_axi_port_monitor_system_checker_callback system_checker_cb;

  /** AXI Port Monitor Callback Instance for ACE-Lite ports of CHI System Monitor*/
  svt_axi_port_monitor_system_checker_callback ace_lite_in_chi_sys_mon_cb;

 /** Callback which implements transaction reporting and tracing */
  svt_axi_port_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_port_configuration cfg_snapshot;

  /** System Memory Manager backdoor */
  protected svt_axi_mem_system_backdoor mem_system_backdoor;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg; 
  
  /** Common features of AXI Port Monitor Component */
  local svt_axi_master_monitor_common monitor_common;

  /** master agent instance name. */
  local string master_agent_inst_name = "";

  /** Address mapper for this master component */
  local svt_axi_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils(svt_axi_master_agent)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name, uvm_component parent);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name, ovm_component parent);
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for master_if  
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /**
   * Forward TLM 2 implementation
   */
  extern virtual task b_transport(uvm_tlm_generic_payload gp,
                                  uvm_tlm_time            delay);
  /** @endcond */
`endif

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * end_of_elaboration Phase
   * A local factory is used for all construction within the VIP.
   */
`ifdef SVT_UVM_TECHNOLOGY
 extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
 extern function void end_of_elaboration();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------

  /**
    * Updates the agent configuration with cfg object supplied from agent
    * command component
    */
  extern protected function void vlog_cmd_set_cfg(svt_axi_port_configuration cfg);

  extern function void reset_is_running();

  /** 
    * Retruns the report on performance metrics as a string
    * @return A string with the performance report
    */
  extern function string get_performance_report();

`ifndef SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
  /** Samples the trans_master_ace_coherent_and_snoop_association_recommended and trans_master_ace_coherent_and_snoop_association_recommended_and_optional covergroups */
  extern function void coherent_and_snoop_association_cov_sample(int coherent_and_snoop_assocation);
  
  /** Samples the trans_master_ace_concurrent_readunique_cleanunique covergroup */
  extern function void ace_concurrent_readunique_cleanunique_cov_sample(int conc_readunique_cleanunique);
  
  /** Samples the trans_master_ace_concurrent_overlapping_coherent_xacts covergroup */
  extern function void trans_master_ace_concurrent_overlapping_coherent_xacts_sample(svt_axi_transaction::coherent_xact_type_enum coh_xact_on_port1, svt_axi_transaction::coherent_xact_type_enum coh_xact_on_port2);
  
  /** Samples the trans_master_ace_dirty_data_write covergroup */
  extern function void trans_master_ace_dirty_data_write_sample(svt_axi_transaction master_xact_of_ic_dirty_data);
  
  /** Samples the trans_master_ace_dirty_data_write_one_ace_acelite covergroup */
  extern function void trans_master_ace_dirty_data_write_one_ace_acelite_sample(svt_axi_transaction master_xact_of_ic_dirty_data);
  
  /** Samples the trans_master_ace_cross_cache_line_dirty_data_write covergroup */
  extern function void trans_master_ace_cross_cache_line_dirty_data_write_sample(svt_axi_transaction master_xact_of_ic_dirty_data);

  /** Samples the trans_master_ace_snoop_and_memory_returns_data covergroup */
  extern function void trans_master_ace_snoop_and_memory_returns_data_sample(int snoop_and_memory_read_timing, svt_axi_transaction fully_correlated_xact);

  /** Samples the trans_master_ace_write_during_speculative_fetch covergroup */
  extern function void trans_master_ace_write_during_speculative_fetch_sample(svt_axi_transaction fully_correlated_xact);

  /** Samples the trans_master_ace_xacts_with_high_priority_from_other_master_during_barrier covergroup */
  extern function void trans_master_ace_xacts_with_high_priority_from_other_master_during_barrier_sample(int is_xacts_from_other_master_during_barrier);

  /** Samples the trans_master_ace_barrier_response_with_outstanding_xacts covergroup */
  extern function void trans_master_ace_barrier_response_with_outstanding_xacts_sample(svt_axi_transaction completed_barrier_xact);

  /** Samples the trans_master_ace_store_overlapping_coherent_xact covergroup */
  extern function void trans_master_ace_store_overlapping_coherent_xact_sample(int store_overlap_coh_xact);
  
  /** Samples the trans_master_ace_no_cached_copy_overlapping_coherent_xact covergroup */
  extern function void trans_master_ace_no_cached_copy_overlapping_coherent_xact_sample(int no_cached_copy_overlap_coh_xact);
`endif // SVT_AXI_EXCLUDE_AXI_PORT_COVERAGE
//vcs_lic_vip_protect
`protected
cGKTYa+X0EbCW.VJ6a-d,3S=T)HM?;fU:C&Zg-DbUCHfc00USeGG6(g#3D#eg?&O
FT#>OGIU9[>K<=J:-L<TSEEQ-KA_T885_R=BZW4R;Y_KWFV<(:eDM[&+GSRb;A?3
>^KI=N#N()S+2e4=G/R?+-48VdEeG:R)PP4eYTYTRHX,U0++Cg]H@13acA,T2T#C
JTENPG4/,Z(ea7U/#JHRDOEFWQ#e7#23P4g-H[IY0810,JJ0#E&+6E_XX8&D7dMR
6Q?W?a]/1ddJK;?EWRF@6-Q9PK45gc/NHODT-2H=&[B-R;aX=<?1^d_=X[WUC;SF
.dae^\.2J1Xf_+cOWW11/3<9)b]/1#1::CPJ\))90_L,G^A\GCE>=b4PCgKDg5Z&
F@-S.1O-/O+.R^1BVL7Q=QCbaQH7Z<0.Y9#VM[eZ_gJJ#1O1+H4)6R]]B827:YP\
[8Y^VbS?D70([BLH)d,[2(4ae/A_9aNE9$
`endprotected


  /** @endcond */

  /**
    * Used to get a handle to the cache used in the master.
    * The user has backdoor access to the cache through 
    * this handle.
    */
  extern virtual function svt_axi_cache get_cache();

  /**
    * Used to get the number of transactions which are auto generated. 
    * Autogenerated transactions have the the property svt_axi_transaction::is_auto_generated set. 
    * Valid only for an active component.
    */
  extern virtual function int get_num_auto_generated_xacts();

  /**
    * Used to get the number of coherent transactions which are dropped. 
    * Dropped transactions have the the property svt_axi_transaction::is_coherent_xact_dropped set. 
    * Valid only for an active component.
    */
  extern virtual function int get_num_dropped_coherent_xacts();

  /** 
    * Gets the handle of a snoop transaction to the same address as 
    * that of a WRITE transaction 
    */
  extern virtual function svt_axi_master_snoop_transaction get_snp_to_same_addr_during_wu_wlu(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_axi_mem_address_mapper get_mem_address_mapper();

  /** 
    * Returns the name of this agent
    */
  extern function string get_requester_name();

  /** Gets common class used in master agent */
  extern function svt_axi_common get_master_common();
/** @endcond */

  extern function svt_axi_mem_system_backdoor get_mem_system_backdoor();

  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);

  /**
   * Function to set the port index and port configuration for an external agent. 
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_axi_port_configuration port_cfg);

  /** Advances clock by the given number of clocks */
  extern task advance_clock(int num_clocks = 1);
  
  /**
   * Suspends signal from being driven based on signal_name value. 
   * That is, the signal will be driven low and will wait for a call to resume_signal 
   * before it is driven high.
   * Following are supported values for signal_name
   * - awvalid     - suspend the signal awvalid 
   * - wvalid      - suspend the signal wvalid 
   * - bready      - suspend the signal bready 
   * - arvalid     - suspend the signal arvalid  
   * - rready      - suspend the signal rready 
   * - all_signals - suspend awvalid, wvalid, bready, arvalid, rready signals   
   * .
   */
  extern task suspend_signal(string signal_name="");
  
  /** 
   * Resumes signal after being suspended based on signal_name value. 
   * That is, the suspended signal will be resumed back and respective signals  
   * will be driven high.
   * Following are supported values for signal_name
   * - awvalid     - resume the signal awvalid 
   * - wvalid      - resume the signal wvalid 
   * - bready      - resume the signal bready 
   * - arvalid     - resume the signal arvalid  
   * - rready      - resume the signal rready 
   * - all_signals - resume awvalid, wvalid, bready, arvalid, rready signals   
   * .
   */
  extern task resume_signal(string signal_name="");
endclass

`protected
75,aRI<0?0<.JX]KTR8<^5J.;&)gS3agf+<_[)TaPPS5#WJ7;>]W7)>\WEg,,Y4O
K^ZSB\_)L7N0349R\bU2/W\?-a0JH&]gFMac5-Q-HCB/G0C+bV5a;X9fcMI3/Q/_
LI=bR/Sa.P[5:)L2)RL7cbDa#@;^Vb_Re+.>M<X<5_<>f&TfXa9T3CC&f[[_8/Y@
/W/3XKP:M1>Gg;#R\c]Q8WbP=)<XQD<U,63Q@O6A/AZReaR(3\1#AI37V56Ge.KJ
\K6SUeN+]>b^9f)JVJ>?:Ld)d4APLOVFb<(]@fS6Q,0bDefIaY[V-[:)g9dM+2@I
;5cVV@Q]&MadW4S:VBY@9HN^]JVg4TG>\,<_fR&D(:Bd=NaYYMDG;X_<\eU#e5(@
Bc0#UfOZ4UAFf:UU7BNN+>K@72.Q9^F6UU\?M3_A.:KUE]<\EQ^FG\<Y#6V0>]T;
DE0Cb>BJ>Xc(SO4Hg_H6>SW3>QEg+CRY+:R+ZYR=BL-1KS])0ZSDZac3M0RYgY:5
_?;VN5^U:;e(.$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
.]7f3].78XM]9SFH_K-#&G\H?WP.,WJE,LgEAOWQ(6<AC1\dWA(C&(#/+PD4QGbg
4J24f<;H_1fd]TQaaF4LRP.9F@6X#ea+V#TY@]gf^4aP?5e,J@92S^UWP#)@.dL5
V#0=<^FdeGGG5D6T\G44@>TXb>,CJ60R?gN<<-DS/DfXC/ZIa](V,P?d1>cJDFTf
e>5P+f^W1[b&fF36bI/TLBM^F]4YfNU2YW6:JR0a]b9U)f<5UAE&3C@+bXJKXE73
1]&LKKHMgdD_dMbB+EON/MFg:NA4<>I0<VE.Uf6-;^/=IcBLL+NZ2b7C:^YI-[fN
FAP)>_6<UI\FJ8MRdQ8Z/)+[;LVG221YD7UT2GE5Of+^#HZY1Cd-EW,0HP<EY(Rd
^3JWR0089L=:\3])=:<5RS6B3f,3O7N3P[-2[HQEUQb[,PM5ff/0^1HLJ<DB8\6Q
8P4P0W[_@TZ\ER#G^3gDQ]He2I?4AfC?+Cc5[#9M@_9XD+OSgb&T4\\+BggK;DCb
96MQO+9CbW#L.bOec4B8HR#_g8?V8CF>P(cE[N\^K^de=<A_RH(]0F<eKRC#RaA?
O\3F6ff[VO--A7RfI)FZ\L_KX&59,3(N5X(\(1^8N4(3P18Z\A^.#7)H8>9D-,<>
gL4V2=f9\<Ae<RRD_RbG@Z>?)ZDCM\cMG7D.Cb\ed.dG)N+Z>==bZ\D<@SN@>19#
7N53POZaAVP5Q5D[LZQC+B(]K\L4Zbc]ODP-.__.CX/FPN3&4KLA:3^.GPT,L,RQ
R74>e1gR:_:K:L]aH09O#XJ&3?:&e/CJ1g+e58WN_MC-(D=95Mb7]F10d-K<DTM&
DXU2-9GML9VYTc]?[=IORDePI)f(_ZI/.K/P90JG,>,Og,gU.ddf?2FL00E[a;C;
\&c:<9EVIR>;^X8EJ,OW/K@08.F;#W\-)G;O9(#c\a\^D;&T=[CP1=#aFV]@-a#D
P,&J)9N60.OfE^5fBaBg[aRg55QcVVdbALbba=E(PRbS5f<NJWfY3C<&4]=4QXbE
,NJO7Rg,2FFa+]b?aITPTNNN+a=B-dI[)NL04S@af3^W9KX)L,X+SSc+QY2^62]5
7b78,?ZM7=MY(_+>,S,gRR8We/5:I(_4)N.VBMD@;)F(#A4M[PL^-B++RE@;V[8/
<AG&#.>)<ZbcD?I-(R(Gc-@8&bb\N0BWMS6gG#A\_#07ScKG+,dVHdU=X[LO[cNg
RNb,C2<L?OL2P<3;Kc&M@b=H;06UTU+N]_9ID8(Q)#XKP(@DQfBJXcG@MdBP+dN^
Q,(If^_UMDX.RV8+:?:+dIf_F(Xc>X/B<(_WO>4;-)X+3+a4RT]9(T=#H,;?2)+(
<NZ]M6aaK50I9[=U6_94(D2fX;eB7<+H,VbT+NVG>MY)9FSa2ZXJM(QPO(L(9KV\
7MAS2+=TF5[7-X:OW6<<<<7LA-6W),G9SdV25c#YGA,XCVf><(7?5O,9ddLgX@MG
Q9eVL5A4C^MP/PM#Jg\HaK:gDKOa5?@JH3deNU9L0YWX7WKUY3e&[RJS#1,)[BXF
<1H0)[>+0XVcN8YGG:Z:3c@7ecae3>T+P93\TRC?@g8^.VQLJeO0^:B4N[Zf_9(M
,.0(Re>-S4<J4=P;\Y3QK^[;FIC<-T8BdBTgEb4.C0Q;9Z6#D^99cPQ()\[OIWPN
+8eXJV[9LZFTD>PRXCJ2V1.HR6SA-,JNPB^cH;/Y041NSVOYP+@3VbX.APJJS#I5
7af4#5161Sg?Y&G<D&aM_0_16Z8bDY>b4PV=R9Q&&=R_Yg?_dJ.[KbaNT97W.:DQ
QU<7UcMgL1MBJaXc,4^5d4:CE/IS11CIDB9_I4@ABZ#LW1\H]T>QR525;aZ6d?/2
3Q[@L[E&?N^&WAP2f#^f=MbR#CE4S(Lb&^+F@>Cg0NQ\Rd61BX#A>3I8?6I=4QJ4
FY.EL&[IbO_deceX2D/U#-(MJXZc;b+;IAD.?6&[Cg@^2M+8QV8d-7OVF2Hb7HR-
XWP&^GaBM)D55&X(C_O1V4>=+0T0//_+EUefd,0M0b?WPF9[+=.a[-J@N)-[RY[f
4fe@)g;6O(OK3/T_]CW?Y#aTR18;=ZG6-aXV^ZL].Y07aAOABC<Y,R1F<SF90dc#
0.K+@8@L5,^UQ(^Z?HQ[7/QRIQHbG?-^L&f=:+H6=-7CK3NcGcbbSU2.AGBP\F#;
geD;(12\2Tc>)BfWNb6V=Ca9A2aCFLN1JSL_X5(e([a:Q#G0\5_7&PeaXO57W[B0
eOH>,B_-\7AMJ)>ME5/H1#JbBG]U[HYS+O^4&&-RLB4If,]:,_(6cO(PcD7[C#GM
\C-BdgG3[/YVYc^7C0D1AQG@\9b<^];S.WHcO#J)JF99#TTF6\bLDB>Tgd5&gfB1
^ffIf2W[C5EM[V]8fG,Lb/\I@J[@NRA/FH)RPWUB3B-]f/;4e=DQIRE>eVSc0OS(
8=4X5\BV3d:E#VUfN:Xd;.X7LHBAf5SM,b]VC-681Fb8,87_6GfeQ\^J&a#g=<LY
PdXW2_.4faJa8.V(09/0Ge[:S<.I83BJ?(>U9D37WcI8e.#)H9NP,1JaH_DOKB&\
/76aQK9AANWP[7fX_UJZXg,=TD2B19ZG.:?&IRVg]Bff5b..(^B,-D]X--+,NK#0
_WJZ6)-fO?X\_M;E:AQ:SN3BI0VOB9S;^db^3^151<aE^(XZR]1SHab,SBA66/d[
SG7aZB\>H81+&<VWfK9F5_B,W1(KA?eB=5Y76#29Y5UgAEe4L\9GBMKHH\NU><6T
0;DTK81XW?#H]a?:P:A3T)WLBfW^OHNYOSO_M=BPB,@ac]1D?33JK@+TQSS#9H;]
E1IJ41:VbZ5X6:HU][-&Fg4^YI)#83>_[S^(e-A>K;7+;K6Og8_6)57QQ4.4?=aH
3<6(I2.7_,U[KB06L#P3PL#[H2[R8)A6H?UKCJK_7LgUMe:]LDC2R7/O@T,W;7>g
Y@8Yb?T00=XdHX]DBbX,R?U#;S2>Y1-?Sb5OM0X9I-bA)Gb3@8:9Vbe[e&R=f29B
&]KF4J,9Q<]5S:PD0P);H(@KcRfD=bWNVWga58M1bY+(D.V(BB_Q63a)Gb]?]d.Y
S/W>_A^WYH+TPL1^>bS9H>>:Q[^3HU50[RON6QJCNc)MJ-.HR9E/aVAXX8fO0V#N
1(2O@BTUUM33O53RGaEdI_\^f-;bQ?04^Bdf?(#SJdCeI=NX;-/.8]/>?fgG85F^
K,K-:Y1[8^+ZGT;8<B(#FacXQ]02_5F3/C6)0&S[@IMI4?bU</RMJ7e_&,-S4V:>
&0E?=Kg:/eMUO:OG_7#a45:-9gVb/c5IegfKZaE<9JJ9bM2fY)O+N3YC)YPYI-AV
RKJ\DNI,HXM7#^Z\g0@8G:4<e&^:K[-?@\:T0&R_VECZR?+d.6^/91&?<#NQAA0I
GGEYBVf9XQdL8T3?NNSSa6)?JLA3I8O@D7H>ACXa+:@BJAKT@\YG@9/Cb?\Ma3J)
/EOXHGJeCQ+GT_-bcO-G6R_X#CR.,WU9)cJRS_4>0DGEJ#@11C;CPVbJE<3Xc2+3
b_=BP+G8S(DDDJRU=M@Q+0[P-Y;(eS7<FZK<45c(PR3BHIfVgAg<D</R>/FK3-eb
&)2B0ba1^WV3HDd3]MADLdD0c5DTR-DJ\1[cZI;f41-,Q5CC8Ge>S&LBdO8eAA^8
<Z.9daQ4NJ-+-D#MW@GL9L0T^#)<4WY=;,;WDEZXc78M/ZP_;6S8Z2c5aWSDCJ--
YMQeV9aF:b,&I@a=f4>9Mc2P?]C9SDL@?BeO@f3W;@__\T?568X8Q9:20Z[\ALDR
g3f,/Lb2Y/6\VL=&YU:N^H5,@Lb6[S5cB4KBQeg1HM@cMgea^+Mc(#&FgP3Q#)Gb
DPbXgbPWAO4g@B-c;=)L0D<=T4(^PNY,9,bb-&S1C(<E]3:c-467O[SNMQXV@@eZ
GHZ2eFW7fBQ\R-;#KgP)U]2Q@++&d9687C&AP\,=CW,AR10\)47MHT8H-b#/T6S)
YG,8R8[#CgV@6?3fG[Eb^a6/YWY[/D8&+8;e7RD@^QeS8=R>9a-\(S=(Y9F+W1<,
1&U2^aME_1c+@:^@XY/b/?H?(;)DgL_/\d@/6\W3)5dKfeK/L(R_-cL,U9O<048M
K-1;EYa\b(c_2XNZZGMP6JR\L_ZON201\:MP.I1e+BR[)@fRE-#^?Rb3MfMc@?+,
ZaWZM28XNEa?Y1Q#NZ::6HUWG?0^cXU9KSI.:g3LS<+AJ+S=@:?f?=B=@5\UN[BS
^KFEH9-V;f/O-MJ:YRe\JHRG>KCOHLMCNg8]Z+KK.(]VOb3&FK?9Ne9I^TS90</K
6J\eM-H>PK/^83-^Qe7/=/A9@e/bH-R/fPb#AY<)/=[OIYG81K7cdBX2,HY,S97[
[=GC(JHAZ/A1BXK]QF9K0RbS#Qe9[g[&0IaC?ARO/J@^HOM6G0I#QL;I<29\3VG#
G8T<_JPUZ^_bS1,-3b2+JO(_):2FWR6R]9X:OF:c#T#c9GH\IV&\Z/E6LE2A2g^^
W..XJJ0K5JV\+/31)OK[8^8?>3.#&[(/>)UT<6&P)NO:e,Q>L0-O@fUUe^Q?e34\
W^OYJSD,#T\J2P_7^8VO@:\=C-@=-#]a3)(+5M25>EE-d3<,\5P7[)95_F@f:)L(
\dec99[<&2D):SJ2(TFc)b,U8=8U@T2]W48ZD8C=LP:NVW]L3e-Z\^J&7RgKM,:&
S#^SRFOK4Je6I+-?:Nd.TT9W,(E[a9ERQ1\b0[Gg@)/X:5;U88BJ[O:,14@[C1(V
45)Z;X;G0NgeE<cK.RJf?[=e/(-USf3J/@A1[QF:6V+\W?WW8-#Z@UgI>3@;aNda
:U?^DG028gE85:=:e84QVea+X?[a]7(a>:BW+6c+c8C:#:ed=GREb9N]b6-88L43
@^S-S^O1I?G\b(V,[L5@A?eJ-@T1.<-?&X^Yb+-HfJc5@OH@H_cL@(HSA=5^&\J@
KcD5fVJ-W/OUMDcJ(WOAdN5T@=K#5B6#IL6eC.<YXB:KY0>b(Y4Y6GNdFOT8S^\K
O-;g#:.QT.;/6:8610TCb94DLf&TUF\JK;9,C+[:)bVW>NDQa.C\W])Q=X1P)^WS
KfG>NKN_.4f2D#3cUbAH+[@SI-a[;)MX,R>L=(_142gY_ZN>?1b_&)-+.X3a.?K6
c^_T7;cS]F8d:AS\fB;&6X?D6_Vd)7P:A6+&L@<,>HEP^Nc@:LEOQHaGPV8eUT>J
H[KUVDQDbD[RZ?CABgNBZ.STV0(Pb,X7cZS+0e/N7-OBEA&B9OR]D_\>IaRdNX>G
&QOc/S]Y8f+,X@AOObFHdgM9D(//7V_:P[1<dQE02X^3c]1dGBV3g4RKG(6F&:;A
KJ^A/abQ<O@^5D=7+ea<RbP>/_UHIUC)(VQ[:TQ^[P-UDG=,TS:#-T)Cg@A3@;[K
agb?6=R-<]>8YO;85NYa@H<L@B/+O=_H>2-c.8X++^2\11OQ,2LUJ3c_(DdM4c?M
+C^M)&&cC6eQ,A1M?F?_;Ge5O=_(]]6ObA3U/fL8]bJ)(S?FS(MJA<0<R_ZXSS(&
<3/>5cH036RT1\C>db^AO+\<:V@T6cEA]?49>R=C;aHVO\&>Q(EDdDdRMG#YG9EZ
RWaRg_X#f]Ob1OM/Ub2CcYD<Z\E?6S(6F:XPYE?;8P3=b7=N?=(TIT>#M#E9>)8S
)CRcc-?]<]4,I0IBG&<WB)+)H,HF5:Te,V6dA<cW)P);Ef=@d#W/:4XegE3]:Q;Y
/Z_L,^U2S>MXNVY6LZ?WT1R#f<G:[1Q(WEdGVCgP/eF+O2g?)=?5IA/^__e>4eXI
?YgOW1CYMK@QRB/7b1Af44K77<KO&Q&+]dZIJ?;T2(I&\A<bX11Q5ee]1XQ(#M5Y
g_-W&LIa2XQWF+K[G//+N0#9<.#@;UFRfZFe>W.&((W.g(Z=b6\LP\W#S,?;M&aa
C+W4GHb.7&5>:NIf<P,b_W0MPg05=_c(8ILbX\c+Ag^eUOR#0?]6/f?11L@71S:A
M#5?)026>,S8gIV?QNQUU.0[,[)g[KK0]2ND^Z[.AWII.T4Sb^DbTRP.EI.[DS]D
5Af;\CCIVQf2.7G61._97D;1EQW[Gd:?DS>aLZJ/X1P6X(J\.?:e\H41e0_fdLH(
8=75\@8>GE,e\E+^aW#ZN83<1J^WWPG,^B@3;5]]&X59:6(^((>gU-TD;=^@D=JZ
>C^XCD1\MJ;5#EG?g-KR9OZeY4CRS@>S<_,^_1]3Tg-a4M:Q^Y2NY/,&):9L9#Y\
UV-&XYJ7)N0]2:AJWNWX#AJF61U=SUQ6M&.bHM+V[EJOMC6:7LC[()H][2GW?B=9
<9Bd6De\Xf7f#Z>)_Ue\[,FUUO#B:fE4AddGe]4;7aMQPM15</US5Z1MR+IC?:Gd
JFff>+0G0\2M?G@-=,KF[X?H8:94bS5fGVb&_HZ]A06Qad/#CUCLCaH>I92)2PgS
_QMd:_&5AG]XCXFU=.?JSYHO?F/MOSSA?\H;_(TFAZ8b,.9U>3;&17O:_.=YV-S]
Z.T=L\3:<cf+^K+L#bO1bD6Bbb?(V@JLT5+EFeWD99?MEQ[B-4V2C-\YgQc8S)1L
BTcee]GD4F;-\2Sb.@[0YKb(6_?1,9D8SWDgD/;,D@(?g]8R)\WeF90YIFe04MB4
C^?F4eC,QP8]Xd5Q2\L/;4\Z4B31Qd0?DQM0XE.SA6VU-/Ed/dF>2>.bHHb3^.W5
1>4d>@V32Y7Ndbe8cK@2W3B\E7@VG_\[\(05.+)De2:ECHDAJ=AN-G3Y9?3<0Q3I
^B?>[(W8&L#3+48SCf6MI)3>E)PIWE;I71CSX_YL5:5I2[@,A0ZJ.+,4[R;^A,<H
:WcTSI^,C=A<c>([,Q9b3GA7.^2+T(:dPQ:#8/Q.<f;L1ff6<HE]=X4]Ae]#cN5>
^3V#SBY@-V]gKAO+FL7TD?=7d_Wg5;H?a<>5VGUS5:LTUCX>?U:ecg\(3d()/A0W
M211Gbd5D;NM_daM>\ZSV\(IC2;D7KP-?^=g1bbF?)=&H;\HD\eY-6E[2B9BaDM>
0?9UP/Q=Y.G_V5X?JO]=6JH3./O&cS;b-S0_\-F>6-<)&?9MG36bTaHD/S/9SDC+
C,.+R5cUaJC7gf0I7=17==MJ<>(f1P[TW:J-5C(.f#6>W&)^HW-AB2>d5:1L).\/
W6TIT#(^<gYRU\BKcJ^[S\YO&,U9.ZM>Tc0Lf^H/6=:d+AQBF+T9gLb@R5Y)H^52
0@]WL4<fFZOcaVGa1fN?84;gXM.[a;7.I47,X+fQ;P+G^WC7ET/^9Zd0WF7HC4NS
/M\@.5T<#JE:d/]Z+=Fge;de^e4cS[6+&C/&L:g1a4e)_d(NHOK]5]D7.XKS<f)R
8\NEA8/[.NEZ:c0#S5SfBD)7B+28X(.;9b?OF-)eL?S&WU4YFF=fVcdO&MU27X=A
O5H=aaND3J6N>Z@aWO-QV?&g_Nc-GTDVXXQKg2/,VNc(<5[82)f=:=.cgNaTL7G#
+T&bD4d>E&:f](0N7Dd,(0.5JPIL6aE?#>?62G.YF-=40NLTUNKS6.e45G0LL,CW
cW66+acR^<H77Fc;M#AMEgVaZF8bA3V0cD;bU?L3UFO&/2:)0e>=\&CFSO-.ZKV[
cZ#=9U^g(A.5ZJX?<=PH0^ND>UT.BCE96DaEV<ac8,f[Q]9(dEAE[4U9.BFYHJ\<
(7G@+KI_(0Ya0;gFGgFggEMHVIAV=7M/S=&CJXW_/DN6;Ggf;W3O=d:d[\1J982g
#V5H9&945_B,,Oaa?=@56eZ]C62RPL+DUR,S12FVJ<A\..Y8_+a8Y/T1QQ5;R40(
ZFZDH<U\[K7D/J)ZC9(U3CMJb^ZE-L5T0g\WR@8H8JKDcZ91N_H#3&/<_7^+O8Ca
R[3Z<65R3J57E]W]B\WLME\N<>P@G?Md=C0Y8:N5S@SVfHAX49\;799Y?<Pd?)X/
V_Z_df3VYVP.:SFaO\,.8EPHW&DY3+&;Y3F1UGa(V:7U0DS)_)[W-EWdD8NH<-@?
-J).RVBUHE&_R36?:B7e0gZ@=(N,QeE);P0CX#3geQ)aa^HdQQHW#YS(G.P>YSFA
=0.H2L]A]+OM5:&0]/.Y81,+))5WGbK[6&CP(eBCY+1DgL55/-?6a)EO>\DQ2:f5
:XDU6;(PSGQ0M+94(>0RV4[gPQ:00)KE]G]7A.fUA-C+0OdcR<6KO.8F,)(40+[S
e][),#)<+AW#1O+.(8OUI[L2:gX8MDG(;eFHCCd&V8481PZ:1=.de.RHZ[U6=A)/
VDWJOJ-_DYB).8d81BC4eNG>bc2L7(R@_\:-+<?@FAY0g_\2._^bKV65c]_.34WB
Be>R&\^;FGI(9?#:/H,S:F/L=(>:&6YIO>XVCb&g97._V-WETYFTN,J,c:MB6#Sg
1]^@[M:ca^)7c3514440FGE7_[<BDFd&_g0\F4d)4.9V@RJ3=:PK#0&2KDd\5;E\
8?b\-e96PRI&8,F+)=b82WCA;R_G>[TUcCXcGN;W7AROY\LZENc-O0E^ed?KMG&8
B1+9><UWIS6b<Gb@U3da7U@4O]4(&F2Q(]D8.U@-U;WLY=1Zeb8+NP]/1/=Y&^N9
BH1R?HM[G,#gSI6K3[=[NH(N+>&>?ULE?cYO?.:b@^CRQ&&gJIKZG(LX4V_<_U4[
9ARMS7]cPUb.K+UddVANagQTS/B@-U;F,PN#dPR=MB6@KQ/@3aY84GEC19TYOJ1B
\QR9.AX_WRC2VU3-[213W6J+D-eU9=7TTTMg9BEeZ6Yg+86;X^84f218b9O;9P2.
FgZ#SGFc^>LVI]/_O:52de@74MX_c[@CMBOIL#FB+b3K-cAZQ1+>b#&8bY15W&TI
R1]SM<Rcd&-:+=fDV+T0N6.3TK\6,<87+GM81?TXQ?;>?OeaZD3\[:S&G=G]D5#+
7D(-OSI3/SUP:&28RfJ9PJEWX9(X.[V2T1:UVKC-W,LAH#[)<[NaEYW>@FH,]8S<
HYK@&+VL\WR,#e9_bE&-XY:c),ET;cOH&FK&+VJ<P_Y,NI<Z?-UUF,.#3KOZ@d&Y
;cG:@E5>+LQ68gDY/M8_7#[8MTJPRO=)2U9eT]f]Z[GS.(gfHE?JFU74=e^V=(52
A+fDHZDX-M)NBZgXFgIdROZX^bT0=#:DET/8[/+K=YQG#8L\,cZK^f<#Y5;?161-
&R2GUec?J,E;gDA]8=.F@XNcV-6;_D2[?V^?PD:6)8PIJO[B[&4@aQMGWYQ.L24Z
R2N5)[KR0@9e]M_NJC_HLM\5B3U=QUb9W?SXcD79=SE891dgZ.HW5(=E]4,+M@1F
T0/75fa-c-[=M&C/(-XI.>cZW[VJ?&bGM-F99+9.JeFN6.O_(>I[Qc@JJ(5c)(fK
eR,[b=8NEb#PA6c4C0ZQSD;\_QGHII?_dff[_?RI/[Bb]AaZ[LaIJ,^3[7F59KTK
ZW(^4[Z,=P\M7EQX@O]+35e1O?QYK6\d#(c?d90N<U(D[.@Ga2[1U>=aNF1:PgK(
fLW\??+E4_e;BEeB))EPHb2R<=&=,T-f@f>/QN2?T,7L(<8/+0>R1)T[-M]:<,PL
3Q[W_-1IAVSGOL13.QfUL:aOgHDB]WLZa;Lb_A&A<]c_d/(<5BZD,W6J\a8fe<0P
@:^#+&KNUL>NQaY-e561bJW:B0A;SU&eSKF/a)b1X13>V(<@O^8d)7aD_?>9P?;@
J#](0H-VH]6-?IOL<X[7K<@W6A]#SLb9#N:)-:+=-KU4S-_.Z6FW\@8VWaZ_aFSM
[^F>5+gW8bSJ6C7EIfU^V^:fD6[:AD160ZZ4=-OD,UYIN.MB7Q:g^>LG\</a&=6d
O2Q8VUd)&Hb5:)X=KFb;Za>AMZ<]-N7[N(TYN&6)U3bSW)\SL/;&fBcO>.P^Xc9]
F#-&N05;WFM2G)eKf\aSbWY-U\fBd11G0;.7AZ90WJ=/eE,VP5YJDcdPZ&(a=^+g
c([-AXJTKRFF5<.<APeT41HA?e,MP(fa]CH/BCZUM::/KXgBMXVYOfg70Fg+E(E+
8#;B:A1QI;.?d8=4&N&FMH)P_34[HbIf2VaY-_3c?6a/-=VJP:YS<4Q]KRcTHWL7
F?36CfWKSeL?M(-225]WW2STRWDSC5#JR4:E2F6X:V^2MWJ53.WCF=7B[P1M/XC>
+CPO:VT741EUD_#>eE^CJ7J\7+L;/-SAQZ,bd60AZ@PVT4.FB7B?9O&^-U;=;F+#
9/1>Q+a6+&+ffe14T<&P>TeWRL?XZA3cRdVe>Q:EKA;/P#_f,?:&:VYH<RVeQQG7
1&3=Ce&M8fVD/_g#@&:/FNO&0gH;ZV8>=CF9N#g0,5::6<+?V#Z5ePe:TFQ1gJFb
<#X78g?.(;K:#da/[(>F>D-bbQf@1\]0c5]g84==?2J2Na?ZWT4B@?6P1XJ/0=4]
9CGPKd2,R70>L<27Q(<QE/,O;;_3GJ,RUKM?Gd[fGOOb)&_S;&922f?D75?]<?@g
Q=Fg394,F/JKY@P280(9:XP:FYWcQ:-(]M2\WP#O?74#FCWM4;;PGP9_Sc/V_WGG
R.:ZISaE&=]ZWWNROZQH:FJ/#R\/U6_ER44Y7d0eZB5H-CQ)J_d0FJK36V?F]+LF
:e<Sc5W-2,G^X,ZH:aA6)FX=gWR&@C1X[?aZ:5bJH[MKc94cUTW?g0:K>RK0STQ:
=N7]ZM5:)##O:72QXeSB1>.#YLGU03#ZT5&LV_#O2/HL\L,)>:f1Sbb(R-RN\=3U
T5O^SAFQfL7\6fF7gH0Qd9HM\-5gfeO,TcR8&-R)gSB(R5R>&d5.^OWTQI^)6B02
R&@#OJScLICU5=-;-fT4eHP8GWd@d1[QFRJJ?09W-Ub5QFJGIIH)?PN=aQ)W8M&2
:X0^7QHdJddV;dZKU_T0B]N4^?I=JKQC<,(d,4MHP&8:L37+fP.^F(2H??DbK+/M
5bZ6c4:FGQ^3g&3[5N)>@B&.](b195dVD&^GBa+BVN354H95U8C:PTX+e</M^SS:
<Ad_gXFc_#,<GCW82DGec[TA=S/QS/^+gXO@ZIb[KE2:;1e,>F\@bX?+G9W_<8a7
g8WNS[;_&5)@_L1+Qc9<^)B_RF[-A5KV4+(VdbM36IECVEa6NP/[W+>G?7Vb<^0O
E199V=A<F0YI.C-U38;A_F/XN0:N[P.cM&Fd_0@c^3ZEND]1b;._SgM16Sd3K.[^
_R>T)><AS]J#/@\_f)GJG?5.9Z_88QYTOWLfFO1BGC27H#ZU@=VWVZ48e.e?U4(c
NOJBg=aKO73#1d9Od..7S8HX&PF#bfbL0G^X_HE334B<(#-=#5CY-V#LDEd#45[8
=(WT#?]6L2U1K[A]CJ+LEV)-F>L_X7++5E0HJ)WQ)=CR17L@]5/B:Eee>;dU[<Mb
c_=J(;c<?a?[=5B2H^K#KKBO&eM+Z5MTT=b@B(8;;)U.O>@b->L.^a;QaO<X@[9&
KMGc=OT8[T@Z>f?SecL\4gW+Q;6WL&-R,4Zd>b#Gf4\-5;#I4E0YC2d\d6GMRDac
^Y=c=WPX-UP^AC-]\f2;LeY=^>(>UN^@N^]Te75Y&+gP?eICP05AR@=7X;LI)7&c
AaF?cH6=5CP^U#[X++#RFT]QPF#aY0:gR[BbB-d<,A+/>]b21>+:HI8?_2HHE@d>
UdZDDU^d[=\8Q1A@V3RKg;gba9NWWDYQ75^254Nf-+/US=&XN:N^_S^HF010VcLU
NC7I,abe)T/G96B(ZM++1==Y5U-<YUb1.\R(_T8FcBK+4/1@\UMDGARE<RM-N-Dg
IM]0TXfR46&:-9#A,ZD8\gdaHC/dX>+ZeHZ_>gVB1Q7N#c-:E[^&D#GNRXHCJF?f
g<M7LW17H4M<N?3#X0-[;NQ7SRI>A)-NEHRg[(DRG@8?3E_0)afgP?JLV,L5GMWc
bRARI+W83OD6_:D0.BZARQ991PCCH,EHTI4T>S/Z)@>V_&@)LT>O.D[_VfK+e<5.
NF^d:gg(L+Af_0a/G:8L9JgC\Z74_5/,d9g\TUV7Q/2SfAAJF=Y7K71g=5dQa0b1
9T(Ka^>B4M&?-K/C]GDNAJaB5]+e:R2YaFO;6Ff1?XVK(PB\eP?Ie=&>W[MKVX5A
4BA:cTf?E><GO,K)?/#=\?N6YN7Y&CQ=WB)+,JN9IJ7^7[C-C+]T.XM>)T;-?J2B
4C>7eO<NC4XD>MTAYP=SY&5J+9QAZ1KO/c>;;GdW+VG;e2@?K9&E76b)+a)SKa[B
JM0MU_LC]R]?MK,+ATT+9Z\^>aaR4U[QMdB1HF8?gRK]]HgVF5aAB)+Q(\W1ARI[
N=3SeG2b<09C7YG>a1E3f-P\M72RNMQ==CfE&CJX.-\N<F=?.U.Z@YF9ZZ[ZLZB9
,7KGE#5,fA#<BD_#<^Y)N&&X[FfJ.N#5#9KaTf1fJ8FE)YFDGcLKYD)3#JcJKA^=
+L?3^D=B<#\5bN9PJRW,LaM<TMN+XRdbI5W3V-TB>=L>5W0=:A>FRTDNLQEfL@Uc
J59KRAH9?0[A8.6)MA[\c(</FLW=(>dL)N.\Y+Z.;=fOLK<c9V949A=,SBZMD0E7
BUQTE:fN&O.8RdMRL,>3-EX8QDe4b?=6/U0YY;SFaD/eXE&9#-5+TD-\_G5=fL\E
Q&Zf2T54LLA+J7?NH-2Mg)=b+8R.IOcC0DDLgBDP;.+Ig:L:\780EObKTfYCGCaG
gAWX4:ETBV?I2EEc(=PgQC24+Q4F[3;5[@+A35M\La?2H5&N\gLPQ&<W6N:N2J<X
]M&ERY^(2>9(Ce@)JDcQ(2P<AFNY?3bHeW5bM.Y>2UHU&M6c/?SB9XGMa8@:/_,T
644[V2d=L<2@+F)E>U/(F<C16Tb.5CXKU=66@J;MVfL1;E\&f^N#=W6&HcFd2E@H
Q+H,.H0121V3X-&1H0#J50U-JGb,#O6\P(WX[\-[-E.=QMAU7(V+E/_E9g8&I&<V
;a>56ceIODYHVE;72^eB(WN9ZD?eD3W:FZ0H(LDZ()7^d8#[_DK1CSLOWFF)D]DZ
GQbLN5V-K^gIag:B1X]ba<+DNO=@V]=&)K4GK/=N]6M@bY#_ZeS=^SfRSQK]W6ZE
<.0#.g#W559\MJgWg)g,6FgaPDX:-=NRD4D-=eFaPWQTRGDC>J.d]4e+Z2e#D\QK
_C3HI\eaF&/@-1<8>ZX[_:@(HcBVe-WU9/?=TZ[#F_E+c).SB>31(<T#d#I[.f&-
8)&8a;fXT=D47=45O-A@E8U1+^L>eKALLIS5&,d4[DCT6ff&<LAbAO<?8R8RG/VY
4T>WgT;K+@&4\H5_O04bY;OaJJZc>)IdUW+XO49?[:EM,=LcaPB?68;Q#N@4Ne[[
f#&:/JEJRKQH[QM4J5MW,@IOTVU.#SQ08;<6c-Z#D0:Q#9]e[Zg6;ETBb?<?719;
\f^<DT@.JWM8/O8?R&TK,21a9ODHaR:.I+dN@TUd3cSR+8,X6>1/0R&[b[Jc[L]#
IZb_&JO6LVCLW4KNf0g<=X:UTH&<@-KPJI.fG6+)\4(I(ADZ6V.P4Q#bSTd0TfL;
e:ESe+;/)NN&K09],X1PS7L@R6-f9cg4<=AG7faA+)+J[d0@HJ\.HA)bTRCTEX2=
?d[ZR?9dc=L,J4C0d]+@G3V/Cb^=DgVPb)W;LYPFEX4QDV_TZ4a7e2&93)/e,D1)
)PV08;c>B#)VJIMJQAR1+QeE##?9^5[KI/\g>NdI=^T:Ze^2V]:d2<Z9YXDZeA?^
KI8W4YcT^:&2-e5<X#/D:d\CaV,+,D/cKN7J8WAH2&-c7);J0U[0+,;\E=3;E&:B
>5BA;_Le];W((Xe=&L:2=>We_J0Y2f2L;1&YA-DdN[RB^ZUIU]#-S-<8dbQCgCR0
X4FeJW>.;4TZRg4;Q?08KDe-^2LBO/>d0G5[eI2Y9>JN5SbIE[=S^c+c(4.OR4-[
&d7g=UGaa)Z;-FRAVDNN#G#4K4R.].fP(CZb[@J<[RJEO)gD3a;@9_b<^\a1;4V3
JX5R3KN,NB0e#NR(DPeVF8T1/d<7G_HAEUN1?B.XPU)DE[EeZSN4<+QcaJM5MCbY
U0340\4UV#-MaG_:fE7Q;DC]KRHbBO7,B<::KgR73_DgF]I:\0K_1RX]>;1PAUUK
d9S_N[e4fS<MF]GbE4BLY_R?\cgB[25D\G?^7AS0M7.7&@aNWaYG38<f8.eE)LO\
;\Efcc,WYX6\[95?.-_QeG5VL[-eX-G:1Te[FCW4TTWaL:34eK(Y&Wc>-)H.HeTW
[OY9gF5VM9;bJA8>dB.;#?FIJ6:b6Vg/EQ+I6]>T8.ZKG9MJ[DS/9KSOFLBB9=JY
]Jc]C.XH7cQaTN/4@3?FJ0:,gPN07IE7QPU=(=a7X=Y#WE5M-X_UAKbNZfJ)YXeC
)dL,8[A3S<eN#4EUa9TcAC+8L8Q9L97DPKA(6^==:F[&CF+7Ud9>11H^+;10=E5#
?]TF2X-EOQ1A-O=]fL0B)78gD2VOLgFP8DA6EK7Q3KF5P##=^EN+H6S]&0TQPC00
egdXYSB.[R;43RY>;LH);adXE(IOF<&_RVDMQFQM_6]^^MM#CTY&S]aHD7#W\YL5
8,>ZMRRPHa0V[RMf;;]:#NH]/2=B,D<[2>+F(]Y&UNS.a-OA@HaQ9K/H[.=6.]e2
9.TS<AM/I7:HIR;R/S^c_->UQ^/4NAcGD(K4I.QR;MWc#&;gUb@LE.#[#Z8Y[g8a
fQS51&IMYHf\XODccI#?3=)M6T\Oc0A^g/aCd2\SWZLS[e)5Tf-4G_0DI@B@4PAP
OY&)=1Ue->:beB2CD9B9UAKMR24f4(RJTJ_a]U-dg9/O\?[E6PL;]G@cd0GPD5##
/LY,A&?]8ca/fPKQP?@SUKL/:U@]f[6MDBX[R2T>?HC(E5,^;WAH:OX;3/A9Lg_Y
@,6;TUWQaf0f(4DCLA\f8D6bEeH&@2NE;V8N0)2?BW49(0_Oa[O]IHQ>ZZZBbWU>
ZW.TfMW17654^C&6OUdL_J,YE\C=g=4>JS(-(+QMe9Ke>,MLUETI6<dZCA8GGB^=
EbVPe;A+EHcH>+Hg@ID2^gc.MV9ZcXb\DAR5&IQbW1[/Nf2OU034/0OQD7:\WNa.
UJ_Ea.:SBdJ^STPIM2&^;d+QaIOV_b\[]/]H]U#9b)aJ>NY;RD,@Od;5>]#J<LWI
>:YA=U4eHYJ0LXdb_[7[QHLTdI=S7,DZ-(#1#aIcE>@DJR>d1\4\(([FJYd#-?DY
&eC[GJUV\)N8ZW63F7&_V]OU?)QeZFe4LV;;/Sf1#;XVFBJVX3]R9G6SYS,WJ.a(
B[&E+P7OcaT;Z3+I6ggHb(.YOf7U90gf5(J@<@E&BUa-8A2)9eQAI8:A_4g7BG&[
E=?,N[QU3.2MVD39g\N21VZ@3<DFFK=LaL##Md4>0]^I+(;U=C.;X<7eKE6R3FRE
Jge0-?Q0W@M?f=+.WN##Q=fXEI3L]I]cL/UP_575&6:e<;90ZU7^)5+A/DIYA]H\
a5]\d8:a<T-V3<F5?GD&/U<#c,8W,c<C:e4d^R0.#I#df^b9PFG/KHAO0MTX&BD\
Ia<+M.R.E\2bVBA2M/Z?R6PN.6FEe^31:X(R8bD1)82E0_)X<HObR9Dc<dHJBXA:
0P5e>Dc[3Z;bRA,F51TCDFFcPA,U<,bDDYB]J5VMOb@MJ52E_9+gb<+I1B]7953F
=I9OL+Ybe1@aA.[e.BQI\=2CK1]c/c^#BLcKU=S<ZH+?6)R5-BBV>LXCdG,\Z5cV
]E?>UMc)7A-baCG^^@3\[+Rg[E>B9F,B,NQEP:c&ZWYcRfdWa-\ON/_X[dRT+_Yc
1TF\G)((WR20\J2_76T/XW1c]VU+])X39^EY]ccT58AC=WK_f/?=R0NXC<La@F1^
DgEW\eL\92>cI)\WA^ZW86QA=DAOBK_PcAC?R<0OJICf3KE5+>.e,OagcZVfU/.C
g[c@T[R,SSY?9YbgL<g;Y/3SSC>CV)V7M<K0Bc=K:2+_IHd>Wgg4&cX;^2[5F-E5
I0<Q_;[:,7N,Kg6b&J(C58K5]:MCZ1PbTA[5g.TH2A31ACB=M.+C(VY]FfUa&d92
_,b#g_J+]-(+TSJE2BN1;0a,#=]CA07O[]N?H8b04[T_JVQMF?eV5LOK/JcT.;HP
C6/<#3a\/V/Pb+GW#^F8?W&#B[?U)4cd>Lfg)P&eZ\:NNKV6W,RbSTZ?=1=eU1X]
11_LaUJ[9/&BKA6G_Of:AJ1A\V/6469e<DI_F;/)7<GV_b>&0T>Q2\\]8R#=AV1L
dC=]cZ1)@?eIZ?#Q?RGcS_Y-)J.MN4CVVd@@M[1FMeL:_KCcaebe2]ORCePGG#FK
/,-fNO6Y[YCE@Y+\D18:Ja88<N<WCI_K#PFaC&?Dg<N)Q5<aBX#B76fSQQ&&BT.]
3@3BF-CSH<QZ?10Ha4\:<\6PUE[BbC.YL1f\BbXO01M/+^&g0,.fb6T:MeM:a^GF
K[O\JUSO2:FSLEYBaC+)3AJ\a(H15C^c-S?-V5Yc5.2OYd<21I4TRLV/Y?ZJ7+4W
Y;AeC&&E4&<R?ZE9RC(@AZa2>L3.\\H5#=f9-D9dKD7.Z]<7c=HZ\3NMTHSCS5CD
_IZ]]G6b3#OFR@b1G.NTK7d6Y+6+UN+8>D(aK(>[P/2@QU2L=/NF.:8KP6?;VVMO
NHc\7##M:5+XZa\,AV1>8U^PKY9L0@b#&<gWbO095(V.:V6e>B2:#/8S3b(cJ@+<
d\DK-6gP6Lff&+\?Y_8bGHDE.Q3L^7fDQ;B[HFL)bHZfI4T0&I@RR&c;eO^O4MH,
#[>:ZGAFb6>1C_@&7[2=9U+IgKNV_f-C\+JfA0\e5]<3,]VYMePd1JfV#30GM^S+
]e1\ELX#Y1R1S38<@F?95=S@I@V8>AHARG?A;#)&@A\,a(&UdUGE>1FHVZcGMD/_
aU00YED02&bcK?N/g+?KA,4=b,],WXU291@-(.TTY<CV@La-=DJ+-\SXV8Q#5;RO
@0C4^g6fTfI/:d?S>,=ac;e00A45JN9HUSZ:(>68@,?),\[Rb,D&IfD^c_S;0fN[
e2IA6+=0VK\]KPLF1)W[Q,AZaNH,@2K_-,[QQFDS\\@:A=X>f-P>Q[P@-V4#)M>T
baU^\C]<08fOXVD_1^SadK8>G_09&WYWK1B]55V7U,+QJOL\=g7Ue5=DQBNP?MNS
3E9MF69A.ba5<23LPd0c5g<f>c9M9477-6T4\#A(f)))?_R&KgNP/>Z8>5+a8]98
JS1E&0,bdP=K,HS)T(LUFVb:QSI,[JWaD^LK6F^L1P+2R18R.EE>&61eZZF4Cd_9
YDVIbQ/ILM(?DfG=e5e=OE0L^VT?_I:^(211-+&;8]3:aC-&\:cd:SAOP@&<Z[42
)W,V3XbO[c/@+T/,gQ@VC,A-QQYE1U&TWfV1Ee/]aOdffV:+]6_4@9)1S0.9J,U,
3fdII4SK57I_4(\gFEPaAM)\@+d[AX]IA].8:6JfQ>O@bR7fZHA\364&B8WfC1<M
g\E>:)1IRQ5P15&L)aCYd\8D(<UW.,f;A;^D\/6=ATX/8G^.[8+63W#cTPbVWDc[
/dGBNTO[#e2/=gfg\_N5JBRWCCf^)^6=O(^-AV.I+e.5UFd;@9c^e,d000F;&V7M
ASZ,OSP>OU(+VI@?4P02V#c;J,?-KK>,2P;SL@O<CD@W(B?&gMdC?;V1J3@/e@bA
MU9W>1M9K4>N:9.JYZ0b4#GW5L>/[f@)1DLMW>@WC[_fG;K8)-eUFBD)6>Y8<DFc
ZN=&=JgX:@f8,J:Z@gWGDHNRgUV_#VUX337,\KP68_PKgQ)/_)HR?e:b1FXgO,BL
Od1VGLbWF<]<@f?AT->bD0NR4$
`endprotected
    
`protected
Idg#/AP8SGS/OfI]ONVB3EI\IR\&U=bb0EI>=P(7ZODR6N&J1b,0.)MP8;4>0VO_
+C]aYM:.?dg/.$
`endprotected

//vcs_lic_vip_protect
  `protected
Lb4O>Od;8#M.gYQ-=(9,S_G01-]WA4:<g[MFR1:.Ig(S31/HC2RS,(LPY?La4CB@
SFd6/0FXFJ[;)?^XVV3^YaMM\;2M;R+49:4-0SO+Yeg9X+5AH(S^K?+,f_NXG)G9
N6X3.AaPR41<#X(@eT<2/SIeO.TQ,(6Ifg),IHF>JF6N-]1f=:]8Q-:2c-e0T)K(
6e[^^;Wa4\4P[T@#.a(KdKED=XYE_J@]&\CLT=d5,@M,[@Y2L6A<VG;KVJcJ+&5A
[B<4bMfcMN(;<88Lb,C<H,JEa[@_T-/\\.QO7MdB2@/QE/Z:_d)DYBMNM+I95;FX
34G[#>b8;KOBP@+L;^X7:TKHaGC&TD5IMe@(f]JOB#U-e3<1GdWI6FZg9IaZa=:.
4G>0CM8J7HB25F=Y<6_e/\DRd7.Ta-&J-gLb49>dDb4GU_2U&f^De@La;+7e4B;B
b7e=7f+PBA;GVHX.WCN)K5gIP<84>GZ>T61=[KWbJ#66@B23;YWJFf/51.#VcW@W
[eUTM._??7g]7N5aC@J.5@b5NW^2@gMVeB+X]DE+#W&JfN?I\./QB6C@?IS#1Q>0
dB]Q3LIXeSYSbF(0]O3cf0Z26F_f&V^K5d=Jb=JW]3)Na<#/3,8&]YK5LB3[#VD]
e0TO(KNASE^6D6K6JX5;#3RHZ>4-6FaV)Z5Z&;@A/b92gFFH,>WY&]:]9PW9R#PK
PN6WMIXX9Oa1TQ5,D_.U3R,^Ke&K8E7Q92XcR6Y+6aOLBTbR:>(Y<W/NVE=ZO<,=
QE:If7?=/>J3ZLEQI_X;AZ(d4L(IVTXN#Q8#SG2OQ(REN=T--:]X2U1GW@43?FcC
.8gD5]gWg]_:3NafdIM[ITXT3BgdS1FK(2&=#-KSUc+BB=J^3CG4MBc]&@aRUT-<
;g&((@P7Q:/d(58<g)<f7XG?Xe8^c59PX2)W?g7>T^(I?NaK^_)0M[Ae<E,eH4KP
E(.aS7Z>PIdKZ]=1YUO[B=B_XTY_8dD6Ff#__=>Na4?)L935_Y-IKP@aa8._3J#;
)S@W?;A_<R/GKA^SRKX[,g4M;aDITN]R[<8e74R9;<TSA#9)M=C8>?4?T3EMR</g
^_244_7<F?OdaI9O6<?@^XFg^D9;)?I(be)29G]eW];:e&b+4U_?;SJQ,(gf6Cb]
L;VaY#Y[:?>#A4W7Kd#e3e.5:bMGAK5N,ea=MEc].TTR9_??75SP:,G9BWdK;J1;
)\OF_24\GgAI<=fNFeGcVc69\f[C9I#b1=?PIC7HG5DFN5K_d9?O[(U-JT=3_\Y;
dY4b?J;T(?N=ANTFcCRId_JX@XfAN.SfPGQ])<03:99##ggdVUg51YZQ;AB&E6L[
>bM2WFS?VXYC>U^PE&Gg=-R+fE0U7(,O<:LgMOKbXN^4((#:NWcHK_=#(cDHYU4g
]7WGN,H]YUFfL/7PL?JX9RVW34LO)A/WLPG_1I4fS5?4Y752fT@,;G2\3MV0E79=
a4a9QE3313@SB[bC.&+2K9a2SEQKM.];eUN35f,AdgWX5)3FC);Ef>C^e[E7Lf?A
DVK<bf3+=JAT,.8d1=]M#:^HY#e_<+-@\@O9RfB;#O?eX1^JAO]<:dC?V+P+cC8Q
\^6Lb-=7PIO[SH[dLH_J7H3>0M^:,4Gb6H&YBG4T>DdXf]4X22,cgHQE]4V<+1I&
De:LST5?1:\DA;)^H:?-3543#Z^6&c1EL):]=).;g2HAd_.S\bX8;T27YdM5YF7+
YZI)=LDd:]CT=L,ZJ5O9.T?FbXfOJ+d90aI4S2d\B(J3Ic18)GJ<5TEc_#US&TS,
:V&5PG;9C(QG(/+OIIXL.)JTT&/DQ1#<G=DfM8PN?<+U56V_K-1g&3NM)P5IQ<BD
UJ7VO,0D#[RG=0&Y29R30ecYH_U1EUQ#?0;&032^V8+XC/AdG>98KaX>_@;4A/Lf
CZK;/=0(G^;G6:J,&]OS^NOHD2JR#,a(e?B1+ZF&9a4X(GZFV6Rd,_@eRSQZ>G0-
O:@RU_12WEX;10FOSY3RA<C0S9D)#cWe))Z/I_VeA\WP@\T>(>[QaGXR2/TS]f+S
W8Z@-/:>:fKU1O+[e48K8c04f:HG.L.8BKLb&AGJPB7a&)FWZJJ8bZO9<MY/<L;X
)405U5WeO8R(aKG@92bLf>B-5.U7IgXR2WB?YDW03<+aTSZAcWV#5?):DLT&+N=e
ScZbJKPXE)Q?\64)_1JL7J<RY#K.N5S0_.4+CQ.(8gG\J/OLNE:3RAaI>a;[>g-b
PM^8UK5].#?fGA9a.<>H<G;K<fV&Ra(FT^g-VE#OSI&MPY&DS#DZ1+F&OC#cD3DW
D?:ceXZ7]AA7d8]]6#XAMId9@P,e4)f)W66/U?=^DN#-W)dXD]CM#_&LTK@;_(J[
KJ);G:bTG5?BfE<->AC/V\\/U=<BODNH)]+7cW@a_CEE,D/7X;JYI4f&4aX11SRD
)_787>6Z;#\cWcYA0#eZPO5VY,:+5W1ZC-]fYF.G@683YeW=YWEANDg<-5&VXMb?
bP]8.MY<8^.#Y>L5>B@g(H1HgdOB9HP9?e[?-X:9bS=2OIJA#9F^X&=9\(4BC:\9
bPB<=_2UKI8CM?gD^e3]@J^C)[9N[b+G)>?<\3S[OOW?76_&2GMU@CJ/41B+PNdL
c9)ec5dFU#E-b;RcO:26(3b((KNXB<7G0H/d]1Ge[;&@a^Q;eOa,?F;cIV>K>(V/
9F9=#&;4[;#A61>+>1\VWFL3\<;eXR#^@2^gb@b)4T@/IL,X7HG>U-Z81PaL810+
-,31AUe4,eN4E4XLeZW]b7]ZaA6:NXY5e<\Na<NI(J0,//.6U^^^Yf3VMP:UOUHL
&WAe#SaMJ2&O@\(bQ73:V,C<&8(E1T?JQ0E1&KbGVCGHV[7(+TA\YcK]&)T\7fFS
RbDdX;2Qe<C:XfbUY.;WE<gd9G[@OTG&Z&Tb(@/&T)^gQc3fM?I2=.>O#U&3]9X_
,adC33.)\PA1:5A</,cJ#.C1\ZKSOL+McgJAZN3X2.U&EFWR+P]9]&D6W5M[LPLY
WVT7XY@&C2X#)YgT1A25@F0G?/_&1eW08S9T1V/&(fCV?bP#?8^GIgR?-^CRNM75
)Y(W/=KIf:1VGU/PQ,XA;)e#b_5RM#[((NLXa/MMD36KUfM6/NM4fLJ&+9+G^B)1
cO+?(=NdF1N#@9R+4\X2dM;OU9=(?T-C<J;AFY4YOWIV/70cVZCA6N&8^2H)>ON.
EMC0;&_:a)R\];\>]_/EJK7ec6STY8H[c,X1XJ>GYcWegSY_C#N<U[/3W/D8MVZg
1=G6Y/+-[^Mg/)Xa&8b6,C\8/T<^C_4Keg,0;QY^F:O?fZc=cD_[H]/67ACA<^Jb
WZS9U&=\:]C6?3.GcBKWMP^3GCY@=A8ZN&RDFFVW6X1BAcL.eHO=93G,HY31+E?,
;WeKdIeJPJf&PO+=<P8Sa+ZE(1V(OR+ge+GG##WLWf/B\DMCO:Q#ZI&_=Z-Qf&5b
gOc@2cXWX.-PJ)RZNL<)D<+c:B[8D49=5.59LU.IGcDL9dEC==NaJ(+YETb/>F.G
[3aJ>@-c_WUdT<P,WXIF/KOL?9ED8-A@fI<fCF3J6ZeAf8?R/gUNdZUbK)@8@VKD
KX>-@#Da&GQ()NRZ?IVXQ_242\AMIE7<WaAS4PT.CFYFLcXQC:\:(#NCXabQK<IP
B<OD3@Qe4S[O?M-GRT_M=?E8?69&Cc^[fNPe_Yg1_O<G]O7F-Qb?,gSeE=P4.c](
;+_)-,AA</_E>FJN;QW>S_;-VS>F.19fZ9#Ae@>;adJBA@eD?4Q&Z0FAMXbgKZ).
=Y:Na+;K9EMO+dXe5#:M,JP1N8+C@.@0:+W\.&F\1[#2UY7Aaf@YD;P<-@7)N7PD
J8RQZ)-P=F<0A@?;L094-?;28B/CdXS\[#_#;O9#DCP=F]IH\D^R=gL,H]&b:g?@
=-]_Y+McH67,cRV=]EV0?#?PQH-QB#\TdSYEKT3?3V:=^PA\[I4,c_KA=0N=MXfg
?_C2G/4EAUWg<@c3CL76DW/CffS=4O.J&1T(O7@A\H?g7E\GAQS7MOQOX\A_WcR9
Q=+NG7ZOIe&76WXLc8Y,],U,R:g:eg.SdY/7^(<V_IY9Ne8L:M&?ag>@4X-OA<?V
G^I6ZEb7bW+EFJ3e?8;ILW9#Wb/1DL+(^cb\(.g-=44]#D:g1G>+9A)5(gLL\QeD
R93]MASX^_)SBDUfa@1/d7SaZ3\]N9GRS^YHCX=ID:c3(J#/e37f_e3e-V>36C^4
T>B:IFf9)TOT7/E,RIH7bU+cHOZ^A^IA5?3(9=K(I&C>PH4Hd&[^2_c\f_,E[[)_
<;^]dI.S3TWY3L-dGMG?A_>4K.ad[.Ze\@2U07F<C:]5]aZP&(E-OeIJ1&H>>C_d
-AgEZbC^]B?d<F?:E+E&G84f-D[/ZEP)ef5fJZP6Y@D=W.BI:0)E:B]#+7<^6T]R
JS8\8bL)e,Ef;EKZ\.gCH_MXF2MWPU@O&/:_/X^bXJ@d2+G\VW/SOJT)@,TPRSEP
>;]DSRPEP3TaVf;WI;GQDTZ)Td5LV)I^+[0bSV)O_B>X@Jd93b/T3W-RE+fg?AN8
,=+^NZX,(O)_g@U<B\2=93cfP8=KWABUUQ#;eMa@7/:dJdSb+^7g#.EdFCAWAWUg
MFJ+)4@MR\PUKLa6]19H)S\=L=8E1>e\Pf:@,gG5:83EEG17C0A::[-1<g4Y=-T.
dd)IBAJNXZI?<PAC0DY]8?eVOaZEdR@e7+)U,_UN@2;@(EGHA;X/]9U<d=,b)SK]
,_:E4^95NSW0BHg0KQQ]P6LBDPFPP[cgOX8P4_YV_DfAg.KCB9]DC00Y\[VI_g)C
7;XQE9WD7LN^B/_9;3=+H3HBWEZ-6(<f3Y^<(H[N8UD?_S^/2\^&RDUac3+>GV&3
]BfcE(K5@R(XZ?_X2K,S4][+I@J9YX[PSMNUD4SJ8(6#HGBYQV34(f@:+P7.I(W^
0fE\X9C(.=I,KS[:N);&1]/HABgeL]99JU8UWReU8[fL+WZWT1S()XM^U.7YJFOc
>M]=K97<_@)gbdF=2L<7(g8]I6_F8RN)TGg+MQ-AY&C+=A8:#)J.,LSBM_]2<MaI
9b6f\fPRX,4D0>Q\&9B7^A9a^1<UVEX4S9R)b4-7,L8GNa2M5e26QB:)UBM##<7V
-cWS9F_,=H@@;=7Ee&E?J7V]>4UfL,DL:7F#C(2e2W/-]?W>5Z..8:c4/QZ=:-CA
=IPMH\,2a,924R.W_+H3T<#U8=C&#(Y^,NR:99LXFDHQU:aGQI-65(2C>^7?=Ke]
URU\0E[a.QXBNeLS9fXIUe\7D:<[8/B2INJD];]E0/BFMA)ECK0Y.8H<7#,8HbKE
BC95T.(#\JeEOZEQS<8ZV_5C4GQd-11UKF2cV]-A3F:aSd,&[:8+)R4P94IY[CWg
_>52AMZ#E65b=D8WG?1Y2D=e+6_4I25;=R_T:ZU>?NKeO20A_T#^\WR4+g^M.#&f
fG,.3&-TL94L-\P.6Ke1VA?6.PDLWeHIeYbAHK9bJeN?Sb9#45]MPHIS4D3[Z(CH
f,EgX.DC1)G;N(YYc,.Wf@<O.Q?[0=SNB0e.:7LJDSf&4EWI:DYfKefB0H7V-)^8
5&;2MSCX(AIZM@R6^(SR:FA64RJ+X\BU103,ePXYTP1TAWU^XZ-[VCEfHR5884X/
#X^gENVfbP1CM_4Yg,<ELZAZ=T&JCJDO=]NT(M-4M0N6;6[AU+cW8a24#dH=e(UU
HUK_g<A:0(#2AO5,U7cG-c;7FDDK3(M&0H+:8+0&<J7205(=@>b;gSNA2&FR;g?A
24S,(&T,>=MA17XMc+DWY9G@,^cbL^6/;D+,37T;@R9,9]f1Z4HKSF;=ddDU1_I:
CK4N.RG=(E5[+.@+[47R>Y8UC+^3MO1A)/A9/-QaD?Fg^,F5^,\E=P#K.KD?=RD2
T;E)OgJFTXH\GYP#IRAGY-aICd&E>&?0@,eRFcBa>A,b]E<^HE->4YWG\41<I771
BUO_gb+<X&MUaaLd;7-&\Tg&K46_=@.P4\,:fGRg=B)S2J2/J8Z-g/H&G+V-HaZ#
e[/MQK30>8eg@cI+[4&20GSQ#K86-_4e,Z8?=21(HA805U+KO>5eL@A0>7Mcbg)I
A+0LPMB;dWcbP&3,&?KI])1[fC:GDZ@bV=53(e-4Sf1MA&GEb0X>75-cK8VU]_(/
QLM5,9--@T@I8KAKR8Z+VdPHa)cK5OVfdG(-_C@K@;6:d>JH<][P43A3b-=QX,E7
93=KfObBK+TQDX^^1+YL2IeUHa>+>4K/6)1(Y\DU5K=.TCJI+aSSMGe:RCILKb^:
JMJ_^1aJ-?A=EDX[1_YX>#g14OV_B@ZOdKR<[5f:B1I=N;NEHPDbaL77EF:-6&Q9
/&C8M6T/@EY/?\><CdEOYd0KX.PKeQCK,6eZD0X>M>3\c)fD--K78f=c-:TBA8-C
_aZ=S2CBb4VI#;J<Ng2a^6<XH>Z@c_?:])D0)2@\d^IXg+HY;+2&;GdOgc.Z/B1#
>[5F(5g4Rb:\de>9HY#,;_O0J.aYWbZ^7U81-PHU=Mf1+.3aO48?Y<_<3c)0TeJd
S(SQcd&7d3#^66U-HVa>.8)A6)#]K?_PEObcV44<N@#B&)D+;@J=d=G)L<d.8SfL
L-.4?F=HCF?@-5E)C6:0PVREFKdg6+,+[T@_-EP^<Dd501F?[fIfP1d/F14DOfG^
A2R;@L<2#g8;A<FEM1e4]=M0VE?b+0LS&f@D3):d>;VT\.5RMN_FQXX:5^^,Q#1<
A+&R&4A)728.5:/CN;_3OKfgXce+DBX_bM]5.(/3VP,RbK&XC/F@X\9K?8#7-JQT
U\?JKe5D;,XNcX&I+(ce5KA/>+ZBXY<->KIN[J+04aa/,>K6dfG?f#0=C.GVK:cS
fELC?AHS1D/0?MN/]Cc4KN4@YCF/,+]gEY\R4]=ba-a]&=Q7L+1&=&:+HJ)@^dI5
b=<Y9baF7V7>?@-EBCX4W/e8XcNL[O[=eK^YPD\7fZ11J>.PCG+b0C?+/<65/?(N
W++A_+fI.dRg)TOHNdS9^@VP33L(D>O82PRc49#?2d>V00=OD#D@2d4YB4P>8g&F
XRe?#BS8W,S6a(C8&W-dQ663\:NJ_GBB:(dN0B_>[g0Y)I93fT.-:W,Q9/aOD4([
N88OXE81LIHR#IeK^S<eX<g=NT]gTWGGOK&22OdCTQ),gL7793V.M[&f1.BKK>^_
Y=PB79)0X8^#MN7B8&]S/c8baBg?2\SG,M/(V?0?5B#3/YA2PNF?b(&d[@<V6WgN
F+Q/?[??7DM5K;g;;3eOQ+2?H&;@A20?afBd,Qc8&Jd((GW?XCNg?8,/^0b5^K41
e0>9H(M6C]2CC:BebHT+:IV@II7.5[;P(/IMaG-[g#]@1(SR@UX^4CZ3&VMZ,^aZ
9[bB6&[:>/dgOSMI;U0S=LFXEX4a]8@?P/NU[Y)<1AZF^[]W21Mg#Y,)<M-/>4K(
E4fUTW4>Ed5-8A+6,/&Ze#8(R0\,WdB9AU-;NaINAQdL4aM<+Ib74>cO66d;H\aQ
5;UHS?5&QP&g+W:+g4_\1Z:Z.IZ:PN-]K73JRfZUPZ6TZT(O/EGW<KOAgG7)1ZC/
#64G]&_<>0,:cP5W4g@Za/3gc.cRcWfYcOTIBdQE,=3)BMY3g,7[2?gaPO]D+/0G
RP2eJ^Nc2H]Sd9=:J[F\CYQ^MOB#B>aaQH5R&><LAeG0F69F2f?/Y+VB[>N?_E^F
[&]FQG/+T[G1>E,fINW_ccNRaTO;:1ZYN3:HYJE+T,[aJ>daG[=5(DTK(?[(-V&(
?R3bHY5J(4<b#Ogd5XVUY)33G0GA6.c-cGR_JF)MW#R.+@=0G^D[(595JfS:U0=C
XPeY+-+YbH/]O?8H&YLX2d^@&<U;-S>##Q1,-RG68P,U@NYP(UcePB.&7gd#UVg<
UM??5>W1)e3L,</9b8UMUXCb\^WA>(43[c2Z+TAf].5.XINU@Bd:]19AYKaWSTF2
4G,)+E,/^5e3+T9FSZ:/2J:S:]3A]G\.^RD=S39PcH<#_Q>;\]03()52WK:Me6Ga
_6OUB(E&D1G5P-K[H6P\9dFF6U]N/N6)Gf_&@U?H?C\bR5S<,Na8ePL^UKK#GMHa
HVQL1fA,D?)QUW=-?8c)HJLFB:]V\1K6@UAM&:)938;A0H+QH[Z=0e36[bU,2Rc>
6._Z&g9fR.]/J_=;?d[(6.7]\S[U0AM8GB&>\ID\?N.2NBf2SC]:US1X]d+9\QbI
JXGUYZH>PX4:)f?0B5Q0Lf?C;I1:;Y8BQT8FS-BYHRFaVC_2OK_G8][9.<dTR>(_
Z]AE=cB.M;Ae5B(3L@E<XON#U.XV:0PGKN5Q>3MI_OYUJA\7[7@<Z#ZQfJgCPA,?
9C;>??\(GP^2ZE(Q4Dc8^UY1E4.0=CITJP;@+N(:/HRGU55DYQ05=K@7BG[B&0)L
e0bOTQ&/BX^\,KCECE,Iefe6gaf7<PUZ#(Y[&=YG[^_^\9<M]YG?>INE#U8]G6EU
C52::0gDQF;UK0R\W/Q1;5g2WQA3K?FOEE5.=56MRYeR9&HO)d<&2geI\6J[QA6I
R;\=OQ^-RG-ZgcD0Pe@8.EJT)[WHdSA(11_W>gL<J-3_0)bG.68.Z)44e+>PNFL@
<3Z<FLDNNBG0:IV@]SRMfN.g8VD[UF[,D2O)VUU1cb7Q30FBW6)T+3TB)Z<6)ZQG
B;\dYHJH7cfEFEccO\U80>ZV=9OTe;8L#O8.O568b\33fTcL&U^7aGW26JZ[J-_&
Z-K6.)8]#]9/MHT0e5FgRXWWIA\7\DUbdLISJ;@(3DWU[J#LNY]MZQV<7XI2)9Kg
39,35bJ6a+4g,e)gO\gDXa<eZ7;\bH[LZ(4:8@99b-HdA(CcM\BAcg\_H.7feXB2
P#7;P+5Q:RUY6AdI/@77VV?3O..3XV+&N.,cHV7,-U(??)\F^XV.9EfJ9b@,D9d0
.=Z25U\3W242]c2B#Ne;1?V@EM6fU<_;#LaL4A#Fb+[POH[:1OL)Y=a?1Q?TG\D;
]X-&H-D?]a].GDcg-4+.;_&V1_]38.bF(9adJee5;d,?/A0S]7BAM-g44H]+b,F;
dDQ&YaD?e_Jc&>5A_=RT,-9AUb9BaI<DUIg@Y?MV\I,F9^T^Kgeb.22PbR)HR?.Q
[O6(8?Jd?4(5S\?R[(1<=2O8gdfN<L;YNXS,=;0DA;<<^1MEd1J(PILAcHgQGbL\
b/++9Ig=#,K0.;@g2Y)>4+\3Hg4S9)2fY)N#1&EFBCZE;d^24d,</0[L5Z,WZ(B2
>Z[R-cMB9:,@B7JF_P(Hc\&.+AMHD8f&dc55[6b45YE;F&)7V[1YQ853)8Hc1JIE
bHMA)L6?XP=\KK^bTf7,2S.)I&E\?f9#3f&02B7GIe^RY=#O^/(L7=V,ZD<5NL1>
/+]DRS6C=A6B/\,.PN-,T]g7<;9Bd,R0=d\+6+4Ac7aG7fS9P\aX)5Sgb49HJF)@
]Q3_?\eL)<42d+BH.:Y9WC(9&0-RGfe0UVF)aW8F7#J4>>V9/beAW73Gc/VWf;5H
)0)J<P=,8EcbXEO;8>#g5GT^KedM@XNI^BS,G(/Wa3a8.9BU@YU>GDAQF.Q\MGPc
ZF=+]#d8-;D<U.\]J,LTALeT48(2ZCRB]:?ZRfZ0W>\;,IC;7?5Q4_.K8g0G3KU-
BBJQLR(eOPb/_DL8F9(BTZd=?O,aN)CP>6(F&:MUTOgK@#DE=ffRKA7,S+KO_b.?
[If9Pc;K.Rgb^K2M1c>7Q]?fGR=@MBDgT873YA;fgEQTFV#g&6dXH2+c4>.C/-2@
,2N5S6ea/RG,[HU1(8RN2:FJ>?-RW^fX\IAEY/-?D32?C;5EU@VQEXBA_Zf=b83O
^<3(&(0c]a:9W<@e3,P0UC4)X[7+W#5-fMV,-H4I^d,(AVf/:Kd?#@&7R]8#5d.,
X//UcOfgRc[X.<I7GHQK=,N0HI\-88Wc=-ed^YgLV3\^1T]=3g7Jb3?HgZ@V3#f]
SGU]TAF]3>>9M(Z8JT22Z>[1)N7;H>KD?/JbJf3+d-U^IfQ()_X1=H8QN)CQ@;V6
I,ED59/3W]=60/F_LgGLYcC-+3Xf<@CN-?QcP/cT<D2M:N]eKMNg//QR5EHH-YWX
c4IJc7H)1N0M6FBEIEQAC;8@XPZ5dB]_@fN^^HGOGZKg^?BRZY5-5Ae._II=DDX7
>(KA3VGM+@+[-6(-6ZJb)dg(.?R]f+c@//TVI,&FPU)\TF4Ag7639G4+fX/MLK48
#4@H<#+>+W)NB_,@1.=ZVcKPd]/-bM-_D-=.U(H3A/9WWB2D>ge#+KN[WSYI@RAQ
AOI6I@#B\>KJTP\)F9XN>X0770X\_PECWX.5MM)EX??fO>N4gWZJ,,@f&[C\HRSa
GE>+FK\<Q85>#40LUV<<<1)/&K(D^.;7Z7g).]-YU_2PXA)=7OF9K&:W]EP#DD-c
d\JfZA^eZW7SGaCBe/^@:Z[TICK7g)(4UP4^f:ZTL;3NQQ1S;OYP^bZ0\B,Z5-DA
](+?EMQCa.L-@#C&7991TRcUR.#HNd&^,(KSI+Z6:F7Q[WISA9?F;>2D4<eAHd=I
>)7DPR>MSW0AKSa.9]/XWS&7_=JNc.0dWg\V5^<LY5#fX-QQY9>8O5=C&b/3c\_6
U/SJE;:4R4N1/Tff-[a^H<8;c>\<.PB7Y03)G0IJV_?#@e9TbBKEMeLUbC.MPFTI
G^f39^]LD/]?<cKZ;9YE0BGebFDEM==;afE(VTAcEM,8&I^&@8/FF3bcEB#&faOa
T6ae#T3-.8ZW(OA(<c0Q;-e^\c>TI?R]17f<HRN^<dfE@cM[+=Pg?VAQ4L>^5ZCR
<+>:d,,<>^d1fXW^OK3D\XMUV#]7=GHXP>JW_GBB;Ga#>&,6g@\-gc)Z1/]#Z^g5
ABVf]V[3T_K9]S@6SES:bO7W:D4IKT43X?[X\1;;G\a]HcPEDaNOKd5G3;N./\_R
8dUL6T(S=3Xc#,-O;Q@DY+X4Gc/6+>6R2^&?d:9P8U(HZP7[:UF757M(F^<Y<5Ad
_9&LGS,YMOg2^+LTeVH2]7Fae.Q_cBaU^g^a=N)>aOY2/5g:g9?6N&23AO27<U,O
5#KfIg=DX]DP\88(DUdfKeAB6G^[YHM\e#7QLT+2e5e=eTWYUDLOV2cg3a5Z:4XJ
8eCfH;15]gJ^.?&M[:?I:##D48BR)I&U[Y<TU9M(_(VbdeO?5Y\(7_0B<6]8&ADC
1_ALI]DXR&G2TGAQY0=1Jb3UL0LeYRI)Jd_&;Y>cH]2F,CKE4@b]?JQgYK,O4J]P
KRZgZQONfATW_g-NWJJ,9&^:(=dbRSK/c5fP6TdcW@YeZ4Ug1G#RB9&2bcNT?#)\
UdEND]O)C&5S4>[NPdNTW+(T+5K&Y\1249L+A@Yf+)Z\),LL;\L_40A>()]B>/B6
DbQeJ^8=?YGI[_6a&3<#G[PW^=CG>FTZD@,W:4e7U(5NX#b?QT]K-,)THU?aWaNR
#f<8N:G3<40SM0X^AKKA)IA.B/?.+),fA(L+^HdY:5:d+SHO\Y5Ned]Af[.DKA)E
C-G0a5OY^X@<BPC>(H\IaHMQL1#CR)]G29f/9<8I9B(&8EM5G^BW;Y->F,N987X6
E#2G&HP9cQU82>/@-B,.=aH;JS&N#NR>/9^T7N&Q7ZN>\,GF6MTUbK#?_Sf,LCD5
@b3d99YKQ6N@Hc:)=^NY:.7H=#Of/\UZ=HOUcE:d1F).K+&,/#@E:7WE.&DU[YCF
XG_daM0S/G?)aS:0QgC]]>77#-6ZMLWU=__d>RY9(\POKA9S)?[)([e8_06)HcZ[
A\eG28:GJ(&]_\B,c:E.2KbMER:XML=G/Dfb<8SB9^923XZ=+7XDX;E_cO2dZ3DY
N#P80N+3R#Dd7]KMB^RPJ91O3[R#d5TX,a&:X7X-H2d]ZGe2&4XI,>@f0U^_D-c.
M1e4.J@1L+OJCS]fYC7c]-PM)Q2+J+PI_Q:2CJR:\2<7UO0,MEgaAQF6D&<__HGK
>;GgIW?4=bRDK(>O/)A<Q6</fY(;??\YNb4RP_BdMG=FG?bP/[6:(7H+B;X\EM/&
bO_1G51gb9ZI\=G)e=GE?2C96P33_QGXV-edW6.1DO:fAP^IUIeB4.+.G,Of?M6Y
/-cDER=U=8d,P+:ZZ@7HT\]EL#5-EgZcDD)<_@8[:.@9CR6_\M_+WV.4@1A[4A+T
=,f2:8HQF3_Z.KVU@L2=@HF@A\;fRD]C),OS#RDL.QF#ab[S.fCEA,U^SDa:Y;I:
&+FIKa-3_C,BEE.ZOD@U48>#2Q9H;MYQWWDd3aJgQ6W(f][7SXDS04^VaZ2S):a&
O[)JHbC3G=8c@MXI63C.3U<:6&O[RZS;IH3R.?R(cU7a;9U-RWU/L?[IR?-S1ZS8
.;VUXE?2F&(3/M&0PC>/.SgE[0J#bCg9#N&0IH;b.9P21+Y1[(N+G,fJSPd6Md^[
a;I2Nd3A[I,H^F):d+?^APK3[B=B7:Cg,Laa4F_U-_UMLU@DabIU>0_&M[3+A02<
5Sg784Y9<1\c<M0FC0cFc6I@2FHK=8@<.=PK3eKHT&eSb@IJB+cK^3K/OIKePN;^
,F[?f/_D+bRW^e<#?GJPY7gNK)MgQ#JG2+;GE)+>7YGZ\)GHRa8AP5a1P6[0GCL+
K3U9?OZ>+eJ2NYNZ1ZUa]Y&M_U>_Q0K6Jf/1TT0@H#_cJ)[)PDS9Q50H=SGLPSEX
gEb/g1E@98]1?7[bRb7V,RQ/6\,ABS;9<U&SfROJ;E?0A)1O=1]RN)IH.D@,22.e
Rg^UVKb>2LVC)J\KcZd/9<>\4ZLN:MZWCVbXR,;6:YH16:CNT@A6DB\/aVWc83H2
#INfP/S)OX#c1\K4#.RU>FL>V_5+f]0R\d&-OCaJB>(59O>g.+B9&SfgZ[.7_ZIY
KWI.3A:b[c+72,>FPQ?\bg3:@5#M1R;Y7LIe2&fVF(5G9Mf^E8VOV/6a2_XZ0)5,
>eG>c?U-V7dXM0>4LL-7K7HSQ9+I@=fVU(91HVbYK6bL.:aM(-TF&P(Z&?3;..bB
\SdOC^L?][F2GDM6#9.5Z,C7a+0@VWXB,NTdAWA[MN_DV9e8e7/6a?gN8gGa\dZ@
I=agFQ,VE1V\_^@?OB_cZA&1D-GRVMZ65A\<:/C]=RZF[eD)V0F\5/e+NAbd&_J[
&:Od/EV.cP0;P:W/aBWcc(TYE#ZRCQfG)187BVQ7:?Dd:7&fD]<g</FO4(YP)bgT
Q]ALa&&f(,0;5D572Z.>WggbHEUP2]+<&#_X0EdZXc>^]a.J(?YVD3<MdS@J)V9?
LE#;2]JLR/;6cT[d)?56YEKBdEX7B6aFOZH,)SG8EaQ3M6KEBXF</-:\6VZae\;8
gaGUOeT0<PfP)L_5e]Ab?Z.)2\C?)73P&.KRgbHS/A7+U(B++&&XN3&A;Ya5^9B=
ZX:(GeSF824O9fRf7bY6<[:H?g-4.T5QR_JaN+CG\geS+e.JSSZ@/\Y#\<-V\-/9
/Uf<KRQA(DPM8#DbII4Q68cVE/a=YE<[4)HO_[N0.0)=fcE7C,gG/dQ9dNJ]G(SZ
50C0HO>X/T<)XGbRaf^-OU.@,/@J;]]bWG(J)-1#.+HPOYE4B@3f]+L]PaMACPdK
@2b]<01J5<&QWecEb9R.Q[;a2&@Na)+\.>Q)NgRR_/]4\^,Bg:UFI?/XfbWN0+N:
Y4WVAB>c:S]]=(;b70[4UP9=C^KMSKHKe7WBJ(M^UA5<JTbId0ReP]HZ-&Y_GWS/
3O#TW(8FF]SIa?cF&&&)B4?Z/<e_)6>X#=Z]PQ]B;A-CRLRS;Ea@46eEFGYJDXfM
GFM)?fI[]SKK0C@PX;fGG=cVcU;a>;IJZ&3RBY:#QG^SM5NH=?+/eS4\3N\\>-K\
3VUOU8SQH.<SDbY>G6\]<^>;-+>R]#]0DgTHY(OWPN79\F=BNJT\CQdg<#OHWB#O
b[5:cW=EG<>=gCU]\KgY:,,B;/8OF/a^MBffG?4gR;KGTYc&QgS^XQB8ELfO:L\D
&H8-dQd>#&gI?C/?1\^9N#eYQ=TId<Jf5PY&NAbUCCO4e30V1J?M7T:&d#L)&.\Q
O?0EOUZ3<0]+T)^c,X/WB8100/HMKW-c&f[9V]GN^.)_g?MF&]?:3W,fgf=JC=8V
1g)LMOJVJHe<-H@<:\GOLXa9QCT=V.#;dLQ-Nd:BPKJ=4)C7^.1/:FP@[]RPe]K^
acQfF8<V6U;5F,3Q8FB:DNe=]f+PBeQ6^]^b>B;FfTLM^<S+6F:@4c@]#.VW6DO)
d_6^fY1O=G4T;7_Of_;O6]1GEfTCL[HX8C:?:3/H7#SUY)\E_+\f#9.UV-UcWZVT
W>-&fZ)b+25BE)>AW;PNOYAXbYOBc_1df(1:2(M2+)g(.MgJ]>DI]#gJ1?-7fQRb
VD6#80EgOf]I)dEF/W&_<S(V,g=Y()/bfg4]eFQP55W,?A+QZg^2dZT8^2aY+R_U
KS[V,.YIL^(XVYZ=_eDO\?A:2O3:];47e&e,d4U#>eI9YC@W-/68=FP5=?ff^>GB
W_@?U:MR@L.-V))3<,3Q;c=;DYceA^&fM\AFX59Z\.QaK(C3M[5=?YdE+c]QTS_7
g9bR++K.TKQIb?&GH/@,2=G^g78ICWO+d3c4/cfPY40&YZ:2EGf;6CTd:ZBB@bVO
,eS[GFNF+6[cC#9:Q)b?>_A;d?2+HEMA:8O<-N@DE&N,MVBLPf?1YQ&a2Rdb(#TC
a.K4#OV<UXYHfKK+dNH<#UcHY](/0I0aV#eI;ZT_F.3cKI?&a;]1KaLdQTCD?&f:
&69H:@^RJc]dd4GedaHYU1;1@R5adDNdJ_77L/I<2VK9dS0XE/(OYOFe[/)6,Y@+
WGS.-@8Y(J0:?=ZYW+OBIPR]Y/.fYL\C5(GW2O4-BA>UAW;XU)bYdF1:A74Kf[AZ
cde6Z\/#&INUPdZ_K\D(#?eUQJPB>@]_eWPS;F@)^WGFI[,=D76&&YN(D.3ZGC<<
_e]Cg2^D[[G(,BXXgV5d7PT7(eb<CIff?b,Q16)]d+B&RD)D8eF5O1c22<e8NN+1
3[FU\14\a^UFL]dFT.@c1GAdR>&bLAF1I(RABO\]T>[#V)2:(W28DZ15Q:#=f-_P
TVbIE(354X-Z1,4:-^a670+JJD(BJA/@-b/7S+eBO=W-abA:8WC6950@(RE3R&3\
7<-)Q9\N/]@2&_UB[S7/7,DQQbFQ46eM\-YM#Tg_PN6L(?bL4<4HDWSBcB48KcQb
NOfJSFZY(B9fM3/AgWTdKWJFbUfb(JNXU?FG#M(FF2B,;#.8?F/D=PQ0LTE@O#F1
Z0R@Qg\<^4\^#eXW6eN?8[PYRVGG,&6Yc_3SBK)-MC1L[[-/G1&BFD/WS=[.C&:a
E3+G>=+3;aV@\-+e_/Of,[CX_T6MVSbR2,Z&\65]VbW\K&f9=Y?1)TW#@NbEV)N-
>[HBZQ1\SAG6aN[V9Ba]Uec;#9f4#e=4][T:Rg@HSYGM5UQBWEg8P-9dL:ZM1>JD
W\U27,QHVOP5/)1Z_XaQ8M185I72,f2<b\Q>K#(JGKTMFS;LI3L8?6eR\(_^b;#)
#W]fMY,77)+DA3gg@(_YdV&V,VSa5KP_:XUWBH,7>UE[8<aFXZLV?ec<5TMG-V&c
9cZD=,>19LS5NLVE^4YD3UP0\7/<KH\(22J7ABV?=57QT,eHGF(6/GYOQRV=0^M+
^[KZK4O3\M\A0f-.+_@1f4Y3Ec5C)<0<1Y,+:1O(fZ+/4eMeH;BRNAbH&V92-0S\
bS^V0BdHZ82OS3)LbgCDNfN?EQ/XWcOf.R3UCFdLL<8D^K5&5@G>DAK7#T3(,,U+
/](aT?:TALYNaXZXZYTI)GOX-Z)Vf0:Q1O)bP1+bJ4L)QX69?Ug#e?]J>Y,[Yff4
2B,@FGb6VQbU&(&Tc67:7?IGFEKX(BgHTO02,+f&#cEd;GC56e[_DPSI97(gY0[H
XX:#gK3C22E+4a2Y3Q,EZ=-MdW#0[K:L^U67cMEf)^LOOFTRI&>#]1U34@8--#8\
E@f\]/8)FO^]>DY:=[?UF7J74DCU84a^R(\L(a7TLA=,26OOeLg8I]L=UaD<3C+g
WLR\.;eccW?\#O+<<d>(@Y(a-J\CKL#0GP7E,.YYL03@.X.4Q:)3F3&-S.49.?B=
#c^.CS1Hf<g-5IFVF/1IY3(bU_?.E:,dQd#6ZC53UYcC&L8;1D0,+I[G7W43YD\P
EE36>?=&=SCR313ID1dLL6WX4C0HULbN=RSfMb4#fJ2VXWDG+QC>ce23>>E4LHFc
7,PI<[]J]W;E,b,G^6[LX(-NO@9RU]YJ_]A1eU^G@)L-+\@?bWZ+]a.R2GC?A8a]
>c1.CUXT/HA/DCO_@78]#D_1PJW0XZ^NH\^:3_ZF05T5046PF;U-D1dMI-@6=f4^
VAVKH&T47^+c78=[R02:TX2T(1A?QY;(>YF>TPWe&2]N,^,@22=Ra,<Lb\>f>OfT
L&<CJ-&PJ;^2D(/LNE&5@KVeK@8GSTYD8#Nc(N,JcGA060fFD\K^T+(/)2RW3<eP
f1fQcbAe4X2GHWd6W)@>4\(9]&g=,<BWFcV_73fS5EQ/RS38>e,-&WOX7DD1OAY^
@GW4b9[NR+(/1^cP15:<KMJYJKd[VF\&96MSd;^^F0DSg2J=<f5YAGMZ@W+?G9RL
Pc8/b&e+-YNB2IH_J;:JL^]DDEOb6LW3Q<Y@S?faegB=>CC-]]#b>@a(DER0:=Z9
.aPCJ6e&FR:B>;V<.ZdG(E]1(N^ca0)+>UMIKM/.(@FeVUGB1X/:XdT=@U7WFc_\
ZD_<B1I\4OO.7HTZ:?ebc,@\,]@NK;4O#G5fbBG\>W?JaJ;U:EB9)TH+W=TJf8/C
Y2APgJ5S,da;DL&U]LVFQAU>^cddc9W=0&7<R\=TF]9?KDXbK@)fb0_B>/R^<-SF
EEcMYN1-<ACKGN9C1V(U-8aNOQG-2DE_F(JBXZ>LZN<4Pa)Z3FUXUQ0THXe)ae2#
+S=49JR8K0+811345H<C.(V>B&;2a.&_[RGCM9X=_4W(C]4:P:UIK;[eG2J@)T1Z
W:Z6:.<9;D(1fAQb-4bMY[AC8,)77).6@\B#\dV/-:J[Q27A.cC?^_H7N<BZ+7N]
:KE5/6WW15XXS_AUW^]X49Y@^@XQ;RDTG+K;LaKV+,=/H&_/^_aLH?767,WLT1IP
S)305+9D7H=9V<A1NU_S,B9,3;<=;JQG9^cG//OQM]D#&Af@e\^>HB?-X3AKE_WD
,QFR=8A+8U0N_NOV__T(Z(f>fS=CTg?;I0D.bP@NEZe6/+FD@aRJ7_8OOKD#6I,f
(^d[_7>UL)Fa@K>AXfeTE?Y?;Leb)WE03=)c0(058\I)2d5POfBgNN\ENS1_QNZ;
g]SRNI6eL>(MFL+-\=D/N;H4A6P4-R?K6U7/a)QS#A5gA6[/BcBGb-17:^UKdT4:
I,Zf_d3=:Pg>3LeJHeC;YaS\PHK]>/NbHfgb<@]@e)2:LcGS(8Ca=e]#>Jf[(9L+
\NG4M<Dg29T)c::.MQ=SZ8[<#1)RAWF:/&La9&-([?U?ZU>4QBPJG\fNdPP0SWPS
L&]^I=S]3I:bPcCI>[>VgE<<&++3MaU.fUAf&1dH<O21SXYH(>52@6MEa@O6gYeB
,7]D?a?daX>bDFW8D/aM)_R-c>@=EPSS)8Q+R.dLJLdN7ARa:U;06-)5Ka1C)NW;
&(UaY:4_b,c#e^8LL>U#2f&+:,-O#L8e5>Y)8A2:P9P)JW@^1C(OYD3CZ]+K-?GI
0aB7]c1<ULIRQJJMDR=]+9QL#HBXR5Y=>_,.UCT_LM_@<cVPVRgP60GR6<)Xg]_A
>GRb#?-QYM\0O7--DF5MPN?S2BNeZ,,9RCY4?Zc4gH5F/)ZX5dRDJ:3CScA^D0U\
_Tg(YMZ9Y7H,e\;+YYX,)?(4NOR0DRcQ1b_Q3faC&YDPKH0-(>aM@>.(T1c_DJOF
\FT473X4GU\UQA6Lf-5-BaY+E3Ea@^JB=fG[GD?R_)B>E<QU9DgCXPP0CK\F+<8=
/4C(+R0F3=2e],FBU4N7ET@\3YN5g6UCbFL><430VI4b5gO/3IN^HU1Y-0(IU2H4
0cc,VNDf/HE\H8bF#@2bNg#??OB/L,WUY0/31Q6\])?84F[DL]W?Be9:dePMgf0L
[:fTNT6P#N4M5>Xe15G.OY)ea-4HY75NTF@1SAK2&.7QP&d;gdPIQ;#f?@5=H#/K
cN(;[?>)&40gCB+?b)0<Ib.La8V#+?/-F[^Mcc^>f<JEO75G.P1g;(+A2cB-DI#.
dbE8L#6L4UDSgBWEG2)=A)=[-HGTUZMZ,X758EQ@67PZS?e#(VeJ].D4NN(cBK>M
g9M]:NYaE[N?c(O/CW0VTc+Z87]Lg186/2J]>9R3[,Z(Z/Ld7LL^[<T-:Sd:EB/,
WVd;ZSa=&GPGf#59-U1#cf&cJ&S-(f<YL1CH9QYE7g[#[F@2SUMMRKYg_&(H)=5A
CE#+5\+FXV7Y_U^]CX5=[f_>SN@7aMH<.:T(=?g^UW8K/_;65X@P145=,[/I=(fD
1>_#[@)>U,3/:^CLTQBgJJGJ[4c=2_22C40SAA7<-KOYgTWeFP=AIA65PV6YN^TB
_(W<77[>^K,<N6SQI3^M9]T6X,/0/&Q#Q=OWCMXe\fC]1TG+DUBRBI^9<C^_N4dF
);2B7880#d=g9J0[0]W?E2EYEVX6Xa^?4J:(eXBb&K3^O7A5dY<(1+HV9/?E3]0d
I2#]\_fe2T(U&B^27Id[&cD/D&TVYT.@&f4BZ<0IV67C7?JD?EUcF-K@O?-=eP_/
)Ke9^.PS:;\W(.N><\\&CCX;d6.UY9R<(FIUc3]RWc<PH\U+5ReWEGFYX8Wa)\:L
,cP8=#[>#T[C/&=6=(:I-=[b95dbCBM;5AE/>0:(UQ2c=9Fe#P#.ALB>Dd&J+)6G
(-2/>MMJ@U>OV4LR5@T#g75=2ZKR#3+bd5FQ@:H?RN<bR6T9])(F0HOXU_:<U@L)
)1ggb1DNP85UX@0K=</1<^cO5La17WY#a;3374db4^X[>VQOQ;QX8d#07T-@V&)3
+]edN7YPc.&#B@27G#Nd[5Ld)B>a?-59>0CZZ46\WeR4AFH0VACAV)R;Z9#5PcI-
@X/)T6+P6YX.:b6<9#Y6[L__+@HSL#aO_,R7_UBXA?B-N)T[<>0g-P(1;[B,&9BR
(P>FM^#Gf)G,WY?fOKTHR5D,cLTFW\#fdF@;.W0LTNK>2fW>NVHXFQGD@c,[V79O
d2W8EOIPa>P,-]6&?#T>@Y7N,c_SQ4+=.0^c85D^40>@J>J:/OTEg-O7JP]TRS68
+(B63CDJ=J<,E6^>89Bg3&U#>g0_2]T1G^RFdSX1V8H0T=.aFa?)4F?HbfUI21^<
=[.#-:,6.1^aAJ-?X88([QcVF3-KUPEQe/#>WD?_-+f,W[03H0D39XC>1K+EE.1#
<D-SG7J=K&TDg&52S&J=a6cQcaWDDJNNSU7eLEg^R[L5PIBcbU)UI1+Mf#09R;;?
K[f8Ma\@Tc3WXEYdFa\NW-]=\d=O[CT[W>;>(b_aKXWTSR5a5KN,ZAUAFRB(BYdJ
XT&6.H@JT<GR\<Lf2QVN9E6EC+P_X>:=7_U5MEFd=bHI1D,V;Y/6Q25A?5]U7,W^
L?YFa17(C90(>G0@SVV4.?C^TL;L8@RG@NIZWKO#&C^V=RIa]gN+NGb5^J-,#E;K
g5JeY0_cGWYD^9S.)ZecU#Ka3Ug_.8F5>S4OA<(_eQ/&7)S;f3H9Q/?Ce#HFER/-
;92<;.WW]ASEa^4cK-GUE:ee?W1#<GdDN^5aZIJgdP]H0K;N^8KDO5?H:dX[[:IC
eT[GKLQ/R/<S][E7+DXb6<FCF75@Gc@^36:CfdE4BcU9HKYZBZZ?4?-[/.3W<#e;
HAZ=B;,I)UPFVJe>H1.6^PeeA_?FA_,T2,&CNg___Mb_OF0M.3518)RNAV456AX:
N\^L_[Vg#aObeWeM]\P;@J3X3JaJ@)e\cU8W^g/N]=dK)^e3I/RKgU1EY1[&/3e3
1]Qe+_97/ZGddBZMHNb@1IAc3C9UE3_I#;S^R7UZ</?<_CaUX(=QVOe4:_c<ZC(^
]KgQU4;5C(O#<4B=QJZ5.=ZG)CF4G-PgM.=M?:>Y<YV4=P\^<^S-9]PM-=c#U2Qg
GcIO,@I,YM,J://aXKCOMKgTSfcO\2#1KIaa@:@10:1SPAO7N8Q4ZV^MeYJ;f0N7
D:A:ZZZ3RRLcKP1bB2^0aK_<NTP]c6?3)C0?[Ia9-@P.Uf74,:)#d;W<>M)5&@XN
M[;A#Z,fXMeg_3UIWB8R-=>#:.HG9(>84DNC<J)E0?N)YJ#JYKL<U-)\^TEIQ-RG
]8OK4^@+da:#FH[K<14T3B1[=FM:<&5G>d/[D47)-e-Q;?-I6fSP)ONETN:-4X<-
C<>1^&[7UEDTAET\[?>@#fBC#9U<a+88:,J@OAKIFXS87,6,SN8AMOK#^[DWG\AM
0Z+X4e&;2+-R8g0T\]R&\W1.\aGP:@Y^R>f7J;W#TdIaVg+:;+?_6^.Va>4-Xc.8
a:1:C,c@7OEI>dNfU<46O1J=<3J6/8G]3#bE-2eeXR>_35MWLQW(CF6VCXWcL(NF
_[,\4@J;c9(612W,8(E5IGGF=^[1(P4gQF1Fg/R6fF=29((0.<L9\J[/&^c&agK>
,_5FJYaWE88EPEa?1N\93d(Vf]gdaHa?:/SBLT;^W59BKaVYADX7=&.MIXG1gb&<
EV2]gSD#WIPH8[WPBbYX:ZU,TZb6X3RA/>[U2]M058@G>4TDTLddb72[#eX(3P[V
c@f&WCCd6PEGUUd7eDI8fI852G9+CW<6#OcX6YbIA+b?LC^+C04;=MV:?F2LBSU@
eF&7G=&cb3Fe=&^YMf/V=?dBZcZK_MWMQ&[b70g()PQC[]HQ?KNe@#GZN@aE83&c
aM@?7&J>S6LL?:7,6@J/8,8J+c5bI2Of,\<FTQaN.^OaI2g@R&^+ICU\XF;?a\J+
@Y>^,TKfRZLIU>cQ-NDXHcXNDXHX3OIURdA-#6_QJQGSd874>AZ/\@XbT/N&,K+e
-^SNIU4TQY5B=cWRaC:)>Ndg\Z7J/;>NO-HU.38;Nf[g?_J3H>\5HdOE;<I<XM\?
#QV-[M^Hb&_:LWMFLEHF7ZXEV@d@1_@,/0_-S#d2O@[>@E_=6LJ?d8<]7DN^M3IG
CI?7b0+@g+a.)_eAO:K;<]5?@I-)#IY4Z4BBCCKVWUSdT##4,c0#>,6OX)ZI:-32
,724?VefTTJ:4Z8E_XIEfeI?O^^&O4K07=>35;3]/N?JPG2d^/Y,J55ZdcZYWC(e
EYV4f/[aGA(\@VZKIS3g8V@)+IgXI8Se;[<<C.@>fU:/3_VIa+M\e<&[e:)QI+93
YVYaYT)1_=aH8eHQD?Kb+H8\>.C^I<F?.X0BD&X/0#_2U:03)^@d30]#]dg]4&QG
dadCV#]Ke1K2G<4,>#FXb;A==4Pc6V8#DM+=&38#^3W^Z(-6#E3B]a=&\K_L4Bf:
O)eI.C3OZG:&3#0eScd/E#P)W-3+FTLW[EH./WT\fW^(KPM>B]+=T&MD4=U=JXcN
=dLaRUA#6H<Q1fKZ5bIZ-H<+@/@&+ENTGUD5_.b<\L+>FS-:9/R;[VNdNc6[dN<B
DcERLB^7DLXFKK(EC7PXef:4B@BYVc7Hf4[_VR2JA@&)NI.Fg6]B;c[>0RU(M421
=b0LWO(d=[dLV5\P0+@Z1+1M5H<,&O>4W)7WD+J/)GYC#5:_C9^5.,<>;B4Q7?XT
Q1O<(:e@<e\C(8KL<TYM&K8g]9NR5HUH(\8b&4_aO1[JT^I^+fRAA]dSEcK\[2;L
b]05+U>@N=(=&\[X_1)D_f1YDd&_0Gd4;:,/b>3Y_AY21T3I5/BU7JBF<F1C616A
0CAE?-L<0^<33N1IabUa,C=)(fPBKD1edd:#BR0-gAMFgXQ_]&CITFVgX6:LJDI)
/U3A\A+(S&C37]Z>A7dY6=FKOceXf6E^I0:2\5>M\c2=7>)M(=@,\<M#VXJT[ZE[
L,OOW^+YC-bNQ^b:\&SB(:OO,ZE8\)S),c,,<L9/1WFc,&VgGe3-PV0&\FVM5S,+
^CeI&^XVXATMC->Z2YV2;31@LPCWK.^2V9V<#HaR@Mf5@c58O)K;V?eA8f6:g&Q>
.5T2>-56X2gIT_W(@M]9HG49g?4C@R;PIUd?Q85^(EAX,ZJ;[bR]8Kf0]B3Mg0+^
Z;d3UGZM9_4@3Q5(-e,57SNAY@-.98Y/cSU&MW>R>G?2Z0e3/R5IJbZd@8#Eb&ME
J?AWN],-E.TL-NN\DfKb1d,EgbI_\0Y[M7)UDPOUb3EV6Y:;>;F&LNdcdeA9ae[T
X0YgFB0+D6BY2-.2821R^KJ\>JWU,aB_R)ZGQ5e,&I9a9BII;>=<T-9[^deU_<[3
G?9SV@bFf7GTLgGL<U=_?4--<L])NR?1>@TcT]NXeQ36@)->^GZHUZCL@UAAE3T2
7Z/Cb-Y6F&.&MB_HW1EaD2RgX)g20RJ^DE6G@?gC2LR).SYSSA^;\WN&6LDGDO19
aEcI+>H]P_=-V92\OJ:77X1cG(L&b,I+LH)caQONc]Sdf]X4R#,?>J,[X1#6Ha[0
7^bJD13V(DO\D<QUX3;12(I[?)RHX30BXETN.KE&&7\A@WbR/)/^-@X8Cb2DR<?J
AB((KG&_FA)e1\;3E55CCfIP6AcZGbD[GgEW0.)]+7=:a:G+4=eeP[6.=CH01+4>
B#R&NO8CI9X6[]&3F-PJGb2QD=4&HLR#&dV3@21:/W[#RIgD@+6g&cW^X<IBZHI6
UO40>b.@-=FN1/3A\[SXGQbZC2S4V;Ab:6AB\>,.,dEYNIIA@Z7=R4.e3TI8FPKV
Ya7EW1D[1D?_JI=)dIU\Kg1:,2(2<=.N?C]<cK3@-SeSJ_QTP,OWbK0763+([G,B
Mf<A90(ee4,^>\5<N<0YOR)V5RMXaDW67SS3T3^L58ddZ51gCQ)e4YFCS&A\D<PD
RL1Ye=b1C8O<](Q--+4D:gd?]>I7:>M/[-L5Aa3D1N4=:0CKFQ>/(T()X\Ne[&c;
?Y\NIV]A<LB[51HUEM[gEf^)TT0C3?5-I9H\(F5(e:.&L?T83aEH_Rg44-8;64).
(6Y^INMOdO_JL#>ODeJ#1g,VI?_AHHGJHI(S=@\a72_;6QYK,Ha9T<4OYGa60ML/
;)S=[WP1D1dEL+(Z_BL_7U3OWG9Yc/=\I5=TI:1\\&A/SQ<6\X[b)#H1T[>9g0M8
>:Ga7/N+cC3[Ye]155VAf>;aU^M+0VB=<&@+e7aNS8>_dSY1I/H5?8C:P)QP#e<[
e,LRP[6CX[E&\#?GMK3]^?I.a,+<=-#RG5g2U\TE@WA<P2_F6Q-_()fA=38Md?HT
LaBMOUR5N0_\e5R8F.FTQ1[4\1&NeE&<F1Fcg\,IX@-gL^#,4I@-+N3;d3DWPaaG
R5)@JK=HBgBc@RTD_.=V:(\M@[9FU.:4<H;^,a+FS>gTTFMX]#NR,JX6>16LadU9
5b[G_6,5EBQ+cgNUO)GT4TY3_V_eF]TEBS;)_)>S,^1SN@g5)b5:XJc&MLB2#XL3
X8C6-A976=/AY,O(RDT+N5R^99.SOf2XWLIZOGE4X?ZY_D(H:<LW@:@H5Tf_C_3I
dEX)8/MK7_OM##G@UL:PC_YTXIH@I\eDFSQ-dWDDBNXB.V#M1[e=Oa)I&613I6R^
[@Qb_M026Oa?R7O)X]^(GOGEcZeP=728afN5a^#O+:9C-2)5MX]9Vb)<:55E]-Z(
K1U9XES9\S@W_<?N>77C-.Rd>g>-M&FX\NJ([)#,HbO30_M]4f<9ZE^gIZ+=R?R7
/6Z.;EQK#dg9V>ZDc53_<TdLKWJOEe+.9d#:P]>=<XO,J><Ve;#H(0gfH#G8EKI\
8TY/M<<R5.<?c],fYf+^;V6.Q.NIeKIWZ=-O(001-VF/\B=B6Mc8IcV6&a)#d:E-
RP)-LZRY/#Ba8a8OH/P4@Y#JSV/-[P4bb6G9I/a^+\](;8.81Hf6T7U<cG8[MU;9
;HCXfM^b)V[^6H>2QC3<B+;RLLc41S<e4)/..12#9;MQ[)I14\;3)16;^1/5?^87
2<VgR5gLS0ec[WYeCP(J+,(NU=d;<<6S,J[._^U&^;NDBH9ZSD(MQ1=1W4V]8X6P
AS.F&fNMM:gbg2.P2B/;Ka9fHAYV+G^F+U,CTMfMZe3)C<8#:e)c9Rc#C<UNS1>@
[TPVL^BM0C7TD5fZJ]8V.a-dOb78MaCd=_TaI3D(6O:a?)EU6WfE666E_1UF2[MN
PJ9Y?1X+VG@38)1TIM)d)DQ0N?66C<UG\Z-T.Iae,I609&7K/76)TVMYJbP:Q231
1:b@MY:QYb20O2f.7+8L(Pa5@.+LBNP@SF-JRQL-S-]FRI7_3+SAN8ceLVA=1Xb/
CbZGCLLOT,Db=JHG1(_A(Ke><X,;XORY=SfT^L>Ae.-.@b2eBXJO;F<0\e_[PF1f
<5TJY7>aBP9;gXa&7b/@Q-Aa0Pg<Y\eH0X8\^RceL&[)#XL7DHg^^X+eJ@@Q;UM:
H1-F^S]?K#W.K\;dGa)0gPa[Q^&<O&=RD;-F8MK.5CY+QW9?(^\0Q/c\ZNe(W8.7
H+F9c.CAKV&?,VY@J2W9>5C\K^Rd<95?gXJ3d0O(,]<+X^CTXPC(L&)&ICF8A=Va
KY0)EY<a9;7;K<XSKfFb2e;3RBH0[+9[BA6[b1gL.9=FVQb0&^6CI9^bb?d]<5B2
&PMe(MG2.E#TLLQIW7H]]Y?A4<J/ObQGdE22=UD[:2XKdE?F:c;B]9SS4??V0R++
GP0IL)JbL&NG)F.OJT,X3X44a]0[1[^Z7GQY)TV:AVB9+Q]E>0=O7cH3;B\],=B<
U#g);YS=P[I5e8KX71g5)\FAO41FMf(\MHL0BQ5O5AB/&b]6TA;9M:.1HE+V[//[
G/L\G,#N]DDAH)dW:8QX?GN?:=a8KF,R5_1AW.+:0Y<JD;@U:N2S]V3=f[@76T/.
3YdR&I=N7VCg^57&cAFf[BN]f=-/aM>L_#?#[W+RTN>;#dg0(]bE]S<DDAD_L.VL
]>XAe^;?+b9_(d2Kd^3&N,A4Y9I_]cMX&13Wf0)9F[=KI[0X4Y_&,^,OUV-SXIJU
ID.:WQb8K7f>4g(7^]2Z(,:c>/I.J,2@?45e?X:EQ8@/-#;D.QY841E7BMLF5@S^
.E-4f2P,8EP)\Y]C<^BP1eXaR/;OY14.6;JKb1B04#M2(>^F#(->9E&?==bdHT@<
NQ_G:84)A0_UXgXMTYL)+AJfZ#U@?JU>Pd(,)C)UK9P,+WVGAM]1OL[V5@c^Ub0R
WH<HKN^J=9;MGE)[N>3@f@S7dGNE3We)NOBZdEZ6BbffH)^AZaVf]]OLHOfRZ+O[
gc<33H(VWfW6+X+dL@^cWf5QNOSaYF#+?T3Q^cR8&S8/(NFGO>:6SX6bA4aMN_f?
FJ(AOV>0UA-(d:#;I.66WRR)B=#36e,Z+1I?3A-&TU3aF:^+K2,LFSc\.-SLPKWb
_eYVN\XO_WU>CHa];W=##VM1X=c@K/dZ7\Q_I_VWH=4+Ma#Q5BeEC7IgD3B,e82S
GOfLJ#8QS>VE1[Zc#U+)7R4]P[B=Y906+6,N0,P6[B1TM\SI[G0Z@(EG6b+K9Y;#
:2L9D_eXLR@.gV-=?_2:G&JDfa(X^X]J_:,BH?>+#6c#,Y5&04ZcTNf4J@+@M,SK
9]4YV:C-&4(P7C);b]<-7-g)+9^d(6ZL)KNSTQ5)RN8HDVKA:P_dUM^L^SEH&\e3
IUDHF#P[,09V4U@BeQZ3cVa1\^9VY_VC^<[gg=4RO(_dR#3.N6Z\0.Ge]bQJNUUJ
[=1f2BZ]9#D\9FH),2J>04WQZdeHZ\L>+#bf>1]R+b0EcRY;<0VLU&(2f:BNW]8I
?=N^Kd82aHGD)C()Qd_LPL3bX(^7e^?NOb39),#-4[A0]cXKfHACNZ&E)NL4e,Kc
._@NQ.>:L>^@(=dPDCPE(=091RfC]+X)e4MO5XD,+O1UXW]:4)Q>D^GXD]CN)cZ@
M,[3&E=.5\-#gW(4&1Xe(gE6DfdBNK)b1FG8d]RIX=S<TRX1#ZC:UP7b52.TI+-N
E6c&5O<?HCI?R48NH_V;.HG/@b@9K4Gc@\?PF43gabK1\>YcM&gOc;X/F-_c-FHa
7=PT^:<K@gB(P[D2dCbT:UW:eK>#bBEGQB>XY5d,&:3AAI2(F248G^&,K)/6J^R#
2@XK1gCN1,^P5USaS5=39.;TT>2AVU<&eJJ:XB-?^OT?Oa0UC9IcQ3a&3+P):WPE
5](=EOb;8/52TQE-2&7cJD<8gW<A5-:.T1Tg.^DF\73YS38:]C[/OT/KI@E<4/<J
g-ZGaCL0a+d\&;C9<JE>GME(G@#9]\(RE25/#<gZ(@g)O[)MEYO8VGA45a7D1&,>
0A\a&+1]1FZ[0Zd5bgPCF-=g+3T:/0W9IP>=d7A]_6a&bQKB/B2JN3e-_a,<\/QY
YIKKCJA:(62I#X[(c>?)<_bIP#T7X7=B?V0gY<b@0#7DcYF<2PFbQa1U_3MbN.L&
U4Cc#,2L^61a559>eL0=W<UCaZ3K]K?Qf1HfWW<\ac161O<DU_I3H/2_@4,;Wb8f
LcIP/)Qa1^13U0SSX1Lf(1T[,=MP.afA\,fQ,7b@dP[42bNP,W1TdOFE]D#25I<e
OSHDRXC2cYOG[3fLKCH10CM[R-,H@KHaN/UCF:UY(Re=G]1Ld?d(gY[(V/#]HCFJ
#ZP5YNA=?eMeDP)NFeLHDFFS.fOdI5P/N24G2_@f/]EJLE\ZJc0LP;<fL1#bPS_3
3;^KgAW@2N2^;6Y^/6<[8g[C&6?KD+\@:VI?^.9dDV01E5Eg<XO/\cNEfIgeBZ?M
I,V=CeVa7FbR,K>CY6GW]X0A3d/T&S:WMG,^YZcS7#=F\@JA1KT;:4KKIc^C+=^(
<7O2#eBC[eB)CGR8AI/+9e<]AAKg7XWde^e&I[e3a0cE=O=eT=>IMNF6O+6)2g(e
FL7EP5+CBcY#,\:D#P4g.eVUA]=C)aW8[YR556JQ1^cF#ae](L5a-;Y1EUQ^fFJg
9cFaF5d#:Cg;SO4,f(3ZY>ID2Y=>.:5@e]PZPX0>@V19IZX_;)K#Fd^[G33^]G.I
__RJ50dGL+Wb82,a(@(M_UeBPBUeIG(:VM9=4EP#F0K)C#^+O/SLPL[YgUB5@I:X
Of@S<K?2TNFW0IVB\aAB>:KfA^^Jde<H)f.X>+F]4-@MB^\X(:T_2/7GdV^[[B);
EbJH5TZFg>4OM:b;dV5YV[<LEYGAT._+&1b]<,P1B8+QDbYXC>28_J5ZJ,NI?Y@,
9U>C:e=H086Y)3TP.cHg/)[PJ(IM36:dTJSHE9U]QMW@ebbO<2=/NK](:Ne:8Y^>
7e&5HJM#cRTPO14Q#XDY;\?AgYPJ:?F@#d5J0-/JaF04b^>&6.g?44OO>6gd??fJ
(c0,TS4Vb1cE/.NP)-,8G,Db6[Y-bb.GLe2\#Y08f_@8^C[RJdRU,fZJ3d&C&V\e
/GIL(d3f[3XG<6;1aF18AZ?e46N.K:ML?^55MH-UZ05P^/ePf0XdGURLQ_GBJFWd
EBGGFYIXbQ[DU1dI6&fJM4?7SD7]9b17](=K^\=WXZ6++1@./U5T[?b>/EH)g.ge
9&J+)/]bfgP[ODY>Ze6c7)gf@g:#CVfZL-aADEY\e+>T5LdJB&]]4N(eZgD_A<[A
:.Bf];)AYLD@]?ZW4[/9^P)eVWeOFA5=8-Y9_<H&CcPS0:cACSY;UB:65VH;g]aE
58+Q78UWABF[V^7T:G<C(_\\\3b[X>6KbD83JR&(3I3a&Ag^0e;-/(^LI^WefNRW
cN/;.F)V9#39U;/8O+-=)<D:E[ML&+K+\c5[_KC+DPT#,NdLX(0KD31]-@N;fUfc
J_]]eL?I&0Q^e8P;;89T8M31O5A&:P<Rd8G&JN6bYZKIWPZL5Ab0K8QR44N&Ce>)
BWB:dBYKLGI:IPH+/LNH7J2T(IH?R/LU7+]47@]6\V,>J#_NJ7)#,?3VSTQGc8K;
WJdKIGVcQ9HB=KOKGMaL#6;J;#,+:O7KKE.UJ=I)McEXX>K]Zb.,NXDSZT3?F>RF
Uf-[aec3LM85MagY3g\Q3:Z#[L].^.JOLE_:_LP]E&BZZ8VAA,H\BQ-P^K:T4c9N
IA/]BKS,&W+12:7e#2cKW<7B8,I_JMVbNW?TA28T5c?7HOZ7SAI31A^fdVF4EGEg
:NJaBdF9912Q14Z(N68P8UP.FFQ&]1Jf6NdfDUb14)F@MGJAJDNa@BdC2XaSceVY
HZgNR4-B^^+V8Db]JEF1Pa3NCV]EAY:-@Y-PC0T3?0)71V+WIPMVF.EXS->=MA7;
Z>JLE.bdB#7):)=.04FdeQ97e3T(e7,IJJ\2\H:8aFegcYQ2K\KcT2fXY/dd_:#/
7KJ-N1JCG7P#L.FISL^V0&DU[T3N>/&;F/d9aI><ZW3XF[=6CYa/C-BM[7Ba#/UQ
#B3#=R;A)@<CCQQ_)<7/^]/Ee(#?0;/GYKR;YM=H:@PE.b;]g)2@<;H1^Gca)W0U
J_L?(f-WF3<,(+.O-g2.H#,83MV6+,N;f(R\(@QC]gZV(&+6.1f,I<D7P6^aDI.I
N3+@+D^[[2WYVY,>(6ROf;=H6&>N4;gP(>/B_=HC]V/MK#WJHQ17MSY+80g4O;1I
;4DQU@982Z\ABDKF0_,I-GW]Xf<FWBCgLK82QZA6U?Db@2I@]FF//Q>RX/^L@,8b
N<S1(4[Z))CdL_;g,6Z<?^PEO8YN1<)B\A3]@6BOJJ5acW<[-cCg>_.WbD_b(&<P
E:J<EZc.?E(&0QHe1)A7S6KWQ)&_dFcUVbe8G+e@QcYZ.E<=P08JP:D<@N\IJ^Y.
MX8eT0;4.6J,(VgT(:US?AfM#)P>e[Xc:U[MaJ5M-DL0CYW)cUO8W,AF<VKJUO]1
U6DgJ03e?6Z7XKP.;e4ae.X2+0O^5U(F@gGQWJERG+&ZS_0LU:R3UJ<<K=-a@4(Q
MLPI)2(2E,H&DZX(VU\CHMA@TG8>Kc?_;3C1KS:(7BAMb[CYCS,gFH7;P[8C)/EF
gC4@H40HZ^P5>JW[@&,7[cH>.8<ZBEdNcDS&PI+@C/[gT.EYH5B-=eU\F#BM_+M7
8H?V4g0Q#ee-T@E67>8;=A9139=82,&:Da995Z.A[-]OXU6KSRc2#.,/LRe9L7-K
c,VdLHBT(H_UZY0[VXC/+.O3]NA#\-cOQM5ANK,+S,-a2:N3::IdVFfWegg<12E;
_J,M2^PR90X8XX[^ZJ3RP6G(RYA,34g,[T@dJ4(/?/]gQL2N(^,?f_&VIXB7U:fW
.bV\]QEP.]B4OX-.T(2/@73,4YV5d8Y@gVW_=W;9?>349@X.:fga8T)gACJ8O)S6
T+8BdcQR:C^;X-8UK;a:P1CX8(9B6(=b>G/J\c-I<(W=G8=g)D-7:.aC+7b8)DXC
)#M2&X826T.Td6:)dZ[VT#^U[DB7(4;-b^c?/EfF21BVPEPLTYJI>7U,V<O&R(D=
BB+4P>9BcAO+2S\[D1f]BJd+K[0N^5a/PSb<:&S55,Zb45L]IQ_HVcOV)>K5]3:5
<;8DR+3>)^13<7.a(E70f/_&VP,4VNB2;^.\T0EE8_3g3R3]J1Ma)SD.&ZL-.cR;
Z^:8&Q0&8:+L:bg.c4>f_=9c(1OI(?a[?R#=b/Keee[HQg,faF7+dT0bJG&]>&a)
GK..gSLXYBN_CD-T\&>C[_EG_W>\Ta]Q<GV(4CB_#59(<[V>7BR@OCc2.[H>BMVY
R-feQ@cL.,UgaD0GLI&Z,X]S:K]/QbJO(_VAQ54#(>AGR^cg@5_N_IOcZJS:8KYH
W3f8<RT[LF4E6&F+_LF[M<=P5&DFZE0S+YY,RJAfCE-_c4\P2c7TSAb@f:I66/5(
P,]dLb)U_OXQR;P[2+<Da3?MR??]N-Gd/KJc;SaMBZX2LR??UP0QaM<_1><b7^V_
]9LNRP)_-/;J-4ZNXg&DW^?/T4RPTLP=Ze<Jf7T[]6,@ZAXW@V[\?4Lb,RCU),@5
9eUBIV<XBI\V95O.If^1MU-gC4^d\e5P]gM3N6bN,Yg>7W3HUOLFSaY6bCC)dIHK
MRQg7&@fTQ/8Ug29V:&\4T>ZB=RWXHL^#:SU3I?&T1#aE.M/X+@@A(HT4Z>HJB7W
E0LG\JdUR>DKW1afF]R[fe.EaR]9.)^T2.e=ZR@PQ?DN5?(O,U+B[e[#&Pf0]L:I
Y8GBZQAJY&6T<BN3#?T^QFa<YHX=Y4BIf]8;DdUNX,=VRe32[6A0V__4M^[2S-UE
PRZ&A@<RZC_;>B(P.Z;&I4?/,.(bJ6K#9HNF_][PMV4_L-E:WV85=RR&5A9e#OO]
c,e:/Z696N\2__,1@X]@+D0Qd\VDCG(Ke-;Pcd[gcS8_^d&KY(5:&^6:+QX,/Xa5
QSS&^3f=cQ:aI2\=9?J(AGeDJaFD:,@BH\8L?A,Ge6@Z@RS<(OI.@H7K5/H5G=4[
?g8YD_eI13dfTCW;OC(+F?Eg@D)[0H1D[GQ0YfDgKdL9?@VE0g6O1K^RUDef7Lb2
(VeV)6)6HQ8WIE[,dZGQ.5=)aH\79DYY9?eP?R:L+54<IGg)ReTF^3.0QbOAQ8b\
V-ZN9-DG:V]8c)(-1LMUDZJX8Q+aRbR);?@U8)DQR)Y8-bbcKLcO8,PgQ1)V(4;Y
L\V[[gQ7Z;#K23-4T.(\2a4f@QVK<.Fe7,U/7RbR5^HSLKJfI?D##),HP6<\>_^4
V<_O<(c_6E4F]D+(6[ZcP8BOI>X1LL_].M1aH4YZ_#N+0>;S3PC=)6XLHIRPX;1?
H-Z1-?R?ba:OFY?eMM54VG)&?^9/2XOcA6D6cVgY]<R)M&R_A[:5KUbAK)NLgc=>
9?O2-QQ(N(9<>U&[LF[LZ>2QY3JNOQI+I;Q5@T&IV2#/=eJ3A=K1I@/[CM.CCPC6
,X2-e1fR,9&H#Oe7D#]&<D?@R0JGI-)2?B4LGH]D?YA-7D:,QBRZ63^b=@RMf-=Q
13?^^/B\8g,MAO\O48T^6<#M0?SdH\(@YgP)>Se3[),E&3]:;BIcO9=&T-^FDZc/
CJ;cYKg65#2A8Af[=Q=M.SRVZ1X,J>L0,[DGOKD/:#[S0PVU#>+/dcM^>\gPQ<5[
EZIVW9DbgIF_06<S^AQIEQ7Gd9C.N&;b8O<.1XXK,:/4KS,#MY.Y_)97a\d&K,e_
F/ALgZZG9F40^_#Y3_.)EC?\Fe?eW)K2TA=\cY=3\\,1g.98UZD)W0@-EW=EM&\Y
c09)fEC-AfGAC,6(A@N<#QT7]&TQO?gH]Qg#DgcJK0PZG_#2;M;ae[c(WP9bJ>D-
PNg:V>]#C_C&gc-V+KOb7=98?3^JN8aS74JdV]5XRa7TNJ+9_bf8@9d\G/SAO(?F
4)L4HDcUS>HUcILJ[QYXRLW,UO@HN,(^-#QV,F3S\QFdPO<A1B\UIf.V1M1=IC#&
<\#bXce.(&[_TD/EM+MPZ)@-J-,QLb5aY0H,2VG5I]4R9<?W.8\A>fEgc:.=I<Z.
)WNPeD9Yd--Z[L_D&EJ;IQ2AfYLXP>]7WeVP[073/gP?0&4+YXZ,eLQX>X1[9d+I
De4-A<U2LY=#F^:DTQ#CDTedNXMLKZ<>J;1(d8(RP=<4Q52FL<XA=dTIO\4EI@=9
bde>,;Bf9X:Q5N(GN)3^eIPO;5XEU,+cO>Q;GB5O2\e3dGKV?&N3aHR8,#A_WAg=
TI?c;)2((Cd6\7UN8^ZUgf,KREe;)R-##,/MM8W3>4I+7<\)5L5\E4W.K330&1EQ
;D=NY+SGdedf/6HI3EFc3N5]^2F75@^U:-D<-&JWNB[S.Z:O,4)N46c8_U5XIISM
=PAe.:b+MO.@<@8UTW-N/M]7+D5C=@62IPZc-J.(7OGP9M,F6D]c,V)@fc22&0/K
bY7A7g?SOg&J@CJSDEYPOP:MD#6#e(P/WaNeVeBf\P\^>d0W_/\Yeb>^Oe3bbgCU
WVcEV89#E>L,6fT8VVXUd2Y8QNG+,XSEBfa4RKg/AKe>b,-67QBe:(#4P^C\[2@#
ZL0c/,Cd.8S8_5@>8+NVZ3ID-NT_M6GJZe/WLYIO?+Ug6+V@583c#6+R(-XIY@JF
Z[8NgZCE2U=P4CPH1B\c9@BWI(\+44:X(E>9=>aQc)1Z0B@IIXJLT\]CAL;<1b]#
WDZX^A/UIU4gC<#a6C<efY1U59T9f++;_P#A&+M0W@MQNR)cV0V>N9f9:/6_AYb5
M-R1d9#DYG88&;CL_]KKL)PE/a<JS4@8D]=6eI8#CS0eX80KYMA\f/I\8SKFa616
IHY9I0=^(RdNNN;d0QHc55Y?JaLb9f00Q0^cXaPTeO-B=C#G4;\NfUVZOUTM:Y8R
Xgbfd-&Sg?,PK;X&\/4A^Rc09NP5@Rc-eT?6^42=aB+R&Z[,LNB>CY:5M/Za^eKW
#cE-Ve21WIW<aS(J3?9/UZFfa?.&=/g+DU&U)CM@+XfW]NV0.HUCfLVbGK;+D:DZ
]\##Rf1g4<Y1VgHdJJ63W^F(\A9IESCYQMUd_@K/,B<M#=YJ9#-&aZ2XZKCfU[L7
W;(fS?R8LdR4HgeI>=?Y;K1.UfeLaYYY)-^<f/3gfeW<<17eDEc45P+7_];a(2YR
Y6;c7gLDVWT.cfVX^)Z&:?d1]8_aG-<J7.#+fV(2N@XXBWGHCNXSAMd45gg\#X40
N94DQ/&..<#89e=#S]7]T[K\8bd>V;S.G8@3)E8=/ba3EX<GbA\T8?T]fJW:4,2V
c?@N5_2BWP.5)bZ9^E6A>9I(T6EMbHZ9TK)09JR,M8IX5^QgJ1:(-#6J1O]QY3c8
/+SJEf1I/Q@7f60>=W.c;/&McMVMB<JQ?\,TXBCQLe8T?-(e:Hef=75Vc4?Y#X6?
2C5>24HF4LZ2MAO(7\U>F,O,Fe<?&&E&Q28-7C3RE?5GUgV+[W9C\ZPTPO>a8>9-
0HDHXd#.a.:9:g9\JgGU;,E@U5X7?/^.Q)M]HM=)+DQXJaA1RKL-=HCb-aW5=O>&
9)26Pbd?.@@\[UFK9a6XZB6_:#X,)YB4X4-.gg]>3S@AEc6\32NW.5HEJQ@FV@VC
)00KcX[S)a]M/C&7MW=OY9CM-;]0N1NSB./J>KPGG:2);IU&Xe/ed5LXZG@c^\F?
#TePF;))MA^(WXK^7X(a]/MO^G-+Ag/XX[3F7e]?UG_,5G73L/BM#A>+Fc(R3A-P
,N)B])/D>eI2&OUd^-GK9@AY>_3[=3A[)[2)@]\#GJ)\DF=>((F:\QK^PKOJ+_&9
NY-3S[d7/5EJ<CK8BVJHgOB7F5IbU]@F4A5deKF=L\UX_=9M_I61QYM?M9A[NI3/
NR?R1gAgY-1g[aTT&^N;(4O#ZMO?87VU/b^aH2F^Y0fB@g4fVYRFUZLSP)K1M5X(
VcFF&eG::I^I3O1GM2YG[F;A#[VKg,[dIe9IdWdN^K>RY<^/-WS]M?aPR#?A>KOD
NU).6P1E_5bOM7/X#EK+KfR.bN,ZR+(KQQcXE(D++LW;2f@dV2fM.EK1Ye9+/(G[
)Cb&2eZ=6/28W9]B(d[60g1U/RU=;6aYe0J[+#4fYBaRbPKQ5ZZ)C=FHPbK/X#1-
\:=[3g]7.ITdHK5B(C(bI6(bQaBdMF_g@>?cQfM<+IfeeDIAEg6(=(?:@1Q#gBXF
8H537K?1NJR]F7H5)IJM\NIYR71O5FLB/gG--70##;^H(7;fMaSE2&?>N5,eYP;@
egId.3RGIb;PLN(S#\bZ,GT9X8cXeFK3Kb78Jb4\9A?bd/J1J+1,3)C8?9<SgNP.
&a9S6HLY/b-AH<=-YBG6(Aa&gO6)DB+&FCeK]Za5JSI[3V.6YH@cf8I\b@WN-<./
IDZM@ZV3Z(U44NVaELF.AdU,J=A;&./R1O/DS=Vb[CT4b)IW8fFS=ZN4gGH[(SJR
@^d<bd=B?)38d+?eL<a[1&Hfe^0=[XLR=Ja0c5SB1B(XLK47&c@M+&GMBC:2@B_Z
0Y[@Y,-1/A]8)=MEfRgeX&LaU36/U2/A],+T7LE.N-gEUS>b4L&B?#A6HM)Qg^\a
D4G[;>@QT9PU:G1J=Kb=RWHXePY./26#H9<H-Q_QaS8-@DJY=4GFGG7f&0-<8VCE
W3.0=IG-AgHdQ(@J#5++ecQNB:_RO.JV/Q7;=J]D]30#^7^I[IEXcaRFa4QY(\4f
U@35LWS/N5(=T3Y78E;^_6)K7#&0V7TG4Z:X]RA.>?8<CgO3@b\fLcbG>E&ZOa[J
6Ob1@IYVd,UOH6B-^[4B^U+M#ddT4SZa[Y\-VdEUfbRTS\S:6[/LIWF<GSbOSGZb
=(a-SM2T&@XK5(XS:>)+OFdUNFBF_=UN+U^O/?EOd3b9AR?##g\^:De1^XOFg3]<
^\@3/8:SC>M=@3Z&MBFecN:8c?5(DMO<G2dH,6N5?,-11==8<HK7T06&I5PPVNAS
5M2#J4R/K+3agPg\&AI@11E?+L9^++LF+>(f,>NEYCHg2NKF7c<]T=];XJRaA0KU
3Y^]aCJe?I/5GfgM0PN#)4@a_PN4\5K@:UC^Z>QR)Q:,0BQR,LdNG]K0,_eRWCHP
ccg?<U,JO@eVD8<^R+eR(ZY2#YS(>>)KcC(T5HXFcdHKG5==EaJReZ7aUFe?@2PX
\0\7UKP5CPB?-3D9<CF3:6U6S6B:Q<=R/U?OI<_F^@+.GRfV>bLGWYKc5P2R/PD6
A8(c)DEQC@&JXP=^S)<_T(3Z&\2AU8KZ2.MM^e2>_?S27@UQKLg:U]D/e/76]\03
/NZ6E@f_bJW4\@T0OdT6?X74)IFb/V/.(Zf?AJDS^P9f7e6AS6C4=Q=@^,,3T6IR
M]&T9G&&^-N^OW,c+abX:V0/EX]Y,8/1Y.9a.Vg8)dM/-3_7J)>N885^0,::MU3T
b^+6,(UZA,0\IW6M2eH:Q,;:_R-]b9<g3ZL40AaWa(>X4JN^54)1CXQVZ+3GE=4(
:WJaM)F9Zf57MZ-M7#=b6?QVSL<QS5C@]#FBM+ND&7N/0ca)Y]@B0I//=:@4KG_@
C\LFd9La@#Ve(EPc9S\]3:JUQPNYc&5D5UV#E-V)5DPK>>V,GP:]YD8QTNS2M=Qb
c7AIG0@^,g,,-c_:dg_SgJ_S0XHNE?f?[]89aWF^\Xc2/^)L.NQ/f:^FWPc8YQ;0
E1)-_]F\&>^5QC-_[BEa>].IKG<-^B53=V)VV.TT<B?dS=K7IKf;&;2/YYTN1dYP
=4A5ZB.P2/(C<A.;ce:]YFU9NS1?7_EZb/]7BX,<AX1[PDMePcE6;EKZ28NI?NKD
9#cB5d>2__RY>CfUF//HEXS&G/A8A^R(WgCEYXLCT<7);DKH(5>T8)U4\;W7)XbN
2QP;A[0XE5WZOQe<83._XfgLZ,]QeB;@7BVIW5a2<Vc[/8.L^)6W_>PG9cCg(_?E
F;f5J<YM::UM&8<+K+K/aAH,PE2((6S?WZ3;.:b\WB,21PZ0c,C#JaAg,:,+ga<)
BVHG=M0K+@-Oa@]#E1_>W\@TdR0&2S[,@.LF?\eE-a=]2F4P.>g4<<e@5^eNg+/I
G>f=U:?7..ZGQ>=gB(CI??ZUIG,fRg;8QAFNe+@X,b..]c]\AYUfF-F85,7JabG4
(B1O=KU,ba-/N(C46HM6E^BJQYTD(PN[)TfTMQG=6>CEcWK]]LI-30\AF98b2/\F
U1Sa]^T^HTSg,U=SBXU?&eV:8G_/EI=H_bQRa-d11GE;BKAPCgJ&5JC49Z4S^B6P
f.fb>7KA_^,UXc<#aT_B8V:O[MU(BJLZLeHS;-@6Y5cT\_ZYfJb>S4WQ&TgH&DF/
WbeeP8+8MYeWR\X^:@<75+E-C&1=L<MNW;8c6/fIP^/5]YX@cZ91;0MQB6>6<+;=
W59)S+_bLGK_].#R2WQ\HY,Ig:Q35)RP>;DU?(BF<5)&ROeH86cd9XP_^P\(C,^L
V33/S4ILg?Z6b,/W-BV/,)>d5@TV#<_/=9#^^?dX6?/NLOIH?+eSe1T]d^W(cDHB
AMRde@7>^SFQ1Y<dWU(S57D2I2N]:ZX=936YU7cF;R;L5?GRc0(W.[&?4:8^\G+?
4Z@0C[YAT:6aFS#I<<@BTHOcBfUI2XBR[R]0MW7-[47B#QIeCP2CB(F>T:?4?C9F
&DMZZ2]Xf[R;=BLQ0Le)+gfK]eGOgc0T>G,XdW_d.G/YWP2XVHc]&BR@SI7gFS2\
@#/#7Z3,g\WB73N?M1Q6ZQE8#V^&E4UJE5;<;ac)f9cV8#B?+<A&bJ;U(;0+NI&@
cYVUe,0B2&<MeG.(2HZA+2EKPW8+bW)SD9GM;L.M>&>Q][HUUdg:OFUZ]Af)FI,\
N:U9MaK)V9U^RFEVL)bgc>2=5/78ZR;<C@YA0NgBI]L[K4Q2^0SHU9N>&DH7OLg)
fG:CN]gYJ)EPF>aS,^9Y]H>O;Kb)#@]4U1P-3./.d;A;2^A\O3#eEa&V<Af:\K8Q
_-:Ie<H7^(U#F<T2W.[]\>KXRdT_E_AA[SR-Ef1Y:=V@(RIfQ+#dZJY=?-;288\M
I_JGRdR//\&+#&XdKXWO0b@K^AYN@-3YIY?Vf,?T^^W5.]CVFg_Je1La@b#YBaUB
W/-E>S:FXVYG=M@g(U1?PX7gT69C(+XLN:&3YH<AFG-J.H:FPK;fcV_#<^5b5K;<
TY9)V0&d8ZeVM:]WI\80_NSAQ3Y5-0Ecf@ER::d5JE(Rf1<BSKNPbV.,/B6;?_LL
#N_X^X5<#S&WaUQ>J8D1OUO09@3)]]?04/1M=Q=H81,;Ed(?&/YAI,I(FTG_#/O<
OMQRSf#9>CJ2aJB-5_5^HH.#,(&J4E&?S[<,,09F>#TWY>?>V?RNQE9^YbG,2OCc
<a9&@R&:\??I9A9,a[W\W;6dN[>\0dP<=aLDJUg@O\U;&G0J]_EB83LPKX^bb6&d
U\+O1NBZ\=K0\1eASbP-&OJCO0Z(b^d@.c-7X<[>.E-.(=VWZLNW9ZU^2R@AOHZa
NN@TNR3<1aQOUc4,\c)Y1,F[O?fUf#X@e9^D=5K2)>0=Qa1?H-0C.W0(YN_b2B#+
/\AbKFZFA)5HF)fb>)a^Q/&D-Z2N025ZAIN&1/CacV(>(.Td)]-(PVOM/T-Ie/SH
]/ZFK.@N2L\C-/QE(>V9&e#MgcW=.SKQ>E=&V&F8W&,;1)CfHegT3&e6)0-[/IXG
K-NBAe7O[Q[2BHOOY+&4LP#;N+L81619&KUd=.GVK#D)WLHH_eOG\_S&1Q0CV-Gg
68J:GOS@YUA/JCN=AJ[Z(NYL#[DEV+21]FKObU86c8-GW4dPaA8g)GaTf(H(2++=
Gd:3ZZd6d&UW:SR5CTgT?TVUT<@&:Ob8^+?e0d+;<EH\T:?+b9EG68D70NY>/8gb
P3;L-U+CWbGQf#B:e8YYL>HVUQYX_--M]T25_,(Ye5fPB9J1H.eJ_QdX>,(,V&db
/-(c=5XOPJ3a(CgbK)/f2U]bC;#_>O/bJ.(>\(QA&f8N+07(1U;RebMO\YKNT<g(
aS?3ZUQ)a,H7)]LS]U6@AVP,D=7>AO\GU>PWL(HSO8?)Nd&Id_KC\?]ZQeL]VSSY
BW&UbEWeEYG3/MX;_EPYceJe\48\Pf_,)IMN_ZI:,L^S<;UG?^\-PO^_\35-]W56
e(Z&e[1I^LSW_/DU&D.ASV.1-#7)V^f._]d/gI)ge[=O2K)g62)C?C)^&fcb;YY.
J#e[@_bN\GZ>QP8F=>;.G;6F>U?@bVU@Ld#?[83+@,CR9Z>?]8JC0cOCfPD:X-g[
V^b1=.,\BOGUY0dF6DIE48+Oc(FA]TRJDb6TVHP<JD/g_T>c^@cNc]KO1V>@BZWK
5<N(EOW[)0ZXS]>,:0<_PX_#=_C_HRfSL[-;CSL7.))H+WFOg6EV.d2gSN(Q6AaS
fg7LU.b?Q:Ba7d(>5^A8aSb:#dV&O#TFQ_Z<8_f20e(GB6[cYDbg]F_QLL-W7+(R
f6g.H0L__LCO<IKH=Ng=J<GbPa;a=F[K2:],8D+a0_)d[NG3B.L4?)P,Zf)=8/IO
\d^D-@S&A16?/1/d4G6QWC6[PK]+O]T_7f3])_Fa\CC_X3N.?G/]NQAR7\EcK8+=
(IJ3(8PYcG4.gX8-aRf\1X0FaPI1>)+#XXP:?X.=:^9#W,+(d,=YNWf(KP)Y^ZOT
RfWM19ga,OQ)H^SdO4Cd1Ha=CWN]0HUGIgZYPHOH)2[S]e:+3@QXR[(2T]c^F)AD
Z4^K12eQ,3bT,8VceR?R,4c27FSN:3D5V;RXCC\;()+ABU\.a75FQ3+1E?Q2Q;+>
,K;b^]5=fg;LG-J24O_Qaf;@DP@Mc?c=S=Y=C4B2ZL5-7+e__;[_d/WHcCGeAS:/
DDJ?ZR=/PEGE73JHUEZcX<OaC82VQY#4\@KQ.7\67GEOS,P()75+1Ye;PEHX\[e@
CVX\:[HV4[bL^Q;?53F#4+5RFB))Je+b#KXDUBBW<5RdB5&#^H7b6IC6@(agFV2c
ARP;@F=b^^B3e5d.^&/Jc^0Q4DM,0H)04\SQ[K)b.HW,&]3WJQK_1^3VFMWTbM7A
SB?;AD#:56U[da1[+?/fc,KdcE5QQ1W(fSUX(IM:EbH;Qc@fI,8T>;/R;,;AT1cS
:IRW=;I<[g)?#-FVP=Z^CfBOCE7LWWd>VceXLZ7])?(bW(1f,ITHFQ_,=B2U8M7Z
:TGHL:W[3#?&5OT#WUUbCe];)5aQLJCW[OJgX==</AW=?W#g[S@IKE;Z&eUZH6eE
UGHORb)bJeYOAf6RD.KU8P:Wa<S04?FD^O5)DUQ8HF[L[eX0#<8gf,351JOG9O9K
-fZ=6UAX;06:N@DXH@Ya48SIg5<-MCD&ce1:PGSeXFed2)SA.)K=>O]8WU9#?I^V
PXe]4.C4,-7^:#@0cEba]+:&JZ?_\^PG@Hce<:e,UF-FU<fI3AWE)1[;2XY08aSe
+ESH:#BKNBA-P3AF[AM80)MBfX)F@4bVIP^T-BZCb),bE3&^2[VSGb3N[2gI4S.T
9N,c>@-c8IRIKH^X52DX<CVbH7WURL7@PM/,ZeZWBAET,.18,+E5Z.K,#/&ddZ&P
OJ,1X18<Eb18f&(6XF0)43@=b(6+XU:JVCKH7dSc()#>aeJa>+LMDH:^\[KQLR+Z
SL=I66V(R\f4IU)20@.QdD1fH\>>ML\LL2bDLb6-UV[GUY950bcV/4ZL&X/F5T#T
(G[VN6I2ZMGGf-Q4S_e0QP._O)BXQ7YF<2YL0<9^KMa3+I17WG.&_-Xg3a=V+((3
cYeJFeFPA@9Mg69A\454G>M8(;RTS[QP(B@d=>_=1U6aZHUbLR9C,Z>LV\M)E:d^
OHE^RP0M<4TB8PI.-I^+E2b20>X2A.6JDK_>g19G.5AUA\P)VYTRbPYEY^D;>3.[
(4PT+FA5eKPggU+7FQ=Y)bSdg_CTZFMY,XK8fLb98/?;ee],D,0V58(X^E1I&2JC
,Lc\>fVb3U>2^D?ZO_Y_GZH.PFJcZX+[8ZLY@OI3OcS)[P4[MY&Q[P:0TEA@LGOL
2.^cTa@Y1c[L)EV=Q9+&A5Q)H.W\<3e58C5b8OT2a&AZfbD_ENK=N],\Ag68U?Cd
W275_SP<[1Y@)dU600^=SG(=a2LY(deX5aTB/:KFWfKY.A2;Y]VcMSA^YTZ>EENC
FO2T6>D[ccXPY4ZCOV1-Q#\3E,5BeO)[=#UU>YW#ddc7,?X;K1Sb^E/^IH[OUQVM
c4#C^+]0-MWUb\a56[8,Ld:/K;P#O):O=U,I#+GC-V.8R+a,<1=g?cA(0S0#X@Hb
J^9>3O;H#SLFLdXC8BaD0\W@F6?\_3YUW0@cc),f>+L#e@557EILO,3SE><)6[6,
a4[71KK-.gN[2gSRc+?dPUMMe+NFZ6JQ^-D,00_CC[N.cY4d^&6Af1?M8RV+g?3Y
7HK;>e2H]]1OADG]de-#cFc3Y0>CR[&3Z+5914Q&?;b8YOK_#PTS9GR?DNNB>7S6
V5C8D5?0#_Jeg(8=CfR18#[@MLS&Re-0IVAZeW>XbNPEd,P5N0TM)#Z>Y/a-^9_e
e5L:adaR])E9eESC[Q@XFBC9;98Wb#XF=Rf:)3#\&KSOHVb(_dZeTTHP21&HgN]\
=e5PLVL9)M]JW-)bM2QQI#M4]4??4b\JW-3N@-(70_4Q2g0^VS3-7(8PcFe5MK3<
VZ95>MEcUg+]D4>8_^fDRE+DAYPBA7T>T^AO@SP/K(gCG]\246F<[B;+JX,EG,F;
=#(\ZUOV[a.7^UEV_EEH1WJI6+ZVF9QI_G0]V+E/FSGPL7be8[BfNbUHL61:X#VK
3,^H<0>?2S^(dN2H27?a_cML-d_-Zc75^2YW+\VdOYTf\Z(P=;0]D@KV@WJbfC33
C9A&.D2b.6FSV@@][;2B.0V=FdOd0f3KJY51#OdLE/PZ6YH:DT3a=G#E]VNW,HDL
5F2CF4NDW@>B:^X?>6ccI_KB0U3SQL-feB-#/dKL:4.5#W]fS(b92AUN8VY/)dMV
4O=XW-P)OU#3&<.d8a?Hcf>NKa;_dH02E/JSNHKRBP]<VW>&_I6#eW]L+B.HfVR,
+8T&>F-dBfN9UH&9=Ga_[F<Eb-a[0)&VJO^N0J0):9fSXS,+PV&;<UaSbH&g0./0
PYV^5G,5a4([,b6B_>DR[G@cZ+A6Y&6>(QPRO2c+)+?-cJc1.e-);25YR2(0VaCg
A#DL\33U;X;XRV1_]OR/.#BXOPZ]Y&B&4BWF,G+2fC4/:e)b+N,7.N<&BdGecZX,
Nc;GW9)I:AIQ9\1@caN9]@\F-82JG;@-N?c0?VA@U3cFK&Sb7A19N.[<6KSFU8:f
)<6XBNDO_J-+-@U2]e^_@Y:f8-Ub18J-aXK,OSd\XN>TaJZ9BOD^8e>dL-]WIT-Y
,_.9c]Y+DWP2677I[fb]-/_+DIgQVM2;V<B9+[=F?dQW0\W>:5R5/:>AFWBW<X[]
1<e-:+/@4(<g9a@Dg^fYGGBQZ_+?X;;F=MI[fWI6>bH-4D0MV_QYJD@OG0\I5LO^
<^K<-3&X-8((#&-)d2,6[:6dF1ZSGdP;R4bd>P8d<;FCM1/+bTX@);AdNHY-;6fA
bCAE<geA2g_RU6b)gTcLa0;fAR0f;dOcAO\\ML)T:Db5(Da31MJaa8=\9a#,0ZfT
<34V56K1+@><:/\ES)bbZLB^VMI?13fbGF--ZfdaGQGd.R3dW4\K=+@3WQ.9Q4RT
UE@FD2_5-VEa?cD08]C^Ec)TAWc)OV_g<2E)#b#FG=[@>RWJHbAKJU]e_c-g)]CH
_Ab.Q/_;^C+8],K2OT)FREK-bdg-Id^5.1NFE3#XWO7@_=CT/aceH29b1R3IZ\R)
6P[SD1Kcb=d=&THHg9#4/A/<eLUTf+NUG#JK#f5:F@+0#J9,6KcQY=]2CMOQ2+(f
OH&dNMCYO+?)KADHXb;g#G:^SSf;+3Lf?)]R14A,QZ0V@978Za7TO&ZAU2^.C=S9
]<6=7Y^<QHdXXV?;RVHB?)FJKb,bQ2TLCfLb:+K+d-+2/:))F]LT49BP(D&PfXfI
@2dLS\Q>RZ+bdV;6T.A:Z-=bY^,fVAB<;-Z)#8Y=3+ZB6gXT@Y)L6T1X=_=aeO=,
g6gHWI>#d4T_H:HPG<Y0eZ(g;M?N/a#]Rd])+^<e35UU&/O+c=&;b21;<9008ed.
#=.NXJ?NIP>3c84,Qd>>8EI)\Rd^UZ^Q_=dWNPfd4,3_BBf2M-2O]]V]b0_1,7^f
c+?7YMA..+F8(gF:@DQ^-@IGgJQ@Wf8UXVS5eId+gWWd@Q]_//;Jbb4)8,NE09[H
JG+V+YM&P.EZY::#&W^T.gR2e/NK;<X+SOM02O:e;;<?FZL8cHZ\R#>ea1H/?,OR
d47WH8-6UXgf)MX\6V0gH/]TF511R-(cD+MQ#T92?GB6G)(8ZM>Y=cN&XA#KVX&Y
X<GAHG/Z_X0eAa^,BC>=TQG_K81P8?@@+<RE2JgcZE58cYe]4d7D8^;4:-dV0V+)
bG)J,AY^TG5TJ3F>O4THYO]LJ;#JATS+/ZUQc:<T5<c5)M=#P#?A7QU5=TTGg)2U
L83JHR?B_B[/V_4f7ES2?XGB7@3?5_DAIf_+cT+T=d\3R/_?3SGD4fKgG045F4;X
fUHUUeHH9]\58O\<F5[CFWN1/S5Y,:Z/F8R)R<:/eG=N4_5LLU-M-.><FCC)D.&N
B&/:/M8)/EeYG,)[F,<@:bN)VN9NdS&70Q6#MbTbPBZ.f<:J7X:b3_f0=X,9d,AD
&&,_+#40XDP0-HV-@(bgXGXSc]<c@7K[=\>:JJ6abX?E2=ZWIB8)S.\(;=C#JT,4
RbgI=\D6IL?SXRI?UWO@W=2Z,J):7_W^ME,IC-BQ1==OJ_fA^0b=C8B<O(D,g=YW
M4ZeBE7^;#]>3:Qe>DU&MUM.WVNDc,Ue@-[/UX]CU(,7/W,g2:6WcZG#LDK?7G5N
<#FYB:=:ag-S5)g0FD>5.;-<LAY02ZS5__J?BJAZc+NfDaJGW6JCQ-/]P@V]=bF6
dL\&3]#U/;TTJM\aLG[4cL^6#?G/-6M[=JK3I9F0Lf_KI0Q2c8R#YL@ZaH/U&)aC
A\@84&U5_d978[M=A\ZbVK3TQdQX;S7T5+?T4a?[/Y9g&1R(GMbB?Se3L6dI3,-_
?-N;)#QWY([[MeQ_76)CdY+QX^VTgbdcc#.:P(eF;T,F02Q()7a+L6BBH>ab&2Z1
&g(b_JTE)^a//d^Y0=X=,SV^HM[(7:K102a3)SU2dcB,a@X#^bLFb?6S]a\;g9R[
^7O8U3:W(4\0AV>&47:OgXf:8?NVc?0g#S1b;<C]?4ScgU>+,?NW,/1AQ#[==PZI
9J./T#?O3K0G4@9@BN;(RTDBKSK\&NP[?9)1(&/_1g-?OPO/SOGU-A^R7=FOC9,6
PD5IOW^EN7I,#>:B&a,)UF;V/T-J1GL/+O)0I0f<e_bG/#P&^.T=aICXc0_aLDRI
5d]K_#:X#GGM00LQb#,V0fc#cDK?UcEe)]J@>0c:L<gXb.3VF60aCH5#;B2NX5/RR$
`endprotected


`endif // GUARD_SVT_AXI_MASTER_AGENT_SV
