
`ifndef GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
`define GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
`ifndef __SVDOC__
typedef class svt_axi_snoop_transaction;
typedef class svt_axi_snoop_transaction_exception;

//----------------------------------------------------------------------------
/** Local constants. */
// ---------------------------------------------------------------------------

`ifndef SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS
/**
 * This value is used by the svt_axi_snoop_transaction_exception_list constructor
 * to define the initial value for svt_exception_list::max_num_exceptions.
 * This field is used by the exception list to define the maximum number of
 * exceptions which can be generated for a single transaction. The user
 * testbench can override this constant value to define a different maximum
 * value for use by all svt_axi_snoop_transaction_exception_list instances or
 * can change the value of the svt_exception_list::max_num_exceptions field
 * directly to define a different maximum value for use by that
 * svt_axi_snoop_transaction_exception_list instance.
 */
`define SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_MAX_NUM_EXCEPTIONS   1
`endif

// =============================================================================
/** @cond PRIVATE */
/**
 * This class represents the exception list for a transaction.
 */
class svt_axi_snoop_transaction_exception_list extends svt_exception_list;

  // ****************************************************************************
  // Local Data
  // ****************************************************************************

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  /**
   * Array of exceptions, setup in pre_randomize to match the base class 'exceptions'.
   *
   * THIS FIELD CANNOT BE TRUSTED OUTSIDE OF RANDOMIZATION
   */
  rand svt_axi_snoop_transaction_exception typed_exceptions[];

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`ifndef SVT_HDL_CONTROL

`ifdef __SVDOC__
`define SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
`endif

`ifdef SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, VMM recommended "test_constraintsX" constraints are not enabled
   * in svt_axi_snoop_transaction_exception_list. A test can enable them by defining the following
   * before this file is compiled at compile time:
   *     SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif
`endif

  // ****************************************************************************
  // Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_snoop_transaction_exception_list_inst", svt_axi_snoop_transaction_exception randomized_exception = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the instance
   */
  extern function new(string name = "svt_axi_snoop_transaction_exception_list_inst", svt_axi_snoop_transaction_exception randomized_exception = null);
`else
`ifndef __SVDOC__
  `svt_vmm_data_new(svt_axi_snoop_transaction_exception_list)
`endif
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new exception list instance, passing the appropriate
   *             argument values to the <b>svt_exception_list</b> parent class.
   *
   * @param log                   Sets the log file that is used for status output.
   *
   * @param randomized_exception  Sets the randomized exception used to generate
   *                              exceptions during randomization.
   */
  extern function new( vmm_log log = null, svt_axi_snoop_transaction_exception randomized_exception = null );
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_snoop_transaction_exception_list)
  `svt_data_member_end(svt_axi_snoop_transaction_exception_list)
`endif

  //----------------------------------------------------------------------------
  /**
   * Populate the exceptions array to allow for the randomization.
   */
  extern function void pre_randomize();

  //----------------------------------------------------------------------------
  /**
   * Cleanup #exceptions by getting rid of no-op exceptions and sizing to match num_exceptions.
   */
  extern function void post_randomize();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to. Differences are placed in diff.  The only
   * supported kind values are -1 and svt_data::COMPLETE.  Both values result
   * in a COMPLETE compare.
   */
  extern virtual function bit do_compare( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * Performs basic validation of the object contents.  The only supported kind 
   * values are -1 and `SVT_DATA_TYPE::COMPLETE.  Both values result in a COMPLETE 
   * compare.
   */
  extern virtual function bit do_is_valid( bit silent = 1, int kind = -1 );

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Returns the size (in bytes) required by the byte_pack operation.  Only
   * supports a COMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned byte_size( int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset.  Only supports
   * aCOMPLETE pack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_pack( ref logic [7:0] bytes[],
                                                     input int unsigned offset = 0,
                                                     input int kind = -1 );

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset.  Only supports
   * a COMPLETE unpack so kind must be svt_data::COMPLETE.
   */
  extern virtual function int unsigned do_byte_unpack( const ref logic [7:0] bytes[],
                                                       input int unsigned offset = 0,
                                                       input int len = -1,
                                                       input int kind = -1 );
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Gets the exception indicated by ix as a strongly typed object.
   */
  extern function svt_axi_snoop_transaction_exception get_exception( int ix );

  //----------------------------------------------------------------------------
  /**
   * Gets the randomized exception as a strongly typed object.
   */
  extern function svt_axi_snoop_transaction_exception get_randomized_exception();

  //----------------------------------------------------------------------------
  /**
   * Pushes the configuration and transaction into the randomized exception object.
   */
  extern virtual function void setup_randomized_exception( svt_axi_port_configuration cfg, svt_axi_snoop_transaction xact );

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_snoop_transaction_exception_list.
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_allocate();
`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: Provides <i>read</i> access to the public data members or other
   *              "derived properties" of this class.
   */
  extern virtual function bit get_prop_val( string prop_name, ref bit [1023:0] prop_val, 
                                            input int array_ix, ref `SVT_DATA_TYPE data_obj );

  // ---------------------------------------------------------------------------
  /**
   * Add a new exception with the specified content to the exception list.
   * 
   * @param xact The svt_axi_snoop_transaction that this exception is associated with.
   * @param found_error_kind This is the detected error_kind of the exception.
   */
  extern virtual function void add_new_exception(
    svt_axi_snoop_transaction xact, svt_axi_snoop_transaction_exception::error_kind_enum found_error_kind
    );

  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and returns
   * a 1 if there are any exceptions of the specified type, or 0, if none were
   * found.
   * 
   * @param error_kind           The kind of exception to look for.
   * 
   * @return                     Returns 1 if the transaction's exception list  
   *                             has at least one exception of the specified type 
   *                             Returns 0 if it  does not, or if the exception list is null.
   */
  extern virtual function bit has_exception( svt_axi_snoop_transaction_exception::error_kind_enum error_kind);

  // ---------------------------------------------------------------------------
  /** 
   * Utility function which generates an string describing the currently applicable exceptions.
   *
   * @return String describing the applicable exceptions.
   */ 
  extern virtual function string get_applied_exception_kinds();

  // ---------------------------------------------------------------------------
  /** 
   * The svt_axi_snoop_transaction_exception class contains a reference, xact, to the transaction the exception
   * is for. The exception_list copy leaves xact pointing to the 'original' transaction, not the copied
   * into transaction.  This function adjusts the xact reference in any transaction exceptions present. 
   *  
   * @param new_inst The svt_axi_snoop_transaction that this exception is associated with.
   */ 
  extern virtual function void adjust_xact_reference(svt_axi_snoop_transaction new_inst);
 
  // ---------------------------------------------------------------------------
  /**
   * Searches the exception list of the transaction (if it has one), and removes
   * any exceptions of the specified type.
   * 
   * @param error_kind      The kind of exception to remove.
   * 
   * @return                Provides a handle to the updated exception list. 
   *                        This will be null if all of the exceptions have been
   *                        removed or if the exception list was null when the
   *                        function was called.
   */
  extern virtual function svt_axi_snoop_transaction_exception_list remove_exceptions(
    svt_axi_snoop_transaction_exception::error_kind_enum error_kind );

  // ---------------------------------------------------------------------------
endclass
/** @endcond */


// =============================================================================


//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5lF2Dw3bPsFItk2i/TprZTPTXPDuDROzhxWWKzXiq3Xl2StUXFnpllaJHC6rWdLO
qeOMjojSttqTGu5DvAY2kiEHNgLTvIgQizPono73rkLKfL/eYtFMDIObJJ4Bj7kB
VxbaxH5khuVcUsNiFGaKFvV8XC+aZcX0CEOdQpeMUvyBVEyFk/XZow==
//pragma protect end_key_block
//pragma protect digest_block
wFrrayxcQ5DZjI4YTROSRLEgkfc=
//pragma protect end_digest_block
//pragma protect data_block
edmR6p/XCBITBvVs5zfaOyae4hJ1vZ70Et8GwG+g88+ty9rcPbWOvMk4EwzF0x2V
iQgGXHfep5CH5B+EiWhHPS4O9OjSqXOkq+9ErSzd6IgHVLic6pR2fes53j2Wc3H3
mvjOKH6UH9sOyRyDuoutMWJTX/hsxvX9KVM6yljgCHJ8HT+wZojR19HmX5YioFhA
epnDq82T7AL67bVzj0FgGIavYV+Q7Jsa4FuwAUN+kgj1ig18PNg6fWfz1UetyrLS
UvEfBBywC/DV3nEx91u+QhhyRXG+ZsTkOb5pWZ6DsKKyX02I9yktqWhCpu2u4v1Z
sfAIC2Vy5dfO7UBveqKZaVgV3adWDXlb/lprxMtV+iFOVr29efY9TUQV1Ir0Mu+7
hi5NllAp8HIizAoBrqXV/9EFyby2H1MKvwksUXrocnxVCzyJrdZWxvhtQvSoTDVY
UXUWU0cQIOUxB71Svlc56C1SL8svLsIFaETXf3UWBQLTPdQSztXtMyPzDDpKGPS3
TWydxLJaqCICM4yFk+oroaPenWLeVtZRIIgg5Pc510gyzhUO0xlxRt5NM/Re8GHF
hRkSovWFdMA7frijx5oFlHmbG05GKNw2h6K4sFuZQ0m4CsahaHKRZ8mbPl3kltmP
ILRF15NoSZr/mJHgKV0Psm2qoIkPqZDS/FKivfPPdrv4avpTt4PVrjdhW3dNvMO0
90jYeThxcMUa3r0rZiDmpLz+wEy1ZR6zhvqbKBmm6vvE3P9f1ZAVAUFW1UAm/MC5
9xTxyC/FEUWZnRQKDqBo6PF+rOlifMHNw+QE096t53DrLSCu7Hh13zkp9FqqJMfn
LNO3/rF9cB1sCo0NylKqOvLGnomOANLzZyUAv2mfoTWjAp5EHRgPSJ7h+0zr+UWb
anrpTHBEOFKduM+y/XgzFgsHAROogKjEvIHMZDemEglkg16OSfvA0ITK50fRbhBH
1BoYVAPCFLdTn2U+kyXNoR2n47wQrBFJ9SlXipaRULo0/0d0TxitOPhplnQH82yj
2Shz9F551kiILjy+j0psF0oC95HbEvpDI3Set15cK+IrmNsYT4YWSys+3Uwwnall
ngunuRqP86nBRf4QCsyrGNpooNGqDVAbtAPlIYHko5M1mxSXfkm6FmH5Um/+0gYw
PNMsxoENyXrEXtXb0nCZCh9JnjGa8rEUu3wGJg0nrXJKaH2LlOsSF5SJFCw0rwtX
iLv21oG0x+JMThIsZ2hbtaB+mvCgLVKqV9Vs2z+oafCO+MtQNpu9KdkSXNu5vLmW
HS0xRwI7GsJInq9san6hGHtfCYA4oOK71XAlcPqgWhf2xOJ4giYQyxxgoEAxGkEN
C7Vx+x9oDjUEApj3LtlvLuON2EJq136qFg4q/9tWp6jJEAj81hVzbXQfJKfCNybV
a11SyzWU5ue/sjITIs83526hfiZ3vEqc0Ms65rLG9jTVXGpXrr+w3upHgT+29Znq
Bfddoc9cu3b+0rfNrjPbTtKhSU/Xt8JeN3GrM+0y+pDBX87b2UdEGjjaAexTFWec
NDrx78eT+ozj1RZTB2oSsw3BiJMCFY/dshi43T6RMKnEE9ZAgLA9+vAtgRMNHYYW
z2Le5rc3YyjEIMkgFfx4YQUD2EwNJlOf7GILLmFm8eyUwxqUUoPAjlYVYsI9XwiA
9MfZoUJEcxJgvCluaMN9BGI5wtra0Pg8Be1eGTA+qlvZRIiPffCJO9HWmgWj7XP9
fLElCKv3rnxSwy1G3TDHz2WPHCxpkU1Hqis3vrMBT8ErmndIuozahSi+X+H3mdix
aZiW4kClX8IW4ZisGCE81MPUpNE59B2wIndlKw2/6jxtiqaTBnoaEWwEnt3bkx5n
9gcDaAgUUjFteWkYUCVI5EhVwXmSW6UD23hIX9qC3b1sXQqHoyNlf7QBgGAPE4Q5
xEs28WskYJpsxZp2kad8n9Hqamwk9B0LqAzBkieK5o/tPaIs+e9Wo9x+nN6Q37nT
g/q1W3qlMe/2aazJ6EkPbmVzD6AgllHMBBLDkV9qOJWHXUlMRRQ4aKOG9PZI/XOr
bY+uc9z1HxAi2eQ+VYFRIYHtWn1XH6+gCVxHTvq3Jdg=
//pragma protect end_data_block
//pragma protect digest_block
YAWzEM7Yi5f+Wzgx1E0qMei/m10=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8mb1anTcKgJOtkYYIIhKN4kDjCaEYH4d0mLxLwWg6afi1Ls3o+if56U3jy/n2MDU
zLaygkZ2fMJe4iFcq+kPRBS3oFdjN052gbJpl3PZkdEBSe5C4uSVPJFBO7PNLKQW
ruY8WcyEvkgJCxyOJG58nmwHAurnKRPrv5/hksmJry48JwJDqoZvyw==
//pragma protect end_key_block
//pragma protect digest_block
3Dg+S+tAmZo0EAhbklrHVckKsUc=
//pragma protect end_digest_block
//pragma protect data_block
ykf/SdsFcaX0VMN5YkjtUoYDDAF74cqAy7xaUbG7At/1buCk2Rq/5l2q2Shav2oj
oiCkBT0iCO5rMjwVdVoZf/xkcYn+KeFj/JiL2JwLN4/96UD7KGDYh7xDJunHmxiy
ketQx4O8UcxyEwgvcQtLrxJAwTnsANMpf18k9SyMWxf0yZEx4e7LrJTX4Gkby4Dc
mUaJJAQqaeAYY4H2NB/N12Ld6zRGAoq2Rdu6zLERAHtAK9G0rXFyE9A8sW4VlnOE
AF7ztJwOlKww4G8oao52zG9Pe/4lGhzi7e3K6JVjUHukdHoWf7TZyhzios9yw+n3
pSs0FUit5/5F0lbZs2FVFqWPmIWKrsXhU2upXhlz01ojgw5kWPpMFEcltbnLctC/
5nLyu4aJAJHPiBmJ8TJAUFLiiJOw4VQZlvsV2A3YUc4xEYriJ4p7kSRP/RIkNp59
BlyDulNnajF0AYGQ0UGU7H2vC1IJ22PylcT/P+fzKvrpvvQ6XeJ+r188qCTqJzoC
1nIiRhj7Dy1snTywB5Y3LH/TiMFLOYBhBd3UBWLvK08+PZ/ZMATCCoQysw07jv8L
nzPs2v1tvJ8SWXI+KBEiuah6HUThC3UWe7fDJjJhUdYkjvTJR6HzECrAXu9fzFDy
HRGzQwan60lSI3RKnzAAfNqKHRov+Uy2DLIoXxaOfmS7PJ3t17gJ/jd4cUa4H6cK
nVFDzZPXShnmvaL6IQRh7YAhL6yvJvMyiHVJffoW3/rY8d2Qxc0OEbUChceRZOix
UHJIsb0FX+qS6Hb2fP6kgNaLZnQKTkc94SgNQjcxtow9L/Tre+N6QugEx+3S1gLj
UmNJjZBPZVyn41amklopTdkLrQl2MIy5TpHMjdR7zsRDarjl4FXB3HN9BTt9PJ6H
jA88GQMB+Talv22kXf23FdmE+0qpRe8j7ILF3I8iHMrAHtyNuNec8gqEv5W8nTRF
+N7sKvd2sZoMHMv4zrvmAvso9puH+lOekRkImj+8tUGQHb4paAC/psUdOQ51Kz3g
g3k3pP6pIN0uSIcmdyMp1czybYGadPiH5Gs8TAboTQOK4hV7VV0k+J0b5IRrY9bO
YyAbo8Io3KMhorcEkmGwnGBEtnCLc2Gtq+G7TvxJBvnfLSlnSSRW0D1dmuDxak7s
9w/73qnp+W3jRmsFmGpPce/lLG+5w2nCW/ukcVS+RO/bp9vmxdkzc9gKRMSioQez
6dgxfgQoCrrK1Mhkc22sUGAldJcdcizIfNcpIf56RYeo3fj9MlRTIpCTYkmJnGx1
mcfNa84ilhZVDAAOrxuqJ68kDLA9uDb0y/rrwzQzL1wRwmCHYZEJxTe/ckNs5jcQ
x5R+zq607SWdYdkUgY9IOBG6xb79kU0DfedGE+uZfBxH+f60uRm95hgLwV3+6OoU
DHdhKHTn+kO3sdEir6SoXqRRzw7mVm9zougQKatAUMdmKHTd0BcyHb17wF2qZzbu
yI51i9ivyY5XuYCbv+856ReNOE1ZGid7mmLSpETsA8jOzMjlO+jcWPM3kMI1nj8L
5EFmMV4c/REpR1TEtzdC2vAdxI9S7+ifZWLeLqrVemI3xiic8gl61l8BHZPNGSV+
aL0WbeyCGau4W/2AXnmJTC9H4BMD8h9LrNFpAc56sN1k1nWINMd5Opm+107oscA3
y6gyfNwnASUECxHZJDVdLKKvS8wGCQiQ8OeLWquz/oxjU73tWwkAJIKMk5HvTP/l
hIU0MNdo5KUFRKuE430CGWES3Ow559jARj6JsMX1+6zcBHmcO1Qj2mWmglRCHRGf
kU77svWubplsPKSPK+audnIBLCJ+ttCjN8clr0mlthcpoowvNJ3vcBMs3ezmojqW
j+lfj4/dZ4vODrTvYPfO7Vdmg/5qP6i9wS07ADe/9wTUmfGC2aMUgQydpbpIOLFm
NhsEGPasc9GA1xgm5u0cehUsoQlwgppkY+NZCZXAXeRuHCf5AB4LGDPPpcVLhJUr
paM8kX+c4fC231WR7adnZezIurgEH9BVIRzIZjMbVOuIwRakDFNb8LOZvwzVhGS6
KI08jxbTZ42CW569Wnhp90GyaBFXYhRIJaEaImKDqYpayPysFOv56X+axHK/RUDH
5SAv2QMxp+iWWP+sQGTvwp/xQnVtK5NIgQ1J/2uovbUfM1tJmJnauqZAucAxDudN
Ai3CcFMxV9NPHpxfNVHau0BWIhwoFcKPJ9mtOQ5di61j11syc0+hGruL4pux29+V
84OnvEYb4EH2cZwsR771+u9f/+GBZtvYjjk+oMQA9q07t2CNRg8HVLz/SAuMHOWk
gl1xJ3WUeHW2JKctjY8pyAERPtAqjITcmxsAqxicT9PtKLqJyPTKRkukXnVQ+ZEc
nf1Hb60awxpgmwhu0qPhShLPcAqyO287SVY4qXSIQUMSkT5364KVEnz40PHeg+W+
nnUS5/t34TOiBeua4uO/GBIOeBAUv665rO1rUt1xI8RUPK3PoT1ck9T2MLnMjv3e
I66AV5wlHoYL6Qdq40az0QooUTAsW9+MAVOEEHCJXlmXVYAq56b6UIp/EjXOPQU0
Y4AI3sMoygNYrD4bY+SNf8PVzPflHvRAYgYKOz/lyv01PMC33TmMD+XYhuVjh5fm
dapLRjBK4MpwzMeRIVIaQ5biPQgY2wwLuakfjT1r/+pIPRqDDf+ZmyqT77yyMTZn
+dA88Y/KVM8U6MLi4r6Mi3sNmMjIDnnXHNskAS6kJZi0vWvwt1IksCFGzpQ6ogJT
84i8XsOxoT/k/Jz0ns9TcmHMDpXL4ftoW+7JUMIhLCKZ5PtLtvZHTvjujulTLacR
vytSm0ZWW+YrF8AhJAq+cuDB+c0YK1ggVSGE6ussIqKFk+K5zocNRtCPvtAJMQLT
NjHmHGr+0SBz7Os5yYf5YJPZBU8XxD8ZzQd6gHpGK3wVv33ywlsA+KY3vNU/74uA
6H3Vc0yz8qnrMV8b1MJwKPlKBZa6zvXarwqWV1sDSfp1O14VIqxb27qrWbNQ5JJZ
JNcg0a1Krp32L0mi7TnclzHJJTu3ncaeDgbSJB08r0/WfmoN/PUK+6qealIx0ROF
tAU3JgChiTNoOPSQGfArG3VpHQLpd90I8BPoF/KDKe6j0vENivVMBklAO+VNdre6
6vQ5lm1OHug0fy/8bKhAJFI96YCYujuAY21P46iFOnYOEoC7rUDzUtMR3i3NANlq
yuTJitqlDqIOYc4sNdj8GlRlHBFsJF9eigVnVToXWVVUdTRl/m7L7NUcCGBXnGiX
6OJIPny+jBqaIzntVS1w/XfxAh0mBMz/nNkAmWmCbTfTMZ6sBhnYpAsyh4Ka9/f3
L8tPOrhhwVTVdYj9yqE0tHVtuNNsRyRFZ2Pp5m66tbGe7OL2dMDHmkyioBr7xeXl
EEd7LNn/jecVlfYca53yFolIl6dDsv3slPtNh9x3WN+sVkYYft1kgIV6c16DD2jJ
dGt+tDS6hanqR6p4g1MTlUBm539T/EeuR/3f6ZA2n+TKcVXsFrEp0qu7wkoMriqx
hANeEBG1ca+46VyYrB+EvVCakfWE9VTnWv1n6s9qQ6smF0iQO+VChAVedae4KaOF
dqt2H6Vptgr7OHqOEmxtLjjoEg8vYjku1/YIAEHuH1sQaiPcfZ4BXs+h44HSDAFZ
oIt4bh1torUNnvdHnYX2sCb763ZyjpP5gqzDJa9S5RFtsHaXDorlsvZvO67ea0Bx
4N95LTKihwq+Gg2ntXb5CEI17o028qQs3iePyIAN9p6QvOpZXIAbZ/6++FJ8h83A
N/h2HtO5o1uZhgEw0vQzjq1c6oha+sf4S2NHDgXR1hZQ9B2p650ZDjYlhhhvhCVZ
cAPVH03VegOBwAWoaKZQlUfMGSTlrr6TjfRD7hZfeGFIb47/XNYptwFz648DSOYC
SJPUNQL6VjBpUCQgcQZb88/IlELHyy9pf3U+Vq9rXb/GU9Zime4t9jwzh+kQPDok
mfJ7G7l68ytmlzLBUNBZ9GhDjjyIOMpZNtzOWM2DdJtuD1IGxHniRkCkdrCS2pjR
CmtxV9Gnb+pVlWqOp96UFRf6Vuz7bMMj5pYLEdws37WGseXcDDTyxJuotNMfKCI0
XBFsdEQbepxDzVpz83gUBWk5uE3oZZ8Pr/6soNcKIupk9CvJSAdthXU2vLQijChx
Y7NZANjPyF/R5hS53sXxIzYTEY97ZHC4HxQLERysj8bU1Cu1L1Ff8xoUEpr0Xhcd
OjRyJGwMTw+T6MbFyujh2SpNUDTgtTPiq6Em+SSzAwAGvJI7xRgs6gRBCURtwHN7
XJ1nAjyqWSRq+VHxgSQ/eQYu6o7EEr0CNiiyWoSiKHc6clIyUHT8AYVsVHVHxYbV
eKuT9wyfVXI+br9MCJCFlxsIfdJMUAkpHFN3OKOxeFmSRZC48oGWSFWboLeFXDTg
O+WmaGU+AGCDUx+/u1sfuflgyvvNtjMEvb+XBYN7i0cXt+G61lI8HvlPY+75aMLO
rpv5yeqCoYVQoOoBtwJ8hOOGYcg1CXdMXPaY1jLjjinR4tO4j8lDT7RqZ94vBmXP
j/OMhxTEbdRzUBMVzFZVTSx+ttlOu20WV7LzHCVLFd/d0rhAjyxcBCWwBiSRrWyQ
sUyWd30sWmkSeL62WHUrQUzlzY+B6Y+8TSfZnOr2kjPjO/4SX7T8c8Kf/a7GBN+5
FFO4XBimJKdmnk4gFwSJTtTR3XRYtRpJajca8iKYss/Az6SBYCZFh6XbAMOv93sN
pfWECvkIZynyZ3W++jI8M4C+uv4ZO68N9SEwm+gMEBe9mSf7Q/eDqxtWgSQaGDng
PgtgTW3dC7AE5/0hEOuWNlLIln2ztxiWhMeV0ULzgo1EYHnyfqcH8VQ+Hp4RKZF+
jXv0DYrTqZ8huKcomJ9zUR2tFu89J2LzUba2VkSa4a9+sl0hvtv7RWfkxWB4AOQ3
TMLtYMF6z4JUUmmGuM2IcPX7MjcoM7Oo78ODmSq7CIvHH2DgFUMjFK7Z7uKJJObS
sqyCOkBBThpqmbT3WRg1AT9FIHnZkM8cFUGaF5rImeNIBw1y7GHR2Pu4aMERTSCt
vlj3tshNYDgtPngtpLIz1kDeDtH5JpRafDUluX203klP72WvqoA4ToF29s2hF7B3
3oveWiNx+WI8JHrGgdfGgc8IhKO48gw+nt2NDwDTij08TzSimb56FlyuVn/ZjQes
cjWLtXzHKYmBdUOfBQMQIWH1zUbSGJU2YjUTtCeauYjC3WO3ohZDuxJlu8xlo1jC
6phMT0+mSqX68e/mUTd4XpNowWfFgApr/P8d3A3wzGI9d//oa5sk4xCpwMnCHm0X
Fae7CBvmT5KlmTybHNr/3QAvsW3sRCXKw2C76mswgV6ht3M7uRHsw5acRQzVPZCh
qUl+GnldL/i9+h2KNMKNTNwCawpbtK4LFCzYpEm8fGLVFnj+qA3C4wb0YutmFtZ0
RJYyyGgHbCCMj5etlq2mrsFYUpC8WS1TdXshyvNvRFaTulev+iOBbsU2jlt9ZTnV
esWqZxXbJsDS/Daa9Y/tsK4RuDP/qktbYsaNQIS6luoRK1c7K1c3yoeDuaHaUarT
/fInhPfVRaz2rj8Whhar+j+ZDvhUg1UjP1Cae2T9oMwn2lzmjsDrsmy2HfRujbDa
npdHbjL5R8dGfrKNwxdjhQovhDKvJ0+5lwF88oCEsnsFhWZvf8UUAniFV7h58T6v
VsZIrF1jNvrZaC89dxjIJ6HCbUsfAhDNAHk+zexpe+twiDs59xnxVMym4beruLwa
0IVrMOb22TUVAeMYV5Rud3LyCWrz4BeDL6Wmk2sFC+AaDuCEvmJzcq9RuTMpZeQY
7w5z2vxKXVV4Pwe2NwwKJWw+BXbaWmejgkNKWZJ30G7qKZScCsBbsI3nBOZPGnmF
OIkNgjHaR7gZIBJM1yoNQBG497xzH6F2JDXIGWzOhekl4JXCjjgupVaK02AcoFQW
a0hbHM7WT9wDYs4ms+RuWvONRIhg9axaOVVy18dKBuE9eo97KXB6CZLWG2cdmtGZ
8I2ntWjZyus3x2DR84HfGCz040+VqTL26h5VaIQNIlLGglesN0nYbnaVCfJFdN+r
1tBaLc3HGW83a8m6CPygs3tItL9RlChxHj+gh+sKOaq1SlMLMxIjIgr2eDOwpDmG
VXgnLDSgG67KEtTXxGKZCxTYedubsnmOxqDh8EiXX/pw0VtzeRIER7a03/O2Cdw3
T+hd60qiYwgtZ+YPZs4F2F/e0qKhwhLewz72w1OJZbJTWJqyRvTzOYYsg/M9kWm2
rmY6aGMz5yQ8dxBP2T+NIzhx4uIAJCoNI4eWlR14rCh08HNlg+B1wyMx/M02RdEw
seC+/DIIS4He57uZocBU1iFkEAe3Qse/gfYlDAFArik4XJRP120iLfYIDm64FxYK
6XcpULSfwECWOLYfrlIh90rySDLEO5VbyELRd9JtbHeMU1R5KUDaDAbiC2xyNxQr
nwQ0trZMThuPnysOnIFntxHfhp4uS+j3sTNX3jPFuwylxVUluezJKkJLWu6AJGeT
ZaOGVJ+NZSmBONjYV5aKHcKIRZ2Y/lnnIi7BHCOFJA3s9njR26+juWCkZBOoY5Uf
OCJ2gxqXesyoHMi+4xRpeZegeJlnf8o0pU6pX7j4cfiEahfkj4ZOw1QU+IlSHVM+
N68xhZEhy4oIdX449nODSTBfj0BKm7p79HNR8o9UO/LOKTcg7QUSIcKfSC8ZY12o
76yGrFjdr9wlfH4SLeIKL0SZGoZQpYaeZgtBDX1DQtGH/dW4OrSRQhkZkfsFHE7B
Bi7Jrr6DBzJK64R/HYz8DHWAVDiG0BY3Doof5iTReU8C64Lf2VlBCqVNoDEAffgL
mxsL9oaBsRPu9KHbNcosgxPnkRLyJ+QA2KLbm+QVeXzDEi8TG+fxyNDUaVwt1bIj
N0HtHyKvPALFXJj8DrvS4mZICUa/cGnejadDQi6fjT34TjT4RRvEvO/Kl2TGGRkP
6Alb8+xLM4nYuPTW5V1+EP6paSqXOF43CbZdCqjrpkNIqoIK5Aop7yMKNWl9sVSJ
a7rTnZSAAKdzDNjW3ZVrxHqUhqGUPvG111E/944hEMGo8eS1wo1pYMQVXOb/7N4C
YLRZMnvcD57JFnv6AlBzrPdTmeJ+vNDa5uC7EidzT+ToAg0geQI8ap1Q07SHRjWv
5hQdKm8JwTAQRFYuPynwnMWRVPE56IInIx/AK7z8BpuBOO7Kji/z6OCuO/64L7NJ
apd3kyj3JNaedxfGDAC/W6BO24JjoJx09HFBmVQ7muPQCVyJgNPM20ds8R4FiNK0
vfbfd8HoVsVrEMISvWXBmzy0WrDlwdLE/axBsMccvA3z1BziRSFE8gh7ep93CaeO
Z8ecWOmLwwYAaOpKVIMExfMyn/ZrCdlieAwup89gJd0UXbgHQMqrLgExShtoAWx5
frEf//QDle17kcmWcA7R/SBm0Y/se96iI3d7gLYtPdf3ZNz7kfgtZlCgvoF+fahI
OHxWc5/6QYkb5EhhUWA553hTa4lq1jH85cp2wHjBDAHlWQwcZYGZ9+zVnmKnPw2t
36rRTaGSCAgBfWV+oRje1tIkVAl+oViiPT8uQinn73wFYlPAt4Cu6KFeLgPqD5B6
FcAElzfKBtJBNy4x/DF1vcyCYjkfgqI2KgLLsVMoKht771tErY1XOM1YQtPwWYe6
jsShBniEk5cAvJlxXxISFGxuXK8YvUZT0R1Kg/d9MRd6CLd5NYiJuaS4E5Cw3Q96
gtevYme0ZGi29DE6s+ZjypPEwocq8dVLc0uciBh/3TNCeHC6sVCNAgpF8JDPWHrE
RnqYdhl49j7VHTI7s+f2iHpbl/L9fVuxEu5yo7rz0g1tmxjKSEJrTX1vvvVg+Ash
XEEsPYePqmuI4vQrldC9f+ru+NU1EEtYZVpxArL8QcD/r4j18yNNsyg6loGqornS
zixiuZKWKeOwBDuKLpq18lvHOaO7vCGOitVhchlyyL0wxmwM/g23fqPFrvVnIfb7
1G2lUKK9k+fGf8kKk5JdW9yFufO54cTOrn2N4xGopUYpSw0SpeYtWcC3Aks8CFqV
kQ/wlLSHjIavtVjvNgZdds93jyJKpPlXgk/w7SjkfBTt10Gplc1I5Gbh62NCFgR5
k+/UZibLn0ew37zDVJBO2anATPcVbMSHCVZDEoh5gTntkE4wezMUGq7HMYihjeck
0AiicrEUK7ciaDDYc8OkTKb+f6Nnm/niwNRRgZ4ZYOtOMR9RMqXOxYG4Woq/mlym
BJkE0GpoR+DcHb3hvzCeGqDC3AagdaVsuRYE2fb79ScDyUY+B+YUDB/w95mThx41
dRILtTQRWmyR3AV7pPwOJWCnEDsovdtJKaHuc3LRo185ikuaLYIJNW8IgGr9sgsT
T2ropiZJATXBQ/Qiw0r9tg+pNv6Wn9LwWi/T9Ehz1sWqhxv7P9asZk6nTA4iJIVB
0W6svcwCtm55AiUryW6ROvhJZfRTidiOshbT6t46wuuBR7XQgyRtcp69MstyhqIh
vXqPxqUbs/7GZBiYQafRrdzFqWYjdZQBr3SGt0lMKORiBnZo9NK37DvoTf4P3DUk
RIcG2tevxRq/bThKZ8COyzhKps2BXSXE6NxRfcOn3+kNDN055qGcIBmReDvf63ik
HylRKLZnurbZXIRuB8oRRVQv226LX8hKm0MIhgur2aYACg2wr+GctTRenzXyRqfQ
uQ4aQ13VqMdkRUfUDjqFdu3Zn3TkqKlwENc3gd+TaAuaNQvYvGvEhEA2mCLk04i7
XdKDWzC+ClezlnDfX2hSH2v/jNEI2/hEd+czacOdSOrPOCIiNZL1qI6Zxq9r/MWc
jTeXB0UdwQxEVBtxHGOzpmNk7Z5TXA9/vDLTXoYNQCC0q0DN7asuY89ZEdZcwDoH
/V3K0ffnNQdWa0owcRh3K9hi3jt8ZX0UDA946QoatKCNBtZGjj9Ub1uUpKmiEzOL
kw4BgcvRytgbwjhuqWdYU/secvMbgRBfPuSCH/Z96DZvzga1UArGG4q67EPBAxO0
ZFl1eyA1wkkWRdeWcCebljMWUvxV7dxtgQyj8v8Oyt76Un8Md8mPfUMoAE+C+Bl8
dyBaKIPS3WFAdudiYDTJozg1LPiGhx25zP+hamol6CvuwctY9Kas5hqzRqpxK9cf
3nvJU8vf2EqQEqIB+ozm97IxsfvK/9eND7SbxHOhlMUaoKBPCFOBdMhcySVRrcAd
40ykrc9PA3iKrv18y9nYUXXBT9cYbvVsAWVV2QR7wYmAj2mGZKBX9WcAGZTD5C3R
yTKTsGbQdkIGrPmyHMTNHCc6sJRfga3EvcYQMtc+HPe+o9vQgOZbpyZQaSrZvopW
y6gufd4SPs+fRl4xOHvPCBYS+Zwyxhm5t8D9sVkvM9EW+QdvpFFwByHC6HOxD1B3
YYE+BD+NrlXN7reYbRKomLzVq40bNXc6+FineAQaZhrbEnm6TmFQv5pZ02vpMaM1
eyY0sKZ05kkuNTJ0dx4W6ob2sXXiiBFw8wmho8/gKOHtGmwZsdjNYwpGSiuXtAKz
i/qwgKg6ffq5As+fsVhBONqlSwhoV8I8oV9fjQnyXVCHbV5k2CN112l8vhfebxPt
s2NSOE/LcInxFpjxV+qdkbt4EI3FWQ1pd5c9YRsGyXkOYndW+VUWwT+sqEY+2vFs
nquyBeHTyYz2pEdMdJYP2TNJQpmICp15yoE387aGsV0u5YOr288Y/KiI8whMIblw
pNNFpeL2MdE7LSthiPRCCfAbN850UmGKPQuZbhflClCcrT4hFX3OekX5Q+Ie0Kzd
rLCYFu0uzmzts1+tTrcgAp5z0LCDWNh0Ory5WZwDeoYYi61zcVbattK6oN3Q7pHs
B2aPLutVpEwXatTlO1j/2VRPqWkiVdDkCr5mbW3jVi6ORPkw8a4VdO37tHAIzlUq
xVg4X+zEZOC+yboH6TOw4CEuX9c9G7u8eYuZDga9dVpV2bpaKFUIxogKISNtVpIC
d4xVs4VaDZRACf3vV63BcHdasz1sKLtIOKi/YdPys2mmdJa3ULozmaANFEoWDVvT
BRNCAy9Ct/adNj2HYYwovLcmn+TR+iT1ccob12eJ0B0ik4SHQeSn29BlXmdpIzt+
23kQNp1DSVFsKnvuDMoCYo29z7QvQ1whpo7mEiWQjv9mSq4qPDfD7qHE0f6cBc6B
wEDHkwGxnDQEtevye/31Ykz4YGNXwrTKad9E/plmvXgrp7dsIpMAtvEg0vm1nxhP
lWbbF3A5RKjvi+gWozRlvMUfUKgDaEOUtRO29tbLDnp2VA8FdnJgEUxEqReEZXtZ
Ov0v/IaP2FjoP7srf5CrJnmeqimoFk+atD2Spk78dtjbpncCoCE56ycCcr1t9mmL
ETTYId6rssGVoNuOiUokUo5f2PxddPM/WQGeV795mba9gI9Vkznub/s7KWCxY4Ye
TaxuL3OO3VnYq0iVH7Z/6ozc0LLUzUieAzzsYOUNwznsaDLn+XZyVEZNmRUIOcy3
HwlnBwpZtBl0cU4vkk7pHenwjGQ8MwMC8SGGPf5eqFSsx409m0FKgmXQQ7fOcjgG
cJRE2I7XtgUF4YtoGxQFw6nszc6dSNfb+RC0M/CVmw8M+/6s1Z4PTKmmjUTJE1kV
rV5HMs2C7jZPZMtT38op0479prwOIERR8IcFVBKEqvm+DhPbSWBmE4lVlxkCM2HW
8ly/2eRxGG//L1axP2tNpey7GZLnQCtZmyaq9DvTZEdC4o4H5IvytoAZlK0yC4Kb
bwPaYukz/Em+JZKJJp30NrZbSLasNoP4xP/b4hPlmNdXV0DmIs+dH22SHmKW1zrq
myFCsVzgmfGyBmERed3q/58uo400zb9iPmxQdMxJUf+vMbhQ9i22SIzJh1Okdgkq
KKdUpQbXb6glCny9VAQbWLZRMmFTmnIM93QwL1JyEeKaYpdnyjptddr5FFiV5yqD
IOclyiTvWHM9LqmCawY/jb3P7mLVypS4keYvDOF06lBK2/FJbW2ipBa40Cmbnkdq
u6UXTICH9Oc9k1ekOvCxek0xwf/95asUpje/ENQYIj0r9DvGzd1bDGvg2gm/Zt9R
wh1YgDdTa4h0Xot4PwAHtc6v9nOsGoEh8YtzM0Sk+S3+KEQlBt3bJR9AsgIzZm2Q
/KDT31YCULh04k67NvJhhcvphl9oPn7M38gT4szL0aUlq3BUv3bhoo09yllZBn5Z
qJZ5v04c2SaNE3zHYgKXdwaIGC62K+mTve/ZXR7oTpBFhjwttILuEhDYlw1Yv1El
afK28JbqAB7H75MwK0OG28h2BcGChT1vuZXWaftBJxEMbZ3uCMyM3pg7GLbyJdxN
NXW8zNr4AIzCm5lSZUGOf0YyTqT2ddBTkKD8cM9yYXgawjLo3AwFydv4u1li1vM/
JuuJd+38Cqa9muwILhSdraJvMANSQ7vZTXwZHBNbgo4y/uIT5e7EIPm9ctW83LI4
7Eq8wv/+lvkYRniN2UpOKP1Dc9Fc9fYQ5LCbgWlMOLT2ctwrOqKFJQ4oxVFnvgQ0
1AmOHrl45CMF2GfqPQT33UG5/YiF+nDi3OA+uwTrJ70WLG+VRL6rz5UJaCxmcDli
0dGtRgC8HnDEG8YurOwhLCxpwhaQPemQ0Sh86KywdXZd0Xbm591bbnmwqm63ABJk
glggiOtiCA9/4OPqLbpcYtxg4QMv4qhFUrBP1QRclPyaUH2R0gVT66tiEyG8bxFn
WR7J2KmOWRybJvZON0LQyCOMOAOMhZ1sybtxV6fTggkWZoJMl5NtEY2M2iLUBXVl
FEyGJKfAe4HPIAOe3/AGxwb7k8kfFuNCvfvuV6SripRl8QB3g85r6umbJ3E6s3R8
Gl3tuI7SJ0cuEE4CRsPxnxOpBHfwK6lUj1yPe/Ed8zS9KBRhGMoBaYCEQhK4sdVO
1uXkHaXhw9W03Jtr5scYz/czzj9YnkusvXLvQeTDGATfbzbuuo2bKdxcdv+H6Zr0
e1rnFsDL8dG3UxljC8J5ZXdUdTFDrxWsbsYoB5mOkg5gR8+PO4kRv+TgXrPLz/4o
X8ZVa9QXRnTREHCmG6PKgHRns/tXjJzS1boaUUygZcKyz3ifj3QnJDXK383VEabq
cF1tEibx7knbOaqQV79DcNSp2vgoo9vB3utqyJn98WJf0xVMkRVFyZ+mRIczzMKX
MFqBVBFoW6meftlCfR19Kkd4znecXp5Ux1ViLq7RgP3ilBLZyzVOse8Q6ty7mXX9
Ni6EZ+exmWD3oBW6JZJjDXRuBEsZXhypuMU2ahCBEFRsFQW2KywYc2VfnlW+RpXL
OL6t9FCi19b2O5MSkZ6AGMQZfrm5j/eOP0Pi8HaEu2YVj7fZdn+E4/3KTvNXKHSm
pp5yliXIFlbaQLqy04805ZVqA630KAGC3R/XycmwSwsUIJ5We+1Jibhj/ThC0r6Z
F8tziOUjwxUh2C6nlHEyX3OhDxYrc8+6Xgyor6OMsArqvQX5IHFnrEp5DRUGqNxF
XJOqgfat/smcjRYfikwZsUGnJBRLMg9pbgTGTb94k/6q55mLJdAJ2F+jGIYJ3imX
XNLgmR/nHjDeSyTDUoBf79tuz4L7nkaagdLglwUzibdzQDbgrLSe8GGC0zeZhjJR
5FzUbsM6lBWYGQWLOOLUtjRGJJCWIynt1wYCpW+wlRkN1K4gdIVAum4FiLsvUKTp
jiIjDJc/vBVM5YcTjlxJbO9yPEqVpiZmS4FgiNLXTdERWrYmczZD/Yze5wwCIz1v
m+VnIVDPS/U3VyU7xfUfq937wh6/UopDBu5kGYwpZU/MTYiHHN8H9l2j4Z+56Sjz
u4dSG+xIWsIvWHieHOGrQUVaBNBB6yOU3KV0QQLCThJt0SrCMjut30ayuw6O/g2J
L3RzmplkIJ6ZN1yb8l5lVxGL8qPRK7zHrT91ZfnqUdcp89oadI9WZ51+Imj1BjbU
CFk8U1TEFj0C9i/Z3k1pDMtGirIycGRBnF+bN585onaKO2SxSjmOFxyB/dmMKk4s
3spjoNQhzNwmBzyPmDDRmqhzOmxv4PIomGVEqLukW6lZchxz1o3xWyoUR8hdffmg
1z0RfVi28y3E9yGuwNIAdMETo7S/XJqLZQPZMnZZ5L4fWWSFYjiF+BwlYYjuV8+n
6OEgj/JliObLpHTr9VLW16T2AzlVyY30XUjBGAzHa1+MxIpiGNWKFxNTG5VBC3I3
cbmvIX0W7zveDs/Jes9HJTesJhqCyc53gEhJNFjmZHnXRkGrK8vWm+Xu9cFz2wVj
N7alkStibr6BsXNVjPJk0wL7FF0/xvmq6vUV3eiwwzTnp1COKV1GOkxNdML/O9UE
zkGIAi5RFzmApvrPtuqRESKYW42iMUFm6Qowp1UCRQzYoHCOQLH5RqkirE+0bGV4
TA7ZQ2o//MKNh9NxRVWKHVI4MmWLWSjKWpCiDD9tL8w9ykf7ULuS6SiuY+Wz//yX
1BfwyXHf1Mo4S56f73TYEObv2c/txJjJCgwSNIRznOIgHgvcU1IyrJ3J7t5iMIhF
aX7OwX6WTUvd11Lz2FTEYSCHjHViqCw7V/WVDmYJcuS7Okj4+ckNJdrzamqgNmNZ
p4/FEuaQ6G2VoYu236ovVmV5JjpPb2Ki+iSjYXZ9jfu6r4tTWGq7NurIm2s9u/NP
owLosrSRF7xnVW7/xWIcPxwc3eekXHEi2dEaRDuOKzb8tU/jB/Ds8F9KJZpBo2cf
WPJew9XaWwnmBXCwTRUYd99rehZ6FB9Y8o3WbXsQvJp8xrOix9PY5emG3rIIBmWg
Swqq6vquHiLw3T/tnrj4IhoiW/8YnHpRhttwwEu59PwcdiKMzXox5sYIwPSNUSNQ
SBgWQXn/rB5Sifa3e3SVv5M1/bSWwYkAdOQJgpmuS1rLIlq/irlgFL7D+puBxYsa
IdWVSmjwgNfQFhPXEFFwvqfoZ9HgCJIs+fi2Sl5SAUFCcnLu/Vy943cFQxfRxT/S
Mf+FX1M1Xq/mcXd2s7ddRN9lVZW3W5vjtmFK4Y14lzafFoQzJcafIGTj3CivOLKs
JjaySbOveEtl9bi97FP349c8oRafcsfIhpSqiJYPQUGAqXWi2+Pufcswv1/U2qV5
uUYG0W+cwZrcY8lB/2VLXRJ99KsDHZMIeM+31rTK/KSQa8bSUguTJgiP7mR94PRB
fD1fmPzNgURK4ak6+Nmt9KMnKhlkn6Q2dlJLnUbO+LPkRS2DY1vv4po+bCGs98kW
rEwLqbXhaYFWMmcPwwNA3EVsle7Uga6IEKaSwm+y4XDj0sqv+6R3Z59Ebip25HXV
OrBHKfKdPL3ASvNgI8P7nh3VG+ty8gv2OBG0sva6ejIlIdLc76kEIY1qUxET9jiQ
Z7fpxEefl1U3Vdk4zVS4aMG0DFYFeQ5v8+j2WG7hkK+PpzcGmA6f4RpYqoeAsE/s
zbYhD2S1X485Jrv+3hAJ3gEMVQyI2QEadeTh4AeWdI+8ANmkGUJnabvXFBWAmoSS
Ehme1nxP28LYb/LfW18CG22db867gmX5JQrZlfdZWYtCuIFFc6XoDNFBsa3e0wpQ
AI9KCN6fLgi0T15WtaJIo1FgI4Jp/xJmpqgdcSgfFqMWrtURJhVj0MoriLYMdxdq
ql43kOj0w3ZSs6K1u4i4n76zM3cWCvFqjut8uixW8TaSXwy5Ffd+srYuk4aLmlOU
pPI3EPTEqbVd+tdpkWflU08m4MQ3lNewOeRACag0/doP0FFJnm7TPb8UlXLCukK0
YquXPowaJ8860bqIkDf7Pa+ow3gsrZPm5PifXFfIeApjSKyJYGGPKn1RDMvTE4ep
ML01LwXuQy4GChXQdaKrxJOoAGctU/6IuuXWeaoTynNbdli4FdgctRxqR5iXj3hp
otR4/Y0h09BofQd1Cul4xWUnAZPGPKQPzghEJXWK8Y9nJv4IWLgdbqc4Q2XeOq+I
bJ6bela5swYUgMcfqymVwzRRhzg9KPHAGL0+fxlOHPPpgwyo+k9hTN0AF5PCB06f
6M6RICvILBf1B41SLCPKbJhoVJti0wOw68TGU3nFpj0R4KEFYETbB3Bs5O2G0RLk
7HVgWmTjaxX8FZTy34ZyxQvTE02wE5ndgYzh+qh6Bzw++CbUUnFhn0OYJf3FLcfJ
7nS+EvLk1/Gh/05tl3cbLVjJCFAxB5OzAnwxqz0hibE4doK8PYyCA83ABPAclM+a
WAtzpnkZZkLeq3TKggpa1Dfh0pllucnMzHuRQtDqCGZF6bXRTNoZy1qq8vjrycz9
FuZA32xCfom51k5LuFuAZ8waw/2Y8ni2PXz/NHbX4MzSB2vwHEf+b84aIDFQaHD6
vWotaShbGH8Nump9o0uh75qC/JyCeYXEIqGouMauvsGg0RaP59hFsX+iTq3yfPyB
SaHZXUslZu4hc0AZAgEun6FkJaSIssBd2RIRnLrdABK4oRWtrU6nZrpAvXltPlre
zACO+YCBjACa0TJ2TNI0JCzlH8rtYZFIAfsptmlpB+jeJTTdao4o3FQcNFLX69YD
IjwDuq4JmLaKpYjy/Y+CwPqMNN4Bv00+mA9CC6CvGZMi2FQK3CdztxjHaLoZd7Fr
BwR0tTopVstooZs/PQalTKDebpJ2YHjCYqZaLlR46oyGCUia4au0l5+rAm6+AegM
c/iJmkVhZXBFZjhxfn+kcmUpBaWr2ZKTmLh9AGJQwygQAsMAiIUIPaupN7bn1nFY
02IzCTlKyrKkl34yT0mn+SW/CxON3Js4E2ArTM9kEKE5rwaWvB8NRV9N3p1z3JGi
MGZSyykgn4h9VdrrHAR3+D4EOjIbv959YUDXj86c4Ji7Qrs0wLIjW2soAnff65Db
gkaMY1dw+l7yUWLGWMnaqPSIEU4PgSIOvMqp8p/2b/z8ggq83kVpi+BTSS+n//0Y
BIY8fSqTBPZ8RKmJOHrBZ36zEOvQZqMu8SvhdGut/ZOOWLmHdRfEj13C9nvE6q8V
0tOtAIiqZYMOxHvLe/Ow5L9JvtRsKXu/WrY3gYVTKaQT+Bay2nU45SJ810+xQQD2
+3UrBoTB/zMTxOizWeWDD5m43IrF6zlRzONdHlfrKsNHWyw2+2aDMlsrkLEIHcSg
ltXF1S16abrAEPxc7h8SYrqsfyxoSYugDkJddHUfXt1aN5/CGTDac5fzoY20wwAl
BKFVabhnzYa6sj7GltbZtHEkcN1przTYGCy09v/x+9unvS06G8boFzpjiyuP3KIJ
rFDJNzwp5SzYC50c4iCus5QesX3uGFSsR0FkydIMj58VHbEQRuNqKFdGUGaUlXBf
HeQWzLIMo+X3Qv5xgu2LCHWFo3TZMiH+yYDBbAxXVNY2xHNErKRAXJpWETYD0DMk
kKRfXhsLoo3adbO78D8bkYwZgMWEnkjm5Zkj9MtQkgVH8Vj0R/UhMLbANpbwyevj
6h8VSap2Vpx0ZSbh0LmqMYq9t1/UZm0MbDAayMrYOLYl+vGsl3ZZrWP4b3SlBPgp
s2RZ0yLrRJYk3iNb9YAUHeFR/vskcEo5vddnXzxMQ2eYBXl+39vxdHb6b59SWfWW
BgnaJ7ZXTeMtMDwk5NnNE6yeyHzCT8tReR+j6p+8IekM0SWWkQf8wLMbtduXSKan
b21vFrduD+uh6kos1sReyDPzMDKPnX9eWh7A5UK/9b0+WLprejaUlNgd85iqoWJi
bSO7dpuUt3yXDuVj9lSGSB6DTAoSrQeCjRcYIzM9Sv5bfdsZTh09PbVjTtx8pqHh
FZ17OkFXs3hlD0Ox+fWeFtR4mkVEcg104f2zbW9/LvoVSDZM8gBDYfGRKVSqqPp1
+uDpSiZ71/OXagHWV/DZNi5bTPWwtDqnY/ymO2Nr9bBfjBJWzn5pFopHvFr6f6IA
CWjcBpbfoiqs7HWqJ0+FVTpzUOJxUY3iBYDFj85FvaKxZRUhzaTjIyYoJHEPAFzv
dKLQApn7xXMF3Gy33ff9xcZyFa8R1ecILW1AUuKSLJngZ+yWzsQnCJQk3cK6w/7U
zxjRV34XrruM6y4Z8havhLLZlyI1W/lKqDYXAAZjc+ul4MGYIAxmpYkPBqnUTd69
KlkmXZ/nBcqbySXZBvh1TF8hCQ8ZhqOxXIQSKIj6GD7wZsXxjVZiuoUQvzm6i3Kd
3BTKfSzDJQAOQMiHog+2LGlCarJ5YcVixL5T5Mre8yVlEDEiv+WDUERKMEKOg73j
rK/wwa4jqiL0ZRrxjesPgqs4n0KefZIz1DFbvfeAYw4qG/SdTdrIV2uvit995BDS
syW/srJQ2ZGcoCf0frpGzfxB4AE5KXAWABmoXF4BW2TfbiH1hBymqscw5yAbKTTj
aNpt4bftzUMEROYoe/+Crx5JC4BNHkrVXJvXJflkC8V3A3B+h5b9Q1GepjE46/JU
o6ew5pU9hPSeA562O+LCwbViKEpbgDFBMf0BjCKarC9ay412/6Shncg5sFRGkkpC
2FLPdu00JKW7kt9Q3kpEnenrZrXEa1kYfjYhxtiY1SjODHSQRgLY20blqQKFmYYz
aLjZ9bXkoGfGCkgKD1XXEdneP3FDDkC4hOnwJb+hBXABzZ2mXz02R3IQk+3PEoyv
W8Sof4apJMmuIzL5iov/6OnDeQBG2063QvP3ZzXbA8qO6I7yXIL1XpyMM4CT4lNt
Q2+/vZhqrnrTKZ+Hin0eSbHvSnE+Sv6w98fkWzvDuJl3DhjC4Adlra9PzADs4VuM
cvYqC5Pvy0pUJwi3cTwbmGhy2cp3Z16aANsF7pmqkH8MfPaGJjWJ+xTw9c70m4Vt
lm4BS8b5gKCqobls4CVjGsSwW2gDp9m/F4hW+pP8/TqMx2009pGk0xPmpzudhUUv
rS7Bg2K4xO7jewy4V0cC9a0u+BNXk3JvHXuxB4Li/JAoFE8JaS0lEFQ2NnyvbJ8c
ebpYaNdyHw/gcuu59axrXnfzrQnN1zqoWxEubIHiLzou9oLK3dpnzHLKvmWAX6CK
hWhGSVyJvP3ZaL0A1nR7QtoIHtrDqIgpoEj7yqnGfnO1lVF1NrcjrPpvRWibf/4/
IeI/1UKF5vuyja5OOWJw4t0Noq8TADkaTVrzxI4Pqh9gBa6Nq/YhC96EA/1dd/dI
xtvSEmF+/yaQJJ/Vo5gHRNURj87MT2iqHdOuH1hoQl601pD2flKgQTeYXTFS6zJK
8cqgXugkPRayLNIaLQjHAF08xD8BycBqdu9pN8I/thnoyIFy3BvI3iUAf/4Fe1qQ
D7/Vxbi56NbWNVOyIMYCmr4PPFr39d5ZkX5HawsFnRtViHOb0o+AIWWKpGlIyAUP
r9yMz2/7nAQ8VPyJjJHpbM8UNADorPkP6YPdHZvULRf7LRLzS6dfXFgaL36hAJk2
pfDKjsQxqjp5P0m9Lm27OrIGT7xHNFDZIAWhnf+EzY/KKMXeh5MbWNPVtKH0Pa+z
suSzIDtPgbm8ZCVzvc/6Wrfev3xIOgneMltGnbUzjUMakzaBdo3Bn5+NUBSE1Sof
BVaaZpijBLEAUgV/FJEURBym0NmzBEZdn94I28NQ5JiatGAVIkXJ0BWPMNVERIel
2w3VB3YPf6TGW9Ft7UQMXKws1UZZYYENEd19sJmlhygo7sqY57A6HoCI1/oxh8AP
8wmciOVVTwPX8ZhupMBZ06zM5Tffxr+b4gy4Gc6I9vgu/Tfdo+sNeGuZqN+7+PHA
aVDlHIIzT3R0drp/9FKr+Qy5gLXoxVT1E+zMgLa9Ta6QdiJajdabu36FIO8RgsXa
trYhH9e7066PuQIGfoszGU9B4xqjMuuxlzHCa3iEsow/tdRMdiX2mgBg4MnHUI/v
QVbYYLVlke8ePTWMeuuACVA+ttzu0OYJx4YncfRzyo5IoV7bdkWIHu6UzmZH6UmV
coDoUFbRhdbNDOUfQWC+1fi9m5dtmyiBRbQnNvvYKCi4oXvaY9gk/WK29HXRkump
w3eAfDNThgUqiXXF4V2sdx3MwgwxDmKM4cOsOUQO5qYOFwU2bYiBnT8N9NPiocx/
h0UaC2LRkUHyHGhDtF1DDAFWd3hTOo1RTSUBSLd3ul5o0W8oxmB9toz9AbVD876y
2hJkmSlPu7NlWTA47IHxDBZ4lPEOF6EpAvrgEEN4rXH7wM6G+D+tHGOT3Va00vwp
2n5ovO5ozINjlWrUciKBhDfT6B75jkN/VbAzAS2To71nVBaG9vDaT8jdGwTXlr5D
A0rDkakKiEyg2FUJBrsJQSJi26YF4tGQKl7FZnwl4hcElf4APgrZuF9ypUE14U0C
7cKtJzbmvj1tr2tuNf1Wj3DuFhcTdLn69ioNUHO3satE/oMQ9JZA4NM8Opn+5q2Y
aTiXq1mO/RXk5XusvFQnyOwzeMrU8m690jfk0uxwYskNFTu+ri/furtvsqDR/LhA
FGEECBe7zUsytVJ6iucNmS25MLA4Ez2yAPZnyjdVnoRq9lEv0eBFtuY11qbd8o0D
P+ccvFq9KHPxdafwarP9kbtN/NpxUFU+7n2anJhqVT9qbfUyOdeIsdobTke1vnF7
s5IpFRPDhEAWwZPWlmMripqGmZV5fvumTsBhCMCzUAH+fJQIdENqDXMfYwljc8O7
DXqB/SaRzTPfFmzLrqK7WX2+MrUIltcDkRWv+7InMQCg9TYGY0mzeOxOk7AyFuMJ
jBUU9ngrhfVecOUW+ZUWQveUHVIQxNP6t/yWr/NYiDXT+g1RL8V7sTCC9fpZHupo
ftLkM8l5XoyHbGqvJlU1mJ6fKM3NyABQPwKGKQqAQWsTprrYX3Gv2l+mNEIZFq/4
MxtXSiaZVkC/MmWzkWn1LPKUzqjU+9qMf5cj+xj4v+CEn9tkX/tKHS8oPcSrqKN4
AurGUCKijD1qArT3IdZ5OFVmI+tJ67NPxVHfJnUhCjXZC7LsLF4XDbC/ddN0QLAg
mgOGrLFvo6000NGA15FAeHSc7xm37L9lAp1Cw0N4xc/Lg9XKYl9TEvRq3oZgHAeh
/xIVZelpZHQQRFJRqiim46hlAH7gxxt8mxagDuJaDs7Q5jyEWnHifPvNKbi3HJRp
OOzC2HMsSqgl6UzKHtYNTgzM8dK5vQk0LuB0dYQ9xwMveWzhGTexCEVYQRbLTKbS
rENUslJaUb/h+3St4JciVn36bd34C1opjQRb4s2CzX+y+vmOYR4ujI5ilDEQ6Pwm
Cqr1i7Xodj3pnyn2qZIxhKiU1BhxlF5Nq4pRySdYw+VzwPy2cndJ19dDVEXKUnLT
aTnQiQa3+QbNixslUKbsCVEPGyFYmphGCGc358+WTxM4lr0RrRkcxFqnLJ+aO0wT
aMYU46LO6EpQ7fO2xav1yzvv5937EOZkkB8v5OxyPxL5gFGAM9q9NKvgoW5rncLC
knC/A+Gz6q89NvEh45XNLX7FYH65OllbiDduob5QmRk5jKKdefQ6Pm9bm1RZ/ybP
CXIu4VnG1Wal95Gw+o4Qe0rbTQe1fv1JZoNwlR8RWNbo//17qLB9UOxLeqvRiJZn
jwUGcEYhJaAcjqalPN30BdIoICicMbXhWDO7bnctIhjKL7nf+svIJDTIoMQf7bTU
DzgU4hHEjGnQ/d84rl4yeh9I1/Qg1hJ0EYA4xXYvzVdxMJl2xgy3/2wQQk+b5kiH
eHLfJLH4nYzKDurrzD1V/BRg6zyNcfXQC5YKFmk6fXUy4GgVcQfpHlrTv5jItzf1
DZgtINFEqnUz+eeahUlGuiZiR34v0cEkTTJPtcGuEw+UOj45aAlnV6Br3LVLGmTC
SNqYZea9i90k5Keedw9PrfSHsMGx6SIVF44l3u1lNFT0NoNzACOBzuIx8J8yrjxD
BfBrKIppgW2xi39rzL6a3EWA6P4EN9s7ZbJgrDwaJ2wIzAVXgYoaoDHqg1K70thu
nhb3R/TpkfmyE625gqNdYrsrfL9Mqo1jaEWqe17k2VoeAi8dhzgSX9xlIg/htcEm
s6MvXve7qRtFfILKCX3mdxr00klXhkoboLuZtlmxkx3McLjsRVD8qMBKHsaJH/0L
M78FkYJEU9rP/BRw4Cq3km4UjCCSqkUGMFzjM8xmJNfzNyWqRfR55hogwxHmidzb
TMi9H6UQbsHewik8aa2AXkWS+Vm9z8pAGIhyAsehQjLUazmDLfsBt1BkUb5Vr1fh
3zrsW/2GCsfuoN7JH+q66wfEjqLAZnGAvqoojwymesKEc184FhETZcflIDXkWmhB
phuHKxbo8fTuro06CjiLGxFqOrJPzl5+JQ2Y0w5PFd1Olg63jFiX0zr2g1uaj/E2
q34uKj7w3OpjYo5kXpq6Co6iV3vsqH4EOyuRCjup0RMpTzQe6QCKOLO8o8wNqSqA
f680q6ehOEY05OC+caGUIYBwqmGr6nQJl2Vs12lDAP55o+gjUAbsTRoKOBXx3gei
qDiH+DcYydotfE6zsKOaOhrd0gBVzGku1n3yxw/Dx+qRV7sHKELxRuGrbiGm9S8V
D77EzzrF+ajZVAHqCkhsOhIkbBPL78vFWkU5/jAkRwW+SEEx54vznsdp/vqSeuoM
3AXtlG1iAfIwxLG02WQNDEDWm/d/w/enYLqxjpRtCDFhAsivhjtjvl3oSJfFRFZN
rkpLmmIrKd+m/hggSj5le0oq3LkJAitiARkSMt46+Tj/M92UojAH3pVRfunTZ+BU
WGUHVF//Mgvq78LQS9QefOmIkDii238f+XrmFhSrxIfiqvVSduEOKmTq1HoDyddA
y8hhlGiLYDqHqshHgx6sZGFw0b9HK3VdhaNFDlCUE4XP8FFzCM2wXUHbzW4fBzIL
XJ+lIyLnlE+cN2qeWssRlKLg6+I7arqEX8I4KlKkciWr24XgDORg31ibsT0hJ6jr
RbJqUplPxdXRs++49w7w8Yh84kbteMuqctl+0TCwHN/wpzgW9RXrZgNiCzzlZ65h
oahtBEx1SN+f2F+A2K6yfUrEOn5rvbn2ctBMkX5J32Sww4EDRQUY+rI2me24EENk
scSxwGXRsQrE2S9w+VMSKXolxoqu+nPJkv7HS0v25Hi5QJEcocJDNLsymf7xAAma
W6pdzRpMsqxgwcRf2yCeUqInM9lS0nG/Co64uvimJq5TnmS/aCN1Lsi1blbxZfLs
MyKb5js1akkBnqbOwMqj2S5oN/m4k851kVdDGicxBN/DfuCuj0eTsjPIL2nBo+dH
gLKFVspSTVZ4/HxIq7YnubpgJaf3oH6k0//0RIV4b9yThmVdBkKY05olNyu4ekYJ
ILk5PwzgMmvivpHSbnUrAp511T01igHhcVQgMRIYf3In9+j23TbMVs4DRmIYYU/p
P7n0KG85fpTxxilTk19c1lZDY0HG6DuZy+zVANGJHV3YFCdyjK+ek4D4Ttz3hWJN
x7XOUWkKmWID98Oo4C8RZ30uJj7CFHfMICVgRedue2U0qQhNAaxwzOqcVonD1+Pj
f6eXddDuxbv0MY8SKxFyhsi8geqfT7Q7OwU7Eu/c0vLF53YS8Sb6TqCIg3ahmSwP
T8T8z+z6FyAZiktGnXk956CDEaEjTInxVMIdnU9TcM2TgtACVa12BfD3X9AsR+HM
NZpt2l2CRYj89e/s6Ortk9bHkQT1OCjOFhzqTuJXa9/KNaP76WIlcMrSdrEu/YiV
MQ5OH0VEOXa5duuUoRYMBRo3nB2dyjvjjHWaPKv9d2uyfSoBTu5zBHJdLbtnlFj4
pl+/nXUWEmJtZcsoklJr7mTTq11w4qrfmJCCutL4t5F/fYqvZZdU8uAssec9289Z
LZn9c4B6XW1yx4teGVpj4qM1o1+GqoEdB9QSzklpPvdWOsz7QMqvXDn9TeJHYHSd
rrvwxrxcvrCtPpFtQl5pgCof4Ycer2fvNxbi8UDW7WykTpMY5C24ccaaAH8RETp4
G2d7qVrlw5eDUITfh3J3KCWcrTsPyt3ZL/wO/vOFv+olt8s7kZz22qj3EksIM+OX
IeCAS11qEXS2aXBGsqUwYA7ZjdIAoNwctcVfDDKUquEa5avz4eM/zgOaEh8Xa0WS
LdDdrQQb38zv5yqKtlfZ0gmyVWiz7fk9Fa3hLWUCTkMFuutOgibaxyqvYLOnTmNt
Olo4wsR6p3YFZAbbFINFYBA3fvl+ehCISdnDZd2fD6ya+g5YvKi7PDjLlHvvHwQ/
wceAe82VnZTvi1OQOpNKRn0AQKBtSABwkYLFC/2/ogFPxDg6e93zTR5EZ+9YnPhQ
AxD3II+EA4Ag5vlulWNg8g3MIlbazdVQIrcTIlkveeV8pMLAhIRRtQdMk5rc4OWs
VYQq90Gi7YFpqd6hSBzIHyBYWoVP5X7c/IUdp1kG4TVH9fwzUL0SulDZbyUIcBST
UHj94byyAdujZCziiKt6lWO38NSkzbwD8vGcY5jBdBDOm3nLeWvVDjXVWCv6tyKJ
l6OG13ZkYdouugHNkG3NEitUsdXk5TPrDrY7BiV49da9qnJK3/i1fEAkwxf/NdbF
3EZ4L4wYuCgBHzzFC9TNQDwPoMDB6gD10VLYLV/IxkndTsawngAP8p1z8fwM1I36
/vlaVLruW86MozKl5gVEZ3aNEeivkz/ytRzfqhGLXlNxuMNzrtxkySQxFJFBLWZ3
rcvRaFkUyDRyoE1SCfzKsupgW8jKDpj8X7IYiTJSsbu4szhC9lgpcPNuc1Cm91Z5
fsfL/Fz2om0YIKn/nyiOWChfWZLUyYxPItXMbJXrRwBy5sVPXpSn2MNwNZoVpaEl
Qpo7lKkSeHU93PDoBdExIfm8kPMaSKJtZCMRHD3eTorNiTWt2AsAyjWffuc3VauF
+S2p5w/kKiHuE2O6qNPacSRXeLLTkQ3qNhY++Dsilte2MA6+1rYYDIVq19UnR+2K
hA6a6NhuKrLl87ZlmoB72y8vF5Ul3xibIJreAZvdjlW46C3MAg42snkVXJLD1APe
l0eEU3v9ipkfZ29TCcqV+IEYFfWXApO1Mx0tUDXDKgv4j8VPhvBqm0IgLNY0LtGS
JNDFMIjpCITS/S5+OXbXhzneyaOmHz+5ny4llX//m7cUmBK9yriGQN99rFiywA97
p1KKFEnx/V7oXXMofjip/yrXB+ygJY3ClPCnItSgaN8hS89Lfawx5SlqZOjQeeKM
V014nKBepmNiMJbZ9rq9XOp7rxL7klbRL5gChRjVENMtON9uT5ZMkTj9ij/KUSVV
mhfzueFfiReojs2EYPYr+PsUTSZf4lmmcmFojhMUCv1/lzj9cE3hRE1Iux1A3j9z
CkEsXZ91HPJu5vbnEp85nUIlAoZlzbdKV2zDt/ghh25douUfMzwI0axdo/GuWSkg
oGoqlOYKiUqXZWyj3VVDOcLc4txAk3Tpu+B83cvFSDN218IH4mC6DP5KQIYRavDA
oUoFutDj2IuWRGvbNIvPEuNTuUAIwBgMzfPaA3+PyNUyaiwv+sq/kFYrZzoaECan
ZNfdBKk+VgTNB9W8jqt1fNEClmLWbYwULJd/bBSgtBNUHnEZOBREfWCx0Wt080Py
nIruqR2PHzuRVoPxaVZ/xhCcVFdsLStRrkQ42e9S4kHPuMIdY1Jc7HeS2NWvpoa+
rpyp0JMNFr08Az0Xxylpg7c5JTN2jeXLgwmiO0dWQcWBEzK9O/ErgDD8Gq2mTZBo
Ud4b84Xvv/wdTaAgfZIWgkY+KuFA9i1TnOtXRdt4xqofXOnutUJPdArTEX2iigVN
EMAf1Bnp9foCZ/dszarO2EDCDnZMXfiD9VLIMMoLyJJtohpQ8XDh12E8QzxYiG23
5GAjQ9iewB2gRWlaZzN91Y2OUN3hADMlSjdcT7Y7A9PFkQMJKLv0t9zIbCqsVtUF
yygjhRa0Tmk9Fat+Rg+vCYmnnnWKGRfqepq4BF6aJbUs0hjYMrEg4XJ8Yo2OFEXE
Fg34IqNIw4JmaBUwTtvBymdpDQkkFFPtGymG0M4Yj6fEIW/s1x8uot6t48hSKRpI
g5pbUWkILDkBsyOHlaaV3LNgrjBj+DAe4Alhq3DsnheYkiGTVsDFsIxBh50s91/D
1MgJAw7XnBgJOCrTqg9us6p/pQ90GFhzkvRTkLShSwXe8rZ+VmNmZNUxjVkj6ciF
Az71Q+poTwPWCtcOxIRVropL3SIErMw8kFe/VPXYlzwiWj6/bSJge0KOdkDtjlDO
agJycTKPJ0Y9piBMykLvZAR9KBxDcPP/YjOzOsSEjFfZHZkZHWxBFniapvIHnrnn
CbD0MQiriZP46s1VXB3NJQ==
//pragma protect end_data_block
//pragma protect digest_block
lN+ByFTIdqZoAtR8mtMHCdheog4=
//pragma protect end_digest_block
//pragma protect end_protected
`endif
`endif // GUARD_SVT_AXI_SNOOP_TRANSACTION_EXCEPTION_LIST_SV
