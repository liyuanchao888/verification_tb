`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Rxq52fbBrhTcguwOmCSZpI7HW8yMyqypV/l9kWuPD18LJ73uYF4kLJOMQRwFUA0i
8HbNdp+V/QQsxVnSYS1tFikUXot6UmEj6nYbSWClr8KyubLTplDe5alpYRxup6KK
R6UHm5R+Oc1A204xuNlMuLhNb5O5H0s9SZgNpQnghDc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 83        )
pgJ35xOcclLovVMxUHI+SdiCGKgrb9tJjxBjjQfHUnaPJjyERVYKmTqYQOdZrgow
y0bGGul9YalXNzDFnFem1oMkkqzOW/PB47OaKSjkJIyLj2ENKtNlWeZBC6clVz3C
`pragma protect end_protected
