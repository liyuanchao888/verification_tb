
`ifndef GUARD_SVT_AXI_IC_SLAVE_COMMON_SV
`define GUARD_SVT_AXI_IC_SLAVE_COMMON_SV

`define SVT_AXI_IC_MASTER_CHAN_DISABLE_CONDITION(interface_category) \
  ((cfg.axi_interface_type != svt_axi_port_configuration::AXI4) || \
      ((cfg.axi_interface_category != svt_axi_port_configuration::``interface_category) && \
      (cfg.axi_interface_type == svt_axi_port_configuration::AXI4))) 

/** @cond PRIVATE */
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_ic_slave_common extends
svt_axi_base_slave_common#(virtual `SVT_AXI_MASTER_IF.`SVT_AXI_IC_SLAVE_MODPORT,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_debug_modport);
`else
class svt_axi_ic_slave_common extends
svt_axi_base_slave_common#(virtual `SVT_AXI_MASTER_IF.`SVT_AXI_IC_SLAVE_MODPORT,
                       virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport
                       );
`endif
  
  typedef virtual svt_axi_master_if.svt_axi_master_async_modport AXI_MASTER_IF_ASYNC_MP;

  protected AXI_MASTER_IF_ASYNC_MP axi_master_async_mp;
  
  /** Snoop Transaction */
  `SVT_AXI_SLAVE_TRANSACTION_TYPE global_parity_xact;
 
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter, svt_axi_slave driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter, svt_axi_slave driver);
`else
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_axi_slave xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  // SNOOP PROCESSING RELATED METHODS 
  // ---------------------------------------------------------------------------
  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_ic_snoop_active(svt_axi_ic_snoop_transaction xact);

  /** Removes a snoop transaction from the queue */
  extern virtual task remove_snoop_xact_from_active(svt_axi_ic_snoop_transaction xact);

  /** Sends snoop address */
  extern virtual task send_snoop_addr(svt_axi_ic_snoop_transaction xact);

  /** Receives snoop data */
  extern virtual task receive_snoop_data(svt_axi_ic_snoop_transaction xact);

  /** Receives snoop response */
  extern virtual task receive_snoop_resp(svt_axi_ic_snoop_transaction xact);

  /** Gets the delay associated with snoop addr transfer */
  extern virtual function integer get_snoop_addr_delay(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals */
  extern virtual task drive_snoop_addr_chan_signals(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals without ACWAKEUP*/
  extern virtual task drive_snoop_addr_chan_signals_without_acwakeup(svt_axi_ic_snoop_transaction xact);

  /** Assign the snoop addr acwakeupc assertion cycle to transaction*/
  extern virtual task snoop_addr_wakeup_assertion(svt_axi_ic_snoop_transaction xact);

  /** Drives the snoop addr channel signals */
  extern virtual task toggle_acwakeup_signals_during_idle_snoop_channel( );

  /** Waits for the ACREADY signal */
  extern virtual task wait_for_acready(svt_axi_ic_snoop_transaction xact);

  /** Deasserts the snoop addr channel signals */
  extern virtual task deassert_snoop_addr_chan_signals(svt_axi_ic_snoop_transaction xact);

  /** Gets access to the snoop addr channel for a transaction */
  extern virtual task get_snoop_addr_chan_lock(svt_axi_ic_snoop_transaction xact);

  /** Assigns ownership of snoop addr channel to a transaction */
  extern virtual task release_snoop_addr_chan_lock(svt_axi_ic_snoop_transaction xact = null);

  /** Waits for the data phase of a snoop transaction */ 
  extern virtual task wait_for_cdvalid(svt_axi_ic_snoop_transaction xact);

  /** Waits for the cddata of a snoop transaction */ 
  extern virtual task wait_for_cddata(svt_axi_ic_snoop_transaction xact);

  /** Waits for the response phase of a snoop transaction */ 
  extern virtual task wait_for_crvalid(svt_axi_ic_snoop_transaction xact);

  /** Waits for the crresp of a snoop transaction */ 
  extern virtual task wait_for_crresp(svt_axi_ic_snoop_transaction xact);

  /** Drives CDREADY */
  extern virtual task drive_cdready(svt_axi_ic_snoop_transaction xact);

  /** Drives CRREADY */
  extern virtual task drive_crready(svt_axi_ic_snoop_transaction xact);

  /** Waits for rack assertion. Times out based on the rack timeout */
  extern virtual task wait_for_rack(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);
  
  /** Waits for wack assertion. Times out based on the wack timeout */
  extern virtual task wait_for_wack(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  extern virtual task process_snoop_resp_channel(ref integer crvalid_to_crready_delay,
                                         ref svt_axi_ic_snoop_transaction curr_snoop_resp_xact);

  extern virtual task process_snoop_data_channel(input svt_axi_ic_snoop_transaction curr_snoop_resp_xact,
                                         ref integer cdvalid_to_cdready_delay,
                                         ref svt_axi_ic_snoop_transaction curr_snoop_data_xact);

  /** Samles the RACK/WACK signals and associateds with transactions */
  extern virtual task sample_ack_signals();

  /** Drives snoop address channel debug port */
  extern virtual task drive_snoop_addr_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  /** Drives snoop data channel debug port */
  extern virtual task drive_snoop_data_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  /** Drives snoop response channel debug port */
  extern virtual task drive_snoop_resp_chan_debug_port(svt_axi_ic_snoop_transaction xact);

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function void check_snoop_to_same_cache_line(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function void check_resp_to_same_cache_line(svt_axi_ic_snoop_transaction xact, output bit is_resp_to_same_cache_line);

 /** When a snoop response is received, checks if a writeevict to same cacheline, or a transaction with AWUNIQUE asserted
   * is in progress
   */
  extern function void check_writeevict_awunique_during_snoop(svt_axi_snoop_transaction xact, output svt_axi_transaction xact_to_same_cache_line, 
                                                     output bit is_writeevict_during_snoop, output bit is_awunique_asserted_during_snoop);


  /** Initializes ACE signals */
  extern virtual task initialize_ace_signals();

  /** Processes ACE reset*/
  extern virtual task process_ace_reset();

  /** Drive default values for master signals during asynchronous reset **/
  extern virtual task default_signal_values_async_reset();

  /** Perform ACE related checks on read addr channel */
  extern virtual function void perform_read_addr_chan_ace_xact_checks(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  /** Performs reset checks on ACE signals */
  extern virtual function void perform_master_reset_ace_checks();

  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();
  
  // ---------------------------------------------------------------------------
  // EXCLUSIVE ACCESS RELATED METHODS 
  // ---------------------------------------------------------------------------

`ifdef SVT_AXI_SNOOP_FROM_SLAVE_ENABLE   
   /** It configures response for exclusive read transaction */
  extern virtual function void configure_exclusive_read_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, 
                                                                 input bit excl_read_error, bit is_overlapped_write=0 );
  
  /** It configures response for exclusive write transaction */
  extern virtual function void configure_exclusive_write_response(`SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, input bit excl_write_error, string kind="");  

  /** Returns the consolidated response for the specified address and control attributes  */
  extern virtual task get_slave_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);  
`endif // `ifdef SVT_AXI_SNOOP_FROM_SLAVE_ENABLE

endclass
/** @endcond */

`protected
\VTN54KP&Xd7OUMC(XPL-5+.C9?F9B4<??P[-)#/4</fg77e.OEF4)PeYcAL0GLN
/)/3]^]=;>PReL<XI@a?W57K@.<_?b44)G.4N6E>=HWT//EYE[e?.\6-aZ_AF.6_
Pa8;(-17g#MIU512?f,Z013&_E6+QI)>eBRJgU+=8:#6<#<cXOJA=N_^?F\M;HP3
88VX=>H;)UWBO,0]L926O#ZLbO\Z769c=1,OZE6&1?D-#@?IQ@I^DZ16=AQDVBWY
#B7MD<VLF\CP(M>=7XgWFCML(_@65>(R/SgQZbH\bOM@QJ]T57T?3IR-6BF^KX,&
EP6G:.Y>4Kge@:O&>JQb1K>9]6KRaSD6XL;Y;g8OOS]=@AC-2F8UAB51&?H^YaBa
eb)N:2RF[A3;27TP@<\5#KF_4AQ&(MVeB_I/0,E+IFE0);+M[[)-_[GUGF8G4R_B
(c3SLKb_[>9e)U5I.^K5cCA=OFKBW0+DMUO6:33V:UY)C4EFL)^+ZQRQX^EA1+DJ
_AIMb]+CEcUge,@8KPRHB2(&:ML92/cTN0HP,,C]1TG=6Rc0@bSX,8@]J#7DC,aP
B5?LSGIPI8VbU;#dPH3MXHI.+MaH;dPTM(-.5A8Le?Tg(E=X,KT0H/=FS6XJ&GP2
_U_W+SSfL/)SeY:,4^3T.]aTb<9LS;[SFN?0>VAV4G.?G&W&;c=Y8M7G8R&,V-<G
3=3(cDf&1&\UL>MH]JJ2IJ]e?X2/^#]TVUU8WfNd.;7=+M=..VGJ,T[:9daQ=0PR
60#+Z)DgM6^)Y:eGE0:NO3N+BfFRK;ZgFd)B\b496=<&3-9\gQU#[e;YS_AcUSBL
DG[G6^&58W(fMS@7H>Fb)GB]UC;<=E8;CFeM7U0(Wg>Ta-(1gEIE#G;/;Fb]9W74
+MfO)a[PP^H::38C1X_,,>)c01XFXfC:eXX>/:O+673IR7]<bbQQfMQcT.bFB,:G
7YIVHD<-\@@7a/Gd6f>fcQ-7QgD7@)S_^H3W;^Ra6?bKFG9PcN[05[K:7G^2AEQ1
Z79f^IHAM&NSGVIRFOQ#W#0WS>&JH@Y7W^MZ]S.X:W4IO@7/a=a&5,3bGcUdFZ3Q
F?\^P^V@;.I#:Y9+?LY1]6/J<eJM=W,II#&bUOII8_1[_-:.2,#/^(GX<OW]6K9?
]<8(IY?_,,GTSS#5?]=cH#He=9E75P8KIC&fXA+U9-U?F_S4>eRH[HC_L_NK\UQA
H_:XTK9ISW>gVL\-V&_<[]#a+L\\Yf?_C^Yg;YXgFeQ^cPbT/VfK]?O:20eK1X@b
J6=DHN-d7IEfU:,889edV:::JF__b-9=.OHF7[7d((+)6b0:J6[_.&78e]XA,F-I
/68<OXGZ+U:ORN.KK\dQC.TgC7;aH:bLfCT@5C-D?d5A0R,&:T=@_c\,:(+==3Z(
D:6Kf\XUBJ,9;-WMZ:W-B#\J\9[(TTR\aWRL;4eWLSVFe?d0E5SQNKeNFGJW.:KH
<M#WY\L&#P9PI85f-:5LAGX_b<[&L9U)(C70M<:&+]^.RJ,KU<Hbg)e-5GbPUMKK
=WEa1QRB),(6EQeP1\S@W7P#e[A[1(FZC)K)3.TYM3\M/4HTJ8#,/5+a0M+Ga0c7
KF-C8V2U];],AR[d^>XUPPXcUUX;B3V[#?KHL)NBdLcBd3?O23QF52[gZaA-.GYP
N7-@ZbFY>?/3f9b<6XMZ9LLB56V80Oa0IM_1ZSV.dg_.R_-SD;\SOYKK#c^c?U(_
?8QL5/V2@3Y_7cS.09)H_#FWEL?40MD8HE(<C>MB<9O.A$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
#,(A/Y9)TS,YR1MPC8aA>c<-W8M(XP.P)M)()1HL1W\dXDG-#QYM7(NZH3^TYKYg
K2d4.6dFAS(e<+8@WR]W;OBf5[H5S<c1-KLaL>+I\H87\AAFL1;EKX9bD=0FTZDC
O+JX3#79bW.a&=71gg7U&+Z#S12L&HP2-ONg/5]gWDf&)#d_HTaUC5PF=W7<&bOA
bG5Te,6CL3+HM>66Q:76IO;1CLS75)(75J_f.6._EM&NA-WV7FbHH\[L6;96IG(,
^][R3=EC7caU4>\8=(F/[83[cCcQ.4?E=b1:?\P,/KfGWLP7VGAGG_):4fgZ3<e?
?LY]TR@#>9NdY:M<Va7AO&<<E12&C([eV4B/@5M0.Pg=E/H\5@A+?LY@IWHS_3L<
bDXbaQG#I2+23IUAOOHWJ\B:RedRJf_.ARV96G5Z9TFa&1D2CJ[QUB(Rd-T5,N,d
DTO=IS_J,YN7FGE^[bAf3,CYQ8_=-^U2eGg5>&6=(AOEF+eX;b.UU@F&QR@U9-SF
OA;IP;H/.62&P;7G9:=?]fZg<FI_bE]+6K(D:MfT?+//CF-VV)OZ^>=O//=;e31A
0Ce?1);:6a[^_(<-Z_PfL.47LK-4cg9(c?TGc[N:-^7Z658IA4dCg6+:-@KDefTf
+cGL2_[K^)H:O>QN/VQM7H9C1+SJE<Iab24-9<[>Z92GOWAZ8.@OP&AU18<bdI&b
:+17&#CbOCaQ/J,H1UOBM1^^-[,FdEHOD?ZM>f9Pa<4/0,b,07>3QGa,Ke,g[>,L
Z@gW7d:)<.bTZL<Tc0c:D\)IA4;?EO)7JZ?^+b)4_]EA37V[)#YD0LAQ-\IUTgB.
R@<^(;g2#Ef,^7V8QBdN=_BTA,3ZVCCbJT98(g;4PM\8Y;OS_UQMB<N,5bd/:3MB
N0^TIH1+&?39GB0U(&,\>3^>\eI>fS>JTd8(0<d-R66\EbXV[O-U\feD&O=O844E
EX;I,,KXR7R^^QKO;AHRc95<&(VH@[P,S,2R9&)E3C#Z39d;,_#Xb+-V?&U-B:BZ
HJTI#KSY+g,3KKNEWWD4d,FN20+8P]b/>0H1NV-dH/dL?YX.27/A:e;0444NZQSJ
/H:GK4bV4cJC_MJ3AM)=C\fBK;1HOC[G=@+LF]L(DcIFK.H8T+eE+EEB7-:@ES/g
85)Z?b[U(71MKT2WY?&F6HU4KC;QWZK[\g4<#C(a5T;&R1^/77/bP;DEM?5,+(:D
g5DWgg4b.71[_]_+GD_9:6fcfG<fXKUM0WKI-g.AXI2.EEWMGL70)aODF>U8OE3V
&@@FDA;47+7_KYa:aW+[T1;4^?)M\ZE(F3I[-F=LIM7U2D<VNRTY&dV3S8g\G.Z2
BHQC0I5R<P6Fg:/_U[Q).02VLBbNKF4JRZg(b-_^GOd?S-EM.7c;\EJ2M(YJ>[/U
GL5CgVHLJ]_Kc2KXKH7d09@X)b-N?>&[LU8XY5Afa)<gYYB8.V979UV]EADJ1WdI
^J2G&/<(f:W_?GFZ:=08^LbG54)-4fMfV(eO3.OMB,),ZbLc?UaWS_<QA#;&,BBY
<28a3NQ+#]FbNaI&:fG,L\7P&]5:42<YH(=;]G[0V9)FYa^3gCS((.Bd\1QIO(=:
74O.]6P1UD7901I,U58[e9I:6@)>gf-41V;MWDBEUDY=-H>#gd#UU2ABg)+FHI=\
/H?<WOaW1(&c71[M&\7GS=b1A+/)Z?6(T2dYeBZddP:UPbNOgKZO04-e@9;.>P[&
LMH8/8cJ[ZQEbIV;40@]50V1+&-2dOWOT3a\[=6?S?C)Mg\^E/3X>>9#9PYN@KJH
A5&OOJ5D5.1aSO@13E84RH]L1299:F_bG>2#WY=_KQ(;,cMfBBe1W?GU][PcI-Wb
92.d9@@I<CTEZc9<g1b+d9=:DHebCCV>Tg0\982Bc=T@H8PJ#[RLH7(=OF5)cFEZ
a3UbXHH+(eb5/4Kb:/d21@G[0F@D#XP=1.Rg?GPR8C:I.L).]77Wf6(311cf?g5;
5aP@BR62+)PPGcKc4(&@KT\\E7^JTNJA?KPB/P>e9F@a+9D)BIO&+^Wc/<_a^_3a
LK5M.LH@#c1KZf-.ZgPdB@VH+CUeEE@M(1_P:aRJ6)0^[C\fC]TGU;_-JN:afa,=
3P,Q-KL#2U2>XLb60B(N(8)?,)=^/:52K;Y4eVH)a7)B&?G)G4_cM2?BJNf12>S1
B_8^82\3T.<\8<<b6-A7_).:;ba=JLESWfQLLfPd=&G>dV34=IMVZ6[\e9Y3>U36
X/FNS5G4(429dGWRQFE#2\eJcAQZPF;cQfYWI<L#NeVLPB(GcBNC.GTC>,0>1g-2
NIbU]aO^SR+:J[@.8aW4;+@IeT/KNRX<Z+L\(5R-Ob\EN\FN]_[5E;R9Ta3M;(C[
aFaQC^Td?a3H9+Z:TB5\fB/ERV5F1\7U<5NL^1];WQ0=f(0<S2A32(=BTY.@bLf7
&(.N?FH#>/3TOO)XQ],-WZ<<<)\KXK3ZUb^c8BgM]gB[U12S&Qf]Q#L6<-PcFDEU
a2KM;b,1b,^NLDIea\@=_7+&eSSP]8R<M865<c[.&EcK]H75Y0be9-TfLI^)eT_.
M(XK(Ia4];^[,2:<gTg):1;-MGWSTeJC/EKD2,:B81g\OCFeC-;HE<#OcdY#CNe(
K2\eZ65:XaWU#8\Ld9^6HGZKHM]bRQUOgdfb27?+O:T,U?DFD>b68e#E/M(g<S(a
<fSF@7],F25Q=^>CNF6g2+g]D1.YHNbF_4\@__AMB_E>MPd[I(\AGHEbRB5^P8I;
DQLA+Q/Q8KgX5OOH((W7GWK,Y3.B?G[-X:=HRYQW^47Sc<=2CY)b(#fL#=L:_U@V
d9+]7ZEN^6\Z)N+<N5fKJ:UB#^,T8Ge[X<\>RZfK?,:E(MRD_)<a-.40?)NVd^fR
NPMOa1;6,;25E&[C#GeAGJ0]NPa(=>86FGH<dWWd<D6(8f6\VRCg75O2#g_a@.UP
NAg(+FA,P@F1/GfFZ//aD9:5\D7U@H:TYAfV)1Qg@#SbdV-2.g^<DGEJ5\De@_]c
cb9@8gcdN5AU);OAY[>bWTAJC1YgH+G:I_cP[:3I9C@[OH&eC;dEI3X&O&E<0+-(
(=0G,BadRL@=PMI<7M+1U[:/Ze2J><YG#SUZb@7],4UNR\N<9E@L/DCD6?U<#gTN
RFa2VZ6L]>)CE0+POWdEE.\9.Zd=R>POQKKWW5[f_c,/d\4d,_?XMC4[/-,cBT=b
@+)FV:U>)C)DBT.R/E)A_0f1Q=9J)]L7RMTY<M6VVYgCBM+fL??SD_P-G7181@4)
<Se<.?Q\CIY7EJ1a49W[<O/,C([eJ4AI5+E7O0E<(?c0BLF>;P@Pb.W&9&ZSFQ/(
Jaa>D,g0d<)].T9Fd5VQI1g>b==(6f4BJ3O\E?(93[Mf6f#Fc<+OZ(1<:Z?GGWK9
>S49f^\\F5F,V/b3J5\G_F8;XFObfDRTSS(@0TZ;S/gV5a.Od?S[?IM.Y<WULJfI
6BY\6Y)g>)FI2A]&XA-RY3@P5OO(Z>D9aX386UM08aC5f;XQ&<9V@21BGYI;(?R1
&)B0b8W6gARZB0BAI+gWK4#Q[;c]C/@7-4b=B]^0#DF8F03<IY1_5D\Q<I\_.a]:
D\FB:-&b0\Id:b_3YC^T<73?,-M,f\5OKOCe=9Z[GH7LGH=VZNbU]]<aa,#<RCN]
;TOB.A.PD<8;G(:WUK2#7GadcP7-OBQ/^1R66:+E-#8MHY9GRPc6EfCW74KPK74,
CJP7=:+61N]]c7gd]=8DT7([>e.;gW=U0X2.f4EW\+:U?PC8S=OcA1\GSc>dcAgE
)/+O1=H)2gEO[fR(N():G_:S61&HT/8WB^ba?O5.c66)C/;46[)Q&(^PACOL2(fG
QNT7(?d)EIBMf&1FCXSG-Y7@^g+XbD]>295,2VL>:Hg-Za#)OMLb,#YQ[?Tf377=
CNLdR54V-<=8.Xa0DT1,dRdS?8P-gC;QA+]OQTe2R..d[ZD2]K<EFX,Z/8Jf:.RY
5TBeO9cb/;.Q8ZL-&JV3&<7e#4T31X>G7T1Z+WUH/e5-R66e--?R=95I+E5]#N\d
\_8J?VDf,O;&F4CJ[@fKQ6X6JXaUKY]7\(<4&B80Mb5/V6^1^;AF:,49R<NRfWFS
QK>DFT@JS_4WJ?CNYbbK&Y;))Z_/<.N&7f;bA@b\bN?[TV=X<[SF&Y_65@-YaWS0
YSVHN6?WC?FeO\@::T)+YL\-eJ&)?/eE\Xg?R[?798Og[24B@+^]OM7b+[A]OBI:
E?[+KM7;V5I48PZD]4,a8QC],T^24,:.NX]Z3.U3Y8.d9^f=L4^;Jg(7S+79&4DD
V\>IJJaZ:MDV=MDTV2aTDB-U;3UZ@/)Z0gV7CZ,O-E.BbZ,M3-E/dcf9+3a&:ac0
7bdCeQbQ@UV7G3H(XGQM\&]#.YF3IS_=KW&VM?#^c_7Y61H/f2Z/1OIE5\b,7I0H
W<E&?O7aP8-4?f4AA#&+G_1^C<e5M:04eSQ8fK0)&>GPO/@X;7CE8#&8BY4a6@^S
A\UG3&cdBGT)4WK)<C?#F?-6LFG19K_M):P+19#UWRML_?J8LRT]HSLC@?^>D9L#
3J)/DYOdM4SM/GS6_&Zf.-:/]?E+B56FNg/@[+RA)](c1_PVL0NK.eV._1L,L#ag
0a2a61V9/R^+d\75LR(64M:M2NB46;>+aEOQ:,3DFB1AT;d4FK?7<I1g-E&Cag-0
bU^Z9(#R,YVQH^\J2D([cFDS2c@aOZY:V)MN7Q\&EZJ=5JQ#B;&@gHR?VEf6bYX=
g06\S6&BQJ8D1:X#LNYD=3)_=6#X==0PP(eONaR/52?VNgT/X8+-0(,R8I3\G<3\
1N6OLXJ]f7PG@R.TK1Z@?FD_I>[#fE&]RO0NRF\229DN?8aI#;DNRGV&H1X\[MGT
<,<63DG#WAPC>Z_c5>-108INegQdGX9G-[W-fB:VC_\CUFDTT-^WdS)+<,4&g_\O
6?DC_SaOISP(C&/.^b>:PO=#65be0WR5C^I&7^KcJKZI6R/#eG69GA.Paa_O_YPa
O+P)<bJgf?&&6(<YaGT&Y>JS?ZIM#UH7+UH\(9337P<IPbI3]58=YR[aJ(eg8PV2
W<>W>PQ[\I&fO,VcL[dWU;MT]\I4^/[#NaF3E67NJa&-a^I1e]B[:R&M+/L.aWX]
FDK&[[HV<N4S8B=9Y;/Z,BV.2\0[TJ<Nf[cG=KE8Be#6DW90OKA9;CIB<BP1#V-(
NFD7S@bf2\#V[<2cPUZ66&KIVGNTDE>\cWcV2_/P>EY0[RNN9M5IH.b0bG(LD+4@
J_dH,C##KbD>aX.B.#KI)Xb(dH..&(S5EQB;O2A54A4II3_b==PD,8KS_TWOS01&
G=.NT@Hg9/;TOJgB\/_Q#PVMX)[\YIKTdA>LQLZ&:@6<2JP2:/N>&>fcW49C4O3F
O(9EVK8bg9Sa2,VHW7]+R_](S25=]?-SK=<8U^VI:#)SRf.a?]I+JPND1/8eQRHI
7IgW1aF=FE4K#>_6eTf:FG@E_2/VSd\L@SGP)gX6d)9)SZ;_(81?:d]T5FD\:;]8
)Q;aYDSXZ-@fe?QSNBL8&]@R0@EC/]f#0c7aM@PgD_-[0:NI\DF#]SQ+J+[R(I8b
e/NK)8cTdOJe_R0;K1O>4?B>9TY3=Cc=HQ#^Y&e@LH\bN_g&QQW6Jb_g;e3-&EU1
,V?f1B@:CD-<27DAU,C6.)X4>GIf.I9>fYB^5];g+)AT@dU=8C5<EdY,^NNZ<LU.
,EW1H?4(@<K/2f-3/#4MXRWX.[#9BK66?5B[X/1&I6P0CUK.bS]#WWdf-/,aXI1c
g@eA61N>65EcD^LZQKWbLD3aOO5Z2=-PLILO7A1@_@7AaC<Rb#Na7)GDGF1C+)J7
5d<Qe<QY;Mf;&1_B?W02_JX,BD1Ba?@CZ18TQgD]0PQQH(55Z.5.MTYD-@X-FFIY
B@^#Le;:=[IYA\Mb#9LNENIIgc42G;[##VWI;,=ZL;Pa=_NT7dfPF[N;dI_NZ,Oa
,<.?U]KC\3@3[3D6<C5Y/4<](&+FBR^S+/1X4.2c\M]1dD7>^?2,+A]^fEE-;(KJ
1CeX>X8(X@(cI95=a;I0FcL(II>)[(:1/:=M>E+F273QH,Eg]H]NON_gS4I&aMFL
45#0[L1@4<]+a<AV4OU0HZ#V=7A.0L9MNBL\b2&8)U\W-&<D0J&Q0KIZ+#Yc#30F
fC)V)\eMCZY]92;g/HNc]/g7U0;X50<8P#e__,O?X#Bg/WNEK0-OC#A__VVXDHCR
CXKU9EEdS4Q@GY9=,(G_]Q#S2+6>R8cHQ2[cd,fGA\X\Qff:=@P<aG9)JU\Ia6^.
T<L/TU4=.]?A:_fNd]>12)@4.NRN8d)+#?<E[)DbfT2LW/DAb(?F,Q51?d-.ASIO
X=?P---AV5TJF8<<UR3(].c_4_PH8..?2_4@a[[4(4dK0<TI;3^LaFZ=:&/;/9?@
_PS_C00/M]]IZ7C4eH_WaBg7dE@84VAUDXfT5^,<.4;#(3Z#V3L3d/_@X>&J+/@^
KWba3116:L).8E-3D8\<WOSMKAW9Y+K</>9W==XY6>5<Rg76e>F&UL[^ScHS8HO>
J2V&<8)6f]b:VKf0(46dXP>VM4>R?G1.+_J;<P@=B,]\Y+=W)^CIa8Bb^I+Fe:7=
+;PTL+H8LI,0d:=JUP.ZG?H12Q)S),J5+g60@cB4_MOeT.64CgLT+T>W2;G_+V_T
/a4B-ZWU0f]U@IB@A1X8_0EJ8Q)P/d#;]e-#)1FdIZWIBNLS:HaCP^E-:A90WXa2
f+13NXFBaR=:Fd,bE3@,MGMT=;]XC4a;V<:CF<6?JQ&b?D^3OE7T0+W[V0f7H5>2
f_UYgdeFO:)OUG#?>_=?[0@NVV20IV8ADJ;JXJ)T#UH,9?S6&]NY:+;?Pd,Ie#+]
cMX;3?4OUG+^dOJ>>K[VI;(Q3?KL<a,OS:c)02.3ggSH.F8KaLF:5K_=]SVc2:=a
0Y6-CLNaLH.]2L1EFN]_#?edF@3>N[VHa\SGR41=9eO0ZL<]R;OB^,]#_S#5-7^+
,4K^.b74?K<<,XIbF>#7CM_>Y4CPFO-]D8KcA3EM(c28YgD@2d.I+S/HLI=)&E.+
-QaNPY?8+FT2^1e(J;F<\b4Bc71R^70I4cBbP#/dX/0[5gdFD6+_,^d\-9]/6CI(
8d<&3?EFI3U?E+1WPcE8M1afG:Z^N7XP969L[C5.6RB^KPVa=4184?gPT;F8COGU
9J&J7b,I5_VKKaOM(MVd58GBd3;)I)NaM<(QL?N\;Q4:7;[JJ2L9UN\cPA_JCRaM
+P1d0J7]C?b2ZRA.,g=b,3KAULHd1<E85J.;GPY&=3_&2O-9#OdCU[_PC1<6d_TT
1O<7a;>e43LHN(2)gdd[KWIIBa+GVZ=Z>DLgQPCF]&HSD[IJ@8B:CH8\UA2&UDDY
&[=ca2_Jg[09.20:?\H=g1-;YTfJ>J@cC+_3;JJ&3)2eK37Zd3Q]5R8,gb+B>&;Y
TYQ;Hg.A7@Y#9.Da1^EWKaXbV#D0cYORQc@L309:gTK7S6KQDeVKF,.GF,T2OQIc
-HHdB6EcgRLebc]>\f^]Y5OSa]:;7J-KAU6,O4,;8DYY(#OOG8(XCbSMb=@N<gIU
aJF][]RD\16d2&35d<P+fIQ-OR2A3L8;0U^Ae^9T,0-E#P_JaHcIV^@+gfZ2C((T
ROBB(BU,2C&,L][J\9/RNHHP4gaUQdUaV-3+[e06Cf\D.TJ;Z=,8UGb=TUD5;aX9
@FI:WK?;f1Ag(Q/R_3=U,;>NTCLb>3&S&;)\)7(JH-OKA^OdR4HM4DI;+cb[[:bS
c^VAB#;]<DeZ1B.O,C[ZC=?d1^49.aHYU&gZY=Ef:AVc+T.&2HJ(&&0]ZTY?2b/]
@,Cb>+5e0;XRBLA-H?EZKFH8A7T1D9d\Q//:;7&OVZ]MVG=U2HMX=&Gb@KVGc6@N
[8A2D#]Md9Q0&dN,FA#8[HN(N8+K(TRSV;Wc@A9\@CcdU[OJ#d4GgEc<fH_6F=ga
,Na+-#G5B\CF=;8OG?,=,-(;H[e+WHLff<Q._/b?/S/Uag_g_&P-1-XG<FOJ&8<g
ZdeNF:?-Z53Gf.+=50@UFeG586OCJEWaT5TQ?;Z0FI<H=V3+P801;;B@\RR/=ffT
N^,B<?9>F(-5c&P)@&QJAe6WW37LRN<Sb-;@A0YB>Fa1A[aX+)MeI&AZMV8CQ+[e
\25VLIg05aA>3(E7,Ge640]SVcH+a>,ZH)G..BT<),f=ZV<Z?QXL>L+R4EY\H.UZ
:bbF[-W21L(>b9@T=-.3TD=6TS5>MV:MZ#&5B7:a7\G(TN/1bS)O[C,-E&GIOEg7
H2PgI8fQT4c=aCK?QD/G@B21N:fP4)]6N/W<A[81K<b&NXfN9=+RGIeJAN,+>G3T
J]<(BG21AN0OSe=+.D/+EadP0(Ia7-IO(1W#BTg#RN35&.GcUAM/C)X;W9IfOVZ:
9G[557(]W/HO+)I\WcPg]IbEEE2PF2Qc<c^0+WAWKYa4GW\W9EBgSVRcfA7O5<\Z
4gQ>>_D#VWQ8N7N7HE6b0P0SQ)\QQ?/]1D=7T4),c=Ba):_FXL?RUF:@XbIBe5)T
1Jb@W7&\Qa/V:SB/+YdP+WMZ944BOHCE3B?#V.J<^Z+\4RR^CF;SN+bDc6GV[R)O
H[Q,W8N0_TD#SUJ?&_.T2@H=F0;ZAU@_8<eUKLZ<IeS_X<\?gZ,E?=)BXKVWa5dd
?8+WY][?1U:>+=)^CD0:C\,<XadLNBN#RQ5[H<NV(dF/JNMR:aH<;J]KKEES1),c
^-J]1UQf+:eIDWJ/E(BGHL[JBW>USN\7MHV:?BJ.OON07+U/K=M)Z#f4Ea^5Ua]7
:Y<ag02e0H:;C+-X=5^EVLEI&\(6EGa+cXfTK/_>)N#@W-CRJ<:HQgDEb@@2\55V
PVCB>aRa44IH1]bdU5-PK/-A9^W]V5I58.7(UD<I+71SB(+P,Bf&H1?f7/7ASP7>
bd-/g50#cLO88_JJ1YdgKFGYJf]d2912c=B8RNdY(V&,QYeJ]GGd-V,MQcf3>Xd=
#^+F,N,L;,8\9NODg=_eRX?\a+50P#=+\K6Y&+W]L#+>@=OLFeC./YE&a@f:4-LQ
&aCP6W#231\>V.=(B]BMXCd7#FIf,YKeHI>IZ>7;;9UMG7D?9YH@0UZS1g;TZcW+
O[;eVC9<\[[OX0VY&03bgFa]KU4-OfZ3IW.Va?BEa+7Wf/\F_;GfMF@M9GDFVL2/
?D/.XgT)/TE+5SLAC.S)6P:)Eg19)_L0Yd?bQGcPFD^d6SL?BAJHC]g[N<NTFPV,
O\PYOV\93<HL]?<3LRKf.)N,4CN^eW0NWM@B1QV;,WZ(D.UG[S[@Nb266I(+XK#US$
`endprotected


          `protected
GUFOdeSWcF9RT8=3b[+7]4U>@\H[b(+@SZ56=EYg<D0UX02_NWUH.)H1NF<33UG#
-;:+AMM/Y^.3,VO>U,V=eZ;C81ID,RW=],Z3Z1a>H+)LTTDSc+P(NAH1I$
`endprotected

          //vcs_lic_vip_protect
            `protected
=I/Y;QIPD/HP.DI@QBdYEAdZ9(O&Z[cIedA]J//;P(,5L@#)JS.=)(NDZYg@BK@<
FMKY#KF@a5g-1#;SY@5cQR@=g>8Ub,5#A.g:KX[F1DbcB)1<:LA^\BfV)#[)QUYZ
(LgV8f6=e97N_N:afL,R8F.N+Id&Z_3gDM?)YP(/#XbV7a/WAF#EFW_d\FKQTKLQ
V93AZ/WMBPI8/#;6_8X2^3NV]4EEd]DeB&^@PWS=5XX?CRa^M@H7g1\eFPc)d@-9
T(QKX5HUS&=4ML4E?0Z/&#U[R>M7?[G-9dU:,BHA-&a8<6F0gVd1;DYMJ7EH-WWN
L(aF3FXN;^/W2<^TNXIO7LI=75D>;>0JdS^/.@QfF)2A+;D^YDR1d-g@0(;U50@@
T9b\83MZD>K#0aS#GEcSD-[,<gMHO1T4F/5F(75YW1MXJXW<@P)a_.68FL9GE_75
9/#^\aIaFL&QS_S?Y]9;O_#32PD6,:#EOT\7>>ZN.(PW@fMTU/Je&.FTgR2>(U;a
M?L0AKR(D1NJ4GLPTJXB60.9T-H>CXZ1JNDdEJ.3(NT,:R)J#9^gP[]W5MIIBNC_
fcKAUHE(.?]#.JF@,M>(A<LNV0(6#>;IADI^8F6O)4.K#f07<@<R8?#90HR^IF_2
K0YABEa:1<CKN\V3CNSP032Y/U4e^Ad9C23?U,bPg>&ZM1A0[\XL@8S<O?Z(LTR]
b0-[A&U=gT_^4cIg;E]dCAF?\@Z=AL5K58\B7+;1MfgDF?9a)Uba5.VRbBbFdJ1E
RQ2,Q?Z,V[RI?.M=0>A&BZGSS:MQ9F\>00a<BH\1E(JO;1J7QQ8LE-=NB,[?Q6^?
M0I&[(C7KA3M74?(QC7baAW&;ZT1,2PB,18\+\HZW3I8ADVP9(8GYK>K&ef:bQ4R
A4c>DU<aJf&,cb6)YcQSdN+K@9SUNSRR0KJ:06aZ;L,LTO>^+^G-Z(EL2I-d68R^
MKRN92;Kd+F6VcIS+IDX(]ZM:a=AE8bc/1U^)&[W.,QT2AMDLG8@]TBe9N9?EdP;
SJ(#8RZ5]1SR-0+IU-2B7=+EL,3c[YDfU#0VY&4D,e2.+Z/c,.K(W4F_UU\c4+fV
DM7OTRJ:XOc3?M5.156H;-D2H>37D72\86ED-W#2D6@=2A@aGY.8+V(EXbEE<4F>
a+?MSH@SJ3\g0M\@R2>7AYWeGM]N[H62-VUV5I2OPd<B/6[CGFgH_QX8J@Z6BGR_
M=cX]f:+=X#8T(,F2M4ccD#^?<_.Z@[[1Nb8@H1VAV7F6-Q1Y/YVM&KNTB6E>3C^
=ITRH;FNGT^4CL)([+OJAV?ZNa9M@M.W^@5&WSD_#Ba(ZeQP-cg0:QJ-[V7RH8]c
8E;/Vea#6YUTC,Z7HJ)P-50+A/(NF0#O]M#:\^2T=4a3K(a\HL=07V-4=V6\[DRB
FbF<5WS]U:75a/EQ<ES627^49S>NQ..R\g/YW(W)B?<_aUGUXQdM67NEZ&4.)RPT
VQKKSX-ReY6Ad74;1TXE0[)-V?b>(.R&N2<DKUA9[;ZZUf:KNL#e56Lea^EdY)RK
[aCff0+X>Yc(9-+DF<[P/T.gG7+V.PK[,/cL-5?&?9MZG$
`endprotected
             

          `protected
-;c+8=U:Q#46OS7;/g6DdKMAbC?K=>Y06YI/\1-G8ESg&.3c#,52+)8>4V6LR1Y1
W3g)a48g)I^Z&)@K#X3FCX.+ef4aVLc(>$
`endprotected

          //vcs_lic_vip_protect
            `protected
G7F9]/\aaQ4Z.;B^KX_55O6ceOBHCW\Wf,Ie=PSWYX;-e<If;J[/-(V/;.GeW;-4
S^_=Zad>&B<gHBA@GY0O;KD1WDUUS(YM9M\O71\/DHZ4\</]/MH/>:&NS<9dHQ6V
Na>XG:ZK4C;9,P3&b?+LDc5^6@3@P4FC=5-XgSZWSRA0d8cDO;/A0ZEg\K-JD>@E
QNe1CCG2O\;)2HMRS3G7EHC\+F@#bS-)_5_a.#7gZa+6D)[OB+R)L+X4>#YF9-A,
@U[2:/UQSNF\1S:2]TKRcZEL7G4;/bE9&SG->M?1,\?CRD;@Z@-D44W,/]WM8.Ae
X8)G.2C_Y-#>a\+^JV,.N0.aSRd-fE]0GSZdN+Y2\-#ObML<)N.W.E6</fK_=dP7
VTEJ(554b05C3bA9bJ[D?J]3.TJ=:AYO?IJ10dU\E4f\IE_g?4\:ZcI6/L>7L6NM
^Z][;U:CUH?TLgN]:MPM5NJYEPG)]8237S7,1<L>OLX(c0EE<X=e&BaPD-6H]H5/
aId5KCeJ-f^46TIFc4egGS^.ON/PO(SRaQTaFcHD)bBJD8T03_NJJ#/R?XXI8a6>
F?7_0#U1MB-U/5d56Fa^TL<J,cPY8<[g6X#\3=^BOdTAdRZOcb_NHX_eQgTFT8FS
HQBTg_dC+K_@#^V+W+X#^.0,Z62)5+<C^.RK1FJN4RIOROfANP.05)/M<;fF<IYY
C:eV1Q0a)9ZIGZ)>JcIZ1Vb3K?>ZcUO0cPcbL:#R.Bc&1U:/PB-;#R<_ggI>K9=1
I#.5R<N+Z[I?US;YT2),/:,Xf12P693J#d2G=137abB82,cFZ(6M8e:[/Ef4Z(f1
/=e)X0+.&_/:NFI148&;f(.6YBC_(Dc^[c]RN#.TPT&D#aN?UX&XWEaUe]e9HPE2
5YFHD)&]_;0(CEd6J#S7B,R)Q.d,eAIPX##\PW^QPY3D18R8X1ZWD&>EU5_[-6@N
R(F5W7XgC-]g\1E<&O?gSR_.Je6CMV]AQ^.J=_eHAD32(WS::PeJCZ^7dAU?Sd_W
>6T25IM3><313TZU7_f-fH;Zade@9Ig^fePVZV9.a3]\<9f^&)c#F3X+Fb/c1DO:
Y,JK78\#SZOfP.gCOC=Q;DB_Kga0[_3=[>.(JcW5RfIOaWU.4T1bOReW7NGG;#P?
#NA0Q9S8@6,L.=&ME=96U&(R[J#BeG?_C^)W;5/24XL)&V#T-WHb?O6-B\8JNZ?F
8-RT)Z\YL.1cG_NXNVDINb@aX]-d-L\UK/<1gBe?/O;;Z(cgL+-AKgQ[QNf:5I+A
WCWE6280;:BIXf]11/=1f#[=HB>A0g-1DF+APMYfc/<6F&CGTTXW//C^ZDaRc]B7
]&&caXD+@5[^N#W<)a^_.^bPDgIOQ1N5NVYA0>D^M5#AWc:Y&+1d_;Y):A=,1cg_
3I>JO6HTF@@ATWV].K^W.c#/>Q?We(=IE0XCSUE+X4=2a_:G#H>7_GB>\[7bZ9AS
AWF/CKJ@-@+fEB[LTG41][>&U&BUH+?PZ,@<JD^aJ\4)T\Pb\0[g+Rf:#VC:F+Ld
6-b7^[;G=7b_EXe(-SZd\#CJJaZ=QKgHE:ZF8_XPO?3-gHT=]1?0\cFMO#DW3J#_
e^ILQB8OGg64SQB606?-ZcB:HOVS^3OKFIH9JcNL:A)AMHE#e,IW.,0F1,9=Vd,(
;HfE#LF\O9PDYE=Oa>IYaCZR,JQD6c]O><R6cO4K,S;(K[RWI>-gLTJ.B\A3J\D&
:+,E7Z_C68/?2B6QS)CTYDTUN^O-;LK?.;,7<b@70SZ_g/3)DE1a?XZUCW?&,8f0
TZE&B8=<\N=#,Nfg0UDKCL6E,N9[M8e,WC_7B_I<<A/RPbC[M7-I86&O=E;<><XG
2/G<-+/^I]e?LR@TBL@b41Q7AfQ6OB.?1?>39g;WB_4a;PPIBIL_@4W2F^VM1;J3
=I1ZMI+_N+1SObUVBK:)\ebg=_S5M\e,ULW.7/[G[=C@_)NgY&K/IVb1;C\YXa&S
L,T9[_a=@ZQ&<_^9._CGMY9JO4HC,Of;_S,08OKJ=d])4S9P5(,;XgL37ALO[MdC
O]a8K#</-Ac.O:C;a7RgEDS<=<[Z[cWc0ZNLR3\,GaK9HE+.dNI+U0W8O=/(;?gC
,JK<0CU(dT]PdI7Q&-?]ZV=g28gI[D/261Z>HD^VJF,MYUE7UXfcZ@AcT)NZX.+c
acR4H\@VGdN7T=&eWMbI#]/<&BcN4<5G,Nc427g^#T+&,>M0Me2D_B-45]egK@>8
OX[aK_SfJLX#FB4a1F^0ZgRd3>6=H(6&ab0G/PUeEZ]]KO<]BTR?N)/N/@N@=/XV
7CW];/1F5SUacXE-+7-&Q\=QWDa40E0NSDK)&;gA-H^F69W]</N60(gRCb[4)-5T
H+_2_bHFOK_JddHa:])EEAT;&@M?LP^XH1+.JJD=&f=.P8VTO-J&>C\a43QgZO^5
A+II(MH@g4Qf1E.gV10P/&?@SbYOIH,B>I&1fHSV\Zg7U410G_H[cCb8_9O,RSRI
I\ONM509D;eY)((,I<[0<?(b;\d&eJU>:4\&Z;>S.4XM,dd+@A3cZ=(^WQAb99;9
PK0@gcOa\-L=#&;46:cd:8V4_M#a7(eT908)ITSP8V]Wa_PD&WTX_bGVOFZdDf19
V[K:ALG7Pa\+8H=]>#PUN>]aS6()JX)V.I)D&=E2+2#&>(EI<0^E/b<U^[IZ?HCb
20(VA3LMg)(=.LF\(<],_.B:SgWX;;c(MP(N_X=+L]UQU3<_DfUO^M-H1YR>[+^)
IW0d#R[\Va#39I5&)]16VUTg0Ma[F-C0V8_cc-?7E\OWF]Y@D+K3<A(8=:(Pc&V^
OOG/HD.(D.#USbJ?F4#c72AILO25C83I5_Md;5-<SVBNcK(UID6(=XB081<9Z)Cd
ZR@AM.8+[cVVS2LZ9U9YG.0,=eG,NW>3Ka4/J1.S>c&:-79,:Y46B=T=B#g-+I9@
;+X/OU+)F@AC]DP)M]J8dH0@YT;6WZP4Q<aPP^c8LK#DJ,)Nc6dJS)Hd+U@20^9C
97IS5@AB)6^J99QI:_ZS/MeV34gR^@G@+<(READE3SO8V14AJgTg.U1L?P#]7bH,
RM&1RUG+?RNKWb=d6KN3PAVJXbN&>#)OUE6dR)(O43[.KQbLXI[=e@;/M2f=B6]P
8&_A[dZRTVAG0;YNd>]Y37^+ad7,:6IE8)aKQJGg_LI+,S^AL,>eHD)fG8JPY&ge
X.Oe?>(1FU:ff:Z=R1@8e1G0BTE3OaN#eRdU;/GXBVUK;8@^<35B(44=(BF;O>6@
W7XS^0P_RNIWO>==CaK/OfAdVBG;L29;bT[);4ZMWCSUGR&_3;Jb?/:-QKV&7B#8
Nb,.4(5R8a8CA3)4KX9^JeeIY2Q>I[.D@LH-Z=R8<MXT&f]6T/cd=757g#2c<S&1
AD9e[=:f9W>FNDJP(#&PO\,DYga2b?:1cagLSO\K_K>GT=&8+:K,HJROa7bZDXZA
;U0IbM@CTD?L1-B]71debRS^S2c0_2/5X\9Kf,T,1J/g2DE:^/2XG3O=@.1B-)g:
eDHA@V9^aa;4Y29CKL;4+0dV;)@;R]HW2Q]\6G6eYUP/\]6c2E<NP)=V3bKaCL9g
aY#<Pe:0DYT)AX?@3P;7MFgd+<1Q1LT;7EB5:+WMF?=X08Y9dP#-ZV0.YM@RCGT(
VH,3DV8=46&N+3c?]]\?PK9WfUcdR/Y6^L.D<XZ]^-/0^>33R5(#b9U?a(;\8-H#
26TbS#CU+F\QMdV&26[5LW(#0FPVPfMf:8f\:&(2]X-:K^1?UQ.##eV+E<56MUY#
.2.YKNGC1feJ8H+/0DB&BgJAF+^;N1IM<8:g/(BHe3aQ7_#E_5_:#cg,cBD1.0Zc
^WH(4^_)Va=Y.7[NRF8>H(CcA46b:eWFMH5gO4Y-DE&5VEaIQZJ3#[WF(eRYQKY[
AdUJ\7b8DO5_fAOHDeA<=?C)+c0L4+QQMLHE)8MW:SP8K6<)[=NC8M[/EW0#(a21
Z?D;,GB7\ZC<-c9V-D[G2A)1B4I?F=caWJY^^D02ca_e-J\G?@5ZSVTeEGF/TLgP
EWa9f&4K_KT6U@9dIf[.J6P-fQbH>_dZU1F?APVOQ=H+UN^13+K=d>MA.9_c-<K.
C86fGM)>?LgWHN1UN-_L=ROJ5QOF+b[>H=5+c8+P,E+LKdf]aW23P?-?g+;?Pde-
c[LLL#X_OSMA8Hb68J(Dcbc)9^@d9N;,JPYOM[X/D-1PdLQH,Z7=8,J,Q:UXF@EY
\N2&3UI,-g14^ZMV17eQ^5XT0RS/4LS^-.JM5PB0H>-N?IM<cH=TJ;;FCT_,b/TY
-)[_KF]ZER(1;/7DVQOF_W@).:;5<7B6D-V-Z,7f4dPLc84#-;N+:8fVL\[V-SBS
YM1=?HU#@a0?a/RK0UO5C1X4ZD]Wd)&5cEe=4^^aJAHEMZSE4Y=[6/BaXOa,GOBE
&>YF+Ed4:C/NA)[Q4Q^-dZE\ST:D#R1,@#U50OS_CD8,?,NBXN16bG\C0@M^YQ4\
2H554NA#?K_ZY4eAf?+)^K-+\^QU:F/2T]?7YRd0+<,,A$
`endprotected

        `protected
ZQS[&9>;\[fd4B.NH0^ZN&-)GELD_0\2K7aPT54UZ@F\gWc^Mg.I2)e=5#,3FQ-8
e6S5VA#g.A,O)9Zb<>2>3(@A78W_&Q=f:$
`endprotected

        //vcs_lic_vip_protect
          `protected
@50g1=)B<)GH;a-S5ND.^eC5@WZY7g-Uf<eY5GN^1VaQe\::HFU+)(FeO:+Ad@(\
Icb]bBSe8T2;C#R2UO&O^F0FQYEBX[<#HX#]]UOL;K03?TMVVP)HJe1-b,\M7&?R
,(O7>GSE1[PLfA&BgV9N4XR(b9DZL(9_XPLTL=VcS9>bL,.^UY3:5,,,cT&=cQZ=
,<.W#Q+&INa39+3Z&:O#X:0cH>&BTe#L1e>J19NB(PKKZ6P+92K\KP3V?X28Q@Pf
[?#Q8VO3KH?d+&Y(R0K.c#ARRW.Y17^#TT0SC(f_9WUE,8U]4V/J(F,=^Bb(G>KN
+(g8@@^FQ[6Qd&PVdV?Xb+JII<da.HKOK3,YA/K#WTEAL9=TEM_Ydg?;g60;EKP]
QX&RRPb8U\9cVTS)X9<8H6g44UGd:=&c8&5?L52TO^PX_P?d[9M[DGbF]_4P4e/M
<TI^7W@+UNf7G:2SXdX57(C8Db@G;0HK5-T/76P-)270]LBeXUacbWS+KRL\D9J&
0FG#PM1X5g/g/+]@Z\YF2E0]f6)@+5ab.V)T3<0[&DRV=,G+S3?-CfDC,SY/7+g#
E?>I2\d1+#PcCXE,7OS&a;?SVIf_HAU4eJ+L?6\dXM)04C50gN<:^KS&]W:aQ9\7
WCL<[0)],>LJaCPTd,I)e4He@@E;6C20IBg4V17I,Z;\[B\H6g.G&a1]M#IO\GC1
F2_JD-TL)B=UQMQ&+F\>OCZXB9#c(>GZH+2W=IK&0V9>dY?QeTN_FCU(ZJ,-/(/G
0/Z@b,JHZ4MSMOU=Y-b9-5JZ&_].ZCA#D25A]_(BSE)4+eA6._FQ1P\K4KIU\d?G
<R13Nd^3^/NZKMcBT:CO_#A^(16d\fR=/&[/a5.2cH@1-=YAO8&.L92?HG<Z>^W9
L3I=(1;M@I#,9:IU/#fL.G][6IR0eI?>SX0MANUO6#c6=3B[3L6\f&OYSgNDHC(1
CS(=dPMbWRSIB<6[O+3N3^@G]9=8<)M+0L?NTNa-&A+V=Cb<,K1B3F[g@\BA^;AW
,+#@fa\&2P6-Z@31#X:>7@&?L=U)0/;dd7UNH2NgAKYMXTHe6;85><K5V_a4UIM:
Z_bT)<1#ceDPA5gL2Q9e=g9#X421Q?10T=@3cdg/6FXOXSL4Z>0ZI5RI@H/9W]VV
L/6R1EP9BF:HO-U5SBXbZ;05#[D9_OdU/=-5aMBKS8SQU/CdLO&ZM)gK59VdU2K=
=XX\MS]Vd8Oc,\Z,#C+,D)8;JXL&D(#V.)_Add5bWRI(HG;==1A#_#a5((:Cf]<Z
DUE&K]+@B;QHSPdSH?eC#B=1^BY?#EeM=KbA:T+Q7_Ib9Sg<&,X_g#<D[H8&YV9e
8[LPJ_I4@M]ME#/==T49H2N-+EQ0\8:ASf9R([4Dd/<QS(B_0gB(d4@PeQ,-T6bN
1\LI#@.aN3#^X(Q7YE;J.3@K<Md3#5Y59&78#EJ2S\UZUcUHaDL6>bCU&CJ]UPH.
,g>1^K.1EHcB8Wg,K+Ag@B^O)efGQB+4^c\O<D6ZXVF,CX@(\VJ7ed<6d+^,K:,R
4D+GMa?aWNL[]LTOI@9)\_;,9CEb2V;UH\+Wb@Q1<_&NFaDAIJc=ca^^_H:JcYY@
I:ceO-4DQCOV2cP[J:6QJBL-+.@_X[+WZ.[3aY5FeUJfcQU-I]]-Y&-ObJ+UO)T6
Le>;L#MfdR(:K6G66T.G<[>^D>;?XeC:85D1Ze/E0(.eF^\^LRd@7eb/a83W?<@(
,?M8bdRZY94-EZ7RSP)6^HZc7.]H)ULBNRHZB^WHN6O]D)eB\FE&Af4,eEU8E3Q/
EOPAJGJN7.CPc3SKaZ&N=3CREc0+6>=dcfR#V.6BR3YZ@>&H1ggOXe)^&M.I-GC0
5RPSIG?9W@@/.;b;:S52NP;?S5=7GS580K?P.e.W<bP]&@(_R6eLeXLS<CQ<6RL1
G=P]EH-a7(:8c.KT+8R;Z[=0gG;PU/F2gaD#Gb13Q(4^ZRUGd:.dO>gZ4RA@L)6+
3&BA@/^aCBPM#UW_XdL4(]cfRSO0MC)Da])=d>U5K[U&9#2M50g-Nf@EKYB58RP.
&2Q<)cF=Oa?H(#I)D^BH0-^<00CS4aQ\^gIT],>33Xb>X@#VH@.N/G)4V0DL1_O=
5A&E)_MP9c2/2-G:[_,?K=(5g>H_G85A:SbP>(4e7/Yb,B457dJ=c:e@YJa=0UY=
(c?X6S<07=Z7KLP,eP1PaM7;c.=dW9OCdId9^ge2^THFJ^7&PS=@]]J;F==WYJPc
=#JP4G\51f_a[MRV@I]H6ZO1GLcUC#I_[1Y9Cg9O/LF90cU=X]43Sc#Ea5CH4(+B
E]IC:P,[<&9#>_/RBFT_I=UQ\4(&X9W?=?cTJbMeW^AEI@+&]BP7BOA^a2D\#EH+
:5=O\^]A>Q&L9X+V@gf5NIZBR]KT9\e)S>/;_Ag=_LKPBQJW9ZL3g#EFGB9K:SP;
4XS^.c.:5RNLeZ9g34b@D,2+DLPYH#ed_&AVRWYGGQ3gP&.HKb>@B_+S_V6ER,OB
)0X=8^LT&LI07BH5]#SZCUMLYWO/f;/b/>/S@a;U6Z8ea,89\SE1.82gP5aYg1MK
R6G\S3I(ZQ6D<f4R3J:);:]c1]Db;XX8G3bV2cR37&<MXE+-/-?Q#F)H6G2NU/X1
bXc4gRgc^_cCb,18-R+>KGE-/&e+dPd)c34YCP#0=9P+(JD\SYU?K;eAP_#F9:c.
WX(D9#[1._HfcHOG:^P>HcTGdcXCcG-d9)e6PL[OBRL^_C0/1[3@1dfPWW(G^5)-
@DE@Dg0a:I4QG^eIE&1D98YL#9>^/F@WI3\b0L-fgCZXD4^8<#c0<aN@I(b1gc87
GfMCK\-4.c7g2Jb:43O9&?Z7[5]d/,C.VNDQW#LSaT:32>#Z:Me)J/>bR]bd]CNf
SFN+.F8Oe_.79IZ,G3W#)A..=N9bC0MY:I38Ide47YN7W<g#1OIFFC)YYR4QY8;)
F/#A>.<Z7T5#-1[\;Y)<4R2G:H>9cEc.^=Y@4SK-]8^7^#,DFF[S^PHK>_/c50)?
E5,N>W>N6e9#8FFB0:#Q6L1D]BE&>?ME]9f=F[73QA[VV:C#:LV?)-T[NdP??+AY
/MM,^a7cWU+,F57VX&cIaP1JbdA_8M3d7^G-O1,Q6/GSafC61(M-;0BG#BBRO88N
D:a;Z37Zbg>WWbG=_RV-8=SfP7VL5C=g>e_Ig3N4HT[-c_:ENf)e8(Z]P3\XD7A=
)RI^]H)FcKW7//,T7CZ]V6RJ8O_Y61aRd\;PNU4<#C<R5CMEBS5.eC5N<GOc2-dW
J2b3VFWa=L/BT.R?C6S6?DPQd[\#;b#09bDH30.7GZR6=RY\8?AI<BSTRNf&1N0@
4d]KEF_?(NISbV=M^cWaO?0UdZ270eK6(C@J..B,WcWe?>Q?5a=S]1^O.g4ebA/c
K75IU,\1aAE+NB\X0\>U1\B^Cfgc\=-_b<[I#L4>8T)A7]Wa,_EN8#96<CR2G(OV
(+_K:-XVg7eMQ196FGPWg,HIT\R6e+K5&>[+/,S>B[\HR#Z4#&);fU4S=d6;#G0(
fCV#N#=18[C93Ea3\9ANZfJ+NE;R5-5PPb5a;.b4[=7FHg4R+DPE_[\2<RFSeXI9
7J/XFD2WZ=:MXX[@DT5c7A0E+adeDBf^;IR@@W>Q;@.-KH;O.(+63GBQe/C>b@aG
[X0Z-A^d2a]d+^MS6Y&e=42G3:U7L_S0Qa3,LY5d\cDcR4>L2J6Z5_<W1OA3D\)[
8B4ce?/P&#S]A)(#JbR&H3#g16CU<VS/QZR-:-A:<YH-?9,3bT^;g^c-=a]eM:@#
CKVSa8+(dO4F]EI7LJQC5GV8J;I+dCEIdJaLH7<F<(2NX9e;Wc[EW+_DJF&J/MM9
2ON:O4BdH=TA94F_B)f?:H9U4)[&1[\4(F>OA5&?-&;b]S8)6@_-76Y3R<M\@:8<
;#JR/J\LP1AJ;G)6#gO:2]K6g=78Jdb=+2eQc&gG#3OHK;Q)73V\A_?=FBaZ:/.L
bO)3H_JP2;R0NL?,:?+eFde2-[Q<72+SegAZJZ[HJ;)4B#e[?_8XHLZd?2Zf?_2e
f[Re;g+UXTY39bQJ91-9Z=CJ,0-)>]cHHIZUR]O8NN_4D$
`endprotected

        `protected
RR+d+8&ARYVP,[H61Q5F9(V[8)\AT#B_O]U#V6,af&+=.PB4OX3C/)Z]01B&>NBW
OQK5Ogf_JM18c3EQT0<7NJY0YMT6U6]98[7OJ&=@0\/UW]eg0VQ;@2Q/8AY.0.)X
ZNc5_0ZE]LP@BfG/>#Ob.+Y01$
`endprotected

        //vcs_lic_vip_protect
          `protected
W&X2-,&^:E[Q+H>Ud@??Ugg<6=:;VR5,,G=GKHc#B70?M3KU;cb94(1)3,J@5CH?
YUAV)UE40gO6[]=N?RYV<QL,W-YMAaA@WS)PMFBfYT_X..(^[UeVP<GAeCX\(,?5
VG&K7_5:ge<KDdVd#T2V@0U3?J<O?&#a,EDg#W)]SZR2)5Yc7:-eA_0Fcg59<WT_
3fNO&22KG4g()(4ddRfA\O<Hb5>GZII]\[V7APB<S=dYV:B.1_=#O/^7KdE(g&[b
XJH,1a+8NMdL9g)ICdXG&Saa[(97HSY&O]&T<f]OQKO9KVe[H#<99E5bYXVfJ;,E
9ICQ#/1_TNV@/9eXTK_Vg1d&LbIVY@HGgR_10a-7fNZb?</Ff1Q_8^a]R.;[.S,5
8^I50gD?4F/5X-2=G1CbFE<?&TdDEU&HVM;(aT#((6X:NNS7F[A0I;F>e2;6OTY&
+BK\gZ0YdeZ8_U#7TO8]PHJ,[1/E=J2Sf:IBO+XZH=2\K&O_SWH\]YBGBE@L5AN0
(]J,ec>[/0>RXb67OJ^D@27&/b[[6G:HdTI(H)@]]47<ZV_4Gd5>;P+A?Cg\-_1K
.[+dD7c@Z#<T(&W6P,<.-e]e[L\YJW4:2C;(@Y2S1Mg<D$
`endprotected

        `protected
cc-_F^&;G&?34KE.0DS@.VDC/:1-^dG7FeJX>>d9)T<dG)ecLMS]&)9e1BSP5ZA,
,,e&cg68Y:,;JR0CIRfCXZ8W@[PG^8@V:$
`endprotected

        //vcs_lic_vip_protect
          `protected
2g)7@_TPaF+6C8#2FIL\#NbFP2,4bSADQP[0N8LH\;(,cPWYGGEB0(X5aI9Y.>#R
^&fOF9OV@?-R;^8E?2V8C>H=aK>3=Z0ebZLE11C(B.C@,P_PL^S2P&0fI:AC&JSQ
KfR4R@=>C5ad&GR3D:<1-<\8Gb+D<g-T#J)&,Ud#Ra\7OLGE51DG]2=L@K8f7VWH
+X\\YDAHG9K:dfF0HMEEBV@Lbe4>]AB]WA.8_^gHc9[9OL7\AEIJR-3>8e32(=?T
2K+Z/.C3T#Se=PM5]?dc20T)>13NG.KDN)S>K=ULI6?4/.?,=4a(5cGJfSN,-a--
ZY:N>LC4\#GfEdII)3c-4?;]+M-Kc+_-1#CBWMf\+ScC=@e8a@FD6ND^+L82b(OJ
0:@)+TLH^I7e;T7OHVY-Yg6Tb_&ePb1>YAK8C0^(BU-eTA)]+DRV^3ZB,?ZeSf)T
XSI#,=CgY+9=9YI?^8RPKLb&7KAH83HIa#P+L^cZU,0=K6Yd=IB.A]3K)8+gLR^4
UPB+2-OT-@VT;OM5\HHI]#8/g/Q+\d]6[A49=4SKL^V/:LNT<N]3;G@A4E;4;b43
e#<&<dWg9<JOJ2cN:Z4K9g<3T0-K0/B8USK/:]QN1CcE)fWZ?SVfNLEZF\1\6bM>
^KP^H^J47KNO&=c:g4GZcXPBR\7)-<WFZW+:;#0+>E5I>.&FFeOZ>gZ,7QQ2E-;0
0F\/SSMR4eL)[bVW6+CG8AVP)LfJJ.,I5f<7?2R-+?RX9Y+):0_#f^PJG81,/&\1
2,W5A>T@RMQ(TW<_L6#2L^1<D<3H34H?E)T9HCcWP#@,?ZKNgD0f&0<9S@1fISb\
Qa4MX2\][00c#G@(7H7Y3Q,P4M?3KP95b83918?f@5]M)#1Ce/N[C,)f6X7;E5HX
C>/V9beROcL)]F>d^egc.+H3LcFE;D5SVK>L7?AaP-9.1[X2WD@+^^Rb4K6cCDBc
./F1VWFK,;VQe_P)^9^E6M,JBXAGROP]QHf64HcII.H;XOWWb3N.-Y#ID&GLPadK
/4;LE8;c9b7)(a#F9SFW/f(IBQ=>ZHRG.+\87b1=E-PNdcJ1d,9DIZBF+IGeGBGZ
VR5e^VB_KR/C9P6OPeeT?VM^,=-:c2L_H)1()=^gaMY&2?O2a>SI0_O<83eFRfB4
Wb4<R9I9P)1^]_E3+L>=KE>VGZ5\^(65KaB4\)MZSD<,)/LGd;NX<I2,()Cc26@9
_256eg,4B774O#2>J434J^Z5=Bc=f]\7IE9@@DXCF3;1bNU,dA<>Mg#_4b]7_9U#
ec:MCc@N-=2b#:5Q>GH]f?f@PV(D#Zc(;:KDFT9:TXXE&R>feg/2\/AHI7^b+ea-
-cI>^Ia7R@XZ,JEgF>]I-6U9BbQ<0E-5)Cdf#S,0O34HUWJ>F2\CDf7Z3-]=3IO+
g:@=G?T>XN1/GMO]TMF^c<2VcRN1@&=UWSb2K3.&,=LeKXV.-gbR0BN;@&Z4a&(1
.,bG;XH#Wb(6Y_B8P6)V+W-(X+9;7>g7XE9RF>L.?+beg[62T84OLV7?5f4<V:Va
:2LLZ)AD7AYbA^[P97#[PQ>bf?^gJ(UEM(JXRHWdage9N&=;OWBX?P^Ab.dV-18g
A=#Ad]:#1S+=NgD9JWRH>RU/g],;4+G6b@Z?S_L3XeFe.LX9826-TS-0YXJC19VL
YVY,CWXed+,Y/U9NKe9PXMNb.S=?L+>e]06,=0TV/[)ZW2=,cGF;aHY[):9>6eC3
,)@S=dCT>>Y=PO?:I]1G4BT+5E7J6MVEP,d>P>+X=5=O/#2Bd2Fa-.;TQYUc\b=g
d\\-#H+RV4@,I=[P:6adg>4-\-S,?0SU.C2#QQ^dFH^F3/]DD.MAE+B.eM^JNPAC
W0UDOGDG1P4\.(6Y:SSbN#T-\<2LX-(W@,c8&=IEX7_J?S7IbeZU/M&^0=L7f?5g
&:RYTJ5H<4/(3fc&LgZ7QGW3<^91_ZKcIT=;NZO8J-N(C\LOd#57H\QUYWH+QJ11
4OL=S9K@O7C;8>0,R-e#,U/ZS7JWUb3N=2FUa]U>D3b0[@>Ud<EQ:]eCRA(Q)fe.
G1ZRC<YR6UJP7DL&+^X.>Nc9HTKf>4g7);STW.gQEAN2IA;]<(8.Xb+/X\VaVM.O
R(a)^[(NC@ZgN(;9O;-9[,W+e,C8X,I?7B=W59-cAT=\,OQ:(I699b0WPY:D]+c[
DbKBQHa#36FV=;^/DI#8>MD7LXBPDgG87Q#D5Qa(fS.F(8^FLHP[S+S)V<-I</8X
3JV(UIN\HW.2F\.405&CWV3J:M]5VaM(SI&X<38/Rfe(=gGSTS\0D\a8_1JL^QMU
_@#,J7RZg<4WARJB(SR_KM905WfHJGR-6(bdb<H(?D)6RbOV>NcDO7<S,E[W&Y#Q
@]<.2U,)5+J,E>KY]9N0WK&:_b;QD5eC^;8HW+aPAL]OQ>7FV(U?38&<fH0AeKPX
:f:SV.9?[D):JfJRV9S6_P4HNPAJSM]1-S+_K8&dS93S(@9_L:aMJeJNIFd\aX9[
9<=.21YQLV<#@#2,N1H(/C(UXI\<7.<9EV)dB=_Ug\]U04&99:(\;6=I_V-0Z()_
>15GB?BQ-aT)f:H=(E>d5C8_?;&;-J/IEK\agbNHc&&eC\HeC)YJ#=TFafYA71;M
#HRFG1_]/&<FOPU^WU/@)YM)&PN;BK5aF1>EO>;dB)\@]88UDK+#O7D7R1;LO(<P
a4aWc^)B)@BI-Ce;bR9D8=Uc(a8)Q0LSOfE@:(0;)6NRRX70W\gXJFdB86ASC2f1
;,.QZ&b;#895B[K5<4V+<0a:ce9@22,PUG&1[\4Y&d^JG\OLOWX.PE/\aGC1N-Ke
)\\3?&eU.D&<c^G1ff5\[X=?-<I/3X2-[-86XgfBcA]dT[G1O=P?-S0UJ4JgHJ8\
[@]Q>]2Fe;JLFTg\aS#JCO8FY1=2dC46N-CV-52f1bRRY=OU#YXbI_;b(\2/89^X
3AbOYW+(Y3VgM,EQ(VN&IBMJTY)77]E&d<b6CAXEQ@\ZXfgX5.QcC]U3Q9g_RaOL
HEbDL[2O2T]/fKR#c=OU#^d<,TDZP:fbFd5/AK.EMPaMe5g56V<86F=>06K=?.8:
X>=I\V:aL(O,Ac.6gNUJd)cK,Ob43M?HFI.X#c88Y@GaO:\C-eYL>Dd<\@;,aRbP
1b9(PS(BV&I:?2bTaS16Y2RLeLYPKZN4\#?R-BbaJKc[.O\#-S/(;-6XO;>.^a5,
Z(5;ePCe=E?Q9^)7?#KCL/AOJ=1&PdZ)@O,KOKe3K=#0KXW2@0(&4HQ8ScgaU[F)
Q.2(T^Y,2WEM^R-Z=76<1LHG1G>OMf^#\(A@Y[&VE1ON,G;.#a#+EXg4X-EEHb5K
;^9^fP]_1f4B;G=YHSB1:e&B<cNX:X7>,^1W;L=aE?c5HX#,+@-G00f.;C.9<?]7
T#I>T1JOXWBFA3&S=B-TbY-P.>N&[^SNK3]UT:50A;^.D@dNLR]>FZTMD<3OF0TO
/WD=+0BHT(1EX\]RSfe1CG&@F4[O@+9]_DGa28+OQ+.-WJee>#eXI,E^_b,ELF+P
TC2FP02W\-GMH0C5-+4f85Qfd^gV;fYe=>g2UENKIFD#>]e&5/JO=dLQ[V=e8a.H
)O?H2=cEG@1)]9V?_M2(R/V(P_c3a->8:g1[f(-:3ARg;1?/dO>TFb9<C<ddZ6#A
)\g@EOR[\C5L#,;[<YS@7f0U0;fORS<])0?KM]_Z0a;_eP]JL4H^,L]2]IEJ=TWI
80S@?Q81D3fR6fT[#SVVS;7CVBd[<@,B>4K33dG1ERBf#2TYR/.HVC<:-/e,VcM9
T,EF[VgMH4G,7=a(OQ<2Z;@LRYX3ZMg_>03d1Q0[]9VND:+@ZWFaK=44cb2?)=R1
,OR(/ZK&JX@F25=T/R_0<+IgcZ7O)Q-,NJ5C9[NBY+73P^D:7X)GIITe&3+L3.c4
B5]:0)<CCSCW^#\N>1a+@=H[a)6]VM^,U7E;>?BP-d_(DS[;KXT)R,ZZ#ZV;UINE
;497[&:-U@dL7#NXf1=T;&8BbR>2AT&FS[8:5&B64?7#@f#+aJ7N2T?@CKaKV[@/
<a^4)9-G.?CDed)1_P82=JGEG=:.0RD[bH<?=5b.(g]Z6:e1-</V&4E)Jd?=V:MQ
U/KN(^f?.#H3]Z9S4V;4,MQ]^9O>:d1[&]X#D3gg4+C&V0](50;S5CJ>4AQ6-X&7
0g</U7T[fcR_3RCPD_Z[U,H3DeQ:HF8aFdW)0,76P?Gc[S/AcI>ERf0>QAW.+AWS
KC8:/D?QOTN?08d/C6)ERGLK92305@2+SEZPgJKcN)364N<:OC-N(>#OZV^-F\99
23R7&KY0>@&J6H-b\&(MgOM707gI18&3(]Lc/4R^MY\.T^BD],K]1#0(N](8a66Z
5=SL+M^7Hc2>)E>f9XY]>T38RZ6W=;(7G8aP@2aB#-FW-(F@;DG_K),N674UYG9F
BOOUaQ1)BA6V&dB=#9E1-RN(1J&=UE+T-B(\XgXdHE9DY6SE8D.Fc+ZVGfC&?IEV
W2R]1cK@4>M2ae.L@-E]XNP_-#gQ8NSa9V2fX=/IRO+<#1V2.]21M<D;MHB8@\S2
ZX#[@fN67a5c-)d:2BfTJEO,&A@f??;W&PI4,762HR\]eZ^8;bd1(8HE\^IFJ?g7
V0^4OY#]KU0c:d3#Q##;3g5,S&<RV8cC-dXJ6?XNaYU19K&)3WDfcM5BMQD72[VC
#X:;G\D^Z=9JG5Y>aM,,:J8V=a6VZ,FK+]2b8]NAM69CS8DF0(EdMHdbY6:?:)J[
2WM?eA=gFR_0:QH>WOGY9V5BgUWZK^8E^B^e5H.DY<g8)YS;K[2KGD+SKD(=W95N
)YCOU2W<&P;\EEIg]S\QB[&HU\Yf=BW2c]RNN+1.X_<W&<LX7YH]I<Q;X][@PLM:
[+H7:H)TYE#AV\[/#43B?A/?A_8:OCNUGM>NQ4DZ<36eJK(?KCWPYW&JeXCKd4K2
F-QF80]e8MZ_RG3#6_X&VfC/E^+DE2MNbM-,S=e4^[bHWOSSY1:aa3afA)Y#dBIB
;:^cVWB8O_6Y1fR,/Q_F@:T:U9HNd(Ia_^HQaDdCQ(K.=-(O81_/V0Y>6Z\=5Z2_
N-K--KRge?dLg(XW]SI+BE\)0+)T#<fOZL)be-#d)Y/,=7D1F;W2IZPc?G.J\bfC
HISLJgI:99MCHTR=P6O,OQJ(U==<+CIQ1Z+9P]XY>G3LN[.1/;>fAP9QHd7RF5FM
SIA\[&T5-A(5):X5e+6R>fIX2S6R8RR?BV]>MHM&/.(<LQ-/6\gN8?a-TLUH)/()
eD7(&)=8@&dNVL0:?57[,1EF(DGcE5L3CI<17&dUe\\dDgH12HPJ\Ib3K&U199F]
^5.OCXP]^7=HPEW-CfI1H8+5_^83=OH>9NQLW#2R[Y-TT5?Q++=T(1[T[BLA_,LO
IJ&0b8>W>U@H10E9f(=PH[O[Xb4X(Sg(,8e+]5FS0G2FS4Q62>b5HP23<cX:P4BF
Y[=<)+-N:])@Z0R3CWA[9I@b@HT;(.9Q2]DeL(RZ5?4L-[+\b9A5TCW._f=4BH?,
EIB:cNA_L>+K4Vg5HNI;J3M^=1.G([5^@V=2VA;G[QW2&Za^JQ0+LS]GP07?8U3H
C<2X2.b.804/c5:_8U\Ub)D<4:(:N#e)F?]&IW\7,:2:T]:aQ^F&0-++B60WRZYe
PPCaL@b]eObM02K:CVCGJaQO5c&(c/cS>M?d]UdgYg;U?KgM&&/#;:#1M<e4B0b[
Z0(Q7R9)9gb>>.a,A:6[7V&fD-\>16\[=cIAc.@F4O(O3R.LKU?>L>VWZeJ6K2E5
fHL1;F\aQ/Jf_E0gEMC4&aCGO73AM.)9]5[a^GP;H)7R@]KQ=4\QF/PKDA0LOVed
,I=CUdA&aBc@OJ-=^,D?]NGEA@XO<H8]E=]-&SS]_Pdc2HH)DJH/HTU2eWDLN,+\
=,K:_;W_OgV4YM6ZfaK6bS0YX8B-=GYaFaPBS.GX>9Ea+G.BS;I+BcG7N_RIVabd
dWKbI^0d[GWAg&]c=<TfO,<c3_12bA(^e1c+407K;]/3#IcaB3\I<9R#_6c,7CgC
T16-5.?5Z,.N:PKQ-6@UN19+Vb4>M]YNLSGUJ4XUcGeU\C:EKO.;&Z6>H]5I_;?Z
C-gM5Y<.=V+2XU&;,\@=CE]4+eFIM-aLVa,@(KKXHA]GGK-D:8>]W_-MI-3RO.DG
(:0+4^]5A@#01Q/6;/MFQ?&I0<+I44cD5=c<NOTd)bQK5cO.:&GP77-MP$
`endprotected

          `protected
36_A-AXB-LEb)JLFf&_5g4>6PeHW3:#GIFBYI7WPJaFcA44#e4B<()C74-D.Q:QD
[?PH:G/)OL?7B0-RBO._&^Q..BE^HSD^>$
`endprotected

          //vcs_lic_vip_protect
            `protected
(^;G2N0073:6aGLd?/EE7Y+dO/Y\#YA7cgESP-W<[I&P?DD13_CB4(SR@CZ.7aJ1
^=QS]/E>VDQC]UP#c6gN:FbN<aUbbD)Q=.>:@LS@390THfWK6#FZ0<EfQ0DXV>@7
Q4Qg3DH8GIdPEcXAV<JBI/K4Bf2VK=,2?N=^)ZJRG?1Ef\2QNN1,[b.#1FHcCH6Q
b)1gQ90H[O\QgddBCg^Q=LDDN+d38<c39](c+DTf,A(?ILLPSO.=#J8C&&SD]S9P
2-2gg&+QB_@#da86d-/g&3E7D8RYId_Q)>ZY3S-94+8c3-M.9Z5PV3B.dc^_^TQA
8ZcQb49\NRSI\Xa<fB_VVg\:AdAIZT+VBV;3L3gUD]P<bYC^@8c3b;8?;18#)1O)
Ddf8S=PSX_2VP)X/MSH<E3+K7fML+bIXQ<1a33=Yg[IP8ENI.9,b?Z5YE4JW7>,A
If;@?,K\fJAP]=@DF.RXV3g-UC3B#3:0,]gDDHQ^T+4b[cKddNf^d,PM@W-cTbE/
+ZEVX]Fa/0NaPV[270T,LX)=ag\-T::dQ@,egMVN,T<M@>L(<J:^\U#YAS9e-S9V
=@Fb)(b_GAba/$
`endprotected


          `protected
5(11.IBTY[^WTJGF.^(UIVF3SGV>IL6&?5Q[9;J=4DT6#(-N=:9I7)=80\28ZHaT
H]9YO/VaC@g?QLV].;LXce4G@+gW^_b^>$
`endprotected

          //vcs_lic_vip_protect
            `protected
46I]S9<K;J69I]DZS2_/A04,YG[_]815MHd?6XD7@DV@FXY1K^7#)()-CJ3dLP:0
M[g/4Z9fRZN]SZ[/^^HK<HYSV.O;\=P/ULF?^B07[FCBV#a0B9]bEWbIY8a7KVXM
W0;-Zf#VGa[>;YH&EHQ7I]A#ZD:PdSZD4,E9<6Z(0d<>SVRDE):QBFKTH:c84W1K
DV,FRH-^adGD0.6,7/DM>0]MbI8MD[8bV<1Lg18F3X0/CT:(9ONG=CQcB_d8gXQb
U4N3(=D.ZS.>H\]:CVO&cJ.\(F_#OAIBKe7Rb<+BbZTT?Pg>Ve[S:5eQgCRQ+@2P
9K,K41MPU:PdTI=4+L-M=685#:dU0(^/Y#6bec,US&7abU6TS.6#GH-@S(6K.=<>
]^0TKO<?G=I-O/5F=F)CGKU&UZN]GO1;UOS2CJ0^S8)B<dNX(:6Q.BB1C>dOeD6c
-+gB_RAI/F+44X@<b->SNL^WLW<X0P]g9#_5=eeMa-f7_d4FFB=+<+QB>2\a6,Z-
P4-Yg:F63[F[?\L5bGD<-^4YV&Za,_&_WV)_1^H;fPc<D[;MC()9-b-\I>[2Le<A
1MSNKIWFg;57P+XJ-]\aPc\O7[N:V\Rf?O2&EF42O,-^,K(P+_[ZIE=7GB;N/^fN
[J^F(<5=C[+\GG3W+eaP-9=8_g@d[Td7c0II\bb4O16a2A=b.V#I1b4C8e_CWQU2
#)dUQWV29HWG\TT8\aKH/ZEDg6KEDHgU-@E\9FaBI(\_e(:RC1YZ:5(+,)FY^4KM
2;71RL1QZ?F7TJ&T\R0;FO<217_RMeXL;8^N<F+Je&Q;C:+9E>UC\<4M?VMKJMEF
(fWKPNNEXK).AR^&cV#YOO:)00OF_V8GJAX1?ZWEC95@f1VIeTbSPT@C4[YYW4=+
BC.6c1M:5>]YAORM3&)+_R1A^KV<5&A1X:&@B:90-9&<W_,(VBIJg7g,J6M@>b;^
TY[S1B=>I>5J92E+8S,:=;TWD[_FN>,&QOZ&W+MgM/,P8NY]b-=:0HLA(CPBcS)P
c1dPJ:AVA8X/GJ0]\E5V5BMD:9-SJcOfRUBN+,ZTHL]UX@L3c34?4cLPb<O(N6AW
L+C)0Gg_43]fAX+eY)U)A/OVHgFAZT@L1?YY[6Q,Y)X911(B^Z:+UXATg?a/5+<3
T]Y#eb,bf4Bf3-KFN+Mb-2@C:Q,=,BUULFfLBKb0ESd#)ZZT<#3A<7+=4+Xc4J:]
0?FZ@8:P[d3H1-Z)DM/06gW;a+]\JObZ#B>9K(I?>GD6(6:@e>K]e5cHRYb/^F[C
TA.^a+A^;CEaRXWLAG\,.UO-48aUPaX\g67[3]gSPEDdO/WM_0V[#HZUS_,.d-3_
eSVL^A<N943#._:aVC4,JN26(T-bOX4+aGZ(d+(ZU0X+BceZ7(f:)C06P,<6Egfc
a;.\6SILIMN]D,\59,K304H53G6-e+B9K0XN\TOe_aM5V_0<0&#ZGRH4c=G.9UQ7
4&UUY>_Xg38<[Yf)J451\V68U3CFL93:@PZ6HIa:+L6NYQ<[N.CcH5EgG2BPLETM
U-N#UR5HgbK4Z6#Nf4FZ_^\aTXQZ3e[IN\L+2eCGD7R5LE;E^H<FDG>T;YLD.dLL
S6.@_C)\eIb^)J,^d:/+4::P<4W.[)[[Y@a7=VV.GF#6Yf)PT/JU&W[=YS8L@Z0?
[1F)#c01-BC@(Bb.WST(X0/Y6Z#\0V1(53QUSDI==D\-FE(?dRK9/W=>9e\Z9FJT
5Xb&X[WNOf0,,V.R9X<fObV1bXD)YAK4?N5)K2e:]Wf_Q);8#Y&_\b>N#MI?/:,@
-30f[.B\32GK]a0(D[E=\dcG7YL-MTLeT1<1D79,<Z\DZ2g:-GJ)@8#/6U#SA#3#
[GV>8c(D2=+=?f/IPY^J2-faGD&)N/fFP\LJaRO-gbT>K_+:,Y^XV]fD8,gQVD+]
8=4?)^f=Z]GM0YCQEG0XN9f0a2fd134:)51;V_UWM8[4:C.IbJfUG##=T9H1Xc3[
?#=:2<F/4&@c+\#:K&)>e?/QJ<MX3-9fK]W.fCRbHdT\AX_OH+VX<2eKXYO_).^J
aC8JWDPg0)&AMdMJ#<WSC?SP(,R5:STPf8LIX8@QE)JB[-VJe[9/>AQAaY3LYd\.
4NQDJB<Fe.VQ#^5S.S?;-G.7T4M0,X60bY>>E2:8_ED6dZ]g1B3\cdTPR^a#<I)>
WGScSS\dY]_<\CA/=3#8b(3#N;-]@HEg@0g9?b3XKXcEF#6aLH5EgX2d;;]^Q)0-
&AC7UNb/QX?X?3&5SBeF3QgZ:>c^YB)&\+cN]0_J(G_V&gQEfE5(F>J_Q-PgDL?F
R32B4Y6a]A_4FK2KX,#-J.BRR]-PdQ5Y0KUbERX>gKLHT\c\=S^\2VB:^cb]XB/U
AffLQX4I6eW&3C\1^J_:74YSIS8=SC1N8<D;7DD_bNJ=WBAJ+,WETH?33eKHI=Qc
)I?RaR1dUBB/1,:.RL.<1X)4[^fSU6F-MPQRE(fA6PNb48^477[<5/-[b4OFV93+
\LfLC=@MWZDIOaP4^4UO16Z=bXR<3X>(_Z6R?_U69QXaJ(3]7faeOP91^2ISF_OB
6],I)80AD-HG0HYMNT&g4\KQ5dRL_KV>O57#CcZMPEX5#^3347g5Y.7&,I:_5YF6
YC0[:LEa^<FA8XcQVZ.D,&:C+@gKFd#c@OO^O^gVON>K2B0ZcdAPNLa7g:8>[_Ab
XM3]?VNBQQ1gB[-<>>]1)Q/B5-OQ2RB^3^E[M=YJ[7JG\:eOM-cI4^Zd/Z5@_@N3
RG2L2,B07VDJWcL<\7SY/:DV:>0HeQ5XFTX-95g6Ed+A1QIaG7K/8ca)#_S9OYT9
X3[RQ2a1G48J,$
`endprotected


          `protected
cFR6BY7^3<XeM.9AQ<TH]bKQ@D)\N-X\^2:fF.a7^5bB[/JdXWdE6)d[;F9G3f3)
M5&2Z2XdN=)W(,4<_8,Ub2GXNL].gFT>#4Egc<DJ(cYBR,J?MQ[[6Ad[I$
`endprotected

          //vcs_lic_vip_protect
            `protected
4C@:+Sf;Be3+=3dd_B1I,C7QfD>GTfCDXYbU^8#_L:Jb#Ub+/85Y.(8bJ,S&_L.9
35WOd1O&.99^A;af.+.7)428g<cE\E(,f;.X@66>9g/J_\I1?15&Ab8G.cE/.IXM
W&S:R7TGcO=^BF(<_-LKD_:JT?8I2?A1051eeFZd6<07?GRC:ZK9][/L&;F__U#c
Y:<P,CL^^DF(^-]H?cZ=\7YQSc3SeV3=f5-cPL5g#[^>-7QB:(LUgdR?#)_Ff2ZT
MY/^=gFfF/[S9cA9&):TJEBCcU1PUP/W,P0-GI6V?]>YE^T1CBWff-5,D(CFY6\G
JRFZC^59:6\gH^9[UV.G4-P7gP?VXPF6&)T6AaA9g9/5N^.f+XI.e&@QU7@6M,0S
3N6aG(G7LOCHC3)=\QI:M20/BZ=Ve:C\:&d>Pa+W?A/=A&[M,X3XGb+9F4NYL0WG
@,beEE=_PXQ<a2-1^E6/2U3V2&E8O]]bdO>bEQYED20d01AVMRaZK5_fBQ&fNF:d
>PIC>UNVO3/J3D(C/7GDc7d7?<-01?>+C1?OGe+)f1QA,K[C/gF4?_LIN0HG<dcP
9RC&/=YGb8?cE=K:f;3G].3)_eC2LH@WJW)\M[+,@gI4TH;5=MX_Ud@gWIW;P;GA
,dNV9\9)U,&Z<\f/>5Q[P#0)/CF9AB]eg:L)VL20^\eDSVe@@I]O)TNNOU84g1-]
F;\E5M6S)[Sf47Uc82c>PW?G1/-<,K?L\MeO+J^O_N:d;]#:.XcdAf,JR3O)SY->
bTEf+)V]fGTP[aXC3)De3&_bX?BdH&R+1N4;Y:DUg>ZUGbabdF^WU\_8[C)GUgdO
.Z9T>2N:DM?BJd5ME8_WMFYXVRMfMV,1V9X8I-W)LR4<f8e/\6P&aRC8b:9EfZDd
CRFQL^&=-9_SREPB09&aN>U=\H.2bI]Z.)F-&-V>#=_?eNP)F\bW&<3?R3=TP]=W
(V]4e+B7;<N]b8W5D.J9:4Q]MVgA_&R+#4?\d0#fBH&;-c>4J\7PN-_32XL36Z(<
&A]_R)C#_\T0K/X7J5:?[V23Q>:Q<HT3Xb3.>JPOE;/;IH8LD)NYN(7XegZNa8#7
FZc6Vc213HRD\J+XZOdW-)a8>[QX?5>RGD7daQ=G/Y(=4=gHP(-Zd;9FJ:&;YG1O
]-BTHbQ;M<>V9dcC#IP74-<c6T/d6>7UOO7b:Z8\5@D4a@_A&eJb64ON7ZV.O1\U
#=O6JX#;#]Q(cgD?465L/1WW^55D)cf(5c?+O#/7.)1(KA5PH)?dI=B;9MB;)JM7
6?^^B>SU,3<-&ZW2&@X><,>QeU5VU-_Z@:f]dD#>(PGB3497cT\:MYQZc9RF4@CD
O()N=/NEcXENMJ<IFYegBZV0:aN@]@;+UA6MK5Tb8>bbF6ALPf>Mf]M2e.&^K@^0
.4VcUV]1Q?;-dP?S>.+@X>N0G,A=SFY)5gF#ca=Q>?EN<8.5WIS5BN&[Jf^&ABAH
]39(HR6#Dc+0[A[TC[PcU:V.@@3_P[&[D<R)IP:1,SR29>5L\PNC^O(dKJbFSBS7
Z8HP4@Z/GgCSOO9B1H#BM\COHaKH-H0dCFRU<0ec0\T:7Pf=3OYPT_=3-B;aI9DM
32Q?7[,5=QZ9LP?=SC^]SF[IFggFFD^\4<]Z5?Qc7d=K5#[<P^-BISKa=B5A#;1F
@.+A9L+MYP#-FCGXDVCHS.2MU=L]73d0,X_R=B;19XMFN;>Of:YOJ;G(FbBUUa=M
A?UWSULgE+F7,ZHHDb)[3FIR\R6XVV[2\.NC&<9DY3=5<AS6\RER2WTQZ0cTefBF
T@V^c8Y:B/1(6^-6(9(BXRV-adU>d6K&Z=dbMCOY.8=a(6M#Y@b<CU?T12ID7JeT
RLUCe_L<CJGS^R22^I;_#e?810_)(_Od@2N5M-bRO7,1ZJ4H5_J[>2YW8BXP49FB
HcCH_4X(X8D)^T.+-9Pf;P]dBY\_WGY&4Ya4:#<@MS.?&;54#WJGSLE-bW7@AQ;J
ZSX_8VBJW2,[K_H.7:X5;LXIO/[97L?/-=:RP8KU#O/@8@ddYDVe3Zf9),.b+:@5
eW9#X@BS+5-<P?:)egW]d:-N@DK<a@1ffgG,F@7&N>\6AJ?G:LNITeA6+IUW[Yb.
@@M#4daXc1Ua[::YKB=>B3@CZW.:B[..eg=/E.c;aUUG.e9C2J0ND+L=\SOVa2M(
A5DGFa=dYA7[Gd2.7>e#]JKO8]/AXYQ?c#DGeVcbXP0FRD26F/Y^R4d:D_Sg^486
W\@ASgNU#1FW\^>4=MSB>RQ<+M0)N)NZ4(25[QBC[&XX>:0Tf0NEUb97=DUWWF#W
Ca5(/3baG9f0[D<2+WaHUa[dI^g;Da.&4FM?d2T^0LYY_#,_BVd<[E#_]2[C[G:+
^[HY7A=O;KZ/-KBX:9Ug:72N5BcDRLVH6G2_gW,bg2Y=O&LM<8]YJB)F/0Ube[B3
#M]LI^7-A6XJ63GMJ16Xb=KK]^QZ)e3X3_S+A>M(H>&PR>MgE\[M3-3\?MN;:U<F
52&RWP\Z4-^SZ/>&d7G2d>9367eH9Ebc.(eR04^f,dPTeGPF3GKN?PIV^SG61;2W
5[7Q30><&+>C4PI?5Z9:5LN,2L+?PG@JcWL0]M0>NdOLP48,=IReM0b_3Zad61RM
5Q,BCHJa^[-[<SA<;\\Af(<N8X+R,LM@T+Q9E3J3aQN_6C)#XV0eNc^6e[M51UUJ
K@JK=\U4K3=5&O5@41H1,XFKFRR-N@FfTOM@8^,:52S=cCU)QU3T9O+a6FJURg_e
Z)4:M[PQ#8W:6OLF=#^d>J==>E&O8bN-]FM,Cd)#FD-4,YaPS>(E_b+_&/R8HM[(
)=^J5T]P:R26)Dc:\IMP?Q7K;\F?572K9L.fM5+?fH[ZL@egR5WeDM^Vg62\IT\)
Fd6ZFbaIGe;2#B3>&H^Bg\JLAgf?4^6=O#P-d@Q.Z\NP\H/PE9.Z1FWMUS-7(>#F
ed_5Y5K=@;P_6-U<)_RWDKQ6QPN+90=)&Q=5RA>YM:^XE^Q\/</eaEU9\P7A1W]]
MQ\S9_,@EQ@,9(;Y//#UCU^SP@A(.B.#dVFWYXBMQ=;4g?/V5J0;@;_Qg03X=U<_
TX;9C,WR[L&cDEG1#4(=V_eJ]f@.=CRY:e23O(Qf:CcOaNY;7&GE/U;\3,8O:DX#
d=>,)ad]c4M3_@.#01\)=K2E?,d9Z#gT0/=5;8CMRg]E@,)>a9a@?FXIYQc:H]@c
c;J:IWF/1_S]dJ.U/\\NP7J,XC1P::81R4MU>MOCK<B9M@Vd(<NN:cUXV_44LYOR
S4M>QWVWYICQeA&0?&F:Egfa--2aBD8adg_BgB>N4>LP.KW9^e9g4A#[cBQM^V<0
12ec>cXOVdJbO_G<9GX\7WIP=VZ5J=TAf9/3>_A-5?Kf3cf4.;0(Y?_WH[..2Egc
d+[#YXX+/Qg4Z3=+&.WNOM2GML5[BS4KL[G^a/J[O5CgI_]-MQ:0Kd@+1WL_<[)V
-/e[,B#03gH9WAP]#Y>KS;?FKUg[DR?gf7S:T/5-[NV8SUD7YdXe1W7Q_H=\/]EY
/R1,?86:,-0.XI78.[Q^8b.efb@A3dUL4YUZRA&TN)T5?_fa&_W_5PAP=<T0T]O-
Y#:@>-ZRS;5RWK?)4)YX_<[Q4>WfR_N;C74TTFPQCD.<CBW/bKOTUEPBCQ<=\W?-
2#)G9;CE6L?d_M8056O7NY8JJMH5]=WIO4YCEbXC\6D,LOBQ(bS<aVPKOL^.,\Z\
1<H(5WCc(5&TS@&>Jg<M.EM3F2Ic=e>?4YbC0ST.4DI:M50@D9M5\8,&WN12LN6d
1^T>FTa_EDMcSZ3^SH-6C.Mb(EbJEMA]TC>,F)aW+VZ0S[<fa#>C(4V.?RDF4N,2
WcES3=?B7NbEAIJ@T7dNCc)F1;OIRI0[aQN(61N&6B<=RNUR>4ELP[X+I#TKFH,N
gT#.[7:H68HJI9fe;.TQN:aA5fWcWM_Y427]]0V-,5HdTdZ1NS+UC&\]&_L3C3I8
F@L#8OUNFV,=<)52]^.C05J-ZZN9LG>Z<>AZ6:A4HI?(KdJT\[?SX#A&:M=6K@+I
9@K@.XG+_\;O_IMD<C(<4C_J?AZ4@.N45R8U<aKBF=3JG)<R;Z,Hg:]W0E?L18G^
2565:SE1?N7DfZ@J(LaG(MF#]M#:;T>?2U4Ca;#(c2G2AI/9D,&N3FLPGXV79/]P
A&05:5039&cOM?^Y0)#;Y<;WVXYFe)/QcDT.((\2;//Wf_BL7-EHS_05O1:R/HWV
NTT_F1ZSf.ZHXSH_:.M=N])EE60Z<a,SBK5U?Eb(=E]W<5^;>FbS.AUfF_a.GePR
Y6@4e0=[fT8[PY#OO.OMR<[(dcA60]e>9c.?f9:c_a6cF(f#CT16J1T/0UREg/7=
G6O\XUHV=3d<O84gdS0H,@C/cT0e1DWV#M_YgGBa<W8<-J-(]Rc^d1LMCD?Ycee\
S,Y^T8&FR,fY[\RSXOUT81=K#d3D+7GXE)2,H\aXJ<56B,DV&Vgd3QgI8O^+dfVE
d=83?C7MQ39?/L=TP.Y-P(4eD@HS-YD)V\\YIc=PQ2A.OIW.5+eL>M^_Ka#.PZ49
,cE&)[a;_(KBC#e0]0.)O(6S[(.fGRWg=_@LD<gc@D?bG:bEZ1GA132>YH5g?B\c
)RgWZ<H]8eVaE:8@4IcG>I=CISY.9N.@JDa-EQ&a9,Z;O#\Y:T#TH-5Mf)=X5VGN
&CVU,SVQJ[.;&.DSZa40-)1WHF)?CaRbAKM5QH)9YTFJ/Y,3VDc_,/C8N@:<d+f0
(S:>>C4^Ee+B2Y6JaQP/FU1acD5KUEGDf:YDUQI?2VCe@UEC[EYLdBb^QR-8,S_]
c;CPVZ_4g;[Qd&=4F[L69\bfM7R0XR9;_Wca=N4N2If9FMI,AbB8_eDeg&N&(/7\
J\(+8TeDH:I:C]4,M,b?S24OD>a@MN7V-ZI?CD4H5:1c&9[P:C(N.ISU]=OZ/(U<
->&F:D;BAJAL6#cA7Y]Rb]9#TNB.VQE1:19R0O.Z(GI-NMYI#XAd-KE-OdgdG&N9
fOC<9KCOZ\cIJB6][^QN[>DHJG4\G5b?>_440IT;SA>AX>Z5]2(g1SN6:Kb5+,-,
UC?A0a>NZ1(#MHMMFJ(fM0HA8P3.6_7,8H:7O0:bD0DDS2.0H]FgI#^C&EQJM4LY
T56M09YBZ.Bega0<:c10+LbTH^-K#W/Y,E3eVM3P:MP;W7]8e6=7JI+TF^30#Wf\
BW):H)J,\I&9,Q=Ac?3D6&JVDGJOBJAM\RLaGfZL^M)b=fWdM9/RS(A+).S[T_;G
Xd9V+;Q-)1TN+<5-4DfbAY]d6;<CgAAfaL>5ER9CJ1J>DH-2W,J_G0G\g7E@@OJR
.\2E.Cc7RBP&5WADGdS.5UC[-,9aGHJ1#+3eOOYH\4e=8?CXC/9GY2:Ge4:>Hf0(
9(:X1#)LMW@bc9EFKaGdIT)>HGISgda?)dD.I@AD_B<RR4\ea(FM>:AY)fSX\:)P
2HfJ2X+VdZ+=/3T03,ICPTaEAb]<=Y5H?EQ_G?.eFU[IW(B(8d_g)FC+7.NQD=g9
e8GO6/;#+b<L<GNDAQB&&BGZ.&O]3WN\,U,JXfPDE5TVfbU#g(3^(e>YeGZ>#SM&
S^AVHa/14XGcCcfdKXFUO\:1MA(0YKP>([DU?bA\ae67A>WW;gUU).e@#,-c#IcS
--]B[RKKU(=X?IV7+@gD)(:WPCJ?&Z9WdLQ3db8N#Tb(g1e&NeK,H914SN&?6@?@
UUANN2#166,eVXgZ<3?2=eNCV+M17T)EQ_,)ZQ\FI3<5YKC?69?Y4LFE19K9VH)b
Jc^R:WB;IV_Y;PQI0R9@:d9H,Rc3^Y<c=57^XYQ=)egUY.Q#2R;Tc7Z]=TP(L-L@
Gg/b.L<B[=E?,X^(+ZZ.@/@&)\AY52_PI>^6WEC]fRf^^GD:AHLS+P:ca.aNV&P6
:).W+7,_^M#\3K-M;3LFTc]e6YRR.9X.)>-G[7DXJ@=BNIT\<fTT3=3S,[^PEJW5
<#9#B>EX9;WGG>XP-[=R8I>T;<1eJceAD@N94CdQEdeeb)G))PFaP7+&@:GD:#L1
0Lb0DQXDfUO.OAaJZ.XMN4Bf@1BTIaC<@U/9M+Kc?K;M6Rg.R+F_,EK^WKE&Da83
N(\DQE9E0Vc[\H9N-XN#_[YJ9^ORL@dZCc)+a8]57YS5bX?WV.>386INTJIBO(gR
eKa=(NJTBb.caFf<W4Hb.-7SHfC^>YV+OM\#CW8&RP[<S\4Z/-cggCHFH8H\LA,=
D@9931PZfA3ce6LZZCR3.ac8eTHP(8HI3XW[.HSB#3bKc+T\G6V;Re69X[d.2Q9X
eA9,I0NdH?Y#D()&-a-;,)bO\Z1<;UB7_@Z)bD<TU7/cHJXFgN9@gO[M92:b[^FT
Y3TF[3U^@Z6dEYLE0&^M:[G?\.DbDG2T+9P>Gc)J,^LJIHT][gU/BW^5e_?H=A4>
K5059\WCUCXBG^b4IL)Ug\,a&d[E5bQb1T\O&X):HgR8TG/Z2(O55]F&?:+P,[\_
(gHP&]/D26N@Gf7eIA7UDcbTdKfE+(RB,Ud0AE7bLBfcDKV>cH(Y0I[A?1KIVL=e
N.PcTBC4ET4<.AVJ&P2cbaJODJ(T^87>@PN9H17#52<7f<2#S@2TOS9]<cZb;[5<
\O;H:WGKaGIBc81EeSCd:DS=M-7F.(I94-PC3fWWTR2=eU\[/ga@5NbGON=B_Wa=
=1LYS;ePf,).:8;DZeE6)/BYYGe[Y#W/Q0O0P&b<g673c-Yd,.A9-+EF^#&Z;CY3
(<\R]1H<Oce-f-#H4;\_^PMNNH5.O)\NT8KE#M5[?X25V<;3[LX_C41+Lfc=#OHc
D=aE2GDW9YV7;QY=\8.+8GP+1X-(L)J[DIFQ]SKUYU>ec\UPX56R=-bZWNA+F_aY
@&IX]8aQ7798^&33RcH-P(\VQgH@J4.8]D<XfJ#A(6JS?HD?/XL]cWUBce7-K6P?
KeJ447;D?MBdQ7Nf)eRY(]US[\dfHQ4a&dD4;f,<#@RePWUK-cZ/)<QP2a:C<L5W
WE7C315EXJ=_g=;V4T5Q6<:NB]KIRM,[cT)Nf2I5^@?&C(99g2ANCK:/Qb52:3>d
;<R+3J.I6[>/feI5\IQBQ5_c4N5:X(TOJ9&BaReS+2-39F:8CU59IAI9.:53H+R3
R1ABOE7_G((XPJ^.bEM_:Z:5PbK=bB-V[M,TC])PY[:R-Lg,27&X,;5XVb_55#:c
7cI@]W(=,TbKKMO+2UIeII3/;bcSe5;f8\<\=.AXA17c#J:\@ZfL86.NUQ,30SS#
P3)PgKRBc1=WK::)3G5.KW5#L2fcAGW>]\JVQgJR,\aNE)SW0B=EYT?;?064=QU\
O/>9N1/Y,/Q1#+dB&HA<L+;#\]c+^1#);JX/_TDD&SUOVI9A@fMC^1ZN+VC0[1HB
/JQ(P=-:J:T:/.:gR6e=daC#S6D5=F1#FbVC72;&X)c@X9YE8V5]R4QILQ)V?dN)
LN-a]6V#c_d.Bg>>NggcY2>:N#1@\8Hb-c1<D<9F:U9\/.G^e9UGKWRO0U<QQ9O1
eCWY2CYFADX<e4RLQ/d[KP(b0XPKE6_G[A0/TbXe3NG5(a9b4+R<UOX3@_61Kb2?
L.a5OXR_/EEER,0<VRIC.Ac3IW=\DL\Q)+d1KP7FLcZMU_]9ER?Q:26Pcg];WBQK
J05E[^>.A.,KJ+JS>#B50,KY4+I6a)9UC:35PKQ61\UWb)N&U+YT..ZMPLFRMT/3
/1dVJf<IF4O_PXTGa]#-3]?S7ICOC:@KRCY=8C;M12<#;H\V_EbMWX6.1Z/]::]8
AJ79>Q1S+-2(W\T;Z30LE.4gQ5_I-;ITg48PW?gLC/Z2&WT]b?VUR(EeM;\5X.QE
2^@J0f\JD&MaE-V?dQeCMbaI>#W.7VTaCJ#]/YB<ESdbEeNTeRY[MGRT(3<X/GE#
G]@G,2?J#=MQB9PJ]YNBc+gBKAKfLCAe1>J9(dg@47]_)ffFCK59WI25HG,Qd](6
;c.H]dU62+N),+ZPaO>\O5GJ>E\&,\BS6d7IL6EEZE2&9_N86NO^S:eC2;cSFWYA
KbNG@W&K^]b?I3396:_38Edf)92EI6QMeN+c10,&=g]H;&Qg2Q8Aa01NS.ff+g9U
,N_073/W-(cdZ/47X1M#W(HZdPTGE5F9XK^d75VHP9\B?O4G#CANe-?;2B/U[9Gd
AdbbH4A?PeKf1Z5J.C5\,T0?aP.FW7=V4LH85+\1cG#&F+UfMMM@X]RZSIf>Q&LQ
@(_=&Y[X4RT\.OBaXb[)=.JT_P=7L4]+(Z(B]C,f?U0cAY8QT_Ec]C40E/@g/R)&
]Zc3<1Q2?I&HOJ/PJ&@;?@AXPNAT^9Mc;9J,3Z^Y=H<URK35_/)1K-)^5IL@7M9N
O^gB^;VH)gFF8J2EfGUeI@=3[c>Cd025=@>E.EcETXQEZD9:8_/LIaMg+(?[]]AQ
90gP;DZgeb)>aKSDWVG_I-Ma_VCL8.4/J>>:,VNCC?PF<-VNKYFK([B;I)X@/ULe
L1((;S42,bAd7TMgP[S2@2;DX1&Q3Q=bQ1WTaHUQ67A4F;^(C4-(9UP],Z:JMgUT
eQQfZ_67;^g?:D7>PO6\).YXHg:DNSfOVX>d?.UdgY::R=0E&R&3dcBFS\7Ogf[J
g4e.S]Q]7faJf/4JXI[gV0:RPVAGb8TU.J,;.2]<E#0/I3BM-)Dg?N(UDa\>P73G
^;#]ESRc@\La1>;5/FB8F0N[0P,\EA]f,.dg[.N<eS-&..(aMBH#>)@&g)c=5>)<
Hg>4D.I6V-D<LDFaPOY4J0aGI\?e;0E.2a:JCFPWSg)D)3WZ0/ggcW.L[1g\ZeM?
e4P_:/@G/T<>;>GeQ#e6PCAVWOYeA&KW)P&AaFbB6Fc0F[7LIJ16/F<Cb-bR.^)O
F91Z<K);c/LSOIa&&1.EEI.),EDKU-K:Y1-6A[1,7V[GN95P=Db.(.]_eMZ7cS,c
K1/7d@[@(A@2UH9g:P_1UZVHY[6WZ0H,aaZQ97[Z@#(dVE)J.&;PVK^VGV6F&[(e
W#@Q)7W+)4aeCJd8EPM_OTZ[3_1,[(C/HIHA:QeGc4F)_6G6WCCFR?I[J4)6^+_8
3UVbPX>D-fg#XZ<DI?Cd@3LTN(/F@dCW>/#5?>K)f<]H>AfH]7Wf1C[.L2=[E.Bd
:ePR_M9YK^6Vd:_J9(6?eUc4F/U.d@0M\VX0&KU2GPQ_R1ENAHR_eFIO1e\[-;:/
GQ6,gY7)IN+\[ILFXJ4AUe?P83CBH18_O5ITOU4^BB.MU?7FfbYOKK7Kc+eRBX=a
]>FU]dDZNe1Sc-#VAZL9#NQaQQ]OQ-[BJb:g^6D<8ALMM;F-K((K+5PVZd9UeDIV
=/@.+?S4.KAT[_3#+TA</Z<W<f9LcDS[DKg>]0HRIgO(SBNPOP]+7\+L;]a]=W;>
XPf/=17b,Z:N1-#O]?d)fM?#/:^P-HY#>^FIgD0H7P5G)=27<.\N(\Ba?C>DKI(O
9H&2:C6&.LF^D&3eObcW06Mf6AI>[R3GU\FD+DC4UK\&8MK&JeP60-ZHCWYVB2YP
7#11WP2;fQA\R(LW(SXbM&)9+KZd-#8>&IbYYIH#C68<\\N/Wa=+0)\M5Q-8+g<Z
I@b[PbRQ)NMGJ4-1JS(T2QbF_4\>PL@Z05Mgc(@MP<XX>7I7_L/f>5SaFK3&=G8+
:Id8P\8,]9L]+Q_SQ^?Wb92KL0E:(YRMCBR:#Xd;1E,=VSF_F\2;9R-g<=+0-O0>
XDMP^6NRJN>\:/_/WXMVb9.0Z0)aTf[5/XB75<2H45;<;40+?CC49VV<1,>F=^>=
;cV91#ZNER.DSB/5H@W)S<a9^d(PIQG1c3?I,ZE_b(Hd?W]eR+WMK>D95>]@9;^4
B09T&;4:f<FH+]US9A(QMJ?)#LP63VZHK[._5a#M1@NG.KH9ZBIU39Eg@:Qe7g:/
>L>XVO_R;Fe_Obb5+E@K0Z3>F,--#&:g\&\a2(R0\^0LS2<eJB;9E<9++>)RF92c
WCH5HO_cBA.HMXbU#7F+=UAD<9AB\GTe,Z+DH&8^SZXbIIWg;H-E6>Q5QFQKV[K=
Sb6JLD:c/_W0&;F)SG/CBX9e\Y)@bcT[RO6=Sf\OFW35KE^]5>ME[I75f0##@DcC
KY9N[H_YcB3MRIU?X&,<SHbB0W&HE0ZD05/?M53WcgBY.ZR2L.Z<-DM(>^.XRRJ>
ID6IL5dc(ea;)?KB<<e5YYZ9#(NgaYYdBXN]S(Bb<^[eI,GN^,^RC:9dcS8QSOP)
#R-E=R637c9(TEAe7,@FC.@Zd7NDR/0:PQWfNOFNAa]TOAZb[320_L:K.ZD^HUO[
4&-8^E6-+VRd:J>dUB9>,B>-bCAW?dWTZ00f^9d\;1L?H<3R6YaL]B0Z=2fdAID@
G5(N<PJ,6<6AfU^@C+QL-]<O-A-9=P_O:L]69;N+34;#XK3,[-Z1K_bMaP+,#IKg
D)e)403B9GZ\MbY:fB0DXdeQL;eMfaI./MGS5(7dQC,#Y4B4?(PX/L8a@047EaKa
?U0HLNaEO#Q/2?/:Fa7,G94GbM.c,ZMM57Ag2VgPNL]AS(B:3]5DB;(QSQ(2VWQE
,2:#960cO#PS\b0P-=>[^\#H3GY0cgF1gJf>(?5RIF&B]d@ZFcREgH?W88Z#<O2e
D/]I._51Z=;(ED68:&5E,<S@?0,6:daO9)g[FQJ[g<2OE;JY55OEe]@L+T.DK+X8
:L)B;INg&K>C-R(6H?:X&_G\9212QW9_E,I=W-^c);D;>bXX)B],KZ>H5Q#,XZDX
U.C1QM+=cDOPJ^;X8UQAIc-GY)(.Rd1.][L3?/Hgda^^+^g&aba+AKWPQCE\S&b_
91@Lb4b,?D;BJ0HCM<JEZdZ\c]d#B3:AF&ed?H3<Dg?0ZgK=>5b.Zg<C5HB=IG>0
CEKUD;gCC+A,C]9>Z=?J2L^aQNQ>Y@&NMM-K6?@,9?K3S4(Qgd(8?.U&RP@PHIe2
PD1)BG4_0U2_7RWDK,Sd,\7ZK/Z;a:.1/S&&BdT.LT&278.UWgC[^7Na)aI;VdJ[
POD\01UFSTUAf4e)b/2:fQY[ZeR6VY]8dG=W^=M6F&1+8\=[[-Ya7&e6B55,M?;:
5N:Bec0JC-L=FT5?[(CN\a_d37KOE_<;\O-3gR6.6>c23RJeOZ9bSSP4ACOFggVN
+Ia8eDF>?PcAW,P(B<++3=J1:22Z11NIM&KeALP@HM4eAaC7:=MINA3=.a/D9B,?
EU:C7T6R]QKW4bN8X8)TGJB@@E_[.STW(,<95b&\XeDY^S6@^?>RCbLb.<U:+PZR
5b9CcG>;ePZZYWIHTF7O)9SVWE5Xg4&?5bg@8c@e5K\[882cOEdJ=+@a.,G&Cd;e
388<1]NJF1,JJId+GVJ-E59QE=<eDb^HOEH\f#PR6WT:[(S3VOb8.^9URG_^]9b\
3[fDfcM#N<K=CT94(7&\O^b-]1V,/J?G#9+7C;V;AS+3<,^44Q]3Q2NU2=g\1aa(
]bGb-]3D0Cb32=YTZ5Q3:N,1bLBN7,&.=O31>@.)FBZA=<<9bfFg)C0]9VK6gEJT
]f.K^UU68^bRQ8X&bR_B&G[0:d)[g=g1PLT@aEdOM58;7aO7Uf)U)O/:WZKYK/9d
A@3ZB\?3:7/eY8TV_^4ONK3XG>=d==U3/):fdee2VYSG\5FI&-\&bC+W]]IV_.VF
eI+XbYU<-V@/]-[NOW6Z5UFD.8DEGPQT>-a4J.-5bDbFf)e1bUX=6O0QJ8;0:[?(
?25K.V^EdJ[F5F:L_#2U2OJ=VH+U4g)1GV[4WCHfQF>.+-,#7e:;a68,@\/(U7(U
<KeeC=bAVT:>ZacIN9@:L8G#A1f@Lc]3I4P+FCDDRA@U[A0QE6,BZb3d.L6<X1eH
=358N.]?g/M8Rg@,8HZRb,\:=IgJKR4SHb+MO@UA<a+^)JBAWb5U.Za5fBg[O^ZY
.Z07TNO54Fg&JFb?2)D-5:[H(_)IS8fedT_=H/b7_#6M^aBV:?[61RP-Ob/C2AR)
XIKQ15R[Y>&dH>F0/,H#.8?DR#:))]a+(WP^10F.eB.C)HeI[Ed>cfM(XCSJ:K@7
JVg7b^+EfUfMCAB]MK.V-R,@f#^U0dMU:eC@?2W0@e@>gb5ODGA8&@aR95]X0(G>
g(JNaW\I#gWP0.#3[7C<@:\.3CVU:.2][??FD+A,aZMP?.XUL@567[0G&g[<45LL
+DOKBZ+dOF]-Tf^&<f+<D/&-_\]7HORZeOeJKP]#^?\42B=LbGbBY<a@PL=1UT1G
2#8X>c0,Q1N:SWTTMaV/Q0VE_Y8A\^fYX(_8#2cDBN58g?)\T&Kf^\S6U3Off,e6
=\:-<Ag?9S\S)D>ES(VfVeE/9BfS,g03ZOODE:F7]_6WY@4Uc5[LO;8QF?31[dA_
X(.M/+cI(e@\KVCD#>MI^M4@6GKP]7?()eG<2OG+M(cF^+N)83ML(fPYZYaRLN&.
\@7RG915(4g^(L,15OMHBM_9DVI>>PJ7T8JC[>N_@Ub7/V2;V]<AWZ[,<FC2O#cJ
H<WSMP>BYeMD<cPgRS[>90B@6/I:K]BG(JHfNI1?^4^V00JR?IR3\838?V^;-eRX
f\Ve2/eLe^f=T1ORVTVdPPOd8[.QS3)MCKeO=-)32^Y)ZaS<XVaa38#g0Wa(@R8T
[&G4XS9,YL[AZ4/(?=57]\(J9KcVbBO14OQG#USDM09AYZ<-;e201.J3^O;Fb9(@
dNgda/^7U0+1/IX=I/QM6a,=6N;/a&XIS=d(Y@d><OPR(?d4Y9GSg9.P(6ZHG(<@
D>dXbODYDB]ZX5.GT.B1_/+>VN553FU_eP)D+aLK88ZaD@TQ>)74IT+]S7G_CP\7
<F(7KZ>?82=Cc+PYA.J+4BJ)]SY#;@cY>bF)#YgegbY(A>d#6VSN&VP&9./+=Pbf
ZbMV\&LccYA;e]BLcV#_0SU:-_O0d[g9MR]?B68_U#:[DY<H?O=>,VG7FVPD08@;
VHCb+^;C-MQA&57c#<CY0F\ZK[W;ECLLDY8^P(Da,/T7LdP--d-9<>1G[=0?05B&
:f>AG]M2+A_A[eI+L/@U@^K\36RE^;OK>1;D&J;bBY<Z;@^>=1C/]f_TU;D^#AGI
c,V7((f6dS<2GZL8WB5HVf<)6<gdf?BV@@C/BcFBE;],=7REA1a&P:K:\EaL0Z=_
>+^O-H8<bHHe\PD=BM+E-<=GV\UT+g5;6@bT;L4J\#G&fY@72LW6<<[&.71e;H?D
^a4,U[T:\PQ^O+:fLdVW2Ke:(UG#&EB(]dKg:P2df=Q#dP\Ne><<K+F?H76Ia;]C
D:>8fEN-H6UI0_XCYHT/</Tg/FT_M2U.E&4GD-cU+V(\#N:;:fO1e?D6<0))/65_
P5>bN8UW)_918eI9@b&Z6P\BP&THW]8FP4;D58J8PaR_[AbP,2f,:QA.:AZBZ9fP
f-JfG@)<.:CVC8F&VD&+C42-FK6cTL1QK;[^LBbaTJ/7^&N7A.][=73K=KS-^C\-
H?Q]Z&e1([;<K#;#&5fN4eWMR.1NQ=[,>e6H:PRVI,K8-B)?f_/0AWL<8C-0Yb<f
^O#WZ]8L5Ha_7dWNG3X]/A_B^)c?MP#6eF4XfXY<#?a^BLEVf,KR-8d-8\#UXbXG
3R1P]Q\X:\Y&KQKE)JN:CCWg12PfYS;eSV7IPNIKe.1R<0bT_=&--2Fg4g_+dU>[
4be(=cUJ[dea]&6,4]L+8U1+=TfY>a\PaP[1IQ-MKVT.=H<C.,<G.F,?<^517dFQ
MeX)J-31-E-gcE-HaIT-8e7P-@2P@Z-f-?cbC[+JB6_gEbTBa2G]R<9M#;SME3(3
8IdZ]EH[R>4))bCBDf-.AU;9LgTg\5Vd^;e8E2I]X40WQ+7I<=bL+&^,SHH^]aHL
MBR[e]/\NFF70A;M&OCGN>YHbS]QR\cHAW-+&[?3?cc/J,3)FW+,C5[>\=b1]&1R
gKdS2-.Q-C.DE8@4bCgGbOY,R8K87d7\O#M?(g0VcR_0K;DKI&W#=FQV9:WBVW/]
+BRE28P(C;#-I&E4Y995Za+&V2R_F0W_42RL#\Fdf[BMS[CC7-;49,3.;XF^LTMd
e=KVUaRd2HU,+=O_f?]E,:&SK4e#RAd<[8NG3XA23BU\FJIV-3bQH>1f?cQRJ7IK
1M>NJJL_4eI#ePB:^<XUW#RQD8KW^)@-BbVCBTFJ7PM-I8(918,HQWbZ9K?(P#,V
e(,e^\aNEWOF<H(5(Q1(OTB?)5K61,<gb<O42;R:Q9W/B+Tgb+ZgYb>78XL&98d4
VL4/Q<V[IOP+1YJ<Ie,5:Ca/6XG^9V)cX)J95([:VcAZGb4-QMVa?d9VSRd+@YQ,
K)^I>D&A^.E1;@C>aJY8NV_2S=5>]343EE\NBPTf2G@bA=LNTB;MPRZ[7bGL\S[J
5S#96H8_)Z6/Y;<G\6fbW/Z/842Lde:8BT?0D.93CPOe-fNR)#J_.[Ad4I2F)2O@
H?D8/,RTQ,WbN+E8e@Y32Ab5/A5OH8gM,eeU82(\GB;=-RJ,--Z#IFbNSdAaSK4)
B4Pf-+EFX3ac]bdCW<g#569-IA-XaB3Q.aA#?8LDMR8:WOZS;bR=/+UU)\#5BdYV
WeI^,_bG,0<(>F.+3X@B0[GW&\NPI;BfGU)ER#67^5H._@,5-\C.R7PHMX=a5@-J
O;9EV]<EgeNA0CMC5[@?E_d[8QKYX4)a(B:(MaIKOA?UH;\G/Dg#1c#KO@Ifab-\
4ARLD_b>O=DCfbe-SK@_+WfIK.Z^Q5LXeQZX^a+EfJE/9c+3TN8UO#3I@eUEUB8:
/27IYT/d=B4Y+(/Z=>?\JE1[gLf7HBY2#24_F10M?C/&3(?,(NO:->0HB.@@L/3A
I-+;EDdZc1.\_gB^;EBEQK][RC<KecPKNc(E#=[#?0?KWcUIZ)UXT,B-))g]#4\<
WL>QfA+)H2ET/bF967.V(K2-Q-^B.b9H/)_CP6ED47#E>F^<1&TP0=7AQ_]K[.c)
?@\KQW2aVBE?P,N8AAEcBPEHZM+H7EC3DM4XE(&6F\c9_G&>dZ5FI@3M4&EG2L2)
MUX4cYR4M.d^9FcF@GWCMP3(Vg8B=EEeG:/2#Q,g)ANFHaJ;,gUPPS8aDJ1VTBM=
01N4&I7=_^1KDf8T\/@>>G1X[Ud\d<_?ZV0;.#bSZb@cRLVVOEJ:@+8edKE^?bIE
5TE5S-NS[X+F,JB:c]5I5=;-_PPf9NJJA486C;&J8Q4c>7B3Y5eKB/CPad#(U;;b
5g1D0QA]I_(V\2LG\A&#(64]Y:3KX10?(G3)>,T?YdbZ;NB3MLP]RK3;TM6Y\\D=
/9KTE7GQ<A+A/9I?]WeN5;3U1H5L6@9O4<O>[[[014e12B+50XDI<8=R-2]/U,,>
THbbK&dK,6<b&77/<TGG>DR&?/@?dM<VAc[:+2^Af/WHD3b_(2e7=^X/2A9a,fXH
1bDMQQfYG4^G6NfV_&7AQY=IDR?M&#S+O6b^#J5?;7XF5[fc:6/\F3@E4&]34d\S
#HCb+21S5#?e_V+&UK.F(5S^6Ha.&Q2IYQCGEGDV1Xa)?]AeJbEg-\O2.>Q>T)VN
_]gJ2?O@X#8DG9G0Nc&bOaLV7\.ZD>0@J9AJRaZ/Z&=.=ITGH?<c3WU:B?1Tba5E
(,?]ECeRFGVO/EB^H_)/J9B?Jg89@a+K)69>/X1)EP?Y8BAO[@6GaV?JRHdL8;1#
QCWRE#^7e7JKYJ,S,D\>@HZFB6b.3ZH-WMW)4=JRIO6#c2P&ga75eKJQ=IE.9GD;
5JRQe?KKW&[.0fce(&+HdPa(5YU]T3=-b9/QKUV2:@W1Z?A6aTK^A2Y=YAb&eE2=
g&(,\A2.11[9SYeXRI>QX;8]^/OCI1.)2CW<YGRMGF[-QAS#04KMdA](M;&98DVV
HR1fO>;Wb\+,MV?&B\W2@.cK)E^8>eGKO-)#0XA)/#NIG2+a^5?;4eI7O4f8ZS^=
E(&S[TG;GI;D&,Y302D.Y\&LB)42PN93)/\9F[<DF9E-;d,_9E;@-b??0D/<?=3^
5OdG,/.><6dHH71&)UO6CHATB3NXYQgG>0G<??##c#e0P/+ZA1OKe.[:O>O-fAAB
K;EUQF&9B@/(E#RI[OJL^#Pc-?1JWg5[Z&_=I=4aOK[BQf[M.)+7WE2H)f:R2<XS
7#(Y#ASS6@:@0XN[^I_B:W^aN[:+f3\XUWGaWGJ.4>_MR0719(Z\F_P_^9.\P(E<
U;UTaPC^:KX9ZWC]DP.ga#Eg:.?FGd/D)504O57@Qc)]G-GCR/ILA7=BF=]KYY5D
\fKZC11\#IL.<UbPB[2ZIdVT?0LWWT60f4?&JAa@D]d&\=+JB0+16^/dD=\O[N4Q
_6/>&8DX>_fODA>]E-QOO(Fac8CbbU7Lb:/7\SK#:P2UDM5RP76NC2WZLD<fb[#+
0BOf4?JeZeYBC+<H(>-/ED:C><-XDD0YIc(0]^0fZ)3a/a[:)a/]A58)7D/2ESZ6
7=AD-,]\9@fCQYK\g6Z:#gQI/RP9SA>Ncd8XQW)BXg(/,;49^LKF&^VbR8QH^7,\
3B-1H,S(XFE(WBOb5TJOX@H?[).5?3<c59):L?TG3C0(VHN&DaYRVYAZMdc26&8)
e3C?X>V&HgG3A?KL#T4gN6&MW&D)JX0d)DP;^g[^+gH0KC?1N,]J<TPJFXK4MOH\
)[3WI,P]/82WaWWB>Q36K\/C1PU673U[GJA<J#?TV4-5,>+W6+]KG#XeccNA6e0<
Xg:2d>\bXQL03Xc<S.QCS._Z,KW?EJ);G<M1@Ne6]&8f=5ab[;NM_fLL8]AN3F(5
6c_[OUQR8RIa2Rg=0QJcSeH0L0C#FL==CICf?.ZAbF(A(=YMZ^^VQT0S,L(NB2BZ
X0M6O\5.V,@>>^+W0@,D6]P8?M/<32C-cRO\SG=6N:]E]?Q:2GPS8EHc^0Ig1)]+
99;CFV4E/>gUKPGUUJ77J&WI6GUZa<Fc\=01MC&Y-303W@eGR2+YB.)Y2HFQV]fD
_P/-&0GV.dE/S6\YH]:Q)#D5@#^.#L<JXH^LCF9Y1WJV1[TVg&Q\P(e7CXTLV<9d
/26>bcL?VNJc6c9^VK(:#@TKF9CJb7_#TS;U4)DdJ]bX1G(;\N/BOA[H5^bc/HLV
([1cJ2)De&N=_4K]S370;gTfZcT0J^E1Y&a),TC50UG<g/2M]AF_;-7MRc]?d##J
QZG3),)PR1/HEB#PcI4(N+fg#U@F3V?B-([6=_6gbQ:>Zb8.S,8ZR:4Z_;gG_d:?
KK[R@ge2gQ?[?&BMeXI;,>Q\P2_U2GKXeBX::F8.O5]N./9&/P5<IJ)W.\J[6@FI
9])DTTF>.gE?TJU09Pf\Me=VeN=Dg_-R;H04d+T33g=FLW]GTOg;Na@(#@^(3RBV
Z#@GC#0+4d6RBJ40g55cI1,Z-197+cb5^>SWC&cc.UeYO&_39gbQC^L0/]SND&?>
e1M:JDd.E5[/B)G#RI1^(T<C6-F<<DY/2C0U&&\K7500(D#GL(WPaCJ4W2B:^8;F
LbO3Z##UFV(bF;E[M;T2?d,1H^,b>M\;N9;-Q(WSE]I.C+Td7fIGZ/29SbLN#fM;
M1c^7D1W+Y1^f[Wb?\;Ve68INPIX>VTJ:XDa/H9KCK:@8S:2[EP5gY\c\<+8UIIK
OUP2\_EGQ);Sc93fO-SOURT5,-BcJ,N4H3_P.[Ld?RF>RdJ6.E.b.f/)/7V?.?_U
WI3L\L1PR2R5DJSSbf?c15bcMO)25IL,3R8X0N[-&ZM72d#8J.ABgS3>VD.+UJ2Y
HW)-:<g^c),B8FUMZL:@)025e+GTIH(E[V-XGT(QO<E?E>aY#^OMgeZ.N=^-YcD/
gM91X1cB<aY0)H,K7Uf;HMf@Y#O((3D:W?5)[CN;VA0R-Y&S;E:a&g+)@BEEAI=O
UT21]9>A715FU?48.6]70UfOKB](#87O0fL.HZ)8)@9?@[@aOF[S:G29ad(dR/-K
XM3KPb)R6F<f50T&<-g7O[9ePSQ;6YBP;(:_bI+E.=NP7KLHaR)J(O9.F/;XG@6.
Da@-f.RcM0?J[Ne^ZB69M-OS[M_7;>(-f\aZ:a(cVbWDfEb<#F/b\-30K/MgU@_,
Xa4/VNRFI25-dUXTANB7S[[;&;>,?YB[QV5K9^:\5)_?D7g#HaAPFH=A[#6Eb>].
FS3M-:C<[7EfJ_NUP2e5J/:J7\4].IM,d#=cSFB1)#-3J5O,UU=a]+,g:O)U2fB=
IR;4JVg4,e^B;^^?BKLe<#Z^QQCX560a6,BdA9UZ9XL60R0V,XN=@Y,F/?GeD6Y-
B=F1[YE),5R39PA4V=I4Q,D@g>^Y/a7\7\Gb0K0Ra9c[b<L.(0cM9BS8374-K\O6
7ceaLQ56DQ/[G>A9EI(@fcYS/[M8(U\--g=XX0XNA.\:T]f7C,BG&61G)W)-I89L
RB5LG0P8=]9OZBHfS8\aV2IXb/]IFUJU)]4O()/DAI3.<DVANS?</M8OGE72MT^f
UKYWWUW]8YECfbI:cNBe+bDNTK,T.VD/1FSA<C>WVR+B1EFC@Nd,GAY(MS4)Sf_L
[S:ZSHHMJ(V=/C/f8dG-C-QR;E^_f^^0.3+b9Y5.8Ye6a\\8[_KCeY=\b0F7e,UX
A]8X;&(44+?^c01>1G1Qf);(0A->&QaAAML2&3dHFd>\GDCKAX5XN21;b<UD+,3=
FMSeRJ)\b0MJ-.:Y>[7@4/M\;A4USZ9(c?XO;+0:<H4PJ-d#d(SSRR)>J.6QCV[V
JfQ#UC?11:=;=Y/AZcU7dabfFE7cP_/YOM9&FWbOf_G&?FHF^AJdZ0XS?2[3DA3e
O74&/P8(XQ,U-V0G57FT0-6WN4&>HK.1N78gK6-9MJ8eb#Q6-BMT8S6P):Fg(E0_
Kf344#7RPO(P(P[b8P9F]<UQ_Q(DAR5.GR5E([M3AA>CU#<;<X)-U57[MNO90>,H
3(G&4WUK1I]Yc6QVI77af@]2]R6F[)MC:3(2N29H\Hf(IFWda^PU,2-c9HeZ5E#X
48Pc[>)BM0cB93)::\G1gP:I];YPI-8^YgTKd,Ag#MZ?<Ugd1g/9[dYC,]:(b_@<
0P[HTR54F8VYR00R&E,adYKR@>JX]@QBJ74)(Dg>IPHfd#;f2-C#=6;+\^I_CU(Y
dUI0T;XVNVA7A??+/DB7=S(FaL)JD6I^PcXD7<<d@+XdEA?[gG&:\[NW#OBeGDM-
aX&<933]-RH_LHPM2Ib\cWGXS;Zb/^BaIH/NQ:?TM?]L7g7(#C_]LA]2QHc8V5[R
FT&d/&]4OJYJBPa,ATgHVN?<CTSaEDZJ87BI?f>K(9PD5>bc4_]^HD5)X#;K<-5+
C+G;-P^@BVLd,MCDML(53UA)=KNT67L(LV25+(K30A-1NOC_KSRR7:cN8RDU7N2.
Ea+c5O_NB0<1c&C\H6#\\1^,-\N[<2TO4)Q]g7M9Qc9(H:/VLPa_<RZV#FHE9Z)Y
XD^X7=cPaA#e>:O,7c-gP8#]A]ZQ(--ZWHN8S3(/Ke=DV)a?O^T<1S<W3W9PHM)+
Z.c^^M.VaJSU7G\4;f[T;[25e:A,NQ&F^ZTcH@T>7E^JKF6FU3Y]6[JM,8aA,Vc;
37V5fZ;V74OVVDBdE/5IJ=a8J.cbN#RbMe<.363^H>MNUL3XC<UQW8O1+4ga2G#\
cH1)D]SP,_>7LM>VS9MCOc;6#0DQ)_<O-DbM._;I_A?7\27(XBL),YgK&(L?DB_X
Y;CLZ7IQ\VD\YB#QF2G76L7&gRCKDI0TO>ETMg:;f:#4@=??7QfV^M]7a8^DRC8Y
DL;PTa)Z[>,-]_BW-CFY@6DW-<+G9PN=X8ON5W<0NR^EH.DbIcbR9_GK#>:6C._Q
,WN)VQS?IAgP5ST2442BL(3M4Edee>?eQ+OG]Ra_GR4(?=e3PSO=[ZdIW8;Pe0Y&
Ac]G-JCM<[:fAV?EXb;e??W;MAL/:917MH4/>F[</]M9JPOJX5TZD#TK@=@51)]>
^^I0g]OOC3JR&R7U/H,/bRA(&[2(5W3]PCVP0F==Bd]?Y^4I28b+/)NNMRP;SB6U
,E62VGZ>+gI5BGF5c,E1KQL7cSSL]CK=SLFHM4[8>Y)ae]59Ba5[AR;_eTgLAC4g
-0eQSEN<^5HV&K&_HS1S3dPEKS],Hb31XO=CfdL5F1)_4W_bR&B\^.e2KAJ)YV_2
@=Ca9b)Qg7(TDCD7:5?H?+-7&[+.Q)4bPF.EX-1JL55C1&I]Q1.:WA8cP#SK+BI<
Q,9PU6W_46P7^:G>J?0gT6e(aEQaX:OH3EZBWHP^OMW#U8T^LbHa].@L^aKXgf#3
7SL[]WFAIa^OZ1V<HJ(OEb2WIId3H:&NaBd<D=6@GdD9@318<.T[J9dD65KC0R;/
PY_(c1?E<?4YF0Ff_b_E0SWH62<D\/L@Y?GW&V.=e#H(Q?ReAcIQ4c81RKJg-S-4
fKE7c2(2U+K[3gVY#X#7DeOS9)>bC8b1+KDfA,4<Eb.1PSAU\\VO[#10Y&NW^38[
+e]]EHC4C6/.+99b2D>e-S]#.8E-HVXeAQRfbXRLBCL[6C&WD(:69a]CF.bY\+_E
&aVZU0)A;00DRT6GC?_=PMe6e:<&</dNgV6TZL6JC@(6K&=Q[@eUGBZ1;)-_:]e0
C;@LM4=g94@eD-B4).fDBAH=K[K&=RR^J?6T8RK_=JZD;^fH;_fg00_J0?IaC<;^
U[+(AaXUJO/::VBB7a,N:4<>dL^^93cP6,f:)FXE)b8AI:IW09OReF[8-0^J,000
N_\NYLafL/87?(-b&Nd[W\XJQC3\fO5GXFK1-\eaCVJ+a<3g>GK32-AQ_^f)?R@>
SD>0\gHH0(G-.#AfM@@7HKDB:NRJ3UWKAgOUBFB/@aHAe^C<.AXVZ;K9If;UY^Y+
QcfXYUXX9-N+29S#GQ]D,10URE=<)gO&OIJ>e3PO=XfTc^SGb9<2+@6X?YC@[V;Y
B#aGJb^<;\+CYM&>ef+(C;OAP8O_&M0]B6:0&-.-<^=2b1bKQ?]+N,CLN/9#7UeO
.L-CRALLfZ=ONRZdc0?Q.<5dbZY(?)eF]0^6VYP>)++H7ZSS.2_#.GZ9&K8MaAU0
BY_^1R<ZG&V/e8,-Z487/MU3,-MBHY,D#YQ/JaO6&\CfF<,Jf:HSO0LEOR+.33PQ
1@+P&,2S9[PZM0RY,HTPK5DNN0/@+.A1BSY8;3GA@Y0G/[G6/>c[^\-efBg5]L7G
=^C1V^QFTZA1a56\K8C:[3f_3V4[<IIB#:7#5b3a4M4AA54@-d^8ON^D>A:HJ4]F
>:NS<a>Vc>_2K@T26:\b7&:dHS)gb:+-e_?,[Y[[A\A/>3,Yg>]^\=<9da.TOY78
f15,;BWO-/.b&f0G?BB)H86,cN,WFZB^5FP)^VVN#V7]AR/GLXBSI4/;Z?#cE?+V
H9-/;7UGWJdNVCW\Jae7ca67,#+>#[OS0:4.4Q+\g\:CHB[7AHS>7@[<>e4M=;<C
D/gJLYbHCR&bK<63<L71ICT.)MG?HQ3O8?GJdGcT./YI8bH1IYKDN\^G8JP<X^7#
;EbAQZ,+HB,afa_7PYI>0-Mga;P47PN/.7A1#EXJK40+Q=L\8#AGcK^IQVB92Xgf
&V-2B[.f5ITG4@_9DRXM(.[1/.P\R6TeWO]1#.I.0d5#^U,=:N2Z+<d,])c=VO2P
aVK5fSb7F9;;HMd:X#gXU;f[L^TH3FUU[E)e?39O?R_FbO6A3HUF@GB#/L(,?f@6
]=IZN.e4@f]-><KFSSUBC()]=NQd=EM_BVC7DHZA)_OIMc/HJaTT77bX(<5>A/7O
Tc(P?40Y+gICOUVA@Z7<LcGf.Q46<-6e1@/Z#T9Q0+Z;MS^/,\--^+NfEa<7BX+\
G>^5aT=8Ca0CVa_Q1T1;5VPK1eWa;V^&KDJ1@+HD.AUaW,4V(,^R?9X<(O+OVDNa
($
`endprotected


// -----------------------------------------------------------------------------
`protected
_X4BCH7Ob2TdZ\K\+S\9a0/2A957R7<Fc0@1F2c66Ce8P?];U?94.)W-J\BaU.J(
XM)4E8eC.D9d*$
`endprotected

//vcs_lic_vip_protect
  `protected
,ERgQY>bIQ+_/-;ZU;Uc@+WWf;[R4^\ARbQZbZW<5[8(7MI6+FE0/(CJe.U89&Yg
4#V^DB:@]7L.1B#45X4RYE8YA/;=UBJ<DE[c0bU#1>R,@G\B1XT\]UO?6H(VXG&W
>((T@^YN?[N&Vfgf#(K&IFdC@RfC^:BP)PNDX)<a)ZS76@6FBTMdbL42AO:G)A3Q
<:\UZ#)FI-gGdHS3?^,fH5e(5EAO#S(d>b4:+Z77>NXD;)a7U5-)8@2H(0Z@ZH3g
D/\d,SU<FaU5B3;JgP2O84e(1$
`endprotected
  
    `protected
#:+Ga^0O.\c7\LNgX#@e1g=@F-ZVD=.2Q_5_.06OO.YfFCLO#P[b4)Uc-UM:AQKN
GHP756W-.fI1Z_g0#&VdgaRBTV>>Q(0-LfFX4Y\<M@I+2GJ7d8g;1Qd#TW4LNC9P
YR[[41?15A=dD<-H6VK67XRB1$
`endprotected

    //vcs_lic_vip_protect
      `protected
?/R[5SRb#:]SeVba(=)_Nga5.JA>\^0+5Y\OV+E1:Pc-[@,4_.d:,(YCP&.CN#-<
++G(;1agL9+A5LE?#PFg6PB-]4D>[@-+E=L>bJPZd6a5BT_P-&M<UHKA<<DGI=O5
B,Pe(5]Z;dd=JY-26[2O,c\d=P(/N;58#\+OCR@@T?&Q>JY@4]-5Cc)BcOG/]7ce
.7AYCOdLO9O<\CQb[eA:\C0X)00a;O7-\8,@)B5eY8#]NeVKBA,UTLGY^&^#[G=c
41f97SGZSHc5;.(#5/R:Ua]\>7g#MLJV=G\@XT),O;I=R.LZe]cV1N#b1#P\,HMQ
P77:)\bO<U1eXSVE1eD#.8fV9?A8gO?V@P^Q\a10C.F4EISQT#P9J4,f4gLJ:cAe
JZ[,99a)VXf:Ed4DZ(Z38PIPd2AO(W?#;9A05A@@2LX#g:^_,b>N?<O_U5Q[LaQ]
?IH9)g\d;+L(&B&OYW#7XDe)a?M;?fVKZ^eU2,J/A,M&&PKOU)>6bA=VHH6NYd30
^R)gB1LKe7H/I;44=XVgf<GIBKO</,U@_\4Yg20cR\+)\X4B=ZV^?N0XH:(c3XZF
N,#ZdM1B;,9eH>6bgI,X5aLU.f:?]O_WH81\##&L<+IKG@4P..><+O2Q?fc7[WGN
=#Cc&=T)E7SO0)H=L7LOd]FE:-3-;S@g3cT^#,d;XQ=UKPW@a=Zc0#TP5fPO&)Sa
^1FP@X,>&TNR8cVdF5>-^_T4/JAJ&^(_[geTeMfVb@0X4TFK,9Y?POW&7<+[>bV7
g8b:.:JfGEC]cOCVReY6WMW]T?+9DSYZ@BW7]TT18LZ3LeIYU_;QWWNbPf_,R&EC
B0d_LC6g3>?cOZ92e+Sc@d]bcDZeVY1=&3G8D+\5@<fU,[]K6fEIZZ_B)O-B+]EH
Y&&J1M:d<,agbeHEK.U(TSYJ?bCYcNG/F7T6TD)YbN?1N;#GE5T[3#aCW[9@Z3DE
e^aNTXfO4]Na;?6_4=3A-?[0.W#PeQ]A>1YN1_]E[NP6=&P>1GU01X0PCKLZ]W(Q
eN-PQ7dGW)ETPWaGNCYf:EV_4;W5D51ILEYE,N>c@--M0:2QId#J;NFKa8AR/N^K
dbOA712c_P?@[4cX47>LG>YM.4K9e=N)-H(9I?<O2=PdJ+O/=A&^E[XX<],3QNc/
7&aMAP5^T1H:95?@R<f;Fb)Y@1^?)0>5f?M9X;T^ZM<K4V4TV@6A)2<ggd6WQ1cf
XR_H1N:]KAbCJ&QWeC5ZU->>NMN(XQ<0326C)Qa_QA(,([7CFA52RWPMIS=<d218
-fJ@PR_76=86BWg[M,-d(2445XBY29+[X<N;XPEP/OI+;4G+-:AIU;MePTf/LM3A
4RW-&W[eY7_)c-OV5W1aRR>eBFFD5B-BXUZKP#6X6D5><0Y6aE0JRXX-c,>JE2-g
Pa0Cc)@>e5#/2E+/)U85c/.c/WJ=RD;5^dQ[.<4R^Z)6IV0BFZ&..KYGG4D5C#+:
=FdfP5EVDK+F/77N78)OE\,I2CVg[b\1)HI3-^B1X5,@7X,#IIgYII:I\A,RK@QK
][e,&b@_?eN8)V_3P-+UYffe=5<&>:Y2P4&4XR1a;/[:\RT+fbf5/-S,cgGgaaGV
(<PXg:-JKPNHS&+AfO<X@_Z9D7fVQ7?K.4_HA,(5@2VEP1?:W,Vb_LP2@(TCf<a0
+2AaQ6&I3FK)LSb0QFR\gLWXPRWKg]b&VM=dW3cPY#/QS?^)e4:U#V\M7(K?E:b^
]d14Q^YNS@edWN_-?D[X#fY0;g.2egdF8/K#B#C4W_7dD5DSC,/O0=WS;O<J1CGd
9)JOUH41S)W8)52^,0I_\AfANZH9_-RbDN>?a4U6&:Cbc_MNUCcDSUc8d9UE(QQd
H[@FEUIO]c]C/:8M[a&3(+X#2>8aG]SS.OeS(&A6UW9;ZaBM#d,aa=)HBeU&VIQd
6@Cg/SFLO-2ZBZVY0T/WdgIJ9,9-VXPbM+E05U8/_1H&27bRADf^dfRW\O0LR?VL
[fAK#LP8RMeV=SJMVQ24N5)F[82XObRX<\E4J;(MPK[0(70JQcE0a)2Wg[(_P.3L
,L#\;SHa_(-gX/X]cR,(0G^1Y6=5((:UTEV/>N,4gH28,e^1.cV.Ngf3UXV7NTXa
LU&4dE)+;g582DeM@YcNUf^YOUZ>g0OGgDfFM(+cKcA=4a8b/0Q)RCR^LZQE5@@e
M84C0I]AggP&NN#[C25C_aJDd=GN,Jc09)5.dME0b?f[2^YB/Ta?;@dMMA4<YGbE
V>[;@-LSa/#[-6C6b)M-BRH8W80a7a>BNH/D(@JJ8KNY6MI9=G;3K/d0<fGKL;#J
b,B5HK7/74dM[,[6E3]Rb7RA\TD1]]/77(Y.5-<Cc]GN-1-XZ3<&I\E\6F@Tae^I
4(KWd<-W6W8DQ6P;;?.0_&:G)&):NTODBQA[II]<&BP9[Q?.+.f5+a0[9>IdD9Re
99QI+HT@ZXNeg0=#,Jg?D#POP0?[Q0/I4fE=ZgO/[D,f74eb\CbE5]U2Y2.c##Q>
9H8O]c^9\H;9a)g2aOTVZ><(2QW2IK16@1AKb._[-5T)7=_d@S#U\4+=NBR=#DXX
(MKdZ4V7K9@8GO0#\XMaEN=2ASSE(8\=&HcB]:]NTT\FVZKgO(,7E\#3f(-Vb)W-
HE&[)Qe8Y[YUaP1d0;O^X:@>JX:NB)eXYTM<419XLRD[dGYF0+KWOU)7YN>=#^&/
/R^/<cUAQZ)>QO,8QXR^+QIT#FMA:;-?A@S]ZTB1WZ1S(LPRZeeWUTef4AVJZ^V_
f6H3\XFT84bGc36XE<dAa,GS11a=JB+XTcN<\a+/?H7K-\b)C-/NVJ@J4HQg0MKT
BPF1?.-Z?ZgLAC,_H.P3EODXPRb+U+;X:AJM>fRe8>HT>5fXW\8A;?ABd;f0;/:3
7<4,(Z1,C<]PK8T?I74\9YcB1gBYVX\E+[<:=/QdbJQ=g>\YQF)eO@07I8b&J5A]
c7g:F+_R#K>DJ62?8@N3^cICVMU;F:]0&XR=2\W15&^NG/<5ZZIL2R\e^IeU;\#?
L6Y-e9D<?CcAL4]+US?(W4XUeOb)0XAGIe_X0Fa?SeW4C@::C@2KM<f>XCASaDf-
UU]?4D2\[T/d_BNJHI9c+VVFDJI4gBT:McNB5V\?J<8K@B,0I]]@X<YbM&bBaZ9G
PKd.RT7.ZMAQ1?TQ[Pg7_8K]_UHeXCM1=6R4)H#T\A<N0e5,HceT]K1F-Z#[FLR3
A+:Mf)ZD_.7W[L<@b?Y>G(5)B.S0]I4b-g:3K\&DfUbJ:Lf4@Rg#B)J^[],TCNaX
0D?X.:54)Jg4)501dM0BJd?FT>e3(=bcHWJX5a:bD,NM@:T@N6fLMH/W_OeNZ?2e
DP8=aL86G=OcTGb4\05@MPTKcSb0\TgP1X@^\^R?E(bGW[&S(B^@T_D94fM_FAIC
1OW<=TaVE,/+&XR:>G(>9N/^3DYCA9WM)0;bd5+X:[;43Og)AF0)e:/U35[S5K5R
;?\P&&;=K?>R&HbA-48A_R2VJRX-W6&S&gR>Q9:#V^?+VOd+<2^F;-A>ZHcQHd1D
+C5[2e\QQ2>@Kd[ZWE0H5L-J\L6eLdKfYV6[&33cIH:NC37\ACSA-I21/_V:IY78
.K/54E-;JAM@6DI+U4#&b(dXMEWb(d2g+,IGB+I>.f?7Ha;Ef9,IBG1BQb]cB_KS
a3]:<^F)HAT5cK^,/8.TY5EP7H6\0U-Y1L[Y^gBSLY,AT<a6+c#,@:dB;Z,^=8.b
f<167>5c#<\=7Y==,>BH2]cBHLK_g&QLc\#dG9-V5+J?J0&QIR-/A9Q)BL5#2da^
gUS\?1N<1OP+78PJ^4YMeN]bT5BS@,1.RQ_Z[c_4_@0V4]SB<DB:V5H7+<@&7R+Z
>RGR-_?)M<(gMS\LD&Xc9d-77=66GaJ6E_XQCOCIge,/0=W_[U(NU&GAaS)SG23W
BQ\3S:OJ^5J:[>S6@<eCW_3S2-^MJ^,?[C^8eHXX<J9R<HG=P-&TYLNL73a9PZE4
XG_^E_3\P<(\-E9/(DPfP7)@P2;54D_Nd9ed/VVM?I&3bQEQ5>XfMRI+\ZT?fX_V
T=3g[EcQM=ea5f;96VO(D0YE-X8.1SC?D1(E867II(D[fZ5I9(Wg-dW];)D@DDDV
Kf)V\RKJ0^eB3KS;4CKID\Z5;L#dTO)=MINPTC79HE\BW#5eaQZPdHb:RSaXO-g2
NBcgGPQ5gC529bXc(3:@T3C+S:_Gd6ERLW3^[RB1Z:PbegOL_BIYI#[Kc<OO+W/c
#,)g.FMJTN<?>J[/V(I,E7WOE<0<_&b_IA5dG8QbNB[1CfNP7GKb&U_X7-]LFR\[
V5WM;2b]=gM=Sd4c:E:[5V3<X@5;c[^c#:VG]B#4g5RHQ2aT_&)3<Aa,GG7_.Z@H
5A8#L7aOIJC.BNF:c3-NR/>97Q^,d.0LE>9NJ+QN0]H0OVB[I-(&F+Z(4Gc_;Z?1
::0d/@f:8(DbXEG]+CU(/cdT+Q&#F,QTWG&J-AJE&EL7)^AVB&#8MSbPe=[6<TBQ
+7+1IG=NdQRJ97ATGg>PX0I^-JV,PY3<IQ01>KP/_d##-(K;EK?CF2=F9[FT.YNW
+H21U?Y[\4F^4<[0[UX_AN5?20UJ[fM(f#8e5+@OJL](?[D?>1SY]MegSC:6QT4B
/LB=2]deZU?78OYK?>c=,(a67fA&OT2?7H+C8NbQbZ0c@Qa31-aHOE3\Dbc5G\c5
8=EV-#9K>32EHO_JX<#9&FU9;M3dg)G)/Y5Y+dV#2a=\BYb1C39S+]ZC>X+K_L,C
c+\VVXJ)6G_Ld4c6XF#df,;I=M&eLU_aObIaMe)7Z4eZU^eO-526G+VB0f5:JX=]
WYcd[[=^(Xg4@2;@7<KZaJUVZ-2160^WQB7FgMKg3R@=a7;RGe?M.+BfA:+J+NI<
NY_I[\1>fPXM&8)9[.N]K7aJ1<2egD>8>c0QPHM.;/B+C]aZdM,4UESP22a+&34X
d]Va&aMINI[^3ecGXKfDBeF5B7[0(\eM,N&TFG)EZb//_BcBcJ.&:Ca6+;C^bTJ3
Q/)LH,.8&79R7DJ8f]EL;g-#H_g9>77(^?cF(IcZ[G29J6.-,OPH6C&/fYcQWC&O
?UE\?WbH;0R[S5&Jf/?0Z5a8@2Z2_&OD)#a.0EW=<V&cW9398]eb-edYIMff@f(:
bA-JJd#7RG)6A9R4;f@<<TY<g=Ca061;Ie0<B/G(TN?9Rb\F#6JaZLg<2RG:/XL?
,:,J8NZ&58ZBZLgbgScc?&:SNGR)HHe.&7c]XV7_Z67ECCM3Y]6@=cB^,;eL7IX_
.IVEJ@7^/(:W=LBfaXM9;dMO[ecA^]RE76,fC?^+Z_K:(U\DL^[&;IFVMg<]fTc&
2MQIOX?X=_F=:8D0:g8a=>X_[:N4)b@bX2>Z?d/^3FYBGgT;U(O3X>V]W)>F;78S
cE(()^@2MJg7gDeQK;(],N;5a_<^LKAQP_3/0;:^8\=[?,M1C[26BY&CM:&J5<e+
RN^5gEEZ-00DK6T/?7C,d7c#),[38B)9&4?7FZ[7\_^e\732=FT8:R.@3+]/[B,b
a@?/d)9GSYT56:E5GWB5a1DY80]<?H/AV-f49W^SK[LI<BQEV>[=[S;7^_GK,0c?
809:fE8HAf;MNg]9/\]<X9=e4[F^2d4d\.1+0&d1S6FG=JJ@aEZ/;BCRMKP.^+3g
B<8Sc<QdI_aS:@4^CG=V30A(F[_[Jc7a,HISGF3[S4U#6)\d>JO3,]TfF[O/4.JQ
<6AK#JXAC#4<aHDRX9d\?.Ng,AIT@]aL#ecRa7M1539D7V/<0&G>?]O&f@K/QLcS
T_9CD+<BZI[&MeMM5X&H.Rda[+NVVa]3Z+3TVG649d]K2LdKFYJ=+EdA/6/&::QM
a#A@EM0NX[:UXXSJL34aAP4Q@2#O-XR<2O>D_].X2<>+9L#1?)XW_?+LD_aR6aHg
93GVJ64F6CIIbTH4.Ub(+-Y=C+HQFGQ21>0f94EYE/-(]b_S)]fF+d(Q\/=,bPBc
SS#0PVXF[UH-,]Sgc6<^[FcEF5B&+T/5L5eIaA[c_7O(-B)L=OD:6+,;_XC=,9ag
dHbH<0W4]0MNJPL[HG?bQ0Oa70V@<ObG7HB_e;LH.>&WDNScU4U7,>UfG[TBcF2)
3FPecSCE,S<7:9PF3f>&.48Sb;9.;Q,bLAFFO>f)<,fF>?D6J@A<_L9)R-);eXG4
S<S6A8TNN#:LC?YERZ9DTB2S7<Y]+,.5<0D\/:TY,LP@40-#+2=W[MD9Ua)aR?AM
6,1_eRR#CRH;AM6#BO[4&Q<?Q7>FP^A.+5&88#KB246PQUGR[HCVF/W#<g4:@FW(
<,H;CP3<06dA&\D:3B=\/M-NPcNAbdAc=9@]-?IB=2<](L]2N^19_H;4L]J@ad8f
.57^>YJ.>P#b4&E1;&C>1bC,UC(4g+)1ZCQ5^T=NM&ROBM2)HdZ4+.M6S&dC70b5
]Zg9d?.:Xb@X5G&.0)N1&<9I[<K[S7;,DY#-UNXa3-aA@5;@7G3G,Tg\[e+V=X_2
eNbbQ[<f1(f08V66DYP[P0SZYY/5<&:85?HS,De,KS97b=HQ?KXQb;QQ\7f_OKIV
4T8P(#82/3+Tc6P-E.QP+A.7Ef&IC&FB+;]7)e#W&&J(UQ>T^WE,cb@U?UCQF[^?
Fg1O^\,<X^-.e8.5]H91f)[6fJY^T(-EZ+I>K6M-SO0_PY6WN.9ZJ6L/YAdWI(IZ
Q9C_:QNA&#B97VK8P9+&45cU)fKJE3RPgZJ?124Lb(J60628B<e[,7&._9WC#P,U
^R,[93b=>#SMK-)FNW?[P7R,@cdL[D^^MOTT/@VF:8EIY4.\^-&54Z:>Md6LEFg3
GfD4bd6=X;QgA^<\MOMVS:e))d6A6\C&:E76FKQaQRL+:+A=B;WF;<6Q:b?QXC\-
SAe@D#<efP9gF-C@[-RIa_,=c[HBD6O4f(7Q;6+Z4LNYRbB[+cKO/FK-ccG/]FFd
M>#5:T][69Dcbeb71Q[@9QP?5>g=Q?eM2aBQfL[5O)aDb\,>H0I2d_0@2<#;9C];
ILbFGTa6:Y-E22J[BdZ5;E1+Ff>ZK@9bIDA:3a\9IP;b-2J^E.?N?MAL.J++6G5D
.OI3C^UM3[INN\PYdJ\?P#D)0GZY23MQQ-YRfe]ZM.HCQW3RG,B\OV7g5H1LY^>P
g)]2@;;PPeZT.,L+^a+^\M.G?\b\[0=g1A,;)-]^?-^XZSb?/_C\()_/OS1YZ<,:
]V>95@/1<[0EaEJ,.Z8;fH\I;.31[=K4T7)\>5d^ZNDd.P&=)8ZZ/??XSXcC7J<]
18g2X1Oe@O3RHY+3I6O#@_<+B>gHAJ4a4Y=+&AYY6b?.YL-g2:DM6UB1TRFFPBMA
KP<E/GbgMYXR=>-OcFUNd3#4]EBeV&_TR>X3Gc(5)RVUM)=MGP:PKSZZ.E#@XeGP
:W3=bULM-T)KN8Te>KVc6^HDCQTJTTQ?=Sf,Y9A7762O#J^92CL[aB?7O/O&4=c7
d&eMQd<5fe&3\a+&@G)#b\:BT_ZXd_3].)GQ@3K>fJSK^e+BY2(?#?+aTcdE>_>:
XbLg0J6LRKE;34db]U@+EZG0@=7:;@1CAJg729<BNH>VY7<J\g.J]4\?U8Z[dL#Z
P(\CB?8+\M;-e13UH:0UO2:dOfZQJWRfeJO_=@(5NU?1c^LT,;d,fHNQE;VGX50H
]4a1.^]I;a50H[(J4N(>GRGVOS_MM&99R9;,O<LEXO7-I+2>8@)\eSfaT2H;)c,-
(RQdE[XdXM^Wa=EED\PgB[Ca^]YKONZW)c?;9+85g9_,b&:GUKKOO2EKdgSR0[A(
Vb.=MKY\)4e37V3>,aFH(1QS\V=0+WacI^JR<e[XM&VFJ7DPBV,ML3?XTbHXBBeg
LTGO#a4d7M(/_U4feE1N0.TPI3Zfg5fWX2eGC39EYLc0)fM,Jg8(3gXIQ3D/aO5@
9)X0FMC-3SZ4DOAA[^O7WO_0Q>R1HHbI^&a<W\7)@5-&3@JX^&TT/S0ccCT:IK\A
E2W4LF7>(JZ(edTRG;d+[bcgOL9L)1U<>\>R4TP?MBcaeINA[bHPRca38[JD5-=?
;(H.Q[=\&Y;^=:IV7M3_]:Z6,Me,QRT>5aN7LJ-ABdad3-b^,TI-b^,V+[0cY8g[
O4gVeO+e8HfRBH^C8(,7T=96MRJ=(N#&FaJSRGN3OW9c1M4:.Aa97S.-_8TZ+\S3
>?7ZT3O)=PeMX:8FN;gTB#(W.d4fLQ(TYFPQ#.FWS5JB0Q,E;cX&_Y[PJ>?;RFa1
+?WWW[:_Se&b@.RQ&+&Re^HW#WKZMT32eW\?QL(<+NB>FGQ@fX.9Z8>>._VfE-?3
KUQ;4]HY_Xa[egJSWd97e-^F74L/;3YVbCaYe]WC<;]53fE0fREeI4(L1cgA@Kf(
C210MEIa=3GG]D7+82VN8@UM^b:GY38XTF1ZRcSXN@4JU;HOEN.:1[1.B]Z;1=X[
=K5TB=:^@>FJ6+1-X(G^AgC@H,d):gC.IN;X&d4a67>3MY\U,:3Z-BT12)W)@4Gd
E3Je[H)YJW_0\L4gcK4Y:d3=/,Z8=M0<O[J[8+(eSdCcdQ,19@Q,.B4AH,\0FK^?
D:Qa.+>KT)7[95Mce((]A=[YGb?f+>M-&C@Vbe\M?UR35aY3IAB:\+RXFUE<K@[/
[7(QQ5&D&W#LB_KYaDBB/a/L#b[A3f>6V8FIcZ#5>6;KIJ<),Fa#gJ0Y8fF,VZR3
A1;EFgS(W(b^BL>^P;<&(fe>c^.:07-M9J9+LNd6+X2.3L[-HO;9+_2a<PIF5cf)
B=A,8^5\)<^Dc<#3#]gUe>-?3QcM)2+aLc]Q5eR-GV&KN(7[W(2C,L+6d#8@S/[c
Ya+)Y=b-=)K2=:,4CC3]XFU;X&V.RQU1KW6ED_ZDN&OK\N.dXB5OWSZ<6(9A53X7
Ue<(C_]-LT3C?,dW3[>0<)=,C2(G=]Q2DH4Q+63O=.53c1>I7Z/YM21HBeD^.THL
BA?HSN2:42G?CaZ./Sd@88Z:T4((G[3ZI\2]2US8YLdXGC=\;/->@6;\;cQ5&6]g
@00#1B1-6a)Z^AP4HRMXCe8FBeJYCDfGPfLFZFYdWK?\1<K_T:WGa.P<LVW4_-a>
R&99NHE2G;W_.4c8DWGL/6L;L41aR2SKg2^e,0]:T.L@>POMF2_8LG=T>6cZ(dR9
OIAIE\MEfX;[g8+_(;<eZdCX#2S7@[JR?B3BC[TF26.N:0I:ZKgA&+CG,A4[DD#5
\(R(K9O[GP:7R_6ZYfY7X05_EY#fZBGS5bBRcBJ3T22-L&7E]Z?-1f/&=4Pg>>=D
F14;^D61Qe+;S5^MT<]LP]X(OEBc4EU&\W2gaB6bE;,OZaS=YN9_AN\S207++.&V
EH#gC/^XccHAI=.S/BOJ[c.F?g+WNH=X),CKF_28=+JgB3aL&Z,@BVE@cg6@0R^.
J>0>[<C#QLZPg_^cAKd;?./HC98K#77I1)10e/]Z^F5]-L:7-OJf+M^-V(XPV/V]
NQ+VN5N>PS>J0KEXe+H7NR#Q)EE56E:#S2^7#LWL)M>Ce>&S@C<bX(CCK.)SY2;c
:@J.gab,H(aOVZM=93U[4B;:Wf;_R5fT+@[@CgR9bK<.;>OLfE?IXbG:NNIUHWA2
d@DAPW;>&0>9_-BY=708.TbSL5DHE.a(dDaI00KQSL-U4SdcCgYZL(RLX)5@Ec\0
2&)U0+P+DM?B84GcSe@Q2MMY\T;/<Q1G?fY5d[FGc,QegL78IQY@?Z1IX9VYWUd<
K,YQW76R9WQ:b3:X;::M>>TWQ?G9>&5XJLEQ_PHb[ZA+M384B6J8^H:T@OgJNf+2
e2O?OJcMDf^YK?=Q<@VG+@@F37JUKHMGV2<Nb)J(W5V=W@6,-[@UNQV#VC3>9^a5
If0RFg4#.HW[QBdbPOg<+.C8aC0d-(A/K#)BB-^a<6R>NQ[57]eO_]AGVMYII-29
&<J(R-36QB9/C8]O\N3DNgB<0;7+ZJ24F_P>Af#&N9YUC+0;VU@=O2DSIOd.G\/b
Q_bg1S2^-ZL)e9;6SQ4+SH(1>):R(D]=&KL93aGW^VLaR^U;6>4MZ8eL3UHaO(^<
?D&Y8A(W#?&e&T7=8^R&T85XNIJgV?/N+3M6[ZJd-OJ\XQ-&#g&A\S,:#&G[&O-;
):2\W3Ef4(dO?a-W+?9dZebA,<+2F1d_8F).O^^J\L@9EM6.-4&U=14HKc@aV;=_
b]AA,U3]d4NSMSOHcXGV,N1L;Z[G,-)AQ0FA)J)d#XWfHVfe7QJK_MP=Hb;?#T]W
I-Y0cG1278A(#3a-B^TSeXA&#U6HfB<@^g(?c:VUPe5\\N^5=;V1EF38Z85d[#:G
#Y<=0:aL(Lf=,[dG0c3\WTQRWd4]SX=@IR0\1HdX>Yc_-)1BT7D[17L[cdc8YT91
Y4X_G^9fbB/3N-+WZ@c#5gMC[SRMS^)95;[.6X0X>\LE,Xg+XgZE3J](B4VU\VAK
837aHgUN4d/>EBC&dO=1gJWAREQEa7AV>NXXYHY_(H?V/AZX,Df-GFgaT\aI-W1B
P,A@b@#/(5#gVg@YR_A)4JL9,LMJ@K9AQMdS&^XGe7FNf]^fW(f>7CU#<#a_P?4E
U2VDeRfTKeJLg9GX\DYO;(8-)Na_cM[R[N>[&9[D4^GEH[,ASfB(f?GG(;cMeBe6
;&YJT\>MFa\T+R61YD^1@dFF.fb\d_GS_c(8a[H_Id=C)K/06fZ)S;f^U8VP0Fd-
-18O;6^6):aW)]K9e=10=:T^Pagg<@X,6XS3=BI)Q]WX.^GI?5&@).V;ZX]GI8>/
L;g5<O;(94,LgQ:;278[0TLfZ7Cg+>gHcX<BT3XZ(RD5S^dQ/LH@]dZM--]>_cXP
JgKT081XCH=.M35B[Lc5P:H@<d\_I@5Y+dLF:;9I)PM,1,WY:gWOf-P#W]FS#EK3
0W66HcQ-=\_HU=-;1WG/U.e_5AWHQJZPV:NFgPD0W#+_K=L#.#)Qc,9b[Zg^(J[c
6dG?Z33S<>.@Zg)Y_6PNdFP<5>AM_US\Z3\9?[)1=YBP6<3IOUcScSVVLTQVP;gX
cgN-+@cKb1K1=dQCKdU_6+I+1_IRQQ>3EM6bSQ#I]c1A8JaRc9UYG-d(1_?L8aPK
I,,:3gYgBCQdFRND&2J4H>O2]L24QcP8_/F0J4c7;J8Y?@55fKfK.(QP-C1H)/8(
MG_,b]G\)U(>fOa>?.TL_ELDXd-_c8.F9\T+K8[d4B^))g-USIQ9MRGBHbd^]C9R
)<cc^Y_5&L083=P0]8e.e+-MM6>DcfZO2:6dg;P-147D]NKUVg]@9B2d(ccf4?J:
d:>ZP7X::0^W0^GEZfcL,5W)g3egOIH:77@GLGSd1OePO#Y]RSQ-5K:JB225\PRO
S\=B+FZ+_,=GL#P+)#cScMDK#&)E>9e,GYDS#\1@DG2,gM7KC8)0Q7/R6_F(3-E5
EL6=P+[-/6ITSJ7JY;D1PW\5BA&9&:I;W,0cC]Lg#2,PYK,&/RPaK-c4:f1#Y4+W
6EIRdM<B+ZFZN@>:@ND;=6-KM=[PL0>Y(SON1S.@L/dYCUHc]E0a]#Ab/b<0-M;G
&.\Q7@?T8Z,MaYX47J=YR+LX6EN1cFY[PWYJC:K2AY(L\VcG;P7L+BXKAdHRbT;:
:2_@>)JVf(3(:QUF[<a#:RL5V=Ie2]BIcF+V(1OU5?&YY7F8aQ^-;D(2KfWTR71N
JBOD?-<83BTPcB\KVJAAP[dD>V.55MKdO,5)VSL)Weg][2;MCFK7d3N^Z<;ET+)2
5N].3;NTIPK0Q;NW3+a]X+KBL@Hd\A14YAJWC>JMS\,DbM/W8DBe;S[Q_4F-Z#;R
=[RBKT\KKY3)(.5eONNW_F\O-\G7L(AG[NP:W^[2]ScE1\[1=)ZTfc.>.OPI=2H^
Y:8(SP]I?VbA.Z9,SP37Hb]DQY6@FO^1+09@^67NUf=F:GMf2\A@aOO3W7EeXLBW
:5VONFW&5_/fKQ)XMJ.&&;LM0REb+5X.D-?2N(0WfBBTS0EgVZ1EKBY<P?#>4QTB
4_X8;fPR-350g_aDdPb((7I-;GFLB\W^B\:6SY@7N(\P;/2U\8D?B?.fNMaR0c8:
Tg7)>bAXDea?-\]>1fO+:fc-0:Q]^R#0X-G[.VFD:[)7P?>,7=V=62V9gHKf4;aL
Oe#aI[LeOUf(b:<)7We>dK2R,e;e7-bHJ&eN3_3Z3->Rb.WKSATVV+Z[:9>PXUID
>I2)3DY,3+UR.SaLg]:O9gJ28.AQGQNNg)G_Vf,a/&JH0./_fB@EYfI&E7e)D0.-
8<a91GgG7GODg1E&gR(_Ab\.=?SA58\A+7+\,EP_D)@^<[JPE=D^,MH]Z\0.Ob,?
]F5,<1?RK])0/<#_15O&SGOEG0FcD[4)?+fa]J\CYf);XQ)Hb(_b2,^WB8Le1cJ2
X?8.)3?8S6e]I&659>PW_8Yb91,]8<G7#8>Mb=X^dRK97f\V4Y;EfAM6/5-fO@?C
7VeVS>O;[IOLAK4628ZNH0(JTd,Gc9gLY5gT[@N4#/CVYaE+Jb<-#RW3RDAM@^RI
G6&(&XWP2;@4W@-c0J7LJH7=J5^AgeR\@Y./b0cZ^[SSg<8_U8=ZQ/.N9&1Y37N.
+,F2GYP=7QV5=K@O3Fe?]28BMg:a>NHT4J-)8Ga#X8XM<]\#_]>GH=P3L+XT.f0Y
7HTN0GeY6NGV_Z]+I4MObd#.3)ZQ>,/JO5PNc/G27RNQ?<:,8_0fYYJ#geN05J:#
+E6Nb7@HSN_1Wf=^^CTIIYTg-fT;J^YNF&dJH[=DL+(.eA0<?fVUI++TTg51)E,(
PL,A,OGYc8?C-<ADR@Z)4USK6?8Z02M9L7)1#LOL5Bb,1aJd7a64W0QbPa\1G9V8
bgEKWX#=QKa_L;MB[aIO]OEF5#BKDO8baGKFX;RHaR6c/93A/a)L@0XX#C]HC32.
96c3QCPCBG-KNOAS=S#WC;CJ#Rag.UFUK+8UTT/<Y&?EUWc8ZUf.7^L0aN<Z7_W<
d^d5,[F6:Q>(T3=H(,WZXC>_ZWDX+.0].9fXeWNLOXK_3I<XTIP?gKDbfY/M<NgL
9T>;O.(Z2.5L:eZ7>UGL7N<cHIGK=KNFXOfXb6A\;R(g-E(@f&2ZS:.LcIFZIIf7
ZUGPC9F;R2V<Z_dFRe.-XPG9g:51cS2gJHLNQfGP#DdKf>BQ_0E_@ZfEP/?RQLd0
>(Y9[f+F;D)XJJb\1^_4-HX&adT#ATG]b]^E;]FHa+[a?aJ:F,V^<(BF&HJ^Q/5:
F4#+:aAd\4D6Dd-36X3-L^AcXdGVWg@(0EJDT64R/06K+WQ_,0/6QW<DXL/>TJb#
@K&Y>ZbRKU;)c<f,&KSC1&-=9:J8Hg8bgd3[PeMRW/=)X2692Z3Q5##R;>I2R_b^
J92G=Ld\cK5H.O5c/W&VY#5:ZLeX)L_+0R&NYgd1AbDJ9H]f@d5^KYI5@Gb21&Q#
+ZbO(aH6GH(#MAMN5\]cN.agZLE2F9\f.PZIRX(A63JMB8E;f65U9B)3aUS#@9OF
#().cIU]@DgdUcG7H?f2)?;d9<35[eT#-g,KM2[>\4[)@^EI^:BQ9#-F-\#gT:+D
&eIA#g5R=<.KPRc3G\;I7PPKd+L.,JNWJ#GWGHON]WE_JM6^5O6ZP].VJ/]X#)0;
VaSH?gHB21FUBf#R)BA1^TP@;/bRLMD6gd\9><?;CW>AOA\J\4g3Z16_Fa\1\f)_
5)9Q#CcPO+VL)4M1TW.]#9?f71bOZBYB7:Bg8?dKRW.VHM;7Gb=C<EGOc3QC:d++
4.Me-aD-3b;M]KD?28ZLI7@#a[dH&^K/DZIUV4g>8UO?IGMc_,W>Cc^a9LB92C:V
SDZeLJA&Fe4QS#^B7/6C+0CO\SNVW9A/0G/AEU?)3gF.P<,LX<8/_&d2D4ECRCc9
==NVUJ1[EP4OVd1=&X^M4;YK?H6Qe/O;RSA+8M#WNfa#]E)3]C.d9RV7I:I_3gZN
D8YS(+Y3H?&Pbf?YV?<:dXB#Ea_YIS+ga&S]W-.&UYeM\E;M1VYUBTS:D#2XLSSL
:6YI37[/b,0&5^,<cT2^#c1_O?[1E^9\O=TB;L&A0<?I=E&\b)R<[&5_A&Ud6K5\
7<c&KOT7#,H-NK:VC:[H8WA3dICE<2H@A/1&G3g3P#37FMK^&faI;9D<,14I+^<f
1dJ650[aUbVO2>++:U:gAJ=QXW3dg:[Y3Bf/OJ9Z5d#MXLe\BVT2BC9;SKP1UcVc
&2f;RGQ8M4MN94^)#fC8TLKNgW+9dQ=F]<-U>JH-K_I7Pa/PDU#O/\XEXb3GaAd:
_-[E53<T2GP@fJGY9<^KCQA2dB.7QQS&TW&&VILbA?@[gCL)P\:cXP3T=6CK4gK)
QL@@E-DW,E[TAH2>,G6bVC)RG.U&Mc;NaJLYU/BA<Rf)8&;46TgaY#EE0/43DC@=
I9CXM4gN61Q)]S]a/--9QE=I6aeD_)C]VECCG,TZ3EJ&0=GeBUYa#[4)&K3NPKDd
_6)&Xa[B#74X(:-gN[6NXH/+BGK&<]],a1R_d^P_H32^>)[_0L:dLVcJ&<A[/E\9
cZNE701LeYQ&JA-<N/UMc:C-#)A?-WQNRgP[]=[+c9W907ScE0#G^)Ob\[@&DWgG
F_QM09fc[JYbY9Mb8Y96ASLcNbaX7Mc)>Qb4XACF9g6P6@A+?-ga-dOd4.2_MW4_
R12C:74:[?55:/VBKX(_W0D3QaM59UH.47W&^&+[J;\TY.a(IA85.Ee)3473RRPA
AIPb>Sd7DefbT#U/C4SU]#PBA\PUCbD)BS=/:9LAgL9Y\=5S+-#W2f,X8>LI:XO,
LU)151a^<6^cVb,X>9cfJ=HTU5_LMcc2M;L;V6LTaJ=(3Dc88Ma@9)b1AZDGO0?F
9c;FO70.#R^FTW>3T\8-0(K-?O?Z_e83U8E]P+M3Ra17/L,I&CM80>QGY>2\0U=[
Df.Sf49X+D4CcV8MUIC,^9KcePF0ZLAO@JIZJS0fC@H_O_0e(U(Q.F?XD38SJe>V
SG@_c]_b<c.8H^SO>T44#+Y/E;aZ_J.&>CdIHEMa.DRc4c_cS-#7J<HdQN5R_K/B
9TbZN?NgPH>A4W9IOLXTE]ceJ8GD]H6<BCVEU/(N1:(EJPeS@716HO:4GK9-UUED
7D2b=N@eW08])0_+LFHISPS5;aZ+K_/#@-.P^T5K<]S_1=3\4L9EN-fKYCQ3IHa-
SIb0(W8=U2eN1-@LNC5ZPIHXFP>X8F9H_d,C.GH_?DA@\QEY\gU7(H9G.)Z[?KN1
Ic:IYMCO+(MXZ)fCFN6Z@0QKF+IRZ9NWd9E7]#aQ6Xd+<>_=g,.4^O:JGQ4&T@?:
fPC.6eCOJ^_B;9[,(:04:?K9;XU0T[:(;F<K&3/KZ()7G^-:AKEd/,JTGY[b2RIT
-O0QbT59,KR(=V1_/BR.<e@\HG9>._^@-\K^MCN\5NALE[1HQ5MPOJa0QR.+@SBB
NB[A?\W_Oa]N6;<>YQb^)ePAJYG;-N?E#(8S)BYUA3)C@YaSW5=O3R>D_97d_N\Z
)IFM,0\UaF:Jb=UUJ.P(SW9RGV-]H8b<@A@P0&>-Mf<WSNUPF=I4DO1T@HRKDY.+
dCM0F599I>I6F0)L6f/6^K=0[TDgNMX/OW?<0DI<+_E_Q_8UT4a?V=cCea0#;^/J
-59aOdXX[(V0S_g(/RRELfD?Zd-4d(N;]Of)dbC&Y77:LQU6GgMYHRSea4/?X^H^
D..NJN[#U@,fS(Ig)_LF4bS5R9<\?Z,U-\^f;LM&Y)2e]SG8[Ie@M/(L^^]]g@QG
9\D,@fQ>T1:5<>\@=fcI3DGYLW0OBLXYWaD.bM[U4M0/K^f&=#=dV<LB-aXGM;)H
@c)cZN\RC4TLX#BW]c5>7O\HdLFbC>^_ZW&0+)gKHJ?S05UW^/-2+7OZ?CZ:Y6N0
SA3?)L?D/PK9@a#WSY4,IG[#TeVeA#gOHDD@@/[f86-E8U=?8#Lb-[HI.Y9[S-LK
\,\N5JM-0QYMB;FGL&&XI-^B,7,^O:_)2=.WEYCKe?:1JOK@fC/(0SWX7cdMXA9g
WX4^P@J7@(]G&K9#X9XW8ZBR2-\K.^g@F-S08#B@a[1fR=.#_UBeSEFRVHEI)Ca1
43[e>)6W>PS/b]8Z5f1SB5@TY3,ME-P6b/[1WI_A+&_?G3&Xe73BT/[I<#][BNRd
bNGJ]=1_[UW&F09?NCN4D+S<#[&>[\b@#T<gGU4+SFH]7Tg@O7_d2Ye9.B[QVF-1
08)JV,f_a>QJ@>JGE@_B^;6_#E6I6\R/W^QLF.F]-Z5PA#/R?EMa=0Sa=\B=(cPT
L^64L7YMC&?cELLZ)>eeGAfeXUO/C6.&:c<6[\DDN-FTf,?5+b@&7LA#0cJCZO6]
\CT@=2;\=#_ELQBV:46(T1?Q6;.4(-Zf[;Ha:?[;3e#fURD._NCA(9GUAVJ+1PNK
I1U>.PL<c>T[VA(bP;&=IB,85RabPCe9+,2ZedA08EB@QH)@LS_&-eAgbKJ5(b3Y
4eUA(Q/FC_.]Xd6L_6\e.SHEAF6^Q7QX/ZF<YV^a39<:C/)ERIY[EZ;?;PBd>C+?
:e4_e)/.DPA-c,-+?.S+NcSY/H4277&3[d8\f#/C-[65F,AQNEGOCB4XaT(^<OPa
IXaHFdP]5?c>^<PG&]^5S)ff2,d(SZ[S&SL\a)G:;AAJ:ZVMHJM7^_FAQJ;1[A(4
X8,eaW,7/d[YLY6GT.-7_G-@3G]+MJW7fCF8-XT-HZgVX:#YcF0>YWAC]1]V@_?C
/J&O[;#B.@e2D69WWU-e04<C.dWGaHZ+gTg9+EF>0Y]Kdb=BH[(fZ^+G\4V7ZbFW
_=W6)0,6;Xba^C,G(0VK62AgB3g>YRc#5c31C<=.d=HA>#U5UMHZadeI-YPCO5JW
]e&3W6B_20If#F(?YBPeH00>FG(\][Q;TC2WG^S3CRXMJ6ZUB=0P>G5F0=3HMWa2
AgICQ<MSG<bb4Tb[38/gHc3UX-3f1>[B2fKX-?;;e.QPIfJL)e5.GK\YDBC6,cVb
,Z-?DNU&,U/PMDL._^N6/IEJ>,(SNY.#g,)3>]E(UB2\@(3V^?^/[Q<DgA^aTWa+
031S75]CYKD,]cD5YK0OZN[42&?B8=JSPT9b4@gQ0:XYAFKMRNgNW5>gI/_B&AZ4
ELPfI@?P]EMDR2=PUJaBCQCF1&5EZZfT#+7Yc[SY1GKR2)?Q.1_aAYPYdJUBeR-&
+[D<1=LV&c0e@Nc[CL:>VFT>@_T\-OL4ZP?:]4GL020>C5?LaY4V9#^K>7N-TH)N
PfdeM4,L;\:/DJdd2[DKeL2g&+^<0P(#-AO[\c,DMYfPQVQ3b.FI)J0<_Z09H_Z@
Y-e/0.W,X7;1>8P]@aJY?UHb>VOdND<NW_3FFE<N^Xe.+?0,WEdKBL2:<8(V:_M1
YX6W4L?AM^WJTLL3OeFKH:afE)1W5S>.G;Q?Y)4]18<FGc,,[C//&gRe<f_NR+Cd
9O3>YEL1e[:Tf^P3-Q:+#4PLFc0EJDVKG6]TOa)V^b@)/(cbNTM3bM>C<<UKM?57
3F(BOaLP6J(L-5W;e3)^JLZfDgUME:V86R<.X4gX#>)\@=2\2EffSE?Z:&H?a?)H
\F?1TV&R><]1?_:/_XTOS/^F?D?ffZ9.a)R,<W=?V2Q&^;CbGffdE,c\-EMS\VXO
M/GCHLSXTWCK>HQeM(]ZC0g8+ddER+6J630R7:U[fbbdYe@]e,:QA/AYEe[&e?;+
=eI:+HV\C(&;N]aegOVbAIIC=)gVMR\)(P;T?4@;IRD@/9W&(MFXXI_=/^:XX-^J
<&K>IZe17C?[S62G.\HcQAXc@X[(<P6#53GUed)5>gC(bW8_.G&A@eLef2I2d=<+
)bB301MLCE0bYb?XC5Z3,@8a6=M_,4Pa&^J,T,\//LL\HX^LfaR0:5eE(Q<Cg&L/
bS0[R6,Q/G)BcbS[W0a:f&deX3Y_7(:HASTMQJCC),6XRcAQ[g,G1RMNG<<2BA;d
gH6/8@^-@Sa1-C_a;25?M.?JbC0&_(WU2_D5OA&4,H,5fZgZ9S.Pb5W,JP:e54\:
5.;,;27EYU7?3>^ML(0MV/bDdYG.K/V2C5#59\cBbU)eKQX8U\0Ma8:G;NWA7@e5
8BQ..[A^.aJe)&L>I@Eb-YgVU=11RIIU>dB:?efgL.3(Z,YX^cKT=^BA>>WBEYLS
;5<_/=:O.e&^fOH_.:K]fX(=_fWX]2-V&PCX-W]SHI<-F,=LRJL6@L;UB+5aIXbM
KNd\0PA?)1>TYTNYY0g8:&\^Z/BX(;7]:AP6XD>&1.(;YD6J)J.P#g)2722,,-)&
gMc?;.>QKHO+)-48]OA?IVV9MW<_bBMWSg_)SDLSUe216IL(FTR1@IC]>ZZJ&b0T
[J5V&/YJ;URJ8+)X_V0+;#,6OB7KRfVWXD#UV?/2]2G19T(HRdMFFg2<L3\2S@#R
ZEEH02gW+(+.fR#Ae<#4fVZB9_29,M\0IT0+g06JUZ#:SVW:2D@eO_Hg-_WMKb3R
U5JJT&OOE/.g[W8=X5DE)FW_M+646_F0g/C(bd/I&Q0MY<U0_8IE;#acZ)WZ=E09
YA,;Ffaca0?/S>WV?^c.H48^I)aC&B[,[S]3#KbK\DBe=P@)A89e#<K&ORLS+<^-
YS@#NRR,S1R23R8#<VJRScJ2/U1TPB4,;[4GM7IZXZBO94J,43J:VUW1P;YQV5V?
J:?AF.]7Le&AVgU+/L[A1XAdI^LZA;(D1\H-:S<D@GQNN.<UX<5Q0D\SUFYBD25a
:)PV/\5P^1SZNI:FSbUO+_UAXGUXI(b+>,)D3GfC?L)X3+K_50g8W9Xb>(;H/Y#5
g4AD<-Y5]^?.ZI@0[08-3d1P6A>\.YG-J2N6YJ5a[ZT\_S?eMG:/N]]>dgYOZWOO
LF_6b=6&\F@<+_5,Nff-(<5-&B/0NSD\+:E=H1@R+90d884K7@,M.QA2Bc\A-FRF
HB5GU]NSEE3_#1);]^fB)P96PDEJB//82BR^.5&cBGOZ;ZB5[g40:I9Z8,geML8C
Y#S7e_de0)SX1:92+VR&RRaY7@:\Z^>I?>=/<DDTc</Qf:7OFP1f6bJ/?A9SS7c-
R5<S6^f(>-J6-.L;X14DY<#VJ9?R>QG&/4U/F=;MKF:_2L;&f3P<bTMBA8GQd?14
:Sf82Q+7X-,f4=Y;?[8eD^@:-QJdCIU/HgG<G:S(bEZf?W;9I_I.LJGA/K9XB4F9
)W=:g>^)Q-U9GWMT1fLADP6&?BNSUN#L;D#?=_&H2Z-K)bdOEbcUU)]+c_CQeM/T
g-08XeS^.U2U=IJDJ)K55BMOJ5#(_RBg(9,QKPMOTDgQ&L?,XB_V#FE>=V@,(/BH
@gK^cPB^c[XPV+c>):W&S<[d3Ga@L,aN]I^\0C9T<4-&PYG:2&:8WYf-HaYVZf#b
V#&]+/3KFFHbbMPJAee/8O\/3,Z.2:Q-LcB#[#UK7J]H?<V3:B8dKFT8)>BTC=DQ
EG9bBC[\H<-E,43G=E2ca>=f-MZ\>)SW&HVEL:&3WML4<GV+5VG4C<X2_M<9H0D&
)-:I@^F>OcG64ZI]X9eP&:_0KFXXDfg,K_=R+H&5:B,<Y#gZ\LHTI#O<#dZ2S<Pg
3]&TWBP>.AD>e;1>6OF1BB\ZaTfFT0Gb2:]]MXAfKC^g7_Sf5^Q5dJ3Y6,;R26)d
DdB6a?7W4FVd]N[E<d0gX::2MfDb.INJ0_G=+Bf-R&JL4D.DZeG;Y8LXbW))X?[H
J\eSbaKU?9A-Wf3M+8(B_U>:0eI9PZEKB5,CF=L;&7W6+c]EP(&VIR0K:4CHG78.
I/7c7+ID@34JHfD#a\&GW5NUY>N7C_/75Bd;Gc_ZL()63V,,:Z&L:+L:U9d=Ue/S
J9^EBKCU_=A.P.ga+?K,UB]0TYN[Z-6X1L1;QVf;GJOUZ6^Q<(f^O[_YTVW[fVT>
4fNL1[C;F671]RWU0JDW7F(Ie.EX.,cNA.[UaP#-@-4cW:T=NX.-fW,)2^OAW8=L
,QXLQCQF^EHQ5O6[O:R/0M=OSTF5ER5<JNL[3U^@3U3:>Y,U/g4ZW)eHe9G9a@\K
J7aQ5JJ36OV,2M-HgaEcUWOCbf>Nc?3QaN#\caYfX&9Yg^P7F@9&-@&(#3dF1U&b
U\4NQJFQfE?XWZ1AJ3U+X5F97fOU?GVC10@@^?B0#gL<3??=9Ib57:.>2=g+]_-;
5)#[.[MYdREAdA\bTN,LGFJ4(<VB883Q#A4IWVg#SL^?JWgJLdI[[OCf.6_Pe[@]
Jbfg@VJ#HKXHB0<f23P7.D>15e0:13b>GDf@ffXN9\]31&E.;T-/2C.)2.0?]+LR
?F2D?Z7.?TP[VX[7H.W]7Ac5C+=)W05W5?)bF1(^aA6^6U@/3HB0_SU3>_TYQ+1c
f(0XL7]@H(:2-AD0:D:X?_@Q8O)PW6)+T(AM\Zdf/]N\5g]\6]e-G+>8SU,MeB&V
3eC9d9]D>-IV5I@N>BW]M/OeEZ8;U(F_937L;>194CfgbD8A57cX)4@M4bDPQ5T5
-N;7db==eQ;CR&KB+f?O2ZbMM3M)IQ@2]?-ecb/O.LN(EeBSVHQcNJXZZEaCP,@R
NeQ,F[@e_UcQT.VXWT\Z\g6A\DH.,;8BWB<FM3E)#S>S:4)6g\4C(8?.9UUL;)F>
1+T:INE@7/1.1_B/2,c\;BY..<XK//[Ha89.WFUD2T[_V+8U@@E9)<#BASM-/?DV
:F&HCc#Z6^V^KgDdVId9S>aXb6b:75P6L3eP?NNe/f(L;-:>N_@_;fM=I\@B5Z+b
EB^QTASYXDMc42;gV)+C,BPC,Q2M;1U&/WBYbLa)/e\_a;gfXD9D63,Q=QZH[:X\
C(c^b\/_9S_8Xe^KG].>@@P/]4.Cfb<</B42C)cPN?;GB,ISW3ZXTZNf4P+NO]M+
6JD\f60C2?^M-T<XN^eUE1_:Y5;5<BM\]K&e^C5IfVf@EZ9WJRHK<;T>e3d_J>1a
(LQ#>.b6FQN>11DaB_K>3gNI5+,EU8Y@(fD7RBP2M8#J0+?3b?LDcT7D4@7VTQX=
NJD7>:49<+,gW;LdH-._9M_7.5g/6[C75)AU/V?FbJ#e4I1^NDLHS,Y-M^\G?5_^
PYNU712_3BdaCM=Z2K5(0L8e8>M]6:aF_6EaJ:VS<^(FK(18OFHbEH(=@BLJ-&Ge
f+=AAVRC9(cU@)g(1X3J0BB0F(QH:CP^,[-R,a5\:-ANUV/A+8^X8@GJ:@eS;Ge/
)13cP#,@7LFI2eA8O/;cTGIgXPZB,Kc4NA78I[]/f\=>W7+_0;>KR\M>^V5S#33V
SJ3S/2_;BcNc=13#JK2ML2NQ\@W9.))c?Y=45C#E=d.daIS4A8=^DQ0OUZ&@GBE[
>22?MF]G;+1K]]I30?8eWLYKQ=?fB+dPI>>2F5>8&T@Re-SJ0FGX^>4\IAN70LSb
H#_aHXM5LCD_P[=(7)^Ad:U0;JAHE3U12H&2Pfb^OREQMY8U[V6fWU;7eC05ee&D
5@8/S9Va239+YgBSSGRGRXA2DAU=+>P:)&N:#A+I+fDI<-YY07&0E7XHgcGO#^5M
f9+R=Jd#TELV@JKI30:@8@#B-BMYYHMFcQa=<^,RdIf>1<3XCX(+5+c9#(=[?eXX
5H<-aReKIJaYM3d/_SgBc8d?b+H.ID?/BGeLN:]<QaIJB&e)MKCF421RL?0984d1
&7Q3MXBNHM=](;LU^O7:eb)E[9:SB6)6D4T>4FM1X2>B[@X#;XcWIHR9f@[2QYX&
U,UGaaXQ.^[VgF0+OJX.[(91.VAReL]R<:Q\4/H4<D/,HPP,Z[,3GGU@aGdQ8;a+
3QF3S7ea=bUb9=/W3KWK8Z\3F8F6D0aK+c+0Y8C6KTT8S:U<UbFb<GJR,7T@O95[
6HTNWUO:X;R419D4(Jc=aBUW@TAf0^b]SI>LQ839g.,AR^J+gdLC(A=[GA#0ISCI
U);6,M2,1,/8?B:RCZVF.Z=Y5[?;.KPW1YTW.OU=6eY#.UdZV#b+fbJ.C]2[]P.J
cH8BL(IJ/4WPd.f7LC_V-]8GL1^3\;B(FB9Q#O;_L,GR=ZE3J,gUI5;#U(XGM6e2
Z.Ld+/cIGVBDS(Za?X4Db(-079W<9<GZZ4[1IT4e?HI21a@:K43>6.a&U]/J9G9@
Pc_K(G4(?c6RP7LcN\^\1=MeB5-K43a\gK^TKf9C]aag48O?64@R_,KC07=c_e:/
NH&_CK9QVWa3__A;9:]XCfN1d(\A9d0.d&e7_6C7KdeaOE\gB0e,6VgD[cJT_7&d
W+JK:d[9e343JSa#1D\]WF;P2/IGW\RCa)]CL5_4=MM/DYJ6[g&41JfQE.WeK_b:
a7dU\VN)g9<-TCafN9.VO81[M:C/FRX^A=aB)<:(_fG(2]&KAa&e&JA[R]\#4/Ud
33Wa[MW1=(260GZdNcYX5T+E7L_T>VR7U=f&d^V3RccCHf?dFZLQOa4+BTWGS_Ua
3Z6)?W4T1b\T+/7)c&)HLJIL25Q4X_fe?e-74Z(QGc7\dMaFD9HTT9-M,B_@UC\&
/JA\f/bD]f,\7B[5NO9Wc_WCWW<#0Y@cR[=W:>)+6,S:&e7[)fK920J.URfKB(8V
F]8HcAS\]cFU6:\Y0-J,Aec)D_1)Wd,3KAVG8^U:L_Ng5UXdOE.ETe0KDAI<-XHe
V?:OX(+g/^2V59bT;O3T[^ZYeU6,HB]XX+VM,IC;\(<;&2JW>?4_8>H2QRdG87]\
,D(VMFHRP9A_4e>De2TZ8(YJW,b+]b.<)V<B.D>)8Zc9W8S#W_DM;KZ6>9^H5Z+(
14VZUT&SAMFH4NH?IdEM;P43NP71WXU,[e+-;6&.#JYg7=/VZ[L983:VD&a)>^<A
V@));O]V&;LOI=@Y<[,^dQG/8^,G9R>PW-NBP)c18gF[N\dIe;JX1:\??+.[-ENg
--:)I-N2cV)agH8CeET<CAFH3+6:GWe4H@53RXPKN8eJ_,:W0S.#<+D.X?GSgg;G
7G<^SA?IWeFD00#5:K1=JIJ=ZG1@#(fK(.0PEffd>]K&Y<#gI.:0D+>_H?)K<#@+
0=.?g[I^>_0aCdY&^\ff6FDO><,G<UaNW:/Qf&<3^G(5^;d/=:GP#CA(KF0+N75.
(@2TMbBLg4IO0/TeG4>7OIKXE;b\3FgEU/GNSbHFb?6\cO?616-<dD,G?.UWCQ>D
[ITE,B=H#2_Ng3[8^_\-0gOO5>e)bd4JY_=-KM]=<eL,J-?<J)EB^IM9K^[Db@Q?
](d^VR\81#Y&O)F/f\CC25/.),M5W<8egKP;00=eDec1D@R?29\UF/GYJg:DHQe+
f?RY2MK/dK(Dg(Lb>HB4e_Be@7U^#>@&]CPW?fSZKQE>N1^Q)YJ,91Z2d.0K0^9F
]e?[XPU]E5)EUM>e^TVUE3LZL-V0[ffT13[YFUR:EH??007:<?2,b8-dM:[c9@GQ
?=Q20CFPOf>73VQEAdD6a(KZ^(=NAYaH(S.LX^P>VFcL@RYJdd6@g>FJRJ#XUMcK
JX_H8ZI1.UKKB2Y>H?+&VD2,#G?^eFU=2A/>\cgO5H]@Q4+QdUEeV\S-L^/3QXQZ
\BI]bLFJI[2MJ:WFeT49P#5I5gaGJ/7FI-48(DXeNGFWLLcKG+FIA7;g,-[G:E2I
.FV4SC7G?L?LQ7-g<<\Ze9;@Y/[P=/436_#621UTC(#^@6S27SF:@5VUd9e)\[@B
bS)V=<H[LH@BdEZ#If,PR@,JMV^0^0_Y\]-V]?FLI5ZQFAV8f5(IcCJJ8UN_.GEK
>RZK)US63S[,TB<]P/VSIUSP9I@HDW4+C>H_&OJ-:JZfDZaVK-K^T7Le]\R8?4aU
+6WOd6.#fM#B&O?Zd#<ObSYfQHSa+GB<V;-W?;EU0+X0_gfeE8.34HQ1A7:c&Ug1
0?.ggL[DOB[(gN405/))VQTFXgJJ((#3OXVAMdL)FH--PdB=VW?Gd&<?M:(HBM,<
2)A<VKLK48C#4D#f/ZNRXCKA+?G?6LdWX#A<@H;6Q-LPb#+[b9(Rgc;@Ga4Y9031
H.^#:M7\]S9(Q[U2@Y_VV1cZ-E9b?11\dZ/?^5gWPCX#93CHI],[D,L]00(@<8,2
BQLJ<C&,6TbG,_U2L9YM>@dQ/)A8Q6S)MLIBK@XJF:@(,V^+HJd.00^U\J6fW^YN
<^eMM(=B8^JXZ6,+[YV-fe)W:BcN7W?eEGg/W)@F136M74Od[C\2g\@@?DSf:MaS
@RP(>eHA[+52M,c-Z>3^)QcA=,&a4CSDY>8c0&X4GRT4@#C//_e<I]+e7WINJ7\>
T18\9+5122NMUK\/,^Ba\3J/&:[E(^OKP0HXU9:>EHaGfTAF5EL?G0??U8.&,G(e
J@ZSK:;I91/gZQ7?0)=L<#AJ9PMBP9@-XJMZ23TG3Q[4CF&B.YRSMBVK-P)9c28<
;F^YKEG2C(O4EaXbS65JGcMQ5QSWL1L9AXKcB2YC)gT4(FW6\[KX6^a^8_RJ:/_7
V[WTG2\7759QEPV9Q4&XK<bMX,UY0:cHT5V1ZS6Y7W;ILXT9_I1,PY&IdI.FFc1;
9/SR/<>B^?4[L4LGX38GI,[&g@Ua[f=QE7P;1.#O_B4bVFd9MMW^17fIZM?SUbQ9
,bf70T#[K-CMY;Be3^98@H?;P[UV80LOV]Y6I3J@S):XT+dU@G^@6QXQ(OW+Yg]V
MJK.14Y<AY#Mg6M@U^Zd>VOO3cVRgO?BFe.Je\f@aJg9->@#eOBL^Z7L><De.5Xa
6+bc_2J.JGH_V=I92+TK[)Sc^PZ0c6_IH2H.)VXF2Me6=B-OeX+_K=M-P8/EZL.L
QD91aYH39[D4<D?6Cc<_JCXC4_<_54R&-93gZ^W6BR,9e#NZF_3/]+6dX:J,1VC[
F==F\S+8NZ\SM0MB6bZ^Fb^^>c_GdS_1811E;g]2&C_cZG[TDPfV6N)g+H-dR(_)
-b;N\;=?3ULPP(J[E;KO:RaAb.UaEeQJdK1[[ZAdV>#&V2^<W,:4A4MaN:MNHL-G
J+OWe9[<M:aeFBDK-3dcOU\5SU>R.bZ(1L#KdQ&K^?XJ5=WX=QdU\2:,U--39M1W
fJ_bZE>TI)TP/=R8GZGW6DGCR4AK[^LVQ@RW8]7Qc@B4C03IYULW4fd4dHa0(10R
K_dB<D5+4g<?IZ?:]Oc,JE91F-fPa_WYWGA&dZR4A(N0NAYYLfN<)R3^YCff<0Q,
G6&((b9NJ^.HL;D:4XZMEe]F\LZ36=]W::4F:A2.b[c3/M.?.WQ8OX2\K0(3ZJ:[
Nd[>Zd)#HeJG=IS5Y063&/(NBFYKVM]<)I:BS,]ZUR9:1/bH(6adUUe=Ea@eO<>&
]]9Xf_ODT<T.F#f-]3.OK,,H:Q4[6TLR9e.^g)T&8<V2.MNDfEZK8dF6)Q:6CVG8
ZO@^&^B)-G&L<V,#>MFCNC0HSN]A5a\WI0:NDVCJ.2(4GDXZNSb@Z;-0fS4K.L0_
+\<d+2<@:P6JZ]L7gc(]8d.-&L9[GC/VE0Mb97;:YSLO6A^=>a,FPL+:D10D0gZV
1T83RIfB3M<2K7]&PFLK^E^>FUWgg)(;1e-?3EKNAQBbI=-g+&fD?1JYQ^-8+I5^
,GJEa9#e)Ze551YBR)A.D=#IY=Z]UA,)SN=?g,eF64HN3UX#9+J=P-C/X#;dUK=O
HF=W91W&-^a:C]I6B<9LfK)eQ&]QOcMa#;:@K=L6H(G@5&d(LCA-@Z2P]4=a&\aA
E/@X/ZJS_QgM9gabT6A1^Ig.,7FgOPZgBHNZ?9INaa<Q+V)#P]B787S.3S;-Ka5.
;F@SE<UfQ2SPRd.@Z-_A,>>,:\O>/&;4fS..WTK(-U<@4N4CKPH=L5LUdV_&@+UR
0^O4R@b\H)TYdg;A&YSAP4bR3N9LJ.KKO#U:H]P:I9[Y^1O.@-.)^-4L?cec[5aT
UVX5/C3Ze0P:e9Ref?RTDA+4[5ObF89UM9D)X8ONdT1?C&5CU\J@ggd:8-b^dLJf
QO)<aSF)TRTW,J,CC/,.\@:cdZf23CH4UF<R_C-<W7?S4b,@0A3)],OaB;Y\,PNM
;aY2&e9UN#A)&J4V5.EBP^=3Ya+IDKUN(A/+EM1<DB5,_VUg.fMNHXWM-01ZY94J
Rc@H?XNN.#PKJB0OM=97JCgL41eNg6DQ#_XX,V>\9/C)N8_ER3(fDRDXI;(K3a=A
-:EYN#W+&)PeQO0<T,:e3;4e)VBR(?JgNU(&Z4^>\\\)YT/Tg_PCQbC=Z>RN9^(G
AXGGVa7Ka;F/d8NP9(B11U2Q(;#J<[UG=5FD0f^ZGZf6>1TBJ=NfJ2_&RCcK6V3Q
>b<Nb/(_d@[XgKF<9dK],g\HHf2(D6ddZ<S]7VVeLQfY72Za&Z];Yc:6#AC]V3eK
aAZJ5Z)=bI=344(cG?9R-,O3()(Y?(QTFO@A+(3ee7ZK)L3UJ>9#?.00c6ee6VP@
POX:AWQNJfV2>S2[bd\eRcL/1+BYN(@RBV2a2JT.QWZTe:_EY89fO.>\<GVVU]U,
91HN:f?Z1JgJX)E\H=S:2FH#EBdf6YaZ<cG@3]g05f=?UL,2c@3&MI-:IS4>WQd9
2g0cWGPQ7Fb.<)>D=];DI;@G#S0Q]7K]CIMaPZR#WM?4PO.K4a,I.R3CDW@,I_a#
5[E-ZO[E?OW;LdJ]cLeD+\eU>SMK5B//<;eVQ=C=a<g87_1B3EcB-@05[-N]]ZbJ
>[.-CTb;#MTT28_dG8U)[C4,[@64QQ1EUaVC52L-@]\L:N&<_Z5>W<=AEL;@5-=3
>74aI[0_+EQ8>[POIa>>)<.a4S;:>/PI<]#b83P>35ddA5UH+\.7_SWA+f@0>SGN
CL6aTKS8g.7]>LFK>:J3SB&GN5b+31Kb5E<(eC2/I27D6aE.b+M7K^GfY;I0CT-B
E6F3Zg+5K#]fReS:E-S[UP-:>^Nc9>>A)>G/QRe6Z<7K^/&A\c[f)5TNc>TeB#d.
.(#:4W=+FC]A#MQ-_HE,)IO@&Q\^I5F1J1(>#8KQPTaIfN])CfQ@;CJ)DNIeE2^L
^.._Y@dXWIQ>0;@MGOUL\C9ML)&VD0(R.R9K#X^AT+:>8AaPN/NW5]Le]_]fGDV)
I(Geb&G=5G];#R<0(KWMC@L==.IJW?M?F3L8LY1-5fWQP5,^(O/8Y.L6b9f#dZ;A
^eD+?AO?[[M>=BK]CaLRH80[?252f_(>0G;69O/:VSL5631gX9BRc;Z55a^a&0)>
eG,d<,>0H?;SK>9-ZOd9JXF7\:8ZYSX5#@dg/B5G)/70-(ab-8LK2.f=.ZK,:_Rb
F&40J.#9>]]GS0U2KDX;5XH+:(U+JB\@^X5PP9F8b2L>S^@Z<cLWFPZ=RHS?A;g8
+HDCX]5V554UL8&M<4]C[_=Q/>PU>#W1CPQ\>7[60e?=FB?]H;^R=J8+E4<eN#U9
0bS_/1V55[RB)dWAC:_0B[Y/R;1]90S9,8C=b(,=^gM)^)6+@=(:>H#C[=<K#LJ<
7(aIfD#@3LBD00,-5WXB,WJL@EIEc/;&JYe71d1agLLQb..A<Jgf>S6WG39E(X[T
f6-F=g7G)LCJO5&f]P=e?2T&J.>[HZQeI3MeA-=3VVN?RPXD9^IY<._dIP.MRFX@
I&c5+<e7Ue\Z#eC.0OX;f4O<LLV<a+S+5-BY\06PVAOL=7e;8FPZ+T5CP(f#2)3W
H-+8;ESeUdb6&HFRP56^HE5d,T[V;BK_&+K7;VdL9I8GJ:#WY_b.b?RN/acV?D@E
Lf8)]PGD6_f08Q1=?HKBFC-Z2DIFGdaFJbW:QR?e,PN<@\&;3Q>,=]/<[Ub<5]H^
7GNbN+R4D+(KC10fSQ_[/;/63N=b)b<<BEORAWf.gH79f1S=F7(OPB^R:MONf_\R
DOO^NT56g\FN/QF6\7P+AFZe5=VV+Vga::aaA8&=fFWac0)DJY0&D)_e,?fFbV96
H^ZR17B)VAYCgg;)J5OU^[:?6(JX_gN:_Y:^<Z>J09Wag2LdTUL)@gZ:#NV9(gR)
GYC?G#1feIN@:=,:P)7PW(a)5Td[[0XeE1#]L;,FTU#>M1,[4>;_;[<,aJMEaBA-
@35IL)<6,bUd:a;,E4M<75QK3aPY5\_?G48CAQ:1BA7bF(#JC>:4/UZ.+G,ZB?W<
<QcV00FTNKH^1?WRADVdY_INAKC2Z28R)EcAY)=aRN#S)6ZX;7_31[E3XZG^DBV3
(CK(JaebM7B8@8S-R5BQ@=M[@:<ZFU4+EC3,3VXZ7baDDZ-C_@9Lg_1)55P55TLF
d6T1D-O&UL:TE0-N5LM95P51J)@T[1KCB87Q/DGcaUJMXQ(#CO8fXD32OF61B).8
V_JL_EdGCL_WIdb8EMACXX7L6W1.;DD=2#(3ONQOW21:K)=Z[KJW[P](e6=?_:<7
#.dJ4bcG?c)9]@AGR]JP3X(,X_4K1R5Mf297@5K/cYVeO6D<1\/7.aPB3W^=)PQ[
F,-LL.L\9HWU)f5-/3DUGR@.:\6H9Sc\=L1Vb8MQe(_WAT6Z)?(Wc9I)7b65^FYa
<f?0PR(5bGI?FFKW1Me+gO7=9R[5A_#abS3b.\Ta4#EV1g8&O\6LR799cX:+)fT[
0#,7=IN+V@,2=72O(d,>LCdV&8B>LJ@-P9Ef]ZDK/OWO_3]9V5J2K1J]?f^[+[RM
W;:>8-+(R?](7:@bIUH,>]I9W^VGae<;U;:7dM[49J/]dPd9?bM<D5594-Bf.I3]
eON<ZIBBOR,6^M,R(0T_RIBLX\ec]ed_EQ\DYT;MB1=3g?ENW.VRaf_P[GO&,S&8
F:WAd9KH]+N\(d1P1J]B0WAdZ9?Kb#YT?.5]CEg.5eOM_:7-<FR&:IO]L;7\35F,
,OAN@0TNdb/93JLSc;EWLI0F<Q=fLEL<Q_e>YbbID8>AR=6EV<I&)1J(bK0]HJgA
9Ib-<YO6>F(_A^BUUg3SI7:ZI3H#V+5EW(A+N152FKF+?(B@HR95_GY-6[S7F>d:
NU]D\fH5M-+3FF-5IOP:bF0OAZDNPZ9G_X4OOeDYOef5[F)8FJEe7B@IG3f2e6Sf
#g7V@dUG9:c7Q=,5<U-,cFGTbN&gQa&THWXIAe[6;FRL7VHD6/OV0b?=9fbDZA3V
=OUb2B0+(Q/:Fa\UBAbUBBRa-:<3#;N1;NG@\9_AH]MS#3NAFE48N)fcR_\.b)gX
[f^0S:0Ae6R0R8DMG3f/L67D8L5A86d7K-_;\baE5YAX7#7OOY>&7/+?BKAD_>cX
DaJCT]S_bD@9E/eJVIZUL^(1T<<fKC)CC(baN?-YW/POC(V9LN64J=4WR=+Fe1JL
7QGLf#0H>b,5F9dg:.^&0^+E=+1WG;JCBF=VC[5XM>@:P](L#7L9@fOGU3(QP1A5
.M4aBLVZ\KeJa)^P=\<8VgTG[H6X^8)CM.6VDOU,=UeT)C[WV(Dd[aeC3M?W:C(a
P1C&eIf>bT,:CI;KYcT4c)db&d.UZ]&fV&43fdQI5YA+^DAYPV9-@LEUJF@>V.EC
:<[Ec+AcB7H&F7O/ZFAeAbNM@&faVeN_E2e6_(:Z;d#If:g/2M1bG(U7(229]a;Z
Y2]:_9O&g04eIG6>C:V,gXb666Sg6OJOK.[]G>Ye3FPJTPX>X[fLWdPeBKY;Y?9(
S>Q#R9PHYdN03-cU@HW.^ccPYdX[:UZ>PO+CGJGB^1NH\@_I1TLeX=K<L^3DdQYR
J,.^edUYf]?ab-1QQZG;b/M=/gJ8J>ZPbUR8ZZ30-MUdWM)SdYLabd.D#1fU(NQa
T8#9B#+?+MVK:<\#3688(fa&2@G:Jf,USA,gd9,F.17=<K9&.a69>5]ca-KR752[
&I36IVHC3Hb2:T=&186X/52@.R4\VgOASfT])9;+#F.R.@U,d]ASZMGb#c@&&.1F
V4Q)NGS/.@@B#M-4Z]01NP/b-Y)Vfd5P56IK50KNN6dR<MD\.b@)d4I,K)2\?2;(
?ZZg2KG#S:dZ6b6ceL^/9MQ^6,EQ-<Z=JA8N#LB-L]2)7)=RdLbSR/,,QV:IO>?E
&@b08(Xd1e.+gcc1&ENT;4e1.O71_=MFAf3+7Ob/AcLbJ;(X6G<#WE3IQ[#X=ITG
>gZ[@DQ,K5P0:/&S,cF:_T3F_e>N/R#ISYbP1Fa/OA<T1g(RYDR^V/N;TcX&N,>+
H7.=fO+-Qc3dAZ\NB1dWVA1DSVP82K?^M?9M8D60#eg3-Bg7/V9Kbbg_(&e:8T(9
/6[O9Qed1L256^0R[RCEV(>?;]F]#eda^.<JMOE17NZSX[NVJAT=TIE+Dc9/^XJc
C.1;Da.ZX+6(JePG7GONT&5g_?BZg/Y#Qd>[?8:=+6[>9,B@K(-.#(&cC6VNHLKg
(\aTJCb-/DD#7D.Og,BU9O+M=4=C,>,fZ@7Re7@Ka:.Z@^A\BXSA2^e9dCL<QIHO
B/G>67F;;bfHK\Z;NgDFgL[[,T?DC-T(@VgG(/.P&9X#f3)/3#SbN5,KYfFL/X8U
Q?3,HfReV,:G5F><8]\VF<9-VV?9&=PNTF@F_18aUBJRTNHGUCU.HVCZc@I:^APT
7b<&2f,3Zd32K3KAY)ZDVAC_LV8/R[,230M[gUI(9Db\(@@0;QOT.XISW-=;#fO^
(J?0UT>?R>&DWFIe=\^<Pc<EO_N1b/bCGWZ:.Hf33Q)b=GFL]&LWHE5Gc0b(,+/A
7c@8b9TNAa>594D;6[e[VRc.c2a@R)>Bf)K5J?\;YR[f^3/5I41L/>bg_a4HN(5=
M.]V4aAR\<?/7WP\H#5<EY8TD\B=@0M]B?W[MSeUe;4[K9]&NXg+UY5ZOTT@H\9Z
:,-Q>_dY@(BCM]Jg?bO.FGY>6CA[d5J2b]ZaA<de)3TJ&6dWOKNU8&VLT?De-2J1
HSYfBW1:EM_HVN,V3eSUAZ@VD5dGXXOFGdEP0>J-[[<J@#@d#>D?.f6CQ>CXMOR8
ARW)>+g&[-b)):L7b07R420?#6Z3/FM_&DI5+HAW[6]DP-THSc;>Z(c0.Y\JT6D>
PP/ZaSDe2E0QW2.H;Nfa?&U_d\9S=Q<MT.DaB#8(R4)8+0cg1H<./[3+(:Acc_4E
\Td=^?CCM^DNK:@0eEC5RO[Pg?4DO3GEQ+51eTTcMfI:JfaeK]/dFK53B6)9@&C0
9R:O3^0L9V8X1S)U,^VR.E+,5/OT__B<X_JCY=#RNNIK-9>@HRcRf3)Ufa,V2?(3
WUadS?.H]3W5M:;_,C.-B]UbGcP3PZ&(KW/Y5XedE;YfNaJAT98^e2\53f65C]d[
&YSB2O/F28fGVU23=Y#+?=]cU35Q^UR<1]^J6ebR1N_fB$
`endprotected

`protected
NY-ONB1QTeJQX+7.F5^KJe_V8R=YH2FJRLHOMg@Sb;?O5fGC)Y]P+)@/VILeY,J\
@b_P8GIgTI9Q+$
`endprotected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
Q@2K&<BgEJZ/DS#GF>3b0N3Y<:f-J2BCb8c(66fIO)<._dWF?&)S7((Z(=>eC7c/
WEK[U\b@U:81,T_3BZ7SI(#:3Y;<IVLC/B;fUde1gCSAbB636HPAI-TTD,JOQR]1
b<;=a;3De86X-E5]f]S936dN1=]X6@CQV>GW>1[KfVB->XAT.K@B@VJ@&VYdJTEN
@^6CO(=_)\e;?+e5+^.K=/CI2Zf@XLd>;I)]2VfSB.HQ+E4?@[W1&52L8^\#]7?K
be?3#X1M1T_P0UN3JEM+Zc[G&?>)bX\AB(6g]X^<:Lc^Yc,g8I>?8<?&L17=].\:
V3fdaXU-0NX6B0:+YD@g^^ZGQg;c<@R<C9>:ZKT@SdEV>b=-[Y8]5DG[Ne?X6UXX
H3GIYf?)V=M@cJ)#+.-NMY5>4bG,.0>A<XfdCc?bFDR?A]?7TSRC2)N[abdFae2M
KFB61b0B7V[BND9]J]1MFKbf;EG7VMD(J(8I7N72O[04e/YI7&Y3-UTIDIP=,KEF
=cP&X(@H(-FY/a=\(_-^ERMT&?E-J<XOfBCZc=YHgP5DTVI^6HXGPf\SB7[N?)H(
-#6RKW646H)>Y_XbU(G4QBf&=W_PG=QJRBN)\K)dfY4OB#:f,:1>:\)E,:0HbW/_
).?0J.H>4_<@[5>]>>BE#:B/N?##H\44Nf<,fV)6/QIY?;][R.97X/KP9W#VLQWQ
AC7TFC(c_bTa<42feeYbUOBAY.R&U=6\1UeZUA[DC+9B9fQP,EEY4R2a<Ke,(N;b
^SG>^)Y-5:@fVR0:LBAWd@/0#g_O(5N-Y:3;WeL7[M/a2-&Df//V8eK=X+?EEG05
:>cS1\bFO#Te\@7Z8A+E7-QJ@P2a&#>d4e60)?PO&,L<41[691a9DNL8d0/)-\P8
0#(#:,[ZW#[7QX).<3;EVF0aQ[E73&dA]VXMW606eV///-5-;R3ZB&(bKH1(J?=Y
NK6dLJE8]:?YEMV(IdI92E<8HT,f5.Z1XJ1JF;/6[-YP;27JEM/P,^&-e8KA_Q<S
XEYG#4=_&ac>8MK_5B)?=3;D=.5gV?c#[4)/N-geLO_+>=0^&R>O?+A;cY@.LRg@
SQ+<18V=FIC249U94AFeAP^#F-=gIL8^9a-#aK[aJIQOZBVP:ca[GICF-)UCUfGe
e=5Z_KCNZ<S\C#Qb+G:^XEPAMWV\<)U?0O.fe[8YfE,PbgL9fg2gDEC8=G9VC-L?
]#GA+8QJU8(R1UE0XI5efeCMHa:=f?97#^;)A#>/@/>\eX(R0NI3]&-R[[NB:\a.
[0SV@N&YYQ&R:O>W9^E4O\.B&2E>\\g):GaW.39/CG498Df2R2FF=)+cW?XRRWB?
N9PN3KX@+Z7)JB63N)6XJc+g,[QCUTWEUZ9S:(#),@:1NB<<P7<POB[Fg,]PW#CG
:46/M0]6^:2=Z>Yg/<XI]3aUc=RCL[I[fL1,_WSA\cYcKTA0L&+-(4_fED6Ib&Kd
U95G,(0cgfL?]?XDWKV>OE/PE:2Bd:S-4/MgWBJVDV:fE./@PK;9R@P^26T@V8BZ
2>[IT);1A?YL/T?,X,D6;J0Ja)^U<?39;^9Td0BH9FD71a#)486^MK/3_TRMf4L3
]7/<R;K&8YQ(]?<4@U.0E0P4U64NNMG61U-b_@5J+;g5XegQ8W,IL5QDgGd57953
FA-._De79H6X[X>L2]]K:UVB-0O05^8,fE6&/RAB:M,/+40,#+e4U,+&MBMBe)L\
^A?MF]>[8K(-0>Q9:b\f4I+8#H^Q6D[M9=d=Zbf@@=7eVV9;gW)LFT1MMXTd_E57
9&6f5f>8=?N1TbE=2bbb5WBY5g43QYO)6+&8dP298/DMF1AVGX9AM<dP&2.(GO5c
08(BQVbUVH]RJSD=K1C;[IGF\fV+.a;5?/I.=;T,K6),SDQ6JLP,1V_M;9W@ZWKM
N04[/_H>K8=aD:Q&a/80P:?:@=BB0dY3=0f0VWAH;H@::5Od0Pf+M?HLF=]KbfN/
PBHQ68_:A>,;b/&R,7cC]J5,+R]PWN\MR3F?U5d]+4P][=T,^,O.T51KR&28CKW7
N58(68F#KIJ]e/eH#D<H[KZIXUC\P4Dg]<G\NLC&;WHDeY:fGYN))b<+H1d&?I-H
8DU,NZJXWbfTUgfeL0K1@DIF#.6@-<.=XfQc8_:MQb?[USJ1c]Gb9NI94MZRR)/]
75SaLET&36I\A80)/O8MGe.)[G97<@^d[74]V5LPQ8+/0Dd1W#XB7beK<g8DKK33
>fYX\T2OW;]d@GAP<EF&C=:f2O1gJBgCDC=gXFORNEg/]2NdfI2S?g#62A:^P\bK
d>Sa;[dII1E2V#F2dYS^<NH-LJK;FLS=5PN#P<,bWg/847=@Za6QPQaC?N&D[[g5
geY:J#\D,-=b]G\>IcFQ04;28c,5SEd,9@K1_?<g)ddP5+3-,L===e)RYcZDB+LB
2e#/#,,V?6IFagVe6+^@3@YV3;T](<OV/XR>174M?QWegM?5,&Dg:@0@N:G5B^A_
KGOD,0A@8g7?fX2YI184.J4S;;?fb)b1PN10OM/@N>2\/b3((fJTb+Y,,7W<1N\6
f@6JJ9g@B14L/a;8L47;ZUR.8;6g?1KgM17(Z@M?C:faeGXR1\D3DKg=Sc&6#]J-
0efL[P,^I>Yf18&0K,<NbM\^J::#1R;A7UXSR><ZG.,-URdOKPd:JJK9MGY/&&7^
L0gBa.=SZ\2ed7/YgX[&f@MTbYW&BP]]=HD.ADZbOK?:)6VOH[90RE-,:<W<6e6=
;T1Z4PF;JGH@:-=#>0c?4>PQ7BX#EN-0.8O\4->JeWP-VTUL.EZ_e29>N#33N5dJ
<(JC.POC?6F5XN:VW4XO>19D5,Qb^ZgV;O15?E10dKOgYa.9&QTF86-]M+I,8WSX
,4([U?g_B0=/\gNDG3-fC]fP1](@L=GJ<S_@d?Y:]c+L_I.&S&6J?N+C6<@d#0e<
^8)e8&11.V+^L;ePM7[E^(EQIBXPW>+(_SR),9#fE_X(RMb(,;1A/#18S#_JLT-3
O:W#21>LLHAbHeBGH\Mf3^ATD6<[.2L#1K#?g4.J3MUe^7Ke3<^afS5dVWg-=Je]
dZR,ga\1A\M._:1D>DEUMJHF_\V7,/7S5)AKa2_B#b-#2bLYM7g8W/U0G>YV4DMP
QSA3dK+,1S:EC3/bK;+DFf\e0dfHR)4UBR<R;]A@gQb^-V#(0c:Z@:^\6X=[7XP/
&>6+d)f=G+e5[AOY,CRa)/X4aPL.>CN,QZT^ZE/#/@-P=U@65Zc7,#9-dK=:5:Va
(E,.QfRIN1]AfNXM?I)9WE53c[(D2@;AR\H3c-.&9^.4FV\[X^>5:5O04ZQ7PB3N
@,</9EV[G&,G6\#Ed(K^A+/.FMJe5JS(THDI?M3/VB<f]AbOOOV:V>U@^AbcSd6=
4M]LY1W+3CS/CMYgQK]/:Og^]:b4XK]c19DFS?:aW>D+M#QE>KaB81e,[acQg4Jd
6.R2H/?1U.NdOW-Pc6U1+W3E@VG1A-2HFT.T6TIK;1_O9BNWcC\G[:LLIW]RT8?[
5cJVSaaNgN?905J1(;.-UgQVe62aCWdFa.HU=VU\IA2^[T2KeTW?9bYXV6N8QH>-
0CWY_+6LQQXYYdOSUX)UB>7/RZd+(H_&(RN]M5-1A-DB6FeP3Z[a_<#T9I[cL5gL
-1Y>@NM0?PVd(9B#@0E@)3K>?P/JA7,&A[Ia/Aaf7XfF^SC@(KfPRJ23cB]#cFAM
O?^QXKg:6SXBQ\0A)Kd2B;bfFIGW=DQE[QI[X<a+JWI=\_[2?,BZFKH)DP]>@a,:
8TGWLX]A1,7@1:3@7:=T:3BAW5#R7cAeF^5a#[.<ES6X9,L=,WE91CUcF;C),-+4
:1MV59@c)BYa_D-?.&K#dZ-7468Qd#.DQ?;-g&EAKJ/H^L=:cJ:;4aWR;UU5a+)3
>\YA41GGg<G\RB@=^,cfNJRI4.;3I1a4S>5SF80B]_XM<gX4UcTWeNU44HBKL.2+
LO^NC3+c2JZ;^]O<f@TLC\;+I>U58>\g-8ZBMa)H8-baDO8U:=UAUT3A^5OU7,^<
T8C_O.2U,e)a5F9M-fE-8(LIbEN9-&FWCcXKg7TV8DZAIT/LS@KY80Ca/WM?Lc,-
#QWL68:JR49KE^TJ?X7TDGeGQI^:D3I/K[LDa]7cTWYLDE1B(\FALaT0TSI6GKDW
;e/=I[AcQ[3.MG[).+_K;Y>(/>O#WC0/8d2PO=PBL_)La5V1C<8a,[RJA9SK7Y6T
]2Y71DIX3E^dSAaDO[01[EKd1S?2_S(YU]IeC:;[Z>bWFS3QGL?\JTgI+7WB_7G1
,L.@TN^FT3cO=QC^W3@M&M;_R<DaT<E[-:O&-2NZg;FB:cH#XAge7.]cTYP>d)7T
;.ZR?(5[+fTfZ3_fQ>Q>7ON]BEI+ABY/8P@&U==>Q.)A:H=^>egHQ:TFG072FgIK
Xf.6_&Le0;QQ;T9cUS>K;3<b163OHF&KT,+.@LI7>1<EY;C.-(:\H2,6efA:R6eK
6&Q22a)4I<R_F3b-K+eT<B)/4]gMNffYR&0G==?D_C:KL13AA?9,E53(Y7J_8Ic,
<FRd5X8dGHA,CfWE3N1[IR)GB/f?FDC08B5&(/C.W1E756ZEX^FLX)dDa@-_dT&O
-Z+P2LFX[<C[;&)S]A3J_Z2[=)@Z[\aD?N@Fcd]a]C7HQ()F6)<4+LI]+&I0XbMM
/=^M+^Rc-QC4,ZK]AY/BfS+V(c._WTT6ZR>6gGP6[V1Y:0D7bBf7Y6JKH?_H)aFW
a&;V=_HcDUDKD=;Ee_2eCW:O(ZY6_4,X>8(I^9\VJJI)B6-d=51G,fPS.6JVJd_:
4EgALL;6=.JYBN9Qc((E>78I)>bUY&IaeE-186RJ^W[(6bD2<,ZV2WVM.5SOS>;3
4)CKaOgB&a=Ja[[g2GZc224ed;OGgeFJMNSe+2e7c6168#-&,@AQGdFKbTgX>(L<
\6Q.F8e(-1D.9D)d1IVQ+2@EGE(,F?QMc4R/d?JNLfYW[<SD&662[KJ/90ePIgZ/
Z@UdB<P;<G(R/V-9f_A4=BVAT^]8,RHFNL<DB53_W(ICUCKNAbCSEU75OV,@=eEE
O3?TAf[,6>#cGgc4TdQZTFPC84O^99682<6dc1-?a4(PMfU(+[9=/AZA(.<9HO6_
cUJNa@d[(FMKW<9-OM<9NC_8b_S<bWYQIa]/W_,#DN[TNTH5ZP&8OESbb?<-8\?5
99Sd;Mf2-<O)L:Y7<@E&a3AESL;)f2#D<H2UW\VM]Y3(fA<123;]8YAMc\GC\)._
Wa3RED-bUCYB]F#+BfcC62/G<f/)8Q2@ECbH9I+-0fa>cRYVK2J+BS],@QF@@AD(
b5TCI0P+=>Fa:#9&]CE>9\&A#X@4cOQK,d;7Ef1REQW#)5fG\ZcHC7R-Zb7(W8##
S3)/M8X7^?_C-^4BYbX)WLRd:eceaE_5dVA/@/4-Wd:)QbR;4#S/9FQ9<(PQAJXQ
a)V__US_:Y>^4S8OLfA7U6fg.2EN.508aEK@a3,^(M)U]#C)?6R,IRU/.DEKH2U6
<^#WDg/(YL?OC2aJSdH4/5JWXJ&dCcc-;YcOG,FGD.R7c62<8GX[)3(SAER8S-HZ
K?V5^f7+3(_(?E/6F(g/gC-Tdb2G+^S;9PdZ7C)e>.&5&7^Ee^=_W8V\(a_\S/F@
\B@5-,_Uf9+#5MZU5E)]^B)(SKTdWbHRSB_M3E&]>&B1Eb79TfIPJ@g&F>SO8#W1
E=Df;0?]Y(c^Q9E:P(+T@P7Z4#L=XCEJG]WUfZBP.aD#P:eNc)+<?0O3CBRH2BMD
?NFV,#(^.>(L(DY;.JW4EG>11>gGQ:9fX4:fe&#<758,S2M:3C/]?XOF#6;62f,Q
c?CHGOQUL2<P-U(AX&(MbKMI4^B9IeM+4S3LaPY\9M^ceJgZN-B8\K[Ee7E5QB9C
7C>,])a4FYSQJ??>Q;8FN[6WI:Z>?1P-+\5BU[A=V^fcKDgA]V_C2L6VCZWA@Y(J
@XS)8DM_?dK7K8+/7(^.=E&SGE80&2M?;9J\SOG\c@G]f/\AC0WXaEe>;I[.J)7I
75]FHfU(5\3>4OE6XU)1)=(IR<X-6GgH+=a79@g_^6&(6CP4Z&OHQP\LXf<2=Z2)
NRM3[6#]FdVcdQ&DP-^Ra>(G=/@U47EbVVK1[PX4/356=6&I?J&4a,-^#[R7.>S@
,PaTc6f^)0XH7\9g9WU977(+:fIY_M>(3Wa(\:0\=_W>>_Y80c:AE;7g.QMW@\.#
f&(L?394./RSIZ79OM1??X].X\X-^SA^3LP2N8SNI]9QK=LKK_#BO[S0)b_^6c.,
^(NF6F51^5A=.P/YUU]4W&SU9YWP1G==\A#Z=U(]S/+J4ZDUZ]N(^,\.MH:I6aW3
:8Ye_83B_J&6=_FW#/P/b)@af6UP,>HeKRH[:NW/PNXf6_2?]AS9c&E&RI)RHPca
RG:/13-58RT6HRJ&?D/6LcJ89QSK59;^SSe/OAI=_])H;;ZZP\YTHL4ME5PWWVPB
F0<L/]5(H6PBJ>FF^ZBJE&OG\>E^ggSZ0Y][7(WU<(WR,CbHQ;=0YYHL9.RMaDGN
93LJaTFJ^:>##J5,O7(Ig=VdW<cZB;cM:HSE]4(J:P[:I/Y<V;:\\M=V^\@?91g/
5LCJ;QGW&FgXQ5\[Mfec]8J\d7V^);WK/I<Ng\\a;a5YJ[eRQ(XAG_&=<ZVP<Y7f
T4aRK,NaI3IT#46W3Ye3+NUg;PHgbMQ(T#c<e^/=cXBU^2T\CQ.;H_S.FV,/1ZeW
[C.J74N/=..TI/gLWBM-Sbd@#.Z981bXPYf)gE4AM6^G^[fGW29#fV&?bC^4LCTR
HbdHKEA8QH4b[XWV0C^?\<,X5NLG/bP3bHUSd(#B^;78BdP(2#6FcNZKM(=dI5O6
?I9L3VBV/3NOEGY..YO9TXW_1Ff,3E(b;AQ=<?GB>DdNdX4^-S:Vb2.<cWF.4ecX
KW3V\g)19N9QF6[/#;]HY/8#5?3eH(c3D?E67(IP?ZJRMd.B7^FPWcCH]/9d&EGK
:[][<C&?M(g93O(c\T7[1G;A4</PM:4e_RM;CFc2M+H>aKR]?^gX7CU>=FWc?EXF
#H?Me54B4WB-@]c6<eW^e8BN]^VWT3WCX[#,>ID@fc)DX2VHE7MbEWYb>0YIYC^3
31NPD5;NI:_CPM#1f9[0U-VKJ=(K[eVE0.]Y[VF,68J37Wf?g+fbC[=,bFaOUUVM
60:g:K=dWSH8G?@@]H#46L(Za(1IW>:e1<H?&,/2,I6-A7+Tc.A]aKD<3#1Y_U_:
]]Q_/CEZTa683CXW]?B+5ac05a.??JcBK6D_XcSVBf^^0_;=R21Ta>4J?/@A4-eI
D8R.D+@?ZGG@33@Ud?@&V<J2L&9-\=UG1#XB8Z>-GMf[LZRP5<7AX7X]=gfKFU1=
/6eE)2HIR<1&cTI?1.^9,&A]O.D->N?&d)M(a#>KROY)S#^,L&@L;J<d7?c(?2O8
RVDK9GOcQbV1=&EIFI(bc-c(@DE#Q@ReLUNUf.7,7=f_GNV8Ea>:,P(OR53,U5fI
DH-fSR:D8GR0TAfK-61U7/T[7H>F5IaWe&[e#^1N?U1(K#_(:^6?KEFLH[C_agA6
#Uf^Cc#6XfNaCe743eLQ)CgZ(V1?9C2D;96EF4)Udf&FY=GM7g?<\QDU(.PI9__D
ZXc8(b/cV_7P.6M-XcQRH;N=/2M3A>][K<E2E+E>9&AOC+38X/YFY@@RO4FAGFW?
H6Z6KH<&\VD,bU6B/Z3Cc2bI^7(+;)YHO>XQ\/:[;be/<a[(=@6UDV)M6_>3M[@[
_^:&^9VY4K#4&0>NHGTVUd\?g.[\@7LeK?1KL=#6PGJdV1c4cF1ccC9-U)3802OB
NQ.TO9Z[:?#UCX<&D&3LIJ>_gAB5CT?5T^aO:>GgeJ>(8+LG3>?O>A.b81L2-J/7
<&#aTJc7]GE]WD76S122QedgN]=)-acKH:UF_[cF?-Jc8:0I)aUGMANcP.A_b?J<
A@I2,,>1DV>c.A=6c9N^,6G#CVdZd?453:2RSbWB--O-AB=d.^P/HD6CY4?[BC/,
/SOKKSDb)YL/^c,2=TDVIL)Y+@aUacOc_O2J2-J#0#:<DCD\cc7KO7>54?HP::V@
A2YD0;#8PNL5fC@JXeW/+KUfc#H;ZFXB9A>:1URM,ZJUBe8JfKDYNQ5J\(MLZ//Z
^=BJ/\b76f;3\))QW4X6TVHHg(Z0?AS>B5#?aDLSUYC7-Y_bN50CEa/0-3P:#A57
(4S&.4e>SQD\a<dQ7]>_a=]1Q,Te?OUDJ+(/T5e8e@@C_DBS_3-eLL_f>UZ2G:Z9
6eG0:P)5E7:gE\P.NYH2Q13=[;:LAIZD7#Z4FaMYY[Nf?9b1b34C,;Ja]@<G+UG(
<BFS-b(Cb[O8BJXDINF8Q<8C?C+(HNO^+eDJ2069M(V4caAZb9)-_U1+c[e^_aYJ
8;dD1MN[Jf3M:&d?+>2]^#J(48ZV@4GKUb9&gd?O2X6Cc1M<G@7J(c]dLb(6d6Z4
T03?g[VANVG>f(W0.d5.#[25WYL6#3/bLFd^#OND?.H5c9a+d(.I-M=/<]MUIMZ(
\56@R;;(]DX3c+OZH.&Q[]AeC>GIW.fF\Ee=42c0>7<<?fc@M7W[8?]:MD&\+U8H
]OUGY\aHb51]Uef5f(/WEH8,+\L..[6FYPGaN=/38X@3FQFKb&EEH03dQ]#H(aT@
55<Ie[>V#d]/+/BJ6U#6441WGXLX,[>b/[UC/eS7J;g@>c((5&>H?G[XV6N/1Mb.
@\E>827EO603:EKf9BHIe1NJS?V]a&2bBb2G5&[+=H)Y0HHd4&\9QOJP_bd6+S[4
E>4-6X\3BW42f.K8W75cFH/Z]L8<#UW/M=E=;11][d+O_OLCSWVeN^<\W/OZY:>2
/F&:M@&E/0UH2Q=<YM1&8W7P[7/.0Ma_]MA:2f[<2E;SQd8&<^/[CD[=K-SCH(e2
N(3OCU=;3>e]VLRM],NP+&d8_4IK533VK]e3DB(&(&-7&Rd>T>BL\=&Y>I=;]V#D
&CgY\=\4<.7S[I39&6,00SS,1D#;XY_IAbP:DJ7IN3ETAEU\KV;XV5S&[cB0NR_(
[4]5F/R2(\\&b\gGeS/Q-W^MKWEd(6OQ/<BO;,<QBKP;AKT6\R](1Ia_V\DJR:9H
&(2VG76<K0c)T7+ePB\bLK44UY(8g3(BfULGTLc06JF9H7B_(BgJcVC@07E.:+:e
E@G<,Og<^&GD0Z8Q-g@c96f9O4+ZB+TRL//Td78442d(a.=H_7MX\Uf^^Pa(&A-Y
K2J/TX3_2I+R;FZWSY;;)57Ac-F\F:APIg,NX&7Abg;3316OGdWdQ]f7@_4B8b[3
Z)2G?/5bH)M77G1Z;I@J[@WZ#.fM5-J;L@I<Y5TPV/P@H\]L+#-e=AcAGTQ]<#C#
]T&)E:=&^V6bg()dg#;[?XL8T.F7(d&)I1g&@>C;+2^]eWa@_fX:0T7P7(OZ8+_0
5V_O33YCQ=</N50_DJfcgNH;?J7XS6cHfQUU#8JNSTb[T2_]U7OS4:[IIfC_bE9^
gV1\B913,Z<4JH6TO/CZD93/3349d(a([=YgCP@f-dXD,:J^B2/^D3c9R8^/3JOD
:N^ZbABdPKC6dVUVFO=S&7gGSVa,/-]2YPC9KbT@6J1aG@T>H?O,Z4<g4D71RVT[
/L[+<>-??NNBdEFSPX[WGRaL[=0NC[_b9H5aO-9YDf\gaLf+ABK<5I<7fZ\Cb&X6
@>E3]^M2a[JfYZBTPQ>^/8#56L#BgQ&/O?gD1eC<e^f]H;;1;W(:TY;^0/7RIFLL
MM=f0MfE50(.3=XI29VHQ+NOW]&AS9:(W?_\YSGO_(aEe\aOP_X;-3>TCMbNT@<>
gOKE-5[V89O30Xb>:KHP9HFZ[KHaLaI?Z,bROK@&<(73/G&)eYH]#d3a8]aH>Y>S
.HaE,M,#X0C;DQP(@VR#LSbIBN(L0R81eN=e5#UH[e@IET6G(HVUfE4D<>?e+We=
]2ZSOBRIdG&FWEVU#[/55c(DK@S(.gTJJ9F:d;?B9CXad:Qc<8ZL(;FUNP>^_D9G
7gOfKVEd;_WI<OQ,AW>TX=b@6FgS\LQUF]gX0Ge2SaO8MfM0TZ5/N<6g#/7VGGfS
FcRId]F=PE\U.c,O.Y6Q,JOC3#DG;Y:K.,N6?@)(0KT?TGB_AV[?N?W4YG@N,aG(
V:d+XD_?#/MZB8:g#&5G(9C;&a0]/AJ^bb3M8\Y03Cc.W/JB(<gR9)]CIP,00f;K
RDS0MZB[HCRQ&R:Y3PZEYECH\a-=9WP?PT#@-,8JIQNCbIJ<9KNN.fL<[A9I8)g>
0MCBbdZa0S)JcL=QC;Q^_9J<<.379LM44#=FAT&g3gT;H[Lb3f]OC+6OI0_4eT[3
@AHe7#:3:NcF.8Xb703T\YRNg9;0aR8_JQ[)R#.KIM4A]+RU+YHGOFOB>d4YSaBO
f)21g/+_\e,=HZR?^=?TEYR8:M>;Q+3C0dDbG?ReWdH0JNZ+52-:8F8?1^)S]AP:
FU-1)B2I#6_381NJ#]7[1K=0.>@5B<H^:GaF,08LPfUO9X_+^eI?4EWBOPW<K80(
CL5]_[S,]bP::L3]da2fUQ_TE,QJ3:\+YAg/g:C<LHJ#M?VLZC_ea&S>S?@a@Qd5
0/BNYVA]fU5HKPDS6Y2JXaR?0,(:fe/b:5RN]Tb;@E@\dIQdSabdSXFVRTP.33LQ
2P\fEeI(#5JfRZ9P)MAQ)\?](7fGV8b\:#,/<;Of?W9HK<X]_+^WLD5cQJ_M>b5H
M+U9Y><LTTf=bSIY_9(7dK;Pa?OOK]10M:c1&2XP-dAP\LR)9CU<B/W9R\;B7JW1
[-6AFeM?R7.3G#4T;>?]TL,H&EZ8Bc4/C0Wa[TSL)^Z9[K-5R4GY_IJcU2ReMU?]
[/(7YF#B9VE,aA8VPW.d=2^:]T_H8F-\bMLWWDcRbUBFU^<S?:F&a(<c6O>Ta/RU
;XC)@RQ^ZQ[;f\MSABc@@=R.UT:)N6FdKCD7=Z2J12IH8Nc(&H=[70a/K8\JT]]6
T)TbQF<WL^5)^]-B1#,N.E5P&J.(NCD9_M-FF+KBfTV^[<:@IG5&]7WL[?[VNLW?
]H2.CE]_4RU)JFP=Y?c8K7:AND4L=7YfJ&Tb(/(WYT#)bI(Z4a>)>@aYZU-&Pf4-
.Q4S#188H8f-]5Ya\^&2:[c_aeH@D@;J:68>-fG>G?W#<3;&S\c&[\YEP6K:C;E_
ga30/UIBG1W59eTGgbJ^>L^1^MddF)&/ONAIUT+gF:HCb_NFJX[-Ue@IGEMB4^1#
AZ9/gNQPe6U5<+?B96HcD:)KU9/UEIM;VK_12[<CQHJ2Da23:<;WZ>bdSJ/P:K5O
M+U&(]KKGJ-A,_dS)_:2\g@FIKW3KUMS^ceCe659N]Gfa]5&b2eX;,(eQ.72^8<T
a]U#?(ZGCg0H]JP9AE]?fU-]e]S;dB=,BO;N>NF^_2C^a+A4d+>LbXRC]EG&;9[a
f=f5@8&4O_BCB/\C^g;,KV,L+/OR&bOgWG_HF2eMBF3#,WLG7MK(X=>1OL0JA.VL
F91f-1[B9(GU>deBbOBUEUE6+.MZ9>C.AOK\I0-X/W=GU72Dd2M^^Q_L&\PRAT9@
\:XUC2<30[FfJ9:EWb#=5fTZNKE\Vb_[SgD(WPa/JR+#acQ[eE7C2M-D[XCOfcX#
L;0f30DQa]DJG81UTM[e[,V8Z/=@9?[J)=L?I0#&6;T=(6L88;0KU;Y/?NTD4fIg
/?@Z)1_5?+^e(-V8)WYePc=H(0a(R(Nb5X)dHSE2e3F4bW;NcCd:J537&W_8e-c,
LeRUYVMX<M/CIaZ:_H(dM:?+2^(#gSF+,d8.McFf3d-^YHFY2_N]F+&0.A\_K[ZC
4,YRSaP3OUI.)9+?P-5?9AVadgTc1?9M@b\XK48X_4)1feQe?gM.e5];aA1#Df7Q
b;+4/AJ\9Me<^>[^8U<J;B-HAIPI6EYI@SP5/(P:7WVBcJB8BGG#db?-c&>PHe6[
&479(JA5+Yg3?&5]>I1]U6O5[(9SS7&UU4ZZT&X8[CHYL_^X-=7RWPTP_I,-\ADY
=:RZ@N[QgLLV,AVc8be(E9&b0^)QIEPUZDUEb+]g1:_<aQ+Nd^N>T_TJ(AB;:+EC
8+VdJ[b2Og)@TE0C2b^0E#MN>YGNX&TDVH?]/KD7/,QC2.0CC5gcg:(R.R\2<dS+
@#dJ1],#(4e4]W?E^ET+X&\+P^=5\5gQK25#]3Z@<;Eg7>PO+B4c5JF/YfMPJWZd
&XODZZdTH]O:+<;\@L@O#N1CAc/(&L_8e<LC/X+M(08URY2J2\,KOKYb72d2R8cZ
&7K]BM>CRSXVNMEFR6R4#Mc<ZT#-=,JR;bM4OQ.8[:W@e3+..UTE1QS0XJb\bY+J
]EJfAK@/P,-X7W?W.+-^TWH@YC\YYZOD[T@g-VJf4Ld4[b921>aR/YSeV^=\O?dT
=1TGDG3ZHbPF1,S6XCWcIdCB4[-7TDOMN8I?4[ZU:PU_&I&C6e0I5@UT4H74\N5-
W:dSA,Q_7ZZB,G(JDEX-#;67PQ-;)gG:,6OCWeS1HR+>L?gF\]6RS?.b.;]1J>B>
OEX=2)A:EEBRI0aV.cW;L&Y8D(?8R&X47;#=BMM2e4@1SM;+V.-P[2P1TYW0XG<-
UZI1<USBWV>TT,,.4YfBG49;WaSQ>a505N7&7eC(([0+?cGUGcP8bCd1XZKgYFJD
D.:(6&[84X;.D]G+/FE)a_660c/(cU6;,aKdLOfg+AEBEHG[]&b_BFWX:Y-#f]SW
F+O\/c=b(L#Ee5]VM+8OLQ&AQ93>K&Z0J[PNe==#=FS=BK))OgAgO<gY<6=e2>fQ
;5@[#M\,=@#S)#T&EQJ2WRH@7/;DRgECE=:A[D9]:JMC7]gQ#9:G6D[Y32Hf7R@Z
?J1P<@ZF8YD+?VZ,ZTREM]M4=RXG3NbfOID.H2M\KF6S0;eQ\)ceQ(EJ.8Fc+XgM
]]IKBDQIUHUeV0Y<>P#dS?U_=GRMDefRD7bOV:49NeF,1a6,BSB2g\aD#AdeD/+[
HW1&W/_RXZKXa5=8#=[EF[C\1WP]QQ=.FE#\Y]G;S96G\I+IEG6gX+F))2/d_PUW
7Y)4<_#T5)gc+Tb7V.BcACK]1bI)JT^M^=JE2IJ(SKM7@6eW1=Mc]f;L+1=Dc3VJ
4=LTeT:MJ\P&?,CeBF);^A&+(0MRdZ=^V0\aW8WBAY<PDZ\b<X8<N]J1VLZ+b+WX
W2DgX]H95,1?.A09X80OV2K__Sd6fPIHBKO+#R6IRR=T^-67TV=f2dID@V_>db/:
c/)LbUaHBL5GTFX^?TgR_N2_(K._A\gW@[(^gX3gFdgF32/X\QeZ:<528)E/:8(#
f-)EDH?:F5SVGf@-F)65b>fTe7I,BQIRC=FE_(ZF0[LA&>+bIdPULbR>&X@/>+/5
@cd0A&\Ec(I9g>dB@+4(@b^>97L;-E@G12K;7Jd&.B<7W+IFSX,?7E[3cVQN6US#
GdPJVG7SV)B6a,?;S4:a3M84_^A.YY]:KN6:fFcBE_XKM.9+ET[a<W+6U@M<5DCV
HP^IIZ:]&fN\OO5@SQ3F#O51BHNC;8G?8.aWa,&FD3,G:^8/3RE]^0G,C.E;[C/^
&eA;0c+X@JPIc;SB=8WPEB=#HcfOgV#2=GR7R1g56T/OI0U3+&TRS\7;JA)gGALc
N4)#]PSXQ-W#MZ]>@9VgG,VgE?U&9IRcU/;WY94JgcTUGg63BG+OXAeN1c,ME/7X
a_QCF^dHDW8_9DS[H=MWgBJD,1Q2SIC\1IdgLga)+9dZN4LZ+3RAHaFfBNQXUY7P
K@JD+^H+<7CSS>U@6:W,=0B2/5eAKK6Y@C.f?&WZ/ENKT+6aaA(G]7/+<&=OZD?C
ALHQ:\:8@-<eL=;Z_.:B?60V,EK>+W/S31<=?<_&S#\g(C&/;C[/&TBEPIf9fdE-
[R(H-;7&M]@+380,43Ja8a2F7Kebc+]_eg8RB^=?C5R8)KF&>F&cIPE4C:9D&E(D
gdf8LP.<&EZF\2&Z:&/+=P-[^_fN_Bd+0(Y-Y3+LfA39-V;a-9gVV9N8K4N(G?<(
>#U\0dC]ReVeD@AKdANY2(C6Q9=2#C3:_J)O,6NWM_3@^E[2FBYdG0ND1b<gQ/,(
d_X2bNN79a:a=TYDIfV<F]:CM/9K=6c[8b31(f@\aJDZ(]ZM+AW.PP;JL=JaDW;I
T=&bgUA9=D=:d;2WA7))N:.Se_--&<b-=.=A0_C1dFQC;9d.VeK&e,0.+O&0K]>+
J&Uga2f+#?<SY))9-A]^MBXd65b0F-3KDKfP)-:MBV5C@ZCQf1?1PWd-bPd@Ec./
K4VF.\=GUX0IN&M&ce2_eJ.fO759L5._H+VH_(8VY@8)Y_/L>N2)V7:d6BL5X\5B
L08A=G..:VN+<+;70aOGN#[(2=]_>2;WX5;\_4J>K^QTN\JP-#3Q4a2cKZ?-[&B@
VBd)H9BQ.aQd.d1O/+.DPQOMP&8T#1YB/eJN]Ce)P942H73T2;@MeIV_\fY29IZ7
0Sf1?a[P;GcSZ1R=IM>G&7^A77D@PCZ-bZ-3H#d(?8;OID56..#Fb0S/Q\(]eFEd
:?S.U9)Oe,UO<?]U+L^KK;f^1)9fL95.:bVDM-D_586PU(_G[KYA3\^_9@X;JTS_
FWKFUf1=SAUP[BdRLNLTMZ]OcOE18^>O&Pg[8b6+M,XCXO@(GB\/6;f4g2]aMZ6a
>719/4]<5#I?bd(.:C#=U0;WRWPa\-(aMea_0EH23Q+GOI64C.-:HQ^SUfaX3<F\
HVJIT_TCeeHB]_[<K[^OHa=[<cW/3f(X.fg@=-75D?N)FR#cCH0[NJ(?D8EZ2\S\
J[[;A8f84;FLD2QT(=&:Z(6f/=QQ0LcEG6^,eF3#VTP@<7U<0RZ;(;&[]AgW3.KO
IGcNVfg_LHA:9a^,X07?_.C=g2Q?_7Of3_I+?Yc/4a;.abOI08(:gP:Id&HcMe[I
R/aX>f13U&2QONI_GPDAc>&V8e1^KdH?UE#6GW05Pg=B3+\]F1L.[V;3YDgWbK55
7]+GcUC9cH^QQS3?e@:d#LHOf5L:X:4R^S)32Ge7Ee3ILPDE5QDA\N7\Tf7EBACO
FE=_,P_[O#@H;M,D^JL#DL+<E67gUcGWPJe=8deYGcg(13IBHB3(+g]b]81-_3Uf
I5P7ZMN+Y3Lb>ac0<T<4.Dd[;_d/c6e)H-IUJ>O.-_?4N6-Z1UV+Q+9P&=I:J8-E
H>T7/@,MGb)D,#E2U4^_^=(&\8/^&6],-DaKgUX9QS_Md<CHM6dd.cX6U]_/TQY8
bXT53UcV7W73E>FHXd+9/EB,]H(Oa\@Nd/]75^UP):?5?4EOZXK+(D.+AO5&O(A3
;bL@:@Z#W&@/;^/0F#N?FZ6=K1:@gTSg[Ve/48HX>4:CI7(&&bN+BTGg6JM>:H(@
/;VTN>V+a&1?\/d.VXSd.a964P(aIU:DZ=)JM-Lc8J@_:7Ma3SVX>A^ZEEBK9/^^
2;1QM1\e)CWg@-0YW<7DSVV2Qb4/?eP5:@P>L4X29)M_LODM5C5O9ZD#,b&]SK_A
S^=d.;<H;2aL&_?LGW4,D\fY?H-5a6g;\fZ\FDVFbXHDZ:;-A]&.:1.86?<NgcAU
,=GBMZ7PJGCgBX)6S4UN[:GMee9?XO/SHAG3-CY;LDg_a&UXYJE85I+OfUaNX9[Q
-f1X57.^=]c\S)CYd7Y/JDTMg,A-V9IKFXG:63^GD_KC1H<ebX;Qa9U74ZJJKG:Z
_6b9_cB;3ZK3@->5WPV-V6(TGII@G3:,;->.&J.eIZ7(H4/)K430<NP\;7>7b&^-
>JZeHG;KgYd3,$
`endprotected

        `protected
P8eG5U+TX@PB.F\?Vg]0dRgA+TYV&NPV1@d,c<2fSC^EfMKO3#P&7)1d[W1YE_ZY
I-<e/46:f0B^/S5KD\CEPN\gMNGPL,?=f8d0aJ&U)>(DfeU8J7PCW1VP7NePYacX
E8W:W@.J/ZeVAbVS_IXXI2A]:@FB(Yd7,X,4^IG,&Q/Y6^/G6.UZG&R0EA0V#A,B
_&#Oe-4e_4BQbZ#bdLg&O:@7;:I])Y=>21@(E(>ZfY@OJ/PMcQ8_,9#]).>@1R,.
dZ_.3>)<GC@Q)$
`endprotected

        //vcs_lic_vip_protect
          `protected
L,^I[V+RBRd,8XW7\U2A:aRMMBP9PJgCPFVK28M=O)E6L)B=<-f]5(5fAcc/K<\W
L.LBY<B:IVP34;)_SX=#A.]8Vg_B:+)I/gJOf&FF_cD_&P<ag2_??MG@@eW=L0=S
6c\IUQ-@^YQV^]-fZ[4fMd(F)V&BIF>=@;FS/;AMYeGW:<cEL99DUB:T_:8FG:2A
K>9[TYA>/)/Hf=?C_Z;8&c:Ob3JWVA,QQ]XKQOGE;H:eSFH\2f@YWBY1Y4^&>fGH
D[d2g1^CIeIP0P^+#cRdef0[V8a5JVE5@DX@Y-g4&MP7IN&M7c#M?a&XRZUO)A-X
N1GMI\LAB>PeC\[=(5^JW(U#,DEL6>(M:]219V_g#3?]WLL^ZI5AXGUY1M8X2IF0
1^QL1XYVVc^IbdMMALb_E\W,P.T(Ld]8-:ZXbNA[e:J>Z[A\01Q1f]7HYI.XLe6a
eHdCZX6ag#-\FceCgae]O_XKG#;3L[;0M:O<1IdD^2#?Z4_7CfO6NY.D>F3-;SQf
Z5GOf3[LECI:-U(KaUe[g_S83O)6W1b7Q?dIc)&UQ=7=;57VcSK][Z[+1fCMWg<;
+]0MU][P(<;c)<5,(K4+]VV[O@:c=+Z)M:KKgC?9b>(:?Qf^Ec&I]XQZ72&A9D=2
#+>c1I791,\@aNdPJUA.F:2/@9YbC+?_5T0,[6)Q>^0QRSZc(BeYB+BCK-8LKB^a
97,)g,P?eZE<TLYFPZ(9^Z^V^XEC\VKQR0)F39>OM87=MWQEFTddR;<gUCT2cQ9R
cDN8XTSTb@)K\R313gBXKM[cP&J>BZee&U_R[XT42C(?<]7AQYDgF4dfP.2gd>G^
VgOOR\2G&?UU7,ZJ)W<+ZGWZGa\)QDVg_E]C+#P[.&XC@>HW@&W0FU(@\OAYbJC=
T-Nf4)>)ARD09)H.8d?C<4-B;3e+UWPT=\P@.9b7+NN?^gd\d]U[0B=ICYP5a915
f;]f?>-,ZAJXaCTNAd9^bM6UL@YUfP_)c^+PQ1^IbIZ8J&/EZNPU(HEf>BZDG3_c
eHc4g0??dV5+&QEgZ3Q,AQ<I-eIY2R_d)bQ1]-<U+#dT>c(f=Z.?1P;&K<@)D,K)
85?/6e4/</fT0(O<5&0D)+?7CL4SFP5DI,+.&=XD76VVb0=KX(Y9WF<QM#SU5]H4
Mfd:?R42+BC(&g3D3;RVbN;6T^TJ@SLFO_V?]0N8\e&M-\gROVE2RaG4VVVdL),H
S&a/c.]/\LFDF=@_a#,E95E>C8ITRg<UL0F6SY.S6JUC))R]JeO=P>d^dfV<[0.N
#KP@d,Be;W]&Df;P0X<a=HEBd_Q<&._gD&g)H82PT-egEW_\K&&X=?:9[04PTG?[
Z[b<-&g1)O9\8Na_[B@[]eX:_=a.>aQOXA0>-9:/I>c?<WRRC0YV&KB+G3^K]4K6
8e11@]<WcFM.SAZ[)eE@P7[#];^?^Y2)\-<bZ5b-V)QE\f-J(M7P\f,G88FV2=\]
8,aNZa2@1_:;SeI/UM7H4SG;/K5QPHF]-WKPbM8W)D52f1NB-&KTe:C-RMXD62(U
5\9V+M3GCbJ;P(D[^@A<G:]bE8LQ62EICd,(<4(cBN^Q\P60QFAHBZ2C-PO(UABH
^fPW,T_WR0U0K/eJ(F=4+@O.WVN>FL1E+U1CM<E#0aK[ac.f(KR41,?gR_Y_(-F[
O(^.AX/,3/d1O(8-8O\L4G]5g821]cS]6HFLed<TZS_Q_J+[-gA]M&8He9)<+Y\8
?^:^J/&53A]GT9M>/YV_Pd\CW;D4FM)M^(NEbSO2/ZG-dQYOQ1UbD(L:=V)./O0M
WWBG9#g[.(:N&e5f;eReaTN=GI()/EOQF,86)_8)V+gMRGO_Xb.0]CDD#W+K6A.V
a1.C5^BUTDG^WO&X+Zc)e6Ff2A@3(4ZMW?/H;76@.NE+\g25Y&5N+M04>.8UN+#<
0aHP68O/03PbPIGN\&<#,Y-ZA[-@_SKc&U0LBC]&B0D=B_8&aSH#a>GWeAS_J)WP
S:&@A:2.;1aCIS3>ZY^B.1PYf+N#ZcfG.TaC2W&^E?O5OSe)U(JAcZ0YU\VCL<S<
TP/W=Ce6X37)0FR:Mc2D;+L[6Y73(>gQaQ@>A?KKUe^1(YQ.4:/_86)0^Q-E+YMJ
X2Z&;aXaa,8?QG.KCU30)^:\XS>#YBXf3,W(]=[:GIPcPE9c(V0KM/0I6&XRO42B
TH/ZdY#ADN/E^9R+Z5\P\KHS7?I0&#5c5EMZDYEfY]42WW3aW04;E:L>Ie-&C?4:
Mb39XTa5gC:;^7F9ZQXQLP\;]D7Q)e7gR?+aL&0/D4^J&Z>[_e?,Cd7e4,0b[L(J
V51C^>f?\63R70T&>d9(EfK+B0PXPP9NR7>WL_O#VD8><-(X^0=2[/^PG\Z.Q\8B
EY+\=+=eb2HKg?-8HNK/0RXP8>2]BZ8@9L3cd9&+1]6>L8VCHS_[QQ=H1&.VUB[b
Vf[?Kdd#c/5]I2?J6#2KN\<=[:(,C)G&B:0+,bSVd(gJ;JJbU^S<QK<K3D<GeYWO
F/-/cLY^F7U5H:#XNA=-Db7;NU@A-ZKG-RM^]Nb)SAbHGcURH)eb8#GR0?;.:2\-
\DcMVK&c6I;ULOE:I&[UV39Ug9C+()MJ,cIEE.556?g)64Q?c7[bQbN0d:d(LE/e
6N^BgfcSQaHIDa9HQ_K=P7;\b0DZB3[@FCIg0H2fRHE>P#224?041)DKYXIZS(>L
fTRd;0/&>#O;PgY:V=QSKBFQ@C[bcEN\QG,V^#Z520I(NW3&T@0CZ(#TNPc0fg-U
IM()<SYFH61IaCU-]J9=TaLNZ:BeR?ZEdD1.G5>]K/[[[a3MLcQe#0-aK,^@cSeb
.:X;1[f_N7TWE8J@Q35eFN+NIJd:>]D^.@FKgU(XJ\a#IRO#/@:?3J4<^+80<WcJ
ITP^)ZOd[)YCG19EgOHSAG2#76KRfd/;:RZ3A;IVgcE?91O2]W/QWb.Zg>?<]T7,
38E&W^_c1Y>U)#.F>0ZX6S6?,6dOFQ>P,fKDd]5_2HWPKNGM1)=FCeV\E,_e\QT#
MD:NHg^:c/04>A=<B-T?BeX48FODgDU.KQf>>CV@9\6&,Y].ZZ1OdY9XIe@_cUER
.\+R9NEX\<aX]-[#a_dKXT-c7EPBE^LRVD<)BeJ/DW.N3+W/[N+9S>@X1ZH#AK(M
^)gT-ScOP7cHW6<>=TB8Dg?,DVDA/TH>=BQS4(@()g1C@R2+^2.1AMR#aRa3+JD>
X9Cg)JE0B42c&Ge&:HgE51>=.D&TS5TG&,5g8PJ1LgBQ+=;L5BLK8P2aQ4A.@(f[
39Q^Q6QN&Z1F(W-LE.A..e^7B?#\A3<Q)4S,>\4c-4(cAY;.^&F0+Q\ZSJ\BJQDd
OeXQeH&]RJ[e7Vf]3SU]1R7F4+8(/V&(-<=7>&S:eNVG._/Bd19;PH&1-:PAN=cb
e)+;6M)?OO)f_:.4EMK+Y]fU(Ye@B\fVHV\]3Wf;>LZ6HaEd(fOX402DD:Q@(K?,
_@^JE8[F=ZJaJCf(P^B>E^85-PHXD78WFH>KYg8@D,(e2:Ne^U:C;cDFD:@dBJJa
BeU]N)^.3db[_J+/=Y7&L+#5LS)D[?]eZ6\Q]7E<b1-+YANAT8T5T_OX.Q/.;HFR
4QV\cTI39L#?0GdSFL2U&ND-H/QU/,#c0<AE]cQ12,&W\R(7_fH&,O7IIP/QHQM=
/;5HAQ2W[Q>B>]14N+<3]P.M)UBbLY0EIWcEB@P5/g9\@.G:BPc[[EBPQg-#eJZF
bJD,gUP]\e(:T4DTJ:VUQ];;.LP0RPV]LUQ1,69SMAeL7A\:F[e[6FX5E):?2]Lc
MJ:+<7^894Ba)Q+Vbef0?>+?4YO\0P+3\-=&-.,+:G5@8;Qa\VNDeRHXCWOa/>GK
X>^M;&=MaHPOI;I()[,9#DPCT#M1VgG=?P>BG5=b+&g84ddagNBCT=e/&DZ&I2RL
\AcVR>K#fRD\fY\<,]P<_.U?6(N=1+7]RcT(9e_I<8+(Q+T<Sa\g01f/&M[&Md.N
XIO5JUP.Q>c(cA>^/BcLeK:\TeG]dRYDZ9_#)#@+-8(X?&PP5E2IcU_:]H&/bZT+
ecGW+Q+^+\84>dW6g9Ld@,;QGR]g,>3/(Eca^7bZ^&O<CX<40=X)HI/@M_9^YI8g
faR]LJVD+:^@90(/YG(,2ScQ&I7_^VW0+NYcbGHA<25.;>PAEV7_YV;g<#N>OGE)
#gT#,fCe64KE79+U^QOP0c((=,UdQ=0L@_dB@7K-(<XYGebVB&])7Md3.KJ;8_&9
5J-Wb&>26NLdP5,@W4>f@N0D0eB.WAJdULN-N2e>O&YXMAPPD9X82Dg)/N)+HfL9
@OXCC.N\NE3BLI8\)d&^>+3(aG^OUaX@FIYIe:g#cN&D,3AIb1EWZH:D@W9RMX-#
7e/PbfY00;,d:\+1G[E;g&f1#AAGaS,AcU9/#:JIeKU:FXT6b>V.2.]45M/_@dG\
g;XM_X=042\;JJVG2<5?Rg,TF>HLED]BDY0OcW/E7AK+b9<WV3N;^]dQG@d[EV6S
aVUc(g>Fe#[1]F2]_3V=)4H8=RJ66:6.L(NZa6bL+>,-g5I46aY;1E2JE)YX-5+>
7IPKJ0S7S+Sbg/F]^4f0KU1X.DVI\3V[d#:/2BB]<C+0dcE\_PUb\J8CN?_FKTJY
1TgWJC^>1fF2/Q54cBU_=8S2Zfc4\[.\8#Y[U6\_S\aGYEI8N4VUa5/,[@bYF66+
7=_=e_6gY;f77?<a:.Wa7_:K_^0.B^FVVUbaV274UfRd<5,?Q0f:fd.#:B=G4T)<
U,CQ)U=87K5#D_8TE?C^Igc575b19O]O_EF=0/De:<XIZ6+5Vfb#c2b<B[b#I29B
eD7c?XF=g#=g5(9&BA/e[?U]/9_\)-=U<A=.eXJ6cO@5NK-?<RNTBXT5X+]0FYE/
=:Vacd?\O)I_&I6D=:<A:1//A2X[b=,?6_WFfdSW8]]NCfb7\Bd78f,^SV<M3+()
];,O0egbCLM4e0S]8M-HQ6cbK=]CJ\[T(F87PMX=+gc<=9/8[/7O,@TH+-_(D^1-
H8Nee[@YOHSJSDQ+a(aMYfQD6C064dSg+Y_d(^\Z;f.Z70YRF(QV-&fJV360+G4#
0_;JK9>S-H;_K6#2VXBA-4<c5B[C##HG99?UPbIB@;fH[ZJ(F<-\V9DL]/bb_Dc+
,W1FD-gONJa#]^TJG,3;P>I=fX<7;ZT]e.Xa3]?0D4/76Y9LZ;K9@J&BOR7O22OW
cVEg/RFFbR\Mc021^10J/eUBc@)9FH3([I1@gaP\PL6Y4#FD3N&1))]e0<a2ON;0
]?8#e52.&f<ZZTf7eQ6L/05LYN&S)=4O&R,Y[CDYb)R:]/gD?0<Ya_]JD+gB6&Q(
XX^AWdd[WaJ+XK@?:H\KW8U?W2=H/-(RZG]AL4@_eAI,N3,ROZg9>/W8AeA,U=3c
.M4XR_7+Uc6@.4(RR9[9Eb&U7VLZIg+cNNHIL1)PP=R[CD;N#]R5MG6N/DHHag2-
2>IC<92a\/G>ZS]:K9QZ-4fWaY>CAgUK[Y:MAAb\X/eN1/(aBD4d@.XDVA8?-3OF
.e+@.M-GeO4QKPQ^DWHTReK-(1_/D?dU\>_JX?HS@L_1d[1;:KEI7BH^Z]76TT04
aVVWN=I,7(E//e?AaMTV5E5(NbIAZ<7</::Vf9(cLdW=QIYf?adUcA^6b9F[U;V<
f^IGL_83LJZ^XFI6JH>=#_E:N?@Y4S:^egbeZN9=_,gPgfdc.O0<X3N>SI3M[7^R
Q_0YT-Y=ZKNWIY+B^CcPbAL@C4IR</6P<8Z@T5S,36@4&_I?]PPRY]#_GHEZ\:PV
f+HR@?@>N#>R#8JQS89S9(@J(?&b]9fRNK;&Z,0<_E6fd6)TJ/6Jd.938POa)a-d
B-S)ZTM\?3J:Q@I/,dA\,Qb+WN/b41cVN_13b\Qd34UcX<_.S2\Ta=:7C-4&/NgZ
#+PGU9&5KgdfWWT>7Q?679M9.\T\3LNG\:bEPR@\VX0Q)+Q:e4<?OWQY+Z7?QcJ[
_9,6V&(K\PUWDXYagg+H\1]2&8@,_#67^())41FfI3TSQ]eHXOTKME\A)NWE&1<T
-NW[7+L_KfbN(G8/S2E>5c^S]e=4\]c/D+G@G?IQ-MC9:aLfYM-Z:B=9=FF3#I<J
=+a,8X(.LU[dQ]T45S(L,U-HJ[<PV8M3=PUX+JK?^C<9fFc)La5,^&D.Cf,CebcU
2-31[J_7A67SX2+^K;7#RP\2IMR;IS<DJ]75.P7V/WW.ES1IO1B=Z+GZ4c8#LPIY
>=8AY>G^W6YZ]?JA-PE&aec<&Q.@A>;\f#2[M^gbFc3Z-YEKK)9aeN/R[fTce.Y1
bgNQVR.1ReI&C>;UMJVU/c37:@1/Y)HI[4Y-&,c<?E;NFN:#.Y#6T?FXGQ8@dMQ;
??HF3X[,@2G;-eYJ;a75cKY2Q6gV=+(PD+W9J]V@#E54/.=W3A3>+e5K)VVJ,0@A
WFe,)3&(TKEGC36PE3]RZGEBNC\;:RJG\-IF0\(J,9[I5Eb=EHB]1\X\W[JT_c_f
.[S/\gf:\F-.(__.+2=PBEN?CMYGOFgUK]X=KPVNAR>?+J6fL\HRQc:>GX<bKZ)_
Q=/T>]<3[K-4aOG^\b,OcN<;&33D+(Df\Ve\Nb>6ZQcLe\fJA5-9V/AOZD3&^+=L
^[5?GYBS^L,@2H<;Y0.N>5VVXX8NBcSKIA@6>DTO)c6;Pe=Y=9gP.G;0a0Q+AFL<
:K1bZ+N-JPFQHd)_DVP3be^WN=BF\8G#D-T0Vg4&)-cVL#&YS86&HGV6,TZZ&T>P
AWd]=^>ME7K8M;06HLb&0.BWK)X(O2Z5E<X8>d7:]Wa@\K;ccgI1XY^K=4BVbU)8
)IIBa#[8LU^0DX6eWOZ?#N(T_]4>\6P)Q]Ng^=ALVB?FGHOCI:CI-)Y0O)B[O(;-
0LI3?E&2(4C)(/>Z^MY(cfBN.2\5:G?K(-P&C;&SZ8>1;K>fE/VM]P@5N;TVc6Qd
@^>FM0IH\C&\XFZedIH8R_c-,6[LN&<Y;<.^X/ZO8_R>Nc@^_NX<0\]Z)4[O?]c&
,E(D8)-Q3GW2-I7S#+,L;37D&>.7+S=)eIVXZ_#DWBdD=L:ZK00C28WVa+32[@/G
HYO8^4B(B_aR(b^E],(fG_W-Cg2K61=5&ATGP+bgJa@YcK6Xb94VW33[5ZROc@Sd
99CB]/9M,gCC,R^d9cT72INdBY_NUA;Y^5I.U:eI1ZHb<.;c2+7-)Z1C.(.PGfI5
/3gUf-5d#ad7X<G?]808Cc^2,Cg83YW74Pb0OC,356[MU1eZ-=:,XY9O__RU_MOE
e]CQg9IGJ_fB?DP>LN3PAAege^e.LPQ[P&&9ME6OI@RB)a\d)[6VLKb65]N@#@,[
?X?_^N_Fd@>L4aS+9e0]I/C5MFQRPXFd<C<O&-H/1-(X^/=5B4Z[M)F(/a5]5c/:
=.I)L12[@67TG)._-TdIC3<.fE2+1+HVe@B?S]BEJT1\Bg-gaS;]FKK>/3KM+0Hb
3,^KR5F4e\VA;8P_^?1&YXDIF65Y\ZZ]]Q]VUNL4R7.Zc4FK.UJ&G@-9KgFQLT;.
f(/E:+1+B<bUF[@9?fSRLW]Z+f1;;a->-:C4F./2X(2/a[,e4HB;J7:g8K\CBE5<
0(E^]#P&aMQPI[#6B/8O8Q#8_bX<L+_9g8&_Ug>URda:f0R(e<X9VEFEQ=OH-):K
X0_OgL16M8;)>WEeJ=-E5Me7ZQY(2_EI_GDGRFSQ+_Dd.e=[@IW=A29FGSDACFRM
3]g_RN/>2AcdbId+0]:R2(M3IPN[f;@B7&.gDOWU0DBOZZ<ME^A&U]dG&BRQB[6S
8HW8J0(A\5EaR&:GXW2bC2LJbdMUFeQF-]BUdNU8A;MC[\Gf][7B:BgJ5R.9AM?0
b^#O^.X26eM-RN_\LH^.E_&=dDZ\.6.bgHg.DB/ZR[)EdA=A^PC=PY9O&V\3T9LK
aTAU?PT^5P73fYF6=P+Ee[Z3BYd92H09e=;S95,Z3WZU0ASb#SL)/?)gZH3RTKd0
.4ICcf6IfH611QZb;KcPMY\(Cb;&I5[/gaS\J(0\d.0G3V54AfQfV3b;Y27f(F5V
=dDg_A,<P]).NaO<R3eK>^^9GGMQ4L.QA2UKe;fQDHYQa7U\2V0+&E9LAD;A8V+9
TG7K>X1LFD1/QZ31W9;8<BXB)CE(@49L#O2[\^@XT#+:R4)8C@+c7]+^_>cAHBAS
6ID][@[(L3<>HXX\-_[fH0HS14QM92.55VMB7^H:VP8WPQ=a9#G/L8+:O)2_RZ;,
\+d4EK2L>Z():<+TJLI88MCZA9+WK#O-3H0HKV<,B[d\3C5[HM<bcRST6K9-V[M5
E\=T_4C.fYCeS&L,=0SLe,I1YC/XHGV_E()XYE_&>c@c\GdPRCeN]>6IA84f/db5
<#]G[;/#QGL0+2>]]I],S2/e[gFc?BCQ?7SOP.AUgXDe>T89(+QRO8S,g8T1OHU)
@T?T0^JF,a6CXc+?(GG59#1I\(;UCSg:OS(c_0<b:+R:]QVA/K)a3#I?@9WDZaBS
,eG?)D/]-bBIVM4NV;bC#-eRYU.G0;;,bPNS/>1a-RDd)MC]5;-NJO2\)JAg2dWR
VNOEaE<M8AFQERI5cBd]>I^7<O1#0V/2-&#H:]\dJRbC#6feNN#,QTUR@JD/-[@L
4X+)1fJ.M?&U_V5M=aJM2c06_SW5,=4d_7(Q8+S0^([+;Tc).M-4VDO>9A<M_a5]
dZZAR=a#eBfIZf7,A1@E7TT.D#ggZSFbCA#1e>OgB@cQJ(IYB/_Jd(PJY@^_GV9e
gSC_#bL4G<cT\BP]S;W7CVQ0=;\J;fDM=Q:&a9H2g+//<W(PA/^Qf3I_gK76e=V/
TR3-,(]WGK(.IJ32fRUEC-D[RHB;Qd0?E[XQ^IPQc&Ng35A#cc.C.5FD8;3Q(1CT
^YB3F\Z5/a:-a/YaYdEZ/,Ib4VH>/B_/?0(^LG=0cE,86?Y5_\\@aUVcF@FFEE1A
NJL7SF(9LN\B3R[3>8PcP3-:CFg2,N,_6ZGBdI-@gPJ:Y-&?VI5IXZ.b3F4Pe;OZ
X7:PTBaJ,QFW9E3@;Y7-:.EV_QdJDA9,3\^@M96De4]&Dd)WDPT@7MEAH.34781T
=YA[JfHW3/B1N<f&8f6XILS)_7)P)?Q4:)>_9)&eCd7H:,=(/):)UPc_\V096&Q8
N3HAC3)_Pf1DV<S1-2N4(cD7M#H]bC<7gGX9)Sa^_D-g.:X^Q0CN=R1.INN>W7,H
P[4MX3_;c:>OM_EGf1K=);3eN]W3#]@;KGd\6;fR0eYO5?c>LNUK&=8c0;g:AY3O
W;G9O+KVNd-OLJ&aZU27R>;^P_cKg@XNX<aT6daU273>dXEIbW+>XCN3>SCTKa=\
(bEQ=E#T:JMTZ]TOH=0F.c5=@Q)8[LU]\eAIZUMKM)=ABS73B-(_DR(JB1f/NMYW
X#(baW7V-XE<:NL1VOKK=b(K^eDF7I7W(:]B@88BaC&DNS3LG,JZ>1JJHI\aBbFa
.&\JZ<\L\IaT3&_;YOb9LGFOK(:BXT?E1LD:H7.@V+S)S)PX8W.bKdX,5:fg7AV5
>G+MC4U8EU.DE+J63^YR^J[80K=KOMNM@TOICF(Z:Sa7^)QW??=f6ZR7FMT@-&5B
Z/&<7YfLg<,d]S2:_W\93NXe4G?7PXeb?\7@?d(B-;M4gbaLZCETJSOf?]@^fE)d
3HVC0.@VfXbO-)E(5TL5N5BFTQaZ@CC>DK,Y[65>HM5NFYAX=]ZQEI^U,H/^V#4M
<b:dJYbDYRd2K.;;8EK_1&126cM9fIKUY]6fR#67;fQL1.cT8J=[VbKZV[FS+;__
\_gBFP<WZWQ.Y64]9W@#c3)f<YU[?:bN)dOgCM4_?8]S8(^U42=@_[;,GDP[cRI^
P:SYV3e5?X&SB4X_XVG-AM?(2(V,;gK?^UY:E4FS.7_SaY>>QW_1FX[U:48,@O_c
:g.A^;cZ/8@X1FA:M?U?W5LU]14B-M\8HG5B0+K1:+d89H,\E>#=YB879c6\RO.A
[0O>WEL8bPf@d;@]4^(9V>Q3cD>^\T[_3,IZAT))EG@,W_Me5)8<_:=>KBQZW]&Y
MONYf?R9de8E/CUM#1@#YB/B,V/L+LN)5^VR=7+P:3FH:3d\LT6BTcD\N1@&U3]I
S<8]g^/O/;cdE;BQX/Z=)b3F2;[Nfb98F@a<N0Xe0fY2C-,[W\U?C.9N#30/NS#g
T,R>G0gO82HU+8aWLg7#R]\O39LcIIU);)]5+W>#6DPQD\GIJ>\)WH--WbcQQT.+
aHMFT6CI,O2b?NfT]=1S,fUZ74JJMUI_6Aa=YMHAMG^^Be+<NW8]X:YQ3OI)#?YR
P39,J[acee]?TQMg/\#2,M5G7a0OgB&2dLV3JZZUD&cH7Mg:Q1>)UMJPZP]AD?-E
fHY-+[Q9(E+EAND<VeECV[EYcK64gWI(M4@[_-Y_#Ad-J;GH@+[QRaAD;F_WCT<O
=J;:IJe<#&Q(PeW@L&E6&X7RNTGEJU8UBa@]6?X=f(:)UKL_Q#K6Hc.05P[>#W?Q
.ICeNV=,7):W+7\Fd;Y&:[>QfIRQ&#a>MI(fW]@A@GP]QOgE2F2V,\2UVYW+7af)
]O;R^-GO2,+:f;RVb2.,]=ID6.(W1G2OZ;&,d=dN.WEWeFWg=@2=7?(E,([D97eC
Q.AV?Ab9X>U\d-V-:=X+4V5g=?V>N,&+RId;GG-4JY-E-)-]W_QN?,EW8JV2e,eF
?)?KVO?ZU+(?&<ARHDNQ?\>Bd16Df)B-^LRbD=3E9HLcG88c,?[fdR<E@OB4F21d
+7+V.<;:e0CF@9[)4S]5,.9+Sgc2FdB<5bdbf1gS8</GN/.>edbf8+(7X-VEB+2b
_aQ,DZ1:HIX=_SX/d#eOY5L4><A<X^P1LJ&ae9:QScCaa^_MU;I4:UeI-9IfK5U+
Qb#Q2DE3cY,LM9),F#<<[b[WM]W?:^O-H@UZD\;U_L22b;d,<E_5:>H1[<]9K@]?
Jc7GO/Jd)dO9,D&FcK5Vf#a9be.D),W/;#3BLHZ3:]X<T2VZA^<cL;E(f^,PIZZF
S:[]1/f/gL,I)E+e4LUHNU53g]W>TIO2aB&ERX_(-adeTGcU;<+5CVVR(gH-?Y4e
UPec^QT>&8J:PX[QPYI)KKT,RPWG+@DdSGd)A\O[W:6-O3[LEK7bX>IdX3(^]1+H
+\YG@]PAR36a]_I[7NYXaLK#@/e?5Z&2DBH.]e1.bcFP.^Qd#bG=\aP<(b9\fC<]
WFQG]L=&O)Q>d3M>1D@gPO(f;<@8KC>O:ZJX/E4:QVK>(D76Y\MQ7:W#R_RP53QB
IUHd[9WCeP2V;US#Q2.f5g5\DMOL]M0_7_@-X33;(-._DQbM2XIS94Z4,KU3^:Pb
Wd@?J4U3-AD[H79Z.SSb3AKI]BLZTA6A\ZeMMD#cD</ENZ>G24Cb2@E)+S^fS1&U
BH^P)_T(I&QZ,XRNG5AdaF]E0N,[ZgWa:IAA3:>:=02DY/@AN\JZ/03G]).ND^EM
B)+BTX4I4=McJ^2R1Yc^@XD5<EWV4F^QA[-#LIJ-CYHZ3:/c,W..@13cM[W=f4Z5
TUSgHUOF>bJ#_,]8Fg_.N^42XFI(>^771L)W@]d3c8:DW7g[HEZ:cQO7d:4[J)(T
K#N/(_Q/eAMS?3<.2[/>T>7HTGID6Z,?=#S]1?&,E;FW#5ga9c#HQX8()2?:;0=J
RB,-<Q+#^0[R@H:-@E[4ZPC>AN7J_?\98WfCR6ISE8DL^1LMNYU:Q_H\_7=AN98/
=,P9eP2E.1_3+,\KF^#SIK#,3#IL-#]?B2Y0/YA>#fZa+[c@D,TL&,>S)KCIU_G@
HMgbW-FJOP1HeU@1119MW.__1aDC60bA[0^\+8UF:-NG=D&.cR#\#?PW.a)Xb+.c
WPC5(Y5>a7CbU,HXI\3dKDS8>-89GG(,3#2C3<7RBV^V1>(<_:CHWX[W;O\4#(S?
>-^\34Fd0JGd=G]4>=[AWeUage-L^3Gf?)/SH_Y>/+NEGS]:JPN6W?8V^fMP]RW_
dd(XFU&@IM1T9+_FcfHA7#UO&T?=C_fQ6ZL.I#R&LM3Rd)DGAC?^3f6]Z>QNE((N
aTBaKCP)?\2D37/)a_E]UWK1\C0Z0,D\/OEUFO>cfWfQ7cK]I-:/V<W,8PZM^;.)
ZT.))<INR=Y:.4dMH_f#b)73W2_^ZG4>VbbPCb+E<gQ>@U9#9\]3_3P\DeAWO<F)
/T;2C;0[K.@.7FN^.bWRaD2V-gMK90adBD)I;[P.c=<PZFE;PJY^6?K.d,YaZ;L@
]POT7FW-0#A7_5Z<cMREQ@[,X2Y3QTB?Ocd@UWGXRDDc)2/QKd9MIH[[,QXMHG5Y
Y8GbQMQ;?LZ;cO]-OBOd[IQ8BI/X07@cNJTD&CScQ:ZF@=YI;,/+3X-fg)Xd]O5c
D+Ug?>Pd[?-QPCY<GCU(R>\5DPcO=bE;0JTZ<41\MW1=(K9AEOTUPCR53g3P_b<G
OFC:(P&5=@?Nea2;R^\Xe+?MVN@.1D:BI;L@9\@P9M=?SgJ&[N-1.D70,THegf.#
\FEb;^P.PUD.]f8c4V.&@c]86TY\;6M5&:/ZO^49FR[UaeA)-e6)V4L_KP^S7?[1
>;4Q@c3KSD]CWKCOA2CD1O<If(/42=Wd&HJb7O(O1cTQ(fQR/AF=/eIC.@^Z/S)R
7J?I.8JDD1WTc=@7,&Y[VSS\N]\RH4.1EAU0UB+BF][S@L<.4SIf@?7<?LI7,9X;
/;L&IR<5P^7e7S@d1:1]gbNU#PNFE_EfJW5)?9A8&)F&1c6HVWNNS@8@QT?M5^&,
X@X96,c#=75V18GaC4&R[,9EEc4\U4KYP<JEB-EMc>GHAM_L@MX/,,eNPR=P?+Y.
WC7T:f0d?3f\)B6gY<KE)OH19-2I)G9Q?3Z:EU+bM?RW5(&)cfd2,D/3W.(f@[8/
.FW#8<BB1?&LcF,MM(4R8F1UG&M+GN2gL.^MT>6/H9E4>X]P;-R?B317QVFYR85^
&AIX5K9FWI1\+6N.F;PQ;YUMSJ[(AT#;9[7g5.Q_I&EB)/V5T>\Q\4,7;#,I_0O&
#I\^T)O<0_F4^T5Fc&0X(08?g^L)BJ;NR:P6K6d^34OK53QS\592B6^5T\Y7Y2K=
(52EU)I72V2TC+6=gR9[I6C_0cNH<66Y3aaZL>)W-5f#C]U\1Rd-HR0>.4M@F:Ug
+T>3=NDYSU.=G#I=AA_#:12Bd.Wb+)H=?VCcU2386eC<Zb#5I2a[9R=Y\_=8[]K(
JUU+<V3PJ[FYTDd0[-S3GGU:),f7N:2_,(P&FH157P+P5MX+0<TM5)QVPG11.6UH
P48O.1,dE&7DCP=.?;BP7,;M,J<7WNbSX3?bX\ZA+S<,e^ee9ObA@6(bN<)-LD^2
6L2-R)8:dK>d)DaULP,a(a,M>JLb]CT;,@DCc@)eQE14HV(Y\:5Q[_E27aD(_Agc
KXO[;&(R8R3CTUT.ET1C^NGG,c4N;R(Rc=(b(BFb?32?Kac+HWVR)8;F_UQ7TYJ4
ULe:MY^>dXH@IRR:GGC&-Cda[CG;F=>_aN4\A#QAdRFB&bMVFA.eB>/?Tf//dQ8^
EDNH<f&IW]S>]H@/FLG>MG509-;LU#9W(4d.IQU>(/7?;gUC01[\QP3FgCK.VeB:
EJJeRL(G=ITYQ:B]=Q>ZG/\<&X(W5^<44:E;/Xc6EDdf5;0+TDCJ22FbN5S]\M90
Gc33gOZIURae1QP#O@O?NbH24&Y>-T]H8([_+WMM@,gC?aUd))4dTDgacBObF<&X
.bQ&RW<I?44_d&ee0]=\+Ia8G1fP#OTCFM&]<51D)VWM9+/C74WWbE,D(I&-P+S]
9@MLG#IN4K@35fHCgCUAOTJ?YC[S>2fQN0NL=,W,@@,g])ANg6-_F^J)UHAX+[U.
[Ba-Q<PPe)/5=O2(fV=5gUZ>Fg>6NN4B<e29HS+C&GV+(YGKF+\)=UD)6b(LO7_;
<<Q=,UJ-C=Rg/M;<L#(]Hf;X_-IeQ4e^]&8]_?PNQ@aeN2#4WP]H,3@73A00&BR:
f3cEe?\#MWH1dg:c#0L3b<>6-GY=^DFQMT^(V)bW)6+cD>J=ZG+3^R(^ad+\?9^?
Je]e4N85UT)ZgBWI1.0f@AI)A6;4L#4_@UIdYD7:/QPg<a\gVXOI/A5VVbQ8YHJ5
#9]gZJZ>=AZaZ&\]OSccRA&eb+1dP<8F7d&cE[=Y-=:&J-VRHEUFFF:eeTYZ#\&;
DEgPWL^@SGg87dNG^9+UPO_Q)A#)SNN\KCa;5K\;Bg-D20QB3VJ^\3dW4F6[KQP_
J6D,fAGY0OBV)+3P2dL#CeW>2V__<6([\Kf]3.][;,#JfPIcTP80&ac.aDZfT-0E
cM__?US\fKE2R4PQZ=#BTS+6VD/-^c+WI2VE_HXVFO><3=0MWXW:C_MBC:d,AQ5@
MKD\aUV+:^Q[D+cVTOOM5<14GcR6aC,]&9dB4XBaUY5X]E[F._DPe\IV6\(/3PTM
dPK#TY3GW^F]GY;7;I:1B52<e>O]b((RACR6)@]RZ//@eQeSJf(]J/<WNSD=\>WS
QTJfJLEN=7dLYGX;M.]Hc/RBL^[6F2Md(A?VAP_XULRFSKYXWQHe-1J&;c83U-W[
.BdB.gF..PIGXJTB_c\aNQ_/0&-b]NE#VX&&+dTX9)^GS:dZ=[B.&(6<5C&2eGCD
#^CYQ;[cXHZQ3U(IY#U_]Xc]8)OHXNZ1@7_ZRG[&,b5M>cE2eP5N@X:,K6VF-gK5
TWW#GR<JWg5_0)(P1:;J+cBf]VG4CDS0QLZd@F/B:,#_;0^L5d&LN](UGB2])C5C
e@MKZSL41#;C<D8N37:D\>PF/Fb-)V=-C>g&&Ede598)]a@_ea,X]K^4@-]BeQ4#
7A.X&G4.C47aQ;Y?8PD3dWTI)QOS6QC>9Z=;aW+:e@W;C@QXa5#&\R5U_4](RZGT
M41_KPY1-Xg_0+g0<)[dVKY5G.bbU8>1D(O\_0A3N#)GEEZ]fT[5QP1<93MX950+
KKTH?#0WU/AASX/#K+?3^-N5=C3_H9:+Y@NR)M=J]BgcFMHNbc/LJP=]MK45D/b>
R,AP?F^XO+?c(U@1FIB@&G/^17/U3f)#L:[WSY(&6)e380UbT80XT(B\/HJ+^LWQ
YN#>)AO)6XF)Ybe^-X=4J/>PP1#-E17O64aT=d[UE4MSO[;AbO3NQAZ&:P2#D-6Z
Yd,<.],GVg3bEZJB[R&JJ^NJ@P9H]=.V2c8WZ)(^-B5,.]7APT9SV]#=ge4Z[679
&B_ZG73;fb<Xd/546F.(Rc@NNE5IcO>KHFPgJRbV.I9Ve-0fbT=<AH&OCMH)7c&@
,C,;VAd<fg_HNSX5I8C\-(L;V3I9W)R.KUKX4<gMSYJTFS[\7aA[V+.9d=]9I22P
TMALTW<Z9675YUZO]ZEM>910Jb:-HWJT76V0fTccT0gD(7+L@4+-gBV7H@gE4J2[
Qg]/8e-(WLLd=PW99J60abWCK2,Xg,CeVc#,7H?\QS/72O+OUVaRI2.gDH^eVfa1
C;-1&eB^R/1]@?LDe/17R&SFAX0=@9VE8K2&ANW3fZDH9Bf.:WYed@c#A1TGH?.d
MUc9?WEbeO_BZ?fQRd3\-O?RCV]>U-ZVFS0/YV^KKeMeZ^#b/VI/:7eABB?QWA:7
CG8]IKYX_U\HCWM#5Q(H8UV^1PIf\_9F5H:dDc&UQ9AK@e/N@W/TDd@ONd23__Jd
ZD/WQATD9-DI]c#\ZgZ[:+5=+N9BCVf<3,:JA7#cL9LaU[SJK5(_:/)LNIS7Nb8[
[)AZ66QPXdW0f;?W\KA4FS^A58B>(JT.=]#KeW9[ES.YJ8G:=(K8:.MWN9eVBfc\
WLdWgSGXYDN@EZ)VQ+4<aMTY0:..1VQN#D-NS&I@7=?,Q5MFY-@R>&b^7a#4#JEA
UR85K]I?4X(I[,6WPNAKUfF;^Tg_M@Fa(#\YUeZR?&f88f>#7UXOVI@8<;d=fJ&K
N+.=fRF#E)MJ08H3aa.1K)b-@TcQG/^P,T2:_X3H6_56QH[CFg]a,U]\6(\I0,Na
9,AF4+DO:JWY0778IK=FMT7H@V^9C,)7e71/a+M.I#XD(RceX;[Qd49Q5SNLG/-g
0dUfOVVL&\/=:);2<DMOKJa9M0Z)A9aKCC5&a>>2NH[:NY9fd1FPKC6))QEW0)VA
O=gI><D(S@J??G7eg#Y[1:YDZYU0_aWUN<ORX_6Xab]a@TPT/[@A;O/gI[A(D?&N
L<K\-S5RK6(f,RC0fI/2A_]+1e=P\gK@3ZE]GHU7,/RH)41f#O1X6SP8HN>RY,5@
\W.2GV0;?A\XGA<C6bSd&@LC\^<+:WO\R[_fJU.&HU+E_>W91g1UT0JgV-c1+-F<
B@P\KC:D<AH&W:gc#Fg4b95NKG]@C^a3f/]?V.3W](g-N.^,HgBHfWU&5+cf=(OC
a;d/F0-12J#5fZ2>T94/7[=ZJWMA,,3/8:Va>P+K<2cG-I\M;\CO#c)?2\N@2@=A
OL]>:]Q+UQ^?W>CL47@Egd5ee@A,0X&F3S6)S?HQO]F?W_(aB7bQ/</.?Z#@,?EV
g_HgQZ^NMY/-^DEc^IO4>5##QAWI)?L^:EYW?GHENffZedE]:&L^\NGT72P8>\(A
F[XXc,D>&]_M^\L&[QHg#H]W3LD>UTM6+SZ2]^T_(9EGH^e6>CPa93DIO6U5^.aM
DdDP0LcF:8RA:WKegFAE1,T_6:g[.:6b4DgT]]>/T#?Q4R<+1MD,A6@a.AND:Sf_
WE_DL7H<A/6\V>_Q_:[;;@OAFK&cR.Z;6JcG#MaIf-\&c]Y=<&MI3FV0+F&R:=0M
1WO,+[PF.MSQYgS..a?5Cg&7Pe<6-]A,;U9#WLY_U<4Y81]XY#97J2gG)J1>2/X(
YB5+#92S)CD)JgHE>F;fH&KB&>OJCTLJW>^g<+;/;D6Q64FX8<Z-SCaOdYbfI8W2
]-33BX1f)/4IYa<,XAJAXJ7]#8/6+3K1YO&-VEHf^DL2?\4M1K;:XU#dK+P:A,GJ
B3Dg##7+IdQ4]/2g--FMXWGd7=NV]OD#OLIHVQKV0L)&gb>HI2#6#T1?4XOFPe2T
Y_^0g)0^95+7EV;,/ZTb&1C)&U.f?11]AT87-ccV@c_YS48d003D27R3@>1M-XD7
1;,(9D;)L\XR(B52g.-gT(M<;#.&JJ?.bfJ4:2=V+1fJD;AB;DC?f#-IT;d@6C+3
F3#9eEQ60N_)dJXB\Q.;T4GgGI;MaT1:5;DW?V]X5.9,NA2FYGGS5_ABAe4I.6g8
BP0f^/Sg:[3eU4E\a6FJX[5/dc(W[a<),_gc-#V)2I87+MOTS(-EA#V#f=ZL^:VQ
]S#/e2PAU\J+AK52=ZN[S&)F>WaJ9cNRbT5,-Q&C>VIbV)0DEd)(J]8ISMUV_P1K
M0:UX(7:+Y3?EPGf=NH5b5M+]13I]XC-]8CA,PPNM6UF;25f3Q\417QQGTFP/\=@
4]ega6KKXD?[b0P+3P(@YXdB9Y]:Af(90>aUS_<M@^(OPR3]<-9J?ZMfQNF;(N(0
03UWX<d1=@e[Z[+Ncf?THbF0g[56g:CI?D+K9.6X<.;.e[bNc;I4+)^<)L[5fUf<
HU8,2HcK8B<Q9US)_;J/_H?>0WAYe?FOY&KS(I6<gB]C&H)d06I-A-L>SA)Ege/X
5a1O6[+WDVcPEX6#A<D)C8cOWf6Y;TAJ9&]0O_W]U&Zff5Y-8,C@3(\(FLZ=0R#]
a<Q]PTc1[7AaB2d3PXT#f6M8-9(eaM4M\6^,2N:FXA1X1&SKOd2Y9\:K+>/72Tb0
7+6]VZ.&-,YUEP&WJf/F/C@?JI_-,gR57YU0R=]gT6cMQZ]L/CP[7RT-J#-ASTNF
M/>BM3a\>)6Y[_B@;[DCe&1K(.bI;P8Da.55HX.=a3Q^f2:a-NbBOS8)6b]ADCGQ
MGP+)Va.NLQ7QUd>-^T(V&>V2e>Q?@(=BT)D^5WCFF;BWBLcc)8HAE7X]<Q\\.;;
)3_fBJT:/2c[&R26QIA.J-_2e)Z#KQHA,>0\,c\ZY9,YG\U;HO-F<]:eV\.@PCF<
,=25J9FO1VP+EV\OP^0M,)SUJJgE7E24:T5(&DV/D0fU_C<T1V#1Bd^(aFcWV(EY
RDC9ZVfGe@R6d]WE4Ba7V>XSG8.c,XZ=>e,<@;ZA8I-+RN&818936]J^8Y?gS:_?
RcXM&62)dS;#0RCN/<WH3H6[??V?2:gB(+1_@P1Yd5:OC/[^>>\B\67U-N4?-f:f
cR#[Zec>TG=c]12NSWJIR:ZPC&Xb1E^DUJ]HYG0d^)@g[M?ZRXKgU8?=D5)655A^
/EHZ-NFQX5]5O\MAf:MHIJJ&dEc<L4VMd-g2CKL@:_1WZTY2gLZ-&(11Y1d>Z4P.
e8.=P6<KYAeF8S6UOD>+V5=@4.TFID4gC-&6Y.Z]N@8KfT3;f,cXKR&eI?FDGd&G
bR-3/T/M[4^6HG4g56[,6W;5R0K><c)QBaRDgW+2bB6.eB/(/YW^Sa5)R:&_#^GX
3\N;1,E,+KJAX1S??O3ONIEfWC8cFM&(P8=U<CP0G.56M/SR2^J]3H3NAE?=MOW/
M;.95+)cfBQ9_a@8EOPLY[7#/;C^DP/@3==O1-,+DO1SW+:(aKM@d7D&D.]+EO]E
S4.GY9M\@8+\EK_I#&2d#L@8E/LYI,HSD,eW/S7^ZZdH27LX.fLKg(>6eO=d)->9
N1:_8f[^O,/],-GJ_IJV:c\9-\+4T,5S_U<Q[g-I5;]7a=-H#&<>a1ZOa<b+[YGO
8//3fNO49A)-KQ?V8@+.S9<JE/:.SV[[9Jb\)HVE@M0I^JM0a7::9(=I>e,CbHP:
\dd\g=C#W[U#B>?U3d2WWH_H&T,5?fXLV75I8&T7UKM;gA;DF2KMLC_SJP8QF_\e
4LBcQe5g9b#XZB\8J^R0(VADERIX]aM-R-fPQ;#0dM_903VWX^:<-Oce-C@AI5KZ
IK0.2<IO@FB<<)=,;ETHO,ZEcgGA2=8,[/RLI0NP7M.<[?/H?U;B9U94B/=TG@+K
I)M2@6\KM]D9+VLGG-E(:fYQP@QN2,S,&]^DY\D9_WF/OCFAdM??S]3VUZ5X&7Be
)L/a.+:#7YAA#[9;bQ9QbAL^/9[=J#SZX,I_XXH0-2/PbKQfee6[QdYS0Nb==Ua:
?@Z1NLA^LJVRgE[;a;9.\=V25WWg5O1B?W()E@<4:,L22FG4\c@0Xd97&e?b.>GV
\4U:MHM=eR2UO+6bKS/;<8:>U.f_@Ng\QCI7D?;._V9)QOc[Yf)E0bJS4&N[1V<\
^JV#Bc&Aed?.7:N414G:1dY&cOdKNV0Mg:K#Qb8W5LL0;1G^:,+OGc,=[f;b#S)E
#:5I2eAObC:Z=,GU=M88&<J4E87g7Vf6SR8?Q5L18P5)L<d1F462XPNV_JdfRKBV
?H@]<;0==M5E;N@JZXaD\Y-Va:\[ebKe]//]:aMOIUFM20.-(B?6B,[1LD^d<S6;
[PZ^ZIIFgfD9G&B.,a2<1MAZCb=fb0&1g&K=70aH4<@G))F__UY,PLERd@OD1c],
e2EQ?IOPSULb1Ug)c5#I&B+a.Ecg5COf=]DDC\WbE]J=LX2Ob3>LL6I734cI)f)-
bY_d6O48e.X-5L2gGY/#NFUeY>^KV=?@bFN25MO)e3(CJCA<4/4Z);.UL>91IUK+
Y:G2GH39A3e@LSaZb:e>@;<#&fWRZ^?;2KW.a8Y+bI2UI#f;T#62,^7+)6dAB2U?
ZX+8C38\@Q4:#.dY+dM1X;4QJE#[(U^0gW8.ZF>D(8aDH,G;ed>#>EO@Z\TUeI#D
04N1]&\FG1.Oc4d_QB:PV>:\&NP+XbB([-H6#]/NGKa/#PHDDd1S?)V-?&L7(:.X
4^N6gd:@W=K8A+Ic=XMK+8+XeOYR-FZ1A6REINfDa)D?aaS/@Z\MV8F5V/,KU&]-
5HECRcY[0c14)g35,aK_HJE6fNSRBb4[\^#HJcYU6UX]XO>FWXea?R+W]]3A1Y@d
Y@XO=X6W&2GbID#7DE;;@/6>XYM9_?BGO?a:(=WbXbIQ6I>CZB\g@][)dL9/S30[
Z<C>L_e\UB=Y?#Gf<R)_6d&T0V1I\Od1K)a;+a#CZG3VH)M<US624G^TVc,5CXb,
:f#.AAG\/<1235DNU5BOTKGRB>]W6=M<5.<JZ5WaBd;<]2.DSfDBY;47cM+S41\^
,MNWB_E5B=64+BB+=D/0K<_.M@:Q-=bfLfG=fQCT6;Nec-VeE0=gf;X6(UOUJTRe
[ID\CGeULHG;FZ4453UYDW\4ZEeB6Tb&XK6J-WHB[4cb+GDfe#\@.\eNQ8C7CGb;
=<56ccM^]eAdK^,Bc6DPTL>+9^9^?G^M/6ZH@5,A@W&&\TMVEJOD+&^S/&>O0\-A
[a^DJU[CH)>#(_JgG^XS^.g3a<;YWfJ6,6BJ7^?VD_C/>_.1>LBcE<:g(Q^Wc-Y7
&Q[R[UZ,_Pc_D@;?6Df]bBT\g)_/W8/W3TS4EU_dHSY(&9L54N2U@4#0HJG2972G
DNSL;>7[L#D4B-_JR.KG)g,)(cN6_<RR.B^@PI@EYDNY=D\gN/(7@0I4>(_<e\4K
PcdQ52P@6/8MBcM+3b;@VA(H4A:3&S4/Nd4?&E)Y=))fHE5KK;0#BM>GBSaU(2^R
QHB1-F@:R,>7G3/ZOV2ESDa6.KGE]1e_+0KMZ\J=NFK5:@1BPV/V(:V:JfZ9Y/#:
g3-3LYB01198&+QHU+:a&DCU48;9PK#JGf>b7TfV/8L+/@0?DeZ1[Z3<CHCGfB8K
:EI&gD;U,fDd9W)W#Q01FO84KV][Z_.Jfd-(<5Bf;ScOXLVW9.[7>Ef(U+EX>T;\
VR(>Xd0EIRM4MST>?bLZROfCL72:\Y?J>;F68:eRf#R]>H&>GZ1]V80_&;>>V&MX
<bDG9#6D4Wba8-c_].\NPbCM/W8?[aAc=?D#A/)PLa2/>ZRfQ4/(aNY@6MF^d:eN
DfMF=;c3Fg-TALBNYbg;B&3J9FA=/,PT#9.dB:>7Q4-AZ4R3f_00@.Z:6A7fZ37e
ECQTY.,:;_ARId<K08DYJWc-I.;:#4&c;:9:)^-^C_Zc4+AA-G_O,Z1RMM+6\\XK
gKG76P?T=NPK?9(Eb\(_Y8eZ@J78d7Uc,\f@/0-.aQeZ..9;Ifa2>M\3#V:O\4BI
BU.2ZGMNL+N0(T]ggggSZG]fYg-=eS\&7AQZ;__;/LbL-UO^S.G3b)35;#ZX;B+=
U;DJO-];GFVSFUNb3-(HB/T0]+A\ER3O#R#UIGJ5]&\]MT>G)NLH732eE6LW>#++
T(ZI<M?E;L6HI.D4@8S6W40Ged)VE5O83K43b-DLYF:EfH8>5YG0C#HGML<<+I79
8>KA+UW5FXADR>P37CWP1GHNaT:@dJbC4MD>7e)AE?#6.+S-<5bP8b/PJ#S[&TP?
3?.fU=GW^KVJB38\B:R,JR<@_E9#eNBY3a;(7/E&b?<W&LUXU);4/2.2d#/GK7g2
W]gaIG/e0K1:b@-Y]I3918Bc@>R](2+GE4,fPO\/T8_P7f+1UQe]-7Qg[L>>GQ3=
a_>eEgZScc+TK+0ecA(,G4?g7F(E-eY9SIDI03T;5(&H7^[3H?.8O>X78S23a?@I
&>T72(/+P)aL/KgOGGNBN:]b]BeU<[?;GY)8(b0S9?L-gRKW)(=NBR&MLG8P696B
cb7gR#G[J)AbLRQL^62)QI_1c5T?R)0e;\>@:=55&E3<P[T/RG:--?7\(HKI0>7Y
Q/V(3?fQ&P?;_GN8H.dR;B_@.;,[Z6)abTe41(0D&VL8T\<LO2A:MCV\]^O8SLbU
TUB=H;5g/O+L/(BP-G__P#Aa=Z5eQe.cf?@&MLIGIVPCb^LZ,K#85fA=([V>AB-(
077R:4W@C/E97NfNDKD0#JO(#HWE-:3:NVU/.\Z^72Q5aUHW_5Z(9Q:Y:(BB.^-0
R=@U(8(/\)LWNaQ7)fLGEU[O^L8,F:JSE20[fJ(1OT3#5eCH6G9g&XZ@+R;I,g0&
2DC7R_=>&]6LXGBCGB[7:_dRPOCaR[V(A[=G-^/a?)_3B5^)NB78OM^2B@FG,6O8
=Pe?G>F9V>EL-$
`endprotected

    `protected
a&S[6\87e/_-A.CQ@BDFQ5e8R&OUY9<c#67^S=JQV-P932gL44Cb5)35+HNP&fZM
+b+6JFdc1C<8YBTA9\9g6MRcIJ.T0VWTB]Q0?INRbV49F$
`endprotected

    //vcs_lic_vip_protect
      `protected
[7^>QFL,cWTV^SO9e<TS5306SVb;>HYGQT9,M<6]TadWTa.I,f9,)(\K[K17B6:?
172f1]F:E-f<Y^]>#9Oe9A)FNaWLg,/S,Vg9]c@ge6-N)IE?3U=4PHI5DH1fC+?Z
IO>#)<6H;=AVUFeW,T.MI;(e.K04c:<(VJ=]C/:1UTCB6##XOaG[;<6gY>#3//WW
X]g,PEQ91]2=8/7IF=N7XB:RdK_-(<.K&7a))9Y5&X.:9Vb4M9BYVI/&ef2Oef_V
=7#W20^73egVGI(E<5eYcR_?7]UPPFM,?PPQ7M5E3U8K2SOff0Ac#R0(;0U#^V--
8Y]QRbPVKVJR(@QL0BVB)2R073Sa0RH9V<_>8>cbU4V(;aB@0?3P]_e].:X[+2&W
05=HL?KgS_a2J(11HY]+Ca(1CPS.1L5VBLX<\9EZH)Mc4+)_JJS+>:[W\ED,HeXR
K>C:R673cd1:gJeaHN#9cI?NQF:[4Pc4(Y/8J@)<(e#9;N#Y>^cW5,>eIEZa#eTC
>33S193b0_+)AQa4;b>NEe#,XE,#+4(UTJYY,D=aZa3Z<L857YK&bCROgV=Y7_;g
g<OQP0#HN)]cT\RH-TcW6)YGQ/G2b0?\_e12,W3(Cf<3Ic@fJCN2\E/cQ.J1<cF;
A+LK2=_E3Dg7;4.2gO^>,\K3-6Z-aCc)c0T15[A(93C:@?a71>=2Q0=;XBFUMaK@
RcJ;5<C@.b)LQX\=91MK^GO3bI8_+@9^PH.6@D7=HX1V_]^:\]gb>0SZ+V]Y29S.
Gg>(>BcC-2SZ,a/CW@cHU@[RBB4.3>3H+;&B()cZ:FOX4?19CL_DF>fB[]GYCK0P
H7;8J^^WNF?b9^^aVJOb;;R.FJ,Y]589eAJd/8e>L<B8(9G>=CU8\-_GcV&:EbZ2
]fDf/3I:NF/H(d9.2N]Veag>c9#I.:\g,L4aC+LO6K^Ie<-</^G6-,)]Vg@@1Ke/
D7bZO],];(/X(c7J@,0-65N4f;?8_+Z55[[8V8XVQ_E1@P#Y9gf#E/0:/PIO7f7[
>1G1Dg&[4J;[AaT7d))bCZOSdf=3a:KcN4+b9#ZKD6XSeW_1MQ0=IXQ@(bBH3eg:
#a[2HZ+a^/X&VaIE([4?f=f+E<Ba-P2Y]0LBT6d2)(OMA@U0/.=60>P#@R6,A2>O
,:6JH9#3Jg:T(Bc\PRMLVc/7fI14GS6N=PK5P]0N9@)=0AP3<OWD?;I5dYMPaH,U
=402.RCS8Q,_^7I@=b8WSG3I\daT)1dMOfH9.I=(0+][0;AFRQgL39\=Ld<U6&J6
[&7:Q6\O[V7;5NX5H_Od;:a)c4ObAcV0AEf)V?_Pe#J1b3U7+;9T/)fJG@@MG?J-
?UV40NP_WYJFR93L/?+()O@@09/[8d4B;c3faOE(/BG3g+E94<:I=9=77DNc+.2^
@&E/SEa:HWX9DA;WTHHE5R4YRae\ASW]59HVAF;L?,S2-)aAHS[JCBL=.EY34?[1
;/E+48OPF1Y.6=ZL:MYQ+6\:G:_Tf-&19-K<:Y:MMRR#IU6-GA@P7TTNR>L?H4_b
XDM&Y/D/9(b2OVfMU;/:V\8J>LENA<8;:IFR?RCZ#>MOSV]NV+I?)QU[Ma/>ZG99
6-e[^R\gSU40#@S6>Z1K#D1GZB[R)PBS97)#UeB5b6[L@_Ud\)5&>&B.)3S?LUaB
P=VLc@78K=9KM[0_FTJKI>B6)CNLWX0CN9_>Y)UaIM3QCHZ_b]c_c=3f_b0&KP6V
71[;FQ->ZRbdbb:175>2Eg5X;PZSRCJMb07>=P+)WIg+69=WcQc1;O4>;fP+(Z]\
VfcZDI^Pd<EJ&?[RHFYc1?@IZ<\VIF?BUd2O6I?c107(PUKF8R.0)#Z)]Bf,YD.I
G=+,3&]8T7YW.[eE]B?Q+1eL13;H>S.BB+e(g@MUbK\a)cf2X6VJ,<0/.?P3]/J/
gQ/71DcOPC?J_A3f1#\dgeFDL6J_cXA]a-P#S+VK#H.e^3XMA.D=,.1@CZ\L]f_=
6Wc=?=c96SV)04ACRMVd[2BQSMWV&X8JaL11&7efdD@@+@QP7W)N39K/0.cFAJCM
D]8LRPP,]=;ZZIXLE:Y5/B9#gK8.Q<2<)HfVe<Ce[,/F7R>==@Q#GW_3VCBe9V&6
JdAc7eML73N\\^4-L8?\1P+bH7HCW3U@gCR+?^_EK?fZa?A/OS;fe:\VA0U.\&-W
84KJ.)#R&08VDa\?UP6M(_HCIID#WGS7?Z10KW-Z9G=4Z7B?..0e[.AaV4CK?Y1.
1@&E:NS#]Gc])BS1)5Hg;^8d/L8@_Q_JCJBI.ga;I\/Be\/0#R:2fD.3:P&#7=;^
:&D;(&#)b(b]<X?DF15V2\,FLX&(=fe3MfD48)OU1^-GNXIc(OSQD#320@.BP@6=
5BTTWSeYX7WE1Vdg&?fWKLdIge+[X=X>SY=)Ycb6#eC/?:KD,.b^8[@E?&;DfQVJ
[2caGD1TCK.cH(1NdW55N#O9&<M0_bU3c0V@c+M;;I72g#E-)FW0GAdTJd47K-WK
EU7V.f,fKI+05I[1^VD0HXeQ1=cQ<5YfAS=E0TU-^SR:M;6GWMGIQKd+8g;X2=[&
,+YZ@Of/3J3\;;/WPNE]KV?QTbeGMBfe;]C9bVN3=AF,3DJB9P8VC<G:CPdf[dcL
\G3eDA=,=#QD>RAa7@OTY96G/9\\LTKSXN4U97c7TF#=,AX]]04AURgTK2+5\.L\
N2=GedTgB)Z5QZ>#a[G[LVC&&(F/IY4EB10GO)aS>VR4V8LQ-ZdQ^IQ_Y:Y6Yd^6
g9/AdGWB>XR=W5MaEKXC>,/&?TM69?U9,E4>fCBb]R:L-\DK3-F9L>)38<FR>9_C
/(_2O/f=<&K(3)IT:8-YQ.#(Z<,N&X<D2L>[O0?gAM]M0,82F\]A.4UG5(BZ7F53
egEI4?[0MPFP;4/\Ha[FEX;>:UV?2aD=[=K;^f#V=RAgJ6eSUg_,>ZbfECfMKH3N
0,+Z\FXT:aIE;>SR7OUdG:T)<cHTfDUI2aF0Y3G+.++7ZQR:F^L8@UeZ)5,>>d:,
[eb12MJ;P=-NFA=]Z1cDb22EbEO[9:9g0+:<OV#=]<c0A3Z?Ib6\WWJ:W]]PZ//?
2D#A(P]M/b9XG&W9]02>K.7IUXb?.dW8dJecNN\MD5EJK+Y<aaPZ45+89VGA7/4Z
3g<eMF8/&(WCYS=PCCR.dNI3:B-7[&&M(TV,3QI0dAF:\B(H5+;#aBC_7Gc^DUV(
08NV9?0Ca(=TEHN:OR=(9FEM.(=K1G-&]IM;eS+;bM#)KeIECg/@-EBb_,)_/7[d
FNIX;3NgDIW:8P<-&PcHRI5Z#;>Bg#H<gAeEK&YH;P1.)G[CA\6gZa=_7K05[g:Z
SG[06YFOZA\Wg57S03F7.]5UIeMK/[^4V>/]c:dB^C;b,J5>.UNOKWN@:[gU&Seg
I0dWWfBBeAXJBP@fO[fd-DV[N>=[(.+A;XA(<-U5e]K=<]Be?46HAK#C:P5[2L_S
0Y:e;,;WM)+[&+K^_VM5OXZF5f_@^FT)SZIA[Ug35YAD<:@ORRB8[c9a@STe&=9.
^6N_].<0PD&/EEQ]M^dV__dV#3)B_1JR[)dR8A;JNBD57H>eWKRUH&KAT,U;1@9c
VP(J1SLWV4S>cD^1YcTO-fE_\1&cO\8CDXf^6FBAaFPS[&CN^7FFaB.TNXR/c:0#
c#J;=P05OdQ4,Y0N(Z,S=cg[P39J0g..X=aAX(,bV+J#^RTV^3g@bDSSN+7-)Ra1
9gVI&7L&d7/P?@E,MJSHQ4ZaY=##BfJLD+^C^:1;]8;H1VG?P[29DJ\dQK.Jbe?W
f/T\O:.]@/\B--]7YC+KI:(AOD/?=IO-X72;).:LTLF-O0XbKfYgdI>bc3+Z?6V3
9Fa.POW;JJd+/4<F90]?S[5Y3UU_&O(F3]M,7&NFF=F::OZf@FfH-O9b_ac-^CN9
+VJQbT5;:^3FU;@d.O8W9C+geT/&C#<)A]70?@@O<.IPBIP>4X,VB<Q#UC\/K#HX
,X\g#_KZ\V)W_Vc44/E2N3DQ.XFKS[efMY@X/GFV6WKW=>2C=ac4Gb(PLcLEP>8R
@OC;LA2/Q917JJ0C[]]RgP+H(DT8:<_V#TQ@HCKS6#=eD.VNW?R;6bNR_BN6>dEc
#DBIYSN^2U2EL)g7M0F-DSRfT,g6YBN75+VD.++<@I/Se/OX2L>BHcfYC^,SNceV
2V:ffT\V-PVRD@RFS/.5V1V(75;b+A]E3,>:?^fXa0VPEF8?K5d4E5SP1(Ha+37P
81:eVIDdT7^Gg>YJSA#F6W2V1,);6#WC=Bc@R@<:7I&JUI7eMS,RPBO&,AJc6=1Q
>KYX7./>W^g/ObNG:f<E+[1b=<6X=9XHM)g/;=D/X;B\?d0H@3N\24<4+IU)7T:Q
+C<Q[gH4_GQ@(3VV+S+dG<.aE\],.0X)=LOI1:=8c)f@NI5g-09QC0771f/TEcfe
^34W8PV\Ub(.)cK=ac7(RV_0GS8SK68SSS/Cg4KZ]HUOfF[/e96aLK7SeUC)&,0D
RABY8G.[W0@SaQ-PcJB7.cRDaYWB=YPR?OSWZ20BA\LV@c1FBT4\#[3C<B:@aJ_1
\PTL<KK)a#+b^NeRDb^:GNc7K82Df,3R6a-L=]H89MUf\0OIO^U[^6862f6@<a.,
beOSaceeX]3_OX&==HXU</8>b1YEXXRb(MLca:80Q^>477FKYF+.g3IJ<ORY)+B1
-H3F>:VPND&E]-.7M:M,L6c\OARS>OF:f&XJEe8f5+<@ESU^(8V6VHTZAa[]?@Y[
X<7F:])U0g^BR6&0IM7]A6gDbb8C(5#6??Y^OR/)15<6cI[B2_+=U2E:cO:G56?A
aaNDP3&YG\_DW6]Z.VF5,>OIg4GP-C,[GAVf\TA]KGHMH1fKI[[:J)Ka#2Z7)4C,
JKf1G>0T<:U+e9UIc@5S\Y(_PIW9+ZVW;I@QUg^EgFCIcF?8R]b\/8H)A8LGD;8C
E<NH]N-,IJdA\Q2@^;^IN1?_J3J,I0#CYT\0QS6Y-S[G<FCH)3:-FYK61Y<Mg9-:
,+,/4bFS^e:L1e<Y^9Q&QF9(>ZPFO:N:da<&c98^=J][:RZU#S?bH/Z8fCB-V_2L
2TJJZ7W)3M2PfLBNcZO<)XYF.YCV+OL-)T9dJEGN0>EX=#NC1^a.K4g23UNPGb5:
>E<;F[SMgQAWdC\4H_UE[BaDf^RO,1<;?0)B]aXXWcG&(E:7e(Y.(gdRf8HV>AeE
#bW<LLf1&bK)5<TWK]GOG-\,QL\DN@Oc7DYVV+THcR/JC^+faO7CTY7D&R^bHgc(
WQH^Cd.V=_&EcOI;#HO/&Y/(a9,&R_VOb(D4=2.EB?.&C7_,7\_gB+G&=[#gIEdD
F#C1U/IH81,LdVcA.1ZW7OD#)PcN\61/4=MEd@T\6=99.+XL<eJN>3W528J:-Y4,
L,-6SKB:UdH?M2\Z^[PKc0CbSNBLAF^QF@aE:,<6JD69=4T?MId)#Y_H5eP8f3Gg
BL8HG.3RFeUg8I\_0\bNK3B(U@1N,O=d,&9/aSV++(Y5-d@)A9-;Q\gb]9LG#5T>
:6TF#F)VSNPV+FK3P/17ATK<BRJbX#36@K;QBea)[>L0A5:gc_^2.9+?>H;ME.PB
c)EfW,gfO#&.B-RW94^]]C7APO@Xd9^X&0G+/?aKOEW+B,:4;/-+_2V5J1MaT))g
\@<E<cP]&Q:UC4L)YD/K&\Sb?\23)?<1=Jg.OCY<cSSc6T1^ZE3E1NZ2a3>H-BRJ
&RH4R^R@6TLT329[D<A3C1<fYE1/^<>Q=GU981-B^J=eTDN^&e=gO1>:K=O1\^.c
^8[2PG8P?S;G_\9dF<;<AOR6=&8^IAC>HEPUg=Y.T^DZU+d<dOf1?OB>NT]7MWgL
EFLO3dTXMKRd<BOM9H2<dN-,(?@K#/\(c#ZT+7?>/^2:Lg?T7IfN28ALL2?c@H/K
a^775FX87GJ(_KID6KLPG7.2UMCa56=.;;F<4I&)C,&=0/a:6+-KB#ALK$
`endprotected

    `protected
LKgddVPXa+S:f8FHa,@a@TE6S=)>4:<3b\_:Z,-K\C<)Y>8Hd_@W.)ST[GX+A@CI
T2)+9BBG=cUM5I+Q_(820(E62$
`endprotected

    //vcs_lic_vip_protect
      `protected
OR8A@&\?[_WT]@bY<d=9XG&G>JWa&WWKCC5;7GMU?g<#UW-?R[^D2(N7;\JK),&L
-JYJ@>DZWAf=Y7NASac_R[VRW&^RL&&@NE,,eD<[XF&&P>V=UIFO(#,c+48L6P8R
EU+TL?J:-_?Ec^LFI@ZD3Ca2ODf.KQL]EILa>L+_P5(^_Hcgfb\d54W(,3E(;0,7
+g1](dV;W,/V-685:0BV_KJ2\1Qg8.5N8dE0Q]M9&g/^10X22KBGF<0DVWH1:IN@
KQ<HY0PW7N>&f7DV()O@VK1D0=-N9XE5a>;#,0&T:.H+AbB:Z/-Nd@6I-4\d2IfU
bQfRcW@<eBIUHfLWKd0B3+N/g5;T(U?+N;c7+I\[Xd-TZOeILGV305+M\A(&(2F8
EIV^CJ+BQP[WAWLa51#^K409\Y0E,I/;0(3WVH\07KU0d;^Y#b=,_\,RX>.04[5:
73DD0EBXf]Z3OQ?5Xb[^gSI,C=FaRA>(>H(bWR(X8&\TLf_4)5\TE.AYK:g^R4I&
HXcU6FbW5Q&\OO?O9;LO#9CAe--V75C:NXL1=eW[#?:ZH9IK[.XQUc=9bCD7,9,M
0>\T:Qe2Rg7cNFW>)O:&Y\QF4]LE^M;dfH<YCE<Cf7G+JMC9Mc?.PeIB,T5;BG>>
B-\g&CBSO<GAWD=4&?Jf[;/GEa]1;+,KR(1f(B6TNZ-75KK:S2&U9YS^74<;6Z&G
70I_76HT:TCR:)_[G6IcPDAd7]VX5^@d#3M.SZ0eWF5@K>8b7QD-45G\K;<3C[f(
=ebJa.\9DY0HI0D.T1C05COJ<+>DO6,.AcJUBNMSKUSeI:ZAf^S[E>dA(EKc?-5;
6JZGU<RU:X2ZeX,765-V.B?8CYY)1ZfP=JKdS,./1I,I:A&NB(=)?JDJD<IIHAG6
3bDbFA0^f7\gEZFUXT.&#<b+ZFV0FD/(W6Cf<-cS>Sf8L8YEC[11=3]QdV-ZV,4:
5T0O5)5\7ZBD.)c+g\L5KgH=f.00L=6MYfKV\.#I=G1#GLH2\K4dcWZg9.YZ71=a
GNJGeN<K8NW4CV<0M0E,Td0?F[g.Y@(X+M)UKEWT/,,7OZL0TQPEANCVO#0\9JE8
EY#0NRaS7fSQ&/NGPaSJPM-)7GFR1-KbAKIN+,43V-WaXI6W6@Md:@IB/bLMc&K4
\60)S<\aDN]c<=&LW2XLJg#)Y5UC>M.f6eSB^a@12O^e;0_8?1-RV/OM_a+<S]W0
=TF1SPWGK@QRfd?&5B5Ig(#-6PX>>d(]HARVJLT\_]4KZS_O/9FI=gYT281_E81\
&E9>9TeAWJUb5U?cJE>9IE(Y#ZcORY65,>HPcJ(PJ^J-eO\^95L0S?9WU+)26X2;
JHaGIXC2J58^G1aNV3<N1Fg.L;X]@b3&g7ES2_3A@GXTVB.=.??SRf+I#Xb3AWeY
E:N(2LX0I\LOXZ]f1?Q&C&Y)Z?G0&.[TRU1C(Z5eKg64^(9Q/5S>42K,5E93ADA=
XVefc9G=dN+,?De8COOa<>\+R0DD)\..2+Gb6XDDJ>;_+Y>#>LaYOKKe;38T\Y#d
8K?e6RCPa@,gZO@JJS&>P<]8&._^8_5e,F;JL[d-/>ZUe8Y_DbR=(.YOQ.EVP2C/
b=S]Ia#?bcdO([^:cE=GXSZJ1eUIMF3RMOeQ3eCR#X21(f>(V0HGR9NPKC(^S-G+
EQDM/Y.&/>&[03TL2.+ea?dI=IDTEF3ba=Q6EC#K49Oa9;:>1-VY;:dM<QDX,_Jd
X/U0;E6g?=IX;^DGQFT@)K]I>MNP5(0K@?f,1E<Nb^]X)4&TIRd0RJR:NdW50/f#
@MK+=\@2KLJE_:W+8R060ZfW-S=e:Y@MA[AVMf^0\PMAF3g8,=Tc>O)RT5KMIP#P
<7)Xf84J@FNVF6Q0=VCDK\8^bW2T0,VNB:^(,#Y,H_TP65^.@=2?+OHM-7E155d6
GE<V2.04NP8MX@ES<-c^Y^4Fb-EV-_/d.M)=JGPFYN&c+^Y.-9d9/CMB_Y>0A>6N
bD1fO+e4BaQ,RS[=Q1NJQ0DRfQ.aS??+b2QJER:IbO?6-bE>Z^@N=bP,:R?]#(4P
0HFY(>]8(#?AY79L;[]N/55D^DLA?Ld474>KR_Wf;N=4[4<=G)S<)dJfRXQ-OK4b
E2FSOcIeFM3AM&6/@7CaIET==eH4\f9WM^cI0K7<#F6=4Y7QBcG6:9Rc9?S>2@9]
C<gGN30?gAFFd#bM9SQ-1XM=;ZWW0WZH=#9V@X.c@L8#76MQa54_R]#N6=:&L.#S
MPG8#PX4G_(\#WI_X^cPI&9,U1P:UNKd\=EC3M&/5Q]3G]ZT@gA1GFG0]#DRaT=@
_P+#D5(c6QX7@Y46W<(AB^,K3Bed<=AN_VYdF/OM:TI6+bLHdTI(A5.HXe0T>WK-
9?^M?&<)a<PO4J6=7_Vd=1#)6RTcYd[;.1?]R=[VX-90dea0=GMOYHfDXfgFTY1@
0Qa\F\1-^;aI)HebJZ=7>/K@3-fO;,,84P;#&U34G&I6Y0)cW#d/Xc:>5-;PQH-9
HE/g)VIFYW[&Z3WE4.1Z<EEPK8LR,dCA6Wb7BUP_]+ST[)6aVUNI/^WA533^c4>J
/29;.?8Z#TXQC:;WgS]L)e]g-6B9VC#4C@faJ2^AMKOFVbb&K\2dcd[E9K#Xd4]g
E6&Z^NK2c]7>8+DK-L<B?(_9:c=X)YT(M)KVMCLW]F+?X@R9NNAg?WF^/Mf?6@5E
W<aTFQTSA_/=.4D@ZK2&,<;b66X3/-O28SF^0^E6D12^DKZ5.8_ANW75OE\K3:P5
Q6Sc0.EDP^6_X3e1DcH;7b/]U-g(fJ1Q@ZAI2OPgUPRNE+@47N)>+gf5.Y+RMLS,
Q^SfC(d28ZOG?.RD\eK[W?)@K\C:]93/\,_bf<gP>g2F(d?^7L@6^,O^(G<Z2Be8
/Z^JV;C>;[;+7;8.T(cRT9.\d?8#TD^QBK_@Q2[f&D7gG#CcTAUC>aEHXM4:9a<(
R.W6L+S&75c5EUL1IPD1@:F_X4&<Cg+[Me?#7LD#EF+GCFb-D@]MaCZVPQD44]_^
e+>E@.aJ/bT.RP&044>C5;.@<cRPYO\9)0L(F&DDM;b?-QgGBB/&>X97=QAH+2_,
#H;PU0LPFDGSK<Jbc4c)@MaLVJSWJab4BF(O;IBC2B\;RNMW4EEFcMX]+.(?2>F3
&b8Pe>]B[K@&gg/Qd^:U7M[F4O6N@JfL:.9K:--6;?8U)7Z^KAFS1V9V5&MIWa^Z
7039;D6&4U6GX/W]T0K]fJT)aC2)-QQC17?_5NK3T0?2:_])F874537U88=42?.X
c3N?_)Y;^92POdSdgX_BLH1b,W:;WWLdNJULE;KBYH(X7F1ZCO_F/#<:1@5a&OZ[
;9_)=EVP>+f\=b>^#:SD2Ld2)FPcM^T@)SUTDIUYW4H0HY3TZ4Y#N+74,7A52VE,
?cIC;\TWbd]0(9a+F.Y5^cBUcDUfOFE;RW+1Q+JCWCcRS.CT#=V?/^C-cG+KbgTQ
1fHCeDI+U)WZcObS-]_:98#9aeXaIX3\BTQ2]LO&F](\R_<W2<-eH5ea)P670e?E
^7=E@f&XDb?JZNfS,MODK.G+X@)7-/9YJ1UVZbH_HCW_D#ID=bd[,KE/\):Nd38G
21)b+/cLD6+6Y_M[9;DJW>Nf0[0U&^F#b0E2FM^)ZP+^ObCKYZM<__Z2?]d5V/-E
N:-@g;9f#7KYJDO<f>27(W0RLTI+I@UO(Z78.L@Q#Of6QH:d:N4T@\I,)>^ZT,bR
]NaMRE=U&JeFBGK,\=HO(g9e-1>+2FdD1a<<D.UX8Bde77[1HK.9\#+WOQ,A0EA\
(/IC<K>V4/a0JRKJPg>[f>-Q.J4:W;F/OIA.+01#JR+;ZGR6R\ND]:7SX0c6(:)G
D7MP;+]G[7RORR3?0aQ[H6Be-RT:V7WP=0R8U7>4cLJ;)8dQgJC-0aXWYI)KZ?@)
BJDLS^IUJ<SUAgCY#JQDW=R/Oe_TG<)aFM061g2_C3Y9N91.3?]HcPdR-1+@8APd
E2NfBMTd>D+0^LV4&L3XIKQRgV/PP;E76T<3</D[(O]/WP:&a-]@T1MNOZA[L>N=
G0:04:@-D_<-)=H?^Zb;[EZ_GB+@-\S<=DVN<413>/;L.;:G8J67@gT&:2L\\G56
S5P,]WSd6[7V&&f:^CNW?4LBDQ=&d>;I<E0-LM^@DU8]L&[4W,eNZ3;):F)e:@5-
H]T:9dg7_b,YF293J7+Z2CT/F6W,A.[G&@99g\,O/fcB;APcEUKQP/6^5[IO[RFM
UD@L;A&(5GYH:O3Id,?d2V;(:/da9fRf_Oa-6[\gK-(I79PB6050?5,>.4=DQc/+
WKF1d^d,U1H=?5>gBPC?<T6VH<dNe#Y6Q&Q?:D^HUQ^S^7>VHaYUUZ4,JY2HCa/B
CML_18G>VYFS2#:V]4Va((\ZJ5A^&8c7;V=:5RQ]NCCO+#WYb0cG3GP4?@FI1=FO
/[CfaE0LeR27WBG_Y-J&ef)^W6FV1;^&4[-2Z8H=8:5OX,PW<JB)]5#H@T+O0=KU
eYE?[)J,-/F@/E2O4ZIK[I;21/UM=+8(YT#@O6G7,P<\a7?8c)=SW06e(^4a@_^)
;>M;#[,;=\<T\))g_7?7-Z0X+WJ;07HG?b_#caYY^cV[MDN)3M76Qf677I?Y()JJ
^AIUE=cT&X,6cJSUWg)WG0ZR0+VI21BEDEfPfJ12.PI,ED^JMH;RHN]Q(GHERfS5
9YEdPeY@?DH1/5F/b=,S74PGI)d?C#3ZO9HCI\A)3,8X8JA:XL;:GbSf\N5>O]J?
bP<^](63K&N9;I#YaS[af3.7UJ))[BgFd412^_B)SddK8/c\MIAR^5O&O+PUe)16
c2LX@Wc@NVPDA.+Z]I<W3XOPDaegd]\(WHOcIgGd5<?TS2c11S3T4<[:#f;X<+3C
07N2Q/B><fHCb,U8L:?Y6WFNK_XD2-ME0_[fCI0X1+LJ,:\A7>;TcSd_:_.RSG:>
^I5<1Y1g&<7:52BQ6a><WEGg;I)H-2M]2R;P,dXHA]18KCb=WON[;DeLeV5BAZdR
>>b?RKd?N.ZbK>)[]9E,L\MEWPF;JW(I?a8;C#?)TS>#)WS30L@4dVLUG6H-,NCd
0VS<L9ZY,_X[f5,MP70\Id+[R_(_H;<Y^ORPTAR.Y3>[)FU(_H;T:T:d:@0D6+cL
PdLeAL/c0(@53BYFW<XZ^G<g@XSF?VH/-P_T)OG58d]HK-&-RcXgRKDeWd&g32O^
[J0dF\AUB4E[MEPeYB?feaCJZH+aAb(FD08MI2D:MBE-GLUg:c:Y1bPC>a+<0S,_
,/a@cIQPeG^e&K\OK05dK>=#:A9JV9EXBbDC841+^-A^@V#[,/cR::[d(RdC;FQe
fOYXb0IbeOU.LCJ9E.fP&B7>+6[3ceTM4.;c_gY<.UK0CVO&@KTGOBL38W]QVYAE
_9?GXd6F6CI#OWf[9CeR#EIgEA@XdPZKF)/5F<LDM4VT_?D^aQ)L?6#T(WfFK&8M
U#a4G<:&SQ6cd;fQ].TT>=U)g,Bc/aWJ@edd4EIL?3^1SVAJ#.BVH9(^36)<41Bc
5BgQ14C#25>U@[-fQ2ADH9O_9X/K9b2,=BA?])8=I\]QX?.3D.ZUSG+V0Q06)UT7
0C3bD\MH=fBW/0L\e^Ba/&HXZO[:IH3Bg6AUKWT[Q5XN#3I[:d.)O\>1,_VdNX7&
_V]\Fb:_8Xc+:7H/V<1;:P>6RF7^<J@fP7E/I?H_Ag/#710,K[VDf6DYaYK<TRE,
U^A5?9XS-[B0EY#I[@\O/[Z)Z\N?[IFcDM7@+ZZX4Z^81&4)];;=1-2JL+/B>W]f
P(:Y9GZX/@X-VgZZBS@b&52YSaRG9Y6T)Rd+9P4Z)P#;4N&=25f)0MGU7HF(LH;<
3^[J0Q4]^V,NB[LJK[(SJY2Y4$
`endprotected

          `protected
bP/)a[:&.0;6A92[0g0f]CQ-,bf::6)_ED[AUg_B4L-cc:Q1?e0U-)+)c_&1V]DY
(c[)Ic5\fTI@<1?ARg8#\^VDQgeZP;],M1ac@-b>Q59M<[6(4:0?]>+)I$
`endprotected

          //vcs_lic_vip_protect
            `protected
OL:UC:GO<E-KVBgA@[J[0W?N@c5@IZ:Ca[0D&ee#YVV\/CHb,>251(BXH16:2ccQ
\BOQ)>ecgG630S8b=@5EHVed<T#_LRY(Q#0(#5bNPS=W[JVPAg(2=V8>8#Xb&-H]
,,b[GK+KWEL:^EV\dMe/2eVbC59W/I](WX+T5#GA[M\G9:;be];>UMf+U8N?X]X/
;SCd.\aW]<JZ<8S1H18TMOabXb>^H>&#IXHO.SJH#^P:c6S\0.cT^JGE<Z=GEH9X
].Z7DAeZT;6B2)f+)+)6[:I8?4ZS)/B<TO=>2R=N0SHgQ)+Vb7QNUP(HYRCg;#A(
^:d3LLZ-9;H8GK74IKdPO(;e96UIO9TZ;4)BB-a-7N18M,&&8a\^JU&^<Y,(B-5\
.JFR>;/.)JESRB\9H<dL\5U:,Z3[@-)?GW]&^X>Y\O1M_gRJ^^<NCa2Q5=THEU/X
6\#/JA8(eJ8.DFg&&gZR4=_e(?.?20EN\M8KbG,@\d;VKfF@B_L50g3T=E)_>,.J
g-cO?dg\MgCDY=EZd6K67aJ+,V2H&_UWMTaNZKFN))JJO41X<CTWJF>B<6EY(.K#
ONCP[\A4Q4S8##c)eUeZLL#a_2B4Tf_/H,URg6CFb=.KXf7KED-f-8(B?TYYbQR5
^Xb>F-a45b<4IO09NLY+^\F:^(FaJ4bH8IN<4MLRA17Q7UAc[)Z>TQXOX:B61BRE
=->fb5#>Z,Dg&b[g-9gZe:EZ)MYY(c8,_EKFaOKS<B(WMTYJ68\EKU,X:S42BQR@
,UV[F;;#97@\:YeFDV3QPH^NCLE858393FVID<Uf\AcZ7N._::3]IN<&Y?:2-BK[
G-KQ?9DTNXT>J0G#=#f\EGda;T(9<1Gg@-FU\7>&g=6PR72U+7b@+\XWfb7943OF
Q@/VHDAdgJ\CRETB[VIQ]ff>Kbc(ABgB\(:OE;O</J/faH\3)^N0[a4EIGIOEQM@
WUG8Se][@a114aW(B<=CTd-2Yd9]dRN43=;7OVL.dPR:d@^3_dJbc4WO+(?(,ZQ-
^fS;QL^1-5Sa)(\+d_JQMI)0b\D,@IfL8^8E?>gWIa]ZSad:1[3B-D>TNTX<5Yb<
1TfAX8SNeE2)8X^IbF7^c^d3H2XQ?&HLE?822[\ENYZ2XVC/Ofc?V9eAYA_62CCF
&(+#99;7N&00@>aI-6e8e#F\[:ca_O:ZMCb0bN40>fI@OA]>TXb545?]LV62dE0>
WXBgT5)&dQZ=R_<\O6a-cg&U+PfE9\(2ID6H;90:0T1N=;_G]3.G?,6BV]-@cAEZ
XS8WE=D7[KJYW_ffGcYOCNbRE^-0BV<IPR:#KDC,.F^BG=2D5BSNP^bc]d4C66D]
5_U6.NMHIGC6g5K>W?b\ZTV\&ND.S6>DQ8VGc=aU@_+2@RO>)UVD@F9@cO\Z>d-C
;/&1aQ_CM(BMSQN]<GG)=JEe/0bZVAHM#5JH]<JK89MYC1M;Y016Tb:;CM9>dHXa
aZZ&;F01UPf3(/ITY=I]G,3EeOCVIG@.ZRMEVT<B).Wg2\2#.f?A,b\]]G4D483,
0.fC44R;DcO;Z\;4G##)JX(a34Y]]?OSBEKK\:BUY4b+c27:eId_3Y?3M-dW0_(2
<?ecNb[_4D+SbQefN-.cABI4MXg91/JO@&CM)D\Z3WP];;NTSd55Y#R?9A#QFDC#
b_0P=#R8A5K2285T+>0__2aWEXPUHO@8]KR9N>eF),V7U>NZDG).;6^eFOd@5E\8
6JYa/11(JXOc-Hd9.FdYI,4H.)Gb4R/,QV:<fb5[=aH5MD(OZ2S&_eeH94Ge:-<\
SRX?7g26a.;#f7aK8PR.^R[###O4):)]NS-\-G]ZOc(H\.Q[WVF3L@?.&,b&#C5B
OPP8g7P3+\aZNWD+_1YJ/QQE;Q:Dgc#NS&Db2C8XUf5GTaG[,g\7_#6_-WcTEWG)
NX&-]+f6OL,GcD<4L]>D1_/BDUP+#SX6NgdRWA\HFM__R..)^K9L29V1TM^O9S.B
+LgCZ\A]61.@OcTP<BgbX=;+c]WNT(/g(0Y[#U+fRD[a34_7>XD7bDH3M0SD:SYd
LP7RI/GJM@YfdUAd=(cDVT4//TT4EX:;4T&_dF>I6_M+0ASU_3gMW7P_^R89G4<J
.V?>g[9JBfc?>GR9-XFaZOJ5FgQEG1d;U/[Y;AaP<2J]aZ0gE2=WIDHccTa(U5ND
ZS??^,>EJ9&\dHU(UA0]Z=dJbV..]WR>JHB5AA-TRU((E^:X.OT8\Y7Id+<5aQ5]
R4cT2#<H_@Z\^a3P.4<SW/[TFU<TaJXd<H&G^^&d];I5WUV8:Z3M</f/Y,Z5b5C:
=F[W)(-YfLc53d8LdKOK]UPWc8XL\+-=1J.873CLFH,dJV#d8?_@S>K,#@EEM-XS
><-@]GIXPR/E?M40E3C+/)dEGX/c/-0R+VNWc[N>9@<EU(MNW-a;.X66XEZAAbM2
<04:-E#^_POA4b_aJX2\J7JOeS/FIJ08;8RS<#HPRGG>6G7G/FIQSTQ.F]QODd+<
bAE4MM&fZO]IaN#7VXSK[TDcfJ0ZRSN0\)6Mc&721T5(/3C;PC]3>cFc,7#.[_>C
KgMg&MP4\1aL(LJ7_JK+L6?U&\0P,H^#0SEM02W1J#8?^9P@-3/,3f)98TM?YgSG
)X0\81A/\[e,0A;<8V<L=aP^P2W-J2UfW6TO8ab=70;4d)7JJ6KTSD@CJP7ACdS,
cO84W[[1+8b:Z:UL.IN>P-c0A#8VK-WWZ8L&b#]&YR6S&<+_bI>fL7gL)U-OgaAY
V?8f0K^,9KTE.BScg@eR9>[Sb5OY\+=<BQ9I/@fZ?\BT2.HfW_60J3C./bK\3S[/
TUMA&#T#G#95(Y?ET+Z2I9YUB+\)T?I;KS]DK,+cWUDVbRJ/2PG5d22PbbP2)RZT
C<C<W5S2YE7D#a;cgTI9OL-/0g6=@7Zf3;/,gIO(^X+790-FYFG(.a-S^.(-D/b]
6]I<UQ-HOJg4RL_3F4))aPMPO)/L@+9LMfKcdNLI/O/0\[OMaY#ZZ#.;\4SWe[4\
gSD9#JW<F]4O]3L8c,#6LM]_)W0VWf^,GK6_bZ537YV<L0dU>Jg/.f9A5+YR5CI(
EgaQXDHcHP1#3S..I0HS0\52c(#DI)a(ZC3FKNQ&XgceE04-3dR8<C&L,7I\7B0.
]Q)RASNG(a<G:DbYE+&79/K&P;(R\77KbC36]V8X&KO(QGBf_QBfYeD#.X@FaOPN
W)>-aW;?04ODRI?6b;QA.>0=Jf&/YO1VCC:7-7M2_]KKVgXPNeZ0Q7:&):7G\g00
:/[C^-@&P/Z(B=>0c\-]4IX?AFdWS\W]KeBd?-P?E_;42O@KaTb#08@D(Be)A@X;
BgZ2KBCRSEUT;7JbW<KQJ#a#Sd(C@R[^1^@\?_@<IF\eYD>g9,<Q#@bb@+,2_=f8
ZdXf\@H4:9(97[2?g5dO0,C9#N&<L3>K2-?P@ea^US(#bf)_:2<)?f(;@W8HBU82
VNLB2b05(?:3OR2+KX7gb&,6_c61Yf14(.0\GX+<0JY_1W2;H#,[7DEc0LXeW85E
^e+>Z8SJO;>4KEC:U(M1KT)K9?\7@A-]<U,eg)L]_VAF9O>>P793)d^#Y0;L=WYI
XbJ,eKXNKK,M3]+^G+7KfgBH,K.20:>gL4KdNXX:L3O9J#?EPZfKCEaa-8c3?G#R
D1)9:Odd3=1NbAYWWa>U^U53^XMgBQNP&,Z/BC#?=DI5]9bIH&a16c&6cU1#O@7(
KCU[RQ,7X4U/0L:1S2[721PfE8S+PS)+@1^B_VG56V0WI)]4Kb68MMDS98A[F>9g
#b]+TJNDfMLgF?.6(2_O=\;1(a&#=e,DHe2UA[[V.F3WdMR3Z1d:NNCX6&6+,]fa
ca1(R?.VG\>.:?I^&X3^7^F/C6+S/c?NFW)\K#e\+]RT91I)JRY\,X<=;3#X9B-Y
^,V\NIYa6@J6H3.FEDCS7X>;U+PXP&>H/\)PZR3AG&0((<\.BH@1?Q2HDR]dYTcR
D3.,.(=+OA:^WLA,b\/;[H1U?\+96[WPK;>ZV(WC_;QT>68JL@g>R_B9Uf3de?Wa
5S=1T+?22.c0E^M\@/TXD]I>VSeDHbONeUOI<fDO7:0ZX=9LE383-]&3U&M0W_-H
gO13&J][T1K(ebN_=NZVICQdD]7LXY@CadRfR?>8:O-8K/R^KER>Kd)dJ8.)_ZNB
P.TYe=7\>)P4900gGW9O.7ddQ(6KfA@Ife?gG6^IX<IM)1\O(#\XP:R@#XP6C(AW
/6(9YP5e:5P,(]U_-B/5S]@WaMU;OLc4?7BB]6=9A/4>#ZMNPcBN1a77QHQX2D[O
J7/DQ?IS]N.DJGXYI3VVH9]X;I^FG]U;SS>6PQH?EKQ75-)7c<[4/Q.54CXC+Z:/
&WH.VC;)L4_)E(1Jgd#]JW\YGV[3&U)2RAQZZ>N22cUe^M)ZY3/9)-16+CXTT4=E
HG>.1Z_9U-D7HM+<\Ea+KE8KdL/KM;\]HbB]@XcZ)2fObZZ3O6]CH^L(PVK,,0:(
V+:+THHMP>I]??Y50RO#,U+BC\RVLN5J_><VB5Fe644EcPHT8_@>_G;M&BD;6f_#
TX+SG=U?\CHc6&Xg(9>GPUISCO>12@,QdK28Ee(8;R8W0F7V1OUDQSU>[PKbM<.K
c8fd1(fH7_g)2/S9a8?6>d#+;L]Je0:F7:TJXIb[3BIQd+1FfBQ>d[3+IJZ&E;d.
FN,23Q+SL5;B)<:2#/XEAd<\agVTI=6I..O)E/eS^2DZUfNcWBZ4aM6;gNI]+Y2D
E=6&[BHG6PQ3<:f:+I],YAM,S9F-7M5Df>aS?WXIC,-X,gZ7L^U+2:LU0O0HTK,S
?Z+?NVg1X7WA_D,;Ra4[dJ^SR[WRXU#:GG_g]:>6E-W.e/;d9?&EXO>R59,e;BU3
GFdH_@g0W6W&UC>,;Z3<5;99^;MI@YT,J84VG2\:dI+H6<2K=ZYU+6KEK[135T=T
I-?F=gAX+_]11fP=ZS]6ZPRJPURgMAYebf8#9ga8^1]7C2D3YA5K&9,U1^O^ECMI
5,Z/9fcY?=.R4/I9T?U24+MKN)OGQcV)KMF.A[RgI_TOR0?[I8N\@Q@FF^U.6&C4
R_SE5S,_W+[G4#YM-0R,&a#_,Zf-TBBCJC:4GE&B&UK);M_>ac.RG-)?f]1[N(TA
W)]>^ENCC8[H4Y,WR1J>_#dFH3U?.2H&&TTD3X@bPfM2<48O6RgIcG67/DV,BD[@
V4O9N>[Q#&]ge+(d6Z>?NQaFER=3g@GEc._7[D]9-/T]L[52+DbBScGI&E\4MB=R
BOG]IIGER[L<<N<D(e.8PU)J30[a9SUMa(:K9d2OK\M+751>FTe.+FI^TJ@WW^=L
QL8^Z&F72@3GHYURc+L-_<ZY1U8cWL]XWOTQ65TQ.#L<P+CdcR@FAXA1f7J9?S:F
MQ-_GSU3E@P@M_b4AI:FBbJ&O64K<:c-9;1Sg,(A[b#;8O6S&[GV/E>S1LM&0(D/
)@c<.I:YW8FeFZ?bNJe+;[XGDWOEP-/,^[Q=3?@=Ze<F?X<Y2UYbZ=7\,X;W^<dF
M6c51=3GRA+#;U#d7&W\+3KNe<b#GR6<QI<bSfDgFP[4<7TXO^DeA;fWa3/66_BF
7A#17NC_KMcF^L&0248;^;BVD[A+__B_-Q=P+84.H3X5(P2[L;1SGfJVW/F\X=<V
J<UM_^PGfR(AUNVAg+ZI]d46+c(f2HIY[B68F1<7,A^b9UP?4.KV_CJ25Y9V\1U@
JPIYDU99e17U,=;XJZYWJ.8/115Pa063LbW#XHZ9Z]2/PPM^]BL[#G4\Q,)WBS^9
P(eUeaeF,B\3NM1Y]&5@Ge8=D?Y[9:;(E+9.)QCB?T[[PK5U_;LZR0;I)\QKFT@H
UcXZcYeG@W5/2-US_7KZC,5>7FN&#+>b^)e2Z;2MD_1SEdb8T.K>fE);df46V<(6
(FS,-GfS[@ALS6fCT#/4;.<L881=H@L>3/W##W>gG>;?#UZ;DdaG.de?H(4LN0Y9
S/+G.gX&9aV8@HV;A0U8WFPLg#BEH=+d;U70DKcgZ78S+0EX:SPFDC9U^MESLY=E
#6[STf31@Pc;>FcAC^#-BHQ[6^e?--F;Z#MG,5<)6gOE7)Sg+BY665>:(?aSWQ+U
f=Uda=B?=MAMJX5,,F(YQ:a(/RWKd@=Z7DYcK:4V(QLGVK-PS2WZX)UM\>>.cTML
H6[-WU&_Q6_ZVgQ]:f3EV4a&)A-,A2Ge/J_c=[T&IA+:J2XJg0B00,eeVc=b:/BB
=RW6RJ_c\>Lfdc7(M\bQIY+bQ1&WSK_[YO_XU\V;J1TV@C:,A^551,a0FLQJe^Y1
We?YCN^1ECL>L&<ZfI,BU39PBa.DFfE;.G#H5f-c[&BRA6Mg&PH]_8I,WbB2aLOF
WadE/Z<+4ZC\;;.Y@d\cFFHRON\U3.-/FB_(_-XH([)Y73+S/3-)6KC@<L(f2Wf&
8S>c=21IPD0Z8W@1P6Ua2-VCeD.>7fNeEe^BgK[&,FOH4EWAe=G0.>FKA4AACG9)
\SEdHg0N&g&72@XbeU^4GV^?;:221[KeaQ3GI;<R_YXFLb8M^A==L?/3L6SXYD#(
Q2(G?NCaTQT->#8K4,:6D4Ua?MA(N>&]6HF7GF:9[VdJ+ce_1R0+1N[/I9LFN3:Z
.<UIFAZa6FF,A(H)ZBG(R^54)0X3K@3W(B2;=TGVVKZGc:E,@DJ8BWFH@3?9gcTQ
[B-,<MAYZf0?R&T@<#VDMIcbCe6W+G^0AIbYW:/6LF5Q1,H@Q&OOfYPd9=R.XOD#
0>X6e#&K9[@6NBQ4F2K>8RRd:RL?P.A7W7]9.>]X5WNU2cDg8F?F,FEJTHI5U83g
[aT:R^+PCY6+/_&)P;RNLaCE[g>J.gM=HDC8d6;Qd#HOYEY^>TQbKMVU(Y86(c2R
FZE\++;dC.#d+C,:;cCGK8M7EPCMJ,9H0U2,P6gKY5OeT](.>=]ZT@f6(MP6g\a+
B<Y-W@=N<?1M^4feQQ#Vg7S-+U3.F>302P+?D#g+dQBc[&SQ=5<)Pd,1NWWAGOaW
B0PS_K#\K[N+=R]HZYc3V;CN7X8f#_3QgC<VKQ-WORPGQ=K^d3OPA@(0dAM@)8(]
W9Y92[/9eb:Ue22#2+K,;?M,1]OO=Q/L)-UZF,ZdCAbPM8@\QggB2?)9>B?NY(I-
/?b==[\fN_a,YLR7@D?X\9-Ng32<3e:-8[_bH9Kg];aS:AJVM<H[b/?R83I^gCP9
E]\;@:OeY5.5IcVH:]/,+0C#[8A6=T]5QA@RHcLV\#;W>YN#RXFRK11I+J+H.b\N
L]/Ca4GdP+BC:CcOS9-YY,E^CVYDa_c:OW9I]K@?UOCN(^MHW_Xg\/U\MK<.Ug00
YKB]-JL,H5VQgdMMSNXS>)C+OZZ@.Xg,V#(Ed6IEDL9K/ge527[2[;2W=2QA4I4d
&9b6W0>W4>\L0Ag^AF[a_A.G08SK&fFDY4].^.DG>0=aEP/Ab4KKI[#cM,=6ZHG-
=f([RL+41^K7P=)eeL48)T>>B4<-dDQFWCdLIS84-L6:d8YJXefXA37.^1E@#2U<
SHY3Xc])ROV#a)IFb3&=C/>5[AT=GX\^:,^V#4F+@,KZ/M[153:&7+d^Ug(DPL?A
Sa):X#AJ[SVdGZ^/?/Rd8N7a+RBB?4?GI/T#CF-a;;^6ebA72YU\NT3\/#S.LUfJ
)B6?4;Cd]?d;MQ)-T8&&.Z<]()&G0dX92H5,K5:.<eEGWf2S46ZJJ[,&]_e0UN^;
\X:)bd[QgUDQF2M:<E?[QYV->GJ0K<-H?P@M>P-57LK9Qb<\L#LC>aSM?A>A&;G<
4I&9GRBV/V&^6D6:7Z#]L]MC2=NM=g&<]/0#S8,fQUU.N)dXN,.XS;ME(Xc;[@8,
Y0fG^LPI>47S3NK:NFOR\_WY))K-4682#c]05+Fb?BX@82W#7IRKL89d+;TX>gU&
MK+J4GTYBKaHB8GXGEX+EGQ_X9R]Y0#Z4WMH75OX&6).5fLQE4_R=PT,TB0.G-D0
)VB)L+ZW9?2#c\75_:IRIa5K)6@]U@g:7fX&B31C6CE)FTMH(025RE]VO0#+P7d_
^^K_Y)]725gMRS-[UIDEH9F^&I)R1NB4IA>9^K[\KTBD4Lb:Y[8&]4J&T+R9;72_
>9APg][>[;+c3KLW<E)V5f9_2]9b@^.OKNQ+=.7Q177_>ARIf89\dV>W74AF&AN#
BRN9g^8F[3NRYZ<DX4@XQc-W[TZGNG927M>5-PL9^UT?:XUSX?0e(cWEZCGZY577
/#EW>@LM]?b=B.P5fV#@1GW9bE?MD]/@E?9N9>T833OSCKO?6XYY/EPT#3=,Ja:7
5.E\Q&VT[d(ZcgRQORcDF][NAASM(1I1,]ffg@dgdI(24LWYJP,agQMG1T/UB&8@
55IL>3(g8_f,4I32bA?aC_<XHQ/ef4/c1eF/]S+RVa8[GG9=F-2WPV^YC_J)IVPB
NM6@e-M84D]CDHY-BUSDf.F2)R&/-<OMM:J]28,G,[P@ePFV]RXUYdD@PXPR:?@d
.M[:d:I(/P(:]],_ceWc2NC5V,/7AdgW>9Re^N;.VcR^4M/EB??CQ7]ab2CJWG.f
bAI3Jc1:Q[1:95[^2c,Dg\@KAJaa+(>8T9M9KR?+IPZXZ2XG()VSRW@Xf><e=0(#
VXVF/)?I#U-51/SFT#><.N)=>7cFW_:0UVZ@EbJ:M0L#GS@TdS]PBHOPDQP&QQC[
J0HOKT5O.O1S#[3bGLV03K/PeLb:J(T1BHV&LVC0VcL+B[P6M5ZgC<QC,Q3T8Y+f
N:8;J\2SFO2=X,9<]?=D)0UPS^A83g8#+0aRdDb+B1C>7LD-[eQ??69<XAKd=]T5
;.5(6EN/N1+<)/YGDbVHga<@@34BE]?1eZ\X.=]Fg5F#\PQ-MY?(5SgcUe@bSUe@
;2@S0-c]X<?^?2:,ESD@2WP;R@<13.I6.[,RDJ1BAA&<)2Y8)6]#<0+b6,7=]T4A
5T^G]bVd/MN>I2R]NR;a7G9EZ?1+>McC\3G3S9#+L?7J2^3-2&0LI#:A@+6XJYeb
Y_VK+0bc4HVJ#WWU/UbOc<Z.K_=DN[.+#YaH_:;(#MCW1d#LC;#f)<.18_(9=A8D
/F(TF:S>)g:GcB>,NQOD;/(:89SRBfY0>=;14B2?O5Y,bE)&QeT\CaSN\ULPX6IG
<KJP)BM_,KL/EH\Z<UBfF^(W_[:&3[.b+/&,]\e09-D(R83DFK.Ab?gOVGDHE[H@
[^f>d.4C0N]?GS;F=5Q8)#@d1D\b]^AS1A<#.A=9?Q:)PbLMLc5f6Af;CaXBZYE@
Uc43CB7RF-KQ;.+\4BeD\A3FG:<TagbAQQ/AH>[>6?OeXM]3Ugf0V3=@Ra9<9I&U
O5QG3;V];>-B?[ZNa8HF&J&XK>QNTAT<_HN>W]Rf&4Ke\^.V)9Da[A7D:9e:P4PP
(b56YeDCA\d?Gbd4+EUd[,5P,2LOTQa_D_aW?f6AJDC]gd@<(92BZ#&fDQQWbA6[
].:AL:[dA4KB/Z.(NTAe#<R/CSS--2THZbO;HKbc=([e@-_KC:-aZSH12_GKF6?O
6>WSeAI_BMVU0(F\#>9cd,7WLMOIY8R7O=SNa&H9ONCI1X#d5NFc^4^Tb9U<JW6[
[+@_++[QM?HBZg<X[[VO3NK.,f2dE\.0+b))#XCA/U>@,eWH/Jb1:fPQa3Qd0A1f
eB.aK)aXV(;3XU<GW6U&V/^<KAC?R=e2f-\Bc@I4B5/J)+#A/+I?WE_Qb5X)AcF<
QFF\;[De9Y#=@bFDO0#T07B/<3AW&=6M.-66^5FG<RYV9<ZFWfQSd6Eg60=2V3<7
0T((d:O&;QaT#Z)NbI^UB95I/?CU#9Z)4&8NC1XEWSgXZbQ0?/-W3Ig5K2SUEY^6
_g]0Q7)(@c3]6T2O[+>U91PU[<<ZZ;O2+8HCL]NZ@ce<Z7gSZX??I=J5P9@b8G+4
:M-WgS1CH_fD_DQ,@V/2d+FZV;Z1\3L90ABee9_K7Q7dH150:.>&RW_DE8R8J<[b
MKaV_]f)fg\(><M(W0?_(c\afUWN5E)W;7PL;;SHX<W8/G]LNDPKC[^^S+WI5CHQ
M(6-DGN68Z+CX/3:2BV>^BN#c2VSVJOADW08<4C_N9_J8:>@2-?C-@HO5476fae.
[JA681(6(N2H6g8[(be9Gd9U^BLV3?AC/,G;Rcaf6,(f?^>WQESBPEHg=UQSU9.V
A<;\=#9XFb6WWV8\;Na]]0f:/HBG>]:bGSgH;K\\,MYZ]#,LOXc)e8FNR-1Ub:F=
<6+EaU2<].-J:Vf9PadcN8A0dC?Fc9A0RC8ET2VfE=0@&5fA-S0\Q8ZTaC3OV.=Q
]DcdDT&@7LFeHX;CA3I=)FQA&N&.L_\M4FKNc^U+-.&RNS#PKe2/UVb6]0D#&-P8
(<:eCL4JT-O)J1?\gIa&ba)[^EMAQR+8UYDVT:c8YMGS&8<[=FCe-WT9N)8H7:,8
<fXD4Dcb@aA(4C9G;VCFI[SPg,NYWSBFDFD3SPd?eU&dD8==6c@\1<VG<+EJXLU]
WMVIYLE:#bB]H0G&A^QSg?+S&C(3P0]f[GF;F<c3-[ND83Bd2318Z/NG9B-\D9UE
Zf1MDWW_O?S;/B-Oea=KK>F;UgJ##+;L<_L_J5/&=3JUbO4P#@A-)gdZbOKVg3TC
Zf>71Rc(A#9fM93^d<O/J==JNQD29/>2G?<96fVV[E_QDZcK-ILERJ[Z6<B3/-g3
c/fA&2S1CaWaG/4N?5/5[Pe-X<6O8#g+GW+O)fACX>d@J(g3?.@L3:MH]ERK@W:I
XGdKX=ATE7^2.5&C878VgG@eTP5(DS_8H/Ie@T>E190S2BF[#\Xbdf-\GZ.-5Q=I
d\08:P6e?/]&G#fbL21W7<IOB_NPgPL4AHOeg-JB,aD=^XJ-?G:fTVCPPZ0HQ:D^
a3>abE#Z143dK3bLCF,2-b,-d>_gHXb99@JTZKUd<P><0_;@652\2IKWb3-(5Ne2
8=>34FS-A3^25Q+H^_-7.97<WU\Cb7Y;AcCYXeS.VQVGC3\AP3FbJ76DJM8(=bL9
\0W\;ggeBTL:1M.<:&H30&If5N^?[75KG&LD^=Tg_NE)I-[eaN^d&T?<gg<)DbOO
QNA6)beP4YcbAKdg?\4PI)V[\?a_G783(Ib3\/PI1V\(;])LgT054;E(Rd)1\8KL
/P[Q.:BWL9CBbe(f_6+5;Z;4_J48H7A.XJO/VA&)QDWYg5VbO;5U\)D0d#A1KW6:
/0>Y=2#e,dUXDQ4T0RQ0RH1@3LedQ,b/ZQE_d;+eD2;>K#(OH7RP3Q9E;#Z9P7M=
[RZX/6X&^8=NG?E9b-cI\T?KI@D.V9_8,geCO8=PJXY.B:2,(U=HCP&TJSNYf@D0
.Jb1X97>/QgPSgH=F1J.g4UST;NQG;UW2Tc@M3E7S0]_EP9,W:+A[Eb<KB0IB/&W
G=cT](5&O0QH]K]WUS0F=YbfEJWR^.?5C(QLQ--#OLecZ:4I0@YV(5g-bO8THB3d
HLcfH@J8[1#?(26XT<g0@ST?/(2.?H)(.LdZgEb.ZCH8fEggR^(5;?/#gCC@@6V[
1J4R1U]/]bGe@4dH974=DK5[EW]YZceSR4]TG;MZ#,D>W?+2+;=-J#781\R_,GUU
7A;.-A5GMUZS@\gMXa(T05>/>IYKK);8)0dZ&17P&QbGO<#5OV5,cI9\&&9Gd]gg
4b2/W@b^ebGTD7)dIOIfVg5X(QJ=)aU08_&R@9+KN;a)WXadKG3L-+SgbWH>CHU8
8HIG^ZSUA_bB.P3:L.E#(X,Pa2<K[FbZ<>86Q=O/1KBW9(c_9(-W^bAFH)SdBe?^
eY>>bD(Mg7#;\_e]LI9HaEXP^^g6=[DSW=0H5JT(<VS=D(^TV;5Oe3E]FbM0^KA:
WC4OE6C/UU=]W@f.#S1C43Jg?eR:,H9K9FHa?WV;JZFKFbMF#DD_B;@UE+_@(gc(
>8)e_LO_7NI=4bf9[aJ?2U8X8NN-5;YA#WDeII.SGdAW.2P<4\/3A6G7FS.>P)LP
O&a<C_.GH7E[WN:W:^edA-b3f3[.:I/f@1+UI-83,<OEgZ]_HfL#M9?(aOJ,WJg/
\dJ-(eN9eE@1I46=[\IWDWQW6c)[3Z4<24Md<E?^f^.9TI_F5\7R.S-^_(:DB4U]
&a5]6TBPQ^4]IOWCW-WY590#[>b9E;KH</\/eEVfdC-[S&ND4O0+&M2,@9Q[PN<H
F(\MG&I/VGV,:#(7S<#>SEN]=@OOFQ+;(&<9=4>2R196AW^H]fVRH_QPEO4/E=00
QS]NQ8Rc@8KW6X)e<VYXMAb5,GBGO0+Z180I.8_8;LV)K9:MA=_N0@SDDB:\I9[+
X1>@E,:We7XcR]TL36N.(=UE3\FM(;6@_HZKBN42fHf<VV<,FP29bZN(3I+>2-TH
+Ng^,;&dc#1Z)=bY8?GeV4@=CO[BBRA1;DYGL[^:[Fc?LXBH;41(US+\>dJMYF74
FgD_=dAFW,3DU&4+[=Pd3H:gYQ))\@A-=2X2US?L_RBQF/D1@Z.25B/=69Q_0K>4
aLTOAg&7VVF32X8C+Xf0D<;2[3_7S(?MH7L[FPYeB/6_Fc(G36#JNLHS-0A?#JLK
+\UMJ>+9[bPVYM.+d4-BK_?<7-eZ5QRZ5de:F^feRc9WRN;P>+5[<X+.<N<[C9\=
cT=689HNR:2U;ER(MTD2^c5=IZ2T@LRMJDc)7QIF+K][fQg(B;&,NLd#gaFG(WC2
)4J?&;dIabE\Fc;Z8f;=^>(aLL/XOM36;f#0#J+XWX=LRK2OfY_.QfaB#QZNg24N
L&ba>GYJ-Q[JH2+4M+^,)EMZG_?FZQ<H]\(b41\\APgC.O.e:1/ACg6,VWJEJSPP
O\M_bB8?5B?CHK2;C2K1]ZWF/W(@29a93(-5YB29ZE67,/)<;^)JQO-GV.cG?/,M
]RITbGB?ZNUA/B92^+KR4UHeVY>/=]Y^USED_IHU/.b,](@_JHF?TeSGTN9MQ2KG
PWOV+Q3:=3=YUQKg=[>>?A0c=ZCgDN@NFV2GJeK(EWP4@U?_#]>V/c.P8U#fHgC2
[Y2V1>MZRfT/5Q.:JNddU]04Q]ZWg^@G:QfMVD5MS[fa?d_2\][>MWd+B=_T0+8K
7<ceC.dfYgJP2a904d^:@ZQUU\TB\^:Y&^WbI.UWA1FFU>2)OO.?^)a&Y2/.4;HC
MRDH>+UPeS>=<L:7L9E)O5O?)[GKfeCSFO6d0KbPD0]2_1M=^e-)LL,C7(>6&3RF
P2Y+^2gO31Y:K9#c4C4g<4I,,H(0),:gVZ5)eE[J(&1D:Bf5DCUCe8/W8GJD0g,)
7aACUD1T-5PJ^U:=)<7f+_gT4@]]-ee\(:)ReA&3S\6Q)TMLZA&gWf(/_XP\=&BX
DP6a?)WN+[X9LFBT;91G=E24UHgEJ6\-:Z,OJ(SLJ5KgI=3M24\]:bQ?P<IU0T.6
,Lg?EXMFF_+DN7e,;NWcG?HUJX\1He[++4LOU1DE<=X];f@WVfG6Y,>,=]>d:.6Y
>c\G29_YM@2L/VHf95UO0E2=<:\aZ/N<S/dZ(PdQ_^BB8@3^U@K0W7b)e;#^GFKc
+O@#N6O.,3WO=QLX[^N4KcXAP#:LdVCGX&C82ZLH3dO8WC3B?2/QM)c-JM)LFQ66
gF>-S:WV#e0#b75JB>R7?/Z19<Z?@)C6<J\McX90(a0W:OJ+)Og:Db2]/9:#(^7a
UD),K522GEff4SV2NGABY8BcfM>4]f3C)7;PPa_6W\.Y:.=A<E8MS+:a+0560B&T
2[ZV/F_;LN[&LHRa#1,>ICZ51H(4.]9GLMK:_)H8a#3R1N2D7:7I/#-E^HG(:K;:
H1[U,I=b?.Tf98AB-c<&DA/NJNIRGfad89NQa3<,1Vg;F@W_&7K9M7P6NXZdb#+R
9#\-]D^#gBb\F&S7/?X&9[d79GA(&II^1dIba_2H6Y2D.6Y08\^GEE4a/_T@<PP0
:7Q11&[?52Na&(3S8C&I4PBKKU2a>=_3D[9JfE3;L.PW+@=<ET8S8PEJXZae^-gg
&3=8<#T..dI#O3\&DBVGL@,=dcN^^.OTFP8EXUR=J[W&Zf\YN>E:2KaHNf:A3^L.
D]2UgYE=RSCPDHCKQI##86UZ#+ddI&,[\YHF7J\YbfOZ8\b6NVRAX35/9V&OCSAa
R^US60M]59]L[^P@PJ2=/PL4;QCE69<O<IB-aTJ(O3-Y+&QAR:c<XOYF)6Y/Vc75
?D_FFCTK9>59&Y:)M@FZfe[4[-H&R(Ta^Gc+S-8DR(8NLQBBYK06K6b4)1)aRXVO
T_H(.F#EIK[::.MG?;KMWEULWS&L=(]L0Db2:ZZ<P4@^5C<GBSa8/(JU3M@:)f8=
_cS2=bb;B<I+E]/4G3^Fg(Z^C:d6[3Zb@E5X,VE_=;d^ScYP0QHB=g?.?.5[?PH9
]72TH_H-:D4cR\,O0^gAeZL<@YgC;-L:^JBU\]W2(T#-0bH+T>#J\MP/b:1W+Y[P
0f.K5PR]4=.X7AgOYM,&IW+.H:R(ScTeZA:FOOL,LcGaX<G>129BHcED^1d^)gIb
M+^C&fF,<Z7+@HD_Q71^eVS.\@&T1A0]g\IA#:=B-Z)_KSG](ILPTY7QW9:ORb-/
IP/#4/D6?J+.JN+a5a-.1_fg5b:JOCR6Vc<IMHTBR:PZNL[?b&OYaO.ef&A10JKB
^^9_O#(?=aPN&)#_VF@1(e=[JMQDb][1;^4;+Lf+f#e.?R.DK]<62df7.e\#/aTN
W?_4f5S+.@6G/(LNg-W,?[2TPS;4#8ZE<Z]_DCK@+d,;JGbFCZ<2Ne+@JWJ,07TT
P0VKZ2L/I64<EQW=+@2<_?5?85^RT/IQa=DWb]5L-bK/Pc,4TY+[0D2&?[8(Q@cQ
R].U1Xc_LC.eU5272g;.)#+I9M;:IIdeU-A+]dXbVA0_:c8WBC3/PDG_9_e[3<EP
[.,9eCEB@_.He,[7T#5GEJfX@]@:X]ZZ><BMP-3)IX>E6J^[gJ-<3[+gc(OH?P6M
J_U_gQY]UdPBb]6c8JT.89H+5M<N[B)Z-X?\Je.3bK1?@faQETK:,g+Z,=f&;:[\
a>JNfSg>298H<<IF,>c(JS&JWc+^=H2ce45P2aFJ,]I=Re)SW5\dKeC7dO=e;+GI
(N+Y^D#X>\ONLe2.TF7fYC3LX&D)M#d7g@.<H6T18J&VLbJTWeIJ9NIWR>FBUR)2
RM)B.?9D78FLa;@UfT?^UF4ZV7&f-5AK>+<LSOH_TQM\JUZd<gNI[LMa8MZc76H\
C]NaCd@@VbO>F.G:S3@SB&E+RgKB:RQ,.Mf-^UDUWNE\FB:S.J08E6;5U?SaZJ+M
:56VQ:cdg?>eB6O6=4c#D[=T;S?;d8T-a<2R89LG/)AdCPQQSDJDLC.NU[M1/\^[
+>g00]T_#P(Ka?d\4fD-G?BLCE93KPVe:OIT,I:57(I<.cAfKY\+C^TK4HeO?gG;
HL(MHE?5^_S4)dIMA9G>8J3Q>f6PcM9Y+FA]gQaaV?e3A,9?QU@LSA#[g]:SN8:5
(/ag-?7JT((c&f9N];,c?_>)0b#Q&,I2_g2c?-@IKC3LA\88OZaNV8CNIfQ;@.7B
1^O0,.H2ADb]NBbYD@IF#^#Mf\Ie2,K-JSbLU>K9@H9M:gE)fXX/VD3W7(a76L.5
:G3HLF-.Y\)>_]RdPJFOcS_Y4SC:@0eCU6\\M&K,?2]<M;^8:@>9,3?ac3NNVFY2
O#7W<F.dL@I@Da:I,[^bMKB/&bdCaPA=_F>)PQVXF5\;V8gH[;16agNYJ6\;I(A?
#c?b^[7@V:f&AHdQ7EQ@B]102/+&f-\O\)Y#[Y&GO(]2<>)OE_d+QCW9c]4S0fFa
(Oa@H3df]I)OUE;G&]BWL7H9AZP,^-.3WYW->.MfS>P7R+FaaJT@?>,G5FcS6?P&
T7SD]E\fQ:/&a;:^7]L9,7QB.e::)F,UF;YWPE<N]NFO,>YS7,^HJ)B/D\P[YAWc
1d?FZ6^RFO1A/6;8[)KL-\T@WC8CbW^\TV6Kg\ZG5<J&Rf,YEMA/f()7I2:d3#N^
D<^Pc0MVFJb.#H>;JSR>MdFEP([ADe,C&:PLKcJbX0U)TL@FD<]/Z4ObH/\+PR70
>d6W,-_]9KT_@,/YL/4P,^-L^ZL#GdSI(MX>_J@b#BF7H)SFRUWU8[@UI^UTc/PP
7M3a-FV)N9GJgIAfQ4Q(TT[+MPMGBKUO7N;\76K;QAMA(NJS+:AA.5(KKgd<TVTE
/?a#J@O=cYbETagUR7JDU[>5&0Y(2Q@N)e1)=JcX#d>SA:@S\c+Xd\-dRR@e[;1D
a(CeU23H;.ZPYN2G3Vdg,e541G@^+:SegZ>B\ETO:g=R2I/X)/4K)fJ>f46F^;b8
Y_d1Y_Q;&)E#)XK\DKaQ^<WM>A#^cG,H?,d5/FUQ/OF@Bg?c,E+0g5@\Q>bUC#86
^bM:_8\FWX/e(9L=EUg0>ScR(#IaS2FH6_[3;FPe]IY,Z,/\;5Sg]g<H&ZO1<Pg:
3DY&#6I4XS33XN/UJ(&?/M/FAc&;e8Uf,g:RdeI#N&RFKBWO#)DeIX^f8(-IP.gS
EbcY,^X.@I6acN_3RD5L,bE?D.JS#&.Mf3WX<BgR1&e+YUQYO+N4WL]GNMLCB1X[
dCVQ^Ga=V4ZK>D>bLF=-E-B;?>P:\GN8UQH7VTW=2>.,4_Vd-XNIT/XF^B\=fVQF
==0aV;&[g<2c>,4bO7>S-3NRN6e?4?.#3;-KgD=HeW5J7eSegDT5cZO=6gW5H&cO
#N\@P^TU#.=K8L\N3E@IF^ggH+2,WP9W:YR<bG3<PLfd(K<c59.=f;/.6fVSHKRK
921.)EE5F5.88E\K]D_=PSaHccM_8BWE#<c;,b,#0?MaG&16J7K<:;6J::0X6XPX
#;./,&3G]FHde:)EO&e;M#O-fZDZLa,/GS_R(L@Z#YL4W6c<?:A[3b1UY=FRR3U0
&;A?)fGCfe:Bg-P2d2aeUA-)Ig/d+ZK<\-L>?A,;?KccC?a4<W8[Dd-PaVM:LCH-
6d,3OHKVQM#b28Q.8I]d/ASN=+6?7/gW?YZQ&&]C(E(1XZ])KbWZ/-3>6JX_+\g_
\SB\<ZTKSVdB=bVf51KcE>])Lc7X([XKKC6HOR,?CISWRX+AW=ATfN3fL/)2K)?a
&RT>c8UGe<DVQQX-@2#ID6)&bIP\R\\3Z<?BaH69LBS.8&8K.CW@ZWP\:F,AO1C#
ZRbGYH&9@MfSXQX/gCPL3^KRTJ6VcS1)&D^L-RaA=KL_26N&Y+GaYZU2a]e,2^IC
f>_;R^]VUF-W+/f9AB323I+/\\2/f?8X0=:)-74-a4(.)9eCXL[^IYg3[\H2UZ1<
PP/7dS1dV./a47YZOc3>-e(I1A2\K,V_QHU9K>JYGd&(C?b=H(R>T^+)W,YX9PL9
S@A\I@+@EHW\OgAC..4YCTgBWbR0A\@7&9(^,6)N;WaQ(:YO>bS)T3593V(^IKDC
&A]42,_F91JW=>=BORb;cfF/:4Cb+D+-YJ?M?QR@FKQ7:Ya_OGOQD,J65\O<+:<;
cA5H.DDPX/5,]M_NS)7bEO<(cgV3M/AccD6VX(68M#9OX/[[\.1Q(864._VBX\@N
W8^C2J615f1E6Xf?RBEfP=W70Df\)<2a\IPT^R7FSKV;W^N^e26K.9XVdI@R\MKE
W;LN0@fFIG2_XWB:M5#4JWQVVF]0)^;Be;5NY7-@TX\5f71,--Y6e]c-aO#DM]5L
+V)&?e\:<#Y4GD\FF;F+T^E<MgTWd:7I;^b12=+OI.9P0(CU7B>7M;G(^/NJHL<0
c3X&cAXM/b2X2GO+/:KM3)X2/(Y<1^,.A?UdMY2;3P/-&LZFAU5Wgc]TRVE)EVN;
?D&4B8/:Q2O6[6_ZbaS\QQe_E7:-SYX]&XO+6,X;_RPQfF9?G^I+39U_:aB+_K=]
:[SXd)ULbGI&N-Xe,;aQZRg>M0D>(a>ZWRcJ(_-EY1+]F[DDSfJg@9S+X5L-[BRK
,^B:X)g#P3;C=+DBJ05#N2TILAU,=SRfKb&ReMg-8bK^H/JA58DZR=cV@0_-VcDa
<D)[]?=4/YC6#d0[];C(4K(12+2I_7A9]?[;&#&C?#K@f6W.5T>,L37L\(3]<#DR
BJ]#C?G-MUBL\P&)YE#_,5?g2-\3HF#eO>4W+.GVTPII3=MN3UHBPcL/>aJYC@(-
:LP01&PJge^-;ac_AA.R&]>72AQLC_7]agT,<5K_<<Vd63P<f_BE8g/?<JVe0b5#
7EE_=gY=f?0FE(9^<cfd][LY3C:>dN59SH=gf<>F;7Oa2]2#LX3Rd5WFA\[FV4PC
[^9Q4<g.a+W&R3K,=V(#I+:-?W2XI[KM&S7e]/fV4P-BTVY?ZCYCbOU9L/#bXDRB
NPYdS.V\,T1=4VUd2Bc9S#R.Ga?g;#X._SGT(_GTVHf?VP</KBQ:184YLT&a76\,
8Q_P@E5ZY=^K1TVK\HMMI/:ETSF4ba;M&#.>Z#P04D?_6ZcS+)B3=fLEMbB=H))K
G2<U#bP7(1Qc#2Q4^1[Y<J&#6Sd)13/K:.U]5XXV;&+-+C>5gKEd5.+d\Z]TI]@6
S_;IL=JO3=GJe9I99R40W<=3BT@NdS3PXCb.KVVIEW32?/:3-eE;>0e=,XIWSaJ+
LYX;8R<.I-E]BO)QM]2E+&+KF[d0<:<?/K=2<(>dg<3U]GDAPW&K)XX_7G)8.D>G
>Eg47f<bV^;,LVJANKB>-/LS_8]&-72dON^.G1PC)DEOR6L+=cT;@Nb<C?.HJ03@
)&,P;E[BIG>C=b,;H,O1FG./A[>K.3\;^,#OH?RFeeNVd=Hde#Qe_T.A&&7#3I61
:YV2=&WO[:SS)=5+-E52@0OQL><AAVdHSE@g<@FPfPAY/-WI/+^WaUU8-bb4W=9&
P6WW+A/B2/Mc?.Y[)Ece&@d4aaYN/_)Q&ZgcUW_e,(ZYL>AN99aE5/;LTL:9^]18
C6I82eA:JJ?>CEf8K8.C8]:fOY+\+]GNM7-A1.8D36FfS,+I;X<3cM(=I_f]EP]J
5RS?<4;U4MA>35].U<=E]#8[X#F=@9MQ0NNI[>M;3[Z&(ge2-ECRgRBA[R&#ddYB
/\=,HY8O@-CR,bJ09Q^b#CVQUbDW3(ec:CEP1/U4+e)85I&@a>(R^/)>=O993ADO
XL4W0&=?G,XGQOB6&1Vc@XcQ_9@,eFB[ebWN+XBf4QVEZXKS85&KFWP6KT4P=H#@
0ARf&;?KNG7<_F\f.@S]0U-F,)=]+=?DW,JY5W-e9@7dfcB@E@=ZdRI2F=)^+IA?
cY>:?[NZ/^d>,I]b[9=W?OC;J-D>VA8/YSgUNa=NZc+Q1.G7^PT42SPbH9M5>MWd
GL<2M)S?OY,NT_]4:cM0TBdg+6-(9^-WBHM))G.RG.Z9-X_b^C3-eYbf_0BJ-DY8
VaC5HN^3bITYQ@Ya[_K)ccUTA2ING.L13KMX>DDdH).UB<KbV]->d;g:BD5PPLH3
,^)g&HMf007KAfbQ-&79VM2J38@<^?DATETE(LD6/3&d4ZS^;Y>B/K]/GH0-CK0X
=SBZ7@G;[NZg\c>\]RMPJ)N)8[S>6=+Y8.:WUbFfDO;aRLd/\AYcUF+b)2UX^3&b
[_19(Z<#ec9TXRC>gB?.(_#Z_fO=#d&^KKZPV+I&T,?4eR]X,;N6Lc5]P]P;W+=X
CVEVHP>:5JVM4UGdYgaU:+0d<Q+)_W65SG7K=cD&IOeTVRO?)aB=BO:ITbb+L2Z1
QQ)UBMIGKc:TEM\8<,.(33@#3HK+Z(bb+/N(5UP7;&8M7aOG04g0.&>Oe2_HK5Sa
_L=GB4_.J?XJ&N6<H.T?7D#,d?59>?,d0N5Pf^d//9TSE)1,H=609#6@906(V,;C
)6)PY,4Idf[ZfUC-A<CXDPfFee7&_UAZGI0E#<+T0?R60W_,@EbIAP7O7O+B6a_\
UcWXLe)<aTO\O<W&9d\dVYPg&C<0)36OU0c(>;9?S=JPZSF[#c6N6K-7VCUUDb8(
^W0g>DJN#[,9OZMM.,@C)Q-42B4G?e7H#^<_T,V_Yfgg\[\:@7@5:Q][.;(FU/6M
9N9XFM0-Ed-dWG)^@b3[QNV.EVeQ2X;8cIcSR^eE^_/^(A#.?)M,-.WF&)_-[+L&
f]CWENWGO]Z5&DV4Q]8TS]Z-\0,6<f\VTJZ3G&TVA+173B1=7U16@[9CV4]g>#U#
6RXW&+7OZPg#&U+Ea.CLVJUA\Z0^eaC<T3e3f>UPID(Z@/\dX(RdXYQd5[63.fbd
UFO9\51dM3FD&BT2WU#O_J.[T7?C-FCC3@<,NNLCff=VH6N4ccL]1B(,CEGY6.4.
X_QEfbg[@]5X0QV7D@5NT>)O/#Og4?bXMVR^?D7;O+DT;Z((/;)R=&LF=(^[F^a=
7X0EF<Efa..Ud/OG]0+g0J2>1KPUJ/GJGUN\59BAH31S^KQA@4eYf1.DaLd=ZD,^
,,A]=22@-,6/4S)S6D@Oc>fWZ22:A::98QY:ZcGc5(_J\?g=B@QP[.,Vc4FP?VB.
\9-NMUUGXO_VTfD_L#D=;VD.=)_&AQYb9Q(,3HPeg156CE?CF@aa:0@Ae,07N/&]
XSJ>R061Ae0)E43(eMPY<QUPZ4_,0JWWO3<eDBAY-[BJE2S_+CD10/37SEMCG(#U
)7OP-AIJ9b-2HWeIa@<f-L@RC4C1LRcR_ROAJeHFe<7.DJ@gFQKEF/a>W+aIX,(.
0=HL9TI3HA]WEH@48YNPSDQgbNG[1FbOJ?a_D;_@Tf^Y_Z.g89&RFPS7S)YPad(:
3QU#g-3TGDBHb9WK1Kf=NB-1+4S),;.7cb7)QWGW=SVP[ebMgVUYV#>KKP.gMd&\
9\)+54H4dF)aHA5PVCET,LCI]fbM[\O#E?IYC<L>9.HF,?Hc=V5B6[P>+:gSM=eG
f.G6._eU)Bgc?:++F(T1O2+].B+()3(Y[LOV<[Z3)^e);KbLae9,E69LOQebELUS
bA;HSH0Jg3W3^/)J^/BX2P^0=V6:?2--9$
`endprotected

`endif
