
`ifndef GUARD_SVT_AXI_MASTER_TRANSACTION_SV
`define GUARD_SVT_AXI_MASTER_TRANSACTION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_port_configuration;

/**
    The master transaction class extends from the AXI transaction base class
    svt_axi_transaction. The master transaction class contains the constraints
    for master specific members in the base transaction class. At the end of
    each transaction, the master VIP component provides object of type
    svt_axi_master_transaction from its analysis ports, in active and passive
    mode.
 */
class svt_axi_master_transaction extends svt_axi_transaction; 

 /** @cond PRIVATE */

/** @endcond */

  `ifdef SVT_AXI_QVN_ENABLE

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use for each token request.
   * Each entry of this array will be used as QOS value for token requests made in chronological order
   * for first token request it will use qvn_qos_value_queue[0], for second request qvn_qos_value_queue[1]
   * and so on. Each QOS value is bounded within [0:\`SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   * NOTE: size of "qvn_qos_value_queue[]" array size is set to "(qvn_num_addr_token_request+1)" so that,
   * at least one QOS value is available when transaction is not configured to request any token and master
   * driver has to make a token request.
   */
  rand int qvn_qos_value_queue[];

  /**
   * @groupname qvn_parameters
   * QVN allows a master to change QOS value it has driven on the bus, while it is waiting for grant
   * from slave after requesting a token to send a transaction to an AXI channel. However, this change
   * has to be in an increasing order i.e. changed value should be higher than previous value.
   *
   * "qvn_num_qos_upgrade" specifies maximum how many QOS value upgrade master will perform while waiting
   * for a token request grant for sufficiently long time. This means, if master requests a token and it 
   * is granted soon then there may not be any QOS upgrade. If it is granted with some delay, then master
   * may perform few QOS upgrade. If token request is not granted for a very long time then master may
   * perform maximum number of QOS upgrade specified by "qvn_num_qos_upgrade". Once these many QOS upgrade
   * is made then onwards it will not change QOS value at all, even if token request is still waiting for
   * grant from its associated slave.
   *
   * SVT_AXI_MAX_QVN_NUM_QOS_UPGRADE can be used to customize usable QOS values. Default: [4'h0 : 4'hF]
   *
   */
  rand int qvn_num_qos_upgrade = 1;

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use to upgrade any value it has driven on QOS signal for
   * first token request. To clarify, when master sends first token request for current transaction,
   * it will drive QOS signal with qvn_qos_value_queue[0] value. If number of QOS upgrade specified in 
   * "qvn_num_qos_upgrade" is greater than 0 then it checks how long it has waited for token request grant.
   * If it waited for at least corresponding qos_upgrade_delay then master will upgrade its QOS value, 
   * already driven on the bus, to the first entry of qvn_qos_upgrade_value_queue[0]. 
   * If it so happens that master is still waiting for token request grant and it reaches next QOS upgrade
   * delay specified, then at that time it will use next entry i.e. qvn_qos_upgrade_value_queue[1] to upgrade
   * QOS again and this process will repeat until token request is granted by slave or number of QOS upgrade
   * is reached to qvn_num_qos_upgrade value, whichever is earlier.
   *
   * NOTE: Master doesn't support upgrading QOS for tokens requested in advance i.e. it upgrades QOS only
   * for first token request made for each transaction it sends to read or write address channel.
   * Each QOS value is bounded within [0:SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   */
  rand int qvn_qos_upgrade_value_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how long a master should wait after sending a token request, before it can upgrade QOS value.
   * Example: When master sends token request, it will drive QOS signals with qvn_qos_value_queue[0] value.
   * If number of QOS upgrade specified in "qvn_num_qos_upgrade" is greater than 0 and it already waited for
   * number of clock cycles (i/f clock) specified in "qvn_qos_upgrade_delay_queue[0]" then in next clock cycle
   * master will upgrade QOS value taken from "qvn_qos_upgrade_value_queue[0]".
   * Similarly, if master is still waiting for token request to be granted by slave then it will use next
   * entry in "qvn_qos_upgrade_delay_queue[]" to decide when to perform next QOS upgrade and it will repeat 
   * the process until it has upgraded QOS for maximum number of times as specified in "qvn_num_qos_upgrade"
   * or token request is granted by slave, whichever is earlier.
   *
   * NOTE: size of "qvn_qos_upgrade_delay_queue[]" array should be equal to "qvn_num_qos_upgrade". 
   *       each "qvn_qos_upgrade_delay_queue[]" array entry value should be a non-zero positive number
   * SVT_AXI_MAX_QVN_QOS_UPGRADE_DELAY_RANGE allows these delay values to be easily customized.
   * Default: maximum allowed delay range is set as [2:32] clock cycles
   */
  rand int qvn_qos_upgrade_delay_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how many address channel tokens driver will request while sending this current transaction
   * to appropriate read or write axi channel. Even though QVN protocol requires one token to be requested
   * to send one transaction on address channel, Master can however create a transaction (xact) with more
   * tokens to be requested, in order to pipeline token request and reduce overhead of token grant delay.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       address token as transaction dependency i.e. if no token is available then it starts sending
   *       current transaction as soon as 1 token is granted while requesting rest of the specified tokens
   *       in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_ADDR_TOKEN_REQUEST define.
   * Default value is set to 16
   *
   */
  rand int qvn_num_addr_token_request = 1;

  /**
   * @groupname qvn_parameters
   * Specifies how many data channel tokens driver will request while sending write data of current transaction.
   * QVN protocol requires one token to be requested to send one beat of data on write data channel, so Master 
   * should set its value at least equal to burst_length. However more tokens can also be requested, in order to
   * pipeline token request and reduce overhead of token grant delay for furture transactions.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       data token for payload dependency i.e. if no token is available then it starts transferring
   *       one data-beat as soon as 1 token is granted while requesting rest of the specified tokens in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_DATA_TOKEN_REQUEST define.
   * Default value is set to 544
   *
   */
  rand int qvn_num_data_token_request = 1;

  `endif


  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_typename(svt_axi_master_transaction)
  `endif

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Random Index that chooses which particular start and end address entry from nonshareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned nonshareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from innershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned innershareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from outershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned outershareable_addr_range_index ;

  /** Indicates which domain-address-range has been used to randomize or assign address for this transaction.
    * [0] => '1' represents address belongs to INNERSHAREABLE domain
    * [1] => '1' represents address belongs to OUTERSHAREABLE domain
    * [2] => '1' represents address belongs to NONSHAREABLE domain
    */
  local bit [2:0] addr_based_domain_mode = 0;

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_master_transaction", "class" );
  `endif

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

  // **************************************************************************
  //       Valid Ranges Constraints
  // **************************************************************************

  /*
    Mainly covers the valid ranges with signals are not enabled for AXI4. Covers
    the state of options signals during AXI4 Lite
  */
`protected
+g+[F?aaN19Ja?Kf4<30G[1a5Da)&f9/)>SV3I-fV-/U^A/.V.EU-)KE\9_QgAQY
5f_?[OBLFa8J,$
`endprotected

//vcs_vip_protect
`protected
VKg9a<]fRM=ML0aSN.e@\I>9(L0EGFBfQcT][L-F=>5;gT[,@3X]+(2^348[ULX1
>>[;PU5=JCEF==JUAM,RJ=@+19B?NZUBHGEM;MQWL38LS<g3IWX>^=W<=G@g0bba
.&,#0__8-?Df&8U,#T[.aHcD(4-f2OCTX+Q,VZ_E^AR/YPf4B\b4&K19@#.-ZMO_
<8,<9HYRM+)^O0.,P^OgUUBJfS-6A<]0TYKX,#\cN&fA.E]9,0gbY-d].C7S]?<^
,#,FWg2GG^8,EG5MWFZU_cG7K(ZK04ENJD<MgeK&0B7+[--ZWG92e8=1.HJ5^Q,D
P9>I6MWN>RXRJ)W2(/fZ-UD=D[ANW9D4C-A2JM2^=;;;<G0RURY/b_D7\FH;9RO?
4&fVX3YT7Lb[^,T,-G]>F<(a:D1&53[>fENcbQ_aS\cW\20G5H/D@-=d84WUg2C4
P_d0M5\_VUXJB=6DPDS4#VH8);O\_5K9>/8O6Z61A4JLYS_a;@&+0;+Z8aFZE#2?
3bF^T[T</OZR8^;M8&ASJZH/@Oc5,eE>7/@UMPI3;,NLY:7L4\B.#3AdWEQ^,A9&
&AQ^]<V4bH5QMGPI5b,.WgL#@6eVMKV0N0eQ0D+KN(D;5@@e\F(RF3aV-A_#+^<5
b>I]QBeE1[V0X69.FQMgR(g=ZC7XE>gW&H&92;4a/PAT0_1.J5/</=_d:/Q(;ZVS
I[_9/8+67&RNR_8\26M7Vf1[B=eUT7WV1,QL>\6IRSC<31X_)9WdWY4@cD,)#0/L
4O&A/B(UTW#c:J/Uf,4aY)8^,2ZQ<U[4]N3]d]B]L(^._[0(CHeAQ)/_c94&U=C@
QRbIOIXZ=ZNIHP(K(.+G^;=b\23D[,a+NOBQ&C?H7\J?1#=[,]W.;I=OT[^ES+aS
D)T?RVO64Z0C@BIUF<fI=]aI8_F+NT@f50&gZ;b:XfXKWg\4@Y2N6J-gYUfFAYeG
V@VT&+RY)83:.TKXR-TIKP[=G2+,/P0R4>>RD-/,2gU,J#IUYA07WE(&B4=F-@G[
F/XYY0Q6d;;88,\JTc3@NcP&+/M(IZ[^ETPCS<4HAeDgF[LPT+@39B:@^_OYKL5N
WRMPe\84SZWK8T#N_,9OgZ?JQDS8TEQ17GPd^]d(FHUYG^,]Xc<VcR]A)84:T>P+
aL0_BO^UGeb>KR+UH29bV>6W>A8.N(/>e\7XCTgKCR\BEK740eHXG&d6MWeG<=&e
3,P@D>#79g)3gN2;\3U+4VS]]]@a:42f)X\14DY:U2f,YH,V&P.6a3;OTPeDX?;.
ZC_]K[cH+gJ@O9NR5[X(MJ[18DOT@MM\8B&YH=<d_N2I1OPA?=M@VQ0/T#JNeU7_
?X6N#PGL]\>\#XaW_Ufge#BY8;Sg4K=9>?P8IdHC_^?KP8B9TXM89YDYZK^-1:82
IMN8F3J6(?cUMQV#;01\32M,\2,MCASEAUe;4RL]W.#XS=A9]8U/:D(fO#P]I=UN
ZDd=[e>Y4b[DZ2=g(_6[@AQXV?@<Z3ZXMG&0:,.[A[PIQIIdg9DTCP20THQTB]8^
522B0g\XGKJ7VO;1;AG(#M-Fa3?31VN(cMg:e-N9VFRXW#\f\6T/;I_NfK-B>Bd6
F6939Ig1X[Z\^]GYBR=UXM:U1+dP]J_P&^\?FH)V&7beIY7d=c_T]C2U.Y./<AXb
)7J4#-gO28WW[YW]XO)EM^UJ[2+WbF.a,:<dJfUGDC)8/DY4E29_C).V&]a>6/MK
JV@[@=-:_R612E)0_WEFLVQE6Z04O[_cUeD4JX6b)fPSO7@feQ[cA:eFG<IT^OY4
QKWND2e[,M3+9RQ@)M9dJVEVS(?dCF7#bgaVa#6&&L1aY205&/\UE[EF4Gg[R=&K
[#fQ2PKg,-(Nb;Q?9E63\&65;:@0HJM?];Z1]5,I/Z0;+fQ+51S=ZXEQLYa1CJ(G
U8#Y=:8<Gf]](bV^G5/I4N5J4(M@#1+G?bKL^^4cXf00MDOQA(E,HU&::^?\<EW#
W#M=<UDYFCLO9@</P/0\dV,D[@\V3UYb-<(2=/OL4EM]XVD:EE,+P0GJEGO4g:I7
T8F^64aGU>bb^2e(O8&-1g1ELP20EMB68]VPUX_Ec:b->T4@RfB-6JD=5gX:@R[c
=0RdCKK(]/4T\IB+[fBa63S?PW6H8db7ZNR:gZe#6DBDMbHF]7R<)1&29]YeSHKV
[[DL19W=]\A_3QPeY&QXBUM+#0Y/,QV(e=78&HUFHW9;ebQ;6H^1[],;ABGe>X^U
8VJ9188Q?.\-;&7&-Vbe[<I;PB[F<\F:.B7FdG7YY_YFAO?8#NMadf=)/WT;15_H
WI)Ia>ZM)=PP.>Q-3:6)#CMQKDDI5OY#bN1S((eaL]_RO+H]W-0+@,0_\[JEa&gH
7?JUc__?,+GO#@4U3cLHWPZQK:)-@fSY6QNPdaa+<NDVa>B)e^e3IeO\\Hbgf4>4
39^#2MM,bc-IYg9QOZ]^^U#-8-?KgK^.g_<&L8F@Y3=Q-#7U7d6-R4EEFCD5HZS_
&H/S</[HgTc,GS4@8>1HaODfbHRfWZS-8XdU5@S8K4G:,^=;T38@]U])P/.MR]8C
3]Z0V4g;_&HXM#H+[.NI-Xe,W8\#T#IMKA.C\_58(NY+Af3QP7a++&fe1FD:(;#-
@QFdC9De[2M.LK&6K_ZMRg2]+\D<E(;N.T#g1GbQ5^PfZOeJ_0MNc?4:Tg6,L_<6
e3G65.J((,&Y2-^CVHD?-I(MXFR?(8_[@WKR^RKc<Tdf-3RD^ZTZP(cK6JIKUF31
CV\bg)dCEE>M=e<<c0Z#-g)23]@VXK?INR92K#+:CgAH8TF:;Da(NFH5))Ve&aC7
g7HU8V)8cP?0UUS,CE(IcHY;)-)b_V#&T6+NXYC4O?0QC2N/D+XD5]6.T97U<2@X
)W>MMB\g1.-B9\L(&9b57g/D,5D.fa8X<U8,2Wd\ZOcHM,a]g;(+MM3dV:?M^X@S
?XD1BVO9;f0<CL8P^C]_X_59[;f07X92V)Y^CT]8eS98-5f+Vd#_eI4Ab?KD@)e7
S=W@FHdPB,Y2fcP2M)LD\^ZP;2-0.R1c^+7B\APb:0W8-?T7T6,1G.P67a929;[O
77OPJf7V8O[;E;WdKWU^-f??H_N6H094;UDf=\]9OZJ/M+&3\U4,U(VA55G[QHOg
(L7H&1:V54FXed74;@\?-&ZEEW48gaK=G\Ng2?+f;OZ&T[^H:#TeJ:bVQGY#5.?]
KZ4d^C1=6;f5d0X/=Lb<AI(BS50B[_+B:)7#f0?fc=N><ECQXY3?,)g3(JGgR7BQ
E5eCB:B2?cOdU^(8dKU/D@d0?F=g^K;=[LIdOFa.PbZ+OP(+G#:[0d);F232_A\9
A^,WH3]6?85^e4Z9B^5,SJI^7R16&M\69^_S;?TDLIfg5R0R>TGLF9TbH#Q3HM>N
];BYVe5WH.>(ae/[ad0IfgI2D=>a4MOK1P4++NK^EIe1aMO,M6QKEE8RaN&<YDO-
NRdG>7?#3^N8S/E>1/TRb,X3>FUcS>437_JKXQ7,DONM]VE+49]]9g\?g@/,8N8;
1Q2Ca<OQ7]^JPI+DQ^IZ>(Q-?6IZ\Mc&ANS#PD)aMQ=@@NfeFWIb3H.6S4RL^<\3
W4));;I(g&^[>:N=@TE+IA>Kd]3a@(e=7fBA69N7..)4e;)_NXd)SXKW5(72P8&N
7=G)@^A;M>NPe8](#]+-_T53J49BYN7PN:IEP0-)^W8N6/E54)L5.L4==^b>E/b?
4[9HZMI?C^>A#bY92OY4AK,8BKP\WS].J:;B/\\Z>K33H.,&Z@Q16_OH07-U\f?0
..cG_Ed/816GWa/I-Pc+UWD+=-?,9g+=L;0L,MR#cK&/4=Sd=;KH2[MeLLYUV.##
gIBT5?91JBL;WJM;E3@IW/f&-H0g_S<^fK-I87Le)ZB.G^^YO35C/Vb^Sg0>C(De
2CK8CJ+A]a3O:gVX13&7?6+CC(IN@MWRN39QdJJf=ed7:8[J.0/GePC)3=N]3)a[
8RL7,f23DOY;_QVA7b@D1T^6/fJ9/:V_5F9V20DaW3U:U93C<(K-R/[[S]/V+R.;
[RA];&VEA+.gW.7K]5G7ND/gC=QGVD&O+cI:VP6&>>DDK0DTW4J0G1/-SC<(O8N(
@G-9###\GFQ_Y<KC#<],]U7dP#14R3^gM-,10=g9?R#e<gYQ;6GJ4/[M9JJXM>M3
dFWdEJZ@?=(Mb/4Cag?KLc2Q8DN1[J+N[;=7d135D6;T1VL1GEAWd+M@#ZY\STWK
32aV8T6S[MLTB)b+FY2ZIZ\H[/3YVC)RUgYOSS\RW;A_CQ6WX_[0L6>b6B.02@W_
1QfAb,.B;M0dQcN9Zde;?&F:RIfHf-RfI@>FJ)H\R[MeF&,=YS]QeSBP2;ZLS&@1
AVD<?9C_[_<K5.(BXE.3WO-DZ@(eQMI;Ff7]a5:J5f^[@,S05ZWI#VE?4eYM;4PH
_MJ#KO4H(YPfZ[gD(L467F?;FK2\.eL[>I=LgDNL1D.JaDG#GcgbO=a5<C)KdL#9
H-fR@I[=b5R4<e0DNN&73b/gU1+0U_&>Bd-^K#+>_HW7K:?3?-M6=GN\G?e@LK#D
U/EXV7]94(d?2YP&\C(S04&?bH92\E/C_3(@F?S8WZ4Xf&/T,>dUb.KP<bEb5a3_
H[Vd??&Ad<2Q1TRe\>I1-NK0WSb-gcPD9^A@\JGDS)MLf,V+N)EZQXN>Xb@G\+OJ
;M@.bH<;cV^NXV,/3c]Gb]RUGO9XAJf)9#+HGH:UE79UVfJg>^d2cQCQC1N72f@]
f=CF9[P0,U9GTHRDXO1\U@/E_:QZ_L3Qb:&YU&7g3-P<RK9MWd(7KMO.SJ7.3G]b
(]aYe^V6W\LQXT@\34,S60Q2ADAf_#(UR(8aCFgNGCa6YF7&5SBX.T]A5ZZd^0K+
UR23+Uadc2d_cfC<XY5?P5+A>e120.T:W.\]+&K?[_gF)N#@9)0/HJ(e#)fHNXY9
DJMHXO+)Jaa4M.D4YD_VH\V>QdfHS<\VbTZc_O3O:9+M-YI/GG.0a^bb=>+U#<\:
gKZF=7O)H,W23bLM#ZS)(36W]Xa:ZX[>LJ4TM#)Z/DddJGH/1R1AFQP(TDBH?(Z9
)WbFbF9W,?bcWOGU]f.OXNYJfX3&6>&(RD?A3ecYP#b;&gc?#2W1P?RcR9Y29;Ra
DG:\[9eE9g(RYO,TAd]_^#SIdP4[B^e.YNUFcFH9>f+DCGEC4X=:g@<f</T<?V8,
RgPMQaU091+-RaQBCXE7.)1YZLf^gZOZZd4U>P0R7KI7-d19LAF160+?)\IOCB/E
5eV0S_b;3S+-5CG#E=\]\_eO.6?_b@7HTQP(8]8J@0^21T7KBae,P<;e@?UL,HDQ
S0[FLIN\SY5gAX)e/03M+GM+=.9;CQAIF&&ENSf-X2KK?Jc8#)V&\G5[U1f6;-T]
=C).@HcS84JA?Yc)(fXa9-;;b=gf#:LI&Qf3J/0XG6-LIgf:)#7@MQ7>)@FbI/-/
T/RGC:E?:RYYNegF[bDW6VCN:W:.RXTA(C>8@J7(-6T/?_XQEKR.S8FQ[dagbgNH
Ucb-1(b]Dd.KYX[21TAB]_,C-\T]BBSLead-46LPI,?8I#Dc.HKMF@EI>CB.\8/4
J@2.2Hfa;9P)SMYJL@]8NN-gKS_K=S6JZ;+])eU)).F(]#M.E3]8]T8Nc.;=1X,F
PN8OX9f..#(P/fJI^L3913:#@R/Jf+504E^?3ODP)2B)KLc24EVX),-,f55CA6/J
9=3)b-7\/(f@1.#ML5D;WTbZGN#AM#JTS>SBO]e=UZL_ZBZ2I,)+H?d:,9=G/I2c
>Mg)NQD^]Z:CS[H4GEHEg_4/Kc(gZ?E>EK#Z=3SP^>;KR>Y\^61O/V8O58;9SeDN
a@O:)=>GTDL]6J\-9/;X_1D2(81WRBFU@UQBT#)V6DCf6fPF&d(+E:fSfaV(MEA7
=Z);#<_.H\J_.fGILV.gC20EM^6&dKVfWaEXb(^f7eaA?Q:f8D)7,(98DC6X18?6
]?E5aZP_aK#AVZUA3eI09[I]N=]@/&B:,QdGBcV,HH5d]Q-H(J?[Z1JAdV4RKdfB
.-MM.T/\NOU60(T+8IEe1[(>NF)5RE=(IS[L9E6EJ=S^-/SH_@YB1K_,UJZ8TG_C
HDOKIEF3]HI:Ef4:fX38CK])C9;1c_QPV9DNbA((HE]W]aC>1DUS97b-O:,.=UQO
?MR@HN?853&I/AD_&\I#6]D2?7B6K_[;ZC,1OAM.b@R\cBb62R(SSW1FAfS_3:e<
GPVF#eI16J7@(6I4TXAGb]&NQ,d@?bY^GU_KObZ0G9Pac@/]N(YO<c&=KP=/BY,,
:(Q/>6L79&c2d]W7O6[KE.1(9J3F;_LZ,cQ>QY=9L5g4YY8ZNR4UNC-,1Wg_g^GL
UE_UF-JJLRBT]aEd+.7BFZ<_&SbcdDTSUV31=c7Q\e?I:KgY_)?U\4:Q/#.S#Y.7
+7]c)/5VPXMcX3>Q?eB<KZ[#[::[g5.bA]#NAcL#2@UA7CT?C^Ma-@g6?E+R=E.O
S=E06-Q5WJ,Q0)20?Rc3[-Sf\5B@d#&E/QcVQgQT_4fc4HJE5WIBYHE:^.]@>FK.
VeB3YfaY[\FYg;E<eeXUS;225;DO9Y?1ePN<<#SQQ7V/:WKHXWCIP),RX#(G=/Kb
.4Ka(YM@(^4:OObN(MaWZXH3Nf;.();:55:SAef:^_Ef@1Z[_4/MeZ7g#S:g#dM5
A&@_MD+KEH8c]eN=_R6dgeAeB[dLRX?@8T5/^T^LDRZ:N#b>R[Va(^b>=gW4Y)QF
](AO7A5D6__2GV/SMdMKYG13Je&1T01[FL6,\Q&9\.0S)a9V))=WC-Z-;&d1SKM\
96J&HDF5e9[Ec++=>XH0XW[-9(#&#QbXM2D7fJXRW6Fd==BBH.+^#=/90M_U+:O>
c&VG#[b&^?3YV.U:KEAfUY<8J86#>SeGa>U791/B0:F;#F_).>QVDORZBVC2L\/[
/MNEFO99f.5]XB]+HX0ME\LD#D2J6eK593(GfW(HIL<.)M.ID8FD>F?7XdE&Z\-b
I^ZRQ]5#[=C<W@a40WVS3<_N54@VYTH1RJ.b4YS617JQ/]7Gf>,AT)\G6T@-g#1A
M61I?ScZ\+C>UT[TdGB1K=H,K9V#7MODLMcUa8U<N.SC65A8d^48g;L4ZNa-M#._
+1Q6Y[A?365E^-WK(Y+QM7[f@/R3,B3CaJQ_DC)=8KS]cE3(7W.8)Q[P@\<#V^T]
CU9/-[7_@]\T.C8C)e?Ff^]VP_5(B@1)dFc+:RCW+<+).a+>2JPG,:1>(NdRP2Od
]=^).Zg5]RUC:Y64<_Y.A&8)X/BK8/T&0Ca8Yda7LCO+AXIQa(1]>Lf,7-WLWeU+
BC[4O<EP[8^##6U>#I)UCOQNf#W=&H6FU/5-[bPTCF))c^DG=DVHO9OI\@Te@-M4
W@D4P8[6d^&#A0]RIWBZR,TTK+7eEOeK2SUY_]2]g4=?cCD,bd6b>[N/9=;d\XaB
[Q2Qg.&e=@/C&)OXZ(bc0K?I^62;;)1N+8H09K1+DK->-#+_A>6eMZ/Bg=/Y;US1
<>>1(=A7O220cfKE5RD7;LXdY7X7#_8(QLMLV[9<]KF.f)>8Vg;C^B&O9b7YW1_]
fW2ReAa_E?=f\B4\U]U(/86RQ=9LB+bS2/:]/6=O1DcJ<,GANJ<\H_FLGW/+6->Y
-=?,OAbWBTebHKE/<Y/)WGDIHa9K^&0M3K+aFeQC62[JVWE&OC]VHC0YSBQEOTCF
6>PC.U1cJ#XH3ND1JUUKDA&@e,<T2N49OW26[6PAQQ)=8cOODW[X>C_2R<?\VMF4
HQ5=<,PI1WIO7R((I[PN:?XP0TZ)W5)V7S7&[X8&8M3^bR]#9f4OA^WLTQ,)L+8]
G,9R_[H68:/7FA0U_C<;-<YgB](]JU/UNO-KQbZ9/bOb]g[=;gV/(fDQXBTZ3L&^
E2U/=?PPaREE?Y\aOO.N6P]Z)ZF4F>SMgCO\bM\UVAQ4aIfK\#59d+DJ9)-^3&ZJ
0+//7>_?0[<[38VP3T>8GZE\c79-_Y&FcWIAG&)&[[+Wa,;?3WGC2C.8@XcEf[,Z
ggLEE947L]:gfZ=.TO/QUe8Se72d:KN>/g&>_HX2d5BX&^/bbR0=K8BX4S9O/NK,
GMF5e#CDY5:/VZP00RAP=+PP+g=WK\?3ZcS.)Fa0gE1H)Z2PJb2L>fdH[dHIC&b\
>O&+geFXCU?g;Ad_?V.\6f;&/JX(685V5V209fb?KMZb&36^)P>V]bXc1B>)R21@
f/c_&1_6K&5HN-B9U/Rd^6=9Y:M:YAM2<g(W-FB1&48_3db>:M[Y>F4aXd[+@[@b
O4PfK5GTEK])=]V\IA^3UV/=1JVK8Q/ZLMBHOGJH?PT[P:#-f/C5R?Xf^e<4G+C0
+I.G1,J3NaO[5M7a1U7TJ.aGMF,<P[F+&3V7&P?_#I]GB37I\M0D4AKD:TX^6G3N
e@d]I+:HEG&;SJFM5LZ5ffc02a54g)PYKeM+7N@+K27G&ISC39Kb(DRNPe/_YfO?
;6U]R-Y0f@RWHL?CL.e7S.QB,^>3.9a3TI:^b3^g_]AVeG9:d5b>UNGZ\/KIC]RK
2;)&0=\[P+K-2.RR\(+Y0eIA3X(PVaL2/:g[BZ=GK.Ka74_QNG;W4/f2a-,G^dA4
e#FX);=:-Hb9KW&J9T)B6GQbPK<M<EGY>5@QIZZ:G:6K1EcTACSL=B.0e[<V^CUC
PeWGI7.D?/\=)9#-/_8e.b/:M4.NU]D[#OK@/O#^,E(f:JMSbHW,YRa,XX8La>OT
J,?Y:9-022]4UYV(FDa\Gdd91E<IY5=@(=NaFC3)0A]?13L&99&,2K/&SIU5]Z[5
@Me?:ZO8RP\D^5Z&::^U#Xf<8VZI@9N,/T(aRVKYUU4#FeY@eN4:3>W+M6]]Ke:R
(>?1[[&Rfg@6cb,VZ#P^+HI8\I:<?Q_.ad8LDZL/^acQS:D25dTAae<aL_U#B(E0
dJ]d+;d@S>RS>_#IFC5@UXI_8WdS&Q;\6SVU>0DEfY@dIP_GZ,bIcIQX#O5/:3Tf
\3OJFG6JF4LZebTYN??+P63F#[]cPge=G)?ESHfY+O3Bf:(K:a=P&XXTc^,S9S@U
]FG-IHe>B]QZ]K8@c:N<_7,+FGfMO4Q1c@7]S(OD)OQ.9b1E:(J45W2:Y:?EX[eS
R(<HeO3D?7SZ>.bda0P.&RMYCPg^\g9PQ3Y(J)-BM.B<(6c0TY_(RAHMBY;HfZ4N
FOFTeaR#OB#,5G(+1FEBAe4A9c[)aCK1ASW#<9&#-f;?>C+H/fXK))GTXC9J8W:g
=0Q6Z:F5EgG[g?CB6-\HeZI[Z5a]]Kd?YG+2@=W+.;Q+bMgP)H(+JZ)g..NKTA.Y
;(J,@a-7FbMe<DT5(Q=HM@f90c=<;;RC8Y>:9X_&Z8LPGVKHE1),:g^@VG6,R&1A
6(NI9,3J,_[-E)3EZDf,45E3b,f._U,5U05S:@EJOX#1FV-dHJg>7HG8+GB1#ED0
(?0\a/VV1ge_\Rb?[HcL,4RaU>1R(Od?O-48g\[)Ya(PfA;R&?^Z#D/;@9-cS71>
>753>ObaJ>aVF[bdGB[K<7<Vd&;Z^1S@Gf6,X30(DH:DC<R?,1_QLU+#W)(J02a)
7;B;<_bWDSV7f?3C>+/>Q<K_Y8E1EXO36>?agYPLA-?gSUOSf.;PB.SaT3D]bD4R
35(5YQNf>#:c6,X#6-Q_WbgdJ0@7./c:#2XXA3\@#a8=LB8OM0@D?P1IM=]>\ffY
0G:GLVTa;X]^gKIfG\+GCR@WS^5f2fa#^KR+EAA^e&(HR]9T7K6\,A/.1a/.1B;I
ee<2QGD+0L998+Kg?,SUA<.<=Q@XZN.<8M6U(EBS?b:(8FfZW/TP&(JIL>&RfX2)
3?Z[IQXN)/#e[c)8.Ae)PTO\Vf8I91<gW@#6(F(T&,,c^3BWgc<F6-;RDG69:6ED
CH:RINV+<4K_0)H],:#2.SI08[A5PXGDH8.?\.+^-&9?0XDV4ZT+\g2aZ?K_0&3N
GJGVE=AJ2NS[gSK-DeD]<Z>CQ3@a;^Ha+2HX@b6bLaCgPdMcVM0\./Y>I;7g9K@9
a:?0N&43#CGb)Y]4P]-a(a>RU&M.YDN3b)-b;OQ3YJ2PX8EJBgJ?:dHWc)]>e:d=
B-#M<3LPF0WE<?IT(1cBA>)eOAg:/21-&=,ZF5^cA2N]CZV:XHFe>UG\d,@EggUG
HTT0H;IO;)9D&V5bgS[\GHXeAHaSJ\W;QMPWZ2eBKK;#>.;S8dVC+XCE\G2#TPe=
0_R>)fe278I]35XgLb7QV0CZ1#B/S/-V(QT5aZX??J_?A5HU\J?c;ZE;Z)X^Gcgf
g</&X3J<Y]a(BG#-[>#/::&B<.RWc#JABD>O:<e+P>V-&cH>QT0#Ta/e6Fb:YU6?
Hg)2QWI^1G^2+)g_C5eg>B,(9P]Oc<9RS-J_F_P.[Sdc)5Nd:^96-L2.0G7]5>=d
I<M_NHC+M^23M?<EILbVH(GQDS@&GN:GE7ACOE031cM9;J.<:JTa7]S(=a&=f@N3
RSA4-P.D/PD.1:dM>PINIDR&HH10_#4A+EQ8f2W2FO2(JP1TAO[c5O5^GXL>B?2B
9(;?O9R_7-Z3O=UVTLNJ.-\#(0^T/P9_b0J(<\8Sg428&)VB^)gG4UGSa>^CFC@@
)Y0N?L&J1G3#d=,=FH>;f4S>SJgX,KD;<dM9YS^K]QR0>_W[JQLY+1.KK2fHO57:
+(LDGAW[O=U:R5@gPXX^0)\7=bg;KE/VS+eUdCG[;<[Z?caKN\2&N7A2ReJOT0Z@
F23=(ae&W3a5S1\I<E:.\9=M/6TE]7TC<<VC0N+^?dW+g,1ag<;W(&QZ?W5&KVA^
?1J\<QJJ]C2G6g06=JW):WVH._YGOSF60&7NV>8)=W01VH64Z-5bDT,[P(8]1U._
QS3GdcK_Ef9<df:A@faY,FKS[&IO.8\T1H<H@9&,HKc6cU->4CITH<R#R(23)S#e
\QHR4B,1_1^8#W2SLJe((<UcWWgK5TgF@IMd6EYUFVIWLe-9Ee[&<Wa[OQQC=?49
D.:9P-4Ea-0+:I)W/b+_6<,?NXNba\H3)d+)=Ed6O=GO7b;[MC))29,4cRB:<[\c
C4L9K[<f>CgR[2[FM\N8G[/30^#OP+(UO>2@^(^P6RCF<ZDJ)W&D\ZaSe^B0#]Ua
MRMRT72S5\THd3X;HfU\,ME_[\507.[I)7gQ<G&&>BXCEC\d0A_G.JaLST,<\9I,
T/F)\#269D2Tg)94QK@>95WC,VMH7/6/>I;<;cG\Xb#8L(ATAS7<gLeQeO7QZ@(E
1FG=O5Q&,cd\WGX/cQGZ?c:@JEbUG@0?HY4McR8d>UL_R>gJF1-2\@RDIEK)GM[;
/OPb8\E(eQO2c;,BD(=.JAAC/^7:FUDa)eT#.S-3/9&==^,YN7(^E>G[cWd_)V5e
VJ8&\:2C/.JG.b@<I@0ZAgR7S.e)d;U/9;P;_g)NR#WKCcFZ-JB-H\fV28\:]I8G
&LS#/]_2;B^^ZPSTWW\T5BN6(12AO]dR#FQ41^1@EX?4d-Lb=Y<c0c\S8W3F_<V9
&L6-@@92+WY9FTFPWP+-#2L>.0+PWZ&TM^RLJ+NN^EV)@LW:V7c;?,5X#IH#T,ZV
_I,6gOg-fFUCZ=e:8-0WCX@Z^AFa0Da[=7++NIb6<C6D\&A/-D9:][eH>&S/4]/W
(N=;#&FeA+LRQ((_#X7,(_>_<=EY,SQ3bKC69DcW_J\NM?5HYV4:7;^/95FVLX:&
aEJ#KLDJP8Cea,Y(bdbb(I.^U(7F=;F;;R041H=RaebGf7.\OF-@)#Z-EYJT>UVE
\;>1aB<2&R#<(SZ#9R<A9+=N+1c\bFRU+NCf.FG]D-TK4^3AP)R=<R<T\9:>6T.e
?Dc6EH;.)@VB(KJ;IA(#7Yg^ce(JRM_DQJR6<RRF0_)e3a&H7[_R[#55CRbH9/[[
U<Q3gFcd]fTLR,T4UB[dYM4H-&5(W0\=6/C0TLdPc9=c\B5@Lb,,L@81]OTY[UFI
e]dP^_2T@F0)O@0ZN+]4D+2UW72X#RK8R@cZMXA&Z#=<CW#(JHF1QN+Ua.NLe+>2
4dP\1MIgWO=3/BZXJ0Q,CBa0;cYLD(G-A+NB)K<cD?TLfKF<Y9=6K2Q;-N_f+^VT
]Z@[D=aUN7R,Ve(e5eX4GG8JQT/:Pd;Z(WYD\DJ0FV5PX.=]@bK+C0:N3C/.eC(a
5A1D(D=]L-\XLFbfd<X1b(V05_R]Y<VeT>J7.CJg<_&T7IOT7ac.9/#W9Q<g9gbW
B?X\34P3#Y=<fBQMSCVL1\2IUV;1HUA4VTf0bHVZ.8.#b&H6FZ]<:B?Ye_/D[e(J
Le6PWN6K:I<+)0aZRVH#aKP,(.fdaI#80dV3]&B(6#O5aY.;,YF;aIH;8[/]dRYJ
6F#R0#+0K)TWBeN?)_b24M7Sg#QS==N/B#L#@;N)75>:BISU&JHTKP+K>bO,Vb2W
?R=RHEf9[N\[Q[WD,86]K2R1#M^E(0W>]EZDU+43aWZSbEULE.D^@6^\T5J-6S2B
J;e)I6H3@bce3\??<SV94f?Dbb0)g.OIg1-FG6RRXW625<5R&,0Ua\=#2@Y:H6G)
I+4Q=Y7(Z/Lc(YJN8^QZ,Ggb1M:6AT6T0,2J79&>NEe)EBA?\>K56V,1Y5.:&HJa
A@S?C@?Y7Ed6[DCD5GKVA>Uc39UZ(4?FGC/bC<M0YV+KR_T(&BFNbN;1Pc6E6.8G
Y.WAJ-^QKM[ecRU\QQ=7A[4-=fF&QQ_?9f&)+HZYTYV@:-2BZfO_D+#E0ZL=(K\J
S<2TL3R)[e?EaZW@PK;TB#DL\Zd+PK6R9)^ZXKd(VB?K^2^.O0;A^P[ab)HS_QWJ
c2^B95S[J9Ua?4?;.EMF,>3ZXg2=T&BMVO+JB5+9&@\8^H##QQF+.5gC&deWd6If
0?Q-XPd2)B]T\DW.:d6X6E@>RDEYRe/BT]Y,<66\QNN;fQSMU=DH.679ZB\\;[XT
I@BRKaYZE?e;3b#T8YPE7-[>^,4(\bc4MSCA4d,&W&/4FQ#-#b@F\ZUSeZ)H<f(<
),e@=>[f4SB(&<F/bZ8f\9&e-a&S=9E(D/JGgc<_B;(4Ug-NHUYTJ:HV-1b(?_a_
;I@S>HU?:35/7#Lba<GTG30e)RG9N2217+#JZb\c9P@AF((G4[##]J=<;R<)7cd\
aA56Rdc5?P-<:-,J]d8g:L5@7W.A9Q1.=]RW9g?fB47f6Pc@DCD@(+e/^CX:fQ/\
+3<<VD#<?,Q2^I627;J4JaNA45#OSEOB0T0[R/]/7WEdQ2(JO&+g>YBg\1WJ>7M<
;QR6Z+:6&3=>G/D19(]DaYH;g2X^eYBG1.fBcR/EOZYG\f<8TP9@U_S1Je4W_/L^
\K,Cea;FgD?,JAT:^<UCA9)9+ggPGBJX&F3)74,@_AN&#(HOB(PA@T]PES@,+0[C
W5J,0LS2<#L4YW+YU57..S7HJ)8c@\9Y;5)L5M_@;V-cJ[S05eMC/V#b87LKF3?G
/-MV,I7g-0D_CK-<\G4b,88#d]Y<9X4Y6/&(6Vc8G]affI#]0B9>&8^84#/#:T21
;@)\B6TMfY?.W>MU^#ZCVV;WYR=YU_I+B04EdN/_/F/]f-?/]^C?JO7.@dLe)<#:
YGP:eY/DX_Q3A-(,7a_Ud)<4^P^WY]I[U7Ze.:>4];][R])MH2^QHC^>R[;3BP#[
P-R6+0:3=Vf(5#@)Wf2g3eG9DKdec6d0=5/:fdV32eaIc1M8?-ANHSMARcH>0S[V
&aS&LK0DNYUHI->1N[JfFdV>;CFEH<M,Nd_0/>70a?VIWfcGc&G&QfE-YI29,)Ub
UWLWOKc:4Cg^:U/eF1R&bfXF^c@JXdZL;#=^(?8J)UESf8F.TYD^Id,7NG&CSGfg
91ZAa91eI(@2B6.H\_&ZZM?)BbbTHQPbBc-_(>4IWON_#1fD)_Z@>,J<+6;?02d:
K;X_#@?bMZdAR\(87D>=cS-D/7W501GTPe^6QK-A9Y9CAQaC-\N6RF(@gP3XTS&F
28J1IcO#VY)T?54Y.GTZ7J75&ZI(VIIZ)UL?Z6:Z8@CHI/C]H.HgZHI6gaHc@?O4
VZWAOH3@f<FQ9@+/(:P;Aa7a+(aEZ@)\6:]]R2W_B_UgHN^D^SFAZKN5#Y:0XM85
IU,W)1dfJ#SP+?)I&T#cJ&\MD21De75Y@dNAJdUT=ILKT,a+0KWLH87Q=cFN1?2X
#1.ZV,eaaEgDZRZU=??EOHd7DF<MOX0cF(X6=P+(^G[=7>8OEcC_0VcN8);5WU[H
==D3O<C)g7E;A&I-[+_Ea3GKNcG,.^H-=X0R^.617=4M&BNN\&\Ba^RY@YL#cJN&
#4J)gPAXc:fH>Le6d&(XYQBOb20RYV(a,3JS\OC(_..U?-]?-<:_Z)6H]YP9AE##
LgPO(Hg,S+NSfMK^P^6I,XD2<P[Nd:E-cHe7V2.Ta92HF)BHf,KY4PMg^U3GM,5]
,74fb7@ID</fG/Q,7bb,,&EVS]7S<_VaZUPg7#fQG18;UPSAWe<3DJ[d:PHHZ._G
#FA4+e5>Cc@Y9W31(IABG6E)Q^<b6(aYa<@K(]Q2?^9-<g.IIIV1e#W(V14ID)4d
/+BSe4LB8gYUQLQZEZC][Ra#,1K_COQ1B34<^;SQ.7W>eU<]/>c\d;L64<>X0+c2
OUQC-[V(^0\f2EFIVg0F=(YN9>Z0@a(Jd=U]TGJgHW_&P48I;F^UaSR\.?]/)9JF
aZ@B=]HIe9KN9&RG+5=C,0S^7Ec8f#g\5ELgZaTcJ#gP#RcADSBbSUaFG;5NS[?Y
cOS,HO@C]5KDQ0F0Z]7A&0GP<[d?RAIHTNV)XB3EeeMT[fT;]TA.0W,#.2gF:S#2
XOCdIVV37G:Y5[0UW]X,RQZ1Q7=_YUCPG:S7N;dVN0&=,JTDNZJP)H(RC@/H643#
=,=1[0?OFCQb=;<SJ/b=a.>BEFI_/1DV9)Q?fMD3Rf,#4L-[0CdP&3?OVf=GMcOX
C0I,U3DSAJ6NO]@Zg=Nf&;M=T_L5R7DPL#D(&?5B6NI1NM/9EZNNG+:J@IM1fbD,
J>L(<OVZX\JT04a&E&C&g\JJ&]+7E15E62(R/,D]bI5#]MAX,dTXef;0W(,Y)DS?
d;]6HHL8EAHOT#Hf5Df[KC7U_fVV?XF.Q^U+G>f1H/\O(]_ZdbF)cGfS1-dV#W-,
L]4.7U1I^I-05[I1D6\IC1H0fVJDg]R6+D/_XG3W@FUD+>7fKd6Y+C]\cWUQ(Ba.
;gW&1;:D9cV,,B6RT]P#_63,S2,\.c<05T^ZR[>gSHPDD>=F0?bPYF(V5-9NE-a&
]]g?G^cE1HI^O6KX/1KF-\EeDba>0N=BgMQ^+bY/QU_JDa6CQB-H:]<E0a3\c.[U
^Q2?&PLL+b&TC<IBWgZ7=DdZabA8XJ7^3B#2ZYUf5FY;S_C;&b==F0d70>AN]/aG
[0/c5NP4LEQVIZ8_N1g1UfC=8&0:c;?W4f6YR#fgE,F34JC;#S6II=1A>_52-1M3
V]I?NQYR:2cT&:+V4Y>AWfGJ_B>:gRO:Idb:OZXc?g[_GMWb7a[P:4.94-]1]]9,
1;)3;0F=</R1^TO]G\DWW;6O7CLYM@#d;2\3]ORN_AR&-MDP;M?U\>g[BGCM1d\@
BKINa>-8,IY5J?Ag<TM;2G85V#[YB@UaA\8[aVI8@7[bVeBBF]6a4,:cKV_cF[3K
BR=JZ4@_AED6da95EEI8)9OOgbd=WSDWB\2&BS;RPG0g91+DG54G:Z8B5:(A(#;)
E=4d&BD)1PDEPU@)P#R-^]E(2([M3G\WO[V_B&6935^K_^W#cJ2-GJTD/=A1+/^<
(5Ug66,bWNC9?dC;Z1/=gL[?3,+#WB[@LL+ASgc4_62LF9Tc0.\F:<,b4^TEAEI:
-(LN>Q&f,</EA&A1AU>;JTNDFCP2FR?PV(fJ9^/6AQ9bC?J/S(fCC5-5]BH>8T;U
gaIG+5X-O)YQ;cgZa0f5<d&9)>PFYN]XXMN+bgL>Q]0.f/&USC<&b=f.M\P7K@T>
=A3D(,=8LJ?J/K9ePBfE5H]A;E0.2\/VcQG5F;/5Y=Nd(Y58d1J]^gbTfHaWI:IY
VTSX1g)J@8H<I_gKeAbF53<:U=5;.@O-cN-12^cdG06D_&+]7:UVN.<e1adRM0fW
GD()GP]F4#f1L,^bMb\0J:DF)^_VT5PI@HU.>=/8f]\Bg#AS?7f?5P&9f7>b3VIE
Z2MYRP\1A>4B9)?JL-L1NAb5YNd-JE3:@-U26@HCKg81gP;^=_HJJ_2&\)+]WFH:
SKL^9MA0-RMDA<L7C5TP3-g\a>ID9CHd91_AN5gZUZLWAOA^-)^Ec2[#B2I1P)K1
C\=1b:^HEP].Ed:g.E)>]X^^>TZg4)_:KXBF?+,AIdIA4W&Z#f8LWKV]DEcSe[CU
M:a8M499Pc/U<A?-RI=)2SfZaXU7JQ3bFT#7[Y9HU^NMKT+d:N<MW?NZCFS-g30U
/0\HcE70Y9f8?Va7T/-Ba6V5c>?OfNBV[_RC9Z=HEE@gV4^J+I-I55RGTNN\W420
J\EPBgH10R4X=7f&I)4[1=]F=IdR7NY>@9)E)7]GUgCZc3cB^DcWYF-gWSK,;b:G
#IYCQ1a\)?Z+UE.5BX5Y@.947G0TH/.Tf=A9(]H7[=&5V-;ZdOODVdPMK28YHL0T
+gfF2c02&=X\10BK-K(0[AV;G;U(1FD_Y0WCK,a=8I7HXL<YO74g)RDCN]#[E.N0
G]O&&]B6/fN/g.UbEgL9;S@g&#\^Bf+Y;M]ce<b)XeDaE3@CeP/)fOLaT,[\-+Wf
D0PfOEa5N:+)A(:EPZT>a0/OAX9^W]0eb6d#X12LZB:V]NM&c2WHc@.]=_57)a3B
\b#E/.(1d)caL^+TgP?\Rd(858WbD6Y+&)?)5L<Z>AU25R.a5F.9<JgH?^[SD?0=
CD:)gOg:1OIM<Y]#4]I00BbRMeUgLM/6F3:&[05WX?0dS]0^ROd3YX4\0)eISRW_
G>XU#^e7Pcb:ADd9NC0=1]MNIG9W-O1Sg?2f9eN53Y^REH-cGX?\ZACE46P[@AP^
AQf3;F8)6QLI-YN<f+<)<Dc_^]D@ZRePdeQaJc5EKY;Cc53D;Lg3cI(gHG5YfF1=
?1SWPA50C3K+KD:]a+MNXA[6;LJ@]+JKDX&B2[D)F?^b&K6E22-W-0U\&@6TT]LB
BZ-VPC\D]XP#?]bKEP<P.Yd4DSSY.<<9a,QF@_3S0<]0OLHc6-[DNRd>8?N?E(/)
KKIQ^W+_5@=DB,,d1H?M]O@()VWMG1?RJ\aYGOgEM_aV>0VY,?,)59+S[^FDFT88
OUWU,fKA:593OE?96^\(U6Z.-WMDGU.c_J(JR9XX+D+I.&_N7\;@U4V_I\+5^C,F
f/G/@G:[/8F..8LJgHUR@QT3=Z)dVHS=^S_]M-&4KfaM9\]=aF,E60LcX+VLKb>M
,#Sf:=J:4eWXE<657Tb3b#@\L2DG[3V:_7e-eP>CYMG,&ITKO^@&S)dA^LUA>2P<
/OdD->dVMG@S:+OM])^CCP6/?AdB@+^(0;\,@^\13-T+NMNAAcNP#MFFVX\6I1Rb
CcObFE]CZSQdH7<^8)g31-0=WE@L-^:-e<>/->VX6&US:/;c4WF[?TPU)P8N07R1
9,U@AM-\P[6Z=KW=I&LNQ@O/0P1\_=9OPeD?MK[LLL#BRT.^WfE/N-aI61]J57V;
-aGWQYc=>9B<4-8eR.BCGBY_[]\T)0^^9IOLGF#7?B?-<)YO4?Q+<TbOWTIX^C<9
,,SC#0AB>DB^@gSZ#PB2gQG=@:WCF-+b/,GU5@O1I&P_\@(eP9c7#_cES><[EQ0,
2ZZ\V?=SX.,AS))P;-fX+[1@^#39fU3BggO]L3:c;1dZ,Me\TUg]B,d+8,01<VO@
dCdeVCI;ZaaERg:Y,?T/6,4E5&:4+EXW<GP,6(@NXO_ZQ(V+\gf;NZc7:JFH\,6-
49M<WD5OUZH^W;;fVHW#cdL1Cb&.(Z].MId:AKAOVVe5++,FgQdH=V:=2O&L7=9>
\-#,MK7M<G6>8N_6.La0_4bg-fSHd)W[R/AIR5=g_gBP)@0fYeQ8]?[8<Ra,F_de
dcP&3#ZVV;Zc#ACR>a@=<f<(T7E56WUB>G)0Jce,MBF9Y>Y2LU+3N6,e[#F^)f[b
J?cMfI1;M<W6SQB31SEE@Q4@&cWZ.+HL=&ATHN2gD@KfC&6c8WHGSe0Ib2Hg]Sf\
;;+59U,:M-/XgW<_K,M_f[#LH^[32#H1>^?6RY=)6X#K4ZV-2T132]NY&9AP8G1;
<b^];(9[_&YcA0cMU^46A/X5aR^D6NFI()R)5-OFH6_e\&663&?(.5N]-8VO:Y0+
e5Q6Sa]aY]>MZI@:=&V4]7g7)U6J<b]?@F(ZQF+:\#](ZF23<#b-<Y]I2f/X^4Xc
X\LI1FHZX8<b[Q(.M=]RFDbS4&JQ7e76>93\:U3635(L([T12CC])N.M7RWUgQ6J
R/5/T]2<Jgg1MRPeNH]=#?OLbMNN/>#R<;-7HW/KW9DN(R.(16;=G6[6a?N>c/4b
[#&Y<W>M)HU40##L=&ZDbO(M6>I,YFI56Q<LAX>g([a<NOY]9IYVRX7OMZ?/Ff[6
B94c;3.gVN^C+;#VQ[9TQ>@[^5/:0<\CQ+W+AAN)G._91MI:[fZ=/>)E)a:<XS@c
0842M4]66O;NZW2=Dg[S4CECgJ&BQ)g,N?Yd[b:OcB[+LcGMB:AB-9beY,G=GADI
.1E]P5X/_8=>dffR8cKQ:@Bd?2+NO^?D-D&QTKQHRL6^DIJX5JX;gED^C&>MXED3
/TP]19E#^_J(a8g?YFNDfO=eDK[O7bO/cf(SFJQA25]^:KT/>\0+,@7Z&=3CPFNF
DCB5>#7[0Jg0af1fQ.O6U6A?cZ&+V758@,#g(ODA=4QQf5FQfF]EE2S:T;=^X9Ha
&N=@&:<F3EW1YQL1F.93?HFKH6)JZ@E<bf5;Q+5BfE8[SOLIJ^L-\T;IRQeYFbHX
[KEQSBB9XJAC)XWf-(?==@VJKOD<X=/&7ee,,O=6KG_A^[IW]5[Mdf2[Cb7._?XO
E@5))CGVWe)&P:H++)<@)+U<7dEeE<RO^GNfH_3[5[cJ([_OR:\:75RI<FWX:&)A
KM-.0VS7L>f1E#7SJeN?[DgLaH48&ZgESAB2B+3LBZ7C]L\eB^O(ELHX6BU_5W\b
0Ba2#T@M1C=MU-SAM)dI^JF+J:NG8Aa;ZR8.AN]Ta^50T;#WCb(9#K/)6HZ0OTT_
c(AYgHT.P@He?gN>IJAF:YJZ2D;94IfV:V:4_cS\_GAgg#U(/_/OfL+(_2ff+J_K
>TALK25Xe=VT8+=-S=5,?Q?Y\:HM&FV]8ec-\ZW(3__,OGId[;1AWY01BC@S0/-C
DeZ\fH^BXVbY3gN>6V&P9@d816?b]Q;^dU3b-VgX>#.95T\fZ(XGg2H=7^ZbSHe4
I\f];e/#F,T7gU?I[;NY_c)51,)\K/NA(I+2MBCVD@2K(De#65YaAcIScQ[WW\,I
1JSJ2W+FB?L@e?4AAV;VI@/-D83R1#f+=G;b#(8O]427B5\,B4M-,D?edfT-K;^2
&VW6cILc5&_U#BKb(QX)<d2U5(Dg45[Zc&+bdX2YIY/+ae4J7-@N)KO/<=HI_g0,
a1DB(JK(_K9;GeH<7XV=R3#=M4]C+&YF@+ZaPR8Rb6Xfgce_O:CR:W+LYc/agb&(
cRLe[I]IEKP:YeGMJ&A=^3)X:CNb]d7EM(+M[9bW&#QQBKbUfRN,NCHCEE#1^P_:
@fJ[U_4,9GG^3JKR-T>,TVE:a0S;2H8(5FdSKED>/NATYO^Q:f>S>D]<?1XLa@:f
V5c=F1S(;#Gf?3-IbZGZHd0?QU3Vf8M>P@L.0(EYIENe-cc&@DCTNQOGN4E21U#1
//8CbEf,NdF7E-#PFLab##A+<Z6c?fF#K^2@9VA)?U):_[L\GAYe8R/@??2/)1YJ
)W8KD\UNJ+dL=[aaC6&b)PS&JJ@<_&:g+d6LG@)&8](OM,JTNb8Rdf+;+Ug#e4fe
S0AZ]cQ2ce<(CQ=OcM>),R.@c@0/Z4B@\[E_[1T<5dSQIY//6JN3GXB.3>9I\1C/
1M,9[8^X=K13OH?&4-4;KDf8NHYGBHFeZ+daN\=0)#9X@eAMU-1(8a=:d,50CD=\
=4=3ETBK<:2;K7_G@_L/D._WJ7eD&+[BCdZUdA9<6);?a+6EEQZL.?f,-EZNKf]X
If,^G-RKMP?VWY_5(+=QbNNTUaJ@?eQ(f^P_:Vd@)@HYYJ-5c?32UKd]W_K8TR)C
WS2]ag-ZF/[48HM.5SN@VPCW&27-BJ0?2W::VVB5\b+9RaUH,J^;+J5DF\,<e(.S
;ZHc5Y\9)cGcP<3J4c2GOSPIgedHXQCN?,=-T4&PF1KD:F(RDL+/5Ba1QSXR3Q34
U=aYM,4K)^Z&9@bL0#Nd>dc4J;ZGNeBXGPAd@[JCQ-8G;&(g8931G/CQWF_YF2].
_@:_3]]JU6<1=:23C&UJDE9VePRW2GH8X-YB=_ZF))3\H(VNLg@2F8_Agc>F;UZY
U:74@^H?YA.=U)Oef<KJA9_;fQA<179^UM28;=EW#7[bg/b/,;T.+:acEf^ZT86I
-??[L4U-X?AGB:QOHeG,Z]a#aJ0[Df+ZEVVH04V@@A,OYJVB##EHHg,U.\_[32J8
dAc9F+=>AHPK)TT>TgI)K&U<\,N3FWaM<XG?&9>/JF>=LB/6RaceVT:Q^REL>.fc
IY@#?6AOS)E_;cVM)J43+^E6\BI]^3<6AWIGHCg+\4MNdDAR&?(8A-7A=>JDbUFc
eLF4QX^#g?3Z66/d(JP55^b]1SK+J1W[cVU.#V#c,0?FSU8\R87LYFAKT(aT>)OT
J_5Xf,LJ7c8]_B0R94GI@f_eX5Y1<AJ&fP7&1?#6AOG,Z0C/5F7OY384R_9_b_PN
&:[/7?0S1I-CI\\W@8PHX1XWF32c/+VB_#BU8FKA[83DNNfLQ:Zf+\+L+M,aL[bf
#]H_73(A\T,S]c=[UJ<W4:,/be46JVRd)#N8:,:9YVOYZ,G3.35W6OQDMW1D=)5<
T?\d399\T&\<U.?Y-4Wg:JX[D_4R?H8J[E-;_:T]Vd&SH<MC;fBX#P[MOL+\V^EL
N_5=.gY]W7)_F<N]CD+MQA/gTDMVW\TSWI>=^;I514CP4FK3O<LNCS=D)@/]MNJ8
00E[Tb:f^C#-78&H?9a/X)B7Y2MD-#^RRe+HOO_Z+_;36XO:L8B]aY>OADdFf2<7
(@LK.HY2[))>UQ[?^e<CcCU#5f<36\[Y16K]cK5GN.BG:00BBXQ,LdHa2I=K7bKF
QFZ(b.C&EVD?V#+4?VcB2DBN4S8[S7-b#cG[@JP<RCCBQF/\:WA629/>]/-WT=H9
I]OL\b-QKK\a2]K.:IbEZb8BG8_E7ae2/J(:?)D+1#D1+=(<J8:f8A(HUb=_,MK3
e#5\PNYaWEGYC1U^1&RPTD?#9O3d<PE,?,agP30HcI4[KE2/J5gJ\.eU8[I-/)g_
Ng\dUEe9ZW(7bWW+?#TF]g<NI6W-P:P=+4OR17HI/9+FSTP7RFdd)W]PK8:S\@)^
APB\J>M,M^.T@WX4_dQ+#GI])G7PU)(B25gH\.+S:J5U(\@AbL,^Cd7XNLJBCD15
&XDb[RNO)UbVGV-TJ-A)=H#^&X#TZ]gcF99U0I@07?IZdFW7\NeI>W&VM5X(P=YN
P[8RRa8<f.Zc:68>0Ja9UTFOgfGaLI]BJ2?XaV;Tg0[8b;4I^LBIACZNSeY\@->e
^P\5KCI3:,eGe(3IgFeVXe@??F;f5)2.1<20(SPa^F\CaAQ=BPb93XXPXHMN@W2O
OKU)3QB;9LO[SFTAW([cc(9,2ZTJX54[]WO-/\DUUU9KLaF\Y;^d?Yaa##L/##1D
ccN<BRQ/@fdV[S8G\UDYXeN6T)+P72304VW&YJ-7Z16Q[D9MRgMO.Vdb2eJQ-(#O
^G6-+:E\c\L6g_M4#JJE@_R?&b9Bc96=GgL(6aJ,7OJdV.DY.g<4=[:A6.J=gYD5
+B4Od^EFE&7JB:-3.G7]VX>@Jd#T6df-<f-NGR8_5>P&,O.eSNea3@41@L=#C?-F
XDCF.MVLR+7b1e?;ITO\TNR+()#5((H2?3^89S,X0ULOe7]2\b^:+P>T>[dXG;DH
4e5B&\[5XR)F8T&Le,c(Q;A=L+&YK7HDS6SJZ=a#.ACcPF0N##<&,PJ\P72X@?HI
;>>R^.^<_QSFg)Z471e@U_CLT_GW[3&1ZYV47U(WI2/(F95WA/KMA\#7#0&ZTe/b
(ZT-/-F[aaQ.K.1JWOIeG;gKIgYc][@M5/DXXSaA+J,BSXb^2>=OF-8EG#H[g:M5
gPTf)QWQW\/d-M5A#afCQa0e>KJaRKYKTcEC4J(/IN;.UgHFG]UIc#d@:5QE)WJ0
_OB,7[#9/^b0-C3[ASZV)P0?2:.-H6WU#6@2^AZZ)N?W7<RFK3CAg>2;ccf3GP=#
\-c(LbD,V^YG87FD9RQZVF<fTc_5\<Q0T,N2&TbQaNE#B4>B:NPb,g-?(0dV>V(<
05d#90^G8DIL[T<[/M-R^-[5I4D8e9d<8;39@A]5LdI\5Y2B4bM3b10?_Tb7[\ZC
,@P[a39^#\D[>0#/;1d+EaJ9VL-MN;>W.&J,3gV+++B=;;8,L[cb06MT+#40S3>a
[#c^3,)dU-J.LL0UfSf9?]\N1S=EUS:;0bCZ?VT;JL+0+Za=APSf[KAQc@WGFcHW
P18Ga39\^bd+I5c0#bU3>0&g0<G4/N=fS]?4MXF39c9+&Bb_)/ENV.#c?0^YRNUA
5EabG.2;e0dG@U7/gdNDE\4,;2WA^N,a#Q_0-b<[VbQ#+UN1LEgQF;HD;<M>B]DH
C?YAe&(@X(0&CL-fLOW2PbWDD0eOW&7?^7O_E:V5)O=e@5,.#HW>3,#[/9#6Uf7W
)Xa)=K-9:ePH:;7f<^aa3LBFM5X7_./V/0/F)1)LV0?O8)A3W(.FOCD11DfO-f&K
bF]6J2S-K/;LQbXHaFgFd@X48?S#HdfL<aJC,CF/TEW6)>+#T294eGN@]FCZX5>:
^(WGb64ZL57[77[@UO5:C/a12]L&J#@BD<-RV,a+d\6,R@-PI-TD2c<<(A8XI]J5
F4aA,Kd1ROYDLD[T;+-4Uf0)D&b)GLBRZ0F^=f2DfDBR)J03BC9\?W48?^UT7PII
JaeTDSc87SOG#_[6^+E>O9K?\4(3YG#29HJ4)f/X^[2@#g+?TRX3K,ZC4A#a4EDV
F-BK3[Mf119S\=beaN626K>?6DV6M]eCUZ)T6B@?VMX9gOY4/ABSV6)f-RER->1@
7)GXeT0dN3Jd4EEVFdQE>X1ACTIN9;4-K7:(gJ:Y8^PLG\B;Df2QZLPRO:Dc3RSH
+_B&a5;?4EAY-HZU\_UVEW^JSBR5OKecHWNb##=/8/TTM]@XcBM&RaSC8ecTR[0S
gXcVMBA-XFgKE:A1?L#)_/6R4MC[NP/\^\XCa5+afX1d#+EDL.X_Id#BAJ>ID6ID
cR0=.LN&b3,.;4E)R4-3M@Q5N[:IWZ>J?c@:dfUe,7+/BXI-XEf]_B(K^O8869c5
>>gOPK,X1Ue_LWEG,,78Hf4^[13(^Ng#:]8\^UdUDTI>A+W:Y[S=F;+O\aF&K#PH
N?N::>BTXNX:P8G88\N4E6+.=MH_F6Ac8&&aGfCMcW90@d]ICQ:N1;T[TV[d@PY\
Y./<bV?1^@,Y0FKUN[>N709Lc<UL]<cFH41e-S[G/gC953Z];7aNQ<)(0Ld49g#d
BeJ[EQ-aVY:.@7cY_6d5RdZ/W<@Fb2N\[?aaQ72R_PfEBK,4JO+?c>84;c(Y.bSO
V.3QP<IPOX<3T09SH87W>^=&O,,J2c1N4TdLfK9dPAR,(aDC17F<=;.e-6\7K82B
#-)Sa[gb,Wc17B-5#OaI=Y8C1PaAYJ)21=+1^HY=CUH0-COg@RGKCSH35ZMA=0c0
TIJ/Z@c;aGB5JSI)NW3WLe_J#Y,X3;^8O^@/@?_[TYYbEOSD9WH2b+0YN0T/;[1G
eT^#@GHbK&bVKQ_M2fA3\[#MVc])7\1aTcRb,)LP(0G7--^=88OG>4KK<a+?B/]5
,IbD,&@Z03OWUH7LJa,-MbV.&,CS_4@I7-(-4IH&,SF(;91;N@.,?@?)e.[fKCWU
3J/@H(9Q-PBO::2&29S3>UW_LL/.H>S)[K@=^d9>7EO30fYLJ6LT-Z,c66(febGB
&M-;D8\\G?(3F&gU-,J]caWb8XZX8&4;bf)_N##UAJ304=)&bU:CPD/C6R]6V^eM
LfND^I;=&;6+ZVdV:).eDHcKg(V1E/Z5YUWV0]S1;_,SVgY<Z9R6S>A.4KERFg73
\O_e:YPgcG>E_3&+\2D0,(KLFATPd/WJd:a(OUa_IMQU;V[VU8:JQHF8OUA7)TQ#
[eHAd/P)&g?.#RI_CX+=SLAH,V\_VbK&LQ:AHN)IL4fS]>4Q59&0Q=2]>O^B+d5e
F?f]]=e_@:J6bgFcV7WTJP83THEK\1e95V#,4A(aP@:1?32G<L3?^ZL2cAWHMP-+
a@T-f4T22:(>KO<FZIVXMSf<6\67:[FBeDK/#J9/[e5&9]SXF/4BQ3_US6V9/-Z_
T8+H)D6HI,I97<R0EGMM5^(f#SXX_+b<ZG[PY,&S+cDF/-.R,0I[0fcgcV9S+N74
5C22<S,SPDe4><\;B2R\1LIc1/4/_J:W^LP@9,<=Mg_CER#UY+D:;^2&H<M,I4gV
XNVRD<C_8Y1^2PVJ]U9?A>K[J9b&,ME8FG7;7P[.?@E\Oc\g+VQ\4=:RANR3QVa.
4HdO47GFN4([I1+eF5T+@E#FQSGfMbULLgH1]:DO,Z[T&8>?+F7+H7<gOWVd@-C#
-eJ\Pa;/:9(C:[#[WJ_WUB(2JIBfe2DKYG6(g7eRb(Z5GOOG4F7>I,>74E9N3/.]
=ONQ9-@f7_TFC0M;\N1S,]G?JgUX-eL>MWGU2OSE&E<U-H8ZO6Z#-FA>>:V-cB2)
;=F^6-MO&IOYINU_1_A4Agd5:-38a5X/;I@D)NP@V7IO/,I/CBN;>51LYIGf^7X#
EDH=KA-C&Y;L/#4:Ke[EIfL))Q.L>>5T(>?U5@2fgTRF3T?Q>GZ?gKVWW4Q#UJdR
98fbA#4XM;f+<d@ff^4a&XT.&/;SX]7c#O_[<1b(DOcSX91#0=@JE-[S=F^+^B;X
ZIdT?;^>:?5V)(2E1&DGZe?dI18-V97QeMY52K<d>(GL>V.3T)PRf@ee)(XXSJHU
0CVNZFRcE>Ld>YQ><Z<4aC6?UDNL&(R5c,<C,>Bb,S8G,)XT.+N7AK&9cT/I?<5/
d4_OYa+4f2#XYIFV@71R-+e>J_9]9TcN)++a&KA7MEA>F&Z/Z^<eYdEeZ.1d2NC0
<>/Vg_f>+J^.&cWdJ:0I51aHKPfP;;e,<@eZ+N?MS8a.>^gD1DEY<VG6V><-?)eZ
)b<8/R521;dA1>VE3K?VQ/L[f2?Q3YDe>c[(JfZBM>SG]<U@EQKOK8K7PDc:G+c;
>S1?8@_]38QAFH;5HG#QR:ZJC<f-I28=-aD9(SZa=.ReL]EP<gAOS(c_gFN;X5</
=7EF7IQ?/OG;TL&7.F:DAY&b(\ZJQX)G79H.?@:?002;;1a[AcQSBFfg]&6PZLdZ
L-@>V&g844,F;fdKg:UL@PUEc;W+9_5T+OH3OY3)>5IgH4?]=f.)XP]<aZYW@5QX
WFdIQe\<,_K_>WIP8f,H,f;9S\FB=3W)S95aQ3)/_U\5-E:MMc]a^L1ZWWZ_)L54
B8]EeU,f&OOT^:VOU\aY,0(cL&NTWXQFLYHdB8I]bHD@VPQLGd/4gdJ:_]OF:_G)
@MC)LdZ38XG](\H,YA[K7^=,_HgAKKRX]MfSS_/QZ+IL,(.fRP7:gTb)gLG3X[0/
.b&Z:&d_8B#[2LM1L#QP@MB1-7^)<N_=f?/^Sd+gK+:P_@12X#Me0^)?g\G-F7>/
&O9]]0Q,Pe=BP:INPI/1P]YCd^1]a9O3>V3/aUG@PO/0V/)CACc\Bg/3a;RLG][f
L90][(LBR]a,G6>A4f.XB6?3##IIKea_=Of(^?D/>/O-7Z96cgZWXc0ON.JaXg38
AMA0(b,PEM(5L#SD#KL0QB-MG>IO_1@BNN_]7S+9W5T)N46/QW0T8V(K_J?g5A_G
Zg_I?NJTQGd(9,&KaR7RZbTX&,DZf4.X/be?Sf]0Mc6.92@R]a1HC9-f38a&b^W)
B;;_9[4IP<fcVeCPce9621g#^GKSLXNK\eaI3-^)2c#ZQ,?WK3DI6L,IQ&T^KWPB
a>GN/NAgMP->92@LTVMOe[aNB@+BcN=YRB,O#U^H9M[TQ3/2U,25XZ]DW:=[E5)S
TBLFN+N]072OH)-d-f02)?.YYKRIT12g/fM@(6d:Z[V[<.BNO/S42/b9:OeR=VXT
0D:#NVO(AgLRA?bI,YQIQ#ge6F0@Q,+IW[JH_d#Q5@W#+F\ZX>FQTJM&DTP2_:/.
+-TWD(-?,A\0@S,5FJb=GX-?Z-[J[R)6eEgAWQaH^&]7_9I13#89JX^C09JXA&U\
88D9(c/;9M:I-6[-E,@,f,3_[deF9Tc49K#8SNdEYUOXd\A);;UPK0PTf5F5#^Ic
=]D.YeHP=;._:cP-F3>1@I&KMXI@;W)a\=ZNM\0XASf_&I,S/5FgEa?>5L4FeZTK
\[.>R3/e5YOM5[XgULdSOLg.1?4:.:IO5+Z_LF88I.5ddB.g_D[C?e+IS[gU5>gE
O@@d/83T@D/=OT1Q7@T#.&E?P0B4&1FXWc9C1e.cBOEIfT6S.Nf/+]TQ1d+W,U:4
TF?:(R]MU:([IU\+H3@gNGD\7HEB)#fBS1AE8\],fG+dB70bD+QM,g01GQM2K@Tg
_+<[FJ-+5^^F?]]EG9GWY6FJIN6C)[9XUcNEBRb_FaJ\#eL<eA1[6dRT[14,C7O<
HWF2&0WY9P;1ffL;0#g,Vf3(DIP+J]P-bO4B^MR(e[\ALFFgUIc/OfA.2_AV#H##
PgHY@_Z,./UBJ5g,0S/dHaY^8?_8X0;^.56.I/dbeZBReIbPG=#0/7_-6&;2W;XP
)YEJTQI+:(7,JXC&H,0)gK9[(KUA][^W@D1cFHDKDV08+G)GL:]_\0cNM_\3Z8-Z
9G\894KW+5;09=00A/ML&]PV#-EU^J0,HY=;5G<bJG#]YQ8&U^VK:&1eNe#9H2<3
J=:75:NAc2Q;[;W/4&TR4#E>A7PGc..@;PQ)Kc<VS@JKKRK3?KM1,T^c/@#5b^.R
b0B<+9NGKFUfJ+4ZO0eFD:aOB.aM48/PW6K<8I=W:WA+e,X1?52Jd8PH?<B-3>TC
JgRe6BM6I0UINaB#2.G^FYT=0@;>.T=?=(T>[EO;IK=Ma]S>Sc;cIEQOD0GG1A3[
AOJ.&:E96,eSUA?XQ^-]ZO[e\Q;SX4a123QN4FS?+0RV2UE\J_Ua\?HDFT+c(O-J
:0R6.^@0-QL(F)\:MYWcK63JH1@]HIYD+N88#a?b>7b3Hd<SPXK;>/TJ(GWV2:PS
S;7U#,ZWO/B8SX^>fI?EMYARH-7:S6PE=;T(_H-D.K.T:3f3aT5SVQJ,H2J108dB
;gJ=E>;+>W2a6(S2\(@?,gY(#RZLJ-[TSLe[.-e]LAA&DYX]Q93Kc)QV:N:TK56R
/>fP<LSe7WLX5H95NXJecM)+fcd;X8R&7N@0@V1c:3@Y9[eK9S#Cbaa8C:Bg^@f:
9g&gG1F,W=PS/d)UW:RF\RRe/:4VP+SfY[93Bc+K(eZO=CB).E.+-F^=GL2R&,@>
881f5QO-U>ZCN2/?YMUFN_#X.467>b?>V;K>Nb<JDEI+@QT]0U?4Ng<.#5J]G::1
@;B2/bKB=(;=FeM]PIZ?ESGGPUZJ+Zg)H+V4X]c(.3-5Ab>S]<.c.4LRPP()O(07
&#J,)11#bPc:6afFGWWQAa(AJ7Z:eBH6OVKcb5+95G<W.Oa0b,F906I<EXU<RSBO
5_4TGe^fbRdbD\W(,0WT0U\LP6US8>8;D/D_[N?W.a/NZ]\Zc9?9#@&Mb^__5/T&
fJS+#VL#:Gg?XP+e0MPMH1S&3JSNH@HdSbDOZ.TCOK57a=X,cR-MRR@[5a6a2eUX
.<cP(IN2&OQHL?ge,4gTCI-4+7fE&013_+0L)]A1f5eI33,B#\A?NW.?X4[9=T\7
1#BWH<e9G/\^VEBXY^/2EJB_;,@D#2MXa;5]BS[T-gJ+&gL<fYf<A)3;EEN/XF-0
eZJK&g41eCBRg?9M@bB&gFWH+eYFF1)J+I<DGbK9X0W)U-aF.7K9/LV1;9dB3VF/
MUMAKI1AD_3baGOYNNC50\0O>?#-^;#@H.BCJ5NP-Wa3N3I)_O/_#&)T^Xb#\fc,
dFBYK+WQeZ,YSSXPB^Be0DJe2(=<9gZ8e::X9_^/TI1^#cSUSLaZN5b+V1_Q83B-
4MA>\)IUJHP7SO1=R&[K(8YX/Q0/4L-O2&CT.C[I#&d0U:#3Y<XUF:#1((I/.d<K
H3edD_2?K\>NL9#&7<?JI83:^d0O3fSYJQ0NWA:Z1X2IRB[KK#E-[JMRT/861^eI
-JW/I2)RGc6[JKP;g(^FSNce^^<H?Z^1&a[^Y3HCJ::XUV8UA-+42:TLUO8DB]F\
2H+^D]DL]+^X;ZTISc]D-?=LDY=b-Gae(DTc&Pbg4XF&I)HSB>1=2@7Ec6Q,9GMb
gT\8#.X@RHAV#84:R=bED+6,a[\T5N[NM#>SR[1BG8eE_C#3XYRY:F,=S<7<6FPb
1g#=5;TVVU7__]/4M03X8YU0J_AP@EIa?3WZ2>\_#3126;E;\Kd68d-6R1Zc^,(<
><Q8IK?3T?L9B@[VdM&W=:<4J048?Vd)^A:2QJfU6UIX=M<EW>/;(2L-UQEaJAQ)
b[^Q?\-K5\(:L[1S\AV=H6+J,&4f.#C7H3@O3DIN#&c_b^PG+2)aOI/7^K)5ALa]
b-O&YH+I89b?#?f?.BQN6gU,8b#+g54FFc>GY2\&gb6T8+]X2+XH;P[<MWMe.f^e
<L.+D2>5Uabd7cg5C5a]TDbNfWP4[gBX^c3V6B<HP56V@=W[[_dVXJgcW_-TLN:>
M+WY1;e-9O7^#9KZ&-??1OQ4S&\:PK1KMVU=PbLJCa]VRLQbHY5AP7M7-^,:VD9/
QZ@N8=0JXKR]:ff77<:bgTUY)NU+-H.gE1C)cGG^UEc2S<IK88bX3>QdHDd/c.1#
2:S?:Ae_36&RTDFJ[5Kea)T>F\LEc3N?GcLUaMA[)PE:R,YOa4)9#_>L]PWbS/VK
;6V83(RB7BTYSCI4#KD:AH@,]VVX^YVEa3M5#NF9.SMYLB.]<W94OCYR5>76V/,)
Dc^:[8:=f[?8@64F6:O\.0dVY5DgSNHQ&:8d\3)^ALR3)O042GZ2_PZ?7<B8##A]
:a;K5NFKbQF(d#;B9f]52ZFa<L]9:#=LXR7(Y5&M<X<R8E>g7\C</5</4V>9cTJ>
7F2&e9&G?/15dJTJ6U_6aG((f-PbBR/RcW88g?+.Mc&/@O\:(,2DALR:?)AGSTJT
;Z@?WWW#eDOb;W@gZedN.,X2.agda(f1A8M;VC=\W&6QLZd<?3>?]U._ZLJA-ed2
U4RbKbYH0>_b?_-\#M0=UNf7TVb27)AdD+6-0:5aDa3X,f6PU5LBZECb\LC0-:L/
L##/fLab@g_PgYT04\4K(T>6]CWZ/^;5UGRK\BX\gTIE-(K:QZH:=9]N<W&_-ff^
B4fRf@WTH.F_X6:5JA0LSWEBb)&&EULG391JW,0+gCA0(eCL8;,230e)M2B]a6T]
&@>A&.61&R/-7:Kb/7Z^M+/O\D>4Jc&DCB/_#,T)&6I6I#KaaS\Z6B2ONK1XfOL8
RbS>_8F5PGfLV0E(gN6DD.E&&O6M(DA^Y)+aRA6#KcMe]WUPOK8H2J()//3;X(?L
&<g)\DJV=O>.fA/a?)e37[AQ]LbB[0@eZ=H&<[>JU3>1.aX@]R^MDEb:.Oe21<9f
3,J#)a6D:#@P?H56)-9MZY]Q>d&Ec2Q3cXNR=.?gR_LGUJMCZ_E-ZX/J58&\U2/c
#3e,UJfL<7YBcIUAQK7DC8IG@U372dN.MSM(9-=6R^fTUeY.6#AG[]9&R.QS82+1
6W^D0Fe1aGd_74-J.HN45_O)>D_I7gAKbFU2g(A[@#aMLOaD>.]Ed;YfB.YK7(PC
9J5N^S[/5TcC(cBI>)e9TH@29E\Z=bL9OJ2b<.a6+J#/c.Z8,S895WJEO]aMPZWM
cPK_:).L+;K<UE.6Q.D;D:\dI)Y+LYJR_K7VfLM:_1S(FbAYW<>;K4;YI#(f<R-4
cPLNf#I?478XHII_^]NWTIYXU1:PJL/+I,AJbB#AAZC.6=gVgKg8b\@=4=3<LaF;
D6&=1[38bXO^&/0g9Q6Dc:WfNC[HN-/CX0E?eb8T;?=PZ8O\f?F2QC\.6X+:gLV2
47LcLf9FR._)EU,J[WG=OJ91eaB-gF&TXZY@TW<NJWT5D3[PV]H\NW4WXY90;>)N
KB=1P6TNU/GeQS,YdWc1Qb<cO&;FRb2eSGR4Y6#KGRV:,@LQ2ZV);0&NPI_^7adB
IX0H]PC4&2R\e-8^I\K,D.2446)/KZPeL1Ib4UBX29e;GV/X3)(HE6LREVLe9,KE
Kff1P8XbCO5M,4<CLXVN+->TV]3fbZ^eU:=IO_WZ07P?0I)&GJX9Z1E0X(49)W@K
JPX-),B)/Cc5TLcTfH#HMOF],P_g0NQ\LJY8P#:4NF3D&):FHNJa7D_TbSb5XgT?
e7c#b4ccH:0^/OU]g5HCYUQ/Z(e97CRcOSS@7O5E=SV_5DM51\3(1:KeA4Z=Oc=;
e&&.(GaHTJ1c=fcXQ>&f2-@/&2ZWN<;aFG;B/<\<D(:./+^57<V>X#\JI[Kc3SVc
^58Z0/C3G;adM12b\5Y=M=bad65ZJ194M?cUc1;P\WB#^_\8gY&W,aXZ7B_=6=FB
H)[A+EO^f<FE8(K<1M/c>a]8Kff@CU#OECT#&OAO0dLV#Bd)UedHTWe#AU>^.9ae
f;fdOXOa;_Y3/A6(.c8XK9(:TV;H?1/TIMff>DN56_gL4OP3QfVJPe,+OJ=T3L.8
&/-f<3,a_gE@Q2&We\P=;3-3\4-((X&ZST:fbY/8HW^<^3/XXX9,:S)=C4\bI\XB
a6W:e_NVD9NF199X5&agWYOQ6QGA1(?)N:Sa>/+.R0_/Z:W(g,7NAQMCR8\\(R4_
XQ<L-[44eUc)gSQ_=7:C74S6gTQ/Hb\.d^X1N,FUE.S?9=\)T[U[&f.-SD3-P\XK
M-223+@+aXbg#JcVcWdZ=8[-RS(6\KK&8JL\U[6(D;+8AG<4WV(Q:gK>>ZS<>b:J
UD-W4-f4a+c/aX)(OGC_2=AC^I5-fDc0]f9<WTG?<;[>Rb__O/F?7[EP&8aJNZ.8
[.YfH)SDgP=9_/&8IaH_#?HON=5T,0Lb/<M>B6b(4S&]A/^c2\7K=@P\BX+1TFUT
ZWC&aKUdJd7VUOWb.^P?NSTHA(4&\0/QOTG?WP9N<Md2]aHT;e]]EB??W?,K12Og
HDFCY(f<@IRNG72_JBJ\/][VW/>2>2DB<B11Y9L][6]DL)TMM/&4.U)#^PJ4;19f
WPMa,KAb;0-=263BXP0I:RN^6(=?+NHe9IDI9BYZHGGa@F#^)PdWM#\De<AB-Y9F
69<P32XBPV1?(/Z,\1MQ4KB=/WXI?K]+N0?U&<JDUX(OM-0JD3[cBIXX#T+Og/A;
)WV:gBNW?/#&PR\SDM[Q>6;;#<D3V.dXc[=DCU6:f\cU=NF.^SRAM+cG_MM[^JY@
6;@OR@R7K7ec/EN04(DU\dSIfA?3CH7=N+8]E,@f-;,Wf;5ATB_@]62(L6GKA:W9
b(&43R#S^94GY:H@KR72aJ1Y0#DSQf7++QVdCAS/_-C)?D9Dg^R,RDd@\644[JZR
XY@[BeFdEP8,IOWV/P;DcRT2)9a[]=f&9B)de+@UMKR&^:R].ZH,gWd8a[dg+B52
/P97]G\aJXNeE+S\[H7Y@.VONMe2:f(Rd:IOc<8WHME,7=_W)_,WMB=<Rg+(V\X\
MF38-SZ,Z-I/2O8;MSNAcA=/^PMC9J5:O.aJ0RW=Cf6QAL<A[1.PZ<cYCIYUNH7e
[RF?(5/^GUJ8CJD&EAP30..f?)L<&G,9K\,\ABZ[1=e<QOfAH#F6OaMUY)BYJZM6
bNQA)?CaTOF@VbN<1aSI6KS/>#?6EO&277BO29XTK6d&JT^_a&DD)-4?M6gf+JAa
\4F<4)N:AdZ>D6VO8JAHbL>8c]().6H3B1L;0Z)dO)FPAfb,4_C?:>)8gI79aLL)
.Q_FH_DHTY_JM\F):2K-9:;7\W4]/^L1<?PGgP\=/CLI?&O-?YS1<GM#7bb?TM7B
=4NNN/X<]g;D8&&B5d#cCER8WcSV2;CN;Fca]I;E+H?Ed-YRLC=\L/LWI2L6\;7.
2;#@Kg?eFXK0;ae/C_;D&_LO9@E>GSG_WC78D23)-#&SV.RB,0Me0f:)/:e>9HeI
c28fBH<1I[^W#:#5H6[O0/ag,9Je)e>>d7J)<Yae34dKB_,ACP:3.R-W#f\R:g9B
C1KZ=JJU6=];cQ:Bc08W,MT3AD[H6=EKVP]RBS;?Zf>M70>^EZ=_=bS\O6S.:fQ]
^.e68:a;-B.0:K<1A9Q\O><#b>BOI,Q6]]R8[ZAN&\FB8MU>YZAcX[&7aQ>.P>2S
9PW?3]2ee;Kb]C3CF_^NbG@(+f^U+JUb-M:?VE,=>,SE&L&e.Q[D>TYX;S#W=G[b
FbPbWY],M)W&@T]V.3]IM\dU(=](g+A2/7000RKeZB1T7?e-+VS)4&ES2RF&fLd,
)@4RCIF_:KJ1QO.API/CKGFF0,T#0:T[(O-dQW[B+Qe:Y;]7M5.UC=4L)^^S8Z.@
PT4/aIR2D9ZX<0RbTbW(O#K7d9U8>>a<XSDD@[8d46e[:DYA/ceO=4TA\6SX7RfC
BFYL;O8JOUTO?M_.J#eS,;6?_PM4TMB)G;YIV8_04gSCb\T8NA&UfPT2><N(:M96
ZJ2-A<@6^Z?[Q^2ZB4H)AX::=].?[C06AYYCW/GEBHI<3.)E(#X@:D[8fG)[<Nf+
aINf]V#W2gd@f4b9D>-NJBD_P&C/GP9c^#]Dg0GW.5bNDP#g0PdB[C&R2OWU9X:D
NCY;8FB>F06e3;-_WbAO-^,Ee^TQ6b?K==KG(J9K0B?XKY?REK7#OZNe8A3><T\]
.c,S4[+FE]dPHb^T<LR-g,1TMO@E/0/-6+d6d^D8AFU)G=L=8:bTI==ZXS,Za3Rc
UP23UP=2Eg-McHB,GWW6bF=W)9CcMeCJ>dEJH5HUS9JgVOJ;MF/+D78A54<;ZURP
HVfH4UTAQP4]NZCJ>X#I=XaXN1=>RfDF?Y7B1B[S+ed83bIHC7YS8^6RT->LY=ON
^bYCT;PW981-6ZQ\dAg/B[Y)Qf\^LV2/[X-T?Vg+?+gZ5KVOG=LG+#e^f7c[\G6Y
(MD=(\++33BbILX(&\YVW)LbU0W^-,A>DTJc0f0VL>E1UAK.^8TK>+GXF]C0/I@X
))67Ce3K/(/(^DY([8.N@Fb)_>.I3dG?VQSVV)(fFW7\[)(a]S5[SC-V(1F.I#cD
cSbM9QZ@)WQKdI7SI&f8@aA(>8SIF^7(?,5,CgbWUN2;&\H_gXKO7c15d/TUF1&e
KM2MW:]f;41:a.R73LF<.ZLd(DLW&WJ7de4e;&aG#C;2LQ+cENaGcH<d1G84A;Ia
+Q[,FQMAdaS8Dd/U()U?J:C(QKPUT0G78]]+^D7f13=<+-c@eC2GZ,3K61a92(8W
1789C3]&dE4J51ZIf2-B9H^[fJS6AYR#gP,V,MATV+HW&D<VUT,7XEK2GbKAcETe
2RW4U?3W)gaWJg+B2#6.],GP=Q=(<J2d7G7^7C7>-6B)8QO_&2R,AcebgGfP5+U,
77?Z_e3)@d:.Z0:Lb2^?ILETK]P(VOeH9\c+Ge]g7XJ:?S./Ic1,JYCR,8K4HBZ1
O8?WbEWPS5SE87DO@V<1#^.aOeN=aJC(]1^?(#f>S1<L_P^eV<F<=;NOKZN]g50L
D8[T-+GGX-=Oe91.H4JfG?^a&5F4/+L>67HHLOJg:M,W\IWVV33@]A@E[)?KV9#4
ISY,Ec,Y2KbRef#KBd(U?VQE&>ePLPE5S29R_&(31]MMaf@S^L>6V;R,^):E3@\T
7YZ4)NI&^>@2]+(F[X>(aaW:S@(I([6H3Fc,8X41@cH/.B50>K[/GPA,CTKNKGRL
2]-G/<XI&Z67f@VR>dL^_7(2,R8Q+7&)9^/.21-I15O,6\M=L5:_@QLd,4OHBYO8
]9S_a0c2(/ELV-=J^:,RR[S8A5)<T&Qf;;LGWgE.YB=\fS.R745Y\5Z)aS+TBVU7
](VS_?bR\#[TUGEX9+Z7g>9HIRJ8FM5T&HR:;MANM)&C#0ZRY_(A<(RePOL6ZDdc
NDAUT]a&TV3[VX;1-C4C=IgLS8.CC(.GYF:AO6e@9H&0TQE5fP.eG-E>V#ZPJGYS
R-72BHeQQW2NVcD7b)1<?90M;VF+3Z9\>G@9O]#N;^;#\f;g@\?X\IF1)Z(A6BG;
1[7WQZL_/g5Q0+E.a<V#XJWg&,R_[DX\/Z[P97>fN[8UaF5d0QHHJSCaY@A10e\:
bBA@ef,BCGI>.(],&7.@^]R[3HaB<eQ[43ZF>d>,7>aK(->QMbXK\aO1Lg7CIM@H
^c(7B+/C=2@]eY&\)V1G^J\IBb-7XS<@N:Tg2YVf#7QeA0]2;b95L12<_@(.C[?;
56=c#=eE:f[\VI>9?(]2##5O5KRMf=cR>MVbL-Ha)0?D<cS[FQV)AVNS6R]JX>(I
af9#U1;c-MBYbNf2RcOZ>f?;#X[<:V;]Hb_L/7YGg6\9A5X4RQK5M_Tf-Jc<@1YN
P=-C=#&HeK)1.#=T5X2cG0:]5Zb7#.&Q0,Gc=KS#^gZN:Cc[Vg&LDf9<:^J7FS.:
>P5)07Qb:YJV862TCO\>OP1KK8Mc9VL\=5WBVHZIf>YIJA?];;TbST@b7ce)J@\e
G4;YZ9]MVg(KK5[Kg\^M5\1:8W2#\.X:O9Fc(ML(^+.X(gdI190^<P=0EA8>:L,)
>JRO0+aU:<HF)KC]P^^aZIL]U1b,A0[7[YeBe\R6VJgW&7cf>H^?2e)NeHAT^6EO
Y4I6?MX[&OLfcGSZe/DG3ETbK?FSB.C[a-2Wa,O+bT.H^cM,MW7)ZCd4(P0/^VfJ
YYTCNKU2_=T;,0g?)Kcb8CI[+dd/.,e;N^7-([1EPd\M;--E^Y,gH]P\K_7a^gWb
:bW4A]><PVSIXTQFU=0=;<eQ1deX?0W.2WKB@4H6g,/I(&:I=94^adW)6@&)N,=A
E2K>G<4Cd.)@cI]gL,MBRSJ:?f0O6<8g:QgVT,NHF5C2^)_&J)-f7EC:\dLa[.)&
=Z>\VeDZ@d5<(55Q)T[>K.XQ.+_U<-]O)DId+YU;/RD]E2g\MB\NR#S.Q4Eg0RQ&
2;PHJ/G_1dVK5>:W6X)e8(HZ1dW/+,1cfVa_8Q\^+74Q+,VODdGFLIc==QC9N.L[
IB-CI#BEf2BRMZ>06?A4YAbea:;4G(@@&@a29G(.a<?@DR23SPX_:[2HJ8EM5822
S9dGG+Tb726+Z#3TTO-;=Q+_S0ODQC=gT1I26LXdeSB2U]MRY[0DRXF7\NU,.fGa
C\R@M:(.7;,,7Yg(=S-KR4)?8\V^#^>8OFUe1&Kb,W:_-]O0]FV3(HcScH>bFV0H
Q(>PL\_FVI[5=D&1<(eEa9(D7fE98=<+XL[?W;c9L<OKA86d&MdZ_AV?gE9c>UMf
[e6H6OaA5ZL<cFb>42TB:&4@G=\]ZS)8f]Oe9dJS(CV^0^SL29O5bcFJC8U>UMTS
HT8TN#K/Qc-f=5U>MbS(;T)BQP6-a3cLAB2SO[LD(;/Pee7IC:E<(F:__Wc7VgWa
BP=>33F8e3V4#U7E9>./]f\;S#\AeDGDJgE:[1P4,\4U[.N<C<7a@42b3Ud.cF5G
AD9[G>BECOUXRbJ^/(0fTE4&@9B&LAGg7;HY7Y1MaD-\[1/)dKHdbO1.;T6f]EW(
K6^-EN5V,44MVI:I-9BC//[+Cd]#8d^dJ-D)@UPR8fc0>[P)850ZQ,978\Qc>R&\
+W=K614R:>b;7-78=]WD.WJ)d=9LR5MN^ZYdP)3L;&<6gHMF<;K[YXd;V(JXGIT>
NCO8CSBR]&Q)@P\J6)=])R2WZ+6:>1>g>,X4EbU6:M7&N^RWb1QQE_:-<=K6aDLD
/T\L/GRZ7J(Z0ECea_d5eeE_d6.#D^6ZRV.FGT2-ORIM_RX,TG1PSQ5gDPg#CM<W
3TTSTO]1ZV)E0LIS@[;MXd&W9BC-0GH9HDP:D]D2.>gH-9VX,a9IMYCac5RZI=JM
)4MgP&N-MW<B&4@:E.1f=U=&=1@Sg.aE;/,Q=&;EM&QMJ5BR5PAcHJDZN]A[&Xb)
#,&.4g0Y_YU]6f8<41XSBK=2KA&d5)O\/c(0DHcbQJ.BE8RZKcB\fI^#NAbAePBU
2aLD\1<QWNaXb?](1NW6((R-WLA42-FJD3]ARE=Lc]/-(^7/V6C#;KUL-LQ=,VfB
>MK.&U=]/:GCdCg(;]G#.X1Of0f10LHc.]6Z4)JYJA-;gAZffFX#QG9/gU-OQGG\
PR,V+#8&5[#ACBQ5DQ9_RcF;<?cd+U.=.;=c0L<SHW9?OV4HeZYDdE?(_?57b3T>
YC#2a).B_M(K9EgIbR#&68>9P?54Y_W+>.Wd-S8:6O:9EBI(RNe:WZ1;WRP:AEK8
Y?[0W1BOW]AfPD2P-.7ab9TLH-NgK3KcAY\MgaH<>gM\aAdF^0S4XdNDcdTKZP/=
52AXMRgD[V]2R)Uc?2Y?.M0WEUCTJ,0Mc):T;)f283T9[?CLN>J4IA5)Qg@g=6JL
/<I,bGZE(IAG/.:H7RMB?Bd511;\BBaI.CV])5K2I7_?4;1A:<Q3QC=Ga\PdN1L<
211#;L;dQN84FGGcR[;c@,#a+A(RR,bE[\S1LJbc.Fd5P[3#]13g97M4/K@LdIC9
H,eHR#[LWH()++3D8/&;&,-7H7aL<He\\6CgP>eg&&c=^D3.K4A3.ZG=N50EGJ,-
,)YF<<B<>aHVDFC)dE?d6/dg:bB]W5T)Hba9:c9G9>^)Oe0)=0=dA4V.#X^cRY91
Z,L)4CX]KD2fD&1Dc^fd^&f/L5&cIKE^?f#__IaZ+7GL_-^/Z)@^KTU=7MGTKTA5
N3KM?@WQ^+<?Y5eEU9\V)cNIaJFF\V[bZWNT=[+5>>+b&8EPS?,d1ITX]654\.L)
=,N)D0L<[.X)MXc_=1G6C<,A.F.BRQ,(:#9E\:[M+0NaS1.4(ZB)gE\GYXeDM)2M
<:aR3MEX)KD<SV^H#7K=E;JXUg:X]G[T<N.16\4@4b:-.bOBg3INI&)R[c?eF7C^
2H5Ob(K5L,.YRRTGfB_[aP.]FI75_-#T#)-826MZ);C0Bc6IgSc9f^,U^/YA0>G;
(3Mb0;7H>6T/Kd76V3?<B0]I_OPQAY2aC>1</C(b83N)Y94?)60QN33.Q]XXZX?Q
f__GZ2H-H2_?5-B6?)K=R1/<LWG5]#):=BU7,VN&IYC[:3AP6TEM=TWf4a]-^5YI
T4cB:-_&Q=QI.B@J.;9H>L>_]QA2YZZ:6(R.S_7A8ISR[;(De/)>?S[.__eUAPI9
HQc3WLf6eb85X.[@-LT6_a9H;#2B?\91@7G(a5^,[DFZX6E3\T7?4\4TYN8OfRV2
79eHSe>d9[]AQW.E:f7];DW]><6JWMc5_ZOWL_;??#L6A+<e@N#&#E6K#3]#6K0b
L^]=BK2AJ6b/cFRI.L<g347A>A/@8CVZH2c]-?cbNTW;B#<BSDN\_K.HA7\WV[]L
KW1@DX/&B1HJUDc[6.(cTd)2+Z.QY<f6]e[?X[72d)3c[:\>_a2LZC\1+8C>]bCG
Td,c=9\Ud>0Z+PBZ4U)9b_;N.5+BJ.;:a9&W.M^3(8Q0H^EK^BYQTM]8c_JN,\D_
B4^/==X6D7Bb3@+AA.E<5[fT+O=5]DIYAIca5NQ\QgDVC4[aGaF@\7e\:WI>/JFL
:(<P.#c-fRI[0JO01C^YULEC<B8ge&H()<aZ_5@=+_eGY+F</G22a],(HG+eX8N/
I&O<AKQ[CXA:S=g]>dKfF()[Z9If-(dRJ,)2@Z()b@AMI)#434g?&=f_93#]NV23
8Gg?aU23Abe.c4[WU[IH_5>U?S2g,C\Z+(DP3Y)>M+[KOE1IQ8)S,g,#3aKN>?A9
E>Dcd=Jg[];c\1.FB5-W.,72B\?12g:<,EJ30eIJ4fBRBH8N^-bAP,7a/:Re>=^O
X5OS12_Y5@aTPGaLY&E6LOQMYYFP-2bY)HZe?dPGKT5UKH;AbQ[YL4-1B4Sb4\A9
^KRgCFM5QFXXC3c76Q:J1ZYVJH0Ca<<G&OD:04XB([@B;GC;9([^b2egK+7c7(+5
NK-C)5:gbLK:W(Wg=cSY9(PL?;<[&QZ>@bSeWMb?VWL3:eT38_G:10VD:BOORVM_
WO\6V<,gS.&JWAWV-2N)C2V3E0#e&.N#(H-/cMN.O&GfYWEO[W@LQ#3(1)6>4^Rd
^gAbRFRYNY^<<I^g0(0IIDW65L(=^YgLF4=ZX&-J2[N=MCJ3?0B8_A]YF.(8e+AC
eSDWP;U#KT&_\\Y-B[J4UVWUS6P<T2SX(ECF/;H:8666/MA+7AP=-6c7&Q)Gc4M,
QS(@Y81ddCE48.\7+K=W3W\PB@A,a4QEL,\e_F3QeST:_.\gPY97W4cHa22@J\a0
&,9BD1;GCW3Y>XM#0+P_:7fMA.B]:01-1eJEA8<=6&ZOZA04:8Q#6XNCe2cdA6QR
#11MWDE\S=)<]:14ZQZ+8[K>6TLHYU0#<g_1J57SaV\>1JR(5d>>AJaYcgVE.F6=
QB9CIZLN1.eg((:@)DG)fS4OLS[S25SY;^\)-4-Ja1.PYcCJ&&(-/^Z<c6cXTGO0
47-4JD49.H.R^=:KPP9@71)QgQ6a4_39^BVKV/LJVC]MeVESA+;I1X@8b1O^X35N
0c@;dN::O)C5Z#ACN1GW0J7\[@0SL7#7/8--[-g>f<80,<[X#eU]-c.>2LeA/)ZB
LbT3289-(NgJcdHO+CZUU12;;J0C.]]B39/2X#U78f0W(YX)N/Gd\1&-f+gc#T?F
EQb@c2E+=eM/LH-KXJSK1FOJP^R[?5IW]\gDW)@BLOFbUZ.DBSbKD]_6N&CV@?-<
>+33WD\M9B9#<&E[/\,VIgU-LKf<;&)BS&dd4c&DFG.\G&aA7[S)_4ZS7N0\&:a3
McQPXc:N\-dLEae\D-eT0;;CYP2(N9ZJ;:c-49PXU.<[IC-RR0_(e0W(X3OSO9+-
G#&-@CZDW9,+YYWN6BV_=ZSU)NT]R0C.\Uc4+F&W(>G6gIS.RX7Nf6fY)UW9/2QY
fWD,9T+1^[7>[cHKU3=IAVCEYLAY:IPIV;&5O5(L9-ZBHQeC&QCO#b^83IXe@QLE
EA(a4-22>D2TL&UK_,]g&/CNTL<eRYVMN0R#225^#@H,PG#W9Z>KbXAD^+dWV1W/
g=eF&DDBWA-ZGS,HNGXU82KNeVX<XYSJFA_daHPM2Y8gcNDOX85I8aP44F9GNY@@
=,\<?G)KKFXd=A.3=3K\^6/1\#(M;:(B6OX<HafO:.;aC4L_3?_0a7XZ3=?XP.-f
[B5,S\f-,F=?.g@,fBTI><XQfd/&V9:/?a32?ZUd5GPW90C\+cK)MfV:#?c39^/I
EJ0W,937d>N<g,VA^IB7Wada>II[7fd52TWE3&4]8ZMH-A4Ma:=_ZHW[M;SLQSYT
\69<(8L.@?/DOIK<<<,ECS)1[OSD6R/1DEWYdd?G5Cg:UW[Pb=(,e6;XFAEAKP4=
/T30_+_gCHUSP[ZR7BCK:3BHO/^TcZHQ/,CNGKONCE)UOU?fDWbSfcYfA;K2aCX1
Hfe/g+GVHYfAY9aA#T,:1:/cI,]0+Q>4gBJQdEgJ79e#DA&d1=[_I+G:MCCeGeIS
-H(gEgIR_a&YgYTD:;H)2MM(3d?<CV<?X)R@=0_\]gPee[2R@PK/2E_\TE2)D<gV
#;V;3BX-O;[<CGL(+Wc0UG-AD2#LBe3AE[N47AU_Q,<86cAf;1AB?)7D4L@S6&b]
_5X+<IB8CXO35c)(cgd;7e(+cW7?<:[_da]@dBBDK3/Z-e>H<KF)#WOOX2M<W+g9
?1U/fa&50MQMO764VK?V([d:JTW+H.41\)D.Y75V-bO<@e?XYe2JE\]JgD_WD?)U
>Ke0WZVAP(&5Zg.A-9Q)/N,FN.d\,\HM4cK3L,T05Sf/_NA5A6TM7KL;,YK,:2H9
.2#P^8&V[K87#3L&2RS[:@QT06gAZ\PFM.KB8,b:XbN(<#.E:1(a5H_DcMC)0;SN
MLE]QSXc<-U:UI0KM8,E82<.3][C+SS1XfT:;Te0e6AM@>#_-QEG/7\#D(MU6:E?
<b]@Z/f<JB2PTM;I>3@8U32\IDP5#fD,Q]_3ZIM4AZ#Z63U9@JG[<<ME7^::2(WX
ZQC/<Q4[I(IPS)Bc6\=S\D/8[Bbd(^[P5G^76A/-&H3>g@bQ:dO#)(TQYJ3b-6PN
U^T5\1\7f.2[<cUa\(+<eG?Ef]&:]^JL&E1cC+LY;e>MC,+X8M,96[((J3#c?B@d
QBK&5HL\ZN077F>5MH/#]0@6HN7DA&67]3:T&4=B0)IQ6:M29(]L1DFfLM&D1LVA
:eKb#J4<F]6[<g-d@_.fJ[&X45PGODJY3\TdU?Z,3\B8MYScYb0ZUfIRK5MW<a-\
O+Za^F,GX^MY^2LCM0<NcgW)V4>U(=IT@Q(807W2PUIf)>5GdY?U\+/TKab?5a&Y
6d<#HRZ6Y4:YIe6&aA<]LQ+@38L[e^0\]=@@G>5AD]MP\_@aM=a5abc<=\<NTffc
OVDT7Ve(8,DP32gWNKHN91WHccUd07+YZ-,#\G:ZO9[0#@WSS:+UE3E+2+1^SCVB
::&&MSB.#@G5^aL;C=96>[)HaMY7F3RP4O<W=-P^\UP^&SegYLANV;afg@<P8-15
AY1d=f&ITA@a3B4>:8GV>6=6)YR)Q;N:C&R093YC0MK/L1=Oa59/e:Pe?\->PY)V
gg_-2\RRKUR>VHP:;&P6/#fX=bJ^-BRE_>@gJgS-P:VbQ;\OB]8_=fJ_QC]#,HVV
MO@6:,Qf\deHQ/UMOXJCS=7K&DX4^QD>SS9BAA3))H.O>[dF=A=QT;@^G+DDa1Zc
>Z64<;dL5/1AefG3[G0EbddACB]>2?)ZeQ@2Ib]c24+EN,Yb+1P7PEV>dDGTdMUS
d;)625[/;@aDM1P?d[&18>A9dLXUb@/acS(>g/a)8(BA(79Qd5-?a6HA2>EBLGVD
;GHEHN]-g6_e6W\&?8AHR+N6gD.6AfT7&aW5]Yg#YdW61ga4VERZE_ZLW-.QXLfB
KaSAHJMLP9=;^.W]bRd7,]]_=B:E0ED@BC3FFSW^a1D6c\&L:8\R6L,]^4W<NJ:1
7&YY_L3NJ[>04J9R756P31\=(Q+&LZ/LINP6CFQ,8I\#(^D=&F]6a00-2=TR1WL2
[:QGEDGbN-OAC8_.\.U6Yg+FVg?S[@,^NP3;f4BEQ6W9;CQC3Z?ZU\>NQW#(8:g+
_d>#IQ.cFV:+8KVO2g)7TfG0KZ53\IZ97/F5W_bFW3@]/ZIU6)4G5(.Q)WH3&.W&
RBJ+[d8Y1ULW:;EV,36BW^,6S(dJ<Yg(\>;K4Ia:GC=NQ]C?7I6_A;dc<\&<C:6C
@Tbg@>cK7:Z-519@c:?/:+^VeD-VJKV^&N[fMFN\HaV=e7A7_VSNQ+BRbP.H/Lab
/:d5.H_?EGZG15[Vb+-#GX2NADV4KN<&7QAH>V>LadC92IRc+7WG&1K^^5KdQJ]D
aU:9(d@P@Vf:HJ/Qaf8V+N?3bRYXUQHQUJfV.Tc:e4[V47L1?5&AaW1?5f;FE4LO
Z=WBAZ_A#=E@@J8.\L.T4a.U\Y34dDJ>VSVfeQ-bcU\T<\Y&TfPF:+Q,&LQDPGY5
#;@ZC>^Na/0Z,(8[)fJ<KA56F:\H;=a7//[-4?^g6TH?aLSFPL\3SA:@R\Yc\S^E
Y@Z<Ie-+>d#-I_.K([[#&U->?9e:&RO=[G9#fC7a^]V4g0;QNBT/H(A]FT09FC_Y
F3[KS00d3/]YO2<RWg9EbPT3cX3bFJY0RJ/fcG,eVR/6D2?\bagK0K0_>KB(185d
IaKCAbNKeOM&.F-]Q6DIWab42&_?bJRK4H#VE#Q8P_RdKL?6<PFORS\ZLI@-#,L#
-^CV+Fb@>AHB+\P=?@<\fE7W:Z??:OX<(SMQYfPE0T^#]Kg1Td,?-YTH-J=GW624
3dfSb262XNW1+aV<[F8&K5(W;A(0G4-/FS8)Xd6Q9H89?\;C^d_^MJ20H2&-cCe&
.99(Z2SPBKH5NQ@HIONM[TR<_IIaD#;QVd7Yg#0)B\b09a-GLM5/3G5W@SPPG[-<
C>:@>-Bg:F4-G9d)/=S4RGLb8=Idd@R=Y4bDM,IBH4I[7,=)NH[]BP1-eOP6cS6A
6(.JGF.K1R^01T\?D>-?F+R01g;HMPMGMLF&3U-a-\GAHPWfdX2(7O#1Cg.>FE]W
<E\/GA4gP@#Xa,e;^L;gU7FO]LZKHW/G?S757L4SD<-,GT^IQagM79[44H:<YLgg
X_\e6QQD9g?1[YV9?U7;<&Da7T&N6/X]&(IDdE9A_+KJL?YKeL809W-dH]_#NK:O
1CS^V5Y7;X-M#<a2<c#_9RRLD;:GZ<:+6T^O[Y.9+-eec;==9cGPGA-AY4c?LDI_
LMD?ab4@./O,Q3R3;a8M638)3I^NMbX:PMN.JMZ-#_590S#U0W=]58ONS._5&S;B
;J\2)6@?+&c)0,.&0_Tf&0dB#5/ZgKAD0J8/3VgMUO&QR@X/K/KeZ=dMdTI3JT:b
I^:?e>C=FEVMHS#/gP?07)1\?J?E>:\Y62](7WGWgQYD=L(&B+EGV+THT]d@6T2;
/aX9=P=:M\gFf\9#-9<I\#^OKW_,N.AIeZE:fK=cH]e?:MLgXUQ1:4cf,YG_>3Ta
BCGDBR<K(<^^O@6;F3CJZERcYAS#3V8:7VJQ36:b4:9XTVN0/+b]&?Y-25fZ#8M5
LT-4QS1E)-H]bG@A/I6cG8^WAHcT/(MP,.GIF-0d-,I1Z=&8.BIQ3)9-g0#6:LG\
CgMY@9D^[/#M&F_a/&Tg#bbe7&^CKb3YIMBVUQ?#DVNX=5.K<38.&-GH<+0/]D7@
/f,?6U-gGN;.MD#OR7US-,=-5Of(JUL7ef1?QVN+;O3b;UU=/,cK<EHfA2Ad&90?
WM_:/9HV2I@UP;B[YUZW(Z+[HS+]bYBRA29\E1@dZ29\TD@+/=]^W1NO-P;+WFZ6
JaK7XdE,_,.7+9^#VgTB&&Mg-\=YYG&N-U@FJc];\0P:[)4&D)UX5f/H\Q#.04PS
<2-gHT#5CCM]NLSX7MYb#AcH(@2REU=abC4_(b7ICL/OX6:1eM=Y&<><X8,X0gPW
?W8HGe,OTe7G@P^dT:P5fDZQ=,>/^AY4^]GCU0\A[(P+84OH)RDa#M.0+J)WY3fD
MD^Ib>#[WRNW98.-<<XA6]E?[Q=0e+.N)_a)URM3fV3Q20X<e]bd(@U2-@1Hf;Z(
Ad/&0H7gJ-8C782ASL<@?1B/1.Y.(_-&6:469ZbI;FNITQ@65E81F0#fEVGc.,bB
R?C1C8dW)3^/.CT9WYT>?-\bNdA=dW_(L^QVWR>?[X?7SV)X]dAc?2+Ie31@VZeD
^IDQ.MS+N>/3N3+QG(]_HcIa9(RFMab5Y+GB0=+TW]Vc;1f]b.PLgN.7WM5]VfW&
45?4&=>CQ<LG>aW(\0&^^?AWA<Ga0f1(3+>O;(RFP,bQY(\M]R@6(6C9>:4IfafR
6\GC;DUMSUS)?(^ePG=Z2#O359;4;\QIU^4)2F<CF:80EOI(8F@5C,(T:Gd-;L;?
eU6eR(=?UbD^X69A4V8ZdQ\U.c:cUEOcJ2c8LH&[c<-U1JAbLPY3<<BXUK&7E5-b
J/bG>DQJ,(;Ga^?OX_F:^2UMBI7KO:e;M=;R-,_(b=&K<4YMb+4#C6IeAXIG)N:0
d3#Z8D]XWQ0-GJ9JPVM-c[].O.J7P;c1TD3K^J\.[W8/Yd0--,407<?.(<gI_&-R
VdCD?ADaIS:S_,Ed/K-KAZ@)SM,1bDRL+e-<;M02TBXeT3FCb;g-L_E,Q&L]8N^.
IS2b6HLWP^A/#8GK2aSYbIW.._;?g9F4SK_dN86R[Y;&=f?EX1>W[\RRAA8ddTT.
.&-(WD>S-@ZeB87f/cNaRZAT=;Ud/)BeBPf:5^GNRVK2NG?RffX3HSY90NDL98S@
fTB5/B\^R><W?)[<acdVDKX0B1__\/(&VZ<Z?R7-8)?1aI^GKcDc])XHdVL?FG/Z
_;;[GHL+b-8DFf4&UU9gXRC,^a^WNU0^WUL&WT-IRHWc8ad.UIAg>KdI8#H,5gW[
8+B3OWJ:Wf#P9I+SIYH][S7^2>1287&)gaX9KM8+8:;T3.aQN7>bN(YUV=c4RYU@
&N&4ZW?PTCG^d:>OfE-_6KO=ZF5@a[X()g?]Q^D<g]1d>_a>Gg&O3TdaUY11ZL,S
ACE,0-T^?-J:[14=Q/?DIf?]&QEU=(?D(eSCgD=2LA,]4NVQZf[DP0@T48]8P2a-
ZQFOa8g?RF2H]7?9]9S=0G1TTZUaOPT=&O_=Ka9P7++K[:O8L?@823M)&-FML6)5
/1U#DTId\CYTNIgA;(TJ)cPc?#8;<=8g5:-K)dMB_bPCc\OA]N^ba07R6ILE:,1f
4/bKQD#P_:J30Uc<SdO;,P6X.3WWY;E5_KGDEWKI+bX^N02^=1WTeTK8E4TO&F]&
P[@cW:;4FW0bA.LBX715RX?<_YFE;(W=(bV4FgaH.L&Z1#-<&BI/g),9AXc&(2UM
66QF_2>7A<d<#g@0:B_\TK#P&d&@Q7UYD^_^:-g-0.Qc\ACO;5b0bRSQF7.OQ5<E
=X/2\7dS_edf>HG1a:IeSJf?]C/UPHVf.cKaV0EZCSBVE=c8(ZXBSR[S^K9eG2QA
729;Z_YNV#,fVS7_fSdbeA3A&?0dNKM;JRS^)Q+],=;?9)d9EeCQ8(,J054^2+1D
LWEO8EOT>5M/8GMX3:BK](A=Zf&[aPR&Ld],Da@,9B\IGOX0^TJ,6fDC^5[;8ILY
098TJLL<2KIF>8<Ra0)Ue3R^WA&/e>Y/S(,X/T9R/HBF?ZGCW9A0b3A-+DYVE\dD
H7ag4VCUCG+K;#@4Sf8H^f3S.L26dWdYWRag0P1M=Z<IIM;N1TRO97.f[ZM]IDc\
3DU:CCR:7E>461+3[U4.390UAN00HLeE&NV@Pd^>?:8/5b?H6A.LP5O7c5T3UA@X
BY;5J&f)fZ8:Cc)B7aR+):KT#;_CKg\[LSYbOR(ae?K;W3,bQ[F9\:5[bW8EG><\
&9B1>J_Ie.30/IQB>BeIJKF82bKa<TWQ=eXd,W@aFB[RYWUegK=G\YG^C/TNQVa#
<Vf<BN_\7H[OL-)Uf\fA/FTI/dH58&B0>Cc3-3@e4,>/fUK+IMdGVQ&&F<D]LZa;
=8GO(7.?20WU=>J]2AbUef(7YMcDQA_@K,?Y[,]Z37),SGZL@N-H1aLMNQXYH_d-
BNB(5]K:]/)R(aF][N086@0<4dab)@DJc6KfU&Z&:_?EZKTCCK5,Zbg#Vg@Q;YN,
XJ4XN_=WdM/8KH8^\dG^,V@f-AB-MgH=a/]).HR:-EXOVZ>9TR2X4?6OD-9XEcDO
1SaDJ,-X4cdDdKDe;d6<5DYW7)T>BXc1(Wcg:V3)f5d4^K,EJ],C3QgT[L:RU\FA
BABLJ/-PDg8VWMSGZG/I+d0Y[8RY^MO+U]V2BH;Q#)@Z]0Q/3C.OQQ&gYYG8N134
CgM0GMaRQES13/LdA:#R+I,/^0KA_7LAL[X)X^@U;HV+3=U6df^7]XK-45dfU+L8
e0bROPU&:Of:3]C7JeK/34PESc_O#9W&8#-.2F7@dcc4b_eYWbN8N_JIdGB37Z0>
fCccHG1B9-GB79LKUfTc1M4);P\75@(Y=D/Fc[-(-VUgg;#?V1W,0K;PBX:DDT#c
dXE+99;JRM_21?ER2OL]McG),;]DaDYdB/IGdPSQ2FfR0[)KS96HCT9c?cH^)>OC
4PJ^P=L5c+P^4#EGb/_2]FF5Q1=T7+e50D[,LGE\/[.3:J\5C&Y.Z,^KdHV5M6RH
5dL]IGB24;XAE7:DLE2LHYWJH0?:I/R>g1<&-bMXIgBDca@,=F=C?3C;J,0W@9CU
cT,)gTOR#\R[0/:2DD>N#;HcBPVMdQK5YGZ@RGK9_Z>YPQ<4/0X_#f-fLgEE7gI?
#-;.G^R@\eNdB?.#(?M1;>?,4V>LXX[e/.;PJ(=N+0THYKBc<JEH?>-KW><5MKJL
;NEVO(-G+8K6H0:1+O;(GO:KeUc:&1:GIaeK8Cf<&O/EMG3YYL+]9IGB=65YEU;1
ZX\Db,H[/RF@4DHQFW:;2Q2e)GJA#=(dARf=0Fa]86&fL/g:F4/_NJ7#3WD]UJ/A
;MN6,U]+CZP3?.+__K608D&R=-V)bc&f](@/g0>03Q#TK0e5-631+XWTK;O=G)B+
g-We)D4B6FI/a[A=B#?bN8I//#;eK+a3D0.8+,a5:gLFH3Q^aMZ6)]OG-VN8IdLf
)LK3JaNN^(HS(H=5ecC9Y,W;.CMOIL(=GP=6X,8RV@#1O3Ye9LJB^ZQ\:=4^T++F
PB;[>QFR#G7>>(R[bP_5Y#XSQ3N[\T7#64a(B6QPH,TL]7Y=R^^-CfEJ&Q.BUcbG
;SJc^DKQMQ^TGJ?9K2MdaASE5U\@^.^e]<LJ8L+8#M078[dE#3KX67SXM\XAOd&?
Ae8_\Y:LSHNI/7^9O#fUTS?eT(;B)X;7^dCY+,STA+Y3Q39T;2/?)c.fP<McO;0&
3O\QK^T(9bZMQ+RAY\/_f-]^U-S_]a1#c<_I9c;>B^;V[LK\U,/;dagF<:P_2^4X
7/;7Z0RL<F&.HA+[#ND,.c@WLdYNYS+:9KMSA()_D<T8MWG=d\);?S_\3]_YeKPZ
(RU153:R&9N@[;g\V8g2>B\YVI/D[<-44]R-M>;C3F6-g2EV&Y1R877a0:=WZ&>a
>+R-G5_Y<=D1_V>)YHeaefQL_.gPY2-/>_/\[cX9V.^<Q/P2Y2Y/de-Q46)9S/T3
X4MT\S8CYf:;NI,DG@B#S]DDgMB;IdMM6gG66.V62<KSUY.F1XD;<)f>D/>2H]W4
K??Tc<V@3&gCHdAff8:T8^M_.a_NUB^MYXaWR]H#NE]ZF2A5C)1KF3\8-E)0R>^9
)<2[T6UVD@]5Y-XGT^6dKYVXLb?+O&Y3O)PHJ6U]>HY4N.8>GR8R\dE:86+E6(O)
00F_7#F]JQK[)1g;??8SA&LH,W)YOE]YC+PLBSbaO><\]D;?S/JHZBb5.V-2EB1M
3QL03YZQH:S-41NR1U-8<gMH<+S3D?P<c[&-/c.f5ZLHa266>Qae5HTVFD6O#\C9
5([]0OXZE<^LE;Ug/b)eP9<).4GX9&<R2&cA,&(X1B=#e;dK))3)HCS<IYJI[+d?
Z1R]SP416b(W,=0QN2&L#W@Q_>H)JEAZ6c1Y)H_\.4);[5]O.](\cHC0<d.d<-NG
Y-\IMYDDKfYO@EZZAYYG+U+@b+\QRIH+?#1TgQC)7XI94NUEA7a7NAX>(W46FNOS
&R#6gKTNSTG9/SWgW@eLf._S:DJ?<2O>U;.CWCWE8g&E8]SGJ,Dg1:]6]=YTg883
gc,&WYK?;,25[5^gW#3<TIUc(-c2P#[a+3Ya=[#O_>3[.VZd>&B+L]]+[Vbg=YFS
@)]<.>c9F?W.WgQV@B21^_9ecPAMXXAO2.XD#I&?77?/O<L\Pf&NA@cJF_^Z]D[f
-3+Qe?4593I?AD&18^.c(TU5]]_PD/AJ5+TPIJL@Gbc8IT)MYB+_)g1e6gITG9W^
0^GIcD0^6KQAgXXNN).+[#8\VK:DY176Z17\2b4@)Rb2F2QD\b1?LNV[QCP4M0.Q
\Pe\Q9)XD(c[f]Z0-4NOa8g@BN9K7S(;19bL\4e^M@1bIf0fe+8H0YSYdf:N[:B;
UH,1]^72JbF0bD0>\Nd8RY5dU?[6;;_<PG.gR.?)bD6DX5LP^JSSBJNAeOI[::8V
=8@fBW4[KW?Ice=@IN)[UZSL-]M-U7@/;-:12P)NYR.9P/<N0.KT4974A@EMfCR?
H_=QH4]Y4KUAN##?&EZEU+R[;HaT:FEY:AHNK<UR8HXVFM:a+Z,\:@VP>>BC./U.
04[-O\EX966.]5,/H].2MY:3\0.;L?f[:bJfg?7&PW:B)a0N+]R^EYO9Pd0,,Ua0
@U.>L+JLV@dHVaD&Y(3M]gA?Af8)<6g&fE0Wf.1Ged07L33BIF,2#&+a:9dD&D6_
=SB]MQP:FNS^98:TPP,^VN87:@f1NZM\7=OJfA@a=+DM/PQO[6LcLJUbJ.8HB#Y^
D/2eG;DGb4#eTUJLX=/S>G@3(_1R)#59-d\BPdeS7DaA=_7Y<W,dM-7]&-?B8dg4
6V,+:MI<3#^7F&:Q7D8-Qc8YKUf1aF]1a<RSV;+/;A<:HJ)81-gCCEge;@,cU5VI
b-D652;G6b#5De#E>^:,Sa\_4J-U\Q]]\CTH-?/eRW2-3PbT>,Ke9e=d5CY_;<T.
8[[BS)+;3K]/J,^+^<Q.K1.?&f-8W7)gX2S]D=G1=/-V:F(X^G/AJA.R2ML2G?f.
_:6bC2+e1]2T:aOSWOg64C>[8;eT1cK#0:JeU\ZfC/8#L<7A/U)CBT?WMB;5):GF
?\6@Qa\3W-1?<MQO^-+<5B7\gZ;7-fAbU2DRJ4DEL07/)gd7U1bR1Q:P9Q2-5Pb7
U^SHR2>2388,SGUMD-=85SU+7#Af&\OM0LP-,K]OEMW&W54a:1#Z9R#>D7IAF]2.
bHL&^;.(b)LZ(:4=^HZf5JH4B:0;-7(V]^J)Wd+C90>VVWMEY-GGgf4U1+cM8EPW
SOaQ84)8YTWI@dI,^24ZF07RG>?9:T,>ANR?_@cB+-?c\TPe.6S;US/D.a9YCWOg
Q98P]GHLD:NfZFA>,46#[@Z2-&0M)GAI(J@8d(\a_2ec+_;B5V+-RXD_OF1HAT4B
2XTEAP(cBA]JZ:g36eV8+eAe2+V@a6XUP.Q1>-E&H]J=_DTBdgM8+aTEc]6_XM,g
f_=eJgbT0S(05X^f?cL4.CDe:]3g=J0]CC(HPW&1-4,:-BCILXaM\I:YV0DX^<H4
d^P_L^C8IA;H]9&LI4G4_7GY2ZOLCR>SQ:/CB(Ic&_P62>FYD1QY1MU04^RB>c6U
42>QTadGT\S?-bEJ\)JJX7/_e:ae&?LcXEW\]B._-BH#aH1[_&-4O/17XNJE)RMD
CVC^#+g/S3ON:AG7NdF6(/VM8dBaaTMbVP-c9J9J+/3A&0HUX]fJdY\eU2?2W64C
0=&Rb@\V:1M(Y=H1>YQb\ca=[C\-ZJFU1&D#MdQ-A=-D+F[JaVacg,-0I;fWHC2,
CD#:Odf?:KMGFM4Wc674U5S7d6WbE0I.H/6OcP:_>MF\1]@d_65I_D1/,CS10OO&
8.UL98Gb0FV_bNXeN\)/CYdZ.<&G6/+3gE>[GQ=6@CL]^Q[G#BSH)S9N7,(Z1-+1
/?/_,Bc2K39YU<F_?BN[5S<>J:?EFXfDI,f,g,B0+DbY<.^U6=WJ[N=,C_b+bM,S
VIT5-@]#1I9N?=(;c):/,(=cQ9[V&0f.7?B(6g\B4)4cB4A+]_ea)?KY/Tcd:R1J
VaB>5CG[(14<a/.aA2DZRIF3=KTd3Q)KGCWS=9g,Ae^eeBdA?48gdG9H:;>eJ,<C
f^(NUB1?&WTBFL(3D_g5d@]@Q5bEYDg1Z6LFeFCPX0;dBYN#3bc]b/F?QT631OZH
9)g-H8eQHYB2dQH.ZL@4a<TZe5[[,461#9+Bg6Ge\Rd+4T(E@5R[&b>7SMD6PPGZ
&W=?H((VVJ\>-W)#=GF-S3QNOI,L8F-cZM:Od_BW^R5Q3gCaZ4;cEAdI3BLMKPB2
^)]a?aaPc,D#[FJGC?PNOO5+UR,=A/O/C1c88d]U-[#MfC/MST-EdP_N596J1?c(
KCZYKHHc2(;]=5g#0+?g?><X2NZK-bP3WQ=)9GF0)M:COS:W,Nd)5D,,d)<dfDE#
/7dO3JV012d6X/[5;/+,TIU4TVaI(e-7QL&TVG0X,?g)B7ICGLIY\40_H@cM3GX5
BfMTeF[>H&)BH;(+@de-F(FDT1PWFSIWB1],PY:[7J1)OGJ>AQ_I@e&#7(Dd?<+M
Y5g0<4a4WQ#^<edW/BNdGV#:5fNA/@@B>EMK:B_We.:^,JaYK7YB(dOa2A1cC/6V
^D\+PeYf]X;3+)a#L(a.8D^O3&NG9\.K_U2>G0#1b4@//Q);,3#LS\ee902WbN)L
:92)K6WH+17LG)D8g^9VOdY.0]eMKR-8#Y-GTD4\OKD@2S/-b<bGXE1ae11C=XX.
]+dPZ)P;CN79H9U-a@+<\d)c1F5abHd6_EAF[a>I7BJ66E[H44^G=[VP@29)85J=
5#E7DT-c+d8E8(QJQWS6S>0+>-_XSCV=J6BGZTH8=S.b+dG7N]=2RbK^RR1;DPAY
9>YfKF5E<O.;c[02+F[UP0XAUT)OAK?4S;O=U3)^G\b]4bJAOT768M[I,2#>)f(O
M2V\-c\S7XYPT[fd9;e,),W?&GZX4ML/@,OF8bL7XSWV:Ab^eM#Y-/\Z2,b.,NA#
6J9A<T]eH=52.6;;<+\[f3A=8U)ER\(=1)I@ZE9T:J25,JP;:L.B3.48W_1<-&Mf
I@8,WJS)EUd@HR/_<SEOHE&G7RO0@_\NbZ(TIc6_L\<RYT>/0=TQP#:]UU=;NAc<
^VdLL.?/NT/_f#-R<34;&K3638SXF?[/0N?.?[@V^06[/g)e,8&\BVUCJ&2-X)D?
/I@QSM.38(RdQ<L7fE:WJJ4</f,8WY)&N#Tc#E36X)9AMO,,6aD,W_NIX]Q/;gAG
[-YM_R-JdR])J@[a<#^KK:3-Aac4[Z8ae1S_3B:,YA:.g@-I[;g5G67+?Va81.5B
H8.;+>T:U&NXAcQ##c-\=3Y+aDT2A1KK@/W[]],FW,Gb599,A?Bg-<d:_7/K3I[)
2NKX;:J\J<\<.4GR-;b>RN8#,=35:;WCHePE.V>a=MXggfa(<HLG>dXabAX#<M+I
S8Z?A]V&G/2AGNR(D0MV:b>95J<cV_XRM+6([6:FbTQA5ERKH92,?VY?<9dgXT)c
IKVT/(H4P#?7b-6G#O#Eg/^<M_T\a;;B)RMY#8YBKL0dc(3-Q[\),dZgQ;8&NG;<
#A)MIE^]#6XDdJ(e,HcBE>OIb2I5/7^,XXWfNF4egaA5Rg1Q(;4a<(^1+0.NTLOF
@=456+<E-;S:1N1#&&W/HL9KOWPW,bPd#RGg:KTTCQXK27b/>FMaWM;\/VV\>795
eB:6\9cK#72H5VUMdgYfDL/R_ZfZTbZ0B9_Y\Md.9P?PGe2#U,L)BL/9P3>g6b6?
g&<I=RD-M1UDd<cRIb(F.?deYG<f@\F6F)U4G0]UBZLIddd8NEA&9O5MD)1+f@:3
fK7:L8TeKEe=Ng[KgVccR@XH0&CA9EI.XVLMc4N_4b1KP6dEdFac^5(a)9.ET\9V
^@GE_AeB3GX8--dd-R>YA(/VW8+TbB96SAT>QE_1T-5b7\c<HGMZ+5NbAIL7U=PP
[+QAJ;[8REI/I7>[-aGPa\LL5:6,,S+7UL3&bJP/XLDJSEBg/W5039V.=258bgQO
Y#CK0+=a>]gCCH:X?LE,[_7Y,N-AN\HX39ae4aCMK@cNM8@G.H.F.\32N>BY&J5e
eH\1_&/-YaUR1dQe&@Z<?g4#X._LDZ167RgZFf@)ee,1_YSPZ)-/;aFVKfVA>E7?
.>V3.C;BZPHK):(T_38)eOILaMEH1FY:Qe<@(]/KGP(@8Dfdfg\FF_S[Y8S)UOZ+
^JV1b3c71.eE/5aFgMZI8<NA7dWIM(^]?SJg@MMFS?aS-1\]8;e;#Z[2c7.T4=bC
5ZY</-R6C:(ZMZHYd1G2I.;g(A7,E]4@K5-eQXcK1914KC7c6D=Q)I\/C<eDO79]
e7_]H;D&.L27:MX8:Z<,+45RgUIDe)C/B6.a#-8AWZ1N;Kfc.VebNb6+Xb6>,V9U
d+108_\1(b_\+Na^bV>d]Xf1?_X5X@L:?J00Yf89=D^D)JTMSbb>73OUPQCKJ;JJ
bFFMDa,=)2]TP_TELYH_N/S@B+<(beDE;&\I]RXIe2Z>I^S^)FU61^e)G\,KEf\C
&g7I_Sa#aSa@(#35gb5V;M?FWOX9EC\=Wg3bP9N/;0HN-,dJ),8HS2>2.2NJTXSJ
@CA9?Z=H03/_DTLgWG[fTT3)D^@I6LfT0^I+A2)b^WJI;.N+SaI43^fRUcW&OF4J
ML9MQ.Z;;#=.>IP.K@5U5H&C\I_2O/I<,OJI)UI=LbM\/Z]Y2]Z6,[OcCD2]PDTO
(b1+3REBQTNaVCU5CDE5d=?N\:Z7CCI(CW4=3P8g8L@9KO?SHK4^#[E;XfMYXeBN
+GS7L0\\Ee16Ib^SJCODgS-1#X),@++ID)DM6JB=eXM</@-+(Nfbd;:G,c2P&[.a
gd=#9UC-Y7]SedJgW55NP2OPMQ8(EeQ0\:BB]f^JNNaA,HD@=D#=R+A,=a2)4R)P
c=JgI9YL;eS&HMeFX>NW:+]XCP[K3RcKP?ER@N^4@8&=X=68WLcOC1PZbBSDe#F/
++cMP@fP)A\D-:gH1Z-TD]KeQ<bWP:@fIX[F#RaU<A[XE=;f<<He^][bS:FgO7?8
)d_<^gK#,7]2\T7L8.N;)BbE9/ZMJd0T&c7LB9QHRDIHQ7IV@KG?(dS_ZF=b(61Y
eYCaO;4Z8T7(R#gPQe(_YZW+W1WeMA9CZB;Z5ETTLb[#-<^;=>bPL(eSVfU?A51R
JE:??P=BE(XH5G=8[c)(:dIZALQA,0L,Ra.EYD]+_11.fJ281I(?\\\)[,UHSSUb
GW.F_cC@SEV/T>RGEQJDWU73/Y;f&,0W]C15+Sd@A]+<;]3Z[9#<BS>4#@#2JC6J
H6\ZAC,bM4P<BRZC@-PE(/g0;+??^./S-Gea(UG/Q1UYAA[PA#OGL1<,ZYJTeKUB
XNb\&TcP7X]P;9;6,5/?45&.C);I;E-eY/a\5^ceW,\/;>9&.6\[2[0_+4J[b0-5
C5=HV<J;,_@bD:VFHY-K7Q]MVWH&5<<F7SR&67I;8JI_::#1#V/P+L7+=XWcQ1D_
D3g0.5bcQPA#BfS]\=(DVP0@g&H]PFf\0PY7?,RQAS6f<F=6ZQ75d2E\#<M/e_,;
^LRNS)e/>?3N=f.I4CV]OX/=(^b0dS),OV_NF]bVFQM=V7BcQW/E3>4TK8#]A(^I
^e3beZSYB)1D6IGUXRcX3YPe].]H1_3/;>9N6<N)>Q=][_I+>.f]^2ZOOET78WXE
=ZbQ85A>KbE?^LOW>R[&L#^2)5I4UR1^2S6FGfa<C#BLdZ:\NRa;Ee<cD?YX.G<Z
LNZ-aQVPF[@=F30U<AQ5N^VDKYS&9ZALV:72+=[(a.VcZTA5F<^g,;?)M-P,c]^c
2N#XV),a3W[<8.NaNPbB\IF2.U24G\3AQbd0@-@0aL,FU:OV9cg#2]dDDMDA](;S
Xc8#P9WG/df[/USXEe1CKS>SaO&GE,5)WDRd2add^/gb4]MNSfK51J=2YS]<;V^A
N^C<#-T5);CJb]^ZIO1cLS2?KMV(T>?PN,Z/2=XFIT^M-JET5MSI0IMTZ0BMe<-N
@ZCQb#10X35Jg-6a_b8eag?:,JMCWIcE4^UCV8QeKKT6C]eQ^O9g6]f&##e=DbD1
GBM=_8D6T+dCJVdN23PDUBV#S4&18;_S#FN,CIA21a_6PF270b_e_T[eHdgeHQDI
gHO&aJ25fM:@L:aL?(A@?63V9G5d,Ffe=Yb??e>1W=[:MfY->7e7NPS4&^05eaSQ
KIBP7Q>-CB>>E-S>c?\+HW9]>OIb,-QA-&@@&>Hf9Ba/\N>R1F;B<\Z&A_#(<1=/
0]3PYe;>(@d7GIbdW8]I9-JTZNaXLa+TQ0=:)E),Wf^FdK+[Y:BgW1:2#?f&PU@:
?Y9ZP7K7D6]/S_S1D4-L--)V#M,,X^;?S.[B&P,F[GZ^N[+VCC1SXG#]7dI\NTT6
fC99.A6[10EF\EFT=N:a#L+<#MQbQd0cD8[^)^f:UB]+8457H]O^&IYJU_TNW9P/
J=ZH>GG8<(SR@E._OI\R6+:^#(7cCQ:W4^&[P7/I#JTO][;,LG(A70:<9gRDS/)+
>G,):M5K6?]/]_<]91LRJb0NKFHKTc&1b_#NEBNX#97@M)@WD:F[H\(a7QSgSHc3
]HAI:d>c,O+UPB??YMOKN.;A23^@d1fN?3M4>[:4e^&GXURd\-T(gQ#,T+^G.]]d
F-F?N\)FDN&.V=^4QIJA(<;[d=<N&a7#37B51MfB@A;C-+3X9Dd@]HB\:2+]bLYR
ReHUZ6GSV[JFBM))FXcS@?aca4;c71R\(eUV6Q&?C/-;9,<T+]dVIE>eO)b_)0cY
)X2LRN>SHg^CcDFNA>0cR^@F026#4P<I_eFfED><(I<RN/UBK><6CFM:XM5U.MLG
\S)=W#5_1-YNG\SbdQ6DES#S[e3XU3f\511a=(H-<J<T,O7<XZ0DB7DT,EQW3;YN
7]g#<-QOQC5I.4c\#Q?4:Nfe9FYG8_gOSLU:cQ>C8:G/>g;#:F8_1C1Gf,CH9TVP
S^.CW.aK2,^2a\S&9Db?@F4Z-cPDeCb.C)/J\Ne]=?@a<3G-,/WIJS=&R_RSAe2T
Y<@XT8)W.Y;8U-+gT^^)@A:[9MKM#b/(daT1cFXc/<dS;O]3fe.4X:/Fa.1WD;?]
GTY:ebF43Ve)/>6-ZLB#PJ44aX4[-GGS2I)U]WI-0dD>827=8Qd:e[N#RW]HT.P_
L2YF/R6U]/f@R_5C,3DD1R.cQf3Q^^5FX30eO.;60CV4WDLdU/X,Bcf^&L7W=HR3
YfW(@8+\KXJ<.a31\E=0=4V6LN),e@_(d/geVCdgH,M^g#E&EFU=]-3OC875#YTb
)+.::[>E26XEY_V:3?64D6GLT<5PdOSX[(dJ/gg&aTUYOLe,S@AfVfd-@;QPQG]1
5bTPL_;W+ZgEO_@<Kg]\V[GgBQaLKHCeTP,:]?28?-5KN_CC(E&WEWJI7g::00FZ
N.fN#S?=7DV2a/U<UD\CK+,#?2O_;1YKIbN+GLZ+ZD=Dg8+E?_2<6Oa:VX4[4[]e
@?R@GcTG)::G8-K6f(fCJ3-F0[[LP4.#J28aQ+&@7@US8)K??&e:ZD1g>).df2Af
TDPf&aa[D9@b)J]M#\QIT<M83QE#.YF(V:[eW240b@V=2,3?WA<E#/5U3/)L/142
>5Y7M1B[DebE]=Z^GX.2L=702N5Y/T1?9^I2=UG@B.#OdTUL1,-\dZ3N:+)=)Z-?
ZF>R;8@Z:::]b#HY_79&?;_>JLTFMM:JKU\<3VF+/cS[aMe8&IJOA.fQLM5M^YaV
_1&2b[Y9SY\(Y&N8>R)=HdR<-,3A1-F:C-_F.E#VB[6[D7+:AQ9Y^1BU<RFPcHN)
MaOSd)_e@.dIOFZY@-TU6/d:,4bV#(2<1.@C8=ATU9ecb.)FTWW050C[4H)g>bS,
TJ#DZDUHOb,CbDI\ggfGH+&]Sf7DG4>=E6@:=D>4BHQ]dY;H8BgI@-VO(;=E9Y:Q
c;J/_A]bA?FXLd[WATK&VBe#.KPDWY@3=K8RX1H8&((Y[V\8NaK.#R3^XI<g#<(I
:OUc:c=L&c>WOY8VcCKUO+;S:W<A[@DffTTdM0c^M]R_D(F-B)S-XRIb<A1?_&g_
D^cEF8Ide-dV6O84<aa[WBfa5c<CV3G,407fLWIF,R5>R&/H_[fWU85IBCfAcNIX
R5Sg]+:XcG.BM(JD3DVg:5bDfL?_NRKXB55:N]VfZS?T2:@41HXI1Y59?U#_XdfH
G,5UX^gB<0)^-R7\Cce&;)7+;^]#Q(7::gR<BS+]J29Le4<>+&5](C3Nb<=I[_)4
\g\Q:X<F+#8)J=K+(_eUTe:BdB+N6FPH1F@;ONQc2.T-d8d6eYTH/gBb6\JB[SJ9
a@^#4cL8>(YX2:2(=G24G0O[IPC6Y\b&L<E]J[^XO488)DD50aL3][?(+R,(KbTU
E1R)QMG^&]&ZK8?Kg-0[6^6H=A>^JEGIBLAeQ?>Kcd&\_KETE^gb#.0):ecgJEF[
/EX0dYF>26J<<2_^I+/J.g@Q(\cH;6XT+)L7gSWX)P6P->=.=.16/DHD&4^8;_IA
A1Z;=[bCH.DOR43\Q/-8a35^>TQ63W@Z,#?OTG/C(LOUEcF0^5AP>1Y;#Z<:cYSc
c@74U(_SA9a3/9C#A0T5+<_;RT6XgHY?4ZNIQ_/<_ZfLfbc<E=#C[A+@+NBLR=cT
<cD0f4db&WI(051R[B&3ffc_]W#>J0+:620PEfC.LBU7.+5I2CdD1[[G9-3(G#[P
3ETY^F4:c:3WGF5,(QZ.bgS>&&4Ae1XGM;U?X-3aT7SY(R@3B40/01@>[,S;]=N1
I[AYG<R?0.^XF_S/OTfV^J7\?2(KFgCeUB/ZR.F).)D>e\HM[=G,0A^&GAQ<F58Z
PR/7Hb&]aTAeGUeR:-&;5ed+\_+>/&3^W+F,gd1\YN<cHZDLCDafMQN;ZX7T:9VM
bb;H+23S-21+3>DZB:6,34RCCb9Z>9E8NWgE2D2WEWDWK_Q6YH<H)7M^aE60g(3S
]AgffA])NAR5(-5E4MXB1W)+eOIe8#6RL&ZU0?PFb6VC#d8M][+<G+[Q\BWb(((e
OK3#4=JYNBEHCN\J2a:4dHFgF\4RBS^M_P6<OR<^[=G[N252c7a[<RO4E[CJ7U#O
Y]=,;e\./2)]X68OgbEA#SV:VFf<R=)^4B5bB=C39#[^e1U\ZfQ_aZTLUNI+-:-F
96O@I@LJ=7Z1>UL(H)KLCACBIT=ZO&G[(aAE-3DQ\+MQ[_Vb8&3U_:@e5Ha9d<V7
,:;[[RDR3:D6-A:[WGQ\]MPBOR>;_@+VMIFH7a&=]8gXDA[6b>BL5JRa4YEA3P^Y
#B4]>5WgYR@J)&0JcCcO=W]ANINMKA=Y5JO5d2&.WYE_LJ>,-4X\UIfVJKeP++cN
fF1UR/W&UH1BAb)H)gKe1J2K+FH4P/U/f=SZRgZ_\_LdBF74bYW1R+T,dIJ4<41\
.cdY(#GRG?#/YANBGP-PC_geUH#HMXU@BE,03+G3WeH+Z@cdf/A(4cLaVW8H&7G[
?6?UHeP#_(-UR92)O/-)g&&8ZbF[@I[H9b^R4[#=EL[VF9I0;)a-=6I)>9HA_Q:.
8XDFcGDIOZ^P0\TgY&3c5LCC8]PS\[H\c.b1R4b(A7:Xe>RQg>62\+f^#PP?:Y.g
0B[8EUFcD&1-g>Y^IYaeUC+/&ZD(@]d__B(b,7S@b0N7&)33B:HBb0O#aE#[,AQa
P?OIbKJ_GZ&PZY12Y<^;eXU[3FLCC-N##VLN4A>YH\=HC=A+/Y>,NH#PKPD+M+H_
-WgWe&73JM]K,)O(dB4N20TbEO@]PaJ7-#,IXB8<g)49WS0@R+=][_,,N^I82VRc
]e)/&[\A#H5B)d.M\L=@-Nca2HS73aZ0fAQY#YY3,/7G9J_-G9F>DUYJUI7X][#K
7:dYI2V>,GXAP\D@HF9WQZ(GK:T+[FI010,8aFK3J9XdHd^#4]49K<#B7\DB;<a9
Z^(baD_)D@EP8KH7]XC<715Z:WMLXVe>7YAK-7+H_64_9@A;]ACaWQK@d#KD[78=
.K+]b1R[BgC<2fcBIRZ6UO,-,FT.1?,BJ4Z6?,QQI1FcEAZUD@?7^Q&,ac(EM:T,
gO3fPFW#cXd3KeJT2,+O+S-9MW,=Eda6O22(?YLTBS.f)Z\d9\9D;CRK443H3+LL
a=^c7TFTB8bCM8MK:EW<=.<<&7[9V(T)0DA[edI)ZZfdK)F#T55;8U5J](TV#U0\
X3\MA.4]17,K@LV\Sg=62PKUMCC+/8,c-;(294FeS)e]2\c4(?:dGPdgPaF8eTdE
P[XNA/3?>)KW]ZJS&#DYOU_^6W_I2:(4OH3005NJ+Q=T2?)M#RK+KN6K>B\FICR[
]];.R[dPT;bOH^5T_OU4/Z?F#0UIC2De5<a5;N]-);&I@G;8[2Qc]W4<R1#5ARXB
#ZV_IcbNfN:-9J#e-J\6A;Ug73F?5KfeBM45X\O/YBCSSO:]QOCU<DbKT.;B8)Q<
Y+Q2_WfLFc3;GcbO#,1+#B9dOJD+:-WV.46+X<d3GS7T\1fK)CXNV_\8W1XIBEL/
5f)VVA]A0g8MX1ED@S1UW&)/2-SHE(<#/@<G:f5YN]#4QZM]G\;g<PeYOb&Q/6L5
V@9._<<JY6.Y/gg&HgLN)8;8]^T,^B.S5IK0c3eEb/\]9OM+#CUVVGR)1#TH[(O7
b5U?U9S@=+XNQ;D7DCT^,CT;a</\6d&WWJ9N,^J=T^-0&ZU@=\7OLA0Y8LQ@N\@c
FHSHZA-Qb6-fOW1M0Ra=d<^L#00e3=1+0UR_BD86VWB+5_HRd@F&)T4OPM:\0BOA
)]g89=70[>\DLHZfOL44\-/U]@)K;?WPEK::9)>ZP7YQJ[B25-ICY^1=ULQS-+JO
H3O_Gf]SIXIA6-@7>V8,W2Lfg?dX(;.>.eK37dL4/ITQ[HJU8G3_E5[c&_USQD,H
<F<B0,[/8NEfAH(R9TX;^@RB:WZ1cW_3>M/f>ePM;&DRLV:KD?7\D</Y2@)T;)-Y
#V7b[K5]#bad@XUTceE,B/1L.abV]#6LdCDLPKPZc2(0>(:,7fB/>RJadd/7EY8S
aA9X\?O4F#Y+KLK@e7NBc-JS&c02T]_>&I49^H2ERBb-/K<EL69NBGaAEWI@Md#S
+bECS9\bbF<@)I8.8ESMRW+.,[3V_J9,?4Mc_d9L@4-5ZMSNC#c9D=5(&f(53;S=
QaZ3CUCSM1ee5#CY\=Ng=)I1M<(=DT(IeBV220DdbS6CMb-Z2/0_#F6gXO2\<2?K
a-\.J&86bE]^,X;/ZXE=6<7IZ^/;W]K9I=]7-#6XCN+a2VA(-c)U(<IJEE3A?Jd^
_SJbN)>:71cUP[,1QAUNE]Q<E_g#L5ME6PP_3UB-29V;aR7:3(N.b(b2][O6LNcd
6=,Ic4aLMeJRHEK^3];7=UefQaZ[K5#-.I2fNQde-BbJ4F5cAWX+-&F#>27_1=8/
PNd60(E5A<4.J6BO_-05VW\_;N&XU6+N59>a1S>_LO=/JGPV?P\DLL(XRb^R8JMN
U5B.LSF<T54-LU[FOL1\FXW>62];Q#:1gTI_CG;D[TN:HL4SZ8\;a5G_3eUL1LY^
;K2&dbLRe1[(@(bH2/Ia,Q\2E1&Xf@+=AOYNS-Z^b>;6.d8R&(He_5Y=CAP=;H[:
JBG^5bF&+7&0JBS<RO<g.,4+BL/@+3@gfAI;[U9QE^L3C,S1^b8L:8<N7KHZSL-8
NDP.SEW&QB_ef9dD5-OL,PUc00#d12SCS(9AXad/]&a^I[H-BX_PI^(QaX=]daEP
G8Q)I^?QP>f_]JC0]A@K>Q.Q]c/B^<S<<(=IN0X4FJ56.RFA9X<eS7bS=;W82LFJ
d.73CJTT\bWR059Yg0a^[;FA;(eBZG>-Qa-ZZe#NILMXZa1Xa;Y\RK)V>Tb=0]M9
LWQ#R6X6SAbT=PG,;a/^>7gZI:g.CF;V1>f.6eG#a27b?0.5[<BWfXUC[CD8dG)V
>>5AQb+8IIC@?S:FE\I)>D/7<_C2D8-VJ.&AGXQf:AC,D;5e]F<WOdg2E5K5L)ZF
2\6PM,0#<NbVZ<@HV#:O?+RJ5M+J.9SG,fZ[PZA;X8.d86H6F@3N??X8<DJgCE[V
)4QY@+&LUFZa),QXW(IAK-1;K9XgT+7419gU2&/2d4BX<X-OQAeY^[SaU-bRFMa?
GG5@@[@,]S#H.FgH_(/_>fdQX6M,DLJ^Y65WC7S<SFG3;3]_K<YD9VgF4+L_?@AL
:4.>LB\R0L8;-YL)T:B;6<1XMV7B7bI0,7S-1J1U>R4/TL0g:bRfHA1EEYd@-Ig+
6]Qf0b.]/KF=#GNMB_>HSGc4N-H\HC874c78>W=5\=4P/&N#E;64+NIC2M_QC7gc
19+)]@MXXFfMTF,XYB]@3A0CfK7T\G#E[;.<SQ^<FP+)?9WcbXLPPT_[a&)E;/?f
8JUY5&0(.VFMS6F@3cHc&GUQHY(15b)Bb2+Q719K/]NEd1ZKS\R9_D3D)c6gP7e\
0)d]9c3,2HM??UPe</8>^Q;3-DR3bg#;BbV9HXUAb(27E7FDMN5^/6eWe[W@;dC@
,G.\Jf.T7(ZW3D1]d?7^OX8M(1YDfI@ARdKbXLbEdJ:8G)@228>Y8507/Sde6P\+
_(#OS/)_8a+NZLR[/B5-#aYO&E0fgg:E\gBa==^<L4;bJ9)cYbe-###@b[f,C8I<
#V<(OV]L>G(Hd[_CMaOac.JIJf?IP-8eIg3K6g;Nc#eaMP[)SG7?[&8=[4^f,LO0
915HZ21K3>]ID[EC_/Je/Yd@?Z>AC991M^g.ED?VBNGcd^Z1QH1#T\:HNf2-=1D?
<8BM&DAP:5E+B=gQ;?NPc;?+B=/A6-&HG7FC8^9C2<1#?b2Y=PDH8EZGg8]RMf7\
M4UC7&dO]V.W45J4g(UTVL_]31AdVPfF3fCR>U9]TJd/J^H(_]=g,4C?+9)-J;Z\
_CLWR30E:\<IUb2TaUSMWM<CEgf8fU3B6QYUMYO1T:=d@>._5ePaeAF0Zd((c7E8
0LSa>D#^G)H)<2DYHNQ@]R#2=\5Yg=T7^@W]1,8^BA)a6L<\[R-0;?J4E(^d?2_S
aQQ.16\.W6XW9\W)c,X-COcJ3JBK#I])P@Y:Jd\:V9.<b=/NA_;MQH,Z1/A\)#(N
/A9OLW^S862dWO9NaE9<MRBG:EO/9]9350A\eb0ZD/.e-fUf+HZ<]=>=W4D3#N2W
]H/3UHDBBd2^TX3/6X4NW<8&IU>XeT<0FFZIc<L@N61]IQ]b0)a0E_XXRPbRJK=;
.9_KTU7IQeD.T1Y.]6,[S;X(V;Q58(7bbHgR?3]#.bOMfe3A_F2b:CB=R>IdWCIM
-\I@-eE5<=eY2BW;4.];2&[.P3]XIVY?Y/IAa?EgZI>SX=NZ>];1bMFVa6(5<JGI
dN;Z/aV+(65Ma2b[J5-X:8?@52/@T77>=DQAC<&RW7>K0-(PU+aB57HS]\Y2K&8/
)APB&4WI;08,Mbca-SLM[D#XBee::U48fLU0PB8L7:44bFgNU3SUd_UbXDC/gYSP
&Dc-dPHAaQTY+HFM8;25W9G.eWYWXdH3_-[#Q/XQ9I#:O/0580QX-J40OK5c.DQW
:XNXG375(.>E7?I36PUM[IS;[M-dLL_XaM9:IOG7Rf^V\fS1&\B31KP=/YDS1LTL
[KLJO/P919I(LZ<OS6#MVT#1gP^9[+;N48gT[,L\[\-P+13gg?21I+NK_A]X.2KN
,EZ4,/,HO4BXPcbQ.3N-2#J:-bZ1<+[XO5=0(:C-:R-3bYW8<X)J^Y3_#@P><(b:
U[,P&HE.UH?g?PP/3MJW,_D77,HA[L_R52UJC[ZN4LH#FM4Q#TRMT+1#?#=:-cM3
)&b6NSf[>b,GTPXcP#/@+Cb.FVE04g(Cf/Y#T&<K@JR,[.ZNaIOGE6>L66dad;<4
V8,_HKF]IQF.8UaOMYC9a99SK#V#L=V(Z6E&SD0LdI.9CGMHNO2#OK1[LfJ8+7@9
.I8RC.b19,/62:1bP.-@]J.I9@H5K/;Fd;QaKI^_N#e-SN7FIIN6g=,,#-cAB1A+
1S&R/RB#)8^[b>O>DDTTMVPGG<A7RJ9PVF.H>F3PT@J]g(P1E/4\5eL.[0_J@N)(
@NdcOC0RAdNA:H?.5.]/OFC)((TA8D:0,U[XG2Lg9)VLEeS[T+RBe\^F1RNOaH4.
7<#W;<BJBSd8TK3eDS6_JFP):\Y+/406&4VKdEcB0Z^I<_4L,I<a#LX1Xa(D17W4
6S2]Z1+Id+eEDGg2Z.\VP.1:<9DH\8=ERGOF_g87#A1(\TP8718\/T9:gA5/T.1N
NC1B&dZ4T=(dKa6)B_-QS#<GcJ=#BfOJe+R+LfH)\K9@?Id\ReV_>5D5M0FecJJP
;:P?(D9V2R],ffef4L1bSKYTNFAERK5B],HY88Ne>gSD3#^d11G-BRN^UfaGV6ZG
T2.L+?ISH(DeDG72U3PCed(75FC80Ra8OZS2cV,3>5N;5X;5SB6SaM=W^8?/_B?O
:c>d@D,M/P.R.(1LfGL_)U^>9,M-2K6OIME-6T(F>e6YWgX#TN;_W@b&1#9TFW88
+8Ka@Ne>5&V;PA-bH]C-\\Q06;77@>N8PHVQ:X]/6f1^\gKgV<EBBSV17-(Oc6:R
Q7_R>gB^?]+aGDQ19AFO6MFOXVW(/T2]7_F=HHD-W-Y>>J0R,LR_=SOD<3bgZ+_6
=,+J8Kb+O14b+EH++MD4_@GMNW/6BBO^X=2?1\AV=Tb=_==A;Me;aQ_CL08+A-3>
;^1&aF]:U1Af1MaSccL;HGdEY@NP-Q9YPI^0A)]K>S=T658GOg<L+-bA>^eZ4/IZ
4Q^3(JSGH-8S4d-P17OOD.;c;cOM>GD,Q.OEY^B8,&#>XdQY:B/@GR1Ee724,H)1
g+EO,+gDdY>4=Ia?f_Z_aL5K?4)Za#F4S7QC-dbbP9UPD7<+1\C2cF-)9>HS8]F8
:U5g([[B/B5W_d9&2Q.M1^_,@4TaeM+efZ4>5)f57(=Mf3RD7/L\X=W<gbC8]E7/
V).cMeJINbe2.T)+S=QX&MB#Z]LVK#1f3B.X8GMT8FD))68BJ:EIa[V(A/c>5aR-
bKcSCJ2\(C\F<@]Sed\Vc)3(d/X:0Q5NU]&O@BMP3fM2EHR>Y_Z)K(:@.X)-g2fP
>7C>NUQX<OY=GC44(6\JS\W9LYU?(fX\H8<c,/aF2_e>EZ8aD+V,77Vf:DB)65Fb
RfFAL0b8<9\?NY,Z#627MF;M8UgR?7g+L+##d-Zg5EG4K+bLHJ:AAObVLb/JDDFg
H=a_d?G/W)O6X_#YU=5aH9,_:)5eBE<\MbY:ZdH4U;eJW>286[CJeZB.Jg@?I8G<
gI\.J^IQQ^TLA]Vf\^<#:<]/Yg]:]QD-K4MPL;4g_I9+-f@FfTb1&([&>Bc]XS&g
bH;<82CEd3<6e(?ZNO2E>==E+32N&0KF;<.EP-AC5@cZK1SPAAT5)G\L+.R1@^#T
/DQ8V4Lag&a<5cYC>SH(c9_HVQBeUQ7K]U(OR\<=g(9#[4\a(2UA[:W5DQSaTe<X
L\8a9cgL/7_Pf;3U=b:+bc.82<\Gc\J&L3SfeO+-_cD\B13V31>?6EO[d\8>O[@I
QCE^CReJcFG9S(gC5_+F.+W&]9[BUJ5MA>aD3YU/aS&TE;)=QIMBE@.=RK\+:0(S
;:Faac@,ebALDb/]^T^.T.SUT&IPA>?UI0[4Y?^#e8UFC20[]74Oe&7QcXRB2ILg
17(AV3daE8/g&I[SPRM;J=]V(IJ4+cY;T1R4&f0#20U)K:7eCT]ecV0J2eg7d&1+
]&17dD0\)>;(fX:<O>,B87VI?S)dH1OfDMQY9=Z<>T20;FHF=f@55@_=/A?1IYK)
;H+>a[F1.dW1ZD0e?fC:]6dZZQ#+^.)23;bV^9J<MeA,da4fLGQGgS2ZXA_V,:f;
EdN#QR3=&f;LU9GOYK?^@a9;<NX.TO6:g0,_:;5FJNDC?G>ba-((YT)_9GX^OPb=
^?PT>08fM?b5G&<9Q01XCDd0dRc8M_[b;/5gC>ID6H/-KS@7MM75\C<e4CgR[?Ze
:;Jd[cKUZYGZ[ECSVT@_E(O>DLY_3/&dgXZ1^gP\_@K-7>fKDBd&Mf_Gb3-R++TY
HH(IBELX\-.B/>QF726-G];@&e<>=[SJ8)]^Rb3Q[:O)_S2JFdQ9;J@g8PYfd\1F
Z61JQP^;CF=e.SYIIgQZ2PDL=BZGNQ.[1YKAE6]H/)?&Z-OT]XLY0)CgAYW,E0J0
]85df\I)9XJD(,KMC8A;20]1Qc&MM+VX2U5Zb&+Y8,Q[__AHNbVa./81M)ZY.a\<
Z245B8=68G&7VWdQadMeB]FH5)bIE1#UGNa&0.LW=eKeFg]KCJV/3>7cVR2WB&4&
<GA:KA2HY0MER@Z7DE>X7SIM?#E-05TcLWQFXTL1/bR:PV>]XAb_GcG1B6(BW@8Y
)K^JT4V7[^8&(?ZDOd=),=LDHD,V7c+Vge&HKNDA2:,=XUXG9+:]1YdD/?Yed:-;
F-]dYPQ:gFS.)b@9W<R\W7ICWDa@S:ZR;^EM&73BU@3,.^6A-#@:35U@CZ4^E^EV
?^>LY5<)G^N&A=_,9N1]\F,:DdT0A+&SQ;<6PH+-O+I?>&4g.<NT3BF\.SZgH<L&
Z(R<?bA#FC-:]M2HS]<\b#9UdD1:cHgS,B_HOgA@58@<[7/O::U<>@C0#8\H3R6a
V1BUCTW8Q:4?UMbS)K8Qc3WJb-Sb3KV@R][0Q^49AF6?A);QE)51#>0C;>LK^LgD
QZcZ&OI4<,fRd51).4-5;(,JbF\-\+[e]:S\J([3/.]c)=edb(0)3?&QL30\X/dY
+<<ZBaU<S#SRO8WJ;CFT[1bNaMW?MgFE&bE3PKaB?06fYXf//IH:>H^D&)@.:ac;
R9Za+V\I3f1:e)0Hd(HM_)BLHaNN4K(X#0N,F[0WGBO)W/)<(YggaZe[>J_f=(^9
[1(UHQV?/_c9GbdWJ#6+66>+Z&\DW^caH_bbGLOd?^L8R-#\]-BE4U.POEZ3SM,7
2c\/\>_a^),A>U.HM=eEL)4eK:O\CMGc)<O1cBNE>^K6\TcEX4A:N,_P7YF8WDOS
R7([VG\L11&gE@a2GWP5d8?YP,IY>SBIg+&X](8ULPNggd0I>V?ANVW9(<0Zg-M8
8)[0<-+>MAUS&S]&9PeW].[:<VJG]TaJ/Y45S]=>CZCbO]>3dRIKTIH:53Y/<SFM
?Y)0QcG0X7Ub4]8N[/Va,1d1J5G038-0B1UTR2-,DL5P7R6f1/#NdFKM?3BPH9V)
\_eOX=X.P?8:RaTc>6I>Q8Z+.[6/UQ^D]H,UgTaH:AI.d-UNE<Q>2:DGB3e/K+2V
^A[O5893^F)&^.F;V[&F;@C6Od?.6A_MS7/-bILG<3.8Y0<RN4BV6QIc7g/@L0HJ
]B5:W__O^WdXA4cF/f<8&QT22RX?f4eP(V?(3+<+0::36B(fD6f5H[HWaC,PECNP
1S(&cQ&EE30M[Zaa&Z>0NY9J.QOc-J73752P1CTPa__&&PUS9cWU-<D.1EBG8U)A
?XN@1g/WOaE)>:^:>?Af_a.ANGBRH+2RE_EO?QR-<(R0O6[C>H-;LO+S\LPH</4;
9.B.<W9UU,E4ZH,\QI\FW=K0Y@DY1?Ka=c>Mg7L5gUK0FJ6<:9cY?)=VgcRK[KY=
eLU0[AQ[.cO8gN,5J.ALaL^1F_4UL^?97KQROcB9DYgEMRC]?6&^c&aR^D5>2P/V
J@&GZ0_640W2+ZA,@RIVI0;3Fc2FVD<DdJI\EM\2,E9;N#_^>\ZTC_35GAEf7^.,
d<-H8QJ-YCLf:5G@>Y6/TB9RP@\B?^/d;Ie)Re(A<+5FZV4PdC?LfFCeH8ELI^;7
Y1/I)ZVH8AEFMMSMM,#20FR/D1:c;JGS.K[RUD):a(0UPY+NEH22:KT=G7[^dUL6
=92EREZM-Jg>.3+4V:+LQ5>\DA1W=8N.RUH[F@fPSP#1G@-N\H=4J\B+RTaG54V;
ROdg/8bZ<AF,bY2f+@\X&e)2Y#U6:6LCdeX/##g(ZIaJ@@I&#,_+)+^DaY-@,UI5
[R(9S]+0F-#FWXfP/=)?d0>aJ/g^H26@;)4Y/W<Z1^bZJbdBUM^ON9_I[XbMZ_L4
SMaG:OE_;<b6Q)\C\<Ga0N,Z:(.W(SH@,F_@Q:Q.=.^+^/PA(CDZM?((Y/Eb.0VW
BI,&3+.BZ0V5K:/N/8=+RYDM>[-4>aG\dMf;9A(GQFHTf9PRY>2.Q?2a7-ASbdC6
L?8GIHF<Z)=HJO;a<Q1#R9))L(B9@A5N@Q7.F##9d)65-ecE\:>D:36\IF:(W=5C
aW2I,PL2g.;\F2^:<&C/f\F/M?+db1RYZ5?/N18Z:d,HBCT/[I]\BA@=XL,>P]#<
GCMg5<JT(9VHBVc7S2LT?5@Ke83CA06+.XN?3Xe#EE84+&RX6&NPA4YL5-(I47^b
@R-fNV<F>+JB9BCWSg5)<)TaP6[QO#2+VR?#F.)O,Ia9):TZ_2W^,)FXRJ3EeO?Y
V-5FbWM:SgJbTHYA+:cJ;\8EL_L1L3A+6);V3Q2AU+>;eMTRD]CUa?e5A/3a4##>
T7LgX;B&S3UgBMdYW2H:V6WS]CUS-8/+X:(f?39dB:?>&fR@4Q:_7fZ36He=KZ/6
=b6cb]+/8g(Z@KYY(<L)@&:/FaYR8gD5a(e)38XUf@?.F[@].H;.]E/O=L?^(ZWZ
eXF?B3ZWLYL2UF10IWXG/+YJH_0#gE(YdJ:UNc/LZ/Z+;1Y;fU/CdRG]<_7@fV/;
W0Y&>SHK9c:)2(O?(NF/X]#A3\H(?+FSYNL=;F?_d8)7[MeHVV2\2ZDZ/CP#fO5:
_/^B.EG2,aVAGHKJ/T4S9NbP4DY6\).+R]@OS_^?+;Z@@J)H\aMC]PI0M37g0DE@
/+;&O.I;8SOZ.4e.6K^2IX0(-3\.@S4I-@:eAaT^6Y0cVB(Y92U6G2d2P6g8?;DG
c2(K2\XH)IFBc>]R_Q4Z73+SdD#L+QLgE/g,7<PAP@L^YI1L6A5g:7-Z-TVdN;[T
SH8S?bF,WGP+YX\3H=KD;O.QCIaCa@=J9eg]NR.<)72S>e+:#U56MNM,GH/.c5]=
H45[;D>B3=Hc9_;A#79/X_U_\?UUM_ScJS?8YVD)G_0Mc1Gf@@<QH,&S?#/gS)#.
PgS2f^BLABAF5:MM,+#gYfcPOJ\[dcO/4K,(N^I?J1<4+<NQE/<(e4UQLc_IJFW)
-_O>QUf;0:;QX]Tg[dZ=BZSI1_W3NW2b@[VMBLCKO<XYa:L,C?B)9]WQ13KC\DB5
Je+g_YNTKU).EN6;39IN8G(58#N?aI_0\dVKOA4U_-0=PQ/bge4@AfS\;5TCA;XZ
d=fB;cH_<=60L]X.LUTO?,>F7S[5SNPg+10H?7]b#FC-GLHRXE_2.FI7(94_BGNQ
_N\JXg]T-2\?MJc]L?S<S=<<deDb/)6)gYIIY0[XbfL=E9Y(.42)K4aUb]N4_a,9
4^>3(/OC#T63I;WESZXHB.KF31^L0/?LI/dH)Y6ZJ3,Y@<N,R1d]c8G0,^6?#,6F
QFg@[)GB8M7MJ--&+Y4KDW/#F.Y>-@<_4(>Jd:<3;+L(=A(gY>+[+QPA<\d7>;H/
8UWX+[VPUeRI)J=b,=L[F[^a^/3JNZGTG=b)O(/1dR6E_dMRIH@S9]I:HX6[Jd3b
8A?TGCYDRBYN3S2aWeN[-7I=E8MK3M22K?.=8EY<@QX]>(O0/a/faV5^=&WRR75S
2=ePT+f4:68-0R\H&Me.@cK)Q9cVc_gM/(;B-Me(@9P;D0Z;NY=Hc1fCdA(].:d7
=?#C8J6f818KY])\D+&(:F9SVUc482f.&gX5G?-^2?D=6MFX5&5gFV:>IT50c.b+
NQN]D@J)>I;336R=51LE1PW>//D6N]O@_/EJ./U8:LH5@(TVRV(_6LJVAWV0&dda
AVOW2E+W=CE[^GB0:/EM)5Z>Y6Y?QL+^-Hb>WTB]A]2N_ON.bJ4J>R.C#(]/H9&O
=8?();^860Y4bg^0;dO?gN:DC[HQX.>G_0NJ-<_C[[-0SG5K6e1_[Z-Y1GceK)[4
#3=B.E)5(&Ygd?I<)]QVC88fUSJ&0b(]U\7K+M&/)^fH0M@KM2N?[b3Mee13[S64
_cd:>1P\Q;+E^,A\8?JO8#<^?F\g385?.4?TBYC&-E-TZ(;5bdE.XY=HV(;N(=^X
+3WG_7&6>f,UL#TEDZO3P8.CORWZT/d,gKPEeO9_DcD>bC6(?@9/L&b+XNN04^,8
12Te1&D#H2?XObY<(LaDRFTEI_(R1@@(ZUGQ<;05V7A(BQ+9TKI/?fMO#@]ZXM[7
Z6=c@G[NGHJZgcK4F9X(@dQ1R6C,EQ9>g4_8/:S</Qd2\B2OX8P>9Y[RV;O4&MH]
c[cf@&1M2OFCOcE8f<0PQ6@>=KW3Tg.?g45@PG/-YS=W^3d>dT=4?EJ.:9>bMK;#
f,gPaA\[42@TVC,+J).>gP=+P,PaS15>+9b3VUX;JVN9PaAa)cF(c9?fW[H:N&?L
RKM+UD\)ID/&.1-<9<5@&NXQ+/c/,fBc)TH(Y<BJ2Q?g;5M[24PORgeNU(0[Q)CR
]A6@(,5M+M9IYbKIS:\b.Y-51/E/d0G6S@_^P/>3VUI/D/[f6>F4U)P9>NP6HP06
R#+\NFH6eZF=f0O-e#[YHc+@@?(bHFFU>?-aXAFeL3@VLEfT<dZ7_KaI=ODe[Fd[
_C\W?IXC8)N5?cV-##:5A&AY(.<7Ua:?Y_XHaM:&,W^)@OC,=d4@&fGQ^HZ&U.BZ
P]9QI[dU)UTO>G9__?S]S\4?.(,;VYdQ;-#RU16UF\_F.)fJM-L?WOY(^XE^V2-(
2b;/A_QP]5Z,d>VP_:94WSCS\JJ)[E9])1[_/.,1a(7Z4IP]BHDb6[RS&,I]gZM7
;U8f:K+<_.-dAAY:HJ&+K4S=M5d.+H2LU(?Q6I-Ka/<GQ^W=gU-RV],]3-C9)TV1
)[S\G/VX8C=.\-K[_H,dQ&WZ;E9P.VIK.Y?O6/-Oe)S<>:a8;g#29WJH]7_E/^6G
f[F_F/.,B]8XEY;D0P=3S)DC[#gaR/IY2b4_egRe<A?V^G]bMfdCe66bO8X-:9[d
4)@6^Hb.KMGH>(_UI,]&KUM;2G4#(4D&<]74#KUDPPbF=/&\AG^;f7bY[JgT?ZLJ
,VH4J7:GaI=c,IA;O:3a.FW,SEa/O)_aAB-cWgY+703Y-__IQ&HIX-T5cO8[5K\@
-3]+PT9CE]\XDYE0UCM[Red[_Z(/(@=LXWKba+V/KWFgI=Q=H2f5+6+,-C\>=H()
Pa96;DSV6I-;JF]GM>b<(D[)LKC<UANgf^5eQCbOM=CCVRc>?KEaUA^\GL=E0^6Q
XACH#aP)M>.-GF=SU3/B)],NN:&Ze;6cIO+AU]M9RRJHA#bY0)G6:&:ed/J7Q05G
TLH(T&e\[cAfeZ=8cFQ9?GYZIOJKQ>;(QPM+PAcNP0)KZZ#THCC#URK&#7HbF)WN
0G9-](e)@GdSG&#2@8dZH-BPFR^[:ca/W]H(GPF,^L#[Ag(WXKa8d)WLIYMIX@K3
C]T,YgAFD[:21_XU&4XU)ZCREU.GX9#[dUBGKIfDH10d.U17:Q2b2U.28FFg0Oa7
\.12HA201#N^QV6>)SHZOK>/@72Y5DVf767D,519GfMQ??7T?b4e\6U4Dfe[\ab)
INA1>bg<-)Z-6GOEPJ/\g+AYO#YP\LQH+MV=>H/T9SZYaf[IWR.6+UPBIJ@DJ9B#
,3J(9Qf1Xb,PZSQCfaHbG4UTTJOOWJR1M8/LTYg]NFYOD]H0f(OQF<=,[VH8BcK0
R1[7eJUE#JSa]ES6BJR=GTC:97B>[CP.LH0KPCUDUYR]2(R-37\9a:F)D#-M16[A
P3\7^dEFYOdKX;EEW^(>ca4:X0+/G2_Bd[].+f4@.a+)^LD-C>Q-7/ON/.HB=HR.
\(/;0X@FAHd=:0JTHSGXc7_S?R;HLMaN/GWJcS=g.&gR8NO83VQ(N=_-S7:;bIB&
SG(@+cZ+CDB[C:fO<4M._cA?Pe-M#&Y[K5b,dgX5[9&U6IUX-VI@bBeSB/JH6/ZG
Qe)HggVAJAVV<-dF#_XOSJ(),0NU@Dca/-+TKHf1W74)a-6]OKZ@T9UF:B#ebU(3
+TIM^W&3JYB64=E7:L;2;P]<R):ac#]5)G+d6,YXKX@>K]R1-Z:FEV[3PQ+<5XCP
4NK81fD]V#E1?FDER,L;3D@TBF03=0;CTKcUeCWR>2Yg@T#6HR+[dN;++#;7/35:
f+c2aS(eC#U8G&bd+I/eLP9T8E^88WXS:)ZZ-Vd.8eJU2,Y:/\C)KBf@X:fg=6;K
DSO8IMDX]HT]C?FTLD+8)EJe-J;ISb?a94O\HJfR>IZ,O<J_;C./OB-e@V9g^[dS
Z,?]&f.X@G_QLgOX+?B,GU.N<=8W1@BTD01e0<.B,YB61WY4944:XM_-&SddY<ZT
&VXKIeJKE,&/.4M?]&+LZFCO@-^+a\GBA[-T:#P^2<8<;0E19NPCX^dBBQRbLN64
8Pe0X&@M:e-T:9XDD,2R5+K+2c(VAV=D5?;8OQBV1T0ZM#-6]b2&Q7.T>A=bUZR?
1O9&H@ZA8SYO)62cS\X^A4dEZ93A[S5g]ZQ;L6E<54eEX@d8AC6f@M;RW@S86#Le
7&J7/.:4)=Od4bQX#6bXV2B]/cf>T?_f6[c\GRDfJ3@CVQRJGDX?6bXB)GZK:cE6
ZXfaKcTE>BYSgZL=&\?Ib)=L?+C^B\g?NQO\T-<0G/FgNV368K[6O_H;F:CCd392
^&;e#_d>N<GX;=4Gc:E^9B<def5R,W67,@bJ/4CJfA6#&4WI0+eAZ42UgLT=Fc)K
c6RZE9.fI]A19#F_@YA:J=Hf,<\eN>d9UA7<8P1/VW]CF6T-=dD<V0)7E?Jb,XQ^
aG/G<a3+9#YZ6)?^;8V7;J&5PP2M57;bFYag<C3,6=4L4JS2.(J.c(-b<VUA,:JX
FD-)DJ5DKL,5Y_P>L&KKOQ^787A/dZ?bUCI7_W#-?BbEX]ZH5,0^;>/eU36b?SN#
BHX[#L7R9-UI=51_@M54\8B@+8<&e/+9V5d<Q6E8P/S88ga2DCKQH>&JR_STEPT4
5,KdH::5D>-4PPGBP_Sb](KL&T-7&Z7<HA2F+)1N1I53GbFg^+-,dU+K8AIdO45F
H@:bZYW[RZXC[?Q0P.H+?12)X6a0:PK&^JYUZRD#)Ae2J:Z6bDVFc3L/gbB5X&]g
=\9LDHYF/+30?CMU.P_C.HP4/F8]-EQ/U8F\)6Z@=B-?TP04I5ZJ-@LeA62V;6,g
-E;4973IF<?;T@+G=&L5N+&N4CG6CTPQ&>KHe-=8EFP=e[]3QP^NZ6)8f#JPMe^;
W<:;SP-(?WHdGD(SW71&b8J9gEIK5/Q-N@I=C\#a[bEOaWb\d<?/c<(X/&]4b,AX
_fXX]I9SNY/]>.8cN<-RBW..D\c8d/e?V8BN4:EKfG?[C(?\FX3WNFf0?cDDSCHI
0Y9V==[DQF-[cAQV,VagC++1]-.HV.&eKD-,4(CYcgd@>5AZA?Nf;0+ZVPX+E4ZK
9[+-<1GTYOb,e\aa9P49Od5?6aLC2a4_e:864+RXLM[bUH&./f?b5eMLS[BH1]5+
U[b&0R6/Md@N.dER/bLX(BQZ,V@WHTFV(S^H>AFA\,B?K>XRK[S4:+M)#&L5Z,XE
K#W:HT?fC_-#0#EX8[XR:aUc>I/D>W(d>XdHIRW4;\>J>.^T;(D9J^7/c5PFGMf>
_7>/UTK89Q3>@Q&IZ+59NdA=+-G)>#&^P_FL1c&5^LUS?==]SaN^bDYL+7W\+CVR
(>8LDXD-0(X:(0H+CX]9IWfY(;X570b-7@=YE+R.HF0S2DA?TU@69bGZ,9I^5Y4.
3;VOX8^N#Z]J-c5/f^6-,;(X<A8D]+(TE1gV#WSQGU<TcBb3NC^Z>R?+E)T#)^Kg
#5bPa[7c0Gf.-DJX:af3Z]XQ(DeX0H.aC[bM4KII8)QHB;#Rg;c[^^23S@56bI(a
WgCdMM9.1Vb:;9GbH8\E)HYFPe1d8+6^deOZP;;HEXLK(H-8,4:UB@\ZI6IEI>6N
Gc,J3g8(2]XFd/4K\XB7N<9T6E8ZP+AS2Q:b2NL2D&gGGBZD,[IPeYb/)&B4f4#@
CBQGIf+Mb3,ZN1SN8?4^)cUO5X0R=&@A&;I\+IU8E)XJ>53XGdW7,X2_2b7/R,KT
5\SePAQ.0&7[K@Y<@Z#+b+^F6Yd<2KY8IfXS5/CY0-99QS@U:674C?9HCRP_1F]_
K72N(?T]N-F5.5B)0YL<Z8NfB;-T<bR=@G,H(2:?-.ZGYPMgaIgGK-eFg47[<]@B
+[MN5VfE]GWce+ZT-T1e)TDA(.a=71MC/];7ZIc2X6a5U7^-P66[]3\VD)6EA^?N
b5P6W96cEBI?dIPT5MJ(S5R#+#JD&e@G#c]V-L#I1)(J/S=2eZ.6TE.HN6c6Fa]C
[-E^N@B]+;5SR.=C:_D7ec]a/=MP3(OG+Y/HL5cMc3^>I&<g5X3=T-E.P&\TL_Ea
8,IIEUAR:@YGQ-CHLPdFP4F7N+10(ca.]J=5<O3<MXQS>40IMZgeRb?OW8UgRF,Z
##aZ=a0DL-KV].RRQ70\Le#@)ZZW:SA9O)]T8agXI(R\+W51HO@H@B6);?]KWU[_
6A+PHMFI,@1+J=ZW00NQ2#?-.\D+>S:CgaV()8JY](3;3XHc6PK_5,5OG&aS]V^B
>2E]VFX&SL(;&\H3,H04I)H<Xad0,AW@>__bcZ0W/@@LX=O:AcU<JP7SU^:_.F\a
/CeEZK?TKICHT,H0JbH3>KfY[_?7UOa6[I43_03f5bQ,J<^60<D1_0)]+D.a,,9<
WYH)6U?a)KW8D]<EEXT-.<[Y35KRb+2SJa^RWVJ8.):gE^/WGRGC.X5Q#=3OGb/C
DQ<)/\P2fb]4[ZCE^Z-C=QY5^HMR=N;B\GKSC+[W[Q(R^>W34J345);b@dN(Q3[/
NUH:;6WE>_.^OaEQ^N(@E4:NaG0?Z=:We@&#U=c;.4T#Sa)A-\>5Ma:fOK_Pf2+U
f.W=@#UNWWT9;g+X30ZM8?1K9-Y=gQJ[WIR#S-fQ(DMPVbd6&.6?MObYS=DHPOP_
bXNTb2?B>^[LKK]dO7T#TFHMJ<gC=.YR@(f>LPfXX]K^#N]2S6;bbd\H(2ac7MDW
UVWS0&Gg@aQ<(@[U,NB4LJ/3KMbfD)LUK60.a1KY]F^^:CRKG/<)JE6T/IWXBLe<
F[cTS>OE))]Q@NOU_<&ZH4gCHN52:^f:,(b<P?gFY;2N7<H#:aOJ?JAD][T57;33
d6TIK&=[E</Z-_DdK8f[WLE>dbTTK+eP0@3a>aBRE\We/QM+,L:4CS(eJEggP\Mc
ebMFROG./MDa9&eK54Bf)7H:bPC[b?cV-SV(;O&QQN_-9\=GUCNAQ4[IgUa6PKJR
L;FVGCYC^NZc,GLLW@=WU(9];f2F]-f^L3[QNWR;TfAAN[:2Tf@5U[a>&A2)3^g,
0ged_:b3>c&DXNcRZU,6M;a2a/&e0g./)>^)+KfA53Z6OR.]IdKbfd^b;;Z;7P\=
L=@@RgaQf=/ZB/4b79FBd0TE1@<M.U(&3<H6R.QE0O5@JAe_CP(/Q^JfFB<GAU,S
]b-HJ=:OE5+3B,g/WLCDA##HJJfK\@PKJ=E?W2<]:-Ld0PNW@KC\bR/a:(UO#_/R
<DaIaJG:])[:03NQFL3=g@eSX:R5EC64,?IVBO^/gDgHNVd,V9CbGD7KMZ\GX94T
LYBXKdE3P-D(ZXSJ/9@864]==QD)I65XY=c/_7XNP8cF8[3=a(WeS9FY>^?8);D:
.20SC;(3JQUa:SR3.S<<B3.[DSgadeQ<.G/3C<43g@_GR/b9DPICPBcMX^4M)7K/
7_A(H882cX]/AQ0KQBgYG(gM2J,4TH8XaK<;O-LeAb_d>,6CceA5e^c0UH?.\5d>
/0gCT&UZK?Q=I:G#V^6c0N.7ZdA=Y4=9<W_NN?>5F.43(f>..OV_HeUQKb3BOcZX
WPNTN^a2MP_HV6N=0/PJ8]N[?/@H1B(QLb2&\T:NH/f/[@_@a/:/_N#YfX\>TD(F
>JUMMEfI<2;F)F1+-:-]Z;8?eU-00-\4^_]bA6HSE:A(e(YG^c]a0\A655EULf-Y
1?I+fS/1_V?W@,J4Q:N#,:dLCP+35e9C0U&:F;9[cFP(aDUQN@_J\O5+I0&eJ^+F
P[.Q2)X?#EX4HR94_KLFSP:ed;Q;3A8/V97^>7b_<.,(.7,2f?<4AeDGC0NCW(_(
DX,?8>,D\OAR2RSE&c46P3KdZP<4RYHBD,#A9COB#KF;a=Uf8=&QbLPff2Q,79A_
05-b_HH3Z&R-8bD4,ZB8H=67f)a+YQX4&4^,e3]CD@?[ee8[6-OAI+@Z.I/.Y/DM
N9Ve0.Z,b(R()2W>)-d^D#Y70>/#Q>6?;>PWK7<8__H:&NDP,BA;a&HJ7?L^6[f8
W/[Rg,]3OTMK64+JP?1S\PM0G\W;J#\B[5@J[A52PKIS/>I-\DC-M7IdgY4f\#YS
cEMFPeU;#5)/e_0FfR1Vf4CKd^8&C;&W7;#8:(W1E8YEDU93.QF:R0[Y,R)6N;VB
;E8H+M.[P+#<KY^EKcPcH>4Z[\BC>/SP78F>^1e6DZC<^XC&]6d.1Y;X+dYZIS-H
)dTDCTG-FE>B2#B]Xf8,VSI_<^>&(c>:3c[12dO+(B6cQeaB+#J\=OYZ#?>P5DEW
4AMZ8^(,YC0TKN(H.a[@Q&M):VVT2,27_(5BNI#:&bE6.Z3]?bX:=]e:YDB\0Z>+
T^<?bNdgaEE&@\WbRcAM5@O&PQCG,\;2f2/VY\FbcM/_9XSH6R]?:A8EaZ]R)DZV
,ScD/YCIg-bg);eUOBKPI-CJZ&80=N62#7_^+DTR(K6YYeB6e1QK1YJ)H+751a:f
.KWW6cG//+03,c[2=,G/GRU57efFS\(MN2b>:)@JJE9CX9c<&g3CPe#DYT\V_&[B
6MZaQZONSXM:N;\#]S[V;L-6aOVKHG(1YRBTgAag1RfYC-7:+V6Y8&:[O>XASf8e
.<>+,>V#HHD1.;_OfD=#F]-\Q<VObCQa:8X,W^W6@CT=F;QQAYCK0(5D0O;aURRF
ZZOU3[&,19Y8<db-.C+P\\>B,eZf2?)].f9<ZcWQ:C^V33gUW?N=^)cP;>B[D0._
^JE8<]85)aQ)HR>E_JQVePMf.05]VM?:AR[)\aI>0e_<X0Z>@.PPaTMVXFJ31+LK
L+,V+WSbDL1>f]59HdMC:3c.RE^B+\&3U^57?4O>.g<:XW#cX,;W]aH-EGS_=3T&
2cI,ga=_9)AR_A9CTd(_.+09\Vg7&T1@_0E9(PS=dKf+9-@)UJKagYJd0.,R(5I&
+F4A\@@ZUMGX-.BGR)caGFYB:@ABD8VW7<P\P4W9(YaF>Wa#768MC#e;KG_J3c):
#@AbW3DCd/&b9eLJdIW?g&&#JPRXJ8;C4W<9>#9I,.CQDd,-YaSAX<O_YG8?a3-I
.0WP2CQI:f&J5IS#TaM\]5_Y?A4.fa8P8B[@7P7T8/GJ9YG]7T6>AJ2ScM-VBY>/
VH;[@5_S[WN_F(F38_KWd,7@2,4K1U8MSLU]4+>3N/V:6GU2&BPBD2e4&DRa\e[Q
F_AU_9BSG[_Y#SNe,3Y+AZ6J/dQ01GXeM0,XL3W5DGa8b#A?[0CG.fZJX>B)2JH]
2cK+C;,JE[?1]5]=dN.;fgO:_3e(=[VR@IOg[ST7g2<Z-I;/f31G4H<;C\6A/N\e
J9Ea)a,1P2BZ+3KP?abU<NP<=ZP,a0X)^K8/#AP5F1BYF5Iba@:MYKFH78TKF,L1
,_+H[aMgVD2Y+YOO]WBQ5TUCdJ9H51H(2]C=_?>-_D\//GKK>RAD35,AENTYe?Z1
TOEe3GDSA9&K(B]_4/OMd\0EAAW4VX)02R+59LZ)GLKL5?fOEUSUdKI.]^0,QRI[
2N;eWX7,F/+R86Q&fbdSXDRNMaC^eKf.3X(L#W_?f:2+B+\SUa;TO7eU8d1J<4U6
,MDO#C2fK&L_TQ(J9[8;?4V[+>Wf[\4;757<W/?QL7TG)W?+]9A?J-X0<GGMg8^:
Z.IZJU4<LG0dZ1a&,G5SP;X<JNUfOW-49O-R>RF#REZW2,aPJ_ER4H#QORgc?WXb
BC7[eH9=5J@XU++RW4gNfFX;CUF2GEPN#+V,M_3UXQ#05^.9I-N)K>N7.A&,=f)8
eI-@0QRHfU9]f.0H5\OG4:<Z2E^[aAB.aE-aA]/<K_Ad]^O4gAYD?#FX,+YVO2Se
O1e#2bK:_gJCCG8bfYa9d+9:_N+Ab826_E:-^W=KUgHLP0]5994g.WgT[6O\-,Oa
d7(f^(GV,g-)bOe::NO+B29O>G0UGRWIP&-]Z83-RX,CN5^Z\^82gAaBJ6A,0TV-
9/Na&,CT^aZcaTc9OP>+C.a3cgN4c-NG=2@EI(eT]840GSEP5<a/I=XbR&ZMX_:[
fb^S-4_AG#6Id<gLUg-PW?5Qe>0e.gRO-Ce[7g;J\aD:=B260Z0VDgbN?V3W+@E?
R2SGF7YDLfKB#6T+CE-/4WQ?ZN,OK?\2-U3.L?+\KE7JX\S,:_OFc,B+@W+Qa4TV
e[H\IH4P-gD/#[]Yb\N]7gfEQPYLKWVd(K,95>,072N6COR0-Y,\N75fbT3d[TFE
;6W9HM>>P@@X/Zdef-.Z&-;5#X>>MH4=L],2^SUc,;SAOGWHP;/=O)77_&>,I9@/
5#1#Z7;9C2/1V^2c3&V:9-,3cLRMPf26b+(14L7\@Q5R-<dZ>S4]Ed[\e[6>P()e
67]<VI]8/@Re0Ad51V_?f(S7O@X6=LdW=[(gHLX\B[>\-Uf(Z(;H06A8.bgFcP8S
XIa=GD?=-R[b\]#:3(_KWO)F3AV6]^E\_XXV>N;GY.(7RTW<+INd4e:X=(_XY>aU
R:<MgG;@E:WYL=c;1gfB(4:Tc.O&X,_2609[gLV08Pd/-[9^bK9CS((NEKDU=ON2
6Af-BC0_aBfX/L#GHM+L.],</9[EcdaOF1cK\Ac<_\;I-H6#].UfK6BE.\^KGgMN
2Fc]0fZ>=U]VHRXAUf\__[N#2@:aOV\KEY^XQC0U5RT2//3,g>Qf7eTba7ENbR)N
CXK7)#=/.CJF/LS-O9.>BQP-ScXg-N@\81,\I4#.[3ML6H9R(P:/gI1Q/YT)/a,B
9cTGB&YeP+6&<4/X-&T>#CLP;(5T_4</0@^))0;H^1MN+WO6Yf3&,,Ig^6&3\MO<
2Sec,E2/E&dLR&N>H&gac-^R(JFHA4>YE^9562XKL\(GIgZJEgK6^+Zb@=O_a,@>
6O.4^S1]6U;\CCE^IX\1L-HE4a5,ZF.OB<6Z-3X.L&(:WLF;B+3Q80X5]YERU?A?
+E+Ee:RB.Aa-VD=W::>bC[.;YT(LK<F==QX](0P#EF=>T:ZOC9=8X>&V;73W[AG/
L:4,W5PRQ/(:#MV;M;QL-Z(/IeZRE:,0AA<VN^Jg+R<;Y1\RR:>B:W^&d7^-^AOH
4+4f#P1?6,]T-DP_d0&LGL7&340DWXa]>8Ia=1D[67/Y)0W8:)#P]R9MS=)-C[8P
R9@W_1&Pac45(\G]:U/g4B/3>O9#\3FgWO6Cb#:eB.TWXY.a)O5?/CK^E+/QMZ+7
1bJ)\3cR]Z34:[T<)B,-6^<F1SYU->7/]I__]2V@PB#gPgcN3G,H,RgQ=>]]LTM4
H.)<7f>O?\[I//AKb0QdRT#1]I(cK?-V9I(B^3,T^LCALCd?\,Y?#2]ZgHXIP\UZ
[,IMe(U=F;L<3-^J0)N-?6SB;LM\<HN5B2B:EU4gf)>+JMPL@P1;QWO(\(09+VHU
)(\f;@5_@NBC8T&:G8&##QQZ+=DP.RdA;EI=UYZ/KWTAQ;@(DP,f,R;.b/e8Q<f+
Z?I^ET?c?B3MHcNQ)/#0Pd^6QF4:EZg[#=&D?XH9>X=.a/eC.>Y\<O8J:+EQPaGg
G,TLEA>+2Fa)[Ue,R8E:eQXR\,J=1;4OWU.QO4+Xgd7T73B[@,[MBd\8:PP^O(.K
L0>OR#gX&U<QC=fD+E2F0I.J.JH,F-[Z9Kb:^,U0+E.XL/8AZ:4)6C0:-&0IMg)2
T8?.+GZIWT&-a?]-5\6F]WTa6SO_I++6C]LE:\YK6Ed+.R9_6=0Tf>(=W;gN0PW&
^LJ]28FHGcXH-AP8a].KPSJa;>@D(?#ISe)&])/@R6G)<]M-^Q^6SJbV1ZS?a,_N
6NET;G[46gb5P<J_:cg&6?bB-G.TWgE@E=@F)7Kc5JYIAcQWAH:LbJM,U5?&-7/#
6GCG.PDaRQa<KgM@Udc2K;3^/:QMNRC)Pf^:U5D#BD(NO0eIFL;@SS(@R45WQ0[-
X2H7J>g2+DgJE0K=:NeFKL3Z^QAC:::O62:CXJL9@950WWVAI-d]U57#:@Lf^&fC
62-K=0W.7,8B+WX9XFDEC?3H35CfD1C,F#G>2eJ5</IVdT?.5CK:SE3JH6)3d(<d
Z\f4bSOC(.WQa[6?KJUCJ9^;^.TZS&/?]b^d7dY.eL+1U3UP9<Y2[Z7RG4Cbd0NP
)R3[]C@38[d3W2^N@\H3@GCbL)]&V&4faS60QD1c4S^b1:+:^I&HAcg<5=:<_1@b
;;V09\JQ&2FbOQ?R)UX1NNIcIT8?I/IbG\4D?IE5T7F\_:NRXcT0L9=c/4U-<1=a
262MfGXYEJ@-edFM+@KTPYbVNTED>S>Jc-XVM7&1bU=e6NeX:W4U@YBbT_<CdW+c
Q=;/3=SUFX;Sb+;A?S7#gBY2<35C=>OabQ+bV_T8N6TOAcJ&6RTbAHRYUX/?P?g,
.<e=ZU&BKC#)IJbId1eKX9]>U3.,K[O7?<97_Q6\]<K(PYF0g>FK@R3?W_6H>)Wf
cV16+XA7+VG#3N=4Z=_;]]D-N[Q8H@/H?(DM;F?0X2]?WW_d0JW/FY]W]>T97=@N
cQ(-GBIcHeg/LE_)-<4OM.@1H6-]1O<dZD=TL(>/WT.M1+X:bNVH3.SCM/I5X,4D
_N2PVF9O+?<4c21UB6OQ#;2gO2W6]_D]WIATC-&=SW?B[OE]Re44=:WLb:B:LUYT
V,G^8H+XRV=3/@>4CUQ#&..WgNW-&eZHX2^CO]TWL+IFO&N>U\eC[@g:IOBb=2X.
,P/KOKZF)KU#BN1[B,BF4gD]08Z9T)EZWMVLFg03X<+AcR>Vb#+.7=d[F)dDT6a]
HfF@;eM-g@]Xb@J)]@b:BGaO1<_9O]G@6CXfYNIM++fA/BJ^YHa\#CLd?#Ga;edg
bAc\c+B;180&aS2g-G-AB37<a(H(V?-2b4?+ST#U4/HR+>3@dTfb=#Ed37]7G:3X
f\Vg4dUE64bd4@[MT6==J_aP^9Jb>DZd#_90.&M.CEb]c)JfQ,=2P@9/E.[7VOOC
,;^D-,LgV7/9=\db6PD4<CV0+=HZA1O&-1#Na]\2g+bJ4;D>?:1.KFdV/<GO.3R[
&L3Y6F>]Ka,gTH+XaU:Eg6D[d#P^92])L(BL3H0Z,dMe5?41>5<L:S7Rd+^2V@3T
1Kgf/<<91,#+RRS@H#&?UD80A<JC[KDd(6R0T=UR[8c]_Y\N9OTE&KJ>,EF=VC#+
IN:&QMN,N,UCbC@LO-&&OXKdJW9P>g>[J-fOf(<QWR/H2Ed_Xfd9+W<40L[(.HZ1
Kf0,(F[#(\N3F,,G66FU6>UXA+8-+)?GK^=0ZWHaV-60JaRR4+RG)?2aB.+G1CbN
<^NfAY8CP&EW^826Jf/48f3#N0MU;?;/QD^Nd>3IM^YQ@]2S_&&2]=]8)c5WecbK
b_LYaQeTMgbBIWT.e8cG4/aDBQI-WT-E0bH6G,@1g,^)F#))P#B;gfC=4^4>Y]E.
+I_^]TIbagD#@;^@-MZ:JKKE)SQ9Ebaga(H;WG0_M(L>[g^ABD+?F65T9c500.G-
L4U8(c3U11;-S1gaF(X6C2^9/5B7R2\aALSeM^ZL87JR_gW\9<HAe>&TBd94P39:
,,GF:J&FcBfg+05;SJ,(PS/1M>/FeA8LIL2/3(OF_Y-M<9];:cMZ#CG<3)^MX@N2
H_Xd0PPNgW?FV)NIf9MH>,(OV1=5R>Q4O?Ofa^NZ;VV@PgUeUca9R#>4U2WLA@2U
^JNIf.32fQ7bUV):AJ^[]5aDDAffURGN<EFDH.@b4#:eEH6<A63N1J_ZP&LW=5-S
Tg;WXC>GG^YE_:?RN^4H8,K:>8VB1c^OD+cHUg05aM2ZJOP8,B)HD)Z7f4^Pg#dc
12.Q\=3:X-+K7?(WMcK(=ET>IEV2K;d3M5?\/RG3g>\&1?V\Y7A24V;g^D^dT;?6
SPHU.:96_-bTH<\@H0LcF-EJ8P_F26(T9>3=ca.;VF,>,cL>Rc?O=b>fU#K&Rb=X
Ade1KU4PCGB>):-L3g(=_3)VCT@_EH/KFD9@]_&+[:_P[=-[/K(\S4FVAB;A,B[N
G#&V@>GZ(ABRA#?cb=[.Yf,U>0+?P:EZC.agIIGbA>P2dPc=T(Z(94SXP6(24&IW
Ta_M2+KaQ=^;Z3@&4Q^6NfE?Z?8V@5eQfZ-O0?RaS]WKJ_^YdL_<K?E:E[/W_H_e
/#@_eDKbV92GP/<3E9A@eCe80K?e1);[;-NUJ-EEJ2>.cbN:NH^-PN2/P^LAT6RB
Fbc9)HF,0gZ>Y<S((U)CA[GIL;>F;;7/(+Pc#LYD/,d<WO5P6EEe9a<(;-_-8GZ4
=LW9[gWQG2d9IG6[WbUY3gRaGQV/e;?3XZ7J/V8F-Od0,XBWaL(-A]3NTY-JU7Wc
(7#DGTg-)^W3b2?5O.GdZ&N^9VA40P6^F.D+Fe+8,C3>JKAdeXZP7[E3Z:6UcK#Y
[VV<-LN17Na7<K:57Vc4cLd]8J)8eb]-(fS+GVO@Tf=3X3Led80TFO4K(B3b@E:,
A9P,f[/#M>gcQD6c+QXT,>RPZ&BaGS)C?efXL.LWKO+__0T)a^B&#d.AT=f1,R<d
UeB]^S[G=)GH?0[YdKA@4c:4F9MK&_-,H+#)JO+)@V5R3d,7TN-2I8#).QggT?eE
[6<U=]5:WKNXR1b9C&7G\I8_+J_;&L:\X35^FCc4,#aeUIYODY5[TZEA2@b;J^aV
f^@@6VSE:9Zg479EcdUP4U[LEdYe?AdJV9_;1dUR)A4I>ga)1cLAVZ5791)aM3UF
[TO9WUFL/McJ=;D([.HIA70b,#N8,6b]M)O=2[TM+PV<0.cfgF9K/a\91;9\AE7U
U6Jd1+2:dDKMVXbE32L\[E660@[P.PG3_L;FST6<H+NSSC>LDgT,YX86(W)eP]BN
O(ZBZ<IK(3R1HVK)UH)3NN@b@]O(gXLKEf4V9#0V<7X?6<=G52J:ER(60Y\U6EGG
e,ZZR3UK_^ZY8X,G0[bI1DL(1@J<LP<IH3fP_gH@)3UDJ2e?5<;b#?3bFbZK:=g@
7_EF791LLeQ-4EgS#(QB_;?X)ePIcM&FQ6@</+^7:T7gEO,LV?HcSPb@OaIPNFUf
OQJd-P)X\/+4U3;UNA>J?C@Y[=J>ScAb^#cFFGKQ;[gc8Q)9M-O-NHe\a8HA(C8U
+^IH0C(/E)G>Zg@Q^]eTB92dAI.U;3eN3##V.XY1)_[K&,P^^MGYVCd=3I3^AFb@
-Z[4D?H.NN#(1bUF:5V-Qa@gS9J3g(bD171FC[B84f@Dd(/#[0gZD;g3;cSMQgS@
)&@;\/Bg;bf8Q+&MTH9G:KIB0KF]E]1^0+OR9Z,R8)Vc0Ta1V43,#&5>I5._6HQ,
.R1:dAcbBbMG93UaO3V66R3SZSaf^XLG-)2X^C2]b;<_GXfYFf;g=,3.>;]e:>=)
0UM1V&G7QHO69aU#)4@Q(ga-:=/Y(5ZL/.@DeEJEf28Eg&F>9\A292OR+]X_RNcH
O+H=]O_,N;91D&X[8.fMfQ?9[HJ@9a^@-b1=U8e0>fBDC:?:^^M;^+4L2-Y[B4aJ
<=,\7-O:g4TLP?6B=?S\(d?g9\:,)CMGVB2G0<)2_F?C/&.6NV[P18Y]WQ0a/3.Y
Q394ACR7K9B4Gc6D?c04#gO@798]::Kd(0AWYIfRbAAD-Y8I)079Ag?Z:MPX3T2;
]M\cc(d[abSH21SFMN5#GS)GKX8Yg.>&,BXTU+_W]J4)cB7YHF0GD4A7EQKb]Z=J
I2I>AQe7BI:VaATg6+&Cb_2QDXGFUF[6b5SB>MB=[2H.a&-X\FZ^:D6EWcL0;]fL
CIG>]HfTVRR7>[UTb1-D&9&d.HQXB26L8X]<]A<;4\&4P>^NAaBf,#>1OHMZ)C-3
GL7@e+D?&).:ag+c+C9,[==_XQNA.7c_Db57M#ZA]B>2[LKGcSc&RJ(GP448[AVN
gP]:0672Q>]21Z4LfRB<#7,LOD4_Y]ZLXMNXF9G3d].T0QM]>/X/P5LXW=Y2F,_R
RTQY0H8PCb3Zb[_3:IJ5P4KQ_Z\(T>:748G4(0,2cfB76)0=CKKg]^B=TTefOSU8
dR33=8<5DJF6\IC/6VGacZ>0JW1VMB)7.)d?f^]LKI<f[>>IANKgVb2G2_G&a(@^
-WNf/MY4f7TCACfE=4__e@MPZ8)7b0#/09YY^_9#dNd]Z9H+NY(X;&JDDG=fB)cG
YY:Y2+A4O613+;2_fe81[5fY:F_5LDT@TfG^Fa+bNIW_5VESAa<@a)A4K],B#6.,
0]:)&d?,&PUWO@_KcJe.-g:@LT9HX=bEJETTc/0fMMS>KdUTb66eKNMT8K[L(3GO
MG6AGX0[>P/XdJ,B&Z5bb0R<g3OI-W9HaR(KR3GbQ,<cc8/UGK_F\L@W-0D,;Q6W
We3(SJeTO/_U3E\74A2@A[7)2J/O.A22G8bE+SIR3\Q_8g66E/-;(,XEgW.4TJ+I
OGNNc_NVeZWgE0Z-bLO@T)\XP=c#;ZE>cYHM35)/=.<;cIO,+G\ZRA]@FR3VO8Vf
\;J2,KC#IR&4=3fFaa8=6>0?OB=SD&=#9GbZO,0XE3B&@(<BR?fcUT(cW:LG&@/^
8dbK-/:I2Ag9(+<30;8e),YCA1AQBBe8PZM0XYYNY._H]cMON.F[-U_U]8V\]5^L
NH2JcFN4Cg4ZdDQ3D=#]/HNW-;64dH>9]&P3Ed5JT\?5^@FBF?[4ILDW#PZ[URA6
JS&-[cKGHMWJ;0HIC,_FEMd\?cBY,R9Lc;T>(:YIb_b]ZJXUK&f].g(+2&FNB<fM
0>-LKO5Fd]@dUO5.+PWBcRG;V8?c1KS-g3KL^,K[B-O]FHJ=c4:)R\XQd;WFO/,f
E8\NJeT5fTC=>BK>]->Kf-^1E0\55U8g=O-8;1(bGF]VUfZcVU(<X]M+(>,?X1T4
gegaJ(2]H)=gZb3DS\\AX+3e,Tg5KM4?RVQFgKfB)OY+ScQU/bT8O-bP-AdS69N7
b5I^WPYM@BWQ7dF5X-O01/[&IT1JGLF;^c73,/^WN[??c7]SAOaG)_5=(Y9a6^);
7VBO<D+L#M+S27=5)0>/QW5IOAf[BJ_QD[?#?Sd=<6D3<L70A6?4JgcR&AeDgCG0
^&WbH1,dKVNc-9L6[d,1-]LJa3_54S^HLc\:DIbM.XXO\bYW?C>eQB,35&b/-)6@
;.)&Q2c:7M\AdS&]46^1)@A:f4,4GPSRA^eFf,1^[JBDFZXK16H_T1P@KH9XO\P@
8]^J(8-?\Ne0#1Z2G_,ASY_9[_XQKL/._:1T/e/TSF8]283)EH>[XD,)DKX+]Jd-
&TfYR0P2CG2B(V9@[XZ2>LU1Id>(&O^HD,^^gf1MC/EPNUBJTG?+7RY;PJ?]6,W?
,:+\D.5TZDI,(9D4eNX:g9AJV@)2&_J4E@VL=)2_bTRPG;Dc^,=&;JK4EKW.2b>_
(@0S4PfR]_WOUBg.)d@eC@,9+5691)Q-H,,)MA45\Zf5C9GW.RN]\Cc/A6\eG)<Y
P@NQ],^4CZF@B.bZ(X,]SgQ^3;;#29Y;>H[IPOBaUT>cY;?DVCDM,&(<NEN8H4,D
UeFb+:Vc\XS]EAc=V;bB/MeH[ZFcT?E5FEG?6cEB3(Z&YSeN<Vd[4?e/NfHBD[;L
a9g(bRJ2B.T[V:MF+_GB5Z&11Y^8Yd7=^)B-D#&U+X:=B/G@T=:=GgHG&E(H54Z[
4P\(HbIA)EREYJ87&/_:_aIM1GOJNg9UaC:3ccJR.,_7P&O2IDd,<,\YI#LKV1\Q
3[d825#KFEadT-7WRIaX;G,[?M\HLS=dLeMC=+-6>Vg1QP?T<6O+9[-;I7/E>3eM
d:.Wc)GBDg8].VH6@6[&gYB]5a#8RQb&7H6\_G(=;U,+.W(@]M\MS)LDGF-TZC,:
Pb7.NL.Kd9/Ea1U+H8^1^]3]10,F2&+.3O_LeG,2Z-1<V:8D<;1>e=2W-4d^X.OM
30VABc6g:6:1=c<d_/3[;a9aU>.ANV09EZAHd8L_]2#dR8B2HDe)42W>6/A896YL
Z0UN83\)T&8:4(M:N?3\TCH:ec3&#g/91f-F[OYKI/X+8bgNQf/E51g(e+0>(b;,
&Z8^LF+\;=B4LQ9bQ(Z@D(RSdXU9T;ZDXPY]Xf=2&eM7&\I9W4)BSR^52U,K_-9c
e0e5MJ9)b@c9&M2OOW:<X5.6[8I_0G52c1)@9\c^;J\Pb1c6&)8\2163A1<F,#Z2
@78^(eV.3.TA(8VT[acC7/\863NL,>N4[N:=Ma&F^^Z/HO]d[;Db-dM<#L3>NCJI
L(9S[.J)>T&78S6c.RQUQb1TL<Z#3S\^6F]?X#\02RG:GLgaDeXJK>+d:V2#)4Gf
BUMeUU7Y@JaO>ET6fI_AMW]\T^E29QcFcI93Q#OZ;O&1PWSg6a;QGdD)(5dVaB0R
)GUCcW5O5M6)MU5CZ_4WH:0:@UY>bfcBfA;b)TO<T4=2J4c-9bMJX@Le<^CUQV)b
V:V&(GUQT@TX6C7R;g,/b\]&UagWfH4E3N(Q?gDc&6+VLN):f^OEKUa]X<\&7WS1
&&@f_P72-&K+&+TdO:?LLD4VdTG>6X>]KIeBM&9]:M^gMWQ<3K8O-]===CIEV>.U
d2IMSc>-AP&+,$
`endprotected
  

`protected
1JVHF\Ig_)e>9+8CTILY(-NB.SJDNP+M.G7\L9ZL#B+GNG43TJ,4+)/JS,P/Q\TT
9JHW17&[?6b>-$
`endprotected

//vcs_vip_protect
`protected
;Lg_;11AWBIFA&T9[M/^KEXT8,,YH?U#9aXGD(L3MT&4276D06166(SMV#8S5WTC
aH#AE?\WC]K67e\J[09Zb2U>bPdXMca+XQBO=Z_D;F_+feT2VSU=fNX)TMGIWK6P
-Q3]f,CBN>9eO-C@4=KJG0V]Q?6M@^+D@(_TO^V?89;fRN^;#7/>PK-N3A7D_^0G
YBf5__;#4KS3OS(=\GOaAG;+S7\PB(0NF_4,MU_OfKW3_WaR)@8,U1-\gO5)5(U+
3Ae/QAOd]>=T0_IL=,7H]&B\?gIR#+40:OdO--:6\#/^CN.6P9-/IKdEg)5?A]6]
A]30M-PP<a<^H\9PD?(#^cf_)L>ST_WGLH6Y_(ULART:K)ac^Vd71:b<<gQb68UV
VU4>31?&a<&8d9XI<688(/EU2OT6IQ(CFe-]>H0Redb<U?A4)#09:=IdZARIXYT:
J5YfFDQM<96cG0J-\BYd@;O?DYC?+4:ObDc0W6<KGLWMV;D=bQ/KQ;R,I-CScg/4
ZZFN\7^bad60bA>KaWfQ1aWZRY,6@-]6#9XeTONO__KdH(HC<]T^>KWER_cGdFTC
)cR_L=E4S+B(d9^EUc@8/J<K/59@C<WP;U2beYCaUgS9NVBF94M&\bf6RFE6TbaY
+A^T7<:;TW(gGL2&P(,G/V)]480IR@)e(e&.X[MMDI^748K#NQ^32_a<WC692]LN
HXZL5_Z>gd/V_98fadB>6[@cD.5XbI+<@=@14Q_VeP^e#3eGTF<Y=g4OY^#>WcPB
0@,J8:8Y8GBYP-U=2[@cg94O3DA(FM14J/#bN;K8?7g+]5F85^GTA9OJ8;(X2ZNK
R[(+FcP+U6M7,d5S)E7Yc7U^T.#+NC;A+gCaV7_&N^@9W&6^Q_Z=&OXXc5NcK:,B
9b.T\7C/.D#S4Le/NJ,7\&RIP^Z4>]\,+=5::IIKDe]1fIF?F=W,F_FL.d<5d1:R
D7c<JI@]\5J#]/MTV:X7R^-M6QQNgQY46efM^ddC[]gM(,T?HDEV(-((cc:eO6fN
JE,6D\1^^E.AW>/JT\ff7H;TUM?@c\XNg1a)a&QacM^RM8.PT5FP[9Q;H&MY8Z<3
C#WVDU[\/e&0_1(>]BSYF\VN5;CAb7=aJ98VOWaQY#M;KRBVD0aYeea<+?&DYee[
N952A?M:FP3CJHJP<aW_0^6&a-.daIJ>A1OSfU>O\MeNE@9FU)b=A.M-aB#QS]AP
f;QH)d4:8F-,>eO+ZM=E.<E9S7XO/J00X5(\^aWPaZ<8OcS/YR>HHUTL[F7>X=UL
,6)V.78b307ZRT\F_N]31Ub)-A:D_AXc^Jf/9AQ)#FW[90QP?\QXfMW(4:&E(/R=
Q01P/3d\:5DZ(_M:EKA1TX24#MOeY8/.>(b1_L1Y@23AZ@aU3cFD,L[DA0bM._DB
;8OA5d8Q@ONZZcOFA5X_\,GY;a/8_O4I5_@[U&[c_OW>:PU98IDEC.3aB6d&U147
BA?ZM6C5TTN2D9#e:T+@4@9e;PCSg6f@@Z2,DP,@BaG\XS;^,c30EC\Qg1QND.H1
TT<4U;191[ALJNF3O[MV0QaG+XBY1Ud:Qg6&9\H.Q#f/Q);@@>7A8R&90MT#?UIG
U2L#:Of#&Va6aVOfc7#CSKNFI;S_#T5TA3:FEH,/cU/+/Z7&42JEb8ddDf5\\g(c
cWgVT6/<Z\S\13WF(KAd<b2Q_)Cb/5=&BD\-#1&_dXEM4Ic).3H6=:SfN(c_4AaK
7Cg:DAB/T966B\Ba#9ZY2)bRcO:W&>RJ6.fM5=g>+LYD7YFW?7e2+GB@YO/7NU[c
Z+/AWHT@AT9Bc]<RH7+/;<V5(.V3F@]O[X\:CZ0[#HOR]cfT_8#X>aeN46ZYaK_^
bE0Pa/Y27+8:M8(dQ.<Y;8):<3S/D,]PX29]MUS^9[C[U]E:E1?3Eb,W@),[4:RM
JI&-<=e+HG>Y7LJQL\@H)7Jgd7V+QS8V1^<Q;b1@N<;T6FY#_9<2-d[TH7eEY02d
UgU_-K;NED@TNT7AcZ+T6;#[>KfK#]@=W2ZTX3K)@CP3G)LegX>).I:WJ+_Y#P=^
B^?dUg_N6LEZff8XL^/5?;<SR44)Y]c(<^Z90ZOSdPeMF(NBK;[_e&/392dO8O]G
O.JEHG?T6O:?NJ:<:JX@;2F0JfW6-#)X_77DBYd<LaDQ2@5RIRO.&C#FL(@@[>37
CgT._B984DF:MB5ZUCM1(Q7O.EA2b;TQcB>J1K5,[G3B??\4[31]DMHIQO&HX<Q\
eK][DL9PgFUYJRG,e(B8P#1_KfOGJCI5L^L#NY<M^EK^DbG<@=Aa;I1U<K>D+]PE
2&V1OX4)0-F>YQ=8Ea2^@G_^N+](>e/O@;QIG;Y-8:I.?RP\:OUMV@402Q;[eg3E
_B8;5Z>&Jfdd@)@QX_J/H9I;RTa1Q@.R(T-TWFAc^^,<C[Z+:Ca]:c3]B-KYKOQT
DdccV=3=+FN+Z;.<-<-Bg<IOI1HWL7-K-4\?6Q#>-bJTfBH&40361\)17gH;e(&S
FE=JLGfIBM5BKD8]X_Fg\9A(-M/DaPG0J<Mf=/Y>DJ]<M>?_U3I.,&NF#FJ+\PVF
,eV0M@Ke4Ra(DT[STVZ=YIV[cU60/\:0ILAb:AG?cDS-ZX100\Y[d/cOJ]XA\7-O
F8+Ie,URW-IfJa2&IJ+G3@_S2K,2AQ#b_W34MBW;LaRO6DV33<MQSSFC5AGe-;fI
.a>^1\B[3P0+#<TJF9-6+O,[R&E(M&2(W-E>GQ]GXL5C5CQ?dKKLa[&GY(BcD\B?
:3-,De<@38T]<(TH7aYW/UD[Q-F[JH;=F=+?C9=<;W(gQJZ09>@Af+#Y+Z)/\e^>
TUEXV,B>N;bCe^+ed<25-&J@4[]G1+1:RED/\PB;3a7LOIKcCW_4GKFYU>;@]QDC
dUH23@<;B60_354WgI<X7?[=dF,926C?/0_J=4BF/SZC@&Vd7(74K]C<a6.N]DN+
:B1X(MbgY::^.]?>ZZP^d_9R9CH/5CU;DX+T-V,_3.@DLRR4,-YL/=EfO5MaD77I
K+&8<H&I8,FCGQT_<3f7O>TES:S[8=@(FIT&XC+-1>C9_8L6H0CA[&K[NZ0_;#2Q
><KDVC[a_#d=CcI_b_=N88\-V^dPB3bJ)R@UY^IQ#;8VVa)&[+9>;_KS4[VR^YaW
C9R?LCf0<0PXWHR?^7M3^)E4;W?>>-3aLZGd6JSQ],fNK?[90PFSBOAI23<-4A;d
FHIS#.1Y1YYT]3Q]75KT-7A/Z^eWMe/d_X6N;JbfPV4QYW^ZRcI/@CO?ECR,0<52
GQX=W.5AAcOD2_f;NBfQW=JM1KQ5@WgMC-)2:UK4FM4X[M5@<F8._?Aa:+_>3H[L
:HJ+-[?MR)34c\=7/aX>6(YNGD??3./5Cfa[+=6#5SX10eJ_QCQa[bO/S@bEg@&C
R:_dM.2R-\E3P.6INS.#Sd=5RR=3QD8MZ_0-LIUNKG.e67T_aR=A[(<.^2X:-B9V
TU#Y@gD6]_PTEc0aJC/3cH),G>NO50HG@e(ABM0J9VL5@YV31DGC26LNdLbGS@M8
SF+C]N5O^]H46=RZ[(gE:W5J5IRRN<1fWd7+TQVH.:[:NAMEC=&aYMENKE2^dQ]L
E)]=DeV..fD[EMI50Q?P,TC0GN3#UfK[3@9RI1dfgQH>CEB6ee.MJ5de#I].c](Z
3+eMD3QI+cZ7FB4H762,LgZ7(=/IZ\fWS2bMX#ST(g/@DS#1.U-?,^P)U/?8-P0/
:UN53B4&+@f6R2<dR._489E@@_5e#;K;TF4HBJ/N1b3]9&Z?E)IcQJ2CU6bK[>2H
>.d.F_aLTY7D\>1)(2)>FCBPJa/VeKJ5KbED-Y_5AgRZ;fQU^Se\8_M5Gf:fU<66
Ja9I;9/.Bf_<5T<((>-d76\G=4[Da-T;a8@+VL.cB_MR=ZCW3RC+[HB@^AbXK[@J
ZdN4?P#BMS/1+SV]S,K^AE&aOHE]PKfOQ@CL3,Q@gG9L6HS(ZLZd)bBVf[(QZ^-7
FA2c0Td9<NO,<,)5OBAAT=K0:e7ZW1J#,@Hf+KR]\/Y)T4?>aG@B09IdUPb@;c?.
A(Q:LX,Z@J;X(9Q,_a8@aEE9g5^PC/R,B\8XHbKH#U#8a?>YB[/e]K&;?Ydd)XE2
4OMVYQ^6+Cf;6QLYM@4-R;9151#,OAYCX@:4VE9RCC^fU-;TXJ/f7S=e/2+MfA^6
QF>L9MWZV-KDd&9a7>Q4ae,D&4a1WP4ME-?[X]OW9Fa6QfGeXG_]TTP\P=Pe]:A\
=8F2,#H5R)gOeHW?WSR\=X6JS,Y@4333]-bA9a@Nf4@g:SF;2,1WXb#_eKBM&B(Q
K(a:^=+cZ\=I^G^UNc=UJ_c/F[W7YU_DcAaMO-284eZ4QIVDNK+P45]J.JY?76,N
?M0-<2>JLNER:YAPO;cAKSLCdW>XSMK/P9-\1N:d\WHA9A]&T<KJ^gX/29fI>OHe
2+H@9IMIOU-deU+Z^F(G66;.PfHdO9JfV</-Ie^03BC5?KDS]A6L8B\X(fgI@&G,
-)[-+B(X51C@cD(d4_&M,JeXI.3f;B^]FQea=-C<AW@H-e#&)DG;?6d-.)f#<KW&
L64DN?e)1eLSK.ZBVM>,X5SI5LC5;6GEW9cI_HPYL2Z_(N3fC<&RW7J/C]TY-U?S
)_<6g4[:>d:\.I,HH6D8S]@1XS,<>P:-0JUR<T_DMYD&Z-R=\ZaJW8(3WKCFTGf/
GTYPHRZVFcgK[ED]b13,)@PM0eD7+7]7OP063>7Ee_)X^Yb-+/C;5NfJ1I8DSX<(
[N_D@1_^eO1=1?B6WaUGe_=WQMO8g]E\7e:\&-(GX3J2^\f?[RD@,9?,)]+T9bJ8
KYE(U.V)4/S2<2DB.(JZ^g?Me?g+BUD>8cQ7W);HDN32dH3N_>bbWc9D;e5.dY7W
.H9=B47>H[aNJ6RbAb8.bYPGV.:ZUb6N7;/8e5Ec>E@^=<VD9(8TKZDQ=P5FG.c;
E\a=5O1?U6?Mf7eBEO-&=eQR:ISPMa42:^/3.<<&I:/0:BK>C6XY422_WPT@92^/
^DaLFYNIKRg=77/43?^Q.LU3)3H^/:&[NRQb9>LEOYG>)CV5#e848a>&=1F@[W3I
2^..>aT^EA+S+M>^Q#X[]aN7ULe1RaB.6SGC_d^-f774AI3WagD-<^[232AFXWD=
AWee8e>e0a0I\;(dPSd/b?2(222T_NO<5a>:2(U>K0Mg4,,C95.d.<Gd-RR(DE@K
46)=/Z/#P37UbAPS^?gKF@GbL:QG4+e<0Xgg3(--eZ?7N)S,,#6R3MT9?.(d1C9c
TV4>UF?4)=>e563eZ5=&7)E(LJE=,5/J^KEcMQ\QdXW(a?I58;3@6Ie[7V1UB:G5
WCIK&HT4+LVUDBNS[P(,?T([/5>&?)D71SNQ[MFBaf9Ugb2<fRFZe.a\,:]_-(AX
Y\DHFJ/K\X\F6c,,0#fWFEA<ZF0N0;(.QbL8NZdbOQG+VNLQbD62FE;5AU6B(OS1
322I[4]:JB>VM<B-OZH[1bEbWQSWG+<E0(L_GefL,EfOMG8W9geCI=?A0.98R&S(
_[&[Q^FCb0\#f9J&cHZ.2S-)4_[T[[G>H<UO1VXeCX/fU3g&&O>IOe35a(a([TKQ
U2LDGaJ3E0KV<9_\=<O]NL8P,T141U-HT^:<KSb-02I\J<+8G5;Z;CF:8^JI,I#.
[+cBY6J6+1V_-EL/]7KYX<(Q@eSg+)4X>=fbD@R&>-,g+Cd/-;_8\S<0:?=T+eZ<
/F[DOJL9Fe+3B[.fH?7#Eaf(]6V=FDPT4P3#Z<.-e]3Pe25>7(C34#E8V/M1a5SA
Gg97N0?M2f,W2d3:P)6#4?7B/N/X:&HK([06_S^?I)6fNPc)1L)[)NSK34E^Ue_V
Pbc^U3/M+bf1OJb:ACIbQ/6(@<abFaH^Z=B>IZ.C1IH4-cb9(;:\E=1B9-W8D[[K
DWZUJU0^]++:AFEgG&?_AddL2#5Hd_[T[)<a][[A,JGfUAeHWZ=cUKJCVHZUVZX4
XcCcLEN?NG.(.e#[]JTB+XZ2>>gS=07GdE]H16-]>b6L4>+V6g5_L[7VM5V(2d9@
@g#DR5<4\UNfd,U5aN6<#P/fbYG?,-=9MO4OY81VYNUOV&^()WB/3,.3D9:&Bbb8
[6>HJ@E+MZ/)5H9V@59JU(G;+Z(<??g&W\#?ZU(@6P0cQRUL1Ye_e-I[NCQXF&@S
\#W2&<Z0_),5gN3+G?1;_5J?A-@L1bReW<4YHDfaB;L&]+f8^<2c1BB+_f;317_?
2MM]5+9<(7gG8D)OOLOgeeUg0^L,0M-)V<C.5YI5/>f8@3[a1\>BH]::QZ&R(QHM
7T7IS@9C1FG[GWO2,U.WOdU:VWTRT)5f:X)7g&-;K_9aZQQc7_R+O8decZf)UR>A
f#X84(K.?5:G<@>AWadU1<:fe033c,dcaPK6LF6T3a&<&]D+^DFf+==L/:afG<2d
LQB]?]YC5#J28ZJ20a8Wd/Q5,X#26ORP6/17.Q=^F:1cKFNe/H,b[2dY#QgM3AXJ
4C[UQA-+N?XK>BCIY2R4EeHePH,L/JEa,8Yb>Fg5(<[TR<T(GE(KWT//OB84]^T<
FbL38=W8HQ+[cc;afJdS?<,4;g2de.,2)&Ob5Jf/)1C[67F;YZ.YbAAdVUBXaE6Q
c_e7J&J8[MMGWa4+\fEeH^WbD=FPPQ4_YWcg2^UHD6./)D](DF5<fR7<3FSKA^MO
]5/3c+Q33gGXI3I1,>+G^F(T/>_W6\<NYWg)@B9[)DY+D/b2X?a-Q[Q@W[b522OI
570.&]&@76A-eXQ/J4aKR=ea4C2GE_6Y:D3]S6[CeCS5eI36?B9dgG2NM?Ac)_-2
PgMZ2:@/1.I>YA(aC1;-KE-T0NXZ4EQKYTZ-19U8YSJOWV_gR,9JWOC;7Q,AZ9H^
cI?BHe-[.Z8G[2VR_)EBAaQZ[OWTJ=fEeB,^8+@KdK]6O5F@>6dD<4IEb@NJREbc
E5GHOEg5+JDSE+fD[)?5&]YT^c^/b125BY58fNS3O6+8O+N?1K,YKP0+4d4Nf4#H
L)?2K+cH#49-F.I;ZWIC<CMKedg8R;3gdP-c.;MYQR=Ve,?Q3K@-#LF7^6g]A24#
g)K;/G&YV]-O7][6Lfe@PO6X_8SM&;]H6X7+D&2U[dVbcc&]S@=GVc)4HbAUY3g0
B/OYT4QcR;5bA/F5#\A73IWU3c)WF6YA(;fJB_YS0CPT]CN)\])CHA.dO9H#<&Y_
,4;).A+NDCQVP,<<:1)&]f4cZFc0IcMb)<S-23HPWWdMa1Y5PS+Pa,+,.\8N1+Z7
gP:HQYdA:\C3+c;9RAd=0A1SFfNXK.K)G(.eYYaJ91]XR+aU5#<N735BIATN#_9g
&/6S13bS-1<(3+Rec2NQF#bfJ@0HE_.SA^GbbX>D+#&dE4f8Qb(9>W^-RX1cb7\L
&4IHcR8SOXC@]\2K>Z1=[L<\1V<eG(5&bTATZ+Y1gOSCJ71Z=N)#WFWd>]+DU^[f
PN489M=DT^/)?FD.D1K_))Q>L_-gJP0dOK&<0+gCO_,g/IKZPEfU(4X=fQ09-(B/
+E_ZcI(G80E9?,H^)D^a@29\8GK@FG@+N9L1QBT[gK1AFd&>4eRQS1JSc#+K0W+W
e:QMF/0@\HMH6a[f3c5D5:P?665GVM9VYRZKE^8Q/>T@(8R[D8G6\PaCK\#KG7BY
:<_R:-G:O(J4H]<;FLaZ(2)0<0MK.N5W+fBU9R_.g?a,6[64NF03,?@aJN;.>\)A
e8GASK&H=d7135FGJ0ea-+S.8>/Re(LBL4K^[\\T,^A]=((ZJEH)&KQ+dJ-:BO#<
L))X&aMUQfa@+-dEU=W1OV>@RO:eK+e#ACg0+4;@P(E88</8S\(1<,U\8M?_E+;Y
U,E,<:V4Q=8<K72C9Tge4U3V@7cRRbK/O\12.RQF?C>9aO0,XWT#TeYV\T21g94,
^=6:F571CKLI6=84N?A_#g0-_eO.+7>Rd/(ZJJ\?GK[_bUOdP)KOGZKAA]5b<4>Y
.Ua_7GX[be[>,58c^M2=GaU>+-9V0>ce9N0#G@_SCXY_2>J+/K@+<)@H+YT@?E5?
>:9?C#M0()7\>UKY2VX\QGXQC,VKHCET9\-#>):8V+-(#56JZ6;IWD0>e9WDY;FD
>/2JNJ/+8NI]QBaIT5>9S45#T+<)Pfb8a;-P5K\/,X1.M7FfeD^IXeY5AfSCJ,g7
[(f3;W/>T88_=6^+A3/1,V9/5[,]HC[<bd[;RFPNRU/8f<FM6(>V\XC=ba0OI\F:
If6IJPQKWcb8,;ACT;B:BCSP[]N11f=1OWIS-&>4/a[]8)d?:09N64MD=A7Z0D7D
)SQG/T,E?N2U6DC].S_bIdH<0HEMTR1aX&5fB,G:eFQ[EC&3\,DC;X?:0/W=^=P?
fLP&-D8F,RI1.Z7Y(9JPdP]c0NJ(Df]+bId(8GbQC,_YA;3V_61f_X@7+cDVaA=d
RU39N=2fZLFOE?J;CD53=9A:5A:C70XZ,>E(SX\[VfB&&/4NI;WGVeC1:IE.\4dJ
G+LXI-NR0UG>P@#OE).+5MMc>E[672^&=C@C>B2bE5)2]FN7Zg-->C@e4-1.B<Y;
@(ZA/H@E5f_S(N6,fY(a;#eWY.9CWg@deHYO1;BgC#a;cIM5:+G)a\GFe0H+X<]2
\>Od7P3X@)RBO)),V#?.fQYETMKEPgSSKFb.T6OG>I^W&cT+aIdcSMF8bX(V+USQ
]#@R)-b8g4a88,WZI3^_JX#CfKW=XV>+d8c.T3K5A@#KFa_2+ZVZNeAD5bf[^V;(
T3Mg=d@M8?Y))\ae-V<b:#OQ/-K;DAMTOZOCb0/U;#EXBdKc?9b0U:d\.CI2Q:a>
RBEWSJ;+:8P3=+A>^Jg&O9Kd@gG:B3#_5DWX5GL[7BeKa1;DH+^1+;TJH]E;>Y>6
Y@T2I._B/NL@\]Q?2B3NJT<B+?>O/g2AK-<aWacE/27L>EeQIa7+<[de][WAONU>
80;W+?XLHbCdS+TP4?KI2fUT?TdR,@A/cKKI##MM@KObRV_34TG,(AZF.ZGLe((D
0>AJdMC,3N45GHcbQTOR>@gLEY<PNJ0ag/H1/Ye2f=>?HFY@AC@?O4)GX8F;L,Bg
_J=H@K[XZMUD(-4<KTEJDS3A(LHX:T[\ET1/[2IF)Y:0V-^a#PV\>AaL9W.3d&@a
9MCVH8Q[^_</>)@W-?bR+S(\1VZ,B(I9NOP6F8<JP)##S@9dU;7I8^56ARZa278[
^T\\bE)3e;O7>KOe3bCcP8I=9d)5;W,9@R)cO=[G#=;E-LaX^I4DA9CD04fb=NC=
.\BSKfea,6IUH_UU/W9JSJa;S4S0gKQHAU[Be<gIaNZZU_>aB5LW&SR:a+(K8bEO
^@Db]L;7]dSWSKDL+6M_&Z90>>D2Z0S,-/T;fdG[?W&P<CY?0Q28Z=Q;:(33V_0e
aL7WT;OF@bB\?<G+F=L,S#QCH+N;D-O\Q7:fdSS\VE0AI9e5WI=SL1PE^OXZWb#T
OTg;B\/HN;XZ[X@Z>:7Q@#\-O.DL]HP_<c=633<MSK<R24bR061#HQ4]bN^H#B[S
e6d&&AALW_)2b;H8Y9Zd/VW,>,U>d:^9DbIS87KAD?cLQRa1<3<[-G9(V5.Ma],^
@JTZR?CFgOWC@V\5<:YfFH<CUNY:cQ-#Uf(+75QRPY0_d/<C>?HO4DE1[f;g1.S6
Dg]:C,9\G;;_Q.0/_RTI#_?3[Sd-]=1KfKH)=M[-f;40&OUA4O_)eAY+S9UK)7;S
.:+L(_EKfFf<8;3HdeP]>D)dOg(^^Z8/)EacQb[2RBU[7,K@b5#&?&JW\Q?&(NAa
CLZ^CTfE7EDO7U:&e=]_eg,@S;MAO?ZSVDB8T,2._cQXRN=B7dTC7-GbbBMH_F>P
,HQC?IAHB8gbB[PZ/.R9EefC>-??/K(W_&a/#eSSBN21Y/PB&=.H5O94IGA->dL+
:Ee/SULHL?3?KQ0LYTDI7a\>7VVMb@g>\_.1[-<1(dYN[aS2G[1e[c0P,\[8RbL4
7=KGA3HPaEC;:M2a/ZU(4DIS-UXS2cP]dH.^V:@G^_(ST@SNa(5>B>RBM>5?&I)F
U9),T/;VJ806U><bgc\dMQ<b/0:F#&F0+TN+KZM-JHA&^EA@D7E_#5:H7&0ZM8];
&RX_B#7<FB)1bAUdNZ3_G1J+\DW/[=d=[0-.A>c<0JZ]cGc(L5;4A+B7e,K09bSC
U/MCcJ]AEIV)Hc]I^)8&;352B)FA&.>#O>ABV-NASb.U5Zf\aB5eMWAB_>>Da_e)
K4NF5K1S#eI=8dS>]/H^0-7\HM1QH))]H.]e_aO0)&D>[@L+X;O&/WK2=>E)98]/
#6?2ZFK85RNYD&Q3D0NX3^W6K)^d7UHa7??(@(W:;X/?a&M?]Z8ROTa>NB>&Hg]J
KS8]_ZIYQEcT<Odc9?_+5OWZadCEW=fbBb,X@<[]J+WC>H;6?)R^>P8Q9F\2@)&J
P\I\bg6eeZZ2ERdY[F^d4[L;WJ9>.]HMX?PcU>_Eb3+Y0_>JQTD=U0V-09J8#Ze<
HN4N0f<A9VfC_]1PP-IW.(M1C#S>Ig=P<>AS#_0SbCcc>9&BB.g+dEbeW8N85L1M
7IgIYSeO.I+a-P/AP,CLWM[Bb2^KCOZGA5@.-fM>)536B1f7=.7eG,RZVYg?gRSH
.IXZRK?J;Y&8KIH47?X:H&Xd,U9.2a\MgPd(170We/g?gf48>1=DIe<AO158BebM
DMVLZ[A(HBN[>\=W-SP/,8+-Zb>MRUD>K7?9JA)AeGU,AL01-D:+g^[(E-:>VA38
M9V64-7Of#)PPYSNPCA?GTSJ#K.Tgc+2..=O<IUB()/H5XP&N.DC^:..9VSJ@03T
>?]\edHK^]2\5;>(7>P4F]07[RU0_.5#+YZA0@.e6CYT48:R7>72a]G/.3=F&#.D
N9[I?/OV=fS,Y-M?)U:1^>CXf48/U,/[2@CPF\4g=?@:/2\Ld(eN=W9DIR_?5,ag
-#-MJ[COe?,,4d&YQPT,R^9FMLe+3e>BAg00</L,:X1F[HO48UVTI0YgfaL8/R99
TAR#PB.#@;aWcN;D.Sc+5gOL4G&_M>a0[<Z9^Y):a)+=JMb0.<]R)+b#GD8SG6J6
AU#L6.4cIDB#3dLMgQ@N\eP5S4X1GZ[I4MQ5_@@]b,UdY674M#&MDBgS3LA&15Vb
YML)3]]I>S:^-7V[2#P/I8INH_bPM:TC766H9#cba1[NNSD(WCHTQE@cd1LLM22A
E8(ab?.CX,<LB;FMUOcY_A+6g:=L>fgeN2Y^\^H-Ed&JU+ee/<B;,G>(9:WG)JPW
HWTO-X9b4@ZFC.Aa?-I2UQADP_(S8dAIWU/EUP293XBF8>56B[dSg0^V\N84_S.3
Q,/]9eN\QIGDI\BaK>dcVS^bRZLeO^g45\NB]K[^D^9K>0+f=aV+WA2OG3(7K/Cg
[R>XSG5G1:cS@a(5#cRdV?W?cd7feD=_e\#@I\[-ae^GSP.-A^B.@<La:((8,/9N
4H5)f4&5IKW@;9)=SR:\La)(IE74Q,<N3B:AA#A>QNa@82[X:(M3N<T],Ve^0&JG
5aKA63PVNZ-U(9(?-F2Y:6#H>KcDW<&4VfH_-]-9WFaZAPGMcKIdTBGD:b&[VA&H
@e^U6@)XdM,RI\e5=-09H@Sa?@MJ..b6Q+LQA(cC+I;@b2(^RD1fL;B5\a^e\0Q6
Y]S3[.K/,ZdTb(b9^Bc#546Z7Db=SAgGCAQ)Y.#IH:_7D;?QF>TEDSHF,QcR7eSV
1_EFAa7L@.)#5#Z(Y?77YKODQBIO](VXg@[BV>GZ;Z2[F(f:3TEZTW<?(,cLYG8]
5#]M=PQa3bKU+>b7YUEb;4ASgI.:36JC=R+,I&\+17]/P#T^)5@f.J./92<6-_#,
)(O>7^eF/BG?\P;NC=4>6A#MB#/cTG,M6MZg=]TZJSdJL0CD2F<G=IBK#Q9#IY/_
2f.@.Q\dYUAaMZ.A)2G)X#IC&Tfd=[H#;V,<LeS]e[&F).4U+8,2>/SW[_-9g2_e
I@N[.d^NFUH#(;BL+G1:F575OPFCSJOQL,O#9E[,Pdg_f[<DDcN_W1)]bXIJGQ[R
6\Q54d4G2CI6TE;8K-J@3MQHAT=NYY^DEZe,OOB7=M^3DM7,IL+(BHcM>/:NUC(B
ORNQ2a;=_<+UaY78;)QLCSR2_B:WW8I1]UI>=32EZKU.Id)]?8:&F7T-Y(LD);f4
W1:RgLY7IR5VF0c,Z55P>cIYP/PE(;GdDA9=@6&I?B3aG,>FL<5=EaG;1H,+5Hba
3U=WCNeFP<<0(1@MRf./a2:6Hf9E7U\6a>TMY)#a9[T/NS@74:;Ue.(H.H<XQ_b<
WA3LXI:F]2-2XAZ]cP[&<\ZRQ7f,+1]+<,<f>2U[cgY@-&]<9M36b4Ve-T04,fT.
SSC=R7R0?U8]I^A@A-BC#2ICa<RNZYCILBAIMZ.]SAfC].@+,PRMV2g98G8>[;H@
^1YMB(=Z=J_N33YBM@f==RfHd):Eg(.bFK8@d^:8&fAcZ7g7fUT_J46?_6TSD;Q0
+Y/<];C;6@(_cBO9@Ff9G&,Fd91.9Q]8eBM2P8+;(dFLW0gH;.e]_Y(2aFZ>1)WI
3WDfW[2JP\U=SG6cLYfDeC<U7I;T+3L64:.[A@>@AY-DfbR\RHKN>W,Y9=;<J19H
Ha\AK<VYA4W=T>AC9L.#5FJ9dV0FS<FJ@,QBGCFVMG?J2/VWa41&]=\8001#b=&8
Y)>XBdgAZJPY609^Y3[]:V:)P#eJK^_#:S<@5HTMYdV=4NDfNLUG.f\VNDD:G2Q9
;>5Vc\PbPa[/OM55fY0R5O[I:+8^);D]2P.5D,]FQRNLXK4UG/]().]<@P/:.<_c
;]7YGa_M7=YBD;+8])Yg&b4[U&^89@e]30b&1GHO@I+Y2T<V=BE;6^eR?cg78-K7
R?H8-?9XO6.&)924T^cK)3X)IFb33IS#E):cXJC6-MQa?e(JP[a>;B#NY<DXTL3e
gg&;ea;;eA,K@K@I+G^I8PB-YK#6<<,7&8-c2g2a.3FU#bUM#N<L.32V<JB9fG2d
0T/8fWN8QLIDK-e/g0\5N4&,<(=Z&TFG:V4b-Q:E/e0_,NKX)2c>Gd#3Ad)GUD1_
:1C#c-c&14-+I8Z:6,ADF9+@P8Fc.)JG?7#HCI3]0D2gWK,]6M)VW,TZUO]Y@2[,
=/T3?R59a31(5J72?>)fV-eDRM-).S+g_^BeHDE6DMYXA\#+ETGZ&;30J-4Ee8#>
eF.5)6B31U53;>g9K:?/J5AUTeLD+DH9/gDBJBD7-(WcT6F]L5YJU7W[RR:3WVEB
-4XAcH916a1\4ecUf7LF1K^6D(/-05P0XC::U/G-3(IO^79C>2^F?H/e6A)GZH_W
]4F6@Dffe8/Q](1c/U._f-3UPM3>1d]bbe4JU/QEG?+b<_gD7D,S[fO56TT2,Q=,
60f(K>^,I_7UAKP3YM81<W-J@26KF/<YAa=3D/B]H<8\IK96.X2Y)I8KDb-.Y]=a
M0BUXS?+8FE<O^4PWM7?Y5;Z0IIP:3WLZ#[[Y]0F=Jf<NR,ET[TWOQF.+UJ0KRDV
C7@R-[#YFMD7d6)H\L5.gN\)-@F6U(@/1TaQ;MEU_ZEGH-P]4b]UT)CL18_#S\cI
HDEa=:f4V3B.?CJ-_<4WV_+1I=@&CN_+AUD-<JD#&FX,R\WB=;MG[E7HMF#3MRT9
^=\KJ1LGI5SZ_8cBc=L<@c#\F4/E>6(XK(2?BFY(].L=;^7VY;AD01e1\gZ.]9Y&
H8_RYOP3]eH@f(5>5#);e&[Zb9b/_f2gJ(^bA4<&&\1P.?C:[@+2DUQ#3CcTK_Q4
8B8NTg]_6P4-[FPZbDWSEO#A=e<M,]VJeRLWH+b=7V.HY_UB4@bYWS&I-#5/&[M(
\Va][>33RKb5KJSP2K;7ZPe@PULW><3<Q-,/U;@[4ccEPQEY9c)GNN@aIFM:9QZ?
TgTYI68;b+XPH7?MGQUY//RBK34e35:@PSKdI^R4Ld5(KP?W:JSHO@CTPJZ7Kg&Z
3WaeY4YW4J\)KM;QFXW:a\7_>DIE3E>,)c._^#0E=#<^5U8\,Q?4EBGC;]&P)L>S
/95c)9\^]\3_\<fb;JX[?C]S@Rf3.YYF4,&BTF\#BXa@E:dWB@^O5[5gTF5B7@Q\
=THHC&\?3LY^2Y2gQ];PaXVL,]4?Q/)(.SRL;<)^1I6[^#1J><ZWdd<Qa=VNU2H4
;dI#F_g]YJS&6T>^gFUKU..2]16=b[a.02@,YESb46T]:;^X5C?g]c=(]W[/8e)(
L4#<=4ET)e5=]Z\JGe-bBJQ1aF2?DL=X-S@Q[0RDQECTQ_W16a),O;bJ\7F07G<<
c1Ng\dKE4:[A&ECO<GggL3A[0GRNId&\6B;5dO5GMYPU3I,YbY?gD+LLaXf26FO:
g0QHI4=@RRTZ^(RRC^-=;?N[H5cfY7,4(-bgTIWR)K;P830FS_P)AAbXgbUMISZ1
R-(GfVc8<B6T5[0^7VWbTI))CX3B5a9Cc-Q@S;B6PN=?b(6fFgI8S<>5c9]g8_f[
EV_=E3G3fBMe:UIJ423-Ld<9=G?[+H15\Gf(F6XE&9D[acaPWVGH8VE>H@d]Z43A
?H(M<>7M#]-^)^dLVcZPd]S/-F=B#_F)F6>,+3^-Q35f5.>4H\P?4EPZO>?+V1g+
7&^,F[]@X?IMWH,4NX3[1@a43>(L0<W(\]d<_W8,>A>JJB9ag=TQ4AN@46C;5a,3
Z6/dD2/d84@&d>,#ee:GNEDb@-L&]RDC_#@Qb>OBRR+-KZ9V<R?E2F8OdZCD4)1S
P&HgbV_M)F4L@PGg)&FE8B<[LF9<dKI/XS5c\I)1W=.+F5<TFIf(YVF29;H-NS<O
K5PF;?F0c)a-9a.0YS>&d+:6f?#ZUTC4=(;UdX.U5P-J)AX4W@557&GG)A)g=[EH
XIeO.0-@MM1X,>:5RZ49SJ[=\FgP&>BV&I9A>@?2I/:Z:<A/1Sc;OZ#_Y(@Y^eU:
_RF/Q##KE-^N7]55LSXe++9_IcI4De)bf]#/Qe<5N)-8Y\fd8)I=C@-8c#P+9-,F
B91fW_dMYVUOGTa7U>4]R+KYX.#-)-F]_/S)C,,0VOaFcRd-G9//dO?GP@JA/a@I
(8)@9<f[P@-QRMR50D8d;F-3N0(BRKBAJ>.AWcc/40WfVe=BLgO7bcbZC6STCQAQ
gN)F;JYQ(;3IJMDOJ8S-DEL0gLA:F8@5Y,=7@@aR\L]GI:ITHC0NP6fHaXSWK2H=
_#g=UAd?S(&cT;J+XV)f5U?FP^D7TbV]0U47T,(A7Rf_8Y1Q;)H3JFL3O--0W_BU
4Y1Q7f9_VI//eHM:>#T)4CaX<c76+QdNW8Cf^G1L_Y7-I/_?dCJWQQ(L1GWH0XH2
7,00U,92X:c/SL-5&\D[b^7_Y+UZN)Y#S4@KVK)f=^e>/USU^We8ZfSICV<[N/OJ
YI)4KZHgd11[-?]+NSbV8?4V#I7Vb(B011([.ZB>TK2<G_FB<-E8+GZ,#K\5g;H=
_TIJ3N04:NQ2J8Q,DG(V2TO/TZCf:1[R/^-#G//Y<[EC+bCC4NGJaR1>0MG<07V=
.+IPY<d@N8c?CELM]]#ZF91@G^#8_ScRS[09X(gZL9HQZWW^IB^BA>RP;L9@c7KL
e9dU]YRf12O?d6B]<aa;X=N]BVM3JVMGEg_)@6G55?OO7D@E)#FC.9]J=9EJF#fV
]4<XA2Sb4b;0_4+]JQe\)VZ\ZbDQKHK&-_#<T&M-S^0OWB^a=e-0<cXNX6[d5H_J
4ID8&HIQJ26CF_?gP-4E.b72AWUZ/N1_QIQ=(QOA?b-#Zc>T54?CEFZ#A7gSK8e7
c5N122:N56UZf]Mf6,3.Z#TZ-+4[62U2W3&W2-491@g_-,DfA9,-96)b__HcU:?G
f3&2W,>5GA@X4S=(DVG]>/Z.3E6M6F1G,6UA/9C#_\GFN=bfI,BX]T3gVD:#bb/^
Z,?KH<+I1aXU+H/>]\0(@W(Kf?Pe-K7Xf;?^^W5dcG<U5<+(0=I]XZD=0RC=9@O=
Z-1f72WgQ5B84H#^c1aM/L_@a9:R@62,gC[YT+(N-GX>)H#aVEGeX:U0(^GNdPKQ
\L68860]+S[9-Z^0]a_]/cbC.?-=^0C;(/:D7Y4&85[^@aKJ&4D]YVg#E)43@WIO
)3X<Rb[OD2WP2\=)W6:c3b]C8.4Q\7F#89/R,.?JODN=CP+YHF]U,^_e]F8.gVK-
g,M_L+EGb)-b[FSVEY3+@?U>@E)^6aHBX?g2THDJ0W#D<5.;V>B.-I/FKcB9KHB[
)D&\<C^VdfIG1&&N]9SFb-fc;e:[V&.I64e+NVWc:HYZZ=f#WVSPTFJ/I]L0>eC9
&HC,3E0CU.I.?<Y7fST6W:Oe0(UC)#P[=e#HegUWUb=FU#6B/9Ac[TA33[VU-AX;
LNgN2[LY),P3M7.]]WK\]3OAaF\>IWAdPA^Q3_@a\B\;,WFU3MG&JL.\eA7_:c48
P6N##CNf].d0ZOQ^8+I)PF?5:YbX1-ATeU@-^Z=/3[L(<fEe<)UG-_3fZfIYP8Nc
d?-fXB)PD:e.]J^L>/gX[W76Z[@?28M<?HT:@I[f@RIJ7MO(LUE1.4+5)09WFKe=
.a/C.+;;M>H>C]7=O3KGEXXd.0DDdGJA.,48=3:PVc)Y<>O>SLc]PK.d\44]a0=5
\MX_S[S6f)HDQ+N5H.D&_OCg:CAE1QW(LYIG&P-OJdR2gEAfcNOFb>^@?#L:MCgZ
e;P;_;6T_dU^<D4#9L2VH.+@ATc]4#:^3M9.3.TAIa^PZRfVPaI&_V3=B;;N=Q&8
G3@V1UeZVSFVZbeU-5G:RB=KW=,f^H3@)N3,WbH(8VZP_GbU;7Z<VSUR2-Xf_U6=
aLfBDC,c_-&LPLK[K>3NGBM:5W.8Y/#HAC23;>GE.1O0P<6.H+Xg^0aD-N\L:)>\
^/gQ>/;&:Z(<ZcZ;(7B7E4+\T-dN3A<EM^?[/UceaBD1Gc#&Y9bXS@HPP1aM@Z=1
,Bc9:9-EF>X<^R816AG.U[Zg29#]DR1L,U&\TMK:J>]R81V\@\9\8bT>I<2efO?_
SX/JMDGMTY8UZQ#?[9a0K7M[d1)a(Q,,1W_UFZJb,X#X]J\@e#T2B)=>F0N]<61@
6I=Q\bNHYW:=H8?DGX(G@g@/L0g+4;dCJ<=_dUX.+H>FLGC0aEbK>/T(8D+)^#gV
cK58<<6XK\C33&HCFERDIMXf;S14Lc5g9FO=]SF_ZdK;Yf@A<Q>8R7c0BEceXKA)
a=UePE5#0-#8+Zeb]dWg)K)+<Dac@Lgb3]B0[KO=^OR=c/\6\X&<<MN3.a;=]Z0B
V0E._gFLU(8g]XT3+#RN^7c#M5ZVfP&LYK0UV_(@B9T-B#XTAE/dV:E>#IdB]J26
W-KOX#O0[\Y_[Z64V;]U/:Lb[dDSfW^191ZI&-R;2G5L+A/992V2e0;e\d?H,+Ge
CV]6.58=g7(UQO0W-R#@/]9@<0EO>HJ=]F74bZ_Z<P@LZQPK\R6H=M(^<&1+RKBR
]6XI\,HTHb>N=bGN4O]c)=e84+2RM?(+:@^<d&IPV3PFRb\PZN+]#e5MK./8<QAg
6ATL[fX@f8#,083M9=#fO/GHa][/_dIeK2I-KH3RJHg.G/MDXC_;6BN2W[^fKZG+
OWcP_;>:Q_T?.#TM;71)D9I(AP6>\>6&14L6cY]<a-H,^^WR_+(SbG(^B:F&L^I]
S4[/Q(JD^?]=Rf&WW@aCF^5.De/(>/AVUAX[:])O-7)A5^Gd(4Q=d>^Q;+M@WEQ1
F.-=,>N&X57M9aX9Y,APCRL=1B?6RSZ]aB^S<=U+EdPW5THK,D;&M3J#]II:AAS>
P1.P_1Q^1F1+ZX&E&L4EHSH8Cc3XF_6]X^FWM8Z\^UJGVL)-95D^BR-XZOJG53[;
?eK:9UA5ZG=^81V?YXHG0:S[P3?4NgHBKdU=-UQ&cDHcbT.VBXDc5LeAbdG.([#C
R\8=>G&Q79TD1LcfH1BPSI^JP@QG4XNJ]CcP981e?H<+I#0Z.QS<PWJ?aD9eNdaK
^_(Rc:8WBf>W@7N_;1ZM#M7NN)>gIeUcc+_&.6]LK;&K)>\WT)X#Xf@JZI<@7KH;
ZO5bSO]bKL>S):=>GBe1_ZOKI^;/[g?BYbF8[GQH#:^L3dVJe:84DSb47HONS2A,
2.OLfM&JZ0]fZ4\_PGVIT&5#Z8R1f+KB;YIDBc9A)P53a\^-=2U26b.edeS9D@N\
6NZBSa[;O3,=@C<eMf<c2EOd2FeO0ER8FBYQ@<ZVJOS1@F)KQ+-=8?Z@3VZT?_R>
W\MT5=\[8QC@UC0O3fQHdPUW1eWE4<V;^VGXMaISc=C>X?/JdM:+DI>#e5dP0OI-
UYNXfTA2]&183O@b0V==b=YUBQFF-de3?Idd:,PNI=UCM6,:L.dVX@V:WP2bJ.[K
.C1O2LP-/_,g2PA75^TWd&fL2DL.K/LD(SK?+N(LfTZ5>5Be53ZZ&5[:4XIP?6OI
4P)d4ef51-N+D+Gg__)//e[&A<+Z.)(d0J\8SB\CSXc[@FR+Ae<49OTP7Z@2g:\^
W8<R(-6Oe_(:2Z^OT7XeDV@:X?G\<cF)A[\Efc+4Eb9Q^]d@N4?UZL,QL,[&XVc3
;AX&EAc,:]BC:.@_X0?&G,e3N/Q^U55XDSI4FR1?1[WFL[F@=fZB6bY9;Mc[(IA2
_72<_[A0N(KeLQ9_.(]>2D;[Nc1<6Bf,Y-FMf&3-3..8&/5bMcfF\H>c(Ig>\3D#
S4B&VWI,@31S&dCG1?&/\^@c]/H_L@8OP=IWMW0\\aR3=\eGG]P,f;(@gX#[:XbR
aCU>:BTA9C;Mf:&cGDbEeB>U5DJX32FB7(?K>L:AL7ZJXX+X\.9>]3S;MeeF>Ka9
G@^D>TVUB+P9^3M,O&fgV/P#AO\=d+Wf1NSJQ0XNg3/78eDNG-ac)Hc3.TB]<T]S
BP#NTKf[=4cS^<ZP/J0G@@@Z@PZ;D>g\:O=C:AfMSa59\_)5EI(-eLL8,:S?WG4T
?[[3LS[e\EQAP\@P(F:#G5TX,NU.1X]Y#2/^8/OCO?T3_MHRPAfX=XGH)YZ[4@P0
F[6E9.Xd131WYX.gP?)P-1MH#SCgJ]><2.7WV9PaWONSD]Q>;.7:=-O/M;cc[;G4
YYcAcfDbJY1]d=E5g3\)-.T@#1bI/cAI2P9/.cNb_#ZNAW(P&G,_X_[\0;a&@Pg(
Y#N[^<(NaYTMPH_+)5I5;:QN8E5=LT?bVLRFW<Hf-^=1>+G^,;CdDOKRDX-3.+TV
?e[Q+;=UHXXI/CQ;M&RT-V:123;H;1#L;H4F3Z-(81])bb7-YQRagT1TE9+W9VSf
F<J49(PLB^Q@UITeWN=4APabCPZ>>cf<(3d](Y]_KVc\/#7R[fA)OG9+&d4)?-_F
V,ESaE=>3XBE<B(AS-7^:gf]28^OPFF3/,aI6X@cE@0M3X+P30DZXC/[M;Q&MZb4
?,<#QXR?F@YH)e-b[0bBF:,@H+XXS90c,=/TD.-YT:9ZL8=(eVaO.eVMebR<W&VD
N5ZBVW>O<Xg>cNaFD3_\=KGZ5A6[bg8PF-EC0_W03JB.V<FY3@ZW,]N?+O4_9U.X
.>,[&]F6D1>HX]Ag<J?7.>=]4NOfK=C:#9d#1<1TT1E9R?b(#e79aV+I]F:\:)TK
N:+3FGUK6d3UD+#.#XW39>N1D-]XdBfI?N#Xfd\=C3Md>^;4NDO5DG5+I1HXP,Ie
(&_EV(DJg&[cS0bJTO3_)6d<,G?J,dHH#Z-&^\3<<BI1FC>aA6-fWH8c5QAF-X:_
-VKX:4B5H:4bT+(&Y(M+]AI((RTSV\JVBG[>d.+D/b7(<#D<R(:7+>YTTN\)_(#c
)G>CgWQ5Q9KgfT4^NP9V-&ZDSVB;GH\cJ:6?Y>((GQWZY_JAKfPId_J5[^4,_Z?a
8JG[c3BEA1@W+2P\=+]J>EWS6MfZ#3ANf=<ZKK)2\PC-OVVWNb.N^c\]Q&dD;X-7
F9G[KVU)@/F\[2@9c+c@F-/[J?<cIFf--Pf1_]=7@\WA@e(S]&Gbf-&#+D1?3)Uf
,0&7_(Q0XT]cS1^K(-;.[Q^IDb8Q[DP9D>?RgCID4\bTQJ<YT/:-;IbeW;2Ie.cO
[YU,Hb<;(MP,7gbb0>@MKaX_eN(H.R]NgWf1D>(Be5UAZOO+ZU-&LY_A1(&:1KKB
&>1@G2;e8>@QV2_8,TPJ:f;#(TXS]1I@AF)8B[DT6QM3ADT@&5M\_HAgR)c5SO,U
;U0S,RN#WJb)#M6SN+cYVS;J2RaE2g+=8b(+2^YTL2[NdCa;^/K3MaRFRHaEUP<=
8J=Oab>+.f62Yd3;1@9<+=:fD#bZXO72A6OKXICE+D5bb[T:MaK0]S:3]+]834T\
;O.K&cJGM3ZXMW2;RWWS2.1B,W7GQ@]#)#7Y9<,A9OS^bGb(]ZMX[68>X[0?]@>0
)@6RDa\F>CMHAMP^\-;cXeH9\Q0Q58?77;LPb.g^_P,X]g0^ES]BC>ee_f.3DZV<
65XaaSGBSeFAGfUO#X6X9^0.\VWM-=>8?B;ebQ?V?>LI4N1b:55d<6/SU/IMLTM?
LgVc50fed5TS37P103U,ZIFR?AD?@2Qda:bA>6D73b[gWgTE6I3_\YZ<T3(Lc6Re
Q++^WA=g3b/<_@b#:?QH^.68>T/S-,<<:2^1?18<(IG;_g1<K4R)?K,,V]PUc04Z
d-V7DXaDB41ecg4&&/M37X>07(.&b.S0)S,6ZS_c7EbGeR&R\RPU3-0=9;g;DeC7
G\(1UG+Le[\)Q>8LR0Fd^5VaCeXV@<f_\6#)UT[ga[+)gPET,CG_-<(OEGCGR>XI
L<S]Ub^:<^)T<I\?Y[[1HE-dePP[>Y/,)9dC8H7RaHW4N&_CM5+38K<c,8XfH]d:
0]2M-QTZQNHc_QV5K\b9K?5\,6KJ<B(X=AAU<[_>##+>N9ge=.-FP1SbHPMU?DY=
b#N[LC@aT-]6fSCD88?Ae@N=-GENZ)K)LR:dQYFXGM8\3Wf>8CSgEXI\JNEVHb9Z
f>b<Pa-NM?GJeY3dGL58]JC:^TW[#R3CI7\NUCcPO[eR85TJW&:,6<;)>HQ#P3Qa
-0cMRdV>]]4Y,E2-)<RWQ>:MIT+\O1Q7B-<#^[e;K&E_X+2C.gLfLSE\\11Ndeg8
e4RPY+@CE=I?d@IG8HHY58F347a4g[??-KHTW)(=3G=1HA)fURBge#0),HRKeed6
^S3Cb45+>5<^#RAHPZKgU/6^NQ)2<J]YE)J]FY[.3+.@@R7(D3>3S)TKBJQBc.44
62;L[eBWGIf4_Ee&.(b(=&2P7MO2(;/0\@ZAI)bK)O.BEHZLMN?J5-,2-cOZg:c(
cWM2FA[D1H?_@eX7g-8Rd0XY]0(N=Q]>bSM07KJGVZ&W7I:)-g8EE3-#f4MY?#8Z
cbE>7^JGN=&55.b\>Oc4d_V<LN=b9.S#[MEMW>gLgXX16@=WD88<9dM:&JE-A)BJ
^,.XW+>D85=7<JZD+[7d_J67I1(@_Wg]be+:&P;O#MC(EU3d\RP[C;Q\+c>I@;F3
;@R9#XS<3ge:@TAXZS&f<D,<.VTD,8(g^,XG>TfcOL>f_6?@1dQc3.a-EgW,FZae
LX6DO+DB--a.e.K40MLA,#]MI)Z0B#TN79+?R&@cF[<cbee@2W:aD[\fSVZY1,)b
X>^P8^J7O(;cU#QCUMFcd6SV\b2^CF,_-4]Lfd&L)C+aa96:LP/1BQT[<?@_:WH?
\HJC++[[faXM^_F^B7O24#]gfb5;g9d&[UM?Y=6TS(I8;6dC;e4IYY9eXIT4JeeL
6O4O1[G54RQ4aP<;A5C4O^d^38(O<?8a#cKCG3@BY7,f@^)PY)NcD[N8ecC:Ea+S
BV^WH:Oc791b;U^7J\6U.(RWf[XJ+HYK_9eLAUX/BfMfGNLLaM5@?>:NGJfIMg.A
DG9OYaT\(_@PE?(L:EQ]TPLLGb8@,7L.<A_LZ=aAHQ6S2S];1)H_1HNG77W-5=AN
)J\7/)0Q.]eJQVA>Q49;eG@IFRKaT(UN1_3BgDDB(WK9ef8C&LD=RGAKe#&G3DRF
gL_Y>T[H0[_2eG538X6dF3OP^gf[+R;_+^ZM#eOYa]W0UJ)eF_=-0&Q_#V7\VVUM
6d=f4E9[OB:]a;@AGFR2?)cPHJ#13,IPKWZHVeJ5WaZXN;>OJV=L]=^X(JY\F2P7
a-A8a:E6W=<XK,TeGG;MaE^KYaS;4B:._Jc<.b#OUP=)T311=\Z:38Xb<R&,GC4,
YFT?0LdUcZ[b+Z+cPN8EIdSXR-aE@fJ)A6X]G0E)f=FX^MRa>@.Y/(WQaN710R4.
.JeIF;@gWB1A.W3/NaRK6=SI0(BL.JIbeO^Q7Lg3JWK@-d1\DX)\XNF=VZX8O[>Y
TKbe]X-AMN]:T/Q#SFUG&4?TS:@ZAO()M@F7Y@F]#&=R1dE#(WM7Lg:@1_9a^.0d
,3-HI:a[SERG9N;U[1(Jd847UgMY].ZXQbM#7?N6KT;cQM\B,:WCN/-d8e6Be-BL
[[HBZ=X58ID/g2>ccI&g[Qd.)W_Ce_;QeI3VDcPeIdJQ7@Uaa930RdQE&.WGDSee
?>NY;)RBfd+U25Z@/P,SPEE0G?D\=\V[8+^I:3>2de,5?4KI)9D6A+:#,;(D9J<[
eQde8MA[U/>)?GF?3W3(c[&W=F26TW\FEJ:fZF7-8<<GLSI8bQX;,/?BMI)Z9]8@
V[eVWGBbW0#:a,Z@;06-&MA8TE0KP4@[:bLg4FK=Q&DL_>ecdVR[FQ6R)QR9YIdT
&T8,8C>0RO1,/DV^U-.#:^U9EA&1#=((AWg6GHH2S^382[P]bT;ITFVJ.eW9)/Y0
0DA2FZ&M=M&@AW\[7TV73[D-,MPZfUM[a[/gNZS@]EJb?aYMAAVG5?YR>aLX.cPD
-+cWRLQ-Q@d/0_]&8(ebOJ6O7?W[-/A[^_eG<_bQ]C&E[^JSLdaI?HfVD?B,g/<H
Y_fQfaR?X<?COge<\7L7]a^]:#Y3dKXIP[P8dZH;2/JK#0D,HH;\Y#.<HVPaNEIU
<KK+5dC.YP,fY5<18aDFfJWC#Jg1J]>M=b(8>OKd[cL<9K;1H84\CK2OWCJK^;V0
fb3Z+/4&D5Y(;;3+=Nc=YW?b<@<FW9@BT7IPNDXeM@9=,gf6VL).9&XN^#OGLLM5
OXA>b@<]6\aWBPTUU<(5SC##K;6W5d-F<&NG)#/KS+V0aB6]+b,GAge(]+V]NJ3G
:Ub/QJ(1c91I<B(9N1I-IC\6EDa:f.,Ad3?\@9Y8OPf_]EPPDPQH(#CT:PLN><#:
V6KGd2HI,6VX[E8BNF^;TK)4=?2>JddfPL:7;V-0T^1U1<Xe/L3DA<UgKT11SH?\
K>X494-]/[93>)RbTR_Qb2;a8d]S/(I340g1UTHNQ;=S98HQd3].(9?+8MH4H79E
&0C@3<C^L;?fgL6ESS.Jb?7U3f5C_:XO0<g9KDN#gCK&@a_94BbZCdL4L,^\8,O:
+PZP(c?^63ZMMQ;g03=^JWRWWL<OMc6;4e+1\:8f7EYKK4Q(U[>UO4;Z&ZC=\P5E
3D#:V]OYB#9PQcGd)6U?FCT0KEVP9YG,OB\B:.<Q=G6B-F8D8Z#\FFN/(;<KJ8.<
XEQP^RED&bTW;>G=K\@gU1BA^UE[0#0IbGV8+f0BY_TH^/.OgA&0D4]M.;^c+^&V
N-7BVG:/O\)LJa-0Wg06C<[H-(GaD-a:Z.NY3O212NO:O&LKZG5CK>,Z4\DFK[dH
=VJN0^()[Xc8dG#ged=D9IXUKDA[5J;IVQH.9T1]IB-Z[@e90/bLLA]eHA__2T<,
_7Yb2V##Q^?+OcH276A?YRMIU>^_NN9c]F,)]a;Vb=bIXd\@LYXCEV6BDTI^0=H9
N1,:W^gKI0CTB;E9TU>@4;#=EYV.Ibc&>ca>)&LCfD8BQd41T+#O:O3:[?EM(fO2
38?56I74B0g/J+C4FEIcJ\cU,PC;:HP--OdJ4fWe97J1N[94F2Z0:>\:);H9EeJI
]RT(cI:W-T^<JHQHW>KTF]9MdM,FaAW0/84gU[?@<&Nd[/f1^+Z,d8\Vb/5W=2Og
H.5WWPDdE,E1V#Ac8GN:5.JA02d4cK:5N/eg9JL(D]AJG>X&9S)b+>:2182LWe@8
)WV+LF7AfB8OKZ2VRPH0^Ped#GW<ca[Qe0;@?Ec<VP\,6V8GFB4#&...dMR;KeG5
F:__M&[T3+Tg+6BL[T0>YJ;SRJ6P3P]bV?6J.J,_g8<B0_^W5K+9[;O8@Y];-KXS
fa)W.O:Tg-e-NO_M.[A7C.\fZ<I>Ef,&:8_dO9Z1b+SOa;NYc@0V<e_C;LX0PO@#
/MIbXeEH<>c\N?I1-&??CRV0[cO-)(<d#T:(0F#.c54EX?_IKN)7-8C>ZdM->;g(
OJ#PYccd;@O?MKS/eV.AA<1TgMTM_G2VCcO?-(T2=O\We\T0cAI7^G.YUP6&+c/&
;>II\2Bd0:MJ9(JB9BK0#GYad/fOC3QLD,X(_ADc5XYb1^e.O0VK@QG(eDfC+VMV
O>J#.V\&OedE=V2VFN>X<)(,.-f/HWY1]5=E;L,#5TN8HNJP9F/J45eM?:^:9>I?
>):E+UR].?I1Ta.ddR_<A=RgQ]b3;)3Q-@EQ2W<bY/TI-#R7E7-9<E=;g@7+4F\I
XN:3+H<VEMCEYBd/bb>8S^OS_f+.e.MP4Qg[;-9.FEPL928/W\P=B744I_1:(#9F
G>\\9^;H>Y\BJJ_9Q(P(?Z3)Zd.P:ZT.6V>Y]9;0O7U+-R335GZ,CU+Od9CL1W,X
9\/SSgIBU4JQARe(g405d\T)9:c#&52N1SRBF/1NfgH;b94H:64E,5+-b^bQKB#L
G]JcI(F+(3?>D&?SN&H9aa8F1Y;Z:AO3+]bB4eLHdO[7?WSC29R4QXBdT.E7+&)-
?:I)f0F;9.C37JMd-DKM^9=Wc@\I[)R(=[<fM7+,TY_U^WKdPSDT(SP-:cU-V>4I
.e4\IHP^3X#g4>^09QdadPJZdSb9P?A.@)L];_fZ:E+<GFZc:[28+^)4Sf-He>#.
&FP\08+^.YQfaKC<Md1D4aL11],dQ//91;XVJ[>36.=fL^B#fE50P0&1#G<AB64g
N/b\<)gI[TeSAKdGKMMXHIRc)]J9M88)XK+]@.TPLE8/,7>,_;)4I<H_@[N9H)O1
FC,.#<b@<UY<WMA;/9TX3;,D=\fLe]d;Z39G=?gL&-f:c2[\5bNb;JLOA2?S<PGa
W:gfDNB0DSMc(U6+H8X7[8\.D0aH>Bc;XP0,C.QaKO)TO0Bd,OZ7Tf#bDJF/F&9#
<L:TB/f1MFAdWRL:+bMRQ<;d3Sc-NGWFDX^Y9N&WT.]9/)\0:^fZ/X)Z5>\-1A/F
&G/UQ4RY.Te(?]R#X.,^dO;GR@=f:4SNd_X9b\>KZeBb/QX2Cb\)P8<JS#G+:1^S
U[@V-0^-ZZfUVfHE=/g>ZWR6?\3f2,4;f=fcc([g@A]#YDC9M)Wb>XY\eSZRE8M&
aNP2.F/369c]O,JaW4K@X828eKdDDeW40D1bC2+U&JdCc7PM>TREcIU>4:/cOQ=V
;DH[aCgdb@9R+8=+BD0^?b)P;XJ81NC,00Y;\c_(5-g@WH-<bJK?V)-E8P,JM:]C
LM@D8O1;ZP@^aN7V(3fM1Z1,b8&.6OXI\VEbe.D8]-C340J1\L(2>\-]J3<B;Xd3
.C-Y\LEJ?+dCA46Z9EgW+6>(WMECJXM&EEK3/11ZAg7E8AF?MTOCac+U?BM@G;2U
/g7-ECIdKLKH6>CE^&F.a@Z#N[S]#4LB<\@##(MO+Z+,(/85Q6V1e?7@<<CM;F9f
IU]Z9167#f7]c>@^EQ;RC&?G8G<2QK#;MGGg?2IPXL=BU]/E@T4Y-KWdXQW1LR:d
)7fLKEZ_[FE:gV&0MRK(4A#<bQe<7#eRMX3)c6IV2c+VV-SFQL6&FFGSA3ffWR=1
89-dJC+ZM&127f[IeAOQRV9a2<M//eJR9ZTRD_52aH#Nb,,I(=?9)J7>]HbA;)]d
2PAR[XEV@RE>aA7=GH.HX[9d6;DWZJDUeL#APN+T<>?\Q(b00fU/.8H536;RgX@W
]Z49f6543g&;5[/g/)F&5:L?#S=A^Y6U<aS0#5NPK=FJ=E^@(1NHHIH1NU\5a+7(
#FFICI:U4Ee_FQBJZCKKVg<?Z[](25FCA_cY7RQB@(IWV5:0P7M(.5@35,YHa,9&
f&]AR]E#LV=Qd,@Zd\LN88f9EOca^eW@\#^@F4W^RY)@d799:96<AN0a0V=_V@+8
7,7[4UBH,V9(4_EA0JXM:PQEHG87Rbe^D-Z+c]+(J\BD6+6W/a1UNX\9@b#PMV]N
c^<R8:ZUM2I,28WE^[NA#33-(cM>W6^]c;T0WYZ8(>^GSYe^bgM=TX3V:[eOaXDD
GIG6&5dDE39OdCNPW#=]@8,NIce^J;bMCfX#OJ^/CBSc3W3>60DF=U7(M:5K@Q-I
4c;d.-\&ddD>(eP3)HCI2=LMg76DEM\(^gY0FCPc5K\8X6NY@#8+#5_8LQd?@G9)
;P[5&_]FA:/+&cP[PR4ODe;;3(5GdBS+I/XL/@VG@d1P]Z?G7<&SN5,=a\.;G6:g
d^8\XFV++E\?T<(M?a73QY^2TKbS9PJWUGgMG<C(MUO;ZAUf?+#46^aA3[E64Z>K
=9/W>GV1)/OU)WEU2)^Y6Ud8@<A#744+;>;2CdK]7USZd<[RI<=J<RbG0Z#/2V2N
=B2RAb/8/HHO@BBOe;MQEe@#:73N&M3V3E]9F<TJOX1EHHH2XE6=.FL2LX:4b,.,
aD).1JW]F\FgCd4e_H&+QLCJ/EEH@9?a8]8<=3-\,E;M(cLV<.-O\ZR78]H.3bL2
M>R/^^U1Yg5^2+CJ/g3LBNR7:REgL9g]d(Y@Y\Wf>,77]:,>0O?E4-UXI91V26.8
7]41:7N2P&;19Ba<[Z9D&8D#)YFGO?OS1[f;[b(HM\f&4W,H.LBcMZU2dZ8^N2:/
G[UMDZ/U,?9d0^e-@KCX0@0XFD2Dd=M,O[+8cZIf0Ze;R.Xf--I-#>U-TQR,Qc&5
4K:-=&WD^7Z>2H01AJV[>H:7=M7<J.M-D_F_+C85EZ6)4ME^XL(Y^(>UgO/Xb/T/
<Ie+Ia7QF\Rc#NS+W880\7gDOY3<@..I/fDIYM<SQ8CQD4C0@b1:I:E[\:0[d96)
D+]RRHU4\E57YPS+H?bV-WV35YG-+0#9R&J?#,?eO,ZQgAR#7O-V>UEJ&a(^I0\W
XCEJAIb&?JEAF)T9-4<EIa@C3AL^d(HJ9Q2;6,VP372.[_O:Ac6aRHSfM<63.\I4
NOa#8E-ST/)HYgV<B=]d=^AO5LIK(E@/9[/&2&:^7HKS.<_0g68FgZ1M7W#]f^A,
d7XGB0XQ&3Cb/8AG_C<7^\5VE-&d=,aN/6XKI/F52W.]@#1I0I5]-0PAH-YM-JK5
aL8?3T-gJ2]E#5N<TeD_BP:9.FHGgL1>Z=1SR>dWGbE0_].;a-2OLFI;2=(R+;W1
Zf>VP)Ld0?;[+@9M4M=?(I]Q:&7QJBXJXYPGD1g?54\K7SR)J0E4Hc50eU9VIUJ<
KF^M.L@5S/J=U_ZN^(3fYRLVaT9U6gFQLed,cMZ6E6UVJOWc2ef41BZ7EA#G]PDb
80Kg)8.[&U#F?aK#L+J[3L2=#0<BS)Q9-6BH\YFeHRL(H7._:.]OJX\]@)HJGPX:
VS=U_IT.G,2R8OaH14bbV;b1ZfJ]03e.;0[1+g3R,T9dGT:8CLaL>7aEQ^[QQP/3
)L/B<Q_X@TT/B&W<4VCIC^=HV1BTF6(cAL.4MMA,@^^.aG:[@8&BR1,)HW[0eBcf
</;>Y\e#Z400VPfNdT872DOOC2A?c-cE=Y^c9VK@OTS;HQSN2e;6C+?.<a[eO6g+
VRZ)6.#LEIaFed[/gQdc-TI6K)AN?7>T-b.#8[J]3PDI.E(2R,<OT)S(<V5.+COT
&?3YO\0PKfQHUJC5\V\&5JZ:ffIL@YO>::O5#^]:G[KX+-A+f\^<FX79)Pg,;e9D
:(T=,>7?&-Y?[AZ9-8aKWRZHeLd@X.dANbBO#.cgeM(WZdSGF:9a3GR[WORa\1K(
:_\>+8+e&;)K[fC8FSC,BGe:TX61gWHf/Xg_+JGNG(S=T3IQdNOGWI3ONUegS_aA
A8KOaV39T2DF->BC1Y_?@/]DHga0bf];f0>3PQd_VD+\,LP8VN,;3P/f_KLD9(3A
:X\g^CUNL=GW+D=5?[Of?,XRA/gOR0O-M2Bec;;G.ZOce[.?^)J<KE=UZ-DfM,R5
?;40I36IDF1(a#cF>S(R,.ROMHC[B:,E)=DYg5Qa-2PgIWZ,B(Z+\9/5]2TNSXe]
EcGe<U4EU99QAPOYe6G#?^cZKZXPTI-P>:[.\DR)MKd0^?a=1K#@+DUCV#8-Z#gT
4ZYY75X1GU>,S(d_-A.,Y)g0e3:081+1,Z?cF/>4V4.K?AV-O-.:-Z26.TbD9&>L
+VJ::GXRg\LI\Ldb;,<Y_](^W4/6V[^Q22-40@Fa-C]A3H5>\a3a5gX5>Mbb0^Yb
XLH3GLA1.ee>)4<9LI-S/J+M1+.AH/9C\E:Y6G8--+d1>X?Ug8/P4gfFXdOJP^9@
9W\Ta?1E&\]+<&KeR6_b6^Z+g;9#^N\OC]Z;WJ>U+c2=,MeL6K;A48_(?VDDaPg1
MD8#e3=<;:F^RKBTB7O.(TQPa6V_YO:[#+(+G>S\g&g[32L]?/Y.#458K8+HA.:8
E\,OF(_EG.(H]^YSS=@C](\ENf<K@D.A=K8LUF#J.gWAY,VD9\@9IZb20_LQ0R=d
Y8Gd^6&TZC?Q?LGW6(>WS[d(;&NVBBAQ6R4V?4S6&[LL=.>AK5=41g4[52R;dEKE
75&OS[/HeUUFc2PX9P;TB4e@KL;F=T,+dP7#FTX#;NF7XQ.H9,Q.8,VE9VB-ZRbU
8<MeUa(P&T]cf2A;b_90Q_?I[cVB6]\aRJ:5Y;a:STERV,9.36=_5MB;M#_QLge\
YDHW@DE^17MY-2/PZM29e#\<ZB7HB?<d_;(+PNe[W^ITI.ZZOKSc(/cXaEI66#6O
S;00@8H[<6(E4BDfb_]Hb[#6+WJFJII0/<I1(gRMea5\:b6+]@WM+<ZPSb>&]c=#
fN11A\P7e:5608dA-7B[N?gMRD:2TDQ,FI/XI(GK=7H=1:_^[+LK=HE9Ug7#[Z+=
_60\B/4U<4WY@8dWLV[TfHPYYCTg;S@K[JLCN;c7:fEMIa^,2I44:P/a2F3g8BJC
baAQX\GW\G@F(RcSMTDaUfEW4?EK_ba8MUgEb8=S2?+E-4(0Lf6O2eB7A(gOa+RV
ZfHR].XL,NfO1]\/5f01094f/:QU93:^cSTB=W]4\N5^HA9?6^9a8TVKa?,]F36V
dgLCb,(B5LfVMVf,<4fO9Pb/>.IH.OV_2VJ2g0gW.XWIW;#O^[23K<>6Pd^PXIHb
SCF1dHHM>McMae7&GN/3b&4<IYNBO_CIR\NT]?OR](g<O<(&IPI_5ETF[U+1A9C:
Y9=,=Wf#Q9MO?D3/3FI&&PW;EHI2T]LA>U.6SCDFf2(2g+[6II/>KXFMY4-,[>J4
3GbD@gLE@&,-.G-&0XAINZ3^^U?I_QSOI/MMDbOEDJ,9g6YBeJPL4D9_QUCL8X.:
.WIBA9^?IgB;\\2AHVIe>VYLGR.S/WL1J,[N:>?]7\.#-H1H:KT9849X)=/>FNb8
^Rc9\T/FL1\0;(D::U8^7f?0a9,T-^X);XJ[Zg]:DP+[@aDZBJ5G>QDO?dFP:C-)
de=0Zc<J=/#C:g0fQCbLde9Vde,S]#+VdH>PCX7ZS&[C1KNb+?d&?[:9eG8N5P=P
0Qb2>.>X;SBOBH=(ANEbC08Z\/HcZGTUc&P80B=HgKCVTRfMS+3;@f?PA&aFF]<P
+]NJT-JKZ#)6e>_EdJ@\MBEVT638EE]\D,P6+Z:IS><eBaQ<g.^>Z7;VeQ@a^>V)
Keg5N?Z4\cV0Z&.a=2S4T&@X8LEY?TX@E2(a&M#1e>?b-1g__QD&UOXAJ\,5IK3G
&IcZ&]K&Z[49S<gdb<&Ea?P.>D2++NJ>HZ]LH+_B+(_6C8^,2Ae+fX,(DU]Q@S(&
5J;^DUQ06/L<])6--(d/E^2]2RG,/R+@6&a^T64WfE3-?BLT13KQ.Gc^DWZVTST1
<4YUO>F<C#fMVG;[#8+-+8J>+2_]gBTcYV;ce.LaB@]_[LO_Z-AWe<Z(2<V;=.2>
YMKA094;J[gg79f?4RE#@;4OIG_4BagJ7M_).\@QGJ<9dN[&GaI&C=..8:2QfLGO
\@STW?HU;bAW&ICf#?+E;@)VZDB;V-/HJ7T=S-V)/B4,QO\R\=7fE20>a=cGa/WX
RH0T/&\9OQ/dH_1C2@eQ039D)\b]8UFVQ#+.X(9U6MH.8cfR]Y<=?c@.G;6@U#0L
2[[UV6c.:ce6&;PT&dAJ1G:f<g0edP+a:BNRDa[9@<gdd(ZL=]>CIQ(2\LCLc&DY
,,_IJ\AOcM\.?OJV;P&1QTM(aJ:S\0]b?d]+HR<Fc:DL+d=.B#]^KA8[]Q0.X;F8
AJO.QAaLV)@O/9VROQ>+=UR]#17)FgCg^a[_&#eR)FEG3],2Y3ZN=g@HZXE<:ad2
R#,aF@7EJL8Ed4AA:GUL[Y3YGH[@JY;?JAD-I;E2-Y)AXGX#J=4\-^(;4E<UHH+)
UJY4F<8K6K&=5O,^H.M^H]=F;3SK3g^SM>O/:2Ye>D(fbU0\H^NQbRe.8=+#[,M+
^+UQS\L6AO;\[2YXUW#@\)LV=Z)^e4_A^_;cf.QL.-S?P6D<c3T)(P]B5OR7&2>O
/FQD:(eOTV#[T._:b.Z?=KN8KBD@P4d^-.(R77eR?2@:2Z?K^2SJ24QI04>2[8)-
5I:(\^>^Nd0L;K0f@@Y87&;N87gf:2M?]/NY?C)T[_KM;0f;b5=Gb)N/#Ba-^AH6
DK.DV_33((dV>a.VG7dA)+2RH^+gWCf.c#+6(?I@=GAH4H8<J##,QcWUWDEHc8@J
G_XDb;Q?g/A&=f3(g(>.1G](QUK(5M>:.^KaTc,E0OM=#YZ?WPI_>c/\SQF:?_g6
Qg]@:2>=X::[<V6/OPM83LG17/&Ef5?#^8^./63d#RV7MQ5QPXQK0S]X(-be0[10
#IL+7QVU(B:5[75-Ag<^WX=c@;1RKQ3\S,b?]MWMA#=AQ#,a[;Z9YK9X5LB;BWO3
(KKEKbID6GN2=cAT7&\0;9A<^.970>Z[PAQ0OS[8T=VD@=T\W9A(#>G(=3:0(0[3
<MOT3Z[3.-Ic8_2bc[_0(JAXDDE5(I,G<MOMSfHYU5QS,Y^U<X9GB<3aPF)4Xb@c
0H>+WCHZG\DL8_+E;;KIEE-4<a6gb1Tg3Z&bAX&:X\;?(P&;FfSGNUKR)gaNcYS=
fSK4J)gFf)EDc@KN5-48I,2&ZGHEKcLE\b(d29PHGNK@bL5W0:P\FU=:_/,PbJf+
TN4Z:E8KZD,;cHODT#<CDd:Y)RcC>K;)bQLVDUO4(+:E6)aYH,bO#aVc\dD\:ZC#
8EPcQ7UBK\E^J2VZABHLY)=94=J+eS143R/BSN55[[?Q38L@gfId4[X)OcL[(4Cb
fT<<?-@(b]7RK[=Y6LJQ[9baH4Q)H.aaE>CMSGZR,-5G8,3NRLB3;5YM-RNfYOCS
JJ3f-T#fPI/=IQ-\Q9#ULg[eVA+AH4ec/3FSHV:LM/<4a]JP?>aabP+bH]A?V&;c
.<>HTId0.ac)+GU7.aS_GESb7X:d?)Vf[>#:LY&Y?g3]Y=eX8d#]]dX.?]+,d=<L
?dOMFQ5.B7FDYMg0H(-6[I_/&-(XDGJfP#4,@7ZaPNA3MTMbM8QE^,fHBE>^BdN<
.S2V>&1<MAJ.1HMB5c\V+Vf@Ld03D@;3c]Kdb+6+P#b?9OLNTU^Q&#\6.DBCP]I=
0ND<E+-bU5IG2&8HOBbB3OP-0e;;;4/J9XJQe,4MIY<>)BQ3H0V,:#_K&\fD5#GY
?(465XCAAE-B+80BF#(1D?^_c&8Q1+WQ=S&4JEM&<0N&]^WEcHE1B9-KDWef;<Ea
+PLaC>W#K1R1@WH<ad/Q@8^[U8UfJ]QaFYAWgK<<#6\3B521R9fO,QB^1>bU7NTe
A7@S]QK4[)8e\>>-LSO&d&9<IF[<geHIQ-T(BI<N(5SaZ.L/EEFDeIQ=afdBACJ8
IHd6))>#L16fJ:(1DCcKRJKX\]>5]abOV_[f8,?gc,I\0VH+LX9T&VQVO^AJA<8R
<?CI_;.;J@M)V4QM4:G?DVRJPFZ3V&&3DSLSTIT7OW5;(BCFfBX-_)9LLD(<3ac_
S?^Xc_e#J?,WHNY]eRFWN+XO8?_:K/A7d1dPFUE]HN/@LJ2#@T)+-eeJE78DE3#[
NHZef/&E>1<\C]8P)W:B+K5GYag.I&;3-9#+=aS1?C?23J<-KN5A<,;ebCF//-GS
[A18WA)<P6HdF0CAd5I=#.63,9HdBNA?OYg4.T#:TS:O/3<1fI?b.6aLLaAJ>U3K
._K2]S^UNQWX+gED[:]V46BOaO=7E;0XHS?c.9JMDNHSI[.8=>W3[MXfQ?)1N9L>
+Y+eMQC#-\JJ@XZ8NJ.[?:?\>)Y=@;-.;>HSDO6&^^gG#D:X94._c\J3;(Y:98b+
^b[Y1DNJ)##?bVMd=1egR=L6FX+BWaeGK]=;^AINg6_6W:P5-A7OT#g+).=@+9Q^
.HX6+1(6VR@c8(#XI9;(XY:aV:Qb;F74e-O@.?D;>3L/M/_aQ?XTB3@(]ZBXSYU>
3P2O](0&?e^>Ue@/e<WBec-S]XcgR\/&G2Ng1>E:aHN9de\-Z[M=<O>:c\4gb7V7
\K]P[:F<JT:[S)5PPJYGP:9,c>U83_?,I/R-eFC5>/AJM7=F3FE,,K,0H11D?N.N
[?YOB);[<4Va2,eH9XCL=6^WX0c(I..#L7R><P&S;1ET-;,4NCJT-A-PfcVHWURC
Y;</F(PW]7-)Q<8+/+1:V4.FUT.9Wd6)4F?6#9TbT?)1;0B3:/RWQ/=;?TOHP+;/
HDPfKV1dV&D&6Z4G@_]2#J[Q_S70cE:K<DT[FJg9eHL-[F]=VIM9RHCZM0+YQ&_R
c\,BVY<fT?<OXWG.;SRK3YZD#A;@fYMKg=HARV1-fP,&2H0P\9RDEBCGY_:RTC+0
/S\[OC]J;SY2-P2e0[cHFNRV4S+=[IgdGL+DI<ggd]..8a6_@9P13f70<5f(Xb^N
1YD9b?]=\W&OL@SD4)@aCC70CDKX@gbI7G_;_YS:L@83Z(VY0(29A@cC>>7JfAAA
>UQ-L7U9K6.P9aK-C3F\]9+X^AcD3@=O-72I[a=KfR0QdW_DMd^V.(XHEB73JE18
.\9>1TbP#;B=<A,g^QZ(K)722TMC-/U)LE;HNYX)FXY?ZI-==\X?1,4U&&b2AH-X
.-:-2CId?,HH[5^<K0&f8L^GB/>,D/?f-J(X\YfF\Bg:U@):W25]<A1GB4)d8VHL
J(ECd,#7VQRYb]],ef?ZDDQF^MZXNKG,@(@[<Cc.CYN=T0ZC0G^+&b6/(AM-c910
>;1#bMMf0R1NAaMI2S(UCQ[_.=,GJD)_[cgI&P3D5O;.@)#CF2T?WTI8\>E:75,4
fg=T860APF[EdW8CQ.Qd235aVA+O6;:&BWS+LT2WZ,V@+68ZdFg\dN[0NcNXRE<Y
P?<Z.&a?^>ET5O36;7LX4]<9eT>K7cJFD5#CR.a_^]>XN=d4V.S8>-eaHg,a0:34
3Z>dVEZ-@c^aR?/I-4UDF,=edKH<CGC[7[b@AEE2936ZP@Te0XVP=LAUgH^0.)MK
Sd&cY=I(LLdC(>FOY>&?bPUS;T=#HMI>(64f-bbBW23H@02?<?gQ9;T^LWH-_8C;
BZ96#MYbc]Y6R@):<:f&E8/,SgRg;+CdV<K8GH82_0DSE5;#66S5QYOd;^^b#2RG
_efA-Ag#.(S)DYT[d7g\?A@H,\b=CL93EF_PdX)d,-YIg1OVY6A@9Z+d(2^RZ7AH
a+(IM^+47O@DG7@P=,@g&L>P#-_,.@.[#84RJPUBIOZAD2(eYQP\3e)g1aLR_E1D
_[LXCT^db-6::3_eCg027YID,<HbaIb<XdYP84&H[T,ST<CY9fR/H89VcHGE;PGL
<)?684=\2T\(^ba?2N7E)[H\fKEc-)7Z8H:MOKWc@@KYM4/BT,EBMc[-ZQ=(;]<7
VUUF@\#>>/9@4Hg,.^aZ]FMSO+.DNeC776JaL5VKM/U#c&8OG]-AM2&50@)GSeVF
;Ic_Q5dL?fUd0Y/Yf<S(fC(V56Ya.FKY8C3+__HF/-J76&K72Mf2\MLS9OZO=[TE
HO><X?H<])I,<?TI6V=-@Dg>P0Ye_Y(S65d^70;]6SWSR]6D=?F248]GfY)WF4RE
^+e@Yd2DB^SR@B^^[]=eWOZ^,RcQ6DV9==dg>P57ES:^3&=.23@[(HU0B<Z;0M[K
+c)_DOg:EQ=Fc])@)<EF[EQCdbY+Cg:ND3SPMD]]68)BMHRa8=>ERc91Q2PfPPXc
U_<]??b/J+BFTN]\<YGba<Z8L#_7\]++\1E;GTS?@)S]CZa&>P1gY^f6XODP7Xa;
A>b?QQ:>O#dPI/<\&F:VIFT79=T4PFe24A&K]AQ-e&^8U.b6GP)Y-)>Q]B]?eTOe
9_.EWQV-ED=^Y-_2-e8BeZ.HQZRGXa.ML2Sg4^EM#ZW>:7SeBB)<gcP6.84(gY3_
\8V+].\\a7L4K.aTU6#Rd^7WAdWI1+G.[DH9YLGP?SDUQS]>]_g48bffS>P?J,4>
]VDD^7_g(W)B+H-cF5_29Z]-,(PO+@D2fQecXXK_:;J0X+[IEK5;WGCH5:.=c.V4
@BK)A?c9;NI^/,.QV^aVYQLH)10fIJ\7=#eUWOJ4A1dC1),_dR+0QJf>5>C&/VE)
ea^e#cJMO9,H8(IdfcNdT=G0:EJDW4J8B&C9,fScI>FRba7))49d&JUd&S4),+N@
N9IbMADAZ,J6U[MM1ES8a87REDJP,=(dK=PS3HR1VL,?^-<0WDgA/>=&GC(Y#Ce,
[;;>JD@fKHJ]8#>5T,WTK_449C7&c-e6USYN^^IOgg39WfNFd2(/B7<Bd9)H\,>S
]eFQY3,Hd<JaVZ>G8C;E.&gc>+H<TT(2/.+:@24a/_YIZ&;Eb3HUU@GAN^M6[N5G
0S=g?XS(Z^A8+=f)E,_8&P<71-VdYISVaC4a47Ne6]).F?K;1)W0T0bW<0-?g/gY
ROHV?N[@V[5b=FA^/^/S7R>J]5L;;GZ<4[(cYP^#67901HB?JR_OWdK,V6,\Xb0\
>CJM.=cRd47(a6XcV+?fU]2I39f31#)4IHc6NQ=:&C:&9PKbc;;N3XS=\H[O.6f[
)FG(1OBV9.g[BX#>&2DE(_2:f1\BYEb17T_G?<292R5KYb^<M@M5g&436Sd7eGG;
eEbgMK^4IEXTYZ:+\[a8@A1J_&W74cJ>J<A7@A5e.5D,G,d<G11;V<<c[7+I&ZdE
ZW1eW?7UgE/S_RFH()N-5Wb5[E6dQ(\@\DM7?Ob4dc\RWDJ=d\RNZ9J;L(=bF?T^
V1=aZHI)Ng)+A2\0KWbc?^VI9OB&4<_2ZR5?:Pg6I_D=N6;9SZ5T>MI7dI9R??0L
^,b(68AYCXL<G_e.TFa]8@2RR2MMR0eQ8.+?e4E&1(MWYH);U8Lga5e[5>.(#D+8
:c?NG&BbTP6&(WE3cN^Q]e@=fbU&Q,ND?-XWPTPG+A).QXI):Me2PP\?U:-[LW:_
f[/?NgAVdSX&+$
`endprotected



`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
  `svt_vmm_data_new(svt_axi_master_transaction)
    extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_master_transaction)
      `svt_data_member_end(svt_axi_master_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();
`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

`ifdef SVT_VMM_TECHNOLOGY

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_master_transaction.
   */
  extern virtual function vmm_data do_allocate ();
   
  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);
  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0] bytes[], input int unsigned  offset = 0, input int len = -1, input int kind = -1);
`endif // SVT_UVM_TECHNOLOGY


  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);

// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
  extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

//---------------------------------------------------------------------------------

  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
 extern virtual function svt_pattern do_allocate_pattern ();
  
  /** 
   * Does a basic validation of this transaction object 
   */
  extern virtual function bit do_is_valid (bit silent = 0, int kind = RELEVANT);
//-------------------------------------------------------------------------------

  `ifdef SVT_AXI_QVN_ENABLE
  /**
    * Returns index of qos_upgrade_delay queue which matches with
    * current cycle number provided. If it doesn't match then this
    * function returns -1, indicating current cycle is not suitable
    * to upgrade QOS value. 
    * If there is a match that means current cycle is suitable to
    * upgrade QOS value.
    */
  //extern virtual function int qvn_qos_upgrade_index(int cycle_num);

  `endif

`protected
Z&Zb1N8e&3?b>IgGaRS9A3LTHOV=3H=gE-48FXcdZ2XWN[:PAJX37)+Y25UD?E#(
:[BHf?8:NS.b,$
`endprotected

`ifdef SVT_VMM_TECHNOLOGY
     `vmm_class_factory(svt_axi_master_transaction)      
`endif   
endclass

/**
Utility methods definition of  svt_axi_master_transaction class
*/


`protected
a>g[g,)ROV<7OTZ2YPeHG=M)P0@LCb.N@T:<N0W3:0OgQa_77:gR+)ED89.A5YBe
8,cP4:@&[b-e2^3K=NGEH/J9#6YZDTM&/P)#T4OV0&ORPW&S\a;HD4;+IN=VT?-7
X<VGGVEWJ&N]^JfGY)D]/f+7b#I@V>)6/b)^0.P^RaMLOA=IGXE;TM-DA4Y>6S)A
fE4Ya=(=FaRgXY3?Y7DL3-;4aB]P(=+F#2QBSH5K^^c)][B06]AW]50[Y3,OMHPU
&T8_bg0D3/?=VXLJ.D:D_TZf=NS@ZAQ4P.;OV;4+(0IgLHHMV2IPZ01dFH1?d(_R
537L#Ce4TJ1e>ee4D>XT0QHL&7^RE1Zf+:K_9J-KPQ]5Z-A.<F:a==<bIb4a,)EO
.0J(.(RAO3bB_L?b3DD-Y4b8,O]-DbQJH)NNG7X#D/+<?8:CJWK_-(4J:4dda]+2
J<HE;GX>51KNUC+_B[&:6:KSNR5@/G&ONdgHKf:3LG.T\5c59GIV3IJ4EO+f::QC
aRA@^4WLOYJ05=(CNH-HFVb5dO.P+JJWVAAT,7([&e@[(L)H=Y,VJZAe-HGVH0WE
<OZHT2PX)2=Ng(?]<P9Y3QEdT6T^:P/O(eNU:/EaV#8[I^^->.Xf]\S.cD82XId/
gf-MS#B7^aHVF<<KaEWgWBLWaPJcXFUH]c_1UGR;;QTY+J1M]#M,._:/N^CHab]_
OPW##^(\2<aA:ZDb?AQG32@IL?<W)S@Kd0Z[1LHU\9@^Te&3Z5<S4?,8&I]3T-#I
R+CZ>d4O,I3TS[8WP>DJWM&9BfK\Uc9B)E\6ZfZb5:/7e=GLOSC-M4,6^KBAL14E
Ze^/BB_.#KPL?F14(SJ?P,)g)Uf.0A<dB?+WFBfJTWR#56CY)e#d89gae\gf7?=/
U/X1A9^^+c1TdbdSK8+LYNeO6;DO+8N;_R84OQ#4)K4MZ\A.-<U5ab<T+<,2=8J-
1HZ,IW4;/DNDPB&F+F&?gS6U#XX5-VX8^4b?@EbLN@Dc^C8DKKN@SX#d20e_b;04
H-+M;7WY^&d,ZE7T@KIFQeDOT]/NN):6@D[=fdbW?^DJ50PR@>6+R1U97[\K#0MB
2)0O(@\.<ZYVKUKG^FMK=68XL7659KbQ(8:1Y4eYKDQHOa+P_C@-b26+&/K70I9I
W-HHf(Z0^<?YU,AX]\-T5IS@ZHcRI82?-;9,S^7g8F9<MeYUJ05P6SVB++QZ_fA;
gfe76VFR=J\-5<G])Tc?0T>(HTP&5SHHf;Q6X0J0K[;.5VG#KF_>UCaR^#PP#ITI
>]N02_]^KWL,J5NV#.@4LL3-SD_c7BR302GZgY4\&NI7@8GFFV4a.GI0;\WP]OG]
MR2.RKcAO7KDFf:419(C\&2W)#O>Y,(dPc0LL:+K41H8XS4HZ<QEKQU[(cb5^PR<
L&+\J)+AA4eGJT[^P:(]^:L\,<ZJ.Mf+&RF:QH=#E)XM-FXcJ&:59\/D8/19Lc.0
F(O)VNSXJ&N5CS2(EC@NcTgWIWQ@EPc4,V>0<>3?(a,XHG?2HIdRBfB[5[J.a>7O
1PM?&6<_0#cE:;_7PA#.N@2QfAM=3Bbe/+dT]+P^A9I:EcZN8R:S\DJXH=:T\T.L
b1S;.\U,3#fZ0LHJ8^[8?e\a2.5IYZXDLNbZO9U&QH<;]\E0gNM0V-#=e33GOZU]
QZOS?A6&W:/AO#P:GS1&b>b.dG]Q<2Lf0>gd?(X2Z^Od()8ba?9+,TG==fb\DCTP
C5+<fJWEXBI6,_[X]dP#aW@(PQ]^+a4b9#JXZP0G-&X+Oad5@JDK)TR<7,\=/[3e
fAI0M^;7:g.KdM.+ggaZb61A.##V3OGUYW_ZRfIaZW)VDX;_b8[cg?6B(&]&>\#8
8,fFcc^e?A9\9eIZ,aO,aM84=?b65CQI4-6T/:Z2XB]A]_+S=,.^aX/V\eZ,&KUE
<-<bVQ1272MD4DDI)U3f)D0_#OML9/SNa6([[N-c-C=##c4-TgG>UI6QFaG3[>_\
><WC4&U-:ET>D.-b9JBRVB8,J40<C</)QD[&91ML#:6V)M_P]U84cHR)6#XU<S.E
U];d\V_d&)=]&fOEZ[UCG-1T,4C92I[&0,ER+c?<8>cPLBTB,F:[M-PZJNVb]T^;
M[fXWK\D@AO/.BG#e<I\g=1T7$
`endprotected


function void svt_axi_master_transaction::pre_randomize ();
`protected
)F<#]?6;NQcUL67DKA?;e&4O)R,?1=2\_XC#S04:4.QTB?_E4LJF()COZf\dD9]1
beTg]+CG(]+]U9QQfDDSK7U0FNDBE.^T-0O&JTKH7#3>Y-/c0(a=3Z/,gdaA+AGU
6O=W3NWaBV,=&[79R-8>#@f@Z92.\2\>e9&FJ,<@cO<=>W=/1g?;X\+/If/DbfL9
BYKGMLXVU2228@aCISE)<H526[fIC14C)+[CP<;ZC;,63LYcN82EB>=Y?+:a&,4T
AU;e>J;?LO+1aPX<]^F/M1O?YA@U>)R]6]0(U\TWJ[SH/;+PI0)E7Ge#(XIGd-1T
d#Ve?[KS].9_=W,cCKdWf4cQXJcP.&ONRa&&:DdFga9bMgQRW_K7]HDd5);GFaS2
ZbXBPQ.C:FU<(<7Ua@7Cf>cQ6$
`endprotected

endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_master_transaction::post_randomize ();
  int log_base_2_total_bytes;
`protected
?MeFgB&W)0+X[bSd;5XaL&23T9g@>QKZ/7IMY3YB\;BRDL?cH=#95)Y#8GgO=@(Y
CGd;1J)a_e:+a(Bb0S0MGG8)c(P9/R29H[40g8UKB:S_Z4db=M83f6?U=a?3_d5@
:,;F@P3e(/FcKU2P4[Y9a;D=+V[LGHYXfe6J.eZY_+g7<\425aOC,c9W@7)a9AG1
Y&-&ee4;^U1Q12Z\;L-TH::S>&\6e;-]OS#B7:4d?SX9<L/-JTY-M4G^5@/7^5=J
02X5L<SK)9UPP-#_f7_]/cI513S2F&+\_)d;SQ-]TDd1_?a06R>,KTQa\36Y=LS<
8.KdNQ_V>[I)2I;bHYYC/9fTTNY>BRQb+5J-7E;P=D>[NXbg:\W[?:,GP/\[f9gL
SL\:+2KLF,MbZ@A^@LRc5@:=8-3FU2Ba&dB#F8<6;/bcE@f[S+LDd>C9_VJ8V6NT
JKgcXDYgRa])JV-71:Y+2(9S]QFAX8H+W=P[^9=9GDO_b])AJ;[]PO9:<78YTVg#
21d7WTELPS/14YKFUQ^(H#^\+?^].=WA:bY[\R-+^4;BY<^aQB+AbL8eIJ7<ZU60
;8)Aecc.6O,,X:C4#Ie,0[DcMV9-.1K>K>)YB_c=L4V7/D43YL#P]&)B2YOGVadC
0PH.?d_WQJJ7ac@/D-c^XJ_XBE^.Zc2S5M7;W0aB(=_>[+[02U+C(G5Q/GgPPV15
5Tc^WIE?gI>?e>]S>-<D_HdGFI&<3Dd,FOHL6_GETe_526&b?EZLJBHBLD2YYTb5
/-#>6J[#BA]Q8a:#Q3A2d7W6JEN(\X-&;$
`endprotected

endfunction: post_randomize

//vcs_vip_protect
`protected
9E8SFQ;A8@C\I8;L=RM4EK+&&6^bZBBS]:#R>#8QDQ#]XPg>PG[X,(O5e+8Z&8[\
=@I+M#]+AgNT1XY4^.)\dU/E<gQIX-03B3EORA(6MgIf#5.9]8gbI&K0R91Ce7QV
R0WH,&bg(G7^[GE@GHS#R4=]2_EgM_.R>,JC5<cF\B6N6,0]V7U2@6L7_47;>M;7
a;GGKTK/eWg;I\I._K6dD-9eKA50c+@(STP[1>?&9R+eNV&SR-T<KZ;,.NV@WCd=
&H0)=PYU#3;bQBG0Z7_a8K9T#)LZQH\BgBVIXWXLLQ9^4ZTOa@[?D01V]\(7=IC^
BZ8GK]-,Qf,P,6\FBE&WR\U>:AT/XXJP.Ub<GGeHCH73\LW<5^8Y+d&O(TF:DF=^
0?dY@?B\ag:Na)ZJP7R4[d:Z;U[P)9SH=X]X/)MDP6[UZ2d#NJIG/)0(f7N.>@g[
?M5B-P^+V,4BQb4O3ZG8F&E+(]Z0BN036ZNT)\GFCNT+0D)BFHF.<-Ic+:5M<KSc
KH.JUOA3R).a,0I_0Q7F@Sc30AaD_ZbA:PRB?8E8M-e3L6LQ3f;Y5-Y20R/Mc+1C
4(Q9,H25&gg7&UPZHT-XMfP6a<Q4PQS)W;[JGPI\-,CaB@A>5d/))9Q(FF9b_VPW
,>aY\)BaC8Y<+3)/;YGGDUFEOS4PDS@YX7#(4M;T-<O3gYAX,A),=?7PE=SJJg.G
QUAEd&\_fQe2SJa9]Y@E/ZUF^3AS>fF&<PE4>c=Pd/-O2]/JO-T=JgBACgZ[Q._O
Db=>G3T/?g(=2g+c2EW;ad=RCf_SBM)\;$
`endprotected
  
`protected
<M(K]VaW_T@c7HL3=05e@&NQ_];fcWYM>d]^YU,Q1JF1]^LQ9(7K0)[<G<cHZ8e/
+ddODF6ZOb6c,$
`endprotected

//vcs_vip_protect
`protected
S;M)[.65QQcgH:3&AbS>0K^]EM,0-<6bIOI]T0YZ47)&3cURQ?G(4(8T?[3?d0U5
K^A;8g01KV\0fK(_UAA74+2e6N.O[Y==VJ2)d75R,H;I]\[7>-cG=Q^:<dTQ.\;(
K?d(Gaa)I1<Ue48H=3/:A>/T+R3T-(c\JE^\B-X\8P_7C#GEK7WC;^5;;X10WF7>
b&#5YC5LD/A+N>W-B=D<f31(:)JG\_XB7CE0>2+KLU7WN>#\J3@#eZ;O\W<e]A3[
O=bKP^.(g]/8@KJ:KdSF^^-(1?9@.?a,eV\1Jb?fE;W3E#0PMY;,0(b&QVcVDEc0
L+@[MP@(Ue#G.(e1)&MR&\#Y.()KQB8c:T;@R#]0Z+-aAW,/6\0b>>Ia()?Ca&11
^R0#O_5#J4ZG6TU+RbfK<SeIWWDc=2\3MHPV7JcY_9N,.W5&(:,Q.K?M7H2dfNd0
)T8B:.,K7DLJX9c6O0<N^5^JL\+WMW=N5DYg^TVQ+-_UML.N,O_E5#N7.C3Nd/4K
EFQE/I4#TCUS1<UB=/<]d1PP=>EG]B_0@cTe5LZ]^LKb<LS=4e8>\fg<2]AS#B0e
P0VX_7E.U<[MJ];OF1[]HOHdbPUKdM##\f3IT;Ja/0JFO&2SLaBUUSOM&_D5.L-Q
Rg-H#C8F]7CEU6J7bWK-;.H[dD:Qa-RO>0f-gQXJaU<&4Z2&fg:/1b[G4ZKRf-?^
UMYQZ\L(7=O6Q];3]D>XSJ1[-/YTHg;eV5c\ZN9bW43U)WMRgA(X8B4RN;g&;/+A
G4.V=)<a(0JBXdBJZ_;S):],f_eZ\?B.:@7)>VaKX-c<\+->M.C/A/CK&^@A4S?>
0<H:9)84#_:];PS[D2ZWb)3.=<1#,cM1BQ_[-92E+]#X395RGE#_+f[3MKb=4bH7
J2Y-3\9KdF8Bc2.049,V>9S>UUA3b(>&##9M;J#gIMTJ9]MU]fUTaR]DgLC>#:]-
#.C2E9E\gKO]1Lg0G<?G[V2MG?a=0N#Wa+0\#aLHN(P6E64;XR?1Q5LdUWDaFS07
J&H3)[5R3,+CYMd#=T&M(]?^1XD@^-47SU4RL(;^bXJIe9VJ_f2GSS8XG;J9RO:W
9XWQ[aQ)G\Q)M@eNb8RYW5C8^CO5E.&UF98H0&0ENc.IK(6\9635YPT+67./ZXEa
\f+HP5ca_g9WN)eA((KGA+G(U\5U:Wcfge:E]]?=1?\A5JBg[U7]-C.c^5O0;@\#
M?QPE@+N><KII>7UeBF+9\)U;#Kd90F13+cEbRf_N>@4Te1\-+.9T34.7Fa+EYXb
g.1?M>.==bJ+^E>2/#.cO,.9EfP].96,AB/K:;e=.O#5e[F8H\CJT,VR,(eUdTM=
f1T[?8Q>HM);g51)bUMd)RG[8^fZ7W,5^+H;LBM::[a_O>CO2745fB]<]Fc[6(VN
NNX815Ma_6gNKD59YE#cX.&g5(RcL?Ia+N>@H#.Q8?1f,B^QO\OU@J=LC/1>2I]K
TI?bX@9d<B-J:ecYMWgFOU+XOD6G7^]U4Z]_\C_6g-E/JEQfI@>f_L,,gK\:CFHc
@S,CSGKHAJ=[KUE),W,_ST-KgaHN80CW,aJS0M33LP.9^WZW#0O,&Tdf4>RQ]@:2
R+LBI+^#EK2=DGZ3CQT_aRWA,IQb6EW<-AD\;3/@N?>J;)F1@WbT(Le0^QIQd4#I
RD]AEXdE0>].OY&[O-@Xc(I=_CT?O==M[7DA+&9KOQ7OPaT4gN_KF^=W=N;5M>6;
dBUR&+ZJ2W#MTf@<_-0_7]E\@eL_=J0S[&F3Y[^D+DX;(Dfb.IMWc]QD5;T@b2_9
B^<HHX>XfbG;_9,\=:_OH=-Q5^B2[^XHGcF154)K5_RSU&GA7@JC?WGL233ddOV(
JE-d?=)dE0Lb=?ODXPY6XE;&:a;I[KK#CWX#H,0R4P9&L6L6aRNNX]J7QA.d5S72
2TK],ed.]#=6>a=NRH1_6N#<,G(&R#CB7Ua9=8=-3I^F4DeH+g+()G6_3UHZR;+e
9429H+XXbN2cAWXWS^:g2#@1PcIG-HFA:6C3+(]0UH68JeW=I(Y:N52E06<gbZ<J
\6S7VA,aQ[=eET.#OZV/ZNfU0J719SLQH79-.]=9J^P8?.9Le/dMJD@S3KDM4.QD
OOBJ5/;57.c(bTY<8agR7Z0SXY;BZ[MZ1fT8JFLc\H-[:(:]K]=X6^DePAb,+R>b
X/Bg=VI=Eg6W]dG)CO3F#;F8e5R<091FM?;Y;,7]5VP56Ff^?bIHZ+QAI3S-Xe-9
9BB^GPK3DIYb<_Abf(U\4_\JcU2e/+YM)c;HAeE\\d@Z1Y^b:657GXEP1,+>U9P[
:e[GAD<bgZRa>6&CB?2BJRgQC=LM?^/1Ea_LZZ56WT<a&T0W(1A:;g=N8]1DV47X
bHB^Bc/@LQ?N?EZ7BU7,>\^PCH@J=8Y.a],E1T\G#b9X>a&^-33\[/DBX.aT:]8b
/7cRYR53Y>U@W8f<WcSY/V)F^]9\VTeE5@+NC=\BT4PUN:)d9(RT7OO-LUMV2;VL
V<4.@#<D[RbZP3>8D6d)67ZX,@;]/,dU5U_C7d02H4g-Z522U=(0?\M;XZ8DfWEV
(8./=;&\5G9@_<TGZ-<Pf(:Ne:UB:#H/^N9QE3RI5_0H8:07)c(bg)HXSOX0#V+=
QPQK@O7LF#R:FNKc82Sf5.]9-0L[1SY=N1T_MeD6<(_>2SEc]<_HY[:73+Zb@KNE
OWS]8@5E]Tg=[7G8M7/R@ER<;P?S3#Z7E@OR?[QQYD1QfR\IH(L1?9]93KL=+JeW
aXdCS/;X0?L\^@YGI5-aA)gV3Tc1dI2dPT6E).KO:I;1QD_+Y64cU7,K(K8(O//\
MW@LH;eU@DLMQWgC;IW^DQN08@?7O)[HFX:)I4/Lg/Z,M4Q?cTE0L@:fHF>SD@g0
^0.KNN(QSOa0]NOY);LX0&QaPcL,GA-@0Hf:B.C4aO_9[8.+S6MWdY:LR3]_8L?c
H8\f:+I4A4HW#LJH7G)B8+F.-<.6e)2WIPIL8P5JRF-T7Dd@8&<KLVKfPOe<.OLY
#PE+0))H)NgFYM:CE<@.\.dde>:OGF\.aG#0A2TSeQYddc5b+<W4YCFL2[@Z(2bP
9]106PRGN@X]<[CHWPedP0:HX67R6C^K)2eHaKAEM6P?M2EN&9/F]5IXLLZWSDRP
#1BX9RZV9B]a_Sc:I@>4GYGZ01cJB@^Y@O/:H^Sd7fb^cN1SM7/,=HcT++b>AB#1
0(2\0X:W9c8&e(7\O>#Of<Ca^:ADVfM.WHe#5f^AE2-H5.UEOae)VP4(O4+,PURX
9?#<ST]3.,CHM8^6GfN0SU5UV+1XJC[&L&\^)]b\EC^7LJG&])5OL^0,gH\C8@gc
Yb.F>aI#4WCP1#52I-aRg:DGD&0#J&E\Feb8[;2I/bg_15YJ7Qa/e_=]deRDa0#e
\M_4[16[3+&_M92\eG:4:O]bS+QCKI/6B-J=/dZ4Z]B?(6F.@I>1ZgdEV.<.[5<I
FOV0-]8N\]]\E,d=6\8M^#P;c(.#FJM9MSabJ-X[2@2S.4ZU^#c^ZcX=48SQT0LG
^TS)9B1VRCUa]P<X0KW;R4/ZOe:X3L,:.Y@P8GI2IAX?H2(13T;;W^I?&TaD)QTR
;fZ2:SWb(RbP2+dQIe^0S<27.Z<=-S[5P6M]WME^393)c@,2>Z^K.cbgB/PU1[,A
_^P:&JUZNH<[JNB_DEegWF?NUb_)F^8EbU/d,aR[O2Lc8UAB_(UCVZ4==+-SY+FQ
S#KX,<;]TA2^G[>JZ.IWS\:(<D3QWKRKZ7e=PZ97W(K6+SBUJ#C)YSdabgHEe\(D
&:,IAXB:L/:B1:cS?U<H<:E(7,Z.M0YN]=A8U;3/RXBHDJ(&P?,-\(d]@]5?>Z@J
I@J33QFO^07<eFC<H-TRb7#d)_f)5?_K9J+-(],.B>T-^G-\E/Z_;0]C:eed1b;R
UWAL9-D@RHd-(-@_[Z60I+6R.L.=QQHXS]\G>g.)OCLB9/,<Zf4P73NIdOB>a)B<
RRZ#LHF9&f?MccT##HbF^6gT\4:Z5Q]HM3Ld0AVZ>dI0F9<0<02a>3aNG-0AKBGa
IC^MU5F:=H[JAaW0Gb8Ta2@H33Ac(8<&fPa&E?<fgFe7RQU36O2fDCdVDQR(JTT)
<DDc+MOK529^gP4Fd/N4XDBOW<\:c?+TZ5U<P;ZX979G8;BV?c]DR)=,9)cT.09D
[=]N,VK(E8^=B^:C,C[J.7UEQL?<?+d&4g8\[@_YU]D33WgMO^B&?@88LK)A,f9W
ZA>DZ)3ZCM6.1/B6b:J+#ODW[dVDVd8_IG17:DF)_e@L(.]ad51bW?YSQIG)Z038
Q8(gRd.+;HT8.Q&<9:0<5;g73NND@2H@R;a6)U]YQU4;62L(])1S?>]T?9@60ERF
LKE,1=dLU54XK#7<4eL4;P.ICR]-C^g,PeYVN(4A7W^UNU(^.,?K=g90f_Q.C;-e
#-A-^8AH)Ob1^M0dRR@R41,gL/^A^,#MSBEUaG:F.cC8?#LfHF)]L+?LO03R1Ka4
f3B?/:C/eHdfH;-ba;#PTL&:ZYPbE[Uf9TPc.XZQ=a5?>7CIG^eE;#E8=7QL)X_J
KW0b0I<+0:M=dQ/D_?0fUGMU-?=1#:+dbf.@L6CNMN^]/1>(SadZK6F\bf?GIFT)
,]ELA5^ZZ.37b1fFA,BcF4,efXQS/[dX;<8_R09_aB7V(4/C?0SV>abMKS0Le@cU
LCG]FD+2SLF8<[.?Re)X+M/XU[^37?d-5ICbZ13=a#M6Ig5JSfRZ<9C,A>.8@c=V
_cQAe?8#5-1GW4,FZR>T(+ZK?gRH1[.fb<&TUd/1>Y&\VQPKJW=TD^HND&@QLf9&
#(2@+aF^-0/074BA;C@/9P&7DH7AaAQ6X0]<9a9EIDX_-^cf@K\YFVS^WAB901=F
9.(Zcb@ZX61H)Ga:^;?5QP;A2;Z5.e1gQB>Rf>N;MB(\?PU\7e)CCbJAcI4N]S5H
,EVZ2FO0[\C2N;TAf]JaSI#Q),-A(e]-8N0?-K2/^\7Y>dg7:,9gE0cdC]ULFXg_
XCFZ4fgI9Ee?\@7/GNfGR^4Mc>W<LB7Y2JeR)gO?Xe]RLWV8,6YGV#>KbNFE\:J@
W#RK#_VCK4,1eBH4bUY7XU5QaD2[#Wg7(;M,V<LJ5_47FaO8Y).HASKSf.NgK(CL
OC#EXGIQVJUgS/J(HJBGb1Tdb,S8O8-TY.>>MOU@UAL+8\5#CI&_5a9PW:8Q.dRU
-2TF\QY/A\9\>5->6[7aO[3WMUEXGfO<4>cC7FdM[0ORAY2JTQRMX&[Rc>d<+/4D
X90?F^,>KY+4OU28WK]YT,W&=3WG@H\U.D8VKNJ_c7UQ64DX+SKa\)cHdd/S+6OO
:F/5N??fcF[X_W6_2dFP+VgSU[_NCW7,N(c,OB.PQg)G-?WQ>=53>G&2O^)I)I.;
VM16H@KM6<SMIc6FeLD>PP1=IC:c61PM2YVN3?N(MF-C+K02N]Y+U6YSY.d78XP-
4X/bG95H8Z7]S>.1EZC02F0ONdN/5H[>=a\13=.V+GKY2+6C@a5GF@KNf:g)@:;L
\Af+f8.CZM=dCU[T^31^bEE][Y1&]?f.\.=#98X<K;B&;9]/e<D)M;)b2Nf.bNYU
IT(K&I2aE;//OPS-0EH7RIc4NV=JTE#<e/_6+RD&FJBHID&eB_dOa@7J(DbJ37NN
?_Z<ZRT_KC;>26f<XRZ<Bb0L1?84)GT)<Y1J;G4X->0g(I272R\2H6cRd\bS/A(d
99[X+)G<e)#8\)#+K8(QJXYWHZT5,X=5a)V\)TgNcMM]-W_=OaJa38g3K.[=]Q;+
EM?>><7b,G_5996S_,6F<I5;,AV<0gC31GK:dS@=d/FA9L5U>:+18B,/:4:0B+UQ
;,?S/E&XF0R6KS7PA7NLe--T+KW[f22XAg=b]R6(Kb[KRd_>.)8/e3T;#WTYdD=I
Ga[dG>EV;&[GS&M_1U5GT,]Z9,aX-](<aQK;-:<X](8#BB&211\S7e_9<,+/9f;]
PL]2;2ZR?[C,/USPF0eN,KO2&2)&,Z[_BQ#cEY]J<?gJZACS[@R+4FBb/A?[5&=,
DQ,A8IFWW33_]7eQ05ES9g=HUg^NgbLXYWZ_W9d)H>M?9B?2S=]_P70STRMG750I
dP__PQ4ZA52]bc7IcMK@_HSWG][=VHH+7,JSM=]UY+_cD)6TYY4WORVC[3(V]X=2
e][Tb)M7?YMbRA)D:Ab?SU>\32_FOWFMX(=[^4<c/6.aC26T8?6dH#7FSf^d#9Uc
Gdf<\3-f/Y-7S).<@A#&d(4g(K//9JT\^(PA/D;J9\F?ggK?@-98:&/2Ze7?F+&^
L0@P/UT6PCHC[7JBE&1.\ZGFg&87H>;X]ga09)1S?^APgc/20KdFDQZYK#=f&5TH
;>a?O<9c5LW0aFcP&OBF#+X-]89P=CebT(5/0C@f,=#H>-#YDb:OOH\@H5c38IBM
_Z422&c-8<>M/?dCV1A7(?g-G[=Q0+c+8)..>B;M1_CECPIW2,U-aWD#ggM06@Ee
R/L[e+K,/cH/Z4)KDVTe4f:T?Z]aMNDf=.VGdW5KQYDCFU8<MZ(YF20Zf;5GI@+(
T9]?9-=T105#b75UC0a]>X,fB:QA<N0/)D^&&=REE(e8,A2LM0\f)?c,;E=/c2MH
aT7OK,H]?@b=U+0JJ0=@A&6cK^6\V7=CB9&:(AfB/T^5J&cOS\@M)DG2gU.OQ,G/
cSLCe^T?X5MZ0)]7,()OdcR(f^+WEdN?P_K=Q]/8H@MXZ23&MGCKM\Q78)Z5/WA_
NYd(@ATR5UDMC0\LC&BGV:N0I\];-#GDE/1Nc@(.Za#3D]aW:)^=M<:1?cA<U/-a
5-BF2F[_PHCU\TCX7YSDXKL;\c9B2Lg-fXYQbdX)add)C)UJTgBX>JW8S7be5^5M
bb:dT-_:X+6CbP-Y@a6cLG&A??8LDb(#B9L1.GG]IQ&3,E<B2(e^A=3<dYZX\?1<
4KLL75dBb@\EQ7204UOd&CB@Kg23gWd\M\/#V<4]K.d+IT^B^512YUT=B(0O^V]0
5e)_PC)(&/D0gb:KIG?:fFTZ@#2P:b+E0ZYaI;VJX#;H)JTaSOY3JPZV+UA#Y[O]
]fSY.:)FX1YRR^FXCTQTO_QaF(??6#_+fF;P_LG>fdUAUg8)=:.g@KCO?O]+NfD;
)<S5Q\,:R7V)HfSWQFDEYe0Q3/WDE/0/^\L9Q03X)[;IQ)+T55-TG1\0;TIZ+bMW
(LV9DYDe;.2)=D(Ea6[H^S_@HNB)/W8IXWW?P8R@/+KXZLUK#b_[Nb&AH8WM[_eN
C6ZRSNX@D9IP<9>/<]e[D:G5VK3?ZD>RC3]?DZcb)NFOSZ6LYI;YCWL^03(d;3Aa
f(G2NQ#AMCaMJ^#cEL#8=:JGGPBb\2CD?I^=N0T?^0d615KP_;H,e1Z=JU=)P_MX
<COCLQT6IA81]?G.[^YBH,:dI\._aLKaR)(HdKATPU^?&b_48CCX9;21fTb=5@J/
a@).80WFg8C74GeNE]JT,2]cg1b5FNH^XC6aXGCWPeQAZOe51(M.KfTP1;279Ub@
&g74eA49V?Y+7.Q2<f],IR)KYJFDf5\TC=>UBQ.XP>X]<_g=O0(.=;67598PT;,D
TcNCY>2X&>[834_FLPN+YELa23^&J,Z4Za=\:\>U@//PXN0LO[-9;UFMVE+=)cMb
]43]f=KeP,CJ>Y4=Y]W?b,MX_Y,8De>@<cCbL01S<,&<5;?0P]8E_S.5ZFSDR+5L
[<3:VEWHTR>1XUF[9&\&SbQ;OB[36Rf0/ff9fHR:d?MO&CFb@3?F;W/e(NN(XF/C
I[ZaM<:BH,;Z)&)39]P2;]HX7Y5\^DO@]/4&HfW84eH;f2O=<>=UI?U8aJBeA0;2
6;M):KUc_OGZ]\9.K#W+UaN4LZbACYWHH:@cFKg51_YMR\5MDPaM=VWgSGg3d#cf
dcb.9c:[&b@<?=f:>688MA^_:J&cHV6N@fA:W-6H\;&=<NX0;+R6V<)(B0BgbgZ(
0^;XD[IIeN@bC@EBPaU;XU1+2HNGZ&e9fFX\<M]T-3;->2T7MVS3(0+UFD8:O?[;
NW-BEBU)affHDE:.IE0T=Jab[G]I4=W@-)2NUZ7W\@N>J[TWc784FP2fK81aLM:.
J<5fHb4H8)YTc63LX<^.\G/8;=)[R=.9@,;8<@b;FW\-<0P.8YL,RK<cPF^H^N0G
:A1[?+afd>_=6&b4<^)K#g5=UgdcKR0IH3JM_8W0R\RRCKXD\/@N7OFPK\V,6HM;
GWcg-ENf8))53&bM<Q13VNA.1K6dg>FDPf7^OLgb]H/;BNe1?:Lb@XS.52ZG,f;?
#+;243aQ/72</<LfR?G6c5]cQc4+cDCb[K<8KL&WF,7EgK@UAcY>d2&^;](4WZ.J
PRGCagg8^e?:ZQ.:E.^#2VbCf@65fTHE^#bbY8R)CS/ZU]R.NBU>+KDZI?J28e\4
4fc-a<f1C@YNb;:B_\I=AO2ELHH&cUP&#1/a_@+J[&,L,b&VNQJ-5)U<0C2ecNWU
(J__N52DM=12[XQ2Fc2RZH^PX#(Y,.L[AH8C3KOCAC^7J.#QAGP_?6I5RE)/dVF#
]>[7ICP.-F/gYJ:,9HaGAT^R.f,GQ-+)f^T@8?;ZDTG[KB05+H1.RCa@L[F&:6/>
VXQOA((dVA.f\G]GIfB#BK6<;VU7e]KG&VZLS]>?6TW[,fUF96eN<6/KNG.X:1^,
LC?0NITN6eaTQDP3E@88W6-P@Kg5HXc8W(H+KgH5ZRTEQ+(^gHW/N@,EPK:1K-g\
UN\T,/\S@WNAZNW9<<D0^8eE&LV>T]+6c<Uc8cFCD5[POe?aHAa)J13V@KXVCZNb
&dHC3eCc&&L?>:1>1=Eea/827P1VV7N;5>GM?B]?cX-Y#P44S6^O/484OA=J9Q0T
/T,IgUQNQ-.[Cg:G4JLLJb+3f37]J9H><]E.:N+ca51eV5SR>]agENM2F54+W#/2
Y:80b/2X(YNBF1QQee=H:^S2SARV//WBO&3>+8McMJ[&J2LcHeEPdUT30#8U\F5I
7?5D3FHZU_ZO8,4<gdO^QLBWa<dH@8.R;O=(:Y\?YD]_JMdDNQ]#?+D5Y8G_51D(
e8&c?+81KO?WXP[IdZX8X<AM&-g[FeN>^QYL2NW/ZA1a:9g5KP[<BdEPZ#M_H9-M
(G)MgFT4S2&>eQQM0H9&B_\K6\gY5B>?BCF4RYa?X5:^JT\S?W5aQgEW[]XW2;@(
W9=-[+LZTW1I><GJZHQF5fN+HYaX\SP2e[&)]QS(Q)Lcd.S;:K=?Ge6P?WL)RHOB
SKIK_=Y.C(E)<;:&:JJ)<0;=V[COg7HW_9O^9SW^HGCf3R@A3(e84WB@TeeM3A9W
U]BFBfGF0[]K7b\>M[[?=V:f(a=F&>c].D]@I2b\T-HQg+6@J)Z<(X?T;A1#8[Q#
YMDYCGPL)9CG<<@0M71/4.b&>T;<E>Z.;2T2b4\_X>=0_^?/6b<P;&P<WU6CO,LY
5;#\HQW7E&]FdVLPFGZaVW:[<IR;\LT);XYAc=LGC9KcQK-d;@TU?B<FC.)0]#X-
#2#KK28c42bH7W6c[CPC@LG<?1O_Y9^^,DA<B;bSe:eWHIH^OJ)P8+.Id=7MA8].
BH,BZ98WW7=fLM=F5-Dce;VNQc:O+>SA4SS(QZKUE@=>E>7c0<<VFAIL6,Q?45gN
2VIJZ,JE;Q06FX[BNHV@,4LB/D.YA+W(7P#78+_,#JHC7YS>51\UU>R<;&OQE[dE
?32;&:)-DN8L.Y>?69_9705?c(IKWGRaab,4=eICK(C?7:#c@gP)aKU&V]ONE_BX
N4D4_I\^8Lf&E7DH)C?(_WW,<N2X>NHCT/_(\7MT(8_JFMW:9X/4AC<GI>3H[5AT
/8Y[1OAM_/U=C9eae4Ff(C&Zed<#GW1&H]:O=?DX:65+TSBG36,>.X.0d:JBcOIF
]/)DF1T&>M1I).D5:c]CXcDG4KfCXK66>^Jd@K+fG[<Z[CaE.W-3(#+->82@2V//
DB#0[/dH[feF3CB5Mc8NG51,5^ZEUPIHUb4_?Sd3g8.XMEA&XG@SS0dSN@])@#N=
GMfc&)/4&;5QEdB7\^3OD:ZH>1NC#]fRUIcJQ8G:TB\E+4VX\PHS93I=9)^Y[Sg5
D9FLEc;,2+-Ic8Y6FCJD5=IOEGD[]YO^1d=DW<2@a:,.LR#1DT22U(U5eF+,&T3&
?>#\N#KP2d&J@4;-PBIV5aZD25b^YNYF=BPGRD\].6CZ;-\2(W218:=+E\/29/H-
We5V).bDVM[:+35Y^2,XJe_QAJ7TEQ>>#K,aeA136[ORb=KK@KE-7Q?\b,VS.M80
f&U^(E:e>Q=gYJHX[LQ3P0MM,+IG;,@fZFOC1,1)X+U:?@0)Q5#g^\4BM&Q:M&A2
B]Ue=,5)FGK/SF&T(:R6BA6&E?QU^FSe^K#&Z8\3G>M4I4Ob&V(9J^VLEO9K8UOO
2^dU/4Y\+>De6,Z/>:PY:3?-d]C;4[<CO(D&T3_+gF.)6(b38E?7MFK+-U9,Y:0W
UDc//[#A+.U>^N,ceZE9^-.Z^\9FL7NK0_O=8>#R[g2=<GeV,6f1PY&b]&bDGL\S
Q@CEQ@I-gDD=YUXf&]N_45D_cMd7N30TWRG1Pb>W>HB75fI=db^[^M<[Z=)26.()
]<[20GYVb3fG.CGZDXG3Y5/@-Z(;F]#P@9^K4_6ZS5]&?60#(-Ha76+:dEP>Q@Rc
?@8(cfS0SY]8L\C0X)aZFA.+1XKf2FI.M:8GG67T:INJ>V&;K0SU.+7J:fW9).a1
&_O0HN,.^FX-T4PL&=NE:a6(R_T)VCVXV;)DF76HGUZOBFUf@eKBgN@1I5_JaJ7W
70d].d050M5E4:MVNR5]A),bb1=PgQD1Od:_+5J3^P,UM6IJfQf+FGU(+TS^a&Df
:9SWSTL#33B+@DbM.TWJ3BE6Y(<8M.A^OQO_Pd@bbT,\QJRG?-I]-]TK/X43)7S^
48N8ROg]IVCPDM,;fG3JUKNN[F_:9+D22B.UbYK;4^G:;UcSEGEK7SLYK:Z8YKPF
,7,H@-<#X0\A2e;1?Q;F]/9ae7V-XQ=FQ(;KZ(KT<U,@dJLZB9JEIYMZ#JLF1/0S
O>)1#:]BIW?)MOK,gVYUR3O9G[H.4\2D7MLR^9KBZ\LHWfF^a7]\ag-.)HB&IXWP
UEM7T8PMf>T&HWC\0_Q[OFO;_,37T/JTZG94VJ?E.a9N:V[-YfP++T0fD?.W489U
:Q2N,M[(7(ZF)Z,9_<5dV1^f#AMB\_OZQIFf]eY@WXNY[5:(0+:4FFc:S50BU7#A
,dXJ/c[G<[dTWc#96\8^UEG)G)EIZ5[HaO)D#)G_1OF^XPGRE+LQF5JZ.#L))[Eb
2;4U9gNC[>8<#Ea/.W+b/7.f:=HFA7&;9XKNKVc_6_?QWNcAWZ1ec_.Q>W&3SKMF
De25dZ-c;b32-gb=UEEgG[H2N#/(N(CZ:1PK>_f_^1/6^+J<&8L4+RB8#+QMW=]+
36M.25CG\LG0J4?O91F@77FZ2S&B@P6@/H)eB/[/QK\PJIf4F]6JY9)b)RJ3-g);
P\DM]d>W(d9\EYDP(5@5S_d2/dDaM;37(-G<AGEIN:/^&,SaA2=R:/4#Fe)3UM:d
Z?Z#BbAcf[VATK=-][QcT>63-UDf]NcT_K>[CQ]X(QKcf;BDX,AC1)=NJQf6)R-S
#^F2T:H\U9PFe/&[TR2WSFd(SLK+:Y52aaO?H_.A-&K[g+J/]aUURU:,<(Y._D-M
Z9N)TW[PA>B_?#bG>VDDLDbDD#P^W2[<G>LR40:gQ_2&BW)-JY,>5/(4J5Qe47.D
(U#.KdTLN2H#@fgD[Cf8#d@f\\<XOTJLDI^RMI@N.+[Kd45LdM<;8IRK4Y54>fP5
eSP1<_afNVbBW,J-5Jc.)8J8,Cc8VL#V2#DO[)UaPEY6ETS(QIBIfUX6Q+LTZBJ^
8SY@]64b,+f]._Qe&O^GFWJ[JS6L@X=V[X85H\TVTA=Q;#a/Y(WfgZ=/]/L1T^P#
f.D5(-RQOBP?6?#3N2SWFL(64WK477>;Qa,IZ&<^B12U-CKeT4>X8BUSMZSe0:36
?B3JKaQa(]\G70Yd?.55+Pe&?5.VYLE5W=3g[K<#N9BRYN441K8eQF\KF,5D0K(W
#KLJZ5=/,.8]H[MNF_R/_#1LaYQASc@KL]P(T/N8+>C+\&7.=_1a;:1G?GS8B<5T
W2/G[^.,OZ+M,#RDLQSP_)E,4YFAO)=OJ5@MC(Db+g^^O-L(:bQ/\7adM&X,358g
]X^dZJEb=)e<??.E\bQB.>2MQ.#a8GA2)7+&X693KBJH-JK6;H/+((cMJM;ZNO-1
+XW;B6MY(A<>O^HdX]e;\c-f5D,UWU0/TOdZJU7(8\&S-G,L([ACDVbRK5P42[);
A9Q/]>;CD3^Rf0>5aW\_)?>4];[<]99d-28?T2ee0WI&2HG/)([e(>)06DB(_YEf
\15:NC0:+G8R3BCOQd_@[;4e,7+3J]+8<#QfI<B9#2):B=OYA,U;M0TE8BbcUK(J
A-S9KPKE.IIF3a60,K<7+>T.+D=41_L>.R),NO_.ce/g(:UW[-CXQ-?_=X907&Z#
H7H?@1U-?#I.0NJX2[,W8G(Wb\Ud^#ZbJ_7ZS]3K(4VVG]3FK)>)TfPf)Y/-8BZO
@WDI15A5<KWTX]fbBbCHO^^=G3CXOB>[R=[@)bS#.]LRX,I>(G83UZE-JU6TXfCD
?#+Bec4REA_:(KM-ATf7X(Q.@Mc;Gf(G>cZC:Nd::XX22D]e<[:R\_@.,6@M2ZdQ
CWKf#LgKN\b[V&a[KS?]Xb/b4f7[X,CFdT-LE:2?e86MO,d&^X2LQ=:_W9UM2@96
9B01geDN4FFVM4C^TC-ISE;L9eM5LHb7EWSf::aE3D>NKB[,I7H+\DV1TF:J=,U)
YB#bd&/?UKU.[X)@]4bg36=?9Q1/cf443^X)U\9<^Y86B0P3.c;&78dOH(2N8&^1
E12[;A&44JIVb>?3J]?7>@W+DS_)90]4Ve33^\.LIKC0#I//W>_\,V)@P+Qb3Qc(
<Y2KW:&A&]]b.;aHVg&8b+6<J/P76P=fK)]7:M#-LL+ATW+LN1#U#K/C:2AFZag7
^7L3cR)C1DBda/+^(DcIPHB&T#9dL>HULa+H7AAF@Y>d7].)]KRRC=L;+]1<A1VM
d>BdQHKN:6:Ve4=H@\fUW/IH[,F4SG=7]3(RC99SH[KE1SeE4DB,PG8Z=PcET2Q.
(WFY,ILdE]#a,)M^8Ud4HGEEe[(V<ZN6dW4&1+T4Rb-HGcZ,DKJJgT(&SYd]W:GU
LeN8PW0^\9c(X?LEP+.18&V>Q#&9#,LME3HTT]fK5LR;(Df2:a=C,[=WRd.K.\^C
&)#>8Q#70_;\<I+4e)X]TISZ?&bc.FbEE3.ONGK9\\^-@TCRN@+6TS#CF#5bJ,^M
NJK@NJ\MNG6a-@J:-K\JQ@?-8:_0R)8(8TVV=W8aLUHMYWMd04-:_U(QPUc?E3H1
DYA+KZMV(22V:Ff<U;DLIg5RW)CP>Kb1&B=S;9XdGZ_O)\;dKXIe\7^g&W?4ZC2]
4C;\#acI3&&UPS8b8BSI;UT=WK)fQ;dP<=_H>^_a3bOF;8Ma@Sg?EV1?VU3@H\X1
8]cJ\6OF?M;cC[NURW6LGaI4_7]PCN@37?agXW?;S]>BgV-\2,P_8@SF3-UY-F8G
U:X_.S_B;/)\SBI)+K:f61M,^4DQ]?GfTTOH9+<b4,@NOQ1;<S-XF+P7QI=a?VV2
LX.Q,0_e/2[AV0IfcU46AYS,2)bJ5@_/E0J?E:FS=af-<b^YP8DIN\d\GA:g<E6Y
E;YB3HZ/,E+Hg7S0F?&c,g>F9FJ41U@D_S0W_>CRN>)6+Md6\&[_8,Z:#B6HgNJ&
-KPUT83eQQ9PD_YN.U.&ID?4Ha@UNPBPd^:B)Q<gN5T6NZS37RS0QQ0P.,Z,RD]A
L<7_e+0+bG+IBN:U#Q?6g2;5>(#1@c(ND@F:(RX1+C.1WAY--PEPQf]G)?]/4RBd
BU][FL(#,/IKMM4dF=Y_:C@YZETMM50T#f\,TJeb_#>PL6K^C-ggX[8b@X;1[,>B
=^K17QY0PbR?-_FQ(],H&\^b_>[4H&.;?<c9_0PQN9Q2@0.?L4NWL,<T,0B[ET/\
4TAITC\^Wd[ac2,W6(-c8:A8MRZeW]e4gO0]4(eVC2cM+=PcM]5.ZQ83VM@d\e2:
XS.K]N]96g2[);82^QH2@T\[.06M(gI(#HK+0\6e>D\73A:&f3JI&6ZRE7XC(.T:
47\QH<X<5026?dW?HE9YE1U-ZZ+b2XHZO2O;3cY_:D-9VAT4IO?J&1^#MV<TCG8\
B<+7H+B_)[KU3UU:./ZIGY)O^[8NV.4&1)^+D0=WAB0CK^JAS,0T^?F0fT6P&D9#
O,)\KN#FeKCX+ZV\,@f@\_[BeQJTKMKMP?BU=F0AC_6L^f@/2<R,\ab7c-T_>Q.P
(V^O5c))CN)]X+<?Pe:F;U\7<5[a(71Y2cc+K)MD[(PDR\ODFg.0>JJ]>I,.)&a<
Z,H(/+&,\RH3cQHC0@GIHK-@RKN+:UVb^AGLHF?4YM=MBU3521dW\C=#?+dUSH7T
M](ecF[WJF96NA?Z4=b8FS&RBIU7/_G-bW/W9?D;B-S0W[ZYLc^<E5B,?PARU=U4
7_T]D@W4=P\FVIY1U2\g:J7P;d05;.G#4K0fU.Te7A(fI<+d-6FQZ3GHBd_A@MHB
YBd1]JPDV=Y_:HI]B.CD4,;?(\0-HF:4fL3ZC_2&;bUR+(9Z74#(G;8MP54fFI7P
XZT4^=&:SZ6]gTT@UE]Z+VXQBb?9)dF?IQR941A@MARN0baKY?f9ce)H\EId9KC8
/50R4[#WK1FSS?ZffED-Uf:+,]ZX0RKbGM8[[4UYWD=/SPd4ePc;<5V.&KVV6g0b
Q4>MT;:^;[X3bE3F45&8T&O+-&cF;PYgcFU\+W(#JK=:U=+bcQWWD?aAd;(IXfF<
<caX?U?8D7HDRKf>Y6DeW?JZI4Lg.3[1=7]TQ68L\NN)Y#EDT(S.2c-&T:JH^,F#
a:FeNe1?Of/B=.4e1&8e0CdEG:E<=(4>fTOa1bdg,T;=@S[:ZR1;Y]A-3bf=VLED
JGG^R6+V&gEWa]g,D]0O#LfPZc4L1?NZ3N-(I]MR_?EgBdUZ?FOdD^\NVb_92E1R
[]B&b9IYA:dI6E6SgRd)afYDJ;\/5Eg4YcEK/J8TAU9A\TI\H&GObTdLR8&f,ZJ?
M0DUgPgFe_f(IBWW+cgTe#TFRT5;&dT:3XY/N+/;_Fg_4]JY&PSQQZ>H9AZG8ZD1
X/>_8A;;JQ6&&ZGXI1WA9U[K[<,9LKdA;=9HFc1IVH9aI@IK=LZ_.g]N@I39@_@N
/188EaQJ:0Vb0JW3@\B\6dMA0,#Vd^?-GH#1-[))_6;cF8YFOLUF_IR1-:W_HABZ
]9&GF+I0caa?FL1@=TX96.b([68@XN4EW<8\)W[d[A:8F7TR(,ZWC:82I2MSRLa0
L1-H0)9P-(a)NFD505Pf_24e(UdN>OV\Ac_YU7]QGg@M7JIWT7d&,e)d.<]c[]QX
3-+RUFAPOXA#R/0^(/V16CXF2[8BK47_g3C+P1+QNUc_\f>-VBIcJdA;G9NKX+Pb
##09Cb3.@INbJ7aND_MC]UggO)TR8@(P#8:0c+R7C.3WRRDV0b[<WD3#Td.@R3O;
QHMJK\?@HZ11?D>EWGNN2V,?>HZBDCYd0(P@L?+Q7;SKWF/-MSGaYF4.T[L&-aa)
&7VXb9a8M8DAFQW17<SB^99P),W5+R^QAX+;8R+#&FA/OG1Tg)JID#;C8O@]+U#\
M571/IB,KY?@e7MRfg9:eed&.:19ZPE<a8GaXe6P9/90C5d7+K9[]6FDA>+P?/@?
a#:f.J.:./aIX&#W?O\_3BY5L4W.Y/VS+Y3H.@Y.8#[-#]gb_O9T;@Y9b&:AZ)cc
Pe[_9d=c2@OK&-?ZAa72f[E(/B8/1YD9\(1<-aKQ6Z:Wb:NRQUaES]D(dKS\@(e_
WF2a7H,6W\Sec_OTIGC/N5M?A[VcS(4bEMK+NgaGR^f[79.IB8:<6;,KYM]9:4Q\
J4>W:D5>2a5_Q)Z=fSW<1C2ZJOLC1.#:EC,G4.]8F3VD0S3:W\SCDOcC=1QM.MWN
W/aH-Z9<?+NRV4M,HE;cgJdbT77T[)&XT[U)20,./Y0@S0FQ#1HP/+A_HZ+NgM-g
K\<9bB=:PYL0A35gS-7#,BGBK7P1X5FD,]gSXZAF7<A<@/Xf3cSPU:VB7C/,#&1d
Q4RSK_2/IT\;ZF5)PR[5DNJY?)(#-:_-&-B^>eYd>QeT9FCN:1J,H.g?3/U<UUC[
.b-==Q>1a-H;R8?;U_6Q_7FbLTBNg#_#DEW9,VdR5Vc-,If2TAdefEYY;=_:K#f7
.AZ(d]YYB#+&G>KTKd_9d@J[5=8A-e.@7.>A@S)F4HR6&D2?EUPEbW7-6gI<>G(8
M6BCEK?e7aL1WI/4W3M;;(aGO((5gNANNQT7H2^P_^.;/K9a_Ne+TJ+)@VgFU\)N
NdC1NI<4g=-g5,bWI)?ggE1B/L1C7(=E2.G-3MU(AE8Vf0;?<OLa>47G#H3/Z^B0
TQ\+44QQA>OX>AKN.01K3H>eREJ21^C#UUa?Ofg0A7<,3/B)Zf1M00\BH[]V01QY
gJU]A9<WPd4.<DIeY#6:KP/aN]aaXDS5A[DW+e/EO@EdO24d\2Z(1f4bJ1NR)7QO
-58S?a(&Y6K#KVcNCc<P=32_[[0PH#,Fce4dEW:V)HBFM@=M;XH=3\g_(YD9H\g7
S73OUR0<>Le(US99(?R7YJGaYIfB4,?U4UbSYRT(D.K>34K]M++_1R#b7.6[92V6
C0gd.dTefcN>_[e1V^e<SBQMH+)-9?NM=QZOJ9gd_BJ1E(3NOBNS6J;cN?1^XER.
PM8.O2_;<BGLCI0H.X1-\M-X5C;S.Ff#S;P<A9?cD_-9cHacL#SQ#BX-R5A^@O85
,;82cIK\3NdEFcA#PQYU;OCFA@>La^F._8Z<BN&(.HR?5-[BS^R;_[[@g:eBF9\@
&^]6_bc]T4+F])6BB)E=cC4&=+I58a_/5S<]Lc-PJIZ:DQ2aSTa^ad2fVII,N_X+
/W=1_cKB,&T1,;S;G^S.e)-TP9<([VP@HD<\f/d8&5?b&6C8V&3]V]N\3&A+Cc+2
V21-:LP\(PHYV7O6/a/04C82HRA,R13JZ_V&Y+;#M=2D,BI<(fT-;^KJ.QL^9.N6
c>8fM4WJ/_I<f([E-RRKa_X7WA&\c/,&.T7-]AVbVfY&/S:DKQb<c#W9Ea<dXMBc
]P5UV=NH-+[?I9-Zd1K47R#=GAGgC7H;A7#1D/0D5G=[HGMZSN94V8&e?U(e:,J&
3.<5?A::4SF6N-MNg]J4R/I^I;\+4J>D;V/HD[ZP3@XMC5\<483T:E<#^UI@Y;PU
>L?C>ef1aURUZRO&dGSaJ7_d+&A:I2#52gVPd7[(ZT#Ad3Lg-6->9^e,J\A26,16
U30+L9/DV?CR9TCg.))2N4_99N=U.V@(&N#O(WEZWB?(.AdRQeRZO?gI6QE6;V:f
B;7Y_RF9#e^CZDENQ5[C<]9a?OAF[BQ:[1:bDE>,ge]6RHF46]L#]?@8-R<6/OgA
@aJZ+bV4gKC->P6BTFQ5V6-B7bO29.^<<S+N0BC0-Ib7_+C1&<d4Y#I:7DD1S8&f
PE9D/&c<6JGCN950b,JDG:]-]Kg<B\]/^6XJO;,^]#2(XK+7VJ:<^EO;5&W6[FUX
dX0Kb7J,-G(]YC)8:;bg.=_Cb7]BcMg7A=?=)(JUPP?;6C)T=1dR509&;-cEa6IB
<+^bbAC^SCZDFE37NgEU-_;8(Q,L,e2\(3)LN1_Q-W@/a[FCRQFH/G(F]5<7H<L#
K\GI^\9IO2+-58a>Y-\Kg@70G)B1^,DE_HfecaC(4fM;NY7LYZZ?(g2LH2P55_F5
SD+JC#G+(.)>6f#6<H4:U/H@QYD.cf(X>3NW>#C]:9X>_/&fS\M02VcQ7dZODC\O
JB>BIWb2LF75A^+g9VP#K(2Z9NTg3K1f=/&>7R6(7_H):V;JI+#,.a:/_:cgILQF
OeORVF0Z-da^6U<TV&JQ7Ed4eaH&WD2YGaK#PP98T98VQV<3];f:O,Wb\eM).(T.
?8/#WD^\IH@O=F]..N>.fY^a#/PQcK0MFe2G&>Q6^J,,Y^7:2,=63W\)#+B/.=V4
PG_\-M=KY,:bSB1PE-BS?+e=^YP92A-[IMeb)-c(+UgLB&2>1D=C23a9aQ9]A@-d
695Q:I-8bWX>cW9,9Z8NJMKK,.3_e=cN4-:RHF3P1G^&#W1T.\R29Z]cCHBYfZPY
WZ0@^?08U5J[fLVO,(MS^<b>.SeT^\/BfA<F@?XV0GD[@GX,UX:WbST3/gaaP#Q]
Y2:>5<PK@-=:GN\,RSI2b)_&N#N/EIN16>OgL><a.(d?3L_)0T&<-50/FSY?NK/I
[EC/\X4C>Pb1B[S]4MOLUFGA8FVSM8\/AM755;NS,-:_6),8Ug8MbCK?B#0KVY8:
-L7^RbEI9T79PR-b4c&K;:2141-Od>SdR8K6f;8]4TOYMag>GJ_<:&OPKeXUU?&Q
T(8&GY7ZfW/Uc_TG,@]R87NQ>9B^PNMQPG-E11H10I[E:.XN>8Na<+75V>H65.9L
DS::6<(G+QU1DY4;QT(==C0;5UIVQFRBVT&,b5<WB?B8MLbOBb)42Y5^aR-?-565
?^/MREB44cA&<^#,_P(PW=b()6R=a6f#RB\^,&+@C2D4G#4N5^++.U_Bc[Hbe\JT
7C];KGaBB\?gVfA<:eB>e3a1B&\P?)W0HA/3B@V^3PS_RN,[;bEV../c]>b0[W_.
f##S1SBZ-b6,:/47EYDHe?PM==VF1]@B&5Yb2LENRLa_<K8aAT&-0890#C\2fXf8
KCBW+TT:(.=BBH&0\X<[<IE\5WVJ#V)FP8:+:0MObeaMb49<=gYI0f)VIe#0]T2A
OC/[PJ)#.aW4NH2HM+-#dF2cb13\:VG;EY=7SfFgF+(9?SG88?HLEH=]0K+1Z.b4
=J[ePd)UH=F3,K]TUABFX^2/:3O#P2Gd03;LBfBA^/e].cJ>Z53KLcO23f49VZ&g
&0?f8;\d,-FM>f5X=&3Af9b6<cg4SZY.MQeX)>U(1BN(d&B33J<2I<PPXC61OH14
+JH&C&3KLU7JB+UTJ<-/W=Q,DJY\Z,OFPOdXK/[]NRX?\c;ePAM93LHB#c8[_g)Q
NMg7P^[DcA,BK>eAAfaR8>ZR=DX=#U(4Ef:&-?g7AY6e25D.<NgTDL/VZW9EF87?
G#-YcVcY5+f4G+[D9F5AJHO@G)#UGSIQ8H6bNb?&U,YVaZAGeFR@&?2YPXV^J49N
8@PfBW([PRW;XbC_8F_a75cYcOI?FU>XKE=fE^44bXF_=(&aa-8\)P_EB8ZIb;\]
5M.#74;Y@=/R15C@HWbGMYN-;&Z<f9Lb5BC84ObH6aFST7[Bca8Y\Z^>@4#MU4_0
NRg<SV_Ke)8>]VbLdLPaEdDNOX@9TWBHUBIKGKM-EOfY19KKL,7Qa&.JCG/A0>aZ
XO1eKY<GGSbN1K5W)]1S[#7Ie_@Y;A;)Y4+;1O&BSPTG)Q^9^4QM@]Ff;@0gdJ=,
LKC;c6.PF8)A]-g+)SET(dFM[OW?Fe5F_K(U>_K22SdJX#9E,4__KD58P;3]g\#>
Y<g^BF<-MF1VDS2LZ8_A</>)>_<S^g2a)Q9-_AMRgS@-^=ZI?Ze<.=HW(+;6/.fE
gXV&J]Z9B96\Tf=V5a4;],8W2g;OTaC<,FDR=eXD1Gb^O]NF@_I,g3IN5bU\1#>#
9>@dW>H<MV1GLGYV1RWS.eJ;MEc656MX2aC]e6Y>]S\[B]3cN1La2ZO/@^/Le,CJ
7He@1UGc?cL&SaO7c<^3?(1TdDca9(@\1&]:&S>K2>R:CWTC4U[-I4:KWD;WK)aK
;R\<AgSdG@9I0fSQ.(gBL7f[b6\f9?2_04/^\L\=UM\O7;BDX.0;^BAKYU^9-(f=
<c#e^([+<V6CcPJVNQf]3e(Xgd5S_N(_4QO0H/Off<1>S(^F2E6g18ATO)^4NbN/
=H/2>WPX,c3VRgJXec/]]>a06NU;a9dMX&OEgeS3E]Q;YDMb)8N@fN,==cA96G-4
:3+eXO2WGS^3755g^V;Ba7U_^V(J,e+@T#b8CJDP.7V4HC(Y>MSN_d1,OT5EI=QU
N451Y=bJ60ffP#A63(TOUIfCN4^\T.8:#g[?UU_VM=1CD,23<J+Vg(JTVZ6?(eYD
]NOKG\26?UXEF/\)<G_Y^dB4cO^SOcBODK,b:f9/eVNSPCJP.V<SKL3Ja;XcONfY
YeW/V#?6S+a@,I/IX#+YI)SUO-<gU<T;XcX?1\=Y1g7&?BPgaZ=CP)G\:98fA@[a
4V/9:0/N(TRg2PB>g;E-Z:5AdTA_,Qa2T3UD-6C-Uaf_+aF/4I?-5Hg/a44IbZdY
1LYF9CI&^\7>RO<cOVS7J1]MG,5DH/UgPEK9;G&_2Se.fOO6A1c09SC@OQBK#Ra#
67&UFN,Sf\J#^(H\b62U8_ZVQQY9SE3,51_L,M4@C<;O-GAUSPKDU;>.[@D@=08_
.8O5AcM1eA7A2[B9d8M75(@Q?,HVY_BSG)R:8L6C([1K[7VSM,]OM=Z_VgG2c].:
JFfSc29>;8,dBC5\dUZe7aS)@ZVRINL7;#N+5f<#gIQ+HEM.1N[YH93[>:^AP0KZ
DW6PZH?EHW2-YFM#e5d)ZT4VgQ05&ZgEb]\@N/[0OW81UdSYQW_32<fX610D/W52
CX;QXEW1+YMMBGR)[8N5]QDYA8@0D\3U37,KF4^+4e?;&M\HMe,1JSHf[dKTJOVY
NYP3QI4Hd;gaW@1D@e?7fGE[2.F59)>F]1--Qb@WM^\BA07:(D&4X#fQ/.d?]4@9
_,FbH4)+05N_e@DAXT:FPRUKf25d]Wa-\:H,12BVQ7HGW-^Va6;4M#VL4GWZ,6Q-
Rd&@HeH>d.VJS#LA#>G^X/R?D4^<g5c+MM)1bMg(3d:41]-S\LK0ZJ@EaA-Bg/)<
88WWVb-&>REa?KV/93B=R;I4PSd_g12/]@a)@^.P2UD:OQX\YS<-Nc17FU35PKN<
\5P(,ML#4bfRJD@R3;TBZe;;fS9]>-RUXUG#TL4Y#R?1LQ#Kb@XKd;Q0d3]([8IY
9#[9;cad4#FQ&RH7f]MB>TVASJZ(UD=g6.4;0@=]T86-Tb[TI@XM1#1&:L)))34J
=BHQ-9?5,LaRFO1BCL_LPEA:>1)V>?bWAS1[9H<YSQT6Ub(E]acX2G,<gZOG?@.d
>5NBWC]R089cCNS,/4S[g9U_dZ>98,0WHc9T<;W<XcW1\JAQJ2?=CB:gB8Id-L1F
YA\@U5GFEM;B^EYd<g2d#_OA-@:12:@-8U;b[79T/^XRHCbJD1T4Ecg<f27\F)#Y
WNXc/&+eG:?HM_,83_U8;+6AgHF@1DV?Qa^C9#01C.N&<g_&MAT#;?&C5<Ve;_L?
6KI:adD?E-#&+MWfYQ)dY=:6F_K&=D+K_68AJ=QNMb/S/_<-W0g7)J]7ZLW+=f5-
bBX1b2LgY=/PLX1++_.U8^?]BE+&Gf,S/f?(YF])/(Bf;7TB=[ZcT,.-H0,?Xd35
dXL.<c]P301DBCI5<=a(-?JM87;+6SPcc\I=):7@aU(QT-5\1IZPO6,TANY..BT/
Yb7JV,b1L\UAUTc2_4,8V+HJe+P@_0518Y@b(3DW/^aG\M#+.Ub842A^FJKfY8fa
<89JDTFF8;d81(<?UJB><Kge#bKgdc]OTUc+DFC+R;Uf-R[F^_Zf9]ZFJFcAYMc,
Ja;HZ+7d34R<bUg1-R89]NYLRgPFM9(O9JgVa2\6ZFQ#fYb^)7O:4[#@IM0M@9/W
c&WUG[[1V+V<Z<W3PH-2>0)aPWR>:NQ&\JgeS5U\EfRS5+M9V>\V@^6:X;UGXKd7
S36c2<05S,:D_eRTEZ=e,&ID?+()JZ7JV>5WL52(Wf<(53R7]N63X@/gVY>cC<QM
YQc[bW9F2Ug[6P7))ANL##D:=+<_0D^RJ]5-M5<Sb;Pe7U#[HF850=55,5334]Fa
KZB;NV#,IK&_52/LM3LYK@EJI\aA3<<,1>--=5KL4^&\DUWa>)M<YX/L]6&]Fe9;
N\Tf(FMOXB<.@U,V/YGQ7d2dQ>R,F9V[5^XGaF5HYF\35IBJ\7;)RM^D?N+>Y9#6
V=R\1b]DA<RCdR5Qb?bR[#=Rc6Z6,FU>7RgeLgH)_C>PA/S^D,L?R,2KJ_4R<#GA
@(\<35d:M@#ATg5OUN^f14:ZMH+&@<4cD()N_bU^QK1RB.58)M/J3I1<I<e5AXW0
>5@#DFLR(f_VM#_HK/3;X#,dMLI\_QX)D/7/RV,e.=9UNN,@=d_51-]@J=f0?5E1
,__,61HTP(L(1W^3T7C_JLY;B73:5)O-Y2RZ:2cUa-SPJBA.)7g(f2_aQ3A9-^04
C_(NX<L9;+dF?VcND-L-QXAG+:CVH&WN[2D9bQF=OdUIDR.F?eLIG(_L7ZAEH_I6
JLJ>VFZ.:LN^e6DY0K:bbWODAH&/72:IcQ(6eTL;P[gOP)8A[g-C)-;2I@aBOfc7
P<fN/J;He_ISAb(b37#,OM49,IfY,_.1(@GHQ/#4aD5>A4E_:C5E?11V:&2.>AR&
e8;&MRG]\R=_6GK/SJRM7N1O.9dE#=F5_:E(fWMH77@bDJVM)5dITI7W&/=,9EE>
WeTI&?Z]-LWVF+b6>>a9?f?Z1AgO-LbUJTa&-e7/5VV./WK]/gVU,LGW4L&Z)?N\
_7ac(2cf;MF[8/e=ORGe^c:g9DCQgVNR5+IY0b9C.VP]YZ2\[HFN&LW#AFQJ=b^]
a[>S3UENKEe7Q5H95cERGC5OOSU8aDec3cc(dLdG4F^(LOG1ZQ3AcPY/+a^X4E^_
Q,W<e+[5BG7W\MK-:G\6\RecO>e\^FG@^TYf5f^_[1AgI0W/F_J?fY>^(&/K(\1X
[QD3Q@aQdWP7dN7#+A>SIG&e^,76AR]f;7YJ.d[0;/S.+5WfZJI3LHB0Qb-0)N/:
FbQQO\3.V9JY##A,)bKb+dCNFFUfBDO.U\^C&:+N_W@)c>@X=[Y+X1E>;?DQ#=-e
4X+0Jc(W&10F.:Q9Y9b8:We<bAU&&Y7?1P2U[AeBdade(0?(=48;ZA))#3/Z;]M=
B>@Q4?d/:<b3&P+Q7^3-<^d:PJOI.V8KTEO35T;&N(.W&61HcT^CN5Y&:^H<5JWM
0@(EDM@T]2cbgE#fX:_#KGQ6@0&H3I/)MTB>B&U;JVOHfENGfNK4L<_.YN-HaEIU
B<;=7R67[1R.HJB1=F+6V00LI@1]()ZU4d2dHY03<Y[R9]c-AA?(A9^62QL;f38G
D-[e(Q4.KR6&?<&W<2<XK3[9W<IL^T_W()#A_4:O><,<UMU5:4OC#?JR-BLD6Z@O
B&8..2^QABH\a<>gFDDLWV9bf#;8_NV#EH??b@aFbS)780aMcJ0Lc<YA[A=)?)<0
?Z1a.2g8g>V\D@#6H=Wb_2(I#1<_/bU>6#b#(@##=DU6&Na9BcfU08Ag55?<997@
?PK3DK9K:M5:dP44V=.Rf=7FEX>96R_<gZc]ZaD=XVM6b_#J<-8503=J:WSU##;I
,:WC+&V)eNL&cdN.4@;R]Cb-Ta\U#N/=bgb=>Q+LT[XZ6\.G4(BEC+eM9L@I9/a<
60A50\;RI?Acd3f4(5#e9I1OM)A<O?HEQJLMM=BUf2ggBB,AM307g]7C61GVAOVc
M.fA)&@?UG@ebV(Qg[76&Eg8PcNI2\45aL<449JHDH_ZHFABO.S5DJDF0eZ9N2&\
(RL:WXC3,0W4)B7dd;gEa8)dBI-@#M-3?dEM\a6Q)^E<b>eGe:=bCIZWG#YdWB(6
SV<80X+3YbUMf#<9Y7./37]Z7Z&-VDdS/EWb6XabdR,K_K0B#YWUAcD&05UPE(@5
>Q.ZDdC]3I.c?PR;5R@:SE4E5M&#ZGAF@f\OV5EaDe[;C78aZ2W70W<?^:-.DZZe
Nd8X?0V^X8eERTf+D:EZd(>V@9S<e64\P(XdJ1ZdMX4HW+b-5?V[9f4cc^N3[g9+
,Y4AYY<(72:/bYCUM#FT3R8/^UASbIY.a:_2JG?)HKGcD#UE,NX>9/NSI57e635.
>Y\<.UVPMDCU(=Q]MXBKg,b2\?8OSOSfU<EOP8QJ/1aU\2X0S9ES^(PCeY1RWFFA
NOC6>\A[_\QIS&a[]VS>^ebLd?c=KD[/cfZ?d=.^a,80=)\MFD^TF@7,/#3A<,]d
b,PG183MB(WNX]0C^GRgI]bX2TZH=CL[&1#Z8F+2TW(g8Z-XP>PBIa>PS5J?HY>L
Y=Y_MV)S5M>BA.^>Xe.G=(Y8VWT<+Haa>,^<9cZL2P@B++18H/6c\18Z[?>7-(a8
]H6,@IaJcQ+9CQF@Xd6K89</Eg&c,>=F>=2Cc5)Z;9&P&BSgD<fcET#<U_Cda@C9
:-,7@5Yb3XE+Qga?]4B?:7D^8/_42>?^B:#Cef5P7a<,NgCP1-IRUS-O[U;DYWJ\
B.((J31aVDW@E)3_-Y5GVadbObf2;B[_>B,\?W9KEMXT[\UOJd[b]:DJU\?9MQZ<
-+-baH0gK.Y.\eA@aK.L_<5G\6SA<49Nd0^UE@1B,8>FFUHY[Y4P6g?C+f0\,4YX
_cG0WbV^?>T@E)2VW?,I9^1-0218^@U)aSACL-4Z@Q2;Rb,+\UgKb\SW7LO=_5HH
=D)VDBE\#:&7c[>SK2K>@I1aWdK;AW7^(@G1DI]2QPO>bPEW9M5E=L#]+Pb(8MPd
(2C+H8d.KB@f17MI0PYY]ZM<A.>^/5=ECZ3NfT=&&,\IPB=:Md)Tb/R&_YHKE=Nb
&QK_dBS.5O8O:T31>#(II+FICV-K.1a5A12M7d(>1dbMa&G1>&-fL1\9OVAW#Z?G
CVS-D1.A2bV&PE7g1KN#g:ZFYcf85R]Z3J(F),A)#WR2g;]O5MP>;B\@H?:^(6ea
-B:aCX\8(+HO&/;XC2A#b6[g@eQZ_^^>RW2MGL?634;H>2X3\4=M;42HF#QOO2L^
VCPFTSOJ?,&/P];bWW_4]f8/9[GWG[;DAQ7bUZb&,[)(.WFWCT5J>RH&?,_O;.HB
^Q.F9K6b[E7V27<_D,[ea)&))BPdCOS+&4F7JCMPTQTC[DW;R#026V+&1Gge36F,
2&?@8M?8Ce_>CW\1(G;KHKK-\J,LUS3@^2B&D=>/H8N>a5Z/LH]f0cIeK8]W9d]F
W^PY?J^#X0.D[dXRLf5;U177983LVEF+f_Q9YaJJCO4EMPV_EUeQ17W2<BZAY]b&
X:E5ab8;\1J1K2?HBYQcG.9.^a-DB1#>H^]W<PYg.1,Rg8P,Md5fJ)DU9[5KeR,A
2U42dMW-1Nf36b37aAcN;\&7Ge<9NFT\c=DBJYG3IU#/71WG1G&JG9XPVYgGDgER
c:&AXDID[V^^48a2QJ8&6<a4W+Q#;;UF@?2D2NY7b&-^AM4E3(=#AW0.9&71(H3I
J@&.>T?f-;T-KSNMaOZZJ:63bLVYB^H<LU(T[:]/A</;,D9^Sc[4NL_F@HBEYTNC
J(CM.E]2])e.R(9CBMaS^>1XL[_KBFI(H].,V&])eH)UgWQU2IC#LDB_PG(_[4B[
:)LO2(5?3JF9F<8BB6]A;@e5_C5,dN?3?+cIg.^?+?e4^6-3bY,b<Z.9EGa<NT-Y
1MSS:2H7:<=O@1V:Y_;RJYbI)e^8fQRW<[8AZ#SFJ^f.&?(ZWKYMLDBM+SIEe[U7
Rg[\2S7B58S=)+ff;.SgZWL(Z7/_Md9.05]3B\Y^FAT3VPg7UDb2LF8ePHd)A<dT
@3c^VRJR=4B=;)AZ&JY,]DXEY^g((6QQ?U;fdXaMQbUgEBBRPD;3<4X9eF;YdMW>
Z:C?R;.3QK,+R.a?4DI107-&>E.7.;e8R=3>T+69G5-eE;F<[DYaD:B7S-ZPPUKN
FcHRL/C^S6DC,5?=/aN>]F.Z[;/3fWFL+.(?7a66G)3DXT\EHf956CAWY_?De,-2
^F)(><LdTZPfL@PP6[ODM:a@/97VQ)8d;DeWa,\M]d4[7X#)G:GARWdAdN-B1e1?
#R\M6G1c#7P7eNg]fFgC.2UW(A)Y.SA@36CeVW;J?bPScY5Y03GO/f[VX2^2OOOR
:IY22[.[.\7V<</7?F@)aFQ#]]HWG4#VM#g0]2-4I69Q.Y+4EScF>Kd1N\@Q+DC,
UCEEE@?BXRY)++VPR.UR(N5?Q/7XP.HS,@@MMe8D>VG#84&V1YVDBbHfF#S4?&]]
_2I(B->S-9X@]3&1&74,(#V>a-bUbgGE]JOSERd2R\f-F+<dAX8bX#>d6:FV??UA
[&=ZU.AH#8dgF5FK=9I#K6=:RA7](-,McNYL6R;N2:FG+3:WF=gO3gB4.C4M(,Hd
:ILNg9&66P4afId<c=6aTaD(]G:&L5X^1(3WV[3AYfB6+S2ZPYc_.7_(#>LgM2)U
A9WL@8ER2)MfS12A<W&QNIgS,0<)RSX&HM>R]f8afLTL_9;1^IUeU26A:=TaK\&D
/g>KbH5=W>4.FMU3^UPR0N2T\AU,=X#Qf0[;1W8\O0H[.2M8UNJBW4D,J[b&9ZDD
.E:X6RIW(Ld:M:R9PO/b9M:;]H>FQFfdbW)&1ccc;Q1f_.M+?)/GU:eDf&RN1G?V
&[+3E#-;.fU7bLgLR3<^7SJAb(&-bI+0;(c^PIO-O#&[g9_]<UGKN&M5)[Y+NM>C
#;dXWJNZ#W3GY28]6-3=;#(.5S\9,X3FX9S&\+ZY6:K#7C]N#G:]FR[S4JU_V>6)
/Tf6g,NZb]]?8[M(1412#WVeBFS<cf8fP0SJOPgbG93?>5dBM#[-M>#2dC2==.>;
Ng>VaV<dbA_YWcT91?(O4E9N=[7\,d=Wb,TI9NWY@E+WZA2XRXLI=d4TS2cQ0TJ,
R/TU#.=9()QFMH\O6JgN8Q\#T\D\A71[8:DPWLE(7LQdUc]I4Y[3;MfLGXea#cL/
+=fE/I.g59fHA^7MDW8cgP]VQ;d,8b/OfXGZX?V6?f_K]OW,VB[7,:^BSS(6MA+)
bWP4U&2#+S\:6)&61b:^UN5?C^RZQKW/5>d8+#6;_gO;?]^67bSUT;ARCYd=PR&f
_MV)C9FC[G.8/2<a]b/JRGZ)eW(X)37Eb71E-</XcbKI=HSO[ODA;DZ6:[GBS.Md
<#FEN1LR3=]J>SYLJ7>4#@:-NCKS5aF9[KU?;:=b=3,]\4AS]8H?G+JGS/F+)PbP
RP_QT7J.::gOZ0:F;c\=]#49G^Ub3D7Eb7;I^<+gNb+Q[58a#5SSM=\cT.7g=:c.
eLX1Q_dCU3@,?\:cGXYIB(Ge+^I5<EO@FK=F?OQC2-.8g&4(2TW/e]@H@2\g8E7U
K)A3#KFIVFGa,.bPU0\SPK&=aQ7bMQPUd\AUZ7Ac/XGND#2Y=)5@(ZKD:VA:f:T?
9:Z8;NUV#cT460];1;OI(0;Xc+JYZ#RL7Q)I8Y&S&U;0ICVf5Xa(N7,P?.&=O=5S
:.@b6bVIYQSC__8BY9-BB1;e:35E\1RXFD5WUd(#A2WE\BQc+OF3YQE7.=J@>^He
PcB+6AU.K5?@F7#YHgDM81RXFA#SB+O/)R:2W9fXfQX_Dg]4bBSL_&J#D-bR?Y_P
)OFa^IDT1VQY[>#+PQ.+FG=:/Qgd)4KK]F@SN_VC69YCWcUaM9De]fC4+ZY_Yca\
NZ@H@b8V>6/?6f52^3?@Q3=Mf@cP@;UD^Z0^7T4bK@OKVEDI&=4])CD.=RZSZ,TR
/fXJ<J>YPI4)@a@^Y<3YK_b>I/+cEAJVT2dSf[ZS+Z[);+,e9&?]]K6IM9F<2Ce&
_P-Rg&Q++^Y-@55&OJPG=OTJ/W>;1AM6#II5b+QcF1)+X^UNHe06&g=8_(]Q9]XC
J&-89+?#e86PB;7G:cDJAdXD[,=CKC\KYX)c^0NGW]<E=TY>I3ZVS&g-;#aYgWA1
+TcKaWOH)-ScG>cO;Z@97H=bAUTc9A6,=6;<&;2Ff.DBb3O8)c=N^)cTd/O?Z[Y[
=KZ/+@LNGXc59[TbfZcRWZ]6)S3V&[4O&_=GJCU_/3K3fD7-_]V<D6@LAFJ;TW&(
gASICgC<09\H#Sd:c4?AYBTV<(_OX7=gJUVW?@5X6]G91/V2\B,.7-J791D\,B)_
6O;-d_6UXg&9#0/L:HLEUM_b12F,c3NUFU4J,GLC5O^DM+/g12-bNG6Rf3T3Ye[=
5#[P958Mf/,d?BE2X51Zd(U-61GRG=NL&][K+;a(T9J4gP5SLA0b0\]38YI_R)Q<
cX^2D]@EAWYb,T]A51FLDc^d<R^aQVV]4d^d\[>XcPf+bP,-U:ff\A]2V6Y5NLa(
+C<3J]YR2:10UW[>#S;TNT-:BM=P[2IWNUT0J>JNHY[bIH9Z^T&I=(?24ae785E;
+[T^[@3ggMEfFT1KWWL2ZgS,\Y<4eHH;=d610E=:VF\E+4;f4HW7.9UM=P4&7<J-
fTQR+4?4]L_[<aJ/W0g.[]bO[K])bMYC_aU3_dgdE03-Kf;,1+&8Z@SJfXCcK05K
5b=J-<0Hb]<Gg,?,1MC?/JJF3S@1,dDRf=4=)2dE4_gcdc(]GQH_PU)@[#&BFC_H
-TH;X7IRSe+J/RabO6+_H:8#/>15IL7SPe603eI/f0cA=ZQNVO9NC3IH0H5>Ea0e
S_?3]Uf?Z-aJ:3(:-MS0\&WaMTY1J-51=Y;]=ZcK-9CXaAMHgK1VTM^[(dc=R#1&
JCMb<cEGbN??\LD32+7]YCe2\)8)aeKH]?eQ6,FH7X()HA[]BgLX,9P>2PJZJ)-]
J&;Y&5;RGH#0L2gf<?M]/S]DQL5]#J.W;,dH.KO&\YPfaD48U,\S<#e310,?64=W
Z^=M.8FG0Vc(V]NT1^H4/g&N(D+U5I2#f<@,53R#;L6,3(55KA<aO6H=Q5e4VXQ9
RcN&HD<N/,2V]KRH8GdV[D=B@\(1C)3N7Le9?28SfLZcO(<_OaIC;<GEK0c]cXBc
fe\5O>g&d;fD;@+QeNTLS^VY/X48CP.6:W=a]_K2_AW_:X4I^]+Q87c;gD7A+CO2
?ag>V12=+NGJ36Y/RK)[I@(_^G9C,cC1Jf2EOGXeaEEZ=;[)I&0Ye@JLU9&/##2M
PWB3H,E/b)3TBZ9GK32/2J5]4ecH3=d8[60/\c:Ob)Dc:^)-TOa.&LC]YJ\03_YI
8F>.6=HD#K=,b@59<7J5R:P,+7X0@I]UGb+MLUAAW;M8@I_/NDd^7,^FgdX9XJJ4
BX]c0fcd3O3T:1?>4:1CZReQ1JM2FD0DMHJA&Ka?/0.1:BNQJ.(S3^_+DD56Mb<V
L_:CEgaV,@7H-?PUAW3E,50R9?QUb6O02DDgH@(4;S(c6I?+ZDT@K(c=TSY829:)
5WA+8J>#XV[R19F>ZO6:bD+\2C6PFU2.f&Gb6>HO]7bWb2c+#fgg,_dBC#-W)1SV
fR=]@0f@35Y:,>bgA>P1;X7X#P:gJGQa/d[K(5AMcG#Hg=?_,5QPSAZJ(87d[d8X
ad,E:_^W+(VSRA-c;?8M>-1QMLXRHdWU)QI&AfbgC[/W26Be)]EGVbXF#OQ2S8AN
;RO,2V\T2.VQ_4JT+-JTa.L_-D<J6YTUZbM#\27HW6@[fYBg(AU-J)Oa\BOgC:F8
\A?.8-Cd&S16+d,D,-KNgD?4:aV]N]QS>=bUb57I?_BP#Se:16aCMBMT((^1?:>6
AdG)JLQTOW@?9NM/\6TgE93eKE/_0TU?@?HK)<dMBGXX0+&,H0\V=WY<A6#B5Dd0
FdVI-\fB?<\Q^LWBeXKRb#aU6>PeNH_Ae?8Z6[-+:.RZYVTN/2>#^e6+V91N_6bJ
;5Hg,0GcG:fA(c@CC]5>?&A8OWG6?9?Sg_(?Q.bD3SK=QNMIGA0=J&IC.EI#&DA.
-?YgV=JA.d>c6&:61^U>H^(]T?(RY;R>30-A7^7SUZBf=EKNJCV9?2.<#T]=62.,
f]Se/cJU)W8UKCe#;]PU-4c/SfcFND6(Cb,MV:2d6],4b#/-O.M@7Z:C:2:eQ22R
c.4<AX(8fHB^)Qg_\RSW:(7(aS0f3&=W#Q&0^-.f])J)735cQW82E;#VRQdLfC39
&g^cP7UU4^(@G8^,@(G_X9T4MU2>-c)K2aNQ+LI\->MLTOZ-+QPSBHgddMNW:_fV
a)\_<afIg6,S0C:DU\1]aX&1L0De)KP=&SA6\H/=;-PAJV?EZ[<dZ76LGX5Y58+;
dZ\:f#;7fQF\,,bLN985?&X9,@_YXQUL[Q/P^=>ISX9.I5W;.>FVQT.OW)8=_EDP
+&47-XWdDfJa3cgf4ZP9/3Y+V(Ff5]GTY@RN>_<OMd+V8:=:BMW>Q>]bA^MaNcHY
#.^.(?:0+,.M@[0?fgE,TaB(4&T5R\7KDP@-W1:+8D7H:7..Y0eSS;ZAIY>OKSB,
+^<R2>YVUf+2O_[g_LVbGWK[J@=L8;ZbP^/\M9[3-9QR[[CSN\8<-[I?B[ZfT;b:
1\JLC50/V5Q2?3@Z]Ndb)[PN3+DQIOIX<.UEAMHD6AA//=aYO<>Bg9;07+0-=D-M
=J)X[e:F]4c_Sd4T6R,gEdZ.]22/cE>_7a0&Ad_<+G/>UHQ4)32OKF56a/12KN-R
d6P-23P:^V2,.=3.^QE?N1=f6PUHT;AK/?@R@TNb>HMVUFI4C5M?)5fQV^HR#[OT
g/PA>^?K4aX^8Eb=]::cUNXI\K,U)MOT^/4DSL]D1L83gX/L+Zf(_&?c/VSa\G\J
c6UR@WMTQ+:QCgAbZUI>_a=8^7FZKW.8QOENa&McZTJKa^^aGg\BgQ@),02;_#(J
0[_CEOg2ES#^Z/KZ?KeX2^HZ22YNAA/_ET_X\aU4\\CDd&PX;,9HA]ZC;5V5>a1P
J<FVUQ)F1?A>UMUGMbS+T[A95T(Y?0DfPg;YA,4FZ6D?GRc=2JHG4B)C1Q&FB^6N
U;HA.96.c<I[CGdU3QCL.=^-)WI;aBWH_HXQB5DGc3d_Xb9Af39:)F^OA.-]P0/-
6D9I_cZPK9SdH&bC9.bMGR>fR0?SHPZ+H1K8<=2aF/T&dQeb?H1S#bQDF;0c31cM
GS92R7#9?B?_UQ.]KJe;(g<KaT9<BH2C[4GJPKZ:_J(Gb@TSf_bT:H]S_;F.2Z_8
gY1dK=[?c5N@S?Oe=G^E^E[9]&3ZH>1LY5TP9F.U^(U53G3;RZ06N)eZ^EYZ^)8-
cC@Z7=:F<9dK9F]P<IQgaT.+GN??>OY77g<CC(.;,gZ,O[)SfR8AN@V?LGQ<EDKb
T-)2(KH,E#EBQ5L2#W/P9.ZQFW[[8+G6acW>[ZSGbTG&\#T\7U)J/e=FYPWI,45X
FNa(:)MOO(?RERMgBJ3Ib_DI;N)J5:f4=/_DL3HR:C7T;^D&E^H5+B0A<L_1H)g;
G,793;gbNHaBb_@AR6CA4[S?_XLAb8.Ke4J:eVE=^S:d#;ERW9:#E-?PA;]6A?D]
&7X?,?ISJ)TN]P8FGDDK0NIYREN.M;5DS>75Q7Y<C1;[@-=UL8&Y#(2aJ6HDUWYd
QS3^M.;-/IW/TC^P<A1X>SAgH6-a;<DXO[VGNMd\IEabJ?8Q&)AD&K(UM2O@ED#F
#/W=.K+BTO<fcddUb)@;_-IW^JLK>@Tc_E.Oa0MWVVT#=3ZK)Y1773YQ];^.PU>^
&gC^[(6Y\.ERQGBDFXOS.#NMN38+0S9,=B/e>O@aINb_3UdYdL\Jd<IJC0c3=RV5
086V_T^R1&Tb?MZcHFF4O46T47IWFbbBC86O^Le?F.7#H+^U329>EQLS0K/_M8UN
M9XNQZ@./L)L^)Ga+_D1a#CSFaW-fTgcN2Ic#f9)=RVY.,J+EH_5-;0+RfgbGbB:
>/SGY-#g6L_<f\5&b\c)C:=TXfN7.,=E#[)(67X8,SUL3:-\Z9)cAf0(S<;5:R48
GgR<TP33:+]W=3f;,EARCW//?PV>>YA5+3c08.Oa[V)9XA=IA)2YZb:gN_GgP8JB
Q^+b4G)1@&fYZ^.693][J+=S7cLY,gK^NM<&Y[g=gX<D@bA8>6CE^FV,KM8;7bH-
.6@CGg,50Fg;>/2VILSPB:#0VI@d>>]Ka)U/XT@f_a;@0YM#83b<0EE/,MPUOQ,R
?@L9LWPSTTU&cK7T[8O\_MLTSQB=g[&)ZOP?I8_g;V&F+U)&PWO21E.GOLF.7Edf
L;JP^V\M@UV61d?.?J\68g^)Q2M0<#A(265<-^GBU(L6C?3NL.-O?/))fNN?d)6/
dP;;;^dO\RZg++,\D@OEg3gK&(<X<K#2fD(N:5-]UI/PX;XEYV+:T#:TX;]6F(fT
V1E9T8e5JO.e<HGf1S0.ZA7]74U,7]::<SH+a4@.dT)aJbJ.<G2^L5DE<c@P>^a8
+OZ//=aDT0RADB/6,8F)bMC.Ga=,MeKIDaU(6QKQ5+D[Cff^[+[BG<8<g&T(A:O]
K_O/<#PC\3VE\KO6OcFB#Bg)RZ)fZdRUGEQJG390<,U&:R0J3PG_2NO)\A^32fBU
E&;S2X_VW2O8_F\-P0a&3;0A(Ncc5P\=:=I-[<eU4Fge6?#TYV,Ug?B)ScX6=H?P
_bB0(NYIE^>&4)BV+TVW9BB3c[aJfTNLPV423J>3EQ?M_.18K@6-H_NcY,3@R@f5
H[\NBZM?dXW:K51N=^&-e/RYBB:L?=I.c1.EO=VPb9Rc[B)0YUTQW(N#1C9Q<EMf
^C?FA<dPOHb@)LM.H[=abML<RgeC=F@NV0+),:aXF,B[PYLA/TdbN(/4.CR06=;(
KNA?F1=(\cQ740^?9+\,0\[_5&KXE-JHV=eB7<9[:-(R8<;gOd.=07QZSffYQF_Z
UZD<P4#<71WW\24^Q3TY?8a,M/,JKJc7W[1>aZ]Gb]^+Mb<,e;)&UBBd(aEgGMMG
)46b-T[X6H)W>G(;_Eae_4/=WAD8f:c87V5]EX_Rf&^,XPQG]NYX&D>H7(UU_0G&
^fd/4V9_W+VH.T,SO[@V/9;NFN6#/c:ZTU9N>/-PARBcS5L/)JW@b:2\b-:E2bd?
MB#@<HSC,_:,W5.]O\dZRe0_5.5M@Gc:Rc=:+CTa_K],L_RZKENJQ(L=&U\O.M?/
+5N7[0HO<4;@0=4A0>-3AdL^#L[[PgdP=93Mc^4UbIZ0NYB,GO-JIDRO<B)/C?;E
2PI&2I@.#+bF8c==2^9f^J\XaHC6A40JQEc)99dOIL<UO<-/?\_bd_fT1^_3QKA(
3J4=4Y8+RH+UdZI7>CN1E>c;\-VX>WFIEgJTQN6(SdN5fH1BbGSaF#],GWa?_8\c
^._#(Z8aV;X,([_)73>AILbCGVab7-7Xf3^<1-N;fJCH[P8R^YU_B3;+ObJ_dU8R
(W1:IR6&Z-I2S4LR1R6S9G8.#OJ0OI++&ba);6OU0F]9G@FCN(7IT;Ed3=R0(c1W
HLF.ENG+Gd6+:]D4JU1[&[X]X)TCD]KdccLR\e6&5:MWRB[QSZG??81FC5(\_;K]
5I2BHb1)ZSCXP2Ja)\>5PG3:a.[8]_]g@T.PVG^4@31=/dULC908NFL#Qe&(\6A(
7.c6A.4&7.F:7-I^bK#=X93OeLd^IIQc[)>#fL+P#fa6fQ9+IJDK\+?<C:=CaT&+
L>)Zb4Kc\488XaI]BJ2OaGK)Ye7MDWC&BIV?5)<\P63AM/1U/YSHI2-)e(dM=62P
N]e?5<?05]TKM]6,?fQ;R[a;/MDNdKF?]?eUB6M5O^PGF8E?0HF<,BVQH6]gLaGF
@?@W8:ECG7VXZ-[75[,a#FS)<X_==ZVI?:+<\)C6?4:ZNfQPQ>JL=;2<,BGJ/d12
fO1;BP[[e4U#QG+b:/;_5CLc9(=+U+/7>)42I98[E6,C\GPaMK]UQ\TKY/94/d3:
a:f(L0_Q?F&#a4MU7fgG4)P/b2DFA59T\aNX<P3b&[H:N/38:eACIH;RQgNRC/C;
;Wgg<>ZL:FNBdPb(^1W;J.2D=:CDdJUTNPND>@UT<U>-#2bXEE_VB,510+TK=4,Z
QCFX,>W6BbeQaH8:1f97JS\#dS2#e5\LIIA:7dBOXbHDG7R8Be2Ae<=_[QI-8.57
YU8H27FP3D<AgUA##+1JHVZC.+5&aN,IU.d+PaX^T_2Xb78-#OM4H[^a&bYUc8-b
QdXcWC+GA6^SMIS<2]EV#;AA<AQ^Q7dPEPXdU05aK66NVJ;]HL#PYRYK:V.e639b
IAGT&[Ad(f]YKMZ-QIPUUNRG(Kd^B-#gRd3NL5c#<[.>#][V0R=WVZPS9-F7daRC
PdAMJ8I^=22\,Ka:c^]0/RNSgM9M53S<3Y/V?A^C>S2V7:RYF?Y3VS.X?=?M>OZ>
V@:D1G8=L+)93)F.@)^e[T,K83-&R)@^A,0Y6cdEBf:^+^NV5;Y-EI.Y2LgDK;]<
?KYFgPJ992?[62+)Y#eFQ=99.d8c3dW,3\L>c3.\USdRZA\2#W)RWZa]I/5A:/13
4@.;W.UY?]-XR[W/P[I3e8M2O./H[?Y^;+.7J/9;4VHL8c#+Jd/0fgH9+#aZ@M@R
cN=PbgN@Q&0aE=R?9e&,3R2:LD]D)V//=Z,Da&A<CUS>X#>RIad>FF13OUK:H.7X
W]MOG-QHFF^,G&QO38^AOGGC3g.IZ9[B[I+H&PW<Cfd^D>[M(YT<_PYHT,ZQKIK_
EfS5A551;YYW:b)M,O^)=.R#aTEOL<:+g94;V3bM:[EDANZEH]9,EL(5H]&c);;e
ag/^ZLH:3d8?4+T1Qc&[:c_NN+T\Nc3[T\g2LLO,C5-/OGPY;dJP>,0/X-)7UA88
WO99#W<@=)JXD<MI8)H0J4;<Ab#5JZ09S>5G9f5Qb#-=[f_A/]<??BKSV\Fb5PH7
O9bcJ6=JbbR;ND)fXX]>;JVPM-KJXg;GCg@C;5>#M]eE+^#2.#3&afJd5TGI6bH5
DS1dbfP,>@DSYX)0KJCD=RW5WFP6[SCM#=]SPff<&.BMY_VH<F8AQ?FB=K7=9UF?
U9E33\FYeRd9I9HS6#M\)KLF330EA3/SGgB>,P_BAecQC4]M]YSK+V</UNZTSEe)
R_+6@#:4>?_KJ3eE06D&,0.IGL6d3A?63Lf_L,^B@0GB6PFE]0YT9bZU[<-3^EQO
-I3PaER0,<c13a,[c5e]EdT[BL[DZQEQW>[4DALZU[AR5&=>Xd5=HWfA4[E4TWN+
;\bE1KQ<T>?Y\VR:bN=O^-55gUd>MM5_PDGOCY-\T(=GG5;?@SM7@&-)G)b/T?3.
e>>E;,35\J;dO;=0A]=CRDH@?0?#C)F>/\V&F<#G:_<D3dZR2]@5LGF<_H@0W75e
:J@@@OQYD+IDI^CUVcG(-cYYKB:d?HU7?#R.dGD>>-g1<Z.9E>>AaDOO61b8&WUK
NW7:R)Q0U2c+QG;XRMcGSG2OH,Q?P4,RbNM5_SVI8RB1^?Sgg&6+NLe:G#)K@6M6
Qd+SXB,_efS7X:280?L5(3e892.F<&[XgF1\2>KYc\a>+dQMGZ,gW[2VKMOfSG+\
[>.bPR]FPI8:aT+fK@W[ea9]67?4gT)_X38UBLfYQ[MZaeN8af,6bXHg7LRe)3?X
FS#P9F5IRZ(+:dJXFd]]3\QTV,,^2+D,HKE=da]ITED^JdX+/<gZ<1FOXFF6SCe5
b<F6;H+cbgLRUPP)VS;<)bMcBbec76XJ&]I2LZ0JFAa@9]b9#F1VWO60?UDNHbXP
&6YJ:95]JLQ5AOEC^K]>a0Z>eCQd22&1/4?G-UdSc#:.Q[;8CEdS0K,SMfOEc.+<
@6/DNAHH&J5/-<IH0BPE1]H+KH/b_&[DM&b[0)ALR#T#N+FT3V-4#6W3TQ#R3?8V
^JXPTK:0)1/&)H)RdJWJI0d]/;W5;<9FR6RJI/-5P,B^=8\^6F]<H,C<:DD?I,>#
DI\fVcAJ5_SE#:O13(L5fGBN7c<J@74U(6OX.ZN&@7cUPQU#?T_MK0C0(I+4Z#HD
IY11W4-Za9(RQ&GL>-C;OMe.R[T4Fb9#B82@0Od+;,VL/g_g@8S.BLPAXP[P-O_d
A.9/&HOP]HPQ?A3_c+.d1<9g6Q_]Gf#((fdb@+Ff(cX2MY>IJ),TZ59c(ARZ5Mg;
/GDBdTb4?XK.?>5ITe:?e9(#VTRe]+O-bT;@],Y)ABUDXRN/0U;:8O3TK@U^1+<J
f44-f)56EdLfdQT/T:IIE0(#4$
`endprotected
              
`protected
QV[gbBQg(A-g(\<Y:NKB[12c\5cb\VU37CG=CYO&beXdHEUUV+bR.)BBXAgdY[0-
&>ZLaJQ/_C_KP+E<>:3=K12c2$
`endprotected

//vcs_vip_protect
`protected
e#=72P9-.>?4.27[=45?ZHCf;B.LbGWeca1d.]e,;bQe-1_6dH:/7(91JNE=\ddW
D>ULUMfOXJ[d)-YAHbO=K=.FCLPS]I/3YD4aNMMI2C\^\9U+HfI@46]b+R+FM>U.
LH0b,V87a3S]IDHc-d/?U(5Uc@-][;1<55O@C;</&OBGCZE&2YKHL7Ef8DAcO^d\
/E6d99-/880+JHR201DVU0<V9_L-P,G5B?Q#<XB;C3/ZcOSJ)gF8=W1DL0A_SF][
D;8^-\Cdb<>fFaVC#Y[>[5NJR0cV]2;4#N=2dE/EE6SA-HMUR\]Z3L&CE?RFgcZI
@eZcU?GcT7e)R+TXeV88?.>PL4P-U1+,=@#802K3W(O7gfCHQf3ZDE#<EL+XLDE]
\#DO7,-c^Q,;G_V>-VQ^,@U)I\F<F8/M7T#.>+RfSE;^EO>KQ+#1O;S@)(H<OdCP
OIKEcTFB+BI125UV)+A&fJ\cHPSW;TB7)Sa6-I>dXc&9bC^e:;e\SQP=4e_&TN/5
/,A93DYQ5\55WQ?XBAdV1LBf1Fd)ZN4^#HMSR]1eQ3c5,g+/:E<XXcE-Vf8,Y>0a
<XO;9g3PE>=Z4I97V3F.XQ^.da25aEAb42dWYNG]^/g^>]NNfWD[B0>TGO8[PT&Z
+?JEdcdKOJ2U3I9XNN?[6J9&&]W-W(V&g;--W_2;bZ8?8ZfMAMEE.S-Uc8#/TQ8_
QZ7BN?;7fJ8M.?ADI4^PUG6_/db)UNS@8XWc<9>F[fcE@^61F=<d5:eE(:S+ZgRS
/;Ube#22F++:O726Wa>/]]WCd3ZYKJMZL)V:SN6YObN\P&NBB<ed<N;R?E>+GK7_
2V)@I[Y<M5JAO)fH9SJf?D4O6G.1;?E/:-A:WIQ#.:,:E]I48+HKAf9I:N^GJc6Q
X]T3\Y,7TbN\(F9TA]gMO=\TA_&Rbg,ZJ9MK<VP.\6gXU91gS0(NT()LITS+TNQX
:\X@Z8INL940L0/=-L0N&^X56\ZM2D2C;:Z2gA,e#6CQ<63H-Ce<TDE8bW=U^&<6
<[?2,I,WT[W?V42-cP/1USAcfF(\<,g\\O<=UDOS];A_WXEQ<);8=-V-U><<(R@P
<+N3eX@E0@@+_H[g0H+Naa8RFT77BDbfU/0Y-Hc5Gc,<U60PcD6#V,0YMaUH8e\[
^R]G-b_;>8cS_40\](/EBJ=M7L6192O&L6XA1=X]W(2W:2(T#J9>J4)^-<?Odg:>
1F7=4HVE..KN[1V>4/+7/#Id86M_8[XZ_((.(H76IV@KE5AJW6F@;.HO1EXG]?F;
I45#:H[18P6)8.AH4#4P9&W:)b<a5C>TZVP4eHIJ:5O)?E+36P068;b7e/G/bF>S
MZPROWUW\aN4GHP,b^DUH[^gT=>e9_cJTYDJ,OW80-QJZFMa_T@>3gX.NcVb))QO
U4\_DF2,-AB2A]1Jf+7#a9VY/d56(DP^)=/3BSBKN7g^PLDUT1GB^D9(Y?0A2G3U
M&2b8^1@1./=U>\>2&GQgM@)GcaNIA<3),/I1T/NJH6(G=J+863ANP7S(VNf;AU.
H8SN:6C&gX<fB#7^G.>TX1a_>)I_H-C44@?1NQ@4O52<c?VTN8KQd/:A?W4QMG?C
C/00QPI+FF+B1/J4d-FP;WfA^^,=@Y[GTd+CX4#G4.b9:E\18;-Y)gY8:_.QHIX0
RB57F(VE<FT+]OLdFLU:X_e,?c7-;(RY&,_;6&S:E(+55[DS>:7^8CIKcP:/READ
Z4CS2APG-ODRX8:<LCDTdNLE+4>=[4M;SPMPNOK].Z9AE?H^^^VN-K8aBR_R6dcW
fJ@C3AW@^BNXgge\XT:##g[HPH<@:UBMMQ^R5I&/;9f^^Kd,?G?Z)XE8BVW&aU5?
;T4U=I@cA<9gfLU^fH#GI^AKHQXE^)S;=?fg8dN6CO<G521]bF)-a48d6bYb\;J,
=-V7(JZOc>M\JX6K_LO_Oc\^/5HQ\efYT@\Y7[/5)-/cYG.S2?5RBS&MSOM=;(aH
;8AMB<Wb7W>GY@6RTMbA?H=H9^eJ<<be^R9KAQ<PTg9T1B1aU(RXOLJ<aN;LV-R1
5>&Dd=c7FPJ;O<e5>N)Q&PTF,0[>N^=)M.+?aSC;/0S2)aN+(6C3Z.XEB566]<K6
a].6(b/T6IBLPQXE4Y5W9/0bQ,d;&f.X&K7;ABg.\I5_PM_L14Ye,1)GIU<XANdE
b);C84gc#+<2:-@ERY+XR7YGa9c9<C)XK<M/VO;+67Dg(D3.#-5M+eMMXH,PJ_g]
?e=a/UX7;A(8IJ\8S(HGaF99a>@E0YcT.]H?aI+6?Ag=Q0JMA8c6:d-XC+92J@gG
egCWXNW1e:DVaAC]7^#.#X:(^(H?a+-]0I?b=5,OF\V.:dS8Q6PT4fMK.76f,MfK
@;2=?KOJ98^7>DE1)6c)._V4:^IOgTXRP.[3\RE]^ABR?O;6GA/e\P2QAEMEe@9+
^Dc1<M/Ced)8MD7)BRUR,&d90MYc,5M^g<9F.ae1F)F#+5O635X97/;?[.:UgGgT
aMEMHRM_:\(&XPVTKRc]eFII+67;RX-S-&W=LCBI7XG4e+(=d_M:,KP;+I6>RIJY
PJ;?96Y\)FQ>0^\5K0VQ&(YB89?&J72?BIO#JN]R[N4TQYPH>2aN/7AR0NJC9GaM
@de<fSg&S/46<PPbYNQ[Bc9d19)>+&@#eVH4P8TNa=V:G(c@E9)Z?E-WS)XJI;?+
RdBP[G#A<,(\JN_eZXJ-/5?71@96Z>DaMNL61#0_e8@H&JJ@NdOfG7WHGGd)FH/f
V;L.&b2;&X_JdY#:D6F6T(E;<RJ1@Vg4LJ\H+^Kg)U:e:I,/X41A70VY6PII?4VD
.6QGR_UP9);<YUBJ^OJY<(3Z(1:3>,2R0a\&.PR:7-DW9C1+eYRWS?W=?JU?4@WO
DCABHM-V&06MBdU,5ZKXaVNbSLVR.]78SQ]82Qg8?@/)AU\>G4b+E#([OE#_P)eK
C(Y51Y?T<F92RK]C[4\JNb7HbcW-Oc&A4,3[44^A_X#eTK]=22afD[]M85C;f6.a
_?K^?=#22cJG[(7b7#^_5(1N7gE<NaG/L+.BRQQ4TK]JEV54Pa<Wb8_T@cTA,aE3
2deYY1Ec/Ng/\XC^Z2NT+=69Y6VH;@DGND5I-7H,Jc:3N2ITY6&^R29;XT0deg2_
5Td3QSK2L<d\W@G;]C<(M^cS7Z:L.0Z)ST_:98-HPROUH3>:+VU>bDXS&GL61dUU
OFWS0#BG;K&DL+f6.Y-TDa\3K8L.,\V#^K03)Z?4\UMAfVJRZ-fR^&P];POH&#\;
=RI@:9,.5I71RKJ6BT#1gAJ.JbR-)3<gSZ:VOa4deJ\>?:[_E.<RE_C;T)NB(WC\
9>FM\_5d&->0+Y\6KagUL]U>cgg<MW_LNWHG8B]CWXA/WI-)J_02U1I6gERSW_XY
;98W4+#SUOL?/DS<[D6afd>G3L<g?[0E5^DfX_:a,Bg58AK1D)Ze65Ie3RCY?Y\:
PLZ5+9Mca9]a,7J1]H\/3@HHZ\c@@bV#];?WM]([W&10BJdVgJe9#2BQN@ULF6#)
L6ZdeOXZNDYWE^\4GOTMQRX\GfSDTKaS)[+cY)B[5gP(MGPI.g^F@R7@9K_c0?,)
V2V(DX3QYa1+eKS[6F&g2MX+PTAd_5<-]QADg3Y;bE<XM]QS(>gcBf>+:J]HJ8E7
Q.I=?5;P>10Z_USMc86=59R9fK5QgEec#^NDZ2]cN&NO/KZ3H0CQ-<4BAe(HQQ?g
I_\V_>23:CDS70-CLQPQ9<a>8Sd./;,fgd,>QT6W/]BFUd>Z@WDB3R,0(;1)gYf7
;#W2M#SPNX[KIM0L8_g>bJJ1P^cBe\8J=EA/.Fd3LM9(aH\@+:V,\YPH.A^=R7J2
#M5U4b[IS,90RMEVTAg2Nd/)4ZC4PXU?cffIRd9;S9=ccBXR>[SP@Q1?L(L-b8JS
:;ZWB6]7g0R#KdcEc(.-:,2_OD.&HgJ&[EPOT&T8RaaJN22HdL,G-?S0VUf?+Q_K
B=?0-B@W(<?aFU(_?Je.c_@DR;VGf^,=eRGRdUV;K<&R;Z;[Q/TGbV?ACI2C,7?3
;Z9V,a,L0ZWP>9V;c0\E\,;18^D&a?BcDDS=S=FVd9IGUN&NI:g]QTFKM-NP3N8b
f]8@?._96F6SNZEOD[]@YUMgE7<PM(4&P,HMfD_e8c0+[a:3dB]LW@?eIQG^<0;:
@[T.[8gY5&aE.c8Q;4_.75#^3@(DV[)])e5Df<X\72@AdZ5^^1dVf45..Y^VI_D8
e/f,5)9AR\20)b4F+g9KU-E<0@9RYU4:Kd[Ke\O1NF/Y;:VAZbFVYYE-I63#70Cg
NaeCAeY/;[L7;(2XGG[C]bNd1gNDTg;4X9COc]3#b9Y()YDO]NZ6/B0[ZV?+bQFT
ANbT-b/D_K4Q51H9X,8S2S_e&MA\MO(;\8&1EP5EA-(gbITX<.(#?-L:V=9V<7.2
cH/CMTXMG@f7dXc5<YP_;Ggf5FF5bGLSJQ:7Z/4-79NEL>4?6;UfD3PO_Z[Z05M(
Tb0:gB.Xe_?g0b\SaUc,\_Z:C^EX/:fa5Z?[:R:SA+L=W.O/0[#A0V0[39UU2?X6
VbbPR91TT?bV_,PfeJQTMCK,KP70</fM)&V>;Yb;TJSb4XASd.#aGEI@-@c>J286
gd>c-W?B&1<0a.c@SOI2GHbKWX(06SGPY9g\,@<^^If[UW.M8O3Q8<G9,G6M_QI>
A\<=6[:30A@JgLg\:OBJRRHI&+1L^0MA)^\C.&\PDL(^KVKGTNgT+&LEdN]RKQDA
\fMJEH1G90fWK<WNJAHMG2JWU7Z,8#f;dP#)EDOa7H0OE3/L(3d7bM1Wf;UF13<C
,NaQ&Q\BB]G6\&O^&YYgZ)RaLPR\;0U:,5_4M&Q<&ZACW\I-@&J_aPW_U-6&4+eB
,dH&<7)1#P&]8IfRQ:2<2K+?P)E+;FGC@\dLaY8Z7,:\;-KJUXG:Fcbf.QK^cP01
W&KT\bUWK1-9/Q/K>,MN[D)dIBa3/OV8T\WD_1^P.,1:a]-Z<NE7?[ZBR@XTA3<Y
a096AFgf6]1bR+CFg:c.I8:2g(FYcGM)&H507<JacRK;HTaVV,.G0E8FF8VaTW4W
d[(V:7V&>NV?<e[;PM4.0gGHZG16GMa;LdJ^69HNMP+XH(_I/6<MJ-eg],HVQHGM
G8]IHP5[FBdJg2:UFHdIDQUa<bGI8S1/8\+<O51HHFF/J>K8=fH-P5U.+=91N0CC
H>V+)HPR<WdG^Lf5_E5dL@-b1EdRZY^HO9(C[GJ0>KUND1+<)SYX55J?#d7WA-H[
F.T?H8IE0C=[CNZQ#3:T)L=(>I1CA?Q)GHSMS#3=c@09?4(]_UdK[1;&^2(J7g>[
6:eSRJZbM6133U7b9c9d\[BDR2;XUQ?8)AX2Ka^/W7M=VaA\7?F,=A.?3>Wb.g::
Af3L4ZffVG0873dQF1WI/c7B,+[[eR[J]@&-(,_Y7RQWf&9H72>Q5YOLR=d/_e6=
PY/c=NN=GHM/MDa3<NSKR#\Nf8R2SY4QcEV5#H]cP;B=06=P8g\.5_LMUc-RDS/J
./ESa:/\8F_3SP[1_e>EKfN5f6bUa-6S39X48>:7?SWUe3T)9PPMI84c_U&7Rg=L
=Cg_eB>6#a^g&-B6:C&DaQ[>CLTa\2L/[O[Kd]=1##SO:[[9(4DPgWK?P.e46]?R
T/M/Y&34aV_S9d8^&BRT^:VJA;44:,6)-8VSU&1Qb][A)74c+c4WTaWUZGd?R&NU
5V)Sg2d;c=O(Ma[^edePAB&H@EJ([]X5^<&>=37c38#2QbCa0I_AAUWJ^TW:B\]f
]CB1^G+/,g\58,=((\X6^LZb?d4U71CH3I:@SJHWe&7O4QB[=\dXJ<HSPLUFf,a/
WAZ^)@+^X8B3CPF1a)CZX;&<3<+;.O/-(M_HH6E?Q7b>6dP(Q,KTB+QQN2UcAH8+
0+&KN35e5HJ5HF-J?N[POZ0Z^gYKe3W[OGCITP&DXM]eUD8dCIBC5^5Q)GcNDb.f
_0FJ&)]PD4KgHESH5O=)F#_UA=9LW7a-Kaf(NNQ1aKM=TbLHa:NA;&6[0<T\A&[V
bcH0RO&[U\KHMTHYWacYKM<DWFLW-\5bU)J&F0)L+]KbEJ2XL&6TPH+;ITIQC6IN
K-H9Q[<G8gO5J]HHK(RZTPILaVGH;9&T<DGGN2d,0/[CAc+0\BM]Pb?ONU,Q+(U)
V65LJEY)M[dI&>b37-T53=RTN:.MLed_S\LY<.Y2Z1L\\_T2+c4MVVU,>@&&L@d)
K)FXXADYeYJAgS31H#Fe-FN:KA-YY&:B[8+-)12TX9:)6g?g\bM1#dg0C5HO#1C9
R^D=IgJ3-23VEH1[=4Yc03#QT[O;973(2Kf1ID]-W;Qa-?>#Uf6OL@A^9.d4\.L,
3+NR\-AACYV_O<6ccJdJ[6M,&[/bOO1Kd+#,<7?f-FAF)N/FGJbC[Z1MUM&J<N_+
]gT#VJGBQLG/\QJ/[ELZ4[X-25OK/3f#ZU7ZBL+.YOV>&g^7OB(Q+RMgT&ADSNAX
_&4E2IIF;F(7bggGfQ:F/e+#JBIS4R5421Yg1cR8UN0fabO2&T,8U+O)&26\XOFW
MC8g-B(VNY40FAQ8T1.;1D4RDbZ@(d[?5E&30R>F:ZYBS;aac\KScfa+)#[3aA6c
a9+b>H0(@]aJ/fGB<-c&]3YN7I9O_NKK,[]MM>@f9KI^PfMQL+/,eVH3HDT(01c4
X9]@3C0ON?f-/fS:OeD2VFRUd&R_MO8\LaOZ=/0BJP0@8fVS_8#2HK_]@?WB9T,H
47?U9_]:bIMH/ZSZ@2G&(]852[S)Z:M-Tc3\)U\WD8Y.J?a.gZZ4ZBdYS(VKg@#0
38&X-/I/Q>@FfNU?-T96T-^Rg94S8ZMH-Z:S,79d41O,_[)H9M.d.^V0bEbeEcY[
2aA9:LU=Mc._+:9a/LGW[6L>;(XI<H5TWK_YEN4;-a-1;cNT4G+(C77-8-BKOZ,#
<P.^660IK]RRc5XW=VAH7F&O=UM,BNRY:4ZKE;GgSNC,SO#V2,SX/SEPXbY176Z2
?&MN=_H#.B@IZ(U;(^GREe1#Q,#SV360>2Q>3g##A:3]XRV]U,.-C(F8/a<)U/S=
XWBfT@[=2,OWMb35C3F4<+-YV=Ye<?A,YEJWXZCId,E34f@<d;LYCC]2?5b8WZ#Z
QbJCO9GA]@dMeVT#^_LPMPMB6[,ZJU4:+84?[7>??^LT<+Za(>2:&1&4=c2g>QJ0
c4bf9R[7(YU)O7^G8/;g)Yc3;6X12Y<C[-(3?YeQ[<R;,2XT-(EYcUALM@4?ab,Y
MDeT0)LBFS@.A@3YA;ZP/1SEF=c0^EI?)N)TYI9[dW8cJ:/8J2EV4dKVb,EDVW>>
QWN#);fdXLPcO=C<0I^[KG.Sc;IL^CU59Q>TMGG,#AJY33DN,4393F@V\,gP2F0(
<03XX;<J]aL3dHD9DL--_bK+YT2[I,](:[R^C8JSF]C:HPQJ.CX#6fM^LcLR-[Wa
b^P#3,T>Z4TUX42I)#f((:HO>FHO./e1Me@]#3/G&>05e2M-JEdQ1WPD[SBI8.YI
1B5_Q/K:bBebI0+)bPec#_1N9<GAO05^WP#(OL5JNbQeXUTD1R9_Z?Z7RbXabg.:
N,^(_Y4OC;9<74#67eNYB1V6KSK&MJ\OLQ8I/.e<X2>,.OB^A&>>-GU?aFGZV#f/
?5&;<X&1ZOEO(U&Y\4ba^_X11S(a-N&B-O<<F0f^OZXB:CH<)L+G[V#\9\L_]ITY
f=>[=FG66PZ[<PKG\\S@YE-^#73V#fQ0F_:FJ]\4LJK/19XHDUXR9SBTQcCCH&SQ
0=TK5AM^.ZgB.>9acDS9P(Ac2Ib?A.M,X758+:,g]R7HC--AcL&O.B,3<B]\Z>fA
[MaedZMTD^aIRKB/:J\_CdO5L2MS58\MeLDH0K&T=I)_a9gJgGH=)]^dPI?JLe;>
:.O4S-fdPV_aIS069TNg[3Y6U0:GUaL>+:&8\B(#6XCaA44D\C,PI^Q6FF[g6SD5
\^d+/43L(]c+MbX4dBZXIXE1H,\9aX:U4(19D&[2?MH:^&A-?;DUT8I?:Bdb4eYf
FJ-CMOQacO&2DWK27GSFZP5A&6+=I=Q4M0gZ_5#CCLMG4,:@<0GfW0M&[0.NWaOT
VC@XK_&#]H+bT\9S_#d3>/71V)Wa5UNOM(T\]#aIVBHB(_&_)KB64Wd.E:=[L,G4
H.3PD;JZH(W=aY95[(aGga[9:(GTQ)5Qc;#0W)FRVM#TVUb#/4,IY3&c_GD=d9-/
4e?gYJ_MbFa:K^XYYA8.>P4>[9Z+&)^d]GZNd(W&T^]Mc3XCYR\X274,Y#Y+2AR)
E.bW0a6C(K3RL916#fJPd^H97R6&857]N)S2N3G9P#7;H,C2:ACYQ49O8F(dc:^L
T2R.+FBC+22Qd3JJHa2-+[:[IADU@ROM7)4c[S8&bSa8(eLQHCT\13DTB0/)NS9A
ER3IO..JN3/bb7\QK-YFYA+[WND6gI]#-3?ETHOS)Ace0->]5/5RZ+\gQ1_IE>b;
F9)fMH/B606VeD.4V\9OE]1VYgX2A#=71S],Lcb,V6b^Dee[8,2ffLROC/c+0KYH
?>J/eI@MCV,:(b]GD096cD&XXQW_5&2^H7Bg?3c8bH^CFB1<UYZeDAQ,K+,Xd16[
/\d6A<2K2+-HcQ<L;NB-)fJWSL_Y?#JZS)K.[RaDK=D^Meg&G[g\DAD/24P_Q^BL
&C+PT_:]ZLB,VF?1eT:/OFB4(e4-=db:N,N,)dI8@K\\48:Y:&>LdYRe98#E3/U5
+J&SJJF]JIXB3W8E5O6Y[9fV0>+J/-]_)]>;QOL_G7C13f[K1+LASga<c3M7?]EY
[\+=\;@VQ&X:G/7V._^1dXWVKN.3;A]c[EQ9SH>UOW<22MTOJ&fff..[9##5(^I7
efK8DaKeN&gY^g+a=U@S0>54(Y[TQ@?1)g?U+02H>a0[+b4#;g41VF=)B,c>@]I\
a(T)_=U+ACN=8fT7.WK6Q-W+[A<@<^@R;Of;e3aL:+@5M)Q(82(-g7](6=;>[X6/
P#KE7S#6,]6UMc0#<N^Q3d^X-fU27Dc63.5BISd^e3[2<R\fNR818c&/bJ55TAZR
8e#B_13(CYeUNFTT^/Ee/eQMMD:f[gST=]+FFJOW,QTIC3<J(6MW7=&1WK_Td3;B
=VLW5(fXHf-SMRG-M+g:RXK@_fW>^(S8FO0eBHCWfJX&:7g7eJgWOMKa[HUc[#4J
/D#@JA/87WAg+eU/PUW][7e7gX(I57EKP:\?GE8Z;PQ:4Be:R(>cQb6KSV[YF58&
I+,^dJG=4705G<7S=D2GVJd0g<6eOdV3NXS>R]R]8f38>5,55g(e-F++O?4T4DJ1
eLKB[O?@WI)POK0[b)0([-GWU#&I[1APVJ^7XbAa[aTEOBU-=HHa=0J-2QMZa0^(
C,C_X6(>L7T1XPK48QG[;aYg=c)gGKE<[P)LB9FI3e)58=HV^)OS7AJYR,aW<_eK
Wa/Gg2_.5:YKb.RRa32d]VPT8dU?<OKPfRQ6CT^4d2/LIH#F.M_<>9]@E?cB@d+F
QSeQ(a^Y=L0>3\<PW;1TAK&T(ga2ZU\I,]U[-6MJWVUBe,c&f9Cfda(X5_NPL-]8
QZ701>FALg_#G3Z>-&K:Gg]E&8X[;g_OP,6g;>3]I,+3OI<W;BFbEdSf<KPBEg=E
E[-=<:H5,Tc?GB7Z3??OHDAF>DcL;:8#(MA/LE5GWdU;KaB8\(PUR9AQaS[X_8N_
VA2CA3ea&7)VE>+<)^&5/5Ob;+dP:)=P8BWF_D)X3bMXg1XL]<6<B[:Uc:NI0O7=
S158edKS3Y@W#B948A#&;A1W2#IJAe/M\bAW)1dRSe#=H1Z8O>PB10GWe=F<c.(B
>H__];T=fFO_-FH4A<ZUQ^a7J9IRL7\fI&<Q,M+:LCGM9\Z.fUU]6L>AW.e5)ff)
cE+PXHZ5[J02\GgPWC>1#/DCFgedCc)EPZZ3X&S7L(OaBH.5WK4M0<52GFH,SM\J
EdS.d8W-C6Mg9eVUe[OW11O7fe+Z7JA#9EJR=BXEOa:P3#W)FE5a74J72=ae#7e]
#4S+9:eO&K[GQHPK)^Q_R^\5V@2..d+FTG?d_@Db0:GQ_?aXE>PbffaS[U^a:QZ-
^b9R2d&-8UY2IG4CP/F1>6#BOd##cE9X5W+WI?]9NX51)>.)bS/F07dT6R#Z;BO,
N-K@@+F,V\D:HXRI=_&[=ON>eC+78)->gWMD(][YU.BX=#>3P4\IIaaf^]8ALJQG
D4;aHJD;+B\:H_8VMG-5gZgT);e1>V4eN+(DT2V#&SWHTPX38ZXccRM2_>XR(&AB
0O&)1JJa?dfe=K4g+&9eSQICY[@+C^CKD<RGe\0#:>@RgPVWH#HeBb&eU\+RAR->
#9@B27#g3V1(F8S55M5MV=Z_cH#IO&OUG>?&V3dZCE_KCfCHb9FaP..Q,/MIC/(7
\HRa=R^gFQ,&P==5F]A8A/;DN[GJKE;HbeIbY.S#][);27VTO4V3YF#M^cW.&ZL.
JB<R5-)aeUC3&Ya[J)1)aM#=G6RdC=Jf+T#Q-EG9d1a/aG2Y+/<KHT1a[If1Z]\-
EDKOCIQ-c.TM===PXH(<-<V4(G0HBaJ(U)F3.RVW2ZTaC@@SM++]93CWP8MPUV^#
0E,EJec&332(52#Y&6@K:fWX7F0gHceBBQ<=4#ZF+MUgMBNH[K8a_dYWWG>3D)ca
_4&&QaKc>BJgS__dR5BN/1FNWRO?ZN>U,IGUDCY@6bJX=BD+g7+UG1#/d.T?SQ)X
]Q\6IYc-EXR(XJUV,?XFQ;^OUJKC823KURLB4M15VJR]4_Y_Y\5JZN;98#;SF?HE
TMPe<1>-CHcXR-,\BYEeKRJ(LX3Z\<.gS9(?G+HQUT5NLQNTeVAM3g0];B8(0=<+
>04QMU8?Nd[JI7,^EF0X,>BA^V<3CC&J\[YW&a=]X?(2>C#VPY]LDQT)f?)JC5W6
1aF,Af@H[EYMX;+33FQ^3N1UcG&,=0&J?0]Z9N;NWP6G43;(KYBe7-_5[:P+KI.L
AB<7NIZQ>?&2A&eN?_A&.]3C2,_5L&7ZN[A5N/Ug#MYLg>;.QfKZU?\836QJKQW8
eBW#P1BZ:(XIG.:DH8NSAHHJF\BL<b4(9d<-/7(&<Q:(1@Y3NBQX\9_YI+^\;0AT
#3MC;#CIeZXW:ADGKBef]ggW4[fZ[V^CE;B[&8g/aCP8-=MDUd\TV/C\J.]4^E>1
cJN<Z(,YA+R<.f?FJf4^5-WAYU0(XdNg#Y0dQ:E?FN;(T[V#-5_1&d>_g_,],4NY
06MA0Eg-NSJ[77AOdEgX6(R]EC1LY_4c05@1K8/O8C/#-UEf)#:\]1MLMa1+/8DL
Yd74b0^;3:gb4-McQU?8de/J(.g,YYd)13L@LE;e@\1VFO(ELb;_C]97BLL)G(+?
?9=R;L4@U_GXTI46\-AV#0=LJ\<#aF>d?6;LNbO]^DPX+;UR?=J+OgcIeJL,N^#@
c0+P(SG:X@VR.[4OFO6YW3W5aQQ6b6SG/cfe@S,)9)254g&HJ.O)KEDD4<=/M;\;
/O)E1J?GF0aI0)KDVMH=M-^/(8QPd5L:aMRZO[(@02)2B8I3f)JOLHb<cM_QGSg;
:BQ9)FBANfH.5NDU4HUSa9U;QA9X:EcWM&SLI)3&HQc=A974@f[NZ#R]UPb2a&[B
6^L9G7TXBI<AMgNH+)<ZPAg/AfWCK2(F[S2aFDC2BW1=8S1946S[D]fUA8\Ng:ZI
LC+\?J#Z\]/1IW/CSPY4&dBPY[[&#W:QfWAa,V6T054L>4&6=)Y=M:#LQ3L126N&
KTF6Jb4NV=4&=\b=6NF[bUcM??48ac>MWG1bW=I2>49SVR0)D+g(,^,6]RZ=[:RP
&/aB3-,f#:<1_B07Z0_a&[J:#7ePUPVP@S<Wg_#dBN0?b)[.<&Q6;&a8/T]Rfa+:
:34[P>X5+.7=6,a]2=>4>U)R7PGU=FT5J&^/5gZ<4YC=6f]H@-R4c6O=<#-Zd+<4
#H[].24\bFW4;g(LAEaNA>:77OJM2H+TBC,>D38MTK?FIZ==\BJ70RA(:YCfU-1f
6#06Pdfe0Ya:E^9I=OE_#1T6UREUDS(VdS8F)[W)a/g30D7+^&\c;Rd?2AX6D7?M
\\37PdLIV-)&B\3L,X9W0AcL-V4Y<N:?WRH2Mb#?A^:R)dE>FJ;aAN.+[U[T\3,.
FIA6::#gQZC&CJA>03TRDJY:XLeb3UE[BMU-d4+X#bGS,SGRH5\.UJgO9XB7<@AX
8IK40JLQ3ZHW&a-,H]=5f9>FM539YUOJQRe4\R37I6d@V-:TG^IKYF2T:D)^JRUV
Vgd]+R\OBJ)WdO<V.G=.d5Z((B<N_U53R.aXSK^OHK^4W4;/1G[LQPa^496>Y0H4
5\]@bM]Ub2N=OG2P9A@W/O/3CbWV/gKL0L[14ZXBAOFZN)VH#R2>+Wc=B#V[=/PJ
I[=cMI3D6KNT:8Q@NBAPTQ2dD3C66IC7MPN]UWdd?1VOAX-/+g8aW/8]>0K>R<e7
V,3=\f15Oe,aHF3],QEc?@H12X&2@^#795QLN30ef_E/0,U.]K7#Ig?fL/?9>7D)
5dDaU,&+V[P/U@^.2)M0eaIE2g[^06:EUfXR2QV/KG]cL22,#:@Q\V86>#^G+gQ:
+6RM4eW;L/cV[G<H@S/C8>RJ(1-NK-8abQIT_1JUCc2Q;SE/E\,Q-DGAe-B1B3[&
J9;?+Fa:#<KNL3(U;AKdKaGdU.Q]Z>F9V2\VCLD>5JWSZS:8@C9<KH^;[BJ.B?([
PSfEK]C#;>FX5;>K3a\8/6NAHL2+]dHBeQc()a_d:AadFSX(baZW2;@5_^#2F2_7
C#WO1T(_gd3Z+@P>K+IFBXJGP,F.Uc^]FUOYDY3QB#8YR)]+\fB45OO<7PMHSAUY
V6N&GO7T39VT8U@dUEC[>1bdN@N67(?BJK2)]DSc60;L>+<J_Oc#158S99G()I[6
fD4AA3.^>/K<9LBCc3<Y[6Xd(YfbOKF,Q<O\_+>MH.2X,?Tcb:I-HZIZLNBN,5)H
?(3^ZNFJ191)+/ef2Lf7I>8NWN-2.U,:B92[7QN:)&U(?&c>f>L:?GD3ZQ1,0?9/
W8>AENU+T[e-1S,81VQ<@#2H:W8-E[,&]]SSQ<BO&=8a7#RPaXZ)_J^WBG1cQg#e
SQQEIUXY02?Y#(IM.BI@c#LY.[>H;cUSC@(A4b<(LY,775<B<>MGcSfPA[e.gE[I
0B?X=Y)cL+^6BI-E0D/T548Pg.X^3BQ<>cVLMV,Ya,Ng(CQ&e#,GIN5D3cO\e,D;
_&Ef:SYe_IMVLC,(BYFY??CD+]K0?R>3R?<8b\2>O<?QT#17VI/I-\F^6=U;gRZ9
=+BB\0E.WG?,Q+7@P1K+a^1:1VN]]XbUW(acJ;Y9c_+Sa7e+ea3\/58OQ@\5+X_X
XFD;<,_TY-LQV:[FFXA;#YEB:g?M,[/?,/:VYZSMUTLW2_eP8:_?))^FEF)7U;H&
SZ3-QJ&OXa_-c3=9[Z#fJT(?OaVbBNTAOK=FR6V^0A_ZEBeWHdN;]RC1KLJG8B;>
;ZTed@M)LSU7NLG#UYSD/\^fZ_CL2)a#\<YN8K>.;A)3&d/,M^8OgTOaWT[6,7IX
eK8Q.,WB+JQV14aXUQfd=9?ba80^_#X^HaG,QI06R<2T9CbT0g#K/&G05N7V<3=R
bTU[^.=#>GJ.Qf_&SI426Z[W=O/]^[)R]YS&V_2NdIUL#Y[_S7OULO\/=ZN&>Q]5
N)N(9bf4C767eec7D;J[S>6M3AJJEb_1gAZT;OA/BGM7WJaPF#[/>VTC846P+b2U
:2OB98[]EYYHQ\_E?e,+Z9OI]Q3R3V/a0Xa-26-2LS@bJ/(-IELHSWSQU;WP9JSG
AdGM^\.X.BT[3<B=.e[WSN,c(Kc[?\,56W[VSL>C&NWW;LBe,(\VD@N8N3MK8TD-
+a(Ie]g=9ZfRTD9.Y)\Q:]5&[bFAJJUdS4bHc2_#eTABOYG7H5K5(U<gIF?cR_?(
#U9L-#f88^TMO,=g7@_;a[RM3dDF8eS24+D+ad[W>f7=McdL8_0FJaO00=;3e^<@
D;0E3?>g;F2+BR,-RXgJ_1Q>,T<g[R^>aKQ3IGDQ/&[b>a>ZO0Ga^GFAL?T7L+YT
8>E,dD:-=W,J1^UIcf_BgQ]S;;eb9\>60;fg0Q#fQDb\7]@d7=[GP;e2+36SS2Ya
TCBO?\N=L/(,EU85[_,,0[/LEG2a^25LL4^&.Za74Fc9L996IWW=f^ZG1OX4&EA4
P2EAbZ?B;O6[/S9Q5JI:@2&SR]XKDH]9:AE7GQNTQ?XGFIJ&(C[Z]eL/Da6Ua0_&
<B;/bK)]FTBIZ#HEIA_fC@3EK3baFf;]#L^-0aTM<eT<6S,H>K7,@bSLRI+CB_+>
R]E1B^4[,+^MD>If<Wa6K3S9cAT#D_AB.\ZM_9cLHQg#)b\Q24,f1WZ7fW]H#N=?
I:SXIL<J1J30\K.IgELB(RN15:^gBRI_O?9HFH;@#-7MTd</XbRPN[?bU8QU=1;0
Z^6+PB3O8Dd]-gW=D.89JKaNO>?E90f4EZD1<^ePFc_OYA@0HU7a2@cb+-,J<=<\
gD#@.S)LFYU-@YL/N7M7B8<M9M_f1-0f9HG(6^W0&R9.2OEV;R-U&N1:^,U,53:d
,,640Q))1KB.:P@/3X@5QU@6eB8:#^[IJ5T7FPZ#7UYcY4PZ(;2VO:?6?3+\K0L1
]^WIQE+X5X,J0.3(9+T/>UX1^9[@:S)(/JNN0[0<TQec,]@62X.SQL>YX)b7EXdY
Z>ZEb;-V8(IfJ90AYaE0f9)+-)S=]&0<fRR1;\S#a(O\0S.;\HZC\Fg,.+:5>+QP
-O6(g]Bb)BA?2@EcJcf><6?d&X<<3(IA4?]_H2,bT,U\?@G0G3=VW5+aR0FKRG5L
PL>g0L@).K5IbH5Z-Z9>@>[2LVN)NCcYd\+-78Y[e_Zgg]eV52^S\Rd6TJ2CdIPL
^8P[RcAXDMc0E.>fRMb6g&=4_A/a(+CWRL.IF6DI2(FS57_&^@)W^KSN(/BGHf>H
C;dSX]B/8efac[G3dOS34fHU<Z)R&c)5VY(G[NK&ZSKI-IaG7a:a)-BaT(d?+[M=
P4LH7D4:V>\8=LU0&Y2d5<<H2N2QfFA0)U<NF>(cAMY0(4^J9c-d5&USfg\DMFWg
ZVT@3,5d_?gT^M2>1<#IPO=Q)[&cTC2<OPgWWF+D+?Ke/;_04:US(aY-dF-I[M@6
X9dBA0+ddd9f;BN;e[G5Z4;V8@621R(OT34V=\YUbb2L\R=<XSI8=66=2=Da68DI
N(5\^BC62a?<9FGYW2,]gcU.;AJ)>f#UVJ)D6=;.>6ScA:@/4<7WY-d)@-0?K3,Y
6A6I-1MYSI395U,CA<L7T7=3EHSC>6<97T82HYM34?LVD9SfN?M0aOKfSaf,@9RJ
6g#JI(K,c62C6]U)HcJ.e@aIVcQaDNY6Pf[DP@KC4SX4HT\+34DHU1Q)HFGA+Q#)
S=;e4;9ZAg(aeZe[0N?B?LTB5E]X]5eJXME6S&gDX5@A>V=fg/3#e?VE.FS6^aC=
PEGCfCBa2+?-J08Ed5TM1SaHUF<6(W\LQ9-2:UYED7)YD,T8N)QG:RCCL1/BI=Md
S?RdL-Z0Qea_V4gN9>?05D=H-L(ECG?>I@JdIG=RC3=@T?=FJcQ5_H(#5\&&CaR/
I>BW9dS]#E3.6;RGZ9I1\/;[RL+J9-ab4M)#5Q7.5BHMC/MR<E3DD>F18[27eaL^
VAG>OaH2;.8,U)/d,8@O/Y&YT^W=8JO4?5#NeAG3?9]f02F6B3E_RY_=E9.bE-P0
C>>X.QCH-R@dG+.XNDSQ>)E.gE.+]Zc9]T6T6;+@ceT)HA4DH>g3A.E]#>_gKU1<
G9]LSL];-1HGP6S+2PUE:XND+CF)Sd13H#<LIa<[5]W/]e@E_d7b_74-5a.FZb@A
N8O+AV7@PYRUO9/^(Mc3+(QFg<?)8U&).,B0&1F0E.Y=18d4@JYc_N4-N$
`endprotected
      
`protected
>64OG5.M;Z&T_>KPGBE;1[?Q\7fY<1Y+H:?HRN:C8=ZL4BZ1I\)E&)C]Ng]:(;PR
.cL0I/e7O/\TZRC[#e-O5,IX:@4b+]bLK<Q#1g=U,cS=U&#A4YfV:,C]L$
`endprotected

//vcs_vip_protect      
`protected
Fa5R[gVH616We4^&FP35EA<^begbc9><7.=1O@PX9)YP--Q8QSe1+(0R^WX]<d11
955?EP98V5d7e1/f9Xe.W-3\=N7OPaAY&5_Y:c2&@28V9W3JC73f0,-\ede^-f9#
9-Q>69G@BaMW9HL\ZMA/9XNZc[8\U;<I)ZbV&&YYHLSg_(eHI^5/8ae?1H3a(3VE
d=bXJ?^Zabf#)_98O5XLdbJCCN:U^VWf.1g5HMD<6KO5#Z(KGVX#>_Y2@;DVG69;
1SQFcJ.>CHO9/)EAA=.F/gAV[RbW(8G>NJf1^J5b,L;I>M9EL4Z4LUf4a2<T;\bS
AZ2DdbQRA208Y4YH>IQJ70@=(WY?d.fUL\RI:7aFT4):J3<#4](6Qf.J94KPe.&&
MN>L>I@R8FC7(Hd2VRf&0_g2GF)g/Y3XR]D>bNLJDg_6a3+_+Q_8O3(#QU/E/F-W
H5c=X2(Y-_6a4J(IEH6MA_A]SZHG7dCbPP]\ZV2X6(USgR_J1G?8&EJec-FE6I@,
)#:[2aBaeX72HF>:aD0Ka+.Q#\2fL,7FbV#W&S[GEd+4gU(f]L25.LOPLI3MM.KX
6A;AaGGZ@/?D=,.:BcA)LaWCQ[B-@Y\L6/VA_[6&B.P7F#)2#URgGP7Qgc,UfYa1
2DN]e>CYb_[YKd>2GGbHLCQaG.EDX0[^(.g2Z3f,:\4]-C@(JSGE4HXB#4bJL11U
\bR)>0BS\K&(RQ^A;([]aB;IXNTg>+(1E<@?#DcQQZ1(UVdC)E?T/JeUA8/?/E&D
R_6R9+SIFeP0^)/6>9P]^La5U#:.>/:>@C[\0H:UJNOV5;MQXNL]B\5(P;&,YEI1
?\TIbC1THdgeaS^,=AFTGf&/VD,(Z[,(:64JRZSRJ<?-eGQ/g_@5/Q4=H^N)[OcH
CdDOWXDHC2DFPN<f.@7W][,;fDEEf/\#^[2CT#F\5Y,Uc=K(<MZ9V(9cX)3IWKbW
c_6D1EETG-?2>4b_1F6=C?YCOSWS[EU^X?KHPP(-FO_1CW2(1fNSH.=4Yg31C[1/
>)X+IV(A8=1)c1#3+A=4M\YFgWI\+LWd.@9\=5?cbd4-I82)CIM;cCe[M_ZPMd7Y
K^#/XBZ;V]\aHg\W=Z(=8C#0gQS5MZLf#L6C./gdL\Z9A239CR^;/++ZRcPP#1;,
,Y>TeP2b_eHPE&#O,;;\IQYJf,-IK34UL.069Wa7AG[(@M/VRc.295?20MdX5;8?
V4P=A(Ne^9J\53?>-EaZ1=Wc63G[;UMI,>fCZC7f<@IRA+g>MDfa<LZ5G?F<1P/+
#_99B2:gF[[@bQ9OV7+<6^<MWIa+.>QJ@<L&1d7V1\?&&BRQ(T#&.dg12/FX#(1@
F+TK5>)0(:Zg[?3?IaUbO+=#MM1PGY9.YgO5ZD7.NQC[bX3WL?^ERFG2HJ5W&_eN
MP6ZA)f=D^I)#YHXX6&)H,DC\9C3@_)=(,7/GFf7Sg23OBC2,+[S<2HZV)?XA-Q]
P7ZX:X2aH4b4Pd-+a@]cKX9U?V24M?_LW5_B;OQ?@)J(I-Nc<GLUeZ+HX5<0_TMD
#NfJ^D>I>--QBB?^FQAJNgA7H\(<f1&Y&Le>I^MQ.,(7MV-U6V(R[OFJOM^-<8&:
Hg2.;BfP6CJ:(B/,]S&N(34=]bU?HSfS8bJVE:^O7X^0\,UGPGfaU2.??(5ZWT4f
77#bOA20@,(X:U5]DDe?DC).SJ+59^=^ZDQ-AGJQ.<dcJ3\FSA_C/TGY6EP?K11[
WAgWI/<_@T:S_0N)8;5EY6B;f((dF@d-TNb]:-O3cA(Y\>-cEVG_UAIPUUF8#BE2
P>7e-e#JXHKg^47F#(&HXQ@ZINfBP3N@NV\gMO=#fG8CIGLRPEaBF[Z26+QB6UBe
ff1OCF:^_4cEd)3b0G7dPg19=4AcULQU>]B-3AX;[N(L/L=RV-(K0.Y?8NX69D:>
DYAb@gR7Y7?T@N7P<YecR?M9BgJH6:X2AP3KV8Q3BC@fe,D5EX29)?:DCM8(NcM)
)a#Z_T4-X0>3]Y9d5ObLC0MNPa_DH=-TS-,d<WT(MY_H2>9_)DG;5Ze,Uc;KAQLS
@0AWRX?J++GHgK.#YHHUK#e:U,<#U+B7O]aa?Eeab_&=YBa&eRZ+ZV+O9-X9@K=(
;,#T,8C/XYBPa#S32]2,If+?6&J>gS@(]NL?F5HM\>K_Q1H?@bLR0,D_02-DQCT6
3?P3@I9M=;/F;d\.833ZI804][U^7LcE:e;O+IVc7M=bPZ0M-]Y>8D(DP^Ga(Y^<
YB&#JdO-Z6>)C=Re]#5OV&A][MKWcUV(e#b<ZZ)I(Z1VHT8\J:(Mfc&1,[,?Oe3T
MCU[HX[OdKDbL/,RQ=5UTBc7[S42X]-<5AL^0_].fHC+C<b&)AG7fDJ2fb\O+S.M
S^26WRU>D1-?Z<K-K>0TOKD))U&6(NW@7gJ_#GD/4W.&>Z?D=0GL?.,GLG:RWUJ.
>=#FL7?eEX]8XK=BJ@a2+X(1#g+a,G_cZIJ:<UQNQ2DOQWKFHWG&bWI[[8cTV:^2
K7d#L/Y/U_2L3edF(G?;;>\P^67/E?CE5[F&B(aZCI4<LX2_9=+=DPP7gJBdS3gd
ZESAb8.:13;PQ25N/f-VT]_4(]5&b2]8X9KKfMT:\D:>/VAE+YQ_WZSDE-(H4UGK
e/R&:DEE(=D-aXFJJg?\5^0K=.W??A21=V(-RM1?f5;9b8L^>KgaICSB_9ZOB_8-
QA8Sd_+J/4L0MI(I=89LZX@TBc^B<VFO@JLMJ]N3I+a@gH0>_7KfS;+DaF(c0a#g
C&47V.D4g7G<8?QSd,/E4IARdZAdeW<NYfI4N#UgbUTWRSLc,,YB\/F4bEf&;CEP
G9[(&[66KW-#G04=;>bBag0#e(&-P,S+[Y.:<FRg96RAB5_D9R[-JJ<PA./G67g=
=@XN;JB]<3@:I^e8b^/PN^3+(g;eBZ(5HffgV>7H@W2E1PN+6M?2&LG0<SV,M22#
QOX50BFKZ+?UDJJe(0,T(-0a0?U<g5L/E<dXZVP^6+1eR+FEbQ_?M;[(G2\.aW#:
]bLYKM/7\#7]0:[;>c+N\dCE]EF-8L#bO1O32IJ46@&ZFPg(+C<E@__>#HM:P(Ef
VXagS9U.^Sf<I<[K/)dZGF&T5Je\UOO;aJMNVI3Od5(\J4I177\X<f(.T4);BBB(
b)PWW2L?@X\N6:\BH,&X=T1&>&B1]Nb6(7eWcAXL9)[C3XYL)H/C?f[&=4&=LJ?K
:_/4LO5Je>#5F,6I)DL@,5SRI8^efN7\4/NCd^MA])-WP6#U_(f>X3T-3&7eM_3@
_D9DcgB&SXcR.KcaaZGgIJ5\D>E=/&,IL:ScW,ZO3Kd0_<@4.:OB=R@;&KAFB,=&
ELV7^(F=^Aa;c-Y/,FO71__M<XCL:Q,UMM2eG]0-WZE.SFTBGFQ=SS>MFeLaTN],
;^c6H@IL\G\PHJU^C=VN,A(P_R2GM\B9f(3@FK6X5LI4(+<Te3L#AM.f6F>E<14#
CI<WENW]XA?\<2==+=<2C-=6&;;NNEd5:[B9J<-g8K?PbC><>#(DaSB9/e8VEZ<N
_O).E@BO>WB<&B#5,d0+I,JGG=B-7,TR?_E+KN(2+M7JKM5S4_W&=L2^NW;[G2f/
W#;5#.,cOR+bQ:.K+cfd0<gaRG1Q7&EZ)XLNZHGaN1aC3VF++I:+,SIP6g@?GA1G
]SV_YZY;I)_7d/gO-VB80P\36MHM(b7^T8P>O;2d;S=GQVM2@WP4Z02/g(&:\7HG
S:f0+Be3_9:ZIM+cfdW[9JP@BPW=E/KVFCTU^K@-Ta1I(CTSeWdP/_T:^N+Ue;60
7V?5I7@)b<HQ&C;F8,G@d4?Q]_a,C?A6e>BTe88bb>/D9O[IK2E#KTG@MK7<ZV6M
#>C0?.ZUG>DL_S8Bf\e.Z)_Cf^<2@acR#;A9&NbCG9D?:4CY)Wfc1)7N0DNLL5U=
Vf,M_[2UB]R]^e?4?-aSS+BL<L@SDT-GHORV&FEAXQWYd-WV&ZJ>@@2A_bR/SMOI
)6SI@=7=0A29.NGSd]=DL/CH?L//Kd<O,,2gf]Eb+QOEEc:W)6J1?N9ILFW3>A_Q
NT?=:/9aDHW3FA3gF?1GKX1cX2F\=fUCD<\F]#90J(ZcN,&&)RgCO#V<+Q-.WQQQ
SV>18d-@JBa;,YLVC?(g3:ddT@J^:#1D8Df]-[4;SBYM2(:KbH[O6e6,eQc,=20;
&Z+H_-0g;E[]\3BMgNO,c#TfZTJK[PVA=H0=L#E,fa^4LJE9:5:P?AJ@,We[US&I
+_^/d?A=Z,VGK_#eSZ=KL^I?UaDZRPf@=WGPAaPJVQTdZ49^QNB(K/X::)B9.[VU
Y]ca66d.3E<?U6RW(EORJUS_Pcb]e8GHTaG<WQ?_[cRe9a4bEXGD.AOcH,UKY[-1
G&X1SI_X-?IK;?^QbdAS#.&C.V8eW:4+)KD[\a60Q0BNc\-=LD9V5B>3^5L<110G
9);>2B6,@U;VLeE><.dP+[>5.eY7<47)\_QGFeY?a,YU&12DL_2gZ:<HWa:)dUIV
#?U0_XRZ7;)WJ8N=U-a-f<CE04RFVC;9P2PNZ8dZNVU7SK]=/S@Z_V@_3Yg4>38-
O_[MPf3C<K3E1UBJ=7HAPb0]JG@@W=M#@,XTf)O4Z(IR^QZ0N@P:<[^]B.,\7]fE
B\P^G4>,DF[7KXa@#LK2AWUCdZ=)B+&:5I7DJ.f#(3PG+<df>TT_OQW=bXD\/8QH
R2XX<(cQF;O8_.-)H(+SfE9\R?]=2A=,A:RSd)cR4,gQA]3aZX4e81(TO#8O9Z_B
ac49\K,?+[A.\=?^17#W,DU/OX^fVTb:K3]I&ae0J^S_>=?S-)6LLZ>/d<Uc2BD5
gTa9WF^2e;c5Z0[[86ZFd\ZgadH>]_?IDBU+W-Z1<:J=43dJWEZ23/4d:@U<g>L)
FV>DL3UN#6/9.-C,<Me84#]Q.G1@(&+-&J+&WA:Z1N[XgWd5Z+?(V#:=LW>J#U[^
FGa/PeK[=gF0K4-8:@6SOXX;L<Y),)\HdI9RT(0D^TPMZI+?SVF6D#VBP7=VPgOA
CbT(B.LO+SgPeQ8(^?V@9#X8_dZK31OPT(_#[X+cO^-HLI-2YKUg.([-Vf:?Re>I
S]\NZ3.W6)]0#?f9?d?TVb_1.^e+VJ#B@8afXOM@Z/.-=<)6NXGB<VgOK67BM3gE
-MA9cJAa+K/S13^^/O;<?c(C5WAOO8NJF^1]_J85c8@=UU3C23B>0<(Q.-A6gF_3
NEd5IVY5f/Y-BFM9L74^/FV54TO@WfG<TbGU+A[QJG^S90([,],0X>TcH?BWI.TG
SB<#\#.fV3/S:YdW+:PN>#/B6KGVZ.b6;?B>(XVB//Z9a(/3MU+eTG>[Ic8<O8d.
DBLUUG?742N&L(UU=gR8GLY=AB2OB>P,b0R4AA>SIdJXd&SO/5=#B4BX[(V@-a6?
VHYM)e5B^,V;,]SUT2(0Za/P/Ya_WaQceX^,(_>1)BaJZ3AX5CFIH2X<LbJ/_a^\
<_&(XNZ5W3g<>R7FI1BXKdd@AZ]Ag?J)<<#KC\ZLa15D_O=(c[CLPY<C_cW&/[3,
cSG#WX[3L/UN0/4H[F-g)E=O551#8DO;FC7]WCaMKH+>5Z1]6WYd:V42/d71X,3b
.WM?EAK5PI3D-ZAO>WfP\+b+<YV76(HQbSNO6M+U0C]H<UTZ0fEUE&)@^^+(<-e>
X/K@f)fS-V#0FE#N:aJO4)4MJIVI;:J3AD=PeO/JG(3S/g&W5[F>M3+I-;)H6->g
ad_T)gG7^:R_3-W,6dE/A_5<+c=I8#YA]?0SZ5d1)BX>IP3O+_Mg&T.NSV\O8IDc
,@]6+QT8\1@Jg6QeRP#^Je)C,d5K8YKJZND0<I2RZ:#N).A5)7&\D3&VQLe)KDKV
O\IL@):XTG(:[ScOK1T:0N<&^H73F##0JA<&VQ#09Q&g+cN3V+B#Q+?,)-VAOUb3
,L2/.#=IL6]],7)T5A\A;E70^&ObdLbB.GNZLW9JA@A;7:Xe2#0SbQ;?JCb8^?+O
.4^-f9/DcgJ7:NAR,(+c;^++38\>O4PO#MV#G^2]B,M31A\XWU34MbeU:S()D.JZ
.O=c;03+OJJX,=C#2c<,[2Eee^XXB^5MA:+;82NM:&Lfd;]HabC+>+g4B7b-\]\[
BL0AWAR&XF=Q;5<99JBL4[c=H2=#LPg9EB]e?_cDAI9WH6]#HRCVP,XN,]JL4TKW
S^_4FU,R<,cS1B&8>39ABR2F17dLc-8SEBFL<6._0H+N8K8+g@SDd>Z@a]aa3ZMe
Ofdc]H&K?D8&?D0F2)WV173b/)6XPL&7:@CCbY@M2c2XbI>V,I^]1-.-G9]_+XWb
GQHA^^>X=UE5O;A052#JK98KWH[VD8IB_7SFSYOQcDT6gBD+bTM3cA>8JJ9R058N
4R<D5R+_#.c,_e(NUR,GYO9E&eVN@&NP?VLJC30?11<)WE^]Rf2ZaIQUH\TO,^e5
gIKR2,WXEPY\^/XIX]C>3N9W?F[4YV&)cT(+W)bX>c3c.Vc8:T_M<M&L;:J)2?BI
+A\.D)C+I+=Y-4Hf5R]#QgW-=-UA,0&U@NPaMXINV@Sb9@bCZZ;A2:=Z-PWZNPXg
QOSV0-A::7UV[WcK41QKNDA]=5#B^91@\IT]]/[Ng-\6TR^VgfdQ.S;L=+YA.\Y6
b.abfdc^.:MESM1/-=dN=__YfX/WDZI91Z[AJI++UM:OR<eX8V1(-;W8feFN2O3a
d</TS@@;fX\.W1;+?+.)@^:X;aB+6Y_RY#:-PAV(S[K,C>(&CBgI82:-+fd)aDZA
&CT&;0C&3+^ZFg^+>&XeGa^^/0&F6/Q_(Q2P@)gHD73+R9c^S+H6H<Q02RAO&&N8
H.&WaXA)bD#ND-YYVfB0fMTO.W>J#E;aJDJTB=:<)&M4A#B#_=+YJ/X,R73d\70c
0a3,aI#K+W>+8OY9d-U:5XUab#73LWWKS:Y46P2)FM4?JL?G8-dEMQJd8)-e,X^a
1Q<Qf=@bP0Y/[-8b:B4K9B>c;JDbSUUCWLS5?/)3F+2TWD_B_W8,YWBCf<JD5R7D
]WHOQ\_8@P78UV8U;bCFQB?V[[)D._1/U4]2d#UA]C?1B<B]?JJPC,@CG]XCZ0O;
MHF]bY>_2G6e,3WC/6FSBAGMC\g(EKNN=C#C-d<3A_M+48O0SX#g;QJAbT[BJCdL
Wf\(^5E<AeT-]V2[&?@RMH@XIXCHM__WF+V;M]\HKc-1>Q1^&,Z<KK[d(>?@;\_;
[TP[NP+82/EGeW==0f?WA-C-d_>BDU=Ig;_7Q<U?e97UDMH>9ae0;RC;]IGDS3FN
f<-C(H@W)3D=G;eHJP(2fMP&X?T,JW.0K#25&C0C;?:#I(-QTHCLaa;N+2Q1[XV9
Q2R[cYV=82HN?fb+e7JIE)@U.?e1Fb][\ZBEV5U8^\F7<[VS1IcVVCG=]D4LZ9K+
YHCdDRGT^O4.=J#KM1?&7_EMH/8);XVI[ND[+fCYB3)I@B1VHgW6C/08;U?&NS2S
IaL=S;NAD/XI/[1VK9@-:A5K?U57<.:BN^39>9(0-.U7+IF0,PD#8f;g@d.<NC<a
eA(CEN5]6b,,f2_7]2ZD?W7^_WCcW0S2PVCc]R]77TUXZR?X^BW.aD.2;0WN:)PA
FXb=:_DF(2_0@PP8aF[)@?)17[L.(7YbS>8Z\D0(;VSOeZ;^JD?3KF0E1UDRNFeO
(,JNB0:,:_PFO^_<V6IIY6\F(C2bK0RYf+23>f>^Q7=;4W#V\I);SDI_(9&>+5TN
68R3=eRQXd,a[DX@1Z4@@JfYDT_:Jc^UI1@B[LGd/C^2O[,M4IKNC,ZIX<XF.:f7
NA/3]#(I=a@39Q4G];gT+3).R3KQeeMY>YXXI)@Cc^/HZZ#e]+>?2-Qa<D._FWd7
PG8g)5YI33;=(2)AJC[WdMbK9^<\gTg4V_[fA##(bf[eJcM)(@V+LO1P#g(.-=7;
F9)9TRKOd^7E-Yg89::,UTEJ#-(.8O:9S=7#Z;QD_?CcBENR4CeZZO,SPf#e8JU4
5c3#_Q1^=+N1JcH1L&SXAMba.(bW=),5-R:J\IZ3JTf:#3U4-#8808[GeOF4(>dQ
F.,5NY1\?eVGZ>;FEPREU;FZ&X=gV.V)IMcfE0)&C>IL>W>OY09Q(6^W.S>d3B@;
(3+P]I/Rb=ETK7AFVH8:SEaGUOF_cV&G@a?02YD],g_J&71)L:48SK69UN2QDbaH
V@X8]->#]JVCFE[8b#.Q2dd/,,ce)/>@(GDA(g-&@1:F(&>1=/UD5P)2=,GeX([A
9\>SW(LEOEEF=gN/d;\d?8H\G?330#T7F,X8FJA;#EbBDR#4(TZbND7MF5[DE5gf
7gfM]7BQ9&JJB4,#OU@c.25gX&66(Z+5Pc5]Ea+5F]OY2-XD))@MU0S>.S(>#3]6
J]_KV@16OIO>TDPU7a1+\JH-MDZC5O:DfdKZ:9f#2W4[5D0E^ZG0;]B>Z^C<FBIP
O-e03We&5;[>LbS1BK41H)JM^<+PbCLQ#+DC);FYUC822e.b4/H5DV1O?2I86VG7
:)I5Z=T6T9AR1</[]5H5>^d:[f+_K\HA(Paa1)7^XLRQ/?ED<GQbS8fS\Ng\?BSN
R7ZFQ35H0ZK3IX?OUE9Zdda_R-2[Y@e;bR>W6:OM0:fC1?ZSL_J?_\eK:;?.8<)(
+]aS_/4P+<S<YN+FBFN;fSQc,\:a;dA(cYg4_<F5XY@^7+YL2ZTOK+D]7\EbZ7\e
M:I,5:@^de2I,VA)Z=IM].=9AE).L_U87_>-.eLXfEE5YXXR@]UF7ENaL-5@:^H1
V54KKK@Ga7]/<J\1b\dXHBIUZN8JW#I.N9,O&-U=?K+&[>^_QS+Y)(MaBJBLYGX,
eITM@CfXfbP6bbd4O?E(,0#)^S7RCGO.GP,SU\?g_4b+dUd:&LQ)IO4.F-J>c--,
WggcZ3]1&]YD1f)#Z9egE76.\1g&@V/:G7X[1\I]-^X[c+8aHC),cdA&0TR^6E&3
5(gQ?;@\3R\LH[b0=IU.J_U@1B9,RA[@BOgbA))g==C4NL_TLIcbJ7^2I<ge_SdX
a@C,QNW;X=QD6@cE<;R/91Ba<+Rf.9EUJ8W&VfF^9KTM=7F>S]VFIO7@,Q1gH[Q+
e)&--,?>JV,)OZbZL8M:V3:^YD<gFAd2JLgW>;\FF2W?NYBc#IN:6aF8>&DS>SVQ
0-?g5JEO(Q#Wf4814Y=Z1MBIN7#I+F5fTN,a,#:@6YE_^-cD9NMDfS&O,[U4-1fH
A\IM18X#gCgfbXOD2KE?6&9ff8_Z>XU=[4=4445H7]@LW0D#)F&O/bd^#/16AQJ2
-4F97.0X6PF)937/^16N&NMXb-fc\^4J/:gXKG:O1YF[R14R\T299FG5D3>QZ[:)
\339aDX_[Rg5U4gZa14:)>#GEC=U/(57R[3KH#PH.70CM\0V1]C6(,)[RDgOB?7;
N0ReD2EOB[K_(C&Q?O]A_OF]C]OP#:#ZRI,,8#4bE,;a#U1g(CBK^b_1D6/,e\XU
[)&#0E9CTW=HGBQS[Q6(eMUR(EXCLX?2S,,Q?/DWQE@74T1<HF2G)d&I.f0=);L;
3A,12Z2KCG+ER5UB@O^YZYTN+Of+KC.+3adC-N,=9)Y4X\<L0]C7&GMB4@WP2&,6
L6Q<Na=?TKIKF2,</@:>48D:><?S_7\bAJC^OO>H2U?/:<3a5)Cd)Q/.WH4]V[F)
09C?fT[G52^f:]?P_O50IF1:#?N;<,RIMMRbd/D:A8dF@W531<6_gF-^,IYKa.N6
Z+8N&&:c[1b^+I_EKdKZ>f)&XUc+A2c&:4]1-MI#&5S)JJH>_CB8c\8DA0:ZOcB.
Q6;MH[\P\9MR?Ofa7V3[TNgcdG4WA/&@2K71+S[N5gd;G[0P(95J795:K\_WDUC(
\2I-(D&^A7Z9IH3<^PSAP96_/E@M\\6a#]+:/?3?;Ye1-+)U_67]f;B^?C?cXQF[
QLS;2Q]U5=.fK>/PL=1)3DC(/b?,B4SObcT:aEbT/(dA/U+79UV8gJfMDdIF..OX
9Q/SCd0?R]d5OS:0G@OO&-0.HPcGcYIbH:b3TdK+c0c5ST.8eO-b_:9a:\WPRe80
MODe096<)0P>02H:/ZT#2+E-9.eRTeD,E6BTUb5V5;8eU;X^PKJ>GFT4Q5Ug:fYS
;/<ScP]@,gce.N<=gAAP4B8/0H::C]90&)LOMD^V@c)AMJOVY@^]6LJ,/f,A;]8-
8;70^IPD003@cJeHa1CY6WLBJ.YO99)3<>6aY_(]ZU)]W(c64da7J&?49]A<#_DH
JRe8#EQ5(ZB6PAS9475#_P6>N4<J6]H>8EJ@d_,=&NHT,#5JH6\]?-aO#FKVKZ>7
R8cY1+>c8L(WXX3>TV\HT4IZ08)REOXSLL4#IOL50c/7aL?c0YfB37@HC>KS1,4+
ETE,H&@F=,UZdMbAG2aZb&4gAC#,@,7/IVZfeHC#G;5DQ33[F>eWF8QfU6MBD6O^
ScCOL[MVYY^gO_R,UZ\f4:+AHYEE(AC1L;4?/c4GTgS016327-NT9VT-WU-cA+)W
R^;,<QG\@=3Q_gaHOd>M6;?dB,S2.4D?K#J.?.^I;#X4HbM^G1OVHH8FA_Gf=<E-
HJK19XRD)VGe3QB[gL,Nb+K,)5W/@^BbPe_A\QJa0@F?G8^/G1bB>L</L0LaLUdb
C,PL#7OF/V9=Wc>FP?-.MPG;Y36b/IS8(aGK8EV0K#NYZ>6WC+[]1:_gEAMb,.>H
@?O6Z^RR(,B]W&@3VMCX<YP^A/.\RO_VA5--d;)<82M:ZC7XSUeb137c?2H9+0W7
_;M)Uf[:LbAELcYWCHFERT;^d;<2XHQ^OSTbC/),G7+#^gI2-@/Y=\)AAgc?Y,6c
>c3QI_?\\EQK;3GTb87@[X1(a:#F@:U?Y^1L&LP90P=#bcRSA-;OE#@YZ]=gCW;e
QBUeJa,@QR8Ze=f@08SR6NND;+FX[OBfJNGOGRe_f9)PIFHG4eJ]ZVaB?dL7J;Re
+&b2.F9cWLM0K<DX=59:04d28C[\XA.W+&]A#N8F,#Fb5f.E6SD6@;];5RfB][HL
DUa44J>H\3Ob:M;N,fM1&M,>@E4CZe8W./0d>@Cfc[ZV?S8Ab\C9<\#9/.E9<&a?
Q[\-WC3R8[:1XD[WJB<U:>KVX)OaCHFa=bL\;^Mac87:4WX[U&+/S+E]MTKbUFH5
\Rb)=.YSU?^7RAQTU,PI6+A.5A.VS]_>64F[NPE:?/eKP3N6A9TOKg.YE5<6/6eU
NIN0JTKDb]:J(HU/f5^Y4+>.\9\]E0@(A)?D\MUFRN)cM80UfIRGZ\Q&L\40]a-@
P7-,\D\GJ#gQMa)W8D)/2)VM>]g=_IY;](E.07KR;NU+);&I7-HWWW7XP5>a;:\K
K.aF)HK@GN:dcVZKZO)TQE#B<D3=CIF)791J6@bEbe1;ab=(,COUCD+;1J9:+B[N
8Z53OJ54@K-TEd,0?3aeQS)U4\gCO:><JKH;/XWg(Uf]780F4HDYD&FECA,/=<D5
X&?Ec&T9,_H>>G\(:;QTK.Y(7P&H,1Qb+9MEd_-Hd\QGOfF-A:AbFZ_(1)LKg_51
)bVKe<QS:PcK^GaZg5fR8.>KYL24?L(EG_GAFMc-L_NbeKYP/MRCC&=^@=(VQ@8Y
Cfc&9KIO=-FCYaKB\R3-5<QK@GTV5ggG/RO4A0]Zc]Gb=,<@SQE.+9>P-A&:G>61
Xb+0/V-ZbK>YUC8-D_+(>PB,#fcJ:Ee>L7>Hg9HG-)1L)BR>0X6\b)XING:;2W-2
+6?MC.#FCEdP>IE5K+g:19M]ERO[?T?2SdW,Xg[d,:?O+eYD41J:#?.&O/TU8?#:
]#C(1\TI9@3>bHb2aY-9ca424B5#[]dG,WDYIB1T\I+O25)Ee+,6,S=K\FH]+2T#
+H+^&]A(2<d1<QJ\N3Z?#S@G1T<?;agH552+M3M8ZB^LQSP=Y:]?E(<bFdW,Xb7Y
J>M1gKMJ1\WBY>W1MV;@g1W+PXTA(&N@b2ALe@9O7)9^_&Q&=fg6J(XI:O?]8]T=
faGe,dD(K5<C4NF;E/+:D8Ba--Q64;FD-Z()>90_L15I<3WCC[JEF;d;MLS9fE:T
PE4YX8JQ]QEUL9-FdfLR-6g4<NUWH:3ULFXMMPSaaV=E]g<]c]X+U[(Y+^<CfL_E
:OAVL\1I?_;8IIHE97:8)dE<JOWQZH8D_/LXANf/IBV8>+0OX)K+aY@M8]J^E_PA
]<C(:;XX7dST-IaGdC,/b6.PGP+VeAY\TNZH^1ASIKO:=[>f3.A/2OZ71)(7ed2N
MbWWd(#d<K)\cOa(@1[0.TT3&43a\F9XINc<L<AHN\gYBFgXAW^dIJZbO:&5bY5e
]:#?MOI>QB+@J7^5N\L,0W[O81X<Tf0.V148>MY_YL&GKJ>EWER.b#[,I/=D>U@F
bBQgE1RTQRC8<VTYW,8WgB(7TQJ12<FTKGg,L?8PFcd_5LY]IaM5B09(^N99T&EF
LF4\_8I?D97)TRAHOQ3.Z_#RB?&d45aU&8HAbbF>=?E6<C,YLgK6OFU,<cTQ:2?E
8J<<8RTcHP>H@>SEZP-53ZCAM?4\FY]7#]SGT.OZ9RCB-+(-RC3\4EQbWAG1B#OQ
ON&E[^8^E7[.XO5/3VC/QO=_0ad]TVL(f7GadYU@^KUYf-7e\(52/P8=&21C/(\K
QZP_6_#gCMWf6_=QE.[)3&&TVCG8a(+#Q4ZZ_UaH(&dBWE00;V=OS]S[@V-3?Q9:
ATY^+8ON)eW+9?P?OBX.<+9K6bJF,T,6FcDaB7#(4IFQ7I+U.^Lg))=696#WL?@L
?I+Xd(R,8KYM.TE@3IReI3A0GddW:EaQ4DW78D)/dGc,6HCX>P4ddfIS5O]G@QR+
_E?Y82AYNC)\&FNTNF9c]0K-<@P+1E&I(QEGEB1L#+99VWND<CU_:>X7.A+&II<g
H^3^4ZbMFUFIO0bV84:<DNOfdY4F,7d/<E>]X2A@Y]3f#^^>:E^I(Ea42J+#0<V^
c@J=bB)91RRDUA=(738L.W7N]W62U20N9&7OUDQ85&]#_;8bU=NY@bIUc9GfBe?T
KNddW\O/Q?L.aC_O3C=,XR?D#f+BO@a01g()B#RL:NWO,R?]P+-P,3_RE?Af<:Zd
T@3fH2?#HK1TM@PaWNJZ@^Le=<&\E^J3ZPd(@@Q=/g;J;Wf0I88)N0C.We,#;TH<
cYM@V]eeXfW/12QQV8g(G>[9aDM&R.]4?,Q5=GSOeWg1aH.cfE\N;Qf&,&a\gU=8
]:ZDRJ^ZT1?S>TbH3:?eBg)L42P(E0&,=UBY0e\JUX/L[>[H1EGNALc4YW#fIQ1c
Fc<6.Z,a^#fJb5,ZbGAL39@d+LYGX>-&,X2:TH\.dRHg2EcUD#F,8a+??=N&LH)f
AD:-\-a\Z?Z]d2AC:>HFEAGCWC>cU<a_GO3#.P(.c^;b+#XbUAcM+gYd+#H8fbOA
UBW.-N;LcHbZ(MQcU(?5ME[V:A[@dPdL63C9ObE3>[]7eD\NU<6RM=<N8A]>.24V
4&;-dY@F[RU^@^>18L;+_T;_M[4\gb1Q,J<T8HGBf4W8M#N8;?K8;;]GdAGNJK;Z
:;V6Bf7]6bg^(9&9aALfbST>f#?ecXPN/]&TGTP@TQ\90Y2(D))_^@\/T&(P-:7E
5#.^1H0Aff&O?AS+NUR)D;9OLSef.)L0DgA[/BB_[@628&-\;O;1CI-F;BBf=X2C
HYW>D#)(_3AGY,U)S]WASXN/[S+J5eLZ6Uc79\T[.(PeE_LP<(+PRY67B12.O+:W
=?eC[6;0N(d;TB8g,AVJ0/-PQ#9:4&>\fQd^<8PB\\M[YWRQEQ;I#d;1XT8S]BHX
,\)XMXN=#=HGDIN58>[Y++,+.^H-?YK=N2([F]A:7W7:>2+T]C-6&TVE)gM]4A6<
FdM_Y6H98I8B4J8X=(=b8?g.ANgb-3#2-.^:S+=\A_06PT(;,_7QVRD2Q_D92.VT
(\:(<<ATPTfbbP_=9=d=gUfMfBB<bZ9;,aJ._^,#6BY?XHGf3fVX]:W;7f]@&&/)
\+F5_.#(6#M,]W;ZCBH=J466DD<dDW(GLZY\/)g@XE#72Z<_[DD1K.J9?]:Ze(V-
)FCWVGf2.OI8&MSg5aR5]eC)K=3A(a.A-UfJIF+cIg-:+dd,7fCg).[VJEG3BK2d
@dA4_B#Q3;E)R;E-=3d9/38,^,F8;a<:g<J0-2-gc<+9=N:HS??-/Y[A@3LTYC(8
3T/A-Md.C@&f^U(@#Q]UW@&@@0eDI.B:#\e3c\7Y[?@7]6TN,TMERC>8Qf@3:SdV
LL3\WE;/Y8,T=A^Lcf\O<>Y7/d152+L@.Hc7OTb6ST<K^?O<(76Ka980Hg_ZA5g9
\e(LWXV/e\B-&e,ad/\4g3@e4A1OU6KDM0>I94S;33OFEc@#P5eO:VL=N04B\#?_
.e+K]:QVbU]__(W\F(fXF8I&cNRE\4e9\0O#/J=?bY@92eTA/.A2@O/9<U8;:L_b
1VB_8\3.Z5^1(4G52UPdTc_R-\aGE?Ja\a+g38L&)51T:>7U]Pd1cDMT:P[:_(,N
4IHN=)--RMc(VR)Y-a;U=HN)<+KRQSQcA#d=(JRXc79-K:JC<BK]#RS+Tg@RK6R#
:Ld-7SJNZ&0:#T3Ha?[+MI_.F?@N3aG]WV83.Jb_MM86#JC[Qa_&37Ee\+cDed^,
Bb)F&?CUAb4)Uf)>)O5_]57BP6,OW3=C5]F<e3KMV:FKgL.3RBN&X:&6-)dB[:1g
IY;5;D@Q[ZCcUJaO+[QQCZR/:?Ib>L(\J2P_]b88TAO<g[\Y&g7DQTPECfF);71?
&\,L4;/]/#VR10L3L[<:ETT5g=QM5(#D_4>\Y4P8U>PI^W_=L/P4_X3eJbF04)/e
QBB-(AA;f37+N3>eLdCHYcaAbTfKObYNG8IaT5gaKPVHQ[HOJ>4e67Q^7f?(9,>V
PQQX87BMO>>;JJH&E-L>11F&^Z^8eOGQgJ9PG)e+0R]QBXAR;5N.]2e0,:=b,1C,
.3d-J)ID#5\bAf[CTD..8\#.G/6[X/_@?D+1WXcLRKG-g[CaL5;Q_U+.>(;E(/O6
???;OIQ(ZB:GfP^[CW(#MUE:6a@V)+8#1]NfB#BJKB_1.?KREFP.eTN2Z)6AZ3X-
EY/+IA4\-@-1\SI&[.(7T[]^MWgB94a4;^fc-S7RMD#Ga5Dc9(SQIb9_;bZ,M]>]
7M2SNHHO8E4#DLKDgf@::S(/9d1cc4+9GH:XY6?\]VeZ)^/#>[WaY^/H#-V8Z/fV
N16F&fU@J9P;^;(8fg<^[&&@g^CVd2Yf(@23WGDHY(Q7L,0W8fS46:P.0MV)49IE
M]WIU7/.#XB/Q4F,4J>E8N[3M=WYg)]^/#_c5^8f8a26OFGSBHR8DN6T:Y#<aI0,
ELY@I101C0Y<cGG7FXC/RQD94b@L)W4?)WQ/f79_b?_Eg?J<ALcUP1Z+2NX7HV:D
8OWFc_DQ,IS&Y7YYX2>EW_Qaf;G-g;>e@SQ@F(BX[H(b;XH:Fa61O8Y=E)R61#L_
(U(8+UZM/.U6;1SfOHS-18>,2Z>-Sb:XQf&1MX/:N<[T/7;9gbQS2,cb20CRB6^=
CTG<47<+d&NWIJJ/8V2Q[RH24XL?bf<SP]b<(c\PPTR;Zd)fGWGd977:)Q9VX+]7
cLaAB\=]]S6S-_R.3)MK3_9)\F&bb;U@P=\Q7,AAf;f>Kb+HZ)[R3-SBL?8W0;YW
B7,R=990)_D?ADPT(34cY/Y>TbD7&Ea]3^REbT;F4a:)WP>:O[_E5O4gb;^9(488
@,07,)6S=ee[S7G)3LVV[BS/6N/Wf6B@R2b8)+&+BLCNH+8N&SS\f:+(=KK/0E<I
4Cf<c^;,28f8R\<>&S);>OOEHYgE)&#,Q_\H9;#C_c>,ZH)f:@#e6SFceI<5D9A)
RKS#-/.cD6G9L3,abH-AV9VX,^]ZV5V2/+?EY2>)YgLY1e.(YK3S^P?WYC_LU-M5
5d=K2-[NTUS>Q,5Q+IJP,8De67GKZO.R4;03eC^7PXMLcA&HQSc7dLGKKR::ATHU
J./IR)A\O^70Y=G@=cZ-bY&USEL-_1[Y11DDN5+CT_+DW-MU1gJgEUfc2IRH?A>L
.(ZU1YL-;,GfMN&XVd1>7aS>T(#E#\Ag(0NPbWg?@4,(-4Zg9=Y=4@#E<c=[Xc#>
FBQ+KKf&-POA#0C0AT@?b-1#A^/eQ&YH8e)/>f]-[:dVA6/d3-fQY#]BaK,GVH@_
R(cc,Mg:RQ:bJRO-b<aM_)080LRF_AFMA?P&9(8HZVZZW8RLeF#>K-=.Y7[8(@Q\
A-OL2bgff?IYPB[.H?OK#3D&4;4)P6D=?W-[.^=2S(L9;=/]T[f99WW,.<LIDTTY
<gX(YBQ@G(F;1_.f@gd.ECcMR)BSgeYg2bVK77?=-K\RdKI==--g:cCZ0J6e_2ed
,DA^R)_aGfD>/<fBD#.P.S^acVF(WLQ_FNf0G<@Lcca,XQXB=3+SBa/_,EU?C8>5
A\e=8O6XM>L^c<;4T<&@N2O-WSB\3@#Rf1Fe[.BS-X:?@8O7Y]2gX=.=XcN;f(KP
8K(N_OfA.B<=(>f,+10Y1(X\J.A@g_/BUF1&4VdRWD+X)DR_>KLTMagS?J]aX]ZH
[&=VO0\c9S7)7b,)BE,SXF.EODC<]S=4<]U:/[[CW[dD&HU0KN^Z^4;F9Y.W.ZA5
-3BFabASN[55>OMN/6;R@AGZHIN8fDW5]P@^N;OYSHa77^QSeYVK=B>D<5KKVd2>
2QCHI<M7&N2K]Y@W6,4FfLU,B2aE5).9J,.WN3b4=3]6NbM/[9O-HCGJfEELAT4?
Z;2+IcD[>N[/;O.=MQJdXTV<N8][5b)-cKN&@P>HPVC+U4S:)3#ZGYF^<?(=GI2d
,\-3-d,@0<)NSLM7NZga;M?24eBQ5(9b(4YIGb#IYP<Idd,=EQeY6O6T7NWTXd==
EKP2TS+5_0<6&QI>6.[4J6cO/L8\#<6XO1NIFLYW0A/Z_AFZK&9TV?>Y+f+S<+aE
0-N(EYV_:&]9>Ld#8P<XRJ;K1cDTRg6Y.))6NOSB?P:@&6E.1EGbP+N#7HY[I^Z;
?@F&8=(+6NeeVNeBZfB-DUHLQMUC,B,MQI43O0^[EPCBHFO\#P/KYHc:I<<B40SY
BWQ9JbE&NUHGQJ,#^G+1/07;P.HTLd>,\V]\e8Q3c3aKEMNK1KYK-ZNe]T)U?&AQ
.d2Eg9YOSW.WfI:)-PbO?;HABgEMDC]QK5PNd(94(Kba422(\e-.0P8e;YfO?FD9
W2^FW91aF1L=^2KgGE[>D?/)^;/.E>IE+,PYa>1P0?UT1#2HRMN:b96/b9bI0<E>
EaNSR=Wbc:-Yg]OF9[be[_@VYN?[1KIYc^_^9W:&P,-dRFf,\0U(CG;+^=;Je436
^PLYg2Fa<:9)GQ&Z_6GJX3-Y/M[g(V&g(.MZ]&U.b@7N(FUcA..Y)?0EL@c\[#M)
Y(b.FP/P:b]gAR]9UJ3]6Lb[2JF&b9^;E6FRCZ_+E]c_d(&J,^6WaTbbdWP1NYdC
bc1a^PYfL[K6]-5D#OGI(]]SO]5OG_/?BK8M6bRJC2D.b>)8GL)7V^H\8Bb5>6_[
^fMDE@eA+B=8K#W6::P_09Tfb?W@)TH=#]3IHCWTO;I^1HE(^U>JEBQ]V;c:OI@)
BK_>g38^IUQZCRa197QXC9^/5J]@I&?.#PM&7BbIC[JAMZGddgA72)(Bg)W\5T5I
T&C1OGJ.X#TA6]DWO>Y17K/A4-[,Ha:2dg:Y5?P(<EN_<dUFMK3E8CY><RVE\5C1
:E1K@4Ma[K0?HK,f.6ZLTQ\+9?Z,cG>_c@TIcC:LKf1b[eV&0IE\ec=7b#R&T[,_
L)C(B3BFe6MS+]4Rb3+OW>4/464_eW,#6(HO4?+69dKdBf0N-NF1WXf-C8CZ+Ia#
7T(cNC-.A#?TM\MKdaK)ZKJN,3/9K\?2R,?[:BbY-\>(AA+0U=6.6&VSLFFN<T)?
8?H)19@_Qe:Q6\Dg:4TMC(..(9C[E+K./QO?:UAMe2:YJ-<9+75+]G8c9&#.>HLb
JR>a@P&c#ag=S9:38HR,&#W8]LL,B]_G)(VM6#ZaDGQ/D&KH4g)+CE(FEA;Rc@>Z
1@b^A_a7Y5(=_5cC=g[:/M)]WW:<(1-UDAa=-B2([gP9D5E6GZB:(#<-aQdMeGXF
\MGU9A0--\87BN_#/_[X4cP;W?:/Z-:5I-A+25fTg]&3Rd7VIDffb9c)@F92CdZP
CSRN5#HU42+WQBM6/<9D0dR\0-bQBaa[I3X]5L.CP>1.V6DNgf0X,5a62.6,BRXd
A9P?W0b#8e_Q>5aY^OacNVR]).FMg<QB5O]4JK(@4J,A@:T[BI_OJ[IIdW[#FfF-
DN&(+AF[M+0TFKcJCSY,IYO<AZ]KVb/aEgcU9[6L?\;L:1Q+\Wd+S-F6DH[A(=V/
C>OXFNNeB>[DZBSdg-9eEa@Cf]XP_EMP6M^\eG#ScNf<KW3>O3@^0)5g(IL8ef@J
8MfFDg?SJ7c1<RA+F0Dd#C)8Z<;LV=FMK;)EN.)-(HZ_c)@,H:&O5UReN.VM.QSB
.Y_.:fQU\@8,<aTV,;4bAKY2V/J&D;7LY<AY#]8QcO+ZL;)EPeJ_b>#6acd[8GMT
-L8C,@0d:X)Y9Y9_W&7;^b:F:3#L:>45FG+1C.10bGT;S9fVd5AF,NZ=5_dI8=Je
_T10F1,MTH?4E>N/.95:F5XVSHJ),.>.D7Ob2;f3Y_OcNTe49XS?(O^EJ29HT6=N
Y)Dbg9D:>>AA,8>UE3S[]F5+K)R_E_FBFK?dAgUQ01-<c\Q,>>F3PS.8>O]J)Vf-
Y9=_XUcPG,MFQE@#=+f1C9M,eV&U[S+0Z;#3=U7\291HgeQ.M]YJ443:^8g@_HJL
K,X/OC<=S0-cTI>5?9&[&\-,0Ya6Q+6/&57g?:/\TXeSgBc<9D>MBT#cV.4YSd)c
BW)\6^dUG/<564Z5;.gZSfPISU:)4)?)fRcQJ#dQSNC)W.L(IDI1@-f:OCVD-XFQ
dT^\-KHNgFW9B_8?5SAC10T;_RVU\?+S<;=V8W^Q+Q)V0;Q;SDGC]H#C>QcGA8XR
M#OL,D[HD9@TeffZOAYg&(Qac-eUXUf@7X7a8Ed9eec/(ZP@+D&SXPK[3Y#SN:_#
:P7>V,FgdZ_WN,5I-O3_GO+ZNJPg-B]&f[T;@,6Qe4+=]09V5H4MEJUJJTVPHOZ9
-C_)/V^Q:6ASOFd=.]1=Y?a(@QIgcV[)0#aHI>g1/Tbe0Z]&4cAc+g7c&41CE2IK
8)=gDI4<OZ)I?eW1^eaKWSM=8<fE;7EL.C,W@b5_/Ie5]^,YE7]F46U/RXReT@S/
^X@TcCJdVS\QUF@N\\:?OFd0[-c=6NEH<V8^+[P@8H#g=UF2MC.RIYA\cKYfbCJf
Z&f.>07Q].JDG3[<XcR>fP\IfP9#_M+W<911=?MNGWC;Q)L,SH3JKe.@:<=F,J)B
4O],\5cbEaL]&bKR+c@D@N,Q]dPG#90XeCJ8L1Z-Dc57eT6</NML.9JQH1M4C/=S
26(,;CX9R?(Z7HWe2:/-\5MCT)eU#TaAb38-TFa()T:6P?>XAb)^DGb=<ZVOGJBO
INZ6A#4ePb+<O?X)[T;A3N>WU2K^8I?3J:3^JW(<AV?V-]XLV?2,<=(G0#KJQQYD
>S2a>d6_Sc@2eJa>-g=VJb9(NFO<ZIFP>eJ4aCR==NXI)6cMF+aFg<7:2<(,._F\
JXR7^Qdg;44gdL-/gLN1XZLbSOPDTF^F?K?WT6DTYTTeBG1FT,TY^FONHUdf=XZ9
.?I1RW_9N=NV;]fa.Y55_^ccXBb0aL,BSMYB@HNWS:B&/17;?d_4+@bCPS8>P)Q&
U6@S(ZKSX(]WKE#E?J4_>BV13:b]c&V+H]F=(+A&X<LE,KD.e03cMX&29V4KXA(7
gPZ3CcGJ.2JXEfgKJKMB)+4[e9?P_aR4:9a0E>8C\@P12#?<d9^bR7[EKIe&_#D@
:\P(dHFd[A[3NN7XV7,)_4^PM,XcI]DAggGL6]d,f,2F48@D.IUdDO\Yd_)EQL:+
8&]F1\:<QHDE\H[2b5UPCVN40V/WH1LT0FISEQI1XL/.0a0RN(Z@WDgQbfcF(Kf=
U0EG+]&HHaUT/S76bL3gR]X8H?5L_0UNO:g9+HEcJ?T+>g-+A<<&?3#,F-H[JCAO
S:I3dYS6=<QaN/_]fcIJUCIgEf&7f?_E.2LT^KCbE?C4K+3K#;FCR<9G++FZ=,MK
OGfUPcaZ2=EMAEA9KdW8SDDSb1TVb,XNA[F8=<G_[7e&B:2+/.#]Q(D[(K6ECAI^
+I&<VG&/067A;EAb:Q_,K-XO.V@F/d:IRe9Jc6Z&Q,.TWL15G(&OJR?ER\2,R\.E
d0U+OA0)M\9TM5A&._^V]GeOF]=LZ@83:[NGA]+#O854bXVaa:@#cS5Y0AKWA=9-
aY^<)>+RO_@:(d0OM:#JIb-9_;?GDC25[C&B1ZR@KDUTR<Jb3<Na5a_+&RX:4ZW5
0:B.&[V5V#0D-aY][9&#++4&\cE7(290#NL;67[<=KY./G3g=62F<\#7,FN7bf=F
)203N#edYD,b@2,g7]=d,]84;#YW9-40OL;Ef^></8(QY7G^\+K#AA(^]_MD/^Tc
_B^JJ4GW4UL]J(^?f4WSZO&GaU9KL?+Z>C/F-ZJg6IFcA(242K;73gMNI==^AP5N
M2Z5C-^COeEeZ?]V+UbcOU:<)@g\/C:YgIf::U7dI<GM/b:KH<1-H-25@&;6fHCQ
[?3=2[NKS(CKC(WUKa05:+L#<Q6.?,/]VMf5<O,@]d>)5d\3:];@8;PED5:=CFV1
)E.REW7W3g\6?,g_Y]XWX=[bP4Pd(f5P?Yf+DI&[:@UPbH--<HUFDdX]&UZa^[gJ
T,+SL@beaLRROgc;)\&X<Ge<.G;)0Q9MQ^=74;Q:B7]Q#032W]gF\4g,M&5@XU](
K2\f7^D_=EI-5_LY8T0K9EKRE7e^c?E2<&bLdPU;bY05D2&cc>2Q5]6&/Q,B+QS2
YaRLZ&bLAK.4H1OD;#WJ0Yc.dOf5D+\AZ3;f:/3Z@WF3LE_QC(24;BRCc5Ed9f<a
g)(@.6@+H^8.@a/c/Q(8<M88FR5-cW5T+\Pc#]Y#HV9/(MADGA+.([E>#M=2\R<W
/D468]g@=:PQKT3H@f3aP3cRcI1/2K-Y#:IA8N1gE)V_E&a1OR.Q1?FV/a<(N2G7
B&NAVC25cE^UMg9JL-HT#9HYB7E@<1K+Z&C,c.[AZ_a]T_5bcKeA^=U,e5[gdL-N
eR#WRHFXA>=8F,)Ic.W(a^D2X2/EISK+;EdT=?[E?M4MD?D^3;NYe5ND/?J\/f2?
bP():62)g]c9g5V<UHXYWF_I_&9e3IeU-#ZdfXEU_I?R\WKQ<T_TRg0<7Mc\FbDa
\+85A_P;eF#&,UZ8?+fUP]2\##V=<S4TWaUe(Z4>7d2Z^.&5YcD(dEUXCK&/S&bB
=0@FSeGO1@KMR(UAI<Pd3\^M&\D#A[<g7YbYE8,:gbH,eeCfMU(MG9QJ]g5DSD_[
X=6VODeOCGg?.CAZ_@MJ.3+?8.F-[L<:^EdZAHSaV_>FB??(ca+e(,=6@H/M>=eg
)FQY<#(4560]][>ILc,I;L0CN^d3W,E2)\E_=Y]>+FSD@acGE2f\/^>/+V_5YWVb
7^L@JU\6&G2SYSISe:)X2:[U;<7Ueb,-)CdCC+RP_^W4:e._Q^7.;b;>[</agN?b
7e)3]C)R3\NF.fG#dDccTH+N/L#1dHSKK)cDgZ?:\BXa^/W0-#Z5QDA09.V]A=4b
+eBFMIO2(;HFO.O/e;[V>Wc?2KQgPJ_fW#>KUT/VT/a1;gS05@eA9S?OQUe8,[7a
BJ1<(,VES9g)Y>Qg]/GSDf8\TO;e,(C6OaGW?d55-?fD+\,,6Pb\DUca@E8Q,R5c
6/_gOGV9R0IZ_a+a0JY?#-aEb7Td\Y&1W_CKC1gT-4WSY@&6]c05B=MQLRZK_KK.
aT6/M-WYD.1SXeU=0O4&J6&;H8a0B>#BcaT+\)dGPO(11dgH]2cDW#cE#6:/E\^<
e9YPMBOT90U>V3M;IXdee,/]44K)9e&KW:JWQE;MZA><,Z&-G4[-\dMaScN1S?\S
2He-.5aMaO,M=CeB2/Y>F.TYVR4L>W>94D8S+W#2-@<5eCGe:e5PH+(L,^:]Cg6.
.b\1H1@[J&AVg#K.J]fY=NcMY2;I;)K]=4VF;@+C61@N=L#YUcP\\=?_6/0[Lf+c
C)X<22Dg-e+CAa1L.B#OWYgH/SPG3S(F?g#O+7Q)]E2\J6DL,,11^^dg:&@X<9/C
X/=S5YNe=g;OJIYAPd-Y4\-bH2X-])(^QdD^cV7Q)B4f&d<9K;=4(Q?7]JcWBLGA
AAW1YD8=-fR9<>c>=7Q/Ca@67bQ6V691W?a>ef8W&+??:dUfedSZ1GJ?d4HNVRfe
^0\C9P9TNYgMA8?3J_1(aZD(JS,1-6=]LH@(4G)6Cb)@S191-G]cJ6QB>JA-4YAU
#g&A/5-JGg9>^YV.R4SAE)3X8]H6McML+/4S#:F0+IB1_Y>GS,8TI&[&<AfGVg2d
5\HX0gL5[&_?=A7abDW)aW[-;/F&?4bUWM5AK5]a\RH,TO7<P3.NFX>H^\D5<L0N
B,9C)OGS\0Aac@HRHICLf:Yc,6RQ&_X>2T@X=\OC-\Q9bKf/I]K]IHIE+<LA12)[
bYLYL3@VYF(5f3_1PW=J07FcaJT4f7=LCD#O(E\4dP&(O9STTX8K/ZG^bg>ZD08(
aKO=N;dW]#WbGI5>T?7T)<.fD4^CDR#9DMT>)\\]/FRf2H>/LW2H/X4PQCeR(T#E
e-H7b#,?A,g^^=H^XMb#YEYQMUG4^,]PM[DQ0>6SQE91_&J79MN6:Fg(,]cfLcX(
\C/\/>K>?9_2dK&U6<^Q/T;1g,_>3@;+<S&e7A5^@J/QO0L7-K9;Q#[H=_6f602B
7&FJR_6S)ZgX5[[X)g9-QXNF^^7]3?B1LbUAI,BBL(3=Of@8cd[K7(?Eb#f)MC:a
Z:B&0VM@@B<-UeSEPS[1O=;XAK=4S5cWV[-\-+ef]]IYTC,AObT@=M(gACTU[2=W
,)9ec6_7H__P_,@:X:YZcFIIXLGGeEG#)Y4IM/FXd?<L3BR=G>)bJP,UNeS18KKX
_@f>^Gf-PDf=bJ&00_;,TCN5YO&1XP[fB\2,(J;;VRN;SE5Ed:P8P<EM=g:)83-U
\_;VLWc[PX@3d3)D_&-J[4:R5YW<]0g>H)f7g2Z&_EXFN(P0.+UH+>Y-Kb&9Y2L_
B,b9g,MA4^0E9(4?__?V(g2>0Q)cDN([3_+8=cGdVCB0K&)Q/4R4T5?aaH2bY^.R
T_/@I]a3R\0b-f]A3K_DY=9J7]QdIRJcW^;KP]WbcJabGEMQb6#8?.:-Ia=3E&:(
_S^R;6<-cB9-CJO81]MRa,c--Da1D#FCJ\S3/HEZg68]/-U.<7Q9>]:5O2TBW8L=
&,5K[6dWa/[&FFN4e[=)f;N.FT__b\4)966/JCAFAOJ=TV@65SI_(bfCa=X#WQ9M
77]#OLU&PY(4dg8@@^YRR[g3W?:T9H]\_3Z(R7P&;ZK[RH+=[6&/,VZRA?R_c1-0
8bCZd1GCeVHN(QK[)CHbB=eLc,DW1;,/gLQ&20N.;bET-[d^@(bd\=74C#W[b,[5
D[Y8WX+70SXUdTS;E:Y?\6+67#[5ZdK#YI_+B,gF#g;HMG],dXKDc\^XOg(-XE8V
423JfW4I#UZ(IbFbe?]7;]_9YULa>=2eOCIaMCbM)+1RY0,<1,..U11\WXabZO=6
/_&8_CMI2eQ515D]9Z?X<1\8\-<bDRG=HV.cYa22B1cBQD0HEE,b/1;[\[#R&Q8d
).?<.P4U=F@8OgDDYG<M@Zgb121@/fDB:U,<V[J#LXPJP,fX2FKC(b@=JM5]E9P=
F_f#8,&D]]3>7>a;I.N?033e/.\AZ@(ZQ2(P,AQ;LDga7:U1L?b9TPX7E]H,-76a
G&N0MTF6=VVZP3]0H6@M#E/IK#;dMfSFW\e0^c]c_Y2)S(g;:]2JE4AP[/K)6IRQ
WO=@HWJKHI63_MRO\/d7(ZBCNBCbV]YS00c5aJf@2#F];Q5WES#c#Kf@,.e2[)I=
aPH7F@>(F64(KN65<)8K9F;^^-I<IdAAY3;UaFB.d6F#bD(A.,^YIO@LA_8U4TTP
<@SJST#CV=cZ^4)^7#b5_Vf[2+/ga?9E+CL+d9J:.K82c:)=UPKF53f4R:CM.7N<
#1_7P6^PR,]E)K0eC?(<b8[4,Y2BfV)YIGK6;aQU3X\^IGL1K2HPJ[C<3(=0UI;N
e)JA+N0V>O-L5/<edg<g7<fJ[^PQf/Pfd[#g&;V=FeQKgG4/>GWgcXL4&.<L75;d
>ITP5,@Qa(.c9W42K0<7@F.^)+Z#;WO;PaH5fTVEKaCGNIbcPR?3&(d&(4+ddI\3
^P.AB4<5X+&8.Q<5J(aLagJ_CbaHA==]S0dAX(W[[,bff7&@aYP+\,f+4g4==2E0
YI^cS13@@QUAf[3PUgISA(OCbXZ3AX?YNF7(ABD@]]0[c5EX60P-V7K2[L@]ed&,
bI(QGK;@8O_fUB-=R[fWEb_K9.R#JY+=&/CPW>C\R^HRd?9J]6,>_?47:(f0^9W4
fD-/bE7fT.D+(?3fX7OS#M9G=)OX#2H:X#-D,\2H5(+fGW18#I?J@Ed0EIAJ?M&U
<7:/;GNQbf1GaG0]>9+S+We,J5^@@EBdC0ZBZ<3DB:K8W(3fLWd6eG43HD3RO8d-
ea,^<HS>E,QI1/_eZ^XaHI;I)@6K]:;\V?bFZ<+T4Yb2=((G4/.Z8G).VD<Z_]I#
XWYM:-ONO6FfbRH;WYJ&3;>&_&-(/Y-4X_6ceG>@GX^V65_O#TU;FZWC7<<CXAKD
&FF]b/:/fJZ2(1S_LTY6+5B@Z;NEOF&/c,#J)09USWNXdHPTFUF]Q-ZbZ/5I&\0C
/B/T))2Y;(9+4[-f2Q<LZcf#&=30U&ZHZ;7gN,/;Tg&MYAO3_J5/N&>a-,F9C/K@
\MaOK3fEQ:VKYG:#)_dOb3c?8fPO.+S50/ZQ<+-=SfV2/eQT[3cORd29c_(>C8cX
J;G7P;ZU8J>g2g=V;C,GG&VQUEOEADGK5CGF3.=CL^Jg0W-)WMeff&?V3CR@Q=8Y
GL9^c/V#<.G2RgLLU,D#Y8F&4FcR_ecN9Ua:L4WZBYa:a46TSbf^>f#>,O<4I0.R
6L,;))9Rg+TUPKC-MOJ(F8P.L:N,d.Nd1VJ.,V+CTJ]-AUg+aIO-:Ae,fWI8JRc9
<T?8acUBZ:02@@W<X-(e?<LQ?3\-2&UV)S8C;d./4M7<7U5Z)I8IEBZ1M[Vf?O9V
?-E5##R&98>0#S<QaFa:<;+EJdT][[eR&a:OdC7=U.^S[VFCdKMW;c24aYe/gQZ+
=77)<LCF=?:JT9LgJ9/P&QM[<BV=P;a^9<SAN88>0:@FNI5VfcfP\8E?8:MHf#Sc
[]WRcF?Ed.X11<b:AUY:/4:X\8cHEPZ.48?+UK2>O(C#CPUDeZ<89VFP5#Q>XYZc
[3C@FW>NTXO;<gV7=U_\@3=_>\JC6(E)Y[T-VB[3S9X(VIIg2.5fFY7C\c+XF7;9
?_I+&ALKSGH)g]]-e;g+)JeRa7(Q?eR2L7E;^b67XQ3N<DRT/?3GO#7Z(=(3/AU_
RgL?EgSDM(IUJIfBf-_H_8;?Cd#Y_Z4_OAgQ;A83-[/4.&GAf<#Z2L<IM1cX1?F6
R5S@TN&Xa<6)M)e=QKEZ,W_:^aH8V,KaPP#0[Jg:C>.S;)ecPNfSJ(]F1TCLBU,J
3IDBQg(B1ERSK>&1TAJ)e>Eg-IZ\TOV9cGOP&S54f[IZ8;/CX^XT?^V#3X:G\[f_
H/JF.>L7L[E,fQ#&@/aP,K-->7S5gX7)\b+JTWBHR+7_Y^[AW:F)^b>@9T>^^Q.=
IM&0<Kb1C_A:?e>KKKC^FV/OG\K=#>TTM_&<5&ZER1Y+GJ9W<1RF<<I:9?B_ZSAT
c,#g=&SL?)S_OfJ&c]#TOP+K3XQb<=VENZPP@12-adE<O8Ce621L)R>D<=DfQBa@
2,d_L5?SeE3C^VGeMcV<UD0c12P+.@(FQ\:)((KL3+Q)@M^)#W/GE&>MHFKU>3.9
_LRWD7=>=\YTAH9F/-<EFO\9N_&GbO2c)M\CS+GXS:?cCa6@ee4CUQ-\b3TVZcd2
ZNT>FIH6KQ\b(U)#OS]/bWOZ3Nb)d=<Ce?5PMP3T\C?T8GbU4?Nd]dK6fG@8@Tfb
H/4XXT)\6Y[0J\BX/F5\6?0_6SF2N(]ZEPCYf6e:1b\PX4R7TgD-DCcZZ/a2RV5B
,WWYb\58fN=<L[;ZZ-?Q?/6-E1)fdX[<[0+KYBLU717\K7aJ57?O<c-Wb#2G(f#T
fae33dS+&BP@/0AHS;Z\/VN-P^LVCWA.fQ[.;Od_[7\[T&>5d.Y#6@],A[0N?CKN
J##[JM28C_d8N/^X[,.;.9.4ee>)6IbZ:ARZQ^c),96-LGOY--6VIaO3b:.]d\;=
\O1\XX>:E4gXefV)_7b.4QeeXb3GTN,@,SK(0RQGFa6Fed]K)O=O3O?gUgWT-?4P
OHS)304&a)=S(MLD&Fc2eGRAMY9@B2ObCAeIKS/ZLUBGb8CLQ3IH29P2I0/Qg:)6
?G8@)Bc,</c;>>=b6c4VQ7Aag1H\Y5V,,6Qa:]##BW>+#V9gW:FdccI&7f==TJST
?LE)PYb3^/74&]C8=gWgg9(9e#ab9T^AJ1-K2.8C4]?\CTX0;&/c@(7;&NN98Sg8
Q1&21f/+/J93e3]dK=aJZKa,fL,)I@:]^>OTZ<Me6(9.,O:54E..X^+6;<)@<@A.
XYH/Vb/XWJ)Y3-A-L56,.9O.754NNe?<#Za6CgG8W,YM]#IFI8EEZ]:9GRGL_CaS
VYE_K+31>6e1N-0\Y[K=HC[D]23I+&(MGI?,]@?KE0Tff_IcLe8X#Q<c2C-=SBY[
2bIEOQ@\_>8][LbCGGN+E,;A1.UNRSLfBSH(N1AF^E=MT:^gg2LF>-7&C./:af(&
86?fc=RNO]HTHQPM#4VE&7<35gAMQ?c#:LPL16BF)aLBNa;X&dI<_cf/]0?8YZ4;
Z]W4(I\DTUQ,=/2FfCeG@=7A)S>M-WWFa/H::IQP^fGRH1\A#a2GRaZ+E68A7G?g
AQM1EfW+O)b@4)Z+\SL68:5I]TbJK#,6=C(DB14]H[?e,7Q-3GM&_+N(YGe2SWC:
0K-HM>6,VA08XQ;<P&DgPId8+]2L\<JYZ9f.gL:-c>d>;dg^DE6KY)6Le5PNGH^#
ZX(A9)I9(g[2[Le;[OeP+2:MQ/gfE^M7>:T\QVMbV)dA3MQ0?R;+3CXBC:3KORQ7
@_>P27-]@SV)@RV7KN,QO)R:eM1Kb;V36KR42^/c8FR_g7[f3EEVU[OHX2O8ELc\
XWH(9FN0QK_T(H4GCT1>+,EJ/7Gf>+fHZ0FM0WbGPc:1US9gAg3L8P,)a5H(fJQ+
dGP&gS,#AB7:7[eOW]2_a#V\Yf#&5(TCUPDJG@eJcG;QFXOZ_6&F>RV6H5_,I9P2
c,>R<M([@a<O#):d^3MC@,Ubg/:NOT,JbTC1MKOXJ1@#3@T]-X\A@IO?Qg_DVd7]
F<VB3Z3H4\7(8I[]aHBP;_CW/Y<_YH7#+B^OW@[&)&^(89ZP(-XZR&FCOaAZ-HZG
.cMa\3=^fM3_BE:cYB\:#<fIVSHAX,DIG32Of5[2M[??aPQK5S+?,^.7L4HWSB]2
2d@W6\N@</]2LSC#8.K8Y)NO?4B((Ba7[UCc&^Y#1bgV72T0PSR#20)R9M7?;L_#
(a0E?P:IFKS_E9SAXP^He^8MB[9;?:I@P@?bNF@#Y,WM7C_-L3D,VeXc[^H(U_HX
Ge;1IJ+=@#;DKHI@63eF?(W:FDPSEE;&CeH[-MG9A7WZO;,;_ZILJ=/8UM]\FIDO
W,&@c/]7fWVK2FJ1D8AaGT97_T?11<Xd:<@@@CP-a(LIA2YJa]<(>\<--b>baS2G
WTJ.6\?3?)H5@LaF2J0+[^-9V5bYO;H;2/BL@g^&;41B:]ONbAF,/C.^0^G?BD[f
KHEJ2MU]KUJXDHK+f.+AR2>LgFDZU,GeDASM]@=JBfD,;QB]bV:X=W]1G#fXd;.T
=G^e;ID;@-CV.D7d<@)UT)UG&6bKBHS6I3\WVBL2fM:AF_6db1O8=HR-gY>VOeSF
7G@.ZY=)_2WVd.6W_,Q#^LBWF.B\TABMeD/cEc<0?^+814>g5AcI8BU1=.(VAVJd
Q<=L_EV(>Zf7DW_P/H^72,3X#.(>E:[fGCSQAR1f#1TTZ@^92]_d]RbH4A3#,+0D
ERI0PSBQ8f@A<Q6>E^C8(8O38487fCER)<#+F2c#f@,KPM)>?WBIUS8LWJBBC,[&
><T07KCA-9^>O7CQGU3EG1/4S,R?6SD@a]gHJIg0HSY(M[X<=-;gdF?gHS1T8b;[
S6II9VATKE]+6X[cBZ83b7W7,LRYJLH7YU;\@9[PaQ<>gZ^C,)UNB/_143N/a@Z/
>8cC[66BTDJ;\G2^fC5HS],dF^NNg-ZPX2_[(YAQaQDc@JTHggX>5H\d_R31^/a,
#&_V.[&a>Y#.a<b7f_aQT5/D#=]dNXL:KQKO3-V]A0IO4gL9C6R+e(X8CRSDP0(d
QZ=g0RUeS69cYB;3CaU2c#PJD;9@B]@GX:N,5X2@:)^Z3/=ZN?=K8+>3\D,+J)5R
T@ZbY#N#[W-?#R^1@VDgf;QNfP_WS=5\bEHCaPZ4BaJ&R..d63XcTE_JfgG5M4DC
aBe.3A9C6ba?F))Q<SeBHd5D>a4M78)IgDW_2ggeZ1ZZ>_@,Uf>-3g(,/DXL&1De
fO8)=Rb39S]G[/Q=;agQT.ER:7aHIbVFJ+fM&cMMWa_N-37OU&W/K2LWV70P(8Dc
e4T8Yb03,B(d=<_RT-aEY6_fIJIUTLD9b#PFaL(@g(^c8Q&PQ_FZ(><P.a\M(.0H
Kf4Jc:0J/6W]H<9;41=5gK/&KFDD>K4,\T<5+N6G>2bY]8I>KRd-J#cU[<D1Gaf]
6GBLC<SIcBE5D_B3E)<,.E?2+21>a>,4Cg6K]\Ce>S/^L]+@A[g(&E[Y95M]\2.P
aM/RN0G_._8fPL@?ITUg>M&\8D2b6N-d(;GAN1SV).>QXO(E2?MM9SWXS/3fO-bG
#A-9QC6V;A\T93TfKKe+W3VLQ&<MM2L]EY:E7^\_f+>bWZbIPIS.L^be22?_@.Ab
4\XV#]K^^JcF1G;>P9A=:RdR_([C72BRfaC0dD4H,_)?]ZSg^98XgF4Af.<MEH7I
SM1\^<Q.]A[].^@MfeZQ?=E@BR=,KF[UW)\))VRD(>=ID;-)P0W9-U2B>[NH8DVK
[R&6/F#MO.,^.H2EQcb[CE?[,bYd]+VOKS+ZCf1:a>HEO=F2VBY7(R<S][:S=?:H
(0A^QB[QV5O23WW/XL3IC_2U_#QB9:aP>ggZENZ8P0Yc?I/^cU>Q_<;T5<g?N+5&
+/6OId25JJ-:5?NOIRC5c??B.7fM4Q)b_,;1&AMb/8a9_RUFeO\c^LI]PM=:b\]0
U6YIZc:#MbRNJ8WYV9RC.LV<(?P.57[<+LdAfegW<W,2HD:GEBgVV326G_5K+PcQ
,aPFS7DQF^gZ](0OR>.1&^c&F(S^C-K6D0a&B(D;9W16D5WJ,Q<.(S?6@/FX16;^
BZNREL#/VT>g,30:K2M&-^;G/[Y2FW-7>P)eS^8b^1[;\]?D+:_7_RaAd4BDVE:<
SZ:QX#GYEG7K..29_WP82&CWAN[F>M=AMU2NB?,&YM0H]68AC+PFYY8JA=+XV0T>
C(6\a21Sb.XPEEf.?D,CK6@aI?2O&fQU_gV5U-3T5Y?1/D/.,/AgW>38@GB0cS(G
-2\1CC+/IE94PVMR?)=9\#G&W)8ZbePd5?X7-bYGD=HWf9FbA;YeNcW/NS(O]ULO
YO+B&ARGDSD_f-_UM>9HR4NC(.G,_^?YDE;R<M^E_/a,.2HBIN.Ygff[PYZODWF3
9=W<6UL4].A+YMWU<NAW4MI(fZX[3+6eOW/0#2#Y7CL7H2cbHSK\:7d+&W?8UM_@
N\E[X]e<S(a>Q9>b.a=>Z/O(ZDBWXCTCL1M]^>KH7,EN,;MX_?:b3;7)49>+V#S^
3\UF\WQ;R0:@W&&>.4TYYW&,Fd3B\b>--PZ_]FJ_bO_CAX;]R_#d=.dC@@@GBUd;
cO=-0?ZV4Tf5_1f1:XA)?O94AXYH43#TT<M9,FR<Z5W:T8Wb?7[9^BRbMPCYS1,9
Ma-3+E=CK]NW5E<T\7XeY7&;,KJU?TR)I/d/51eAIO_AZH#&-cZSUa-O1_1:8.PK
O6<[9XA.;<DXK]K;T-]-_F4(U.H^<V@M_/6K#3ANO/@B=;\:45>CK@B;>[1dWfIb
N?PAg<->4eea#R#X<1-aFZ]K(,-6^O/+A;)R3<4_d4ABUPfW0R9^OOU.LKQ13+f;
KN4TbF1><NRJE3L>/=+=^/QQHL;OC]^?T<)Za?U_)J#,&JD1Q)_^MU15D^aNHNg[
C]WHI+,a)f-J67^45#V9_6Y]YHMZXXT=WEW]FeCMFJF#f^?+BgU-9EXTfc<G(<F9
+I_9c?^@&-4#ReIX:V0LVOGI-^EgY=\Mf3:[:>,;[R&J#=XI5^QeCc@60E;gH18X
5f7XP_T437\_aRc-dD^6_Md[6N:U2[^\HM/HM_IOSfIKHE5)GY:G#]^P#)b:KIRJ
=BJa:_]Q3^-8e;-SSBZZ/.+R:M\JCfPgK0LOE2)LdfW6/@=GD&:]4(IK:/RH5OT1
BbT(31[466)R;@e3N8.+[TX8ANU_9c2GP@7<dJY<0=2#=8&N9fG\+DZ7f1GXW_g^
&A9N(<LDM^Q.&]_;d\Jb+]]EC-(T2\QF_d=RZ4QRW,XV\ObH>0]#<^?-TD]L(caQ
U3d5+GeJQ4-;bEOJ:=bZQ4(@)]NJd7:SAABTU#GP3A-,4/aNF=4[=GYFTP[_+,A^
G8H(e6WK/DW]@WAR(S[NP2H6(K3(/QWL7_K],)D=g[<X(,,LPgEe?=&d^L,K)B>Z
IE=PB<FcX7H4.0O[)J^>UF4Na#J4#A:YQLLTID,EM5YGF#YSJNWO_GR>]b/:f(TB
_LfVHUZ.f56-a6Td]Vd84?c#INe)_4O)6&M?E/&EE:6,++,SC\Ic?_B<B1IIF(Ze
aU+;=YZ46&IIeU;Zb9I\W=KZJG/e_;09YJ)^C//MVg0[gG:YX?LVAT7[.T10cb?0
[Y]b8:XNTEK[6:N9E7Z+JS5eB?3ZM]+gP^K>9K&>X9YY=d2^&.^B#5T/(^cSX[R8
c\FZU,G8gZIUWWB0<Z:PEC4F./-fe1VDW76EcZEJ\COP1If)72aNMC+]PC<7<gcA
eC/2#5@3J5/4#0,3Ve\>561IGOA]#1a@]?8aD9Uf_C;d:A-^WRU91>5X-9-O>/W^
?D.O,5U6ZG2P2_Fg<C5,Ze2HV<N1^?4M=@=BC=COg5><WC,P\]b8=(^9f<7K+dRJ
YP((IWc&PF0N9)#_7T?dg54GVDgbYOJJGeKaL;HFMTZdR.#I:-./;]]^ZGZ3C_DF
AdQM@OXY(4J?G;(X@3[Y<e1[YU.IV4[N7gF,W#)XY3CP[J1a,VbaS_5LLV&#<VL#
BRB+M7\^UVTF0\Vf/7g#5<[>4=;g>&?7ELBd/+RI^.K]PXL<H+T6MV_KTWRK#,T(
5c\eNH0<31=aY<8I5^AL\AabTWH6>1_7;O,)d?RG^K0+b=V07+Oc9A-Ia01&_(g(
O./>^+8ad/KT>]KA1Q2^L&K4_VEN>,a+KA>K-Ha11EUI+32-_@^\Ef]>@BR#?+S-
GHgNO]e9<<,9WJ7N+HI)W0Z?:9#&5GTY;/;XOKM,MLS&1TU?J[eD4],=6/PDOGVW
^4d3?S8<_\6XNY-ZfZ&\YF8(e8.3Rf>a=T<@#//E0./WL+5^K2S9&CZaId8_9fGY
<#GR\eT.I<=A(E/=9Y.PQ:=,PMPY;A45?6d/0)325/TBS0++dJUY]J1c/,W/60;?
E0NP#69N):AK3+DgPQ._D3-M=IDAZF(BIC08P\[,^[=c\O,IVYE]C<S5P_BS&D-C
HOM1</eQ(de_&@f(d7S.K]&3O:HbJ<^\:fM]2D?#T>W2+.97PK4N>GIHFgVO3@N3
,gD5\;_Z>B9A1,Jb9g=1YVFV5ZQ0KA/?U_W0FRFKHgO;-R61BXF?CebR&A5EFe0g
3>FV7L=(_X,2N0Yd6Fc]CcIQ_D52IEe7Vf<31NQ@OM1Q35O)\)L1VQ;=+)B0,=(g
PXX023GYL#g=F016,OB)4=WU(0,[<P\8MQCPC-GELI7VF2N5f@IL6ESa.P;?efWd
>_92XT(5J.[;&/H]8Q_=-E5>2X,0_J\-^DOPJcHDDLW<RMZ4_d-eb4,^MbH>,aH9
ZG7W^E,P?7aZe6<TXD-Q-NUKQf1Ke/FZVCKe9+1Y[:aG&,#QUXAeHQK8=ERYA,#N
C@BMc\5ERW>gN\)BV79@eZI]/PGO/=c-.2(?X#JVf+?8:b8H6OE,gbb+6H-S6a+6
D3FP8);1^W,(4/B:U5W)?7)@d#?#D#W3efCgA_@9I[L?MXY(4=3L.QJ,#BY];91E
Zb)G47e\U3J.Ec<,H:F?CX,HT\94+b(2-O\[OD(bAZG:<3?=O.>D@-8HHT7M]YA7
ZZ#GK.<48+Rf=cP+g_<UD6AL8OQR[-,L3f^dM>Hed=C&O_R?dP]H[).f(Ng<QBbT
V-L5.VJ[2J-,^9,-<N\<S,#,b9X#4-L4Y^8\_?0I\A4?=TC#R+8eBgJd8IgAb55U
5f?MID^<&:U0):PW.fDXEI38AOS-BJYEW1PI^2W\I2]?;8]/(&@+/^X0JP7Qf\EF
_dQ1ZS<2UgLF]@A,/O^([UVQDCNJ)R0E^XeCQ1Ka6a?(:>0>WJJI[W?Q+4T.MEBa
f&9CD-ZYRXT_QJOK(J3[DV\4cdF,6c&_#1KN#1B/M2=3gaRN0[ZYba_5THDQ+Ug6
dIe=JEFd)H\&G:W&V7QNKd]c(20dZ75[7f34c_b3/)6FDRLB,U31TF56K:LAM.CP
J73Qa>/OX1#c]&(1LaS_[Me,F93@&)>+8F?&[U]eI;f3\+@E,NO9\5W/:-Y)0Z?b
)?UA-BG:7&9ee\Yfgg_gd9c1##FL4LW7;O,>QQ,2>-2B97J/Z21J^)-gdTd+c#4Y
If.[f#/eG4D6^/.Q.?OceLOeZ9>&Y>)3I;,&D2/f+f;MWR<GWdCca(G8(P6N\U0)
-/.-T7X[DSX(K./@I2[.C&@AJR19AS6IC-?[g/X1-<ccM.CCWC::P\ZAE?c@SJVP
4QXS?IC?YTS?Y]_V7)CW6R>4b=(]?+M6=KEMbIb-AVA5C/_1HS0J?#dSFTPaPP+/
:^\<_B,Z2C4:/XV493ZPdPJX/6)A.Jc;)eC),<H6d);11F50<]R+_:HYT\G+P>GF
4dI7A1:/GfP#ceg/41KE5TbaE4[7d,2,4-X<a]N,Z31__3TFT+7/R5KfC6Q2FecK
9Q::Nga)DHgF[2?J0P+8H@=W9W(5bGXSeHFD.gIa/?:XF.N5SY14M?);0Dg]c]1O
gOf<VK+F7J^RPa>KHBI_cGQKS8O3Lc177>]]8]?Fa.5MWHb@9D0Z.7&If+HXILa[
^FKc?9NK)=H6d43(CDaGa;@aU38_\?REG&-EC.(YEEVUGY3eF[B;Xb;d[Q4^5;Q2
LfG,\V_,2\aDZ0K-N6TaJNV^E>@#\[FBCfWWe./X(D./XARQg;)SHKX<E@^Sg9@O
LE)bJ^/9FJb1QKJ3<?^-e_]Zg/IU)8:CIS=fNH/O1O#1+94^O,@P.[PS)T4gFY5Y
P9##4A&T?28R;Z:/PS0f+TdY&P^:aIYcD_&Zd)KK+K7WR,6:-#1?,-ILJ(G^WP;+
4H5J6<GV.</-c1&ga-^Xf5O.LU&7?21_X;G,F?_c>RL(>UR2JU7SC(2CDZ@_,.aI
<eLROgB\^d,DJK/CH:_W)<gV#ZF4D/8[.LXI@AFPg6]]U\O3_.>R4/6@5[&Q6BU-
():)fN#,^.HNM,>b0P#6TbKgLZHOBN)6]E;4N0GO8T-F-O#FZ7TCRP::T-HG8X0-
??fJI@_UAKg(0U_Z6M_P#FSLT=X6A2KG=N^c()X\[SZc(I85^_[eJ]He6f7QLX2_
TAG&??RNJS5eUO3]W\gUKPgL0;JYE-[Z(\B>QK_9W7_69A</)#[;-22HV1WQ+XcV
,&6]TX+cT1-7:?E^+?A^S<=7gWB,5_U4gQPSDb3Z=5PV1IZWfgS.Q3Y4;URQaZIR
[\3:7(\C8>ZWPFHKb5JZ(_JG=/1;O-JQZJ=7<MY<_,2gdG)5]Q1_,d3RC1<(WVT<
IEVJ6GP5WX^9_[bE/;;J1(K\]+EY&V=^V]XY&EHJP;Z^)>8XANO,X_3](64EXB.K
ea38A,L=gZ>[3cg<GdOgSS-TTMe^.ZMeMc/86B8(J]0-._5PXUQ(N<b5SHU(4;V3
JQ+Vf<;WgTBI[?;;<cb>#>aMDDGM7-J@XCQAQ:9R,47ZWL>6\cMd2K<,3V;JXU[>
,1Mf=U(PDGE+fe(VCLa_?H,J5N+(ABH8/LRA:Y,X;QW=Z,e#YGOgM(\_T(FM[&7T
4P>TTB<)8C=5U&0#]bN5?Jc@f93EcQFDg@cX&3C6Y)T,^A:-EAcS7SON<QFSF>K1
>e.7Qa<=#KV:<PG#I)W+)XZB]Y+(Ng_\Y6;BLAcP-L5YIO\,N&;?626=TXMb5eN<
:a?WX50RUeJ+[dB&a:cQ<Gf83XE,a&NX0U^C=^5ZJNE5(DVFYLRb4>LMW/=\;f3X
R/&1GKGd+\M9&Ef865IKSQ_^&<?2BgW]N,8>ZE73K.6ZP7V7@JVa@H[d12@e-V>,
DALDJUXbBcQ?G.KN[5AU#^?6/]D&LU\>c6FX)IXQR[OIWacI_]75X.,\fY#2BT\)
dXTZ&/g:_LF,;bK+[)bcYFAaI8-F(/,\c&46:2e5?],a;Gb9]YKEX9A6?2FQD.EX
LS]E_J?Rd_EZ[B^C,D4RdY9P\,WY3TIc#P)/:=G<A<6;?M[MBFKQb8+Z,1^NL4;B
QN+WZ=45UX1P(&_.5DG:\f)Z5KD^OLC?<Z0T;)LT\DF&a^M8:^NY5(K.E?6CR-N2
4Y2\51db83[XH5T><2V4T:)_WM;dUD011Eb7ZD>#M#gY^E+#_4)V(^EM:80cIQ_8
HA#eJ9YSeKK+Qd4_CY=H1F8B5.IP7Kf1g&(<=AU5Ie0@R[VZ[F\>&KaD+3O(L2X?
9K+d.^_]aTN>[3^4:Y^HW?-XTTVPI1N^?8=A7JZe?XD(Q1eFWbe>2]dS-b6b)5B)
[Q1gE1)(OPDTN1ZS[[AKUfU)/@NW+X6T]-<;;1933=+N(6dOZ.TE<>YaNd]<YdgK
g[-X([2.K+53XHDD8T)E.BC.LA,UIFW;[/;TGPU]Bad#RMBgg#TEAM#d5eZ67ScX
/E1M.^,P.A_TcA3+5_5MeN)R=281;ZAKgR+)_;U#SUMZZ3;UM&<YE@OC_;R,U6I[
A537X-ER>KBS?)@,(0,N57VB5L,Ng<BQ0R/gR-O(CQa<VPIMBUVTYE,+;MA=0J4)
\#/bI+/1Sb#Hf+U(IAVX.LT)(ZPZ.Ed+4-g8f7?\L)fJ9M.-\A-3&]X[,Y>4A6e>
]_]?bY-bZ\bS3LQ944TdJJ=b/^8<]LL6.)bQ\OB2/:5\BEBB\?BBG;/VF41#b@=Y
I;E@OD5BX=STH)+)<a]Qa90SLO6^B+&2\[Ga;?PU<X&2SeWU?=JYQM/CYL_YE-&D
2VN;FP7XJ#JPK3F@WCT.)ZL<JQH&gQ;de^?R=Q0&;HU2=0,&.^;9f=1P7?L.e+74
=S_V<^<e4P;/7KQ9O=VBJ2B8:1dC]@(]F#4KT7Hb&Gfc;]Jbf_Uf,G?=F2J&M2aC
?Ub5YD\TFcc&gg7+f&+=Q+T/Bcb[\M-g;5F3EZY?VL^2V:=>O1/a+CN]cKR]=FPL
6>W6)=e<YL);M4#S@U[cP_I]AU3YI;\?TXFW6LIL50#6NL^-cY/AVT.O;N\L+B3[
,fF?WR7-N8_DX&2#c57f3+HgEH1E:a8?/U)-fB<dNPL6KVE3e-P0A0==Q5)@9CHR
6=.g4M-=DM6HE2fYM\#>[A73OC^+=b3JKA@YY2)OR)3359Ce\NG8XaDA7b]41]:d
R30(aa2)7bT3,6Qc(Q<8,b9=RG-dTS=VUQ,IAD;:CFUJ0>5A2Q>+H@B\Z6[g:KGd
>KG25PZ?[)O/F7+8G)Tba,4:>cHS+YV9RL2Y&4b[fe@L5J?HEGf?N)\<;\X-+e,R
;9-[G,bI5FF-:INcK+=/G&P5Y33Z@C(Z.b<dgJ^,/27dc./^P)>9_CHd9W(ABVYT
\_BN#408eC[/=O,/5RPA;gXV<I>&#M83^eLK7\RY-cW&K]5B4PD;9,KOWU(aeKV@
VW+>e#SAVO[GI)CP;@(XS,P-]\/[H9a8Lf3cgcg/Yf2&D$
`endprotected
        
`protected
3VBQINA&R\P[#0\C/a\d.GC2g+B-K_25VI#ed>[.eG+0GN4d4.C?,)AY#99MZ5X(
4U/Z5I\WC_>O/:VH)1aHTRaNEDIZ:UTN/+HN+DT9TZP6H8LA6>N&UXU;X.gVTJ0/
f2@=LR40_NgO0$
`endprotected

//vcs_vip_protect      
`protected
:F5U6a&fI^cC3OH6VSg[a^M,[@R<D>HU(.Yf-SfU7RB;XfaHMGQI3(&Z+6VY8)L?
+F>/3-P#_cW:e^?MDS[^UD1+#a)8C[(2E/K[@\5KQTS2-GU6O1CK@fP;J0f&;0B[
;,@SF\)CF7T;&37[P061Ue2MBcC;\)P,SIFf4LN&OE;45,1&5/9+ZNB>M#Na.NV.
6[8:F\7#+738X2CI+VM;__.^S/62_>=BKdICRgd3^\+b#\I;1)QJFcLXR\<&_/16
>M>K/JZ7C[W,PAHLJ20B#6W7IbD#F.WGb=8RIVWa,Z>bUe/<cNZIDF(,S86#M/Ub
\V,&&+TM,BS5/d&F@8;@:SAg@gW_D,TQ?-(M[V(=NUf)gTU=&<F/UW^;6X\1I=Q1
YJ0AVH.6\(DEV&#_fgI>#T9<Y\(QMfBW6Yb/WFT/bW:\,E6>\N21/()[DJRFT\f&
3.9e33+RH2P6APfeF8>-)5C_H3A.d=<O/7bRf7[CE66/+)V<H[,41f/RNV9c>A^0
(4K<@X,cSd4b(Ja^XANC_fS&7])J9f;f#]0;[@3fVIa;VWE?-db[RD]/f.6,OOW9
G+LV&eU(FN[.O_(J&GIVPW#Ea_>QdJPeBZG2@g7T@7LLS&R=YS8QWK+bdY@[\B<N
>Z5V:Kgc8:M<3:&QQKM,.40N\J_Y4Z6\\6JD6<P?-\1f;AW;&ab[AN@f7Q+AbP^A
GJ0:3RcgK[Z(7M@XbbA<)#Fe=a6EXg\.[.USNNSP;7?G96aO:eIHIAb+-&f^&NG(
F(fN9cKK#g^0DX:a?NAVd+SVB2M_b2VL&(9[UAW(Qa^WQW9V-<bU7=7f;2b0eaYL
_^^E,VN1YCX/2.E]cMNH4AR<^F(G0T;TRga31J4S_:CL,4&J.5/X2ObJK;@7/fHL
:g4]-=QK)4@ZC1L/4eEXNWZeG;WJ7.Y>M?OAOMIQ#e]U5(/P9UPI,)9L7X5gP9K8
BGE_/,TDY4M/I?MAB^(XWSN_&4WN)W_6gV^S-RX/^ZV8Ccb8TgbO9E]f;+J9Z^NR
).bIMa7L<\cTJ?+XR4.0=;J#\N/G1KAZDUJ;RJ+[G#F.VPO.ebg,7&38(G:54_[f
g#38KX],B@-b_J^J3U)/Y&f:O#g1D]2X(X.]=e5=Lg=8gJCg)0c51&54M9JM4@OZ
3/+8+F0_I:\9.^#__0NR5C^P8&O\&9T#)C]6D(NINO^c89J^NC@aQ+fG-[:Tgd/R
OZ=+TeFIdA[,OG[c>-QGT;FMg-CC@S3fM]@(_f-#)fAA=AVAPS0UW<7L+._:/-CC
>YaV9.\,>2E[HRggeZ-TX)=5d(L,VYK#6W[,ePTaP0cbB?@\WV03gdf#ZeZT&(3M
#gU1V5a]02(+B_@6R1O(W-<R/)a5N/dbf;GIHe)59X^V;H+c5&8]-W4FKMHdM#]L
/BZVfc-DXe:1V<=\N0:>57TY8+gYe,#8aeD33+g0D]+c=RG0_UX5Q.0HQ(AJ6a6B
.FJZZ7-#S1A]2bKP-RVBG@#8@gGL>WQ-2e,#W>-AK&NP#XXH7<4Q-N0WdD-\1(X[
G4=CJ&c,.)I@E)1@+S:\aXRbV:VIT3E&e=3B&cGJ1IDd+#O.,#M;IfdgV.1Kb>Cc
6]_J5TI-D@;0g-4;d;+dF4T^H@.de&NY8.D:[JcU(\08M5Te[_#Qd12R0>?,^]:0
[G+25X.T2a\AP;12IE<Z+e=b;+S<H@Z,PU4AVZ4/E@a[6;#<ZT=\?B(&AFV_@R]L
M](d/_=CH/F/K,5O,FZH\(FECI>)8UI.f)JQ_N?V/5;B^\bSM,-ZH-X64HT1Y^g8
]KcgK0a--8489D>Q^L.a@2eEQBJ4gOC]W;L#Jb5QDZD>2->C66M]C8N<3_D?A+7,
G##XOK,P5gD@?3IbQCMcRK=<[d8G=VJ?IB?]O+=N454<2L(GH58[YcgEX,+:9BUP
VL92N27JHW;1-@/FVJFFd=V@bIC#7L>9gTZA;JdD6<a>W&]/;=S5^f9PZ.,3f>P@
?c5@fV5)\GF2P>daF#NQ=dF7+?;ZFECT6&)DX6/Q/\)RG9EX2D&MR(LFY5=;0eI8
K2G1KGP6bAf2;90D+SCYgSW[4IC>bb,4C&T_0SI5E-K8:)]ISY6>=4Uf)6027ZPJ
>&^A@E9?XR\T;Q-)NgfN@I^Tb[^MUA&8)PG;e;b3S=PV5>L8Z3=,X.C06;V5\5F?
+L3#3N;OG[P:,#0116L,X\]=>3[RK0F1&<8YPVQf-a].N6+]6SP].;_7:[[0HM<,
f\#[PJ#GW\2B4E#C3b7.^Id9/&DY+=]RUK;X7fCX.-dR/T-M:,2)J..T.fF.0O85
/DZIU&>#8M?V)K(IXHYe]@@45&6;X7:4]_+/KUaVeAb,=MEYP3>#8K5F/_dU)@RG
eUM/\FJ_\/#2dSK]6b2#9dX-b8_(=3G-.2F@.1.UA)_UPXHa[b[g[=7dU&O;]5SO
=6CUbYQ>5aIdb3g?><Be\W4.)UZQ<;DY:->^b,9b..<:I]AZUUIb1T\>YX<D^R9<
dVXT<d4H1<JXS6O/fVSX0<&ALFFV1Y7-^DW>H3&/<@G7JZ::Gbc1;N@.V@D,62GB
3AFC6C.4_MDLKH-FF#cKGbRT16)^J3H59.4a8Sd17Hb0GIYJD#RP(eIA+YgfM>WP
\eY1SLY1KR8I^V=7dC98+Y=A^X6M@2YXa;X08a/a34V;#J.XWM(HbP?M#cDSS0/]
.9>K=g=?+L:NQ?eE//1ZC\BcHcWSSL,P[@A&8T9:_:d@K174K64Z[a[NgO6YW^NF
)>45&RgIff98809CCd_IU;;&-_&(JV>=5681fS&g6D/]KW9gK]aWO=C?VSQED:96
(A59<(23a2FLNb(gaQa9d:PG3bY7=,Lb8^J&g><HP<;9eHJ-E.KBU47d>51K45:3
_M9FeMOUA4=BZFK#<+PSg19#e6E()\d:fU;834:[\9@H9DK6B5FFXV\8S09ISeI+
/8Se^0Q)(D1/28MUSbEJ19Ddb;G<\?2VM:537a^3,_[aOJ/g&Kc()ZDQQgKg_@J7
WD)NWX,bFZP>(b>0M71cE2E0?:dYZGOR>#:8N..fCG_K=_QJFM&8#U>XMg\0OEDZ
e0-Qfb3PX#c_L)7(JgJFb-J145G52,(:ABfcP.0FKLNHQ/JI&OaFW3Z^Z=+MRL1H
?7@WDQD53<1S7[FZgW.R6LE&/ZM]E=e8&,c^]<L+F@@2=/AKC/E&O[HG8>6_b<9H
=U0d0=YOS#B;3VM1]gKdd,(&PFf\8DbONECSPSERVACd@NN]2N[[6&fP]d95JF.1
ZH,D:K8\_SGST6_6^@G>G7g/7@NZWee9A7[d73;=L2A)U\S57#GXc[Y=4+4,dUC4
O5<c#>c8CJJ7\#E2S)O69:GQJCM0_-&3A5fFFP;]BQCD.8N8cfSUe]V10T)\&R4:
>Z9X3V6>d5JfIUY.;<@KV0V9XSQ@CPC[_,=(INeG@/D6>6/V4S#E[;??]-FKTG.]
>\)GAF84V_)4=/5-K<gQbKD\@&[LgRYe]03D;dK,MNf[7FgDR/2#gAF8G;V\DFW]
d0.N.DIZM-b9/99J4(Qe50G[4c_SWDC@&SR8<TB8YaB8IPe3+V89.M)&[^RU/MX&
:b@M,)eC,#QJYFC3Q-4HD)Yf-5;A<\4,Dc)1O4)5;&:57gM=+/f11K2NLeGa24#-
9N;:438L(Qcag5XF_[MfGK+1G[V(cR&=DX+_4(/[-#MSEZP(1[(25O/.[)]=6>_d
FcfYI._eDe=Gf\==TVGXWM_gX>=D@XCDY(_P=@8;KVZ&3UGS)C2X4J]W57;3EZGP
3(1CF<P[)R&cRCbf98^R1e8,-]]CPPQQZEbSBG4H@7(N3J.D^T-<Jc2^YB,];])?
PbIfbC?9CR1KOKW\,5PbYGK?5D(R-K[)99.(2+NF<b\SHWcY<P.5K^ZO8@-8/Pa\
.fRX91OcKY@LEZB-K++Pc0Q3QH;QJePMJVDK\?U_0]?_<W2;f02QXFg9E9EKQMDA
/e7]/RO9W.g8Y)f=QAZ<fU;fISBc-8Q51>/edO59,^bg.PR?Z4I&AG0>f:c:#FMT
\Uf/[OUC=LgB4Y??-^ZIOaG</BgA(\<\\STK8(2G[@]5C;SIJ+5JbcO:TCVASfG7
<OT<-LNR5HEL9PVQ,9ZG.DCK7T=EE-7_.ff?]df96Q[9aaJN:XBdW90NBObT)[dg
+f(?Ka#4>Z079LPPD1fW?]NZ?DO.8?)D<O::2Nf=1G\>99Z-0/Kd02_W3e;)8Q7b
S@e_I3a?W8[aE(]FU.cZ6&LSXJMO&KO\R/&PLK5L6V24<G7HK6([gbT?-O;b<=@7
DNIE_8eP/f?IQ+[WE;,SKb\F--cQbR6F>UJO_@R?,PC;P1LDe<eOV:5?K^FWbM_/
FI\e&D&2AZE92BEH5NUN+F31T+@M7+?Z;V6-ggYb66C,Z>,_g:dEY7UJP#)L71/[
V/B-_,0d(]5+.b6^R8)G82)DcRZ?D+CbUC)NO70R6\6,VP:VSTP=A.QPN0VF^LJI
Ze\K3EFV\a9/\#KD__HC,0<<:PY>b_@aJ72gN?RQ@J02NN4.H0)8c?K\</d98@V:
NP:H]#9:\FHA7fI8@ALc,P^3YP\Ga8g6X2HG9<Z,a=76[M#Q<ST^O8K>Q&:++2\(
#&1I-9N[FTF=M5_2TPZ0P_5^U\?97KZO&W8b1J_d]PA[cHPSRfY\Nc&<IM--=GdZ
=CNeUWJXEF-@e2;2+DE)U^OC<(I9Ye;b;\&NJCZXe8@RM?Q[IAFHR-c+Y>Y9NU\c
CW/EGRL3<9ODa=CLW>5]gN3JbL)1^JdV6ZWXM2A_FLY\@Z>7,ESHg2W^Q9\e0^NQ
aO]V@[VbR2>ZL&IFf7=+ObDVU;Z::OA7CC^XP,6R/AK=He97A.^=83X+.282cPf&
W3g]5COQQK:ee-Y()c@RFZ+LXE]NQ#A-B1MeI>P[J9_91b(cSUMP=O^2PYT6W@(C
;/SQ@>[;JcQ-H\]CdUWW+P5;EYV#8XUYc)M@7:6)L/[J+YW,8PNd30f>a+6c0_Za
5>I7(\gUP8g5d?&D6gZ-BSa)V<Z>[f=6T^PA2_,E3DH^FQ&/E-ddKOD2_>G>]C)O
^f1NEBB2FU#>DW4UC0CZaeT7,?B7Q]JHK+Td8M7/(E78#4)D9?Q350VVB3aNg:Q3
RCB;[RKLPQDaKG&DVL<@-^H_a.F&K7\QM7Sa&MU)]_52gUM,^ec2(7FVAS#_9.I[
=&dOMEH_RgYPPM2C7J#gYH@WdN&Y,W6(OcfL;L4L048XMfIE(2(E([f>\&./U7A)
N(C9&\VbX>@Wf^4^2V^J/-I)3g]5O^GD,[B^47e](e>=:U+gH./I5,Bg2#U4g,@5
ggfG#F>(66R#UF[;5F+g/_#-BWRBXHGM+JO#TIg-Y^[g53VAPC&M@g^:H9gQ)_1+
<\.=T>S+FIO&f=7SeM+.fGF6gF7JLU/VFHEbJ_5fc@8=R#]),,XXPbB]2E1;RU0H
BNQLLLSggI)0N@^_4+XCFc=Ha87)A=?DS)d6L[.NHa>P1JVZ=)AW;(VacQ\FIOPM
_I>9?H^-B8J#aWNL,IW/]2M2.>9Y&2I=A]S./#E?^cbM-dY[JATY#]c8?E6=\QVL
Ca<P^_\Gb.AXJ:e&835-fF)QX@(R)2dVLY0X_,Y2a0\-(X/#FJK5@MbR-<f[-aN<
2_fLgJ@O91^VQ3e__JYXVb+P^,F/I0-AL98Y8L5U#)[-Lc=cQ8I\3<>4,ETcC3A3
[^g@d2a)ZXKaCERA^dS:5-_?H.ZMa2DT3f;VO47-WJa..8c]TcNX9Z^>Ub)Q(MCd
-Tg_\O<Q.HS/N3AZN.W]g1#9b&e/X--.=[UObXV>BB6(g7ba4P_M3/SG,XMASX-:
<,S)^3GQX#(6\b9BYc7eA)Pb,b.26(KQ):#(K25T.1Q@YZ;U-S+_4MbWT;B@)aXL
8b)Gg7^F8?>cNRL)#L.bc>7#NT+1=Od[_)@NL/GW?K@TdUcLA5I44:@9d;-]GNZU
fA+,dD/86Sb(/:a.=<-XT>RZVFN@7H(,_\(>#CC501gDVF;<T2HQQJGWdO+8TD;[
I_;#c;ZXOZFPT(23P<JB?7(9KLA(S(8#(842-]N>gcQ(.d>.\/E3fZ@.M&P_P1.K
HCTGSPc.<<+@/.6b&73Q]Q==],<>=VK&A^<C]dG@6=\],ZLS6MO]<<#Lg8L;;.N#
E.&(=c;eJX^fG.+I&R?&d?b)_H4ZW[1Y403IK07_0c_M5A@g/WVY+T=LbY2)KF?b
dJDPDV#)RZQbFIF^]aP/O2EX@TP_gEQPT646EC=M6GXY6G^7_2Z[>fY:_Xe]1+EC
;,F(@?aJXS,(@:HA9X([Id;,+^,beA<G,WLDf)GFUfc,8G9)DeT9QK#JOCP&@4QR
9Ve/BV#&bGCF4+GP3)5:##QR9IEL_K7_Qe&O/IY<:4TGKY>9@.K;^<FYJ(;IC[f?
g(;9:/VAGHXRRRZ]4/#YSITXcHe]ZcPX25/+bVgb(58HHZRP0eG/30Za4&bb#Xf6
QdIc0fXS+U,ESCRcOWJ48AGEZC>EF=1&bZJHTAHYM?)W;=>f2]c@:[R2;IET+6X^
SF,DgD23cVP#5W5QQMQ9R=]3KI\2<V8;=X2>OaL^.5:a(15:VPdOF-,b2S#:UQ61
GI]7M[0G[9@>N;gcK:Y4+4O-Q=MRNNH/@;+?:AKM.-;>0K275gSHb4ddX+S(_Yac
()_P_KF&;fLN=UEa8NAcWWR_9-)[e@gf#6S_2;fO^KQ>8W-#^#<WG@0^6MSS\DMc
M2UNZJR1U7[+OfB9a8)WCE:]#bXP/8>78)\4PQLM#BC<H9UZgZ00GSc,E#QWfY;?
SNfIKX@]Id8)+S)MT&6a@7G,DLc&,Z)7HCM3b]BV-.?f=3?+-J#NFHTf@BG.S-:T
9GFIeG2F#F>#^T4,FAMAD[cK@#B74Ef</S&[,Be.8#&9/N,7?Bd@EB9GQQUa]Z5F
:F0,U=RGO&-gb(M..?G-HMQ0a4?O6Q?0-O+T##]>T53fJ/Z[W-0WgSZL@b[;49G7
SH<1;I+U;<B?@A+8f]Z9g&?K^&-1#H<0_,)U.KM[834c6H93^Z2#eJPIG_7K[ATW
^\Gd.TL>05:bG(#F]c@;3IaZ/?d5E5?fb&IHaRDB@A-=#=+ARbHPDD5C+](>)g5W
9QccHFR1e1^f8]0(B[=MI1^.Aa1U78K;c1WP>/eGDB2=)NP]ae5.WIAPLe_.J[4b
Y.G1CW^LU2EYc99IIIF&W7<K/NE=0H0?b.?Q1NA3cc)0YAP2.D),<6I;W6D_6be^
cAS)9;7?/<5&3WRV2W+cgb2?R^JRC4MBV&UT,LXA5df=R1e\D@(4eLHQO/H\HWc&
:^7K\#YY75.8HDG3a[PaeP+<E[>BO;(0:X1R(&caP[^T9H9@fF4-RO5+gB-Ea#BV
U(^XB/]=@Y91=\.ae.Xfb2bSV<OT76#AB5.0C#3[\c#A+;bG_Kf=O-S55C3bc6C8
IT0@bB3fO#1#AMZ\8>+XG>a7H-FS=,/L0VL@+c+G5=b)H3IB-EKOSH;6_MH5YBJ^
-[1MaS3#g/PLEU1)GJW3N^fXQVIH@^8]:UJP_--O6F>\/BYQ2K:d0\^Be4@QD:(,
C4/B8O?,^f,gdGfW@GMbZ]I/.\#NRJ16A0+X^H^^48a=NM_6IF4D=aZ(QONFIHPI
4.S@?.Bgf7QK;FbN84U0NANRKf5bGWfMcVPZ6@C7SQ,aQ:b;4O2M&^>@,GcObc9H
IM(BM1HM5IMGL+.H\Bg>]ZC((-AS8Ld0gd6-#c[KM@Rfa\(Oa11Z.4<gBbJ276HT
S+b3cSO0AFAHAbQ@GZ/N<F7;AcN?B<)2X)G3#(#X9NVSF]>[c6@Z[LfIRe.=:JJ/
)?^A<7[SaE#\#T]CZ8/bXMM8ca13LTYAEZVRaHJ[2UG&+KHa4JU?V.W2.S=O9#J:
OL]W.4WSP6Le#Y_8B/EW@G+\OXd,>.X8&FbP[L>XL&<+,Mg](X>9gDNO1QAcO^KA
[?DJg2fBMU&?U+LBCbU#LSFBH@g3+S(VCK<5SWV\WH\#c;VZWFeJ#F[H@E:(&K-H
1&gUEUB^bR@7SQ&\XAe)+S6O977L?>QD>dI(6(Pf6d)6P70Gea:4KFg>JUQZ3gd&
XE6#,d;Pe,,3BLBI<WX#DCER#Q9J(5[Ob_VVABI5E-O>^3HSDE\R>CNM>WAHW&FS
eV,9\56f:-3<<+K.I1aeX7],cM&[[/J3[[7N;LQ1[4FJAa?Ve_F.6(b5]b5Y#2((
SN.V;7,P6C,bRL_aRb+IUP,H++7d[2JScSF0OEH4c0==E#(+N4b[Z4^RRNN?I+@2
&ZB8N(.7L>cB1=6g.gZY.R1^JU2OR9-7f+WTd6U[XeJGX[=38.(eSHJC2GCcI+))
/H;Gb[Y6+;a7G2Aa1R?:<+T^B;cQeBY?YD-RUeDdGFOcJDC(\6BI2d+8?8HE&7\]
LVg&9:QV^+_PYXXKD&C?X[_UgWIE+6g0VJ_72:74DP[SWfadIRQ)R\[<8,2+UIDg
E#<C[9=:V4CY9:a,fa2([(K02]2>6#UM-gdY5GeMJaX)N=d/:_eaPF57Ra\2NW0[
7:-?AX0YEV3g4.4)LKKS5RF\M9+@9b1.0([-63OJSgY^#<5L;ME_4dS4=DRGL^O3
RSY@\LPH)e27-Q0H)IQ0WI(BRCZP<2D\.@7UIe?57/N@:GbR.U8N/?(JTH@J8@4.
dZJ]MB\X(2EOC(#5SfaOR1e9\GcMa6#;6\2d&UY&1B>>,G5+Mfg=>QK)?):]-97)
-]c9(.EDGcbZW=eRA_S:M^WEGQ+&LX<?6@?JHN9GY^Wc(\6^DDOa?Kg2dP),)fQ(
6/9]86AYS=QD_c2GfVM^CGPIa5eU:+Y=dA]fNAHLP5Gb;YP(f;;K5?d_?D-P]SDb
AgC>b=#)E#9eW>SMA9_&_\/C0)@@AF(;@KT<6A3[#;4-65FL[98/O4MS37QX,^@@
FS-9T5HXBN1g=e,dc;GT<QPC?-70M<1Y0JXA3OgVTD0&4[?#Vd@+QCSZVN]XNF.P
FEagGX@#<5\@e#-?J3Fggc0VbD\EB.C/N_.>?/\C:L_e@0[VR>B?A?M^7E3Y#L16
OW<7]Md4@>GafKYQGZ6fYH,L1RZ6Ze1JTU3R6.G=K[Rc#b,03@\9Q8LSXK7=:\[&
[>-)1SU&WRfF,bL)Y@D[OA\a80gYK3>/9adeU-W6BF>?^2@J-e72WKe9V-]]e[&G
ACC@:Z8O^cUFKCaXU/\g(?P2.\\S9C\;a^S,)U=&K(EY2VK]>U&I/[,GRdA6OPUd
0YefXZYG35ZFU.29/R[75-@0)QP)f3;X\TFe:TB_YR)[5&ZAZb=H&]UbLT1ZG&YD
\)KZB_>?147WK.ZD2+\>OP<OG<7<V.D+J<HQ#L@FB[JU_3c#3QJc?5bK:K@00N\;
Q+149>>8Dc2Q/cc,X7V^@7D5BS#G/C)d(C:&KF?;0E70,aW92B-^PTCe_SQ#BA#c
P=e1.<TS\&UTLO/OSF6+=Be<dR_2&?92eb@N:4]Lddf,-;I8WEM\O\WL6P^:8a4S
da4OI4OaI-gM\;TK:dFR0<)BL#,&)F[VcTOdC_89]bf?b<\&E/1XY1&HH(SGS7CJ
38GL@WA0784/M@6HT]J=/d+X_F4cX(0U4YN>8cfg8\GS9CRGH7G3<:0,UOE-bO9Z
BB+)d;]7U^0:)AG?7EQPe1WN[:Q\c&8V:2G4B4=@PK,EYR6RU8:C):XSQ/1[bXQc
E;WVU0KXZb9383c)cO.S70(C9/QOU>N<N6be@A.F>cNL?\F46+VD/D/fHIaCV.57
?)KOYNOA#)#J45;B-Vg?8B2FB_6g2LU;_L6aRU1>FE7Bd:FT4DYP3gY4aBN(=.YF
eWVHE?GBD)a9>6JfeVXY+4fC-D<4#8_77]1.I\7+(gaY5X9GRE.=IF&;f2^;+Ncd
?I:LTI8V>\g&J#,<LOKNB[J)e3+WEa>D[>K,=\2:@5\I-_a.#YO7<_-<TE:[Hb46
U(A4K;RFX>b@JJ1S,7#:QVaLXEc#9^@>O)V(UCPM14^N[7e:]+b3eCT-L[:S0\AF
&S5S^&K-JNNCD9D-P[U0T)JIW-T4de7O,]D)3C3_6X)T8DJCI_C<9D[,@I_-B9dN
12BaB16&VW0f)#CQE=RSGO5Y:4>8EIIA8dfN[)a7U2.1/aID&dT86:D&9(O-Nd#W
9RQ>_e[:KR/1Q;638;dJg&?.=>5\F[M::Lb9ZP-R\ed4S-HRP?VFcA0Y(K@<Y;LT
O3cg7#@S@Ydacd];gK@\.QK=AD(DV+/ZOAMTEY7NMaP8>Y4>O#(W_1&Yc#d\?gab
BWC,BgCU1:Z9V1a8AD7S_^Zc@R=\f\]\RW:WU[3bQVZ1USF:a2LJ]9<U)Y5/e\A\
7L\DHg4:1@VYS7[@Rf;2bF?3&^U<TX9:_DM;)91T-(X[Gd]VTVE#4Q151dY<Z:cZ
&>4K):T?)a#C=#fRKTPR@P)EL(CT)837XBHYZ[Z@cBLK6G:=Uf@R4CG;LL5g[<Q\
:MS>JfG#\J30#E<7Ud<fFT(0-=JQ<&^5D64I1WUB(Lf\G9/JP=<MRK[>]9FX@Xd<
fZ7&Y.+.bHfZ)U]^<3\LH]K9@C,;8K]5gU/ca42)#D/La-7=NHMCLa^H#1/SN9NM
YXZ[5I6O?NAJY#?K5(K5XBD_QL87TIN<D.b;64W9G7T3A)-&2/D2(d/;?a_d[S/K
fYVCL^F+cQbaa40eff=cU;0.Bc80R;X+4XfC6JLG-TE]HdT2[+=gC>+&XQ-6JKIE
C<;f+P^L/=-B#-QIbA&acHU-[>0U.>H?0LFd[gdVU9FI7MN4#gXaY47=&,1G2DIY
a07A#99Q3ScP8LX@@\DYXQO-07M+\BedCG4bZ=/>GMP<<FPY+0W5?H<CKa,d(37/
^MW>34+J:cXDLSd<TRFFRSQ+:WVF4C4Lf=ZebbDc5TQ#a+Y(Zg^Xf7.fY\3FZ11&
Cb2+RIW>^1?Q(IHZ62E73H1HNKH@SH+5dMgd]<XM:,W)IB[=4RE2HU+4RLEDLf<:
FHZ3N(Ef>_TT/<XNdHE8K/a?G#b=_7V,HD7S1/V^^?O88KF(ZWGDD<^,@g,Kd_J;
SR)[<e4:Z?S_>f&\IQY.571Ka#0AQ]-](ScCJ5.M8Rd)0ZCSVT_fCLAF(2YW2:QV
)[X:EgMg(gOVD;Y;&B,cCC>ef(J>GMFQ:^9XCZ86:\g8>HL@54cQ]18aA[2]D8??
H7=H<K]\eE+e0>0egc(FVD[>W2()cP-X7,4FL]>G<^2e<PV&B2,LL<JS]9C.(9LZ
=@6&[M>FV(LQgG2RdB@9N37@/.1N6Y5gNM]VCe:cR\2>2B[BG7->5\ggVU_0F:2Y
7:X7287RFcb3T)2Rg-;0KCAQU;>UOV.MIfdE#e7b9=^aX^)<OU-gHScE?KKa9G7c
U70J/J2g-VBfQbfWMZOcEdDM<;:H,HMGOYJ]Hd:OX\Qd86/_CaUZI.Sg:bO1.1?_
UF9+g#=MJ5MN60>0eO6aQB7R0(.bB4JD<Bf5>_)]#e8c,QFXC>F+3\e>WDaD2T4O
YG.BI;&-_TWI&fLfS8\EQ@IE?_545&bDg_I14_#U?30N(K@05(]QK@(=U)@P[,5=
0918<&W>2KVAO+2TBXQJP>9,(_2Z0\f()W?08N.<9KdU^Ne)G]a0N1.PaV;<KOe_
HCb)_\ZHcaC?=UK\^/5:[<M7,BaXbC0e2-Sdd-;28J-F7&b;]P[JZ1DH4aRP2/&B
^T^_N?I9=[=Q@,4G]9(V,AGeQ()1CC@.c,WH4--B;S0;b0gb?S[ADgH&7Y(8-]MO
d9_:,^#H#L9+LBMT22e21+3[9)L2,VPST2-)O&aIAH.=,^?98K+^2JXGFY3Z@XIY
.Y;BRQ;_#H6WBg(#L]3fA2T(9BI>H+MTA[/76[SF<Q[NYS)b0XWV4S[7S2_b,R=?
<;]&A7?g:)2=:>MdG&C=8@DeGW(T11,g5<W5BYG<(G&;4GVGAKN,U6YNC1:KK:,R
4(2T,S6Y]QZCUKX;>T5FAW0^RFWL)RY_LPY=F,c/#0216R3F.9]X9<C,bR(.g?fX
-S+Of,>L9?R[bNEVG_c6OZ2@/fG6E[A4dJ>U#1Y[CFc?)[MXZ,[WQ^&8PF1AD(#d
OaEY.D=NB@^\Je1MIb0AHO-9\:+b[3Sd13C@g34+E_J:DLKF][N^^=MOK2A[H&fI
N\^3PX&E0;_2NeCC]f@^GGH\9e0V3Z(N11>DL>,_8eQUbT\Z]Cb=>c5SbE7F4<fR
BWNeD<6bb\JR0O<]Ae@5O&C7SUe\O1IKX/-UXG:]3eE-62ZYL<8+FEH5:\-^#+AM
0K]SUG;A;A2fL?/Rdb9V;:@U5[Md?Kac#DKY&//V081D.X:H-OAY55;LZU/Q4?7Q
Q6DK)UZ2=)[O6g#8G.OEPNR3:515<W_FV[T-[Q@#6@Ud/+TD&),3L.NJ3U4B.L6,
J5S0/-W5:^59GfN_<G_AEJ2b:Z,A_B-Ube#Z;+8<@Q?WcG&ec86Oc52Z\B).7<)^
F=KC)(/JM.65,0<c9W9@4S46<)U:;1GDReW@4]W>LZCR,;+cPW/53JA2FA@6KL3,
^/)QG3(e\T0#]GY5.Gae8),N=9DXG-M0@(]@T?YcA,XW5TM11NDe5MQfT):@/,Pe
3=^W\d.gJB9^d,2RR68F.Y,WDfVgOZ;55__</e2GD4E+=NIV@/9aN>G:KO;1MLCA
AT74aPe[bR]d5-Ue3bBYE&C<K[c+?WU.R:OVDcD/SaLK/AW4DJHRLT^a/R:,PV-X
F6B@cK7[a,SY2J5THT._TDJ[0:RE-e?]NE9+gg>g#b+3YMf<CfPKC)Cc^SA++/@a
C_SPCeNN08[C45=cA??&E<[2BWMH[4VbZ?+Lc#D;FCd=1MBd<AfGGCc@g4GWAbFB
BB?+QGI7II/CQ^:fR;]bHNRX_4>/)5)#?bG01CIPZMVOSc)CELK^:eL^Z#M_K27:
g#f#<A?\,E@5:TH6J2+6&PgY;<ZHdNZ(KaN&=4g^D\&&<.gaNSL;IgDKCCLO_[8D
@a#gOHO_54adG121a+^eb?0GC2eSS7g#bLH4_#9CU8T8+/I/cdXH9ee:,YL]XX]8
+?/e+7^eS0T@e4_>&<,Y]bIMR_ZD?<7@6H-5UGLeYG.9H/XbFgRcJ5]1N[@&&0;,
2RG8J]SJK)6U&)FVG-]Ka,P\BgBKNV@[#UVS[T:0\@N.R]X29VC=DaF2=fO7&\_?
<g:N:KU#0Y:T()-DF/Y@4bDAT@NK);#R^V&D:,,dWPKURCXJZ_AOBY862A,fC4RD
_]0/bK(BRH73KX\S&=<-/.Mf<,T[\C,d(8WC?-TD:fa65?79\aIES;UL[\&4,C3S
J2(:SM@M&IGG7?Eb/@UJBWI[c2ME>PY)0&:a6F-dPJ^1H1d.<c0H]:Q_0IDY,#S)
==?TN5.-9>e(,V9O?_dF3.S)_1B>g>_QS:gF,^1O:^N-@G+ILTE6.Je+9>JPR.F&
@[MR=2>UDS]2AcZIUI_eRW.4>Wa.81fTJF26@dT8BL9.Ua>d7O0,O3cZgL,E?)HQ
\F6FIf;#&Q:H/:Y9Db11Z:4Ib-De=9NgbT5A?C77]^fHH<M1V\ec:9^7WF(I0>)[
I4bd_BCTC07V+c/IQGY@T:Q@F?Y15W?CV0IFbKA:06_,,YZ+NE9)SR@DIQCDI;fC
KW#<AR32TH]9+S7+QAVJ>YZ@.HS2AG?eA-f/bb#c;[R-][,DES?DYgP.XJ[BFAb]
N^QD[+5L(>ZI[D+J:@)>7XY/gDW>HT:_2-M0E]4@-1?Tc6Y3Bbd9fD8J/IJaf@G_
EGd.Zc:E7:9GKEc_A\ERd=J^WBM^^I5;S(B:56J@K;>&<XC>U,3cMB[c[b;ID(^O
4MQ+N(]0)_8e0>X6F+7b7#cWL1:JdPS#BA)TP.V/)70?/],(MH@8K-X\97eG?9b<
8L]=O+84]N@H8\SN^ANAO?[P#c-N+f\J.2[8].fc:@RFT?e-^gX>,##HR@-/YCA]
GH8(_f+=>^/#,]b)ME&N99XM/[b>G?Q)HTS2VNV\T-X]:KSJ_L#A8UAHP:8Q[69[
eH0=GU+M^7;)@gaIcYX2[KAV84a-f121G&N:45P4+3D]#QL/0I)@M@.a0HN)O_eR
,LAD;e^Ibf)#fXC?.<5IdYLX3?GISX,PK&UPX?[HUe/:)d0<8A1V[4Q3^J#_._IN
;H+SFM;;S.,J@c5gd7IP611A;I#cDX?6dG4YM/FML;P)gG1]F5COB@bZL(g38A[=
WFH^4?A9/D5NIEPX4O?7D6T\T]UDHR)[Z\/Z9-<I=2C&/>6:?/f&O8CM51A3GA,L
KC\)Jg/N>^bGT]aM5F7W&V0(X<KPM8IIFPC=]0:e\=0cZdg210,DJd]F-)E?c(^P
>AOKT6)_EW7W[Mf^C;QQF]V9SHOJ>U>DN&bZEP6Nc4+UX)9E_I)cVR(FF:4L.?&V
E[aEXY9-PRC>HD6]GN_JAJ8cM,D;fA6#0>L#HDWM=\FWO<J+N\-:b@YZfSdPf.NF
OIg)SZd6L-DLSJZXKWP:afbJC)Va0UeAK@R@X=5^N\c(d8_aI3AX3c/&),P3EPJC
326e-/#C\#W\S?CIIGW+OW:R1fU[^R/?5K1+g?2[//_J_=5Ub\+d2RH8N[37f_b=
0^&R_G\7T1^Le,g6eSWO:EfJb.DM_e8agW#0]ZcQ>G(_VJe&/UB8D2AG](C:G,GK
AB<dQ9/(N^b[+7Pe0EQ>KMD6V;:ZI0@F[#@bQC-D)1;;Ua7YVZ6A>;U9[5A:Nge)
CU=H4dMQ(EZ;_)eIJ>b/YSf@L@PALE1PS=4TK[K.[MY=H@KZVc1\IFPMDW9EL<V]
cE9W/@Gcc^6KO>;)bOAU3]?:1?J.aHYX&Y.1?7)/E?M]@-f=RK9ZXU<>=eIL#KgX
F0\5B;>X?/d5X:cHcCdOd+ER]^H^)Y?g/]>5U/?.A?:/M3#3fK(I^SJ(0#9\,1]b
AZATT&=P?>&X6bB\00Jg)7[BP\+_X\JA]7D0.(ULF;Rac[Z8-M)>9&WQ:HT>/LKa
S3L[E+NFca6[a4B1A(C9LbUE#0e_VO?f=JgFG_;YfgSGD2->-##OaO/1,7LBR@Q2
\G[0LfeBF.UW?6)<TgCWBM,;c;f-C9]IK<?-KRBL(DPNN6.1_O6I\R(?XF4^f>A=
,M1VgB=BOZ55,MN^OTcNO]YP>_gK\g2^6c1E69)-?;>=Sf,87D<73-Y3Pf:ebM^2
1T@N&^BP3IXFLQTH4a/4;]KJF/7TZX4>^N@(:R?9MDf_DM\Q-0fUVFV95\bWg&9&
T9:MO_\&RKcLN-[N=O1S,:Z:?ESID7WVY5.UH>KMBHHE^M,@Rc/;T9fOC\/37T/P
AOX>2N:ce[XF<d2c.KP8X)77LZ?gaPVXaRT9HT-EG]GQ^1N\^.E/3##&-0CZ:d5d
.ID_M&>+JR9-1+KOG:[c#_T;_GADf4J#gLaT+1@D+JUMCG_A.<[H,J-JZJ9H4DdT
5GVcFg5&ZNE>f8KRN1AM,NP4NMDeMf1EJE6.3Q4eYg/?Ff=UXI1V<gC7(]N5E-_\
6<_L@S-H+VgdFC2=5<D9bgR9#G2E1IFc^HI;YK)+(X(F5d@(1SR69BQ1ZJ?ScGV7
9@7F5f6?TH/#?-&[._4DaEKA34W2K)dWH;1UX_VN\ed<&dSDgUVU&N(X<K@^NEY?
cL4eG,_<^FTd^9+NLULZHKVeRfISGBL0TLf/37NB;&Q>#/LPQYHPeE([^I\;1.[D
7fQW2[b>047.55W<H(?,&F6FI_=16@I)6@7g+0Y6Q+7B#_Z)f55?gF5Ue9?FJ<C=
B<S3-9U.bURb3.EO=<4V-=3C)8eN@bbN1AD&W085:C;QQO\d3O9B#97AO/JD@2)a
&,PKS]7>=cdA&U=F95KC9J2eeNX:XRgO5)ULU]D_cH3N24H9Z>V^.=3&1O.MNHOb
.M(2Af&S\gYb(BaSYdb;-Qg&/MXOM7]6^4U6Q^Z>&RA0W,H3/Hf7IgL@(T;5?-+F
+G_I\JPCL11fN865.E+eUMd@Z8eGVA7f,HaI&=6&C3#(3R^/cG.5AF.5TSPJa42T
7Aa<VBOBU:=N@[MZ>&T:Nea:A,.I3:C]U]^\(N4IURA]/],b+].H_b67]bWT3>DJ
X5NWAZOF(U]7=39?7TgL,>U#;C+.V@A:g6Q+]7,H-Y,GK[fC2&^HCW3a_5O-)a(-
<_M&\0ZQ1X,e#]^a:f.L.+^RGMS8FfP-T<5[K;0#2#<BYY,RXV5]((g&aNd2::/\
_J9I)#Vg;gd4/E^R-bL>VY^99WDT7OA,@5<S7e\^).#af[CSB-2(==ceVT7TZ+W)
:Y&,YP24#=3GGG>=-#7Qf7dA+YcgWZ&b7+H?&7(>P5OBL)@3UEe(FP8Td?K:.cQY
5F<N@_VUf6&bgDf2T(;3P9@K1Z)(-CW;DV]:[D7\Q.TPFJc@&IVaDJBEVTO<NXe0
G;;QUCLe2A>;4+M38A#OQa(Q6EQJV_@+K1;@?L<]GV.PRYCN2(DWU4dEJRcSIdVc
YXDF,SdH?e=+,U[4;9#_;WKg7MI5W=[-aJWF1.9(^a>ML)E_JAQ^MR6-^Y:g_\6e
F[+^_fc(R5<3\+2>27^aVVJHF.U-/<g5ZLNT(e#OCEPdQP#683K9;/6Q,RTX56U^
4HT?)LM1C(d.XCV^gLRY[8Id5X?)YR+TTZ@PGc;3a2E7R]cJ:-B-[@TdJ)\IKWTa
b>c0::_ZF0\KF41#:?[WK1#/b,V^PYabCO,H\0_M8NMg47G9T74.bX)2?cP&dA;d
RI#-0BB</5<],Od[HQCZ(Y]RO_0=5<ZP1f_UHg\GY/Fg/-GR(afddL/B;/7Y.4H]
?>bC;5A65Z+[0JGE5=6P^=b.QP:,:NZ3B8,#6@#M8+^IHLXT(M^>@(^L(CM>>Yb3
gP>D;[\ZET@NY=MK9GE-bR#.3bH[LQEKYOL54FZI+GK]Y4c<5@b3SH6gE\b^13FN
2^IS)UYVG[>BO^+0Z+MZJdHQ1<#6gZD[ACP(FW,QLWfQ65)T+:^_gfC>?&7U(MI^
eTWUbbFN(Z\JOF,N;g[e_L[WV,#FWPLHfaH7=ONFP>2(.D>UYAZdK)5\ccQ(eK_8
61#g_#OK&UN17)Z.:S<FBY&9>MR,-(2YJ2G4T7Q^\U_-)gKXaS/KHaL2<ALJ_C<-
EZFV1<-5_I.M:^R^;FRbg\H;,[@a]3P&<]QU;;1V@5d<D6UDgAD)cUc1a1&+1+eM
._4C-TdNYLUJ.F(B\AgS^A??2495+SDJ4g(]4SLTb1dT6^[c<L^6QUNcN?d[fQ3:
?4+WT=V&HTd?[>&QgZ(,T1UF&XU@4\C(HU9A9WK3K2,;0Z+6fJ-9JRaK@PL30W@R
1gWMDQ/[\cSZTJBA]D3&9PM5aBg5+N241\f.ITV0&@0W5db5b?+;G0.S,=M)N9A?
X^fM.KJZKQH#TJKAf3=\O0:d90)&_CSJ]:Y.#O>9P.cdG7M:U_HA/51)LdGK2AUU
>-E:S[8L=e)R8B6L0cd21NDHH_f)^,dO>d_7[:cCFdM50)SET7VX9\ZTERD^G3M5
=EDM?]_&FN7(b:WOUM]Q0Jd0@2Z0:52UOTf@:e7=NOa#XRX:ZM1I[cP5YT5A(g,Z
.\YaTd[fVbd-\:Nd9/T+g5[L67?;^;V-9]_[@dE>49LZ5LR:+D/X:gY_E5NE>Z61
JZEL-8S([7U9V0^X@Z)DK0+;Zff[bg&/N)TCP[2)I#WARAR6LC1,fS+1EeLC>7JG
6Xa0VOX3L=?4NO@#]ZIEW)OM\/f(7C1=DP8FAF^02N^DLFQ5>DGbC@P\@7Q(=-7D
aXY40f+UA7Z\/TA:,\:<I>=TZH]?g#GH-1Mf_<YFC(/,C.F=b0\]<=LZ^F>N+KVI
KOP^AQ3[P)[(6S;7FB)NZ?F<1K1QJfP&)T>#C6PZC2C>EP3L^.#/&HW#),YF-I\2
V&aJ]DBY>V_?UI>5Ea[_JBMTJ9BcQY@>eO/P)@>#Cg,UaD810QP=Y<U_L./YF?[O
T6T0+4RaRP//0:2?H(U\O=,2WX.1NU,gJegK.V4bPd]/gXQA@gH<_135N[9b>/D4
@5(F88&LRYg_)@fb?HISW9B,#RU=K7V8VF+bXS&b@?H79HP.0dPOgF/SN1^O&H[6
5QMPH^=Z@0MDZS>&WC-A;ZEgZee:ed)QR]O77JUZ^Of&9S024.;+Cc5gDJ7d<.K7
IRH0[YY]a0gcTGTM2<86[-#D:YU/6559a@WN:Qe+GCD@WY+HE@75fCNgg?3Cd&bH
d(K[/@Le-)=>c?XQW4U?[4RRA&2KUOH-TQ<SKW6CDa1&RcTI\:J[,A/J/)WDP+.Y
NBAb,5@,c;Idd(],UZ6RZ?GB5CWM0TU1eAL43L)QL&RLc;#P1[18+9;5.gdNZIGG
LM=GeTASP\eE67?BIfg)MHR5V[g^ZQRg&.OC0<FZ#bC&ZM8=L3O:eE.ddSQ.XSUF
7fVJ/cf3G-eB8JA83g^D)]^Tf)fMR#:P;4YN[\8;C_T[6cg6N:8S#<^ecY^QRA05
WD?]X9?-K4G6d3/F=Wg0Z)N97_#/#:6#;E1bgddDVa,&/ScDU2)@eXYH)^aH0(MY
FgIRG50AY-_13.eAQ/1_N/O^:IH;W:cZ]@bU4d/9FU/g7ETTf:]W:-N[N_2DA,]C
<IA5BP9V-63#L11<93B^U\)O,)CSN820TcXXPaP@](Lfd(M.WQ?LJF=LK/Y#g3]c
)D_7=L-,RA;GCa[C0=OBERK=gNR@e]W>PC19,ggeL)8KVN9b/=Sb@Y[NL&Jf=C1,
>\ZD>]05a0-HfZVI;?U?^HeK9@<CTN?I<=:2UD#aW9V(\2E:V7^\e<G/VB5c@ML<
bAcJd\@Xb5g4TeB^eObV>^[CE1MT:3N<#3(M]dM<6HOQMa6V2EfG&2,_#&YJ1R#)
Ng_AH;\#5HW#2bFS8.LO:L&,0.?F8C1=(gRKZ.fQ9+I^]2S#c\DRQgL]M&a6e8G[
4UII<YR1+:XKff[4FCXN)TXdK\d8M-11\g?9FHFH7C6_A6],FT0gUPPP.X=Z/fG:
P4:/:[K=WAU.WLMFXJ5aB3QMT.b<O)c.fNMaaf^Xb=75LT+,d3(#AL7LZOWb??C:
^7EA,6=8R15>gM^22-@J^/J:U7MK0U;TL[]\aI4&QK)J:=V36>6T>):D,HMX6U#S
,^;-F15W=ad7CAg&RB=.</@24MD)?>TJf]Y8(+D_Q8eX&^E==<&L6WA[>TH(e7A.
E?QA6A1HI^COX=3Dd8J/G^>^XAaV:\(R#:JFOKI/F0&8\A(6OQAXT.=(CV\O12:F
)S.>,5)LUFOFea;Q1@Z#=0-IF1dfF3E2<gNZDgP0C)5L@F\D\HI)_+>6)-[b+KB_
GJW]e[<G^AWRU-;7F]/g(\bL@LSN\UK=#5,EBMG@MRY^TP?<4e=[e(.I3_IS/.(f
_gQQW#A^=B,7e7]N@LLAHT1M.@>Jb8cUN:)a=YRV\S7gT2/;,b.M;(-W=V,7S#aY
0f9cI#?VH:XW;HB>>8,[g>;DQV?@e.I7O/XZ[RYR:-;KII-4;]7[MD/b-^B8eL@3
W?_XdEEeZ-:?)?(WZCH24/8ZGO<4?6NE5e6S,Z[dW\[<eKWQM\/F;)AP.S5:\La-
IMYSH(8X[+Y-7b;/37C)5\CS.)2@)S,8J:<UXOFEHP\6LQT82.8C<I:D:dEb]B4F
VRQS5X>eU4;JLP0FLcRDR7C;4E/F-P/\)1/S7W(W0^HE@SRD]>J:,AV3[?/#YB2I
D>4TXa2SGfcD1P+F3G8YBQQ[)210)IX#CO710EH:Mf:\cHQL@5eRDL0,+cQ##(3Y
&W&gRPO?g/)8?+Ed:.BfS:^@4>KM(-IaPYa0I]#JTCeR=&&:J6&5SM/7E=g1BB,A
@6&5K=8+_-;O+BXJ+[JU;6-/9T<:TNC@OQLU;5a]VTCJM#8U3^L31.38)JFP7>5J
gG7>A@QHE3W.@,2O=[9GNJS_B14T;31=?XN#M1^4A<[Z/JAMIf&Z<B7R;7:gU5_:
.c;G4[T\F1P89:HDHWKRLY3&5(S[<2,J7GZU9]9M0dVG\&SIPKbPWfg2[e9O13,[
fZ0dJ\>OR.L[&e(H(KNKEL^[[N?R05)I756b?+0eV,,4^-V-dE^AGZH+2U1N+IK8
L_FI>1:K:Rae1ef>VdB::1<50KIZ/@=VGD0EOKAP3K0b)YeKCGSZJ]D/FfMU/NYF
-3/IV;DK0(@aEK(P14QBH#Z69]&3.0T>?KMG::<JVVD]MI.[GPO2))9T(3&Re>;/
],]b3VDNd0DBFFS;bf-LNT]6K:,4_F1>-C0,Me>d_[1\_4=J9L\Z?S,;]EXR[R6#
afZNGW=Ibc]=3A3@Q7bZc65(NeN&G3PCA[;:WKR7<G2K[b+aYC/@_H5Q^CBK;9UX
T0@0??@gM-:1N<A\88cGSAH33F0EJ4J)SHdE+K\3YS8D3F67a[]L7GR(ZUD-g/?@
HbH&)QRYTd+S)T)3AGcC[=;DRWM06,]3KO&61;:G4Z)gS&];(.e\[#fc2L&8P>10
9g1/>>TMG-L&+B2ITC8.:WfUVY14SaL>fN4N4Kf^]ZZHa;4=M4F;,4ebUM0Y.1/(
bK6DFJ>?EedO&:>(/HI79?MRa1F7+9Aa_44]+5+672^,G<ANbP-g;9[;W6S,[e4V
\3ZAT<4,N8XLZ#1]_<0?P11\f4XegR?7Fb+5LW))0fJLB1;Kg4#c>9I805eeUb1?
a>Y1Z.;g#?4fNHOZ.<(O&[IaW3O5K3P,W)ae@cNMF,[a)WaK)^JQ;UZC()<be((7
Xa>+-:LeT@#NLTYcTcUb]P17I<6&C.OT,VUbNPLUFb_R)GXORbN5=eHeL2-4ZXKY
D??]R5#L-G=<bCAf18a0TI_S1-8GJ?BCY]9b^;+;7HcB/dccP9-Gf[Fb6,\RC];F
X>=51UG<W-NR7@309bSX7PT3_/,.SEO\B<d1g2a)L@XW:<HWSZ7?(1Q-A]Odc\9H
BH2]](;7]CPE+Z4ZNE(LTW+KX>)&KH1OH/?3fDF&S3c3&W]+#Q0>@&OJP]PUd6<9
8>0EB?:d+C;a[S-=[A.=DW6+-C_&GWK4:<7/eKQU9TY)#29dA,X)LXT+Rd:YLeWb
CXXW/&/5/E7OCGUFB5B#AQ4Ca\5\2K1FN>@3ZAdd/TIJB730=V/cG:ZgJfTSYDZK
L5FV(^GgV=DWA&e)7@d[AE>A[H;F4+F^S9d\LAb4=#NSA?,IO(]VUYA-6FF)D,22
)3+LBC3U@\4\Y0^ZRI@Q+fOI,fG=)bWfgR9=P1JTE>]9NfYDN=4\<4ZN3/&S?@;T
:-V#QHXA),:gNA69-E(M&_THN&/+,/JF,_>T.OP0AG:PCQ:WC-BY-?6UPgMV)[QU
cfZK3f4NcR#dL6RE:E8]X1=2>5,VKL/&?;YJ1?3[b#.&a]7,AS=SVWNP4AcF)8ZH
.M<\ZdL,36c?W8^N&L3;Dc.#EYIE9P-[(1g?M#]/)HgZQBaU[FT_^a_gg&AcS0:-
B]LH=<]Za&PR,0@deg8]GOJAL_K=GD)C92AS+cOe.g+1<1bU3^aUbZ3Z>UO89@:U
&5#^+G1;Yd\K<O;G=E?a@B5/B;=)^W1@#>&aQXe#10QNM4L4DKER7B5?<1FA9TXD
=gMU22X:(gR4G(UUP5D,X@#ef]_PPbO3X:[,O3fMAV2g@MF<;M.K/C4e4+M#OfTH
O,feY=_K#:ZM0KQH3NY>d:<,G&P=,#c50L7U?WABO8X]LWTL6K[\#]gY(5UG?Wbb
.VUcW)Mdc_]\<L<.bNQ>0)S>2VDNY;S;G8<L[YJe5Rf:_:?Xd770VL?FR#YdV6Q7
:]77B0RHGZ6a6D^LW92bb(e2H]&B7:?@H8QE-5C6B#W<6P4K(M6EU&GDP]GY40QS
XZU7\E0c^Ig(=[T0/0&,U?g-AH=JGB._QHP.aLdSdK@/OE,DfdH&7B>^&8Y_)LU8
bb-f)Cb,c4Y,VK_C@6=&N7_<^.BeD\?_B#^Y@S>RZ;deNXBC[[R=RXB01D?Xg3@M
?2ETGaI]WM[S9O.d?KS?c,J+>g(bNS_83_3CHg:6.#4OOUT1bJcYRYf@dGcG>af9
@=0-41Q)J6Y]>Be4/8O=KeddA.24:S)M=EDM#(S8M1>Q9A4Eg\8JA8J7:J<b\1c[
M2dBBFKDUgQ.:eY1GJ<R_aP(SZ>P9^WfD8Ee3#()e3HN+.09J-<5P6g\Q/W(0X\4
;G_V?A7]b(ME]c:C?YeV2KGZJ_7\D(39((7(f2D7S\]4R_BLT2+EB=KDd=^fL@Nd
,LY9-TU=fU/5PUEO-<EB=98[>XD@LT:/8A0V8JG[K>^&Q55R2fCeW^a^CQT]dA3:
/MaJTZ[&b0e_JC/]MG/>]26^RfA(bB;b[@/RC1,K.G:fXO&,UDcKI064--;L^<>+
(=PA]DO<;FBN[0[a;?O@?eRX0][=L2/AZ<R?]eXV(X@U>M3H^?@Sd\E?/@8F\AKF
:LIWZNZG^c/_MYb[)U[P\L&4WFdI81?+X&NXf#53f2O0>cEPfKf1JK^0#ISXIcG;
9:&V?0H=RH<K:a+e92.?GUgLMSIGT.AGE8b<ZR52=\Zc[-B0,;1E(HN7-+;S?6O.
@G_f6McNNQcS>;;6(RB6g4cR&VBR^D<(9ARHX3@@RO#-=)K/.0>+.9TDcec^(RYZ
:/@9f3>=N0cUbF2):IU.K:2ATT:#g>4@dKCL_af&)E@R>>R7+4=O+\PFCcSE.F31
Aa.[6WS_?RM6_A,/-@MI_3^;O+EPY@G#.>59.gbX4+]N>]@g]1WM2CLPJW,AB]-]
VFXfT6KK[P_b7eKdD8,IP/2@UK1fT_#7J#Mb,Qc[Vf(YH&&DN(;-&Gb^AAS[^T?;
K+M3f_0.<2#RM@>^b-0f1,L)Q9NI3#>O/G6/P4_:7cNZWKJ_/b#&NRDK&=NVe^e>
:.d8M;.^OEFQbMP^(fQ&N<Y6:D<bSNK_BVVdc<A66/FcC.24fD:0b4><aWRJe)E8
U_AaW\^/G&@4W<1UgV/QF:J1:N48L4XVR],M_N)VA5FD1PB[6Xe9ZQ5YW:SZ)f.b
1NGR(fDY+129J/3]LPH[8(9YBSc/S4OBAg5D<KR(:HbZ[EZ&<JWX?0]@_SZ1.=LN
gU51bS<^,S_3(Nc0HWZL]W_2[3>bNgUH0b/[RPRb4XB#J(_=<gO8g;X-6(_6STS(
F?GL78T:d7Pga2eJKL]BUee@=6ddR9C&H-XB-B3#1FGZ[e6dTP@F,U7LW=)H?]EH
9O1TdI.EEA]Nc<Ya0;4QaIaZbA,Pg,<^0dA/IO6TfQ2.K]DR4.b]RK2C,LOL.7RQ
HT6<F&D(FdD9c5<(:a6;K7daR;FVXSW6XcF,^(C)+F#.H@,/I7ag7>X#f<U4?,:b
RDHb#ACd9\CIPV5<.CW(#LJdX?E@.:;dF<;TeKO,]5D=0HB18JS5.0F1=HbMOEf-
8R66TD/24?/(.E)^G>>2EH.R=G>6/b.;dC[1>DH:[^Kg4d5EY_+e+g6^(F4IdKWP
V4RUM14NG6cMHUF=e=V-^e/_TMd]K12WKRJ5+;[5[S?NV(&@2feFT9126>-6^XZR
H9,N)=.H3J::AU7Q(A]Qa>],,JKHL,a_19:XQ7c_MTW<G3bd39KdFES^LcQ^H)F4
O;GRVH[4cR@P@LHQD4..F.5C(AP?]:\XDR#?Y[dK^E-^.[YM/QOZ2O:D?NJ<D(\B
Lffa4@(=]/EYMR@P10^]KcbAPSa/4J4Jf25M+U.WVNf462/Q;2X]#cO@7DPBXg(#
4YMW:ZAG(b,fJ=&G#]N7J01bRV\bD2L+,6PAZY&U8(11Xf+28A,]\Jf>(3.\GN@(
AA0GbT(bE-TH#2&6&-,HFJ6X=<:9c8QMZA[5ffXD=IeX>Q,OK,TJ.ZY\T\NU+V45
KVbKHa,M@80T8EIe)gLLW]C<eH&^JFP\0[>Ua(bJ]RC<RG33Sf#[AWda.ET?)e\4
6W+9TBA/f@B5gNA_2&C_[6R=Xc0&X1#5XTQ(gSE/eDODf6^#U1UMV-&:;FX+YT-(
7UT/NG>1PH-IIX9.IKJ(_[>UgZ#E-,7A>f)^1<ID5.>OG_fLFV4T8?53&VXe?,>:
T#E>9g/XHNIP^WNX8L?MDHPIS?3.ZYZVe+)^@5)e/4H.#0Cd4M,Qfb(2ZVW@+;G9
J(e\EG><4]4O52dfIO-A@.#Gf)addFO,B:=e#8&1<RMg]P3f,&d(>&^//X59d9FU
>N[UG[^8[W-+7_PO\QLB5IPaIa-ZP1Y(-##(X]G3DeRgXg#3?.KQd)Pf;7O8gU;6
DX7B7B(WX&I\-@_@g\GOE&=B;1CCWN]b1>&\2R;C/9OEXPTJF+UNX;/=S#R[2<.\
O.g\W5A)9T.5;MK,N#5MfeR&UHTQNRe5Ce8A7NVN/cBc.,9W)I?d\1Rb(:P.2ANW
3HL;WQPVL[V8OL?I/_5AV8_P2OPFGU9]8<AY#\H^DI=T;/UAVF12C^V^).8JPeZO
Q/398P)8I#M20a:SP:/aafYNdKWU;2\3\8a6(YQ6^;LR[b:\+1,?BOf&g=+-d()b
7F9A#6]TL\I?;7f&BJ,NCCe?g0WLZ98(7\K/^]TRH0cMP)^f#NJK@7MEJQc,@e\&
MTc[@SQOZF?546NBO]6L]I/g),));/R:?;FN-OW(gRBX6=C.T8+&.AK0MR74QC+;
^aa8RJYb#gb/a^6b;=8eHX2TPVZMB27?0]^=20dcdd&d2Q:09.W#bb\a>7,JMHe5
c88d5f3S<73:<e4H_.UeAJbaBCM&bN9c.N0M#77@46>)R9]Kcg&cJ01b.a@f#<+g
M+T&D.@X=C]WGC.cEC_@^H5-S&J/)RFW)OeR3P605A6J/)K?g((YNZ&:Z:=&DF,W
6]f/DB5_Eca6ZH;)f)X@R;6>geMaY-MXIJG4<[aP\:^O@&:dJA3dL1(_2Vd\QR)B
3>+XE6VB@)3M^D+K_KUd&LRa_<ZG+M5>7a+@RM/F^_O<+6(ALgG\R1f@FF-H7]<Q
f?D=]1/+MTY)FTV6[V.2b_@C3)#Fa;TJX+D&NbdJLH(JI;;MIJg_;.SE[;7d^BA5
LJB?GYdE=c7eUgSZgSW5;c[RHYB6C/K]eJ\2[/B?1NCcO-Ua_WXWWB1/GQH34C<_
EV@3f)a_EO\R)8MW1A6?MAg<=Bd^d@QKXM1e+K4&T#M(5XT9=)GcGL-_)6IIc,\,
#2:27?QT2_?e&]ece;EQ#077Ecc@XX3(/<Xb6\<[Mf:N3NFR85//P>f:W_TW^5Vc
,.1e/SRKX?O=F9E\-&ac03Q8FVf\#8K(bYO(OfJ7QGD7;J271HN?.^a&G^CeS_&:
a5:HE?Aa-4fC4A#cIVQR21Q^0XLP7C+>)FLX6ZCTfB?_C6+H@=_ZLS[G)D\FKMN7
CeX51DMP7]/C)Pa,VX[Z<Z4,OI#H/(/8HA)/NJN(8K>LYTB&9JGCKW90/:LB9ZfC
5.6e)<fUGP[e1E.:[J\I(F1B4gEI9&/gC-NSGUUcLL^#cHTHLUeSD?&H5W^KAN2?
0b#D<eHZU8M,:YFGH]L+T^_?U8-TZGd@:<&DZ-bBOSZ_>cTH9<0A6FJB3f0:&?[9
?+B#TIa1e>W4R]=[F&U((C_&-Ce\7W\)3b5<24M3D+V,.S/>d./##-\UOVOMRaBK
?/71#G9Wf,.;Z[V_dEF@LdJY&WB[8:F=U-.Db&P<g&+O=YXG;8[HHAZg])#UZ&I/
O&0?;?(gS8#R/I#X7,9AAeJ8f#>ZTV7BQ6QdNHb]b0LMIUSg\EU/?0_764,]8B\>
OH.9D)UE#G_Z^RgI4@P#c\O0(2ef>QFUT:gF>;[,CSbU#/6ECa[8V&ScWWGO-L7+
^KM0Y,+c+Scb?d;7G9DDC?Q=OW[Rc,E;?2,gd@.bEA?7GGU<#.21-,][BI=)YX7(
G:ddd@E/,L]#PUfV3dG.aJQ)ZP32N?NN26dU\eHEb+JQ6Z>.1:H\Q\cT@B45G6LD
)dF./4&^.BAJ:.H_<_AT;:VaQY@UI//U.&c27Le-KG&c:#O&.KTRBGN>U+C8(6IC
JX[eR&?+f,L+cD]U@4gF(IV?3L4A8Ae)@5C+X[6LeWP#Z+MS<_e6(^)1J([6SHII
eF80QO/SCddT7H-0KSDbHaV?8$
`endprotected
      

`protected
5>F^dB5FEU,9[&)7JWRLR7T>1@9YGR8ZFEEH;6G+#LRe/>F2b[I@/)&NfJX82.(c
F/2E]97;f+/Y8/a^Y:J:EG6D=SA]VJT1L2WKG(^IRaQ6U(E?<9&aHT^0ST:#/L^0
_&/[C_dS(HK0_>NP76>;69TU/T/O2#I2GafMY_F1SG(4H9>I5aY<:.MS/MU\1-:Q
#E3>c(,>JX66T\YXEOBX3L>g1OO?J=Ne)C:aB:SU@:\da#:ZS84]40P6bOdJeH+]
(/bUgYJC/=:YNNb6/(DNEI9M.3&93)a+DJ=3Ca90We;)+/&995g(SYI/>#_bJ_+&
fa0&c4,9.^.N)^L><OJ)_PWE4G1FH:U3A6<W5KHZg>IW]eTKO8:9=JQ/@:G&T@SQ
;ZD+6@XY1XDTHVMV>+gX<+75HVM1g6Y)>T:;2T@\fAPK)3f,9TLAWIb.(d+7)#N(
SK?NHe)+T:E9)Z+E68I@[,]bV>LE+3E-_Mc(VY=aVg+UJ]#b@NYQgKgG[FP@[FA2
K0@_<AD_^<?P5G74B74-QLYD)Q):W^67G-81)4IEPJQ5Q\K\=f;eKNO/Z3U#<DWb
##M@M9\gbdP+b)LR#\#F-_f4RcKf]#UL=$
`endprotected

//vcs_vip_protect      
`protected
/QA98-Q]58:b0GSA@J7cJH[]LX^\1>1]=cTNM2ZMF.TDec0SBA5^&(#+b(B:Ybb,
J<(XA2/-)a(EWGe-:S)>6\#I=U[M?/beK@e4N1.a=Pg?f4H^++1Z<GT9Hc/IEIV/
Af:6Dd^D6O6H9/[NMED\MQa+HY>OeRKZTIHWR9^W-<\TS(2B6f:O@Ie8@K[5R(?+
Y]^W?6UMWCE.)GONX6&\^-U7H?L+E7aON5_)ZO^4(<2ANPg4gZ(RF>4<BX;bIfaB
C;Yd@80fg]&E&U,0GZY+Z(R8;6c8L_WTa)MQ-8L\:40REZRC(dFKH[&CcAZEP5_X
R;(T3E#9<FPf,T4K>5-Qc/fAg;f)0J&@>ScEXaF/>(40A(]c#3b@EA+\2MdPJ4c]
QY5;Y96MJGf-(dZH@9e>)(M@gF7UQ=@).66;eBQZ(I-)N-=C24OXIA8M4[0?EN2T
^FL<PI/caCSgB;?=&69[Jf@C:Ua-Cb,#R_3ZY6/gD&H7DSb3)64J@dZ/ebDB08GT
,P]e:T/_PYI[(62A(>0I&DRb[Q7EN2<Y;#YU4<DRP1V-]8_9><\_K-3d^I6M\DCE
U7eJc0N=CA[7Y]2+ad7+\:WZHe1^WRQaYV6:JIa]<c1d-5T?:B#(LJ0:91FVWSOJ
GZHZWSf]T-WA+e[#G4I>;]>8&6>E0PXB&BbDQWVH\=,S.?+Y9g#T7g=-5;H3699A
\W-0Q+bN>]2g=7-6^\)I50fV>QD.3U-.f:0O&1VRP^Pa_(cLS3(<-R(e2#PeN=5,
&g&]e]K\R)L9#O4HA;#BCa74=L#XS\VUW1K;54e/9F64A67LHT<eL??K-6]+,cCM
<E:IAecP##d4].Z:&g,(cb746$
`endprotected
      

`protected
?UV:19AY(\2W(e,H.I1T7DB.Q?0G:WX>FYXW7,RQ?/fB(Y-QJgfJ))870:W@7e2Y
M@a2GF(/21<>&G9?L8^57dB.8$
`endprotected


//vcs_vip_protect
`protected
:T_>HDU>([OBVO,,293DZK4@U]6SS(ga\69PcN5Z?@D3&[5#bf(D&(9OH@JZ2\,d
2,O@fN6@A[SbbU_g_<DGVS)[T6\9b&b[,,LM9+H3&3^C-;^0)GG_0dG@b2.)]f<K
#KI06\@FF/Hb[SCO3b8A4JEECN#/^U6a9Kaf(6Rb\1HbBHW^L4G[Y-KDIDY,UYG)
\;U3f4(@^f//;dSb,6A>A1JKeH\K:Af7#DEZ8C^]BU-IRM_/2.M8g<3\M9(4E+>d
<baDbR8BSQN?;A.0,#;9(1CXg.ddX7C2GZUKU>HRHZ/\]LfWR^a<JQ&c0dc.Xb=E
7M(^/BTQ#g-(O-@:LeZI\PZa@g2<W00=W]PY=-SG1fXS-0)/&PAZ(dNWJV4);GP=
D>Od23E,QA1L(>7DXKIP8^QaD#4]/A][=bc))A/7EZ:PfV32;=gREcUUO_\8GEBN
R;?Qd-H&LYfQ,=9@8<C3=gc#GI4D0>OT=+R<\>VZL6XP49(D?;:0>K[PgDUM#6,U
Ad8.GE2XO(9[PEJ>^W^<0>CJ3BB1<-cF_QWFE;N3;];a?Z#O)DWB@3)9A5U@<#K4
ZQ6:>DAF&_@,9+Jgc@#VJdWF;#_.L3F/J2.DDN_;QbWC_-Gd6aYG^F9dHCL6e+FZ
72))&F\=fYV;I?XDR:6WY_:>R]&KSD&J#efK/IQTKd771KgUX;K35cJ;bccME8cb
EV/N&fE.K/#\\MT\,6g]d)YVZRg0T)@:<Mb<B@E(N9f@QLDO3:^)B5>589<U^>AC
YW(^.K<F]#XV4030@=g5JH2J^_(+;5M[9HA6,bU\d>H)&>bPYePd,Z[HH2PYQ7I7
03WO]V&=[cQ:77AGMBU<Mb(/X:B.PZY(Q0S.#+RM<g/5#&+<YYMHGUe6NZ1?XU-F
6SIY>[_016C90H-;39R[[?c>CZ69Z7Xb?ZM,X-JgN3_=.ZO\_?Q-?MG57UOXDQb;
f7(TfJDWN#LK0IJL_TMAV96E<9;b)]&+Sd8I=C[dBA,Z01eN>:gFF2(MR5WNKL[B
.+,S@IO)UP0fNI)FQIa.?_X:V-2:.LGWY>g2IZLa3_2,]bK^^O.@N_)Z\(a/TKE7
Z1[2GXDE2:S[]QBJWS4>3XgIa1#7gNHUa@]R5(;Ta,->)?6E+2c#A[?IA8XM\0FB
,,RHdSVL9GLc-dFT8&J^U_a69CgG&(;-DYfRVf#G_f.47.;=ZID?,F/LJDVb@Z[0
++UG.ac6SB,)D3SgQKZdOIe9V=+4;CT)&f-\,&BT/5:OeYCP/7I81OP]I3.<D2<J
[_E4J_64_E,PAQWVgKW6M.bZ3<]EV1@-P+O@/Fd@\+SLJU).#_Zg3b.]WCc:B_[V
]I-UL86D;V+TZ_VYB9KaGdJ?C:>4::KE4^]K]J<1P1I3G1(P\#CN0<+H6(QgI6JV
2H/8JSDO304\bY(_cU0ZgWcCMJP^ZG[7XA9IUNf_^]XUF[(^eI<#7=6UE,3V-,3;
.NbBW1:]0&-NFX;J7&ZZ:P,?8Z:2_eQ.0dSGS<^^#(g]4DfF7BP^F_>)(KH1E@9X
Mb20C[N0:2[HGT0O\?&R]WgONa5ed(b/gf\f8=e51BNYFIHIc(O#(LJX8&@:^\;P
cB).Q2H#=Y^KD49Ug]TL94H40D26FGLDaG2gHWfZ^(5KM=YLa@WNG&WX78Lb7/\+
AS]fH0DHO0A\a6VP_YbJf5G5AE&/L////b@RBJNd^^,Y@I0UfVOP78JYd3KF3^-.
cY+=A2P4;b;N6+@AT1_7V@PH-Z?,NWXWZc^L6O0G6(AM=2+LOY.)Da=<TfRU29/W
NC9#dY15;gF-_?Pe[3>?3])0)&CACUag9.Te4E:#=WJg5@_/Y#S2YX[_/>\9RI9f
e6?#f>2e;HF_(P[ORLKV?Y+f#75/56<A_:;@F0b(IP0I>-G2Ig._]=8dd[/Y:]b@
^\2);H<(7N\K]fDV)T-P6\4_DYGTTPWEU7AI[=D\/Y0f0_e^[V?Kf@M5F:VA6Y@)
1[G^Ibe:?N/8d^,5[7C5K.Q/3_4a]0D78b=HVV8708[,HD#J3T-)4PZJ;87N44.\
gEG41e+]6,;9],T7^(<LgLX@^)I=91^XWS5eWY6J+,A^Y5eC&P]&N/7N,)&T7I>&
LIGF=TZ-fO7VDF#+@^84Z9cIJ2_9:acOF2X06Pf[(IRS9(eP504(-DdDf]U=:NgM
:68_UeZ(:B3T-aYN^GB(U5cYf5EVSJT9FF9#F1+3]+>V1YM[R&;#GX_a74;K5,\Y
Tf5WHV+-Sd)TNM6NS8,acZ(R65YM_<6T];?L&U)#]TeJH1U_._^[RSSIAS0Y^&c@
1:<VT6@D]K4V.E_cB<FE;)EDZZeSXD2T^D(N&O38.C1N+8=KO:H(2b<>TCGfJ@eJ
QL\M0QHbP34;ffP\=J(b>T63+c;Y],Zd14fEAH0JUMc-)eN9^65:713P(M/eWf)-
TdK+TN?fR+b;:I[6WH&AeHNSC0[BLKdgTRF<fC,:SLMF]M)F1<Q(I0W(U;@<be?[
SJE&8].X-0[I=b7Q.\8UG+LS8=7YCBC1LA>0VC1IgK6^+_RAAV<=&8SA(T.5?>SH
aRA_AVJ&\M+-05d?cb.VH<.9TeVMQSS3YDN/<7-MIG0_W?\VJX?(&&=J^R>JZ3Sa
+D(37_W/0F5[N,&<5I05+,d>TUKJK?\\KaQ[5L;KY69__WN.>f_&S#6X.U_Lb8T9
TYBO3SgVX2WA\.agT-TRdKZ^f9:9I:Y9&+?)6^7-MA#T,2@=H4>O.UB6]K1bMMRM
G2>d-5^6IGe<MSa/c<?4^]7(5SQO]1PUc16;8e[DA.-2G+_WN2PTc0c8LYJ@^/B2
&IC\</4d[MEg>?5)M8;9)VVA-+f7\P6Y>afQE6NNE-6,C,WPVf)1b-=,U@^N6EWR
_(bc@AG83.5<>9UBa8Z??PZ:,IS_]Qa_GW/X@dJe=)C4e6W=2TH9/^5^4A+:TL/H
WdU\M4XCWGO9D<>cA\42V6dX(B_dBd-fVE/8FW/ab#KM#H=.DWe6CUS#\\L2ZAaH
=EQ@eH0RMZY>R4TD03c[6^b>JAb1#gaNVg#,-d]E0<^.3fN]U:f(3?dI2YbJO]U&
@]S[)P(.(T=8,H&U@2H.TTX5VWc\ZR)Y96/=\2QR/3,aCM\0MOO3e<AL)\dG;=W?
Q:TM@)7/+FT[=LR(<fXcMJb-S=VS5>X]bfO;SDQ13;R4.GKZ@B3OfO<c,PZeCG/_
4aUGL9Y=b+Ja+8U,:4Gfe43+VG4MDGSINI>CTW0V66=(cXgG5d8GE^,7d3=QSC1:
Ze#^LT8@fbg&._DH&PE/+fDIMP4(OWQ003N7<E^ebF]O;]8g0F/c^T[cORR<3T:(
]6U#ZZ=.e,5e2R;\I\NPJ9XEG_3UD[76T?6Iag[NCd?YF))W-ccY@JIR\[gR>D]S
.=)N0ZHODgd2gUX-W/:),b?X=)adHWd=GYNef^/<O)6\?]\T;X&GLB96M<OI&OJ2
ZAP2SPHCG#;OZaO4Y>>dO<AaTY[9C\XE&3><_0L+]/)+c4HI#=aHJ>UUYUZXXd1P
T#MPZ2W-Z^85?@HXFb8=1V5P@E#6RfAPV?1W<dT)G;e7]#d/>[L.__XN,Xe_N^N4
YI+=g(]B[9NAcPb7dJEJG)eSHH@\EaY7BJA;-E3@AS8:.0;eBcBZaWT>g+?#L3B(
BVX/F6.F7L1-/3A=bCTC7F&4YgD=2\L<]3LCD=PYZK<(]LF/FIcCcdgKQ5>b;KP<
&QcUPA/02-;E)0WJ^F<Ha,3=[NGg=7A[)TdSDBeTg]O(d_4,\+FH6@Va[Qe2bTLN
S3<]O>^L+0V6[10@,-HBQc1U8Y73RH-(<8fNBG9D[e-X.)BBBD&]WVYfP]TaFS..
/D:9L;1UY6SU-.O+(R?2Rdc=b+(\R)3Ya]IRD2E&c8bPD<Q99J#0:H^>YR[.=T7R
D6Q]9^U2;XLS[,NC/+-G&HQA:(gGgaY>AH5D>=\:M3SEELa+^U^.Z0_U567S@97G
O/SR,KY^U)XHKNA_NYN)OJb[-&(@gT?USS6b8K:[-/K;AaQ\^6A<,Q[T6]O4J(ZZ
eHc/bN_YQ^^+W<X&85M#QXT0GaI//UH)_Bg_eV[V>MIIfg?)7N2Z+9<T;4RIa<,P
?N<3T4O#AcgY=A7L6T((-HJ091KB0eAI[EQ)R;1T?@G8,1JN#K/O693bHK_Z+7QO
=SR:?gB/Q7:DQCKU<@2@R;:75TZUQL&+UQPHOg^A70>1HY:+)D/7(HZM>ZZQ(Z==
?^/V_#W+Y8e\IEW>6b<WdZ6LL[;YU]f[.H;QOZQ?BN^Uc[9,MBM6Z^P.[WCYE<#/
G[SSZ9K=/:HV,/]#LR50YgDJ-Ic-TL6TSd@2gL3.AAbV-:K.T1fc6+XSNT711S?d
C<NM&fdGHWf?VMB7193=AJ+@.B=ZYT:-?B](a:3ZG[2QVTE5=44-Eg(J0O?Y38R#
Z);_b]TB+=7d>B.G2F,gaR6M5&dSQ72Y4K-c5R7gd.gf6.F<DZY#XgaXI]+eMIRe
XG<^4UTM:b(5,Vad@YV^L1Nc_b3OO3KR^7]RT=/MXW#+Fe37)++;OeBO85-B@LE8
/50C1/)E[MV9fA1L0]DCH@@5PU?/JOZUBA4Y\/0YII:=B;U6cbV(a2.ZP7+Q9f]5
eET3=#;Ae99Re#.<8HeT@C[6_W3)4>d5(&U:I6#+-B@c8[48P&P+eE9-KVIOZ?\C
]22W\4YbOB@]4CdT=<Y<Z-,2FaBLg(6>J@a+=]fb&C2D39bI>N5LM3;K.A,5f:O(
U[FY\N1=FU>&_,gMDg1.Q(;]L<E+9W17@0Q0aE18Q)#J81DRN)O&b(2K<G.\VWI[
c9PcC=I9cQ:A(AZZ<YUD3,gNIW=W_1>9XKG]C-PLT)9\-]C\+5:IG07L0c(2\E4.
1&D;XZG1[]FIEVDA+VF^+:b+/WK2QD4)5\;DZc@b@L-T#LMQ[I-Gb<>4#4fc6J7J
6.(UK4FfW84=6()0\2S<9=TL@Kg<Sfe]GS(LN0e&/WQ\;U25?(5EXDd&FUY4V<<S
R@#_B\5N_L(+>RaAI=H=0:]TK;1EF#Md;8EQ;QGAS@MFMV;Ea2(G5<8O^gJXRDQ8
bc^cRV<16TYK?#KDC2[53R.V+5Ec:gaKLeTY(-@]0^#]7I89S6,82:,fPUZ(T>e.
<F7HL676>Qe[ZDMV2G_HRDUR[#T2_DCT>\ebFg7B?Pg/OEGW^BNP[JLgO,dd.UgE
JY]O&Ee^W#Ad^]0BHa/EQ/]#0:?6/@NO4DJf[OPVfD&cGQCOd??:VH4&B5<&9Y_5
K2Z:eHJ>RFV;^DbO1@J>bf^8]E=D\?=5fcdD_BL>=LZJ>0UQ_gc8K5[g8Bd#?FC+
)3FE(2U&?Gb5I=3+_M:J^:E:bKMOW>cM-eT]-G9DIJ4]U^H0W)7U7HOL^g:43UEA
cN\B=N+UWUgd-FJeM_e[]:AdZ25#N>:X;4PgHW(N8RJe0Cf\),5^2M8OX=0<4U&1
[&cb3@R]B;-3>aT5M/:L[UBeAI7PK0JY])57C3VOH+a1^L0JYc[EE/K<&]VgBH)5
C8XF,b)8&9J5a</YWGFI:Y?X2T.]<dG8>N#@MP_MSO91_Cg1@?gV2]FLU?1-BW1=
93He8>4:F6,.S>_O_^W)CJH3MgXF5L5K^?FL9WY8Rc@K]=G3Z#;[&QC,4R<gcWKQ
-UdDCU0:6agAZ.3BZOO8C9bJD^#/:B/3,;T_7bHR[)03D5:7f+</G[_=JG^Df_KI
^-fZVe-(Z^<)>:#1Ja\91\&bgH(e8Nb<4:KHA74eWR\.@89XXD-b3@-Wf(.Y+:]]
1Y0YM;XGa9<9#O,;@,UI.FSc5UF/-[LaK9(T?FLa.1\2dW-F<A),60YM6;:Zg:W5
.c.(WY-D30LZdGL;\W@=;Re<UCG-@[4Y@=M\H]<:f3S2KE^Ka7V#ZbHAME</?(O?
9)9,9Na?N-]8(a1SQ@e_0a=bL:We._b-L_2_F@0,<-=6g3\cF@+?YUaK)E8dgAQW
]gF\9>?)/aX+8Se6DM)RU<CJ=6CL^Lbb7dRZ?Cf^e[&7(JA06f[O0\OY5EdM-R#B
TI)02XMW_G:6LP5S:\(_9R5X0C=cS@Oec931Z9S)G9@<Z7_A#+f374+()TWAS&_0
O^F60A+>.2==G&Q0g#&/AVFT35DK5g/.Qf/RHaWU&)_>NXCa9BPgWUC#L=^d^B0e
X#W(GRW9-D44DJI9e-,9M8FcSLLC+R;_38F;IB3U@DJJ\WE2G(5GJ(/e]\R4TP?U
R/[^_E:D>;ZMQQ_;>/5.[JR0=dTL+L\VdTC5d,,aH-A^IXU?b<U/K3?-A91\FBYB
]f]c9B>[/J:fa,V+I[>\VP6Ya)S)>,0BX:5f=W.1ef?B;W8[ZfK7I+R^KfWQCK8>
4O6a>A4-Q(,<>QgbL^g>[4<ZT(#;cOMaD529FE]V9A]Z=8+:<;0JS\\?gXS)g?7G
f46=R\BE30:HFL=/I=Tc5EVX\.c.+>_R5_2(G9]f&BHJ/W371[>XW9Z6LA>Y?LUS
fJ57E4XgCId6V(^>#D(A-D?&a(2O5O=BaFZINd6EXeaTW7VKcEXc>^<BUM=5#S<_
:3-S1S]J:>&9^2XNgJM#)cBaF?9>Pa7AV[,J(K.)CH\CY9ZNgG_:BeeU<XW2C6^g
b><6?(#@<)02a[f:GO5<6;FO#:)>@-bTNLV\>9TQgGad.RJF=CFBYW.3-fE@Md6A
YgfP6KOEHWe20=d2e+C?6V@2=I1DA9/T1&4:2E>C&?F2RGZCcdcT>[YSVcB#8FVa
.2#0V^BFFDe,g7_]I.=@:;UdGRF+ZW(?ZWB[RNIUb:>01C>eFRf/J(F?1;O8A66a
d,50&>D+aK_5Ag3L/[9f)@/S0^PN1#_a/>)ALK.&6MEPQb(\C4KR^BKR,+,7,gX?
\.@:T(8TKM?X[_DH64#K;_93a4@N(2WgH\AG7/P16MGWIL4HE2M>:2E\GQ8,)6:I
e07O^IIc=CdWI.ag,2JZG7S?g;R<b7JQKCNB^A@/,.N@^dR71(]2FJEY/SR1b6QB
M=VNTFc=aQUOCTCeLQd]@_e3Nc7bL2cANfKI<>\\UMG@RK=/f+G/9SBR6J<KZ(Rb
T_Y:J&#ZSF(?#(GN#=\;c@#g)X104W2>>I^fM0\..a))F:/T\)]?d+>I_eN7]e(f
4ZUT/4bcPEXT7?dd&8L>N)K4Qa,5g-1DY1Sf.,.c]RY(8FYSD(72;[U\758]0TQK
_a-BK[d>Pb\#+>3TG>E->U_A7E[7b(c1(;KF&K_DA:f.I]cS>;_:V6O]c#O:2.WO
TMKUB-^\U&DZPfKLE2K+)P.G1HH]BM<:[7UDUM]&\;)4ZINbc;ZQUVEMBfGF2OQL
g8>U)fb,UFIP/,;8[E0b9&GJWGK[69/dFOUAReU3N&-]N[510W>T3NE:L\+Ad>G^
#B^cQR7B6DW+60)FO0?N1f+NVZ#6KI/F2#L?ecagcS.P5SGXdMg,N[^H2TA#(S:9
.:03(:F2V=U2WD/)&]4O5R+OG(fce)5/=1&+GSG])WZ@C+(^Fg#1]I[06W\XN+Q@
UbSW=Jf/O8P,_AANbFBY3W4=]b<c;&,Q/]K#70b_S(B7<UJ3e=0;WT()G(^g(#5J
aTM^/fT^#ReC6DXS,DKMS?PW-[?E\.W+fHF,YMGgaGb-[>1#dH=]I/MTD:4PBZAR
HV-W+RH;+KeM?4]RWgJ,/-]>+^-d83UHR1b+SKX0\FB5TV7W)2ZX.;8K,T\D8GP)
cXM7.:7)6d2^)NNYRX9(]fAf78EMf9JH=?GPR]<=E(5KC&+bI/f)d.C0Rd:W\47.
7PgS?H8#1@(KYMD5QYN9AL0&e3UbfMMF(g[YAPD<GAcNW)M&AAH]]cAfGd0N8M;f
#_(:Z]+Ac<gJ1J;^IBO;&B==+YYEHCQ1OcHb6\:bgZPW:OYD/)7\O^>XD2THQ#I/
E\R^C_ZD9+VE?4VE8+I,U[6TWE6-/<9DNb01P26OF?4X5HHEKXOQ.VcZ7X+=_50S
V#SUc;5H:&RE5g4,SOLZ8U\G.HQ>,fY&^>2SKAa>Z&6\I>6J3cBeCTX>;TY^T>Z[
XJ@RW\-6GO(JODM0e,2=AWFb),Rg[YI6E@;^W(M,-HCc:eX_W/W))(TUYN-KJd?Q
B=CFfbTd9X)8Y7c_4#Q<C1KH_AEPNSZfI_SU?DOaW\fR6,AL5GNXe[\A96/1-\f4
L\F[](:M#X,?,0=c6JF]XO;a3TSAW3FB.@0J^X9\5RU96H^F.E_A/BdZP[JRPCc1
_)4-eHcH:\\80-KH&>A1=5fVU3C:5AWAPICHI8(&^_g80@<bARNM?@]_YdAbCd&J
K,R[b6)HR,;2cQEZ#gK,Re[^@UCMM4^@OFb8Wd5+FV,LHG1#f&A9D/P\+5?U\+-B
VLORE^ON4WKcEdabU3Ke0XOddfI=FXKg10&A#EPKCg8=7Y.W:bW&cb\X:/WOE\c&
OFd+.TA16N\IaVNXR34A)_CF01YT8e(3@/17\XC7)Og\.?cZ@0R5?f2\A^dC87N^
>C0bYO+KQH-W8.71\bT#D.8#f[>DD.^c6]YfB\>7f&/YN@^&cQU0+,J@K=V;ZNK(
X7(b5CD)\E#Le9J5f;U#HTeY^f0G4E2cU88<2JQ>?T0;9c2C<BUfF=D/Y7JH1XY>
4V1W1.V-d0ead,KXOd,5G.Q?[7=7?EN8.KE-_cFg8RA/,\J5/#Cbd]J?AM7TRWT;
5U_>2W-/1GGDK&-?OX?DYV@)S1.70eF&M1-gADc?.#>b0=#7UMDc/NcE6N]X#B8#
2ca&+)TP<faRVZIPSb)ELI&V[(a2SV0DCKNg8BGK3HBe.B#0?M9;)b,.ITV<f:2[
CAPU1<Z+Q[G4M-gd=];cT-X;YNW-+/0S_L<bSR7;\aY3Y\@X[<W8B7E?389Bb-MK
0Ha6<AG0RcN.HWCg(3]ZSY.ZTZU6,@N(Zf4OG5cWJG;9#L>4AC0MFX_Og:eTOdcM
_/Q442Z5[1--2&M-]^QKLSFPS-LRZY@]TbE#;U5[71I<XU=Kf<GC@5HRJ+g@6g3>
W@6F(0X(fDF4?Q_egJLHG;1](#>Y95XOL+HeUX(&G,\H&L+]ZVI=ZBNW=\IWgT]L
K;WfcbIfc^WVHUS?PEHcG;IE:H1)CE)a4d\;CTE)7+67UXOHE#(gLeZ;)Z=WE,H^
T65F8B[X00U@DbeQSJDQc227:<8&O>c+C=PR:IIGE^O:J#C6I5N9;-+f\91TP_e/
EaagXR54270DCBJQUW5^6&-0)]NF6UF?X8W?QU##WG7a<I,WJ(8>X<I1e&C\E-1B
c43I1O#XCUd4^,\KUSNGRGFf4=2Y1Xf.fAc#,(a3&)8)BXGP-R#3_/ZH<gE.]Bg9
)SFeV6=G.K?,(T;@V#Cb<82?>V3>Lg+H+]Z<=9RFEfY(1U1XR?2YYN?:Z2]GIX#/
Q;3)(+U2f^#Se?=a^aFW+@8E=JEME83ZA7\,BJ\1=^DAC-&f]@]EK,g6CS,g)U/Y
L4dP;\M.1U;PAGR=0,KD[7Ne<FbVY6:VVSHN/=dN)@L[V[H-Xde\87O8A?1c:Na1
B8)>Ua/Wbb1;0)V#\UWE@H0ZT,;2BPXI.<Pb.5()g]@3c8Q\5>T\V30.W3I)fXdC
X/;_LPM-;GA2(;9O#,e>@gdfTW.cG;SS1USA8KU.A:/cH/3EdC159aeT,d>RIP3c
5XfB\\U)HMbNAY:^S@5N=S[\^5_HJN#d>18]UVYe^2R.D15<DZd1aV3V(9Cg1S)\
a00e0#/E5,8^_c_36:AFMaZ\+@9CN]_G-M]YAD7c?WfH7G2ZNL@L5AUH6dD5dJ\T
(H9LQ-f-4]G+8&;<RCc?UCJc8)gQ&UI8(<JfQFYHS64LKK1_6=J=Y7e+a)edJDA-
3T:<&/O@)bO5J762gJeRY7@-Y(T,PSe+MM;>b4&c0<5]@DT?7O]#F843Ka@^HI/a
:H3:9NQ8DVT)OQ=:WVJPGfUP2Qb<F6L/32E0V2[3#/TCK9E#-;:JQe?51eS](8>R
BI7ecLD\T)61b/\6SP;d+3daH?Jgb>AN/3L7E[FQFa)96Q<MebW0#QD+3C&eUP+N
/8[dcV&S_EP?#H&#.L[Jfg3)HR<f@#B@YgJSQ/7GQ6W4.K[6g^&&S@a-#3]\aJ9B
C1gMEWP#\RFG5N/=e[3VLgUXedYQ(&[8S(.)Ia6;c0?>&EB-F5aC29WW8,U<MQC>
M>&EUC:5>5,NQ/:>bDa@)0VRe&<0CF(>@4@a;=VOFBS/85gC<C>W(4b,W.U_aD;M
IG<(XGIV\SM:1=IP2e53e<1L6I&)E#4H@_6+>660YLX/YHf7VQ5Cc[C(6ZSfNTXd
?6JN@L4V[gF-?7TOCR3aG-L.8K86AV9.Xe=_BM_SYdff7I?9ZNFMbD?J_=8(#IDN
@1Y.^7<.]?.1K+(4LAXZ]EOJA,(Q2[].4W(NH_g:;edWYF[cKWXDc4@:>O4?8A6I
&AFc@Hc[.+5Q9,<^U;BKST9JN6S9AUHUY/<5I4=eD/-^PT8O^@->2>eBLBO3><1H
=8M2a-R:fZZ(VY@8<X<)bO(]T9V?J,A?7:+B@7AP:<:+eN)]QS(YIX>MSAa4XOcc
NNBX@B9?39-<Cd#BNE[4\,JaGM=(<8+FGN0/;S6KKHHa?AUR&bG7F1QZ5E/d3Db=
U&-Y+G[#bbHU)IS76-A]?Q4I(13G+,I&Rc=9EG6O)=4,aW[;Se2X6:XKeX&P<SK)
FH0#.UDHU]/,gfAHfb0I9LWE2>L/AOXBOUQbX:E6//@aXUUPD]ZPW_cZXA1Q<R[7
\#X\K]:]d_EBFgL\4XN_6?LX>B.0-\KPEPQH\DbNdf):_H-P[JFT?[<Q-C_0XNSG
C0;H9[YNJb1DZ4?>MM\I]PISE7SBbW<P6<SO2&\1.PIb#N9MD^a2FU#SCY:7ef2b
KJAgYYU.QOC=?+cQ<J0^NVbS9W[bf;SYRCMGgLXK<5PNcLS8eL<6a8:+^)C[a?,]
UPXPYeE-:;;58K/<e+I?W3KK/;B.^Q(F.3I\96/)VQ+cf\eA1cWBBQaDN93@-\^H
ZL]e_W+7f^bf0b1\3?Ua:(WS)3WNV_P8@R:c.&Q1d53VA_5HW<HWZ-TF@UWYg>++
eF.9:P(X5,3g<IMfML]a]>\73?eB1d87XS1QKFeLESDcbEOgG+>GR2NO-;&aG]bH
e>.+\SW:5#<<2eI-W03NM[079Gb]M33E1\G(2VV8V5+Q\?>c@PSA?#fX[6VAP>Q(
(,M<0D]Ga1W]#WOaf[O97g#2cQN^I[&M)4=V&=W_TCG#d<GZ\5.Y64Q;aWV\c0/@
D8[3cEVb7bF2J#?@JC-HP,VSNKa+-dQ-LO_4I<bJdbM)b3[1#L1/5&\=-U;-PPG+
>+@;\RXb+G8+3LDZ)\Zgf(^J4-8:]@(fb=5]O<\3QQQL?Ze5\D\#1A=W-S#NgT>7
WJ3-.LDW6[PFP:46\G2cFAf:E^>#YH1YcWcc<)f4;5f^Z1X)1LU1&USGF-O+.@,f
-IXY[<]8DLVV:-&&(,J^WN+VfH\&V5NZ0H]RMJaEOd8GI]Ue_F@dfK;]a--\<L,=
GKeLHLeK/[KHdSCF-PY:S]aNaRX]8UMHDW.\A(M(Z2MK^^HT>__JHY>2c39WBG2L
C0T0/FGe;_F?TF9ND1>[a1>M30(N5.K0+Rb7J[/Jd=-5\&[#?M]5fWTKM=J,;+70
K&8^McC+IO_GS3+T,THfQ_YM9GLJC[]>B:.A+0MaDI;3b?9]/dbL9];,<]^T1cd?
(\4^AZgR)Z4@f?]._#S/bO#b]A448H-Jc>/I.C32c12^7FeIDHH-QIc[@4DZXV5O
6,ZJJRF&RVbOBPYT@I[[f9OgZF+5,Y=?@W,RT=_PM>2\8)KQPf81G@AMF\U2^2;S
JJ0D9E^PQ2EVRMbO/E8IV](EBS4DTUF?>M3_]_2^5a.UMBgb0=XGB?dAJH:W<)8@
;5WTEZUFXd8f:<Z5g0E]S7@4-3GbT4[dG[.EGNN#;[UQGU6+/I=H;JS_:C^]=O>L
[58SRD.7M050AIZYb253bO8WMA5S,e;KSfGK&9_W;I5FfC<a2E4U0-[88\a[OD)O
FU2?bDV;ITP^GUAe58e2Kb44QU8(fg@P/KA:G,Mc1[Id;&UR&4;\KWKH^7A7^UD6
(;PQK[4]Q@[A92(/PX54(cP+:_A]MV[;35.?.AbgWTB=GQcD)6.?QXD1g;cR+5,G
d=\BNU:AaVfB>@Ag]79;9Sg/9/_QEc4c:M86e+T[9:7(],cAQ0GcMHN[Y)9C60B,
b;5C#1]KYR1S,RaA1g4<c<UTGWIKR3>U/U)2WS9Ub:)[S6&DTD5-SL5V5_b60bL8
-L9EYIbGT3@]85gR/]WEQ7S\H0R[]HQV-]#.IPAK061(0QcJ/0eBO1WEL+:+:8D?
NQYfUGG09X.deDII/J4/R\T?B+e5_@eJS]gVMCc=NG-M_\^0\C]dW>WW?b,V=g6e
2(;BdL05=UC2bIOeI]SJNaVT8a[BKOGg\R<<><&2RX#7b4@bQcg[8<eAMJC3B0NF
DE)R6^:/YFY&<a>XgEYW)._+_cT,c;/HZg9d35D)[RT#(BP+]fNP)NZLIIdgG+E3
TfV7F-Z>X4W./bG1;Y9NN0_0C9>CWZa9EV:Q(=/PT:/.RW:L93Y&CL3KG=1VO)BG
94TPFG^U,;ebg9\IP^@M(.>B0(XL[I7Va6(=AG)5V,A8>f(X:TB@/-e.]+DdQ>bH
UH=bIUgL8O;=J;(7ZICe(O>?A,6\CLCQ>=8g,P@KS;,C2+.QIF)NPa1c09UTWJZE
MHX117(7U1_(g^-)RV7I<)#2f&Kb#XXU\O9O8ASf:J;[J2c#.PXMX8HE>g@0P&VI
)>,?]>+>D5a4_[S=N]&)TL/,:Y=)/5>-<<H3R4UMBC_])B@57]/H&[O)J<_&O:=c
_4<+Y_&^.Y]7GSfgRLf8L8f<GU<00/)5C?KBG7U/O/b;51f-XA?:\SR:df_8bcDF
+/8Ua8f.(EaV,g<^36Tc(?VN-3W1)f#_-cN:&@;F4.XI0-EVdGgceX8PVRDLOOZK
>dH[AL6M#(M1)&/@DVA&8XCRM;V82.fPbFLfIO@Q1b5faZ(Vd;BOgE,.RJY2Z?PQ
/1@>dQ_18,CfC@>GCQ/cXQK6\3LZEf=3[XO7fA.P7)U&:(>BB,Z@#\/J,U:4_S=0
ZGYd6[D1_=adM?KY.HP:&ON7JO:V+4GMA54135@VB1#1BBH#?1I[JE.)4c7=)gLR
,7P9(H:JO7cXP[N[a4Dc568ZJH>,2Ce5Oab3=agaHD[X+37e2aG5(_AU@L1MDBWW
UV;.KVZ2MS>6Z>VF;bU\RH8)<6KW;6OSMGD1Q/]LcWB^IfE+f)a;HKQQNMfNOGEO
B9M2PR=N)TX3fT;U.I5XNXBf[Z/?VUJ]H?4[bC;;Dg^cP@,JQ4ZS1f7.HEW(Z7L0
eR(EIJRTXMDYH-EYAGGZ8L79JUG5?A:W-#5I1++IF8\\_UQaSEXPKFgG\,T)GW.L
SL@)\E\....gS9)OeG:BA5Rbe1D8=&JZaP9&C440DNcOLBM);;[&+:ZB@S=CD]1A
L+V^CHYS0S7-Y.Y_Y#GBX?Pc:_OGY1;cUb9YE;7f0SGR\Y>7;?OAYJNV)/W.JB//
RE7Q6/B@I)[g/KQUY(OHa(1<FNLJS4P@f:Z9B#KYJ+N>:egH+MK0b-_Vg28-LEZc
QX<6<8M>KG?)JF67+Q-Q:+NAD)(=a.UcR8S;2EYLAf#\>[]VZDY\+(P^NY:/CNV5
LOKcD1@JJc]13);e86HQ:2e#&2e>R7^_+aaH+d>^:eBKB.60U58Ef\2>28,Eg4^+
T(5cB:5.UQ/fOS^MWWV63B&E-JFE+e_X_Qa0LLd)L=b61Q+UER(W02M#OL05<5]I
TFY-T;FB)>A@>3Mb+eKH\9&M06AE^&_a/]G]AQNNBFRD3EDAa(D#H8S)NP=.9LW;
E^AN[#620H)]5/IGB=)=L;5T+dYNIVX6BQ#Z)\7(cJD\(><X5YCISSd)1f=C]Od=
2Ec,KPcXJ&+BQ1YgJDJSB.Z3MF#bf9M&9;@HJ7CB=5/Z>>:WYK1U]KZ?4L(<<5gB
bMb@ASD^gWQ]+VgY6_,D//\R=6<L9W57?22)@=C<89MDKDDI?&=fbNO_O7bg7BS4
?ZC4eMTCXZEWe6?^dBF&]&9^-+CIf;Sc(8@a1(da^^\3b?d9#8b/_U>5+RGAG.f-
;0?CN&)M6NI=HeA1XeNMe/J^fY2QL3N&/X56-13#g1X;ZD-#Y_H1Qc?RaG)\<:[B
8K/^6J:X3_g.E?D-GWB-Q+#YJLW6g^,;6Z,c5]V\Y+1MM-GaE/YLbf_G\b(e2PUY
(9(:@f_Q#VVa_&\bA&gR-@K8]g9M/#KeP>7?]WNV@=PO8d;d3OcGS>a_bHP3-)@#
1A5:K8?61X<XFLW)F)=#dN^B:D#(WM<E\Mf_LG;4KfK75?-1\)CJY9S)Q5#g1N#K
[f/RIJ5A-g(OU4WU\:LO++[GGVR;VYdOM8X4)TDbA+(X:K&09.(IBZ=(>WHFa50@
Lb06)BAK-0aEY>UD:M3E./=?Pf)+?0bM067<XIQ>XO&/TP8SIN@>-_Sg,<Q5D9X=
<ee9/C_//:5I;=U9C7K,d[IT_A_dS\W3+YeK4aYWFUK^B\/1U3/(PUQQ0;.b7Q>b
HXQ^TD:,@X3>63A/3Y;YD:7P-d]agAYNH@WA4EL(^d/^RO?.3>N->/R,,^SY83#V
R8I.DQX11<V?,S8Y77d)g4ZICEHVXA\HF^)V72.6:X<#=W[@,Y#a_#3b#)LP/;J5
=>BcC=gb.?.+<U<Z[&62O60<P2)G-&R4TS?O:,7Wc<SfW+&#M;(a^,JN237@K0]Z
PNJR4>XCB&[RUL[+Sdf@^N+]T@7\/(d8.Vf29^Z04a92CLPU[2e?#,?G,&De/3X0
2MG?X^1_c^T=^U&Z=OP>TFQ?d6?^^36^bW8FEK66/DC3(4T99I3WfAK9,L_E\@XQ
N^;:,JDIOQJD.4<BHAbf=>3c4Z)cS-0S:GAc02CO4H#QR,1QY-N5[[<Q63L;d]9U
b,b(DO=bAN7A[=#9YB,#U9U.[XULNgJ,\=O)4QU(MSb&b?I#]Q^[Cd;X0R0)J&1a
5DZ@f?H3ND;:MSd/SM-dPXB3ZT@e,.dBg_._:-f0-;999/Aca5._V<7P<0.CW5&4
ZC89?ETRG/1?AP?L,1OJ\VG>1K?\JT-@4d-NS._YXA.NSR7T3NgREb5[#:;PG4QQ
CN7Z,TZLe(>P[C,9VJ9AXPE/XM?eY3;eF?;\=B7XPDc7T8a/20<<K=..-P6IQe-H
_)WUKT6=V(^/Ie;@\9VC^F8@S;S@8A\4gYP-3<JXY21<,d7.g:,]+HB1JN.9F\3F
Be[^JMRW:09KEYA-[69&USRa#R,cD.TD9,3H-W-K<+Uc@16^R1]O:]_&/;D)CRYE
Rf4L6aQG:.RYbU#__._X1/UYf7D:VMa40[DN3?<N_X2+cD&H[0@:8@c&G?&8U&_N
25=D=;bW5QJ8]#5_-ZW>a\EaP5_]ZfZ1F.gI(NK_-7EbN#J82SU-@X;(fL8e(Lf\
d.b_Y)[8VEfaW>Q3A@@=d5fDg_>I\DFCb?@bTAG:8#QKN+ZEP24#A[a)B<g\AH9g
34963/3+dg4OI]Z/IRVW;^CddH?Ia9Y;<OQRb4@.Z\=J5TFf8bJggI3X3K,:ObE_
-&AE@26Y#4,@;=fVE1(GG\]LDf>C\WPOccf\<Pa]]M4OL)<TNVCS/Ge2Fe3TgI3M
6J,]fE9R]?+\SQI##;CLE/)Y0cCfRE(\_G4+[FRQ6#2/dVgA/5bDDLB>Y,PI.C(e
[#?C3B;L^4[Xf2A/g>g5bW#0c-d+L-1FIAd.5f7#FR@aTELB27]=f<Se;XE6YS6Y
<<2NZ4eg6Z0:2Sg.=J84-O0&4a>6.WAM45P\)@[.KH=S,.HCIW#]RU2fU5g:UXF2
(U-9>cgg60@I26,IW)RY]X\bESDXAHG)agOL:1\Ed+B=?^c6^?MfCI#Ce;)#g\E\
ALd@S7+)GdKYW;7JZ;)SA([g-TP:/-.5dM\X-E42b<5^YM7?__-S1=<L&d8PW#@,
]DJ73#aC),KQ;#EO:T+e7N>Dg_5Q,b<cH_-cA;JD&PD>RKMab6OB@Oc)S3eQX\6?
PN9TG^3+?O[N/E0PV8fU2N,Z_#bP#9]SO[=b32R.E6)J94S#8/G=89\OK6PSQ^9,
3U4LdSMK8>K:;F.9c^?c>?d6V,Sf^48KY+LM#IY/@M9[B92&Q@NO6HYPg\-9:_2D
4A/]cGb_?S+TAEZOLEDX.-_\#(RMK>f\^?5_L3S)PV+:D9W5:2-Q@ZO@f(38aL)8
bB)RY[LIV3+>;2WaS<-G3-7L^cR&#\aEc1Q.0,S<(JY?ESb_Zg-Q/CYXd>eaGUH#
?\SS.3Jg6Y/D:Z5FZ)(,#>Z+#^WSER+c@M-60G]04>21cDS#g+VJ[[]+,7A=V,LZ
\RYW#78SQ1.CdZ9B[R66JMG3<6<[3(J;C:d?R6ZIW3@Y&(Z&QU]&a0LMg:/A&f]0
)+[Ae]CCaAgNc_583@+?_B03=LbKMBD<Jf6)_b3<OM@Td)=HATVSMAB3P:?\aG;T
WeN;>#6G?a6Va7ZC4)_0UGDAQQ/SS.cA73UGef5CHTdQT85DINF@IYMQW&::]A/:
-V)B(VEE#9,A+dLR5&N&R9=5QF.?=Pe:_]b;;#Gc5X<a2:G/:SV/<E];[8.P7W&W
DD92[IK,2RUM6c0GC0O+KdSc)&W:[??eMO+AFgY([[Xg\Z:\TV[?QZ3<^=(<T&JO
PBD>4[b0;/G^YH[c8>M2/SGW+TgFW;\?WfFT,4Q<9^_#3KFS5U93L67UeDb5;NA<
59WQ_=b:BQ@<8P0cMedYFZFA^FW]G45ZM+1UAcT.KVe,X)&WG^@U_:+)+ZS7L9B@
]a7W_#)OILR1<WaPe=#<c4#dPTT3O(E\M=]VAD=a-LdJSgR.\gO30@DA9^<^U^Ff
,Ve>?1&)FG;)P+OX36=+^IGMG=ff1&IJH,=dIa:]WJ_@[YEIZ/?LbL9Z:a5+[LTJ
5V6D7#e^@;OJV.R(DeLXScbN7JN7F2X?6UNd#ZSH0:FaL6\0WYH1g=&@B@^NAQ0X
:fR-+2KaPf27,G/.3af:8Kd4ISBcYHP4cd&HIfIMRI:<O^EbEdXH0A]QgL3cI@eN
+-)H1A&NV>2PS\4Wga]Wfe:L#ffGA]AC1IC#W).HZ/f\b.HU\UQDf8Y_N(5(:=(>
XH7PKLJUP4[A?Qfb\X6dY7O&<ZAX2P\(EBc&&9fW;Me,/2H).08\?,?88@F2b9(;
U[NI:.B;A_&=d66KacF+.O.9g7U<;M[QcNf33QBf9B6FQ/AdL=J0C,7:aDNU(aFH
#Z=39d0?S:FS^X[eKgBc@KK&B0(aAO.XUIW6Q:-P-<,BGPRGY_D0<VgQJU1XfZ=c
,R6/Lc()AIB^gG@CS<ZXQHY]OS[[BP-<X2<^UV7XPN&\3?d@Ye4EKI:Z^KWaET[5
XWPc]8.PRA?R-eIO00H/#214&[;_d^C?#aT6Y,gJ54:YN9#(P,b_cV4K<<RI[.\#
]-]WGYc.;B7@a,7_(;W0Q[A7I)S/E@FV^d?)L]&fEKdgX2VRBD7c?O(3(PF/2^4D
gVEAW2JXK[=,4++B2DI7b;Z(3_)A\@SGF2<I&cW9(+]4T6132ISZ@FP#FfY_S-.Q
F^OffRQLYW>ac\.NN;ZF/)[LTEF)+,C+[3;@OELNR2eY,JI@:23IG5KB;<);6]4B
]6MS;U)Bb-d4F9b+PLSCJ(MeMebcH@9^7gC5_QON:_FO16:09.)D&e2E1cXK9]^>
FUI,<Ha2e;K^V(^)T(bC9&dPDC==)+8bf#HZ@b@;-/7YQ/O6GJ6>^T//J+#K8HL.
:(,,Dg_KNWI3ER65^(0D:<]BZbL@:;/1X4-@R[TKf^g][-UcV0gL^MQ(=+4N?]EG
7?G\(be2-Q[LE7CB[W<\4b@(E6Q6cg(1Fb\Y?1dS.Hb?S35d,eZ=eE@.=H3+EU5:
fXL_4RMN5IEU-GJ-0?e/Y^?S9_[+?G498WSH:H^)a66Mg#Ve[-@8#\#bJ68\LGHU
=S5LE<&c6JHK)2IL=D.AgZ7K>UMO)#VT1)W/R)]e<G^83394d;WP+fUf1M<a;d3A
A?gP??8]G1cCF1=1Hg^LbcfgcF\?V5Q/L(THafI+Ba[U^aC1,cWfNZXAPXDQ[9-X
UNaC<]8Sf/+/,&3@fM8S3aD;--4:DC7a&eS?R-AO?<bb[W+U,;\ZZ448VEN72=HS
T_M<M>IB<&=D(O(TUOI&aL[::@65/IF-8>24@3Q.@N_XUX+LDU]7K]4_&fSEVD+V
@dLM3\X]g;C0;1bdC/FGIS_V\([Y-CdV3B?KWJW_#+.gJIc_/LS>)SDW0/E_3I-M
G?EG5R4--03H:6BL92=XN&:T[Q<<#L^@6DRDTa#eNN^dW4M,RdH&44X]<1,4NFLC
V(I6bdSTWSc2B-B<]8N-C(8^9bD=X#S=#_&HK48McPE8EJA]F@UGN?<4Ae[MU8+g
EH\DKR(&KeAgX(d^@]8eQV7e9I;S2.4057UA_(HGI_bUWS\2-:B.2L+7^.-^Z8\K
TdZW-&[TcOXZ3Cba5Q8:?@E)-f4=GeJ5a,XD@dSG[<C:d##7M;K6SD,+IFdXCa[F
C]DTEJ?98G9gI^?)^S5<]8M4e#aKHRQJfPaSfM]:1dE:PZBA;,#eU?)H,O9/5YVS
F7b?.)U/C>UO@I.<fE.TRLT4G0@?9?[-=/FKWbgH5:RCdKHdeBU<;/QNJ3S8V0N2
KXfW?LEO48(<CM]-YN;/;[GS?XW(8DWPe4g(M^a=K)GE=N4.<Z3RL6a+WC5]7E/f
BGL-<Q#@(3M;F:7ZdSEV.e^?^.AO-=G806MGI]OFSL@>E<KA0>HB3gZf:C?\FRcF
G8(5>-KM-HN=2CGXH[\.^M39[-.CK7gQ_f?4BY8/MGc49=RNZ73-&1T[:FHG]<e=
?,b-WCGT,I[ZcV8_HeTKT).\CR@6M:BOg\E2=@AJD8)HGV\^=<+6GaRM-VbW4a[D
06[fHX&TC/U)JT9cd:)JKLEOJdQB1(aS_P=GdVQCOd7UT8;32T427Ncd2XKV>NCI
UdBV&I745QHA>/UWB7d2=&E=>WKB]6#IM#4\f]7=;Ff?I+\D14R27A/@Tc(;<KCC
AfY?Z0^T8?GNA.?6)U<=#,O&aOYH17)]>5<+@a/#_HKY8CQ1/.KSbfTMdbgGXgV&
9W:VAIAZKg_^EI6,V_ag6aI?RNCA;-(9F//D2L<BZ/4J?(_MY;bYNTR,V7?Jdc1.
g1>J8I:#7A##P>da9VTF4Ue/B.a/-UY-=3GfW-dP^:?W[f60Eg?\4)#7T3Y04C/)
1Y>C^Ha<7Lg1495JcK0E@T1X]L[-8;MUbU^g\c\T#gdEPAaJ.cfOYS>+FMDDg@/;
?XM,BQM-dWd)/EI9;O+b72ODaEKHJP\g@@+L@Z\)3G@bPFP([(,@TKK(E7Y3+cXY
c:O0b+W7b/a1Y4cS&\5?65_WL1c<,Cg@1P2@Y?9?TCGBPOc&[[OXJe1P&=^>dYC.
4#5bcf]CQ9WU7L+CX6+AF>[P^O=SKSN>>7#dFPB:=b-/W&GaOG,W#aO)7.&M4+FR
L_I_PX0J34/5^9=1/B+7_)8b@GZ()].[\:Ud)(^15WX61^DF,3I=DAf(>C3^TF#5
]S]f-)F1Z.=))6J?EPdWAAMM,a/66IU]0UB)8AV>a<P=B#2bZadE:&;3<>=8P0;J
,,^K+O)?Rc(dLXQ:X4>I@0[>fRA:K0KQ]c6@Dg6WabL1\<eWWA;VUIMB/fE:)O5.
_N\C9+M7K0M8,JDD&_H4<&8/F_>eCE(W@2QDZK-QKU4RU5.>RE_AM=aUPbLgN<T2
c3V0N]FO242fFD.I7;W9+33)a=Q2IGbR7e15+gLTWa8C<]Q8OY:JI-U\-A89F6M.
78TgL9EESG&_9)#9&5-)0,4_Y-b#b<CeF9[BMX19H/5;gMQYKe.8F/SG-5.aQKF#
HS&Sf1<#Lc7_+D:,.<2JYgP)=QgCePfORGR9O0Hegg<>;9<(J]S6JNc38,^;D@=,
V+D^.V0Z7X(@9\9D-CBSX1:9O)#6DYHDA-_dX/_cg#K;(:0&fZ1K@0=cHfIZQ28B
V>d5GfM+VALB5ON6Se_NWNLT1S+]6<-CI(1C^53A6aT=[?cJ&&FXW?6N4CC(ISTO
AOAfeZRVee>RAGQQ[L>GGJDAI((RU6J<R<C>T;;(.J_G3E:(MFc27]\37Ee/&_;H
T>@1OI/,FX\YM>aVc,c<H^_MXXa>^0e#;d-PNPD84H4F;].93DWNQNIJ7a2&;Z/R
JUeN<]WK;52X,9ZQBgeFH]FP#2^89#I0@^7/>7C(,Q;6,AGZ&:b+<&/8B.5<DW[(
?]]4&SQ+G5)YR&O1OaQ]CIY2T,B?@EEAM(&WEg=4X;FUaaS<HT?8S=3^6@KI1W,g
G7fEc>).Jg664L#W@A:7_>RJO#G/],:3C@>W:<ZSO(31#,YR/[C#K]>CP-c@=;Ia
HQ#aLE8K]J?4LdCgO,g,U]G+LX\@>,IN#7#EeR),4d(R#R(I67JYM/B=-f.04V./
^B,[bT13DY84,5&MV2N;CW/ZS3fX8cR?\3;F.;2,eCRZc8^-E]3GT(WE@.NGH69Q
:]&;X<_J(RI,&.C.PK0BR#aVD>4Ed99A?f.Ha<CMb;a.1eg952VD_@HNEI+9[[-@
)K^cGdWf^H\.&dWS6Ia93e?A<dJV&,4T@b81c1+aO9Y&P(1&1bKM,709C>Pe0.I#
?Fg2M=GK,\OY1BbJ6D#HD4R-5TN1^g;DX0EB3E#,a[BX<ab3eF2dV8?5CU#M-IF)
=/,30,HcdO>]VRGYD=]]/(#V?E-Y-E/gARQfXPMSY7)/CZ3KeebeIDb8)P)^^7TY
9N.Z]R+ZYV3WFDP]4/:2T]gR[IM:<g@-@Qg5;UYe9Z#L)--@#6@GF,^,9a/\O8df
C9]7U1XQ1]&791YI&Z&;?).+VPW=U92QV@71,,9&Cg-HG4.W(1WOa9gMEL4BLYf;
0>:Xg9^4W2bOB?=S/:K>:e>=-g1\P<EPQ#>WA7d;TQcZK]T_8VU2,I[\&XO=P[_@
WV(<JQJ6b]^1T7A:D6>]#:eWBFK;=.]@H5N+W92R2K@-=P&,9-2ZCCMc/BJ58@g+
ZY1.A(R9&EgN/^EM6ODbE-:NLW+V91;GgYbD0)JW&&MLOJ8b93P0_>,)V(M9\9B;
:,Be#,g:L8NG?P^L]/ZAA/^7E;6P^&\-dK)#=V6>EAJ[4BOE0BMEG=/d13&<\A@T
K#L\?;M41(+1P@6HAW<S@#>XEU<_GJCa&K9AY>@DKY1/C^MRa<d0VI&D8V:]FEFJ
=BE&1HVT:>+0/F;6?Lc6,N/EYD[1W@GF<K>],+b31:MS3b#04@3V]J7eWF;SKSaL
-BTBER,-g^U0g8=c;Y2W3>gL/.2P.P\@_+\3E^60(acTC[PHNaSP=(Af]7X<?PB5
W8(_7NN8T3/B2JIKEaEKO<VTHeg_V)d4)<V;KIPZ#QPZG&7[J-Ld]>>7-<_UHf,#
.^DfcO.(fLKTP5>aUYG7P[NTG-V[+5E-K<6?2N8(=3A4+4O1.KaK3K4-1MOQAd#J
6#U);H/1SUPHVC/:cXA9TM]3S5=13.2?F:^&\35e5:b+F)TQ(W2<(Qf5&7;8\W:W
:Ng5.L/_ZB#SC=9D#JY#)\P@C?59>?T;R:V@MPILHc.^BYC&PA.F<(cZg&K#XM4J
-5X7_YC0cB5T66YPP#5Y5V800]O:H^-(>^Q+46MC;N70CLJ5XFffaR</d;Q]J#O\
ZNU;E2MW@MW^_O4S\D#X#]T4EE4M;CP7<+9=L(69f+PLbg?0X?cOTQ42JE@QaI/7
d_DL[I#9-d@DLb=@0BL+(/<ZHI-f@SM6>-5[GW#ZE,0c=6>gUNYRX0&O=\0-5LEI
T+]@cFU+a25@1FYYO]V,(e9Rd]MR;1:P[2C)VS0)8P],>,;ZPb1cN0+0cJ]V0#U2
WNK,SCJ+aEK(6D6-CAHdZO7\a6-EbTN066eG]]CV2HK@S[32E.M(CM\#[E\#<(F@
PT[6(VH?;?W+L.ZN\d2HHd4S(#<cdI8L:P4]7=4c#62FPFJM7NfQ,-Y975b(+?cP
YKPG>\MY?-&RG+>O]?E&5AZgaSD_L?YGIO[U2_-#EYOc#3;AfU17Q1[,PG43U5+8
1(V>5(908:.9?7TT<;X719XY#CFQ:;_^^V=N3QN(]a.@>\]1\KIE=<4C/9Mb5N]Q
Pc>^8c]I>P>aPNJ<LT?7ZH?78&&b^&PQaO<bTY_bLLN(>Q)XDS_C<dBX]V)^R@M_
?Z9Y;g=DCM_U5TPO,.I]74[BBNF,8L-d,&X3;g_4KWENS;[/G<Na)F97TV+XGHLR
FM:IEH;=(f1UWfKKB;4Z]Wa@ZY=9:/9.Reda^+L((=UeQW2#4dLQJ3J,=ga2ONEP
C-PS?+U^<\e2)VR?PJ-5=)S<DANL]6BS>CcL]3G=KLX4<3aXfafO24=JcK1Uf1Q1
^O;QU_SQ,,MH\AQX.KF2=&LC)>&+L@D1#4-DL_-WSgGcTMeOaV/5L;I)H.M3GCCS
G(Y<-=4Y#UG<,O0P<HW.LG:KI(BI2?7/b^G]2Nd2>W><Zb0:L85)-N]>PKA..9/A
OSaH,H/H6T?-/afA(L3H></.RYW+F_Jg3?a;ND56CM3Y0P9GbJDE606ZScNV\MCN
cSYKFUH#3_:&4/T&SSP#6dNB>_QM4944fFU7FV&#X/.T&,9DcUg0<GHLQ1,:2)@W
PD7^&f3dLWR(fR4U<TD\ZUIXL=C<2RaLMgBDg,@MfJPSEb4LM7ZO:J#M7&4DB65A
JZ<VEE0ZUfW=8HKSNB73EN]cH&_=Bg^g;6\DRB6Xc:A;,7CJ)\MNcK#B)NUdfd5H
S<E8M[F[+.K>W&SK[Q0gZ/Sb/9&8OaX7>L47M0?QZR_?9/,ARQ)Z6CJc[NeYf.PV
9^ceC=MEeJ9#3Sb&]\8NC@5:[fF-SOI.Cb((M(\DT_O@CJda(ff8.8<JZ3>YcG#=
V9<UUOR7[.He=P5]<,RY@<^)2GBYf^P]I7N2LZ;WbXMdECIYT;RNW4OXd/e8J_@T
dXKPUP=X]eeDIQ<.KLGA;R][TM?B^T_)b\N(@X2\[WMK[ebF?^(G:LC,aUgeFYXO
#\]SRIH6G0^^EX#gENLG])UgeJ_S<(3PO1-J27-B#3FUS1]#c+dTcgb=;FZ0.N)b
\29dV_OJFM(Ke.Nc,b^QV3W?IS,(;Cb6?GFX5Cb?^I_DG)2PD_dMU(4A;4d,LZ2N
@JMA;HCcdE-MAFTV.D,d.2QgV)Y.Hc>+cKfWX0Dge;Y@)(I/E6-7&b=L6:PR,P,Z
-2Jf,]a-U;5P1)AdDST.c&,Qf\)&a=gcX9GbOeS3gN)F@I7bELF[W+e..T(WQ:b7
d,N:AE(AJ<-aF3B:P_^aV:(7>D?ae]GS_H2-N4-@0,Rb>8),aHX2@&X#J;_\_PD@
65/f??F.P(B\Y<;Bde?.WRB#:6P00_V]aa>W<\>J,X:WY)ZM#CYe:P#9QCRFAe@J
E2Zf-J81ZU5B+U)daNOF40)IDg.CF\9N]_?K+^<-X=LRTZ6bDL631\<76&RF.1Vg
ec.OY:1D5_cXBaTVZRA4SJGP5P\1cR>-/a3M-UA&f9_6V)6#:=Nb)Kf&BE5UQJE8
=;\T8&7JDg\E4C,@:N=Q09=HD67G\FU<GfQ:ATDMCObQ;SD+XKBO_]IA:V6HCZXI
A=g5gJ5L_RQ?cP@6f]YZ0E=X0=X6)4M^L(D_KQeX),QB_aYX^Q=[@H#\f@@O/4.E
O,e\[].<:S-ELXL>Yf<:90JH[bW+?ED;;SJ.gZKXS_P-5UJe;RV,D[f_U^8+I&V<
BTSIfF927:@LN&S_LD:.TW<c\3O#W861.].[9#84F.aOfLAY#\=7/_fC@>JN6,;W
>3?O4^E<AG:I>H:R8S2T=(-_@A>];6X[Q:3O33Z/KG0EORJKSCJ@/X39MK3[6-]+
W2Z2OXGX94c)J2GTJJbBNfR]cVNON#>BfTYTLV5>^-Ig:2FZb2Q.J.FXXAV=^bLL
FYRe[KC(;f^-(V>e.fMe39>^V<G-\U0V4A5)7D])7;VLEF7L:__VTJCP/7fO0DAf
4P3Gdf5;<Y\X.DM.=g1ca[,8P)Oa?:\-8P[f6NFSOV(:TE:6-^/_TH;(cQfS0K4C
]P\(8c:IYYWMP;0K7H:X.e>?b]dX4(_QIeXL75JC&/<^QQS8F6<9eIJ[/3WG/)TS
CB#Hg4T07f.J66@5T(cfICI7,M/-N#:6412OT,[9)/<;83?H=b;Sf0?8LP7W-G[U
-c3DF\55F_9/:=cUO&#4.\B9<@/^O2d1=E5;V&RW_6?g02N;)F4.UR+??R0aS_0;
=J()WfG7Z)#-JA#1C@]OL+-e1[IJA.?Wd_c5-XdM=g6GDgKa/dZ)ARSW\Q/A_GR.
=N]eV&R9R6eL9-?:]//QQ7,;aQZ&(#3RJMFYaWT:QNaHZ^JEBcgKLeL+\O@AGQLY
L]FTSJ^W8,8A:BV:IJ3^)K+,;d<Eb:86>dW&X?C#?Wd?Ba#+\cY2]D[M2NU9f@c8
@&);WO#1aK/bQNR+_g),QD?BS,^f:6eUP.<\)=P/(-<49>R9^/(bKCZgfBQ11#8]
bZ+Z--?EXR9YCD14H<;QB4C^(P\#K@a[_;g&GS_,ZX^[c@&9/?GB0D:&GCZTaU&Y
7N,]T/SKSR@d]:UfX8?TP>ACe+Pbe7KgCJU1Y)M:N?50(5\MYHb3,E,.8+HJY,L;
]0P6@.1X+1RV&G2U?IUg[ZRZ@8f=I[ULT97Pf;Ta?V\AQ<_NO>38AM+5e?R8Kg[0
M7@f9cFIM6]=0@2_gc1OUB1.1=6?94[a\cZV]2AZ]-<.6U1Q/UF/dT;ZUV\>.RfU
80KK9X,S=WO9;e8-^_:?f]LOKaG0F)6VN^aVW6]&=S8>/(CePcT-B9_FP#W#+<XL
<^H^4_Gdgae4\=HJ#IWG^L0eZ3MV/aI,8D-H(U.F0&XW]M:fHcL_HO;/bR7(@b-6
YT-_YW[12,8>g47QdS[&KS:P-Ig]=0GCcD+R@6[V4O<+aM+VbU9_D4P0>_4&6e2B
H0,[EHfF;ROE-RLYIaL=9@)HBd:,H8,.=,;=X++<e_1&6&TH5]8\B(Y6DJ.f^1c7
1.>>]#4ZHDVEAH2LTZ2,BG9>dWP-U20SeZ0@/)bLCQ16Q&;2D\1[+TOKU#P=XHX/
1@6)-(-YDcBIA<@fZA<,6[<gQZ9E-A&(#NS-c-FKPe90C;)e58TCY#?gg_BM[d(Z
bc.BY@P1H8?DFRSQg,)0_OZ(bSSUQGO5^79S+/#D&#-W_F=:>2#^:d434.8bPY:O
:V:<>VU@0:)ADU^=5F=KLQ[2/J>4Z]7V0(BJe0_4g71<)f:;D+E63;Q-CJU.[eQE
QC^UN[P6IOB4e2UDU.#+GC(N/O2JK?=4\1dM8?b[\.aWT(YF1)#2gC[(6/,,5#cd
ABNb+b,,#dA5B-IMe(,dgI>4\JDg+SE8;JK=AIWZLY36N^aLY<HFJ0M;00K<:a1=
;N_J8e[_Y<JE8ffZQA16QLfEF]IA>(C\MXFVPgZ?C/fH]aS<RX7.\G<IXG2/BaQ]
6THX>S7ENK)fZ=4eP]1bGee3-0-3JfNR)X5S9N0@eMK(25,]KYYM#8[]MZ)9U]-Y
P_7+JZLQ/=egWeaCX:KEBX/F>+/>&9_eCHOSa@X_cc):G.:C-D.A_-@6b-g9B:>,
#Z9GXBQ7d:X)Y]>W<,-^810?T3aZMbQ@9d5J)J8ERSC)I9+8P>92LbY?72X^fR(E
AMN)<SLX1W?0U,EV45L9N1Te6KdbE7eCag.[3YRfPRUYG,+e:3X7[(FI>PW&3dW=
f->C_OEf(47<_TH>;0,O^c,AZ+Ze0SHXGGgOSV?eK9AYd(/a@XMUU0^Z<G5gWC9[
eE>,H;1[Qa<,19C(d7eI7<3\\SY[ZVL]IPU_\:F:+U8LMNg@gB,S2BBALUa<^:>&
fPJICF7I3571ASXC-dKC#^;AZ^W.WT#G@VC+P=d.@a2)O5B_#1YSV)I6QL2EcT8_
L-V)AWPB_UCO[YXb7T2EP@6\SY?DK,S=O\Sc57G-f80Fd;37L4O.EeS[B^TIK:KE
6]HaRW.2^UTAeYQ=DL=L:96Pf;Q3LJK8ZWaeS2FVPZf^0,.ES.c:(L[-4#/Z4_a.
F:T\/MRJW@GC/H:K.>&d<PaPY+>FL_]gK6?9=,:[GQ<E1;^d,BJ^R+Q(7D\8NF9S
6VRbeB]9geF5P3b5=H]/J4UDBVL\IH98Z5J(LA,eZJ5\2I[?eHBJe4/BRU5[_RM;
A<DgO;S;g+\AH3g8b?.+[9HPE.Y/<EU4cTZBNZRS3-&CYS&5(,[Fa]9C0d>8b,ee
]T90#0_^^L98ff/2-//?[:8U+CRSP@W;4B1:M^FOfeTRN>8+QRe#FY6<d=N2O1MQ
S)T3YE7Fd@QR[;#XBXT(=]HgREK;(Rd)M(d?&g5O=JS^-CW0/4X?-L]L(ee&fKDX
N(XYMX;VO;&D(X&22RIT=/;6:@1CODb277S3TV,(8G-3=bQggWS,PGP=<9.0\0U=
2d[(GUKZ,bSCd)Pd_98US4VJ8W)?@M?RPF/]aeDgF_K,W3LPCY,b5HUcM0M,-66@
@EN4b5,K+/Tba(2CLF2C8E+-H;?2,--[VUg4R@^GM7:95M9B[&:bRRaf?YN[:g(N
1^JU)a[F?Za0,E=b4D(E^L7.1O[Y_fODA6Pa<^[JKJMc=e+Z4;4G@K-O<VdD+Xg^
^<P/=bfV+CVMX(VJ9IZ[N4(67AX4K.WPM\VZ-gX([]1TbcRS;a4.5]7AK^J^cN5?
VEDca736agWZ)\:](3\6Md6bdKJ58=G+;VCJJfW]U[+_9LN2>^/9FA-OQW<FQQaT
[U3bY8B^[N:P+12f+NMJ2]NQ;K/^YAT3K+V=<f@9WU0@T6X-D]19O7GP?QOYNT-?
gEd>6>P;)H/+B95;?^>T[f,-Z>@=\8CL=19]H)a@&?<BN?P?gRXUWbIBJgIa1d4S
C_3;cEODT.6J]^=]E<Q6UWS75dZIO>1F>X.Q\#0I:.B8R0B>\,fYO,(Yd8S1)fZU
-a+d4>QF=CC8-=8#=DYOO.DC20eS.,K]#ANDbKc1.JbM;9U5#JGXEUKFZ0B@CG&I
(FA9g@3.X+[?YPR\(&-cAPSO.E9HdDW[@K_H3F&<.>HT@efWH)SP+2_2ZN[ceHIg
L0]91FV\08N\,JSY)<LaND\g0_[-?)A#1&gd7>/CZCfQY57a0fMH8:CW(T04&(@A
fHGY2_K9D;]#ORX0X4JT^Y++@7AaO)&bH9@&7-J^/U=MS&B@OM?><?-7.d]AGZP6
R/Q0HU5bF,O)P)(+XL-O=UW++Sg7NVEfT_<(1WaU[\77<)9+,@SC:2[3,E#(D>N5
4F_OPNCc54:;D^>?7^FZ))[FK):UMJ4B1Z6KO.(]PW@S(^&BNb5:\HMD/d6<_QE;
,NQ&(RU/4#fQ/M)\ZC^^7@3+aK\P_I>cF70(9&(PK2^1E:9B9gG-WM9EN0<7@]PD
C^4b3TA8E;5[;_cL]90;,LGWaSA?4.MEg=7T7UDN>.Q23GH(6gb6N?<-f4fb8M2b
;Q=a#/6H\,J,Z3=->da,BR&=+.0SL<Mb=Hfa,W=>)_&dC&+3:]ZJPTY>I&+A:eSc
,FEQ2fNaF+8,2HC^bcN5P_#YG#_^FI#=ScDKbU(YQ7PW&V++=JY86]0X#RQVU<8/
ce2De4L&:b^fDS6CgHH-WeRG8^]9[5:SSB#B,Y>@e1&PV;d+0Ac3T(LDbEC_R<W^
C+#Q#0GGDM?<#HKRI87IfQO+S8K\<\1YR>U\8:R\bJ0]686)7+g#F1?,(I./ZD-C
OK5Z1T0c[92Dd?=722C2VWQXRZg?)(F1e]KcM).+GI^DM_[1132c;??-+2C=JX&O
abN(P_.;>-)6A3;_:,<KI))a9c4_&YbcB:M,Ha/^f?[PLbO4;X2V/afFYO^-G+AA
-P>0/;ZW^aILL8L0FOaZ#WL1/.-33U0(a)5+YAH>G^O/NG3/(]Z7>RQca]>YRM5Z
.?B#LE0FKP4L\ODO2fI_NAb(=EG/)Y=[V=1A:5fJag^T.LAA5DFHFLK25G7BJ?>L
@U35QL3W?,D49eA)+N_gN#8^#dC(NdTD_OIA(Q:+>f/+1@B21-RK9WH8IQg?<b5V
?_,H2\PQ>/(H[G3eO(TQ1;,F(A<R]KdNOB?d0EZ9ZQ.;>4GS&S2f.N)7J#[&Ncg0
W=IYe[ZN;W1Dd/((K<]S+Vg2^_;e\W4>VDg>dMU^7Rd0REQ:=Q\?&#/[aWWbR0Kf
11\+.N39eG<D4N2ZfgER6YScWE2#gY6QN9/I.YSO]BE;N4aO^NRE41&?c5e@L/TD
[:A((a+<LX/BPK,QSIOHR+E,]>bVHg)S/OB@2/TNPX4P_JA</MH?3F1)W5D8B+^)
Z;>TP&1R\W^U4&2g6D^0DXS19-E]\WGK\DCT4XdED5YQWaNc1dC.C[5\Gc-S8_7N
W43K;\>;A2D][\>05D^b[#9>dc>,5V[^TYI(V>Q3,UNgI0880,TLE#[ZVPa>;A::
-]XYG<9K:1]ZB:M[\I:^[fIS)g+4&3F;fX4M2FdEC[Ze+6>-41[?d-<.+F,YQ#eQ
/@--g7f102\+0)LDUbRM_@@^_^,00fP59,Zg\3N-b36VF7[e+0&eJX4?fHZ?88=9
;[bB3,W?(J#SYVOaES(c7+dE=A0PeDbd\P87N4S(e[Z+KgG&AEGCRe3HK8T.gB:A
/^<+##((/\M2PW?495069R(dYTP^c90=QW2Z8):e1Z0/V/EFA.\_bfRNFaf4/eSB
dWH#01A);9.1O^O^)K70cT[5E#9Fg,IQ8(5)=/.OR.C3(:<>\_JA#<2A-DA0U?&>
DWR@U11E]\YN5KWe2___RR\8GKJ3PR@<,&&MU0EYYbFUCP&[C<2.)&PI[?96fW(5
PcAGVdVg1)b)QI37f@KI^EF,9H;Y-56B6BV;5\E>2d[F=bZbZ8K/FV6BeB?KFS@P
BeZ+OCR3E^X^F\WNgWVI)fAO\1KX/#MPJWHa+e#7C83:gRfPNE]M@@CSR7#]D:dP
C:QZdbE^O:[=<X,=>@1cUeS),WY<B.:.L\^aa+2WI\b+J\27;.=2G3UPI#]Q=M1c
,dEOTcWXS&\\JCQ:5)]-_Af69Q-&)+BK\F&fH0+48f;gJQd86,KBT[BJ;+VFGZ/V
PI&TE/9?NT4CPDR&D/[4.:.57aAN7#fTR>3-E4Qde?<>aC6GeG41:V]d@c-_-^.R
U0GZ6EYF=]Q/Qa5eHf8+X8^6@cg;G>C.C5QK)(J051R?Q,_PBcL?c-WCD#/YL-[d
4R[6]U0VAR:9NQ;?#_QS.2,H\6ZN,./>_A6VU5J;8LTb0;^d@V;.C)FPLG#)8YMS
SXccPO22e_HBggOYT72E&?S[U.65\<D2[bG?Wa>@D.+Y&7Yb#9T2T([95C#A7(_F
_:#9.9dJBb8;.cCg1,M.3T+G9,DRA,]?>=IY#5U8<C+9:-V\..H1V=_Q<:IgON^N
Vbg[e(+[8_QWfJIQP]HDC;fHZ\UfWF=2GK:eS^I0.)UaQ]+<:<M;c1IHcIM3#ZW2
1J7.<a]0ZcBf/4b?7U+S(J,Y-f+g:_b4FG4-GTKF\=>;:C6PI#:QA4O3QS#gJ/^/
g/2g(=04=;&HJcb1W4f0cN&?NLC@.24K2ZddL]LSaH.^^a?Z>0T7O:9_5=??Qa;3
BY77DCEaK#^X6e#;&1KD,N9L\-F56L6[ZWbR/cV,?=3(2?4Q^4JA,fS+^O?MVcI2
A:/a[6CT_+OD4R88T\X5c31e(+MRMA--I@3ZX1.DReZ.W(ZTHV2-V=@^;d6cZf4J
@6A\O;1L&8YY/S:@#[MV#XHDSa:dd2b(XJU4]Wd^T&Td(OK[@AHb2T9@KcA)-ILY
38PeW?C]P?MHSKBC8&(8)a5.H.HgQS1L/NPeg]NcVE0Z565a9OF:9a3=@RAO:fS4
PBE(Za)N#dMg7+D4NedA],gV#Z>:A)E5H4O11P9#,?[&cL=B(XJ)a;XN1=XK3#>6
GI>IC;1gR>c-?YWb;Gd;g@NOAM2[;Y:U9[+RXS9\_2)acNP_d?^=>-M/YD];=R<1
W-,.U/N,g._FdCUa,OW(1,0><>[700U6X>\>_@MO;<-&77?J-,(+QXZVCIC]#UTX
71QY<KE8<KD<LOg/+95R-)S#HUP4a+B5LBTK\N>0+?V2QWCc^#VORY#12\Q3E11[
Q#SZ]>MPgWdNOAf6d]_/\8[1/LeYE)Y5Tg&AD5W)M,c9cAg7bc;^DLc#4OUT^+1M
fI0.gIgdB,6FZMbTZ/cU9G0J<9a-&=#T[BB,=O<LZGcF1.__a<XHMfe?=SH8eGG&
\8-FUSKU9?J0EYNc8.^D2@)O:E]OaW9e;EE2UVB0V#.:5fQ2(W#[2Mf0#Ba5aBHX
23XF7b@Z2X7V6\f[<^WJ_[_H8OL_L[CSRD>1STH]T.35ES_#</QAMNdId352YegK
c((\0A(g62JH[e(Ug&EA:KSf[B&(cBD-aW:?g?_XPG=@+Tf\+L?V#Tc\SHeAeIXE
^)YD>;@ag:>A+D35>f/T_3:\&dK)OIL[5Kb7E12\=4FS<KEcRI8LI@RWHN3gVE]6
R@:7S85Hc)9dG(W7+PE]:]JONLLL0Q-Z61g2;8&6:HR::XW3R<>/7Z.EP1\Z,2(G
f(fdSD809-Td[1T3ecE[5.Vb[Ub/ZaXC8,A,1A^Z1F?=EJD<gbKdW5^bK)O@C,_F
cZL=b/7NP&)??f@M)Sa;IXO])H6E&X74e7U8B3-9,GH)g2D+R=HZ1bSJ/EI+,/fJ
,K?B^]W9NHU8Ec/Hf.[(a^>_eC(4Xe0YH4WUg3S[1P=c:O[9FUG39QL(&)0O+aJb
Vb+OV[#Af.V.&1B,-CDB<HTRV92/.WB:OfIAZG@O2fQ<<28[Sd;^#-OBA[_M&AU:
PIfE&]CBMUbDHZ^db?5X:f.Va/7\U._TG=[27OLJ0WgSR+OW>GZW(S3e&Vbd1<G4
W>@CF>HIfXP)?Lg4PO#+Rc3-@[BH,=^-/D5-EQ(Cf>W&1<BdI=DZD[=TA(@;?]c7
@95Y.I27[+F;H\XQQbef7(aS#C9C3We3>P>dNOdF==NVZg0;d3N2cEK\9T@M/A(A
1_)9:HUC2P_R4Y]VLf5eg&(bPFHPK;C#K&^AV[&\PO>@+g/TQBQKDbffIebNMWQV
3,?HOB0P2((G)V[TO/==g67]8<[/./_DM-@RIYE2B@IIIJQ_e4(e;JQC/GD/HAPc
Z1F+1,_FWcM^I/T(Y\:R/]Z;.=)>TUNHYgZcP&1H@UK^3/JFG(_^Ua4X<([4\-+T
d]1S?:8LdNA9\M:X:AKAD(BY47ARZG;6U>[:<b]e+VW,^g/5,AT0D]V[JVcW1Uae
(N1X#<+g(4:J]FD58a&.EM.E0OVDH3^@bKf/V3@EVc7I8WO&G_7;A[3F4gfe4[BV
\33Xf8V;LIdFe8EHb1^;F(K@F2[6Q0_#3YOg+aT->DeD:e\6P=X,G9]R)\2OX[8[
@KL40/@BFNO_:U2#@[94[C.(>gBaf0\N[&K7_QORM-+)_R]<78W<0O1E+Wg^(XJO
gDO7NSCf)&[;Xd;T-1E8PC)XKIAKI,SI6^QD2JV@HGG4:M?@2C\DB().ZSg,TaJ_
;((IZ&VS+9PRIZI-Db3^YZZ0PHFagZRM])\7V<KD0:P>,VE,E\W,\efYbJJ9NBS4
PTVL?gTW.9N79UL:f#V<=ag.7GfXRL9]15Q=)LM#>-06GL4,^MbDY+.UQG/MV8S<
IcIBM_5X+R-I2f6]WG<L1_-Ke4.+6V.MJ+F8S9_5B8M(L?0KNQ<g1ZS7<TeEef]M
@MFU:fBQ?^7^EF,ZUY7d\?M+I1H+>gUa_.NKPS=^MCWA))R]^]-Qc@[S9C2b1?>N
:2.R0ca6+?,1WF^>dTd5YeB)f[Na\2E[O^X:@_^A.MgV0Q/OR=.>[:UGWPdBW&#4
]9+VC;HD4B1G]/@]2I;46fD^I7H7BNGS:ZS1_#?5P@OS1]Rg-:7C:>R0e@DSZ+IG
H,P)?:SFO46JRWT7P?6CXF\7TgE3HN78YM1=6GgbSgVMbG5\@]UeU<_-6UD?[GXN
Y)(/f:;_GYON\ca8IX\>]bAPBfZ2LMOU9Z+5^591IS##,XbUUN(EP,U.cU3bR6Pc
c/Q=UDXe4KIW^6.R?X\Z/K;aS_A@REN&g[&DC.[JT#1+IM17>b6)BN(+E2KKYP=[
aQ41)UfAT]aBY+UR2+f\(U)CZ);UAYSg45KM]S\-J#F==7\M/a-606WU\LE3Y[G/
_T/POD#H\@=84Wg^R:OHY_X/D7PQ(gY><0XH2M.W24#8X3PBTe#1Hf/C,/D;VCO2
:F7C).OfQ\\bbS=EM2@Lcf-=F=-Q4f=435XD_J)F_Y0<_2#.&[3.20cVHQfIa2Z]
;^7VbU?-MS[]F+<BQg#=B9Kd0R__0d,@Nb._#B?=>/>YNS/b[\;1^g)cT_VZ-2+0
_-XK-=3PGM)+P/E2J6Y\3]AV4N=7H?_g/f9b2(89Bg[#WXa1AE84FD+R[S@>+#DH
-=G(WOO??#1,C-A[?(=9[?X>F5A]HZ.68AO7gJ_R+_/2LBM5<&;W5K,O-Z)V98GS
Ib)],^AR,Y[36ac6Q:D@,WU+26VEO#JFG[,O6V([U1Pf[)0GZFKae7U#40]8MS==
5_^A@QAT,WH\L.C>,eb0>R8c(LCFAY40)+fVP:,HJ;eaRI,.T?<F#1#B[@gf0:]A
P1N;ZL>[,IEa2/X5_EHdW2^dFZCF3dMD-,E&I,CN./JC&UQ2YDS+Edg9US9CfBZ)
bYca[5;gK)B][7+3<G;WEYe?I5#f,V.WQbOP#JA=A]0<;L#e;WT<Nf<fBK^bI+GM
+e12&-T3d]]4ZQ=&0U,59UJSP@DAdUgEeJTbL/]MH>eS(:.HUX@eeV)bg2/@e_b2
\8I+,D7,23Q@9dG&((MYIND[fdAb9>.=F&A=-R-B^P=PD2-bdP28T4Y3TS]^+SF]
O)f(@^L2BV&]R#YK#1Z&&4f(;J:4cW0S#aWX?]J5WG.A9aLF(?E3/-,9Q#U\d0,a
M+Ygb/=F=&7X\NcPJ?R\DB0[T-dP\>Uf)OI6;B?4F0AM.[VYKLU.;K[U^JHKc]C2
/&1G]fH5D4-=L>=cJAO?RcE4]<Z+H12?4gA]]BQ\558>;We.4d;V.33g72IH1J[=
B@PcO>^72f)RSUE;8W@^b+Wb\)3c.cPY3-O\db#:9)R(bLOZ3W+8^WK2Q+0KV-+_
>8_[..[][W-_[P8#Q[DKb\fY/DS=XNfL034/OY^HWVc2DQ/WM\1Dff##g-AZ2)e[
4HQSGa<,#,8WIB)4QXE0NL=LF&9J4A+<B_52;<O6@WGZ++^L(5NPG,(2JIBgf-P5
Ib;G2(A/(Z,G/W/)LFe9&6V[-UTJSNTedH-H,V_;8_)e;A1V<\[ZQT;BH(+5\SJ3
X<&-^V]6-3C[2B82&LDBdc4XT9&M/2:C>P+^OR(-G4<C4-M34(^YK24,5e)cA1?K
PESNKTK\D4g8@eegW)=b)N5VL/#N@^+b/6.LT,]A/ObGSA=T.DI-Y7721BQR;;B,
T2Gf?gM@<N(fID2)_B2MI(/D]]0f&:C#a8_3^0A5(a4([GW.f/<)GdbQA-.]XcZW
&5a#AZ,[eAIca+4P<baLX:]ARf2GYCU#BN2,72,LOG_=JM&<B9E;KH;C;PUHTW+K
89)Q))JF+O(G7JF=D=cWb?GdAb)JdIB.XUQ_8dI0L#Qa<207;33^ZU3E1]0:2D1C
EZFK.d-\0OLW^8,+8YU>8Q5BCN&WDSQG,2>3=VMEJ#0OZbKdWScHJ7AM\:(R:2Da
_bgW9#=:39#\b^)<#LP,R8@.B0?>K@4YDf#.eZL7BQI_C]4UVMK3gR?F<=82^Cd2
T\964..66;O-CHVHO8E28ITQF1\<J]J-R;+?X^AU70H)cQ&O/A#Med]_cZHC7QW-
:X8FWPKB65PgH^LKA[eZ;^:MSLH#/BP<0GUddO;dV+H#,b+FM]=)WFaI-g6a@_LW
?dZ^)8<3]L9.]F7D[MM)DFdUJcZ^F6f1&4OM@cM0<8.CW^K>Ta]2I1+WI4F?PZ?R
>IGg=8DUZRT],P+K5OC]TEFg8DJ@;BRcKD?d5L0RKgL8=U9J0/McbMeNO.-3^AXK
NQg\]/GgW+9&Kb(D.UIUfTBR+Nae^B6QDWPVgdA#5,P=BKbJ</-N^)U\_KG6CP&3
^W0H.5Hbgd8(4:fD5YE4eg(?D.4ae0A>F)aWSP=A4UJI@@47T01[^H#KY8>]-@;0
Q9_0TF+8/\ZKSG?)CD2.^(];HCda_@Sa^fGM4Ac#.g=W@;DL8M=KffSf3<>Dc>OJ
>>(8L?bHU,9584[(11<]J]T\-c&1F0HU9?0,bG<A_0TPT>FQ:FI^7[(7DLJ[D47/
C-TKYD;MT5:B](V9F=^FK9TL>O1(/QC+]ICQP4-07:P?Ub@>K[:2]f0J6F)9@^bZ
@#,)\AX&^WC(6H9Mc[9=J:86MCB<2gW5OUTGWW9+ER@)gZPG7d1LbUcX&Z6f[<7G
?6#5[Qc2_AF>.I+8@ZN;N4FH0V\TQ48LLG^K:4Qec@eHB<b/6U5[;<&bJKdGf\XO
2W0dC:U(f&@NO#&_788>,EDbK700XAXI?/NA.TSV]L#W(8[.MMSFIX+gIOH:+8U=
f)XJ&7+>+@&=@Xg\dXWI\1GRJaVg<)/=<PF4MB>>H:^93B>/+OY[IL@\G,QN5YbP
cC_\]CYY4I<)5V4PL+cS>LT_R]<_I(N_&Bf/L[UG<4U6>1L7G?<^bZ9;._:d1WcN
(PHS9^f+&/JV-]),A[g5e_Dgf;I,g7g-BBBXfeMJMWR@5)V.Z3)7+^1gcfF<fF,8
dOb)>/7&MAEI\<_37@.X:[[OAAZDHJ)&?>R1S08=R6C-6J]F3[L:)F=aWIV+HELU
0K,[+=:WZ(#2/SWWZL1R3(.e,ce>^(S)2U(VU0cdR312/c8EGV5KZMg0O8EV+a0-
3H76FI)>]NUSa+PMRL),[LMX?2.LA6GgO^]b&310Oe@J(eQc>-6&G:+d.(b(ASOU
ON6?QaCd:e_>L>BB4R45ZNE+df\&\XCF<12BMH.+Y[^R/S)ZbZ/EMEU;[.G_]S6P
OV@-NP^;8bMf:\JQ+?[I1b[c,10)OI:S1^+gV\aV8R5DHA[2M<6-),MGJNGDf42B
Na;W1Xb0=S1W9UbY>=PZ^<^WIQV\W=P6MK6P80EbPdfS<:gE40\#C-^SJZP;<]]B
gbQFdX&;#OT+g+QNVWFfS?/89W,]3O-XC5YO)Z.LH4W9=4Ab&KegE,=2<RJ]ObX<
-ZK<GT=T8>W=;&>.UN-_EYc(FMCOa:HIf8AfKVW82(c;6+IM,F\NP[_Sgc&\7+e#
T+6S.(QXP^cH]<1g]+Qa)A^[APNT6(Q=>PZR5&27KRB:2-ZL[CVKgS<PU4;2)-2C
:dN@b8]&)?E-5DHfQG0FF.+.?bX(JAS1B1dDR\gYUA332=/_#M0(Rc((&J-:47fO
K5=U)e\ZcfT@O?<EQUTS,e412d&I:G>AgfYUf4FO.NAI5##GA4M/^a.7C=M?d,cU
EAX55QACXfL)EXYZD+U@L7[O.>g7LYI4UH,(Q^842CcIOGP,VRc7N0W+75)4Pa_\
06:\<0-S[6fc[IQPE2A4ccX=4@34WFfH\P@)b1WJW3CJ3L=^#E\bYYS5.?KNBEB#
Se5cSA+B?5cK:[I^YRNNV,WKM(,\KXRfU(@7ZJ3@-/A-[dL]RNYOHNV1d&+dLEZ,
3(HF1]JAa:c<3T;BP>eRg(Y:?IggeeXQE9@D10\O0;F.IZR1#K9^cTW+^K[_bLFX
>(914V&WZW#gde#K.6MeFYLB7efcFI4U:B9-(aRKG:\N-b[)[f9g\fg)NQ?5Xc[6
U?e)T6KGaD3,?XHTG:gQ>C@.gA477SQf)_5Mecf#AdVfd2e#)86:5#:YM(48O<<U
bX>e<Zc6A\45R4P<a_SfN<N,Z2/9^HC-@a)b3;G)(ZfHLB52DD>3ZEW7bTB9Z;<d
PY9(C[])P+VQ2BZ<L>B7;L9AA4/P]0OQg8eWX+&c?0c-LWG/U96-K_Z&eB\L-X;S
1D-8_#T=LXgAGBSQE8I-fBY9:UAaYdA_]0R.DJF_R;;dE33ERdR1d]0/@/V^GIBU
\g^GJA&[=:,UPHdEcO:#G8E(G1beadM@dUC8X/4GIOf](N.>Z8D@/JFY<Lb,^(C@
cXH@D4?PT1&(WX=&FaeV04V\J?Tc)8HaFSK^Y4AD_:<8;R0\C&EWe2cZ-f(?[dM_
Z]<@F8^Y#S=^1X:OOdET+gFQ.1WDNNZCO]<3MS0+]X@.)CZ.JR4PZR8>KE)#4e)A
:AZJ2Af:<a\0>([[,G3W4P^MGM5Z3=Ua/aH(d+6SPVa]SUT=;KQY\0bN/7WN;K/1
S9FdPDA_U939A#^[#\/CI+H&@Fb?9=S8X_?XM:>58M8W@W>K60+^A3SK=LM)7J+L
fLR60[;5.\H7_VQX32Z+:?^<5Q+]CeSG<7fTGXORH##W+&IXOcY\Xg;@b84>3=:C
GL-e\[5<N3/0;DPY=QIdYN87X#Yf<(^URF/#]?cLLJ3?A&9]4]Z5^EP/dYE@I=Gb
\cTe4TW,5HcKCNQbX6T28>B\GM>]<^2.)&0X(d6R^#F3/&]Sb1D-ISD/YX[X,-FU
6SV>:X42^2+aeELG[#IW[JE7B8,C_,-VAR:K=ZD0HKOJaS6AdcFAG8b&(,32W0P5
CUYaMC/@;@_B_[L<He4N[GG[QQ9?Q4A[;N&g6;L?=4IdK890)TJ15I4^=_7W[N?;
/)d@R]EY<(U^+cXU6/U<d.C&PIDd)NY<+Dc83A7P&bHB\1eb9H8YSg:TM].@KY.&
g8a6#Tg0eCWcO]/ZB]+Ud:TVK&X:=SgGSSXdIP24R8\0KH9<KIQcRLa82HSPIV8V
=)4L#SAe&0;U+>d/Pe-7/UWOe\<4/PVLTOb;_0)VA\^N;;RFPBPIDVWI;b@/KCXc
T/0WJ:+P;^JI0CTU,>G#\?M.X@E2e:4Xe>f:Nc:>@(252+[b6gLRB_</5bX1YXME
O\\>LWc]>/PDB9@8D.)52Pa7[_B5@)?5QI9.@&&M@32?8A.@f)?#T2YUDR?b8N4,
Wb=(6E&^f(:(0.;M[5GQg&HbZNHAF&RBP-9]8D@I7[DDQN=;L7/^[]L_Uc7#CL+/
]]]:27\,NQDXW<aU=f=3AU7;a:-F_M5,AM[N@/Ae1LPO[XgM#+93bH(AWJ-QDTS>
VG_NG2S(Ug=J^\TRV9gSg^X<=S(6Y:Q,8[&X84>V[aWQeFX0PC)7O1(#\OgS\PX#
1H0-.;#.<;&)1:M@;,A226=,1eg&)(+88c-;_Pa,?c[3ZU9eC1=A[+SB:+==8OEU
;8:S3SC0gL&R1L))#[RUI#;f6\G_JQ(YHP.>b1<FQc-\[?CFg.JFbcP8Ma&H&^fE
&V4+&UYXH<__,82e[SP6C.?&c]IOJ:.\0A(7>XA]Ygg+>6::752]S>BNR20a@24J
g,<MT.(-)EAB^6@OKBf-#>=,I?@6/2.3KfcNZR0[Og<TG)O.X&BR[2\(V6LPEWc=
X7)U.Z)==aNAP7SG:?2W[a\K(+a@W/2X2-Ya^e8/7C&GE]=0[^5Z^bT@-0GZ+NU@
KP;75\U)=(;0E1+>WS_VIg=-+4F@c+>B(HE8V.QF+7J]M0FgQ_/;UX.\9aALU\AF
GaS1C;OUH:\2).MCWB@E<]bN+-c0Ne;#,VK,<P^G]-Da_H9#BN7I2U+d-.bONT?U
YSaV:V47I5FV_b#TPTQ]d?(Bg8.T0,P2_\2N;:/IAE)#c1FeLYeS[23P^65c1;TO
ZPbR)0.b&Qa647YY:12a86=2==VW=Yg2^T;^Z_SM9MRI4GLA(6d2gLX=A5ANWd(7
NIX7@GBU7EN[6/U<9^CVG8I39CJ:DD]QDU\/]NQW)J8fcA&b)/-X_[=1+9.4]/[#
-&?=PK/1fR-=^BR#/V0XRD,S,d1QcX&gXgTNa0gY@XJ(#fK/_9f[#>C7G2(+Ng/E
Pd-c)_S\N0LF3/YJNDQ;GG_&^Q>V6@eeJg5&Wf=I6b)1<YRU.R4b2>bN@/V])9cF
0^D/-(,fQ2:][HXP2:b.(>X4b9f]+Q(OJL5WRDd:,gR.#1&T8:,[^0+<U52FWTBa
e^NOYURGA9OBV@1LKHCJ-\fC=(4(,IUEPWAT6HE1H;E+_YJMS8S/.<HIQ.:Rb5OI
T]/_[g4?&\1=2QI9U:(-6M12=.@cK2eZH\3VS^BYDV5P6Xc/&U.gGC/K,Q63L9Zc
ba9G_J3#Z[fc8<86CROS<?V7YDYaY5;B?VP)G7#<HRQJB(Bd056NeIPB3?HgMJQI
;^aaJ9C+[:=<aO\\#-TYTD)0&G\a@6?D-[&1?N7EEb1MJJJ-E6IHB/4Jda\1,eH3
^8_OQ=C>d3,Ke](g[#>f@g(QMQA/-Jf4VL_)DO+fdNbQS8RC-RV2MJYD-=N(O8M]
KU+YIQKdN6ZEKZ;S^J</Td-GO4X#\:V13<;eJc_gP8Q(D#E=2DcJ;Z4>?CBI93D[
-N[f8DcO=S6FQ^G(Y]VU<+B_@34]/6#FU?ca^(FJ0,#LONVT@1BXXV29S59Y9b9&
@f^28.dDBAa9#eTA>Meg^8&.VNPH^c:YI>I6GfG,RJFL]5M;URPbaJL4S2H=2:IV
4H-H.@4U\(WX41/]N[.4N#^Y.\<P:[DUcE&6DEE5K=6e@AR5a-.?C^Oc+XL2,?)O
FGI-)T5+T:d(=923J/+9170U?-0#8Ua-C<ZA1e.>ZVa[R+9bfNbKBN>dA<:._[bT
T_SE]eP@G^DDQCE,HE?VgV3+M&NGEUAF#E\]&(^2B_>/B)<cfAS,Fc>T_N9=&F3K
@PC/We[<-P_JY?EN8JbVgL5f<<bRCR@J\6gPad-N8O_(1_VfV9S&Kd+RIgR2S0L8
8_]LgD0+def9bW_HK4,;R_,29[d4+[c8]]42a&O9;BZV4R-dCgG2O9S9,]Ze7PO@
#_&._34b\[-=-e&.e[[cI3dd;V56<0=Zb9WBE.01#QU>d3d&@-cZ;^g/CN^LEI8I
9cW9+<2Ic.aR/3eK.&J@3:O\E-T6(#?S7a,2DW6T5<d8gd;d,g_2^&R>R)=cTFX9
P8+U2#7B>RdLb/<bb8PAfLgS?FcJ3;&;W>OIMJ2Ka#7/HB1EZ3FP&VU-YFVV>cbI
f9d(6YBD-J]:CPWQO>COQ,H1YBU>GNXcFRJ3S;@]V3=Q;JV_A0Y>)B9aKJ29]]=/
3[NHQBXL)7]B;HM??7]AM<&&)F<QK=C&R@JV(MWQX#SPTbQI411#)YedF-cD^&I+
J0cg;X#ScO1Le;+<Vf.?^?DG#b-;5A+M&aGW_8<J8V>G[HZU25[#TcN,][&e>&J?
N_PbaW[RHLUQJ)d?Ud).76)Q4(BZS0:=TV7&7#_UA8DC+XAaGE)\9aWWZ<;936@R
UL/YX0Z+?=IA9J3)83HQ=7FI;0WFSfaL\Ed?>G:2;Jd4[Iba<YLP93#AV>ZY+]ZZ
HfARe2B_=FWJ<(d#:7f/CTSB?Y#XL\D[;P?1_+T;B=L@X+^\8ddZYWe#E=Y-CSV4
8C<T?BX6D0IRQJ-TG<eMD0YGT0M7Z0+-6/fYNV-5.#CWSS(_6Z:G(VA,QG:L,Pa<
/TI2b95M#T,ccB9&b+]6<U9f+Ae9#+a>5&77HW@;>b]U=N]96d^DPL5]K>,eT;K=
(8K&<I)1L=&eG1,1=<JS,+(e:>8:dAP=2IgWSIaSMG<99X1#D?e:4Rf0Q9BAMU^<
69,>:MY9X5AQZ_?RBA+/eX+cVUXAf,9T_F=#O&NJ@a-3<CP)E;Z@06b]+3MY<W@G
Y^+df?882,T^^;24C7+O4CB@_[A[?NU<4d.>RNDU#cAdbZ[W?XL#c0Q;_);>O-/U
G5gB_D[f,/W>[[-J[IM?IbR#\DKO1g7747J-(]#S,Z>21BBO;PC&@Q[Od3@,8)aM
8KC/Vb9@QO:YeQQE?LS/V^b+fe14L+2SW;^8VO+EA0+0OZYKX9+/Y8fN3&e^9D83
_)6,CXeWP).5Ad1HHH5/-cAfN.I4JBX/+5&>bPHM[S,6N7BDA1\OM0[4;\g=ge)K
;NTSOOFC3.#5)7=/L,E[N[59(L84)((MPLELQB>0:Z;1)ade.M+9&NW>#.DBBccT
fGH]gg7:GL2;YOP6^06;7T.ELC=/Uc0\B9MQ/@C2M=b0B0Y)IM7Ie&2BM8:8W<H@
RWV(90AS8+;EFeRL-U=?1)=,J>4#V]JCBH;NLDKgJ\[GDe@2:->6G4_8Y&]>LG=Q
D8[FA=_T20+IT;EfJ8+=K(_f6H\MbbH[46]QB;[8c=H:-6TV)IY_I.NSK<L<524X
a1d@0=)8PI>S.MA<3=<&&B-8VWL\/J@;>+W#LIF5BBXaU2(UT,X^+C=#DT@R^JD.
?H-bf-85_g/P(9eg3_5C]bR4:?3MZ4C6N<Cf?7\9,&.L/ZV6OTQL<1?=QT]]gK8W
dO53-6(Z;-b&D@8[H(/SNDfWef,\NY<]/S,B@+WBV[^D<[PWaQ6Qa)B@[5fT-RM3
8H80KOc0UZZ<,a/B3[30G./X+b#,1aNFW)DRM7J6e,bbAA9XQD^BL44JO9=fI#H&
0@LVZ+B[_)]U#W<(Og\HB2=WRMLTZ+H<f5Bf9?8_A)0eePM+>cKKB.L>;-44CCgH
b7e:#I53IJG#HN;(<2-R#IK^O;OTaS)K9Z\_#OILNKEC2=>?QBO,Sc<-:Z#OIO93
1A;UaZVZ+6TC]CVRI2?S5dXcaN,8KY]AaG6O5a:#REFCKSHVQdE8KD?.<BK2[T(6
ZK;Be,ACBFgb;W#4VS\cc_MVd#TQ?U,]ZX,(D95Y8cP>5&U<Cc@c4X1V385XV_^/
40RfG4HU-B5Y>WXU-H[R-WN/)E#&^>.@bL&R,SMO2X,KZ4[35DZgF;e(eUK55XWb
8ePPCfX2BbJbfK@@99S7,X&,e?=:V@HEF)Ra7SOFc8A@EWIBV]TA5^32X=dSg-)e
@U8.X4:=-L/##_+WDZRHPS7NPc_+P;f^Y+]0V7-&[H@aW3XDTW#)egB.31-GW2)d
0/)0I@<_=VZ,=?.FURM\KKF_;6JU#9+6R45.M,T9AP3&OfW]HO+48CB_C/MGX^8>
&[.1TP\;]B0LG9HZcQ<HXDGM-V^,1<.9cA#/d,f,8CJ[Ze0<cSdM:,=K-/5)1e(P
b@0G8P.]1ZD#0f9Nf54Lc[72F[_d<Q5IB]9T.=Jc>7<C127)Y6ca&F3D1U//Pe6^
XR:\O/c;[c[AH]K@:>3\B4-H:1(3#9cBcfM1fLXL,5E-R&-#OD,3)8R=,W7/bea.
SHFaE7GeJE?NdRLIa,QKV?Qc@.[SEfED1&[=L50>Pb8L0Z]e9\=WPRPC/d1++,NJ
+e3&a5,9e2:48A,#;PSNE:7Hf6.Ug9dWAe+:0b+aH-g]95,6.J\TT](_F]G4cPHb
K(BT4.U+5eR?C,<:L:cCYIW^PC[T#Q?+(@;Z)J]63\I7fRY]-&<>TG6G.XLD@[HM
gQ6,Bb[:Z8ZS/;+JBL])T>&McS9[P,XXV8>W32PQ_OUC<W6/-L?6+6g4SdS;5^NJ
#Z]EA:E\&A,E_L<bf7&\\/NO#:.4.^?NF>1=UZ=T5-c];NFM(<3d;eSa8=>c5:#9
a#KOgC5:8-GARZ]?QDO5Q02b&QBgEMI+QcY/(Oa#KP>fMSa:N@D,b4KN@E2=AS^>
aP-VBSfAeUS[BYAD=YQ[8B.)ROI&:?@GDR^EdOZD6(SR=bRQTA=W,b+75FHNNE+:
I[GVfMBTUB+1IE/a=363(<B/_L?U1JO:._Fe9f1OV.?a@SGLM4Uc[VM>D7aD+9.[
41eY&I,8ZER4VY(8&S,5UIT?<U&gS1=+@NWJP.MI:aEFSXY7;0R3>a2MD,VZ.(b.
H\K#ae5e7FaF;R3K&@5aCc50)W=X[9.;ZMO;J,&8Y=fDFYSJUKHKQH);@-9XT-b/
G;1=EO;#=5eH#JSD\>6L.I>e-&W4<MfO<-.T9d1Pdb15295FAR(=ENR3DF]PBJK_
eF1-NZ?7[#XY5>96@2E)FL1UD)M5f>@)XdH&a>OFPHfF]C.-JH+bYT,733g=J;bF
_fWbdVF?PPB^NLb2J3IgeTeH-1LX4CW(768CE5;H5c;_@:GI:E#)GLZK?6E=V)_M
W^C:_]7)[PKE?=:bf(^+#YcA.V^7aFSEY4E0^2Y_aO1b.Be#?9A-N5+<fD6b76:-
@I@E.0BQU=VFO<>;cA5b9bbMX3Wa<:]gCVY\-cA0[[#<J[cUU8T12W=G<)F&PH22
<OOO0]GD;Aa]AI7[MQ#LLC7MQN8U2[CKMV0<34Me(.F?gP6J[fB=@R^+ZPWAE:8O
]4429OUP76[GX=G_@NX8E.OcGI(G^II>:A=^8IS2Y(O9:PI:Y6S,_FBX,S&<,7/E
2.:,NBfcC.f;OUCYdF&Ng5F6OU8:.BBH[KV3dR7A9D6BQB(=IAF7g2&9Dc#-[Z.S
8Lg1?PE@+)CWX2<RJ^Q,>\DUK>b.e:d\bLI25+/72]G-I?4G?\e-NZD<&DT^TY#B
>4WHCY@.NYT8]I7B,K;0G(6eX=V&GHGJ@:H41)BW]T;fT);\BYHg;e1053=ecO#V
A4N(X6bdcJ_DZbDb>1:AGWGACKMI8/FKNMVB6XEcO47>+9^CPB;D[/62/VM@^^Vg
2-GL01f)[FI+<J74=3aYe>:/WY)+QD3Z)Y1TR4XNO0SL_bac5A_QDVbPP,FG-W61
V/a_RdXK\e9VU7?;L7b@>8T)H=]/HI0NZ<\3=PIYbM2-H8X(Q2)OH_9F>3_LQ5?>
MQK=?:@?3JAJ4@:D.bW60I8HT6c,EV+R.CD_<OW;g63-DII@OTO^e6_G:USSb;+J
+Mf^,e/FVcJ\67\G\LR=@cV.+4K5L1H.B5<WNV\)L<1K1f\gd]:e,DQ<#N8LaZU5
I3X,(/[Da;B#P-BeQ(P[Tc[9RDL5?M(Z4OUbXZG7]M?&DP-H?fD[0<Z1TNVe\3e-
.C^f7W6>=?RG>4B,(5+^&\gGPMcVOI=2A--9BE7dR]VdMB+gU<:NVP\a9^].<W.b
<bUT.67[CJ7]C/I/0H-E6QNEaK[?_3J2]I(3@#_dG,bN@D>L(D?MQM@83+PO<BgH
M<0(].UeGF\YZ\6PRe]g.+J@0ac=O[FdJN3M9^7Lc#>:64KKJ>4](B6gS)V=P?D=
?14T:0B\2L_b.D&#>M88X.8CMWe+:YQ>ED<@4d<WHZBF(;3L8V&=Y&^,c3W:9,dQ
d]Z9fWb:.a?(3,^S]1Y4EbKUd&3?)d\<E=Q]-8Y6T=(3<RH4YNW>G6^,K(V<:9c1
-_&=3-]#_XN;fTA6/]_RIN7c89L04A#=0-Z,fOdHUK,TZ6#dSUcBSXE]J7VN1RAY
^2C\UUB_<H.5;e.>23P:IS4:<,@?,Ua4KNGY-2,?+\ZcS=?a27]F[Ig^154dgO^a
d<58+=;dR5fJIN#+@@X/.RQA,]GU_8^H#L\K4[8Q>eE9A6I/^AL<UEBH,e,bc2[(
_3/<d0@[>f@/)bHJ;[^:R--,9EPMI_3<).?LKK&/LRB_fR_UMf;,-[S/_ea92PA\
#H]O5,8d^/JT[/FaCb^0D+6MQJ</-LV3e=B6K_e9MLEJ;CVQ797\4[DL1\f>N9dV
9cS/JQC&DP=2ONg6,N1#FdTZX0B4_@BTX^^6,8g^dfQ^3H09UC4374YV8YS&Cb<@
4<JHACT#P76LaG.g<fR9L)Ne=Z7HMU@7RFc/V)N>cUMfdY7QRI0S).RT4WT>6.U>
?#dQKUE[)1MTLb_/bAA1R:N:^N^;LKU@9THJ^^&=X.6M7/(c57M:>,&7D>5dBf_<
d\7WR?Y,B)+TGBZ4#/Q2=dTEYGQVR,<@c?F\2:+(1aRL7TI=;>@53_,5?HE+L/OQ
;E;_\8b86]0UJ\&Q86#UON9#I\-?;4L[_[XdY=7\U]fZdEf.(;DKb/e&.e-A3K0S
]ZV=@3V3EXP5/^Z4B4c;CIfZ(6cD))CWY/0faZK,SH(XQ3aUXCQ7,+78CS6AI^_.
//0LReSd;9Vd9BP-d4B2;I@a(:CJI^L-7HFXTUQ1>1-CcIRTXP8<RA\X(NV9]J06
;@M]#Le62SS17\J4e:K6,7R,BAU,00&5<OV+4e2;^gTg7Y3^(cfL:QU4(6);/LN6
<..X;W?J=RK<^d-dbe;YLgA7YEZS0cPQ4^[&(aN8Y1/NR?JI5a[ED:E0(6]Z11NE
[?9_Xb\CV+a=>&?e]&B,S@B=8ZRD^&H-4P1MfabJ\<A#geR_^C(?Lf-6=K_4UaN)
Hd<P.U8f(:O)]f2(WfC1Pe<0?07&6VEa&64A>5PQF,NbLfM7CX8S,;&3/));V(Af
5>Z;d?J/POW^##Z482J129D@SW@C3QM3S>_Y)[:].L,Vd9Z^J^#bVL>QN\R=eQ35
CeeX.;XNJ/^QdeQC/QUS,:);)>#cM2A:L]19J21f0Z87Rd:2;gHc#6gY5fO=,Ye_
W9)U(2XIeaNSQA(fGNJI)34f?P,OJ75F[2ee6==6D9HKcX;MA85QJRQG8/@5^,>\
a+@_HEXVSP,WUbcAL3E-JF/86O1Y:Lge]F0617:?40;CD@QB/+)+U/g^Kd=;<P#g
gMH#,-44@JMJ0_eQ^5_GdCA_.G2,:2(Z.5KH0-O7fWXDST;)E(LK2KP@-,SebHUB
Edb\O:&43E_JUUC^ASb09B_&>Tg[X:7.d?+Uf:4;ZUc+MVZUL:b8H419g,3cT--:
\Me&6\^M&N,-5CE6YZDX(E<ZeS32D;>,@FFRGNK(G/6T3-=HFYJ2c7E^X<B7IVG2
FcB.P1IJHD#AM>JS60?3c,e3g^6Q53A.IN&Z\Be4(PQ(4(4A6#:.5#,#Y/).LRXW
KF3W)(5I5gK7f4SSK(HEdWc>_O=f+F.Y3N^M:,P5:S1YNT;@P?<CbP6OAZXJ->IS
Q:cL9ccG+YeG@^HTa&LP]c6a386EDKH@I_P5FKLLU8b0L_W(6>)Tf(FSKaL:=9O^
9IfMZN-5L908eDMCY]X,UBSc\[?TEMSWL_,AFS+gG0>3?7KAS3D3JgdKE>^RQWeF
?I3Q+95fMF7HGR.[LL/?H#5O4T;[bGM_ReZAVML5P?,\,TGSJYKL=XL802Z4LeX>
-3/2YVW+C<=Ue.RM:aB_U+//#XV@a^E];J)LXJG1=Y)EF;DgGbZFEU]B#<?b)HN6
Y5b?JcUe8FQ&LRbBdLL2MF(G4+.F#+;68TJYURO236QE]MRSZ&OgVgRS\(JWP_g+
7#3c8@I]MHM&9G)\?9?KA<=8c?7^_WPM5fg)LgK&[H9CfgX.<6dd^^<fXPdTdga5
OB4QNY75McF;EW\@0LcUA7_S1OI4P]+S^I/,M8/MT&)6a@Vc?,:U&e+CA@d&f7NW
>8A8S\4#NZ4LYG^ZGgKfZ@^aP2BC[VXc6OZRbN0XZDgI1X[X09,V2gXGBRcFf7G8
?9+XfSE10O8baW^/,(67SK9>GJQ_5Qg24RNN_.:[23c_)=?d:YN.SY:0B@:8U-2T
P4a;O[EQOcPBJ#QZR18D7R0ZA&NOZDedS\MS\4#2D-_DZC<QJ2;NF1\a3+G04B=X
Z[K\9@&CQN]?TQ)_Wg8OY.ZKEW<]G4dNAOY;#fZ<EgDF(@R#/@_W:OVPAH=QF#a2
=8:b(AdfP90?d(X7-ZeE2O?9bFO1?\D0d;fDBfOO(QX;]\0G6@JN@+52+d05cIC5
LeGN,?8HDW:(YHaKb5gf^Q4Pc_P?@.O=BY3e?4)E+SC\4[-SN9>VVAV0X)VT&c(:
;ZF[)31_SLQg1D:Nf&Cf8VC<_5&Q:V<(A:(W06Eg&VW+>NX,>R^<DUGEB1TUffCN
be5NQ6GV68QS>;^Q-^I\O+GXAT3PeF#F=(=8C4Q)+2c/7^GK/B)2:X(N^9QLfB/;
)RV.-OK)5T6[dM<X&.C/^BfBf_Q2gbZ9PJ-P[dLL:?^<d>19#Lcegb2Ag:)[Q7Gb
1I^T,-g2a6@C^+U:^?M_FYO/UZ+B=,]-aA_\\4Xa;>d#_WKBN4,d3dBM9.EJDYQH
Y3]OZ+Ue[(5Q@>-SP3+Fb&D&=_^a3PP^>GeL^TUZ+O;CF:&1dIeOJC+A[O#Kb-<_
J8/KDUX9JN4O#c/<[Q81aJ<c))S^K<D7_)(a9CE/FO@/UaAgf9E9O=5gg-8WMV+,
(\Za[BEf]3=U(RIUUQf._NOP\N3)fb[fGF)7N:+HR5WZUH)SS&BFAf1WFOOE0J3g
;0LA@QC9#^JVZT<Re1/7ZNe\_VaIgf_87d(K)0N<Kg8V(MER36[3R<7^8S993QeW
HLgSX&#.?YBZR[dV#Y-eMf_V/#LN0T\Z;,gdVdD=/Oc5TI<ICJQ=3S#67FE1H9XX
-<feZ<^#5@=/FO)MRK.R.8<_0S3JLA?)1ECHOH4/Be&F8YafB:2DMGd#(K2#H)5)
-]8-ULE=e9-8&_YM+2gVC(1KFeM-.DF?W0W2d4<fR?@7N5\<QHK^NYN:ZCefTLU>
;1:519RgK.L[b0,(5e1180YD2Ge;+8:KOL3IQAL9[E:/+#dE.T<X]L<D,ML(KY_V
E1>Q(8f6=g;^.N\0-F:&T4C]YTOO+dCRX]:Qg@:DYdTELV6\A,g)S3;D^TdI^c3U
K[B3>-KG2Oc_Z;5CTIf:4.+9.Lf.\#1YI0KG]53//J^(7#DKSbV(/P<:Gg-HWV\c
)B7=#7&6ACWKSSIY#D;Y5<^43KGa=33VER=fZf]]7a4<g3=U10/Oab9K@D7A)NN;
\Z>1K,CYd/;_4a0bFIY].FgX/:T_S-]C[d4HC+0g0W3#:3]5g7(HO?gCWX4SK8fW
0Y<d;=Y6&O]D?3DV5UYL+eC0IK5O;KBHe3^D&RCPWT@>Qe6SM\MMJ56]SVJVEb(F
4L\\3[JCK]NSTFg->N:,7@A8#d(MV=>F;D<D?=0E,#__c(H&ebQdNGVUJR-ETWS#
/64=bGbFF3bBQ?K-:7T4f^]Uff:<+UKUV884[\bC+0MK0XG,K]\.RS22DTF0XE7;
^(#98b<^Q+@-0ZXWX>E2LTFW\bP(bIFb&2C;OWWeLH9g[f-H[<YAeX-(7GS.;3T:
53GARbBg8e;Z<T#EH]?B.?H;/Nd()c6M\6?Nd.7INXBG=/((E5cH&(ReB5e0.bHP
B[L4HEKeZG9K6QYKZFZN>N4MHEQOR6Y@,J)(3GUSF90CZ?/c_A/E:@90e&+LTEWG
AY?3>J9/Q^1.0MU6]E^A2<K5\GF5)8Y8DS.EdT,(;40&\IMN\9bDQ07fd=]bf7Hd
+NV4C#21^dLYM]GU1A\XD(QU09WeY3,R3&).63&Xf-)QZL#]X?B:.;=JbAc5E<1)
O7&f.+Q3[f2A,?1>8K2L;U<X,@E8#g#W<NAI?\\g\,P7MWJ/Ra>fNGbZEaIHJfOF
6CUZ#>49O;/=b>B976;_(ELc0Q>ZV^IQaV;#A+6J(OS^C&WILB^AD,ZcEMU0>STB
#8NC3HC3JD/,?F/dL@N##,.M:>CYE/?IVBY@aQfRg:>aG]9NX;/>W&CX8WF42RO8
e9M@GU23^^Q/8]+@Z^KN?MGIPNY.PJRFRKN,A-,3<^K7LOg->AMY:5C)MC36[G/7
EHVAT7AQCX_>_W6\T5H;Ld0b3.2Tfb^D\HZWCPIR\HX9@<X_:_^R?91?a+c82LND
J=[#eJ4E\01+I9KB0&3@IC2<7fAO@QJb1PGA4+9eUfQ8Q7&OEb^.g0ZP2?=fFACO
gQfK65HcQH=[;f/=c(I?b7bcXK2d:?:G::SBGAV^GLI&eWI(=[I+;O[P++(0]ES(
YH9^:L2NTDdX2O4[NeIb9N^#c374dVQbQWdHO@38<\7M.PFGcdVWaa[5W-gAIBO\
=5T/WE4.IUE=4S,;K9>>H+DZ=Sc_6THMLD6PZ[E9[H_MO5A/ALZ/Q8;0E2RB3,</
^L0C7g7IS<TFT9@V(&e;K,^OCHd48I.<T&Z9:.@[C2-UQDA#G0J::\KU2(OKNA2Q
=Ig1JCNQB7?RUW:/Ib&=)=4CH9ecSPHCO>4U2/>]A:SX5;bWUF96N\VWNA+fT]4#
N_>GF5ZV2JB_HF_S-:O^(L]aHWa<\-P.&\8.DW1M>(=P:MWI5X#H,ed,I2e#3NS3
T/g\.aQ6GD^>+NRZd:?.cYD6OSQC&MI(^;P.DK^MVC,.35^B9S6f\Y:b\<RYME13
:=5T:<VO;QBXTE)DP_V7XV#X^B;DJZA5_>3)d70I&fTP)Y81@D_]P#<bSFZ(_<FZ
S-E2?O.M5IAWLV)=C6.c=1S(]=1dQc:,,=L4e/VR+J;KIUGeeR^QAcED#/PK&a0V
FLW<)8XXVXG9^/&=]O9Q;/<c]&f:_C@[>If7I2:E==+4];,8P1.FQU(4MTb/)>&Y
]GB(:.?/81>d6H1<36F[_&AeD/gQYf&,^RSRKE#Z6V^EV@UYP:<0-_<NKOD#PXeD
S-[e29GM].Jc8427AcO7d)=;;7PT\bWUZOTS(DIUK;RUKYPBfeAb8Z.)b,;:aM5?
T7.@_N7g/?e[-[N347\gUAUE+,TA>;<8CJ@QNfJWMYGP=@F-@@1&Q1P0-W@C_AFW
C\LW0c^X.>2Nd9#MGObfeJ@LVU8MLGAX[78?3G=T_-&eGKLDN,])Y:DF82ef;eH?
A:K#?TJ0DfMb>YIQOPF;e+>;EHIR=PSWc491KYKW8b(e=HL3^XHN8(=[6Td\D&=?
f&MdB=Z@@,LE7B+.IV#F3dQY8\WUKOWKX9J+?8N7G6fQ#A_6^aC=\[19K:SaJ^:I
,[[#K5.Hb6>_D:OX]XUCeYB2;Af=SO3<GdRJV=VRaC>NHR)XY6cL&:?N6KaQd/gQ
NEF)(\g/gfB5,,OD761G(6NIUMcI.=>cIEV.&ba^:3@]VE6RZR]f>T]H;Y6KK@7B
Rf2b<<CfaV#^EL6FgG=K2WH^NM>M.9L@]UG?c4[gIM->@>;9NKKBBASRH=aI3_HA
d<5A7_OF7ESM+&]&[HbHg3+@@DJfEI/]K+bY_P..O_Q0Z9.L^8fa,>.SZFbS.80V
K&gBg;adDT:)ZccZX)b=MQ--9)F@81&\])7WQbLOLVUcMJ37,XC[8Jf+^S7E/<\0
_D60)f^^G-EMF[J1>0)K64eWQf[.d7eU8f7/T<[4J-;Y#4+-YRZQ,?,&_f=0HR:&
.U5WB8^\S3TdL)<L3]LFC.X&_[0[719:cFD&8GC^?W3SbCN9FX(DccM(B5\(#2O,
@.L@ABVV?c>aFa#(eA4aA,c7S9&0.4(9d+@L#<>]SG.Tc_859=0aGbBWbEP.#e<#
HM;@^8Z]#>0YZIEFX\geH?YY,f<78G/[Z4AP__;14^7Fa<1==X,?@Cb+MD9Ld#^&
X,@OOOD62A5@1FL8W;f-MT).F_NY@(3[H<^>A=I29<[XdS^/4g5f(g,-37#1[0:2
[+4A]9>E31B8A2&OYb,@8L\S1Ba?#Q>0?^\STM3D/,2LOd=ZfU)D81?6@1<XJOYL
cENA^W+G@d1fSB^.CW]<0X3.b7eaF,_LCDd)^Fa(AcM?8G]XLWT3Y,K=-Q4Pa0G.
0SL3-;)6f4+74H[&;^]@#(_LJ^f8JRCA_.8[NAU0BWV@S5KHFE76Z==L:_\(;ZEV
.ZMOV7OM2N8FW7HEDf;WYcI&5Z@R1)GII[&SWNXHb]UP.V2be.T;8W?J#E1Z#27-
&K1NaSc)7C98GV1@1BF:A<_U#29eEgMJ,/dgQaGJ;f=84ZYEUV,T\33HZ[6C)M#?
9?6gNAWMWKI-WGX-Q?g&6=,V[.S@VAWK<)]9-g257&R=b\[Jb>Tc,+@d)_)=_>>9
@3\FGIAKDEDH;=9>70Y:7A=OKL?-+Y^NED+574P8Sc[ga451Z-ffN-XR=aSOTX;E
[>+:W0<CgfG.?8#]44C&ReRUVF;D?)WURaAURQa>0>MH;.+_1JA9&@ebMDg,5DH^
V?<RN]<PZ#Q>_-N>5D],?CD@54;=d6A3+_,L_LO]1TadQKYR5YQc9O3JY4YKVA3.
;^c42&4L6@c4ZKIY8,\J.=9ad\,(EN1>ATIaV8Af)aeXHMGY5I;N\=>eR;d)@=U#
^cI/M4UTOc9G4Y8fDac\95YDQ?V([;WdOOY&#+7@]/a_XK9@+@+EDW2#]/R.dId?
9XfNF:?I697RDOR7Z&2JZ8C0OH<W(8DJ9UC^bY)MH@c72d-VT);71XXaYQNOXC/>
+VHZ0.==X=b^8/RA[3A+@SI/,SN@@@>N8Q3(9MBIgS3gOg]@N<CLY?H;/&0U,Ad,
b;Ac?X=(;:&7D8<FK&5R]g_NPPKM04X,dT^=@J?L3Kg:K/EIYDX#5PNcVCdI@2ga
VWeS5)d+MN+8S?#X2(1fT/T^=[bgN1eM->2NH6YIeB(Gc(&IQ#+T<W73U8NLZNA5
8XLR/=3POS\I3EOIJ[J[JY65-=A(WPY\G1dDAH_0L_61Y5+/)IVIJ<9AfPPHRCA=
P08A:6RCb+\gE0?7FZ(=(SUJQ@fFa8B6GJ=Y5W4C;)/LQ8#cT9T>@JNXC_VQ_3J4
B&+SGT>ZWKA8QfScdCO0cDJ,^=e;J]Wf3UP?>&Kb1bICJ=2>BUXa=5YVcUb39AIV
.?4YC5_?g6NL&7M];IMbE;>:6/ZMc89)L\&f_bGQ^=Z9[N(T4&aDXA4YDdFTDf2S
f?eMU85FPPZaH#</YT.H62,b+F6]<J48)f[MJY(,(OF]FA8XHL:6e5A.LM3H4/K6
RU?N&9EdIN@)ZX8#7@&cVQ5[Sf=@CSW-(Q9T\?dI?8M08YK4T?8]F/_e==)>4,(M
CCc(Z-dc;>9T^g0aK=Q@NbMdV1@AW7g&;.Fd.ZC_;0J3,E:(BIAI[]E;BRJ_L=Y;
-2TS\6)>>L=,]D=O_=(F8gf#662A)JaRDTMLR:cVB^,LD7[IMLIH\/HK:E8_C)+(
N&0MHSc:I5f3ZV-90?ZN7#LZ:#-f:APRXX?B=-X+TY_L_7Pg0&C>6Z>dPbdgHODU
-M\3+d13DTb[]>[c2MVTWFA;D13<==+cQZB)M^74,10B:.?BD@+WO3fMS-VNGS,+
>b4HW]?#87FRWg=<UW-<?SUXEGJ_AZ=[VVLOdO3(X9.M1fcc]LF-#B\7EXAJG<S#
[5QW4eA:9-U);#4=E68R4.\RMA9<RCS^9-9,Ec]G2U:11eF2Y,78BTVZHM37&7FJ
PC3K\LMJK.R2Qe^^H;>M&CQ&<1[ODbTgbO0Q<e;+b0SPILO1:A&af[YUUd=Aa,5<
G8IGEYT+RI,07HDL;Z4Q8J>1H(,<Z,Aa8]6V#dZC0T:B:]8D69WJL4BV=3Z3d9?A
EC#OOE5MSL+WY0LGCC]LB)Z22)@X#LOJ@9J4;:@ODe#+6W\NE/XP9Fg8b8?7N#gL
>(#gMDL<I&19eb<F5I@>ZT\NPS--]+gJOK[A:&W[SAg[V<EU._T6=SP,Y>7O9#^Y
Q?)1.dPQ6JFC-dR&]G<N4/W)F&@4fG+]9@5,7)NV.RE)4YY#[BBa.e^7I=)/W7^.
_]\D8dW09L+deeDI#C4b0,5(b7/9=#-N#OgSOdG,MVdf2\T4.Zc:NdJ?@L@=,NV3
7=HIN#&+487_e5,H&(V?3[LZ<>EOF(@7:48Dc:gVSS27VMR2bZDeWC@\+,1&GL1?
e&.FTX^N2aaY2?>#Z1K-O?SG@.[Tb:4cgYPF#\[/BVP@3J,\##0/.(SYS4Z.7L;c
YGUI,UAOTJ?<YR=6Z8-U;JALF.?E2:71\M6EDT=FY[^]4JMD-^\1B/;94R,fX)/8
:c^e<56N9D9D\(:6)5-Y<8If@)J>D009.bM@Uc=?OFa3>9GN<A:YX^XDUSSEd1<d
^d]c)B+:0e,VE722,L]BF28d5.e[L:J3/.V_&UdLa<&/J95[C/6]+]>5P+:=G;LI
XE?G>PJ5/D;K3[DF()2ROJ<X27GIGZ/#<59(>C@MbSC)D&X6=\:3A_,NUIS>PS>@
<WYZ_\+6]=aMa)]D#9_BJW_H<Ye7a#aD64Q;>/=7[;4?RKQFV:M9Jd3GYNZH:eWJ
)_,.a2BMA4,27B9_d+g7AG_QXW-FKRWgd#QYS;#[gN0dWUUDg;6g1-]:Y:YBC\,^
>P@EV?(,AG_c;,PAS)?)9IQY-L#40GS0T?5a\U8CMZ)cTaYF96E>NcD[6F24.7XY
3ZRZ=L(HJ/\c;7R>P2[ReQ=:PSY)a_8,//28YCOEcE1:#2J(f3?[cTA]4>7D)F[]
b=-K52ae1R7[R2Of:\6LT+6YJ,OZEb:4c461I8TN.T)6g_9G8\^e2A:A.]6-egE6
Ve&<:][?ZeMT:A,DRV[?e;X+)TC?I:E-aLadU&5gE3Q?5^X4P-Z)Y6AM#<fMU.]=
1O=9:,P>K1d0.KQQ\8_K&#1GZ:Ca5.XRE0UWNCQDdZ/\)SO[.\H?HJGWXS4/)&?P
#E];F^Y:b9Y53-0509R_6^-;AF([=7^?:C-LdB&2.\RHb7GcGQRGWfdGT?,dRN@W
39KX+2Z(6+J=4)J:7dD0_+-KRf&43cZ3Rd_aBf>DCJ=IfSRVO2J<XNOKMa1][Ue+
CD2O?#)afdU#I],(B]9A3JF=BQ5XX4F2^5D@SMeJK&\0-Q0\\(fR#[A=ES+BgVP2
eNdcE_4__Y)?7bQ&-2/8KVfS^MTa&/8fV-L,_Q7@aT\4eX&\QQ?.BBN1X-S)+&\L
A882[-RR6WT&?]d9Za>#2&2>K@H-([Q_3+Z?[GS]7T5J9L(091@R)BB3/gZJB[cI
;f6Ag(\D65g@K]1O-F6ZOX^X.X0c<8)F^E)?)_]\2W6XG2,d+^J?2Q,ag:;IA_@@
RZSO;U>PfQZ>-N_\Mdd;HEM=KI8fEPC+N[?3d(_b@c8d3[Zc=A#ae1V2Z5f>3DQ\
V?@V\TdD<JK69:[,77HJH,9)NUb8;b,-c?d8X?e6WGa1EQ[cJOO4WPAOb7F014-Q
=\QWFT#ZLgLN&d]L#_PW7N83ID]Y6RSN8_8FGS&g2/dJV\ABIf;Y#B8AB#[;?.fQ
:]YPEYR@JfNR-R]G-U,]<=TOK3#:&6X^57-:;@QOLQGIa8(,c#2N#HINWaaQb1MT
W/W)b^^Y]<,6)QG0)K3M1d1KTYTcR[b3P+0M7d8<2&/cOa>2A[:/f4dJV32:)M^2
]4/QN\;Q@:9/Nf3-@Q[Y9:R2HPQY;UeJTa]5Y+=(T-.?=WH?K][IGb7[Q;5MRL4c
#NSQdJ.:6-ee@]&(g?-2g:MNJ.YBM0#=P/<M;].-WbcR?(V&e(?24QZ#\39:g7E;
=a\?\]/O)UFD(EN_N@VG)AXbZ0UNaZS10OLD>GTSdbX/MJa[BcS/GA<&L]]_=?g&
XE2._29R+2b,W;1BZAV&\M:PedOE@(,#W]@E)2;PbV5^bT:[AL;,36?6gIL#-HB=
E2V2EZI@B0_86b8\BMBYVO+=UQ+BW)L]&:c/NKd7df5W;0AXdZF9OX<SWBfc:.<=
R\PSWgeH.LVNX8Hd7&1Qf1M3TWT0GS-P6N9G,g/J9<)_XL4>FP7]]N=S;<1EFMBT
8c,>Wg:64.2e3FZQV&7A-(7PcdD86XXBY61]a7[OW9IcVFfYaP#)C)>5cZY;3>U5
KEWYTI085V5,>JQUe#PJT\HU=Z+,(P&>Z=XXd6Ra-W]1?Z#:QSf6\NR,:;XU9K?\
63FVE^^W.W+M.[Q_3M,+ZRgUX.\[TV^dSg+VZYYR[Z]8PCWb0/FQH?3_EgT/>C5.
A2gTJ]]8HW/.JLE\T[QVD/YTMU0f2b=I?[-Q<3P8Jg?>E5Sd8e>A8&K-_.1.(8;K
R^HSX-K\:>HHLH:7/?cg<7G-KGO;H,Z&L):6ADVXZX(O1;<R1O8O&gCE@UPHM)(I
4Zf5T^65G\M>;M:/-S73F?eB)X-B8@..A4(e^F\LE6N:CWO=-RLeDcH.S2AUQ0,0
DZMdX(dJaaWQ0CLH)d6Ad^JT93I/a8QIZ6.M#WDZ]0de#\aBceG#T^[cf,ZbWY0f
Q&1/9)H60g<3U,NKO)c64\JT1$
`endprotected

     
`ifdef SVT_UVM_TECHNOLOGY
   typedef uvm_tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_OVM_TECHNOLOGY
   typedef tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_master_transaction) svt_axi_master_transaction_channel;
  typedef vmm_channel_typed#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
  `vmm_atomic_gen(svt_axi_master_transaction, "VMM (Atomic) Generator for svt_axi_master_transaction data objects")
  `vmm_scenario_gen(svt_axi_master_transaction, "VMM (Scenario) Generator for svt_axi_master_transaction data objects")
`endif 

`endif // GUARD_SVT_AXI_MASTER_TRANSACTION_SV
