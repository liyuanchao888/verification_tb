
`ifndef GUARD_SVT_AHB_SLAVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_slave_monitor;
typedef class svt_ahb_slave;
`ifdef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_slave_group;
`else
typedef class svt_ahb_slave_agent;
`endif

`define SVT_AHB_SLAVE_COMMON_SETUP_REBUILD_XACT(curr_xact,hmaster) \
  svt_ahb_slave_transaction new_xact = new(); \
  rebuild_tracking_xact[hmaster] = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact[hmaster].is_trace_enabled = 1; \
  rebuild_tracking_xact[hmaster].store_trace(curr_xact); \
  curr_xact = new_xact;

class svt_ahb_slave_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                            type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_slave_monitor slave_monitor;

  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to slave common parameterized with slave monitor, slave transaction.
  // For UVM, it is available in the base class ahb_common.  
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_slave_monitor, svt_ahb_slave_transaction) item_observed_port;
`endif


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Slave VIP modport */
  protected MONITOR_MP monitor_mp;
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_slave_configuration cfg;

  /** Reference to the active beat transaction */
  protected svt_ahb_slave_transaction active_xact;

  /** Reference to the current active transaction */
  protected svt_ahb_slave_transaction tracking_xact;

  /** Current beat number */
  protected int current_beat = 0;

  /** Array of current active split/retry/ebt transactions */
  protected svt_ahb_slave_transaction rebuild_tracking_xact[`SVT_AHB_MAX_NUM_MASTERS];

  /** Reference to the current master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] current_hmaster;

  /** Reference to the current retry master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] retry_hmaster;

  /**
   * Current and previus value of HREADY driven by the slave.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit current_hready;
  protected bit previous_hready;

  /**
   * Current hready_in signal value
   */
  protected bit current_hready_in;

  /**
   * Used to track previous burst_type for error detection.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected svt_ahb_transaction::burst_type_enum previous_burst_type;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit active_tracking_xact = 0;

  /**
   * Keep track of number of transactions since last reset.
   */
  protected int transaction_count = 0;
    
  /** To track if the hunalign value is changed in middle of a transfer */
  bit initial_hunalign_value;

  /**
   * Keep track of the addresses seen on the HADDR bus; Used for protocol checking.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] previous_addr;

  /**
   * Keep track of the HTRANS; Used for protocol checking.
   */
  protected svt_ahb_transaction::trans_type_enum previous_trans_type;

  /**
   * Flag indicating if we are just comming out of reset.
   */
  protected bit first_xact_after_reset = 1;

  /**
   * Event used to trigger passive monitor signaling that a new beat has
   * been detcted.
   */
  protected event new_active_xact;
  
  /**
   * Event used for handshaking between common and passive common to
   * inidicate common code that current_hready has been updated by the
   * passive common.
   */
  protected event sampled_current_hready;
  
  protected bit   wait_for_passive_common = 0;

  /**
   * Flag indicating if this is an active or passive component.
   */
  protected bit passive_mode = 0;

  /**
   * Indicate the last transaction start time.
   */
  protected time last_xact_start_time;

  /** 
   * Flag that indicates if hready is sampled for the first time.
   * This helps to figure out if sampled_current_hready is getting
   * unblocked multiple times in a given clock. <br>
   * Used in passive mode.
   */
  protected bit is_hready_first_sampling = 1;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked previously. <br>
   * Used in passive mode.
   */
  protected realtime prev_hready_sample_time = 0; 

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked currently. <br>
   * Used in passive mode.
   */
  protected realtime curr_hready_sample_time = 0;

  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;
  
`ifdef SVT_VMM_TECHNOLOGY  
  /** This is required for VMM where monitor needs to know when the driver is
   *  ready to drive next transaction.
   *  This comes into picture only in active mode, however, the slave monitor
   *  has a handle to slave_common. So this member is added here.
   */
  event          beat_level_transaction_done;
`endif
  
  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KDCUsBCgo9Kl/++cDs5YqoLnxrUNq1qR/bh9aVIoYgV5Aw4dnB1CF+W8DTepNmu/
Ek32eYoeubwdKasXIKPEf2Ab1EIrUTtv6SMHKweh4ruJTmuslBMe/NR1qRMnaESU
Z9TulZf0hCmM1fRDe4zWzEAC1Oi04NBg0oDLvJ6aBfg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 644       )
DU4TPMlfaPJU6XVQ8WsrS6fAfLnNtLiFstwcq/ddMUU/kovRwJMvhkFDvKrV/FrN
b4jC8FmOQ20ZXJUxvLutZjI1+Jtl5rWkIWsis9sQa44oD43t+gBZeM5cGD6nTUFU
jOZAghzFBprCKaxodrZUS0PURv5uBEIVQHgGeucFyGUA2L8M7Lm/wcpVxDseLnMm
2il9ZU2zaPPTNENa9qw2wLKnu9mTcxdvb82b2sx1/awbpJTH8gHVffk2FJ6buzIQ
oJKLJKEeGw/c4KCWavOuqYl9pLqt9+PHBbXBEJ35Z96sJnQn/kovejT1oAcBA5ND
kiZriHLdTSE0O8XRkG6Cr8Y1gADAb5mHzekWaJa9aR8jNlzuzhRJPAfn1bJsDRmc
4QkdG3glFx7XdFqHz4v/jqY+QmJDMLJFCH/wN1yKgRs9pddmasN1My+UgWoXdvWa
tm3sF8Jo1L0tkPA3m9Un/LE9zDotwe1KuVDNU+9qJbt/eVeE96ZvuncuDgqLuxjS
OZwKy73F7ovSEfjTTkIhmIDTdu7OCprG5zYKUse8ZJlqj0D21PnZ4OlbwTm3oGYZ
X3+zn9MDwNxu4X6Hc0RFz9b/M2KBTtu+++Y4YkkWF7YwhobkjHUK/zUU1mry56kI
cVZXd4HTnHm5fxOZu+uxTHOuKX8VWgk6JXR5ClGwJKpdBge9rzBttkoJ+6IABgxZ
fwWzVRyYYHybC5B+aWH7rV93/h1/NDdnP6JDjOJPHRlOy/swLk8xuyDcpykIONCK
sgV/0GBCs9HVRdggW82nRqu2gMpBMVRnIDgI6ymf7ITG6ODLyjjOP0KUIbrrjoZh
UCXH3NQh6FRzN3I2RYgGOYkZozkYvXi9lJ3GEvtCxbc=
`pragma protect end_protected
  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();
  
  /** Monitor the signals which signify a new request */
  extern virtual task sample_common_phase_signals();

  /** Returns a partially completed transaction with request information */
  extern virtual task wait_for_request(output svt_ahb_slave_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_slave_transaction xact);

  /** Monitor the end of transactions to drive the observed port */
  extern virtual task complete_transaction(bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] hmaster);

  /** Checks to see if a new address phase has been started. */
  extern task check_address_phase();

  /** Writes data into a slave memory */
  extern virtual task write_data_to_mem(svt_ahb_slave_transaction xact);

  /** Virtual task to drive hrdata when busy is seen */
  extern virtual task  drive_hrdata_during_busy();

  //***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IYAVeJnGkvFu0ERwZ5WI4b4LQT01QXAouJliG66wABIKaBq07/kwVFae4UMDpVvV
iFahpnJJdAZPL6ZQ0aak1cLPgo2wv+a/8exi1Mx1enfLSorAfPR8tsOVBDbe+ymc
8UeC6pHYT2CRD9bkKuSu9mVlsNEJE9hnlIrSVvv9LR8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1906      )
lU02e3KSBdgcUhxBOd9Mpl4Am6hJtSZJGUENvNVeg04CwRUUujYhJ6OuIeDlqjVc
6rQNCaBPr+wEXn4iHkT+OQD/CFakVCX2roDs6Vzeqtrn1FepDBQH01iUL9J9fwxU
OVbe2SKfUfzY8V8UQN/KonhkaHGN5YRVuk5vdkTY7Dk7Y38NwCd8nuSpTRJI4oTd
KfiALIy0H9R0FGqUizYEgjR9eDsKWy3l9mXszeaxMTnBb6KZlv+cvUy4I2uvMwl9
FCMw56sr08iRY+VePc0uXV2t/Pyb9eyzG+SHHSndhNPHB5TXWiH6069eebZ3HX24
cCADjAFENsSiF3b7YE3QNk7QO69nlZiRYAIrul8st1WohoXKvfl+mkTxiekXMnt+
Geu6iY11oFNVinYj5iMk1wDI8q0wopcLPAXTZAOswacytG6NML9WlfDG0VeNHrHx
OEt36c3frRZKVbD0s/k1Vl/IWDc9eIG4nGOVLTEaJ48TbjSWNMU1rvzJhDi3l3ch
Rbus29G1y4YBNesar7I6LuASgr0f9bjV9JvB5bA1+aaSoPb8GAr4dbcDpOEVD0/a
82jlLdUbtYS+naVJiTs56f4is+CrSdW0FOSYHrCY3UCK9M/WKjrz/8OJwOrXGr8O
cpPsZT8oSWrtdh1nstQsbF4taX2YYV3tuBYrj0akqMol3mESJ6sXZ+NyOMXlCqce
BhcntLoy1LUVcowrhY2szE+UxUgX2+9pdTQUQpY/gQw1nfQ7RN8LNC5J6WkiepNt
EJPqEnmd15mCA1rzZlelqxF4sP5kg08/GhlFP+W+nuUdH86T3/yfV8d9vYO2Er5K
0bltUqRvlDpS/51OuyO86qTBROyS3bZq55SCxKmnf9mx+OCw5mCLKAwEnr96AWh7
4R6DeMliLkQZ3s6NwcgtO3LFnC/dAxYfz55+9hFLWlVBEmf96Y8kLw/gMlhHASjz
gEEpibk21xvzkrOVsX4TA36ubaOuPVnIh4UBUjzHUTCLLb4AxzWHwDtHDHNnNuEf
+F5pfQmPdkVmTQ+g4aC6feJw9iq/FTvRTWzeKAidnBvGepjgTZ+3AAzmO/J2XHnE
/C+zW7G3yCwMlxP/yUTCf1VUG5UX6ZhJ9AqnOpnMwBZWAS6j25OieTPhhxR6wIdu
3YXfYXx5ffi6uZRk4/3B6BA4Uitvx4gGoCz+xb5d/X44gmL8wF0DQDBLRiotnswx
I8UHsCm6XJjMZfmmZ6aV6PoE6GIkW8HTExjC341yfOB0firmI6v46MNow9POiZWb
i9qCGQCSfAcZbfipjOMVqjyqlic0qgGA0VbaWIj5Wg/BLGspIepTcHu3x/PHEkxc
6IsX/XNvrFbVL3I2C43YLMIZh/OTDltrH3nwoF3kjGiJ8BdPWmYAnBjOO3dEfymv
/ebTrjjXuQkDv6HBb4NUG6HIM/qgP8GyqJzkF+odXNw631w+lwJkL9hHaCi5D7Vl
IcQ3nH6bVy9WYOMRfhrtQM1g8J+hWflNFOq5BkW4ANrhG0AwkXDgy8Mx6/2y2PO9
gf5fiw/qboWYz2vgHKuTqoPh61CNbF49IHf22jx/ZCtOCOFdv5nXP/5TbYZQbHs2
+ufCRpYhoD5WFSKZNuTzQEyPYbcJ31s+3SgMOwEO0d5w2UFgbW+8Zo5X+vq6TtN1
Fi3Xt0zcKw1EFfmdPJ/f8Q==
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
onNc2P/NsIP8vA0XjKfEq52TSOV2hXq57fzB3NrVTpFcVNtgX74vIYHcgOEVuGCm
QMvqAPgz6Yq3XeY8VQyPGUsQy4aBOJ6Yv5rudeWUMR4Sx+DPzElGDWFPjH6OEFKG
nd5tcTiPr5dJS7+w7xJp3CzmhHjUJEWEpFvzVYYmAiM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9102      )
CZ7e2ZZ/23SUKgAEALKGV7f9f1+qanL2jpLCKgmbWlcXQZc2L8Z8WCE5GAH/3CUg
DN/a44tcpu8vICezscOoi+LHf95XCJDaUp6JNeqvSPgjFeiQczgFw3LFlye4Nj4I
0k9w05KKXF21mK69TnD/wMozBWn7mmhuZNrEbr1F+i7yHEAkln1smHA3QersEHk7
ZusjZA2N6OAOvOznKm+LDDhefXIGif+ypFSYwBzh9J4902Om8N41xeGVqV4T18AI
BUOiWtgbP4ZpAKbHYRFZC1i5CYOIQnYPIcnVMPvLE7dpTUh9r8qwGmLRvUIS8bPs
XPaSA27tkVgM0ERyAwj4I1nifpYqfjQM7tLkiPlY/oX9YjOILVccuzv0Bbrx2WdR
XLChgkE0KigqhCvbQ2lFj82TWj2TNxkMIgNuR4zBbK4SayOiMq53p9j+h5+hvOj+
YWJhPc4krpJY3a84xTr0oWf6kqD1Y0EuPOzxwoLZC5CtiQR9AlZ7usfwyDKU4u5B
6IImqn9qd0vIPAiD5Lgsokhy+zkOpLxJ27XGlpjPGnUSnrVSChK+kIf8Kf38nO/o
ldwSpIDRSl0oaoXbo4SgdYNilWhY6isXOYoJulWMAUqxEO0DTo60JnmrTZksrtBr
0HT3cYkcA7Q49JvLjwyg7+pTMKG6DkGMDi6SqGDviQAM2huQtFsJMiyuicjbhZGT
sBD2c8Uet4vOb58f/Mp/aq0BePZgugYQ0nAz5T1PYE8zz/GjApPRGIX2lsFTlw8a
ULG0XRLQBpYCChrrIMtoBTR8NEu40/DqaKvpGA+SZtWNG5BXNJon0agBg2T9+/9t
192SmT3OTIOunLCu6MixW8BY7VSCDShcdbIvTzpbwqmFHeQOk5XVTPvNQmlRlsM8
oBqEXolMDOq9RiaORp1aSA4IdVkM5FhvZp2mE3t2qAhtwDSWG1I4yzNSJ+otPT1I
krSFOhd2sbTtSoaczCILyJf3qo0mob215pOhZvzegIMTkcxKJiZpWhdz+bXGopR+
FSD+yU3wV/dR7MWLEJl4mJUiQcI7Mi+Oms5lgfRTCByal9tE/cykqVdfkYlufrdC
0DPyHb+ZNZixouYL3qsYwf9rMno6SzHA+fp8/GB1w8YHsLwoqKhijCke9B9OsE/z
OKwV7e/s4ON1O4iiVt0O0FbWSClpStea8jKNsBh+43z2PaTf7wOy0TIDsZNlNbkU
8ofXOZgxp0diJQ1sbTZXle9aXcbGgR9InckCUO9xkOi91kA7BJqEtnOPTY/sEzxR
oUkuuXzdmZzdb3hXK1RHXkXJUVsUQcQ/M9FRbvxukkOEl/aYqEWL+9j0hdfRHiqQ
ssrRP/AO/HaONTi5ylQOD2s/EcoTAJ1MeYeL+hvWhBRDUfqcbjWhma0xn15kWuO5
PX1yB7YlcfkP9uOiz54tjbxlvq7NU3O70erndmBjWBIWXZCfn1JAZ/uTBoH6FAWH
8LTyl87zd0IoSOiI7IrwmcTGxP1c5F2clx5Sctqr2pI/CNls1B970e12NxWicWKK
MxxWfGQoVNz8l6XTfjnPvP4jEcyskdpbM2e/Ov7X/X2l7oZrkMffvPFSvLlKhvR/
aNHjmhbj9HpIkAJEOQ4UkATE9qffGdC49J9uhNU8mrpxoocUM/9P3Fwa4yBtFbdU
R+pY99/eEHks3GEvyhy6dd880dh2sw9YYcqdK6bSh250a/kqsG9B38ynb7lE3GzW
IpUaS7mrM4LMELg1V4vHjip607J4Q3dxHExtOjatESvD7Ba9Hhnunp7eRWy75FRK
KzaoeZ91I7ttPyg2Hn8of/X9TKbiWky7eR5w9WhxzqGrV9XcB/w8JU07hUrnf1wp
FTlwbZwAkV32ULEh9nKc6Bb7Xc8SMxSwm4DRq7r7gDAi3RPxE+CAFevNg3vph0tG
pSL6B7dTDMubWR/bTXtGkt5c5BgxSeJRL73m6OQqf1PiV8OBFB3NhI6I8kqsX8Tb
abSMEl5Py4FpJryO87Ft27deU0toSL4gEEKZi4ERqd+6F+BqG0v3gy4xcAV3mhQr
VNNoY8fPsMDFsFoyadbThl+K8XgTD4t/RFtctuuHI1YPXWzIh/iDJBvp006VG23l
5edj8pMpe5I9+tCfd7QQZUWFAAEish4+g2haBGAkR1nbyQ565gVgxFP5FgtB6EtW
65G95/Pwcwj/3U+LvVySpUzVrtEFPmRFiL2fadq06Zz+jGfjjhhL8iumoj6Ldtwz
EaxxXWL/kJEb9gbtD/ihuG5kFxBHV5YZf5/yjIwCAt2QuFD1KMkj3rwx7oazujiw
eNaDjqJss9HFNgm8eOeELxP74rHnWVOisDlCjyBUzuxymamKlRx2TTJghnlLx+ki
KtdBpED3VV1wSak348lDxI4EqLrWILHEA7vUD2Nef35OpRwaBEDZ9UGI/pMIXq7I
6l4vz/kivam+TaKlBzz1eoF3JhUt9w6gg3xYEf3jIGVH1FGoCEUX3CFM1WGznEAM
iWSquXPJ/+uxp+w1/kAMwYYschrUJH9wDYINbhe+U/T84d197LNwQ6kJ2KL2KurL
M2H8MgL/DYha2nPBUMX6ALvwReJcTvSzbOLVIaHcTrvhzr5MZwEJgmwo2U4DOP7Z
yErTaHmnMpJLLJJfwIrzzqH68af/HN+5vYieD2EEydyrhzGbpizFROeorEdl8JZF
Orn/qwI+ohw1Cb+3mWSQPvoPE59TsL2faWDJIXoGaSexTjXyTAHkH5uBrMZiUA+z
QDM4ZHIOeis/pv9eVz3RcYWFWcUELSLJcZJPpW+sC20EC6ksPeWAU3cT4GbDkmCJ
cBH9u1I14wedWRmeLPaWRKmwQiZrPOnkhLbIpWsvbzl9+LbY1wZGE2lYm1RlsUc4
SBqsr6jfjnUNlq8l+B5BIY0pYLLYK6GdVjK7+Jo1REknI8AaXRY4LWyzmG82RR0x
t9vgB/GIOqBWE6qKKK/gNf5Px+o/1pwebdRGTViPbmRwqYc+tWgag635VZVrZdqq
QMvuQHctKzLY9tYKqYEqVa6Ha7vCa0fGIp/8SjA81FYrgQQolLGInzN1TJonGDb7
ZzZxWnrpGWTezc8R610l4uyU2CHPfCk6J9MJB+/65qTHyF29ntoEL6g8R4qMlrdb
t3QN3ovw43K9vXHb2+0fN2a+h9Pd6VGEMa33Laf5HGnxNjEhcBqMHOC15/l4FAu8
ryp4q9A0WGXe0umchyEY7D5wV8qWXTfk8UOg1V0JgDFSQY8pxLODU9t6w5eEkD2b
I5PMbiAnSHZYTkBOdPnTatZY5MYeaH/VG5sEwrQ7wXWfBoLIvkk8u7p5mGDrzoe/
5vQkj0xC3zv2syjyqcf7KKfUChEjuLFnJQvIj1akrF+tIbosmezVS82Jc77btzsR
Oeztrgn9S99nxeZwoICTv+upOgENGdl1zkm+SqIhfJu7d0YQkYEOT0QGCIkHXTUs
XN9F7fYfTPZfnkr33TuPm/mqv3NtVSiPX0YBeOeBOeivnQPLfPm+prXBv2gcZreL
KyvVi6GQ+EDCZQhxMi2d/M3FYiLCp+nC6s0K1OXFEdXe0wTMYxTy6VcpRqqzAVpn
slha4Qvw4s3QyK0SmNvQQc5Iv8HGSgtLv2CyGjdFB4Ar37Jft4LCQde2UjejeFoc
qAktdIJcL+4/BEQwX3eEivAR21zv//FQdP7AjufwUN4HgYzIXZ4izKTbuTdU00T8
1mhl/WcCR7ZQbXHDHLRqzga/HZYmji5AGXibkopzASLNKRAHlJujntsQ73ncCw4z
n4pAmNbZWRZBD3dKSmfrhWDTEEPP23A9N4IvhKCwZ/FHBXpwEpQa231UTa21XOXT
gS0e25030lwV/cUC3FcGu7Yap1ygp2jUwclfnEAzJDdE8sxAIyu2ztQ5qroYjoT6
IlA4x6OZjBOMu/gCfTUUsMZOBnpaf7/XSnsTaLpgAQ1n3h433k7kgcvdI50Vf7P1
5BacOv/1COFQsFoOlYmYOCNtx2fUu8HEuy/RZ6MUzj9J4D7D646HE+doqBDI1+02
pmYWBl0hUyvz1Itu7kdlSS3s+8Z2G3R3FFGCwlRS4IJo2nbO+QMUbFGF0Yn1HNVy
tmIpSAcuODNr3dsIPrWxDnso36dQxde7WYFJMsyR2GI8NvaTTLOD5Zn3lGXRAze1
1QIQIvQ7RNRnOCmjVyBMxLtC0KTSDlR12zMCOb7PI7GE4Uhgpje679oZbIlwa8/Q
We/FRQViCuWq9Lxn4bd5RO/hmQgEq4OqcI+CMPs9rDKIEMEdtJgtbT4RH8LR1JIB
Y7fQ57i/7nEpAs/53v2g1N6LBaCn29Evb1z8W3FeO41dxuCIYwHjLyhB8qYxcEMv
XFuwAVaTbwjPzMGgU55BHZwhyZamHeFua0bT2KpLUi6/IzTaMKKAwggLccDS6RAl
UCUoU6KBC9jhosdvUWHy2MAAkPlw3CapnFj19V//Lr6l4Q9nsQJAJafyQ9bkXohL
HduipjnCAUoZWpDji903Tt7v0qG96gGLOrHE/ReEGaMRX9KWqPzi4KTl0ROiiOe1
I5oFIR3l6bDQW2hWXSRHcmuOCyO9GUp5hfPtbB9uwueCwtE/JqLEfsiNCxohTdyC
ElIsJJIqMrvR1CcOZVZxiTat5W+0JP4sS9KNwxJK1SnOZN9guQPjeCfEWDQg0fNG
sSuBepXbAr3IdZKZEFi/9V8glQiGEyqTw5woIQRiX5RvH0X57UnE8t920UvK+xSz
jegzzmsTJ/2vjXJF88pa17Gv4/I+BjIFAwD632Y20D95pL2/e8uUgSrkoTdKw9h9
kVA3th9tdxncnM1S3SZ8BwEcpiZic+v//yjiOY8RbwBMv4jD/jO5k7HJqNC8x0Rj
HLX+p0FsjJ8GxM7yQZPB2IrN1kgVFhJOHM2tsRfZlbjX69PuYglmPIbqX/KQFdox
yVszI5ryDRdXyMfyWqXqG67uAUbQvHMIzesvYjdAulmApFNjtnBytb5oQIG7b2oe
f4ypLigbdqGDd5cleKCSUOGAReNXIRVj+UzVG0z9jUMaY34htWiLZyNbBOf480FA
wFpveKBfWeDmn1Naq8PB5I4cNqqZSSIf8cco4GaYu3J6leVNC/6/KO5x8UYthmEX
6q3brUT0BKFpvBlDsVK7NvyX3X3QhjX/yrWLo8+FrrcwbEhjqBEEiRf/IbJ4aqCB
Sv6oCZFskcqEnNqm3vubP98ZSTXazCMk+jXqWzL0OxM9tUFmQa7umeYy553v8Tjw
/MwObZ9gob3buloxbTLpeSzkCC4cXzokyfBHR2UQfs82BnWPBydO1alu9fTI3LxJ
ZnSQAyrkzYyGnLI+/dAkJenWi/6DVdI/bGTYDqXlOv0cqqnS7sR8s6mXhDfCtksU
+oMUVMDBstMDiMBSiL8y0TkBajVcy6xHUtOm/D1jYXqBo1tsXUCT+NC7JPNmgCmp
KkZsf9+tvH/SksvYgHxsCxM5/DrVLiN0wAN1c07j0XaCthYTCr/MFCaiecOa8yug
CAvqi4hap3Z6lxzcAodqRkxVpgZcF078cdksdPM5jyFvV1SGEVWaT2js+nP/HhKk
+L9gaju9NKm1teHJewLLGQK0TCwTYTV9A+8EwjufQUewy20rm1YVuGuGYJvn+oIn
ZgOpD0yPYq+DLTJWWoVgFvapPho6LANDiuo3ESLVoVF2a0HaEphH4u61V1ECzI40
i9ttVdp8Z3stLRcUrFS7us3zvliTsT9OxXY+mKuzrCbL3DL0LvWSLeP0VhzWVa1W
Ifiym7WtXi4x0+rG9qmmcrVQuhdIBwsF/J6QxE6ns4zxc3dMiWZHzCedJKHxFjw0
6+ScZMZo79M/seH0RWELIaMSnuWYth4hwb2Q1Dm2GDFgC5hx2OzSFBG9PKBV79Ks
gjMXAB1LIQxSR30+7uAh3xIIAaohP381gQw1RCqbXWzvc9LwzhlkzHcTstJCRv/3
n96YpK1+utV/xWkJIDu9OG7zVSNgf+qyaTDECdLwuln21tzBqq6rG4GJ4YkiGk7f
DexqmXnKdOzOzemVUhT7ivBwg2ZWyAQRJ8iZrwPzbHYHBps5TDWqWTjXEl1Ayhqc
pIcCHA9iQwkYjF687a2YBoEHNR3hDBC2bRXC8yFJuYGzphaSuIUO2LSAlpFQAx8L
cXCYPXcYhcpfqeS1zfAxHZVE2CYrT97RKyz9jT/YCY8kiKoPYIl58TiWUsZZifyw
Y5nHZBNy4piV5IUloHGI9mcn2EJ1oko76CREGfOqG15fSkSoyYo+O5qn8YtzX6uQ
jxTIA3/4QZ9nj+f9AICWz3Ozel2+f5w95+yzUW1Uq3aILseH+FknIwXQThCZrVBm
2Yilzetr3/Qt5xBWhEuYRI57YyXqtVgjmRxQ+gtKzbyaP9tY5PKM1pJNhtK3OZLk
eO3X6AXe75QoPj4xJ7mfneBn9Ep7ArTi8ILnyBHYhabrUGNKEkoNzkQ7Th3mGy9S
SKitQJJELIZoX4rmk8oKeyyxEnRQ4jbz4MRIg6MsJQ9fdC6Ggg1TeXJpIMYNRhf/
U8X0ZzRdck75Psx0gKw9ueFtoGFArUaKZ4vdk2GEoUdHnvM2mFVXyuDL9bHv8WMW
3KLXkPXNA5woIjSNyjsmtgF9xmeam3UdcgaICJpKFe1OHZSGAnVUxYsm/7Y8xYK5
hyGVg3ImM7S/Uf9mNbV75MyAo2OZNj5QpJUDivBMy/ZRJ4Q1rozSNa6sIzv1v0Sq
OiP9K+m0z+WkeTCbDsjRz+jLgIktiAO840Gc1VVDXdNTrPHeaEIzwYed/C+0kL8I
lZE8MbYZ3LIEmxHjxlmrphZQfF9iXnn/ckMw8kZ9gsEp3E/L3TuKPKOrY1nF4NPf
4tAl2ES43gTIMHzaVXF1TKwRuE7HaTh/viKEVQJMh3R5SzH+QaOJIcGgVv8IzGCc
jOEOsC5tLNX3bhf98CEJyobigKsmceaQ61kdHab40jaDxEfHExHZEsTschjLPgFC
9xmJ/M1cRru0Ec1azkX5bKmmJKIb4IFEVRd8ZMQPNRrw+9AU9fe+JJANseA2WNFE
OeZ00jx7TwLAWQH0KPAopJsRuRLBTghgtHQm3igedvWqvu32CvfxJ1l1nQs0r9KG
zVVhIkCLw3CCXZvBQc68j0LK70aqbKFc2t/K3J8LdmF+nNaalY5rtp/rShLkEPsc
6By1YoziPm9RtVeDiWopJbNlTHZTfMKsyQfD6hwAdWMvoI0Q4bYrW7tU/81DWx1x
yGZWrH9S0AR6MjrQcYL4mirrPCCCVnsH2jx7bUrHrIodCO20Vs4vAXVYyLg+nfn4
2Pz1nsadpCFwHBuaivAmCvW2U/D4kFR71O6s0dbhl7bSQnNSpPc9d6wV3uAg6WJQ
yBht3SQrsHY/uoqJOIxEZwmqcFlKf6V1xetj/oB0Jzyxb3od9Lx9GUgwtJ5gRY/q
Rh5iSpbm+sH/FrbFlHmuyTRjg8K3qf6zD+Uc8fdM2ZNeo812FTd44R9XBsH0OsBn
IwqKSYIFrf7xqnEBR8cqIGn7/2r6GNRPOkrS1V2qOMfh0Q1MHqiBWKf+zCLBUa5A
Rst4UUPkAYgmsN4xiqrWdXfrirs/NHqXOP+ZctSznWmQU+qU+Z8lUNUd7XfevZ0m
5AtN9GVuXVafu4YxQakxV/xzAJyrfPSFel7F8N9pHpDAxAtJyNA2VcTxcHHDdUFZ
SQ00YqMJy5KDUrRDEKOk3m6lFKluR8Ho0QZlNt4EVMhf1tD9N5UHH1AVxMXXRroa
7Vk3lTCt5l6e33kBXjioWXpjfPvXpJNpSgmf6Z0xWphjr/KeO50D7cnRDW8t/zE6
4HLDC0pjXQVR2vSB9Eq7M8cYSw3oRgSBwgM2La+NRtOj5xod5u0O/O/s4A9vD6pW
KiQm+cGHggeDwIKUzCJ5zeIyCUIECa2ky0fKySsdP5J0IE9yTIizPM/0ELeDClTq
FRZgVCoOytTdRCcVXDsZQ1VV3eRa5gQQmj1My2NP+P5E7K+gtI8Pr5u72avn4cE9
wicSh/NyycEvOthX2+bMXnRQt5C587+8qVKcld4DKcke9W+//uMSrAIyAjmiCwwn
DxQMjSEWsjPVTpKXgtsIiQ/wlDxP662mqGTaFUvdMOBE4dyZJg8U5itveWuxInmC
zoevAcGsSyVYOu8ksBqzV5QO2LsP1HVbklqObl+Mu9HrgRSsPpdoAZvHXEbog45b
QzTzsqIIZYWZh4D6fXZKvXNEtr9rvgXKZnWV2B6ssOrgKMucj9k/ljSsHe4lgwAp
p5lcWidtZ93xj0TMkUL2goatmQ5flR2/QWavz8ryb2lFdBN/0YlFCcywtf3DXlnC
PSb64itM58BdntlR/B6N2p4ubkn86kh1U3Ns/N4Jp2u7UfMMtgOROOGxcCC4hh2k
2hAoW96jr74C02hQjfNahbM6/0u1NQKTLYFVLdF8bEC/TKsJ/g8r0AES+X6B+8IZ
oOik02wSFXnpQ3BjF9qw11koiIoOURi/4q84xeMI/oqIFh01DLn7REdWc9biq36D
Y2bXVcmMfl5HXYIRuUTR/0S3OUi+SK57LjqrnnipK+0axEtUEgnukk3pMdTcluF0
1zlhoYPOsqHDYFd+joFYjg6nZBRTMdgIUSdAIL8UJIhlnIue8IRVjLLSbofPV8Ik
BN9ysvpoZMog1ngLh20g0108mIbApzh7N1r1Hv3mcTQgMB2o4yfwwoCG6g0+38it
tt2yNHf12UkRQSlIlUPRI2QYSt17h0Y03NM8dgfAd91jWDfb865tcd7AOolUNoGj
XlYIA1NWAjZkmNO7AlnR5AqGSFfkr3xiqWalJ2VSSSbQ9idIMuunqwOCjg9RodJ9
22c0o/hdRDlW0/opvfDLt16Y1h7+UA4LSWgAMAOddO+BnLOnd4cq64XcFfIJd7h6
VFjpQorszMyncKuQj8X0xZ6rraPtXBXjNUImZSVhh2sVcLD9kmFBdF2A8LTCb5QA
5NfcSQf6jAiTKLU5xwL8GUBbk50PhltrnNqO9NT69vZ6+OQTcQ6tRxwLWEpNWJEb
FedFsdHgbaoSwwU4mESX8t4OpVvnt3aNOKQW2RMRWOjswG16CBE4dcWB7NgL/sXn
LGVPHUPAGUhsvKTsEwCVDJkd7TugtEkfZ/8jgLI+2s6kgPm9+3YHLNNmOlbN/kpZ
ST6OHvqDfQ2RKgzs7NwKiL2itWgXEUt0sCQrXHNGsoAJaT/gE722nvAwTr7XYjun
mGs2DFw/3qdJA8GaQKykuBro/fWghoMNuyT1AZjNa68qQnvxrxoexgOyqBsQdu/O
y92Ve0pG6nqrxShhRzR2pxsfGayI02J1s+fRYPiPcmxjFTj8zsP46llYPTfv8FV8
AEwFge/eOQTMJYz7wtg5uLLhz/evvvoR3z7DCGy1dmWf6tGWYI8BaW8uHyqnG/1z
FjKdE2iHJuEmjaxSkpYDZ3bAPP/vrG2Ek/E0FVsiGkThewuD4SLbZet/25QmrSW+
uuAbPbko+Xit2hb3vY91R3BO6KTjbcJgt7EOYlGXO91Dh3IBs51n8QssNRmkTtsH
KeKyMEKXFJjTR0yt7K7c6VTFvoxApNauhlVOa+0lozVgav5TZn4M4FLCT7dnrCaZ
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
SCXii9iMyLI7vi7Mfoq5vVAxBpJV20LnJkaW4XP/yPMccN8c8aDDSsTMNkDHwkxf
bSA9ZDO2FyjjMUmhtolnnWsVJ2QbSH8NqJ0TSw7E2bS/DJZli2MvF9+stQuUGNvI
cz3ZcE7nqrJexsA3iGu4XzBwYxHaT3jKi7qzBAw/rHc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9293      )
8sSXj3+LTKpiZ+y34jMHEQaF3bn3guhYADh8nKC9JXs2KUiR1abR0+CQAE22r4GN
VPHT3Tuki53CGYLnJFEXL7WkFT3hkfiJl/UlQYvLQbRfWKHGmnHmLldg/NHKW6Nn
smS7Qk0XmvIhibvyDFQUJhjon+VXOYZfw5odYjD7g3YuWBa7UjZ2+kwn/99Mf16u
nPdABhZ1QUOkvFVu2gs3INUGCLToGAGPq5L1l3/ajWo7NXwO8OrUEmS9lmPoRAmt
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KGCvy/aZFoVlzCLo9UKvM4pFfJbeyyE0Mav+XwAIu4iDCm7siSwDxiw2389L/XPt
yO2WIpWwANFm8Cc1VarDoeVE2sThqXL8m5Jn5WpHZCSnBxksoQ6ATYJWZbFITAVm
dpULygu+4ZF41UEtrwxabEkcFClh9aSqZyEYbJ9PLqM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 18945     )
Hw6QDCrk6fq070rPVB/KHUCaU4RTwXQp7QF4cOrh2c21eDGzDVPt0OIo3mXlUOGM
lC0q8RG9l4nQhGteY8HMkxdRdlgSM85frPSszIkR502wV/4Aa8n2r0RhUevTq8JO
nsjIzFOFj86+UEak4gX4geufV7gUCjipZQqEhXr4nTCIfcJvVuCWE5zkIAOvDSIJ
52fVu8uTJIG+71tHKS/a7d2NIcs5hdk57Rri/t0NBrdldv0tL3hPFEvSZOG88Pkw
32WPcTYsKw8L6je84shZOuviMRwx5TWdzNsS6uvCS/eQCDVqvOs/m7tCFW6DpchE
G7Dlx+gkRTzzaNewOerCoTiie7mJq5VaX846wHc6NT68Q7E+7fOxwVu+a8wSg+EL
NSVHktqh7oZAl1MoshMUJLMXcTRIUuhinaxE/Ly4Qmm/gKeuTf2PyMACRwwoIHH6
xgzknwRJl6MPwlrQcwoq1zI104/tpa3j45t/cv1YwcT8R0O4YWFayUVi/LBpJgXz
tHLXttEJKwEq+A8OeeNpFg9avpIskrfjZlmT5H0SSyoIAtlpUAC+OHr+FzEAWe4s
hlm5QuWF+B2lylAQyPRtA5fSH5Sc3tYeBiVEIqUnoJ9AZsqPjDjNf91TM32Hc0mU
SNUcf9oeNzyclPpqgxlZF5OQL3tglvJ6Gju/OczT2HmiTWPKFR81JIf0oD43UOPc
sGcW9/g0ITZwrCH1W5E4UBXMGdZuYLT651OdOZDz3ZpPXVBKDO0YyfQHV7r02Lch
4KSkRIKFXmwH49bJs+n3YQSMLguCz8ffPrXWc/XNRpSbjO9QsyJ5uuTiyGmBOkGb
8eI8UUu0Uj/Gu8U/lAQ3mfJqrj5vso+9RI2MIM/ZVtLuc60JBJb4jLlnOza1FL/f
Wwm0kzzz/eMRbynm+yT8fZQRTPOHGfZugVPTQPP3X7BOn8wNxFXhvaeDluqrYt8+
A2fOyvHP259HmbsGEQZnYey8Zxv8WXg+k8eBMmLJHx8qePWPB3SgynLfwaV0nv2o
juMrQoMolhvZybBQRXOq9SNnqES0exact5ZK8LzhMBA1nPiYxjm1cHA/2L6gfJbL
wrxFQgZ6zfR5hEqVtBwef6AH0pcvKQY4Eg4MhLmOD386b1I8oEdJ7fOs34SQVMiZ
2LWmqAQaG0y2ty52+7h1qeYGE1OX+TjznIScSg0GznHcE8qQglocLf6RSl80rOzq
LZxuRUL5JUNBffsZjLN2lao+IWPXjhfibzredlPW0ONDLmGLitYBzWZkRIectKL2
isyzSAzv9go8Clwvrx1biedH1Wf9yK5pGN/Mvcu6abgyrrbeUIKwPjGlTpbeZF2k
26GT70lls2HyIYn3FE4DDqP9TvaPA71khGVWrE0sZevk/djSGrvCfUc+Bg76Sp1x
I5Nvj8gwwVr2Y/ht0YoUQzZorDAtNY6H03LRCTv+WWUoYt7AQq2pSBguAbDwzFAr
M3FrI0n/hW5lF60kdEI1Z3TkBSRsbm6oltNw2+hz5YDs4L/YIixBQ11U6+AwaOfK
LsCen3NVbJfVwerC8k8LLqJ9Lwae44xso4Lrp4T2KAzUX1IabaNhGBbYrStpfB8B
NqMfgGgooBvAfPkkKa56xeIO/idMXjnwS9GC+xvV7AqaK/A3nmJGeIynHQrFNBDh
B6p12SNtxvECCcxYb2yu6as9ARTHddWYhQHo3+cIZK3XE+bG8yHZIwjhAgcGyzje
4tQLMUszDK3dWhYezdKvJwH9ycgTkHAuOWrqCx4fzq059yXP0d141M64FM5aUjUu
Ll79G/QJ1ZYoma/Fjrn3amqP9LAvLGaCYhNEgMSgVkKJuTU0Z+Pg6EoOEGo9eS4F
3+1Fs7r6WXgNkOyU5U85/kBv9VxQ37dsbBqvuWq3eO0qRSuP4dy5u/1dYiWtCgtL
GpLvfW0D6PbfyLH1ldOBv92Xo0yMUuavWXev+kq26lKoCuTNYpgEi49T47FmgVbR
uVuW5rsj3Eleh0XYtT9cmbtLRRzHWe0v5jdXrja7i3F/g3E4ETbleVUzoxVBo5tr
qaJ02RwQfceX9OcqD4THoKDxq5qLCUi3Uc5vRS13TlIuMXttSMpExpdSR7aYbPnX
oZ1AJxCTZ3aCCJkcZVqJKyBBfS2QWorAN4DWEi2DDURH3VvcALML+iMK9FHypZw1
QpwmcP8i4+TPRnAph6AWf8xx/CDxddDszmhqg4cvRcKJPBr8wS1F0OCgsIM7/0jg
vQ4+VtaHmXjoiS9zzWMVxmcKH5HvQyFWwFLWr5nfCs6jvxL57w3mf1SByEgkw9T5
eToBpakhGN1B42Lyo7pHdBuwhtslbmjYH6btHU2tMBin1X8Bn2FMdSr/h2YkmfUU
iQLG3UMdbuegwJxfs4uz7Ixsf+Q1D9Yk/9rOkfyd7RWsPpP/Lcl2dHkdsCLTds/h
qIhX4beU1OE/e+qzp3at6Mbfaru4zrLRS6VxHs4DChUONr7XNDzMvPqlFzGx60aa
P2LIkG2vG/ENBpsO6TAMZiZWfedV+bxS4Jz9WoE8PpKQLIjK7xtwkJer42tc9aB0
PkOh+mujBZsEiwtEVehDfx+m5YHqB9nkbfqbgIgxYFeFU598asfg83TUjGWQOH+k
bajQlduiQqhCMRjiSwkomLKs49Rv8yfqaimS2F06g56ZyTHZm2dBRHJ5UkKl6lhi
2Q3hjVOOuD5zVNmd/acJgZ6IBPRoTvNwjAroAQjI2zviluA3Hj7oiMORMWrnoGzA
0niM54FtLxg7DBpH9DBxEYaaXd/mi1gM2JxUFyk30aUrQ0+0dX6EtnO/gsUY3b4O
h6xVxcakLcGOIcrPg6yvHQ3JtRvUhuRk/rUJCRF5PF71ahfg9qVIhuqZHVyYcwdK
N8xZqOts8KJmOlPNTvEzp1uXkf2CCl2NkrH0d2Yo242oUEs8wnHy2GJPyc3rCqhz
xaC3QkNmavjoEEifHkwuWBTDMklCUYzzO7YNdLy4TwGf6+8Xgal9/Drf0EPnoBw4
ISMlqBNHvaiil6R29Pz7j2NGUbfcPdSVn29t8dw7+7ShdujeJxUM8O0rXewr4Qgx
2P+3OwEK/1ll+SOv+2VPl6aDOFeC77MO41e6N+m24OIi8S2JXjVtMqZ9Nnl6gxp+
zqBirMa22ECCU0a7AnYDnKL5Q1LfEe6JOc2dA+dGkaqnHzgR38ts909NZTAsMu0E
vZDDp7Tvds0bOCHr2qJfnAEdTbuLnYdrcRaVj9l+CdSdHs3CC+o9VUoPQ815kFGC
8QDrLLb0yg11HEA7FXd7JJeilZLpEjT6OHvM/Zdvre2d+w/3q/WAkgbE2z8i/9sp
lOUva4hN4Ocy+CzThTHMvzYd4/YWJf/1Q5OPfvjMSl4xN63xTl4QQ3aiZnG2Ux/L
+++C0pEvNQTPcYz1m6Vi8YnDymvNmzekmrLN8CBDvHgRhB7I9QWzC8NSBDyRN28x
KJkef/uIAwzKuzffYx3g8TuCUsK5Nhk8eCEWYira+u1Pqdeh3QOz4WoeIK1XuGF2
+KjWS4De0fzx+K1t9ERfxsUfokKXcGruFJkQ/+U0k6IFkfw+bUfgeGMy+ov0/6jT
YwkT/vJosCAs2PVaf6+a2s40RKgOdOQGTPzf1qkigTqSk0UC905urLZg5FeN/AWZ
vBdubrnvjGCE14nWV0A2+V+wgJanT0DdQsdSWpGSunD6qvOibIQ8JfHbEp4XNmuu
CN140W3/Z5OT/pXYz9TGSX/v+jdZxwgC6PQwcOxyiwYDncrKYu9eCCcAut0m8z3x
A2g0xYVi2Bl/yZFAbF764aqvT6zEgCisEpoQ7+r0ZwmceiQvEHvZw2kFQKiGcSys
JGzVQYz7lRD0gzO4tTsj5hxCdTueiUdyUsX+xbjLk+vA0d9Yja9k+aXArYS9ROTS
2iGZtRA4YdmpKsn0q5rIZYT1fHINHKb9p7M2S8G42bSb4K9Z/CSeGdWb4Fz5iapq
ulK4tFhWgzOfpaGU+waWPRAfg419yMeKZPx2KD26twMwLbIK0Tdc9t1kx3pbaeol
ewHcoQ0WwQxJJDH3nqaOFxt/VB645MDMh14ii2M+Dhnl8aSfoQgOMmmeACaSvqjO
8ESgoM9EKr0m/k/SJ/MvqCfk1UTaSXV+Es2ix+EnCixUJ/0TacuNS+1bsLw01pwa
SK4B5WMIF83ENh6kqHFDxCcxuj4klKo4TQkbmaIidQRqqYdwcJHQVj8/iWgolP5s
ap07u/n9bL69kheok7zah6LDmA5R2kWY1N0CKMgEV88X5wc/k5bguYC/N4GKiIck
iimjjz9BfbKO/YM0QwOlidtahF61FQBSJhttB9C/qqJtk/7YWaFamWbtXDEXJR4L
Txet0+s+jjd3KcWWdTa8jWHp0TemEmrGYD7GpbEI+FUYEv/ilkjffWZJ4mw4LbE2
ZYlof3xT8h1fSa27GFZQQV4aLTT81UUQbKdFgmWtmROB9lRbI55weFOxj2lpMRXq
mcNSo3YXfubcLUixlTvWfnoewyiZPQ5zLprAlNCgW0z4o06fQno2TlQsCMLUiDrg
LxZxL3lhOA1fKQIW5olCcS3/9tP1QepLr7D7It6zWSOHWMQ6mCIsmtT8ZMi39oCe
8XTHXYon6hPInDGXBgSw0yR3VG5c/0XCZzrGMdhB2QedxnY33yjoRFH00sZOjfYF
bpAPE6nHnHBKFkkMKalCUzQF+u5a1NwP8QkWqU5RbizzYCDXLRpUzYwSduaLDE46
X7HL+HaMrBSQpBr2JMYmeA/Y6sHveofM4B/G9G54P9uW3R+z99JGbvQglIs+o3aV
EWjel6W7KJPYNUZIVdQXi3ts3QCnbJFa9v889IdmNrORFrSSFTQ5ih1nvOo0ol7M
RvxEEmxjDDSjjFnvVb10lS5f2Nl/8SGzC0MaO2KSdKdO3ZglfXlN0lHKm/zRSyn5
H7BYvTMsnDn2ZvwKRymlSRAgd8sZcNYr3kJLZK9ltdSNjri061U/jbLbvHtw1ViO
ciXl1eo0xQGH7WOLv6es2EH3ZbmBMBTVrr5WNz6DS+g3l3NvcF9rEczIPXKyTksd
YTR8aMRGBX2Dqkws+0FKbiSCYRAFQJKqywyBQ7+4FVuDekpRa/JA2cj/RsgnTSY2
jPjRyIoUxLPpbwOwK03CbgTSPvgqHsR1jjtlGt4YIZ/Wzver5OcMFQSDmiZQWhQc
SyiXj29I0akdIawazU20gHXG23judRkV1jIXx4F6ZC7CD2JU2kLtmjDO6XPyJ2ZS
3SjVOJycYjoCrO00dzQX2UjbwDxpExNuuZwhvq0lnEod87V9a0WNUTkpRSvJaCqR
lSq9aRSE2T3F4JbA8U8NCoaGuuKUbEM2N0IMaDNfE/vehiLPLAQxsnQytoKuh5/3
t/TML5dlR0wGhSELpW21e9ZNJ3FNG2GUxiNPSy+BefdwbS7Oia2lGpuBQ8L8t8ve
2MoZ3DvfnuV5JhFLONbF2sFV0cAqZ9RvQ4nTjql4qfL9aHbhGpP7sQoWvPJRkHnR
YAP+bIIEHSdH5JDouXKZUHRwqoQMBCrqQskmKUd+9HJ44hWUxfdrrA4XN9lJBZF0
aPzRJnI3z2rgvbsOdfXYr6IZ0Ar96yzN4dP5LfXHMaCKZ33hQk8dEtYeRWIaDD/l
Q40EXWZ7dTgckE+r41yo73pY2F/6wybx7VLj6FpefvvytlSb473j0Mm/LKUkEOcZ
Koq3WbmdOPrHv+Nq34hZzYlHgNcL3xuSlXlcrVXsjEMwVQVcLl9XsChiXiTcM4Ub
7Q/wQvEk7OumygzlAbRwk3gPhQxSIY0uAmE4NagdiB++nEKHdDZ+Wt/fNmy+/n1v
Vb1yMxRisnpYO3w5Bp2xQ3knWEXGAhNBK+zZvy60wIdbz3ctd3ADDuhRxL5npeC/
64VXP/xBRBwwvy+QW15iwtNawwLj+h+jsP5q9yexSFOLirVyEACMiP1s4UIpZBPO
NDU/B21+28sG4sapIT2J7Tm87yRuNVldRlsUHnKPF6yu92rpJbuD/Y4Zfj4jrD+Q
VZOzEldQLcY4VqwyNFALItp/ruZ4XKygBAEwswWoXuMSFc8DVPsknqtFi2G3Almz
c8R9OMrC01B4u4Y3X1ngxcv+SMxKDlx9NcTcJ03Y6PlPre7Q5t3dsuMCsHqqjbtX
VVIcwII43yo4T0uqKZG2kp9Nt9U0DStm1mf1mqKN+hbkzJEuFsYCyZFzBKobiMFz
p8QUBBTM7TlVTyLyIkeebxwjfFyOBOkPBoLMAANGH2IhUeUD8INsEzsg92fgj+o3
87m4SWr7H3DW32XcNcG+5fHMVAVILF3Y24Ko/wv1Bs9nmegp94aUx9EaRPQCUGsh
qsEMZh2cvYucFow98W1EQ3sQB/NAhgWBWd2a61axolwRBc+qpc1D9gEHxNV0Nhqq
y05fsdxurH+rzflxDtZnqnFcHhwrJpyuEmVOXK07mo0yEYPyI8EpOXMulYH4O2aU
/pGfLMBzXmJBwF8vNR9quk3JVk3cMMzUcSwxT5+zZHhS+DB+nhoCuhpFIolKfhpo
5pgffoZFkbSt24VllR0pWX+bBfdR4/gDdgdTT5XLlLwWV9Enb7dwiby4RTqO4NYx
fA+u/5GgAv52E/x2h3dMqCD6LQHo8EItVJkjetkLQMCgo2hX9uMnTue4hYAIBcTN
FYBRgJkpWqeXUgUTcXCO40Kg2SR51H2aG1gtr5hIZsJ45ihnRYQwj33m1exnhwci
4AyPHyaHGy4vTBPNquSq0UjX/0p+YiAw0XlQf8RVO+OjbIFFf7Ggx419x13oXqQo
5hhqJHYXmI2mWN4aSrT2gMYZyA5Z6/26xmJb/m/XhJbHLUp7/7NCY73qX+Y3YEbU
rXZoPCHchqMY6Vt3Xp21MGLSjCSQ5pqBkkgwgetfAN9oKliB9ncJiT4Kz8EOIswQ
MC0KLEevcLlAsdY3lcGGHgWxF0+OTeFw9zsK1sHZ5DHLLZQ6hBt75AsQfE01Dmdt
kLCA5/p4cFyoKP30a/p7RoljegU8njVhg68bfuzqcc9Cq3dKHExpaDaXXKaSU/0E
RsZkNKefMlHN0QcuXskfoJC/9RgVwpt+z8wlRuTv7oE3MDFp4LvTfTDc7wDZg6y2
oEl0AybORjTDUV5lclITvnmWlHrfDZKYa5jwMUJQDecpaSwiTC63DXavgcL5EINz
Vs6rywaqHiJSRhQBw2i+cOybqXJdleF/fhF/fftgjJy5OkefH2BIh9NTHgkzfo5U
pQsrXTUiWK50/WD9/PRGJKj/7MGy+MfTA+VAWj8fyohIAAsL6dwJzpqoL2COg8tl
GXeFV6xR631t23EZCouspG7bgyN/n3HJAj7LWogukalOUSv0gM9K0SplvUPfAMAX
ATpAajjSyLMgYWKYL/oFbLw1P+jQSFrT6n3BsHwuoTVayv28NRgIVdFR70T2+L+3
QjQD22KkEedaPx/5wD4DrRcRA32WXvjswIiUR7TNC8eON96YbODQ1jRpIkjIEUSy
SVLqhri1V39cPF3QN4y5OAYM5BhKlzD07F8dP3eG4rpCOpk+k4ghyG2ZTQvtQlH3
6jDI2Ts6sXo8gn7B9rceESWlFvPCQnTHO/HsRbAFN4c9aV6P9fbcM0PFWyf0kGzR
rnHMqb21/OILIiS5I7knVgZFTf+YWTHIVvUpDktLmN/N/+wlveO9vw8QyHGmxpva
00QmfGKDRjvIjy1tIjXH9yDNg019txos1CqxZrGY+EpFJF1fumouHrLBq8g4HlUZ
ybYKak584b7i1Lj1sSsbRbsvarU+MiLHvmZhFduIEtbkW89Rf3SYksr41Q85ljKB
bQVpo6f+dQfI+xw911ZqGEYMM89Cych5RHJ7xuiUsjfwjxSwzYvLF0ueIfanuO18
fv0ZNpV5AtFZDnRJDtN2gVHhM31CvW8C8sqKYY++2tebQnoMiy5rGQrgJfub/D3q
bXdOVwjSSNWDj1n8xqhJV/DuGH18QN7muYMIQB+mAoIMhV/znsQAhdozmePu9d6B
63wQLIzVaQ6xAGAkzqVq0t6xrSCwMZsjUKtMv+kq2JTQ1J4fNpmMRyOdFtHf67zK
P1Bk/j5f1uK576x0aATITKzqrmh/Z11fYiK5dsTAts3Veg1891fmhEctWRF+OZA1
ez54Mv4Mn24g9G5Vggzs1uqMN27dPJX1+ztShF4wGQHTsTWr0xzG/oQNH/ofyZ4B
JdO4GdaixCNWkyawZZC/W6u+S9BDXNTVvz3qMNJ7TLZLLsOqwPUbF9PVlkhP3MUw
5w505g1ruGHpilVGFbNUWJvLSHi5e7vXY4R9TnSOUwaoj5B2L4Lip9Vsbebocq6C
hU838Rl/7AO6eY575Hz7Vd3/h8JuYoPrBOKuXaLAaH+NLJU0j9Wy+3ftH8oQCV/U
JDzxXVYgCcKIJBmEl2FlcgU4WUDXfCwXS4JQljUdrUwKCy6mkQ341T41wkRew19M
txJiAi5ceU35T6OaDsPdkmU0MdhvhxYa0h4GbviU9ej6RsP7ZxzU32GO2VVJHRon
y83wWY+A/bzucYlSRc5zYfp301FzxO6nXibZdP1nQR++KfWHmJxgldKfKHUSQeVb
nXZJ0VDQ0rXiGdOwMqPcdbKh55OiyJ8pANo65+c+HJQfqvPjfGc1hSj7iWt3Ftjp
aSwrlgzTPdjIABUeFYVFSoNbggLribx5mX4VZtqEhbbu5jhEN673hlnH4IjoMlSL
HeQiJTCmKhJdpsJi9oeDmT9+EMUY4IWvTj2NsfT9nBo9nEn1P1LQCOIM0TQtyAwl
c7WgR+I5JJhXCSk5zl4T1VbUHiOpETt6v5/0chKCZSYmvzBEjkAUaPfat6gueeVV
1IYsXRtknNe51pyQlqUucpHwcC5Wq6RVb/iZcVC6Nxj73ko0Dej6ms+3PfDnXb17
y5/FBK+NAzVARdNp6venzXS3OPCP4caJY8BOPI88bA71CRgb/8JquelE7aKv+aU7
wKS1MQ2BdDCUbW5bqQeW648MMT+xuOh33HwVqPP6HE9E8yFgZ00EWqPLb+TG33lz
EqSXx09rm/Yo+7YDm1sBrfctzM/8fXP7j7y8aoO8xMnUlHiEur29yWWNtBAqrCyc
PECiUxCdReW5tOUd2ik2LuEdPmXd/7KgRe0VewxPkggKhUAGJEJd+BhRZXKPOcmo
tSc81nkJo5AOPIO+pYgQGriKsJFlHlRRqzKdx5JfAUywB1uwBgnHZSikHNH44euo
WwP98yQBazZ8Up/9gdg2k9D+GgvM40tGikN29Ylc8AGsBN7Z0cQCFC4HmP/f2xY2
8efJsmuBwYwN96jtRzXK7gw9nFtJYBD7H2k1ywdiVl6VEV6btSPnNQAHIePA2m7n
bGlsdrg7DCmU79sNA8RCQGESlhVCND5JYsCrgPbPiIVMpXruCLasM/Dh49Z4MGpN
Qfgm3EtRY8XAjI+krjPnTxzWOTAeCDuFSO3xOMwTa78vvTh/gwy7GZhQt2WtbfrS
9mQTPvEL+jxI3OlXM2rjwUbNCGlna2b6tg7rOsqcAVhmksuYnuZrXFtdNHgvrH8F
rvKnJmJWU+QhvPGi5nOrlzbgariX/zBKx1GH6GSYFbDL0IgOQWb/MbobuWM38dFq
qw+h3LDnWKJOTrQ2MlPgZi5VIXkpwiov8AryNscq6zgYXdCmGd3ogquGhZLjirPp
udpqqx2H6wCwui3Ol3fBhTS3MGPrKgkDdLpmLMzGuLZld4FRWYaqp+zwnGkbtz6O
cQbLVkObYSzxhbyeXw+3Ql/JrYcGTWZCWXYFENEeVB7d4x1ZLcWx0h1WiSMAsD1O
dgT19nC+pCyX2XG22plRLa9cwakwfN835O2d1tzvAMp7FdQrdVG52ywpuQ34GhVl
at8ZMFfL34anFYJu6LJIcVq37xaCYJStmCUoCfHyQhS/RJiC8oqRb5so+gvbTC71
QJosxoUZvL5ENk5/E7V/G/cTzds5XPXf3l+cXwwhUhK7hCbYJF8BPrEmVHLpkTkt
RGSZgmGI9McO6wAkvBv/DlQ/JN93cPhhHSLhkzp9miokVc9qLqWV35+tAjUpbQ2p
xZLP8BuAX7nR0qvwS2jj+wl+9WlOMfeQHE1B7vXT6+fe9EC3S9KBFCcB54i5kvPH
/eLZQw/6JY4Za6ZriGqjYjJK4B9F1wdM2/aCn0e83FPUHHawi06dikZ0msNBXAzH
BNrMGBECFO8sYctB8haMygeiUcbS6xBWAg2AkbjvmPz4O35HWcGc5xV5AuFvt1bb
+6YqBwk53PRSZiihMDRqgXEC6SQr7CxHQ8nybkLqGLiRKUr82tsdazkiTDp2dqGZ
ssXqXuLibFihWPCdjt5N8/WT1ZgResJAUw1iZnda+JuOZ7bLeaqlVGSpNwE1sX4F
taRVHC8XWkKkocmdiDP/TmANDPqbC9Kdz57IvTp411uIQ4+9wwzj1ksU0X9chVnR
j3y9C1U4mJKnGFYiK3hDo+Paxy3QTehBCMPhSfxs5x1ezRNsEtYvEzJqbIVVQp1J
Hk1YsSPTgDgAINPSZ7UWAp06voWbn5aJNtlKnWcXOd56AquDnSTsgNUx+y0hbXFI
xvCXmWUIEd+5pblxO2vSM3xzzz78Pbklfk+XZzbQjquEsHZoaVwgoK9eMShIJw8h
OJJjTB9a202paLc0sMLkaKR+tXb+YYYZNB/jF/S444QMy4gfrvbRA38tvKExfrgE
gk0cZZKyGpkudQj8epYoRvDYl2h1SvJLWI9y+IvWgNEC4SJdUde3Kl+cFJ5G+4m7
0KKp1+Tjel9NKenk1NcR5tKGhVC98kSrotDbgEu9x9zqTuMJ9XgYPNdxsYR6BFtC
hzIYYA9422WSpuY61vWOTg21+u7YAo1aycdB8fOQP6Db0vywWzTH3SMxt+irFAVE
xjyQkuHcHvWqovB8/wIPsEi+Sm07RSk/oqmtfw1xZtxJDRiw1f62+98EfuiKrxyH
i6rz1xLz4Ct4eMrU4HtnEi3cCeA5qRHvC6jgO/l2KD+FhVggWsYii8He3LD6L/oq
bPbPqTGx3ge0MtTSewz+TgMLcXev9ETaXKM7H1tQqz/sLZiDgAFz6IttvrPQPLx6
nT5oSb6nYrRefl3FVt7v1Fskadur0tw3tXBDaoww8+hwj4YHtk/PJcWTgqm0bUdl
e9dMSJ091EEYHSUskSQrEMLhsjfUAbvtCKIng2Py//hzF+I5zM3xIMOONiY9alyQ
YevfVXL30H1S8qj1bUtx4YYSFikhRwWkfDSviJbdECkzaCn6ElUFM3ml8QUnBddy
+gwPv5iOPt8dmF0YvHdDYOpVNL2C6fQHP++MvcUS5cSYAb3ywI8rKz9FlK4HMOid
6BPK949kBYa07aP8YASbU2IvD5tHU02Ek0GJ1sXNikGrKtRJdTsNXJduSQyKQkQl
BviRW66n7OIzBMcl9y2IR7G2dRx6KKmcdwBjXayMzO0BKOofAjY7+kqj23PCUM+a
Llde2lNOo9sJAlfov1D3fPhESOrkspLLW4AD7T8U0RKuPtGd5E1FtTQhlEU+nDZ7
B5e2Ij1rUjgd8KZ7MOKgO00vvMbK7mIATIHMM3pp0eIiK+ZfOnH5TuSVzJPPbjWr
DwURW9Pv/AbDkFnSuVwu7F2Wu0/zOupMCulsdDWrNBp2yoqcatW8jPvbjbg7zoEp
wN/lgysE3vO9Sz153vzNpeFUU16rAJodOyWyNAauMuVemBDbZEe/JmbFwx//JVRN
LD7McNERKOyAjKcK9Wth82LQINslANub3nc1/9Sb7XH5OsYfTLE2IzQkCUZ4KFeA
pogEZMX825jsAzkyX5bP4Ke2cWGHG7vso38nc3fZOj1alg36icgKUvo6TeOhr199
YRqsjSEPVzsGw6E4OondS/6U1HcHPO9lg7rNBXt21taY2YhlbrctuuEsWcnevIGQ
oePOCuPoIyFvCe18Kc9GeAxFKIKTNUdEKqkyFvK4Cp/Wdm7Kr1Uk8qkqVDWkbGTB
2ocTgCh1ykVLdtX2tt4PY6Ax//ywncOgB7k5EwPWU23qJgktzSw1r548EexaCEEF
qN4mbQlG/ex3HYasoUGSf0MQFdlp9nn2iIs6NlDlidhPJQF+3YYFcFy69jWud8Rp
F1mwy8viz/5Pcf43B7SMaFa5CYJa/uoXEKwVQioGZgCWDXXluOSWlXDkkK0MXogu
OQRW3wkDc3b5ms93jwXaNpSkRZFSwEG5Be2CDXrm0OxeKZJrqTLCMZcCaJGyG4qe
cpAbJ9Z0Y5tzphL/G9EYULsLSNRVKY41vG4dwB5Z8uOoYjHLdP/YIFGQwxlNYgIA
JZvxryVCjf1M5NIBw1P+UZjw5KP9yP+AVXIO45h0tnO0BZ/kZ1cNzgBJASYk0S1u
fLheKJmkfkRKmMO4KLzrFkkz4qsB6t5WbmBBfWX4rp7kFN/3P+/LINYuF9EqMDSR
OjcOldWx6clao0Cw7oY6mvVtURG5p0+hChDAx9a9aFdp3Y70ofaX24jS3+sxxveb
CyfspEfxuzI7g2soe4M3MfbkmkwLLbI8nW6zKlaLsJTqVVpOE8RtYBBoT31HdhmU
ZgxwJZsVov/AjjkfFwhFsc4JC623r3llPZ2DULwqYNO5WZ8BSF9aUPW2bgaue2Lm
4gQH15ZEtMdxVrsDMNgsqeUEfnkLEfCyh91QfX7ItoTAWGJGeRyHnIonnLse058t
5dF0scM+V8cKg26kAKhccSnDSfd1Y7eOAd+DixNGhVWZaYYV8GuOkYo2M6Vzz8ot
Zm7C/haoY8eyfjJPbRDp2lrG8Aaptr7hu3wDBzxOTQ2PUSc+1K4zv43TbVuaVz/i
JDBiE7ahwDkgdUsbR6rlDewpoVv63unDdD258xJPiAh1exGK31rQvTamVol2p2ga
FaGWEzcPKZ7P0jMqLK89ww==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DRZRop5J6NSqzpN/NrJL3SOZG9sP8JgpxMqH6m8dB9AMuIzpp36v1Gs5mRsX0SPD
wc8Tzi9pNllw0RDacijuiklVy5iYilvSNmDS7AnMDVgSCBbhjzIZiCgjvE7X6OVZ
CPWAHA77+1uyxMr+XbuHnyKXWMCNzlz1zunEockNmzo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 19116     )
YBG8U4PtUscz/Ujeexi6Gd4AyovVQIZ8KoyTvQzIgGcBbRhYDSLG/VFXwat2VxsU
3xmAJv4cryd5W8pccNghiQvlge9G0my/JgXIhMdkkzNBPb/ZY5Mx4kmkFlV20Urq
qN+ZrL3OGqghC1CAYiSG+3hP1l4ISrY1edompl2ctI5NsRguTPhn0WRQhvv6ZDO9
o6xwdiEs5UYnJw/DYPZ7T1pyWk8MSs5k7Ud2mabfGVw=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OF0xxPprGdMF40B/ojT481gzMgMd+RhnC4z+Mwayp8PlC71LqmcSyjadFRxAR18p
sOLCbw7kYJ9aR2rEl6EiYTdQCk/GHUUAKUpjUtZtjnVmLHPiIn9764bKsF34ynQD
6+CBxt61u76SZAk27xRSkX5/InuLXateZN5We/XC9w0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 125776    )
LZS5eHJkR9cvjqnJeQmzRzAksRsYBS2AEN/awtxHjyNkqRiC4o0rdLcLGglMOYAZ
KKW+Ry9+IteFJ7Lgnzq/Qxlcep9/4wIOhXpcj+5oyfcxuzyRvZ1VwbK9eTHEkdJx
lbr673j3v+leg6G8eiTtAz7xkmmK+VlXNi4NlLGr7TroCh1lIjAWq5RVGGEqkvgx
7Yf8OgG6fwdUuIe+XpfhWCrJzH4KNYFpYThy87cmpxW6IUD45S1qeugeiXPzQFTx
S6A8qtknd84cfNRjVdJ7APhdkkppn/Gmnd6qaljMJ1thEC/C2yz3dS/EChURsUWb
zTWbV/WxwSU6PckBSB5f+SZGoOpHMVRgVeSP2+U+DoXxsE+pLlH0hjptDj6t3myp
WP33ObyKU0EHAi6X2dAi08agZ3K3cNqj++4U53ixZPLn7WrX3SUOqnyAWxEhdun3
gscxE/e++sGKlBRtnsFftzuk6G/L1Ckpjbq85dInyAsA2LzlHgrxCXYDHbQPPjcx
WEOLH/DROzhpgYfupvIN17GRQsHrqhcet3r4iUThJQrr/dPVcsIELjMDQQYKW+jN
Yv37JgDaCqRlaDYhsLE5cq6xrfxMuC42s4LyBhV71jWeluZDxtyhm+rU2ltNrh+D
1fSGn4fZDYIILb1QdpBmZ7khhlG4LmUg+E2fSHBQOXsPbKoEJtmJSW1n5qHf1Kdj
Aa60rC2K+a8HA5TIlj5CYajrKvVDoZhqu3ULZQy1W5FuaHs5Cb8+Vz5BxqLynhzS
wvhu6mHr5raC5j0XGNMo2ppN3XaQ28btrfiEV56JObHSwLGmwgA5Es4vW1PXPSqY
ryD2GAaJsWD2RxBAxNPbfC+PXenK67BsepzvcG3lF0DXzstOcOWsAGSxtinwBZOs
AL82/QEm22V4qYnZUuLIncIhOSNQNGJwfUS9GR2fMavyiXBbDylR/uBTSz4aUItD
YDMPJ8/Zfse0VqBqD0jdwDYMbppKiObFKPkJnsboNjh1REcM8aL5OoVcgHusp3eV
MNbyUMf7MLLPAcc65KrX0Gy/7Hbk4KiqZjiibckm/PrzTfOpf987NPJwMxMEzpw8
aGIzGEyQDQBAFsuj7w7qF8UsUdu0Yd5Y2jIaKhc4RRyL9Tz0AsYeHlaNqNVvxZGl
8EZJz9AOCwMCQSz30KaSJkxwm6IYZ+Or+2igxjfSPCpXUd6Y/c0wYPC8ecU4q7oo
tdcjAAJkxcUE9zKbt1WjHGv3naQ1ZfEBuIFzrZH5guRSCzRlgwJTMiu1gJHc2Liu
KnS0TijS3R2eVEZu92+nvhN2HKXKQBQMH+8qEQSrftkN+LxEqIqy24QFA1zL0Bbt
3bfQqcy2kuGKHP8pyKSPsveDx6osRa5aXt3RiQSCv5i1C01d9Rpq71VLW3yRc4qY
fvCRQhb08CI0Ie1N12MqHd+ckZeeDZsUB44ZY7OkSRXyzTI/3mXmuHj/g6hfY3gj
/n47++XmwnWSX4yhE/qlKhc6nt7FQemmrlv5IEnvhCKjefNUdeNQ4M8+zkFNNQ2c
DbwwWTmDu/IwPFCbux26EmE1J839BqnsbupQ0e2kMCuU3fd0HWv0utDuTirE0onI
G34dOHwSSXK+UUSj5pfF/LAg0J5hCg4WMO/tseDmVpneU/HCcpAfVh23m6EJpX/O
PcZ6jjS+2criHhYWfrbcmq2zKVQ7LGOFO49FL+JgPSpQ97brLjSXuiQo8C73G4Dy
3+DekxlmoHeXmjts42ArtXIQ2TiXYQNp8eg04G/1GWoH6iSaxWyh0Q37qySOsv/F
SEaw4H0Vd5dS4NQHuKwX9bQ5nK8U96k9xuFPslSjxq83sjFSw+us2IA8STMB5lLY
E0pCgZ8AGEDb2lr75srIDFwrbDdIP2j1sJGdjrQNBgsMqTfM5oiH/Qql0OKOXjea
GMn9aGWwwDAwsbb1LO0GsFrbEYvAlt0DUkQNXX3ca9bf4iGmEf1aliEW5FQ/EMgX
PzS6NbGHmeH5EuL24OxleEPGz3k9LMtaHjeaPMJW08X9YFhFQO47V+ATMPIwYLTj
hvK+Ky0PY5B7PwTTuawDI55A6R2agnRxGwYbt4gSGKREOkkInSGt8jMNicu5l/dO
0qAjvAcG8qe/T3/V1MrgNxS1Ck06zFkTJlBrFig3vyITJi+tkOvT+Ay/gGqIpOK7
6D2R+QmPAkdLj9yN9vRrTk2Xe2MhpOi8FZCLd291QT77xO95sqkxU1vOlU4LhDhZ
jlo+4WuKCgmi8XR8o1ZPkhOUPRL0NlaebDM+NLm7O1lGH3j1mD9i7hlkBmDoeQGi
CScPspZucvgsXzegbKBVroXwq4j8dciassk3iStpYrbI4HTDIsjKkkiwgtKWnKjE
s3dz0rT1OrK4Q0WFDZLINCKu3vvYKUpLhx6BToB28x1vIU9v7BfagoiTBJ09RYLY
wWTqCl/pkzfWUPvLlMULK4u0sYkgDqenAvOHq8GpxVrTFUSAzSAzrrj/0base82w
p1T5EDgz4ZxiEpEdG2lNqJt4AyHvjz31WKNF6O2nd2Y4wT9t8BErbR6HSbFQ5NaZ
LZsq8DXTwxstZ1V5DVPMoovNi/njKZUO21quCrFtKqDChNqkMw3Rq94jvEXpuUTp
RSgN8QXaLznfD6zdyCFCFwsMl5fqpxZioYQrQdgmH3qrDNh2e4AsSJiHO22ZpqUm
v1jU6eZirrzjINwdgmHT/mv1yzT0z0hSrvvFxgQCv8uxe7E7mQ7hFHH+zzwb21/3
ZadTq9fRBxjsq+Mpxy/WPCNQV1MGEbctXASJMFsLSNJ8Zi41oI+Mm3ZSH6PcF053
7IvJD6J8tmMPZyYku5x7ZyvzP2gQSQffXQCiaGnM4bUhJOp7nCPTx/BmE6AzhrSW
xEv5+xIsxGyn1PeBKvoLKJAkYCHKGw7eHrsdH2nD4tClROLkNSi5Si87Wyyvgei6
Z4L9iOQ3N9y5EbHelCUKgyw0maJgG5r+xEvgtyG0/kD6bAt5suNAuOP1snCecKzZ
Caq7mQR68KhuqPang/1IBWx3ieKPbU2o2JL1ZpS3ckb9+jGuGlj3JKWyNfEDKpaO
vCYb1aDI8AVUk5mxVDD27JyTqwIBqA7UG1Z8VgvdGw/Cel4/KS4CNGTo4xoImgr1
fdADf/HKUp+rTPMqRnD7ay7gMnfn5Xglh4JckLYzqVOrEOo8gHCeFccrWU+cDOJl
ywZnU1GJUJAFQ8CAFZOYrwFNbKc9Gtd3b4NBehEkESGkNG9b8dvg0ULwDBNo2ocR
yAqAp6uoiPGmpAVFkH1OO0Ki+Sb+wHOVUqtnVUzSFD74rAzWE7yPN9Fq7V2lpxHv
4LAdXYxkrK/VxMBt32VbS2vL/vYAXaoVGX13EqT+nkd6fCl35pXHFixnXUF7zeSt
/URtZ5+XHBQXMES1aOzdZ2QFEWTccSEGuARiGGvSwjcfkEc7DVitfDTlhdtFcnJj
VFpmrvzw9rzwR43z17UJkvl9Y9gZMkI3CX7PvISf3sgkYnzI9dCvx2xQLjHVPRHs
K+9zTdkybm2T/YnOSdhb3TzjtiaELbDRlKaYgnfDO4Yl17UCFvWCf8Cj9nP5Ilco
pCS7L5Y4PCmPnuV1DE2AMi8zRcUg6Xl7DnonWaly3Bxz3smCjI/CfngsH1oiP707
I7oMHYHt0aCLjDnVjUA4pFtWJQkUJI7X6fRvcZ4T0C8QjQ4Q/cPrhTBoCFJ+XLtu
Cx9yuseRMy3d0vwt7BsQl/l1b2rLnDOvsveQ+wTcx0WxoABl9eDIq4grsfFxBsW3
WvFyVP1rzGmtO5Yuq7l8hVSRixj9Ak1nKE1CZs5YUxA+NcTZj1Is66eZWLGba79J
1e3qgcGTvav8TOXNqB2ZNqI/6Ccn5cJPcxalRQ02TR3lk1Yh4Y1ZsOgIUJ9b/ybb
MyXyCLxQhYXPY3IMBV0zNJ6MKW1/zne+LuXNQXFTv1teDla7Pb0xzXwSklogdXe7
llzg8ZIPzPc6Koedage/u0CIIxcRoOq4C1bXIMhZNKz2ltl/vRJPy8KRYN12JnYj
oq1ZAPcLsK1MUJg+29x7vDjo6nzbEj0XkhyG4pEblV1O49COcvgWfFLNGRu0/ZV4
8O4MEJgQ0WIFN2PZkOg7wWhh8v3a4tJAyw1cs7/+HZLvyDjnM7OJ/2Si+9/Xi1Fh
gfxULx/YOywOKdpxuedPkR+VBvdj+1udzBMSDMu7DcR4xKepbSqdN0aMlniGsaiv
+r57DHLJZ47roJFGiUqX5X5wCmd2Ir8d4N7Mr5ET2nRDdrNPWszkPiDn5teztRi9
peX9msz16wePWh7m8830tla6+46GeJIPHb3cx5gOMB3SOdAE21qcjKYpR6H3XpF5
c9rYaRiu8lcBEdNMGae4HA9+FTN53l9e0X1UCENJ9K1aSSdKbmg4heDLhZsF5SD7
jsi+hsPDB19heIueRw6dig7ISy10BDGd+gjhpkCneWzt8TM09fuHZ5sqhTVWNqp4
xAFWP0C9AvV3sqLNKI05YNntEHtR+PQx66i50Beb3GI3iH0jpOHBUm3IWMrzWjRO
CdPErPzRLZ7NpK02g+W5WyglTXpAKmzLR9G4+S3++Rmqf8IxkMA4hpBweZ1wjGih
QGSa5jXDz/oH4Mr9EQ4b6GYqZExKPFWxnyCvmCXiYYgrBhs7MMTF619BvSFr5kWI
5EWsc+uRMU3WfYxOTgO0rErST1M0oAFTEtvi99ZpfhiutDiOeD72dLBvQs9aLK2Y
mtS5hrFDU8t3pO0P22j9QICEhmi7VR1XFVjGyefVYrIa9C8vXMjKYTAT4dLux2VN
3wA9CYv41d9Vp2ai+lJVQz1ULk5P+nymjnk6xScx06jQ86w3OZPigb+JfhZ1mAmb
Pl8bMkiINVOP1Vw3LZ/+1b6mr+LvnkJarOpEqaulkeYccyv2YaFtkkJzYQp6T8ai
QJ85JEpWnVpwygOGketVHKHJ9K5HI4SZ9VNAOMJg9rbrbIpFh0NyZ/QhRoc9Jg9S
MPM3qNxvxXN779eptErJHfEZd84wUcJgvrzoDwnHYb0ZjBVxy2XJ6D4awF0GaYSN
gBKrWp3ZTlWCcl6m4y+zDmg+RclmxSwqm+Wa2+ClSCuAIls0q5JBEdlGOIAPxJ44
LDSR8nmULJpqBkYGC32urhcblgDqnbtgie+EYwLt/qc5pup98HqagBmpJEwFQUk6
967s/EAcUhXbuAVuonbgYCwlDZ2QCpPACATiK/5PDS9oznL+ni1ZYN/M6Ow15ozj
lwBMFRHYjwvbiN64liOTFGAZmmdxeBQycuLQ3deM3ay9IrCQ4xQpo77XAyjDRyEp
mPMVA6VUkxVZxmwtgIiOsEy/JTA2aCC1v11hKvLeZGW1KLST+vf1h5sgk1ujGDuB
YCvY/X3jdOBkNapWhIBPYmT2lWPwlyNa5kODfngel2eMxxqgwSqGqjdlJjsj5SHC
8bzYwWC7Limcj40jY5M6xe6hMSrspn9YHTu6W3+ceY2TwJoCeQYSREhBsHY5twiD
wQfz6I0ssoJEoA9C5IxPqSrflYDQpcCSVUFeHCGB4ZkjyoPpSWecBMQr5w0Po9lp
7u/VuWn0dVlQNaoQXVuA4/TGg/E+Qz/ylybRnha4vMcEotTp/JuJxV7mFKrz8LSz
A6lmdwht0bPUAAR9n4ZRj7aRxZHXBcGtANmRkaOe1DWcinwpYlRqDlr1wdFQZFoM
W3C7zD+4iAfQh/SMwYuYpoWhM11Km1TNPbKtQZ1SUvQ65+4edHkGb5XnsA/5SANv
m1Ss4qL0i67GHSe+dvUC2EtiXivdPXyZIwg0jx2omb/tXyKUpxHjWMtuXqVVfgm9
JIk2hjnvvEfo1BqP5TxcmRzP3DvS+Kjr3ifCxhGJsO0f4205kT/tcW+W3fvQy//p
PHGta2HDP9/ZrR+ptBITUwKc6zu9g4Kc1UFVEWgTbPJMwPwC9QtIjW9p6o+WDGaL
4LTOzztyN2Fxcn2Qpk3iTH6WpllCtvft0PgkIpu2marDKM4jmPSznEH1aJqoWqpx
cHkGEbmE92U4NC9HYtc1tm9U11u7aKK0r7OIbhZPkIGLbL1gpZklYbUUbDYiEOqY
iHp7geL73o7hAWUT6SDjwphgsHT9BQVbyoeoli1cbfcLI3yNgG7dT+L9RyUny5vh
BM/ZWGEE11KphuMO7Z7O9HnOKCiggf9AWE2gWLNJucNmnl3Y94n1vwceV9sMFHo0
WsSXcvn4dxyWHZG2en1W507oZYl6rVJAPqkzKTo9sMYFYSaj2GtbAVvwVJcFL7Q8
kS27sFmb492wyqInNViiRoK0N6ZZ3FuVSR7OKvLkW6eNRuGzJX0m+UeNnNS4dsGi
RxaQD1PrX2v+Iknvrb/wq2shsbpd0fxrcHLfF3xaxj68TmjYsgh5CKBGdgh+nBNc
o2asEjz6mrZpXOP35CZQ4grNavlvHBw+1QpR1a52MkpiSqlBGwHe2OafA8LN5iKQ
EQGzlzZadP4yuLl3jpVJ8txjGLXBY6e9Cd68Tmf5ecJ6Q+PoaBEtMhV4P07vxFPi
CH0HA92QAgENOZCZ4SKNXqV6nb/OMBXZkq+O+ysXM1W5sYjB2SVAHG6UPaoVfIWr
T+Dy4BQsr5cJOOQar1e2C7rXjIqrESgC+9RmXaXehawI/AKbuvhWM3gE2ohtMz0f
gKWoqwwSGda9ha+zTOIIMw3jnNaRtxfYx86+yxxgAzzL/7RcTT0xZwW4bk628RKf
VJ8R33fed9lsdnr+KIOkkFUtwNAHFc9Cv4yCT4zVZj6sMVurJCy63Tobbfr0AM1G
7dy1+lQhvd7lwoTcOJnrsViejs+VnSTWncA3yQchxWpNwOTzTrXSsimIsA7xeWET
v0uYtlE+9YpasVTtAq3Bs1Z5KJk8vyPwgaqManKu0F2KA6nkKu6NAYW7LRJCjKAy
EkDXq+XfpSAlAEo4JKgA47hbD2eaw294xAMmkal1ZQts6yzKu3u3L3WdBsiQaQ9c
ApWJzh5cAoCIMKhoe3UTE9L4tj2mmZKJsb17MFgY4OLZcHVPXeT29SFoyvMm9Qp4
QxuqYlwg/scequDK5JMf9ERC3xQgPjWPYsbsvtKWzhVeladXyY43bDpfkWystX+Y
PpIyUOohLi32tATQA+D4OSLiIeFjqOP9HoTh189prjQ6eerfQA6MuuVpFb0zD0mn
Z5Wc0C5FXdMUk9HEQItxvWa4Rk8gxSV2b7IwFrNLFZp8FkR9+NL+3HGzhAehqksj
0e1kUfR/EN6TzOdmWDza/9Y5YHSoNbXpqqmN0XxbjwgotdcfBM1kIBMPQDsY1Cau
j1jasBPZvmsnpYKVKISyJuWvgF55CNxXa0TabspPDpFz0zKW6ROZ//kQbvv0ABqL
Z8wpfqFrpLoqYe5qZ0UERHQhHx8Pn/dqLSnm4V6yNYYljLU2s9AAMdeAXJoiSHN+
5hZ1ljEBWXvnZ24tEm/Y5rHJVq0Vl/9EVtT+m5Ir/zaSj/cg9YlhM8NQqSv1fSvp
wV5ZD0/5xt9jd0xWKfE0++XCo4C2ZstHoKmvxTL7p5qo1jblVXfias3rRp6GFq6f
PKGgiAyiOtO69KhXL0NoIx4wJQx5YF5to4ME4xgbw+u4VeGVH5660eaX8OnIswPE
8kGMXWNycsgq1EBx5fm0zuUXt0WovfQCgmZcAQD3+anPIBs5XJcKHzEuwFgomZyM
w+pa7yS71QzPZeFhxl+ePnsDltB8L2eP6mA//d/0BPKE2DKtii5y/ZW6JdES+kcm
gSAL8I3TwnqCLjAZKGFcpLjvThAp68j93hLWIs8rtJiPd2129pETc9wUi/rSSh5S
IoqseRf68t+V8jh2p3Qvca0J+sOJtOc61wDePuGbiXesqJncWRyThGAFVo7iFJDg
kEXB+2MnBxre9/Q3V2xZNaRQ/EsTxy2aB6I+UwgZL2WMEt6waWXUqKhWvjtdW9Jq
Y1ja0hkmOi9LjeNFXTm5GCTY2gX3sosN31PC47tnBAFNOkm8ioVF4jgKuHTbeJE1
ditvUqbNmIoDa7GMiJg3xkNHYcK4xZOinsG0R3juzsOaMkdQf/3RD/WHZT5P4E+b
amp1gXFNKLTGh0drAYdBQL5w2dDHD/Ibh693oT1Y6Q/aNkTx8EK2NMbm1cPCWhHm
DffDVDA4FU/UcI0uDNBTtpAkeZ7BRp6vhJRpvyfQjV5DEkeI+MvEpqkd+zXri6Vw
TJAcVWS3ACbSJnTfKIpHyzgYk+iE8c8i5e4A9jCnEuMhJrYzwcZqJ3LYX0RHO4+m
AC6dcDHmAwfdG9SRDsskR/Iou3AGXR6P1ZN7Tz+aLcm/QKcH2RbQpAZJM9z2yikx
SI1rSq6rmULK80BRnhYbg6l1ybqRlQBwFPJPw0oLP1grFBVp9iJMo2vybwsMohTc
ruHMunrYHNsGz85RANE49vY2dIyOEzkAc4huNW4nIH7GnnpWpF7k9qKq2+HYyDoT
nq2LAW9mQDqjhVM0bGDnSShxAZSLIWXkjuXguV5uwsvpIw4Iyq63iyGrEhjNoT2d
oYQiKMCS5gYH7XpwKZcnlikunRmVhyzHH6x2eqm7R+1EQx2wPOIgsnx9wM+dQHWQ
FaKk1dz1lxA6SKHvg6SKsH6pEODjeWN9IuslFInTX3I+FFf5ARo7g/vgDZYXe/V1
2nRl5grhGEwG85pC7T0MWNRacSi5xtu0bbuQMEPn1+zmVPTiMCD739oGik9AEVBm
Z94BJbVh5VAEOPx0siBv7EizaXOLVEygV3UhUvEp34f+bRYQJupwattgnep/ibwr
IAaojn4/b5jH5itMPvKzIT2BsDzR9KZBrL37G+xO8d/avfVgPS6bT+O+UIs7JcK1
6gk+BWUwizDYmvKV5UBdvJ1UekBUtFy3SdG7nAO3U+5ruSkhaL8PSkOtDyYyegps
rt99H7/O2JRvzhcLPFQJ584EBomgkzQaSZZ1tSGQappNjJZxoXLqP2VFQgjy1FIQ
9U+hC5UpPjU86qvcjFBEzg9nxWx4t2eQw8z/IC7EdHsad/LFR7AGJbshKzDdOdMP
BcFw7m7tIhxHxw/Ak3ij863FoAO4uiqNBp69C2in4G+iQsdyguFlb+O87gm5S/4H
tUUB+9zIBGRyJmL550oEt6Hu/RhsYrOOTyGSYfd0iJ5P4KF0WDlJbUPavrHXjM1l
eV5EIQ1whdoN2h7zY3pSJqjC35AGfiyVkwQo8J7rx3uw7qTyRJXZPIQdd/ZZYtLh
jFNCnsX1dVfjptR4L6pP0Itavn8y+M7MyS6rMDYp6K41MEmr0aBBv9IL7MZ0sLHv
/zbq1OkQ8XrbLXK0RA9e8KcOyq96SDjC3G4E20SKLmM3Bi1ELtUsb9IL49lFChYe
EuRtvhFNWngo7i/9LHZxxn1BktcuWNEJbfvdpYgki0dzqB+kaWFyhzPi8Zm/UQ0i
mHGb42tURHHv2z6C6hMw2+IEZwe26f55qGElled0ZpMkHHhwqkfCm77xhVjTiXhT
3HVH45IeWB15A+xBGcEX8ewitLNx5yj1Cx6BrC417Stjcxx6ASgpGr7VtoP9Yn3A
+ns6aQCs3fwZZ3ounMkIzqq2hjZQ88PmzMSO7RntuIC2Jq22Wopr4wdnEPaB2ui8
QlEcNEljkUZbGeNBGoMU3CtfXDdISj52ClCDIxwwIXlpFkN8pM3j0sgirweBI2Iu
i8yAEQmNEZWf64GFtBGikRvCSLPk0hrllrKcZw9AUNBm1PB3sQFLiB3PTpgPizOI
cDxtlOstFmSLaDHk5Wr1ZRdIgogKSOSKctdbLRbkxRFBG0gb1klizcsoAPKhhvOr
xLXbyVSe7GYE0sC9gbkfstzKb1BeN/v/JFb0KNVqb0UvbddYXMAVYx02gPR6yKAM
IFb/OekowL8mKPd6uVfjvJ/BAyffKMp6Q+rcKOT7jGd6rUlVlGOx+l/1FN1aFV4B
c2kn3vbLFeFiTQa8aT70DD+Q7iehrHSselAFlJkBtuo4I6nLXhz5+ml0+hMZ36xl
ojP9u8ZnH5Sn+cLnSBJtOluB3n6cAlhorMgqQXmmOigwYfDu4EoJJGSu/oLWkMEU
+5fVv3MJbBfM9NjXVcJCI0DG/6XsmeJyfNULDc4fxgPWNGZ6IeqahMHloimbEGlF
2O9+eXxe0oPzA9dnbcxiWasGTlETfWtRPI16Fn77x8epY1TEzudNWyfMr5lJXRce
rmv6LdF4425Sz/4flRcLQfZwNVidmHnwpcKFeurPhLew5dRStpO+gEXP4oXhsZXk
VtBGFZQKUeZlogJUTUBYRUtbKZwiJegrWoXCuFz4TLIM9jAy27JChsUoxyQHB/aI
JsuXuoTiRKflWp7yZFq2HyHNi2WegjJjC0IN3I0n1WD8u0Yt4BFKgGgnnRWgi8NV
RuCX5d5E0Adx+az2oBU20pYwIGjS5H+8z/1QP/NcLZKxmiwBJO3UgnkX5561X38R
TrdlnBlYeojo3aruKoIIXJfMimFMzu3wvrM57Ee9Tcu1bjPdYkAWvSmuvSFNcn0r
c2FTf9n2hTV062jgkgXd0Vom0ecvXX43xhhKBu47FwFKRN4Yp8IV6DgjHVsjThfe
F048rRPpujIdl3e1dvWBojayYn95RWfcquyMTEFeNlpdfYOjBDrb1VH34JItzLHv
aedK/Qu2cY5QCa1o0aL9psPfqFehYT8YeuZ/9JhuaPwFmpR/QGx8hklNdpugO6lE
UxGaCr6bNYTllpPAMtn3imJ9nVfHsCAAiuQhCoN7lH3VEsI/vlvRfsy2/p7NuwbS
06jNmmpXOHqwvpJxrM2KFHhV87J0OqJtsrv9dVCH1oHRdJ0MukWGhZSzOTFXIxeO
E8dvfpgMxo+wC2oXWcVDHFqGx3I1LjGJCHfiRQ3ZWb0QgtpQ5iCwB/ursQuBT4xb
YHcQWZSLJF3tKohgJc4DOL7SQ3eNNEONW03eR2/kn+ZMuxuXSn8cf4BLYRjEFDns
ItWiPl24Mey8VzMj+FEBBAAOeglq3mr6I70BMoqSlN9BRnVHzA+xnLPcw5YEKxdt
aI2vBXaERKnN3aLa1UiezXgKxppb8UNU9LsaEDhKeAEBb40YH3F4wu3VJHnZ233/
vwCWfTrvSLuhsZDlKT9aCSBph8PgXFXpslpz5T23ItHFyMjXVebVkgs72gB+RqmJ
KPFWcmtE+yuNAKbqS/1d72hUvwZQz0VXDVKkPj73EtEZylr43pZYbG7ZMK9+5+ym
HuWrn27CaUI1wSWSY/UWfoXBAFF/iPr6vgJH5UjkkVfRQY5OyizJ2HTdlQIUsKv7
onGVKda0VRJUtQ6klTJiWHmcrjJJbwz4KNq/REPf8a+6YX0OLbIDyEnSbdOKKx/E
+8voqS0jBDRZsR9JyG/1x2s/Kut/wwJedpcK0Z1kgAq25YRrnw5WspdNZP2AwF2F
JlVj5Rle590I8W1G9FyGGtj6aVjQs4rRTpvCTCo7yhqNK/72EDgDaUXXUy27woIB
2GkglG5K+KwC1cFusVj1n+mgSiUTqcpLJVCM2dE2REd3Jan65ObOAzRSBSnYaINx
KmLXqvxwlbxx/SWfGyLlyV9oAiUYCZ97MzC/sFvKyKNQXMWGEwYaFCX8dqiq6w/o
rm1yf6UzCaXcG6+VE0xmHCPHgAH8NmkObEh8pSlCcQiPoXVtqsuksqOBKC7tKOnx
zV5v1sjPX11QiJK3/Rw3cYlgDcCTtxPkOKhI6ivplxKPJWvddcvZYEY6nYzzr3fR
Ubnnq/IFV6rqsoG5Vpdfm2XE2jCo4y3FitkYPH4zFOxhZIGxUw41eKmkjx6CsR0z
Veyr3A4hZVC2beYVKG8I8nI2qi+6Tm+W+SrQ3DrOgauCjkiWbP7WlfGl7bHNLbV7
qEUtTLlDQB2e7hMuXrZEYs2vSL0y43tcrfhsE7x/lXd1XmQLHfd9ygRJgOk8mUCZ
XgHevBOqm/amg+IN8Rx02qke/EjkQej+3r3Xu6jFBo5/ZqUN/Kv5TemvqWtRKOlU
NLux2v8s9X/z9njWWsjgEtm/DA50KxQSpwTvdUwm1PJwNziqD26sh3YYsBPSiI1A
90dm+1nCO87PA5JKVrEZgBgfKfeK4OwFd/q0hHn3mRl0kSHfFi6pRjFpJwYKvl/9
QxcGvcN4HMOYV1reoXJccxwvH6CzfUyxaJFhgc8xA+vrb6pC74oJ/5bLU/npomxG
wq8seBpFmX6Z9vqvtDOtUFQXEn3mEa4qaXrKzqzlXYeCoCobNvEHbPFl7H6A4i6Q
NsR7uPaLtzpvqX4m7UDF4zw+gAOqSFcMWXVoUjHy1yg1lLGDGasey4DDcesZtkI2
vl58K972JBLOKVAd8GlMp5wGMHnEjKKstu9CA4OHkNIakxEu3gO2iabiUROWzDLy
h8V7eCA6pherhSUV8+uL/y1DV6guKXOtGSPxdKHuvLCIZRG1xNz03I/0tPhqFM99
AelZ5X8JWVE3LUWj/8QQYD7kM13jWJabM6MtzdeV1ALrJeVM+P0iXNw2M9kDRnlF
73lrnK/vyXPexAeRVo8OW81XtTGQvxfSnQlxzCyMunzHUfZHXVtC+lf6vu/ZbelL
CbzFsbw0pxb8HdlAgvAl3xLvoCCpfQA4406fBTwnA1UHpv1a5FZxGW73mfWhSDnY
4navBXDc+ohtv4NqlsdYBS0TK1PVqOaA0yU5aC7XST+05PKtgniU9W+ISC7ZAF6t
OVspeo7vAzW2mjYA0gqP0t1KGGcBwEIBbO5+vHlP0hGH82L3/HDt+tAqozlu2qQy
U3dAFC8RJQGgrk8ualftTHN8UaSNLdMGh3i2BqNfCgYJIdrH6p06JIBtq0rcOJQQ
OjxNaiwQ63aU0AvN/TA0/OInSLIm5G0xQ/K5MSpAdrKwgEWCtr5Bb24pr6dFGP3S
PWLkTX1bhSeeI3e8o98RuW3tDSdTbukm75/8VW3UQSdMNg1KeC1mCSoQv9jySQT/
VYveadegveHHB6wNa31pxtEySrBCqu04gtcpIj0uBlbIT/orriZCmXD4wNscKMwx
reg7vbW1aGYZD+nkXrRX82p4CTcyX65awjEJpug/gwPVyGf4uU7k7ZCuMDaRYBws
TmtJ8Outn7yW7NFPlOOQF9FzuIHwTMGVMmSWdTdp6813GkYIoLM6X51cpG2LTfOA
N7iYHxfCmRnJUXKNaaQWPy1103jnLAoqGj4HGdD/lK3VBAwBy8YEPFAPfIQ7Cyix
hyhzz7L8aU8uWktd32X+5y2HU44qC6vlFPeT57aRxsQKISQohycT4qsdIrr+nrPt
54kN+WahfGdyzeRIek+WAzfWst8NfPA54Yt7e3UBU2gJQwvJ7bFXOR8HCZ6/vscT
tahxDW8UFQyuF/bUCLakU7wX9rWw1EkgaHtLzYMKzNjBoGxpQ3+1qQ8vDdmTLFFG
Kw/HssprjqkC/VT8ey0Ctj15JWmT06FYhh3MVGd5oWBVpFoksKGRXjpTuBHersRq
VV7YqNQuFHniUSgNFkgu5LO/+jgiiDWxHG83ipWEm53LmEBsA85VteAbQK2TvcgB
9PTlf/O0csT159t1N1R9S4FM3bAecqHrIQbinDSJ1SnwWnHPiBXFXo2nRgS10iUg
BRGSesBOrWPCzGDhmJzqNyKch1HQYgPpI12NdSLwiX+QT0yn61vns3sOc2mT4NsL
c7UB2MZwAQFpmr8+UQYLCu6L6b+ARYtfKi8IggvjE4Tz8XR5zPubFMsWOwGQ//86
6OX97QeVbvWei+rm9jLxOZDudnA2POtKM51tjF4FKtF3FTXA4ZwIyJT1lyLUot40
Rus4/O2MHYMH5cb9nBYjwsyxz7Wtc3mmvOduN41Fuv1fXaljzajr+EEPmazDDhDk
RfW3qOYroGsnuuwG6DxJ7FuWf98SemNfQYseAEC5Skjoniiv8Z8a/WVn85iOve1R
IOMoPNO2ScSrSVNcFnJD1dF4iJRM6jPeCVFmoCl3t1BUW7ti1yUhAQCqGVDo7M6M
aro507FQ011ufYIdfYFRnn8UkTg5yHRddY1gYQXq6Lh2VLRKkRZIQyf4P2Mgnhfn
1soxQIWImeOsekPfHs9il6a2NJ178Xd6xKVTpwHkKODqFD6yagCwGY+629gGezOr
TjJ/4Udlg/Wc59I9d2v4U3q5M9uK15PT3ZuhSQA/9cAhjhEs0sUTAwhosGkler0W
gowL20cMls9Qeknx1CSUmPrVlIH/Izo57nKO9cZw+3hOePEw2ganoMHYClhpdUQa
5QTKaREuGpE2VPpqUmI2e/OFIeh9sQVnxH4QiUXCpJ/DRTgw5TxdlmfqNlkd6BMT
HxO5BRB7G86JtH7dv1ZpxP7ylGFnPs3B9Jb9Fw4zdiIlxov0kncV4NFqLRfEVJeK
OGUH/QMbIBNduiuoBsw/I/orW3TgR9AoqUuYo3//fgHp2bYsSIXwWPwOpqdlFkgM
tuJK9sWkiHrXCKcOnqTgyO50J9iw9I8q0r+v/3wicAjIvduWH+goIqmvSGvk4WiR
yxBx9W+tszk7J/7rDUQmKlxSXKoMtekQaCEH6Zo/nmEKHw8aylPT+G7DlyN1slMd
L/ltcF2lO0nfmdMGp/756YarDYKfNS0x38IxDrn8NpoZnk7oZ1FvXW28FkyWnUDx
qvMrkeBEt+TQvXMkFy2TGqZ/vsjFPnGo5Ohnfi1DYQuUuJ3ZU6KbXSmiUSooH+jb
sbkacLfvOWK4NqyhsExxQOtuODhs1E3ZJxQMAMCy4EBA3mEoYRyjbPolOAEcbc2s
qvdKof42dW0KehQm+PzmK0XdyOUn5Bz6WcoChDyindn9QiwYBepp086kGMje+zB2
amRDGP24XMz2LUlbQlmy13kVWP8wYFDaZwvKDJFUGXFFV27FMcLzPuG+q7nOKt5p
4Q5M42lhhfS5SxouVUZHePmmTaqQohGKoSmTWbNk4Js+2nB05uIXAsAGTIVxYYb7
YWQQ99KyAMEQDxyguKHB4toHqXrE53pRcRdiqgGKvpnuMsdMnhoYClRlhhREOHGn
Q6lVgAqQ0WYGw2oWXsuWH7bQpQTS843nPmy/OyMXCBxdOLnK1oNpl+URJ2jbeP+e
MwrAu/pSaqQ2WjGoSoaV/uVNk3J1xqUed63DSnTa1zN4oZZaOD9+786IHOUbflqU
hMrboD4eE877LxNhMcaKrGAEjtpjr5qhWF9rA2GBHgqCRlYBlmgrchxqxVZEfLpp
Fn1Wf7sGUgWE8K8XU1wupS9XvtrydVfhOZ3H1bbf9uTP4sqQU3MV60W7FO1dsM5u
HcbGSq1UN0Pjs2kmVe/IiwmMtJVSRR8XzzI/qFOsf7J9NAxNQedeXwSXkKKLYSyM
bv9AXAY/Z6yq3nDHpcUnLMMPuMq/2eMlk1z+7CBH9djFByYyj2uLEmvTDEj0Z0kf
F3/M8uvn8NDj9QZgCVxo7/IBizxqW58ckss6NObYoyQkkZTSao9MYs0HXr9gdXHk
BlPzHkeODlcJ3lVWWJ3uCg8pNAbkB/9YWhSDUttaRcWVoykeff2aPGe/45AQQ3KR
BO88Y3EuEljW6wSUyYTwCxt7n7Afcq8AG2FGQOG1iV5tLqm2hYnh+kOk0YNy+7Br
Bp1Au35gVg3AtXtproxuULXtolgsyrfpvqj6hETG/c7CBluu5oF+snsE8FwHBVRO
+LIoiP3ZnyrBY4kVkNA83u0cV3CGjpVFSzicN1oe/ABQvnaO7wJ2z65/mWlL+XcO
ptXXgabkVhUvajeMeXgfqUoFPFk/663VijX9rTEtB9bOcQ+jhAi5C525s0QslxuX
a6NNDkBgEf2gxforLECOPe3sawwXtYcNl8U8O2XhItyCd7dfppCNDR1M7hKnB2D9
RN8hWU1SJTBinFpmI+g8jtUn85pkkjO6yzGvLe9tmjAnD4m0N/sBzJw8FKFNgLgE
q38hqG6GXZ6wxdQbpBJ/fiNzhEisArFMG0eFIuWt1pQAInUIPtbddFXSBSVuMMnK
2Fl0diYEFlb7lwpNYmbMNBl7NkONcLVM72K8iA2FdwvL+QTnO4sYaBBENs+pw/Yc
AG43EeOjntSiSfHzRvDeD06Af1kc1atFtnQxLOdA/zfI2Ax+cSv8ikXH1Y5hKYhi
xkGBFl+lE4SmGsZ+qH4XtVXmpzJXUYryu9fbIiYI2OlgCh58+lXd8uN8qSUD4tYt
ha0aLI26Vhgf6yiEgTlxhqFzobyLkYfjr/oLNbU1IJfmdiPKC0cReD9JURPDEUZY
x120WStAv83R0byP/FzCAGyn7mNQtq+ulzfCTGLom9vjxh6bQOoTNySBjeMwzrZ9
FNj+vZVYIo106yyJy9qYgTNogrRuZFg9/4f9mBIq5JCsv/QpzFsz9SLdC/UWBh/h
R77t9BcM7/vWQ3z2Fu7kFnjILyYk8DGcLHTfY/yXdODOuIQay9fKuPqoiZ7eRW7K
+3/Jfq6S7litJXjy/6m2lOAwPGs7I9WzRzZzp0b3iZeWiordLNmgArVu8gNYX4OC
AWShlLa8MRq0OV6RGXnYwjIVZF2zdVCDzzxxHoQ5cVCb8cqdnIsVbt721Xkokv6p
PQdp7hhWjU4mgYjWfUUbpg4hHsi2R7b7spyVa2ekABgeX8fuDgNJsarU0mRJoujA
23YoOH1clY0rmV/4L+AeCyUEoZVMoch3nEv8WCZUTgqIpGaTRsJA7vCXCE6CoBHj
7FrlXUyIsZV57/9QFoig/4AXUX9zCunJjj+7jMOmsbv5M+xjh+f8E296olimjZsU
ozpDIhldFDcBgOCMMRy3HI3cimW5hwMzoImTeuy9RCW6/Gh6lQwk/VxyndecPezH
mS6swIS+wM24hDcpj84Ch64UJ3NExr/lazbjlGKcWbekMFOiPpzbO3VxmwbuOhPo
qWlAom0lm4MOC4rBrFaGQUODBjKoKEtw4w4SGq3+NtWNzOBocxE+R0Tpt1JXNBKa
CKlTfhBytnZSjequUZiwwGEnGZsdOigSW5xJNgquBeKMiV5Pe8a9b1i7cLcU1uQB
GM3yEtYl6fbGFCEGAPboV2nE4YGFrB1QErjamWzdRA3ymNWvCFiQeiB4VyCOt5KB
PZN3PiXDQdPEutgKqIGmnY3B1UR5lBAc/QbXaK4eQdYz7bu6gZhL7nbfMjLvcMKd
t8FvRceeJyEyn3rOdPXZTwkmfobwEfA6vLOnwmBzLN9/tAvdfk/3LAtBAY86KaiQ
MGs5AFAPkj06V9Xc1CMORkWAupDzMhHYEhNgj/Ney/teQNMkWBtRSf5/+nUInhzC
DKLSVyGmWsbKM9boqVHPboJ4HAFiUAbj94miNteHkNjo4JCtTxKv/9JhyttbPp9i
toBK4di0jb31jkpVIXZVP0qau9RT9jX/M/ER9aQIyZeQjgvuoCP4PO+T6uXJDwLS
p11Ym5HTSvuYkbfMLSrYpJNJSGOYTNedJf/OrZ3Jw28hYLFx/QMC9j3qHm2fAiG0
Pk95OSccaHrD0QgVBrdZkauCAackBFc42TMYaOGMhbOgC3Q11WBT4E/pmbqyODVp
WsAKGmxPZ4K6qvY7d1BZtaBQUTlgBGSWYPSIi5H9ptjHXqrOpBWMGBRT96ofONZU
cuVGw6ti05jH1qGhGhiGm+/Wf9qJRq7KKVtXdtzo25eD5tGnVSmOu78qkqK9qm+H
bcr5e9rQY3bEDUKDs7ufaHhyhzUrOe7QFYHH5IDiHvchpw8enhmRA5RtMUSGF76R
R9cvkfHDKPxEjs7CmgKJFuZrDarOqDWLBYVJqG/sxve57A6pUHTZBK6MSJGNAIJg
CVpwt6uMGhWsIZT4IgGyOcqELYifYhttV7DO5ajhsLz2ARgqD3e01J/BgxRFZYJQ
LoJdvru2HBqrHrIN0xnDfWNiVlTtcKmKWk8ycz2uPSqYykoHP+6i+IFmCwW7ef94
fjtLH04M/5a557y3iG6lNukzk5KeUees6z/7wzzlAIYMnE7Son6p2bcjE2wE+BPi
hMOvuwBjNlXGDYkcuMGEeJTsFe/MlZstK2fEopDQzDRKpI9SHM4T8Sd4Hi35NC60
MQOfuBAw8iRemuSqsUB+KnUup+yPguo1nOJf0OQn8OVQCFiHCfxv8EqsZYnVxuV3
qAl7N+8g2BWjOGfN66flkBY0y5NrYitr4cm3qKO3YaOV0VGr1jBSliyBKx5XUc/b
+/qSyJYUsBncuw3kbA4AlUTdpkJOEPTX12PZTR0n5PKV6LVKy4xdXP9RGh/Z3cBp
FOk8hs9jHLrzT+AnffXlZgKxJiJeyIJcAHXPpB6VLqvLMGn6Op3+UdxH4bzybtYP
IQPuRm/eubCfjki43MHxfS6uJrwh0FzjJNCxc0QJWfHUcuPtVYPq9ei+exrcQG8D
4bJ3/wcqvWC+qNrl900vQ/84qhpKAIY/pfDmabErrOO6ENB6CjgEj8qhTqqrr3yD
scTW2nyxzah4qr4yaWbdAxbffdT7h5hCdd3n8ONjoUP1pYNqhVYpfFJM0W9GMsLX
KjtB2VdS8CVw/Dz8HAwcbF61gPFXO9aQwOXWGRwdqXAXoBupVRF6aHB96s/Bd6qL
/j64kUiOIDLnAZuvHHtCYl0GLIBopyiRAqB3dxQPm9QxnTGzPadMUoozoAMaATog
BKrj7f06bwtZJrcbw/AhabyiOEoK1w3TrcUPYjK5w6s8nG5S9vYADCXFuCT2ThEl
Ob5gVIBZk1+9vZU4knJh+xxSaAVLR7acKfbmXzOJ32+9u4qV0HzxL/Dv9i6+XKTr
LB4OeLncK53AjiMwU+qBIfSQHNnnOg3l67Okr+ToaMJNaqEdVMCKxDRGt1Mn18B3
+DcpQOkLjHTKBLGTTVkpQ0d/q30bD3IkJvdtmZTGxS4eG8+1djuKAxKmtLJFfd6g
BDQWj0i2qTjLQBA33mbXcpXr0Xlw8xz/nvzttgffhXEUpj5A1izJa8ontoQFiDXV
Zt0dtQWPypQVpXqYDV4BbjBzseF7Db4ztdn3gRlO+6EdfHuvLFceeduDXDcl/nYZ
G34XffjJSluZx5q97JoeQOGrgmI1p/7icJQ5t3PMIm5WH3E/HW1D94sZ9/yXbRFU
NFiD0pY1OJgMdmpNUPoCUkWEs0rCo6nJ5htmBv/VKd3TSq7bwRu/3+pOZzLrbxGN
7KN9F36aWeQk6R6u2eBHeyYwkG65S78OOUzuRmmSsJq3OzQeadsqJboAAF+uqkgR
Rm6Zb2wL1BOYo+48+1OMUIsx3LXUW+EyA5vYkKmD7LpOoGr5MqpivTGIHplpaz4z
T758cOienlmzkoPFVp/jT1WWeUHekAIEvridBmF9YvbhFfuIZXbdOA0s6W5T3QJk
hVMQMw5Dfi3XWiibdQnFM+Ne/at7THaKBjLreWsn1C6DluyHXrgKNlgoNVuK14IZ
JtpfuZccikVt5E5KvKYUzuNDqqdMnawqx8WOxg+GL93ENO4AXrYpJvKi7mmUPvfi
W7Nt60tagwZBLG3ds2CE1t5zITVqevcqwPYp+UqvumtLv5jXfjJq4WAQ5AoCXM/K
T1pRaVTFBN2XAboFWAEo2U9D8m7NwurV4lScMEyStOYpQsMFMSwbw3KkL0YMEBHW
Rm8qyxOcLyvUO9uxSibYhGFOrXZYKZlgQtT0HZTdwxFQgIECEbEALttOOgoocvIv
Wq/WSOIHzODgj+/sov3vQKaORSC60O6pJNabuJJSqicZ9Cku0nT5NsaRHwE1wd7z
wF7FUocaatDRWrIsnJMl5X2a2SAs4Wpr3bpnrAx5H8aDBztTCgRBjF5zav/qm1fe
UNCn5Ggn51sy0ZmWhVlBs/BEV7s3kocPABNT8Q6LiZ2SPA9gZs5tjny7zntur817
YjlEWAugVc1oaPj2r+ou9tAz4jQLdTGnz6l6Rj7S+J1+tEia1sN9p0NE0geu9W4D
Egl7jRfyIcu8Sma6GgBZPXKsBV07FylTIQ1IE7qphYfAjK7pKJXtCDHy52Q4hDIp
1VUST4rLhVEdJQASlgbAFk1YdcW6yY/JTPfOlMtQNX9KtElsim/nN3UfCA/6iwRH
Ylzmy8oe9jGF1dmCkMAZGwxTkOvv8HxrrAinl8w16rmF84ffE/EbQ8f1AerKDGYe
Yhv1c4UsLmDW/iJKbDqyNPYCEme2ej12eNB/Gd0yyQITFZrY0frWF92/oOGzEwok
CqzioBZVz9U+2Wht08+FB/1Vbp6W9kAaK29aMYWuN0Vhqr0XjbWEFbZaKIFdZjIj
+maekjCZ+pGiNpWLd+cg2W07Td2aeqZZwsXWHrcqmRl+ZOjmUDIE2BlA1AQP1fBO
u0gre6FSjkxWJVV+af0kEdx5rq9pnDL2c+OogJWmdNPGBAM2W8lLMhSuOLOpkw+c
cZ8M0i04PWOlRcTQasnyf87EkDAxCUiB7X1lFPEgR06luz3FEIcFnI+mReuxYJR9
Es1R/7UyL4Zxttr7K9N6aUTu0O5j2H0RAv2Z81AsH636Tr0e8Xk7/b69TcH6rz4m
HDHJWGJiUBB7Sj4sv/CbJKR7HtH5aygeFkWhImdGgmm8nN2FvaYgciVJ5uvfNcEm
PlWh00r++Ku/rt/ZAMdHCrcqVVVoDhdNn3UMSpIkjfxgt4U+aQv1YDfN+WdlMNGo
MTsXsLxwKzQWQkhALlrMXK21xB4FOJcGIapcpT7AtVmN9lremw3SiLiUGV2oe3vM
s3E5PxzZfLgEgoTaOyJV21DxA58wu5chJ4TtUxonA8AcLvJELLnKbyh/IYdADoLU
nLEGXT45CN6BcW/Wg9qknQWKZLNLS/75FmAxVB+FrsUfbWYgaZdEhbzlpe91d7BE
PhjIyy72k/FMgV2INECxFemid6vwIE51ZBol1e7di/A6eaMD15E5/dCYfLKDIUNQ
TIKTTrRY290tpMhaI/9w+fFVnbaMlHW3Upm/e98q5xDE90lhu6p4W3VwrMkRGa5f
YU/pzdwWi2+SjWZXgzQBK/DcBmSAXD7OIm6cRBBiRYXB+ggJaplOLbw3blBLKirg
iAn7gGHz+xreml3GHOB3T6yLUEvhP5zgMHjgSqqLn2hKf1+EDmwtlTWzBiyfMfDp
EYYyFAxyXS6pkICwjzr/TuhvkfSXHFcNykHrhlunCFIRA38Wlx4hRJGeBTGOEwwq
LJ5LZH7d26abdQJEcYdyECMSvFsqz9jd6oUfy36lW+fGgKYu/Xkbg4HehhwhEIaY
wKB1YChBnpqclIb9t166cDfdLYEYvUA+DfwaEWx//sQ2jzJTBUbYkICUlFNs1PaF
PPOBsYcEtiKXTV8bekH6TkBzyewGK6WFCFH/1BoN1MeTAKQLMZQHKvukjqrw3ymT
82eSlMbR+wTtTXtROxJ9y2BPLr5ltbDMFN1eBkFcpiNYa9P99iyyMJNyKKpyM0YN
NDNByEPX7ebe4dJ4v8BaBnanW7ZmVwYC7/WDJDvKBGUQaVunHWByeRIwwJzMK0KA
gWHL2QrKLZaMGLYuaBk1B9DgQWyXjBxLANDaNw3TjA5kubhWD662mqlaOiiPwJX4
6SgNxHQK2U98l3cwsavIZaz7qK7et4vdfkPAlny/VPRkF6xW82zwsArImQDjpY1H
7TweRF4SIhBHsC0EcyQdGfR5vSjSk36B5JFaCh0rEkYI/q+UM29gYo+ImI89rPy2
fJsVjFpv1W7s/U+lMpTs2tsR7Sl3a9TNILo5nh6yk5uuR7UC5kMuVROnsPFpmI5c
wNMi/dR8cMV8HwDnrR5AurTpR82ltNA0SHNO41peCjZoAdiLPDxum8DPrrhsLRCr
9NpT6qpvPJJHHaWojUXbmVuXnQHfD9W7ZB0t+FXaXAGO7B8Qo3eVOgvXQfkWUmfe
gVlzwjWy1elvdPHJQAHOrYG+TA4YVuenDoKeD27yyUIxG1ez003oCghCjPLrIPqD
r/9UwARXvZjjxQyczv/Afu7NinTk/lu2N5UimEmMqZAmHFr9rBmcCTU0AoBpql/A
NIg4w5XfQQg2GOuCfzKz5/zWPgucFEezUulUmI5zmcio8EjgAzORac5EbsU38F7Z
SSGGgRyHZW8UUd4lUfKOibZbZMqW5xPXHypujrya6CHdVks/zVTUPa4EvVdPS+e4
gt7iZsEnZKyTWiyAVFTjGhRxbCjKd14MIOvcjbdaIfzOnVjd96VazOliL5hTdSVV
t9IxOPHi2jCP72tAPcrw4MUOfOLCKaSfQVIEVnDjz09pXFWT65L0RRSBU0WBYYz4
WJD1Q6LIb/VtZfKIiMzTmhAnGxnlHeogS5G/Zslyv/VhFAZLtJMbSREiX3+FWpGg
YLK314OqiZujKDGmNQKAoIb7sjX8XVj2k6HUXIUy4AeiiLS6ATzWWFVqkff6ZfxD
2u/1sAKl2EWXhtJEFXXhQRrIFZIyNk2kRiYVfC8OJ5YH59WG5di8AhWQkLw5vTpu
sjwXEnAQijSp710FlOHbXEgtN/mYD56dfgem+JzxcfPdCABtPR3sWGpzCP7ukdi6
VrgUJUp2Z7fpjZ4C/thpvCvk2q/QZUyl7MgwyDnCUzW5ZoTc+vxnWqN2LaXrmkYi
ikrrBZDwEwyYehZgNLaP356heDRYzPYOoH06+B6sEAc0356OAlwDNk+KsgWm7vpm
1+lCd16lNi7ZS8e4WLlrlLehH0NcTvuEzvzNiHtnyu95KCkBcB4/2lbOHAf0yVNw
RXAO/vDDg3lJVsJUlxThDjDO2uBfTcv3ZblaPiUjnPNtpZ6MA/ACwcY/ePwswh0F
zq+Nff4A2urvk0peBPWW6kkn4PH73oMvglw2iPyp/VmcxUniZ+wGzpHkmSEFgQnd
gL8tkbEOsvmVJ3Q5XhZ8oAHOtfB9swqzpenWosNwtLQj/N/jcIkMHdxfl+VTvlFe
GJ/74V94XbE9PMUndZ8UF88/riOkiZfRgo85oPR3dJZjFGg+dqrstxPYjwUFvPPC
98h7xktThEtlRhu8Wd+vl3HnhCwhnFcmdhgV01t8+RsekxSrmDIH01vNqa5WiEwU
zmtYUCzbPBBZJnsiDDcN2V7qSt80hN+mNCQ58mT0OOw7VYtuR7hpu2XrBhyRj+qI
B9an1yl/lBpJ1AEiqsZu/wv7KStSYAx6mds8LXYtOJJaMLtobFbhPha4tztc+ACf
5ODwEUlp5OTxNo8sLVJVeTltqxudyK3ptJSgP9/3OW5M9tDStMykgYOJwfONV5jI
6xjPFA4dBjpQOfY3Sb9GtZJDPj1CQcW7UQemSE37l0uNOVvujpMnlH0MOSvxFhWU
bkQZWDYFB8HMYI2dUBXLinUlBACmbgNCAwYjW3KsugoS3ctLG182GoEpimpIzakB
QsuqxyqjyiHUDHdA72os4coCL4L/NZUMkbsmSnyLswd+tXympfvSFXZT1ORBAYmk
O933OvR0hJTxV+12szM3zMfqqSPfC+BcgJvnp14iPAVowyldpO/z+xChwIELCvFk
YmNTNhlxDWQqMCd5z0uk+s2X/dC0/7dq+o1k+BAHeQKKc1RcFVJ4Vcw49np7oh8J
tYDjfOPpQY8MYcHgvh7hfbPLdRv08bKw1Vy+Udteb1jECJUXq8qXB3eR+JNSzOGq
D01ejCT3lYEPqplaofw78NsXB7gbSUXnlnv5/TNoO82GhjMDsYlHpyR0QSw179J6
sSkQP80W9TlaPVnGrZRIkbRPfEymCEmd58hkbZTdf2peioeEeE/pKA0KARx9xS5O
fFjwWZYvZHAqs5sBv0UMDb6RCeQGdkhstSueOqQHlOe65F64CRcHaTEs9DKlSZ6q
+eYeq2AU+oKBdLLNDKuNKmXcwDYcLpinTAcLGA2QNao3TKTWTQPAUO5Jl6FtTAhP
UJRBYtzmFSWID9byPD3DJHJxYk0ZhhV9wNB/+cxCrb7dCH42azU819zMO6bPs6cW
fiE4LEUx5RP+2/qQqMhANYwDdsqaq/r8y+EawCPmaca4JO8MGnaQWzXPjX/WafvJ
ffNWmutG/EAUuvgCMd9CksxulLRBXJevSpLAcejeufEk8FQ/eO51kJ+SVX8BoFGF
1Nm3ePoNPWnxx8YE6jJh7h4Qp0iid5gyk/5G7+1mSYDyitNGgAT4ICJY7FXeMkPH
os5GoA41QfVU1ddl+FNGvRgIf199+CWAMXa+eUSiVWNN2ZhF/MO/JtSHjG4XIF+D
OJX9/rYKVy5qcDajtCDS5psGWJwz9mtds5W8EIiYjBZ3y89fcFYXhvDp1n7Wap9v
lZ2AFcc7A8t2vwzdBvRwtQgxkyuSIjKKrD1B5+8Zke8Ahc1fSbjHFWVdcD1mUCE6
gb9KUTYKmpipsQiFpTow4XZ9n5cKdK+m6s4M5TTWGk+MvQHXSjNmW5LtXFNZ5yce
Dcd2zsD89IXTSWAmXomCXIk6ex4cM7hbmbtySBhQz498WUxCBSU6k5MUrGxPLZre
00vRJZyJldYQz5I80B3Pa4F2wmcUksO65P2+hBC1FfGZLGa67YdXIsGtA21u4KUe
S/S1GO4yWMqDMljJvyGhaqjLlxI0O6XeD6imtdVnp6uhw1hIr11020HJukUrETpZ
yUJrmePmz1fSwdnLciSeGFAddxubZenwj1PcmFab5LosomofhCp0U2MK8ktNVWrS
L0/3m6ylSJABDLSQ6w1aEW7YG9lDv94m9dbYxEUwFd+kONLQjpmsoZC6d4g0ERGk
c3HwSC0OFL0Ir82nju3yrFSesvXz6kCYWXNpsg5Hl9o6rK/bbfgOL1UPCCS9kLS4
IOOTvGJ+YfQkQtU+X4UhxFgxFScLMEZE8FtSK+Ob5qy5V8WJeul4YLNMWfeksh/z
v5Z1thEr+A11p8DdpxeotfBjG5dudoHI/38VbNvL6eamxRpyY6gTT4B4Fjt9qKF6
i1HzmHLfUON5FEhyeGk4/IGaSth1M7pLGgzBqFZ2MI+BjiFtzFBdub5vg16yuWrb
6ofOLhxRHeK5uqy3GtCX0dTGDgN4XVsgOTHd9nA+Fl7LU0Ne2FCuZrF/k9wzZtU5
W3dWICGgs2bQ577ocyXkb9MHnuVSTHDvBvfxXHzvu/J86FDnYoPYyVp3sUGAjJCv
TowSkqeR5rQ33VHF1We6u5a+jBOLtcjWjJGXywnDzgG2iapV/KQGF3nvtbEKg8dQ
ZoxphshVoGUNI6BDDubw/6o6a1C5y9Osuh30wjyvDDRaKw7gcsMreFzAte8bm9tL
gUp1S9IaN9Guq93sFzjLP3sC/esWl8YJkWSGmk6aDci6KqDLu5xuOK6GSRyhyj5X
1qN+yqjjcCyZcCRvvVpZ47qHLXXcfNq/2gKheCi7Sx8m9dBQqAswjcgstDDZOU+6
6Z2MMIr6eCzbh/IUWClhji8ENKZBpcMu1QxeP++i/bEW0jFTEDKG8F5Tnvs9Zojd
1tNkmmiGeTsfyX7l62M+erR30aSRQeyt6cqyGousLQTcSuKSPSLvp7ziTnYhltrA
rvTFpsBcofLogeJvBQh4vePrwXk7lEqJ0rbHT9SAxGQjFo3X5rTgYjkEiBS9E5OH
dgR8+HcXxKridfB2n8V/d+DL2j6QLCn1yW37dziifCI17yEd/JD1Btl4ZnHPqLfb
r5IrhXKsbSL1TJ2RFdJo8xCLFmw+RKwyHrnteJByIB+To5h5q8SWRRHWGUK4VZCg
5TOW4L0BkvXOLSL7RDw3FTSxVcfJdwGLDyQZpqOKMrabawI9S+cFj8nJNHvTCN9K
QhqzFlJLT4xqYYypluw9PvvMM7BcLrpDd+WhTqqj4eSjl1ox5UWP/MnT/04IPAFD
opxHu+ulSdQFSM+iksmzTzJr2K2rJpUsXrqN+SJ52bOVQuN2rmIowem0Ez5nTpN8
AwXP5u4JIt6Nzsj9IXHL7C6pctoAsz1G24h5ip1iJTf+XA7/JnOj9gNFFi/nXm1r
wdqdLYYDgyDa6vvsKtSC+RcnKpTDmqL1qcqGdXhUEhJiBi3eohMDVCA/XjxNeoCY
2+QpEQhXCc0QXSLUtS6w0mO7XTonPtQhJZcMgR3Vu09ynS9iitMZNpVmty1KDTfN
It7a1uobm21iuwLo9zJG8/a2K+nAvKZlRDKTIy+e3oUPS/UeQpoLSO12RhNNNM4o
ukD0hnpSWSW6XAHXul9cbUZ3c46O9bxKve0IPbZ4oTXeZKBXTd7Prqx7iDe1R9x2
xGm6s3YzaW3ScWkOddCjEDaTCn0Nt4weJw2AOW8xBC4UN8DYEAJ9Rov7YiM3Ie6a
y9rKQSCkHlxcWHkGJ3M0I6Qu3rVB+PkNk742HQNLy7uKwC59M9eT3PhY0qZBB5gS
er3RZb/JMZol/kffGNLmq5e7MW2YQVJIRBJH9rhQ+51DwNMN6G1++iHBYz2j0vuZ
skegySY7dDDqdXjyu8+OBBvj1SZMuK7Vf1frLACFSERZzyuYMdNBxz3BLSVjOTLN
mf7E6Zc2kYgmxisDyULQOopPSQsHSSBaoOwJcYm433pJzVM4A01LxBfNdolZ+Tg3
5nReMzuWjxIC9z6ODpJc3yzpsE3tH6X97+z1fZ4sczCHYxYWngEagMwtKdKZGol5
xr35BUWrDUdt7RoxOJNDGFW6WG7qWvBjVwNrHfLApk+jwsU9wPHshOJRQlgknCiG
WxJSkrJJP2Tb5kaclv30ga5H0Wac0h77un0MFx0aLnkWtr8zj9EqFMBPJKTeEGsA
YvV0hhPCAzRNnUHdJKLSyv/mY5SWYtXBu+kxlaQYm6mhjAe6sNqBfkt0TgyUYV4l
/lK5eMh4MsSPmhdnzKUpa+4v2FouDerzfyIvMYb1+U1YJOYNsHrLRylH1Wdg8P2g
K8hIP2cF1sypE2wb0wQfedCyIntDFqV9Hz2FSe4UFnYkZiuygIRyTBY/YR9DqpEl
AphDdDEItZ7XUIlINcAP5ozFKzm0eZ7mAYL6hv35VEXJqcd/ZhJXMrhnl53M8kjP
16zxAam2pSbfv2AHJHRYZQ+ehDNbcpqQkKivoSQi2GdgCGpaE2XkEa6Qajfti69Y
8BH3CdPHTqeb7n7QP0MpNBtcWZ7CamLT3/Ux3cEtgQw7r+VoKyLW36SZdJul/8FL
KwDNMOaGQOCze3rF2LUwelauy20jPyIZ0LJJqUCLiFYS9+lRsjGm7l1oWCAaX0nu
tX7A8zbVHO2HY2J71orp4ri7oXTKPwr0rELt/JI3PONXja+5V3IvHWgV0gqQwDs1
ekKvSQlguKmm+SXT/Oyut3d36Jzxy3CnDxSPg6PV5m7YgPaddiFYXTe3m3sq+ZTd
uTrJqy96ppwBCrW6zkp9hz06RdsLzi2r/aQLcEZwcGaeFJx7qzRNMoZSXmfwvtBr
xe1XPgUq4+YUp3LeKgfH0g0DqkmCPhl6cfSocmC0d1X7O9Y2SCFppBKnjXTRvTkB
7w+emI3DXEfvO+O2DXkXbpL39MMUJuYncYd0Sy3VIuBYqynOTCkkQtqoWCUSmTR+
LKHBoYc00mxa031wmcftqu9XmTJzQ5jYaNWJXjbEsqBkJAbkqBEgg4L8eFw+XrVh
kcLef2Nz74IGd6Y3LsVJCiaMp5op/zBmX13KGpYjStCJhYbM/mQ8x3NBHO288DTH
cZ+EoBcWMWB4JpZ564Wi13AM7xvTkKxoxg4YRk/wCWPVaVtcighDwS+nVApdJgQ1
m1cbUZqg8aRdgVq2NsIFbAjaBOEquOJY3Sm8GKjPl+2+cvEdslRypak8tVMbDF7v
a2IOgliHP2iAmxTBHcpWKRT/gGAFnsZOp5occlj91oQ9dvHU+xgNzH++uGl+v/+a
km5GJ+UW57Q7WHHQcNSaHJu+48/CmZIg7Ool7EIxRyKaVlLpaP9byPAGsBhA9uNt
x6EmVMs7v0ZiD2af1k3a7CcD56xpVWw5If9haGuWu9SCeqOKg72XJ7So32XMlPZW
yF4ZSXYj2l7wlMk/6mkfOBzWoywB4kWEdxlNyL2QIsefyRxnvk2NcLB+WbiXJIId
SRk/tp2hbayCkh+a+jX1HvmjX11zOBc4VCTLouNxtC6N+ziqD56aldxTOXoZx0CL
0YXdsEEcfbsl7wxB95MRFoX4NAkcfRPr+PNB+r6dRy2VcOv3TajKObW408emTDmH
gN9GOQlZdDoLZ2Y3IaQNwaAdWig4DF7yasRdXg+scpVjiKcbnmbi8BdjWal5cpjL
n8FCxFJ8dIT/pVdpfYv6de5BG0E6zU5orPYIzkNtVy0g4PxatJqFtRTFQri3dMxF
n8jYu9I++KnxvweKwF6Ua7x9bTANdkHM5jISNGeyOZD7/G1DynJIFL36lekuehu0
Q9wTerE+L6Z+oPRlr9r60sFtxBDn7np98xcVq6+OEnS9oqYkG2Wtwt6v+MQqkGBP
yFhSW9HkAQPCc42bVHsEZcsiHpJYvT+lyS2EuqSHzR8Mju5IEPt2SABeeJz45NeJ
OTxyPwqvQu/vi63N9ApopNYuSjSXew9Z8dMes4ndrcWVfpxzhnqHycKxpC1qB1pS
G46BqNFgDw/FQyD6HswvEIcnkMRKq22Hn1HbaPjcbwHWC2ZiER5GB5PoAZYglGWo
17u5233A/lJdFtlu7mBybbbHf/6XJXb/dRtEnEAmVFGc8jfeDKt8UswadDCHsTRl
HkrUjN4IG9k/Om7LT3h+zs7PGCOhUjCecaGmisuw47RQ3ZC1khoomfTVANodgxoZ
vtY6Odq6ArL65bIbPC77SFE/IE+3deE6zpfsgTiYKc0QxxRfVa2k8ngeULi1zHcE
+m96EU+W4aZdVTg87RvT2KuFuOC4G1cp1Z/xOePuRVBcjyx44ZcRq+in1GxTRHxA
8NH51i2DA3aICxduCRzjyGYe1sVbj1TL7+4YMqLI6j3/V4a6x2nSIiT4pzabcYYZ
A6tLFjZPkzHohTbaNQKrLRpUZLtn9xk2ghOhy04x+1DjoTnvkVPg5UDLIr54F9qj
AoZjPHP/KAtMLfIGsEZo5olO8FwL3WK0co1uqG3kBsGoFxhR+oBES9oBCOFCfpgS
z8LYowypISyRG6nw5W908YWVfLMOEQxvgaBmyX/tNJNzX4353TH/BhnsmK4q3fhR
4DdAQK18h4Dv01w3GVp8B7DgWeIO7D1RnWAOfifUKpJRAE0bLEaoV3FJOkizAL2I
wqsCVOtBPx/31H4nito2wQk4Gvebq/mHTb65cjLLVbPl75hNtz4xoE7oAU+no11K
OYGO/HOYrSkKnBz4Tb5ZywcvL6FKK4Fw1SQgeElCFWHga8+6o4Xgsuwd6IbA1cDk
B32SsjKDIHPMcl9V5B/nG5KXefEwyhtG8nNhUNh0tZ+JYGuR04IuuBMYNnUPP7De
vktDgQjAd27DLV5d0/v9S/MTCAqKu0Ux75Cg4hegLXFHnIOFT15TZveOyiv2hk9y
KtpxNJ1dQ9fNUvPWRI/1Nz0xezIWDEPHFEXvh7ZWmHMPwvgJvck4qQVG7Jcy0zFH
gB46L0ESRtD6QF5AiXpgSETw0Tp9HElIRT7yd86GU+rVEpiSFGEFBpwW88cRfQxy
14TUo3tfxoOhTrg2bD1IcmC/Fj2s1RRPPW2150b22GhEP0q+nhramZdjpMTiILC/
4qWnTrP4RuseDeI++tpc9lVKWrHnSWThZiSobDSvgr4fpUdpB2fdj20JJtRLSF8/
SL+9/1aW81k3ktQ5920IAIaOax5dFNL9FUPIwqjP1KVFL779KOVryVRcxMlZ8xRS
JF8kO0OqM/TFnCBsUxriKKpfuU1mnd+OHN2JXwoZiSjNKvIUgK06oV/vyK2Vv1MA
oT89lG/At+wX7H8CibQfH0IA6zcmuhGxqhO1FIAl4cLvZDXiSm9mV0KnZbxpGlZW
M9ePE7dMPSbYAJ7lrYMmkb6j/3eHYg6GvRq8habkPhI8+yKCRqVYfmMylU0dUOo6
jKM3qXyeEHZ17aK1QlvXPvzJJgpYHcxSAanm48h0KooOl+dB1c4Kfa3F1kMBeLwe
xPkPyGnYCnC9KUQVaUnDOfKjuuDI+emCbAqGgJaWtFSsHCiwk+Ejw5gNUMbnUHEC
7rwglkE1KsLgUFJx1GdE7VXKPMk+xFFFHiWJSZR4mMdem1siipM3RAiDZAy8+Xax
DnF9YN/xYQCk31cpnEdctpLCqldhM1bTvyPBqaLo5Kvnds1aDbTIdSTOyJMOhFGP
FaDNULcTlbCmg9bCpXa12hONcLt7Qv5FO36TAplvEjfwn17UJdlOCWee/J4iWkff
FR6tk34rTZGhoVnUwGyC7osrWH2gGSV3snqr6TiyOSRsx8zhxKu/sy3Z0pnuRxo9
gAFVQ0+fyAYnsHKwPapXZPqTs329pAz03iexcvJh8PjRkLSYjdy1oKN1SBvlSwBH
aYhJWAzP1QsR/cuHHrsCEnmZkm8Idwdy6yqZrZAB5+GV6MpETE06a7PKQAkuZAvR
d33QgFC9zH00mFd+gkd7M0DkhNDE8ILkqkmp1V7B4RyVh4rIL8ExiW01ZQgZMKL+
0F4j4BvxkrRh874N7KGtEM/TFHfmrcbcl9Wj3ouO43dQk9OOpZakl5idHtyUp481
/kT0Z/5+9fQOZLeb8Q4nMnoBlWBh0UrGQOVdHBXeEeHY4tZOsEajuAChetHcDHWM
9eElI6u+kht8HhOrpbIRrA8SzYjHQSlXhIS15e2uE0TTCjSEoLltNZN9iDRD6ecR
bjX2vMGsrxaKZFjcl86OJ+ZKIMXv/9pD1f8+TmUdnLgFhwMn9ZzxjhmWXjOH/zKD
GIMJ2Q1Oc7XMhBH0i1NKd8eW+0q6AiyY2V1djVDWRM9Rc2XuVM4GBVIHDDie7udE
tXOGLFdB128vRt/b9JbP+vw1KY0RFMCi12XauME4wYKGQANa+GQojHXnmDQPyMGl
V2WbyrRhm3B+Z0DkMRTJDzeTuJTphs1GiBoBaUHvIMQO3XzR+/F0maCQVwO84X+q
AQQoWaZvRDJZ97a4lCj9Kc3QbM96GFKVUsITq6inDhWf6kTeeHUi47tahHqz+hP8
jyd+LS+WvquqSVDQGW0RCJtMq/kBkmC3RLpzxWRLGgd0VcMjvDE3ldO3H02H0hKI
YHaCsz9tDf4R0HTUQtNgL+Ad1H6oh5dehgQ6+X7Fiea57eLqx3nHsI2r12fMGMTw
N6voTcoI3poo/+ui24ajDqa6JxN4hfwUUct5sz8CIKcyOPMihANiTWXKpg7ScV6b
sn3rhT7XCaW142wswXjilKj5gVpOZgZJEtx8SU9QL3EW/+KlNcItiO0IHpVyHNgm
LGOtz4jVFg3Dnskks/ujPMuML/bph6/Fq+JiaYVx7geaWpqpS3fa8kClhQx4tNSp
0XUpRRUdajdBQqBVxBR4ll3tHQj8HOStZ3vpXHYoCB07C0gwe1H2EMC5WGV8cfaJ
LMs7KuxXLoKGaB6WPDBQYg0SXlNRZkGzAApZJhRAhI5cgPdoOKhg6ShcGWu6sYOD
xVDipN2G217jFZ9uCbsOA8YRr48WMbNOafgzxD9fsySMhKNK/KQ8fiadXsmiNPLO
Xqr7jRvym1EERUB78k32/64JwxQ12KFKUumtJ1GK7HW3LFXx4wkE42+cX/FSRjEt
da1TALGAv23k17cgqXxQsv2/f+/ooJG7XmUvetPHhznkdcbGhvg6cV6jzWFuz9CW
2TgJxdVgRKjXuHfeh+tQb0qBtRv2fsutVsN453gMT32IGKYYZP/ksc4JMzvyZT1K
OHyyWI7CU23J8oyWrr+KPWxFCjYrzR+nL4kq18h6TuOlY1G2ySQbOL2gYmyWR932
WeJCjPrOVCnTrFdv9x9DitlrVyH02avtbaJY8M9eCQ12JeCpmkTbPuC1SdMMB7Lx
8WZLa8q0pzmr7sRq9o0xsgrOL2V0paPTITZhF68AFFMScErxKjOnLg873/AAx0WX
kUaHE3i8oks4fu9Rpq7XMOl0CQd1wc0gB5z1XqDfqu28UTB2UBx3HT7wx63+oRR8
chRgfWIHSuY3SiJf9WT6kTWNnbYv0BLV4GqBH1e5OnsSKQ4KFSeBLWM/oK2SCQlC
50IxjrNhFQlsU48XvgMVr8V0jZo4LfnnHPM5o6xc+Agij3k+G/uN9edYj/8ioMof
lrU3yJ4WH6lNSaWZO+R3SIFrN+IsM3ybvGyoIL723VPd5j46zUfU+9NZRPFLEiFi
3UFUjIqMn/LFVTuBA8OaV3rHz0ADi49OLFf2La2o3VTI8rnzpGJGbqnbkeKCVwe/
W2BicqKyRJ4YtrIha6She520704oT0U8cYfiiQfjcX3aQBCIOk2itCbB5OWPhF9O
k1KVhXUFJtjPfu4w5Czz6oPXiVOkhbSohUmxNhC8K7th9S2VKqu/bCGBQpyJuHk7
WXoR2CjDxWnYil/1QBbtXPl4EJfVrHYGKvQZ0SkkIJUymIzcEHsHzMmVM7IfbVOr
96lTmagGCB+6jlpWkoma2hULTDXOUN22mvi2Fy/3kX7RalQn3l1VLZ/FLV7mSoLy
2ok+PU/fEA9JzTgEHXnSvAJ+BKVVie9TkEIERc2B7+6Qo51zuOoGRsKvRlFK28vK
Vo6deVA3ghSmzBPjOFtkDtstUsezsDmAra4cuEE05doB6Tv5W9+qsy2MufEyOfsH
5Ek/kN/NI5m/A9HGeY4p8fuekYcXUYAorwnUQMB4IXxYmBnJdLfXuZKX+zcPabuk
Gn7MGm/uG6sRH87YgXvJkSF7jkj/OggvFKOAraWulU19j17DqZI1uWqHnz4XaEBx
RimWgmAUc3WU6yHeFLK+pj4iK9vcMRWBE/nOv48FQKjKUUfiAM1PfEDImQypBRFW
580o4TjuqwUVTgEFZCzDGRzTBjTMd5PalfYhOO0KulMwLR1HO7OLxuq0s8cRtj9W
fEl5FLokMBEuLBEu76fDvZqvT2BHiKgkaxglAXm2/LxzUXtPALjufg8td0aJ6gAK
GOQ+rB1fzOv1hUBhSbyzCuYWO52kqgHsnIkW93BSoXSsUoBrObc7cCtfRdKFasMp
Q9t8J8WNm4A+Jey58NkTmB7Uyih/vMldA4wVhVp/1r9U1t8NqANe+jnndlzocaMb
ldxVlRSIH7oQPuyx1mNsXnU5aOt4F93sHk/6i8ga6jFyLCdFmsDuFJ4pyPR5Tcl4
YjAvM1iznW7itY7iUgzkdjF8uxkoF7keqTMh0nqgDylgttPVVQk6CTsgCv9pJfnn
Ij7j6B/cfArNquAavQvrzUNmzLODVK6ccWT1twzDNpiPgHpWLxVBNqvazysquwZ5
9+O72Srj4t2wYaIFuRA6OCY3b2o7QrmEFu6xAQbUIUyWw1PI7v9tPb/aoRFhLuci
8Z71DwaNifAw7p3ARCuO+qBwili8GTgsvWqGWPE/6EMtEHxATHXG935/v3RAMta2
brE9bmpCOFsyBTzLxV24Nqpb5mJWL/ePTSszA7DJvfMqZZb5tS1GyAIH6esj+y6x
NmbH6qNwt6TMQfEssj+JxhePshFiZol77jQ5CPKogblopI3mj5qurnYR/Q7BiKS7
WpZazWqtFaELIl1Zo9bcTeE23AySFWiFj1poS5Un40FJCt82TXZafaYFvq3Fx908
6UkKLDBF2h44ZjhAh1fdNbJk4j2gpCpHfZCTLH6I8Q+eHnPqG3mubczaII+Ma23c
AWOIT9tOm4HE/bYRzSNriU1DQaRN05aUa/ixG8Yi9S5aqwqS0S4vd95MrOBqLP1U
lXWXwN1W8+gjJacocsacFOIwtOaOSJ+wpvrHmr3TXKgKEOhPznkKUTHdOlKCcP30
+/lIASnLePF/4PleabXlwh5geEUmhGLBoTEcGlo2Uhs0SLHN0HWv7ZXQ7KdBtQwk
UjMwk+sM9DJq4UChMuPFNGpLJgMTTZtARbcl1iyPaw0ZEtxShXa23XXkCHh0cy0i
U2UGJdQpRvG8xy+STfRq8locZabJdceFpGdX90nKt/cqH+z7PCzcES/ERgsUgcAe
OTaPXNv6uOVowurkA5uenCcmkrXChXpyRs1Td52EE4MGnmYaz4/kHEVOBj59ZmAA
4MOIZD9epb4J6WjSUbPCQej2dPr0lMdbKJeGBLfnnYHo/dsoq7O4ZpCcThZ6hBVN
TWON9uVSuYb1FUOz8JXISR0iF9tAqgscoE/X6kRHRwt8Q8CsKrayjwBw8dW3cf23
gDRSybcIi1wJ1KiaixV8toDdhnptC1IKBLsADney8pQjsCKT7VI7swQR7RTzUxAl
53Ct70rvGkaJj4kvyLBfB/joTbjtFi0W8L3zQPoZ74QYUUqxbILZBdY9iD7DQH11
TprMhsyrH9YTqqrqE7qQqiNAWF/0Bd7kBi+zP53MqiUpggZBgiPSi7roYTFBtSuJ
pG58sAvFADk65cG/j024fb5UTJb0l/gzPB7Cyw+hhJMmeWLEIFlAdlRMOPTwUwhO
0UCO7IEl2GSd0oVOsD7vcNfOjSFxziUvhEedfZtstSOROPUnHC50MQ/2sKvChukv
WTm4+kEPjBbTkvZQav6V103LrQmyS3+nTpWr9PhpQAnytSH7wNsw/qbfyGY5VyRn
AdCTTeAFCYg+53P9Mkor/rOb6sOWv6rgxBfbXJBKJ/lMQ1l6kSas+tbfChICqtSA
D20egnP59PJnMiyr80Kr/OEE1MVgcKxo1wEGpQQPWCvn1U2fggsmZV75uc4iK2RP
V4NRHlG81mqcAvUOeN+kJ6L3dzXVSZ7QDhzPflfR1wcZ10Sd3SJf+c7HWz5mNW7f
ygKyMFLDE4C58KHOxmoaBhIiU08uWkiZ8bz/M7ohIYhBR7WwLqKnwl0U0KXK6qOv
mhRzW6ttKnR6/7ypPBlhayTUeaqneEH7LpMul6ciu358acz1KUoB9PInc81Z9exn
KvRPso1bDYZlkZrYZkR1w69yhtSVXhCvuHVObufptJdYahbUuTx+gdrdaSbiawpZ
1mXahE8XxowyDRh/BLghW/N4LNRiyCb/uAA7vgDNYiJip7HmnRu7M5d2kYZYQc0q
ubFDTlijb8ZnXHXQNQa2Ol39Eu2SOQViy39grJxKq4swPxOp7rOWZ7aRaFJ1xE63
5dJmXX0dZVi5M0hyJwWWGbJPSa20sek2sv2urPdh229YRPtevQbE5C5P+1dsOF60
G7JoJyQ0eKXwRfohFa9VO99K30XsThQ14bAqD7Frb5i8MS9JjT5YGOeo+UvFXbaZ
W0Vn0/vfROL4uM0lQTvSrEQcyh3o6MVBRLOHux6hfJPxZAT+L4wGiOlR4bEiwa4s
n6wSXxUEOoQ3g7MywiQAtRxCw0kkOrjUbgmLnLyjDTLgGtz8LgIEVu+nFgfRuu9v
PzZU64iyLR973j/FmOCYyWKRYTh5ke/EemZpZTaxn8NjXLCJ+mGbPNCRdWs3JPy5
nFM/tAwXPkFoFNVaTFwSjrfhMCYOz1jyRBYEG6nxIKt3cyh9PgNUucieaMbzhq9P
XztW8A8FsTECAh6jG2gdoo489dFUao0KSMXiSmGNXyL4N43eFyuWifv0D7PFH4t2
bxVPfXAduz8V4Ul5zuxkRQ9iqwujR1TiFtOrwr2kMosrugLy5lEweMtzxl5TwFNm
n+i1EDeCBC8R5ZyfHddk3Mc/kaiN++Ei36R/q9TGA2xvg9TOuhtA+UTjRmGbD5H9
jhAobc+iM2BUyD6razpB2rFQhuMNXN0iiQdCqdEtmPmYug+GZ0vQcRMb49hLBndg
hG4Inx4MwXjc6On562Hj7r8HfX1RY/W4/kfhd70XzbRKLoHSq0seSP+A9V2UOOER
iV/X4HPk/wkHng997fBj8BEO5aOEaxB94D4nZQ0lCgrPZuhY5EEeiDK4FyM3TXci
rI59r8ZGLdot2RLiz92wiusuqWWT60Yvc1v2kgeStUvPpjDMrwmQxTD3eziSeuCZ
Ro2nJ8a4Ki2UVpUahp5uKmbhltWJH4qrukd8/b9fGKxVGLAT5Z4l04ARgsxh0Lpy
LyKgwWadEBn+231kW7EZDnLyEfY3fhsdE3MrBdBgAOaLz+QfcPojjNP8CQqTENxd
9EFdl6zOBgMbWkOxx4lz7utNgclYJ6eqyGWTdIRfnM9e35QLtcyS6+T7Ch4tBHdb
sL3IphlZe5KHgX6Q9E8gAcoj2f8nJTd6l5XL4x8YXdYsQGiO2pE9Bibd+FkJCbd6
Eio3aO7U/XwVKt9MSqWNZe4hacTkEJUluGRBSDiNExK7aUMCHrY7O+H+JFHp0sZ2
Xoz+h/0RFs7uQAtt1zqMBDxFaoTiL5jhmreRPWEj/pvZNHoAjd3R3W06fsGT9G0j
1UOliEMNgzQ0t0cwcDkwshUCNEYakL7LFR4cXPAQJ2ckqB7lgAEInoW6g7mXK9hT
OyILtGntNsdsgZ6o/ki56sSQpkuYsBHS6c5tos7sYUk06bKAkHMpsR/gL0y7jfn5
Ql0mPx5ylh2Zri1n1phmyQpTaViMMxOuufCRxYTgR2HaeUd2A2dht3SyHEHzw9ZZ
GKXEjh4VRXG31i+1u78b/Yc/R1K3UHVYncbuh4g0pW0FgTV/OiA5ghnPu3R+pFuR
NFZypK1ElT+SSkY4u2Oqi6zEPYDB+FUaamSgMsFuWLeq0tR6h+kNvnP19ZkQLjLh
kGbphhIbdfkUEuLP5HzIgnW32lEgjSgoANC7F4tnI4ov4DcQX2DNxJZxFD3nGmuS
VVEawv5+pLOwKAnZjv4UkB4fZ1wqG3TzHlf+6XNqFDfqEVrqXFXHECb0eWfvFOKn
E4tO5h6YVsAcc5x3tZAl1LChWOG1gqELS/3J6ylq32cYWNKQE7wdCW/dTGoMkXtL
fl1HJZuNbE1JI1mP6I/xlK2D9u7Ofqd9vdIsT9tsR4dlAKiNIb0pRmR6ze8S33Ag
vNLwPBba8uumKraF6FVqzyeAunA8YfDtnxUX4XIf/CR3WGqR3eFrWZZaO2bxbbQR
Jq0eDUzMvRCuzQ5h1wnzNT7i7+qKMdRX780/PS3wVHXs0TZDTfBYOjOsrvJjN8sW
L13t4ny/IXWNIeGPO8+MbPhyr8nwlPgg0ETH7i4riQH6gAZhHkOzhVMOeEU/94Qp
nmLSEGazzQb7nauAk8BlA8CxXUYKWFYmHgEiwFh6oRQvnmr5y/7dap1LuL/946+0
asQCVaxVBaIBD+mt8zcBjrJGJsJ0YrmFpzUlblHqT3OR3B560dXrBvHsMkLBvKyE
FbEM68VnmFZl4LdSsUqmEVjvzIjK+TUZXPzU/EkkOvJ0eTpKwYvcIXdJXLXB5hF+
yFPF2ng/a0m8xWO3N/OGRwXC0eoztPa53ihqpPWoxy1iCHIqYWUIb1lr+CCNCEdt
JvoYrysTvvLud1D0/YoRdkV38zn5SC9nhXh27Eqq4q7E6ILQ3nYesrBPdb35aaaf
mK41IdhgyV4BQ+oHzrRH5DYtzFOZ/AZo0trsnV7gAc3Y+asEtUl3nC2AJEIK2sw4
GGB9tXuDBShWZyqhdggTg+hsFcRj4wbpSonO0eNr3r1VlsjXembr95Y9bIGatJDj
9uknk12lBUWG4BUYr9b1gQ8Lohe3fIAd+ohVUtSG8sfNlRZec4uIX2yQBSD82El6
sEdwZd4APAlf9c2eoJybgmlufnMVxK+01haQlp7Rrg9clZ73ytLaCjlrz8K6srtp
Hci1isXK2XmdvC0Q975yHzslkxm1CQ2gIqSjdrBsMMksAHTIwLoAxfDnWh1hzO+t
xg9INCEujR7JfOSI17DBPEBXUYxiAshoXrpa4E5T3thCgnFC1mR0A1WkUGB+keMH
BxUv6JNzjJDP2kKYr70ieaFE04HEY4nIzC3sYvtRjCEpP1I7teHMZ2omX/fyaT7S
hgv627Kj+rb1vwr7cnyhNHUwu+vhkp7shxmmMidhlMROfLJrP++lfUxTa2rQCVnp
znCmeYT/jwcuLiy79AJNwcqwRSmVqmaVG27NBOrY2eo5wdkq00cy0K71jaWIukGS
r0XCDb0wt0GQtWUpCUPs0MvTqAZYbwOsxL2WMWgunuFtDG0fk4v6gY5j1caagspq
C68SKMJxMX3ctGdRoMOkdz0MRbJKJBtdxTaE0iBpfz+qdMP+RgAoh1yWs1z3zTSP
GlG7HwzNaO7FWjZPQLX+wmoSYvhNSZUon+nCqaAhBmTrWnmUeodYlkivIHS7WCL8
Sdv/Lbb0IRD6kg3vioVZFICWB8vMa+/mi1u/QQWYagP0XO3HJ9ed0g44AuezfZEe
udw1jqfoFt5Mbc3XB7IvZR/2BnpSfmj+sIWSZVRgDSPYkC51l69WJSaJeBM5Jmws
DR+YqMl+1LgA/g5skTOiw4Lt1NChhH3gA7QyucGtcOzIWf8s5voVpBpgZJPXFdOu
nVsCqB6zpSWPdZPwsXQ994dSzn5PrVACZFxdm1gSmbFX0Fw0qicplaLnlqrUdHG0
nJ6xg0NfKjEByh2ESliapQ9agFJHNnworDquqzAE19FP3p/e1/pesbUbx1hPDU6S
AR1hB1rAad/bRRW2VOwyaWOSGgCN0ARINzfPvj1SuFZOWhmoSvE3kXvWTAiTk4sM
T6Ql2WzQNQjboQkPUUdm8CgQt03cCtvFKpdQkCC4FhDDfLZw05qIu9r5KBbuoQe+
gLiFb2PweAdr2IaCBUwgp3QOToHqaoMaKwy+xvSbbLV48yERh9RUfXyybzNC++74
9xOxvGBfh2QbhGdbh/pLxwV1QHhRYuilio5NyLwa+aonK83YndRuPPNu3kxfCguA
nEmG53RZ7g3eTOjFKUlX10kEQtCNfbsU3NkgSZkC8IaFjioDIn93PdmwRZjRuB4z
R+P0NBCltC7DxPXrSJoGt8fHS6x1FKTXt6zEZDy6M0nfOuSHwiMxPmi/bgeyXA/V
PcVYUi/1fO7YK7CBFnAca570jGGZpqWuLxAPG0y9LkfEsVSfebo2az9CO8hOCa5x
viNUqdF+1AiyMmH7xsWNlW1kr4JWkgdr2PY/GEKEO6TJM1PQD9heMTRdfgAMDDUF
AiKJH0gDP2bHmqazq6cOBiPS09tv6KAD3J4YO5O834oDvbAQwQRKewTR1TaUWLRY
p5W4DAU+nAP9GCGCQWMrBLE8iNrFXeHz9WMmUf3Q5EbD6ZCp+X0ZGwMnKLTvwjGT
DOau5eboGQBSYpFHFbQNe1ZvgZoX9U4Oub+0d9Vvsz4jdbyIqxD5oCxmw/N6q2S6
pXo83/j7Nt7VbN8ixYl4/4hNfeO9Jpli6636+ati7KQfbjc9/kqh89ifGb7LUVSD
ZwM7Y4o2bV5cPLw+rFlTI2e60sa/zNkfX+po3zHXv4e1OZoBfivQSXsNHiArlUZ8
x2zn8fNsuTkgopeLyZwb5JUm0uRMuYO8oCuRonRJbaXKMKmO46fUzh2dfwWzSPlD
VKIF18gMJIBvDDpGxDCzEbGXpuUapiQAboqcSLnKqV1OIqQZ75H+HS/wKYxn6rrS
dt8TG2Sah+Q7cT/2/cqUHrVTcViWrKGaNJUvPe3q/J29+p+G4q0lvZK3SCT4O9ob
0cy+xzISpX5wHLwkMusT61lU9u55dYK1gWRAIEgzQjnwBej1vGzCTGkSVb94Z/Jt
/JzIFiklPFW35jBMY5yuNV+IRottVL5EUQW1F7P0DJ3OcKr34ZfmB702IZia6muP
/ynqGjsOlkf7o+CZPf7zid2Y7tgQbTFcW5H/zP2fLmj0EtcE0kZwRP+cJki3bWLs
HmJY0zetcrGjQVhPwFAePHyNaYMyBe2TFzJwOvL0DVJWVJiuZTN3U5wocI2cMyfp
75dxBOV2UP+Yktsq0EuVh78fKNUqxVzcP/OcIEuhepSm5HLbT07O7DiJx/rD0DDM
PPdaV850QYGpKtxQIKOmkhisJrk4MsILoRVrhn3Te8YcgdTsvy4l/KDY2MAsP7NB
Zbw5208Joal5a6dOTAX81qvDjuKKf4pyXrBYWRugCi/0yv1buPmtwae/87eMteZP
/5OYQxsejwSLbdGrZHsEx1oT96VjcIPOW/In7sOfKdPCso+j8HAQL/NdlmDr2O9K
RPwOYH20/jlY7aPe5Ez28NMhd2C4sZT3eJsdfnQ+n4IDJqWhvD+OQhWgCf1TMc0m
XwzBKYFMOwYpiex/3W5TNMQpNzsMBnCDssyo0+Bd01VIFa4bvwQVtabtpB50E0GL
nu4x2uOKaWCO6qKgy11ulJiJcQoW+Plkv8fNNxuyvE0LGDSVBJ0qJaxhJU5noznN
EYmrFn5fS5pDZ4j1R9dEeiX3kvtC0rv5uvyaOXy8qd8mSxSAlMNjw2xNrVL1NzhL
veVYqe6NoyOGDaj09IWSuYyXRZjR60Ioa4wClgu6hrgk3RDxnx+54nt2htBRFZ3m
SUqjFIPTic6uxZlIufYcgA8lw/emeRpcBQSQMBTutpg6qGrhtwaxTDrtBFb4dsNH
4fX2tcxlYp/bDydVsJlC1dfofXw+f2sW26Ve7F/kRY+YUC81HNXKGNNMIxkWHphX
lm3Ox33zTH/qy5AgrJjySa85tCgHhCc7KO/pHrYrC7/wXx9cSRs54NpwOlDFaM2H
aejQPni14rvaqzz1BoQith1w4wnkpuhvsX5bGYt6NsF6zp7bdJ3PgJ+pRKPc7GNY
UfosMY4GadLrgqsJ7QHP74vhrpof00hEoVet1Z2vn0nksJwegFkiB17u5c8g4Fkb
/kE48j8cQXElW435t/ORgxNS9qkXWMJjtN0owid9Eq1vc7iXXhk2HqZGZdPWAJnC
ls2J0DJhKDwKvfNBMoN2WyopnFkTkQ3X5wZ68zbU358/OP2ygefZatKs/I6Cr4a/
hfAOxpLztr57YYAF8NaKW7SzlRBPJHvhLzFdrR38PFzi0JxyvGfr3rYHZH3Tcjy/
cWowUlP4z3aoCFqlw17fZvfQd4xgtCQxOSp+VPzFCSLmkAb92iIfMZkuTJGIj3jK
DAI7VsFmA9TMiDUkLHuDZpeoCC3HMxESTF7yzOZU8b4wD+5Dw6xmfNsuMdf97aN+
lK5R0oFe7TkKUf3EBHiCrr7DC/SnjSzOwtRTr65A3XRz5zFqHOfCvYVwmpCs04ai
0LaIxZfQsz1l42vLwn5Qtq3B1zK+kWoaYx8zLapkXUwPzVr1x7xWkNXlphR4zeSd
TwJngn6dA15JC6bWuL+FeRxjavonRKhzgh79B3J2kvhRu5yyg0a7ZnIEX2iSJTff
AqTcs9l7r3+9F7g1vVAiftlDHvfT4B8rTEaRXjHRVKrs600iYMP2Re1czLM5FpVE
SANMV96vrQd2jl5gOrqKnujRn3Rw40HEpNhpUBmSlAiw2PKTUPQGRSejSF8h2iJn
wGVLcBl5W5iHJS3diLyyfhe2/vKG4FpC4EPyLo+i7YEtpwC1eq2gHP3cVjZbHZSO
JlZ+DEfq4kIJvhHGF1v3MBpPG67tr+Zwb+/PqT4xbRdLI49gRWWUJz8MkzOdAt7C
sYL6ZBidC/Bj+JgcO9VB7Gi1Yg8VRiQvXMM8ZSA3ztOs3VXG9cyuxJ7BCjYqOSsp
bYeW0xpOgVj/35+ex4x0xWvAcVKoypuS2ssMKJjRuhzIzlbQS/IAHk7fyXnVOpxq
2Pk0hxQgDsVUXH5FKWf3BJEAZFLIR9T7ERUA6oEX0Z84AVafjO0MW68lyGIvXNzt
AYiwRFjlY/yiaWWufm2ndQx4565sZNc2VzTl1rRh+NhP5nnWBL0pc4QjGnp0rAMY
UVKbn7JxWp+Q1sXx3TBZvcTSrObxslA1Hcr6Qa8uw88xpIMZGh4lvByVD1Z2tOas
dqSZz/6G2beBmX1TEwqjxoEO5quRNFDlSCRl73P2eYrq3ubL68FWjWKoDmaTfvXt
u8vM+uZRCfhCDGiZDd02HhFCA0fTvl5HceSNfGCLRkWz/41nNpfbnU6WRtHI4K+w
RdqmBe0SvaadF6zz9doGFkYSetljhXif8xBQk5nhamxCHc1V2JfffEMlCnXaqQbL
OnixdgyXOU5etkMWdfDUKWY2SKMXWruxozKlZoeodidaPb6bnZTDL6iuU86Di15p
pvxTk5AOC2wd3oooTujHolY0Q9FUgKb0fBtop1BmdvCZdzsutBVNyWe2puiUpyST
fLyuyzTkdDA4LRc92Ns3Y/yu+gHuv1LXiP5jNdfi7bY8HrXkexQCdwq8+gkimVGn
5cvwZg1hUS+bgKwr4lOO7AGfdSWvJ10DZvn0NSiNIfWKgGm/fg5u7NNiOADCxBXB
KMT+/ViuNP7VovhSbUFblhReuQxGUSHb4fRGCTOgP65rHZkzObapdCz45F5j1DV1
jW8wV7YmXgw2TxB7BliXPeKE8o8zgnQqNjUYBuE76XE/X6PheRP8Xsls7/2nvjKr
ufc+1xoJIhDGep87uZaLAPyqzQKsZ5cW5+vOpX6uiAWjq+kDQywQeTIpJIXEODXd
oTJxS+ntdEbwQb65ImbPBfIxgjJ1pnfvp2oZLwopNKzXVRXI+TvFwCVTUsWyNZi6
c0+tU5fvrHFKo2MdUotMaQAZmF6iugLD5wWohggKuqX5zZCwuarhseYopXR8d36E
V8EnFHmoZpLIJn3xCJ9kIV/Gv6L97DVD6+k2dos7xkvsCPzOPWPgvJsqf1S5X/cE
ij64j7TUliM+HwCmYRTuS+w89GlzquAgBx4brtQ9TBzW7wJf9FUePiapQ/eHrwAj
p5JeRx5ldjJHE1m/b1kBXwt5FEUJaRPpmvg6RtSecd3TfXhP0AiAqfyLOxjpID0R
3RG4VmHobiXjIViBffJnSn6f0qRW121+l3YXDUSVS0gSE2J8cTosyd1SWH5eC2JU
UWTTNwSLWhT+Os23m5nr/wNXO1KCeVcS4a9nKDbe9pbgqzB6snO5RH+sj3Aoi7P8
B85EpIbz7Otsc2MKfFqmgYhNDtzmB0rn51YHnmxHxARQH6FKFnscqmaHZTLDhiNN
nh3GBYu2Hsq8WPXQWYeEu56B0Z0cad+t/ZPfrbX6n8D/UC2qv1ZuALiw18Xle3sw
0Hh/lmj6jo/3i3RTFdfiZJ2ZgDh9yeolk9ENO7A//d17FOvuJowlx6loBdiATSxx
HhPDXnjThW6kttM/cYQ3/Qs7vKj/W4u0o/uHQFjGX/N/HyxIYoMZH5XXe/si+I9a
7XFRIqENB7QV7PsRqP6rrFrhbE2IUzuSXwAnRYFnsO4pCwbBEkByZ6JolSGwb9us
MsnhUypBlfXg0T1EFzkECFWf3+uGhrNQiPf80ZWu/wm52SEJAI3gHQu45QXP4OYF
vwkSnHn/lB8cLSJyjZ3XeCq5H/qpBYte5sBPWoQ4ZmETGG5H0RR8N7VWi+2aFiUM
pW7KC1k4ic4WSn5EXJ8H2/G4r0v1xL12z1abbViR3Y32PW7MbDKVxPNy9Lu693RB
mnCMDhvRO0xYn1ugbMy0OQNcXgVHadprTIN906cRJhBTo9YmHhEph+6hta9H1eIR
ZWfxAF8HpA+SXvmvojcmBqu+lr6OXAcijuaJVxkQ4XdF6s3aRoBRrll/reYPWsoo
InAsVLKNl1uoIuNQTft67O/jPg/29JKNKWvvQngd6YaUf2tsumU8fl3XzwjwwW8U
hspiczcgnIhPLfgvxM6t2/9YsFzD9Sp0hLPljqKaYvQTuzV+DaWV5GYtTZL+YwK4
8oGRPXHLBw3qEBVDUY3el7p33XRhezxgGy8Lo1Jm4G+2vrbHHjSBhP9m8PMZlLVg
tMFCYLbFrwdC48sf7KieZ1MucZI/sJEXIkytNJZINYWsKfj2y5DxlGiQ9dsoqObY
jqU0ByyF+2sczNQR9kRF+7SoKVVDfl0vyBkJQRYbHcA2LPsyazFrj32JntRaZTGd
nqX5MyOlT4+HMu+UlOnSp8ve8SGKs4Las+R0KUxBLnoNdgfmc6KFkCggmSHrgw8D
jKMckCq52NgAgYqjUlg/UDm886DoGvK6jXSJbGMloYaUoXl/ojf0zK/++wzZxEC0
RQOji60R3jCiYSJmYpcCfQsSPv0w+W0GMbGI5x11mMrv3h7VipU3qG8IM610THof
r++ZjF++ucJOw4zVU+5TtrSLD6bPWu1aIjJFx3XL/gQX6GpndWKciEPvZOvlA54g
xq6SFNljfMARXb4xOHEkI+nifalR2horWmpW+neaw/qQoJ3pzbkpAQrwlM9xICM0
FCijZq3/luwRHgrQdxBTTHXpOZR14n7rOR3KSBo5s3phF4YCiYCM1giD6L7tFdqO
7Gkxf26Eoh1fWy03lPl7xdr5zb9xkVH2oM7l7kB5sT8ESHPALhhKHPI97+FZpE/Y
3XwtDy0SHKXvfmrMUfpyFxsLX+YvGfg4nrA9KMOXtMIgGSm53K2T/43b8iczPVxI
svaKCLPIgDWqwKQk5zhFH1cc6NR6WpMSrbx6j0X/Q1DDSQiDDANKKwzRqyFi2VY0
xZvzG+dW32W0bTXTCE1Nfaork7mrAAHHv5RG7Vs3ljGIfMt7OQMFeKNyAXwegSli
471fFohm4SKL6WdscVG5KOj5pn9HUI4WeoUF0HhZb0uNIqdvPjjagHTFjHVxYJ39
BcsIDKKRKPJLriClkd7TMr8bfl8kLuxHfzIDnzK7+SxjWNYiQeQxhmV4/RJkXm/9
KHC6VxgrVd1WGqzroIcxmW6VEnrpayCk6sdfFh7cshvUuSgkMh+vX0u9ozoDluTr
BfPv8b8bzDrZ4yQ/VnfBBHnmDEvAHET19sZw9JLSD155ePycKu9zb9Ik6ZWwkeHo
SwUL8JHInelmHPdWdXIVd90lQaRxg2M5wsa0M0zmF984U6Bg3kjWnF00YLZ5Zhk/
Fgsc2b2+fwejtTdaGN7ENhDYZTbdeJa9NW+N/iChm5E0W38ZDMXMj4hX+VfHYU2A
HU6h1qbmp7v6Mx00bxKfdca/+aNdQ/EMH8CnWUXmnoxf3oAcisK9mr/NUhHYogIi
bKP2qmz9J/NVNfs6ZkJDNgzss8kJYz1YzV7t6MBYjmyob5So3bEUkyMDz5kqpwOC
Bdepi9gJIL+GPK4NdptlSj3IKOMJKFlfu2jrD3m6dITh6Uhn8MvrHUwgPSSgi7Mt
1A5x9uioU9LG0jLy3a8dLzff/a1GXZqfX/gVjTDcsfyspAEkNnA8yvXgNSFTLv/j
A2K7GDTol4DizvI3cd96FST4wMK9edYKqPO4LXcpuN82etBZO2UYhks0fXIlzkTf
JGXAoRTO5ktvQtdFpTDXqrviiIAdGk8+761Uhu8TD2D96Awk178OhbA7dyGtILF1
Jsdg2kk0wUBfJQv4mmUvzlmVYYD4vt920AzMWPLuRKvR9oY7BnMPodWmvbj99rjt
2ODUS8EYe47DWkfOo8DyYve3I+Ikvt4JyeEZXWUf6X+szHkZp0yrvCSqLPENFoPw
EVKxwZ230GYe66BRWXxNe0hzMdxKhOGhBW0v/Vf9bn9btLsDVjQEm7mAdi2zX3B7
s4vt4IPSnmafw6M6xGohaS5bv3w52nTn3EVeaV21HPek/EQE2d+bQS2zs8zWmBlL
DmxvELsluHc3dyuQGX0GE6p4XgZEvVegp/zttCfWhWt5fNGKS9Z14swF/+ojvqWf
RuuJcZkM5iR9MiLTg/k+9+DPsts6hn7ti87824J6uCP7jfcjZNKlQPfUTme4XpJc
GEvpS03aKmin76n42DyBHe+UPW3zvWKFr9bin200L5snKhVep5vLPlPPw+EHZur/
8n3QeBdfgkGdJxUADF25uAKTNpoDMPtvCoNewlufiH2iOGyFRrIJQ/Q2beJEQgw4
0QX0ilKl6eB2IblnPUy/FKcIt5tDeRO8wx0dCNLqoKNUA9V8ZSAYnFZH8+L4a8KR
YY/Xk2X9MZWbr1oPJoEnS/4hHjN7LG4jn5rE1yiehwvHj19b0RVFl0xLoMRdXipP
DXWeusQuDI1+1DVPHwstPXVrTEoQpI6KtQX8yVIWHbF5AQ9PqOuHW3Z9lu0+mEhC
M4JzbDvaijH0aGcjqimEggKsJwJgjQyfePQ/GtLPj10Kkaql5RgVVvoj6jFzZB7J
O+ou9jN92k2tNJSrDhxVo6d1yKZVZvyOoOJhtZqwm67bhrsrHBqdMVeOmtt1uYxL
4nFiQxGIhxZHwjUz0prPXZTkhCuAnxKJcMtN23uuu6EYp9su1iuWvD+KtT4Xix13
PDLasVXVubvVxkmYnKVnslE1MWMONt+39+DdkjuRl/0ucetesPNVyryRAMGbvfol
wM0+f4hl5+Y12ysKOlMJOeWE2ixOAKipvrG88omMGIdhqfCJPBnWo+kaOvMYBGap
UBwewkTbw5PjQ+pw4QrE0LmvHlNO9/KfRLVU+6Z4CKMz3DK19B/+P/Q2E7GdIo4Y
Rpjr5NJj0N8n3MGY6dXO96AK7tzQaTxRD9Hv+QdnHwET8fncNh2Em6cVr3xZr28J
S2Nvt7+uHuAyEjM+5c2iorkxWVahtvtUAtFM7zpJkLDP5ZQibrTGUc+xKITJ5V/k
l9GASBhd2jxFYQl69Vh/F9Go8tSBuXtm6/4WGStJZ63yt0UgK/zpGINBs9JUWpoF
4tfPZ5assjjg3AWCN3Znb8NAxH1dgf7lGVt307qL8A72gsUTtk1debcSZfRGUau2
LF3AZM0u8gtCF5tQcdpes9P3beQC9Fy8a+fANl1/TuB+nDW5Iw8BbFVEq5W+efB4
oCX4yPbZf2W+T3pdNHHGzPWRgQruqDGSvfIYcYCElC6HZ3/prkMrHUwkc00DRZNx
1Y0qbDk/7XIoSUNwQ0iXLjHsA91PtaZ84KCx0pfQLGN4Iay7d07eEjPhena9fBQT
eV4ZVz+l6WjpQnF9nn1DFxLzhmqXNiJNC8eCygQfUlQavse3rYRNkStOerGQBAxL
wfaSB7cA8NnRx6GF8DlF+jVAkQvmgrogh9NnEQBdbXU96DMJ1L2kqF+piU77amQR
2fH4BMPenLW4sEGbLWAQmj/nP2jPU7Lfpw7nxta1amjhO85r8aH7Oadk409qg8Rl
cS2hKuns3qV/zbzJlktmsaWKf55YAVU6rJ4d8hUx5VhAqWlml9Qi+XG2YN7ByxG6
iBtt2bKPFL9xU6EfvRgyxtZzB5Vhcy7O9Tt1mSB32KYoqUYYcT2zHLWVbEiNVZmc
LFZhQTJYnP9LIQuGu3aOjIknhK8SGwpMV0qq26aWXwU66I6pVuszqiXMzsLwaG/h
+R287Fw+m8/ykY4b3hQioKvx1x3aCwg4ZbBlCN+QJMKXs7WMIwXORCzKQEynJN6P
mrKwqBMTuUgqN+4SeN5uBKAwMQ6u3LdP9Q1Zp6fXtiXuG+w1oc8ty98IYYSV7pKr
XWKUWvrf2b/pAoru4ng/JeAlkWtUA/LgUsit16U23SFfVPRGo4z0mI7xi2wW8TGb
7C0OSFWqOceoXUXwQvd3TQKdjwYpZH048Eey16JOaoMYypnFfEZqsQXJxRozTIsU
XjCAj/obBNrD4V49e3fwQ1nSbzvPDWwZkkR0pObqErD5jWJnZAfTOrlk+lGzJtlq
UBGKel1TctCXuLmaejkKiZ3z2JFZxR7MgGzNFAFqKwrBvODBpk8nAB1oXUmNc/4M
YWvRW/NGeb+LwTvgzh6ODRrTi8+d3z4KI2BCJg1egDLNrRZBlk+r9SeV0bJl6Ey/
AUANLBpPJsuf6JoRkN5X4qIzTVGuNIcQQr3Ctju/IKeH9RwQzy4A6LKx3edByRMw
veaqCor/f4IWpcF55a7RQ2MEo8UYO/rdVzW6sb5HTZ7sbm+WHDhpuClWRPI5BP7o
f11s4+tF/Wx+GX6TnWc/2Xpp3cT2yv2ouO7rX4TOMNPdRIzBbM11DCLBNIPD1ZXY
mgwAbTjbyhTsE8o+AL/SMMgiXnKzWDH2OAmWdqSgwUqy8tvptw5VNZoDzB/ZuwPp
fuRBOqL39LyicYAo3cQeTxARdg6T1+D/m81sl8YdvPntG+DHItHfKsJ+5NYmOpNW
GYzppSyZzlVzQ8Olhi+JDm+KA7IbDdaLRD1AZDc2qAE+6dQPd320vB4KWS8NBoCI
4utZvP9Q/fsY1oBFwD2DHUB9MU81YCdcP2xKPF1vUcY7ikJzRZ/axOcd2uDU4BuT
0ggtbNWIbW/6D8SyETvQH0A8qKNSY8MfKZhBrib91qwEMjWk2QPd+VSOQPJ9xuiK
VHbXYXVwsJ3JPwGRHpsCmRQs3U81hJTTYCwLMKOtN8LXve+oQFROnNIOXsjYpPNN
ExLHccJ5yDP4ZH0WZBIUQp4xCwNh0WT9bHtyJXbd/BmK9vbHX6eP+1L3XTXLEXBk
NJ6xOh5uvGjejMKc7mUHg7r6SU9Yc8QTx0uaxzUUt7Ho12CQpYJvZod8kJIuSa28
2LfFB6qK03brOf68ZYU4YLqa2PcqFJ4tT1k6vnnUl+DIhCUfalEAi1mfbE9t2+Hm
aGP1TkF97cs96il/vUlOkYutWR1nAjqfB03vCvkysn2TYYVxikX9HHRSMDQDt1Jh
eVnVf2q1qawyF8HTXbcvq0X1qXG1pY9PZ90BsTtL4CeVaerFroHZFunWpPtyAb7F
ws+haID/TNl2m7ytBvaiI4yQ8LI+h4kwJ1fiGAh1TCrRuTlA27ceHOoLw9GuVaKl
lQgCT2FiofMP0rpGtdAyvpCQG/MgoTBp4PSFnfj7Nrh/guo1p4fvRW9Pnx0nbkjP
NW22EeIXvyz+FsJnFx+XS2kdt3X0M93Yix465/AzCJV7jSr5AflQKYFJLh4PC+je
vdVCvMbd3SSbG3ceyLQX6HmdvsEgPLLXA4iVWEUdA1iXBdQslQp4Ql/llglXYUBB
ewpixmVNzsfaiIpctGpqg+QZKScoY41vQfjkso93XimVMgEgRZAlcDdzp8n5Psah
DaaByReSn1QLnPsWeg+84Ry5mERVqMWByt6e3NZyAo/wXRfRil2I2HQWrQd0mlKT
FDtKQg0PNPCjNVrIE8x4dOEF/n7ov3lwXpNyzJOSjfxT2FDQJtvd3+eWsMIfmstd
GnWohY0rLMEKJ/zLl01ZFNeruR8wGsuXwXpCEyRztNRSiIp+/7i/PZvC5+n3pJye
gZJekFhCLr/nN8Yq0/4CUDzVG9T9l/5tlCZA9vwBTLAEZ/iwadLZ72TZB4h9RC/Z
/F02LfAW9q5uea5kzDXN4m1IUy0KPsoUmBXJ8G/qS2V1pysFwnUoTJb9i/teJG4R
r79geZRPu4F1fyX6KZDd3znQTVxkxw964di2z60evNvZjvSnhJ98USzq58LfoSf/
OwxyNrRXn9bFrbFrGPbTx6M0Zwz6kDDZKfT/yEgj0qkgpboVH1JO6eGtKLmPwgWm
TfpLaXfS2sbUb88VuQwRplLDlcPaYF4cmN1mGiegSh1imgpuJBMsJBClRvYNCJeE
5MwhYEjGlC0E1p9gTtQAuyVvi/OJeyR80OyvA+8U/Y+xWX3nIU+GAZiYPMDVDImH
kmjZs77LHN9qq9X+82ago9bl72XCvddWs+rIO5WUQLHW9JB5fPeb8i3blhCsAJpQ
Gqo5sUdVIj5KQCnJFV5qOe+j0+ETVhcl89KMzlJr0LPsexDIs0ohfptKd0yoyEcX
wauNdGoLgfyVAqa72ef+a6VOM6TcS9UL0xuZB6NgXDNJ9cYWmfmXwTxchehYSDqt
siBZCNq9MTuwS+/vGrin4VHTDYyAXHb3DAKImtyEcnELw+mZuSxsG+Gcyu6uqiha
7wzlESwmM3wgFcgT6GiPVR13YuJpxaFu7HYDcM4sUgLJKIBcpjiSU79ow/o0fBkO
o8eNxTubzBtAGiwI59cdqVslUzqQATHQO1i6q5lDLoAkQv4cdJ8Vmyirg5G0YFS4
93Jj9d28IvsUc6k927Zjqc2x7WihOcO/LWVsaLMrfuL0DhVmXhRC1NEHjFCd/PiW
FWVvFP+LwfCNfXZOMCWjuyOcMOLrzuPDkExx6LiUHX1wr+kZmz4ZKpRCWDu5Ig4Q
IEzYB3bSE8hQ6lW9ffxXURESF24PmSkgppSGST6bTuxCbw329yGytd0FvEI1x4N6
V9+Cr03IaVsKbwWxxC49AiyrgdK3sNT041uyjYng5o0Lp6AaQVKJ+UOwL8i+0MNz
Pn1aYSrreY3PFm9tKt2/sZlo0xMo7qAQA5rvd7oL7E8Om6U0Wgkl5YIHWggoyvzB
hyy790S5aNtJzT/MeSxng8qpKaX77nf0mEYdWrUjAUipxi9ZhBrFODkERY6wqkYg
O8kF2yovZGLlpDPi7WCDf9t27KRkXyAkC1OTZpYr1EbPIrWI6TxbXgpU1zz77Wru
rK/FTpR4ibKO9Ruwe5CqtyxD0xAEwylIRMAu3GkPZ/LOfNiTGZkSH9PVS+BhNeIL
S9aYp6PkG6cXn1gmnKhBNja3KNRjrCdHVP2yYqBWVWpk+/rrX5by/T+HWTm6pvOh
w5qi0RnLABjkoRgUTokAo0LW+gaK4cSVqhHPEAKqO1yvtCiBaypBAenPltOxENke
pNv+aZ9Wv5X6HvHTzxs9FktIXmilGxmOQXIFnjBfVZcfhF4VGGAJyQIX39nbCFKm
i62clp3aQq5v1N8dWbYUjX61rLiKrbOXs2RivNY4ME1d/OVwzq1OAMTYmDI1ZjJb
iyl72ANfOvMug+YXvv8eRrIo1UUCNRa3N87dwI0gGGkvrXeEka3CVKfpnW1hq40H
cVT4aLzIFoHRw6j7sVAW6pU6XGgBiP3qmRlkJOlPgXi9Qe90JLDpPx3jOm0PhJit
8PzG0ha+62R6BYcogvIud22LAM/rSqbqmVxyJvAykG24MhCwaTuiQdQ00hbKyzwa
vAcd/b1ZfrfVV9NzjQ+XpUTQsg0qw7VN1xJv4tn3W+UQVv2bGtrzRbl8ou9U640b
OaBBmGNXTRLwSG0qm3mfYYx3Hs/K/BBoWgSl+4TR/M9QOji2TiNozyOUQCSpNKhR
BgXxEf/MTfvxeBkgPF1/DOIcpvDDQjKBZDXK2rgNKT5xlGNkKdK/Py5zP7HW7cxd
i5W8esjmvOE8fqBgv2Fs5uJsHFfDsyPcaarO86fAsrSMPUO5K7Bd/tobgHRF5LBB
aUDwh1wchnXDWbHWbsB5YaONegDk+PbgEi9PmAS89lz32QrHzVHcsf4KdD01sss3
TuQQK7gwiALlgbwC/u2y4zC2Sbyqf9aNHTk4ovVEOx9vqGBzfOePUzYQYPG7n9AC
uTjh0HHjZp/KkqXNE7nXN/YvN+PbZ6IyXFepYwOlQD0CbjVO66/9yH/e+3dH2K2g
LnruM5DYJ2Hqd5vLN/b2v0RCL2ezVTshroJQuFouzWwr7Kpto3lJZUbrU/xt/Fry
v8RAsZXdeQagj1dTfmImkby2krzDkvNwjvtxl5x0uQKchIiiEhH53rQMIDkR+kiv
NBtp5o6RUGzKBcMN14+vSwgvtj+cDSNy4nStRiR0wgzGpjhmygh2z4tyKsIsfsF8
THAlvY0CcDf3ZOq5ltgIbQ8hK1U+nLe96xLmn7NtC2JsaaQYaxIKDJofcPvD1Lfl
G8NYJbPt8afsull/Knu1r8bZznk0MDot4umxTCQ87HTA+KBVMuZoDdr5x0m5RZoi
Lof6EGqKsRWlEcch1zPN6FvpsfH9hKFDG0canV1ka+Cu5hVttNlgfNusaj950WpU
ggJOLLmE+LpkvsoNbElBoMIa0dwdzfVb1YRdClD4bV9+of9pAPhWgY1fBj+LgoTI
lPABdseDoyOe/EgUTPc7neSDmnUNcp0OA/7U9fWpSfokTXxJN8MLMHJ087lInncB
+WAYCMJ9tUTCsQvWg6Maw8Ky/604s3jc8bzY/+S9A/TZ56lAPPvtKmJrhTaAsqsQ
DSlPgJYdckwu5d0rqqJ6+Dw6l4bmFPVj9qIbemM9Ybyvp0tkyMw3X3br12ixrOFL
Fvm+/T9zi/Ajr3LQt74OgsErL9Dq0xesiuQuMDug7sxxw9HNiIw2NNsL4OrMeBMA
qiKJtV2yz0hozyh95zd3C5UyMDTm4um77YJ/+s5RsfUQlMoL2MjzaVxtm0vtLa06
jFHnzUdcMEDyx6K7h3XEdNWgYEiUbHVSQLe6vJFlJzKQrK6KXjyh7XVMeO8IotHw
dETyD3DbQk1QSyEWTuMiZ4dhHELgN/zsg1645clhrC0nw/V+YK1HplY6mfE73eTZ
AsWvT/+droFY6RsBp4M6jSJidkLSBz13CgQYnlFEsx6fZymVhZNz/tQT0TWLol6s
jCdGTY0SL6rqxSjeMywesvMIGnvpIPFWRmb/2UIR1LCudIqDmF5RI+64aM709SEc
aawEAXXOm79te4948pS5RdmchnhkI1QQcsfaGdynW5j0ER3FysZHizDAKjC4cY0M
m/y4oRdKwvzmbx6sP0HlrR5N+WHRNdPNMubIPaw6gQgy75K8MNbJO4IyM5K4xZ3j
HlrxBimG7VBLkayBG+IZwDuQs7igPyy65iUg3jMRwywTbhdwhoXSmv5oBkEpFFQ6
uNjYT1+PbDV9V+FsxItimDPXkGUHEHPeSn7qAJDj1mRHw3Dw8m1RxICbASW5Vf5b
qovMN38HXe0EI/1K56pnasT1/ihQn6a3LKK7h2Oj4oyHm6cGl9No9JDOrUNH819t
ikOMjMtfRUHfoGAr9TONfSZUU9Hyu7A3Za7v0gU4TcDOh7QZRNgQbnRy5Qg4U9eS
98rv8SKshzS48J5RraBG518Tvbx0JXHp3xIFyVUSDVJLZvHpPKIcDjmfGSsW0MyR
/O8/1ecnOnrpp1R+FX82nYklS7h/MVWx9R098UnICqQowYq/b3vHGWsAMUdWHz6Z
vGlhgadx9IkQfx9uZ6eXpTdzz57C/58KnuHskOdPP9QYPo7EcR/H5xZVSzu0jBIU
SdblU7PwWSpZ3pbccn+BpjzW1MTpNnOKTiJ02q/FhbwiHD75b1bQoueI84agI7op
VMjYcvncXeZoq3tphiRbrdwZeHyL0Ac3GE9RtKqDfyocZUfetZFvwXrSjHc4DumG
WBnjv0QKQNIisSLv+3oFeZZR2uvOzHpNbg7fRaegV5Kyjb6FiCDiWgCRSkwyVIB1
FX9Fm4d85/Rcj63l6alc7rEM/EHnIOAfQVxFK5JWw1f7W+Pc/iKiMHkRxXkEzUpv
DssCHuNWFio66kzObGZ8Hbg/SwyNx9PwOFpOlP+dAG794T+40TAVTWeyNVIZMxd1
UefeYUD2XBtyIcskd68bJ7BiQcUuDBMPOSgwltKdPeXPQfKPlSARKK3bazyCOUSE
Rm/MQKEcbI0pryu7arVC7cGMTol9qdcIBbf4dWIDM04ncyRrVipx0tx63Bu3AkGG
ddEIzvfMGHRGGraimwUMzDNLdT44QD5Kp6M901mswPKCS8sv9JAGVfVv/83Q2gXM
YGINXP2f+FH+xcwvEy6zLW8xIzTK6msUH8x1iPIZBeUd8UJdpROFvMvxLjXGnwKe
zfPR2aQy8CLN5DrczKiQdsMDN4oCAKRTJOGk3EScB7Rkvo0rJZ2aPHavSCfgX45O
GAT18FzsB1kxLp2goFPK8g0NsQKJrbBWHT5apr7J51BOCMmqeqVZxf8BoA9f2M2Z
a7z+aEal9Npud4FbEyS9QEJchVO5i60EMmEW71eKeuU2NuOHD74EaR65xztbf9P9
rCb5i8dusDwTdNlrcE+YKJZ05prdc9I5tg/Ad8ouWlKsHcuQb5RVW64Y6MpoPO37
20uyl3iieyRIUiJzWWLERY1oN+QEtPrjqJjj2IJGTosVAuLvoILXtI0/kZWLyafg
H8R615twYQ9T9eRVWwuiCjNrNEB9b72L00ReqcstrcuXx+Dxkx3ydzGpC8GoTUS/
nxCDYUBKQvjF6HUtX5kZxCeRCujLcRUkqOI+AWorcRNOAOyUrBawAmd6f6MJELim
UPVPG0/ZAltcw8yt0jVVthPKESFzvxUA0cawEIRmUXacwZH1TguKppP28ITHhcDZ
4kQiWDDcVd3FVqyagNjR99nFIgA6ohMIK3qLVE9pfYN9yut9j6d7qrGG7BnZ9vgj
UPtYA/83o3i/dIp+oVw3wUvW4o4CAauwO6OBB/LWxLi+BR+gkCv63THO++Bm1rvH
F86/cKuZswyF/mxU8EGraKaNyEjVqQYgSM6zT6wGndOc8KvO02H0zceHtGisAfTk
7+CzIpxo7NI5ksIYPOI/WF90ixaXoz1kLVxPFNQmiVc7SuZkLiXvRx6iRLqZuO5R
rj/SxNKAKhTQZ/FW3RSR+qh6pR5rjsTRdslS/xxrJb/6sSUhPCUNnrHn4y4H9TLf
6pndrjwUXIWUkf0mhLEVbod75xrj7emKXxLSfeZv7vZ6L1P1vxGZGUozng+h2Xg4
Nh8UgigBkDaHGcKMLWYkShkoV8ZxakKqNpPEiHpYrD8eV4xXA8NxJ/CTwmdyRbFo
aMLCrvaY5mcXpDbgxYaWEtImoOOIqBSKuZszLnbLeC7avYwj4VUxXbDgpYT6I/ub
hisPRxeSAfKwOfgNKyr7C6zIq0DJXF2HR/Zo8OV8yqAFx0i7Vuy5u+ArsnxZOmC/
Xw/1LVqbB4vipsc25DO4SryUFv/BDFn9/KWgD0gwno8nLHCPc3C8mbsl6b0ZOvSx
e+7gLLsTchG6mP/XzSKe+IpOpR5vbwff/I8WfClQSHKtOmL4ZoxzNa7m5MC+NO+h
Q1pVb+dqj2dXLDu/SqhZ56pmrUxVYbfKSUSZ0LCJ1vBl8FRjUzCYE5z/pDmrgTt2
pPCtols3cPlt5KsSimMqtLWEijk+aFZN7w7+LgpRpfERwoOB9S8Ip/nDZ7KxtUHj
snaAN4PDzZxSpH9PcJ2oh8Prq5pbfclhd7K/QjZSB1Ux77myxH+oeGpGtGdTXA1C
psQtcam2Dn0giCm1HFnMhSEnsslmgvAR/LDmNQFe3h7XuWr5NZGZqDuPuJikW4hF
/D17OGVGxj2VpZMecdcx3XUH7KMi9libnsJkVsbeI6FnrwQkFtkO+Tg6LRL9eUi4
9EA+Bhy8O0CoXCbOMf+Q5cfiNyQX6Wg3iMgOlO4155XeuiStdkPvlqEZEI4f6C31
3HEGEnE10Z2yK1SLHik/xLJdfxThpCsOSEn6NDHRkY6yAUDqh0mlewFIghP4CwmU
Wkfv7tE/KSFK1o6q6Unv3eWysbVZ3un8ArcEAd+YnG/puDwPlqrXWVKHHoNGrOwu
xLjhLqozoMsosCDdw+UhdYY4snvd+qPdS7ThnFVqXPwPFGqcEfQM4+AlpmOZ492a
HIhHQWl/Y6OdckJIYSUHi12Kw4+J9RA9DneLiam/nAgDxwrihE5LnDTth52uX0ER
hBAYqj0pXrnPe+PSCdJAjMkUY/gV0BYr9zGB0BIJwdcmU1uqZg229B50o42NGeuk
Kc8VpPa0gafsvev0A4UuXVZuuTPCqhFqAqDPDyOrQLJ6QCAdVzrlOAlmXVqfgMwP
YrKaJfpwDNrsuyd7jslAZKQbn10WX7Tk0O32v8egKTaJLV7sJqAHm1Mb0on0oqJ2
FcFgnHj1+qcok4LnR6mC3Qi9Sdu+bctGboakYn3yPWyb1KjZOKuvWd1nk068qO+/
cRRY4liFQdzUdDt/X8xONNGMfAq8wNTLMKhAqeMoipb11L9aZ2PYjJvucXusQFuB
KSZzjfG0WsbzAk8QIwI8Kjih/kuuCkAI57AAW9JXcFnCexxidmAexH4s6UHQyqtO
2z+Y8xq6yiN4PjSe51vsMYORcmW3LqlGAx9/QrmoGk1hN6ddGRU4joIMjIUbPE+q
FVCo+BAldHu2JN9aw+fc69JtKtB5jIjqbTRss7iyvF953ecQUOh/d403rv+jjADy
31kRcYt7kiEEktsRCVIO6dstS1ZoNuSYkzYYB74mZsvn3VpUrOMcVbXpDbr3wj3n
D+tCAdu+bNVu1SA8ct5pmfNqk7fC6MxrB5BPEZm7w8EdWAkgaF710wvn+Tv1ko5R
Nj4thYsCmUCwSIoF/auZBxaPUW/Cl5f76PTQBHCPokQU4KEODfVNCcYE3L1x6XIP
btDR0QK4JH3GWY+fJ6zI13p7JKui/sGqvFcZ/PALOMUle7NsGo5BrM94+mbazJtI
UqmhlCmj4H2Bjg5mXQs9NRpGros5kSLalGgG6MouVvSUPJJHQNkKETclZZUXbfK9
ihpItFaJx6hT8AAaB6v2JiqBcM1mR9dah0HMhxpYnVkQWT2x+K90D6/6jo/VylQl
+d3wa1kg/HDn28oqGIu3l06NRFnuFlaiGnH2EayF4HNSv9k7V7TR7hhXyJidHuNm
ZA30awiDzbCysfYEW0jAM/4S/9SE3sNyLED0Erk9TJulcj502E9OrqB4ZTiJ4EXV
12qdlpX3zFOc4tSyZPSmteR51ECXxURnX0aGyBORLp7Ftv6l1RiMNW+upiwUcZfX
rG3axPmoIEXvl5yO5MSU7wga54a4sugUA5T+RkUhuyY4QeKIpFMa3mDJ9jR8lYqK
TPd2tH6xn8lboVl3/mIzIFpRgnkdWMVcPsIR0XblQIARXHoFQVoO5JvwIZ29EYwI
fvxeAylUxMesW3je5ycwxRJ+/kPwZmsEk95xTnaPJFCwOZ9ZhGjJJpCuP4KqBXDo
BgrgxiBjeD0iiezrP/O2rkeADVXazJJGuoz8lhr0t1rov6CbOs1FlN5mhCrU/yRS
+8ACSsuZB/M3T0U29J8u+W3fFe0Qc7I8ChCziXA6rmKfNbFJFsNQHt3yktFGdA4t
XqgeOgvl0aryo3uXRX7dPEKCnc12UPYC5eyOBlBxx8KEEaxblNXpk4/OyI3/hx5J
cXJUMNJFoVB3/55kmqVAzbE/NBL/Dgc2QbeOyflXNgkg20EXicbsMldMnB/xdcbA
ZBdpGPp9MdNDpHfGdmoDhCtH1dQCmItfZVqxjdLYhgxTHyzLMeq9KfBfQlapqPhA
NyD6EcBz50FpjJH6dOl0WD3nSkQDT33TiLVWHV/jazOF5BVOc30XJgnR2/sHVwit
bGQt5O1rJmxxc/waCFOkU2xBGQwMDBjRd6ck7PzhJ5f/n1y6KnQMx6a9+QhhRton
yVudYG/rYd6ZhMarMMQC+J7qAcvVrnc8OKrukhvFDrRPIlonhJY/PgFkBy03Ux1g
rYJUw9WciplJX1vSiqZf/V3uSjLkmI0WoJgRvnNKSkUti5gLhyynUJkMQuGD/+KQ
tuH/F+IyieYnqo/4xydwo46A14F+NG0q7vMkzNLotb83t6r7lSwlSF2nhwc0oxuZ
xyfvfTZ0tv/ZBJXSE2HkGdBKQCkGCQyfmVyeydBhc1bfNtjvxBaHTuo8ln0tgeGR
CfXvoOUbQC8zUxzxs4PsoQWqhw/rhyBuZ1Jvn7T0+KL9ZfRbaLYuzV46S8FilPhF
cs5ZmZ5VZ6dCx/Zg0/vPUYEHDhnXR6GqjnVDLARsMK+Vg2x+lBnkKKQtJR+5TWCE
7orIbgl/XqUSMPnC6w8moWExQImLgTfMBba2qM40j8kcEi3loOFp+ZBZH8zW3WOx
+kO0xkwUGtT7ef54vHqdz/qHBME0IIDaD5WH78GWd273KlbNv0eekp/Y5Hlx2Juv
Yf/soEwjDNp9bgx4Fc1avsIZIHI8nCGQZsRFO7tiPnGR/K73i8N0Tz2gsmfU7dBs
4p+YTBMX6ZBCb0q7mfKd13coOQi5ujnSckDO7kBVnDfDYLVPw+dTwAGj4Lhw6FFI
nMnDVdoVxVZYS53JuZDAUihglPQLVQlXUx7GP4lv/2jX9SI/Dv5HEBstbKWZ/+Hw
IBpd1iwMJAQDbZvjDuVjJsxt1QsreBNBOz3xdDmEvlEIyGOo5CVjX6UYOTeLYbAR
GfPRYySK6TASPxOhrfbaXsmzYlm5bOU9jPlyYYyXVdow91fuPQ0ooSFyhgOpEkm/
rY5PpRRJnAIVF9kJ9frvvLz4ZX+PKd3SfTNahMEWgMpp+u6jGbGOsBZnHbduC5EC
k7dOt3QQTJd28xr1anXb54DA5Yq+Fb0eukuGbeQFJ17pztxU3KljJvhAXzNHV43g
GCtSHgczRf52lDIu3ss5Ctaoilsuh7B4LCjTc7uNMPMgzck+QoBywKIdesuehh1+
fMjnqbBxdEj57nkikIy9WT//PdHAPnD8VekVwjCTA5h/rduBjAXkStBRbDzH6bS7
8XzvPPtx55RteOF9DSGs66foizve1XaehdhdVfWvWvFH+t0hkONfMj/b7T2hSCH+
ue7bf7occ9HuA+59il4YPACdp4n5XY6yJY5W94NvWKnhFv9FALAi4lqazhmNb4yU
7OHSwgJWmweEhslP+w0X/allRJNrUAgqwG0W/75OlQ46uVFI8RB6zSZrdE8ug6ox
7x+6KMiKg/xsxMQwMi1x2n/akbiFr3NY+MYR3JFwzyfnyWhCSlM+3N1VDJXMNnve
2qlbKdnbkjU4p8urtOyfCoJ+aZ1jhmrYb15mM5dG5qITfytl7CdgRrlths1Xn1DW
FV81jEDTSH5f0mv1P32K0htvwnvjQmXhafaz1bHdqn/fPodm/CXNs/GFXmA+1wvQ
TKIbLXOfIOFiyhUg/790uU3cr47KCYkNxoVMQ8k9Q5boHDYVAIKnpt1oMABq6MBI
kx0TBqjipdP5k12JnU2vMTN6M4aNxM0zY5Bm0j2QH2MYMEmfgBoLqAf1rb7+xPHf
P+1STRix2b75NwzDLdr2nL/lIJXI5HaWLJD4PTVIjbdJuwg4WSBF35atLcZkD4Cw
v0DQ5QTQxOyPRlwBBvDsXr5chrZ1wk4PoIW7G6acy5B/QN8DH/rl9961A6dTQ2EX
3sPvIkee+fJ/BghFnbyObJYsGR5aQX9MJMUsvkzdzswk7dLRqJiqLYDJi0b/79hG
nh2IdEWVSM1RO+/cDQrA92YoWM07Sbqfxw26dKu/7otk/CPiIke/35716SgbxttC
zlcIrqvQxmKb9TNHnqJ9WukFbCHYO/xxBGEJu+ae5Gi5tSarZd57qtutmt7/wryy
gq164v0TREQAi+i+t1NTz9WXRIOXOY9EI4VzywGz/Bcmx/bWtNi1tnqKRkEKREOG
1+3TH/E+d0A/cAhQ5+9ytBAKPUfNwMbwiJJ7g5+2fX8xNwYnt2Of2ZSjEJD/VaID
IYZbu+1R9luaWJzeAJrPXZlTbtpk1rrrAlrtI8mGrt+LZMwRBbCuwzqwB7ExVkpU
CSA+SR/ddx77Qe1X6zi4a2FqCA2XLNSNsKZGHld1lnB5VfmzW+m5Em7hvtFTARkl
MrSKMKFU93bRyo+C4qV+TZqrwqpyKI6IYaHE6aq5La13LkI2BRvzkqcV18lPqmzO
AAbovxH+HqV1n/ZSqjufRvJ1CAyCnuR20iYuOEhOcDqaWpsPRZ25qOpKPcAL6Hk+
Go2fLqFzNYvTIgZhAduzVapAURCKuapUNq2wtqG5iDyoqzXOpXC0uIhKsDVIhVx4
N1GdF72alhOQP1K6zQl8jRdmLmV5HLo1NRC+A6TRGTAVqE/5cOuaCgCthiXriRzq
8jK6BwH7jgKZWZGwVjjb+ADoL7ialxLaLEmDYoa+wAPLxoChv9nCVDBJbTk9gwjK
sSb6LyMcTNyYeOzNtndVFw4+1b/PUthvn9S0LxxaOkSG04ep5+pzXzd2Xj0DtlSW
t8mmXPqJyy0DctyWIu9QHsSVYSMoeWsj+UyZ8uWt4S834E2T4fCBsclM5qmqiZsA
P2DiuaY/3VksrgPU89mYGIbYWEubjjuEGh1sSEjoYNPjfCw+Sqk9Iq/MrTXV/W8m
hsJ4HAORLhtCQkSYbFrnu8LwE9ChYntQtdSXYE5Yfu/kUR6Eo6EnmfBjI61/xcHm
6ODHzMkKR0yGvoWUPUDgxSmo06lDffIuIxIx7MHNytl0tpxi2TbkSs7NiXplSUjz
MOAdkBi1IKRJFr2merF/07OtA0JbfrIpmCRFlztkmMvBDKwIvOWuQ1pJCrVaKggL
dSvUmrHrqZPO3uUjteWLTGLV97/LQWisuGIe0y1pkrUXDPg+w19y3iqtDNhc9BVo
/ZcDwQ7KHQi3DbwHZVD+hj9LO10nHeVZoFclGwx/JsBWgoQizHXBY0bIL3qiSGK3
9y/F131DPxZTayCleCzgu38e/wYCj/g9NZuRA+e0+EDiFo/UOuMJtswSdTuZrte/
Sk6B79sPJLgZsezdCzEq3FAw3GWke/6s0HMLv3VV5kbz2ZMYe52tZ6TimUGpg0GW
K4wZMKxl1B2ch94wZlFRhXR6C8Yq+cF0NG9NupHu8r3o/2hO2evvjDZOoQoKqpYs
+eOWt1tYtz4WzEJi1V9+TsxSZzKGZZfdP2bQfQngw2NGIc8s4BOb21tmegxjcrud
pF1tmbW5BQ1hfp0ZOI/4iWlwh3iYjn/HIx0YqSYrh4R6DffL5hs5sCWFVmUZAg9n
TtO6PyfPsxJVYZspkFmSrGe1gFgKz2fPAgw/o2fzdykfKs1PSNY6J2JZz10ui7l9
KJlXegx9FlqtrUuFGZywLtcOLAvpEMd6mmXXiA43CnqYh3mGDuIPu1Y1i/fe/Y2H
uyiaqQ3mWMUcJkWsyU4vXJGtUtPIzGeAVmDfpZPoFDshBHTZSXh/hbF89rGyK3Cc
BgXVJ2kAu1La3x9esEaBgV9pmj/Isv55JoQF395jfXabB4ro1cbRa2Jlo2SEY6p+
fKlXI9MItQ8ITlJtNEce1qAm7SlZ26c2tVtwablCad4qhtvffEhrKBCfSPUOpmKY
r8/W0LDh8NqPihiwChOxDX3HJYShq2Ln1H2VnQQWfQ/BuxXQdopNnSzi0QgdCqrq
W47NFk/PdVLxtuhVdeLGgA2JkSZa4BVDcp5YvybwUW5v//5aiqHwnCRhTcrfJVKi
goOxRmQhieJqE9ea8k4AJSfT4WhYb8Hk8hO+qHy/V5VVzJUJlKBSDFptx7yOG7w2
lGXEzIf0SYp8NqJhoAaUnUiCq/zwmgDLXBbjOooqXaBpfX4nyn8rGZltcHxcOmX3
3DjLqWj6rH6ueZqyGrzOlfLhXpA3ktkCUCgqB5RpYsMdq92Twzq3HcqK/5E8IJbd
ak+rfjO+uauo6kzjs2ClT0H1fhVdPu2WLYZJ2rO1NXmf9iEfjBc19sAuAc5UKx1n
+B4GcquSMjG+eraCMs4k97QE0XVq/d9Y0rJqgqbQNCA5Kguv0FDDTeb7DCy+Xn9q
+Y2mwKWjlkiRLHvmHCLQQY9sRr87lNeFUny4XFbM5NNhQ8dzL4+HLwSnhk7YpWOJ
FRZOWxN829Nue5D0/azujY164c477lKOUKkfu3T6af5EOKCiOnXUWpQHIj09/743
L3S6uaf4cHpVJeeVBj2aPeFmVL8D+iHR6DSNfMCrRs0QYe2jT3583EYWr49xc3GN
JKsCTnFvajU50gKwJ22d6kjYseZ0S/0DXrLH+zImTh5zFGAYyzJwcQn0Ku/y6xPe
LbUYYQJNS2U+7dQ9g0UID0wWjzqUu04UjFieqAzE5YQhUni5jB6X5rwmHWuM5gbN
9GehCyBb8Yjrp+X9wLpw+qfMtaguRrBkYqDLs56YOWGCAbUSZfB+38cA424GKDJS
CEx9ZNa3znx12a59fFUhx60b6W7D486pBz7Ur5yTRg4vAwTSBQojMvoFo/fLNPAk
TrphXrMisStB9uL3m0kAQB2BPkugF7LKMi1VbAHvEjQ+/6GBIRiSrxm/JKbMw1Xa
Ok69aF7/8mO5YZ52FUIrBedQuZ6glu7LZMquPUmhd8Xt1453nMYgX2qfs8UCisp+
lYL5/85RLrFtNtfK6pJRR1wzHuQLHxJ5TIx1Wj14kn4AKg8J/dJBADZ0tHXb7NaR
kt3OEVFJoEVLNOUde8EKjwZ95Jy2gZVgf6xrZL8tQshQaxvFwFun0hx8AiTy/ofj
VhT2/uGc8NZcwCXm2/BM48dwUuiyXZ2x7K0Ml6SRpZ+dY72URYlg7bxCOUGmXCni
OfzVSl0lDkC6EGyzmXeMHHTmwJCt4DaFIa/7trS6+emIH/S08jsnFO4OyBGWxGFK
tVesjOcZlFZkrvA5mB53R3Gn3fNYVvq8i/MHmMY96H/4dA9edqG664j49CSq3y3D
X812G49Ofy34UxjyRgc7VNPl26Oa7Gh+WDgzKeUuiccnpWiXm+RFk7ngzuZugXvh
4voRoTTvnu4JbBSsFAJr6Vdo8B1DdEHHfZRiHXrt6cajkGlo69B/aTAse+5h9uc4
sDrLyFzDd0C2QwxZmJEHX62Yjsb2IuYpiZnhbMG+iUmfx9/PdafUYdQf7zN1+oYb
N9nqm0dcN1qdiVxWVmlqJYAO4WW89LRcsjSCZQFJXDiPJQGg8H8BmtIaugsOn9i2
nsZArymgJP3wAHbiSMr4EHoxIT9A9al/BZSdHT0/ExrXZZ8M12wKbDHwVYIHesr8
NdAUo+DvGvRrNKgXfn4lRNeIEnxAV6RdjbVkceaiwXOsjrL3TYCXXPrwiMgSoWF7
5qKpP1qbDRn2OHSzfbL1KLlMhFsucYaPqDjIM6Rmg9TC/Cx5JEMvWTD0K2J3B9Z3
Njwa83+EVyrIF/+7qOTccq9ThYQwZmwbyfuGs3m7/SPgWc021NkBQ3tm0q+JKJhb
y1V+p7c/bOI7WlA4ZqzF8TpXkg/TCfyBzuXp/rEk4/R2JR9werhed/uDeUCEuuY3
A4mnlXa1uSC8LIw2igdps2qGh/68d/Eua0x5jRrGLdUkpDiqIpFbl0oGr7FVh/ei
yyQ46NkzUs57IkYjcvisvAL74CdgDUWT3cSeUPROEt1gQwlUYeNCuHuUZx2B2hRO
6htDAwBoiZmQbQTO2BOLB3XyfMapK6VlYPuczLw45r8Tslv38yXrmUwF1Lldu1ER
FyU494I/nkVaTYoLjDswKwqUUDwEOYxOs9Pxn+q4VmvQPGdUHqdht8zB5XVqO6y/
OexznH0oHqqoF8JTw+iezXByRAWd+NYmYxJpT4xrx9xUaP/lX64e5qrUENG7B1sy
/HnYSYuEdYB/1yETvb9/qnV2S0yVITh4EI1sSjgzpuMdRZ/3JoV1XMAMIqXbh/tv
FwZ9hl8kw5aepl0VPGODYe5+oEagTYbegoM5597Z0d4zU5lGA+cFd1Da1bH5eR25
B4uWDPhrezQZNVguJzX4JeR3E/uqbwh1PFUycHQrdQbxKdf5zHtoe339n2eospBG
Sw46td8kn0X/ZjHtqDwBkg/i47DPrs5dgUAPcEUQ7p4qktxFTC0ZyYg5qG+TGPpm
jwwy41fEzjSOGPXBDlT/ilqjFRySFOn/gPb+Ay4DLlW+c2kyUKVoLFt47y1r7iBL
KWt/m9INGIv/WVBXaZCfVfrdl2B21mEXp1G7PC65B5gtuFy72sKQrkpvCkMy6g5m
EmdMJAhVUrfxm2GyVRsi38AxoIU6huK+SRyFBJYWDpD/bI8wo2XL66DDsuWOBFjq
/FO9r+ekgvZ4tmQjzU0sBVZIIz2im7W4G+adUMPTsaCK5RqipBeiDv1mj3jmJ8wG
TbLpEOD4wi1PtoikD0F5XhfRqdBhLa38YJCtrE4ZeW8C3OQGO2BqAsZYmPRigJfH
Su267BHBzRxXSz5KSYVDXur+mYm7/XPQkaDLisdpeJm6SZ/pbWwgsZHXj9S67md3
FZwDFAsMDKYUPrnVJNSD0P8BL+V4iJxVf4Z+xH3NYv1nSxs1xtuO0wUZ3SnjI+Gt
PFN/9X3OsNMqMvLS0dQIf3oktVVLZiuzB4YWGT7onpFqVIijyRywltrXvFNF+oOP
9/lWJKrEMzizAabK8rtEd5XhtinFC4QjMBNqnHYtaKZjJMJhcitLD68cA+sini9b
Xuz8ANBdqVp9ALOgPagKPfsXCO9/o8qOmH2WL6eAENZUB+CIRIapeP8qgcKoUqN7
a0iL+wgRn7IKUbMGJeqqm0MtdnXqYy3VuLryuBF5SpfibP8wIznyFkg0KnYTLum6
WvgkNJDUwsUwAxEsw7UThv/p7TQhWFnFlMU3Z6r3cg27GYfYXRRQ6jqVJ8y9gRHU
Q72GNd5cH6Vy7Rqhzicko06zznor5UTT2KudACVdznxC68Y8iTMh1YJncB7fAbiw
6mhHM+Axzfyn3Hc32cf4yCU9dUCk8UorMQHKqTv3jVRWELykmnRNx8SMnA8cqZFC
jZkkbrcDmzFbtqr0PwVs2B5SCzucjJWdb9MBWeW4671cwJg1sT4v12ew6O/6idfb
zhUAS7wK/7LmTAwHyWmX9h/RxPVslB7c81CH+NfficS5nbSchHlC3tTtRYZDJ/U8
8p3NCX13SkClLHJD6Vg7flQy5Bd0rlPlhnFeLuyqJlj1FMMQ8ZNs9G/GjiU4meH3
8GtjDNTv4mg0Z6bKaHCw7ffJQs9v9H1cn9lPczRdew9XybMsrj2GH8cZlUCF4mHn
hGZyVq+9Bp8fmY5tlLPlx8yVoUD686Weae1N8Ed6ciR2CrWOs9Ti0lC+y1oiwrEa
t+G3F80ChPInvu33BvguI/evQtaH8vMVbgkpxLfurNJNGpQ2Qd/80EjOU1duvVWU
lr/rv+7Xt3vMZDFtLrSaTeu6R+D98XKtBPzZjAEzyr/VilMpeh9PuO0x3/y4MFUG
5s3SKaYDAALbj7V7w8gZJePBO466rjQ32jeUKFpaJAAinXyXeW7gtrqj2Nn2A7qM
rcf3dizU/JlxBozWwZXAKxuXbXd2zVcTFwC+h96XclVsQm0EGL5bevG7gM5t4Vi3
0N7X/OEIm1muxqg8JOqNwhS/DrfOgAYx6g3M5zHsCpxTCn05oc4FjNiSU1MirQJ+
+5FLDJDrnWPF3qGTpF/ko6+sz0tPufwT27uoajR3QT/Vd7H2WpsXWx2yOz7FczIJ
G5kpBhZYe4xb1kfdDEF/f4Qmw4Zt4aOBQygctcbqN1dEHH3HEPSYj5MKNWdliVVw
D/uVNZpp+8phixTpP4KAmEStsdbbXtTmfVYgbXE5Ew/5lyWE6N95gIfidBf11geb
18dO++/am2dFDXt3WZ6DkIx5IAr+E2Y/JrIRdsnAd/sn3pHTEH+afIlR8PMWJZQm
wXIpV5Q1X2vwjVuR7NbCEW+6JhXqX+ODWQUhJWSqoZVKHORSXBYc1aCw8AMOwoKQ
pZbsVfcSn76CzETjSZHS2CAdsCY6RQ6w1CSGj/5LHqvaJZUMyKKTyrZ7KAozX/6L
Jbem65tBskZiZz1ccvcwJxF59GFEw9RLk0SsAg0LDKaTLidWBM/NIkeqsk/FTJFs
DRz5QjHVE3TElcVlnJXjKYhWWqveTfiJA5zQMaredsKv6SbHydzAVTCcyItd98Hd
j4REo3WnmhOw5TpHgiLPvY2ighvj8E92T6Wjc5wnZQscaxAbv0A/QyVgCTZ2jdks
0apT6B4fOdhU7TrYf1I5pqFCVlt+TwGp6RayV3o+JY1SeIG6uoMQuK9upZAxFwk/
dtha92mo2Oo6fzz81lgDDJlsaBumA8GqnZ+LHNA8+TZc8L7YWrYm0T+w7YO5vNxp
tyRLStL54y7nhhMeG7y6vQg3OANQxZTu4dkvT5GjshEz38Pl2By1w6Vn1R1N7NdU
nRi1JvRLPo5JP+nbjSGlSxs90fe7A9+KTE0hCwX/7FQJjFB6caEDv+kVLlIvTrOH
+VgyR+8Euy5DRxrICMVQQRtlkxuf9LBUmjT9D7qCqwJMqNQqaKY9BvpGCsOLdqws
ieFrEQitwEBiFACQ6DEc4wGrE/dpsFKAEFIWLKq359TucstK88PPS3X1EyEzJccN
RFXXM8ZeOKFLB7gzpFOuqfRe8Zk9Lg2EyoEosyZDyJmhpBkUG8oIpqaVkY9dEUHY
ztlpjhvRwhzo/rQ/0ZVxSlfbs+lKq6OHNtKo8jsgY7EG1NqzWktnyy5v/WbZQ7BZ
8qpuAPf8vU+7wY5Au797odAEVjNrnweb4uufUFRwR+JdzdawvwAE1xEBeW30cZ2A
61+FZdGWzyqDzFDV1Y1gm43axgI65Ea3NnGlwKFdXBaqdwtWepIMu9c1hSZqotZV
GtTPPZZb0FaQwZo9fLliWKLNkAG+833rknR6dYnvlhOcnK68RRnauFL3ftPcEBdZ
OFTtqsGfgVWPE0MOeoI04gMMIjsoiFAI0SsjMd3gKvto+uqgOMdmPBOB1RT40I7U
xRbNLWiKiEYI1ZdzYjIb35a1N7kytjbp6k2nk5Sn+jWCn0dM8M48VbYxrrmQDdxZ
uVaMyK6emOUNA715zEHZ2O2FBPjNP6Tve9lyv3TWAu3RNCL5LLrGZv45eUR8VE0H
7vQBCgmMlTV6qBt1LvHKpqKY8jI5gxrZpAia6SoUFRBtWVSd0TvslER9Zp57oV6R
b6+Mkx5H9v7moxLp+NDcjIcfyndS8DGvwz4EMUlmBLL6HFWkXfPXsNHIDd6QQX1Z
BxnMnHUlrZsLC/NSyJMEpO42Kh6R3VnikJksGiAxpegTY/RC3O+6dMmlKoOEnLkW
9+91hZEC0PuuhjgZjEQLsfI+g2FXLYl2oN9weS5VRUuTb4hz90i6rX7kSIntpBY4
64cZT5DP4bk/IedYRd6jX77AbZXtZ/WiAl7rZch4Wus7QId7mmo+33lHYaosQNO/
B0rtw6HKB/wHOheWkMMOcSOFXKVvCgIB5fCz7+bT6GtKbSRx0WD35ny8suOZNYpn
oqpYojfvQzaj+PWhY1ZLw5mjPlibpV8zAEM9WmhyBQwGgNBXqmdUT8jzmLJBFtmh
71xcDDbODiYSF/BaUgk/fQzXwxNGN4j3XITElgeGYFTtyFgxR8kJl8pBxXm8dbTY
Copm0P8DCez4EvwaQ0oteV2j6ePWG/iDEaZ8BBvRsjHfaKXOyZvCFqmMxiFTR/8j
D7Kxxxn3EOjn/faLwPlW1rz1Jn0b+PCCE8UjjQugiM5g3SA3slcHqx712EmW1So9
5dOwPHI/zz0LVoiKEiq06RTWRIyV8K9NsZIImoeSfLyvCvtsr+6X54tLkn8jaGBs
mQaXtN+lr4XJwS1Dd2QNK37mlBiAolX4MOf1Vt3lGrV/8bVEpOFb5n0qcC+8zYkL
Wg3dcP6nP6841CD3Q90wa/cb8iyTO17EQ6iywcGU5RQa4iSYZcUrV4eeFd+ZN0pI
3Ao5NSnizSMnmnWPht8T6+vyQZZ50tRdxWs+FA1rEdVLSWuHvxJlsI30SpSDqlT8
GPScOgQYEyBkpNCCy7CezvKHoiz8/P5ywFXxFpaFCCoTVbX3L8dIl8+exvtpZ3cD
pUzwLW0TTp79I2jV7CFDSJaEgKRUkFvUrBK1dWPJnmj3pWINqXkTEF5d0PXOoGjy
xLmgYk1+wd/6Y6sMAfrhbcjdgH9UbK6QkH5Wgu0ZhO9saRbBWzrEXk6fakRgkUwJ
dMtU7RmGKXnTPWbHvKHqqIECx00AqZJS2Rnm5CygceaiqJLao1a9qaa9KBIi2e7D
q+a3ifV9SsiUnAoPPUHf47kgeI52j6hmutMmE2XAvZBE+EoldYggWemqyLXFOskT
fdolO52mnbmoTjC5fd/g/pcp+/nhnRXX2IZvjOOvhXQhef7PopemH11w6dKXz7mh
MDIL+MBSS3ku589+HO3AmbIYZeUveWlWxRbZtI3HI7ckM8IntLNDvGqyhoRvr21J
U7AvHDWOOPYrMUQXPf0oPHqTXXZy75chAo64qprf0LtkN2g7/MsKwUN+lSj3UlZc
AkM1QeHA/deTiD2HNPb4RpI3GmanFRWk/m4SIotV95wanj9c0du9j/jmH/XpKlW+
5GCRj2ljkeYktse47X3VRkADuuF1b16RH1M4GoaDp5ZNtQ66pP8XlZfPfGCRAVC/
2CurU16ZvmFvWkj12QN7RARvLNJblSffAKNArdtmLB5WfC+2NQBa652wPlNu3/Q5
InIR3oAv+VVWWiV1EkM6XmQYhNJvePAnVgtAba/gq2QPZ7veT/bxC5WpowoF0Oow
qe4TXz/k9eZwFhRsyzAgENqiDp8PQdwdyQBuWgQGPmR/lc2z6x0cG74MX91nfQFS
r9kbx9aPP6OEdP+FZsupf5q6aclerXUJM/tjxwVvvhMyCrZG5uBzQzsbh/Sj/g8i
QUCGE/OXLTJ0VWUUt1T9QAUIsFmpyDr4wsFdeCZJHyGxVVI2/HFRPX3Ze0cCvHRR
zRMLMRri3D964ALOaMqb49pcUdo6TIeaVc9LcAlAFaLVZ3iDTEuR27wzkZ1O8YnI
Qd9H819L7oAkOIol7+eWQlmFKu7l5P2QnqjM8EqRHDlkcXiVWEyzw72FeBL0+xq2
h3bLPG8WuUewEOVRMqwruhKHeRH5F43jcXhvFeq2B41V5SPhHsxkWtCP8hPCtHeE
/R2gkie5TWALItTelpSz26/cJgxU9U7nLrfUVxACPyv5nbLf3s2DfNIFWOYMxfzJ
P9Mh+jQ+lmqjdry5fAgraSZPp8xrZ+Rw6fwUhZ67shjYv0Q8n926Qs+VK/H3/rNI
Xqp/o9vzRoJtkmCgP+QsXIR+okdh363m0aSo/ieG4wTxo/SNeze/GsouCipvITi6
rvhnZ9S6GOgKs8vf1iqUcUciHtUXPN37i5XqjKjclBt+lmS4Pl5mPxev1ftmQ52C
OW9o6sKsChmcEl0wOyGe44h6FuiuyNJsf156A9i/AeQrgYYNUfiy1TD/e6TMcW4p
xvYH7IhWadhDLLJLXvkMFrdL36kF4WHG129lFGPakTTLgGdR9dh6b2RbxQMSSJRu
X/Ue+PhbAmWKaJM2ryOD6AYD7ApLuq6B+VtTmQ9nxopfiXbJrx8jOo1Yv1X7r6NB
PddgavPCbfKTwJuJJa78K1HtqBkJvFosNnSFnE9o977KJZ0Z/SkUBR/8rQWf1C3R
1hmH9yFA5xVsYvW78xraSWDlQ9h5eIRaqmHMwuRuUWl8h7i8vTsxYmHAWC1suEcg
W+cjghgRQaPjnj1TFN0TbSyMg7uH1/8OoQIo9QxN6ebwztVte0DzAzs1SMvIzYr+
Th3w18NMGaUfscKseUK+15uU4qA4dah8dIn6FqP93lK+YzpY/Jfk5sNcCgBkY+oe
KzpQBX44HD5KtsIf89RkBtVIDVULuMe1WCGwO3aVno+NNnuWGQBGNW3rp2bmIy7w
jVK+0MTjlPp2M3hGA1Pe9N5ZFPE/yqeIGvG9iHoiDTbLHYJvthtBJyby2Fw3jhkn
WoOC6SKHfRk857DOE6WHQl8f41MIqyd5ElvRdDlnTSHdsA1YCEZ+FNdp24Mz5Sy4
VLUUVFAeAiXr8tEz9q8GpftL2I65SYZiCb5NjODYjpzghLHQ05a2JwcZCjvBJpfD
arc6XzF6keMyujV6dLGbUwXuYenVbpMlWUq3LRON5Tns2tCplRCJRarB5yTEjDBS
4t2hZVx2nThWr11/RJJaV1zHYn7+4g+O0/yWJZij8N7hATZYd66WgmW43HQoLEJ0
HIbDBs1jCk3o7jxkFB24AXm2BRTsho6K2qcSAShKjoCZJDUCx9VhXDul2kqK7GBp
/cMvFilouqiGPOoiepDkn53d20LxqjL2B9HI2DZl4iUQ2u+7Ur6xSyN1VbcXDXXq
AXuwMyppvnPM0LO5GnH4ZXP+WPDWwQD37doymVwp/3uVS9GbO8+c7C3E6caNB2Ki
9w5dWnAX+aTZ7dh8HjqohaVfxFGuzeyoLVf+C7lGhwu8el73iAq05dHkKCar9DT1
neIZZWZ37BBC7P57QuQFNHFa70bt0Ql22n9ajITg6YzSRaQOSxy7lwFjnKue9DCP
TqRhKeQFasXtpHMqYbjHrYV0vEiazJ/9siNBLb6TA5b/ztc8SHb4arArdFYRvWbA
bRE0N8LNum2eErLhNebkm6ljNZv5erqfPRg5fYitvnYBuISy+rEw0pXamq7LzS87
QlbhmxA5lB1l8QYjnJKiD6wixDs+ueeT8D1isKtvDgHm6VEGptvGqkYZWAzRQTfQ
dVp+DvT+o2DOiID1yotmPBjKJL9obcPE8+851sQBLz/nY3u+rCl1EO4ZvymCZuU0
qnpbE7Sx0X1MKnZUOe9Fcj//YHQ41IOY17V0VYCUXTwI5MvX6WqQGAWZlKQxQ6LX
qHn6G+eOer5Idwsel1H4ua7e8Q5RNI392xeHw5omswosGbUevNzPGEd9f+9/ebYa
8KCG12dgVEcEna8xQju5o4etXfCa5HRDG7YnxBiu2/vCfmu+rKeF8CwtqC+zyjas
WZymXjfsmA/AiWyq1RrhHyxqLnd//anULMAuOQgH7FZgsIbn9FI/A3Lad/0vfOLr
1trZLOi3OmG0K8s+7vnxqX176larKCxdHcXXjgYg/yOYHvTaLEz/7z2td/LAi68T
q4mkAyUBqn0iTHh1zJoV0EJULtuilG8/ujvg3c7RIeUFL7150/waDrir9fd45xop
0BBV8gXj+GSbFxJN6luj9rkyzwjxrC60gXxKRRtYrA6VZOuLJpdLwUfqXH+DfrCV
PiAJFtgjcABcZ/JGqlUkNFgetaF/idVcAR8pt97CBgbry5zB+fzw6p9a20hvLBln
8M9zBJ3KedACR4P9gf5BK2fGeBFjUdokQdk5B4gW4Dvrzc7IrACmGRKHsh6M6ktF
T/GAT5cDPGMk6tHNU6pKNMBTKCn9ZQYvjnJKzyWvWZsqWs6Egp0tJJ+YvIXanzD8
HHnDsaYAcWlTt1ezqVvPheuSMdrFqPA2jurOCjHaFsCx0CAHPG3xB+HfIxITtLVU
+iOWXtUePrhMy4DjyKbWBlxqqN9dK+iXRc9KR8+xsKW36GakDD692XI/xfSNUtnt
YK1ZOOTvbREIyDzSEjL3cKhDRY5oP1cJABZ2EpCr0ffOLi3DWvgrxlOrh9WOQ3jw
QKtxcIbfg5wIoDrfmxs47SYiU6jIwyheE+B2Scc5PnAArhid59UmDhjU0U/wqF8v
T4B/SZ2mir+CAViu2it33ZnptBW7uhHRZe3HdFZzPZnD+nwhlrMkAnqsIJbqTRXQ
vCw3Grp/Ycj6KoEE0mGI/uOl59DnObZgis8NS3gW9Zfn9O2VD4Od/2/fxvmLkVD7
Iq2M/7Xr0hi8zSkzF5G/saUXsvX+l/amvRiidx+AelO1UeUbyJ2FiVsYWxhmTwhZ
9cu6M0at8JdDsyO+Bp0rQ8bIWYJX59H2QcpvExqjCbkciVnR2URw+pTT6lJXSGL8
JqFZHKS1J9LcuFOQaD69Da0JEPBml01xTz/VBBIL8L1i/ud3j64419Q4zBrPKy/B
kHPuQrjRYrcRj5hgbvTHyWenD3xolUA4hd3wfga+sqdqRckm/Qx+LdfSQ/EQb2pG
Nj3+YF9y1locifsoFMryVr+moPHYHd8K/OjR3WMV+zTZBjXRxmPbhSNT5hUlRe1P
CPKs/RwtC5Q2yyhNd73sQJGsmiQfjA9R3jBdUykO8yOGIjGthPRIOdg4HsYJDAkV
ukppe9Fl9r/oKuoC1Mv7osPFVlP/AP2MCgflLKOBe5KKRqHRxWEtLn69wl5eWWfl
asn5Vavo6p36VglxjNf7ngpT4ig627pLeVG91m0F8CZi80DrsDf7y6r61Ue7b6Gj
X5cXao3Ak/XvjnMP8VdmG8E+fHKAzBOBuTjpSR4Ick423iEa4OWQ0UMTZIJcqeMb
MswQJ7Qeymv53S7nxJxrWrTbqKhHl9p0f3jBdWi1VVqkY6wPuWJ+GMpKaquBYRHr
48JzdFWZCkoX7CimNvpb5Tmzb+qYZ0m9Ivv9sUtJIxhBEO3iVt9C5UwmGPsVleXv
kevly4tjtHsDRH2BrZ9DEdf9WVL5bm3BMgvMUjHCxEC+YbmqVdSiagEegkeWCtlb
cyFlsJnmUKB4ncudEWWIdjm6YRB3dEVL/rMxFScyeU3cz7+od7uSulzywmQ8m8+A
GMQmEDM1NBGlNmrBU9aLzzJdEhg6Sw8qkLSpr5dxII9TWSB46QM4jj9Jf63mkjDQ
Ng5juW2TvTb9qPnukwLsx5FpHxcMLJmiNvxkcnV51GpsGwPJKaM3Z89Og/LVBn3K
XW8e6Sh9dLSKp3hwBPF8xe+UmldmKL1sAb364DlFm2nCesEA4j3MZLOKGHf4mWja
26p10xaIwEGqpIaPZd/u3w9TdvHL4adpi/cRZNU3G8KEjvmC+DH2lPvOGXE3JQRt
dI2+pc9iyq/c5c4NwXZdKQSGrGfnY+DH8qb/oWhyG+IJLT++U4v54nTKF83GdYo9
XR+AHuXmQ4ZRbk7/t7jnxZrHE27TVUk5iapLPL3VepFvpmLhJRl8J2IUCmm+22kJ
bID47Ek/IsYvfVNV74uSCM+LPNABwNnuYjfik2Kk6eUNajFrvIK2uLFLXZMPQnWP
I1UsxXw4nkP6X6RuuUz52kcUj09oX+tDXDGtso9pnKyTAShsJUXvDAIARHOIGlBc
e8vOIYAayKf/E8r095wspOmKTl4vPoA/Rt4ikTaEOx/u/FASN8Wa4GeY+w5sSKU2
5ThfvPBVRUdY9ScaG96tlu8z2KEgYZ/asIkT56iGrq5DBqEAtAdbSVEERCRGajfP
4llFRoH3YUVTQmdzKhrler4D70QnGs4dz6870qmbZE4P9szFTWj71P26ed4nCLQQ
xUf0kcapyl3xAZf/H9j0GRcF+UYhoupgExkzxOqOt4Bn1v169s/j72dzcUW5tgf2
M4DOGGTEKZ93PFH4voe9bZv2hFofFKydohYWy0ZRUgvjiC7rDpbjKYCENYhP0K1B
8TlJGMfvNYz2hEj0oY2hsa2qFWNiOJTMCWJAwYhtkb3KvnLU5YgSBvAeclIBVqlU
d0mJFb8Ghg7oMA6hGtgY/fkNR4cRPjb72OPt9rFr5gHveh/L7UYgsiaV9s7bEYgG
hL/Qzv6fsE9HTq7+Kxg6CHfchGg7nKlhUaXJzqe5MICoyJVpmYPi0zDyIvCNqDB7
OEynuYylc9GnSPBfK3fVRHXezEeMAB6otX5nGCNBAAE7XfX2oyjRy1tWo4xCZrVy
znvpQvS0emu+kRXFvMvhuQGv+Wor3hpteoaVejpBGg5X/oFeiEk3JACoUsyIOYiG
Jwj3fDL+5+aCR6lKoxB8ffoWLc9gCJr4ABnaFIVolHYUzPj7QZTaJZD+cm4mxdYC
CtYwVzzkSxwwJ7IyskQoM817FcRVU+k1qJC7eEQx4NjyrdebTar9D7Fuy1IQGzkN
wNuXW4Aeg8//Y/GBmW6K03Cmu/dDD2g5ljwEEtFppO5PLSZyDCxkMc0w5o7rVPYm
r+vAGkYbKBNj+dCkLZKiBqYe3G5BD2PapceilOP3jUuZefy5EBbooQOVPQ+ocmKg
l2kSwvFSqZ8XhVMWMi+dTfV5epRvIUQOxDZwqeJvGPY0HH6XRzClAiQ1/as4vp2i
b0W5he6hRwm7DB14dLA+3xPFF9T3RHXbrY5yOTJWoxSsNY4EPzsHQhU7baDiaGuJ
wn+YXcrCklVtcaUQ0S3BySOH3RrW4mj0Gf0c981OQAau0QL2U9dYgDPaCGVHPaU4
bkVBFuXyR3ILMzOF8ZDiu5IHl0JyBv2tGPQ4Xmewb/KJmndJZmqSYSjjRxaWGU5B
x5WFfRafc2t2GFmE7afdgT9WzLTQVeSorYXjA0MSLysFGE1EKTAdV/VF/5uD9EQY
H1Fgggb87BpQxxX6z8B4477XXFrn0OXtbFUbi/UuCZ6r3F8GZRA7NQD8z5UbwBxJ
t5nqaC5R55AOaFtmbMkfq3So1tETnGX1z3tRo6XXhKUidaLX+c81K6SxYcoJxQfU
FklFqdGfEYqPUjUU1SeDmpEiHdOG15TZ2dVf8vxgOugTVb6rchOPv8Ov827H2ph0
STvnYmB7DaRNShNhdlrBb3yFxLuCQ1+fBeLiYU02gn9uvONQLJ36IquvnVhznh7H
tsK1haNmSBdA6oSKzoBcQ8EB62YQDPIvgnuFdugFnm8ocVBMUy3lmiNVnqS6sz8p
L63QBqTyWT58bmcyBDZCzzuggP6TSzH9q37UAJ8BVnWGx5XWqyeiGXTvlNF0m4aa
BrE7g8PObHkqiEwzlSlbVtG13KJFi/sPEo48Ou1uBMmZ2Y/fwn5DVY2/mpfCdQYs
m2s8jyBaM/QETtLXTsXnAIP7T1NlRk5Wvo+KLATgXcjxTqoWe5z69elWxwsdH0tX
XS8MAUdEu4M+AfLD1ua0R1QXrRtDLmcbJf4Nys86rR/YRmq0bS3OvEcGW2sn7yQt
Ay0UntIqmJsCZ10I4zgrfhePJhzVPV6sQrwEG26BR6yGZASF6Xh1iISPFrNxcuK/
4BqnA/Xk8cEGSEueR2FxxHzwthRv5eKJuHo/qqw2wp+pBCBQTIge3FA86HQHeSvx
Tx7i/kccjRePHYyeuK+1cFwfstDncAl2YUoSmpMR/Tr7V301dnKez8VR4wbyUVI+
DKfMH2bu0ssOw+dJywzD5l9FG7y9V3ZoEVT3zUMA6JCzh1bi8NZU8uLCA5aC4Vjv
M5TEBiP7K6i1zsiTkJvquE4ZrHnO1oyOBSrjG6tomIUwvFLY6dsqIkrlzqLaoLfX
pDGAtjSx8XkEE4WrGNkB0pc5LvQ6ffLMJgjMz3Nds0LYV3CtODvyCXMKf9QM/+SA
gOEyqwBvSLDC/1XocxTelsZCDVbGGWApGow1wnm4uVrF82ML76rcBK6VVoaoGcdj
473n/ck7ChNpZjPrZEHx5DfAI+5atnJHoSeBq3ldWKo2nzLkObMR+irjPWMTq5x8
Fj5UGTe5JTzp6MN0XBTPkAZt1GFTkFazjFkG40GVJGaDsf2Fjf5wTWne8ADF9/W1
yieLa7BVPqOKJoYCL8lwd/NTc34ulhTKr/tR71jlCg6/HGJAbR9SyyglohcU/MHJ
a5HCnT0fNEb7RXYEUUxt3OqdnKCGnkeegqrpmxIwbF/HzSsyOC2PE4SKcSUkyEOQ
CXVjgoc9JXgajJ1txiD4qVpiZYqM6+jaNjXUaIlArEfVg/WN4Wprew3q0d7XGIlT
hhPqkLTn/cVmqVjMrW2r59niPVbGHdavRhEibSjhVTjh0H3cFNXTsre46V4x9JYZ
nORX7GejIXh7puior84ilppGdIsbNcwXOsfFe05zSxE1+L9SuS9Wf6tq10ldrgke
RBL2iLfaqg6XmPotIBonLHGLnt6JuAU/K3r3ZVm0//PGLF5JlQeBPYfUqzqqLjkQ
3HEI0VWWcfFkMK+Ltf7DubLtHe/R7SyagJQ9H7jRD+prXnFlKP5dhGyUOqwp2DAT
XPVb1iGjoNSrqBhCFEHFe6OOYz/cAGiq21p2xbpJXGKVlTIfMu9nzkfMciPw6HUb
c6Wp28TW+8+eZGgYYTjfnwiiIJkKxeTSrzEe1AUikTLmpwMXTgKnvmizqbA/LjnF
qBI/WkdRBovHziXfHTaX4k8Rfxe6OPnhCj573FWzcHfmEwBqNO9piBM68VSkaWBZ
up48hYQyJ2uSn3CYBU7h9568p5CLhT+Fx16YqMCCE0yiX7zcWFc/VTyr9IA8oe7N
yXbE9m/OfeV5pLJanNyntjcarbjplvsgE+pgNs3XDETshx3wdqI8vyH7y/X61VqO
QXAN9tq5OOEk1aI9RRtxH+kcsxohyd06TVbhNiATb92C2ylYszrOIxsXiAkMq+4U
INBNnxVHs2cbSwzX1v1Tt/jwtiKvv+K+fH+2n5F4wgM0mWO3cGQ289p4BKBXofF7
2T6yBU5BIXEeaDpJgDIfDG1ergpgQ8wCsexskhqVYRxJRVWbxog2F0bql8qviWLL
CkfJqqM/l4uvVx39xz00v4cJ9IfqwzzWq+hP7lse07Lqkb3A3Axiocic5iJnrmyv
hIPTJ4xFNgAORUSrUoCW31OIwegEdpfxfnYpPdD8kGT/Rs+vz915rwYZVuagqKrf
RzlfQNrWLsdBYl6J1VuN6MEYXm48y9lVlEewzZDDMzllVHXF/0+atJ5djgagevnh
Y2zLKPAJuVbBSDcsfIyO/2YFdjFkyTlb9H5/hMP+6rtu7kIko82L1BU6jr/3MZYt
VT4s2VWMd0twfBn9TXBbQbWf858XJD0e9OYJRzyG+K0NrLZqj9yra0q4OVOwD7fi
fXOcSem2nFHiLh8BsBjkd7RRPWjPiHf6jZ+Eg7Mf4olhgtZ8F645zD4sk+6iQG4Y
f9SYLsVW5NnYSNVhRac9CaId+3YIljgS9kBeAg7hfiPbrj+8PNKUW1uCxptdjKPj
rBXcLUrg3ml9Z4kMHG35BbTZ/tdEQVI5KqXz9xh9L31uOfoU8CdG0b2fQFbQEaid
rpEVmlsBtianA394JakzPjyA4nLEEdFie3oHHQyBZ4xVlp/3nre6BysNbqTrYXcC
cpyAzXtnI0OyUZnE5K8lgJRFuPsmpYaH1XFhkZNspbhfrIWGa36yg6U6NnfHcs6E
heZQEDBU81qj4QsZz4u+LEdWWOLQRrHaJ3KZboBlIsnwcxbXpvOzkaVuyjxvfTHm
wl3nxlNZbD58g6/Em6wVU65bijJK/jFkAL7WpJwGZL62ftvcTIFE7J0c+l8HrTR6
5yqJmzE9ctZE2r1s11lU1e82jLDlNWZzliexnl4uSO0LgBoNPcNx+VY1K/K1Kgvr
Hk4DdQUUiG8QqbzVvESQ5pZIGFQIMT2f2RhuNHsmVB/dym0Bnsmk752lmFCztOSS
KcdeTK7BHzUu6RHmHZZW4yQkY2f2+E6V7OV5koj48gZOa8hAo3wB+9P6oMLgF9jV
F9WAMYMK1ccnnzJkzibaAqA0C23l4qEORiGjs5OFW27fp2Z0XGXSu8qK/9d7Bj0I
//hzwHUjGmGDOXgjv5d9Vf2scCPDWFCggKTcAs3tOgyImkuCkzUzLfRqUGqZblBF
TYelJ7FQccTYCLos2jQNLJLKVQ3hxrkH+OGdzhQDCIsw+/036NZ7LeXp/nhoBwJb
SvjyldO89jEs71O4L6dCp3WeSL3vyXkCz28Ckx3guUnw/phFqddjSKNkzk6WBUy5
x9n4v5rRs0u1DhcIFS7fHNiAr6RxZfIDFQ1NThSxBhPJ3LvhlgTPhhKC7mBc7c6N
EAhymT6OZia/mIgdLfhAl2ano3I3JhaNUhoosY6ErpYecC9dnlvpvbqoGvQcsP8k
kGXqjKyLS1qN+nG8+ePnP+sOLzO0F6ZmbvOeYfh78BOPHqreoeXzC3r2Aw1uTpfd
O8z08/jMx3nwqw4ON0je2cO0GuGoNTqIXHRfWWYBYAPehMQ5BjEk9XRr+MedcmPJ
P3fCErlkWsdWTxjvJrp46MX9yXAa8cagYw4gINKTCNPAXp6Kp63dRik4IC7U33JM
vUhgLSHsGRUvj2hCiSncGMCyJtgq8s4GJw7a+5E3aB0/iAUpT1cCceyPrIT8crll
i/Wti2EA1W8neZdH0Urgd3ZcQoIJVlaU8Muh9zt1tCuW+4Azc5U33WooLIe5hpH3
kPIOG1TBEpKnn5y2flTCTLoDHiY604BkCOribag9PqtG3dl1FvaS/f7i5I0qhb0d
RWjH3nP0SuL/TFYuseheyqkOQqF4AYQ51SY1GCh468p3iyBmsjNOe6ZhUbt+A/+V
16ad4ux4Zs0zwG8SY7gdoY38FsHpq+6XF8m3E7uPQPvWpf9boQ8ShA+ypKq6lrkT
USMS1t4C82ER4bB2BLN4lCSV/d0fA/lkwys9iMvHxreV/4slRD61RBWmZ0NNlgxn
aV9GDZkJ6bzfXcbMlUnMvDyBtR3KeX9z6P8Y1FyKYlizgPneOOhBJhx9uVt1Tuta
T/aly2nzurNendHAUXBgw0KGQ8B6DhBGRdNik/eqMs7BuY8CQh5KfGf0+ajfeoOC
hARZhYyZo9P9pG3VNEBqaEOzdsAoTGIE0GmPDjx754TrtUVba6rvUZdptJXgEOMS
c0OCW1mIwIeeGfklQ9WMQY38WFQr2i94tmuFqHykIfeQMA7Jz0GKpd30Hd1vj+fM
NNMzBDkH7RdtC9w6m3qI+pSzOT28UdCVs42qLw/oEDXnCSvqOPBfLJwOQAdRo6li
S61yif3cb8FePBIrHkjBmyN/uGuKRa8jjATb7FCkSUiNWq97d4xak0qGM/GRZFpo
Zpc/t7dGqJjM9m76ErDOIdArGoUD2WQF0DVkq0g/KMu4Yn4qZmBJ3z+HAkf+mktu
+nTRYUE5nuOLtnV3lCJUOsudMq3T0LmujtrBzsnEKmPoojeOOS13Er18+elL8xep
fZEG1M017yiQP3n2DI1x015rOJ+sbIOYegPotw1x+k5QpYZ7+/MnEYUOmVdppWcd
Ky+y2sxlUUBCz2zpUgEYz1lxmG2HPwQykw5udbNP2IDgboQ04miNHKYnHfrCFs6U
+KexwHlqJmdTlSu82SgzvrquSm79P542oLkTfIIViPszV5K/LYBKEgCC0YYp1V7N
LTjj9+QACvL7PNmcROrW64FZjVNsqMJQaNLeggr/ZmfMDGBWvEiwkHzGZ4gbHkdE
TzBgKuRm0evkkuPKBteefwiEjJfMNr+4wU7aJUE7ebN1ITVHg41OpyjOTMLTNklj
/dmYM9BxGxSiUzYc4UDHc14fOgHGnot7c/EWWuTOFMCD5vsYIp6rFP+mgnczE3D/
wN6/scf4hbB65R6weBMJO3tbJH75GsraY/Su0ztkMdycDVKuRnf+6UYXCkv0ow9M
gFgANVr+8jZ8+j09O/Czr0x0R9vSL9ioFCVMPE44uApFbqojge6j1FeHvxrCLuuI
fr25jc4xALu1LHFMhdvs8w/bqmhiUg07SUhBieQ0PmFCvG/TPg8+hi4bNYCZEY4f
JlZeVl6TvxYzq8byEQCukzRHO8Pg93NUBro0EHUq/XF5yliHcYgxBu3mHbQMNONU
fZcrrGqHycOTmjrD58UHiBXE0JABiWoW0MKBrfcMuhbUg96B2+YRnGT+MjwkML8T
98Vki1EXH+g6XVfY87d7uzV0ksY1pZPZcp22qNjF3iwWejn+vkxOEBAvhkWx7y+H
SO4OSwTLaKO25GKm1BifKWH1a84BVXTFQEA9yA24LWNln2zeBg4Ld7wb1TWDscm/
8piV6NrLWdXt81GQY5nMqQMbtvwrzW09ZE4SEJgG9ZS9vtcr7QaBMMBFQfCVwK9y
KLJ3hMdmATsNnnAauEbRSAhTBJclmGx4LUoRrdmHKjs1NZ34CEDycCFDx4mqpmh5
cwnUJfcamk3TyLGXK1jdKKFZiD3USoz1EOVJOPNFNRj2vmXcN/bZiF7BZNYjzhlL
vwXmZf+yp2Def/FJMHrsdAd8wvPQEbcYi7g53VH1/0nPFp0J/9n9VnWQ/Md0vScX
pACbTnvLlgvoB0DEGN6lVqbYk1sqbqJyd8rFpadVmJ2FWLhC0A3IzAi0Nd+nilOO
W+lR9jVLhXpUA9FoDAKsausitv1vLlM2J9TSHw0VAZ+m5tc3izP0h7EfJflqmZ90
AN5s7BJkG/Ok8iblk5n0st4Gnauj+dL/tg7tWL7494u0pXV9OUsaSifWH4Yusmxz
HgRt8Z2xcctV0itGWtUjpl6+++1S19X2oJFwrE2Ji65PgM18H6CJfE32mY5Wmfdc
j6JUoJJ/BJwMJdXbYveQafhCpOnAIUPZ6SuQZS0jN3L3ErrgHgz86QWKywxVt5Dy
D/E2I5bsvp4eFU3LK0NA+lCyGMcoiq78a71hlc+YCSyktkJLMCqyJHzZ9INnQAuP
d6lDPFeY46ucoboZtQA5FhuFAeLr06ywz6lQfkNeQfVOItIYqLNx6vUw1Gb2wI5G
on8c2vUMHvN4PAioqRVsPf3tK5X/3dtYUEeS76gp+nmLLGSOGhaeEPENIDylm6Bk
1nr7QBPNriOi4mIaa/cV/6oDcfM8oczzIMw+REnVjNwuT5Nc5SbNXWXk53xc1G7k
VU4uTWG9EXkMqH5wu5Ry+yoX2dq5geE++v3F7Vq2NW4A72uyC6VRx1lFxgi5FfpN
aYLVAeZt7UPpazTs1tPISYEmxBuovRTE5XeIOU+iS+zV/bbQubBnHcbRrONrbbm9
uwjyR68ErAm/KGoHYzSUw9hJayWaS1LqEPIpSMLEfp6Cs/gNiRTrsC+cmnm8nY6s
/HejG45Zx/sHcwVouEyE47wMxWR5ms5a8cuCF2RlIpb72Yps6xWReAzgGu8OAQBq
nXf7xXzCljYrt2wSs/dUZY7eSZJupW9pOJvmitsqKOk0zgSo/c+PrI6q3y/rjHpD
hmwPoMiEBYgsBb4CDkVunjnZpuNrYZolwAO84UZ0YPWNt4rQg/O/f8M2hG9opSRw
+T0ZrzgiRDyMbpNnZ/iS19PZuFd9xRFUMDYyxCeGT/1Ot4deDjIC3+O1E7Dufgv9
ZhuwqBhSC3hxSqV3hmGMyLCc2qB8MvAcDC0HaEOgTDErxK95W7s/bWioo1uafdgk
Wu7+xDLSjuZqc4hiCcztmYTPsCcT1XAEwKpAo8NWwOr63AvX402IZ4vtd/RiRNcv
dWtT4+F75BqcPCt7K4psdksP08f04tW/b7oKXwvYay7FoMZpWER7SRIxMlTMh62j
lUFKv3FY4Y05fULK8J73fOIzPCZl8ceBN4BszYKgTpMIM/zI9512nQygazIJ9nl5
po4ajF/h37JN6VHZMXjmAf3XLTa+vR/1vRWl5ifnUOxpTmcgpgszkKTykDZBqgn+
hJZbb04jlveycvOvhwHRND3Czz+O5ejGT1Gk03A6HrqTu4LeiMq1MbGVE7BsY4hD
fZjqd0QyJ9P4U7psmXo5qpwHobUd0FZnaRZRNs+RrvIC/wS7w6buOtWv6BUTppRA
j7q0pOc9ii/VyQ7hrEFDUHW//Zwv2j3qnOCyVHXnsWUO4FfHxQagve0zUojOJYdd
nOebYObuxPawPXyh6+4vDyEJ+J87qj/QdOLm4WJRt/ulpCnbW4lANbCE4aGUsyZk
OkW46UujdfeaXozxDDgNamD7pCJVhYJobe4S4vB0lQIKeCeJpXCXOfZWsVJKp5jA
RPTcBPGlErTvub03AAHIFPHN/EVZ+HobrhylgBazYsBN0gs6yhbb9YUbNOol4Bls
I2yDOw7kdH1YejDTNj8Khro2iWcIv55Bo30KLdC9pEcFWiNVdjSOXO0DjhH1tVXs
NUjhfDytLp5AwC7mMcLw7lreLlscg1YlrxAi+tcCRM8wUO0575Kp8jFphgH1PKcC
sLWAquKt58pAdLoIxwgy6lkwgO9kXbiF1WcRkthcINggCcbHm/ivfMMfqTyhzsw3
CvGghaO4NSf+yp51dHAAuWabK3YVgQcURVbfJ9Gwocq3x9xPki0vYPpUCFyUvaZ1
PG9lJVvWkAoxo+rctrX8v9W+gaTj3Ur24q6QVi229v1jL5uO9kXQM2GZXN9Y2uVT
FL7SHo7cLQeL280XhuFtoenZUTxyelQCtYiu0C50BnJXl12u6ghPQRF/B7TtWoBD
UyxlTDSojGyw41AX9K1i3euHdyZF0idWPTc0uelMGzgPpVEOl9+WYiZEONhQ95ny
sASh2zUnhr91jRWheFUcAYmXAgOuGCu3TCx+XbQSAI6imLFJwNPEdJM802USP8O9
aDZ9DqhYTOnST2/suUGhbjBshIDeCzguSZegvEmvE1c6n6HB7HE/5tZj1bZLNP76
XpNNEklGQaMZ+LFotJU1VcJzZqpsXdoiv4xSKCbbw/qQyWQMliF7aH9QAzMR2Rpx
Ws8EgvhbkKBVKzi41GmilNsjDROJHcJsv7hAAXyh+papVLbHh3ZEQg74C6/8CBiQ
CbDIJuUSrr5I0iqV0WzSVt1GT7PSEqjKAflI9RjGtTes/7SQsm4eC7/Tzakt+EWr
t8RY6uFlKDXKCuvlvQpndRg7DBbdO2MZrsqKj3GU0iiYSQKnK3hfF7LtzG0p7YXh
z+AY1o3eG23hSq+uRuWiCtIPXx8y1phdM/tnfLcS3gmBIEYibT/HqLwj0hu8UOP/
i0SwvfsKobUkgWjVrAyLsK5GZokteAH78g9b53mKEQVuLsjjpvOWZavgh6JpmKdv
D7CZSku7iSbXOCTawCe5yh+H36FwpA5j4MoCTr2nCvgFF/I1uEVcRF9E9z/CxcP5
OxAZVnEXLQ5o+Z+dKMD3ZCosQk7PvwovZTx9V0+qrh6QASeI4H2MWrouaZNbRW1N
gWsfg72hpW1gM4JscvWA1M1CTRpjD/od8g0sOcy1YfAjxtnNrbgaVDkAeuxQ92MS
aSbVBKcSc9vWaZzuy/yKHjgXhs1e4E7hgR/KNRx7UGPlxUi4IPg7cWU54I08LV6J
2z+rXfCX7sP43mfB0eYbCS7rMI+oSL85vbYsp1vZctfd6qp9PLX01KxH+bjiuIOv
PfyOSPv7Lb+XMK24WDInMff+IPCUUxCChBDRVNjGRuTshqOO+M/42JRUaFFH9A8P
pGhE3AVWGpOXCkCKCrPoVaK14sqfmHB0zheGK415LrJ8qj+P7ZjLDiJu3A26X36r
qoQzSASrhnshl7iNCjjnhONqQn6SpYNHS1F5jEQUMXc1lRzWcRXhItvJdPmZtjMT
wcGJwU6Brs7NadHqovric8nCC7/X0iafRnEhWgdgA6vcZF+xMEuO/e3ueJxvOI9H
nYAx6V1h6X6vVHLdJEq6zhPT0t0NfkuW9H+j3zqX1at8AYkiyBQ7nnyl2KJd2SFy
dq6QNWEo4jHBmEOWUi1liskisAPaujcNE5JEwTPqpsIayFxUJdCMPm1OCqvy02nR
C36Qoblmv2Xk49dqf0bEKwCXVf4pr7gim8+lWqE8I3B50vwDvnHcLqaSAX0mC0In
DBe4Cu4Dxz/bepFm2o3He9s0yk8scgVAacsmDZpoT0WpxI9BSPS+FLld4gmSSSFC
f7RvwmQeaU8PvtnGLTjas03iOO8OUiIdydl/keG08IK+s9OVWsLW7sjgG7fNKkI8
mN4xYO+mfUnXSLtLEx0LzU+oIYexchteFBYRmIdOb+qKTSMy48wbMD/cwx4e1Aoo
B16APixle/oJDuPxJDv5XnPiNhmU/TIjsGhJcNrpXYuMypBKZarzVOBJUo2vVoL3
H+NAo/lsJQ2rqNi05dJyOaYe9U3Uv2fofzGGc3EBm/Wm94xVWqgf3iz6H98amvAt
ydGQvtp8NzT5PlG6D2fpSUTsEK5B4VmUvpQATp289FI0En34oiJj+qPlzLYJOdql
9pnCTf0CPC4Y9y/TKNtbjDHID51G2djoK0NOFzeylVgYW09+wqavbXJHxBcDgN/V
Gyk+evm0PHznxK7j8ElGCSh62L7E64LaKY5HXpvcPwzxSZ/893jrwAAA6Mh3vyho
iwOxeA4xJ+60aI3M0MXFH8/2UD7UiENZHd+VBZpdXgy6A7/PtCarsk/AnsJSNoMs
zBT9YdHS61M1gI/tPiGsyc4RVOMNgLGdX7C3eRmkcM/I9FeGSlPDNHsrnTIYZTSB
xtzcmoJ2QsFwqNC5MmErFFEQs6tQ89ex6Rrd0L83sJnqKVz3FoooyxJP6vQ7AuXI
864VdijU9FJsEmX1OyA8SppYwa+xrAbut8GW9Lpz9O1tkvqB9PRamxfXIm0kkCdk
tJPwxk4A/ip/seND17fnpB/8m3bQhIRWhsrSeZkYeKOlJw7gKo6XMbdZgSpaItuO
kKKdReuvPOKz3rc+P7N6HZN2ZpabwNOq6pfezZnRz2oeHAnG/q+deNUtNma76kMd
EiEMnOfdqMfbM3YHfo60YQnLQ8xyDjBoTpQKfQAaXENWwUyFHlOrKmbZF7BBIH26
m1AsKq5QMTfPpzvZ/R8NMulFiGOe9+VhEERtxQdVQBruyWjes+MTCdIKxCiHpl70
KN6kMdyDKngshPEcrXyefT8ZX7buDBxYyzgxlYOClOfNUgDtQMa34qEPTvWc10a6
IwAJ6oDTBPWF/+gtIFbaA8wElOdsHxWCFkslh4MviY3HFAkNlqe22MM8o96m1TkI
FOVgcYWeebvfLRGCRiNPUbVTFSVOvJNJ0UjZ1eNVxZkr+1fVQA99LJ8OmbYGTcGU
6rkZYxo52/5Ei66yYzc4Dsv7dBAAiFE1Pg95IeaiihyEjJ+boMJK5INvP0okvFB7
Dtae8tZDc0NC2gf0zVzOtRxFVDwIY66v2nv6tjaPcNBwyAsiN0jqmunhv7Z6dsw/
SEqQL8qttsVF2cH37DvbKTL2dTfjf686nvg1ufWnNYcg2jYkhWjZnu4P2IiqjcMe
mKcsBbUi5Y/Fo+R3n7fhrA7a46zlqLYeJKveXTMgDGo5TT7LaHYGJMXK4VU8x7ne
GuGzHmXUZkvLt/RczQXxKTgROGXDLfNXn1bJV0sxn4x3VRa82miOrkTkwwFTCzSZ
wHGamy035+phytjcxDdJ+T58xdIlFg67PJXNxwmKra5N/BuBY98TAHlG1bbv2s9v
iM3sqaT0VWNluPhcmGxxlweA/vzA2Pk5irZ+D9xJOhBo9POxExnzLiTMkQqK5CxV
2t5eLYnEEO7AYc74RP0tVoxZdsc4a/VPtok8HChn9zaHSOQvPs4aa6ivZQgGZKtu
DY/IA9j+sUDPilAHMJEaCUq36ODbOz7hItNEeuyVIRHTXOi61foWV7wJ5htmop0W
QqkH4xcOt95WQIYkTo4DMiabX0E3uN40WJjK/l9+8FecJ6F0eq48lHuAxvTsjslW
fjFHnG0O5R7B5mmZTxnF3LOVRs/ytV+y42eFMazefI5PpfWNqm7scOjm17/+ovjW
fmPf0odO+5tyuqA7J1hbBq8rJ2Xqhh42BBZSKZByNFRzgvBrE9Ia7phr9wVRvezl
ufCgxdbvVbArXTjzAaKZgcj193oRxRWv4BH9lPXklGt3SLycOgUH65sZRPMR1Pw8
UvXClHp7D2BMUB2lWy4I+HgKc6gpvEob96tBO8sm/1IAy6GF4yU9hW8XRxkUbYEM
RlEnGy9D4xgM5fTqFELVmnNkdEME6pWPDIcuO4bB40l1yzBXxcSEDcOlEjpBWqns
KBIuAFEKzbIQR6gAMsnDqaPdaxi30HVqB60woH5HH9OmRAEKz/gGdvrjU6gJO9wL
fPO7LamHKbE0QDKcVznJVQDe8zIS80yavci7ZiGV99NWbjX7h2u9+/6cZQfSK7uS
bBdnPTRql2GfCRTBlsNBMNdc/wyzZt1lLQ4JpKFbancGiu+MqFMLXUrcE83IsIPM
lZdphlIOy7tex6wZf8dyIywr+OAS3a9CitLbBwbwJM4PBXNkJPgqp7IQ1k46QOj3
91QWn7xb2pOdMFLoGbwbluU6exXF9P30R47tfhddmkftGNizptu2UHQDDPkMTMEQ
MhVI0mUalX3TQraeE8Ee2HmXvv48y9GczJyIkCUGftEFdtoaApf8aWzECL6BOOtb
rc1w3tMz2reSxUJ686zwFI97NurXDuvwmvWuPEQJHJR5Aq3Wna4QPKw5su8Wie9S
mrgXmkAOZqqGq2Oav/sHq4GXUSvcHjk19++mGkjFp7BjOKlR/e5lXEKpt2UqBwwJ
gP0DlRS/bw6Ju57/b7OQkrlUnjwY2QLEj9oisI+pJgLoowJhoj2m8lgHn6HIGLZa
8vZcCtbIrMO1NAH3c6dC7ONljV6fAdb8dj4qwHMhAMT10LEnUx4HyZUIZiHnDC/l
LGrlIDNORM/qkNvCOpUer1b8ZM1AjVhPAiva0tntJqm1nIQtY9ZvMJ18etN0TsDt
50b+qdWgmWw1i2DSjn1Q/Gbi69yoOAn1JdIimgSHOpD9RD/ycEUNncxlWm0Yc94G
Z5/GvVGWOjgj6QV1WB1C2aLETlQ6Ky9fPePIRQkvzCMa+Max0DmXTCAiTNlWYnx4
G8r7B0yUdRi+LD3HhAklC55H4QrAhibGTp1EFcp9jbSIfgL7O62/lAyXY2ehsviS
W9qD7sID8OoaRK7sna8XHumvZpxG3qpg7HKeCbv0ylUG4qxioW6IfiECH94/jGW5
DwMueCyPWeb1pYoEk66NspLacYJkMmLoyUQ18tHndHZr+r3BrY61zxQ+ExK6BvgW
rp+a/XCplZqQBepuxnOBve2e6M0+cqssUY49QrUajBmNUKnhKa8Ff8hEq8OTUV1F
bHCny1UI8wNFOllRqFbhhxH0xaWhPgk69aE0PkAXPulLJbM1yT0ud7ZzWRMrGxha
YhK/xZrKBvFLGmdkMP0opsRuSlA5KopQA59L+Au5xj2qa6pxKb9waiIY92nMzG+a
8eaIvmZp67kCW9ebW+5cg6owmBodJ09klOfjX48INlUJv9E8d6Q1jh9FujP+WkhE
Tf9Qrl2SnYIS1EHStjPA6q3lf6sPZgnsFLxPEze3k+MvpRExH5+2Zt0iNgcO1fY0
oe8VQKdY/O1MbOnrgzrKZhzBi3uodt3PbdEXNk/gAPmBe6/6Fa5BgGMpyD6AjOq8
/c+bA+RfypdfdOC5IVox8wv4YGBWXxmI+VMEJ9gFXYHmQ4Y9kwM6ArhWeU7TgX3d
g4HKZ9JeAyQ5XdKXE9q7FgU9iwqk8T1giRjBckeBscGm1aUYScPUa02PP8MNSGkz
qdy23rxIodOBwkZTzO22LERgZPIhQgudD4AUUv6F2gRbjMW0qh3S4EuKMC2vxcU4
W20VG98Bl3XNp9E2lLLSRFM8PEEUX1iRYyRAyaLBJWhc/q0Bm+VUdLS06fH1pusG
iFW973fv5bt6a+zwUzSHXFAvX0OpHSWzFuNZ74ED4X8j1lEvAatrc4zTxu/3AAob
QGd2mZqP9s7jG+DbA5mwY0XY7FUTakDzfL4fVKQRqjd+/DrGcWfuRoVMeE+WgmH1
Airt20ZzeAiyH3PSIsTAvVEjV2LCOaWcRp456Eksjr4lqPuxU0IlEbeXFVp3EiQ9
JzDKpvMQvaIABgXxqXE9QwRzBjXvayhsvb0SKomFQSWYQtsFHiut5UH0AQXaVVqN
UqLVA8W76Q74f+2VNxahgCUw7MuA4Zp9K7mmSXq1dgUOUau7daOFUKLDjt5QZM5v
Ty24l7qaPmWkB40FKkGyes1X8rYWTCFEbVcUOAb2iwZUpW4E3LTYybl/W2kiWqP6
sgpe905ALMgYBpUGkwLy0iUD1tG8EU91ANy04HyJ9g3SpT3CpldJtxIjaq/BNf+w
9G+FZ9PiRrAgYey0Kvapluc5awbEnZ2yASHXdu6To38boZjs97vqUe4ohKIAay22
6mhk5lF4j352YAMNytCELpFjAp83CfGxoHCWwCUziDWpPsAufCaS2mMDJhIpZ6jf
bLGrpv8ex0afLb2rEPMn4stedYVuhNqduBUH7p7Vidw31vt/0JkzeQtEKY62Y2aS
WDbGB3M9CjZDUFHVx2SmEVayWZQI2vfMaeBftv+mK2bBaPUvLQdXT8s302Pe0TaX
0OYhgsiF6EjvLonAIz5BUUCVBifLdN6P4N17DCS2EKyo7JywBUdFdw5uJUe0h/hL
myzqi1lGSG21wO/fzGdyFAl+J6+yBihleqRBF9aiaHTb8bf3Ty/FXVc8flV6/bse
2Ae+Nz4nU13r1rXfnorP2WQEUSHcVNinGU1UX5qXLOSL2dFRi8TWYvLlqH5ybu4p
/eE525Vn7OSJDeU4hcQL4fboMIMwPjWF6fUU9KNMB/16SgorPtT2UzXTibjKRjdF
r0uvvt7ppW5Iuu/Fxyu566tJ9KZCIWKhRxwQPtRUEzK7TduuvV9y9xuyL3Nz2v5h
BtbJuty36UNZH7sXImgzygz50+DZ5Yf4yi209PMAX3KU+TycJemO95V16HYMTCx3
++QueArNIKY12hvOO/hBkj5DkHmYt785Zok7vXFxiSG23GDQejaWUUdmMOWJqE5Y
xu1JQ1QQRkThH7EJKMYp40a7UyF9xEfBtW8oLW6wI9rn7YxxBZ82cqAkMDKrdxqj
CraRq+09w6XT1Mct7mZ20S+cBd2k3fdcrc0hhmtkimJ4Amqh/XosmpQ4BbzPgV2A
HVYOJr+7NySQHFa+Y7QmMfJaDRlx+rvRZL8GfYa/PR8Cqqw8uFzkLdGNkEfGwJPb
f4ycyrmBsWfsIFPxKdVElzL/dNGmTKX7WDw4VK3y5EYM164D8xe/Aa/FZMrzxong
jPbwqWF9kVnCp05aqNOhLOiufyb3dmkNPJLqVpNbQo/UkqK7oPfgbQDJ0NhVsuAj
BJn19VkFZ26/cSYHAtwdOCBcc9aef3UyhUrm8Nfos6IqFEAbiM/8x8/uMMq1qkDp
0ZygaLrH88mvSaeHKMtGqfl6R22WK59Bt1XDacV8lhatUMD96nLW8JmRWZfjemvD
8KTbQDWgvzJu+K70EutCp4FCZhJQdYeM0DzbvPAKqOx69iOhvN1o7c53YlAiPgsU
8Z+yYeufXpQAOeUfd/SU4CwjKAek0Ynei6TmswGVB7rEpZ15sb0kd1E3BMn6wUtf
apjNxmczte8VtN5U6WkzhtLFuqXPHXcvIgGnpKLzKOJLJkfoS3SiB7EpVxPiTXBF
2QM7Lj2+r3lfaynQxhU05MOa/AFv43YFaIHctq+IYmWu2PUPnutt3+tprKmsj+lf
p1Y/o9bSzuzB+ms+w0R1hl+z2quMx9xEgOIeyTmvW7pszfMV62fXVJ1/YCDrcHfJ
qROa2M+PmvEAtyjo8mvnGBTf4gHcvNXueELbRzazaAZ6iqyqOkwJv7YMWmCJcx0B
5AvEz5AdS4zLlaKX0CfjDg4rD4u4OjEclQ3lU3N6UqrD2kiAp/mbrL82Z2OLSXvL
dDDE/+xewb4sOpfZSOcF/NhI+PkuEgSrIGSa9duLBcxYqEU+ynK92TE4477y6rJh
9bBMk9iDQwmDBj1Ue5VL2RoxslVp/CmdATy/uBt+pejxnSn48m7IlXmc9XarKcCp
7L1ObDp1tuqL1itsh/u4Ce9RQmkaEUspb2aLCo5RXXt2jmj039rQSiHxVhZRcAyd
c/e2RLY2FfXLddFkp8GtuaeJHFD/C3c72XiPCuOO5yYhvCtTsLkqRQ7XUNxax3ZO
hJ54maOze09W2Cf/4wzBRdQhYk5xfGaz2katHQmI/r+FepZqYxiWRE/HVJ+iLLjy
Q+XLZ9O2l+SwbYAiuORl1G+jDQ1eqWRQ3NzPUrCVLZljTKx54AxiCfYWsWnSlM3M
jnJNUHBx5hXo5z9dz2856MoWxNkg9RHctVqPl65C5ZZOS6DP94slvkSe40PyKOPI
g09x/SQEF0DAXyIu/mfRLchAnxd7v5deeDEu2QVgzQc7ykGTQiAEaQLKdTGap9ek
77Q6AJZhsCSaEWo+eCJ1y8ez4ZEx+d7OcEQ8l0mvHUzHZ82anuU+j5IE4LnnOAyg
1DZjflTkqc4IlBtj7Lw7UK16VmPrCIAChYu5mZzDAfZUN4AxvjTV60O3eDPhRh0U
mlBQVuLPJ7a0n1KEYLi6EZKx5hx8OJb5ealk7m7APm0QNk73HlM8/CeLnIJb/i+8
SbBhro8J2BTejLPAfbJaP/QiL1vw3sQ5NNFKT+E/kQpmSywytpH5EFw+uSSxirSs
3ApAA1IQxRBkb5G9X0v9juwhWUMzGHK51qQGoXu1s/CzNYi02a0Hpf3I91am4Lbe
FiRwatmMYLc6UfpSH4YuDVDc4QhGS0c4l0djtax3pDO+mvGamTowai9vve7jRe0n
XlZw77PoD5gbTzA+dYqOkWGQncSkz3pD0D8WoRsBo/LSQHLXRm3+DMU0DTs8+kvn
zO9zNoyAmVA6c4Yxb4h5IziU/HQ3IFTxFe9D2nQ4mp9mhVSWLqLsfiPjsxqGRIde
MeYumZjJLwRHopXyBD4AicTGmYuV+oYdQcr9gx7lkglDnLiUtzOc0qKfvhUoV2dN
XGYh/8ShaDsvxB4JlbuxHK4PQ57ddHW+UfyekS94oP0xMrZvHKYAPQyXQOXx6I2P
1Q1OxlkxdA0EaCkIO/m58u7V5gBdwH2jOzzo7vpClNDqE531E5eATpKAxKQqxL8a
NVLDuIgFj2iD57scECVC6Zwjon1lP48yXOsR9OomHS3UPhgcwO3sWpAlFYsif7r/
vU6P3C2vVB4Z/AtNe8O20/1Q1UmLUjz5COgfEIGc/hneg2UXUhWp+PFqVovBenXf
cbDmjNwb3yLDJOjGZJS1NFBSDRAWAg0Es/vYUiQhG0/2M0Jz7KRjF5vwvbgYJWUs
AAoqeefOeF7n9H3yFjgdWs1OOCajFe3q/rhHED+jbOAffRTAAKq6/8QIpVhEYpkc
vJTppySbvqPBruwG1rZ8iGd/O25P9dOx78Vwub7J13vaDVKYshgxSaKg2N7IZpYH
z2uv2DWJLyQ8n6vVu3VHIQVRDNdERG1e6A1qHzkmoUZQTQ3Ep6wWAs7KkExV9BmB
iPUBx9LAfDf5b1FpgsgHQmbPpN6HLssZCdFesllCDKStvvHLS4RhB6VcQyaSk9Kp
v7YIdMheUx8HHt91JvyaBOR6olzx2f2FmZPlMGb1vSsJKam9r4HFnJjM3Fy8Te+r
FfjkGMDtE8TaWu/QtznEF6LZLbuer59pkkS0dXawhWGEnkOOxvpcFbTY36iJ3orG
60hfoiACbnmaQTYhP+7kC57ixcucsMUaj7GNsffla4s42aYFo/CLOfWRwnkpyJpI
R2J0YBAB3zkQiCsyCvCCQOU7AvIfXYQO6ILIlkRzmvNhRlO0tVOV/CFhKaqgjtHJ
ur/OT303HEnKZZU03fnAivNb3v02QMbzqrxx2iHzUx8jOrrChXNV/QMolg9IdfEA
KgARmdwF/5Dcv8k9c4ZUdzPQs9Nz7g0lneB1qsV1L3y/JK2OkyC1zUkHRliiBZ8V
W092yf+VblMHg2edS5+P0tenXHZXR5texZ3UmtCENyp/+fLl5OwR7AXC1hHtS5Xp
leVaLn8XjdQNnbr+NFEHfBUem/9NvHgInwwk/iSHIx88WG1OH5BTYUG3PsugrMHT
bkqKcMxeErf0rp59gm4MHchQgC1lfwYh+52YdX4tTVOzuHIELZEmVJVOUcUh17kz
RHJy719qysic5VkTeZUfbHp+nm56mbluB/1Heme5Y+i/UY97/pH7enYaLQWh8anN
xsq1gpvKLYq8UAqU+YUh4ZVg4Afj+Dsf9rBtzJ1NDeMZJX/obpw4GoCXuwfF4Fwo
IVWNulSoQHJE6f1nKRLD0t+aMSX3Q7uUmzaGP9HfqFGx9L/Jqu6gfApOwhFtYXx/
4ipu+f1Bzam2pbKuL1HCHFFaudOwHYXlw2gex04OjPb1BzLJJ7dZujLdDdwOFNmr
Ys8tBjy1AW4wT6rgn+CWC//2t3L0/zc0//85DT+stbtWcWwZtpnnqMs36hqbxVq0
X26jn4k6fwKiGL6MIo0szcxVGN3yll/8dCWGEJmJrmve88StbCWREOIQYFo0XBy0
7pMjBJudpKKVsScX0vtCATO2wqGu8rFnUGv4yi0/hsbOrGVp0Y3S8I6l/+wRZQyz
n2xAYkVdq+wYmE0BIFXemTMroEmJXSAtopSQtAZUiU/yKw4gMQM55NJf9CqdJYgq
6JVSxXPBeXpngf/BPQgdvdX+85CTt2cdjuZPRTCN9UMq8kPE/yk4KT6m8ug4lpj3
spHanA9mWnVxh5iF7QNnkcRlWbVFO/HOHAAT/pB151dbma2K6pRpQlJX9/k2dqHg
ZdRxwuZXWb9PKttTd3xqMFQK+Vjc4h78eKLsr+7F3Tw4EcMquTYzkhq29Z15Jddh
9uegKkAYREuRgNIhNEaLKbPiz7vQJWHn2WzCaPivjK3KcXdLpZU7/HxAjzchY0pk
SPHu8/TGSTCGYKOB1P7DOfxCVjX48KuO/+S5JhwZWEV6KfWsLUpBl8pqe0BzjVv1
35xxKuATvwT4exq/u76Go/aKOQnjAJnER4QN8BYh8NRAnWaLTqbZtaNWsPTOdLfx
3xsns8MXdeXhB1nfaP4Gp4hylHDfb4wIf5J2BcQOScKJV/WMrZE6UrrA1c0g/cfe
2cKkqDq6Q78Y/EJtits3QmqgEEgzRIs4kNaIGJEmPRZUPdBAu2icfy+5lptwbbmJ
jsTXs5pfUujk7lw+O9PhHgTno+qo5WW2X7U7QxZgtVG5KY+NCrSxYzj8X4Fj/vc4
eQ5OswLS7pD+/6P29hEyhdjswRXNjRgp8g1m8dkN+7Sdw7EWh5GTxIGMFWFv1akk
/hOwzcbZo/DnyObsUQ4Iea34YXItJklJciuCZaIQVU/zHdQR/nhnbyxiHxXGaTNH
Usl9tjp7Loe77xTsQEO+auO6JmzuPsOw4E96dROgNB2C8/gJ4kk/jNuVijUs4Wzh
ydlJ2GHYZEfJ7Xa9NBODFvHo5avFXjdEYGPGxcwXIV1Q/RnFdtlmZcqbt7OT+DhB
qJ5PN5iCeX9IakbRcrxjLc0NTaikJQPcn9EV6cOt2ruoqtE26ZL+Uy6zm1oA0i8j
NjRzjJoZqlZNVbvDHr2WhjVIqk2Q3bWEl+i2DdxfXcDnBvXDqxjRRSuwVQnTBuDy
ugCz82gLZ+3lhMvqxWDqKDmk/WuExxAjDNA0mGNSu7SbSozdqHIOeENrL3mpsPNn
F3d7Mb2OzZAHsYginrt8ms0PQoAY7ah/+kKCfsMGKrOjlpOyEow16nIITllf0Nod
RJa5tLZmBEoXT0LH2baz6Qx1cmvjcWHS/QFZb7Di7tnRmong38ooqF+qvlr9xHw+
fCt2stADvvjCKfqyiuLyAHPcTIbtlyO5dAPtEvrnv/9WL7K4Mvnb9/jpdCXr/KO/
O/OO7d0pzHz6T7jg10s6r5oEWdksVDyJRM6sJLLtbMkQt9Of5g/LZfjIlpaP3Eey
sf0CcShYjEYgI1napGbKnc9xocnsnIo9ZHUY2/yIn+Yj6Xb/AkaejlN2xYIxHEE6
y5GJoHL0aBVlfLy+/F4/J1rVFmUNPaMpWNNKBxY5ylf/uWe+L/GXsUkf2PyEgg9J
JIy8Aec7gpRl6mgq5MTe3M7z/DOHfcwrXCKESS4bmCP91tu4r1oqmAUECLPMHKNl
zHCMV3KKKVc5LX1jGYWofaT47RUu1pgK64O/Mvr+Ac5fqYWijk4y+oV8SohHdWCW
bvaLek9Z5Lp7jrlgtXf9DSrHfjo68RlKlS3fPIeC4eCalFur4DqRBQzeJ2GCfMTq
lwZNBU41w1jvWsj7sNDadficlhENIdhlptffrHXQz1yE8OAgZ7ucD6wLSUc9Ki5I
xB7TcF4xahjdsgtNxn8I8+K9I+4eohDoCyRI8EMSuNq7YOBmHoRz01lzFlK839gH
7+lETDm8kTffwLNV33+ssq8O3cQeAF17vHvv7HRv3EMts0idSd3aTYBSP4RNrkSf
1SF/afTujZWM0kvQ1/ZGYFMThBS49nofL1HkPKP3ccUFqoEpO2cYJ7/QBk6uKSGF
gB5fGNpH1LLzifEapz7ZfDm7TJ7ELhZzs8q7RPomjIlqgZqCebClottMqCxuOJyq
VSFenl91X6assxN2pIqJZA9YLGAybp0DN1Pd3es0q56hycq7d9caclUfuluSnV2W
XhJ1hVBDJphIFSOyxxvuwG7qucs/kEudjTUIZRm+ujltbens9lwXEeSF9DC6BXUS
WkMyN/7Hqa5WBKHUtcnkzEH3aO36L/tBZKXzKyu8eZmWr6By0g3HhdWfXqUp++rH
yID1ZWh+YJJHj4XRYzs/Ad2FMzVYjVU7SGz5esUxoBmfLJyDXE5aMIaO7Jwt0g3a
YmkjLi6gSy29wlBIyTiVri+AYA/n6iTGzljdyYS7yYWTCqBcjXHE0PrN59jRN45u
+YaRoB/3Ip7CjbTraMOG0xVA7CqlJxW89lk4qS/0tkBSbanPScw38HNEZyldFTtH
KLE1O+Vcenqr2PLWb3ffYR/1R8U++dZlCQjMxg5CBQj7WdGv0Q8h277BClbmaruy
b02S+nA1hsoRdm+NDBITL1o2PB2eEVpVKu+RpJeA0HLYpsVvhBQBlnBCtRKGXm8Z
aSCDFx2vctmZ9QVQGXF43dBJS8KMimYhWt/l/H81niI3D/X/mUsxSi/zhjOXAgCT
so+Ofzowau374xtd2TDk7/UThz22tr4dCmZ0tYnm6Wu+X0nOpwD4GWs2QdVUWkmb
ueJDm97RQ3I+4onjjhGJpuBCObbAK02WNSvWkvZyMktVYnSQTeuUSmln1/kW7OC1
VgYjnIaIeeEKJaIVzd16eRFu/8tXIi9g7T2NkPaNZtWyGtBE172InGqFu/vMb5/S
I1ZGBG/G+gasl1ak/eVwTHuquH8lW36Zn2uPJT3S+PXSB7KBuzDzLGbsF/ojiPpn
lr7nh5lFQXS4NVc0FVjNaewTT8XL5rfvpLlRLpKfZTEr2R5g/FJSRoxRwQSVAGuC
MlRS0mqKx67F5312wb8Dfr+h7qSiMJu7ajh7XbM75pttypVKDNgASDx6b8D8r0QX
HZ7A2tW19mO+aShPcWMWUItoL2sVQP+faHsKbFBREbvLXgdt2NvyKT/iyzni9/Qc
biZyZYuqKFO47I4bw6TtvwK/9IfSghJsOF8HXcScJY6g5ffw8WBlpQSBlHphZGzN
rFJKF843DNER/yRFH1bf6nONtBOcaH30+TTL91sELJ4+c0h7t6HKn2w6jQrKIT0o
Dq6sBqkyXkHwpeKshoEoFVNdy9nhj0v6innuCFFwweaY2ETGBvNLTsqyLOvSEFml
AR6+sPKdF6esjseaqH5MvtnylyUDpP3yBELsVJmCk50MjFXcSmrv0Tc4UOvmRimP
TxvDLLclYEtD1PMcVwRkC5L3cgQHdumZmFpyv6ShVdihJ2evUgbxCqMQXjn+eopt
Y8e2zVC1sHGVL61r50hmH6gJfqZBAX5lGtOl2IC/FFdcu8+3st13c4pzMKrhpzS8
vLMjcAJ62HYh4F8x2rkhqHN4Livin1cO4t+tJC9SK7TDFl72t/JMmlgLCm3+1qWj
JLFN8R5qgye8NqcWe9ixzdAdzEBmgn1ac7wrmjV3Q9ZVdj7D7DGqLlIn6nOwP67N
UFsiutBvOviaeOuQj6uWgsKNaTd1LRTmkBsEmHJheVKEnvfi2Qeqxo5Qu1Ko0w3K
vvo2ZDykw2MdHmx/K25pjLhCtWLdW4RENEg+kYF9Zs2zgVSRJGunRbfVqV+fcMCE
yf8G9aFRLg71ol3K7HFu+xdVPM2joMCwhd9XvpPvu+tphIMg1ZVum6d5HRJQp/yv
ERBoC4JHWPGZ1OGAdO0ROew0H/x+gPIHevF78MU96Dxpx/+vUnYQeFqt2DR16zud
9AQqL1rbgIofmohaPU2spZT8f2y5Kxfiq+dvoA7qNFGEd9QToR+dR5MgZdc4Q5IL
7mnU/oOpFTxU0ttSbgT8Gy9dAHu7HiokF1R9M+BmOJgZm6mc9d2rngEFx09URpeU
sz2sQYgnbN1s927kqc5z3UgwsHGe8zjOhxNvQ1EWY66agoxXtT6ahtzY6bPmxVfv
6hVSSClo2I0iMsKHf2Ud92R2ZoxxcsdQO/Mlvm1UDAkPxVfOvQ6HbKSf6azxJpyn
Exuy9IXgGVgBRmTA1QoGh30C/UkzPyNWC9iWF01dhWiOT1+vxfEQTOF9HVTON63T
mDi/jZechypb60RTeLNYNu01ZUROq/5RARAeNS52shmiBK1Usud5d3QUQN2ZJuPd
PB92M8iiAzAoMEzV7YnX7Tz5avvmevKgvkd40/IDomzf6lrUA1A5RprW78WcoeLA
LsJRSDL42hKJ//fwJqEoV7KUcZH8FxLHJXjOy2G2CXyRk+feY650ruKNdWNRbGUL
Di0L0jREo1y5K3o1/SBb8reQyoNLTTmpjENy/h5oItc2T2r4CF6LYbEj1sCs+jmx
0fNUhWyFNQU/bQmsC+ZxW7smBqKiyl2y/MvMAXqJ+Xx330CJt1dyZn6zRkddue36
aAXas9tbOJvobHX51FBugxk4/O/eRtOklowQPniC24iDCrNM7hjzHHRMyljQq2/C
CU+y/WsNHgWt7gmL3YI3bQl18cdYsNaBj24lJk/IAymGnosjrssdY9dhXX4sV60r
Dc/KiKXxwBuPFLtDyXdgWdKKYAE9XC0uPd4QIdcYYhFFQCFKGJpQ90w4b4ViabWO
6UeULUyY5iELn40ebw4Mw6uL5TrYUt2azn4ptA282sW2Sggp37jJg/HyksxElYL1
s/TuNOlRBZJ3NqBLpx5Zp7+4jr+sBnWrSJViaZ2e4RcmlzWZW9JlIHlWiReaVh7m
vsyVJfTmoRvUtJl55m6Eh0KSMraJD2YXswHfbFXKrPbauO4oF+4IVnjHCya5W6eI
FVSkd6F34ypp4MTkI3tnquOhTUZodKd99rdvY2BPqyE2f8Bu2ieGKIkirkwWsLsP
Z9qkQr6ubqq6VmIF3W9jSdgzLSx70C1xcqM7OLbihdF7iJVvgyfGr8PN4zbsNIaH
8yFyAdIfn0LWkUQWbMrwke17HikSRpuNbJI2qHGpY6KjWXNEoEQfU1OhI4QEiihG
86oIVB6Ni1xJLRgP2yIp+iGgb4V+Cp2tn5qDkGNKQ3gGZpuiLwZn1LGdNBkqOm12
7Tkr3DakspAJKczqAlti8gWI2ySBwS6f8D5IB3FS6ra4gHgThglpXjaBdWpR1iFd
Tvic8pbaKFbOpdKRcoQW9JsnwbxHE6A1smlttUdl0Sc3SrwswpDmuk4VonmyB96J
bHMQST+LI/tZlbSbXzrpDvcvY2psu7VicBHzJc7l6Gbagbwcxr9jq+Pv3KOlW3La
sik46bj1AX7wcfqwpMvJzJX+LtQ3n5iFh2Qti2/667GNcuNd7V3phZUzkQ5SRJoS
RI+IblOroHZ7eXKWb3Vit3jhrxJaYHZlbQoDrJ/SEVtHkQQX+pLRt95S/dS++QNh
dD8eNC7koIYhUXtYXHgsKSfGERZd/Ljd6E6itXBkZJE1i2QybTWrFZbYphJihNTO
4/KEJ9X64QTV77WIO+OT6b1M516aSWIOYg/gMadiypraMKn6jJKi7AJkWL7mquAm
tgcY2ZlLjPmO70rNpUYTjmA4TxozmsJo95WqkwMJnATcuw+MQEfaB1u4DJ34z20w
msUq5XCVB+7nyHF0L5ML4teRfdOirDl2ia8Urvgzacez3QN3bKdbdYcgnsenRZW7
ZW5YFJ+Vj0DXQ31c+B9Rfry2XP6i8Kz+yjoEonU1mC2Fdx9UGWrYS5dTYandIcrV
Xb8M5jL8hxy2gjTgXkFFl+0QZH+l4vKx/myumKYbh/LGLXlgrgIz7tVvxe2umktN
ahOpwj2Oaitbgist5Iq3LYoaffjMAgbwaQ+PuBT0/wc0zAwS9lhxLMUHttrvs8BK
ON1qex8I7KW8bi/jLekVQdEaARfxaD0yU9riWKafqk+p4Cgz+o+x+jVU4KpOAtxx
gbkkDPVt3/o5TyIMLEbDGEbcNONn6fYxQx4RPS8zytx2a9VE9un7XTwK0tmj9IyN
4dxiY9H+87to6zpTH7s5J0VFBGsqI7F4twm2Nq7dIuUNhY6Su0e+HOnK4jNjIGZx
LCsYEAAyC+latzwUlyQDQBQW/m9rbQlSon8RTkhHpNUgnjnqJjQAEZYOrWcjZopy
SvRThLgaZEseM0FmDXX5MPEU5ELbhhPdp862OBk5PGIraDuGb8eHfEQOxzus7s7J
4kWn1zP0ORhxbHrzI3VlqIGouRrLN0kQ4PXq4HKK0y1QKqcF/SM9pM/M7nfG7tgP
R1zQsCp17383VogJ9USOHn6gQxQdVSJJ4MS+zlTsyBlHtGckPSAKmbAiW6GFXt8T
uF38W6iD5UXmb95zHrobkBWig97vs2FVswFpuf+diFtoeoIvx0mjcCkJ8b2hp8Gr
3Vr0sIkDt0utOGSklyYAHKbjkF7krBa0ksgTOyvxH6VLTTLikfsQzX8xEf/dL7mc
r3n2Hy+ugkGyWTjPsOMboTXDASDqz8ZxEf3VBj4SpyeZ2VDXot11IcmLri0J/h+7
rqFJs27/mTgF+Ld85vQyQjiAv1Vuy4TxIWjZvl26k1m1DgaRYJ8aUXz0SiHWIaT9
DvUx9M5F1rgPu5Wo6AtH0WIRZzn/724EIqIdgT/RWowupqRWPYH0+1J+BsU2GeXJ
xL8aPXCmG6092K2Fdl7+dz7MB21kgb1rTQImJtT/CJs/zgRerwry+IpZbO5QAhPc
mMxDV8tHl0YUtfA4PLxBe1NyfqgRKYn/6iB3CK/H/XfZ1zmXh7CwyG/QCrf/WN1l
PRu15oGa+plFfG3A0T2W8axuKcX6R/IBeHfjegf8d1K8z3njUd+o1WcKtZ6gLMZM
CUJ+XPNfeGABU+26aC1q0gVbaShpbw9b2e6qxQnuRBKut/PX4H7dNnkyN3ENAicZ
c9Mllgb89v3+31TyOTd7MMPYxKSULzvc6B9is8EQZ4kJhisBTGM50JUV7ycx0RQl
GbrZjXqfxgIUEGD4bYNMbEDmtLqUD0/VzuOxK+VHK+jAaotHn0Uda5m/AndLhBS8
9bjTx9OIyXgZHKCIl1m9PiL/9PrXXsTABZhRtO6mLqRSwt7zQueQAfgmW3tTEznC
rqPgPaXBDwAbwVk3fzLhI/YLLBw3s599WCvEQ73ZdDZR7dgmoTT+CYmHbAO6FB7s
XtHiFSVGv1SCRrBrdDLt4xzNALlX2xE/I95teKgr3EyhGvDcuaPCsJtuYDPWuc/A
AQJS9IfcAdEwUU3XITOCSeMcnBnXN3UEVt10Ile7f3NM86SXwYmm4dvwoKHYKYSQ
Jcrf37p+adMo5bYSLEw/I7NYhCMNZSFgkXeXyKdedOUz6YeCSI9MlZbTmPpxmhDd
QZAfi4BEWTB2woW5F+yDxinQmhxzn9I3sHWhREw5tgl1FlxojrCiFrtcji8A2wh9
Ki/8MHJqni3OSxLXMrCQizIRIZ0GJ/EHcNeTfv62wiP8FtpLugAFWPQ8cHtkwvyx
jqGllAqymTk+FNlUJQjUA2FpPJcQbpsfYuKEmvu4MJRSIZADGI/lg4xEv+PFXUoF
OXj3zPOP5GkptP2c5cmRaiMdJgPTT57VtfSxjjPB1A5s9s6CrfL5NU5UEEwEHrKa
9OvFxSvtIHkdAl7vjQyGGr9JnJhTxYjHORlwRVciy0V2H76YueozWVz6npQ2S8We
TvLMg49UOq0n5o46zFhj6wdlK+GORc1+3CxJBDIuNMd+yrtkqB8Gx8VnwdtT2AgQ
5lHaGgCUrfN6kJ/jZiAjh9G0qnQr19U1oQpBbl9M1DdWhobkgD9EeLvdO5pbTrAb
zyCW2nwf4IQsHYVGOjq0abIOc3Hp25qeMUje0919JOxSAYY3Jp3YtGIlY2JGDj3P
TSXpWGPI8ZGm9NInurMvlKkbI/gBpe/YJQnvMAMegCq+CaH0ygEkJZeJ2sxxnTRp
SdeI1E1t/8xVypfqTjsz6ZGKUD3pcrD7HeTGpdQEs3RGQMBt63u1TpLU1Z3epFf6
y1chhEEmob11WjDNTsRyMd2WekeDKOzyfBT/XytGGdSn72UcaBAQAb3ns2L6LqhV
TtVCq43no/vhhAcvzBvykCBP01bqs5iM7Ib+8Xou839AKiJj+or5QQMmqpw2CXmn
0FaUu90Cew/uWAoPHarM1NZzz1LXwZnq8X1gBU089MsSFFRuJKDltvvznMwp31Rs
QvFWGj+NkbKOBGfUEqYt2zleWebg/XCXzEO1+1qzJNYa6FYKFZcN+vqHD4mx+192
bcDCS0Jodlg6y98souvr/NNfR/tUTMo20hh8IuLSnTDQaoKn3FXhxy9tjeEYh6Qs
lHrVp/31FZBJ6++Ago+5/193RhxjcDcagQDkVdufjNmcQSUTLyiYA2o2NqdcxdTj
pLreTAAOOhnigxo+66EWvMtf4JMXUQ4yL3IF4OGe1HyDi/UIMCBb8P1uGQccGdQs
wfQRzjdjqflwI+yqlPdSKSG8zYNoCl4vAJiuoe+/fDW3BGDjqBx4HwiLF4aFTwGb
i4jGqk658WiSJpfz9Y4hSpmfuwMFspfgHzH5g5j8GFtZNyyr0QZVojzn+o7jdmGh
RUH2B7t5kiTB3+ns0th96yYzjmY5i3I6PA1dccsrRxxggrYHzziD4pOeXER15tp5
pNwntzU/3xpRNtlup8+oD6TkgaOH5HDhVRZhJhNN21turJHElLOdFKZxtTyF+ENo
akF/9t3vEvXHMJVAqeO+xqfp8otQFP6YiOAH8ME0mHrUIPGH0fRZT+a5erBVyxwP
bxx0e4H/+A6xlM7g8ezbpYRFjsiSd6dAEjxC+KTNwsL7SOIhPlSyT2sG28RFiQY3
rtWyGJ8KM0rMkhzkPbBVXIb5BaHwR8P3eAaB1Z0BYsNz+CUhY4Mpzgplujt1XiRX
PpXn82EJdyN6I94vaMYFxFKA5dN/CAxoUR5jiLKKB+Y+8rSS9D9d6IAaDM3X3E4G
QGbVPCy2O4twso+1RWwQnLXqMOOFFNbXjmBCPrnyF0LuyyfxUvLq19wI7gpQoWAi
l3zKq6zfCkpOEY3rqG9jC0A87v33Np5pOtgN7KdZWKOlb8kkoGH+/z+V7muKSQzh
GWrbTStjY8ZiR3UeDAN2rnjZVWQW3lMFUxxiFJXzYUCyQUm5dknLmWpZU8hdaSat
5dbe1gjamIGIi3+A9GoTE26eMde2PRzFO/6Gs1FRcAeb3EgT51pwFtMgu1ZEwpPt
R4unBDXRShPQ4/CdDyM5XrIUMdaBTsu+KMZi46lqbhuG8GbZyzVlrI8bw4mPzOq/
dcu9B4uTWbzCMbIz1I/5RtCaE7EsnIbxmVuVPVWLlOuSoAzOW6ns18MMMDr/fZEp
UHFUWuPjySWHvXC3PMYXN+/vRDNsYQqNoFYuvCvrKWwbmpDg4qfZPWRBFn1fcBuG
lHRAgF9cq10sWgF1x8xXuDoi8DvItDH/Ua8s0c7i0ozo2zNAo+/CLW5/aZCpAyZg
OouCULae4D+XWedtitcRn/zo7uskdcQ29uetepKj0QEX6Id7oq4PcstHo7qTlFBP
JyEIUckQQsGLbqzbZjZLerch77G2MgLeAp/POu46PfmW5fQZecYMk36l0VZgYW15
IaIzFPUE2aClEfLL59qgQ/UzgzfrA8CfN86S13xmeZe8M0F+gvufHPOKruI5e8Ff
+74sVxzILpRaY1zKKJbwNsRrXQ/Cz1WFo8LDPkbuB8FbvYSxms1w3cMjD9wKxvBU
ri9jvkEB2KUPaMc05UpQ5xaX8009zuBm4XbCOTf+w17rhBhAPpE8O2XdmRSfm2PP
/Jicp2bSI6nQ3mc6tsrTyRxXLOSDzTJFPMDk1ZuvSMyvjf+aqi3G9Z3nWZeGYrc/
zKOlmFqfHznPXWqlkppMuITu3GcvKZ54WQmDyPYvdWkHTAEWFVgug6rxW58BN3Ay
NSKBCryCTeTD5tElpWr5Hn15ky8IMsCTjhu0MdPRSSJ68beFadZk+GWOgHn7MRjX
oCt2nqKsifPiqe7yrYbGmAV5YAbcABykvjt+pGp2RRl2cR9dpdw3ihAgBgW/0hm+
VGXAFv541uCTdv3cDdxgIeeZh2ItpztiLVQbIC1itcAp538R3gDOxlm+tbUXTYSW
vmEzGeYwFwEJXANYSyF3Y9oVh91aitnEAYQaAZcTBBVeehwN2iPNnGydI1uWETsy
DLbhrxdSu5h+cTFZh589Spz2/aEXsqQNWgifSTnP58pQBKrgKJah5DmLOuvvz50n
bo3F/35iqyyYX9rM/loGg6llfbP9Wiopq6zXc5Y/hHBEGa7EqrOH31b+u/7jVwPC
wU6QXaKw+FlnwtTi/14LPhceszGNv6tmZQSxSRfqQOVv6/ypXnnXdrBYiHIvXeww
odwDzS50KSynOLLEDzcwpshWhQavyvODIR/suSg/39MnrJwzgUtY3qvWDM12lwRU
AGacQ1G6RfDoyDrMkHDBVlTHv1yEGlZXLIZMQR55HbQaLVm2VT2sMliVJSksl3Qy
nMRzeiTSjU/bJ9Bpt9zPK2nShDG1gI0gojRVsLhRPvvN34wKSKEGYoArlVzIbGNB
zJF+4hm0U+//ipLCT+2hc1NipeV3Pbh3FMWFigz1qDfCidKov/nlm94IQbke9nF/
RCH6ZNo2fF+eoUol5FkVujSmZ6dhTyJ5dyQ/XZpWUyuMhR/SLepwzYb1q9p0E0TH
dr0Q+3ikwNqyFI+a4mCYzpc9ACUajD77WX/AeqH4eEdF1XPoekkU03WPe7ew4V3j
59D17lq1XHfM8AhzOXY5nxn9Igb+PbW7uaBN7FyJqk/sVX5mKyratRqnyk2eMmQX
ZmLIWuq18ygBhcKudodD0FevkRYD2YmPAkxED4jqNX6FQsNg6WKS0plyW+8Ft/vV
nN0ZlJKiVNgSjwPo/FIezWMZm0WgM3tGy5EPVevln87nozT56Lsnd39IMlN983cr
hWIbShmyB2H62RiUXpcA9aBnQhctUh0+a6WZOkbC1tlQYfBKdK/beLzi4HuZsL9q
6Av6Ijrg3uSCZAkE6ilRtnRybvV0xLdF++z8+0z19Jo3LAOo8JSabIBjFRpmotwC
KDQ4fTfL1j78Wcw3VFgXorRd7qva87qFm936g2U40lYEunC2jQGkQxNh9oW+fjdt
k7TFCzo4enWIdrMpPZOD+zjHIEOFCvsYMpwzy+rAMbmkw2eeMiZ9OZZv3WjqkXj1
hnC2Wm9gARIExLSR9a7ysDcgtVUqmqIpJKMCtiPw+rKOxjMef8Xx0m+TQ+TwA/Kf
tu+onG1p7DifsGgOsR22CXMKlBgNsYC8w464OAHSh7+SpAZ/mAhS/ouu8/Z+cNF3
iQWQgRl+H2diHsEqMb/7xg1cfK7HizhS4Jr5Y0LacQYydelBqk9BCjcjH05oTm7m
k8E1HVEvT81VQQqGc5pE84lcaF8G31kiudjHFsAlObuRjlWpls4tsduOLuiQ+ytr
TK6B/Elk7SvAWK41BUxC8hIlefHe6Z0Ow0sVuYUjq0wxJ+URdYODZqNmyTAv2qkj
AoRn1Tlb6ZW/CE4gDavXBo385T1rv6FTBCDsCTUeA2WN6peSgq2NohnYtIpElfaD
l4JzzFwUAovrOR50N2xqLMv4VXkZeVrK5cliX5GkJ3rpE7hOzQ5EunncmPzqIPdf
GBU4nqcEIntmh7MhMQ+ppmL+XZQNvzHeJ8u3s/+B6CSOzCJCK6/iqEm5jzgkRODF
D2HcOdxQOFIb5yzqETQ9rwTfdPCxIZfS1lnFRtaEA4ABz8lYjKlpLvZ/vxEB1DlE
a8/tW5cBvJjAUJqEoUF50k1LE288uVZbSmfOCbRcjfdK1rbM5EzUDQZBJhQkf39m
jJSEbXHd1O4MIiTz4NRGTUNOg/s7ozgvLLTEkqpt+lom0F9XZgO39O/C5Ej2qghO
HgVdue3oZB++AuIV5xLnGCmU3BbyHWuy8rjkABEMrqTGwPjhCs+tkPewysQACMSi
/xIvmUR5OnWoGDkAgPm/+GjEa9fEnaNsxejYhh8KqeIQ6A+cOPfcDKCTPmwMqjRy
LsyouGIAOYtTAGGzNkZGQUq4qilVcNabN3GUwMm5573eeg3LycFMknbUsr7smUuD
OmfPaSVaAMJBjm4krMah2JluSknLgrb/9ANC846NC6MDEc4M2yQOQBbCFRffB4AG
H0O2CMUIMKD1sMB0wkBCa/kKf+/isM2LNxVds8WLV46SxZWAWMcBj9ybIwYP5DFI
aOxveG9UAKOOJXbeV2gntFR5fyXrqs+5ge6O3JXI9fea8b7sopN2jQDp2P1Pn9En
z4PEhyXXg/+YUxfBzNZ59O87k4P3bQ1i3NaIYK1F2ITdGhMma1s2q7uWJw6lnZDq
o6m271oKn7oXBYojI9l3+hHCl5Q3k8aUddHtA/YHuEiTWgE8cHkPZofjP4N8XbzO
zkAvTQkTqJJqNeDfHpoVy7Il7stQv4TvewyRK0NbryZ+x7w5Kh54DH3wo99sWnWC
vJ2kFKscZSqPcvkdp+x5prsapqR8TSAXh/9UWPuPSi3kArLNHJ6JKp/HHGXvTkUC
hQb49C+M0naT+lKI7IEjDBbyapg16Bt4ItJ4zM4OvbDeLvkgUlH5ZTBrhsU4k+iT
rhGEzjhLAQksYb3yIZ8W+u+W5syczbI9fBjX8VtG8ArJDRAnX0M+LnO0DZKg5bLX
5FM4rKMgdIcSmktV8yrtsC3+0hWeY9w20mB6tJ/GDUcV6z8JeUcX/VeFkSHLRGY6
lgYCgr1noNFs9mk1N1DBEf5hgaUmgu1WIeNGbWmR/TyoZagLxO4CONnAPWYCvUqw
ZG4MirisSIHj92QLs+c4VYd3Jt453QeyRfczbf+Tg4PYzhme8nuzypdi8w7apMBK
ozRAIbW2Kgrz6ZVbog4GP7aKoWJQLvxO9kRSFJuRlNLP/cKY8olJD4v7ArF2RGNJ
jyIRN6SztcUla0jIsFae1rwWcsvTki2vicLnm0rrQ+OzQLG8ka1YF8bkblaIdOpE
Za9fnyQBT9FASlDjMCiZptjvNxcTDCR2DpTZTnb8mGN0vIiQzKsi6pF2jbDqEgBl
mn0gd2NUpWJO7H/ZSIRfkth2yq+1Vx3OJoUVcabCgtcH/2KDpW35w3DuGR6OFrOQ
DYDBC8bqDaL7wMTYDWnTSQIZY0AUSYAmP9HJkXbG7rauFOqIyZg2Eh0BJvNSKgTB
JZjTcFsRjgPGB08cyZL6qLJxwJpMPYRoNDeh0OLN1kxBGOaLviNvn1u+Ss2/SlXp
oY1L3iVy0OQppXQjEa2YxfFNKNpvFwPHGpVJDcaCu1g0H/oMLmtW1Afz7NhkI0x6
nAUWP6U16Te0uveT2AlmnIAYzfATFC41opTRshZZSA5aO8iezK3h4AIX+AIwudZB
Pb4LdSRyIxySjFx+NTwE/WnydOD3krsUgPdSIEsG7soJZR7mkQY6fXOhN9/upnTg
gpx9Q/FM/q3QXaCRg61i7CEYNf6bCEUqHl2B0mtDcl+EH98poOHzZq4cgSpEzM+j
kae0qbrvfx9ExPrA2ju7F35LsqBH2zzGab7NKQBrZRpwlabkqnF0wUNtPS6+k077
HMjoqyyUu1CHIqoj0gT3SWaDh4dbnLFnfUpZeDSR78qDWMehf3YbtyBvqILfKAEQ
rtE+YvGg3NQQ4Hwm60HlL6ODfpq4kmTR7Xi3BT9S4mGulXSFomUbf+Bu73NotKmV
RBFOxZx6lfPc2fW7cNxZMvm2tljAId7SRELW1+ZoE3HELdv6Mou2UkMOcEGXLj+c
gtvgqNEV3X7EG5dM1xuUA54WvTCT9xDTqMuTyDq0W0RqQ44Uqvowyf8I8bQK3/ZY
+xs1pvI7Qi9+8Cn8QJFSjD07l7bsc2JqSb86ij7wfcpfsTxOW0oTWSBqCoPgXXp8
WZykAFhkO3fiml2mvo87HxaH49YJyohv9s3PqP8KOH0ipCz2aXJAKNaVKttlmJyc
4/j5evftVkLkIk6MMhL53Ce/uBSdWXZdG4ZfML2AC/ie768AKwHcj+7PmvNjJSQC
5BttIIeyDGJEmBqYkZ7f0zKklE9RO6SWmVZyG8h+2WJT8KFU576KmkMxDfnIUNgF
hlN8Jk4e1Kx300lMUQou5yh1SH4jjRlpr1uv5SkFtHMwKPR+A4+yH/t0dZtKYU8H
7UD7yHiw2Pjf4CCh+5q5/++cdKHphD5jqQPb0whjZn6hQx1gt1S3FotjF3Go7buy
DdKEbxiL2d70AeV+JpmrRsks6u4QXZ838P+vhha6kG19oslDBZK9Apxvg+0GnbZu
oa/u3HLuEoMAUkYrP8hXw8RYKBKxAol3hMdfFchpB6lqqHSkC0OoYO/Z7ScBUlTt
JYS32RpJ3zrpJKNYLyP4qqaEFs5Pft15kL3RliXRH2jOR1UXNO3XhqCS8bN1iVlG
Ltby4QqGGorLF1vWNvRnlbNAz5MZbtEshP0WipB2ay3Rvdd45UptE4O7XLUEZQQK
I1Xz6jSQ3cS1uqjKHL1q9bkHHGtPd55ZeWocRIM5s9FWEeuaOe/e4S/c530v79Dv
g9MSKEZJafIozDkob8j00yr76xg8LA9hAcJX999+YPnyR1mwa09rlk0Uds5k45gz
NDAh4/Iwp7tvn2rDURP1oCKsbJQ4TEmnJklEBaqDx7lBuByQLdEwNMgq0rygohBN
HCrOrefL1ddnodVK7dwFRtfYETk7xuXOSE0jkczEOvmN88LkVS/gyhT+sCFPhpFw
r7JhJnhY3GC9iSiIwAbShVvIypczL3YfBi8DkCjnYzikZ7hljt8uiOCuQCcfxr/q
06F+kKO+UlS6QA1dZoFziBedtuD2YAy5PPWIZnudl32z0OZ886J87FnA3z9ubAUX
fzzj3lhvazeJHsYgYQ/B9t6T+CMmaj4zTZkSyI8RaoS7/6V4tMPe4m+JRK9amwzs
NCwLTZpxpDNjkYJoz82+AicMIyp61lB7skpevnRYolYKACePNAYSYf98XiBW4a5D
y440Y9fsyc6MqAogN1mMqbF8fZJwnG75+w3Ny4Tf4qHv97DOXKdwNotVuaCx+WgV
310+RecUBgKaQDKHAg4wSWx5zPuAWGjLtnBPQbb6Z07i3WdGmFgZTR+AJ6+MtiJS
HDikx0CLGyicQjHRC/BZfcEC9iU+wtF2d4tqE5eCDjsvtX8FC/tfV6c2EaQHHvcn
Tuck0ohxOhCS0Q/5nDvll3CGgE961z+6T5YkuRHdwhyAO4JN28jmNFWalaubh+N6
YC/VbuIR4aLYyIpL4vmDogLONraPO2P0BqZDbbd1xLeRbPh+Nyc0VDDZS1hnsO+t
OoLuEkIbH4aW0TVdShW15TJlS6VzmlOvfgkEDf881MyCWJAj5nrh2gl+n9J/H+oa
ZdBaMJNVsaBqcSscmpICRiBQBAFb1b2ObqJ9L676l6ZmjcyYax+oh6Y1Qiq4w+CZ
rxXH3noOwCrVFRgStKFTi/hA4Q/aN6RSKNM6TpI1i5JmxAs2maeodY95Cl1Z5ptG
HTWLq7cy4tYtGY6Na/5ZQFUPRucHuYpOvTbfyD0WbDw0BPPtZE+99zJZAUPMmslR
2PEeLtGgD4iAlxPkgwCXNjuNM8D3TYAIch1E/4QU1UvT7uCK1+SpQMMiNxwFQHc4
jBct8QBOq0NBeZl9pdfnPAFuD6j9zSnVpjY7Tp+J+KoEZlMlCvAIEwc4sRsFXX0i
eQC35R6cTzeSjlH8AB0M9oFqGndL3aZbtE9sjZyGoKgAbgnqsSWmsQDqjW7+2CCX
Z2YlqvRDxBYTAoqNuzPBiK6Yt/c4b6b9EACfbPecsEf/P82O1mxprMSpsBoPcnvY
E7fXv9KZdX5/BtSS3H4JIPqY+kq+StmSHrdrEivtNOM620lAFn0qQfsgGV/+s2Tj
vwkXhbOXO0Yp4g8dIM454ze7G5jSJQ5JjL1oj6i62vSue9QRvSJ+2H4zkSoQvPMA
ra2/2agivU/+TyEPfQwoaBbOGzvTZO1AQk65S1NojWni7Qzm75tOl9x4Xw43IU/i
pIaGS2k8U1TurUFtY+r0h0Dj2Tilr80pBqL6SQjMC/S9gDpNSu4soWagltFUh1CX
uPXL14WcSgSFF4zKZ9YwPNkLYqftnDLWD7UB07r5JtVdFyERKEbBy4Wt9tA8T/Om
aJGzABVvM78XFnfv436UhiD9dIFZkNPV+utbH3oppRzDj/4cE6aNSPHsnlA7vS/p
bRoCcztx4dK8KvHM7MNwfiNB0/UgHAyCcYg/OzZEAhI3ydge/pivX16xWjbmxocg
vRho29XxI+scaUn+t86arJl+r5J8w/J5FWFFm4W2vnE7W0pCy2zUpHR0XoyuY5Zd
cevpHe/EjwSMyZI/E+FtCV11HmTE2chMIevhEiKNycPLOXshJ3rjbmztVy1chTrT
HS2X0WwLzCvUhtPfJoccg48n+URfs0DggwcF18+uQ3yNbaal/U7n+ZWHkZqizX7w
uD5HSRUnSV7L7vJIgmXKSuLo0R7scNzEupGHpg9in9WIfeypjBIezpv8QtTxt++E
kn7XSOyoXHa+xtLnvNwk4I2aCa2+Q1eUuwMqAFm0jkHmnxz6RRekBJ/+8iYGoLn/
EzS70A2sXYalNjfGWMlTbP4gwFy2dXU2XwUchjEVzfDMkr6CAfo+Dw5WmRfapAZf
WCU7/LCD2RnUdKxDDDav8KNYD2D886PAgYnt28alR4EOHnsynBcwTrfiOGeU9jOj
GxlLTJmzn6tIBfyQ+6ggTtTQejN6X/WHFmeejR44i390NYwkyQHx+A0ay0FWEpfc
qwq9UOMPOp63wBYyNB29JZDSCfUFYrE/6ARW4g3cCpM8WcfwDvg7pHJCFcZPu8/n
GDDe59viz5eGkHTOS436nB3el0a2xhkKzEAOmndReKnWx8YeygzR6LsCNXvSD/FY
v0OutKnaPuL8uRg2jiKYOf9OI4UdJ/6hhpFmTSi5772d1VxOWvb7qdLOtOJvXTL4
+s7nl8thM34qeU/bgqZ7Sprj+SW1CD2SulzIZi6JNU8sbULVOlR8sopSmNRzmdTv
NByOM4pqL2z+7FmYsiDHtz0NVHOn6DQussnEfXurFIqt+LIQ3lbnJRpT7pah9nSo
cxU6GSU39V9WUJyLi0TbarVAdeWxdMcHJkpI52hAxwyQKqeAHCYnwwEg3UsWYCs+
GwRxEBG6ylgAqP/BRAcNrKF/wfZ+0kicSqT8rHqtIfBL1GNrZnktb9sWuAMxKd5Y
CNi+2B1Dbs7a+kzrgX/zm5g08Ysh5FVH4YBFN/9NgjN90MYlyN4f3KW0958Pr/7J
U9Ht2X8G5RMttcWHyH3Pt46o5qJ157EQpH48uOb9hMaYzNsg44PusuTHYq9VXRta
re8qjrlCq6dguKGHcuwxUrWHqSN+xHNhNR+6g/9qyX+r9+tBDup5ZU8f2xZbV46D
NMwUWsohxchKLKfC/WhZGJj9cRVdomD0OjPWJnz8tYexyHMdcqvxL0s0LDaa6CBl
B7eX7uADe0p4efguWwkmTuuAcyOy4WycdNqBEBWknzemAIeyfaBZe6pF9lEVKrNk
w6EFJOeX3OXnfEcFF/phaAxN1BCarDRs6KOurwb5xDoV9C/c8frcJ/Welv4IUjVL
AcutdAZ+o6TgD4Phfis7QLVRPU6kyb0oUl5kAnI5A2q47/AcU2CD34MxusyTyHYM
qz+pbj7X+6Go88qf/C4a3ZenT40tnL7Jyx2eMljpVYCX5lXIwjHAX0FTdOWHpy1v
VnsZ/FpwXYbtfdl8YmigKXERvgXNKY6ffRFo8uYbv5xLmRflREpFevDb0MNTyUBm
vAo8ZWwqfEOPNlhYf6H53eva6v5+EkaYYXZjTo7aWdeADuJbYxh9/h8d1SPa9S9y
NJj82cMLTY5F9oBYsA7MJM9UL4CyonlH/6jjqAcrgtXHUmNwKYVuRYdbO6mRFEoy
qD0C11iOoeuOoBOF1wL943hbAqidAn2O/7lPJ1aWwKe3u+6/RCuy3bKIACMzWSvt
KwACD9fG5nAGBI2E0Mzk/19i4hKEBpuIorayBPlZY5tAEDlxOpTczyWWLskAto8r
JXtsAZ4QyhjWBSrCNuefwQVN0pUYdROunvN8M2cMg/6MRn21dGJt1znpTg6rMWAa
Sf98l+RspenWomLblO2S1uCust5S9hYsilbgiZmlofBWj0h1Uj72AVYUFho0izfO
tU11C48XsIqFA12fSiJAfA6nmmNrQyVNZujVQJJEPpRGIGElqQq6tEo0VCHiLfro
UboQCn7rWkib72Ti5BGOwf+ntoy1FJTDW4RFUy7kgJV1hvSb41JmqphdOp8rklcM
F0mt0SBokyiMZUO4dhqKw/qRuupIAG/bUcgJZnJ+AaDI8CXvVpS94queP47QzTmQ
tl8/a3Fen0V17SP4gFfA3kYqbNqvf9nLN5ahTpRwX8JXX6jJqf6m8xN8oDjDc4zl
AAEcsWrFaMg6pbhTfxXmunY4iotX43duK3gr5xFPRa2BQDOxq6//nas4dQ9IO/Fe
FKBXJXFU2CXU0qNoivePgPNiC2DjxGkDwWGumSFZ1ujpoq2j7No3QIsFXe0UFe9A
WAQ6RGT4mq92PoPmchMU8pvnyaUKwy+LOkMIlrDnsozG5DvdxafjI1ApCB36NtQR
OLsGr5wsSaETgT6I+wul0PbJPc4vAxt7ioRt4RJv+NhhNhZwNXfKJqr1ee+rMpiw
JqSufVghK5cX252o0TNHP0wD4/ieip+bUTxTt2KSkVYNovmFw4ZrDGxWK7QVemlI
Wi64a+B7B6nUHfySWY2qNuHdjhmeS8uiVJbs6YkV19p45MMT67IGgix4O3P2/2kT
YJzGYhUaPpHxnWOMAg6R/IaNebos5q+GCc3sbwUjrDoJfcsAjEm/MjGWpmVH1DqQ
4Ar4cVPad8WhJ8NGRKre8UkT4kK2ZwWus5IzEgXva3qliAuV4aQ6lH3nkYH3P1ZM
guvSOK4gmBbEtfcVdk4MJA6guTM2Js2i9Wnn2J1gihN16ItxBcK06Xmk4bUjcfJP
gjUtC/YtECuIn70oebWEkHajbwRwA9pmpWCUualrNo16jhxClQ8AcCM6z+fZfdjz
hqXEglQlh2esvBLucPe9jEmg8feSD3ImFcuLJ0yV3YGu2PSAXs3n+9JRmBvkO8/R
eTBkdwA89mTws6QMEthGQlbswhX9pdv7RqwBQlwYZB2/+I2FUUvVKbH/1h9F4xio
5wiorcToN6BWz9C6U6LDIJYTx7do+V00e3M3AbGe9sXvebpDxqq4xc+NOZ9/TdqW
/us1ZJsXgZ2McCz20hO3ZVIHAADZy467G7+5/CtORusC3dMCZQ90qpOIfadKE7sr
fbVG5MSWh0Fhor4cNSVHziIFUC9mgOyomK7Av67rWxs4Zf3WwnTtRfYz7YU6TBAr
DBFvXz7nbIMj6Ry+WrZSpCFTKOpuvaUPnjfZows591IBcYZ+/To5//tkrD9SW977
KTy12DOkKQn6+gXbTfc6sczMn6NjxXdJHIUrWOqoGVyqODNbQDqxlxibHNWWPVqQ
x8PBJEEpXXkV/YnoITzvwn6X5hsMwbTSyitdtCCXAMuH+hbmENUNUNyNgGm3KTGS
PQNmxN5mV/7bUzwZJaUIJtP1kW1vR8WvHXAPTFHlRS0Nl7j4r2KOaAU7R6sAUiMO
UZh0LmQvt0RM8em/TvBTlYSrVSTai5yM/mxvUXYO1qvzOTFlOfZoRGGBVO89UNFj
eW9iW1JSe1gHMXfMRAthK0y9rRCqjjtOSF31NVH+HakMWg4EGwnrXjsPJ+cMzGtU
0N5/xbsbhptKkvn0xhQxI41cIIurC47NAbiA8kfbz1ZmcCdFPQioBgetzi9a7oBI
Fnz5p1sJvtpZQpk3v058YuSsMLrRwWy2dUeEDSm8q7uPpgjJCUTgJPFILqBZKsWZ
v1XyGq9RIrQ00enfja/ipaWb+yNA7NAL8suLsUptN7OVlnY79tecLofptSCMnuFb
Qt7ljlQS3wUePOAFKe2pEr4wHdu3vU9mWRwFYIdmXgrlc7HUYuh4uEZf0PJ0eGy4
f2O/dKBO4I4mxhRkH/V0JZNLYaC7/OWUBX0ePsUsS8yHeMiiHkyEkjuqDIUxRFal
yR9j+JMYsuTXSqi+FKEsHp92NePjrTs/ccfOlkHVI3faeRJ503uFaRUrff+Mjq+t
872024DL7SauPN3Mew+m9eu2Itb35b4jhj++LVzAXyeMpPK9P5OvE0z9qvU0IXZ/
leghfckJwoFCYixhTLg5eXO6MkVb1KQPNbLLALJyrBvf0cuDFSKaQ1aDEZDZJUbq
QmS4hdAqpVrlfte9ar0oAKJ/BY15QapdJgVLfg+9jMrYQUOGRY6gUWbtTZPTwR2c
bAsMZkI5gS/1jLG7DW96dpWgOP1PGxTInfjNXia9QWaPZJTRuYNfe2uU9UA2GfAI
1OwgBwIRutMqNZ5cUoIGvSWOIohciazB9MbnrXAHnhebTIQL7xFQNGzmeond23Qc
FNk+sTcnk5MRqJM1P+lZB6OoDsk3cXoX0S1AWCvx1q8jmPaglpyQFfR8vQq5kany
n35wWa5ab9fV3fLapATy3ul3biMNwzZ4RMCKGUJwAYA4094ZOyzldAOXs/az5N9L
YKS6mNXFJ+0kelR3wVMJmGgy8mOx9YVZBG6zVVwSXqKe1I2SUytcX8uw4VQTSCh1
QdJ0/IolIHsp4tjX3Ml8A0EGT3XW/JUxlF55GOjpHBkk11zMVav3t7CBgDIBzhms
b8lZKbkpLBr5fxjKKTWiVFEaZjzuFj3Yfu9Mcf09W2b8mSN3IyN5dTvMeBTf+zVF
L1L9dRS9o27WEfoO6Mkk4S2qEpriwCzyfBGnD4l1Ug/PZiUKZi20wTK66kl1aokN
ofTCoUnVpEeeLFnfZXfz5H0V7EYwwHWNZlOFDnh0mAE92+NPYR0cfVhiczWjcyav
LFbZDQzWdAGKjbGWkMKJZyw/3m06qN/EWkbHnMySf2EspnPVYPRTyCRChVLu4Qw2
Bryn7IKcunaKtmxvyhXD7uzy5xR+UGoErZTrsK1sa0D9wPKym7ggbrqeN+00rF+P
wW68vVuovDxDLCvdT+w6n1Whsw5YihcXfKjwTV2Qy+r2Zj4XGU7VmPs6ecao4eo6
9sFfhgMAsp6YMpEk1+ox/7AsgxcL8p8EpjETiAwvE46ioW5QcAvs5kUTgOQIjAmk
8blVpFgjcmax3cSr8Ksgx75U/8iWC/Wx2yN2LiCO4k1x2644TVCC8c0wHwT8pm2f
5rC1VWIpkpxQzcrhpQHC9CHf00uu96ivDUIi6a/qhjekauas3megA9EM3rAPnZBN
m9qEKq7vcTPg9+hUDoTdc4islgzHYI/aq5pSLoWptv188/lld2dDltFPKAWThJ6G
JEtBe0tchTyMEIPouyL6DsNXpCVKPsRwzRHqeqtM52khvh9gSooMBRh/O0kAXk9J
iZ73E+1MhkO2baj1ln/kIQ4sBEHuDAaDoRiEC7bhQrMTjXMk1VWg/ttBFrHnMoK7
4oeaZZAPv6soVWMrsInK4kt36PPv6rHBLRb0Y2tOHV2qSwAWzr1e+YWfwYP/IHxv
pRHChSZqCy48ZbaPUl04yBMqNxCkdMsX2hpAi2lkU9jzszVtv9XVQBAv6K1/s5J+
ZV/9KJfMpdx8HWFScWlhR/T9Q5slI3wKXvfzED6tLpAIdDZSUv/RsUXhGEGnH/Ew
XJqjswUdyp6GVZxKksmgRBPeZIrDub3qbP4NL/F9EDZJtF4fS4uzVmGJoVlb0hSb
O9gtPatNGPqW0mBHOTth7tiZ8MYN89BGKpIwv17Wgz2HnbXRHly4uiWxK+G4G/kk
fqq89ywe7TL+F0ZKUasaSWVa1zkQfUH6UmGNFl8KPWkSZJdZu0K6zLAMOzRYBQ3j
rpn+cor7AyVy8iObTYIe8KTT88hYfU7llmSdHjo9F9G3KN5VSUKmMnSNogfWKtSm
GRxz0Nln3H82+eHW6dM+C2VduDDgaJ40f8WXMC76BFp9GyhXqyLChvxQ9HcK7Xu4
FtNlt8Tr1+HaDxnXpLhBpGIJVNnewxX9AlJeIYXqqz2kSk6g9vKkcgVwZ4eAu7m9
zGW1BeYNU4Ds71OFmByHLMx8kbmv/q0opQra9OlrkGzmfwIZi+6a5Glxou1ELqPl
m8oXwHckFDZkm9Dszck1fTotAt2SFYj3CJx2L6vdnS2dC+ZKA7XN5sLOZCIrXLVA
YJogQkNeib0LDo1pELMO6csgKXqboUcC3M7SCiBa+hK43KGjUbaRUQhE4TyKURzs
FLq0U8pEnVp9fO8akHRxRgIap1xBGnkWI7PpBKufxL9y9m0amELe2OGRbQxZTlzJ
Y7Zn/sNnPCTuhuutdqLHeHVEhlp1dloQpAXY8Av8IFAPsq2tLwE5tK2pLeZdqqeF
Cdq1MVyTPkslfRl58h4lLx3zZMq1AG62dF90ej5tFZYa2J0JbtjvRwihjmYHeRoE
7mBRSkDQc2kuyE+hpWS309QWrlZ2lmf1MHPY96umWHuYpoMI3JavxUuGl1AZ9lCm
bbGs3S2pp8sDyC6l9qYndQ6G1Lz/tLGzbo0+/52aj5Qxdv/J42EkXnLAJMpV6eT8
wB/p1O2aSmVx55p9yEZ8H+gbJWedRUa3UJcyhl86dlf78U4m7EQlJRA0NKrf63GK
CrxSSImpZG3HgpcXCxFbmVplS9P59fI67o4oUMRffaykpcMw4rlL2txn+ADlDlwK
W+pqY7CxfgzSrAAA1iFES4TyhYax7pVkxFMCmA6h3UqRl6Q+PardGgbHBBn3loON
PIPTlYzNKHJV0u73Q6REdi3bXdMLKBGkSC//draZMWi0l2T1tmKLlbG6gHswbOOu
8VhB8PGIwCQLVOHjvdI4WUEA21+DUG4E9LakBBPR14UMW8qTTCp+Z+DbtUBg+7xm
R6IIZ4ACyrvPJJMk5na0kcLE0EqHlGBccdpFGRJNKRP+rUMlVwV0azjwAtTvE3Q7
RvpcJTQs+lhp11MU5JUpiSmWfFeCdMr8DlsGXK1/TeYEf3L7/+VH16HUXmKW7Ldc
TLoRmETlK2C5nHk11iXWCoPE7DULanOO9wwhyHCXdRVRf7gkpxe46fFn6vzsrene
Tq/pPWrSlAf8z4IX/tu9hj378xwir9DNZqO1Evwb4cFIhVseMrAJK068zM78hmPP
EHj6aIQOHADXLcKZbBzBl/i8QpbEWGRCyM02ojZ3v63kFGktG2nnoBScs3b+KLhW
gube9y/1PpuCZ6ZGCCwJX44Wcs0uY0iq2XvgNOZ996zPYgOXfluam8uqPMJAaUfp
xRysKRQ4IECU+w2LR+WTs8uH4h3L+lxsoQZBRZhDk0wR0+LfOQrkKE+2q+X77QHA
yLIlzwAyI7gFObD6o52wHtBJNnAqRvVrJKXkMnR9TH+zhAONPxIThn0Rf+uDnG6T
nESPpKg4tD+LUN8kZk10NQlJVhuqD9ChAQmVVm2/Tq7JhL5loa7IHvJ7yDVHCPS1
Ns4C2Z8d68nlQL4WrZD1WG5TWeFdZgsasA8Ax3aD8J6SgewlvB8M53IAIP4BfwKE
+VmqqbidfoCId7una/uKA4Ki9JrojD9uj4u/O4y0IRcvVxIvJQKdrfE8gSjLFfaK
IG3ArU737fMB06FQfIlxvLw2A77ajago8ahrOIQau6ru8WHJVLfmxd9XLmg7HqSv
/9Gnnn0Re+4b7wLinHwt+rqAprZl/3vZoHPXhhdhUjN7bEjHoB41oZqgSNllJcnv
xgnl5YYjcZ4BOyAyTdAugO3zWb5W+vPxk9v78tiwjA2IykcWlmybur1dOZK/q7NF
ohchMyZ8vid0806DTn3I5me5ZUIqRZh7olJt7wN6vW7CV/eTQaT3XCCDmCGoUQDC
aZZOmOuNqQAKF7e8q3Z2Bs+f+UInMgVk3rhKWq8Z+tf5P3aZEcmdrD6vtjlihz6m
AhNyuvvLoq+qjg5QiZ7SQ2FVKxcBGU+gpixMP0sTgcYQhDBuzmRXm/TmQrMGHYnS
PY7wJzEWli3myDZWi1TvjSGVtrblPcvJ2XR+3/RnXxA9Afe9VQP7LjRyb9/ekKHF
T7U9fbASRfDd+rjgrcQvTOsU57uBdPw7LTtg5v5NLVZkhYXWFOFUeAOYNx0J6HoK
GLl6wuotiMg4kPyvCrQJdgoZIL6kyI7yowCXSZknT+hih0+5iOtxHP+uRcjhL6rS
KPcCTDbMkf/Is8DwIdJzBjBGDvXmhakB0YCe7GBbac9rPHMQx9yo3m/TNvT+hx5/
aALU7nbCYo2czbZ9LkS0/jk/Tn4xvmCcAN0UqMMCdoGdTUmpoqT/LViGwdNRzczS
0DBBNuJ4LjhB/q5csXjuoa+9Q5cPbeE6dLUubThZFngHk3omxSy/bdIvIWy5jxhe
ADwytC2bi5dsp0/hx8SQTzfFAr48xB3hIvolWfO2A4abvEV/t4faAli6Suj1yW3A
AfZYA6i7BKLZmY7r5oLLlkqN9F40uFxHVa7nHDX4NHmeV89w8pc/hUjmh03c9cNy
63V9Qzww+96Vy7NJlStcXt3srWzCeIu56RdFq1Tq/Vm4Fl/FDemXY6kpNoDx/IwK
Nma2e7MddV7RQK4dL4bBaha5iQ7GijLm5Yl2+7WY/ezVgj1s0Yr8h7TC+dYPqXmV
3+ESgIbO354gnlnd5FhsTQoixIKGB+xzMV8Q+jtfMNalY0VXm7mEdj7UU+wW/m+4
keHQwvbp3ZjmxqJ483RSgWrbuGsk+doB8gtRSA1nx30KC0rAZdWvTH3hqcD39i0u
TYg/BHtRHMV87biUvcqDiDB9Chmgodevq9d9GitsDO6j5HH4pe1esf1nFhh66kh1
HU8Q2UWr36nrvcwpOkzIbw06AeEA8Kz2aJ8k9kG53+ANCLnfH1fqby525u4A9daC
M1Ltff7T/yP2EVrhVMBa7ypJhjT7GG31xfG+EHwnt5x+exc/PsmF2aFswbkL7OGP
lvM46wSQrV3yYgWRlZjD0cpX34joIXNcDvd6oVpzrM/KWeEkYacqeRyi9tbQQ6vm
xfHLNfY9f6QNWU1v2jGYTRGpCI5W6nVDULTenNJsXX1wcx5HurPQU9288cCeWriG
E+vu+kdWANVtHxgrUtzq5cqS+Q0TYV6hX+MsWD6+r8St5U7t8PANiDLxIlcW5/sA
KKHwVm37jO+bJwuJ8lXjlX91yNrys0Dx2xroYx0UYeSfCqQhFza12OfP1BiPf/1Q
m7eSCQzq9gY/rkAuJR+/ieEi7mEzuKmp0Bl3rMM2Jq7bTv0VubuIfjrCjhCqzbOv
+5967wFv51yOiJVk2AbCJN1xJtGdI8z4PU2i18il6RgLD4AfARSxJVJYJB4uTOLm
MmYintW2dstl6kIFJlJd2Re6DtFYOJsOUp0nr9cUAZ4W/gkJZqRPF4RQs/FH+Wfi
XtarrmGawxJvNkXxDLk8uG2vW0KK2AQ3TSvI4ekzu1SlEuiPjipl2TaqNwnzJtvM
hMvge+VAmxUP2y+M48ISycUOZ8errtemUNo//xVbcNQpoCReQxzGEXNXtBDKn9AI
oz0dnp4pXgt1iRYsC9DhRwx9yvCzVyhIOxXOTh7/skVSMscPzsmK9qPSicXL7wZr
PKqOW2/xadheKNA4dFzZVnFys8Im/hqH2d6iDju1b49iNhonqLwT7t2c0/uDvpZN
ZtFmwkV0IT6UO2pDLYz0HO7289/rPRC9lya24iU1RKP+dB+TK14q/068Z0JUBJxK
HM8zcNuuwSNBx/e6WcyStQsXX6vJLgvx/2yPrFDmR5WkVeBkONNvswQLU3YkQ8ib
3RRNIopDZb/uyhHptzSAjJphz1lTveGzJ8pL7ad4zlQTv6zLDw2SQbcQ+7GXvS7n
QuBLF82vJQa+HgxsL2BqkclRA8DMGw8EqLbDeACgLU1pCs2XxU7UmQYALoN6LInz
rQOZ2nXmwBYTlB2nUnvkWhSNtXygXpzT+uRK6bx34041CPpa51WtXzm8CdgeEpxa
WeVDIE/5aNPxuL7jqAPjrAALn056i4PFXWI9xmifZUqBuiixYlUr86BJgCYOBx1o
97YeVIkVMU2wtxgdOSSO88/JApoCOH/AGRQWE15YfYR+ZOUvCatvl6GbsasQ3vsR
Hc6YPFvxmDW+h5cRS6ZH/1C+XbAS3WW85BkKwSmf2EdkAUbFGM7n0EB9/nrBi6mU
adl62YK/gQNhv+yxQQpWUHHQWNhxLzzpTd+wn3ZkmOYjMLfTwHtj/e1I/gFN2BP7
ISDZ9DAvViQqkqf9HfD90J1G/Abr2yAlR2Qh71gLuoYcaVOjUKWlju3cfz2eTSXQ
PlfiQUzHkKouDrWRUYQKwnnB5xHI/+MgOSUEIVqzcz76i3B5BP1c4qim76I+Std3
IWOaYSPl/KveUGzybPLPFUixpYg0pZT31qWAgxsTyTmyU6kFKdk2X+Qa2B6nAvOF
Z2iAHoClQ9lDKhCmlOaldG2iyXw5V+6rw7BygpuBRVJFO1Rhx1Cm5CEuxE8/nn26
3fUJLa36eblGHEUfCf+p+acyX8kDFX9siTPZuoYdLhBNL0e6S1d8SCHCnXYetmEP
YznBuRfa6R2OTbsVji0snOIW5Gb/J9jQFGfWkLcspW1BawDAifVICPvf/y5TkP85
dzV2krG3m8VJyQEE2CBY28AJ2/muPsk9Fmi+PTtYV2IAb2DjeLQ6T9jfUzMb2o1d
LnJf+12pT/yPLMRvdDlRVCk9FBn3WkQ3+kbbRhioHH7aKdcYDJAuZLt4nCzukiSE
quvp8AZNcLJFkiA+uAXF8XuF25z7jJKTIaokk6RGUQVU9VxBRMpxdDGji3NuQEhQ
BkytTqJdNZqFhuQNAoaKfOEh0SRATTxPp/CWcpTtNk1u0hidsp2/JS2QEDSNGPrR
884BI5MPkkXI2B6NypX2zH9piHNFmhU9HvSjI8d0CQ2nPNtYiXAQKOohYdmVaaVn
NGnGN6MDnOYamVQNyKQ9EAhrsKgHQIgOcbsrclgoU1cYO84/2w+Y+5irsvGilwQP
CPjdbkhjars3+92QbH89Vg9EKec6IiQ9qrqZK9SpfLzyosFeXv3hF0rY2NivhD+W
6QNppBi/Nh/oM67Bh2b7rTTNsd2x6oSG1RDVHqcWw5sHejvFlfl3S6DJNk+QNwO7
FXWx8wSvWzRihhqfRRddAZcCd71qYyhQM5n+IE03XbnpmcVyD+jOeR40efPL/DXQ
SAdqgnkIYhtRKewGMG0fmW7f0IPmTY7ojM2KbQSAHZfcd3j4Sl5xCDqEn+419dcZ
qmSy/I4l7bTebX52ytk6uE2DByUIyPuYn9ZvSUJS1Jbu5OPSjZ7P9nSf1M8pYLVy
Tzp9b9oXU4hEQZN9BfPCGk9i9e8TLALpPPg9ER0A7j+qY9UGTJ1MywDK2Y2dJmst
8rSLwGfiTYKndOIj8qnEdnE0+Ta5B56FgAf2Zx7clBcbld+9KifK1ACvgT3awI7W
xOSBKa/ruFmHLq7mqntknQeXMwZbjjESHOiqcPQ9sZYqYuL81mId77QsvSlKUrL3
hh6FNAJT5NUmPZAstSvNfL6J1vq80AiPSY2nvDVVCSJmCoyZQmNb3yE5p/xBZ70o
46QHzlRli9wwtY39ZdPCQxBXW1zoRQGWf37hVK8GlBN3/A+4Y6pPASpl47Pytedk
91gdmz3DzU+7LtmGS9/sN4ajR2RXacVTZs+pJWe916VgyTJjDDp6SqbdS8vjD5xW
zVgz1vCjTboRmOgr0PUGqJmDExrE0mlteilBhe2FLC0CdFNbRdTR8kKm4VCiuXgq
C/72mgmcU3AGnQGbS3kKxu+9Ukp8jjUlATlCGu8aU6CwswYXF59T36SwOgdu5yGb
NGdkwlBei80rWJn3WMdkZjvdx75GSEWyTThADWL0Ty7bHlPjw0F6P4ji1ZPl7IAD
CaumAjnP7oi7CRfvb117X7aAtQtkBFWFOS3I3WXTHs3dFVwWEIEtCCEB3UfI92uK
g5EylqB2+dYsG41MS4b3qD+WVIKMM/yVSs4ziq1bMxFQ/UiqLXkv/vRHoSNTHZi8
uqXW40cMHO73DKpSWmexME3OF9COzJ79e8/BPu/3ZtDNyBm3ZpSyH8hF97Gd8WZo
cXplXqPzGKHHrZs5UwJd4HIR/k4X2Ta6sX/99Ldu0LNmd83csP++ogYkP+hCFyVZ
NK+ESThI67XR1SULXCRq5VrFSGjnKV1E7EECIPWToBN5SRwMEC25Hiz+i+iBB7wX
ZKDBV1k23kUC6DhCFvnry3IqzaeUHy77c2DJnolwuY8GBYOXfpetcwo4Cm7YFXY7
s7fwSS6BE4lbXhHhV/wVKRJ+5bFCPA38ybGO3MPAiTykgphxOrrMPyUVQbI7nbwm
3ZcvN6M9XRSPVNrLLOPltbRTCDU8toJzc3bhuy/c03zuqivN1yyno3TceqpL/KSm
OtZEpUn/WJwVaPNylCR/oPPt+er/mUffH/ZRvcBQA+nvpEZC4gOzRsMjAFgeSxzz
BEyee7tyNN58RejDmBdAgkS5qxtp7pItz6qPGU385ZVGqaieJ5buXl87Azs7FaFY
oCzg0K63EOV1CDA9RTdTlXrZySY+G2xpR34G1Ej9adaUedvH9gXtXQODHc9f/2QW
xaD+jIHtNloJ050cGYgjgLdIl9jUtRa6TA0ukF2oLpRdOlvY2pzJE6sEIVT2SN2K
gE2jSbZv+2+67WTPr4xTBYbUmeb9K+blRkp56BvskchdxCyCCDrnZSflz1BEeaeq
Xopuj1vkRfp2vlRq73zNnh5B9vyKjTWFBXdc3Pj/TAckRpB8bChL366w48s0qmNh
VGNBX1PRRnRVbWFEeCKkfr5MopK+LKgOcDfVD+ufLPd+uvXVvS2wENwhojuUZQU/
8ilui7HLXRWMckU0KlnPD276GxWOtQaSwaL4QQkp1uBqz7Hvd/H8If0FRvgsPXwD
FrhCVyjsu0n9kxTp/c2NP6UXNwiR1rvvDIzRc9u1PDgaBbCR5BF8K6kd6Grw5oX9
q7omDF+58BNQgArB+bnWdTIo6xrT4nDh1puh1iNSydHA4irqsZaJLQbZVui6JEiq
Sk5TSMf/0uM7QdwUmABvPm6eRglNuz2Pby3+BDWxWHh+jkHx9Mwwp/Sg3W7l/zhE
haGu+Avop/0clQzK53ARV5OZ6z0rv6gFnDw0RkcW9uvOvE94pSaKD5MJdm1wn+CC
EgEQobyoPz/KGZr2Z5cBgwOE0HqzAGqrf5JTO8ZxX/+4XY+NTApzJ+wJs3fkP3WE
B4MpjQHa+LRtj9fKeLSNkaNH5rsb4gUR8n9LU+Q0wB5p49XuHX2QG3dsq1YR23Ih
vgjnXuPzbx56LGHpFHOxxCkBAD684h3/MEfg9KKSQM8w7Lm6cDqbKCDu4fvWPo3N
k3qWTIHuqCL+8FNypWkucVZJjrIvBdMrhoM3+aTJZDEJgPRz9rVzhOczY6Zac3JE
9R2G2Bo6ROJ3NTPw22QrsTbnrDmgoLIxfHdeLdnHi3ma+VhzZAhnvx5NkmcwK/95
nbpFnWWZYeiCphZASXhF1IZwbnzy81YJmjP1OZKGHqnXU4Dbp6oqU2FoK8fgt+3/
TuVjniSLQ0qF7pY9ySNAbpdviQbS0CjDK4QM6BQpCLooLAMnPrGmtcBmN+iGbwxX
OPTU0sd0SzPf5dRCsi2hb4/rKp18Fhho6b/Wv6lfof7P6ain7oCmpPg4vx85ZQ2M
5hFiSJmNhqemuNhFC7lQnzRc5B4awm+0XI6Q6ve+BDztyA7zp4tTUrsSrxtFYowb
wO0Gy+3qYMXCbxnmi+Pb7w3ceZ98zGfKSc6glUwtx70ULbsbovkT56THgIdtaczc
kTn9WcIiIC4a/alvFkOgAZSZuOJxd70CXSw2d8wq9p5oE5GXKzOWFI5uySwKerdB
tvS6OmtR7INY8LRuMxXdSTyH4a22RbnuLMiSQWiv7o77l+Neqkd1riYEmvFWi08I
tdwvytHM3xlXnv3sx8Wd4zBglEj2vpm0b6nQ2nTMGcYUQGyW3mAHuh8w1e8P+Hcv
9EgMDKaLafBVMwLmLyVQBtm5WJoG10zfjIORHG87Y4ptL6SV8+84BNSCKrkMRlCm
DkOzcE4gC8z5JUW8UhDRmrOmYEQxZQmOEPrsvBrhDn5GKVbiYguOraduKAAH0Sev
GD9Q2sEE3hZ8bohsyz+PdALBwUisI01FXPu2qFX9NkcWT1pOBaViLlMrc1yMpELz
enGQwF6N4K+YD1mfuoSuBzRwwjoxzB0Dw3t6eU+Vif28ohlVBGuxhJd0eQWncxB7
/mxAkSKOpWozs4uZH9NCsPzIVfmDkPFj7VWmswYrWnFYPIGnEa4LeAi9FUH3LRqM
US7lJoE6/aLJ571P8YwH+f6w3uu949ppUT/zhVA/PAgI1t28O6e+9OOto0+Yn5uo
JhtVQfMOVebP3SNk6QSTSRYJZfp0/XFFo6SmKucuMBb6VpxeutKvbXSphBrYPV1x
o6lzdc6RX62P8+lzVDNLPTs5Dfw+ruK1Z7tC0hYYK1xWvFsHDf98G8lHahMJgKRj
o8vrFiL3Xk+NnJgHGfKWrgJryFLzPuHMaVNQ+xtEeYwYQTZvXhkCES3XvAEzWf1o
DZ4LpSQpVih9Huky+PuGPS5lpnU42uCLSiLhuegTDz0tDvSObom9upvM8D570Prf
k9dyBCSHr5PC5yY1HiOTzmq7vXtnlLieYfSF01VdFcGO8/PY0sNRyLBcJgHCQQkC
biBoahNimpyWgXHEQUEDf9Rne2ztBPYtWH9lYpjp/FTT3TJFuW8F1MpvIriMWagv
z04GpZB2hvVKHsp3Zi+DkFV/SNsEMwt58AfUeggpVyrryHT5AyLlAKLd09Uk/R4J
FP/PDX7n4blqeg74OpRO/JHlLEDFvewGrxfi1xjANHXNgOikUhZHCww1COhoxXxv
B1hXArK1fPjh/Wa4qiRkeImjqJb70L1kVbpNxoyzJ5TSI/SRsNRiRIyQEzaggq1n
1jn1Zm0KGWAHP1Q6hWUAyJjbkGPVfPSktRaTPK0fqmHF7d7J5JUVbOT9mKDbVYdc
ylkHOm29vmC13RX5ka46ZAytwzjbiWByslgg7gsRV1o+7ZCarsxZO4NlLZSrGoXB
7kQrGkijyVGfN1JNpwj3x3Dtb2WBQuPtjUaX8Xk4uI7QpzIEKlqKzwoMr9pTaqAt
nJ/8W9FTW+1Dj/7b8HY2u4IdUDG2qZnPFuufw4jUFL/gaAbAlSm6a5UF9hRS/enL
G2Np77kyZrNtYNKtAW3d68320FC+I4BY+DKLfcd1gzstxJb0ApL//akbV9z2jLZQ
v0sRyVULZJHEXr8j1UBKYk7SYZCXHXEcCp/3QW1WJomgdaunj+gPX4uPlujM3Sel
1qD9buy0t5qleV4c/CYG72V5zVRzi3MKoCOAphj3exgGVgnJm0UUoGbonq7+ZjmI
9+FVTaRyNsFhudVdUR9GdhNfZ6Ucsa8jJjKRqY6txHYGIgQ4w7LqPT1qy2xEF5oO
EC9UsbEpUlecfSgwJiSs+LY7QJsuWHTRVd7H1V0nJTaMaM2SwOGsppg607LHWXQi
DWz1X/bP0ZVJUD/VVsoxGQcEx2gWBW+wPyE36M5BGQaAFn6knKX+PMjcnhTCU8ai
APG7yGUF/JtPFQULYYmuhOm3pd6ZBlrYLhV26gGM2gvPSDHfy5TXJemFztewsy9Q
iphFBz5rCVwsFfcNKlxLxnKEBjtmtxuk2ITAbo8n08By+fMgVA3NYBWUQV9s9XWU
oHBuD7Amm3xcJW6PBWD/sM1thQbg70vmxjRr8pcFhuqYEE9K6VgC0uCkQM/sriRz
SBH63xLLdDwSaujcOPtfr6/ocwVzMu3yvW9+iW1zKBVIDgRQX45L8VqW+XOvFK4E
hpNzDcV00OSG7+0g49rJyyWWC0n9vT7CXV9rOGfQw5d3oyTcrFxbb/vxoUqDRw32
9nQ5mAxnQjFTxgFHG6PuTJtRsxUuZjHDSkC4qWmNJyaBAa9bE22Bjhdj1bCdkiaW
gzuA/+8Z3P1/0JyAXSPjKv3lVDb4pDOwNhQ+czwo0GA2Sc8v10mR8WJG7yEhaMg7
+3vu38bsEK42lPE4NN3R3V5HT+cgO6YKPZWMKsPzJeo6hgrq3PRMyZiSOYHQLEWj
L4Le2lbvvgyH904Lsl82CpO/ue/LhYaw+Am6xOnZRbH5j/mdQKiqNogXL8xpsCXY
GaYfq3KLIp6qX5Z6H1S9HdW1d94phTnoHOMT3Mw4kLcmbR4L8qQ0oao6LoJODOW3
Rj99tLvlEbZtLdK5fg+6RwExdITnl8ENOUGWkDjAafQXPYSq0C9njXu364gbsQUI
N3lu42/0rqign6bn+efnwDd3rGgaxsEMHY4aODzwLPYli8r+bGt/bZyf+eama5LD
wHHrHHgLoBUjOHuMo4gsHNDYQLd4RbdIHqinGr9uhI5IHwMhdkisvKymyMg0EbFN
PSI/LIreC/t4yC5aHfWntv3vC7cFkprjfxeyTu6hd9MOaCSON2jCshUZ8ixrvLCJ
tDUeozV7zW3liJqZm4HapUpLzuoUZeeXBmceTqovzvX/cmLqTVu2h3Pbg9hdTARk
bHq7FyYH8mNFOGN+gaL1PpqupVhWfo5K+F1Vqp2OSsc6vkWSjMbE3Bg2jIT810lZ
1eNcpNksstKQYmAzawD727E6SqkP4+0/KSplBAY5GAn7jf7TRVCkubfFl8xkFl4+
ONNthnhv9DCf3yMyDkjKhv7C6D0UZctwmxiEkG7xVviFbQLhtyAY5BEezCbt/2hP
9I33gPVwHwk6lX+/n0mVhOj6Q96ejQ6xT+e4Ilb7fwkaLdUji5bZIEsWe59GCyVL
6h2AaSEcQaFdtyPwHf9iCvwLVJfx6PzfwPXu9dzyf97lTlShCsQpxC3X657iMChF
rzDXjmKPkVQvQvI2x0A8jH+DUIk7nahOKYxB4uFBCKj5C7xKUmFpQInioiOD0OB3
w9auPclOVdZt+yRvVPQIqcZMN9emYK+PFJWC3CSD7XkgqNFJxCiaj5gr+96bfyI5
knFaPfT9d5T+yODUHGeCGPvZm5gtr2SKa7bCp8GIB1cyPIlwyc+laZ6aunTzPzqP
GactgQSyFKAJEsJ2hFaIDPqBWHXVkKJzzphBlKLSp2irty68GUp5QtL+UkaMVuzb
pQM+VeUUo/7oo7/i50Z0DM/Q6+A8eK0mheMkXRrS8Uw3aDgrlSbimpoKUv2kDUEz
xC90jtzapX5wPliHo7tvYuw8sb7/PUvLHXhrkTXj0UBxzUQG1uASVdyUYyMV4j8Q
dLjNsO/L+FmIcEyaUCDAocbeoxmnxEhseTt1aPDFWUtmgvqPITgShalRHk6/5QVG
D9gdGLAaUnT/lpG8GaURm94aiJb5F7EXP/in0Aj1KKnNfXxjijxT65a4P1d5rBIA
/WmtLMMN1wj/tegMYNr6ycP/aYfj27YgPHUEZEBnRoQeGocgWrncgRVBRpdYaYQY
PPPMDzm6GQXwNJ0YlDDMxSARWC1WKfs9RT46kG8hlbneIyAbPoKt7aIeKAnAh+jn
heCn7AdT0ZDLjqoqW2UOv/WZXmg+6otRLEHWbAAzNfwuiRxJshqACMMu8t4L/m1K
Hm3I2sXZA1kEGguuOj3OygaaFgO3OO6PkIP63rHzfc1zf10gtcncpq60X54Kf6FD
XEpCx6XUek9JPdXezYVzcuEmMxha8SZW7zknivFmwzZgqouMDEnKw4/LCKU5yuN/
eIpWERqlvYmnPP8MQOv8Z9h3frwXe4NX0FniNDsapOFqhiE7cr05hUoUTPnFJCfA
Rl4R0ovY6F5c51dhnViiiNwMSZPxJrELmDa11tKC5P96l+v+zTfHKktz9WVS9G2B
YKAR44xq+Hw2mjeoUAo6gemvfefOwBPcV8/p/8dGClPvNm2HAb8eL7cscyLWrOW9
xIKvQtz22EL/RgIwHALMAHI/Bz+IJR/mAUtXxZlv4zXloKE+2lqwox//yuIQhN9N
3z9Dp0pGubc1tbxwR16mwFvuTmnEuRfNAOiL4WTQcc2amX304bnMOFX1z+OBOc6T
TVrmU0HtSP0IpNudfXr1IBtCFOkCXPpVwxvAFi9Z/rQj/dHOsl9YkP4qfsiKsxjU
uAsJWT6LYaDwrruoz5izoBLw7mAFle9EVkgtfO7i09wI0rN5flz7G6d87Os920LU
pClWaNr22cy6GOtWjOLeaHYg6uFxwPCGate8Lgn0moxA58sVaxUIxwOTB0NNR4cP
EhKRfbIG/ivtaTfiYTKW3N0WGfVR+7K7aTDdP7JwGLOFC1mlPq3woX4iZycbyvZ6
EI2FKor3RyLPuATQOb+EFV6/6JpDoAzpPbKX5c4LF52YWuajdzbEDUrKuIAg6xQ2
p/25G05thjIt8TdCJ/pYSossteMhvKRrcJgWAut0rC5OpggOXh3OEbKkC1czin9u
2rInNMIdWk9o8a6yYPEKfqPdgfyVgumhMX5KhLW8n55JvvkwKapTbm4F/z8rvook
Q0otTIFTmpUvDcMa8XvMfmfa+eK67F+mpmT8pLFe81syl7GSIx78AE7a3raZ9+4z
+YM0sh0prG/eKpuaTilzUwFhqBu53spsitbupqB7dez7DA6ud32exWR5xrQ5MN7Z
ibAWia1uVdOIKxXw/h/XxaIfCXu+RD/u1uCOWoOT5wJ0kChbNXCG/hIht+VafVNQ
kIzl6jjqkAFoH0Nu140XWy0tNHTBPKo8ByzF4Df/flP3VcWgBq43wvevSOm0XVTV
E0df8jj+kjD3cnzjMpmqioPRHjdPbOf5GvkbxZvwtMlUAuY+ZcVB6/dxiDTFYzlx
kiZ2ymfwhfjOunAXZlVzjNHcZuMQRxNrWfo9YA8kG2a06G8T2EEXvpfBHYGFd6m7
ZmHBGd5aA/PD5iA3UoM0MvdnOrvqwlfxgslIjgp6ubMiXMsOPX5Xt9Eu1+V7wkNg
VQOSYh/7FbFAqSO+KoIEqx8Y+31UOosYHpqydWCsJ6MVaWUqlL4kFxhHC2jRqm7r
3SyVuhK1Cfsz0UXHU3ZEGuETChZfzWevPuMkW798/rXY077QfxUmZRJ3XMWZzijN
YPdA4jW6ue0FYyaRB+plDLF7yihhZ2pArKFlSy1/cIjCzBTWhgYZrd/A7Y5VvGU/
5qq7qyHEmcbc+St2k1cU0R6Quzft8KmreDvpFKMWuNekkid5ehiYCizonrbytezQ
0ZBAY+O1lO3FUn3cYmNf6vQiCBYDDudRx0KHmUYac0s1AZe+qQc/LKCr7HkAxl3A
+9FVp4aSHdjIWoK0JaCuJ/khZCu25+dKqj9dA7/q7+4RSVvEx/iqVga0FJ6lgFES
iLZOkqY5v36iMQyaTntsMaWxw1Hax4YmmyoYXA3XM52uG+Gd0Zd1TTV2P+bNXgqg
oZgBmeEsLIAmC8xFhvtveVOtGaczDdUsyfW9XvVcmSpr/ls0v78EA18ubtlDt1fu
AwhNREVhqIi7UZ1wRhWnShZWVzvBuRtdXPBxj9KxmQF8YHy0ifvCmHz0xpotV7Kv
JMzoWxAvsIVEgNQBZMd6UusiKt8fvzPuNzIyLkMacYTIyAKyV49uXl13mQgaSY57
g8AxU2fbSqM89/aqkFBmCTmmq/Z8BZXsUX4Dld7Vasxv/KXYJvsp/+ooqmvRIt7n
nyCxKRIoi03cXBMFSpc5BjrifpdV9zBaCMOmNsjEcFgDD5JowYN0+OxbtSwC4qJx
myj50EOGNKxwh4IObeFLO5c/9w8QHNZvl2OYqG5kd8NEKhypZlSfEwcCVw2UpSNm
JKWZB2yFmNnpywPDcQ1LdQdaomZRo6wpZPIsyZe0k6T9Evd3a6tLbht9KPyhK+/6
dTOQX1NjOfUokELrz1A9qmh27zh/U/ZFRaD+ayhPR8jYXOAWRaAYrO+hq6UiStvw
Nr7157NVeft3ASNb+z/pOxpz09Hfx86tItFALvz2Is1EfDLwcuSTHFK3EuLZYbUD
G7YBiknRnKRcMs6fa8hV43KDEuRnCyK9RJ9y6O459GNDi++z0fFNiABDQomnFJnr
ppOAq+gHD39Jj4qNm1DglcDExKDYzV4Ov6Nic2DtHC4Ag/gDrBG3Ekh2bjsK0QMW
WTd7IpJ+6/MWXoIjrr5V2QRSVPZhoIXNTejFiw1dThtw0BIkdpoRa9OC88me4au8
hZITH9BEWgaie6y+6ww7HPgiCEoybK/4zB2Zc2VrUGSVmJxn2x8CL/rO5X+ZenTj
Bt6+tuYquCX2M/5k0v7NC5HMIrQBnrE2msqJ4yR+zWOyctjCiKKj+ee26A37tXSt
bw5bMbXfRwOWYQQ2hbsiNWO+bcnOjgEo2FT8gPcj5KvW1xckwqHpeW3V3yc8XnUS
9XAZwgDr7aEKknuHE2YWKvjXbwmIDQJSwD2FNAHizOQQehhaENgrMMek/udg8G82
TqLZaAqR1byo1QfdtuXIV9YAU1ZWweZREsw+4pS7o6hW7PhVV5swlfjRVYhcds10
AEikJiUyjx5ysa8sUFjLZEd/VIWEiBgsLaL9w5uhN/pJ0YMA6ZtRAI5LhM3X/xqP
szYOoKYklNPA+LMpgsXbiFRmBo21WZLjW5cCeFSTHiGPnhta7FLqHxA5nofD9yoL
yacLEacwNgrDegwxeqPjilWL7jcm99cM91wmhVQyQsoHqpsOdgTdLA+8KG5nXsv1
bzb3lvHdI3FUiEAA/Z+KdQqTGesJMgQogqt+HfDEjAczekozLBev1FLzem5zh5zx
C3tiX5r5n9uORFY0MM7tnGLkBixDxAv+YsRTDsmrugToiBmglWo8ShCQ/3MDz3lW
UeJZmUDUEozKt5FIEiDgKa5Y00Mw2haYRV6oI4pK8Dz9hqQx9v0YSDwwq5JARscW
IHWAA/lcgaAuzYL8yNlUuN5nxY78V4blEb42EgNbGu2F3CGWKPdKtXvBZODyK4Bd
XBvMYiYZDCQ2TZJGT9Y1gfDmW+ZxDCKzRl/a49uGMgc3Nq/r7qs/7SJlOls0PcA7
w7/5lmm3UVpf66/3uGSFk4zED5iLPT6k71FCw8bHIJEoxvT/CzMuif4wqZA35XcN
6Ht1kDOKlKWz3K+rUD6nfY4VN+amo3VNNmecB8+ufL7wvOb71NwtoJvWnZUFrjd+
/z/URQ52bSPXwd7nf3D0vnt1s2aTF/2KHZls+E816yduCxI3/EsrxffERoGNSjg5
FPN+YJLayKNB78cVJ17+eDgVHBQWws9T9pNUqmM9Eykb83jqw/wAsqaO1hmr2dMc
M4o7YamJhvNv74twtcPb+xoKmhXi7Lkdu190C8CDojEtVVSl3HrDAJMJenvEf08F
tct8HSWAll+NJgKBnyOeNzQbNoPGjiwoVJBcyD0PU0ML/BATeZgDAH51u+FUhO3H
L1ph+6ekXtF0GzaKpRzNTPxmREbcUzjtW0jo19mIcXFZMmscjl6zBqa0/FTUZaDn
G0TLUB5jUBtMCSJVzPtAm0S1Lw/MUY2Rb5X/T0Q9PiTrp/QuWSgYpUDxvr/W6yGJ
gE6F3e5fS+gCR0CJxHmaRP4yRW3AKWf8YGtEkNvBLJMN2FFqwtXEuyyx5opX2nP6
nvxWa5WlgHEDSuJWc+yn2RPhH48COo+6bjkORCwCnpslHNYAflBORLSfFrB1Dkhq
BPTM5M85c5p8b70MAk42uPe0K2jsGWUzQso+YefZotcoUgFALG4jArPPQ7ivBhY6
WDzzdsqEqq3OMv3eXqLdRF9uzWsTwWKSoEZPll69lzMJ63I8tSyH7v/IB1+DoJ4x
7a8qgvXdTqZL8RBzb2MRjIok44Q1yd5oj87AD6Wiox96Le7Dud9YnZzBY0fWuSvG
A7dhYm/YfN8N38/xSNCEEeuAeiaTauX9Nc3SqNcy5f/M6LUfObuFswkvjybgIQjD
a5Fs/m+ZsvRk4sJIt4B8xnVEes4A32HEip8EOXhar5+Ca6mArDtG+oEerB2kZHgj
ZUzborPnYEF0iiBt+ndRO5NvWIYl0KLNh8nBfuu9u7JowI08qIS/CycGjXTFnUNJ
nXad/GFRCCPN1QPImRwQjV6IeRi+AT3fWvPvNwgdzPPMN7MNlXu8PN1Crdsw/6n7
Khan/ae16YisFOt2XS7uNaT8c6xuxd8JzcZFKYUeEYL/Lx03+TP4or0P8cH9zgam
/uSurkVoA0LFnOK6E7Cas2U6gvxrZl6u0ohn9glq4cxKrYIPx7YutklhAsCe1GWn
Ga1gkNOLGZBgfVfwXUOPZyjA6zkxBHEOOb2YQs0SP9sLyp6bkhxCHoR9YiQzJwNV
2RYXvWfCQwBp4fQtJDP+o1kHluji030yLVemL3buKG8Sv/mLjucc9BOczBs0oZeq
RzDvcaDfJelGl6EZm4D8dpbyHyQ2xrstungonk4zk6+94HFZtCOv+7OjWefNHAp/
CnF659Dn7idDBACexmGFXPrhZulyybM1fThLOEbBqismgYOH/EmkLHoNbFLXZMwS
KslNyL+BY4yuVLCyH4rO3bPYJUkNR2Pt5Z+5pLkWrkZq+48dQ1F95xhxr31xRIIj
lEvDKS6QD56lPIIxC2B9pi8tdHVeXC+K3g63om6OGXXCEaYd1da88/h8X0V60du+
dLhpaGfXoQKWB45LNP+bPCMTDierIJLjuMIiphbfTKEsvzyRK6kDTFSnKC0qfoEt
gb4Lwsz1NavzaA6m/6R9PdnwPlZK2cS8j2LzVSPmuvc0EosynNDXmZjub9Tsghvn
nCV5zHrkZlRy9K108NstIAA75/Wqa+e3MegvyQR4siDYGG6nHPWKgdrEb8Qrzqrv
+w99aB5kmWM9WFSdQUYbkF5nWys+toOoRd6vF4Gx/gKmy5Eh764bday2mjJQBH06
LUIveoYEqwoeyMT4Jbe7y/LHCDiGkrxEJYhILquVDEhSMrGbqT852dAO1WYgWyMY
Znt9QFSywxAJUH4EL93cQRmOevLzTQtVNCLfZdYLj/+2aviBY8ARqnWEmIjAbrlG
JUMyMelvDlZq9N3kH8JW24+y4iQqgi29FjcgK6lsd9xcMqfiUugWWyYdpyje4laB
3JwryXutdJglkSSs0hcsB0E+em+Ogs3KMRgvAUmaC51rvhKpX0xibhR1kmZBBGxj
kVCe7fPdYgoDVFt38VxO1OTRxfMXsokOCZzkXMozPrmkB+SNR/6FfxbTrJHzckz4
xK/qbR+oc3Jhwx61Um+AufKDhwzHPipojxBstO1Eb58+xMriBtxoe79ILvZFUsxV
gAC+5IYAdrHsBN4yiwOFN+boMGcOi6K7J7I8aaNtX1h19s9mbD0j0jdjOPS1IPeY
92ZmYAEORLcsUaCr4YjlE+4A8Uww0GaTyxFiToigUWMpepgNs+nklWsmao59K8y7
e1Nab/hIE7H4P4AkmBeDlkPzyxN7bjdaOnriI+6eOphtbMFlU4SCfdveeKDKmkis
NdH2AJLAEiJ1eTQVB7ETWqjhYPqxle+3g/0ICpkaeYSZ0bB2oh9UJmUMEK6ngUng
IkOSvnZdjGNehNdb0LW46JtC43iitUO4nXQsNoBpnIunhBfmVRw28T2uvwFfuUn1
KDCamhpsT0sWRiuMjxqnhlCT3EyDEHeV4X5uMsCb2uFOsrHYpNOkKW9OnYdQIikx
Erqn9vCTCrV+PlG3XKlNC+jDLAaa3DKeiJHk1RPCZX/FX33KXlp8DdWgxHRsU9SR
ZRLghFy+i5tqivivZlNIKGuWoM+Ls5n4nGA3U/1mN8ls2DucQ6NhyDbSGdXSmbVq
WGXUhK2clRaPQ8v61Evf6obrHAEAkBNFOZfjlywwVpdf0qgw/HMMTexJv03YSezU
M1LlCtJLYZQ+nTDAVXZODj1LqIew45JR30yJl0VT+TxkXY2mFbIGdYOcQ8LXVsAK
figwIQZYF9+3R4soijRDasUI+aabvdplwpBhpuT6bBZTEjEWIpd3/KoLF0UN706Z
+ol7yLQNVvkRF6fYH2mnoNs6zZ5T4GSegO0DokKWwnCX4qzsapgWHYDGufyzZu3s
AoV7jZqcKZjAv+SxoI/+YtQxABNzDhNl57PboKvrw0TJLEbOdRFkOxjJCR/Gg8/d
Zeeem6qL+f0h/bec5FGGYkg4vEDm4/KaGNRv9orS34NFlvmED8UB+tVg0Z1HDPA6
G0fNEcu5KVIIVaNgEVxL4yTfwVwZpDdmvC/R+0HRhp4SCH8YYzDe981souRHQ3bh
ldjtMcz0CZK+roKhk1yE0Nnpvb2C6FxgElitF9K3QWklXBHWsUO8deIHlUxfc9Vh
6cpORNczhC50qzzYc15i0mY14FGZymf529Es3TrOJWBgP9Sg8WvH0A9LHBFZtE7P
OBWZ6Ry9aK/L3KVjcYotGQw2Hd8uPZdQpfIFqN7qcfVQEE8ijTU3wn0nXAFFTgQq
3uexys3Qq+8MXZLx9uqZODyXKJ541MVXUDe5f5/26kzcxWx9OIFcmn+Cw/fiYdH2
oshIgso+VnbXDWtQI2rEpBLbZ4davFHlXm35ocWg0nVQkuO0DKSU1LMl5Ui/Svc5
NRMjf2Jwm7d+awjIHjWI+frlNhUFU1BzBME9tKcaTK7hDBJ60kdEU5DvJOBW/hyf
tuseSh++dnF9L72J49Fsut4xLXvPXCKe4aG/FiUedtH+1KRrGBJyOB0h0YhK+mcR
WA2qYhr/rtqdVtCrLP8xuaobQapNoymzuyWsHkuCTHNMu511ZX0a/+yuXRd4xmAc
UjXJjzNSTk9t+w1iaKjabPUEY8vlUrFmRngSG19XXoEciaJDtJbpghimxeTfXbz7
xudcE3iPIZvdI0Jol7V9gCtQfgDTlRrb3Xg/aVUahy7OOXLnLE9Fuy7XZM/hMxfa
hL3ETRU4dR02XQkKISWAu38QoX0VeMhZDCMtKShpvyl39MpcM1bQWKmcb8lDjJL7
w/rGU1oTvPonzref9T0c6WY6wI4tJpSFfCOmmXVTKdR8x9rD7TZuS+/3TW8nqY+4
ixYJJHlFBnlGpiA6LeOa+phCmcsQyjjsFC9krB0C4OFtAtOUAJZ+v4mFxMwrCEfQ
f0h+BSIcHoG4tkChfE7ZuJHHzMOrRE0qS4nGK31AtrLlh1bGJkX07X0RxtpGnSA3
Dve9D6K+p6s+tOBo84QRRzK6sXmLtUYNL36na7PiBHmMq0gPIN1bafg3f+m9AdtC
6+N9ddsD2pFZjr0oBl0jJK+XaYSZ/hmIBVzA6/3o2dpUcbuPeaWhAAwC34qteK+W
YNNTdpg6a8aguuj2Ke9pcmo/HJI+RIgoLEQe4ZLjUOerOJMGjqc3ZhEmIuq2hhDd
Y+6QqpmN398EygZpjMpzb6yCCAF0tODYMyRYlA64a7ZfkHocffiBioaSQqMsQg1m
vpF90B7Rr61PKCdjZLAttB6gFQNDmK/92kLnvGif/WugAvou8bXO1YZW7eXg6agw
+CVCz5wBq9XDVcpY8VLAoQsWLo7m+SDK/cpgHcqAxmksAbQ32ljPl1P75/EGN6Oy
q/z9e0f3DxYDQyxMTdQrv/1IHlE9ymp1RFEFA0XzYEiT5j/czvXvgSeONYxbU1qL
l1Ah5RlMxsCuw0KRUp+ukl7V1JAIhR9NpgMrlFP77dWv4KbFUc3BHek9lXxym/EC
u5XkO/2jU0Kxb/cn0dmB4uSoKn3/zgZeszGbHx1jDuSObeyjCc46E66xsGriAaVe
YafhfFC7cPDGpYK/aAD0uFldagwE+nGOa/JLAf2Hf67g1Tpn1FEpDT5MLM/2GnMU
B1hCq8mTmnXOH48EQA5ujRayglCWJhBCi2TUSjh3hxET/sPMwpNR6Ftv28cPOfaH
SdHfZ3uTyS0sbd9yOIDfN54DaB7Vqs9oQzH67ncLfNyU4ebQBggrelb8FHoXEU3W
hj7VUrZCrwaZw+VCe/qVnDvJy4L7l3WWjXhcL4nI1s9LwRn1XBdvZXvjf0vQVMZQ
72s851Ixcv2rAJyzxlxPhjg0LbOVwcTfUsu3QiK2APg3flXaEtzDgYiay7YPyJAv
KS0r39EraNCjQtv3d6EmfOVUagEEjRVxfoAz1HndklwmrvwEaUYlxxwIzuiypBx7
K8UfLDefmJUu5j/OS61wPQx4uZHUCJF6UOncsKwdGNdA+ZULq1cDIZs2iVgOL26y
mOc+sl6k2yJi/PrT/56EPggR2rU2QflVswCQnTRh+eU//reSoPmNqKrWpypvqvTr
mgogbw4vJRQ/OsK962P0I5q0/7BrxjdVffocLrNW20EojdxTjbpptVbeVYOGxgAi
HgY3AnaqT/qSb9MykrqT6xdlMnj/OZNekJBN2bHFvPURKj+Pe6mgjBSfvOdQEqKc
HPS8ltKbTm9UxnucI1Bu16S8lZe8cViYBTs1W5Y8M7r1fD3TXHnqpZuuxH8yU5uW
4SXtJPDtdCpOx+bTliyGMAKhFlwxx63ZdqEx3xnds15xUGuXKwSIOrLq13Q0ljWL
DpRyR261BQVzCNUJEWhE4TFDnIR2DQb27qSKDO37s2DXWE5VBIZ8XoKIAoxVHlOv
jG4UP2n1LlB8wJ8M92zbTtHF2S1F3QtjfKKmkj9KISeHCo0EYehlpLL2Jv76TJnF
1VvIS0wtL7bXDYsIIFpL4WEKFV0ZX63YORMBcwCpNECH7FFSE4sluyUTwbH+H8Tj
4/6o4eptF58Vq8iWlp14z+7PqQtQpbasC9/2za+wMNZxjVG+e3v2xgIywLOiMQ8n
ISLtt7LDTXcstjumP3gRac3R6Ic89+QtMXcC7CvWmFEyFZA51UQLpWW+6RLzK7X6
FtZUsCkRc8FTpSM9LPREUfWvfeBlTLWtUj78FHix5tjmxurw+Azq3xtpBZFNO7hV
qGw/5kKdrtNRzMPeQTGzvFhomQ6Sol9e9WPjI1fuSnreEivZXHgL0i9xHgRK8uUm
OIyogbPcpTwKv77mkDwqYeW3hB3rM5/GhM0X6bPUE2MJq/fVIrub72NIp+9SMBpC
/iIWbIohMu7GHnNVv/GgrXF5WpgrKp10YhnNmph5hWewVsUY4IekxPdRN2XMOfi7
UM3X9Lsf+e6l/zojcM3eIT54P9Rw/kFFKDO08AFF3HbnKmUYioRhK99yvgbh3n7t
IODwFjdpSVKiFzgK7KnH/tyXaWn0NypzE8hVDeddY6ZIfclS1wH8fjJFFv7Z/F4J
KIuT2I1W6R4aZSk+GXz3b5X5y8CJXh9cz84sZ2Jr1O16Eskc9kD4YXuozGrztxoM
QN8AnfjManP40uyHL2pfT/ioNDJftnkTe7MQA4HhZ4IKAE+tqYXHVPo1kAPzgjCg
gmqwvOBGPxkB5HkkMQsI/ToTfPPwB0tW8X3RTyayfOzv1fMw6D9mzKZF/vyNrcAZ
li0TxdXK7EZzGCpO+nlIU7nWIe4eYveLmJQz1rZsa6i3AOMIgabWfwNDzjIvR6B5
l9uEb5VeRoHykFzpqpcrRHcz3FQxguO7cmQUgwrNHWt5tYhDWePqj8CvqeZeVZjH
5ObcbwMHGhTQ17Np4c7ydS/3pq/itxyDrTm5uKgA8yG3YsRDi1HmvqpXziXf2jBy
8nkgra6xzUiMn7Ao5vfb+2Lwdpi6c+0+fUAmaEqpPy/ZZxnpEevgmp+3mfn7Bjik
yPtQXXoNQOINoKMz6fg11pWHs4+6p/+Bxhrj3sAATV9JNO4HmLfpnfi7L4OlEE7y
yojB/LHYQqg2Fimjisy4igSLmRSU3QHs89TyoPZz7xMIIsqRaJmvQsjevZT7Z/U7
J+5gIJaamsrDIqXZNDOrZ3KbYCadItI4MknTQJJIAW8Qjh/YuyEZNrS9RG0ch62X
n4wikQOynf87CvptUkBB8kscv/kroymC4cOl4W2UvprnWUhU60jGmeA8a0ygkxOR
gMDynRrb9E/39frRKwDQRG3lQjsuELzOVY7z9wLyuhft25q5g5syQnW79irIQLhX
lbIwIV6klqq6Ybd8BDMSCRQ/KnUxUYacEVGzOUy9CL/FEksfCnIIh5mUBJeU0yQN
ZUWhz55PCJopCsxKqMhfOodMWdLGD661+sXbFANhzoxokyAlRzAOjUR4+w2EfqkE
F/JAIL+u6GZmheMMJaXHGWzzE5hrdISyJD1N0h3NjdOtYcdrRfYkyPwm45P7ywYF
SZwbprKej/uYBRW2TU7bgLxpegaHdXcWaBIqotg0nT2+W3rIAjCqP5lvSNFPUe9h
oQ2QHBhAIFstrBIorX1GGJ6Wy1zSKEFj5Y1x2L0TXoIV8clWD7qp+njahaJ65c9i
MZVKSefpSO+ERd5OZ92MCK9PffD51ZEt5Rc3nV+bSNPreW/eb74QlI5OIoa6hIso
uJkdA8UtH3cvbbRZbRNBYRVCfeDbcR43RTm+avTWle8wNLqQ17nr4jRRvgE2jZMw
tNQwt6pocgm55H5oteAkdbKitcjr5kH0coFacC5DxbfoAJUscwHNWFyaqr09y6pL
2SqqWGekkv7wHFBpbOLfoYegFobf92EuhovpNH8KMRw4YrcGzh0O+prhKfiC6vka
kMl+UGMY8SGumQ5GMJzTeExwn0uuvfHbxK4x5V58A8yI47BJ0C4C/cO5Wl3X5bbH
n3dOyNmrAbRUa1GNO/TjfK8iUpPfSY2y9czdwTzkxw8FvB0bU3RqFR/6cNYK/KhW
RJQqFX9xDQ0d7FpMGCoHFUoeRsr/iu4CwH6ZaOtnNzSPsRyUDb7+Pu/rbY4YZ0tL
umS+XMB/t5/DsNtzyZVqMVHfVVTecqOQl3mZDwNkt95q112dHYs/xpstBmm+UlEt
LsSowOS7s+4T90v3bM4JY0wciUwWdfiDj7RN/XsBDL5MYA9PRC+cT/7YAhQXZa0q
KzKQevSvKLSmDBF73Jjx5qz2kk5jViv2yuDqDOo2/PnpTNxArD31HYpiDx09ZMnx
jYEB4kjm8FD7p/AFgvofBUFzOntZ9Mdfv7YCFsrF2fW45Z0SQdsa9GXgymSeM9sn
3KPsLxVOeg7LZsV/ehvAXT5bwPYmlkqDXtFAnRd/HTujb7Ig7ceDRuF9zUOtBvFV
tvsIHucW3aHxB+kE0byMqDlehLyoOGUczfP+YyU72ePeKkRvOPdcZJC1D3ksRNpT
X5/76m7I45E7N7Kg5ptIi0THVFTbVYG31JALzmd6du/vE/xtS3yTG/6/LiM1BJui
DXa9nWjXPn5lqJHMQg2MoGX0GpLCQqWyGv5jHPKnE3IaPqtneavSQA3cTYVMR9xZ
s4LB5ifvlbV9gd8ZMGHVctuUmlfJO6up/oi7grcQ69Lft4w5ZiHQxW1po2EbS7ll
5mTVsPeMpscP+CZNOdUKANZ5BihBK3WVyk+8mnmie77YxMjy/XhBtkYQOyfxLANn
9GYJH1xzasGifL7dGi7Obua7+us2axNNTV3d9NPl5xLRQvPMRNZnqDY54a3eFZ/C
SEmS7kAPrqFMzoVppKly1W9VQSNqHW5RELd4QQaVscxP0YWUpx/16psy/vYZqWnL
qnwD5RrabqQgJpWXCofzzancHQh7LI87bd4F1jDH0Q0BiLAg9Zjshd2f9hthMVk8
4EoPBu8cGZ00uDQlU0x4D0EnnIwgTOqmwVqy36jVN+QFWVZARN8houEmo75FI3EF
z6NkeMztW6LJCFXNqt53g+u1GHwxCudKFd9Sd5u16PtEsrHjp7uIBDU7UM4bCCz6
tyUbd3tX45wQ4QusDBklIWU3E3HWA0vR2z3WguQE4DMn/tc+dAuYGBI7N+RXBVgk
tLiEjvLhkzq1ir9rWZzUcDaPMq5Nu2olA7n1b2WOHEnE17mFKwYsDvgvbs2+iLTZ
aL2bc72hAiwXFFOeEoHotMfR73Ii1YCYwD7R4Paxz7r4FdJ6OTl7jC5t+rxRdMTq
f2Y/A5cvFK86eCQ6sTUwQfwQHmDeYjtHc+HL4m3t8RvYDJxoflR05z24Axfxno92
q2JcFxP4aQg0ZA9tWh1gYRJDMvux/PJkARQNJEDH18l1+vOShd4axWI2jHDsV+c+
lv/WZE8x0DAWffdPvE0otueUi9wks0fx3zuC9x+0OfoRKv9YEs3SH3CcBkwJBKLe
8qW+4XsGuAqPf+RES1BXAu2YJ/iRgbXVwYzWwQ/h/YuLB3Fss+UpRh2E13GTSpLB
GdhxnU472BD99hUPxJUwMC8TjTb4bWiqk5d3Tl4KS9hv1zZ5raQKR4ZnKfiJNHEC
vLzohcu5kuBR1RukWYclzN+4pEpbGfXbHECL0/dBvALxWbyO/hnnT6f5a2r++i6p
XrnPRDxHNslyKPUBJqTkFEGzwpkRWGDiqZU76FiVzqdGCedI40YBX75SrIzT2Vp/
o8ZIjSuXAN5ASovT5bEBLssAag96WIJKpZIzw266OOo7gqL8PME3vpVNu/dYp7xL
mep5dRfAKKndYC1LepufIlL3hzudyqku0e65JzPVRIM+jccuU+MtdqfzRKrk6WWW
AXvnn+Gto+mJKVl0Z3GX3zLIOA8fZAbcZr8LEHykznlgJwHOGY1gtvDpYUnob84O
P1j8qM6miKzPfuBwNCqbLBPLQ6D/HudzTg05WAFbs6s91cVx1LA2L0lc0JY+T9yB
ncMPsN1mtwJE/mOwzXCUWJ9b/apkOJ3+AM8+AKfYsEO42YiDVcUXesorxP7jADER
7oW5QJevh3V2ycuAmVyWi2wAmeIFz21bO5YPO/HtNLzOSf3oD/zILH+EDyHuv6GF
aLsr1KVAYX3Qd2wgO+X7ooKo00qkqTSLZ81W0FMHefKNqCzaQtPL0S4dRQnxfz+W
YxvlnYR3Q2vULZsIkCgrKBmttQ9uDIRqv5K8fypa7kavCByXOHqcQj+BFMtbjCMy
iWU5gbzl7H/JTfiv91tI1wERl5aUC85XLNx49MdmZJV1kv3yWON4rIxBY/LpZZvi
J64caD8WiiYXzyQ09lAzQlqmQb2VDtNJ6hL2jEYmg5Cml8+tQR69dcRMZ9ahI7FH
Xs739+oOPTvBkUQDbmCn/e+sveUfq74m4XQ3TCjw3Cw++qM84bm9ZBTBAHcl9tk2
9jenPNKZhFiC/JlK7ZvfBkm4B/FglIYKPDW15ArV+oyp66A+YPghT0mG1qh2HGlq
2VAVboeZHEToLPQQlubyIVL8IucYKwZkhcfBXNRRVce2NZ6PSoCRaHZcHMauUr/o
mmbFngeltPk0jurW/NTLXGtt/diyk5RM+haLG6canQuj97+vLqBx7GlsFU665E8Q
W6E9zb4yyd6RcAmfQB0XGE0I0gzo7I49SvgkKsFetn3TFjvVtLYW1g8YxKJdt2D1
vDWO31jQi8v3JeHuS/hOS7o7cYNfDX2SgEH1f3k59TQ0AcqAZyA3wP4i9/R7HpQ0
24GCd1mRoF3ag5OmunkFgf6zh/25eIp8kMMA7SAXXrdKfFrlOGLeuou1xpD9wWTN
wJl8kBwjpAKHAROMvaZMzXwE2SWPsix1ZDo6cziBosiv8dvropDyAZjfRE+apc3G
OsScBxOlBpK8CGQ6ZW2fmWhQdK0KoFqkA+vCz8a330MEXCep3tNAM8RoH2ktAbgg
0Q63hSo8JSlo5h/jgk0Cr3A2aKkg0L0UxLHolOvNm2Asa7Vty7Pr0r6K+HSxbTa2
rONfxqDfyiCfmyb8CFx0WyUNpWl11dThXdno81GgHk1ekdfPDHl2ap9tvUU8OXa/
itjX/RpdPL5+uYdSdVyLFqDQ3Ql0uQEl7aKlItMtClCIGjkPsAzTTUoiQ8nYJ+cd
OAjcUnOcA5WqPh22b1V/MVNkmuVANcfboY94kbKw5y8wWUhuZlEd0DiTSNDDy+TZ
zZTGMjjLimsvuhLxnGZx9nEvzbS5i3XCpJeTIgNK7WW44PuL0uv6EEYAd6LErKw8
gyO2oHHkx0Zo3DwJ6IB9DmWrvvPgfqwTGm3wc8/qWWVtIEnRNcbNSgzDEVFUDV7J
/Ck1DSzpQg+2iUOGmn/NmUeYY17MdssL9tD2oMvcU/NV1VxLw/QdSDJhAvgJA443
4N2b4i4NN6dQ6ueWKvl97nhZR1Hb5hTSCL+St2kVfV1p0efrUrKyz2xOnVNqCf+o
ItlqjQaIJ6DepABJGx3hk5RC/MzD03E7YYZfmkE9qSf+f1N71vuL2n1Eil6g1JIo
odb5zqQiIjAK/d29TR6FKemYZyDq7Sjc0PNig8FyAXGKwzxIK74zCbjUvXHGDRzN
wW+o+bmX3vu3cfJh50dnOPSYNCA2FvK/9X5vwzxn+VAbXsvmlh60AmAv++WM+pbC
KYbZeYepcea+7ds5z8e8offJinuEBQGJU4CxZjGpPyIu4aRTmLEhLXUGj3wtnWFs
B/PkK7m5G47R0TwG7fX8cmfO9iEy/EFlpkDkM9LvSX2qtq5AqfTb8WPyaYKWECI3
tJp/zVsI1CuYzcMJh1p197hnLA0wltQIzjl9GkiddXKwDme23Zt/rA89eWD7KmNe
0zosquK94bBoV1F7k8OEIRwcjCdaT0WytOk9zQ2ihk09tIt0iklpEHwOo+A9c5m7
UuKu9HQ6Y3e1+rgG1AfwxHFssyFx8BxSesNfQHW5uy1HUz7e1sDXNf7WsvvVybjW
XnDl4n24TxDVEGMQoyLJ/Orid5Y+0VlMxsboCB4n3h4cjsLIKU7IwwWMxWL+j1S1
Nu+AFQ1bEd1h4UFtLrgKK4I2g8Ca5jK2HiOSURBjp+9GRNOdrDFTpkZEJa9EEaE2
dfqseTT/CI4581T+k05MuZ6ZiIX13zkjhuTVwTHR5siubTGDS3MhZ0aWXPXBEQ20
7JLPH/sxKaL6c6QDtpIH/Nb2SrHdNMtxE24q+kqdfY54fkcGdGxZxPtOO3askiHo
DYaEIrBeAOZ0flztix+OPsEbj3Cw2kWOmAOgxkoaZSzy9wfG2Wsj2d9OG1KdW5y5
1ulu+Ue40f2WkgGGokXN1MympDYPauNP3qVmRmhTzPMlqea2C1ec2zdMk2ojS628
7uUNS1HI3OEwmW8uRlkeJ7Js8AyA1SjpaC3ZxN/wl5SvBDqig2baQr/b07hLVnOk
YTQ2cK/KMGuM3p/1gFmrbgStzv1U+Wc9lLNGA/4iU6VrtuvNmnhtnL3gpBtcXkEB
StrDZ1BVdzA4JnVmqTYU26T1601K0WwadL97wqivDSUXjugls5rkqHiDrHa5vPBU
e0qjDb/MLIZjHlAra92qVEpMpP6XPbEHSzalOJAmJPqCw1D0rftQjufbJsSF+MUz
AFhnhLhCqCPg/j/96jGocuOwRAUqsmgpn1IUimxicbJWaQj9ngzWicV0m2c2WP7D
yf1kv6ItmUifOnGJOH3+JMhQ47O1CRIVgvVO3oTqzHXqTPQvbYgDhsTx9i2o5xrD
7HM6fF3U1XWP9dmBisSw6QiCcMO0x03M8arkGkzfXhaGlOgI1aw+Bdp61BdWkK2s
uvt+ZoRX7267v3A9OASAizENnWcVZ9JL0ZZ540kiuYRN/EXU1shDQt17HEMPiehR
a9zO6JB5b6wkqH0C/iEvQ9A3Dju7ugV6LkXJdNjePvDAPOUeZvA+v6slP7SzaJ0O
WaMn5ogxgKnKyQP4FpB/FU+h67FJWl7xhJSOQGCBe91NeewFBpAI/hQzmeqRJZW7
6DydoABM7Q+0cTaDZt/M90s2BqerHx1OKCubaBYXVHgrXana1hQw60B9vFpS0Q/1
Vorw8Fq/402if6h+CQWWzKj8qh54p5weVsvnp03ToLbDloIcO1rNkNMQGcf9iJMh
EiS6xaE1iUKPvW07ixLEMVE3IfzsaDjIwD/L8mYf71c87NwG0BM5EIg/Wi+23234
T/BqQifikJE06PhuWUSu+/K2lDUOogyCPXyzvPSlkQ6aOjn/2cvkCYnXZDsFLvLZ
3U3fQX8M6/OeSy4iTq17V5fsZTOipubBauSrnA6wme7oslQbk4tSjOBrgtw83igF
vhCCGG2ebdLmuGjKAPJ+4Tg1AEZIluT6jit65gzrqRlp5HzN6rzsQfHE0xEB+DAy
BImJhkFcPZomJOeFIeswdPgnu9FN4UGJ9ZmbXIoNqkWqP8BnOpop4BpIrBsBWrOa
IO9qPqejXham5x7iz2UcKL5Arc4GURn1tj+3IdxXbAdC6YhcKp+sHUlZzxa2dU7O
2p74Qegr6bcb0otoGFy7JIx7lVp0kTY7LTb6MK2jjS4atYqlfISSEA8BqN2Ujkwp
yfmgbPVflzQxJGJ6tFoMQF471h8HBT+7YqC9B5WL6VApd/LWOaiBXaJCrr5GSC+p
86hYlN/dDsUfapvS0PO1Y0hnz4obyjQnZk3K8qa4R2aXzoYmjSP3sHt38xDbOQ2l
9VrAQIiT4u5AEnIwuiMiwRktsGUtscrKkASSpPMYB+GGkvWQ9VKQ3/2iN/QC296M
IibmAhuxcJqM4KWhnengMOVwMW0UcB4TqaoD+1GCeQjk8G9LsSejweHLXYAp9y9h
blRhU+CGeif2KY1KFGXaiCZFvB537DoHTSdRN79OhUkf6QEaohFM2EV5OVgjXT5Q
yifXmhVzhHQbKcTi2+/Jb5nxROu9cbmjV7HgI63SRq7k9/TCcnInUKo3VWgvxqfi
tEtHCTYJs+nF3y1qzFjii3tFQVXGGZtonNXtvfLoWCYV8UGaFkHHz2XNbryki0AD
aBR4ANCrE5EraW8YYfVuMUZ0sVNS0nWNRnmimuHiA0Iikd6dWFSJ8uyacEGIlgXC
hO4nAzQNEZ0wd2JJ0tMoNO9jkiBSb/i9UsZGXPmtNpBoAklI+3/fW/+APsv5XCJO
JirfQ8JctoLmtfaqEmbgTyNs1mdpO7CZTfmBxXDya7HN/zMg2sDic4g7uCEpHx/D
ocHl1M8ZkXHPB2PuDTI0vS56i3QHsOpj033ud8jV/VrZvM2/ciN1U/RKHeLUBeRS
Uduc78vtf4f2Y+CFzvwtAPjfGra2MR9EJ/OGvBWG7+QzU9iAk0GUYqOwEUqrE6Df
NFRncmz2/fS1n75zO2aJr0rH3RQ/8rZzr4xK00pDaHHfhwQ3+giuY7xTrL7ZktiD
VAXXLJhcp/CHvGYczO+39ns/9ea8p4Ce0Wu5xyqS0rRtYHCBL/k6GnM4yqliU2y9
B6OWbivrJBxZ77aFdQE4O4gC9FOX/ExX+EaVjd4+Vg0+DKTsTkl1vGLQj0qOJups
IH4BxO0qOZpApKmoiMJ7/N2QQBQK1Tt/DqLnMd2S917NA2gmap/j7qdXwEtwycu9
FGqhCSlbq+XVsYm2qEMcZrcW4Kw0Lmk7AXsysIQ941HNd38cdDYDbm5cF/ZEA+/u
HLt2OVR6uvWTAD6HlQaaIjm046jZABNLokgY0dy7wb5wzH/zjHB4GzIXCmptkD8o
fQrbE3e+n4HQRZogcka9kObFgX4xRYRAAHg1ryI2fBJWIXwlYocFeChzvDMcT7XI
MjrT5hG8RgFxurb1I4aFzB9PQqT+/CtMNsI3Onlhq3wNEzWapy7Pt3AGVTghR8wh
uwfhlu0+gh9sGz7Exrs2toiG+yOdjEuD3KUjcNIsRiCNhLgAFq4BqZMOpM6cA7Q9
dUTNTbD67Tsin0MGXcsh4A==
`pragma protect end_protected

`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AZQ99ZROEuvG0M7tIxrW+DnR1FrxR4IDJRgwOAXsuL6/kdviA4iHW8m28uoknude
EiXGFFKYfsqd9xMvbfipGy22/Cp/RaQL8N6vwvDUERf3dHzNU+TaCXKozvlmRh6W
DCjIhb8xAJPfufT7bOubAsthAp4SsFlQeyxfh5mGqMw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 125859    )
mdD8uKifJvedj0dks8cBFnq8CIw+IGTj//yJwhMQW+iT/CT5ndLweXenJJiy0dSi
Pl8IDKjtQpndMtddhk8a6/aID+91yGwpmAUMSde8daf8B6DSLfu9neCzn9o57Fxa
`pragma protect end_protected
