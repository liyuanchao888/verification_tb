
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
    `protected
ggf5+(L<RQC7R(KfgF3Q&]c-SHN5IXFbKM_+YSe#F;Yd49ef0[KL0(KgHC&2K,^,
T3>Ug:MY<.U9U6I-4.WYY]0\OV(O)F@7C6c0P_:fa;=82V0CL9GW+HY2\gYW/L.6
XdO&Q;2@Ta/V.H7Z\\)O7<LQ^f&:6Wg4-=N&OC7e46856,R_[eC(ACA.FF^1)EOC
LV5TVcH_+8EgQAR36@TgB,LQ&[YaAbH(Z;;S8dCJZ45)B>\g:&0[,O+g?M?Od)S4
Q=X,FF\EXU;[P/>-TRNa)P8LN3#&7V7&;e+(^^WMH>@J\gc[7bbR\L8N4L+^T/(?
@HQSH]bX][[HLO;89I-,:gKG.c9808Rg/;M;T=)K\0cHMK8<+U:F93<F(LDQ/C6g
X)<cT4T8VB^CSS0<g<039,#&08?/-a10(&+AfY05SQ?]MF90>W;X7I?_J-5\Y8.T
EVf#OP?UK2)c_YbE-+4_X[G#J[R=SEbdUg-W_QdTPMM(64@P+^HX6>F4Z3DI.TNA
TASII9-;FeX?S47ag6;0YMbQA)T6c/P7dc:WN:/(:N+Vg]=8gM5b<<;Y?T=BG?>I
^/>RacKEO+60H=A8S#fITYN@0(O=].VUQ7Xb\Y.Dd];6N@H4L2?[EXSG9eSPcC)Y
U1K53@4;C@V7KWE4f)a@4K(/\<d&XB_I)1GST:ca@4O;bYVC/M[T5^SGM$
`endprotected

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
  `protected
>@d8&)IP,S>gK;?c-4RXCfY3W2gV,MD:DL^;_Tc0UX;>4f/3eH;9)(gL?C35g30f
Z6C1HKPGWK2-70S[TADAN7/Y7c&206AR1Y0GJHCFfBBFI#,/C7[.5<d@2TNfc_(c
X-CA>Z<(Q]_C#X5@:AD1;3Ce96TZc2:cWM;f)AJ<OD89ccEeXX>[NUVH2N>:4^N^
CX;MT5BL7NXU/)N_Nd&&9TB1&.Q)c4V>fIE=c54]]ggHZ9^8_dI3FE+T2VXcb.61
Ya>LadOcY/B<<L;g6@E;YXB16$
`endprotected


endclass

`protected
@4S7C(8e+D88UQ.4]Y^8P77SIZZ>J(9=GKSG(Y_OPW1TF<MG;T8@0):80H+.ZW:=
:MdSgM6,FY:ccLf5NSN9GN?BOM4H&Oe:d,eL,<Z(&??W)<ce\_QHJJS:(c.):;-0
bNZa#(#(CVESeA/^4F77BCa6^&Z())Re+aX>JN>C<H9<(bYB,?6,U,LN(S6TdP;/
C-V6d,.Xf+2C4[:P?L=^LM?,&;T,DY9.UC[^V+YRQT3?H9@\_VeWDGR8f@R\6KJF
VM4,)]H&FRIK,6I2E1Y6([Y-<+1[YY9>5+9W7Y^<U)X<<OH)28#LX_PE>@EIg/)T
K=f.e(bT/5QKA?-^g[MQHXY-7$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
a6HHPZ0gad&+eK>aI2-/(+YAZY]&0d2<X2R?X7AP_L08COdI2Naf2(1Q&c;VQ)=F
=&YJ/=)bR(K4=;N]S/.6bJ,fLDG)1.P2C/6EB-(5M>@;Z=Vc4BFM351-/+>#2SNB
V32U=+8Z7]#_X9JbF?HQLBAS,J[9Ug7aYG+_Ea-RO)\KH&10^dUdNg,XT:UNdJdZ
PS\OLHcJa4V?=\bFX\:&=:TTAHS?R+Tf5@3G6#1D]>6)fb(G4b54&?]f]7Sc)3&#
cHfb5dX+:;MM\B.GRX)3.eTAI5Eb2/e+OTD<&&,cKK#SC)>.K>L5NWA<1c4bS<L;
W.K@?aNBJ)E+?LFO1SISDI^33^[U\\4R=WASN8NAEc_\1eKFQT+TLd_TeD#PCP:.
LeXT51W\]e9J#>6;.c3_[<\OVbUU__bQB6Q<HVa(X6L6WXAaGaB,De+/ccZ/,N(=
]c.U7F3c2_7^DGd3KB,^&/9(EA@-gYHaNQDWPV?a6WfOLHTaC2T)@2J9]^\7>NCY
HDHFVR/Z:N_0AVPL]1Y,aY;V.d#OS3+^>&3(,L/,SC?DYZC)A8<=dK2:KP5RT)(6
A;8M?3&E30H(5>[3J#[=UY6P86XXaXd>5O](R35HZRM\T^51RE=X_)fQ7+NVdJAV
\XecJ]5W(f@7)CE7;AL1;#R7-E&6ER.^=+f+B+R=O25839DP[GSDGf^;(MY_TCGI
d[]&0g:-V27OC6H@Ud](YN;Q5)AIF@WS]]])[dX?&NY+:0cAXff;W\F.<<Ze8BTd
^P1Y,<_+<T[f@<4S0f_)X3UQ\Kc_e3?@T8]8=?2bZf@Cb8Z51_7+.-_d28D-<<HY
0aN\9W0.P47;>c_eX[&L1O5I+eWD.HafWZ1J]IeV=I^761ZJ1:J16Sa4Q#3T0]ZA
KcDNd9XC9F@],;ee_A_eK5:VMGH4a0>=E],)QECIM383b>.=gG<(X_GMda<4K1OL
R)A1SCg-;a&6-(WY6Rc;4f7>Z@Z&T6EeLJ=3QH0c]7fE:=EKcB^?R-//6>99bXeO
?LFZN=B6.:=^=6bb4Sg.AERSWHLMT27Zf^#Z53A.4U<J+bAO>)J4EA\-6)G\a:(\
QQ6LD9H(5-23fI>_OZ@#9\((4?E9][bDc@7:XUb+(24U@?GF/H;d<R(BK<f9M&E8
F^TH)YDg9K7&^A_8[5Hd+0d&Z]CWNaTCODH?M.6fZOS4eZIH2&<WY>J?C=9IgW2B
_,deG&/g,(?R)(2RU3cBfD7]5P>U,4?TJ+<Y0MM^/ZDUQ).@S#QEgXJL4?OF?B5[
P&8>XZIFU(.4Z9SL4QfL&D&\SZU&A#cZMP?--3OJMgS=cgL9&-R4[5_;QZX/@6^(
HLagcJ2ULeB,Z=d,X<4&=XZ?N8E2;P4d:#e=7Md+:6+373EIMfT07?,?Aa649U-^
K,@b.ILJ0K.5KV[+X\.2^gN,O[#b.\]Y7b39[-W6Kc+?8?g/TcNNYc91fP/g-BB@
E<RgdOLP81S0<)&WK0]=I1CSS1Q>)@c]SQ;BA6K&eTJTGT^YN3G2NQ=EA8E79fOa
@-&F7e.P?YgSc)_;MGd>>=:#3UGQM5==QAf7@>W-cPa2\;SBKe8a;NG-H<UT6Ua?
[?4DW1(eI_RFf,CB?KDV4JLdI.FJ>]7Z?d.d8Q(2EGS+Pe]KcaL1.JAPcG\b,(Nc
Pd6GCf<LYd.>4MaQMF11ABcI18#/P.F_XbSU>V>T7,(\R&_a-;PFXTNE#3?O=+]B
Df+-?&.-J0GeI7W+?@\<CLTO3G\DWSOR-+]2_&]_HCQ)d,6XRJ>8FZ<:4I/WdIWB
]f:4VJP))/B:AF?IXfJ([_(K@VP@<R9DI#c)GZ.9WJJ\VVOeD38Vf&,X-VXG;RPV
c\5CaE5^c@TV0US4#^ac]>4f2T9S)N5G76^+&Q#]]S=E;FFK-Q2NHE23O>bL4/Wb
_DSJ,?Gc@=4TR7A<4bAF&.Gc:/=W&KML/EKI+5b&V)d([HCCRPMXGF;a5,V7X/_C
H?,^I)4D=3f6FX+bM-UNL+E[HP49FVaYP\5&@.>&B^dF-BP;D[\4K(O;;D/VY\g?
KT/H?^=((4=ERQD@fGBFGB-8/S5MTDLFWM;<bcX7;;OFTE?e7GA(1e-QfFG=Z^T1
WNKUaR[TOA<;W67Bb5Y7(Je>-P(b-gPH:\8YHBI2VL<-<[4eQV&4NB?FL)IJK8+/
67KHd:_,U])R[<3(C>(/[U4gaNA^8E[E,Ga7M-07e\NT05V+ZS\G4#5/HSOJTT&B
7cIbR(_PGY0RHc(7e.\)(:5#.SJ<=:#SDDJS\_JUU^AKPH?XTI<W7:\FWcE>GU+)
?JH-(]<S.VM7O]36E,NO](GSW#,WLTaDABZ[g[E;R->6,^^)KR5W3NXZ=LZYM;M?
g9S+ZbZf]LDPU^/g>4FFG[X^.H#g1IE#NcgL3<&18J3/S/FA3-GH3Rc/2#T?K+0V
4D&4J9]K>QXGB)0)YSG<YEU-KTZFd5=0fa.\]Q#Ne4/>AMSY>J9K8fSb:EbKf)MR
;W._/P?G4E?Q\3G[)&Q1gF>OG@9-C03[6@U<K1.;#Q;gF\4f(RcGR=:56c@F\<^2
9\83\M;X#PIJO/EdR<F9PKWK@8I@b4<[c_6L.^K]2[TOW:G=?BYHH_R_<^eWW>f5
/^b[O.#X[+YUO+?GIP5HP_W29c2dA[@XL^Jf[QLJSbRZd01b0V@3O:,.&<M3B.e?
>_=f:,7TE:^4CR:]A44C?+BZd6[DfX(>3baM]<FfW5cIY5A^7VLB=9Q\[2R?G//[
;9FLg?[Hb+OS=MgIg0-/eMJHFA>B#c-@PV4_(4D-7(4IAAAB#8HR[KWV_)(4-D?C
@f2(NN2>dVPS,Bc10fSIT90X&/MP8KT/AKaZeM.HFINWFYf.b[f05LJCVOe^RNe]
TC-F8;UORf\Ef(544MH4NY=YMXR@1LKNXf#fGQA/,#5:R7X?:g2&2[@;&#aD?95g
E(&65fe8+g<d4&\+,0._#.NX2[)_8BRYK1T4CB\Kf<c0S+-?6]?=-A[+2_7a=>[Z
EHN):QG(RbSZb61[].Of-F0P&gW<dK5NI57HQ_OFgTEG?K)TFb^\<dNd0&fMKLYI
Q-^1/G#.c\Y#T8CbAO6UE1N\IE\eEbeK](^W5g]IG_-H9_8-LJeUAgHEaE6WRSOF
:4T)Y9e;)+b]:3HBg+CHd55S;,]F]8K,2ab/SYH-aD<3\Y]IR&6_25B^(Z(=TFa2
UV3(+5@d&GTcf2WD,WT^e^W\[)b?I-JQDd)-J[K;DE/gE?36&6c30A6S;6L,/:fY
F=FLQcc^K#4S);Mf7=P_R<g:TT&9a,;X#Ac3;2GZd09AQcJJ,#L4]=-f_g5>;/RB
4?_/.[R/YKL.S>b62c^]X3.A5N?2Y2]<e.Wa7(AH])4DDOM]I@U>Z9,2X39C8\>)
F^<A=K&f].7F5NXf58&JV#\\7S&S#?/REG+.:Q&A]RfT^PR[))6M-1Td+C;g+4Q0
T^\b:U@W#8fW4[DUGM+A>V?-RM<9XRQ0_F4&&^V42JZ6K3[-;g2,/IaC0,#K&_^,
I3[;a-UDC^?FBFMY/P1SSJAUV@FIHC994Gb[gSc#S5,KC3)^88+M0V<C\XcDYQSJ
L:0:b(c.^)=14D67K#a5=>J..B3(;EP+8=@)Jd<8_bH(E2M2U(@([Mb=_^T,CM31
cTLVIH_70@TaH3S^;CP\4-/)@a>\C9KOSU<S.0J5eVO;JTV0)Fd:5O<M?RM4/49/
M>GK&.d/3BTSYTH;0M;8J_YU=BcHYE\EBPf?g64Ia9gN9YXOK3&#2\YSaLT#4[[K
bM=U<P^Jb=89T-/,520Q@<4&.5@5)RBPLeT(E_S[1Ud-UY]ZOF@P199FK,/^3JO]
+S;3,H&]H]+ag?_/S5cWd=PW&[X-#^\;B:H2NKEOI.CRQg0Dc<</eA1dBb7M6X#-
D]=@<YW-T>6[?[QJc(OBC6149/^BgZK&G6GcMI>@W#[4SK9D8CF#HTf):;K\H/L^
(LGQW(E04[T::FDOQNd;7D=S(+E#Za\^<,JeVBA7:T?J>=a1GCc8?T0K>YI1Ga7,
7NK^AJO67_-.P.+eAc-YaY>&e5Eg\?/Cc7L];>//IR1b;>^\G,457,P)]5BB5K;,
#G5JIG[aP-dP^^LA(DD_NLSY1@F6#E9C;X/7W_8Rd&]cEM@4C3MK9/Agd:5g3eY,
O7-TC^7f//g&D8CR-8.4d3^NdQNaYVRdS3O32JKJ(.L,L\0,\N-0VHEE:=5[N8+U
ef[].NacK\JHdf2[W>I5_M+DQN_W>E(_RGV,b&A(]g6a):JFA>:4_?aMFMcC)LB)
A.2T,e3S-Y70_OAR)fNdTA?-KSgCV(G#bEa4G[0e6IaKa/+[<GY.NB1a+3MB6T]@
[J.d5MS:d1PAA]IKVYV8eE/^(,&/-7fcfN?aP:eb2=MM.,.JBT>c6NMBd6g+JX.X
H2/TD8/Td5UdeV#8&/6-X^@Z+A/46YJ0ZO,ULWB\_ZKcK8E38LF]N:QT0]>L8;=_
D@2XZ^YSBLBbOH5A+88J#L8f<-3EDY146QVU+-(:,U7,EX5b@DK#+[BABQ]M]L9P
8(3F1R3g@BIK4J/[G,B<.=&DV](^fXZYVgO(P/=;\Ng-@)F2Y8DJM/S?#[1O&G)N
;bU,aP2#T2A^LEM^)V<A2KQfPZO#?WF4dg2CJ1:RI3_7/BR0Z1N[c,OSg(=J54==
DZ3&A0Q8RUQPD,(Q;Z1)6)1RJ+5@DG_J-D@1McNAOg].fDI1W[g5cEJ2-P?#.<&d
7B8-;-45^XfG@9HM31[2)Hb16T&&1Z6>H#5_G?1DZCVJVP_OR=e9+?B]Y^ZgPeIX
R/:/;J0bDKI(0+0FN(CND;U:5^)705B40E.=FM,KUFOOLPN_TV8YD-@#VP]HRT_Z
OGP)UVPSGR6.3@,2OFPG6O;e>O)a31^1gRO5;CL^,:ce<\3a,)DZ-Y@UWGB#Z2+)
W9E12#>N2_NB4SO)WT\@0)=Z1=4(W#@6J6P8]5##SQC2g)5K2gfEf@6<W]BO5HdV
5@N+OV=FU.@W7/ccK-VVIR1U<HM1+T.K6QA#_OUegIf3S09=0K;.J:PQX4<L)P7I
2:5]O@F:JYV16TgJAfT,EWgAB]<EQ2d<K)07cP;/Q)c.2#\e7:U)]C>&_G22#CbF
<JI/W6W^211GORJ#EQX-+,1)]R\XbRfdZI:RO&Q_B;JK/[;;NGG,10-=EG/Y:P<9
VYa#CUKIHV0=>Y54@0/4Ia_1P(V/eL,[O951KT&TX.Zc@^4H#9(IgO3:_2[OCE09
CGB<L@64L4+-#SXSa;57NC<11].#K5#[3>M1IE8<E=Kf=,M2,0V=FE8<d62e6#(^
X]e^VCgd=@,a;.gQ9Q]F42J)ZX:7Z=6.ZV08<0dRQGM_fLNYVWb.LO(a+cR+#+YD
8LR:C+4&5>dGA^H<5)2dJEH+-QbMEE@f8G49(;H<CXe>H@UOd;(=)NQQ+^aH1WOI
?Id8cg-MZa1(@.X()CFN(HVJWP1&g@>@S8Ye7SWTFb^Q@1dO(K^0YC8TN]N[L@SI
Q5F.<1,e-XDd^T\21W7B4T4ba=FXK45>T^aI03N?:1:>9/XKe,;EH(YD+WHF30PK
8G4D2X=WN(a5\I\7NBXSe1Yg(U8H\M-;G].aP.SWI>c;+A.#&39KIP2EP5;_:9RR
OOPIO=;\5#\1CacYYVEd&N6KOeZ+U,;G?JdH4J\4ag4fNdMdIP\_a+WXa4UCQNPe
Y>4e>:V5-SRK^V@VVHaX-:^eDO:(7?cYYY4B\S0N;&?T;G\+V5M.KVR2GM0Z6[F[
a4W2(>cFLW7FT53C,:C5gV&JI<:D>IdaJYX9OUU)2,GIPGU.Fe7fZMc_1JA4TE;J
4>^@dSEA_&.:&g2=C?IPfUK).2ZeIX9;)(=CPfaJF11;YWIgNEMK<-g]4@EL>7+Z
S9/T-CGE<a)B,0b8f;S:&&,BGPG=])>Sg\Ja(bTGd\C8(?5>AJSM+0Dg5^W&e)@V
1?0AM6)MEE+_/3Zb:+Ib=4@9:J8Q,c=d^/FfD\7N7&43(NbSRbTGO+,fF6-)G_+>
_Q+>C:KIB.T1=F/@4VP:c:N&\U0,+:@?K]R\\Qcfe,3[g6?^A+:Ia>U1FDGM1:[+
P-&I^YCbDGW\4M<>Hc)^5;_B/]d8W,>eQ.cR:6cC[^BN\CF:C#V9U6F@P:SDJ7I5
&O?&@a^W9e^?15#ac\3BC7W+AG24.&e1&fS&=GDR7<KEI]9YH@LH]Y@eY,L?YIYN
)E0YCF6Z,YJ6E_bJ)Wg/VDd^/4.[FOB)\>:,9MbNIeaMKI;T;QN<X;AaO8..?4VW
\01(-f#<4-K@ffgQLRc^cMF#93)PW+^Y/M_)g=X1f\A,2(SUJ?@(4HD#Z4./.-4>
:.7,#-fSA]G,<(@>@,[;PO[VOcaeIY[_D>M6^K-?_-^Q+;QM=S,+>1C@YJ+D1,VH
>),H=NaH_Ec]OTBY&9RCfK#EgFFL<XPAI&_PDGA#XaTVSDOTC#^H6+=fFFW>(C4O
8YV#f5>?J/KW7A&DE0O>R)a.H@:I5V_=a.6@HMBOFY2M;X@BXAA:0#&/aW;0O8Y)
fW@-Z.]>(R,=)KV-8NQ[W[V9,=#:=0cGV<U6L-9\cRJ;M:2)R#5aG=>;Q&HP#EZO
JP]@PSVTaM#VdaEPBYP8IJ6b</IPGbU?4MVCUS687W:dN^U>/cKKU&gZAK7-W[A,
[>OF7Gf<E3C(Z(;c[C2DD(-;\]0IXa:eEVMbE+5FJ+_V59fIRe8\I9ANO0G/3?Y_
4?Ea:8+Hc8e0DR@Q\L@<#Z8_a7Og9H9&W^LL&+,XSOM+/gKWc#\5^fZ7AdM@fgPC
#Da_7aQ0JZ59?=bVPNHXC=NcZIB&D5O_UVS\&c&3T24QRM3=&,+4OUbYOMYCaGg=
_f:5:6I6a>FV@@gN:DBD]6+4D>(.^D76dL1^087EMca7WDJ#GZL#]<H\BP+Ngd.O
Vc(b-6M>fV5#IZC3->Tc44TPf(2UcJ.@8cAHHV5@W)gYJXSQ#1<W9E8Sab?MQ7K=
f]M;ZV.G[UbMLIVgP^9f3I9X:T^\->a2RNPY@4-g@5=XX_+C3Mb.-gg(1^A-:G9a
g-9F5VQ>E)a1QU-GN&-eHAT>b>#Xf-[Wd[_8B\-e++4X:XI^599O8^179O7.>\/g
H<&[IFP]N,NM59^6a5)V2H&@VCFIgHMe;[JgJS09C(YYe5bA=?,K\YQ(+PXg4(d3
,@9PY58-fZTGAB&21[ZS@aPF+K<\dE>,,G#P#fB3e@W?@Eg/GYR.8VbU(C\bYDg^
_LRK(?]:\]R)ga8dUU(9gJSA(0SaGAUF^;CLG-A5.SI1S]8-U^VH]T=TOHBYZ1^D
@,93Y@WCcAZe@[YJ2JO9\@7;0FV-M;0S3_9&PXJXRF_f+^c3CY<X?7^A97fLZFGf
:0T9WG&-NI,3KeOWcQEZK\@gF)Qb=c.e[HZEgJ^XAf>[aQe5=&>&?M720a^4fG,)
0O<^L=8>]BA\>(C8;LId+-\\;^Z37d)\#\:4):NC)aTWZaRc<B:+#YX?88_/?1cV
H\NK?&C_#,+S?0K/@dY8PFCFD8fb0XXP--8[]b:1GbKK7R_,Ja]U9/,:dTAI#?M_
VO)@JZ:;cAN,\)OQIDZRDG6.[/9VfDETFVM-7KBgU&UF0T96AQR6a?@G)?HMMS1<
E0H.(43QgKF8[=O6ZcaS>efQT+A&LT70\POE#[3-)@NR8<UJBYC:OZI2KW\0G879
cI4aW_)>dVP8A_-JgAR_9M/WRV0+/>,-N7)c,Wf.PF4[P2O=M/a;,=NGf&>^8BMC
GJ2YZ(T.LRON+24@IC0FeV&BQ,DBd\=,(MYa;[138QcAV&4O_.YY/S08>INYKa8H
4Z7ScK1VZ+H]0H_B+P/:gILJ634&P]X[C(e[>VZDQg9L[]++;8E]JM.GOCIH)_Y@
BH21>_/+A+R][[PfR3]K[SU0G7dXHbFJY/8Q=+c<IdDOS14VTSXH&(=Pf&f=]V6>
e-KICeSR0&[#O>[9]=Eba_:T#CMa4YF\fAC.)EI-JPN>WVPAKZ0T+[HBb@GT.@8f
D#3=RV/TTEO<^]X93;7&+A8)C6C<Bc75>.B_ZR^R=/+3LZL7:f=a,VK)gU)9F[5T
;4;XJZ>#?87EQ<TUV/3:bO_OIgdJ7g5C?2((=a^>c4UH05#,83<QX+[Ve>-Ebc.D
N5J@HUL6ACT(;\L+Q]JY7+EP^I,II>,+)0)A5C.AgdM,-e9X9Q)[W_>_c4=NdU@E
LJQP8+R?&H&CK8P.gR)g7RNRAG2=P\K5.XACJfHN[c=8T,6](O]dgO2@?c^2,6]V
Ha2Hag:JJL=d86:+eaa4VP>=X8.cTCR:<Q4CB.RI9Yf7A5+@G],S_]-Y_.g[-Fgd
A9?(^V8Wb<M\;VTe8RU;c[?S1ZS^36DPY??DX9A>MR#7,4V1QN_1cdXOYT:g>[<J
7DAQ#b<L][CF8?HRf\^5aD0-FE>T>gY_>1\O<bgWZN\4eT6:G<PCfT]F=D>2g^\R
=QUKPg19cI5^]AX^56_M_EM,E#X)GVT-a_)_Z7(^f@Z@>7gOfd?fA9^b9VZXNUH>
.GfV>E5)K2)Ia[S_TeTCDA-G^VA<PR-c+--\0S:VGU)1?A^(S0J^&2?N__ZB\aXU
5<a2=9M0AOAV/d5YJ1P<NV3N]7NN1N@K/TZT<UG+dQe5Gb]/3)REQ0,EMb++1ObA
K>F4?bd3d:;6JA2;b#G#L@5aLb1;XW<Z:K_5ZET\UMS):a\0/MG;HbW1@K01V(KN
K=K/BIX;9Q<VA^34^)S?&NP\4J@5G<),TdA@-.4^=V];33?6_Z;<J/09B+c=+V,0
V]]aPT:#5.)g]]Z23HYeRZED,NAL2A]67DPZWOV=5,7G01Tf_SWI9bId/.b6=@2G
/R=C1S+)d>P^8,1+U^416Zd-8D&c8OH(WSc_&LM(Y.6.&]I1H4-#K[N@40fG>HI\
9V:KWB]AT0U?K>\A8AN3.,ZBP>5K_F7]5GG.+M)cGCBbffI2J6);9O3bAAB&^HM,
Lb57Q(DZ6>FEO.C.>Dg480UPAXf_86Ye)=NUSSL0e=EU3:cXZ\EWeBSfC4(+2V3g
F=_O-UXF3_QLTga6F&AIN:K.9HM>A2]H^CLQEAZZTWPR&.EaY[<Z^TA>YVKCT<Y2
M)E-#gL29RNKTdO6R)(E[AgP9P9M=Y#^V(^O.?^^fHF]C(-3,7V]La9Jd.?3b08S
de)?42\[]O<g0)9Rab2_BM),-Sa0/>_5eNc_/QaR^g+I5JW@3@bMZNPc8GFT1M)H
9#5e:B,Zf)Q+H8>YOR<<0R9YXdY&N-B[<^7f<SZg#(38@d3C8Y_W,EWSb.S<V<A+
U[g7VX=bNBJb\:4<M8F^=X+G;2[\X)#Y=cZ:K@?7D]JX)/SHg9e,X(BNM>O@\]:N
E9O4gT??,YH_SZe@-E2G4cRc=KX:6IP]9\K@R(TUG9:cZ846EK>f7^C3)QN/EYDN
J8(&RJ7&1[[\RBZ.T_];4;9A[@D@UCH8ga\BX4W3-N_QJI=_81TA)GJ7F@>Y>L<6
F1Q6D,H<W[7DWBGS<bJ2SI,?<NFcV<EW6&II8PO).3_96EXXURK9Xd#Pf1.Be+I9
b;).?Zg>+HSa?[eJ[0-SWR_4HXH>eN>&gJPc5[L2@XWH4G<Ef^C.:TKY]P?gdU^D
3eO@\2e870YVI_;5dWR+R)&2=I\LdTOTL.<\+2d;0/&b[&@:D:MFT5-]Y,J];.]2
I<D=_]Q+)CO=\f[c1I#SNYL(Z3)IMW71YM+Q2/;L^e)Y7b=]1/])CU[5C?K[TM3O
fR3KWF@TW,_7R3<N:4][MSM;L3]Z6Y\IA,DfH-d/Mec(-KbJ]4OdV&5EJX<UfF)/
A8b^L2LcGY#[<EE_SBOgP699H=&E\<U.Y>eH]EZg5VVKUCeNZ)ME-2a(Me8-@,=K
LRFE24:9bEV=2e^A+/A+FVHG0UC_T_be7=[cT,bJH#=\D4&8B#E9CE\/ZNT6Z7eK
IXCbPZa=<LQ>6gff5.c]87R=HfS:RW^@E;A.3-IUeDV/ZYW<1IF.GL&8PQ&G72K5
W(]SCU3&25fCO\\MN[(VK-3KZ/;g<K6ZL=]J<J@?H97N[16@YF/bG6+ZPUVc+95@
;.+Ug[LZ]1Q&AM==K^^\1EF.TMCCVd=3K2d;1+Q?L5CaVd0;dDVN8,:/HA<@N:XW
[U3fQIeZNOPO?fc7S>BNEP=d]A\-FQ4OX5&bcNH.0E.ZP/_7H)Y^bU&@Q8V(?)3<
.4]&6E?efXX3M[<M:[:ACH05O#;K][Vd]K)@ea(=R;C,J4S,1:\GT#Q&>f;+#&C;
.)=EX;Eg>S_1#c@0>,ZLDK2f[-cJLB:I8L\H/4\]aDNE^gZN-T9:^&Q83#>A\NUW
@NM-&?ZWBNEU0RZ7I4H^3KF+C]#?>C.3f-2ATELOCMX8FZ\H74bJ,3EfeXT2L4J,
)R@:2PQc1P?AM)FAS)KT]&bI>PPN[1\=L4]_DPT8#XU)35eZ[e83Y14)D90FV?2D
Kc;>Ue[eX8=gUS/-8H&?UU-(LaE@X2[;Z-d^GWC(OL,0Yc>__2bE>)<\X/NfgBW2
KN14_VGOW6<3\812I9P(VAZ-AQIFd/7@Z\6e]_FLP=[DN#c+PNWSC3+NZO4O:B+U
&Ne-\CHCX-</?Ydb#VEMTL+af.-U7TF-AS(_aR_Q6TW]d?Xe8HR/O?;Tb]I]VC^3
#X@AV+E]7+T&V_fX1>8c9faMO<4A/,,0PG[f.LO(&^c<7G6ee\7bO)/=-U3D@>#D
?0OZH_>=H5R8)E:2[?QgMg>A6T7A+\)BTOHI91.PZ;b0/cHD@D;BKA9<H[P8#X[<
F,MW+b\OG1BR^=YFe)D#5\SHg#:K;fTK0>)Y^80))2]VIVJXQ(@3L68R3WddcML-
VDQJ>KE&-?8_RFZEaaR\c)g6d?\43I.&)?#=I(VaSYa-]YHOOG:&a6#C;6/:>YPG
P96e#<F.A#ZS0R8aaP<138\B@>WKeL47ZB6EE@d[X+I.(2FM69/.BN.0\g7[?/V6
EKQ^6SbVegDFBY3KCR/?OL)GN@N>L8aW)1K31a@S(/1CRT18?RbP.2607cB^?3We
Jg\[B<V)--^2D6>dJ\0=eDeEfN[AKCYZg\86I53ROFb6=0;#a1O\AMTc,;OPXfNV
14VSL\:\(Z:^OJScW?BFgc/L_OE@<f[ZfZ,IJ95_;(&5:>eWF.fN\64BM87d5Uca
&5NbZ=JN-\A,A[,/W_0AB2:8@KS2a[D?7P4V[>/-FVcU(V,;,#J?F:f^_G5MA@+a
/ILXV>O)QV@W0Hd.B+K+:8SUIHVEG(B1??f+X&E?,LM]+LVV-MQ-BYVd+BRZPZM[
[775Vd-?I+>a?Ace7-+N5C1TVSL@3TS?)WbIG50ScS8+aHa:J@_5N==g:Hc03CX9
8>U5RQAF&6/4DN5?<BW@CeL-e-gJGV2?O[8@P9IH9FYH4(6g=LI4YHSH5.;J;LcT
K)-W+RcOLScGUHf)d>(O0IN&Sb/g^<DAF)U&5V3K40=g?VF#.1PJ2]+I>9>e.&A?
HM_V,H+Le.ZS.bZNNEGDea,-A]\+Z&=Ab(7Tf\gdS:G9O\MQ4?e#Udd7/[+?.N)I
LC^SUW48E?@.#BW7G>Q)4Xe?f[UR#(9XHGMG^FR7,G0-U7<HI4JQ?dL@ad+\ELAZ
_T83(6>>VW0CDNef0,N]-/;f@+DPL-\,:HVX(geGO<;QWWaZLRf&)^--@@d?/Jf2
<e6;(869I]ET#;U3(?Y+^7@3AW_GFQaH3+,+S]D4Ef^1d+FQ+,eC=c7,=04Ad@AF
#X:Q@4&X)<c>H^C6;A5X,Z4SV;d9@T)++146/0?_,CBQ)YYT&(FHfV^,<C5Wc,FA
J[N#G##[:NSKA2Bg^R7-eHB(UR[\?1L-766P6Db;7]b?Tg:698IcCVF,7)]E2A@U
CK<DNYOLN57RK^LFX^eHI3R?/_&X3X-&U.b#&;SAGV(AMTHS]Jd&_?eCD>:C4M5^
4+,).]D;H^0I(RG7Lc>]WY65ffI]/F21b\/P(_?J:2<2Z2H+.+4dRJDB;,0.]#,S
UR1R]0=cSg6)3Ec<\fDZ9Z]L8gF&D/R;0#P@OC0O8McCWfG@.#)Qcdf>K6C02_VY
(WdQI_X#_7^a_Q)g&^d=4H6/-MD#e)0-cT2?gV:]^EB#T?bIc(B[Z;KXb;bcY>)b
e4\\cZ7a(H]\+_R>8UOCO@bI(BeSMg^1d8<-4dZ8F_XX9(RUR&DKI:+eCY_LJJ-Q
d2/f68HQC8NI5fYFQ:++L+#&==/TYgPQ+B9FZ)E5U+SF/gSW,J2LX065g_MKOgA-
gTCCT&M1IF77>)UX?JO;CfGVG?0F_8AaS3)KSW1MGW\;:Q9X)50bWR\f.+C3&[79
ZGd;UPI,_#94?T<[LNNOIE8;ATXO2BA?<D3#:?@f3b0H4?OI9J>c;,/XY,2FO:]U
^d(;.>a-;4T72@R@aVQ.V<U5O>)X.6ZcAcA(Z&CL?HU<Q@d;RH5?._Z<W5eG5QgE
_@E;^K)D@/V)<:MXT81ag+U5I3#7g_LbPB2.C&6^bRfZ)L/]OgQTCa,M5J@SEB=B
/5ab8PU7,b_=b8,FE\G[,gNIU]4>+b=B@QGOF=dHMN1341eg5#.3_W\XdXM(34bI
I(c>7UGb8X<G#g.9>fZeM&R9?6O\T0>63dO^b1RXO4J8;VU/D\QT#ae\\c,@4fd)
9LESJ[:WQ[)HHbVCIOg.EF<6;HK+FK66.&A?AM4H@Va-2-0.NK]]@c[[egSK+-;4
g3TDRbO]PBJ?EGaFZ@f6WK2S8<E@P,:<C5>(:@=W42O?bDJHbPL#18F?E^MVEb8e
:PR+RV+5F+DX8c[I-3/C5&/Yc2E]I:)0AC\8N5[.d\G2DR73=3.2(:YK2CVffN?O
EM(T<=1J98(424_,cW>+9=O]G1.d</,dHCdI_96(D:QKe-_E2M)-.CYP\G8MaS_f
N-FIKW)a7-JeESR]NKI?I:R-@MK_B^dNSPa3GH>);FP+F5QZBf]7c:H<G[:\,>Re
1fF6_FWV2F<b_H9,c)>#VOY=a6//ZN-8)ATT;4Cd0XVf>YZ&+<dTP>W[4.6dJ136
+6R?=ST)N3^^#e)-f>TQC9L;fONb:)CE-.[EZW\76,-K7HScC)9I/9;(MJS]62=B
31d;5H><;=8#NgY2G[0B@0:F/-X.S[Mg05I)/gfCgC5>#e6DL1##;74?AIa+C(?T
]6,OC,:0CL,[;,EdYO8:MD(MTaeUR[b<,+\fBd4_BVJ53B<S\dB=.ZS4bA5+Sc+\
]Ad<+FW]V<cH0(AAO\@;S0_@04N^c8/1:3Pc.O^MR5&H6T[8W6K>c79b=:b?6#:K
HE:7>[aLY#b8/CZE#.(N(<CU=CCYY1V@Sd;,T[@K+T62beS);RO-MgIG.Q^ZM&a/
NfB)@?:He/4(&#L,8fOdC7(K8O,5B#c)YTV23Pa;)J?#7^3,R@>]1^Y6CY2SbgfD
[0Ug3aNG#-aHgUSTS&a8Q9GN/;3^:I;[R]SQ0JS]H@fdW]+?WQ+DOaIDc_6_AT99
M7Z&DL@J3>.(INM2IMPR_@5#2?SAf2F[[ePObK8C>Y)cH+AVACQ72]QJ2TA@^I7g
?8JB,O0:E7A8.D5V:SYa^1::<03<[b)_[8\GV^I+D7=)4<P4(7Z1PgSDB,OENJ?4
A\LR,+9P/TJcYY[e[ENb+>7Ta-KR8#JK5Ed9+0;XBJbZS>VCD+9Q>bLNDe/ZOT8)
a:CdDdQ=0g[?:@J3]7RA>WS9-M7X+@2@^Ng^S#R7UQ^V-c#&R_32EM8fE3Y5T2W,
?.DTeD([f#=80X2/(CC_@^5_bSMN_UdZ]FfV;EZdX3=J1YS0R6cMe7A<c85+TOZU
R:R40.d.#<+RF9/[&<(>@((]M>bJU\b;]L#E0ZLPAb//1eLW<Ea,/]P6,4Sa&+2N
RHNPZ]M/bG.cY(5<.E84e#2RHXJ5_?V356,=EZgYb8Ia&gM8)5RG-Bd:;;M<WMcW
3;5eJ;]VgID\Q:?JDGM1;&f5JC1&1XV^_W(J)>dVG;L2PfTIGe,)G=3M+O7Me8M>
4<62c+LdG:]X.+RL#);2[AUce5T@HJ)24AU3OND+)VB;KfQb&aU\U4)OT_LJ2M0c
UFMQ&FPZ2)DKg1-PBO<T=9H@^G]<0TXG)2RZ.WX(:DZDUT-BR@<A/645.:QC#9-_
]>G\D45QR9.#X&]D\)V_8N+XgCCg)T/=c0X7G?K\B>\;KZA/F[JQ9[<QO?B3FL8G
8.-HF3UF7R</TfaYGUgLc0(FFJ^>1Sa(\BOB0.P]R.R1/&@SWb.()<VeG;KJLc;:
>dcMKCTT9@eX@C^)HeGa?Qg3SQ27b/GAabWUae^LF1LEd,a,-:-EGX+^.fHW+<[e
)XK1?S/>6L]\M0eRII_9[BdFAOfG0fdQKP&eVWU^YbOfKOT:>DF8;TH3^S_V>Nga
EKT;@V2>AIP(?1206A@PD1BBg\4Ad_a#D&LZcM;E-6N56,/2^:RZG3QNHe1S[I+_
=8b9/@fe\<60<ATA3BF5C4O\L[O90/5dTU/6,>-#KD7B\E;.9&be<^4<@aG>:I;6
5M?2=<f74?00@_U]@5E3Y2<04JPY#,O;IVF1KV1+_D124T-8LYN#\/LQT#QH32L^
MgSO6Q@UMg4U^bH;2;#/Z#VbWPa=_@CE#A3QaDR:Pg]/XbX#F-N&+U/]T25X1ee;
X?BBF[:_U5)]0J0Y6[BQAF+0GTYL&CLL?JPBM)LeU3)KO/WCbDd/ba;_7XJ_OH)K
-TfLe1#b1TO#C^<;;(3Q9=4dG8/-PJ=4:Og2N.0>(RAg_PW<TJ@>]D/P=7SAQXB#
7L=MfO;3eaNa\?g?_d]BC_fW6BA1?7CdH)UMCT2ZG;-IXWe/HZH+ea)E,,(e+U:J
AgXT@6C4fA]H-19HdCf+^.]D@,((Q9@^1gN?dB-F\deARda_FO,g2,/4c)d19HI:
<8U+XHBG,_W46NTD/]3\7ZL7X[,;M=c3,b\(N\LGK<:JFa4-gYY?aM>YB3.FOOGO
6-&4/\VUI7Q?,(O(1eb#NAT;gZ6QHe;[__B1b=&4<K3/()ZA2cS1Qf\Y4H3cf63g
X(,&[5+K:TV\?E,Sb)KbeVdT89.]eAJ+\(B.K:7&?e4^(V=G+)R3(ES<Y9e=#(60
K:[=gKGRF@Ob>3a-.4d8>M82:5KJD#6MQRbSQd<R&;417#&G75;>#)0(WZ]\/P&>
]I=PLKQ>GcD=7gGU6X;)QFbVNS&U;:[35M>;#8a35QB5LO&G?MSU)U(P8@X/PA1Y
9/?<Y]G@UM0_2:(@gB[6NIN(#@#,>[g?CgTN<]ZYPQQP/L9P36aBNdMR(HE9PYc[
-@5cWL[Yb3a^(3GXcMdE4@c00ReY@\Q?F=:DVJNS,[M0IBDZ\^0PH^Z._CA\+DV/
XX;._F\6K@=H/S<2P3;/a10GQV</9H8g&DLMN3g^?6J12I:2fGR0;([a^8GO4\5F
03Y3Qe7&AU>N2>S5HeLZfM0(92d?-,7CPEVX2fA>Ff-89&@g@XQ>BS3.X:ZNA9,.
3XZOG&C?BF9M5#DdE7KDdY1JeMGc1.TbdD^06BV0[G4AKO(,+d):#QH[Y0bGVE96
7b<X[D(5eP1XYRe.(1)O4/6D#P/.CMS9N@,DV+S9#JE,#=1f#Y;_<Lb63DR[Xgc2
5gH9I^NN(1PV_@-&Q&P4Y>LK[PS]eeZ;TPR^(4527JAFEK2YL,YWQH81T_bIWcbO
FH153R?Y/0d0^+bTY4\JO=+.8[-Q:ZcO)YS&82N:9UR\/BUV@(/?/X.;)O?,Z<HL
_)V:LDK\J/83EEMRCZd0d7;4(_)-XYQgZO>3=JR3cT(e[VE;80/<UOO)<,(;QZ)Q
?C.8M+N[S+=N/+H(c)XHg65^>JMd#fEd@_YD[O9]2&96N4Y79\.&<SCK9L&a0[5.
aVc:^1\;_d6&D8#F9@V];FYKcJB<Jf4Y3)=1#a\2RJH.gK_B#D,]0@8M[^_c?KTL
,(?Be]6KOcc@g,FUD&<YWb;gL#?G>=>UGSP92.S,^ICI5#X&KRP2+45+d0-XdD\d
.]=EIfSCcW\(K4-8=X=O<^/:2:WLQ1EM\>aH>0I:4Y>H(VWFBGG.5BNO)K_;TS.7
7NMIY1g:.gXfV5>FY=)#62I@G9IQ<VHVVc&fGM0=J<JM8XA^C)ePOT^H[W8P.)UW
@:8PU4/53)[#V3HV^:fA-=Z5QNT=8cW)LP^[fURPe87-R]KRI;#WYPW_c.dI)ED2
1c24bOP/=LMLJbM?=/ND<</0<6TcOddY^JE;+VRA>;5d9ZX8U-HU7)J]/&.K-\O3
H(XcH\5WI/C#:X]H,=X@];+f[_9a=DLXU+>\4I1:?Zf4#[6R,^>,5C1IG(S8aCLK
Hg.7e+PcgASL?;9cML5YdfT^7Me-&U>T<1QYeQVDA^<.g@&V-f3LHILXKHQ5eE+F
]/+W0J\RQFOL>)=PLg;H(O)<F14/09E5=)NB83/.DPH,EX_JKA1K.gbW,@ORa;^@
95^/F?KU2?2/R[aUR@0@QDF19S=Of,]Z&;H)>B\1//U4^U0+ZMa]T,N93XC)+S/d
[,B+UgN[D78&e?K,N^dE)/7D55UUL2D#eF&92D9O2)N@W^fR<UQgY]5U^Uc7fHJ#
SZK)Ba#\Z-ZW<2S8+T8<+@?+0S2]8;SDd:QOB_cd3\U^PWN&E&FW?XH]&/0^AU6A
e+^XW\P0gPCLZPdICN_f4]-&<W@G.17C>4[b6#+FLZ[KNFfaXQH5J)H#)CAFA93B
UJ(YCdQ(<&PU;&a/HS9QR)&JSM:LC(T+)HQ;e5Ng:@X1HZE96eJ&XQZ-D2c]EYP^
g7&EQTJA:[MU@[):LfC>ZFIA/S:e+(//YMT-JMUa_R#X/efH_EL<P@--M^RI;e0/
S)E4XA0Z0P=Ea0H@\c\,BWL[K_HZbDf._O0efXZ+Y4#gAI#J??U^7eJCF&+P[9\W
HQEB34/=J\JFI6UA>b?\^E2b2,WZ)gL9S[C(7GSYT_8BC4?;0K+dBR-)]FC@fA19
&Fb(?K@&PQZR09N:.:6_PN=9(3&YE>9_F2D8ROD9Z[eQ+)1&=5Z.Kf2F9.@;&FJ4
4)e6[bA[2.[f_O6Se^RgGFQ)M#O6-G+fL6B0NEb1WHO@=c3G4T8TQ@@#AVRT#UKW
T#d-6XDMQ]MRaMG.FR7F&DLH3)9dQBZ<?L;V??Hd4GTB_dWY2e#5;]\?bOV&Gd;,
L@HSf/)&+K4@@XTLH(\P4&Pd74\Z<SVGCT5+/cD^[A2E@Je#^U..+CJ:e13;.\CK
LB5E_3#_PPC<RK<G#=FOW[&8Z3UPX@ZJPf7aT3(_->aO_3OL\14ff;[:BS?U;;8@
^;:DEa:E.N1Z6/:UX@E8Y0#(aEB72G?W<MbJ;04=GCe9)c_dRQ;I5(KRbE;=++^R
IcBI&5&MJJKFJ39-)TQR/AM,P)+3&KD9^<d-_5:3>>SVCKb&NNH>ae5Ea_A_]I<Y
S.0IT?\>gF&/?dSdEVM;3eCL=a@Q;/DCF^6[U]CWeK0@W.d7c08F1aJNS@UXV#H5
9Uc-XSbDBGa;8b4cB:e9QLC)5;>7Q8W/gV>E+g.(SH5K0a90XY4da.<7#VY9\9BG
Ta(3c:4M6)Q\,B1f^>/XL9OTb/A@?2bUF##ZHQ=>C.YGVM^D^BB6@2]eJ&@dNgb[
MM?eTdTJf2=7feHY5PFVN&GF>Fc&Uc,4?J<10P2]g7_cHOJ,TAV.N@?I\>MS@A;I
&6Gd=QJ)/X04Y(,e3Y]8f5b=\4XfU:L?2A]0TT[Ied^K4-B.:dAbSB.UX>d84&T&
O1@g09gO^YB:B)5)X)6GJJQ/CP(G:L52KYP#W_UY_[32W=-OT;J5]_4&dd2NYK/&
LdF;JZ@405S[#O+fZZF\75BJ25:-6I5V+=HAD#3:C0.1C.DV\H2@\FYC1ZR5VfIG
6P<a52.<.B7>7&=SW<;IOF)@75QbCG#O9T\4[3cVXbd9+:O+7=Re5eU9Y7+]R[)5
7@dbNM5d-554CJ(#Q(^<eH6#-:D&F5I21:,MGFQY]\[?T6f4/Nee>DR[dP1LOW0S
Ie&:@Ubb=gO_d[DdJFOL0T0-eW^RYU@F&SIB2fM?MT5a0S=0H9E&CHNeQ\]cT8W4
B/5G-DKR6]A7b3Wg378A4=.T#;RZ5eYT4eVHE.;5TfUWM:GZMEKgD5E(EUAT=HJ(
AF<+1X\M-bX#8I96aUQ0f55BAcA.EDCe[3Ne3(,#1\eZ@\gJ=,GZGV^YS?a7K)Y(
U];,F&_CQcL\?&3B5/FMYH7+7VQdVS_\gYaC;=XW94FbMW&S-.#<3Kc[P1R2a)2E
LZ:J&d/_4^dGO8PJa:@<:4,@O6__Hf-e2Q5J3,2#?<d?(=O):^?f/=ZL@8g4PU#&
,<:]I_@4NK,d8)\OS(OI6e0abT])N\@]W5^<7-.:V._M=g[:S#f;-W.dZBQQ9.:P
<91.T[C@Y2V1T9.@4a.F(U:[OIEXV?1e];(V\d@E>>JT]MePbH<TBC0I?<QW.@-@
F<N@]/CJ>2?E2&b3P;_N/<HJKC1/6?d49.d_?BGT4IMYM@U;HE7?Q3;5D;X-2:D8
BJVQ-U+V0AT6E9#)+VBZD<[;]./gRU]/3.&/aDF];YHU,?9Zcc,Y.5_J642,Z&/(
\K?_@3XG4JE-0Sef-<Y[aAWA;UEJXUJN)g-#BAPg+0?(TABXG]e<eMRa6c_PdNX+
\;-L14O0[R2_Lb\+QU574;GBF84Z=5:,<;XcY81][JI(DNXcV=48#YIEF2ZZ[HLQ
#DE4.[7D>6=K/fR()a81VXZB^#S4ZLQC:6.P&9^Z0f]C2/X.J\Pc7@gO?JI#P<d>
Z)=6.,1cA>=b3A=1/#3X?DF[^60B,(D?ORF-)F=?(@2)/X?>6Y;S+<<JMJU)K^8a
R2eI@bZZN^+g7K)g@SP5Q(fWM1</6G.#<f()1[[))K\HFcf#e&^,Sb1]+\P(XTe]
=;>.\-_/DgUYT2KV0SGI,@LdgR9eK[BN=bg:Z&2OYCL7L\gb+F3^_0#0ON3ESBeU
U68^JK(.a@7fIV.3H[eGQc/4.>X[1\<7G5T:cZ]BgY3fX;CFd#e(^;fTdg@\gdGe
A.fBL-d)98EBMP?KF,P9^7BG@TUR9<VTPD+4]gfC>)K./--fM\_BM;/=dYA<S4Q,
@5LC+:,4I[RbP0cBD0+&<BGD1^eaRac-\0A.+e6-/-1L@?=N+L7cAbM?WXaN7?Be
aLGH;gLFQP)+B5TQdC/EP;@J3f6@g=SdKS?JE_UW6OXaI]C\7>/Xb/8@PCM.126=
c-X>\[#L3:M\#I^?&,P)D^BBAD6MR[F/>[UHbY[=M)YbE\JYF=VW.cOYegU@@\Ng
4R;e^PQ7T]F9[P287IH>X.1Q70dGc]TG_.3Z:K8eeJLgF?ONUNe8,dP6F4K9.FGA
(B^ga1;Ldb2+19O[H_ZIE;=<9QXf]^VU?aH_CD#AKcf2H<g.SZ,)f440B.II9(2&
T/+F)RB+GLX<g]gKE^ADY;#3@^T&H..7>BMEKcSEf6fBMc/\3cSU:==P?OMe;F3\
f\[/EZ6[61..[,>KAQM6eGHb\EV\[#5/_31B(5DNHg0gcVg=]^fAET/@MT^LaI1c
<(5HGD>B8CBGNQQF6CJ^gROL72(feVSKFDSY+?=_C)>\MU-OS2ZGL/L>,MCJ@V9,
[eHOAg</IZ?5NANGRT:>D5?;X<d/c;/<DaT2.QI9@1#CTC7V],2PT[RHR9#\6K7M
DGCO-HI7@<TT2@aX.O>fH?VVX(V2G_b3B722H)4>MHTZ<Z9DQFSeJGPX_H:XQ.Qe
IG5=X+O5:eX_.#]e,@CZXg2d7OXZ?;B0M&K/JSO;bX+6_?GBPX[\F(_LIGML_OKC
RN/E(.)6>g>NV1.7H#/]VX=]P+7D9#M/CaW^b&HFJ@ES:DY)Q<>4T<e_G#7Q@Ec<
<f@MS4C--5&65CBCYP&]M[cL(O9LAMIT[\-f>4<)Q)1Q0J1N^W/Q+[Be6G-fPF_G
1A_;#5<FOUM.(2]\0OfG1_@TPLDW:QVW:4K-9ZcQ^M@:/ZQE&L/ZDZ]O?e#X+bWf
EZK]/HTNOS)50U)RK;AIA048YVT@PO9KG53>^D)0g/D.<@;F6CF@&-/#3;P\A7gZ
D\\2EY^(),ge_4Mb6REVNd_Q<?D][46164/36N?PPU>g,=f#FX(V]3Ad?eVZ.=QS
+d,SRF#0F-BECcKMRa\#.G@VZT47KaY[4HMM?@O?.P&SB+94CY?6D>.=@C7B[VaQ
Y.QUG>(HDDQP)QcUPG(X:\R[fHb_2ab/)<-V/aMDdN8<EF=<)F4]c<F?Qe&LW5^>
@Z8;J?()F8;\QPaWR5JQ>+IG#aU5I=b(B1^Ef3&c]?UScAPL<_e#/]E6Kc<\Dc<9
fcD\SFVfF_3;R.Q=;,@&Z?V5AdK_]YB_LRZS;@-b]/.0Q,RSLWXf0bDaZS/,B_^&
;Z=QLON#@IJ]g]FO.bBB]RSCMFf:GPdQ;7(:+]M10?^_Cbc_+c-W1Ad8P&],.5X]
8\8fcPC3[9NMD47A4R0])Z-VW4R[9Ue?2>Vc3FNS/3ND4VI;6Rg\5ZdQ7D;00g(>
+HI0/WD&gMP<(_3#?b1@XB:NXPe<_0:ca:.PIHcYWS.NGD:P:S0W,^Eea&H:aFWK
[,U&^5RcCP2\5PC(V,eG30)/dTBYZ_cN(AGCYZ[I0g6aM-E<e[,LQ?BR35_5>=Oa
)A.@VI^_9IU/YLXI;@A-O?DC<EMG+0N__GZgg45aGJIc4W.WI2_g4<5FH7+NJCPY
KGaOgXHFW3Y=K)geeO<]<PO?=Xg2:81e;0J&.eRT_XSB8F1)1EcA[^#5-a,1FEDX
T_#/33?_^01Dd,:LHZ3H_ee^8=N2O]eLTT&b@,ZH./9Qb^_Zd[.L:MB+S[0@6=LO
aU6GdAdc[Bd7FUU2EN/.9N</C0b6UC?DAfXag^5L^0[MSNF&Pb+0[?KZ6JA)Zd8F
;b+K=OCgIUQ,a2c3#<>5e_VTEKgRM427RdV/X4L;PB&]TS_c4BNQKD\=[O>?e_^K
cO?fMN-WOGI\JU&K-Q.9UEVP.[JCS@T&b:XEW2#^DgJfQX&@aGHbQ2Lc6_JXUA0@
D:5VM)N)W+Pca6NO2DE[57)TM/3>7DZZV9\SG6bN)Qd18/C>GOI,0R:PRLF70];/
TR[NNfb:W(VK=Y5d0I1+3dWeg3[[T^H5d9^ae1Q^[\F/eaRQ_T#)d&a8RLW5648V
15FQ:(b?:<X2bM\N\@4(9^&\BX/+4D_#RSe6Z6B@GE[G.Q[&Q<IO8T@7JWe5OcKA
cX]_QY^MAWAU9_#@Z/@R6Y?WF&^SXZ=\G>3gbFAE,\=/W,-0gZ3f[gKgW3+1,JU^
7ZQ>R<-D?&L#d2dW;DCIS\(B1AW9VG[[[QbM,=0LNL#=RUKOJI#DZP:Ob4OD.>]<
4)Q;fgd/X.]N[-<<>#^M;3AP_d)4E+NE8>bG&CGJCJb/f[FI.\:Y/QHSfdZA.6aI
C+G:<12F(.EEETXLWQ=\;2Z>NC=U\E]#DG8<BPYU18g#;-M2AQf=Ib9f[\V>C^#g
#I^P(KILY1L^D;=>T/#A<[GQ<(4Z+G<7HOcZ>>I-7QgIS)E18QZW_\?[>@EfNHg:
f8EWd44HaK6@^ea:T1P5LIcY&3=JNQfG(L88:0Q/C/e#Y_GeDJA)JgHTZK19e.BJ
@0ZI@>7P7^CV8KX(/b3HGeg/^9;Uc=RY\fdHK)@OO.<f@b/eBCND.cC]3b#@3^1W
5OS9O8eI:dPXbC]f^D@gG4YeHI+Q=[@5N0UG(?H2(:#DV^P._eB>KK3Uc@H=A5Z\
[;==IZ?60d1@^77ZO;VOTCaK.=<bZ]c/cbEgDU)BO,.<6b.A@U3C4Z_J<V[/&?c8
GLZ=Q@<LK3P&N\#Pe2GYB^b[^86F1N<P?F:D5-HU^14gGKK<+K&[VWP_bJMa,5Q0
Z2(W)HQ]=2bY[4IcaW<[([2F:J3FOLaP4W]3<:4Q;N;@\D=aWXG,NNHfCG0:PDOT
:2C>3/UP#9_78D0QdU6ECO7Q]9T&TDNS^+c,_,&[:]U1N;=OG)@6IU2MfID?V9,<
LY;G]<dWe[_77W-C6OU=U37]X-MU&Ya:fP3@6)S@&D:+SH4/d)5LY?@9>D#38Uf_
WUJe(&8FUcYa=[EJK6])/NJ:DY]ZKO/FdH5:YaN#^J7cWQ:&N5:].e]/]Eb2#X([
MfMG=/f-9:aC67e^eFOCQ=#5,4d=^TRAZLGHDQ9T,[/WB1PK#5QVY>E+9eU43;Q>
d+<[g).WFDN[[,8JSZ:fMETDF(ML.fZ;)V<,EYX51WJ3#?Yb2K7N4LP3bLDY(M.K
CgPb&-K-;/ILBa@Fe2KVC7482dQBMQ-A9(GT+N33F_)<?@?MF3TTIT,WY,VEbQUT
>g_98GgDQ])^KD1WDY61I6V0JDg[HAN^RWRHLGCS6RF?7NHOPH;.:2@-Q&_],MZB
;3S@SP[2L4FU.Se_5<(P^;A+N9_96-ONY;Da<5Of/BDe&,5O713c^/D?)bFS/=\+
KM8e<KVK8E3[3@\;WOJV&J(<bNV^34c#=F&a3=6Z<GD0STYWVNEa[>@S<<-[f7J#
bKbJ(;ES8;)N:-7/cAB5?DbZX<7X_.F>EK_TB0B^<AA<PR0HMD_2M/eK?\(D\Z^3
<f&S&eb:G2@0FHP)1-Ne7VB:W@Q=/<^[,]-6WZW\/2#XAE1@e?Mc(Bdc;<+8C11d
HZSB5NB&^,J^NdQG/\NSAETZ;HI\[X734/W&>BO9/B_fL\8d./=4[XJ(7=UN&OS_
Q&b,9VHP7(-@g2^V3SG0#fY65YLaZPT<8g8UL=<G)J\Sb2Z0:0W0cF6GVc_T^_)S
CfJVGTT70DeTWIS.)\3@/YX3-IS6@LWM\#@L;4]\(Tf_-<8_b]\D-^1b;QMH)Y]K
2KR88U#M06Na\E]KNS2P+UCXG3M4e3Y.]OL,QF?DL^;QBJ4-.UO?HegOT:2_(EH@
F4EgWBI<:1\DJKX)HLN#+G>G(W\8dW,CcK?S?AZc]QO<4B5/f<UN34eA(T,F?0Bg
S#PF.D;(?B)I.P7?.>:1?ZXU@WUbc8Kg[e^G4cW]D7;21e]a9>4c7-R;e\LSU-J@
=[L?a;GAL21d0FQCC)@Aa]/O1Y6ICcFH\-A4VF9c1_(A\/XHJL=/(WT61<4+FQS9
Y==?HY_]c/K+9.BI#X\R<.>0=/e/Cf_+7Yb(eGC53=/O[R(T<9@QK0Y0=?\:5<KI
)KW=Q_KIKfABS27a@fL05O5G867RTD2_f^R2H<df@^Vc,dN;[6P-Nb8BL9_&aJP9
\EL#-S@5Vg6G)R7]PF+Y=TT,08OXFWBdQ3_I#S^1:TcYZ1ZID6-^S;8Nc^/:g[A4
P5RcM+GRH)+GX(c.EL>Sbbb6RV8BVS&7TV6[WKb(I]2UP\9[7_[UBM3QSQA8fC(:
_I=ATOJZ+;XcCXU2D)eZ?:G+=0UT1;FFC8#@-^.e0eICNcLLV##K<JZ7Y+-L)O0P
_:Ng;_V)fD#QEMEd0T<c+&#a<I/7\gNG\Q1,V7D0dR&TN4Z8f@S4>LdP,#RKbcb5
5SB(I+gBGe<X77dbVc#b:^6U&0\fO&/AV59@TM3c=X<31d8[G?Eag/F8TGW\,J52
c&KJcKI12_dac;M3C:WO6)dG85^6O]aHfK<d/NC0=C:)^-fB&G?,<4>D#B6[_0)C
aNc(A/_:1LI#).C13W(CU4@^</;70K@N^3-e&)<>,(T(af/-7fD;ZRXLd;#9?Dc3
^E-P:.=U^9eM2O>[>/KPZf4Af\[9-aI<0adM33\62)+C]&F7a=)W:T)9OG3GbQPV
#Q\IMVIU/1dW?c:IP.2YeDJ,.9#:837NcaAUfdGQC?C1V,API(2Y3>IC8,<Z)73-
SdYL4Kf?RcdIRf)8)cGRGdVWOO69b(2)S:ZdIZeEY;WSdGA?.>@,;5(N^#(cdYaV
21G]XLM;CK\2]S.W5@YB2X87dc,QbKc9aGSH48B_eFIKZIfe4^F:5Z+I0.2-U/N<
M5T(T/7@.>N<8(CRcGAJ64#MAVRI?0JKe_0QCA]V3&gI-gYNOAB&AOP03DS]-,2)
20HJNN=G[g9>T)YHe1:#5&(LJC]LLN2bP#L1>M52K4<RXg2D0UU/IK1G=C84A#]^
7Q23#J4P)EF,PDJ/cY1KDJ27O>&O;bCG7S3W29M^JEHbK;MO32X>2]X5Z[f8+9TS
MY_L[R-O^#\_E=7U+7LV](\;KRUKBEY:1[3Tf257R=V2CBBJKILe_&A6b0?9ZbHR
I=ID[\bR6A5bA027B[.TS^MGQG>:@2EM[U-]A:3+7I;X@f\3cT/F0b9JA>H=4)96
BH751VK?\ARFf6:41<^F5Y/YQ/3+YCX?XNed9T9O;<Hg<00Pg)DbgJ0#>_K[(_f<
]0ZZ3EW^4a2c(eG-I-V50fCbZg0(?EIB\-#<M)L7ebS7VfM;\B?L[QJ6UVQ\W4MG
ZPG8-J(+K-P?Te5GD.Q83QV\J7/?LcS^_TKE0VKYa?5\170-:H)^ge_BB2=YL;:I
87M7_10W5<-E)b>BU_,gHL5UF>7Q_/CMH6T7\)MGdRW.4P1S3,R5cN6QTX_?\,ME
/OKSIC_IUHLeD2b^a6&^YXG_dfZ+T5OUM#2HO[C,Ag2@^.R@=/GRM>d\0M_0-U?7
M7a177#H7]X\fg7D]:Zg,NE2)87?:>+@;KDM1\/+R\NR<1EW3#:53T#FK/Qe\=:+
^Rc9Q:@[MXS.D<aeAe=SAI[F/Dg5B]7A\W,XI@5d&]S<decU_LE/g)IBf]MXcQM;
a00BFD#LW\R9EMcDY?Ea9V\PA,MT]R4@HO4c8Va[DIT])2AJ\S/QZG,G:MY\Kb>O
+_Nd1[8I()Og@90/]=Z##,6M;=cO9IVCOSR=/87Z5)3cMI0N=c762U5^D<cK]ZBN
H7)]ONRKNM\8_+eDC]TS;KR-&c3YFF/=]ec4aM5G,e&e/S4A8I_C/N:Nd\6fG#,Y
+F-?DSaII#M6,bEZ2JGN2^[U<#<B9?E45O4a<IIbaBg/JYd?BA@d5Ra3Ec6+KYWO
[N#[@I7GYD1:YU+/W0V?K:G5[]2?>2[5CRg1_5aW](CVDD2-C]CbRXSZ6NZ:&>40
E;b&ZHW==#H<EH<cPAKF+P#)\15;A0\/aQ#CLQU-2&EZCM\9^\RC,]=+CSF_BYZb
?W7&E49gQeHNNRMJD.:&Dc;PA;UN6--WFQW7GO)0)P=a?c]OUY;b.1[^+1gZ0f:N
0X?R-Z1f.5,IJ@.dQ/T<R0aMM<3)/GR/6+&=F<J/f)5c/S=Ecf]eNg?+SHZ2,&b4
.@5VD=J&N)[\K+AY:@.+SY@YfF(+P8O]XeT+W_dZXDE;(<NT,0_)O@+\UPH([D4&
X1e0=\FF0LEc0-^#V/V0F8RZF]W6&3NMHNQ[aGf[//FL,TY<f(b]Z/#cd^QD[QeU
1OI08HC3[#T:4[Xg\<Lg^?P(bMMJ&YUS2T.XH+-1S=C00f-^A\??^P29O?#R_;07
d9I,.J\<8\H^b))6OdITFM;:&]9?@H9W[C(9DX4\[>bAU13eXY)f)MYeU1eDG7)-
F?__(d8S5PIc[a0S,aMQ26K=91A5fU7\WgO=gZ>[LL<;R[42BJ.A4/>CK.0XW@H;
1#7K<-a4VP<g@\98Q.a6C7_M^HOG21a3^J05S;Z:8-9acPCX4PWW3J/ZL12\[P\U
C,H^PURZ,Uaa4b/&V)6AG4g_T>NH;c\5U5M[eP3AT#eKI2Cf29+\IL4,?,9bBQ8[
T+.-E=e]+XESRI;c[]J59=26U2bJ#ca-TaL,X,b1N9?-DKC;,/X&_=e274UX88Xc
\;).2^(-8ANa)9P_CB5g4EGP.MF;;IT/L)D.C@WVAKF-\]dLbMSXQ>GQ^77@.&B+
gR>DS;U[-;&PPTA;C-4P[KPG3EE6+5^VRR[N#6D1cUd+^M7HG0g3]YSEO2\?4\0_
=A&>FC)E>.-]G@[eTEMA@#@J)?b@+\A3aF53-:OL10;51@Jfb^41.bWV&-K?1G\V
\eDXc8KfMaR;V)69A6,/1CT+Y[GU4bd3:LQJG3^LL?8[V0#8O^5XB[9GQG8PG#Ne
:c^RN&95V)+QggHD<5=2O>Ya;-D.gF+=.>?W#gWbHfOZ8cN@6SJKO_Q54G:Y2&CF
g]<:F^36@a<6<GRP&7E\FR9KSb6a30KN.O:cM.-;[)OW5X\S\6NGDaDV9>T&P/B]
:;+1NLQ_D0d8=JGO3L-.3@5I=d9+SL5[+/f^JCOgX_DAIYB,P2DMIS(LI5_K/PY<
8Y-DK]Y=>aAZDSX6H4C2.\V3J,5&?S+Q.2eR-B.YI3DEcgWDKQWTeA1(M-1,+-Bb
5d#G7>D<KJe.X35DXO9TL>)BF<UE.TE.]D1+0MO7=G:63AQR3)3:=&<g\^gU\&cd
Z0^F\O2IKZUCc=?EB(@(O/Y3aTJ2<SO6A;,07J\#9)<;_[HQ?9&<cLUfH=f/OW0F
=Y)U6SK,UE_]VIbS.O(]5BINB;<;:aV8\dC7aJ5-gAKU/,O9^]#VbU&QEO18&.JC
Q=a52-9M4#=V?K+9<5>(2@3]US5[;]B4/4@UU#:TUM3Ic,O3[L>Y0a/aXITXXS;<
Y&4326]S-]X<R_0N&BQLVD;,UdD>8abYH?/KBG;UK+KNfZEC/e)Zg1cGGdT5Q&dd
E#T7;Jb9RC6aGS>c\<;<Q^0Rd?GSYa\J^g.?^>]=A_<Z5Cd?[T/cQ0a_ZSXcC@NV
b)^_KY>LAUT2A3Ub6d_>FRIO7\[9;2,[eCfVQY<?.@)NcFY&W,5-I>JUW=O.VL]B
QN^1GMgf-(R<)?P\P?ccK\P_<J,fJC;?gBUKO-C5NF&4<4BJV?SP7FCV:5e\PK@Q
_&64g48LaXaEA[=KI#KUX_U)d840\I5P;>4[0fDU&7.ML&Y<b?J<ZRME<.HT@:SH
Xa[6WT_UUAZdD_3LS[_Y0U@\F(UGR=HHeYMQ_N?;_bH0))P?8)W5?Q1bf&3PgOWf
^RN[>)T5=#LDJ0VEOE7c,FLGC9N6(+b_G=I[S9+&JA<XVc(8&U<L_92e?]WL=4,3
Je-=XSa,CJ7;OKXM]CK@g7fHf[E(B,JPFVdOcF^_0,\0.Eg:?+5HE_7?>/K(3dAU
;5LefXX)[eV80\UH.CF3EedS2(d8_aPZ3H?E6_V752VEdJB5<.1FSWACQTL-b_c-
DN=BEO&_-W2aP(IXe:f2<W:K,+OU98:^1DQ>@cI#/)e-I0)S+XAJD--KBEc,O&YP
#F@&f@/:#^=9?JCPD=dbH&,B][@]TG5KQdRODY+MfYP55EU5?PLc]N8a6Y@;Zc&O
-2@a&4Z197^cQ&45C6DaN74/ddGGBa4c,WH@[SOT\eO5+HdPRT/3bd-5c=R&]2Y7
B,1T8;ee^5D2W/DAUB.N>,EO=[f37//KR^KSI/F60,^+aWMHDHg/[Kc,TMJ4GZG\
a7Ub@(;7C.C[4DB7TQ42eOK]fC>Q+KGRbH;g;_S4;RR_Q5T:c]X_2aFJ2?.;V4Gc
2F./)W:I.;>R@a@I_ALI1Gg+0H#H3FXbQYQT;WB9E[&<U<04<H+=Z?[]e:67>9OD
I[eZ=&9c:Qdf)Y0TRRB;NUS-/:^6QEf.DY-D)Ra/B)IP44+CJ2M3Jd3,FYM(f?(;
XL430?+-8a\7P\]g[^OH7db&=C-&<&Pc\#(_GRcHGZ?@/?Sb59\H[.60ENGO>]PH
@#&AH,JZb&=RWZ1+Y5;Q5FGeJBQUF-eZ\;(gE,;P7\B=\@OM]<G.E:Ya;eEY)61Y
6/c(A<R.PFY=FJXUC0911bacfNB&]SWHNZD.V0.@4>(0YIS=bS>=:HMY/^1Q8S1W
c>@(IL)0L6SJb;6=8JaJB81X\=5eTUcJ#5+QD+a0-KcEfV5]97]baC>UePP46caR
+(FY2G4#>:MBWCEc6H\+O&/F^=B:UV#Kb9)WW18>XUHf4DCe/-B^0TW/>=O5Ba0K
^fb=SgG/^U6=8#^WLd3\C6ZO?6C;d>3G=eD3eO-S@B>WRUO\<-TWO9#aHOOc^5Fb
].DIJ</I+?UTOb57PRBNZ>\TLRY<114NW3Y>OZ\V2GQ43WGP,KBKfNgSYAROF?Z1
].-BMRZPJ2I\GAA)<60cYD2<bOH8SJF?CSJSTH(Kb1G9[Ne+<QJ\IeN>4KI2X07G
#L<PA_]+&M\I:]VS-.E/I(O(E<X/CD+:(-e3@P,_fCP&#S@b32WYBHK=(MbK#3g+
N(b(\@^AJfAV]^?VX;a7YY+6]@_cR>eCd^?@L3ONd[eOIQBP_e&ZFH_K=Z(/53?5
7?_5RgeD9EUQUYBV=)Cb_LI5aeBUX)bEDA:;R#K?AZKEFQOWCMS?8&Q-#-+A=M_X
746PH9CO,J@S_SWL7\/#/1f^.Hgd5^,WWL8J]2cHTES88DQ_84(1=/B,\793dJ83
6AK&7FCZ7AJAI6gB[;4Eg;Na_^0D]+cJ>SC7e&c1Rf:1M4I6_[MYDegRQCc5#fRJ
6)GIV)SaXAAFZ[)MG:6VS_@67aU[fH[gDbRB@G90Hf^_TXb\5g.Ke8E]e>#+,fC>
B@S[KK<ET(P_Y)M+bF]/<(+LYZ_FO5316X1gA>^7O3?=ULNV(H&1,JC3MW.JP)@9
Le:^<0eL/XAZZ>&D)S-9c05.Z(GR-G\@IK&B27UP<Ug(RW0_G,V]/a(_W25J#6Lc
-8VeTaH(f]K.G6WIJ->>+aULFfb<./@YE^\cTc/7@^:ZYONKTdZY,-]&/XNg^;O?
LQ/&BEa3Rb__R9B@Zf)dKU7L]#ZbM/8=WBc+II8(gXR_^\a5@d\PM3C>5H1d77&W
#gF/Df),A1fPAGJTTF4J37]8B?[A#>AbZ><eR8(:J+/bKO0,Cg9JQcKcVY6dPOV)
;>M0DL85@U(0Y#bV]g7&f0ce6Nc-/-IeNK90,](g<)<ZX@^f4;I5YJTP0+#<1;:O
T&SU#ad)+OGT_20;F;6PEA0ECE0[,G,;/V53SaPKSJWJ6^J5F[?6\gOJ:e.U-RA?
DFNCeK7C+KBfV,EPG;B)<I1ILZ+S#47L^GS>0.7P,E<6//)Z_LOE&/H?b[43EN9(
^VRB1PPG;VQ)/1bI<+YNWF^DfQ-E:e9QKfK04S<+P28X@?+7Q&+Q1g/33Z_Z4Fe/
=3Ce:OG96:^X&&?fF=A;@VJHg]2.cQfJ.QI:-=^^K4>8<8JMSPUa2QLQRB\CYeGA
9]FLfI0]T\XTH?S7CfZ-<HE5SRTRg\b4fbV0K)UD+SLSBFGY_6DNW;YaaeXI5J0Q
\[RQQ+E]-bA;)TD@5KNUDMBMN&KSQg<7HG@6(74MF,&@/JD@:g3\bKMeK4&Z<N(&
/a#5]SMX.<<bf0E.,d:c-Jcc\dO?4[[WA#GSS]W97g(Z_?/Q@77JCC;404R16PL.
4Z:(0]LY7;WQ0.fIV_(M.+CYG\3V8L0fb/@G[N4]NQ[+FNW<f?BCXbT)AU^@W<9M
JAg.dU.ceHW1+-F4D)VJf_A0a)WVF/0:IZ:>WaAb^,;0DY2J0>EQQ7bG,AA91/O8
?ZeagV2?gP?bP>9f#Y5+@<AV4KL_\1+Ff]<NJ4Y:Fa5aBC>)F+UT<-\_XE)d9Z?6
dUcWQ#Q5aL\b3DY(#,?gN6dQ9/(/SA[0-OFKf_Q0_4BBcEQ2Sfg>RL\W],Yea&&>
E.MSMC@CQZ?;NP-7OG6?]49/M:gHP3A2D>E&H4S\ac0:TRd1WXYXag&10C^TeGM2
[e8;@LcN&Q.[4L&SWD7+&[GZPCf//<d_6H:7KFZ30>FA?B3SJD]Kd9bQd-cDIAQT
\LT@E^=eMc4S9a\WP9:ZX;JYBD96IPL>WO/M+11XD9,Z)[UEV^>H:-fDMIAf#@L9
453B9b2W@Ta9@G[]JHHf6:ac_;XM\Wb(3/#-a<;HfYKQXHa59V]a^=Vcg5HZ>(dA
&QQ(;K8M6:66KLCOd(ae5/EV+Mf#>;U,/e\;DV&F?D7WYO<+U=,fK_](FKe/FRNP
N\--&[4V1Od_dDV;_//_F-RJ3Hg;1):E:T&J\(J^Gf#.[87Ha]O.G=SUPAK3W,;J
98?M7QeIeTO?D30(A71b3Y7?>\,S4f5UMQ>(1f(HK62PcUQD?d6gSaEg-_01,><4
f?_EAP4f[,U7N?>6N7])D\7f<aXF;L):7,+@9IY_NQ=bAHWH84)PQM3U8]M5]0R<
@M[0+Q8B;B>Q204/QV\UJR5(8X1885(LX>f;8MW&/&>3fed,/UZHNc:bAQ5YCPW&
a(X;E#IW^SALJ8SL821T.c+J<Cfg_?-)HU?1Ag]>=K/Q(+?E01E(KR(WI>\H<(HD
_9D-L[5:[3E<0d3YU:K_Pe<Ab/fXD;^;eH12HI/6a.9TT0-P,07N\(+1NZK,\ZD#
<Y<N)Af,V=[a=P),N@#LL9KRaGM1F.Q[HfJX^d7d,SO#Tg([RQdSP-@bgY^SJc+^
]>_W(d_Y70g_;F0G]90_Y,6@@5Y\@];?EgS8+0KZ^Q1?eI4)Df:[22/ETQZdf\a=
H;^<NN45e+#D(,I1:[YAW-efB:UPG4DZEX<)_7[L3)bRR;=&7TE.f#@LARF&0(RH
TV:(1]&T]gX5f20?.AN3b]WV5@A?;;[VEX1,J>,31MV(2ZH2R>UC;XTC^C)\KGI-
/1O)Wa&]=WVPM,=S8g5K6M_W,9MK/&C3,bW_7WdSU+a=:(ET4DcW/<d[=K&DaSfF
Xb&YZ(b&VYQ:)B[P-456ROg\@d+5@Z8\FK]72_08>Y8:WKNY]6_&<B^Tg^dHF>IA
UNP2O4H:U+TMO35_V,UAOKg<IQ41J:f_gc.d^BcPPV&D:4EVcMU?[9Q.Y]Z62_3Z
/+4R@+[L1&a34A8dZfeB3e0X-IbG?YF[Z6K<P=1.L/1G4>V<_eOe##VRV?XW(L[I
&O8+9;G3<a#9ZR#L?[2R^c.U6A0Z]PI2QN7W+MFPeDV>Y#-[QEVM_EC-0?B9#GH&
J_+X&)[I#d0+_g^4S0\I=0&/gZCV3Ug)b&EG,7&AQF&eK#I2(I?-;7QT_e[+I9c&
7&S#Z-e<O9TXfdeDYY;HgDgGHCW)7.Ed+G_>2].4I6Y>WP9(a3@:@5OT_I]+;cS&
S>YP3c-O3>\0(:F,8(#P9c6;ZgR3ZZ@]=HE+f+OJS.D,Ob9ZX9L28L)\3H\PZ@^5
Q#,#SeR5Ta8:78KW&BJM?0JYa84BTFVO<fYHY9^8/e\HO.J_=8/8=d.fQg+8RH9@
Z<X9YU68dUO)X=X?;\0S6MG9[3.>e2XW>R31PBV)<EO57H<@SQIb6V48c+=S25Y8
5N+/:LBTUE&VG9af<_#[_DHPdZJMJ\C@=#6F4?:@_VQ49eZ0@6^<<B0/^#?WX,#1
XI(VQ15>L=TIB3d(M&?X.T62Tb/QA;Ie26QP:LZB9]#]L-F5_Gff04;B>RL,]+<3
R<TccBYEJc7@J69+<;U^QN4^1;S-+8(Z#5I^ZNNNeLG/W)+:87_NG8+&)g[TK<8^
bH-9DI+^GP&C<M9@BG>M+MeZd@g&S_gdg^D.cfY)TEESI5#:TgQVN23N&d(B5S?b
8PQYLMIOET.WMVAEfCCTegfH&;FT4aORE&_/,abRN]VXW@YLZ)aY-(_Y>\<2c:HP
8S?;a45,KVIa06:eIH:-cK0^>M4,\^96X,5NTF3AI=^9(9X4bb>79A05(FSF(\D:
AT>#Q()8Y(A\A9XS&_Y05Y[6(NOHGH-DgN=+T?=MA_50;g.#=1,\&H.:;3+cTY0;
9]dD#QUYO=\JX)QGc.e?KLf2?^E&GeRMd?MYRg?K:3?X-7F4_IMB3=:NJ[.URPZ^
Sc94^T#0^<=_@VQ)F>^0bCAGf+BJ2;Ed0&0BN?I;/#-#ENd<IZ@J_BZ^6XY#IEe/
EEaZS/N8g(WJPAbN;,/\V3GY@e<a5YNC:@b3GGbHQ-,[(.3Gc<HfX,C\-GeTf-_V
Gd.S;&baOX)WCI62d.7B_ePQ1KXG^G+(2cBJIY.C/WUBNX^:@Sd65XQQDZSX.MbY
Dg>8&M<WO1:./0601=TbGN.Ff0e3F<)HAHZT(/0D33AUc=Zd<(;:d,U[ZRH_c1.[
HTc0?AcP[-Z_Db#aZf1;gQ@)R>H6gL()OU3E@H9DHWI&?&e)YT_]:cCTNUY/VN>A
AH.d(<MIdI4?I\O8SbeG]6WPT[Qb8GITgQ/U3>:?@(M/9OadUA@PYOgDA.,BO6:#
aZeZFANP4Q(OJACST)19A[4@5DMHTVCZ3++E/.DdLSAA]=YVRUILW>IG\MR3bK/3
[;L3TP<ENWLa(X3U@4IgZGHBQ]RYBXZ<:M;,K0)a#CA@AfdCH@>]WHIGN$
`endprotected


`endif // GUARD_SVT_AHB_MASTER_UVM_SV





