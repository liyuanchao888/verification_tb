
`ifndef GUARD_SVT_APB_CHECKER_SV
`define GUARD_SVT_APB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 *
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
  `protected
#^ff1)g&69Fd.\C\a;8D?N?SR97W=3^],E@5Z8&Z/\5f.bT#G)>#-(GO+,[^;HA4
^ecH^,AB#V#I2V/bYT_J5:X:(U&g[b+@7gN1PQG2N9Z\C#:YM@E,U>egL+f2O#GO
\0M-0f(Dc8#,FLT8eSG)(9__3(7(\4f4QY]VH/6QQ\+Vd/[PHLQ-T9d/aPT;_><9
Mc-P834a,F&C#VNM(</Q[Z+,/3^.MKDH5L75(&<WP_L8[]EZg3K/Ue&\]L\G+.S]
:AE6_D/FgE7,M^Q2HGa7bgO_.-:53OV5\Kd?646fSDZY6^H=Ba,)I=g)aF04:gHe
WHF07U6Q5g)[@QgKS@1)6a.fA_99)2NV@3.RKO;1_:ES2a3ZXZ/K#W+TRcD42gPe
GO8G=^>R:(@J5d&[=Q_&Fe.JG&F@Db\7GHBBLS-^8#NG&fPYLELY-7e0@1E[\c:M
eG/EKX^82ebJVS@cE?[Y6.Y4MVe7SfIKG)55;#:&QVf-3_^(_#\V11F;NO/R]>CS
;.4#&d5/,MOG;E&6HZ_&4B^N5J4HO(HU2J@dLVd&g=90,X8Sa0&R=Rf4aT:\C5Q;
.;UU+(4DcZM9RJTK_#OH9EU\@gUDOXP/LG#Z&)NC(\TFPAW3GDRB4BNMgFF&HC,^
A].&U,0#\MU[aZMb8:UI4P..(D/Z>;@/CI(1M7)gc)XBdb@Q^(c=7XV_,>+Xf&,>
e7gf6L)]N[GPW7dS:C?@#D<^,C@^J_NOTGS^V=W[8=XY[[]A=[-S[^<\(>>_^+Y,
;3NITIV_6<P&8fAKe.g/Y/b]RD9-PBS>(/43+\J\O.VMDN;_<3DF;HP1a#gH9]A2
f^YbHCO:8]G;eHFH^BUJg3_K[STCUa<SdU)_8d_:=<08^(PZ58RfVKb\a\Fe#-GG
?,bf3VHM,Pc3EF21d4b3W(UR:O@5\8\CbJON+6NOd,@fV;IYbLdYJH.D92X#H5M@
aY^UScEWS4ZPS5:fYAPXf#_=-@G_N/#?-I1f+I)DLd]c^6>)SXc.1>T7B#FXg;)S
Nf&HBVI>:Y=VcM(M-TDUD&f3-L7#QAeFPT.2e3+1EL>WLYfW8JII-5+QS#[(DUIM
B,\D7#]f6)M(D.SRR^7_T:B;Q7Rde5B66,#FAIU/0-:7(5e4D0?c17G>YVTV<JUX
G8?82^LY3V74[@1WQ>YX#cFE3b5IfP:D5E398T@Y,C6.5R1Ibfc]Y)Q(K(/T1-8g
SX&D6OD/D,,BWa/H?NaXT7c7CXD/cH(:UCQH5.V.WHZ[E,K5B:32@QWg8Q;H0HYF
3fQG](5\[\A:]ZE8fgP=PB@c-+0eCNUQQYHNSF4:>#8XCO;]?N/C5<9.f.PRD-O+
J)1Ig.(Z+K/ACa+ZY)Ea&2S:GZ&9RW.2.R],[^_]E2_Z.dZ)-gA9dV+fK3<41Z1^
?/F0?gTc=Ff@eDAKW[R,0LF5Z&ec0\a8E5YK7[/RISCPSc4SB/6]-Wb&MD5_Y:E&
+GE)MEPIN&1/:TJ_T#;A]<5)R^BS5XOCV0IB2,_8-g29&#8/GP;[a&-T)Z&>)c@c
eM1E5#]:Z.aW4^T1Z4(<XK_\BGJX(g&QX+QLHe/2b1Qf9U:-@R-ZIL8I^1Q6@GE&
WM/.2R&Y7L\B&e8)cbffX_LU2U1?eWOZ&aGg\WA_&RQ]N0Bd.Xe\[XS)8^f99&4>
=B>S:&H-[A,.(I+(gX_[D_WEf=7;;0ASS3gGYTQf(VWX<INVXMRdF^g6#J6+LWL[
L58b;FPG40BV4aKH;>&>SNb/,AQ)DE/:^-<;cfg-gP4.]C6_gXLT#b+CH\8[Lf:W
S0A=RS3U^S_S>+7(8U;VV]RBKQE;/)(e[AMa,[N;>0;-+dQQ^O5)WX1SPCaLY)eH
N>GPV)g_2=WOBO<JZ>]VWA;8Y+2#@7,Rfg2;;_JXXA[>124&6AA/3gQ6[c<:77Ve
Y/_D(<&YKHQE::cO&C-H:+-d5:AH[bMXY[/g683<S5^YLLa\UA35_XJ=V8A<S(]W
d(3g+KBN^A15(E>8RV-R(1C@\GLWCWNNSUERW0+Kcf)<@EU:fKAH/L9OJ1?\4;#_
KLWLI1OFUN)=_3U)33T1X/]<Fcf2&A&D&LUa,=>J9c/4ZT+O1+\O/FF2=,IXaB9:
6FW-NF7]ITQ0<>1]g^20_QB(bI(1G,K=ZF7c6M6>J9V:[^bR2PUGBGIHO^,8:E5S
UU==2Z2M0B9GUJ4M_E&7IU@239#JN1:BFGCdK/=-_OFM/8&Fd3TM57XKQHYL5QE^
TGd(IAg#1d@(aW(c]\P?QHJ7X4(Ff7OAE,0(Q>E12KV]^;^[&g^S_K2):I?,U?13
3YE[R:Z<Va-VgY;?/dI#YW.cf)#(>\2gG#^MeWP=WPB:12\edIR=<RYX/A1C\.,3
4=a)JXW53C,>9dDgU?KX0dgJ==@.B66PN7Y#YUKDJ@C:a1QbW/_L5M8GG^LUHPZ/
R,RQMDKUKREgP2?7,XV]GYe;#>AU0@OS&g)BXe3g2CGX[)[?b#gf<L]QG#IYgW8,
\O/2+QPYg_=RBO8QVF=>,LS)BC5__[#B(8aa<4M2:P=bad4>QS@GBYc;XILB3Q[0
9)4^1F+=4<V;H7+,EQYPM0UbQ=F9+9:.@VDFPUfeO0Rg^,5C&I/#EB?^@X9CIXWN
IOBL\NG?..@HAd>7+4CLNc\2==#a0f/-A62ZdV\_VTP;_W=AQN]XgZVGf=0fEL3O
CV-bg,e7Hcc,Bb0c/LSHf^_EF/\A3AKQPf-AG#.b?c1?C0+fLVQ7N#3ec;9&9K6C
ZV/:RILP)c3Y.gLXdTUBIJ1Fde,/HEA?7-4Y:GaAg;0L@4M&HT<DD[a[7[S?:fQf
-7U&7IPeg&O@=f2cL6:4)-1F1$
`endprotected


class svt_apb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
 
   
  /** Checks that PREADY signal is asserted by slave within timeout period
   * slave_pready_timeout 
   * Group: APB3
   * Default severity: ERROR
   */
  svt_err_check_stats pready_timeout_check;
 
  /** Checks that penable is asserted one cycle after psel
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats penable_after_psel;

//--------------------------------------------------------------
 /** Checks that pstrb is low for READ transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */ 
  svt_err_check_stats pstrb_low_for_read;
  
//--------------------------------------------------------------
 /** Checks that after reset deaasertion, APB Bus is in either IDLE or SETUP State.
   * This check will fire if APB BUS is in ACCESS State after reset deassertion
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats initial_bus_state_after_reset;

//--------------------------------------------------------------
  /** Checks that following APB control signals do not change during IDLE state:
    * - PADDR
    * - PWRITE
    * - PSTRB (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PPROT (when svt_apb_system_configuration::apb4_enable is set to 1)
    * - PWDATA
    * .
    * Group: APB3
    * Default severity: WARNING
    * Note that this check is performed by passive Master when 
    * PSEL[svt_apb_system_configuration::num_slaves-1:0] is 0.
   */
  svt_err_check_stats control_signals_changed_during_idle_check;

 //--------------------------------------------------------------
 /** Checks if psel changed value during transfer
   * 
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats psel_changed_during_transfer;

  /** Checks if paddr changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats paddr_changed_during_transfer;

  /** Checks if pwrite changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwrite_changed_during_transfer;

  /** Checks if pwdata changed value during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats pwdata_changed_during_transfer;

  /** Checks if pstrb changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pstrb_changed_during_transfer;

  /** Checks if pprot changed value during transfer
   *
   * Group: APB4
   * Default severity: ERROR
   */
  svt_err_check_stats pprot_changed_during_transfer;

  /** Checks if multiple select signals asserted during transfer
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats multiple_select_signals_active_during_transfer;

  /** Checks that bus remains in ENABLE state for one clock cycle in APB2
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats bus_in_enable_state_for_one_clock;
//--------------------------------------------------------------
  /** Checks that if illegal state transition occured from idle to access
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats idle_to_access;

  /** Checks that if illegal state transition occured from setup to idle
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_idle;

  /** Checks that if illegal state transition occured from access to access in APB2. In APB3 state
   * transition from access to access is valid transition.
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats access_to_access;

  /** Checks that if illegal state transition occured from setup to setup
   *
   * Group: APB2
   * Default severity: ERROR
   */
  svt_err_check_stats setup_to_setup;

  /** Checks that PSEL is not X or Z   */
  svt_err_check_stats signal_valid_psel_check;

  /** Checks that PADDR is not X or Z   */
  svt_err_check_stats signal_valid_paddr_check;

  /** Checks that PWRITE is not X or Z   */
  svt_err_check_stats signal_valid_pwrite_check;

  /** Checks that PENABLE is not X or Z   */
  svt_err_check_stats signal_valid_penable_check;

 /** Checks that PWDATA is not X or Z   */
  svt_err_check_stats signal_valid_pwdata_check;

  /** Checks that PRDATA is not X or Z   */
  svt_err_check_stats signal_valid_prdata_check;

  /** Checks that PREADY is not X or Z   */
  svt_err_check_stats signal_valid_pready_check;

  /** Checks that PSLVERR is not X or Z   */
  svt_err_check_stats signal_valid_pslverr_check;

  /** Checks that PSTRB is not X or Z   */
  svt_err_check_stats signal_valid_pstrb_check;

  /** Checks that PPROT is not X or Z   */
  svt_err_check_stats signal_valid_pprot_check;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
/** @cond PRIVATE */
  local svt_apb_system_configuration cfg;

  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
    extern function new (string name, svt_apb_system_configuration cfg);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   *
   * @param name Checker name
   *
   * @param cfg Required argument used to set (copy data into) cfg.
   */
  extern function new (string name, svt_apb_system_configuration cfg);
 `endif

  extern function void perform_read_signal_level_checks(
                                                         ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]  observed_prdata,
                                                         ref logic                             observed_pready,
                                                         ref logic                             observed_pslverr,
                                                         ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                         ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                         ref logic                                    observed_pwrite,
                                                         ref logic                                    observed_penable,
                                                         ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                         ref logic [2:0]                              observed_pprot,
                                                         output bit is_prdata_valid,
                                                         output bit is_pready_valid,
                                                         output bit is_pslverr_valid,
                                                         output bit is_psel_valid,
                                                         output bit is_paddr_valid,
                                                         output bit is_pwrite_valid,
                                                         output bit is_penable_valid,
                                                         output bit is_pstrb_valid,
                                                         output bit is_pprot_valid
                                                       );

  extern function void perform_write_signal_level_checks(
                                                          ref logic[`SVT_APB_MAX_NUM_SLAVES-1:0]       observed_psel,
                                                          ref logic[`SVT_APB_MAX_ADDR_WIDTH-1:0]          observed_paddr,
                                                          ref logic                                    observed_pwrite,
                                                          ref logic                                    observed_penable,
                                                          ref logic                                    observed_pready,
                                                          ref logic                                    observed_pslverr,
                                                          ref logic[`SVT_APB_MAX_DATA_WIDTH-1:0]         observed_pwdata,
                                                          ref logic [((`SVT_APB_MAX_DATA_WIDTH/8)-1):0]  observed_pstrb,
                                                          ref logic [2:0]                              observed_pprot,
                                                          output bit is_psel_valid,
                                                          output bit is_paddr_valid,
                                                          output bit is_pwrite_valid,
                                                          output bit is_penable_valid,
                                                          output bit is_pready_valid,
                                                          output bit is_pslverr_valid,
                                                          output bit is_pwdata_valid,
                                                          output bit is_pstrb_valid,
                                                          output bit is_pprot_valid
                                                        );
endclass

//----------------------------------------------------------------

`protected
E(M?E_5_V2RQdbIS3U<-H^G\KE[GPP)f+7-XV-K18:R3KX@c,:Q#()9?Z8fSM=[1
8Ve)-)L8:?-V<8=^fJT1W16Z>YR#@J0N2WQ]N_9Q7D7aH;bcVS?F0E;<2B+7.LUB
1\M7Z/@,gf@E+8/f9,]bJg87<S6ac8;bY?N6bc@SPD.d0D:H./2g-VAK]3A:_QS[
b&R[+SA9e.c_S/WFf&BaM&E3_QTH40cKD3>\YEdU4<YRT/Zc\:R8CTAd9Y]^RGbR
7;^[Cd\,5#89&O#bC7:Ae)EEOe5SeII?^E-<_e+a);NQKcgeS0:g-2HZ&:JMZZdb
UY7V@1(EfFb<VK5UBIO89ODT3<bccC_XbbXE.9d4YCbD-0RH@74S-O(5R)R+E[aD
2edY0EHKJ12APdUa.B#MN1RJacSLfF:M8ZY-[-R&R\8G_;dG1YQ(-W+^T.7Df\5f
+E#L#/RX/HD0X5UV.:FR,>ECI-#_?W<bf1F+)J8)GH,N:N\+<A2Hb6#?a?K2\4_R
+YY?\+\IE@/Z7F4,g,;cREg/VfIS?MYfCUAd<#LI_AV^-@9+;ZN9/0bWG:@\/GQI
SUA5/.(8?D7C&Ye@9:=(.BA48?W6g?9280g=QW/+;HL^@d4Y89aA_NS\,V5<a+H_
DH5-@ffB4Q5JN:cL8.+:;U&VW3N+=I5:WM4UE.K>MMWQe),\TX\)(@^.+;+F1Q;e
ZR,60S?ZQT&F,4fAd2-c&b[gdU0f-<&&+,OgM0&-S[JM?ff33gOa&XMWJUd7/XB#
BKFKQBL]-/KJJ?NI<@LXUBWP0<:=?eW<T9(>61NJ9T7?]@/F52JX/F\55=ITfAJG
PSIBEdCSIE9:?\Y/7VdWFf&W1Zf(?J;^V5d+,b5L42AgE4@,7M?#KZSN#=-PcBFI
^gAb8HeW]aZ0&&@D@9dZ3PQE^)9deU3:\:K2#+T&(@QP1DZ?MI(3aY/g=?\aXd=1
HdZ[Ke;1TW.e+00d]:c<(\QH429S?HA6IVaVf;T#VUBMBDdSHM@OS=3Z8,CHR[6G
T:6g-2Z1LB;aSBWT:]F<O]#VZRA.8L2McL&;f0)#W8F:\g.W/a.c(A]54E_9Q=@8
Ze;O4B658L/)FN(^fYG,M9HJ,^NNA?D=Rb4bP+;.M5R?FYIM4ND]dA=@2)K;?5N2
:2EH5;Z]Rd[7GXge.&Q;A)/#C7c3(QL7NQgM.#@N;W\U:2_3WTR[\PI^)Q[/5)8H
-7L]+&[S/J73JQM,=Vgb_3=740bML\U69TD6&3]/gGXb3I(#SKPaJK>8H1D)eE4f
2+[U,/#ZbM>bG<Qd))--YMTF3bA44LC#V0Fc[7A#V:fYHP=/71dA;L^I-\H\WgeY
FR3U]&WT4Ud@ca>O?_EEWB=/.^fcFZ<G6IMfK9258P1\9E/M@X,BZ41Q8T#3JRNZ
VXfW/][)C62HbIdU2O-edMLM#c?Y6>1]E_8JaDHe,YEYKYCE6[N.U>FCe3OG<B(,
Y]/0LMRU<M:K<0,#Lae[MI,NH@IISE#&F;.7eUKB;DA18I:/;7#,&:.P-/LQXdWJ
F)NO\2Q_/b1XZ_cb\#dVeW2@e3([Ff1b-a:-6fVaK_>IFaQeOF[KQ.J4E;ReR9-;
?RQd:N#EW+5TZ;CC@1N9]YP7(2XOCccabA&gIJ^^/Q;TS.OecG#U+XFZ4W#b.<.b
\eNQH5c/EeF.CUWQ4O_1Ha^IW5bC<DJD,+0/0ZT&[a=,LcYTb[];ASINH2^Z4D]O
R6:7BCLF4A,WI?;R+ZE#\7dC=YdW&0U^B+JULOI&X0NGTM^B?^B=)(G&[dZU6X=C
WADR&c.2ff,>&FOfUZK#;P33F4RbH=I2M&EWNG6<JMI-?O5(M0Be&IOQ;_Qaf&FR
\Q6fD:=(#8C\2S=.:YbF.8e]CH_CG3>=_fSSKP.RX-&_NBfKIG,D//5_(Ba(51>+
^:_F?P+BX\cb#=[-QZ-g4JR_V+OL-1afgL=G5Cb,3;&1_W,X<[^=/;,f)XJA=+TN
aF5[QXFTbce3IU65GXgdD/5S;SBL?a#f=#A?N,+8bUT2A4Y>d9?3\#UJL1b&14D/
(\g.4?7fT]IU2EVebE433:FD?H7DU]3e6aH9,/>_7Z1Cc?AeJ<;N,YC3#;18<#6I
GIC5T_-XL7A[&9Od(H43.3^3_;HWe=]#\K_EVW-2Vf_eBP0UaKG@3-+N2J;B\cI=
Ga>d\1ceM24IcC43;gb2-4G?D10JBW=84f<fDN;(A64(I2=PMG(PN>,+[L2#Z/B6
9G9bB:8=g#5PaTT,=X5#76I]WG?2)EQJ5L=2Ff?^e^;<d2OJJ(O8/LC2E0NJeQAO
8##_UBYICB^#)8CQ<5cGVfF0?E_D(-Q=90Q;cJH<ZPd[RV_Nf2SH+5W/]P^Z4&O#
JV]>7BC1[@JAQOUPVU85GP2]b:U])W9I:QL1DX.V7gdM\W=YHG,G:/-)aaXXUI,P
;9TPbFd>K&2S<LW>T47FHY8f\GKF=RSJQKT0eX+T=de8O)>Yf1K-@Ua]VEO(>Fg,
DZ(03D;,EI?ZCP[gd\T;@a9=5L6g8WAZ&;2]ETQF)IcI3[->IW3H+VMYe2/W)+-b
JUG[<gKb7BRX3bBBP:QbDCJ1f&C4@JH>>M9bV0^W._#a.1bbE#&cD<,f]NbdQB@J
,c&PT_8bPTU]UIdf2ee\/HA@S018WacQKYT/S)C+a8&C7XdWa;[W,YTaWKaAS90;
J[D4^ZS/9MKT.&+&R967ATAT@^4-7)?8YFQfVU<?4KG^X/(JP#K>MeL50MUDCWN+
((?0f/HOJYc>X8^T;)2FZRHCfIN6AYgbKM^PP/HS/ed_LdFT0N)S,,F\f>PdNT^/
IF\79^DVIHKbJHS7ZI?_.+=;W19]:eN=3BO-XGd&4fCSMeX6aJ<HKD#bV/U8?V7(
A(e6<bGd0cAbZQO-Q6D#LGVS6-#L.RgFFTZ?W<LIYJ<P83RJ[^_\5>6+:305F:bB
b2;(/5#,B_Tc0)=6ga.P[e7J::_BPAbZMVL446)+&9_S:5\?L2]b<6WLU@aVbg9#
&.bS)/bA8S89QW@:E2T,2I?E9O+;/KQ/gW,:RXG,M^GP<X==BfM5YeCg0bPD@33N
-U<^b^O)\SPAQ6&8Y@Z^3e7T+PNZZ&D3.S7Q^R^2LA(\+_fWc:9#GIMN8=NX]P#<
aIM;N?/@<N=_(Z<2.I6Ra+ed]g7U5Hg@D0+R)_:?cMJ@+a.47];9U:-/0,-AE(N@
(F83;6[Y=2_9SJ,[Q3eHJ):SDW0>,H;YNE3YeL@[=AYf)M?2aG(#<1HMFSF2(X:b
+37N&Va-DbT-&Y)Q(R1.e\?,M30.ULf.W[f&-2IBM11GJZ0(0[C_[S)I]3+O/RcT
d#b7&JQQ/AXJCebL&)HR@4:]+3M^&f^JW(eDggbBQ][-K4U]I1YeZUJ(;BHMbQf:
\fT]533]M1X8VLW,R8bA[JJX6]K4c\SZ6=+YUSf<CG_J;;e<AB]J/_43]X=VE(O^
bHS@=([02I=(SE;L?8Wb^R\[)__F@5]1SJ[O9Z_V(_]C=^GS?&B44d&JV:4gdeA1
0NJ.7NGBN6E5&+KA<EKQQ:C0&2W3Z0E:0>JBg-C&YCSe)O<\D<K+bPF]CfR&bT7K
<QM72[H,S+aQR4X\>0e)LDXccO7&OaQ&b212#K:cOc27aZ?OcPY-U(8GB(UO:gNZ
+/10X>6JVKPE&\39,XC4J8<I4)FFFQ6CYPBaN36X;&(U44++U?U9.CB;-@S:-cX:
H;bI9c_&<.;JL[31D\W)5DH1,;H</c_>=P0ZBb<e6N+e3K=LF4bbG^+3EIMYY7>;
25,aXU?^e#>Y:QR,eO>\B(02S.BWGW-&-;ID1D6?@cfZP+2:efT:JX5J(<16T^@d
:91F_[VQLdHe/BJ[+e1-dGBJb9AX>faA#:Y=R^WMAR^a;8NbdSFL6<&,Tac:ZYaG
H;RIM8)ZA7>-L35Ia+,(L2443.2N),5T)Kc,<[]9XSY1S.5ZVULD?aU.,DeeGbYX
b32E-?#0-aPJFDaA3aPA]UASWZA^P3d:L&^3LJ.cX+OVQd^[6P;T@2K4M^B/QDfW
TKY58S^a84eYc[>ANV-2N.,@c,Z1BU)Q+A+O\R8,cI6CI^M\UP/[&XN.,_0\@@//
8X>0F1ad>Z+>D/6^e;NN,6Lf005YDHcP:1\gJ;@NTZ(PY08a2Lf;H9d(,f(?3[XK
fH_1&;N?)B9.;bB27.VQ_g3;RLMXc&:MZ9E-#<Id?aCa_7bZXE:JYP3]<a]a7^FH
[]9(T;?=W=4H^=K1f1V=2,2[GB6KcRDbMf\E[,g0,J>+,S/^6E9Tg/c\9,H)1OPN
XL^.X68g&T7J2&+e<-7ULcH>_-=?B1,6;TZf;_)^T-[ID<4C9VZS[f;.>L.FZ]a)
Sed0#FEXGe,+8WcI3ea>7P>>)^1Z=]PcX1egcYe9UVU<+#b<OQ5WBc>@PA/]U&F;
4H\RB=3U4Da446H0J5d><F:;E-EXPOL9..YLUMgF0T01?E<;1#9d3?N@313YI#E:
_,_M\fFdVDOaF]=4daMG7##0OC@?F/]Tg+GH6V.T3?F\A.>A?f>_?^GbQ>E<5b0+
Q@fP)DaTM-Z<e7B7XAI(NbBIE,HM9@)_CAMHO6/A=#cDXHDS2/&U^1Y>V(1KH6IM
.gOR>Z0([FgM4G1=(,/7MZ<MfVg2&197DB/W<G\]:ZU.,@2_-0DKTUWW&,/TM1&/
K4#H5;>)_=N?56PFZC6O(VK6US;FTAO2W(PNgKaOY.]M97_.#Z<_L.A(]1&a29d6
RZ8<FZc/>R>.HHdM>&d<N@0QV1dT-SLS(YUJ69<V_CIc7]:P=4B=,QU>MGfSLf:^
899gTgKd=7(U-NOe9g7&D4_?V)a_:K&5Ob9IN1fe]Q4Od6K;Y3N(9A[2GdYM.PTe
/YW_]IZXMffO.M@=cFdSE=>eL-LX^EE.=8-MR=X]=f&#bccd=DN79H,O]MaRTJ5Z
(+[c1H#fdgYY&FQQS^3daQ6:H4G+]fF?gBC[Ag6R1g)H36DEQ<U.-73;#eV3PdL2
NT4+[<?bbaB6@O3ef,?c<,^f?J.-M3c:LQbRRDGH0a>gWgQdXFUVR4U=X9TE)<b-
E^AH,^YQd:I6[(&?.(@LW)JXfUHLMZH?POB8I9H1eL9V@0,52./=XMB-fG0Q@R@>
R&R1O;\024RbV#8_A2cF9J2XHbZL3AKS7ITf)+W-,@8XYE1=L&C;,bDX:UIENf<E
^cB3dB8KaB(_:^D0T/C,JJcD_IKS6CP.:f7cTM)P65b^J,=bI>?.-+_+c2UO0&5,
U5gCDWHRT#)7[1SKQf@Mb)Me^7C_Z(96C#;O:eeaOUf[B-Y/):&Sa:R<<a#e[4F0
^@4)1JCa7XRKMB],#GKcR5J]36G&8L1\#/]D3NCEMXJMM/1Qd82#9N7HE1a#bK4K
@a/>GG=7f9(P+[5[K#GX0:Qd>PAeId5,(_Kd[,A#WHg;dADV74F;E6/X;@AW0:]9
,D(>80X0ageF:E^17QKLYETY-7D)2G5&,)T\;J4BW@WHK1PQELOVK?7aJ^/,RcD,
HK.BJ=6)?RN0:g5#7MA\DE/F6IdSRdcZ1(]ZLM;?0f3=b6IKa;0>fESA\OK=3J[8
IWa??B>Q;PH+T5R,fJ,a.>U8=E/)B/?/-6J/Kc+(:C\H7=HF4OL<OfVUe4LZRG(E
H38,8IJA)PXf;/A7UVc#L_3S>2T7Z:(S]Gd&0f,A=K+H:BbYB+TB8fMQ\JWc:4IQ
9PT,U6DG&dCBE7]_IHL>S)&Wf(>72W1-Q>=J][I8>R9#()deDf=.F(V:&V&7WXGb
_55^M,1?>f,)JGdR\<LE0],H)D]>Z5=O5LIEEF\X>,U]D6,(REe,b76a9MWERI)D
@G/gPR<e2[Uc,>+a^;N[VO&MdFF>LHbDIE?bZ0#Jbb#:],;6B=LVMHefFeGUA^0S
&R&D&7Z1<XI8?V(ARA^Q2V7X)+[bOW\_B3[YA?</cg:ZEc)N0;f2KZ=O7Z>L4@L,
1X,[ST3Q9&>_>/JL-4Ag.2W[/I:MNXS(=F=:8H\MB>f:B:ggaK+Z^9VF5,/OY72K
Dg3QP4KYS?LJ0:22bdWeTX&OV23P?aCS];T<cJZ:-K1:XV6DcRQ;/I9OW9UXY<FR
1_ZcJN[><ARF0E?O+4IC&f9)H-<XE:=]/<2@HKJXNQP2+#,9+W8[.Z.S@9B.f31P
Z@@MEK[6Q[;Yc,73a0-]MMA3a8^5,/CW8)017I2S:CBa2\:9^Tg>]8C82;.3a9-9
3P+Ve<O18&Y=PO,c5EO[5+6,IW/@+>VRB/Edc_YT-[0aLQaS>^72cVRGE-a(_7]/
,-Z(f-0#(+&]W5+af>fJIM0@:+F8C+&)9SIRFL#JY\I]T^IX_FPV&IL:Y9B(bQ;Z
P[89^6aVO\7SRX87Z29V=WF?JNB4g-?AI^Y_T]VCT&DfB)IAY+@4=MV(MP1OD:+H
:Aa@I_:g_0;^,>4GM]<)Z>PP>dJg7BMX\08KJ,-;IZcJI,WM0Efgb>YB:0PQC8L/
X8M9NQ_MHI<16+>#IU@I(a>ZIbS3[H)MZ_8(e6B]-\>c7\M/>1KfS@(CcNL(?1>G
Ha0=b/<?+#@];cYU0V4E33#S83c(>AI6M)Y^R0LAJNdTc]0\7I/6TUWg5-^&(I^K
aLcG[2O]AG/]]Sc\LKbMY9R07D]D+@N#KN5KS71TGY4:4^Z0D=;RLRG9Od@I\#F.
=4BVBE5ec<Z@\?WggC2GK8&dQ1S/JZ:N#c?L=X^0Mef7<:,P+\DD?KLbMT<_6UTP
e];YVC9N+M9?H=/]A8R(.3DcDdb8.QfE[ge@^CJ#S0K__.>U#48d0PM6;E33BL+6
(Of]ZC)CG7.M>A8?G0+,RG;G;E,37WVd9>fef^+0O_XWLc(24?9FfZYEJN077BJW
R0-C@93]eZJ-.cX;?04Od((2g-D=4A\C0L3FHe=FSV1GA6eJQ;VOB#DbA_5L0JMc
=:UQMb2P89Ud4]G+?a]7IU=b+L(XF91cZcOUEBYY_-OPNbdQ>I_a.[c\P<M2ffQT
A[3L&N^9??4.J3;(FPGG5:^eOM5(]&;ZJ+E1aP/T+BVdV7\R:&+&>D4>FP@JcCf-
0D6^M[bE^@32@4FJaWX8ccVbHc9NX+=LRS/N#/3f,^T#YXH6aGAI.LCf5Z;M(0Zg
2T;NZ/7c=M\IBORRIJK?P(MT3LXY\)-5S/-,-S:@.J]>Wb;-bSTe^9A>EXe+g>C4
K^dGW0)Y6D.2>Q0TacG5BbG0eRa=/VH+DA;/Y1?g//_9-;]O&S6A_A1?JI0D?]D#
E/g,0-<Q6g^[6aO>NE1.dg],,F9K>B<1O0J_-CS6RWMXP6X+\:0C))M4LLT5DH/4
9/b8_K+CcI]fE:c;]SGJBa_PZB0gac-Tc+fA1c4;TfX]EPX9-^H^LM:M8d[ZQA0X
LDYN)&>0eQP=#^K07K3<8Z_=:d?JQ-SSG<]8J2YL(,EJIU5P-J#_O.e_.N3R,ge#
BaV[,Z46UQGR]]7/3<0KVK1[^Y9B71F64a0_:9_@A4S+&4J(,-Zd^c[9KXD+DSCK
1)ZGC4\(]GBDSHG2/@KYU);G=P(JH\\AZaE]0C)VeM4-KNPU\WV9,8UcBgcE9Kg,
R]Zg+</G-^a71IJHUR)TcgS.7)aQf,.8&COgf607P.]L>@\X+R?39M,\b?d<ZS+b
<[[Y>c/VJ#MBaS>e&Kc(?DJ\HGMfTXGO0Zb3_cQ.=XK0L<@#+Fe=:B/3#D>\IBd,
U1:IIOe[K^(=^MB]6NL52_A^/-Y-T/b2EbYL0MH102SX[(N-?)M9,77Kc4H3;WB.
7aRW]WD:[]7Sb5)Ta#OPf\b)KdPH>,g0R3UWS31#ZWROFK25Rf=)N9.b)XObH4d:
C1c?9Mg<_U3SW.ZTS819NOQ;,gTJJ/IVW6D-0#g0HK.5(GJ@gV:IWVMcb)RS>3cg
E6#<<@f9=.,^2H(PdT+9O0+9QTT1+F,f7I7gQ/,EG1<>-OOCZb/W59Jeb;3N<YEA
FNHd+&)Zd3YR0JQM2d+gV9,(U8>=c3]<=[00B?PKC-ZAeAQJ<AaZP4Q4WPA3A?=Q
N]T2bMHWe:c1?:IS^,]G7W.fa;HJ-AY)@H9I_,]14L<\,.E@eH(bgG#SC0X]6IOV
P;_?7I6f)998gR4Z6H36fJX877:UMaV-RG7D1Ud^Bg^89-RLg=XJ-b;W]+_+W_]<
g__5]]N=UdRKa,#9KC,>A,BVGN<]e,20\-fB5XfM<[J+/+1d&F.e\R=c<^1]cJ]b
bBA^A7][fVSJ0SEQ=FVY1.ZgdYG-,GZTKgDZML(GNS)AOCX04f>--OM2K#Y^P\O;
:0>WQ12(O935X<E5KO1:DbK@,[[=\b@]F0dSSG+GV/f2BFFQR]cc.V<E\V3J]4M=
@V5.(W_V>?T<)MI;#?YY9+&R/aZ?A/T8WPgfSYBPTZAgL,&/IUR40>eGO5bO^_?)
>3?RY9V&]A[7+Ae^.2J/SJ^BPM_I(J81,OU4T.\C8&>?ZKa=L1C(>[U:7FfS93\f
C]3D;2K\d5[28D_M]_AZ-D=Ga\F[R4Ug^@FCaVHB6^A,&_\]aMfQ7])?FQ9SBVQZ
/VGTZC&bW0K2F]:L8-\_7I93Z8-;]]@D;$
`endprotected


//vcs_lic_vip_protect
  `protected
5PM>&#Ec^Y/(E=3LBFD:L71a-].7ERSG()cD6S87C\+JQ5067&22-(aPd6>-]HM5
gTM/J60\_S7.X]R\_H>aM]+SLYa:]dU:[VW[P37FaXMCL0\U]Ze&e6@RVeHb2:68
@X)@UJDIgd50W<ZEN7-GVI&4_3CILA\SV&[&D@VB1LGA22MK2@^Mg8dN)..-N:Q&
NbU&JN>&>cPZ1[=C@-Y-..Og#f0_48X\8U@a_F\d#fa]?K)Cb@7@B_R1I<OL7/6Q
WQJAXcR:X1/+Q]I&(Jg__UfT#S(]5:^3(&aJJA4+AGe6Y#PBI]LHG/Dg2[<=U?>F
=EEedK[LZ<D_VQ7R\/Y1Z3>@^>+^=@4F9#INQ[W@]G8(/Y6-A66ESO<^MQIF78@I
D4Tg<XcaJGWR[KPPN5BAQ9SIg>9H&F)#99.Cb7XMbgT5,F\;SS8:af<M[JF0>Wg2
)M#0.@NML_73/HH:aE3C0T27W7.?L:3HQ)XYG4O^Y+,[X>BQI=#Raa&;U;H4bIQ:
-O90R,7N:DY:EdM#U6B:J1_]ebR2;78/NKTQ9^)QP&,gG=<VK&._#D>K<WYMN^6M
#?A#/:I>60L3GJ[^@>_@3JKRPR.//XdS:ab?H55ND:8cd_(d#)5RL\/XI(?N0@8U
8.&/CS8@gcdJfeV312^:b#P]4Fc2?OXEA&<5MDJ16NNWZgNcU;aS5A+7)7,:aaF+
UUf[6d)d_.[6>;-=/Q7A5[=g.5Oga^D+LC\,BJR+TB9J42K.GQ4KG6,AJ9C#8]J:
gN,)D>=^ZgWFK;<+:9U(_JQN.Hg-\>b4DV=+P[U##f\4]1\\^d8LZ]KaZ6/>,?X(
DX9XC[DJ6JY:b5;-Z7^P=5cNa&;3HU7Ab.R&N1ee^ZAfK=UfG<P+-RF@O^R\+F5S
94&#P]<;c>,2H-g3Pf;bbDZG8RIaI>J2FBaLH-JUO<^)HA#e(]3+)5]50@LG+f0P
EaA\?MGFI&WDPc6H5MTYED8cF4Ub6cM09]HE?6J6YT9cGU_ZHcFY688>U8=ML+:6
@fEbF31c.Pb(\_6e.AW7IT#]X&U@[X-+H?WVK[L\G2IC3??]8dSUaD;62M1T+;JS
93ZK=,;=>dD8<:d9.UJ>TXL-75GKVa]4KPR\Z9XMec@DW9_\JC];H>PN0OO+WQWF
BG#,:O/J21Q-NX,_[OB>E2C+Sg3ES?>ZKgeN->,\Xc83bc.=L9XY5\SF38A\=BJ/
BQQG0L2fZ+b#]b^\EBfWU>25,KK_GL/;BdZ8bggWQEXI^+8DW4([BSY8:UWX)aeg
YJ.J,G-)g67XWM:_P-M<^O2]N/=:PV7\M-R1F4;H[c5NEbC=HQ\ZURUZN>J>LXK.
O5T22e6f;&NAXBTE06_@&RS/95+;gIZPS_cGZB<LD/Y@)<0\g(eI<gMc@>785>LS
ZgKb(KCT66V+c>8RZ9OP2)8)cK@8N;ANTgHe+2Ka8JA;/ZB#agG\U,_YT2^B7D+a
[b\PVZY0EcOWdX>8QI,@;<IcE56SEYKB]E/>Y,3@39JMc0KNO=eT4/)\DT?]2Y<(
F2+GcY[P#V?_/d<-LN.3bTa-9DF431S3eb,dEN=(8RY=9L(PZ)T6T[2[.;-_TAI2
,CNJ3.L(,fDV^4Q;]AfMRQMB?UO#6A1^bKgX8IWbade\dK:b7K\<8U=^fb&=fY8B
Z3MT>eAWdb)2,&SNWZ?2RaFZ4H4PP;[bN<<&#+E&K\SX1X(D.:0Mc3(T8^W]0B]T
b6GW<\-aAN9aI=-T0Y-YOR8K/>>1554GL3:&?\+PdWEMdP(>0T[B[.gS0:,Z_[X1
&b,3C^&FU>38bY(F:g&ceB4YgN6.0C[eg+Be#WEG-Mg(]2Nb/gB+g(P1:8ABGcF@
?ZBIO6PQ;QKW<(c:4>a3SN_L7FH2#GeA(UX5(@UTDSN;7gHY\WS(OM[5cNDKV374
R@\=FA0fK1f>P&1AcI[0^IFD7>(T;b8OOSZVf^VgX&:7I<V7SR;5[gU(9VJ^cU]B
GI4^5IKO/IPUb40-]F:HGLa41-B7Y5c]H#cD#_)bOeX&8+H?Id:9LJ[V8<f](Y;&
M1GT&A17COS?F&1-8_I\>S@X)K#&:#dUQ<cN;HK:5_?<X]eU>399+:ABNF<,0#ab
<Zb:\f&@ac+2_1\CY4c?+RV<3ET(O93[P?M]0E#Xc3V&aFCSe=+<:Ng>,&H&NMOE
EBF,26-F&]UUWL=7/BD3/(#4-d?[<#H;L\4NI/R=Sb-S>YZ72<V#<ISbS9WOO1Q4
C.S0[@,0+0FPc+GG7O(^,?W-:V=2?](123P);Z91MSQSU,c8FBZ8#P#RafFNYQ(-
VcO5<OXCR^6UdFgWWY8Z(@WKD(B_eCYFC7SOK;4UB2M_Y7BfA@7M4Vb5gY(/H#5d
cY1XWR\^8N6)-X#8T]]Q<ATB5(1XZdM&SO/X<L>9@2+&0WZ&6>-,6(^cL]8DBH3&
8_WeHf<=V^+IDQH5?-=SdI4;/bI=LM&]WH3RHI-?-&f)ORPWLGGD4]KWB>7#/]\@
A^D84]S?:GEL2^F\SfTR->/MMDI@DA(a>\WIRF?BYMZY2fKdcdPNb=e<G;P6-^[c
P\M_YR@[g?H_+7NQaG-e(FDO##JL3J]P-L4IQQCGW[g[M?<<EI9(<F-3aZ&ee7Uc
WKY0bL59#+D7#2@PUF]g3VU.aR93TIg_\NL\Y(.9X1A^9DSJ#?^e8X>U#+;E6bUA
XQ6e7N[Z-Ib3PB=MHZ)aV_+e&_Wg^T]Y:JA-Va]H6Y)4XX2MeXC@7b8=cI7?&d4d
[YHZD-0gfc7F=_C4cZD4dI5bH;J04+^V6]EcOO/J1KESb+LcH>GO:D(L2RdZ+EJD
O2+OZ)Z/;O\?6^=NGH-b@\A=Ig/CI2.ER7ISU:O.RI7e9?293T4M\WKJe:B25;.+
/&5Ca?[[WIN<2cX>6)YNHfSA+1YI=PY^MbM><^A8QT[e^I;P46M09\L8O@N?3&CK
@7UZ5O0GWbK1R5TS+4A^g+MF@&\+\\)M@Z2^]Ze2T<ZfV\H4YS[AV\25K3&afD/C
FD-(VP@(XME-L#G]TN#L&3X5?<,(][+^Jf@NU<BQQ015F9?&b-Q/:UA\dXb)6gUE
aCYA8;+c<cTR]R8eBMOW>0]T)^O?J?/0A^[F9ID0FOPW921f.=#aBSJS2f>a81K0
V\fU<W6M.@a8aaQD9[(<SS-L).e(KNAG6/2VK,IfDR-=LIK<08Z3,>0GU=eL6BWD
:W:\I?DF;,aXAE=BP#bcRR(YZJ&-QO^^QI:+C6;WK&,(=O83#KYa@3,Z88[T65;L
c,G[,<Hf;2CE_f7[.>N_7J@Ie8[Zd\YcLbUD][FVB<DH4EEC1=K\_b>8fdg)fL@W
B<=c6^M?:+T\U4Ua?:S]>36E+g73:M=B8^8KT&Ceg=H:ZRP,Xe2Z(CY)+0D\E9Z3
CB/@1c^>^Y^WEI@BDV<K(NAD<QXN#C#Z,:7&G:_28a&Z-Z,@@^^a</LQZ=Q(9NZB
_[4_&GEB8eK4<+]U^N2YPQ=K_2HM.],X80[_AALB)a0V&cHe6af?@WK@<-3R=-R1
9]7d,L?a:@H:ZX+=HWc(DP&_BdTXH4-bE#3Q+.[\)RIW&LSN8AQ7f-g9afQ>[B-@
OgGRZ\;Af;J6Sdf8J3Qa&);<?(+,);@b]X9e8/?.K1(U4ENBC(RXW[&_+T0cTJYR
f1cE,VPZ0QGQ\(@W^SY,dD.c(J1:S+-WQd]WKE-UGU8O>JRMe\YVFN].<ZC[R1Z;
=)<BWdIe7<9;b>b/(IOXfFS/&K)O]d&bbc>;AG;J69UfF9-+@X07SO;7QJ(W_(-B
,bRI6dF;dPS8M#&?TgHPHE9+&\,>T\XG#HT<=Y<WS8-CX@<&)\geA:e00>LCf(C+
/97H=gX/,31;&+(G_K/5L/G#9?^bWM_9?Z-1/(PSK5\&c\M4B1GN?3fC?3A.<&1/
gD(([b59:XN>,0R-C1),O7;bZXf)3GR1\2O_8gGL9Q5Kc]88a3G8aFM9YQ/ZPbVS
4/FZLVO^:]]3Y=JbAM<eO>B,,F^cYG2dJUF>Z@bQ:]MAb@AXHT3AGHb)^KMDL?#c
RYeMe&Q>Ib,#+MJ.cW@6OL_:^E=0LA5]];W^4#>VQ6H6A(-[^8Ld?GQA.&bLC#>L
.aG2-^.b.:R;:8B@QXC-,<14.aTD[^4]\K:78g]8>&W1#f^ZL)G;E\UK:5.?]c5M
4ZI5C^=TSFd\XOfW50824@Hg\Z-<.X1[[\dOL#N0?bZ6XMWES,DS:XS_L5OX96SH
E\YS2OPO_[FKT_\PC(g+<496NJ5WB[4,IEVKFX^b>gP[.H00BC,H;TagT+C5LVVS
g3I[>TF/8eE\S.K3SeD@#:TJA5YZ&1MO-(:IBXY^\5;O;TcVJ2e[_#g<2_^FL[CG
1W9ea,e4L[4MJ23#3N]AHT51:N_ZT6-WZMQ_)g/2KaWTd>>R]/dcSLK)W(^eDS:E
,N#BXdL?0?(>bgK18b]f#\BE2(>eH4;3]?)Z3E2?Lb@WO)W#-g,J-bA7d<MO8A@#
_IH9ZX3Cfc)Rg6V;+O3c4PJ>U>/IQJMf/(Ue7-cG:fU-B_e.[T\;+A]K?aRELY8g
DW\IHF\((@_4eP)857fAN>>][8]]A_&#=_1J:2)b<82DcL93b=<DCHP(dDT:9FWE
CI:SNa?E6)IeQ^-16gD>[@S29?@[QKO#gY#TBV1;8gRFbNGY+eO[0\73TT@)LUHR
>ce,G-/1:d@-208+C17)HfBb<[f/2[HH_#2?35XX2U1?/4J#fT52PfT?.^?WZW&D
W_]a=LC-2?G:I6O9:V-f:VTO?NP(.K1Q+BaXL),4L:]@\79eQ22HT3ISdPG[e7T)
^9S@2gW#GA0R#P5@/[9\S##_9P84FX]OJE;6OI8Q3B+=B:X-O,K@eCXP[@<[c7-R
NHc)39S\,C3+)f:13gXK^V=Z2IDBEdTfT09WYW,38VO./>6ecdN,a8-#a-.^-9PC
QT\L0GL(-K7@4/1B+,M4&GdV&Q>F\Z>Id:J?M_G>gfg,C@/==QNQTU_:S<^-DT7P
=K[&Z9X[GWY@5-.^c;+HWG^eV92L5,\\(JN@#?MWOgGa1K;+BOS4V9fQDgL-LRP8
9L&gEdCSI9O[#86dF(R+CKeFKK7G290S.S9BFV,-A[M8JVS/=#U+ZE7SOX@d7fEQ
\gf+1IA\\,?,:VEUQ:Y&gR)BI,_7>LUM7#PY(IN?1R8Y[9CWPLSNS)OI#e1P&OD=
L724C5Q7g9CNNA?=1GW7=YGb3)U):9EHP+<_T<N3RL:OJO0463+BZ#NO5UZ@#/8E
;:C<\HHQ7,&E8BCNQ2\V/P[Oa[>#_8@G7QN^>2O^IcN;A-+(=UB-G9]K+[]Ea.2^
GfK#CcK=H7d&9B]@5V-1\2S0eOTe6O28N)Wbg&ff).c=Hd)AYF8gHcSe]<G9_#)7
M65G/d)I5(IUB[6I/EK9Q0ZQ;7G2Lab_MfTMg6[=&e@Qg>#2QbG1SGJd9,Me)&AS
8T8b7N;7-04Z7+d@E29X<7L7/)<<5NM\H@9e/?S:O^N;=Pb5I_J<,E.:V:S@5[O(
5.DODH,PK06KR+J)d-(3AG0[Z)UeH(YdbMUaDV7[T^Z1VTd48>0MbOPK-;[F1G0@
WaMQ12FH)0U1X54&Q8b48(Q^3CHSBf85>W+B\A</JB2-UUI1?DX/=]4O&A9PY7>9
WYO_4c5TQO[eUHcOcGR\)V2GP;XIDTa-IB;RV\ON0a>P+AdT,[^b(Ja9LBS8.[I,
bC]J;c\W,\KK4(_9MBLFMN)WYVT^,=gFNV<3F]_//?WcO@H@=/YEQA-f5=1YW]ZI
gP2L-.Ae#\&?R5>TZ>3?MT@e/[I9bXQ:#/1W=4Z+FT@<1Fdg:A?_f.c?S:Q_1e/^
OE5;5SB&)]>.5]#Q)SK.NU_:CeDbd;BKcFQa9YM_N2-6.Obd04:2:X0B?J,0BLH#
^-MHGD<dWV&:M8@&;Lc5gS]EZSDX^c,8&6T]WFSJO3_Y])8H/A<BM-=-c=dN(/aG
g0TQ#2AWf4KB2dF&/efK,N4N;M##\XC?HS7VW??7.D1I<&[@&1?VX6-+225O7dHH
?H3d6.:6EXV[B;cD_N;F^LC(YHHZ9SED;C/e#[&acS\b/+(bGH(e62BK@OTR_9Jf
Ta(9+WDO>54e;dYbTJI/(cO\NgO9N<7,B_LIG?I;d?/<[4Q0+66UE#Y]ZKAVaVYg
<;\6bN[+?P<@&F=BT]V?0C#.DRD+390MB#VGAN).1YVb7F6Rd0),,C:0f,40S&BO
XS(F4H=+=>#0&;g<4016[?=AY_L;4;Z+a@JT6]QB\UM;?&RcMC]W\:_]#]Ld4fbH
eIVfGY:7=aK#+P5<TbI7#@N9gWV=(JTRJ?XEa&U[0PT+adeE87De)8@-]#a&IZd/
;,KG5#&9;ZK([F95,45d-^1OgTR>H2g0e^16Mc:Ic#:aRV/_E2B5@4?b+7I7;>4e
33LNeE.\WQW.VFEOfC(2DBK]d_-a/QR\_^7MOR2N93/P(;0&#A#=FSS2Y\[)QYcB
\]bV^YJ9c-)[H1,[0d@I9aMeZZ=35abP<F;^S3)CLKVLLTce_WIVORD,O^CVXad3
XHT<A>9#@T;[PbY5M2BQc(-C@3IP1Z4K=E[ecA\c;TCT\9>4-&;@L;J9WR8)(V>F
+&_4PA?\ec=>Oc.,]N;@=)\)=#,@(G&QH,f041cYIK>d=D(#]7<FRbNAf;U0^eP\
/=+EC&10ScHW9e>\(W.<&CQZQ1#3&:/X9^TMKc;ZP&YJ@&G)9C(EK-DDe:,66RCF
eIgaCa_WK0]F\O+Gc30&,(SH^C2))FYL4ZgH[O;@43BJ,1bW&B1RaTT6f8gH52U,
5b0@?32L2gFWg=b0=Od:_8Fe0+H/@Cc:AF7[A]caL3?GDH3R)5C,D^3.\@(2X>IU
7=F[PV/)=NgP9-?KU_fEfL@VEee?g93J<JKa+U;26D2PB5?9FJ@BY,VLN=&,D0L-
6TQ2UUZ#c&S;X[EY(W.];X:BbaW2WQT.IJe+PcWT8H+M_WHDeA376.>D/JPQEGDF
H&YXagUPSbVP>+GJ+ZOKR4UPJ3#89/=]]K3XO#c_7ZGJC7Z+ZYSQ1HSFE+[L2XE,
e(LV8Na82L\3Jf+<VY@JH1a:8?FR8NW:Q-;K(>d0XE(b/\IR_9HeZ\28d14NFPVa
ZO4c;E5:HcgXE_5X-B-C_:BKK\Y6&OA\#C@e0#=]0ULHU3K=;W1=C>c=\H4b.?c@
4Mc6ge36MS=4SB\^K?gU6)bZ(=5ZM(T-XH=EQ/?P4=?_;ad\5+S[DKf39/ZR,-@2
Y.5\XOU##YI^GAC..g85>7UaIaUUM@b9[NYdOeL>W\^M2+8/M/]7DDb@Db^B=b4.
@L3\Y3#.+&.2]]g8L4C2#3+K\RI^[##QI6P19Bd1;\K-3FQLW1fWQ#K0=7G4JN8S
C^Md7YY0(>T>B_8DTMONa0PSJHCg=+#4_?3.3:L>/#5WdV/<fbJ&O)+M+Q3+>b6a
7XK]52(UJ4]a_5Q:)K>e,AgAJ6;BP]./--:B/7g)]<#)<N#=.?GJb7@HKN8WgABO
?A)Y1-X\@-\1Me?WA1709[0#>7f3a5.P<ENaH_H/;bW/M1E,)Y=M[VJ2W6I5)VH2
\.=QMfN\\-XQTG9egOP-UKX)fXE2POReNPQPT_OP->S\E1gWK;,J0F.G3[HWO+V/
,I-[d7Eg<XDc1-Ea(C?Y6<&eTIE0-HCNJ11bJ[c@:\4d7QFGT+1>>\9L4(Ua@RVL
;028R5Z)29).V>^(BW1\E-:ZL9==fE#D_QM&?G(HEL(@T;5IdL(d=6PC<g>H(?SW
-_H-M6[QGL\0X9ZeR]^5a)/^2c:\_71YeV?)L27?a6M82]M\-a2<f1>bc=C#:(X\
UX1@WX(ML6B:HZNRa:08^0dg7Vc7c8U3dWGYU-=5[DO)fHV<,Q)cE<F1YN^\75_a
fW/#6Z0XF1b/WKgg28[7)I,9\d-A40P=9/9KF\IQ_1.bKE(2YcWWbODBX.L,gTbR
Ne2gYYW33DM7<C:(I@0P@&_0K79(:X5[B@03H+,CSD71>)[+Q40GB^fG_:aZf3)W
\JT<XWdM7#GLEfgef3G/)_a+eCOT?9K/abC]^702;D1XO(FBa6U6b)?FCC(R1<7E
8KgE\3gOK#aG\B3AIF;MX4g6e[TI,;^7)??<I_\/TE^S6)V1/VP:YN=<=.>81E>_
/J-23cF[:9=>#E&T-4J[E:g#Ec.P0_O_4.HE:TL2,9<^T<@K:+#O84/ddc6.d_8D
QAJ1f;=JP,;8b:NJK8ZR.OI#)R(JWg:+D<D&.dGKF,;XS5ZG4],DHDQ/AQS[g77M
)7R?F1/@E6f9F]DM(Kd_b^YZU&aA/+F<T2@XUSC26(+;3R;JeFRH,IGf\.g3++03
c=6cP(J<YYc>]&BJ8CP+V+&818&_UQE#/\8C.dMCa_gY=JbY3-(3:(X5[NEUgf6K
.YD0O99[5F7PVKKUE]T\V9N\/GY&YXc076&aHKO?(E.@4IJ?_c#+)K[&,Kd-BUBC
-#OPad11bgO4:e7LVe\6LN&-1])7N\U3XOH>/aTT761&2;aSVXWg8[?&;O>,TQG<
W\fGWbR.0E^C:N@,1W>f(,:NcJ_2K@B3V\;):C?;)W7-69[4NQB(8I_+.O3K<(40
=<M(U+1:LEeA=H+ZI/U]b61gOF1GNU(d6]b:5PKX3#-dABJg92;;RZ5O5(JNEU3X
N36=We3+9X]f[R?6N7T_ZR6(,RKNK>Za^ES+6,7>O5@V&AG4X57ePA[H^P?TdI-a
J61eE4Y?&7SJB(#O3:<+D2W4Na7+fLX=]XfDNQ_b&#M4[RMG,QQFO(;N2[ZHPO&O
5Z+N6>#:EJDdf9<>&0G?Qb7O77#:7^:F]e9E[_>c4.gW:<e[_@7#]AA7LM4>0/Eg
H#[ER:LL08P2]VK)F&XJDOeg0Gf#@_Qc9X4C7P.JZ.VAe8:fG>CCUb,NZbJ-Q9I2
KU@Q@Eg++a481H?5-6-7UB4d.0FU#Z)((Y@K72)/Ee+/6ecP=^,8-8BgEe?-eN?K
M]S]E_bA,/VCEEI3#K-O(FH_KMXROA/DQD0)<P5a<>@J/1Hd6XdZ7CgI_(O8g8Da
Sb9)Z^T#Z=H)g:QCcSQ58eFP2&@-+3T[X9ROJCHf8&7L0KANRWd\_+:J_5_[7;-<
:F3:@eK;8OI=P@;X?@?MfOTV3a[d#G\)_SUQEEXFO&H3c&DD?AK?:>LdSTQWT>Q.
D4=15^a=(P8GP_^d#W_80J=3C/R2ZQd#OFaI\Q\1:4<ZE-=?b5(OC=c&?556EP0]
<S_DNSaABVJIdF9HaZ@S^a3;Rff#UMB[&+IQ5e.6_WW)2]Na\^@L;.,ND/B02aSX
#[E+Me?J_&gWf=#HH&gcCI1a+PHNe+AVS7?]4\e&fDIfaK7MN]U9AV,g<N91]]QL
QXIN6dKEP9a\X<L7&+P0\J\JDMN).OY<4]MU?Caa]Y(3@9EPX;CL@._<1?N/PA>8
OaXKcVM&.Ld8VD;K=Z?Q?Rdd>4M:2.M^[<b2g3HgObeNgf^;R,/TITWBPW#+5VDf
4Dd>]]ae<ADBVeV<EQ]S=XEJC/HG,TgP@:3G[S8Reb8a#fVBdBabG?WTJXC+8^N+
-3_HPFAB&X-8</Y/eWE1<[(aQg@J8P/PMaN\###.QUJ>^F088-7OVJ?UY&X@AT1V
,BK]X</8,5LU^]1F@XFMCJSgK0(MFe3OKBRHVM&4PW4QLGH_R[aS)E7_XA5M]770
9]G4/^4D<VQb8Ca3b&?F-e-3/0C,ERM3ab)g=6G890.F[0BP^O5#^LP7SJHDAQ@J
<48,([P=c=V5E/Y+9b>)DF21PQeJU=T<?@]P_\3:_\_YAe7;.@^)bNVJ?gT_(c,2
+4C<E4(J#/IdO-]EB4VYNaa1,_XaJ##.eGf>>W4LUX^+8?C>8aLTDf0_;_F4Q;c8
F,@\#[QE;>e(@T6_cTJ&QQW#IU,dEFZ1]QH[YB7[^NJX15OdAcJ2_-T,:aQD],D)
BQQEdQ1V@?-@:>D0G11Z9Q<+gK63+Ygb3<01#d-SCC]R1Ie.S&GeSEJ.C[U7bb5X
_be]<eIf1>[HB5VDCBff-ROG:G57a3V<WVOd>]F_#<bAVH/:Q+D5N01<<XY=\_D&
76cQI^#J3.VR:?3T;D-0)L&>K_aB(>01YS.4,dQQD@=OX;D@VDK:DO@cYSP6/Uf?
.GeL[3@?f<>;]IK+=X5G58TV[&JadBY,7^O@a_2NVR)#2Y&?[6/VKBU:7.[J6DQQ
\K&#8b(HN(90Kg8N;[THL-6<ZfXQ\(UFH3<(d1PTW&MaFG,7JM<URWKGG-G[;;Zf
X<Q_MH35_CJM1g+84MSZc?VOHN_K\]cB7f<XCbO<+PRZT=c=b/:e5CXa9Abf9R?>
X3>X]-dTfcUPI?cOH9C&()]@2-1OBI7C#5R0<A.cM#beS.<BG2ELB@NNgdg)((^GS$
`endprotected


`endif // GUARD_SVT_APB_CHECKER_SV
