
`ifndef GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
`define GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

//vcs_lic_vip_protect
  `protected
0PXE&8-6\2//3EO,TT5WN\BJEDQfa197/YGdPDSVH#g&##6<4Ca\)(S_gW>+JE2E
Y.b6S=7E9X-0/:&GEH5,\X)3>6/#Z;=Z)V@6&IfL^(T(_:gf<S(4@B?b02FSUgTI
TJ,B1.GI+)-AdH1UD,.)d<[0Q^HC##a-TBEaR=]cFCY>@>#W5\A.e#@,-E6JbG+J
),LdG+V_dUf1XZ6e1UQ(MQ#3=#O/BI?,OS53WLUJcd?C@>f7bIcX4B1J\Q/:IK&N
NX4C->>,eF[CK:[JHT-LJ1>&JPM2(0Z)-C5=E3(.@=PC^JQ)E-8\_bZ9)Z6S[6C_
HMI0MXf^D(AWK(^^=:0M(g@#(P&a)B]C#G#9aO0AX+@bc@FTbDTG8e=_Y4G(8LLb
QQVB<U9eKR6@J@;U?X-ANX3Y448P.PeCA0=XNcFXaI=g;Z4R#)aYX>O(JH9QI#4F
cF>^/ZN]#T)?9cIPO86GCV:V1OPYc:U3<aA@2BT17dN:&=<+eP(G2T.M9PKEC/:-
R4Q#-&P2=0;01H;R)_+;8@GK6[Z-[PC9M((E)H<3L]Q4&MP^e3730QAedHa>ea4P
<d733)65OebJ(e].GOV21(AYYU97DX0)<8H6gW1I7-/[?=6.75>;IM(@_#LFO3E,
=H9SY>aE/g3O6H[6D-:&SKO=a.HXc:a=612/.JbT&OT^CP?/HPB72WIP<aCcPSU&
9UO:MB1A_A4aM-bM9-[U8B96JKO?-2=AJ94NbJ3]fRH9L^SCUCKeANg.A^0c6/>(
]GPg?0OaAGC2K\&+^&g,-V:=XdDQ/OMX6;;ISO1W7GeC1YS\gT]3De[8J0[7SV0A
Gff3SN<fBgGZ#O>Z2RZI2[J/(S3_FGPOBHJPD\^6W,gE+AJ8S;8]X2U(CXRA0b?Y
a&&4=0d/edLa-ZJ06D/<;?FG:9W:3]C&RZV?E-)@(13aa<AG#=2)ef#:@a10082/
K59-#IBJ4@KZ[&:GGa;X6(E>OH;L:QQ]P<Ra:Re30OIA8<MZ+3Vg1X]JA?)W5_49
V]gTBGGA12bCWP1O0/N;Z;&:S,98NP.Q-E:B1EFb.D/E&2fgS6@#=0_]TA2\a);_
35,(2<14gg8A4\\OTA0bBABC68OPGc@JO8[4\L8[DYaR#T>^^JE>#4,=;cNLSVIS
fW;NBLg<]#WZa<d9<;P@Q>1T)Pab8X,LJY4:[b0H0A14@5ZMB@HbJcd,HB<@MKJ_
2>dI=a29,,@XY0C1[TF6MgEc)TLU+WQ^G1[7,Y+[bOJ1ES/;C:904R=O]]5LD06e
<W(GdJYD[;YY@g.Q/d<-66[Ha+/R>@@=TV]\eK2F&=^X6/28)X5-MNBJ#RJV\-N[
356A9\C1EgXd>IL6>ABEJ9PY(R++GWI,12LW-@JJCLGRA_gA<ET?TV8_C6HA[bOU
:40.^S69c,]/4JZ@&0W\S]MM<LES:?8?1aYW<+1JT@,&PKWN@b&^I@Z[#4-1Z8Dd
?]^Y>[Z-?:-7+KJGbdNCB.aBQD#;JY[MceTc)0-2cZ[I3N.>O1,I=-g/DC_M/@R-
IWba:,<NBB)<^7Z22-N9^#0MDMcS+P1eO9:8TYO6(JYWO#[-?c1;PcUg4-5?42O=
]U;d+KcWI86_?)V77VF3?b-]9]/.1BcRe9YSfSP83Qd)J8OUaGE.=(IO9F,3H-E;
[:5[X[BHd_SG8F@P_UeIa&U2]<+YGS<EBLHHU,)V8[5@dFXLA?7(>A>)8X2<d#,>
&6J-Haa0D<LI,bg[P5bO>42?)AHW,;9O4OG/G,[]MA,N8,Wf8:.PG8,_WT[/6I6a
EH1JDE&U&ae#>)C<7&&4?MFfCXJ_6G^J)]5e[5@d8-a-V,C<A<PQeQBD8dOC./AF
G[Tg86K1T3GD\PcFSFJ8fOM&XP;IQ8AK\(>L>?PY/<H@BZg]4R3E#MJS;L+&C7]V
60X?5OYCW_HJ4Pca,I&/]YN=6UTZb^[U]PcCXDX_7M9E)@M8#K&^=8.)=N2K?WVW
&OB^XNMe>UAZJ@CILJbB?D@^^>+Z<c)_9,FVab)b<EYQCddL3>:[.2LC<9Q16fR]
EE@P1)+FXdR8cbCL^Yc8[7+\V7<?<&SR4[;1=E>^JSLKdLDOOZeA;e[K^4cdB43L
M,fPb9/UdJJf7UaGaNEF>Z5#OR7=>36?TBT]HXM)I<Z5[:)/@Z13]Zf&46WT6RXM
.2Z,S=+PMSGK;f3TQ\G)\A1J;(.1I>dF1:\3FK)OU.AdIM)49)-193PUR;S/?1>L
59T^,[gPZ\J9]/RbGK1@BbDMeYDE/L#3RYWI[d9MHc:CGaCR/Z<Da,\?N5[7ZILY
V\L)U.<SQ.A\G-DgYST@&_#D_A(G(T66HPWX18@3^YWU&V]P(bBWFU#>JWM8L+b(
5D,L/RK.(M<SXd_gB6;WPI2M?GZb)G9b<.T#L_RKf=4]a@I^;YdT8L->HH&eAgf:
#>?eE?N\ZPKd24H:7Gd<IWO3OaZV=A#EL6:]7UO:-WGKW2Y13LW>Q_3#Ea@)-.S@
6+(UTYI+1?RX>W2AA[_X#H8Z\fP#JY+&Z5<Y]/0][]\cSQNX5,L#Y(U,RJ)W(aa7
PQWY-+2AOg:O+8^.cR(,8+5XCFW;+>:;<0N_]&Fc\/,+\POCWMM,^D:bY#1HEI0S
@NcFEOUQE:I<>ZL-H,GV[IV=V@D0A+R)]BcBgE&,bQNe;T=]c\1CJf[)2@>Ld2U?
K-_RG(UHbUd=J2T/1Va662R;89EQc<>KGS6ZL6QB>&fKSadc=^dSF:/(>fFE.>E2
(L2>+FgP^^(]EFKOC63MaEHdV?)M18BS+&@VRcKb?QKdYDg-[4@Q9,QJW)2/K))D
W2e=b<V;Nc=Y.6CU;IcXHfLV[CKFabfG8EM/Zb9VV2S/dXL?(T2E,O==QVHIF:4A
OYF0.UL#A4_X?Dc8IH\0K?TdcIT#&bIZ_c#e0\g+7G(He0?I;,T5O)J9]f0UUPRB
26T(^4Z&K[LS\(.))AWJYJ6=D?2I[#KD\]J7GOd.6-&M7K(CLT<5H[?6T@:Kf/Q@
YIg?c([gON(e92Z&Ua+2Y_5A.Y\P+f(:J+c.VRIB-,DFE\5MUO:Y/=7F+RS;,c5P
/36eR_WgOME:32JK^&MX-cP4dT[d(AZZ<ZU@;X-EdLSQUNO0>TA<]1P;GBF619M?
Q\3UgN,2[+;@Qg96&8\J=^\f364ZA7:BWAc1BZX8gTYX&g=M(bEbT+0M3.PFd(-;
1O:ZKJI5Y<^=Sf(b5efC6&GFF-CcYSA;LQS9=NF;_Dd<4+?^bJ<eT-?YcT(@G[I&
Id+/:&;:e,_-5SS4E7P@R773@SQ\HdRW51(MdZ98-2O,8U&/3Rg4#B-XN0&S+-N8
+e--3/TdR+X#ANPQGf>CKMS=EG5W;<8([V]3=MA;900?5/_L/EC3:SI>V^NXFVYN
Z@Sa+<80S>SE(LSJ0F7DY<N:71W/H@[TY=aHc&GY6&fb52f)Ie(&6H(ZJ/KXD;@1
bM-)E55?fDCG=YWM:d-RD965SS;gT7PQ(GZ2HAa873@SX3]&Ug+;H#VgX57N]W@@
/)Df9B5I06a03f6^M55_6<]RgaSP,MO#GFQFZ#G5EW<KMYZ3IT]P42_9d:^PSNdb
Z.4EC#./b14:eN1LdW3\5/SaF2=6)5<GCS]._C&BW_G=V_\5&+:)[?:JKMSXB:NI
Z_gRf\E[4_-A>+f+_@B#I?3?4fPN6,CCa6;>,0(J(82AfKacb8(Ze,&)\4V(#U0=
0W?Og6MD0Sf&TCROH^^^-.dg)KG,]_Gabc3<]e6@1MFJRW&WIAQB^1Q-A)1(W\J-
J6Y=/865gHR(P0@79gTANd4).3OU#O7Q:<90JJBS-fIBPDJgf4bR?<-_WS4FN)Wb
LR_[\:(QS/T)C@-[41-:)5C4(TMZK)eJ;(Ma17;YDJRN[Z6FGL#Ca3QURH>PPSZd
VB@TQS9,2&N;;>HXe-X_;^6P].H#Pfg=1K0fbD?WRJFNA3H>KGcB?O6+,:bbf7MW
?750/?BeGaQVL,KN]QCQ<DRP=V35704G;AT34)AWMGVL_Ne4WE)G;,7?/7T0c_7)
UA/D<O@+cf^M[aLQ,SSSSHX3U<e[9EUD+1]\Le.B.6aQ&5HZSDTOB8QZE2E>\+?=
REgZ84F,CN.@7?3J^]cCZgQ=D#I2X_U/d1BTa>&G&cg0-L+[dL?S2,0bVZP]K0ca
7O5gSFIF8KY]2-]4eWZDe3X1?gcUfSL3]EB(A=OJ,AQ]baef2^](A]&.<QNcgL9/
b9<B6d4P7K,bTJM&E3<fO816OJeaa-+91+Pa@7CJ()gg=]90M]06?GK[A8H,(C65
V<)SecE2AM30MK0@g\04Z&F9a,O]fc:#Q981g)M\R7B8O[@3>YEgbL<@_L2J9NT]
46g;\1^g?#LHS/c-P_K)dTSZI8QO(fMTTc1[T[UH#P^[X(9+X8]Z6G@^K0+^(TEE
BVK;#D22K^\V/VHLZ,T8W3VAT0MGaQ041OgS/W8Rf3+YFEI=@Dbb\9N)PM37OS_g
2FB5FNEU]+M<X5D,BH5)Ab^=VfH5L+Z]_;6B]551KXAQH(gC7ffY=HK+AZeKG)aO
H&c]8#)fCWI<fFA#\[5bA,G2S]A<dW1^-V2MT]E(YJTHYOH/M+QPKa7<e9XZY70<
RWZAG(D7^[U-YINW7(<GJW#BS7T>V>[_?+/>0-20;Y=;Zd3^@U-/SA56_YG=QS9XR$
`endprotected

typedef class svt_ahb_system_checker;
typedef class svt_ahb_system_monitor;
`ifndef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_system_env;
`else
typedef class svt_ahb_system_group;
`endif

 
 /** @cond PRIVATE */
class svt_ahb_system_monitor_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_SYSTEM_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_monitor_modport AHB_MASTER_IF_MONITOR_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_slave_async_modport AHB_SLAVE_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_monitor_modport AHB_SLAVE_IF_MONITOR_MP;
  protected AHB_IF_SYSTEM_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_MONITOR_MP master_if_monitor_mp[*];
  protected AHB_MASTER_IF_ASYNC_MP master_if_async_mp[*];
  protected AHB_SLAVE_IF_MONITOR_MP slave_if_monitor_mp[*];
  protected AHB_SLAVE_IF_ASYNC_MP slave_if_async_mp[*];
`endif

 typedef bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] ahb_sys_addr_t;

  svt_ahb_system_checker system_checker;

  svt_ahb_system_monitor system_monitor;

`ifndef SVT_VMM_TECHNOLOGY
  svt_ahb_system_env   my_system;
`else
  svt_ahb_system_group my_system;
`endif

  /** String for storing information related to transactions to slaves */
  string master_xacts_str;
  string slave_xacts_str;

  /** System configuration */
  local svt_ahb_system_configuration sys_cfg;

  local int log_base_2_slave_data_widths[];

  /** Report/log object */
`ifndef SVT_VMM_TECHNOLOGY
  protected `SVT_XVM(report_object) reporter; 
`else
  protected vmm_log log;
`endif

  /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;

  /** Event that is triggered whenever the hsel is sampled for active transaction */
  protected event sampled_hsel;

  /** Variable that indicates the current active slave id, using which the 
   * sampling and checking of hsel asserted for valid address range is
   * done. Also used to bypass the data integrity check if no hsel is asserted */
  protected int current_slave_port_id = -1;

  /** Holds the sampled values of hsel from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[1];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[1];
`else  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[`SVT_AHB_MAX_NUM_SLAVES];
`endif
  
  /** Semaphore to control access to active_xact_queue */
  local semaphore active_xact_queue_sema;

  /** Internal queue where transactions from AHB master are stored */
  svt_ahb_master_transaction master_active_xact_queue[$];
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_system_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_system_monitor system_monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param system_monitor A handle to the monitor class of type svt_ahb_system_monitor 
   */
  extern function new (svt_ahb_system_configuration cfg,svt_ahb_system_monitor system_monitor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Sets the configuration */
  extern function void set_cfg(svt_ahb_system_configuration cfg);

  /** Sets internal variables */
  extern function void set_internal_variables();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the data phase signals */
  extern virtual task sample_common();

  /** Adds transaction 'from AHB master to IC' to internal queue */
  extern task add_to_master_xact_active(svt_ahb_master_transaction xact); 

  /** Adds transaction from 'IC to AHB slave' to internal queue */
  extern task add_to_slave_xact_active(svt_ahb_transaction xact); 

  /** Gets the system env/system group */
  extern function void get_system_env();

  /** Process this transaction and execute relevant checks */
  extern task process_master_xact(svt_ahb_master_transaction xact);
  
  /** Waits for transaction to be accepted */
  extern task wait_for_transaction_accept(svt_ahb_transaction xact);

  /** Removes transaction from the active queue */
  extern task remove_from_master_active(svt_ahb_transaction xact);

  /** Checks consistency of ahb transaction data with memory data */
  extern function void check_xact_data_consistency_with_mem_data(svt_ahb_master_transaction xact);  

  /** Gets the memory contents as a byte stream */
  extern function bit get_slave_mem_contents_as_byte_stream(svt_ahb_master_transaction xact, output bit[7:0] mem_data[], output string target_slave_info);

  /** Gets the address banner string */
  extern function string get_addr_banner_str();
  
endclass
/** @endcond */

// -----------------------------------------------------------------------------

// System monitor cannot be supported in the INTERNAL ACE TESTING at port level
// This is done in the tb_ace_vmm_implicit_1m_1s testbench directory and
// the tb_ace_lite_vmm_implicit_1m_1s testbench directory where we mimick the
// behaviour of an interconnect port. However, these task need to be defined
// so that things will compile.
// -----------------------------------------------------------------------------
`protected
W9.LKTG1]cD_.0cJH\[<RWJAdF.P-WY:6MGO^PeY--g@)c<aA(c7&)3F1bf9G6UZ
WCfbf=MR=[/94&CG8_AKH7T6G^V#b9\IUY+gB#.K0;B+eAAY6<T]KUa/,]aCL7T0
5,W;U->QK@109E\=\#<WY^+P/#bG_c6K[HfLP<0@<ZS8RPVV82_;>>^:#8GF?:1.
LRGQQ<f<3[S;HE))dR<eg(6G5<#4YSLPQZV3C[b>&VC6&7?.OU:71711V&V[<&[#
R34V^=K-aYDgP>D[aN_94O^DZa2GVL5?&\.gO;5KKIX]]Q3ARQU7DGM>+:ZOZ;\V
AW[LVH;I)?SAEYWE,Mf/2(FE&aaH,F/Ge,&:83AK8NP6G=/8f4-SAeFG(d)<J\EO
QV41GDDY3Pc;Q7/Bg.T:R_f_d](XQ3daX2^(.R\?6W:[6T465:N_B/J-J<J/._9e
<Qb1E00<6f]2^OI[)A?1/N:e>If6)6N#;1P?+/+^:1Ed+dR^J1ICXb)MY9b&5F_c
16c+)S#d-3;LSK&BEE_1>H_Fg:S)a8G0?=gK:;D:@^;_@)cOYYVeY4MWN6)UWAFD
.B\agK7AT?[8[2CCH/)Y,71=Q;FDd/VY9S1ERa3a+b#4_^@g2gFJZ^d05;F)Q.EE
Q@JdW,7&./fA/:)LVF)EJ@,A93NLe+=eTPJ1,d=NB]fb=BOHUGTT^6cM)\/+JRE7
-dg3016.SQ>U_f\GH-ffg^S[Pd1QTK,e8Q.cH)<NV1YbH$
`endprotected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
IZ8X&M4R&Y71(///+_4)85>bH9#eW\8/Z92.7J?ZN<>5QgSI]b>C+(XE/.OPa.[f
P=4Wcd@ESY0b.A_N7GfO1GV_ECD;OSZNVcHPP]_acf^9ND#Y+V@0P#:SM[C2b^>J
E<e/\+8=eC1cc1V?8I&VA5&5&O)g8H>dgAEG:9Uge/3))8L;\3VFF8X\fceJ3>/9
MC:V>CJ^cd:YSP0W,GY=8SR<c@N:ZYbc&[<#E9@N#/YPEBCR\KKZ&(R&@f9gL>#N
DBcAVfF>SJZP?C3MdLF<<>#(+4Z;VgA1?Z0ZAO^Gf[T\6_aSa3f\,ACgT@2L5g/U
f1N_\&Q7\W<]FW:7S4[RJ7WZ,]Gffg]+;#gO)-,TH^dXg\e\SJMe/,>@SZJT#J<8
?:#9D;SKcXaQIP[C2V3USB;fY2V7d.1HT+c:Vg=QW7WIN^+VS@PBB=D2ScIC:;&e
aed96\H#LA:G)(80WGXCX2>K0J96Zb5\E_X+C(&9A60;NfYWY81W8.G,fIL3,VQ,
aO#(&NB0^,@[XW2HS3?bH(f>;N1fPSg[R)=c10d(7P]S^XMYf6UV>5L^X)<2-/5W
CA^U(fH-WERCIaP;K>7H2V^>&@1Z1d1-83O7>2]KK:)H&SVdb55W;7N,R9\cK6cQ
RZ#W]B?G2dV=[#A8<(K#6Z=F4LTPP&0F+<\c\8+faWB>T\&R0+B_2BLG>6]UA>[c
R\\XG3Y+KU;?=QVYK:=UZX_],.6gZRE-0>Id^=K<(T;=VAOC_fR(N(I/M6UR32:7
S?0CF4[&)(=7?(:UGV+#?A<Z3ZVRPgNSF7OLX#HU=<BTGBQFO5,4YEW0cb79<^3;
H+Y]=N#?a\H45=&f3>=3=b^0W25\031OZ/VEPWGB3HL@6QH;NG[6aFfMeMYQ<T=Q
\9(N]c.2P3T#R;FFaC-S^N-O__.Nd/^Q(b.EF#_aCM+E3eU3>2G>+@1dK<NUH[9e
e834IX:cDQ+?WNEA-7K-<S5M#PS&O1Z-^#e4C?-)&=L^2Y>+3E8B:K.LfF[RaLGP
I-<U,ML#EM>@E\Q9VE2SBEF9YV8J9N_?]^]4GcIa[-LQ(S-g[[6gbO&7@+CGN3X+
Z#AJd;:<b1^4\OR&9,P+Re^+)UDUS5MZ5U_WB/F:#6/?:?/=B^E?(S>W,#4T,Eb7
=>V(171b4](:+3<I01bVd1E\RMG](>XZT]0LN/CAROB7a+@Kb/Y.a(d^g0]>B,Nd
cP2PV25LFK-+]e.b=M\L:5YA\17G9FSV,b=LO4-V(GPYC>AQ2d(317<gU#&^_(?.
d)Y&O1/R&1KK15.9;,=8)..L]<Q7LX;_YKDDAAK:.^[gGePVF\aO\KN:,T\CYd]A
3KdO9I7PDMHd7f<K?dD5b0(-48>KQTIfd&c:FX1.:?8?2>0Y(4)[B&<M5-b-R52<
(=P[Yd]O&@SA5SgUXCfSCM#C77ET\RDPeR.1A<)H,dL-UC/Ob1L0fBe>LNAcE^8=
[XM<;,SdU1.3SMfCeZ4,9+)ZbIUGA)T]7OWYO2[^&@Q-[gZ?K.VNC:+F=Q.11ecE
3F@bLKA@Aeg=7^2.cQ#M^#OY/@f_dOg9:\Z<&;4RH^@^,?-Q?_Hb>#<E43HEe<2Z
,SSg;-//\CReX[eDB@3Y?RO\:dC?NHP\FPVE+9^_KT9)QgJLWe(XLFX]9PU>gK(a
99Z<;PBaB(FRT\(_S6;Kg8QLQRC]BE8FEM()_[7f/]>&bZTHT3PFf.6:]cOd-[JC
Va&f>PCM0N>bZ2=U_TV9]K27C,1>X<WBO+[:#TO/4X&1cY2.6R70L4HJORg?,82)
=^X0e]+AP.(dV1Tb5@7UXTSS2]U53cg=GRKMeKS=DSd6&QC68(+[,d^Z8+cVE,S)
=eX9D#Z)+LD^^A1>bJ-^BGA8:/c&O]#:Fe(2)_?:D;<DXQ4^_9eZJDDRI^UER-TS
ALc9Y<,@9IR7,GP)BP;4N8V2#&^SV5IG9_10[.HGXIOEC^N(V;F8[4eJALHG:03U
6QY+N?[6e6)e&T+CL0@d#4Hd_#A#RdA&K/dR9\)S(^#U)&PO)f^LY,L__dE,W,aP
Y=4(4X,YY?Z)(/>BaE@\FE,.GBX4@V/7c5fE,[JDUg5K71>AJI5bcBB00,_ROgN/
UF=&D@f?_+<F+P_XUb9PP1J9TWY/a+:P1,6PGb5X<:TcGA/d+d90(_I931T4ZR3g
50^2+,,I)M^9@\SPV:Udg3K8V?g9F9]10OU878/5QQ#VX4_ULRC/5O_aC0RJQ3H=
6LbV_70C/>Z?;CKWYA)bdZT9\Rd)LAa6M<\@5VT;f?@0df]aUW]SE_#PWNYZEF]Y
,.^NeBNL8O;:;@)B@CH=K#[c,bd]6D_6])NXM>T9L(PCEG@X0NN.+EV_[?)8TS10
d:?f).GaNdDPb2g)+3E?:+<RHFVOYPL9Sg[bIU4g@YN#Sg_8F?aNXcbD/3[OW(6_
.d3DGe3/eS:=g^E;=FHQB0[_V5Ffc?3OYLd&,06/:[=_TSI5CMBISG(ec_NR7f7H
D:&ROeIIAd[5_297?c[8ZT+=:8.a+W3bd]+6\0BUN8U>:dG^WB<,M-5S6dE;#HDG
I^_BX)[QQZe<)2T3K^Mcb(@fbZ^CWS]9c(_3&,/DNT-Q-3:b[(9?CE(/>.?d5@@X
]3TY:I>YTP/2X-/3V]6,WU6+MDPJ4:4N4RV5J&L^8/<G?@gOV62Z[LYfb:O18Z?P
a4;##,=JVY45-;D3?&H8>RJPEf[KLAg(6\F-G[?b]K/f5KZ&C^E95EI;=?JT95L6
MYA]_\_d=e^S9f:bNdbFBV_B.P\MGIT&??2N]XJ4\/]OgYad6LV3fL7_2Ne=>,C#
#:4R._?YLY(?6W0QML]?FG<W)G]&>=@NF8?>D0VfY6H5)?Ka5+e>+A;EMK9cAd_L
/051<Kg(d,+-1V3I\@MY<=&-7@(cF^>4C8J2T1)Z0&DKWb,F@=J?EJ6=cc<^58D7
];g]Fd3;\0cUJ(9/I-,5ET448@ZK7YYHe,@0[XHMX(X^2EDBU0L8H([VL0D@QDNb
D0M53N.I^d)\R3<BOe8cfUffTeP6OXMVO\(P3@e@[&9-5a_bTKN-P21Z9@WB1NVX
X.5]Q4T;]OUWIIBU:3\E9g-\HE<bW_23ZE&.RQ2:M^G]K\L4\2T[SXXP#FK7LB:)
5O66K-UY3fH5+OKd&)SM;-Z8/#/XebE:[O5\4FMWT-Z\?=Y?0H=-0+9,;f]BJd)E
C>-OKL?1<3YRa<N0eMEGH@/LdUgNc6[R_B&Y,4MEO[_RX^>TXX+G9e6\1H4K.L6,
#fc#BB-eS2-/.-\.b9dHV;\L\>9:J7CTJ0\Z>1aHS[1I:IMecBVZ&=cUAH<6[SJF
(WPb.]69&.<g02=de<^K0T[?-a,#<2K+_cd8@\D1P9PHOJN2(-L]H35BX<TCF#>^
K,RBO0;,1(&-+U/PHe@&16?AT1(3[DD45@2CLc81SY@A.N#/F7OBQ5SG+4RH>X0W
+TI@VCIN+eYO+N4@?X&g:RU#UY/Ab[9_PZgaf25SRG=cS(6&\dS.gHF4bYdUOIWM
&1[B^BSC/g,7Nfee;7))N,.^JM&F-CJ4^e_1U;0HNF3dE7.gL[-K6QIPYd<;UKHK
XQ,0ODg-cO0.^bKJU[UK>^eVQQ.gI>\:L]X)bd5fOV7;F9KB^-6bKC.8Gd3D_b(d
I6K>YSZE]Yf,HCbF3(FQ+?DebAT+NUH>VCQ_R\YNFbd3Bc)ZD>-e^#F]C_:)M,Z.
J?_EO8bD7B]DBZPBK5IP7IO[PL9R3aOAY.OS?:MdGO:T_<IE=R#3-99VIKQ4F2a>
<0W@7).I0A/CcOCEb61W81.2KbT,^,a@d[Wg2H5L&&R3KEHJ/[;0+NgU])?K:O5W
9.caL<WBF4e+RUX<@D<6d2AUXTYQXW#2-H&0KT7\FV@Q;]@Z\7[9Ug@Z_>@U9+S+
G+2G;IP[UKR:#EVOL&J1(<(1US0AH?(K)=KWWO:62(Y73.f1R;73H5N[XLgONd_S
>HC[(&Xb.G2(1GRcf(Rba/;08bAJ1B@R,X/cOYTIVQ=C93R2)eETVQ(#XD\Lf]GJ
-FLCf#&S3Yb-KZe#\;^I.9R_N),W0S^;I?cVgBBZUY<Sf6H:0S46_:R>/RbFL9)U
3_/_b4aS6-UaLUK8#2YWT>Z6g7,b>8R7&.1SP=[>D#AIf7Ya(d(&,fJ^T=2.c(8\
5f7)N658g=GZ#OK;LDO_F3YE3U;f@a&T])G,)[0?fR#2bMea7EIbb5(-,@[fVILK
X@]>NXQ;QY,ZY=)b>JdX)_:/Ldb9W0CCK=Nb7#WVQ=aHI;g(Ia&9Y+0(\HcXSF--
7V[d0:SZY78/?d-QdR00TYJG]J7QLO&+S[CDXd96cXF]V#.+1cUM3?&-=gE3FAB[
R25JQ,CDg[f3\Q+I#)eE;AW6=)b;AI=[FK\/S^U^KJf?2cQJ:+RCb?4/dODQCe&E
d89<WE8bVe1b[=:)0:(,279W5Q1gcG:ON4g-]0LCO(6VI:f/^MJ)[NH3Je3W)SYP
Kf)ZbVC2<5(]A3CL-HaK[a/^d_RROU,=3Kd-BG#d_5Qg]^T>@c5#.B(,G8&5.>e.
eG3PBT9/;S;c)H_LgK=R/7J>#-P=gMN,@.)0[f@Ce>gW)-0K1?U^Q\6HeTR](9@O
^ES9[7)<\Ma(/B4AP6KUfA50ODbR4VY1=bV]K_6(BY;N3)>LOBPA_b9G?/0McQ1H
O#g?E9HB1GH2MU5T9S[Xb#@5=fJWOcC3Pgf5e@3<cU+T_6PQ]_D@863[1?5ET3Pa
KdE9+dP58O][3P19T2dP=^3Y)9EQK_,;1S=QdW\56<8/EL=P@@C70WP]?9J;+._G
CS<gL>1Fd>8bc+4e.UQ]ITL+KK4G;QQd[T^#=(N?cf-H_)P#AgOFV5](7dGVfR7]
2XZ_Ub_C.+LIZO&#(1L:)VT5gH9Ne1Obg(aM.d0ZK2/cb:N)F53>>dWC>UXACeLS
>5Q>HPeZeOLWcPLR0>cY;5RGg]gGg.EEMadbA^VYKA3D#D(84X^)3IQCd0;+TE3_
JR)1FN^a35gF3_],aK5).>?;TCBK&O-F6CYUOMHG527I.[b+Z4L;aNf4JVW;B;O3
1af0afY<BaabO_/\d?:9=T+]O1THRC[/>ed3Z#fO:RO@UgBe#Xd6S34>^bcLe8.c
\aLY#BY[QBOJ0(Z@^;,[aDWW_dL=+ZYB_3-PBPR/gaVK4S=\_(CHB3_ACZQ(Kg+:
G^._DT2DgcH<YYY(ZWD[Q<cgQ:<0YgH2b&#/FV4(_#1F9g7OXS/3e/:)VNHf>SX]
_55/bMQ?gQS]YGQ7Wa,1KL<ZgS:/4X=[<//FMXQ4JDTKGeE:WK@2JCC.gXG19F1C
->c(dWe)I;^SYPYg4@aWOaS^QNf_/<Ae3RPD7^0:1H#VB;TDAW\?S9A05#J40BO_
]XXe3DHaGF:=FJEf<:aK4,<J=K<VR0;?+FGA2P_WZ2N&5dH63+;IJ\1@;W,6><Tc
-gWaDZLPL8.GFGKbP4/F\G6AaPQBf(]FXQJDQ&<)8GaISaU^U1;<,R478#6aHVF3
1L<gD(bPQ@P0H.@7++\U(0KCBO-/=SV.,a:NTBR128-Nge^?(E007TDgE8H&#L3N
A(^gS[<X<]Kc^ABIg7N:E;_6XAU4M@/NYKfe?#ZGcBX902G.cc(UgNQMcPc:ecP,
7aUIZRZ)6Ff&?(9,4UWKH5F^65;Q&</@,5@0ZP^YMdb7<8UP_>6)3,Fdf)KONEK2
2W&JaU5QP/g?:eJ6X2VeX[2A3Ob/-&QO9FLeKS\B;>/XENA_5..NJ,I=>?Y];WY9
AW#X(&fVGeQ-DbU)H--aUe=RJS/\S6Q.7YF+.8b\MV=UVP4@b>>.5A0Ed,Z\[_E]
AU9[Q;K<#Q4E\(\5b,#+gBg=75B0BV_(Z)/NM+AU,JZ_5aKVD@;9DP9]\UOKPRJM
Mb9<?D5WN1F2^BXN)3A\ST<;D?TX)bc&9CLV_gB:7e=+X&8](L<91fbJ>g_)XY+O
4J(S/E0-eg-JL=,PZ:?3+42+^P1?H>I<7L;:BTY<=GM\Rd?[3c(EW-C_8E(]<67-
5RY\^B35-=[W28E??ZdSX4F7(ZE?S(G\NIaOJ.d92dU.dETU5aHYI:+XEc820-KJ
0e0TbV&USFJ6N&;T)I#+3e/@-L871B(bYE:9#14F/]E?IEFc<N(M.YTJLAERSZZ+
I[gF-AB)/@Q9])AQb[3U?^8fC>_H\(#5?.8UF;f9afIEaF\7W1=[_68Q\C^;gO07
TI;2=QO2\Q)9d\3\A1-=HNfDH>5bb;f/VG>],Y^f5WY9D+5Zg4gX?8UFN8U69Jb=
\RGEOR:Z)]]3L)b5S.W:7U0f5Za_P[A(-3R._A[YIUC8KFBJ5ZTD[d(8E)/:SeD6
@@IX(R5EJI0+QH?W,b+bLcd@8(A^73,YD-Y#7@\]Y]IYEc=3f7]E(4Od+-EF-[f9
HJQE@RU,AR2DW,HfE8cSFA5#>TT<W:OcX>VDHRP,e]_N.&UU8EQI..JPe_KJKCW6
_1B0J^R+20QEP<].6>A)NSG</S#Jca2-#FYfJdLAIYKS<MI#/EVXb;29ALZTHUaX
HXCH@=MK[1Q+d\UG#4CPO1a4DEDQ+3^0:0fV5CGN(0/L(T8a>&UZ=cRR5b#14V?W
G0be12afG\N+>=4>)Y)WYRV5G2T84=]=^+T7g/)2RY@+G>V=DcV_XU&UL-a;+\^C
gG)M>;]T]ga[\+KA4XGY8b/C<Z=0X[.\YLQ&2G=U9P?bg5cLe\He9,M-C[Z;\g_D
WT;:OSL\&)G6AQa;?d;OdN]7NB66G_;=;;;g2U.3W4cY@AXcID[J<@/JI+]\,eYT
8:MG/-bA0=V[aTH3DY?Ba93IaH2:GcQ+)RN.54.P^W(3\\QbO;?3aQI^WU?OU<I)
3D3-\7GDcX:FRUfIf9]/aF68;)Rg+5P4RB[.]KJV,aFE4#8J,0@SRHf_61=805JH
;C_dUWG0PGM)US6VVQ5:YQ1W)23,S,&94X]8C,EEKbBL3\;&]I3,QRd.g)N?5VE#
]58#S]f7;Q:b[P7Z9P0ZL36895?A4U43NL/]1/G\GHbcM&:<UbK.WLf\QS7WWDVS
KB3WS??gOg;01Hd&WAS^IRUaABa0&W]&_C69X#FCM5&E(2@Zb;IR@IX-<LV52#(Q
ba.:>6ZV4F?6F^+RJR>>=I;80II+e>g=JAA>aaX8Jf98;)Pa5FBb\N<Y4SKCPE#H
[H^YPHLY;2J+DGU(^6Z&<A7-MfGaZGJ[b4EW]]eZ-fODBY+T>bPPfG^aRS(I]EcM
+#S&KQ29,U4Se8R-I^cU>Q[Tf\dOd:UD8eYc[@XIg\:@B#P6CZD,U;)1\06>VOeZ
,OIT2,XCMXWc&#Y1#f^();<HbC3\7H,N+/-fK:,+2KbdR9T1@-^#MaH13CV#?KfT
[E#Fcb-5ORVf+6^<=..T^GSW:bdT?3+\O,6Y0GE7+=:XO9=/Z,/:ddd^+M9)+^X>
B#OX21W_bTY]TeJ:F^<_((O1^@F1<]0XW&\AU[FeWge7ZN50YN1_<YMLe;[S[&_J
T^PP&G_=(N\[I11LX.,X_QS-BHS?(b78[S1=NATL9FZ;[I0bTDGcQ<K&.gUg+e-G
9aXP<BJWeN7&.\?&=N0CI?10-c,>IH&?2@3L83aV[eSKcgA:G,^W5P,/fX4f:_J0
MQE1cGG\YW@LPT71/,C39TXY@c[,Bfd=E)c+Z.)EJ\KUE]PB+S#/2;>f1),7fT;<
L#5X/dP(GWXV2G-R7#:JQ784_7Ub2HcT.TAZSf2B#(2P[YebAU)_YeDZ].^\AV^[
a8M7:[UUR.Z1.H&_>)4=UZND_3D<6g3G1OS<:Nc_-OCGBGK&G44gV4=9LU8B\4)-
24K;6C:7W:7/-\BQBY&VE.a.,f+H&_R3KXUW><,6;16,U8<gX.e4UFdfN>F(9aa>
#aFFf._EID@U]HgAY6?0G5JIK,=7TDT/cDI]^67UEeW[E4M,\\b8E>Qd3d[J;_0-
7P1_MNE3VSV\;.1g+A2-c53[7,,-6K._A#2,[UQ@aM9+VeI2H/CM,f48@CO0B,S&
QUd7ZG_S505ID<FbKBQ)2E#[:-B,dU>XG=,0ef73Y>NJa;=N/BMa8Z6Gdg,HSOK:
C\gL31_:7,L2dZ4CJg.cDEF]1e8R9_BX@&-7>[7faR20;B0VC?V?W]<R-;JK]R5#
]L>-(0gQ0<KZ^DY7Z\]9<IcU<KU0C>d1XNOG2SY;J1]PM#7,IG=M1,U0W;E).BU[
0a(D,P)>.FLc0J>1U:S0f7#E:-0#8PC0;cUL]9c/9Zd:#7SO2_(>f<#^3?0=EH[)
CeE+JAJcFO>;WeM3/CE[a>S6_\OT,36:/QZ2dQD48KD(N>/B@BS?U4#Qcbbd>H?D
I)8Q-UE_CNSXJ:WGWdJ:c6B5,\3(K?LJ0238,M/MT,FERYTeH4.6&XUeTe8LEB53
A8LK++#CRFa):=0b89SIDAX.d/)UK&TX/X5,<X1R#GB1d4b2N+2ae9>#/+KWZ?^?
1OO[PIb2]BKN,cE:SAgP9,5=-74N44T#.UN,e&&9Y0JXI:HbdSf.3F=cM/BeOP:#
)+MFN.JT(gfWP-N?>#a(5Z:@8)TSZ6D[Q&L37R?HNS:+[F^9VMK1LeJ<ZTJRCBE3
V,,<7QA1TFWCGC_?U(g]V-f?CX@PfdZD8VB?aVbN&;K#_8EXTZ98^JB^BBUJK0X&
Q4E\1TZLU.WN9<&\2^\C]98&A?f.)CAXR=gX-9/FCKf2(8RFVOQ0gUX>+PB(a:)4
N+57-L1,b6UAXF-L8^GaC:HO2M4(fT51&D6SWF6BT1YXRb##D<0c@#FZE4[0QN1M
JX_d<=7?/&B=>TVDI9DZ_&Z:_?.BLL9R:0HAD>+PRdZ]_7\BfJ)@/g6^?bTEYJ94
L)^>TDNaQG-_dR,<<U?-OYM+Y/<N6NTcJKP/UAF1Jcac,</\fIDGA\@=J^?>f5b=
d3EeK.Ef\g+&Q/I&&0L=T71b+a<[9EU()M9H_C&dX_IeT1G.-]0PEJTBU.I,gM9)
[3(::^4ZLFDV1-O?LEf&WWfI0A8W_Z+SO^65A;XGL1&97;aePWVfC>=A47c\5,V[
38)VYbLI+IURP0+aY71S1[:gB97\8U<P43gEW6[>N2.I16O(+@[QVOAL4_#-\>V,
Ba)F40M8?<D\<[9Q,GBa6F<c._\]V51M56,9b@QCT4.aJFcPR^-GcZA.,Q\IPg&R
8Y\DXcIM=@IdZD/I]-2/IdeB4IE/QL?9U;0aO,I+_Y8]KU7U96I:8feP5\^0F<RZ
IX#^54OgPGN1WaHe_cbX0>VMg;JDS<?f1gMXbNUeN3d9[a7f\/O=TgXO_=BB:^B<
[f^HUZ3c^@&4VT^f9dD.=C+@X?Z[MN:.IY(D2[PZFOUL7-#e&7ba&7X6C_N<159Q
N>#HHB>^HSd3=0/dN1&R)>6]-S0Wb#[\H3=eC>]9Q.g;B#.DY1#NcXgL[EOc,P8W
<TJ3]I.)=/MIcM/CE8eW5g/9H6-2EIe.Q-c0CT.ODFe9YJ\F;W6bQ2E,&;P1dXH:
E0#8011Ha0DKb#@:-]LD9>e+W@Q^N&Q^)PBcPZcCY<./RZRH.XH?8^-H1K0&g7_8
[[.eKF/RM#cR#-KTO76.)>XCZUad>-(&]N>CVY/HA-1/O47F7Pg=J>0I5+CNg\\K
MdNI].1@(GFN83E0-]5#4B)8G1Lc;1MV]CMe&cR_6A[T9F#IEceDcXM(a;BKb@=D
37dR1WWC[L8-]@DF[BH#@^1DY07Q58]G&++dX3?=UE)/E,U371bN-MDKR]PFd+38
DTXVF9.)7HDH.Z_ZfMUD?II6aJfdWKA#Cb#feU)K[2/7+NADDD/^cI58?R3WEI7a
g2aFbCV4JHgQCE4_6U^35?Cf77bT0T\a/F<]\XE?,@LfPR0J6?[Q1c.cBMd3-C2a
M_6e6KK9RI3MF+?/8]BG;F(+X,G2V2/M_/P(1d9WMAUYLL+&Y=T[6:a(/+@_UWCY
<F<NRJJB,G&S\/d+;fb@40C[)_38FY?X:0G9-P7H7BNMGQ[;d:HWX;J-D_CU\MF(
926HXEWXNVcF3S_+UVHVS2P\_eVUN33)b6[:[b3P1I>]eMEEPWI:.+TGc=8aY@[)
>c.PY)9E\R(\Q\G#SFFS];e2d(1QSU[;N?&HA\U@IB>ZST/S4VJg9/)SX+W,EW;P
0dM/BgD9<WQ5,)PWU1C?f;&EBP,QQDO02TK5//2T36^\H8FOaD\g.cdR&;)O&<;)
f/8+,gPK>^4f=SGPeUM?(4_<+XP>f_/6A1/,G.,U>SaO8>VV6Y)<SES@L-SI<X8g
8+-3\fT0ZUFSP6O]a#ea,P,FSeSAe9:4<;_WV4-.=WEH];^T-?R6bD\EYWE.63eY
2M=d^GId1>MR;,.]KL&>KIFEQ,7BOIg+C#bQG7>^2[)B<OD7V4#WMUES8cW=[/H>
7F>UJM^0AM?@g\36U:Bf4-dNd=3Z/5N?-CBEO/DV\9L;,7XVA9T_D4@9Jf?MEFEN
T.D+-+TdK>1O.\,_,VbWaI+]2A\]bD3TJ=B9/VBgRSWX;X4/d=:[UN/a>@fgf/dQ
2;dU:GW/J?#b)?H4=,@@FU1PRT:4VPX<Ac>0Y7gZZP.46(8UV+Cf=@[ZKfYA3^8,
HX_+@.0K=M8^99YTT_CZ7C])UJFYYDXF^0)Dd>?a6[9+bZ\Qf9<?&_P-<.^HH#AX
-?R6LOd4J+08P.1TVPge&/2)84b\:8@1>C(R&_1P.CaC2T_NFQ]@=Y[A:cD;HSB:
e41fDSXOGV#&faI:E15.Ba5C\DO_HG?V6S+7,=b,V?-Sa(\O&F;?+H4FUY2/Hg;W
g/&Z?28(FYT)WPeBH0NE7b34OGIWN]&:QaCbW2WQL,S5V#?WP-C4f0MM=^@B[^8R
G3^3T?.\XH@eQ[6IGA[cVb2S;/,^3AXHUKV3fE#VZWIFbZO&IJX3Gc6/e_5bFZQZ
/M>WPEMHBB\&eM-Qd-77DY9/?U=ZPU@ORFb:W3g#?T-cZd44>MM(4I:V\JF>P#C^
+>ZXXDCW/b\FWCcQJbM[dDK?/,V@DOL(V#2fY^e0g=L[-((S9<)9@DRMf1gfb6T2
gg..:6cY.);;5>X(f/T@8(PcKb;4[UY4D2NRIUcL3/[]I8OE+^Q#IEB3gfWa+MOR
+eL\OV2_+?HR<Scf;b3>NB+Jb;<_QcU6/F]@C>cOT+Bfb7RE5Kd[\_+dX.MV/ge;
ODWY.,.OYC;,-V._Y)PSg^PD1+43>]S1GRXGe^3#KD#gYT.0(57;f>0.0/)0^WID
\a7E6\&d+J,Vf7)Q]-<b.@502F,2=O#+<DE(92DPFQU_)\/]4ge[J^0)MFNVA1:#
caVFS-3B)MCeF2XMQN-MR^21+(RNQ6O?5.VJ6QD\2@Jf5ad9^Y=e&NRRV0+HI&_R
3YgGMI9\<:4#3]^KV_Z[#A83dHA(TW(Cg\1SA((3I8#c>GHaf?RKCIFFVB3ZZ-[S
6f\HeR_I(PKF\TK:YHMI=Q2a\)J@3e^^ZPFR>;R9gIcQdXNLa>3&dZQQLbPJ_cc2
gQ1<:+6&4c#c?Z;D)N:IM7JDP):PBcK[_84O2BPAd8?=Z^#F-XOeg(,eEU>KReUg
;W5O6DYcCKfXBYZ)SNM#P)M/)5Y+EO@DQ)LN6^d(Q]C>8eEbCN3(P[M,CR34-K0L
M_>0T5c70E62?1Jb7J,eA3&/BTL&>_^_[c7(9Y+=^396#N]+@b(a3G+N^2^DHPW]
U3]7U@aU1^/S1@aWWe=&e&)Cb=XCHE(7)3;aBJ8bMOZ.)]DX<PVI+W67:FVRQT,Z
/DMA-]LJ2[E4UBRMaA#OHfE3Sa[W::[D0g^MQ27W(<f1)X/+DIAT,94=0J]()U51
IYU,DP#XAO>Y)_;bHg0,<YbZ7-W[9Q7B,GPa022[&^GbdIGGGC[MM(+5-(5VB7A_
L[C7bNcHF)X<A)fA00[PZ(1&L9PTG)MPZ&Y#EJ&<4#:d][^MN.,34(./W@D+AFT<
3Q&PYUb=QeQUN;2T#g?J\,7#(P>Qb_JLD]0Ee^)REQ==ab>(N<D/VZFZSA8#8Yd.
4V0;4<[a+b5e2D0EdQ#Wf+UVHW9\CTXMc;MGT,8eeOLM=CJd0<;QVP<=bBMVe]^+
>J\F[CD)<+N^J[J4Z<W)_FbHR[TW?NQCFaSKX^JCcM6D#50#OaXI/H0dDP2<HfPW
(,NIGIRUZUba35#GW5?9KF?;;aYc36(@<ET-6BCV&[(U>UP?aVZ.]-#Ce^7.-U16
cXTMN-6)N0;W^[7gOc[G,a:IXQ0>&N4-_@/5cH[#\3NYW^YgJWb@:M,TEge&8f<d
)Zc>I]5>V#_A?QTE@F&A2ZKNI@fJ.fK.P1PX_O15[LD&G_0^)g<,g^B>+T3B5OL8
\C/0\Rg2-H5/,Fe>;TT;,Q5-(C(PAQ:e&&N]&9RJ]e8.<)9RN;I@,8?(:YU:BXf6
:c9J1.4-D^+Lc>0MNS\c[Y;0GVfP#K-NYBY;[aYG,BD0Gg?=#FMT&dcLK>;61#E0
eDUJLT.C53_C#@@eF^O&R&2J]g.OHZR1NG11@aDPS/W4P)<)0YLfUJ7MM0NZ6WQE
7@:2YU96TOU_47HV39K\bLN)(:?&)fXLU@J(:C/S?gRE/T#0OEA];G3MIFH[[1^#
^-?;-E;=017X\SQVZN[CGRWL2M_da8)NaTCg@ecRaFD?e4<412e5J?I+L63J3WWP
dF(G_M#[1)b16T2H0PFdV90-@W@X4WHV),>S+YC:aHK1(Ba6SU2,O90f+@OB[_aX
D^a8,/5g>IcN?TNE&.T&Q1,[[AFQM6NN0fJ1J:4ZPK=?),E?L2=JO2/[J/0Id58b
):)?=SID457FZc><V&[CILS25.CaRIES3\b_[HG1gSR8>C:egG]?ZHH1C&;>3WS/
DUPXHN;4@UV/T)^@:Y1d-I.2H8ga^Yc&d@:&g,f0V4-:6K8-;(#-48NQgE42[7cP
R=@:gX_I2:YJc=VZ=1?7Q4e&9#b=9Je\DFXT5YJc4bM5>C>?bfe/8L2b9M0Sb4Z4
IRa,97;65_M]H-f7<ecNZ&aFIb1N.g#b<I)HLY4Q4@-B,CNP8<,\_D:;8:^.YU99
JRUH//d^B9H;b(>J_DbX<df@;3c53T=;_ea?X3HEQP@Z(C0EcSSP14R5-3:8]7ZN
M2e?XYCVRVCNTd]I\QS0(=?(XcO9H\eUfK5gXQ.T#X8STK_D<f/X1Pd_PJ/S+^6(
)T/NK@PH0,PZ<V5\C9\b,V^RMf5b;6Q-9a#?9?,KZI,@IXD^d:T=-^YO&DL2)dGU
J4):.:2Z9M[7;M(Sge^<L:IQfd:=.=5eN2>gVM3)Hge#/MUbK0E6_a8b5>D&#BR2
1g5H<Uf,QLK+.eQ\8#-._fG<f,_H,8SO8LbOF]M7B9_ccJ1C6L3&WaG2fLWfE=Fa
-Q4.81d4,/J5S+R:9USE]HBSX5WRZG86)8O:1BVU(,B?)ffg/(HXaF=7GNHb?c>9
F<3(\Ea>f,0@H;]Ne(6CORIE#\I:-(.7T+07EEL.E5#SWaOP?_L7baBRg^T7E.aV
M;XKd94ca4^+C]9Q#/dP;PA2EVZ6:a)A7>Q<)J8)&&?_@F,;>[QE<SGK9IY&A5]A
<VLPB;C;5ZPTP5:ec^4D_JPV+7JDeE2gUP6NN+LbZ7]TC5>FJ)9C0_3+?3VG@HC;
ZKDRGRQ.U52+3=(1d@26f\afB.9S5gDI0=M&MgNCIgZcBPGg8KW(\g(;DV#INSCD
.O[\:9g@N,^DB-6eD-K.AYMGZ5E#aFA&fIBN3aKZD6_TFgHAaO&.J)JD+ABAK:9&
72\(8-]5CF&?^P+XL;dC<&^=DF4--<4BS3E+?R#?5]G3S/2XYb0NSX<df8M#Z2^]
]SR,(_3QR.Q4E]g1B,CXBTN#U;Z2ZAKd@cSXgeQ61STSZ22Bg7e@#E^8<AO=ALeD
(NGT_,^(RLaKXF.P/f>;<Y8f+T&,0@=FQQSSIPW5HA/\L>?\+2cBQ6>?3-e+,?0;
^2d:MJ:?K&6=P#e.c:E@B<^U1cFBc7&a4CbA:<@gJBQK&NC.B,OEP;80)MOaHVL2
e)]5.HPY^+XI,#IM<T)Z@,QdHK/S-b_E5Md[#DPR]<-..LdCU;f1g^U8O6^.K;?F
GM>D-BZX]gafb&A[^K/-CJ\f/13aA)VGE/FH_HUSBNY;)&[OC0RT>8(3AWBMR8XQ
=bc6DD;-7>&#198dJ0RMZgE:SZ-YRL(aOH9ESTagKCcU=[cUN#2UK[JDfZ@ZZ=gK
b[>LZ2YbD0]B<f8aa^P1AQ_T-VB@-G]0JRS19;+@:cE;cO7.B)&JIP^I;5fZ\=GJ
8W(,bW0e^UA3,Yf^^ba9/J4SDMRTgVFVa@dZEcIc83_6;;/#D5>f,DL(fBYUcLZc
B;,S?8T]2J/@TO0adM\ZA(dA=XH(J2JND(Hf#QD@K@:gL1LH,I6N=[NQ75ZO&DOT
L\-:48g6(fIPO>cFd/#5@Z;MU09fb+8TYIEJPDP9[-A+\a4H>N?1eb(YcMc8eJ>4
@P/6262c0-2M./#Q#e(@Ad[K\&6D>;K&cXAZa,cC9UL>0/-B:/.dcIVUg#aPR/GY
-W=gT5P^Ec_O)JO?B^PdY&]V<03K+g1X^T)/5TQZCI(?G-:_0U<-OM,;03K/)C50
&:S,6-b<,4X(&XI;]@EWCb_-QOTD)4A1-L)Da;/)V#61dY9J&d(d#dE,IMTATa;X
B[a4IVf4_OP.2L[9V.?<Bc7X)8a/fO^&E;Nc?FEPAX\FWLD));-J=dV\Dc3\5dc<
NdZb8?ZAO@acSV>@4<&SO,CLRR/1VZ7=(e[eaF=VTOQ(fcgN7GL\;B.I7D\T6E-/
6dSC+HY;9RE_:\[XP.b(M4FYDA+0K#^I6V>3[)[BSY?4:Ue-a,X<8#&)MPQCX]DC
RUD\@N/<ICWcV8,[ePT>DD&D[D4aE?ZI<8.+Z)dI)/4.ecF#7f?7RL,YR@f2F/cO
54MF>N+HA;2UTO)4f[2DD63V;gPMG28DFC:Q1R90VD78;1aNX062YB006J/;L_=c
/ST7X01NF-[XZ5@>a523M#;G,9_F6XR(&,\?.._+U;8RJ&JD>;e<P#g#(W^[1?_T
+d;c&^GE&QU-HY9fV,^[WI3deJcb;^VLDN?D81<S8)Y5;T?#^8f1<86JOONa-;:T
2EDTZII?aV<f>2,<;)D0V^DZK)KC7&;_\F&O_.eL0f[R[5O&RRcCN4,A3eTR,F,>
F3OIP/.A8cS>/Cd-4/(0F95GQg-H6@;f8;Sdbb9g-@1PeZJS3>QRJgX&J<QM<A_+
P&)]cMJ4F70XZ)1UJIf9DCAN^LaI.8Mg5]:RVR]]LDVdaTE@a0CgT]5M^2ZdPE^.
..;/4/<?JV==Z@Zge,e\GTBYBY=HBOXe(T9806FfVeB=bZ,4X&T(LEc,B<?_cL6Z
<:OEcOG0f?/9/Mb,2f(76W[X+Yf-U_QXgN^Q;U8EZ,^[1#4/@F4D5P_[TSG6A-.S
1X3g4Mg77PX8]edM[1TJ^e71;)4(eKNcG_dUEIMPQV5.TL,R)&#9^5C7C8FQ_W3F
MD1cXIKIc2e6aDWH>1MbQ>9\fRW70P/_-O1]^CN2G0U#R;8E.0K)g,D>S;D[I]^>
NI8LgFF4dR9(OF)Yb#30gWI(;H;4>^8Mc;fPWGFOb0:Lga1CJbA:/GUTCH?_J[,,
>&Z^aUd=cNdY3-J?+Z79ed/dJ)eV3+.-B:CbGbQdH:0ec]PFLD(W\MeE\LFO8N3)
@6>M08@N2A]U>RGY9SE0.ae&E_E^CRR3,LUbK\E.9F)35b)7U=f=]5O1Me,^=gM&
)043a3.eIfQcT?&3G/(&^aZAb7J\&0eaA+\=9e0f/f_a)+XegdWYRg0-YEE/2&1a
d->2LJ.ODae3KCBPcP?[BX5T=#/2=@54gb_J=H6Fc3gaT+IgD)C)=5YYR:R01;eZ
7>[=(Y4DOUbHM^3<IVCMY50<,?Eg:NbWQZdS^MXE4H^R2AR1,(6RS8JL2e6WfgeE
c)4/I582),gZ/-13Ga>851D++6\9,e5McH:=XfB@,g1D-ND.\7G8DA6+ANMVAR47
/BY0F\U(37JK1TV(XT<K4;,+R65N1TITQ_>J3L9:H[e9ZDcUgII)^]5=cE[Y-\/5
3-#]P^f\dU+N;S5P+/T6&@)0a6GPBS\D&V9R<TGBP;4_G1@FR#0cW@)R+QX@H-GQ
VB1_?Z8T.D&:DUd1Xc7,AbgeOPW2[>:Tf4ONTP6+8dH^O^(DBcZ>A(gVPaESKJ>9
HG79(S<CB@F?/]^Vc6CDYg;A?^42S18c\O>?a>IaCU\G/VNUOMYXIE\YLSgZ<_?)
J9@F=\:bL75VW;^Hb^Q(MM8L]DeTa2+?c,M^,GJ=RJ_GeZ>03_4Mae(I\<^Q74F4
PPYID90G\E7JdMHf.7-D6A5LKCSFXW6J\PTZ1GfUHN(XX\-+UU6:1b9BFGG1K\g>
fe0<(<(#@RPYU,,W.[USb_4d^)GXMc#I&66c.V:W_I;P+U6g1NJ=HL8\^WLBIQ_5
K^;(K^045F.+2Ya-IC,WPX@5ZdWa.X/0)RRF]DEI]bTYG0a<e#YT7;.eV&YCZQ1D
9c@:+3Gf=(\,GUUEWcVRR6]#\]#fR#-PXd1>/LGL&Z@;?M>0213JQdO.<7c]6Ze1
(c)K/8T_;J]GFgR/[65(Mca5P2.]S9aM67IcZ6c@f.G<&C@K:f)TD3TeR5fY61G(
0U546]U5]WC_9?.SZ]eE\@]:8QCf)VfJ(C.KBM7L4=1N;4_==;R8,27=VOJEgfbQ
?QY,,7)]O.]UaV#YfMUTMB/Hd:RP:Ha2?SR))e-Z+0<Ag;\(Z6[&7+];Tg[JV6^I
d45U\eb#(;dXU=POBQ?PA4d-2/)e8g3_6X,V2Y<U9be+]dISIAVN+75GGQ4X3YQ5
f;&_C+6X&S5W\RGIR99K<^^/KF7-52)B#IG#VI9I[;aV[5EFV]UNM6TN\He[^<:S
@NSM);>S(0@@1]B]\&)CXLAO(:cS7UCESa@X,E5f>b/IAJ2?Q9Z/MO4DX[\W+#76
1L/\Tg<&X;[PT@U:M8cNQFUR?AZ-d)\g]D9UaKFd0MQd5F&3^dI+X<;_\0V)0g17
H:]]R51FN4&;5F;G^(fFXOQ@PJX9YXd&R,d-#/93_)HU(@V,I@V]&Re(+2_UF\KP
e@U4>=5I]L?&SKRX@L+PF7f9JS,1,W[X>G#.?GTT6^JYJYCIWa25AA:KNa\bRcLI
MaUJ@bd[#_U76bBa7aO?5R12[U)G-GPCd##:;Q5a_8HHP<AfcHRV@RH50HPRT:C/
8WL5b?=b8NQ12E7Y9(].G>\b=IG-/D#U^S:C+N1Ke+U#R@.d@ceFIV133FACE[PL
^)7>9RS_ccQ42CZc6E88JL5@+7#T3U=-G(SfaRU4).)3P\T+aTG<?7/:ISJR9E0&
^dG#XY-+ZKWNc3\,HZW&9-KDZPD7P\-\BHf6Ue&?)af]=9S-#V2EVRL:RbB+/>1<
e)N9.JH9@ST<;WJX0TH/M9c5HA/[WK0=>/,LRaKG1T&H_M]UALeZ/QTWH1>PI?Fb
-DfN;3<ed<dQ,WZ@\R6fR,?&5bdaNDc3Zf^VfP3-NCBPNIV]/1_JZ/<:bNA)S^SI
./2c5c=)Q^<M(.GMH5K1g)2O<G/McfCRDCERIAHY37+E]@IPHg_]-K_J+A?PAZFK
/+[I6cd@)F\gdP_).;D63Pb4Z@H4@HJ#.S\CTPc2E+Y0E7cT\907YGTW0TRIWaB4
/B9.\UUgWC2e_De^5G&aY97I=TLUeLAaYAeJ\UfPIM:W2E-/9?Q];;B]^b2M\XAT
:f@>1c14b0g5ICUU@-LOc[6Z0?+_3bI/.3)ZFS[F:gW@C,9>^P#1X=4N]fe<gDIe
U7f.DAW^_U4+If\dM7fJg.SbF+(cZ<b+:J[_411aCIPW2H\1b]b]2GZ0)2X?E1:7
#+BA-&_CDAQ>E+ZB8-^]\&1B,NR7a/]43S&XceNP^b>-&2=:;>F[0T&Y.=,;8<[(
UO-M-D_[=V8HQd/Y0C9d[NDSD,J[9NP4fXQ/.+cQ6,7;/&##O5D+M#]LBNW)R)#E
\I(f<XKId_YW#:65@B@GKF</BFW&6GPJMS==eMK6^dNPR>U^D9.[(6K>ca;0RF<T
)ScOQJg#_aWO.R3^gM3?Ld]TVYWGS&eZ\=2g,Ib6OFfabf\A&ITBFULMe4<I7DFb
Fc])X3PP>)2N,X2+VE4g9cJDRYD>LM-_?#=f#S.O1HY@#F]_VPb2V:6Ec>Yb,/N#
^GaPEN7(LJdd;I^<4Q]>Q3=5X#g@_6DK.=@F6\M=#+3[P9[/7Ka.f],??-=#])bR
78_UcB1g.E9R3EN8QA-=\LI]Nc:Qc4EW]5OK/:?Z6e.b;]+\M6f(HD&g5R3=.QJf
GUWJ@#WX:>fP2E6&/P5.NH<bO[VQ.cWZ8,UeBX<1SV\&UWId1S8.ZGeKSU(V4@87
gQ\OQ)Uf[Wb\9aPIZ162YQC<0U8&;;d[6FOT;;@_B0)O5^+@G^?RTR7NNOZ50_?0
,S-7VRDIJ<OU+)0E7+dA_8]LYA8cWAGSO25AS5B#78G1FPFTDXTDP:fQ>9gSE>73
Z))N>HZ-#N/M&.::;1\#(SU@D]d,d7]LA7->CdK+c;RZEN?=U_:U]f2D93^IYLGO
0#R^bNMC3c(Y67c-+,E[TZd1T2.UHW;C99BV1=.DB613MUX<c6^><BH5J(+JH\bX
g_M#J^Sg0-b.3<:Y\F.0V?F7\P#UGcO)9I;Lf,#/:PCEg1&#ZVC6)R=7RIVY9W7b
fQ1IJd4+S-A^()>LWX5JW/N>K#7U^C=H4L-V5>K0GD^F/<1>\T+#Q+IJ>55(0eC?
?SeMNdEYE._D>C=K5XOX:\LNBB)XK4@^<_eRg&?PG8,Q?GMJ?UU48A?1\IF<eWF#
IIMaT2f>17+^V^Od>-g)QM(bHH6KA^M-7FN&&9GL38G3Xc<&A.Jf.?>O22U0F2H3
g]Peac6U0Ze.Z9+=:NXX4R3=AZ1HJIF7Z,ObbaM[[1>d,JY>gIMb&Qd50&4(SP.,
^J?0FJ81.Oa+;F3JFD:@NL[:SN8/6<M8Wa36?_;g<[TJPD,B_M:3gBKSd5]?Z6<g
fD\fT#P.ePOfKB_/5\[4HgZO6=LDEgSG[4O#3HGbfJc9KY7aQ+4&IHVRbaO]cHb/
36&4GE7-WVc?.CPC)-0ZZ+V9QRKM)4f5=KP8GBD.TEgU,#?^<FH40<Ua_6Q#([;a
(bK0X2KS9]5T&):HMG,1J?aD^-C_>YNV\RdeJg\/@H]\8F=d[J_?:gQ]&bA>DLY\
V3^,VR5E[HM0EY-H8:]ScP_-6;,UA2XTg-_B8gf:+G2T/AZ>QT.B9B?3b,@B#)A6
?TZ^8.I/d\VYCD8LJO:94N-JGc;4;<HK)B5##KE,8e@4a1&)1Mc_@&N,K\\7[^6?
1gQV?dT5LXgKX-70L0KAg/+WBbKIO\MD7;:;@@SV=Y]?S4K\(7<=:8a4F,g8\6fR
GZXC>ee#>HGT)adC0C7FQBB.dJ3F8WLVX?/g-O&2]g(29A,b=XUPVc+S[2?g=Y??
A34_B(U-IT4TgKef(>:4JCKQJZFJ]#1>X:T-?,-Y;]Y4<c8&ggE4e29HgY@^Q:5g
aX6_D=+]\:Ef004B)4[Sf;&a_0/Z;NIE^KgBYI;9Vg1I-5FP<<0H<-=^GF4D.&]Z
a+EI4@4b[7\dDA2N+J-HZLLfa?QYQcH?)YH9A58H>MZAS@?R\JWg>N]GMMO(M4)f
JCIV?[./2B=,TTdO+bDg#M7c0cZ<dJ58B<a@94dG=]RH#H(BOLe_>,#FIX\a&@-P
a8(,I6OEW[7&]3b(_-/SdA.,=6VGg>(A6e:G+FWN:4T4^gE\V1&:UGcZV4_c40a(
^PII0BWN,C>/40S@63GWL1L#T6ECD?3-W5Y0D;0?Z:N6OWegHPTB-1/6SM/.D9Z(
7CD3MfNAP3[L4V(ZF6#/SLbdI1Xc8S=aEWa,&PVJB^5FT3GR<@399eaBQEI:N+PE
UDP1TS.TMV:<J5WD72cU?ET][,<_c/E\M[<c:ZKBEEZ@,g:M-YNR)Y(CIJJS<O&L
<;cSJg+[3BBD1Td=:O6eP_8+\#]MB52geaAS<3WHKS.IbS,9D1Ng4VQ.YUR:^K54
^g8EU.@SN30-I#6I2I,(+21B@9T6E.E>-WWD;^@fQ0EA2+(HcBH2.>&EN-4D:&;Z
,>dZ6T?X<g&TI(08fe;PG7\4;ef@J3.)@Y=71&KK-G(gfJ]BG>Eec<O#OVP5C/ED
<9.gZS2#Af&CA2:NZCRGYe0eF9+B,F#Z4S_<<4W^_c\ZI<RNA#D&^8,XbR@dXJZH
KP.^4GENJ.]>K11ST<=DgR/4Tc)JBKT&(dP?F1,;.d&LZTUe3Wd=E.a)K(Y@PSfH
.D&(>YF.TGa_S8-V_3UYP&\6CO<,WJR7A_?Ma=Q_FC^(_d/NX(ffSR>60IH11XD<
a]d9EE[5KNb/c_0H+XP.d0WWYc>T?#c\NL<EOGFQ@8^TJJI&:(Gc2K^YGCCG.QGf
M.=F4/2/SGccb[b?Rd8KU0gK0\,;edbMT8MCM7505[?D>Y[]M;(C:g_&VcP\</2?
+/;8gCJ@B_8g.OBd5PbV3-1Z=:.Zae]44@/7LWN[^Q-bZP;8_P^]@7Y<C^.cLQ_4
2DE1/;-YU==B5F#<_8U2_8;US.20FNG?UDI=E2?LSc/8N.gN)Q^VL1]JOPZ2)KIT
X7H^-/W,/R<Oe:Y2[aK2IWd+[Q44OefT\RJ#eZ_9TTJP1<@0cPF^gC6TeP20B>c[
YaYN^&V2<WEJLgdeQB+4MgR+6WD9BF.::)XH/P3536F@AdJ]eI^G8U@?^#TBU_G5
+HIANAZ>=2>38/f^LLT:-gQM_gdR@KaTQd.AUgbMCeW1<>7KAHg\HO\Nb&=^B87<
&cfN<fbL/,<9L[E9\&B-:_\#8ZADNA=NW0_fZ5QX)a5R[,N.@WN#7D8.;E?(L3F.
^DIWK:3KT<f7VC3Q((76)3BXY7>+,PP5)J>8(?312XYYG1(2?P7K^MD(9fT1VV,&
g;g71/=.ICIcH:D]UB>RTB9U[DDgY2WV98LU&:10E<G[9c)CfN;9P_MRTg2M+B^c
LJa1Ae?T]YCA()cS:PV>P,,;2:KUebAfKd,>M_T\I5,TLA6]F0JAgUV:QUTB(_UK
2845QM8eTPTYGNB..37LU^T[Q>U)[f^fD@:?<+g0[D]aSLK5O/b]a\5+Xc>;[8N\
3M;5&XNBPVE+?V4H3KZGbUO;.EXW6>=99_T6:=\gHC,.(Y,J@gPNc),3I&Q5S)+R
>B[Q^bVDX;MH<-5/54]A<VIU7D&6DG+P,c7<B6:eYQad-L3]g>d@@0JDXF(@__K\
dOF_E7.^&7c3/DTCNe7X(9>>Afea\OR>P0S)E99H,=]?g;FBTGP))a:W-8-7??UN
Nf5BPSW)RQ.FYKX4E)L4KJ:2cJAe&6L8A)B6W=2EU\DMXXeQP:U9N6f9P6/1VSf\
N^\L;&?8ce\PPOG>S_,K55)-R5,[;SS<R=MK)_Y/)B1(I3UN:6<4dT;c5TA4b;Bc
IaJF(fb6;EH#^XY?P>T<?FCO\#NRc>A)=&b0((PDE5,/[3IeK\_/BcZ,.]4/HE&&
b]@6Ug0A4aK\RR)J/f/:\&ae^,+A&dcKMFY?+0)]#8^.JJZ?V]Q#I0Y+IbB8&gR5
#;N]g[QV[&eT7BT6(_\EJC]G3JN)31Y;d?gCdYT9BO55_c/KHP:BE8g\=)FfAYJ+
Q<\-R&Yc,cPZQL#?R;K3(65@YN8-DV/b<S[SSeb>Bgga/c0-Md,Pfc5Z4]PU./9g
&JZCTdfZ,V1+3;d>RO9J1P1M?9T_EXPX8@@([?5F)JDK+RX\?Z#96D_P\aVDd6e_
?O@Ug>-Y^>(ARL\09/O6((,_>N6#5e<bT^6JX2HO6?Ug1Z)4RFPJ/+.7:RNTL:>L
E_7?S/3_T_>g5fQ82Y1L7-#eC^TLT_G.R@U-28(UWHZgbGK600@f7RKU9D(QEBUA
M:[W-\>GA67C<3?O.MGe;/-bD@<bE[X-;e=>IcU7<F)KcF1XD6U8;=/A<fJSbBFC
+J-],]V;Pga9=9]G_AAcBF6T2OWa^G3=aR(fFN+F#2g9PN1OWd9DFeC8BHU7-3+0
@C[U+WdT;AJWR20[.(c9].eKaX^b[50GMbE\&be(Acg&fTfS4EIT-/?Y/HO3>Jd3
Z_5L.,^=F0TaZYYb/Q]6IXOA?D6f6KK+MI./V\CAU#?9TJ0;N-]5<L4I,\8^C9]>
:166D>)FRa<H9c&4FLeKd@-OGT,MRTbKg#T(0EQD#)5Z<1cMQ+]H.KQ2UV#7SJYG
]e\1PSYd\ORJ=^Se9g;>f#/R?<Y4/Rd1,<2B^[-1Cd<RJ8)K-72YRKEV7)4<)R/6
4Ob^WJd#3e/aWe;21DMWW,f#OC+<g;-/Td3YLTZL]4+(6T/O_1fJfR&0IU/OI#Y5
1O9]HK@Y9YJZ97@5]/3bU.\/FPW0.ce4gE0O3G64@35f22g9:GKVOAT\FJ^P9bY)
AI+P1GWDLc;8bSMVTC\9WV81M82e+1Y=eQaJ=SCSFJ#B[5;79@-WDA(594cYa>@W
RfNZF#V1LV99.E)&)@[_-fC9bg_.)^/NV<\?BXGK7KbKeZ=DC1LSA[?^)5,F[A??
0U08IEg36.:)2-0E;_IQ\IQc0;-SO1S[636F8g4F.3FC(0-_fEXQ;=\FNP0,582K
8g1WCWR=2N7/2P?59AV>M[G(g=Y?N\1We>?V6gB&;#a.9AM(RY8Ed98fUQK?L90G
K?AY30)0g@QSV=@;7O4Id)FdQESYX\c)PcSS_1NHF7IK(CJ[3@W1).d.V&F(Ra>^
6;e6:d,A\&RC(>I+3B5f+Zf-4/6eeXQ-KT94S1=4J)4BX0cKRIL9^P.DJCaPc=:T
V.Z2@AA-c3)FRDPgMe,>:f8>ECDd#+9c[OH;d[dF@L1EUA)LKN3Z-gXQVbW&&25_
JL\Q\7HgP#LT5,=A[Ze+F\EIQ++H\YJ70_@fL-I-+e/Ed3+PPKYQ=b+>70ZOS-\e
(\a<<bb0#1)->D\;DN5P6[G?KbfXRU&ECQ6[WPZ1NKA5L)X4)a0RgJR,-L4bcT2,
U10A:;(I9L6S[20H>C9.eS?<EDJS?FQZ-4)ZXcDF=f0_/W@X4]_IMc)Q42O+7b@A
@bd<9fGENV\+f5.IML:D#&VIL(cPJ(Tdc;ER/3V7TK:NNZGP-UY2CQcXGRGfSIV;
4,L9L_-YJfFa(]I.?>Y2_600R7UX]3NGbgIQ.b(DdN5bYH>bZ3L\M7VX0UB?R4(c
6]ccD:g\G5:&#9_<)CdNVMHH^=5N8V<O?U(BOg73Wd1KcQ_Y=4BAP=c3<X/\f]C[
\f^f2FT;V>L[\c262(6;IcC^K]J7@QT1=NV/G]KeD)eUg=IDV<9?9^6L]0<-YgAU
SL@AU@AF1b95.G]QW_VB&2<;;,dKCf<&@8JdX5OS.YK0H?X5ZYTXQ<)g1KLb2;)J
@\c[9,<PWRIQ4W\T2<1LYPECe5Z)a2(4-O]MMPUMWD52TNCJ)I0JgV5XNcbK>2\.
]W9/X+;U0^S0ZXN0O)Dg>2Ze;H??JEXg]1)G<36aYR#e9D/P4Y72cR@Q^D(-PUQR
ef63_ZI;f.G1P=WM9Ff_b?ER)&+f3\JJ:aEZ&a/L#\H&d9XB3L[Y\J>cX31>1T(@
KT>/e+.E,KJV]:SY62,MN[)A?d^[?Tc]K+/#B\0RH#8:7]g-D=7[8V\.d50FG\4C
^GM>;^]FZQg^)9g0\.g>81GQ3VKd<+7Z6E5Y6_;FA[GWD?c?fbO@RA9N@M52KXZe
_gEM73PW4;b-:X2&E;PPaJGHF[+,d]_S59C>Ma@fY?M5X733>U(ONPFc\Me>;<?/
X7-aVV832V8+GKRa9LA5HYM<JU1Z;N@Z,NTabS&=eN=g\1\HWd3QFcaN27Z?]dDZ
UQ8b1\[J-&5:NB<<?IaP,=^H^#]/Xf<I:O_1MJW\KM>DJeVR4QC;I/@+VO8:7SAM
HE]^ZU:U&gRSE-6_4IP7a04dD5PDY(KQ(X+_E>f4a7YgQ>OWH^YaJ=a^\AY#MEGN
N0cG4]JB.2T++WGBG-5L7CA?[?gXSReL4SgXFdFeH]\[#Z=4_c?0WC-R;.7dKc1G
Y9,,cD^H0;?L++S24MQPNE.C#0J>1=f>ND+fEW+UEJ29SA+QTQJg]cZL)=OIQ3/:
P<J>2-a&0S\+;-QKZ.UL+13-=LDIaRJ@eVfd[Fa(F#CCZ,Z,c5D@Xc3)#F^]ZU<<
E)fDbQBgZU1;AIZbU;CgW8D3&EPBADS;XB2gA64=(#69g]_4IG5)/G=a:8VG>=?-
Y@+#OdL-JRQ^]UTMKN=5?689E0-5D-[C6B_X8d[cU[4[57cgB85B2[;ST0@S&d50
4R,=G0gJJ9Xb.&B642>fadX\7JcHLE2J/]f)\SMH_B^VUE>I^AM52D/7Wb[-;c/7
__RZ-60PM-)RV8KgASfeQ_F?I>D[M<W&4\2W@)d?F+T=QI[.LE5[PV&7:DO+4;/9
(5a74g(__1=9g[-F>.c++>KAWLCSgc-\La8>X0)CO(3&8ETJSR8fa9DW]=BJ2-dU
GCS(G6##DfP)O8&F.b:FPgIAETU(BAS6+;G^VVcER,c(T6(;-\\YZ2^(UC^HUPX?
\4aE=?EJQBB[@#@Q72^V,<_,),G/?Y6GFN84(?If5XG3cUXcJBRQ(=N]>QUM0SGF
OcP-bRI2Xd?0YV2Q@)-4UMOND\O^8T(O(MQX\4)&g<3VC\g516aUdg6=aK6aDLA,
JGO]IZV>LO1ZVA>61@b_CZP\5?P]gg\3(g=?E2TCD&O_eXW5<f73@UYWKcD6Ae\(
J9UGg]I0R8(UcEX^Y3D)JVF3=1(2_;&@/W(W8b:=GW67eW7D?+K0/9Pe>0+[.-cX
ZVaWX#_?=SgTK++g3g&OA<\+DLX#B#^S+QE7H^#_C>aMZ7\VYe7X0XfZ/Y\3RHP>
7Ve0[UQN-^9f;:_?T?S@B_fZCC29,f?0[\_LbAT3UdHN9>b/Z\/#T-dS+7IN<df,
<5U-RdS++C9HMAM-FL/&FS53HP(c:+L=)Nc<T_aZ-&>F]R&DL[<ebad8dL@V)>aV
38dd([\dONCN-0Ja?5f4_GBI,JeWJ_O0MBEYZ_230K-8\-E:]dQ+Kf+Dc;age=NZ
^RQ7QQaOP9e+&4,J_AcZMb1>fJ>e7P(EL2N/TL<DHWO8?g7.W.Y\\3a\9N6V,,9X
DW+]]]6.6<KVfINS7X^I3cO.#Fe0ZC+XB&eU3?T_7H(+^6:]I;?)E3[DJW\2ZdDR
\W8NSV7:G5,NN>FT8^9=Wd^e26_I[.AQLOO8&P-N>Z8N6E\MI)V;3YT3-N8OJM2-
^J^3YJ6baD><[.&5IC52H\R_1/X=_;V2HA8_=+b5,HfHe@WX:G>F<A3NG=)+N&.P
SeB++Y45?LE4XK1>IV2F9=^X1@<XOCEPFIB@EDGf^1O6KG@&UL8O<3^2],TS</X;
Ca>g(?Q,Z^N8L@P[3NVKD,[^0]C+W]A2/:KcM\;^#GW&?;FQ1PC1.D964Oc[P]HD
F.;WBEI:B#<9^e2YOPWQ8bC6.3eR//b.3AA7((3NZ6dC^S),IIH]O^90+De33ITf
]XeTJ/A0^67A<DSe/f8H;SAag3f:OT<G9_,V/_X#N#0XKVP@f9;.X[aB/(65#f^g
0P5G0/a6(WY/T#>#fS;,9A=F/;b2]9S82DNf&/N=:<7XM/JAVR:V(#0:6ed.I:YY
;GT]5)#aW1_05HC6S?9gE0<W;CM]U93J)R(0E@9C(PQSc6O\LVDY=RK85dSQK?fM
CB11&LGO@(F^CdZJARCV-Vb>38@Q\X?A_fQFERS-VbXBV[_XU)?L-\8(AXU-#.6c
b+2@5c-OPO/EU3XV\8BV^e.LO>ZY#@^BNN#]7/>10L-Y:>W#IGC-O3V;W@01B)9,
&#JA=\+XL#[++PYW>JH\d.2MAc9HCg\U1T6Re7./&@#Q3]-KYDdR&(GA\9Q.C?NR
1_@KP/3ZgV.9VF@^fP5cW4bB&g(07^<1I1DEYbY+OQ-E:J9<;FY^f5WQ-5839(\[
=.QK_PddL8#MARAb+R,V?^Z/4F\2PCCNR6@=:3bb<UU7d33A8TG-F@UD.AXT2;I/
4/6T1GS=<bY04-b4FKFEbQP?AM-9ZaTSK4_K(BgMDO]BLP&^+0?N9+O6Cb#@_)8;
;fSLL(;S&;bYgVLMR&=6BfKD3^0]99\MV:J7):TWfbMfg5M&U7fO+14E/Y&ICN>#
f6O+?K9::]L0LFN4<c)K&J(Y[5X(CT-d^A;N9-1b-IW&-I#b;L8R(^TDPT]A#3d+
[(AbTO?RfS8FO^7g3RNAZZ:AU:Y9J9IDW(AW^Gb9TGecfX\0B+;(5JXTJD)\Ue\]
7<+Q0S\,:eP@LVG.[CJDCg7.W]^TFQcL#2TV2LAR)PK-a987Rd6+/P[?D60A0LU=
aVH,YX3(I4aE;M/GKYV_GB?e-7QCQfC/118(RT\-^UP?EU@PE@f(fK-MOg+cI8ea
9LaTL]#F]OZ)a^E=7a&&R.-2MY_+4NRP]POV\Dg#e1ZO+TA=-UbVVVLa&\]3g,0=
a,X26f<1;.H&FK9_#D/9ZN3X=<.ZBGM&/G/\LSCZD2I@R4gPOA:K^Y9R\0F@L&M:
?NFFd:-V^HJCY_5B^L90eL4d#MIKC\]PIJI3.N2O/6MEX-:1K-S33,,IKNP)LG.U
(T)Q@]JDc4f9,6U;[8P&2fQVSCC:-Y8Z;gI4\G\fA=d9?0cf-GS=A_ZTHT@BC3.E
-.07Lg_VCQ:/Z;&.<X&9D1)?@2AF9&NX=LX6#@cTNNf;eJ0NU5?JdLRGT>Ge58:0
CO-=O_PGM;[UW+(fW;=?+DO7?ML2<aA6c0D<1?>R0L[g&,ZZGPVcZPGZA7887#_O
X+^c+WZTY7E/8?]2-N,1A)FBKd=B1eS_3b[&O>:.:NWI74dZG,[dBJfJS4.L#NQ_
Y-(M85SHI^CL[fVGaQ2^<63V#X:fDPc5D_OBPeLYX/O_4\LDA&@)S0XD,E-JQ]HX
TFFNT-WN)S/#P8;@7[)LP:4N\HY6P\C=PbB1O.>^-?15?FEe<E/#G<V=8&5GF])@
94f-K56@FaUbT8#N\=F,R7CXcGMFE>Ie]V+O2&@77[@R84C-]#>[gP1ae#RaUd,<
a80S;(NP:@NG]Pa/O6KAJUC;C\WBO0PWYSZY/MDaS[YZ@UNQ#3G,P_X7X,6=DYW^
B89/=B_-1Ee)),M-U15/Q=gIXF9bNVAF+[+^:QC)&_Q9H#;^7GXU;;\b>J;:_,6\
\A_SI-PZVbd3NO^OY,078&398RdZSQMDWL52\(I1).#;5Z_;V7V(E[<@_8>+@d,[
f^><Ja3&V0+,KQ#Pff3V.9.=./ENWGY>V=]#_]+)bQe<VdS]BL;&V;:1AM_\52>,
\.XE:DC@(;:4I7<0>A+2Y]3DBF-O_38Se+K;O0X&??12OZ^9,FMKS6DPX65Q-TCL
.d4C_HZY(>8FO#47(&AZO^8Q-+5f\D/[a\B_5eH-PS8UBOK,dC>=Y78&BbW=26NS
E\XVI]S35PF:Ha(C<Ld0^cN3.N7VB+bd?]QA5ZDDTI2gA-V#T<SP3cX],#XV.&e=
[a](S=;A5.N^3<5RM^1.,eg]0J]?9N4)[\VUe_NBBNX^eYH<37>UB,AP5d-RTJ.d
#be9X[Lg4BTT8:IWSO;7:MXMZWX]D-5:R[]g]&<DOUJa(HL?a=>?b^TI&[aICe,Z
^7Gc&_\I>=,4CZU(e^IQ#GAM8-\N9P]8bZAa6WO;3?QKGJ^g^XJO2L6RGKQTBE<&
<dG5LDT><@Xc9[CLB+5[6UY&Uc/QD_3GPS(OVbN+MM1S5\(N6Bf[DBSJ#g5bI?ee
3-<<F0+gWQ#=KFQ.447(JOR7AM6[GA\O(DJ5L9d5R5:TW51E/aJXHUFJZ[.1N(/S
cg>LE:@^6ba_gLAL?R@Lbcc.MdZ3+-5+J/MX-+\FM.=>C3EA1Z->CPdg3]dL-J7T
5JBO6/1eVBPC;YVZYD>AB/=BRP5^\>Y(K&D?/]4SM(BbWe1,LE8IC_Q->#<J:WB,
:]c;NF0-gg9K?C0Y-A\A?UT^Ef6?=>GYGV>71,fBX3C47D&LF-8:#ZPOSJJd28(8
.#E_B5]:3H^H4Qb@HD\0(cX^96X@bX0=)50Y6b@XJ^8(a=N<W:BY5QcBQNTIDEd?
ZSRV110)(,<KbNDPB[cCIE.121feMPBZZKJ]KC@7#,K;L3FO@EP@NJTJJ)69&CS#
FSLQ&PQQd=C>^AZ5,bWP,V-73(BQ]6eX?=CAD=f,G#N+da[UW@D#XO&TB:SX\b:>
NIgGaH9COZI;B76f?]aS>S5>LEP[TbQ:+030O5>Fb^4]a[b._AI>/MD./EDY#.F/
TIZ13I&6Sb_fd=W[aW(@ME)6^eg?KdD+Ua0^9E#g>=^3U&/H,:C.5>;+<aH_AOc+
B8d\,S2H8B-\FO[VeY+O6Z_@e,PVEcWe>d,@d>&38d0_=<6H52Ud6H_fFH;F0]@:
>@YMaOSF&RJ^T)^U@RAO5O6#V-N;3FJ^80-P9^Nd[3QgU6R8)aJ?S&]=(?MbV4Xf
PaN9D74eV1KQeLC&X[:g1g?b]WAXbg,M0)Z0&c_<5#5YH1U35\BFMZdE1RQ0#32;
166+Q:RGQK4+Tge1&<:R;.8HYD];IC#Z\0:R.[Q;W88VB2@dg;JY^;93.L<04W3\
.5MI73X/I=<):(c##:+B72MafK+3(TZ,63Ud&D&G[Z-fT@M<&SFfJTRI7Q-JR>@W
,OW#Tc1N>8BLS9F307M]T]8aD>-R0KTLP]UES\(:WDBeIVCcd_3B67\c#,0O462B
YP=++F-DEf+1OTKEc]Z=[2>MZ?)Y0+<70ADRaIfK.JDYUg;<d9-?;WfF.E>@2QA&
\7XS::1aD(E,=9gYLGLXZZJdCc33(G#Oe.IR.J?Q=?MI1fdT?b#K/>B[B:@4I?d2
A&2H/ScgH9.?dJdQ>@F/AXIQF1BKePWQUQAX;cdSc.0PQ:bFaf,bXY4&Q^LD?G#<
)C1JVgcP#/A7[)FN<V75>[-D1\B9FUCD@LITD=UVI-c?MIPL/c\8EW5UEK.U&8RD
X753S:EG-([64[)MZKETKT<RdC(SC^Ng0MbSB&ef3W2+8#79,(+=);9Xd_0O9>Z>
EYLF?0EH>ZQEb5H7]@S&U8O^f&.0ILP4V<>C5OKI,74dJNH=^c=ZY7M)=Y&]-]@g
D;KK:e730?/X+3dKE:S7[]6&3@<9&PLd,.UIFU(.[)991gJY5P8];LJ+O>=YI(3_
a+g\b?7X2<F5=E)I07A&)]HM24WJ>9:;8GN@F7.aVGW^_#V/_52G<;XbSY/Sg(R5
LcN,f:gSA,EK,\f(D2f47<T;<<15XHOL\+6A([7MP@OW._YDP<1[HbIZ)F5^(>UY
/A-Cd([gP1X/;N=;337,bWN25;cb/^J+d3@dcTE(Y6TPZ9-GFA-29QVT(NH]I]Fg
d=UY0B],>BCA@RBP=EE69/U?E(+&0?#Y_8&?]Tfb?8IZ^F-5VegBG\Qg,0eK_D_B
QWSBb/GfK6@/Z5\1>>ZTbe<E=L\^+aXIf^XaB:C:/NUJ,)[^HdA0N_WI;EEaC<-&
RH]ZM>V0KR&9RfHd7\.e^6&8^?L@eVJ;SRZ=E4f4N@J4cDJ]Y1dRAaDWb&VD8]C^
1RZdCa\WP=2E86Q\?7,@c166#D[dF)-aJS5I-+FaU8Y_8f^L>2-9V@6\W2QAX;H@
KXJHT.;)Q/9:<E(L&a1[Sg?JeR:U,DGe3KP0gA[PHTRQ1c@Ge/a?EeDfd&.M:VE(
])PB8H6Z7&WA:U/9dM;^U69BJVbI=eSa9GK]aI1e]PI_Ff2M@_/UC;R&H0)&bPe5
P3JBI..5HZX/8a@8f5.a=HXT21]-.XDYd0Ibg.C+PZ-aN4)O@=,<K&>13TQQ=>FQ
(M#:AfeX7[-.]9O7g;;HE0BV/b+#LR)=Y1/G:d?f?Y3,ZeFM+g&/aeP_8IM[SEPA
;^MC2D^,<[A:60Id1#e84g4.:fg_K^)_UG@.4FEc5\X@gV<g:7G./.F.eG=g7]=S
Ia@+dCSCL@12O1SbD60;==?<@#Sf4.MZBUgG]L#:JJT+S:[:(D65QdW@cE@D8&S(
_N^HdeBPD.:\,1?cb^(#ASZ?TP^WLC[F;Ea^)(8^aMe8c]AZg-O)GR=C])=P4052
+#f#d,(P#[TMY>g//7]V.YR-.;./_)P.YdZ5N<#L0X@_;XFXNZ@<YHY4E8F<H@U6
,Q)bN&54+:c_VK5:JKAS7/D31[XZ941E?c]P.KY_F6T/11YBE(+EcUX9.U5L;ESa
N(=]1fJEXH+-f5[2L6VM^)[08P^0Z#-C?Rb^8Bf\<-&@dW9(-MS)D?5G<^3dg&,:
[L6&+XQ-LcT02d\:J@24=-RC<B(G;ZL70D+GC+8=6)-],,fTf,:O+TO/84RCO:I6
V57cT_RZZS7C6-4#SFPg6?;H@B)=41f6.eN/,=>X.16\^A;\gY1)IS\O2@9,628Y
Wa9&a.87)YHSKL_18\]gY#H(T\WeB/c-K]U^:49W\b,f[U;Q;XZE?Xc#J#0T?I[#
5H=GU@?XSA[>G)EF:\H:FIL85He+Y-<RIJ5bNaAKaF#D1U0K2T6/d&Y.abA=LK<M
0F746.Q>3[+3F:D0)(D.#]fS5L/T/^Y&0X\X:b/FR,M7fReF/,G7#e59He,)g8I?
S/-F=\X>ITW(ERd2AJWXC]RH4@-UMa._@f;P)D-K]-O]e,CUP0:&3.R=UQ1#SLD5
9Q:M)@R<MX7OMOX9=6c-g]_gb@9T;gfBAUKYYK&:R0_7V\:5=QX-2cc(V/&eZ.\4
d>@5]RWVY>1:G)_U+f91(d#KU?87Z=+,aG/POT(ZG(QbP0(cU_bd4NcGCY+B9T(&
HU#LS/,7U+J6>b(:Ff;a<DEJ8RFP<&L>c#&.,A>G@B&4cEFMP>\Ya24J4cEI6^Na
bg>T#DT2S]?YI]7bT>6XaLW5LfD-OKRIKUA1=K9Ig]X1)PFJ7^Y;&e8:1[:XT)OR
\:SFD/gV;O#^>4IU:T7])\Q3BgQAIB\T8YV;K<V#7[)6-#KE4@b0#f^[FND0P8QI
T.;Z-d]gZ([\M/0E&aP=K+D>,,1<DKW2R24fH54#W4NNJ48>:@GT2Ub9N1C0af7f
cK0I2P:]0WNQR0R.T#.J=0&V+S19/;4dSea5=MD<gLa3H3Y0/3.)]R7X5<@W:06/
YI3&V+NKP#bQ)$
`endprotected
      
`protected
/(][&4S-@_E8/1RNfceL5b1W>Z(@;1f0.N,VS51I63L+3Z]?c&?&/);7/d74#G1>
g.6W+&Y=E^fYbXfF<f0\cYVREP]7[T53:$
`endprotected
      
//vcs_lic_vip_protect
  `protected
.T)]X@R8E5+>eE\GOfgPDK(Waf.#_KC3HZ>Bdf\J7<?P>)0<EV9S0(\b.X[a/A>#
Y0X@(57YOR__@NND<VH4EX?B41U]dBf38U8/3)5d2R167B=Y)R+97X:f_W9P>D</
UD+9VEQ168_H>UY97B<SWJUV=](a-S(1aRTJ<b[@L1^aL(5E7HTOeGEM8B;_17QL
^MFQIM8K\P>[V@)U4#\dEb2f@1fYdJ2\9d2JT&bAY]4f5&a.L&FXG_-O#_OL^:GN
eZf\]0?f(42;UO(;WL]<Q;bV;2&W7>-,U1WAI2E-EH2Z,5^_U07WH_ZbNEH=_bZN
CPL)JR8Nfd4Y;8=#0=,/TD2A2CaQ#B6]1[\Kc:bB4gQ:KG9PZXFWe)A2MVcR0&#S
?@0WRT2V6G12G+L^Gc^:B9[Zb&7:=H^<\L.8@/e\C[L#PZ:<:YGAODZ9ADI/J1<V
E&7NFEXFU2J&7GT].c]XRB8(\FODUg\E00NVaGOL-68TRMZf2(Q=f&eW.N[NLPMf
>Ic/^M)Y5QVZ/HG),B&X\A4&2Z<_&0f38H1+K6Y))Cf,;:2FQ&U?YPaWV)0#AcP;
bT>]1WE1,<^)B,DL#^V?E)7ZIMS<EZ>H/.S/V5Kd)d5eSdV3+U6>X<1R5OBb,RTE
^KC;_,R[8W?,S5fS;N&1GgP@U<5cQ)(2J)/>Wc&HA0&/Y8e;d&6)0M3OZ-K3F)=N
J,_HJ/?Y.E-28_WI@P[cb9I[2Jb/\(\\/+K->P9a2^Q>80&+:aPG^^IC&Wc-NTH[
75?<NG3H\(8g(S:^7>IN(bABJ^LV/_^&=0fST]eZENeF;?(d?=EB7=7bgWVJBHF1
(Uc1V=@@U1B;=F5<6f[(3Q6C(^;GZ/H>U649_&g(LA4;e&<6E?\Q#V16WF+[YO^_
+H4QP+2B:1PeWCHO4PEI_eF77?]Q(J&JU_6Ff3<;&f<bd<#OL=g4Y1Qb)X<W^6<V
Q[0CMLG6,,+XWBA#DH5IVO5IZ\+KBU=Y4+(J>g:V\I.3V4FO)RT]=4);:>I]CRJ+
J3c:R/7_#+UZfb3d]-.dbUNJ[f#,P]L+&2\d+EJ,@RC,\F\W8RU.[=3_?GaMGMZ+
XZfe;2bV:I.G.+LNOBE47gT4;53<bRGZUF;57BZCGPNK&;OMU\I5fWUV/6Q#;<&4
K+D#^f1aDEQ^-4V<)+CQaZC#79M_SZ9KQeF1==<C>^1ffVH_U0W)_E_+;)FaJZ2<
E;<X3K;.bW70ZH\RB86R#^ZPO>a1D1X8(3)PaFG&B:T9PF2/8#M5<>NW5R1US)+5
O#B1[SGdX8(0RNe0:=c]0+1V(,O:VYf<:Qe9NU8F6@NN4/2EC:DBCM0YU&_ed2NJ
?T>RF2B:ME6Q@.VR@dJEH@V?(\:7//#O?79@GDEFMRJ5PZ0b]aNFeYadGO9EF0eS
,(Qe1FT_fPfJ5GW?/-,ZOC&XM=;VN.L2C3Ve]DbZZ/f6ceR\a<Z?)X@8-+Q70e;+
;YR)][)8+MNPKP0cXO]dBc@#A;]_X;3&H089]D:1>)[f=7N\g.;//YMX5\,7W3:c
:0/M6;M0MG0e,?9eMIeF<[;QVd8<_FbCC<^FH.1>Z9T)RN8I\.#_<2IRX9C/c@<B
/Y(eUU##VU+A<:8W^FJFLA4b)^OXGUa^0b/HZKV;NS09N=UU5]4_6_/8Q3HI/N\2
Fbb:5</_@bC?FGM^ECB9d4V/.U:AJ,46+]0XPW4V0^;0)K)gDYD1R&D:(<LERg_Q
AQK&H?]a]Cca.[,+Y(c0>4ae2<WKD)#0f?G2ENYc6Q]Yc.69MJ45B,=5T&DcN6PU
<9#]<8KZL,I4OZ,FH?@N,Qd0<<8a?97HMG-/[KHdL?7)#>9L.&gWI^:Y2#A.fH:1
V:B-@1W?V7<5:5>LH#ENP1^XY2Z#bL+:8LIUZK3.]UA/SQUQ6[AZ;>QO)T8g/;06
=-(M2_M3[M(S12e1AVKB_045,SQI&eg;9&f)/:&<d<KT&MJgC83_cI>Y3/.(W\@G
0b\RK.5FMT);?K\(d]5\YW265+HbGS6S<)\1X3.]1>#[3\>\BPTO<M?,[.NV5H2S
A@c/V25?Sf&S^C,FM9XH:JA.R2;Q=N.@W3eB]JdfJ1a7fRW#<Mg/(,>A(G9a7)Z-
\URRH1M8-W)gM.JY38]Hd+6Ld]VcWbN]d0]RVJZfA^=AcZZHR3?T?f1W4c.T.[;e
f6c56d5Yf;6Y,NG9R24-2D128e_Wf)1,#K#Cc01#?HA)RJa@&O=W40A2fUY#D#aT
48[0<.&F48fDSKE]E#J05D=EGOaA@HK#<X?e99PRO,,+1UPNAbCS)3SJ6G9\b=d+
&@RDYU,RUC?HGKL[39O(KH^-25X2GaH3.I#0\QP5YL(.Sa@WWQ:>fU7WaT;B04>f
cJL7A)K#g??JH[<#Mb(:d>5?FS]?SJZe3PG@J)(7Ga&>Ce,5g7CfBY?RcFWbJET9
.\PW;,VO4/E2b),.[H:=N&C=@BTBTaU6_-d3Eb/N)JZUeJB+gI,&+g>Q=5H-R=b+
)I/MX?E^4ebFVW:V[KSDQVAQc:Q>)P4]_:(Q5?X?e08<8S@9(-O+>c-8^(#IC;5c
H@YYaG5])aO0JIL<6-gF.JQGL0_+[SD9_DaB)7TUO]?fdPD^9Z?b9f6g]#7M#\Te
fcX>\A?D,GeZ?+C/;XQ81E]R.A>X3P?DB89S<IITPLEaS2R;A?/]CS_NYUH0JDU-
EWaT3_N@62RDc1(-fDI/^>HA/=I1A#N5W8UW<7\RIJ.eGWL1PI<5N=/cg(@g^0?e
T?,a#OHa.1/dHgF_ZIYC;#0cYXL[C.Q,bHP4OFV,3@5JgDA]a;[UQe^T6g<4T2+e
4HT))QZF@++>2Z^Q3-TGOb_8EYU=f&S-H.8..)E:N&FO,.LAEQfCQ[cSRU<:b-5I
-[\S@F0_@^;?,Sf0XR&S4b,R]A5NFE)fS/R=2N1@H(,LR_NGL2_=)=[>AI5SI492
BcX.EgIGP-(#09-67KPgA9)b)<YOV5KFgYXcMV]2)UR<(1b.c?gHfa4L:[>SJ@g<
ST6\=JJKP8Q@EcRLdF>HL]DbNCe>V;WdV9U(WBUC/dS,e#(MDHCO,9[U3,;5K]bM
,?\e?=/=,-/P^E]-,7ZDXN:XCd<()0XNW5e;9==#W]^.?-Q2.Hb[fO1NHf9#XEbZ
O-c@>1TC&@S2HV:^+2VG_dR2[2[1+QB.6&-<D,3WX[NT6/<D_XAf5)e84>HZ=>G)
HHNTVUI6@)Za1=d>J0eC;:0;@AJ1gLg0NQ3NO9&ELaNH/,3<MD-F>BL(@NHZCZ06
>7AJaS&;;gaLSIK[?8+[>SAS=1#E=,fUG)^e7M+d,/e-SMRBC4&ID6LU6TC@0BKX
^9b0?-\<,:S=^+LA&[X:+O<,aMQ583Y1@MWQ+KVe9TXZ^aJd(7^Lg=67Ug)f/7;M
+#YU>[OZU(c#-2Z.6#_\dYZITgTfdYNRSTNHP)effdfcB:I9P;<fA1X_O-[;3K0L
Y8K@UW@D@<<;EU]FR>1]YOGEO^2bV&C]?5gcQc2YKY&LGP<f[W545-A&O=[cZM,4
2dG3a^SS6MdXLOGP1-JA\:)ZTc6TJYe.?7+R>#YC.aedE&;I:?&==WNP6QZDGS0c
f>IP55M7ZAI>bSJDA0[daFB>\YEX1OL(=(FRV/W&<-?UI<+,CHZ<D(QOA<gf<+0Q
S_U;bG3J?6+Oc2)(S5^?CeY?REB6MIG^G_]FI4J\W=dULYOgI00A)e?QB-KO8B56
JKgZ2ZOC7(W-=#Sa7=[X[@ATV,<1c#,=\>2X(f9ZJMFEAE=QGL>N^0X-YQ;5S@KR
I#O,+MN\T[@bD]IE)Xee8,efWE3c)&#4Q:QR?99TP1.URB&.77X;E4G@Ba^<5ZMM
_WO=2+e-g199=WY\Z&<5cYTMaGQO]=EJ_/bY,^&)7LC^9;WF/I)QLd-Fb)>+?[9@
>M5dX6=f)a]^MI8&,GO_=I<(Ue<N5WJf.M_O4UHD3g#NBQa;5](0aQ,#Z#R&AA2)
5EAMe:N._Sf#BJF7BN)WaSdV/AN&-cZ;],77e<eI/[5J2JQ:R:,D[.:?[IGAH2PW
&S)2:.HI+A)#@Ld#HET-)GM50(HOF1+f@MDAg).E-V@gQC9J1T2C^+V]KQD^_bCN
<,A95^&&-Q01B6G;X)AM\6fIc5+Z@85f8@EX0f7\eO+e@W_57ONL:D>P?8.<S(Ge
[?PNe[3g:4:RM0Vf^(9L>9W81?H(M)gJ_-1D-HQe,Y+0MaBZQ+X&fCJ6WWNI?4f8
N:a+=?\g+.WKCJ9E<X8X8@7\6g]?>d]0Q+@0NI\Ng[LN@8ZIR4>CS3FWPdC?aVM<
C<2>2AY9FAHdO1NfdB(:dY:e7H<IfD=a_3SGa5V;:2Db:(8#F:c,IbW]N5<7gS=G
OMIFF/1D78N\bA>0A4RG0YL6A(7(F/[b1\[>;2-a8DL.NSba7Yf<f];N?2)c7XH6
&+c,<1\fP2K9(adTKPOGYaHdXF?DRD_&7Ld>2LgcSF6)_c2@2M\C+X?(g[SK_bM3
:4:_@S;<?>I;aLJAPI)eHL7:T2#8943G)3LQ^K^^1\59()DX7R>Cf6(4ATZ^)2bI
EE+HN?M7[fIU<Z\[W_##&[S+MG]&XULa+C#70G/XTKc;GM2eC1;-CFfTeGM]^D8Y
H,C=M.N?RV[\]DUD;0a3cK+YUFJASWU#fe8?OS?G>ed0:_9Q=;9](R8/cR11TQ6,
C/&d8KW:HYBYS(]a6T;gG4Q7T>a8U8#2HHFJCCEC^]3EK+fY9]=R8./QXA>[>QF.
IL\a+\:Q7dC,4-PB^,c<+_&:YcdSdJUTK(;eFOBbAL9e5Tc&[GCT98M/<5afa?-N
JV?ET^0V[PJ+VD?W42PaP4L#WG2]Bf4g8,VC/F\@+TfFbOaJ7MA/aPCSN#.F?^gX
^<18^I4R=^IZ5-#;]Ee1#\gWZ7:H[1d0[JTPE]#<5B15K+^@C6+[^+\Z7Ig)C7V:
I>+E<85;7/Qd3X0g-3E@9M^8<.#Q+CPaR)^2?)8XY9#J+AEVfFUHFJRHg^KS:\#0
NKgN-FE]>WC,ATU.9d=]dU&ZMF]f#6(Ig9BLc0QA0RQKe0OC)c(a9N=,\&;^g385
4gHA4VLgWSZQ#a&4S:&?37\_eGMEX3b4bW0VWaSN&<]1G:OO\+=@^/UUAW&ONVFG
8gA^F1(.YVYFOION3,WU@QG>RAM3f#U&Y;RfJQ^P(bf[,,.J,^3KYXED6Ia+(:dO
+I5_eAZDBc073@<=@_BGUO-eI5DaQLK(W_T6#>R0HcIJ(EdG8[;U@R_PH#FPLMFZ
,fO2aQR]cUF/J[I)6HGE]Q6Pd?JcYN@2H<YY(3@]O--1NXD]4b7<GE0UF=g]G7,^
LS?P^\DL@7+P9fAQ5f-<-AXCJ1FX,3;@SWNA[AK/-H]HF_F;1C8N&V.<40K\.60-
1J6Fe_;I4GcSL4RgL;ba1fY;]8OZSdd.+DeXScFHR1Y9c+<BP:NWaG,/\E]d9G-#
6G,cAZP/;9Z>1??,41K09a0-AL4QA829#Za3MJ^?N)N16+H0-K>R)U1;,9e8O9IW
Ig7W364#5):E<G?DO\Y)--Z&KC[1[XgFRR4LX6?eL#NHGYD(:&O@.3>;8RP&gI@(
E&REHV#Q8[\aT+[Nd/S/Q-YRQA4-0ZYL=YIg/7e&]1>59BF.39>1GOOf4c1fF+ZB
^\b5cSBdKIK9OEFP3BFJK8Rc&7BE@YF\F=e<F)JE5Had-eIV;4)Z58EM6GdJ8M?U
aJX(Y<Y_8F+0S?1:OCGfgWFK8/X70BRIJR2#;VDDAOc?7C+&D9\04Qc:bY#7A\g^
/B5]Xcc.:PTX[+[a]Tc.XDB<)9BE./?D=0UQDG>H4P#TD=0^[X1;QeM+()8WR#@R
fB>FT#G]<d8@@<T79DERF(Z@@AP#)KFE]CS6YF(1a9:8?8/X=HSS]NZESYZ+K1FT
D[aCESdH#DJNO7gEGH1e[O]>\c,#:6<CK0adUK8LO4XgN[V,GIR,#^(PceWH_QU]
acf7M]bS&IJE/EJB//FR58F:<\X)</AOYI<Z^U.f_M,#DI)HM<A=2\E.c7+YI#U-
).(.(/L+BK?]43UBeMfW;;Q&N?J,g)=Geg>[^WWC>==-^eGAR?)L>[6-Z16)N)Z\
E/HeXF9/0^Q)?5dCHf71-a\]I=296U<(&.G&I-0EI:=]8^OM[</1GGfF(L\<.5U2
XHV^beC+;Q?QCeL:1MJF]X-RU8AA,?_62P[+bW0;4O]>5FH,_^/g3&:CDc?^6MU9
aC0RRe0_]dNIAJPSSAO0?Pf]g/[Q]=(3<ERS1Pd76,CO[g;OdAJHIeXI&BSL-3S0
b)>N4;NRDYR)-Y\;O-KcC444RdWQ&S7d=$
`endprotected


`protected
DQ=fT,8,UQFVWJNJ^,bM?HJ6VfDN1,UC7fE5^_]K9X,K>)(U;.Oc3)Ld-?P^Mc0@
6_(R.S/#F?@+@IC^07XC9MW9_V?R#;OOMgI)P_;f/5+a&O9Ofeg/6.<E>8ZE3^5&
($
`endprotected
          
//vcs_lic_vip_protect
  `protected
>[VG<g^1,PbgX?e[CbUU[YCN/GHP2];4)ZQ\VPLd<gFR7)@8>C>=5(g5//baD[R<
f)F[U.+UNf@6T#]5?FXW[P/(e:^HN3YLIPf]1bI0I3@G6@)P5E@g.\Q2dA,F[aRg
QEb8.TL?M,D9_e7ePc5:SMO[a>4AN=I[A.ga??96U@0OKTT,TX64[XdCbdIIK#/L
:ER?a?PU9XR@&M^]EeX:#8K:5=+/[]A6K1WFAC&:Z?88G[_0<=3V.]P.g&)9+&35
cMK60)++0#5RfBa8eY9XO-7>:9)^L0:]J-/-L#Y_\-]&^@JBV5H72TGOC@VG4\M;
,O#We5bUVb1Y+@]M@=7HZQM5SW:6^HV\)PKPUU6W59.M)>5cgKEg9^P+-fIKbID^
+,3<S5UD(>[((=Q2FZY8LO<d5=>a1G3Q-ed]97Dfb[@JX1DgHGN5^5+ba0/MQ/Dd
,)/PEfN0O/,I1#e=A2Pd^g2CCbE0[NcbfBL)SaX+Y[TM=dgKW>.:+gP9H=dBD&:I
K=.f@V6;A+Y+0:<7M\+230[18.O;Z1&WNg8H(3GS(:QWI)QF<^0+,3#[H2&aOBbS
0@)EV)D@;eD<)(/<)^gac8@RI<2GaMK99;a#-1T3KJ3)C?0W^=PV?EKbZV3#QCgZ
cX.dKA3:U]Hb90G6a4fQcKe28e7>5a9K)FWaG8E7Y+IR#5(^O3ZLL,RL^ZO3^e<A
3B0,4;bE]VDW]#M<.-J8^<MA_>G4O[YXJ#VPZUA:QZMS+SD?./+>e#<;dPZGJVT?
:ZV+:00I/TVVGfd?aHJW^QX/.AR]MOU_NED36-<)#-eTgD-[9SCIJ]Z=7HKH9E_Z
NY<BF82-/:8AOPbU>]2&R=:;P?K.CcMGK/AVIBg_#cSeF5C>f>U_:H3YX+34;Z=S
R(a^8YZ,2N((T?L0S0IAUa?7@=;7J3F\cZLdGe=BO2aFV5/FJ6YF+-:+_VOba4H/
@GDeQfa0F]Z8:MCHJ<aSQ,T42/7.\HHO6[-5W80QUW_g:FG2fb6=4X\gcVcQ70GZ
CfV&854\MbV.&c/YQ-f(B)CdQ9T6g#f53@]c0c\UUFfH2]2Lb.HP8#U/MSEJf3S]
Wg\S=<TLXd8JA/9T-+TYC^+)=a0-G,C?d;cE522/gQ5ABKENgR#/Kf;)UK4II:)3
Age,Y@.,0Vfe-(fOAXVLR4C.MDN^D^bS9GHbSVg8,TWGY3SK#)P4;\5)_Q73P,9A
d?RMM1#Ua4a6HZ,T7b.9]3NG/>FUL7a_Q(KWL1K874EPR<9R4GZN<5bBAGgfWQD&
fDW7@b:4daBgAd44g)F@Y>;USKZGIV:-4B/BbWddQ/#d#Y<.E]GHN;SMgfQ4)GFJ
L^P?HXE+X]d:TR?Od\PUP_7W.T)FHOBH&,c-d#ECX22[:BS>=e]75#W[>9X26\83
=78R+T1^>OWR+Q]L3AgbB,778:ddbUF<_cd-NRfaM;G?/Y=3?gVe\aeeMa8(Eb)L
JWI0II-^WNJ9)D3-C<\ZAS/2,@RG/K8E?GUF1WJDKRA.GTC3?Q)[=]ETV:;JAb\+
L??500A5WS9T4(HF(LVMOf1LVB<g(KY&C:,O9a9[<cXY;UGQDe_,L@DHU=96S;MN
e.dZdG_,J<AWg6J:e+YDd-9Y<(BJQD?Q<B0QRXE\;J?N+gHHWAXaeHR/3D[^O;2H
YH=Y@KfU;b?;Jb2B&-_9Z[:5R[.WLIWf9>VVO4KI0aYgc1D-:L\e;(2YC0WMY+WZ
9_ISXMR/d102]M9,.;L/+U,O&+/[QN8:N^W<dYTLIJ.g8>cSLTJ+Za];#&HVXca5
_C65[9XgFT\8^d7.E&O1BKf:K.=#-fN:UY0]+&@(@bG-I-7:8+].S0Z3<JPQR;#@
MWfgIXR+>:<L=3)8\@P@#OVDTHT=W0@@O6SE.f3gW,Z?a3KgLJBJNT-_;d9[E7TA
b7=TRdcXYB13R1QQfT7OGCD4KERU@N60=YF:gc\^9M37AfF^,P7F?G[_^U-Xa0gS
HDTHQJbc&)SB.0I+[X]F@EcdP6K.4<=4N)5O:a<-HQ8?4P<4CV++_.ZG6PZC/6K3
?6+]JfV4VbM?Df4CG+93&YCgbb<aG57\]:8c<6Cf+KMAE6AZQIA8#^-1a3Q&_V9[
O\M]8PKb\bd=K0^Q-EP#A=;CQ0VZ0ST)OZ7<<KLgIRPOQ<:D,?14PWVH;+R?:\c9
4=_3B4]4GQCg:=1^GW3AN8\\[>4^C:<A.4H/POJ::Z+)U),HKeJ>Y\Sd&Zd8]J^Y
gSO)Bc&Z)A:YQTIUGKFfAXAIeVO8c3G(g#RO0&UDQ:J;9GVJ<?^HF(+M46K,eHWG
1T0/RS#;d2J@&1M?#B1cZX:-\E(E7G_47Y^]5D5N2G5),,O6=Z_I8XPfRe]:XFV9
3QFKReEbfOHHg3PRBZe4ALY-QQ@X</4YD9B[LBW;af9fEIVO=faTXdb#MA(Q.bRP
2[8PQMY;.M+gR[?L,W@U_UKbdY<Z1F<)[5UJP..;1,/IN;+70Z=Y91^0SV&3.g73
X_1GG_?f0\EW8McCB5I,>GR^:H6cN1IY?3Ea_XXR#?K7Nad/6EQJM?6E/JZHb+Q\
38Oe0^Y<&PLLZ^+#KGVC16[[DD3#O+Q?TT,OQ=7DN/,#<KgR-=Q,6a2f4S=S(3PO
gVXaOEFfE]3c]S#\SWFYMZU..94N6VB[MPS<.,eLU-V4<8/1QbC6W1?Fdb,L5X>.
4H.KZM^T0=DM9fA9TWVdN6?[]UK;MOF[ZW,9,^R@(I#T5[<BRNKCcN,e\2S&I_H:
9N.#gO:2&g,DbY3U43R8B[OS01f^E<[bdI,IE]Z:@<P)7f;9I7]5^#GDOL<g56f=
G_(4Vd\1HXRW7.B#6GHgg/FE7SH88:RF<6&aPX?GYXP=H@JUO7+F?c&2BU&ZD:2b
VOLI>=5T@FS\L1]A1cKNf/Za,E>,bY52=P]H9T_);W,^9bV(Bd8MQ/#\46I8C7>F
KO2e=FdVTJ\(/a#cO><@P4c#ceI.6<Ca\ZC[>>:L86RJ(N:YA:^90\^?\[AD\-+a
c/)AC_2[L2Oe[aZd3S>LINS^7QHLeLGOQH&#WZ]6+Z;d\F&fH,MJ<W87,+E\5AJB
b92QBA6DPRR^KFRG&=fDgBd9[_T>>-\ZR0FZ4^dDWg-J6#d^<V]O#12W3Nfb]Y8.
94;BNNa?c+SNa5+]_eYF3d)_6M:W_:1XV#@Ec@>^c28d<,\+;BR&377^SX9S0</@
TeMdH-eN3E1cFc#gI@KFWX@KH^5W<SHfK_J7WVUMc)?6ZKcfPD#db,NBW1cgRUH4
@,d0UJ77+HPOL^3+-5^#<>\>).Hb5JMCN6WMEZbf.aH40dJ?G0>Ka#+D/@:Q:]V:
KGQVNa(;+PM,6c)/A&4RE(._g8@I1;1W\PgDUOPCa:U6LcD[SM,)a.&fANL4L\(5
4dVPTWc/]7X+RC(.#M\?Kef6,W]-YIPZ-,8=\WXg/;E9(Y;.=IHNB&G6bU>4-Gd;
HNFO0R2>dg6@I=fbC)MY?57MOR&)_M]508F+:e7XMC.J/@/3c;Oe4MN?I:GNWJHA
QS3,<Y6&D[E6.b-I#c9L./eW#,N_@S5^UXT>2^Y[AW-fd(4D<dE+a5@Q(DZ6V+M]
8b,g&(CIXf+?ZS6gOEbT.RXM@4BI.(LeMUT\\F)B]HBNI;=TUYcM@M/2#CFbH=_,
NTZ766Y-#)Tc0cF>[#832LDZc;]E-LG:2S8D9.GX8+@UId:;#]-JdCEO<C=4:6)\
@<&<KFYUBe)b,LH?G?;^.MMKP#D.DA);7QZ^O5:,d8&)d,7bA(^]#N(37O3_5D6;
e/<<\IE[0V3fVX7LOZ]):]#-RI@d&&(U[>K1JaF5W^&b)_;M2LX5\dZBcY]TBK3B
0QWJKBY>Dd,,X2S_Pc7[edF6IP69<Y&=CV3T:e#1Cd_X6Nec5a6<Nfg1E:N<E)=K
7V]><b#P92&<].J>eF<Qg0d8/[LEY=R?+CTYd52A5B^(\<\R]a,/#aGEUd#9>>dR
f,H\L)7MfB0cNW+L#<HAc)c6=^?,EQ/<gH,UScWQG@Q2)VLN9[70QG2SC9LVC,Xd
BY98<F0B40E<AD2]1KHYNXU8K91/)=:XDLT#De<b\e/ESX7?NCSK,Z).Wb.TXdYE
=aEVeHV_/);Abe-<Pd?gAc<]2MG]9PJL5/7+\\12;EIO/BD;ZJ8#JXcI9->N\GQ;
;MNWZ^&_/fZF[IO.[N86IC\R<MP5DCHc_eI91T>FF/MK-KY-GHMO8:6dVfY1;eG4
;UK2O<<:IMSPRYFA_YaR&@8fG4J_<G<&LCf(-f]U7E<F7]++DE9:2LM/J/P0BT5@
))MP]/C/bcSL[.HA<1fRGW(eAdS#.C&M:+LdZ]UZ<I(@XcS<X:DY:)FOF#S.&]N?
Fc7NIC<_=;JAfM0TW.KYeLO-\#\>65TT;VYZX>4A&ATD_DD5bM_60b[U\4+1\5CT
d8OXWA3O_<8IU6N+)LVbZ:RB5-XG9W\[&S2b7L]QCH]E@J7JZ:0UKJaMYS@aaNI+
MHYaf@W.9\\1+013&]4:G^Y)]P6(>)2.>7W^#\,^T4+&4;;_)+dHRBI>SMK8G@4T
@4J:a<(OV/bbWX\EM95fb6bU5\2Z4\/M.[58T_Ye#Q+OMIKaSdG.KSP+VFUDE69I
Hf7^Z>SQY7JK/eQ@R-ZOR3FAIaG6W^Ha@/M6d6S;,0W#>dRNSUPYNBLe(6BES>6&
XBS]Cfb8XFa0+NZ8Z]XFVZH_IaZ7AU+EaG[V+IDOgaM=GgGB]?B6&:YT^GG6;V=b
4)ZI,dN)]R0WJ&;S:JQTB^.cOZW<81fVC]LQ^UdOgG03,:602[V;=1G]00W\AD3f
;PKF5eg7J/CAfWCRT5J//)>Y3/OFIMgKbC@VPMPbJ.0J#6;Z4T8^@:X;?Of^.JVR
g#TD-5VXBBN=4\NfI<^8/:]+4.Z^#RAE,83+X?NO-]K(=+&8;@.U7(JGRW2]L74Q
)P1ON8+1;XA2KF86YGOTM=@KKMPUD?R=@UM6A-HS?8QJ(C2(CN#1QW@7e3g<EZ97
Y1.U]VSOe:SA8HKa)b=#g)-e1KI)9L2cW,&D]I.(//cR3@HTQG1UPTXQ)f6AgIeV
e_:d-\GggUcbKU^d3Q^A-M6KSIM):B>OBFZdf9[2^\f-TDO91fd1?#5Y3Ib3@0c>
G01,fOILGD\//ea+)e4Nf\WKbOHKPHJH?>f8]/;5XD91b:I=/1OXGO(]1A5;BQ(-
fUaY>;<LW8cHEa\Cf:-c#Sd971cWVN)U(K+QX=DC,B5b_[=RQe5H1Ta7PU;?DLQV
CR1,/baXYZ(cAbGTO+QZ5H0^EY2?W,5=0Q<M/Vfb^X&2Y/gbD.S@YeUb/8-Oa/c/
XVg5J<2/GT&Jb.,0@M[P)V,XE--U.4SOKHe_ITB7LSFb.W(,@U.+2AYf^d-LT5_P
^.U8ca)Q&J&R1-IRQ(<6,A=EA_#B0<UgU_-U\3\_Z91DIJT7_#<&0WEY8J#:c]=G
.&XAa3IBU]@U1AXE(_E#P\OIC@=79D-9W^+cT+@gD/K.HCQVbe?c6EC7A#A(^7:R
g=d3U-HE>PRNL=>HJA6U8T7X+N]9ed\+;OJLF3C#Ve>HM,TN-L#HgfU?X?XF\Q.^
GB12WUDWCWZPIW\cJR)_1<Fe]eaBd:GC+]DQ>;G7..OSLZB2Q@bB=a685Z2MIQY+
b:NVO)(b-gEd@g3#HB+26KG(XVZWdBTIJcZ3?X:eMUR_MTZ,<SGb2G^FfbG4E<0b
ZYY[9)T(G&M;\43G>)OQ&(YA[;R71_9.K68d95#/X#T_SE#2<0+\>,#)b4gaJJ&g
T17C.B7A#9b<1.AgEQ,OBb@DCA?b8Jc1I];c]4,]Zg?56XM@cdF9,7>=MLX[9=F/
RK@5KDR.>ROFS&[L;E+B,V8dSDQI[Xa(5CN5YR#D\SVgd^KcGD^.8ecAc7MXAgTT
PSefg,OLVETB947,a6U>I<JME@.caEN++Q\X0I<&]=97:24]2P_EC2+J/d1Y]K0C
3DQVYFP_(5NNGA]7?GbMc2,Ud_7,US6cg[K&RJWf)GYJB@>=1SLWJ&6_KRFgN1+e
&Q:M@Ua_I6DO:dg0<B02)?N&>JP&LUe]N<&N>2d\;H.=SD]Ub]<N_7dg@3,b0B1R
O(2JI>++32].EG@L]P13KX&aSU85.79<MYH(&7^3B&T,2fHcDWd7BPJW<Z&c\Kg^
AVS2Q^:V&M,\/GIBIQ^fS0LY4HGH&XFK81IFc#9:Vb5IPF>CN--5U2+VID+I0]N#
2^A<1EN\LOTcfL=Le2YM-Y)7/UV[UDM=4GK=EL></A)DZ9FQP/ZC-R[1&b.#,ADX
cN,.6QFA=;0M2d,KaR>G<gQ8?6M]G^3:,;J/-dEP3TFc@bgX]9K90B?5?E73&M5f
?TI31SFDa6Yb&U3f7-GCHaXL7fJ7K]05D<1_Q1DSB9RX-1SR?@a?W0E,-XWIOeRb
BH57FBM&?PZ&:SK?;>A.-=F\e)8F5,]]^gF9.S7+-:BAB6PO?&[P),3ETQ07+d^+
2(:1FEb(];/R<K>;CA#M1O(Z0&T\-@2Y2)ZL1^DC^;fd_O=7>(AORWLOd4NB;2]:
AM-3.I0+^JCdVMN+R&\=I[DTKKJKS#ac/N>N1TY)?X[dC7I/Fg_3a5;RMY1(BB^6
Y;#Z,2LX5X9?;GU5H7S(P[AT_6V8LHce3XV]=RdR8FKZ+2)+D#TMRU7edD>=_#Of
73+f4WO,WY,ML1FL7T).NUE0N?1H74</1FS7\CUEDW<+c&<]ScZ^/#__CBe4a(Ke
3I^XX,b1a0]EQf^V__U600d=S:0d@/>[K^-Ka)DSM&635c_3a4MP:QBGV?ac9@0>
@.;KUXUD[TAPbTM#1]WY&2GGPX(>U=X>f]EQC6TFgG5AK)DaE?E=8W1YbMI40IXC
.V,H9c=EO,eZGc1e&/-9&JTZDT><--cFdV@8:2M:,M@JT+]2Ya:B\B8W,LTNT]>)
Y#&b0GGNA[L_;/LHV:DcaU6-^4+P#JS+UdZL9c)&1fF53=G,U7I79?YRHgXa:E>=
2,2IG4E&)CCYO7F3##3UB2IEd@6L1#\7X8@?X_T,_QS8[aVW>,b3<=S]Y^QZ5T9B
/I;K013E1P&Z-SJ28FJgX]-4,N:CSM<7g#ad@<fb)g6eU^,CW2-9[@^ZV7cMHId^
K4cM/Uec6^L#Eac+gDKY-Yc-;44@?:]J:KG4T,??R,B5<.@FPEU&cc<X[N_a)^Y?
9?a=>7#5&?@-C4eb[TM<d]De@XNS@e4-a+G+):D\@^7e#2<GZf076]e>+EI#X-N8
?]?W^6,-Ace5;DIN4U\a,PGVJ/dRCaC7I2J7VS;^(dM;(#B+)ZCeZ->\F:A-2<Lb
Pd17Hbbf+I3_bEa44CR8bRP];+9[1?UW/1WNc[+F66POF+0PP_,EFPf,Qc&T=:,Q
EV0A7K.CN_eZ,adPDJPC_[MU212FTNgDR(Q&(dEU><,)BV^+P^(:K_T&Xe6Q/)FV
P9CE&T/6E3>dS)bQ=S)99fW\F0eab<78I289Y^0;X(Q_R6MNY2:AK8g=Ub=bg&PW
]]L-7&#5fcI7CdQPQ4VV4QE4(_Ldfb-/,]5fV?0fB/79&HI1W5#8].d<NY9Z:[d7
2U_FSgKgX3B1WUF0+UXK)L5Lf(Q?-^=fG:<g0)K46GO>]H^g-)J-dAf(@BZHOXXa
NWgK8G[aVRJ<(0)&Z[1F9]?^3\VROAX[+cdOd9HY)4C5WJJ4(],F/@2<bFWWY32f
)GLPX-LdW,)3B0P6X#RHO\/e\+QEH]E+[S6fT;TZ81\>@cRT\O(,Ya7<Md=T8/b[
)#<77O-GU>gLgU?b=I-U@D=]H+C<N_1/&>31H8R6IO#0QeL=W&c??+3UEIgAS01D
1XI)Ib<6eE]/3.-ZTf7N_^=295TC.V77J/71^Pb&2.W1;-^/bD,L)[620AL^[Cag
2+68P+54?QBD23(<a@?TBNMLe;G0bbb\bcK]Kb,91WbQD6bC=4P6V[_[C9O.S?L=
&;f]\cE7U2Z_PP>J-X92SC(2P[M68R7@BOW7+CE;:b2APbZ[7+6KOG1WNP]:ba?G
95_U&(5(I5f617Ca39;\-5#MQd9KF=.9?07f@(_NU@<JOPG;[-WWPc/(FC\2DV-J
;4C_.VB4G^ZZU7K,M9ga<]\Oga&ICW7\fg8d?,SH59Ya(68+bMbI44=:CGD<1).G
JS3,aQB&XQ>IW9^1(Y(fI;OCd;X2JcL,T+Z.:)N/_3[gBfFRMFe&[],]WPW5\.M3
EC=D5W(=K/a:H6_7<G1D^RN-.#IM_N\_G(RY?)TQQ#=6JW/F7?14Q/Q2aTM/=:O-
L14gbI[g(1X_C=<O\0;S[8XEFPV2Y;94T[@[_]Q4L::6Z]_OC0+P/(FF]DZ9:97Q
FY8,-;P<J/A\/ga:[d[)4,#/cPU?9=cAb<ZRX>Oc@OZ=0G>D([)])MR7S>:0DK8W
4UJFE<?^I>(8CCc06_#Y/_+.PK6K;)UaO4H;E]f:1?X[J)RE_;32)Q5Ye1X3ga6]
Jg[P0]4Y6P=M,3[W3._G7Qgda6>&U>g>X^JN=a=(cf7,V?F@E#;?(?ACHXIT.SW(
+0GI5A5FOI(-J)N;KWL=#/#TRR4?]5TVA,DD6N(H#FZ3gMfJQW42.SgB)c6PeIWX
XL5EYR),?]C)Ve\VQ^a1_M4#FSE/cH8QeeKH9_dYQ0D7WB,d2DV@fD63XG]3[_>@
NM&BSG-9IS\2fCf>_R\Jcd(+^a^PZ^5=AKJ0=g))+dN6<MV1Q0IBFQ4[8GU^,fH1
1L[LNd,,,fV/R5J&W>2,GB=]36^/>aK)X)b#J7b2U?;Cc=0BB9++799\(8=,/G+Z
cBcU#]K93,gMVZ:eR0RT?V&.X?KK#;IfSeSK4N/MH)X8Kb,&@S#8JH(=O;E+T:,E
]DPRA[;VK3X-.E^VX0C7Zba7)1KYBBK?EQ2.H/04)bC,N2d#@AcVKCW[37MXLeSd
g;7B:H>:eZ76YQS.OdKFFL6#BZAMH5N/J/&S\+a[8<2J]^V9#&#T[9EITY=_13d7
].?AIG+E=-=OEJ^MR-g\8>6R]#C@P4B]C?D&WL^,LUW;Q-57Y)5#2La.\JO/_#\#
7D.F5+4_QEZ4KPN@c+MP3<UZK5&.Ia&2bBb:@CX-O2e>>,:1Ba,SHeC52AAD_dUf
J0(D&d9f0^d1&-O3[X5AN1d4HZLAJ:A68V/ZHFY<3S&A<OgYA&9d]f]^JJg_Sa)L
L5NK@PHH&(I=VV4(C[):\fRH82F:T;A]4XWc)_4#,+a]=DT0_/(I[(U(9Yg&aO@C
SFQO?GX>=V/@#aIgdO;^)aa/,<2EI>J=4I]BL5LCeI7SX>F\g<:LG.3+_UP1A-F=
&R:\&G>XYBdZ2LG+TAbZ&H?L728;)a=>P-^M3WDFNM7cdD_,>RJV2&-]>#+>OVU#
+?+CCb-ORf;HHCFD.66\9?O6@:7^a(:(.81J6EU[U)J3=XZ_;@PDZ^FJ:?R36,TL
bW2^Zd,]Y.JOU1[\3YU.+/.H?S7\]0W[&JPV_#-7@UTbUe5dC+Y]/3-26@GW]Ece
=MfR4;[.24a43b1G>_7G=;FZ>S4GNY8#dEWfVF;#?XLDX&X?+L9&U.O3+6ZE<,C)
ZJ3<:NI#dY01f6d+6/eJFf)+M84;&6I#X-+cag;95\^Tf@8BTe/cQ()f1V84He,C
)?UDLXTa9EZ(2VJ^;EE<3X4#S)Ib,W3\^CV\FZ0a?(6SU:eVb^[C3d#U^PF.NSSB
3Sb9#+3f&D.0+Z:\42EXK8E</d#2G0?&@K4&DAT=&&TCd,N?HB[VER7ag>M/dEH:
AS+b,W1e(gN+fQWW+a54R5XO;gRO:2Q[+U:aJ+QW5-(,1^FfGecT^?.11859S.K-
E4Q2=MDFb6]:(Fc<_U]K4b:4#Q^X06R-<:S2A,\/TSa]IRDgIM.N\?d)#=\W6[.K
5<D]0MSaCX3(XBEJGPfW/#F.2=#UUJMJ-a5],?0DU4P:HQ&<<a_S<R9H6RPXTJ(B
(,Q[DJ.W>JBB8GY\C^MRBP0O(X5/:/YQK,I+^ebC]3JfU1+Hd?UI:@NER<dX?6A&
:0ga((bQ1GR_^U?DWI#YeM#L2SN\@gZ]#0E\7QbZ;S^3c&1@+CR1YBGc.[7ObUG6
XJKg3AWP2/NfOdaO:WZMB.+J^71^U]d_<?3D1VMU:;e09Vc<>:>OT<eGMT_QL=+;
E2\8>(f_^?U&D.eU<P,_PVc3C;b[&.P?75Kb)/^5O41bEL,<Hf@CaA1N/<QgPH>f
1@-YD\;J\KCZRN&7)]Me1_<e60#aYC5WaCTS5Pfd;2#JD.,P1eBXX6FdY#./DOD;
L,))87;<aC/AV>HNIR1fRQPCX]Yaf[D@+\3J&)CK#caJ^f3B&T8+P?&,8cW?#E@_
]C5][UG7(c]3d3I)#Y/@GF]80.Ze<#MQF,B=O,=\PQPNe3PF/dER1/OK&NTe0(CI
g[C:BV(H>cIW&U7d-BH.P4&]bT6JFG3^F2Zg(b;?@#HJ,-7FX<;WG@Lf<2IW,cLV
($
`endprotected
        

`protected
-X^L,U#5d1.WZ)?;#d=&6f0FU/E.K?Y,#L^fXFRQAZ@IQHC,;JJd5)9[TU61+V59
3R@DZgS^F):7.gL7YA1WE<YcdSJ7+?SfNbDN9WJ7LM)6O<.97?Z\E8UWKGHR9\\W
BW1F^8XR/_7a>g[g2I&#I?I2;26F=QS-C#OZZ)4]F.UKIF?MD9V0XB(D;Z2g8KV)
aCJ&;_073JM1HbF8:,Q(9=4D3LE4<-KbP]NUY#62gAI(I&SF0D?<8Y(DJ$
`endprotected
        
//vcs_lic_vip_protect
  `protected
TAg9&@6>FY+=.<VfOcG)<T,-ZBW=U_0O4S]^K[K)),O206fSM;ZN/(Pc9LLB(M8F
1_d^bF[d/8a]S<HOU-F.CBcfGNWA\IDH.TJ[[S[F/#9@1^4L4VBJ;=bXIgH\)g]9
;)-=c4+6Y3)TRAFS)^U95?O#PQLQ<_3IP]:FI&&SJPNQ+QD,RS)QRLIARJbb>V;S
@L[AD+6)C8GX7_/C5+ENNVT7]TcF1I>]@N:J+A/A/M=GF<7P1fNd,=M(AXc57Q9R
>(W_U1]gfZ:8eL?,UgeK3:MWI]@2HfHG#Z0;c(:c60d<;KEcL=]WQ12<.[Y8VOYT
\IQ[Z+^./T@S@:G)LX1[KK5;g>DUVb]T[YQMQXJ+Z=#=X.G=)<2DP.H#5)ANPg;?
ON)EVR2b8,=1QE@H@^Ke\._<7Z>Ga.H@=bWDBd62fZ+OV&)T0T^W<2:URfC,C3QA
GfgYPXJNf.\YOOKCBN(E;07<b9:fI5E5X]=#\4>HgX5LTg]Y(.3U&8DCLgAcQ-H#
PL8F[Id)H@##ZK#KSK4-XZO815,>JTQg3Q;&R\ed4<R9S5+f3WF_WS_FcN+=9S0+
>#f(Q_H0.c-+9EB1H0O+4-A&dRGD(Z>V(]UF;[9)^aSBVIAfg#D[4:YQ469LI#0&
J[;(aFUJ0Z[M\(b,UM.V<A,Ac5c.c#a&fgF89FJ4:ES+RgVDeZ6H7OOEGQYJN2-b
Z<gg.]Agf(MBeB\+K=G]c,-6[>]8@G/@(WWX33<E9L/@e1bPNAD@8+8b8aN[4_L.
6LQ-=-\Q^<0-B]JIG@fOM)f1a<8\[?R=Y-.KbN0SgTKIFH58),)e(7FcE^C9=LRe
N-J.fW:#9?B89K+dECa;aF0LMVVVWY@R6\dDd18KNG.?^#1F5Sg]Q&PF&0FMX1Q?
D&GYBNDeDa.?25;d;UQX][]UH8@)H-8GB6O]be37<F#M>7fO(:U)9I,<S:]LP_Ng
PW7OaPgY;-57Z[Vf&EWa6(b,?^W0D5D,VLad[O7(\F9R553HNcL[0,#CP-X=-+Qd
F8>^[.fe2E\-.BV)G=#<e[U[(VNVK\L_?.4H?f:@2JM.^87#)\\Ue+.</OZVWS)5
5b^>I0=9T;]4K?0JRQPUP2B9]#;C,Y6C]01C#52<LIb&]/U]\@[FKZZ)e2ZP]+ON
BP@S_1Ya#.F.21-UgI3+BQR1X9bE(RQ3MW_WZPe_2)c3842ZLIWKc]fB;:P[fBbW
5;,\P+H.eV3-UQ]W6ec_JT2YA\&.:BQ(]IKU7,Ra]BP+7#KG_BgKVO,<XFc2\Q&M
I,KCD.&9eD??SDW,^T>-X3GKI<f[8[]D0(1R)F1T^f5Ggc]YQ5X3\JE>BAO>8a[K
:P+cJV4^9WL&N^\BAd_,)4gNHER_T7<_?>O1\_K1?1TC=#2I>,fSYGDH5(g6#56=
=_MEW^[bO>CbS1Y=.DMe,+&E3JO-13,X0Fc]Z)La-1,:,)H?gV>g1]>C>5VRW82T
9HUKEe,3)+>b/gG)5ZIS-_42<>)DPP6a>E+6+,XbH\;5J:/P1daU65aJVK/_W\2Z
I,9\(5#Dbfb-]X(,9>eNY_S@TA-N,L<5=N.UL#LaEd;R<&AgN=Q+/:<4&+Ge1cZ#
IGX):121d1NCR01P:9]80S,)/8L:]-[-RK<IR5VQB;2HgdGd(RI,4=V_(2J&\eK=
9>?,fd@VBCVBVJfb<;4R:&:)aT[M3.+#9ZgRfWOH-/DS>+@_Eg=[JaB0a)30JM62
ZdDA21[&d.;+<FPK.fN0(>dZ_,PN/N;e(IJaS\;VIFTI[cRQ#g&O_(R^ea<(BDXM
/\<acT.R>;M?7=XdN@3Y-V(/1(>Q\7aTgKDPa@]>\D1.cYK0ZbK(>[@dTXZgJIb9
OBe;Ia_TN#[&NZaC2WS?@&eI.c)/#IHaB\HDQ)8AbT8V+6ROJBKf4/D,^)3/=?bI
USAA>T+AP1#?c=Nc^NI#)BEWU_1bEHb1FZ8fX/[B]B\f_W5<1461DId<C&/-4;8M
FJ)K1L?9[,E<\&C/[&b^e=Pg6Ef3PC:g-D,59J>9e2FPdM8Da?;e1KMMcN#1I3\A
3Q]VX#-Qc8UGSD^4#>D#\WC^[<YCY^+=(Sa0g&fc<U#12?cX/d4.6Z=A/>C29T92
cbGNW(N/Ac5CG0.FI1QWbCC^bBZ.TG8c;Q2&eM2bNQR5QU@gPB0PP^;Q/]df\/[O
5B19B3bW(Pa@0#3+\Hb@F^Z=5W:A3ec]+G]Y3#\+9>\GYeDN+7AA0Ye<+WZF\.be
I9C0]SbZ&b3:+IABEa]gDCAT]HcFSXJZ:V:O>L73;=548ee]FR1IKVD9Rf]QbgZg
B6U&U_4e();]S/MEUPUD9)e5dT<R/Q)_b=F_4gB@^=fQ#gW6f5;L;C?V2db#<XKV
cG^g3=0/Z1:[4B=13_X[,.KbKP>7&\CB#XaN;8UO6?KY@/#Pb0?\IA2^AQM^<[H@
4M9B(MNY98P[2495E3P\+RW3]\\#]f,2);K#_>3#^3bFaIK&-JD5/136S(>KX4YG
1JB?dWaeW<M:(G&M6e_K)=SBSLG3UV<f@&cF/X^L=ELU-e.g(J5dU#gXG>V:_NP\
5XK]^_)[SFT:_dd]=AJFbD^8EF?9)7PG,2H+Y<6==[+K^B_dJ11+fP=A-c?H3P\9
f=^)B@1K-gb4W&fO4Q6:J^YJ-ICB;\<dcDIXOS/Z[:&R.S,GSSNG(+;CV5]NS\P3
R.6<dN9NS0#a:[T#c@E8(1CQ6?Y<LVA2Sf>LG.[GNE<0(-9K6/&EcH78Y/A>-20B
O&<O)/A)WP\fA/I]H7Q;Fg6HaNVRHVcO_#K>6@^/Qc/]Z0G+4OG,49/NZ8M9cI:5
)SR7+OI2<F8MZe=LJL1Eb(TA;R=E9E)F)I^Ec#O3NUE<0Le7_87YLK&)R:@Rf/f&
D+/1.^R78\0H4L\\:LQ=@3H)-=-U_TD89O,Q&49<>BKV3E(S1\Y&>2K.8N9?()ZA
3YQX4Zf)/=1b4^1G<=.9c@cLMR5PC6T@PR5\L+KT7f6FN(Z5,[<<Y,4@J:EP\:Aa
WAb]eRZ4K<>KM)bQg_VGYEH,Z#:5g@14V3/-00I.P@KcJ1F@gXY]U><\Q.2?c4]<
SNL;5K<+R#_+&V#IODSVW0RM7RXHZ>aE7(S[3]?b&Dd_JVUGZ<b6Ag6=\IEaQ1PD
HOXFB87:K9fS#HY[MV:]F0_:B^/.#@SMWQ7<31^ec1,6-\OVcW29<fE>2EDC##U.
4GOB>E3[&-W>FJY86]3dMKG-IE-KE.MY4&7bSJFKJXZK>gb5:(+I8TKb:-.=?LeP
d_UcVQ>KELG824e\C9WMSQebFQM^Q7f/F/LQdd25d<O?@B[&H.I[/b926@0WS.>g
gC=Nd<Q[?SD12S5?@T=.\75?A1>SJ<4gP-_N=X5G/])N_1TA0Yc)Z_>DA>HCQS,K
WG8EGL0RTN#.;<aPae,fLW7<T^>+\+6.=aeV4LXJWY:K\Vg?E>&KV+Q=72F4G@b9
cK#Y#VW]]TeLdST;7M<IaW8I7gONBJaJ53(MGAa5]<0X),BG@;94]cUO>QDD3.T>
SM2;_dBb]JXg2bL].;@_YME7Ec^V249Y9=T2I+8E=+<59D,_.++b#\ZD9aHNPOR&
a@9Q5U:e_KE/C#K0GBFYcC[>;.A,0a4_,^W8\[5U3YZWJ?H7X#>=V/40KC)e/Ff;
,PaM8JUZ-a5J576G.E_;@.(\MGJY7JE+2<H3UXYcX-bX&4GdP&F5\]#K&Z1=8P7e
T^1QN].K,6><2D(Q\UQfGR@I1]4dc?+ER7fEa2Bacbd#.X_YN.[GVMLJ)2f=,#P/
B<Kf>@H67G/,84&5:IA@BOZaJWCBG<V&^aX<4ZIC#P+GUf/fE4V.GG[-6))NHWS&
JLX,de&\AE>-@aG]JFDYdWa^8K>eO.UAE[2S]6cWCgT#E:fcd;2^TIXb:adBAH/6
W>(B&<GfM:#\9\2A)9aT-^-/QF9e(UZgQ&KHfR(18f&DWW^c8DWF..8gc_:82]:-
63Z2;ST6:=DMO29fW_aDJ+e-_N(_]OR^3<9_1g/^R;P#.C;IS03XEf1/:CIg,K:=
\S#2V/5aKBcWEZ.ZP@^IQ.3VL:BMJ<^]TLgY6\XM/ARY4KfB5KF@5\NZ-V\f]-6H
_Z&06F@WDPa1BT?^/UCI-O_M8SAP^IO/aE+M)d?)IM]GQ]XJ2EP0&BY^:3Zf3fQC
R+TfC-]/@#gEFB.MY8TcUC+<YHD12^GgPYYdA]6UTAECQC2<6J3ZE)R(UeSF^-^<
c@D9)2C64I<<FBVd.Pf>A^2O#,PS9f(UcLPD5@G((B9^5<,MT?a7V/SL-EfT0Ra5
FCc<Y#Ff[?US[UEb])7V;T;/aG&7aH)=.e/I^P/R?<aP4=-@)eL-g83&bJe,?7BT
^.WdNSKbeLH5P;:1)\XgII1:Sg:g.;D>#X_GAY:_<K/TMB]R-#g7[O2C</fNHA(4
7T::(\Q)CR)[4c3^N1H6OH+.DG1KUU]8)0K3(bbZ(<D3UXX#P=^)Vf&X.&[^fE&d
+3LB([<A2-S^Sd:ed#VU8^4/LG^dZ_P.5e+H#,/FU=CJ8&(T-KXF4a(+EQ2)F(9Q
PLYT39e@66aZ8Gd><fdR3/(L&.TUe[fIUF)__L+#dDE>3SEPU;S&6?Hd4:7G+GV9
C)B&OBRdcHO.DU3-4]Ge9QTOA1feeXQC?@B#IEXO@NGaBRL=P^^-4D\V]W[LI_a@
Og=.<4FUQLMBT:#S@,N<\B#c3QL<WK2ObHAF9AgRJ1^X\^<e\Fg8\4?@V=60<f];
Z<WWcY#5<+//[?+/,af3Q(=T3RMH5>4KTb79_^CW/QVdeH_J><S=^C(Q;LD[O28D
BV,[OUX>S(W))gP&,\A4gae1_CEP2-?I[U/6#VIT77L)X_.UG\KRPc0eNA;U/b4N
cTQK+dPN;gUV.FW8B<&^;D<<N)deaQb1285QW[bOg[g;&C_c?[R\H^@.d,6G>f1a
bc6BX3Td3IC>J#PZ=N6Fb:U//V8+S(Z9C)b.J[:C4)@TeC<3-HFG6^O9^B=6U##,
L?3LDTT-#]N9+?U,XG1fCLa89A_+M622L-IFeXS0cC+@S\VS:6WRFaQbYGC&_JNV
N@8KX<U(O=;Aa(W_Z2<dPDa)Mf^(:2X-JOTQ)-_S/4,;e-U]67TSQ\US9>A2d4Q?
e2Mda4&=H2;Raa,BeT6Kf(\[(P_\/YJ5Z(b@V2.=O>/_b]ZLg&eHH/CDG#BA&^@\
DTMbbFDWU_,@[1^TSC#VEH5ZF_\9^AaYf+>O<_D;Y0IOQ>a9b<4fWdb@C,AWI]F0
)5Te1H4b4Xg;ZXCEM5DDeb02?1aL=>T,9R^cBFO.,B+LL,].Fg0-aL)WVY)[;X_^
?e8e@17CC48Vd+]UC\>=fH>D<ED.X3g4Zd.,cE2DP@(OaddYdMbUB2?a79<DWK<=
0XfBaV[4U?+7D&M+<U<?G^L9g=\:HB=\]/9>;Cd-g=]d+XNKg;Of,T1.9EUSdgA,
#;BW_VIP7,G@#X(X/.OZ)C)UNZ-]>>U<#XO.VaW-d-c/7N^=6Q-3<CZEX4E)<0W]
[5E=4Cb2V5YZLDe@T-E-\Y)C;f@Qf>/bR7(4D4fVc2];&4RU8[Q;SP+HYf=<7c_I
M)1B0EGDF[d_[B(2/CG;G.[896>6DE=e64F61DL/KFL^]0#b4QdQ0DdN+?NJ-CJH
^43R-D9c2A^gX@0MB^QE[]YQPf0\-+d#S6X:/Q^UJTX>?Y(Q]()F&<Q4c[.;I>PO
@]8b&O7P.F@I/d8+1If-]5-[I<^OAE^eD:X9-g-AU)):Y[Q)N>G5()ecLU64=M70
R^>UGMOCZZ+02:83)YdMCGNZ\1_3O;a6S1?I+ODGIKK.(c>IQ@0BD;<NgR/X4fGT
PUI27(<cbMG7_C@fX(=Q]XX+3GWMT780gN392e/+_1I(_AHHTY;.W@T60cN]EW);
>+,,>eQQ1WLPQ,KE38Mc#-faH0TM5\FFAYc@6VL/g>eDcd]KX@e5)3M4c\&JKQ,0
B8XcYJc(=AfA)fUNGI.T\beRWEQGB>\NZN:Hf:CJK/WeN=(aeC<>8@)WLUB1,SZ[
b1R\fM?9]@7>-FU_ffT,c+K1Q/DO7LR8GC+1OY<=CK@f3c24@G.&3QaU1W:AR\.f
fcR=:#E#[OLQb(EW0He3#N9#SZW3?/)Tg;<]HAQ3M)3T5BX6.TK53/H/,eZGWEZ3
\b@739eH)#4gbZV7f>LV.-BF_?Xd/g7.Bae<C>LIQYF=);T+NH_&BPWJ<3Q+5-V&
\BI+ObQVW;D1CY,8P1aWdM,9IBG1E5Z>42[BE:/2O=;Z[KQ56Rc<Va24-bINO>W9
Y7V[HY/#=HHgHc[YJ,S5dI79S^eA:aTG3JPO4M64cLAPOF(0-&149&)-.2gT5==1
,6OX0@KHXY3RRfL(X#]O9,d,@dFL:D9eH;>Pf)f\4&>U)C:UI-_KD9aeZG\[IZB.
2TJ-X7_a>)d#P;6aLcO8Q9NE7,_YO0fg-49)+14;C5[C0DP_GN)^=@4Z)Me,TGDA
UQ;2d2(I/JR]4P^]aHE=J2Se=T#[LH:)W]^X-3E^Y_eF31ZAeP_,1?,J48Z/\HJS
L)^@4(/,.a4LL<;T)XZ1g))df:Z[2;]24K-=/d=FA:c@-3OJXBdT??^S1d7J/;ZR
6,YE>D<MJJBI.,R9P\UX(ga#Zg]UGFgd.57>T]/4^@+.G8WFa8)e/=GcO2&FI3ZO
8N^ZbGCMgWM426VE>&&RFacT5B?PNVP4MN2E<HLGEI-1GC)PW_E<?=?f].8@A<&J
[J7(:QK0\N7Y+S157-+T227MCZbaSX2565&)W^E>Ge](FF]QUAg5NG1f>FRWUP-5
ec9:RCYICFEMAR[aPd[a0Z4UM\[fOc(PA:#>L=;I0Jd&V)XVS\^N<@7AQ,,4Y[+J
g;,6=7>9\8VD>I0]]]=0UYJLb2#59c=<N5#D4M8?)R;\Mb62H(M0&UO>T)MMK.#T
Z7XI_SLE[SV(FgM1JL;RcD^5LZ&I.@O+XgcF_G9:[c-S:]YY/bX5A&>#,^9[Sg67
f]-;MaS=g=6XA>Se5SVd6CUTE(U\_)bB&YY0E<Y.])3]7VNU7.,6J&#6X?UAZM]a
eTfS=XOeG=Y,>[/E\6@)Zf73X^]\<G6_S7+_]a,.=6=dD=++A466_CcfJFREP:,4
?]@3gaY(,TB(=-PQ9H<UB2IY8_7@I_G?5^X.SMTLR\9+HR.fX#IUI>C+eS;8-0<C
b+OG<5@4C(W/_;?-2=@T+9e55I(aT)/0768cZ8(YX;TZ[cFcfLe&C+68eU>C(=R=
@@;]<9aTBGHL/1:HO)T<&)5fSd-[W>S=Df:U,_,:+.\\>,E(OFJY]N_1..:4A#OG
&(2a/Y;cLV24;I9&=[R=7T?aS?K166R6gX<1Ff,1[7PX\@]NT?[-5OW-__W+7D.D
TTK(G8A:2P(09Vc<A\FM8abEP;L;GVMP^PYcDdS+_a_M^8OI=8LQJQN@6LR35S2>
[LL50\C+LVZ?VLQ))D0VQ,J)PUBJC?UQW8AJ(OaDH<PHg#&a-8T#V:4&BC=QFb3W
T:PWYYCb,EG<_I3AfdgKGO>;VJ+GC[E#d,=Ra:]Ea;]-+Q26_\fF)E&?b78Z83(R
BI]3(2c=e]C/DH@?JF#@:C:;G4HAag##16VQN+b>M8352WF4f])GDY1?2&[[Z<()
)9T\\)L4C-T4M]:6FEJQ8DI^2WCA&AL<,\(EBET>L1aY4.gcV@@M-0L8NaV=1KNJ
\4Q>(AP7aKcR\3B,/PC69GC\RBPOSD+bb&&cL@=6I[TY/;SdAQ]3UbSbLF@0,?T4
BbW@,=SJY^RWd-[_8G&2;_2692^OGT>(UZc:ATdQ6F]6N,41aec6E3P02e\\MYT;
>UB)CEP0JGYHTNeZ^;bYBJYVH+B=@cPRae[f[#9(,VB2/c71@21U?P]D5SBSOgN8
OORGD/161G.Z[GZ>#(]OadPGZU0Q]_(X-gRO_]=;-W4]J5EV41V]P&ER7.OWSbed
.<DLVIY7f\AO0T]3(:S#Y+Ba<1cb,O4&[:#d,T8PTa6Cd:8H4A/L220dXUFG=C>\
1gQ^#d.Y0.dE11UeEY/Y>f9e\9(9cGg.^b3d?9QLNATF]WPB3=-7K39J9^0UM,CH
Q#GU;>U/T,AF8<Qe#=X3MZ,9Q48PAFA&d30PH[EC[?N\_KFdWK^0DWZ@3X)6MAEA
]9\(H]<]5AfV35U0f62-Wf6W110E9>Z<RAa\RWYCA=+J1/1e,;LaTSWe2SUHCHWA
Fg\;5DZa):LT>O5Q>#<dHS3DC)T7_)781b]3ge&g4,#<Ig4KaJ)ICCfD&S3,/R-/
2(5-DZ;Z5QD4a,&fP>VWCM=aeBCK@G@G<DDKS&(7SdG>QeB&E(>,c?Qc0O>76ZdJ
V9HD?(:BfE?8.:f^Zfa]OU+aHK=_a<G[?L._5g3<YX;Qd7QC/>XTU+<g75a#B2GG
00Z7Gd9<3MedQ.O@bMP?[T;4MN4@A=PBacH)MKS)0?eR#@Vf-I=e.ae(/F3YATfC
WS3UAPeKF0gbHAIK\3\=PN1W)ZN/C+ZcCUJ&\[B4UgHSV[/U(QNf?gC>:F63R:gJ
N9#XVb50VdZHD@Xbd&ONa1a?[9^\T6?TD6Of94?5&=Be7J(.7DBgd9_UY8UZZd)4
C_[GQE6=2Q2T9)6(?\Jd4F080Yfb6O_@fAR:;O[PV9Q5da+6Y:37]O:Y;FE=DQ#G
O+2@<B=9g2TFUGEIG559E/[]47OM:HOM,[/[X:;NZ39&;P[[BT\M.A?0^G#GIA#N
H[8ZXa9.AR/TCGH11:g]7>@FFb48S\Z:ALabFAe6G/ZC9T3FLD#ENYOF#3CHXMP^
]da8?\O_N>S8BZ2G<aT:HbSR;\Q\Df</5J?-.+#ORZ+&U#_.c0B\_Jg0S[a[-&.S
GJcFQ,@eQY2\]gOdXg28([7gfK5fAF,A7S1[S1cR?@P8B6A=<2FD@B_282)^]5VH
@AVa?_=:92L=,g@^+SG:=<Q&:UU2=DK=TT2:BE;bTGL9ge-WL\,PeH+>L)4GGX0@
?5^5bN.6bLQe.<Yd6N:gR\MNf=+1Y1WC9b32feNNe)QB1PJ)4AA7._)<f0QaBPX]
(29f;Z4C?RWD[]&Wb6fQ@#EI;L_BYNd/V12G^_6Hf,bccgD(,,JG^eBP\V+W<1#c
+\DY6T@JAb_1XF#/4@OFc/WL_?bJYW+5C>(d,8JBYBBb^DKJW_/R(MU..,4+KPaD
JS6;9MfO#NTT#TNKP;f30(/5A4L\^\(J46#A<M(NU#TDEB_[YAITK.V;0[T</)S]
3@5BW2AQG+^)H7;3HDM?CPYJ7DWSI+;T+<?-;DFaA)_bWg#8CWC1E^R=2^fNc=<U
;RL2Z7>4/BTBN:[XOd[@.f+8=g8Ic5.2X@/?4\+-:@QI&@BGSNL@[.]43TM-97<S
FZ3SOE1)7OCgbg:.>@ZUY=5-M3+S42D/K=6aZ&/]G[5DKW&&VQb;,JFP;(CBXU?R
LI-Qf,^PJ.Y:&f@Ndd20/<7e@TdJ=f7<YL+JR@/Ee#@(=9+Ee[Cg,DEJJcdNEX#M
+eD/2=8<EQTYDaeM&HYTdO((9:9_fTQEU#=5)1VWREWAR]?D,[,795@Rf:aL?MR&
_)J^Y6FEcdQ&&:W=J<=TDMPB6eK5O\/XXCFf3Uc.3-2;PH#d0e+#CfH31<X,Q(@0
P.-:L&LX57Uc2CdaMZ>UU8JfVSBG#S/3e,2_^U6\Q2G+E6e1][gdGdU>,4BW=2@X
S;F4cK)CU31I4=S^6A/bXIDe9Z8-U/#a1_eEMcT(7URS+e8VWJ(83P_IWG4RHcbY
KIN2+SN_d<c5HGOYH(.^TLBVZ]Q_f-;K(3Pd=IW@LP9L\=\UB;H\6#5J3P.B22e6
>976A)]/-T=MdXPc#Z=EbAX2bZM2=IQ)3)^4.O2W:Z96S_Rf6ITEH5aFRYU^Fc_)
RHQE.,0aMQ.^_7H6LRCZbC[/-^@[_+IM_GcL7YS<UY1c;dRNGHU#V#f9HSNFPWX:
39Y2d<?KNEGE&P0c,28f<EUPc6>RJaW2/.A5B2f5Ba>a#<-M544OS&-ARYWbX:Fa
&J;gV,N-J-=;-CO?25C>-KL5ST6&),QQ7D6DN.?P=Ac1a)D1>fX(0T82=_KODP[f
P\E&[+>1?ZW?<9_)Z?&-6I8-8XU=071Z_71G#FO1-O0&-(HNQSd=cT3\dTI))5>=
->BL>bR0@IFWNV^AEJC6a)BV^1.36d,BI=1SGUPTR^<Q2&YHFQeG<QgUB9/;JB9S
N8\P;Y1e-\U:I5@Wf[<M2KE<?Db56g?>K>V1MV_FDAJSD<0&U,OQ97N_=@JG;_@M
+;1c\1R)c]FV:8IICOW>fSeMS>af)ZS2S29c,PH#4G9]96HPM29K4d3J_<PN+9.R
,)Ta@,-8HYFE/(2RS&JNMg^V1E]\EfA(0@#]B;[#LX4I(FTca<YEB^?)9<B[^8W]
OUE/.+bBN>&GP^W2^F5A1Adf04#\NXd+&N<Ja(WT3T;U/.##EV(6cWNY1:V=-YY6
&0dHE-S,LBFJNGO5d74H:6d(O:5Abc4KKaEf)g]^f)CcGG1MN;11R\G.>g3RF^GA
UMb83+TP?XL3UFLf-<aA,,Y:KAP(ce\AVRHE;MKHbHVN8R6P993FIZ<c-ZNQWPEE
2SH:1+H_,-N+#:92d\eQM]2AX+V;UE:37A:N\T-,1AI)QNMe8&H\7_?HeHK<C#8)
>GN[.MO/&gJN_d&d&>VECU(#L&38Td1QV@Fd0fNRC7A\V<Y8.d0CdZ\4;N\.cD2W
9<NST^2;>?(FQ4BG?F@B_.FfLgC2D75>0XdJM:/@B0YIR3K=>-JS/BQ5]51bc3b[
R&YC(<_S=I/XW7G[AEc4T;I90L+&1[?gI2:.;@KbW;H\2;)M9HM,G=cAY,<MVXeS
@O\KfO(T>IG]GS2,bFKIOD)].2XeOBMB9RQOPC>Bc;BBWPZ+RGD9?GQfVJfC&&1K
D[(+e[#C:O3a6/J>R?H(/BPRVQ[^&MEYY;UYHC_;L5#9YZA1R2W)=]6YfXY;HH/<
(<NEBAHT2T?^+Q)f8_gTgU@^-#@[SWe(T;O4;NLF>]6405AE8WQRTUUGQdg&G-6H
2X(&9]&SH(INYW#RI4.0(#fMB0_W<d\XG3b]O^M[C=XTg;S#6abDK@8)]PdSF[/_
Zf>;N0#+M(]K.c]0+L983^f=1R09JU-RL46e3:#P&2,,NFOdO2IFEeWa7@JBf(S\
@FReW)U_YHPJ,=S)JX&]U3LFH9D_a:^fNN.1:d?@VG-;VMaMBYV-g4^J&U2K_AgE
J6b;3@YKfVdfP5B4A[aVHL(FRLa\3]gd02=<7\]1_P.&d@S>\H:8g_:1121)K2;B
dCKRS7>,X)_a@a9LEeC4GR)LS9PY0D>QL[O64235g]5OJd@=:GU_O7;)L4e?#9g&
g&YJP(IJ@(dEbAJDSP_B81B:N>f_ABeBISMYT7R^?KC(&.Q\C__YY#[&/]#27#-G
:L.L5K-Y9e[0]#)R&e6aMYW/@5/K^,J713,7g:dY]:PO(56KT<;CZ+H6V<bf<+a=
4M4FO;231VJNbWJW-Q4&K28AVdM/QJ.#=4LafcB@-H#BT.HJZ:Z@H6.K_OIUXb^+
Y))3A7]IO&fc\b]B4N6U.&I=FVV4RTcbOc^]7]GSJ9[+9gd+ZYKVKM(MMU].EgB(
Z7)#fG=O>Q2M9A/egKX<8R1HRFNA\5K,71V.;;1fX[H@C#1dP#-B36C8;217<[5\
X/11?]QRV[JU2S7eHHHOfUf:/J=+^6(E/_Gg/UbB2X?()N8L)UaO2&1Z<_7M8KIa
88b9.C)G1R\c8G(TQELXQ@D1)^0H4?,2<I?8eQCYGfS9Z1H<K=KQ8X@]7#,/)E,N
^B[8GS1a8SF1O2\^P)R#D^.f3E5]\IIZH>KE3eOS[f>V0J]I\]MZ/c_ae?)+Kg;^
5K_R.\Xd</c3gZ=347cW\1#Lc:O;[/g770J;HLE5(LVdfJW^,+,[We(>=6RD:7cW
TU51L:<X;8e4MGSN:8P?8D&gJ7.0\T#-0=WRdQAYV@_2-933-XHL1cK\HM\-=+Y-
][0Y3;f;(e61RW8=5#_7_RXY)+9]HV^^[.93+)C[^>?-V?.b/.E^9/H5BZ29[6g(
3SY\I[H.M34[L@+:MSV3[\>7+58IC89fY:HH5^F_g4S^2HOcN&KZ+3CS@^5gB2g3
:V]DeU,:#&@RWUeCcHB\1=/6+K:e<2KVR^]+baXcNd(.QO2P1e&X1EX.^R@)-TY5
KW=9W,,E+BKZR.fQa<<-0B;H<_JAM5Y)CI0Q9WTSM_=U&UW28<f2]&X&b-AO/6Ra
a9FDe\I]EMYX.QI)8E.a(D@\A,Ze1UH.MND3c3>W,<HUZ<Z^K7B4O/g,:I][cd]=
+YF2FNR,G.K9@2Z]WR+45^D:26S73EMQ-?BQd#\^ZcgM(]f2a?0WWVI:aJfQ,64@
JGEZ1-H-/F]F2M5TY3aQ3QPS1fOQBK.cF/WQ@[YHC@&deK4R<SA.-))N(H4,HK#Q
WB4KU8OJ]UYgD6&^gfV<9=W?OCXc3;AbW--P7CNZO9<_d0OeV?bT,SWfXQ:cN78=
[fP_3+>09N:XV3CT9J6(4g]>f,06^+X4A&FLX_E4JQb<<OA(;NCgdMeO]fbV2a3<
#eMd,DW#=/C@)+EJBYT9U18_HAeG@<QV)^AAID;.TMb9=8KBGV4^CKg<aRO#\<O=
Y2:+4/g=]O2YM<L:5//N^WT:,eS&gSNOH[9RF+1\<GC=cRaBOXK<-BV^0#T[26VD
BRBV)N\fS9R-,[O-T=#fTObE&baFE?U[+>0B1SI[H9<@88^#b,\/8#5NSEY+0M.[
-87Y_BUA/g0KdYf<XWWK8a-A.4?U6cFM_7?deX;@?><0:)MMdCfQK#&2RdXU]eE6
(LEJR01[a<>d8#8=L9)_4.E9>LUf,;,QR[6?bbV\)\:=\28?]ZMJM0QWL^G,4K&[
BYWWdbZ7RKW]WFK@H;1ee>>WH698P==R5VeS3&7d-K<_HEL90YO-X9^b=D&=Jd25
20g0M1P6J^G2TR>LUV2\>-YeJHXH:5.)<SN/2)-^P)=b9WPdU-65Q+F(KP1=P6(J
^BOY;._F+Fg@?P&T^Q/Lc&VB1K/F)5_,=DMT9D?(WEfeXPX-F<./aXLXfD;,03:[
FcW(c>(?]I[/-QS/f;/CK<3B);PC41D-c0E>+@GA,H^1V1S@Q8.M,F]&YL^Z2J?H
O,RP]\R6.ZLg@f,_::aF9&Pc&N]/]OdW+0<MWFKDO]51P=EP36X.55.FSD,G7V<g
^MY^,3AW?/?TTeX(8cUB6-JV5<Z7JFTUdM;[K\C/,#]8_0D-03J,aC&\KE^3[;K]
VdCDT7?&86U.^W;@0-IOH\AP#a7U56/ddJ=7;?eM@_I=R;?S:)NY,Z0TA]H5<bGH
CaQF]E_0@4_?ICMYE2>JN8AKgO5U5TJM&c+_UJFg[,;KF.K6+aI5O7fF\4JE?[e@
J@@:=^-ffIKc.6AOA#RMTYE;M8>3#K<g&HIK(M:_dNT.8c5#Zc\a<^9MXVIW)e):
FVX9L>4eSfCBceRR_cG7)Z(2Yf07b1]XI8gK81-^;aOYJ:JJ:HGJ4_N6_?V^E(YJ
169J?JP@M.,SQZF7MRG(8VWDg1?H]8;F(@(OBaF&VAgN_DDL3f8O)AGFI@2cBM=O
C==X_4bDSdJDA:8&_G9T@DfM+X?7AN7Cf+c88)9ff[B\7IHR[H:7M/PD<Y59AOe8
15ST9db5\\MXG;;0R0JeC;2^PA708MINJc5LC/c/6+#IRf_=R0(a-_)Ug+JLUVT2
KG)C-8+M]J1&H\2Z,2M?GWbc2(EB_Hb+H,7eQDSB:3Yf?T2U2HF_-.O-80#EMg4E
.C]PU9JAH.Bb8MTS=R4@e+@=gPB^^f[0^C_ZF\W2e?BA/TLG@@Q4-X8A10V.1I1,
K,9gUgT&#E-#ZJN4>5gZBGBV#V5RM]_D6=>J5R8BJ5ZY+c;U9J;N6KZ0?+8b/X/1
RC\PDVgb/cQ(=)?QRZ4/b>[N\dL(&ggO(1UdC4+B];,I,MG:<,c;./MgQ8g<\033
(.-VKbe_7&Ra#aB;I8>E5e(+cK+B4)C+F.27)QcbG9MF8NZJ(7Z=GOO3^7IHB1S&
ZV:gX12,Y>2;DY9C)G5>MWBPf,-dcF@A-2:EbNfL:VGPSO_:C_MIKU,W/[<1YR@Y
NILb[E8RbW0:6[KUH(YKXZcH7NG[=P[-,XbQ6SI2R00I>dV7IHKeEYY(QW@eH]@=
<@0[459NIT4+Zd\H9=DL<(0[X/I)SfUZTeOG4F04,N=]^7FQ3Z6<@fbO3T>,K(@d
B;f9IeZ0AP^<RN8I^4:X=(HR+1&dHU+<&]8D40)RM-BA\##94N3^#6NP_CE&0Red
P3,N5O4-,g01c3-eIHTR.3.0;+W/PRXe67-2/L55=/[-;2@O1+db0#H#BHB&>Y/Y
@8>BJQG\Q6Z?eQ;2GP_abFI(#HR55We408E9=PL@=Ye=Eg4QCF9J.c@;+Z>_>[F+
D2IK10?Ca6#63VA2dR:gcZ=TIZf#9ITV&)EfGAMbYIL9(1#b<[>VSVG5D?B?/T?#
U/#:1f4Q\:8<0]5W+QeKJ]I@.K.WX>;JJfM0U1GM/^AIc-SKIC;Q(?2&fZ2_M,2,
H#3G[5^SN2ZGXNEA&#2,a3N#f3DPB(3O[BQ6-Jg[eQ4/99DQI:Wag5LQ\1N)5e]d
:;d;I^7/DA0Kg.2P;G0_cO7>XcLC)(=VF11RcBJ4^gM5C2E3YS3OJ44JX_<XW4YI
9,&1,IG,]H=K&0E7GgG;SMW[+V-Q+T5>M^DWXE[5K0f4EDaeTOH3F&AdYXK63;;a
6Hf0=:VP0<C-b)ZIE=#JO4C=-g[AD7fJeA6aOKd\ZfYZVJX2c=Q8agaV/+d,+cdF
)8a6Z,^(fF8A:?GJYCN-^7?)YIg,)J];c=+,S/4J(<.#MX\cS#PUfSSRHMgQ.1I/
?O4<NG6J6C,H1/=QC;8/0<K:3:Q+V+GPg:>\d_1de)EN,ANPZ<A62;&=2a,cI4.1
g<XGE6ME#,OLT+d?M9-2Hc[,51.a329\QM#g):]/#5T()]1P.S@MG+0G+3?#WJg6
([;#bW:dE4[H+9<_d<T=A,G=NZ;c)\87DIE/@F97+d\g]Q6,LMgXK007\2(K]N[D
F?9(Q.RRPRSI5L?Z</1ZUVMRN63c]]G3>G1@>-6]gOg,X2fE<UEH1)0T-@7)K^B2
=\FG)YU2[RgY.SM(b\&b_7&M^c1W;_Z+OcWW+8Id=<UegU/9(+H2J?>[_E/EfAbZ
?D&X)KD7ecE1DF7MV;gV\4Y&Kfg,8N(=F;6H4g/:3;3GOdI)4#7\J5@+//XR)J_<
&.Jc)Q(c:XV/9/Z?SNDUIc-9D>&T/(L:U;S&g_aA.B/ET<<^80MZ,6Z7+S(1XBaL
MT)9L)+7T)O\+R-GP.=XL8+M4gW1<U4X5D]dG)@SZ,[S7cES+B(=SE6SFK[,?6I+
MGFeM0YL06HZEA2TY2\5D3<3N#^GFS@;+@DOSKSc75d]F-ZfJ+)[8P^CN0VYS8a[
SVFZL:X[49N]JOA.V]^>C18Y4KB]bg78D]Z(7TB3UZ.<5__CJJ52570=3EU).^Se
R))9T]BT>>;)-5S?B/cg;(;?O&<DXHQU,8;.STF(g\]AOL:I?TbRO^5?SV1]6WQH
N5-9C4e2D3D5F7>-dCgEIg9AP^GVISa=gf7JVOc-SJ,>0Dd5/K+0LPFNMad9QG0)
4eGe^8.N4Z6DRV)>/,MKE0X:/CS0W9M<,@/KQ1PIX7>L(L@PY5ZG@?c2EIO1M\2e
fYXM.#D^X.J(3,S&#@T;d>(W?Sd+4f/cD>+2AW(b.bEXN=ML4=BD.QV&Gc1AJHW<
Fg-LeKS:P.f3<^E]40,QP:I,#)Seg3UXG,NC[)3Ja/Fb=[+?<RI4)5eGHcSQI<fQ
RS]d9)K^U-GNgC;N1WVR7_+ggV\bBPa(?)F9G/FeGU08EZ5d>cD50@N#93NBYUeH
W5\J[X]W;EdXe5NB9>Z&HUeH@9a9;AN528_Q]DK=J=GX]0\5A4gA5<<U-4KC1U[b
;bZbfL^9H529Z(@374>ZKZaFcW/I@;ORQHQ@IJ^6QMRSegTD>,[E,6VHEH]U=S-,
P7aK&H7PW2\2LU.;?fSDb8g4Z51ZN0#IQT[]=R0R@GPI_01=1C,CK7):f1#R@YIg
&^CZ+>Tb>Ug[R-,g<ETW\=+&XAQdcdW0SC^\H0^FW[P]W0\FeM-,Jb90HR3\a\^#
ASd8F]XD8V=L:;DD<XR0JaPZB[Tb6;13=V)-H+COb>H&_Kbbdc2BB5\Z<?ML&EYa
ZW@HJg6+SCaU4aB<gWKQO:@/(7KC_c(,D5HHZO/J.7N+M>=P\@d]+J-#4,O9JP46
(f2BaJ2M5IIU_c\gId63-.FFE,UK^bS\M,aO1U;6^9.B(]_agM#f6a\&YNLbKHUI
-c[;0XL1/\f>87GLfP<-U>)T7[(eW-]_WH0:NF(bGIE97Y[eD)9=4f]35CZc&8bP
V3\#-+?/=/db/OY#fL8@,cd9bGK4f<eYEfGL7aH3g0ZL2HH;^61^D;URb/b1H8Jd
4f;E9?;NbcNURFKa)AC_4;BcW.):=/7gLWaRg=K:bCM(g8AF)Qc>Mb\B6>d4c#W/
@Xd]@6<+NS^9>W6cU9;FPaM8CZ(_+@HCX^M/OFC:#GS#4^YLF[B?&dXTM64F>_+)
PQb,.JA)A5#(e8\afbYa1YQ)CYIU^2_90Mfc.RAA(S6OR8LHMIB\=-AF2?)TJ#.c
9_>84>5eY,PNa8V4PXbG=&TNHg_8V8IbVME0QSZ46-B)EP;D<JIHP#2<E/#5>6H/
)HS3(M>BMV_L)7K[?++6P];=8bVf>&1Pg5X[6NK3HX?D0DB2<:YD&/1<;A.-b6,;
/PX2^D=PMU(<HfCC_6G?ID/fOCF:H.5;^7,N8fA1K\E7:fJf6g_c2(N#&6O[b4VQ
8Y3=d_+f<LA61+#B.2PC_Qd=;XS0d4<[ZBBQN4c.@ZX<fDNQUU[<gb#(\;/R&D:E
]8,RQW;[<b(W#U?g5A\R02b8[G]K#F2&X@QK44KC>Qe(+VcD2[/,3L1=(+5P<)7I
eXZ748ZQI>CIN]?]d+;34gK\8=AYX]/#35Of=,P>G,:IQ_W(0I/6Me-bH2MgQ<@Z
d47M.4]910<?9RQVS[IR_7<M/MdEH5>@Ye_<TA(GWYTE:SVFeZ)EH#UV8=,?bD@X
?514R8<_TD/b4\J:X.@Q^=[QO<YJ35OC0\AbHObe.ZQLMeR7F]P9JD+F.JS@HHa+
/g0;_B>aFEZV8+^[0S\I_-6N31U2(Ae.:+0)?WQV6><RcVNCR8cbaFFfYFBeO/0a
,J^NdaT;IY55BbTDG4YN[XMf\D-?N/TL:UBaF_dd7&-WV#_&VOfdb6>/23M:([&-
#D7B0S(3M++^]6EfgU2E.Yc\O#6A)B.;8;74KH?9_0Mf<4R@aXb8@R::3X.^b5MV
O:G87.J@O2WgRJ\+86c]AgaR>X>FdTY[-2^6^6C7&RA,)2P@Hfe57Z-8@R?Dgg)C
DUa)>;^):>H0.I.)>GOIK-8Ud=8)539MWRPX#B^CQBe^3.Y_&,8226HC;BA#G2,O
:9aV-UMQX]ENOJIeOcGgESBV1Z-^98H#AWXC+,+./bZT&bdMGR^Q#ZMQ5/FMZc3G
8O/Y2T.@A/Y5g5)FH_QN6K^NI\K0#b?N&QAg8Pb+E#)1fAGOCQD/U-ARE<Of3g90
52a?:)Z#US#8_JJ4;M:ZfB.YfJT9O<[Z9?dVIVK5(VM7K:&K0Re3/:1Q--4:@5?6
OT1U[6gb1^1&NcCLf1+O26.HKV.[34QQL;UdHSY9AT>>JS17-9)ZTL5&be/b[\X1
E\)&0><\aI5@0=LHP53L23Y7_1ZPEbG8]1a6(W.7^D1eU2LYH>;((@a[T.-S6Z31
dXIEa1C4[1;FXGd2-<^4MALY)B7.PV71f3.,AG]QNYR-C@Taga848T,SDQ57D6LC
^XMZ<#>@cG]M6HJR0/E<?RbWISBKfQ#ELNFP[gAe]H5JE2E0=cFP@M_8N++N+X_I
YK[PU;C6)Nd+:),V<4V>8:::PVc&>6K,4XJ-</A9&\:WEPRb;<N)K>R0A2b+\NWL
<+6Rd@Df2e77U+-4STI)SNW3\0O6]D@)d;F5Rd8?B=_.DAJEUK.VY0;T;.e((G#X
L0@?URc#_<]C/\#a1<NDDDcV79]gggd01<P<0\QOK)/a,L4He,+(IA4#.>/RR;gR
)6@\a[S.+4d5\Q3\YZYQ0aLa/KO#.?[?]]1d<7?VF2(.E+(7VZ=H)M9a(b)058[.
RINTaYBe453#TLO.I\e#Yf[X)dJ<b@&</#^6dLC<I,,-?SL1ee=OIU?@DS?ZXdDP
D.DL(G;Kf/5I.bD6^?(1P#&3CC(J3&26eVcFDC+LU]2P29edIM4K:=OT?Xdf>#7H
(MXUP)(EI]@V5,WHUU8D:8)]4^T&NNG1(IV4SJUY#&MTZZM<V>NA5ad:6=3QJfH4
>.Q=M:_L?15]3fd@b7e3?UT2P_OK0IbJ4+?Yg\-?]X^cD9;f10-]5AB_0):M6U4&
57BS-PPXW:LEI&YD#Xf_cO4SF4,6Tc/_A\#X4a8F/8VJA_PgN=E&>f3T=>Zbc+1E
.gDAGE?X(d/RHfQ2:c[WD.OW<TZe8=DCe,TQ-0f-Z<#&U:SGZg.QIQ:\X-dM3Jf-
eF?K=Zd4IF0ePXV/Q\&L=RE@R>R6E=WK(TP9fX@[57]FX:GC1>OKQ9Y6Ea.D(Uab
#bSKZVa<E^^V8g=0QT]ITSVKZV/+:B28bd?)eA3Mf_558];3<&E#>TW2=?3N2SB2
I/X<>CcL]>fQPBEg95.QHM?1F+=8_bH(D(H>WNLZE([U>^=,-0/V+(Z6DA;I</1<
@ZN>2e7:Z;[H5UC&EI=EdUDG/Q]S=?;&;?4<>M_eBg/./XQBTg0PS>7HVd^>@<Y&
CgfCGS7G[XR@_<P.>E/.F/gaeJOB#ffI5<&7F6(Xd0<GK5c@S#dOC5g^?4919638
;ITTaNVZQ2P=G@O5B_2;a:&.aW4;f&6ST?8FBSc@@bUZW,1?C&(0B3J3?;&331ZW
cZ3XB0=4#W?)Z>&IfT;aEL+3[.dF03A]0]52)^>;^@#7?]2;fP0\:.:;L:)<0gY]
Q&+R>6K2XE^0gabNK:4/BMM=-?R,V&:E]XT\0SVb;EdW4N<(C^F:?SbP4K-J7D9N
EA2#8DgRDF\)RaNN,bRVL;ES2DQQ(SY5-2NQ_b84[gDD_UdZD8aHf,d3C\_R36Q9
eBD7+,B<SV=E?J8ISX@+<[7f=XeICKTaI>J_=1&H]_7?fD)Kd4JX9;D7_V:_a2Ye
5<=^gU+:OOM5^#?(<G+[I?U]-R4#,ASJd;A=C[)@JHODI]U^b-U.=.N.EW\XL^:;
E:?JfBR3[P7N&(#A<:D1P>8@DRUD7JB]X.X(-d5Q#>c^:T]KJb6\IcRF,.3UBD;M
H;1T:AAD#2K:@Sa_J-\I(AK2L+dT_<+EdY+X[[3^c?T=O.3&Uc#c/M\WW@d>CU#5
)P;0E4]JU/JXX9K;G8Q41MI^GBDA-QQb>>a?:/G^M>EC[HNPZ/#P;Y?YK+9-^.FS
f(S=F?X\5K&,KO#a[+K:V>;ge#/MK4I&#3><M4U^8TV23RN+XQZJE#@#/W\dY=S_
,QW?6<2>6Yb9)a0:[Dc\>3:G3d(^F[(>M8RZYUGP:MU&>I6OOKQ)03]S2@?MRbWE
Uc^&=<MUV&)b?&BSWJ\4JD39Q3)b/L>83&Y^SPc:J6I?NBZ^.f(7+(#g7G0CCQ_:
T]XL&aG\YbVgf#YZWL_R3U9.K-6YIW+65S,BMB3Y<YAQQdc2DGd/JDQL8<ZT[>V6R$
`endprotected


`protected
V7)OJ/]PbgN1<BeTPC(BbVYA?V&VecN?_^2ad7U1eUK[>#B@FRNS5)<?7)V?4BE1
LJ:4Ve>]KX5,MN^RMTfJJ0f?OB5N/cHK\^B?c_RFLVI/LIOAIP<fg4317E8H)>(<
90?8XS6Z\5+=)fBPNe,K#02UfMRXF\6fW)O=XH9?J350MI+fG8SN-B<bQM;]9VJ5
[G5aUJP1WNNHOF]6Lg4GAC_UgdK4_8((5-K)0T?7+(=g4;.CFOX/K9ZPTFI&]@_A
e#Nc?Y7UWSO;6^BCd?6IDL=FYVMH5-cE\=8<fXTQ;BbgD$
`endprotected
          
//vcs_lic_vip_protect
  `protected
-E)(bHPK+BN#cX4N=aae;RZ:Ebe4f<:H4T:7W&TST3Z)>,(FK+Ge+(O&:JGcYF1T
=TP7KGP2?:M\\F2;)Lf\JaMXD\)O:H-g4+/RJ<5QfAfB1(Z^+FHA(?RKCQ46B-F)
92XAV+GB_?EC5.RaY=<aNf@;7\Z=R-0TJ0-YJCQNe3fQ.5DCcQ]EMJX4@U-Zgd\a
&JUTWTM/)ScO>cfAC1H#UU-HRWUG&C?XSPC2c^NA^b(G_.cCB.Nd=ZH(\OeFC0SI
59WVV3e0(ba2\LNJ2)D&Dac+6&B7b2B96W3Y-X;dYJ0?b+IIa]M_LXIa8&0#U+^W
QJ^QZfgBWP+P:HM^dH+V_Pc0NaC[DI]F?$
`endprotected

`protected
,a^CM=46b6651R,aH=7@=4K?F/M5FfI[E)&:acIBCO[1.Wg^Z?T32);#I8Q/4P[Q
;S[g[FdZ][P[_J#,;?&#9c>dU))bfG8#L?_cAW=T=G)X49g91&e2BT;#M$
`endprotected
        
//vcs_lic_vip_protect
  `protected
PB=QK6.9Xa.Y-8[:FRBJc-QXa#\AUT3T^LD=PR+1a:fP#]..5.Q=/(AM\7&g;Z0P
&dOAE?=VN_g@14&OP8g7(c4fC.XL0C[b_6Z\XgZ-7L)XK1HX/+A]LL(d=TTOP0=A
.+&E.=/O5/2dcGD)S4(-d<YNF[@a7]PHI_D2X@cQ+d+&GESL0./A_D_d1Bg:?-Ub
9.Mb^[A;>3\LA+EJ04^E:;ON4X]17(.N:FJY@QFNVT](C7D:SXKK=fVBTJR=@c^.
71]=U.<(?XcCA5DPb-U3/OF1ZUQN;^LU57]K]ScA+BPX6Mab=QEKbLYZ/=6f4PVP
.)Ydd1CFaP^#,./D9_c[.#)(T2>7A&YOSd;C0TTR<e.BDaNE8.ggbfcbcQA1A.8I
<ARH0ILQbEd\DHV5S<[G[^3\ZAMFH#(Y,1IM;A8-4]AQW1AFRC77FRJ+8Ke,dF=J
_J:C_b\0D0&I45FY4^-bR[97N;<F]GJ1QR0>I9.06_<HdY(JB<@[QE]LLM&Q2B+b
^0I@XURgFY=cY)2N@I):Pa-e=;.W<T82:7@B+:d^Q917fG06D4#g2?-[=S<8]G?T
/57b=;V//?>Q>G[gK;aF=5WZW^<>80L7:Q+f8C5eY/acA+_F)7BVHM;<&DWOHLC<
&McVJYV?I.JX/RAWESGYKM7AK&G>U[-Wg@M<B&,I0\-3Uafa&N[V6>Sb#]4<D^1X
>M:^#f.9Q/RC._bP4L9\H\RT<<QaWS.:R>M&T6.XLB+.0M9/;ce@7?TEB+@d9S1A
>9R/_),C)=@ZbA<(SaDA0I#^?,9CaDN+W\SUcBF\6LVL#0U10JA)aA-aWd&a^V[V
6\T\?;D><?DE&F07D^HB\M4A,NK;:Q@72gZKS:\-+4KU0&QP.>B@Lf^J4AaZc7Y@
TEGdTL,Ce_Md4=>\D]_YKGJY.52gH:?.I9[6,07=<4&DTY._Z_@CMW=2ESXO0549
B3N,XN[5.9fJJ^1U6]Occ_adTg7dU(KK,_,7I@J#P:+GMdfRT.?6cH^;ITJ?9-)#
LM]A(]L@O_O]UW_HF^:[e\&P>-(U0P<#d8Z><R1OWb)\-;4:4M^>I,W,&#,U+@\8
<fcC@EgeAIV?,2:5-1+NFRM-c(P06#&V-)Y>,e#:D>+4?EW(+Z7UcS0;R,TT&A[.
+0J1Y].3V@8^5]E+34^KEPDJ)JTf^?JI7JAUVBY.D5JNS8#,M]g\gV28Q4AH[LI+
G,XO?Bg#:=+#)0DaL4F7O.FF8XT?I]&LeR_1:J7EJ5SBD5EJ1H<<_9.9,@I]a<CV
6DKBb7eEL4:TWCPD?ZKI(2TOJ.a,/QG1K#1(gRHaCBCSJ))+V3_._b++5]0efEVe
X;IJ#0JATS[S/6&CD/M/OF]?A)g(F3\^U=[M?E0H;SR\Y:F]<g[S[-P(d0@)C;,8
KFccH@(e(F(S-$
`endprotected

  

`endif // GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
