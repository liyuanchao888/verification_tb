
`ifndef GUARD_SVT_AMBA_PERF_BASE_SV
`define GUARD_SVT_AMBA_PERF_BASE_SV
//`include "svt_amba_defines.svi"

/**
  * Class used internally by the VIP to calculate performance. Typically an
  * instance of this class is created by the VIP for each performance metric. At
  * the end of each interval the values of this class are used for
  * checking/reporting as well as updating an instance of svt_amba_perf_rec_base
  * class which stores the performance summary for an interval
  */ 
class svt_amba_perf_calc_base extends `SVT_TRANSACTION_TYPE;

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Gkwa6NyhYFwNGZhas43ZJWCsOxyuCw/y/KffK8Py0GFtrZCqX85vSs9xZVvXy010
KGvpfYKOisJ5LOxrgp78C7lTn4Fx2N2xAa52XELC2pdqk0a+1fCH3X7kIldF/YjC
2fvLlerfmLtovfQ98UtlcSLCwlQrs1tCWT3zqI9cbM0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4446      )
AyEMFXAjPoohT5d2/au0+X3aT7WvTjKPx5wjB3LwFdzzpgtOe6RNnnF8g6Qx5mLJ
YVMetHDpa5DhEeFfKysV3/ZLL4oa17jJKZ9ECqD9m9H06EqzdgvXFapsIlk1SwwD
d6bf1hrIv55w7Xh8iEH/CHM4WqnGDxLobaTVE1yLI/JwJ/vnprHTJnt2A9wBInet
X/UUaUCodVmUj2R5P2ZcX5Unm4q5P1P0/c6FB/qtUU+RuLg8sy/Zj/lys9e8eW4I
YiJV5AhtfK3IYr5MTIf2fCfqLS8+WaXqAFyHy13P60fsyPfmfxYgOa9oO9WMbf9x
ThfmCfEMO3UbR/VKRA65zvR8sSLVEl0QZhdeMCnlOri77p3dpe9L3CToATcLVt1h
u+xjtyasV6fOs5fpCZE7LhDRKYGZh9+mIIzUD3tz8DdbsORI68GDGWfrhLXv9QFd
Cmwv8rpLdYlNlM1gu9/yeQU2paG6fXDIZ8KgF508b5amxhBssCycmwZR+rfSqJ3L
SED+12TkNVXkLuD2JE6xKfpY4gSx9UXjdLtrOUXGuPwaLGFY392DbeIa0Wij+q9m
z6TXlPdO7dcfcgaU/XKhnw9tOhL0AX1u1VWlf7oRdNJ5eFTPOCUk45rPZ10E3dr6
K1jRU9E/M4sky6blpb1EjnYE9MA2gxsJGYtVv+N8EdmWDfsf7cUH0AhvYLxoE7Vn
Tvcka9r4gCvW0mcf9vs5ji6wDcKGxYxwlMtdN//Ky8NTCtp5x26Ghu1sa8SrH6JM
faT6GZl0dFJ0Idxx3kfYfnvdnpO+QTkWriUdDGQcgJTuP5YaUueCXE+TCWvEuFa3
x/MGyCSAPOXShk0OoS07fnClqx+AJNOxzr/fMJRhB2nDx4VhYqikRIMLb5J1gwmT
lRxKXUEs+QpckpFJ9pp6HSs/swXwh13CtCCYLu1ts0q5KLpxOlXQlARLMtMmotqg
NGxGvjmZn+jVfaoypYX2cpwQvpAqPiBexQT+sBamcKGoir3+SvQhFqdzls+k1HMm
JU7xM4DnLG6PY2903v4er6AECiF7WVhfbKjgbfPLo7v7odP7wYLrcDaBq/6idFzt
n7tmTBkfq8HyTGXc6L7cbOqRYl3qGMH6HzU+4kAuaN/V3xF0ElYHFdvIdoyGOpMe
ji5KdybnWF45WR4oZGjR/ZiAza1Ged6zb4MOr1V0WPM87+H9V3KNTRptXOk3O8NP
2sXa6VIhiEpYX+blt88fA166hcTWzt5FFy9DIY76m/gycSB7jYRB4mOVwJEe65TM
zwuixmp7AcAPNhxC7W1bHLvuiYJ5CgLfbWqgzW+bzKk1eFtcnudnwDzWply9kxIQ
/ZbXGLOHDrF50SjSOpDu7g5ze9yIGLlHH3tMUgi8pufvZ1wzdItBqT9qQgehLmnw
sFT2pAc6EVqYTSmeFbDwpBWmRof75RkfsizWWkEYvzerKMJ07tF7r7P04rdIxtQc
l7mQfu0mnALIMlB3p3atjX+py1fhqagHvTtoLS2KQJ1hQIcskAyHV/vjNSM+ggyP
tDbwb8XE2ZVvVYn17rYFkPxA9a5JyLiJ/l9FOItRzHyX+ryoulXX1MvzCb/Vu2oe
1h2BFappIFFkn2FvhmL2RzopDztbjLOZb+7+hbHK2Im/V41bTVdEJKqdnQY7YdxC
W7TmFR6fvhAQXs9+nGXkxNz8/e2D0aEFDtzRfMuqItE4QPifdFb06eM/L8cisSzt
7vLYY7nRKvFccnKK0SyaP0iuUoOKno0bGl5WnLfUjnPQLDdgw7yYpSi3ovKkbHXM
A2OFrcsVkKmlfhR07VEif38BR6hzg0Aiw6zjTCEGPbammDHjT2UP1WnizwCPQ4P5
DHGkOAt/NX0AK7avYxRdGIr3IofwrmJSaWxaqKMv5P0x/nCBAFo6zWLkvPOGmwHc
wJKsCff9nzBuraxPqcGtXxeWecdAlI22sCAk5+/x4+bKqtlj9wuDd6k0CnFHIXVQ
Y6eCW9zqyEeAk7cDRQiLZkxBhXXvXkckQAGDZbyy7EAJwra97EA6zLZF/u5R/Y1E
R3FXyoahrxaoOrmVYzu/kU2qHg4misdkowTtBtxDXNFcv9ogdVWLmvFYYeKRa424
xP5S5tywTO83itrQNJJxRQw+DJnkR+2LMpx00/V6yvXxL0WHlDkSbAFJU+SO/npr
Yc2WMMQ1Ftfafwbr95E/ei4jYBeAPF5i6lrK/Tg4U3O0OS152KIQJ15xm6YitmRQ
YmfNsNYsipI4m78d3/7WJPy0OsQNZUj3PbHsdws0PLB4dcUigFjAtgAYdCZ9lOem
2bVtRGlCUUD7h3LRAyUpAVz6g4rIg6m9nm0EtYIbsgNAXfOkD2JLwu9sBfuVkPMf
D0IBv/l+vG39HFsjAa2MQZWUE5eQXnS5ehSX+BdcvNMulkLBcRnQsZ9ZiSaxNeow
1JyCpz52Uv/KizswhEe0/ytYdsaZ1+EUT5RyaCS30qofJng6xtSCaaI1ZRRXOZIf
nwceezyjcsjr7jIDXWXKAHTQivv69Ungs83QGtDMqlrRhP24isPe8/M37NMgTcOM
2/opjMNe/KY2AzSoJGjYk7zyF7BEIxmZFv0JN+Q/KtGKZeJfXEe8+Ip3Y/eO5In8
s8eVmUGZ52Y+kxOcjcYadL8ZvMj7NTLW78eQ9E4YEFbGHr6zO40F/xayFziroR08
DIOqARU/jN875Yw/12Fbgir42OXUoUS1f3zGCmtYebwx2gPpTyM1+PxsrHnkmQkZ
PnfEvxdCiX+BymlcsgpOIwy0KLQBt81eMaidgPL+eoUHYry/hvrfW/TcGUpVB4aV
vofxWRhPfdJYzv1d8nqbkwUbkxURhYmeLZ7+vwJ2SILMN9l4KmuttgQ38azMHt4s
MYXsuL+PfI5uIWaLcPMuB2eI/I9hYQcvuQpG4EsvLVVQ4Arm572iYoY18jQx04lu
ZbbCtrLWJPIozYFTIsmuvpwyvjEWzKanNLpYZyFoCOBCJPx4mcAZmMNUpdcMns4m
sUOEgSSG7opM1uTF5pu3s/hMK7s+OpMkmDS+U/MZT4tS34U9kRFQEoZFeVtEHOfD
Elpet5p/vJhlRWrYTIHXSRGmLid9AighyM2t7Gm/D/6G9LaGsX7nZubRzhtnAdR7
2fFKth4oX8/C/QUXbu6xnHhCj9F2WjZoNWpd2iw6sAgbQdY4gqEq1Rg4UDf9YNF9
B4NSt/FyOmjg5AAysgmEgxy761h3j82fhh2c5Y8K6NpuQsQzm2fEkB+3JCJCPMIo
UHQfK8IdbKMxXhzlDBFZ4BIWohLBmjqeMWUXEy+rWK8ev47f3y1U0bSJEx8XNq70
5wz9kclFhdmL/q1X6Xcezl3K3ngEoDXRKkSqnMLzdIatKV1XwIaq6uxTm4N2hB26
gMrX91ir7nmFAf01uuZvEju+Vn0NfpFOHWnCKtvtMtWEd6+cqRX9wBc3qqhqfovZ
3fHBXi524rWnwn/XaLbP8YI2OhH/ATGJO+Fq75spFboLxyRTImUrC6xkJGQiZtB6
FcYZaYbOMS27+mnzh4ERtUEfYj2vWXlTjlT8HaeMchY1R1cuMLSi/g29w/UNgC42
rGRdoFLchl0JY4prE6YU8dBgyzmk5c+pTNCboYVppeYpIpnHBTTsCFNmDJMR360N
4LzJzT0tCRRSmWbkxhSFhiD39BJFDOAibzSJDcOPLBmtYJCwCK5I+iqa2JaLYuX9
UR+6VGAurOG4hXq4/VZrqElf/oAMllGL3D8OBPMJvDTrIYoSHqlJHMgFQFSuyqEh
oBJ2SNRkaf6CO56+rwWl/6W5SShSFTMR37Jvg67aZMuEHhOZ6q7BXjuXriLliKiN
LZaxInp4Z1gV6+UMSvwVTlxAQimd8/zZB5d0YdklYFczqm3fi95cK1kswqXY3Cmh
bUvC85/WUo9NQv35mYrrieCFALOyIAHkKrhcn9Q0zTvhSAzg7tIZNtgtAvsfCT8l
MrZgNoU6IM4XtSQuwb1Y9PWFoGubG0SjVL91LWp+6YOjKLPqH6sW3wsPJkwW6iLl
juRkz4m4eoFADvGftf1+VXiV1D0tTX0fM12L3qm9OCZwmsphMO2Xq+2SVX5Aud90
uO6sbyrZT9EKm29L0/ZCGj/lMZaQzi1RMnciyWpkJhnhyVBMLe6JXGFwyt2qOGsd
HizNzuloyv3neqcByW9VwyOU3SF1JZv1sEXuxZa25N7E6M8VfB29SrjarbEJA63i
m0w4lp7iBeEno94y++69OF6gdd2LnMhAFisW0XYM6Pae4CUsILgMShSIXJRiwn5I
ns9cpzgtGMXolifKojl10sx/oufR25hyHaOzQc3jWh2LlDsiTzYCLUDLRx7Aj317
V98aSdYrXSEo39x1Aek46WtObkHR2hT4KLXWKWnL1kWCvW9nWrlyWZ/idcgRMp9V
Lq6x7mpE4nlA7gquanP7InJCz7eg3sWILXllVbfg/PQEhiPTJXxrG0olwvY8FkbD
u3IswQUgL6iDqcVAJmjqiB726lOC/77ZD8smgZyeys7c6tZUoklXQw1wI1bltpTf
J4jlG8s5KpB7JNTydRSMPeyBlNIVEqVQMxDaRt+aE44cFtj99qhZlhWo1n7OdiIy
u4EKVmM2DRZKTEH+YkXZiFjqh2X4JoByMc0RUY0PaTIYs61xnkqBiVb/8npTSxIf
ZxmQmu04hvo8VKWeVrGXCkM8KF8aBH8SvyULe3jajwHWPl3Ikh/wXwyKWFXmMvdd
UzH4BhjlJRKQN7lLTEaJSIMj7TLxoRwT0l+VSmiYTNkJxofZAqpGeNtqRSFU8cwF
IolA59n8GOOIuq1UV59+Cs6tYVq+1h42OSLPxw9sYctFOBAhmUyD9quqmZKXd5xW
1x9oy5YyYSxV4Pymuj+LGNSWq5QD7oMUug/AFq6tQySz1SeE3HMGqqTCarQbvCtt
xZF7lz3uNHT62sZJfqsvpyLvv1R3LASvzHlZO4ir28C8Leg4WSr5O8081RnaikQT
fJJ4G3vv7IC7GoCiDdfPnvvzWbNsvdHlj0cmKJXOZD6n6Wh/vBeNgAu0wlLt5bIl
xcwzByXbSqs+TW4paUJLBazJRXuunz42g5jw65rpVy2i1bzHwwZk8sTX2Q52JR8G
Lic5eLXXu+POc5Fn1QnL8FuiGB5WykKbxFG4HdS4B/7XYms1yQJrjtrfkT18KZvk
DSOK255eB/qC5Z8hlumlRH6uiENcs1obM3nKf1O+PKgUBQE6vZo/Cu9IZw85905l
W/lryWrIKhsto+x8BwrlX/z212I+B56tHT2GkCbdwyTJsahhw+Hkbo1A+hlifnjY
flHkQyh5RuT5HG3J6Mk8YJRvmVAkOtJgFx/Eimd3yKxdcdURsz+89+88H437gTHA
7Wsmz3PrPitg0LypmS0zWtGVU7LnOw/zffohtHj89NjUKeBWLS5/m8wD+x4Gr2e2
c6VnMspAx437/pddNuqYmjnCBIHmyp4BfhN1VT1q/J6kUErpRcrlPS6bdZ+jEBbZ
ci73uwwyLPZ2Cbde2GGyZh8MC0R/V7pE3mBQgnNc0bYtTSWx78ml8/JY+SKKR+CQ
VbY5y6GEO6fvOI1InKtTxGxCKVXr78M58IKieIvXrK04HPMa+5EZ0X+VZVQQL67X
hbRAfIsry7t4rtpGF4CBw8ahSiGyL4kY05gYlzjhFBxHMKKybm0Y/2GlIeFVhJH5
wpspCZYniM6g9FxQYdCDQ3jPxfqQmgWcVlhRB3a7/j370tlJ4AlCQWi7NHHoBMUQ
k6qCNqUBhTMuK5cmJ7AKuUIBs5d8h9IF8PwBMYgW8D/LiOCdA1WyIYqkOfO4X8el
WWCNK8Q24M+LiOagn0uiok6VR2ecLOb5chfihoXyqC8z7qiqO1L3kRlGQ4Im90yZ
tJtq8ewCIp48MPiYlmO8X/zNu4MHo322NcE8dxKBikc=
`pragma protect end_protected
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
NvvqcvccOdkXutknCWZPJ+wpISVP5J4vnDsLCWVhddfGZZaq2ZyzHKNVzHLIf7aQ
XKSOxUnEpBN3G7pyVPi/l90OFUH5EoHiqPaJbmijh81LrMCn6iq8peg01Te031hF
S8SDugFN+VLLUxbWs0SdCIsAVs1yeAvg3CahV3sm1rE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6816      )
AMbMz5rURRKSy/PPXU1A1XzxDhCJp/gjBM7DsHXBhEWaQpVmnCSj7iMH7S+M3UoQ
xWec/yflcEVzDvy3EpsVqVAXHzWS0j9PncGlAklLPxe+rFK5MnXsLpfsCc1vr5G6
EWe2WZRcNY36JJ3QJS67Oy4Xrrj9tEOIiOmNPaBc1X0q2V6Iz4HbicbjJkYDwvJx
kU6Xufepsf+OSS8Fyn/d5K+kA8LlvreA+iB0Yc2kYDifE5nGjqJojzkjE/pR4CKG
G+9gFNANhE+lGisdpdIValEIv/qmZTtB52+ROS4UtG//s2lRHnirtH69aLOPOUf2
PWk0YOy5D0B+fA8BQ7gpwoWwpSTo8bm7WejKmGxMG7Jec4NdrN12vu1gkYRcZ2zH
+SDqjFgtEfWxn81uVn2a3srDbW5wLmJnlSvy7+TKFTMIrb5oqKXGXXrxKDYGUs7u
vlfpP+wtT1Tm1c3KyOGucua3hNiY5mr8B8vuB+BdhdhROBCbmcJQpc8T2CPia4Lu
SMNNs833WWV785JVN7M9+8QldNOYjs2EJ7jcwGwXrtdrzaJSGTzfdUSVFOkJIkA2
zVI/Z2R0tOdtiBw3tG3nL4k+aqG2LTwqqSyshIHndpv8eCJ20zdbUl9ac8A7AcPL
bOzZD08edtyXOlHMTPYdY1GVMCIKQX1XNbev+xJbd1d2lIN3S6U6amfAUPM/EksH
oeok2NfHQnNesmKk3Hs7A/V5dB19xGplq0WeQCJvhw1Gcer3bs5aLcU/8a4fRIiz
Lg5fEJ71LtnHrh45CojYvbTM1r6vUS5kQDNP2j2Lx3cXqNgkfDWx+BrvlhPwF4xD
zTLSEWcCNf9gWbK4uAK1hcoNnSmlV2sov7pOkD3W3TcSyT9mIIjkuxxEW4ECHrPD
wDz7lND0h9hMD+87I4vbMaoApjtcQwZ6d/h0gwWgnXJHXqbcaCgYId7+BhyCu/0Y
DhiAZAyyAjuU0GvcZs6PCaERtVnSoPdle2VOyZGnVzwQRRwN6RV5jZdCMWedGxEG
FwPi2vXpsyGm6TjfqVeFzKSqDwJ/PUAb/3L/2KKY3GtBFJ7720Qj6yHxbRq+YXdt
grhccuIh+G67SIVwy3NAfj974gQz4wJoiSEsQI0dJ1FmV1u6ZtSrc4oXn44uyamv
0FMPXV9yub4QPt9l3BM+JJ9PCzaaWkzQ4mqf/dZ85emrlmpZksnesvI2ErbllVeu
eUMfFSVx7svl992iD/I33+U+86HFoAkSgJKFHaQ3Y9ZUXgvatqGjcKHaaRaLLo8Y
T8x1Pbl7vb38MhgMr8PN2x2p4Fp5i/nCPSb7YWvHZfo3s3wzreozQp421PjXG5zk
K1m74moEvjLFB33XsW3Ue7Qh7Jp979AxTPwd0hFuXQRDfkVK89KE3jiNSXRHvz2h
uir6NVxucYmtFslsHox4h4qQ3PiOcFvqNhYthQ9wSFoU5DtcLBr+0NdVTp4w0ZFA
qGei9OOYDKQ/0ZA9I/Mo3rGcP0i4d7hj5PWzMQ9NcNBJWgFehb+/adBhbS9iOSP9
YueaOcj9NTAyMh1AtI6T3pwCi64DC/EtAueGVKejSTEYkUiBNRnYFZ1Xan2f4Qvp
TDj76/pKyX7IXIDkbAqA4keglf0O/zXk5wgGGKQBHqkF22O39L4CO7XvbtcBBBNE
s2FQ6ld4K9xhWOlrMetstWG+aMZGPoPiTQqhG/+u+mVpI1gqblZHvRPgHrYk/GlN
jvwPpeTCMCFDBxUBkjxmiFMM6f6VqlhC/bXVKZlSeITvvcTsQEKE996A1D35EtVN
T/MHBp78vcljGLVS/fVBrj/BWGYVnz7NbDpFjMf8yAOD4ErSd6S78+Cs9gyUFUz/
w03DYh0lmM3mYzM20vrbKIhu9NB34/gvC8vma5Etdc8KPcCSHA7MM8lTh9TJaCDH
la+3gWzP7io2PueUBDazpKGtBNWQQIfV26IoWZJh3m2+X409Qn8rCwRUr0MCDIlW
zlMQqP5JYDxhBSeXtHuqRTpvfWiq1flX3INn8RMspG/L8zJaXEmSeTtsTIkU5nYb
n7zxkIWn8O7xK4vmm+UbLBKyZaTtLMharIsGgMo95b2e3DzzfRtZmBGCwi7LcwRO
ko4ejN1Izsh2WxwLvJDrJXZ6JN4ShWJgzLJIupcQK3kIvCV56Rcw6+oThTaqrNEE
tymyoT5tToJn/HZlUyOr4kMmPEl2rYFoFn+ysjA4VjRS9a7OTCGj8RuzTxllG4Q/
xHif2gAfbR2cL+YBLWmEbnP8CC2xpCfL6HISafzPuZFbiOut/2pwS/ypB/c627uk
XrJLrmOX7XW12nCEEvMEmkEcUyPv8LkDiYSBCRoMPzzHdjZ7WlBRLfJQ4PlNJLGY
av8MFmR6KRNCC9MzAACmNab4cygGdgtfbRxlIT+IB54cN2CIxZwcyguUmwma2uXV
y2+XpoHGcwH/oTppLsVoLUywTgdOzLqPqUWgBD2PT2lx4dc/T3ZuGc53NLZOT48c
d5wzUqpTrLKVG6qmuurMXvVf4WykZWzx0dVWQYNkOShQYVCknN6CX3T064XDyDDJ
gLlhsUJjFtKfME4ieGFpX7my1Ms4Refqtr/Gy0uRK8SwbaIjHPQ0hyv7bO16yO+k
C+NRsyS+uFs2cYsXdtwGMsmkfkZctNRKi4K6AZeT/T2d0YcuSL3ojvLgMwqSiJaD
kxFmLjK14o1NxhJs1LzUAbISSg2uStP9GKhlb+zxWiunxzR6CQXUwr/W5X+iq3q/
LDqQsfN5VsfngiseH578vHOEDjEM1TYVIAFetSpvXZ2jERLObP02U9awNsgic3nb
5KZGKT5MRnqgdnWAYec16ktSiImzSIgFnRAV91x1E+EenUfF2Jr+4ncklP5G5CUy
Dz/g8GpnXGbjO++ybmxcFK+RlC9b+rYlsnf3IPQdMn0Fmbq16d42NRpNVdD8w/oy
Gi/XMc8CHOKnj3eFkoiUv5Pj1rBT+OkHLeGxqB/fObVZ8thiFQiDqA8l7rLNcHbo
hdjw1b+me4stzNCFHPKh9keHzNE4rLRhRy3fATuWk/R59Gw9dKNED9Qzb8XdoJeM
5Q/xCJMwwZIyLVX7AXdZA6cEp57i7WJ3szPkabricQl9TWtpTJ0LlmL7FRAheYug
mRc1z84TDNnQbj17BmMV2hM+M8aAf4HQ9UEl5sq8DzE=
`pragma protect end_protected
/**
  * This class records the performance activity in a given performance interval.
  * Typcially, an instance of this class is created at the end of each
  * performance interval configured by the user and is updated with the
  * performance results for that period. This is stored by the monitor for
  * reporting
  */
class svt_amba_perf_rec_base extends `SVT_TRANSACTION_TYPE;
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Oi8Vh6oxJsUdGqBQn60Hj7Ln9danUuXEdu3ObBB+yZDDCfBR1qQGqvPX1S+Budhv
LiYkoU8xdH6HOi1kDSDVn6VdcH3gj8NtVoQmBYKONlK8cy3GRE3eynbCOC2OHfEF
3oJa8UdDLidVcDG6emWcERrqFSsvFsUCZAkf7/hL7oc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14691     )
r8XEOnrZ3/UYSGzADL9eKACCapPbzg5H4Yi0xQtRf4DoX7E2hrKHwUXz/e2KNHhc
P1BlrgrM3eT79LZArjdZf7PdwPnXXBhZrQTSQomCn92FCVm7XPT4DdX8ICszynRk
sPhlPy1szHsOxSKqCmVLRb9eOsW3L2Uyrw1AH+sNRgcGvpGYk/kZ88eOlZsDcit4
Rrp1aRQaJgnnAZvlT6OL0aNxmh3J5fs1ktmOJgzfHUr71CYfEjTkrp95o3CKmjMz
hBX3KJZGt9FsRCmmEBHLzP0z3uaXm2nnLWzr5svsExIECHpo8IsX/ipLp85Koa7d
Fh0s3geKPTUuZL8wdBX7PyUFlEBw9bvmMmolHBGAE58hixaoKJ4/YxgcQ9Fgsjnx
BCBVE/D78xIm5E/0tPmZQYTvOXcCaB/WCSpV+gxrAP1ZESxGIsPldXcM5fsiKg7z
eysUjx+oMcFZf41k1k20w8zvoPrOs4HTKNpZiDHjIe/DKS5W8a/whhYj7+P8JnG9
GwieeF75R2YLquAfWj8bEaqre/PlkTbuPafC9zRk91qwvXY6/oNZbEddEj3YpARj
Kt8HBRlYoCgTxNGkM9a0MYQNSk4q9fk/DNyn0evqG5PwSHf+lH8e09hTk4GwuIEj
pGqD8IqOw5tD4Yg5f1yEfHtJWw4kQMdCF+MsJE/b2OlaiTNjjNN/+xgO8WUNOVqI
n9AXhGoKZmyL1WGIDrvN+qjo6NbujrqKEcmekwV2g/k/q01/ZK+pApaAmX1+XMm3
YR9T76WL4T6QyDloG+nuaExnSLp5CaQoThYswTUMSREi8XDimXS3JW8DVg/314ui
eEdnJdUDYoDf+Utcq2uMnNMvAOwmEXiD3/qkt4SaQmMFmR0V01gSzuIyo/Xmnmz9
WJH7dDdXqNCnNEvrqzv1iXHSqDIE+xzmluMAavnDv4zcodNyNJA0WEf/FbDiTuup
v17UzPN0jWW7rL9G8EUtlGyQvLKBA0ei7pxkA0tUAFtDHR9zzuGAhd1qPb3LEECd
+PJ/paiQLkQHrUkiZD+0yHLu3cOzH1z2Trl2VNoSWzCARdR0Iomrxh4QbJTU37xv
HvWLsDEuFwcsD/ZBEtBwQd9wtO6nrqbGIN/qjy1GKjzCybxUSm/SaJfifpr2GWjh
E/go3b6OhjnK7/GWGFwDXey0F1R1gI9vDBchIIX8LRwdMsENF/kDEzQkskn1qCzW
ba9AJEktUoIaJRzdZ26+BHNYPT67HIbzEN5utX9QtgstqeSQd1k7HZtULgsQRVkw
ZsDjBemJIWm38ExeiSiPJJ4cAU5xtoN5Rd1MmFbNQHcCvjCxlDLyn2Hg0N8G5T7p
Tsyo8ghIKbx9vEq3+bdpPGNcps+JvsJS7QHGIS4spS8TAaoM3N/rygawdzmsiBtj
70MI/+7+5plp5nOxve7VOoTjAibniX5Nz4WDHblfwK9VHLtHTcWAeFKAXzCfYtFy
IQ0KbTlDzHXXNuDylPr7Scmq0KGpvfrta5dt4no2bEwr9OYzq/8720tpm7SeE8NR
nIZQibbkc1zxxt9QYQzQGMrMA5aJ+omGjbJtdtodCGNjQgp3KANtZNXDOfDWgCyv
PRQ7Fskf/7qEFlYFMmwAQBES/ZkdYGAKtMurofZ0Aufi+m0vtHvIkZWYg6CpN10H
YXUYduS4IwONq+q2y3YuPSFOIbIZr8PZzkdMKj5vyAebuy/9xmTTNFnyiWEt69UD
fF56vv3xtm3t4VOIAeY2sOnufUzmTJYhMo6cUQj22lpM3lSWunLpYr3hk2BU5ELz
RE4+3kq6XBBUPWGwdhMRmPquxv9LrdHiHM3UiLCR7CPGB4etgjFQjJxDtVXWTLPm
Su0CCk19s5iqtcCXsN3tpYCK7FRzmyQaOGC0DDDJd5s8ijO0G9rdIWjow4USxuLH
p60dpE+70SYVhxtQjg7MfBD9aoFoIFQzW8VemUQZdBbOH46lJjZAx3UKQnAmt5T8
I0lgXloIySjWjzHgHrQqgGuN2ZmOA0VH7ByOoHMZx3Zulk7IulnFdzaeS6TWSqWi
CZ4Ervb20Gi3VQOhuCbbitH18tQY5CJyBLWu0ZRyLSDdpbeKyKj+jidKPBe6Q/bm
awbNJEZsc0bj4CbhrUW88EpoZUCDU/ZSTWexXAv7Ifpz3dEu5KfKHyI2xv1ETfQy
FJo3LfqtJ74TGGhgchpxOsn2KK651s3cPOZWxXHjZHX+exe1jnueRnQbTlSw8Wcx
Ekid9IYKvJ1QIhKmIQ4CSSbxseV0Dh/Bl/qBZMkbQ616HLgOw1HR49G+Pr3FjjDy
Hof8/wLZx+Nm4uPDcYjeI1SN3/G22AQ82LrxR3jzJkDEpT+jq8tYjanatnukuCFc
3z6mcrlISWwn15yXAvgvDqkOqSbMMU1nqHyk2OlVCeR8Pf87IWwC88Ss/aH8VCMa
cP7TljjzwhAA7P9bpjUzzj8PMXJKWWFzqZKMxLFmfW1+WZ8kSh6CalRRmLDz8Czt
C7SZ5tO5pjlw9K4ti8LqiKGQZsFw6Orv4uSY0UOS0XHFyzDAsWfLPNBY8FP0lfM6
LLGp5GLIXnJw2SnjJQyllCuNmQ6aPiTx4r8oaf3hQoELTO3zrcTi9jMkmOL/uvQU
T0tk+lksJVgWs7vT6jp8dg74enGcwxhr5eEpiyKnhuYxXmRlzPPy4sq0RiogSO0r
H+rx1baSjMHDV0JuunZ3fyScO4J5OoAvP6KocFIwRt7Ui5ygJE1cpuDMrTOiyMso
Jhf71ebG+DCrjhGHIfTS8KIaCOC9eN395/x1f5HvAIXCmyOEvu+0mmPZj4ceShvp
tll5IO7PxHZw1WGl3nd0wRwvfxCBmXaN9dXIlv1lBY3t5ymf1sH9uDU5+kebwN5W
7kTFzNwR8x3m+auol00my9PGMYeK6Gb2gvT5TitEzNxj9IScBT+MgPh433Fpl3ni
9TPGJbTHCs2qPL8gNqArFJ7DRrWGVqcez10iLtUgniU4mQlSuYvSVlQ9ums1H1dE
82Tea10lF4L/LhyM1vgTJwtotKVCqWLvb26RTh+/GpvIbKnI6NURY5AsgR+6RsuK
gEnkbhDgAKEy3DGI1+aL3NtRUqO29TRXXDZ7L6uGdQ/9BrzfDPS5TDs5L1WvnDWt
iB+K7zd4ZAT1qVYxtqG5SFjffXqGKEsC9xktNv2kQIhwA5mRmJd6fV5oy9El9v6d
DW6UqWu64MxrrPnw66z78FxbQXaPgu9ozIWIMk05xbAGLkoUMFVqYDeDKmxz4OOM
kdoHO5YVwxi8CRJ4A4tNNwUHzQfd24Eb68DSrrTNBPMq3H9uWDR0sILCx4ZVNkl3
DH30LG9RNUlAtVqRRw/GNavX1IGK5N0BjdqPYDczu9qxEezFnbVBUf9h4ORAR2s5
tXsPBOVX7B6/DKAVerbrJCS80osJFvk///Tj8uyk/UeNrbY6/NBVryZ4PI8rEtU/
wjvoqP9zdI3Q6ePJGMgORKoesrz+fxXCw6ZdFZniUsK9Ff42FL+cSY9mwxlyc1nW
dayoWIPqBlearEq8OYRKRa7sa1o+0gxYpn3Lo7nHQyTnjYFVfEYp0ITsrjNisQbU
CVHal+QBgsaTIDcVmFQdOnQljohqHHY6uQ4hAMLTKeh77kXs7qkBVDH2QgzUE7fE
LWWxXoFJ9VqJbq4n2cjDkhz+iqqOuZLXih9IDwJrKcDMw/wOF/j41PYQNKZQg/iu
8MPNYBbShX6/TuIZ8jhVsXcqUElmnzBUFlrJ6cxfEb6HBG6hq6WVrKDEg2jqzoNL
RO+fUnxwrUwaY2VmUKpcfDiW+57lC+gwjI16/+ISvAVtlo1lhE1jXqtiu2PkF0Pv
cb8QLCKw6LyrJocMdndc+St3hy6So7WGGlEOl410HTb5p3nMbsAXwkZUMaoh7ZFm
dpsV7fA6XNl4a47AOFkCMXCWtzY7owCf9AS8j8fra9ypkSkq+5X914pzxhToDr2j
CFtbSCJt9e3PpD27CljDCZnaRb1Ewe1nzWyHe2Z7Cj9EH2Mt9CbqShub1t274Yhy
f7tBLlhVnCQ1GvXG3nDvImX7ButbU74L82txn7g15hZgxIRgTZfFBaoTkzOv/+S+
z1tykdDuN/1YwSA4x4Shyz98oQBpNgys/smxCRjTu+ilv2j11ZsszIW8IJwYrjYs
iKCrYvjFCZfLBupScg2ijKfB93XBu1TmJiOAfKSLXNl+0jiqgjAb0FUknGJL4c49
L65KGzyeXOYl16NGFOzEkmUKuXlM9jiWNbA6BvblseBwdR7eUR5wQeKEiLdIOOxs
GR5YLFe6EkLDMVHnovz59NksZvCOF+kY4uqM+3LZsRrrgwlRBw4j7EliIWWAg6zm
BXIfsUlKjDbEHHnQ+ugtYm6z6cTZgcX3NcI2tkap/xdOLwJCeUmdm0uwDBXdLGqv
XhIwWGYZV5BXODbzBJ/Ms/j/WNdJAVrO7hNbItCU2iulwcS+gqCo88K5FqMBZDmS
tXRA2ab/5mXlewHBPNqzO0xfh9M38eBG1vaJQ/R0hBy4vt2xKhmVfvNPuKykyaDT
iJJpTt0NnRg07jTgEAez0s0qUsqWEUAuCcO1KpjovsJY9598jsV8Z4xvV8cRRlxP
QJy4XRyDQBtppq03N7Rrc6jsJuNWSrajsRLiItUQajYqDbtMmbTexSm03/qhDFZh
hVXQRyQFzb6xKzWdnHaUQgEZZwjd+xLZQGhl/ytX/AyXPie7TtMu4btFQOvZCdYi
3lSoU4FY1g9ydjJmy7Y/L38TvT1lvPoLiEZu6x+aQWh2cJw0hv7Wp/SxTOZN+JiX
J2TEcLdOkQ/mkmnNA/Nm6GlEqLpQQhpeL3PHb9qGn1v5rgv5+Ku/XdMA2cq/MyhF
141REw6UKYdbsuMnyiBLOfrVkrl6PrDDbrEnVfcVOJ1sdFMaZR6ZjkWlQG8EMsPE
UR2b7VFuI3oejHpcLU5GlarWtgbBLo98PQeqrKO3Lzq/a1RrRI/DsLjRkNVSM44Y
76QlaRAZE+tHpRSWZ6Dhq2+/QgV4UGW9rxkok7OygiAbhNqQEVk8uBh7+5pljZI9
UsZ7uTpgBnq9EeqqRg94QtbT/fgjrvu2Ktv9wF6wUnXS1rPXNCUQZvbFuRG3CVmp
G9EC4BdS7UecACS5Q5ppXmho5hYrSddFgYIpWZec61MZsekd+4VimyjZxLRoWWII
1UlCT5ShUl1mmoqwmX0wDE9knOuovU8hOncRhzHpQ89oxr7gwuiKQmb+PJQrzQzG
LaLXCOSndns7LSjOTMJiM/vVnWk3E6nQaWXLTd+qHOOVZdlEpM5eygrFbGFTBZR9
IjVOHbUCTyVP0adlkRZwY6MUjcLNMsG5cN6vPbSBwvGcci65P9alEyaEM+8slM3Z
l0Z6a1smCZWAF+jDaVghv2zUQ7cGCUxzMQ+ooRbRw65/Sb0hqcG6WrkrVS7lX1GV
S9eD4zCRUtxbanGMEZTtbF8LgxoPpQsPAKA38WCr5a5tRUlnjkX1F1FEPC3MTx2P
v7a2PXIq+msC55P5BCCmg6OxZzZHPQKt7DaBg6pJZNiMmOBszKatff2CMcIqCPKO
gfl2czYqu2vb9uhXFpOETwZFtXmf7Vkq1xpdgUB56mQv6g6X6iwi32bB6faPQ3dy
hDOJx0A5ao3yn7QEaVxMphF0tE+ghkT3P71vSC4BaGjYirqEHzCoEnOff8xNktYw
0P5lwRN/zOb1B7ooH2L7L8JuVIx36+pcrH3UZlWzePmzn38w4bCJvOkEH1oE0S6k
aYlE7fEWByXYbQ46D2mpiBp3OD1BO1UrVgFNyDYa19+D7yET43b2lN7rMw6Iq/gF
AhXUa8c7553HooC4sz33/+XEGkcrwPZwwch78Lwq5mUEjCx82gq6gL/5ydsuEG9X
jgSxly7pTQP0o46ohPzSf7VzBgDeF1yRui6CAJ7QcLT/u8JBW+EQqrVcwmeHvKNH
xfxzBVJIS62z/cwnWNrKo2vPm9BJJ022lMCMcin7YRmsN8MxBoggAkHAoJwDnXaD
E3DWs0Ci9Jca3qxcdvBxkZqmPhU6Uodg20RE5AvglLxVImkpy8l4/+uDw9+Mm8sK
mT1Kx2bFxnvKKE0118/AcHAbgNxaLQpaPPRY/vK8B+xfncoZMF0i1TH8DgNNO1vU
T8wHqUrP+3W8ofapGLSiQIs51eQ/p+o12fpVVLZjNnn+p+Q8KAizPz1vrGbHj7PP
BOMdKPBdS51wlwcxS6i4833GRP34q9eW6qzUmmd+SlzNQykThAfcqnP91Ok/+9HC
fASS+ShPXZjMfr3EOlZYRcaCF87pnnNeF3K1csaLIZeWnw1cjwz2evAmGeF2gexQ
U2Ee72nMnXkfXuROgafZWorSawwr7MldsG980RBsF5+5kJytDiEjQmBanupIZGg0
vn8CDb5oexQyc+ZTCzwUP49jzvj6B1PtFlqPA9jN3dI5QvsqFxBV/HUyk6h2GY2G
5s0ytTbFOXuqKY+PqIqawQHTt2+DLY906mHXfbvHrmBEVvdQ2GzpUfne6tFtCMt5
y0zu/QVk/cDeGviUnd3LGamPfBtlSe5gCxC8jtnkkKTRMJDiXugldMJ4O4n6nmfU
dBXogCs6KWl3ramGkAgG4Zu4IIzS5rZWPr484Bee/bvOAfuxb22xUPqfo298Sok4
A1z1rKDBb6JhgrRHMIFjJLYUXpyq28VxRQQHA5LcQNqv3R8bcKUNvr17swNXzT56
KqwGE6egkzNbhfnxYxFLy9WBFxWev5xpsRrFRO8uuPxSArTYf0TghWoie+yNdzYr
jP4kFOCqHV+0AjNrg3KKOO+3qwBSfjgKa1JwaHs+o6RJbZAUKfi/zU40phhDPwg4
SgCHYiP8z75zdwobIlU8xZ2urRR7U9HInS7el3w60ldck7zQbOzAeJramlzmRc79
ZQI9uriGVBC2lSBVm8vTTRobFAnJIotqlmak/5hR0k+iNHpbawO9Hee8C24lMjlI
kfKYmd9B8G6iccTIhn10siIjMdabb47aezNYMUVCLGz0cAYcTgXV+gPk2+sbzxFN
tQbixTGGEhCzN6KuO0LjgjjmJoY6iXRJUbAqlMv4LbjeZE12q4VK45TbIImwS9dM
iCv5eoF9XpKeS40V3z0OYTSTajPpW7TqyIB/1n0iV/wESe7TuR1UCFDo0rkUQY/1
554wybK0q9n2bOLKA4ovl3YyxFtb7H6SvkzefNqUNytpWeiLmFzPEUZadooYlbgm
JOp19UdbvObWr/xDXT/jfEfNwNKgCzE5xbDRW8mMyX3Jq8PFwU27FbbMp6YqNj1f
nj2eREl8uWy1lGR4QAXqy8kb2pvT0WqqOXnzDlxLzTiSjQkKlMbaOvnzf3zmXpQW
HhnT7rgG1tJOLjWkFYUyH1kMGzcWFrZQ2JSQAFoxCS2wj2Bt+0MecHXLhnaC+Rjc
vOSwdwrtwMUU+j5joSeq75UZhRAVgU6uJ6eCz8duu0/dMu0EmAHVeqlg1K5xYqKM
n5j417600Z6GlrsfRCINtzsAy7a8bazwKup/WGCrXhZNO7+y8N4yMsML1N1QslSI
Y2dzNqLnmbQMV2u1c8wK8VcZ7wzfd69J53deYzv7WS8FEYUdAS9H/qA9+/3WVwEd
2WxhlYxD8nwewczbtFjRD3kbLGeoh3rd+IT3pY4eKOI0wYj9GrdsLJl6J8aN9UQG
Miz5u+bxFbZWsScJGnU6oiKSDqy8zmCst/MfykWzvaEu/mlPUjs/goRx4mrLewA3
51kTbVQ2vVO2hpXcbtntDThWSBpf9i2cILX+qYFwpvOSiSdpy3i7iIODN7qYBQpg
G7oJmK4zO0z+8ym1yOBSbiiz/P5Pkt6NpZx+V1BcC5ebNBV1fOoSfADHCE7OelwY
Twd+olPIUjwJu5hz4vv0wk46UFmyCZxhkJa4gQLZ/FezVzu2UU24iZ+NH40q/tQI
WEO4xL9ZL+j70HKJkVnws4Mm/D0lF73nnFGIlVkRx/xc1ADq47wBDekVnf4gDwR5
xHyAvv5EYbAJaxoRjovHRrpOFIHAIVYMljYa/mpb8lfra+VUg8wD4oiWjP1BCIwH
FbvQVITvKYObYcOrfJuJIAsPf0PS91rt1k3UEyLn/+5wHOvbl9m8f/ynio47aKEQ
Y0/ebGqv30WGpFnsXOWF/F7ENt2zhoiAk2MCTIZLj0YdVkQPsCJy/D4vQu4lPCLy
eQiOx0xicRqc9iq1So+eh47wl52wedAnBHDBFpNEhAsfMPCfvm9x5PBj1Z06hxxF
DKIL+ATESACz0xlo9fAB77SzHavHheBeWsiiXmSUA5yDNwnPdQaha6iZfzyAk3R8
B66MX5JNiM8CPKy293I/IksfOwAtV+Y4fi1hpJjkpqnG0m3S8+PawGXVaRyZGL/q
XSnSkH2RnTP2IFjI44VLMgXMvENLeN+lyrbPkC7YPTX10ZZL5CpVg2wNwkU3j0aS
mX00NmltmAbkzxce3SD9rQ2mXjB2wKRM///ZO62Ue7WLxGn9ojjGUTaAZ2YHFL18
SdUjCLCNKY9Jt3zIwLSgY3jUC/uVWtRccs5OpeUrbXDVcwOWiX4CmAFzUbnp8GCQ
SWXIsCEK4ZI6tvCdmNe/1GU+c30B1XKMDQwfcRtP9S/loSHGznvHAxJH7Xr1xsba
yXkHvgufBvUo+wuNmBJSlG2rrWc+27vslhqHUQ6tTDqVg+4DItHPYLcnMlO3pMHn
ucfegZMSeSyVPLy2TW+O/nc5zUDds31625lK1E657U/b9XOo2Lk9LKadK7PnFPaf
pxew/NNhzd/UjDB3BcCFFzxoJzcLdKB3lYKeSi9HqAcCi1DZqoFo29Ak60rXr3Nz
WN2IKGM/24qfTuVCkErdgCANXQJ1DG6ENBZ82o6aFcqMs5ubC5Q6ZHTZwQqhvqVB
OZ/e4VeX4gj/Mn3np3/CBiAqK4hVshXggcsr+V5wOi7HeZ2J6g5PdrNVI1iA2Hvm
hO+bM/UYJJbyy6oVR6Pc7CZS4CjOKyXXgb37t8j4WBm2hnnNVdYgB9fDKpqQLUX2
ww3n+iXFwJZJ7a6vBrZJ6fpA6Jx2TzKlj2ZDxK0zIrP17utrWcSfTtFLJ+H2RY/w
+0WhWi6vhpl39WBpKa3iAwTzNRV4iezhT0R4idYTnmzk32rNXUGsLW6JfAtU1eAZ
KG6oqDgdm6EfmbX55EdZ04sOpN9Ik+Q3uo0V9jpoEdlKhOa2YeUpt4M7oyuLEDqu
MI9MTfqnvFvlp5nugwswo6cGuEDQrvdzeyzFmDB4xJCl5NQ2hq2VszTruK8C6srm
QXiGk0SUUbgpt0jJ3xKu4KAwDHCOz9+WC2w7u4m7bjU6W8v9ds85h3aVIKPdbnJx
qAVdamid3AviTJxnh2RgSk8NDByTvAWPC/w138DdUH4aLHC8gB5H57g/ySORsThq
iT/ovUvWrL740frJmgJ2S/WCn70rMW26CkDFulcKdPGf+8HqwKcw1qNma3oO1/Ci
tFZ+y1PlOcaTvRkbEjmQWdcEfEhZihdHuVUHY8T6k/lUHQRQtZ9x8bveYWygQ6zE
0tLJs+VVkSLb5AWgzUPHJP+Mq8nx755WVF7vNu+esOUZNnXuliAvRkfRj9KnQyER
c5wAzLMtGfKSN0t3/peCt16pGmlEVhLW3UYahOhAjp4GqHIGNWXaNuAzl/dR/WCL
CFYaaH0FNk+gFm7/ml1JNNfTbL2jNyOoRYn+JGyVIZxbR43AM9TEafV37Nu0QPms
JLAy9kisJnFY7mkVeubL538FoARy5sCwolVzdUer04iZzXoawmwVfgxUJYjWOcvu
OsdHSTyaNJjyfUAiRjK5w6MdQ9pGqv9aXwd5v5Zp36QWPOIcyh+9Z/68gE97KWJg
XpHkuFox0c2Sleug+LA6uBrF4xgVw2QW+PRcWm20oHMf3X9Vbxrkqj5Inh9Vs4za
1tMHqCJ0bGKzdMWIPhnj8yVIu5S5M9jtzfuu1Chf8fBCraSEhyqnPv8WD+GxrEJ/
VV2zPtyVfFq0ygRCyg3ku3elOkPdIXc44DXCii5bk7JR0SUWpH6MiskpDVagrlRB
SDi01m2UqBPP5BbrWMzhTfELx41WX8LF4CClTjSmF5tERw0hJV+vcx3Qo+MOnFpy
CHTQ+qszDC9MWD4wv73e+opMNp7zjIQe7K8RCaoJouz6gu+TnYKxPuig62BCnRz+
IpRA2n4OjT/lvDS6azPBhu3U6uVE6RFXshHhOE9qXw+pgnyyrf5P1ww/Q2Bc/ZQx
RpxrOvk8fab+W7SGuKDYJnqNP53mxTshq6M2iKkStS43upcmcgg++sKhNzuPlh7U
8BUwB0y3G2KZdsrGmLUmd+q6pnxFypTdJ1ucmpxkSsWIJSwUkb3j9kOSGCbQPMro
46v3FubLuWjZ/JSe7mIVCwwLcjvQQwPzSH2XnUD3pC3Eq6yfWU8kmAcHIarzzsW0
ZGvNmabfrRhA9vCUzXn/DnTLCrBXoQahQV4txDjYVapdU5K280S9ujbazP5fYZA4
D0o7rRcF5tTReHPtn4jHow==
`pragma protect end_protected
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Ao7cWH3/D2aG1B4FXra6LkVB9mk4ARAKbtTS1Zgt6i58Crvs2KvtCtGjID3lFaUk
E+SUcO54B1FSOg1q370p5B/LAoqZ0fwMOP8wxqyrMyDuLfeHcBFGHeR0sQ/eD2vd
NlI7lvim6XopiIPzVEJ9jiEgAIg+QncOEPVN5sZ56+4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 17363     )
du1HJsGY5TGLffHhTzNn5jee4ciHBK2c2pUgOGCTdkhEbKJkdKxqwH63Uzksd2Ix
/a/RId8quevf82E9lVSkjkjfgUqepqeJQEPyZwX1A6sPM2j4Q2O7MYyMnteYAXz0
xGVeJClr72s4p/3acHpZbvfVBMFO5aUmNYR4JUKah9rEng685R32K327+FCcAvk2
BZo9myP+5s5LVcxcKbMqnOX/7INHIRRZ6xr9v8k2ethqUtqLE3HgABkVyOdV5k5h
+reul/K3tAnJpxUCl0uvHuvco41oIAPEREGqiBCseSZHYYEzB8JgIh9+X889WR1r
SnkAk7SmVklJRIN3i4zjiaEMcElRLmiFVgntTZqQpMiTXpW6kD1DC3/y8IBZD22i
gpze5VuuZLBX9XBCPXRHmYwHcrQd04DfcQoZ2md3q+7onykcDtUzMx9aE2Z/UJoW
4LJBLa1DuZX9HAn08nUn6rPvDJTqo+jdRQdzmJGCjodaircmtGva4RjirBpxneSX
DvkCLv6CSBI98jRFJ2UXboPPW0bw5EhpQq8gXx5M7yaqU/AOlhHz0M7yrP2S5h4n
4nyCCfxMJuVdxGxC3u9Nn9ihb+91TmvDJb/6P4NkTUOQXRZGlYBUncRtrG1LcYwh
DVnNjGrPXhph0L8QkKHUmmKnLwbw7ncD3KwgdFXUtYpBkQtvjBFbs2jTQJvkLhTa
D1p32XUsh6pTJgLti91os/N7xlfZD2idnhnP/PHpaGeobBEhZLKDKqkda4KWuNw2
yVRTxM9ItBo1bP1MfmnUNlXe0mZTuAjyijr+eOJMqDS2mkRhj5S6tBbdhOANNr92
Et8R7/dxfrNUFO50JKFWJYPh2vPzzb6xQq4HWu0VvopEDJkGe4rmp9ZxSDG2rgEc
NTQTgLuixbxNShG93bi6/yahRnDWQ7tFEeZOJlSEJxfiYwFx/Zw0Ra5XX5vTEp6/
XkuuqfMkFItdgp1/q0yZ1B9GBwfGHTfva5u8q0sWykHZM0u1X2tWkCBWAzdUCHGz
Q6Nd7X/IJD8G3mKyZVa3cEOcqrAc7GoNDwg3NKimSwFl05Ss0tDB+FpuoepuS86g
a39Qhc6v/McHKmtOi+7EGuLGTwXLKIsZyglL0ckRJzsA/0pgu6ocwHPrvMKfztnP
lYqNL6BMut66mT8G4dL3vXkeQKvXtSp2WPMJQB3lyFggxII1fKRfwCeempHeN4fJ
ObcsCFtS0yo62GLQgftMdfs5/70AEjDRG7NQAwbXa/2IswxxmCNzXeayGzZBv7VT
slbRNt5AeIq7OZ/2FIZadv1CeCSeW7jzupCsoZQn/jlMSaYoKUOpRvhmUEuhxjVt
8uQTZNmRo83Rfha35gQdmxQTYccQkvKaUF4GTMPnt11tiePt8FBL2VvkJCLmttAF
z4tvLS6UKeV7mdWVxYvLDYs0ZSKrDqupHCey3E0ygPwgpBlCrcbXdPmvoyZsYbNj
1jb7JvK6tnJhxmqwWKEablnzIp6c9G+/BC0YNNMQS5FxPNS5qN8qAT456I2xbl+3
Sa38peOj8mNKiOwpY4XPWjDVY7XuP4SqTyysQPgya/ZW1XPevRcDmIAwFdRxliSZ
dgpFd6MOft/+5ayTeoKSBIWeO2r0goXWC6c9K6/YcWFNP9GXRLVEE3TxofNtsapF
gqMzaoLxDvHuuTMudpTgVOl2+J8gNZ/aU4CIYvcpKro3fRFbh3GcEJnbJfa2fTur
ir9SL/DG8TTZpzPG5Y8/KVdmn0rmgwKrFXzoou33v71C4PFzQwQJBWCILiiF0wtD
1O6VVZogQkWCbeKgHHotkv16B59s6c6e/+Ho84WYVopgPvHDgBnzpIlknJnCVwu5
wv7S+e7t7edRiGYTt3xjz5OInZpb9CkrJ9JGH0BFz1ZDrcFYDfz8uSDWI9nAo+Vd
S4XqS41hOa9O1lqjNkEdeabHms7kDtn3DU+dwmyAZPYzt2yeg1hQzNgNKLjqPlwO
hlAZ4IcfpFiZEJbrtOjZGvF48w+ltFXXw3NOp8dyCXm3XNlT4Xpiw8KOEWLcGzfW
Ma6PRhyAs5Hki3/N09BKwU1QzRcyRfZEEb1RaAEWeT0Xmi8a+1mqt0DkRrIaz0Es
K3QgT+8yw305L/sANfdfEPTUTF0Gv8vlyXHPvNzWExs4vNSwEW8zVnC8tk+IY46M
LTD1pHvaEoRJSuVwCPiCqXpgxJ3XYJjoP4l9LEf2FYWtKGI4PAzPuU/SirYld+oB
JfIGfzzk/YdbXB1oBYmEXpf5cwF86dwahA/P/x2IFSmk6CDKQay0QVaFCctOHET4
eK+R8BliSrOD8YPYED4rqMQC/u0/muLShrr3EtgWWNgQ5/vzb3I7gnVSyEKbXWch
JRHkG6kLDZIKiw7IAN+C/1iayKlEfZdCeFbQF4mGFcr6GxHKJVZKrChBnQZWLVTs
60G2dHbdlyeary59B8oN0dC3YNVu09Te9KbHUtP9IfAhCcaxzkH5u9Wd4QTMHeCl
9paCRAXoaCBFcyHqfE06RAE26YpUt0ZG8aQBPEL2MSpSf1FEhRb62oeucPz1cOLz
EsPn5qi06v3kgvdJuQ3feEKQnTtYhAxkyAM+PweNqi1IwmI46IqXv/hyMG1dxwMx
Rd8B4O497Y66ZGDQAd+UDtb4StHF+VYjpxb5w9GaDm1OH2UapM+24T9bVFNkl2nY
9+fZoMoXpsDpllN66BIIaTfhwEjvHG09rF5Kc92bpSXw7M0Q8ymRybTtwfMhTLrW
hiwO6sN8Cn9wFKH3vYCyQ7OEHlpxv0RXsYAxCxlurhMxb1lC21iyWZIx20xFi1qS
aN6WAXNHk09Vv2G5OdOdrGhOjo6m92CgnxjA0rM0UHtoLNbB/uKnITk0ykewDUUf
14Lbp8ZsuBDHJOv3orknA0OGx1A/4eWxIVPnii8D4chZ6qGO3nGOKONMJE5FGqnD
db5gQsfYKYgvvCGpDcUuCLpLtL8aFMAmumHl38HpOGlbuucQQuFoi4lUbp4U0NaY
zJ0WbFbpPFN+JF2QQyUX/AgN3lLG6xi5beDxYj6siFJcYJ5k46sUvMVLcRD9rKM/
2a/hATCeIMJdp2cHaU2AWIVAPjnD/EcIgOulcMGVeA2D4M93nxP1m75/1yQz6Eha
ZiLMIaJatF0AM3O+bBzcOdpsYC+pm4NNN70PNG7jpzU7kktHrGX9HcTLYFRfDlcr
OPLIDrkm/Bi2jgdxP/Q5zBkeu4v3xTBYCZxiC91B31P25unXwUTsVRGQmWK9GDpZ
9Cc2owEh/MMgLEW8oQpl2vfM6lhG0fQLpiEWs/Aply55rrGE7PGB6A9cZEsG/6n4
GOhWFHz7sgQoMMeYCIms2qp75vlE0Bjw3UX0uwIZOI9Lq8PKFUqRaOqfLJsF4yJi
yUlHLO6YlWIQhUiKRkBrBMp8iJRIOiFpETML6fVXbZ/JjlJpc9l2XI5fkY5npgQT
Rbx++18jGMGUM7yH2y0gaZAakDfNPrnVZ1lhRdjyv+bzyUV2ivogNpD+t9y+lWSd
dS3+q1S1JB8AyqetYbhFRUh4wzJTgeKZFqHW2kIPeHDsVpDJ4k7p8haRYIxH82/g
`pragma protect end_protected
`endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
lxN1swUiEkIwz1jsFY9H2oPreC3qPxeA22Lb9xIE+sDKTegpFWHYaZnFfZxkvvBT
W5bOu5Pc8+EYtyis5TOX2iMt5t2s6d1BUAZfPyQ4J7MkuRdF9leH/IFOA/m6lU5e
mMAWayo6IghgAozijjI5RmGEd+HtEY5JiJskLp242mc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 17446     )
BrGmxuAio9r3WvMcEhMXfmK60Wzq6AlpTyFd+4IF2YOmhImyMbvgg1QAv+lt074/
OCdL0Cy8FZjJ45XLwoZu7c/L9Tui4SAIR3pbur/X0mjiEP1SygUNkgWIbcWh7EA0
`pragma protect end_protected
