

`ifndef GUARD_SVT_AXI_PORT_CONFIGURATION_SV
`define GUARD_SVT_AXI_PORT_CONFIGURATION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_system_configuration;
typedef class svt_axi_system_domain_item;
typedef class svt_axi_slave_addr_range;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UhZgkVHgMhDnDpYAD3Ent3d+5Xnc5oXdxX3KR9ehmfISpOvoV+uJE3Lpa3qcJ0Jd
FN/djJNlDfOpIwrZK4sSUo7iY/Bi8uJVniLHFTS17hDM+2q5cr3n8VfZRUjSAs6f
tSNLiJUISvh/pW+CtV6Do8LJnf4gE7TWfpOC5I7TtksLd1dscXyUDQ==
//pragma protect end_key_block
//pragma protect digest_block
KcYnzxjiAy0ZAch7dD0iWF0CYpU=
//pragma protect end_digest_block
//pragma protect data_block
9KFZvsmR+/h/J9DkjSQJOLqirKFPgt5sJA/QPb+z0e37LnlV8vwMsiJiUByPEnif
zAj3wonsW+cj+jyQJjgReZH/3Y6pDtwSO2CFrZKr/1JCJHHbADX/Ovqz06jiJFSk
lo/pR3valYXcM4Imf8DSFp1G2ivbA9p7P1auHMIYh9M6t/MOtbQlFGpQpjJBM8Bq
/RP1G6yH/3UnQdQX8UowQQVci/ZwZze3AsiQv68zUwWfnlptcoqpg0ouatCGHnNi
DegTl7oVjMYjERkEDXu2SfXevWHcl9bgUZkZXfxjjPYvYsMsubIbUKlbfGr0Lg6H
a5liDtiqv6KrzN9radrmjDDRDmBg2/9IYHT7vhZuGV10Rk3gtL1UDx4llR6bmAoa
hgnSYvJ79OrHBk9CRemqPd+bEOCIR8QmzhAxQUBaSVdF4aqJqlOLhqQ60ca7HT++
AvJyH1yDol5QD2QZUCYK0nfb4D7LzhmNfRcq2zgvM4lmljHR9Q/GjCvjDyLt0KHA
POrAqOY3ADxb5refmu7bSiyp3GzTrnfxv5TWpCZUyAcr1fFsEZOJ3JhvSSnMWVqt
HVXcjsSMB8pVnG9wImRwAYcF22zk46NrGJTSkJolFdUIHvvYonLUTL1mzvgLJ+dO
ysbvwwhqQbyMv+kcemA76HOYsqq1dDFn12GTp2CZdH+tODzLRR/jxn3V9E/OxisW
k++9L9QlhMrKn4LnSFWFz+3t403L8/fOvpqOxKGKQMAOTSc+Hyis7CY6fyoyhajh
5mb6iON2wLwJ7bMAbR+9gNpzbvzVncPI5y/W02lBk2ouVnIWKt/3P7Hf1vPfiZEf
hw9Vs2UNDGyngP1IUqjM9lLgMroAlIPPdnR28MNHsTnEQbAc+uRHSWQk8CqzFMiN
e0TXYixLP/mSJ2wHoI6c0fYAqf8kLEGm8hh3hwaFReZthH9CJazKmJP9PGS3g9ZJ
DTQhXa8mhQR+vBXI7YHYw6Qq9yPxkRgRvvWbxx9qLDu1PdkbJrvJ+QZujmITyaif
+K2golUCqHtjhwvxU1vta2dsN4ERRKJmJDL1xOdAwmK3ZYxFNnvUChLcFsLnA7+F
Eb7ZY7E5BwI2r5kk7qyNYoYPkIiUc7d43xfl2dun79Ypn4xKrEXWmomjNqQIbDfT
qenoVJ7AlbKtxaCTOuLVz/Z/5x412/ExY05TmkEZ5kQ+koN/kowIFmMNgTTRDNeV
7R666XHvxI0UTu6zvQcSil7kkaMjr2c9IC8MVhlpvxPfl2/+MsPZ39KGCE/YU45p
5/jFQS7jefEhO4xsjMTwc6VIoFA/PBk9GelwK9xbMdI8jYrHtmmSgxvvnKxLOmVo
EeRJDOkBoFtaN3iwgNwv16GQUt36gSKZEWv8XW4zYssALJXecLGO37dKORFZrgrc
lhWuKQZ2WLagD47bKYqqRAj0AOC1jzy8ZyLpjg4bkDNlzL339w0fSW9mpG3kYnyy
PBUiCUUHI65aLefMTUK5E1wIb0INDrhKFZZR4G/Uvtm2VM5HBW5zgAqS5SKqAMZ9
ohZJ44qbWOK+3c4gM3MSZglHf4ghIU8BcOGIg4Tp+Mg=
//pragma protect end_data_block
//pragma protect digest_block
f/LxhD1RCoZMjzpp33tj1WHB/wQ=
//pragma protect end_digest_block
//pragma protect end_protected

/**
    Port configuration class contains configuration information which is
    applicable to individual AXI master or slave components in the system component.
    Some of the important information provided by port configuration class is:
    - Active/Passive mode of the master/slave component 
    - Enable/disable protocol checks 
    - Enable/disable port level coverage 
    - Interface type (AXI3/AXI4/AXI4 Lite/AXI_ACE) 
    - Port configuration contains the virtual interface for the port
    .

  */
class svt_axi_port_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
`ifndef __SVDOC__
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if AXI_MASTER_IF;
  typedef virtual svt_axi_port_if AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if AXI_SLAVE_IF;
`endif // __SVDOC__
  typedef virtual svt_axi_stream_if AXI_PORT_STREAM_IF;
`endif
  
  /**
    @grouphdr axi_generic_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr axi3_4_config AXI3 and AXI4 configuration parameters
    This group contains attributes which are specific to AXI3 and AXI4 protocol
    */

  /**
    @grouphdr axi3_4_timeout_config Timeout values for AXI3 and AXI4
    This group contains attributes which are used to configure timeout values for AXI3 and AXI4 signals and transactions
    */

  /**
    @grouphdr ace_config ACE configuration parameters
    This group contains attributes which are specific to ACE protocol
    */
  
   /**
    @grouphdr ace5_config ACE5 configuration parameters
    This group contains attributes which are specific to ACE5 protocol 
    ARM-EPM-033524 Version 2.0
    */

  /**
    @grouphdr axi_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  /**
    @grouphdr axi_signal_idle_value Signal idle value configuration parameters
    This group contains attributes which are used to configure idle values of signals (except "Ready" signals) when "Valid" is low.
    */

  /**
    @grouphdr default_ready Default "Ready" signal value configuration parameters
    This group contains attributes which are specific to ACE protocol
    */

  /**
    @grouphdr axi3_signal_width AXI3 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI3 signals
    */

  /**
    @grouphdr axi4_signal_width AXI4 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 signals
    */

  /**
    @grouphdr ace_signal_width ACE signal width configuration parameters
    This group contains attributes which are used to configure signal width of ACE signals
    */

  /**
    @grouphdr axi4_stream_signal_width AXI4 Stream signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 Stream signals
    */

  /**
    @grouphdr master_slave_xact_association Configuration parameters required for master and slave transactions association
    This group contains attributes which are used to associate master transactions to slave transactions 
    */

  `ifdef SVT_VMM_TECHNOLOGY
  /**
    @grouphdr axi3_4_generator AXI3 and AXI4 generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for AXI3 and AXI4
    */

  /**
    @grouphdr ace_generator ACE generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for ACE
    */
  `endif

  /**
    @grouphdr protocol_analyzer Protocol Analyzer configuration parameters
    This group contains attributes which are used to enable and disable XML file generation for Protocol Analyzer
    */

  /**
    @grouphdr axi_performance_analysis Performance Analysis configuration parameters
    This group contains attributes which are used to monitor performance of a
    system based on measurement of latencies, throughput etc. The user sets the
    performance constraints through performance analysis configuration
    parameters and the VIP reports any violations on these constraints. The time
    unit for all these parameters is the simulation time unit. Performance
    metrics that involve aggregation of values over a time period are measured
    over time intervals specified using configuration parameter
    perf_recording_interval. Measurement of other performance parameters that do
    not require aggregation of values over a time period are not affected by
    this configuration parameter. VIP reports statistics for each performance
    metric for each time interval. Each performance parameter can be enabled or
    disabled at any time.  Monitoring of a performance parameter is disabled by
    passing a value of -1 to the parameter. Passing any other value enables the
    performance parameter for measurement. If a value other than -1 is supplied,
    it will take effect at the next time interval. If the performance
    configuration parameter values are changed during simulation, the new
    configuration will need to be passed to the VIP using the #reconfigure()
    method of the top level VIP component, for eg. #reconfigure() method of AXI
    System Env will need to be called if AXI system Env is used as top level
    component.
    */

  /**
    @grouphdr axi_qvn_config AXI QVN Configuration parameters
    This group contains attributes which are used to configure QVN features in a
    system.
    */

  /**
    @grouphdr axi_tlm_generic_payload TLM Generic Payload parameters
    This group contains attributes which are used to support TLM Generic Payload feature.
    */

  /**
    @grouphdr axi_traffic_profile Traffic profile related parameters
    This group contains attributes which are used to support traffic profiles.
    */

  /**
    * Enumerated type to specify idle state of signals. 
    */
  typedef enum {
    INACTIVE_CHAN_LOW_VAL  = `SVT_AXI_INACTIVE_CHAN_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_CHAN_HIGH_VAL = `SVT_AXI_INACTIVE_CHAN_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_CHAN_PREV_VAL = `SVT_AXI_INACTIVE_CHAN_PREV_VAL,   /**< Signal is
    driven to the previous value, ie, the value that it was driven to when the
    corresponding VALID signal was asserted. */
    INACTIVE_CHAN_X_VAL    = `SVT_AXI_INACTIVE_CHAN_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_CHAN_Z_VAL    = `SVT_AXI_INACTIVE_CHAN_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_CHAN_RAND_VAL = `SVT_AXI_INACTIVE_CHAN_RAND_VAL    /**< Signal is
    driven to a random value. */
  } idle_val_enum;

  /**
    * Enumerated type to specify inactive wdata bytes of signals. 
    */
  typedef enum {
    INACTIVE_WDATA_BYTE_LOW_VAL  = `SVT_AXI_INACTIVE_WDATA_BYTE_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_WDATA_BYTE_HIGH_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_WDATA_BYTE_X_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_WDATA_BYTE_Z_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_WDATA_BYTE_RAND_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_RAND_VAL,   /**< Signal is
    driven to a random value. */
    INACTIVE_WDATA_BYTE_UNCHANGED_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_UNCHANGED_VAL  /**<Signal is
    driven to initial value. */
  } wdata_val_enum;


  /** Enumerated types that identify the type of the AXI interface. */
  typedef enum {
    AXI3        = `SVT_AXI_INTERFACE_AXI3,
    AXI4        = `SVT_AXI_INTERFACE_AXI4,
    AXI4_LITE   = `SVT_AXI_INTERFACE_AXI4_LITE,
    AXI4_STREAM = `SVT_AXI_INTERFACE_AXI4_STREAM,
    AXI_ACE     = `SVT_AXI_INTERFACE_ACE,
    ACE_LITE    = `SVT_AXI_INTERFACE_ACE_LITE
  } axi_interface_type_enum;

  /** Enumerated types that identify the AXI interface category. */
  typedef enum {
     AXI_READ_WRITE = `SVT_AXI_READ_WRITE,
     AXI_READ_ONLY  = `SVT_AXI_READ_ONLY,
     AXI_WRITE_ONLY = `SVT_AXI_WRITE_ONLY
  } axi_interface_category_enum;

`ifdef SVT_ACE5_ENABLE

typedef enum {
  STANDARD = 0,
  BASIC = 1,
  NOT_SUPPORTED = 2 
 } mte_support_type_enum;

typedef enum {
  MPAM_9_1 = 0,
  MPAM_FALSE = 1
 } mpam_support_type_enum;

`endif
  /**
    * Enumerated typed for the port kind
    */
  typedef enum {
    AXI_MASTER = `SVT_AXI_MASTER,
    AXI_SLAVE  = `SVT_AXI_SLAVE,
    GP_MASTER = `SVT_AMBA_GP_MASTER,
    GP_SLAVE = `SVT_AMBA_GP_SLAVE
  } axi_port_kind_enum;

  /** @cond PRIVATE */
  /**
    * Enumerated type for the kind of inactivity period for throughput calculation
    */
  typedef enum {
    EXCLUDE_ALL = 0,
    EXCLUDE_BEGIN_END = 1
  } perf_inactivity_algorithm_type_enum;
  /** @endcond */

  /**
    * Enumerated type for enabling a particular version of ACE spec  
    */
  typedef enum {
     ACE_VERSION_1_0 = 0,
     ACE_VERSION_2_0 = 1
   } ace_version_enum;

  typedef enum {
    ALL_INTERFACE_TYPES = 0, /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE or ACE_LITE interface types. */
    AXI_ACE_ONLY = 1,        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE interface type. */ 
    ACE_LITE_ONLY = 2        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to ACE_LITE interface type. */ 
  } force_xact_to_cache_line_size_interface_type_enum; 

  /** @cond PRIVATE */
  /**
    * Enumerated typed for the memory kind
    */
  typedef enum {
    SV_BASED_SVT_MEM = `SVT_SV_BASED_SVT_MEM,
    C_BASED_SVT_MEM = `SVT_C_BASED_SVT_MEM
  } mem_type_enum;
  /** @endcond */

  typedef enum {
    RECOMMENDED_CACHE_LINE_STATE_CHANGE = `SVT_AXI_RECOMMENDED_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE
  } axi_cache_line_state_change_type_enum;

  /**
   * Enumerated type that indicates the reordering algorithm 
   * used for ordering the transactions or responses.
   */
  typedef enum {
    ROUND_ROBIN     = `SVT_AXI_REORDERING_ROUND_ROBIN, /**< Transactions will be 
    processed in the order they are received. */
    RANDOM      = `SVT_AXI_REORDERING_RANDOM, /**< Transactions will be 
    processed in any random order, irrespective of the order they are received. */
    PRIORITIZED = `SVT_AXI_REORDERING_PRIORITIZED /**< Transactions will be
    processed in a prioritized order. The priority of a transaction is known from
    the svt_axi_transaction::reordering_priority attribute of that transaction. */
  } reordering_algorithm_enum;

  /**
   * Enumerated type that indicates how the reordering depth 
   * of transactions moves.
   * 
   * Example:
   * Consider the read data reordering depth of 2; R1, R2, R3 and R4 are the read
   * transactions to be responded. The behavior for different types reordering depth
   * is as follows:
   * - STATIC:
   *   Once both R1 and R2 are complete, then only the reordering depth moves:
   *   {R1, R2} -- to --> {R3, R4}
   * - MOVING:
   *   If any of the R1 or R2 is complete, then the reordering depth moves. Suppose
   *   that R2 is complete before R1. Then the reordering depth window moves as:
   *   {R1, R2} -- to --> {R1, R3}
   * .
   */
  typedef enum {
    STATIC         = `SVT_REORDERING_WINDOW_STATIC, /**< The reordering depth moves
    when all transactions within the current reordering depth are complete. */
    MOVING         = `SVT_REORDERING_WINDOW_MOVING /**< A new transaction is considered
    for access to send read data as part of the given reordering depth when any transaction
    within the current reordering depth is complete. */
  } reordering_window_enum;
  
 /**
  * Name of the master as used in path coverage
  * This field can also be used to specify master specific
  * slave address mapping. Refer to the documentation of
  * svt_amba_addr_mapper for more details
  */
  string source_requester_name; 

  /**
   * This queue will hold the names of all the slaves, including non-AXI slaves, 
   * to which an AXI master can communicate.
   */
   svt_amba_addr_mapper::path_cov_dest_names_enum path_cov_slave_names[$];

  /**
   * Enumerated types that tells ERROR response handling policy for AXI Master and Slave.
   */
  typedef enum {
    NO_ERROR = 0,/**< When set to NO_ERROR,vip should not report an error on receiving decerr or slverr response. */
    ERROR_ON_SLVERR = 1,/**< When set to ERROR_ON_SLVERR,vip should report an error only on receiving slverr response. */
    ERROR_ON_DECERR = 2,/**< When set to ERROR_ON_DECERR,vip should report an error only on receiving decerr response. */
    ERROR_ON_BOTH = 3 /**< When set to ERROR_ON_BOTH,vip should report an error on receiving decerr or slverr response. */
  } error_response_policy_enum;

  /**
   * Enumerated type that defines the behaviour of the VIP during reset
   */
  typedef enum { 
    EXCLUDE_UNSTARTED_XACT = `SVT_AXI_EXCLUDE_UNSTARTED_XACT, /**< Only those transactions which have gone out on the interface are ABORTED. */
    RESET_ALL_XACT = `SVT_AXI_RESET_ALL_XACT /**< All transactions which have already started along with the ones which have not yet started but are present in the internal queue are ABORTED. */
  } reset_type_enum;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enumerated type that defines the generator source for slave responses
   */
  typedef enum { 
    NO_SOURCE    = `SVT_AXI_NO_SOURCE,           /**< No internal source. This generator_type is used by master component. This specifies that no internal source should be used, and user is expected to drive the master driver input channel. */
    ATOMIC_GEN   = `SVT_AXI_ATOMIC_GEN_SOURCE,   /**< Create an atomic generator. This generator_type is used by master component. This specifies the master component to use atomic generator. */
    SCENARIO_GEN = `SVT_AXI_SCENARIO_GEN_SOURCE,  /**< Create a scenario generator. This generator_type is used by master component. This specifies the master component to use scenario generator. */
    SIMPLE_RESPONSE_GEN = `SVT_AXI_SIMPLE_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_simple_callback is automatically registered with the slave response generator. This callback generates random response. */
    MEMORY_RESPONSE_GEN = `SVT_AXI_MEMORY_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_memory_callback is automatically registered with the slave response generator. This callback generates random response. In addition, this callback also reads data from slave built-in memory for read transactions, and writes data into slave built-in memory for write transactions. */
    USER_RESPONSE_GEN = `SVT_AXI_USER_RESPONSE_GEN_SOURCE /**< This generator_type is used by slave component. When this generator_type is specified, slave response callback is not automatically registered with the slave component. The user is expected to extend from svt_axi_slave_response_gen_callback, implement the generate_response callback method, and register the callback with the slave response generator. */
  } generator_type_enum;

  /**
   * Enumerated type that defines the generator source for snoop responses
   */
  typedef enum { 
    CACHE_SNOOP_RESPONSE_GEN = `SVT_AXI_CACHE_SNOOP_RESPONSE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, a callback of type #svt_axi_master_snoop_response_gen_cache_callback is automatically registered with the master component. This callback generates random snoop response based on the cache line status. */
    USER_SNOOP_RESPONSE_GEN = `SVT_AXI_USER_SNOOP_RESPONSE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, snoop response callback is not automatically registered with the master component. The user is expected to extend from #svt_axi_master_snoop_response_gen_callback, implement the generate_snoop_response callback method, and register the callback with the snoop response generator. */
  } snoop_response_generator_type_enum;

  /**
   * Enumerated type that defines the barrier transaction association approach
   */
  typedef enum { 
    RANDOM_ASSOCIATION = `SVT_AXI_RANDOM_BARRIER_XACT_ASSOCIATION, /**< This approach type is used by master component, when the #axi_interface_type is AXI_ACE. When this approach is specified, a callback of type #associate_xact_with_barrier_pair_xact() is automatically registered with the master component. This callback associates barrier transaction with normal coherent transaction in a random manner. */
    USER_DEFINED_ASSOCIATION = `SVT_AXI_USER_DEFINED_BARRIER_XACT_ASSOCIATION /**< This approach type is used by master component. When this approach is specified, the callback is not automatically registered with the master component. The user is expected to extend from
#associate_xact_with_barrier_pair_xact, implement the association of barrier transaction with normal coherent transaction */
  } barrier_association_type_enum;

  /**
   * Enumerated type that defines the generator source for DVM complete transactions
   */
  typedef enum { 
    AUTO_DVM_COMPLETE_GEN = `SVT_AXI_AUTO_DVM_COMPLETE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, master automatically generates a DVM Complete transaction, after receiving a DVM Sync transaction. The delay between reception of DVM Sync and transmission of DVM Complete is determined by random member dvm_complete_delay*/
    USER_DVM_COMPLETE_GEN = `SVT_AXI_USER_DVM_COMPLETE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, user will need implement callback method svt_axi_master_snoop_response_gen_callback::dvm_complete_gen. The user can program the delay  dvm_complete_delay in the callback method. */
  } dvm_complete_generator_type_enum;

`endif

  /**
   * Enumerated type that defines the snoop response mode during memory update transactions
   */
  typedef enum { 
    SUSPEND_SNOOP_DURING_MEM_UPDATE = 0, /**< Master suspends incoming snoop request if memory update transaction is found in the buffer, or is active at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    SUSPEND_SNOOP_DURING_MEM_UPDATE_IN_PROGRESS = 1, /**< Master suspends incoming snoop request if memory update transaction is found to be active (addres/data phase started or about to start in current clock) at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    RESPOND_SNOOP_DURING_MEM_UPDATE = 2, /**< Master doesn't suspend incoming snoop request even if memory update transaction is found to be active at the time of receiving snoop request. Instead it responds to the snoop request with allowed snoop response while memory update transaction is in progress.*/ 
    EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE = 3  /**< Master either suspends incoming snoop request or respond to the snoop request while memory update transaction is in progress in a random manner.*/ 
  } snoop_response_mode_during_mem_update_type_enum;

  /**
    * 
    */
  typedef enum {
    SNOOP_RESP_DATA_TRANSFER_USING_CDDATA = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_CDDATA, /**<Transfers cache data of dirty line using CDDATA channel */
    SNOOP_RESP_DATA_TRANSFER_USING_WB_WC = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_WB_WC /**<Transfers cache data of dirty line using WRITEBACK or WRITECLEAN */
  } snoop_response_data_transfer_mode_enum;

  /** enum description for various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE */
  typedef enum {
    NONSHAREABLE_XACT_FULL_ADDRESS_SPACE = 0, /**<allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE = 1, /**<allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE = 2, /**<allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE = 3 /**<allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
  } nonshareable_xact_address_range_in_systemshareable_mode_enum;
  typedef enum {
    STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 0,
    DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 1,
    CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 2 
  } source_master_id_xmit_to_slaves_type_enum;

  typedef enum {
    FALSE = 0,
    ODD_PARITY_BYTE_DATA = 1,
    ODD_PARITY_BYTE_ALL = 2
  } check_type_enum;

  /**
   * Enumerated type that defines the modifiable and non modifiable cache types
   */
  typedef enum {
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK = 0,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK = 1,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_DISABLE_CHECK = 2
  } master_slave_xact_association_cache_prot_check_enum;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
`ifndef __SVDOC__
  /** Port interface */
  AXI_MASTER_IF master_if;
  AXI_SLAVE_IF slave_if;
  AXI_PORT_STREAM_IF port_stream_if;
`endif

  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to the master/slave port corresponding
    * to this port configuration. This ID must be unique across
    * all masters/slaves of the AXI system configuration to which
    * this port belongs. A master and a slave may share the same
    * port_id, but two masters or two slaves cannot share the 
    * same port_id. If not assigned by the user, it is auto
    * assigned by the VIP. 
    */ 
  int port_id;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Name of this port. This is used in transaction short display
    * to identify the instance. This is copied over from 'inst'
    * attribute.  
    */
 local string port_name;
  /** @endcond */
  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to master/slave port corresponding to this port
    * configuration. This ID must be unique across all AMBA components
    * instantiated in the testbench.  This is currently applicable only when the AMBA
    * system monitor is used and is configured using a configuration plain text
    * file (as opposed to a SystemVerilog code that sets the configuration). 
    */
  int amba_system_port_id = -1;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether output signals from master/slave IFs should be
    * initialized to 0 asynchronously at 0 simulation time. 
    * - 1: Intializes output signals from master/slave IFs to 0 
    *      asynchronously at 0 simulation time.
    * - 0: Initializes output signals from master/slave IFs to Z
    *      synchronously at 0 simulation time.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit initialize_output_signals_at_start = 1'b0;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether clock should be disconnected to this agent. 
    * - 1: clock will be connected to this agent from the testbench, 
    *      based on the svt_axi_system_configuration::common_clock_mode.
    * - 0: clock will not be connected to this agent from the testbench.
    *      Used to disable the agent as per the test requirement.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit clock_enable = 1'b1;

  /**
    * @groupname axi_generic_config
    * Handle to the system configuration object
    */
  svt_axi_system_configuration sys_cfg;

  /**
    * @groupname axi_addr_map
    * Applicable only to slave VIP
    * Address map for this slave 
    * Must be used only if the svt_axi_system_env and svt_axi_system_configuration is not used.
    * Typically used in an environment where only one slave VIP is instantiated.
    */
  svt_axi_slave_addr_range slave_addr_ranges[];

  /**
    * @groupname axi_addr_map
    * Address map that maps global address to a local address at destination
    * Typically applicable to slave components
    * Applicable only if svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper dest_addr_mappers[];

  /**
    * @groupname axi_addr_map
    * Address map that maps a local address to a global address at a source
    * Typically applicable to master components. However, it can be applicable to
    * a slave component if that is connected downstream through another interconnect/bridge to
    * components which are further downstream. Applicable only if
    * svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper source_addr_mappers[];

  /**
    * @groupname axi_generic_config
    * Indicates if WID must be driven for AXI4, AXI_ACE,ACE_LITE,AXI4_LITE interfaces 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit  wid_for_non_axi3_enable = 0;

  /** 
    * @groupname axi_generic_config
    * Field for updating slave memory in request order
    * When set to 1, updates slave memory in request order that is  even though response
    * is received out of order, memory will still be updated in request order at the last
    * data phase. 
    * Default value is 0.
    * Configuration type: Static
    * Applicable only to SLAVE
    */ 
    int update_memory_in_request_order = 0;

    /**
    * @groupname axi_generic_config
    * Indicates that the monitor will check that recommended number of transactions are used      in the locked sequence 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit check_recommended_xact_length_for_locked_sequence = 0;
   
    /**
      * @groupname axi_generic_config
      * Indicates if X/Z checks and signal stability checks must be enabled
      * These are low level checks performed every clock and have a performance overhead
      * Often, these checks are useful only during integration phase. These can be
      * switched off after integration to get better performance.
      * These checks are automatically disabled if SVT_AXI3_4_PERF_MODE is set
      */
    bit per_clock_cycle_signal_checks_enable = 1;
 

  /**
    * @groupname axi_generic_config
    * If set to svt_axi_port_configuration::RESET_ALL_XACT,all transactions which have
    * already started along with the ones which have not yet started but are
    * present in the internal queue are ABORTED.
    * If set to svt_axi_port_configuration::EXCLUDE_UNSTARTED_XACT,only those transactions
    * which have gone out on the interface will be ABORTED.
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode because in passive mode
    * or for the slave all transactions which are in the queue are already started
    */
    reset_type_enum reset_type = `SVT_AXI_RESET_TYPE;


  /**
   * @groupname axi3_4_config
   * Indicates the way VIP reports error on receiving SLVERR or DECERR read or write response.
   * If set to svt_axi_port_configuration::NO_ERROR,vip doesn't report any error on receiving decerr
   * or slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_SLVERR,vip reports error only on receiving 
   * slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_DECERR,vip reports error only on receiving 
   * decerr response.
   * If set to svt_axi_port_configuration::ERROR_ON_BOTH,vip reports error on receiving 
   * decerr or slverr response.
   * Configuration type: Static
   *
   * This is applicable to Master in both active and passive mode and to slave only in Passive mode.
   * The default enum type of error_response_policy is NO_ERROR and is user configurable.
   */
   error_response_policy_enum error_response_policy = NO_ERROR;


  /**
    * @groupname axi_generic_config
    * Indicates if VIP would use separate address spaces for each tagged attribute. This simply means that,
    * if a coherent master or interconnect or a slave attached to such system, recieves both secure and non-secure
    * transactions then both transactions will operate on completely separate address spaces and result of one transaction
    * will not be visible to the other.
    *
    * Slave for which separate secure & non-secure address space is enabled i.e. bit [0] is set to '1', it will accept both secure
    * and non-secure transactions targeted for the same address. However, while updating memory it will use tagged address i.e. 
    * address attribute, in this case security bit, will be appended to the original address as the MSB bits.
    *
    * Slave for which separate secure & non-secure address space is disabled i.e. bit [0] is set to '0' but, configured with secured
    * regions i.e. addr_attribute[0] is set to '1' in svt_axi_slave_addr_range class via task /#set_addr_range() in system configuration
    * then it will accept only secure transactions for secure regions and all transactions for non-secure regions. 
    * With this configuration slave will use orginal address while updating memory and will not use tagged address. Hence, secure and
    * non-secure transactions to the same address will affect each other, if targeted to non-secure regions. However, if it is targeted
    * to secure regions then only secure transations will be able to update memory and access for non-secure transactions will be declined as if address doesn't exist.
    *
    * Slaves can be configured with secure region by calling /#set_addr_range(<start_addr>,<end_addr>,<addres_attribute, ex: 1 [secured]>)
    *
    * [0] => represents separate address spaces for secure and non-secure attribute if set to '1'
    * [\`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:1] => RESERVED and should be set to 0
    *
    * Configuration type: Static
    * Applicable only to MASTER 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 0;
`else    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 1;
`endif    
    
  /**
    * @groupname axi_generic_config
    * If set to '0' then Master VIP will not drive overlapped coherent transactions on Read and Write
    * channel at the same time. WRITE transactions received by the sequencer will be blocked from being
    * sent on the interface if there is another READ transaction to an overlapping address which is 
    * already in progress. The same is true if a READ transaction is received from sequencer and a WRITE
    * transaction is in progress
    * Example: ReadShared started at 1000 ns and WriteBack received from sequencer at 1200 ns when 
    *          ReadShared is still active. At this point Master VIP will block WriteBack until ReadShared
    * is finished on the Read channel.
    *
    * If set to '1' then Master VIP will drive coherent transactions on Read and Write
    * channel as it receives from the sequencer as per other coherent rules. It will not
    * block as mentioned above. 
    * Certain scenarios that involve a store on the read channel sent out
    * speculatively while a WRITEBACK/WRITECLEAN to the same cacheline is in
    * progress require that this parameter is set to 0 so that cache states
    * reflect correctly. 
    * If snoop_response_data_transfer_mode is set to
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, this parameter must be set to 1 to
    * facilitate the transfer of snoop data on the write channel without
    * getting blocked.
    *
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode 
    */
    bit allow_overlapped_read_and_write_channel_coherent_transactions = 0;    
   
   /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP can drive random snoop response for
    * WasUnique (BRRESP[4]) even if the snoop_initial_cache_line_state is in 
    * UNIQUE state.
    * If set to '0' the Master VIP must set WasUnique (BRRESP[4]) to 1 if
    * the snoop_initial_cache_line_state is UNIQUE.
    */ 
    bit allow_was_unique_zero_in_unique_state = 1; 
   
   /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP will allow burst_size to be less than
    * data_width for Atomic transaction.
    * If set to '0' then Master VIP will throw an is_valid error when burst_size 
    * is less than data_width for Atomic transaction.
    * This is only applicable for multibeat atomic transactions. 
    */
    bit allow_multibeat_atomic_transactions_to_be_less_than_data_width = 0;   
    /** @endcond */

   /**
    * @groupname axi_generic_config
    * This is applicable only when interconnect VIP is used, this is
    * applicable for all transactions. 
    * So if set to 1, then the interconnect VIP will always update dirty data into main memory 
    * if it receives dirty data from snoops corresponding to a transaction from this port
    */
    bit memory_update_for_pass_dirty_enable = 0;
 
   /**
    * @groupname axi_generic_config
    * This is applicable only when interface_type is AXI3 or AXI4
    * If set to 1 and axi_interface_type is AXI3/AXI4, system monitor will update
    * the port_configuration member axi_interface_type as ACE_LITE .
    * In addition to that system monitor will update svt_axi_transaction::xact_type as COHERENT.
    */

    bit is_downstream_coherent = 1'b0;

  /** @cond PRIVATE */
  /** Helper attribute for specifying solve order */
  local rand bit primary_props;

  /** holds total number of enabled tagged address space attributes */
  local int      num_enabled_tagged_addr_attributes = 0;

  /** Supports four state memory
   *  Default value is set as 0
   *  If set as 1 supports 4 state memory.
   */

  bit is_4state = 1'b0;
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  /** 
   * @groupname axi3_4_generator
   * The source for the stimulus that is connected to the transactor.
   *
   * Configuration type: Static
   */
  generator_type_enum generator_type = SCENARIO_GEN;

  /**
   * @groupname ace_generator
   * The source type for snoop response generation.
   *
   * Configuration type: Static
   */
  snoop_response_generator_type_enum snoop_response_generator_type = CACHE_SNOOP_RESPONSE_GEN;

  /**
   * @groupname ace_config
   * Defines how a transaction is associated with a barrier transaction pair.
   *
   * Configuration type: Static
   */
  barrier_association_type_enum barrier_association_type = RANDOM_ASSOCIATION;

  /** 
    * @groupname ace_generator
    * Defines how DVM complete transactions need to be generated.
    *
    * Configuration type: Static
    */
  dvm_complete_generator_type_enum dvm_complete_generator_type = AUTO_DVM_COMPLETE_GEN;

  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_scenarios = -1;

  /**
    * @groupname axi_generic_config
    * The number of instances that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_insts = -1;

  // ACE
  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the snoop_generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_scenarios = -1;

  /** 
    * @groupname axi_generic_config
    * The number of instances that the snoop generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_insts = -1;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_LOW verbosity.
    */
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_LOW verbosity.
    */
`else
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in DEBUG_SEV.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in NORMAL_SEV.
    */
`endif
  bit silent_mode  = 0;

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`elsif SVT_OVM_TECHNOLOGY
  /** 
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and 
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`else
  /**
    * @groupname axi_generic_config
    * Specifies if the group is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables driver, generator and
    * monitor in the group component. 
    * - 0: Configures component in passive mode. Enables only the monitor in the group component.
    * - Configuration type: Static
    * .
    */
`endif
  bit is_active = 1;
  
  /** @cond PRIVATE */
  /** xml_writer handle of the agent */
  svt_xml_writer xml_writer = null;
  /** @endcond */


  /** 
    * @groupname axi_generic_config
    * The AXI interface type that is being modelled. Please note that interface
    * type AXI_STREAM is not yet supported.
    * Configuration type: Static
    */
  rand axi_interface_type_enum axi_interface_type = AXI3;

  /** 
    * @groupname axi3_4_config
    * The AXI4 interface category (read-only, write-only, read-write) of this interface. 
    * Configuration type: Static
    */ 
  rand axi_interface_category_enum axi_interface_category = AXI_READ_WRITE;

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a master or a slave. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is of kind master or slave.
    */ 
  axi_port_kind_enum axi_port_kind = AXI_MASTER;

  /**
    * Specifies the impact of svt_axi_transaction::force_xact_to_cache_line_size 
    * based on the axi_interface_type. 
    * 
    * Applicable only for ACTIVE master.
    */
  force_xact_to_cache_line_size_interface_type_enum force_xact_to_cache_line_size_interface_type = ALL_INTERFACE_TYPES;

 /** 
   * @groupname ace5_config
   * Indicates supported version  of ACE specefication by AMBA AXI_ACE VIP
   * Default value of this parameter is ace_version_1_0.User need to set this parameter if they wish to
   * to use new ACE spec which is ACE spec version 2.0
   * Configuration type:static
   */
   ace_version_enum ace_version = ACE_VERSION_1_0;

/** 
   * @groupname ace5_config
   * Indicates cache stashing feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cache_stashing_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates if trace signal feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit trace_tag_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates whether the trace tag value will be directly reflected in the response packet or spawned packets generated in response to the received packet.
   * when set to 1: The trace_tag value will be directly mapped to the associated response and spawned packets, irrespective of trace_tag value being 0 or 1 in the request.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 and svt_axi_port_configuration::trace_tag_enable is set to 1.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit loopback_trace_tag_enable = 0;

`ifdef SVT_ACE5_ENABLE 
/** 
   * @groupname ace5_config
   * Indicates if atomic transactions feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit atomic_transactions_enable = 0;


 /** 
   * @groupname ace5_config
   * Indicates if write_with_cmo feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit write_plus_cmo_enable = 0;
 
 /** 
   * @groupname ace5_config
   * Indicates if cmo transactions can be sent on the write channel.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cmo_on_write_enable = 0;

 /**@groupname ace5_config
   * Specifies the number of outstanding Atomic transactions a port can support.<br>
   * This is applicable only for ACE5 ports with atomic_transactions_enable set to 1.<br>
   * The Atomic transactions include:
   * - AtomicStore
   * - AtomicLoad
   * - AtomicSwap
   * - AtomicCompare
   * .
   * MASTER:
   * If the number of outstanding atomic transactions is equal to this
   * number, the slave will refrain from initiating any new 
   * transactions until the number of outstanding write transactions
   * is less than this parameter.<br>
   * SLAVE:
   * If the number of outstanding transactions is equal to 
   * this number, the slave will not assert ARREADY/AWREADY
   * until the number of outstanding transactions becomes less
   * than this parameter. 
   * <br>
   * This parameter must be set if #num_outstanding_xact = -1.
   * This parameter must not be set if #num_outstanding_xact is not set to -1.
   * - <b>Default val:</b> -1
   * - <b>min val:</b> 1
   * - <b>max val:</b> Value defined by macro \`SVT_AXI_MAX_NUM_OUTSTANDING_XACT.
   * - <b>type:</b> Static
   * .
   */
  rand int num_outstanding_atomic_xact = 1;

 /** 
   * @groupname ace5_config
   * Indicates if Memory Partitioning and Monitoring (MPAM) feature is supported.
   * It can be set to either of two values below:
   *    enable_mpam = svt_axi_port_configuration:FALSE
   *  When set to FALSE, MPAM is not supported on the interface.
   *    enable_mpam = svt_axi_port_configuration:MPAM_9_1
   *  When set to MPAM_9_1, MPAM is supported on the interface with mpam_partid_width=9 and mpam_perfmongroup_width=1. 
   *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * - Default value:FALSE, is controlled through user re-definable macro `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM.
   * .
   */
   mpam_support_type_enum enable_mpam = `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Partition identifier.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_partid_width = 9;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Performance monitor group.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_perfmongroup_width = 1;

`endif
  /**
   * @groupname ace5_config
   * If set to 1, it will enable the master component to support deallocating transactions.
   * By default, the value of this parameter is 0. This means it can not support deallocating
   * transactions and any READONCEMAKEINVALID or READONCECLEANINVALID transaction initiated
   * from this master component will be converted to READONCE transaction.
   *
   * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * and svt_axi_port_configuration::axi_interface_type is set to ACE_LITE
   * Configuration type:static
   */
   bit deallocating_xacts_enable = 0;



  /** 
   * @groupname ace5_config
   * Indicates address translation feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit addr_translation_enable = 0; 

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a interconnect VIP port or not. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is a port of interconnect VIP or not.
    * .
    */  
  bit is_ic_port = 0;
  
 /**
   * @groupname axi_generic_config
   * Indicates if the port_monitor protocol check max_num_outstanding_xacts_check 
   * is enabled or not .The max_num_outstanding_xacts_check checks that AXI master and AXI slave 
   * are not exceeding the user configured maximum number of outstanding transactions (#num_outstanding_xact).   
   * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
   * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for read and write transactions respectively.
   */
  bit max_num_outstanding_xacts_check_enable =0; 
 
  /** @groupname axi_generic_config
    * Disable the association between slave read transaction and master partial write transaction.
    * This covers the specefic scenario when master partial write transaction is split into
    * slave read transaction followed by a slave write transaction by the ICN.
    * If set to 1 association between master write transaction and slave read transaction is done by the system monitor.
    * If set to 0 association between master write transaction and slave read transaction is not done by the system monitor.
    */
  bit partial_write_to_slave_read_and_write_association_enable = 0;
 
 /**
   * @groupname axi_generic_config
   * Indicates if this port is interleaved based on address to be accessed by this port
   */
  bit port_interleaving_enable =0;  
 
/** Indicates the port interleaving boundary. The value must be in form of bytes.
  * For example if interleaving szie is 64 . It means interleaving boundary os 64 bytes.
  * This port will access address locations based on interleaving size.
  * Default value is set as 64.
  * Applicable if the port_interleaving_enable is set to 1 for this port.
  */
  int port_interleaving_size = 64;

/** Indicates the group id of all the ports participating in one interleaving scheme
  * All the ports which are in the same interleave group must be configured to have same 
  * port_interleave_group_id
  * Default is set to -1 . 
  * Applicable if the port_interleaving_enable is set to 1.
  * Its value must be unique across master and slaves .All the port_ids having same port_interleaving_group_id
  * must be contigous.
  */
  int port_interleaving_group_id = -1;

/** Indcates that DVM transactions will be sent form this port of corresponding port interleaving group
  * This port will not take part in port interleaving for DVM transactions 
  * Applicable if port_interleaving_enable is set to 1.
  */
  bit dvm_sent_from_interleaved_port = 0;

/**Indicates that non coherent device traffic will be sent from this port
  * of corresponding port interleaving group.
  * This port will not take part in port interleaving for device traffic
  * as Device transaction addresses are not interleaved.
  * Applicable only when the port_interleaving_enable is set to 1.
  */ 
  bit device_xact_sent_from_interleaved_port =0;

/**  Indicates the order of this port in a port interleaving scheme.
  *  For example : If the port is 3rd in a group of 4 ports .If port_interleaving_size of the group is 512 bytes
  *  This port will have access to addresses with addr[10:9] == 3.
  *  This parameter determines which address bits to look for an interleaved port.
  *  Default value of this is set to 0 
  */
   int port_interleaving_index = 0;

  /**
   * @groupname axi_generic_config
   * Enables port inteleaving for this port for the device type xact.
   * The port configuration parameter device_xact_sent_from_interleaved_port
   * is not applicable if this bit is set to 1.
   * If this bit is set to 1, the device type transaction is interleaved like 
   * any non-dvm transaction.
   */
  bit port_interleaving_for_device_xact_enable = 0;

  /**
    * Indicates if this port  supports the setting of Poison field. <br>
    * - Default value: 0.
    * .
    */
  bit poison_enable = 1'b0;

   /** 
    * @groupname axi_generic_config
    * Indicates if the transactions on this port must be processed by the axi
    * system monitor. This configuration is applicable only to the
    * 'system_monitor' of the instance of svt_axi_system_env within which the
    * component corresponding to this port configuration is instantiated.
    * It is not used in the AMBA system monitor instantiated in an instance of
    * svt_amba_system_env (system env used when multiple AMBA protocols are
    * used)
    */ 
  bit connect_to_axi_system_monitor = 1;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Indicates that, if this bit is set to '1' then user needs to externally push
    * coherent and snoop master transactions and slave transactions into the port monitors. 
    * port monitor will not automatically sample it's related interface and hence will not
    * create corresponding transactions and instead will use the user provided transaction handle
    * externally pushed into the monitor.
    */ 
  bit use_external_port_monitor = 0;
  /** @endcond */

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates a tlm_generic_payload_sequencer sequencer capable
    * of generating UVM TLM Generic Payload transactions and connects the
    * master sequencer to it.  The master sequencer starts a layering sequence that gets
    * transactions from the tlm_generic_payload_sequencer, converts them to (one or more) AXI
    * transaction(s) and sends them to the driver.
    * Snoop requests are still fulfilled by the svt_axi_master_snoop_sequencer.
    * 
    * AXI transactions observed by the agent
    * are also made available as TLM GP transactions through the
    * tlm_generic_payload_observed_port in the monitor. Note that the TLM GP
    * transactions issued through the analysis port may not match one to one with GP
    * sequence items created by the tlm_generic_payload_sequencer because the
    * GP sequence items may have to be mapped
    * to multiple AXI transactions according to protocol requirements. The
    * TLM GP that is available through the tlm_generic_payload_observed_port of
    * the monitor is a direct mapping of the observed AXI transactions converted to a TLM GP.
    * No attempt is made to re-assemble a set of AXI transaction into a larger TLM GP.
    * 
    * The layering sequence that converts the TLM GP to AXI transactions is the
    * svt_axi_tlm_gp_to_axi_sequence and is available at
    * $DESIGNWAREHOME/vip/svt/amba_svt/<ver>/axi_master_agent_svt/sverilog/src/vcs/svt_axi_tlm_gp_sequence_collection.svp 
    * Transactions created by the layering sequence are of type
    * cust_svt_tlm_gp_to_axi_master_transaction. Any user constraints specific
    * to AXI must be provided in a class extended from this class.
    * 
    * In passive mode, observed AXI transactions are made available as TLM GP
    * transactions through the tlm_generic_payload_observed_port in the
    * monitor.
    */
  bit use_tlm_generic_payload = 0;

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates an AMBA-PV-compatible socket that can be used to
    * connect AXI Master VIP component to an AMBA-PV master model. 
    * 
    * Enabling this functionality causes the instantiation of socket b_fwd of
    * type uvm_tlm_b_target_socket, and socket b_snoop of type
    * uvm_tlm_b_initiator_socket, in class svt_axi_master_agent.

    * Generic payload transactions received through the forward b_fwd interface
    * are executed on the tlm_generic_payload_sequencer in the agent.

    * When this option is set, the svt_axi_ace_snoop_request_to_tlm_gp_sequence
    * reactive sequence is started on the AXI VIP master snoop sequencer. Snoop
    * transaction requests received by the AXI VIP master snoop sequencer are translated to
    * equivalent tlm_generic_payload transactions with the
    * #svt_amba_pv_extension attached. The extended Generic Payload transactions
    * are then sent to the AMBA-PV master model via the backward b_snoop interface.
    * The receive response from AMBA-PV master model is then interpreted to
    * complete the snoop transaction request and executed on the AXI VIP master snoop
    * sequencer.
    * 
    * Should the AXI VIP master fulfill the snoop requests natively (i.e. the
    * default behavior when this option is not set), the snoop response sequence
    * should be restored to the default using:
    * 
    * <code>
    * uvm_config_db#(uvm_object_wrapper)::set(this, "master[0].snoop_sequencer.run_phase", "default_sequence",
    *                                         /#svt_axi_ace_master_snoop_response_sequence::type_id::/#get());
    * </code>
    * 
    * When this option is set, it implies that #use_tlm_generic_payload is also set, whether
    * it actually is or not.
    */
  bit use_pv_socket = 0;

 /** Enables the UVM REG feature of the AXI agent.  
   * Applicable only when svt_axi_port_configuration::axi_interface_type is AXI3.
   * <b>type:</b> Static 
   */
  bit uvm_reg_enable = 0;

 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables checking of wdata/tdata only on valid byte lanes based on wstrb/tstrb. 
    * In a disabled state, whole wdata/tdata as seen on the bus will be considered.
    * <b>type:</b> Dynamic 
    */
  bit check_valid_data_bytes_only_enable = 1;

  /**
    * @groupname axi3_4_timeout_config
    * A timer which is started when a transaction starts. If the transaction
    * does not complete by the set time, an error is repoted. The timer is
    * incremented by 1 every clock and is reset when the transaction ends. 
    * If set to 0, the timer is not started
    */
  int xact_inactivity_timeout = 0;

 /**
   * @groupname ace_config 
   * If this attribute is enabled it will allow snoop response data_transfer bit for
   * MAKEINVALID  transaction to be set as 1. This behaviour is permitted by protocol
   * but it is not expected snoop response for MAKEINVALID 
 */
  bit  data_transfer_for_makeinvalid_snoop_enable =0;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /** 
   * log_base_2 of \`SVT_AXI_MAX_DATA_WIDTH. 
   * Used only as a helper attribute to randomize data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_data_width;
 
  /** 
   * log_base_2 of \`SVT_AXI_ACE_SNOOP_DATA_WIDTH. 
   * Used only as a helper attribute to randomize snoop_data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_snoop_data_width; 

  /** 
   * log_base_2 of \`SVT_AXI_MAX_CACHE_LINE_SIZE. 
   * Used only as a helper attribute to randomize cache_line_size.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_cache_line_size;

  /**
    * Indicates if the address range of the slave component
    * has been set
    */
  bit is_slave_addr_range_set = 0;

  /**
    * Stores the log_base_2 of the desired data_width.
    * Used only as a helper attribute to randomize data_width.
    * This parameter is first randomized and the data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_data_width;

  /**
    * Stores the log_base_2 of the desired snoop_data_width.
    * Used only as a helper attribute to randomize snoop_data_width.
    * This parameter is first randomized and the snoop_data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_snoop_data_width;

  /**
    * Stores the log_base_2 of the desired cache_line_size.
    * Used only as a helper attribute to randomize cache_line_size.
    * This parameter is first randomized and the cache_line_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_cache_line_size;

  /**
    * Stores the log_base_2 of the desired atomicity_size.
    * Used only as a helper attribute to randomize atomicity_size.
    * This parameter is first randomized and the atomicity_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_atomicity_size;

  /** @endcond */

  /** 
    * @groupname axi3_signal_width
    * Address width of this port in bits.
    * When svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE,
    * this parameter also sets the width of signal caddr.
    *
    * NOTE: currently same address width is considered for both coherent read or write address
    *       channels and snoop address channels. So, there is no separate snoop address width
    *       parameter supported at the moment.
    * Configuration type: Static
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE 
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH;
`else    
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH - `SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH;
`endif   

  /** 
    * @groupname axi4_signal_width
    * Address user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int addr_user_width = `SVT_AXI_MAX_ADDR_USER_WIDTH;

  /** 
    * @groupname axi3_signal_width
    * Data width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_width = `SVT_AXI_MAX_DATA_WIDTH;

  /** 
    * @groupname axi4_signal_width
    * Data user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_user_width = `SVT_AXI_MAX_DATA_USER_WIDTH;
 
  /** 
    * @groupname axi4_signal_width
    * Response user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int resp_user_width = `SVT_AXI_MAX_BRESP_USER_WIDTH;

  /** 
    * @groupname ace_config
    * Cache line size in bytes for this master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int cache_line_size = `SVT_AXI_MAX_CACHE_LINE_SIZE;

  /** 
    * @groupname ace_config
    * Aligned size in bytes for the snoop corresponding to starting address.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates the size to which the snoop corresponding to the starting address
    * of a multi-cacheline access is aligned. For example, if the cacheline size
    * is 64 bytes and the coherent address of a READONCE transaction is 0x70,
    * the corresponding snoop address may be 0x40 or 0x70. If the snoop address
    * sent is 0x40, this value must be set to the same as the cacheline size which is
    * 64 bytes. If the snoop address sent is 0x70, this value can be set to 16 bytes.
    * This will help in more accurate correlation of coherent and snoop transactions.
    * The default is 0. If unchanged, the system monitor will use the cacheline size
    * for this value, assuming that all snoops are aligned to cacheline size. 
    * Configuration type: Static
    */
  rand int start_addr_snoop_aligned_size = 0;

  /** 
    * @groupname ace_config
    * Number of cache lines in the master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int num_cache_lines = `SVT_AXI_MAX_NUM_CACHE_LINES;

  /** 
    * @groupname ace_config
    * Enables AWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default AWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit awakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Enabling this feature will allow transactions to wait to send address phase
    * until the previous transaction's datahandshake is done. This will result
    * in unexpected delays. Hence this parameters is disabled by default.
    * 
    * This parameter is applicable when 
    * svt_axi_port_configuration::axi_interface_type is set to AXI3 or AXI4.
    *
    * Configuration type: Static
    */
  rand bit prev_xact_data_handshake_ref_event_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_max_delay_during_idle = 5;


  /** 
    * @groupname ace_config
    * Enables ACWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default ACWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit acwakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_max_delay_during_idle = 5;
  
  /** 
    * @groupname ace_signal_width
    * Snoop Data width of the cddata port in bits.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Configuration type: Static
    */
  rand int snoop_data_width = `SVT_AXI_ACE_SNOOP_DATA_WIDTH;

  /**
    * @groupname axi3_4_config
    * Acronym for "What You See is What You Get". Applicable to the
    * svt_axi_transaction::data and svt_axi_transaction::wstrb fields of a
    * transaction. If this bit is set to 1, whatever is configured in the
    * svt_axi_transaction::data and  svt_axi_transaction::wstrb fields is
    * transmitted "as is" by the master. Also, in the transaction object
    * generated by monitor, the monitor populates the svt_axi_transaction::data
    * and  svt_axi_transaction::wstrb fields "as is", as seen on the bus. If
    * this bit is set to 0 (default), the data must be stored right-justified by
    * the user. The model will drive the data on the correct lanes.
    *
    * Refer to the documentation of svt_axi_transaction::data and 
    * svt_axi_transaction::wstrb for more details
    */
  rand bit wysiwyg_enable = 0;

  /**
    * @groupname axi3_4_config
    * Applicable when #wysiwyg_enable is set.
    * Indicates if the VIP should consider validity of wstrb in transactions
    * when #wysiwyg_enable is set. When wysiwyg_enable is set, the driver
    * checks that #wstrb is set only for valid byte lanes of each beat.  In
    * certain applications, wstrb may have to be asserted for other byte lanes
    * as well. In such applications, this bit should be set. This results in
    * the following: 
    * <br>
    * Constraints in transaction are relaxed for wstrb. wstrb
    * values will be random and may be asserted for invalid byte lanes. 
    * <br>
    * driver does not check for validity of wstrb in transaction based on valid
    * byte lanes.
    * <br>
    * Note that this will result in a non-AXI compliant behaviour, in that
    * wstrb may be asserted for invalid byte lanes based on what the user
    * programs. If this bit is set for the slave, and if the user wants memory
    * to be updated based on the transactions, the memory sequence shipped with
    * the VIP should not be used. For VMM based testbenches, the generator_type
    * should not be set to MEMORY_RESPONSE_GEN. This is because the APIs that
    * access memory are based on valid assertion of byte strobes.  The user
    * must use user-defined APIs and sequences to access memory if this bit is
    * set in the slave.
    */ 
  bit ignore_wstrb_check_for_wysiwyg_format = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal on byte count calculation in the VIP 
    * By default this configuration parameter is set to 0 to calculate the byte count using burst_size and burst_length,
    * if this parameter is set 1 then wstrb is used to calculate the byte count
    * <b>type:</b> Static
    */
  rand bit get_byte_count_from_wstrb_enable      = 0;

   /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWREGION signal in the VIP 
    * <b>type:</b> Static
    */

  rand bit awregion_enable   = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARREGION signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arregion_enable   = 0;
 
  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awqos_enable      = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wlast_enable      = 1;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wstrb_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bresp_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arqos_enable      = 0;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rresp_enable      = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rlast_enable      = 1;

  /** 
    * @groupname axi3_4_config
    * Enables AWUSER sideband signal in the VIP. AWUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit awuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables WUSER sideband signal in the VIP. WUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit wuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables BUSER sideband signal in the VIP. BUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit buser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables ARUSER sideband signal in the VIP. ARUSER signal can be used when
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit aruser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables RUSER sideband signal in the VIP. RUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit ruser_enable      = 0;

  `ifdef SVT_AXI_QVN_ENABLE
  /** 
    * @groupname axi_qvn_config
    * Enables QVN support in the VIP. QVN signals can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * All QVN configuration parameters comes into effect only when qvn_enable bit is set.
    * Any parameter which is declared as a bit-vector to support all Virtual Network in the
    * system, is sized by `define macro "SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK".
    *
    * If a system should support a maximum number of 5 Virtual Networks then user should
    * define SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK as 5
    * <b>type:</b> Static
    */
  rand bit qvn_enable      = 0;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Read Address channel
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_ar_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Write Address channel.
    * Write Data channel must support Virtual Networks same as Write Address channel so there is
    * no need of having seperate configuration for Write Data channel.
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_aw_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Read-Address Channel.
    * It provides an array of bits each representing a Virtual Network in the system. Index of 
    * each bit denotes ID of the Virtual Network, represented by that bit.
    * If any bit of this array is set to '1' then that means Virtual Network with ID equal to
    * index of that bit, is supported by this port. If a bit in this array is set to '0' then
    * that means Virtual Network with ID equal to its index is not supported by this port.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 1 and 3 to be used for its
    *           Read-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_ar_chnl[index]) qvn_supported_virtual_network_queue_ar_chnl[index] = 0; 
    *   set '1' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_ar_chnl[1] = 1;
    *   set '1' for Virtual Network 3 =>  qvn_supported_virtual_network_queue_ar_chnl[3] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_ar_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Write Address Channel.
    * This array of bits also indicate which Virtual Networks are supported by this port similar
    * to the array qvn_supported_virtual_network_queue_ar_chnl described above.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 0 and 2 to be used for its
    *           Write-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_aw_chnl[index]) qvn_supported_virtual_network_queue_aw_chnl[index] = 0; 
    *   set '0' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_aw_chnl[1] = 1;
    *   set '1' for Virtual Network 2 =>  qvn_supported_virtual_network_queue_aw_chnl[2] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_aw_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on read address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */

   /* If a Master is not able to use a token, then after this timelimit that token will be reclaimed
    * by the slave which, granted it and Master will remove this token from its reserved token pool.
    *
    * - So, it is important to set suitable value for this parameter. If it is set too low, then
    * most tokens may expire before it could be used and hance leading to increased token request.
    *
    * - If it is set below minimum no. of cycles a master needs to use a token then all tokens will
    * expire and none could be used to issue a transaction to AXI channels.
    *
    * - On the other hand if it uses too high value, then due to under usage of token or over-request
    * of tokens by a Master, there is a possibility of accumulating large number of tokens in the
    * token-pool of that master and hence causing possible blockage to other masters.
    *
    * - If it is set to Zero then that indicates there is no timelimit for token usage i.e. once a 
    * token is acquired it will remain in the token-pool of that master until used for sending a
    * transaction.
    * .
    */
  rand int qvn_read_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write data channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_data_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Read Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AR_PRE_ALLOCATED_TOKEN
    * Example: if AR channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_ar_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_ar_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Write Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AW_PRE_ALLOCATED_TOKEN
    * Example: if AW channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_aw_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_aw_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Indicates if same AXI ID can be used between two different Virtual Network or not.
    * - If set to "0" then at any given point of time no two different Virtual Networks will
    * use same ID for transactions sent to AXI channels associated with those VNs.
    * - if set to "1" then same AXI ID can be used by two different VN without any restriction.
    * .
    *
    * NOTE: if same ID is used for AXI transactions issued to two different VN may get
    * blocked by interconnect in order to observe AXI ID ordering rule. Because of this, a
    * transaction received first will block another transaction with same ID received later,
    * even if transaction that was received first, can't make any progress.
    */
  rand int qvn_allow_id_used_in_other_vn = 0;

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on read address channel. It helps in defining how system resources will be used
    * otherwise, a master can issue large number of token requests and once granted those tokens 
    * may remain unused reserving system resources and in turn blocking other masters, if it shares 
    * same Virtual Network or if slave uses shared token for different masters.
    * 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_read_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write address channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write data channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_data_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for read address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for read address channel.
    */
  rand int unsigned qvn_ar_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write address channel.
    */
  rand int unsigned qvn_aw_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write data channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write data channel.
    */
  rand int unsigned qvn_w_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];


  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AR channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AR channel
    */
  rand int qvn_slave_ar_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AW channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AW channel
    */
  rand int qvn_slave_aw_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for W channel for a particular Virtual Network
    * This means Slave has this many token resource to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Master doesn't have any pre-allocated token for Write Data channel so, Slave will 
    *       begin with same number of Tokens as specified by this parameter.
    */
  rand int qvn_slave_w_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for read address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_rd_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write data channal for a VN, 
    * in accordance with slaves acceptance capability.
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_data_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

   /**
    * @groupname axi_qvn_config
    * Mode to control the assertion of V*READYVNx signal. This allows QVN enabled Slaves to assert
    * token request grant ready signal for any Virtual Network of each channel AR, AW, W
    *
    * 0 - Assert V*READY in responce to assertion of V*VALID for token request 
    * 1 - Assert V*READY before assertion of V*VALID for token request, subjected to token availability
    */  
   rand bit qvn_slave_aw_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_assertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
  
   /*
    * @groupname axi_qvn_config
    * Mode to control the de-assertion of V*READYVNx signal. This flage is only 
    * applicable if v*ready_assertion_mode is set to ONE.
    * 0 - Keep V*READY till assertion of V*VALID.  
    * 1 - Deassert V*READY after some time if V*VALID is not asserted. 
    */  
   rand bit qvn_slave_aw_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_deassertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};


  `endif

  /** 
    * @groupname axi3_4_config
    * Enables optimistic flow control for Write Data channel in the VIP.  
    * The flow control of the write data channel is determined by the settings 
    * in num_outstanding_xact and num_outstanding_write_xact. Based on these 
    * settings wready is deasserted when the number of outstanding transactions
    * reach the threshold set by these parameters. This parameter controls the 
    * deassertion of wready when the threshold is reached. Since AXI allows data 
    * before address, a new transaction can start with data. When this parameter 
    * is disabled, both awready and wready are deasserted when threshold of maximum
    * outstanding transactions are reached. Note however that this will prevent data
    * of any already outstanding transactions from being continuously accepted
    * (that is with wready continuously high) and therefore can reduce throughput
    * If this parameter is set, only awready is deasserted when the threshold is reached.
    * This allows data of outstanding write transactions to be continously accepted
    * with wready maintained high continuosly. wready is deasserted only on observing
    * a new transaction which will cross the threshold. Thus, setting this configuration
    * assumes that write data before address doesn't come once the threshold for maximum
    * outstanding transactions is reached and thus keeps wready asserted. 
    * Whereas disabling this configuration assumes that write data before address might 
    * come and thus deasserts wready when number of outstanding transactions
    * reach the threshold.
    * <b>type:</b> Dynamic
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand bit wdata_optimistic_flow_control_enable = 0;
`else
  rand bit wdata_optimistic_flow_control_enable = 1;
`endif

   /** 
    * @groupname axi3_4_config
    * Passive slave memory needs to be aware of the backdoor writes to memory.
    * Setting this configuration allows passive slave memory to be updated according to
    * RDATA seen in the transaction coming from the slave. Note that the passive slave 
    * memory is updated when all read data beats have been transmitted and accepted.
    * For an EXCLUSIVE transaction memory is updated only if all beats have an EXOKAY response.
    * For a normal transaction, memory is updated only if all beats have an OKAY response.
    * <b>type:</b> Static
    */
  rand bit memory_update_for_read_xact_enable = 0;

  /**
    * @groupname axi3_signal_width
    * Indicates if separate widths are required for ID  of write channel 
    * (AWID,WID and BID) and for ID of read channel(ARID and RID).
    * If set to 1, read_chan_id_width and write_chan_id_width are used
    * for setting the widths of the ID signals of corresponding channels.
    * If set to 0, id_width is used for setting the widths of all
    * ID signals.
    * This value must be consistent across all the ports in the system.
    *
    * Configuration type: Static
    */
  rand bit use_separate_rd_wr_chan_id_width = 0;

  /**
    * @groupname axi3_signal_width
    * If port is of kind MASTER:
    * This parameter defines the ID width of the master.
    * <br>
    * If port is of kind SLAVE:
    * This parameter defines the ID width of the slave. If an
    * interconnect is present, the ID width of the slave should
    * consider the maximum ID width of the masters in the system
    * and also consider additional bits required to represent
    * each master in the system.
    * <br>
    * Valid only when use_separate_rd_wr_chan_id_width is set to 0.
    *
    * Configuration type: Static
    */
  rand int id_width  = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of ARID and RID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int read_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of AWID, WID and BID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int write_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with barrier transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit barrier_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_min  = 0;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with DVM transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit dvm_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_min  = ((1<<(`SVT_AXI_MAX_ID_WIDTH/2))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the max ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
   * Indicates how the information regarding the source master is 
   * transmitted to the slave
   * If set to STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is static and is defined by #source_master_id_xmit_to_slaves
   * If set to DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is based on the value defined in svt_axi_transaction::dynamic_source_master_id_xmit_to_slaves
   * The value in dynamic_source_master_id_xmit_to_slaves must be populated by the user
   * in a system monitor callback issued at the start of the transaction.
   * If set to CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the user must define 
   * svt_axi_system_configuration::is_master_id_and_slave_id_correlated to indicate
   * whether ID requirements for master and slave transactions are met 
   */
  source_master_id_xmit_to_slaves_type_enum source_master_id_xmit_to_slaves_type = STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES;
  
 /**
   * @groupname ace5_config 
   * Indicates whether data check parity feature is enable or not.
   * If set to ODD_PARITY_BYTE_DATA, then only on data check signals odd parity algorthim is used,
   * every 8bit of data is calculated and generated singles bit of datachk parity bit.
   * If set to ODD_PARITY_BYTE_ALL, then on both data check signals and control check signals odd parity algorthim is used.  
   * By default this enum is set to FALSE, which means data check fetaure is disabled.
   */ 
  check_type_enum check_type = FALSE;



  /**
    * @groupname axi_generic_config 
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If port is of kind MASTER:
    * This parameter defines the value that the interconnect assigns when
    * routing transactions to slave for all transactions originating from this
    * master. This value is specified in some bits of AxID of the transaction
    * that is routed to slave. This value must be based on the max value that
    * can be supported based on
    * svt_axi_system_configuration::source_master_info_id_width. For example, if the
    * interconnect uses 3 bits of AxID of the outgoing slave transaction to
    * specify the source master of the transaction,
    * svt_axi_system_configuration::source_master_info_id_width must be set to 3 and
    * this value must be less than 7. For more details, please refer
    * svt_axi_system_configuration::id_based_xact_correlation_enable
    */
  bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id_xmit_to_slaves;

  /**
    * @groupname axi_generic_config
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * and axi_port_kind is MASTER
    * Indicates that the ID from this master is passed through without any
    * change when the interconnect routes it to the slaves. If this is set,
    * all transactions from this master are not appended with source master
    * information when routing to slaves
   */ 
  rand bit is_source_master_id_and_dest_slave_id_same = 0;

  /**
    * @groupname axi_generic_config 
    * Applicable only when svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If this parameter is set to zero, system monitor will not do id based correlation
    * for any transactions initiated/received at this specific port, this provides the option
    * for the user to avoid or select id based correlation for specific ports 
    * default value is 1.
    */
  bit id_based_xact_correlation_enable =1'b1;

  /** 
    * @groupname axi_generic_config
    * The byte boundary at which a master transaction is split to be
    * transmitted to two different slaves. This must be defined in cases where
    * pre_add_to_input_xact_queue callback in svt_axi_system_monitor_callback
    * is used to indicate that a master transaction is split and transmitted to
    * two different slaves. This parameter defines the boundary at which a
    * transaction is split
    *
    * Configuration type: Static
    */
  rand int byte_boundary_for_master_xact_split = `SVT_AXI_MAX_BYTE_BOUNDARY_FOR_MASTER_XACT_SPLIT;

  /**
   * @groupname ace_config
   * Enables support for WriteEvict transaction
   * Configuration type: Static
   */
  rand bit writeevict_enable = 0;

  /**
   * @groupname ace_config
   * Enables AWUNIQUE signal 
   * Configuration type: Static
   */
  rand bit awunique_enable = 0;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of outstanding transactions a master/slave
    * can support.
    * num_outstanding_xact = -1 is not supported for AXI4_STREAM
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY/AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * If #num_outstanding_xact = -1 then #num_outstanding_xact will not 
    * be considered , instead #num_read_outstanding_xact and 
    * #num_write_outstanding_xact have an effect.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_outstanding_xact = 4;

  /**
    * @groupname axi3_4_config
    * Specifies the number of READ outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_read_outstanding_xact = 4;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of WRITE outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_write_outstanding_xact = 4;

  /** 
    * @groupname ace_config
    * Specifies the number of outstanding snoop transactions a master
    * can support. Applicable when axi_interface_type == AXI_ACE.
    * If the number of outstanding snoop transactions is equal to 
    * this number, the master will not assert ACREADY 
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_SNOOP_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int num_outstanding_snoop_xact = 4;
`else
  rand int num_outstanding_snoop_xact = 16;
`endif  

  /** 
    * @groupname axi_generic_config
    * 
    * Enables a separate port/export in the slave driver
    * (delayed_response_request_export) and sequencer
    * (delayed_response_request_port) through which the user can input response
    * data in a delayed manner.  When disabled all data and response
    * information related to a transaction must be given back to the driver
    * from the sequencer in the same timestamp as it receives a transaction
    * from the monitor.  When enabled, the user has flexibility to provide
    * response and data information at a later point in time through the
    * response port in the slave driver, although parameters related to the
    * delays to be applied for driving ARREADY, AWREADY and WREADY signals need
    * to be provided in the same timestamp. 
    * Refer to the user guide for a detailed description of the usage of this
    * parameter.
    */ 
  bit enable_delayed_response_port = 0;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of exclusive access transactions.
    * <br>
    * SLAVE:
    * Indicates whether the slave supports exclusive access or not.
    * <b>type:</b> Static
    *
    */
  rand bit exclusive_access_enable = 0;
  
  /** 
    * @groupname ace_config
    * MASTER:
    * This is applicable only when svt_axi_port_configuration::exclusive_access_enable is set to 1.
    * This bit controls enabling  Exclusive Monitor for AXI and ACE Masters.
    * If it is set to '1' then exclusive monitor is enabled in ace masters cache is updated on successful exclusive transactions based on coherent response and exclusive monitor state.
    * If this is set to '0' then exclusive monitor is disabled in ace master and for exclusive transaction cache
    * is updated only based on coherent response i.e. if it is received as EXOKAY.
    * <b>type:</b> Dynamic
    */
  rand bit exclusive_monitor_enable = 1;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of locked access transactions.
    * <b>type:</b> Static
    *
    */
  rand bit locked_access_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of barrier transactions.
    * <b>type:</b> Static
    */
  rand bit barrier_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of DVM transactions.
    * <b>type:</b> Static
    */
  rand bit dvm_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only for active master 
    * Enables automated generation of DVMCOMPLETE transactions
    * in response to DVM Sync Snoop transactions. 
    * When this bit is unset, it is the user's responsibility to
    * send DVMCOMPLETE transactions from the sequence in response
    * to DVM Sync snoop transactions.
    * When this bit is set, the VIP master driver will auto generate 
    * DVMCOMPLETE transaction in response to DVM Sync snoop transactions.
    * When this bit is set, any DVMCOMPLETE transaction received from the sequencer will be ignored.
    */
  rand bit auto_gen_dvm_complete_enable = 0;

  /**
    * The minimum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int min_auto_gen_dvm_complete_delay = 0;

  /**
    * The maximum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver.
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int max_auto_gen_dvm_complete_delay = `SVT_AXI_MAX_DVM_COMPLETE_DELAY;

  /**
    * If this parameter is set, when a DVM snoop sync is received, the driver
    * takes a snapshot of active transactions whose address or data have been
    * sent on the interface.  The DVMCOMPLETE on the read address channel is
    * then launched when these outstanding transactions are complete. The
    * parameter #dvm_complete_delay is not applicable if this parameter is set. 
    */
  bit launch_auto_gen_dvm_complete_on_outstanding_xact_completion = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables speculative read.
    * A speculative read is defined as a read of a cache line that a master may
    * already be holding in its cache. Consider a case when user generates a
    * coherent transaction for read of a cache line that a master already holds
    * in its cache.
    *
    * When speculative read is enabled, the master will transmit this coherent
    * transaction. Also, the master will support cache state transitions as
    * defined in second set of tables in sections 5.5.1 to 5.5.11 in ACE
    * proposal 0.27.
    *
    * When speculative read is disabled, the master will not transmit this
    * coherent transaction. In this case, the master will only support cache
    * state transitions as defined in first set of tables in sections 5.5.1 to
    * 5.5.11 in ACE proposal 0.27.
    *
    * Whether a transaction is a speculative read is indicated by read-only
    * transaction class member svt_axi_transaction::is_speculative_read.
    *
    * <b>type:</b> Dynamic
    */
  rand bit speculative_read_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables restrictions in the master for support of an external
    * snoop filter.
    * <b>type:</b> Dynamic
    */
  rand bit snoop_filter_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE_LITE.
    *
    * SLAVE:
    * Checks that cache maintenance transactions received by an interconnect
    * from a master are forwarded to corresponding slaves. This check will
    * be performed only if the system monitor is enabled and correlation of
    * master and slave transactions are enabled by setting 
    * id_based_correlation_enable in svt_axi_system_configuration and the associated
    * configuration properties. 
    * <b>type:</b> Dynamic
    */
  rand bit forward_cmos_to_slaves_check_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    * MASTER:
    * Determines the permissible cache line state transitions in the master.
    * For each transaction type, the section 5 of the specification provides 
    * cache line state transitions for "expected (or recommended) end state", 
    * "legal end state with snoop filter" and "legal end state without snoop filter".  
    * This parameter determines which of the above state changes are to be
    * used.
    *
    * Below are the supported values:
    * - RECOMMENDED_CACHE_LINE_STATE_CHANGE: The cache line state
    * changes as given in the "expected end state" of each table is used.
    * - LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state with snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 1. The actual cache line state change can be done using
    * member svt_axi_transaction::force_to_shared_state.
    * - LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state without snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 0. The actual cache line state change can be done using
    * members svt_axi_transaction::force_to_invalid_state and
    * svt_axi_transaction::force_to_shared_state.
    * .
    *
    * <b>type:</b> Dynamic
    */
  rand axi_cache_line_state_change_type_enum cache_line_state_change_type = RECOMMENDED_CACHE_LINE_STATE_CHANGE;

  /**
   * @groupname ace_config
   * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component.
   *
   * Specifies how master will process incoming snoop request when memory update transaction is in progress.
   * if it is set to SUSPEND_SNOOP_DURING_MEM_UPDATE then master will suspend incoming snoop request and will respond
   * after current memory update transaction is complete. This is the default response mode.
   * If it is set to RESPOND_SNOOP_DURING_MEM_UPDATE then master will not suspend incoming snoop request. Instead it will
   * respond to the incoming snoop request as allowed by ACE specification.
   * If it is set to EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE then master will randomly decide to choose between
   * either of the above two behaviour i.e. either suspend incoming snoop or respond to it.
   * 
   * Configuration type: Dynamic
   */
  rand snoop_response_mode_during_mem_update_type_enum snoop_response_mode_during_mem_update = SUSPEND_SNOOP_DURING_MEM_UPDATE;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component
    *
    * Indicates how dirty data in cache should be transferred on receiving a snoop.
    * As per section C5.2.2 of the AXI specification, a cached master can ensure that data in a dirty cacheline
    * is available to a snoop other than MAKEINVALID in one of two ways:
    * 1. returning data when the master completes the snoop
    * 2. carrying out a memory update, using a WRITEBACK or WRITECLEAN before responding to the snoop
    * This configuration indicates which of the above two methods will be used for returning data
    * Note that if there is an outstanding WRITEUNIQUE or WRITELINEUNIQUE transaction in the
    * queue of the master, then data will be returned with the snoop transaction. This is to comply with
    * restrictions on WRITEUNIQUE and WRITELINEUNIQUE while a snoop is in progress as per section
    * C4.8.7 of the spec
    */
  rand snoop_response_data_transfer_mode_enum snoop_response_data_transfer_mode = SNOOP_RESP_DATA_TRANSFER_USING_CDDATA;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE and it is Master component
    *
    * Describes various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE. It indicates what
    * address range should or shouldn't be used while randomizing axi master transaction based on the different enum values listed below.
    *
    * NONSHAREABLE_XACT_FULL_ADDRESS_SPACE :: allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE :: allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE :: allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE :: allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * default value :: NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE
    */
  rand nonshareable_xact_address_range_in_systemshareable_mode_enum nonshareable_xact_address_range_in_systemshareable_mode = NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE;

  /**
    * @groupname axi3_4_config
    * MASTER:
    * The maximum number of active exclusive transactions that will be initiated by the master.
    * SLAVE:
    * The maximum number of active exclusive access monitors supported by the slave. Attempts to
    * exceed this max number results in a failed exclusive access read response of OKAY instead of EXOKAY.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS
    * NOTE: if it is set to '0' value then there are no restrictions on maximum number of active exclusive
    * transactions. VIP will not mark any exclusive sequence as failed because of this parameter.
    * <b>type:</b> Static
    */ 
  rand int max_num_exclusive_access   = `SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS;
      
  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Number of ADDRESS bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    *
    * It can also be configured with ( -1 ) to indicate that address ranges for 
    * each exclusive monitor is defined through user specified start and end address ranges.
    * For this, user should configure start_address_ranges_for_exclusive_monitor[] and
    * end_address_ranges_for_exclusive_monitor[] arrays in system configuration.
    * A svt_axi_system_configuration::set_exclusive_monitor_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,
    *     bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr) utility method can be used for this purpose.
    *
    * NOTE: configuring with value 0 means, no address is being monitored by the 
    * corresponding exclusive monitor and hence exclusive access to different address
    * may also affect current thread.
    *
    * <b>specail value:</b> -1 indicates that num_addr_bits_used_in_exclusive_monitor and
    * num_initial_addr_bits_ignored_by_exclusive_monitor are not used. Instead address
    * ranges for exclusive monitors are defined by address_ranges_for_exclusive_monitor[] array.
    *
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ADDR_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_addr_bits_used_in_exclusive_monitor   = `SVT_AXI_MAX_ADDR_WIDTH;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * ACE Exclusive monitor will ignore number of initial address bits as
    * indicated by this configuration member.
    * Example: A coherent interconnect can divide its whole address space into
    *          multiple ranges such that each PoS Exclusive monitor checks only
    * its corresponding address range. So, if it allocates 1/2 GB address space to each
    * of the 4 PoS exclusive monitors then num_initial_addr_bits_ignored_by_exclusive_monitor
    * needs to be configured as 29 (1.5GB - 2GB ~ 31 bits).
    */
  rand int num_initial_addr_bits_ignored_by_exclusive_monitor   = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE
    * INTERCONNECT:
    * Number of ID bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    * NOTE: configuring with value 0 means, no id is being monitored by the 
    * corresponding exclusive monitor and hence only single exclusive access thread
    * is supported for current port.
    *  <b> This feature is not supported yet </b>
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ID_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_id_bits_used_in_exclusive_monitor     = `SVT_AXI_MAX_ID_WIDTH;

   /*
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Indicates whether Interconnect uses seperate PoS Exclusive Monitor for 
    * secured or non-secured exclusive access.
    * NOTE: configuring with value 0 means, interconnect doesn't monitor seperately
    * for secured or unsecured exclusive access.
    * <b> This feature is supported by enabling secure address space by configuring tagged_address_space_attributes_enable = 1 </b>
    * <b> User shouldn't use this configuration parameter, it is going to be deprecated </b> 0
    * <b>min val:</b> 0
    * <b>max val:</b> 1
    * <b>type:</b> Static
    */ 
  rand bit use_secured_exclusive_monitor             = 1;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will not assert error if Master sends Exclusive Store without sending Exlusive Load.
    * However, if Exclusive Store is sent from the Invalid cacheline state then VIP will still assert error since,
    * that is not a valid state to start Exclusive Store.
    * <b>type:</b> Static
    */ 
  rand bit allow_exclusive_store_without_exclusive_load = 0;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will respond to very first Exclusive Store with EXOKAY response. This means that if
    * no master has performed any exclusive transaction after reset is de-asserted then the master that issues
    * exclusive store will be responded with EXOKAY or VIP will expect EXOKAY response from the coherent interconnect.
    * Note: reference point of first exclusive store is reset.
    * <b>type:</b> Static
    */ 
  rand bit allow_first_exclusive_store_to_succeed = 0;

  /**
    * @groupname ace_config
    * If set to '1' then Exclusive Monitor will get reset once Exclusive Store is successful.
    * If set to '0' then Exclusive Monitor will remain set even if Exclusive Store is successful.
    * Please Note that, VIP will still reset Exclusive Monitor for failed Exclusive Store attempt
    * regardless of the value set for this parameter.
    * <b>type:</b> Static
    */ 
  rand bit reset_exclusive_monitor_on_successful_exclusive_store = 1;

  /**
    * @groupname ace_config
    * This control register indicates different modes of error conditions uded in exclusive monitor.
    * [0] => If set to '1' implies that Snoop Error will cause an exclusive sequence to fail only if
    *        either data_transfer bit or pass_dirty bit is set to '1'. Otherwise, if snoop response
    *        indicates error bit as asserted then regardless of data_transfer bit or pass_dirty bit
    *        values exclusive sequence will fail. 
    * [31:1] => Reserved bits.
    * Default Value :: 0x00000000
    */
  rand bit[31:0] exclusive_monitor_error_control_reg = 0;

  /** 
    * @groupname ace_config
    * If shareable exclusive access needs to be supported from ace-lite port then this parameter
    * should be set to '1'. If it is set to '1' then VIP will allow READONCE or WRITEUNIQUE
    * transactions to be of exclusive type.
    * Default Value: '0' i.e. shareable exclusive access from ace-lite port is not allowed. Only
    *                non-shareable exclusive transactions as READNOSNOOP or WRITENOSNOOP are allowed.
    */
  rand bit shareable_exclusive_access_from_acelite_ports_enable = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of write transactions that can be interleaved
    * This parameter should not be greater than #num_outstanding_xact.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted write data beyond this value.
    * SLAVE: 
    * Checks that received write data is not interleaved beyond this value. 
    * An error is issued if write data is interleaved 
    * beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int write_data_interleave_depth       = `SVT_AXI_MAX_WR_INTERLEAVE_DEPTH;

  /** 
    * @groupname axi3_4_config
    * This parameter specifies the atomicity size required to check the address
    * alignment for a given transcation as per the atomicity of component.<br>
    * This parameter will not have effect if set to -1. The values specified
    * to this parameter should be power of 2, in terms of Bytes <br>
    * Default value: -1.<br>
    * Allowed values: should be power of 2, in terms of Bytes. <br>
    * For example: 8, 16, 32, 64 etc <br>
    * <b>type:</b> Static
    *
    */
  rand int atomicity_size = -1;


  /** @cond PRIVATE */
  /**
    * When set to 1, enables id reflection in AXI4_LITE mode.
    * This enables the awid, bid and rid signals. This allows
    * an AXI4-Lite slave to be used on a full AXI interface,
    * without a bridge function, in a system that guarantees that
    * the slave can only be accessed by transactions that fall
    * within the AXI4-Lite subset.
    * <b>type:</b> Static
    *
    * This parameter is not yet supported.
    */
  rand bit id_reflection_enable = 0;
  /** @endcond */

  /**
    * @groupname axi3_4_config
    * Applicable only to MASTER when axi_interface_type is 
    * AXI3/AXI4/AXI4_LITE.
    * When set to 1, accesses to the read address channel and 
    * write address channel are serialized. Thus, awvalid and
    * arvalid will never be asserted at the same time. The
    * address information driven on the write address channel
    * will have to be accepted before any address information
    * on the read address channel is driven and viceversa. 
    * When set to 0, activity on the read address channel and
    * write address channel occur in parallel.
    */
  rand bit serial_read_write_access = 0;

`ifndef SVT_EXCLUDE_VCAP
  /**
    * @groupname axi_traffic_profile 
    * Enables use of traffic profiles. This enables the use of transaction
    * generation at a higher level of abstraction.  This feature
    * is only available as part of the NOC product. Please refer to the NOC
    * user guide for details
    */
  bit use_traffic_profile = 0;

  /** 
    * @groupname axi_generic_config
    * Enables FIFO based rate control. 
    * A FIFO is modelled in the driver for read and write
    * transactions separately. A WRITE transaction can be sent
    * out if there is sufficient data in the FIFO to send out that
    * transaction. A READ transaction can be sent out if there is
    * space in the FIFO to receive the data of the READ transaction.
    * The current level of a WRITE FIFO is incremented every clock
    * based on write_fifo_fill_rate.With every data beat, the currentl level
    * is decremented based on burst_size of the transaction. The current level of a READ FIFO
    * is decremented every clock based on read_fifo_drain_rate. With every data
    * beat, the current level is incremented based on burst_size of the transaction.
    * A WRITE transaction will be sent out if the current level is greater than
    * the total number of bytes of all outstanding write transactions + the total
    * number of bytes of the current transaction. A READ transaction will be sent out
    * if the current level is less than the difference of the read_fifo_full_level and
    * the total number of bytes of all outstanding read transactions + the total number
    * of bytes of the current transaction.
    */
  rand bit use_fifo_based_rate_control = 0;

  /**
    * @groupname axi_generic_config
    * Clock period in ns. This is used to calculate the drain/fill rate in
    * bytes/cycle
    */
  real clock_period = 1;

  /** 
    * @groupname axi_generic_config
    * The drain rate in MBPS of the FIFO into which data from READ
    * transactions is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction
    */
  rand int read_fifo_drain_rate = `SVT_AXI_MAX_READ_FIFO_DRAIN_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the READ FIFO into which data from READ transactions
    * is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction.
    */
  rand int read_fifo_full_level = `SVT_AXI_MAX_READ_FIFO_FULL_LEVEL;

  /** 
    * @groupname axi_generic_config
    * The fill rate in MBPS of the FIFO from which data for WRITE 
    * transactions is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to send a WRITE transaction
    */
  rand int write_fifo_fill_rate = `SVT_AXI_MAX_WRITE_FIFO_FILL_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the WRITE FIFO from which data for WRITE transactions
    * is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to transmit data of a WRITE transaction
    */
  rand int write_fifo_full_level = `SVT_AXI_MAX_WRITE_FIFO_FULL_LEVEL;

  /**
    * @groupname axi_generic_config
    * Determines if the READ FIFO is empty on start up
    */
  rand bit is_read_fifo_empty_on_start = 1;

  /**
    * @groupname axi_generic_config
    * Determines if the WRITE FIFO is empty on start up
    */
  rand bit is_write_fifo_empty_on_start = 1;
`endif //SVT_EXCLUDE_VCAP

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, AXI transaction phase level information is
    * printed in note verbosity.  Messages related to start & end of address,
    * data and response phases are printed.  If unset, AXI transaction phase
    * level information is printed only in debug verbosity.
    */ 
  bit display_xact_phase_messages = 0;

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding transactions
    * per AxID is limited to 1 for Non-Device and Non-DVM transactions.
    * This can be further controlled by configuration
    * svt_axi_port_configuration::single_outstanding_per_id_kind. 
    */ 
  bit single_outstanding_per_id_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding AXI4_STREAM transactions
    * per TDEST is limited to 1.
    */ 
  bit single_outstanding_per_tdest_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set to 1, all delay related parameters will be set
    * to 0. Note however, that actual delay on interface will vary based on
    * outstanding transactions.
    */ 
  rand bit zero_delay_enable = 0; 
  
  /**
    * This enumerated type controls the AxID when
    * svt_axi_port_configuration::single_outstanding_per_id_enable is set to 1.
    *
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * 'MODIFY_SAME_ID': If AxID of a new Non Device or Non DVM transaction matches
    * AxID of an active transaction, the VIP modifies the AxID such that the AxID 
    * is not overlapping with AxID of any active Non Device or Non DVM transactions.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated
    * by the user sequence. At this time, another Non Device or Non DVM with AxID = 6
    * is already in progress. In this case, VIP will check the active queue, and modify
    * the AxID of the new transaction to an un-used AxID. For example, VIP will modify 
    * the AxID of new transaction to 4, if this is not used by any active transactions.
    * 
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * ‘WAIT_FOR_COMPLETION_OF_SAME_ID': If AxID of a new Non Device or Non DVM transaction
    * matches AxID of an active Non Device or Non DVM transaction, the VIP waits till the
    * corresponding active Non Device or Non DVM transaction is complete. Only when the
    * active Non Device or Non DVM transaction is complete, VIP adds the new Non Device
    * or Non DVM transaction to the active queue. This ensures that only 1 active Non Device
    * or Non DVM transaction exists for a given AxID.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated by
    * the user sequence. At this time, another Non Device or Non DVM with AxID = 6 is already
    * in progress. In this case, VIP will wait for the active transaction to complete. After
    * active transaction is complete, VIP will add the new transaction with AxID = 6 to the
    * active queue.
    */
  typedef enum {
    MODIFY_SAME_ID = 0,
    WAIT_FOR_COMPLETION_OF_SAME_ID = 1
  } single_outstanding_per_id_kind_enum;

  single_outstanding_per_id_kind_enum single_outstanding_per_id_kind = WAIT_FOR_COMPLETION_OF_SAME_ID;

  /**
    * If this parameter is set, debug information is driven on the debug ports.
    * The transaction id as well as the transfer id corresponding to 
    * each beat is driven on the debug ports.
    *
    * 
    *
    * <b>type:</b> Static
    */
  bit use_debug_interface = 0; 



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checking. In a disabled state, no protocol
    * violation messages (error or warning) are issued.
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol check statistics collection. In a disabled state, statistics 
    * on checks executed are not collected. Enabling this has a run-time performance impact
    * <b>type:</b> Dynamic 
    */
  bit protocol_check_stats_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables toggle coverage.
    * Toggle Coverage gives us information on whether a bit
    * toggled from 0 to 1 and back from 1 to 0. This does not
    * indicate that every value of a multi-bit vector was seen, but
    * measures if individual bits of a multi-bit vector toggled.
    * This coverage gives information on whether a system is connected
    * properly or not.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit toggle_coverage_enable = 1;
  `else
  bit toggle_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables state coverage of signals.
    * State Coverage covers all possible states of a signal.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit state_coverage_enable = 1;
  `else
  bit state_coverage_enable = 0;
  `endif


  /** @cond PRIVATE */
  /**
    * Enables meta coverage of signals.
    * This covers second-order coverage data such as valid-ready
    * delays.
    * <br>
    * This parameter is not supported currently. The meta coverage is enabled
    * using port configuration parameter #transaction_coverage_enable.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit meta_coverage_enable = 1;
  `else
  bit meta_coverage_enable = 0;
  `endif

  /** @endcond */

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables transaction level coverage. This parameter also enables delay
    * coverage. Delay coverage is coverage on various delays between valid & ready signals.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit transaction_coverage_enable = 1;
  `else
  bit transaction_coverage_enable = 0;
  `endif
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checks coverage. 
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit protocol_checks_coverage_enable = 1;
  `else
  bit protocol_checks_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables positive or negative protocol checks coverage. 
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables signal valid check during reset when protocol_checks_enable=1. 
    * When set to '1', enables signal valid check during reset.
    * When set to '0', disables signal valid check during reset. In a disabled
    * state, no signal valid check during reset violation messages (error or warning) are issued.
    * <b>type:</b> Static 
    */
  bit signal_valid_during_reset_checks_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid. 
    * <b>type:</b> Static 
    */
  int cov_same_id_in_outstanding_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Set of multiple ID values used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_multiple_same_arid and 
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid. 
    * <b>type:</b> Static 
    */
  int cov_multi_same_ids[];

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching back to back write transactions for
    * covergroups trans_master_ace_lite_coherent_and_ace_snoop_response_association_with_specific_id. 
    * <b>type:</b> Static 
    */
  int cov_specific_id_in_back_to_back_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables valid_ready_dependency_coverage 
    * <b>type:</b> Static 
    */
  // When valid_ready_dependency_coverage_enable is set to '1' for IUS simulator
  // the function cov_sample_``dependency () of svt_axi_port_monitor_def_cov_util.svi
  // consumes around 10x more time. So because of this, the default value is kept 0 for the IUS simulator.
  // valid_ready_dependency covergroups as performance intensive and hence diabling them by default.
`ifndef INCA
  bit valid_ready_dependency_coverage_enable= 0;
`else 
  bit valid_ready_dependency_coverage_enable= 0;
`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid  need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */ 
  int cov_num_clks_awready_and_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_wvalid_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_bready_dependency  = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroups
    * trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_write_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins each for 
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_awid
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_snoop_xacts.It should be programmed to 
    * a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_snoop_xact which
    * indicates the number of outstanding snoop transactions VIP can support.
    *
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_snoop_xact
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_snoop_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_read_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid 
    * <b>type:</b> Static 
    */
  int cov_bins_dvm_tlbi_num_outstanding_xacts = 64;  

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding DVM TLBI transactions for
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid. 
    * <b>type:</b> Static    
    */
  int cov_same_id_in_dvm_tlbi_outstanding_xacts = 0;  
  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates if user wants to cover all the id_ranges of the outstanding
    * transactions. BY default , Only fixed number of outstanding transactions will be covered 
    * <b>type:</b> Static 
    */
  bit cov_num_outstanding_xacts_range_enable = 0;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awaddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and bresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and araddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and rresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_rresp_enable = 1;
    /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,rresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_rresp_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,bresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_bresp_enable = 1;



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen, awaddr and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awlock_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst,
    * arlen, araddr and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arlock_enable = 1;

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type,atomic_xact_op_type,awsize
    * and awburst signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_comp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , atomic xact op type , awburst
    * and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_noncomp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , bresp and
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_bresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type ,bresp
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_bresp_burst_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type 
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write transaction type , awmmussid and
    * and awmmusecsid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmusecsid_awmmussid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write_xact_type , awmmussidv and awmmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmussidv_awmmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type,armmusecsid and armmusid signal.
    * <b>type:</b> Static 
    */
bit trans_cross_read_xact_type_armmusecsid_armmusid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type , armmussidv
    * and armmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_read_xact_type_armmussidv_armmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_nid
    * and stash_nid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_nid_stashnid_valid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_lpid
    * and stash_lpid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_lpid_stashlpid_valid_enable = 1;

`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awqos_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and 
    * arqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arqos_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * bresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop, awdomain 
    * and bresp signal.
    * The EXOKAY response is permitted for WriteNoSnoop for NONSHAREABLE and SYSTEMSHAREABLE domains. 
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awsnoop_awdomain_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain and awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awbar_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * araddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_coh_rresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain and arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_arcache_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arbar_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between ardvmmessage and 
    * ardvmresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_ardvmmessage_ardvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acprot signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * ace rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_crresp_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acdvmmessages
    * and acdvmresp.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acdvmmessage_acdvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_read_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_write_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level meta coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi4_stream_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level delay coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_axi4_stream_delay_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_read_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_write_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI STREAM transaction level coverage group for cross coverage
    * between stream transaction type, tid and tdest.
    * <b>type:</b> Static 
    */
  bit trans_cross_stream_xact_type_tid_tdest_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for axi outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_outstanding_xact_enable = 1;
  
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_outstanding_xact coverage group for
    * axi barrier outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_outstanding_xact_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_pair_sequence coverage group for
    * read and write barrier pair transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_pair_sequence_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_non_barrier_xact_after_256_outstanding_barrier_xact coverage group
    * <b>type:</b> Static 
    */
  bit trans_non_barrier_xact_after_256_outstanding_barrier_xact_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_read_burst_sequence coverage group for
    * back to back read pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_read_burst_sequence_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_write_burst_sequence coverage group for
    * back to back write pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_write_burst_sequence_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_same_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with same ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_same_id_completed_out_of_order_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_diff_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with diff ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_diff_id_completed_out_of_order_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width48 ,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width40,trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_tlbinvl_modes_virtaddr_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width48  ,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width40,trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_branch_predictor_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for  trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_phy_inst_cache_invl_modes_modes_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width32
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_virt_inst_cache_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_addr_range_width48,
    * trans_cross_ace_dvm_firstpart_addr_range_width40,trans_cross_ace_dvm_firstpart_addr_range_width32,
    * trans_cross_ace_dvm_firstpart_addr_range_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_addr_range_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_secondpart_addr_range_width65,
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range56,trans_cross_ace_dvm_firstpart_secondpart_addr_range32
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_secondpart_addr_range_cov_enable = 1;
  
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_state_RD_WR_burst_sequence coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_four_state_rd_wr_burst_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_excl_normal_sequence coverage group
    * This cover group covers specific combinations of exclusive and normal transactions
    * <b>type:</b> Static 
    */

  bit trans_axi_four_excl_normal_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_lock_followed_by_excl_sequence coverage group
    * <b>type:</b> Static 
    */
  bit trans_lock_followed_by_excl_sequence_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_fixed_burst_wstrb coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_fixed_burst_wstrb_cov_enable = 1; 
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer coverage group 
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_cov_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_wstrb_to_signal_unaligned_start_address coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_wstrb_to_signal_unaligned_start_address_cov_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_same_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_same_arid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_diff_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_cache_modifiable_bit_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_same_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_same_awid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_diff_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_cache_modifiable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_multiple_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_awid_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_awid_enable = 1;

 
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_snoop_xacts coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_snoop_xacts_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_enable = 1;  
/**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_enable = 1;  

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_arcache coverage group
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_atomictype_exclusive_arcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_awcache  coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_atomictype_exclusive_awcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awsnoop_awdomain_awprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_writeunique_awdomain_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables cross coverage of  transaction parameters with slave port_id for
    * the following covergroups.
    * - trans_cross_ace_awsnoop_awsize
    * - trans_cross_ace_arsnoop_arsize
    * - trans_cross_ace_awsnoop_awlen
    * - trans_cross_ace_arsnoop_arlen
    * - trans_cross_ace_awsnoop_awdomain
    * - trans_cross_ace_arsnoop_ardomain
    * - trans_cross_ace_awsnoop_awcache
    * - trans_cross_ace_arsnoop_arcache
    * - trans_cross_ace_awsnoop_awburst
    * - trans_cross_ace_arsnoop_arburst
    * - trans_cross_ace_awsnoop_bresp
    * - trans_cross_ace_arsnoop_coh_rresp
    * Basically, it covers if the transaction properties have been covered from the master to all the different slaves
    * .
    * <b>type:</b> Static 
    */
  bit cov_trans_cross_slave_port_id_enable = 0;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arsnoop_ardomain_arprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_readonce_ardomain_arprot_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awprot_awbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_awprot_awbarrier_memory_sync_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arprot_arbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_arprot_arbarrier_memory_sync_enable = 1;
      
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write strobes 
    * <b>type:</b> Static 
    */  
  bit trans_cross_axi_write_strobes_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_narrow_transfer_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_narrow_transfer_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction coverage group for master_to_slave_path_access
    * <b>type:</b> Static 
    */
  bit trans_cross_master_to_slave_path_access_cov_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_enable = 1;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_coherent_and_ace_snoop_response_association_enable = 1;  
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id_enable = 1;

  /** @cond PRIVATE */
   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, for non monifiable transaction cache_type 
    * and prot_type fields are compared.
    * By default this configuration parameter is set to 1 to enable cache_type and prot_type comparation,
    * if this parameter is set 0 then cache_type and prot_type comparations are dissabled
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit master_slave_xact_association_cache_prot_check_enable = 1;
  /** @endcond */

   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, cache_type[3:1] and prot_type fields are compared.
    * By default this configuration parameter is set to SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK
    * to enable cache_type and prot_type comparation for non modifiable transaction,
    * if this parameter is set SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK
    * it enables cache_type and prot_type comparation for modifiable and non modifiable transactions,
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  master_slave_xact_association_cache_prot_check_enum master_slave_xact_association_cache_prot_check = SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for snoop transfer
    * <b>type:</b> Static 
    */
  bit trans_axi_snoop_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_read_with_same_id_to_different_slaves_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_arsnoop_acsnoop 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_arsnoop_acsnoop_enable =1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_enable =1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_enable =1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_write_with_same_id_to_different_slaves_enable = 1;
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transactions on
    * AR, AW channel waiting for snoop response
    * <b>type:</b> Static 
    */
  bit trans_ar_aw_stalled_for_ac_channel_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after nonshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_nonshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after innershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_innershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after outershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_outershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after systemshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_systemshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction ordering
    * after barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_ordering_after_barrier_enable = 1;

  /**
    * Determines if the transaction trace file generation is enabled.
    * 
    * - 1'b1 : Enable trace file generation. 
    * - 1'b0 : Disable trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_tracing = 1'b0;

   /**
    * Determines if transaction reporting is enabled.
    * 
    * - 1'b1 : Enable transaction reporting.
    * - 1'b0 : Disable transaction reporting. 
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_reporting = 1'b0;

  /**
    * Applicable only when enable_tracing or enable_reporting is set.
    * Determines if transaction data should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data in trace file generation. 
    * - 1'b0 : Disable data in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_trace_enable = 1'b0;
  
  /**
    * Applicable only when enable_tracing or enable_reporting and data_trace_enable is set.
    * Determines if transaction data_beat should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data_beat in trace file generation. 
    * - 1'b0 : Disable data_beat in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_beat_trace_enable = 1'b0;

  /** 
    * @groupname protocol_analyzer
    * Determines if XML generation is enabled.
    * <b>type:</b> Static
    */
  bit enable_xml_gen = 0;

  /**
   * @groupname protocol_analyzer
   * Indicates whether XML generation is included for memcore operations. The resulting
   * file can be loaded in Protocol Analyzer to obtain a graphical presenation of the
   * memcore activity. Set the value to 1 to enable the memcore XML generation.
   * Set the value to 0 to disable the memcore XML generation.
   * 
   * <b>type:</b> Static
   */
  bit enable_memcore_xml_gen = 0;
 
  /**
   * Determines in which format the file should write the transaction data.
   * The enum value svt_xml_writer::XML indicates XML format, 
   * svt_xml_writer::FSDB indicates FSDB format and 
   * svt_xml_writer::BOTH indicates both XML and FSDB formats.
   */
  svt_xml_writer::format_type_enum pa_format_type ;
  
  
  // **********************************************
  // Configuration parameters for STREAM interface
  // **********************************************
  /** @cond PRIVATE */
  /** 
    * Signifies the presense of the TREADY signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tready_enable               = 1;

  /** 
    * Signifies the presense of the TKEEP signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tkeep_enable                = 1;

  /** @endcond */

  /** 
    * Signifies the presense of the TSTRB signal in the VIP. 
    * <b>type:</b> Static
    * Value of tstrb is consider as 0 when tstrb_enable = 0.
    */
  rand bit tstrb_enable                = 1;

  /** 
    * Signifies the presense of the TID signal in the VIP. 
    * <b>type:</b> Static
    * Value of tid is consider as 0 when tid_enable = 0.
    */
  rand bit tid_enable                  = 1;

  /** 
    * Signifies the presense of the TDEST signal in the VIP. 
    * <b>type:</b> Static
    * Value of tdest is consider as 0 when tdest_enable = 0.
    */
  rand bit tdest_enable                = 1;

  /** 
    * Signifies the presense of the TUSER signal in the VIP. 
    * <b>type:</b> Static
    * Value of tuser is consider as 0 when tuser_enable = 0.
    */
  rand bit tuser_enable                = 1;

  /** 
    * Signifies the presense of the TDATA signal in the VIP. 
    * <b>type:</b> Static
    * Value of data is consider as 0 when tdata_enable = 0. If TDATA is not present it is required that TSTRB is not present
    */
  rand bit tdata_enable                = 1;

  /** 
    * Signifies the presense of the TLAST signal in the VIP. 
    * <b>type:</b> Static
    * All transfers are considered as individual packets when tlast_enable = 0.
    */
  rand bit tlast_enable                = 1;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDATA signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tdata_width                 = `SVT_AXI_MAX_TDATA_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tid_width                   = `SVT_AXI_MAX_TID_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDEST signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tdest_width                 = `SVT_AXI_MAX_TDEST_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TUSER signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tuser_width                 = `SVT_AXI_MAX_TUSER_WIDTH;

  /** @cond PRIVATE */
  /** Setting this parameter to 1, enables the generation of a
    * byte stream type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit byte_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_aligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous un-aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_unaligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * a sparse type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit sparse_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of user defined 
    * streams.
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit user_stream_enable = 1;
  /** @endcond */

  /**
    * Specifies the number of stream transactions that can be interleaved.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted streams beyond this value.
    * SLAVE: 
    * Checks that received streams are not interleaved beyond this value. 
    * An error is issued if streams are interleaved beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int stream_interleave_depth       = `SVT_AXI_MAX_STREAM_INTERLEAVE_DEPTH;

  // **********************************************
  // End of Configuration parameters for STREAM interface
  // **********************************************

  /** 
    * @groupname default_ready
    * Default value of AWREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_awready = 1;

  /** 
    * @groupname default_ready
    * Default value of WREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_wready = 1; 

  /** 
    * @groupname default_ready
    * Default value of ARREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_arready = 1;

   /** 
    * @groupname default_ready
    * Default value of RREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_rready = 1;

  /** 
    * @groupname default_ready
    * Default value of BREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_bready = 1;

  /**
    * @groupname default_ready
    * Default value of ACREADY signal.
    * Applicable when axi_interface_type is ACE.
    * <b>type:</b> Dynamic 
    */
  rand bit default_acready = 1;

  /**
    * @groupname default_ready
    * Default value of CRREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_crready = 1;  
 
  /**
    * @groupname default_ready
    * Default value of CDREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_cdready = 1;

  /**
    * @groupname default_ready
    * Default value of TREADY signal.
    * Applicable when axi_interface_type is AXI4_STREAM.
    * <b>type:</b> Dynamic 
    */
  rand bit default_tready = 0;

  /** 
    * @groupname default_ready
    * Default value of QVN VxREADY signal. 
    * <b>type:</b> Dynamic
    */
  `ifdef SVT_AXI_QVN_ENABLE
  rand bit default_qvn_ready = 1;
  `endif

  /** 
    * @groupname axi_signal_inactive_wdata_byte_value
    * When the VALID signal of the write data channel is high and wstrb is low, all
    * inactive wdata byte lane will take this value and valid wdata remains in the 
    * active byte lane.
    * <b>type:</b> Dynamic 
    */
  rand wdata_val_enum inactive_wdata_bytes_val = INACTIVE_WDATA_BYTE_UNCHANGED_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_addr_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_PREV_VAL;
`else
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_X_VAL ;
`endif
  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum read_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write response channel is low, all other 
    * signals (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum write_resp_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * Enables toggling of ready signals when corresponding valid is low
    * The exact manner in which the ready signals are toggled depends on
    * the values set in svt_axi_transaction::idle_addr_ready_delay,
    * svt_axi_transaction::idle_wready_delay, svt_axi_transaction::idle_rready_delay
    * and svt_axi_transaction::idle_bready_delay
    * <b>type:</b> Static 
    */
  rand bit toggle_ready_signals_during_idle_period = 0;
 
  /** @cond PRIVATE */
  /** If this parameter is set, the master checks for any outstanding 
    * transaction with an overlapping address before sending a transaction.
    * If there is any such outstanding transaction, the master will wait
    * for it to complete before sending a transaction.
    * <b>type:</b> Static 
    *
    * This parameter is not yet supported.
    */
  rand bit addr_overlap_check_enable = 0;
  /** @endcond */

  /** 
    * @groupname axi3_4_config
    * The number of addresses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a read ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int read_data_reordering_depth = 1;
`else
  rand int read_data_reordering_depth = 16;
`endif

   /** 
    * @groupname axi3_4_config
    * The number of responses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a write resp ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
  rand int write_resp_reordering_depth = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of beats of read data that must stay 
    * together before it can be interleaved with read data from a
    * different transaction.
    * When set to 0, interleaving is not allowed.
    * When set to 1, there is no restriction on interleaving.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_INTERLEAVE_SIZE 
    * <b>type:</b> Static 
    */
  rand int read_data_interleave_size = 0;

  /**
   * @groupname axi3_4_config
   * Specifies how the reordering depth of transactions moves.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_window_enum reordering_window = MOVING;
      
  /**
   * @groupname axi3_4_config
   * Specifies the reordering algorithm used for reordering the 
   * transactions or responses.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_algorithm_enum reordering_algorithm = ROUND_ROBIN;
  
  /** 
    * @groupname axi3_4_config
    * This parameter is added to control the reordering priority, in which svt_axi_transaction::reordering_priority 
    * value Vs reordering priority scheme.
    *
    * This member is applicable only when svt_axi_port_configuration::reordering_algorithm
    * is svt_axi_port_configuration::PRIORITIZED.
    *
    * If this bit is set to ‘1’ then transactions with svt_axi_transaction::reordering_priority highest value 
    * for this attribute will get higher priority.
    *
    * If this bit is set to ‘0’ then transactions with svt_axi_transaction::reordering_priority least value 
    * for this attribute will get higher priority.
    *
    * Default value of this bit is set to ‘0’.
    *
    * Applicable for ACTIVE SLAVE only.
    *
    * Configuration type: Static
    */
  rand bit reordering_priority_high_value = 0;

  /** 
    * @groupname axi3_4_config
    * The AXI3 protocol requires that the write response for write 
    * transactions must not be given until the clock cycle 
    * after the acceptance of the last data transfer.
    * In addition, the AXI4 protocol requires that the write response for
    * write transactions must not be given until the clock
    * cycle after address acceptance. Setting this
    * parameter to 1, enforces this second condition in AXI3
    * based systems as well. It is illegal to set this parameter to 0
    * in an AXI4 based system.
    * <b>type:</b> Static 
    */
  rand bit write_resp_wait_for_addr_accept = 1;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address to be received before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID is received.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr = 0;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address handshake to be completed before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID-AWREADY handshake is completed.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr_handshake = 0;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This parameter is added to enable the structural dependency feature.
    * User has to set this bit to 1'b1 to enable the structural dependency feature.
    */
  
  rand bit axi_slv_channel_buffers_enable  = 0;
 
  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write data buffer.
    * The default value is set to 4096.
    * This default value considers that the AMBA AXI supports maximum burst_length of 256. Since the default value of axi_wr_addr_buffer is 16, a value of 256*16 is reasonable 
   */
  
  rand integer axi_wr_data_buffer = 4096;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write response buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_resp_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_rd_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read response buffer.
    * The default value is set to 4096.
    */
  
  rand integer axi_rd_resp_buffer = 4096;

  /** 
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * Number of FIFO memories to be configured for this port.
    * Each FIFO memory has a specifc address and is given in
    * #fifo_mem_addresses. Needs to be used in conjunction with
    * svt_axi_slave_memory_sequence for UVM/OVM. For VMM, #generator_type must
    * be set to MEMORY_RESPONSE_GEN. If there is a FIXED type burst access
    * to one of these addresses, then data is written/read in the corresponding
    * FIFO. If there is a FIXED type burst access to an address that is not
    * configured in fifo_mem_addresses, a SLVERR response is issued.  If there
    * is a FIFO underrun when a READ is issued, a SLVERR is given as response
    * <b>type:</b> Static 
    */
  int num_fifo_mem = 0;

  /**
    * @groupname axi3_4_config
    * Addresses corresponding to each FIFO
    * The size of this array should be equal to #num_fifo_mem
    * <b>type:</b> Static 
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] fifo_mem_addresses[];
  
  /** @cond PRIVATE */
  /**
    * The AXI slave currently supports two types of memory:
    * 1. A legacy SV based memory. This is the solution by default. For more information refer to the class reference documentation of svt_mem.
    * 2. A C based memory which has more features compared to the SV based memory. For more information refer to the class reference documentation of svt_mem_core. 
    * If the memory type is set to this, the following needs to be done:
    * a. Pass/include (as elaboration options to vcs/mti/nc) “${DESIGNWARE_HOME}/vip/svt/common/latest/C/lib/${platform}/libmemserver.so"
    * b. Set LD_LIBRARY_PATH as $DESIGNWARE_HOME/vip/svt/common/latest/C/lib/$platform (or prescript file if using dw_home build)
    */
  mem_type_enum mem_type = SV_BASED_SVT_MEM;
  /** @endcond */

  /** @cond PRIVATE */
  /** 
    * Enables the internal memory of the slave.
    * Write data is written into the internal memory and read
    * data is driven based on the contents of the memory.
    *
    * <b>type:</b> Static
    *
    * This parameter is not yet supported. The slave supports built-in memory,
    * but this parameter is not currently required to enable the memory.
    */
  bit enable_mem = 1;
  /** @endcond */

  /**
    * Enables address generation based on the values configured
    * in {nonshareable_start_addr,nonshareable_end_addr},
    * {innershareable_start_addr,innershareable_start_addr} and
    * {outershareable_start_addr,outershareable_end_addr} which are set
    * through svt_axi_system_configuration::create_new_domain() and
    * svt_axi_system_configuration::set_addr_for_domain().
    * This establishes a relationship between the addresses (svt_axi_transaction::addr)
    * and domain_types(svt_axi_transaction::domain_type) generated in a transaction.
    */
  bit enable_domain_based_addr_gen = 0;

  /**
    * An array of start addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_end_addr to form an address range applicable
    * to a nonshareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_start_addr[];

  /**
    * An array of end addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_start_addr to form an address range applicable
    * to a nonshareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_end_addr[];

  /**
    * An array of start addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_end_addr to form an address range applicable
    * to a innershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_start_addr to form an address range applicable
    * to a innershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_end_addr[];

  /**
    * An array of start addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_end_addr to form an address range applicable
    * to a outershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_start_addr to form an address range applicable
    * to a outershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_end_addr[];

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the protection type (as indicated by
   * svt_axi_transaction::prot_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the protection type properties recorded in the cache are set
   * for the auto-generated transaction
    */
  bit update_cache_for_prot_type = 0;

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the memory attributes(as indicated by
   * svt_axi_transaction::cache_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the memory attributes recorded in the cache are set for the
   * auto-generated transaction
    */
  bit update_cache_for_memory_attributes = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * the cache must be updated for WRITENOSNOOP and READNOSNOOP transactions.
    * Currently supported only if  cache_line_state_change_type is set to
    * RECOMMENDED_CACHE_LINE_STATE_CHANGE. Cache is updated only if
    * transactions are a full cacheline access. Transactions with sparse write
    * strobes are also allowed. If transactions with partial or multiple
    * cacheline accesses are received by the master driver, existing entries in
    * the cache for the corresponding address(s) will be deleted. If this bit
    * is set and svt_axi_transaction::force_xact_to_cache_line_size is set, a
    * constraint in the master transaction forces all WRITENOSNOOP and
    * READNOSNOOP to be of a full cacheline access and FIXED types bursts are
    * not allowed. The specification allows a cacheline to move from the
    * invalid state to a valid state only for a full cacheline access.
    * Therefore any backdoor access to the cache to write into non-shareable
    * region must write into all bytes of the cacheline. For a WRITENOSNOOP
    * transaction, if the cacheline is dirty and a transaction with partial
    * write strobes is received, the VIP merges dirty data from the cache and
    * the data in the transaction and transmits it. If the cacheline is clean,
    * no merging of data is performed. If the cacheline does not exist,
    * allocations are not made for a WRITENOSNOOP transaction based on section
    * C4.8.1 and Table C4-20 of the specification, since there are no cacheline
    * state transitions from an invalid state to a valid state. Hence, a
    * WRITENOSNOOP will modify cache contents only if the cache is already
    * allocated either through a READNOSNOOP or through backdoor access of
    * cache. For a READNOSNOOP transaction, if there is no entry in the cache,
    * a new cacheline is allocated only if
    * svt_axi_transaction::allocate_in_cache is set. If there is already an
    * entry in the cache, the status of the cache is updated, but the data is
    * not because this indicates a speculative read and the data in cache may
    * be the latest copy.  Cacheline state transitions for READNOSNOOP
    * transactions correspond to section C4.5.1 of the specification. 
    */
  bit update_cache_for_non_coherent_xacts = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * data must always be supplied for READONCE, READCLEAN, READSHARED,
    * READNOTSHAREDDIRTY and READUNIQUE snoop transactions on the snoop data
    * channel if the cacheline is in a valid state. If this value is set to 0, data may or may not be transferred based on randomization
    */
  bit transfer_snoop_data_always_if_valid_cacheline = 1;

    /** 
    * @groupname axi3_4_config
    * If this bit is set to ‘1’ then transactions are only eligible for "write_resp_chan_lock" only after 
    * both address phase and data phase are completed.
    *
    * If this bit is set to ‘0’ then transactions  are eligible for “write_resp_chan_lock” after
    * Address phase is completed.In here "data phase" is not considered. 
    * 
    * Default value is ‘0’.
    * This attribute is applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
    *
    * ** Note, Eligible transaction are given the “write_resp_chan_lock” according to the “reordering algorithm”.
    */
  bit write_resp_wait_for_data_accept = 0;

  /** @cond PRIVATE */
`ifdef SVT_VMM_TECHNOLOGY
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals spcified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * <b>type:</b> Dynamic
    */
`else
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals specified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also, min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * When set to -1, svt_axi_port_perf_status::start_performance_monitoring() and
    * svt_axi_port_perf_status::stop_performance_monitoring() needs to be used to
    * indicate the start and stop events for the performance monitoring. If the
    * start and stop events are not indicated, the performance monitoring will not 
    * be enabled. If the stop event is not indicated after issuing a start event,
    * the port monitor stops the performance monitoring in the extract phase.
    * Note that any constraint checks will be performed only during the monitoring period.
    * <b>type:</b> Dynamic
    */
`endif  
  real perf_recording_interval = 0;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a write
    * transaction to complete. The duration is measured as the time when the
    * the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    */
  real perf_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a write transaction to
    * complete. The duration is measured as the time when the the transaction
    * is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a read
    * transaction to complete. The duration is measured as the time when the the
    * transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a read transaction to
    * complete. The duration is measured as the time when the the transaction is
    * started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis
    * Indicates if periods of transaction inactivity (ie, periods when no
    * transaction is active) must be excluded from the calculation of
    * throughput.  The throughput is measured as (number of bytes transferred
    * in an interval)/(duration of interval). If this bit is set, inactive
    * periods will be deducted from the duration of the interval
    */
  bit perf_exclude_inactive_periods_for_throughput = 0;
  
  /**
    * @groupname axi_performance_analysis
    * Indicates how the transaction inactivity (ie, periods when no
    * transaction is active) must be estimated for the calculation of
    * throughput.  
    * Applicable only when svt_axi_port_configuration::
    * perf_exclude_inactive_periods_for_throughput is set to 1. 
    * EXCLUDE_ALL: Excludes all the inactivity. This is the default value. 
    * EXCLUDE_BEGIN_END: Excludes the inactivity only from time 0 to start of first 
    * transaction, and from end of last transaction to end of simulation. 
    */
  perf_inactivity_algorithm_type_enum perf_inactivity_algorithm_type = EXCLUDE_ALL;
  /** @endcond */

`ifdef SVT_ACE5_ENABLE
   /**
     * @groupname ace5_config
     *  It can be set to either of three values below:
     *  mte_support_type =svt_axi_port_configuration:STANDARD.
     *  When set to the above value memory tagging is supported on the interface, all tag operation types are supported
     *	mte_support_type = svt_axi_port_configuration:BASIC.
     *  When set to the above value memory tagging is supported on the interface at a basic level, a limited range of tag operations are supported. 
     *	mte_support_type = svt_axi_port_configuration:FALSE.
     *  When set to NOT_SUPPORTED , memory tagging is not supported on the interface
     *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
     */
  mte_support_type_enum mte_support_type = NOT_SUPPORTED;

 /**
   * @groupname ace5_config
   * Bcomp signal
   * Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   */
  bit bcomp_signal_enable; 
`endif

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname ace5_config
    * Enables unique id identifier feature for write and read address and response channels
    * <b>type:</b> Static
    * Only applicable when SVT_ACE5_ENABLE macro is defined and 
    * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 or higher
    *
    * This functionality is not supported yet.
    */
   bit unique_id_enable  = 0; 

 /**
   * @groupname ace5_config
   * Enables Read Data Chunking feature support in master and slave. 
   * <b>type:</b> Static
   * Only applicable when SVT_ACE5_ENABLE macro is defined. 
   * Not yet implemented.
   */
  bit rdata_chunking_enable = 0;

   /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunknum signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunknum_width                   = `SVT_AXI_MAX_CHUNK_NUM_WIDTH;

  /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunkstrb signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunkstrb_width                   = `SVT_AXI_MAX_CHUNK_STROBE_WIDTH;
`endif

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /*   pre_randomize does the following
   *   1) Calculates number of tagged address attributes set to '1'
   */
  extern function void pre_randomize ();

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3sRE1AICCkzyjmmbts6YxnAy5oasUehUXonhEqP4w9ojK6+bvq0ZMt/vYNUnMuaD
IvbpOSHQCJwLRvjFluAaDmtF7Im56SKAqxVaa0hbST7e2TeMrwxxtir3qyGAJigN
2Y9QDq+3cK3MK4cGnIvcpa2+erfV014D8wAHpvN36Im1fGn2IedJwg==
//pragma protect end_key_block
//pragma protect digest_block
SQbVvKJCgaEjXKNHNYGcAICFI2A=
//pragma protect end_digest_block
//pragma protect data_block
Wp92nk9J+vANtizv334ZVn+WQGswx9iIDt5ZMUo1NZwptSb+AO35nytpDukoJGy2
uWesSf0X+oCBFJmIYra+8qcJflBw+nsZQrTklEf/3sQa3xCSD2Gvu1uZrNJ/ZRMz
M1FH1yRUxATVhAKZB9Dj7YE5rrznv0PeXFwo2ivaN6GjkX6zSgCvg5UmWpVXoY/k
51xCTbaHDXj4P4dpaW0BIMbkkeHtCgK8OrVkNrEtQbvzHKSEIcm3/ghSJXwCfz/a
BwVdAmZNZ4FDKhn71WwJr1QMTeVMgk4va4vwu3xTl9KTIBi3eJSm8WhRXAYwbiLX
/63jkqudjbX0UcIQbC5eeGGwHkpBhO6ohMCqbLcdOX7aaXVhOdsITXqkqn2gaxiS
+JV+C+HOH4SZWLt/C0dmBp1PdeRr15GV4aHB2n2oa2dppdQeAp8SRRkWqlbLaA1J
d8AasVDKtwdEAdhSZBDCy0BRYrbol7zKeoSWF2/h0oi6b5yeyDMWJHhM9xIiwqqL
rAYTCvWGSFtOK/oq3i6wJ4aMUml7MidE9/XzEJzf8cuF79vGSKOavEXmFDR8hkyB
f1xjcZxe2GC0KX/1FqQeQA7miPpFIpsXQWegLC5M/DLtrPQGOu9oIGn95+oKAZX3
N2QI79G9q0mhWHYVvbxEAHyiB5YHMaqkIyPIpCtl37R4bY/33kPIdyeO6d67zpHA

//pragma protect end_data_block
//pragma protect digest_block
dDgqfRoZEOSI2tG5kV1UitbO/hg=
//pragma protect end_digest_block
//pragma protect end_protected

`ifdef SVT_ACE5_ENABLE
/** 
 * Returns 1 if bcomp response is applicable on this port else returns 0
 */
 extern function bit is_bcomp_response_valid();   
`endif

`ifdef SVT_VMM_TECHNOLOGY
/** @cond PRIVATE */
  /** 
    * @groupname axi_generic_config
    * The source for the stimulus that is connected to the transactor.
    * This member is not used.
    * Configuration type: Static
    */
  generator_type_enum snoop_generator_type = SCENARIO_GEN;
/** @endcond */
`endif

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GDZ9kV0XjOPvK0sddtIlelE7Z2X1GREQD4FJVzpKo1uoy87/zDZkOdLopzoWUCyF
PRFMytu10Pcb8RONXdHKk0txGiSbD34q1hRrqAw2MFDhsXu7vLeGbEdUM9Jgay4e
R1M2A53+r0ueNQKC6C5Jo/WAM54wGcQfWspKawNXlok//IUdI9CC7Q==
//pragma protect end_key_block
//pragma protect digest_block
DFzHPEojtZS+RHrU9hULLsI8Lfk=
//pragma protect end_digest_block
//pragma protect data_block
p1eLFBbCZ7womsonv81LUHTVQdIEwURdmdUynx/Bryz4Czq6/YjQtnUQLlaeFZ8B
4R6zYHwqO7h/jdqZbHm3fGCCxJ1rH4cSzrDj2YiFboTCT/VYpxdhiU0sSrmWwblS
aCazVfV0vUmkkL/6cFA7GoubRGEoQz8YpPc+1g/3ffMvq/dp1MW7GxLZ+nGtikC9
O9FZ7Ffo7w7cp0llyiQ3ja5Bgo6x4Z/C/mIXV3eYBAUmYSdByj6G/uyTMKo53wNP
86fngkARfVy9fXhT5726g5DQa2oYGyO95EE+upxuMIgWIdPKzS7JJsffOj89Dp9m
61DAO0H2yRq9raBEbTsTfSpSQoEGmFe/5UzG6lMnpF/cTiOfg3r014oyw7NHzZw/
xhb/skzK/cQLFOAnagF+NpQ6Rz630BNZ+t7gV2XGddAIuoEaLgQyMgIUKPXWMUUh
seDWQPdY+npjWYlEZeppWxNizphDNyMTwx6slYyTIR6eZkuyV+ychdq3MUgqrHLo
TavJwKonEdlFBAQYUqZV/2giukCbTv7aluChMMK6jJcWzq4jXxvodfyoVAbZfZSB
cw0Mt8izP9CD3zAD3d4/Pd8CWz09VFMwT/ULsBD6ASuQ26fIoJNVvZ122BAKghzg
bio6/Pcb0TTZqIyIg5EPIhoVcDA4Y/RkR351qimmmCWrRZ7mkYf3czmWjYE8WM/E
KRnQ7loUJcmaqm9iOJehCas3U3pQ2Miw2DoJ7rTiG9yr2eUt6sTeuKzZT6OeKvP5
peiarmUxS+mVPVavIu1MjYcZ2NT/1kk6e4T1W0X6LrDrvoG5M58KutEFVhmwPOwK
4Un+cZXd01ia6YaGHHKqrQBKkECEm0u9Rf70kc+CsyoHbpMansqqo5Dvw3elRnT2
8aGAJKyZuiajbDOMX8atbV3AZ9wogKTu8ELXdP3VFXeMZJ6tozaXGqZcS2ByPYJI
MTVn312N/8LOaMcRUuO8AQfx99Ai1o+7kFhXjJdfaw4QmlIS7KIbzmsiisLt6ABA
vhhJ02EW8MXFC3Qe/DY5Zzuu0OP4ihVOJWO3i0F/Uig2zDaKRpiDIAvMHux+/+4U
bApQ56bwsKx4y3xrfWZACjfKtHNq5fmuHOZ4wKwKc9XtN5mJvjNrRd4mz9LhEK5L
uZ9ljshyUO5UuLVN8S6dpAu9ICnfg7VX4ke/3w9THMsRJ+HEUPiY7+L0p7vp2Q5N
QauB5Ve1uwy+kbU1xvvKgplkJhje84I26DgVG+qcj2tmPmgLPGsKoE1XzGQkCL/Z
PfuGp9WqHJjIWWuScfEPGT+nWGZ4k6/TEydHkXnLQ4qshtfncUcTnJG0dzvCI+ar
vYdvZNJwlW0O74H/iwcBEIxWITdBjQSFL8P9LyF0CoWUm/I/8zWx8eJujLPFeqon
I5jwlTWtBodKSWV0dLz/Kc19xADXewO3yVLm2ysQzhWYy4VySA1Iq4p3nnUd5xQc
HMcxPb9FTOL8adE9G8UWdr7WZgNIhda4gBErGh7cKcpD5MUeYoUlc+cIgTqNcDSD
LrUidA+WJCzGWu7q8B0cC6IbTPlzYARpYrgACafZQCK2GAuXGMM3YWxdgaGhlp8D
7ukDMlVfsMVAoFRLvn5uwanihqr4QzZxDTreD8et9i61wzpJe8nFrAZKkQT61WdZ
6Rf6NVFcP/a+6ORZphzdjxmbZ/3Rr+VNNGe+X25uGaox75d8Ugzl8pheB9VBQMwr
NnYoQPrRAXGI+H4NJC3B2ai37GdL5VgzWS4mFxHfa6u2QGESEdf/vSMqGMzQ+wXJ
1q1p9S3sqz+qfuhEdtjEtQDAdSqkRjKpbc7ok/QDB3gyFm0moRjsALbqmTujUQb/
2ptRZdWboaNfasOj5O2KbOFH7TwvVjr8NJhwKcqvQ2jw5MnbKJU6Pq0k4UOFVfbz
BC9ZSpL6VinMGbboP7xwb91Kna+eklWnw1XmrB7mG4hJOgNe8ZBTVtFGVNn8TkPP
x/kOOKq3arByEVwlEyGhaQ3bFtBRe+I1fuCjEa+21c+JAJgw0P9W8A+5Lj0nr1fY
+JvdhD4b+LSBLJ9mUyv20I0+zPIET9zFHTpN7qNqgRhQDhSCKjZE8+FlOdxWuOxk
ZqazExDH34U2kGcga7LobS70xsaVvKw7atlzZz0qEuWHZPphqrXothEIlijXEwUD
1xhtkHSupjPglraaahq42Usptc5K63aFJ3fDASYq7HbRBhwHw6MfAlYWMz6eJuwG
1YHomqGZ7iiZ3Q0UT4IqKxr1en+VVbvqYVjAvN0DXz6RquYuGD3MZWT/P/5ud5k7
QLF7V7Bm5X+NmRIJ8AquFD9GE9VuGQkyH4rY+bVDf19JAtOWnu6mkDwGjFSpxFc4
H6imDPgdJS+Tstc82l69Xy60t9KMB0Y0vhso+pL8tZSSCMlv+mheKQnyZOvmHg+8
NiBCK7NcOB/KY6ggI81vvdOMewY/wLLchhlM1B9icYOiYiYvOouT4d69rTAzzSqJ
ptXe8/gDeJV9kA03AWPd2CjbcRanYf0kyfNvrWqte5Z8az41fZX0SHdAvK9Z2ucN
9Y4OdPjLbrO35kwgWNSzTCuoEnNzkJuBG1ZB1gkshxxm2YRMfKVQi8NOmj58qEdX
zHvsoIPAtB9k3qYAHABBJBpLTPWO4Bjg9XsuOMOcVt45uMqZ6aRTfMBlxvFufP9v
tooiEfbEzBWWzGvCEASsGFvFzaMGKkSdDPbGtL/r8Q7R8ItQ0DIM0lbmhBGyftG3
wGPJkxbE7tJwQ9s6lwLxeD+Bsebfc2JOTr7cwlwP3WMAaN6eABkH+JSxj6tuEHu6
g+TUA4VlU3cGZ2Kz/QiTIymarTZzfkMEomTjvaQ85e7xhyhLrmPlbqCkgbE5Rb18
Ytp3uZk19eqS9JGRck4+xKU7AMcESDcSyhX6tqbTvFAdGatwGcup3k/th2LDmufb
0nMv33u2mtrHX0AP0axLWa5sirH7BwdM2dZh/Rt8LgZBKHXq/FrnHrBNNZ0ZI/tm
gMQQM74GxGkWAWTcbBKnQKnIWZClaXFlw2ZTqoF81SlHZk66EIBWaJwsZ+CWuovI
5bSivHN7wICjMaAswLbEf15Omkf3CFtIIe9+jLOUmRrzSKUV/7lVpRnKoA4LPNxc
XCKmtoxW5HYienWx7CIDFgq1Hd8RuiV6MOggNtDVLQWZYbfZQfpBIsLOUFgt+uQy
cSHeYz/kltZpKpB/g9NQDo/x0f699ebeA8c9qXWH681awJK9XsmBdH8xOqwbLpvc
DQVPKNfjDSoN7rhoThwi71/piDx4cdhcy4HyjkSDFcWOeNLP6wkZTAJRBS6Vr/qJ
hp6CrEhySxg7Btk7qzhnUcnENdRfRlwQpO3UPBTb7ExoVwoVvp1vS13K5OkJ8a0q
W71RDq5wZ3BS3YBw7v9r/j0BjBzYAZIrUAZwkaXSX49Wu/gBiAB9krgzHPQV9Za/
m4JQQTt1ggieuHxt1iEHF/tnYHt6/Yj8CUh/hOCbfo2FqNQlMcL8LufdfAude4YF
qMClwJb1p2zto4/0rSbYcQOa14fVofUvEmY0UPzoi4cq3BRFTzZwPJoZ9Abqb2qy
Ynu60oeAhurR8tkVz+YvWeccQv+TSSI6SIDY3Mpu7BeCs9A3fa4+t71EO02tRcZn
LVcJCgOuEF/LEXXHovlgQiEEuk4MbmMRPhZvw1EgpK/693V5cHA0+udMvoznps5E
HMaIpZmRKG3WkibSL2UI/XDaT3PjTHNSHDsx1VgqiP/4NHRnMGGUFT0IuUINI1MK
2l8F/ais28di/i1uzzXNOz656CVUnDVCYETihcN7kO94mVykqNyoVxFeDyavW8a6
6yiIDl5mRAKmIrhln2WEgWjtamOt+IRSaDQ4IMtIMlfW2QkBbdmW1QLQ6whW4yMa
2HmAFTPpFx6rYi+EMXLLYPE+FHDTLILXa2oj5eetji+K6o2AFKw1pY7uf0Hexf55
yn9tYjJS4llXTr0ZL15UluZFH7RSqqzZobb5W1DAT1IpAawijm/pvi7KHwukos/2
Q0jJPOtkdu8kLneLu9YcUm3+ZX+2MrgS619T8mCbcO1JOhyYblxO9KAQCpojTTQL
WbkxZ/ZjWLgX0YMHX/KUkuIO0Ujy0FWvPWNZK7IYLetBsa1LEenBMOmaoDWHI3dU
UthzHnMjqIDxBff8s2LxsvcT6qAkVJP5P1SFxOKqJr1gGJ/jvcSyXEwFPfI75o2m
yDeK1/X5TPvoAvlubuH+SEu6IL6V3aTEPdY81mAMpKw4o8O2+sba36MuSl+93+8D
de6rX+KNprzqpcNAkDf5Vf4ctcmNKkoK2VLVTfWNDPcfBZs7vomvLLVZRMCxad92
LeNTgucTrT562Qoik3q2OS+9y//QTW8an/50a5MXvMtDoV7ToI6P0Wg4+qIE7dMq
31bpVmseTXG/WxRpd78EZt6ETwUmgYko95Qht3McEaO1hnvnS/kvaT3KXd9EDeVE
YTt/Zfbtsw0E246a7IQLqxxU9UamzxPsuRJmlWtDwtPa1eb3/8XGffugTzD1uSs6
EuZq/OfGbXGylKeBDWoHvIVQrZPgRsu5mMvNFfBWWq7H4rrAvYaSrrRX29p9RAyp
O92m0SriDhO0kLQK5yGU1rhV70IWYPrtGh4tnIALp6iaCeUVG9W6MzEeSZh7sL9l
sHLXrkX78dj8rcojNlTTT3LpOtjvsIIfNx6cqeJmqi2dc33Pnv6zMxfUJKa0tR71
HXOWzm3kml7Y/NfSDEmG6CRAEjAaNy2qvQlpcuR3+q6ZOe1j3DqqkHJGATxrKYo2
YUo+9PlEjoTRrVQkSDidV4TxNL2tCKAnkdDXJMZ6e4ln/jQJSDZQhlXg78iB7q6E
mImACsKglvvoWNqxsG3hsCHW1YIkX7bMssSU77eQE8zBZRceAD4BY6WjVjGXgp4C
EjiCxa0t1bu6JErVpQ5LPHVDzzAhkdOaYbIT9Z1rk0rnrWAlNjVzm/SCeHpP03Nw
t9rZmEz0PfYB7hmnbO7TnrkNmcAIvNWSGN6qbeG212hjo30F5rY7i8/9IKdT2Oi6
XESkoKXPaHkVzEIUtpYh2nZ0tVOn8QlAfaaKGn+PErKesAwtFNwGIigYGvQo9h1t
scodJ5iHD/SKrY58frBMJ/WJ7BtWXBednj1t2oG+9u7Jx3djykBguhWgY2SaHoPC
T+gMkfLU6B6zzwcDrW0LHfJXwoNlOTlKWYCQyP1o7E8HdxWYjvgzKu5b/9qXvhgo
y3p+AS41H8jOWUWXALep742hKvjNTrkWZebpRdVBBZ5sXRqdnvd8191mAkERNCpQ
gz4xeC08bBZI/LpE/+3mOgDVq7AL0wfRyt/dp7FwTTwqGwydRaQKmIqAmESpo2Gr
3rLnIkmXoiNlERJ3KibYHEukMAhuQt8I4XHAIaFRMz49Rljx7rRqWHXIiEnf652Z
lx8sQdds+nIHb7sevDzQeQsGWISqrYQtTAqsLoTXwI+eIHVqe+hlOqBb0Xx2NVW5
lGsqvsAVFGk62GgcbrFEiANVuqVqOkxQM5+0bVDhd1HzgYalBDbGhlbrfS6FFig9
DFwkWELxYdQFzrft2SNCgtinNa920hvjK+u4WrIWcVC5UEbwN7/JORutW1audBgz
IL/kRl8sZ5c/EpsGSW1ex+9JyxRA20fBYtbjtEkrFCefRe8qgyY4N785U30d7Epo
ebr8xOS9NP7xaQdZUDPyZamr8NaqPfUzcgmgyRh46Cf08myyO32LnF7JfpYX92YB
tAAXuIWXCSF25fJNp5JBMoD/qcKwVyIW48C2Iu35/qoxiJoHxzThkYufzHzFMVss
n07bJm5/8BiWkf69JhoFTl93D7lbpefPgco7+6XTfBF0IkzCvqdxZGXLTwQHEhP1
WoTX7Vm3Z77DZyP9MxaxnUIbX/rveEz8f+AvcAV4Fxw32kzKXcWiX5F9trTeZWdq
VP8rb13+ExbZC3uUYYzPEAbSGg4MeTTMOUZmEw+AwlXpvLEIColbs9TPW3d7fXlM
XlMiKbynCdyclbEsZtCaGCucVNtHQfzdrSSwHaFXrTLkMx5+igwyxNp6zZviv8v2
hk5pcqS5MkG8knohz8VwwTlrUPDPDaCE8wYJHTVcmKqRRb3ZRTVVcGM9p5W1w/xg
+Z8+vUyrkGCWwU8gVSPpebnXLpio0N5m8elUJ59fTYT5D6AD10MnM4EoDf6vENAD
soacQ3E7YMrwHZWnfFPplgO2kfF89Xi6agsmOxD8MRfCrA1t4gSTjMfXdYgwSKFs
TygvV2eGdejNAsRx5hnb5dJKAnfUI975eEDWChQys0YlFXIRUVLvfZRyn3Tob2hX
C/nyddWLdYHp53/0A97OCMwcM5mfcQBDLwjh24ALpmVbRQbfT8pazm+8ZX4klDWT
CK2FezTTnxZ1RLG6izQFaTan/qOo2tqU9LH6LsbboWnygtR4EcCQRznG+AkLGr7J
ZRDzi5qOzepzvRo8yxWdccZixTSOA5N5vJ9uCig5U4OnTnUFumnfH69k9N4c3B8v
RQgIywMMus3kLu2x6EBjV9ndrpRlbIdS/QfQ0yBBZESbbs/pCjPuYFBn2vY+WQAf
1yINI5mVPNUoQvpTNHsKTSufO/fF7J/lZqsfLuheXhxobqCAP467bHUg8MnuEp79
EjXtdDchIzi6n8Vu7zg2X6HFm+LU/Hp+f6MolcW0wkOWrq/ArG17SF9sy1LshGEC
u+uA4LPB0H9w8rZlTlW7n07HjR+Hlubmrs57nea57KdOWiWvH2E5eMc4CSa7n6tP
DdsfOKKxLw0KRdUDGMir4f57nuuvHPeFcMHVC9A/YGhnqt2GvQ3JaNAZa6g1WQtj
c7slqrxri63suoe3gHVysYJ4MvyCBZVD9C2frOuSNsoyxeoyi0V8lD6KeHHC13yH
+RPxuF5cShO5quoUAoe3etaUbs8Zl5Sxrj5CrUBTGjmFvGjs0KjBjs5c5OqPxlcY
JPLwPG/A12SFftNA6QulExG/sus0dsS7B07d3zQQKcWS4U+WylJ7t30so2q1ark6
h4zFxVQtebRW5K4NzWX1xo9nqgFDqMVkhfPLT1fZpfLf1GX7B+f+CgJOcIslN8Er
jxEOz8VG+rc1v17dTEP/gd8/GbjiFQ9QQOtK+xlXzx9yR/eFAPaSbrRki2HuNXNL
vXi4z+3qr6+Tqz1ag9z7Cn55klCZp47LDgrb4d5rhfrqe5oV/S08zIpYP+2VepsH
0i+jmXevJDfF0PJAsOQwf920Vm7Abj8emtIZiNCtQ/E6FieAMQ1lNpo8Tl9/pdzf
YfQ/5f51wzpJJFg/SsDIbbQfQcp3EB8CtT+lo3npBVh2tFNzX7CTtbM9MCjHQ6ln
beFjzDTJxitFkpmxhrqG9fQfTdRkQnVEdeuqB/CxAJ0VkA2qJ8zjYax77v4YfrnG
o1v51x7zDbakp3YwinQGDWYC10U/kOG6aiucMMW/enCIKc4LQOlWxzjPOSCft0qn
scCrbTDLZIPR5HmDpSpmnMm5h1K5kuDQNGxFazsI3YhHbdNpaYmADqdWugZARbGB
TV6cMtrVVR6TP1qppLOg57fdCxD9FsOpEiGS1LRP+vQEoGx9z5Y8OWBzyXwZ0DX0
YzsBgyWPH/rF8Ajrsy9BRR7oipwJ8/uIHmAc89UjJZtnIovFphAS8t/Iev+018k/
aFnDDSMEItXkuabBPqfb2cu1mAGi+rBTYPFcUHjamfGkoqkSUL4lDcC3c4CPO4T3
7htgSIb0Iys11OQoTleXrCuH/dSuvYL8rAde9SZQ0TClz0oF+lpmOqctZLDCIx6z
JaTquspKpf34jVorMKglhQ/qQji7URvfYBLomJTLJtoYLlqZNiDn0bXJVhpPBqcz
V+tbtaDXum2iAS4RZDXBu6KqJwamG+CdlH9EoKixVgVbPb6xzCZQ+5/apvf306cG
geJj+bEpdMsyRAfsq8pZ9T20mqkDt5ZplyBSTByXOEEVKJf31v2GpSRpbvUkes6D
4CH4kqXfdW1NFRIppMZrB3WW26Ua8z6gxXj21irhYH00wPWCIV8V+qCYW2gtSwSl
kRdWnlJSh1Xfqw+0Y1NQ5QlYrVggutsKke9gSXUrBq0iBmZAy2Q8E5SEeNBa/eOK
k3cbp2LiPljKQPcQi0uGXB7HO5RxybFLV0edkazS4Ute+TNhioJ7P7KXL6I7mcIG
RK8RrPULAx3mqWmnnix5wI559REIMSW6WG12R/QOjIH06hMfp1nQYXsPI8lpPw5O
Ddmc8kfR0iRaDcau2bpqmOYtketGs75bE7VOWGyTOuLfqFk0ub4MH6H6nNl7ef2B
lVpHvHDpFE/s3z/X3118k/jBhZDG4PsPWzsnDbajIXYGKOHZbv5nbGu6TzssGPbx
fF8nugtSTUAO04g+C094ZPOmUWKKWD0B4n68Qh4PkAU6aeQUsgEBY6g2JVXaVRce
5WCvgmdEWMrxi1go0GCGbQIWJfgZWcXGLqUJ21ToEAEj41UD9ZhUX0IcjeScNT3g
MhfI+43BkON6Rq1TuvLLV1n7APL2kIMO2t6HFnzFpqDoVX1LPKGLpSLZxi6Cx/LX
P4A2fxj+Epu00VRSfuOk4ftVvu2W8mC2V09VDr/GqxMnz5sCojT/Zki2LdQmBGBa
VmPJw9bl2KFK4i8PDopgQh7VXKjCUAM/wLFKYxHG2MGSx94guS86dDmpNwSdphoR
Jzr00N3WCo24CNvu3zsuArbqfxpYmdJx4LNNO60ZiDHT4HQkBK5DXNtgeqtRm/Xs
KDknI45VpEn/MolU/vkwY3j7oDlK4tTf/TBMtm9e5ktIWHgBJGnSAPaNVOn5HKK9
4++L3Cis9Nb+4aPIXwjbzY7vxQ5cNQP4+ux1pC7sGRAmLBV7MutLWxxpjOeZ6DSv
TOOiHI+z6/O+ZfFJL/0K801o+sPn7SJO+4oi/+AV/nnzso/f24yvWX6FjcuDYOY2
dz62fwonXKhUXs/bgWXX1lyNHq6HL6IW4j+4eAu9O+yvFPNVJmISOQhZy4mIfaFX
ofWTijkZdu0NqZVV3WbkPAoh75S7ZrADqoylpnH2J4A6kC0csb5GCLUP9Y3o6mY4
AUNoUMyZ0GUkfLHvACfuF/bdXp+z5jy9PFjHxbM9nF9L+MjcB4xgySdG3HGx3nWV
5k3z88C0vPv1/wld6ZbNa5KLsJKAXuHL2anSoKSDC//pFaGFHU8G0NFRQoS3sRN/
IKrU1VW7UHt0orkVr4mszcowNrfiuTZoPOuyxs87y4wsZda/GXQGRDPM2jaMHQAK
WcTKIQC3SdTzgFMd5UXeL6PDTq/r5ywwQmuY2agvNayE4FyanJ+3XbWDB0j3dAUh
Tde+r0Sdhb1kKYMAPoG4OkhUUHRXxFjOKi2B0wrTKBIVdESXDDIeFzcfHBYRcSXw
QIQ8wALBce3cyAnre0l57ScNom7Fx5zaU8sKwpV+Eg++qUvpC3VD3PIqs53MFbek
4Z7/qcMIyMH5qHNkQpNMmttUENAaXCvz2fdDRCfHI6x9v0hWhoKDMPZdGUodZuZQ
WWoP3qQnYxoSIQq/nHbXYb7WCvO+XKNI2GpbsifBu9EN2hQRVJndWWoqj83S7mtJ
n5Jqs+3qYy7eAwFZtRec9RB2nJ8rIf/FuSrQ232nGGmz5BTiAJ38uldzFJK5DuM3
M3WK7/j8cBQI66SYNqmB75vUmNA9KXo9AGZ2k1THG5jzjGhEHqMwHMAdpLOa897l
3m4tvNQODN6ZFxu945fyfDJ2BIwi/wJEBQrLb4cDIf8z/VWN3cTelxPAGQUWeoqA
Jpi5loK92R2ymfZoO2kL0mdKbJQnBHTBsXgmXnVhZLdvg6Uw+kpWxV441EHZkxKz
OZMia42R7YdouLA0coOqMqaJoUnIsgd0OWpuRRv2Oy7h8UZqnEbs5sNphiaAzhfc
soGQYXnHZRy3bPLTT2QDOf1YT14A7rtIsBUMTZR80pR0xTZ/wpqao+QSTpyAd93K
ASx81e9Knru/O1gGagO2wOnQz4MQZ28wxf8Z8REa6hcGPSjPyiO0nvfz2zcfpx91
f8TID+Xqgz4KdAOCFvOz+24SkB46L72QgriYlXqTiafzV9xu81W08tzZjT6cr61X
2YUq2vUn0KdiZyEHXOi9jt4NDhRE1M7+D/DdxQLrgTLA8PwynyeZ1JLD3fla30XC
66tfVmGFErZYcigN8n6DZiQGpVleWPHZ6oKjtKFKv+XbPPznkM4uYYc30WhulwRL
4qHRlC614sm0jd4FV+izw5WKiCLWLVIESHrw5vj090piiPOJNAONSEG2AzEF2mrr
ijq5z12PPdK3QM0JkiVYtsG/wVpge2WV0frBbgQBlQ+aXCRdoudQQKwtlelzRunC
d65LwC981dLTfQ5QVVoPefIJJzKJidDrmimhxsPjB2CIBL0MURILS1xN/smS4Hxp
uLCzmU9l/7Y08M5lGqxln/t7OeqEBCE/z4ydpsbLWLUfEqPn+XR2acP4LcBNM4UQ
DmSO9UlSYF+Kc5k/FwlHGVePWnE7scGzRhA25WgTyfmonohWtCAFeOYHCtxJ6MmA
R4NsQ3xixq6iS2hutdhRicLIHrhxl1zt4E3VOc6OIbQKlt63WIwZ8uniz9m2stZt
jF8p43K5ACXrvtGab/9dX70hxmrQw2H0iyi0YZB+ZM0Sy5BHKpQCdFF6vzlOgHSt
3BQarVM/iV54D6frJRIxuOrtjqyudvkS5yYVmTJbML2jQ1r2P2fGpB5Etw7p/6zZ
o+n8p7fkGuWkB7o3CI6rUVywEvEVHZVMly+uy90MsrYV9wPINeJDsc8T0AY44mHv
SjSVvrOfn+XHoPWzDHhLpgs9odQGJdy4IAfn4n6G/xjNYqJ26pafQaQZnwZPeNNE
zNJCS8RvL2qsVcrYi8X6B5oqub1oMRYSeuOxKrbikSjpCTpDD4OT0nP3zunccoER
YhgW51NckE+2ROHfyn/fKjqG33iDfHf3/G7Vyp1XSCB8L874s3Ct640XbGGpmFX8
L6QJaghEF8FMatcAThUER+LvEXuz7vmeM9v03Ww+Yq3/VGSvWv6om7KykppXn5JP
DVTtGiOw7GpRwelpkzoFryO4x+DqncIxi7aX5nZ2WCIEmUsgn6yswVj+B/w4bFrt
EcPioqLiP2KfJ6J6L09y/+a2N34H/yvh7tm8hxX6k6JZyP1d4/V5z9236DEfjsjf
pfw2K1jFBDJna2Z+NLL0BO2JOM5YeveGlLs+8rQ3d8vCLW5tjuoJ+HIPSrgp0SIr
AOCvVjI88j1th5Qpy+LRT6uhgxCdR5Sy1Q+ig/0aoT+qIPI1XNpiOmEyXpEZQKAN
vgCG+6dnOh+fMHOO4vgrpBJi9gTdNS9oqrWZEllxdWIm8Sb3ZzwxBq5FVBJP3xeM
F4t63kc2/lpNJU+O17TpXpTMkQZrbj7yIBws5I6nTx4vScrebThPvZOLWFmxfVSD
bkQ4VdrQ8ojP/6XDfwYTR5q55URJQ5M57m6IBzQq43KF5ydyf9Fyf+6IecoCqLdb
6H5rFH4ANZPSgZGNeYeWtATbttOOH79yzr/qqWBxL0YCNi7IDy5nP6YR7AhxemvJ
lZDecFZ/bqqq6ErekVOros8nebSwkcVkMexPzjonbLeiKLxohtMn509WgFXDPots
R3W7u0gKJ71g04XLPNIv8yGgH4MuEIm1No3ZzGqsthUM3WigsDVED6N7eCoPS5vi
pvOcNSeIFPOwbFmhWtewr9ZsJjrIsls9ga3a28eeB4OdCm/1VkTxUyF/vdI7mVDG
NEOwe8hnVmvJk7Yj6+ISwsCF1YvTAauPejRM8MvmE+6PLb4eZdCYfV7iCD5ggI5w
ql+DoIo7Rk+qNM3pIgt3++jwFs7jZaZYzMF5uHj33mhbxt+2d5RoAGwK+0d9xVzL
gztnP53vMmpIup96eFvkFWde4et8rbpKPFoB2BbwcwzbLDYXwQb0ATyQzyF8cBw7
dNOG3JJMpsFHybzvW6TeeHMPlNgCa1lt1oX1C3jOmnAL9P5za5cFw4i7VdbLgRoc
9rp9H9Gyy1EMqGl1Gbq0Q4vpgEypBMe0gwGSaObDgXCIR4hcjZlRmca5kJRGJk33
dgBRHdOgMVIiqgghJ5CqpQhVoSktlylBbJQBeMtHvPD/jehB+a9oWEVcPXJ79Cid
jf/BPw8u5Simh0WUrA/zrr3cHau9P4hqn5rJEDchDjCXX2bZno7uZi0K+Oo5xDA0
hfdfecOZD2XBDLJZQtX75H24IrpT5ip28Z53RuZRc3x0GArSVQt2P6npSc5Sae4S
Jp1q+qhLn6N4yhWmYZQ/Do8TsdxYYNH5eGo0ICoxldsIMGtLuxJXSPfweolweyDd
u9DKqa0THiiE6ea9iccajY0NmK2bWiY1K5wv1unf6gPhb78Gpzk/v+qoM1xrKcuQ
A3c6Pnd2Xqdv1u6TlF0NjZ4lWk8i5Iv/EOCArEVYZq92mkaxk/iWOarmANQNGD+n
AVkeeMp4YX6sJEVn7CyHvNObdqbGPS6A2WxN7vISNEHBW723WnyBlJZA7bDRnz/p
HG81USMLTgjbABS5qRtHabPxDaGzDzOeIn3VmI3EbL2su9rjZfgACnIrpOnqrb5t
otDR6FZrFElyzVx7ZgoDfGb7x21H2PDZKE3IF+QeblaojghGCPy5ADzuDB5oZ0oi
3NPkg+Mh9/fppbuJIs7Sq29SzOauTjPPDopnN2ym/mNJtk5frQ5+2A0C0wtEKyYf
P/VVLDrUsCExp/cN5ikEShRW7TCPI7TPO7C/6N1PoS8MyNLzIPfZpQkXS67NaNPL
VMZc6X7RqisyPkwUvJwkdydOXIhn0QPVzH9dLK2UjBr+yMqWgrl+fMU6eA/AYPE9
F8BD3UKfhySUY1YCnya992hh2XoNp92WeAhX3TNQPEaCHCv7zitFKFH55ZBsFGrO
zj1nTVki/ecyK+VulzQPTrRiAXvj/RZ5eKM7TEyLsXFeuFQ1sOtOzNd1ZJ24Weee
SqPLeAqiGyV+jY3NUN5SHTrTmkQzEFCX10samWQLR5odPbMq9VFWRoCs+6GGhY6J
XIokaAGJr521I4gt7HdKU3vK50NmvdFewIC2t6CwM7fUJ3tH8qwkrU2NQ+lvCUxH
9wbVwYHrkqGrziZrY8wyQW1ONqwAQzSZSEfQ1Jo53z7+ihtaToBatTmNSk9+a+Jo
McSNtLslav78j9m+F5Ba0yOTy5jTJRPt6JfS2HEqS0SuUGJmObJRV2Q3pN1e46tn
W+lG3681PcC0p99VpdZyYlQa6ygvw+JVf7VreFDMYOPuXutjDSqhEAoJ0AMhI7zJ
qqGOjo3hoO72zW7Hgrp2bhIhgGTlD4I+zivenIBK7aD/LcamTukiigQYJSnzeyyt
+H1F9q5UvHJ01GW3cu9zPev6tBrZ+ZqC6N7dOjaK5LI1r+wsA4UeaBx7/MU/bVqj
cue2okRu66vKZnB4jQ9a+FUPQODUx+Zboieuiy/WrJ98s3soiv0Le7U24aUa9Hlo
97Uo8K4f5rpZqYMHketsaVIWjK2uVDJZrYO3dtG4rc7lNISAGWzpwch6e7hwZgLN
QBtG9Ma/OY9ZCc1p9CwZAIqe5AfeLjh8ltnsI64LNfAD0DNky3PjPsyK3Pm2t/VB
UAflgcluFlx1IGnPlGeDzoorvCKc4UQNbb4NUECv7ytrtGQAoXNEsxPBDG/1mCqt
3R3CO1CxVpbiKe49dU8fD9CeX4cq+n51+QS5I+pfGZsaN/3GVNMCr/t0XIHoHwuD
/YW9Lab8bVdBazIJWfxK2d+qzn/q2Uhk/isbyvkBzjoEiqU11wld1hhVkoqvMEMZ
Ch80IcaKrG1eB41pE+j8dhyGyHhk46+e085iWkxBJHcrYBwtPZgil7ZhS/qBgFJ1
e6F8oZM9TJNnz4nO8V66tBdo7yzfC4OUIniN0Mhdd3+TNVsoYXoTVzEZIMOngy3R
87qUZKPCA/G3KnLx6atFp6PeiPV7BG5q4JuM1SoN+tS9MIRC7LXnH4+nFnSDxIhe
q0yBx+gQZgck7gRMaVo4uWy6Cp+h+hIfsyWuVVI6kVv3NZANjDX4ijItKnoOipCE
iLTAsWgPAAtsJqyL64dicEIYzYdyZC2cuWKQrUME8mXqbR1VxQ1Jr6qcvXpR9bBO
gdJPVPyXxqzSoeHFEjP2tdPe9P4xemnLd+HdZzacN9PDyG20eUDdazOwEyKYWMhb
J/cKWRU6HJkBa8GFVEOL/zXt0jzfkQ066RBvjP0Htxv1ff+4vHNOnGlgd0JxCXDD
KvoOA0qRuwA4xOCGTE4TwTCcUQmggCN8w4bQKep1AT45BqWZRayfJQepyGuXuzhG
b4YNQe1ZUqtSitcxyNt2YLrqKU27aMY0Kw/4Y2FNA5z4QoAXKNBPcRLp5KeMnkNr
z/o7Rn9SDXynciRpowKqaM4lO7hAwi3476hbZjVJPOw8mNOUw4HDJ/rIQuY4Akae
zfHlu5vfC8sMRkn2yVQV3sN0qkE357FhuRZLEq9VF5S+er3Gj2EVHJUiNRGHUOdT
/jWEZxnUL7R2LblUUyUxmZUFZaEZKYRoRn4s7WsbPa9ppIkdhDMwSCjFTyhOZc2a
ijQ6bNmEZCSB4gTHqiZs6duRVuaJythjjIldTb5wkpvIHlJSuwdovZZDdkaMKU6o
p5we+WlIf11XfbYrgTd2K64LEHZKBfMmW0Tx7uHN2hQAVyb/wdHvueiEOPtfRmB0
njqlD0KosOrI21t6cKcnces/hjeo7rwV0d6mtJX77+qV6fLC7xU0SQjxZxWrEE64
zCO9/TYg9Wb/vVZPBMoPbjJdLRlCIcDAOhfFarXFVom1ua6RsNW2q4445VwAzNpe
C0wLoo8yW9gFskgp+hgYn9Cvars3uvwBMVo++eXiEemIezaAh3rzN2YXk0VoXiKL
qARiO94Ra8Qvj3ujyD5P5MiPAw/hxiAvSI1kdxL7HWt24KInNKcwgPSGBQiFQKiC
6Acpremtzfg5RYpWKidyZJ92SEKYftvzJ+PWSU3JBvdDV+2XsBGxPvq9cG4YJUjB
qoUltgS2FRmXuZ7fkZc+AaB7rn7WgpeQMfwVtSBHgqI30cl33G/CsDp9HhymC3my
uSWSxmmqzEkaZ/YS9DCE5ajdruKtHSJtSc+KTzHcJt+7PmH35wYe8ssmuw1g7Pp1
calIvSD3SLlSyJA3JC0/vfReUdR8T2ypog9Ymys/Huq4IDzQ0aT4U+YmYO9drfUB
X0+VC1isfHqVTc6isf8pHiO+ltgjW3SK/QoxxApTyfA96UXC8VBJuMO+DalzCPdM
ziQgzJzaxcC5mVqfO8o3l4ifOim1XuPhcYuW3jZdkAwzd5ih/rZkOP3MJWPcpqCu
1frRUtqBuXYpyDsHBL6BCtCepMlqj8TP8xx485EaZPlzpvSJSW4SbQUPlkvKYlfi
t5X0jsaEWc4wCVQL11/uac4ZFQkBowtL2/+xBV8ql2RCJ800hhQX6eIvQ4BX7u7S
I497QmH5r+qhieCX5EKLd0+Yv1ZDHSaOnz6jWw+YSg4wymgydk9gS0b49gDln2KB
OSssOxKx14Sr8sB4qIs22iif7HtST729DNKDSjOk5TMN2FkfszhLgjg8FoI613Nf
z9qaW98tX9m+iNNvVZg/ilwUruSl0p/1VR0etTHkytax2u8fBCQNyPgqsFJz71gt
1xEz1U5TKJzdtSxvkrGnYN4l9c3kA1OgtIZ1cSkooaUHDctp4NJG/rqSgvqGzYF/
8SXQ4rUz0snUE3M0cZaFGWQOlST5fS4Scc1qv6trWQdVDtnFH6nUC5n/NfVWiZew
aoItpGC/U/uTF9Q55wq8deYM4rfzAg2d/Sl76QycQkUJNEI4QJNE+o7fXCRtAIDa
fTOLuRbwG3q4rVA/Sk/A4eh6coxKGm+jNoaCz4KlEyn0x/2tUVmgKoc+G19lAgcT
LhpIQ7RtdekarcjJ+FCPOl7QW4WfhGwH9lWIgcjHfBidqXbpnhFmlKz7Bu48mWm3
LF8e/sxeaCwHyqj0oSPxU20huo/D7Pt2dGJ8hBZpGW9j2dtvovQCAKvBwfmzVbBY
1PQG0JW25pfnKlU+WYxicu8njIk/Ev03+ZEMI2PXKDRYLjbWcsi/04jOJ3z/rcQm
tRV3HcVfTE5nEFv86zwUljSUxX6QHEVf3a7ayNnG4mJxH9Io66PrC5QQD2AcNUbg
RhT6TQUO3Ni9BOyLHdSqQnlOaU8I6IqY2L26c3qOiLsSSF34K9TU32dR1K84gzuP
AY6qJ2BmmhQGx00HuPAvtZ2LjGtf2COSfgKwfJZl8ZC80qsZNF2pIILDHN7FeTzx
nfuRBjlN2gnLCGsFFvf7l0jfdO5Oq10XU1IiMM17Gg0bFvN2bMkxlsEO7/jBXECF
NSVsmgPW903Bhot6UI9xBmVX40B2pyVXr0aMhw1NS2Qgx0BmwZKiw88m3ur8fj3U
AfjU4CaGyQGYiV+eN56uLD0eiNBZNCfmxStUSwTeQViRruPvaxemR6IcTxayzueO
GkmG75yIWpPqvnM2PCKzIOTTLW9ohFg49rVSIWAwJfDUktH/9zLnLikxyEbXe79Q
A20g8OjNNN2wcLP90/R3XCsfzFySRZobx0YOjNDcSEsY0QGbZSmtiNUITZXpMik7
EFODJGESe4rSnrVb3Nmigw1lUwHS7cTd50M0AmOMljgyxA9Tmqt4vSWgvXSQOAHT
KnAC8sIwztlHf7+Or475jqKejy0dfIX5CYFemdh3uG3wh0EhNQu5Zh1/H6ub/fyT
R8j0U3zrjawXqw/HuzJDqECgw7/r4Mrnx7ozg/HotaD0m0pSoCQAVjes1zXUnfj2
WRiED8CA3237XudAtIm2AETUalPHrLy3iY7nZKGuihhmINEB6tx81zx7aFki2uXr
m9QLX2ecctgCtpz203sjQvlxRDSQUC9+7TefSFGpyNnEZUh2B6YyLbPDHlMkwJAH
Ml2UromfscEMPG6A+iY6Nj5VXfewo6rv3oA22tkFWYyJZHEHyn0BV2B4yY/7uFmc
oaMgI18ytzXd8S3X47fjy2OPxt8Req9UiWaHSsxT2Qsnglr4BbXhJQEX+KWLtRrT
AoB5e0pJfqykeZAIScg1F9Hg3oZMs7I03h3VSpchcZSoCenO+KQfIRz4RdXq0F+q
VzwegZz0j5FKr5tdqlZxN9inTQCkDb9Q1d9f9Yn6fF2FyByEJwsJM/SpYTUUni97
DyKOY01TI6L8UkHXAtguXtExVnH+RHarf0ZXQEhFKpMnG7me6tVpib6v3rfEW2Y5
ymVpHvltuGMT2svLJ5VGN7YCKY1BNIwI3RlxcBqiKdtJL+Z1VInDWoVeJvbSLIJ+
NKRoCEb1kogvR8wkfDlNEzn1Q5bn2HcIQs51MR6W9IHvo+DD727TwiUqYAXTxzGJ
0OEb6KfMP6gRQr9UuKVN2h+bYZ7brXGT4n6NV7RaVACkshqFYVMR7py9jRJb/hU0
fSk223N6ZEwLbV1bfVYMxpXZrJAEW1zBrqsK563lt5ajGDunwQbPuRUZpXBJlo60
1oPiDm8XQEI3NErU7spBJ3R26/A24D/qJdK0km7NqKFQi5Vl07c5sl8D6nr7NfKX
4KkfcnAfthcjkT1ikoWiKiPUFzveNXpxM2Dnbkyn1iv7/W6/YSYUJOevFLRzyHt4
gBDSiZcqv82DoRjI/Rl2IszBme1Pt8QA5gX2sb2mHplgzjfrh6L4XHB4VolaXCUH
/A4h1PkDhZL0Ofdc9Ksvbx1xGezKjmun76iTB0gHVOOxjPjVzZYBAa0tc8Hf1VPD
mBx18zYSqNxjHvz9BgnRQSmT2nzQyvFclOvt74opWzfjSb/bNS9u+pJPqlh4yh9S
l9efacGsQDj8a9rubXEBT8CmEx0H8Qnys8LfP46CNDsYiFMiLnD23mqTrUNsz8y4

//pragma protect end_data_block
//pragma protect digest_block
SW5PJXif5he1Nzvb5+2pSvsthPM=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KjU+/Z6J2rN36kLPDBG7iCecfczXawgMdeH2r+7NoLC7TcfKI0cr5FMxZ+B8bObQ
dkh3I8islBEuKk8PezCfJZ+LLdvDfoG9AOnmEwhhPDgVSOEtC+4l732zJ6BP8kW1
HBNEbOVas69ul26/X2ts8AgzO0ZcC7/gNVCIJGOKvkIWB4OmcN20ng==
//pragma protect end_key_block
//pragma protect digest_block
BWNLfHgQrOJnQ/fZuGyj11M24N8=
//pragma protect end_digest_block
//pragma protect data_block
vWJ+2J1WCPQdQuifbqd22WInP/ZamS9YZvNjAnZmc+Er9KhhOX0LY8/ZdRtRm/Ez
Y9m/44ReFo1XW5jaKH8gztalo6mW6k5W+B3kROicE5uxrLqRL3Hy8+LxFshsPBSQ
xgBsSyB8KTGE7semHFsSBWZcxSHtUn6RV8hnLypQT0qOn/r2r9wws+Svggt+8TLB
2rhG7hI/+qbfIi/74jjrqUwEdiCgJZzqKShDB+cNu3C5BjmmFhLvV5RHacfbuDUf
xH5GFlHxc/gKzXcaTuoirWzb1LfTTIKy9D4L7i6Q5jwZX4ptVGIw9pXaso/RIhsy
lxwpz78iy11BvQtSZ+or+IrVMAKOifhaSjgl55V4IiUMBLZZ/z8SHFp45196fQ83

//pragma protect end_data_block
//pragma protect digest_block
RVmbGs7ICP9p5/2ZgWJwzff51tc=
//pragma protect end_digest_block
//pragma protect end_protected
      //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
I8y4RwCjan41mTEc11lu2/sTHT3cp2QbQXX9/iavdOhNkf3gly0Kv/tkocoHUbQa
hlEZ3zj8Jg8AhL9hv+TEBc/lAh4lkbTmt/1s7Pf1fX0c9MAOzPDWWWBs4itF7FUt
bE3SfF28WUXbhsdOrFdt1iebEvSzG8TRsq9yxls7MATA8HOVJCTAOQ==
//pragma protect end_key_block
//pragma protect digest_block
rFhkEj6VMMFZN3Yu4tdqmQKMJS0=
//pragma protect end_digest_block
//pragma protect data_block
cGZqDZnTgHImK24K5r89ECHhV9o7GU8XHKtoDH0xCGYd2OAzKeemD6AzQcO6/xaV
g2eL8CoGu2EpB+DU6c6pBVl5f5l2XZCiCjTWagzLwQt2WAY9AXtACOwwao6bb+sZ
Nk4crQU9SlJ1W31esSTNTxDpCks+fd+zbpjUcwqAWSHj6xICxxFPuegk1RM6O+6m
uRP8SuNj6daxqhOxuGldPcnPJN/hy06c14OdagNUYf/jxGHYyqhej5Quz8hdu9vp
bYlNekhC5eMDAor0T3NY9vti2Y9BcJursnAfdh9V7raNJT7387PV2IN5VioOTNsu
hVQL0I+GTB/QgDs9L3gfLwHnwhFsGAAyIYjQa4tjavQU19hrh/BC0k/IP9FdjknS
mCzigBupn/FG9xGxv6TsesKio37/d5jAvjM1g3OjJHzUEPioard0D5szgpnQ3szo
andVdx20sBKd18nam3D84u5myrYycaSfoCpbny3qFsE5ANz08w8Ex/JXM5ydjKX4
k70i4whtIslB8veb0ed3znOQkicfmRn0kqH+UDCd2FCBTL7BXjReoyItrO1keRth
S5HzVlZ7+pjORz5XwtqOsB+2DLdaLwEDYXOtLbindzjxBlzRZsCkom5idWCbPTcj
t5ZFU9dauPZmnfFd2BflygKPoc5TKBMuljio7YU/jxneskU2zU9v6BA8HnmdvOA3
4svT7w+BYr6ycFyblJOR5HX1suyX/K8Y77J2a+9GOP4NBEDKdNuvUiaEjEFDrJ1A
48l1dKoThJYF/ykDhbiBBjkAYpmPUxnEDqAZ4XWGqxbcxReMOxxymSeM2HtV4Sza
xVuX1BNaqM2GwL9VxE9ip8hWdHaf8UZ9sVMGW2l1rXzTmeQy45vSInnbbMm7rUO9
oFEtbk6Ggm3nWkGOCrY/UmT5yjPEiDISX2HDhKFhblzI7OAj/ViAk+UMqV7ADduK
cInYYFjFJctic+90CboMuT16qrBNLt+wsJaYNnB63r5DAd+jwbN35vxR5hZZYkME
P6C8BHM6YA0ZvgKRuTOf61ImNzy5gDrNmtu4aTD193SLFBVuus7uITPUVy7YoCN6
9noYNZOQhglfqT2j8zmu29Pz5ufILOHreEBFITBQnVoNuY9C42oq5gj2K/7NKD9n
Upr7vWZ3/Hll/ox8ypkZPM5j1z/gjB4NSFtkCzS8YUPpj/id4yKFnY9M8OAgGOUi
VZ4SdhbxgnjIepyVcL8KfuBABqv+8SL67p2vwTVvkkj1HJ4/xqcdX5UPWXv49ay/
CrcAmTFjqxh94GKM8RPz0KSOMWjSNsUL/R0xETrgoONwJ9nlM1+n5HAtju7YR4Ud
snvQhRlEL/7ZQ4vdqvKjW3sjH+ZgZIik/SssJVLyGTJrsw7mv82OJs4YkBDaUSZZ
K9WOw2rYQi/UBDv2j9RMgAOdlIxDXKw9eGV857tcB27bp3wUl7WPdlneWX77UOgq
soGSUzlgpGGmQDri3H81ik1Y+3ZVCcgJ1+cbMMq1GVPGUXYSI6elAbbEmWo+Umjo
sz1XFP5T14/g7/A5WRmRQt8piqJh1ezu+wtqtVYY92FE2+Pl906ab3+jWW++seuA
7zg3o+aNOuYGoTL4WwFvOgp5UAo9xdojDGL4vlxnxHD2+oxnng6D0XzfldehHXvW
oXIzxsvVNiD0bL94QVVw6U4L1omtqSMct3fQsKj0lYNck8OD5PXD0M7cu7to3ygv
OfLXX/1ji3qtt0UZHkNXCdyTi3e7tNQIh3wwOpiDsHmc3WzHJrlmud2GTuI4aRQN
JzKSKUWrR5KJFbFioS1LWi6iJG/GN1HWBOVMsTG6XoF+cS0o9Y7wF0vOLyGsAkAi
v2dEEw6TgDL12rTftzk0OEHM4FANjWQQBQidkb+AFgznoIIQRL/QxYg1mTJB9htF
ipi6np3ezKMxi0T/VDKpvdstysRJg5S7ZAQuFJyvaZC/9DNNRSC7dd+2nS4mG/yP
ezCaaVAGA1imEWNFcp+V+9xCYSX0v85Vya8FrjLmYXlF0ddG9l8/UsJDBQLrah3t
ZvxLQbSo+Kyn133G5s0HjY9ETulEgrVnRoAFfiCsjGXwqUUhlIT24iq409TH+rJ8
bbY+md+wGcKlCFg34PDOwwZuIkh9QLXFCMAgENDglE5whaDvuZOKW8a4tJEbBOGO
9uGQxOI46V7jgunmhMx0ARY6Ih6N00d+cUT4jjMuKoEKaA/ST1jjvgolgQKAyLoT
14WhfGcXIpRbolMzMmmkGVEC9Nnf1ogIGa7h3jqSnQx4tSW9AcSXiaedJs2iOC5Q
9EfdbTRcHAH+WdNAaGlRNsj0EtbVz7kDOom3BqYMVdDFzT/UilXZASwo4CzivWDV
Lo1GhQtIXRrGkbzLVT0vq4R1NrIXzQcf3EC9CAp1AgJpDn7+icemO7RyhXrkoXuM

//pragma protect end_data_block
//pragma protect digest_block
ckkat2UJHJGeFSu5qn8JFV5yLDs=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yUn6OrXj9n5ShFXfd2T53cnbWSOBmBi76EqxgoGQg2EleAbetCeS2hQnkgALXhU0
1HkTpNUUBQOgML/TtHgbOOZgDuBAR+vyqbyy8lP5OkIKdmLEOe/LNA+J6e1dPeed
4Y++zoG2sMUwNQ6ylPI5CwupHK57/ayu+rknlB3KQjNDDybxwQH5jg==
//pragma protect end_key_block
//pragma protect digest_block
Qx9q+BTKzSf5UsPEETMZQHuYeX4=
//pragma protect end_digest_block
//pragma protect data_block
JNaNtedDcQqDJGErzqgO8oQT4UYcSwpEMvEn/1lxqoybMqosc1H/ZJyovLXoko87
JT8OTEpO2txPjKLxl0nOP5xxDUwZGI7HXUaP4W5bY8WDN4PNTTWSGNtRY0DqkHYu
xj21YIcK6CHZwcM8qXgxcBYqYLtYea6iy+3Q4WZXyG2nCc6+VaI2ukMHsof84Srp
2IGdI3eDWIzG6qv5ESZn98scKYmmT9/PNbZDwm0fgX5qRZt/FAHTdWYUtqW4c+Lj
T9URs8cRrj1wOpK2nfHs4M0hSBWzXsdb//fqbfFsARFUO9MBRfR2qafGBP/YQxtu
u9gcX/BEqOPvH2P7Xxz2EBXfTW+GopnoVMR2X0G9MuopyWryU4txkHU7m7hqVq8T

//pragma protect end_data_block
//pragma protect digest_block
QOANfQ6WLTZlklkCWJez1Sn1y+E=
//pragma protect end_digest_block
//pragma protect end_protected
      //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
u7t2vqIkKUAMeVxkdY2D9Q0XfIuxwOSAH8KL4UxRBsR5g1kHRcy0HrUhDLZl5ABH
Z09NTE9HPNiXg9/mhD+EJ5UytXBjQce6OLvfUk6Jw54vhrh+Nf6Bj5iEFnI5rIHR
jK1c6NS/n3iDfCfx51Jsb4orxPr4QgBU9h+haSnwJ6mJGGoDFJBWFg==
//pragma protect end_key_block
//pragma protect digest_block
Dt1O5WrwknfCUo1JB8Y8B5tj3XE=
//pragma protect end_digest_block
//pragma protect data_block
XUuaL8cTVs/iokumUCBX4R9LG+TEIHbAxExF5sT7Tlyr6ZZivwYQwAjfXioZDbUD
jWRB0rjqfIYyolVQl97uLhBV9IdCQOH65Hyu5nB3t3J83FVwWZyZ0FCnWZg8iIr2
UtzsIwT6xblSHmTlzWp/ZSUT7DGQjnEMzcy+/KpV3FAFMUr7tGKPlnzL9t3ElJ2i
UlMliVFLpG0g10C4LadcEhx865moB/y22mtlDHJPUXgtYMgqrSfQUtCRhgqpuQAU
8MZ4FYaQT8GFheY2gmWLOiaDSEy7qo9Zw6+hi39rK0mTnBhEVPbpuwGI32IcGnDG
Mpuuo2S9IwWYYCI12obFQvHtYe+edr+AnY2T2GyRhq5PbX5FQ2cKqbGAbVCO9oKC
pgSPdtSxtsTn28hawc1yangdXmc7X4WWIR85B9UNXttwazVPUdS3nG3ImE07eV1K
jJv+Sqy6JsSpvswZlCKB/F8wROI01sPgwx0iBaQJ53+Wnnt17XaOVfPlsN+CyEEt
7iLcp1qWe/u9WsN0chluzh5XNCOQmwEvbRETwHq1buEtwfryuGM/jN1zfEDgyYki
xqrM48bwqSFQqTG1vU5FTUaZehUuJCUuOaRDL8k8/PPOf9M/NJFGUr6fkC/LtXTh
HRPTkEXFEEWx4z/CjMmfx4ee8eiqpmNG8V3pNSJdjIhu3y2R+8LC+4XjY2lESziz
OqUYJKzhdin2W7zXBU6YoVJWLqvET9A/SMJMquPH+qt9ilDqEzccZMR/duTIqNl2
RKqm6RDjV//Wuj9tupI+HyKWY1fk4mnwgoDrrGjZn89aC+/BF31bx9dtu7Nx90Ga
Pgo3AJfQDknzmcJ2rbEFrvyuZY8Bhv2AUKAb5cgWAk8FFK76KIeBpbweKDqfeiql
/wPiK17z9djxXyXYrxOm252+M0r3oNUxk2qUQlf5qWIdJOYxZ4JeK8BERlU1oupJ
4amt9e7064Lfhl9FipUJqpBcoP6OwbzFrq4F2nDYDsUtm6B0jA7535OWEBdg4Gjj
IqO5IXb66WjOyG7/UNl8yDDC94ktSfJdwOfvzuRnv7ON6HpuptIf17NGiHbAUvcR
tU8QMhncdFwD6KiFJF9dkdm7n9cBHoh6Qc77+2G8kMWZBv3Ywr+Ouf/GCuntBnjZ
hIgZpEcx9PVgqucA+n5yIuLNDdg7Gx3laGeUyapro5sjYKOsM/sdVIwgZcFf3VII
quBCnSv1O2uhP1uNlCzcpnsLHcSZJlbEV4bvaDUN9VP8bDEHGoAhOsdjUb0WMb2K
yc+6qJU9iIqjPULalZH3OR29WbqD496PvMuAiid2VbpntwNyRYOU8Xagz8TQcEzo
gUhLESNu2R1g/GLOZEmTWKYgI8AHtDacIejRSX/neu7saGXYXipm67+GEtZfLfWr
S5aoVnXg3kbIn4ig5E26rz5YWoE4QgdI6E0fNvMekvDmiMYsdTktwQlqI8GUjnks
b8LPZSQAoOQy2CDW+ZQad3Wjk7C3t9nk1BkGIJWDqGlybEL5nswcCzfMT96JBpWg
WpUvXLfGNLL29snxjK2rj5wMlmrj0jZiBW2tjPV602nS/MLVnfEmat5s79wv99LM
2oR0TFFCjTx476B/9Eh2YNk9Df9IVUH4s/IZnD0EzIVBrx38AMsZ21qQsvNmdeLP
0OucOB0Nkfho46iH8slI5U7bJaWR7aiONAGgsUmbT6Ql89zW9wjzsCfFjmvl2deg
Kfc06dRGyTJPYlPa2+OqQsHrnBSA1pGguZbCpph+pm7mWyQPK6ezOoKqpzA0jBWH
uonuBWp4h7HHbt2r5wHqWiAM0iO6Hmap5j86OFO3/7uO6ANnbtJCip7Yk8BIoEXg
jZeVZiz+xsVaDad4qRbfZLfvYjNzpq2LCOOAXnioup232+bp25BYhYj+s65KLadV
em1HFpt6a+5NkpXdGOVZf1PzGqcbwZQaRrN4/mHdFOazDh2nZJg7XpsKFndtsxjx
0UqfPrngtV5F1DPnlJUqKBD10FYjqfLOQNvJ4LrScPTdtudNRKPlgutIaV2PFpRi
ZxWV5IPRMZcKwJjnp2Mq9nioG3lPHl5A/Q4/6CGsOPh25yG21aDwhKE0xV5TX2I9
AACLREj6xkx0nuSffh7Bd7DWpoosMC88h46u02rQRUzNfQdicgmqI8IlPsBO3d9F
l5RiQcBgCFufg3hb9syZaOq4vc+P0QZnkxU6aHjc9BB1awmBhlydGsA0I3wogmHJ
yTUN/5go2YL0roxp0i0Lzl+2fKDPoigLMoScZgETEp3fGE2sgrZQRiQG0eYtJD1w
fmFqcO33Z7fsowUWTWjYcj35cbM2v5qp+duLhAtQUlqFyMTbzs0+lCzc7Etua0bQ
RUCr8KnTW3WHu3XeRXD2VMTAxAsB2QX45kuzMW8YMKuKCub9e/tF0Hu7IKG7CLKj
8jgkQf1N/Tjyyr6MpLoXF11kzjssvGYDfni7u5VIJunZ9tvwAByNT8BsEsrWohw9
G5f90w4VfqUsRLQR4y/h4nKRWJYWQGVArXovSav0KJob5fHNthQQuY0fOKC6G9r6
WeS0dHJ2hNE0G1SWqvG8U/1TCMNJNCaJ2LFawrUp1AO/rOEUN2eCLMCpExVH1D1U
q5JKHxk2HbO5xiHIVNGXZ6rEogKAgXNXd9LJAnrlwuYfvFWrulNWfkRIqfKjMicX
WhxVvnyhhaQYDxAZfoMVtX+wX1IS6zCN9geJaHQph2+Hzv1aNVyOgTPHSOEAAZct
IuWtQUAxWmVgqDVmXZcEqABoIDJOV+w+oqo865AVmSmcIY2vmEjbuc5ZBpSeJF8T
JMoM1lUVCFcYslpvbyR40ipiQ7Rqo1anzy/fdemLi9mCARaYqJUi2lQKcIRPJ0ly
CCkxxFFS3sTiu7L1T67qsWvbSgSZQZWqRJ9TetJqeJYe+/D5YWFH16Y0EQa/LCXQ
vhk4Z0hHXQi0s0djizX2pngFTYk5Qo60fAkOGHl3cPg/7GBYvVl8uisadgEHu2GE
5/gPDxFwKLW4yYOdX2ZRmIEwBGxZdAlB3sEgWzLT5C5Q/4fRKJ+1z2SrRzJG3+Gp
BMWw3A5Q+vynp5bW7JxQvaOXQNrrWeTDFdWRz0alCsKMDOVPzzwsaA1GBud4Ync2
QPrDCjEndu3I5Acd5MXq/rURV0xCiaQVmlLVEySqo1vgo2wh5C/IMJUtWqpIQZVV
+fFp9+UId2hDsZzZnVBPjbpFln9hoC5ED562ZbhuBHMYxn9K0zUHU7Rcg5qcgwET
LUbSl78Pa7HMsgBRRar1YdH8+zI3mheY3f4CECLDlv75W2+FHd78h7zJj7o3zUNH
RohfmikBQZIDTibG8i9BQ0idEtoVwC2FAk7mK1qH9678K1JWi55RFlHTgCh8UOlJ
lH3IW4OoXOxhPIImP13ru6NllOKF2aUGB9xGG1fYHnFKAfh6yc7nSgv4luzLo9hM
x/qBntxdXqxOElEDFbE9P5V/lqCmCTAvJbENWpgIKH/qy9GJVHwfwoqT+s3RJBC6
EDrFXp7uGmvw/Z2+BjEICyMjLtRLRQOtLROjxF3MrJEu2OhQtVc3/NFfEM5MYzt+
yQOGcjulKste9c9Fbwe5plyvrushAW61v0Lz490DjeZ1Fm1MvDW9mMVl6sOOtMBA
HfimnX2m1XbjnDuPLY5eW23m4Ot/qW/nT4208gLwjQAhCAN6zTy27t1Y9iD3S4A8
cX+PqE1b7sacbpkCUXzvbf+q1nascyHiafsJHvtNW40+xV1jPQvLIuhrWW/2xf/u
Etg5gpU7qOdCA30gJTukKtHDOnx2tZY5FeOQ2j+o+QeSIv6XpX0Gz/s/AYxAb+Xb
Wf+RfINahAr22+l5rXoSQCsY1oS9Ixw5ziYO/jsVFSyIU3pcYTBaSmJtRCgieL7E
wsjYNxuf7ClZuSNMbHxWUdQEauQEsMYDvRTbTUgWP0bZnOXjHW2baMHzXhzhnWdG
/W4/CcLk3F6Y3mzAB3murxDQlQW5kbKRWVQREwD6xZWbnboqA+suxYEz7ztgEnlO
n2jDtz/sGTWPTbDQnrzeQdi9NIZb6nI5dWSjDsaiiUpaELgqZ3/uzxD3qwqP7DFz
LKlv1tToQPud/xq/G0tKZYeVuvK6jj7PCN+pAOV+yJ8ro6C74xMUfZ9aHs9ydKIX
cpgjy6HshuF+sA1BX4potwBunWC+S2FOn+78WMlMjLCO6WS8luzLnHVh56AD0O1P
97BnrAwM2OwZk1XY/sj8XGkOk5aYwHhwfLWsNemed5cws6N+tjF4LYw6UFNBqelu
5WNmSX8rKw7Iykggc2xMKGY1UPxBNefImgCaa+YYNnyPi5K6Fb61vSNXtjj1oApK
qK+sbIOeO5724sSZqPjBVv7QQxwAexL04PPnyeuqi2SKhpQuAuv4WRvnyvwxrCxr
yIa/JwLhdTjWIh7er2ctB9SX2TB7wwGAo6xFy4PNObadbNdcc3Hh3sfTCS2+i0fc
j6tV8B21/l35lEqRB4nyyMiaks8Ov4gsBaV4gPr6hRkauTYD0HC+G3ChOLa16KPy
9ukKvALule7qBLr5OLdEG4s+xxQpG1uttY69e5G8XyuSKPAxyiPQb+yP4ezHieUD
+Hj7CkCJtfSATFP6j6fKGqOdIPUVouKo6zSSD9BtJX2bl0BPZt4bJdmew0qZr4Ks
hd4+AN10c0gKY6ZNNu1a2RWlMP0nnQUHC9/v4TvAEo1QJN2yJdF9rk3mg20UxdO1
yn+++r9bgEyyj35zlmzhkvAX1oKMh7h9X5dkfFvzUD22fOUfzneoeYIIbzGzHye9
pW9O0VEHFFyLiNDmDdVAPrArjGqNbuS2pks1yn0qYUatN5w5qZNSVfh/HJy7xvpf
UiO7XsaNrP00wcFe1yv6Vrbw44Y9Bi0N8z/FmLNO8zEQ3jaquCfXVRQWioOO9o0S
bzcTDZtRH0pPM3qk78Cf0cSt8GoZNc6E7PvWT402rd2cC5hVlY4LXo/iwRegbVQf
IJsTSQW5+xwG+BOG/fhPJ0DmNzpmMLNMZcVXdBUoogcevs+JL2yplR1A2RWbDlen
3S9Pn1akIkpOjo/f9ZXT6l064Bbkp+Xf/T+H/EDlu+9L888uKVQyuvajBVZrJneG
8gliEj8le6VcN2Prxc0Xb77N2ryf1HsXXBh8ZYdjgDnsF4no0VVsuW0hFY9aVqDL
z2wVoJ3jVy0Lc1FuW67GLN54ag4u8W7lHqQ62bDcTSVa5bCC6681NMWOk2oHoWWh
6bytr+N6i0TaX15WzkKdECT4xZPGE6B0vcMACmgtRdrOWzj68P4DiTnNB65b2eba
qgFSPCbaTJqIs3MMnhJJXUrsd5b8B5UZm96AkPF6mU3mnh3nkkvLsP+ZW+mZRGKu
HnL70X86vkkiF1173Lt4FhGWWmbHJi0M7ZAKwi2a/KMsxargPK0gjIrtdxzvprQs
uv6Wtdu1GLVcPSwCfnI5/dVePSCSGX8FAP4URt1JHApEkmKHjNbMUFJgGHDmjaE9
92YqGRQSpO+qVx0Mj86Et6Nmo0VaCeD6PwM1dq8PJaFQSvFFU4g9Wj+J+NXMeTHp
ucjv8VWNOYtuSh9GJGbTIjTaKmUQNqgFQq9NzTBwXCwW7Tukt0Uv9fJHibtqyOK7
35qXiFbyhFAZofSaY1oIkd0G4eZw5sgQ8m379KyzJZX4PoeQC6N8ibmiT16Lz17V
NlI97fHymqqGTXnAUO0wQXYWzUhk0aVHnh77i75ylQ/a1GYJWDSiY3qW6RUIHF4j
8p73XYeZlkjrSFnrr54qF+9cv/6eGcuosS+zjY6wyy4c8VsmVTX6gw65gXWW2rLO
BWhIuGI0BKvXWSaNgcMbhnxTlIG6kvT17HqXZGtE9VVHljjQE+9eRb3GA4yE4DMi
WgcVBiwJE87sVAUJSaFnTTkURkCjBFtccql8z/XBIFeW7q/Ict4LMZAJrrZgKkxz
Yrkh6MHiDjOFKBvtib25VSULDdDhdjc9+tgw0qtWbigx6dJcjjz45zszMBA8IpcA
EqoCPRDR+V51XhqJiAhlckVDZHicr/e16V58cKD4Cyr8eQDg5i8CWdHcQRivesoo
o4dHLpHIWabkuR1BIFE3CgWY0RLAJvoKZ3Nu6/o5K5w7Me11ybxT1C4GKKwXb+iD
jAAPgsI3hkUAWutC8/whP/alxGjObkl+6G8xfUnKyTcmiJEW4gtdGddaV6xyx7QI
akQsXU+a/lURUeWeOnW3F1yGbwWHBesxoPaSBESz/2HMR/Yod+UGkMsipPOWGFi/
1FTgaHeQplGzUmroAjw9WN5pOcZxdBTShRZjlO/xOHFX6I5FPlvs79mHuDOOQUcK
lFvsFwIUkh46Mu1SpUO7FvZGITvQhV1GsmIPfNj0UotKtSX4zTTib0OoaHVUMxox
ePLeQZw1lDLVCgGdonx3Zg8SqS3SMQfrYolp7ckdIVAERSkj77MYIJbaJS3Zqb5J
Xn16JN7/Uo7nz/fVL9tQ8ZErXFYmFbWohYBVyVAmWHCtZpa3eGo/3djX9wag4kYq
og52jb7yfAY5uFb9PXJvPnkldtnl+ERO9WF1jP2+mPvuoVowwz5ZcZSomS7RLXLw
ZCuF8+0lcp92YEcOT2AG14FWesoih5zgrjD6ziPIpWib81PxSZY94NQfH1mTinzc
2z/Pos/SsglEOfoYKmlhV2RzJLXuRop8Zu7SCG9O8ZuNIs298vy3V2s1QAffbNPu
MTjd2JTxY3W5LHeEHaHsAKkltMMfdj3L3oXI/QmqJZpNkr7cLEC1wFrOtb8MtYDe
7RGLvS6tjBU4aKuqu8hv21I9eynZlfpzQUXAVjGekuqFZ0h9/o6WUH4/N53IpX7u
GO90ax8eVkkTFPRgIZBxAoCaV53fhsw5ZmXktPRPVjyJnkQrN4Z90DnE2Uv926fe
E8pYUZNBD6WJrY633+PP8BBxHkJEhLDVr67jlx6byVC67HdYM0+r2K4t2s8Tfe90
UGc/jyrMa9npd2iM+Hu7mcQ20c8tOwwtJd02W94pbpI97dzg0lIadstYLLHHIJLp
gxKwgxAmuc+nYFqbcxmu+3tKWkVt20Q+U2aTwXWY+CJaGrkPtWsvUudzDFIZaEug
D9r0CiKRB3plt3o7Fbg34Nigup77MXmcqDuMgtUzY3JvVIrlzn+BanxB8MJN8tnK
eV2UDuntRQz/kZaQ+XnBKDDBJP1/dJiof0EZ8zWmB1iO1Us4z8SeBQzZ4pOBgMAS
iKhFMdreY1OoAAxh4PIniH3t0njiNSJC1e2Ath4kRL2bVw/V3U7I82ccBeo1pP89
EXxX65xe1f3HB1CVoMzINKsZg4w+Hm2dcf393FeHPX7emsBgJ9BNKuia8XwCbjqC
iEzQ6lk9Ur5+9FHD7ntZjr3Co2W9ozVkBHmE3JGeMY5E/uOn9VCQPYZVVLIalJoc
BhZ6eEUdWqM0kb3IYQyUXSgUMA66CpDy86sVMQyRLoBxJJvGzRrVKVlsmQ/n8XFJ
IsRF7yNI2tPcI9J9p19kYTf4DBMoffRKnd7r4PAeRINcuHztrQthpCbp8nl7fk70
1Kxow7ELpKxGi7zJUH0AoDfRsmQMjti6JaZHZCpk7kQaLIb3NfIqChPNk/DzMLjt
fsC/qG7ezmzrVLVuaFo6Kfgw3clYhBJvzInSIqcTUfoSHjdd9n5uDgu73rsDCsUc
smHAhsxsP4I66R8xoXayjWjyW1C0Jblgxy8ulbtz5gBvdCpD5AyfW7/OxyojW1dQ
DbO10UQreWhunTYfHp2nr7vI98HRG3y+jD/2DltH9LvXatK2t9aNhZKgrd/Y2Nx2
IiAW7GYh80sRVJSp71e3GBokeI7Tk/P1RZ7RKIzIuJ9oBLiP8pVwzp1BZB3jit8n
lrlupruV1q+qSBRo71nfH4K0k9uKbfyFlwWX2+MKLKkZCafAA/SjF25+LERI6rV2
o2Tfz+eicZPimIMW6vTbErZVbjatv2fuGYP0mMdq4ybkd5kMprAPQXS2QpeMfoaB
2MOraaE9RNXMjyCTP3t0Pe6u8ZuE69mM1tqv6rl0wK8vmFWgSmCbOuISGa5Y+mNf
6pyo6KVn5hXllaBEMscl6Muwy0OoKMixZlK194A459qjkxJ6nFBsZAtRdOX9b3Un
hw6rlFFZ2pCq18os3FcXWys7ugB17Zogrz+ox6oP3ybP79shhVjRAHYMelUPb5Ov
aBjqYmhOR5MqpIORLaIiC0e64CXJH8Kyzxv6XduLQLIq8p0OdKg332evRmvVNpJ+
q3az3JbfsNG1W5u1o+HqhB1c73vfQVCcIFs/MtvCR1sL8bu1PyuqRXKu9rmi+b6Y
28ScrFoXgopzh5K3ZLryC9aDQSaFPBiBoRVTTPnOR+MG36KXBlZdrtHs79ggcuit
48TbG4QKFd5wkXnhXnYBDzFAlqUUwx9p1LhSdKLgrxMQjLzNztzuOD2pVaJw4mzw
z63exJ5m3ZtN6ERPs2S3oeynftiMPLf1XX+octY0dwKa8ZxGrnuh3s3VDUqMt0tR
mmkiOVwt5aDiYnKuBHR3a+nR28OS62mLWB9KXW2qPGyZwoPtnaUo8Lne585iCQVq
R13Nn9tp+MfGWhH7Pnv85jEGngsUa1ASY7Okdiqkr+PMOvF++cbpnEpZoWkTpCCS
RPgf71dNXeH+Ejpod4Zc/3JUK4hBce0Ra461QNC0YoltLJIqXZcut3XtHZrfF2zT
ffPLT/4/EYnBh9+kxsZ7bgekW1/E7Mn+T0im8yf9CyH+euhxORaHfJD0ZOaRKHkV
LCBumLg+lGpRBen7FTV+R4HPIzmgfn10gnPn5J848gXyu8Oh6wyshaf9EjjlaXOi
1F82Dk3Kb1+Pgk8ZLkJKhJCGxIOzTE6SYBnC9R8CA1BIewsGSFs/4EUAXhy738pi
VINWGUL4OmUkH98Fqv3DrjMS4FnK2D6hy3iZsCDHRkGQM556b81ZNE5a7RZ6/vc8
uktb+9uZS4WJT0w98CP582lFGQZxqshBO0lAgdfYg7j8c3LI/bXyQ5INNARkc4nz
H3wfp9FkkscNSfpf2li5iwKEHdQxW/Kjmrwaz0Nt9ESa+rVNkjT8Gw+D1wwVxRuk
s3nSAbFd7wq01AuUNGM0yNZWeqFZtbmI59RpKftReL6yd0TBAiitLhFM1tYUB8fP
B2AzhtUq4J09tp/YN9apkHQYcGEwebMPHb7xyMXhr6L2N/Fo3LVEgxAzHMJexG0i
jrQyUcneL/O6cY6ECY0zewhQY/UHwR2ZwAv7jbAMeGY5VmjqsXxdaN4V51xkZJxo
EqyTuE6qFPI9FmML0EYMzMQD/JTeR5pDVPMBIH2dfhzG8EHCO/mqR8PiCpGmvScY
YCjLpwUGyZU4iGPlLooaxqeL5hkdIq6cCFe4t5pcywLj6N2Sok8k9MtXn0KnjNYs
I48QKIQqAIznGTbV+TLI/9TnBhIrNFB+qhvwp1GTzGD9mx+xjBHz22pfMuj/tuR0
VwiXGCM0tirSzvKLUyDMXAVIMhVoLTJbtl3xSbg7+XwNdHzdnf52G967lDdjvZvx
y4HMBMWjkmSPLMyKkV8bpYWEfaIRHgSdurNLiUxSx5MITGpAy1xNk1hes7ot3LKo
tuQ0UVZ2dsi81xcolr15KUzDUEN89kaWXCuxyo7YhRQGnbM8gdE20z4ekfZRnOqj
GGEhUeOseyqFnFVJHDtkWrbBr7B1RcY9XZSA+cV3X+dKZnh0ErOqy1W9WAxOMnvf
dJQdyer6Wtz+4L+DhXH6FICzANekDHoN4uLb++XzxgoGhBoZgDgmgnAhPYXznmzn
irfIjjQXFkH8DP6sSlHJEiwqsp5j81lGdxWw2iLhHQ5FhRxYoM00+mBYtztLBcbo
MVxBQ4b4wQDXRMiU8w+9QDNVVv2WjXZuKDj9CgrwX0wK5QlLbvq1zhCq/q7m39In
fzXqoT6IXyPNk6OqzHCQ8mwZKAUgymXDmEHncv6To2hcv/h13M1U6CTUskhMbGb0
rLBsxLQmveB54gfTow0yi2ipf04OyDFlTLY48V8xV8uJLGYN1gXwtLOhDNEjZ9V4
zF6ishf0N0E4byGxvv3rGDE5cq1CDgpCmIeZczqwQJXctjDtlT/l55AQ+7Fn2tUC
kzLTmOI40A3ygUvw2Ltgsw9X1tMrLIoFmDXu2ACH0moo3poYNd5nEjQI/qsS2EVx
4Cp/VuoAogbcvpquF2qnM+AMsmAMGTPz4QQelDHpz34o+sa2kLPxntPP2LazIo2V
L3ReJxrvZSBtR8iYPvL7bI00xnT8REPq+JqrWfbnfLsVknTAHaidKgldNof1Lg3/
cEVoX+eXM0GnRsdi3oKDrKuQIvm6yzVg/TBKYmJPy007q2gkRBJCbMtiSVcKmrpL
DeAjcsAsS7dTwFHMjcJ+fZBEKzRJdM09GW23unurgsFdID1ZdmPysh1BH0zBgu40
sbEZpolTc+Jle0879xsq1grJmuI7F2S/fDvqKFDaUa1Lmq/iR8jRYv0Hfka6aBgE
owbSZhSuy9fONPV0imITwwaoDxzVsGXborLDOSyMEy9hp1QhpB0SeBiXz59VM31e
GwBOpBHdAVRPBzPXySgSud4Pi8wrErKry77SZMBGUl4UJCgmjxw5iNh2BlUyiFvu
OhRz/XZoZLpomhWE+7IMyiTLp2zGs50D7B/f4q6xFuJ7cCGrw7IvzUVBOGc/f1V/
1pBk9reNVIFVlMxwSHCYWZBukjUEG8hOyBltshnVe6LwvsVrayGTps/n4CJJK3nJ
3711s9cbylKmeTUGe+TD5ByCmGMPlq9w05txXaW8u9UK9A6Ck7Z2PuakfUkGOJby
2NKJvpSZamXoX4dLNalihMYbewbugSZstMFuBVOuTrhSo9qLWr0+m5EV4QDncwAb
m5BC9S5R6ZlmunkhebcFhKmcv9Mei1WNobwQ3zMHh3UyRXbTVmrRWylV8TmyYhgt
tU/RWjdkVxAWGBXXnKU/mHl7mUBjowD/UqjJRuUJ/lOLehwszznwxReZ29GOLC7X
cZDu8N+CgwIIJzsDj2F5EWt+xIqR6vcrJts3q3NpDoTGKnoSt6NCIS/xhWhH7vdH
tgTSEH+A4aRHaOgoqGv6xjj6TRkT27jGUnIyzYHsq/hZkTd1A7i+dS7CcRwR+2F/
N4sRLGg5aRRIYWV/eW3xLH2TFQw65GXBR8aFBB7RHj6wEBzJn71U9SoayLBiLbMY
iYsZYdsXQ1eq/Pl8bEu2PxbqiDVrYkchiCl26v5C554aLyAgeaS/7gYHRTcZBmQd
V0nhHUZsa8KP0JYAzuKINusyJtaZXcjKzRAAnEqW4TzD6XTQWPeahzI7kHTEma3J
wI3fb1iM215YlMrMoKD9t9RXN6X1ObDUnyi1bVe862FKM9c+2E1U8Dp7mRM3LF02
JMwWqSQuIzTn65JBu0J9PEfY0oyYK3P7AFYID3QGuhtUuLD0lBlMuH4QjEwQc01h
ED++q8QC29U995drOg1W3Op7TSmZju23RObttlCXDRv34Y5RUL7sRN3U+dW5J5sr
ID78G1dphrCE4TOStK+LM/tzlhawTC+0LozZ3WNfTu6+ErFmLLOKm9SJFGeZ7XzD
c9DooIFYpLt342nPvPtoJXXQleyhACYp1tnyuPOdzuOtQ7k37d8TfixtJNgapNf5
VFk1alcSFRHLf14f5IiDqAltjWcy0sqVMVsp2SgthMHuJXpaE+YdlTbqCd1Ty/qp
xU+JA39SZzW+8bKZ/1v9ZI2ZU6eAeGvDhwhzRLwPCYdU2/wr//IeY8mH5bL1hTLz
28Vys0tsKuWql7RLX0I59lLQEijCMtcHSXJFmEVL8hqTaiw4Un5ymTCqjGLgmVm1
m/0/UrtxdXRXUUJqjlqrJMSJEsQpi6bmqFPaFIyuAvKlx6ZJXRmZZHxbGxaFJCSe
VvjbDgD9fBTDS5kY0urVkW40ob/AGcI3WO20OcXIl3AL6KICqZREFddS/quZeDyo
34H+1jd/s6N3D+yQyvRlU65fG0qtO2XBz3ci3o37tzE/Fwdw04aW9A70Dr8nKeFO
0Fn7ADyFyN+zr0NjSJ20eOzxD6/yYGj5zbqkG+o6mapKY+AFJDB4TfZZPgDKlLF+
ECtk6PF+UvUEdQpkJHu1ejVxKSh5oFFlPcRBfCr6CqHFDw3Dd4fzGWcDLdYzz62/
aJfuiiBZQJ4w+qd2C5acfXXmBvCJy042oZwdBG0J2UoDTk6X3a5ztjZtcK+E9yjL
efkl3xIwuLqhNeNA7a93XlVuSyhRJv6AUpuGO0gAH0iWLyGMI1wLY2yQXRP2P0F9
Hz3M2oN4HXE+njxCql+nNNGnNFwPoWRFkspOCHIDBlOWlTIiHa0E5IpA1o02AcJI
tnL5kJEvhRHmMwF/HTPZ+55DB9jrB5CYNY6q6fDm5IuHaqB3e0D1OKIH5r7VJ4iM
SC2IfSq5CWRk9/3WEma90ZCR8umN9CeMn92ZEV7dZ5ITV+/a56+cP3Ickwjq84l9
Rx2oCYJG5qkWFQQNbmQ+g3P95c/sdv3BWIdxW6niFxv8Uwgpy5b05X2c1vHbZeXS
hgJuXxSqK+j2anCU3aVRT4mJxHOALMP1E8DWsdDlOJBmhdEgSWEBSjB5/Be+DQNR
CMBMBP0ZyLDsqB2VLZWffqesaxle4z1pnKbnPhmxApHZ5Mj/o8EGJK3MtTfXABih
ZRckcwFuw8ZC/d+Qf59Vn1pjJKaDLOhWLniDroLG9t4KjGBf7gahOW7utTtFCGpJ
RnS/4Li3ahiLieOYoY6JbqTpmYbJdGmZ8p5yOjYsdP8Afx4nsaQ5MLJRHngHqfVp
r3suhedhmOWiUo9JiFsqOF6y41xF584rkwAIs4kpnd+xCntkjgl57AbbcOAeKIQy
45j0pYc6y4sS+oGzQhwRckZCJroxXqpg/Ve6IiNydvUG+iqnH6CYSqZOQ449xFJQ
2M7vRHtV1pNHlbtebFRKBIbhHD8akfZ8sbOCxqXu5aOIJIVW50CCxVg3YU+oac83
A674QzBjc4vk86cvMe6vPlCK5VcOHsNn7ECtIV8bqnRTJ6nrhMGg6yfd5w67zvek
UPpjagAIA4aFRqWp3PdHl6//IWAYQRid156hQAEBvUbfow4jTebdiBJ6rq1URcU/
fRwMV+MQmCrAou6YsLgY2/v6+ot+wbtZ22B+pGH6nIKLAKi1LCe5ntAIlYk/crUz
BLmLmdy21Ml9AFwp9+FqV5/i+d/va5KxVV+RNHWPhaf2M6B+JxDoWt01hK1u2q28
+Bl7zu9vbS0vS85GD8p1j6Sp+oQKDGjPzbswVYzUf/aXktBY+jzX2Nqk5C60twIS
pVYRxEMm8+EIEQy68Bu4CngDHvjQ9WsF3PIDHVQlpyiLeHS252DiLlo2/89cWfix
YKZILn/JvBLpWbjIa+Bmdm1zoJn0XPq2ink6UWu0o2GrchqcZopcEJ0T1i7YbUYd
D5npMKIeh2YPj6/EiMrZu5ZHMGgWF1j5F2VGsFAarLJET4N7etS6RmukHHdvXApC
8Qxo51d72MinedYTTBLsQ7INiMwfQweWLRzzudlzVhqUpOYIbt6uyLXtEdj0NlSs
sCKSqeEyyvzolPRjfd8hskMfypzBZqMOq2e0AX22F7lfENgkOeGtltFWQT4X6chm
eexlPWDS3Mm8/BkdZFF04xHLmjdj70zb6GRf39udWurjjZl0oMUoY6JjmpsEv/kh
khv/QuKCJFomCkBWmXOJ6HktlXLLY3ztDAODRC2up6WzKAFGpFnKlovz1AkW5wph
F47LejHddFWXuJVPa+hYoOgyNH838M+UaKfQs1/lf/q6pmTZlgd3VlzW1fnKVE35
/K9RXOcW2HDlrrKsghcTFjVjyVTjgtT6zE/jn5qNS92v/YCvR08jdkZWB8QUjFnN
hGHLbWTkRNgKjircuFd1bEeSEgNS4ihvnz601hg0w81CKrvGmvyQmpQll8JzEx7B
bMj77TpnAbhAzNKMPTrYaLhR1w0fOlptnlG+M2BZGvK7W07Z3xZR0LMNQz7D3RVp
UcDXinvYwUcQ9Y5FYjUHBNai4hzwU3tlhxluQt/xopTOXQl/xaQrL8lU9oy85jzc
zklWtq6+x/qKfiNzPONRY+eRDgaTwly8h7TsWd+2o1dlqA5RirdX78X2j4CZEgId
K3QMcZV6XT3tucVxRPHRheoarNbjerdW2pQRYp1XUe0QBJKd+N07V4NtI6KgoesY
8wDai0p88SOIjrzzcrQfPZ21eaHLwy8K7rzCq+vniWW4F1Gy/HaFqPMboylTeCTW
hhjocaNrVw+vng9KvirBBo5RIE8OP3xMW+azmskh43VpJTZm17TOvkn2/FUci/2K
xMgptuRBTnumkDjhZ5PhB2I1uO2Z3zBVGyMJEbBlXD8BOcWd/KcFuoCuyE/soW4d
gK2DwupZFmzaMaxHEC9zd4Ybis7z1q0W+s95MXZxBB2jI8iDqsnaygq7+yJpzYQz
aC6EHSvun+W9IXATrlfQ/S2PFcaGpAeMiwTAV0xj1kEDaYsjl4KLfKcbfNXBvwQl
KLPUVv148rz0gj/JQ5a+g6b00mt/33cwhhHqPWku/5d69QAnSA63n8ooRLnALmZR
xjZUFzHBjd2CrHBirvVBMuPgqOoIQFo/G4ziGYsjv/1arMjl1pXdesGN+2VGCB1+
JyDOvJrYfRh4ddKq8wTNJK95B9ake7mxQLrPeq0estOrAJGHJqLxu/I5XPfTsDHl
dFnI/Bml+CQaI6ckCgilo2OHptal4qvrsGJ4K9L3CoQnJTqhmsmASQHU5swWN5Qt
U8VsJunM+/jHaH4yroJC9Dz3CmlGuqJDGBeyF38s1rTHNHbCqWYCxYaw4yrPSQrl
XNBnQnhPdS+6Ney+TrqsXCY9gDXHy93SeVGA5WElknzY6OWC2MOg6Wimmz7wZEqE
blzBBXNifL1aK4MoiNWr/Yd82Ngc9F0o4UmbCfGrGyIpQBRJl+62vo374g4Bauin
NYp8P9npcv6W55y0e6u0P80fl6zaIk6nTLXGSzyC4UjbCdVA+ICRm7GAaaiin5q0
spertWRdIM/fpLoV2gatzhzjXY8KSFMa1lcI5nKG7/rJGM7qJKgJXtsxAcTLvlW5
y8HBWRxJSQGBFd9iLXsYDVI7w4/QLZ4wdKvLQx8ZrkVkhxNpcOG0LAXb9oA9q8im
xrmt34g9SZ3TMujITU0sZQe+ZWkATggTeHfU1dGfXk8uj/AtowABIDITrxlvU5Rg
iMDXFD4PaVO8G56vCYGH7sib5kJMP88mTE3AB8L9tFF3ToffjdX0+doDB0ovYUid
hxtktRxBPqt+39NIHNojYfbsE7HwHWhnXpvRmQyyZYk0kuFx2gDzX2t8LpncH8qV
ikEBtQppIY9Zd3QhtWwkGvKk1netR7KnJoB/HQ6IfZIIVE8UOAkD9FicT2tC5rVM
SaSp/aYSpqL4xcK3bPiTa4XraeciEYYlztxVprZpA+i8IsBCWG1BKh1omOvzNrQg
BmUuDYnhr8w4KWImf0UKC9wI2KthFSHgZwOn54VdoMZCsEPjA27dbQoL7A0kJc0C
3KInD5WDnJ5QGtdqen1XWuS2PNqE+YgJJR/D4LZL5SpPyNvT9dlljSUf1EfevZjB
mRm0C6gDhb+KqWn4xo+YHJPgObXWGy7oLO0khkZFBgvvs9/JhV+Pw/iLGxqAYPiS
tQ424Toxyz25DToDqsL2XNK8OV8yUSYFwPphmlTi6EUj4woeTlj6SvrrKXwKp6PB
LwEiYT1ocY2t8prAOHH1ZortQ4iofIQF4A+SKZxFAVV/LOvUs6tXxq3Spo8k80yW
RcwP0CbkPjH7tYHestst+UKLSejRzP/nefXoIh2WbGUdDTyU8iBkqE3LnMP3n437
VLd7T9I+Rh6ertt6KPFwkWj9VW6j17FoSjXVVFckPewvk0LgRewF/sFpWh4WSM9C
K8jPN3kXtdwCCrn745NLJ1iLkTfUjwvuhrmHeu/cXC7RtweFDmGWBVdpAQqSQxQG
2xJHtzWy0k6iNWCxc9hpIF4dD/Y4T8c1Nbr61zmCxe3jN1/NzpXrGLJUi6a1cokn
JrFacjl3fFFiFsh6fqqAbE3M+7wj832PTFBJIPKDOGbQJxUuiiV2lNbztl3YhG3j
bw1lOfS6Hlre61ADJPssc9UyAStVKC1pnzOR0cv+Saa9O2NN0d+OyciC5r7w6ePX
7mcuhIvJwGlVgKaGgGluIS2fET1ljv5gAuhXN2QZ92/r7sZG7o10CMwn53B0+bf3
Xqsgpn9dL07ndpCX2l18e8aVxdok2H2tF7jx+S0+9uNNBxJemDZ9iItYUdH2BWKF
mEZmqeiKTXNHXOqmhx7b4jyLWBBS9H283PkLsSd/uy6b4DO2N/fNBFh1YIT/I6IA
F00JxCvN5NAimRD5FXMHhr77SRuPkr4jeqFDkwXlsaiQIxnqs8ntJjn89kRyxJCr
CwLChjSBSpE31jJLBKCv9AjcyXqt0PEcHKcUMsb9lE5FE5fhNTsD8qNwIiVMqUKg
JrdB/8rpZxFsNGKnTJzSyFfjTHpuLYQxL6ebOEVMvUWCJpRucgTD5jEXINbpvTSu
CH1OnZflS/zyJoM655ervgDPlYfGE++5LBXHXYx3CkS4kogNqSWbY6cgDAwt2hZm
NVw9O+sy27r5B8mGfO6bhWaeEVQHXMY8sTlaFwDZc91NpIeISovsRkfWTBrKPYIZ
f7sROoruzH2VY/bYMNNfREKrR30pY9mFN/zvPknjME2oihlA2YGMtX1okDpNAmgQ
TR+Zu7fQrLwKC1cuX747CYIrlnw7E2fEIMX8uS7d3FqLP6QolzfcPTUJ2zLdySLb
8ltYo046jn/aOpUEfKCyEr191uuY+lUyF4Np/HQdyc6RAHlI4ys6NYOwbGMEssd3
Dzsz84TQ9aH/L63rJ4kv/TrCCALhc8AqcFXohBjOs+KpDS/Q0ElAO/Nl1B9y7oKv
2kzeBmQrrWoj4tn8k/WmOPTRSE/NKg/wrM8hqAq2vtlYbqUVWyRhqXYRiAu2NaQi
5j+i45m8XKffonCl5dMaoJPs9rW+9Ci3SURXLRd/LDgjT5GX+XGsJbcZy8ccmhBt
QrdKFQgUnL0Cdp9zThL+p26W9n5SV9mszIQB3bRzCJxxwAkdKJxxSNleXhMR3sG8
aClOTFOu+uEL3tNzlI4VeCg4Mf77EJl8HpXZfRFvRB0hBlECWPp3dBK+AsQPSSup
gRUw4ClYNr2a6RcY0u3RQzsvJJy3k24GTvnPqwTsqRacwwwqzBm6Tm4Nz5TexrmL
+T6SJlvNMO6Kzm6EI+/nAmNPxJfbAAAPZv+B/qfh1hJ5CVMdBHwmRGVu4NQunkXz
pXVDpr5+URKrpipF6dc6XGSFwmB/L/3tln97LqR2h58QfCbCH8DdkmdGMTqvfTK1
8q82MXnLJuCccl68462n036Xgy2aCYF0NV71BhbSrmvPzpWDKU0TEV85F6O2e1rU
679SdLD0LJ+6OwzP/kh7/rBOgt+Vt+6LIoKQBfVaW8YxglNMlo2yD+YIlN42ynOq
6oFWSzB+n3N49L+ORPSnpMG3s+2cXjXRb6dRgxM2y6uw16E+q3GrxZWRyASUR3iM
1Nyn224MiozU0jMzEHJxqhMhxr+5TdYqkxJFoii1BLT2VSnooZIs7H937sy+dug6
r53xBFQL2CZJH7lFCzakS71Ljfv4Cl0lr2zaLEOMarRRVx8SY4jisttzuddV866E
D8jUfM+gzwoTJ5BltFBS7luj+2PD5puwTHMS7n+4+4wwudBDCxiLYu3FMeRnYctA
BuY/n4dWL9WP8D4APmzUUwbwKx9EXGr/x9a4aMKhuVHWJT7MuvR2SFQ60+3Iwu6r
dWA9Gbv5+LmAKV9CdutCYDe5VgIR9FSCpGVZQnHAvvaWmKViGWVss/ucw+j9Pnp2
tDj9wpXlUT/6kN3ERAZXKl4niaZGs2UlRhqxz/1O0zmf01QBXQYY7hHEICRNjwpZ
wtBjPVFTiGr7WipbQ0XVVQqGbBh+//7oMMnWWdqkaZYi0/JWYr+gtTYfYN2TSSAp
YZvhZdlv4HkPpxOtmyFcSktBY8djIC1xpwF8DzhPuMsg69yeq8JwfozLVffFUjOk
tyNs4xYQqfS9lpYpgOYi6CtVjnNHGY6yBw5dgXtsONk56X65xdMMsfir9OvwnWio
jNOeH4cQFSg/IS+AijfABAPUUZXOvC0dB7Ph9MfvHFtGiOroWMCPeL1diTGbEbQQ
K9C7cWEusnesD0en5ZK0SxzS8X0rJq+t+zWpGOJqlyJmWqhDrd2Kz7DaeOjeMMwo
OFncTjLSfkiCTyMlkDf3Qv+hcE1OySx+ySVXW7l664gdUS21BkMIG7EPYATOtWlK
HSOcyxY6dhWV3h8FroXbGmuX4L5/gzu9PEgAkE+SBlSflqIIQZ6fI9REwYY5kdAf
S18b4/ugb6hTPs1nStu4Hxzc7wafvLrXJpMfXTeJu5JJSzyzTPG9nwaLIY+bkbVs
j3bZSLweD4VUo1BqOzBp+0amk9e3yksF9gHsYOI3jSc9GCBtdfT5oWkoKtTh7jaK
KPBwZzBWqKT2bt3raIlVa+kWpUeviY6Fh7mS9wlsKxWj9u1Yf0T9u9OhbUzeBbbu
bcQRYb33qnsUAgwhtedmH5ZKBqakpc/ZFAxrBASwsgmk3+HPy8ZSHCOdz/bbqXDR
cQ6aWtLtPaPPcvrzZTX/9do2+EzR9tUfeagmGotIaRTGdStyH/ygClnaCf/n5Alc
b7771kIHJ0WP8iIpnH8KGjTokIaZRGL2h9+KadDcVtkzw9GrTDzOSCWM3KKXnMHm
4BUCA2N8gtBzEPdphlRHWMGg37tsLxmVWk1mjTtUPMwmNofgAMK0p742SegPeIeZ
rijQ2U69fHW/GLXe+90wl1ZALrv9zY8h6tx23rPrcDw8uv4loVpnojZZSUPT/08e
4gP6zmUggNNs3bQgG4xRy0sgwg3DoCa4vJF/P7uRh+v6K8TxdJIqn+zpq2urnmyw
njCYpC4M7eDi6BljAnzEbkOf9c+G2O8OZFpNCMM6XBRq791zXy045tSugNYPgulr
hvBy6TT47ghjBM5a1gXihOvH1wd7gaXI+gkkHZwkhhQ1/Gl0lJw6YXLjxk4CDSpR
VCALpgVJj75BioSq7YmnFnVi7xzmqe+PSIimoI4EMFBAy90mMIkcjmIai2hOT2Vz
YAR7xjvQ6Ot6U3W/1mohqeFvl5Ux/82lfW63bDvaaBLac+uuAi9xYQ3Mvlh6UAkZ
7qquE0VNMgyj4rmZ904ugvd6sAopD0dd8TqcNDEiObgZZUNz/re7YjqQo5UyMw9P
jdVOU8H932pg3L9NqewaaYrDozRa27estX/aJxA5UDWH8ySPQKhNKXKVJFTonlzC
otMRYTq0MPPtjQyFJGfaGdwkaLqBNqHVjVyrYhCpzghZSiweUfXNsckTPnp2EytY
ga4Z6RQ8fd6VuKx419Dsv2dQqrOEjeiv1+Y1iqz2+2Y3hRzk+aRLrtJq9+itF8Tz
WQBknijTw43SQwjOmhsZEL5Fz7sy4qnyF/GUGsa/8Mn83iDC5f2UzPUQA3Iki8B6
D+3NxrYB86Am1aScj88Je+vSxPtswDpvmRDLUvqZOy4T4xTyofMHav1Hv97kfoY1
fIrP9rl4Wvx/CqujsnR0DTE2uJEU9VqKNjQ1+sBDb7to8njGj2EGd1U19cw5ygmD
NZIVu42g6Itbau199pLd5B6gYZ+ac36BPH+N0aYtfG5HfZ9kk0drHY0WADSSSuz/
Le2b0U4+3qUoyikbzKvHMGC6RSL7VnfN9pa/Av99v8XP48g4MV1EAOA877tVW819
UMtlXXrMxjRoWoz5lgqf01VyBJMkXZe70BgHYUlx3x2vOGUHqD80SBxv0Hu4OeUF
Ah9GmOQqedbTWUWQup2O4YLCOLM8rQxoBfxI1WyZOOCXcbVMMWnLAkpEp0xxT3Qh
yBRIgeQcDGJNaUqhEbczoA9dLDXaG8SS6Sf/LYEnG6jRi3dSAs4LxI1P3NNchoVe
dog7y3RnJ1Z4ClzSXs2fV0IDhAx0+7nkz3YXCFAXUjRO1Nz+7J0bEElV727K0kfg
NrF1/fkWDfV/iLSHTuQQcgfEb2NSOKR3zb18Vc6Fnndj8Bbbp88UtHTF8I4iXiQ3
xFc/5TsItSzVHhZ1IwED+6peksdamSWD4mQM/ExBVoahnqG3MLAyrrbzVTCLF1cy
wFAEj8niAlx3k3K5FaQL0y0ct7p4YWrf0UIPeTNt4Rg58sYxCPpdwSKbF+TzkPMl
xLjRtUqbEoN5XksvJ+nZHItXot+5PHVyRIB1/YgDzvYDaOLb8u635w5jNhK4jy4z
LgWEoXd8L3Dc23ggh1Vf8uPo+A1sJxegIwpvZwWemcXXnHm57iHdyVMXAE1rBs3f
hDQQjkOqrFNGhK0iHZF7XsxXxP5JWzbuFvbkQMjjsoNG8tA9BRl6YvZUzxl8AMO2
OmK1O1LvlnpfCWm232V6/TRT9FLGUxiI4thBzC9IaTlvUFx6lrVfn+K/LlOVbjgq
K39o9rbdK+iOtdTTimR3ZSfHHoRp4CLolGkaNQc+3BzoW7KIAoure0iu0/VXALBt
eyd8bfYhaprknSEgSmI4Upfirzuu52U0hHhUru2S7v0Mr1++FUWWKtkxIc1/shyR
TKJHgoSNqwYHPvD8D+4/R4dplo8OW02vjQEIvqYFB4DanRL8zSusPahtukwxk4nk
KCUztrqfoM2luQg7Av4BrbMYx6HJRUguF2EdZLiajwIQIBg9+MbvtxTpihTrqpjT
7iLf0xia8/w9UxVnG+JDL67q7hBpu12CPDaXE3PcRh4VjsG9etUfTGmczbdfV31s
1EtnatcokIOC8WFb+uG90tRgeUgfrKHg/qo2Eer96WXKrwLqiIHEONbCv8VnU9mu
GH0qqUtn/r3fSW6RNdCcVhBNsBm2uH4sGIznUR597IM4cKR3fl6yHr+zzHmiSUpI
t9I0H2G10T8RZSzGGESCp8uWklRS6WGufJ7n2DcWCdfeBGcu8C7pT4K58D7CpnMS
BU6MPmgR0dfIPxai+5iQcxuM/89zW4PkKZJhmEfwpsVJzeC2KcNEiK0tggwPDb+6
WuavLqHWKNSUC00jOLrBOIF5oAtgdV+QYcWRb4kiYwdv/qZS+0xBA+pOwU37PlTX
0qOlIvCjh+gxGgvdah2LSYFoLhn0AwyZeWD5LL9EGycMKqlb5yP1e/YMJmBNHTVc
jIW4HTttLuAHqML2r9SH3k5Y2WQk4ztoPfr2YuJ2kbrStCVeNAfGAU0H1h9Cj7zw
ObtndZWie1wPCMhQIBZQnSWIu0rcd8/vrJYQL7LJfY1qMvonTVBnJSKcX+36GHms
PJbuXb5b5ScXwwHkzvJk32ejvAUi9zNPnmu1C9pMhzjPoO+e2sKIZWlQMuaSLeT+
evhEQJKnTvajHpHu5cPkimG3967TSNtKqWg9RyXP9x08I1whDwfy7LqI2ZcnSjZI
N1CUCBV2okoN1TELugYlm79gpbPKZ/r4cccGV7R0V0BYstsUYwF2um8KNURaA8QT
y7N+5QPNjY9eUuz661H2amv2+N2W1sGqLju6e47J31rT/+MwWxEgVNy1rQWloDpM
pBEZ5M3UPZEV9JnDOFYYr80ixiqvjhUVz+9CcWzJQl1ELfnfrktOikuIpOGgWQ5N
V7XBO+GzVnO3C6s9kIfLmuNMBQ+zm+8Z8xmsMbu62hBwQicnlAgyROZZvtZf+rvE
3Gv307vWczuL6SZspmA9O/zP+oiLSjS5GQXayMzWOqm1G9qazSor9yq9PhKWhCBl
TUxWvY0ZmFEZ73nauIAwuIfwInHHoPTfxvTJ8OrSnqcj1V4fmJy5+GXkHaqNAc4N
aYFGPf4Uk1dWD7O1G1QjieE0t5xy+0qsTIQJ54mfq7N7XbK25+Fy47Ekf85rRwFW
04KPwq1O4KpUPntip0+iYKw69pXWN0mYQY6qxVafo1Sl4dmXO+Con2vcm8Q/27Eg
MYmScZFrt7eLh7Ib9uNTGN3NmTe+4sretgIm5jNomJtMN4V2vQnwYaqcmgEWHI9m
bziBncwqwy1tL5BG5ApnXh+mK/Tg9shBna+ZKV+nAZCd9KeZ613VZlghbwraiLmm
Ao4vKweHfXAB0/viCKKeqstda7jMfgu2gldMUMSXq3H53ohymHSabP4ESgHh2jPX
oJ1N4l4MNU+NLVcMGint1aYWllQ20ZDRIpaeeST8b8JdQvCMdFrWBgNz7GMPVqCl
ZtLMPTobfNXH6MbaRn+XKutDSEDmczvi7P0XPOhTwpRy+3Xo0AKswzBz/c8LhDSa
Gl3AnUD2i4S/yPuznLY+6e4zoVPXYDzsYsiCgrm5ewgHQsM9APGEkNyeerJV793S
IpzMVbphAs0c+V+hyZCJQ/c+FrINJp9INzqH1Mks2evgBW+OVv6DymQKtNDuJjG8
AcYcAS80HIXuYmyVF5nKteY4TXsYprvRHvwZSEz03AWNTveGj3sIykVyQckK6OvS
YXUw5teuP7d1L2XFxZWqDjLOKaM5UeXc7vUKAVka7AzvqNZb5/vDYb8eLupcZRW5
KX/1hTwOfm7F6EEQ23LdvW+RjT5Zyn2dKvcXX43qyGdzlo2AOnqDlL0S8OyHsVUC
lWoU/SD/hiPKgFvnj7BnUqLZF/wd5f2Peq143vQwLEtJAUy39Y/s/bCfmItI9kHD
DOtxaNomt9thr5ZY8H+pSPrqW5wQYQ6ci0Jkk7m/fjOfR8bba04ArO+IFpuiSoQ6
Tcjd1Tv1L4FACBDkMOEPaD0BfLXaktL5zeY5k4W2wHOi+SczzxAO/IQrlOsOszJS
7jO6jPk51sGNfdMq7Q3+GqsgA9evutAUQMcZTkOyENP1x+DEgoKyMHfefiwQv/LZ
n868SNJ/kOFWg80krEsnLvEABmV47YUjgJwwg8eEslIHXMQA/HsEZAakTHGIgRfI
Z019cmbJz/KB+jF52rr8vjSHiwDxyjSXS8JWUCAeicvNlQSbpnlHzjpvFonReT9Q
LcEw53kdiytPhsvJk1D2lR14Y09jfxR5fM0MdM0ZpCb49sBusHX/G1Xlr8QL2ajP
yhXmOma3gaaHs0A0kBL7cFC9lG6JWogWvgeTGwpX4OlGzqZ4uPQvfdmDBahtZmQZ
thKB1CK7Gy9F3OpEbIgO/2u9Id2YpbJLmWvovPrOaPz847G3PEGflAnvwMk+jgEg
cw95uNuZFFA/iG4rhnz71eIlIjY18+IWY+Ugmkgqpn/7p7+XbwY8ZEiBNDYY9BkR
bJNz9r131CMuhrHC4BKxbPzLZ+G95rLzz46A0Y/UJpe8c/blF9AXpSX/VVYOqjeu
guF2f4DT2MSey1xvsLPWTuZyK24BGQfwI3KTEuupYjzMMvm9yjzI7kQd75sdPx4Y
83zm5wsBnxQdeea5Jhm9bVyzg4hiJEi+YZ2H0SdseFN3PJRIDoLZRvFmTxa4f59d
62/Aj7WU8o3oMNCYQR7YA6Jkw2YlG1rE0qavkgf8BOWljgktHKSDyUHlE+oSlrph
Fl0QLBpY1E86G/wTQz1ouk4Z//XCj15rq61Za6GMuJXoHR6gcJr0mvXWUtR7Xxwc
vYLaDYnbdsRLDAaUTRsFPRkBl+dmc8RD6/HxEZf+9l+1EaPvb4k0mg0KoST7Whm8
gyN8YF+6fmhvA/errvse6x1jmRE39nv9hIDrg3mPzFTmRSdd/cBeuigP+LztlL9C
0AmkdM3zcoqVOzBc4eXMcmuA0B6RV7QNZ1Hre9fgOrReVOEjNf81yNEpf3a46KBD
tqaK5iC5Q6KB+fsfjiQUUTlxfy3ml62afxBTuJJN0774Qx+WmOPSiphEhhk+SVI9
iGwWbaWEJwXyC7pVJMbko0LJbZ+QCRAW6aFxaFGFZZSr8vHWXMBsDghjek3aeZNp
as9j6pykrANhDcyWgimq6CC0bxjPT5Yh7TkV2oRLDhZdlFszWv/V4XuylouQVQPD
XFHP8jAOAnSZwyQl5EnBiMrbPlj/ReqyYZhC17hF+M3gdhy/foWXBg2JvtHQFy4X
lvge90wB2gTY12+WLBBPTkdjscX/H68Gq2CygLKuFL/IJanORxz9HTjevZTEtA/X
I1Efw2f1DMVIFr+FkPj8gRZH2P/PC485g+CmgtwbLWDNjJ41schzQDRGiRSuxWpv
OZa771X9qIDghX1dkKpgIs+c526ro6LIuddF2uuW6ZnmOR1G0hPjkU+KS4Poz8CD
7relRz8rzpntDY7VviH5LdxS5oRi+g+sjm5gk4vBVenhXPMj60A4Y3yBDgTCRAu0
R3jIRLGXb56+3OO2LvC2/rYyzrT7b4hPzfVZPqPkysaoxttx/KXbdIRdL+xNBfPz
clb5d2c+QDhs55VeId5HHgoFJnGlW9G2BDIUQj2Ni/cFSG+ljjJxgZkebmeI/kxe
4Oqp12rmhhKJY9AIztEfEGytBHxrelLFEha+fg2Vc8yc10qMUrO3CbCew0mzp2v6
3SqONZJE6xEOcsCLIM+A+WZXLWYX8J0D2Kznkt32TvCOiMPW7y6AWmjRPU5h1xHW
8VLrFTQAObdeJssr9tkbmWWj0+2IeQmcBoXPDK/rXQc2b8IGPYbxSc7mWKyMVXJt
jWOIusjiJ40+zzFQPz1hlA4zKi3lgtgs59Hi/Hf37pXadaSDjb1H5MTTYRETGnnH
zqUYT98pDYY99N8MseyM/CNWkJrijnU/9mRwD3sPYigW44q1lMZVUYQ27BwKT+Ai
l+viKH3EdHDp5fsVSizndgDuMyiLs9DxAexzGYa3K5YTBm2Yo4KcaNFtsu4bTpgW
d5plqLznCAKd1TZPHnmSvQDMRJ0ZmMyAXPgLgJ9SLzh3LtZWqaSMtgc/psLi9ocQ
ns4sJVIIJV3kx3atVBhX38+e9HtLbPiLXvpJzfKKMoTCltzVw+hx+YZCYWUfk3D9
848Qo8UJQ98mdJ9TChxYsJv7K2Z5zEHsEk59oBKFikATIfg6b/DEuaFWG1IWrZEu
G87jCN8dD6U7eOvKFt0P95Mg17+lDquc0I/ACGMahwBjy/wVOfILp4Bt1cN7RGzT
MA4KVbn3VeaDHChazUy9QKIWZU4ZmIUsfceme0VSNv0PjbZEJD3y7x3x1ntq4swr
Itv+/5d+PZfDzBlWhJnO1Fl/b1WLmUlADc9Qticb63v5GXknp3JSYB2VERSzlk9t
ocHS/qUz8so2d88DMjwYAexcptMMUsfK7p9VVz7PZ9OIPVY037yU+pUPhl/hRwKL
Sx3wcxBixqr1FlSpCOv+QewmlIbiTVUTPd4iIbmnHc24It3EubZb7UcG7C/itoSM
yLnU4MkH73RHtuXaMa4G8yc9S/Vx5PyoTbWoBsQtZ9r76YRHK4a+mA4KhlpRgd5U
m6/OjqN4+2F0UjjeJdpnWLFZ9ruUhpHK4T3d7Ar0z/to+P4YSZXePCnsuWdFNUQR
Jmzcgga5bEst7NcWOuOfpQyaVvyFOhfInV+ES5jNho0pbeWSzwR8qvZvROq9WEzL
qz5L02tyXelcz2/xhCULz7p+wRKl3PAbNP1menKdkJfpQc3q+7+zKDFfhclkeCYl
eislKiR6vS3svZBNR81fKqtN2dOw6nPb/2gRJwZYUODOT+jFa12gvaA4PJ0zyS9Y
7a2MGTSs3Wdw/OePlWx4OY1BNDY9p9D8sdQm0BVY2aH23MvIbMVm2PDwf3/Jpd/6
Ph8MLdj02VkhQ4jqjG9evYZQfHBSsNUPtZePoteUzeKHj82ppMboHNSnjojo2Pd+
n3yt37/5JjixPJoPSOk7t8ShM6DrGeeMPQBt6bbReh5y3HHx0imQMvVtI1DwIG6G
DcnBG5IO0lg6yMMhY6PrGH4bmWLJfDIt0RzYNihmjTzCjb3pof+pfZqEkSK7QXkd
hxwH8q5xxL70QVrXDfbbYC2BUFU83h0Hi6CiIt3AQHHcQh8TNzmmjACOYoiUsCGS
WmVfrCLjzoaEkVW5Sr+aY3GUdaVg0Q6YPNgWGkHOolGPibksZBHXVMN12bkPzFVK
p5nRiTFigpNFpQCJS8PCT53qX25kNsEsVZxGHQqk2lFvxe4DJG+ViwpJayC6wsyt
L3FrahYX6DFJuAn8uPAKSI7ECrmPL3TJUV5lFi9q0jgy2FUaP0hBM4l4iNvyhgzT
2Ecy82gy3w8ZI/NGnXvrMhgn0MbKRhQVuExN7c7WbEiD/ZH+iqGmsWwXkqQXt9n9
JtVi1P3jJ0y0NQV0kvYpv0BzBVwpXoj6/qS+ZHOTumseQDiTh7x5VKUpfzvAHJ06
zNc3Fvv3p8V2EaTlFkLxZe4tEDxBx2vaMLQOKAtat2LdmSnA0jgl92EallufDxVp
P5owKf9uqhVYVaW2TsG92ZUOkJfslHpXvtINZR+QlwAdIRO1lMpWSyhH42yeq/r8
8BbG3pQUlGxUqOSoG9DBSu1BaB+uZJhEZIgYhyjsyqg39GAeCCxfm6HgwVhd2Epw
wCKfUxSBYSssWJw//CJ/uzx3HPbOEBudNDQfO2LTvHoOnDvBjxybnLu4L3y4WICI
MLMaLFflA9ki65EO5sY8xXsjIbNlWQhFZUIEvNpU+7ilahC8hFGYIOm0LRDX0DTW
ZKpi3wFfzZfL+0BuBym+0kskHJQ59KC9f7UiRTOJNQlLYnv6uA+Lu9cmuI2KIDJW
iHw53D3U/wpCJdoBDi6Q9mNDfbl/Zo7NoZA1BEY9H+yCZlJMJ7v5Ud4SfLSZYraE
A+0HkFpA//Mb0duxAuwtrq4TglV7pqOmYJWkSS5OpAlNKOEY1k/ytiHvnQxHPWuK
mdsekLaHSvb8fsX1ZMPEahlWVA03BAkIy/Leg+7LrB+E2Z7/7fwgH48yVyaX6M2Y
RZXB9pTUhAjMj0GmScCncnXy4c5D0ysp5a2mMUoNsuVPSGNlbvV8rN0AKYvIbWVI
zuzGaro9PIvLvZuvl5bj//hOTUD8shVpXc5Z283SsOWZfmDqQYreZSKQ5uxfLxOe
VC290nTfzCSFxOCfnqIxHyxRil5OhPZ3p48eRGZVSns9NiOxExxV+EYFBDaWGMBB
VGJ6PEZ8yzwH5xkeGN6XXpTmdo1q9WWIQGap10p4ISHj6iPzqZ1Eq2ccggQm/7vq
yW1LYbq8qgZHqmhGlpY2qqs/Fmn7Mx/kpL+YrfzlAyvjNuQZLXAKbAWbElcM+eMF
sMw7rounClPaheSmJrTCSpoS08q4VtJENA+mppXQqWoC3dj2MT6bhP8V3GZn1o9+
UtzvzmB3dXJ4geH+TPQ838Up7aFvgZUlt9Kwl6A5izoXd/Z2HWT2I/wlIVoqtNry
7lS1R5Uh2Ny9XXl0cPqFMPjImVR09yLVnet+SS2Yocefj8ypzXZxOOqzIkuz14Kb
TvM7mZIqTuBLXaJZvsF2loBqvAUwwsSpd5utxC6f2o/HckRqgrOU+v+S2QfKAFHr
WSSIlmMyhi/v45Xquj6zxPSP6Bx0jlHPf7KVWeHx8pnEWPr9Zpym6wTq95W9QezP
hH3wC3PliS67BH1r3Xkc+fUdMC351F2CIilzARqLc7g8WbxOJ0c0O+xct1k/s0Af
jxBJ1wDx/cHJdgmFT9e+g7ekhK0y1rGDmIKd18kmd/D29aTk/ih1v8erQLnhj13E
G5bWvvtJ186wpZtPtJqZOYJ3hhOJsPgGRJ60ESxifMdk7RdprjsYJzn7HX0pcGHH
5+/4P3IqVf6uJeftGpwSOjJVU7aJ6WQYGir8PU345TsNo7dk40mB6FO6EBc8EDTo
6aVM0dpVroVKVouFbJyS5APuyH5JUJNq9nNGrLoj1+M8pnhWciEBlAJJmINt4Jyf
xKXvJBK4LtdmfA+N1LRNk/wseamJXKxW45h4gjBveDg7m/29v9YX4IubsxckVk6e
LPME+zEBgE9LWOmoJiQp/9kbD56lm+UonmSXD4Tb3mAg462NGrwYG5NBOw1Ys+eu
Uq57mdBzVe7q25XcNGwl6Wpjlb09pXMd1kkz0kg8+UWx0VPDuASX19SsEfbCSyCl
JKqOFrmKpSHTU0ov9tmvr4vECaDCmYi6kCDX9yinph3hjGyKJVHCTjePF07rrqRZ
08jj9EPMQ4UizhB547Nih5SXD+zqKpOhTWj8EwsAUSnGqRqPDNx6x0FqYtXonjX6
VbTN0R6EFare9s2yEY4UwqLO8JWQVHmZhN4AzZlZohhMlRxWhLPFaYYn0MLoXQNd
j26x9EMD21VpMKACNF4dtzTHT22eR+EqLfa8BP6o71GmCwbCC0jBuh0UMC/pSqfk
pMrOwClPuUe7pOzNje8Df8r+zZucVah9LHitmsK6oxmE56Ln1U3vnnakNL1MTRHT
I5F5CWJ/NwMXgu2TxByyLvfsgalxR2GOQDPxXxegeKxfJMSGfGUbSSrC6lp2P57T
bq/qFNNmHFbbALCl9diWJUWvBP4VpDSGA4Qc5MPq6HwWm43YPqmpmqQ00mNIM1nO
wIoSddkbEzQkpmMAUTYExwPmqEHgAjxWRpnCmVvRicuckqSrq7IcybMwqB4FviXK
yPXppHLtj4EgEt0zumKbCdtoaatrBzVm2tT3//0/bIljCJecCro1STQ61fJ0jTY+
mxDaTXklmPWTmB9bSu50R6xcThRZgCgYWo1xnpfVUuKSQK9i6cTOy9yKfYbiL4MQ
JJx8IdeGdZkyKZhNaOK6CKcWsRk3GqKgqYPsTKTwndE2JzGPpxMBCJENP1PKl/IE
X68QR02d8h2B17ecR/KMzZdWRyrbrF1dFmYQOzNVYGJhFZ7dd2tBePNuytRoOIBw
Wuh9ucFCGu0MGXRGmwpIZgo1LOvmzjD8RfbZSsf/ntTBST5qJDdkBwlFseh4nm+p
mWa3JPSK7/6sUlP1WilGmfh4gVUIWjS+l9BaxYQbUAPJ5KjhAbSHqV59Q9Yusdt/
sFPGJOV3BMl107nzEnnqsirutyFX8C2PhaZt8Fm/tACicJEnR9KCGzb1LZjtRgsS
kao9BXAfZBK52hVWm+kFuVLYs1sxNnJlVSnvbtJsnycXCnu98gVBFazEthlrZ3Ay
RJLLMylmHJrRa9B/bNOqm6pHxOWQvW0QOKbpIJW0IX8Gdcu/lHnnONOdzw7OVPag
5+1+hXLFXjBDXhUbJSwe84vqxFnKgi0zQWp5f5NKlm7bi2SUvF/96+DYdnauXdE3
4Vtc87zZy2Xj+TJ1NL7z+yMXvbLVu1egS5eKYKe3L7xHbvvNA9HEkDRJAv8UPZT9
zqBwt/pJE73ks0oGVk8KlnC/uvielVljK1Tpza49KNWtesBD/ZO9KzGxapBtup6R
ibQQlgGDiXz39dNuWx8xXAHm7lhcUAyKtqB0gv5LdaKzBmOFWqWD9AKg0+RCb7le
DkCq5w83dyi2TNl9SSctDHj3/yhjf7mohj9lCuYYsd2ef6UtzICjLG0PmpaPYJd7
qFmDTX+/7DxWv01tHTTMWkavXelXDwZz5eI+KEmVXl2OfLv4lFVr6EMJQ3nL/CHE
ezbxh9HuTwx4mGuANfOX3hJVNFyLtTDdFAiseaIAQtXtpBk9VAkgtF9zQo3Zkay0
+/NUZtaGUYw5GrFTShKbR+gUfMojeCHNU589weZbqPml8rGhJa0HdigjaRTWo9/E
W6C2rMf2bDdsvVTiQ+Djj1L0D0a56cbCWZQQzPM3bBqBXrLZvITzGeFfYKJt/BuE
rWXnAl2/2gvHS59P2WnODQjtibvnb+LZoBgVeew97yPSap1RA36wqhww/mg/GtL0
gcmjUb/X3a3lNZ63iN97DI9pwsongzf2nM9ojMyiettSP+nj+NKS97Ce7EV79gqg
F636XzEaR6BiLlK/ALNqe2QPWWenYdAqiOcjDuPvH9dIjMM5BbVXYAv9S/Yn6qiu
Jh0G8tLKlKPQUXwZNQot2zrEh3Hn5DLeJ1VD1XANfIIGyyee/KA3TdRmKMwCLQD0
bVQhmwpJK+tkaQ7Ee2JhKq+5ogfuOGLnq04zZ6TWmUt9FvCGaFqN8EAWOuQgOVY4
ZAW24lFmOCrugACvC4g1rwWKcLGdPg54ZMDa/L/8M/TPYIwVF/nOdKR/WeuVerTb
WkUAO/l25Y4YYZt4B0DmVhIU83vXjL5OSB3pruVEMFPktwxntlYeJ4VlSXZNUQxf
zOMOwcrVHGxGzTTBT8eREC4bezsk3/Alv+7Kk+nHjhMkAathuYORlgiP4mB/0QlM
zJekO9ZbtcHtqputo+mrqILN2YJX2YuaYP49K3hqOEsnBmEGMD89swCK/eaJfWgN
Bmd+3EQfuJ40HS2O3piJLee8wTEGZ/Po6/vvd7DCIQ9Zxnvx9d52FwaBKpM036Gx
Ogl+hS5LBLt+FThFAMmVvz0+eZWNX7nrDtaWEWhzjd4sWP6ufLM06dvhptUV7tul
8dACnWnUfwKhXsxCl0rVtYAd1txAx2nRdK+jq3CL6xQq9kdk/cNkgvg9NVXTCZ9j
V26H6QSLtu2UKU+iEbnyQXKbRHrl81ATuc5i8oi3NasHUDkoF0Y+1A1fO/MlTsWU
FkwD+VorT4pLqP0G3z6W30Miy+qAoTyispXaSbssnS4xwN6PxHkneEC5xXg8Nzxx
6NXM8SWyiaEQn/w/1IE5aAzYoo0c2Ez+ysEj+P4SwdLJhq8o3CjY70WooVeYU+2w
p0nkuh5DpY0o0lQn2n51+cGP06jRrJTRmWzsgwNLnYd6FLYgrED3MreZ1G/Q4YW/
WkoK8GMn3F5SJe74fk7hcmLhnW8Mrhex/9yuRDO61qeWRIy/1p4JNIru+5nZh2Ho
ytleJiSSX1L8xZumX36lJKCkw8YHvQdfbeswkGSaYUu+L3HS7WM3AN91LMox3Yfn
1Mp6US2rmQYjNhQOotQB1uZqQSmOFVFGtdtsrtBy9/IcmhvcMRPN66yVED4spPmY
CvHUJfe144qoGO/LbjjntfVZ6hNzpCLkmhxh5JxGxAwRzrjTHRTxzet9VyJ4vFTS
ApBBZJtL8wkZyiTvPmCASgX3nIsOkdpkgULczXSBHXyuloZpDKi4o847G3joTTVn
L2sT4v6GEXyCy49FQNxIqmAKzGsDFl4az7S1rz4ILujnkOHaiNHCaJdU4aDTQ9rG
QuN1ue9IP7+kifG0dHubmKcTle6XJv4nLJOXyr5R4aXTcTfTnnydPFBHID1y4258
Wl5m5vEH9y0rhgXZvBB/gfEmCm1puSlFDX51izMiowUDDyJKMhM4Luj3x9l8Ay20
LizcIbSNERxGQBCZq9uMl45tpNrD3Cef9arxM4lVvz9Y8AKQ9x27u17BqjQGSNkV
h/Mys7geGknJecz85elAfV7V3v9jVLlvceHIadEDC0DP6KnhxGGYbMwiYmPRtxSK
85qPZVx95/KjNV/YBqD6D272qNhNnf1uw7lhCCpDNKUofkHNu2TVtka88k7tHMiP
sklcAelnn6wuaKteUYKqAoEUEjt3kp7A5MSF/Xl3qD5TXt8zuHYiIRZUnC8tYBdC
83BEOCN8sNqf4+5kLBb00ACZX+J2LEpVl/Xq36Aa66J6FqAab4q33jBoWwRMD0tc
jA8Mi/kBT51f1HE2hPDc9xtP/eizxNONFD+YQWSnkFLqhuGUei4XoR5PFZ1Trtuz
qB5yT1COJaBg569+XXQsV1TNzf9LDqmOK2LV59gWRB0KOb0Yr4G0ig6iIqQMWqRb
xCh0iIubPevxXf27N7bJ0dRZRESwKsfW6lMSnONDX1jqVWqmpLSjZRcpfZN5rlYJ
w6XFtZxtYhhG1MNWod4GSximSsbdBkCBikeUz14/WBi/JKSgwaOKl8+GRujggeDx
diyYcqfZ1aYUHgMDBRQTOLUK+2U+qIU0MNzrPyTv8djoBUjeIRZ+HdHJmd13dZ5i
bWa4yP1CY2U1JTXJ2FVVDYiM/FjkcUaInInIF16SLrNJHkhndvGLxCzhvldyvCBQ
lO4Mm3jQi2o4bVY3aTwpQpPyrZmJAKeZ2BHcG8kiSpN6/LHS3Km+wqo2GRQ7xbwW
UyPDZ8VB8AJyHbIGTW4MB7Nvoktkpm6/wEWo6+fAOF8mbI8cdH9h1ta/6hUh+q2l
OWbdIk5XWIzSIZF4Ui402FjIW9xy2+/4aDPk2plPKFHaDBIjR59AciBSUBcaAeRl
sDN7DqKgpj0JoA1NNPobZqvNfeKsa2otdX28l9N2B3CabRLaMPIHHOeVd8wur0u1
2blqEZqgm7PTSBNS+gLoCWWgu90ot9fvfwWa3UvX+tN8y76gKiKKTvdqMTRlLH+u
UQRceCcGcaJIE4fYYyv8OfFhBKyBW7XutpKoVTgayXbLidPA/u/Fp1SZuIY1fs34
G8qhWIHfVvhqWX+2XOOPf9Pw/6ZEyJZXx6c/DM3eey8rW6lyjJ3IjbcR1Q/rIcRd
pcA9RpFlenznD1FtAwpruqm9OPicTbvZH+/CZkHW4Ma45ThOBMT/vgBjndn+C983
3Q1tqGevRrBWyWNT3uhJY2gPtcr0OOsmpMBNXsk/fRw8bZ8C7UWkShvqnQ5YFlpB
hPr8hrL7C/GYg9qZiyXdzwSebVcKvqEKxO8xVLz3OcyjUwLTf1TroJdRfyKW3MNT
HIOtnUxKChzUzxKi9koOeY+Kq7/W68oW6cMxgJMk/xLi4lTYvhNHlOWY3LwrEvtg
CqnVRckorXbLi1HwT1X2RK1ZrxHZdIHmt4bPeM++LrqqlKPxeCZBQTDfrda9GvUK
bMbNEpaU/nQH/nNZAEtqWoQClojxJFeKqUp9bYD/95Pn9yIcIXbCCtxlztcUcMtJ
D5EjW71m5DevwtrqMKrrhpky19qFpEl+0m4ST8Y4rJTJGRGKcP7ON1Zt6tf1E3aB
OYzG2gsQ0vC2Rx7ku/kDUcbHUusQnnLoO03HxyvaA1DZLtpjarWdCgilT13wyG5B
nmF4ti8mZtcoZebQUwL8QnKpXAk0aTZPCaAipdbl5VDx8d77eSMo1LnHVyrDmuoM
y0CeHhwILwwu6j6y54cyPeNJilmjqB/DPxRcFHyeCf75rqSITvqQw642sy8FxV9t
Gw/m27WWJ6rP8HgWqvuhOpeDnN6iRzz9tT2+0ZTSewWWmnxsyaBOwxnAGa9WVLT3
5DY7yQpyUHIfXUTuVwVfrHthRLIMjnvXzy0uqcSk/SQZgARRjhFMOZoZkbm65ycG
brWRnXFSsf6tfmSfwlx8zv3a4aDQOejT4sto4rc7VnTGRDF6GCmJjneJM3XNaRJS
AMVHzVVLYU0lCXPnljQkiExBaZUG0xaZ2AQYNf5NgqgGZitw0oQgcdG6rOuhZtfb
mMLhFexYhOvC6IhZIDQig8DeiapSoHYh4o5YkGrtN2l3ajWM6X5FQOPV4BPwDTcc
zeBzrdJZWBU3A6n8+0ZnRZGYd0FZ463aP7C/0hpbNnpH+Dy6wfQjZzghPp/PVpk2
TFkV2ywWsVyC3SkXyaf9kyXAW4rCphFPAqLS2ADaxAaYaIZoF7yNGlK9Aemoa1co
/iGtABtbchHL/wKEbd/8+Yh9Yk3j4hW5FYiyVslqFuggdICdVTGhSWe2Bcx6lG77
2OvIwnGjHupO4nuoMyzVF3O4ef+jpbdRzU8RHgkIEmrGtZTsfsMvhhH64ZHo6Pl5
rBj9RSHL//JI3QpLRd/6Eh5+ZGfKZ0CZoNRTS/xTWQzKClrIfEyM0wiUedSpasMe
15W3b74ZnK9iihoaUWhDeZi6JooqyYh7/BrBH0pt+ENrT9UKVA9O4pFNKlznBbQV
cso3SFEwONwDqLOu/2Urt2FttxMwsKQ9UVM37BYGnq/b56QbzXkSRuUK46r4G5P7
xd7XvAvlMPjE/Ntv1WeUrvUsJNmyOBVBeXci7kbbW2OCexZ5Malp84gh2N/Qlf4A
0U+NkFe0MxyU28QFBBHCb7JZsPLXUENVUHi3YurejwKA5y/xQm5ZeMF2KLPecXL3
04rxhNDOY7dfl4hLgq/qjMpNnIWFUMjDtumY6eUcLKMWsbR0tO4lihetmkizc/27
u8o+AW2kal9Me8iuGjTeLGM6pefOSxqDCAAfXGtOu2KrrHXCREXToEBTMKk3ERqb
1WisZWysUiBIrm0ta3A5pxjXbCaqPCXMrKOBlKLXxiaYSMHt1kp7PGm64X0ub23y
oTRAMi3+7x0vxT1py8p3M/8j2Yjpe1XcyhAIw8ZZnMyHxkZKCeOASL52Z6s06Ez3
XRohABjWNschD2fvlaGi1DWC3emWZNdCnBWCgwBzqXXRpo+SEwt/TUyC6tY/+O5g
Bj4fnUifjry7qVzxaBwwtZzepOwmgOFhWXTolH8ZPxCG7bnNOOW84weJrvTfkkp7
fSJh2wsxgejXDDnZIbRWvoLHvVMHBdVNk5LbRfkv8xZz/gZBHUOtLWlZSuQsbXtb
KH55Nw02pc60En3b1q1BMMU3md4L/NiXVxstwXTnvEgx78OHuC/tXi/olrbuIpC3
VtCt6g/N2bx/S9j3set8kxFw2rClgcEKkZ4Jow1vES+j0Y0LgO1XE4+TtBXablR3
Kux4EKDSRP20wQ9cmU0naFONL2Gz6PVXv4f2KnCLVpJa574rHd+VQJzGdShjkJv/
t1d4m1CsHhA9bwwQV5/ekMibPfBFOgyF/oNmo27ZLIP3KTULhBDn2qyMQsBBFecP
Y5G5Xw0uYSsWZ4na3WNtkDQnT35IBlwJw563OGN1YBxh1TVvvj7YXqboKlhW53dh
5E6DkVMbHiUIrX4q0XWqE1WYHRrnh9WZ6hSFFvyrqr4jEBDvGLRsA0Mzbpz2wW2r
6/4PtqYjNz2JGsJA5AyPY6CfRno7DfieMntIdRpPVeOyvbWmRtbDOtbrF3kZPv8f
+m4Ok1SCAtixD4L8FVGKSrrHACwOJTFLqDX3gwV+6yeK7RSHa7dMbe8v8CFOK1Xs
C1J4uhnOtRLhP4x3j6J94G/fcBG5f4iHMrV8n87ZaQRMTYZwtX3zHYGBNNHP0+kG
aJuwnKJy8OmJTCC/FeolhpD6SXqy2g4o6IBD3o+cTGspkE63Ghjy3oF+sT8jDhZr
1BDAOcOXd7i+xwVFd4NRo7uj5Rids12kudGdcOIqR3RmzL+KuVbXaHn9miFK3IZ6
LXUfHUNIBTlZCw6H7TM9+vlJXbSEB5Ajn+If1JCuwyb7H0Rjw/Es8pRuN1yHmcfh
AOGhs/20n+M2jNS9si49IPGzC2UQkiVvAkiyWEN/3PazyxGfYeqTjgTBqYYKZ+qA
ujVlOOtthUIYeHOzNcPMWPllyNwqYmZtErqXnWl5RrtTOBJg5msmCSf7OrH7BZaa
N6fhMynnyCN8MYRnNx1zcyfXRrYd0nJlM9KHFqBYK6GGzK6ZqrXQUjXTfs9fJLBK
1aQbbfhJR41M+0ZvbyBQhL3vEeJ9fNolzvDSKureWAXRXNoGvn4P0bM1FrXqL4to
zDlRcQOx4TSVuMjmIWfF0x6KeTTjl0dnmtdxvjJd/+OEABHcEVV9LjlzuIMLihoL
Kb4nlKdfujw6c0KPoRb4SMG945zuVr3ol4y3+kKzGUyhUoRKl3AeBGlNwaj9RfeV
m/tf4lnnaXTnk4hEjNnXVRw1+J34pa4NnJLKuSbJXMFBgVVpj3SluZYRRnQ7zFDX
WCJmKromo8/2+aWPyP81QqVaQvjZR40aW1s/FiGXG5TRzwyDgBmNfcU/SvsR48s4
2qpEYe8DOeVbmOS9wrGMoGqvQUSY95/sFx8GKBzHXsadx+77vps1ZC9VOtI+civw
SbXKtc1zxpx8KDuYbPDrwh1+WJveQksCoxX0H+cNAUzWjgNDjmssFhq14kYCHa7m
+KvX2W8/OETt9sbOXaSTdUcJ3SBmM0uz2THeDqSdPbj5ZdnLE/stf0VQ/gZKnF2V
TQ0PgAR1wWsAxPEbO0xlNnO8XuJ264WdQZfyEFvereskKRpDWFFkYqZAp+PU/5bh
a/zy3vGvOEtSbEjGTwX1hL4Z4LbEHKcnTpeAv47X/EoJ8bRfq/SJ9joS8ySiMHez
R2dBjdE97I2021EB20UpeBbIzry/AZePeazWgDSBcsl783rsnhjg/N9wsIEvucMq
IPay1FnCc+JXy+rLrl/YwCj85hD1skMNmttpFKfOK/jpBfF3LeJTgVGX6QcAWurS
ITRzh+3VujsmbqZzm0+X5Qhc4BqX0NejHywwpnS7bRWKZCLGtLsmhEqs4VW9AiwH
3Q/Z9MRvKqg0ySFYUAfXgrJzs5QIyPQB0ePyKhYHETGxMSE0Ey+0voynbTNTuOCq
08HPqp9d0Fd06/SxMqRn56tb5SGShkymOq7oUlyAQtM=
//pragma protect end_data_block
//pragma protect digest_block
peBI46imBq5Sf9+/JKa5QG3JScY=
//pragma protect end_digest_block
//pragma protect end_protected

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`else
`svt_vmm_data_new(svt_axi_port_configuration)
  extern function new (vmm_log log = null,AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`endif

  // ***************************************************************************
  //   SVT shorthand macros
  // ***************************************************************************
 `svt_data_member_begin(svt_axi_port_configuration)
       `svt_field_object(                      sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(slave_addr_ranges       ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(dest_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(source_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_string(source_requester_name, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_queue_enum(svt_amba_addr_mapper::path_cov_dest_names_enum,path_cov_slave_names,`SVT_ALL_ON)
 `svt_data_member_end(svt_axi_port_configuration)

 
                
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /**
   * Assigns a master interface to this configuration.
   *
   * @param master_if Interface for the AXI Port
   */
  extern function void set_master_if(AXI_MASTER_IF master_if);

  /**
   * Assigns a slave interface to this configuration.
   *
   * @param slave_if Interface for the AXI Port
   */
  extern function void set_slave_if(AXI_SLAVE_IF slave_if);

  /**
   * Assigns a port stream interface to this configuration.
   *
   * @param port_stream_if Interface for the AXI Port stream
   */
  extern function void set_port_stream_if(AXI_PORT_STREAM_IF port_stream_if);

  /** @cond PRIVATE */
  /**
    * Updates domain related information for this port. Relates the address
    * range given by start_addr and end_addr to the domain_type in domain_item
    * This function is not expected to be used by the user. It is called
    * internally by the model when svt_axi_system_configuration::set_addr_for_domain
    * is used
    * @param domain_item The domain item corresponding to the addresses given 
    * @param start_addr  The start_addr of the address range corresponding to this domain item
    * @param end_addr    The end_addr of the address range corresponding to this domain item
    */
  extern function void update_domain(svt_axi_system_domain_item domain_item,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);
  /** @endcond */

  /**
    * Gets the shareability domain of the address specified.
    * Returns 1 if a shareability domain could be found, else returns 0
    * @param addr The address whose shareability domain is to be got.
    * @param domain_type The returned shareability domain type
    */
  extern function bit get_shareablity_domain_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,output int domain_type); 

  /**
    * Sets the address map of this slave component. This method can be called
    * multiple times to set multiple address ranges for a slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * @param start_addr The start address of this address range
    * @param end_addr The end address of this address range
    */
  extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);
  //extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH:0] addr_attribute={1'b1,{`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH{1'b0}}} );

  /**
    * Returns 1 if the given address is in the address range(s) configured for this slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * Note that, "addr" provided through argument should be untagged address i.e. address which doesn't
    *      have any address tag attributes appended at MSB.
    * @param addr Address
    */
  extern function bit is_slave_addr_in_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

  //----------------------------------------------------------------------------
  /**
   * Method to turn static config param randomization on/off as a block.
   */
  extern virtual function int static_rand_mode(bit on_off);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);
 // ---------------------------------------------------------------------------
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  //----------------------------------------------------------------------------
  // Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode ( bit on_off);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * Does basic validation of the object contents.
    */
  extern virtual function bit do_is_valid ( bit silent = 1,int kind = RELEVANT);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern do_allocate_pattern();
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum value for range check done do_is_valid().
   * The max value will either be the MAX macro value or parameter value if 
   * paramterized interface is used.
   */
  extern virtual function int get_max_val(string width_name = "empty");

  // ---------------------------------------------------------------------------
  /** returns total number of address attribute tags which are enabled by setting to '1' */
  extern virtual function int get_num_enabled_tagged_addr_attributes ( );

  // ---------------------------------------------------------------------------
  /** returns address prefixed with attribute tags for corresponding address region as MSB address bits */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_tag);

  // ---------------------------------------------------------------------------
  /** if tagged address is passed then it returns only the address part corresponding to the configured addr_width
    * removing any address tag attributes appended at the MSB bits of the input address value 
    */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  // ---------------------------------------------------------------------------
  /** If indipendent secured and non-secured address space support is enabled then it compares two address
    * attributes and returns '1' if both are identical. Otherwise, if indipendent secured/non-secure address
    * space support is not enabled then it always returns '1'.
    */
  extern virtual function bit is_same_addr_attribute(bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib1,bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib2);

  // ---------------------------------------------------------------------------
  /** Need to enable enable_tracing and data_trace_enable */
  extern virtual function svt_pattern allocate_debug_feature_pattern();

  // ---------------------------------------------------------------------------
  /** returns ID width based on port configuration and user requirement.
    * If read and write channel ID widths are same then it just returns common 'id_width'
    * Otherwise, it returns read channel or write channel id_width if rd_wr_type is
    * set to '0' or '1' respectively.
    * If rd_wr_type is set to "-1" then by default it returns minimum of read and write
    * channel id width. If use_min_width == 0 then it return maximum of read and write
    * channel id width.
    */
  extern virtual function int get_id_width(int rd_wr_type=-1, bit use_min_width=1);
  
  /** This method returns 1 when corresponding slave port is same as path_cove_dest_names_enum  name 
    * and is_register_addr_space for particular slave port is programmed as 1
    */
  extern virtual function bit is_register_addr_space(svt_axi_system_configuration sys_cfg, svt_amba_addr_mapper::path_cov_dest_names_enum name);

  extern virtual function void set_cfg_for_rd_or_wr_only(int mode = 0);
   
  extern virtual function void set_port_name(string port_name_);
  
  extern virtual function string get_port_name();

  /** Method to wait for next negative edge of internal common clock */
  extern virtual task wait_for_negedge_clock(int mode = 0);
  
  /** This method returns axi_interface_type as ACE_LITE if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set axi_interface_type will not be changed.
    */
  extern function axi_interface_type_enum get_axi_interface_type();

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_port_configuration)
`endif   

endclass

// -----------------------------------------------------------------------------

/**
Utility method definition for the svt_axi_port_configuration class

*/
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
j5OBsfhgFLO3dui5+xWUugAW2j+/hF7TSfRwIKD+zB5rPOct4SDYF/+xmKUZUHcN
hVdMqfPqRFgSH9+NxqXbwGQGysQPLszNq5gWKvE+xsYVdNGGuB6ZdmY0Xw5/U1TZ
AleBhHqw5kaXF02DWxgoV95+hvy6bEMkktdIaM5E0AskSekJb3HjGA==
//pragma protect end_key_block
//pragma protect digest_block
23leOV4MYFmDxhcOPuBusMDe/Jk=
//pragma protect end_digest_block
//pragma protect data_block
CNEUw2gIRag94OfPZXrEKHb6ql6TRhRLWt4jbP8zGjn5AZyv6Ik/WGBXBP/Q79mU
ypQMUQlKpJN5vHkT2VVrsjQS/rqTSQewtIyCKFTFmeUaQlk9xraJpOp/vd1Vf1kc
s7hBYxZNh/D1ni5AjTVeoi0L5iuuofD1tAFXiZKuYTp1wpMOJpCFFvsXKDkWnhxE
eHpZLUjxI8UShyedZELoBhdKY598ZoE9edMCL4eWqeszIrmFaURuaJiJG+tG+hSG
ppyUusxjuo+36dV3kcJm8R6xtPt8IKg+E9b+zI7X0236/gfzCyQRkwErVLtPK80n
hRD35ItoJbuLGjf7drIlrUhE0+3klXaZ+8oraFE214cZk3Kj9LV8P5K7gxqRNdiK
q8CyEQ6wjgHnOerjQANQyj4eJMtsSY355C6mskOLuKyWl2oI/hE2+uiCjTBWBBe+
wS1h/NPNOt/60ZWP1OjluPhD1dJQs7Jc06bVsfi/KA10ypgFGJwdVnd1IQjIWcLl
htXCzh2ZPfKsUWZuvSJ4qPZ/Ysk6Ha5Xd9i2qoXl6eFulphUAgYU3iGneOQ+nZhb
l8PvjFxDF/rIeiaoTz9RA1GG7UDQFZvjA0CelFIToxBL/CuZOCWlK117/E5ZzxLN
zB8ZMiEa5zHnBOtSMkM7M4KAyjq7H3jgaGn5ti5RLQk4FL5+eJNbaJozsAIw6Ckx
zMGWawuEmtDops8sQV2ujBt6bg8Azwxf/vXSXRBZndYZEnKW4h5P78Eu9Pi261xJ
K9dXug7urL2CV3Yqv5n/V8oEp/qib/ShWwbE7LyZzAZMBbL8TneonxClvkQSCbgs
fs4GwIbaT/jlGQ+EmoyNvbyz5QzUBpyYoiiSjF7T9SwprApPo7CSTjW7YcdYTHXk
X9BciIM0/L4SvYF1FJxraAkAWHnx7II2hsMa7pj2BoE/1SDPqeSjQ3PRpLWEx12Q
D5K3MVnkdKa/5Qo+dxgFzxVMKP3Y3qoAbMfjLG2kLWi5N1VaxqN3oOL/2tATNuv/
QRMU6SvclkV6TDSZH3hP71efmRQypNdDF3+w/a3bzwtfiYpBwsq2rOBwfzDcY6v4
KrSMTQX8WPAdYRSLM1DTLHRs+bBcU/2OSeWquNXdJDwl29LjrXSb4FSARepDUsrB
osR46STnan2rdRkNm8lVMAkr3BqldLbjkbirGp5Vt/q2cAZGnxV90GdDBI+63yUk
Ilod8YqDV+HKUVFtX/5kW1ovJ7YmtDYF3jFVjnKBaiKhStkY0IRdcaGdmLQnBNxY
9FhMU3msf1GaTjLwHXiIY9FMx3+MjYcCTZjRmfmJT1rinMSsqNj4uwDlM4I1o1hx
BLIWWSQu2o+wY4G0xBkHOzEdRgX/+VAWnYglYJqDFuE+RXqvk/uwO1KPAxENmlo6
oHJLRzsLueAiDAUC5vvNMepClcCTv/ANtG/A6QWMpmKyTucd2VcklNAsrxLpuLNQ
xqJESmiN1ddp9zGdNYJ2pySvRgF2kVOwkY77awM2+5Q1NBkhFht4WD87szBHE+kJ
IxgLTcWgFtic7tPyZcxWPRtZ/8LjaoGkkMdR/qqrFgob5NqMoWOn71eTM/wDZYSl
lqYesOof6llFaoawNmy9Yd1v2x5x0T+Sa4/pjg9D/Ow0S9SNCfyr1Lr2U/irK65f
6ORpRaHzTsMgjBxnXGSPaFaziiLSlDR0u+iqOa6AnabTCuvM22hmbBxmC+Miqbtn
TeJo3x4yTqZ1fUQI6pBAstlQWXVkSPWEuHR+UeiQQnsAjrWmb/eY2PkLuZxnNT8G
rrjEwZEADPmpLI89DWPJkIHQUSNhXk9CJYDZZEyCz47mwzD+07aw+/213vj1WTVG
m6X+/f5qc60QT07SErx1w6w7yFb/cu4sC2jTFYlc0Dii1Uth1YTtLaB0dYGm3vmp
/eMT40kuN2S8RGcQvnYVeD/vlgIFmZEwrhBAyYsKLsbY7eeQg5QEt7hj41a0bOmn
O7mNrTlTGfAahn7c1d6ZlWP90xk96FlsOlyuAWm79Y8hG9ieGheJ5eEObsHrPa5Z
sFrdqe9n3awshll/Jlg8q5in5xkXamnix3tPQwAMT3mOqeImERSkMmfsA1S0964j
r8QGQoP4g3k/+X3SoKBtxQpoLHmp9J2KazIcMiwqFQpAF4F525BxxmeF1IoIH5PW
bRgCQDCYb7pHXqvk5+S9bjSfyHpVjw8ZXpHEApRuzOIYF7yq6zOEwcMjP/OBwbtE
S9g6SxwWG9DYcQGzC0DcvYpYDMokMuJfA7fGWgDgnNvZ2l31NbsJhTPUG7PG/xNO
Uq77KFaZIk3FDi49F3JSQ77pxRuvch4/wMbR+Gd8Zd3rTpmR2okk1cRYT5X12gMm
nPDYfkw4VhGQDWJUPXX+p3ekGGED6eN+/DH17ocfktCc2P1s9icemxLV/S5Dd41K
MsVouXk7qXHdUkNSTaVAC4KvYPmnxNYZqO/QgkJx0e8k1eHyrtWpRmC8gH4J0f8D
puhW+HVL4m6b/YsFbzTJckh1erv+9+DE6lNgueLm9KbF/Kiku42yNJI8tb6iHgLt
PJshVXcdMmMYW+u7B0tmUTLxQjR8IhczELIZzKJd9rjCeSjPgTwrXx8Wr3Zksd7B
egL3f7tEKxFxe8RmySq0sycgEgEfV37h8qZyu8kTKczm8QaAUtRkbm+fPnUpBiZ0
bPkeM4Vb4OXqq7L+S1HyfRqzu5iT9xip4iBCLGTypdSpoR8w8xHM9TRnPmLOnO1q
1Xnh3UFNQgryJOyNOy1OJVPdWuzpso84uRWk9Naxlkrla/wwJXYM31mZx4r5l+9K
SjODIoR4rp3k6L/1vGA7DtM9m2yPhrdXse/F3wFFVok7tmFBGVwTfXXfQr5JhMhr
vYvS/Gmwb2VruswSaTkatUOwB0P/RNcG9VMN8xoCIJxtVZUFZBGQOrmehOiVRYiL
sLgFznbo3VVsb15LINeFo8WU5q/SjWzfo03v4s9gF0yDpc16/UN8QNk6wBmWk8Ta
c+9tWYipzvhU9NAGwLlQbvV65EU5MhOgkzgL0HEFhoO4cNMYY9e/6DMyxj+9Fjnr
7+uajdukRBT81Nb4fJcRJlpNIWzjEX9SzpcB04MUhbMXv6cI87ki+FherUcpQUXU
tjYSKQJp7VwT8yPaAEKvspy+z0qZQQKtpCSYPnAGtsPYh0eEg6SGLM60boWvYqQn
FhGefqEmKS4Jx8BF/38dEo6/Wu1P3OO109HWiu8YydgJYYYpaW2qk6TZW15Ub6Oo
1LAPiN67PPyGNWPHlJChlrrNI75pG9O/r1F93/gK+cZeU3M46QGet70pB+X7sXtz
WKFy17S5jsYQuoE8mEsKWaeguwq7Mv0KF9x6KhwO4m5ZFrpaipk7C3iHjuBCwRhI
FWpHjYeNP705/QUlemmNSmUL8tTMqa5343KyLRZFFkoNXyWLn+JDQ9eVfLp7G/Pq
h6aOtVi/R+8ETACcatAnSjy0YkQQ02+5xotXnVK9ch8bsTUuopCjddQT8S9dBO+V
V/Aln0jIHP4Y7zxd+hHqLgo9H7YIl3EEoLSKVlmS+5uKitCCKXXy4FppnGE3EcOg
gYEY1YiDy/WdVnKEc5yN8sZeOGuCKSAEcgRa6xBV4MtOdJ7pDfzHTNc4nYUO/MEr
1pu65jqWqBUoGysDZYx9R5y4Id2ImBLb+rzby20I/wNoqDgz6foHJU/3LfMml3Wn
aftQZdsYDlAMldjx+CxQivV1h2XC6hgugiUnAYa3Y0/MqwkX6aQ/HiTH8O4u4rZN
nipHKvrzWg8InME1J6QTk/BPtIcDMqkqwLVU5cSXU+yR939eSCkaaE5i+tZa55j9
5M74xEyfx6kZr6SoInlBe1Q522vn7A8xTiwByAh0hKm29MIGZZToiNHHbYsQZ+0n
yBVNXmSFjihXbfwo/kqCjsIrpNqAIchr9Njjkl0Guc9HG368bmX3q6jGg1ZRw0LP
MfBfZL15m3YY21G5YoOJ+KJFgGGjOkb/kZWaGKn1dsoLmLqH1H/d0OUb4YbAnrVD
/tiSkzD3yHAjDCfT1Wbcdyq2QWZSEXviq9l6eCi3SPJNEmT34e2juT7offxGViHP
X/1ZUHn4EjF9kjh/hx3v7Nr72cyhG200CITLM3LgzcXLt8buDdUzb5SevAwoMqFR
EVYknrgrHaGXkjYyVdJyNZ0aO5subgX0e7X9Kyk02xkbdVmPEgMX3CeHb4XlRw58
4fZvys/rh/Pd562fDQ7ZIiXjl5esdLtpys3QVCuR3vcpQWy5RzhdytzmldP9xQ4E
GpUBXc8+4kppDvDHEjiamqnSwVMKf6AYiuXJQ5vRqDa+ZXxfi9hA5pXfYMBxONrE
G88c1JDBY8wwi/IjFvWWvfdQQJl5PyP4dcsZVbXYd9KzS8NG4a1ys7kK2jdHUm11
3kGHPEmo4nDO0ybYQKy9Z117G67A9uRIM4y5RmHt1wgM6MFWu1M8eI7uYvF9xT1j
GEdzMyZKa3f/WYhFcVUHHVa62fOLVlG8jiqp0t00wi7xUIFGyK6S5BXW8LL43Nti
0EEkCr/d4u+ZG5YR0Su5tZMhrFEECOVr74EBFJTqnRYOkPcnx6XLyU2SweC0MRyf
u/iVyfXw5S90hfDbqfJUi1KpdqhkkIgIEuVPWlrOsrVSn9A0f4rXuXPbUrNA3n5k
AZgQJ6fc5ord3pFxyCyNWTNrr3yeon2nKYzFoTjdL+EwqjFVETNpGIAwiikI3OZI
yiCKxSAllyMPh5DRi4f4MhuaNvUsoN3a8TU2Cj4E/mw7mxZdLsahnrHLotiteg2h
OPIYwAfRvRkGahtH0qoYCzRLyJ4FBLJ7Nmd++YCavG93y9acPWuEURGACE1N/MxE
W8ELvymp3fOwYKCRniRHYyZb7xUs6/jOxC1WcFYXn2gnhny6tc3Kv27TxsN3vwj5
Yy2vTiGrL49FZ1KqJwdFJWSuv3P5MDHrlIlkgUiG2RVipA5WUxICP2DESDxFSuMq
Dqc7ZUSxEDiww95/ZFlBMnojOeRgO1WOC/XnJ4kSMqJerEpIGz6ALq0j3JNoq9vQ
fAo3JbvqA71hSFhDRw//Vqe+tQF/Auig5I7TtCUnOpg=
//pragma protect end_data_block
//pragma protect digest_block
4p0bCDGZIY/vFETTR6iLYuH3eII=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
`ifdef SVT_ACE5_ENABLE
function bit svt_axi_port_configuration::is_bcomp_response_valid();
   if(bcomp_signal_enable ==1)
     is_bcomp_response_valid =1;
   else
     is_bcomp_response_valid =0;  
endfunction
`endif
// ----------------------------------------------------------------------------

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CV/8Nb8BgqE8MB835DeM/EJ3k3GU7nxvsqA8mQEmIqb+ZLSUfdzZrbFXEdf37bXa
6ulX0AjsKLiuVE/iv6QyUij6dp4VUltcFPLa12rnbd/g27m5+szDDMsefXld5pIQ
dpnm0WKUoYlJ050Qcompzhw3JG/Q1BD9gWJZmMZkrirv1vWxIa11rA==
//pragma protect end_key_block
//pragma protect digest_block
ujOVJMieri7xzXAsl/kHtoc8CiI=
//pragma protect end_digest_block
//pragma protect data_block
YU5alE4KbB4wHYZ6loHJ+mThk54wvaEEtBA1sGmY0qT1eB3PtpdSQixtfnQIFiIi
YkNaZMHZsC7s0XIGi4r7AIfQMVXYANutGsTPzgKPojbisO6+kT0JDeZEn2WioHpP
jxfwyFrMguuiOKLUH+GqQ2pKzr5xXQv7WUqgYE20z7ob/FecHbPr/pOhcTHpVOuG
1LTzLuRJvjJFnCqcQCWxIKfek2LSGv2VT/pn5WvAq9PqL9ALOmUj84sjH/BT8dtw
IffDq3Q5udX1rzIs00BxoX4Q5x7752q6ImbFrokclmeNOY9a+pAlpVDU4377F2M8
9v3VHg+Ki7ujK5mmYpzJgAGrH07d587xYSqIra7YkhNatLOxdMHF2/HaVwI3V4t8
U4VQxHCrtNmircT2FCnBmyRIoR018bgn5ZVrqZhHqNBSiYON04GwNVVk89y8ZlB4
L1EAlGu9GunFuwBtbLw9T9VXRCfSuE0DkSsbyqnCJqVfk3N+puH/GY/cAtYxMLk7
UZ4pA1XCpgjCFbmLJu7pEKY0ZJQGuCEnFkOWUKQNG7IMLnzKg1GbfdUGpWXaIw/P
mXuQXfPOEJpsdLNwD4S/ljpl4jUYVMakduOCfFIIBCUaYbBq9peWjPH2MtXQy/Kr
dGPqKCPCZNY5s8dTSS7ga/fA9Sd8p+MNv2Pt3ci23CS8kBl7TB/r/1cQBDvqotjT
nWC0JN/84+RMetx1VkYIJ36un6GXB60uqy6aa5D0Nul1Dzg1uVOTxbzpmL/TLe4t
Lt2mMRSFpJrjKh8kakxSlylAccLlj2BqG1wDPzzbxHJX3acZS0hCIBb97uiZ3hwI
CSOSGNE3Ld0kL74LookMb3h++HfSZo+sqP/tXyUhP6ZLDOpOFeEsoTXURzpeHryg
ajV/uomeA8Wduor4x8z9Ht/jiO6JEyQCxkmQ46/wcxYU+Dk30mPN11yA8tWqwcjT
OR+UHi3uNdX3IJ+izeANAUsUgnLdyTgyKKgTzZB1uLct403Yl6b0BR5VlXnKDmSk
DltoMbzcyElGW2vyyDaxjU/D6ngOOoLV3tE19AHM2u5zI10B7skQ0TvfKTYlsXK6
zybB12x17t1Togr1qwu+I8tJXV1XHVoaabtqgpvhH8IE5934Depk+jyKfNNJiG4x
z2mFWd+3l43Wfy3FOKD9NnkZ0w1LDUAB2n+zclg7+HQgXSCqwM2rjltvrPelUBQT
m8M7M//E8us4WvIq6HMcIiRaZN8bNl3b9NYenIR/O4p6X6oFmfF9EB26BPZzVIY8
iOHmRT98peK5eRzj2NGpXCeY+aWfUG2XjYAEO+EdfMn6QC+paOBcd6c43MElUh8o
dNECeLBkvys5QjOiQ8e3HTRVWu4fLHgjmW6PFu4bbnugDBOGawzHzuwGfjugYKdF
P9xuB3AIKA4EuBWXF/M+flBnvXMMDOW8bLN2fG6mMnIXi/RJ5d/Nc0jsNVUO6hdS
1KzNNBemHlceGPDv+L6TQzrs3rruFwhS0hXhXXpNfXYxxXZuyBm2Rl+d6bSAxVSZ
x8VcafNuqV3D/b4339JX7YGv68j2m0tR0nlTHMKd/KvngaK6VsAoODLTg8kX0v/I
71/bZgcdBn/TC3kEI+oj96UNLX+hyrLzmwzEOxJXs7aOmIh4xffa5v+TnbwRv23w
I2a5K/KQ8XFPi+JiKyM1SVNNFkeD88mVIFtA4XMj/181QI6roXZAceOH01P6t8VD
fvoIF3vbysUPEV0nVTs+x27yCM2nJZ8TTRL5PZ4v4tDcwjGzKQRGBMoxCMBJGTfj
lvcQh4opchWcbUbC7euLi7GBWmxCFoaUy1sfyYIvwIGvsiyacsFVh3DqCZXedZNf
5g0iW5g4ls3nYXbWY3hpRzDjDFKRcdsPTpei3gHV5lNs4lVXXTa2cWm5fbWIFluG
AMl5KXJsLLw0vlRNb0wg+8yX1+A6h0eJaXYEYBGAUfZwuCGCwkBC9mi60kW2ds6j
Ow3SxKBbo2VdJAyHvWcWIXbMSK1qbhUoEG86omO6rQjSl7vv2JgM8vpja/L2HBKY
lUJgy7q7kpAK6ez5ay59kkgGnq0MO+cPWqy96wDw+pITdlAA/3lICBZlvso/L6E5
jEoF1/TmPV/6QR6O5YEnY3utMj+CD90ffWd6EjerLLgGL7sMycUCwv0xdn4NQTqr
lNlnXnP/kQkHEoEL1bvdHEeQayIzjriKYQl3cAtZ25BO0BFMvxkEwI0sXdRe8NST
z37pYWAmfVBa2W9xVKFnuP/T0QEz8uL8jxzr0vIRd3ane/Py+k6WcZri2jO+bE3j
ZCDw0T69UuSeWk3gmU/edwhslXxIMCFjwxDydv4RbYJpdFY3Y8iZp+gkvDxMEsuG
H49R1DGGpFzo9jhqID8uVkzAJ1NOCQxxriF6z1aLdzgPM3s1yrBwI1jIrs6jE4pN
1cjy3gSX+ZUgu/BQgJsrDUsOiaFfNhCooGIRBHayNiiglBHcy7QarBrlUMMNot0E
Ogsu9kAnLkrIOPCIEkvSoRhImWji42aiOrG2BZHwDlnAXJ3+gdy+U8/gUSaxfTKh
7B84m4EQjVrjZ3wa4FYeEq6z0uV4xG/l95DntVtefl2pAT9wXSL++Rr/3GyRqRZe
QPp0Vn8FJ/4K87kqH7CcSrEjQrTI0r6MFryKK62+330bDsnF1bL0ANHcgI+R/hc5
ygxxqhfeckm2ogLJPGIXSkInZ9H82GirzHLrzOp7LCuDfaJg+9MLhL7EQRdLbU5c
b9s5hEtIXl6mdTCQmHW9pOhrMGQG7eyRFnCaDIGlRaZ2howiTrPVESfkgVT9jIQm
UQkl0RXOVg0tEEdgNCbFKDAeQmcO3z9opHDgVu9EHqm6l0N+dVWUkFvCWrdzjQIL
EidetXH4W7Z2m3ndXbx2LhIqfiUsrkXKAht5v2QSyyreBLfR/TULsNVinMv1/DGl
VRn1alN/LnPKcj3rLMp7bywCrOBzT0uyJSOEQQhJUwb9Ay1F/0liTBUshJn2I1DK
5d5IGD8Ni8qYT6RSG/Sw20yclw2zVpzKet9r0ARPG8eBwFTb9wVq5KQpe4WVjQ+X
5WA3+xBZabDQ7lDrRuDCqrYnTfDb03M2nSFZw5l5dJ4BpKhvrf1FlUClh2UD/yut
eRQ+B0PyxHf+rMcmj+eYBbC9vcn7WT7+ERkhb1ZtxsO3QDA3LTmBlw7yuWdbEw7w
hmDGt4PcTzbEXjdJrWJXIAEKIXYoB93Ce7RNmC2xGMOXut0BP36dRu2ThJfJlG87
mTVHshcLsphqk6pRfBQdseZhTOBQIVOol/6dgPM2+hPbatQ7wTU+xjX2xf6wyqSt
4PDy1NjlOSofyMpUdjkh0fyr9hgnFqZqKVKvrVPdksVGgMVjSltWa2pyRTUe8fjX
b/LG7+Yxa0GMUYR92ddI37f+Milsfquady4N/q2rYRS3XxtfrtHwS0vuBX0WJjbi
bcRv5cXcVaU08Xwg31no9DDufTvTSzgwAl8i6ClH16Io7e5K1FFsU8DEr5BXPNiP
KuBxlYO4QJ6g2JHyPb6BmesdyRp3WYxSCyt0DWGJx35SOn96e89qPNle0kbIoGPD
0xA8btSZBLrnp0mSzJSSL8SB4sKu7cMct1WJDuEqHnmwjS76ycttbPpHjWc3xNg9
SFw6l2bY8TbNAghHoLtIgdWJsiGBgBE0qkCIHLLOTWdAsFTUJThuyGXV8fckHtyQ
6epV0q3ud2PYGXnV787xxzY4/GxObBbiL29at5oS6nNB49L9zPAMGlBrL3kGdqR0
GGjUCyDTFIO1c7+lwyTJ1fhYABQj2eSO80JFRCDXOBuJSn6GL9hUZzcyCamgYO5e
ktt+rqU6/XiEHRToNg7GJDQmiOaMPcUbixsJiAmbZAaX3D+yh/+gdPJQd7NU6ebW
mrLbB/jUbllzg9hsSidf4VC2YfoKp7aJ6ZQZyxdeACHQfYpCO6WD8nxn3BEDP5vM
a4lBEpGV2BWiaV9i1fchIA4vPjqRPlYkHmMD5QVLwcDW5FmIOJcRoHGFt6fL6nwD
e2by0QudVm0bYA+wVryG+PscC/sTAwbCTNYuAN/lTQRTnX/HBAgRuv/T+BXW7PTX
P9yPbC92+1y9ELRcG3nnWdLLcoKIQOL62Gu3MkNDbcXoA4UHb4wdI/pzr/bZAt/w
01EwrxkqHVlmdUXLGfpUkUYasovpM2b+nmgX4XWIEN9EJ4ygs0t0aGyN/kR/sSrf
VRrtRK0Rqca+jyLKSSbcTxIKOBCni3gn269gptEqX1e7hD1Js8l3vZJZRSZJaNuL
UV+bhiZLCNRIh5KA1mK8tsRNmWHU1hPqACWjs4j/fsLwyRyuAnv845EBE1iNG5Xp
DvYewR3N6/TDjhpOmIEHoSFxmqMTYK5VqT0K6942WbFx1zDp2fkIk0Ii4ngqN1wB
19ztsqOrMhrdoEig5UBz8wJ4FI5dKDLb/DEFZOyJKxStRcQUMQlKXfX+omr++swD
/LNAlxu+mFS1O5JknuWalaAG3x4NrCCyYLBM9xhI5Bdo5y8w92G3ETxztVxSCakg
Cc6ux+WwZX1o//eDZeXUVZqJb81NxLZVzk2A10O4VAswW5rs4ePA7XAxTpP+aoTt
FfUopdLQxDagIznyrxHRtvSPuEnozzstVAJqkSkplBVPNqQEqGE1v5SjaSW0L5m0
X2zhPH9OSennkY44lRXcbBajKIrN2xzLfEzrDqaRuw53qEEWS8I4pp0suzt3jsrx
3SrFp7T1sHi1Qu+Lw8PEUbqD+XcZRM49excwnYUXfNOwhBYVOZOCwpmM4WEI5u1E
BBbtNrxmcO2B1UunZ6Z2pTSw3FXsmqn63i1tMeb/GzoKNM9mK43d/SofCYG98F0n
Uxzitp9xJv2Wl9z/xn2HabSxuWrZhf/b96CUF7eS0u8AuJL0sDRKS4INEkD4sc3/
QnqqWalTRbLL2SIrmq9d1lwWiZ1diVC4ZohZW+nMziT/fBuC7mhErVQG5Wl+BD6u
tgjU8sV8lrDCCDS08xyTATrF5Ng/mRHIsBh1an/9Wk7ieBG7qKz3s0N/sTpjubIu
v1CxUR/3yKrmL9/kqx2QrMgqszLHSt2zHqSOSV/QqJoqbtEC8LeXmLn04guNpoUk
T4GellZcXe4jxfpoml1jbBJ2PQxXWSqEhf3P0yfjQSqDcWS6TfT8pFH8kfS2FNO4
ulnm2J5tqTJtrj55aoh1cY/0hYVwclCyqP1i1aCIlFhzawpA4MmE1MHmuJLAYchJ
OUL4Nx9yLScuG49v507aFUULJpyS34eaN3kN8qKKZ6o3DDv0Wk7gee7E7NGQCjiL
ud/QQqvyTyjFZQ8/+CzPmevz5HCH1d07O9NCMgQJeOccal7xELk/phgLzU7L8+kS
1QEqMePtvVyIdrOs9Gh/rfQtx9NUXJh6p60K7vf15t/LJsS65K7YJ9fy7fxNneGp
ebWSfb1osenBCYVsPxFHo+3h9jXtHvi0T5XqSTmVSwRaIFTj3mV8y6HZ8FhoEYw7
pWAQQENTErskw7qx3++Nr4THs3FGHDrI8WAO7ze6Eyh89yN0FS2B6ZvavHvxOASc
bd0P6spTupfeuX5xvPMD4qeJKk3NTS5jp4EN96NBMvgYTcaFktyyCWvhtcS9Ee94
B/q/6ksIeSNmB1+Z4IUzubUlDPSiXJ1p+A1vxTFJdf+PJiiSulISUWIuT4Uu2ZvT
LMn3dhE2hBgwNNIHGq2NK5M6wIUrpdiSZHU1+GPwB3VfILHafLg0rnBVWn8laG4+
C2mfuNRSn+gxHGPS50XVP0NKSC6426rbR1x2b/kUG4OwgwJq9WeVN+e1bZRQUZAw
udrGz2gEU9Mo0jVN5xrXnakyR+1Z9Hbkz+lr1bxmFJPj5siesVBFlhaZqLz81tOs
Nth5mVfi62kaoVgRxRSsR2kGhcZ+OR9xWjrhhTIx5H29o4fhJzvYeY2Y3FJOuQuZ
SaopeIN3m34QqM6vymdxegB4xA7rtyig5gUfww7z1wqyr0R/GbTVWBwYfK+95ria
mZHJWYxoH+WKMV3cVoj4Ai7mmtcFbbGe7BOsMjDbEqPxFxLE7zIfsUaXyyZDz/B3
XDDVqEoF294XyjLwxzg5XUpfRiA06LCL8ByGV2512b6cAOZsBU8drRCYZ/mNiQBT
bRHWtDdDELw5mtdq4+s5OXt5PAGF+d/GnvTjbjkuQ02ur0tVFHQxbxfEEctYELng
3DQhI9qP/e5dzkZHmIi510TzYkSl6z7u07Z1xv7c3soXf+LH6bHyZvmhESwvas3J
F4OAYodnuzM1wR/li5G1VhdaLA46RURh8D8VK8sM1bOKqGevy7Ug6VlMzC74pyIA
iy59KAfltLkbhOXl/Ilk1Fcj9HegsSW+OOYSsmnKWnvtjyexVAxV8zx7XSxm+vLO
kuGx7qzHcHA9k9002vIu4dMb2KFuGJJx3qqgb5cbz6IKkGCjT/7MTP7CJvn7Noy6
at6/MfK2me0W1tNQmF+5Ihoo3JgDQN5CtTnDLUUVWwNDKgS6df4w7S+4FqfWCKMS
zdXqG+APE9qndjVjK1DCdJ/i6KGCZoMNQpsGb86BZC/fpJygB1Wi35OIt4fZ6GLU
0Kfp+sZ35OqlR1iaqdePTLDu+S+dXXYEOHEvUTV2r8/HBP4Rk1dceogsaw5ydgGM
e0+ObKomaHBu0wdwPy1SsuyZ/wPMoCsKFTLsKKUenKqWhk4MoXRWG0p+hdT9wmhh
6uqqZUXfVtqffiGRQBNZALjuABezoLXULZrDGMcnYeZJzKXESDe41k+8d/2vfKok
+Tat4cKC5G1Ixq0x7XGJzChy0TAEDuJvcjodBFYKV8CTtn33XVqwgUfFqFfKiRtR
MLrcPmMrxG7pT+InuPFPISDB/v+1fuOlax1WrHxzaEIr2DHYjuRiWxgezAyFZ1dC
2ONKvyLWcInQ9zzphRuEGgrsecVYyIbR7irVzgMvwhKL2B1ekuDBC4SsrHy4QsnM
BFYX1ndl+NZpcWSBi1oeMOl6G87rjjqE2wWhvyvcuk3/X+TcLblkCoGXVcI8CpFJ
yfThnysFNNBMZIOHLFsfKY7BOmbCy5QkNeNQw+ESFasPwRUxzPufeYzRFOEk4pyV
ycNZtGOLMpx6oQQHHU7Jz2Dwk2ffNeSvXnUau+wIbZ+p509DwZfNieglH7vDpo8b
MtC4HjHzSCjGU4e98nylzkrnmDaPGMxioVs/mw6NESELtSCDCiqEYXF4DZuZOSIM
hUjc+peSMewIgzdJ/k3QY1dnXtgjOsloPie+W3E4769aTqpHEF4mFW4TymiqUG/8
l/N90eAPKlwDn7GhM/rMX7hy0dB7kDlfdEKRBDerXFyH3Y+KzR91HAPa7Xi9BATH
sO2Pxe2X5knplk9RbiBHf+6Oud1nPhDz8PiZsn4Pc9gHgCY/zHS4rHIwZmhHVSu4
t+qdQnkXYrqmfWs6iVdoKUGdITWTlqI7wyXBYQKHQv8eRfsehJcqhVrCW3Qu2rcl
+n0YZB89h1M3ixXsz32b6on8W/HsFNbzo/fgMdvSolGaUcXDAAed2K9g/hdC5D/z
gXTT2JG0yBbgl5TcE+ne5zfeYSDOTrtdE9kBKgB/9bPUzcmF2QpozTQWmT/tGKWj
mCUzdnafaaIWTvW9SG8TVorUnpDY9c0yZCNmLA39coAfKOSkcu9FcysrOQrIQn7J
kdJT1R7apvdnPHQBwJB4Og8OmeQhmW3T1i64d2kdZHBXx0w98XSLEp/QGA+5tbRR
gOxUjFdHCNJsc8n4UtRlRd5rKcsvI6Um3RSNjOSv9l42xk6uxXSf/d7C/DS9j8DZ
uzNQQ7rIonxZLNS/L3mPr4TWrNFdPrXPUWGOt+Z97/CNTCKcGJx6WUIYdENSihrk
TLM5mFOnhvky3OVRQnX0PDJgpWsUd2yPtt7uWCXMgiOqukMeTzWBTxuuOyNHRPd4
AceNgjwKNx3Yuasj9M/E3orM+LkjQte7qTSsFvssi2P7hH/NTilCsgFGaiDWlMWG
spBtJ80M0qodyoHIlktXEvUSQJbHPk//JL9wgkvKd0dva7Y24BFakLXeZ+oCMiUr
olVnDOJL2NPLPWxwwp3ySobUGrX/AzURgdZU8O2cmydSZjqzwyPTixl8HkVyEdgw
DJPe+hjpJEtKtnF32nAYnZCsKdLe3uekhhObak+OtUOX2/+O/Hwh03bsFRcfOlbW
S5U7LCfY20Dne1MsGaSrYiHsnpfdQzpFrNK/l/MNkje1+1WxpffMGPxbh4w3v+7q
fGIT+TRrNl26GH7+YDcISoOr62ZuOaBcfP2Y8og65xg2PEdSNKbmcOsmWKHqweyU
VTMItglBP/H04Xqiaykkx1Mpxoek/P92a1YMt/iMAA2WJtEy6gTTWnUpVCqf56s6
PFaNIWFgCP/1IFaJQnfE6qJkDv7oOiwkoVyrxqIhy2vuS6SAkmOBe3c7iKdMW3DL
aI8SXlJYTU3uoQUJBQaJai+O7TCzCYUc7n3WKNyc3WUBXVBxe3Sw7vvxQhkIVTyr
wasTmYzLv2SjMSLuTBAqefkAj8mvRsabnQIye/AKUGXIvsTewu3FEwbgKto0pBuF
d0yD/hlXivAZ9hkmFNx2XMFLhzIXc/x00iAbK4lEMCR5i0ToWwgO3KEyLgNnxMmU
VNsXBQ1FSDRptuGCxgebbG81DAYxD3WZKFhKVj02JK5NIKUtZDsJdBuCDHJFs4Yk
DNWQkYdOMTwY1LWkaelT/PKPHhthU9X8PW0QKx/ujccPRSFsAJdZVeb9vzb7Vzde
uC5KX9Smd2eqU4f/chUTfNZjGBH1OUvMDu4skDbJda9DA3hICMG7PTFiamLwgyOY
0dWYWJvKTXj+vR26KKV2AmSUHdpJ+x7Rs2a0XNshCfloDdLjJ8WdwJLd5byIkxcv
E14GP6614jLx4yZBxvu9LqXyuQJ6R/1XV5CXLOFo4NywCmw4RYbAO5p4vzK46dc0
Ge6+D4OiuQKJyOEXFyBpGnliztm0pSEXHogwTqhmR0obsyBwumOTPpWKRVQcyN+k
gy/PzIE1hljcCaTPbqij3Sl2ekPkpVLRS748Ug53FRcPn9YwOPT7TVsCgRBwxvkW
YZi5UVQSDW8oOfoxY7rgNeUclSg0/FD7uprnla1ccv9tTMumQ50gPEQr5MCeFqtl
oRLJuHhpsCDi+dgU/Fwtz71fwGwKwZunyBwyWb+DXyoz/KOKPiJYaNvnvy47f4fA
4zbwFfVxqEhKFmT2hFmcsLnoeBoQucicS9TdnLgfFreZYdIZganNil1bH7xKpsq6
jGgOz8R8EdLHt9FP/i27BWTC2UqRGJRBkmWt95+Jpg3CXFG8cNA7LCuzPUl02OJU
lYW89kdmoecqV+DX5dsAlItVg2tNFNTpCvHLjIuYAVZmROOQaLBqEO8mHelnSPhT
DKJ7KabQbMoqE2q9Yb6yfngaySD+xfAkvuVJVLzM77pv5IutxBX1inmVpUGa7Y7Y
qClbKZiA/PUaA3qZmVq4uQMgvGy766QQ6ro4G2CRgRlcgoT/5z0ojh27Jgh6Z4bo
l1UtS1V9KLFS5XsHQdBz4lrWaEg98AG7tCZ5ow54N6emXntFrFiDY8bbEgqejDHm
/OiB2Hevnyw6H4gQF/OvrlZDx2ajyYuHCnNLJNGrsb9DOqzWX0B6+idSmW6ZFP9t
7Z2anjC30ve3wvnc87hau+Wi6lgpjvSFno4ppfO18E66rJYQxDZU20UkSGpuiqrF
DrkZE4wPK+e3ZVgFQvvAKCLSXPlJdQ6BZ+N8UL8tFpgzVWM2qTGo7lvrSpXbO5qF
g8yT/EOcDk+3nyalCf7w0LPz1a1wLOrCKZANfW03vyivx2Onhag/BFtjy9HGQPuz
KQret142NXbyPojTA8cMXXFZGoiGZiak3BX+MrixtA5ty5Qh3kXnzhMTQjcPQsg4
D3BuoHUzV+5MpUAi/RlwwCgNeUGunE1mnxATP/uy88qQ9LfOnGzHocCKhKkJf+dz
pvAeGkSsLLgRjEQdIk0YIjzli1x7hUPcHC+fBnW30iNqBzMwN92YLT+TP+Iog0cE
168hD4hDIv49yhoFTrd6GsUaixP2UsmuyAs9ka97ExBcJAH3YPKx1VFzbwFJRI32
yhiNMrBYRxWSrHJvqKrXZF36CobcGVnY2N/z1esoE283HlxBJcTLlGDV0VqscC3i
EqfS4J7zNRvOo0lTMAm3l8p0i3Wsde2DV87v7dnd0PlDu7/PWHlXSQlmcIzSJvQx
+ID1QfKXt3l6F4+KxIV5FD085qdyksIioxAWEqgFrjEIYpah+lSAgNTWe4WBL/fw
N6tYrRV0u+Cy9nJTf+AYBwIFq4CdBJ8F8gII+IokpGK99E850/Pc+oIew3q7ndMP
XmnpEOtlxPxTflOtYlp+4Z+5EUC+JXcfEl3+zMKraUY9y4r6XHYBixzGwY5l7qF1
L4zmF4eT8fQIhelOyV/h7iXgGz1s6NdFGl3J2xUt8ak21HWZfUuzX1I93m/RzpjG
rXYFd389GnfobyzFuwuaXqMdiooKc3+t49ir28NrEPr23s00P/oFqd+FhJO1GMYR
2My+tzP9rEQxNZ/V9uj7DIAAvfU/4gqA1JMShsMDrmGOaNtNxdn0J1dpwLpWXY0r
658rX1Zr1kUOD3m8awYZka0dCXxSCnTkxiUg3sVsgs4Mqk6lK1zsANSlICLtYCyu
IuTFjotqaZQWyNyRllvhZ8zDet1O08YesLe0uICrJL7uaxpZWfVQcie2//IcEVTv
AGPxn4PKxr3c90ZCPST6WccUreqW9gYVyJVd5rKdWJj4k9/yRmIOyxJfC55BaqA7
nRYF0C7W6E3fmgfjgAjXYpU0VxqvuFVDX3jcTbCIgb3qDnO9TccXNFRGHIs6lqwv
JFbmYIDjTBQocFJPsJoJcfN1cpx31xsE4Vt6JZeBnfrju6u+Sn/IfhMhLoLCpElZ
JL5dadujGhMlPb4FBATPzWztHWtzXcboyLHDP2MmvoqPQkn8+1zcrkNKwMs/Y6pp
/nx2NxvWdK/a6lsfjZu10bQCyuGJv3bKRGBBL2C/+C2Ln0xXKhysgXp/JlyTOYPz
n1cCvRYtygOhd2S+HlzPCrVnqz0nH6rh6i8hk6g3ILZYBeK1KookrV4OqsidahK5
FseIlA+p+jUt0Ff/3a057jBekqo/nkcabg5FlBGa2rO+jXf8nCQj2ynsi9wHTBxD
j3YXRQCAHDvrk0aQ4D2n8AjBRI/KTuHua6FtOKoUXm/0ijbj6Je5CRjXN7t2bR4g
Q7CdKA4fs7GoWXGLV4CUVU88nrJ6kvjNWVqiOHKWTiBppqPiC1xye0y+jk5wypU5
dsE9T8Dx2dXK6ZmZasMJ5f8XNORvjVmzPsNO5t1JfR8HsbA4T+RNiWEU1LSWtHWV
LVwugbF/1as5imnLER57noyV/7gqDH74tr72b1GURnnVyYDG9wIuNO1ZTZvOTuNR
ogSeJNaQ58m8iMEkr2HIAQhAVNZtwvKHu/vhFb6dzsI7M8JvuXP/uk0wTqtJGt9G
QmVABNKxT2IHcNTxX6jdlvgTEnRUn0Y6DdV8XUyy9FzkG08htkVxr7xD4HuOJCED
Eye43gW4LFmawTW7D83clX3oDuOAxi7SFPupG7FVWGftfNHzcGPVwuNnZhS2aoCG
yYb5uUR7TF8N17GElWfOe+kNmtsb5HjnZpPQssccBtyIy/ioL7Byt6XL5mqH3OW7
Z6LnejlOaocqeuj2CHpLm/xk8wbTiBsJVYmvI07ValhlJMdoFGQCCOTqlhUUS9kb
ln+AREiMLvt98aJbZyQsD4Hx/OywUuJ2cRTC26ZPSTLDAVH7M1ondXx73IPR00f0
mn21IH2Velh27QjUtlIG+0TOWbjhjvQBOVQ0KyUXZPjxKhnPMp8dfobdeFv/7kmK
iEBEQUzVYfmkcPlNr+KfYKmp4UH30ylie9Dl6KGeJpI394xRY8JMj286QwA7HbAe
Hd8+yaj9J9uSYbD4CNehoogaSdb2sS5eL8RBg66zfAcbzGTPjuht0jLfuJur91PV
eY/Jz1m73uXIDlWSCK8sN8joBNvvHqfgWWpjwf5l6S9x43UgzEvV8PrjOtHtjz7Q
0b6MMkTn5/rgwXAgNoqVkixw/FOvzZwDdG4mMNndn4TZbexzh5ThX5xn5+e4VZqj
/PFWLeiUkxk3rogOR/elbG/T+qt6S+4mlr805F5DIugq3pWcVuSD+me0bKKLAsaS
G19Luu3LJW+t7WYfldjwOhWBNfwHTZxd8+65mBz4x0kGMsl4nBDIFsvkvrbD9zQb
yo4SKpC15zj0l2GN2BV8VBx116C/hQBrHi9WxfbCU0gE0ZlUSdVvonb6cg6Cw8/B
qez9u+cPgrt5Ikjvq6dQ1okb3a2UcXmwOF2BYlMKQMiar2Sqc9k86qex4pQ96Kvy
jnKS+pHp4FnIxAlsUGHrzSj3lROpH/vV0u/mdoNnbczTBAYYatRtvVYIMpdnS88b
XU06molaWMR3aeCN9LsARhib/PNIJN+24pX10jjvZDEJKXKxLqWTRhlTmktnioNr
KvfYUPXEN2mr2NxRYa6DAVtMvOSXlmTVT3Vw3R/RUrX6ViRa6tyCvZgqPPDMG4Ir
oMf3nDWbqJCbFhYH5RMU8w6j8xvchAdseeUwbQCCL4iDTT9+03P+auupQCY5uwi3
ndRrRJ1WE/R3/nWdnj1SDqymvRHoiawiPJZLV0cuWJ9ItU3fSsaul+PoXQSdIWFg
A9X84nxLh4zSkVcNsSsJTJQa1F7gUBpajfgQIvg5HNN9Jklk7GEQDcPQZVRnW4oE
oFO8yWJ70/iezgITe/lQf/meJus5rv5GOqN6tpQyOkknrozFJ3Yma9IppWzwz6jS
ASm5KJISdg5Jsi3p7wUum+Wh0B4v/4bS+6HM2JOyB7CXCbN9RiAt4DK6o9dPSxvS
3DqE40A8OfZjpUnPiLqBq6Ja+xut3H2Beb+xE5mw4ZB9dxQGlTFbKllQVupmCHwR
8qA4yLgfETzLly14kRtxvaCWjJicRndrpP+uFBD/Y/+BGYJjBsAN2kgimCGuY7fX
sNjK/UkxQal2tX1AbLMH1ofYFBAQMJxDH/84N3aOlfDoBHkE9vQ90uSdE1X2Ds/6
dU35u3mx2DN89dACei3vLCxHR445F5IxtzzhUYeCp2a1VLn7MB30Ie9AplEg+S8O
ysG3wPLWuk0RJOUjAy6FaipasjmbmbOSLIofF8q+N2WxPEgMwHogldPxCbBZuSlT
gbVL0E27qcZhvQjMvLMhj1iCTVgAcnQ6Cv9QrWJv2+0HjSuz2TAp2iGLJiZN7/3O
54Ek+NEk7ClNoIX2w/lovew0/jqjTxHpy578DeKXjXLCCLPVFj1ibgA+DkeS/lad
J10ziOBicClerofgoY6PGNVLq3duQyi6HdaLG5GKYIqOYCw6TPrpJ5fTz7KUe+qm
OwE1oGpN5+5aM77dfU5WCPCHBEFch9bq+S+w1r3aVSgBQSOY3l7QY4kStcLH977r
VGAGk580/dAhd96M24kf1lHV25FX1hJgKdwCVKs19HTZy5mHb0qRM33gNtVAXoXv
/xaX1wh7Cv5HNg/473tdY5wBS0tDXG5RpF/RU0qJSjUP/i3M4SUioXnSHhf7eNCz
ZGm2uqIoRmjVYgGL5lW7eLf3Tgfjz+F4RXkQPUnsn6BfUsxjM1Z5a6+Vzm0gJkqo
m/Cj44rOZFddmFqyYHX4Z+Lz6JmT8/nyETTYjfJOoGwU0R7P2/M+zcdVRXuu+5SQ
PHZOPOB3biHppwObz4ng4EU+2eLavO3pDhNUmkc0Abjrm+x5Nr6nAqJDmFeU49Fu
ywjtW9BnZCxSYRBaey8UR1iyUbS5ZSTNCHDsICHSwQ+ZKSvNKU9+tzBjNckXX7eO
n9IDJOLid5zQf9X6SngcgnM+VjFziWpycjNnbEvZeyDtt+9EacYjmpHJr86TbzS7
AiVve4G1q2o4ffQCrDltG2Z1rQFUd0rfwGfheX8QXwjb83RAGcBWRq5/Ead7ZjV5
6DLlUBFlJSozkCtQVL1PQpXQItbmrXMdxGq4tcEl+9Rf7wRA7A3OdRlNhCEICvP/
cfAsPgs8FOOt7y5nKNvpyNQ3o6DhXDA0rPRFDqloZN8zTH0zIxyA5gKjzNqP8LeU
IIgm3zpDIvvSJxGVvb4/EPwDPIBAq87eHBPv8VeTYPtn3/e3uMT895c2MdjkR3/V
eEem5wMdBKrZ7hCUYhXnjzgIwQ9FX9yBXCQrZHB5/IFgWm9mRo+pVOt7Dl4XwTae
yZTJ7/WjiZWnWJ2uuSZKNZKYcwRLPg/+S3qdb5u17c/ZCYn4ECbv3Usz/mv/3Val
xac9SavzDODj+NzTtb3afpnP712g6H3VerUHArrUbOSwNyJ91M21rcn3+qXdEkLI
9Pmmtcf1yhgdgIFrDTNsfIGjimAAOia2N+0kgTKBPmWN7/1d33iI4vXQshoNVcOl
Dpow4jE9/aCultkM94Hbh/L33IpgV6FzT1DViqMTNoTYvj2VMKVMdiGzhwM1n+8d
IztKXDbKlN/KVtXr20CYY0KoadxPobtFxVkTPlQHjZ6xpsuqJaPU20MIpBdsyMBJ
o3RYIdXmXzKE56TSDii9QUJ5Mop6soPe2c3TvxVCARfwEX44BpVV8a8ZH7oYbUdD
tH6ClNcwuAXUF/21FQxZ32qwFMQKyB54c5iNn/Z5+TZbkgkUaYD1G5eger1SlXPN
dkBnMZU1Ct/8kXuXWBP2atwITkivyNll+O4tnQ5Ss/wLux71GDfXYD3+hit9LMfA
VFEGjj2hh0gOFlW4giuv+1IVXraJLOFbrL3sp4w4NzU/VQfgiJAZBtstq/uLiiIj
mWeNK2v3XTV773nSuLO4m0t+WEtZo/nipwsmt6rK0Lu/f4Ad4tLBGaDyzFWGtBBl
kNPi7d6+CyWZlWgEj5xqV4n4pNxrzx6VxF+kXtr3eni9IJ6NFVozlcNhHiqxotgt
NIHsvjtg1cgrmpmpPWm6BVenZlicZwpmkkUsB3OU7IoedYTWJWFxpF+RmPZZftm4
vJcpOoxE3IDoLfSv1pLgIewdMSDrpGtnwgqMObHMhZ7OWSA/fKL7U2PIsH9dLB/v
f54mtlEodMyHbbqIhTD7scHgj3lhwQno5CSOV/Sbl4GJCs9p6m5nvayZ2KThs66a
LzuMJjN9oE1P4p3rlvKD6NvBNpIJontYBV4kMR4mKDCNxKxpt0JVSvWwfI5bw8hU
/GGYX+xHUsKEXKnWR++W7hjZH/CPz5l2mZx490gJX54ZPbTb1ip9NEqq3oPYt3zd
+bQVPSjCrsyO/zT+AWzoAo4T01hIGmbt20ySywiffoPG0Qi+D8ncy2Afly0RA60B
YDKFMCfzaK1Qo0Wr+T1gxIRXV0Ba2Fon6OMBftgifUOlmdVh+sG1Dpx5Q8F/zY4s
LsbsaF6dDmCT3JM1xoxUf1eDAXNZ3ty2ytzCIp5ATDVGc2U3SrCvWb264rQIp41T
RbvkIg8aWHNLWhKc5l2SQMuq14MvsYHYPNY0flleWnPOwO0uuh8gFJI+kLLO5vo4
VTaQmw+ndnLiQQHxX2LklVE3QAb/gbBIgaY0bRvQjtyCW141Zc/UplTBQF1E5EmU
LJsVnEmeQl8xIsqBa3I2fbG2rdKn7OJRglBQFyk2THY5G5ZEiOBLN5oUT1oplTxJ
chkBSO7kSOcVI5xRZ97ihmoqggaDruwrHkT2R/0dMZ7ZOCh5TncA3CSmmHeQ5U7R
HnaYyty6aOMFjPMbVviiwmTebdROHX1EOM51GNUFHz5FzkK6ZiYzg+dafkG6PWpZ
x5M48SaTLmf5g/F5BwfCfQYOGgQpqP07R8hvrvaopPOsxcjw/Xoo55hFKckyRZai
skva+00ySOXAZAOpunCoJkNhXyKzELVHBTNGE1nl/okCNcxSngy+qqyVp/gx+P26
9yAsijj2ZTI4iepFUGoidI0JFX16FW62mmQzpKvt/R7CX9I0knk4U/tLQjxd4R0f
36Zn/jY3Pv+IJi6EsdDGQO2Ol7KOSREXih07hF/aBH78bw/Vio1CK+wJzqsu+FmE
v6746g25j05Xu8LTs20MbYw9/gTXFs2OGpcvNGpm3a3rI/UiH7N8lE4c3smF+gar
dYN7sZCKPDzoH/JMhRNtk8ikUnq3+hIznB9F6ihXjlVqQa6g6bG6gjr7jznrzAC3
xRPU2XaR/IiYPpLq+deuh4inPMHdHYShiMOAYWH+XEmWfF5gNITykqb+0SYJOmVs
fwxLjGyEBie7VL3wj5MxlrZ0YnXo7vKInACO4odXkJvYJb4UGC1vslfQurQG8FEQ
kcCQI6RYCXr80pk3/7eOaAnrkt0bDN9nL6uoDCvB8QPQhtb0npkga3vO2L9k2v+Y
8LRTAcYzPPfoXhu/n3LHX6LKfAvDJH+VJm7d+4ue78WyBuc8mcP44qsKxC3eXWl1
AknY/vdm904i6HRSTEo5P6dReq61yqQmv0+woPWKh5V3GTHC1zNYdCw8M/sLR4Lj
apHbBKrIMZEDcroJlH2dNzOyg7XQ2tYikIihtsRQsZk9j7w77AHQUhVD3DcE1JNk
r7olXTvfXP39C/0JvxZIBxTQJ6peeMdxPcvU1Gb3+WZNJpuhRVxOMaypUvgsiA/v
G4vWNgV1bpzsM1SvtePY3pWEeu9GpG4AUJy1/Ec6hf3HAOnzF0GFGDnlve56nEMe
eXMrXmmiIefOnQU7LvcLoAoHsWeXb56bUlsk9Fi1wg1zNsYz1Jvnq14+vbBqFFGo
CG7F3J1TEwePcu534gjeHr/6FYuLRaeoreHld8iOHB1tWtdbRHlswJs/YZoKgHJ0
sZgjcVU0RLoDMhnihKKjAIPgbRd4mZu6rDv8ddyU2RdtfOgshgmyg1W+ddNq6LTT
lCLuMPpTOczikvr93zzzU+BKbGY3XUq4r9Vn/MAxYVPYSQZVbRs8aoEhDnmVQ4As
49kpPcrZxSW/ajpzJZXlD4rp25dqfU29X8w7gckJ5q7p1Ks2uC5BusD0M5M/XYJ6
EYIzIy+/t7frp7Kr48xwCcxRfiB5Czq0WMTcElCBLxEDLX/LnCcjwrODZ7gP2gBb
R6gi+PsUojsNAkd8xQAI0hv8gse7B836tDKlbZDoIQ5HBIp8TRnD6iSGjdtRxDli
Zw0E4BfoU1MAWFxQe8++WFb8ikrN+K8PUIRIWgziFMdn+x9gRfIm+dHh/Zom5821
IYIZDj8ol8QBCOh0aamhO99NlHA7xxqfI91w2o4lHnGvl5NOwNRGUnLATKt5un1w
L19t4F39JsFUWwvZcgjfhjawDUzd0hIGyb9MUO+IhK5CDwg0LRqb3Qzrrsjn8xO0
GcsbayOlhES43sa3+DMZsNxJWN2/xBTayI5h3qTY12nw5Z5oC8xx1glPfFtaTzyD
zQn9qcxQM7MQt+XtjOPBwFvEJyshQlwp+D1sYqKe6Fe3oMY/m8fKP7cd1kRZ6YpN
PuCL1nzPaZBBdh5MLA3Z/XF6crCodNPHErIVGJlGZzMASPrJlqD45yaFwDJYo1hQ
i0ITHo4v+zxmQtgCXtkwDaP6UakhVuzilTpOBYBrBr4M7JGAHLvodmHMWvNNa788
wr1nhNpC3WFBMEICp8SPUHQJm9uQKxdCKeUrXXdK58sdbFhrN/nzP9UFdRr0IJsM
mi08O4XzW4hRfm0SfKGxjFmHdRu3GwgtB3+i3zSLXYtaAd1E4hAXnx7JSutn/jl5
V66dPEh5Pp/Qlc2XzLhHLmpTSDgS/aHLCXMl9GFpSQxoXwKAx4nzFE0Kn97dIgKi
ldcMnBmoizdi2w3JL1FNLpTxtu6+fFHj5t+S9Oafq0AEob0/yhcjBuhsbqWtFxiw
tCJZC+mEBxO/f4/IIocWtSwXOAlT0jZYELVtKgj0czyejZKvH0iYD9mdyjOTkA9o
99a/e0/pDoRH5tdUmPfhK1rhCKAMB2WKjEK6ketcqgL0oheadqajUny6oBN7H2N5
KKSzCJusD6/v2fA4IOTSyBGEnNeMC/d4PwFXWjOryxcwbgeDBYLrBsJq75dTmmjj
h2QGE2gVg1m8X22Yc5LoTP5V4WP8tLv3CV8V/dW9KtgvT7L2LiRSUyG2iP6WyDIe
VeydYK2GObFNMZWnnkYG0jvOjzfs/lsQaKL3E+Ngq6y70HpZTzMNGEhb1t1D14YS
Zb8yl0DFkzJF04jcbbe2wzLBHUf5rDlUZCUWs07YQWBP2CpZrgiPoypc7raYJdQV
VpXWc2s9Pvegg+YZ1WPhaTu/MpKvNsSaSuM2w1Tcm/BixQ6Lop1FIAJSlhUDNn1f
bBOy8tgAXJIWxFhaLUDkYeVmGd4gG9+jDueDwWeWoHLQmrL/lWDQbU2BgZyq0Clh
g19n1xUyn7x5Lcs02yPRcrlBFJO2mI7P/kdvdYcV1Ho0DbtNF0ePZtI+fFlHHItH
/lIkMNg1AjIj0b3+jOHmkqONjHFmk2BXkpsalCAXZYfyoHfcRSePQ69zMzsJsA8a
MfEdxnIZiYCSN0K9tKJKZ3rVVrZfj42Pb06PYfyAavrJ4UOT/RKntqrfuz9n7aSb
OnKLbykzpsbH5utuMvUXE7QMWemP8f1CXw04TW+SwCCoqjdUSlUb2rdja88BrqzR
/EbRWfMrcP2R+ACYiDxNNwSUVlJ6r4BtEWCo8Uq86O2WTtIow+HQmxjfu0wrTHuZ
+IN6wM7rklq3/9yTnm5bQL8gjNxWYosGrCr/77is2cVCZtDmDj7j4043TQ2/KEmZ
Xg91eqkWyNLCD2UBYYKBcihSKit6L9L27yJDj70kv74A//Hih8w6FfmeFJyM53yw
ZZYJtboFK/B9hYIIbvI/x5M8QJPUVMhVvecBdr4lVpBvlNqq9kBzuyzop5BZqacq
Y3ARulabokZ2X48fk/Wu1nX6GC1HC9+wAPqg5zkZZYqSC+GmhxQ0Zj6noum9g8rB
5tCCobyvYVQI75tUW4a4+c+UxYmt8tk0zPvoBYWjFiVKaI1knLSsYM2F35bUjq8+
y12ouz5RG4x/F82Bp1oXnzAc0MYpWMixaLGVcgxnhOX0Lml8M/elPpzInlc3dnzg
K9XyYCItH/mkfTK+GvkRJuy+192IHRan0+0JhAcGaEMpL1/ZEaqVkwjv9KWtAuLj
M/IzCOUALaITTQMTGtAUKnUi78fyOvg8iCLaHDq+1nnidJa2/+fST16G/3rpd/tT
5CzsgLJ5flPszMTtmk7eSuoRv4+NTBmdxCaGY3IMo2VovMwHK8WevPlfUgmyYdKW
wk6Yi9NFefG6sSeY0bhNaxUySK3oWJcqrSk0ksk2wGgOYYM7oe8nzOpYJ822Vhc7
muBOGRuWhN8d1GwYzwwskxlsLNLAMLoNrAxTHAP+aWfdxasK778UPZ+nFDw13iOd
PUCtWYLCh8RlwgEpAOFSH6BFOFq/Q9zvHbT8rJsDi6aLH/Er2IsvKcL0JXQ6NLES
tl1TUsFUS3XrDboDImCXcIUFOjESiDyktzpy5nSmt/SdlOZugXbKjDJKXIsPLY8U
7RvksYXJWIPpPAzEMd1K+8Z6B/zPdVdicp4vPsWcYAZeSEpiixlmFgLUpLBmmmY1
Xv2RH2Q5MlaZAGfpViweE9XX2l8ZUUyWsWWR5R1cV+T2JMHLa7+RiclypZ+7MI8a
GifeQyOpOeB/UakD+d0ZxWBpDisHr2hj9os+SD4ZVswIqg6wCHAuX8GG0eoOJ+Bg
6S2x8KkerWbdGEWmdCItk03m6Q/q3uXnw5s7ZjWJkjCePMXUT21RgDuHADi2FfoL
I/m3pq0W6v9prwn6qoICweO12uvUFTxlCetZPLW1xraanpkbCcV2OYZHuk7ukKLu
6nYtClEHfuJsUzf3BL8fGPBWCoW6MPUEzQ+r6Dz1kkrVwzh3Of3Y6i5XpRLivV91
5TuHADx6w9Eb1reJ4Cz/4lUbzmgrVdLh5hE4Kzpbd0zim8WNO2nIoy1+qdOntAaq
oRXE4Vd4aChgDnTN0Sx5SGy3EGO3enTzQNBHEKQYaJsnjN/8x/gtBvnL5lB5UEMG
Lw/TNs1Z91s2CUFDjruOpo+jxNSs9wAfRpccD3HpTo4Dct0EcsW7E8W1oV2jA9ul
EZsbmiw663C85FBgUH5pTeMgX0L9MrWyp/+f7O0PoMdxoZ6ZKE91SVP7dPEY4tYW
yoKTPLNhRU13aRQOlVZ4EMPgci3eLCdrDQPvy7EC2WUKB45tyX3T44t3B1PW2LRI
0iamxzy0lAom21cr2VdbAcKApQfYGhnITGW3JWIn+tx5ewagcxHQRyPzrqAg+4Yl
Ki1FfVugJIygJqkrTsM/1eSXUw67Vg9m51Wqh1ghzmQ4+dF05Ew2le5iZAtI3pzq
jYLdpXsApHjC4b8WaAACEIAFYR1NQfmrQvGgFDC8V7+Sgu7YlG/0+vALdOwt7stu
73EqdzFEi1zM5NHVTJP6NSjz61yCvViWo68q/1UHsm3+jV+Sh7pvQ+vX0eO+tBKZ
kj1Oi5eCeMNsae9kMLd7KSRiODCPxUgT+Nlblcu/o/hu7CPfBx2/qQtE8K24jq9v
7FHHEkwdawb6wB+8+bUNQVQiaF2pFJRBzgKUmw4khHamj9ui+fs+qHfV4Fo0xm7Y
1huflEiDPB/BJCEs0cOibM2v5sZUWuoURLAWLD+l7rfFJzP0ge2fg8tHQ+mHt9JK
IveaBfC0sOsB227OuzxsWk9/VwEks6BtZQ0++qqWPSLhY+k2+L4TMF6QyxH9P25k
UfjF4chmQaiczlVq2GekUYLXoyZsvgB+lfpfJaicRTWRYXewBR55IrDR+V6ZNSrY
ZZY2wp1LxqXtQug/2vkUXoFRIeZKbrJX4UqXyXn5ggdb+CEf84mqWzFU6y48RCAp
OUlCMP/lWp6GwLhHL2+2KbX/i6uOhvjuT7bWAgDlyQJLbbFVvotHWQgqJ4srH6VZ
hukIFZD/lfe2xpd7obyl9N+LVnxjY6THy+oM25T2SojWE7vjGtVOjeeT3EJ1qLdd
b+el9r46iSoRNQFuHcV/PYKOVuo7c2VgcLQ1qk9HgGvrP2NC0srd5HDPMdHnjo+8
xG9GgD6heUh5eobd/qvn63qJQXGXwsUQRa/3ToTRtdzAriLDkj6uwLDm6v1NWDxS
ZYvQ5PGfinzdHghyhaY2olfUNw2PZ0TY8YQGSKwhqPfM3tgNYzFFMcCiKrFfsols
OSBj4CSAi6d7u9I6kjAsCEUEAWBtQK07fxUstOAOgCROxLzH3UEniSujmmpeAbLv
7ZsxIfoB5YXjEuvQ6QcEEO1WNXa7fbBCxYJdDKK0ZsEA4ffHHuJZCTYzGdJBBw0t
Z/KGi6iVLwsn9rSaLSXsyrhFr/1wZyVKppDbw5fqWk1LmyvY1lsWgSrybR+rH4AF
LrlVy/e+pPg9M5cxRqBH+yKREgGEdYVyHeOWmWkYGHXzGbusK/Es0/pVCmoU8l1x
dsQJXbU1z13BIepwh0lp+TsTOCaL8O3WgdR6n8gxZ0mpfbxEBFLX/ANfiCCI6o8+
aarEamvcy3kr8SZhU456EZ5kX6WwuDDxQ0mpuNdjk2V+hUMHjFcOPEojRM2Krq3L
7JKRwp3iQKVvvDQEqTHLfi9seCaNglrl6gPn1g8JDRhUJGs8YfaDotf6jQyL8T++
C125+hbZKaNlSmmj2iBkZVRVS7FNFoBR79yMkk/1DxtSbMRZEwc3XH1cpR553gnx
IzIio3bQIlFhClwVGmEExRoeCazLtpcYX4hsnMu/o04XOA4EfvnT27wQUhSHlZJ/
YmnuWM2SOt9+4OscnQgu55KtSFRH//oylXCQM2gDBAGHuoW2IOHuevHxfz1mh3PI
j0+SnIq3UQrJ8vqhVBvWRvurs4q90GAO57G8FNhBYPNWETxqxwIyWPVT+dtkefWw
Q7Xz3MxQFF5nWRyOUKVj4K+adoH0q6UuKgQWM53svqvGSjndPgReM14Lj6doY0tw
vEGxL6IiE1cgXxXW47wG+Dbd8AoJtAAUDW0MJ2ZgGD+OD/13lM54TGfppOWiZ0gQ
kXgz9mcHDNH0iVdlgg++3u+6ji2EomkSgNiRGSrzEgLKLYdp9uye/CvMx7EeM6aF
fycWCKg4M1SI2r2SSwnBYVOuK1YndUpE4OP3LNV0lBScgIIF2OfFvkFwiJzPbpOq
JG0CCex/zXRkiPi0ZS0Jcjn3/Rn/uIRM3w6Wr9FO5o2Vh3MIMi/sQXo2DKvGgpBp
+hHRMdB43ht6F8hCRmEof4DLEM9ldZklMcRml7v6nYwJ6sWej4sRrWd9c8pOTHWa
gppfSyidAwqwPcDFMpq1O9PDd3uo6i1P9Dh4CDU3ExlNG3da9OQ6o8YZIAe1RuDx
PQnr21d2geKPPA9BOpIJ280uV+3t6JNcyMKUdIDAICM42cNMOKbm4TjQsdTYUKxy
twErJeIWeyelZ6zHb+NGtX0OLhYgYCpdk0CcLfzx43lboDHq0y/eTT1sh5yfYgoc
MbEl+T4eqGAn+sNe1pIOMxWPRZXLy48Pm7eKnjL/YXsaR8O5rzDdd6YW7sgTkBJ2
9lWegG9TBgXGiXVV+xB9epum1JE5d2mBtCc9cO48q1z9HsAOdp9vUyudkn8TpPm9
4JpWhCb45oEdAzjT451R3Ukp6BhntaKXGABD+tnuNBRKbuZZ80rjmAgwZ0JXJo0A
QpcT5EGF5Bqous0r1Rx6sxYbmUAYD9/yz1WRKIjovVMZFpgACphv8FKYtoOrQ4O1
OivqxL3L810GTNFncfOdatbgWastIC2TT9DGRob6pzjVxQQ0/eNK2jYW+b9ZIDeI
xv5m2gYDnZ7EMdKFC3g9AVJrzu2JE6ugy/K2erAHYWptsQjN90vuBJK6hwgIP+ax
Coyo5b2e68GWNiRQDi2tjLnbUftXaYo2XWIQUhLKPVLhJDUG3totYdk23Sa5y44c
cKwONnhC3A1oWj/kVna/+Qi1KCE8M1XGOW5oRi/efVFZIsCkH2kjgTnULSD5dMt7
iQ8+b4uOetp2GcKGxzTHtFLDgwE3iOn4+00XMu/elD+CxnGphEPcyQemQw65ambo
s3DuXej0N1vhh4W0VmvgMCYFgKDeHApfVNgix4vMRuCoSipVqJDP279ZADX4MPZ2
wfGvrem07akTk3CULaAFPINnbaF9yOGexP0woDPPMVSE+prvhzzwifCgzuAVb8eD
qJNnAg54CKWkkAXcHrTdMfF8XZhn40JmZv4PQrGAP6fEVLAxcD8Em0nMTxRWV7fz
DWl+rxfX9z0tMeDA9B9avbLXHLcOQAXy8clwALQ2AI7dBdPeBkNCo07v5x2bJW7I
GfGzMAsxBLlpOkgWgA72eN4GYwVU76Hw6b4gNEHVJ4L795FgkAO7xRKDngphn5HS
HVBYa7tsDQKsWmTyz+2Ku/VpwCjrKJv+v9dPi5uS8NP3h/Brzd0offzojRRtgr1r
x6Ud0DvEjmSXZVEvX8bdcWwgjlLX4kOA1CvjIH9RTKVZwnF9NLy4xpESL5i/2NER
WhYYsJ+wHonG5FY3X7/3fbf/1T3OQ4XZvkQwETJOFRBmVcDCn+f8lK0VcSvtLRUk
FJ4uguKA0tbiv+zkwUzxAGLwbbakNWHIIUOG9BHGtl7gzHBb5p6Gi9tJIqisnjjf
ZMMfsPdZ/SugLeu4chpaFhbrVFe+0oPP8yUsDHNfqzwH5CukuuFeIgEly9LkMCBn
aNJMNo1xqLqwBZ5EefFz6H1M+5tcikYl44Z8wgpMSao/RvbN8BCNzPgbQKpoOoX6
M3eHjIJntadYGU0cCDC4a6AK9JPmPIKb77h+8/hJoTp+jEQRFHSogFBDXgJTGTXD
7V0nEFBgHoKql/IHUIROVapNTgXQ5GCfArPfB2bUT/1IZaosRJoJowC3FhFqDW3K
RwhHxMjSN0u41r53weWFGqjj8dlNrRo2K7WnEcbAJDGuck0V7wCcw1MJOqCNnl4q
Z9D6AEiTS0DsUfGzROD1JQGrCYtuOAl+BGVRh4djhHIk8lFG/svdaqBVN5uOXcfT
b5xuHdK/5fuuQDRvas10pfs+u8K2JrPkKslnftEH7Yk7u5o4aTH/KKfwxk3mhegT
lmUgb+dtzK3nsOL/SFflgP+Y+bkCT6vDY81BoBFCI4iw1MbIXhZoYADHdFrGzBnF
iD7uO25ZAGYYXD5kVP9qZe9rxGXbhEwvjiLlNx+b6dMAMrYLbE4DrDRaR3RU/x1K
uT+5AwZQ78Z5KQc8aFzCT293keM/G0dMvhp98VrsmazHyQO9Uem7DVX8kOdP5+/X
iQndqlzOqADDtuEjALTlKZDNJYuDkCItThMtvWNyvSsY+d8kN3uIT+ZjyBY1f+Oi
A7CbszxEGP/W8z7vd1cfJwLtLHCB6b7vAuOKoIxr/ghhroNzNXjk+pawNNA8SDsc
dH1tFSZjZdIjZs0WPW7P5x6go3yrZrLZ89tNRq0tQJRzdM2iOPVyn9mrL4K9mi2J
Irbi8v+V8jKZZ8fcqMbiSINSju9ZYh88ofUiejn+4pxauqd7mVAZG4vbQm63vbzm
cFUHR/GA9Qpy9NZ9gSVUov1A511DrIpa0ey6u6sXFuo6LxZo8CHcXHJK3MaFh0w5
87O6QCYmXlHjdJrHZL7aJ4j/jk/83UOJR0EMdR48vdSjl24xE0zM1Xvf/nznB6Ry
3V23m4nsCR8RtxhFuKgE5hi9LXM8sk20QEYuGvYUbBK+Nx2cEqAC1/HiNv9cE5xC
AiRGcCn3pqyFoT5J5qhYUduBI7feo0tstRMrl/7kbmcJIk+K9a47QTlfkNLIoUAO
CLG0SERvraZXMIIe7IJSpJwyHBtErgdiO9AlUuvGO5pJGkzWVVeG5WUV53kQfUxZ
Zv7tG47BzmBBrqPa7NiB3gO2gca8/wfre7wC/cQgycLczFBQiEfQxjIFHBMfcb5h
G3w9HU4pyoidn6EC+tiVKkdscokOeZLRYXRJhDAU4I96Hpc40g687fkfYMj6Cas/
tWaF8pAaw9bYE5P2YBQGpgWMRfhBZmOUs/ANQvaNLR2Sy1cO2Cy9nXR+15f/49tX
MXYX4ksOGKU8i0No9VZyJdAZAAXPWQVjMEiFS8sbaLdl5ihm0Ra6gTwvygq91Tzi
3c3PuGtkjHp5HIpxUarDrIeotm8+UYgHuS72lLWYKQFXCDbOJJIoKmbGDEVcUZGs
bMIr+8BbyMy8+Oa8IvSD6510WNq1RYr+OS+M3pWHrhnvVW9pGri5IcJXnpFeftnq
OKP8KvViULzGtk6dktvPUo2s4czeOXjP8nJiyrp4cCdNQWwU9fIPBQWiEYAVrGZS
h4B8kCpAmvHOko/RlAsxV2g/ihrCF7H6VIhLaluTc1C8H8UU3lsc0A85bOLqOUF+
6DmvLG5KNVKXjByMpM4awxMHe8NCQiZtAtaZ2khAkYdpeyHZOYbcK19aP7EUEFZS
mAJMZtD9ccEZSDtJvfq/q09LJd4Alf9B/CDy9zcgxys5uVR5e6Dw6GTdHDsLqLc3
4eCVGdUch9d82brhkv9qOCuZHLMKJcmURopEmthTXXrXDWrcGuQS69Yx0+RJwXMk
OtyU5xmYQWBjsnRLJaFNk6xGBRCXVS7T1LNbkhLD/KeD0X9Ki/n5+rEcV5IJGVe9
f3kWujuGd/fr24ydsmylOLlmeFIi3DZEOj/9FQXOWR7WSIjpatA3eiiwjScQ7Mco
M3vm6YZvY0kHvN8kSpEooPb3IrzlHQedv4yZYjPwELpbFkHNFN7Tw7ef8e8BePJX
X2slEfNLL7X1Rtowd2QzSMhD3An+t4PKmW71lNxv1DBMI+LDF/rpIXw68vkU/7JM
p8J6OVnSsy54c/rsCMmm9wEWGwxxVAQXsy1zU94QFw1kJJO/Vb9LQ1o0AkAxFOkD
s28h9udZ5RFiuOkOb5FuktuQxZkO9d1Lz7KJwn9nMBSbnUDZxNdbE/zl0411ZdNw
5bUFd5KDP2JUMgZTIuQY96yfuR9vCUKFShzbWi+JEgFlX1XUQJ9Kf/dPXW3myp9Q
jm5Ep1VfopHRYzgj9roZShSfO96U9FLe6Xem4GxNUsWp9/keQAkjvY8c5pRm+iF+
8fk4xuk/c5FioU+17EFKSpQJ35hdC47DAhE5xsCR8AS0obo17B/sd0N/beahquvf
Qvx7Pway5gXS6IdAIFI4R1MwmnBUNGWdfJu1z7TeWVoriYJ8knZlgV7KePqQoFnp
zBVmaBpEPnOEYuWyt+o2LS6RIst+O+baC8q4kE3i1iJvSMABRxNUgXO1zGnvsVxg
zgqCLabI9vcumBMLrLYqhEnTg/Ht2ydtc5yDVqHzmI12NZZpPjp82zf7WGHjRTkR
BJhL21svu/szqmkYJAuqFe4r5QalR8qGn6DheJ1YOiaMi60Ew3JGbNxlfXdjcVjJ
yAbuA4r6XfCS0d58yFpZ9w/YnOxjxBiZkA32+xYfZGSmCV2dN7ZXWANdDy5P7zdj
q9IJSBBM5cOEKOHE9V7HmdEoCYcXPURHOoSzW56SoeudFttgI99r2qE7osNh2pdM
WDvtLfXhRwLeRFRk/9nTxuVxHAmpFID+CxZ3NA7h2vhf4f0i+zmlL2H299+kC+PS
jVGUWNJmKd9haTHjmWeJJNGmcJ5FMvhd/0QxOj6veZw5WrNsHaY653gHH+1nDvtU
m56YSUSlrQM4IpPl7TtXYkN+A1gWzPi+m7jBDiqmho0Rwxbzdb0JHxKdD/vOUmF0
SzIJ0N2j0sLUkdmmVZM73b1B5gTcAVLbmX9FV9VbUFt94v9S2hKRDt1+0NHpxMSS
RlGOOueqEk5cDHdOwyM6SncZu/mzo9wjpn7IgR/2zZPgJ26dxlgfo4O1W5LmukzP
6caPSbPHZ8BuXoHURMz2FvZEqg1y6bhNniBQlKP57GVBzPGcZ8HNP5I8+KhslysY
pU/bmkoUPx6t/HXkrEumcEMPNWTF9C05KSYf5tqQRVY9ejnOTLtA7rsx2GtQTqTQ
d0QDWGa1icg1OKAZwQgG4IDdQQihNwR18LeuNLuUkpn6WFvHF4/GyBcxMs8ilaDM
8K4qPG5vGn/dDvq60NGJ2qwtTkmD1FpzQiZ6evYiud90HNsCLdnNRYKwd3D9dyJ6
NzlTQvrZkbY8rK2BIVPWFuvLtkwhTuOcbnwy1VqtJ38ThduWSLenRAFWq2IrSDk8
cyq72tbjQuxob5eLjjE2CgF0qfA8u5B/urn4QfORjNEcN4SUTEdoVUFuJBhSsmn9
uoCDUv9+NKLo+LbV2d4ckbk6a4ceO0wd/qD+Iqsim49ZaqT90GVKyHA5ZS050E+L
0ISxTSQXhfqSYVawfe2zTAjLX9JGkpVJnT8foFYi81rHCfuT5GmzeKYc+gZa/rD0
0/uqR8QQU/pIFP2IuoSMWB9GVhLEVNgjEbobY60Wzn6RK0ldD9Z/cMPpgPVemKU7
gpC9sTeSl+HWuQmwwwcCNeYVMVMEJSX2AuoZJh6HPaHKGgsaBkoM6us5COw5CBY9
iplWxjc5OhyyDdpWpSlhaumXarGRQTH5Jbx3T3ldBGuFENQRBOvGKweLN4prpqTh
HJZoJTmPIr1sf4OfAbViveNzjRI3COkd9T9gvmjtMnaYE7YwRcowNGB4Afw0getV
U7LqZQFtPwQflsKTqL6SNkRG1pxQKB92CylIT8Rx3/sVGK50WGKLs+PXSPiAP/LE
e/+bSrP0CFcvh4o1CFRaIFP1k3sgXwu9T7NxBtBUK1LIvx04tqTvCiZvMhBtDpbN
xkfI7Ih0k7iq5PcrV7/3W8wMgtO0+n4ByD0anjFxyVO4FJONl4ykNIGgT58LrziS
/Aw4dBtihlqk7pltja+gJrnDPLwbXgcHElAVHijw5ovZoeNvmjTyWv/n7toKEnHO
i45hNy8INMCmX4Lz3uNDMw/iZD8aEjqAGS+RumZbg0I6zOK9H4P3nu0yFWS9dl6P
6/hMDsOTKabMmZOZahNvHICnVJuR5dDbUbuUPBm9Ay1TJGZDb+TXFj2ad7xOCJr+
GaA0gd7o62FazoSVtXf/BWGlOBxaaEO8V6tzbmm0z4NzTmX3gML5gthR0qYcHyWE
O2hxXyhQ9A8vqf9vmL316B3TlJOqZSrxFiqV/+1x/M/V29KFshmK8fTL377wF8q4
M2KOMKjkUlGsgMYMRgGLwRRyI0nEhLrWNyQCQOgqLnCsSv9zRjdY+ElwJ9eQwJES
ErSa+uM2SoIpuUWzufrX49Hq5mR6sW1QEbq4et3OpwC+NhT9mzGelYDw4CyUEHJ7
iSACeyQrndgQbERCpqska3fiHQ9d3C/A2oppnwLE3tKgMeslCp4vUsSv3/GblXPf
XimNLBygKhg9htcBJVKfH9nYaH8ibkuXjNBV3oH2xf23jr/9LvQv/jp7AX7j8cZq
5AozqzVDadkgjcmgcg+KtJKbcf2KcoNJjJ9xIIsjcDOQyz5UOjOUlaEbhg4wDU/L
cbvbaFnpcYrD9S/hiYEW/fesijU81SKp3OMxIkuMnrMvaBNhm9BhBMmFplydqBM3
9jipWV7VpSYBs70l4wjwZyfsqc7vmFGbe8njDmnqtEEdw6bKBkrSCRHFcIiUqWiB
/nqY4lniSWUgyI0SlmT+40AT0YYWu1tU09voGXSYcngN2QAkV8zxsWQnQA0yDqAz
1v9e0KNM3SVm533MhBphpwqiTj1fu2mNTBDuexio0qMGsTWpPQFSDDIHVHZnVJUc
EuI+DEDvfyJ7sDacB27InUuozVWxO8lZJrcZSIcZk2AnOkDP7arNSAcUfZdubKxZ
g7fA4oMtcima1XlAj7QhGJJokd/J8p0Zl8dqFo11+knP2FSDIgeYGmvJkiwFGYfo
m8t+r/C2yTMpHdt7XmKLgwRUbEnmJ7pUsFzo2yc1kyvf/gIWOUrXa+DAk3LyrqDB
b4CiLt7S05y1KiEXbBM2UQNSRdMaFtebqPv3fEVrfHJ1VUIbMEWYsCucWmz6cStX
TCfqzNq7fRXTUTBDRyJVSq8Agehs+5Mg0qJ6A8US+9mAT48V+hfZkT48wte6wBUQ
kpmqB8TtA3B+Oq992Y/otCKG3hfq8B+QK67XPHfiSHWyzSH2QtRXLhJi9wQiCzcV
Lhv0DrLfB/7/3ZU6eB33y5y4wRjYfcM7eVdJAHmSgNeZdkMAMI5ttY2x1LZV9dkL
76KGYqEG5gvXNJkqF+ACPOxgSrNZ057zA+lso3as48MZPkTPW/tsdZxjgJecBg4A
29bfCdZ0jrunIrFCR7YH0vyvCLP8CdN/gxvGXP5LCangVqGO2KCAIp5W5haLr8S1
tSjWShlWVgc9tINfLtiCProhJWV1qMCgJZnVPE0PSF+tN03pRDok9hs5E705HC5n
n2T+Xxs4beW7HammmTw8/boOGv3YtmscZxKoljvLFe0s3KWMo79MrHX5mrWZur5Q
8KCe284gub2tWXtWTtLDGHMv2owZPn2nXp7xXz0Nh0UbH9HZbFC78hDh0AlPeKj7
5v+zhpZc46Iaxqusc+ZWFiFPR0T9AZggEt9eTwZC5KQM1sgAMgVlIX5TlMhY2yau
ngCuuhImTLHVsItLIl5Wb7fnfkwR/q0jJLOBNWiZlXULCB6tcdA7ZWuXWTMNDkxk
swEYP4wyjitCbocwrm7AuL62GHRkjPdsn+omWsD/3H0qkZxTZKFqBJZL+kASDLov
2DBT2fXu/t+CorDxFt9Ks612vIIKk6qL0I7QzTncb/X3HU6uRw1+CY2zlT8jGjjI
bbnwgZlTrXr2vM+KNUlctcdc7ZucrXjUUa+8/hwOcGStWOAzSiJGr6m8kgHJ6JeG
bHUGTp3Fv3+iRSD4+V3ZLeqANesuJDM7rP3yMCk8s3eaGy6NbXQeAzarYuz5UrBc
hgniGatL7tD1tVZ0RxkmTG4A84n7XmOzHfHA5bDnQQDxhdCDn6D+5BpE6DuLKzri
xTVI2B/EkhhHyZ0/P22r5fUkXg1CnsbOLRw+JqUzCbxPXptBlXP4ltEXm+abv0YD
Uz9Szb0Td9A+mjqCV5UO2thc9OLj2xGtVih5OK6wtCyg5gkfHtngflQQKvTWSSxe
BE5ZUGtNLAHhepLiITsGRlNGHi+SSsW9O9cH1KvYIGSLf2UGNPRMh7Fjft1vY636
Oo7OalGE47fp69/0tXtMnQZWhOWvoGgy8H7OD/3AXi8quDzCcnJ1Om7QY5M7xitQ
iS69VGwkK6ZTczNXKHDnfANhlzmQ/Skaz8l/10PFvsWRFJEqD1i9t4a5NUfmctRB
qe/MlIUF8HW5OPzfv74AI8GUfFQX2NkCbC9NAZcKiwtXyOnGf1EqDr0imJ1tFlnz
OhM7DW1e3MWePdWq9tcd7Uky6MCk9p+MOfaqEZobY2OhGAd9OaJTKNt0CV2kXdiY
eCXQG3sj8G1RP0altJVJV6kWlhuSoUPqmM9NqYGkD/r+hTfSrH5ktpenfx6bf0p/
aoO9ICQ1hJfMLZ0oxyIxUSTwaAKPrRF68rlcffzKpWo1VCeKmgrCHHkQvAkQxqj4
bMZ6q18yA92xsaSTZ31NgxxenPyI7PesfhDIPmIIyW8OettbHQvTIYq5kt9NO9DK
y96Wu2CbyZ8Efvg+enHSIrD/hZezh2l59+SJ8Bh3m8oh7GoBeuuwH9qjAdCDGXpX
p6WiVA+vf49nWGDbuPQhk+avUzZ13SsYG1Hu5Vt1uiVPuSGDKbvkQ/3+JCcElSt6
oUKs3/UcKvXmhG1/OxySY7euRP+0XSo64TpJRSC/qKYW8gBVzfe7n6z//aS4o4+M
c0ZJUITgIheg+83bZ6pKI7MBMP95aHGXqM1Ih+z+akSxCiRJHk6iXlba/bccVBM+
pQ+Zn/9CSrVzL07rZh2v5CzYHX5HZzdbh3kUne67fdxVPCAeccBztuTZ3QY0WBSt
Tb9vV/cE88pkXY+rzeZQwT/U0I/G3lcXLS+mnmXCrYX6xugB+bU7l9M/YKJEJL2x
mCtBsewlaJZk/lfyQE8l9l/tHSTxOT0EWR2S7YV9sGH02+wL696CYmoqYBAMdbzX
aBhuOboKOKBlxqnWjSYEty4+iiRtUzX0NXTbfdDCogL54WFaNYNbAVjkrAlxAweX
UVZfrr6ntZ4TuuD+vzUIGlEM8sW+uIHZPFktxwQWsZkVjcSLQBNTknKOYHpf6p3F
PTKF1FjbpvPNJlX2b04F9lsdqMBCT8koBUaSROhWHSF7KtUp9hUoIZmkaux5n+An
YDH5L3/aGtp0A5pKT2DtiXavEdCFJKFHPrEy1sx+WelfUg7MYF9DFgXe0RCtg414
fa4VyIyiAnIU5H/0CvhpJRX8fcw/WImz1ig11CGY5814a3NNkC+REufqivOyyPWD
TrWDDHG3sCI4JWifXfR+shs65q43gfkedY2ExweUo49I3GuG57f8/lQDFHOOUhZL
0JbtlpzDZ7wJPlrGYVJwcblr/gPwIwB6aGPHCd3j50jJXObAOzWzpTSetRxeHtCt
7IimEw/GHseR1TZsDbPk8WGR4ygGZM3+dzOXQp1GRp/GpbpSAkpvtO3d4cqljvzP
KFh44U5njYj27+QeotYM6RKi6bOkH4QRCHN0N4L0Qa3T1DoqAOdX75kfJ67xR5jO
xajhvScYkIKoffWALkANILWlihXRJRurd1YWQ6pPYcZSKYdf+apQqcANaRkqOkYC
DQz7S6WFdq68eBLEnhzjf/hIhU1GRO5mBLxlbiZdrm3RndH+FSsr+v1Wqs+dAl9t
W66U71S6+MAT+qWw0hh+GU2gTgX4A8NzWJenFT11/4LENy5ez9tmAQ4GPOYUh5wu
qW2H4i4ygoMVy9P6OxV5onwCKpxJvOeGanCWxFAR4SJ80VcQBlPLjBFPpEl0EzAW
WITnOQNTVU3nQKnMjBojMC9ZvbN0hDG4eyVHLVlUEVIjChHqJAgw4J+p7vFj0Wmg
/WZmCVVE29zrLzBKT7xW9cJzJV9w6f/QSj2tGThknb1H89ltiM8A+aSSrm4o9ktu
nLROvO4rOxxdmFQ5oc1uA8hOikxnttb5PqldRwbFVdKZ18SJrMmwufDdHsPcjD2x
OOL+9h3zKE4L/FmAqvfy8pbScoVdIXyxhdGbs/PX7BLHbqL5RJCUT+99QX/hcaj6
S2uZ/5o/JAr9T74pW8wQ98HmXbuTzDAs7efcfngOuN14/ntCZ+aR9odQYlhcg6VM
k+6szrYRy8BwZ4MmMHw2je4urUFmaJPugEsU0X8aWk4Qt1/daqnAh8Bc+yketTAY
DMHM8zEz4o5lWaA/+XFubI7SjmSgySZJVTV7UzvLgF+o96ZXEEM8cu2Nwa5oA0r2
+fvn6SaOSrgt1lmXPdkoU2LMrGctuLu+acJp3+uXcYAdRFPy0JpZREdW54daF8Gs
H+1tj61apggmdeNP/KjznGCMxEHuZoL2rw9bnhcyas6DAazaGzqX/1WuHsYP1T/2
ZOPk2HRtKUqddyEPkcmJjWmEOpXXwYDy4aJvKVAbJ0DjDi/ktcV29OCQr0aAzuVv
mgt0DsMieZm6g+9FfPIOyqnX4slYu2Uw2tPDtBoqM7+/okrLwLfa/G4o96V3n/Ef
qR3lyK2xNZuMZJAcdhk3Y2zbyG90Mtu3E5owIi/zAagaH/S5nF7QVFWmivOUABN0
13gli26KVHhLUUn3Qa5BNEzcma8wYvCl0YCU8v6XMeUISf+gnAX3Xgc/tWfLO59w
osGkJFx53VE4PnjrEUCosbsy2YwHmkJJk9p4p96+IGoXSEpW80nCXSzSX0yLN0Dk
3eoIYF3pPoFSOmdPHQ5Nx4/xqStwJeKLTpuxlKrAHeH5dtT2uYvmMf8u4ItIAKvZ
1IOg9Uotz/zffrs46LD/Fzt4RnMOvCDr3mMYMaXw8ifyWTcxqvivYY8bLeijiTeY
4DkT81jVohKHI4/9MmDZzUmVOkkwnLMcqBXsN8DMk6xGHpI2rgli3eemKqj6wxVn
LrjGyvKNIAzXFIn02Z6IiLXuFvxWpFWS1NM5WarqOex/TOz7oGCIsCKNBC44KvYk
yPJ/kQVSJNFkqtFanZ5Jwl0YSQHP3l9Wo7FPher2GONlM29hLFfP0ek1MGKzoJJJ
9Ciy9iiyP24iJAkHEIa12IgkEtGDagPeNZLYaJIUXse9Ph/w3E4TXnbo8fnP4JFm
nciaYJanmhF8Axu4MaHGJpiXs1YI9Akw8uqRsi/+C1KCQbuBN8/ki+PSBlOvfRNN
K6/zm6ZTball8+njKwTnTdGRJ+E4plT13DATwuuh7DcYnpb+6RENQRgUz/4wIvjz
pOYqTGruBFaYg3/Vl+fBgbsuY7mhz+7jjfAjrGUdXx9A7YC/aJ36Xer0zOYpepbx
YyXv85ZHpDpeLrq/ZFfhJMqwBpAXQGxrMMELKGVcpdJmQDXGLnaXmAO2FXpo99ox
e9cOGQfYjpUTXyFPl2GcSTrsqtqatd+O3ezaUlZNN0AHesu/0MYHbFqrpFMspqjX
H1zaX8UFic0T6Ls1zzcIskFQ7GXu7P178NUJL0IWGv6NA/RCxK1ow5JIrmRSg4m9
ohhB/S7vbEAiHHk/FpCx1qy4IkMo4lbmqmQOcxtkyeU6b41+4UQrnWKfxcenvGMM
REMCQ2CIvolv+TYRlXUEAT1vnX6dkRvb29Xg2rG9Uuc9400fjW2Oyl1VHpqMaMkb
x4GKvjAE+lwUFKAdUSCvIQpr+7ndWFZLnBNHYpoASGTj95VZJ0kF2cPZEkQEdG1L
s5KDb4oHldcYabjn5boX90PkAqsUKEKx9p7y2+iKLQnKX45Obuu9GYfkvZFB2Ov4
aO/FrhKSkTKKjDSZHvcy0baN6gEU1gPoOv2STrG0+UmHRS8gmzGHKORhzPO+K5AQ
KazPQOf6dnPHXus3GclYT81v9A4S8zGXxNZAy4CjIte5cczjF79iiVy4P60u+48x
87rWkm252DnoyzAX/HxOXtPyJ7tJmLMa4hB+fMSSj6RqsdYXadppa4tfWZtHOIop
w8aYS5giDjQm3QWFRaCCALclQrLBh5onDTsVEoJcaBz2geplBjYBJjj8XElgVOeq
5tqHdpBoZcYCmi9/RKEdN11YlQi1LiPdukebF/Saqa68B2pew1cGmHrrico9fW07
jx5Kd7WjKFmRN/MZXJOhtzXv6AkqSoU2yx0VbIcqa/7wsYDieHyAnAOJqc64q5Dr
tw4hskA2dAva4B0oEy7sEQ3ndG00MQ0DHV9koiNdhDkNKn79ufkynZCTuL/xwzIw
OVgSVBZZXOfS0eVijPYQ7EVKRNyYelpmr4LL+aL/SAZDbo57c76LFm26q6pBCej1
uxHgMXvQS9V8acxGt7UowQALtIRh9LLhM4HRB6uQxkvzu9vmIG9GELgnF3O3KFu5
pB7Kbmf7X/lSpH0YtBAo1RGvWHBnuFzfXxS2En08ItxKQ3a7Xdtg5f+tFRVQmiSg
X/vXcFdb08wauFSrqeM8yRszv3HS3gBsWvEnZyQWXbHqH+d5lP+1F44S0ItTtTiB
XuhP5xzj/eQyD46BQjLIQufsSFUmVkIVrtuU0BHWePvKrfu1tLlfhQ6FNrePZ0UW
S8Nfto7zB1KvQSNk6UWSYwCW9qCDo95FK6HY0MAyWFkxaPn3uPRufbNyT2a8oMnX
pI6I9sX+pDK8o8Anb+6xoi4x5OkmFKWkysTkDhyZ59ljDkQwVIAMiOHzSjLeSvU+
T5RG+wZY63JSH8R1DCqReIPdr6Iy3QbIl2eckKQN3qVSpNL5x+ii3ZcmUmu0CN7Z
hxlvaJFrIDCuMRLinMSbcgupRWAISTRrAZfdkfMxVYw/vgO2MYPjqjO8kN9DHu36
V65KmiIs+wX/vbx/HARv/TUW8/R1cjfPqR6jGzgp0UhjY1Y+b13Ib4mmzeF4Sl7P
nTG/aopqrlYNOQ2FpabsIE6KAGzJAPYSB1B/KtldFs7SvCslYYOoXQ51iDjhXkzt
E++k38fSEo6Olvv3A7HTq5uii06Wtjbd5zDN1+rhsnmyztWTISn/E4qKznPMiEfY
Rqi8xjYYmS77m/gnAGrIMJdC0CEFT40LsS9IFQztGSB7fEqrz3L29MpMMsNX80Yg
M/AJglnY5nYdXGdnNxA+huFt1l+UVjSzNcK+o/bOCJKcWsHBFtiTgaReMBDCF3cy
/B8HmRcJ54FyQYZPaULKLkCRjHgakJ5PB5wbr/2KVfkVZimIl8PlxO7DLBUSQ+AA
6AJYN8WPGdslTajJhlLq4ukKniEOtPLIRT80V+TRjuAsCqPlvu/1fM0dQ73zHU5t
3JsKmEYlJlHSRnxhsbDWrwopEkwiwGkWGE5x97zSKsCVuA3AWL/ZzvATUZpZKXJP
FlpLdkNKxjmE1KIREeLaFIBhsk/T5BhBdN0ICnv2T9eLpQmzz7gHOuHsCwNrFP3J
ghHsspA/h9IWKNSjlQvMgxYom/VWJkDDAZ3bWuNHFNSbgWAtAKZ5Mi2jCUqX9WEH
rUqPmer5TPKu9lKgnaa29kvowJeQmdUsiqOawZQCdVGn2mmt24LXAg9zST57Uw0N
ikIl9dqQW+c7VkE4p+fWf9JdYsrizIuNsd52NMKiFY+/HMzzeAZERhl6Ry6xuTgf
+YUjsjnMrcM0kUT7QQayqKyfVZKCj++WdRrZByyrMrVewQMzl9pCsnorQZlrlmsy
7nw6tHwtiFGQgUXDHO+9Ety4SId9lTZNlU1NtJmSFsZbgs3cT4Rrm2y72OOy9eTu
LaILMDltAjvCYNH10KC/AYjZ1flUGY8yqOlMi4BQjtFSwwo32/NKpMTMAlYnFgOu
79Eh/W5wgZmESEY0HURpwWRqii8YEMw/JFVtppbm5BqE/tXooeqhjuj4drVDAClN
CRvdBAXcDO7TbHveqR1KG1lMt+kmCdWCvG/iDvi3zmIKSjF0gvZYXFMqkWn0XLAX
vCvv0mpj3443CNExFtto0rInH5VZU1XQDuHDeBi6V8OTgtBgPsYJxYcziHJD8ydN
Lm1enOkaxs0t3NL97GkUYWLtc3Ump8Hhj4JHAY3oYU60T7PQa2uhd/oA5dKPhzMK
mxaVZDgBZeMUQRLsz309P5Dk42t5EAlrS1G6EnslvJvLykM0oOGAWWVEiItsrDn8
EyiEp2HcjHd2Oy3iHb1xLPOGHRkQwecjy2WhGMva4E9ygWzCpulA0anHSyUcZ+jL
k5RuQpMn+oldj7OxpwSoNNQuSuFRXAztr9UPBVF/QEXGOnRGOdO1TW/dcy5NsnLY
W0jivMBQ2aMGdj5WOJ8gJPniLOMrbz5Wuj4apLVeMwxTF9Ut+TGYZVwBfgfe4AIe
2XZT+w9H2tOYx3GXF1L2XbfLpw3UdtM/c8s870iU+wiGEsxpJvs2JouRGEzqoB0C
bBVVik6fp6PxZrf+A50/F/WB0XpTVDaLhYGqbjF0y/7P2s5I3YanjJSU0Ja5RVPK
c/c+i8++kCQFSA7QtnwP6fMt/Bu/wkIrmd5jgGM2b2GZm/Sv+W8vITiQhgKmeMcF
mhdI9BZwYmYrzchRKYF0jSJZIKV8qWDzbkaBSGXQKwN8jC5Gr32FZD+fLhk9KpGg
uTNup0v40krMZNglr8MWt4hdoGCD20tCcKNOOK9dclSLEqPYgKGJAbl8MLJeGgia
TdvCeNHyun5xs0X9VJouaW86FelQoytbBUtCn0XK1y4mB2Kf6IEzBsu5xu5cVd1M
fOj6UVfuQIp0bspbeMiZrrKY3GyHJYKi0mNdSNWyXmyGvmW++E62EmOGNU3Y72p1
moBOGLgAhPJK7Y3G6Rw4A/4OBWMFNnW5+u6Wn5PDXZo9ypeBbfjEZGKvrz2iezPI
bTt9xobMvOiomxV9SSl8s69mvj0aVSYH4sgNoZJQa0JAle4yltwALKC5PTeH/K7L
WHaRCiTbjvpUcW4gndQZfYp21upma4W9U74Rl91572kmdi/wShTlXTa2EYiaO4tn
xpmA4H3+8ceAFz03F6Vl6DURCf0EDN3wqmDkAzLgLSJ15mCwTn2LoTmPTPqBdYPd
J8yJwmdz+xZgj6OdHA+VzrIoqk3RwUBk1PDiuP/fP8UIu2888AQFFHbyrCNok66V
B+wtRPYZzE6bP+mf7e4IakD32F//ieTqQAaOkXBSkuKOgVFOXqWdoVE4rdnvZGQe
kCzh5zRdwEtuwGmxRuiazS72YDdMABHmvCj/LOza50Kc5483r72StHQOtbWZepu6
bMcA3wT0cwPooRHmj0yLP7xPTF7bej6s1+1aySKTCwsHgD4kgVVj0egkEEh49zQb
hm8yS17mTirEtBvE84Gy1XvCL0w5CTrqae4LXjURt2es9U3T/XmMYFCJp7tollA2
mp4z+leA24kq/1hdgUM/ffvVN1WpL7/y5SmYQ3se1bNl1lbJDad0bPMd5v6frNj3
lokjBp6WUZZtUWuwNJZLgw7HZB84GNb/WcvWU66ChUfjfektDWLL+1FSb1DWuoIe
4/s/1SUuNPayIRMaZWuNg2SutXPTm+H2mZrw2ekqwF6lEn+An6W0od44Pr7ePyiX
JjoWWCY/5X+g0c9XpX/iRmQqtTcN+RxdebVLwuoZuqHpScu01CHHhRd/Q8ZHq5cS
tOdKNzw62qZ9q6kqKZnXr4SvxfdrovvRQFm74nOg6IVf7F9PDDJRgco14XL+mP1V
lzMU+4hk6PQGzS1wWK8z/vZbtRpqj+WY3eaVYeLR/sD0hrE4xVAlMBwUFrA248e8
mA67IKoU4Z4YkmjYgoq6k78dld6Z9XAMFnn9XkO5WDpoKE7OjTtrNYxXRG/pJW/S
KO5ep0UpcuM7wOug+lU3RQrPgqwcLaxHjIbxByxW1gJizosCOV0a6ydNE77BCx7E
jmT6vJe2SWGLBr2Xmc6B07Tk1Xds0ayy2pVhOiDKmjZ92Bb46A4B8E2MaMfSssFf
GnqSqQtMVdoohfXLcawvelD0UJ5+XihIeTWOP0O6orYen6kmXBFahhCwdRWDGuDV
bw43XeJsoCj2PEqLN/TKKLCJ336SHBolQkQR2dbdwovJuz9c3VedvKvWna4Toy5V
G03CtQAsULbaKMgRTq6Byg2hbnse/U0Ig0HauH/xPtsjksKibGRgsDJAp5C33Wc8
1fRPpZhurMvrijHNu/VoKUSEOga0vJJ5VsMlZF7aO3+cu1aCu13lriPVUGo3XMAm
WyKFue3h1T7UAlG25Idt5/C1EcrEpKL2NT3ysJ0pDMh+3fBKC3jZbv/4XtCdsDfN
2rNQpoWcCtL6ltiibG2tCeT/ce2i6VmAo2kr1gNLct3Ek+TicINkxL/gcbwz3oUI
g04lUnrmtsXBP0ECC0UVUVCZAcjYYCxOV/BvTISQDRoQSXIqvM1j2pH5wQl2WiKr
wbUX+t2+FyVth2KtD0ynHa1EaHVk9uTHLq07bot/V4y7y/C4VYIYeBVRBkNeLEcn
phWqKobNjvdt/5pavQ5DOfM3Dzi1pugNoFVdjD/lSn/2Ih5QTWGvm9WbsD5h6uzX
tu/1MJRKfwVywEz2a8dBDVGX+tHovIu+/kKSLF8AUwee+LT/u77qPWFb1GMIel6O
KA5ZWcBGOsQL9X+9AS5AdE3YbwegawM3pummhSJtZiRRMVKHvj1zY8FPK7/honcC
6uxnsCoAU/b7R5Pk0ju1/THzbgp1c0aw6Bvhl1NsNWg51WYzYU6Y40lSu2YIuJ3j
8cRUepO3IPHtCOifg2ToxZp8aMJrjXm76N1ItBWVVJndxJ+ZEiTrLKsozdSNeaLC
QV2Yn/5+8JQLdEEIREZG2DAo+Lk5W+53GuVMnbSgpIRFBLMwEKOX7qWDrqYZd0bG
GWFlpmawH8bAvucvUpTkpALv/RWZKV9YkH9rEms6IQgkXzeAs1ignGLMrMLD10Eg
DUQxt5AnavhFlL/ddc50ZZtKjZVLo+TpjuyZIqFD3l5JZx/exaBuKNcMe6mXSbGX
OCnUwded1vyRy6XY0evfZxemnXMpR4LIVzgygtepCQrAw5sfHrUs8UUD1snyKlbw
kSbhGibI8sh9wdHQRu6dWnXp/jTEv5OrVrMHwueFf15mUWXin7ILKyE3qgy57N7q
g6gOsOYpSGhq2zya3IRiGfabuth7/Nm1RpICB0obeheect2D/U/8W6F7eR20x6MN
Yf1onk+XXZATR2eAyo2OiYk7DMqRrmEhrE4XC2B1FeZTt057v8ocuVYDcJ/uQfes
x2Nk9fzaqDWL59QcJMsFQLscfvDC6jLSxG9fhnCRw6yUzMyywjTFAoJGHShwrlD8
faJ8OkYg9mB+KncMtiG2dgTzXRfCVmpL4Hh1c14tYC5j/+KOGfXA0p62pipKYbvi
gl56cfLw3Rbyjl4rx+M7/F+91xsTLAQ48TajcuD7MWwNPwKF3qmGAVgUlxHYYMkN
N54tdaYuJVB6L4GUHGbm2vJ8LuTrclAJ1iHuxJx/A3+ymBdRAyty5hqdhliRFkeb
OxabkSyiC9cpb14aAylTLV3OkM36wULZ9FywCttLLX1UjC4xfXHl5Vl9ZYcOl1Q8
iPv5y+Ubgl/SdqyfMtzPcaruBM3dYvnFp7OFtqUmrddZi9NV1ADDRNW0cHmctBH+
6w449IgNZGTR+YHV5LFKzLYwxDLlTEiSUow7f9iN2sN+v1FmnsC6/etQsawg7tWV
DQ37v/2cF/PwJ03VHECcBB3gVDijGt3QAkKljKXIx9O4XMIe3s/03LCbh3Kfrlxt
Ki8z6wuYinOIVdzwnBQLMH/O0S0nWWcsxWH64w/rAubWrbnt/VE8wx5Wu10CmUSy
IuaqJGT57t41acocuhJXjgsAP7dDu0TPdQ0JkoBOdlf2O/EeAsQq93tQykudrQzf
vRq6IvjS6gV9gi0hSeMPgl8ZPHX7yjM27g4Dm7ILvWlEppYz//Af7Ny7pQ4zwIPF
Rw3MymynA9jw1KPFTrMG/Q9o1M8x6kehVlFTcOa0jRHgQHGdAcZgILZr+J0FU9Q/
u/EDiFuDLyIWWOM4YwXAGPpd0AO9mugL/xjcpUIlFuBZY49A6Hqq31x8QNg/OMgR
qurEeovWxkZWzfnqiRbdflMgKahKqYfZCVCVGnY0N47nCIuwpbAr6ywgKkNWbGcv
S60Co0Uogw+OzMnLw7GUmknwB+HUy2slg26xYbuuT59CDyCh3CdmxvvqLVnU5EGl
o9zuC6Hel2Ac0uNDwhfF3QpJT8rg2kRPvsuCX7gDT+ytcoT3s7oZPj9WdGZTudSr
XdJoCeN45JoFvMJDYnfd5nwKQdVHlFirPbKzRgfTCg8xRIm2WAVn1KzO8uKvs7AR
ccEi6XL/enBAQIUyhkrIo+MvhTRMnMOHy56GrcQdO2h57HTrh4w6jzSl21a7FWAy
/GPFKYMgjL87AV5HV7U7+uB+DBSoVr6I5cW2swypBPWW/IgXUiPTsKglyPAcShZV
DOSLoX+q4K5FTRQY4QA1lJUuLvfB3HdIGwlyaRTO/44CDGMNDrfdN7GdQ7ASDWOD
sEgdszoKsMIubuj3MvCG+EqUp5sBfqlA+28MKXNfovE14cCLEB6FcSbtbc6UYOY6
c6IzVwtP8klkZQ1Ii4JD7CIz5zgIqMdxi/Ir/E43cWqbxEQ/2kBboda5p5S/qtmm
kZq3wdwFrIATp8rbiZgAlsfZtnM7CU4DMWQiU6mUoBcqJ5EQ1l+JrONGq+oof4Tr
hXux8c9B33g2CvvGYRUW5tDFa4a/xlHVNm95sTUEkYd/6G0j79h7ifO9nnMqf1Op
4QvpCpnWxxA7awXhrNMb/uohBXS7hmBu33e4H3laihi6uOUhzPW+Fn+vSfkv/Dy9
IbLWGB72YYmkpZedTd2x7kcciYJL6hPc1lbBJF0hDYTIe2E65f8Cyhv3y1IDX4qV
umz7VFxOG3jZcK4Qda3bOeq1G5eA/N9MVsFFa4WcmdtU3rNvixiYtqWalnsNFjC4
LUKgk2hbh0OHQ0ij+uu+d0Gfn5VcLpeBjEY4CI1xjm1qhcjzQ/URagBhQ7wyTWd5
G7B+9opewMIJiOkUrKmZh02EJEi1NOceMQOqVye0HQ15ySMg9r+w9oDXEBQ8tXjO
SAzmCE/EXiQxibcDQ+CcCdH3vAQ3ZhldET/2OzKdQ4OSXSkAbZ+OGSTKsPnWq/Su
4FdyGna0FzfI6ka/Jyjqdn9WVlpxLLUME+MlcmhCD8AEXVOMeZzqOjuiAGnEIW/k
LxKSI60wnX0IZ0z4ib4ZG6u12kGB+o6Ew1o8laqGA0+VTZgNgtKGdYWGObaKJuV2
TKWZzSqMR0qvOfNScB1XCfNNWDJ7RpHwVODJjWyFPdQcdYTFP7+OmBUD3zVArU9T
pSSX20s1R+1w4d13HfccfD7AdbUJWkeYOJo1IxNPTPnuXPTfsdM1SLcY/WF08Pey
5it7y6Isowvxj90BFfssdEJi1WXDgsRkZLRHw5S1U+ZOIE35Z7GaKAkExz4gghil
fpib6x6p1pZcqnhfWkrI5ZPAgNiWHTT1ehxt+gNsBJIuxb5tiHZpJCzhSekahUwG
nBoX3SD73zCTX4dIbxRVkSRCPuoEvWk5WQtnTPo7UjvN/5DRxbyBS+Hk3UiI3lPA
bS19baLlWMpoBpSfdr8T/pYRsqP4HPDphvi28CkKT9tXZMURWXKlCPl4u1dnaL6r
krkR77QqgvuZ6BuJi2YGjcBlP1KEomjhw+Ff9RClLINDuSTnz285zOOkd2kPv2ZW
t4zKljiOCreJut02ZH2DPpc2ecJoV0sQ0u5Isuhs1hFF36GJGO32mqoDY1DU7ChN
4z0cdVo1SPvtle2pljELOkgHcVpcsEtCEQ83t6XcupxKlXCY87Zn39oaD07Vd4Ob
3+rh+vkt231aCWhcdLxPF8m++MLkreV9VkNlEsLG9XheZzOlCEVNySRLFL2uH5M0
lzc8hRfceuHQbYoafmMfexJiGeM3BIfJtxr23WhNAXV1VKhaJXeUPbKBR52CZMaG
82vMSZQR7Ov3yHHFGPEAK+AXQi99S6xDGg3Q8QGJenwbRiu6o5cB70Cm0Jq8MWpz
T+JAjCSD93/YyLKxm+aUVsHIkKAi5U9sl9tRG9Gll09hu9chgjFq6mnpfzibShGL
WOWlVZjZeQY8zHglwMSEodDQ6lk5KzAy9NQJGbgv8jAKHvcJo6VceOasSr6WH7Z9
BhVp8J/VBz6kDkvlpdiYFBYIMAeMlkx5TaRsLy8gY0GRaw2/M+i3tu8lQtn2jaCu
B98iwDedcbs40d2pnkGYClrSNFVGA8eLJCajGybHSnHhge4966pPCzEUhJq4U+7f
xYx4vgpTZMgOdphIwtx+xSLnsERtPJQ1oBhw3ydDPdoYxIUADRcVysDZ99nw8Ybi
DOTFDMZjwE7vHbKAwk26s6OiUHbPdB5Gj9vG9ohwh7yo1/pqlkF+KqB/ERmfijPp
Yy7s8mt3u/Dm7YES3mPL7EIjdr7UmXOEEFxek9sOmoNiAQ82QFqHEQC3aNh283oD
nQ0jsSN6GRPk4dIhEDvH7OLhsbOzZyG/OAN+NnE5P9WG/WExgWSJG4YQu8nUfveB
VIlshHUb4VAT+aa2bpxjj4kRVB9VOT3qfbz24Mr6BLvi5r1Tq1uB6+dvQ09jCeqp
/zOpal6P4Z20RcYUU4ASrYQqbLIICxV0/Sn5M/6ILvBwKX9zZIeL2RsXHtMdXUb0
F75gvVAvBdvkZ9/uKWtngbPvhidswY2e8YfqYOKJuEMfQ4o1zoLBc7LZwbGhGPwn
opy56XvB9miFfrrNIsW/L2LnzWmytGQbD5A2wzIK9GSZe+WC/wsvd02fcOw6ZcWd
W6Mr4eNYWOXBjzorcpb2KHkdIrVLS6qc3cm3hLdw/E7p/rcpIzNi9TO1ExEgVVZ7
7hDagP2vSNIUD/GdJrgCI/0XBAzF0BemPrVh94RvaboJOgOs0R9K0vdWB1azp6xq
/PX+YB3pYYGkaHdN+GR3zhS5jCrzxPkI8EV4S9aIQzjniI9/vv7fpTAB/Y8HossB
yRm8q+PPf4R1fEbBWJzx6j9N/Mmds3y8EagWYUt9q2DSew9Vhk9lBhtK/HKwf69E
BZhBJR+stfsray7CyOAOpizANGpdMrPFm/zvfJQkWNY7TozZNnrrLdBMjHRSDqVQ
UN+Do2MiSTbqZLJR748L5TbSi7hrgMCPxfs60ychSLYAUcqhE736V7tAhXodZrJj
mEba8HU9a+/SXgxGy35NDm6qWdEI7MpVHY7oRqPJihaBw7jGUCZGSh+XME5HUjQl
2muZ8pO5r71N/KuidKaMKm3ZnvRvuHTX77Iu4wbxj8J6EWYlbJbynPavNtOuHPA8
bT+rQSB/AuMDBqTF4bdBamHWK4zP9a8atlyXX8vNRiMOCKTY5f2yhzP6v1hjJgHH
TcmtyuTPSAHtYJBAQNV+3MqtVqZlyHaD45ug6wIIE+fx2kFW3jQlAccrbagIVFLX
f/uW2I6hOkcPI1TJACk1GmV8I3MqX9EXg9NJI5EB01LjXpnA5Xbyp1ADMm1EBCOT
1xWyQQIMgLILNgHvI85EqWTfu3GPEZclvthbl8aXkCKmFx1ckwU5Hmi9j0IrHVxW
2Ch2woHAVR4wOumwtFajf0KYFFOqelBsdFtxUzwHzUcOQwzIBaHOOtxdn4aFZ0mM
FhfZj18kazOKdtCQzpY3LllfOZecyfXSJ2hV+pjFbvNCLCEENfHoqCxZHGGIv4eo
J2NG/NrvTsoF9SJzFNQ0z4aQoeUA/yxUlYjX+V9jBrboORTFV7VhuqeoVjR05m3X
Ipbl0O5sr8SvWWozZV9TmyPxM3TWctWjZIpjIlsECYlwqs5FB8ZwT57zV3ujsVWz
X8SH0wi4+QsyQY9L7bcjKH8jurPj7o0DVmjhZC7b7WLyEb9pkJG+wh03Kk+YsZWm
hZdZLZHi6/QaFJ2VQ6OmpaoghnvidIU0zlR7MFa/0zduMWO6jFoabUyVayVJyS43
jgVhakw2+AabJBi9eXXZo40K2vbxLm0cSU6VgRr3sUQMTC3hwe0pV43Ln1M0NmcP
AmrzUFTSS7f//LQuinWNzxZl03Dv0Twj/u5H+HeLYe+KWdhnUHYeqi2vRwWLbApE
boPgSkrPesFyUGbBg78pXmcwYrIboPQOMxEMVSoGudtUMHWWh6r72u9lVA0oPmPn
SjD/wyflXov1inGmghhWW5BQQ21qXhOLMO2sbCuZ9qdnR7bq961ecEssqx4nRkkk
rLD02vpKzziz44Th5ERbTWiwRFH+i+4wpXy+RA07u17gnn6Und9hJi0v5S0rd2xf
BFgP/Wg98Qez1RPWq7baAUKm5NeWnVtIyuqa76wB88/UytWknBFn0FqUyeYocSHb
yLbx7omQ3MZYI6Az5jYJ/MhXkLtjOQhhY++JULqgShMWz3dZp1dBryPqFhxZCDY9
OWH3698Ewa6VinDh2FSjNL1ZW/prqWDZ6S1tmjFWBBURza5FcEghD5mM4tZx6Q2f
rUrbRYrXU+C/gkomosVSnNqaGMYrgYMinJxJEZqOg61+g6wGNxgsEdxLifQtMcYu
/TGrw/8Bvzo802qQLcbUc1sednFGhhgPbys3LgKNcUly2/k76Tsbb40hYNApt0kt
h9WmKXiG536roV9NZDQgb7WSv0bqkCV0e+/LJQi+LDG5rXcuf5OFSaiYf5RhhPyn
uWD0FJ6sSezbj/muGQJRTT6f98icGDeqXSDgdRwe44hA+58Jx6hAMtB4xrSKHTDn
xsA9Ho5gp7nWbX9u5IbU/a5Vi2FFRAJ7qnemit/xoHi8EAsxkr0QsSaVhEi5tkvi
Mu6nLtWbkD29opsmxqwGws8trAfi7QbTC/5h9Me7TVMZviI/ZXevxpg+hhjuiMWK
b5LK9CsRC2n5HUzlro1/nqYJfOqy0wdW642gasPB2QUS9YQUeCNboE6KUAyPxf9N
BankM7SfUsTcl1MUgNgbYUQgvNsnpxxbrosJuVYe8k/AQvG893waP4Z32WXvNwSG
dH9JX9kthY7XMPEq3+iGnQFR6HElma3vujqquHvJatF4l1OIXppUBOnuZYjn6gGQ
SwwA63ist1ZxXd8oPK+K5/v5bKg0eJ7XELxyydsOPn8X0cy6ydag7IVqOrcLV4jm
aiTqkjnouBMRPAKiQ7DzU4bv6lL4oShyEqr8Hbu6SPyrftEwdaQEfeMsdwWZk1zM
FuiTfL5lzAJW5gjXiOQ06GyeztLc4MIIMUDTSYEokRg8dLzliwd/xz8vkyzVngP8
cip3rdsuk54uNr+X75KMqLUSZmgcggp4sq4ZA7oZh3q5xb4K0CTf7zuMK0sl35IY
0JEHkmVZIXXedMsIwOk/3cvKoFUnSIJZb8gYrpKhj96upr6me9nm6o0jSjwXGZVq
M6Pe4FV/jXskOZz/YY/GrzC07DvOSk+xoYDLazCnFhNFxmJPOqqZHld/ywWUvP5s
l1ZbS+1jSUIO3eqNCUC0Nh/kzQe5T8Io2DoTI0ErJ0h+sipKAqgdCX5SCW98Hc8A
wjkyySxnPOdIJ/DP6TqkOIWYzWy0u3fG647CSl5VrwZyX7QBmwqQRoEJbw+jYm2E
64w8QevvE2gzMJNV/562CIsloXYoWAXPYeNHL80YhxEkSLKo/tdeIBpmgWFcd7bs
pMpLn8DovAV7p7VbMH8TZEE0XSBswRz84LvBFRr2QmZrAUBty0Ht1ZiYCMj93fig
GILcwr/I1bsBelFYnqDEPAMx1V3egt5rk9AJ8JH/AuTW9xz/adw5YxUUZQR5RCf5
boYZryns7tDvLwMXil9ushq51Y55yyB7+QqWuNMbHjt9l0Y5UMEmD6k7K1ymoZQd
wiA5BpvJ/PW3qYKJOUZTFWcaL7zJkvyjW82ZrZ7AilP3ltkapUMbZbOp2OoHTX6w
HrNakYTk/eqWiEMHCotcK9zfh+i9ybxXghSPGyNN8s5yAQ51xnf5CDktyTA2pplE
nf6Og97VGHBz34+UmL9PTnv+mNaNOfhCIpDp4Yek2n+8AIBUgkt5m4zvIxbqw480
+9L+xC2cvP+eGNQEhsrxMbTHbYrrWtLOJBCUj+LriAKbHg2q/uHdPoPk519b0t9U
tMhqQv3QzaKUEkKNNmgiZrpU5wQUm2imeJw+87VZjnHI4r98jmfZbFAJfH0y8KCS
pvQzYRqNm0g3oB5Z/BO0tFpiwWXRWNDy1NqDMa7dZPTSh8FwyxdwPn9h4j5wLR8A
a9cx5lakd9VU+GJrCxBV4TfxiSqRZPwpYDPC584XpomcoMDWigbAnef9eMy/Ngrz
ghgkjgqVjfGXHN1SLkOsf9xikYy8Nmz0I0n+BYb+Y5zzYyt32mAewb034IEpPPrF
cv2jnR1GT0v36be6+hE/lJV0ZgcWGflITG/K4y4SflRUWobCEhWaKmOyfQSEHNJg
8T11XulNhtZESMhmxbLCWK6LoVwvoSZWJjNY6SkNKso+PDYlxXphqP72PZMdfEXT
9ItZuIJQtP/b6oNFzYhb25r9m7nbNpqYbLBTBi5pCPtVzDp8/ZWGx9povBbxJge4
jTMVthSQSqrkaRwiqEXGw5r3ictbgai3kaZkRE/TJmoeZTyeerI69ERcnVn00qEV
TAWJwjWWPLS+i8s5XTpPDId+h95Tk/X3atjQqe9onjwOTLv1p8kNFXM+nm8A7lIe
Qqz9glUdKc2HyEB3yHGvxV/w16QPaDAWCWdahRRQdleGPqDvm81D3Oo7PwDsI2V/
DPHghFoMlTIcjUoqEbWAKZqmCuJh31+XNlu8mj52K1/nxevAXKS3O7qesK6kux22
SdmNCbp0U2JMNth0A9D8WKWtJy+l88UQCN5G8iXaJ/BuO0k0WO9tshU2sgfqu9L7
Lcuhys8clXZt+b8fiy+OeBxg9mdggpu6HWm/3F3GCdwbGfeI2r5FOmYeiUUrONCV
iMyeJG67pLLf0i+XgFkAAiXqww7qqpv191Qqv6jE9Yfy3mTpkZg3Pt21juxJyn1X
adXB30kbUfuTrcUiaAmci7HRXZWpp9iE3yzL4M/XLbGUXQwPQovoT2DbVrmal1+l
0xpYzryKvG8/pmtNb6o3I0ZrHc7CwgjH2t93nl88VxPNroAng6OQIuyxFTE4KjDZ
iQC9r9wznXXzmkOu2xf5PDjfacRZrFGh/udy9mD/IcQQR2AuyCZlSOY7uCpv94Vl
XOory4iGdp1NO+UA8D2knJ7zYTjY8FyTyZbY5Jbf4WF/3ZXVB8sd9MCeISx7h19X
eScIxpXv+CjHAv3abHwci773yEesZe7jnGoYbcAQLmox6dVFe7vCvtyf50S00IJ0
549nU0PYm60J3Tx0brvHXGTftQ3SjLpvlM+FxiEyf1aZITjt2VmG1EIazb28t0uk
7wglvrEbm/c+NwMJ1PUfluIJhKIDnemlBmC3F6cMQ6KCx0+u9mOEZyvTQUvp4q7z
7h8xwMmkYE04PTgzwU0R3fC2Y6Fe7/TCpot370NYQsktr1Rgfi7V0PC3TwioQfjk
gZiId2sk0qEfqPF2RoXKJigdLxwQ5sMxZt0q6DflsnSAn62Z1xncqJxJ7WJkGcBv
neuk+OmZwJNahG/PldJTVLUySv/Ahn233iOramd/lo59LxA8i2R9RP2tisZGmlsY
Ke+3OaAU83VRfi3lnP4B6gt7DznCiYKmEmruYRGmX5L06Ov+nD//HfRdPd9acjBS
tXxTWbnUkSmaULBRN3JEsHs3Z7XX8K6u8jOFtjpINQMgpfsNw5kHSDKIZtEM65h7
QJgAnXy1ItBf+rLTAfXcLIYcTQ5q0vrLjTEapv19bbVKYZiFe/0R1AD/4xZWUyh+
KiJC9wUi/cWn8uyAWhJVXoUYNER4v4urD4cxB0SjcCKDDI5CV3pSPXn3ZbzCkpfy
65WZkVFf8s0ErBrVM/Dk8oXNQx6kjG+ZrsNIOe0ndOag1nb/64r6tnZx2Tot6isU
t8y9HSqs87HuSZ0CJySy8sIu1GDjzoUCPSA3HF+2ny5NmKeaG76erjbN3Xx7CUmd
NxshLLDG0OFP4Acr0H7g5ekMpMFZtlvmCIakX7lT6eVUruPA7E6Ba7PAt3E2t9yl
8Fk+yNqvhLIm+kS+jCAxL408Zuj3gKBw2+B20aAPsfIEe3HycmeM7++rO1gj3adc
XEf4hFR+eA74JKc+L+mZo+6vjf/gJXyWvHaO9YN0813FiaDvhV5qPgV24DRSYlW2
2VpZXi+qMgw3g/5hNvwakZPFFzwxP6ORTLRUqxBpvWNuIwkWGii+lTbAVxSiJzla
dcNk7f+fcX0DxmfbYF4qT0FSk+QDrIqVkspZRlMsRnNzu+BVqJzFrvE/K16UbySN
ZkcAGAGgsQVvke8vN1spQ9c8Vp2ww1ObuDI8bSjj8AAydNxwZn+L5kVSh7JcKFU5
DFS5uSG8w4QZYawlKewHv6RC/CXI3p5HMHpMAP8Jy1DrQ4oGqaEdYWcYnkEwzCVc
2JLqkBEW34Tpo1bNu8Bfzm15ZtgHlq7HF4Jf8egKG8XRiZJujopAcd8yL1pZVbpb
H6Ve2k2jwNH7q+GHjNxc1qz5/o2gthOzvjv9otyJjfiLaHGXZdBwxQsI6mb/o/x0
iGpJtPLu+HK2QrCiBx6DamtHA0m0xiyt+K0HoPSdSq/5NkRAUm3xDerQXea3fmlZ
dkzQJ1EBi9Xdn0EcjH/zunTaerpv4KmAhpBG150sR6QB+sxTTcNSTp4Q8x714EdV
kAdm2GFri9LUmDeUKh//iPkVhHBhJAQs30wKtTKPwxcD15ZfYSelrg5ZokZtzNFj
ngySWpzDDsO/9gOyPmDkVoO3WHBY7Sdio3A96HvCmH42deIMXbPZcZOLD2jk88zB
g5YFfcb+W0EOx1ZB0MXm94F34S2KHp55CKJEvqYpd7lB1+e4F2INPNrp6DWPF6or
wCtFrlvR0/aaRHHUAhyXea1WIl7NKEMTY9cI2myumzhpC4tQhX+k164b1DACI5rR
EiFLDeS58eEtts5F0OeZI+sg8syrDmHW/o73ZO+AoRHhgHHdOu4jMd2o/ZnzhToE
3UVY74UCu1GE1zckLMO1UHCTDSSfPLI7Qxcoi53sIT52H5356uuEZqTyd2eu7oAw
QDkTVSE9Rj7psR70JuQ+EmSQZcXiZt14QWhGjBfjQWdmOTLjICTIv/vWxfH5DJk6
qdTumvU6WxwnISnWjArIb9l2ES4x6TQDQSanUR3ASKJR/FxhNSTJ4mEVnHy6O6Wl
H2mh27GqWA8MU/loafxr2amrSYCdoeSEs/93T5ncbNp6hJmYXHn4FOT/LJx7Y1q3
S0NQnjSkMgjr2YbrdBzTkYtJ01MzU4dBtNKz86FTlJHFERIASq1KRHfGRH4X8OKI
FzmlacuGRPRNpl/87L1lITX0xC8zuZxrstw3aDxKiRzPN1vWGj9e9Ly4LjMizUJ/
6ctLdHHB/4RsSUunMDXIEzpa+vVRNJbfi1LLijf4JAXT5NwRLKy+EKzq1fLrhwpY
tQ8rBRN1/cqocCYTPodtPTFX4eKMNjfeaDeNZ9DgNyi6HPiQ+3qhZO+91K9SM0XD
AAXFBYzrpWBdj0gMZUJQ34R5HNBJtlBStWrrXx6lrOeNjtKvQ6nxf99ba70Ro79F
RI8vDvI5cYXBmM1m4fY+oGC+mUmeNrXG68I7Bh8rGkb9CaGz9pBYH7fq9ZTeRbcR
lSnraUTcBKoxrOd83T64fMNGrESlQGFxBtMBgoLtst1riLsbQJZAVIAsL2I7461u
LSb8/TdJReaa4wJ1HFKCXoH8O37aDWXElFHmFUhlI2ZV4iYUdw8lEsaFQBoV8sBe
MfCKao4aJhv3qmxSJb3yoM9oBRSy2Gt0V/kthk+fTDE2oLtogHq+HQqCl6mZ8/LO
szFGyzKqpwE8g5+JcuLkQForFTLkZf+MnBnZHnrNLbAi3sIezRHNGlkIOTi6wKBk
Ux3q0IrpyhgWWfrV3xpKrOAFp+xl3oPWj3CPzsBOOI/xAo+B22xFuvJYGf+DWodV
QI/yWDO6OCTEveHh6UXXwnXnHLE/shuYujXdAPldBWLf4ZALBQZQGyVGW0bsMAfg
gVZ1hC6RteFMiRR6yOR8EI0ddqW1qiqsKM/nEKcXo/x0AwSYws3IqvmRwDaEGeXu
V9R0DLRyXwWmTOvEQiKTAa+gCtYl+Kp8OFSm1HVpTMb7a9GTjCbmwHYoqzinFXi7
lRS+X3DGgWnK7sT4xXU3kkwMPp2VR33w2ubd0y/P18593+5cK0tFYX3Tvam9zCW2
mTBisSN1ufMACgHFZQ95R/aWyUa7PZKGe41SqwGz2KovZ3mo91F+zZzVKZ+WjQ1C
IxJpVIrSuMA/ssWxnkU+eJVo24M250Fi8h49uYio2u8SAaYSD5Dy8lyfbfPqWwd+
pyQpkWOeOO2GEBQ1SLh1zYL9QCWZgrK1hhV5lrZ+NC2OIeJmEqEtXq9+C+pFzArQ
3LlYcuLqsMNxH715++PY5epi1oxARg4U4yRWTA0sZsJ2I6YQLooRjaxC45cQtmT9
sakXy8GxWSJQluNrYmXD5Qr3IHyrl5tzhdT+5qQh73K6lIDIWsoFH21zKbcOZjzp
pkXlDc2QdRnOCkkUc8Rkso65WmFBTwjMTAwjvyR7jjNUz/yl4Ex3odD56186JnYC
sc0aNFB6ySYFSx0kODhhZMnJTLfvCppDOFdcBPQUqSq9Dnm8s9ZtF7TtvcOmDO5Q
MywCEWP3JR07UD1hO1JMi8A4mYrJ33Exnoar5Tmu1VLrbb4vW8Zuye3mHfXkzAUe
0b+K1H2p2bcKGS77uWOXVJNiVcTtCaQfvvQvWpsOLiir1eWqmOkQnbcTatRRP0aJ
W/L93Ob/TBeJ3iOjEStz/2/l+DXZdUbw9dkgjvlD3+brMCNGM+H1EBv7tA45MexV
EHDFp4/VibzbtFVwgE/WPi2J2O+CoBuUJjSUui7t79es+iBbwSupHtt22CF0afif
Hlz0aZMy7rFjJ4bH4MO2ZQlqi/MC+gtKlU6bISBPfrC/arHj2n21NkAOEIkP1SQw
wZ+G69qTHnJuZOcuSeQYMPcOoNN1eL3wRQvgaBQ8+PhPaD524Iesb+VCI+04xJUH
rGfH04nTZ0H9UMvyr0WVLGMkkNbeZM0l5YDzCMR88jkc8grE752/D+vbbtJKJ/Gq
vUGZ/M83grFIqr7kX3B7EYOeAYjIonYB7xs5A+Cx/mNQt0+gK9LkZUA3aboTID5U
hMaYK2D1mu33vLznp+r08Vla7LUr0P/J+FeexHyfsQfJL93Ot33GRSeiJXZGi7AA
DCgObaEkl/x3swX1cvVuYgvJX6VIOqsKzzvzAMf2487BunIADQN0Ge8VDMAXAGu+
QJfVUq2H2uSZwJ5KRWyD80bVoSDPp7+D3xR9k7wfGUIv9T6vL4C2CJY0oANnkhgU
c20KQ7oCulhtGs1cBAigvFfQLp5HJoMXRCgmRZRtegn2Mp5nhV+xXAUIgsOI8pNE
EzcUxfeoZ1pQJOUn4QRF+U9r6em3dj68d6V3SrcCdaNnem0PWBdkGBNNpF3tEk/+
frlGRWAaLpqiAIW/W1kJuWnnzqGwMZcx4MEsTES601dbCy65T+6FDg3Rq7Xkdsbz
tXzjyu60LK36cfpsxvmEgHCHE4Tbb/Uz2t9ftyIGp7LSM+GZD0bh8Mh3cq1rkTGP
TmG4MqPAc0T5X1Jdqz1QTwApldN3Hu/u1n+PTEs7G603J7LUur3nZj9Dic3aLLpo
luQr28CKE7eplvpFyX1r/6OGw/Z01vY4XsXdMU//mHwqS26FHMZvb0vTIlIuGtrU
+KdSZvcoFXL9pTNhIUfGpBlgkp6mMXm3DbGZJ5u4cI3itBZ5FDrqDFJGRGP8maGS
4zXjymQ+wy/amj7R3pk6ufEhKmH+B4xt6gfuNR99OgAKNqFpXYiX5+SQ1a9NyH6s
nd+Bm2IGTJY7kJ1dnby0v2JRqJwtjowVIyfAgGn10Hi43YRiL1HrhnV6QSvUcSfS
BdQMIjuDsWAuc/hHUaZpgKnUsfBIu0pbmaZMMObZA/aJxLIKhC+gBGevuB8kUXpt
tuqzbbIv8pygSVWE5TcaCN9Xjgv/J8ptF5HsrgyYA1kiwxxrfdrDAtQSCvDzRHtt
L0Emmu/m4PnXkpwug6ziSYmoiXew18/7duCWboyg+U3+b5LpCRkITOTjt3BVwICi
Fuzlq07hOtYF6NbEicZO+imnHqFlhKqmjKIDRYq4Mo03c0p2iCzvos3ldl3YppLO
EJ4bncrCvA1ZrDp136nFubhDXzkTbn+EmjLMw1cXjhU5xF1H9+7eQWoVOkmjiWjs
kDmxYEN8cMMaQv4edvRdKwkb09F5lcOgtl/EpKjbeDCKWVUpPxtSdgdoNxNVf+KL
QUOfzpmpROQOphyR7V6jUc4H0Wyd2ZVQvNZiK7JNlCrMgdg/reg80mGiCJf5HTL+
QvFbOemMfOJ3uPPhq0byZYE4+YnRTCb1rFrn1Ag3bsZGK35fDC+LztB0OUil1opi
WPgAboJhywGLS/Q4t8FJhM+VSMoQrMD+tH8YwUSSobgOlPapFYdse5SYD5g/7Ut/
SJCDKQJ91ZaIBbpM1mZdOK7iapswKQdR4pPr8XcdZRCOyJ6w50AcMgjz0KUOHf+g
rcjFnsvgQMkeRytl31zUdv81JBR2gproRnVC/YMKIxGW6T+I+6tGZFYwagikbhAN
qWNj4sSIJw8kJZM2kpkqRnIx68oPLG/8bkfoxRGTFEINUcjN+d7kTjYqAQ4/A11/
dymOqyIIRjYm+apda5Qk0X/gbtJXd7PDaF3VdrMjyU/EWA4EIt7hTPcvSz4ThCA0
m/SkwJ1A8Loqh2rOjEqSezFtJDp5JYDSiXRYuCeXO1LYGdvMQvVEHgVpT91LJp8Y
TRjptmIUPJPZ41Tgi+OQn+u9+vfS1HpAOMb4g81wfCi8/A8K9QKYzNBHxI7JiBX/
1r4aKbNQHAg1h8S2H9mSaWvQSBPlxzCaeoXtw4Z+AfW3zNKsJ0heMwarqXo45ZS7
JTf+xEosyRvCjZWywLRBXSANk7uTqZG9d4skYZ0So9BEBEmD9snKCBZONjn51eRG
8hSnw3xZahTWJeieA8uUCDaCCnqtbwOu+dcE6XAY0krvY0wtqalOCf9sM6+gJsEU
MkQFk1GAR7CKj+7L+n+sFDGRTeHA6TmDDsjbEIzs1YuPkEGs0177xuUBW7LnLtW4
1FEaVxNAMWbW0tSA3D8wVjJ5ycN8lS76w66qtN8Vhup2ANEJ8LWJyCeMCxbcU/fu
XLZnTdCWA+sRVBks+rN/D3wKea9e+5o/3C0ZKPIrm6ka/QTQMXHxgiVQRok1ENG8
cjIoDqYG/eDjb1lT9Mc5j18D2A38GmwJ1nW+0p/lUhv6bJKT24CV3fOsfJrTFNZq
R8DkTfuDR8rS3QJL4ExGsFC3zECeDMJP++c0kDr5av0gcntxHlEVYPi2bqnUuy60
WgSAT4wG0b3Wkqs8BcjqwRfTNz87QBQ2U4FPy6Zy3qIyZGjhAGvky8F8W8tQ2kYi
h7FagtfB4rwTFlG93V2bSz86XFO8r2qtr2XOYEHBIi9eGFDLipQq3ovmNGpZabfO
ZcMNpgPKkTuaYOQkNHiH4dFXXFdE9d7+OnyzbZZetAyZdw+eUkmjmRgEfANch5aP
IuptSh8V/ywK1FX2Esi5x1R+IpNt8GRH7fERVaRHnp8a0yBb8U82zbry7VJwgxPI
wD7cMrrGsBvZTU36oDk8nkBu7XDv5MDgtuexrag/JinJYKZtNSUP0XpKF2+aGrwj
QpX2d0sRwnNyXiUMqAf7AD1y+TXx1ZnkstXBl5wuwE9p39E+01DErTesa42qYuYH
wRe3jhuitCsI/nNFWkn4VLFkVgjHp9tamVHhbf4CZ06RmSa1TAcESikqV+5qSKGv
8Cq3kLpUh4lm1hReeBbce07PSzw0yupKUP+A+ELjnc5oqzoqAEMO8emKHVzvK9Fx
iDDwJDKCUlJQJQA8Dj9OuYWljftSrzipTkftm/JcmCys+2vOIsUc1BJ16LGlutg9
5WWerWPEXVRen9WseWB+BUe9jjPdX5yn37B/U/N7hdY6EJECxeiniuaMkbxGlFn3
lZg3u4XFc51A8vfR25sKCuVt5Twa0ny2ZYr02SMfOOukLekuOh8x3o8SaN+wYxOK
SxHxI0HkMJ7ouy29ZjzllNg65ZhUmVi+PFIcoGMyPZAH07bJCSrj0zvgI6ZB2u/H
jXNwUVMkgxomm3UMN67Bk7PcLI6bwzlTRygdPucJvUtqg7J0va41o8BoLQDNuHdE
hjupFCkjuYJ0a9/TWwAUiskMOzEclxUXS0kEcgM4h4C9cqI4aEahCZFAtx9HHqFK
DeQQyi4BnKj6y8WCjAidM7PewDtfjL8HNCou2jkRL3isIln1R0v2VUgFPT36PJJt
nfX+HlCm5lOyTdn/sc+VxMmea4Xlb7fYf0LIU7UjqhrhIzz27lw3VoOEwnD5/n2l
CyJzI/4inp3NetkOgZs8jP9xH9w82JT/xdaxH0k9X1i6O0lGy3xcrjXOzTIOT9KA
IlnyqT5RAPLtJ0OSmUC8GIka3LKm/sD2UOf+Ttkge8lvKNcNKnCi1sYZ6/TkuPdk
uY6iR9RI4p8b0THl42pYRP6mSowL4U47Tkw1A0NzNWsQhngJ2UDk8daGRWQ+Li4S
fcphGz94Ip5LdlBKdUNv4t3qa5HssT6U4x6NxQIghzSbteCtOfyX5aHNeF545x9j
+OqE5NxzSQVOZ3k/2Kx1h8kB+65eGsngKUH4obv5g56KKadFQwNpPCKXAS7PUrtT
mQws8ir8f06cFYvncWUTlHfQrKgO1pFPrEvkIoatQ6Frbxigv81Jh5WC+GOo1gDd
y4iaKAJz/BfNnfvhFWc9TW7PRuogO1zgsLIxklSJUJ79qIzIHx5psBoruJSUL+hl
KwVoQJlmUJlfqu0Kp3iT/uJHcjjr2IgLUan3PwsAi3pk4yflLjUXkTKQa5LXm7fA
MYTzvaUIvQ50Lq38XtbbDifx67b2HItDuJBGLPhBn9nCpLQyaencFiYM3hBlG31Y
mnoz8UAqvi74pUcBRjUjRV9XHUZLeI6EAT5dAJbwRtUhqeBx6uy2CnwIsbQ/flE+
i7x5h2dpMtTXJCeQwwD77CYtr/UED68E1HWQSoa9T3ijZfmbP/gBF21yjyZbWU2w
EPI2kqFVD/kdC2qgDSMaj18AddR07viJF1c/mOAPgOMaeyq+yNiKV+jYoW9Mc60u
ucGa8LKBQSdSa64EtkoxoyqOwwxPqD9ICWrSFim+h8yoZ928ZgvJkyll3ngL4iJW
48xVOWOfLOaxHcoZRk+BQmWxqdRq+0DCfejhXrIL7WZ9cWA9y0sQVsj+prV4AnbG
guqmzmaez2JJT6Stq/PK5kY0+704C1n1gzcXVXRajlRtztLdj1dlzM2RIpMWzix5
e9sfzObeN2xxlrcFuTat9wf9PMOutTwwq6q5OTvkwZVQd6M3aWVknnVVNfJ1Zusg
sj4usr3XWN8W27MjkEcVAFCBhV/2GmoYmoENivhySQgqjVsxo1FLei/b5wMachWo
xDpZ8u+zO7w/P0rHYJSPHXWDulCvNCYq95qrno/zhPBo8ta2c+hwW6ILBpBJyQHp
2ku5IQCMJ+AuLgbaHFXSq/clI3uUXCYikOcIYK3fkaWkkfWBnvKBZxZaZXw1/rYn
JeGw09GsD2BYcRhWrEe7QoCCTwQr5iAKhDw0/BBTOH4EJ9K2k2h7o1rZI2dJjY3x
ek6kwrizGwmf8xvGfxBJVaCqaUhRXG3x7HnfrrYzUOoT9JZV7xoKlaotg9Xpa+mR
D7RxPfNHa9Q1yNeLTtNUYiEgoklcf4YbYuIMgTf3D85Z3Ky2f8uo+mGBZm4vSfsV
z5obXyGsNX/yznYtZAeHOFn/kmQd+EVjytoF0rqKXvEHsGEDe4MdUrbMJA7CtszS
4QDrY/vxmo3j5yJcGAgXlNC0UQ/9rc2qWWuA8hqJXa5ESDDLK4nCRITDgxdvQdKl
3kbBOkfG3qp0HJt6rh06PwTI9RhtBB0k+zFjLyKFQj2EODmmOXR7iCpqDl8UG2KX
Gy2Jyq1yl1A8P3wkd1Lg72LhfvMitqKMDbwDdFcWoEtUCxYBAs9IuwDeUPCym8bK
8xm6T0k8gBNvX5ayqtuKQjYHTRER2aeSUPKub//Jzi2y4itkeTAOOZ/4PodpgTD9
BttPCNBYM4rdxjLk9n9W6VzBzSbrX6Yr855rSEtJKSqG6mdes5l5Gqlr4h0IadBC
78MvSttDPdbBL5CDzW3mCxa7AkYNlZJBKzkvCNjhXY7PFT9gH9892ukZtLtHPfVo
/xZzLbbyDF4SbOfjCX27eUP9ajNrXh74gOpvrBiRd7DPDOkEjs6MofRqAPaqzXcK
MeAnP6tJy08iUWKUb3csUIrLlS2gFN4zK76aw7sULO16InTtrSh4s0XOOOjLzmCk
yF4gT/YKM82dvF7O1phUaWDa9OPXCRjmzTGY5ZgwNaWLBM+KXhOVX6LHiGw+rylI
faMEjbdeg6BmZlXMSmLB7vqAO09gWQC0ZI1XWoUsfo8rdPw9MttEzfrRyVSPSajd
v9JuhulWZgYCSjPT7pI7J0+EwGrTvh16fb4VYQk09uufR7+ubL0zI2SDDLVItpOD
gL0xf4OGYwhaemm1hJYttMDGtyrwefzh5xO5JtySRTGsu0sBTcyt94Q9QQHJKWHD
GkfbNsKcFDbUQBgOHNIm+TtVDwFDTyTCNCeexBQ3FnXgkUQlNuHGPo7bk7+KATcA
Z5OvEI75mhhV8wfGIRFYU85q9FEnk57M5bu0ZhrtNntZP1Uk6QyXz9UQSwybfjgK
sVaf/Gac7gdUMKdPrFZowW/B2i4YQgt8NpLiMBPc/n0kz5hyvXmCP51G85UF5XkN
tsTDC9YWjsIscjagSEO6OWEima9mZq7M4+z4SteuErIIVgEmuo1us0urTA44Nuwa
+J8tcBn2rbHdMvOQriWzNQ7shA5y9KjPDz0d7omiYaOJIrNojXHu3KexF2vqU310
ez1NbJCFo1yxwYQi+Niin662Ctw46DeRQqUpkxmyTjZTL64AmAIB1viib+4HLa19
p+Kgl2sf6GbizqxWh0zJpSTdfcWWxfImLpGlcmGnl66EKQjuuLxokw1Qg/tXXGpz
Im1Kj498h+dMdFJ11Yp2IDvS/sZ2tmKcF23zML/8wFkf2tBwcUtWAtszXXlmjo6w
vxFdW3vWYEP0irBvrX2mr2fKnPEJFlCyPuLjNZrb/4FuCzD/nEzhcV11Kh7pNhFz
EFpkiJEmnWlzJ98EJZKV9qE84jkcqTT/UoQg2RE+JWEXrqWOosMubWkDRrBd2LRI
hTNh5pGUdPWwsxLpBixnNxX4S/8TAYc7IuxgFNZtt6Cj83g5GIsms5rDlw0gH/eV
B/xknMpSHp4Kip0N5kcCtnsCvxKqrFXEGIsLSxzBUU3gs+4k087BbWoK4zNKPE/e
8CNNOv5FijC85qmcQdrBvFVnghGMfCV70cg3xHgImFk/7yTy2DyvdiDxO+TApp8k
LxSNziDj9pUBg4wb8jfUkGvPiSyM5JlkXJj8lztdvVYkU0U5W5NvZ98Ee6on5/B5
5nGvhAd5sMPlwMs7nIb4yolAKMxOM/3DatWzRet7Mnou2cvbEZhyvIQhtNCDWDis
oQydKE3nIccdBRA3CC1WoMBdbJ5UGYd4ivDb4o8earWpWYvrQ3OqJpeNHpSxVpMC
m4Y2aybk/QXBOACd/564+zYgtPvgsQh7V2HV2rtT221HA7s9iGxBnUXtu/ZOkDm6
ppQxM7AbkH7U0m9QlFfXQxfm/Zxv6OD4jJf5lHLrAfOPkDpgaECgIeO80XI6ADKe
apfFvvx65B2629I85P3aW9iqHtgR0H16HWgg1JWpRH+Qk4ENfxB+LVjy/A34c2QI
lzVheLaO+JLt+IqlUiyshS0/xr3iv/roGIeVxtGCdaVhAd/Wf1KYfNIbYAwRvOT0
8v3IIfj9fZVUf1BHhPgaAR211qIbXc8Z1HjiFe3ydDORxJ5vdPDSWQ9Isp4AdRGV
YyZBMVBIYQtlDl4m0255VAWoCgG8FfGukfD1XeskpDzqAqBbRkxG0hk5+NdnR2kk
YLgSR38GOVBfpUMRKf8lohZIHF5mvCvFXp4YYD4F58jT51/jPxuMt4qmDF+YPoze
04LGlIsjW/1NEOUzUKegEM0byRe8+o4A++QqT1B6T/uW2H4p4Da4luXPaWbepMJ6
FYnTBf5vLPsEYkZkIMa8eBAm4+PuyvOLsMG5wFSAJ8QOqNAXdFPslHjwwkALXkO6
Hp7e5n+D08edW1dfEX1OjEsIhlcHbVjdFr8FV/8M7+vpjuoCfOExZMhQ5v0fBmQF
D0vp/igkfXcAqIlazrqGSUEMKr0R17+5KCqrTIZPexbVRF4e0xMyJ622+5VZ5rrG
DZ0d9UspXi1lKmyg6W5CEJRVqzFMzBVT9ZwR+iSd+IUzxkD/A8cJB1Vp01ENYOvz
PGndghn+uk5FHgZ6ioa4K59eWYDQuGGlVwWv0PE5cf/fbuhacSWqCAH+f6W7Dah/
9QMeKZNg1uPpEVnkRXt5Ow57DsC9oKE74xWelc5qkVIA0X6Q9Pok1oOnf8z3532G
1BvH117z5OcZTPS4yAhN5O2j5qTYFAfW449bbHVOHLmv3EkyCp5CqTYBQyYNLLDB
9zsG472SbnnT5p1uYlFQbw4fYViTXNrCF4WuuhQy2hZo8r/hCIUMDXiXW/0YlniN
b+Cf9iWo5D0WQayROX/Wk+dWd4+oFWI89E6tbgfkOkLx9D1LWpL2kf/bpT90nwxW
zItH3NDxr0WFHP8FIQYgR2GC4DxutzjgZfJu1vd+Wo1acVacoe2njUK397014Ts9
OmmboJEd2N74fON6Y6QYyoxVv0JxLuZgt6q4iHv9Gensdtn2Pk0HuMs6txlXceYF
jxyTcCF2ONgs2DQ0/v/a0B5g8iqTH8lMvlkiK9qugKitjOaUpdqOxXaO/U9WlGze
F6BA9Kvct5501TaEEFLFEXK8brvQhkU9ZcqrZ46ZFSbF9zUALZCLGnIjeC0wSpoi
GNdlENQGu165Xvz5r/emOk7DQF3P/1kHwcCzENrVAtAri+MDFCMB9Y36EKTzM952
NZag9SQLJnZP390yK08nbJFU4/FvNgSlM2FkZUSxml7oc5Vix8LpEFubNK9+JX4M
IpV0+xKV59aqJeVhJ7d3IGlHh1xLca98uSCkHhli2XZpD5boLcwT87k3jkFl070f
3bhrxGCuhNdSkP0LX0N9CLmdcxKvOU5bNhv0NjDMid1tjdCIi6I0a7Caw4EwXw46
iiSrKDltzw+ZkQ3e2brfI6Ud861FFgJ87s07DoaffMEzvnFt+/xh3fF2hMhymxqp
T5wuiwwz1uSYYORi0w3+111Ked/E22CzP7PImqqurd0eoBDLU/lexzME/FKId/s0
aMymqqTr3Ww8T1GB37S4wnPi+sgtjTkX8jy3zAFxqE8n9UDy5e3w0GHUN+krDG/g
F21Z9FKmC9wkyeYHUHOoipfNI3/irm/yNJn9RHQb3pgdlmRmI9iT1Wga6rh4hbxl
firM9cWJxtijjKkOM8/WWrH+dEkp2KvmXw2vwp875/5XMboa4CQMxyhpXC6sHd72
bExaEPYjmSIxzgKNLm71Z+Sw33mmbb75RgZB2P0MvD5ISQCKW2lIQmdKFYhjjijf
IzFeBscfYzN8dx2mrchMvqbA95HdvSNCQzB814CIoHdfPVz4oqrOlUVsKkVE0iav
X3M5STzjUbGAbpNJEstTe1NjscYYXJ6KVhMqP3VGcoAzxkS/UxiXcrBzRlOMdujo
C5qhLYNi91mHzo7+qTHMZRzKlpLj8zb2BcXiXSrRFwY/rYNgneeasDmVxFaEhaq6
Agt5WST58+3Q39t+bGhQkwBvnGYc1lZPIfWuKgBUYg1Bd8G3c9jM5u9ClDyyA8Et
J+DtDssRnTxMh6J/Sr6dyI2xL9hFq0lp9kZ7vIzPDD5QUhWLn6ui1SFyj9gZEmbI
Hye2qSd5EF55bAO1tvK86Y0AEBU00dP+SMHsBaBAOd8f+BOY6QxRQzMhMcFR19xT
9js6Jx6vR/lna/yX8CgyCZQZfBTo/weOVVyarwicluc5b6nZZGZxOnRa2zo3uS8I
3cg69L/nlQxdifshtvcpBCRPEy9HX9IiznTDHAlXhBU1jkHQmBmmNsD2wvtvk8Ea
CTwyzi0KgeiGpUgT2UgtVDMtX0VvMiPfshpJr68H/eXGF2h7UHOCjQycPREKL36U
Af/StIle+4oRb6qqG1CqEgF6uFwZ7Re60m8hKqvVLJUn0Ajt3da7CnyjoIbMZQ8x
ZMdl1NzkEIHC4ceWJ5b9OmTgz1mL8NqVSYEEoRLP8f+2R1hHCv6mIgmE9+OHGatt
vnR86tMiejJpwxuN2zcpx4styTR6W1E02+A496/05jt0Tupmyk/1klPxt6IhRW/b
kFQARIgWDpAQAQdVa+tRxQIw65HkhnnIpWutWXcsM7NPlrdoga8oLNyJky5Jc3he
Qq0XtHTqwCTxUuuTDSS9Do/OEZxSuWtDYXGiYUmu/af8EFAB7Ur8mnCJJU/IHEiD
1Auvs3TQEdS1dt7hQZ5xQs+qseGvgPgwTb9qyRfN1FXAd9tIQvmdE/0Rz7wy14Jg
48SCikm2eVNGTt1S4WAJAzSMOuO/1y5nZK1xTBdfmCOywPJdFrDC55Bs4SRx4kcK
x9jxMl9Y1hIB9kbrUZR/YlvhqyuPaZa/iQFgoboWTQ5WwrFJORm3nVDSJlujam1f
VVQAAUlAJEB8K/DgwnOoqajGwHr6Rj/tTy/Yl3nRkO3rzCslqKlnJPGTZ908Py4f
GW6XB1jxivzyiBE88RvGfseXN0gvq0Js54PQNGtPpYqsg2nilOfDcjmeiZEIVq8e
4N+utmLiPZZY0iorN6ppZJH+J4mGW8zuQepXdpj16YT1kX7a0XQ5mGJKu1lhG1l0
x/4KG0ICMOehuwINa8LnOP7S6BQV0rBhA5ZaXofSNnofV/j7VSHbWoPo9dV2yEpQ
oi8F+gNSYC4+TMQnzcC1uhuM8T0I8GYJWuRafNpxzxJWqgOEMyAGHP/g6fhBgLDj
Z8gm84ejC+WpG6k71wpqeVt68o9SOrb8UiwFET6PhmdcKBFTjFi7PlY6ZpconBde
lIJVzBPDr5Yrk335qRKVTHC/IZqAiuwhSk4vU43Kp7e/RjyfXuDR9sGcy5+qc607
EC659sbVoJ9oZD5KLts53vag4rFuMYW/qz7qN+SV/GdNhHozPpQwRRdWOaLp7dmm
tF2QuVD37geTffUeqLhx9Gq4eBzvr1dEKY7nmN2VJHzOuzuVwA/j02Jm0BXeLOxh
YPzF4euXslhgUkTR8JLHPwWOe7SQCq29Sywq23tIgnkZa1r2kj0HugEwY1S0tkND
SRYC7uF0FSEO/9UgOGG1rJWYyhKhmG6GQjR54g+Uzk26PRzSRWdCpMcVd3OoNKCT
WWLi93pQgeEj9udu3sdGBh2oqNXY1iF1cnaJq96tNykxkIn94h3hl6Ns6PnFAAOh
dKXz6DLY+Bc/UHDPWSjwpRhyoTn7VPLHbuT/RSCNDaL3HyzIF+6CZXBYsX9cTHAk
ZYmMmkcM+I6TfoUCDUD0IwNDRVnnscEKL66uVxGyOVOYmd16Gy7JZJNbUcqjL35a
GlgPAkgezc7yADaN35ZSJJeQ/0mmvnBHWCaelzz/8cDd7Hr0MWW1kQwFb19AvkKg
kADW00VWM2aeixqvHAcAFYXuphNc0LdvkOyBIToIpH6j1V+aUPHJQyik3y5pt3lS
bVp6BNY9QOxRKkuAZJuwD23loDoEnNXUvTOBHrD82MxA2oRADA8bnz3yaw+e9Dvh
eDgCfQEqY/kOP8s1IRTAMTdcyn5+duhSn3RQ1mvzeuL0a7qle5Orz12YzJiyw2Am
aBEpxCWWqH2REaA1ChXlWrz5Grj9fuipoqfOPaMOYFbBA4xDzooSK2DVhj2EFnUT
6jbGpXYNfyDczrg6XKB/Fat1bcN+nxysnQ5Oy+a16G2k3TDLSv/MbfXlyU2mOEZa
eo0juBxGOzNRsfXw6m6Lj9EGRr+817q5JCfCuwmGFDb6lkH7eazPvZwlVt16BQO2
gjEXd7uC8a6qTLtk0Q2enygRMbtvgWxA9AI92EhdvF/KL1Y2lWsTshqQ2j4YWDWy
RzjJIL7Jh8GlvbDU9SaqtFuC0m0ZGkQI6XE8XjxK7jwv6+hV+xyFgf0RHKAEueaF
xpgH12tw4Dsj5W6oTKc8HfxrixED2AnAn9u0PedAnrpUrZ8ajwYTtG5K2BgHqYEn
sjUEZTdjmOiILOygetgBMuxuMDL6djaxqfzReOvJb5zNCUcgqNNP+eYKDP1GTKdw
mIJS/PDf+tjq8+O5Vuw+r5J9dewQjfx6RKy9mXde/Nu0H0CU8GfWf78+0BlSO9go
Av+J7No5v1fY4iVbHHm0ujlO/zsMCriomAoem+1NBneFbOCJ5WozkpoP4kY5/eln
TtNjgwM7ozqT/ocFTvxMzsm+RhQ08Y5JNQXfiV1ToeOIMpzxB4tHLLepSQVZoJLm
NSbNrH41VMy8ouuZYHLiLUM73Skbvz29hrDpaGmGkMQgE91G20CD33m4/kgnRsQF
IYkuTRHX9sUmUCVC356dZVnvSbfqb6coCd27u9/Amx7VQzoXMAp+5SlX9ixcVkUk
p8tLdbkPMwvqEsYJgKxeLJMurFF/Uq77uwCgQfdrjhS48ycx5daJn8ZjY00U/wWZ
yVkB9qoOXkmm4Ls6h6gGZMQxFhFoBIPNA62rVIUNSFLQjh1j2oo5PDXw9xWW90J5
KfzA3HeAmI+ElCJp+p8faAplVxU0nKFw0ZqkEzhOljcU2W2S0pHUx6AiyiJKxgDA
W1I2goPcLKzFUFaliOhX5TOKSLUVUz9O9OJQOakWLSYV+Lu+Al/OkB+Vh0Ld/teU
jN+Crvhx7K30VioUnJB9x4fqYWHQlesyBSw2bqAUCAX2NC8XJufwW/6fLjT5wvhJ
7/GZRhKBowI0ScMSQ1dix/H7EI1miyWHpWHhoF6wzSJ4g7PP+HMbNkMnyUvHOVpC
KlXfZrtFjGRzOimPbBasWXXHA1GSB9a7TDiwS1NzXsq6+enqIXpeQ9jb2HjbBgNL
ozte/TXgjwr0wC6NGuBTQsLPZQ1QYaF5h/TUeD2LjqOODzwrAweGrklcGU7xxpLT
n3oW4Hx7XXsuy+QiAFkdDVRMVeaPPYNTflGyyrWMf83MmwUOCVW13u0b0asQz/LZ
/W3SVEUtFJ4o7DeOcLDlXuibkjD4GmqzdY/Ja0J03ad5y1wEXESO5lrDr6gPoU49
6F0qjxjnpwBgGYUrLsD7GHT/nd5GiozOvq/CwTS5AS82cQLKgN8EmKoPToOQXrgh
ZOWrCe8h+CD3/TglVnXbUBbfxzbFqAU9vbYWiVH27aORymFxWIUiGLy6BbI0/eTp
AZIy9LB99zCp5eXs3I/t4Dn2t8e67jcfeGbPZA4c3HfXt28K6P+Z81fPvXosl/rG
ppwLCa369/+n4v7aCVS+nHizzupVTfQJUbISgBmfh8zhxsErOMJG4/YTBvTYDZx+
iHI8NNaAa6SLkJtem0LiiY0sHztnGKtMbMF5UPNbn/mDRJ/V+8DQpPizJsfKz3xh
Xh48KgqsYIdhL3k0Gsun+2aa12mVTHp6tFvGeQ0sJLWmwewPPCO9QCZ3EWqQAR6+
myiBzqwW9tjDgyYs7PHza6QxBcJ36x9DefmdpT6NWnc6F0fsOvzXFFGrce1+O/V2
fryu6wYSiFOLOqoMgpBcn4RXnYPSN2Qkyh3nTAt3joMmtywF9QeH9eZLpm6yiuzt
0wWhjZUXUnxkksjaf8uhJxKnmRD56mviGBP0ytYyFAHk253nLp310fy+EGbkkGfV
0GlEApEALnkUR5CQwAq9hufujNvaF0vuwwKSINbNEg/bGsp/asHPJs8q1OulhEoN
0Fwvy+RXzRu7ncyEp1odz6ovRDJFLbkNW3pDq6a0femjursrXVH7Td63IlYEyJph
5kkU+pu/bzbF2xwdgEakGCMYac1Esu91fN3N6BbEK27lihuN2nsEiYhIbO4eW+jM
BGgR1NbR3uRmFMDc9zeCGIeBQ7C9VP97LcHywQZcft+7awvqldIqVkBG9zs2rB2S
pKoaKPSIo3Gpy6cWSbFo1wjFOLy1YL+tS3M8HFmQJ+J5n/jJuYoL9J3dV+KAZrmV
NF/Fzg4cAkVZ0E+DdxzuVZflnxkOQ8WFi3+BKYlTVm1bzE3ZBsvztoQ9SLKNPwGr
lxjv53yJotQFA67TatiNhrZrqAmhb55c1QLAqt9besCANAEtW92x6CaKyn376Vnw
yEVWn5mgTnU5L5EOo98xHYZQlohZza3AhE9Pao2O58yzCRb0iHsMg0W0QM6xvoWE
HV4uazWz7nJm2z6+B4Umdx+FOU0mrAUaFmHCZG5146hvgngsAhfXXkfTe/E2JBGq
GIKk7FhWPiLaQnFfyiicNU8vYB5pAPAh1du7dZ0EFybsSMYI2DAovK1YzhLh5ra0
L1Qa8kwXKFccZlJYJ2+BPhtjFw3bsfmrUgcA1zTo8FTtBae189JorxLW3hDpJ0kP
EMpoFcxjQ/9cUsmFhLYDT67a7XPYc230ccnEjmXd6nuHPRSH759jigVrUDY04paU
Gs+dPVApRhsWSEtNxATdbSqSL56QN+r9g/outxhiUAC38oX35eqyJhjeI5A2Zw0/
klvTGIbzzkGUP3BdXqZhm7HzyRZQfyQX0g9fftuuTWfZnjW8xdjlvClUOpEnODAM
KwWtMe1yICNewZQLWgzv+TPni40JPWemGgJEYZ/fGpWRopys//lAwUfsiefJUpb+
QvF4yoHuG03SPAEKSZGLdxDFkRkaoDeZMMtKpyksIBw8Am0+aHmQXiRa3xnH6+S7
EuRUiHOlX+CBOce0/c7yS3QB8ZB2SVzPm6OUsRAv9GLaXlGKPQSkfXItLuJEWoSO
H7xD+isXg1dhNPw858cVwxD+k9I9A5sb2kRUF/Frw7dhBnjWkZGtDaOIUIFE7err
azG36N4Iry+QrgNx0EvwBMqmtWrKlzKwT7a8mqh5gjgqYcsd8s7wBnLGrvKAEwWT
Pn0DiUVGYnNkNXtfd9H5+PM1NL2oqfJZOppUCkI9HAbSYxj7eQXvpOF8mPuKi49l
/PVztvfNk34M/Y17HzRwO/iL2q66z4+kRpNLGeQMmVKWV/EIoahXnNnm3xA34Q1G
THF1USmlu1KQaXHX3un+0X+8Z5zbMR/3Vn5CsAqrK0w4yg3O3Mfmd9RR8p+SlQRM
m2dGt1FE/YCM8KDEKauq2oIpLKfMvS9fcIyZhHqVoKpGXBMV9R6RTWGidY47sQqp
iTIi4MCDND538blsJtkMXqKDogXkiAgCEiCBIFHdhMxlOXmmbpTr8WQDJzPkyUtc
0dxc/q2OnXE2Tq03H5DgGEr2SyLeFOLqoduFwYtDyqvY2AKj7x/UpPtYydcNQvgI
8bIKNFAT4N94FqIlyfMOyf5yNVwbmadFXF2FHR61VtCksJW2NDvgoBTzQ1JcqmVQ
2yrwo8nuTqkjWBdj9ucoe1YDkPY4BJMhRz4Fpkp2shmN+pJknIrRGgJkUUACUx32
s2Y3BlWXi3Ql3psU0P0hbhBEoDCSv6D/ZiX+HX8RouLxW7Bwt5uRy5fFIHlDkJqj
Xwgye9pse9EGa1cvaUUKO5T9JS17jw+FeFZ0c2FiSB146updAVMzBcXn7idLDwsJ
VeIUY0u8GqP0RmpRA+X1zBy8p03kxeXp+pwAkq9visRyt9Ir0GS7+hHmr/O1ej2l
v+/JZ6Bzg7rCmThX38fVI0pUsWxj3tIo84jsuP3rUo+k7GFua1FJ1T2OcA3OOK8G
MyivHzhRgJZLFdAl344w0bG5+PRWH6v4yAFFZ/MAo0536WN/knNYglEWZiFTULew
MSBBiOOEvUeai2SsT1C6guzwyb/MeiVmWZe4QUsqKITpbtp97jdWVbqxW0LG/lpI
rG4HeWC/u5ZutE6eTNKuwaHz2y7egO4pzCqKVWAOwMr3lIVCPCmO8TfAjXJt17RQ
8eA1bp2gNAH7m6DzpTo2Md9P2+SriQ0rQgRBpSuGqnTLPVjW58qXe++Z0Nlq61jB
LghPMZZHM+yEYZDfET3G9X03u3zwnQs0YRNTZLcguITGez3z7zl3dqcMwOIqlFp4
OKVBYgOwaTk75FcikEGzEO7Lkp9CGE514dp52zR/LtuNZNpQFv+HtkisYvKm06qN
Pusvk9q3H1kqxPdKgPfTIVaUUaec+um+ZKAMitdPyNL2900qWAXbVDi9lq7lUcTp
fa+jVwlHJZ51RDm2DQvKsVRuhUoCP7I2SYCyRH88CrdHXa1dzjekIXqirHIP2j7e
2imQEqenkzQLv5okt74MLeYXZBCc4HffGrleonI2EaMoPyGD0KIvgJ4nBY6461Tf
oDFvssUkr2t1NbqgZOlan+sHo8OupkKMSo0k72fbSk/n2qOsS7iTB0mBcAwbr7uO
0cfJp2ly1ri3Mxz3xBZEvnM0Wq6h83WioE5K3vX4eoURKngD91Xv3i/Vt1YX7+Wu
cdhLiOwzsQWu7NIG1PrpGyxe4aoklQAq1MaEFwnrnui8OfXMstcgkJ+FvcqNWEy1
xiQO8Ln3/fvZnzHj5GXfAj29jMz5M2NDElneQleFPRBz4/sxhwRYkQSGeop09zGv
1m9i2mkNeVQfYTK6Wq2QP+4Y9w5PbC1HY8dvXghavsahFhmOL4+OumJdwSz+MZzd
snovSfIEPpEwgw8+s3kQ15bNqMVYyCwJbZKplQAr0oK5ZTqaj+AiWmw/9WMwwbyV
tL39ekOjaTy7B0KAGtuJMzfjPMssBcQuWO75ez1KwC0uV9IbO4Ha+1S1u/BPxefZ
iLLofjK+T88Y9gLoDhPz8QRPOlS4YL0JTyxCZUZz1sekeh9406DWLK4iGtJFWef3
eqwHDPZY/gYiQP9EMViy5PKEPR+60JAkafdQFV+JXRTlLZpAjvLofwkx05MFmPJl
1k9SW3WhG0WmPqN7sEODajgMGPus1ZEcVRIlV1lFZw7skxZoUE5Y2pcvDczByjTV
tv7nJFqJwSIpwdWz22C5XKkPOVE8vG2z7ci5IiXClPHZQldpRR12mQGzE2VqOy/H
UKqYqfbcA7SoRazKSEVKHpqSt6kw2BbX2GlTlM3bvU5rmdMbmzQXRcCKvgtbs0ZZ
YiGxfrGYmFoyMxvfuNQSS4qLRidyOAx23ZfGwv2jlwEmIa8pMT/j0fYwkBZC7k0B
QYiCOZMZqC+6BewzdnbGRaNLrVwpt17zFUc0sIyqM9e1od8nJ9LNAmElIHrpvdd6
wt23yWxbyGH6StxH7PkpM41G3ulvvBA85aXqwsF6HGih5DNrQl/qXyQac97hq8qG
rTAjKYHYdfvMvw7oY5O5kewV9kKcWE5KvORtAD3Oi8ussRAHnafQw9OK06DIGj0o
wADGcGDB80tgg2ZDKR/KAHtIbeOYJDyjjKU/+S9/KLMzI383q5oP/gEhTZwc45Hc
Rwzu7KTAIAVyE9qDmL9pczO7SjrmoP2tjX5mMOzTWC8IOiM5340z9yt0B1GX0+/E
MsmLVlhmPXEohUWrPqo9kx8IWwmuDf6HlI0v1m07GVFoOfz3Htnj5fLYl+zSf91v
4Kx79aJdXEbppJYWVoTaInY2N1fyZ/DSHxA/yaace2Zc7MRJnJuWdvSKc7bhhMnf
QFLEKHLwP3gPr8wCof+aEFE7TUgHjzWn63iz1K2EO+s2qOg+znHBWf/lSGF/fWhA
oMB8oGfD3/9MqT2OYp/92vtC8jokZWiGoO3+7/kQUev6e8d46uLzSrCKAmmsisUh
0dcN/lB3cLPTFNBnmZQ3AGOdo8iCZd8NBTlHHUM0Frr0vZrTU47AyuXgf2vB4buB
+Q1wJnDQctoQFLygcmGSp4M/pVSZbRhTn+6pHlWIV7a+NpIxQcuhg+hn1H14xKRh
EF0+bFORBmWSw9qrqTSEeXbm4YIC7uw1kcHLw0jShyjxS64FSggeMl3x3uCf5MC9
4bBiKAnJ3qLmK0FWJQeXrde2e4+IupHjfHdyiJwenomEF7miPE94jqJw4bK+R2Ga
3HyVxvu40jtWsNTnMOSOV5lUI9b4nb6kcI6NJEupBskp1E4wwU+vnz3USQWQiz45
zgK8GiQR5PJn36iFeYbxGBSPsuiH/24ry49jnqp2vm53KNg3+T2ayv9eyTX/js9Z
WK3DrIlh9ueETDeZDcZE9nOaKdYxRVhRWHjj0JO21eQVFpYMnn9Xhr5bxWePFIAH
Etxh1/7eQbl+x9bHXM05lDZAGhqV/IPq1E2LOjJhC4QY9nOL5MWSQvIp40MxmMP/
kPeY85URigh92WPrcGtyzrrWkD4oI978W0EhW6ijTHtSr9buB5eruqTRgkxWOyaz
lPRaZxs+SQ7C6KLlacmoWrfWjV4Bz+qz72ZMNlxzyEueKe2CngWcBWnRUcObSs7s
/8TRx3/FPdeveoPrOK40+hXUB6es8970oOgvwg58qsOJrYhIa3D3HPRwmTvIR/Zn
O7S7Y8Fb1bm2w0Ijo0CbYeNWJx1qs/HknA5c54CHYXHvuiLSb8V0KJYdJTmqJaMk
msYDs1kZsk/J77fKNkM2hbKevWow28EcwsJSe3eWYHxgXpgLyMfJs9/iNXIFPV3i
gDPUKFka3VvsXlYz2HKi0ETz/cwoGD9OK91VeFtN7SHaEqyPf1jQHRH8/SWO4ecc
YA0N9IiWDzobLomiUE6vhMFUqHhTc6xt4+jASRMcYHlJR2Y0xVIigTN+Nt2TG6SO
kfK4w++ZcBDKLAuxXRu1oE2Ycgruod8bfP3VCrFnOn1n4DJqNRPPbKrTnu7RgOkj
sQC5rxMSQO0nAkGLASzKmPrQVQGwyHABtPWtxFjhFZpQrvNpU/Q/Lgps5aSRPBFw
z5TeVYIXCNy0KVWaeSQedFcfWjwIHqAvEDQNW/v0LXFkmF6gppFjZvgM8nsRlefv
2Ldjvh4+s2RGigKlDwcanaAsBTExiAczG1ENdWphiDKgS3eKPAk4bD9K15jfA0dT
FlFq6iF8U7C1zerqkzcQXOZ1p3DSlCRkqr4xGrneK6o0Mf/tQGFlCnDQEINg7x1H
q7nuMCb7h2g/e0tGq/unwYN891tKx7pWteYEwoSoaoa8iIKvN5MkWhR5IgCSVL1y
Yz4Z4A/pgvAgPZ+/hxUIEiFHSg77IfELY5W1j+pSF+qX1hUrz3Oma1nxaeqM/JqI
wC4JyEMNFNY0HznldgNbakgtRoy71/TBeWVLpNzGOSbKbT2tiQBRW3ujZ7D9z3iL
0nAXokq3Vfg7+3gp9wrWWmW1kV9RpcRUrgDCsv59Mqxb5hGE2/V8dEAulxD+M5Ms
8arAio2RtCIdZeVnPutOirxsOEKvXnw4TSw+7TM0aNGBp8F1TULm5aD/mzHF8vpx
wkRtLY8cp4qUPstQSxZxLqb1tkIPohC2J1qB5T25I5yPdc54xKytz1+tJdNh3SSN
VqBQ4UVjTFkH9Mcceb0zrTExeKGmuG7yrBZ9k3gaIjznv0yWT/wsasIQyWFBTMeU
JGA9RcNBEaZ7rAXgr+h+EOg5fj+F7IIic9dh+T+hZHiH1V6A02EJjhRPeB5W2B4V
Ldd82c/qUnoOJ7dT4Wf4St0Hkt3WD8jlBMx9VbyzQnZyubXlgXUyLX6OC9aeS7Nu
kNFSeK8BuPFLXvr8TlYYaIG4XUBsX53RSO6pe5/ATNnIU6+IR4Iy4WGfvzApW0S2
ncof5HY6upTD0SNrW2TEp8mbWOMSLu0iDGsUtm8z09kLCfB40lzVmzTEVMYkiGWl
32Q1yaf79OtMiN0gNQgEprgn/XGTAtCyeKab3AxToKOsx4HkNT25xT4DBvmIBR9A
+KUJ+3foTyqa6oDM1l8KDBBKmRFcSiA526c1wOg+hkNna67GNWOcKIzh/o2/uIL5
ALYHcFfMCDxSKWHFjCJWRIuhoRvuniaiVP0zoxCwPbwYGo/gmDbCR1MiACQrRJyt
0jDPM7KzFwQaAOqqxUTnZ/x4fKxwer5WVyW9OE76FMXWcI4Qyx5wyGLA5JHApsBU
+lY+DDViCg6yMl5G5PYZ6GSfHLt3Z0ZKOgj+ikAFtl1kNzTshGM4qQY075/51i48
oWK6sCCgaY07LMrTTrUzJZXuER766u2uQm1UcZmiYkfkxOAl13tdXNYIRVrlfB6P
6o+CswylcTsGRRLCN5vvrncXiLED3iGvqHO021akHof32sQCykWP4Nz/iQQtVud0
QSeMEmLP7Jua4n7ZOs1jsHope6V0L4zK0DowWBsJwurlh/doMSW21kRGH4T7dj5N
o9nXqqO8EDhA8FdWBAURJiOzuM7hEFV12UekIlMdDI4ogvmP5opuVaacI8hZ3I60
irxWpWc4PNfEnoBCVQm1ZyhMEjs9vrbzktsxIPyM8UMRraGLIGbs17FIMNHfHD3e
Ie+EtL5DGC4M810M5tuZjdwwsn9SVpqz+KX/mgVE5sjLaRu4aupxsPbTeRecmyQw
l7aXkJcmyXX/izCdDAyjUwxRRsdZqHaTvPTzimZmLBdmHIeV4zcoyNl2uM8kTBUI
Qd1BftPz4PQXd8Qt14y9cDkfCDD0MtyXXoDM+zOPObIcrK325j/0x0H7fhEoUBrq
dIPAoQIWfXaXuEeHPqRzakby1bdcswexTxBLTIGKo3e2ioBk3zi74Q6kjoBW2FpB
BWEZcMis87tUgo9sEV1Ecd+AYyGg7zDIeWtdyr9sAaCKVWja1V8NEeKtcH989W2x
3/uEQwVsHC2xz+kddUSF2H+Ht57j+AfrP/iE/LDMO+47xlUV2hCaRhXTLzCVqIcM
OsJ++jL0RZi0j+o9LTH/2NbBRaFBXCRQybj9UhbxjB++RQVcEMP25PTImyDG/0Oa
PQ5pOSHzGuJnKMV4NtBAZvesjtJFckmDVxRi4dVbJjYkn/NEtplJLBDLdCyzulbg
d2IezEz6Q/vhY5j4V4i8yZ6V/ep4vqHJ8OoqFJrIMzbpft/KUL+a8so7j5CcIa4G
38betZ7mYmEqRSZg/AVWCwigVww97stplBLZMkeqlrhXriTGmyklZQL8XFDJ73Es
IKJPxoGOMa1eNXc3Fodxx5tJwbOAa/31WamHoRr4pm0n7bWjXG0v2J7hsTKvfAPe
RAzYye3d9P7uFo/ZFcVsO2kqI81252tT4i/R3nauvstQcE3wa6ahB6G5eO16+YaC
oPKiv9TE45NKuk4RMs6F02PjTXSE0LJp/Ih9/PujTYDkHg6EyPbQY6LyuZnMvrDx
XWR/4I1tNd8AlmvjAxq4jh+7x8iKswEhJqMxNfQO0/U3a2Aj7xEp+bzYNTYuWwMw
6KDuAEr7tl7vpWl95Kah2/HevEiPqLfwp9v5u3/pW6CdwNblg0hjEhq0suRzBJwR
A8GzC/8wNXQiUjyl1538DWgKqxhep7+t8JIBmqMQ+QpHbejv3w6OG+ZR65bL1bBb
vAI65GQJSVCG03Omdy869TkyChCglraa3U+6HkG9kXkLTantX/hYHQ4I/jVpMaN7
jY1FROLW9YdrtlpRZEgDX0asQKCqRwN1nemMaT3erZ3qxN6rd3V6svCedvFablkl
M853Km4HZYX5eLSSLnyMnkjNSeRc1DT7uGruhEYjjb0s1CP02LABirlVM6cTxQYd
JDqKbpxVyPq9m5FZ4utNoC9gdEedGvp27wPuC8h6pMtcRPqFIu9KWGZ1/meutA+6
06up7+gQNbRWOi5BEvh+0VMwg1w7ZOG8EXPEig5guRBsMau9m5S5jDZ8OzDupp5Y
bxQp2EWO/gJ22dW4yqC6PpoiMYJjPyoo//TRTTELdDCEawBZ262W26mAnBQeq2qL
/PKNDyKGA/dKauyYT4D+v+EIPfSm092E2ZVsiDa7A6O+KClueSwSmAjn+0GFMcnO
jexQc2UUpRZMb0N3+9Jj++ldlTUzA0E8sMRyQsuCaN4E1iLSNPM7w7PXsdYUV67j
wKTa2WWnOxETsI/ytfv/2IZjPpKjLnECW9RDjaB9mTdqfRkj2G1dxqC1ePd2P0ya
rY189oVLnMiW3C5GRwoG+edIgOrmuT36Czszntm5aJQ2x+CQ443xyj5ds/FNzKuu
cAOFKFQ9XodQclvbjTKErf5x08WUFzILiiKyeW5pa/wnDy/VNbWmKj9IiHIjOov3
wQE2qMJOvgyUnNoPRtfA2UI/gTOu07AtrmBizRJRbmC6WawkXT/ccfhzQIf1eNB9
AsPsNLE71NpFfY44/X6+3P1uwZVRsIg0Twqlds3slUAWekPZgjtaH9D7e4YMbMsZ
b/CInL3iGN89FcjebIK/TwJaV0pw9+jERElKIjXi9vrciWN+LeOHIgtlJvTEfOJ8
8bR7MpTGDyyTWwTD1PMK+d3f7FJ+1Oev+NZmQ6HPuBH5SWyyLtsMiv4TZVwAAguO
5jEsQ/cS4nZzLOnYfT0+9i9bcQT06VcYvTGUuY5u9CjM/ND94BGr6XuflK/4KCm0
oD5ZfBUW07jztzPAePK9kJn7mgul05xIHFnhibC5Rk+13YmY3knCjh+9dxZd79G+
Je7c2bll+ba0e/DIjz4LlsntrxmEtu3/C6PVL4Ts2awJiIn2PX5T0TO/ZuaIMLXl
xF0xGJY8RldyIREt1Oo+RONwarIgZDQISOJOEBRUfXL1m14mA0OqpULPITTnMjaK
iGz+zbl5IKbsz5vDyE5Fxtf4pTOQMVLMyKpR2+S9AtHUOVn11+6k4EtrvcY1v5j1
w6EMQD6qMGmMyYXW/mrj9b+mC0CcQDXeEtDPY0rmJeWMEtwX6Zw+DmkkMrZXfg6f
+pip1sss63qN1MQWt/eJuW+ZMntmtMpkrofvEFKacpu7N0dyEv+vR+9v3EavLSl0
+qdHAVXHqPu3kN7l+VjA9jCThuI2DMLv9FvxrlT3AdIqyFRb5KzLwfpfRb3n/ENK
suepEd9l7lgQ43ByQIjjyv1F+ICbOrEw65OhAwnOF7tRpZcAKJCuQ5x6gY+f0EVs
0RyKE04orUFQEL9y4wO2SDNRudpUlrtj0aoxyxjGIwMRUGvkw3Z4lknQh02lhSVz
eBjIREmyOkVQJVPYjW6PwZi6TFpGwjYBooPJd2xVtAKkap/g86RZTEVTTEExrzFk
Dwp9xa/lrwY7FTjKblqwSW/wg4RRoTvqGGgUIYaql622zmj4Dfb/fx/OkPfVCT8k
fD3YJXFgVvh5kMHGWCrhWwaRLPf1H1JfPRYM6+kEdEo8aH6OwpcxQPdk/NAK/Fm0
3vkuwsv1lsyQXiCT0KxSL3zYGkNwhcaPhrsZSn/FGRocWP2Ekgz4tIvLfc/YxLa/
y48gjoKaxaqst9G4ASn4a5K7Piwb4eeHvuKztOZ2CKwxvpqmbj6uW1ijZk+eklrH
vpi1B+y8r3I4akRf/WG3ATShBXdEYesAKw7OPo8qsiAlua5kPddhoGfA1CKzgXFf
Z93joQZH6mGMXwoBHUioF+li/SJbJhGaxMcBcgiL4Lf274OP8GcKmg9x0Xj0bKdV
XH1jjJXellxZNTfJZ/ph1adOGELQGxvb7awGyBBSFlRvMQIftY9brdjmPFHsfzct
I6VwnhcgJ5VF/blUo3mHikZa535DiRLDoZ5iCyMyFuP/7x3LaJIZKYdkNJzTSa8x
KhJVlWylbnLr6ikA3+JX32hWwrMiryL/PwsynhZbm7UUN8IPhVhcR7kQ/R9ozsrN
o5muxHKLcRY0fzHTSxzFetZcqkNwGrm/58g4pqDhuFYTtYjiXb05Qzfwzn+Kf+5a
rzyyeEfOVrzB4tBLQ3tEwFguMFn+it9eZnoZPwfyOfIeJnxAEBtiZ4P4o1PSKrFG
uVD7OarUmyJbKE+qgOjr6aaF5MGGdGrBabNgM8Hbs1THzB742FoH2+w8GbCkN/k6
ATJvuTAwSIGOdizUY4hRdNpDk4mwSMB6C0By5vwqGuX3W8LvDINq9WZE0EL78u8E
4eJEovJQQL40QnmY4596hE5uKPufPpAF0KNibGX288YJ59SSp3j/dxxl8k45HmIz
z+YnW2FOyHpbH6ZMTY7MpkNrS40u93sfpSB9k/nZDpM66+HjMJNpnN3FmLVViOnT
LhsdpwnSv8cQFMNKKU/FZvAn7UvAcAxNUAxtGyQaxku7ldlP+GcIqaxzd+DG7ZTv
m+mORkRRBOk7mr4hFj6OogHxh12oyjNeFjtiogCjyXz5JIEvNJdyA/hVU3GNvpMC
eXZ3VVqVWx0VDHu1JGdwIUAPv4OqQUpsf04jhqhxfsC8dJjbCXH5X4r+qjyfwYS3
0Yi08rwWxY7Zm7m4W0CsrZArqpaQzhoJIbDJm1NS6YOP2Z2HwAQGHnfy26gtZ8QX
HslAqXponxQbeVQ6p/YTIx8u1qzjlfdFOdD6fPkNrIprRnAeBYRaSu//LTLPgldx
iedjRf1YyzIDBQ97fu7Hn4C6Kd0QpHEroBn3+o/7n8xcgW97BIiy/HUm/N/vCuat
9FJMD7ZfW73wAbjrkkGfnzgtwKhoDzVnRVDbTEjJ0V+dJAt7V/LrTDjlTiDndDI5
ZDNvA0Z/76MPQE0CfxNy3WCnvsEY9pSVC6MG3KYc7WCUr5wq4Wwgnf6ELX8LYxLJ
Sluvk/EBsQVG7GgJoCFBZ9iQacbzSdIJTYjgqS7xNafrCrpdaOqe4eX14a72dCpy
//kvmUgT5OEwOb+9gOBVEnGeEELt9yxGqh6LgJmMFrYI4ORguoDE3FqLm5B44QOq
xws12kgL1AthDHeqKv5WxJs58O9tvp7cUuGAcJgnM/SMM193KPcH+8CyMgizClFs
sq0IMWfp+2FEGH4mN3IiVMi5laKzbCSumgbZwzRQcUOTGra9NU8M7firybtUYXND
thSkVeRR72hJAYEaBXRxBN73wvYENLLKA18l0+IdGcBhqM1xnVBRbzX73S+WDrHy
kt8qyuAu5LqYfii9rA7Tj0G/ucFKHrB35VTyIG5asDyoSkqVikpS5K4NI0uSk+1X
YjqHJIz4rPThlO0RYa/0aZSOGqcGe+KfiiOqmAODCWWhLEwKUWeqwR7OMFeb+XoG
JfuawDDcnYjioRHvsV99gwYdr540LH011ZH0JQIKk4Ie51SppqvGYAOtSKuoB5+s
TGUIXSj0pbo/z98iAhvx/nvdSu3zG2hylxAzfsGimHL3xeES6P/e40jjJBZTwKoA
SAuXcQMHRieOJQWdru5c63McTIQ1/gC4e/qdbX0k6jVA3B9VYomdKV9i1YMu24TS
PQous7M7qRN4kWq8XUzFmIr5Lv3AL17awzxX7IoRpQtSTcbTDxkEWNDbHzooAdo8
l2PMxEXAzF1TD0+gaWS2uyJrEJ4OhZ8Jgtvfo1qpWyAviZ4OdLRmnRC5/rsQ8Gff
2falaApPdKwHIHNztKm4zdCBvnLR6/zXcsfLhP8yiOF89prLkHmS0uuCx0td8EsE
G/Y6UyfyDZYbQpt9R8h9J8QJz1ABbr6tnNVa+/LeFghdIyiCOPuYGKDXSfwwiZVS
umtqAlRG0xz2xSGl7jMgXnRRZPKDGy7WYuobXs9Ebr/2tCNAPyEmy/zwM4hwbQqT
A368QC6ZLStsfrb/QhU1QigX9FcA7zEGyzXGCaO+GSO6PfxflUUts0q9KQnvSid1
p6CVK9ozmFFr7SXgftbRCpMTr0Zu8DTj08TBCxOF1jAT4cNV1EYywqgBRiQsCZjn
VlxqRKr4IWD0tE0DUEgM3PsIkuvuJvvvEmb5rQ7fnanxJe/sHBGu4I8W/vt0ku/X
oIh5Ih5g7p4896DIUzZLtQIWSyKPaKf1tFc4tGtk/xG+JKf0GqIefbJyVJj6Jp3Z
/PzANfaRAEe7I7l3YJMBlppp3+LCZr0YuCd8EG3UhWd+za7O6YsiRpG7p7Fwt7Ut
DoqrfOuxIM9ccqnGHAUlq/CiNw95ufmn1TrsH4CSXGV6qv+mlx9ui3tC1oU2AECk
ig8EW/Sk43Vt81e3P5w0tppeS/K0LyEcQ5AdT9o3YnTHwylYSMBHm5YSKZIksbIe
opkWJwSVzUzZcviKqzPs+YVMf8nzxKFYH0MmUrJVAMJ0Q8cEh4N/yUeQ/qcjSBTG
SxcYitfTvQUHeU2cZ8+nS/WgCEc05yzQkCDL/nBazpO/zNIPgREmDcXStSdPK+s2
vJUTeuNn2RN4x8cnjT8MDy+ecb/OWTYVNCySb0JaY+OKDw9/eWpR3FHRt/UesLe/
nzp8zMtf6QiBa/rjdZAHbiGqnor+ErPCc0bVHMqC6UJZiNHEZV1/ZOh8WnQSstNL
QWC/6vPWXY19axJXqcLpQ+lW85gpvGjXt6aMyYFjav52TbM5mOLhR82SmI0eoVo8
cweykwdjzpP1vNn90SDZB7dstCYpZhLlwB0eWilmYQrXwvOoKxFmTePBF3E03L1Y
Bs+Ce3Gx7bzerwYf/0X4z5Wd39gpH4J0wWW73ystalcao5oBFpkBJy1JWMkXA8AM
rW2GK/AaFiFOfpUgWbsuCyGrQIotQsEcZI1G+3i+Wm0ryFXibeaoUI8HUEIlWDEc
XxcKQOzmiWEQX5dOTkMRPsXlMfAWKQ0LMITFf9iJpUzzeu61WsVJtehE5nq7m/mS
VGJFM1BdlYgr+RfC68/JJOBNRgOimZaUSfWFjXr9ur+RK32//XWbMz4X4dveIafY
w1z6IpXceqw7SWC5J5/D6GaJ5PM6qjLHIarGW+rTH04SHKfBQmjo68tSuviH62x3
UZ+f5iO57Z0ZCjOWyI9k+QEjYHXRXj4+mrtGYmiOqE4/R/FdsNFQiw0B3zY80nW9
iGkdqAeAYS2wsUOJ0v0v0g77clloczC9ovenWs3P2zK5FVjwRkZpIecyobdwQ8S6
LUR1TtjqmkCFy0BPri8ycu9WRdP86zAI6qK/I1mHdcsLp4An7NivLlj/BeK1Ljlv
fBH1vpLXeg3hWTsLTLbiA5mS5G7ig/niGB/+01HevxsEagAVmx6kL9LujdrMYS2Y
LjtqxiMPlkK0NhhNsBZTx4RY27R3Chm/+1Rju37gykV8qyNKoiznbC+y7Cr73nTK
j4ca+fjWPRSgCeq8EZ9LpDVLC6eBJwFhXTG40OTulLhkTyUhB6687yCZd+tsn5Ay
tY4NESS2gf/nO7N1/eDqSYZ3BniQV9Qdp+O6ZCVi6miWWTntGQT5k7tOgDL0rUlq
AHdZXnGXUSDehYV5k9A/b4ApfvaDhWj8tOWhfIcmr1GTdB4QtTwbEr/t6ckrN9YU
nWy7XozUQG7oOqdOWH/lIcHIFAsS2OzOWBVa9SZxDu/RwqSSw7rMQf4O9SKVi73B
jed9iiIqEji+attHpOUA3dg8G4a7IERHFuRlRYOryk/uPWKryrlR1ZBP1vvEegRN
Dc6CHJ/G1hW3v4QjVM1d+/SNN6x+tlNHyM6CJeaBc+Y+0VrCxqvDQNv4A1afKA45
oJZNKlpxAPBqAqLwoomNcvAt24zK5InHEBgGCL+tSLdnsn4O8KeAMyiI2SksonAs
3UhAL9JcG0NsnDQDoDDXp0n1ioIBJgs5jK3c4QmuCAEoI6yZNMnI64oCVV5ILYdA
Eg6qJJtIaRTF1+VZga9Z8jNEvfFgHa6XLZxZY/pehuxMjYlbEzbVKqbDYum7NwIb
LdSdDlrdDOQ9n/AOTnwQ3CjfCDuqaLXqTuXPypYXzGrs6jxa9UO7JV5O+L5qKR3j
42D78YU5RMt5RoxI28IdowvXaBVSib5It5Mve0zIRwa9g/zNaTvy6kLcobHst6Ka
6OwzhUv8wDx2/WHzc6zZB3bs8S2kHwDTAF3fIJ5vdWSBxRb4EcznCkDzvNiV6Iej
LawvfOMgfJtsHzO5x+94LTQwIQ4exKWx+zQfJ3yeH/ddeOI3l5YF3wYWjA/vgrKV
Uov5Hn6VttpvxR7M8K0MCKbr5pD8/GiCP99v9rx7qt4P+U0A411o/+WgIDFgxLfs
xf/qIsIpx0KEqxjBcuyTslzkYH5NhgDY7IMP2w0Z3k8smVkDLYkdfmuhETq9gSlc
QHnAzcSTCTwCzRJug6ujsbbpVJk6Cr/D7C7UzDqw2uehlfG1ILaCAbRHuJHKud65
Y8qpicOEsXQLlWgbBpHnNq8oXOz03IrDlOS61H/kT/oTReuXf7HK46Fp29OP5Ukf
2zBilnM9IKrJt6Q6NLaHUhFoDXeds05qwXdw03hoF+S/IHaeyMNqXGDOvGx5qHTr
NzVz+XYDOu2qoyyjXFJdyYOGDSbfRzN4nR0Iijs6uaB4XY5XRt1oNbS7Y0zBKqnG
04uGI67LuvMA9R50iGelbAGWhzytR2GcORvggZZLc2yi3/0PqKDU7KjrrXqYJ0SD
YIHW8xWSpu19HpYHjq6dw0PCTx8P1usFIot85UCE3gk+NykPnV33Sj2gk6zFsTNJ
1Lxio0c68kK3uyLPqfdnzjs3++XBHoT9y2F3KI7HS4q9tZsxnfQ2hSZXiTYo6Qed
W+5FsVLrmyssUFjc/esZvD9R53oCJ4lPA19ZkKOlWPjpXn7meKryam+JE/VejKSC
jdqcusvf+ojJFk1GPZ92/Xf7BhalbYeeId1SZUDUE8LhxSkJRNh9TR6EhHxaXdci
kSeshA+sWGb9EadM+Z/rgkQyK2F6CHH1AXxbxdBK115tbFgx3wuDOLO39EAaJI5f
Wp40zYRYflnpPbknEVX0xttFQKJ1O5/KsxVsy2eP8vE9k6eMe973ZvEW8ZdhSr+p
Uw98jjZJVRLr9xFkZsiLBkajFK3ZQpGFcND2dm1dYItOG4iaYCytuTSvfqDem66A
vDp9t96tQYZZi2m0IFEdqb57gbRplxf9zAnW2QoLLJMI28/ONFiLwsTMt5jrvRJN
7TYbMZLYDMJZsjZL+uVF25DEoXL2In3uIK9Ew5HdCsrSaORso8PUb3e4dqKZnXcs
v35+2f7s4ITWeNFuB156/GN1i610MTHsSMq83fTP8ef2JEUbKZRLOBcfUPQZSbSa
9VgbsR+RZwpWP7Gp7ljk7jIfdBJFHOUjTk9YeiL1Bl12XpeGD6ugKlDwUBbmrMg7
rmaaNaP9GGbmYUkY/XLfeqdqzZMX9bW+SThAwh2q/MsAxPds3OCDdwqgjt+eC0KR
ZXQYAwURjpdRqGlrms4UYdTiXmqxnPdEW4HMoUEutgJ8/zvAshn1I5uykjaWMnDU
sgdvY+ohIrii3yZHS9qJvC0IMdu78QyF3pXx3pIJMYav6gDXols1l7HO0rGJyJDo
cnvUIzqeaT5VfvqCd+f1WSiNF5udEpQqAIErFH3Ip39b4eQXxjzXOMqR/9IpssZK
Rqdg0pCFeIQNgLNBFrIrtcprBYAU5idLNEF0y3/RIpDg66PEF3BpVd7oKXTaxeus
zkkaDJny9uYXujg1LW3ebep+/B+X6q6UFyPZjoXGI/8qNWYfF4IDBeIXh+odZmoE
Ty2Dbr+lG1DAdtYSXHRD7xXJOASzcMy/Yab49hUsqtwt1Wrwv8a5nY+wzIjcUnbu
lc9mrepOUFlWsweG9zP7SuA6Yf/LUQ67WBX2xc11YTfkK6z6d9HNWct2ND7P3G8/
tpprL3JDhUSc7jK/ztvkFQxRB6pOyLLv0Y9ZFUkf7JEtk+BttGbdKIfI3wlcMsmF
cKCQmzWfaZ0mpHvij7u4MOcce4RkXoA8t6V3H+4HGGBnUtPETH38U8U/uyU2QZhc
E7MGl5BvmReVoRSos7jqVtx3u3n63IXHBKe8/+NiOXGgts2aP0Kr6W8zRYU7xHiE
IWLvCijmXhLDK0HIocZbOZVxKL7wmp1UIRAGKMPDNIz4EhY1KivQdQG/jsz1r/AL
0Vq1vcNcrmQhJLCe56LEug8B71RXGuFDIPpc7o7ok82t5JUfTz7cUtx6DBcSHLQi
1jOxfGkXQ8BDoOipC/i29oTQDQsZMF/d7mktPDE3/bA0IBM5h5uIXcjiNAFxTCmc
qDqlzIY06Yt+MrPVL8yXrHgGRm745XMOlDKkQsgJHg775zIk4sCLW3BSfh+t2P+s
x6ocFsQv+XVFZ1FEbKL8rHig5YYPt6vwMKL4zwFuJzCHSoeeoBI8u+mcyiVs9Mx8
nUerbzCLFFQOabovhnB1I4coOrgEJAfy4f/nubSNGQ/feVrDyijN4C25wgS6YnJC
p7mjPUc1e7aXGIpDMEpbgaDx6PEYz+n99KGR79V1awLObrl9KXqdjqQjHJRhB76D
l3LGUzZLSkpxnXKo9eAuOChtCNtBof/3vBi5oVFx5QpMFE4rci8q0swKewVv0DkX
h/Ltt8+aA5JZ0slTrntjCz9uDYfShWnL9qfQQbasNNZ+TQmo4ni/EufjAWUQjZGU
CduvcpzHj+TVutn5FFida7kfDbKg/8nwOOz8SXHYl7QllmdfrtMTK6j9XbeWt3z7
bMIkZkmS1HWvo6Lg7KcFcm4DhT483byzkX9nSO1IOXcL/lE10l5RjaQuZPz2oPUR
ZpJMsc8UBxBYqXoMbte+ihYoUIgrV3eZTJS95tn49uig/r1aDf/4ObqJJEOdV27V
Xczl1tWPu9Yt6Y13NAso/ERSGUhew1H0G/YRqXmlTmPGLZacqALJK2oixtWywhzi
QxxvMz2PSrNAp1r3PmrwqBOtYYVaI6NUpGsHwhxz1vOXSFFpbqXBJLFhoyo+EKad
GtNiqdiD5FLZOalAhlSosc04gUv4uhqsEtvff5FJ7dFZH/ET+UVcLTiPNmpfo4aE
yWvscVhbt8q5riDwQR11xhqo5RQvfTmtjUy0+uF9hy5zS0fXbzU37XBMj/t3cuhD
EyLUvPRpJnBtRT3hnd/7JWmGRBOWaciOxBmL8RYNF245LaByTr3bqmJ/DNzgiY/8
GeQB+OskviWoP9dNrUpEmrSgXCk6rQeah6dgt3641UqIfUNsZogkyXzwhIyQSZMP
45PkLhEe6pgM37qZagZIwPg9CLCJKvcoKEL10NilbU7ZLugoVKX+hBvW7okOkBg1
FTCAI/iQK3W+gUORJq9nWuoMyzGZQsNduYrvtVn+kXLcgAt857mLeZYE6tZa64LE
yljNt1TjnWda3F1VxUjoo4FVq+RR/juGro32Hx8scUONFWE1FR69ue+74ynHvoyA
/koZRUG2Hb3Qy7ZVJFZdtzyaKRKX0nWizQM9UYtDlv/g3e7jcR8WL9zlUaA1u80D
lyCIujJBlLRo3SwXPA9LQ5EZ4LWmYp+Lwz4RkyBcjTZ2Cpo7It1sVOVzil7gOH84
NDluhVNOqnMHsh+jRIMZ8WqoqorRmQK8EIo1dawshXv0g6SVecP+VsJtdzMZ5KBM
pmNQEH3TcmQR1dGckxMk2Y6z4/xUUKk2khcd65hG6MPsFPf13uZeTODAn/Claa3d
jZpA2J0vuTbtx8Zoz1ueeP9GYFe+OXGDTmzCIdeQKIWuQ5uqKpIOxZXyBLwmtHeR
3GGTbIs3JBaQ4Vzyo1j67koeq+BOQ29q9/M/KVsXSHr9PaLXYRhwMJzJ9yCpAHeT
+ujLHrDD7+1nCWGz1xHv3tLXz6U8P1e/c55i0Ki/VD0KeY8M74hW1P9eKuLCr0se
2zGNKSpOReOf5k5kSeLLAEL0SzvNpJOOuz024wuLGERKAalrwwE25ECnHXyVX8s4
iOxyLpCkARDgPh1pxhw9/l2fVrjUR29gQT7mRfUqYAHjWF/UDMIoLQjlrkFhbh/Q
D8wEq9RozB+s1iqBOPysZwrMTouyquez//5kmyyrdls/k/YL4tZnM8Zf1Y8JYjgp
mpAysL5z7pOP8UgUS+NxJNs0eWboeCKcRoF7U7OptoDG5/UR89G97AY6Chcjfo68
zxXmrNE1U4L/CPW6bNd6GP1ZgySpoCTUoMXSxrLCMwxMZFCvJe0CPe3vOEcou1f5
+NiAF92T2z4CKEc4mHkDYOCtm1wdA8hx2jL+w+sO7TY8gdjwjUwcHzebsIyBhuMo
4BMRSdc0oxh7dJfMZ+UXzqaamacuSYrda1XE9AMk/6yHMCuCEX0s5qlTfIVlTMqs
3jSVMm10lD3LiStysJFn4Av7YsRmItZI6HQRiBO0zXWzp9vFMr+PhGDXMnKwFysR
4HtKHtsfa8nWxYO695lZn/dZkC3oaieQ/3LsYvvegfP4d+GQk9IAq68e864fb7iH
8DWS19kpzgXGcRlEv2wXYCBBeqdjoxmkOLdX1CQilnpogGmC5RT/R8nEvghVOOKY
JwHDnWHsG4DdiaEWRifjO1gh8uLNUeNv3s8Qvq49shudpAgc/39pl0CgMEntnYpp
V87MYJQLlGYj0e55HQZ8GwDss4BNgcLaH/++XrHYsbDJ2UY7YXL1Nx7CQFw8UcKL
924maHEV+KEzfrCzqPCHyfZUTfMdwC6dJdAHDr2q1JJkMlxnaEjeTEcSB64XDFLK
zQtS87P/MPNXMcLJu1gu5ReV0AATBfIzevgI96OVWqbgBUmEjZ5peBJGmukD7yDy
r8V9iDmQKgdAHarsD0FVqbBsZ71DDbEU3hKVdqwdplYtjJ6AL7iH4yG329X5nAvs
Y8ylg7/EH3z+RYJu7NwfjUCQEWuGLLoDKCHuqmYeO77N+RdkGOnEKkYp/3x9/Ymf
n3qXgKUxl3AZchihT5PVhPZ6jj0APRPWND3MTzP8RiBc4x0W5/CtSYz5RP5w07km
sCFcbfk+2I8A3jGiRrDjckZ9dnXHN+wBlQWmzQBOCo2Z5qsMGTXnyEL5WBQ27w5s
Q0Ly1c3CEEKf1VEjus7MvDjR31lfe6JPGyW2NS2pNp4z6QUztmZOBdS/KErxog9R
syleuS+9nKBKpUIpCv7QsPoLbJSv0NXWoC9h7TMqbm3lwgYn8/NXK/C8ZfeT+fRD
yOvtqxY6ah8nSt/hQqMIzVqpEivJFpJZaCxZk/Pi6rcCmrt3cBHhS38KpKHPQ7/K
g4ioyR/p47KOaaIjk/PPOf821DLwX8QJ7rncy3qS03BB/MpukYmv3zqlaXZGlSWM
I9NqSA2aTcHdPe1Iv8Sg+0OOlCd9URUmevaFd5yrOU1avgLE2NXLJso0wYcw1ewp
V1ctZyKC5m48w7l+bubgoze8A36pY4KGuOnD182mLS9Nl7CLGXqpYK+PQV043KDa
9RctCrf59a1mzMU0JPYnhHYeyd267vLxKgI/P/4099QSvTzJvPYCdM3TabRmLZcf
zfX/4R2dciIbNPRKbD5OU7/OtYwVatXhgLxbtStrQ/vKHnU/zsQlrW0fmY3d6+ZZ
hgCwCPyOObdT1o9pClbBZytSIETE3IMmUEvoEPqziZUtYmVk9PqJG+19oIcmUxnq
WHBuQFCTJbWnwpMuHJph9fb5xHijl647aq9HaF7HWOm4b21i8SpkcA745H7LmRY/
0Ya4XpHPcqE1Yt8y3ImPNXL1iu5C7P5OVnYc1a2XwBFDTQQpItalJZIsqtYV3+dA
gmWrPLqPKrDQt11KdaAGVoBbsWvcmbwR3zfhXz9SZCWU8xpgV8g6fflmSjig/isB
F4ivRlso32uLs86E+MhKZkwv+iYFj7wEjmhNfOUsbGDq19xnjSCv11W3WUJbKPWX
PqszRXlSMkP6qF5fAY9rrRz1AwjJJ6zVpy0UdPX2dYp1gSLMadTEMFZL2YD3o72Y
vv884hDC4Ohya0oGWFiTjNY+6EO3rQlfEvSjXw1htoAsX2ouEoSJIu8ntjQ1kv4A
VCTqLPncPXVzYuO5VFJ66uSqiaLI0opM+ieRO9JYC9/gUvEwfFw8gBBDKDsW+b09
XcVZKPqRAsJwU3/g+plHv/iIujIsKDYONDlkUgQ9XLhWQNgdInrs3fLZNUwRJdKl
cBegd5tdcBRyUds9HYrhAc19XMPp756kBFDKQigMOpoAgzwvyoBuYp9oxkV/EHJ4
Moo7Ht6uh1bzhqxVfrPSq05I0nO9wwoCshySlb6CoezIDiNUjNYhGToiZ5zdVoF5
9t9TZEqwBooD0Cimfak9VTC8TLv3s55zf7vhGF2C4gu4oVJtfinVlMPbdNrBY7pj
unl/kycwN7q3jS0J6jkBxxiA7jGsk1d3bmsovhLotFGK5lv5p65smjGX6VZJibqa
SlpeU4/0m0uycysyHpwgG4eqBeP2UytQxD/PwcwDUm2QDB9M92BL5Dd0/JqW4rPL
UO+NCS7lKmx5O7w6McdRtR2m7yr7D6g+WWfTFC+HUqKYbvvglM6u1a5FhK6UH9EW
CS70833uCd2zzdGFmerl1QtW2i4XJuuCheOCJQFhlyhDbF2i77JpnM+7Yv0Bf7PM
ucU9kNSpx5HrHMOWYa97+dbhRq/wsDRmwdD+zFWLhxJnU6nYm8qMNxfXRy5FUzst
63zk1D280Z5L+qlAH/nT5tQpBZgkdZuGiHRt0P8RZGXPfkNEJh5x+IT/LCDLQert
VPyCQ//W5dYRNzy5MlA7kN1eKOXZRUVkfgvH9tWJvKZ39RhZQtOkhRlmTZAAdWnf
hAYQYvEMBP+zqm2T9tLYHKjJ/OQ9aObk1ZgnSRo6DpAIIYS3ii+jw4asqOdUKv4j
QMZaiDXSi2fRAVtCbCZ8hs+O8qsC3MdyO0rs/oF/d8ht4YrkjucnQTqPM0wA3v8y
VhPtJhheOapc7QPwKxQRb4qn5xq6s7Ea/ABJXai0iUGsLktVe04LGOIxbdlNQaGm
8Ca+cIoZSYqgRDkHptfYGh5aYcsgJgEKb4JACI5Mn+o2mamljN1FbDyVJEv08ArF
r/X4Qu5Djp8Ji4AKxbbjnHX6iHRHnanfszfWwjY6mHLtRqF6QYYYAEWFsE3PFSPB
SF3s0yA4ANpKL3eCh0pH4c1uI2Kx8XtiKPd0Ida+DR37AVEpMbT80/IF7ooMx5VV
ligcVjX+cFZOzkkXrtRBlKhmAW+9jJYRF2cmATt0wHUVGU4zmyY8lm6WExOPKr2G
rdifdFvh3mqw0jm1XBsD6fKCcQVfR2i+rbfRCjSWqnmzW91VuaUxmy7hQCy8VWqW
zUGsKyYv8vH7Yl73yZWA5pf/SkT9e2Uelvnbyrn+gXMPeLH0rlSX2t9TVcQbaxpG
9YrULA8PvHQ3bv2Q+e0Fj3GrnsDQXt6cC0qUMM/whB1mW+vkJUYxpL+14Sg9G+dR
CWocA/3YSpz7MY4uErXMp9zRM6C3ZpEMBRj8jpIyJi38oKNx/u/gCwboE92HT0Al
iz7SkSwZx4nXifXck3d5S19YC3fbnReiVpqlsL0xFQD8MA+T0ejySvgUvxZGoTRq
sTZNPqHHKYmiCTSxdgmksaMoVqwV3zBvH6GKP6j0t9yOMKMB7vJrZww4bXQ/Tn6F
qzwt+j4BYj97A6TSSOAjcmPM25FHGuUBRljlwF2jaBgYu33OrTfWoL3NjrNcFPKa
fQjczChF/EfTJ5f9x4daJBctFkr4/rCi/SLeF7R7ji2LM8zE3A1i5LkXFZWMHXEB
UqShPxA5xk3xDXlrpJCHiRWZ31mdf+OdG/I/7jSz6qVNzONUnKZiPTGLfvkuZ98U
JBx4wv2kUrmoghcLu65RsIg6fpw0EzXnZjMo87Lwwrp/73CDAwCRnaf5FcxAtBf0
kqB6wySb3ySyIYfElzplph2Yjz1GsoLxpRqK3VzW1KWSLE24foQMw9Kr0DkXV0Mp
6ZsAHPd8wlCz3gpyB5JSFhy6ZSPjI2NFXyjIW7BegOTtJmLwtE29JAwwborBe4nn
24EWyX41K8cX37b3qESe3GvH6WRhrJqghhSxQY6N7DQqpo8nFP0sFtZ3RBG2G8AJ
PYKtVCkLS5CLbZS7VPMqteMQOChPoqZX0R5S0UeVZEoQ4VPX7kSq8q4hHx9Z1sxX
p28SbAyN7pHm5rOkRIoFQsYcu8s94VIw873ESXOqaCv1WJ7BBDwSuPOqCs5XLsil
m8CpO0mFDVk81wxwVvVk2pp8LkriuK77qoJQmuwPtlhmW9J9gVHJPfmPkUARl+ur
c/uuyubqyQa6vDlhBIYaorlnsDRKujlir8QSz6Wtmd7gWSb7PF5SV13R3uPs/MU6
buEMfH9monwzMTgZWPGM85KfmnVu4Gljd/vncBCoKeO+oYP18bPf7KZXp9/IPtb2
xeQjRez9GsJ5Lp3UzzGF6j6MKS3Qac2OtmmeQ38lBNOA6I24yv1YBZtq/hRvTmAu
d9TpQahs/LC93FlFTaOXs55Rru6iuQ/WtDC1pdxM7DslO70pVKcXr+rElP89MTXi
pMykTOczzrRFQd1uDe37ix11k9NppTLfKY+4CP/dHdLPNFxiYhqVxGYhr7S82MSi
41JS1tHSUZ3b52Dtri9EnVxkJHPheEn5KZg20Tt7HQLzxNIjFffk3IkbtjnVnmFO
TU8DZxcjOnHg9o4SFVNrnd8lzubiZN1yVdvkerEVC2Rq6wZ+z2HQM/rYSMzi5YEY
xL4hLzsMGtfxIcuT6aIYNMlfia0MkLbwO9tuogX7loXddYnZ+gd6FremJczqvMTg
GASwJciMxs30MoND6Ykdp09gBPMm0MHI9BmwSIJeH+yv1EpUvOWAASBkUX/76iyh
POM/kTGyuEghHZLQq3BsYAViiDrsqQXboINnupaPTjxx9BL0GdE4jnErpFc623ZG
fik25g0dSGnJJWPFMTSFfixI6w/+tf96c7H8eXQeVO56OR1aoTpvheUFB/EqeKTO
Ib6JZJWgjhXKPwGuYrbD3lgEF4AObYWQbBr5IuwFEwOOJfpXFS65224vBFuOVTn6
FvyVSe+nPb5KkhASula/QPbPcMNuyDj67x1w85eNbEh5IuhmFgXKZnRYraV4I8su
BIayr8NF0Zr8kEutsTsrdZd7Pisid2XnAtYW22FulZ7PvcK7qwgC2VuroiASqPdx
EUtDtJgdjGCrt0Z5xHqvFKUl/cPNqijjHHSSLi9QmwgDm86OuHTBtHTa/kfsWTbv
n7NYs83GgnqhsKwqREt86VNq5mljkVByDhBnemC1fiUncuDxq+HhGh67B8MIQe+e
dHQLDn+sf0gADf0Jxn8KQ1LAx6RiRHsaveL9ayvv7YywcEcR4u+Um1orM0v2r87X
AQVJt4/m9e76+NJPBmBJruRxcAugRnpaJD3fmSB9c4SlZQ2SBd1+2d/ldl1t1GsQ
1Ed8pEOB/Av+ZnVuidUpRCMts7jQyDI8VetdCFvSEjhukHE19Z2DF6tS9VXA9JfV
DA6snTfCHB2bZEvjolgaj4koRkdBf5BuH4S8dXovYvLf3w5CbF03npFwrfyFlRHx
ngcklJXCkJszqrFlmEZp8/peCQFf9c6oIHp3zRPv2H30fTem4hlhO8eSy6ULG4MU
OKfLF1zK1di2pXB8jMz1zQ+0BczYGROXATrdhtWp1SmY3U1ez/t+EeFZW8KrIQHG
Po0LhFHXIGmkl9a/Tcn63/LpffnIb5hzZ+ELYl4kXnOMArf7hfVoEEztS0cUFKX6
V5Vt1PJQle+TtOD2+aFjlDSOaUVDIefbIm8nLmPym4kDw/utzy88vbhqlx08cdJX
SulQjAdHAsUDpF4tkMGQEZ9425qMEuRJuWU719FaITfeD4cIz7gDnhHjrsR/9Qni
EteOfVBFwFnFzUu5yXANvN28znDY9OrsVHy69SjcG8KCc/GpAG9Vq2P1fzooH7KT
bUh28TYjk1GXOXGKIlpQpuIibdGXJ/Vj279HLBypuIoV+OUShHsYuG/ltCib+qLn
OqOTPeAYAIaGk1d4aygEdpcpLT7k9HwsRrzGMD9xbWjUx0BwdJ0Q+AJxu/CrCjYo
V2+OCpL9mMWBmQfCKGD6CZn9/nlX8lNdF0h6Tb7DcGToZJpMiSZGECQEoXtjF8QC
250J5TtZPW2zXSWXicdPNH0GnXG4pyiadLV7ViKSJaccWeO0fMPEkOMlerKwPKjv
sL9XlfSqp0j3jCFIrzrSMVh5bWhUYJTCoosK+Gu/1+4iBExY7IAyKJLBCNkXvyhk
KXA7fnK907cXjeNDKPQQjgAUoRe6dhGi74benChdBWFlZbypoEPljz6U/0CDy/k+
4CgZwbczr49QvOO1KanGyyujp0YirSH/9FglzRKvoZa0M7RCBc49Ad25HAolYJHj
fbjAOoYX2shX7JffZUklB3lmpnq45RbWfB3Oy6up6Lp29zWkrnt/hHk0MmxCTY7U
3rlIzE4JhzXTnCg9109iJNpCweSpax73BQxr5Uk023uSarK4Rx6bOni/6FcW/Xgr
o+CNKyJ4DMij5Pmg1wfYz2GGHwY9bJF92JOD8dAaOyJXUrbqG8Fe1PJppIqDFWgb
klgndT7qFWDfnnY4LNSzK/HvmrN2SLN1NU4qrOhIzyKqPivpBIeWLuoQ0eH+Vk3j
J0rJ4Vt7xO4SvpebEWxgnSKejzUELMqf5PqDEfTbKcEOfZojc778HY65MCyHdccv
tHCGzTB4yTA2QogTgaMpiAs0kaMNKCXIWLq8HMdrb51tuSeU08q9G++XhNyYKQbN
vxswMr27Fz2scDv8OTCIc+2M+IczEGyVxf+o5w3EG5ROWM3eRmkWcfoyKGE+lvr7
arcqV8k2eCQqlc8wNGulmdrN4gxgU1AN100M9dFPgZb0mGYcKZZJAZ7ILjB6xRYF
76u/1XgVW+Q4Eyw5wq78FrR9UUqG2F2dy6x7TBhunPqqZade8OleFz3MeqZXt0Zn
l77kbAFrryGkiPBEDKmbQUwcPbC9MP7ux3XNw4Y0z+INOZ1euJ/5fibMFVr+nRnJ
z96f73XRY2HAsrEy/eC+0ty2mdTtDMcQQh96q/7NezmUQzTfYQDxmRTwWitHrNwA
KI6t6NYkn8uIr5k6kwGgfbl1AHl8lqzxeiH6pe8ZXTTMriMO5A27DAVxcYd6md2b
evRiwY+BN7eXo2CFbsi/gnSygtzyB1rGvAvEx/aeBTmNKuPh87ir4qSjHHxgKpp6
t/B8iXMzzaNhDUmWQBvpu8TI5J8BcEpiOjpFWnD/8sHGM+RNGvhTLxP4bVvaftWl
soBn2nYeNhLXBV1Dsl1D8WGR5d8UBnOdGu+P5KBBTiWUvX7zTZ5DrHTKUFGNS9hu
JTo5yNjRaXOD9aL1sK13Mjx9HhhclrDNtspE2YXfBY3CKOciiakw4FMbwaY3TfGH
zeh5Ml3o+vVmegOT9LXUizqeKWrj9MjeRViRCku2Zm7z7FONFvnzdS+pwSMDZQ4D
wib3S5I/khEIBMjFbZIWSfTa0U20SLl9WZjY9E11meRCpHcK9cqPkzTdxEPQ8H8P
O2cHmeKF8YEj1qa2Xe8zXUWD5j+29d/9sxiHLXXrV6U0W01JhDYbfjcEQJzGOqGF
wUVeMb3yaisX0zwpoRzcvms0hjJM+bAYJHyeadwc/v3w7x775uR+/uXO9ADoj9oi
lBQq4AntyR/TTJn8wWsfv2/JrAisHq0FU3eMijKgHw46EWFiLyDMc2C5pwskWumq
r4ZUQaGisHFgwWYxzHArWC9+EdAi9Iuu+stX1jcc9CFyPjMVfZO+Z3IKrB0ipmTS
Pm4q8+p1+At592QncwZmyoXhs99Ja7rPUNotgtZdA4N3Ew1RBqSyKWKE2MFZFPJ3
DEesxB/oEW3YTvnugX4NwU8fc7U/R/WcuuhTl3M4mFcO/5j0eVaVvDeWbEiIwiXt
SgmgM+4ZGgdaG7d/uIpH1ruC498DN4p2epJqKuk5ofnJTPsCywi6ViY79te7P5Wz
zDGOGGmhRsZHKK2je5eNjXnRS+S5l5fdKHrCo8tukwlgWEsCTDx0/8r++j3c2nQv
WND9Emg6Uz3YpP7nbruHPT/iiJRuiE1Hy1v+GcX1mXnZi81ajRfCvB7D4vTxVUVq
X019RyZXbIns1sdW0h7vcqE3EANmHTtoOBUQ+JeventuPqy5ytE1H1qGBqJyKyqP
3flLy7Soli3EG+eWWEYTa6hEflm4y3Q5PTCK75p9R0PQ7OK3zToIXEG+eAzGN2Ub
9vq0Q5nGd3Ps67rh+x7RBXyFxiTPWn/BXVj/Toy3Qes8eKnIdIelJQj7egkaRTnm
TeT2tQm6sFzKnaXfYSVImjr4MfLb3pm/MFKGNLjGh+4dBG2Ablc5U5G55n3u3y2Y
G84cc1GL6nu5OpssiY1DcDyT03ZDEV7R/5ygVXMYcDKR6FrEWtNdpAszz1+ZtWic
e4bXhxhkljtBsHEXmwK6cbObetXQsob3OWmDA/V29yd7sXA663OhDxizuhnJmYcF
mfT+HFUbmyNoY3pYslQDVTpTu/Yaywcp2Qz4D45YK1/Sy3/KQDkDKRMMq33Irz/a
Z58eP1CeXDM6h678UIttcyVbVvnxd9ercVy7ekgudw5cPzg4j96OQvVs3ArnKYC3
w+KqObAAEWWyovnG5fqWzuM7+GNXwRvkbmUC/f9ehe0md0doFW7xY6n13ukdqUlE
m1DSUvLvsv8DB85tXBry+FsNtrofmgV/rcMEd8wheBytMaDPE4amcPaVtmB72GHP
YL86MxA4z8U3Xf+Qc/bkAzugrkmPMjKau9A1nM9ptmWy3ItU9e26lVW5B9GmfPxm
gORT+vHNDlF6D2oufYLOGxO86YDEgk4XIZwOHfjWDCLeYzRxnBXPRf8MlnmXLocK
cpCfSbL6h3/aHPhPsdof7TwPsZ7NYgWGjxmjJKJBgYuwQAlWlYvllf/cpuIvL4jI
DDOHBmB/RFDiKeB9G9tTCKUY2a1frV1dOoGZgPE6LgDz3vtqVbdkUqSrZS+cLUg3
J9Zeq/7hlpo4c+llMozMM64h1kVGPKZ/09it9/yyttJReDgUGAPASHwtMil27Ofl
/vTmXB7ICl0jaWnkv0QhOYY5O2fPmqziSME0mxQ7+xBeLNp+X1fw5U3aSNcyRTqo
uQpKJw7M0kku8QjOuBUUT+39OW74gwEGYZ8k1VgeZiscFRelpxZ6tNV1cM9LdlcZ
gqcZoC8VZ2XnHEDYpqr9aUHrjCZIvggbxQwU3iKHvHWiHSAcTtUo6b0sbY6T4lT7
cqlHDftQELvrWEwr+vs+elomlQCR5vaq223Oh316yaXXI9B4DJo1kC38FzDwL2fM
AzdqzywbtqPdtcXgDimrI6/lqpVlGNoptXfLpbuPWRgBO8g7JpSECyhuQyGEU4Qm
SOwwpRWtCtj0myzdsOH0nFfKYbJpqYqat1R0C9F2BhtY/TSqkI4e6BqYF/JPjZVW
FN4B4Nh6sRWc4maO7r7jBNPRM4lDvxdPHA6oBBFFVJH4JrZyamcSFFLv0ZV/r9Kf
U73q4ymoDKL5qToMS0MXswE62RZ7owgRrSsmg7pRGrGk/EEAxZ9+HNN9KVXDvRbB
L74caRxNNIGhFTzQMCsG689zM+JCrgzeOd6WUrR0PM0LiY9zRn+t60c5nEQUz1Fk
byixurSaZ3V2Agbk3pSA7Dw7e1dHqTVuEN6ueyMWN/vICupe6/KfwcSCBp6mizx2
Tmiufc9806J7fKWuiQItvlgitkdnvpEVAjzFycckGR/dZHtCpJAVRFBER/5OWeb1
TCebnKDbJotzpwTdN2pY3rrYXUW67TKFgMCQJlzcBNndvBdz1OZxP8J2VyLlli37
g5IBWz6+6hJtWjN+ojqEJ5J/XEtLvVpghp0MAvwuTiSmd39VcMe0KBFLUhmXJu6L
4/SQ8Vg2eyiHOkgspwex5QbR+UGTzuWQHc+YCENpQ7EZ1ODIai6sCGTb5WnTaCYj
ahV7XeUOEowIintkLXkx0xrFbOyvbkLwip77suvd6GnKHMvEWonsJpbiDYdXthbv
xhvgX4OLgXPiYOzH8SOFftNcs1Iww6JOUgpNih3shuisqtj/4cpFoCjvbJCG3nNw
jJfy253oNajDSTFxdAXgoYtLNjhbCyZVLOQiieCDVmdx6nNYjHzNzXJZMTsXIJvb
/RqZiHRAvEXbJsp5IW7b8Oi9PthryMS4ONnYZopMShyEV+V9mUYoKp7j3+FI8OMD
XnhDu9xBcihBq9UXTb9e8MCEuBFkfk9BdM2iuL/674qVMcF0UTvkIJT/IxJVipjb
pWFiSNzKDPuzJKbfKU9CGXbFY23K3tq7ESOkrwQ36N+e3GhuAJbLuEPfb9FD05vT
SZyqFk8CTvdCR9jS7BprOm4P/coqt14CMbvY+UWeuXbk9cxf3mtdIersD33LmwWp
sjO8kAzAK5YIZZHjyjRT8kv/N4q8qDZyr4nd7xh/uf4qrefLGHslVhdHC76WMcBg
o5S36AO5/xk32oNb0IRh0XnQzsdajuUuC8hDUTHNxKwA6KCcSq7l9Zp/K8miSKya
QErTRzFlVxNQ/d/7bOjaDxS2L0Ykc7p4Whq8Tg0A9sqGaJ8nk+vRQXUS8/OpdYKh
mtUB47VZEBdYzxdZiD7cm+ViNymoeUsDp4WRxhrVfV0agpOjbRavPO5fp6b83A2G
ul1S8GwmfmKOOUUMvR95DMUQ+asxCeORPTTAKxRsCQbCSTVyF8yuBqnNwrtJBWov
w43jLw0ITOoK5ZKp9WCfmC4G1j/IL8yt9K8xY2S3W6Mypb2lWJM1ipy5GUNeZm26
iLcux9LbOL/0ugbsHZNBGx7pWQx/9ZSetPFv+1JJbRjDFdqEp+wvuUkfHTbeSodq
nXWgBcJLjhnPe5h84VQOa9Y1TnOWlrKEpT8WrRw2hNxztLxvEWo0R0kFxnu91xsK
SNIKEkJULEXuToKtBfLHViyq4r/CNtUubBNXcj8Nrl0A6RzCiqcpsWiEtYmsc9m6
7oPjwF/RyNhZG7ZflBcmOCYraDWoLiq1tvRatQACn6gS2c2EjO/AZE245P4Irt7g
hmURIYmn7LQpoDRjXUgSyPiM1sbkZHtt/Dc0mcM0DzckzMaXnFT2+iSJDx2K6ctk
ODcx8ZwBmd5T8M3I9WJ0G6O/cU/I6oindCx+mR3+/jMGuQIJw2HLuKLjshjEFqHM
3Y839PtETDblGAGHbvZQTDQz3odJNF1R/qq0PDfE9kSfRRn1HkeF0Q24pMdx1KLI
Hx+LX2hO58rO1UlaUMjDwfxlV0avrL7fQKQs53UBS2DL4L+gohPBmogRR1rZ1I2T
eXHDxcumpWnTAAFG0Ms0guOu1aCJme9yBO+fpEtKFcVJW4dJk1EUm+cKEDI7Bacv
Gxz1rZUonrGxHKnmmM5F1DahtOMTIqf9KOhj28xPa09aDtBEoolfunKi6TU/N64O
ioZ6+xkSS1bRPqEBB3XVdBN6jCfCUiWQRvYx515uum9BkYPKdFDJEitVkR2Loll4
PtcLpcg76UZsV8mlcx+yCWF1BEhTlzzdfjmGypDmlqE3oAaMlkE9BDo2Lg6er6Jm
V8q98ippA2UdGsseJYdL/s0Dc93jep732cYlODgLO1yyNxHjPIwnu4WMvZPuHuWo
Cu/Ax1ja8AwmYDFZuxcnA4iKWD7qPjqIFt3qUd0Gb3z22M1c52AYEkD5i94rJfpS
TVQNXQ+TMkiC2CAFNhep+/olvHe0y/pmMC8posbEqY++8S4x4Nm1xXrOis+hqSaD
lfxCOUIEqdtPVo01DNFVx8UZE0LVztQ7aWBKfRaWUMgFH/dah6bofbA0YaVAAjkj
nT3fCIQLOf8dbQjarfqcGEFLNG///zt3orKY0+DvQmCrbaiAfZ172Qnt0rhqXv9K
bhL1L+F+6Dg2iEpYEw9v9rimYKHAKA/vuqQIGRomYIB9xgAxV1MuLnS5m8ZSfYHi
IXBsAkYNMGjjWgMwofX4xvMws4iWCVyWf7OjCl73uRkno0GUmWyfOwtb108bKKoh
nIBJTL4JKyTbpP4jRma1KxYC6qxWpN2ywkQwGa53JdO4e+w9lWZ5+hoCraS/h0yT
h0POiVD6y3/CElflGpsJqjG3P75d/aeynG70mwUBdxti3ludKrbzgUbYpVaTxi1f
GALAV3q0f49IDUr7ujZg4tn9kADmN0re/gArIQCY5rk6k1qBqhYu4Oe3kfbThCE7
NyTe4f+ZtCOVCrUqCPxryjb004KUOcofm+c8YSx1CSf5otr98Jt19g9kETYoO7d8
MDdkI3kwkQ2m/+YGo81NIkpNXt199GRzERU0g8rEeAc4XQDMsSy+dLYBWsqgvsg0
XZAKl2dLPYF/ll+y/Vupb20DAkzXp9a1K8QEVKORWWEuoVD8uGbgNK3XVLvmP9gL
wMtDmGOWHuB9x7/BTvourNaO3DZm3wAuanIqAKMw/p69ZroTbki5fAugRTWHUI6+
BqBpkyX4aT0vwsJ2vUkxzsEBqGF1CZm1jbK27v+sK+phsDfW5DW5G5Rlm3YIFrnQ
+hFrQDo9+eYkmN8u20vQl2UlgGWnHX4wNvtLw7nxL+uUw5dtistBtnJ2qW6UHdlB
vbFiZsa1W5gxdG7eNniuF88Uy+5MZ7wveFDBpXVAsgNSGYdd2ddOv9ID6yT/CrDS
jFfO4sNJuO9fZyxAUu8C5yl6g4qzt7YhDgB8dpeqKq5vDZcSwViCBAGSg+chMi3D
MrbAZouKcIE3YXdsxJu4xqMqryx5heDF/nXgPJj6b2nMGoL75/7EJ9jFSoKvpeFs
8wBV1KWl3hOkS1RsbSgjxB8v2gOLLeXI7S2OL3E5s7GWYITmq2QXGair23fBK1oa
SEKEm+mfcc3sU53fZXdfLPa6eIkWfArAOLE+dNcwWEIyU687mQERElXbu5H1Ofy1
rtmKKG2TaC4xbRzzzJMX3UiOfWhu7PFxp1qvPJhfJHAFfE0yVX8h17s4xNCbhfVu
DL7ZQS7oXaXfqHYSrleSKjFDCahEeemF5ZAzTX8fZ3rXLeKIz91h7m0rJatqXMvi
jMAiqZDdEdLXTQYq6ySHRXx9HUG31WnUhuncj8IwRHKQuoqyHjkiAHhkIDms9XmQ
HYokrjuIKGOSSkl8MiHBDFwG2G+zHEbMnwfLmTQxFFaMAc0o7eAbf0hpJSwBq+kY
iiocKO67cXysp9OU8LEmi1VGpYRUEj65Fm2uxg5FFoP4e0sUEjnx0DagvhndB1Y+
Exn6YZraF/H7HonAP0Vjv5hY+9uOtJnptOPtRpS9Pz9wtsf4S664zwCVnexvxGpJ
AXQQP8HcXn2SULEkKejd4X6MwvRoozqvxReWDMTocNziGAV6sJWKXrpce9A8D7sw
nZwgFkBk/t0iqxEs2nfZQ3we21v/P0sWrxirbt/yN/mm0xOXZZJHx4sJX6hV+Gik
O7vy6ZIVS2hSLn8/M4O+9hdriyd3lfBNGoS81USGoz6Q5sgxRw3fz3MdV34lqGCw
4oIPDxRgLzzqeFYExYEcsCFj0sUlN+9ZPqwkXCr7Kn5bGUUYIhoPpx/i9ByJzWjm
53CBkVUSySKW1LgGh7rMlh+rdtzVvMDTV6xLlm+0Sjl1taScIuBNGxynLj8nLNXR
/LfWBxCzH/evbzSQfvI6cm8QoCWHEXWN2kY8fhgCugxFkWiu/wL93Bfaa/r97vPs
53qiqILrVI5obptX5am3I+smwuQEAKfZZ6jzE0IloioN3DY0sQmGfO53V0W7QX0T
je/06dS3O+t0niUe6fX2i9RSO4aiL+PSe+fzcT/xhJgOtk5QZULTZRVeeVAAgY83
9KolfpHk7zSdI1WOf5WcFjHv8yBGkDUTJmR5tTQC7ZAPZEJBAhvu30iZXcVNEbPX
BEcPhU4JpLD4RyWqALLsu9F3w/Rd27n3vLZ1wEDFytfvR4Gl+35uSuCNAZJI81Vz
Qxojm6oJx5KFyhdyU89RJYbjOKfvOEwe8Z/wbKawM8HjNWaXAKacketIvvm8lrWe
OuZzY31P+dNcEJhxITAWc0jAfJOey5d1e0ikLrGewI+3yG027/1drcFnJVTIInXB
ZKpuCkA8Vwqiz6j2N7D0AiPLuMDFr3PqQTITYubngQVBSRijecH+UgkR25LjCF69
G7YsD/lQSRUjPYRxZ9AKPE1UqXI+JubWbB/Zuj8mjIJ41o5Jrs899T8Ozd8xfJVs
LiTDnq7LLKzE6Ly7QFjlJEtzPoeSZorlYBQlMsuVdxIyP/0wsmYIAVfxa3jZmU5M
7xCeQWL2ItEBa3pB0sbY1QXBtpDPU0Ij/meHOuC9rkA3thOi1ob6jeUPi/SanPU6
ti0d96YeBK+AP8IVqBbUhERhs2j13u2f8qVv+yV0xqJ1GRa4lQ+PDvLGWeqnFC2M
3RHo6vBs23/qyd4HaUAosgc+9O9pSfjnL/5cv6c3TSiSQ1n314ed6dSmGnVJErfr
iEQBhWja56ccN6JpB8PnHipoS3ARJKKkkokHdln914LxK0mIVbQpl7LOet846G5S
qHvaIhWzWqNWmsPw+eaFQVg+HiozEUmNBnapihJ/ZeqjohAWCmw7l5P8lMA0nVAW
xHSQX7K6VFGWHBj4kg7TJND/H9jpN5nxECbkFWONKLtAEv7dtdaKUpPpOE0ZlFhX
PZf51Sx/5eVOlZdrx00XW94w/OFchORnIbhnmtKJhWMc9glCzw9V+pZb4VTCwIDF
xtU+4qgMdXSeLQc9l6Yxb/APnKDbSbBcl7IfWkSFHu6LU7OFbMq7ney+4s21M2dY
eL1A4iFV3NLI0ci31NKcWTF5i4dR1epSmc2MzKMHfBw04zsROfHeDgJAZhNw8vpl
AgCfH/vq+gRwH81iM2treVXJ6aLn3x4XdUWPUhvXZEtZC5y0ckCUTXrGzPLcu5AZ
bTPeyb7ZMM3yB6DVFon4ho/NJiBnDLNZiJO3Ki90buxCWdr1faDrxdVu1nGyIyXI
sPoy7zdUYm5U1NFp7Cv9Nblw1Fe647K/o5suWXi52tXKCi+E4DWplSJwy9I68Ixy
nNv8uR0pfJ1pFG+uRrpztnfZeupWLRO5Sr9GGnfY34UyF60vSKETabl4gu7Wlho2
Mk1eb0AAThE3v1+DFOddkZ4ovBMglYGoIpexjjrMTN+iz4zQG1qX7a7RvE2/d+82
Imf0RoJmtB6D4ijEYwhyveodX4k//9FL04sdQuAAuJF5PP81dcLz4WbrS5gZ8WM/
e8Nf4RqQ4Ht/LZvHcrpOGs5Pbgb1kcZH7EDcitHjX7S3pvAu739KaBjaqOP694/8
NWctCh3uTtT+ugKLBBMN4kw/fOhyYIjWRkKTITKvt5uONtTrT7jivw1zixJzwq29
fYqSqC8dHHGuTNWwtE0fm9GjIWR3WsUk5P765HacYqedB7Ea6bdMspMH0Lz8SPO8
hTrsCoMfL2IgPKMRGjlw/qjSJDTdBI+1o47A5lxwuD68AQJhrHq+1JX2OI5okHmt
1DjFA7uCxpRmpgKGwL2PHFY6qQUwhv5XMUZAy2XhxWToPrfGx5AZqwTlW7yVUC1w
hOyNJ9M93Oim9oxBE1bAzT0ix8yisU+IYNBNecQuf3eLVThwXnP/g8vugUfZ83xU
Uh2jFK1cVRj7vuVVtDCe9k/ciyOGgPRgAilEqsi2DLtRoimTq8i4NbP5FAm0Vf0O
30iC5D2wXtoVTnZtHhdPzNoyWBmaK8BLk+x0I+VbITUeSwJLkv02HaMUuUTq8ZYD
wBaBv7FqGHMa9SHtdHomtRtAJyBQqIaVDKvAPhfld7iH16bD9VTZhNToekfMO4sf
2zQCZ1qbm1GiNkeqMihwq92Ds90c279Leq/bOeYCptwCrOyuIFqdILo5BxuZvpcO
5QK4zgll54Slqoa9Prwgo0sp2DpSYOXs+bNuOw4ekBXGQ/kNOGnMCPDmX1asqrKk
9xrzODVr0qp3dLy4K6Ev6WDNQxLRN4BgYPjnn6/RUMKla9PIvYSQCbKcgKu3VQMm
MRl0b+5GohhjigpdsMeKNOBijsFCX/TjrBYZGUsdH7bTinwwM3X+l40B4zAbEbzR
nHOGYlo/AVE1gY9Oo4tDwN2tKCnpIZgDkOysdkTn42c0Gkoqt13Z5XMJk6+qVXop
mfYHVeqMvVcE/VwQXhTL8FDEOIiKmV5s15qytfilNwZfcaTKaXZzrLaYwaWsHdpW
XF8pP0qd4T2XBqFatpDfQaLgO2n+8L5Apu3GszSLeT5SBn9XwbpHJGSW4+NYBaCS
DzhYRrsoTzBhggabt3uht88juAQsHDVlTcHE/GHt62qruRldkZ6NydP2Lc3Blp7z
bp/J0cP+JZF6LQ1ZZB3uG8PZFBz9bOABUlFrpI3sX8gmAdbdFlkQ6bSv+11VkSPu
uSsLktsOd1h9/Zv4FOFfkMshAItdzcjowM8MktYQfRnKVpcShZpEp/N1D1R8w4jw
Cbiigcn2j6jYCx6TVqd41BcNWo3IRJRvvcAzXC1ULLRArmejLlqxsuLBuuNLA4IY
+2LjbH9s3LzvChz3GU8bsE+7L27D8NkAQtlp+S8PbQ/UoJb5k9H9enjdFTj1sd/K
hCogT+kLD2qblbbnyrioWui6b8noYxOhuT8OxKFWFip+iQeDG7D5K5PdwfflVZoM
RMdKzh5XmzoPc0NMkHITeV1zOC15OWKYTIiN8dVkciODthuP/+3YgDePuImDk/37
6kuwz09sT6xKVSMOwHOmlgXjMRAKuhMAiEd4GWiy7gM5+A4cQEABebF+FSkCnAJK
Xt5k7VpiA3TK7obd+QDfbAzhaXj50C1U0bdti49amNQIf/PZx0pMDiqO5VfLcb/Y
vcxBQxuXnRDb8dC6o+yGZt7HfrM7eeSj54YykZKPuJJfqq5qmzAgQ3+Yi5KCNpNZ
FB1ZITPVR/cQXo0jMSFtO2S9Q9EgnYZWtUUkA9NfBzb6DsMurYmxKLQ6X/wukwOp
T/wpHCrg+HaR0O28xopy8dol75InYocAbE56w6hXKqLDrBTrkRzwoEkyNPvIaj6a
134mUwQVCSgZ085J5phoju8tIUV1VslL46pn/G4V4hRH1+RRVMOeUxZvuX/bMSlI
fzxr8eUCP0VG+6e1x4moKBWMKISzL4HK0ED8ks7YU9tsA0dhUTC3u8I9x+oTcYib
+leEgzy7p0kPQFjOeDbbUSNVWYWcebmj1agffG7Kr2ByewuXXflbsBTuWzg5bGzr
NAzNSb2uyZCPSozDtl3PmStZdCDpT7Cgoay08dOaexdboqBjbN7PBfbLJDGZFeXw
0ESzUfXM1utfsEHF6bpX7tRG1C82dBdRiVh0fzD6zrh/ociw0CS9m3YQs1Zs2uom
ktV4hOSHB0n7LxSp5H5tYyzjjWBsQCun0ExGxTjaRGEaWr+hDYctCO2dgcIUyyGh
ipm3v5yxq9hjYO2SblRXyijoa9O4e5k89luVGJaw3O/RmlC0baUVHZhXt3CmkERD
1VaRDoOxp5QENWnWhHFG+FYq4Mm1cYrMAeDYoDaztY1hs0LWaMIEZzA/ljZHhk+Y
sU3wDJCzl1zTcqpeV0OqSggR6AM7muHnztoypBs+v/X9P7IDnBTAWRB/992IA367
8quAy6QgpNOOrntOzXsTalK1HS/7AGjisSWEnB7GyrR/49XIVr7exZJlwO3XaEMp
NjKHIgMv0zr+U3LwLUfzo4hJJJWffvy4icLdAvph1Ue29SmDLzcl25Anq2OjLrJt
WwjwXbooAAv264u52UVXh/MDUEqzddbgBvMrJx6kjaGoG9Mp9/OZQt0rztH/E2tS
BcEj3NGJSbRO1mBVUVnQH9wwQ5LoH1Krk3ckGLG09mWbXVcwVM3Rf4gsDCM1j7kl
c2mrQ8D7IOPMUTw5HvpeKPuzrflBLw3t/jj7nrAXG2e2z5XWdTq1uDCUgxf9qal4
GuUH8yZp0ZJZUesnWeoqPsulNHrEcXW/4PdVC3aLfVYFJxvxdZv3ZM66tZ7eRfgA
l26YVgtxZUfXCCw/tXSJfiTzsDW577aq4XAgksxt53hZtFuPm2rhvzTRxAKqVlHv
1UYhBEHxTXsOeGOaW4Jm2yhC8+6EKCYuZLkqrMNxZc9RSvb4dADYH2SM61EA11KD
BZlGXErib9tadqJrcjLxIZWa/dARKm/E77me205MGM5/0ibCQlv3xT3dh/OWowX7
6FfyC5q8s4D0kVQjanAanDos/EmckHkdiuouR1PMfd05KUoidZxASegCgOjlgqQu
wgCR3sgCYQXmb/ApkzGe6csgS/lJ6EAesjDz2IMoAsA6N9ifbAmD9SGzkPVFVFu/
Q53SHGkRpitAl0lU0+vwMFs0pd3jl+EWqVJ/vvUsyg4DWPmu9GqgePqFRXClP/Zp
zjySDt4lcmwyFJmVHz/fcGVnGqnnLnoUvb8Olmeg0gj6W00YOqgrDhvYjmRgHA32
cW59ng0RlbnFcV8iIBMtY/cQVGB0bXS5EaRwE72XB/If0hCutHamqrNV7ETuJg5T
MevLAeTMcwk0ZuRvSTAb8svjPdsDCqBQ1EU2m4MXATUTnptfbMtH/Y8jDwS1Jmt1
UMAzREnemdJyVbfA17qNhDC3Xp1NNyY8wD+KlgNaINpjwMbTFauLZgdeHlQuEwmk
rv0bQ1a2E8ABNUT1KBrP7exXKvFCzi/WmXK3dDdH0/xjCOSvsJVTPX+y2Rbl11r7
HSW7WEmPeSr81aCE6elJ1pHD5hriXgsJOhbZEcBAbScBqEa+OaONFXtKakBCvF9K
iyJGeRF+4ui2O8Ajg4598N2hIMXeB/1EA6eK+OW5gAJ8Hf7U8QE9cr4qG/AADCSc
L3yhyNutcatuTUjjGUuKaU3qnqRoInqhipNrmiG6OQ92HqwM/vMxNIvQrNuEMssK
S4yRi6jTBaUhedBPIZfTIlAokrOp5n2z14Tz5hsb53oe9UjbOi3xP2LjuaZPWoNm
r/O148Wj3m6Ng9qQ4xBdFN/d4R/NBf84Brr/3zanf1X8jETM+LRRBNMt3xqcYbXk
AORm7AfUiNyqfoqTfyJfruOInwv6XGkKjHLxKrXdoNm5zZrwPkdbyYr3K8P7wCZ1
cqbwU0Zgxa0VA8nkqOZZhb91czGga4ddrey/tluQmQcrUFS8cG90ib+4zvoKeenV
LsTuVQsTRWhITAf2Rqh6qh5gjRtGRKCf0Ou1fiSdyosyHnlB9rvlZUarLJdic7Eg
mwNqhz0zKptK5M0GC1S4VbY1jl1owSsX4S74GRrkRt3ubJRU7Eh/ZD3y03r2xzMc
4xy56WW+01WWvq604bTSuntRamwtAb55p/GTeIxoTy+J2A9h45QHmyEPv2xLDayh
saJ3jHcJ3iT05Aztc2VfwcMBuTTcG/kEJ1INXpqMaqLcohcMtJ2Yiglu4dNfaucA
lnqH1eIiiixMPc3mUHkhM44P5OrGXRcWNjF//Xz16s+HTbolQ6Ph45Q3t59aQuWW
2IdrZP/OivVYo0Qwp+GJPJVbnQynZ9CL9lJk7MR9Gb8rUEZAs0Uyz9rEGlvc9Wwl
G3NPHHqPcItkSgo7suSD2HJRvGZRUZKsbjpD0S6UxNbxPdT9TG5eY3o7UShIK/HX
Al7aA5IVb7g4xLWMW6ynFYMoUs0bXR+2hJ2MoK3eVop6bJMoqs+ve/bd2W+0v74s
7zD1W241Yqddjbdh3txkwEX4mKCMXKXg7ufZ7TvTuLPT//UxIzafITSmoz+77kWD
PhdSAt+AcPb/9ymPYdFHsQtfOcQBFW6n9C6xV0+q27Ia8FqJBkTSM76ttKnFC8P3
MoEidVnvJzPFCXgkZjyhuMh58Z3X5UrsZQxzHX9dqIAqglXRIrVYAGlUdaKoCu/y
A8kRbkeHBoCwbG3hxQgKUhev2MglEqr9cweLuitm8nmnScs1Adz3/zm7gDDmfd3Z
0F5FGfXspeJZzFqrwkq+S9SpRAfYMNtuYDjwamMb7Gp+CagS3cS4hAPh7+ujLyPC
mTMnD6ZgY+XAFPB9orRZsby9P1YRXYZnAwMP6d5VZaridqvcRmQNrrAn9GC06Xdi
f4OJ4D0JkMVF0Px9o6wYthN4TS8iG6AxUGXplLKIHKq7AoGUzGxUtr7YhF+j5oMa
xUztZvmEI9Za6LT9VO5wNI2QUfgdm6YnNJtYeOpGt5OYECulEw4o06g7D44QwSdy
j7/ATcB+apoY/hdq4fd+B4wYldXK+wnJ9kW90ePzilgvxX+S6yXRH5JdkCfCcVBK
SdKnl56VqJeAz+5MMnUmodv0nZGUISiGcnH6aCHMe3lKqEottoZVqrdFh3DmHPgp
z82Z0bHPbKnqc3egAEMEyBp7XWU1XbxBIkbi0I2KBk2BBSePasewMNKT+/jeQbqe
FyCFCacs59lQu1hE+4lqaPdgZHlyoWMPdnBzNhr9d/X4ap8uZ+UK72tcVwfOS/C9
dxRIOfzhPWaF/6i51GSz5+NtQleKWzDGBUHM725fCYqXC0DhKS6LMmxtzafYIi4D
TFREwWrrPkWfiP9xOwUADL6D1i/akVqnMgZgTihB+3u2erntcG3CZib53Q5Z7Kj5
FzmwqmiNpxcDGyBtDL80hxelvo0Hlut8vWHwmQTcyTR2XVcMqCtQBRYgKQH5YoaF
sTAKiPPBdzwSYh7Y4xtD5XSneeiczT83PcZofJRErOpvXSkniRLsL+FbXi9u1pRO
I6oIc7inV1+iWDS7bp7BDu8oJDF6WAWQnVF4P4IIuNRL2bBiyb3aijoGu7p7dgny
UTq14pPo77jHnG0pyUI45X5blsuJOBl84ZuHIiIsGAfqYCbjRy2brGFkynXNKcoS
4Gzq07U4sARMtVMPFEQ8wS5oX0nIcoEooAO1G87IV1cfrRlHA6NbGCEYZuweC755
z+iF0IpDDUow0J3eyWubyE+r2fDOMFCJv2hhkRZRx5YsYuYED3MF1f5F6UX2on+J
k/wvotB5WbmYQDjSRGeqOFFpTkspkmuqPW+nsPSdDtMkMD3UNcwrfWDgK/BZpf2k
jkjNaIsmr8UYtdxQLWZKFxUXG3Kb1wL0VjfFnUx+Sx0KUkgIVMvrTE4O7gkv/d+z
xdlHTbsbHDcxNmzvdNAjsJ6F5FpCUjCwu1ioYF4J8xR6maIF136Qs2RW2gWc2MvS
O+9A+qAD6pf10UMPaf3/j/QZg57cif6Bkbzwbw5ItKSjpNbGxwWIkji3WVZLh+Dy
+0m+/xb/M6/FcM39JOS8Y7Z10O3GGibRmtOPeMbqUZuTn9iCtt2aNwBQ3Mez55u6
3Ah0bbPxziuHZER3DScEdLy0znK+/OrIURBV0G3yk25ENpJoq1NkIlC8FJsUdGGp
xBzxcWZ4pl2wUvZMePC5kJDPg3aQy+09VbRaTvKOnXE6TGhzg7DL8jEvBx6UuhzF
AevFhjThYQuPP1MZXL76bRYp/3Bh0bbSUCWHMW2YZPPI1siIzGy+jjsjpaRhSnF8
+PHKiEpSl0LRScCCs15IiKjCV5uP1V+8xS3ItNfgjvW7i/4V8noyIACMXt7dPmm0
EC3ksBHcTPxDYYAeIXM4nMyL1vf1UZ1l0v0fnOP1SQR+1VbQuYUrGDMzm0oTgAJg
VCnSkU0fi9r24sWbJo8JEmPydHKRYp/wxfWCC4TfgLaxmG3ISpR2QU0+dw83fhFT
joN81ZUVGqDVjWVWmiLo+upRD45FMYHd3hCN5ZTy7lW+mpwrgRKiWt4WlvCKHjLH
uvkd+86UnG0k45Zuldb94/sfC3Gfxu63nZUoln/H+waY0gL6nJpJG2h5cDvpgvn9
KZZllaRKo4muQy4x7QO7miB9unRTkoWyjHPFkx+9P4p9BfHnFQAYC1iG7hljxQFD
GwAHqBPDpxPUs28m/ZFCO9KbsngEc3b1onZuCc0Tkp2v8gHKccPPlG5pBdig9hFU
wj8Pv0vfZMJcNj0hq6nVFfrzDcTXh8t/O9RZa5v+5nLd8P8H0dQW2iP8/+diJ3Sq
zsmdhQd8zdgcF45R9YQgRlKdWLuXujhhwMEpF4XyPN4/5jzJ4Wkmxnz3B6F89VHW
0VJPQAUUpdzqWAsRg71/1ECYI7cddDqzBNIssc2DnwBHaHqj0KyLT9uMFUMy+Jcs
l+6W3axJ/qFWlVT7WW6cD1UDjfJdnTnKVXuQsi8iTc3fsBQ3C8kr9y/4QIhgJDSi
ku6ZUfbEr0LU3gMT5ZYASZdyJwxP17VwNgtLH1jg9NatkGeaEhsdJrkI5OWa61sU
HxwO0ezz6r/VCm/lEKQXpRrwBaJ+RayoL9Z5E9M3cHztZfEC5R2x2+0BZ1WOtT71
2R78SAOVTTpqHyCBg5ydAVfEY65iJTirOo0CcZ9dl9NMoAptGRwlbscG8qefHJeH
rw1FRzzVyT0HjusFN6cSgYD/UFJw6+3hQXkFHPI6wmV0SN6KlDUk2JisFxrih1wM
STGTaThltBeG8HV4OnilHxE+KXkE5Utv5jdz2jQVpW8r7BLSsGvvmeTxVUqrO1WA
uXvSaPjCJXnxSrfDB2z2fHpYH43DCqf4AcNcBh1frWXHWZf6+kZ20t3AyfgOAQbn
Xts5ctpeFEjFN3YXa/PvpKFRksM9gPCm/jcnUFZH2MDD6rIV6e2MNemAvgzBmXlb
pOmGIeiqNfoAHQ1qLyCOGO4FdEzNyxjGXrkXBxzJI8Y0E3sxRzCxruIWM3yCIUyu
nv5xiCjURRaJWiLC7qDxmvtaCWMIlAsrhDiHlbIV2A+oxotwJKrfDvmgMiXNvo+3
UqXsPPu3sCg2lG2JUmKjRPTV5qcnzTgFtNzvfU4OVwt+nHZh/uHb1YTQ+jBzabD8
zANESkQ5Pwo189fU5u8u5I+n4zIAeQUp9aL34h2PByYsuY9xKrAEZ8vHWJqtI2Cv
naYhoFD61rb/HwvZ5h9O87eYc7vDXt7BN6m0udjymWGyvUQvD2Pn63H847RxZevf
L3S20wkv7NY++SLQMd/rbigMsoFda/g6g5uzag4l+Lo2CS7A4HEGd2TKVFpxEQBC
BUhMx2g/gOJG8PSzYYrn87+oWFibvOus4U5TuBu0G39+AAMFqiNAtV0EMQ2Yzgci
YbmCD1Ir/4QxTDB515J8O2B7BV4H/IjF9ZkjKCCZRH3WB6BObHo6mcnJq1lYkwLh
u6qahVzsSFCuuYkQIb27ecpp9lZq9xLi0AUZMAZNeXSamW/QBd9KxR6Fy8Y1X4la
+pvsp2IpiL93e1bpzbK/qxabWhznh2FEAV2mbNhsqFOO++amlbgd0Afv7CG1MeB3
e9X2KjBDjnQ1v/l9yM7fscZB3hM2S8W9LrbeXnpjG6TBzxMpyuWeCdI1dfPa2J04
zckY5+irFvoeXKjkW1mXge7td+ddEWe62fmc+5uDdwjnRM9eT4asVH0hr3txt2l9
7aJOZt2MIP5HROitVBm7jHY1Sw6/vVtI+7e5qkqdNCVRQAtJTuUQUP05xgaoKjLU
LAfys8Jek46RM5CbUDGDc/oKWmseIjIF3eIvE0EFa4dqmKy4XvG/JjuWryLoxgsa
phh/ibkgslaacabqqelSJyKoF6q8LnweuMfrLZc2U0G4+ldD/Xj4b51UrXWk+Ni1
I6crxsOTHxFCWiTtqW8UNwoDLSkgzjbQYfVCpUMSux1I8FCc0nT7aTFJ1ns92vKw
g+kk7kUDzA5bOMg4DpBJArUwsKdcPkzrg5E7ybjNvf5RvUxzwFfWH2ijXlF/Hqta
InK5VbhtbX/vk6RQnpwuWBjBC+J7Iq5plkoqrNHhwBEekToxl9uhzukqQk+uLyts
Zkes/+/v9BdXOVZQ7LyScFu4xaGqna3CVkROF0nAfr81EyKgGHjrYd+JR4NeRTy4
NEHa7rlILZc1Yb89lHoltEpsZYH/9TNNs8MEvTR79eZgQqWvzNY6FhlD5NzcE4C7
bPURHt+EamphINEmpfIiso2oFjZOG3ZxwbO/mlaZjbtG4BlYGYIySn3MGIjDNIZ5
8oS5pKasNe1VptRCrfMmwzvw5GQgtRMLnJLGbvtamYRfcibypQ6LNGnoyT1ESVPE
THI0lm1W5rsJoDmA2QmjAzGOZ2y5H8C5iN1Q/hT4xt4aq9fyFYFV9uhMsyLBuY/s
/6nht2p+QXHewmuFKowlpenT9rHT7LXwuWeOv5FzheMAdP4uuDucwjynz1V4vBDL
M6JTwR/njCUGX/7GVfuNMwL0BuKvs9vXaxU+63VEPyCU0Ai7UP0m+sff3hQsEui9
nM0gJHlv/MfSxGG+Gdee6mmvelqNC2PYJ3kXyAcSb1YmkYUu5Qa8g021+bNTT48J
jRiMcdhy4DAyctRiz19tvDj/pgCBxjnctp6eV1yrqkWwi6OM1znikCGGw5n8rTja
6FPvps9UPnRVy3icFfUduVYH98Lk5hwNhGuqBMn/SMSvMj+oVYopiz8i9VkblEoT
iN3DokdEfzjiErJ+pOPnW6luToCBwUyKSap2aw7RScgNDFxJ8KfMxIilIK22pyJM
7rCKR+BxUAvJx7AgJ10fjkZxui2P/+v37MY+CbDzAsQMq7ns2C+8ITjhfqJ7c3sJ
dnyGXhsGVicNZyKwvflr3SutLB/k4lqEHw+TL6IOL6J3jOrMR8V79WI4SaVSvMgf
HdLtzOmUB+v6hFJ1bDQu9cI7Tkg3GI98TpxSazqBsuI50+HYhOyhhLzNcqZb+Fbe
BsIlOXHAR2H+OVIaonZzEmCQmfHqugF1joJK6Y5TyUyCsiy7sx0k/W2xyuPLR2Vm
UZVuR+R2vF9hK3DHZHUn47hK+63Ou4ZUovb1PsuPZQmTBmsi0ZSVckTL4xXPM4I6
zznzWxykfSPf+VlIOz2nQNy8SDR6Y/nu8y/EKEq0Z7Q45BgGpl/pigv9CuCHVpok
WG3dnsjyUsOs6/wkAtzcrvmpg3rnxROjt99b1Fa0XsfxW321rdxyWwwjZ2NpTlP1
bdsXe0JvVOkLKKoGAfGRnMxhs6kZFZX6Ei+0tctagfx9P9K/nWGxkASr506+f0w7
d7vEDyGNoXyO9vmeRh9uPlsS/7ipxFp3QjB01msi/2wFTRXn9ZY58JpArU6GQT0a
LhvtbNc2gs1kd3ieaaSrIs3pyJleYzZ64wARAfEmnAVi2Wt25K9CaIKawgLUMetw
iRQneID0a1QcNCCfzgcGCe2F1DU7+RjsmkOR9PT17IMtg6fVNeMjPWbcNGFmEK7i
eLoJuayk7v3YxkW/e2dfbFrgI6xJxrBXJlDuuHgcr7ZwHAgw9885c9qXL4Nn3gPX
2JW4BrBvnwYHJtyDO05NwSAr7rosTPfwrat+NvobVK+bRvpdC+SXr794bPSrVx/D
hYs4U7jcxBU5hxizwXIQGq0nefVTTn0uRcIQEpHGiHWEgw+pj24NfnxgN7t9IDl4
K+JcwDV1p/yfll5X70YX9sTbzxdGDhBTWDnD7eyxfsmBrq28tLIv2Y+EUxK/+5Rv
OCfXyAX7aEdrCak3r/TnY4dJcWKHmiCL1m8zZQ0FiZxAcRzv5SJjoZEZO875W8Ao
z49ev5YjbyB1yP7ZSpvniqYevdJC1PgdZsHsBXq3FFtsZ2hgU+iUGxsoDmqyHgO3
5DAg8Yxr5g2t+GCXv2KNugijbSTkifNtExTdq4TK5vYbRXLaCt2EfyUJSKlFoiXv
TPN7IJh0tkG4wOL+HuEmscX9B8wbY41yHEwAvyC6W0tv9Td6qeoGIaSMwhukpCq/
49D4OYg0Fmi7BdP1/AHV4Db7DVSN2+ib8WgSbKAHmuL2h4cCO4N2NxwbmuZQ1pgN
5GnSa+tSnQxDaa1AlBhCuXMdTDwBP8dunuv8dZ7/qeRedU5TD54vb3qPIedWeKun
njWAqcOVial2T2XmYEPEv7Kq58JT+Lsgny0GOSr6pCkgN/esK9t3BTU05bujndWP
eqW14fpAo5EAqOf8BX5dyIxbb0x3qfeDlMvIQNh9UyDSjVqBeOJpi8F0qLHAsfB+
KDeUa8uDw2/S71ixLv7cy9Pp/9aTsjxiHfBOW0nVEKUqeGo3nULW6WvP1xxAGmhK
VfzaOarczDEiTprEuJd6Yx2cPZyiRH11jN0SYviCEaQpc6zKh+csHFujqDgu8F1C
nSvLgSkjRK0drHds14AVjLRaDNbUbTxF9e1/9ADCUvz0eVdsK9AaF08dFz/YZbFM
9ZjKLH7JC/KTKqirHMim4+yXxPgG0VTihg5fyoQWiPmc0rpdq1fRnOeAbsVbDy8L
M3QQc+0xP080uSN6ImykLhLSUN92O/W1JI4Efz5sP4gFfsdDV8apZmGKRhYNlxNE
W8ACm6sqfSmB8X31Qjt3UNWqiK3hq29P4y5FvOfpBjajvCjSe46O6Odzbky05jRm
46BNKtEuVuC7xjyfEPgQHyOiUjUR44cPY5qR7cbruSKwiMqZoceRyYqImSv60XKl
/I8+qEnSwipUC1ByfaNqzEjddsn4ouKIYg23+xkN1Mz+0MSkJ83KexwiPdKuWILI
V+Kqjic/vgxkTokxt8EM+KOqznNJ6m8GF1DRV9WCYzTnG1lIdB0D32EL13VCg59H
GHKwGzbgodTqiYSpY4CRoDuRtxhaMh0RTO33oSxqCB1iNThTrUr+sYc19Nrz5XhQ
6NIQxPbcorJM72oQSN01LbXw9f2hvMiClmZnQEg/j+UygnE1/QSEqIi9DCqqo6Sp
n03WOx2qI5DO43WlleYg2NpkTpJtbUasUpyu0evAxWknZElRN0j7ecqn3LJ5S9lz
gpdGmnE6rGdTw3goRcxDf17iMuL51NPOYj456ZwX2q3Omg7cow0bt3Np7VmEVE82
LFpHyVoTx1rTIcqI2NzpNzSeK0g/xVhFRHFiikUhg0rJaMSBb9za/T5hiewlzWIh
M0VBxFxgxOEJyTKW0FGtmZZF9C49BLUC6NOurxYxmTtMOLrv0EKA4OK3KIIMMtCZ
hUyluyUaBMYvVWSykMrlp6u21rdZXBAg4Ny2e2VYhbnwBO6Ml5f8sgsMYC5dHjRq
6qazmPXXTus2qs+Q8bKnWBtyNi/gL6pGOirkFxbLKvhL0b6xELjraxY2f59RQdB2
fkmq0vIFeghdcpa3x4A0tyVxedHrmygUdj3ylpmkuxcxAW2Ar/TIjr1ObrdoBamm
8MJOU2Vqnvju+1PvPdwxkr9tuSYL6VXm3xKa7gORbPLT4Wn9W8oxyu838rc0+iMz
gz0K1cK79/2vWK/rWEmzjp1w6fKPrmPb2Fkfyga6c8LdYgJ4N/ZHslWRpQgjMDqo
pyXeU0U14j36SYxBwqRKA+o2maeP9kbZp4bWwE1Yd5ZgP4HE7dqWI37uKPiEvPvN
AqUGfSliiPSr+WWCPN4gwMCnW3f+1J+MitOsYNR1rUeB3nv5qBR+QyYJ0O9mYTwI
D6L9VVnUPYj+GR8152/SFiQaTLB/sEmeyVVW3K1I71SbbETx411bIB3ICpuhM7ro
kCeat4AAksd3KmlxN8DkRzycjUAUHKuXMrDb8c8qyPREtIaLWcsZGmHMsoVp0rSg
bwit2hGbS55I2G74GC3K/nw1C6vIuykuj6WSJ1bcNOMge3ouZfeMVYAemMEKvWMB
7ctKI4vIwOeeID98Q1ivWD0fAmXhgCEXqc2Elf0xzt+pay7ljtK89S4Vm0hmxnbd
AL1Ir9iDJ/jwNjAAeKjv0kFgL0TPPeKhr2gHAe1Qb8qq2p6XM8gt/iSZ+hrec5cw
0R/MplkLrKAc/Oy8p2aiapQWeNxWeLsnV/thBlM7lgkzMcobZKRFguEa7Gs31ix0
IsJiqGwhA6pWlf6vUEbm21HT060lswKXnT2TacNqQbbKY6UrL8ebDXQowj0ykMzq
HrCONws+54dp0/+waK++/PSPFItLyAGe/UmDbDtqn2y8nDv4QXwHLO4VKSxUwRCs
Qszj3r1+ln89/V3MqCUdbZJH0KhA/nyxaypto7tJinjZ1KoBW01cxSsvmwyd2W4B
fL4eqis85lowr/kVWrZPkKrJI2nYr9hTL3km8bYEPRW8aKFmTx/U4R7yv4ZsKEy/
EIj/dV3V1KOsaR2Dof/QyO4lqO5LqVCcj+0RMJtZJXvvQhwdYbvTjPN+ZRJeoMjd
WlDWVClGSZTU2h0d0Ucz18uvL+X2rpKLJ97Kj477B2TtCeyxMz+1r32SyjWpTPI0
QsgdXcq4xItFSFBEpLKDoTUs9n3DAdFu0eeHOFoMl0fiR19vSU0YHy+KKj+aSHJ1
77bQaev63MmfAhDKrE/yaORqK8GtEtTKiTZfkYYomM/9zWVTT5iYmUGa1cKBEghF
iJVmkZffWYTze0kK3UkSv2Mr05olY8xYXZwj0eI0oDRkx9a0B9R6YLrWHZSCDECr
2jieS5BpjWrimRg/emZ9oYE2RLaqreDUC/NqWs43cMhwYLMku5ahs7O/HnPuF32q
5FIhy6OrVsqHiHuhdn53Txt2A+lH3Eb/UqLr6WiOgubr3WmU7o41iEPYaCE1kzQv
mtYeZqPtgZB1rq0HGxwTPQwLOru7N+QykUxb9jUsI/sy0Tj4B+akFlgxB1FbcJtN
bXATzy3SqBdN5rNP7DvA5aV8EcRo8/arJrpFB6EQ+Fz1hWmucdKFlbjmiiCckT0M
aHQEdI2xoIqFOBiaMbXpX8ig9T2LqcolLsidqR5Q6txnge1nDh57xUdoQhJE+5wJ
PbyUVjz9aEz3Nc0djo9A1ZbCb2HMvtXL0LHmzqgpcpUp339TppZqFw81r9PEfxtT
sJh+scQmlh3R2JQKdoWOHnUE7mAGJCKFS2hohZCvECZ/gN5Rz1F3IyK4qHcrca0N
iPMtN8myaaUpAxTktk1R6fcm83CJg9LIwHDLcbW+AOSurJ/Bisq3KwkJ2MUD7plx
7InnH6JFll8x7in+0GRjj6jLHfDI/s480Lq1OKbEfCZXV2iM/ddj92SyGj13SQAk
XWnZ4xRLMVpA+QvU1Fwd6aRZd64cQEsZ8889FH43J9HDwovUIO3t8Sa3kHt4C2Sx
RMR7xr+M2UTReboKL2Ex9IEF42Q4lgEzmkfoJ1uXvYwmz/IiYIMq9UXpNdC286lO
DvOt1jSDAFCErG3PLcJ9JOle1URZfTPWad+yskbtIU58HbT0LnKHrW5sgBqtD/BA
Rq5eQAvK3FzyKiamY8bL7/t6/esyUmk5ITJ6pbh0+PaA41B4Qt1ydKpaYTJleznU
HdXvaEe4j1eHl+rF33N0rbPpcraNhscuPZ8uHeWQbsOl9ef5PXDJBslEkImwzByI
pzkLlMMkm6JACR8tuhYWs6XZnWR6WOpOGr3lSPssLc31DcXJ6a2AgB1YJ9IuYx5i
s4HR+jsun/8E2pGeekU97VbhBkBSSP6Q2hfRvFQ2FuoKRorHilNJ4v5/ABz+h8fv
vaNd7A29zQN1kt8bVayuUsKEtQzYTy2QqE9oFLr/2HF+FRPj45nm46UIoS5FVjS8
O0FMOUcJ3jtksl4dpauugqeC+wSflfXXgoFC0uiGd2C2vJk9pWcaP8uOTOUuhcuq
5HThG5ljaqHUPqXD/6vd8TsPRYNXblT/59X0kvkUEPOkSt7rznGZkw+bsuZf3sFB
9SgkIhNDDAhuGRg0KI0EcSqN/h6OHyWmKJRn8ExpycBFkgcAgl+JEgkmurHShf8P
x/KEVxZhDCIdDrnYYTzbpukHiGyq8b17SGJE9AeqlSaJLhtI3/JMrTg76j3ruHs3
q+EVj5Ny7uFKA9HsJXP/ORY3i2t32xGlUMLWo+kAmfktMyDJ33Oy+Z7YEFJKOTCE
jV3/V2vll+BJwqlY1I3F+N26oZY+XD2W7OGN4zYGccqR6lBsemOzrhqvC8G8EnUC
kNtGElAeT05iBtoZ8U7B0llWrOKGMsPK+uIU78ecz1kEM5Wss+GRRZ0ZUxEhxTiC
mk12+bM6Eo5/9vmjpHaO479eNyRXEQs1SpBxqFgPBXXvo7eey1iE/eWPa+mXeokB
nQ5y+q3yhNKTItLtx+zYa5I56KP2Gnz2b7taYcpriGZifW9Moi0Ta8t5535zHZgO
b1KIR7NSNQbGb3W3wBCrmXkuCHIBM85eWGSD03/M6y1xwYQtiWapAaigJh/Ox+NY
mWTSMhnd43fa4Mdib7DAMkPNEkN7K1WEzGV3EavO6iO5K3tL00gVzspFmLfZqctd
sViBEyz0k1FqJcAwcYOK6aivkN5x3oe4UGNfp4M/eAN9dqBtaly639DCWdTeVGkk
ZKXNbLzmDISOlMqeNOvFy9+qzSan20/FZnVn4O0aKEG1+neI9o5jWMwOpieybnSJ
mL9X60GUrhiVM0iV9nBkK+6cSVQIk/sF+YQpocQ8sLdLereeikJ8Z1r9HZBWnZdt
49Kug9KtJIf9DSua5UEktGS9YC+PSlRAC4uEUo4MGi0RrAxkZl446UIo775A/KTm
EGg0uyhDECi4oEPTJamIKy5ljRPBXMUMTFIYqMtDVh4+beH3uWr5lsOIoEQryx6b
VTBhKqk+xAjWPmK+0SNGzXCjYdlvu/18f84DDgtBzBduVgqUIv6gXMWFfiPzaTy3
qQM9igkNW07F+N0K694UEQvLyF4wtCM40ufjbcfJkP46k55+4AF/euwBM0/Ltqxb
J+aHtIB2ujXB1qTF08Z6o0bJH2dSAdxYTmFMlAw9ZWEyuS+ktQ/JNpZQMKsIAtPs
XHQHG8jPmqRIeapTBjzOBYqo2zJX0MMdfz7DfYrC7aYLxiC/TGssvXKxF1ID+zlD
V1N5ZD/c8uFQQv3hBu6Bs4i0Lde7xRf32jCfpmleMHCr/cpt4rrq5tgCea3JfGaA
F5kLEYsIGvQk5Lkx1JBdxF8TklFL+Yz5nM7+fg9sQKIws/ZNfI7ujwIHC7ujuBRe
7GABRsKqId+Q5jw56uo5XYQomAIEeGYLfmSzcUAt4sYIqvuj3UUuI+JXRriQ2Yxn
yvb1W08XSeyHuL6Snpd7M3VGYOsWIovLfag4SEvakzyzDQ1cZcYF4mICt7jNf68K
UoaWC4B4jpuws4XbqmGVEh6pLQjS+oRzU5drOEF5GuxzOGAj6Zuli6OcpE2vL09m
MOW2RcpZKltrpr3yqubDIfWD64byUiT+DXy0WRMNXHDQ8xpsCeWKZQprlZGSmhBh
vkH9SlY4DGtDWl15Z/vAKlVFgwgEpA+fA8s/Lvo9PZKo/Dj2AH2C4i5G7HtzLz/I
3m3FSFQCovFMwom6aYWyvc/WDfhxoZS/GiogbV4CLPiOtZa6gxTSG0HFY1VL8ThP
aI/uoHiYa9q6iX5FPgJ41OwmI4tOVuBkEvSZ/IgjUMXyc5Hi/RhR6msAiZpbi8S5
xjFEy+EdVG0U8sc/Z4PbfEWB5iUIB9AJ8GD7whk5XlY4RZrx6egMfsOae2WXsZb/
HfPAy5+ystfFc3Dhdy72oPc1DU+9+e/XRZz2ge5djjJ30UMgNHvDcshcUrEkf87u
UhgyRdfFen3svkn6oJuihZ6MA0Uh9iz3laDhFgapJIKVr707vsMEA4lp7B1fWvO0
9C4IGRiQKNzGVPohiY6V3hhIl5bb4PLV6/aYOUITvGIE10QMoiiQszPe03y+MNfj
lAAf7hUgSGxYgQCAsYc+Z010I07MiQ/qBkIImiD23aGT5cNqARVmWHEH7iknsVaP
U8tjC7Y/9FpYDDz7x/DhXwfSKPIwd+wuFXfZ+Uk7NcHtD+csWubOuTGUINcVa3P7
LaYd1ULK0Usc6Jeo0FP5Z3g9FFtfw+Z2ad+5WqeLdYsiElngkzMSuEtA/QLvLtlG
jqPjszHlqAn25jbtH7urNMfOZZE243DaLw4xbIW9Y2u2xT4+CukDeVn4X4ZP+On2
P/GrlJsokBYmN1rsE0RXNlZP3fsLPywplNFSOAuhL/rIE8c5cvt3FH32kKiKrifR
Nxkd29HIuucZc65mGld/cgzGvUncgMUijzLLEzrw+1snUqMJI4IZbAh5kW/fiB/K
KQYuwh/8O51FASxoG6H5l6k1WMTCtjLpVrM7W32/O4rN1GHo7m60KuCThjBEakMI
Zlnp3iXp/Hy1i3Ti3G5NIklov17S/bjPcbSPBqFmpxnCh5FvtCbBI4Jw1Hp9drgC
62JmcWI90a5CDLGYAf7PuoM4AaoqBmvZkRCZIM/yIidePGBW+kcjEKyZZoI4ZWgM
BZOZa8aTAavge5YpW67tRp5WSQnYEO+ISFPgggyo/qYqn4njyOx31RLD/+kC2rA/
VCYTZOGjCLROioWaE4K549qXLHY7fqEt1EXWl3g0xtuxdzQBFSfG/4BS3wQulut3
LEDpnpm34UsrrTUqUMNhAU1QtgfwPxR9B4bzy5Xx6RLYzE5tZ2AVu4PQw0gj60tu
pCOLYxLvzB7e0sviHVBrmNcmmDh5M3fRlTM2KOZKuAxIwYPwnbo0/g2WcdSh8LEB
cxz6zWh3ZPLPYkNR1V0+bmlNx2pTeTNan9O06z4vOKRwCsLcKdLH+N3U54Rvhx6v
TXZ8YNrwF1yO4/rFTpIIuXe25o1QlLgkjcVb1iAaAAuVH23+qrC2ilty20eXkQvp
CLoM9G/J9XYQSCH6jRZGglmxaly5cpuK1I7dNfLWYvSyEChKptxNPQhnx4bGPGhe
G7BpCrXgXcmnHXo1qq0S86fuQFJtOAw07UV16sBnhTKJ7EEvWw3hSinJm9CnRxmh
YZYaQBFVuGtggT5jUgSWf5z50+2+xLHwnaCNPrxldjTjYT/OlpxO8Lge5xkyN6n/
xMYSyP6138mGcf+PQ31Hl6m+o6KOdFuQU+ac8ELYj3YcJOKITNAry5MkDZ4TbdFt
Is9iT66mQTK6r2zxU0ZyGDIEYcgBGNgenYYx0+Bl0pMGS2Sqz6ksSkVQNckwFQsF
msiNLgOzyvyFD7UuDQC6mmM92TZj/JY6eYCEJXCzYgAe0s6eXvKfPH4zKYQH/UrX
F/srhzZgRFYY6S5G/p2CfP1lU7rzKtUBBwS+REFH6x5ANhlSYEbGT8yADxGO/06F
ANIVzGuiD35vhA4hkdsKqYSKxvsbuJMxSEr+x0Cm/A6kE8l7uhy6I9j7QqmKsgkS
3wvzlbODRqgUoUX2dtTaGbOQqU7n6GdhPOC+bK1OwFNEn68mKZZCiVrxSmToA008
NfuKbZnf9SzGVxHcn6Xv29o44CpWa/UAbOkmWCF5luMtN8dnNUXn0SgCLAD10wvi
0UdT3ek6wKhPv8ajdASBL70XncggGWnwAQbkYc+1+im/PB2Zx9K1e4pIfX2YYfmx
NWJb3pZ/eCGJI42XQQTIOuUNyTXAUsg0sF0Cv4XjRCSZo1JVhXFAPzoIKOnEUzBK
8NBs9MzK5CY7RWbo7vQugNaiYAsFjgaQmXqcyYMC6YQ47Nutb1Gnut+OeFgvxfUd
DF8nCiwTNOf5QCodDfciN3mySW1v86GqVBtLLhuSuxR4e//RT2Q6X2TXJ2IXlkRa
6erHlFGcoyl0/8mdKMMaze074gFPoatKy3YDpO+mRwFrYfNUTH9fPzZ5ukD1aZtB
HeCIUkRpUkngYtE7tWex/ww7W1SnZ7/cx16gcntzki5imTBgLoH/1govME/4FflZ
YVi6WadF4c7F4/h6pwtpBb6a8wnFgBASQM+GfahKq+3noJjZBzKaOAYDkjLnusMS
Pc0qDa0zg61EwDpCuP9a/3nxjteITIUzkKpbOf87Utgh26Yd/Gr36SF5brW5Q8Fk
immQaVXkp9EzNiG80cO8z2xjg7aiPHiRHc22o3LrKhwUnp0PyIzxtgY3AE8LNKRZ
GTR/w5cP6ccg/BvrXjC+DaQxeO463AGcwdHStT5obk0LiFimf5b/0KMr6+yrneWq
JYs+HFISuK3nN8cJG4gq3aUOrqvG4Yxqc7GA9HD7GYOw5+uZQe5Z6Kd6/Mt2fprN
Okz7XVGI+0bM8nQfP8kJLXamm4zvGjWNO36fLjLxnKjkYRMYEhmju/QgAObDnm31
u6DDd4JhKVNcIrH26ivFhodUROhedYvEfUyft6T8dp5iNxk67hptFMLMbq32cGuf
Sz36mectaUbWwmwTNsIU4MDMnbjEgfQr/y967vu2NpXK5v7MCRr0SGxZ5bCDORQB
eNqPS2ONCUWF+cOvgBGQPtDzfMnhLGmJJ00Yh6d2xodnjEVBw/XNmztE2iMwsbvt
0G7H0OvcO8dvDnvgbS/y1PWBlGLiVCKisW/nG5kAljr2ZLX54iY9Vo6Vq/iECK1X
eVPeFAf+8O7B3xUJ7iTNVEbsyq/IxsQ1NXMGlYQKwgMocvjzWVmLfkESdiK4pjLA
epDf2+yTEYPInZg5qVF6zztOuKfMKhLYN+XyK4HTFmUEpXQE15C9eWbjo8yvJBaQ
3vs+97FK7jgyokpdbQqqY36y47nlHX9jRmsymptaUCkRaQS+sL8DP6wuMiydfgBJ
HpoKZ1HZ/Ai/kYnV3E0qwdx2Pplp7Syy2eEWyHESKVJIn47OK4Uu8HkXr6lEtqzJ
sBoMZcgiwMtzUprUhiaRciCqfwaGR6PSAzzMeW5B9lo8TaGx2oS2FkSjj25LjXc2
0bSsdqo981O6pFzeo/S5u0Hi3B7ZdaiYgUJxtoOFDYzGrEh+N5/rJY/rhxCsWEb1
lYOFL/3NLKhKV3KqmfilvOyun6MkdhCJNnmMqOCTrMmsHtf1czY2cRl6gMj0n9m1
pc2UxfkQtyxDbSGRjMtJNGJU2pQlZEpPfGQe+XNFEsd8fxRtZBnrQCKPScHwAOMk
oNYqkmBxOjpe05QIDv2wmII65InBWhOAj8H9sWQ5cgj1qZBBoThMjniO+Xfh9UqT
4QjBU5mo/My3uYOLUTllGK6qcA6PX0CLOCORXtY6lVvlxwYnL4uB7c+R+9/lZ1BT
gvaCYtmIC6PghxnsbX9Oljr71Jonz+vDJiHXygN9l5YX/iQdM+/0ziGQQgRP9pwx
sd4Zta2OvP4yjpqu+HJ3bxiMpiOx0NL9W1hoQAyGrd48noFBWI1v2JpNiCsHvYEo
AnscS8oCajyBpQWsIfOHU0C56YTuxxO9qkcsjyWbt9I+5xBFnveqHTO6FcCIZdxF
vQN6j+/jeeiyYdczvJs6E2vA+Beu5HB9lH6sIiXl7IWd5BlzTqfEmJBDKn2LRNS1
5O0CMgZ1N+RQxuSSv5bELDHrT23USrQrcoMHGMJWEYLyZZ4MX+IgIdi7KEypXHot
LXTuwzUhGFuyM32XkVvIEvQwT5yXHc99WbSL+pW3jkHRDh5kPuy2j7tYbvoFAvIn
wT95B0dYwp4MF7OQbDgty3wy5/tZi+9L870y3GpsYSj3mI9YNr9icJB3IDEz32uD
VDQOVzeDsgwzhZCSRG3U3rZqFjVCUNStXUFv1vc+aHWoZ4CDd/KDZTJHmADptlst
3kaoSEeRbuYmHWeHZ7CgSvsUvrudKjF0ycJjLLBzWK9DlIhikez32oxx8SLO7a+b
M0aHqJ/9nMHqBFzW/ctggwJkdZ/Re+mNhagvQGL/zdyJp+65hdZL9GviNpBxzEsF
HNU9emi+bz0P/ynX5D33QdS4KfeMKusdfxLEtlji07QrOGB2alNxYYnKidoeTDsn
zfxx1m5XK8ZqvyKng5EbI0+3A/rEEp/BD/SVu+ahyi23VlLR9fEPVcRcgob8JY7w
PODVjTNxKWbLMbCzQSvjV/ZI5kvl1v41yA8mOBLn0NYV3YRx4lFfnDWuudg89k39
TddMXvvaXOQTE1yNwFgjQKhMi4ly7zR/dc6kVT8bz2RONPi04zPM5FGs9FtXRN2o
bCFHd86zjsYNkd+QpWNSu2tUfo6oB/oWVDpmTxOIX/zoXl8iLZLM9cv5fnWvgLt5
XK4EWeSkUzOVca/wdkTed8itddlsG8xq89BCtt5oSmHWvL2EjT2ug/vybeguIYbs
D7RYiagF15jWurpZ1Lq3g8N1hIcVGw2S/WbNgXA90nDSuKkwaI8zksYaxGqLZD9j
3H6KksCpbL0WcEmDEoipqXP9tuplEmh4tickw1sT80dQDL4cUbCeetlKvRun3X1x
wFN0doogt0ewzo59MPelIkePFSYWR/L2PK97pqV/cAv9f5RSlk8StFr6h8HuvyQs
bPLzJvg3KStOWpTqikQQZ2CodjFogiBO9vmzdq302z4wrs2Sjg4TnJf+GKDXYQEk
cmGjJz58pAH5GSFwenjqDVkCh4zQT43AItkhghtjxWXkYDbQLNUy5hKZF6fq7vir
fUIdWKK+9Ucqg2dSQHTa+97CG5JH+e46nuiBaEvkLiXVHw8pBVD4/zXyao8A5wWW
yB++gqRJwEUIF6eOHOIfflpRyYQlAaaOj2VtbLNMX9rBjc+g1tHjHhmzwIELA89x
ILrHphoe7AoBHPSWwn0g64xsI7fZj7ofJjNdbPGUKvC39xpMLqw2/0Tadmxuoqa8
xWPRLh0Hq/aA6IWIqy5TjfOmzAFAqOCMzFlJhGBmyAd5jkH2wQlt8zyhXCiWJBzL
lblyTMkYWCbqlkSNq34pmnXLJ9UhmWyJKp6MWX2ftW75aNhQuodsdAO36AOyBewX
qcy+ldJN7m9fhw+dBG6J2yJvu8GOczgeCKgDEpQrBmEgnGK3y5OFF5Jg7E1GkdZq
ZcXy6pqeZbS5ETRI79Rxj1rN07Q8Y4Wvks9EQMSOdHMt9tk4rG6Ddvj2kssI/uCi
kokTSVvTvOuI62pwzwgjJJfYCn4ns09sPuRpRgg9/wC6bZ5UWk0a0uMXJ6CULzVO
Cc+UjnB23Zougk9MBKffDXpnx9A+ZMi67wtsWak59rsa8JutnTtpYShyvFWgUKZy
Zo1L13GCgHxhXjx3qaBvfKtE82wOdL11F5uZid/ycXH94aFyYWOuBHzPaG1Ieeia
TCI3WkebvBBh521CI/FCzl92/bbu9X97oLrUTKSLQayPwtKe6oiGeNXpDv+/AJBp
fF/Hz3oMlgDyK8cc9z4fPNj2PWSTXDYnkfu75M3+vBHsjFz8oLD/XFL1GhQTq0Es
SzivN1OWAKXO05o73v5LMoxgmUV9wb/oOwPShtA7cLId8xomAhRnkNs5jGO0unaz
wIiev8NWM2Mpo/3RIFGKngO2oKz0F2b+dPVB2ziVv6fkU31katoCwT4ihzOhxKWE
XHwwxgG+h6EM31nJFIsbKm3/xJWE+bWsM5VsilN6eqwN+Gp1+uELDlFCdjXgS5fd
oZVTZGjwpYzGFGOOijMmGEMC0iTPaJcnDEvV8Znbsjd43zeGthfeXnchXLmxEpus
DFAfaz7nWvNilGrdmpkz4QtzdAnWq+HVWhY61c2LwLT3FbIgxUYjibYhKQJPNaRN
h1QSofWdz5im1gFuMaO621ZbwVeMsIbJfLuO873ywJMyEk5cEJQ84W/VDIjJdK2R
xQtcEsH/+kUBxfNVHEdBGau9QDTB5ow6AdZiqL1i48+VwzQbRXlfoArRlv8z1s3z
Rjt9Zx3jnQM4Bywx/GW6/gYON863jmyQV0WXooTnHKXAZFVUXqztjqt4KCEyplWr
bClNDP2+ci4wMf01kQBI38YRztzSKAOXDd6v2u7TcwnG5HNDyhqbQNCt17UzaZsz
WI2QocfCMyHf1eDmlPrJ5tw1BzkYGxpDn1QCUfkeAeKwW9rZYLlts7/xIcUv3t52
OHJj3e7vcgRft3l9vsEqhSIh1CDYUT4lPjJBctfb/XwHWwYw+9/wgMOdp1Q6fOJc
AC1+qsMwHjlWC1Asv3pHuWKzCvvjLSCcY+Kq8aHSwP/ocIT8DzWRTgHlyNvgr/tM
ypDwvEfQeHxSlIc7BxnKz7tcLKQbVcbkx88BLBRR6XRp0AF8KWXSS16wt+7xJiYS
z69Z6g1GszVEqSkRjUwns21yvNr1Q4L3TMvNW1ciDHJ+wSVexYkG/wIwSz0ZgnJj
YpnPhIMLYu+s7Q4AEXmdIwbYbBa+ZsCLDAcw7t1p0FkOV7DILLTFajkYzvMbq9ZS
3HmE6GXXH2JzEos1bGTU+n8rpTtp8NDO6QbBgntVGc3kzVtx9LFG9zaBzgl3xaYF
5S8BTUJM5ex7JaJnzuT4AKy9clF+shLRTO2HIkfPMPOk7Fqv4YBiglqCdJoxU9vK
EDv1Q4NU10cMetxqB6c79GrJuzxeEMiJCk+zyXvd6otKFjf1zL2rNgvg/NbzmJgU
58GGFQ+wAzFgeyv+SJTLys9vCcefO7/CucuNigLHYMHB3GGRBA6QlPdKaYsytGAa
V1V9Van3DgW95Th3p8csRlQlM3DHL/FnfyT6Blggwd1FJYAF9b2WqvNsxq/3X7Gq
fq3kBbNG/SH/i9DzvyXC3jNuI8r0NoLE23QeQjxQNzq2jLTM9ITN62AjmUcPoYYU
GM9NYFpRYcO1TJW2Wo7gsKQISj+HgHt+UcfTZusU0wNfYqpbQh8HMwsyKkcujN/S
ZrIdJ3IuIrWe+4uvMYNjECdlDS9aWURBWHkXi36Iu0IOYp5EfqwTPQ1peoTrke6g
mNLVWTt6W4hnFKFG6vnWQXyS72YJIzufSs2Iy/GpZ1p1oKuBK5Df4LHy+TPFvPzp
C65Gj0pWqnV6rZaIK40KICXUqsFEJF8TQP7JNlis7SK00PDpmB3rxch+6ydiGVD+
j19+LXlWW/BGmAtimIpSLb6miFXU0oDxC1okJuS3uwSb8Q4Ejj3Fnep/GqEjTkMn
nUGlx7jf8SGBc0TFVBviOuKbA1Z4GzBZUbXLnFDFmG0OxaoUU1FrAzUrAiscGK/8
VmYe2j9Gp3T9HcRn+uhWzzUR9v/L0cZFC0czx5GcIwvAVinM5VhU4GomDoxne35l
AZsKrDo0TQw4LGhLvgvQNCdlcyq6Dw6jJ0Mi9yADirdRPWma6wl1R6reh9pmxObg
fNFus45rhwT0z1IYmlfXQhQUCUvRlm+Db23GzABh8Oh3I16+UtLfwKiJu4u7cU3V
rd8FbTdfDCRz7gnUK4LFOKGhTldBHuCpjvMZGs4btXmlBrSbU5mDfVvgN+CQSh+W
+5/BtM2MzaawCY4O3qfz7Q0EQqCAtE0Wq8Mo5+wzEht0Lft56lnw/kmC2ntBmR84
2pC2o7Tx2RLIb6SVW247txbhvvjeKw8X6BY2WGRFGOdiXGGbFnemtBdP7y56ZlXL
omPDf8gR/RJFt1BJMYDWpptbLJjL0EKfjrY0w0htvmx/C/lTFwt+3SqeZzVB26OF
6BcMRmIZ6C/f1djSHRIDy1qpDV4ORALQ9gJByM609QPlSWnjNjO4S63b273haAO8
uPInqsMAkhSzlcOAqeGtGvkZMDWcHEieYPbJD84KOKtkI44y427LPXJqRJbF6BIw
frAjyUM7kt+SjFY+w1UvutyIZfv8VtuN7ZTYTAImYIwK50hp25Xdr8hepoRTYETs
xpXjkyvS0y72y+Id8DlthRBIM48dGoY5EZtOCvxTNM2YrRbusW2gRVh3KuM85e1f
4tB0wAWgMnXorUiG8FLG7f4rj1TyAUy46zTf6zBY7pJjZpJaOiKYvddpx/K0stBS
69CHfJ8hwNJBdt/dD2gUEH+0rK7KoLWdIRamgVxBBfAiBignQXUzmB/vDI84uczb
/f2cSwjVHE/dsIkJNMGdocBcQVlizdr1D6GLMtHuJeApmNlr3XyIHqUpBQ+IdPxr
VGj33zzs7NQE4mHGOD7+no85GjIoxZsn8R3SyfmBKqqdHie+s9l5RwHvdgTcjxtg
Z4vdx6lcJAT6xnz0/8gFj4VfFsltdU2p39LyXawfuHRmH75QMT1D4hL4fYxSYzs9
/qs7v//V2GsKEnajxPspQMBY1z+Ryc28tlv4Dw4QhDxaWv+mPGbE7csxNjDNG1eh
Bd6z5NarLqkmjUxPRsB4TcEuDBRRHRmjgkER2Gi618LQ+XCcewCk8u9tt1DxsPNX
jSsYTvzD7B7V/sulvCvgUJVClkKmtMBR30TGKkLjJcZpQUJFepCK40y128gzQLOB
imJRiICGxTK3gVxKH42X8Kx0Jq1ScTho0umyhTGlUpbreG5kVrHfXxDAUP7BEHRJ
nh2bA8M9PtfuG5YYcivLc68AoiN8/GAEFM+kokLiBC7sXYnTLqatZ16DTBPoZVaf
6E020gd15sPPR/0SvK4MJPCJ2xbyLaZ0AOtd5XA/vkSuVMFojSuKsYWMrxYd2DxK
UYsp/umYj1t6atrEvX50AN2V8U0DbjSJQUbVWS0JFqLMnGi18f2Ba2Tq4j9e2rR6
Yct6R4cwG6R352TI6iqxXAO1H81nTgiUindNfWOtDiETrukFL64mH4YDNbOsc4D5
QTp31zQNxOvk45hsnqNioz1hN3Jcrz2Qq2PfoaqxEjkGuuXQbK61olnLyucJR6on
q3e51Z+H2AwUpoC7pBiTY2GiwCfF4MneXmgbjsEGynWUM51sAliVTVjL6KQ/YP1j
USS1yMY9q5k7zcTokTo759wHsxBePYymPZUv1PzPdPFwhkTxUF4irfm17ZrrnM8/
TSeyDeQzbnzi19E4ZR4VxvPXG6uv1BN0AdHIJvN+iR+AnPWwNlILBO9SOyWZEvap
eZNg/Q/3hvbIiPRmuv0Xcl3zRdL3LLkodqf19yS8YL+TE3eNJ3kqTNDzkvRukYxS
mGfcVRX+Sj7Ll6x02l/8I0PLCNzJK30mE7Fw/lZnfOmzebjsWsU54C0bc3X6h9F4
J38/qSOisxnZW7BhPvdQK+XYo00j3DLaHbGiaAh/ZMYF7/gkMoQzToqYJnlljNR5
hbk0ObWvF850R26b6ablZql3wGMsqaPqJbZXSQDIS7cC5D6tYj8cuEa3DXtYSpcu
58W892n9fDLNvMUVEI/Abj2zm60bP2GxY9C3pxmwi5MXAV/17HgDnkN/4gf0/i9G
sRmJtf420zyi/d7sNyUkIhD88sSkqkiQvJv4x9k0zkVvryTZAVE3iNm+q7QOKwiu
rdv4+c9dtglwWvwtaKmCUBNmZ+i74BeSzs8EBb+SjORyL+S4P+yOY1xWVdf+VfUz
GLRz2223rTOEKyuqTMALdQql/xGc6EZdo2ePlDcQsjgrt+FmfCDZ5cwvPgTvTl40
qriA5gnRbiPx4vp7XeiojHl4REND7A2z217qYCPLMWD8NEDT33EiDwMgOd3lzx8p
XSgjmNR1PzlFXA0cng4I8rNDfGnTze02zw4svY8qOqOlF+5HYUXZ9p/DO1hnvXtv
N0YGgzw8ohhL+4a5VHMozUDP7xA166AQUcdE+IvjC7dh6K3btLeTil6KEZl9EsC8
FkCB88MsLTEswJatf+T6iP6nro1zWK/yoA/3AHNm0JQzSqKjuvqSIy6qp99NoAE1
ayq/oraixXrSIyGi6FSDMlZe7Gv/gVy0Ojl7TjpFew73LnIeEhYsi0v7N6PB1kwA
sj0rSvgo5YEgSdwqgUZetyK2emfuMTzwYecs0fc+aeKi4te98sq/C9gSXpRl/UH6
Xf/7+Iqv5Bl3oQoaPEUd4AYwgPyiBB0a0o5GfmbgPPKXIoaTod6J7NJf3qvKYmt0
c9Cf4xXf65ApzklndMZ20fwyO0xDm/jTBCzyOFvfW4BAFTKguMdY8Nj+X7FeD+ci
VVTOagA1RJkRhcuboDn1d7w3WfP348WdWPZZw2V1SCZ4I2NrfOMyLMJF+W4RW9HW
KiHmgBCAWTm+UPmfNyx6uE07LYMc9u+0by567l0649OUbk+exdzLT2p/CazsvtxI
hd7OF48F2e/ZdFZFOyGRQXvMZGi0l6a5ty/WsmpSL8JQp0Dpkq0PAdNHXBEBgBvf
FtwYDnipMnoyZeO5vKxp5Yel0espUbV0AN9yJEJi5Hy/yDetU/fi5IpwlhGHGVfK
OyVrgRQmy+fg8Hb8McsaZRroGVE6u9a7auhz+S1+gRKSkjxvYw/dcf/1VroQRUJL
55QlmC8qBJ/oLkBVa7WVvLU0i7MxcLNDg7WYRYruSGNFqlS3sVnh/0p+Rf2SI4Jy
yyeheuKRsac6EM0v75dTvyRHFpcD4SpsSy+DYXIFy3cp2lq8NK8sNm51sjPL4jyt
MlpqKEJwE4SM6WvHcMX8oxtUtcPCS4EWAPUlvvBWG9+6Q8OOoebunlTemn/RQru7
o3Qkd6pC1hcZzKsCOp6rFQyD+pBq0eXCY7mORQdYkwHzSUwTq/GfMuKYon8vTZ1o
1M0yrB6EiRzDPV5HgWfEmEvv5XdR3mLu1YksQOxdg7DkS0vLPUNaYQjd/HTjLxhD
R6bnH9FPXwB2mwH3Rypw4WdqiLuqls5LI9/Wuicr6WG4B8M8yyybciy18fTM5sH1
GQ46+hioAVPL1yLb1gZ9W9PKRcFk8sSIsz/KzjuoeqhrrtZ6aq+6qT8n8JXiatza
26oyvylgVTo09noSkQ6UHPQRX2lRrT35b3fPEyQwZ7HX1fWFsB1KZ7Yp6/JxsBJ7
SWxZGhufEmHOSiFI8MCdgYspjqYjPwv7KFRw8xk2NAFVX9y1VpiZ2KWrd3K5IwkO
x8FoYrFpeGqYITMziYTx37cuWlbCK2NSvMBZuwdTM8nWjuJBocM7fwZKpcZe7Bxx
WjlQpiobv74GiqbQ60h2lH8VEnsKCdQBo6zC33Q4j1o3P9ah5irgkUh/9PGYoXYk
tDH5Y48SHrwZdx9VF01aX8oWJWs6EKFYhk7iEQkoPYJ3MFWua+2luvNLegpUdL3P
q1laXNoWJMSSWfVOqFUjY6avJQgHVb6loR0MZ6K6cvccVMkAOmEOoysD7GsdXzb+
JoioPyKFVp1xbnXBa4QW10XLTRYPi4+ueJw1BA8g0yw4P3xkPcqY/bQapzE7P3Kq
syYGob+u60DmIAEf2NIdbvvfQWQaVdnSrmJHWSvNb/0i6g/tcFjhocf5H3bGdADQ
NQDcf7UbJFsNaYDSFk5pN70qqCBR95ueElxANlSAoC2f18g1aUzl/qBePGRcOUBk
P0nkOx5+kc2+/yiZ8/TwZ8YKO+KkWppqxps5DKoRyzxK4XjklR9O8y2KquTJG8Rl
qZHcOHXglE3D77XdbL241KOdTIZMSCpktDHtYdSRSSukwvoZ8QzG8eD6EvbLR9/R
Vh+AliDs9etfacG+Aenc4D+bvpJkz+VXvG8nVoENp8QDjRR5qUnBHb5nzavH//GY
d6OCO0UmOk0oJJ1fYo+XV0efQTBvNW/T2QtEv+OTDIi7vEXP5Q9AzqxTRyI974x9
9s+8xXchwDul/oHiuybufcb98lfbsKYTcx6vbUfnnOS4E5oNMMCdrswJlUpy/qMn
LrE22AXxgBwABO1uKgLidu+N/DB+mPKNexd6i22YKv33hCm7wYDZxL78OPiprSVa
5aUBsY6527wKihyiSIWUBt0uZDP/h3BoL6EAhG7l8m9uFaeItFEPxIFAGpw5uQPO
nux+RnodAAo3FbwncYbrWu2leq6qXwRg4360Wy/S5l5O3u3pLkDqYTN6buvO4orY
apV2iOuxM+4IRQ+TyrUtoN1PGzcbmkl9onlDAoJpp9GNRBmZACfuIVS7ULogtlIZ
x/ehWNEiMyOS37mmvBkWNrzvgznFSuAeXJqk0YeNf+KXaZVMLMPqKUKBbv7PZT8B
WnMGWd6zVgXpCqdsF4BHEmNblF5gFgFYOPOU0/+VRdEIUqLFkA5boKP6YK+GmJtC
WVVt0p9ucYPKBsfZ4QOBHqhS2eUhmSDyNy+Lp85JaBS5q7EBcpbObvlvKZLLy100
WTBab8talFJBJcU56PkYo33SOg23ELHVYaWbL5I+VZurgWj22xcS5z48D6D97FX8
v3m/Ob7UQfNN1+xMQsuIDKOa4jHf2eSQN57ZbS3+G2zs5gk9mDwY2JvPZ5tHJVUQ
QOmhie+PdSF6fDdl2L3Rj4JKOL94NAQdOQCNSnZCA0IdO7VDZCFLTDptdaqW66MQ
KgU2BFJaUDKMe7qjc325KpMCfILm7fG866afmhJ7uSq8QIzGGGfRPeOCNWUD2Bjx
15hdF4HTIcoRbwzdpXraqeSrJFWuOVUyrKOgytwIR1/XpcubnAkXNLKsJSG3fSaY
k32Av522DJIz3QD/nOMAWzi9OzpyL2fSu++wYuF/rlfJO8gSJklzlg1W8rdDUKiX
oj2DozzEFlAMWS/dUArgKFJXiefNFwCtvr2vJUo7jPNy6U4WbMSySmYTmIl37zUX
kciuejxeSMeKRzFx51rIDcdcHXO/MpnHJXfmEgcp23X6RUKovx2W/ixGV1YIrT4/
C6cBw49HfwFA1/R1MnYa6Eqt/WdC3P9GQXGDPoN5F6r8mVGjJR0FLsLTuwl6xxLz
RRaJy/EWviH2WPcVagi1H/8B5ts9BEDzDSmvU5vjSaIRfjem16+4AaCef1/K6pk2
k10oggyt+mYYOfihKRc638Zt+QJivqr3bQm7B5rTEZSOOlT7iURzKnB8/vQva2O/
8tcXqeprDGldxSiSojIwa8+s7ZFy6mDIO5CjEeCxTC7mylklZxDMEBeQdLRW1MTV
Z9ZzH7G6M1e2yguWBSNhAqbwYgPmcA4PNxJlmVQe5KnPHHfh5bnKZP+PO9/9Lr5a
G0tJqk7/9i6qU9OBnw27b+BEsuNdWqQkWPy6UGXfNh64wpe8i4sXgnsZgIss+/Ry
5/ooQbemlo+wtJeYE67KiLp53eg/epLDiF5XOo3dmYTCtGbuCTdOcPTA0dc/k7HZ
k0ChYsE91D10xJN5Fv0VA6JqqziKx95soqIPksSH6PowgnDD7BuG+N8wyZTssw/h
mw4YxB9/9YGLxG7UB9t/Sw9Kzz3FaRnM0skZiMEGr3MUMTUlMP2MYwTV9mxTlUTW
VhEiRJNaKlZWMvtsvnt2jT76zAoGHCZ74VXeXy8dEMP6CSO633fsOULsXZYvOXWc
uwojBuzOAN7VQxIX3ay71AC+87+NOok9uuqkufDBWXr825UyBzGxQSn2epngUGCt
awUICQ1b/9jFkR8wYQqxyxo9KhV7WLAi/dPMbsY2IXKoYaYDpbTfGue8Zed5VtKq
6SxmAMVrNFQkavj0mcet/5ueYEGpbSACgd51IEewy5Md+lOuCWg0Rt1oqbumv3/x
sMNwVKwXqj0HwlQB7TyWI/Mgiy6yXuS8TxKGT436+u5I4+RWG8tVvbMgx/DRTyEU
JC3/ILG0Q/YdW9Ff/53v6FAsUmv6SLidmSkeYWza0uOmEmlIzl/Grl1OqokspUH/
bB8knSq4xSjkZDbA3icsnYtn6b2Kk9B1k/HGgVmBbtD1yboRmpR35S5g23JcKvjQ
pYB/YBUDwFwIVC+QMpDyGTitmCkJfUng5HOEHK2NCNHtBgyawWdPGSC3HodcPQ9X
cZQrv/kKCWJnPrkvNJ+wOUbRs1up2UzzTAnnmk3QMio9QhiWHVibqlyiD5aSLc7B
vg66ILLf+TR3H9cKaW4q643d/toEGWMVYgvXAhy5/ju2YJsYqaV+qwZqnt7r3ams
EJc/ZbVLbvtuCAecJJwd7BqyQ7Vsksoe7F5Zoc+yuRmWkTAZnePpsD/k0DIOEvav
mA2o/meuvoU6AQDwq5ax3E50Y8u3vp5ztb8cWQ7LJoxwVk2fHfFHXMsZKhsRaxme
fTSGs0tBE1/zDhZ9IPEVffieHU5iHFL+gv5vYu82jNaFikGoo7YDz2auENbEqxLV
t/2825xdGjM0Fs36FuVFIfeo/e609yuQTc4Bh1jNo0ZwR8OarNL7W04DU30zw1N5
dFv0CvTrIFjLJ+3YUdjPvhEaMe9mWeVn10R7tUoT7gN7z5brtdHjpXESX7Yu+og8
ktPEQZMFONlLg/DbJBpF+cKHl+ix1jciISO/Baob4YVYHbu68AQccVnHtq6B5eMz
u1/pRd4B0QXz5A+R5bZ+20vJ+ELc7bdyCV5JVrJcv/XQP3gaLe5CuWnqeFTzVY0L
DOIUvKNxTRUTMvLGmLhDXfJfbweM7wzevBCR3yB63cDg7yj/ZwjzQnGTd6CPpy1o
cRG4vOtOqBK3HmNdrL4B/7o/QpvsKslHJD3exrwcyB08GUH95ONAnSCxZIg5T+ln
WqGznvei0KCLBGmrH6ES1Zw22M4Uu8GcNwwNdddjFLHmcTQozn8Gip71bbWPjXuY
Qp+6KCrBiQQBCiyi/1vpLp9rrJe3k6aZ4nEFkY5d+CGmeiMPO1kBf8T3Qa4FTADB
E5uXv1tHIaKPfF7Fm19eF+vJTeAS8oZkC0A9/MMYF3vdCu8D7eR2/R9QN5UOYnkG
oppvoC/HGig6f5qruhiWv2dXKmU92ctuDHLscTCfvOVtKgBq3BEhByplENoRgAee
vAHhA6L0p7/wCYj0LTaUPmBJNzaKkKOYRn5Zpa2Y6mcrhOWZUUOj0k73iIeKnPWa
YxLUdummWlQGvKHt9VwRwUcllhUQJjnerr/L7vixKZ4m5ybPoMduP33Ia3XKP1/4
EehQkPIGSo6d955X0Mhcg4yluIQpNsJA4chFzAu23JT8TXOzWlNOMRwd+t9GQuI6
tzO+JGXE2eelNmKl8SUUlIPaphTGhVigI45JCTLtZo1vsAc0HfGtOMWjbFk6USpP
4vmmaD49bGAmxS4E5GPIfRoyGjf4ywSHFsZRZ60ruu02LO0tRnwzZhNoyuTvvHGp
wbWeAPeEDwBdrHTCMdRT5nJSfAvd9SMIaUIFvf/mBNIxGRRltar1qOW7HceX00Ad
J1gK9Rsni9roszl9EDtfJSAcLVpJE/qv78RAZ8BhhqO7LGfsT1mFX1upslmPmBgw
5ty8J03rR5aLeVckguTZR33z3T9oBgfekE5Vflw1/drLQ7JwcKNhj7Wm8ntH/Ee0
RI+gdvImy2n2o9Helg7/Cl+gi8e7JVMmJhVujyNEMQZ67f1uJr+PAP1B16YuKOBW
PuTAaYM8FynqKaqapNWS4HSqoO5Yw7mn3EK2TzoFXs+MSkruTuoHYOARXvxweXZJ
keLLS5IJ68YP76tADGHs2DN47F30Pj9vBNfs/Dsxj8E7iibL57ohDJEDKaGj6ZIy
XFr+ZRl5C+lPwlnzrVP8AAIjR4lwS+tZiSLPytiYHMSu78m6U2zZwEhITPBLVyay
l2cGp5FVwBVdmNwM5fhTKB4fEfkPfvu0XVdSH4ekuGwFfFfViIB+D1noU038MSEl
2D6+wKJN4AoFRHdb0F/5J4BZzTmljrsd95zVIE5m+OcG2Z5zARVlxUkhnxv8jH1G
WCUpRu0Y4Xdzpuy+3s5yGKRIDj0R+3X0Uk5DFh8vV3Blp+n/7GNNTt7lb/QxUddq
DV0+sLGKTRJRhIGgoktStFPFXysbT0DBp8lRh3xITp6ipiV1iGMD2z0Og/BeiApQ
Fy4W4allCaxsvxIv2m0uOh3FzumcBZuGC+cB9RuoJR+1GloUgDtL94DxAYb4/bqy
NzZMgyzYib1THb/nJxglZJuYHnhQbDqfS7DzhQMU1STrvShFRaKEkHyDlTwkJXKv
9Kb56W9qdZJv8GopZAAk1u9LEjPZ2p+xBAqs4YCiURB0eqEBinKq6spT5YHoCVfr
gCpckG0f2YBZRjSqSkivU1QiTKA9p9zaijxb0eLdDqSI8cq16bCWwBftrXdB04q3
sAXvloa2WSedVs+KukSAdHhbqUzY/Br7VJLLzgiHw2UUdzTEyMx9NqqMKhek2pOv
bM4OPPKC786cAQuAaM3hKsynvUMOgLvaGqxYBP7mB2p4/VfFiYLtUegLkLYiw/AV
RF4eGK9wg/HvO4fP+ksD7hlCjmyIwZ9LCyiQjQ5s/E9nK0MlrT24MZIbQkTz/Fjk
yF9ZgVfRtyWWEnvhW8y1vRVXmmZJ6orU622/sf2N6cvD2nOwuE7GvT4reG8LtvaP
b651B4r6zxKDF1VozIZBXxq+57U0nQW2O1ONRWAFeV2AJN2KByea/46CSSNOexoB
kRbPNyBizmCgB4flyJA37xU3M9LDppm0JH9KWogigQJB/m8jgvoVbJAXwMEvWZF0
wi7D1h0k3QwrWZ1e8J9ogNLEszEyuVL8PvzpXaYEUomlIfv4VnELpctxNoVrahuy
mklJvb4Ig0HTGOKfTPR+WFgwqzucuqn1fkyxWwiUS6Vfqh6Ol4iYOnt5nbxl0H7N
RUUFphBQ9mW9sn+VrWG6J6caFXXk/KGHV9FRAnq0iul5G7FMEaZwFXPye6g4vGdo
77TIS7IOL46ucsQsAQtGMhsfWdcQ1TP8VKi5RW5j9mykEScFurX8n3pngQIOc2+h
3/JDEkeFsTghiIUFYfLCbcAV3SnoPcQJ7xRKYNl18xlvrYy1gCLo4jsdjwxlUFKk
+DLDVAT3UEcakR7pT5gseAkTsiLutm55w2UtfkB9woQ5qlTtdZ9RQNxyC5rTrOFO
3OMy47bAXRCA4hQwp6vcOvnofynCGygIhfwc0eKlgtc1T80Nlkq2xvyX3A0kWuaH
z5y6OleetBaOh5+8HYx2h60CpGA3T2Kq92paV29UvTO2ksxBPXGFAXHVVXQA/nlE
KmKZn3DuLqFwfqsCyVSpDLsiCX4qK5q3PY0FaAxzqx59Spbhmh6R1nRT4gbpT2Ae
ZRsv+mivxNj3RWcqnZvuYfwxg367uTs2MUvI4mCzDh3IgDGoayn192C/Euylt9J7
zekbSIiLgPtGOlDm4sYw+Q0idsGucR0ps6psfbljQWxajoOFp6BzSy3DkA4yX82j
2PxySz7qj44eiytNTMERzhpiAAlpdnYXShm/ECqcpLTCQ214DbGqJOzFPMtQCtGx
36pQv1h4SDqZ1sO/oevz2K888ZNMzJ9DC+WqwHvB03CZefJGoAUj9drpn/X1/05T
I5UTFqtprEN5Eepg7v98LmBwLPqB6enZeIhhwERCnu7ZPOLl+tYD5Hveb9xrdqon
fDrJg89W+U1HZGbIUL27TqG2WStisF4+j7Lb6bIhtW+tr51CAtVTPzAUATpEHCAB
nCBkIWi/t3SpNFeR78btcXe1bHUy8L1uwJqYX/0SR9WrOtFbvoFGzoKDvTCTwKkI
RzPCxyXb85iFPEN08K9swsfqyZDvBQgHbZXSebKy5w3UXShAPKwAQsrUVoQTcXvR
Zx+e04GNSr/HzQjwUtNVYSQcckxUjl/n12V3C29zdMgWVxqJULBY9GZQOAZLY1Eq
u66xTwjereU0jkdR1M7fH6vCiU+rPMtzvY4F0rtv+kDnrhEKvA2VrAZc6A2yUrZu
LFyxCHa/yo8VdzIW5L/+Y008CuLi1zPrtbB1DQw5YuGRhkWmwXVFX438hG1RydBY
WmLkddUXWZExdRlIVmqPjdBSHFjwD+yKe+lShTRMD5LpOO4Kli+5TJuuE5/b200O
fYh1+gpyXFqq4bqDpiCNN4L/YSTDK5M9BF05Wr9jDfped+JutqtmOx875DXij3fT
E8Yt9TcDSL+G3QBmbabIeM93ox94GUcnSM+e0Ri3Ld7RLjr5dyqrdJjA8kjImpPk
2ZjeznywAxMmDFPmVZGueByfZ08CqsVPSTnHdF8Cf1o06JXGwTrSoIWsm/KkWTKt
feZBOHl55uS19whrhGDbbv0h7e4vR5+ZaiH6yZnYvKt66jEeWIwjGMpqBSSD9gAS
gI+mXlSDOKAXhhPorN5AuR8byOchnHRhlVXfAQRj0+7Fby8viZJIfPZLMuTN6ZNg
XjH8PuizvOg0XIvzQFgAxZmG9NlgcvHsZdtN8Sh8eBE+jbFaZiZejN93rhLOB9KD
IqcYaE7+MKHNNXyflW1/O7eNRj5nMZI3ZYs+S3vBvAkimbhPijntNqhQBOpy9Nlt
NPM+niecjxk7Ab5ZchQYy6oh4zY02HV95GUlDRtWob792hTFGX0p1ivp6zY+0VQ+
ZavP21UJRjJSuRYQXsmpxbDDQUZiNV7jwng85IebsJ0sXZQgyU4wQ7Nh8Utl4ISp
+QXjyABktsEQsV13H8EpQimRp0A7sDzwO0RTyN0vB7RCkPSCK6McA88ZHZxlZJ2T
Gm89uacxWxZ0rymojqu98qglkgnnoGfC2+yVBupU2tze51aBZ9US8ODA3hzyyVs4
4UHC+qmfqfaIEy6WHlaT0l2bIlIlLnerMLxD+DA2FjpsPmtAhGvvwItSigWCw4Y3
C+zSYquMq2K7OAWazEi3fwZ5LzgKd7FYFx/duXQvGYrLZ6r1XJeejsbEqrR2PeEi
pZ/hG/UKbU09w6IAX90bAeNZqufH91eIzjG2m36LjFkTIl5YK69xuHmlo8+uWYp2
Zt9OazNUss8Gf6JsAMTX9yEyddC/5fiIggIoPs9AignDLeLbz1aSQTSkrZO771pF
Vajx6DOJ0kW4pHczixoNLNn9HXDSUs5wR577SDXA2qAA2MX7D3rtYUnzyX/c+bMG
p3u7JJxO86iJ8Ie/tlAtUN/cYnNcipH4XjOMHCyNUJFAIWHIzbBfu6Fyg5w18/pZ
hsdcnNUm5hbXckhMVHCalc+oavn7X6y+N4bfKe/U9ea6VwkmsCUolxSNV/AaJe0x
fRXr5ZC6g2jtrxsNmnKnuhst9H2CQtenGEGo3lPNiCwZYXLKSXrN4FvT1y+Yk7xu
eNW+1Pc8YnVewp84UlnxM4URAfpHMH/6e9yX3dK9FFHQkTc1e6BjDVw6Cmh6K725
3+cl7R5TCqRN34D/gY7I/pdl/VV/vuRKcfEGVQBiI6MuZ9M6huA8rFsb3Np+Nsnj
56CLkZgdmcA7cD27n+oEOeiRFpSmdjKCGcg7TsPr+atZgGp4pIUT9FwZFnE79x2I
nNt8yZgOuspnVa1eyDMdOpzwHuuH6PBkldvZ950HmA+XM8USsDh+yFhkf1JUemqN
App8i4pizvEVN6G7+nnEQIeM1/dE4QrPkJUB1gf8fvCCRuDkVBfW80cyA4ByCRV5
UjdG2H7rvlI+1cJUNW3yn7r10gjZRHv3qTAFAkMNohrogBdN64tm3/Sc7D60BQea
bOv1qNmjWZMYpULByWHW92CcQVuv1peHPil/s8MO0gCIYJ52EateUpG/O3qmb4WD
ByuWA5Uu/A0+onr8HMQruEOpv+bwHy6ii+n2HytLot5a1nOoNrIoXYbDAcClC5OE
C93PGIs7FWtfrV768jBWTB5JvVG/gvPrAkFqYa1GsRw+GCn3QmiRUcfYjWsKiw1z
4Z0zfs9iZ3KTzlRuMG/XnIrfov2D4V4hMvR5ns2APE7bg+G5qJo79duyIU/hwYbh
5WZuOI1PH68cSg3XqyFu9TyWFtThh2QtgpbAsqZBa1WStUCv5SXW50xG1mFBJtRw
Y2HU8ZpcLnaB3GhCDEd38+5cQyoBBV8Zk7is2tkdwVPLaFGUm+xp6pBRhPCShTre
AGqlHkQXN6q2TyriIpu+56bfCRQhb2e6CXElTPwG7ddT/bYyd8OUa6iT/AYcavub
v9HVKKgG3cnpkPkqkKKgxKHYHZm3VEo8Oug+TMjhA9uL/7a/h8810l4X1get3o2M
GQ93SlxcCXRT76aM7BE4biQeMEAyufHYkEeStFI7/uy0GX8XL0GzKvYTVZR/TUqm
RSzeycE2ZWdZjp4vUcWeF/vJWL0ILLMzxQc/A18uWUpxDTsygGm/sy3aIw18pQUg
D12cwcAKy/JWoMBFVxRVVwASR2I1ma4nATMAHfYtVIAfo1TuGD1m7yKgKGlBP4Yb
ctbNHz9p6H2Vwwlx9TgGmid+TxXEu8jCGL14v7EhCGhsPdctjIaxcgZ7+ES+Z+js
8fVF4h/Okg8oQ5WtUWSDR3IxjYXTfmcWRS3GpfYrnhMxyv4+ZBkVYdoB8udAPN1r
5LoCwQKrBa/zIvFi3mPuc9+ze3j/k8dwns8TVDIal8L8/nCxYIwGAbVPfpC59JkY
vA2AezpEccF7SQjthL2niY6mht/Nf62+gNl4Znf+njne6bBI0hrTlfRW7y15QBQB
Ov+ZACGgkMS+AN8PNINx639WBC4L6dAYRosLOHS/ZL8cLSsbMHpKlShsUbDnV65D
kOG7LrbX3qUr8TkdzS3lWIvTu+pX8N7WusKT6m7aXPqKeTFY5q9Dhsw+Z8I8yxkl
saaYaKNo794qhgSxFnGIEWDd2kjRnG9PanAWrdAZDZsMfxYXIqcy2Tt9EHOJhtk8
vvLk3fI5sj2+bV3I+ZLJ/t+cBw+PpnVAkIoJgwtXpM8cchVUlJFslcL8QTlu8sPa
cSHcjX68INT6fTYKXxp9h+HpST5/0heU4FwdEviKtKUDkfje+sB9PeiUUjkcM/PQ
ot+ybgdtZF3yxMr2pj6d+ZTaV2XykfIPe6xGBhNeWqoWCEdARi96TyoVustig9j7
TxIWACvJMHsZRahHLz4A7NNSD0bHCee6PfRdrMAimD9b/nyeThAtMyE7CvvS7gGu
PjrHi8Y8xPhzgwZcSX3bpdhy/daU1xitVOJ6YMpysUY6Td2RHAL7TU0P/YdHb3rR
huJdxroOj/X7akABmNVOnPuw5x5/AjZ+ySJJaOujpVWBJCUy4sOg2K7HB3RIc7dl
NFjm1WCSI8IA5iJ8EGHU+5Lb/ZYYTKIBrs0Euh3/0tdsCpkzXT9Pw+is3mMn43+o
pYnZv/TMNs8ElN72jUb+9PmvGUS7/tq6SEwgpXRfjBnpXI2CE8XzhDwxn3o23dbq
s8k2/FblmNZ+FF/PgqHb4YSvu+X2sp78ZIP5jz62zFnRbM1sRPS8YGDkX7rCGNvG
zKMbJaQRJgFdC2oJgVhmwSlwQdY5X0MsOh1WZaowIewI55gaVNYv/RhrOsaFbGVf
7a9SfpsJ00DXX3QVHl/+o5CHL4uY2MPZq7RnvuBFKAYznsA95Hzh0xpYyU8id7SA
3lg/l+DsD97oaYqXQ74LpmFS5aw4QSz6+0zJp+jNBnNopWBXc5mpo0HIKUKDwtnM
a+3eQyLlWrTy/JjXKJaSobJeLwFZ+wA8FE6SOCBXzY0kXtd1vKFLAhGB23lybZtO
ITslEs4BhtTQanpAiJgvW21qB41PV1HpFOyi2WZnUmXofGsBI+RYGLYnpXu6YfYM
LxBMFCxKtoZz8HsAIzqNMAn97Xcuwkzk/DaYB4UulFneis2QdNEfm0Xic1v//2TG
3TGrZncomW3BJAkqhLo16Zyg6d5aBv7XS0WjbEB19NTQppH6vMhfSQ4Mzj7MUlP0
P+d27MZO88nh3tQYaqkGobeJyQbbmWqhfwQYPci8wvPTzIssneSQ9ftx8fiiFi9u
uMiGozYRDoM0M6aV+WFF8P301n8BOmMeJQfmaM7FIzrGhvTmOtNkLVHlCjTd1HB1
16afjFTiOK8rUvAYG7SuuK7WKbsB912zNsiGSd+pqJ79z2KebOQgYoFiQdSWskaS
WnHiDOwUmlVFcyATtOt5vAdXEDXgn3eSrPXK5VdwaqDhXEhb0SYQ7rErPYPiApcK
m8Diu+5L7rHIQAlJFqMsnxU7aushRD0IQZQmSfqwYKD9Uz6cxeUa2BlRHy0hNk64
2b4v/x4346lCsJl5syAaHu9Huh87rd+KfaOylhFcxgFUdnbi2JKhGKDdC3gwdrEt
vyInzU5M6MeNVtihrxI+Vgw3plzRBuam5I2hW90JcqVFWXWJNYrVJA7Fm2lQNXX+
NeTLJP6zHHUh3AX52KqXPG9YdodehFTRGyg1r8A86zFF0HdNREeQy/InDhmfOngi
kieRZPI3OCXcW8lPEeqCZLp1BVfmRI2VHiskKQsWEhQ4Wacv8zyuSDUB9acZKi2x
ANBifBnTU/W32uHlaDKOP3f0K9GygJQeNCrRmhz5fm6l6pP1KYrDys1wZqfGMRxT
vmcLafsB8F/xamY6GUWXrM91vfmk9oueIR/HS5Ip3Y6JP1UbE+FfGbj+bCXEynkt
XYoBXyOqmzSqcWC6YczNm4RLGqFppzeY29QiqwJ7c6+jOzUhfQ0MC7sIae/Nm8WD
HI4GB9mP+Id5FZtbicSD/IhViQBbHXR5R7i60D+uB0QmTTolynJDhNTOHnC9MqVQ
TAPC2jf7iAcuyITqFxlFBDTMJ/B3Y17LGeGWCmtyn/0Bi7KOnYhOclwKuDKK4kks
tcc0iNKZbUqw0970UsesZJ8nWyHa2TmKlanXnsg8iA+lGH4N32dZX0Jpx1L4sd/C
M6zxbLIkOEZ6aaQuD+mebswUrwbs2qjWZxlEfmaavgS7hVVVrK4WxTDCeQQbjHAN
Vm6pLvCBEX/bEYAp4lOo1aH/xi6cd0JyhJK1imT4fHH7MwAkA2YySpHJ9EKc8PlC
ohHdPZjAjsgWLFRdZ6priw+/96tRx/5iFoHTwgUIhv40FPs2UK3dM56C22WDLOXK
JzHqIpAF7kdmRilWAeKGl6yTxiOyN/WpmkPkU7kq07gWu3O49nlXJ39/al66SWni
ko3LrhEkVQ6WeQdPRgUTmcmRc47yp6dGajhdIzPk9CRWDLyHTdkbCfTDQX9y4TKs
N7dVsL+fhWAe6BC/TtI/Pm40PCCoGe77IHpRFWD1K/Emu2Ecafj8oI+76QpFUL5t
dbyVMXSExXHcUORsNU1upda+hzt97ZQIEKIFwRhtl5GJtC1GMeLLcCSgKPUfU+sv
IV0kLzbuw/PF7lh+RyoWIQfM09yVEXb821WcXTcXYK1FLQ5zYjXX/bYkVs7siTy7
F+mnZMA1oHOIzvQLPOkNfNKypG50ysUixKLOalpfZ+BG3JdfvLjogwgJfuf3B/Ej
Bt5zcxLy741wrrZwYSiJEy62+f5XIKJLFFUoo8HVzdhmMjjG1ObKALGLf1iuAbfg
ASuSXJmkoCAS3yci9NXSQRTCwYmETI1KolOF6JZkogRwpX70zhHXapkc+BcP+5H+
x8dcKDvXelFt9pbBwQARoeRaYa8BEXxRoa0NIJ8eQeLkzO9fSpY2zRmpaToIcgzr
2s8bxj+1EMX+A+ftBbKLlNt/G5C5ViAghLJrYr45MsaGyfBuo3tadEg4zAlHFOww
SN6cyT5M9Jv7bH/mcu58INWxQcOsJJGrmtX1etsIFSY6q4fg6pTFGnpqcf02Kmo9
Ahk0jWwkqgQUUwXerU0nQPMAo98Qu2bUnCZ+0rTdJ53BLG5yGyc1Ybg+EOJ8bNSg
mBUhop0BLSSBXUsffl3gYZbV8VMObJs9Ibbc/XKioDvCo4PN+vJ3ZU+SCuk6AVht
VCV4/l4FRhDzhc4yiaARVZEEjbJFexiHPweZGdYemNJXyxjylAOsYNBetur72dq4
sLTnyXiFUIa8KxA/nIYYciU2LHTMMaf0/OZ+Kt99M9QLsoN4FeebiKraYUNjnpuj
6Q/an2TSVL+TTeZt0qy4SPfc6/ySmYUFjDLrcf9zYu9xymXX4oRhv38tx0WTfpuJ
fEAddSSbf7Vs6Ooikl3yHH/RYqKzlJdOxKMHm/0yi+mc31uFY0o+xWnwmOzpZ72q
V2m26tG6VHekgfLXiITbNRcCB6ygNvZuon/PSQK9Tn/gBGCRSSqLDZxevzVGj/y2
WU8upMsJtjlXVUitypsNgBl3BfJpqVFCb36ezCYkxNyym67H8AiK9g7izYDRwe0T
uhuaP+jmtOx/Yp4idzGX+JS87qxcWhOfLThUdmi9sTd5AMoSy5U15pGmRW7u4v+M
pMHjXulbnBqllV9QVjm5TaBIn51b0qNDRFcWWhMSPyXKOVSZsN+EC/jJ3y48DL6E
k3MIUxkAWK7mjWjzORF1mvNHrBp3yNWWRuHlzGGrfr0aaoJRpwsR/iAsku2K1KFR
SshKCmIHS2VwZe4a3wNIFnaohITPE74vV4HbjraJRQhHYAp4H4mYe4NZdi2CpYF2
bh4aRGIdNWxgzaqi0qZN4j7Tq9f5J9BILszu/oW917HmGjnCHTbJJbDm8rhek+zP
bCg0M5XQoqY7LRGWFEPBkuQtPK5zsl1O3x354mn+YXSueSkKO9l7ES3SMTeJexLI
KJAx7s62n0cXDuA9NHGBF83Kt2Cd2fp40LcGbaza0mkyVO060rdRUuy3Vk1Mx+zi
+NycTbG8Fw05/tb1r0+7FfIaZ136cBX18pEFaLiqSf/ojccjvCCOvJgNC9MU+AQA
+ZGobGSz2LJcJOLjJsileqC9bFgNEtLLizmPzadto9v8W6x2UR38vZihSkZ77MpJ
efdehAFCMsKOWz28rsqhjPp2+KYoJBZX1mlyTyNBWsAoHhjRUJTcotN5VYTcYN36
U0XvMZ4pvtEU07BcLMHuFmxUp8bteK8dSQ0SF6etqVW1uXwqTRAhlsYuZULOoj0p
hPf0f/HmGY0Y5eohN5hSXliQFwl3NcCvq6PcmfZa3qy16yeNGpdLcBPsW16ojZ2a
+Ld3aYxXrAGUJHf7i5GAv/86CmLEx/IAFLT8ICsmcMs06K1csRwCh2dizdeBByP2
pv7RcQ7kDrSsyZtdBD7S/mjx7+Xnaakl1bUAU87OYnxS8cHT+4MuZpPEc/88y0Kk
870l3nWdzEx1HGE6JQQowvtyFs3u6a/M5CXcu/MrYonuBMFXQH4hUwO8eHwB7XJK
mHfWXZtZXhR+fNGz95iINRqttUnbUO/FaPwPR3M22n3sOiwS/ZlOE/1zOhXlq1Gy
9w3mPMpSQWvGC7gTbg1cp33ecXijftOpU8yeOq3Me9lcDWha3Y3HVBNis7OgpJhz
Rk1qlQDc9TE1zvQvc/FWAhqnneINCb4+q9QTsXqUC3lK97armeOW1tPcSbhU/uF3
fJASEc/lGFTnhHoPVac64HPvwWV6Sy5tHfwCUhXzls/I1Nig3BI+811Uub0X1f4o
vK9X0vxsEHpE8EmZ+L8ZZgFdE8yg2q5pe92bZaoe8cyj7qhaz3BlQnNneKmNAY+z
HY3NlUbD4gTVlqciXjO/jx/B3XzXfk5fKj0D8AolW2aG9k1MlFTlVrFVk43Y6neb
VN9SMddT/vyO/2mCcWh8t1dCh9Ch3cGZmXDi1E3WokI7G0rbrMj8pJN0uL8gF0wC
BrGTkfSuw0P2GOGLwxjygLwl6QUlckaQS4JV/VgsIaBPjZS2NzJlfrwCK4kbiDLn
ypgjC3ndv16Mg6Bd5zMMnVqNZ8X4GfOeSnOo/NHJPN0GkaPyNdVCXo5QlAeRuWqa
rlJV8+552FGdP8zabBQHS7i7kTnZrr/3TpHD/VZsxSYTHS4k21mvO59sj7LRKdmE
fX4Zq/TpekmIhVWDBGEGfQ74zre7+/oTlf5yJF30dODUylrHLKlrijJ7a0isTD4Q
9LCKJiXAGA8y1sM6eqIKLymysUqhFPAIqfuVRgtaHbpBH/DAyDPQ2m4tElL44msb
5tZdGOCqGAc1AMEPvSMVlqGk8zZ/ZK7M1iwl9vsrVanEpARBn0b2cKaC4JweYRpL
E+F/qv/22+S21S5fTF1y4S6utC4eXIR2iyK0h3j94RgRySY168Sfag5NS2XyUJ8F
pdMeti4Z0JQbOie0nELtEzNt8kYnONKAzxoQVm6lcpJDAY0gnrD9HwWcw5pwI8lL
nW2YREW2L25Z6u1u60JFauLTrFJgr2s9NJH0nWfQuTo/z3nBkEpOFPxQXF7x+CnS
kI7+Qt4jq8MX2J2y17VFEJp8AWxrJnCp6BL+5cox30KUIgc6zqv1LNwCX1NxQVjl
VjJcbjTFAr1biYgqNZ8NxDIeDu6MT60DsiwYLeWZ/aQ2FqvTZFLcP7ZJpWs2tEJA
//EKgzBB/tspfQY8AXic+LeGbU1bLGtkjnSjBNhMXQPAOWp+j6LhrFecvbKjnUx9
3UUiTpTr46oOTXMdicqyBRtw8RDCegHygHigSAILPnqOz+j4asOJ1g5WEd3TCyy6
Hv8gb75aQFIUWIZDqkdM5xlFDDN1+RK8XHsiH3yYSPQoENmXfLJSd486Eunusd4a
0tT+wI/D0GpoA1M6M8b3ecviLnlxtcU9BKXy1K6GWDXC7sIOtoVRMMT+C6aFT1dt
jukPeXR3G2kWRYHwOPd5escPLIwnmmZKckNFujUfZnWgILFLNS7vWapr9Qc0/2cX
EaIqCBhV1KaBnluxlPWugyHH2Ryp9UuA+t0XNaRmwoR12qo+EOKxMc9vewLwenRL
5anUi88s/kPetCqQFatu7470QprOf8tR15jy1bPtUJdPrA5e88c2plUD0ahiuKMi
dwIVGdeuJTA9CaJYWPS2oz+tebXEMoEloaiOt7uOZg4hkEbcyZzXIv9/5cSDuXNB
NkJo4X/gUSER9AwruRMFJ99lSbhGA7LzOwOOoSmT1PXlp44alV0VratzVS1OufO7
m7LMR4/Aijbk1lJZIDvl+lpv4YkqzZZk0eg8wupJH5mFzpq1ws83v4elUqI/jgWx
fUrILevX9Vs8AFsPP4xeZty6NThTqC2zxfrF9sD56g+kt06uKyK16cuj3neaGzmL
POF5vbdQJvpDc62pFehs11fQOm68e4qkLyW66W58uLuswcpNJDZ3L7NU13/38hXU
h/3/s9sQEpIumS1b9lQvL9HLkDm3uQo5Llig8eO32d01FPjG+OSCpGXDtvRaKi+B
vjf9wVy721PZafDcL9ENJV6vqYFC0e2Wb4Z7EEVnLCuNc2QPGZ8NaQl0pG7lQyDA
bsVlTv/S4oQ2K2hTvQRN8ClLVIpesGXbvd2AVDU2VEsxRP+AqnIEoq6LQOAGvaYE
b5gqO37vphS/qDnOUXg7Dy2/J4igOoKVM2E6j9AShaDjrqk2V6aHtZRi1ebBllFs
m0YHjJWo1gLD0sHhXcBtL6oiWm1Kmk3SXwdDbfLRlAqkfZkzS+Sb57ZRCKEYcHoO
kM4grRNbZr/+M9Qus5m6+z7HZCphMKr9vxEEL+6AgXXJoTggeNB3QYmq5kRkVJ47
WDjVad4O7r4PQUwh6MjNa05CdXG7Kxj33UZqCAtKDdhECfb4hX5QB8DZYky4sMYq
D3WA6npd2vaABC3Eo0dU8mWcy+xolDQLZb12lBTzpNFSlbNnYCJB3+CrdCOTsRaP
3qF/RpiGvJcMDDUAvTC78Q7TQGa9qS3G0Y+UCrm6rgJQ6wYUyKtkzX4eOi+0wlwy
k9t5w7RcNj9n1dLDfeVtVcWDdsbG0We8777B6W1pbJqoPYvsiupQrIrM/s6YwZzs
wXxhXI6Dq8M4kd1rZLZ2iD9gaVPDzy09GShqXqGww8B0ls/jS3RpqKjIgFq21S8M
rsEgCbRJvz2OSJ28dzVGnaIjj/9AfLZNEuxh90s0n3J0xjq3qhRwNhgmc9Pnkmkc
5XNzFNZmPJ2orUbgK6GGnZtukEnIL9uho2X66shxAcYWvjTrxhR7asDddhwS4bdh
6atYqfDs9m9/i6Q5pDIle/QYkpjKhLmvTMKw2l7Vkhh9sO/gOVPw8s5TKql22AZj
8zDfulFX/yc2wBAffspfeM9PXKygaxk2Om9mXyU2K9edePYrdULb6zMgac29XD7L
wVhEc/CdbiSKxOEhhHWkj9T6aRJ1fb9Z3tD02kAuHNwHxbxEABuFR7CT5ca9QXac
0gU/0ZABqyvcKMk7eVZY6dAoZHPqko1yWBtne0muJAHumlPWsIIZjVNjvHQnat/x
camb0JYWoAkfArjKBqgEqbdncJj1eP/2zyMalPSOK9yTuPc/kDzxTB/OrFBmImY/
G84PX5AidFawe+YEmb4/7xZZr169Nw6g35OzKUcIiBDxqpMYdB8djecrSOPFpvQV
NcjvYs+8mH5H8/rgMYzoK5RSB3ARYR9/haBExjKlU1WxMRDUxEFSXH3S2iOAKayp
46XfGnk+OEC3qc8hr5cUecTwhg4I6c1Jub2U+rLsq8QF178dBPtSYPaUtwYOivbt
PrbT1xL8sYM8lfPVj41UGr5XQbLzF4zrK7+QHfWDKhw1yuUXWk/uP/c2Ug5TkDsl
UcduL9EI4wanARn4bc2B1zbNW2sevVlNMwhsUkwV27yocSIZU3fzmc+hmg/i4nJ0
NjyvDrOPg3q1PRdwfL8IzOyP+tczicUrxqidWjc7KvkqTv5HH2u7jnEeffZ1Rj3i
1jNoT3IambR9UrtdlbI5gGyB1qTTeC6ck9VVhN48yicSjw9b5y8LBA18tf7HNex0
j/JFaFml2W6RgAtn6+u8GW5WQpo44qd+ctFVHlFVJ/b07XLQEPTii8Mapqavjlsj
ZtRRspVs0jqXXF1HCoswKql6z5jMC06MYROia1QQ3wVuKuKw/qJnVTCwmY+0zPXD
Zpc6b8uhKXBa7RKqsgtPwLXCQtoAFfpG+GVUs1yueOA8uCvXDxkhVk8HKJK6kHDS
t1N0LXjfU9uTVU9aVFoIfiPbYga5KanOEdR23Mm+9TXa7oEZ370PP+Da9h1dllQg
QjVL7DhrCywQ3xas+gaEH0P+ejyK39YtlwH1FKtq51f8FVUeMHnhM9J9jco8FUgO
Kr7XRshENEEc5IPlA2ZgtCx8d2sDYUDIP9zultZ6X41eN1HPlxRQwEVE3+dVtIao
3dShDKbBdKZ6H6X38CZxCasy+aNtH4vlULVgcqoYwi5jD4tpgIiuknqqGujEgNVY
6E0GASG4Orgj84THqYX81ev7AVAece96SrppyMXNeQj2ns7FYeC6YlQmMnmS8e/3
uKOE//Ag4a2C6D2PRivmR2U55PEzEBK0TxGSCqMx+gKdfbAC4aSgz+O85HWY2skC
Z+Czk507JggZIEiRmzwbYRLyh1q6zSKAs/WVctbSLVl3rKcw8gIWZgg+nw8tAlTq
XzVm9T7lk4dllZNvSNKATLfq3sXKSdb3VJ2Mw6buNYLkLZ4q77+aDtYKScd6A09G
dbiFaBt3s92gLwn15VxsI0sG066Ze1t+UaQ/BdqOUcXdOzosecwLhCTWmqnOLm5Z
EYRxi+te+1sF3e+UDPIYSD8WpuxdJDT07KSizamKhfnlPl4bFm6hk92mcnH5tPVF
TJHrNgPJ3805rd4Kzz8aNMa8Vufev5n92ym3hR0sTEEmXNepycxwp8Z49Ak5zRGP
csFd0Pvnq+vItF8TVa1WNXbv2NUzgE6kW1rv1cKKg43tvlr8BKXVAobhN9n2+yTU
hb0QlUzOptC/Tse0QDTSuRKO2opoziPl4QnL+oFqGc5o30RpHC+UxwwUEWa3FZNB
yKnAv3kCNUBKfyVsJxtGSFf09W6S0g1ecdN6N82ZClZykeT5LVqDBWUUF6dryTOU
sfOfIywYoYuIqFBBp5yURIIwVYlipac4Mk8AL8zlsavm/hfKJ9TT0jfViXBqGIPp
AuNpk2UE05x8RFX4vJ+UhOuDgwwrTWL57zc9BFcJd5+EvHwhyCvv6/O5ziw3cGIw
s8P5RzUSRk5RAJ0ua96n743VGszyV3WYl8n6i6hgOvNuBWVsKH+pSJ6o6CnlmD8r
zOiIMBCZJISDzHHqxHeWrzKP/XDBco/p0gXgjFQU56ayWDBIL/DYcAIlb6KKhSTA
oTb83xpB7DbICT1CeeBIkWsRkdrgxfoKCjquv/FUnIUtSmTGbp6QkjjIjdTLIiYg
Znx8t1ACarVxQRgP5BL5uTyiCVlPJEmMvTRuOmjEi1KA7xHvaOj0j7HyviSTK9ZR
P7kuoQVBM6yZqe32f4yaLhLLT7HBhF4pgJvfnvFuglGGvgQnEbdYNvZ23vWRNCI5
Q49ULBeuXQ1G4Q6fQV4WVY8l9HNxTCfUGS4P8KFeK+615+Ot7ITrOmDY0rqT3Sfl
cMnCXghu/twr5BFmkUZ/ZzC/XEqsA+gk69kwDlaxd/s2DIcK/B6ufTs1YZR+ilCl
DDthHs5zcsZROA3nVBDaNRab5YzXNXI+hTVCYCxXjrzj+ej+prtobUM8yWpUaxjF
y6kV9zxFDyco5jsqvlbBrb7glw2zOQkXQxcNOz98MaWDctnSBlUajOZFqOpm+PQx
zEl+dSNbMnuBmQrqB/spAo5217Yk6fYdb4dWLe8Nb7eX3zRA6SfZUepqOw+1Icud
xhs7jmQ6mrTd+rfBOZdgI+Sx9eD3nQf0J5rkDn1mrJMaahtryMvKi9jSfiorUQ/X
0fcDIWDed/ee+/Qa77nzswP4cPlBMVNn82+I4HEsjFDN3P5m1j+AFI6B/C85R2qt
p7+nYhHCqK825mbeNELat6QmrN81DQO68FDN+6sl5EzFO5h4ARIqggdcCmE8lxg0
XToyD407jSj9vOWkQJbOTHzBOzyK6mEBD/edQXBVaMUkmtwYmz2b2W+q5SI8CGzO
B8GSZurB4MlELbFLNkbt7Q5/8u+7emk/W7RV1FVXGtbOnb2WuGeUx1AATBFc865g
nE3gXKZgXgHew7icLAr4URlOY1KQEAdNFUOCb0Zqmcc6ED83iSZgryH4cOceR68H
37hdKFMuqcszhkGl5xJGzdrFfvziMC7p322k7XCr4Ppojp1t3IBjdurxPcQ/EOEo
W98T3q6FHGPQuIoINkl7yWhl/HIKlIGr8rGV9fVpV3vIZV2jeNjbJLBd1METPUIk
9RcZztvSMdbOCaT9lJ1Fk6Bj0eQFxbp6dY+5lWEVqbSjSsyULrYCnlXD1BFhDosQ
NIHbJ1c3b30lavcl3zV+dVAh4AFlhXK+8wTVqim79fzrlTYeYICD8rE/zqavRL6n
RaukGvK/AR2voQ8mI7P7tqvsqpMmqE08lWmfdfCSxl9lecAjoddI1jOHSuEOXn/s
Xc2/L6NhS3BKWH0LYnvtSoL2GL8iCl0mLpZusdsSjIui8uKJ3u4kYMlOLBew1h1k
GG9hIKQ5ab/CEOOmjscd/N3mkWw9S0/j9YqtzplztWgI17i8fXiOTAsIfTTydTRw
xM5vKeNE1SVecxPk7y66zFCySKspqTiIp2yJvR64SqymCBwjXodO05Z+7/cJabVM
wQ3pEx2e+BByczTKN4wtzCPm1+HkD0R9v4d8gxU5FCBUy5vjOU/YxJEmSOs+10hP
4j5uKw0J1Mn0TxLaMM74aXyN/nahiBXK6mz782Y6jTI69rDqsa8miUJCDmBnIE8D
0VN36APeFcBz8l1rUSgw8GReK2n5zRU2FaRXAjziV3klUWAoZDjgFdUT2YrrDhcQ
0rl7s2nK8Z/wqI7GSGtsc/cIIhAxB0KU1mouSygVaV4zEvbJDn5N7VIeqlGksMQI
0dkvq/fVRaGjOQBOf8inODbzomQTUz7TCUpFrBxpk8dt0p9hu6YDDkFFINc02Hol
h4f0eI/fsBADpkLdmxLtPb6bwrxfc2MBWljWLQz7V7cj7orwaftTUKV7PltYSUmW
g4Y5s0sF6dzdtH33xkwH9iNgbpxD+IOMBRTZUxsyB3sCOktU44T1ijGGDujjARI1
anS9sfYDqHP9WVDmo2oBzL9LsEUA5ZYrRIjrquzv2dEvFeTzpgP/K5D6ZQHsO90p
pXbwVVkjL2DTmRrJGJwoFcjjQLhe1+iXm9qx+0j/u32v3ykPpNAmp0teTQnjAMIr
OJZRMf9QtyGCwbAHYRlWRybupCi8ojvkDaeHotFzNIbbQQYy7PKgX477NaDfLLzf
ujknoO9bfTJHWNYhU4LyE6z0JqJl5Y4eD3I7pT8O4LYWZrHdhYjLUKFMipX5+U4Q
UweY5l20es75gNp1mrDhe3qRfDXwpmN14lTxWHRVT6KUJKrgm5TOz7UN87JudjBs
M5aAzgEwOOrmf2yYBaVOV+2WMf1vw+ErZe7cqP/lrDHlyBylZuTubZrEjoOyttmT
q+tM4ZcVfeaoQloLZv61GDkP3OaiB1sTyTOVId2iutLXeotsguGXEjwa/ZkMSQzB
vXuV5IKeEDLUoJqmP86wVxSiXjwecBP4rbpuK5Sc3XAhRBt/3NKEghN770sSDSEC
Jd+G0BSt6qknlMsBoiIZnBFSeltA5OpmoBHwJ8HKh26vhGyMT2afIZtnWMa4MB13
cBlYnEMx3ql3wQmW6moaZrmhs3sWHsUdXicGs6mW+2Wr7QZO3Gbc/cvxSgT2JspJ
H3qBKcyWwmSIVuycZkHBY0zSwULnTf/w8ZVIxkLHE934Q8r12BkzS+KabKMOo07/
IgCNQeIoLOPkRz0G7lRIq2dP17BdxwsqDJNR9UEUVM7FadCQb8xIXO2xkncT51UL
O1zG/Y74AX5ANomUvvqcv/4ISTOPWyILDtAYW90ydNrvdfGY/nUUsv4ZvMw5jGqo
nX01j6cF/GUgYeaN5ptwGXYSgVRxDZ/XKpXOR3n2p77YNRR++owRwBrugXLwNHiZ
Nb48gmENFWVFQsxz6TMkNkRM+9F6MV5zr+ta7tQz4Id5mLZIA4PFxHEdbX/HrtsC
DyAkWhJXuWK+6aRzp2WY/XTkLEG6gYUKYuXUv3BEhsl+vIDEsDg8jyZ+2pfaDI+L
w0VN7u3+gPZHtbmIkTryQ4GyF33HQYDzCJAPC/pyfh53+ZxD7EUFTr0IkhR+yeJe
3xcv1Jkj+QySxvQrUReTUeyUzSRA8a0d/CCAsk72XNeeukSU6Mvc9M2A8O18BoRB
ONItIa+U7oXpDjZPpobALdq23877C72aCGlJikKEhqy+QhITLWLkeG4du0Gl16b+
bvw8DBO/GKPhNbHS58hE8gsn/2rRvj2gS6dgNeOA/zrYh3wppBz21CvyKYu9nO1O
2RQ7q6qT4QNf3/Z05e1kT9XSF+oJ5GZYSxuh575w4YYN1BjwZKeJN23k8Opqwbh8
FDqWRBfrcrPAuJuAcd7mtMBsdBAIZFKMI5HqF+c24RZ2Q/rnopQxs9ySG2328Xiz
V/ZHqgtmQeBImPUF59sq4xQlExJ044FkhcPusE6vR+vpmP3fKuKl1ebJmcao6PSi
hVM8Xjy1ajHp6bTo5957xXyBeexUUptcklP14gdtZVjVMQgfY0ThJJwABzpWjWV5
vcciTQWSiKNclJ1GPPt8Eh605R+FP1dYeLpxVmXcGOnOoGFDIMAPcaV9rZzXVtV9
Ya+1s4WRlgUPAnrs3l/6PPMRlIHx0oeBXGizJW/SLTQHIz4DKHuE2GkFRP9e2J6q
EUBLjUgpKgfKr03rt97XvNOF6FiGH8Q6Wn4GcG/06qLhzWRxLkZVGyfiUUwwGDPz
hx/OLaNMI06llYLejRRzem7d7rQd7ue7im8wXw2MmhJvl5dVSqSTHm50ANH7lisF
xuSsfa7uCGXWE4xalqTpPuZjA35QCsMwNJGZoheg+VbqUlpZnl6aXSVEV3iam+Nu
UpQlczTWdJWOAqzbmWdJCTV2Rpk7evgPx4W+Pgh2eZPpyHTeK5W3IScOYXSXZW42
ZtSeDGVD36LZg1d7tLFZ6NWs5sB4JcDEX4hzMlOX6kA8n9W1QMtFSf0/6IfSEg45
xzD5UQkiR3f+8A9FU4Nl6Ap5bxSQdqVIW4QJFqXBWiMNGLRL+WXKLAJvisnM2RMY
LDT+eCWnh9WklShnUAoPBh1G7OJQLeIIj0n4KRyjb2qhfU2ICyT81U0Air/VhJRT
G4tF+wm1yhz/giGZOduic7FCmHos57UAjGg3AWnq7UV2ZW+zhR7Pxqi1CsCLRSee
KofXklQbVKrd1knallPbTCxF+gaYYoVlVDAW6D7rQVdeflozHSV3bxROxp5v3NpR
P4dJ3tiMBwzpIdcHdEXPjy+EncBh5QMSh8+HtLnSGXxaHUP9c5Bd1rJ+WzkR217Y
k2f4PtfduJYTiAY5ytmu2Q5RCVO2j98sn25xm17IsYI3aJHpYplBiUv0RdOQGPYt
xEsuVsdNSk2n8IxKEwFRhaWr6+x2RH5pyHkkxJeP23sg6iT8C0kC2c2Xm9ft9Eyo
Z6F+w/0JJQ4nbH+qP+b5L1xmIQL0za8o0B9tSctWgf6JpLtsBhw3DPq+H6thqIeo
qwC3JDNifqi53tR3iwC38mhUX+urirZWgZAKq2rOV6oXD5+l2pr079If/oWWJPNq
6eB9/2q0wPdE0gHBQNBOEW1WGDvdP9NeynIAhjy+KfDWz6+XWg9bBDkF6T1cEmtc
CRGy50RuN9bylrtekdraxnrZszUyncY7HWdrN2GrQWXQg49ox9qKqKrcoIJCWJ0w
nllH5K1t1E4iLbTi8S/7rv8DrIcNfdgVQYTN4b7mm8jWEVB19g3Z9V+9UfKFED37
QHcGHy9Go1hphmjndq74GwOjuEA+MS+NHYnV8D9oKX4KKEplzwLxFVOfG2aS7Rg9
e2+CMG1Q6bb/j/Vvg76r8NQtuNG00G6Doxiv6Af6C/fXaPHRVrt/7O84nWmyGTy8
G43GUp6UroDhJaE+iInGmocA0iU8+wFSJh3m9i/7NTgOgT1xO/dqmA23zZOGKXF+
1/LzFwrNjr/0RUWzs6SxOVPuWVKl2oADwlRvHVM9OJRri+dlsA5eXSULLDXWQzpI
5p2v4bMFWw8lR+C01fnjE02EdtozFE/CNHQYakYMLu+YvNfSWOxDKFUS2MA3ibdq
7pqxhm9q88HwBBtOxxT4b0FfxQLangOaK7CrdVQvFNP/1ewFFtC18cNp1pft2hwe
RWYcwuY27bBMItD81RRZGx+MIb30mPex+zzv1gqDSDmPbtrJSWOOsX0b6wy4pudI
G8j7kAv4ayx9waVuSXpIdp6IsZqwXG03XkjyzP2LD+vpW31uRJqbfMZNO/vV6QDH
oDwnzgLG7NNhOtEnVtqj6MP78o+vMk79lBu2gfia7R8wxScW25ykW30JinDUEBB3
4/SBWIYkb0aCFr9LFHjAc492wTmVvVcWZbBgB54QnJh7twW+QAMEByRisZ2ejtuu
tlGF91rGI80mlpcIARhpIUastURLQcf5rkI1/7S1UZP6ddrp6BAemLHuA1gpyRnN
Jb3Y5hgURKtUH1ou/0JmGLdEfe4FqnuaR5Aaj+4/H3hdvKz4prHwt6rOG9gegJje
JUfFGXBUb8VrNYF2d5P3PLs/9BrCD6HQNagZt3ilQr30AmGzfi8lFarBFIlpuf+j
3cLBE+xvaScDqggEgiZRnNYMFjc2NSP9pB1kDAKupFgorS5Ch1JmcdChTIeYpwQj
Z1tePTkWNc5OQvHBtqqQBm5iUG+rKwOWGNYx8VUah86ABQhm4uRlq8MUvQXJ794F
YGwMMmlrin8RkUz0OXXaElULUafwJJqDT3ivP872N0ZPOX0I3HKsiwYmnPi8CfoG
4MZDzzKoVKvnmUtReYa630/H1mXrbGd1LdTWlwxazMm+lb5eGoMTkulzBnyzosmT
UcBxMCU3cGPw4xxbi2adBspoyIvbmegTKeXEc6T0jtxPufqkW6PSbSfWrtpa3yRf
Uu6pLzzwS8g5VHkfHdUIgPF54TJVTa7HS0EiOiLXUncWhoVK2YL+10DCLtB0AcSv
Ds+EDfAl/xFEkdIywu8KGUU5rT/0qFPLaSB0ih9B+fnH/sIZPlbb6OVKDGF13KwH
LZs0BdwRSjaR8lJq5msENrUCtJm1FRpXq411uSh019sHrIX9eiG20/pm0Ns+BbgS
+1y5YLg/jnK4Pp85JyslEJ2iILqbEvu1DqvPnlIbjsjUcAqpy/WptjgqLPhtis//
1YNaoec21dYqcnBvywjE/rOvwin+YoEXQzr0WUNJ7dxedJdt5ncMMXLp/+ZlZWEi
LDCoPQErzhRUsxERoqexeASPYf5SlW8suR3OTs2NrWjJVHqmbcutaUmXRYy96rOr
5TOiF3FL4ol5hlk27+8DXXGacM5+duc69ai+4kv+2DnujMsU22KvcFF+ekmAvPzO
ssDBg+yXxPTZXw7WQSfcwzzn2Cp9V6EwXASOqUrViYkiy4JoE0tZnHkcdhQYgKY+
EdJwOqI0JAE4/ZKQT8sZ+DeifGDGbgh7dZBt/6FZdcPTZ/9lJFTIP3shGF68hpfK
MWso/rpJudwvFZtmwmVFUInsHDYG+swXto1Cg/hzLbLqWFGeYsJn52mOO42Z4ZIB
O3OaKSQ749q5Toybq834G7r9uFydShlE8TLFJSjNLNjS4An6w270lGUgqbzqVwcz
j5YTj0TTGW7T72PxTXKTRTWckJPjee9sAZ2YBKmxNhRIN/3upLkh62sLkymgL0l8
5kMepIpIXctnaw+nVaPb3JWiRIht1dF5JTbJYyZ+LpevNyT7w8qFVg4w/s4odV+b
kz0smSAWAIZgNWI2Pw95AbkqIr60I08Q4+HxUgrI5h7YMvfjijbD3CSxmCaGvIdm
W5p0xPJs8Zo2tRnHZVv16CCvacxjYCflXy5FsWrRGegkdgD3fxwDgttM/tR0SDtr
Eds1dq555F18CQIr59H9tn+DwtK1iCc/7v3laOGVY5rkXGmEqBkv6oo2y5KB4uiI
Sg9Sbjknaw0wz0plGq2K9/ol0sGF/g9uSaIEV5FhJMe6GgK+ADx0jysyQEnC9HSM
fN+k0RD09yiko7tlTllSNsit8iKmLu1oD7SXakJikdazg1wrH3vbi7GBHOL+YRoa
6x4uDlxTcgVP4VG9Iyiz0o5dhKb0vs5m8ZI95xCPh1HYeHP0D65Dy6avLCRRfGMj
4wbl4+UaFnVsOosWqnRFwdSyZOsT985ZYWUeDV6mY0x61g4mu4nnry9/W5CxgYdG
m3/fw9cv45I9Ot1R6UOaStrILRL+ZZ0xswJ47/blW7YYNX02fCrP7pAprDSMYMPe
BfmZFZ9KPs2g/BI7jr/I5rFBUsrPcH8B+6C4LCl82RgQLrR5KI75VaF7CnGikes5
lfnyr7mUsSPlqrnzBg86hvw3dQru86705YCjZojb1eYpvHb+RLRRNVGYVZw++qcn
GCF2VzPORWoNF94O75VcfZLvKXM6QoE1rfUtWgW1zcEVf8uaBDMVsx6/GWxKlA31
9p0gDkjTlEKVX2UKemOLld2Yje4c4hxvRX5bzHOPS8mn9OuRkCwmybeJE5tapFGh
My5B2EKzX93QgMspdaFoLzWJiOktvoEu4KoIy/0hOsj++LlPaSqe5/+rm0o2OAOb
BKblp3GMfgbgOIsnUlR1GWub3GStX4ZVUArRR6QJ80weD80DiepxmFf0t0Oxn5FI
sHgJViz8gUcOkdcIHxbLOXokTSYz4F8VyzFuZfcxv8e3KhU9hePFHgwp/B31n9Li
T1FIXda73DRtC7RbpeucVkK0KhE5/SctpyKgQQa9Z54PPY8RoGOW2YubHmm1suNo
/aSzqqvqdy6XkUnhEulWF81cnYxrv/RRDel0XM/b0G8+AOUX/uN73a1ZVtGjPhIs
+M0E8lXJ7WRYR4u+gQnIFhCtCp0kD9YtvJhptLp4naMmcmz/HpiJPYviKsQzXvtS
wY0USaIivLg/NDT9HlMXUII5KdGgt5Xnk9/vM8OGRJ/IMNsQXIMXGZtlGsFNYWGY
GPBKhsK3llxbUPGuw8U/BwdpakK3DVGPW2naVvIIqJrPzk+noJ8+IxUnreKeBZqR
zhioQuMBANyvkkrzoKMpEIhCjFMoe1xPD0vQyRyLjcX5lychB+YRh8SAMQDARlYW
kKAgHas9KQThxAw+mZ2H/vM0CqmJ0b9WPBaSWBuZ2Vc7arb10UQBNPm1CD4Xaps3
pGrXs9ZUBX1YadwVPjtSt1B6CoUHRlFktcsEfd2XU1RPG40+bntDUyiiXuiB6F/a
qxFTTmxoCJrH8vu23PFtY4izF1zmj9LMQCbiMFRo1Wdai6MnfTPKdTgirlWgHJL4
9PRtb5WPxRxlrz590GgK5XYK9+NYb/Xa4h84oVuALVLk6zPOOqd/HMGLCTGNs8WB
4ym9nkJDCYx00BCiwVCfBM/nHKFkFEOsREKFI4643T/tQDlV93iNM14qTOQNtGCV
AsSHn+Eweg8MkFZTo40d+R4PNwnbSbi3BlCgtoLEA5CWPJbPlS2QXbk3YAeDQQgl
zTF323yN+iV9L8X4UW9qF4yJzWd+95VZF7u7Lu7fyHvqmFrJIG8F355qQ2EghBxx
81l/myoOxlHryWqkTfgq7VTMTqZu1EvfHE9vIIMJ4IAk1YnGd+bxOUNkgAF1DNfw
uxdvX6wKorB56j+momuU5fbuu2ekDRny/AKjYeczU3Sde0hq+zoWatrXG6fYOpeD
UDfgN0UqRKbbn6JxjiSNsg8r2rQhwbxDR2VeooZus88oXYRtdbzKQ7WOKCty1pks
Cv8L7LtlhBNTl2ypvziwBKoP3PDBR8vn3nIYoBu9sgNV8JMGL5/G1WY5E0eDyK37
t56kYZ7y3+8+dlfhf2dMY5jHPL6hyaBM8mBwo5evszoqnhlXU8g1uayCG3RRNK0b
JQYYbkJnN/CdHdXbnPZq2EoATATEP/Ahs4kP0zL8ZLtntuYrIaSk72w4UizNz4GA
WZ50RQ5JTaxAF7YGPcSDeHgRMuQQvVVPOoURNu0y+AYe6ww5rh2SRnCEBbBIhupk
MH7AqkETCSLHwBajlLLfrqpTEJMC8mf7pN/l9NzQlPBXk7Xcpc5KamINxd0Pzaqt
SK+llC6K1MjcYatdV8cE3HQkyiMow1AvEL6XrhmSnmhkmi3B9r0iDXuk+Mdm4Jm9
nI39G3EB9j9p/KF8MSizcd8jjkn3kCZibqoQmiYW2+S+0E7w4H7SlCTV2oFh/40b
wzxnNluvXuNulvv/9mlKfSjmM/aYQl2ZcgM+r4DCccORdAx2bwUwrm5C9oWzt/Fm
UJNg54R6XqSYMdsIwVZShLgG6YdLGehjbYLtLtt6e4xE8X0nAd7C+UYnrHvMrs25
VOoLWqZhL8Oz40lhg9NQlZYwM88cQEZRKQh/02e/63Co+AEXEq/JHl42H/m4MmPG
XUkk6D4OhzwcrRGK1jnZzZdCmPu2+LtOXN6y93BNY9abVt0ZrwwKBmQ4qtAw/tBi
LdJWhc2FdQru7ITa05SzgCsOUaJrH861SfJ1n6UG0+inRMI326F+ECs425lPsRxS
LRh0zXTiM86JIbOSZ0n+8CnYMPNBojHlruU1fQ34HadaZG1mRs4WS0wx92Jx2zZv
kqXdUVzAbznpc++dt+5fagn+Ez8VoPgCgrniYRs84JZFxeQfovO40uY3kbMWWY9t
AOY0ZDYjLLGLnF9QFI9O83RyJCLbBdeKtIPnDb7ROHqn0iJ7h6/WYs8H1RZoyToO
vM5usB9653c60AZENFsA5Hdv8XB3haFwQImBBufBW4seysO2lGEM/iK+3Oa+UIF9
SnUXCA2N5AULtVoHqwEvb3JhPAlKO/Ilv+r4MYWr9Qa3XpQtNbaD0q5wx9SH3Syw
Eyi6zUQci8yCD5G0vOVwNiF40Ra7zo+GDCpuBM4xZ0bKWQB52yw0aump7nAXC+KW
LSVOEvY+WqL4UgXe2oh4ZpmvD/ONBIEjBEEPMYRArFpuDLFJn6GGOHg0mynkNW2Q
UFxBFj24bk5vKJxj8w9VcC8eukg50I7CmlEtqbqCIbxp8JpFb/llMgVkqnb1FgZq
mWzXDGMafOsgtYBrgHnaIF3OlQK9FmnO5NYUpbURay5deMaC4vUqV/8lTO1yMSf/
TjuS9sQF+fdfCa6jfrp+UEAHtt5HhGEFXqmNCNMf4M6yWbS+g4GfiMa3OMinQDIB
VshjjwscXkc/3P/jrkvKFEdXEW3YJ/SMWDm/jCVAEn49zrJzPE1fF5vuBcuq8ngS
SxBMbUuS9Bmn+UH5RNvKYY2Nrslm8uWtGAUVtspmt2K8xVc4fV4cFn1dgdh6mCy7
W07DqhqCBhr7KRT2pt93o72EHeZPGD07JCJBzoT+A8gn2JmeCwbM0zcEbVcMDzJj
TQRlsKInZcTBa21aXdczAaLZB4BN7697vVRg7F1QFfmqBndWN6sEuU6V1wNg4Y7t
FwIbQbvnmwjHgXjqGxHU9L753L/5vqWPTHiPEycg0eMeuJKn6s8OcYAtwTTeVKeU
xuZ43ED0XKnxCBhd7HQ7FfQDTEC/M0W0sFRNNhcYxIMabP37mm9tYWTDlX/47+18
CcElhbpidvgn0qf5dtIFkoWGS2Ph2As/Xhi5WH7VJXBhNq/fCOWCoKJW/vHKB6Tf
NFpKPUd5GQDS0RwrDaCMBWL/0ZyZjFimkHDb5R+h3qiTLp9dDLrP9stx/tyXS02y
zxBUGEgjWlulv6hqsIHKFjLLev5OnfSelL4vomsReKdv+F3kEkBOshqzumkvS+ZE
JrsAWPMQDtPMwjTwUwtDn4d/Pa7qEFURNWugonWcbMxt47afa3RnTzChIdL6kmP4
eL3g+AphaZpYgvmyD4rrVVfs3tQmBQrkkENGi9sqxByN4kC+qS6izmrq+LG4x1xV
sW6dD5wm9GVIkXBhv+65cmacCmXi6I8J4H9tilq1oUckhKf66tiFAboo80g+IAp4
RG3cjoXF9EI/mlyu01lx9gouVdQHqjhXcn7hDP6fvGrWYulynFYnGbHUhEY87iwu
2rCGnLG7avhVBGfoOLTIw4vuKkiqpC97A5FaoyNdWL+hKwn28r9zYOasuScPHwFc
LZIDx6lPKYZn48Uiy+mDEq2G1Yfxe+d+GVFWyrkIWej1OD62rTlXtDftLO1XgP3I
AmD7uVxayZ3Ds+eW/sdUyRotiaU4MRs4vLMbq41oSL7UAAI5Lxc68tiQTH1CXe3I
Mr3gsWUo7PLrCKHw99pAioI0nUqffntCeMeG2d950Ug40Q9IvM4EjGqUyeiMbFiB
HtAq6e52zRlDoEVLO2vaoMdSreoMi15miN81rzGcNROXlDbWHBnNY8MYhMGk8ees
MbNxIQtcgMvYCvxFN9/ioI1UQ9Jj8UaLlEuRobSF2ipkYlEufKJ/JqmquZ/EuHpR
esndGyFl2DFbRQS5zBgVH2Iz388cdCNAXlMAhhE9uwvvoWxIKhGNn95dUEFjAt86
oQQp7+oPDjKqoisBTVFPSwuTFNZa4Z+MCZMdY3KtPCfjc+MFO580/U1fanyjA/sR
lNqGDSogf3vm1unmtPVhaY9IiJ5hL5nZz1Cn7RRlKahdvPKLlO9C6iUs/Vh/TyW/
dE9JxlBw/mzucvk113Z5AIZOoChL73jAftK+qrkuz89JC7IB1dMXliP1xKhcT2GQ
BvyCcqBJ6YlrtArTb2YVWQFr2b2Ayd/E09GfI4lgDpBOZ9cw841L5Fbxs6BPhj4X
pHOcpwtt1ElHI4rGtwpKMrLJ5hckTmhADqcv3yE9MoNaDV/GSrGU45B2MWNA2DWG
B4e+adpZnUOtOD72oHzs0CmVlCpqGKg90eJEoNxxr3+WPWS2oNFTSLTxZIMqqKsE
Mz1HXav7vKXYBfUeCdDkqF3he8QQx+2y3RsXAw+G+dbSq0GG6JsmPLxWZx4nDtfz
U8U70DuJT/p/YkSdyVPr9ECj9aSuBrBgZbyHtugizb7DWzQn+f0fo2vWDwxy7/Hv
Qcr4/tpp9bGWKUX8jwG88oVnIkXEXeq5YZL1pnOuaOViEQTHZ/+trB043jg4d1KY
gzqjVpG3xhjhOU9MnYw9nTv0m8qoyLK0qzGWJYFTULCelpYa7P4j+TigBeFGw6AP
cCUHc1sWbdaRM+XNJ/wQGv58pFzxWl7Hpmvb7Gt6rhccXX9kfhNAbyYRU1D/11Ca
mdiFRSWDWNKyiO59wqT2He3t4wzvZHmNH71liTDASsCA9B/yNiEVyKxGuNhnqzSB
24OQLAgvuHHYguLhpJ8IxlDJtqKdPLZi+4I2S7I7b1JyCeyGqMAQGbcdQ6PvjK7q
ZtaZco8R67AfCa1Gy9WizO28upKV8WTUAkVfxhXmNfoLqMOuPOw8kIzLmLmlLDvv
Fxc88m4EmHSIz37Lbczk4VvEm1ZHxOrpsN5r6H4LRNlpt4nEVt87zudKhVwwhqZ/
WMRyYpMhN3BoneGx6QyiqyEub+yuoNAiMQhrZbY4usv9Y0tG9flDqjDHiFP/G7pX
9zxneb8DFKw8iGRCeO+D+Erb6siYiQtqGx4gB2seGKrdKu3hWEr8ftV+14QOdp9f
4bD6sBftOG3UvvkT9hshdLWLyUVBHCI0e/3u0duIL/DXplWOj/OHb1YT4UUWZPxs
dZ879XT2tXju8SaFIdlS9JRrSZ0ii9C8B2WlAiIt0jMLtwNULk1H5yOH884wD2cX
b2OnBUB609hH8A06yluEdCPlr0HZWGHbR8RPFkTEpTlHORQ7dGWgBWLOSip16p/d
9evNe6IK2aguV0G6NNLWyFImCurojYuuBYKo1N/qR2TGO0bEXnF6MUQIJMAmlZ94
DPmE4ywCum9wWIzaUAesm17TqtdwCDTMYFWjP4jSMcNmdBVqU65w4knF7JWBiSgY
6iEgwKFvhGUe+IYBTHxyWA0dkKIxPdNmqR/TftApCP7EyKragIyF50JfDVWzVb+i
ka2iIuLodOrlrB/T9UIzbnnaQ2/3Loe2/nbdLQ7RZvMhy77jO3N+bC5U7cXHrMo0
t7AIoX9qOFtOszEtyztXIFSy9zKb8nHQvZqph9vYVihAW0rY3+WjvC75uua/EaiE
2DT6tAgHykGclvrBgi9pzgHkkTyCM6JHrmvyuuS/yx9ZW0Kngimca7BfkTRhWPGm
VDn1C8tcE80JpNZkUZxIBLsqp7N5cP769C0Gw3POiqsgrQPAUtNEvU75wcPa4Xi8
iND7Cj2GGPbXABOzgri2yJbiO/iSKI9hnsdiQREErtQALc8xClqYttfQzQ4jc1/S
0ckdA4vSZpkyZsTIir/HiBFuiPghWD4aokjGh5XSGV11651Ig12SvM7KabWUBYkq
QiLOtRtts2FfQ3+RZCSppmRSx8Za1f0zmGgDNxeoj2RN4LNUYj7NX3BhMEZTq7IR
0nI6gwWXFodcuIIvEJNjqo1i7JzyMmhpi/RrjzrUtpwLYSkqRBLrc1yMbij0JzoO
h21VcEkK22Dc7iL/RyPAerj5LjPPkDylwAu7hW50aRwxKnn+/GpxwKxwWSHz6Vdd
0bKhP6cs3035h+D7dpBF3D6eJFkNb4CJzlOfQktxF1EgDNb/7XZSQmnuU1aMwc3i
dMvoPtwD+MMsO3Ua4fGdBIitU8RYiVxCXhX/ZoyMKFd2wCogPzj0pJ4esBZOj4bB
CJA3x1Ed8ezBF1kNaK+DZgKG5+QteW4BfWYzTkUdA1uduTbQDmOaSs9LAg9dnoNq
BtFNbGVM0bnGmMErKGGl+ZC9opAVs30KVqS0UQ0octzZKSCbBz+5eEnnkzCxuj3w
l3KOgGtyQRNt0N65bWq6xFC8cfvz/Y8HLcs7SIXrLtm76b5UnUl2EP1JVpvD/H2K
pURQCYmmm95wfnyBak0bfTYDmsixBPoC4r6dzOkD4zZQpDeJI1etPi6k7wEW7D8c
B0GELSMZEHuq2QEgfIJlTKHZqV0jnV6PgOJIutIdOndvom5/KkFOP298u6zZyXfV
q3iubjJfVtM/8ClfjV+crhSYE4ifJN1WmyS5/2VLMr4kZzhZkL0XzgJAA61z2N7r
3BANgvD/oMj6LQJ2FyZHeQMgXU0Y844ESZ97/kZW+ESf90xJK34LoXWRGa6T73rK
iitZBSJyqKGZTKsxr5wON83wX0PV6Jiv5eKg4a434rRUCenNAhhG/0m7LgHJuwyF
HrfPHEOOrTH5Vb7j1CmgEVFsSTHbfMuEbT16W3yItop1fgDRTASLWTYGXTLPDJUp
r2J4Rfe0nLLMERimuZ1DHmRyCw0EMsLeIeSXEeEFjeJfcsFVeOdopmXDZY1WYvS7
jy9d0UuH44O6hOSQrSi6RmorFWki+WHKK8Ugb9+6ihBeGS37z11+eBbae++xhsj3
gCeaKEKoc1fPaCrtaTwD1IEMmpvjebxOdpM3mkaA+zXYIn/DAl8jMb9OcKw1MMU7
BhHQ/1ODdMk+hjmrhWCOdotUmwvg3ICEnxinAlZ/rXwzDtslyVzX6ML8fFEJuAIn
giLEn6b0ajwn/+sKD6czVNv7Xmp6kFLxFySxHmsiZ6ayu070WEuMfIu2Q1JFaXwv
orxB96CPdZ3exzUDn1cw3W18/uafsgsTw3KHk/VMjwHcgStTMAWO6W0U1UkDnuE7
g5qIWLRXvFqJMC+QmXophYvjcsX6j5TFpgRA6tNRiphdYvQ50NGFJan8hgHmzBk9
9JsUFnkpeZOjC1SvluHxs/J9V6kyXEwSBHiPXf/vHAltEMxHB33G7HtGN8MGmrBs
NK24BchjGJhI2O+6waAkFDbdS3IUI8wZvtQANoun4FmdZ5eMXjFay9JYO3p8S0Xj
4Wm3p7q76rQvzYEprCRf9VX190mOHzKfeEzFmLaResWRFEGG6HBNh6j0RMv3wPQF
WgA/pEC6TOYwD+ak7rD5Ls95GA3xfFfELj5nUhjVQcuquy2VBig47AkXxImVUNtA
5T4hMenm7liU5adncbv3hlOxhSuokTVNH5yKDX1qsTNj1suMLIbVwiyzvwqkEs+H
nUvop1X9Avq6Hzl3F8eKl2X9ck/kZZu+2zACbVUMt+1/XtHWLyeWAXNcKgGC6PYY
4qGZSwc0RN6Nsnk1JaoUFEDEL7cf4G0pdIdY55QpnW0E7wkVC2jx3CZs98gXEdnt
MYddrpI3qAmqIsRm/3KppNJI+k+YBlfz5UQdoN5q4Yn116BD2VPuuw+R39cGQXeY
BFmrny5G7OfUbROnUWvm9FUE4NJRRZOUAFGRSK47VJOr/4n2RA0+RWWIToZ1mkz8
cJszfiuu0Oo6pqmjHAJYF+kFn0fr8/lRy8f0KK2VNRtjc2lhlH5wpT2jZwXIDaa9
bCpMSVI01N/LWlKePOn9/DkOV9+ODfZMZhxouPhTa/wspInJD2A3I21bOHS4mur9
LvQ1nvZ7F66IcazI3g+C/OdsQD45n3nVFaxeGVcw9xKLKQC006atBrH6EqfwK7zl
3pwXmc9N3j2N3iC3Lkgphr88dP3a21zKGRjQ6CiXXK5k6eT50SOjHzFWrLZApHIi
oeQTLguCHG7cEIG+tsKNcaaZE/t8mOZOPSMEhi0PlFt5046Clgnp3+uWdTGnxkKP
5Uv19tbZvD+mhXnDufBbhKQ6KyVxF7Huxiut69L4unSOufW7laiCBz59mG2OtlCH
Y08OxgOM1Baq2zA/s5w61Lnufo42pPOoy8eZbJ/J5SNCVNXuDmc4Qyo4ftf43bhL
RbP2+faymeo9A4tE9VCYhTsfCgWdNQqgnjHOFnRwGyRxzlpg38sXR4e+qElV1OhQ
QkUiaxrAx84lFyB0ZGoaR3142yL3h+n0RDQDUOiP0FwAGMYK8xZxfnFTc8Sxrh4n
hLRbCnMtFjgG13MgjBhzF+RXNgVzY99Czh0UL/S2hwtb6uNb1cfNWFA+BPCNhI7z
QMZ9fCAUkziDNhcrAzjiwKsUCk5b6/4OwzPlFRDK6dnLnek+EoKJhPRH9diuDQc7
eLHeaPgb5Sz7IWUSIxlk22hTNxkMn1CBcLiThGV7kYsH9mvgU+CjnH69+brxTqK6
go27X/DDp9xTlk/Sx0ft3m6EF5AYNvttcE7gm/Lyxp4dgiMN31FFhQc4o0foRjng
QM3Ir3dF/wljFUrgUgHckCDnjzPNc98bGcijwjljTzmC4rgbc9KFv80sdXPd2NBs
9LJES9IzYoeiSwEQ0FW1AyrRNoLxQkwQOEhtknyfwLzF45U19moEYWXTKnXCO/F7
A6WRYuRGMHbDHe5d7G+3KgMUiepANV5Fw+ugvttAtMxIlEWsWe5GA3PwW4vP7UIO
ekVs11uQV/mDfxwwu75J7B7HO1XlCZKLYZRJKx8CyHXyNBZlSH9wrYxlSos53BMC
x0wZZlbEcV9950bZdsmYK4IpcN88mWYWx79rvLXSoNnpf86zZ3PdpzTtTa+27R/C
1ZjCyc2aqVIBgrp9Su2LXb+IgJy6KdYdkoUJVh9453AE9+3714XmHxjX6nVgvVbL
8EumwI0UvufQCc77rejJ2MdmvzO2qDiMwink5pf3UUx2LlNb7oxvi1DwXpK9eTxn
u7K2hQHzE7ePRyV4G4b24deToM0HeHneflCzOGpHQgXcyFMQdxgZZS20KVxfZPtP
83EmokLpu/dTO+ceJCe/I/eJMP86lElL/BN6r11zva0GG8gV5PnP43nwp8fvUmmt
SN+9QLsEpLsoTZ+p7Z8gdzrklv5GgvnYuAKJUm/3ZJ4zIVWX6Er5T7NpmPyxd7Gh
+1O2Hj9wzWRfwW8JfLrKnJYVy1N1E6XHOCrBTCp4m0VHjfnYY8gEoNjpxV3oKNBh
4J94fGzWIGeH2zJd0QvMp/s2Cj6T/GYdHOQ1IXOfTdH94heGRZO3B0wd50g2OP4q
srsZaBp12TrhteGMq7Efs3MlOlF9Wb4lDSb0QOXLUq6fX7moYo7oQAHco5zZIcuL
5sReFQyZlP8Z1N3kdG+R2vZ5xNfrOhEkno/WSXdXG0aEvcQV0MZ4+Faog/98eVvL
+WhnbdSxpjj5b4tyr9WFLmE2f3/eB5EKLf/gmK01apE6Ds9Ykbj+873LPSwevVNN
IgLtopbEWr3jb+F9AJ721A+OCzbMJpJTZH+5K4z1UcgfDphGQoZetsblEUPC1fNY
yK5zyM88c4WIclSPqx9k/9lvMKZeaT8fMnK1kNWdbL+s4x4JTem2BSY5p+Sx8SMU
qPsSezT/fHTXVK/KnDZP+Wq0MY4FdoIRaa0PgAuc4dQqNuN9vYkA9nUq9eYT7yVK
h1AF5jpgVArdJ3PA7lZyZwg+7a6o6Sj2H2/wb9YvdOH2Nn89eSXf+oGBLGv8CDvx
9vbKzTbQa227B/98fB6+P4swCAL5R73cHRodlZq55U0ftPBDGiD3nNihxQNt/UKr
t9HvBOzMY2XpYYsZdUIdP7UWLBUnBdqkGVdVAnAvHlz9hMCEEygVFwA+iV/SLjL2
Dvb6e6+ejF40SP9hC+U+G8YuGtDMgp2Lk8IdleRTzN2UtqNAMNXN6qVn29g1lagg
dI+iyCqWnMfvl/5PSCrh1Ofu6s6Nm/TeA4r4ZHxKcLRFDd7QmW3L6mvc6b8G3lDB
lDcVJnVkhlFVJO0+Z/5qL4um15zxPyULCwOd3iDib71zZ0qHLzChR872FdeyNKOf
TnJHuNBShjpKI5VkZCQgzwX58gNHKMr14/KdECD/WBBR3WDwKgMwbX1zskCIlLeS
fKZdCL71oNO+tWnJor5zBT1bzTmRV0FES3+S82HbQqzcRWSy2WraGqdMTO3+14om
0/kBAsT4Ng5TO/WObEqPJi0P63clUJfq7mbN88MsfXSyEWcWVRIGBEVuwThg+mML
edFus957NV0yfmZX9hwqzriqbx+8AoP5SGDxF/AXw/AxAQJ5jWANyVqPCeEHZmxc
RvUpYDeLsH4eRmbq+HgVeHFi1oPhlNdKp198Nve+2ZDe54MkM9SnVxSMkf1A/Zhb
iJjETO/mtMU648EusPnGcnO7sI/ML2Umu/rB41dX2DAXjSR7DlJakZQIOtG55Z1B
Lw0+VP05aO35KjoghxZlC2QfWeIjYD3VMg7MDGstabeLu7fzvArN3anm0YRNxjTx
CBH/6XHt9lDMvdFN/P4ortdHHPN3NY1nWam0eUJF6msga71CKw+/8Oa/jNWwYO7l
w9KheWyn+RQzeEJdR6+wP0U4gsxOgt8efXnKnfrwW+N4ir1mzLykj3xcIjLMZFlD
zCHAsgPHaJhnG7eDzdQE0wEPUJbNMc0mW3Q020Btqj4wiy0HpgPK9JyjlR4sLYiA
LFpg/YLUcJhbvT73asonZveuyemyMU51FAAfQ0PhlQBGGM+BkLCa23LCmuDLeQbC
vLu2ZzVglBdzNVVyzIkpoCqbtWetAMzHlvIUzWSfYJo2TcpSVcHCS+2hm9WiWbkY
XVUiyG+ZZ+UIKfm3+jkZ+kGI6BRoS6HfcqZ8aYPtvJP9fjHOXBHDN0Zcx63ReCf5
8YbeauzhQO9fC032EuOoP6Hb1WdHARnSo3eV4sJ27bu3Wmoh6QcAb58ugMCgjYun
pUfHRMmuU3L2zgDk8eg5wtQL8tfWj9JvO9LRfR5B0OpeiGzRVZt1YtPY7rkv8mas
JkvdvQHBNck5i0ANrj1EkY1plQtohHT14A7/sz9JElEYnP4JJT2LgDuLfvDh4m36
Ka+FFz7h9no8QWWeKaknvmzGtYOQIQLFzzPh/heNar9qhuwnzNR/Fs1XFVVqQKLP
uYAAvqhf0JJOPK700R8hUMCTJ1NFRcH0fW3c78gXXbkCovvevX/Y3yZKD7hSYrb4
htUNq5Qyax1UeeNMZeYh4+hiTr777EbEQ/pPDg9EQrexvE2NWDdkD+56lHljBHkb
iv/TWQl5XiX1IhOgl4hw5sqOPooBd+ubGkPU/sl1ILH/XOQduEt4WISko6XmMHjz
8pW9CCnMD42hkrXLotdPAmvrFjXiFurhSMk0XBvNocIXGGvd1o26cko/U4Ow3gg2
DYLp2v8j3v98eAjcFEfuPNleJ+HYidzYfk1q2MuQ7v8W97MbYYm8HZcKZMA4RAnu
LaEwJFfLKKHAUpcKoc34me0GhSoB3+BTQkcNN8wLQw+ivB8P3qQK3Yr1/zBwXRAh
C8UeZLZqbZaWFNQc97KvRn+3z2PzLwGMWsNqbJTXWfLCi4eH53gcok53MG95cMIh
PglSpSriBJBI33aiuLYm5sNRU8i+8Ikrdr4A1p9ANKC5OXENDQSOzjhBvpyYQsLA
Q6xoXIwc1TQ2IPULdzyvIVT1a+r1B41yXZfDVZ8djAQCYsg24Le4oE7u7PeIIHCI
l0AKEOW4+bjipMlrVIsKfyJcl4tclcEZlA7/oCtPH37OC2wMQMhn4VUFU5wHiDKA
X2ylznxvd5fcf3yozblFcaoGIWdP0GCdRDatFs1VvpdHH03iUW9J7CVSpsMNz/Br
o85XAsOdbCMWtqxTlk4WJfEwEDUUP6pbBa+/7aVIx6Xl38+PE4T8wNVhWKI9wWVg
OAwHQuA9XsFhjOe+InDawvE5JSaCxpQo4CATuh1/fyTA2C+7tt6djd0rkUBJONF7
q9Jkh7tvLGZCDruph8b6PztICv9T1neBumMUKsGNJ5qxJuTgrhadmT0xSCwD+FTd
bD9BDQ7aukEr6BvsF47slf6tThFRU+q8aUJhP6eMPtiEbCE5mVMCjYFxvtShlpDX
nX3P/2WU3n8JwOivNdNuV5bMvsz3TCq2E/8H/oDZ7og6UnB/a9uLCLaMY30DAtU8
aWsRNMfr1SDka8HhaFhIajZlEMBeM7bT1y6seUt1nsWnTPeaCRQUoVoSSWHbJyNa
rSUTN8dTv6kpKR64P0ZQatjl6hc1tUnVm/NG68AQbdK/k936Qc1QfZrlfJZC4kWO
c/2SEBRjGCfiuN7w7+TdKhIUgkMfyjZSLFru11NLHSMN4wd3+e53hc390vm/JkAD
MUKh6AMwNs8cJ4JS8O1VWn5m+k801uwWirUSJzZ1Blf+7+J0EH1w2I+NYPx8LQWt
Y5W6KD+GjHPSbMbNwHdMDGlii83VUnC7wBZCo7nEHJY0PfAqzqx4m3oE6chcGGFD
ZrGRex9nazOhzVgIau+HeaNRHsP5Lu5WpGXrofE7Ic+sqnmssVW1eA9m7bgGaFaU
oMgsqiejlWztPXl0k/VVWx3/WFOCZCuLIW3z5YUAGszNdj2Fb5XXqDuGVblSsXVe
d7jqFZmv6rE09Xs03OiX7REALpJZ5tGmFFD4toNdfDO+VPkiXceYMSth1xBa79oZ
KuCB1B9JThf5nzi3cKTY13twUNn1JeKGIgDNMuVjAdKxp4WwQ56/AWN0ggzuYteh
n5+Npca2qMVFc+XzwaWGhhi9i2I0zhyYtoW/aGK3zOh8aQvsb4Iv09veM2aAR7MY
EY0GSEyA8OXhrRQm/OYBq/zbOChfWJXnsUNCQaGC6kew+tKOsnDm81cMQgG9Sn4z
XcUa19zy5SVtDIS9gEtibMexWq3vX/iXP9EkQ79vZuM+hJ3MYuroKxBZXpVHXHFI
Ku5uZ2JK9w7KkSn0XxZOrcwnP4tpA7+o4pIvdaFW1NDli8zniy20mUo2HRIv1kOd
LxU/5/2cMfSf6K4/3GG5SY+DfVPM1nQ8RzWSEoAZgeb41hhIRvBX8VLayx3KY/cC
v0gnlYvAkUmtGqjHfAB6mwRBo0FjU/T9alNUp/0woNx3KfAz4SEz8hUfjoIW+EZF
irbEBAZYWp3nW0rQfvosfHQXsRXr6yVC1U4Yya4rDzu1tIujKug4VCZI9D4vgI5D
TT/GNRDcLVSY7dusPkSPLG20OgtAq4n8nD/BxJ90p544JeBg5oK7hxoIChja4L+u
AnizCl98mor2wQ/io6vq1FkRifUHo//lSu28oLWBFNOj4RZzHQsvqAC9wL19tALy
xwxpUbJwpqjNdueBhSyXtwjOViKdEz4aRZK1fgidsxpbRQ7/o9Ain9TJBBEMaAKy
oYPe2uoO8S0kbcpPzMjrX9Q4ImJjIr+Dp2rXufRYIk0yl9IgnU6C60sp0Bh6X0gY
p+ZAwJjjwC88aXO8DgyGs4ZqsdP4/4wTC2DhFXtCa6NfYp5VMXeiiPD/jX/b4oQm
txK9yzTxSVisB5MJUU7RKRltmmARvOYbE3FowsA81fCzxV7ZZWL+hor6orCAdhKR
YuFO8XnjkqdgGVHSUCcL2AdrTfGEHzd8rznNNlCzPaQH646h/injQTk3y2BkXL/E
K7RZUsms64OqxApQVLbiXTaI510+5oqXw3QoltEvyeq1Iock5LhgwixZtuFxXpYz
vZlqxzU1IYR9nZ64wcnZgrxFuJwbub2gaHAimdMQKZ30x/r5EOpDEsQZY2xkbUnl
Kx2MQxcN671oQQnsOIQ65UVy/eXhuuNiS2trXO2vI4aEl56DFUlmeUx08ocmJ5e9
CYOhpp2PsRD6k6xs52rEVkumwxkgADx8bgqP8OIqrcvJeY8pfMqrltP0NEvcJbot
YGhNrckPKxJ3RBz5b79bFmsdHVpX5kIrvl8PygoLde7yMgQEuGJuivPON3Jcv7Nd
Qp1pbsTK2aY25UxowQczrkoOD5xcQ778nyCzBTTYswqe0Rqy1H7oPCNkEtoXcwo5
yNAFqC3WwBV5NHHlRRJ2WBaL8E+08wDYK1B4p08HF/Q5mvllINIR9knDSL9aW9bn
TfNWpm9hvI5dD5/8iYezM+EWT6JtJQtUp4AtKGaroPLfTCloOkzhP5lOdmJt7wP0
5/prBgt7qk7pBg1fjVTrnwlIoC4+7/awwsaL6RSS9MdNzVrWkDjVct4T+Zx5tUNO
Tw9Jf3T25loVPcqqyr4R/HKn0R1BCEz0cdDrEjlnfaGoif6lk+p4fuZMGAlmFclf
OXwUCn4s5JcxeayF2u8lvj91smcWmFVRUAkhipio4R6sP4AlzNxf0cGcclYx2Z7C
Uue7CC+g6ymYUvmbtaZFMbQ3DYN826bMeFaTVBKhzUw1qdzbtN2hkkLuxJTHXKuz
SORRU7PMtdTFOT/HUOq76VFWtm+bl0JGtWXandyb0w/85hi4frATcKNn6AR6yhje
6D7aAgegG62rCxb8jOwZ8YqQNG7OqQbdUtE/swFS6X8FykwxzxhKrzlQq5PTBccy
738taw2mE7kLf65W9VMXxNlHWDGqiwq9IoJ4qkphFGC5VWqYg7yeFKO+zY0F1A9h
4i1JWOvqZJ7pUOPH53VdOtI0NqmZ3V7bQS6YhRVP1uwHocecP6+y6lN8XP60/xOH
WomZM0FWq5RItpyqpRCQ2fWWs+J2l7Sh7hF9FJNiJhX9OhuvyQ7e0QE8tjMjR1Km
1wsDx9hQLSfxOk7mHywF3jLmZdfBDw30yiiauUg9i9MmW4jzbUiles2OzhJjWMLs
2K/qg+zZurEbYGMCN2aVbVliJWL1RWWLlJmL5GuIJe6rijqvkQK8MkDx1Qsj/uhn
CeDIPyFlIiztWZozdZjyOk/3nJUW26z4C08NwMqHwATfSVEbIEAp+iucX9zHn9KM
sodyJ0PnZ2mxeUDpohEVeoFcYiRSiEnfh1YXdxIikumcpvEYo6YwJpvLiihMNpSG
iLI/zXNT4ajy5Xf+dDmH26w8jwzwNwW1+ldWEP2JvoV+F97zUf2G8D/geNmqvqQF
3aIQWNznDLs/enDqFgbsSQpQroSJaVk8ZC6XghdfxSMh80Q9IJh4y8yAm/gvHCSY
ayJVdO2EvYXrn5bhtdgJ0N8TW2F3BOz+bwZuDJsLNyEx/RiFWnoK1nVZUoc5idkP
/UuIYJFhMVlgL5k1L4p31U0HVEmZ7JcwB+4yKxJdfDl4TxjZkOURlBY/FyeLGY4b
y9pEHVf3RET4NBHbzvHnZwz4ir6+S1Y13zuuPqeNIVmBPIK2X4lFTHxiA74N35Aj
/a4PTGG/TkO7/r5y/xHyPmy8f6J5M73wreuPmR9lkY4EK/arpFdLw8RdyYK0SZmJ
+vQkoT+KSGzi06g1gEtBpV2ntzKr4ygCiy7HmTcr2nfjCSbNbPpij5rw3xlu+x93
lL872jw5Avu1LOL/0fKw/cY9rKuJowx5TRxK+MEZInZUi5a5tSw9wCCgiBS2uwlD
qs4rTGy/Et626Qmyap/frzkpA4CGTeedbyvq4tmPWQIeTrJpdcwMsSUHm+F1+LpB
JtiRoOBINbUszI8Gm5XsMtayzcV7eMQcZrFkAv+QvWS8rNaVQJZ+WqsJ5b8JVUEk
0c/W5kvamPNKEXQd02jA9mSNxMpc3hzUfPQRVTK1OnOe1f4XkDPlY71DQO3pcp1z
cYu2nrVV27C1Ee7yeadWxg8GHoeefqkFha2HHeDFBQPPtxAmSCKqBXdmRo3Jxu/y
Jr2Hq5NE7F6HDuM96ZKtNi8/5VjcoZJF3wzWIJoxLF/kIs8dxUK5hJUuTXUjhZ7n
lRuJznOSKeGElym3rKRP39/wYFLA6AVQ3kwmLk5JkJGwXepUFNdwZyanrmEsDYY+
YOKvrvyONzERr5mMNvtBict89A70na/6oyBVs8I+xqFagPs+b+LwUTPqX6/ZXVen
gNy+st8MOS/JV5JZP7H66dq9MrxW/sl55eLnPpJKr0GVTu7zu4Q+syel9GKGsOaD
w8LbdK/o4zJjUbnSeQROE1H3KtjpMnakrEl9DyXjAZfLdqlK9EC/9e2G5YNeds1S
lH1u1DP14ojoQH7Fcnj92imjzx597o6mnydKFXf4ZMuSvxF4ihG/ugsLl03eiy/s
veGk2tkzgvf7i/XzdHpGyUxOsKe3XpXud8h7auUseV8T3/Fguzk1ObaIT3AMI1tM
T2wiWr297rZB0hNUNtSKRVlVes3icfKNclq+5Qe8lnZvtbLrbqlCxHTwEfuzEKd+
G8GqZMIkCVckaDy9u08SdTDD0YGFhgbPdIC0p5aBjiXqHXInJZ7nnIxaxD0HnF6y
B1Pp4EUWlkmY2T8p3mJm/Twsa13wvdnvWnGYbqpNvxPM3qtONdycLNW/TuI+RxZM
wJwajV72E0+OVaCQSZ4W+bhSxHzhxajNmKjyutOB5DjJJMVp37eeggxoNr4qc8fK
IPdugWRoJq+hr0RsYUvicnsSUX/MtilD2qxIXGg/xLLe6w6EAHuVdV8ModJchWCv
b++1mPTvnYQemZtredNRYX57GbKr1EMqt1HBW1887TXcE8VJCCtCFCwI2VZZE49t
9PaifOAS355CfQrHkQbkioN2BpPvRVnU+P9T1RqHToOT4v7/E0Iweg0/4u8uVpju
2CBln574fhDvi1ZlmNS6fIhR6f3tOzFpkoI5ya48N/sp0GaSNFrcJx/G2lCltBav
EepVBV69UI8Evzit3UXncG4DAxquFCD/SdBXsSpCtIrwVe6586HQo+gBOCtwyuFi
DRsb4NDgQgcR9PCvd8jh819xqDkZhg3guZMq1fj3Kb+GOCFwLkFxtmuWthl0txRH
3Q7KVdApXgzXrhqLHBo7Hx1HukICQKMt3bAHZL7Wxy6blJse4hrutiORupggwLR9
HMVgFtyZb6+OOBs0veyAAnYgyzP957pt6+4dSeW6JMDEGttmfzseU5q6llxWsrKh
l/X1siOpp1rEl0xQrA2TfC2qBf50YLzkd0Xz4KVVJcpaVnOVt3gi9XnABGzO5Mwe
VEA/5ztFDiUlQzlnvwh8tjse3o5+WaxlKlVbnlVduNM5pcRgr4BQvkMs3LOeoRzU
1lZ0sqVvIOCErqfkJTKSQBQl2zsCwIs2kSSSg5u0YzMoerGwIJrmn+fayuvej+uo
j9w6nVySebJ75VwGFyJykbeQDW5MKJkV/RV3pzvzkQfTVCvQcZTB02y5TXLFGQD4
yl00di1eKADCkEm6SjZjpsMA90jY/TZgh2V1Ay6Y+v+BOhtps7A8WzCJIn7LOKiS
usUpuGPFvZXfQHFy3SoPv20sq12CosdbyvL8RNxhsib7gbE7YSzyGlZGCOCrlDh+
ABfWTo7drKgBaHxjtiKN93ilW17DbeMeICNBNy5PkmfqLD4wS0ExPSqEH3pee12b
NyjmJqfsHtiVcLDMT3VITH0tR4jg4gbh3fUTCixsSp7DRvikHuxHF1LX3B74zyEm
4E05OI/WVdYI2NLhSZiJPTlZwOPlsVy2jZSGdtwbQSKnkOIXSvPCBUrcoI1j5GKP
LettTYeI3VphD3bK1Na6gJddUwvYfgbTJusa+MxLC8Q1Uh5dyX3fEIgaeyCKQCYa
IzM+/3WCAkSm4HB3Zj3gFgdzZHRYLwNu65V1ws3Ga2Sb5wMDd3czHcLrkgp4Ih3o
bPzirFv4x7sCY797QqiqitgjVPzn+9SFEfQQwsmwfJ9zkzfPbYHyfJdbWHZAk9kf
gCVWebIU7DXYdjtzvpMp2TiOMYYfTeZjlq3LhqDHG/MuCc/r54RY6bMbjMGkSWy8
S1YRVdPaq3sErSATlOLr5Xkq5fPDWwvkc4xeRcns6NAezC0dl+nCZ20YNlcFYZep
2eimiVTGUWWbnDeOEAYylivTXhK6ZiENiZyymu4pLPSjyws0Vd3dFEKPVAYva2JQ
sv3nvNhc8O5ynZBOGJmsRm+iQmo+ErESih74TdZM9sgvECT6ZXl8Pi8RbYKOSvnt
Dvi7WiR4tKazAiB3krNW74rUDI3lMWoACFMooKk1l4WcnwsthAG8EIStzuafmF1L
Tlzc9J6QteCAJApNEa4yosXVtJuZ2tYMUWR3MblmSVEjlsJYO3qnWkRbdzdzA2RV
BiD2+RSYsUihQ/c6MUpjv05+o59HazsiezkKBBLp8S2qLCg0Rt90ODPFDaHlXQZW
TkjSQdO7yYCrM6wQ3tetYTtZzg4r8PfkZpKjGIrKmPPQoaMzMW2sqBAK1ShVPhvi
pfgb4R2abPWy9J0Dg8c1vf9lyDRno4SnvniM1FqWcRJTCl7JjrXVMrCp1klg7WmV
31TRA/m22dT3zsUZDvyDGTe3MUTJK2KDhnLY5JeNvIiu59HrWh1eG4bm86uIJz77
rPpvx7Y4SWF9PE6G5x3o7hkI9MTf6DxpsEYHfg72gXlpqy20aUaE66Tc24ruxITy
zwrZQZ9fQ/eBSuuMfH/g5lQ7RXYo5P+MWF0ehFsl73xy62IqcIRFQmTsWNdENl5Q
ayddjQa3Yavvd9nHSddQ5LKdFsJxtA0Ye0Jbmw8IoJYaJ/v1TUauprRPHJ+IqMvF
2Zh1iKIZfQTxijEPaTJw4bvYJT7I/TaRKnprnrS07x4CdBYiHhvhTmj9rmB2Rstb
cHPB/pHoYXJs1cJ26KZxgTqtE4NmA9wcMK1u40q5sbJKWZwOJXwG5Erw3AAUpbPF
l9WUpwVSQoXaSXVou/Vi8eAezXxUeZCWh3hod0c6/RQb1VISKPyxZnqwglZZWLZ0
SysG6eX/u86p+DCCmcYA+uE4XwOTTw7qpL2CAY6vZA2EBF5s/cuCuWP51loy7xiJ
BX59s/dH9liy75hO2cyrfx/Hnioz97ZJ7lJka/f0rZ1fE87I2fuCeN5O8Z0MVKYf
nrrDoLwHXsLzq9DwsRHYm3/NUAwwer34O1jT9oh3F7+5wM9d0Yr+2No02izaCAHp
RL4VKRGZ8GOS52US5GptU4zBef4p6ImGFFD1Bz1HwTqilbQawBeCEXQzL/ntoXGm
TkCKv0t/NQLaEY/tCaAyxaY2NYhGeAnBzQxzG+Iqj4XHb/7XCNVS3kZWoLwqMJyB
Q+CcxqRRCVdvX254yU8cfUTmjseI8gLxvhXJd4aWFPTYdci69e8uk7BseRvzVfCC
akvlEUHkIrAG0IHDHb7qxo7q5eR9gct2cGYUFLDLA7HA/NETZsAHz/sFFjSumr4P
EdVGWIQZBbyF+jsNx9Xzp3X6oz/U4iF2/HQWw4rMoFJqv3EnvwQEjzBXensHXvWR
dQCszYiRYDy/eeMMosSkg2GRYDcmPBcdzEtFBpvFy2EL9rH8elHxh0Q8Q5QexFg1
okp9IzcOOVZR7Afh21wPsLqN4tE/j5zdC+JlJTzVr/K/BN9ufeREFwRB7MabUqNU
pNkDXfXcLnDRie27noHI7k9LUd9ZoXuNtcnUEBWSFScwBZCSSmgRyFC5AoCQRZMM
bGbe5f87G1ab1u9LUy9++jgJSVDy1KxVLNw0N8MM0tkdn4TZYPAtBUPxlJbVs9zW
JQmh3RtHZQDykSI+preT+TzF32Ttu39UHVil24GDhA4PpRSBDIUCap+xnbS3xuKR
71CO4xklIUucJ7OFiabGa8POWM3t5EyW3s4OKYbZp4s78q603o6RGk0pRLcbauQd
XveW/bdD3se1QHEWz4cxGF586TNpVB0/S/vkqGSUM2VomcyVb2SpXJF7UPeztX5g
xMEwm6vqnrV/7ozalZB2Eh2+UiUiO3bYsLfOupYBjY2tnuZleU3lh0MNdRHsXsM7
Klfxc7sRGcXlQxX+fsI7oi1THxh5Sk1IPGkgTtimXFiVci6usiFDfmMXE2e14lMR
Q2OQHBokwvK1p5Cjyi+/hdw1YsM66bUUGNYMESgjLWgirqxJb/V03p7GnQtyovnW
tvxUDBBtb+vFI9k7VPF5x3zRp3hCLT4k2ESs3qL7I8Uva//pEF2YoyUw2Nu9fC87
JeS4VBFy4ciDkcoK5yt14x043JzD2yASpbW1qC8TtoTQW+kssQxWWjCFzdWYn9mU
ZztSXa7ifAN1llMwMxJZY7ploGY2mIQ3PMvCyBxcoLj5P7x35L+o8RfwJXapEXLk
mckf/9+bd31qZeYVhxPBKi/AanYA3sh9DXJxIsXk5BrzVX3MJ7bj2iSvPk+/L4RQ
I33e2cYbO5KBOKpSOvbHLDE08FtlfM2aWCvEiegOAi/6FTsNgC85keCDwbAzaku6
PWmGldb+9nFZfJ8Z+wrrRS7/ofk9fdOb+sKtzf6p3aJgzmZjE4YVl4HQG0uiaXkN
ytzTJADriEj6gMROKvthQRyAaogDtAsBWVfND/tWr/Zlq12esvTj9kk8mNF5JbcN
8w4r5MX0/jHuev2eDnNRTISUyC+V2na0PbR7PKSRDzr+vDp+GK7p/B9ZxSyvSOW/
/PLA0yZtWbKWVsg24eL+2WdmFju7SPrw7Ndf2H9kkCMgOP+2cW+kcrFp0jiHgOYv
pFPgC7tV8uYUjATP5TKGMQ9d4j2Emms53LV2cLJEEMmQPAoDsQ2QIdee+N0tqnQk
A2M34fD82Bu/NIuheXL7mUlhK7+AzMQOzI1bqmrf1OzFLAiIdDTiP2uwnBt/Mp6+
qmdAbTaIIbPXoqLv1rr8oRF8lryRzbjhm/2SORnvvWv5WaepivY4FC26bRufRM7j
n/4Vi2SFxLM9t5RZ8wSxQ3iv0gIG9Bxo97tOK+Xynbe1BtAXcMlI/z9bTXob8kJA
YYaq/3x1PsP2IFLFNUrgIMUv6bJqnRHXxFHL9DucspJTUHYo+2TNSrLBJq1wXGFJ
Gt7vNcL67h4g9A3pla/uicWqWaCvETgbwvfCdr1gjdae9vBEbxTj3eVUvIRFuJAS
rNxpnPfYkjrVSvJ9AkPP+QM8qWkOwdgseLZJe1sKQZS0rgcgJ6wfy5SSFGUso8w0
9Z+Zakg4Pr0ffdxzEY+9o8uTj2BuucheE42ugpCnJCCVi/wtfA2+Ta/3UOimfFVw
vnwofzfOyv7ermsXu6WHU9MZMnizXvcaNy/Fz2whPSxYUnduBpNQp5Aafq50LWh9
l0gLwZ71mxyO7OKRdyrE5ut4o6LSH1cKJFElXTX4PRvshIC6dQQ4INXtEWp+Zpu0
UbXfCohscyNYJoWXhJ/ik9wPH/slDJO54DBwtXl+0MupXdRtqv2zO3B0KszjLcac
sQtFLQhwq2fS+4iyTJWEzBtg7RVzdI3i7eH8qqNHa4hCI907umrU0wzzIJ3jOP3h
fLW9MytiKNPEdNYQyocImQ1iR4+iOrqzFaM7pypIOXjOP0rCjUSI4uMqD5Dnkk+3
BNfGWIserU4zr3mHYMvmjWmzxT8mpBuaRdPOf9ihn7u5uKT0MCI2JLFbtJkHmSff
YXF1VUiHEaraDmWvToTjUEJLNRt9h8BACMmhympT+QMeqtnEt8Z65zDoNF68pQ+P
BPG2zXkciQ2WiDYpiSSSDGZi4edLsiqPiKexaLcw0fRRgjryIhb/yqZl1jCMLbA7
L8//u1QgDZ8rZwg+V/ToKbecA0mJxbdImbZqkbftyl3frkuyFMn4tAJs7i+97qTW
OCe+Ad5PHkbkTg1iqu71tcRDHu/8cPFvAiyA+BSwqo3UqPRb7a3DeKPfheMMbnBi
nEWpYje7HSRHVSel1CSfMCi9RuofjLZRwO7+GqXvvyOrNwj+MiOf6jq62dQZhMaj
8LKeOIfIu149q2rFUliPAvoGODVeNMFlJ6RlbFJf4Qm9PB2KuL6YvE7xPS/cY+Iu
3OcbmIu5SPeyBH88vE/zwYAUytnbzYf20wCf1XGfXVZE6Xpu8oY2Z4YngYxfQOyX
SUouYf1hUS2DEQWMQZ+7xJd32nS2kYiiSLygtq/RfgJJit8+qxXEq7I4zP5sXQbg
rcopwrisYFr75EfdinkWsTOcfjPMnzpMxSIds4Q5tm9Hmv7pbpt505tImJVBFco8
WlBCWrJVlqInTT3aX97x2kw+e0AtSEEPZMkDQmstlDk49+DUWRdcW82JtjS1NZg2
Ijhau7u6oVlYUeV0u4wiAp/k8s1oNqkJ7dHlyBs/S9i4PsWFTys4ifDeDq9IDgLG
pitWepztldtT+8s7uJS/6meHpANFsBUF3W+Vi7yqoY6vvgQewNd2AhzmPio/C5WU
wN8C7o52U3Kk/4E9AdANSRTjg5bSzv4DYoOVFDcJPXFUDj3bfxr1W1oKHPzaLmcG
LwNot7Y/jKUqqx27b79lDxf4/IY/BZnlfNQiNHZFj7KcBb9mMJse43hUnjOr/+VU
uhfOxl9AGd5yzmbwnTs+3qOQC5ZD+UQ53aAv1SPd5HGysvIrLUY+1ocwipAKvaBY
ZZmNcviTpyWp+R7LrV8Q4i+Wrq5JaAu6lMRQ07L/0Jbl2oLTTSOnzpMDX3Jzfzre
L7V9i9pC5ClS0grGaPNGZH59j4+wYsjUqmRlXuR/HCHy3hQRLTOLZoBV2do9Toay
+fH5KLg7s1lR67++K1JcgMelc7k0K5VRFB1wkSiVQOAK/r3xGFIS8q5SeN91YlsT
XQo7yDRIaW87IT6XCBtgKoucLXNHzHT2a5Jv9+9rYoUd/WU5GNYq1PW3KucjE8vP
VvlwDFfg2AWTKzzNTYvpbcgcX93YQQPCo0Bb8SEBj33IwdEefUpNzHT1pfluG8eL
2YRGc4SUsMiyhHlHzQJ7vkZEnvoRCA+oMPmejPhbGYMZuC4BwdYVqwxx1wQZve00
NdVKfYBiLv1o3PX+SKFvAvbqHVuOb+EPvKIC4PJh9oETRdhOcW/BdKvU2uYe8+aL
5gOTYzGN7t/ADfuuvj13tyK78lI0jxknjN/z5tn0035qp60ZQd568l9S6M8fK349
12oJG/Maxwmd9W9edTZ03A9zB1KBuS+Q48IV+jjoA4XZsH5j+FdfccG6nWalPKw8
huOEuMY76MQM+CAy16oPbM+piQlCcoEfz7ruDWtdFdcjl37DuGEf35EtUCE5kTHi
N2wG6zzCQo7vsRCwlv5mJcviZoaEyuFt0zEXgKWVHtjCbef/tNdhQ9DgGli3Jl9A
FiWnIzeiQ7p+DNBNMGT0JaJlzxGlqiVgce54k5Ho9y1Kc6YxWhPf5YSQBQMtCrCE
VzfsEkPB7htJ1laiOrLfFfATbvhHRoJqzxBQpNwiZecQQwyFptamYFLzQr/ofRx8
BOhY/Tc3OXyRUYIYfCzojXsHCsqLKpzDYBnk4TZCcsOPxe+Q2qD6F71HlgZw0PWO
4nNi0fEyys6/xslDVaMe6MyMPrgPJQQsLFUoxaY8x6HeArvBAywNdaxMNNBcKsZ8
2D8RSI3JhUB/KbAJiNJvZscPc4YE6OFHpv2NnvE/pKon5zh2H9CWJ0aPFdMyYtCg
kh3ypWG5l0WH37/IfNbAOaMU7r8vHdvCz+3esVeHmWQoIRhL5Qp0p517Au3j0qiw
bs+gAB+Soy3/KdWkXpCR1LI/ilKTzEu1AadyKaSeTUyxJEoQ7W1rtinKO3JnJ5zN
BlyUTBdrAL9TXSajRpcWfOIn8JFOdN1TekgiMsFYm08Y4jszpzo9R1Vniw3zlXRs
pua02A8ihvDgRhrqQZgqlCTCfLkn/DsqU0tqK7WyM/61w3nepwOZgCAbe/hi6Vmd
lze/sa2Ser9NDtErrSDNUxFtQhOaxDzxO38yzzkMqtMKgGt4miZLzdpQh7uLe93a
+Ade4G5O8UMHHocs3OttCbAwfCZ62hhr9aDuY1g9VQUOFUdzbIlFI1xk3VXLcM+i
vb90jUfTkTw9QnlG7FKBQq0zpSm540lSbBDPSsTWTFcE/jE43djjb6VFgV6WVuOU
4uZOa31VKVcnCxqnGXxDT+8XxIwxPokJfQVGn59ZDgp1cuc0/XsMVz4lpaT7qZn0
vMQTUGpa5yUtfwHISOMM8X7tZwE95+ZCi3DupJOwe7VKcsMBZwoXPTR5tPm5MX8B
0yWe5CjF+tYLEcN4aaBYSJG2Pkm954Srq7refh+5cNT5UpZ8CMYUtRhw0pjOriFD
U6Xz29DJBJX5yYRpKc52/tF5TMb4jsVgYmE+wyVPXm+uJC8zZ5c+vpdAyIox8LPY
dUzc0pJw6q/FgUQy2gjkF+piVneS0Du6/SPnNvpOcXwqkKxxY9Q+AnlRZhakmHX8
GjImNXphzzwgDKXxsYtzCDSFnFZEVepitmfCK2aJ72CxpcLRbRQ7C3WNJpfki+Hq
7e+jKK8HwHaAB7gThoqDZejNQ+WAGFt1S7rC7hlqQXfdfRJKpnpTCEDkGXy0AJNk
/856YqFvB01OtcBc3IUTUp+PzrOrGKqzD1OVtC3WCMVX0eScjuPJbuxLYr1jZMyn
EQNWvmDjlo+MHSlC1FX2b9z9drN1a/g8rCIQECdaps1I4q54J7INTiVVyp9leAEK
2liZwWIgpDezSes9aMkrXWZDjevVix6MbNqfsga7djNpEXYjlbvbOnF0Y2RloTDH
i92e4yGkvgqgTP0+lZrZk3E/dC+YchpUG39eNjtgrHtbpIryE9aeBfhwbRchnDCC
fCugc4IznpIgAA8p53XnltmS9BIqidJaAfM38fFPyL/pOzagdkbilMp4FMI5C92S
Hru5ij10QpxqffiY+tFzT5Zw8wZ9/nFbOp6JqRCQ6L1rkvBRhJi58FcbNhEinMZy
QriP2s4aKjzrWsSexE0QDgQbP5FliMUWxwjCGmf0M+0B8M2sSZkOeJc9P8AvPFgo
ns0YVa0pzjSmMQDJIRnuTWltqpGC2eWqtjwxV3nKuqE7ZcD+Byhemz38dTrVGPz9
QDeWWvrpmhBT82fuAAjwylyTaIb2n/h/dmCLAUNiPBlGo2Uv2V4jkC+9ebAp6vH0
VUhe31XkXfnakGkHqkec6vapPoxcDhCodt/yw51+CpXhpgMo/a8+T9QpMVELZnJz
SlpdkESl5GgXbgAP/B+aW4OpjtzRsnXhkqwv/NDg9v9qp1dEI1g6LRKKZhgzT/y8
NatCeByiF/qz1DxIobmE2UFeLQYG0yvfT2VCy157az/io7YNXYkyBU3RJPu8NTIf
CbDwpeIKrAuoxouXbcTEDny2PAH2e+wWLCRDJgzh7TTPXtu6x8TKC3iMjl/qXYZ0
HyjHbXl6z2A+2rG3+ikbP4GPxDnetlN2wbIeU5Y4E/3I4KA6JNOkJzZac0sRkXHk
0yImPAAcap1ZTDyTfsz+ZrXWdY/YsvcSvwj8+QIqp0r5rLh7i/EKg2L6e/ugJapo
2SPQ2gRpzFoHwDAxvlPmMB92/APz9VcLbMHLVUkH9LGbQMZVGfmpiagVpTm+ZUPY
fXDqIlnlSoAX1O6Ucbo0Sjz7Z+G6Al737yZ/ogkQsPn2bhNVzdwac6/zIdyDawPy
9r+izvUGafhIGxRM4Zx1s8IRgCEbpBXFQ+iU7WnO5QAlNgWNfYw4ww96N43scq9H
Sk5tEfWX5bfVZ8YMYkpaupFCzOUp2XHBuNOXECZ4SERS7++1RoGGG9Yec4kFJ44I
qoVTfmfO2dNAAUbGGl3VywdZeSJNOwSwjmmHk0PDWp7g+1a2oUk28rKpTYiVrI6N
TBOstEvuRt6fNKq6xoF6y0IMm9DvXKRYyN6+GbCMMtHjTV7iTTT3S6Fp/ty6l0Pu
9vabEYdDPv/2BTZL4DNzxRdSAVQ7fhAapIiAjZfVrpevCq8AEJq82k9yCyUlhUcV
nvewU9GzdXgeA4SrHvoppy9sMxPRsGyO+IqPHshnVBxGbNpW1tq88oodedcmrzp4
sLRYNqgRl8iyXc/MqoqgNEMeknvVI28C1YVcsQ/EDWj+QEZwUb2n0dLnuWv0Ng3h
kT1XJ+DpMvdfXXuGTQwQz68UYzbl6l0OAOqWDR6ah0FBPcW3p+fNgIOVhHDsqBAH
HO6m0IOdwSeTdGBSnrrMNLezlOkQ5A1pSpUwLjOcDDsmsG0bmJLNOzGOjZSLKiSp
jBclgyf0M2iAyIqJ/UZhzcst3wYe3963CzbkPhglgRBf4ZWeqcx6Wglg4TA/UAiD
Ql6ffmN7Hjyk0jPw1wrM9jb8t9K18EIqcKSlbI9M0W3dJHOvUVoT9pxU6Keq2tXD
1PpkMZNJ4Mo0pnMQO1FYXalwDTaNAf9xCjXpApmRnwkB6z6alBY45rEMFwg+H5sf
w2UKgaMvAYUbI+mubf3I00NIjfoVxpSMQjEPsnFDghb6t62ZopA2z/QTmaDYhby0
sMzCMrHFHtc8DyJsjC9Ymowq3+zzbWinLDjfgf5LSYToWBSwsDeTPerq8hvfzwZx
tCzokMmJBfd9+QHsdLOWpJR+AAleAc0ZX5MQRcZMFXeBlE0FCTG3o0S1zJQt/U12
I1q3Zw/jfO7nqfA0aTNHSi1o1WLaphYwtiRzPRNExbMgMJZSqEzufPxoUMzJM+Md
VYnPzB4wt1ljSegqPAImToGPYIfWknaLdZLKfmlYYWbOIIQSdWoPuYYeV8EQvfoJ
WAGZ1q/eiMW0OvG70dtBg5wIW7l0tRx24dt16lYeVJOOSrPWxOE6n0XDrzKtiFox
+6gAZRRyy7l3uWgrk08Mq7fw3YyFUzZi2lFDeUb9539XMuvp+djPhQ7qSJBc49QR
H8frrpTamto7HTzldUj23fOkWrHkvXozKo8Gfgr2UTuROoHsAHdZWbDugz1at4GM
t+w2a00HCialvyf4gTwP0SicxvwCYRRXs9BXKcna9a9XhoYrFgLDuEhnUKGSK4ZR
ydWARectMyzAQBdGPucsIELuR7+Jih6mCNZaVrLahmk/HQ+3Xqw7PhB5FmS8c5LH
atZy2LvCyqQQEY2q99s19DiL33E9j25Gbwdn36SZQDsoNqxKhNAjX6DlgAa+QubT
Lp0y5DDw1+vHFSC3RxsW8OcN+cQYbRpLCsb75WMtOgkKhlAPkWyYnifsTthkbb5W
g1tFV4OYCrYI6LGdV5kec1c4IuF3Z1b5haRZw3gHysi2ElTXv3C5URv9yCLl8UyL
80wWLb0w+pfhaAnftLgsfRF3DIctQeulaRAtKcKswDa5Tt0sioi6BreyztyK5DcB
AZhyCpjAHIkXhG1Edpeh4tvaILZDA8BV9FrUL/Pn058UJEQNiAENMEKsN5mk6qT8
jAt73kb51wW6UPkp4dVbD0jARWG5d2Xoov37//wE+/PqmQMNjLXAMZqZ1wU4tCd5
FeGJVAgtfM1mP/JccOLXz3gcBUM3RVdFHbTk98rmxn7tbAfeeiqx9Qo/qOJ4X3w2
1l9BRpcHyG0tqUNYpW0Pbp3iS94itWkOcRychdbQZOn0v+18dwUIafUvH2V4iVgK
20qzmQdkSDyAWIsrybDweLbUxFT7J/I9jb29e4osgUrcW/BwEMcnXS1PAxpp+vGE
r/QrrlPCrtS3bnxAr9DsnbwyMiKUSbg72HiqgSJ6DdPtRWuB8BvbxT8wUxNaOUvD
M8ZSuaZ4NBhSirVmWRFJt+HD/Y/TIp/VyQfDR1ShapjCl9zInt4WfD/4bkr8QTYo
5fq/RphC+I1rA287JfBEAs35K7rqlGCn4G3ukFGyG8rTnIuJ51jt+ncxzXE19swG
TPo8MqLoOYVzrYYc9Isyo3jjHGoISq/i6m8ywsZbAq0lk8WoV4awIN6Y43QvOtE5
c3OnHgIHNP6BM2jK6HXQLoxZz/wGh1klsk6cV9Mp6GEOr9mJF7oIwi7czofI/en7
3RiloOzus1HJ2zTYPmM4f+M7OHr+njUZ0XmiCWMHe6eJPwmWAvnQpEfqVpAO1mzZ
X+nsVUaJ8T/aMbulO7+vL/e8n/AXeeBOs7Ge1qQmgUwpkbyLqfF6V+lbNP2zFqBO
SaNxG9k3ZyL0G0xTpnW7Wh6J3wmfnpMUoCiYEah5UjHLybVnBLOmBhq13N9FXRxQ
/Xqf59MQRjY39WZAOCnIDJ0DrvqKZt2J26NWqhz1pRWnhEOKXroAmq0vCA3Lmpet
drKt6URc8C/qxRhM57MJifSJi58rhWCLt09MG0VHTmz6KKRaNwWK8wyx7dfMfd7o
ABvGdlNE3K/s3tAWN7zA2c3IXT0K9dPNmtlJKo11Er//M5YSCCVT1rxN57FYXMJJ
wO9m5/QC5E3mbpPNrFSbRAM5QxHvXlbpO3pbFnf1zM8eq+8i57wIC3XwM8p969eP
TqqJudnu5d1IQw4jnRRDeXRRYIUP8Ve5dUKOXWzqTCVpjJAWPj71wcfdi9gUXeLB
UAbhzgEq08kil0Lvuxurdng67Kqmi+qAH7mEjZnsHrh3lO2VViawcQEJoCfGVDI0
b+L24GfP9Lzpd8PNxiWwB0YIF/pOzg8Jst58uSYF4oQ5y+S6G/8SZlJtr1ShVfAM
d35qOL2Q6Y19VG1OCBCZqWCad4/MV5t1yxdVE79eluUuGvfICHsBMo8BoA3zPAy0
edR9Yix9+Qv///MKPAbqfvYQ9jBdA8fvKmK8liZisXAwwnuv+n1UN9WoaQiOTjGt
5usQDigkrsfMnXLA3c9iQqvW+Z94IrG5yiz82Eg/YpitJzsRwBXUVFy4VVc3quE6
nDJs3s3bN7ynXjDuyqOqw4uFEHYR7nrzUfWKbpFv+opNZglSM/EMf5hzMOfhIFco
5ANWwVwwytpqeqcEu1bRp8a5eVH2uHRXR9h7stCbptSDGOZggpVIRzRRCqqfhp7C
/iNaGqauaKIewkTP5mRhcVbYuVLNbII3S2aDOvoyIHfyzCO/X6J3d9vHbz2uqBF3
P5n1ubICXDkJ89MIGjdFLSscRgXIytxFFPMXdwtfZr1UzVEkFVPJ3neRQs+w9eOL
ym+qdInL0dUXs2an8TMlAYuUHbCjN5Fx/BRcVVSI3QZa5NuTLWlk+6Q3Vsh+1Pmu
sXmgit0aWnksmZXXq+sWXXG3l7lBnDz8SiUGxopXBtGOGkR80P/mKABgu6XMEPUh
rQMQQA2FA80fjTckYN//oEg9CptRkKE5zMXM7aJrH7QPqmTc8bWEWhbMdSol0lQE
rdQAYL04gZeFfw36zP83053mVMsrKwOXyk7C3Q8CorGiIBnUqhJ0mqSI+1Dtwy5r
mt1WeLv1oMTgpB1NuVjgy7S0CwQmqyQKOeXAJZTPHpzXYmzWQfV/zViMhpZxGp6a
dCNa7h+Xs1AY5Q+pNgEsuoHbbudD1lZgglx9cduEcVe+MCWrU+fnL/Qy+9honzmT
SoroJ/OhzCU4Y0f3B4+QnmnZbrrjlwLUkQnJMeDmpSaMWrqDwHFesLyOkWuM1EuS
J0MpFYFQST7krV7rdNT43Xgxf1AOxwdzTsZ6YIkQ6bli+2t8+tdoWm+4NWRosKJU
60ywICSrnL8N1bp9xVsDYzvp+cETrpSpuT1NPiLmRzMpUvIN2NqXwh6NvJmBZMTC
MrH3/2GKjYOUpMo6UpDzg3WNAjxsj/d/pP3UnwmUFkc9Y5b+sUqV+5krymIBq1Og
Ji+AquauzuSSzoQNYyXs2c6AQ3pb8ftC7Wa4Aqp9qHAMrhIXbm8F/w7tQnCTPq+p
oxKWHH0Ht3eTMnmcbdDXZ8aVHlB7iOH5mGL4VuAuZ7EntE+0hwTv/DDCUmWkwYuc
vLt59egAVi+Q6QWTNDVj9aVr4D4BDQIJcQSKPY1jpA2/kYW2c2JBkCccF6dLnz2e
zg9Ax9x4+DUU3e/0WUv4UdYAojyg4QIRornbKZZcZcA+9wOzie/QGxoabWNj5kqt
V5aCNYw3B8XqPUlvSW6v0TNX26+EEuNICJgzlzOy9qsZpVxdA29OuXib/77YUWb1
CdLxkLR9U+arRlNIcO5UOwt1PVSKHqK6q/NO1+Kxe8We0Zc7TyB/8z7ptNNFodPe
0NeXmnS3r28P9w0vm/ckpR0HBc8f8qkJCFgoxjp4JiyldO4RPcC2RBx9c9KUXcyU
baFSztVe1jO2Ck+Spurb1WOfN4lQDgChWUaP0tgzYec2UEChipmiaYXMQlOGdqYb
rweM/3w+hZAA+RMH0RTv0BX8+KmHXRcuVoidoXLEUkRNlGW9JppG1I8EIw7Y2GQn
fphMxoYqWKQC2YNDmzf44o2XZOlBGlX53qzhvlc0w+BULkdd5H5dRtRsKAyvPxyO
PX4a41LXmnB67sFjSLRkiSP/eDcCXi1QOsYlH+SttcWQdgveYS1qytrjEy7AH4EU
PZj+ZSb0q7ZD0G53boyBCBNVU3ihyze7WTGxc/2uyIKecWMm4yz8D5VV5nuG2ylT
gkovDP7x/F0DXQ2LICdxWUgUQOkgEwUtGsHco20VBVQJWO58fOf5OYWi644mVSEz
IoCjZFFayFYWqXUL9x5D3Yc9PbP3X4PPhGUuSULZDXnmSzx3M8HveCncz/hyHgOR
gUnpbNqRaBVlpxvXt7rz2OWJLhhQEKvAAVr9BZ7KgxMtqxVEx25rdtXh9m8+S0PW
AEruDNRsCrTUUOZxxOAQoyDyOt56YxioPyZFn62c3ZqR9J7fJW4VayLQv2NBWHtI
FsAWv7lDuGiU4kqT4fZ5+PQTflQ5uOLC2ICN9EtX5n82fjSuMNs6el0Pmmx5UYay
Quedf/4tL2U0zgXo18UzKnhg9///tL4/WvY6eeWK0zCyOyTlIqTWsNCOGdJco6Au
DCE0KKzqWh7rf/ZjsyyTpsJiqXQ1cLr6RA71BQ+A53QzL7Dxs4pPFAsCFlWqieD0
ISG40bNHRZphKh8DdAZCPvl12Pl2OJTMP+bhzCadegau79RSq42UNfsM+YaBVc+a
Cz4DWayuHtEMauK6n+yhqRM3T8JseqRdY7YxD7/BNfB9/AuEfI7mja9vguh9VN+U
tniQmGTbswVLCRavN3LfkLJswP5jsFUlsi6aoXyN/fM8BX2BcmRZbXgB8YW8jcJ+
XCjaMEXbMF9lWN9ZS+x0JmwdHamrepznFAbw+d8GXZaI2ccCkcSNdT7lMv4D5IZr
FT0yRT5dxZ59mTYzdVwRYkjzq62UOsW9fpxdwfKmON4ikH9xqLGP81W9dGApTte9
1ats0fNj9BUP9BQmB4fWtnkAIAiMuwrgaGmnvr8n0RRvkdIPORwBDRZ6lSl5Q4nu
x2tjskW9Rf0vx/0NT5BDY4nveAigG5yflifh+VIY67oA2nYuE5U3EZoLrGCNZJ2N
gVd2pbzypkJpzI1+VAURC+eiOalQnV7w+maLSCM3G/ft7i+if0cT/qJeRIRV+CLX
UYJQn6c/JK7BoEzc4ho9yme7WqjIsHR2NjCJS8Dw3jc3PRHYJ6XsuOE7/dijvfaj
dA1Nvy9I8meyapQupiwpNZApNNtYtNuxcc3WMayc80VcBZyPzg3mOZaW+NlYXN6b
I3lMN2D/hNCn0HKE0rzME4QSwaHSidSHLs4OTbX37CAtFW2prkzuP6l+moIXR5ag
eaKMYqmeHRUcotF/ZyO3bthmgYpOl4ki6JNpbgZ2S0ynEBMn9Rdi18tvYx3R/vAU
bWbIs8pfMiDS/jfUyyScW1RYYBxAgNyV5ayl1NdjzIgyKyRxjQJO5sTDctrmafZ/
+dlrJoVfqyuP+me3qQ3le8VYHZWzMhkHXri9cKYneG+P8a/Ztf1hxreU0suQ2Pyo
SgdvnTjr339TODnvWEDHu3EPPZeq9KTOd0UmV32oIdO9Pwc/0flKpCnNPi4h1Vvn
G60wJ9/E4jzyOqpbMSgJawraZysO+f3M6kHc0uell21lVc3yyztYA0HTZHTHuHEW
OwBUAqbkulf9xPZHlRpVwHqf1kCrrCBmtXZBEur8WMCRWBj4Mluf73INgYhWsqF2
lTIk45HxKm8RkftZX/xYQThQvjE9mAEli+d4N8SS48lgW5V2F+rNfyB+M8R7ihPf
42QLQkfKUgBZMIkxedwm/GYfuGik89+0faCUQEO+Hp8/2N8jhMVLORZ2UnAtm1R/
jcWfSCkGHJK1OoVNEy+05/ojBfEGW2hVRTkS1H9pwKWMa3ENmmAoCvoMVT7/Qc69
yypof6IoYsGgG0wLLYWvXEwGaBHeBv6JO4D/cU1EDNO995snb5ndlIsFLEuI57yM
C+rtXTOorsssksEPtGFUQiQ3QO5ISfuVkI4P6Kwcb9fwW6UQ55O7U6gC9uX8IxVC
qAIE6lmTBdDZta8gdwgLYixUOQnY7h4EpDQu1qqk1EnRB9glwSb9OlynA+1RSO4P
rH+cHXzEViq4QMAHUgDSUTrazvlEnQlT4lBazIUqN8EDO+m2KIQ2HgXX7XB3rJwk
oh/YdgcNU2rkrXjGw1pfpsqM5THM1VH5vyOeQVM5D9+45Vj393nbqR7Bz8KnaS4o
yyOre036sWX2/oCTQA4HF/iX73tnkCutYuCGp0+ZzZgSXtN0ErS2CTYXE5o7TJ8Y
zEg2lV5QXmLLV8P4EnsIFVOa5dFfkmPX9OhsqUqVqt7lJStZbmaJ9JqedAgGzZHS
PGF2vYtXa/Nifr2dHUplBIEbBRUnZJRJvP5mWf4L6MZXAXxYBpAebHhpfautRcrp
wEoDLfgP15uoRXiyrUiUkGHRrWawyzMbfim4huyyPFuzI3SC0/73jx2em0a/K5KH
4kHccIE2yDFeOH3OW76eWEaL6vnZ1bcGS6tLvAAW6yyr4WgNchyvy+he0tWxrUh9
r+pxtKWEANkpW1vh5k9I63rKI4LrGjDoS2rirgU6a3CSSd6c9xyWbdjIjePbsVl8
Vx3jdBIj6e8d7oE3/AACy9S27Wil5cwaCWwfkYW0sNI6NiBKUIJ9wS45olbEu3ku
iGv2fe7g9GXJ0rb4TmmYkOvUy8T+4GrLM04j7ZeiBohAhRliYL3AdRMdju5i9gwu
18Oukw+xUqDP3z8Kekepj2Vv+1G4wMqKpEktqhM6CDYiX4JNBZr0KKQ0I1j3Mfcq
TFKl1MHtCR55HoqekiJVsMGptoUXXtzaFifoG2859VyQNMJ2+qZSWvIrxFtM2sdH
jIq6tM1B8HB4PWK3J9Qutbw2VHV4LHj6BvWUN0d7FNfMpQjMwuNeYGi5NzEg/b/K
TYyECJyIrP3xZlPafmb6hZYE4c2OYi7Zx5bRLtQpFsnvIoI8G9Wzb6rkgc20TU1I
Q1fcVniwCnIVmtKRHCdFs8IDOgBcNCZn7hxZctoxcU11aRccVBl+zeZWHaDEhm9V
MlX1VUqCGRkHkH/KE9HV804OdYY9WKtYNudo1B7as8TrrX8wVrWAS6KwMXNvHifM
vklP7LVmFJ0ghiZ3ZiK9fU8j3oSMRds5GsRzF+wQZYx5JjmlJNZsY0RmupHlGMet
y0oz7OqoDfCCtBxVO6TrDdxrbxUoDScw1S81LmedPU6uURa7gmb/A8bXtlVr1tpE
m0+XLRd2KAuI0Pp3/m6C5o8MPv2fKtaWds/1BA7aiKw6gA1RG5Yqde2O1u0lX5M1
ihl78GRLfWEjBhz38PZ5FQQ7lwOinKb9VMDyFCBZEM9cFYpCmEYPRbPHjbcU7sb5
IENZUWmMiFgT7eZx2daajKtf592FkE23HrC5abgID6tZ+ag8Vf7NZJt+IGhS6HJJ
iYJohE/Wbv2gOtAUrw9Y4IdbStm4YWVrt5QCR0rvSJHBGqjpMtgZY7Z/9i+uDdCy
k1/vizrqgBJEiFfuPuSgihEUZ18cCyzzxudXwKW6gWfq4PA1mypNspUM2rcckzAK
3ASZQ6j56UEp203VAekmwtV3/ZIKTlZarGtqevkfFt7WJdQCInHwXXFFwcQUlTAa
G2lgxCvoYtf+ehQLilsitqhG6NqjhYHr7LMWVI1UC8VQjp+shQm8YQ18qV0Q3H7V
Vv2Zo0xhkwxA5+ID7+PI6pO1RRXpoBYSY/yA7xfLpVB89QB71rpGXgfG2DIGjZmH
L0FZo42/TF6iakTFtilKLcQ5zW81tS5guctnygGpzeDzUD0HP5SjjZIWehzyXM3X
zk05Fy1VwSZ2MLL7reK/bmnnycOIFfAePUFXfYazn8UgxursrWmIzRJyERvhpoxP
uL9h2TqN00xa7WpZkqAUiMO55kEaEBayi5Z0RFJvgtcuCzd15sUeUivhPjV7YhVr
063TgGwMS/M2wIZhbFZsNSE9pukU/zoQ4m6zO9lSjki1Mgo4IpQAkwGh6SAet6QF
BwsDYG8SPqKCMB7qJYaRHDwPIUZKGJpnv//lClzv4na+3Ro0eepf/ekO93FYI+Xc
VKx+CkM018r5vaRVUrhmQoo4UD5/JxE2p3ZsnA6YUfVTR8v1Vn5rmreBSl4yPFMO
tfhgEhgU+Fr6kjibtfH8KPnKIk8I4w8Sgw1Q4fK0FAg0QADNFtYqtHFyCg2Jq7MF
DEHfGgfP/fMOqldsbiwLWhxt+jf2kRzy3fk9yB+ovMafcBSjg4X2MVDxmKLjWcDE
G89R9vBX3QwbQli2UAVmuvf8OKzEOZzC2T351xm+LTdxT7jR8XnBBIUMPPMguurF
7y33D2p0GifeoWz9aNxhfewr5A9cHBbeJmxnsb2B09YLOqPNSPotYhizUVVShznN
SBBLWjAt4V3+/24J/cakUPUxV2xhEGYTS7kY8N2ShaxmXm2MwKC5jpqJ5hs/FAQb
gKcm+091jqb60Op3gJYhCHcozNT9DxVCAwc3VxzTJCXsq+qZgT903lxgqLVJyBzv
Tm7VCPBFgOEHqYsQ9iFbsi+DLu7W4nLpe7DKgzf5PMqJUbcHTuQLb+DiSW95gpWm
M5i9uHgXYUk6xi81zM1Zei+WrKLddbRKHjsCl8IwB7JB8O5aU8Ld9HPUM9EyrYuE
LPrydPZtUw3XMog4TEGVcleHY6WTmL9txsY2VM50O+LrLF8rP3CY9TxoL5axjgkd
sGxNv1+8SAW8rbLK1mBojadydws/YdlmoPd22VaTXEj1B7OSP3uBdbTAjfR9AyEY
FqFZsm6UGFOCuG9IW/jw98xWx5/4C+27zF91fcmH+12LG56oZaeTt+G9taMC4mKC
Ki5J6EsGyIHxAPaybH3rVcpfg9GYgHKYdvZLw+euJHg50K8q2cO506vio94Upsey
bP1SGqaEuAccTMM8JAh+4xmPPDB8JSj/iwxuhoMHlF5Or4UmmYhR7+LZjBmIa4vM
Pn/EMIbWkRgfmwQ/2JNNg6CMYUqHUg39UIbYxr8gJ9Ke1wMoP0RVqcsYLPA6a6hx
wIwrohALHxfIFIU89hRv2yBKphexjrdU50tMJIIcWsLlvcbGm7TWBuH6xNRSCHQH
hLQFID5dAIuW5Z6suwRfmPAOd2v3MfRhrg40saJtogQVl9yLCZeNqWLhEKcL5skV
wBCjl0XlUd4cFmd4kUBZUdiNNwkAXiSPNf5dH+QT6gb/EoEowNkok6HMb5ZUzxor
swKEC7d3WpZsJO1Sbf7Ycarkg6TgzK2igfJMdUJnThS6xYLmt2pdnkyn0OGbhrW4
rAY3U9HaomexXVewofitaaUmJMx3e1pM7VwUmvk8cnXcCz6QUPvFe7cz3ZrmQ+gC
6mHjsOr6u3Tsg7tBT56c0DLmoQj0tQC00X/dGpQ+prXcMXzhqRktawAh4J1SqJPB
nknvzSkHtAQRvHs0CrEhsq+9QVfxene6WtdyXFsna9Bbu9Rum/7KnyQ3PnDvfgfZ
oSGaYGd8e1thVlxHOKJUYSY/9Msxy+qn2S7kRqE9mosCjUKEUlq8GLmh+7VEl65G
lFY8jupvwczgx6LRO8Z9Vtf6TAYJph+qzUUrg5WHTxVHnnG6pv8H5bFdPouV1x3D
5Xwr5T0AavNcSU77yxkwMRIjORB3w1NVCHgt+WFz65R98gIs1+XVySlDVr6TfrAE
0zNJLw5ebvN8/JjZi4W4Pz2+y+P6t1iUyCxQYnJZspOAXdF0ldczrucJJ81a/R6S
KcsSweyGuxWz7PhEfuahzijFV9ciKkkza7nzeXw/Qy+MFHP0DJ020HONg16xr/UF
hwMRQCBHittbV0sKYsQka+vJgjqdjw11Vnv0j7uhbX/ffEOPzYhoYUO2gEzbiZRK
5XNFy21jzwWLWZQt4keF1HkZ2mB26czdkUmFEodjEJNG5ut4ASsqMNIo8qTvihFt
Tbp898HGkRSRP9L4CfOT+W0rwTxtEfFLNW6KLs9xBD/DPkd7d0PelI1yVXo7B4wf
inAmUQShcZ1RllPVR7+nPqERXKhdlx3pbmwa5z/htQ911Q/e2jyRBCyiskHw4Cn+
GstBvpKw86WZS3tJY/QBAoBdAxIP7w/sRpKxvbn/uj4X4vIrS+Rlxsgv6YPiASA8
8ES92wAeUMgLH8tk7qRSVTHmb+haLOgMjikpMFPQYmm3tfCzebVl+IQttizp1808
MVKRHYpG6FlmG+JcPAVmuFpBwqaco3HLmPAaBEtuev4It/kKSeDtJTTon3iKAXs7
iPHYEeVmUtEN44/ZfEYZhb3tBD/LvUoI5RdPY9EDueO3SBp9f8sKg0Gns4Xpb2Vn
tboGg/T8k7uiidtDONFi0cPRMlM6IlBRM5QDuE+/KnHN+cMFKXAJ5zC4WyaOpn6E
bwp2giPhVd3YKcdNsdsIMKgklRM4K3FJ5cVCKBPEOZGRZ0ThFwn1gI2Dyi6htDv/
Gt2SsULKNpcAbJwBr4SL2YyXu7XS9aBtk/X1YDmZjKtW87tZ89CAkFA6+JYj3+gS
ceixNMIB4rM47ix0tD8VKY5VHWAuOf2zTAOZxTLVGuDS5FUfYXqyY8vU1eEKgtrR
XN8+9GHzP5HDdLum2zXkfg7gY9eHlL2bzsDMG+kyxNOyafMnxcrJNV6hfgokeTIl
Xxck02NBopzzW7+rTIXMAlY2GEayYyStXrgYN2CYELEaD8xGL0QALkHhmRlQ52Cs
LyuVCWWa200X2qlDhzZb01U0K+hLww/C1O4ezLS5EZTeH6Dh/xAMWessD5E0uq8i
5po1IqbETd49orU8I5UVL5t0AX4UbeBtg2x17kUHTPLW14qdxNvpfyL+8P9m/2od
SLLFSCafnXF5Rw1Oujb5p08Aa4jfV++4usPRR7RnHtbHhQqEZhGM4sflAycGYYVS
h3OK8XedMicYp2LNEYHPVSAqvJwlzhd5+mHYwM0wik44cJ6XJvrQUD6OpeyvvDqx
RjoDKGC3iiOX89X7eC7SUQQnzrcPrvl+nYzh43sRVKlW1jzcf0Ky84pveYOdEccT
/SZoeQLZVscnOTLclF+pPFuYSICUqH9YYuwwi6IFILd6FOfH/9eep4iQ7va//XkE
8LJ2ZRNptoouorWcrZlBqvckb64TuOaNQrqQ/Uq5GAEDCyTw9KKL3rwLKvQWycYo
uxgcGNDAwTo4khr7RdHd0yjaeTlQnxu7DfzEnva809ZcU08inoMcNb3cVOyAojQk
sCYsXte5/nIBTi/XQeE2YKChOy1+WWCsJvWDxWfpzt2Hh5wZ5Wf21DGhpki706Os
xKBs7GCkRM4ESSRBQ5ESI3Sof8Iw/OWWwwIWn058z1O0K4M/RKGvPH0UV1m9IH56
c5DaGJgApJhNirGl5JH/R32R1otuKxt8v1yuAj/j1w32Ywh609/b6100ZSdyErA4
GyJWe6+C5Ye1O35kRGU7B7P/kftArlGKAG5r5V9nV+dek6C9aLlCUkllX7nAyWsh
WRyd4UFlWV8+JA4u2l2qzY4DRyP1lIs9pxhC20BP5Ph33ivnuZLqTbd7boQptgcz
Y1+xCyhkWEvcpNH/xM0Y3cyVjG8f7zHmINi+E6GVk6UZxmRQWWavvwRq3sOlbzID
jp0e48o/TahnvH/mf4uawXW9RsqEaAWvNgTRKssstoL/JS+MMipn+Z0sQGeslHPC
TYUw3BIR62WEXNqI9+sJi94cEWeR7FYrMOrhaQAvzK+71xl6qnkKUTKumw3AbkXk
hwOzpiQo4J24iHYpTI6uK5A/CGgsKVeUi/Oqv6PA0nEMOD/BXNt/8zARsW0YhZrR
Nv/FsMfciIKnvEv1Hsuc5bofnxEAPFfcgOi+P0oqBi110o41GJwJcf+uX1ka7j0z
NX2rUebm4NSmCqw2xE/JKb8DlbivU+aZYEMfHaTC93Y7Eh4CQedDUxbAIccjSt/1
zn/PHB2TWG6zjgNQsQZ5eEGk1eqtf2AvTRyiNBGkSVowONDQ3+32XNFbpodoSC2T
PZ62S6/V7Gk8oL9PzEHmhoaCwOUYdSq8KbZfYY1D8ZC9F0QafPcTeEdYJY5wh/yV
JZpBjIn68o4qWCWN/wc79Kii7HqGmqlTSNJulURV9OIkeZgTgxAv870d7tjqvHuP
/lSfjnfY9J6gfNsGcs16I5cdu94+QiPzf07Z2kq3NMTlq1hZFTqYlg/zgRejjF2X
+M+mlmiy0fyrKC68bosok3uiiplMtksacrqz/ca5Uiyp2uvgb3Aku9wTX9XrjsA5
peqOdRX7cnIcmv9QKMB/N9vVwZYZVRKQgwySy5168CirpIFXVVoX6cpQuaVzG8Nu
FITe2TdqJQajuFKjj27BOkqIgeEz+Ti0h5rddhB5urFOJh0PAJhBbo7X7Qdi5EC2
kfQsPlGKirLUQY4rIRDPDRngQ51EwJbfs+sMOOcYZP4j63IZSo2tYAbCH2GTdI1c
ZFoFfPzsbux8L0gQMzQscgAgRibdEOsEV5ivNtI02vVUhKVkf9nT6CwZVfHEZ4XT
xpGjCEFAtaNBiODFeqapVEWxnuHjwEgH1iX4WcwxElln7pTbPNkDhKIjVSGXwFe2
ZdOUFcA/5O0a2G3iFTPacFYcBlb9OlsjYxRAMGyMyzvwTS0FaASYP93wDKR8YjcO
SasDfzkpoZTN7BdXhm4piHUpbNxdmxfPl4uZN3kW34ICt4bcB8N6oHnwAFHMWyCb
f7q+JoGqURfZBwtZlKeYNpVE3PmMwSqsFgd4LdbnrwDzILmwEb4RFssF8lHD+p04
2nCDRLRKjMTCUDDKf4v7au3oF8wTaeditnLE8utFKHa0np03umYn2dOm4JqKup3P
6AfoRJUjWGld/wkFBpTL4a3onwnAXib57JMBuKOIrvfnXQ74ik8ePMRsBcXnzTSz
O/Kehw/pNfHtjx2pLsm8lCYn7fJ4pkqPyvIcJb35nwi1EtFICEjFTCiWxCZsmNdC
uHsjrf4Meaf49VcNXoGIM/Mx0nNzs+nCp3WQVAZ7csJsxuLWVm+gG/OSu63U0MOd
lvcX+k8Q/yBaFWIvR6NT7urzI7LN2GUxQO9mQBwTO5IRS0vL+BkQzRFySXBlKiOj
Lnjahi/DDukCnDm9/ot0AZBQEAAhS6sRVM54tvtGG+wiKOzsxT6V1JgvKYM0jAfu
QpgboaE9qJtOjo4ogCq7wQRabm9BG5/HJ0pjWfuv1FaatVff/k6ox3WyotDqqaVY
DkF1SU/rrEGyv2ODmanKd61Tk4BmW9ZkFbGMAUxB8uZYV3nA14Vy2Jz0tLU/bN4J
+fH9/4b6ltXuCUkce8MlmfPW6Z4e01vl0uPsGT3zDbEZthf/WSSr1Hrw/kpW6cDn
GfRDudm274s4lLzyPhAzTo30IAgdfJfIx/kVzu0QXgHWwW25rPf6SF1rNEzM86h9
j479PGi3brYne1dB5qLZD+38PWKypBmmHnILpfG/Pj0a6jrb+v2k6SCmbPT/sQ+p
irNaeoqFjCJkLJQlVjXuUYb60fQyBHJqmSgi5l11t9GhKAEpIM7oiq7ZdcZmtn9L
+pKbt0Y2kjXedRyfzIHbNcNxFYzrUjqPjCUjgYuBQbW0F1uoghj2i/jBavAa98Pa
nXYyJiLUWuWEQqj7s4z2GIVnt+9/XrLcNkRFOSMSzfiLAQwYbxsBeIwwckpmmmCn
EjJg0n2IBBBYCqfOOs2Lkw+qm7redJlsGFsqzqNnOIYFpmSBYl0kC3BGhydT/y8u
J3JOPWkSMABxHztqzb5Jfr95BxW2aH0WCZBTuUEOcvzg3LiURFzKIRPrcKqYyfvs
VCD6vzpR38nQhaODJdbhA28u7ND3wEF8bsVGSEHVqPbcNor22+0WKx1UUEzkTnxG
oY6h2tD211/WIP0YoGdRbvTr6pqQpLiKRxB0+ar4ltNeZTed0EdgJatwQzcPeMi1
ZJhcec5eYwl5BT+UbSLkJJjYCxlQXeoc0hHfhqC8mSZ7c6YQVb+OIJBqEpeQ2OAN
U/CJxMOf5SddRXBI6tZItD1nC3yd/PT22sogyDOzLWWmEWQpR/HhRM4+GPYMjZe6
+OWg+xOtmHgrh4u4izrRclmbtaFjUDUAdBO8ALsqPBqerL5W6aIzkrPoFuy5TIEV
it83gY4zJ+LVzIH9gSCHpgBSjxjq5Cgcqdo+P8nomFTarPSdAZ0x2nCVkR9rw+qN
cdvsUGTgfpAEizj9kOWYobONiPNMmEeiDdNI2064yJT0bKJANMGPQYZTzjteYche
O/dpzCIC3GnBDC9lo5MMsUn0HA4MwQQlQSGOLa/RoSQl59Xo+EeReXEcLgUckdFF
6HNnvDuq9ZOYtAHJf2zBQwmRPAHjAiMi+yotvTi+4TZ9m22eEVQDsk8xo8Fg5vNs
jHECtxAmoLu+6qn0GZ5KfU3j7WWnXtS+TxOwxc3FC9SpF8F84IOfPVHTTEbPu2v5
WgHAdrTBv4/O6QcIO3onyIr9muASHMcJUkPChmfJ++iKDuzKPOiCVZ5eus+QWDMj
HJWaXn90MgeJg3RYD3Q6YfwISQQPV96bSEEOZlLFY8xMZm0sCkQGugEtgZc6H0D5
o8xd0aSLlJvDXGws2P3tL20LomIu/g258n7iLc6vXgEyGWQvRB5MFLIez6v0dwm2
J468Vwe3FKkMvpXpTFXiou58eCLPIEnYcm7hJStyEiH9DqWw+TnJ5Uh0dQPumkGf
U3td3FON26RTSGbohvkvZzU/O7U5UO7hxYsCmFDayVZ++NLN2VYuhrpqZcUzYhB3
+3tV4TRDfKkVzrlYZbdC98GQwSBxQ+Na44N4pd/h4heqf4ZkjtJy6x/XXJLeEMOx
asRHX7oKem0SLuMUkyaTQDv+QQ0pO+ZNj4eU+01nJOf5yTYRii0qycl396m3c1e9
NTWQS976KnnVycoiSOboJ3DxzDP2XabZjh3CdfsGc871fgjquw8zrgGOqiLWIkJ/
FjSWMn92eARohmg6CBJwkOhf0GT2x4dQI/U68qUyYQ/ws8SsDyjz1kv6XSU+XAvf
e2tqJTtoe+6B8S2JuHz98UUUHAEsMNU79kOu6mBi47dqN/wHxQg3m8rBjWBHJfQW
O8sofYxJJAMEzRURSNFzeG3YRTu3s3H5ryPbz6p1ygUuxFsUc0nQ3BrbsL6+RrGi
dwrJcFuxvg1PN6MSgzXBm2Mr8FGWKsffeqXXJA4pwDHDi2JQoxUreWzmGPzhJYOJ
rXv0hbvje3HnL92NDcbM2qPKb2MPfuZXGtkC/rZv/AnkQ3NObB18TgnQ7yEDD9UO
X0VDu5fy5u3wsADuRXKojWAyWA7MAtJJAGMQug5jauNPVEX/jUVhFDBbSQu8tiJu
8J1Lk0blIk0guz9lrOoGYJDhb9r22Iu/AAvKQO1la/VoczxzjfAPK6sdPC7FA2P4
iba3L7bhYTRDyhppDtnKXBMkUkU91pxyQCOoCG+gYMtMDCBGkWzc5ZyCjNCKuRaY
ed8KuchT5KQv4LOD0xQcDozoGvP0uVMpqscFZmtRS4rSHPrTJ23lGFZd9PucY/A5
PFj8pqBBWEdg5e/QXQunaLH61FSISmeeGImuOHQB3tFJIdvEtBxVeWG3sQlxZxVW
6oGaoCtt+D8TlFrYLw7Xer3K3+h35Fa5tAI5hCkYJH1xDe8pd6ToMKealwqIx36F
AIs5GjDJRO6IJgraTycMeX7hFNTEF6QhWIxaOgir1ZnvGYaJaz7x37MGdB+QwIrz
TPJ3B2r9dcWrzu3SNIgSfNriR2KEDzlojt0NUHRHM1G8reE0Fz3xK6OwhNMh0X2a
Yn4uVHaqQCvIPUXttYRmswzbP2Aj4U3N/7jG6a4SWSrucLh4QACOzKgzRNrnGJny
ZdVcBmkQlyXMoyqQmOjfJuqNLAaRI/x8g4jwehuLxTr+1ehQfL4KKWrjw/VCksBr
za/h+6G4qjg9hrnQESRvGp21uyyuPMGhQYhxrh1S4Mk3NsIOF0Kz478e4oakbaSa
caL9+a7Jc35qXm78rKs8pLmDcu//PKCkRId0JYS+i3o8a0U5L7qEaPArCajgh/Gr
KJ/TcXUnjoPC22qnNtda8qIC3pjfPudFtyF/IUmiS2nmdhpKrVBKv2KU3nLKgSMn
qu/IhjTasYcwDirqgHgepGQRRbLXr8TBSrkJyDbYCpT7ZCqAsH1tT9YEoRw40Ik6
ueIlXUsA+IMB5uyFjrQ3p1xgDxl2kFjhSqk/wFi8r4qmkpJKB1Z/pVLoxnfnJfOI
u7QDnHTJFkfNsHu6x9lchKO9oie3TuqcTAqP4o2gjD3vwcpxzDWCC9BvJilu6yn6
JzdAHgFbFQGGO8jrbGg/m/MvymqNwn+6Bb8mfIWuw79b/bjF5hF75qYyw5AVktin
z6EllGOB6dO17u4OoS6SIrw90kdBI9x0yIu9rIST0POz53NQIZ+af8l4ERPuxrSd
7gbscNDfs0YyIOpI0n/gXDTsNgNnsJynnZaYBwywDOyojtsgU5oG1n639e9cdrqG
aJV7BoiXgyoxZd+j9s6RcsudR25z04pd6l+54I5TpZ+fX7bOt9UYYWKhT0NvtJgj
EXu/QPEIEQuk66NS3Z1gwKD6FOWbzsLzOxGpVeyszV1K2u92Z0Zv+CayVW3OTkiJ
G62OvdfuCkparhrLb2IZUpOqSRd7BZCOghBkDc/DyMoKYRHGRJ++r5MX6SGNU8a8
d5SvPVkLEs0To2BPDksiDd/Gau4vPpo0tXsqRPA6drnWNBJ/GqBAiOHjL6AGuzxd
VZXktgK2vTOlp92CDszRR+N0dN63KmjeECxiEEiAuf6qJkMqVLd8XMWmNS60VPxX
Eoq0U8toh/gvpDMjkjm9gkoJchP3NndlrPfOmLqcgwJmQ1hwe7LAh+Lbdy7MjBZ5
lW933NDs/6ttg3YoWY0pVjBlgOYj8VAujniTwASAwSOFL35Nw651f+9wsPfmlegu
nEsxTD75Hx04FOq+J2YM99h3oUJSmXPLJkQrgkj/HqWxVjOjPMBXuYiSBQO4XFUv
GCU7ddv2NbgCI9WWPb5iU4/P628rqZc/szBv+bGBiYcGZD/t8PGM29EEOAJLPUeQ
bMi1QQ1Z38Fcbcyd5znwfHwrXQFVkbBQbdjYT8eVXfyF2+6T5Z3hk81E7e23NSFx
4oH3+wqrEBFLzEBAtUANk1AEi/ytCFG4YG023zhSOn+AAhJAeKMnbyQy0qe/gmFd
h4+ajqk9Tl1AGHI78UJYEnHIFSpZYnsQKVu149v3WEhLYybdzz28CSvzg1iKBWBt
kLWFVeGgo53rHEaLRPK1W2f2yHjcVXA08Iwl/cwFeuVcww9zzW6dh4pOPJEOwqgv
6lBEkgoAtpwXqy5erMxJbPuLhuRREgxl+5uiMir6Qsv4eaurPGBIEfjXvMqiMEnr
CBxe3RHM3uxnSb3GMk2SA1QCizP6uGK3LkyhttFytpDACQkCV/Euen8/Kq9/B22S
mcdZJjgTej3UjQDv6HIN6mRudLmumd3l15O5GNrfrgIJ+1Zetjdk20F+pTcMxG3s
4HoC5+uKqW6RyDB9Azdem0CLB1i+9WIQK0IwFe/kItKEFg9Jdg6S2jh1IrdlVdDt
he2si5bnWGtURy/egZdzYF1uGtdkki2LuCvVgxp82mbmsJ1FBl1exUpV34SFa1rI
L0U16m1WsiP4d5/zULM3DRJ12SkcVAlpxPZ/nJhmDbFHnU6bV5A1h9xfbs3KyJjx
/yYbisa7ZvoYqzz9rfgsdBFnCcuLzn09AKnlQ420LpsuOLgEAcfnkit6OlSIrr+j
oN0NuR96wEBTMYOp8jT1aM2jNMfUZGZiyJvfocBJWNFjIXajgGd74PiNtUCgNqkm
ncijPIA6jMpQzEwEsojrF868+9Xk5G/M6a2oGeW0zzTR3GqTBBI5RicK77xbD2lY
3pOLK/GLgkQlS5iW8HrFtRAr8EOFJmVUdLV1kfdN8ccUb3vXnrS1u9MMhkxv6xmw
u5+vfXJV6azGwotMBnDvTkIcHS9uoipph9HSJzhIfKJXEOQhTFfSZOjq7HevC96z
HnwbcoN11w9RzS70+Mc0iAPj58PRCJVk6Eeg+4md1sEDCNb63oTY9Vboiu0/Z146
c4GwMgyO2pLcmG6wHtj7q9tFFd0gyvht2OzRb6CH0N0I610KWfv2gENXUddKwD+K
YjZ09eKcfowq1QEdosQ4HeoqlkBLVi8mY55ipYSXc0EkhGQTWtgtPm4aRgk4OMXy
t/k6VGAv+WZxqKYFDA2CS8AJ9pYu9f4+lse2R9GaMuocqyvvWMtDZneV+dCYvK73
3JXj7H2DOtu9syXAwekbHbOLwbIQ8j88lCsgO/wxNFdkjmrjXiBuL4UBXhS/5qXD
Tm65Rahmk0Co92mpcG+ZGcjKmPM1CTqDgvsCAj65HSERhTHaZMJXwYhZszj3ZKrO
KgPvz9cs9uv39TsldE8hHpxf1gfIDn3H0yUbXbHAEJ4A7dOvFRNgHwzo4nE7cCvi
mx1gLih83xjpGtct1MNVd86e24JNGwC3PbYgprP/1fpwJciaaBqaFI6c7/CaSxqH
JKmCBVeWhria9p63654uWS96QLjvzzmbFEpylY5z5mtwJ4CJ6RjD2eU5HlqucQvg
U8k8/dVufw9viX4nBv2GavlKST5aaD0hHKwNhC24SaoFjJ+axHHeN6RwoNuZc5X3
yGCojVUfFXm7aRUYKlmNkmk/xfbYwYpExzLWF7uG/TwzcUp/c5MbL1Vcalpe5TBA
dxJE1Rpi/fgRfpRn1W2jS7eF0oD1MCpqPeRMuEIu2IfrPvOeyRvqSMsN6arSBTMx
l8rSq9IHVcGWwUhFJR0OnbcgSSfx9y4bwfaZHaaSPsh4gfZS5fq5+sUvijSsUUCd
rzXp2kin04GA45gotGlrmex904UUOn11RfS4Lj/1pII1ZW4Tvnqgd8T5Vhn1GbVz
68ILlErUaW1wojCBGlxjngD8bQhua4z6uil+HbeEgfeyNmG6BQfPremS1A8992Fn
0CYdXEXKufxeNQn51pHA0FZlZ0gx+9gjOOnHZHl3cKCnZHmu8Lq6NFdEk1UQkpso
poT0+Fjo87HZ2G0kHwMpi++CAuocoXiNIz4kK7+OVL/3PwbwW+daVc+MnE5fCZ7b
etagmlvO/+Wm7064/N0u/a/F9Z9EbjtQZsuC350MXxtH5PwLA3BEAIgWIaBzJa9z
RD4Sa2hUm+dxuCo3ZKaoqxXzsi593eiKSZT1iVztgogo11zfh27JtlHVxS/jWIaK
CQNu8jEdikoFRwi9Vjb7wtmzl4nQHztYwLG94EcyI/1CLM1XhPpuTxSuUfsEWekJ
dBZJ05s+OY4EnOryp/1rBq8DxxF7nIk9xFuJ/jxfWSFeP8bjAi2GCvtBid2QJibe
WYSt3wCuNEubS04XTWmzymsE/gR6jqVVkhk2ABpEKXHUJobopj3LSIvlHEMDnCL/
2iqGWU1alyEhrGNxYZLTsWkeAr+bdN2xZQWeIqHMNS3E5Lf5qGoiLT82W1/yMa5N
BYbeUz+q2DolV8zV/7fE1CZXyIX7d2hcBzHzdGlQO3MSGJMhcy8l3rTHfbhsI27/
ulw3cFuDl0Jb3YproRRf/K5qepw7IOsxG0KF2yFPhWXk3Jc0tAEwTaBbb2V9UAPM
XqXU2eiBzfgogQ1/VV+NwV7QX+hORfntjb7rAH2gYy2Q6nhqneW7oeDPNHsyMDyg
ES08G67K/8iE7pQuIh8a0O+C3ZsRYD2myDZTUqp6y/qPpo+ujgQaUCgMoFua9/pv
nGO6R1mAH0zpMWPgUTMTMRfimvz8c84Al3a+JU+3rGXwjKDV6xTrK17KqnDuJZpM
iasRzy8WpqvYD/oOIpIZOe55KdiCLSAxgMctwY3pM4XWaRSDhwzb/QgyQWbHUBkq
Ol1sYb3V01qhzKAMFGfVYntOCNU2o3VjZMhDhoCoVohtFscDi5JXPHdC3kSRiQxo
kxmg1ZDKUZ7bF5OXQqqnTpR4ZSo3jDt8R3MplBQKHxw0t9gy8Vb5RBxYrOSSbugT
Z93U9Kio/cjDaB9omgc95/FI2xFuswxUH/c5SPvyHlaOiowh82L0mJRqXilDKjoj
vOjXAVzfF5ttkX26TkRkpOEPcb41z48CoTdbJGhJaCdrXqw7jO0lytn+4ejQuPmR
wnVZdPWRP3KLt/ZtbbABYvCCDcYU8+XGxrEeKbK5Fl2s73byUZiM/dIzPuXLBmtl
U1FU2UnOVoD+Kps9jC+zljkHO2lFTQ3p2WA7XVkB90hXu7OO2bZCtn2giVNqjp6t
naCknomNTuzd18/EFcyu6OdCeXpfwuHSTncPZh6HMZheFKh2IDkytnSqLTGlhiyL
d7M37xrIIyOZfrKs44c7HhOAUbCVvEUgKZ+RJ9IPjynN9qCeKPw6FBV7Kr3S1RpB
hkdDwqvLSeiMJAyWh1yKkIuNCp6nqpze6SAg1pzqCx8agCzk/g2TwncEqln4lqKw
OlX6GJsCWgz6+JI7jWso4K++87/7tpmO27NqPOT4nnzU8ts43xXqCv3Pf1p0lQFq
bEc2cRDTTxwfqXEFRSc3RLfFiN9l/S2M/gGhSqr9zashJPcnnNLFdXxRzP5KDNKB
TrPi1PnGo4u0ADZXijU+2CAFA42v5d7Rn09z4hzf8MG7j7InEkxskmPFrsFkz5UW
+ILPbXsuLE1HHAEltg98gQkK05j0SqxbQCy10/N0E4ihMraxlsgaxlEFrJ5x+6+o
m2PAdWmlbXSyyeC5qS6wEX5ThFQJXykjpKt12EqJZreOBjUxWSkVxA87dX7gSpqN
AKIVnxZCZeASFhAiBwZsRC+Q59j3AAuaO3YMDnBH1QZL0vSwk0pZr6n5eyTY37LG
gftT1fN5ve6l0HeufiTOicsIiylHLpqpwHzmq/JBWKGB9Q1WABZoERnms236Nssk
5rnHZpnOOcGCsGZQf/QhQDFPyiUM8plLuEK0QeOGzdS1KSmXT0vHIEQeYiVsnjEQ
lueakGUdeIb9IHu0ZR+P4EOEzDr1BnB1nA1n6KL4L6nFimzyFvBXJf6bOIH/K9ls
0sHn6kbB4Ygf6QQX60gewRcDPukKw77xebSnHKVsPlxQm6PZNmv2slp6t/KFieYo
vGa0RbKHHyOAIN5bNwlYgPQljwU34nKjsM3lseEvpFHOfirWrnHHi0MNf8ixZVgM
aKBOtHauNlLIX8VBSVZE7s7gj5C8VRxnvSNUg9RCE1KwH8lUKgT8Uv1QkcMmvmUy
HsPxftJM1HWmTlpNM6iwTUtKBByxwYOUo+AcZ7I0ToRvEdWkDi/3VKoNiJVjXz3W
M1jr//Qq1ggGqBUY0uWlxBkyaQcP/tHOZMvCoGIkAbtqnhAlp28zDumqayqBePo1
WngauGE/PNn3C4FfzTUKS8fp0FzjMA+2mLhmCN2tPAifPnNE0nXITTJC+yhp4yrV
sUYf3AZN7f9w/N0drFh09NLwW8e/4sUFW5X0MFY0HvM+WTDju+GaU7EWx5qoKe5h
ss8adLq87PLf/QXi67zxCbIf408IDe2cfqemKaNrdl16LzHBwo78/JR9RZHHt/L1
HvOOvaD7yNw5ZtKQmX5naWdMalQ9MsK9qLKhDCkytnoSMTiU4qxgP8a5wjfisb1H
A/aChOw89vG8n3fiuNloukqoMGyVdnx2LUGd8N7KgKVvgRUzCLs3vY8Csfb5dh3u
OtqRlkWVSKRhu/rUBCacgyDhcDr51pw1Noq8GKDa8rt9trMLp2QTiP5aM59xs3pd
vELiy12UpFHOIAFh0Qik71F0w6J5cPOvbbQTDZZq6RnuSbicBKzLNXeyb2DgISaC
vlOX6mmbBBJxf8hqcz15/lswIHCygmhXZS9vIsNnJug5ZkUbLkuZWVWgbYM0X+lm
UiEByJoarFeYbOSeocwF1Ij314pTVdcy5mpbRIhggwsO+HKJLPTVXSUd04ApFIBR
hAuKTnsD23AW9EXieoctzM/NbXC/IDtOghkVcKnyNkZ/kh7QuXW1yKHVxrvS7N+n
JL1kvdXjYOIzCnlNq47lZHGwI5dmQ0BmnIDTP60zX/qdYQwuxd8hXmo6m6y3rkui
YVbS0S15iIALcbmQv4FZopzuzS5w6lDhuZg3cQ1M4gr4vTwVPHtAagzskV6+cumG
NL8XmCb1cC+QB4l/GmSk3nyE+SWQqW5vRsBvXGZYMnlh5M7i4yel78gU3jO6z2yR
zZdl6Sw/YIrFyySwTRaxgBniBAaI0qRRIr/TjLttBfC7epv2bMjoTPJ4cez7M/Rd
Pyz6WOEl4RFaW750xmwpUnClkH4Ai6U9V/wqiQe5bwRZAsEXffQkp3oplwROmE7a
lE5hxfVU7VuYXzmVRYEBfvTJol5AsgCVRw5yz26UA+Pl+XlAUHVzAFkLK02gU9y/
CMoj42HgQpq1XHWJHWb4Gb+rZg1+AxfcKEv+QWdMMVYQ5A4Kq2KBERR1Cw+Gyfvs
PEpd5pj4+jDy5/yLbZtGj5mKyVsURgSq9roNeZggipNI4WytYSUNAAD9jA+ykyXg
TnFpY4IhT0ZTg4e7OZ0DxCrMzu8EkDGIvShkR7PqdRzRuF+gsjZd++dEbhAgYRcb
/UNhYP2uT/7/UQjoiCKHFaH4n84HPIExcYQbc3qHSuS4s+JiE7mA1xm4Uh7UexGx
kxO8L/y+G/B5xcxe+M+QFU/p6DyIIG09U+y+mhQk+/rvvroOYwa+bhn95Jdl0Kvv
104nCgbKGIiMRaDtl6AHgjzoz4VjVLxwSyKADtuQFXZAunj6JS8/sF10NkxF4Tcg
eGfrEDgIDR9WOKCmvfiBf3IbodoUDPXGwr5gG5kF+haK0+TWxE8llz/0WdFOTdr/
ASxRSVwOalu/LxEG0Z4v57DtUmF/Fszk0cOlJOYL1W7wYYh8tffhxOBQRyy6rQd7
uznpWufCFxFJeB+XY2RBvO7LyoClqZ5yd+LrZtceYX9u63DT+EMwsGjqNc0jK8d+
MNi0HVcVtN+uyJ0J8ol0UYm0LPuRAn558qidcTSvYWIeXa5rhQxjgSo/JU4uzFja
lKLx+SnkUjQ7GekL1Xs6WwbMj7MTLQwWKgtz7OVQeMPyMU7TmneeUxulRaTe4vk6
8RWNHVlpBK6mf6Cx1b9GtGv4wXZx8ClIZZraYxZuesiviLWJLJ3e05Y4T+koXeHR
AHasVYDAgwlGThuABlwAjCTOgpbrICEvGLTRltbRCpigSW0EksY1UtYG9Q0LktrE
WlRD+uK2FEBGZNutnSSmWNrlIUCemln+3p5AdcRDIL+SuGUYg7ZjVLIvjiEC09dO
RdjkS13gF7R7C3sDviERht7+N9cRO1TM6LntBy2sG7XtGAERUFeFhpJetLLep31l
uRjTOkgOFd58EsDe8GHDroMSQvz7IbUf1cxDmM6V6eb36P7uxl1fEU7GOzkhh38v
IwDMAi9O9ReO3/uCST00gXC9XTahQK5p5apMW5bFl5l33SPI9+EYlnQP532SkebH
LMU3lVzDt8ZGKOL1FySmYvRDfI+yjToY2VwyiRQ4IDzzBh4k29AoI07vH4NGR0eO
IF8ndkZkAjPlgbdl3Icgo+QndPRhSANv3Ak5I1RBIBU5myR1f7a/zrSLJM/nq6F3
IgFj8xxvKcycWJTteoCLYI1HbVcp+kKW1NmnVsn434ljY7LhIzk47miIqOaHDwiU
0zLeITqFLOu8/SLcM8pGiOxwKYRUU/yLNG5Lxa88Dbnu2xmFsrrb3jLCbLK4bgTs
MJMHL72KpSYr9ML2uT/W3PMoNBdmsvgdZRqgVx2qykcPM2TyJHQloYPCKZdwc9Km
9lPnBPbpB43rb4DiJKy0rDj4OBc7/hhnsXfqvzuiU1wZVy8l1WoBlR/jJfvw+bJo
CrpoLz9LnARcNRsLz7X9M7SzUT9EZPwb6KwTxw2TZ8M+wFRgvFWOfL7scGgf5pax
14mWHz5vNvu4GSwSaHSYhXFPuFN3L6PyFpMtcxGoSHqBzBHXkhx7uLjr43m0GMO0
zbhZfYqtj2i0I6/j4CoVSMMPRHXYZEq01qmbUzZlC7utfIsfO3LPvYKM6ehwtvtW
uhxUdIlNJVWgzzSnuagAwnsHC6cgqRHmv1bOVYE7czikXURXdXkla602hLLI/gJu
+PlpH3KupuDucY6iFwmFVzUXZPUtc/LeSggfYt/kMjR5cInija+9u9gAsz4K3/E7
aoCW1Blul6C2Y9DaWzboj1hOFopa4bmXTnQ72+j4KYhYNy4d7e2u2MQXgvWJbAeo
Kkw07xX62W6cqu3gpY8ljS8mfdYpXZZm1+FZugq0b9ErQiUR5tQi1lApPRkTSwDL
lRDHzx4u1NM5O6it1Yi2yM8ob8Hs9Ime+FU4uhiU/3YpZG2CtySfKfMvlIKf49dL
xRKJ5pqpeHyiipjgf0VhcgNTxSGMm2cup6NRq9kvT96VzCMNRuOOYtJm94w2nt1N
mGK1rdJRgs+d5VoEcHZ4K/CGPOpzDk0PzrwunMJm52jD1a+RTXMBPvQxHf+tvP5q
MRszQvh/4UYm09swXyMY2Z9RltIi9lgL5zPSbide0kuEjQd7A9bhDWxeeM5A9EuE
bpcRAf12BOCAI455HVDE2e4+/3Zpzu4TC8+qsvQfH2Y7BNNHfbm1TV8uuAeMws/m
D1ZDSe8i3pfqMxEK35g64FPBjq61GBg52IbS3bFu7VawVfkEwAaIvh2wXTjT/Xcm
woD8vY185cx3fPouGWq8MzM0J6kuR20JDmzwIrrn+9gqDb5jdYsCq6n9X0ci9OZj
Gsx6KOKlaBsDLZ0UVpETBVdpkPJ6Hf2kCTwgj62d6QA0UkyEg/tbLF2rH78IzHb7
OT8ocJPIdSvZmNC35am5rcuDAgvgEl8LTk6SCt368lEQIquQb69+O3l9Uau9DVJ7
14FhsAjAI7l7c/QkiC8YVfOKGQY0UIW1hsKPUvW2NTgliE/WKfJakJh9AAg94z0/
ayNsafLuGBxlIqR846XjwBO07+GHT+uZb8BDcPDi8l1P/ZEZhjOGfC6Hhtxhyb9A
cpDqXzs7FFyN1XXXLlmcCUS3whrrEe4URbRhETzscOYCQYd9ZOypgI4FoAaFXu23
HhzK+DNqDOVDcckheN9j68y98EGvh0vZTiaM0gpVfanuRktZgJHzJnbsAvvs8sQl
bBC3YWtEWmRC/kMHYY06FlO13LrBygRiZRFjIk/5+mEybwYvjOtbGSFtqW4AoL8J
uISxwW39k0R7iuruCBHrtT/2/oX6XcyaxqG1bJlRE42iwLV7fLaqT8qzrhCUUeax
qRx4IHFrlrwDoC/JGW9svMMzVgYrZ8BvsYaGmjBi0Xm2CvLjiAHWqgX1vR79mwbO
xhyvV1ozLIUxx4jIWdkSYVTfvBTwIykvhpn7d1Tt6ScsrP7HyY+WunZf7gb8cJx3
G9bev7ohQKvN6o/y/Ss4dXfnNNKzHSdR4decbZk8AB65j6EgmmGBn1hz2H71mLBc
ks1k/SbRe00qZpK5liTM5Ctc7xTDhH6TJ1KZ792GZXZBposfP7J+3uu28WX9W8ub
JCkvfGalgGBDU4LOfZLwFeuDXzYlkIvZCrNt8tpe0ClXyZqGlakr8AJXz5znNeEK
RepFox6mIC0WokNlf/iZG/BZBDi2iSxjE7tSQuj88tHxJ71d9U0JYwliaL/vRME4
HtPacV/FOwlIFLRvniVt+QP2F1VKmQZmnZOHzqqxyDKfiTHO8q3T6bgRenZZCGEG
NHSWJZ+E/MYcObQSEm3eba4F0nCnbZ3rC1mVV32yuZfYCsYMrVjzx3+Y5wC9UrjI
oI+DSl+XT3nRN55aRyGHHUI/NA1f9a++Kf1WIZeFgZI7ntsjfEQKvvPD8vl9VkY9
Go1CmEfrnDRcvwwLSFeFrLlxFyu9G46eW57oLJ7mmzja1ra4mDUhvtqy73tRHIJj
KgjV06+9dvm4VaFH3DPcw5V0uWDjIRpiYDxo5kDxdAGnx0w/hSw4HsCAgBnODNc2
BFSiHMGFG0SI8brr+U2o5qypBBit9gtPoHl7UjwzZSdtfadiSIk9zot4vO4lS6S0
J9L9L7TazVA7ipK0OfzQKT5WjB32d9S5rVV6XLn3yRxDBZqKSmZZiRsjb/0IHXoM
aE5/Hocf0EuWuGRb4Xls2N2HXM4Z2JynpX92C/uBjRPzGFli4eMEaAFyNX4RqSke
RAxKpGoT6Kb7Zxgw9OoUN/WwNVOelT7m+QGu5G2KTVnzxTW1XW7hKlKuJ4+Bidpy
mp1XPky//AbO8IdAbmxE2hqc3XTXIfS3yxVOY4j0cGnVoZuzbBF/4yxLts6Cfkad
oStb+JBkFUPzJRDx33kNU9VcjpIDxDyo6KhOTWZuSbCkox/ovleILPu7lBnh8pIw
R6adrSTuBxCmQbfu7UfUFolZgZhHYyQuOoyDzHBENTe4sKFC1FBh+8mcDeHpMyK0
wiStwZI0beII2Hfe8LCPY9YuZXXs5Ss5iNy+sAlH7mCeb7xHqfvvGF/zRsoi/H6m
rZdvwwfqi8oFVZQ0Jvx2DBH9+JQDgQyOuYy9WFQTrpH0W4LE+/Qn0CEruigh8FNV
UO4OC86YBBxaG7p3OQGSUTM+sRzB7bG/ght+758V3j6n0shjO8untMLjBrdtU2AO
LY22eAlVOPDHv4wR/BKc54v/VJ4VnLSSvAhPYqKTTzb8LokBObra+1FwBPr3Fl4S
705fvrssFjMDdWI2XxOQVB4DM4ndfEiCUpb+RvxyWTxo1RlrqX8qnqyb4Z1XLwwv
QYBEy+ps3qMZfMTKbL7mC0sUYgDp7DY6kDl795TGEu9PVVpa08evG+hzlPKwLFyI
/6NxOUU+0kgTbCCke95DBNcmwNgiRlO/nIe2Jlhnv2Pw9XZy8w+avg4wllAOrSv+
dvoOjVIb3TNVIgAqCKzLklhyTZ6JzI7YAAwS/4FW9YzWTniRwcyPeESHeWPqHL0w
GgzHm5LBko39ylnMcKAPyHXM4YD0lGLk22W1ZjKNYr7FpHFMHkGF5qmdW3vB2Vsp
YhWXl1fQ9eRzih6mZ3MkCih3GyQRt3eflv6yGbQZcNVMjckxEBcJi3jwjrU4Icp0
owGzLvftIO1f+zF0Ly67rHhn980ek8Kwb+riaGe+/EXD5QtCGxFjH2GuLkphnwIw
79xLIvppkIaDQzogfbud0QubyXiEhoOJUEjg6CSx12eQa8HtBQFMLm7RoOP+RMzt
69JjTWq1kHfRswzFy0h0F9Qq2ck/QBGJCdkz2YwUoATLYyjjD1+UeVhLjco4Xs5b
f5I4aRFZ6d1FiZJwhYhEj/Oe7xGbc7GYZW7gNb3SaUdZUtKVDO7AJJMQnyYWJ6Re
UfsqV6ADOlM/TkkxJihn0C/+PbplLvzNj8ZnKA7pS+3gJWIHHzTfyCl9IS3oo05P
II7sIMEKoysFjEUZopemdGGA7Fxcv4GOOKt0i6ocrUz4a87PQiIs3lEFebvP1VR1
94AEY06Q8odxb6eDCa1m5bG5S05pkuvPh0bX2z82J5DmUUNWxccBvrzAkC9YG/hV
3nayAenoqyWwCzNN278QL3NyYqxO1/zXeNeUnT7lpO+47dEVrR6btV/3MYJ1zCI8
RLLM2GFObHIaC880WkcfPP1l/wq7eMYmJu9VBzG1yWYHx5Dj7Mikyeanj4rLUwqs
ZzyXvrSG8nIM7ilGVoo5jC3NXrQzKFhvpAslUgswjK09195jne3BkW1KrDBhfhfj
6V3tGh7g1ORBuf6sXb8xCwH9xpEAWfF6MyYrgTwAVUqJP3XfFs7q6xbfPz9KDkmV
Z/A9DEaLV5Lno5G92vLvjx9BSKj2NwYaOsWHLkmU4ObJzfcMKSczMZJjkZ08cMRR
ZlGvGYOKVQxOma6HI5OH0rARlPznkSFuMdtEiX2/QFGOVwLJ9PGXwk7s2ACfwc5a
8sVgQ9rdLKSu3qSaO+z1A5lcVpfzOK98vqjSI7NQoo6/SfwQ6g+0y6ofV15g3D7C
JVo/66N6AkiNYjvXND3dRw/wDdkfBNXL5nj/SocZxvLtmpysFUOiuqSgUkGYksTQ
8GIj/5PR5xjHzdmaN8krWy1rMcu9zU3xs/O1DeAc1Cd30bR2anbMFm7pL4jzPRIs
p0JSSLe3XvvxJP6SaCFKgYAjtToD1yfZdutjc9xOedLMS6Y1Oylycnu9hhw45lq7
7sawKCDX3WBWuVjMj8rH+r/jveblcuFzQ7bhk8AJlz3wch3zRtQbPOaFDL/oxXqA
ql6iiQgQTNcrruS706b1smFLcL6B8C2BnFvey9UeXjzkMsB/mYpJ1u4sGnqpATNE
IS7iwpn81HwfpCzWiHelF7bhGH7DzCYGAzpXVkQWB8a5JWjRgm9pgoKfD7CSkpMi
bHVcK4p8fBQwG/4YOMM0hgL7XUlc7lp+upOwGgsy9EFNukk+mD2Yza+zcQoIcAOh
dxNTF1+2GEaIwhYPw2MhpaYnNbu+EJU4ww0JuhfJ2I9KhtL9xgL8CvYKhgxpeHvt
oCGNkWw0hZWFe5pKh+NZ8f6LoYs4fy4r80mnDLWocyu6+jWsDjLtOXoIwwZczHQr
JYds0ALSmyui8jD3SYGP1fu4Te0ktJtfF2wqot+tnY9p4pw7VWvSTiP7hzh4Bygo
MaedjHFgJedN6GMxTSt33GRwD2LvFupWAgWLMG+FQrhQjL9PJCduyfUH7ku2Dk5n
qXAeHubwup8SHYYdSIzhS2lWpL3mjrbrPqyjxQocbj/PeJX5RNk244nAyfcYIelL
r29WG3Vfm0H+LEv1jRefQmVlHeMzNz7/xgQ7UwywAYPrh7PD+iGeZtnAjHsRXxBg
+NvyzHCvb8R6UJ714QqauiRA0hS5m52Y8K0GOPO9+L7/q42l1M2pXezt7L/7UG5t
vb0vp87raId4obBmThB4mqSfUxQ/gbLmYo229uZ0aOVqvYGTarmpyFvhMBlRm1DL
oB/Xptj1xbM+jd7/idLr23cm21YWscHX8iQP/ymN7K4gCyRWCRS+w563mgEbI7LS
1o1XuHPn9liXiDbUPSJ6/v/qUr7ukmq8e6Xrt6bdlyH/9R7jO1Y1NCZpOXIg3KyB
ml+7sO86GIwa97AYxlAr45Oymu+2WBPI/uGCwaljIa36v1uNBDxu8z9T89mJfzIE
GMQIPJaPYAfDjSFcysM/h//Cuun+fOqlDqSQHarIUPCtxWEsmE2f8mN7yNaskNsa
Lg2f06KrvSgRGdzO+wIX/Z3IE1W4U1SyoiWqJw52EnkEFRhsQJY0S9A7TnanVpwK
ABuJR1EK3AQu0QcGu2h1yQoYLmL9SKpNJTayNFFHGFQ+LtZMofwWcpKfwt1AOrT5
3qCuJ0qDe7CxgxCyGwje72NtACtvQGXReYs/HPahMQQUdBm6gUtnthLfPp9gIHdA
XRrY1OfDTs0yIHdsir+5b1/eFy94Q2gkQsuX2uxjGcvQZtPz3Cl04PLkerOWphuZ
c78ovIPbYnANaDErMyazdiOOjIIn6EwLWDVH6iitFE/AT6uo2dJ+ilngCN0qmf4V
tUYgnSShrFoO5I9ibq3nstMXQHuodd8TMa+FeqTXWMFOvFy8K9uEgdSkJM9NMWXa
aXBRcsiS1OlgavJf22q6bUBF+5SLjVKbN2qpZT8nwHH7tLQbN1b0PXKsJMQXG5XW
KygYISfAlT4JE0TU0uaJQ5T3rvX0v5pxBoPGEHNv5vTOgEMzoNXw5WIGYWyXx/Ql
rvZWExNH3QSZ5ECcre4XXk/nq3xmYNR+nGukzq9FkMIJUFZUUOxKMvAHIq5Dim8T
sYoEsLinaWopIdueEWCum9Zvhm7yjAJfDGi+QHjtnQGj/o84xGYS5uX3MisbwBmM
BkCoCoLoq9ea4xUZv8Hlpi44jkKQUWEtbBdXeueILkEoOwycu11ZL3n9mxt6vLtw
e6wtd/Fbq81iYGoboBcCBPiu8yLreYwlXjAAdAw6isY96p8IKNsSVSTB6PwQ3RsL
jPEtCpN1Cmkz/X8705t9ragUETPfs381b9iW6b7vxmNwvDgiDeiu42WqQSM/jzrB
QzScnvHaLNTefoSSmCMqusNqFkvCW61GzV5J7ii9iclRDITYSKetaPWFaGY6fH8b
6wPRTRMFSP1qICYHpm8IX+qb8a4trsT6aW0m5JiVt3GE4SgNuP7Hc9e6MaYDUP7u
E7KQkWKzBg5wHAomth7aa/cuIEFUsfGTqAy0LilbdJHllGSRPF+Yi6GBNRZjk1Wo
Qga39qBJemOlWTJlo5rcikGkmhfu63qufO9VlKljFuUwLLPR62j52siXpLrJs4CW
wnFBL6kVk3y4oF3LijM4vry/tkShD4WaHYJ0NzVrImHwI44hP2JuYQihMAQyebbI
E2v1Q0fZaWL91EtNqS18ExQYclgPpheY0Wh/gDtv1TWoDwsJVracxjD34WraZSVW
nZr1f1+AJ1AoWdpWtWJzfz0mhaz+EiEYcTkhIGwl6Y5VlliK5kRNaClDi/yznEgW
Lsv3yf62ZBcBaJqGL6/FA4Cd9bUSbS6V0hw+9c54eneSPA33iZFy+SfasP48RGt2
OwTkNJudLsBaIhxatNtENYqLMB+cLPo3TwBn+thh0mt++4km6x9ATEF8W0y3gjft
T3c1goiy+gKZ/+ff55PX2oNrRx6tAGHRf9zfpURGbRTwyD6/qusATmx0yiJuG7AI
65vSjbDBF7XoDOJop+gQJ1+D4lx8mmD4an3OdquSxR3z5G2tkTeEEkR9FNUpNFn/
ogZ1MbH+3kcetGhr4MOj5vlpDcOUAItEcnyDFxbKGVL8nHVJ6YYxsS+dUQZG7pjD
4cDpdBU8H/o67lVVJOK5lFR5aFAKvJcrzB4ohHHRbTKGxnQ4y0ooHKHC1ldJa3hO
Jkk8A5UDBtsnF9nX7oK7uGV80Rbz8TEBeqDPzxVJ7Mzu5hTcm+L7Hm/coZ05TEgR
ISNHhzfcb/JSMW2OMDLQh5A/4K+tU+mvaCrxtJ77fd2ng4H/r1qZkYood0bNDlEI
yqTdEsFfzhjHSYauMqXDg846znfbnM44nikl0EOlUyq21gk7fhMc5K5B+jf57coy
ozFOu53O7qtUF7cGX7yjw0MxIvOrFGRrO/kA+OVJ7VJoXhsL/GAIac0AIDnuRH9J
1+yR6Ml+zTFJsBqYYmW25NBhlWuiM1KrmKTIKOn0oE4MRo/lK12CVPpvR/cWeY/r
aALh7FRDseA3VSwK+IEXKYhAiom+PD3zcXXdi9JLUpYHosjdi1DcI1E4LvjNpk5u
Hof3Rv4Qwiut8FdUQDMyY2/Pm9b5SMsfbXeTslIckE6plhIUWFJdoDNUC7j3xsni
gZ6ZpV/Nj95mAA9cdFEhxvJ94TRmm2am1+lF55QegXPumONoj29c1xE2O8avd5ZW
MtfR0Mx1z1N6cdOAaJKAR2MVva9GCSm4ofJ3XbW+19IxtkiPHXb2YAOwLA14MwAF
NvJiTmgOif0qGNbY1Yeh6wJaJB2AXE9qs1wTQeWVpyBxVy1VC/c5sq7l8mzuZ7lU
+72cbCNNzd11fLzPwa1DVa5TXDFaduDG/K2Yhp1iXx40o6HFaZPvc/YLksoET/9o
86UiktwhCgI0w8q47rA+7PzeVKDXHeIh2e7VZSNdJmfTOEOafILi9PZV8xeo+wrS
33jyojAe0iUPYR3Vh2oQZL8zlpFDiN2+sTWGF7qPhlYN6z9+XSWrDE21KV9AwbPP
KtBwYgqJWD3gIWaY+5DnhiRTZywVElAM2ruHoqupLwXDCejJpEoqPmpZIMXevi5S
VaoWMFnedGWJqprX5QuaCVlzHBCTalsEXsFLVSLD98gljSInJ1jjLBHAxVvBN4+b
Au9dtu6acCg389UtXs0cJlpuz/xUsvEG0Kllz/Kq7Z0BfqJ/3T3o9eydxVjonNPh
MLHB/YTnkb9t8Ty2PaIe08RhnNjSIlg0QQ5E2mrqq0FGQ38PIRS7KVv2u+PwwDf1
8tg0O799H3HEksMj3lyW1a2Tx16+FTWL/WtXg6BC979g76OvCUo42NYMv1RYBT2d
0cyD6QJtCYCTo9NA6NrZLtRFkoXTBMgZ4XMajRCu9x2x7htIEW9lF7uIPMeyfpYI
zpdXDLyqNa2vQ8Y8CbVAsMXYAZzCixDdsFzX/aSP4y/coMETdHaJlgHLF3OK5qn9
2DrBnV6aTeBTRcDB5PUR4A2RjtSu8p/0pP8oPVIBx9cWCfZzIDDORdmHWGXKg7mV
wbWaLC2TqsYrpHERaD+IROZUIn+5qT/M7Ex9h4LfghFhDJzz+wqTfToTGarKERxQ
kK7SZNYjQX0FbEsMnCfUjSXEypHfCRrzRuFzPkXxuT5cxLBKbld+8DrFdXXXKFJ4
xbGDRbxMTbrSx5c06UlQdgoidxNl2elRe9ocnyU/Wn5WSQSDWMTFkKExYXW90zN3
qLFBYK2TZT2ebV9jJ7AzVDd8OYsxMeLORerdmsd6BCOvRd+GT+g5HlqqE9voBF4L
98Yr3cy3wyo5RMRUfeOALTT+ba8zHpoVp4M5NMRJQh6FBsbm/NpUKZt8AZzPruaD
iq12DwTLnGE7jhBDHIPWV6vmNaJXJc6a+dkez/6sZ3rbgi6KAYVA8M+0dO9EluLa
yoJ+7LNFmEgyZgLXaM+88vanGV+EKYj6UHK/Kdtk8GYAaRRGzGXzIPibrfvZxU9P
eqvUvuziSxdX8IpKKl3B1zPpXXiQsgjjZnjdPk3Me/8lBuVZQmRQJeuLumovHW8i
k9adJ3h+kbCX/DEF8JiTVGeyuwPeM2qOkaOAsn/80Z0LW6E1eiiRhhdk0M7KdScy
jzntjs4Hi5Y//DcQlylrTsu7pwIM4XyV/aJRGBtKLnUq0qgmmN/Cr4ONgS/2Pnpd
gnDuVwe5v7WZ/Dd8YrRoX2P2DwmWeVLLYwKmB2ZPiPFCIbfg6Z0hdcBaaG5q9/SF
uIAazLEz64oTqzDOMuCBZoIGFxzb8bG5b1LbON48GaKJLLEbOKpBRzAkdUHm+pur
u/9SdIiWzN91HUCQ5G09P6D81ZCMDZfTrSSjVeZh7ikxchhanYkk37bufj5T3HTQ
G3K6azCUQFwZ9OjVZ0WnH1qnrvJoGHmWxpsAr57kroJLXRMtVKW/DQYruNf3PO3A
sLrGk3Le8SbLz1ZaFPu3lU/7l7h5xBwAtD9Jx1bs15SBlh7vYyrLPsUp4YujH3YF
swsM6uvvglALHaabCydYuMs+1Te/KVjnkPgshBg21ArVCMekXhNIrCf+24UzQccU
iZSqWOnLwJVXRgPsfz+eBcl+RQ4iWgb1dqn07c4IJ0zOueJeM0xogBDz7CsDbFim
VeuwWCqnAT4e2bFR/N3S1bWx0USBKCJ3+CRsHtkGfxPYxCtZ7ob+EV8IumT6lYi4
bctp0g/0ZaDPBuas/svmu8SHXxpaUylTBzNMvD2HIwsQnqNH6CSpl5hptOTLCCzt
KYsO8C5/0ZgP+A1tMZju5KcJoJAMLEKcGVpGclx6So+ACm50K7hF45zL1edmQeL0
htJZVWgqOAIobsJIC59YahdsGMCzvSR6Xn28HD5j728+P36k/3lgWU547zqYd0dR
3Pj6F01WcQBW4WFPGzE/m5SpHGpZ65YwrNcyxZwnYM7t1eM0snuWgZUGC/FBi3fu
XfRRPSNRfW6ENfXeM8vRg9UUGkdERMEoofnW/uipqg4colNZAyM4JzQ8s9LmkKVo
1u8Pj3S8W4H7PP+MLz9Sg6Elcx3aIfrL5XdoFkdBy2f43sPDrBYj9K7klgLDjBnI
iPVwDHdQX1oRrBkhECXD34MHw2sHyQahrFEkZXmFa83rZAFZY6aA+230fLJ3ZmAV
1IPvYT/XHDCwFqeLlk4NNKqDI1f2zkfRIpaZ8+LRGOZ1nQ7LeLWCVwhIohmJHC6e
d5Byjv1lJyPqiIXEue2TePpOZK1PsO8u/dr1zoMNwj0b3OsJuVFlLI7oB1PZGNjo
tU84qSVcMDi9hiza+VO8w64JeSokCOMGOYutPVO8dWYZ0Beq3774z9BlhYnxYM/2
rDD1BUflKNf1TKDkmZ8k69baimhLlsAT4ZsCfA3z8SLIe+3qkYM6BP6J+gJUjqmX
tv8m1SwAxZWgZz9zNPaDjwoXSUzz8O177kjxkgwSNiwibZ8YSbLRlnnUFG8+5KFz
/D3MH4q5s4gzYIjNoFkVmMpOOAEk1+xgqr7P2CPziAc2588ZYVnSUHwK54D5jxvN
HK9Ztol8/MIrpKVfHZj8gam8eK2p6tXGegQWAgrm0JzCAWgm52fF6pdCFSleiLcg
+Bx6H6vlxWtzd1AGbvM/opv18SxlzRH/3y5qfi8Zvq8bYq7PM+wkMdIUwoqy9EDE
sqxbH+gFeIZnz8iYPXLvA/tTeSba1DVcBJERMKv6xx/FW5C//O1TfT4SryCkEqqs
7CNYYfUFAZm4V/v7N/oZaj4HsSkPcss0Rizp5iGGmRsqipjH3U6hqQj7KYiS+K+i
a4G31UVJGfi+aGEU/9KNV/egi3CD3fT/8PryKhGEMFVhA6bbVwm7WIoLtJAZg/Y4
5DI4hzM0A7RtmG53NUeXdsjbzdCEZIQItW7RafRmdIELGOm7BYFfLUi8zg3HNN8s
FOK0RpZWefWZ1TZWQzEQ2Mw+WTZWdLHMRQiq0xdrO5sanyLZZIc2h/DfNSIjdFUg
ZwWjl2OMX1ybBji/9jsQy40LTQ2gNZF4m+05bgBd48Eny7dc0NkxWWKBd+0FaiPF
qyri1QUkPt7kgf9QjPZv41ma2g/Zngb+6Db566qHnlADfa7b9SOEsEk6vAYqCJXk
ilFdbkFyEvEiljyppfoy9ftMOAzlh7IA7t+cC0UN5XIoUoYqgjWHDFDE4IUXDG0L
Op6QZGJNqZt/x5N8Y9SrQMvzknhOkZC3xd1nHPeZ1nXLrDm3jyZTdCkzTDk7OlVo
wiNYm4/WlSqZfnFHntSiKFpalmFYCTdVlsSsx51Cq3MqIOlC7CJ/q7CImaZmWcS5
5Uw6jSeEYbAhgdDnWKbv1VkmWN7DOsIvlust4PZ6QL/wYqn1Lw2CEy1kRKzrX7pb
QF6h331HQSyFttbo/SGhE5/AErL85sDYMWiVg3V2iKaNYogN+hE4P24TZEX4NDMA
y8Lj5Ie+oFKmaG/P3JlmBVKY2ytHmAETQfaEzeGmCgk22Zhufgyjpsp2sjMtnCYm
tkpz8EI1fe2/UNHe0AUsvnYva3154jv+v6JZIWnJBCgP6Uj/O6Lm8W+WnBWk5QTI
+ZUsoGdWuWu3fVtNa39vZWOP0+0koU+7mmclg0ZcSf1aHwpYbCbIl2tekiMhFzAl
OmBhpNUi5cXjuL6+GOOQO0hmOX24yTf3USL81oCM81a7mm2RemhtzJStsTLMxsH8
Xfvn0yydPPecVMDzojN+MAgvcbLMuiz7PQZva0SEG2fJGAxolvjiBDX5TrLFB71v
RAVi20Bp1eJc95BgHpNmc6wn9p+jYaW0mI+2oend+TzqgCG1424RQqfmt0Jjgh2/
5BDXWFizz2EDyqm2vP800wStJgjUSjcjW7e7QBQuWALU5NErTe6JAQYrcGiP+ffd
AvZzAbee6p6wvgobiEdlgyrHSYXA0cSoVDx3qSpQVyh8+Fyl0cyb2TugpiNKTLK0
uGNvSfqJilzQJ+THi0zz2ZLWP4XA5vCKPG7ZGiqcZ6iMHaycYLiqVbO7sutJrCHq
KkOxlT2mZPjBDlQpgE59QnR5mbaP6YknfP66oybWkvQCl65kHIpICKfhlEv8ng/9
pp3LbY6rZgHLrGWWAdth6NzEeHlUFO4JP+Ko4OiJAEr0pEEGNsNpa7FijuMuTh4U
bHY7Syx0oSGa8CWfcYezycq3KDZ2fM4NTCzKgk5S85xDwrRvA7VnAOlT9osUEYHv
wa32cRtcBnA1wK3gbVi9vBC3UcFxpJ5ZuyiRcuBv+aoHs39xUHubGb9P9Y2dD3zU
b4EE4qk9gVhBwx53TlSU4NcAs0UnXWWJz2LBXkXM4qoLEntE4wYW+hIjkfAKMZgw
LYzDy0Ysh3EgSSj2AJvXzxFDAlIL7jG5DEP8a+vCF2DVSYUleUiC03TnrkbjZgZk
pE1aAXHV3pialGVGL1rRQ6Fiq2H104G+ZC16EvmTHiCVR27mdSxKZHX4ApzqNlxW
GTCyBk5txnyFCGQGCWJMnQztMvILb9Ukjpisddmc9C9WdIN72YbaCx9gKHCCrv/N
vkNshShqjyKTVnzglUuYdVRP8kSdUNhZfSZ6nUo3FhxDi3A1pfHqNWhqsSzoONOC
yqMLQ2WnNxZywxMZbjmprgzICe1P2bxF4wUxO6WIKImBa1zl480TowGiYbS4lh7m
+zapJJ/DaCFsmWlUPDenNn1l4lDrlQGrHJISVAsR+il1ZtNUxiKBgRw0tqBhdsuw
kK73r8wOXP7aLNdPseFDmfab+mWcYSO6Uy5ZbJTWfQiY8dPvDP6LxLZSJ9oKLHk3
/FdoEvcQ2c01VfYSC7dLx2gTHxk65igQRmOVSpN4b1l/pi6iU0x6gnI0En5ctrWZ
wqTJOyJzg3OQICRZ7UUvP2eCnRXEwXcIOnBZG0t4vhonfIkxd+IPzL2dNPWbuNzS
97RNgno3M1sMjplapz98+usLN4lNorRV21wqyhEukLSql+GRufuKbjeWLEWF/xD+
JxohO5+3d5jYjpuB4djC6Rpsb9peqk96BVdp64vMzrWhhoZ4aX6p/zWyr7yf2uSb
I2OIC8iQGfNu6JQuCHkjkFZ7CW1TTM2HoxT/5ZKqMnymdIovqBVTOghGPRg1NI3H
Ub9/DaSos4Ubj/lWu9cBgIp73xazcMvWGJTzPolw+BNY6p1VlrDPIy/wItsqhkAy
s8H+9MGq9SWLLvij/SBmhkeprqVp4kUmFxhnwZft4c5/5uQ61brkK0hFRjeFMh9w
yp2t5VEdcPeMToCFXT3B3Ck6mISvNB4Aa1pKeDWvHLPVdiH4EHrwPOq4mt8H4tiF
xG+bcYLOuVw1u5zVSHCs39IRdz/OVC5ZZ1XN+5z/1cUb+merP/6GiW0m3JWQZP+K
orgeI8r+CUV1iEwTFBlJXxATtGDtpdBPTqaiYAY+H0J0995BvutnJEPKSaUIKrCe
NoWsXMbVQc475/3zhC6sTywvgmimA7LqgCIVMoVXCb9Uw0rcUTAjamZmC6hJLIy9
fu27UU+mQnW5VBxTRTOdBMycps5Twly3br7ES4tp147vxr1wCaYt5ykd1PdHc85D
UHyKwHRp7ZEesOiXzdqdQSTzRZOQavCkWq8sDEK5N+2rLgTcRSrtaUxBEP7GKEC7
WUJSj8QBvLtxvTkAlPlZ3+tkmozz1BtMErwug85ipe3kdfKtW0yWKNAnA2f7hSYv
IoyRkX6zJDD8dj5dbfVLW3ZLKVT5YZKJYr2JuEk0tTkHWzUum1xGWZMjDA+pf+N4
7NtQ1C3G/KOirxyhRb9CqjAoTB+ERakpewQLq3HNC/8PytpaP1DyD6JjE755o2u3
EkxdBh0cgcEFGp6TQZceOfFvQuJFQRmdvepdwVCTUPGTjnxq8FNfVjfQDq5sEV0L
gv2cagBw67EDbXShDWuAG4ED+pvEy+UJaWzOMVEmcOR4V/TsxQ9bQQ17MuLNYtNi
5Co/2dr2XvigwnHpdQpDNk6DcQDWe2M6kIlJ2VzXR86eJxXV4gw2xdqpXkjwnQB9
Kfr1Ag5znAsS/SOIkHkzxSey5KSDYPtUkRZsYGqElxGeewKTZ8h8VRQsh8fhD9SK
JRtTQaizZUDT+6zKBZvRemR8rSeFwST/5kqfEudbqmP6hMDMRJaJch5p0TOzojNO
QJCXrD/rQVT0nFTDNIenyFHOOm+HG5+LNwv5ccbU3ofbU6mspErLH01TamOqOq27
FwiZQ+08mb7SzRc7Gp4d34C5KkJNEaH75kMMYVv+Td6s5mIg1X3CfIdu4hCpUGTM
WMzXsQM42jxBRZ2EwiCBbDva0+nDlq/0DjRKzJRgDUOGs5f9IdUgDTY26scQ2QNN
2DHXAhINSwnbS+9kx+cTSnokhLYhaTMRLOnnZJo0q7OBQ5u2RsOiklGq5JfM2UpJ
zaDXmHYILHfW7feHl+ExuEgIPWE8qPCTiK+qXeV0mGZeumWyvVo2+zWziVK1YKSJ
YLKLLlQIbNr5pGkqXbnSu6FP1dPb0BJL2OKXsfiUdvZc1jhf4qEZ39RBjO6OGai7
dXW+TmM4AjriWElghX5D/B9/Hffwmjt2gQYABufOYC8t0wslFZHl7xH+Ju9ZHYTp
xq3NtEO+/dp2ktzCeNEGYt6JP0ypr6SGJz1/Xvf3iFNk1HQW/8ktKRcvgusBFK9h
8S77d1TkjnwVKfsRKPS2MPLdNvf6UFCCN9Z61TuOM8JtWEeycthq2WJ4KwPJjele
Eo1wbC+kJM5LWShhBNUOwJlCQ68ATNnnsf9DKjyKEcGiE2KOtmiRg+HRNfNLNLzz
AgdNR8pcqAcE0doXfPI37kxHhkVI2GqxhSPJu2E7A5Aiglvp1VMCDfmyO62glgrt
RxIR/VoOrNZM6ia5OU+KkAohcqxqI0cA8m99qYQf0LZ/7IqRXEi4fL3K//i7mCFD
AWv4Wfb/oblEB8IE4jFDeEhVSpmQmY4v9+CK9MvB3HD2uRebco20/Rqa7Ji2o0Gt
AndSBCq+jZ+WtL1hQPR8HydamNFbpno8JhLa/WuACfP+jRpf5D4QzooGbEcxCJLu
pbuirB2Y2zlWZYp5ymmbBmYlt3UIlGS1k4NsDspoSe54WU4POmDPXGT0WQovmcIm
CEM50PquGuN1NSCD2c6byEqTGuOhZH5byPbuo4K0dZW5xWg5qAfc52+vVI5peB1y
9oCg7m+sXTsbqlGQpzL4P5vxxiTB/OEcN9WHBz+pkXfF3mXy2lqz7PfhC86JIlmH
2p5SB5mMs7bhTE/QUnvePdd8Jc8dfXsQJCVYTdm7l7F4QFuK7m9VbeY6YbtQXxsc
1UFc3gBWTPQYeo49xIymkUfJ49HDEXoW8oGUEMcIWMxaSY7Zjb9ahUqmRC3xOhYU
QSQOGFS7WF4Wcs9Krb0aq4A8SvGswRtCdEdanakwBlqVHS4PySdR6n+er4kV2Crd
A+CG+NxsHFShzKSRMvJNZbHRfY9tRNKJhNUsGFV55rdn+QTfql8O6M/4Fn219BZ4
z1NjbJfFR7IsrMiAyoA3ebhPMrH1sopSCUO9L/BX5wJKIwTN9fzh8cN3u9iYAmBR
82sWFkabqZMyQSUFSofw0vgaqqEONr106FzXrfHPJNMfmHrqw2WFapGY5nc84IJ+
J9oE0W1JKGZxTPcc0ssrsmY6W1+lPZuHrGn7PpSm+QXLw5Pom/aherYaW7NriD2T
9EbJf69XI6oE+aT7uAv37/IkOPaYVn42oOvZxRlsin/9aJHIZMDUaFAAwxD3y0Ve
t1SLw/OqbBHXe5OBQgSxMTJd1DHCApvxmNO0hLDBtnSoe9sFsM5BWJA+hhLDK9t8
HdwaKCAP+8ZLMBJHI09/9Ub0RlSgEHy6StAj2Aj7TMvj4nWjeY+rh545Tf3u58/N
8bckxESXTJAgtllWR9Y340lEiBdAxg4/aT3+EcXw9K3OSeDc6yH6W/9t8HmMKLJV
mUFbCOZ4V0e6WIWl5WWyFRj/etE2GRY5rOhJ9tklbfYCzIib57WYZ77oNiFXDcrH
uWV8HfcElz+VwMgy023YeCsEKwmcFXI9Hk/Z+VVO4X90PFMQiS6rExyU4xJyNgmr
un295mYWYSBWlrlV4kunSkHtzCyMH6laDu1ACT3iq9tzV+sdd/ZFLJ/j8x0dAlLE
f92vDfm0NdfSylR84IY5jSC+rymFoS0vPiP9JMHeLQyOQLncPRyZnxoyAFB+YFyi
7r+8xGuYuLlZUPhVbmKZXaLRNnpUekci94dd/WfnNZmHjCNqtzivj+bbU7rng7GT
1WvYPu9dAfLcKV5S/TQ3jlDFXc+bJjDAckXkIS2ca5ZGTXWa/kp3o7+7p2Ym920G
krtPiSkVdcmXhW+iLToeB4RAhMMt9/a/WiiV5NzYDFGHwbU2s68dmw/pBfIdneWa
pSycK5AFhtjK9Ml2f/fvZYoJ5Lj8B6f8KjCrG3G4LbQMNSA0+J5LStDNBApTdCU7
P1Z82HNE1JjKnCVQ4I6g90hi2Oe7xDZ9AQfmcpwP9PFoWuYgKYnpLqKp2gO9n4Ib
fli5YHupQjldEPoK5YHryFA2Wp0ONWQUNuig6WlDRN8JDhkSRwDoGd+xoXz+5rIF
dvkXbCI7lpApI4WEEt/mGiqUf7MJDlVDSTYxgEmB/ltI6/gckAIp4eWf0A16fS+o
+Lul3H+bF+dQsIw4IjMuXMWpy+B548YVNTLCkSYchTg9DlIrfqKQLkheJpAkTUZU
ENWrz5C4UNunm212hCLfdFBcAtmrpfuQaWxUnrdtsmEzqL1KdwcADEiS9djuc0Xv
EXy0nfteZxkuT2jsBmtyhTYV4Sh9pglPSgVNzQVpy7q3BgKzAOIEyiAtdbDdlrC9
LPHyDiNB0Ff7tNyGmlCWFRYagcLV5hOZVp0IP55PkZSN6UOA2XFHqwmTvLmSmLaQ
bz0ZIbHycgoOiUvhQVDw2lfzv0QPkXmQDjETuJT9YAgvVoFwWa1oaLrCRaVnRmXe
amQU64A7f4Vygx9fUZeOT5z/6eAyuOcOElOQ7ct5uDEbhcxqsKIbDKtPDyifwywm
yd397w31WQrb3plZbGvMSQd9+BIU+Er6sAIHim3Bni3M27af0qd3E7MvGyR7SCPM
VYb+6BIjqKh0P+2YKM7ELGjLsc2VEJ3B5cYkAYh32AJ9muGxCsAa9G/iWlGvgvVI
NJ7JztMEX4w9hsFYL4nSo5fuRsBsRM5WNl3UbekZlbz0TFKnnqcpNM6JfnxGZYDl
MbDdEXrckin5j4mp5YyCzQD6kPNiTNryJTrxn7hoc+iCNct/Q29KWvXE4WiSzvcR
Gci4TRPB0Ym4qlnUUfsMZPCxU4ID0b6F8RALNbhdrSiIAnWLnBwXK+1Z8CINs8pU
6VTPF8/lLUDLKzaqicNST6AfwmbEM3iGCsUGbHxsPtqaolCvotKduqgneXEKVkyU
lJqjhWBOB0myAcczE8opQ2I6pp6OnFirkFqYWU3z3PkoDl5M3XyBPH9Jg1YxfQu7
6gptP+doDNgd1ZgQxXKQ+Q9IrqG1jTycNFoVLileVlda1jf88YrwHaluEseI5vZS
kISRxVeNwlwFOoQWUNY/APosKxB9XER9EuTDYZHsbOcdXkJTdyuFeZb5RDBtE768
ap053zdwJ2f8yBBvXkmpkjaskZmbvon4DPckTqH5Qf//eZNUn85GYL9C2rKArZEq
s0gPXISym7naHDm85pJaIW02g0qTnI4BuLevRXXSHVlcb5wfrNm5mag4My/Vnbar
ksTcm9MyeP+4sFEJ3R0bZ1G/za5/SrTWkUd1ywqnND/jN0k2Y4BqRiSTExtSt7Ff
dDFUsndhEaxdZEKGh//p/0SH7NbcMbWDsQk1IDxIdTldu0qLsHIJDIhugTcBCqbj
D2VtzXySEIay+OdwRBsPekfE5DbengCMTUtVkt5vagJL0lyYZR/7O7G5sdpMSgjY
FJwDJFKSHrCtFx5OKx7EVlGcEHCKCcou46nKevf79O+IzfjkxUyCdkg1H5pDbm0L
La621lW2+w2x1+xLCGgARN3rAvQ+NdW8JhHEBJeF9hBURk8YldMHqYbrKjcz6B7r
HMboVfn7f6+9lE347iFkUadu7LXePg4jos3tpHnoyq4aqqFf2INLz0ZARwQnqgXR
0PC2FOhaBRDT4YOHiRaWo1ZHpTSfEIX6GPrgtiwSRfwaqbtKha1pW2OYgembNg/h
qq9H7pfvLDHj382NeiPb7wsHYXKT1G7b17JR5YlPVymrU8JTqO6bL6B3SrD26eEK
t41kf4fNqZl9IQYQEseMRGJ8ZVcRh5A8m+VQLglnXVXW93nZB10ZUPam+DdyqFZl
t3GORiHjTF9Wi0ZfM8MR2urVWuT0fmeCQXOzPfTJUgh6hta18kKw2aQC/yDQvusg
gnpqe8XjnSuzSbIZ0NmBmdC2CNN6lkVLIK7BFrHQzNyYKhYxcX7D3B7ZTRgb5wWt
y58kdwohQuLNvmngvy/BRv26J0BgHoZJTZ1+diNL2SOlxILxx0nOuS46VbaGOsFv
esk2Yr2WZKZU9+zOiv9I6kCwzm+tupydcDT4wRNYFfbmSiJOZ4RtTxhArYn88rLP
EUHDuDYTV/A8IrbPTIQ3c0FVHbxRzyA7MSMa3JVDJFZummMhvkyUMkEWfP+61vtr
5hkaNGsL5mtZwaCUmpa3W9lSj6nL0URYtqJqoSyShZrbDuBki0/SP6BxN7ZTYVGf
SYwVdl2eY15kfeV1S3H4gGgVBNdNuc9Ugr79npJ97xzlmxScD77WAoB8AHJZnHq7
Naibo3/ZfM7hgm9Y4GOoLHPycfQJiV3dGKODzhVxBwOqQAUYD39e8WHCgSi2tLJz
tDSzYBYwCRxtAGzwr8ekc0nT1iWwrx7YddIvNQ6jOnywhYor3yHOu0ZHIc3+26sn
XZShzINPyElVHWdqGVAXPcbPi+kI0tVmdfHBb9JPtBLUvdMef6OgndxRVWObgdPM
lbYOuSwwdTd3pL2fdCD2WYtC+Kt0kF0OxMDAvihVj4POLg4ShPncla3dMcTpy2O9
XF/IWcstCUprDOlgISnLYVK2gCypJwwfENrP+ZSX1GOTy6CEq+SXjuQ4A6Adm7kR
W3CWmqv5Jj+cB9RO/cTHYfA+OQ222VOyGwsGaMT6f803AXjBVwmqIujArv50q7/c
hiKWGxfL5IJrh+jys10t8MzUidKkcn/M/GFZ4GNfjosOA+lxfE+pgJ6124FR5srF
yp6ksZQtYraqJgcvmUasvQSPa4Ddst68X29Zkl9Z7Wdb0uXrv8I7tPe2dY+ftVmk
FbntP1XuxskQGdDkztPGRMlkwplJSXzp6g+PP6494Kfa9D4iU30GWdAh8GMBQ9t4
Ct3T2uLB8g9WOohO+DKtzX/6VDUQrKGAySk+J8ySDFLn2S8zv184H5GKCj5NoJfu
neYVsYYW35HxcMoAs5t+dKYMtLufZxYIBVl5aWRKWX5WfkziP2KemAFrlO5dfaII
qlGt3zhF8vwyQSaMQiJeK67jW8q25Ky4ztoXh1EOIsmzLRV2un1PoulmBZNfrc34
QqoD27XkJHaHrFjRWXTaNhL+j1FsqpCwspVkTaQm+6LFxs8+H4OrHWmOEekfDqQZ
+DMMVatwaBPlU1RuRMPgPgLeYNxLSR9m5ndftQp2TROYXqg1pEdYKvTz0ToVNebA
yrSRl7a//ddzGCTPSXmkD9B/LBW8ahArSAS6XxBqDeTDTDMYr8sFXHRMRXXfG6aH
HQgEmumdb2NikeZ/+krg8LxFxlact7uGXvptP66pBuWYAsytW8WMg1OLi7DxtUl/
51IuDPwpWwjCZRxsm1+o1hqSh3Hp78a2uP1zn4ZMMh9iBuZbWx1NsJopPY+ju7rg
prYDOqo5IpoMNJhyAESwI26EgcIJ3rRqOhLmyQZmMi7vjRvT9f33nv/FJcC5kr++
xfiL+NGozBOynIO+uMNs5B/PKHCwBWTGg9twhgH4TIQd9Vexn3/nKAU+8rT7kefC
KTkVi5YnGp6M4UqiwY5le1fqvdK4RWBMBVxgYSN2dOSNzWuUyVmtgRIrzYjraBY0
z4x+W34mRnqDirvTv+eba7g4j2/G3hGmvPVBkiPOkcta23WBO9Lv3rZhiMWJTo12
HErKfiKakWqWiBJqDQoqvcnE0tmEfQI6jBEJcgKv+2yC3xkh9WVj9o7tMB/QZ3OW
BWr3L1zuck7TGiGdUCWTXydUHufKAttaG9NS4J0e6byUrY81uagmtZe7hQg7KnO5
YyxBoTEDF8191dfNxDJyMnU8wx/pRZ9EZTzEyUWadMWc3unKevsi4CiFSi95FFjH
bG5a92Qs/P/BV74hnLM0YVBdZY2Z6FfkP9gSe6TH+5GZgfDKUx01oSTmgyPw90wR
e3RLp0X61fkUmhTz+E8X2Wv08PIjZDXx0GngK4HZV7tyLzWdcahzbJkevxHonA8V
VqWlLaV+IxpbMIgijSHzjhoqY92NaDGCBwJoqOu9IupuB3UhM3vwAmwSKrVZ+YGZ
Q0+rME7yJ6w5lvrMA1Pi5KN10JjeYYrzwrJxFX0W5v3Qtf3Wpigy2GvNaoI0LFtn
vUGL6914Ocyz29plHq88BBcIXJ8eOkVfK1KkTeGAh5+2W7GgBezqF9Nxu6Hp26ot
NgsAisqzKHOjfHL6CumXjnz/8KTUDLQ+b26jILZ88wtL7JONxQVcuyCQUlJezqTi
nJSitgcvUwGezLxF/jB3i9NKIQb/RgvyT50DSZRNBq83yJzLxZqEZd6WGtM6XyeE
ty1Dh437iIzAvYxbUX/Yi7GWiHGkC/DN1N3QhUnJNXjokLq2xMoaQp+mP88BPnzb
IhlmQDNd4eBbIx0gOUwTwkLivMvly+QglS8zE9aBtCYh5pGIHKdoj1++U/bVTXBB
sXxMrDqzctes1onkEgaPYg+HDkgX+cCNogiQk7R4vAPE4GOUwHcNGmsFaGK5kM1F
WQhpjQXd6dVgai7gcCp2P7UlaYMU0kxDoOBJ/npdnzk2cG217wVgqRtQxB3k68lk
Qz7g+V1VqMrO6Jm+aln1szE4FeVwvITpYmu9zx4P7RM/+hwhG+c2EUSDy7R4hhLs
dZjuH4mUUaEfqTi6TQF5a3G8DxwiS3LeR/zbgabN+pY0VZM6D5n0i2q96Sm9jAo4
S8MHRP6qc4dIFxXVx6KFM1AtsCkzOvym3BD1hgwFR5raIeVpWd3EuHxjfaTe9wPw
a95zv2AgtnE3sxPkoC0chBYiikhVQkwMrJkt4YoQe6R3ZVX2BgP/NZDui8A4jvjT
Ch3EcmP0uJ60yVGfjWjuzEOZPKaiHLgOEDtl+dNUYkofDyXHtR2kAS8kFcMTbbiL
33NQHfRHifgKBYe6YyxS4cwX1GWGL8CCps1aTMMBZ3ZczjxtNH0dySyGqj1dOonI
Xa1UoZFXJkwjb2EUY/+kGgUDdrYer5N0AvKkREoMwf//9UgFgzOk0YMNagXNqBe7
LprpdSR1K+lhWKW6nhJvG+Y9+xRYGnqI0H7gixeb6PWvGoggwIdVudcedB6kkN8c
y7XE/RoYCB8o5bSAlR0wimFTzwFTwBojA1l+FsHIcGkOuxD8TmmvTzlL0VWTYrr8
CSxpLH34oUm3NwRS5n2Syiyvr285lPeLQHyEKhSGAdPrafa4sT0ixzlSV5wRzpZv
pW1LziiuCrUe+Hab6ZBSIBkWpVtgi5mOxn4YCYdtHFxX+yUhtGn5X9yemIgnRbbq
jFkFvgkir1UPHVvv7WmvSO/hhoneUBoyHSOpyVaKESxwWuF19SJKn+UDMyKZdAUf
vN7tvmfpUbI2vfHRJSlhYni2RP8Knj7QMV3uTU8bFPuSDE3ZdiTD6f91ILa4JMvR
pINNwMzWEBIwd2n1scCMoJ/Wx+tQeny1oeQwUg36AH5JA/Mr58s3q5FTp1FCvtX+
3TLsS6HYrLoQFb864Sg0yoyaymWTsvMEF3KbNZjWhRg5GchzD1khcat5jZGj7pcz
diAWklgo1ozcz11Vf4Zsmxel+7waW4xsueKpHNptgpoY3zYXUee1j5dYrpUqIchp
WqVtuMZa6wV0ksd9LDKc22g985DHSLVuOlYIRdnMuenTnjp4KIaQqUCSCMBYnGCY
B4IRpeRuLQl4SY6RJUcbg6OJXU1uxq5tIldpSIo1wPJH6RMu51XYXsnbBwB0nd6k
B6fEsLf/vXx3DIRpTzUgvEsejd49/mujeY5RI569BtbiWQBpwFSvhku4yeJl7Uy1
maBmZ4bEK3plIJUHxO9nA+wQuFa+NC+lKhgxMW08UByjwClJ+xDO54BPeiY6gw3G
jmDsHQD/CR/n0gXPas7/6ta2nqummmZFgslwEwpDIk4ZvGdzWfSd3DRzE6PfRtT4
xI9yVnWFRBBfu8D9HZjsLkDnAcKEKiM1mPCTPUYE9U/PeontznnPrtM/+s2zISL5
zLajgaA1Xiq0wGciJ1ZiHhxpKWrDbhAZm1lfrDduiYsNa3nCS2xVnYfhu9Ar9La+
E3zEv43T5xMTetYrvmT0fcbYiNgumrN8Ar8BUsHKNBh1WCBKBlVB0ha4bqthJ3zY
swYHS5SyWxgP32s8jlo1WzN87qVWRhwt91lS6BTq+Aw8Cc8X7gqVJM23ggNhF1if
uaAwbeE4h0inAVzLr7SSi+gN43whmHIV+LTyx90yLPgYkxxMGwpqSFrJDTy77lTk
HDkWYAK5vbEOwLXjbEP88aLsI1QLyvAAZDIn5/Iw5durJurAtKtysWvg8goFYld4
8ffaTxPUj5heWwhVmaELcC5OojIy+4nYHqk+81Y/rrDjp2quRGGmqXZB485MAcgg
4tf4JEz8pXT0w2BU5CoWkZkrsEJWD58i/LtxOfR5l7MNhtJcZ3dThlKjVpZmrWpR
HQbb/icC7DPT4/8oMKbP/PBaO2AJqDNGOstsnuS7t+l/eM4EhvXMnFI01TW0Fj0B
mRmbR8woJSNlwt052TVRr5S9h84EpjQFeqDkyQY3j5ouIcUYLYGQ/SJpK177l2yx
dQCS1F7Dfi8RhOqeKBph2G7G+jT9vVaE70SN8+nMvXkzNZmnFNNflHPusAY6TOkx
Ybi/fgxesXOwKh7uE5rCoOhyVXfyJNPjj7SII7klwPUGgzDbVtgmWHUv3A5iCi3g
RWZ9veSjZCuWBcPlAD5K9lzK/QPxMJJ7iTvHHrL9kRSmmtRgjbQoAmx+mgwF7oQK
YU78CKDO7EeCyUBBwyGP1/RcHkPOZ7Y+IJE3bjbSxjgHjEeVljtGhIOH/ooC0uvh
REs003DTVCp19sFAHR6f85XiGHw/s18U6RxHElj8509Q58tvEeY8vUdo65od/WoI
FsHVn9ev7gKgtZynCYVJInG0V85Q8Rh9Tdo61nwtpmCFKAwxYziU6B4ypB9uisQ0
yvBWjH9ZM5R5zICdYtjWQRG/THI2nZyZrIvumvxfuAi9woPJ/RIIQvl6JI3AdtfK
R3M5Pbu6scE8nlPphpK7VEGRfxd54fKnKehH97exGR1bmVQTzDrpoD9dAkblubF3
lL5gR3Bu+yp65AsVj4HzjNYcNkJV2jOW7SYJur7Rnw0ZL79IQ/3ZCF7L5wsZ+Uvi
yRz2Lg5v81qtu+SKZmWjP+ixdwagaqSLi2fSeOE0lyDtCrCGJQSoCn4KP3P0pNhe
Yr/3/abIloW/1ysNh53pfKruXuYDdccQTf1hwkq628mrDCcKp/H8XnVsu9uyt9/A
ghiQT/nGvImu1NS5CVU8rQN7Z7KI15RjsP0LrVgclCu79gyBCxUh0lMFyUi8SFN9
XKmkU97TpWqxQy3sqI1ofn/eDhOQdumtucE5nLhtGpUglmft3Zrfey8jWS+wqnN7
xz/87yeotAbLDCata6aBn0gGoqs46GinJX9mTCuV/4pA7qD9/q74RR1wM+ytryPy
QDXG/yx8ca+lMv+QP1e1BF9cEvQ41/h2KZflxCY/+zcA3Na8uTXOoKJrS5adatvM
rCpMlnPBabc+Uzw+3P/hx0onDP4IW43n5LXY38HHGVTR4TcccT5BFogaVCDEKvFI
iU8mEYYpmFmRYTjXluRrzHFVX6Vkwm+KQ0KEEBXnsWdznjmhCMjMC2Dm3qSKp3IO
l/Wc9CvTx/TT1MlsH4ZacFeqKPfRbNz0NDGERnXZwVi86CICLMO7j45L8QK9+7gX
JUHa/RTusHGwWPvIwVTWW7OIfgeKnuw1qC143zEDVPx59PGGmRYWlrQyvDwHYme7
bAa/ODMczpnsNk2Ts+uKcBndrtac3YLQEz3jiG9IrECJ5eFxv/aUBWdOPOhLYOWm
5GKqZM0au3UeTdDjiORZAxRBKYjyr+SSOaetccU98J45fypUeTHAtFIc0VkTpwuH
WOjdCamQNWdfpjmnxaqZWbzJvYB/7wQaZCWx5R+5PVHuNSVE/UxEJWOfvpNylLG1
9gnNuAudYdGkjY1ByLb5+DBfkQvAdXdjqOGXecb5p/YOjiOyCp6nAbMP6JnbUFgn
lInmehbp1EabeUiqZAObxXaprfF6d3VsxrzUUk4HqV81liUF64v4lF6u1FdXwvaB
4cgkLRv0POW7TCERuMROA6PZ1z6n8IGMxJTAK9/vTWL5Sz2dbzgGCHYRGQ/BIbow
ettC7LtkrvNP1BAcyDYBKaEVo/GLib9YBNwVdjkr1VIwWvY+08EytrOBRIuRWC/y
P1qii6h2Gc54idtoHoIUvs8aFygDBGKOqYq0u3k3mXhXe0F8fUbV1tGIrtBAV5JQ
HJfHgcSi5IwX3rdln3cRF1b7jKo0x27XQvxMLJw240wFESwMBPzFDvFhVwQbxdTH
F8rKEVCVhiCn5L0UkazkMy/pD+FR4JvY1sO/9LgrhZr4Fd2XZk38Y+PNxL+oTzFn
MimuN4acZekmTD/hu1Grltj165IBnaW2GQd7WeROl8vvBghGNEAPUeWOluNfTU9k
6TJzTrSBunFmloDUNUM+pFy3KTl0YcpDwWFy/s+TmMDT2yp0Jjl5WYU4e1q1eAd/
oeQIBuDR7InIjg7Pg2algrAGgxCfs84whiOGjfobrc21EVTE/5sRH6PHcb1WdByz
zwRrYH5Pay1QFm0MdJfoxkhB7g9x32/UP86QBhreUOnZVSjOKopC8Njqe9uK0BB8
xuJpdYdOlt8fOkM12biH0iy5tLSrJCbCoOoamLuV86Cww04P7VnrJQ6OQyQoYqQG
MzpX1ByTdaGn0t7pVaA3YeYjR2MP6ZDJs60okh4XWUz90x3Bgj5lSGrquQi/GxEC
fVS48c8WE5cFFM4BEZerDNn7V/VLWrcr8tIxsSRjDYnopLW65clAs+aFXJgx88l8
5wSxhlnm/jCP4uxzeUOOt3QPaGW260t8ddBcbdqFYHOZ9qrgZB2OWjWqOXzJBsYh
TrFNWF7VCD3gOq4WFsu7QXfRwC6rB8gtR70hs1x2QVNapgzZNW83eyCDTifZACNG
rnbDOXXIzbGoGEy8rMqAQmafuECT39TCQgH3h/3FvHn+vhoywcn1vt3iWDfqnDsC
ouM+YLJLWDr3sdpIF+ibs5FJk8WQl+dDVfUzywlhsNvj3Br52mARRm1XojREcnyy
7GEKiDJaZn/TTunNYv0u8dcraFK6htFadwADnKtbOnN0WHgn/wJlC79lyV8gVBqt
WzJ5O9l+IwzwXo32I2BWdMjvtVVsQtyKlciSGBxngI9CYeaQTVh7VO47+qPNR0tl
hNjNonaQJkj4y48dpVT5U3vtxOvtojsuYBSpiYel3H5KuQzfxDf7Ab48pbHtu/DE
VVlMqjxprQyZKgA6zBXftBqwiWz83L2Y2d/V1Bm3yiXi5ETrh629F8qaILkZsXK/
PyMvrkoYtu7zg935CAp+HPqD4auV8lLcR86ssN87mSVmWf5GgP3MsFnCdWHjVBXL
OvvlkHNxzRvcWBCa+AmYSpe+UfZ7yvM0BBI8LLsB9XRxY8JrQaAwZO0v/egJtJ7b
/fM46XDs0T6FwyJLeNFHM/kCzZW6tKhvKVtTPFE3bnmqYgL4URj3IukgzkxI/Te0
ety9XNkcu4jANQgBwJcB2GOjVvCFTMwiILwgpSkj4lULw1bq5bdRrtoyGpwrDCk2
Odh4ORCeJn1tTWz2o7YEl1u45HmdscMoXeAfKf6124Pdd3eFrwWXJ4b78178/AvY
r903I0gfVKKRJ7lO8cr9WQMuyEf7jd7UgU4Ra3wVxpfNS11xP7Rf602DnjanSIto
DEMPwxXIvlU8uBGqeBmI1KHJROKDmyikG/u2dwW0ba6EZKu6yaVQBaN+mkmY9Pmp
OnTLxzzY3Y2KYcMS0QvLa/tozzsyNI1pl1ehyHQe+KCWsqF6J7NRXRgZ/jNp12cp
j6q11RG5tvCcvbGPb1bIPQnNhkL0Mh/Z2ampZGcQdXm3l1UJCnN5AsU1rgcPMP9N
tYTuTGYgyGZzvbKX1EqM/71G2EbLPkvWfcs9O8OzgtjukG8ROyBiWPmGmQVCpa+x
KS+rxL/HWbfbOpbTVwMVgimZIFktGeXcPnuHjFOSPGffbL9/fh4AINZoivuMga0q
CUiGjEQznCKM4VJJWj2JG/I1GyKps5qEHGBUyb6xd00gmaIxi3GuFBMq7zXkei1O
3B5fFli5AWIgWFpHEZoQfJ+0ehsBBq4Km2LxLwOs2H1950xuAMOGjGfQSC+qysU5
xz0fNrLOlXHDAiFIDC9RDO+nCD0RaJVH06K4cI0WTt03MH4lRAbB6PPUHTjwAB65
g9Q0CRg/0bQJHlrcxsyIQFyQOcSJg5yJOGp/BhN+Dw168H40ebs5ekDvNoVP2k0B
3AhMwkzpgGfG+jm5/63ObI3iptS7vZB9O8Q0Inw6JOegrk4XBZBBo9xwaEr9/jW8
PaJrTSz1mLK6yzf8wxO9vPwkW/6lTg8rHcQOc8xIzgwuCAevd4qbanYh1o/8Ew5S
95+AEriUPJPAXv8dcTZ63LmWx8UHgtCJp2h92AKcq2N9J+oMJdLqwXgsLoD+F6ko
dasq52abSkB/GqWvc9ZpqxZQQLHq0pJ0tevAXUxloLwC4Mc81RYz5GoCO+l4PYHx
Wu+P2WFGuEXwLhdM3b8TWm3uqXBwbnUh317XCDj8XKsPf0lRRqVYAbiS9m9xyacb
zL1iQLy1F0aw2gnfQGHghd0pXI6gYO2wCX2AKo5SotQcjWZoDsfki+521IkmrsA0
y29EcyhGdvmbC1AhvPsdgASxN+R3RQY3g61BZDHbhM0J5rEN0EjwpolK1JxcIj4D
Ka0FdWh7C7/6ibVBJzc2/pvWYKHE6dPWXsp6LYOQVppNq/sX05J23Dsu042JIBLG
5U02gpJbPQ599ugVGtAzxGjEmfLOFTEE+4Mpg3v/GnOPSOQtcSYM7s0AB88AvEle
aCjdCVMXPlgajQegLg7XfNMPWeWmmfkr0SF+b+1Eb2S1lDw7G4zXvhZIj/B2g12E
KsorijkA1QjThHC5Gs4oK1BKRb2yic3YcH+lH5b2FcUPyQHjVTgWq6DCleboyGcJ
gRwibqInnqO1FkJkXEFLPfHKx4m7VLWGC+NPPUOt3rgGFj5PU6C6yQ5YuwxJ2hUM
DmfDxCJvsGQ7Oj0XQAZIeMfuLv54T629W4XCc86GaVbPszMIWrKl/9diKhb3oIFm
5/BjduT/69KvPma1C4axuIuzCGqgAjefAY6y8g2NIMPs0h4jwPWaTJwz6LaSYD8S
zCh1K3Fbw1lPrmEyiv9LTdcOEY2gOj98qAK5b47d/gJgKu7DQcZ9UnDwBoa3byx2
7PqJ0JMkuZYAUty2JxaZMNnHLtulQilLdB5peDpcEcpcRKcw52Ni1dJUgrEP7HXf
WEMtM370JEyncMcqhyV4q/yzfNEP8EejP/mUFr2Ki3Pg0dNMG0UUCM5jQjK10Dmb
B7Aw26bA6dEwtbnE6oRQL8h3rOcM+jn1NkqEXg2kK4+ljVQq+BaJGVhlABS9AEQx
PDYxRKbed81mRySk5/7pT5iZ1gyIiHOhDDQpaWM0hNe+usKbKJnKEoSxzdX+7y0s
PHCWMhpax3QjnrMXJPRYNZ6AK6gjZQDuSzx9ssCNBrm8JCEqP7UUIFSlwW99EDP8
YEk1zEjmNPHuM/bu77MOdYZ8WBn8s+rq9b7xK18PITyFKLKc2ex08r+ZgmJHWk7G
94WEnZRAFlnY7nT+Z/3QQ1nZrGAizqFvqqOM67REIrMJLbvAG1K4OtyjhgKov9QV
+vYoumuXF+Yhmbt0y+giyyDqYRyV4II+Igyqf0UOmLzoSmZZG3KUpcr4e8CdqaKb
adNHuFldDv8X+X602xydF/ePU4b2wlD+0P4qrY7a3F3XQZw8cC/YN7Ncyzl4oVT7
d+668zQmrQoobb6aIVzKWH8RmLDN9GfStLL6+2/z5AwPonU2w0QOEQZa9OH0qQWx
AErSrbP3wb3gwUzp1LQUjfTjvn3jk3BpIctBAlq5VokGX8GtGEdiiRbDrsmTMgA8
wbfnqakWUxGJwtgPMVewd35bs9KTV8UFqrKzI0OXSVVnAyWznLYusCa9jLlL+Z+o
jcs8YEZDlYdrcGSc6j+BspCmnEK1HqwSxw4cZbGpf9g9FsnWe8uyWVSqLacXT9sd
7RvYWGCl6fgOdaNgSmSZjPT1v3EqDp5tRmpdNPiTyPTQQByv0OJqjZhKu6vwHPQf
e1IjspAZySNGdCLYRCG7YzDyIXiLC9bzCbx7iQqLsRWZjFtoWptRDHHm9h0w9TvX
Fa3QzQePWgUYM2ePsZSibsIa/1isPqvazCfeLeZ0Hiw9fQ6vzbHd9UawiRZx34AQ
AZ4t2QLeMAYJOZSwlWGlOvt5xvxSgMukA0RAnMe6ZNAvAJ0ztXjED0M5S+yZxako
nYO3FRpRqJ27kk/5GmVS1CAJKU+ckMpu7WXsWFjEkspe8tSyGedPD/RMtVGqA/Yb
gL0ttX+zjLDELVbOoQ854LFU++PlFF8aP9YIlvuv0whfolX3AQxXDmJu4pKOgMzD
QJWX7CqWpv56iMFJXIWJs598QctEAVZowrFTaPJM6yQIULQnUGpMQEgCuZC9qu/y
my8AOitbpxk/YT8zzYVb/DTBJT+fQEs3U67eujWg4a0CPyBBmwtZA3QKDuHSIepU
vskVEYHPXP3s63aH/O33MXjkdEk7YOOIOUR9skf6Q4tzofCP6kMiXyVaNOJeRo1T
LlRHZ887FquSRkC0uez4lk7E0fXlxj/c8lWzXvrx8rxRHhy0WjpXW/aVVVG0XhLk
x8JfC+ju5hTaFPg8UrvRQ7BBSSIbZjwlXY5zFEmcwIY6t02f3fs6nKR2odszV8me
WzQHK19YSgi8qVDmfMzoeuypWd7sFX5zTk8xVU/zOBFq3jtXc2TxB6UiKFCbWUId
NwaujDUYVeEK4gjYO7aSj617txoAEv44SskrAuYoXcfUbDumsZRH0bnVSsh6CR9g
WZZ18xtmtE6W/NTKC9Zv9H29IukN49UCNQ6PWaX4+LqgRxDj/Z0VmZFV+LjKZiyE
JfuZC4LIh/xxRFdBh+zp1QBO8oRwIu3W1CFEqSjFW0S/EFL23qaQAoiJM13CdIQR
G+1d17Hd9KTXJTtlWIvQHNcg14OxA+pRH/gkPNJ587oQjvNUjCuV+ilM957ZFQRn
VjjcUkZalr/3uit/o17wU1BuAxf/ntmlBGbFRxpFva15WOJdfXrmueD6OlKgqplP
Cma3UYOuiSebZ7AocXqkk+IHpuj44bZtGcb5VcP9eSaFAYvy4Aiht4CNfRM7uCpK
+Lkb2SVYVBp9e52AJLWj4dsMHVWreLhIc+xYW/x9mQ8qE7l6bEyhSpbdfDjlnxha
Rbbei+h3x1Qf4cFb9NF0rHjordZdecCHiB+Nea3fvtiOSmxr9v5HBZAIozryZcWC
ORjSfmIc4+YDWxpj50LMRLo3sIA+PRKQws0v8QxXEjVn8ti14d1cERYmfBuebGeY
7V163mO4lNfDnoPJDd+oomCqzm4wEBXZ831TVH9I3enTzfwAEZWp8RU0yRwjdchz
eUKHibHCcsXcVH1wJX/u7V5aVS7yN+UubE/0/5s/o+tB3PQde0lTsIHAXGg6Wc10
Zor6/TIPO/DsYW9pqI2H8Y0m2/zpbXKGhCimASVFS7fS/b1nr1w8yjv9p2EteNEs
9vbJHXx6nT428HPeyS7+oZr2fk4R18pWNsuJIgMH4oRZlKPv+766otmZ1rKHEeFm
1DsAvXlu2sUTf4ehf/D+7i+TsUB6LbNIO2FUn3xCwygcb+WZhojCPsivnQJMhoYQ
6jP8uHI7gelP5FFPQ3fyAIquX0MJC355+Qu5LzQ6kS9Gw0RZ6w+ZoNFZYrUf18dz
xCWOqqtlYz2l1AE28sou//6KvKvf8JYRGtfx11oVZPnajS6q3gQlcNPwHmhoVhq+
LQBa/9tWhQWYul3EVw1fhh09SSZuIXgyUFq1jRH9fWSoPrj0ZCCJvF/8cTGsNBnJ
1lrgy4OjMYoHhcTIvwWKsBXxWqr3topManBzOyQEP1gP9SqeHVbL4bav22NZK/Ic
6nP98rc4Z+PPHDz0ASlDQZckFlG9AUzZOmO7iIh6C8nY0PjDewId+a2Mw5puMegE
LAY9PZvzmrPPczKGYoj8FoQ6dWAJUKjTiPeil8QDe0kj9RQnPtPG2LNlll8E2fOo
nBBiB3GCDkhAhyPaVmP7VcpWWGe++zYDz3W9cP+dABxgVwBoQ/UeR3MtH72gPFa2
B5dBK+zx7acBrNtaWZPtCEtLtMFb9uiYsz0Q68qCleEkgJqMJn0911Y5pkBhdtHK
LcNMeSzYwctytWwcRKzpwi7cjfWFQy1gjNjNJ/68eMspMBSI5I2f2yU3isekVqTx
knjBicmJrdRd7gda/VEMhtHMBWEQXsbIuTIK1qX3zLIm+ZfyDFdCeq498WlBJ9CO
SqU2fXIyPE4iN1l7RDqymV46zOT5I3S2xzucoMYOiZuceGb+qejMMIF/2CE53knS
vGsvMpj2RyxMrcX7uOrcwykambnT/csTdga6cH3anXTWth7NRcjOAUsr1QTsnM3o
Z8t6mRiRTBsEl/uhTsIaRFb3UL00+KCUV5fZpnbquWm5PlUJwGigZ0kQjM99x3yn
ewvgHmpn2pewkogBUWcxxDGre8gSqGi5HMUli9LKMtzE8+mEGXQasQPRNuc0L0uW
P527z+XeU4iSZyXaA18QajFumd2EuwupaH7cJgg9HFM0wJJL2Am65Zxu5HfLlQrl
kNRR1zduVqSCtLVwX1psFCnJnG+hk0SbBN5eTbQLT++RxnN5InRJz/GUD0YxB9aq
wpFrhQtDmar0uwqaEu55UI6W/71ijoG6NAOWCI4RaJFb50wv/NgjBvNKrXTKSyZT
9hihs/GItZrmqCZc/ga0K2xAzXiVdib41qHQz8eBQr6Ae8rw/lbu4inl8+t6DZeM
S6TdGBL+bCzFysBDnNWyDCM7PZ8Yzlqn+FCGOdPYsSt9RUS3Dm/jjfKvQT/WL7Zl
B/VXWaVcPBPMhReHgbKjkEIcqou74QKRJJ/7I6w3Cs/jTPo0xh+ESMJGvN+QCRZQ
/bAunNlfdtEeoK/UYiPHq3flZRF/dcksDHNrjYQrrqNHchxiUyl0eZXCWy/C3WxK
o8RHr2ebFUbk57ieVbf3UEjeGte/OVPlvpuKkmAGXwEwPH0hMjiYUvmFjDuN9lk1
MhJeHmUl442ztCEdtxa6iMCLLJKEEwtN8XfZ2tClDBbM0SQkJtvqgMOQ2X3Kr80T
3V/SCZTk4CTDo9M/um5W79lDRvyc4M/Zflv81ELavp4FB0L2iFAOvhkvei2Dtz9s
pt4tddCQt2eBaFl/hFWRKeQLnmlb7hsmcFFjgIKm5YzX5nwCM4wa2XSdtLunxWHY
9+YBhDQcW/qxCDrji0VKN5pL3D15CWnQnosC08ekybTaWCasxSbeRk7Ag3iI5jP4
ogfT1huSoOjfv4TMsu4/+qrWgq0y8POo2EKjwnJr7/Lw3EXLYBshoiCc9XnWXXOG
4azgqvCZohXJhNXPRjNriLTeuLoQ9wEKDzZG385Z90qVgqgRuYCKtmfb6GABArr5
R02mMUz/G7B1m/++XyfyzfpxXmx7TW4bEkUUsrhhi+QdUab0iMAzWWDgRFNmSRmP
MB1CKNCBJsWbQTIuGb5IhyGfVk1CGd3DALI3/3s5OumhFRlERuovkPwLv/dN2gci
aMSQggS7XfA0zmhelWwdy9IY/W8fBPtJg52Es4JrvraViw4HMPffi0ED92lts5F0
Lb0qqyiHwVZrrqrh2OBbpmk8DP0yYvYYI0/mTb+cPztB/IMIAgBSB4Zm8cEI0Pz0
CRmDGWF58b37ygbAaHRpI3Xm2+0uKYSl5rR+AgxXTUfi8dlI/Znu53S2ZsUZO6QV
PB+lOeZBt/yDZScyV6XzX4enEiBrak2PvFhZ1hMXKDoz3eP3WfYRKgqgTxLWeCFu
aGdP4+tCRhgAyrd2tXI4Pj11k3dL8tC4og44Px9VwYvup5qOeyW2DhoN44FJ1S5R
7oyVKyI9RdRQMWRh1t1kJQIZuHQjDZjrAObMmSOohVe82HHjXn6h78sRP5exPEKh
EXV6ySLwdujTtIP12/dkl+YZsc9bAIM7C2GIykcE6ZDTsreEHr79DzyDddg7J4sz
/ClnmP0J6d0YvqScIUjun6+WD5KP1WSpxRsJ3QZeRUtEYwAPtALeYYbMQTLPM0X3
5nf/+ODfoDwwlgMlvgw1GsdH1EBhtP/08f7s2v7PBk+x04xRooSUU0ImO79NgLET
WSW33Hk3rlS8CZni2pz+rNI7CQPSDnWKSlyFcSUb5a99qnelPGvHlv77FyENsY53
zTroogecE6G2qvdvxx9PTt70ttUGT8aSMUNsGSz/sv1hf9WeHnWZdYYbFZJUQ/le
fpT7jymj0RrQHGfoI3ZxJV7Gqw7jqaOP5wNL2GbcxO6x6GEIglPNFWnefHyxyaqh
L61yn9Ui7XxWl5eIHn7UvV8Dwn1tVtdJrO6y/3qa328/gcdM+iJwO+u6zeXa+5DA
gBDxPHeRVPhSPyaZOo/sulrCAJBQrwm9VVfMnHK/zS27tlk2d5zI6jSkyyDnyOAo
rXaWPK8rbuarhXTqvraYGpoE9qOlikgFIh1WxCVyLmWd8F4UmtDZvOM4Yyi48UM+
MXuC/U8HROc4lFSIYTTpP45cdjVE2SpbaWaEB1kTOFufxYowC4gzoVuwJJTkCbSF
5ZK+aJUz7QvSckDkZLMjHXF3wqqjScByuYo0vNcuC4kWkD3PEC4FbOZgrM01AoWL
HvBN1yyLLpAWfhjhBTMgSKXEjSBwUbZgh/1/FGhniokVovQloPgmcuePlE9t/IOi
Du7fBSFeipDX4gan8JkmwW2ygG4AMG44opGCPz3dwRhdS67SzbnylCQum4sQ1Frh
UL0jwWsWLrYL7uXASoY52cxNP125+tcgBTocJCV7NIBes4Q21+aXrbetp5snnej2
2mefh7bQ9xhtZ1M/gJ+OJGsXsRh3gfdTkDUPC+UwQb9qNZ5s2ryn360v9bjw/ny3
Kje7YH8LroJtPGot7Y7IniwawHbz35vl2NX7w6S1OVCmTKEadHnxmFswoDaoLGqU
yz7UsyNUMwBDUa1KlFe2xAHuT3c2jLbBjJSIZOGpaKzioIE4cvxtLK+O4vawbR8q
yHTRAGZFiKU3xhryLQrDnXie03RigsQRj0nGsmZC5eM2MrXx1yzYzAPdIWt2lLm/
u4oofdEzHNTpToM5rMluYV7r/eR+iNdHmKymntFizgenSxD+8kra6phs5EzBPDZl
L2EoYgPqxwR1H8VoTUMJ0AqNRXadIH54XmvGHK2BnmH7SSmdZEM0UUkyKr9QwD4h
H4TwevVi++diU7rhPF/AV0qsscPybySmARHt3L7A8YA4uoxanOZqy0hw2G1CLNPL
3IqPt6T3y7paFQ3Oj9O+b4E30QlVPrujzDrdrASvbzmHr/4Wb2eh2Uy+eBLpeFO1
7+tAigobUO5v21iC5nk8iJ2+SNegSfn1364EOfPC/2HbfSPkcL+aZPbee/C01ezu
3xmVkOvRE8cZ8qIPdm0E2IK82x33MgFAWnPTdyzamkPi6a0V8SL8iL07h73CS7Yx
rHeRfYUeEduLYlbPgPKsXsRjTzPiHHPLzlRRqQIixzlyUBlHQZjpsT56FEuy+GeC
z5Bfy8LpKNd37uswJTXplzA+l0JR5xmcxupFO7sJpSf9tpCplp4VM6yvpj+YSXFn
aftriP7XmI9Y4Qb1ObX9HVfmQCDJ5xIQdVH+kf5TRk/HCxrmtPGSxEvOCQQystSE
zJIIDeafOx1laSjrWg2wumCvKCck2b2opRQwbvgWOLdI37Y3NGeQ/luk9cxcWRkT
JanCjnEIsxhuVrsHlfPHpxvcaw+Gl97v6J0HdAMFgi3tV8mpFAr8UROhLrs/2nds
GHa6IXKEO+9PYFxRPRUXcMkAftIwzvwAbhC7gHGwMGLdoYPFU7DZ+sEE7+WNtsG8
dnAu7QomI5Oq3EXWKzcyr+pZMUSrv5giSkChLK8pl7017eZW9XQM9PsD70YhLaSo
t9WU1Sd2mnHi8AqC4cOS8fsSE126JOVBzHQYXKwqjhh/nT2vjty1IbhB7HCpBR7y
EOINJifmQkU9i8dy/BfNBwVQdi2l7vxKx6Q5SFFLW41FwjaW42Yn4TNAcDMMbaiL
VtHLsPkgqs8acFJ/GewRn9N5gspKQorMqOPuGpLV03rg9wXY5axZRLflk/xAEyrF
jQpzV2MZP3W6S9SKRs1WRRm29r4cqxQnA011sWqu271IRAO6L3vR/+X9kFb29yYi
NGleFZk/5+tT08a0clN1jvp6WiHLT8YuTD2IPJe8wYbBi3Ev5XJkL0ZU0+Wx+wjU
h3nfa9jnxHtBpkHZwnA+Iumc+LwkaF2LYKrl3/2prmg/sq0rjqMT1HybHdNU+vhz
bHUNCWrfQMZeKn9rZMnBKuJqC+Y06O+vUe+zDVb9Vn6JkZ+4OuHNLGMFXteN9VQv
zdX+QFFa9BhDPCrn4HYqGQGM1uyauFRQQzXDtqHjf+Vph2M2HyqJYiNn6GNUGaXR
BoE/40hJEdINz4aNg6j/1xrsljw3v04VekkmhqDd/JdKXNg0SbOVESi8w/TGxjL0
cVUUZwN9YcVCk2dvnxVXbAo/Y5gR5K8n9jq059gZALkV0eUf8xuEOM66jv0CktQF
iYftLYzMeeYgxtmZ8QK+hL53+tv1rfig+m2NXrt+VPsVTG6GO+rAwgfCztSBnTje
D8xHGDraT0ZqG3u1AsMflPtRhiJAo9HNNUSY0HaA4XIA8Ahz8vAyVaVYF2EFnqhs
UIcBm3V8ua0lsF2KMM4YAMJCQbOY7ijLjKdVoGqyjVdUG0FcAYsogNC/RCJtb3Sz
OOoN5wRQH9yXLCL2epuVx4s2hY1CghXnAn84ueDm6HMoUY7zEEmwoZEIT0/k0tk5
sNwG+12dTJAZbIHSAuqwKbzoiHZZSlriQQhai3DPabDh5xXa/wQm73wa262ga/Zq
EDaKC1G+N5gcRdYnAwnfXORl47glegl89VoX2l8Aa8/3kF4xXGi1cNmwAcCLDtJH
vRogendHVbNkcGSaxxNNlE5HYfwGyx57gg+iaNpXn8NEMUkge0jToZ85kuJU1d/L
0LjJPJH3NndVTh65vwpyuBJZYy9URTCeU2rEVW60ze74i0XT3eZCg/BLqMP5KmIX
icbN5Yc1nnX5qzu3rSqVUpYXvlurXYIT+/4y+22xBe75Cz8gxcH6oxceiYaZAMBa
tWzAIqBS/2GwIUIZLzPKNUMn99VBSWrJubviQj8ek6QbAQ/N+hKflTWM6AAyyTfC
+krr9OWkm9MocnLBlaY+oHXuPmfHv667V7ejxKVTLGC3rrmMHjAg8pis7MzRtwZW
4EB8BNiV5To/w790Ad5K7oMWFg5peB8LwgMUZiGC2BH+SKlgdoBfHI/GvL0D2fuh
jG/YEF2VuAs0EbygZwbpjypdy9/xyh4kP+J73VyV8l8HYbEBBjaYBclhy5s1Bw0X
G3UdFdsyV07wRCcnHfnIkl7dgJvVTW7Tln2Wx+T4iTzD6Ejcs+Cio7q4migxFePA
/67Qgafc/3gFaah6KWzy9q2TVJyrlMRwTETNfvCfbdSaLhaYBnENZ5lFhQq2Gxq2
ZT5xGZ5/9anm4pNJSr1ROmPp1B1QeF8K/AAws7yCqeyK+gQWe5gSPOVxGJXh7Wqj
LSTccwi+a9finUO3AsSItt/7Rv/SZ5H5D6PtTUBXtGV+R6v0a6znXeo+0bGZUv+F
N7ukw9eLpe+Cd/AGu6llnryxFGIk/IdeFX5rTRsCFc4gIQyNRnuHNwe68eAcPJxT
Za/3maIiser4DawZdU399ItFLw2Gvustf6IhUNu2twx2bv3pJGMhcN/zMyO0tfCr
BfA1Gi6hvQOkUVJWqSw2hZHOQw2nYwL1HP4FOQulZfOOndRoMgCn264A3jDOG9NC
eRxfdEbJmO/+mn+U1Olu4aeweJDBnAEObr+l2X9elzNRBBt0m6Cr/aCpjN49ajzz
Ohsi58WD60q85DyGmwDhuCcYoHA26Y3g9eGJf8XtvJn9lzCW0uu8cKXD2FbvL5GE
Zq37P1F31ld3mOa0E8LY4421BVYcGh55ImHOmNR34+q0p2IOWsTNNWQTo78tj6hI
TKXMrmRjPj79FqSjQPJmurLlRYmnjUapvxCb6WH1OAdBl5PjvKMvQPoEOx3Dl+Gr
iiK+53V2GNNGkxNWjY8P99BOjJ99qd+mJmiY9dsMhRBma/3q5KPy90RF+8uQ/UgO
kh+QczTocsvhRM0DejlBpb3+ltF8X/F63V41ftWqBV33WRJc6H38qwDnLz3Z6FHF
w8AbwVq41FN5RTOqNQDfiZZNqTiGd4N7NJRkEg5xkZt4kqGjubWndwPn8E8AHIuE
lb+xt/lVxSv+i79vL460A9sv3z+DsPE2or9n7GrBa9pQ0nreH4D76e+ohpfJu7u8
msArNu7xOR1DYv5hAD9E/KGUwPaypi5wnz0McZxgnL/BtRJQTTwlhe+bVdxMf0B5
AOCI3KfXtxw4qZgjdmcKI6jfSOX4qGMahuqIF9lxQ5aQ/edBm2n7z9Byj9HwbSI9
Rpmr2zKtR0Icq3R9I1rA2Gjt/rYtyIIREOl+xbCKpfxf1a/Shdl3lJSioLZN/Ui/
cMx3QR8LgzipkVF/xci9OBLeVyhIJq+yZ9MvXb72iQWD6WW0OR/iAwU+FBK+3SN2
KprfdoPnbVpLaZAq158dCn4cekO9VXAJrRd2EoUZI/cL2ieqjMQTaZAL0Jtyw6F1
Cpmq7DY8XK/xmOW63CW19LBsr41yJyfOacI81YcuiJptZUgOFoFF8RgCmGA13yOk
HZ+aCFkb+coOwGTxQq9kiT0ArvzGGWwrVd+FyF495K54LX7lZXJzRPDXuHUf0oR9
Df2fs8sed6dAXr1NU8zX1lBaQEU78TzY1L73K5WIf0iLdQSKnxhbGZvz85nLdulv
YLZBIsIXn2blK1QqCpXH7my0W+wJ19lAJLkC1JjPysHjpo0pNMzH4GuH9I2Z3HBp
z84TPfZdQRRPYVVj5xxxhiClQSmvabgyBSmWjl68T6zdnIuRBvY63DvUP4Acq9kv
4dMm4T8CUqgYoaha4nb9h/8eDO03aBd/6l9CSCMJXu5TzCPHZYoE4QUQj8m3Lwl0
sGM3x8FjqbIjrahnPtYFBqNQO3tvaNgMzi708lDXteIBpKN4Q7sdfmYoFE44xU3C
bFHQisfix0dSVNnvcyyoLpklZMnHP0epVhrvuLMMyNxfiQ6KiUNJdh5KwDVzVELn
BGSYBcj90eGRvbxvVpVPcWKA3NJhcpeR8EAgsXSIeqp8eaBrHMhIaJ7XZ91YN3bb
zQA0Frk8fmRRYbGWaRn5GAsDnjrjqClryDTdHFbbKU8BZW1gUQSnktWg+okbb04O
4EKR+loL6G+SC9054n5bljwodoTQzWggbRg6zkOhIxGhmnRtcmKuGFYdemQQc8t8
U6WbIR3oMvXSc3rzHZjXEwxVR22pwU52XKjgNsPJq1eN3dFupy+uSa/74w+Y0Us1
3sYj8EBKWgm/B9T5BP7e06C8cHzFsVKoQBNyOARnk7mGBjNbckqpRtSFhFFXU61y
SeVgFleEdNYHXdwMn/kSpnlnWxFDYoWoqM//mBBN4cx1XhEvmWLvjxl7w24dGxNA
+o2+8eZ4peqNGIbY25jVt6iX90wn2Zo3cuSvnApc5+abbo/O9gsUMyfOdgOQAbpm
0Rn81LDLb50mrjkQLaszqQEbv7QfM4aARZ8jdgt2f4w48pFDyjGsOzEzcAR5iFtK
1L7Sv+GfPIbCJnE87ORUeG14ci3Bmd9OzE5vUbFoLMUvSSEDLCO5v7obT2aI7PBY
bzyXTbQsIUVLHjUxyz2bGJ4eURkHV81i6hmkn07zoHsZTgN7TdvOQVkpNA50r6ot
8MwTDHic26532Id0aISa5KnfFw5GSqyu02QmtW1cGkD8JFofLo3G7oCKi78TJqdt
+i6PetSUx3XrsYnY65v50T4GlqvVw4u54JrYPMNqgE4BLaePSXsSDx5ZLGcDn78E
NQQjSV4j7qjvuQJVFs9bZ9HhtFN8kB1t+hkjToSCyyv7xnB0UlqrhKVOcAuAUNCt
GYiNHz3/j36j4mWOTU/0zZi9WXjkwrs0Gee/M4QNGHstUFzzKnUZG/EB7Tl4Im7f
LcLhGqkaWa/7/tzypdXobqYmIM2UwgoFdC2iAhYPW21Pht4JyYTSheHwtdAVog5z
CvRG+2+fPk3JaeWxCuMUuG9mLbKVLrklbB6KWs5DOGctiDsIz/5m7tc2x8ZDQ+Zv
davukyP128gL7YCqgdgmevEQwKZsjHB3bq0SY1KzqUFK4uAFi3jtgSqtdG4qizzT
7cqP5W5J7p1z5AoJDUQrwnlL5yi+RWikpQI8Z2EXSU5eJdQBv0HsEA2Sh8vpEvy9
QODCJbpWhK3qpArtY/03NyIu8AqRCsiGrhIB+HqIGzfPfa5Mr/BT/CPo6EqpSckS
hA4aEEry3//Tmr1dm4W/HyxcAnioukugujiwKs724LEsveD7Jb56q9jXox/9Y3bE
5s/7CGP/QG7/1xEAtbE6V7rb2NgJtej00f4ZsNkHiCbUaWqOo5QzaBxR0KzHqW4Y
vyGQ/Se+YqiqxeUhaWqBkkqycYoIO1ijQx56G+KAkuyLrTTfL1BSYYiHuDHP0C1c
8vlLrkw+P4K9e8IP7QykYs/Sh2IcLiVYLPD0xcZ0wRmDfe/kSFIqyccKqJYXr0x9
AD5dcaQdmuShTYmJZWBZeaHOGfXqpccRXi3PsFZoMgh/bUGMmkK+24y5aezGggpz
SWFiBQHw25jBkkGI7hZSoxFhIyBtcvzgMgc7shIEVeUrBNSFQyxUzd3HFSBOqj4K
fIfuUx3Gm6rbCR/9myGl8+w3ApNaZ9TiqYthaf+8IYLFMm3JcI525GkjW6RRCVf+
0450NFibm9dSn808JEcHap7QciA3m4sBwbPVeLMg27HsaBjqkeUCAb9tX1pCRvhl
piZdG1wQWcXOG3LRl2xUQqTHA72UvQQAgxUiojRPkIt7S7mY5jkFwdD8M6TSIuci
/Wco0rndRMjQbpOcoOF8oIy4XSgP9FTCShBgVHQus5nG7l/Wf9Gzha+bzStCzjan
v1W0gVPd7PF5ODNxcY7nqhdslM8w5aHHt813snYKrwrzBla8sYeHQ1LhnjCKQfyG
AAzmpdN3x86WHkhZWNZJIz9oNBcayxU3vHcDI3vJvzTui7Ag+RsHXs7EXqCQASdL
u/WQilu6+wMFDgWz8aMEECuig7Dq7hoXsjKInnPUR0vaXtCEpPNZkWGBbVyisS8I
xbQAN5GMyFyfjiM/q2a8UDo5oAdGxvmt6w0/dR2l0ohGTgK0jYsPxyq7BuTxkj4Y
zN2tBSb3AvihHzdwznTLBjDsE53kq0+EhxoNj/NLB6lK+6KXo9Ck6NgTu8Z3B7Gc
Z1B98mDqbR1QaiO2rnJ9E1RZ0UaejYFrshC+hxynpEXC63CY3nIN9LcCG/T/Ov8+
FpJw6X8jLPtxm6KFbzTu4bzGoYW1HTQP/nkawzbJc3lrtQBy78OGT7Yk2Bum/u4Q
Fs83M8U0W04PSqWP3CoQ2jmHqi2zwGV3mwv3tpjbD+Ve0UsIHIoxDBV7hgcb8dsk
zXltwCb9zQQncK7Jh0EBWMkCFaoRxofr9BFzOpSgRUJWinBL2Rr04NO2Y83DvaAd
c9KBHDbyrzr3J0FHImQ3VD0Fe3K+NRli9KVP7cXxghDYj9lBsu1jkjKuR/gRD2/e
ATKAsf45/U1KPLFoOx4tgN5CRf5iR0l+pUF0cxZr/b7XWmAjY/jzOP79eIsVHrYY
CFNxXC0ajb7Uu8IcbCgrSrBm9OQjAnEtfoAZE9T7U9leDu7AhwZUIfM+CnZQvdYG
6A5pOR8O65WpEdMb6M4zCvSMXV7Sq8qLAYzZpwkygKJ2Z+TRyw6RlFJmpOxE0nia
qzQa2wyFFUnSQcI7GapdeyFPV7kZuIbEpoZs2MRrQVod622YR3fX5gDrciWb/kT6
m0cWvsJ4+SXbnoN3TtW60h/XkOBiJgXcUz5Ca6gTP07Wd3nP8VHqZuV5xNNMIL0x
5paUNZKZgP34rYcIlapJMGC0lpCSbZpr0Dn5G60F+MPHF4hTJUN8dnDjgoDGa3bM
5eE5vsMkwuPn0ZD0qqSx17zlfmuuPK2OVDwcAC5OXCoGIdPO7gwsSNlpYbjHCNH3
oCP2hzO2YEwGdBP3NE2NtbyfNNWUefcch76mVOonEguaRxJhyRDeQhy7oK2/u/gf
sP3KISDuN/nFcPkc82+0VhYi3sumun3BRmoGb1yKYdn3/4wyDxD5GYZDMY/IAn5D
cL1UPIwbI5hsQuFEqV1m4wvFZYOGYCwgTqizwzvgzNWxkPxvcBLt3d61AZX2y0E8
iMkUwgNkgDyZ5wDngeTALot1QmXeaM8+9C3+c8SN3RTnsM3C9EJ2z6NwZphCD8oV
ETkReBhXZlKKgf6cKF1f0FbwlmfWgMmdtiJ41WY+H3Q85f+BT4lWmO/1udOzzcLQ
qrAjOAWiZgQ/lgCOA+5HbUwO1tYVSVpp2gtR6zoE80VUHtUOEAiKkg1hvdCiw6Bw
mFKz8ee97ZDiR3/S0iHFAFNMNY24Kq3QZGpKc6CFzeunJsVi7M+w4NjmPYyLBAVF
wG9yb5IpPy6G8SpgbOr7g8LVZIJvuEsS/6BW7BExp7m4jiMS9w0xPoBDLdOrufnG
y41NpgDJp0YlgAK3no17dg1cXEafbsaJsKzI6xe8LrwGMVdhfoBDtj39/IbpN4gv
lkvsWpWxbgBVogFMEoAf37Fsb3PHc8xbHstFSvhbge+mlFPo9p5f7zIPITnYaiOp
cnh9rBmZqweJHsguuBCeGAU9iZ0Frt2tOK7Fg5II4jL2exe3Qxyi8aFeKkTXHUEb
r+P8XCITV+uujQ9zB+Pfuv1878BjSQ7k4w2hh3B3mD+LwIWCQ08/cmjzmbyOhNQp
smCDAkR9agSePQPs3B9kagUevYPOJDy+Tp9PdIij6XZkk8N/87N3K0LdB3Imvek5
i0K5j/SBdHC3+srNUrAK2MX5DvxfK/LzU9tNO/T4GZzwqVoCgEKqcu9pIIMJyTAP
ZKgrnDKa1AVBN85kcTaicFhejrwenBwObsNf0TFGmyJaa6fEndNKg/sh7HEORQEX
LdLKv931crvuOWxltmWj4YiN2QA9tC3EVQ63B+91lfJVesXWF25euhTf2Ryq1XDZ
txvUd9anD435d8HogXju7FWAOmt48CXIa3jev0e6rERAV36me33tAEmNbo1aQAIy
ySjlyMmVBq+e5khVXG0BVhkISdK+gAykQCMNFjAx63XRiYnT+eBl975KZNgBA/WH
Zv9TvOOx79ya2NDzyqik2hI1/TUpCOD41V5vs/Sgv9Y0uquwUZQgqhfvrVrxLjPx
ECGjAduVNNQfNXiNEbWY8mrX2TRXtwGhIhU/GWwLZFX1NAOiC+llndw39Lam0iLt
rfhShw66mwOZbL7hUrBSfPhQK2bt3gAop1ZokwTuQssoahRZYxM/iA1gYAL4NB9h
/Rcx1nKAFo1SC6u7keweqwjINpjeUH8ni1VMY4DOiwv5Gg/HqlkjL3SWcOzXyeiI
Cwk3qPHD5Ku5ShpsqL0z964Z5S91eWOCz8zSI/i4sXU/Be4cXSmhuT8apo0zEjyo
Nh1qdEnZerzv7HET0uzeFWkpzB5hT+ThmvXZDqdBKIFBuiy1RwqxEcrtIi4UCmuv
wAgLxIQancjokeAAnuBrefWI0tS6bS4X1YFgsKCeQPCJoNwL/7xIyCpEfP0Os79v
DimFOOLSivmg7qD4ZRcBE/myWTusVbhTl5yzjCHyBxQpDAkFgh1aGuPM5zUF6Gyj
FYWVmk6jvtZEmb0ImWWI4qeZR5qkQhVaP1SnfwaUnIpnOiDWbLogjLE1WyqqU5CL
ZsZju7A+sE6PUdjsZ9Q74OtoFz7APJVyp3cBGkWh0XVT7qZtXi+y06uS4sBStf2U
ESNF0sk0qXIwQeFMbIZZvdw8vMAhSsLpNPHmR1vjfKAg1cI4pWaW9CgcdgEjVRnu
HB5C/+/wpuZse+PCWKi0brbUQJOZ+QGBx/4TXS23mg+jsyJEh8Uye9Xd7/9a9DyD
x4+soMixEiNezKjrtntETmZOxLGbQzJ3YfnnF+hzNSB14qDTr4D0pWfmIbZInqk6
3oUheetGf01gaBizwnOpUKQzbxn88Ch9v4njDE62FTOayLIs0/sXVMC6kGMVxoEy
jnEIF9ExK5Ps7fkXUWoVPkhwXoSXvqSSH5HDgWeEv3uDsFzdqZcifqIOcwMsq6Gz
JyqnSLCw3qZMiPra7rHwyJPLUoHfwB6FMMA0MA0E97R3+lckE022hoVjlNyZvugU
k1SZ01Yk1iC6mlV0A+a+OucraUMoZdM2EMFjn8cN9msJFPMRQIhrToqaZu8eBLXI
bOPLRb/H8mzqFHq/6tCerPcci7oYcGA/g5u6aNx9tgmsHrIGvB4KAzjjJdZa1mTd
4KIWOiaTtlXnbXDMzgJE/nXyYWVPD/doTpzGnXN6B+Wr9p24+NddHX4zTwwjk1iE
Uk/5CZs6TXr6DUTqM72PdAhwmu7XEfvvqT+A+/LXzXt4s6YrMpu0FTJt/Gt/f9VT
wnr7JAZu7HtEfAcusk+A4h6CyJ5SNeo5Sxl33lqHIPIAew6CcTbWhEOgWG6G0Zr3
vsVJuUbikVfZP01q7kolcNB1K9SfHCBJ8/ZorwBXmf/7Y4mNxkf3aeiK4nBBD4s7
GNkO8jijqmrF37u8r4z/0BTrwb+Z7s1c+sn18vDlnPZzNiGpOozOJ/nEnjKjEyfc
dcgMDqFVUzLTDH/+dYGS33VBIzmhzqFIHbQOaoljaA9lmtZOcyZJaljPkA7Ui1w2
vgWA1Xp4xmbKM54FPPc3JOBuVBoX7M0I/fN/+bMdtMwaDoqTGTZoOigb99REZj4j
M+3v/mY9/6Bj9t2hOC5X4XjTaS1cx4K6C7aKNgDWtVNU0X+d/Ajg23wR2qWyZ38X
2nMBuUvOgeW+OQB6hibCR0FEw17gnJAqWFgEHslunY5trbhibmDVPXbkQiYp3xne
aYc5unZ4YWvkQn1wskTD6cRpTGKmy8r5WgXcvclW6RzrSuTCBRw3/nWajyJjBTCY
xqoElmjGOFQ0H7xv/A/VtPjpDT7mMXy1JnQMwp8OTI180BWvWGoYgArxtkv/pfhg
kedIFmki24NSHe9DNnFCuPerEDGmfU2ko3Xq+KdWdHHmeKl+XsBcL1u+5JDqJrXF
kuufGhP5AdjOjyvmRJhUpCn5wd5wsmwmF03AegY90kLph2GVsr1SK0+RK1aNHRR8
MUXNp4y5zd0ogEOukoXxI4Dj76aXI5qb7K9u3PQ7Wc/aQRIBmvA18xPMC1LmsGc+
5Ljr9ra9mWfydBIeqzpHmk/JOFALzX3vdzj1kkolLphtKHDr1yLNFbiB8HPpEin9
YwFVz3y/UshBBv8M4loqtZNHJb1E5nRbaXz+6b0HTitlpRVEa+nRn3p+XgEs7trp
F+jN2uYNt06PU1MoRHxh5A1lbY2hAUP8iijMLpHElRjc/KdrQVH5IISS7QOJbIer
ws+0tEZSpIZu5uZukpCQ58Pqyg4SwQc+hl1yUyPSzCDqhrmTmSfxK5DHTAFE/BEa
/K4Ilv4zjGV70nKx83iJjSmuSYTbZ8hmp16DkmBh9IUFbpA3LMquYM+HoUpEcu+A
5NMtpmvOA2Ym7bfrC+5VkQSK6LvPE5JXJzScN16OoYpl4LcRopwoqrXwL+s7CFev
q767sA3sZ2smhHElgKPdGia1M/KFAmw6CZTmk7U1xlImDuIVLl0LMYVtBUX9b22d
Yh1+uXMnZb1qsaXud6/zIDGS4MATH2R2voVvDXRWcQmy+gmLUdsGgfJ+Rduvwlro
1ya5TLzumpbt1VZgmmc/+QaEqnWuUvtBtwCzXtFGxdWd6KM+0HHk4S7P38t9EHOp
IBE0ZDr2Poj6oUFC4zHH4VNlt3KdsxLaKY0WSg1uZ3QTEdE4E1MSALkhauxc73nD
Xo+n+hdLZFclfn6E2NN/kkIM/YnYBitUIBH2+hI9iDgnHXh7qA446e1TOb/O9fbw
KQd6zKkOT74jxYdshXJW3U+716Uww9IHvKP7vldjQB9WOTBMoyouS3JuUXTeifbT
50bJ2N3baIxsije9UGhDsa3KVOTd+HU+o3Y2TGJ7H8hkOGoJM3qOvTdRW7EdSExw
daGHK6EveRM4KyUZZoD/b7lYwQ3fqpXm2DCmLO2/HIrTdGKp2C1G5iUlNVsmzanw
Eu9/nTRD6Q5+l/HrT6ayD7NIwBUgpHFJMz5ASd7YXYy6TS/uFmXDI1kmWxT9Gq7q
aCk9qdi/fdjb9v8Ck9xsoKKc5rMTwebJ/HjMMNpybWYHXkf2Q3P95EDVSFYByhqk
GkzwPnlrRX6eTflW1RhoFVxelcXNO9gtlmh1wILgLtkeEUNoLUL+/uQfjYoGjtlG
FZ5sNCiqX7MwhPgFtj9MzetRWC2234KBtYFgFyJ3FXAl8rKETzMoJA1cmmSpYbab
hkiMriohklyQfVYnZILA5Q6ssY0NCPlhhyBeI+UEu4oBp2+u+17dl8lS9GWH1c1l
IIZkliXhAK+dtIBv5AypSYZYQZZv6gJ26pzEin4IkchaybmrUKl0ZtfY405y+H5q
TJHUTgMvHh6F304ps+x7yza6NNHJhOAO0LOA18O5+it/j6wJdBpSq7RA/tc+RDBb
NY+Wh7kn4wFccXDdOuo4kP51b5YqfzYVN4N0PPHMSPsBvmRzHMJpWXIVT5sD1A1t
xS22DhBEMk8vdO2R/hjbcX9lFj1NkeJ1L1dmBPHl5lDto4Tkeioer/gXCjeMeCOo
JNWPigU4drrNJLTTWlffN138L7GCoEP43zOVi1kU9/pcLqMpFopNMwxvTJGYLVJ3
KPj585NuFvcss2YI8o//muJJ4G6G+tVBsAFqQmpHOKaWL5DgLksSVQwuKvVZtIZB
+m63M5cOy4RJtUeq1AdhtGGApnoVvcNF9G0d4HtZfijfdBWisUNmoNQp6+adwCXr
BqqGBkeepeUa/ThsZDfNtq2zRteHBJrSxGrEgrlLbspXhas97s3D6gXG/XytroWy
XdxzqSqvbWuFB8+ntIAXEgvlf3Zk4DsQjmpngeklnOZDli1XlOvaluz6bpGznTo0
KCG5vBQcbArO4GOD509esPixwS5eHiDu5eU8UOavjenXayC6xMBQ/ZokDvM3B75T
6i29BFSSx916/6Yiljm6nZdn5UPeiUqQhz+eg/AC+kY6D6Ti80JyFx4x14hs/MGh
rvyFJKzxQ497zjcxY5al9G/7y4nJwiU73Yk87ynyf7BeYSdg0GauexPOyHtYSaJx
LfcdM6bOhvB/PMddF7nvcKRs8ZQ6Akp6M0d5hsbOoFzkdikz/FnB3LWJIRHGIgEQ
QoSQVEgS5X8wXmkQZebEKRHdYbGyoGDLY7TXEDXJzuY0Vbre2iFpYAsfBQAjoPvS
NrXPUOHCv3BshjBa9UoAVQiLLpK8wVT6pRji9etATdCqP2iS25DBIhtUiut6ne4v
lhGwwc4kBNbF6mvUN/gdtEylPMChR6yaUQnXawMm1w1RylxuP3iN8pYrhwTJNHFQ
5k1qyHsLjzNwh/Jb2wVQ3pMoslGKAlzM3G51T9TlkvNd0+vNmGjigyLgGDpy9Lc/
LAtVKmEPFwt4JxfVlnQacymZmGHZh4l+XyRYP2CfrbAQ1ZNeskxgpE92o4rmG719
rcsoMVDAgnFb9GLdhO/qYv4i3ydYTKfLYh8l/ixM0u7VYJw9EXsP85eaXMESyNCp
NXTjlac5ggjUjmfeIOfA0F0XS8gxC4ALZcKcDbaqIBXc63EC20MgVKrAvzUIyMWj
zAaCdzr9Clsf5EVLF632DvkOoQ0DE/0yTdbWbRPEe2TonsYAn19sFbWtPvPVNoHj
dG2fkD3WLqUmjNYTYajZuN88+QyurvJ1zgbSohjI4ilK7crzSb2Lok+kDeaJsDpV
PM+taHDe6Geq7ueoYmRe0ANFyw3gmDh0L95jBRu2fubgCSoG52LUeR/kw5ZNh4Zi
l4ovz+Y/LWxd1/LuR7Lq2TbTAWRrNBHZNKL+tAFtOL7csP3MD4RCP/cSRrHqz0cw
17KIltgni49Akt1n7CVSQ55oDC4sMniQ7Uf+bpQ3NjgUZvkJ/a0vtM04Bfko6AsZ
/Upp3hEY52xK8/OXEsqTivh9utvM1RX/JS48a2HuAQ5e6JMOEvji+HtzaT5pYie6
FIFRGhznH+4BcyoovIY3XFBoEVhO+uQvs3+NHoPR6SpzAgvg2iYekFpCcDTqoXyh
tLz/7vTn0s34TC14dTDQTR1UgWadyepdGCRInC13lXhS4uW9+7zeVplyCwAw5YZD
uaAGqFj5e/chL/Ovzi8ohCsZAa2wNt9sv7D3SdqkKowU9zrC+sBkScc2yR/xxwFp
PQ0QsdniUWVVeBTMFgeIIjrRDGswkrH5eo2Lm7GUdxSoL1E1Gwaj4U2GjfeBH9UM
euX69ji0LFkyxgcAg8lcca8v805HDU2uyySpMkKzQoqE/qYK4g6V3W9ewH2/tXGO
ZS2iF9WzAFnKNSVwfvOljPZ0aaWGR89WLgSgzd6Eagp/OXZEOFo20i+9WgVxzwjg
wm+kBDuyW+Xk0w2sNLeS6lxAuzhNNSsjLKQ1/3Zb2zGU+I8wp1+LP4mbZ07m5t8W
ZQYCIAyzSh++v9nSvQ4ea/D6e5g39wWh5itrxpUp2ZfvBXaTk6zUPFayiDyMFE0O
N9FASbN4/8z8VAZsHxMb/o1BdfDBCdp/XG23zSNZP0NBcwEw4CtLFwv2GBGu/C6k
3hwUYjgdeH8sXwX62kxBgNeAts1FzOL4upK+gmJVa5CPa9hwjiehqcydbnv5Vsv5
/dppK6WjTbfzc5HXkMqJP44XlasMy5ojX6pAo2Xhqj6ccxbNvdb3dvgY8Hu9FpMm
lw4vbHf5Gv5TON1Nq9Iub7mCmeQNgJR0K4hsMLYxfQUzLSHK6qJSxnIHSOLIg1eI
q28JapNy9vX+Nd4j7EBZJrKTO3Rz6qLnqEW+dkOtOhz/myFcVUC3/9gMG7OpggXw
cOuOmhCyawXdfn3mBf5Aigvclnw80sS24Wg6+6A+n03QrUfTx1VlEuBjRtNiWd73
NsOXdVPVLwtpnMYDSceKKffLTskok//xjTaEEd6zf36k14Vdibeci6eiQTaU+9n/
uBYCCJXUCTIbamDx1dXyBVmVNiksheGwIO+v8VfTTL7B1DS+Buj5+vY8vlgVVtV5
KdJhPeml9YPoZvg5U4vByZHD83DQRS4vUl/xbYcAXRxU3GdffrYqQbtO6Qdd6EPV
gxU3Mc23LbKJ3tf7xC963LvuFj2Wwji3SUrbt8Cv1s/KybBOaJMV+HuMtu9NLyfZ
5MEmM2xmZElIiU9mopLBHh101hlBM0IuBupmz+SRWWhD75cdoH/PaqD2xYCQmOje
hhRPE1qEnY5m7J6OM2OlqOTRknZaT0EQkS27f8XNPta+Smu67Sdp8R+uy5Wl5PA0
zEgw0dCvmTMOklxG23uiwiiWfZ5e6T2z5OXUCqAiD9pySWpSmWk+jubAjc+RN51x
yXH9UooBmqnghQDgEDXQuofISKRic0hGy/cN+otGo90p248An1cRstf0Oq4SO4s7
9qwwqVM0fIoUmE/eEVI+/cC7BcrlD1H7C6Fnunp7Kwlk7YJgrlftuaMG1lwmpA9L
QJGwoE2vSwnqEyCsKI+X5qRnfbYJEll/3X8G+VO0vgQLp8NNHk7AB1TYjsHqQVLB
SjghBG/SUFv0Zv1HxqrPjqRsGWVKa19UK9TdY2trxrxWUovJPrboYuuWz8Z84/xs
qrVErCWkA3TmFRkwaLH5SFXSvesWHGTt6qUaiBwW+iTb1473N/8OSIj5JxUQYpXe
ogqPW5TxxXOmaPCU4Ph0MLZ3M1AQZz/BGehomwE5hTwF3G1BwudOMIBKsx7ss8BT
I+C4Tq5pUA9kYazhK0EITuvI4hQmJQ8paJqGBvOeHEtzIQVsRJfjBIKYvu+iFkBY
uuuGFrIbwkEtV6hRDjdGPGbZcRLI67e/TwQawUendGF88/latzOqUNWUpBlt4Kg2
RGqf3kNpMoZ349GQvblagHAA+Xn+RHro/u9jYXB/RDQSjqTJ0m+jSPu1AKgebraf
4y7Qy1eAsgH3Cu/mNzn4Lrd1/lnF0bgC17lKyEtWJ836W4l0J/qICCZ9WPfszybM
mu1BneiyuB+jgEYGsFiS1odU8Iyfm2yvfjzow/XCcJRbxrstYon7ITl6P3xjPXqM
7optQlQYipiP4lGKbwq27fBbfg1eCCNDuQ04gvYi7rrY1fMHiAMphDoO+t2Fxbnp
/r6uolI1cgLI+9Q7/J6ADXwRmA6poDp9PeO/xqJOhRCSiwa0r/iMHq5VcKuPK5fZ
j5aHFuqWGvZ6951h2T/6JAaOEQEyIVuKalVqWMwihpsLQ7dxOkbBRBbkn3s2QUlA
myWfCuK34qeZ+nfD4n/JvprU5MLWSLXWbq1Xz15cFiE5ZzWA3nr0WQPQqkBQpmZX
x3sjfClB7JPU7o9jHBMU0UVMHn88uWF1Z282q1k9zOcRiAduuDafpwB0JJfFcxuw
QufNEa9wccnLGfZn2gQHSjwWdha4r/1MneHJM9gBBDT99+45dEnhJOMcQBK0hJ3v
egCzXx8dpi/ygzocdkRxhSuakWMvIUideHrtEtahSWH/DDfcuw93akxh6lffWLSk
VmzBkA+Lz4LrTAzv9b/3LenAc3NkgG40oY+D55PwCAY0LN9KU8QK5oRKKbZNNwU6
ibMpKHwXJIplmStnAk3bTP0aAKq0azN7MjaRbStxxw0ENHLb40KRS7UdS8o7ce0l
k2F0CNdCc5RMwwJyWKGOYz80Kg7R6lcsx+mdUd0IxzyRFsiLIDtpBWodAhKrFGTN
gy/HkewPDJxI83ezCAkivQQ2JqD7Dul2rLC4BTQTTvrcqZkHovv4Ixt1/xeIAuvr
K2+tQYzVTme/W/Lx6u1DUCkGcwLBTvGkHvKV1RVMsnW011rkgJvMlzdNjNv3zphB
ae+oSE0DSyNrAHbBX9ncN/hhE1IwMotd/QEP9D1sS1WtZPnWTAwUg9iuSB5qsE3F
r5ESJyk4OeqMlrpOKMQeY0AeC2kTt2yvpMvevtwAAH3L/qM9NbUwhSvxsOKfIAUs
H4Ffdjb1fuZw6hTaKe7XLOasgB58fDe/3cU5LF4lFMyCMqnBh1JpFr9POCufeA2G
CvqEBMvNEETadw/LjzZfma4c9iy1yeW2VFEnD0MhYGoCA6c8mj1R737qhUhHitbt
2oLBpgAEWOqj2apz9HjUHXi/eT7HE4oZq7oEV8x/f+b9wEQX97SaDWD+GEABsypR
cEqR94ytTodunoUJWRfqRvuSqRNSYVoVlrDLZWoH7OxWAVQTFGbQNbRjnmjTDpjk
tf35POIStF/C1T6voFNV6RKY8C0XPQbY5YuOEB+lbBiwq5JlvGFaWWzQ3o2qaPp8
+31GZF5JMcS9RnOit5s4KWBqXrNQoI9kTs+F7N6+LKB1u4GeZY2lBN4W969hC+yw
M36e1bXWenSQ7O/wHmWq6nLi/WD2Wvb2wP4R1POfJqXR2oYtTSOI7rSN7BEtWCC8
yuZXSn3YAXUY+Nv9IdDhV90Z1Q8o0RYK7fbAU9F7mhhT8poWDP+BL1DmQ+zAjK3d
Y5BHeXbwbvLdHkvAU+19PSo/YQ0jR+w6BsySZkteV2LQHfbqxugfH8Bge85jzUXm
2yaNoJeFxNpe54dR/tWOhlCwaQN2IAWQrtebIIKRnAdb/c7U2dvVAo2BwvRtSHHx
qISlX/BZky0lAO/Z4z+pf9bqjAqQwR8ttglUIr4HwxU5h6ADA03SvWTOWfxQPych
YkWbqNGN81p1OuvR1cnxE5AoEm/6COeiro9lxuHiXWRdxW48vCRMdwIx7sRiUnze
bxG/apulGAEfn6TvbOGxNZ8M0obLh3ARXOlXByAh3EV57KAmYbYB64NV42pIJ7Jv
0fq0+I+93pp1SBXNgd+cR9TT7I3Ctb3kek6rtGU69AE3M7Xgpv5OX8qOZkVOKXgN
Ea5oputznD1mugvM1L9XpZxN5uocQwz+CKGlvzY+H/NG+hZJQxr1E4uZjYrW18GB
hU5W8nO7G/F7q0wRHnb6XCKvJ8eGcr4MItF13otexW0nttDbUonApIXw9Ip0gb3i
bgAKUBD55lC6ZdOwDd1ZBe1PFChsUa98iWEi5H5zAJ7JbkT3tnJ14wJ+5wPmyCCv
dUSuhxLFXcA4XsStorscKkQRjOoYFKVUgGHxDIzZ2HDkdP94P0n4ad9Fg1QAexru
pvOmovhq+pJpnBhKoCutkX8u+XKvOLTWq85NXs3uisNUFBC4/PHmFwwnEu2WR+L2
t+qgWt9bbm057mMUoMWP6TkZdrr/+FzDcp7imRPb8awUMkC7lK8CRIwP9khC7vSw
mkImc9EOtYF2mrhg5dQBPTmzkbOsPQtbiSOSCytJ1S8KmbJe0HQ/BHApahb1uM9U
zLASikcXkJ9T5sRRbve2FVOX/alWdp6P3s2X+07Je4mgiNHoUNFuaySS+r2Zc+KM
ZiZ+kTSsdlEIhu5naOmG/QlsVkrOh2Z6eFb+3/DeLhBMNgyp8muP4t/h4hgeeVa6
5P6Eduu4IrCA91KxrHGIgSF5J9cd+Nouqxsh0Ct8a7+FUftnIlElDd5qVNSoJxKY
TlM5jOxwa+/vjjaErc91EVfqcfZSmHLZus5szQY9VV3D3Yj6/Ls2vtqPvpxMPJTH
NR+XDghdBEHpYFq909u904yKEABS5T7rrtEB2ScjmMwNXPD4aBXW4k9NDCYQfkZ6
ZZJKzs6H6QMEHkAwhvgCLGoPQZPebOiXz1tuAO1BK0yYPf3TjwwlqvYZy9oGvJPX
4U+BKEo6xDkEfPRvaEWkpyIq/rU20kZYDmVE/Ic7Ojj3AHu7inNqC3ymY792tLjg
7QazfzRRlwARBCZ7RTGyuAXX47kS9wRxuZImzVTP+dC/0B7GsFE8sAhB7c3akgwx
8KFnwA+qSSGZZS7SbDgaZ12VK3BbnV3Cy2J273D1/Jk9K0cHLkXDQeMVlzi3J0ID
WzwOfU/JBURtb4fOrne00633fnozHk0gUWrbUvf4Rwb2mb0yaYAKpr0nATbyrvef
szjgfcY7KWY++KHx1QOaEerl7RlPDeohVE2WnDXKPCwzEoiEsu3RuRBeU1WeIqiV
qloGddu8EyE9BShueYLqNZtOfoWpvjMHQLrIsB1NuyEpD1BmpEUhEj3hpUyxCNPr
okC32H2os4Xm9P0RFyFbT+peHcXQen1in/gps50K0gPU4jAtr3fFaBSHqgGSSydO
rpBRs9gf+59JT1H7ezVNx57YmBQASK0u0lnyUb2PsmH1BV1x9hBaKteHIZtnyXRm
o5ZfjL8XcXbrynVcIj7TZfMgp1GDjvyBY4KNQQ2urSROnQMj7SKF29nM7gjNlvKC
NPs3qvimrkz5EmCTYtVkEGAv3rDsu9RTlK2dPge2DoUYe+8UyqxsOXrcpwKSGqZR
3NkcnG+JsVHbCYuIR12bhi0Mg/FlqSsEHL0cDPVbzXNGAOdXhDWm7sOpgvTz+4QO
3WznbqiYcK1x8CJ+E+3mP8tpGoc5hzUhiZvr5BLK3dpuDhDNO5OvWgqevsRyY5z3
DAVb1man3TszE/BKcgIEsx9eyWJBHqTWrFDloXZTgXb5eHUtnkG97YV3nTplTQuc
YHZj+LYoDWFSTmrdMXMl4kkruwlo0yb8KO/xcLbVrVRa/KpOkrItyl0SkIACEW3x
5Wt3sHyAtlJOsAlaK0wbJAXeAM0vupd1K4uvB4aSHjph8ZKZNHiKZKZ9AVNP5IdP
XmuzuAdC8XykKywein2xzqIGf1IddlCik2hBWad8LVpqDq3sb0Bjl0wVYHH/khpB
epCEgsazATXNSIkTKcbYXSVZZMpV++S7E1xnu1vHHbMi+Po+f8c/yBFWHdaAPs2K
vej8OsR9mJR8Pv7K07RLd1iCfQ18cEtN5VNPLprWf7lkbs9BUlUBUqboKWcCVsa4
yW3FAjzhOla9X1i1H1bR0xkRpfBji6hyFNsIIMg4LiHK8TqnaZvhyA7rntSuTc5V
ODgwNOrUvrhHX+xA3hZ5m1PmfkTJ51FC/YXqn6uBjb0UV1JQxkiWbzxGLvXuJGwh
ZfpsEiukmTHA/Krj9lo88vyJjYZkfvEZH6t7W/06GeG8hUYf7f1CS+lNJKT8zPic
CdVmLJIB6jRnPER9y32anGZvOXGuki0E79UtQ2RcNyHNhbRCBlfcC9IzzZ9Hbb0K
8PDB0ObJhQThmaks66d82S8J/I9grk5Pq32Rl7tzq8HeOc6I3N23NI/Kog/Aqmrn
KaKsnPfGGyEsVY9PIDW7FgN1NvwQEYyefF52NyAKjXlR0l9lXPaG19igHfzHriSZ
ZTLMgR6eByfDJzaM8eFXxcS426lcpeeEVscs4938H2eWzyYU0hSSzhMiUlCPTOpQ
eAuuBO4LAk4dWyAbEJHe5a6ez02xe5YESxAluqv4z5jXItWujeb0tKQPi7jT8pxY
eneGvhen3K5uCdQXD4Qv3t8d9MIUpT+6aujxmP+0VQuBdj/dlgOoQGNooacwBgfc
zdzTQMvHBvgXUQ022RqbppiQTg74Ksd1LMxqXo9FuHjZVYU380IUnNdNpX+Jj63c
2m0LB/3nJqpO8OvlW8zexu2x3/WCODHJ+HE4Py8WpLqKBruro3JXMjnKaGiey6Fz
LYTAxDkXCiegcEbkNIU+5soVWPE9B8otc4Se90CkGM2xtlVEoqirtSPwBuh9vu6A
hSCNGipW0+5AofR53mM5TsIGkdKGvbz7NePoL/n/nRTJhJ+2Ssk8mJFiqheHSJPr
UwWNUQFmW8S0erBVvmEyKKR5orING12rkRw+ZnAwYQIU2PnTIAuohENM3n0DtxB9
gPvWT65owi1R915cNjdz4bPJAB0S+wl3W4l3WC1Z+FREoim/tinE+irykdN77bZ2
bci/t3ls3wxwNEAXSzahlgQieT+ea4sPfj7fF2be1h1Bm4pgOgsAbTLMopPphsMV
HEmZUPmpjpZGAI7R9SmPOwkCK8uAbG9eYTlM23ZA39xpqq0fxvpsaoxJxNolhRsE
JNIQKIxXyotVdhi/N7qcqV0z2EWUJdM0lZUKkS2LHZBlZ6k/+rIQd3iB2LFwj5Ev
FidVESckQ3q6lu9bgGpL0mbMOGh9W3+S9Kk2IqDNlNIcf/HWDfBHb1X7V9qVjDF/
WSms1ES/NPs0q0mLCw23MdpxpG7MdYmrLY6labYxJwcypX/yNE6C9tU8KNBvxEAs
xhHSDiZQwdPl2sg4jp5spK5YLun3s9SBRgVGDq+yd+aI6xmIxGnl2F5Pt9H155F3
pTSL1/JpAp9M2QB9KBlr8N29an52HlyIVpqsNuPdPM2EwbrI0n5LzI225ALQkZWp
iGSOkBySe7qDnIDNMQN2+NIG3xL+eIQnlUBEPRvLW0x9b5fblMcYd/XkT+jwvsAU
MRo1yOwdFRlV7QI7r5zTBV6aW4n0gnZU7+N9KMuDTlZRdl8eRLfsVZPIqnYbwZLb
e9mFXb8Q/xtSMybB6DVW0N2Dmm8NrxNWq5gPkczzwuhGclvazdSpJ3l+E0ttjtvJ
qMgN/OmtHYP3aTNN3L1ATH19DdUi6eaDQJxuTu5P4phbtalkgGQ0PtNCnnZW4nlM
VoiGy0MLT3vGFtAURTgpwCXdvMTC4LMJu+M9MFwPPpdYl91oCED9rM/jq+JYgO0J
0C9qvbjUkmd7b8TpI+obmVX9Ml94U8gJ6oC2SCcRdKbt8XBhYmbjX3JPtqAyb5X+
9KKIBWAPPRoROw70flzITZd5HVKOxc2/OW4o5iqHXVTBa5BFa5kPJwdQF4OO7HYc
cZb5sqi1HPsq7wD5n361XVq1Oblm3iaE+jEF4gUfNw2yClo4g0BWkcUzJjYtpsQV
32XKHJfshmP6yNaHCmF5rsRP5YKLbNUpZCHYQkMXfJ3CUuYuO+kqfzdXsy6VTH8V
eQUbZaX1d7lvy9mJnqUkaWzEEcVjycpNJF72gZt8kPj/37FpFzP/gz1PvJAEiyyF
LgFXcjiDfi8JF5OGBN4WxU1FPq0iHGr8HpU5y0KzLz9zHk8IS8mKJNjCG0AqoYz+
8L3LeRCpZTvdW3qDYfGelPhcX0pQOqBoTcfd5Nxqg4gl4YdlP9PwsWHGv7ex0dkz
20/g1yycLLehKAjY0+Ce9lbA/MvVZLE8UIsPTI2GAfZUQfY0iFan94di12qsoyiB
v8wJ4QUm3Biyz2AYZ1eDSDZW0XP/V4Uft69RoyVwPCRo56mRrEfgUcbrNd+KpcuL
r8wHIDXPgEaBgc1cmoXBFVw7xwjl/YNbMqtdmGLywIWdt2I+8WVSeLN2nh0ym5Jw
VdOtPakq47vQjYrqHsKWR54oV/hG+34zA8L/hnoZ5Fb6rAzXGXF6GV7OPM9gJRA3
CxFk9tI4vNKa3PcU1CduuMwB28SCle4h/3l2d34VXBnj/5z2CjkFNdFg72yCBvbb
Sa5sF+aEl8q/xP1qlxYNLRivHNHUy/wgADKUZrA1j1W7NSsp8Fpd+bmHOPfi2Fd3
vuNaIulDcM/yKw5NvBKhbLN7+ZowRawHL8fKlR2jiuspjM+/uYjWz1bgUKpfxE1e
MicZQt47tZbMEz1TecL78/woQobtWG5hwtSTOKOXkF2BcWdgagtYR3teqZUycEn7
coITvB9oarZD12wMbh+Mi1wfSOeO0rTraOjo9ZzuP9VEUa2JtC32e8GCLmyIrLkZ
xCRlKsUO4M5vfIT7y96g2acajDOqvhEiPRk5Q+NkDdGjg/6gFFBRMXGi17gIEQCA
2I4hy8AqNWye9KihquyhCK+Sngy7A3Wcorx+CiDrrSAphlKgcGAHKtfJPu3HiXug
RvXJLBp+IRUrFClVTDlnvuAHrRo+fs6dxWW0SyiIyXj3HwOJGTy/L8Ksgq5wpEwF
anPjmVtjhHgaGEl7Eq5ai3R4YSML230728xxyW75nxrJ+bi1WoYziUcKRIXmbyBL
W/Z4AK8X+rsM5EtBl2TnVZzIZua0/D54V6ctF3ndc5QekfzeoIG6PW+ys0RlEzkR
8Ty4IRcY7MF5ddCa7Q5FAQJa+PW2uUODP4yn/a09C2QaTnDFQs/2bX7RMTn8lIjE
Osny8eq3dntVeeg9PgUkAq2CcP1UMgC87ROEj2j4SDl4TIrOPfNdxmMdozO1PWq+
Wpq619fq9fxaiolT8XNl/15IEJmKPpn04aGGl2Cqd3s+G2b05EMsB0T2MJf6oN0r
Q6nz7OVGk7emM32zhpSLJfYpSj04NrR4Ts7qicz5/4rgqushHhsM/nDcBjhhRYCX
HUNLKl6g1LzHa2JXBVCOmSU0ccFbyEDTFCDuWyLdqMVeGZyVrMGQrqdv0EEoc1e/
iNL5tPnd7FwACzXAMQxmE2GkYYMIMcyJ3w9y0zh+q1WVxBhMc1GJsKvGNPQcByJf
7eeWISz9x/M8RrJtTUcCx1q+/Ega4Jjwe1J+Wx3lDfD1Hm4r6PJ62wRiEGoIvNhY
pWfC5y/TP039/rWdWcO4qxOh9zmsA/BfC55IoCq2Jdg0mPtCe0jNudKHaDCBJKKf
YqElPlb/4UbPXBt3K353IFigE0OfY+TaPcTfs7OP7zSZXKERM3eU0if+TwwvPBz8
oom3+RvljKRn3XQV/cYEDsI/kMNMnagor1/zgIepTfolXwCwi7+K9Wfq19zthFQk
AJm7ZWdur6UIucIRggogLjs5InsdgkERomi1vVoMjMUOuL8T1QNInlmtK2JNrTFR
Yfrw/RdqkVkDnp8ldxawwgm/u8u3JZGU/REkvVlsLsbel2n2TAb5TlktTyjFB9Du
fKKLPidEil9n+NWMyKlcgM3hytwPre2bBFrhSxQcLQSAqrWB5RCPPY3khYsX12ga
LcOGEBG8Zzy7bgSw8RsafAQfJDIs/w+HRr5nDnnAdTalFS6ALpD2KarA6xpTwbfh
QXMZM4JBBB4ztvn9Lx+C9I0xgRD7oFGLLNOLY+6p2BwINM9Xqqsf++BtxqR6dnEj
d9MNIsT59n8HXBehCOC6D+wSQV31xLLSxZY6w12RAbhT/nRy9PBzT1sEfYZAIyqa
aTTrPqxadu24YIB34Wl20wwMeT6P1gBC34rbXE4LBmohpUd0L6RHZ/SkTDtLeI7f
fmVb6nDqb1ZqMdXrOtdhxAbcONVPUnYygVe5qXxwpA1xlGqvo4DXUv26SVww0n0+
T7kOq1nlIzDCxm0VmfqBn3RK/t+HsZNtBVAN3uBk0IKC57E5y0LPGDVCmzveZFPB
gTkgSUE+PP0Z2pJHRya2vOckyv6lvZc1J68M34CYqCpLypjqvNCHYp5vcdCKvkkM
ZGT1YCITr/XznP68K5NozuGJKdt4OFMKe2ZE34HilhelxNYXQbmuSF7OxBx9zvaN
PplqVNPpgqmRv2LcrCv9DW3++xOk3Ai/TSAqTNQcabK2R0dn/hqUl8IJVU6AkpW9
Tmey6g9U98ev4FUfNNZajIafaHHqa2uwnX2p4qtYFkQJOZ+7o6UDS2UI7CIQiKRI
C2Kxe0qVQFy3AIf4/dKCAeL95b1Od+DDm5CZIdDfs08JPcgMJS+Qn5UnKO7ISdxp
mQ2sAcxETJXq8iuijOh0OmzEIe2y7jrfB8JYqD2xbNGyJ+8AKQ7tAHrXzA8jSQO8
Hg2za+A813Bor8gP0QwuNCrwk237pnpu7fYec+Y+l6l2nlpJj+YWbOZs+t0MrEsg
j+zWT5oDx622sEQpIaWuGVsceAr7ADFxdh96l1iFIajo6Zo4xyAlb5+xP2L6jWK/
LFznsxGTfIFn97QtlBkAcPlyIQ8Zbzo0FpRzud88+kr3gdwMIrJc43tai7AMtSdJ
4BgDwPZ8Clg7HJVB+Am+TLW/MuXOTuO8YmyUozkshkFj232nCDTpAvsLsed5xJfg
OBmqpO0/RHs5r24I4PV+Ipe3V9rBf5hf8em5DrnlLghmtGt3uRugeeyfYcCF9SoX
AewuqIk5cwl07biqCTPHiBTtlx+mO2kiPMnJuc/SlLqtU5iH+OF+OP8I53r6yhb2
XRNfRvyYkXVxMg4J3SQfsiv/uoKZ/BfkARxmqDie8S9qVWsLU28A0lx/cLd6J3Fy
45u2zbwXchttFVofgOj/HbCqjcsEw6qQhiNOrtEwhEIjGhUla0UrWP4xddB2p5wr
8EVK0TpdE1U2QuZdneBhvRaa1HzoPzOERnAfRk6/A0RdVwCId4r66FTy9s5XSrtO
k1owRdQHXG8wZN3NfHoJxuDQ1YFY6/3pCaabh5E3bp1WJwikFrKxQhczTrTHcrjR
hthCpMcFALSzImAGt0DwQUyLyGalnYcahVuTDy106fQfSBeah2zN/Nowzm1jfXwB
YaviUsMoK/fAP5mQ98FgW43vmPZYpsxNCviZwSKxphg2ZdCH/OiC1DMDJK+Jo0YY
/+mca9tuwDXOZHqwSAzjghZ9sZKczoHrlPXkmw/6E4y8VSdi1VzJ0bRFrvqXS3ZX
Qs8czqlV465wP6P9ss8wvDMLHfQewNfwze333K6iJgZzLdAdrdQP/pgEteBhdR9g
ZlfBTNrjYNRnxa5Oj4+8WSeVZldQzQXc44IKbFBkDu37+dCoz2v+CPBuLNencmkr
/fIvq1GLzadqfLpVNz1xWvjyJPtYBJK569pGsJavRH7xC7t2+FLL+J2y1INySz1f
MKR29qD2QydZ0eJ7xW/TSJPHck2TGNjvhyQOKtaaFgLKVKU5QYqyqviLWerpwaKg
35UrOBnxomgBwmFuDsbW7WHIZKh9CZE9gudl2v0DOeRPEx4cogSA4pukMRgu8G1x
xD6mIsJlhKa6uvxNrMwkr6WCRED8drz/LV9ckW+IJZ2acbuEg2jZxdG4qUOaoJGM
iUaKBSv3lFyq7zsqvJl6ALzLVF7S7jenHb3paOtFoLbGQubLld42rm3UceyKx56G
oovrihmR5l8fxGTSOwm5KMH7sD+EPrN+z51SiYoTzhN6brpUGcI91NuNvQQAUZW4
ab5wvk0u+TpY8RCZgSGxUHgEK9bf//3pjGU8TAmqnnp9x4+gHxmZlzKPeWq/XnnL
Kq9/cCCyg0Myu9c9GCQUGZEJ73D4Pr4jWtf96BieuaPwU5Q+LjZ5LZe/sh2+sERK
/IRXB5iO3ovfLfSH7we8W1Ci64eC2FTbKC3RAJc1fOqeanLwSlbnNG/PhQuslPEz
pdxrTnjQvRMEDaPHTnW76jUCry3409wmRXis+pvvzS3nVl7ByXLvJd/tpzMwJXgn
OzAevbFltBcpBD9IBaUmWn9C0OOUhvgsfVSXjJuptZ7aEvU6wEoBueWxPR+rtKDK
W4870HppwE+pEqmW6RBorfwxwRMBLttZv+b8fnzPkZvEV1++JdVGCC0mMOpq3rNm
kMPpL+cjN0s0yQHDP3Pa8ZPjC37grJ7CuJ87B5dQvbyHQ0vHNgbDqnlb6ExqQtvl
1zRMxY0fHm/Kde1W0J8ejFV2xezGJdnodfSPHahZP4T0icVJJvmvKsOuEHChLcGu
0Wnnm7BNpuwC0d12Eiz45xLeWnIibseYsuNjhloP8MlWlUhVZkuia8js36K7jPsu
ij/P/h6VwVHYgTyjczaR0RPp/vSbwiZYi9ryXzl3iBl3BEpuBef0aYfhdoPOwuD/
ogklZ7BWoOBeR8Df3bElOk6XOOvv3JDNwzAGZ1hF23hQVL23zvqDbn8opHNoQxkV
YNdUlQA7lwNClM+Bv9W3eqv50dUHrAITAQ07rRLin4EeZ+hPxKweNXILaqJFXcP7
s6oNZeVBuSTFRIGx91Rmty2q9pVD4SYrIhQrDYQKB0S8p4OG4T+Ac8+Sj37DEE9P
dsY3p9VlB0CTZgb/5Nr3Os58XfWTRIIF73P679lI4RCCnz8kYjtooIzarufNi9c9
mYNg1DI7xSEmNegqiTA+8nJH+nZsaZC2zvclrBHxXbNs0cVmr5XVNtHQyUMO9PhJ
lm+y4lNFOQtfVOe/hjr5cLpbMjdNXn+kDWm2ta9y5EqY1hCsTHMpKeuGXTc3BNTF
LQhqDaYlrk7RRAoTJGt9rXjKISU8NFWfwhCK9biTGR9uvd37VaoEMKweGczflX84
IP3wvt1tw43mHiAxaxtCTBqce0VJ2tshZmLbTSaEy6wYypQb8HKk96/cikJ3w87v
NjHLsH5lEthnixIWC2gvw4wt8KWhEHMkcQrB7juSGEFj4A7ysANoDuPGPxp/vb/3
JX2Tz7usvu8v1xry6IAMU6Si5DzRa/xDuDOfbD4ltppPGTWH9kvJZrzc/6CBg1nQ
tzFARem5aho6GLSxJXosu8Tb8zr1gGDsP8sSPNuVnWhYVAd5E93W8Ymak+kXwyGJ
u2KKsyVmjsVMzMpMrqzqx2Q4hNTRw3wp8B1afFXMsLjiPBt4s2sNgWUI6GFCYAYV
TSFXNabTx89zCQiTtt9acuGDK9s9ZvXqsyNs2MJ/Vy/Y4ODyRzCpq2huzQWLeym3
pqLYhNGrjU9JdsNJPXZlUmX4QnnTCddhX4NBml1GTuuE7vP4pvitgjKLlopO+yhU
N7xwjRRt+Q+qmBf1lnQ4YxZYrqAzGzwLSQnzPjyyl2gqy67cT6bp9wzxyXyZBfvz
H5GW6iIQwQoiI9rfUa3C5cC5861EJ5N+iX0IJJeFtv78ZLHu3isaIvasdCvbPhV/
wdmNF1nxl7eVmGZ1+g/jhM3Z4f8y5X8bhhs9w9TGvnk31YrJ68E59usIzbT/Tl3Y
MHGMU6WfEHRWLo8a3wzMLPklx61P334q4C8JeBgwtuCJN50NqnPzZ3JWuWBq/CIA
VxfRHaAjtiluhm7yetWiOsfG1V86kpwD+/A2NO9kWAf2O1jQM+C7zdoWnZBPvJOS
2KOGtaLu0qHxsQUazXFxqnwNpVweKk4h4m6QIIb53wQKqlSMWfJ02+cDbnEJ2h2p
AHV5+IV2guJmY4QrnuBvlGLlG+1nlt2w6HWufdZL88xumg3Pkab/WUcOqkEnkBI5
+O4Q99dNbUpwoqJ6lf/WYlyxyWV3Bnknii7CT+EfplRQCaipqfTJUSzsdTq0qeYt
1fCFWEvgh61Yh/0dvuKQtI4b4ieNIwlamt7OgtF23XJ7QGFFxbrD3gHCFT45493c
7ix/J7vmWKwH9fpjySuLwa8vO99Su1/HEPld8V470zJGLEGiBnSBwtEymsBvZLuC
LR9Eo7MraWKu9fW6i/Ad3cvjw6p/7/PC1jJlMO0TyQhH/8tzu/QOvOcYHM4koQFM
0ieuMDyyBlw0htCNaZNp5DjYbo0vqknY8jktLYhC/+58g0sgL6++ZQ6NXQ0dQvlE
9q2id11uLwVbBI3DOzc9hy6jJOatj5zG2MSAGemZwX+GwqMyPMc9TyFjfmptrIIx
MnMWGvx7cJ5IkeYCSOtj8EHXEt+Er2R4wWSOkG9rIwfrVJPw9j3GU2JNXX+UqbKj
g7k1BDW9cEds8jTiNF7YU1PbDIP6ulmzxHrkyFeMa28ZcC/ChVUB5D8cxj+qw+0r
R4ictWT6P/8QrCC1+7bI6Rj5cTmbpyOntn2U5S9LkM6BWhvjsEP5KcGhs20gO4S+
lGMs//eNjLwMYxLUzG5aC7Wrk0eF81TszIhy6eIn6Wy76rQE2h2zqDxOWLYi5NWG
+sgjFHU1FWPWEGs93euk9dxNBb5QL/qZI95B17Q9T3Qq4dx8uYPh+vEQ3lBdzD+T
1BY6XQB/3w+sBXM3eoaaMnjjI1TfGCN8IudyvRxBvKtjRSXELu0zc15XLmc64sLc
jNDkMvezbYqMFG32K3iIhAmZI5jH+s6SX3FGaWZM1hFEQl7/kOviV/nZTayNF7gZ
wBnJJid1nAzxHibHAICLHnsYOwsrB5nPnWbeHkRKLyKQEZTAnss76NCm+/vkYyR/
Wnut3uCkJi3aCQxpYzTWdQrXnFBnkoBMy/C4pwrPPah1Nwiohf3vPU6yoqhc0QM2
7h0e6fPk3difaSNzGJHnJsrjatZzXoR03njhDl/uyCt+1yv0DhJvKjCCxE1Qv/b5
ZDx16G5ORiQuE/3heNuFPGAh9XFB/j7+O1t9/blS6QjH3JgtWZ7oAitUB4HsKeBA
XxRuDtlkraooHlW6h07wtjMXuzSWAvxokboG8xPI0IWj6FYvCI1WcTKTscbkenyL
13IKZU0KJh9mA3fd+aA+kFrfQGgM4SP2NJ3PgFe0fzeW7Qmm/fXBcwz74VfvdcTC
bvC8Cr2bBsvMHaWLwUR1tK5FON/Uy9k94CNTVESXWQRjb83h83iwjj9mGYCuMLCZ
s+klUtDXi9w3qwRzdTlgIP077kIxLwp9g2E5HwAOHOVhX9zzu8O7+9T375G6AWz0
PKYmhbPvl92qdqXNRSxXFBNiJwOGrkaQY+JQPVGSNucKDfpoInz5BP3rionKZo3T
xCIv5Zwj+JGxxLMjxr1RwttHy7Rm81Z2bAfmmJWm43+aNpvkqe4BVnWs6BF/CHcz
rP2BoC/Tk2KujNLkw/jtJRefApYRxg7qH1CC5k1HCZwH/8WJBU2ey+oObnGGDTod
ba8pHO9iIyh5IVpeH48E+xWx/Ns+D8A4O7xusJnToTampja3UtsW2WWFpBFb5y0t
pVhqTn6la2DCTwDVJsvzjAs++sLSk+zB3WVGnr5ECAtGDb1Ln2t57b4hCn+cKf8J
+NBLdAdM2Ki14XZYLNw47MFKDIgZ1upNYsvfN+GzWui4tjLjtDOxgJR5AGuO+ViR
L39WeoRK9r3c87o8r5ultkAGJaq+b9m89CtrnL3F9H0HGPCHC6AtVqDXCPi0gl3N
6lxNs6PlxTU5sPD0KFKCnoAA+am+BYBIre1RQdv+1GP+ALXSEzQV17FZ3eL3xtZN
Ly9Il+aqE33iuVcji95OOTKS4+lpUKVyKdY+PpWt4m9Mk2RL1jUy39EL4j5Eocf/
OTdcwTyO3XgioKD0jND/T34n2lVDoQodwa6N85/Qfjnc0phEBDYPOphJ5i4cR3Pd
9VlxsM9wvpUQ0Rnw//QkvJ20ZGLa8G9s6I/9r6MziKFmTZa0laT5DT/SX1bjB6cD
/3kG/X2OQFvrWklXBH4vvUmz8eEvVR5/05UpqXQa1EnJvhXtu4sGQI2DhoEedUw8
gly1TfF9sEsiPb6ZEOFIVNFFjKOJGFaLrKEvxmLCGSNjMXAdUQiImWIfkS8MebLJ
bIbe52qRs+vZ44235lUar9scwrGEX8QAQ/jyxT73IPFSaaUmSVXj+EhaGCUhTLDo
vW3msqu94ExshJUl9ttu+xAprTN+ojP0pw5Cj6xxJP96W1cyU28NMNMFVK6l02fl
V0WxYn7lXvOh39/LLSefTM00rEavfnT45bFlJXipmDWDkJQxcfTeJFvzOpjOGHD3
jCVx2u0Z8TjWnIOMGu4XOFY2sAVBBG4ch2xdmT8v2Dr9n3z6biYzGe5us1kbsmzL
RdizKlREjePM/ll/Hlb/0oTDi7HbjIMLweeIdHMKnLuYIqpvYhFhwELQJYmV38Zb
222j/XtvZ99sa5AyG+khPEKXZ15yR9lJ6Kf5xgUorkC+ySBqcczRD0P2qUwwG3ej
6C2qFpYDPRYq31lxvE7RQ+g6Dw6oTdv1oKzaqudkqIMQ/+cCpdh4aFK8bXjQY8Db
Q73TjQ4oJ2Pw69FdFnxhKsMLU5LgylhjSGrFDCh5rjZy2J8USj7FhxqnfJunNQzh
5mQOXdfR81hJp4TWFWSbGm8fXxQj8tYCXeqBJ2b8Ky2iV7lVXpx6mINpS5zMBEwU
Xb/4P6owN2CaDUi1b7G9eZbH3/Uy4GxXFKR0L1VGAVk3fs6JBqdBHJS0MCOGhQas
U+TT77ULuqsyQG7ST3cviPT5qyD5K9Ks2N3iegMxmpGT5TFi3jOp7SIbGvb0Izu7
dnl4CujKjEih0vzuFQ6VCPVU/JqxT8Z39GpYc61Q88GKbm4wOKLriXYJ3oYt5uXA
dbochtzIv01Qbj5REcWq8szLTeJQwKV0pOmkMVuaKcE71h7/wrViI6u1dBvJQOXA
6lMDa7KYUCX6Q1ft3ro/D7g58ZlHRfkeZU9rQn9ZCgADHGkGtv8NMmbQm/li03x9
UM8rft5K9jT+0aVn3jSKc6vQALvWB4rQMGmP7TQ7uPc4ie/1KZk5cYqsQCX2Q2kQ
ELTQA5Is5l2dnrrASGPjx4iGvWV7Z14Sefi7ZpSseDoDX4Kjn6O8E20QyvGhv+IE
aMq5XbfG8GAKG9fKEdmQLbbrSO44mABR9Bl3h1sqR4A0ug7yJ5fkXLXyNkCfVHVT
qs7sLISg/IGSa50hHKExXL1qDN6g1Ve/n8mkxjqmy6zaDQQbcq/0DZa8Rx3PA35T
+4zMMpI4JkVd1Ff0jhDQLnys4OzqjShbLFxwFW/ehfvynI+51dqDZEmRSzAImrbm
6SdnrJrXSG0AW+QcC9zRpV9meYR8r6hjOZlbPYQJ1UtbzCc9/7dqkebZqhQxBmx4
T5d6aa/WdC0Vkoa/QuKm3Z7H1uShCuqLM/B46t50clw6tgG0OOwsdd7zorGnw8DN
UJ2JSlrnBxbbE1I4erfDHJEZ7nIzIx1qi60tGJnXKKK8Rq0vMhaatzgp8s1F/5WY
vlRodHQ9TcdgJbMs2Xt8F7TCiZzrHNWwb6WgsOaOJFoOOvw7/QDRWuWKz6ZmRExi
1VhgBcVz10+sR6CWk3ZLUl0NtY6zkH4XcdpQL96YQ/nPxX8irDKALG1dlCd76Swz
lPEJ3PLCesXwyLx3SQxAZCjWhqdT6RmVepBKaqhiiAVAAsXAPGC98qNq2/j12t8C
nHJOhin+mZpH1wyfWKEOF7WVurg2wrukdS9clwbSbKtj7t0fmbS94XYK71I7dqme
5hPTWBRSd5zbw7Rap/nycB/LrMrDMyipWiPdJD+qn5+wyB6hHweuW31zjGc0/Ion
5/nUhICZ+/hA2CwhjgXSYqK2VP3u7nM9mzm+BJr0/PvPdsciszw1QqHEz+afmYOT
l17aNocNNRjG74ibDEleJdEUjitzeIhwWGFm0CJ2MrGbkT/BcK5LHDDzfl3ZjQYc
anPNm6Kk8R6Olj/L1hxz36j+RyNL0CZiqeniMQ/hNCoDmxwvXDUdkRE+xJVo2gMM
hx2e4MxylwiAZ2jmdYGCxmGFHI6qkAxHJcl697JNrWbTNIcLcA314Dp9nf8dJ7ZU
6lnvkx+NXelZz7z5yjwskj3ThThMSrABvOApB7DgNUgxtRIUxw+et3IFO6QKW3z2
yWA8tsVU/PX38z0LexpExSeXyAOhTDd9U/8zlf2ZMea5ueVrpLyo6On5L/j7PBqY
MTw7K0lx9fYkIn2KfrWO4pFvy9b2O5sxXmbqruSUYeR3S4uI5EW6RD5G6tX3mlD7
MiH69smZrQ7UawuwP9nnA0mELbtXaqfzgHt3a52Ws47q0kzLXiFDD9z3RABSlc++
6VMvXri6MFECGlLfMlP/ipWc7EhBEHopIu9Fwv3gKwfNI/DICdAHLRdne7FhaJbp
BrF3BYRyIWGrljh7rk8xDPpC+RKPHtHEhHx17A41Witn/Ko1LUIOLeP3aSnwpF4a
9uzsFOGNcBCmZnwenXvXat3aVFAhoQj/63XzkcT/Y58Fkp5SF1emZPhrC7M6gy+H
+mvJjhWBCmZv7H0+k7BzeAE4Uh+HDaasfdCxLpW/zB99pEEOkhKkGpxAmVosVdH0
iabFmsdp9YwUE8kAMWnCrYvUv6nDSjFddDA4WxjnDdQEmS35wIQ0lppuF0jQIHgh
Uue0an4pLBraMGkNZnCRW3dwfXzwObpzKwlqZqtQQspUS+67fW/T3ydBxFa6Mupn
porvuy9iR/8rwGGxyjx6/ha2kv+Yq/7Av61Cl1ghN3mhQ71SSEFAw8Y+u/DtfR/5
39BvqjMaBN4bxehZ08fw2Zr16UwFZSfIRB9DwuLZzrEh6XyT3RaZP/gsdflb0YHb
CakYT+SMWEgE6Nf22N+8Ye7F2kpIjOhT01b1dydBq8Zxmm/iAIQUVOmcBFACqNM/
XUcyHi8fHXbY6XGd7ylB1BRJeJhiztoPsPodfYdjw00RbirigVIrZ/Yx+ZlU4FYu
t3OfHi+AyGuFWnjMJy5qJMapL0jHivgufYQpwnLu3u4PNAZ5KbPh+s+PPZgUZPUK
smwFyVa7pSq4OjKMfQJNZ53EQ0jUiO+cT48swRVIw9B8x2MXkJ8R8kpn7ypmD8dW
+LFIUhfFnKLxuYCUMeDYzzn6vdzHS5Yt9kvBYDz7z4HTdg+l5ugzTTWhOZpniHHQ
ZL9L/Eh+XcI8srvqBwj53u16RXe1BSKl63dC6Y5AQK1/pcsLQWcEkuUqw+BJGgnm
F4SiPfkG11q5EhJ4q5mCSjIUvCyp0wSJvA/oU7T2Zj7r7QrfoYJ/dDVxtPqczWx6
gTSjqAguRRRHXe+PQi6LHiJn1ua0BvdZu7KV0QFEiiYCsIM1HFwWXjZuTJV3sZD1
eD/uwdqziKcXZqA2SJMGwHS2w+s+6CIi0fHMqcnTbK4wldydjImAHCENqBpxvk3r
0aLdE7UDLJsz3tCcMKhaMMP9iMMOmYUy79p0++1Rcx97GSxyHobe3OGsTZ4EYFb1
fUgPpfPzYCzqezb+BUC/3bZI4taBPEz/4omXi+Kg+6L/NITz/+z1eyBktcFxNmpa
FYNAEBGMHQ+MEtWp45z7c2gVSdGVy7iEkr2QCne4NHrBqJqhUduG3j13aI+oSxAc
PYlnD0Wx5cG06y3yS3TyqlKOnK5DrRq3v4nnfDfusRXy8PTEvMk9jR04BuG6wbS7
6SM/Bmz+wQu2dgAHxiisxONNkVeOrdxivo3+8dzkZBzAZXdnFvYbZ5bssm+R+NRa
YysMtz0okjB0NrKJvBNNBsuohpQn9xW5beLNnolVF9+d9GKR6GuG0pvdakQ1o7td
8FySikx4K03uuaSzhUz5UyjPg5i29ASn7PcbLKSXUykf/uW/arZExKNOqMa6ew9A
dQhLKztcsxhgZ4Pf7yBGLAOX3PYbKE+EneK1CY7Jc6PpQ8J59NHBxKTXEVFpH+wS
8QEkDkbriJNRzArRWNMAhh19xYcODPlOpyiOsyN2O5sLzMOxVl+B6xZnRhVkhYz4
1a+XI9UD1QN+uOMYydb/IfSjD1vH9lpw6NwFpaanDTz1w67BzZ+A84Q0Mm+y/RgJ
y8K0i2nhRp9oCwINloJbK3qX4OeiAfYLyYgXlbxTGMHds+MhYV1BCQOaLNG0zOTQ
HGtcVRTfoXZ8Dk1nvyY8esuAyrLAwzTEJ2AgSLWeYR1342dFdDZzSNjS6ODbUOUD
BBXko0MlTklTp7TqcoYTVSRnzm67YVfp3FSRWu8e4RKLsEkyRYXE7hIY/2T9W4EZ
t6b+Syx+NqZ4SovmA3gawA3clOZlFMXHo943mqS/XHsXg5G/uLiBGhIssUvDMu77
kc/t18Ccuj3fXVm6ZPxCOab3FS27rJEczJ3+Gdipdc8HOX9QZdDdfpljw4z4hMmx
Yf+gex7O2oTPjBvR0zje6EC3xX6SwCcRl+VhwSpVWjhTByz2QM8dbBPROfiQsG3q
LA1PfHki6QI2czPLdSR14cSKwD/ASDYzCPQjhWzlBoIRz2fKHNT4RpObSLjnafbU
3V4I1C081m/u0sUxQKgj5r6ttNByguXKMK7awLCu7x2E9OafFSASC2Vu0tPYQCle
XMEjXW7U5zVvBykN0LeFKZ2xzXJJ4QFSQI4dGQiZNnw6k7BhlEZV/68hvfeetWKU
CHGgoDxO2nmbWtxdCfHFhydGYYik+M+ac+6rnpyvP/ROzTrmxwlN850CG76xuXJ2
TmHoLoOQpz71EbbYHjbkiTHTBLhOZ6h9TyzYCngJV9IORe4+Y9//plu7xM4vSByD
4ckcFt/gYpft5RNEEv6nLMFKmik+ziBsgKLuedn07DT93fV/RH943Xc+gNgOHffS
cfUyaVguI2JQGIHQheb9Zv1phkwaV0h0pgctDdpt7JuN3fz/qJfhRIEX3z8FtUzu
qigIcQsjzTjVPuwHdfOEioGfIGBnpuiF70IwQxQeOcFGMML+4DoTdu9fSwUSzc9V
bg/IFsxfy4bqscZ8khWQLXkU2ZzJJPaRJE+DoawOYX9X/VQvtpzpOZQY3Q1ca63i
DMpHHGWJVqI9B0hO1672b8SbIE2SgeoNHqVqK4jWf+PG8QBnFucbjAmi3PCENqvd
jQ0wkxT89dJZtFxb4xbF9EYx60q8Tvv5TLMG9by7iPSrkPrAF9j7NZ6R1XLqLpCO
x6NWARnq182ZNAc4M0o1oqZqI4XFWVRd/BXUocwYSHqbgr44UMNBg3fCwB+OvY87
Wfoh28WERgvOMtkE9PLzXTtYhxyTQTh8B0C5FWmYnI8qsjkHNy4Gew3xAinP14k/
GpCnysRXLXDW2voxU04jwbQMMvI92YOQCe3yqk3xLyAKlEeti12kzVeHUnqMT17B
2wV2Jmv6qDmZFODcXuZcFbCJ4EXJlU5lT1S/TemnVOMV/l0ZQlX/adKk/zH0YSh6
HI40WEY/vAaj6RB2EMFpPzTEn83NuFBLa1HegQBcUDszUe3tXbE7gWAWV1l30Sa0
plyItS8Ktz4tf/uJe/iFCWT/4nKxywSsSlUHggc82wbMQvxnQU2irYGKOBKEnFuv
2OKwvqKxSIbOhJS+Z079CSRIw4YzqdivORqtt/mxpdZ5puzUug+m1TmeHg6AuccV
ueIhEup1ad25u0yKKELl1/lzzdBgcwAbhpglClF2t1jbg2MF7tLbI9lq7a4LNpOb
RwtnLgmT7WgXoRIYz/AmPZknYh2RoFALm7yKo7SbnGqqdgfeii0E8Le2RkWXijny
9rejBDAPvPAg2+6axXa/m9ReqM9SL9dPPm4Y4c20xQPaEc7a7hJUirS+VvbPnlrC
oFqMlc2WYurB6tJPgekec4GdCOMxwZgdiTB5/8n/bPRihQzRmBJfjg+AqGDHqbwu
IpjLwDkMvl7iM5DyhafztDbeB/Ckuhn8BBPygI0fVx2wI9ndhmxd2vAzd6njcQr/
VmZr9L4ESYCiovCjDHZtZRBLGSNqdHFGMOgOaz6HOD7szwUWnh7BEkAe5fOmj0zH
OVms2MCPcFo0LlrkuXn33xG7b374YyD2U5+6lEOuPEIuCrYLKxYsKCAu5IdXE2v4
j+AAa7kTNlNApQw2MK7ni6taQviD5ombBA5Ca3vh8Xnn5MbxLyRskur9xhfmMSrB
7stClacE75gvjgc0Ob5UXqAxQMFK6T5k1BCfhkAoCB9dDo3MtaXdFxqzzKCUnJDx
RZloTbPUPhiIXCrPnDLad8lIgy03GQEaTKERDNdYhXtvlWH5pcMcRqbMdu71sSol
Dst+6qGWp0A2tTbePaxN6pRL+vYQafdzchzdMCvdGmPbA1+tYVFu1NS2k3aupc+5
0cw+SaDsKKsweEDSPTBYfz6yZOMzJWAtVVPNfFq26mU6kra5mlxzCfAWGQKE0cCz
Xb1CpgHlYyXZZi3sbLqEciiIHD1wVahOzDyPCjgfBwB12JA0foJEnjMnU4cQ9R5t
IKnDUo6/1cEN1l6kJenJ6m7nfQI7YkGz+MKVKprD09Puwb3Ni+h2jYrwrx0PLAk2
hgq1YMk6wDi59DzsUyFexqqeF1AIQIlJ1Ts/cyajyEoSGG8tmcPKPaS9jkcC80E3
bQBWyt0Oi2SEUNBC5xiMDGSh/tQBF8cIQ7dKrPQBMSgwdKM8GTa1tYQR7YK/mJ1/
zcY4qdDKBG89ImtSt68aL3jNK/63a4+RGMcJ/xm+XREogNHXsXbc9ZVko7rTwi6b
ek7+UhGsn6tqSef6wIdhg7gzBNiXJH9PQRgHUrjMxD1BKXGJlOEHS6avnadfrcTc
gIexoiQDZl3m+2zeGvBbSrynMyAQDjwCuFnQ6Iv6xrELRnNk2BBQFTkD9cHfNC93
BDUYl5WhezHH1eBPh7XcZuuQR4hfWv6Q9ldn9NK7PB7hEt6y+cr2C9D9CLA+Syct
cpR0RD1xrZQ7K6dCQf0/5dl7zn/4Sw4BOlK6ZO4vyWFQBcyRPkbo4aBRaH3GHu0a
l/o3LrETv4ZsArRNDaXC/SAkwd80+fpXAxq1YGIabR84A8ayl4SKKYuN5W1rFEVL
A5USqsTHDWgs+1BKHiJvsQ5qMs+nK9tsdNCA2DEPrTmc/VOUZUE+bzWiJSVFO4Zh
9VjEoLq/6uJKcBJITK74cTfGwz0g+FPI0jWSieOg7Et+QaxEgYXARvJzzlG4w9Du
msxGUxu6/2jumNehoI9n2felQ1JySbK9A0VcLYVBqXL2eAEaQBxjg3bdblGeePI0
BmtZ4cugwsRFL/e/Sb0hDLqRMwOGjsWT5RdaBe1r8Sgkl5zMIFCJDBHhyrNARPXT
by1zSa8nGtuoDT1H+SED8K+DSCnFwfUoUC3fW2OuLTP1/IGipEkOnWTdM0WDaGyW
rLkOdkbq54wZYWnQ0YoKE/596ZTwn7SWlPBe3Ag6VgnWiW9E/Lk12F98ACiRsDEP
TjGwZat3GKzITU/t3vCC9cKihLAAqU6GoRBiYurqMFzaMzeZkpu3aYOtzKV+r7oP
TWyhxUoEQ2Fo5q/XELd+rzfR2yXSCs141dKAtrLMGB8wI629pMWiIe58T6KIuGt3
bBMSpgdJhCQt82c80x3znwHQ4qwbpeouanL117CxhY+HXzvg709EkbayWPdonroW
GIKeJmMvlMHAnf2HoPqZBr7yc/dLYmsKyXXHWBSB8tRFf6cGB5IDNtlLDcnN2ZNH
8+zDe3c4cqObNB78RVbhwwflv4X0ce0SpvgXPkb0Qzru58J2+L0n/7hdJMEqCCax
F3FsJdKsHY+9DcA8tUWACevaRgpkVe+K2yOwFRZB3qLlmOcib0V7rU1wwujNz5Jm
8VAOYIqJZQBQmxnnYcV+JKhzzrblDuUjc0NFMiPeRIKy9HjiKtZh2MFLO8b6Mn3s
T2q9B36aXmYYbRXSSx6SfzqL9yS78lhqnwNFc49S1amD60L8A8+xapqrBpghTlJ+
XWA51crHkgkW8d+0wORC2FYBrlQcOvtWRoaTkUGcCBIhM0IR2nrl/D03zDafyRno
m+NyOeqENFrs+aETR8jCiDzCiM62w2faIu1GEhM96fxcxKuWHrFCMgrt/gdHN3UK
6bVEjtjT5zrm3QsjEuy9/b7DkpwfB9OqTRZmIXrW+aPIwUEUhhV7ZUCvZsh79ZiS
GzXSyUVhGklOQrO6zadKCKC0Ajr/rGzL/OzwWbzNISyA+wiBV+xDjOJvkfYegcna
p2D902qgeyKaRU7bj6dOq1/uod0Cqj635hyhiFOR/cN5Ep/BPMbgh1s/bjabq6PY
4nwdolabWVN2G+Mfz/4HJLe9jKJgdHQWALAg1iIgHZ/CthPZxjrBIT4upbXdL05b
phr2RKcz4COqsD4nU8m1udJeiqQheRnhrA7fA6iEzhoNR1GGRZQcaIFlqieJOHrc
HR9TdEDNtU8s8al83xJkJB6/fEt0BErUOTw2/ENj3ic94CfBDJJSg5cHWDBsnvUX
X223f7NTnFnwKraB/vQNI6GsakUqXrvHYZXeIa6vKEFXMYSj7XYvSfLJ4MHFF6lD
e+M3LzCoqcZNH+GLe8IXk8Ej2qnnhR2/5AYN/gTPYEp5JweGdZtHk01AaO6UHnct
BtCSzk4ExL3LdCUC9BM29D22pWeJ+Vm2x42RuT76O+sU8CuWswVpINP7BoZ9Ffdn
PJoYkz7JpBKMH6vb2pYVDWG48MCuHRZHCGwQauoJ8OarhMzjQ+SnEa7ndL99N5cj
FCXW6cdsp3v7CE1Nq7eRCs7bfCABjYPWftN6a7rPyoLjSyNvH4TMfOYnwNxRcVZM
tmiOqA0u8hxVKcyvYvJDySCcBO+KhC9ksfaPZSM5VVya/IH7ORFJRtPKTJKgvVD4
GfxRP61DnbqXQJXJ2g5B7LXfAKC6gs3Mr7kelpwdGw3XJxgFJuMLFZ6qmJQS+XlA
qOcvBE6cjKPX0dNOnixnwnQ9HlQOHxiNbaFDMNYLNI9hrNbFCT62tKBs8XWa7UCF
l9ASn8gLqnSxUDDFBVMLvKIlp5hbEUNkrGVMjfSMN9WypBTrAk5/pVqQ1QO6pUEo
iPyvmTMDTMwwO0e91DMapvMlLZZKXm4c2ySCa4lzhWgJrFUgtroATQerCjVRE4p4
icdJIKqqWA7nv1E+xElhu5aRaJ/ohPopY851Y7EyDGKCWSf/pt4j4KBtj/TT2uQL
atOO/pIYJE2ygMsUB7ftlq8uBtkJjMTMS3NYRcTzrVtpMLiJ9OWaB6d5pR6fB+2U
AjSUyyHvHluoCQ/7+Ih8262v6HosewQ6V0DF84kzj4cysDpJRgLS392VYOY8RD8e
qMcnJvt8U0h5tKsgV6cdI3Sb0wmwjWAt9W87jkTG9LvqbN/HYMZiV+XDEhTKiRJO
0cerWTsFOqRU126dgx0ErMu+9psbmZpDVh4i1AsbM85Tod17o2MUixJ6hRCso5q0
3ukOtsNEi23l/2/hiVnMl8hYj5Dp2HYjHXiL8L7OLgzLaZoYUEjRcPnMJm1JNsIn
4EV5KEU6+8n7LHZAlMhQerR2V0fSkmK2WJDEWX4C22Z4MSUnhW14LEgEuhG2nMF6
FkSc/FvlIDdBM4z01nKUgQgH4jju3eYxG0cla0M55eU2+W616EcHZVt0LZ2/Xp1Z
oMXRh32dbNkXjQFtBnRFVo5z3IdZFZ80JwymAZfeVTuFRT23/2YzM348SaJe6yB8
qF2MnkVN3RYUel9c1WcyyLuqfV3CAa2o1jjcZnmWoYvJhb4XcAEKR3YlgsG+ogf1
O2UYblROMmKemidh9/Pexq+DVEwGZNNtUFmf1VQbNE647ZtT8Xu4Uq/fUgumQkY7
UQqlbzSHrrggtGK52F5QAHrNmdsMGDtaKf9cLCEbcIlSqocTM44+QBygx7Xe0yu2
kYKoJqCYVHcCe/Fuz5/ExIXum8VpOz8AR2BUDnyvqfBWuIpCIZpnqy420WZ6lGqA
kLl10tZLKVU16Hj7If4GhB/AcbZn0dj3236L1+76TVDH8UQNThdfbzA8so1lvgc/
cfGxR6RuNMtwyLkoZfzJ4/nnK5TatFvakbRGLaUEBQtJPNCM5/FI/jkd5OS7IPdQ
GVsOOBWQtNpCF1FNFTcKXmPD90nfaIjo2FFDHZlnOtJcfg1EbaHusHl1ot/0k2xB
YjMqdEbyAujwsu9eQwEYgAL4Z0e/oBiJacJGduhMgmM1uIBnlnJEHR2Z/EIWu83B
VlZ+Haq5b663sWYzYdx+T/5masBROtARbYlB+be4DaxI3QdxpoYtzADTkij8hGm8
RH+ApKCMBV9CYDacWu3IEF7sz0oBdv8mjHHSwZU8ldM4Io8EzrLssnkhXjUsvyOe
eDTr0uQODeVtc1n5oeI03RsCfCYvvGlhcc8XVN+aFS4LuMtU3qy0CNIHDzXmZPmV
P522iF4kCUCEYr8KchBGJKOKjT+erFkyAkpKVfKukQ23iq3R40EHk/JGyyXNnOvU
CyRpp3AYaKFqD+N9GxvdB5bER3NvWP/UV4esseUy/rZKNxU/gCWwY8LogLc4BJFa
/SQa1A9pjtCjlqzwImsTlzNJtPjJtjA1VWSnry5RyEQkMYMCfIAcD6IQWK9WxCZO
Bs/GqBqCFZcokBjvlwphxzVA2/X1PrijU0fh1Wy1g1LPj7wOyLKPs7qsvw/syZiB
NNRWa9dqIDRNnXJy+OJvcoZAILcXHfdG8X4bVqbggRRvtaDP0A2CKGx0oCuj4cHp
kP32qshtEih3Sdk2yTDaIEZS3pFMxKOEB4TBr4/JUuvUo6zA5r5R+U35PASAnUy7
NWQyU88GzGhsH21CZCU7QTKwNXuoY///Y/Mc4EzZmfj/dp5tQ7xlWoe9uuVjxCjk
THHJwB2p+kPiOTKStoWaCU4+I0NweMRGwhY20hIEVDCPs//Ur+K+j6qCp3qLyyKV
GhE76Bvj0BvhUMjYzhOTB5+i3zHEwGrNuyTpZtcciNCOj4MPMMAh4bJSy9h8yNaX
7O0zvLZvpN6RHGtsCefNL81G3JG6haSw5wapupIHBdvVyXEMIz+MfZSDCk2Id+SY
E8LxnbT6fGvATjUpZZoN7SubsaPrVwdJGtx+P17fS+nWMx7biuN5CQ6ViHlaiWek
Hj9e1CfIU4t/+Vo0hDmy4nBtly+DnKepnXNuwpGKJZ766h7fkP9a1zqLxxwMR3Ps
UrlmhqLC8PPvAW/Pd5iB5P0hg5G7fB0Nxsb0apEl3EGGWzU0FhzJ9wcRmFOGzXZJ
wjIUwnL81in0Nze6uJoOWqQycqVPkrAUjdM7JmLkNh9UhW3psFEN6FV/tnr93Y+w
U7Bfu3OmRVOMgESBh2CBY9NJZC+AqIPeWxJIzGqhF6oh7U8FCJh74mN+P2j3nhFn
7s9gU5LaET4OvVpWsj7oTZrB/jFcnT0XC3pFzia2PyMtiaYRVbfG2ic9wa9pyyVn
BszUOB8MK4YstO9Vvly1My5i3Tqiz53GRW4Qy6F/5umQXWBhWVtXLhjmie389CiZ
XTw8EMct/47aCDVYw4/FTRLhlpFfdKMZsDjfsHxUR9AiN+R9iZJqbmXkxlwlzjoi
tv1xPxeT6TttbZFWrbz7iLiEPcabjYO+YVfLzZgXXga5PfYSM5dqoHTpaikH94B3
iZznU2WuM4MnQyyrKKXdw22yd/VOObuK/Z+s5SJWl+umuW0oQ/ZyNRvndqtLkpS2
qd+DEaVsXUde1iEAaQxoCIkScL9RyiQoQ7Zft8ypKaqUBZAN1e2sFjMjIeoDgtGD
vOcFXlm9v/tQD9OMcWV3thxc/GYYpKw7D29BbhB17nvV0P4gpZnzdsTQZ5gI8feK
f7tnQkAp+XszHWbtsFZDmBpyEgrjh8Nccxd0ez1howN3gVYKBhUBxrKEsn7e4V2Z
XAXTebP/mB5rkrQeQm/pN2w5lOv3JyXvCohlZ9T9sQ0EWCAaUOAjDSE/oScFiXYP
v5Rs7ACtiOXdDtzSWB7sSwqW50QvyD97I3Dvq6Q/5TUwWxfLA0cwulhmbr7Ffr4w
dChAEQIjBg6N0KLn/2VQ3pz4OeMk/q5FS/PMHHIWeorDwxqU5Z9qu1/wL20BahuW
4R/UtDPBMMpkiSxeYOJjknScSH/twYg5qprklWnUnw2LEypG7TC8fWpd70UO07vl
UHjgegXQd+/rpn275lWrLYl6lgCsYA0hE51Tt1mROE30I99pTyblyMuDubUp/iaa
6EQwssC/7WXZurDABhhLogCs9QQpQv0GxJ4w1HCcgyCoSB3UwMXls+150U/0+9Mg
8bx7bf5Ksk78S1oQguMh7jprJFacsNpxAGjCZbu0jnJJwXZUDlV/kEBsnJJWFCKO
qsnVkgiHaUOKZZ9VP7mOB48XEdPoiHzaX+UBcdKeyHN3GiHaPYW9M3OHpRgXxylN
kvXIZk/CsdpUW3KbbxEzoQVZqnwBETQdooUt5Nl053/KE/a1jPGAKRvqwYqj6E7V
y+rSGJNcsi8us9ufSGHX5Dutfoi7d8tX8p66IukDwd61lqRMh0ergerdKyXQIgOh
my6Me62GYJl4urgGcl39VaaW6txnuxWQ2vdPhOAh6AifzOfunhOGfjgsMJw6bP6E
5HekSk+SsRqGIy6BDT+vLE4khuodZEg57XAophxoC0VF0zUeQ5zSsYCIt4Z6ZtJr
tj7gGrm2l1pfgdTufVo62FTtZgRcWHN2+C+LJRXjS2V7eMsb1FT/sbDhlLJDbkQb
1ihVSfStlbciKgY9ePKA7Cb8N/361lOE0niXdUoW81rZJivqCa5Y6KAB6TkExNZl
Uzs2P+ZE4OcONugv7H5+PvaVkyTUCVNn56p6PwFzUYUxnwCDJWlEbDGEt+gdJf9H
q0FgVAyWphpt2q43mG0zOmyNNeZ4UNyjp6HBFzRgoMI4KE8UviYItOWEQKh9d7W/
o0n8toijjFxMVMsb2B1MwHZ1lQkqMvEQYSBBNkRMBecZFk5qnDlPJg3LdzM0EgxZ
NwXqFtRocTnBkRXGgADElR9RUmT1HCbW5ytHJcqMf1tgJ4V4sBXwd1LEe5NFz7f7
jWMF+XrdCNThV3sO3LrVMgpkfauLids1NdXTU21/HXj5mjX+8ljwTxjNrfKNQUDy
7CTGtRtEgQUk0utFZpNmNe1zSPV7Csj3Pm+6RPmIBqmoetrZOvMrNtC5ZA72UfIk
t6RwqnGsiuNVY6dxDsfttwy//MyaFL09g1Cn+FboNrq22EzzwM97ELgikkNwkqj0
GgdYMLB9f5E5JkOn/W3QB3f1Ca+Mb8V8G2TwWOOotUWFg9o7+GRXxFfPmOInOAS2
3tyvXaftN2t1Tss4n6fAfDdo47TzZl8zpN9Nf4ftZQznjIh89pFnQPzMfKdSs9TJ
5ys2fbxfBtBqKHtRgHYySK+aPxUlMakPeDIxw98oJsTY2Rgg4hSK2rQMTE6L74sM
Nif4PtyBb5T4VZ0B+ZbJCxZ/I3G84xEtBwKyf2VWRY04wk7qNtRbFP69Kn6T5tK6
vAJO3q0WdB9x0ablfcezWXlVeBK4n78VwQytn0TKWv/ydUhicStGQvidBZz2Nb6c
X2P3DpHcKm1F1G8zAy2em1UQL6swb1uKeU4EsXn/R9EzoQPEY2gjGIh7WlF8yLvU
4gvr52vSiHSeCQ4HB5h82/M03ufW/GASxgwBM7VKZJUIfSC+gi5v5yzxkZZdYC3K
RG3P16BqLpi5ISDCK0D8Uovuwz146wWKNNTQcMPDMDcwNtYQCuBTmXZbGyn8ENgN
ewODInGmaWv2MK6srj4NANVvUFj1+fhuKxNVrvbYCDjxbuvU7t3izb8TvWYQQEdP
UAv1XcVhH7ZRpRqIM2AGbK7ymzrsTB6jkTDgZwT92KdaFQh6hSJFSlBMXJjZcJoc
p70fZTA5MLoLHTKGLlFxPvZfWZPg3MvTLW7RUBcQCTcYmLWRms3V7duWEn2fL229
5IMg6Dzx2PtVXE4ijqzMJ7CfXDtDD58gqc7ZRY2l1RoKErZTBtSKuuX3R2k8lAuj
DuXPlwkSeTjzs7VVfH8OMT4aQPXUIjWpGI8ya+VUlcodZgElo5C2oxpJX9ZYttOg
LBL908QB2rWbt9KT02x4UJ3U+Bre0qNncSWkAsfvYbeWA+i3B+RnLEmDkwQtj6DG
cPyuLvNb4qGUtXxjnYG++sLCRsl5wJd4uZ+GZiRIJKHsygGUE+dT4MJtcqZEAApA
SRTQblVQz9xe3bnrD9z2Z0yQVlMsj3YANvjcd4BMcBa888j7OdtIg2/isa7jgiB4
nLcxtRaFJxYKA0U2xeeR0i4Bslix/+enRaHWtdItr986SOQaojpcI7EA6tEDMElP
f3oQHYMIRyAPEp6QZhmkDysIVFsb+HYiVSgE5TPuTXKL0cwcNGftpV/JjaTCjGkY
zyQhNs4wEMf8g+S7B1mkhKu80Tmi0qzLd2i2GWwf/iuCWYDbEuQWyCRCJ1xb6eF2
BCY9PbdimQixHd4UzCpe8aqVe+oDhpUGGUTDWLUpjJtiHu4kAv2/+8CI3I/BdHpf
o8vFX5uKak4s+eV73fzJiX47dEVZWbJA0k6RoqiElyXx3FQJ8emZDjdg9b9sRXmU
+31H8uZQkd98kmsbgqxnwfWe40AY3XoaffZUeUSupLsHhwMLn0b8R6m/HKXzyQJ/
M7jbniQ6g7VEW890KZzMWKiMN1ZXGxIGZsSvIWV19DXamFioDoXBtVNpsDrEnLkS
TuW41AraDUf2yeiL72hX/O8NlfXeJURIojZqEBDAiGMeyYsssQHL3d7nuL5IDVRA
uRH1R7walIVUGElwShPcPGGrSVES5/PxuuFhdw6jVDRYfm+C8DvReQzmtE7DdLpq
Of2+XRK0ONJZRPJMalSIZ1PTbWR8qqF4DcZ6FkVXYnWLYxJmd1gZrCIZ8FHIBide
9BbbWRP4OzSwM9tCeT6T3L99A79Nn6Rv7jX/s3gU8qZngyjBQlVRuW5DXxFphGRd
hQSo3NohqbwDXCFyZxOIDIu5RhLx4AyH6EVRkypSBNRBHmp/saAlf0F3/4zzsE7J
Ji8zc7ezOCvFCh6Nq8uy0GueqyeGWdN2NZULcTs3RG2QeUrj0h2MuAu6d3i1zQLq
QunFD0X+YhN8d7Vo+cnhYW9wJSq5B+6OK6svV4xDFawd4RAKFdjAXoF2oFEpZu6V
xpZbrg5lBAXAvl8H6HVdtX6JDbtb4cLv2fvGn3UCk49WZGmOXDqWNfpB1/nk/wmu
+Q7OQSbyZA3ARMUtRJxrnVLuirlB89ejRNzqy4fEybRk34XybSn0Q0jtXGOtKbd+
HTVgk30obb+v+GXm9/3GVB0/F63iF9cj3663yKHciU6axnRInuWxxj9FgIqk3rIF
k2R8CVkIUZ4Dyt4Np1ofeeEzmbn7T22WIh05vGe03HnaujgF3pUnYO1PQudSRPDd
EfdgrluM1TRZZlvFM3FrR8PKkMI2MAhbf5BeKgVNF1Lmej+sOWIMWqaedtreNkIb
sXbpwLy4IW/9eYYQpONwfKbx7/gp0qUvdDhfdiImv3S1sw0eeJbLqxnnNwKIC9BQ
+qxQch4A0nm1SL103pHbsjGffvPRwDS+xeUJyBGLJsSvrpVRjzqUSi8DdRX2uMdW
mj4l4gef5f7vi9h2fnT+YUrsw0SDTaZGzVzeW0DjVUlApxFI9rNMVv8IENg0Q3m/
Us1byAcED5NruaywRygJ48ht5UTLxQGpzqvRiU0vVlzbLccpNvLqfce0eWN83bcp
0cQsSI/z5CfxheDErzmIO2xnq3J8+C957r3slGNAlG/NB8d+NKwb5AC5MM0w564V
epDfPOogPnm9kovs/+b6sSx5pfp2rgFcipahHriHVXlahZpfUVbx4xcmA0Evjrtf
KjFU/6Ou4xPuY8IqSrV/IW+VBcxwSfCCNtYjhyyAhn+EHDECB7KTc7oSTatzNRP/
Dg93ZQuiNRCKoFSxeZNHOF4D+/E5NmdNq42C9KnAHtfM0L2PGxWw8p0UoKEi3+M4
uhcPmkMLqNRUzVUr4Dn5rnqj8BLXp/4yHBRY8uTXaKq5NAf0boq9EuqwwbmISwCW
8cjKFuxKpFtbkJLNv3/uGvVMP6eAN88TLEC+tIHL81QNhABuDn8HTZDgS+s1Brv+
dTp7Ke9AByvu9YF7g6H39h8XGAaPNNLIqZaoWtGCgWazsYnBFiYFX6fyrT85zj+k
6PuZgw9BDs47mSk3mvyuG7FBTe+miynNvRi5sLz9lBtzCz53AdN8aoc9RqyzjWRB
qdKbzlEiXGEvPrICQeBx9gbbZXHc0Z+WBgpZQkPDC0j9G258l3gk+1ZcgNlxGD4O
XZJaEFgdrjYh9VeDtTow+ka0E5R3JaAxF3uptkzZzEy+phSF1nx4ztyGy/qmkLwl
2M8cd8AjFo+ALJMbawZ+A7yP4xaNFLDuOh6mEuZitmPhGummhfrTb/pVzZngfmPF
69YQgIMaWsSkGZzPBmo0xMzbAKSW2mc7+Lx4y3/z3w6bNxmTIlDzk5WJNP/vVTgC
+JMTcsutHXLQKSSXkkzCnT4Ipp9rTQvJIQDIpjQ/hdXvOfb3jOnNfQk77P8QkOQU
jOUZo1kXccVNVCJL4LO5qbIzxLgcnlZnNR6fEF7D/cI6yV8V86SJYFL9gkQsZSsm
XGEpEedFLurW4hIIS6i59+ubf+00734KJabKjqe/TFJbsmN1pwopAHYO4j0opWji
QsRg+4yqfeLh2pHHOZ66Wa34QnSUqu7XLBrg6iW7JFS8ixQtzi+ouzXo92v4nSVH
Ro4lfis4NkrgQX2FyITv/T/DbSk8eO5pB7ft14rfvHAb3pwC61FLDyWybym5Bxeq
TcnvM/2i2DvW43hV9tAmPRwAPs1D3Dje7YX8LWWGEsIAmMGuCBQUhPa+v4CUWypk
ovedlE3XLV2rwQNGNDbVtCHgjGEtz0Zxj0UyRLtLqp1dDHt3k9OmEb1jI+TpQRFC
7spAyTwxaDvxytC/vSHwonaB2zpcEgaG/yR8u8QClaQGpMkGDEmvkQLadGFTxfDU
7qtyahoWum87MryxAt7VIe9U/i//6/D8a7Ky3RJyW6/I3W6/4GXWHr+uF4dGhU8o
H74hlYBQWICqMJwnZUxtLiBDf1/cs9Tb34yEpdx7RHLj7o6b7E3VRjGyJFzmPV8y
aG74sg+7OIa4OZM7YvAfULvjAlOADyV/u0egw07e2hKO52PtJAA3qzngAZBdqLAk
DztnO3WU81nOMpmU/TAfhZOSQArJVFRATXrwNzObUYz+9P7LoGsqhX6kyWT8AGAK
sNloYN8nIZH33fgeoUy8oQTrQKvpKca5I5znmaRtNEWXJdQnR41eqAwoo8g1zCKh
OQBwhtAgqUqdtVma189QaUZzjW/lyf+jpAJcGCUF6Mn75rVXMQo3oljFKwCSgH83
3zYZPWtXxNLfASqCSardJPDco/+Y2CoS9yFBiUhvALI8EQ40DHu5XX6rgpQuCu73
7dZyAXoD4lTIPLo4oj6KdoXV335IYfU0CbMhs95YxdSZq/iqN2BpZvIsGCfWMpVa
SYWEVomGuSWJ6a/AyBQX7fU/1cIuyMm4n/on2IG/yB27CFgUWWfNTyuTo+CP452i
fSVFwkjeL+rmdgOATfrlKgU9l4K/EZSpUsd65uILHXpwE7nrUvXzIgK3TeV0Ap7f
fvXVqI9vHkbroFkgvDmOqppm/fzv6A65lXEwOoMB2phNELNrwXuJO1YQ0QdB97t9
esJqk3DJwFN2daPOrUD8YWy6pQl4yj1P0DnzTVzkoaW9D0BOf/lCmE8tCKNwewzt
meq+3ZV5sE6EX6ZzcQZQhrGqURZ+3SjERXxGH+RO/KJYPHejmCIFerCtUWi0Kvmh
j4xvaTA8LVZmiBFpCW9PhuYqJLyvUPjC+vsFppELJYRn/oxp9XZe5sMNGP0FgHB5
6dGgmQyRfFgWm+5Ij93tEiCAoPr6ZMnsMUwuL3vpYQacoNOqYjlLDGwwCIL7rqmO
MgFlfBBoufXlsoIBwu0Em2MYZWtGW+ZKBbMPLZoCkuiDVu01JI0kdF0/EuMbLnSf
8y4YjRSaYoJntRijzjMQT+KcDipmVyRfXUaLt2KXVaRGVXnA+LqoAJezxAnn1LId
eqkKI0NscfG5d/QODQzIj/0r4/2Ak939NtoNC55Y7HjQBF+laq2JFcsb2Pr4CXAu
Gwd2j+33yAygo2yVyg4RMJFgLmz/jVmocASzdSDYBn5D4jkNecXmmhmrNjUWIK3z
Sj8XUaB/hJdjRTKg/P7qR9iIAMY5diCrP82JEpu+EXyNkcd/gj7uVanrmuiy/8eL
5m21NhE1Yri2z2APc2+l1WWYFgHSEamrIJGlD0lkiCoZ6COn2hDzJufO/iRRyLoV
8YL5MiJBzFZshN5K2D1jKVSF8daLfqAcgLTeepaLZszERjkQ+hDifUTjcu2ri32L
gYGpH15LxAOgRr0idK6xb3EgXvkQa9oiPDCWdNocUAF7yRe51al3sP4aCAuRw3yj
X3S1F0yXqA/lvZcKNetX3I/hvB+/O7bzx5LLbFE6fD1WraSVmRBVO2s8csIf1Bnb
hAE0IyNln/GGty3ay6JdI2T8jYmgplIUM8yIrmTENCTceljHH4OqZQpzjlpJj1BU
+aGubk3UeewUwgGQLq9lp6lHjeDw0PaEdKPHf1XYu1nBavYFeeou8pi5IkzfjJW5
BLKOWMdvm5l0wO1/Ms82HwJKYRTqhhBjc0Fx2NhmLwXVJFES5zVoaoCbpOSqpaDw
Z2uJN6ssPZrXAJGQAW0qXBmuCvXdbRAg7uM9y0rX3ituB8RBf7lwLIJjrFXGLtN7
yrsdqpKVjiwcsRdYGPHlFmPgHYaDWEo3RBWHiRfERyyRybL/9ZjBr9rC9OxtbG+J
LPQRMWf3iQPzLckhziSUkrAzMWIC8hMUMZq9q/Btl8bl9wXG3GG98WZju30SLKdU
psyxOZFvdLydlOqX1Xc+qKr2dmZsFvjgBQbYM9fnA4AhQSX5Z5uN8h6RalOKNz4a
+q6x2hDOO6+YGsAdXvyAB+V+nk9oNSYaXrP2vjDj/EcwLNViDn6kx0uyihHuDz5K
NtDPl1YItg8EDrOZ/GUzih05jFQ79zxTEZPgxUBTyvPSggTNxMTgCg1uY0WAcwZM
ipfy6e37ImSH2EhOgVCxHooxZeylH7wuab2iPV918IXIo/ncZCpZpz86OoDt8afo
Ob+y73/hdc4/cOX+cJ3WGGnW0wAtSPoX/VQVsjW9/sW/rwBkuKkSvg/j4U8o+aqp
T28hj/Awpk9PyhfeiPmM9HvuqEM6ZSbAXO6x1vNQ+OEHBgepE8ON869KdDkiSJdU
rXRatuDfDRJu7UbvkFZNVnEa5nSiuYGq9GwXReS/Xw2Ocz+240KYAWHs677vlrMA
i/YzIcHwYyiQCiAfU3Tj48kgwTE5mZP0bsZTj/Fn5hCcEE8Z3XPppOuCJGf0G48B
pB/czTKHeXDeW/jA4XvUJ97gUDTHn8my4jU+7usXhWVTQAa8n6VXca8WrJXR7H+e
4YfRCEG6jxvquAlsuJ3AjajUeiPWhWMiGUU11FapM/n/50rjesPP0bbrwkQ47wFw
xHYfPa9i4Ht5klOIQulVmIZK9uYuY562HT46WbzsEYA9W0M8GcBfjUJrK5vaR5Sd
Hc8F2tP/ijcABYCxfkshK3+WkB5kGN12AbtcNN0zrz+P+13qoRDyaa9zR0ESCnwV
aBlhEVPdTH3q/57R6237oeUV41TVi4P2u8xxg1sGmWtFdTCP21IinQdfCKYYocgj
+Rvm00RlBsPUjFqZ5L7qmCMjPC0CZdHZMqAWThwO0gOO4IT0rdWfmrPFVyFhosoY
JM1cP6f5K6HSOT9qtEQH2mItFxzroJW+6/yk2WC9XN1V+oJxv5OfAiCIDyeNIrnC
PtVnP9GMWnLkoSc0L0kCY5Yp/ja2Ixmc2TrTDOYyiWxipBErLt7cbleLmdit7q/O
TNSzusOi5FcYXHmil878p8y7QJkUnID31FCoxR6iE7L6crRo5W1GSQwj+l8w/6gc
yO3Hr582fDo4gnesgIOFum5bZwkFJib+z1ibDEerQM2cV062S9s1kJomWWXxW5GD
y8/JuK5rHvt+LDwTTWnu0HhHPUrljukF2EAZXPrpZoQq+klGQC3Lo7FquKLlaZKa
+DeM9Ekrk6X9GdOUhrnSOWD/UpOeCr9DW/GGbGxjBkX1Ho8bl7kcusOeeAo//byE
opR+/U5Pt4AlsvDpy5Kfh0pSoTvz6qd+155X8GvUNvtH8NotyI9WXvIQlI2hctHy
DS4mw5bPwVEC80jZgP6G3Dzn8wnB3o13n+Elyhs7RrYUzDlcjGYmIzVlgd4w1ZEV
GoTrkkh51t8PXXboa18H3eJ55JgUT3g3irvDpLPuk5xn48kd0Uhg4ABzdyUoCwyy
tHqXtGE5h+5Wm10PGAw/ZFtg6C6EG9Hfl5NUPIzoWDu3RNQtYBeiKRGYqSG2QK9N
KWKY4xfX71GtpDVmRhTs0OWFOq8wNHtZRMFWPqNId4aPN7WvPR3Hke7Yq8v/LdmE
fGuPXwpd3AvH6CvII3YxqnVSAARCkxwqNa0w5x3ShBVCA0inOVi5rS2bATg6if9c
HYKyVt+pFspmm6qZluo48EB0AuLU7j4+eAIXfU7nafrhZPc27/HfJ3wJvOZh5weY
dE+ANGTWASCr76bHNue54fwEwRI6pkPT4mp5AmsYYJ5nbHLy5AamTngMSzuLrm89
Wo1iS5VtZFQzAk9sewvRqnDIDDe06H6VU3GAOjIc5WRNy+JRDU6Gdl2UaD1Sjcsi
IQqa7OKdOuMUAaS9BDeBQXPKJFHx/PkfqMtdJPo5W6v5p0lSpE+RPRuFuehz2A+8
Z+Ypev2vyAmN1hJFNuEkJ8YVxzrosZrkb8jFG3i9s8GAnEkZGYid5yzZZNSgOlPD
vYIbVVMRm9NnC+Bj5mdgumXgTO8H37UrBZ4KBSmSkUHzxcQnIh+/QtYLKZnmhGFI
vRjo5QkiuQZVof6ApkVkdxqSelwEp1VRhTakfuC4L/1IIezjEPWXAaMgMOPx+3Kv
7DG+wWUCON0OIPj8hSqBL2VuxLwuLkYgE0FR9cs7qgl3JvqcdBP8ZmpmbYHbNKma
ba/sYB3TzQYlNoaO5GmJNuxGZH8sZ9On/2AmAt/9QO5HvcezEHjiNhUg1vTMFGgJ
6TgpwWP6Bm0Lhu4BG0Zgiedl8pMvbkuBq7vz9QL99R+vD+d+L3mtzeRMBIYujKp+
BvFm/f+8y7iH2cNfxS+sUgLuntF5BUEz+qRXHK/4JR39V5ouu3oVL7pWRdO1Pncg
97Qyd2keLRp6iV+udHM44BHz8dz9P4LppVHFRJR7RWNocp5YflkYF7JMA1Of8Yah
N5e1v9x+Rep6yS+BARLz5mpRx/GqtN6ZCOFXXX0+XnUEIWiInwaARp66N8QCI8hG
1cgTCtZeyDEb0ypb6IjGYitt399e8ruqKMMv3073hsRbz8VSEe1UKvxNqJbyUnfe
u3+aKjDaS1UzZN/awLJpn1B3yOCgkAmdsW7Se/4wx6FJVyXeputRNa4/pAygiV8D
y7uKyZkLB/STXKnESU6PdFoms5pfrKbVg6uiVoxVD7LNMDFcXhQaVh/wK/C3zYMN
t885h+8Ic2ciWipaKenxQ9vdOypgnoGNHQavVM68YVUHBEu2+Nqy+33dE3zIV6vT
+pet10auj0jTg2aMJ9TdOWT/5bm6ptOljTTLIgDWiEgc6+GPojduZzYfrIWr5Aa1
GYoAnCpZUg1wjLXCPgHc4yOMWwEaNSs7bigBfKIsL4OfhOqTXTId9sodeR5HSck4
gVaq0Xgc5hJJojLwWTNU6c1QVQr2NJ0CEF4T8wwk8AeCUQIxOtibZPH0Tred9iTY
Zr/Stb66VOTab//yoeGAO1ePiO5PGexuLwuszwy5l2EvhD33b83EVn/n6dXIfysN
f+2FT+WVGpmd/fCTq57XaaQxKWR+PWC5YyDy39/DJ1ebRRBezxH1NnkUIF1UujqH
ZMoxwPvHn0qEVJ4Ab1Sk+WwpLZpZZePAkj94T78pY6XTC+L/iHbi5XmLNk+R3Qsl
LnMwuthvWaCuHaeNYqYG74wZepXhy3YUBUNVtGFhxuJ6xijuOTPugja3ucz7d/Xj
5nuYv2A7Oq1TVQi/g3JZ2jQsObOixK/xR7qqObpm8sJ9Ixvhl0faHEwh7+qmbZ5K
EhZ0P2UStLgDYlxiNSczll08161j1dQxkwpPoldyvtg+rhCEAhROOqG6x4UDOYt6
CRgfJR+Ml1jLDKEwWL2ibvnn8GZuIldovysIg08A8jqeXIvppkPRC2OYUyYw2+xY
PvHuq9tmFwlGTa4mnq1xLJw1l8WFB/uwzDJ4ZSIMA2fOfXR5qMbq5/VWtSsN6FBv
cww7WTTHIl2O6+gKoYeVI4+6oMshlZRS1GX8lffZtKsQ8ITu+f7JsV7IQCRuKmYj
Y97Us2ix0rccuypEkpJ7d43jY1V9Oy6nUr+3vyGvSQc4v84JtefI8CbBhqmaPU9/
D+NFkAJfUx5yVA0t4GRsWQ4SnyJcol9QB5o/gkfQKwFxdriTtfCdFkcRYNHsxxPn
ujlJU05CIJhqTlUz3uwHbSDQRgiNzJfJkyQVpRmvGxukOumbWODx4s2yLZcAMxgq
9bpG/Rdz7UftpxypGtoyntT9yW1MlKUa2kmDf43az1f4y62fZTvGb1JqN+6YBEX2
puby4DoluiPb1ZZIo0XGaTObkoH7VhQq7WczuYuKmM5AX62GRE1F++NwSqFaace6
aW8AXiF4olNNb631fLCX32KOZCduRpoILaR64yWh6T51nEgApovlzsj7M7NLGmkm
imWNwDpBIP7j1qDg7jRT0VbgObb5dqJ+M2Obq4KjeydUSB3Hf+Ga/Gq2GSyKNW0Z
plvkeNqRnScbeB6wJHgQngY1ZKmy6r2qa20TErJFjhmY409YyFYBlDatCmTd5nTz
Bp8ubDpxI3ieZe2aq4sKIhOoQ/Cwr+2k+fEF6vBOSjf/moYTqVf4wsxWheP6OXaO
8tGaSxS24Lvwj9d212iNfkIjcjhyotjhzt0rNl3afKhQ4DhPevzpwYH8mY8kppG0
pilOrSHksmt0bg8LzSy5waiOOF7jnpj8XMJPEbsCaG8kw/kqs5Ej9bfXNgWr0G/u
iRFrJZxNxbYpL1/Dszh0IYOhXXuSUbXBqpuioqPX8xzUCS1iB/D9fRgjbgOgKHfV
ghCKCbD+zcgVVyoETkSqiJsStZvtz8HVYJCZ/qoqozevFQlm4PRVWgDSnpd9+ZDq
nDDKAd3xV3L3z+sUJlOCLrxofofswX6hkKdPuXq97UWNrj7ALxupXMz/u5IefaJn
E63e6xgvqIhpthNwwR5GMgBl8zmk7EENy0W2hGxra0he9B2arJr3hupiBMuc/aqr
dlingXjbcfuEiD5NjvIBhQskq/+OM3M+ETGwQdfLcGsUHgWdRXHw499TzbKNmcy8
fz8m2+JGM0yt6oaWFUmHv4M2v4VP5wxzFkASDla1RaqcWYuRwKlY4qsnxgm+VIdO
dyKHmuGawPnAlO3g5GvDSO0a1MuBQyLlhS8VoGaRhI+pJe39XbnHk5Q1ByF7duzZ
R78QtDUdm8OYoJV+uOsCLoFpc/bFissEXot8WW9KyYD9sD9qvnAwn+aHZcI1Mnrw
lAzKHe1cHmNtkJDm4LoE3Ah1l/XZfFsHvuxTt7pQ+3OfMX2Q7sn9ttjc296cBdUm
VBYFly6DliLZfMWoRx3eaOcgjnwVEhVsWM3DGhaU6Pjie3xnTXD/jMY2iZLMfCel
iEzSg2DOuWqR1JNUSXTGo5i4S8gTDn2lLSYg7e6/8YRVxbFR+j4pjrp65CwMoJPd
yiiyndzH2k3dGMDdxgM+BcXjKy1g34B/w8U9P8NIhrejYmftRXNLQE+4qM0ZUKac
4TxPl9BC1juUd8n5G0qO9ATP4pp2/vYuntxfpKCoWp5adFwTdIxksqpBRYwaourp
BcROhpzuqPax01+Z+QgBFoGf/IVifadl7F8tmauMCppb98cAT7hmeYBmUcwb+0go
c7bagAkMvtvm6Jjxy28PK124DOYqoGGVczm2Sj/jLRQR1xH3ayJb5dhEaJLaUQg/
ijciDelquofiB9GdcKy8DdTuKv8zQyMe9+LHMd3FRjMth6yskY5ylRay3YS7W6nU
FcM2xJUmLTwuTIDtpqTtWewO0N4Ng7Ayjh+HtexxaqKrJmtMIOn1gDwL78DQjE9R
gW9gUr8EyHqxJSBcqYbJXMfJRfmYjaAh2xj8AKr6pCfy/PTYCkkbT0k1UYjHXg7w
C4dA65ejJnqrd7pfJH6Tlm2xX0Cx03zQIOxbVcO6cTVl/EFcwGGs1SVgwFyjL+vp
59+eXx9xL/2ELrsTyHhBiU8YfpDRQyY5g58UEhW3dtl07B2Pxk2H5DAk9YPbCl/E
+rB7cWlC5P1ODzvcthENxl1+BAjFXkT2lNV6JuK6zRkYrQAVq+YuizFgc3fPho5r
Z49F1EgbbNts39Nfxu15o8WQD8sEf5yPt7c66jZXmZGEq6IL19Nv6GBLXhyxPHae
35KLNzSdJbh94EP/7QqtfM3y/KNmZRaJysl8O4uIgSKf3rwRA0Eh8mxyXhc4zNgt
H6//I8DhrtzsRgd6JXJgWZ6loSlsZwII1WDuQQ9OwXB/jGxeADCraa9ZucTA+Www
QK318yPPfwI9yVjjelR1CzivOBQyYGUKvE+wQziEfQ6u23FpOPg9KL6C6/4GLkEU
CrRvqtneS3qmnp+60JaNrNDfQZ9oEbwEXmsUSxLk0OENIBlOyDlJzED8VMFou0jN
ZoVuhWRAtBbsWbOWvSgNYOMFHnYgsPnXYJpRg09iUKGUFpNBb9+zmFysyxoWLB+t
egsfOoizeaVGlcvlfb5tJHAfX8LhljdIn7sH6yw3Q1twHnsBNaxFft8nmt7gZXQf
pUcEby5FM5kTBcKKxLketBLdidPDJg/lAaDv2H4amRz0GTlkvTpaO3S2Z/3f0T+l
5jwgFrQ5eegYWuFZhKH0MH6Nml8St29d7VEKKJgD20wyZ1TzATyCgJDjLBAJk5+x
SkjXlg5/Wg7NpO1UkS2Gxt8+mYMW4lT8fEUHx+IBKrTgoIp0JR2KOfMUkRdaJJFj
MPRGcqJts6vJOuwPBEDFcYZg7BD86gBKFkIJUlj/YSnayLNWG2ryfwZxWm5wj//p
2Aui+d4EdRuw33Gr69IXHEesoJmq2ryTuxE3R7sSCxNCYagzNE69GYiLJFNEnGxf
v/L7GWGZLcDZx9an42Ciy52dxyhDEFbg1+mlMOIshK7rtaOYe9gs3UYwaoQ63USv
swxYs+8J/ca12oLRgn3voTRGOvNENJtw+9O7FowdtaXcjd+1efClN905MtLXEW5t
lkbdlbOpxGqNV9JISdWKyVyY0jCgSkPRs+a/SHjjs4lfkuMvWsoOKXaw9P3B9MzD
SkvaagQRz2B4Z8ZiorEkK4mPcE1a1rYGHwGQR7M/M3FitUEUHry4HYwjyKlV46D2
iif9frZ/9aPt0FzpSiWFGNI7GweIEn4p8cg8FLjkgTAC5YH5iwHIJ5juND0AxbhI
y6fLjHmDYRHPeIjrJwq3CiAMHkkF3vTlZG4h7JuxMKEDKPMA4My/2BKocUJRetdd
H81OES2LrXDzcVjHolKkoGhr3okeyzawkQoaf176iO8kprLEUrd5HJvxsqUo/Qia
KmiBzu+juaKJx3LzUoBZebyJZQeNT+ZtEqa8xstWlIYqQZuiKEkp5Vp+yLwXaikU
eT4tTZVOwndwNqLU1DFp13hyLwnRT5rnQJaIOIPNBWeYe7h2LyDPlg/nIJUjng22
uiYAPrcxEqy1QmvzDQfdesUIFYNl3ZkLbGPdrOycE/4/7NyjYCGYTkzvW+oNrfa7
C/vd9Fel8NQJAEY94UKUCM6wfGUMmNkQX3lA9EevYGLF35MaglIlR0WCQke/vFXq
jAzqwVtHCEtAwohQClU+m9+lT6j68GXuqe/rPS8rKQt2vh+X8UbTaJtvkpTtLikS
VI7jF7UJ/esUYWKAbCWxuTWzoGIdzjohbkYsTLs+YpdRF5MftsM+YAB2s2C2L07J
f0DsL8rYzOWOqCOE9BN+YBV2q2wGxl0qIHXr+MSsiKL+daPinq6jXirLpgfcE8VL
HMuQ3aaJymzkNuawALmRCxh2uxIG52b0I8JSeDLeY/5xxaDyhewZEM5UNR0ZhcBN
YmHhhWz6fwUlJE28Fvv/pFgOYoEzv38y1Qia4LYNC1eDt4RmLhZlZR1oAOnJDVRh
qDXpXNsJyIooux9WCFTr1MVAbJGAYUkZEDYLBEzNzkCuMMpbm8DnfVGGCJhcxiU+
tn6yrUsPrx/AS7d/KOYSKdLKsXUF1nDkG7SahTGNw12yrnEgdfMVMXXIKYzsT8sU
9iiFq9YM6tzl63ssmNIp2JqDMcW/JZUCqP5gpQINIq9PQtA+niuODx0a4tziQTF+
cdiQXMzE0ahLTMVBsNHctEfb4GZmLo2NK/TTOInWUA8F7po5b37wtmK1lmWsYanL
39rHwCeGpg4LCffEzVFugUj/hFfmJv6J9vGmA/h3Kzk4MyWm/ISsw4HuWhrt5/h0
BfSZCe7fkXgGvzvheWLuKOizQdaeznEUhro050mY8CV9JQH5HQ0/1CD1KDl7jx/C
wRdcj75MIBfw3JZxL85mO5ZKjyQYXytskIUZ2NyXw4oLeHyS0ybl/IINEv40prTA
WUtsVIh6AWHkRyR3yK/pNB/VdnkkdXZI0EMdZFijk2PGyegGuiV2jiuqN18wVLGP
NhcDZObXt46G3z6Y294JRr/rxzN+dUOAmgLLpgAxOMgGHRWy8QLlLADhKZhUGWuc
QcKD4G8++40LqEDwhtkLCAJMndQYToVu4Qty7DlCqDl3t7lY3QadC4Pry+Gy+BP/
ZtvbjlyROlxqZIgGocB/yO9/AYvgm1EEJnJMRGDjVG7guzhHq6BNFkOQj8OFyXX8
Fc3u/D6Hjs30s0b4Wv/msCSdFo9llmGoHWV9YQtZdNf6PWm/5qhFgFgTW/t4ljik
huELeFqDLAY2h6mmDJ5+yNBA2PUbk3J4ZVNIsc947bRFyCh5VmWMgCNe1lKKLRGH
oySWP4iW7mzTw6KjXKUJJQcrS03dr/obeztXIRbDKiVTw0CE0JryFGSFkAAeMnYk
LTQ7C6+LsIqqfuOVEVa5s9SPPZ26wI3ZGQD2Ol4ocv5D9QvobTw2SVJPNT7o2KVi
m2WCgrcR8b9W9TyJA/JV1eHeZ1ZkNDdp5CD2jdcSXGyHO7qUtAI7LnXstYdvumdY
QIrLf9taLwYCN5CoAJd2OQXKt4iVwswOQIaJqIJ2wdXMA5F8LlWNKDkEBPH6I0CL
UeC5EdrDiog6bTQVSk0cgKyed+T5dtO3X5HvRzINlV2BSDzzGzxA+Jbr8csGxvu2
u+Be1iD10k9TeGfvwNC6xHZ5tmG1RSV3dWpgAP2JZ9T1EH5v6wGd3BxFsTpMriy2
Oj6irPus2KdQjcXWEbr1PnxhsFLWkSoR+cXxZC0W3Q0tlME5K3GyHMP6oQai+BHV
SYKXufdRxeumCaRozRiQy0LQP/6CHrJGG01APNp50vGgNFmTRpkrh33xeueYtVNa
FGWTKL/041VITDOOSaTIF7B5x1EB84UEXCWXK+BTbHqc37I8/bfPS48VCXDrD5SU
JvmUXoZwzyT2QUWsgzfXzKbq1THiG8uqoYo8IcBpYdji1nFVKAUWM5EOqYrOD84X
16BUPPqNDJU3Cq3bai8UBDYYCxb59Ey48tKLXMEsHF1m48XgZ0z+W16Ljlav7Zou
H0jLd4vgR4o+B8XB6sQYKOZcRal6bJWc3/JkL/m48gg71ZxjRQ6iRYz3lcLTwh1P
TwWMnLi5EHcnUQosGU2S0fkiVoRSzH47U/8R5pB30GnsxEmySxDy4KlT68dpi7IZ
z1K7PeNbwBUU9XBbV/sM8GkKUAAzYZNlD3AZBjJmHmp0i5sP/G3aleXuLYihzgmU
dsU353VFOYkEVEqNC5uZ3vMoRv/In3ETK/j46t/tWJzDQKhgVp83/Y6pNTJpiIBx
c0AspdwtYzdhDfc+MW3DiRAOqnw9X2m1tJDxhMqktqI3/sd4Dr0kH5N2d3ZXTBjl
nQQ7ZiYz7EV1SlhYYEo+4UbgMiZINpAUbeaZCQI10tnfhBKIUQHmmg9myFwAgJOF
lyll1N3xO/8xGtWQ0z/AvoTh7nMoT/bVXzYM9mnWrR/WBfqmMnrp3H/E7T7XXDND
/GmSKNZxKqC24Vh22JB8w2K913krXLiHPENcAWUF9KzO4uBEij+NUrxz28K/ve0r
aH5/fcJkwUnPIxRxQXMBc3YOLirL5nfkIEL4l+390RJeyOKutNJBTBwETD8B2Okw
IS+BfMd6imcEis4iF9+s0cVFk7LJwMIOLFd0IRwverNujPBtlT0NYmxuj3jCWGrn
02mYfi3yQO+mEQmxk+piklK3WlFp2NpprXp8XNoxFLaFI10Bb6g3u0QE+r9Yh2Dw
+2c4p20bljhLDBIAMnNd27rhrWAKLIKWYxO0LKUuofE9o4CNhSiyMCfTfe3mT0cn
W0A//1P/MECLU9y+LvxD0Roi5wOJPKuIe4pXWu8D+Y2CPvRammnS4iacw7AHej1p
NoKVClrz8iiyUnTP4r+1Z6HKCL9uCNiNFTenkz2FidtJCPXDeus8uOp1qzbGR/r7
VcqJDKBszTIjwkjPoI6uYw54T6B2jgKEB4zKt7xtiy3Rwh3vwiIbYgNb0MQlNw3o
7E7oAOscPV+Ghb/5jvuS9deGmrN3T13pZyWuQc6Zgx30KeQ3IaHWKgSfM2VZcpX8
9IB0A65xmB9y3kKWrCe0Z5riJhBQ36Z+pa/1EAJkPZWc0skOfYv0kKS6ly55+NS0
GGapC93BsYL4JJyvJqGhnM1homrl5qKHK2pzRrOUDA+2JeP3+N+hC5mL97nPECvr
+zrPDyO9+RE/wBrPp3jbGYebwKkwAeoHbsLc2ww9RqPXyf2cSMDj2ifgIyaqe0Ty
sKJ+WlyOqkXyVIssUZECHP4phYeaL3IorHzdXdRaD52Kn+p9q7q5ksoY1Fo6bnVJ
jWQj8LUk6yVKQV0HIsHnIZryZ1sdvjJpUFFDoPVU2d3cTR4lJBiv98KWouzKBRgn
/ZZUxdsPdRVi3RkUPCzHYxoZFrUo3d7dh/GIw4ZzZvH+4aUwI4xwO6zqQAlng8QY
d/qQz7oXH29N1+NvgGL+cyJBGrHIy+dXRJaZsgBZVMAsYe09QLoN+V/pvbKe2pPB
I7AhFV7scc5Xr2Vr77+iy+4RUtkWyEuLI7DHsIX+hgWP3rxGnmVt1aq61SEnidfw
F7RTFcc+ZEkNpo0QVb04y/GipzfLVOz0Hs09pihoPznbD8fEneC27P9SLp8BCqVT
p70FFDGGCJQuqqdbdN6j672J4MYl6GzkwXYM2DfvIQ/IHRd/mffQ3YUaRnh5VyAI
q7LtwuWJq2KKVxA0VNk0jFGQ+71Jg4PYDzwqhRYYJyCwj0siL8f0ZsKdz/xgmNja
H33JzW1QGt7GScXUbZkEEi7R6ibk7zDFhDf5epBxfvlBFbGmJ7wtIR84vfevfwZf
j7nyZ2z3ERp4G6SuQJFtKga2Mh5mQPMaD1jlBtD4+knXlAEkuwrFMLpQ60SzyxQ1
VnpP4PQcSpFx0emUC4DQ8tuMjcsKZ/cdgYMTCY//KeoeSfHKUaLBScbIhONRxf0C
kNuNa+E69WBCaaw7leMPaShdp/emRrMGf/BnoaR4CUu2meohS2nAESXfsGi1Bgyq
8zWrxOzV7SsrNc5GidwOcxB8sjRj6E5f/D/w8UFCm31opzhGGh2pokOepGHoGLig
cr9NHzJYUvlK/m121MCH/12ZIU4B7Nvkdw0oeW+r10Nf3/Skw9UEK1BO7NDkGcBk
mXIBls0hKZGqeqcZv0xv5M1XoC8CzayUNER2RnsfRw/VdkLwBf2RiiTmPDzcjhRQ
kRrFNK5Z/RAhpvD1mhyko9iKYrHyZ/qZY5qREN1la9uakD6qsCo9KFEATB8ZKoyc
WEuwbMVXaopIvg/xVEFNJXRMBJhVVqiy43VmHiyM629q8bJVW7761XY82wTMHk8g
U8SafkUp+1wgBIgXonMKYviB2eVX0Jjv3rsawzs4/4gNFIafG9C0xWutGC2hrxhp
G2+bV6S4set2iKrmLFlRlC1gyOQ2E85jCyzvBrp2ybmnxqEupqExulqEfYf4OuXW
KyNmBOiXFMrShvjk+h5jwmjiJPl7/Gt+T1EBtY/3GmSiRbNSVlylor3AXYO56s3v
id2R07EwpuOJdHsfmisHIka/1v7eP8iSvSLkxnvaUarMuKFioB3F5iOlevSL/CtO
VHn/CJcpyzK5jSGtIElOI2HN1IJo0whUW8aGoNMGdzrQZnV95f9s8aNpmKn26/Wu
bbfoIHPBoKDeOwQ15DF5RPD4GcPACK4blaxwLGZ8jxoyHHsx7QavCqrwoqYOvCAe
oWxIfIfgi3FJHoF3wwtp8pCwPNAZptAaw6zC90e/FNVarpi2QqrK2AePjLURDN9l
3d1LeeukeX8yV2ChTOoujH5NwwzzoAu3PNHC7LVOWlyWB7WBHZNSngwlS9V4rqxI
XL+TKZkQ3pLioPnAesYvIRlK2YeRpLzuz4vw72M4LyoOv6r02CGuYj31xMZP1B3f
MGqDGlGCeAVh/o8xsuQjzK7oPepYoYoy4LG7b0Feml5nT5yZ3GgPAYpLB0yKhigU
JQAGlbTFzCZYNU+s61jRxuJo9NeaQ4nzeaM5mFHZk3d0K3p3lTgFjWCRL0vTHg9O
WFzhgVc89yQOhCsaRpRGoR7skk4XxcgOjXY8Md4u4wS0kaK/XbI6iwOG3PM4Hm7n
uUiZvy6mtyJUTC3BJQ/zZtj4dGi5aVzRAgVrjtG5myy7UXz7zSmRgbmVnyIwUZnA
7kbds4mprskTuaZBk9GrqJXEvfahL1qrRytBxYR4k76nYNjTSozLNHMsXaOZiGBw
3PtzI+qsrDzgCMGcGPqk2cOlZyDfhZmpRm9Iq8sL5R74okkvD/5ARVnCPsktWNzb
Kmsry/4hCjlhZJUmpS11wirhrx9KxY+qKfntrJMSJ5fWgGgeCOUEmmYmhkE+8Wdg
JFuwDZZp40oKt89DdI18jNIpr8NYGZCRecaHDNeA6eDEh9odmi03gO/2NfLd4Wrz
+oNyv+f86uTMMYD+dI9+1gEkfLXTuV7zUSss+bq4OSVUX/6TRUNalvc1aS4y8oaT
iwpf9fQ4xoeErr2pQRtlliLmQcFdy6EhquoaWWI5WBmWhcLiDw/FFq9m746HBUZ6
zwBaukJPq5Lsgk6YfGg6afFGPPN5eu7mPlp03VjAoj5Ql0oEHfsu26DS1+I/j/fP
yJvZM7nLpk3SgVmJKvuFhED3HhlARtVdZWpmC1jrflQyWfxDAScVEYdXivNx3ZZa
qbRvSRDA7V6icxA9R4yZgMUcGjm/ukhWJK4nB8QsQD9/1lUoWVR6+95MlZs/mwkS
u8SL60qcuKHRpvsJj9yt/5LHKb2Qtqsa8xUSAC6J+OAD+a/JSQ8fdha5ABCWnfRU
kgsvPz0N5mUVdn3dhrsmZZ8d5RVQI2n4bSiMXoxVRHRVDJBjBK12RqqmYTGWuTv4
5JJWYeH3PP1Z+T6348e5eTp2ln062yGTUbCcskSbItUQfk3C6ZwK+dy155RmeyPe
DeG121TpylWQvGyobf51oXNCyZzPMqRiUStnQHQXpoyCDi40mQpUo6Ib9ByV+wOk
Sel2hIxzmJiomE7tInx546oqPA4vC6sYDqcIe7x+xNGCUMPje1eMXf90rIbKRVpo
DtqfKYANzE+mmnLcwIvJPbrfiFuBZZyCFvi25miS9cExAJVSd6oGEe+8x2Fpxr2f
Pfaf7LSSEIXbXZ9riI6j/XrdR3D6EKhJSRGLYZhQUORAKwqh8rmP0dyNBKike5IK
k2kT8XjE0cYfuimdJqmQ69B3NHwQBusweJw6ePP81n5oGwGOOk92efdt94Dqvfnz
rmprlwyEkx7KkPWrTfAf2DAE2wWS+ONAQVOv+MXOL1mpgVdmiHUwCDtdZQ2mfeim
GE8zOURIjJPWoiGHKQmYblWhARjSEZRr8e1For4HerHQEDfXlSw3riBou0UidUyR
/JfKYJcuWjzc7Ub0K4yxQFXbv4/MKk3J/Gjhfh36B0WoDiYECH8mzD7rcMJh12EC
nwPlqv5aB1knYmTE6FlsomqRc3zlYpNvPKjQMvex8/Op+Wa4DHmxomuWZUklkaCG
r7XLol0nhx9dbgHpWerFxqpT/t0o72RBgf3MEJs9JFJnziIJG0EILxTN7XuZsv+v
8xlzRY2xXvPa7dsNZ1xAUA09jnJFBAQA7gyipiQjvj0Rh14w2jlctc0l2LJFpFOQ
Z916dSVAIMLlk47pjHfTWoGFcqkzZF4Ltp5qnyA76+21kJeLlm4l0fioDe112yEB
eB7Fw04H1IJF2ytXTqMf0VxUye0qb+2fUVDmTGfAjeLQZiL4A1S0hZwYe74dSzsR
vX96n98FeVn/3eWd4hsGQnauH96c0Lu7RTkN7E+w7I6D5AMnMqJZketjpfcLZObv
exVJR8fc188k5v/Wo1cIwvLe1b9cbRCWcUFhBunvOj/6Rbo6grA7crts1x7gU7M0
jZLaSwRMM5+kwOhbYk55/JjKsvEh3O+orF1v9sRtM4DGG0Jb3U/m+4PsH1+IIlAq
E8p5XBIWYrQXo3nnFtMxajcC3fAnkvTT7sOCqCM5x/oHiIog10uwOPaZDi4ZxA4E
6+J7mrM79pomwQVy3Y1xwi8jz6KrE24ADVzJ3Qw5nOeueHFBNyHMgg6GKfBPKa0g
DEqTy9q+EgbAhCnBziIQNKZqLjQW3GPO15sK00CubPn3586KUTAWR9XSNmESUKHp
pBbD1mUZd4RVXfek4hBIe5KbspKOfGE0XYTSUY6A+zSP0Gm8r1m8KdQTlW+QmSxD
Tt3xj/Qe/k4QvpooR8omqZ6P2baGmAl8o5rAvkGPkwXemnH0OsCksDn7cgdJgrzD
6eOTt/xHQbQW48SuKVZBtg3aJL4pMWyj3EnanZO0VTGG8wm4tfA9gkSJcIqTVebL
C7Rm8mgUuPcc8wiVGQ8iAFRs4FZ0iG7vxMA2jySmiZyhpQd+3bpgzKhNv+jCRLda
tCX/3GwmG3ODvXqKNAAKP5RhC9uF0B+eglva0uE+oqMha/Vvtk1VyLeG9UoSfTJV
/WTJ4J5dVRe1LWURSIHDpw3FMN7UV9qLYe/UScOedj1EweiQQIrWyM6s94Xf7qta
r6BFk0zM0MWwlDPs2UaHWH1KhjLmnFwwr7liG75JxqvVFmdIIwsbh4Ai5yTlmhNC
/Z+CdiSaq/RAJHjKL9gOdXAoHfsDN3PSkdhQ/9cXlJyYlIUE5JQgPOPzik+Xa2Mc
xdJlhkF6jn0/aoHRtJZT6uQeh8J/nF3VsSRlmDtNH5I7clJzlVxlRjT+qwgZZlz8
3YqOKIX6J4F13jynaO3N1xIMr0i4FUgkdsU9PAAe21meJj5lQtnFkaGYVOJ33E1u
NQmuxyQD2U0E/onJO4PrsGezBWx4th1bL014odl0aZfs+MHG/LJtl2L1Ut27eEfB
JY1/F8oynuIN2g3ZSnvDmtgqmwQSeCEJ1noLb+5UtEWRnZfXJDPhduUwNts57Xlq
wRFwQsxNp0emor7hS/THl3bIs5Zot6FoXNjVY6h5vnoUbimNHm4vOWt8Kjs9WQld
CjtHfokkNIs/IdpkFxMFgjEENKP2Xa3ajc8kHpAvJkxWcuPrtXD7CaOKFAiIpill
GVKgsscvgQCjwKkm2l3pUmsHgUIqTpxs1N5zVx3xz0RpCIQQP3Rqrmv0vqwRe/Nz
7QRcA+78sS+y2LmGwxixZR9WD8Bt6qylQZfHzXaPAJj95aY5Bn9axnn+ZU/5jgkf
wa/AoINIl8CyThx+4b6J5ksn3BXyLSvrtOY/pSf96iysCzdppbkNtXGQAX3NkrJA
+4hnmuANXnQ8hpGsVSR+5ez0WEnStZYIW+hjCK6CxGs82io8Ol3DPSGLsx5AsIJv
ny7ZwHovStW9afUJDP8XDL3kQugXxlEIX2wB9FViBFvOPZVZR7mIEJD3vxIjTs3h
a0Ayc0+W3yE+bf0BtKDvS54+9MZHEPk/R7X0qodNqRlnIuzUlInm03Ue9PQfSqGy
1FXgtv0QhWBeelLhcYYq++rxJmfMc7DcCzkEb4RAUXkf4pcGJZscwfChBcF8eKVk
2G3QR61RL57qGFUQFoM5S4uwp1wkbZC0GYW2ecpi1w0dr19kKLWIfhBuoGeTMoVQ
MBlHx2iEoS0h78TdgXpc0KHNZi+uhHnO3weZjjnHZxBKXPviYjHeSdv328LSWuhl
ASQ7LQdXxfjiQZwTHxDjo9fuwxda+M+VBoE1H1nJghAUff1MdElXHg1B/xu9esHf
A1gQqPkGcMt9g4T6cUU9u0Jk7G7a+/8hOcVl2pvtUt21PSO6syYkGrTAwirrFSry
06PgH2FctiCyKixx+uzWCRNK1/jE6sfhlWERDW9bNpmkya2oVnlxbt8UQEJ4HuRD
KwrjWvEYfAqPH0EGRTvzY+uV2DFp2aGyjKYgJ6esIvHQGqQMadUIRhG2f4uiYg0H
eco2EL6JZ3Z7K95ZzPcPE+IUVyaqflrX32Iuh/iYauAnABDsl5ufL6nSbP6R0EG1
v2sIAgbXvyLKLTv+FNdhK4agmFqn0xhnKfDc6DCnR4sIJJXLq1Hczd1FAXfVdzib
0FgCH4xKIVbzgmA8P1wVwlNCyfUlXLwntHzBcII86R4doFWfnvGek5l2kO5FENJD
LUBqlui9p7e2GOYCbH2PPtatOC9heHLKtB76ClijeEAQ9UFiSCXJGw+8kwrmrN3G
NUQjamvvEzlBl4JU/osOqeAsGjd0ylC6B7sulWCldXkpP49WeTmr897kZ4sY55S3
SEd18Me681ftuiW6JI4EmXE9k9HdG+CgZNHaz8BP44AP1A17YY2DRySZ4w5UmeQE
a4uXnzUzQvAeZd6i00daYZgXYxxGKtoi9Kealv6zWbFS+O3Fuch3VqhgdaGiYYuu
ymsU+9cxMjHv61a1F/4jPs5ihmAOD5M3152VJSttzNOALunTynKJ1gE33cuNQuc+
if472ySg10OoW3pFn1ulidXUXzEc6dEoGhFfNeaxb8ktLhl+3C7SipivBXnolnWh
p/38r/i4eM40TKYduXsvZZql3hcLlt450RaKOjWadd3deMNkgO7/jUkcoMPfhULq
v3lnPin2LV6UI+pHdpivQ41rHNJ/r4ds2X9+HOh9HLZ50BdE+u1/nn1pmA3GSzRJ
pevjkd77QBqL+cOin5HiJAJx2FUrJV/4W4/IA1YwsGDMLpRTswsKj/EWWRgdyx5K
1DsgPkCAknXdspfSB22OSmSZYzEc95+8Ydt5Ug6toLrR3DYKrPWdqJsYpX9sVh2Z
Wzz0U9vQGdHMwpYn/Ty3IF+Ok/0PP0y6IfeBhlwU7v7nDV3lp2mR9EvU5g/LtfVr
ulQxTmRLaeLHHa5eG7VDiLXqE1ryaGd19Pxhfue1XUU2XlFWYjA8I422bkD3YLwH
YvxXeiSdWhu8doiM9V1gyBlDRMVZgV7jUEKdSbUz7MhJkOjypOWzpw/msO2lfjGu
H5GoNEV5vLNAasQ81Mcb5kHwnJdZ5yRSXr0G2NvCPZA2XCQAO+M54dl/EYiNPlM+
jw/0UVuBwmWU13qLtVEhTcmomP9JokavCbN29GXpuzFc7VzE9wtEQ3EGT/AqXoQd
FND5fNUBiLryLxv9HtwGqNCU0xR0dzZpPt7lJ/EFXVKpluMb+qoXIZtXqQCn0HZf
J0V72LquPofqX5u9BOv3IKKPfHnoBYeHVL028vXN8vsKD1zY8R7rt0XFELzkJVYy
H8OdgMZOmqFlO10RwpHh/GF3aDhkzi7NNScc27XDHuZ89D0TuxX03yJLFEyN3g48
2JApVyT5na/dN82aVTMh5ukokJkU0N8o1hF3OECImZUO5CU7NCcq2c8RLjXXIofL
z/U5B5SEaQayvX4KBKoR7NkpW2Y6hrkqACA3MV8CjgnMsTMdXRo2C7GUzig77078
61fEtO8wrn2jT2+9/C66zdg88XvV3vtxTKavxTXjV9ayZ6g/Ev/E/p42L0Pj4s5n
oFbzvL8iKVCEgx20d/WEGk+LXPEIvBGTH6nF09nqppi0owf4zg1xClVmxFU89rB5
YViBE8Ed8yw9H7y/x1nrzq80nlm/cgYcNaK78SUAFK8TFM6b7zki3USkr92RDqqn
XJnOFoujFjB6FcnBefrwDfTpkCw9H2TdHA0O126IEK+goRk7X6Y7skZi2A/G2Cgs
M8dSiEZ3MjfwBst6gT1V3QsEzlrHYfmIrH5KMzUOy3kD2ZZguCCx4XlflMnmi+h7
YldZi1sno8KytTxhU8lnukDTxkvYfxczLgwsw4wtT9NCZeuzXjd2cER+qPSFBSoZ
duyqLDAQCxO+WKGHFvj5G926jz9ehjiRahPOfVaB5FrZM9oEHcOlbDMDD4h2shrI
145vzGAO3hHWeFxwBzJortXVEOzq3XpBL7goaUZCR0XbQ6prnCXHSrFs3sa/gXMI
GHUrUiOV8kLjwrckd2uOyOXfQJgsQ3yjSSrQcL6FSX0HgelWfmkUQrRUWQUIVXyK
4POBLsOe2n6DvvpJ3ngpgcBzGZZOybAmP1IDK4GDbp9oNE1XjnOmaxn9Zs62soD7
6bcZ9moub/gnyguUCetG7t8iiUZEnrX2VuG8O4Mr3REgTJESTe4Efbh7+sl1jKIt
45AIZzW1InsNBTTAHTfa74HEY2MFprKzV7ze5abokmGoQ0m8FhG3Pel3nFH8VeiT
KBVGNY3fMpMnP0IDU0ZWbG1+vLYqa9CEF24NN2YwFus4L9D/WG9pwVbUgr5x5nDN
VCZJqeI1UX+CJEAnLaQmWsuVgdDNSHTR2E8TyImc1lNGQbl5/sCBf/lzsTML/WLX
sWYwE2tmgXrMrkGi/HeEuz/MJ+ztR+vHID2n72EFEStCCmGQd8cVP1d1ifAx1u/B
ejFfS7iEcyfSYAarO9uwtXYZMAiJGAnCUCrY5Z8kdGS3oEW4rwGeD4K2nX/pb/Iz
Q/75+Q+XqMsLvS3XZiVJpnftXYwNqPzAZf1aIAQ5lpmOC6GdOKtoYmrkLTyeHaos
LqjNq72s1LwAYkm98c16Hbew7oNmB4/w3JK6M/sGiuS/+pViD90U0qfjXz9LJLU2
5Di48FxRzJ/hzRxxsRDuHqoHphF+gaiyS5strHeaDTQxLDSDPoHR+tbLfUP1EIna
tfGny6tv2Zuwb10lCXK9h/13aSERarxiIY9YBzxXdq6Ivf6xJ5RoHbY6vTa8838+
4YqMVVpZ+qgIFIzomI29Tb0Pi1JgTux8l6vB2THGhKv5o8xc3jbyMMo9+PX2Yja1
UFgGln5TDIWloadhO+TsA61XOrV5jLq7G70sa0ejs+rmQjhxrau7cz8OifHyPeDg
Ro75ZD+R9wxDgrok4HT5I7KCdu4KNWfxyTr4XiWCv0gPQ65L7gJ6B634lxWWDcxo
kSTpL0KSgddXC1DqDkmUA4U9AbXUblHmZuiFqMCZIoKo8/vXoxmSWq3jUvg/UDXW
+WgCyS8umPOqAPezDYjpzn8UczN5C4TdoZ+/+2OfSZBDBL0TJeO/Z98MNqKR8pxJ
CQxC9vfDuJkXfNMvs6+33rqlptl33Q5eqLuCLBqtaV1unhD7nkIoKUy0BvpNhUvb
nPMG8OFa2n7P+DThwHbbXrwHbrwABvKS2l0C3XzUOVbZA9TnkiB838b5/G2/gMXC
BVB50ykIX92PI7cfsE9x04h6zx/RY9fFDwwkoRJK4jigJy9q9YfPkguy3BbGm4EC
PkdirDml0LQ4KrUv4I0w7K3EWCDVBQx8kHqKPmZPfJ5IcBUlut9jdFJVy2nuM+5u
S1lvnzjM4p2hZ4vngIJb4UqiK77VFFs4iWo2dd0MOHHuYc4Kq3aWt66L3yoFp5y9
91lUyRvXd+bTNngj5ojAUx988CBiYRhMddEPmEZi65qMvWkS35WseVYKjXB5yJAu
Zw8P/n9lHdSLgDPopAPZyT2kKQgdbMTrxnst2pRPn8Oa9Fmm9/+STkF1cxxZbIXq
X/SQ5cHZSQu0oyrgZd0t90hVpHV474L1Za7Nb8xMPV2vSy1de8fOgdgK0Yr6MGen
Pbc4B7XgD/jQ19esqySdp3tpK9SSCDAVxtQr5GIvwLDf3fIPfOEkj5cXEVIMNc2r
kL3sFnGeGQbIsh7CQjiYYC2pq5XSETmVAYhnZG1NGunqxG63+vT+nBCm/p7AUa8h
y+7h7sB0Sz/ZiSOcvNj36s8upf+LNfWL+3nBHn5ZKPiAlmhhzRN0xNY5X3Ojmlhv
QZMszFdwAQobaQqVMTzu/kBq4sBe652A50NGm75WOBxzn+6J14PLRaTiy5lDgv2U
vVepIEh692L4vub1SNpxf01LlwZjU6MIlaPAczYmpw+mKtBfcN/+NzJbbcyUokZ8
Cyr3Wu/w8+Wpq0XK9PUqQRa0EkUGzBs0ornrBE+CLikxiBnRRJRxwSg1x0KXFwf8
u66MWYvHwIdPAOhytdXluf3oxRoYsEZOYJfJo5fG/iZuuiOQkGgKT9RlSXOqB8jj
xQ0ntUWZNcBZsaIR1PK+lS0RBqAELgcciPkiISbizMc9nWcSLNJioitMi4oY3Wtw
TlQHNphQ2AefQl314EuQmfoFuS86cJ3XL6c9nzqFh5ja2YnVVAmLsY1tDgQslKTF
+mqv9pmJtOjPcxdktXlC7ZcYyTS3jgwsKK2B5+U7iTdl15x1zpc8kf7tZrrzFAYO
MOUd7aE/TXs3G9LPGiWJmZC7O9ERTBnw8dArS63GOJJY9MtyLFHRdaCHskGd+z5k
ZHtBrMeHxS9GE9xrZU9bR5bLkhUZOArbTgUje64jZHCjic6gzDkwUYcCG8KOEd+P
FBCrDGeo/KuLIl5sCucvbkAGzqSuJRosM5wsntXXlMIdjrfSXTy2GYWob3TaJFnv
ZGblL1gtugJyP28a6rz3/QJy6rks97r548+AYtgEtUgmhpe0IDKTwT8CJP/VPRzn
NDMSdlr08YdBt6i9OPAdHK6QyFvBXg3eOl8kurqrsb0GNwJD6sljNzx1gfTGjJbO
sv7fWs9oH2YUUmhk8gspH59WIpyAd2J5SDMHPn2RsyBOIL2vO7o+D7V1InQYnjT4
49+EM/MKeDwzCrp1grWwscEKdPx+rbzdW+MGp6PcwuKCDHP7hIu0CNH+0YNQLIPq
c9jQVezDfrGaJGKA08f5vUkpBFOOKt+rauywj3+coc4RQmIR+le5mW6xz9WOORlR
1PLQsGu977P19AiYbQMnejdfUlTPwlN776HmRhm4PLAnIB1cePoqkwDXNMgMAIjB
pJos14rwnVzRRMBufsF71pmwbx0XEWB4nx2NkJCfJtIYRl7WPLneD+3O75NLKobG
wgaDFUCEcnVNq8MX24TCDDYByVi9LZAEvX3lOAUWEWpJWGa5DiZhL7QzV9OlLMG7
R58La89rGNhxDEvt/57a28KxMzIvoXcMKMnCBUGyqu0E3f5gkDgtydQJEyEWNfrd
/ChArfXmuwivtNFs3xO2c4fwXlu6v5hzFsCcZ013S8g1BOeFC2OfFJbjS3ALJVex
rgsVaIY2pPtS49ucyRt6rLT89jmkcQSSjWo6UGO00M/NQXcni8Emq8epL0O4eurn
P48h9QWy9VRbd/nD1TzT685IUXdzQx4+zOQaTAaIU3hgGYyj+jcdU7PbTEMFKWy8
75v7Mky7fR8BEl0KXeAGEkHU1CwSN0oZ1r9HjRQtO57ygEC466//aoWB8PdisCaX
n53gjrhkN7HapMhTGN/TxkIrgaLU/L+qLaaLyRB5Q+Mh2IiIbSr/Ri3tNDlE3CD4
NQuueqv+VjPJ+0DwW64upEsKvrjCMODc9hpxiWanj8AW3hxejamzkkuKZmJLn+Io
LJr/7SMsfQvESRvI4FMxUdctifwwUERZwqEmKMjUBRJWALcQNbYSiXEgU6sS4/9N
Vm7nA0tP1IS6ZT3usqzBHPm1juSNztNBAayErrBbKaj5JJ5LLybaDA1c26AAYkLA
arN+Q4sO7rBg0iGGbgmUyK3Lq3aQ5cwPjWewZATuR2+nq6++Ltbo2rPnpDk20dNn
kXGEj45oWrbqz2FOA1WEcsZcAHTbtOJCDZgbmUOsOMLROU/Csa5XhdGCBs8Jlvrj
owvO3Wr9aVTF5njvlPf9MLoIugf5fL7iafYaw6v9d7bjU9rfgtMpk1gER7DICIpF
WsFbC8nJsEpGVIqw++tH91f1QvrT5B+/3up+eCUfd6kwUqF6egRfe54OdJCpq51u
ocibpqrHPIU9g7+S8w6Yh1fpx2nfIuqd0ZwvhreZnkNeHWSxQpOab/8Al5NcYVxI
pTAkjKkcfu4MLeirPCXXhydGDoVskHOY/wTt8y/CZ9KhvNutavQKbvioX8fleo51
lx6lLerYAjPMbvP2ya14jlpNy6xSDcG2fuS5+ezesf+13ID8OVU2fMXSgbkaB8x0
CRap0GvJ1mtiW3w7o47LhzIAImfLyZ+t2YuFP+PYii0XA8qzV5cvonYzfTNwkmtk
jygNAtzZFvVxd/yF2SqxD2lylYYK4A92ZfoXj7sdqmj/23A72OLvdgFnlsZl8thd
qeG/kBId39fiZLKdSN7SNXbti//jcid4zwgSkh1XV0mzy65ax77pothArboUVNMI
NKevUpR77MkPuRrb/8Ymmouz8rZsoPyaUzRoTxeDoJkfE9oUD+up3BUVo9Y3c5i4
kTnci1WEVOoqYG3S8mSI0PWknU1cjRapg5AZpfdoiY+M84st8XFa/a68eMEidb2b
bP+rmEuWszlq/BWTSkQnRxBOljpnq4ctLLd7UVp05GF3jIu9w1nIHx7gmEl/Yy9m
Jb1Z0kWEVhGUhyzWQwqNeIYzzIhYzrVCLIIaT8z/EQ2JUal1/DodRqeBUZ0aBig0
uyq97E6FNGoJSdByCjVja4XQfyA2NhkW9KQMLQ7LGo5Hu46xnvF4ri/3atw3xElL
eHOdfbjtY3xrvvvng5lxyycqtQR9KinwwRb/XcMV6JHKfSxqd+1juOyz9BfhnaXO
q/IjYtxpdHBtQvCU6upea0NGerBN4Ri3HL7VizQmgSvbFK+ibD9b3wIouEXFc/HG
/AHZJr9XFpqdt3+sbcqTq71T6EDMJwebD1o6/kHtYjK5V8uVHtPCt5fTX67pqInY
bmxPvTN2BoqzCLJYXmfCJR9d8eJ6QtVwM8YyuUUbbU1AE9mS8WIprdBUF77Zwo3C
1aPbzHecBMrwpGdRFGOks+Ngb22JBo9+KjB9Y/KIAFgXHxnnESluVtyWn+lw6qc1
A86/gk4kojBhJGQ5A+LwFxTIFTR3dI8hp8iTGTlDzq071W30n3UpkfsSJ5+nWG09
ZpQB35rCUEhA+HnFjSKZzIpBzALJINQGgc+wR+rjMWRhTWMDZAlxogQrMJ4HtIw6
BYkl+8y6GEYYdhwtde20bp/bCayMFY8d2p+tayKUIdnSpOaS0nWsqmMDkbVi8XBp
o3xPco4d54hFBZ1Gy3FYCg4lyBT+arxegIG4R7NBbiqD3ZHkTxcH0dm6fgfAD7c6
7se/7bGNUJosimrrcLrZDkCZyRkks/49najMCPYV5S8ozOv3J1/h5GEQy9WK04U3
KHtJ2IPfO/yYf8FvuL12S9m8eZl3YQbdwYGqfe4yhmbNnMULKS3n5HAZ4NieiJmM
2O4sZOy3hMDewOrhGTTMaouSjXon/saVIW2GamBJgLkQiu7Hn5G3mkUeJmu9bv6g
UOr9ys1lmRzUMUAe9pYP21zNqn7gfOJkXH1UpmSazX/w2Bgawv/chkx/CB5WQoUy
ciOXAo5/IDgkRNHmAicbd19JNSLqfJO9LYcGvY4rfZN8x4+3w7RbZ/XY59onqGbI
eyQv0yEo1HuLUGiS5SgqPbkGCP9t7DIla6gX888uApvD7nuPGb9JhUiDiPHGRzU+
THntDTp5WlnWK49AS/J4X/f7T05nqE0O+upQVpG/ymJNhUU1sWeehjJNBlfAafjX
dH4f29c4C4DSCQl56HUtsvzd6TTUhjOVpseUJO6CUDPihoZ/t3CI6Ho/ZW09GR8c
d+j32Gdg3YMLk8SRGmnVFiHu89/ZVeTo3SVR+8o3x8dpKqlbinW3w1iiwLsq5iu9
2oRG8jbo2GBfXJ6YJN+Qg0endfFIPksn0hf8lD7NJkZvG39sJgnQCr3O/SuTW96d
l8+VF+Fz6WfMk3fz1qJu6844NYMsnPt3wfm6Q/AToeqLpLgWUUL3KOZ9ANoq7cmt
mteE3rFRzq83A6hKSr+2ymvQQsiGMsftMGc9XweEG1GMZ0dJq2sWfwvZmKQ1018a
5O0w2uPqyjuDPAUp7v/+LsI6yG+SINJj5iGtzD6yJ/2Y0MLGdk5dCr3IIgCDSXzY
Dac6wQugJXyueNRIjAVm/hmsihFBDk3d82f129hhwq7mSfEqDHIlqv/tDVGMygYW
/RIu3bof0XPrS8CbN22K9urGaEIqlqHr6IgcoY/6Gr5UKczQpQYFt7Arzm9GWOVO
KlWnrWjZeByMPCRBstKuaMfhFFbPMm9tFkYail2Dl1a59+ujIKX7GK8sPu8xWciA
wWuULbIIZKOsRpazaRuXwpZm7F7IuClTaiMpARsN4dnjT3Cq2GR1wdrEmUayzssV
6fF6dXx4Cijd34mYj5g4R5NiKmmlmd32tLPZ8oFTdfN9ArVSwncKLokb8Z3S7Pxq
dhsXS5Fgo1irvXfOsz7u5c/J0H/q1ink9gjmNYgc8zDj34BsFmZQJGrqspcd+9PM
BxX8cu4HveNQQ/C5w1j95pbqhtROhsl3aXhUtmM3vXMpDzPHliYmKuJCa8olaHYJ
2h+nGRjGbWvXyjecL/bAYrCWKqrIh8eZV105fUHDOa+Gh7edrOMVvOmBH4toJjNb
t/Ng8RcxSdRC+5/0UJvdweeBJs0h7IP0uhgj5/EDQyZ1fkvSOwC44O0S1LteAsyM
4Xeiut84Ql3lNXKnpJRsIwbHvopXuCUPon1Jsx40SavpgVg0Mcx1F0+fwRHMVsiF
3uKns0v2tmvmTKyvq8MSXNMahuFLD9ibcRIH58UpqG36BD5+O5RsukwXVu6cIDzO
4kIGjMml3uC7xRsmtOLPRNbLYEjsuWbp3jVH+YGKcCa60qgOKIKeUnGE43ulr12d
5DDJxrZQVjVYRhIYzMBrbTlgp0GeTepPTU3V2CpiIjPfw3gQl4oWV/b4KLEGAkN+
x0sZpRCeZs1JwgDwosnWXmgFeFJF3qNoMcE//heBEcYznkZSrgh0DQm0ZzjlDkj/
VpmM19M1Rm//a7+9/tj+SZkhkjq4bMm5J+dwXHwezVWnRxvV9NMx+edgzGeFHGGa
l7d2pi3+/U7ik6sr4z+2wG9Pt9FpTWZ1T7ZC+ED8LYb8wOAYnEJcr/FrX8WGubr5
uzInXeD2xdyKC1/im7wa7lT6FH3SBMKO9lK0cwmsOe/ttAAl6tHBs+Hr2cI9m85H
xkwEdSgwi85Qx/U9gAlflbgP12bU/F37PtJO6QeAhgugOPlxC6TyZmhSN4dRdczW
eGQ0SsLApUUpecuchc9OoYhPPstPRX27nt/8c6okwgaryjGlBMdSA+lOvaMaODV0
zWaB8Q+U//IkoOh/tsvjCtBUxpKLJkL2yfL0vgfASkBkqyHCNFGdvjANE2zrlw4w
AwScxQe49fKhmtR6lCXgpqjQfwDpfUyWNuTcrSj9D5L7q2cnLUf6ibUCFHaxXJi1
6D2po4/357B2R+1Dg/DFBeyeejScToJRfdMQ1K85KnnIwd68dztLtBHLIyhnf/Jl
sZyB73E6dYw907FhJoHD+O2BBSAr2aTT2c8OyVJqVBIyGL4zcIu4LAf3tUWGwsSa
3FD36y2Ht8ok2hyb0lQpduzMXSuTzvig2n44H/BC+/T3nRrKogyYeb0x3nc3pz4N
fAnbvAtCaQHznrMGNTO4H1GYz1MPLMhlMJeOnsd3+g0JLjtzz0FSQ13ErFDyWln3
IURhkuWBYerf32OuxnS2TOU6wtU7W3mSogM4sMB00j/zKh4ZcncTRU0SMeCniRXZ
HqUHWJSwlyICCeydncGlkgsFczeTJ7NiFVCR11kkFk2fZifhuHUFhLx6wnkD31hJ
FYtGSFYfKW9ZCNBFNSAcY2eZtBA9KCDdGzh9NB9jUtxNa/+LAZCsmOErqA7qKW3h
wtljtyEkntmnHJS2NHe3Jkbv5tR3+W8qofGAAQpY72i4jyF5IkddgzNWidCLRPvu
v73qMj6no+/V585/4ECk0zD3cuUXF2r6ca6y8JxKd4IySF/XJm5r7zKCAh9aPMju
ROj/Gf1eFS3diByNlRXBICaiMoybKTCdvIReXTDmZlX7E9NJCb7zjZ+zh91J6Cg6
1fahXgzsekJo0EDyGNPZh+7mphGPTbv+CNw0ISGneFWExetCogQzP+TGtZ6v0M6F
jaFWAmyAQLYtmnSTO6GrfZR4lGq2UCOQfvD56hOSexCty6NhINDPZdpg+b0jbP0o
ajeGX5UHMijpY7AZkt1c7zS5TaVtElMjtWuJSVSe0G07WSa5h5TuHEonCIk8wJQt
QGh6ZmqjsAVWyFY8gs85FtrkWW3s1dIz53eq2efTceZIE1gON0U6s/SXIVHa/nGi
Mp1lgub7ZFsIcHluh5HcM9uzMaBEZHlJsIS2kcNYAIQGHCDZwTWpj4rUwGqwcZA5
kNNnnnOprVfRRmqhBdOCc0GdRtRYFB32K8x4UOsB5O7emrQct2kQ+Vgh9SOO8IdV
AB2hA8Y+bXZ6ZzhF/FFjZTkgQA2prjT1C/qQRfSwMMSeU2yW4HbrNOdQG4XkEA51
9cY8PX5qJxGfJeVo11R7JQ0cURytq7UG4jluJLPgn3J5Z9l3UV9F6C6YWKSaOWza
iXBh05HMrDCIgKPg8BbRPoekI+UO86M/Es0hMbXxl7zuXbCnyAZ4dvecV7WJXIB9
ZooIWRjCjVYURUt43U7xWHbPiXfOLilGzv2Tp0oLaumIPsXuC5wF8k6WaqET2TUz
hVTwv1Nk4MShA3zBKjAo+SBcGI723N6P3MQa4jy287M+NJ572SYJa4wy8OROE9g8
cO1ne7uo3FW83PEYw5MFtL7dZzl9X5kwF9X/OOs1f8nuC4AmRKBdwAq6IV0diEdu
/TmBktLj/KEobRV3kAi6046q8lL7DYa/qtK455jBMyxZREOFEHNW3vLwF5R4dhd6
vAt4EIFkWj49pHC0CF+odt/gsxQmkb30xEvvSobpKKz2NZ2ZtXwnRi8aisRiJzhf
Xcbndalx37Gt1XTCgLiQEy0crJXk9SRwHI4iGS2Ws4ioclv6ONpecJLOHvZMIQd1
PR2zoaV/SUQMOqXlGLw2KpxALi9DG0eH3I8JL3Mi0qlKIK5Ny+0waKtfFmXlg9As
XQaas3ec7XrWm/2rFb4yexItYEQnYtGV2pzXUL9UJNiSQwm+m65Cp0v7XzGREsai
ZxKnnMlETs9wSRfr/ZOhADZcHolzjQ2aP1nj3A4q+BHp9UYBa0mZ2T9y/i8Rvgsk
3Hm1FofEkd10AlsM5HJzRvPqTrs9tZhZ3Jxz/SXKOUEecEKlpRNCdM6Zo4uQFqTF
mgWL2AVSXSwWxKGh8vJJbBP4vfPmhIEwCUReHh7UR3KmBxFiyaOd/iOjeP0TC76f
MDPJZb7J9ezCUFDMuhsqLjEa5TuRnT7Zv+Fn7h/cs1eefe6SWwz84emWL2Fb1Yrt
GPCKPqTzxV1190jq3w0XS3ssSZjjiej84K2Va8gekjM8uhkxLsw9TsAdun7b9iwr
q1t2rKmYz5otYZ441ukFadHN/5hj4t8LSZQJVWl9oTs8noQiY15ku7UHG1vTlFDf
KfCxHJytUmpeE7RB6XmSEBY17M+NHaZz7b6ivgBZPX/SFlcuKyfKPp3TwqcX1LTH
QFP7g7bkHpfb2YdKChKz7v2M8i/V2ttwbqshqBUEloUnDaiqyk5JInQ5L8NgNQEe
tqbMVlSj+Of9YS+vRq2LijCalC2cQVLQFQhiB+y+XBGayrFdJDJYcNRdJchi4Q6u
NkFgrmRJSG3ij3ey2d7IWXfH6zp2eY8XKhC5I5G8N8L1fal0mpa253aMwyIxyqcJ
K1KANa3oSwOWrcq0DF0Evn6wbhdsXsiIPRFjhYWQsOAMEnCVHdGWjBq/p39wIzGC
EWaKDR81YYVMeIwzWc9P7/y76QVyGueX9ElVApO6MmBtdcE2EUFk8Qh8/WaRMNfw
9AJS39x020hjzBzYkD6din8l0VOXlVU+4HvWXI1wPBp+42h7aAweFqOacdzZx0IJ
yACsZgCtgszpkflrlAs4e0+SOO6ggGCCisBGz1Wyd+wn6hWn2GeQbciQ9qxYYunT
F6cHWQqa58ehi25QcxnEH1I1m/Hwn2fHdQsWAsHXkpJ7Nr5/HSdERDof9KHDpEuh
Ekw5TeoimWhGQSX9LS53DaG0VTfv4+VzvU0feMS9eNwLomDzn6dwHcL+VfqFjHqX
oeZnRFSUY9Q9N7GDEhXDGPcuqWpKYZEAbGR6UZDqi2D9114aeeefe2YH4zdTkBDh
VHonJvHZ7RTLjk1MM13Yj2cAYOVCuWFSRYq6zMZfwakx2jgM/jzBnSCG+ZT9ilUH
X6i9PKMYSQej85KkfdXKbB0/QGl5Roro+aAQKpDCjK06DJckFwZextflEu85lt3K
8Tu5UnwGTHCb/Snb35IKeDmAM18djs88EjTm5OQz50hMV1ErLHey7W++OlNbCPVl
lrqL0LU985FiDltLZt/IitMlefauM4t3ZmCyGz+CPyg/rz9Dymfk/zXtl5IbScsp
H9fsimvIbjhObjsc2AquqykiyVGLs+HvFIRGqMT+h4TN/LU59TXTUD8vz0kmKS1T
iomPK1g0UNl9TaG4ScJHvtzkU5PLrf3kjaN7GgcEZGsolUi7zwW8a0J6DXTFDYOZ
U9sbYmxOkV6rMtlIpfJyUtxNSuvVbFSocKhZh/2mcJ0q52o5Z+9WnbWkS72SWm/2
4Y4MmWAhNtX55E7FPN/W7SeK3oDb2jXxEkn8seNrsFTeO9Z+DZY7r4PPQ7p6foY2
0Kn9HiVHYtHpjnrEo9E6PTOyokdEV2e/TNI6HJB5CZy6uC9gYq8msb8VckUOe9Ur
BMN1/UwQiREoBx8t0a8ZVdhpgmXy3KTyzyFUfbwh9ueM6FwN+zzkDCTvnGsHlcRf
gbpBICSv3fDQLanBPCcBFZrJNoSNmoc6ZjA9QFvoT4otA92koy8Okw+2WEIui8z3
I9Kk9rpQQlYwD6IFAD3cObyJ5erO5p6UmckgMcxtFtG8GTmZL1DoqtxrmwOcC70S
APKVyNZ2uo323oDsbSZ86jBL0RSsvQpq4rUk9OFv53Y9XlYZE2rgAPu9FFgSWAI6
fWFdgHkYVQGIjwprAhbj3dSHCixbxRVSveOARYVmNCiLqqBDgW2i146fhTUHVbIE
EJwdGLNtKKnHjhp9gABK3OvRNZn7WzP9hvC1xFLmXxX3K6Y/hmt8tYGDlEDbgDJg
yLPqIUDdeD0VluQ3L7wTIOjBySR8+t7NxK8y4w1hk8fPkGjQAdeCT7V/gu3ET8L1
P+Vn+bKcLY7tWeOmbYgqJirs9W7vmKj7OwCvT/4Pc24hYKDaSHrP3NDTdn71aH6g
bn+APmJhxrgzpLLD2a67N8FLDsr2ownWsyQkp8llzwkOU+5FLGiUZfxS7/FPIOuB
woGe4s38ybTPZJd5tlZQWIULkIJtmVdk0TqQwaYzWl0GGOjTiqQQYyiT+ZBhJev3
/PSGJ5iIR+CrXhnfoWfa2GrCB2vAfYcpfw7Xh3V+2LEuZQBrcEhC9GIeW5/6AVcX
o3DFyGWVElkVqKyiOgTsg0VTAnUaJC+gF7LHG7ZJYGuL83iemzVdofvZKRKk8Vy+
RPh5NPiNHcKi+isJKnvgPMWMiuDmMtX025lEjBcQi+UocWKyyvVJB1SMP0E4DCFY
mJoHBcW/p3qWLkG1bhA0C197fe8ZS+izC4Osh6Zr5drqYEZxb3O8qFkB5HQZKluX
jm5C4B0gPaMnB0nS4hEvWyc7xNi81OreqesE85RSe2wOsRbX1wcDpZi1P5uWVq9O
KUEhIFAHHXi4OyO9E9UP8CZJ7KLJtAnzKjB9zqQ2vcTOkbpkBqASWT0f3H+1yIBs
pHhAN5k2QjshHukZlmU1tNK8TM58fXuwR5MQ45Fb46GA1g4A0fpx0fFJwngGjOX4
gnhIw6Ek18j5X3rete7cduTW5w52Q2SkmBiMcKKZFg1P2aiR58YqUNGEvLs22vtv
xAq0sbalD70pgbhY5lymLCTs3dB/FcsYbq+7CQwQhwT61d4uOhLrEashzmPaCJL4
MKhybcPmUzuRaHKVTKqjKfE4lI0Kuz5jMZszV62uPYTg9hMsn51ZzqBZWq6pQ5oU
nNE7buJVgOAjoz7Cv8Wve6nfD/bZ6+Uvc2ihP2HzmwaEVcECeivI9mYGmlGt4pYN
DT1ORXr3a12BuMXO0xZ+/AJeJPhVLKP8urLNAqJBabvCNapM4dn/chl4/2qLlhpL
B54e/xHfbrJPwTy4GPIlu9JQcizoxMTAL932ICR5XpJIQLjicQoQ3iN2vj1O6LyV
2o9Oz90db7V22f7FnyxXiesrmLZX0ZPsNNKxqijHCm+7Q4dZB6po76UiPDh+Uvtc
0uaO1LEiU0b+s/eD6mMxMjD/EzW+XF8f1xJOy3uAhJZk1U4+gWT2gMF8tiyuWhcu
ea5xsRflpZ8Hg97aMlX4c77FxhiZYO5Gl0zJS+Sly/14lxhy5VKI5r18LevCpzQf
GnGWwYFt434cKqc2tXn/vC5kR54DO4812qAlEQzB+IpHXmKPN4MaKfMyitpgazbI
vDNe6bumrEuPvoGLCb3/5bX5HD2WcZQLobTuAo7YS+PsNAWsbuBdeqjGJmRlrJ2Y
cUMw5mTG8qKoKX+JAX9Kr7qMwQsJ6Ahz2HPVDhLET4ECRXiyR93UNSveFLh+HLor
0I7ps1u1/qNYzgnc7oqAnvxzP4c6VaW0Wf/ZTDLTAKORmF1G8X4jqnNk4Pv5VbUr
pSBeFTZ7DyLyE1y6eley66bkSyhUjvRXiaerPQgx6bRZUFLR9lecPZp8gcmwB5K1
16z11ZEboftl9YdodP3oeV3V7y5VxD/DqDABHYdb/KxigKw8GeWPi+2rpBHK8nC5
3AxJUs9Xg5MeYHaCKR/Aq2jCFP2aP7UD+goZOzInptYjn3GBrRczMa5cYWfF4fPe
nUp+jR83ipinCzPSAR9WVkE/ZgAnswHHKyr4u3xTxWapFYt5gPERlnckRl1GXQpQ
CbNlC//51FR/dQf5y8MgybR/vOLKIJG/g41K/uijnd0JxDX57GbD+0cNgQBPZPS4
DkxEYE2OLxLPCE8Tvy5qr8I6I1cYXItPlgYwm7eh2h9yqsz0pPuFlsYv+CYhQ7uF
fcSp4ZDBf9h8ZaQnHORr8n6Jr/uNulEkTpbRsTcP+miSKNa4s71uqGgJaOnWEYhz
bnSzX82DQyn+yWmejgkSUC/IljXpWS4mG4GiraQXGhQocl/W44GcWJZIB6zUblO4
1Hk6LryGvqZ6jpOepAhbp3nLm2W2ogA9MT+QQN/JynSotKvS36QIdR+31oUDEWMk
1AL0mrZaRa6Ci8SnXCcLLYBa64ZUJljjIYh53cxAKAGrExhG5NCuAHJQA9IdWLNB
qGIY/MMF0ON4Glqu++eimzqaBIRmMixk30OJIog1h30Gh6JYhI0AYwjyX235p03V
ONQG1MZ7ibMXFJSdEN6SlYgB7kA63FVsTNgW6Abccg0JSE7tIsiR8q4i0LIQqo+B
2UhCR+x2DzJ2Uw3iNqUA04FF4PYRBjRREM2nFuNQXPPl+bNmRj53+A0deq8v2Nah
dfciM9AAyLLGxks66eojEFz85sbU9slMikSY2woHUtBR9sNFGio6PN/9ZMlLL5wz
IeJwiKyFn12DYy8Udu6pMVsBt4bD+eRmoZNDjiCAMtrkLoB7OYOvR0Jl+m0Q6k31
XIr7GSBsZOwJlFuN9LmO/00vDkGQI3efL/7Hfh/+a9mdAkAq+1QvEv49RkxhSPUQ
FDPAu7tz2tfEOBKU067+CNFsFDYAelZHFyv5I1llhv5vboPxgfe8AgimPhcGZrCP
TO81rwfiTHFI3IiLLfP1postvXObb6W3RFAga19mZ8XVJt0+TwSp3dXYUopO6cUe
N5TW1PSLzm0CiBIfYh4rPV2CapvhKQRxoPYnNfzaWsWux40i2PGKGxA2V/rJbtdG
NTs8l9HECR5t5lQl+wqjPvb225m1Kqglg1aISt4xeZVDuvQFrYPToXwczWbekMf1
2yaStjU+kJDeQNrrqGfgOeqP9Z/+CLho/I7FAoPzDUzxHdFPCSZdo0b0nau1wrmu
9MgrYcCTXIEdLHaDVLsqtTRHzHe7pPaiVboAPqB5T4hSqxQYe1/hfza7NJiGWreF
6C9hDSvixYkdVGb40h1vUnvI4HqCPI58kLrMDjG72NWbeVajh1bSHG7+Bpu6hcFI
kq4+n0CJcRqYZ3HAjrT2pJuzH6+o+wGB5b8MYIBMtYWUoNvGfE093PwRCBnvlCKt
iZ2cZTPFCwfQokn89o40u8Fxp3hfy0PxAsJ0+CrvGMqWoWCmTlTVtLcHdp2Djl/9
sjYNZAfVMaS9hS1ezqfnWaDRtpW3x9HzrPG1hQZWgIUZ3Gvspy3DBVrWgfHDI41/
8v4efJQqSVSO0o8lmMKeM1z+GCcW0S81LI7zonR8Si1W8sPycAg0UJacI02Ll/zE
f+0/D3C38J0nny6yDN5v4gjUeRK0gE+1+FZo5njojabvdGOMA3PUFVdNJ5whuIuc
7A1edk5IJcaxqvh9uJrpml0KUM50pGFsJS4UGO5Uew3E982Y6G+jlGosDavbCf0n
N1kAdzS8HrCnMEWqjac2rqCQ0jfva8SnYUs8aVtYXRZz3j3gCsYpyCD0FrZLBg2W
tjjMCUjFNEKQ8OVUntJ1QC0R49PIGaVtCxMjJUSJn2nvtrXfLnWFAqSi9wM63uIo
kagSH2ZeMH/CbRav3WMiWR+yG7Xba+Xx035vzGpCXAN4yqCVb3Lrv4CZQLc0/88t
6VxC4V0dyd9kKEtbx2hKd8DGr/g5gMAwA1g1Rgj0wmYxRHgHCKEAtCr7gQxSuy36
ppY7yWDzfEpaCiiob8/kzvS+HuduZaA5TsZDlC0zXugIXbXVATVEPfIFTCC7sGX8
nzEcp7i2NFO0La7A2hdJc/6yi/W8HalVP8AaUyjaFis+19eq3N2H/DuSO5Polp2U
F+pTJbFgLE4iGEY3yNWGv890xhkrn9mVP5MKCGT1F8iXsLtRF6Xn+HOFDNzTXPQU
mvvKRgJo+YcdOmQvyJQCeQXccHjUN/apDsWpiD+4HVkK6Y1CBYptSjwuNOJn6Rhy
6jOCwzfpSpXG0QcHwVpt0Hf5+RoYYdFIv1KD2P5NB5ooBvuNfzJhb9n4p8k/LAEV
mPEwfIVMYfqIF1d7Wi3q1QPDPs/la326EstHbMp93fJ+qRFPJQoyWWQsE8twzE6y
7Jdjg3pQFbiDh8WySRoWOX7x/BiZKHGTpgI0hezB1e0dAEM4OpCJdmxFzIoNNnDs
Ay/1v9uPcvAFbpvN41ZQw/A5LuaIfKUr5VIuZXyR40VKV8JtlDTt2PTBRhb51yon
BmhhGwnwUje6fjfYV/pCdLsv3NtOWdmraoATIYzMT3dW8/KQ/QfdacCp1j/HwKLE
zSK5J+Vl6WqUTtEy6lCIXNjvw7jkzIMkcprEFk2p4Q1F/46BjEARKaKlhynqXW0T
1KDZvbHIrjYQynglwVZdZknyvgUyATOvTMh2mVlczhF5yC+/M4KIjFegz+tTiyaO
8L61y3P9qkMNBMxaqk+F+HONlG3qEASw4hKcEQgQ+rjUCDZLa+jOZ3fPeb+kWMfy
gSlAzTaVFhCF372nCl6LhQUdz2m5wVNAhPWTSzN2gozECrsFnfyMGEDQDLNUM1y2
uAAfwGlCtg7NC9JRH1yaMyoWj+AlLXnz+l1I61hNqOCD9cGprfLKrgsVOfH9LxQS
t8tHhJiliKCb4klTQd9oSHXI4G3804dnCqQSwgJjHhMQkhJ62OHQPHtF6UdHpYMy
iMqFiTcDzhExKhQND/wLgSaRRB8ASq0Qj6zQMUJ8pBvIE/NV5iBu+Ld6yevyHBuV
Jnsg/FfMY6UDKS6Susdast2FEan75TBUwca2lNC9oF2klr8+3pHi3q2v1NjlicKq
nEQOhwl8HMwDdAhqwn2ta5sgprGn4lAvwNIMp9AkhHjNm6rv33XAucfoxpL1S+pg
u+7gntDP3+G9hgVX752rBM16u0RNwLItKlGKFtFKNISzOCG4h7kD7eFznlV7wCOw
6iwx3PtkwqYH0Wwdx8n0SMCCgdyqLyWZd9WvyjcOk+PeCUtwdFvmjcbeMbns/UdW
THAghP4vDSSOZiaiqUHcbb0JCOmCqleebfJ59LUBDjPIfq9SH6B/Asl9QXxQXdVR
yaCxwa9q6E6ttUXp4eNGM52AaL9ecIXRuG2KBmieRP8G0/hFoyqeZCgpYDJvxDqx
XivtyJhoGYnLnLN2tZOs55oSHIHbBFbGGZkOpopOcX4tN1LgNPKe9AhJtRTbVPto
xNXJjr0YE9G73YL6GwCDcOwA7DwDeutETC/fG3z42pcdQA1CUCgSWCNvIF8+KM5T
9zg5oGyma5VAzCsjiqaJ95Ct13oNGJWm2bDAfLVdKrqUxAvoBThbjktoLY6LsnmV
kgjmewE7Z5YSWRiW36bedXFmA4onLv6SNvhEB4W+VSOzH7g1U4wGxpG4TNWsZvfg
yEV/WbVVJCq5+t1AnXf46hhppr2p/Y96pxIj483bnFWi8Lq2hNjg2IUvPJIjP1JF
Hke9r2wQEdrYWU8XXOZMd9qAAx3IrOQM0yYbEWCnPz7TH06ziN19Li9Zm4nhG6gn
bsQneYQA/BcnvpttJhns34mYWG8c7TnodSLpMNpUfg5fc7YCEn6ieWRt+QDv5Pv9
/cxOc5kd9EUZEgpTnAGq3u2D679emS1avI7k4gfMfSnxWYfZTIkj34NWgInxNutj
tWRKHmp490mxlwfrJdPtj1oh1iqlyTHzCXJFWpYDkjgml0FOi4WRcXyUrpecLyOi
v91I55f1+EBC3O0bY4KJ63odwr9Al1Z1Qtbt/vBlpt5AFRbsfhka9qNr3f1DSuvL
ObRYiVd0jFkxfU8M5d5yD6dMdHx4Zb2E1FsniIxKrCGBMlY4kACMW4vzNXJBr6Ke
lP5VreJ5r8nijdfa7T5gFZJhV5PjR4BCxuybAvJmTi92w+ioX7lYqemk0q6YkJeW
jEPVAH+tLbOtKITYLmPx1lTiXlgKGNfXf2pG8OTXboHRm7jtfG357BDQdokJP1Xn
9H08qSDObRr5e7S/gg6YHNTO4O3N9c64RdLBPfNBKADBXjxkH7euvhuZGsuNXCAU
Gxx/W2CQvGaLXh6Wh+YKJxFWfvJEBJTUghNtXNl5bfsPfwUNmTje5REEnZ12aEeg
EGGfdL+Yh/LAbNNAQtI9oLYFjmssmAHHTf0eEMttWBea6uN0QbPYZiV2/lwr+6HE
i+aYw87EHewdwHmqi1N7bBHc+Bky2+qSJVZd4zXxgupqdhTWQB22Gvg6Xap1PJiJ
ngK/64ffUesco86dQeytEJowz81QweID2bAt0reFoUqPu78IJDTFgvbMfFa9I26g
NB1F0Y/3O5LYshXBJyW3e+hVgg660dMwqzNjRay7oejTrx6fe7R3Y+YzCNOBCyTH
sIeoLNSmVgZ8KzKDbaA/eIOca11IXP/1TZ3S/qSIzd2Mm2SOIegmvRvyZ0o8qRSh
0tLgc2oQj2i4ka52OLRAy+o8lGxuxfhWvWbAUv44vi5ykRVgiRklMYiw55td+4jx
K5nrxP9VnqR7P6NKopQpsdJPZorOdPuiW8EVmigKzzq8W+6dMJ5mGMIJolsA3nLC
b7qpdYyDL2d7Z+2fo2vjH+UxTZf9ve3TBQdxHJp6Pvc+iYA9hdteqoHlwTqIglNz
FVJMe7XUblSVnn1b25MI/aTTnKW/PxMWzG8muPvlw+DOevGPOSV56ys5QTz/+e36
t3siDZs3UuEYHuA6UWdxPaWaW9vJeU+7WYDRjCDz9W1Ub03Kz80ysXVkImAbFEq2
QZQBsK2c/fhs/ELHlAH8xkNyRKTX540LsAOGAbhkfQz8ylNBFfP9t0HU4tzqM7bw
MFTbBjZiOODcIa8mfRc0jyB2rNLEKA8f3LimqKkVt3V0Ps0vZFTiJ9A7oQeYdiCa
CdIvJKQLos2/sVWrZL1Gc+GmZSb3XaFhPzbecCYUlsDCmzMZ+QIEXc9MIRwnSPnY
swbYstRFx1saXSVNRcO7p9hkNSFhyzo6A3ycDCVaCvArSBaL7Y2w+/gbB2L8qg87
N1htpHVdlZbIY7yd++Pm5BDPPricPx3XZ6Y5D1j3TNV7jK7DzeCT7zjtT7WBGQFo
2fcxPWa5IRfbevtBfdARHCiXg7pI6o8ctswHVkwqlZyVff8wHCnvmw0IMeMcXp56
MWHq/Wmbm15QWTnKGBcmqWOuJyeQyCqlzTQ2jV9voJ5zVT7Im0VjrKT9rnOKX0eL
Pug9Pd3xORWsMPlqJv971RaXl+k3iV9hiu/iFT6lbjzYIRYts4Kq78SNdZLt0LiG
gtArrX+GY+gzJrIoSMuK/jjzEFzS8QA6JZsg1XMlwXpGzU1sI2DpKV6wacL1ByFu
TBBBHiCNZIHamPNWg8kuBucrLRGShqd74+MxeM8NPo1Cngrvn+EBdjsB5SKQYB53
LdjQ6eL8UNOtdI8X2xd1w8tmSZQcHXt5M/s+1V4enV/Mb7zrU39FGjE1S3RiHH3B
UsWdlPUxGxvEnDehLGV3LZ/x1rNUAr2aY3MGKrtTjFvPXKvobolcdo3Sd0il1Wvn
iwgxwQCMJfsZ7gOK+6+Isax3FOhFzKirGu3ngSNwAt0HtqEFFNkD3Gm719j8bTHE
sXtcnnSg5jC2qkd0asKqJq0MSYJREXV0/PQU8+RPsAJNQoS4y/1WBgPelPfMMDIQ
qABwMgHyIWVGtxNyz5KbzHf8o/ia0jugrqZn6rNfaBtxOFBw6jvSpwAMWyRwvEX4
+ztTr7UsMJJHysArKbxj0RkHZgZhZ+FyGcjoMx8ozLkt6+69QwQsY83e7d6ksGpt
crzraPh/NV+zoggMq5hKV5fv7TBwr4xF847OKMqlv4sBKT4WQD7l9nCu4GlMQURO
b+tkF/KBwuXDmZwkGoQwrYUcBjEElbnQ9FLJenzOg6FkACU+z6kfwzmbQ9/vV4p4
BdMS3q+J2enj0rGSA00qr8zx+S/bMWIJ8qimZ5OZrC5VkNin2gVWZDWGezg6GEFv
famAL6k6QmAnvT190j1ZRN2G10fR082BA6vPRQ8Wxb/1Jdws3xde0LTXudimHlqF
aHCPmMaEptEKAmrL3B/xS/uFM4e3Z9Ud0sTQYg5nnBKcwCpPJUtHKIJlCHjG47WH
EC+G5S9DadZ94cnXFPumaqUxyGYJo3kwK6AOL8rvRWOKa1lDl/pj2ph+6mYYfRvf
gHNIBAy4+fTzlTf+wlSVSi+b4gGiabPaqZ/zdJXxVmpImrj5/qolSml3sHvYC0HF
qqT146dldLzSb9tQk8/lSS0r7Z0G1KWU6GyVMTMvUeK/+c4LNslfaP7tE6hymbFN
zmIUBV9JP51G4qf1iXVUEcyC6apawpyq0HeHSLH48agIOzhlkmOjo/1LR4kW4FE/
SNWkES5WWci5Z/9y5utKJk/sz9VK0MSgPcQXjwW8xG4Istb041AsCHayfy1x0ScE
rj1fdInDTMTjWECmUJv1S4p1JUkkvnLIPUO5XVzlNNtjvuLWn4JxvzPKyY9SlU/Z
dCCoNMJROiUyxE4/U66tq6KCrL2ETTvJFLKVAggZAKcKAlnmqfoH/11Gd3z4XOOw
I2XMc69mHBd5y13cuHj+o9mjzK+iWERTKl1GGbmyVck8FTYxm/tt7h2Ji18dv4Xw
d/5EJaLXJlnszosaGIT1XFuxoalUfmkzJjg3DnC6k43iwYWYkSBTUFxvQGcfO0Be
bRplZNqKXxrfqneURWKHrLoyShS6TXaKxofOUkkcGW4IjMxglkaBYg4lxFeCOgcv
3xvG4PX5hxBVzI5GHMHIXWPGD6DeugXRIeixZHFIZUE5BoGbq2YPrry5oYiEeoAW
m2tSHWsfGPnmupS9JQjR0TyrffIkOk3/+JSL1kBhWV1oZnMz9hpQyB6ixMapIW00
RNnCJ+U4EU7JN8En5vIPy2FvXkdBvyuc7BVWkFfds9PYA4HC+cEyf8yf+GSuxCI4
sLxN4Vs2+YyUu3aFbozIzBiWKdqUwfKEUP8QSdp+EywWFdW09fiCkoVSioOSO2Xi
92efhEBIx3FBhCVt9Hsf+KKO9FMjQjypUM2C9PjruUbt5d8hOqlZnTpKNYJqoXyn
vD4Yx1rNObpEH1a2xh0n7Xyw2PdtTPnWhD29b78TC8qEZfu9d35Q/QeNiUH50QhO
liBJMzrtPtGWj2OSfRHichQo7B4w32JpIq+7hY0xPvMg3v32kF5tAqquBzczDd/x
hPLIC4EFB0p843RohvPC8G2/aHj84Ejn0O8oA9PQ7Vj13XcPzKlqWzZNeNVhhrCo
zYGV/hngHFuUrmyOAJqSzOzCG7+0pvlqYi4xTS14Nv76kMt5vL2YnuVZdsE65WF3
Qpm8d8+tA00X4eeovLa5Hzri2/9SQSfvUjcXFqHz013rfCxXrBTWCarX8mCdGwL8
9DkqmGvqYEgp5fvVfTX1XxlkOs4+PMDoM/70c8Paqg3N3E/I8tMXDlpQaRIMO2Uc
n1rb6t//K/azQAB6oDPLELbsSs7oqkJsO+7MlNLUcGdsNz9VhljD/NXS/2kyvwUt
+Cr/d1K2X5mGcYKiuFccuJU6SPq0+ann+7OYqzZTuVT148DvOzIU6N2Ge1tTbYPy
lwmqjdM1Q5IiXmo1M2CiMhExgydxiazWJzB7j3utmZ/+XjOiKNAKmv/XmFIhPoLv
aPXGrfS0EIrSGfKnIlB+ExlXFZFw+FtzNoyDC5uOGlXZZs9wa/6eSiFu5bUU/AxL
kAwuDHWTMAy/M1O0C1PuR8w9xilP8CaEk1gxF2+xk8bHh/JBotJe5ik+fkuMHgM9
t5VU1QzXKeOv3ysxFBQARINfDQa5Hp0Q2siLwGlchXTGubhQZ++2sZUZ6p7+C79l
ZvMnpgkRrhro7iwv26UMsAiOB8uhDotk4DQ4at757Raq943QTB7o2Tnc9efqMmYA
/auOwM56pBRfU4rDzcV6eHxuekrACDR0OVsstwjc9ZpDh/vEr+g/EO2MEZjtKNvH
zXhF0oHl49cL9ZLvouvAFdrq92YWhe2wOCUzenYDdvfrItZhCoyumvgJy2mL+l8Z
4Jhh+ktUnVL3swNlJqeO4yAOSwlIG7DnzsqRQFnrHaWsI4H53IDlxJG0Rk6ciQpT
stniMkkih4gHbIyouLwdji22QRhfD+rn2mPu8qxcciVbKq7Bc3OXhQW/e9RWWTi1
SzILoNSgSR5Ip7Fx1cwyUmlsq90mGqRfn/okuglD2TYW6EgVT4nzyZL8iND9CEFu
WXPXCpQX/9h1O6D0hWinYk4YdXzGPP03V+izNZ+pBAHyWWS1BsBdqCCuPZoxXBlh
/5G8pRCy/lK+6gQ1zvitI9Lb2WgCznpQ4yGzS54K87E6Ql6WHihjSvs1/ZMpdC2q
hUkfe4ZmjQfo61ylrpn3byAy8QxsiqfnBdz8RQ7+AFTF0FiNlUNXXqujVh95HYdV
9gGnTpvfKdomoXGKzxSwjy1PAxduexmVprGuNPzlxKSSiNd264xO/3zAxYnsBerG
OnMk1bj0aJRjrjRJOJcA2CsHkMmQtG1JzGPB94yxperbVQuHInEDYqlt3dCWzVu+
bK97IfVY2ySsK+3NraYkxKe47nB7fLDPSiuHZF5MxoHGqor8KzTx1PXCuAdCyRdh
6O1QBVZRBs4+SAiPs9SUeEKzn6CU7FuiKWJqT01tada/S5EVtgRYSMq8bF0P1ivT
L/HYC2PrBD1oZHkWk4Ct3ytrm66Kvo1HpWG5HNmyUEZ6gmul9T4V5oVS0SH8EU1c
CQ5Eqnms64wS+8xVFCrVtbj9j97E+e2BMAuy+x/igMXBHpmy5s4snMprEeckRlA0
GItDXQCqCneWNVfOyCBw5/KrP2JoNsXN8MYXJRPjC93mG0ud2X32ujhV/hrYUD7i
3wyZQ+GIdFpiBdOlnbNKAn4RDEMWuJDAZaMW8tGh3rX+WeMg4MKu/sF/Vf0IRgZc
Ta01prQ4RKJzS0Tark5ucF65It0OaGq2nt5Yqg6jBhyW9OvZpY3rU0JDaoevpqN3
uiVCLOMvLZdf6ViU58yo9oqaaT6RkBMjxNuRBWlD3ddlGu3p2WmzFDjkL6wlPxd7
pZgQTonruTS/RDyDil5bKvSpriqKyz0ev2E9geYuYHKvDIVWO1M8XDHq0LunuOJv
9ccbQd3ujvLBD3KjHpH1TUImmy3Ho4KT8GuubYhmjgY9OIwEXyRpM9ukwftPTMJ7
smm7KJelXvDSGPwjSGRY3c6hYjklxSxFxlC5nLDEuy2HhyJhEP1xPB3Fk1Azi/SV
mcyP6T1OX9nJz1KtGkQP8T1FR2HlL8DXmg6RnsDVgsEsV9AcumJlkWzNmVymBOZV
7sK21tZ4sPvUnmSJrjxD3tEn17EGyWy2iQKNQ2EJDr5lkeOKCgihrvY/ptOglei/
3V0tTuVFwZ3pQkpT2IJZQ0OzXwt8ZkCE3Il1g34fV/HFlCHkTEqGYoURzmeKDSdj
BJqYK44Mq4IKXBYTRnEOru+fLFUwWWDUxRQeyWSZYxtNUKme/rRwltG8K04UnMtL
9nrnwRUCbd56jip4aOdNmfmIrwXmXK4b0LdWLyY5lM05uU7yE5BrZfIWbwPo6JGz
BSCRkzoJFEJBNV19A02wMpBVA17BUVf/DoacRsxn5zmvXrup2KMgmM4/fAuhre+9
j7reL6+XP89ItjdVY92OQg6NGnS8wIgTw6Y6Ufujq4plIp4Zolqv8dLezJvtj1b1
wdAVjdRtiNqwieNfRi9Jqe4nN4lvVV0i4n9wM5zVW4tKyLtI7j0tgiPagvJSbnkw
v9NSEs+jsrQGBUrn1sUhOoqxxAtJrfEx9lLw0X5sQ3u1kmh4GUCrT3JMLCUhSrgC
SugQzQJnhq8G8JM/OUm34kqOlg+jmxhxq4f6TtBfy2wmrsNEj61pR82m/b05HLRm
SQPnuWKrPndQ8tOPnWnHE2OYxv/hHqAGvEjP0eSSV47c0u/B6hfxv94OfGC0HzwA
77qere+0gFtoHSDGmTkYX28U9/WqCth4yJFHf9wjteSZy976kfJH6RYvD3mrRn9U
+frQ+z1loEYeoznPFUT6d2jcq7t7NX2gqZNC34PkTbgRi14pTS1suo6mRCPy2Z6G
Mt1VaNpYO/PhujJnWEaRiNdH8Iuv4I9+hHXYW1Fsss69zIDTC4s33IRar7lovj/W
PZr/CsArNiGRgGbOyW0Bwzu0dw85G+UYrwrBbrGWrt3sb2DTJVsgdcewNfUbf1C2
z/Rx1EyjCur8L9oY13rmvjZinAvHZ/iOWd/BieTWc5E/4mvVvbg7X4LPklBxRK9F
4iw2eZkyaxtzLlSHEguIhMl74fV3XQmZjhcFS9PdxCjfMxsHcev4G+YjVNGmi6qA
M4OKjtUUdMkEQObn5fvDuRJT+RHtctLqCKgoIz46TRUkiGVgBQEbcclJfx7/YBvU
MzjuEEtUnWQtqq6QfSfzrSJQvR1spBPGOCzotmtd6e2t6JpfztuHLXwXUg2qk8PT
NHDhXkoblXWIPAA5qYRpChB1nopqGn4Z20NO4TXKRA36IB6OmcLcf9+Cyx0Mrm72
iVH/DOSGfHmP53heoDI3cfGUJPEuZVMGjxDoUn1gAdH80eRcNNNHyZt8SLIcd8nc
8npRSN+zBi92edGK2d95xWJGvMouMCIncP2CKtMy/kZ8tC6dFLjz9cdYSEeV7bCV
QcIYN2eZbLOUZAJikSdZwbUnt7tWaEWyc6Y0pTZMcmobrDgCFdqFuWazAAOyQDH2
72bbS4mNYUEMs21tuLHnlI9IdJNKRx07DQCOYznKD9vXsXKxb2rkVkPehpdB9YxQ
+AJL32UxNyGHGJ9BMb+h3M+IUP+hOUFAqGcqt2Dc2jFc9U7BjE1osqTf2eYDkFFD
B5SI5hiAKpNxFvpBihxrd7sEUoVLsOIsHIUl/cV+Z54B+M8Czp4+5zUqCFgO2o8U
HipHGg9Iq0DLNwmzQgVmRxcYH3m5DXUDZfS7GdDzqotrPQNz07sUWkCrK2hpW4mw
EOkeHslQcILG6b7C/k72zya31ntOKy6bJZbZlRFdBrftNTbVhmup/KUIzW6P81Iu
2Zo2xrRNFJICMfEzwvu2xNZiIbIz9d4zQaRfEb3qO9OCq9eCmhdXvd3EBLeoOWpJ
Ep3PzVnxPI6CH1gidJdnMvjuKIPWCJ9A9935EgRNmGuz7N27I0hMiuRCPpuswfJf
FOlLYGdPastBl3QwZygi4DJPterqQaw+eElRhwB+gIjJQJJ+VQncrrUX8qIcZWGk
mXEPWKpTFYIUjMG6s++yN39IY7qSqN1bQz+zKDbqRBjxZkuW4sm6gEMWbnsGfoIG
zmofuiTXop/q9KI2GZsomURfGSb548ymAKERgmapIEcmOBVfXo6MmALVHsAFfyfO
2BZJ9tCtAzsITMBsrbUISFIB7qHVZ5kja7XNJzI4wFLN57CDcBFC8gXfRwhbjhId
SxnDAhtS66i6msek6Y7obtcL7YK5SMAf3SW/rx80gvBDjeEsApuuWyri1c9Q/gPD
qn/70C0Ci+xrFC83l/ohjM6e80iaCmzq6OFnKa1dNvLPEWHfGjqtmnT0qaIisAX5
tt9eTVkQdNH7AXIwjKK8FJIKu3jNh6uf/aqOZU+bOjIIkdl5EotvZeveU/MYfkXt
9zXCnz/APJBpCLPAEz/VxU8dqNkxivAtiIi8RZeE04KCDpcby2QVA6jxVrNCIbHh
nrFc6cGGogCWoGTTn/DDgaZBxqAYc+DAmZXPg3wTomlASkKqVhdm51im8Nbgj1uk
F+gBmECxsLTBWJgiI9HjtYySJ/NR3Eb8MQv0zcytGzVZ/GqgAmxbogsLtkemc6uv
55f2cCNbwysaBD3DV6pHLg7Ud1DAee3V6VL5EwubOZX9NF/9k960ZQMfGLWXzKSE
DVEPEZaYarQ41LG73to3Er9XQw9jJd8ksqd7HnQ5FPtO6I96HmD3i5ykFuUxJdg5
Uyh8LSNnSQ3cCEIwdH19BHbQvYFy2P+f7ljIcnAMsJK6QvZK4o8XBv0WYC/hbR+P
35zI225iDP/6QSrkpqwVnZGcyVM4qvdfUunN5fAzqcC5E0F8nPJj9htkJjFbpkn6
nUSur3rPHDrkbJa//PcOEw8UleeOUNJqT9d0Sr0u4gjrb7wyPYhIf8ChZuMcboXU
JMtLK1cRFKpW4Y6CaKPZn6GmoIHseKk/t+gn1DnaS/DZx7NSL9IFWG2TR7W7f6dp
3U8f2s2f0NeVzhCt1GnWKCWHqy6MGbC+zLnb7XU/oYugNzHrqBq/WqQoT3OLoTdI
onEeRkC+o2UdbeWzHipma8H5JTthb/7nDtvd1wNxV+gNzhBjgVQ+OHFluxxrLb3l
V99xsTOLpVpl6vqWEptxVB9pen2m4rslhXNqcY3QUkXNGZvq117ncedIEr6cRf6X
2ySyRjNM2jrfhzAsQ7eiSGKGJ/TSoxgLiHDWA/9k7wvHu/pr7/kRVvN88rN2eabq
wyhf6FEMfK8gmU6xhgXMz/LwBi7/Hniqjz0NhdUNfLXLCWvy91oKbbdSXlGuR2a0
794/ZRyCD42w2tEWBCsedAlMx84CRNVaXR180VeA2fetcEGclKSL7d0MNcRSvlpk
NpRrikqV6EalWR6NUbWqErx4V4jehIPR4sB7Zbk1bc2wXEYmPGLMVgCOq1AyvvJI
IGmgq+wQj8W3yup2FDSNtJSh07+r3xVCyG0szjXiZAzYav/iOwIyFpV/Vp6FAnDt
6cdfhN3SFJc4MvN8kSFxAIMyf0zJY+Vs8S9XXZkqVCcBDaMJCqzvBIBydn60QC8R
uStwWSgqoUAJRBkdsD8H7obXNzFeqmMGBqtoogTP6y8pnyNQF5D/nJOcZolDFdXJ
Yqsw1qZGZ/KG/BYy1W3VlDU1Ukz0M0xyTI9t9J1bQswV8Az9tIRuoPgVk0GD4tYm
31bkj15pskj1F+Klwe5wFb8co3m8oR5qgEKhdPtBFbd+feg+xiRRgmdZCAVvZEcj
tYZhfb6URTs5tE+3Hy3z+snmWku1lmvbTDCDakPnVJCCo2ej4t/Sekj08dUZXBXH
Mb3Tr1qShRAsZdwBCwE0YFgxgGcNF/D8N7voi4EdHKOA+EHT5Trz0lmz2WO1d42i
gh80oOEvum+Ou5bsQ0wcEe9jmDHg6MQhEXKxveqWo4TDWkNOwa1QeYxQLJK46Knu
+0clezwmBnOdGqPSL8Wtuxo6BGUqdtsrixJG+C880u/nz3IxYOcm+rA09ReBxCQO
/5A+pj0ZFXz5B2duqFVthqTwRYdLsBYjqWBktFC2It3D3o1hBNlMAAArcsLsRhUu
k788HpQu4VLoByNtWqGX8PL7rolQEvhJXs9qB7orthxbQ+dyOZAIurvRKfT976fw
BbOnS3gLdxyJe31KryUsaPyqeyKb1tfKdKS3Tsel8IMfbHUgdoIHWTcN1XJQmSEO
XOQegllMBexB2VrFwZcqXKKKEYLqL+XfWQSmSb9zZNNQYCplnmQCCxaMmOoZ3txI
O2OD7vTNju6DiJ6bv4SZq/lVuSBSlaw1J/epSbodgMIVkW17Bx2jm+pLWJn1Ij8Y
8zSEMaxMvZlP3tubAD0x+qT94Pa9I9x8JnVDDgLUwQUpokgOg1Ke6oAornGrNPBn
FYGNhYbNUZc6qTgKeur+IP43+S+J2HzRXwJxDXPAFGdsVZoTStPqFUxZKKxLYva2
n/JhBI7Pzi2ENSDFl3jO2VVucMyQ42hQieRT+fPH/fQ2dF62RAHzxmC+4wERPD3E
0hod/gCpfUffQQGZWrLxSTJrzOy0P9e8UDjbLYpv4IdxRnfYm7WkaTnpYw49tIZn
meAt8D/wBfmETjJ3F5hy4y/1f7tywf10Q7YTo4XOUNe9Nrzr5fZbDKGVXOivoTFs
9Gt0yJO5LSerPYtFb3DAoU1Ub2HQhxy/5/e0aA5milczQdtLwqKsk3Cvs82/M39b
5tIVfIyo59efR6VZnTZz3YniVTT9W2vBJwPsQJ2aZ7cDHzZft9m+Ie2eqAR+WBXO
Vxllmkeayp/5kNjAuPE3IlmyXHIks+gxzsCLflK5CpTtLpKr9dyex2bHnS28B1Lo
DPZXrtRBSaxJR0rSGk7b66L/jjuNtKjvOVR+zJLVQx2HTZ4Vs4d8AkN1MlfjQwqh
bKAYdodJZvXOqvg6/oBT8p3gy18pXcAdy4yjubjwwiRPfk6cDYWvOVIM8lFGWXSz
zW/H6SstXRlAjd+LhKZWgACu1aWBAPH4mIpY7m9P6fLfzztE20YZszpSd9MI1JyT
RxKEKAVStxAmoajyghVm27r5n4un28pZSIySIKM82TFv8F45SzMsu0QKYZehVn8N
D3FIdfi9wiKR+7cBL2GivYmKh+/YCGK9BVPVsLCtZ4X4y4avmVv6QmUVjUqa6l9b
lx5gTQy7MliivVXdBikuGLu2tQ7ybjkX8uBFlM3gdTqUVRQBOm9YnP3frFvQdAgF
GcBijxU2RX1tlG+RlpqaL0vACf4Il1t+4Odk+E2kW0M7Ur+SE7Rud2Fl1GXHX1E5
TqmkRmFf73lNjjFiQlDFrin1OPQ3We4h0Z04qdll/NnKQdmQrrRjWvW/9p7LENWB
p5qjQ81Js+fkk2KZjQdAGtr5HuCdWilGBxD3c+2K+O5mKg8UywfgIzOQNGUgdns/
usO9WkQ07w9s+6V0YFM4jQ9vOAau9aztdompVDsBUMaBTJYJiZLSCUi0n2Y73F+Y
e+fEiFju63OmHHb5qTmuwffn6HFIWbdPIqx5YZK+P8LmqORwTQXHw8j7apAoPfEm
C8qf1WsnJgTy4N/P/Jmexs8kdWO066vTg9ir0kLMgSsM+lpb7Q3GSIgypEfe5OGP
jFqTBkVGYxlUiYRYpM09hsSwgdrq8JSvgvM68Nua3dw6NDLGV2RVj1/HAqrQx06i
KDa0iJI2ebTSsWpYH6jAQiLGS4EJINj7YAQYpZ5X66qPeXWBxDdB2XodmZvpJy8G
eL0NCuv/lLNPu6f+Ndr2txcrwyAobvY8Fk/RLn0xyWw2V9ldSyTGvP7Q8h1V82sm
+Xg3GpsVLclkcgCeNKNRrkwvApg6PbwyKiGXqyVNxnltCDg2LPFw0OlWX4fa5g4h
cx9zSYorYYt8AJ+KJawhnwgUEbf0PpoyGwMyuS22DbcspOqsE7Rjbu2UxzjABN62
ZemuBSRiju6lCQz7RPzIKbSorUXeY5p+Wf9Votd6JxBJDp5qXeJgLAy8QvJrVK7Y
VwnFi7fbTuycC6xI8xJ38FKcCDgEuJHKM/ZjHhiJyvDDnJvFOARJlzIVCpAKt8NJ
ihnmyrFiYO3DlGHz1+WWFwB1KH4Q9oQapHWSqIEWYmEATyjcijPudYp//5SXw3Qg
kzp1Z7hi7GsumOuaJuAEt1nw0Y0VuXKlWFF0D7rcX72qR5WMCjrgXzOlTObDc9Kl
WBRofnqK5fqvz0K0j05nRcnPHoHpc+nXbeV19tcfgseciU+9ObCakcz84/L7cLwf
AKAgdrqGyHMmkGIq7DfFgqrDZLqn9wbWSTLRbUMmduLA/GB5ESWUr6c6N9vkILFZ
9NZ0CzMZetRmj7eE+k81jT0yvmcX70LO6qetINQNWLaNkhl43YmHdXHROdu2/R91
uBC2ONYOQdX1KSjB/ehDaXM7EqnTnPA8Bjh0DfC9tsxmvH1bMUCIBNhjQ0nRdo0l
8bO12HyAcMZ8LP0LoyflLTPvnEotueW7kDtnkR4dKlbH6Bodp/sPgcsHfDJ8Eb0F
ZEOKipqq4X/ERBHw9eFyy/lvw/c25Gqw9c+SL72cTkplOLJzqkCQizVWpfivPr83
sPU3sUf3wu3zdsYS0P1FOxxOkFDzqQL09HMMVpKD3akzeRSuh6P6c6Q0llpHJUR0
ypYFNEqq14nyalT3c2VFk4n5h6jRsXgsfnuRi1PSEerUEoEsz8uhPYIDcHFGehU7
/ctrPdu2aN7kqvVBd3/6m8iUOJc18KammW5ptYkhFiKxWbZzyvFUc/fLdD+cMig5
QJK5nWP6g+IhAsT3VROQc9m/r1N8dqFPDrNk97MyF6wzWbm5qpyipfl2b1pi7Ru1
RgsFYLt29wmi24hBvNN496PXlb6KYV8ms87UYAYBaZTHe45ws95oW0WmzRSaxupw
dfttY1dYF52KIjq82hfzYX/4DzfvsDd5loof7pDZSWQHqw2eRqbFWC2wZqq50Wrt
4vnpyiCM05DscM+Cs2C5WSC1C/0LKeCKXob7rfY6SRHi4vaPwg4vkDxHoWU4+QX7
MiceVaKtZzI42OHRlKBVe81Ik3h088hubwFgDGDDClnLzsNm6yYXlBh7Ig1rQ6xF
psIncJZN7BDM0PZVrWOMM93xoNIG8LzP9BfcKEnv/3E0Wuc382SQf6GW7eFHCmlw
J1pNVKGLniCyc74TtbwQgiV+JjB2lvYObLVTIihcjeW+/anH3pNxwOGevX4KxZZB
LDMJpkZiI7Vfk6la6DArtp9QMbnLkAt+XfHvOSgxr/N6z5pFzFDU/fKhWbeq1XiB
XX34XEGjGh3WM5+LgtiN2AB7uGElRaODzS+TveYkF/wX0EHDNrxWyMKbV9srpLxx
JBvkAW7vKn8vgaBvxGlR9lcKmJHgSSQfkyVjN1ZmXdqMTKKnq98v+cGci/oWufzW
wKE2+HzkPb1GAK8HWWqZh0UZBhU6xKTZpSoPdnqs7XkqYDDo6Q51x+4OR/Mg0ANY
4a6jLdByNwvzoZVcmqnYCIJxsFjmpsLYXZ9SwMUrQwlz33xa1bcAIBKsCRBI05Tk
xWUMYap1lf2C0Aj6C/sHhc+t5CWgupY0pcANpEet59eJnjov38hJee5YO4yUOVwJ
wXQwMJjpCQ38whTYd+fVqYrAKD5ERnwRfu3HDAo2X+0LavhGZDA8owMmz4S3OuYU
+Y1Xh86bTrQpQnoSQJotbZJdYXSPNvw2IAORrRw2h7HOrJQaqjq9GLr10xscnURT
ndiKOPcM+EQK1isMd8tK2R3JAiegcQWCj6rTG9BZaGsIdmVmsnxny9OnjeEbqTZY
6gEn129MV9XmoOY1afxbnT84hCsph9nP+PnWYozNDcDjWyj4MJN/cHekcG6zMFyo
2wuMjwbSSpb+mjTajJuW6GqDioaY4u6L5vn/0w1lR5kS6Zba+DoDMRfsZELxHbPD
vDBWUs6WyqDwodrcZu5z1QcOjdhO4RP+DYbdhdSNXrBBd+Pb8cKSOCIfvyfXuusO
kjKMhZeO7CDX82IJjZwMrHiPHmJIMwemFFdhVPWc8g+YUn+T17Yr93T4qvIhbwh3
4nNFMFlMgOd6EaEF9HifIh9qJRTeUPg2Wq6HrxfPGb54VPyfcgl5Bw8qyURoVdl+
Vx3Pmsb8doUqbgfGvlYGG5ZFzWwTLPccNQfiAEkYIXe08tQn7OgVXFAL0ICqT5O7
NItK1FYQ1EF5Fovkjed9ykXUDZpoZ3csBCRhn5ChZLb3PKyyWA9Na2r6tpMmgJPV
hSTW+DW8CPehFwBdm3m8C/8d4Sb+P/A+0/I+PLVulFYaKQHpPTW6K0hrOfYXKNbq
Pd9VYJy/shY4BynHpL+7bJxGuSz3J51W+WczTaWRoLmy6a940cccpGCl4nyzDF0i
p5NHF3bGCe09H7Cl/B87sVvILLM86M5B9FLi5tmDzWcDoYoR8UGcBNPwXlA2SrTF
JHD1VfKrL9O1Uua4QnGKyv1cev1c7ETU6eITRKCGQUDIIhZksHExeo7FZYohUtF6
cy2PeMhgYUr6VaX+pgfk21GOd/w6cfnvGuepvIvpp3KF1Lsi60nBSo8zpZ3oqZBY
kqM8AzbIoRR122yXm8RGK1IbvP7HBlW/9kJVRfGvOXUHCBo3kMQygTRlAFgEpSH0
wSmpA6PleLECcm41D+dD3qPar8NNq9WWtQAEyEhAU//efC++BbziuaAlCVv1pjNL
SWRcju7RFuAOB0n5ryieD0sP7vYimZNgRuRi8MC/DPQH74BymwQgoXpoBiF7rlBv
gZmqbjCRntFNpKpfO4rPfp1DEzG6ni3wd28EobNnMH+4Ua99ghkJYRrQRIbFc/mT
Apmd52mYDGpdgM5jfEyhsV9zDJJQxuH2a/Ep2Mzgzn/w5i7rjEqK9H9OnrUUwaBz
7zogCnWpzJZdy/JrrkX8NAIGCjWd1Tzvs8n/as+kaJgAgTlpfcSLVYmw11ZScTp/
7meO6PyFTi8ZVgks8ZRCsw1Nbmkrt7j8Wcq9BEFrQS646B3UFjBu48CE7i5PaVst
xmoGwi9CSqb8DODkvsgjv+TytKc3vYrC0T7v/XfCr4h/roXLEJEU5ChH0YFNkxQ+
qBc9k0/csNVfMza+rCIwECJyEcExGcHxB3VjOesFVOiE04VBsb/Gaoe6BOmuU48c
JTralGGINViVqD8thqO+rRMOSJh4lAonKHtGWDNcwCXOS2I/rDx0l/kpnBpBQM4G
iRwej1fkGQSFOxYidCkhCtioeGMXBj1jLJFCL2441JkkLNtQr0SWYJ4/vCSKJgvu
AECpKRg3+A8fq6AXgPwRaXAKvBgEG+m4CoaDNM9CLxbw5mbh0SMh+zVWijbWbSLX
95csXJ4obvrtbvbglKomUCnRrgudods+tzSxbnFrrGyxBbiTYnx+3dGITJ034aY5
Z8kTr0fz7F/H3Dk7G3KVlCmehCLF3jK68rbZUxyIymeU8HhCILip6SvXXROpk0Wa
QA7tNw21WQV+NWZ7FKqWEmbCNoYV4QKNzIxccU5UmgctD/rcdVec3XOszB/NeFpY
hz3gqOBYkZnQHgpvsO/DD9xupFJtbD68mh5HU30TxVffa2yXLPO81S7DpjGVqORK
yLZ4hFyuTrx8qbkodKuJfT1GGCfrX9ucxchxD5LRm1LAChRLbFH/ZTgHUIetF2z3
D15nU876ixYShkXg0FGoRvQT4uuSZp3ZDSNbeHHd5mpmz+GIe2aeVXVTa4yVI+Qy
2UgSXz5YFyrswhSLQd0zU2va0ACe8G8blfYD7X+SpWkCF8xpCJBQ7a0Nuex1apHN
4NakyK4vm0KoNXYNEWJxSrYzCct42u2m1lVL8FryAl2O5JZBDVN/pPjS/6fLWAQm
8TKTffI9u14Pwf0SGpnczn+kFUTzSIp/WmLa2Y86s4xyGwAU/kfRnMcQACo3yGNJ
NozmSiHPLscB2Sy6GpX6oDoWVR9rXMhhgS9t8YLU6Y0EAtL+1f046S0lIgpuuKFb
D4/WwfGRfiQ2M4boR3Yil275NmdP7zttT9t0CKk5xDGRjvv7/0V2EpuwiQKj6l2t
rDQ3ncgUmNTdfmHYdzCfvv0/eWoe6ozTK3RUmpevvv5Oe7OLFp1fy1b7+dS+ByvX
8r/YpOrKDnlAKj6Bh8fPbKjl0eIk8ndrF6ctmDZtBn4aNeYidwLzzQcwNHAQDjvP
+2OPZ3Gdovuua0kvmspmHjDRJHuarcmRYduaBStYbuvDTbFcm9sgLGe/rmgcBB6e
Q/gpPlwtH1xxHyrS0gKGAk+7X4xE7XTxW/seYymSdFcNbsJAqUmk+L4Cvjkc0RPx
Znj29MMlzClAji8loFJMw6AQVsCrTGq68w2de9pAU2GrKkyC9iVFlt92Fn7RfuBa
I3LvL61O+14LJzEk4wDLpWTFCVLWuvumkNNhAmNJ+SGxKf0w6vAW2vDMdYt1XRQ2
fFFkdJrCqQAYd1BWNveGQ+yFvWO9rmH9LD0EZUbyfEhL0uY0J+lz47ZJGWMG9M1D
YEudJKcME3IVaNDRQEMIO//37lj0YRH2Us0k7+Ptvm+FDBR88JYhb+6bgBPQDzHw
eWjA/yDQVFkYZRc+s6r12ItvYoxjVdPGD3hqBPEgqCFsw6IIg9nYR3h/I4/8kLbP
FjOihuKZQDPQ88igxY7zlbB2VOBJ/jbXYrG2J1u9iIV2IEtXE0GG/mIbNUG+C2tv
5CP7wXZs4fG0Ccz1A/47/2QmF4mHmJkF4UzvBlNN24k2AoAO3Np7N+YTZhSLjbjF
/Zg9ZPI08mPgkY264iHy8vQvUfNfgV9TkOPxkCprGy42xgN5fO9jIBd7VnnY6eMG
f2jl/hfWgteiFu8cM3w5UfGu4H4DgzL0wxY8VgDyuICVoCvFjv4GiCPRTvPy6+17
ZbcRM4KH8ATgTGzZAI2J/8/XySEZegLb3OgEJKuC6buJDD85AgyIzvOIuhV0TmD+
JG52A0MiTssg4U9wIc5ONtENDz98Gnc76DkZ2ePgijRo2+rmNJXqlDsVeUnhqmHz
7I1UkASNbGheBa8FKRpb9pvrLIZkvncXwXYbQ0IDuz1VNNwZB2aPTdh/thleeaEA
U4gXjRJv/rPgWqme9KFMv/z8xdF0zi5Der5gJ1ON0BNuig73SbOBKNLUXUHPLytu
FVpB52Dh8gYGVnfmbdf1y4GbEucAfzrQ0vlWE8GThnyLHJrTDY4AHanElt+mexht
0s+ETIE1Ny17fPfpZ4oxCOMlVrhOcgUj2O3JMp5UGsfIfNS0p2DufjkiOMYoQQhf
9cKKIDnPwoFbzbEwT5PvjW0MpAR/QeJ7d+SbOtdzVlRvcAJ6lMNg9cJ90rneAm5C
0aFeRJlb1g1nt3yEXQS+iqlnjdTPi2MDXHOMGES5xTzeUzreZOdcagJR/9XrdwnD
FxPgx7mIDU1QMHOVdiPSpaKnchN7YLSynMK63UKkel6ZWRiTOv378ecUUQvidGKx
SJixHmzGqA9vY1nG4Y+qfChtJiFnEJZd2Xa3oDWc7kWLc2Rvd5evjlfQM7opNSje
QVU1N+c+H7ZFeHqytJNYBHZDBFrOSrkOEqW7EUJGdE91jRuW8S65+/LWmL64yLay
1uJC8dbQPUsMh/v2v4gIqOxHJqTO9BLnZ4t8gkWXyBJ5geKypws1ok8Xr9Pry/hU
Wz0t4+iKavAOQMuzqQA+hIAgFqHEW8IQ2PyMn5i0Jkx9t99uYiWsD81easfUe8y6
lLVtwxdl1PeV9EoZLhxBF9QjZb66THSPxZwYy9HZX2BLglVWh2IeD7lu+eudadPJ
+/n1rTOaxTGJ/CNh21xact9Rx4DjVPHq1SlkMnWOXMRZb+MQ17rw/WdYv6rKG/Vf
M0pza7QUmS8Mg+hMe/+DU2/Z1RouvVcICsnZKqm3OYtnJeOi1dADQDyKNESIlhBt
y8ovPaagdPn2IFMBbRXECiUKd5P8Yt0eaYIbHneZ2EAYdMPqfa1Esgo1AwDoqZxR
nXQ+NMeCyfz3OBodp2jPDVtSvhJzEXY2/1+1zSXvzDzrGItLo+nOnF3liO1emntU
VGNoCeODD5Onx1En24UXbzZIipEhdOCjqIMsk4uelt4DVthIIy4UA2W13wgQnbcP
8h5zxq9bSgu//1aeIraHXAE65qFuk44mr/GEq3aTAPJmLKLVvouUB6fGRrQ1Ik0p
pS+DqUJZMz0xwSOUPFPobD3QNwPo7afTdHHsgr50UrWko3aYL/294CKnLcP/CqkU
93xRhI7Fab4l8O5VbWFSHuTA05OAngBrlbuHYufBN2fN5GajZ8dboAcpDjPed2Az
azKFcJN9407uKfTNJfZh1zhMF/LBR3xkvOuo7yC71i1Z/q6sjQtM+L7csM5flIwx
qmALHd410VajqVsimm8b2ZKgI5vJb14KFPRaDMpPCbdp7fAD69muBFMfysmlOHVL
W3l7sgo5uYAe8RpsD7FFyIuuaMqY4uxXMgIxG0Mms+/0P5H6Zr/m46S+33mjqRqw
1zqEW98V434dO1MFnuWIC17XB4hN0G8wHhrnUqr+9WL8ay7SCSn6NjZ9VUuf+Jqf
R2fSWt1Qj2+plALEbcCwHqTNt9s7LDukim8sh3vCk1LNci08OGAikPF76KiswXBK
tSabc45x6x2Xp8jQHixly/MnCWW4uNK4JUnidhUGZ2F2uYumRW00PaDsvRkNRJ9B
QOFaEaHQmW6ThNT1Llz2RyL+aywZj9y+M3YWwDGtkJRf2JIQav1rA6b7ID1+NbcL
PABpD1JFM5Sd3/CG5Z39XwcVVZCSHCNcXvx/kRhXR5WY307eWDdPVhpXPA3zo0/V
soQRbOHrNsuIwlVNrz/dIrERpe0K86Z9uwczW05sQw7hdC6j83BNJcHZ34JfWBcL
w5ioCd5rhanpmm+2fD5CMHi7ZWEGMHJtPn/snbA15QxsU0EvV9TY0XgN5XC2GVX6
vW3oS5MrWsxdFe9xcs2ECwOI6QOaZqgq1XhcopjII8xedRXXhOnn3gs3Z/A1Xjkh
LptAZcx9350VhZGiXRZCe4oNhcA02rriMxvkHDac0+s3weoao569voAX5SfuDvd0
oPuhi51pzgO1EBaRclRIRAJIDW5tBFYyQ1b7HcbfMvxEaymtm+1SjNfO89VJlsTh
mD0bP4R4ddVUGdnlcYm+DDRglmFgAuMELaSqjVq/PI9vcErZMuNAF5mUkaC3fB12
+Kj5bm9nHyoSMTwaHOIw5UXDK9SJG8Mn/dd61enR4SYi7FXGE86xK7s2xAO7/X8g
67ZaE6WhUsx8Chhw4WBPoV9qOHIALHNOpZCpd8MlLPZlWLFHPDtW8B9ZxumJ/YGK
A8Qw8HE+nDgTjMCYYzwvuCBVnX4mbwvnK5AjWyi/te6MPDeALNnnerWvDT42IKfn
fCZNuIgGcOsPxlkTaI/qdSyluUg91NGqqckBP4z1pGWnWCGc3JVIP5ZhwK0mjMSy
quEa8nGGNqiLmyXbP0RUNPhUPb+08L4Q4swEccq9fMUKSq3bBKlpZ4IaeH7MnyaJ
gylYcr8jcJF7JBhWr7IUqdHGs/CKMQZI3SphG+yK6apFCGodOJaJeMl2+xRO78HF
SHoa/LPS9cuuFEAx01Vju8M0dLUUdpZIWkznFWBCJhWiwlCrn1kBsU1B5jlU3r4l
WU2uazAYdQXCYX7NUaNhVKXVmY99+vr3ukFmq+/60EBDZHzHHfZtG1+h9R0AwTnF
NIXzjScKal6ZUxrEojUIqWxtmL5RhrLmmbM9xdpeP+sNqDCpzQulGpevWVIxvljn
ERhLcCt4+lduK9D7lhWUnOhHg45IKLbZuP6JN+ACdYmBqh1zPkSl2Flym5Dh/IV5
yXiSvYNKGDUuu0O0VsEBBb6MC/RQjZzUs/MzkXE2wMvMBYCGHV6vie2lkpePem/I
uO1gWc9lZTanW1gCk4VekfSksOSbYqSRE7KwF+DVwAK6uqY6Jpz8yqayeBKwxLuR
0aNIU/SsUuiTpIz4s1yWUjDd6TZkeH9DbDXiCmkp91kwG7TE8CQyn51l+Cua4Nug
f6J7Ye2b3dxuWOgiTXo0u/nBahy9ihXeqrjb0GnO1lgKBZf8Nr0dSQJJ87CPAVuS
1AEuvXfkpEtHOqR9bdke8sh74F3EKqZA2NPXOjNdpUAjFH64RSX5jMBbE8ffn22E
XJRnz7W11kEzBGkME/9icFP9HYF7CLDodllYgBJiK/48F8UemThaZOj5ctUEVtWK
2y03mUrxJZE8506Jzf7CMc/hwD0A5JubCTkIkhLOfIpJ67iTF5VPHTCwH6NGludQ
F2HliVVW+7HwX2o3KTH3d6Zq7n+maPFl7GraTbSFRX5OSF0ScsN27JvRiKHDSPi0
pnMKF4XGaacdo7s6sAHCHvVPdBaBueZEH7NEvGdSz7FkLPh/yXlOUuAv7rnRi52d
aXW0cojvoU7xB9Do4S8Wcm23d/6wotOnuqu2UUOESdp4b6vcP+At+nJlKdbRwJ+i
WqtGOGcSCsOhIgEBR2m0SE2C5E3oAOERqN/e3ml24zoIBYhd/aRicW0Jn+tla95B
cdZIH9KJFrHH4Wagmpopc72UUKtHIW7VEnWOAEAyx7kp9MntQtoPdaiFvUAvOYt9
6xov5LL5sHq9HdI+Fdpa162qB5Vl+vLWNpRce1x5qUmZfkQ99R3/oNWKph2v4RQw
8DqJB2Js07HqWx1Vp46G8m9R8/jqALZoVf3jUyUfoMiNATdn3J+QWL2+xY/U4ldH
6LjO6xqLJFSj1xPDEbUEGqckU96KMkpngMRBCrapZ3guTfbv95rdMDCgkgraQa4S
GQ4fc2C/5MX7Ch28YSAyVtCD4KmIuZ5uNlCweD1NTmJnAiDy/OHVJTTQh7ODLi1Z
nJWSqG0Fp0phLd1FzmoQO0kXO0RFAcCY1lGWaQ+0qGi+LmcM0Vdhp6RkMuLZDiJ0
knA3SQWnJwP8agbOW7dRTeH0FvlqsBiLTuIYeGrjEYwoDZvqgwU95pHPQSBS6btA
1SFrpWqnWkiHq8vKiZjCqZeBM5A8smOCDqp4nhr416hPFNbUZ6OKNFuz7gT+sBZ3
gnsZFNkF0QzACPy4tuNYL2+n3kQhx12XWYYihsDD3usd9y4vBSy+nk77j25yad7b
rWKwqYYBkGFAHl8EkOW6GMwGJr1FPJ0Db1qcE38MnQtO3db7dxGXjyXUvyQf9XUa
bP5ZWb6BQ1rO/M6A6f/QUwhnEbSCaPiGIX3Hk7ZpIa8HprYoKBpg1llS2rZ5czfz
tgvrKq6+RFnyjbmIc8tYoqC24Osvi9GGwRmcIZ1S3fwDDABni9fMFZb5KpVR3VPf
XHhyJfSvy8DvfnPU8+3TvbVJK23UwdQwrnzNitYGJLRrl+K8ugENsdDtOzwjxUXr
cDjGhKUbr3C6KRq9DH0xB/mgUmDebjppTrW7mrpNazkYq0kwoNsJcWNTaXYOfK+4
UBn1rbGJW4y0s2yYvQGLMNR/8HWehfY7CnSREMIiNxI+5D1S8FkbQlIk3N2d5kpp
tRIj5fOxkVHyu60HjWoLXpfVj9TXzAmyphcMWmyCQ/izowHaxtYWr07zz+gJtl4L
jdykLLtIfSewsAlXpPr5HPEJXytGYEvOQxB6AHexOYd68lvDZwPDJg4bgz/GIu7T
6pi+spo1JgYZ/eOwZiyG81OAHembqd4O7bcuMtowCyCmIbebTgDqo1TMEwYSgdmv
fQlUAvvSFh0MhZ9Cl0/4oYl3Yo8oAm0OZXeZoQu25wzbfI7/eTLhpSyGVh7sz8M2
WTsdout6ZxvEUhry1N6zhPs7z1oD7oIK/wdaegc1shr5mn/8UvLl0ObMnkjLgHkR
3S5NwIDf9qTpfmxHLgpk8hVbk2VoWD6ug3X5TVal6DSOY0TDj70rhoNXLJbQ/PiV
53HOsW8FHIU9R5iBCOKFNA+mmRw8YXh9iKzU+A8zsoHR+9AUczkLsALd4/aKS5JD
hg+7VG8Vj6pscpCHdnRrR3JiySFolJ4rz1lTTd8jvxrvkSncVhY1eIbQvjsxkI9C
RI0BzqJ/f4NfK56+hSYVHKoAXV1tSaggy+IuTaEU6FEwAAb2RSWxQ3yKMAbkbDYl
Zwt+de+rS7Orayj/vLiV9fcoytMa9Sghwh8OJbTyEnhQH5YFP2pyL745UkpRllEB
R5dOQ50ZY2F1UseEsI122CeZK+R8RNaKvacwpWPnNLZtqPfe0Cq9cwdUvt5X3k9B
kMf5mvmNHLyeI1WawD3TpAW/a7Pwzs2LYmOWVElFiwE+L/o3oHNY7RmDnxeK8T0l
C3htJBvyAOT4Q7Ti7vAJx8kJXRWIYz7AuAENXF2dJDut5dGxbpDfVrmsFGrpaPSG
3sC2FPMS+PEZZbdT9UfQ+878tKRVXcgkojaMPn6+eVAXhGtEXerz3zzF9mwn1jtq
2+6b8hC/1BxxnbEQkPRx+tQrtZfetFMjOAduuE415MLelOO0Sc+0F+LRUp1EhPHU
JZd5yM1n0MmsDeSIPUi7r7oGUDqwibjNX5xCL004jOQUUOMcjb4F+rJN1evPhFP5
Bha/jYTDY9lp2f8jr36odOnJFKmmHvWRli+Rz/uS1fHcnlt1WtrGr5MqJGOTmpMd
bHp658Z2NCeY8oIjgOaXCo3RNl8W2CrGe2wd0YSO7J1gndCWV8XuXGsJyXbe33+V
l/f4jcKjZQz22D1AGfl2kyKfKHYhkJXTh8p8bosKmPEzpuppzHR9V6+rbW+K4BEA
qgNehmpb0Acl6orZWCuBA7zO4ICtkZAei0U2uvsT6I6eMWsww8ZvzqyQH/yPKoVE
/RhcMgLzFAGwDNYQHpuBRIevF+Frul+96uOf2jh0f/Y0tm2OYiCJkQz0vWqDENFh
xkNqpKmEJ5bqJrA/q7gAr6WGzslVzQmFcLTTIXDUkd3xbH+3Zd0eFo7o8BP29rrj
LFK82h39sXqnqksLTu3ZpdecLFCZYwvqOF+YDcV7ZbvWH4jV94FdMaK7TLWEgzjX
o+AAdZnTwvKxSfaz4fcwNVmCQ2AV7cOJb9bCyYYpf5UHDq10opKMnEVUidBQ1vQa
ZCXx1KoSIFuMf0lbGkz6INdBjfrFwl883FpEPqjTIlr/+v8vRfsBFPxTVacfmP82
89uGRgWOFey+M/sPngTk7xbiPatGzk7/ppYLloG2qPIH8OfBszre2QwEMvMJba9G
GBXkBfSrXvf2KbBH/xE2/dvtB6uWge7I1tdjGbmzMp9MPh5N+2N2iHSE3aDvvbCK
fi60dRTXzx3N8s5Ta9S68o/ZBwQB4gQrdkLqf9hI8BC00U4G79fILM0GDcfAxI4j
q1FxfvSHL6EkEZ0Y1hUcZzFdYASVnAPamXbRCnyLfreTav4xMVne3LCG2rKV9HvO
wUUNeiy46RhEUyT9II49wduuLLj+hWBgOGpE3OFkGtqi7K8DxOPwXllFgYk+V/70
YYSNLM84/LdC+yTQbcQeZTWuIFqy7s9xiZBQqUcsZq+yKaneZW0iuqrUV+LHUAjJ
MFu2wZM7XlI+ksdXNf3H5tiIXK9dRDptsroyoOgvZGO9DomDXWVpRfQO2YTfU7dV
ZioEMBbK5XN5w1YfcCdDJKFEmXs+M0t3zEyEao/etZEH6eA1u1DV6Z3TvgR15Qw3
miMevy2G+le5Td2510wfGZd9kj0NQuKhco0IswB6vPS4NcT00eKI7TDPZOHK1tRB
U8OSWXR76HtTuVDDeYZeOSOmeAeN/G9xB7om1f1ptA6iCXsiBk6rru6366/pQkUl
+IhjVzFLogpZp0bOW8rtCrXyxI/Bf2Rm1a1ccMQMzTL/YM2W74xNgPXBcaiePAga
ruu6kdPNaOp6D9pPjoSBqzYN5vAatg8NHljtirJ76wyPUlojtLFiPNfzxf9XmkiW
TH3OVjIEqyYNlJqqKu/Ee+n+AzyMDW1lfdslK0goRMJuPnBNjy10A9vHei/G4o8L
ThUGM2QUss96Wh2QiS8Ja073O8LUFS+hPAG2LLmbEXK3iWwNciiS/3aQArKHM3J3
V4PoIp3a2sikREciCMRfWWBWB6HdmO9zKi/DgQHeays/VWLDK4oInflWJdw7oXF4
An1LSwrmr+m89pLFKtnsJwCf4zjf5eox81lEGMAqDwxlsFojmcET0I1HAH5VcxAt
JW9M+F12liayqDJNx2JbcVreuDzgnMQOuS+Z+cxwYPE7zWhO0mTjvhKt+Hk3jVqH
Ilovow7/hVGpT2lzV88xpP5A4SfCjqdz22+kSgnzaZDaKmIZ0CyDrRqovlI65qA8
rjVj6p8tyfcmm+DvLiSJJPvoZTN6DAK8rv0muEFrA27uYpZ8sjHzgw+Z5Y+nKqba
DwxCoZEztv4cNrqXlFHJHnya+WnfYHBV/UZtW/Qg7qMsiz30PUTw1/ktos/etZRX
UHPf4cfbBbpuC0vlUGEMZLpkA1vb0sEPvkEwd3P6Q0uZVEIfwgi8Wxrk5R0spYY0
qL4P/C1CefQCKMMeo7F9jmS1amY2RMwP5jxqSi7sh7Af/KNrdP02vBEflsEzGtOm
KjkgVl5dKzQrf2jtXiCDk1zNLB9Pj2PA9/8x0NZvcl3IoDZIJ/nxBPdguaZX90hC
PjfTdA5N6hwOtHZmoCASh74vlg34944jWY6RtRrPsPRNPxGsGVu3msg2Qhyzy37s
oJdoCuq8wnonHvM3WvXqnzlxlOlHom/zlUfAg7xbuFvMYif7q6o8YABfOyxrFHEn
69cb73mzIDQS+DmV/gYHpbuYDYbQeUyAwGpsEcNTt9gyrhrzaClWPNKEQHvAfRmn
rxaEt9FPD9R2gEdgKaNQYNyg1eCpu6jg9H18mksg4GFpM411mW2phloBO23yunJS
qaYhtCZi7gpjQ8PFSnSefTF7FGx0afq2Iveez6aqASuf/rwsnXOptXlSwtI72w0S
4XPyCkjjSewWTOl28QY1yPKbTqv+zIZs4Q73PkUeGNvvmM5B7CdQ1GU9bswAN5RP
br28fR7ejYBEEebmEQzJbn6xfZoX8fGZ8pA8GvfqoKN9e921fD6TBe/QZ2Uqh3ba
S7FANVOiPTo7Pr/0smgrZ/ESHI9grcsRBUP9WC7KWqJkVPXCFeEVB76hR7GhmKXu
gwd1XogRl18m5CJFJTn/lOnf0YTFhuGqMMu02jwfURV78shvyIWiGc4isH0ySmSn
ped3bAu/PQJF8ARNl+k4OTOu7MgauryaXXrTAaNP/JeVqeGJ2T3IRLKu2WC2aOul
8uPu4NdUT4Os7R4gJzXqmU27r7KFaMhoEg918ggnaq2UNkKtT7JyvsfkwndNpdxn
wX7mHFwnc1n2U/SvYC52DJX83n3+C0zHJ2gag9zYsIHEaOvAOGgdZItLrlOr/bpC
ORQ+0igxGtcZ2AdawlA1kMyzHyGRWkJQ0oqAMkpWO6BpvtjWd9HiCMGTvq+kyXCb
AMGh2/k2k1ZSPOPgC3xu1ZpkWLQBTsBJQcEGlLeUsKrUTujJGsZznKJmtoTxqrwZ
zisLGkHUX8wvuUWTOqY34nG3/BLfL0D8512nz2UVZfUcr0SRKpnB7oWVnJozbVGm
/1dI87tlYQN/yMaJTOO1WYexzy/t/J8NSMHKKIDe4ua2iHaQMU9srszVWfdovKeg
Y0dh7aFgHpDG9JW3EQnvDU5xjfhp38986xVeFiYeoH7vyETShi7tj/yioGAbs1CY
w2CW1f0SiakOMWybJX5B4jbMMmtKRWKqbqvO1rfihxTpMztewFsqg/OvoTJlxxl/
3A+3npE/OLT3nfwOEdn+U88ylSbO2wYLhiGARz7b6ZGc66K/SSExMGKawK3RzpZt
e0o/f/g1KLw4YoKnBoKDPQxh2gP9X9ouyL6ku3AJsx3UckOEHsYPQj7Cn/UkyYVe
fdGhElJfvNyxMoVhZFlr4FrvSrqx1ENLsaBILo5P752wjnjl9+NpeDlh9gLzIIr9
6t4K6p4wUsyHh3pPaiPfslZvG2U9Ayrbj/dTQlXg9ftvBKkxIDJrDY+kekjNd0Di
vgSbqHvWify4bO7sRDCPGhfLHyMyy3ceEje9AdrvIzZd5Io9GtumpunRMIDYApOY
mLEwHPrBzqJgEzTSKxw2EJXR0whMQAGthiKb4tSjzekkL8W040bQFS77VJLpd0+y
2MHM9BWA8NeFbpjDvfOR99XlaYyq3syzE/cRqD+6Jon1IpI6aRtYJo71yPgUdavN
jB2ijvXEA9PpzEt7pieat/V51fKwDiyEqh43WEND8jD3zURsy/8UPsRFxm5E81WK
3chfuPJ1M7wMt2kAHwcHg4ayXSQbTKKYH/mRJrJ+A/hZJ0WpPG8kRlJInPNB6CWf
T+5TSBtYd1ktLb3iz2r00LKvuLhw6IGK0m1IKgs5ea0JeEV3MxnKnVjs3TgZm7tM
xcHgqjMTiAGrHGdYuB3Vu7zzhzPrgjkFelx01suU9kW2o8pbEprWRcKpRgoysLht
KzIFlXg4/kSGtdq269wKAGr7GlNaOv1zkrVkpR4Xicy0CPIdXrCjQdgiTZFJ77le
86LpxLhqsyJaVC5KWi+JtSoKEgmWYFT0e9UOJpDsP3FVueFanu1x0t6GNuiRk8vy
DZTCHw2lQL9a/FrtWn/K9ODn5XnnbbetzcgDhZcIefzsa5f0GcUkWrOSt5D3pMo1
Rnnm/Z+znWjs4NNNQHrf9Tt0sxTnVB22cENqEFz5ubGhxSLP8MztTDc7n7aIlcQA
yHiKvEwRIObIoYTVmPiADZEa0vOKDy37Eoxv6dX+7O0fr1SUgO8Le17fX3/ILOAI
hGfSGkL3v8ZRiGqemiL8cGwRQYBEGlCYF1CSDnUJABFml/5R3ndm5aWUrrYC9jMj
bn1Or6VpdecYh6+cEZwLd0xvtGkgG7674/4h+pL6KWDEqmGIbP8JdLv1FlBTOFgX
NYMXf1Lnk1Kqer4MlJpJuL09XciegCdST2XvBRlj9DIeI5YpO1As5zztBkSCb+Wd
G6B3jTr7odGFjvrLY4z2LcU458Jmq3a0sgPUFd/7SZ9/4Nm4iQma2kCNQ41FZd0n
XbD8Qmlkrbddyu4yGVrfQ3D78jStGlRYKwL74baA9Q/8yAuCE0WtcRW0q44p5sze
SI8nDFaLcxpvtMlXsiiywMXZ02OdC/+yyrce0+/IkJPEbh7tWBpV+8ew86jiuYHB
X6iAHyrWw3l881h+8/CyjNfMgPsJdo5zpDXjhAW52sa5buqzRBaVaJrUEb+ijh+j
Zi95YMZOTv7lCy9o3/X11T4mfgyiAV0dT1Xeb87IHCXr4Bz+8qdDDKWp7KQoMcgv
zxKIJJhe4w6dVgbQZT5XY579TfTdfGknMlKe1YsbJT1hrDTddRvxtp4SAKe5aSF7
rQ+RBINwoVhOOusWLpywslofyxVM6dNaUHt8aVVMl7KRnVToh0ZO9MNfL2BL9htn
zYINWgYDXLqb26DRPAZiad+CPM5SCEwAVUX+J4tUkrHhIUT8YxPsa/GfOPreBWIw
VqX4w/i13Q1P5mnyp+QUVNQt7TgJ2aHePoNGan19tt+XPnuEgr3IJucA1Rkkm0JT
rHJGT2UDqPMTi0L70aZp+YJGwa8E40A+fozpPIaedjXcBMq+Y69XbDum6tp2rp8V
8dHogaLxttDYIFsHqAyfuM0BXqtwhFiIbTJqj5/gvGJeoFnOxz4tGqwFNoqPg0so
aXAvTsWHjTG5fakxIggak1mQZIKgNJT80KANjQH5PXru3ipqj77xjlKNVP7AvB+6
N7x+cdNAfbphdh+L6/FqHzgIxfRb/Js5iXdvprPcRH7QMspBpsIlTOKOPe1VLVnh
2fypDbkkgHXLj72x2UnaOrXTbj4w2HGzaA95CvTqyPoR2C99MDacTE6naoD1yIGt
/3aIjbTNI9LBopHW5W7rjehuiOSBkMAUMbfvv6XvM6yv0ClUDzItfS0eCdY0ka8y
MP3Hxv4IZnLWUGS71yN6TvpzBHkjK7Er3Lv5zIXqoJAVcyQ8ScnKRaKwkLx3/szu
rzyvEM6RSSwEVCekxWR8OP4SAjSXBprc3Q+NXYNaqfiVXm19sezcYUwlAWOUp6s7
r/2AVb+ccbBsfo6cqiYLw6tOHJ+eW4YGxnG9yGwAnyAhPpEMZsEBnJ50FN+5Lw+a
phIKLV3nEFc0e4jYkCwzpnWzMlu50PRljedsD4+ORd0pnfjT+8/KfTW/vwGdkSoY
oPVM5Wv0PaOE8LVIRBTHrv9lR83UraguCETdMbzPv8daj7jC0XzheK4U7YL7tlV6
jepF6mxIyvtuXTsS29x5SuwaSp0kYk5d8nElhkooNKBdwIDTHnkhpU708MBexNU7
LfKhIOzeGB1BSi1TDSHP9iIEr/Z3NsWfenboLHLaUlhI8oNx/7RvUVDVwIxMz3gZ
GUE6TParB/Y7cAxY5Ml+hfR+tT1o1t90yf6lkoKgwArpAE3hHDDCtRUPlq47g6Li
Uu4m7yqvIv+M43Hu0Nj8GeX/TOP82qIrOYKJqJfQ8epNbH3oTuR/U6f2nX+ym6Kz
13/gLbZr7v4gXltncOE7Xk4j2JEIEYd4jB/VLIQB0FHKL8jIHRHvYAn9evz10msn
f8VROhAlG0dvfcC61lE4wf7jY8lr8RhOFXNr/Z5S+ofvFxZW9afJscrBu/OqJSwN
Apldsf8gW8jv9EfFXO6KTaBXULyzcljInBcTMBQ/1bPu+Qc43bOxAWwAVBqt0Adk
qdMTQ1yn03iiUoZwSnsXBKgMnkfJe6bqQsTM0tmEtKtDkrKadNSbZZisFN0UBsTU
9fqt+2NaTKKOEqHYeMO2tnhjJoTkM3Nb6dZ4262OGNDGE+mXxHbjmmftAwLXwRG7
EULQGkgWDRqpKB1244UGmZAiKhC7Q51BVoVHqUsqSmp4KjzYtmey9VzOPLUAaKF+
NVgqglfgIm589snxoHE3h6z/iQsAuk2Qd9RLRRCmyI4qqH0bu5aOb37q64UDOCAL
dmqvgFjDNQUFI49k2QI4CoSiDEi6QnWjhI4v9wfbjhOlKgGI/panecXlXEUP+ttP
1U79r1QPtjbceelyEhMiYM86k9WXwWDkSwYyre4gy0bgBA2hyHXUHcuKzjazHvdG
5SGZT761zCQA0E/8ivF0VY4iO3H/+gD+7P2h6SNd6ykgdpx9px7bS1uHkcZPkzXE
v04nbjpGXP5Ct5ay+ksvACe5E03Q0jecmaMx4lZUbj6UZwRO0QnAiUGnFI5w7yel
LnbA1eY69TB2hN0j/5ZArxy60nPEdRh04wPCa/727LqCgdrpeyP9KQsRUYWWEkPN
Fqio69iqQ1icDEkQPOas5U3xYJUp3mQeEZ7Id3lkBpcB1VtK0n8lD+4jWeMu5O/m
HJeJa5wtBz7113PPxG/x/VewKJrVJw1St1H8+3WrKM4PskxRiWikDsZl31J7uI4l
5O0Tl6xdxqO7FKMkiV7ksNNvbyxh2hu587aTLlGSXu9MEIKCeixHbFVWbiP80VKG
iMc/UaVWyibN9+5B2o+FYWVdbhPs7ziDIjN34C6cGKWet1tg/Z/m5R0NLmFB9tmY
c9m7xnRKNKZDz6v3QlJetot20jywtiHkfXnhiWwYua4mySUT/iInUX9gBku1lRI3
yRLgs+4fD+Jn1Ti6BrjQvJJ/8mE/Bk+uryMq1rbnmNLPKSy6tyOtfb5PbAeWtmM6
45UT6FpFF57LWo6nKOyFsZNQ+i/Nkx4QQSbq7qcBNAwMvTniUp129pkqnreKmB1P
/LNBEm366ZiZHN8pUp2p0gpyxMpRbL3OM0egPQVtLzoJqlVkL8sxz/VfYoe3fYz0
YTHPt2cNya5YpXb6aJUXvYv8myyTiSDRwGUpUzJAsUpTQji9fbLugDW3GppN9d5e
USiGxBL5UNUnXAQAJQsuRJut10DsyHILwwrv1b3wFiMISQYOHZzgix0oUL5Elugy
SVr0sALYwka5fL/VR5EIlpbKAdvsBCmy/ZBFRwsspv3u+MGgrqQgzZEqu8/Mz/aw
efzm6GevMK++F6sDPuW4Dh66RLv4pmuLei0/f+cIgo9HdKsVhWDt5A1tS80qJlOJ
BD2s984WanHS9O4/a2TozLlFXX87JlwptDjU5Nat898LxUKMXZQRv/hxvEJk+6Hu
r7poFghWGkVKT1IMJFNFisYMEo1bF+ZQSPkeT+YaWlDRzw4/0fPMqLRm8PZjbnK9
Dt4UVY5nD8PwbJ5hpXMxWq9twcB+/romj6gRkaG0BGFpOc1L90I+EJnQ/VMXNyaL
jPcEtoAeaGKkn7b2Gx/g0Q2O2ANw1vWblkgh+R/UGbwRlVG8zCZoQZhsnQuUwf8B
J3T7uDoPsnzEn5LD/v+3JO0IFipKAoErQ5dnleI/55M91gt4Y80fKg+fVxtB1Kfv
o8hzcQnQF1jIKir1dE0dqYlMRMDAy7KFU3foMkiPVmWdcMf5FueQb7KC7AJC2d1K
JCUogwO5QeL5nReN7haN7S0qSNGV83b2n7CQF0U7JDf6ja6QWJXZicbZIW5+N82c
pq/QkpPat/5HuqNuZaPA3r9MWNGQ9h+hvwCefo+ND1QDdBenyevg+uDIPI4TRuME
M5htgQKsP3JJ6EE9a9/ddHUIkFY8MYCBtjCM5qOhXtqmVUEJJd/vLvnuZL0mKUNG
nvAmFxUxlHSya9N3h958ECY9xcmMsd+43lnQVoktQCrKOQ8GTm0QYGmmUaY1ShEK
ZVli1evWEEzR1I/6bMN6h0ubJqLaCn3HO98u01AqlkZRcfkmUdIzqJxOyuiDXnDV
PX3pdkbzrMoonRLKieWUkKwBLppWMcdZw5zcCns6NGoxh4ZFUPfyKVouMkwpCW0R
QdE4XrTRBbQZwelH7vbkhnDuXnwPPrG/iXzyBVB+H7zZFtEQw9ThRBBHUFX35585
A2ctbxYVulfkBLMF1u4U32ZcM0LHgWol4LH8LaCuELgod/qzbkMeQiu91Mm1Tfsk
owQZVLANtlZSTYhN+pzXyX1MM36KFhI8EF6++ccjV4wXlIDszvF79SxEsJJZlyyi
pyha90F1jzWAwpU7UAVKznBglEwt7XGR1URgVCDXwCfDWx0y/Jvf6LAGb8JrFQ9A
K/yLT/0N+nfifxIIrGGaM6/EiJE85HPzN5M4xKwphoqcXFeMygc7SMq0wi3gfWjX
isbcPkYgjscfmsIPcVybsmbZn5NReThKCg7mnP8QDb9TL2YAM3r6RCdLHJHZdnSC
nIF/zDN/cHmDgnrwMnVyqboHicANo1lS47/5PME/ocf4Rq7sKCJzlZJsakgOx55D
/RHUSKFuLsTlDN75Wd0/+gp7NVzz5A6EYRBFebr7DntyyJ3J3bYhLJ/vy5GBnrfs
6ocmY16EihVjruGrJmaO6Zu4AJLgoUE4bEjcOMaOZ+h8S7tnSyV//awT0OF+uTrg
xMjFyTErGxVEmIHAPKn4Ejcoi6RRGRkkJ/xDZkgD5uKT+tdUbuflpwHq/vAWGvmo
IJVYMhSIiRahrSTlRDnOxpczk6UwlLYj31FAkUbeWGykZJ9xZEpCTb6V1OxK95zj
mhBwSyatkT0dGK5P9i1+6PZB+OUoTbDuEo7DEJSm3Q47IStN6ceUnMA3JrkGKYg4
LGMiY8Rm3P1Nhu+l7vQm9DZ1mRkpsXjFSGj+KDVNxur5Bb/ijDO9jVOHDE7zvnsq
Siz37saktBNrHuPofW8bF9mzqUDMyTGbHjW7EgO31sh6Pf/5Ccc5f9QIzCRpRiQO
3kyxEqsQMdlRL8DcoN4pJqWl8BdwmRNa9jxYV2YcqZjEKWBmv20oRyZPe/XFbtDn
X5XpXZODo7YauMA44wefqjbPn95cf1178bHEoT5MKl8hWKiK/uUtai5DCLwOzZUU
z970gKfNGm4KXP0KQIl9NTEedN9AOZhWZy7nyhTuOgGfIBAvJigDHOwHf2Mcv8sj
vdYCjGtLcBBBPh9NHq/DueOdcJ6jv5UBdMTyQvyl852Ro8Aj3aLDBUyy4Tl0V4xm
7HCBI53bp7TpfnsQgh8RTOPIvdACc7WTTxA+4UE/9OaZxU8ixwpDryEnVsdXb7EZ
AsG1XFb1jUa2MClfSQusr6Ptq8BKrJ3K2hgS82inXo4EIur6Lg54kyGuhpeH1rIE
su2ae2yzmPYG39+hAFWQJSBsLlDF20VLTMHrMoB2D3H9LHubKVO8kt8nB+2v3z0g
yqNeYcUDwJ7LNs9fHaU83p8DLiL+NTjJ2K87ahHSi3DbLxLhNJk0d6rn3KcatuAM
ZwHbdOGXg5yBHNjKCYMq/HZvmbsDQ2V86LR48WthXLZQPDw8rR8xTKLLSjUgqzt+
/PSWLbckYivNmTCJpO3C/CaPFjx6Q1VHVHsFYW2GwDUci4SURF0lSYQtrNdPOZ+Q
LZ4M5TKK/7520+VLHHQ+F4ITpkuH57TomwhS8BXCc5+2C8V3THorGptBMAtbfxxR
cGblo+ZvqqzR9clsqXbY/5ICKM+BvkqZ79fymwLfIvIkiBYriMw8X68Dp5oSd4v1
2oydzasoVw+fntBfpAMa7HFAqqn3IO2TCHuGGNL5+6/n+lKfla2HCsIXlYtHoS34
+TrDE6UFuSmweQGDHyjVMaw+8sT1jBXVVTHDKHttbTbSPyjkIskKwKjEpwOMLbx/
eANU7yjDIg4Cql0rJk4Or5TMs5TuCa3pLUuB4JitVxdQ2KUuV15Jp5XwS+MHnZb3
FwiQCsbwWYQCdTM1yEt81k3TuGMXnr4+yx+Lz/TnXGYEqdv9JbTa2SSkGOXtuBSr
qznc53R8s6TCvj9aS/+zQ8Y/IyG5QWFXGSrDTAHl4O3lmn2q3v1obkrWbyF1iQvV
jYb/GTduDq4ZV7RaamvA9OvtAicfE2qVE0YrkSBdi+IJHMaxPjyUcNyG+7jWIuZg
kxJhq05JUHaG68o3kLQnZsQMOrkSYpX7EDMTj8H8QZ8s3qmaBidPJ6CzM6s/lpIp
XMIwuo1Q0tUaZTxUj/dtc59qMNAkHOx7gEUKWe9IlKsDXswtUJFAW3b2hgrSlq5M
hjQtCVCw7j/0Apkojbz9l1v1xxnxb9HHARH3lM4+x4QhisE+nBhvDrRE8BI1uYAt
Fwo1R+JUYmpCY7nNsa7OxwnuQwjBkmDqCeidG+e24eVvrHbXRx+4ul03ViTD2Bn0
fVFf8tYwWgV5NprspnNBle27VVEeHqxr0Zbo03MIEWCONzcfwiPZ+LYjMtatLa91
LL3NLoycm5ZBh9gTfWgtV5lAL+uzp5rL9g5BGAboiJ8sU+kgpp1vhz7PfZGiSpOx
wTYqCT+MG3XJsMfsfoyJaKOPNNyxmFUKgK6c4OUy6XqI3QGDAQdGo6KoED4S1qIp
wN+r8WsSYvwSPhep5yQ569iB1HiX+RREjg2d1ZsmymLGcgybu89KBVURX9QqiYhb
0OjM3fyoFfp2U4VsEXlrv5wP4mpw5X5pIquR4ekRVgOE58sjzurExmrH8CfXUEoa
PyYi6iQ/12pOZcvMMDRBLQUH74uC/fH5ZmeoAB3mAMUC6aBRZIVnfSiUlCewQ4dw
gMbul47/bO6dd9VflTk7uZ1op+OFQaIhSkZeybnQj0Mr5DIQs1WYDXnbpDLcnkNM
vWhoJt1uY7JskHdcBN5532IYlGI3xbix9//FY4orleMc3AvmkLXbjg7vK2EP7Abz
hydDFC8zvvkaZHSM6VumRP3YN6o9YWmrmMVylaiVr1UrIk6Pk382Zfn0tJNqwNwh
tPMY2okGvHZAHaS19V9f+mvWvSk8dKjLO6DLD4AiuSschX7SyV4s90cCpp6WjJyu
HwguY1hqKyIkqt/zF4J2AO4aJjRSI05X3jnSXrM5jbGFmRCbngEp8Pidiu/MtVgP
eaHSilGhBsTukZQOS0l41EZTqpL1LLcndoeUlb8cpB1A3rEbckq2fWf0l/VN+K78
vJAhCEDrsIKpUkCGoShaE2FXHXxGuXfZWItBojnB9cSUekrkXvsGLLsqFG9IIDPw
OK2hHo86qeBTaxem1V+3xG56nOXxpmchg3zBoPl4j4fFebnYbYBWAjx+Y8bSP9X1
oG01tFFVsSAUhK2yr+leQyINswcfYFInj9Z/yKmQFK8b+/1oG/VNK6Qs5Axmqb7C
RdAdCaJ1ym2bpmMdleQGp02o45GAzA25SqV6DktcAS8cFhOWt7tOb/tXQgEGHPQB
JAbEIFIZgHo9+w9qMyLXxUaHYz9zgp1LH2aVJ1IOJL7McFv5bUimzGQxOEmBpYqd
MB6zC9paT30X01F151moALyMpdFn5hPduL18Bt6FqmAWiupUPfvX20AaT5pX5wJG
jzlff1K02R4IXv9WdLgyZ+GOQxWSV4+qTqmPlzfQ+hDhQzm+xwqAbZ05/xFLRnGR
jJlpMC0pFEPMPUQYV5hOHZ/bnW1gut9jBS0aviOITSiU2BWqcgZHNt1l20t9fwpP
Zti0qkaXfDvYv3oTOXXhcCR3xuc0Q9dSf/5ymg1dFDuwePXnyF1WLPWVmIF8l+PZ
WXLv7pZYo3r1evh2KZlVzyGJCK+ZpIgoTCSZdKqOMf+LBU0zqlwurcayVNpgCOpO
85QrhPF01kkkkDy2L/+3c3uGcZsHKqRONHFMHnyuvhyQ3/w7Ym/JDbuEyvVBlArg
/qapmhDemTu3uU8ftvlEiSDXHyr+zBzMw51UI9GJQLhcVWVe1nvZIU7IWDCIYOXu
22AoeKzxObqU9jFeDkga2iTg5NK5BI5Z/l0CyXv58MNAxB3ziixyo07/yikIP4Bm
Ff3BAFMGRr5T04rfUm/D33ryMZjzSdSemf9QeNnnK4a1Lsawd5Orlgxk63nhj0az
L2PDjBzwvY71LMcGyXdp3LIHDiLPpCSsHmBYUaaYeMSYPvjhm9jDkFPmhtz6m4gd
qm6GEAyTAivnjF3gB6obINs6a5P8Ini7NSZzyLl6doFTBoKwpStKIsY7r/XQs1Oq
FiPyMIkYz2FdHmynyf4OyUUJ7V4YJAUKmKEC8WgU1OGOu579Y8Z5F6QlGE4mtSOn
KkPkPz3qFpE0GfGcN84Y1s3EQGp2VnRI2ojGMlwwMPYv7LMcbL0+qUuqavGoXmmE
0mI+NUN1n7EgQ2hdLzkozJTRiV5HHbvPVfzuPY6Zp0J1XYPg62f4sH72GNm40NMs
KKqXn84sG0/1fIYh5MMNzFTqO3xE4NFq7SoeiGgOL1K7tPUp/hkaBnYPzEHzuie+
opxeNrN3+BDEZHngDP1mqq1+PfU7eJaE4824EzTC4ZTnQJEDmImVjf+2Fepb6Y+2
YoxIbl41/g7qrjuzcCqKPsKJBd//r0shHHhojzH2pmtQpd2Vt9dj5/xwev4j1ts5
iZn2QiCgaqkIAUIFueLnyZj9yzM5AgHrFEc9h2BMO16gcmoEUG3g9COI8gcGxWZS
WkwyMzBd77Jy8C5JSNCDyrUopiJ/Au7onuoG9m0YRyg43/C4/mEJCGGUainWmkWY
9uBvN7JjmqwiO9pXrPqzvkTsIL4idq1J2/XcBcXAtiuTNdPhkttO4xTe/td4MG/X
DNIXz8dH4R900Adkv+hIXIT3R4WTlAYvAe47ZsfHn+wkHtOiz1IVShAePeIMQE3a
EGv1wNGNR6YzupFiv8/rk0ilx8a/UgRscP3VIfTKFTz8jnk9f8qQrBsr2xjTjMJt
h8J26P+63M+r0mCYB544AGZ+TUHFwd4VMTaK2dNOHaEXHFktCm/CDvSm/dUzpdRm
BE+H/lQXnAm9CdA++TDnDnehdhzamOxRhZyniWhij0rbsytdS1jseSsixcWQjNTn
vfgTml1uP2Bc/ss7uZCGY3pNaLxjhuosyVhPuois6RsbuFopoStWReO5QtPSNM+T
ck/Ca3mCIMhcGXB9f1dyxkZ+isHkQ10hbISho1lo0XjOFpHF9NktPZ6Iz9dV66wV
NU4vxsx12jPjAjG1CU387jB9n++pYwdzu9Ny75JHn5ByMf23AvveRg6UL1kveRrs
uIn8bTe5hslq7MWURU1V+7yOKuxWGmtc6P/wLDRaRlYj3u3zqzXuzdy8doINDeHS
Yv+4IUVRd94dd/v0E1wBhCwkdZ+ltS7B9eb3P6tTY9hOGfm8kttWrDVd3gKmp9f+
v9cOAlX6TlD0zF0Q7Hmmyvn2AnqxIP82pFLEvomVdROa3Nnq6NCgNAgwM8f40OuD
xgO991Tb0gs1fjDX9E+kCGAxk5RbLbrBTPv0Kiqtv/rAa4azJAYUkdW995zjscah
lRo0ceLipiirPsIFBS1x6n4P2kqTrJDY30iOyvej+Hp1FpxwQ4HrJp87Gu2PKRYH
OZdhJy8QNmk/JHw96C+Uo+Wonf9q10oOD8SG+bTf5UR2ZqVIvM8ev0cgCKG6xCei
Thq0MPTYqu1Oc/8OmCopSRH0m2SqYCCoivFWAkw1cCpQ11ZcVYXeh6dyU73+Rcdb
kiQZgr4ij7dGzJJoFVZo5Kjq3SDHcdlRs6gGcpnv3Jbgu8abr4q8G20IWqKSzILm
Ysj6244vTxLbelXTDHCH8A2YQm74X/h9E56SxkOi03IChiJ43GKed/BdAfuKISuJ
aVrfs9AXz2EABQeujlgU4X/DrbzSYsIMueFPpJ9laF2b34ZZUnBx0NA8xM8BmdjC
di5pSp+5tNcy8yucAbAN0h3G+tkwX4ItlB6fS++3WiXDomyH5yiGCTYGPkgkTpMU
mePC6UCSbnYVLaQ/EuNC80GzjsN9f74bTWGdHTnog6f7VvDVAito4q93BispvBtu
LaZWUknqmlW9iyv+6mNlByAHNPPdfsNspaahqO/hhoQaKxDG4nn9nQfSVoX9zXFb
Yw0RYnkS3yeNzd7Za9hVDmpxZDeEWK1RISBPKf4eWXSw2jlnoOwRQpSqU0DZ8UX+
Yfh51jrE/htCFCp+hNGShFfwtYfWV0pqIi7SdNPopjt8OmgETI+nwHbZrtRStOkW
p4vAtJUAZpF66CDPZbN/FIxQdP4gtAhkxB50V6LZMmrECw6dC7Olnreb1uRfPOHf
rtIXteuwRvs0GDMD/0Lqe/Y/19VZwPlCgF0SWVwTzkhlkagH0XFFKw3dORGqpuyU
KcgLVZg2Xv5zTyaICkfmh1ECc7P3GFXCjzqhvVxfadONp0nECXB2TUa4/L9xuk9M
ZrQaNqWm/pwNepZscyM1wiV6kLerJe7KohNieb2b5ZRWQaAuUAYSSEQiM97Dp/3D
w2hEoXPUQRq+8MyxPgnnov+wLUFZznbm/ylZJuUwDKF0zOcVjxtQlaGhCCplDX2G
UNnunQDt6MHD9XOstWb/7/GkztQjItRmCP0QUZn287/VpiGsz0kXJsspYVuN0Xi8
8jTp/ZSAu3CA1img58mlAwgraMS4AAdM2TYmsPupL/7NuZYZt+dtHRoHWS8Iokkf
zx4BUPH184CMqOJbbj1jWh6UBgYyak2YZhiEFf+EzSymrc/3FdYSIO/rds/yiSWU
ghzYZKNUMZLpTbwvsvXKj7a9nmkb/jtj+pCBZsnFkfPnVmzcyTQ71WEVmooeBEHQ
ibS9ffhJlWv0e7M4Doz+8/eVR0dSGoQ8V0R2teO3HrdaxzlddUCHFqjY9jtZlOG9
c2nOIi0z0FwEUHIZa22PRJhIlKKdsFi5t8uTfaM9TMQ+pY9cwvKXCI51naX7Yomm
UhXJe2Jkxs9O464EAd7MF+f34eFx9z8o4E7RjHI8wmqBvIjVMa/ddLfj0AhHqc4N
9b09ZHlVfE8swIyHIVejVg5LUnD1jz4B/e3HwhQYbJ0jAqitoau/SSDeri9QKck/
4gGeZRLPUMJV9LI1owmjerubABraH20oovQ4wvnQOOlBMeDxif9CQhEEOmQWfmZT
olUl8yr7GIYz3quZm8r//ckFpiaVCNcMwvLCUHD4fD6N2Cvy4ij25ywWsO/EJMkY
niqw12yEUEBfdny5BKgFlJfSPNuUu11DZe6XkB8FOjW8k7Pw8/6Y3ayc6Q7u/w3j
tb7auFpJutudqOQBN0stYSljav7FN9tWvFUlrZhURJEReeIahQmWvd1AUkTiqQ7w
8BHImAIoAFYFUu3NqNdE3Wh/XwiaKOvJSsLeaKjz/bUyZUtekLKHndil4wwyBmec
MInZ/i+UtXPkcTrqhYY+mcP5b21zV3Ci04vXSg8LpQgNCjVv+FFkXl/vTCHP5U8S
H7uXg9joylRVhSvwNUvfwCcxgLGiWuyiTWgT6kxaSlNh5Kypi5oUV0BiZuxrTl0j
wpt3bQlGz8HSYxhpyVwb9d6suyk6eTNo5sbVFh+nb9TF2maFC4glnKTtSi2IiuPC
Xe5quUkZ6GWbpASi99Rk1egngeIf9BivsV3Kt3f6N5Ne3CY0/cMhMewAp+CwY8C8
oFhi/8mEXv4DZxlAc8lpMa6MW+D7yJ/RFQ6tjgFjT59rMNZR9oJ+eQaghQcgR7ou
WrE4pQkcUfdZAVmLRM8hy4KH/rVjIWpAZ6BwImaBfpxqKX7vjI2EEf08Ie4Xlynt
oSKs6OF/fEnr/7HISYFdy3u6NF4HMkSPag+FOV7Wqy9Bh+V7z7M4ncVwmy+jzFBf
Sx798Q/HbKM61IIOBK54YWzYIKxkOba6p8542118XbHCa7A+30fK9J5s6glZ8qTH
SnvAZtc25hlucniY7qUC3LOFBArBR7vjaPSJhiMUU9ezNEq29NR8XGDPPN9xOCgn
zeUYh1paivedS0MASX+JPyQCq2RGS3bnTHeOqxpJKU1pWZK48nqSbGj+VWhMt0Rm
jJCCveppixeiObBaZEUarY5GvVG8wQytWZRib1z/1KjdKMqcpoxMGrG85Xz3WIPf
2KJnLv9J00v3EJXy5mAr1t2J21yGhgui7yjUEhMpZHyUEfWklcLFgDdtbyVEB957
rbO1mkdyw+NkEc+pqLBdX7YLlIc+IX0++Rn8dVuwNTPWOrmXR/UzO9EssXXx+cvD
ZYa8SSLOYG9KjNDABpIHDRInavWoNbdcsmh6IPyF518M7aQweVW3QGoEDDI2TVTF
CKE+tWO/QEU0LgB3W8qt4Nyn9DPZj7A9laXuUUbEuvivFmhqtzH2xU25I9GBQak9
7pQ5XMGOISYOLyZQ8Yqn/HxRT7sqZ0+zge7vd1OuOgFC+njMtwVKXMDJtKuD7/hp
6ncd3yucZJGs4WIm16fAdFiT+VwxGMuJVlO1jkIWuDcdc2/b4U8pVsr1OrxHfFvb
s51JQx7TGRU7+qiOA9Wlbf++D3C0GXamRSyXVVoWWSMWHEu6B6+5n4dLI1I14Frs
m8uF0koDUcXWdNjg0CU28khmQQaQ76CbSvNvfi791mw2U/22YYoyoC/CH/JpbyCl
Pr1H/nJy1nbOGSduMLxQpp/opEwD2eaaURoK9U7wOTEkf5PrWd68JzFCBKy36Ltl
qPBEFQcvol4odFNamzaPJtuGRe8l0Vg8XwCtuP8etAFOUalzi13Vkh1TM4/t88e5
n3nPTt16qBjabfWW27hxFZMw5LcKY9GAGVq6P9BNBLFUf1ApEJy5LO1/xcotU3ly
M3iJ0oSvPhyJD2qSKDdk9gSwecjhf/gNj6fYeGit9LdY2JomK3ECP1Nav55nmWTS
cJDfhFkcFfGWx4WrJ/GEKAz7Ow8DL7x4nAewJfB2FP7OyEUcnKMun0doGDz0pDIs
QOgkh2p8OL7pT9PJKBi5TD8We1bZOoLkZ5Js/d2h7hvNbdJ6Vs3LGNHO5LEdW+26
JZVF0qJJ5obgDn10zWq5yrsA9vrYg/pShHx2xi99mAGCTbXr1E7nJiPGhaYmCryJ
c9upc9XGzdqmif3yJoIDdAHrA56lZtbcF5vm/PL3tl80GvQOi0bvkaYhbHQTbF/Q
1im03ycW7aQNy4G9p1hoNgqo0ZGYKJVedhZG4683NPj3bPrSwZtXONu5o0DhxMeB
KlmWoT+dm3LuPA1pf+j+9W3cYOpPkftLfldXAoAAzkn84d1Az+/mUnfAX3NZqquC
vUFyjUS5fP0DJM1lsft70dHXUahzVhfoN20s4McA5IPWMfXudCPyi+MmEQts452b
plTLqpaCB0DS+Ghv+z/d0HDxxT/VMPj9+91MfCS9H3UTwa5LrTyywWYmouKcR66G
QFgmh906JG3MHCq+X8XLbbOhWnBARRVl2J7aiGy7fPuy8EZB2Cpq5DDQKH5FmlWD
C+M+z+0+lZ8pewUk/EIDkG+SnHBgNJgJ+dhl8rHZeL0PYEZcQTArOZupIP7qgHFw
lhXisfxFJayNd1mc0wObskxdYeWI3qsq4+Ro6EvrHseRkNuDdn0NJbthpkF7SQ9y
FRY13D4GcQM+TXA2fgXJUWAyGpZaNRsMzwdP9TYj9I5eIAO40m37tfR9VPzpiIP4
Q5mRo8H0jrcB1GL3+MBpaWyDkjnWD4I+hRkfHl2NZSYttqVj74uPZfe1rmkUv83P
I9C7uBbEYcuy8OnDW6WS4Kbp3rUe8OrFdY0tR80uMSmHie4vlAPc2Oy6uEdlkhuV
j2m9dxE51VLWwEAuY3HpO6M559e307LMMIIubbrFYzzNamqtqy+zAp/qd9/1giOV
VrAn5iLZ3Qnr9+LkutRuR+EmY+pXyYiawCcEdDzglbuJ0iawudNX6dPGGEkKxQ6R
WcRxIukUHxl5ZZQIFBuo8zzQTRIHVdnnqi9/4haUryejfmAZfyfm0vzA1+3CjHR0
O9tDQvd5ETUZYHGSDutwiuIBMiCmBm3YVfM9PfyCJJ3K+49zsw/OUkCMWvAgU6dX
JdtgfhVioS7eJ+Y1b2DuLMoL9sfHcHOVhGVUxsIs+cY+znFd2m8+Cfe3fCBTym62
P50OljfaNRpOgjPDy23xKcS+RClP9tIcf+HR9HH+y8cnde1+A6GqFfP1KUOWzOF7
/3ILIrsMt0RttMuutgCfx5pVixBYqK7+mKixSS04JrtjUfeu0641imNvJKKUe6vH
pKXnbrd8HmWtSFasxwQjiR3BVWvhs04zLlrMbNASOviJ22Og3RLukRUf5+/7+Zr9
iOYIlk8PsYF1UivJ/h6w0qHbeI4znZw7MWjOp8lJfkoG9ni1rI23+qLiI4CO/JNJ
+K3BwptFkOptk2VlUB5fdEtdL+9ooEn20ySJGuCecCYd14LG6NU2PwjU+34Bu9pz
w0pEozet1za4JJJsxvSRrKMj94lUS7NmfyAP9v/A0B4xy9OoHjZG0BRQPplq42qY
K7Rzz8lZfgXX7aJLPI2pnUqNTqrbJfrLUUTSV3MQHIHOIGrh2AA7dZH4TQqIj+qg
9n/iht4FdseKFCKkodHKt9TAZiu3qKjFSvjqnL42Aey/nDDKUbRNOXUe01jGEfI8
poRKNq7mum4zIOX5uTecyEnTAjManX74vZJA7MNYjc9LWuaXAfOrgmKmYQxJEgXZ
Zg1HKvOKatRoz6b+q2WvinZjJrsrIDM2oQ6frOetq3ohDMvdcP1OSLL6j7byO2Jk
kSGktbbviWS+pM1eHhCZ1SDwKsGJlwfeEbhuwpg0QPPsGvOVObGbyHGGS/qiy+OU
SBAncfRDk2ZrtX748XMrBUBwng3lxnsw3QaGWw+OrS8MKTdGewA4f2dHOSgoHecY
+QV2typndhiPyuErUt77HHSKJM718kW5b2MKj0bwIC8gcWOTMywga7TLracMNvPg
8CC78G7mJSBUvKWGLQzkyxssVKly0bwd1xh6Osz7l+nAARIDcsHY72GQBpI1Voxu
2W97/cQoWcLXfO9fcYaygNf1WrhfMK6iHrPNV/m/GZw1pABeBOFhzabW67pNUfGQ
8u+3a8jn3+Zf0Jten5kvJ48hWm3855DthKaroQ6WURgqPr06XDyu+E5DOP+4BZT0
U6TIaj/htRQWELZ+u264PFxjNy7ksUqshv6sQXBNBlDjxnP3xYZ8tZsNRyXhoBhh
hIxxjkw1Ft1lP+TdGdqJ7MVtSEaqYVugBjLdx9UeqeOF7/bkOczE35LChmKyBfQL
i5RlNQZXWpRQ8WVMaJGLOM99vOKHmpbaXy1VzRB0YQnEdiKKQeeE9Hgfj8uCgQYL
A7FM7MX5UUyf09o6OJsZcA9mXnDRDfGt5CcYOAaJZNLlcLjQb0EhdeHJuk5BUVuB
VnA/5+4Wb2fGhMUjoUlJeHGUlj14K6EVe0V1+dMpBOEDY6ozO9J1KQ/Qlum8dFhB
ffRlipbfB++Qkov+4BxbpPxVQ9Hci5Y6GJsZF33A2nxwLOWRcQuONULKkASAmRtZ
kV7Ax/R2Fo8NxhvcW8nIzRVQJiyuCkNT2s5xTFqIl9I6yuRBAZpYt7B817T0SgZp
ZnO6kP49CbcokWWtQIOsUr6vzYuFNclWH091h6Fxuho1POTQWUnW3oyXmc76AJHs
AZoepIJvOw7USLQLsk/GztHYoe4vDkNA8EIpgSMOzptLU1jnL0VtasenAFS6Azho
7sqnn+OPtPGt27aisnPtk/v7qe1+GFHs9o9cCH26SdLEzR/1yfkQsubQxmPndiJr
/TCG3S5ffDSgg9/oOxqXYrhTDsoEyLHPjCd8tnKphHN/kEr7q6KI3w61lf1NcL6Y
/jlmtU0hNAenbbQjLo4uopjaCqpM+PlJgovYCvLlCuUScwvSDbZwZGXV1/rTeshS
uDDDlFqWYFNTj+fX9KJHHD+0penO3Da6fkvqAukQM4Yrq7Iig/rIIXElGBypo4CN
vVeBYZcdHXl2+FCFsU1C37uiqC0w01WXyy3uowMNEf8iMXH+k+K5PYQ1eOkBi7GU
IcaXyxKs71XZEZ/WsIN6WPBzHfrWNbQItY3p821qo4nJAJwagzMbsArhaMDkC1UD
spz0ojdCPml+lDKcKEre4VwbvGS2nTD7oUwTs6ZWpb/NTAuwuSy8pHC3lSq94iMu
8c6DlChPJU352E3xcvEhaxEtuoPDAtGTXl9oFuS3Tke1Wdjt8Y940po2Z5EfgGxj
GV8Fwx5gezY69LjotqsO678OGphS4Ks5i4yvUUv6CxkSpkylMhopldLjbCx/OWyv
ll5hTfmcVpwkCSkcgZjv9k4HMU0FVNwtApoa1VDWijlKfpNlKitN/RMobtGmPZvh
EOKLjrlHqoVknaGIc2R028rVhcNc4remfGo/yE69CB4fVZm8gzZ5tJBcsgER7+Wf
iuyj1cH2/RMKx+U7d8iSld3LWFqCwaXmtZLCfIoOKqb+5+YC+rF9MIudZ/aE/u+S
9HB2H943fxn7jXIYH5cszYC42AzAzLJOS3KkNOfU/h7Gd/RltTwkpofQDLSzaBHD
nxArFz070hh17E0nTrMDBM26B7IL/dDAGBX9/sDPYYFVDI8VklGCf2AlTO5VIjH2
tvAeoM2qb3XvqivtYyI7z2UWIx7EUJSLSe80/p+OFz8KAUeRQrWv15JupKzjw6bG
ohI2dVfFX7ewbSiPToBc9MZ8a53liL8J/K0X7Kax7bK5HUqIUhvC0cr0zfGgi2Dp
kUA7qV55aD75SUAs/LvSVtPbH88SHpH7AEBv40W/0uyCZJLxyfnQPwjSTuf/kpT4
wOvj4C4xMpBT/z4zh69eMQmuXg7G3IEjbbV0z1+r4FHq6aTr2kpvb5JtN2FeN7O2
SDpNtG/PjJDAx+x8vRWsVwiDfhP9+lY3CEdWee8D3Nx6JcTVM/tweLHJqEkTwwO8
b/a7EqJBUUV//XYOc/gvcBTbqkAtSJmxRmqHj0EVmXs2ldx0b1Sw/CWgRKBADU4q
Ld51ALTeSiFCGnGovzr3Usbc400UVunpzh7AWFn2y02ElQHlzws/N7x9mU6cUv7b
4ZSSgVRS8qA4cCJtBRUqyoEqxe4xcZu11RkfiUerR2871WqPQPV1FaJfRoPw0R7b
lNwiAB22a92/SzypkHngCnTnuJgdH+s5iHVJnHdPyQgrLpVm6HU1dfK4zDYdisRR
7h/swerur+KsOu8fkaX/3mNQsNl59MQQGIVXQKH5aYcyY4YOPzgW8arGYpiwd88X
aKK73u2WOfAI2mK/uRWnIuNTf2o3In3Q3+gYe2wkocznWf+ZBim+Wxb3K4Kx0QFX
lKIHvJFSG4hAjeYCTmvkzpNm2MnlC07j8RL+lYOTEAoc4ad7AhTuPWVPQWimCo3l
ONhv1mJXGa/hvn39raYCBjALqI8mKmTsrZlew8KJSntWggGuM2hnB9fiO89frjR/
L/dqk/AD/B/otBiqmjtTioKaGJwNLozJULKfzGMksHfBd5eivaZH7FzjiKSFqpCF
988Vzv1AZLQAQcTiU1EG2n7uDOmHWcsLPctg4Ml80+BGDU7ch4eG5MQXJ8xJO5Ld
FDP1FCcZ/oROl04qKWIyelFZs4onMpYv/1w5Z4ed7gOddyWtJzHAN4ycImwKlOH/
Lws+bdLiSGKfJt0ko1q3MkV3E9xrh0X02/aRRFR4ETZPS80F5DezTd8moVyrNcEH
+9LDa6HUmbQZ0KJFg1ccmBHS+yi/aCJys9+JZYoeSBURtAmcneXXXM/tmZ9zHvBK
LTXe1o3V376ndeEoijmZyPubNP/6MUG/r5z/JP8xtF+bPmmEMrZL8XQ89l+3i4W0
1RWmS4KDNNxBsUuwWtUlVmbWHzeHeOCI4L1/ycP4eVhlNkP8io4+VvLqcKAjwoTP
3/dP4Tetr6lT25WQftHdgfnKFbEG50oKfTK6LagyWp79TLHChiA0iZszalnAn8wA
YUCOz2+U6bcvglytbdHabIQxe/EwQfCoBeNYjbXYum+WL6bTFM28vWZfIgY6aDln
XTCQrVp144AgNweBnegcX/LVHWkL9al71vBhOY1BOAN4ttvKGoec6PXhy3l8h9SJ
t75XTDZM5klkjPLHhlvwOFP4jyEI8X/cEN2e6x9EBGhntX+xHe1TfBws4Hf50x6e
OXDufSs+6uyH3IusjNuKRVPV/Pk0DQvc2aYT234wsX0efQV4JdpVLlF81Sq8dNq5
SDxOB9V5nw6Plag/ioCJ6m6cus3NzsOFggLHUKfVe8akQSgGSZxB35bj5/TMi5i+
GGJLjryUvNa15tUw9DVkmjZlLuh3V2Zmiu0f0y0BvmRUdQmXYffn4/k5H48X9czm
Qo9wwK+dauLDE+Is/zw+Y0Gnb7wiy52+7Kuo9rZn6uDfNeO91gZkPlczpWWt08eo
LRjr2y2nbfrF83/EhgxwhLdJDI6f6O1h8nXiCr2o5kpNI3d7e4DCX3blKKAaMwDz
+siy0sXZaQ8ikMDGSQc2jHronG45vnet2kbdjR7kgI/NR+AB6GyiZvf2cyGkh52I
aU26Vql/jkGU2lgJPzCQLjyXiKcAaZnVSzlKS0IE3/BXQHdihFGqV/JJYPAiNubC
X6hLZ9RynLzjqg+0ofMX67kZFGl+uBSiKvZyCx8moNriBm7+/UFDPsF8cI7FMO5T
KwKqr6Cq9zwLyq+FqHLkU7M6Y1NRCgXw0Q+isQ7HFlHXFc3ICZN6NwQGBcqlqqhO
uDMfLDySCIfmTqaJ7tTDN9DaIT7I1A8vMj8W0vohyY2BvaUgZJAdZRBZXfiswJWi
BlKitPsua3PHnuRyNNQgPmGTroc5k5PbxDGiIUvTwdplqF3NJoiKRSZ0saHUCqsl
omNHr+uxpdTC4awyJ/aSiMzfTcugQaCWiPWhRAPKB14YV+L2P5xGYssPgBiCxbYN
yI8N0AIDkIE5C+PRfo4r5RRUkAn/oHdbFvnRmPJOW0uSqPjeSDLYmY00bTRbwr0u
WIoXX6LFewVqsv7peeSQW/nflYQIVPrGV2wR3GN9emz3WiGsruIcF0XvvBFhby8e
7HsjfC9N0dePq06a3Z2K5DDDk9Xk/B83fZpNbqlwbAqVFGGLirkgI/6pN49YninI
k8ndYNU/STlJMRTt/ZRossCSE9FFObMX+IBBQybcCMKBmwIJJDb9FKnzMdny979I
mF7SwWvK7Ydl8opEbeWMVXMZXgwCi8UgHCWPr13TwzLHDmNL1g1omjb5YXtyl57l
6EIGdOpJo5BUqnV8qe+e9g7eqxSIpWHvTkvHXMeNca1H2ceFDFzggUZpCjy28f7J
7XaNnz6FlVLKGPxSt7ixOM55uy8MVwRnn4t7RqhHtOG+1VjHlQgBl1F/8/M6Y0IL
oTkzQOaIZbx/APOJ7MBc+YNyvCFX9jeg7Stz7jPy2zUm40O3ybOVzYaONpCuKdY4
FNmvXJXCdlnqVk3ZDukWAQfJRWCSgFjtPCxFmTRbAlD67dcV5OC64F9Kd6WCz0bN
bqKOKM4DM/MvDKizlZp3za271mQUi8vzxT+g27fcBPhDkcLac8gKPinJd2TqjcEX
bcjCVKlbqr8/i9g80Lt8NyVvLjQWPm4zgsqk7Gi9nG0Lj1XAIGpJAbdMrxsqQhuT
/4a2ToyesQ71RHct6xao/nu+a/mG0SOaG/6BvXTTmGpb/+5KuCiCCgGD3zIwUuuS
KHcn6qNYz7H+/UUyGcjJl6PtUxG/38uud3KqUu/83gD+poTLGSUm8jA5INdeLLOV
klhHEf7yXh5Z4A7Y063cNIFWJ0Lc8Y0ANT8GSJ4MI3393o9dhEU7grhZTBZssejp
VfCEKYMkFsJfDFZJUJF+95DU6Sntf5Q5Ai4v2AnDQvZuNgr/Kh1vrUl5rx7jgFmA
08H5CH0EVzCiY4MP8hK0oJxlnABEfpN2PUK3ya8tfy1xiztjSzlblW2+p4oMuaRD
+WE1+b28taed2U0LHQHOSqHl0PKfPcQOjl7NdcTDRTnQAVHPAsDWRBkLe+bMpcXf
Ub8XZ0ckCdalxXIiR3OpwD6YGmXQYNwh6f1KRJ6QNdFv7CT0AjbDxfl4FdJB/7lt
r7WJ3Drz5dkW4yWfaFtpE+jT+1goRsqvf0bzh6GASJ4ypnGp40V2xXm95FwgSIBb
Pg7nMpLvIAEfGkbgqTB1GlNIZaLJ0g+omi/8w7j+JHajp/SlLxqnibomYKh7QAyK
Aq9vZy42Ru66t82jsHCBcSQvPk7ycbiQlZjOgC/sCS3SayPNsyL+E/YZOOLGAlCV
5DbBvQug38t+2M/wwPzdnhCp8/qkSr4+KRw3HaNnuBHMv3MUWQymGNNJsqHwdIjz
s1dsEKBkh/9UtFKySCy76wWd5sb3FbshCuHsRYC29mmhI3ggAMJ4h3gbT9Bh16sS
ISVbDNSkVjEUbMNi4SgkhUelPqWBItC9yd9Mtl7Uo85EpY4xkv95Vh0GqM0yyUoH
2QYgK11n/OwGwa6jl4O3lSU847oBxy8Ud2DKxcGjI+6uj2Y82c0/oNxbwWgWmeVR
+SurngvmPr/wem9Bws5lD3rM1tPIItflScYiXKVIK9AeZFXggR6B+TnLPmTC7NmS
FC0mLCGCijLXYJmwOcuxK+FdplnSxCteZKsu/fAuvwx9dgyr7F/BP14d4JVBi7jd
TTXUHxtFMXGKg3NRDxs7syStih0oRmPOJrRAMW+ADu/4GIbKObqXpLHjbggcGmoL
v0oTDI75baDrdFTIDdZfVncIRSfVDS6luU5BzW7CZbiYXLjXRMOG8E9ecJ+MjCkj
dFE2MxY91gLDKK6TKWl7UttmVVRfz8QlqMfCSpS3wQDkLlgPDbGiPSbYms7XVrye
Nb5T0BFYYbNVDv08dpujc5rQ+xRnZKDtERx0UP4vX28jhlxdueM+kN9jYCx1BsdP
lI7jWTwPF///CT4UaEf7bFyIdYjICKVePrebbx+toRi2aSUUdm824ij9E2l/EHSc
wDQkMAXEFWeaxlHuBz8KYDP2twdAy1j0wdO/ARtjxKppZZK9n0Vpn4Fea9++zEnN
IqsVPbWW0sL7Gr07N2P+31cdiX4TBd9v0pe639w8+mZ8q9DnDRCQZ7V6iRJZwXNg
l/FSt2wbl+fSUhWD5cpKlF5HhcVr/7hTjQJqkcugH65C5KAu+lNWzmJr/Qzbahwt
VOUU0nBkVEETwfhP8lFbtw/fyU/qu4o7m0mhhBp+NuP3mxt7ieqT657lCrlQsTPA
gxqntDCJehmFB65ocarnat+R7rg/c0/1Syg3nAnRzlEqVCWaGGPSumP1HzI4ivfT
+V890Kd2vu2GcmnZZh3sZeiUDid6qiZZe6cR1Lvw+MvJ69emjNHVAbEc8cycRnC0
qv8J1t+PQZHS4duMTnzgnF5uwAB17wj+Km1YCd51cWn8UkdAePUmpQu6jvjRQMcL
cImHF6juHhrNXrjdH06LZ/8PGa0JsYNVNtl5K94iPxUykP/vGcz2bwlHm1g4RM6I
hdgOKb9Mm+FJ4m8rYRDUVUknVfND1lu+GG6fS1lbVhqwtVgImxlmrs4nGBon4fI3
GhTpkX9Tlk255yVPS1l6tLEgo9otWke133PrOJgM9naS8iUjL91j0MAFpOS7SEBa
7emJnk0Yc6NWguUN7PQW8kZW3zA+EPyl3GJalO+x8AEKlYAMDkMjtRCsw07BOMcL
zSpcrqfYXK8yQJqhFEDOOBEAEmat5l7/sM0GpcwWzUoWf5c2GX6Z8GP2CiPnwsd8
bj9aJksdbsxkqzVjv6qSKVTdQLm1j5Ewk8sBHAUFT0JzIrLLqVxx99oVurbG7j/Z
b0Sjf6Jouo6Ua3M5tz0tehIIJFcC/OwNTukIkblE2NNo2MuqXaOgS1qKTpws0/5T
A7dgeuTOJQjkdJiaGczmFTp+FQY7IUaRWZf0pyN1PH3GbxJ4xxhQVgFM7peAbW9M
iCJFl3SoQNnfezele6Y0ed0280p3TguNAccDHV+0QizPa0tOrbQPH+Itp0R+LRuI
WiJJejTTGnEcqdn8M+nkHoBX4RbRtq0AXjhG/pF0idnj/iaZPtBXqUJxrByjPGML
cUmkbHRYwzDrsMN+0xSnbo5TnHu/Vtwo6W+rAck6RdSg6RBQnv9c7bDmobJ2uLaN
3At2rl2d1lXyZGVrgJRRl57+GwGG0mjYgNcseWZcIa+nUhC72rcF0GEfuSsYZz05
KI/VG0WliVVrN8QpzOgXWU9utVGvV4ZoJ0tCvLrrhqmnnUC4bLpgKFaUu/awOTTh
RyVb+p14BEYLlqT5zFoqnVLCYeZB008USqO+wYI9LR347mEHMOIXPboNRjsLcWPR
0CGzUaFcpu1EOXO27rKEfRoxBjhpuTzJqWq4oveCVqYBzTeP3lxyVHB7LTPEdxXB
yR/nVq5irlYgzjrKiLlGLgu1PgFMpWSHi/Pco6jTIUs0e+cvQzmAk4h7DPSFjltY
Zk5CDWODsEiipjjHyZ3iaJCQyUsNf0LmUV8nkA9QUzO5zFcQTNrE7Rx1BNq5P7NS
tAuccTS/2NA6Gmmfh+L8YnWoxX6bi3bNdqbw15g8T0KmUoYS5bTrMW6J/iLMQ3F6
KYqpydSLhgcmIzi89d4ODqcSGTuaP4Bg+1arUS5fx3BF1vEoc1noHJvV9HvL81nT
TQ6C/r3oiKj/BHbNTn5wbPH4bTJzsv48sPKY9G/35KBBKH0GyDRJ1imQ1SdLd0jS
m9OroHm/ZEPpwHxSkW7A6I+B/fnhUGtBGw10M+5Urx1cn5vuvGgjkZLoTPYiuDI2
YC4pCsbptb1alvRvdsKlwTEPyP9cEzBlpcR4dgEXCkLPCaXP94+Hka78azmlwcoq
/opF4oyWsrv60kOYxSC6l0s1oygWqXm3aIf5PeqnT5bV9o+6tTdOrCcAHO2jQKmO
Nvv7QVzyGfIpBzl9D0NcBKvdhrJI8QYMRRlZYyo6mKi2w9Et26yKULrNDH3gTecc
ooYK3ZR5BZK+13EYOALmNoZ1hed3Pa6UAfi0Aog8ic+Oh5KIT7OErVru3fz6EVkK
59/ee10SQny9YECtxA2jCHampsH8kX8aclYRRyRVuFbFrQF13zSxqNxwBEJD8FU3
ftxjAOhjiQmRrq8T1FWikCn0RoYahiNu1CVXLz8ftTMLTOSygujQ42kXEfMbqEks
kaFZHtRovVBB+hUwxpa+rXmPwDS+7hpAAmAX3VjLRGRkxee6X1zVBaS7KavkaZ4Y
/2DWNKohfJhyxifmbl2Qm1e6FMf/hzateG8QtM1kguRBPkx+pGfYygMrsm7KuqrE
6irA/PtR5JH0mWwkN2mnB3gpdjWCYwPRB++KRSGM5isH/I5F9ANo6lTSJm6XmODB
S+NO3D3Se9m586JVsAAAptRcTrjfeVVWNjaA28Fz/deznyl71JtoD/dllRPH/MWv
ALu81A769AXPB5dYxgImH7CkUKmCP3T0fIYgyCUye5i6paqlEfn8bL8RVaB0Z4CR
QtZzwEckXAgG+7Z3VO9RSAP3nSKKpUAMwRRR8hNr/VxyHJJaya7ZuWRpWtHr2YUG
mZGsdep8V/lfGFBkMrWdFytBbYMkVg/PbSnZsyL0LpcCYNS7t1FaJIShoRI6jI7R
qjm7J9sMrFhcsFIARWjZ71GolLMmmA16/n3Q7xGeCkoqDugKGXWVCeJ8Id067P+A
TG2/YczZ/rLmXt0TP7TB6aulojN1t5rRa+5uEjgTCguLIXPwrzn72RV4+Xdv9hjt
qvpM7KFJ/dbrw2Fr/en7r2ibz08c1h8ZlBZuWCBnZbPUP0Px9Q4DjXNcBUfvZDvL
vNXp9Vf8Q1VS/j3E67nHNS1IA1gY+bqQJLTJr6eU6cgrv7YB+q0opcmL7qL5SbwM
QH28sfGo7f958akkdvbFGEUcWUAyavRn4yJtY6FNA/m+CqJ6B8bpaWI/naMklIcT
Lu4/5fAY9rEZ/OswsZkqed0bOxhRkm+CMXb98rqQcgCfJEvPPyKgbZb8wASEo2PC
82xWtnvn0P4sCoQdDF0b/PnrdIyXmp9puUD/F50w0I/kzzrNDFiR2rg4dgYyobyn
8T8tfDWc7+bpfzuuNVlJ+Zysm9DaXMCxnJdxYo8guVWyuo5jk9sl+ud4Y2L/4xA7
6pAuXUU/+bDqfM328qeOuVTQvKtcDRhxES/WnTEeia9tSYpGqJ+m42alWcLmQ8oQ
xl2tgvS81i5rCRSHATg781An7rjcmIpPR0507pozS4+bw2b2lCM9BwYQ81gDdmRg
+IlwqETQaYB3WIl8VDUzEb4fQ9iixEV6yQM21q7Mb5V0r88xH5v9LIdzR36MmhNv
SxVTXGP+8c27By8Ny14Y6cAG/wAKuKCpZbt0tf4q3LIStjKwGW8AKdLu61vu9ri5
CcraWhQ3yLsMowaKAM/tLT1dZzABojGPpNAUizBWohAj2k06B5BQYBV5+jjrE5Op
jed9LWtB8dFhCeprciT1RW41qzKFNypMcuCDkSc6nH14CMzmIAB1KyfV40RbhKAM
BMnl8d6xahYdeZw1LUJqxEKe0/8FuTzlO7OwTN+e7JmsknPsqtg+hOWdVmNIuEgN
4dYBt6JUPX9JxR8d9GajLDXi+IoW1/VN7vGMyQMnYxJ7O7BSl4Hd9x8tbL3qbuaW
eqMuGSX8F5OSkf7o9MY++K59slHvuKSwoBfZeWHK9sDNF2vwRMyiRboMo49d/+pr
4fVaAsnDCRXlHnVFu2UxwQRIUdhT85iqi3xs3lKw4Y3LtnJ2Q0WhssyeHhnzjXO2
zuPTpdvYUf7o5pQHLOZC9lGdxYAmO2QCLwFO3ZmktnTKHEqVVmTvz0GWlpIyIoIQ
Uw1K9aLMpCo5s0xnW3Lgq2gGWLBDuIoZGnp72wN5drA4zT2GMB2zvrxScz/CH37q
MLSaEOKmrX00UxBBTVPtbCN56JZevzsi5Wzn4OCUZDVWDBDkpNLWTE5c/VjbCkQf
bHSW98CiJpg0sKYVRtIYCCbc0zRQSejbrgcp06aqhJ/W2NkLPJsyrfD45BQ61jkD
vUG60sqA7iNJ1wqKF3b3F6zEyUzh0l7xuWS8bSU8dHK+/INQTCQeW4NjCbUK/66Q
mDMGbU1GwNcWilyTbDEl1Ztz5kfNfNDYFJJOg3CQn27ojbUpNBakn9sZgBbUAG/2
4/UZIZOzOyTTSls36CL3lIbf+2SKfK6xva1u4XnCnjvnB4AaJ+Q65Xf2F3Gl9J03
9fpe77/oh7bDupyqaulc1xXkGn3ACFUa1LYFG/2ecPn7X5NUWg9DGq3vmGPaGh6K
CGykNf922PXX19Y/Di7SSTUZfXG42RBg9zxGEsA31TfeyzEQCn6MntiaHSgpIACv
omLx9vL5ON5T62r3HA1Qih2+T7eiqtkhBUwM7sbmK340+egq2i5d8uMz+/lNCZcc
NHfJ6tLj4fNZ7/X/syL3cQDw2Ws6hsqMicn/5Tj+zzTzrPR/QQpWhk1PTIHdvbzU
nL58tKqM7K81Y1kk8CBsAriLgzZyB85w7ER63ehe8s5PWBt4BWXNqtamGgQi2gGf
1uwgkIWDZeRvysNVwssWYBzEpKZ4Gypkwv/s6BUWY+F1+xRa0jhvEUQqgjZ5rzUz
F37dCbuiPg50Qthycu3YTUobKZnJVNmNOIg8L90Fa8rhGpyoehXTIo9q95b62W/U
+0lbCsAVsSlVIlBJxgemnqoTeUrCvojgYnxxyKHAgawf09m72lm3bW8Y17BjRX7W
H2uP0SuCHdmUfj5oRVWoLNEIS75gCf8tKQwD5ypTh4f3y5bjUvcm1UuFN7uVlb9G
SA3H3KstwTWq3BQ6HTUoCQvsYZ8I42DVTJlGEm6hQatQAkzQddmIDKnirmvr+MYt
1tWJ7JxP6s+9WipjqFYc5onFkVZOnFZ6hBJBRMfZz7xey5b4XmnwJWsvVzi45Ld5
foXqrZTUFqFSGO7hbi0YYdA9VhMZdlpzxSlsFIpzYYd87mA3jheAITtzfWPTmxHl
5qrQVdjZ39LjPSvL0gYPL2djN22r1q/2y1mXpJ8XyxaNc6neQBR/6WdiPX42bT7H
YLeKofkBWGXZdDyFAOJ9ku2ZaLvjJMCuFZEcu6GtXLVY12I+WOom5SP/R+0BEFoP
giq+qiOD32e+7Ue1E0sq1tutYZCF5wGKGxltbt1rfJf8x4df5IKfi855hOPRXBEU
ax718TdnytlM+bIENTYDz+//vySN5ikXluLbFyDH5GYEpQfe5XEv9qbVWAZ+mU5z
HBRWkJOmx6zy3PmyVXM0UQdch2pwLHgUDovkAw3159XPHL/Nja4kqElB5V+a5Yqn
6ewRDi/YTuvPEYnWPWRMMbLUXxbZmU33dtCHJDHZrJgqGrrwxPkE7B+IISlhrmGf
Z46uugPOVCEYFxQcRzMCb/bzsbzGMujJRRUdD27KS11T6p5fR/K1iuIHs66uQekl
8Tci68bgW8Kc2sGZX4jPt/c1mJD1yBC6cdNEavGbptSTPsEN6MS4v6Ka4l3i/ZEe
K5SyLO5mbPbYBhaewuj7BGP7YNFclrMlp1CcopC4/iQKBRxY3wZ9F3ORKcPabohZ
CpdFD/5uhNgGJXfg+kG8e/gXbji7FFd4C1xOwm26ZzQfAfFasRyMCuZ40G4DiKPE
05Z4pZDLdEsyiW66kKYBU78WgVe7kalavKZsWVfQDrEHwFyj3N7drZfX9e3r10WR
ZcbLb7PYYf5m7MM0KH4Fm5GqsrO4WXn6VfJTmwg43emkS2zlVEq617vUwF9QfzjD
I4zV7I98CD2GuEp5PmznE/YDYdAmpCdo3lZEQuK8zFCEndtMXHpdmd8SQDTkQrhA
iYw4h4UpCiS7kkV7KRgmjY0CORnDdvd99bCSOveboEIj15BqIoqOroN85W0ZQ9cB
kZuUTvlWPUNvNc69GJLU8mrTHsAQv+bcZgQsOMV0nhcyckW6PA0hLIWdes6px9jU
5IrRmztyCSdVTRVfDiyyZ47jSijq2ZODksfJAEgCzQTx5cRtqHjR3ixSyCijLRNM
LkG50WuOPAtC4LSgWVBsYsNwyBa6L6IYyWf8VGiHJlcIwXvwJ1Urb2XOZHxYZN5G
AVxS+RtDf5d8OqENc85r4Ru0coOQd84xlinIU5m6kGOot0Yar97bnbI3ecSghr2w
6P4l3I68xHiBNruigfoswBEIirxQr3UvztfoFObWzzjb3b19qJz2UXHqTfKyb2UI
y3QKivgzRQqo8LuZKdZhWHhRUGUXmOOwz+yqxB/ROTeOhi1g/D1ZxgaeynLBIUC6
E1u/li4SwyVjJJrx82soF1V804JK+MZCP/Xb6hgxblbXFdlrR+aKQxl2oEOnF5sO
L0u4yA8cwUHLtdok4sfUhdZoq9XIpyaN2l/FgHOBJ4ILsuD/ASbAhJKbuEG+IpQG
mIjDpvw7+ZT1wRKcFZ5dvPE1fKAcsNgK1IPKe0ntUSqOiJofYxRRkSWlFWq1cuUW
ImX4aHjM75QOeHSIkKF9cgxfYhlJx+9HbcF0fs909C7FSAg6IpzUjveLDH2oeSsA
07CA6HTRzIU+nRaNJXn8HrtK/e+42UlnDMoyaK2hV2K5Idn1KljcuEJde1QaPUJc
q51s5EAT87i7iHz1jz48A/IZHWTItPNEjTfK0SHC/ILgrkeVoL0Up952SetEPgry
CnpBB6it+kPiiZeXkCyyj+PnN43FRsYRClUYy7Clc7VFUk35TFFa9Ec4R5vE4f+k
yzQA/6yk1I9S7taSqe3tHM5bywv7bpiWCvbOHOKydfgk/Tcynm2wj6aZE/xIsR+S
PqyYiIUveM5h6/EfJul+mwyq3WosXeDJUi7cxWIAsVVvJLMCURgjuUbaSF0waGPq
gcp/Q8SeGmdeHA6e/yysgtiMIctpkfybPeknR6xHtJD7kvpgyD7+T80k45UHsegP
WyPxY78Fz8E6OpYn76i1jENrZlwcwxPMfpBfnm9RtZXzB1yUC9C749qvmAUQM2ML
42iYoZkaDeLzjboG7pNxIC+GEeLFninKDBbiN+nr4uMFqkjB6VGqwkptVWWGkAjg
BzcSh/Gv8GDEsBrZAAeata8Lr2FBNR228Ifaj4JlLKvVkKFGUvkQJzR80nquSE3q
8gY89Bwy7SZoL2Tzvd8FbEzJaQ5yZWuarQYBH8egRiLrpbj5J5MQK+BsTS5Esopt
CQtLU87ckOTU3a6RYdewvQ0r6aRe5ytcrh0eZPQRfc8m0dW9wcxekQEsLVK1dZY2
c6rKcJ+fd/fdo4dZjrl/HyiRKB4ZtgoY0H4ocl4truDcCHr5HU9+QWfqF/gUc/5l
CVBYX2j3adpbNRlDkgpao5i/pWJRAth7eGeQxZL/ogo4J5TRiruRgPrTJbMGPPRu
jqXY4hmdKYqh08UBDKgED6iHUIvOrbP/SbD95yLTFESRDPYqrmml73YXph5hWzi4
iYqT1uNY1mDztJrSWYVaScKNKqAGHVwzYl0bKQXQ3hngUo/+j8hj/h0xD+tv5AvD
QUCoo619VHSWB1DIME5Z9TMdxwtK9iJ22rJqIybKvGEDQ+2/TOThcjK7Y/OtfD/f
0ThQDuWwqCfPtECxawaQwJsGO4R8EtwUvF/oBGx9baEUeeXW/F+mNbLr0LyQG4rq
PazEmnVWuqjRvbm48Trb4Hy4mGdodvtJzBD2P5MMUidkGgAfP9cZjiWruoM7TmFW
lbHZKq4H5bJEHN8E9uIsso0WzoBEJjp/Z+6tgHLWymW+qxJ3Y6Etxf7hDTB5QAqV
ToxiU+inbnZKcubtGS6aHZKXUJb1IUb1fwv4ALV+UJ2sdadlb/6IGKLDYuqu0EFY
bv2+TKnJW+/TGW2kvOqpBKoRmNCkZ2iy9eLMLd2tnsdAv7SXrDLrIjwPvmACe8Zy
iFYYcpyMZ+uLRep8/Euk/ImnfH0t7iTIU/1ZV7EyvhnC0qHLqOxR2CdrB/3iwh29
SW2dPFXbU5cvW6370kiauqdx/B7gFeP05i3odMTLjwNGvWFnZPfl1UlxK8xgILu4
d0UjZB+sMNlpHex+hpO11mn/QVzdVBnu4UvSXMxGoy+OprGCBqfj3f0XSsj6m27J
vLMg+YaJaQ726Ifv3J7AjMpnYEsG87e8VRdpoJrwbl+xcMv7kGtxmf3WSKlV/Klx
HxT2w8zTXmAzrDvz+hKi9oDANMEjhHOb42Yr/v0+c6vqiLT68yfFgOXjppj3AW+i
p8YZDchdhELtbP3jvpy0R2/DkK6lT+fBp+DEIcAR8saZLNblOc88ArSUSKoPEYjK
2VJ4ZX23XYlNlpMoCaf3dF4p1D/pojJcqtNJQDyOrEkO52y/CefyCbRPYVwGsE4s
sZmVywG8+83fsCfLmWTNbPFbMZzBsrOvGdZkXKKvxzIYCMbCE9bowzlXgQ8UxqbO
1m9bs97BQhhO9RX4/6cM4JLBNxHxDpuqfcqn8PHwSjGvjuAVPByrLjv4gANFAjjS
3LyKuo63s4arUMQI3t0nFGRu7/29kSHikpZNTTv7A2FHMwwk5mqjPxUnfJIUW2db
U/rQLP8ZJAsUWO9s6exWxyyRi5DzgHCe6J2QSgfU2Y2IhzWXFW4TsqKaACTttbqu
qmtzIfg2f9wX5nrAGqJn4FjcJb2J3bUaTfXhuU4n3Jq7Yxf2pXP/2A3mxBsOly6K
NWJiEIHZZpYCW2M74N/ojBLsYTjwRC9Gh1pSCisVP/l7ceK66W5kZWVtWHkO77Im
ODZr4JC8EoSPaLNsBmuWereWwwHvoHtskFvC+nB6VxvxM6YMZQRxeZiZU5JpA474
QO7ZqyI8iE3HkAIUX/y2bMft9JQFxs0RVizDEu5tfIDCHEr6V5Lj9R8s/C03Rn+Q
CTLieucri8Jbt84p6Wv7QeT/VUfyblx8R9vTUzDzjfDvvp8G3wKVJ3iDvUKyTECU
dmj3k8FUm5xqXGKqTpr8wqX5w7y6Ad89N7nUDg4w3uyFQ8Stbhudzq/vskX5Ijkv
IdU02xf9DbOQ5WRTyJRzoDdAwkkyXOYCZxJxrNivrgH1oHo5/h+5f7xTmOn5F4zQ
C49xkNEsDecvBOgF3GPo4SBsLUVpcW/JfKtl1sMqwZYnhbbiTpqFi4s3lFxkGUJD
9vdPdh71m0Hc7m3CP8dSaswdgH4A5ijaT3YkJO6zTZ5KKY0l5OwTXWwsC4wNMLOl
Ki3JOfojjz+Insdl3fA4WjWqV6w3RobNqqLUX6ZDUuGjeXMsE0ICp+yDq1XUymTi
16XH1psMK+hS/v+rNkRy6+DdOcHY8t5aBzEYXBwWaFFb3hsl1l0UVY6yuefNM/Iu
JBs00k2CljoNmmrxpQYmU50YBCtbk+vMUylu01jhSE/4805TjV5vqT2gjv/7u9mQ
T7OToRPWuRJuLAXvzFCCL/dWWQqDTx83lCPkobbLs/bZmGXfOa+DfsUBsLx2sBJi
0J2YCAeCL7x90RzLuWaVsMiiOGnAMRk7tFdWr9JR0nfsTGHqEy8MDzMr27PH3t1L
boOiRdKR1x5V2wZLN1T4MxWw29TU7oEYVTmV4pTu+/CeBfsNt8PazKEL6diPbA3C
ZOoSTp4v5iOgTXGnifZpW+Kx0IErgEUxx6/I2vkTK9sLkWVc38ESHvdXE1BfFhXA
3CQgrDWjQyN3JEF0fvvK+1zj7gNdHud1KpaEkuEwrlEVZyWYEhPiaGnN38eO+BX/
kIzRCNxgL7jqDbhI5S46TRS8qQRPwXTBiS1wYX4PtczPvLc3mGgrM/uf7RFIvLhJ
n/QAn3IIV4uArrtC3LKroVLV8rAqYdgC5j8GPocVvnNrqQqtwa14fsfKut+Ix9ha
Yzi1iWITyITlo9+d+RRhE6cVIjtBaY3y+jzwmAPRfkCHAdX9rl6VuC9PwUsbbIXo
5YhVHGR/SLbRhj5oW+0D/HntnLcphVNyuTsFlH/WYBz6gv/LTd3K/ZOq0/5/hxtJ
3DFIa3K4h/hAoinoZnZUXJ8wcMM1xpmbD6mlZ4QCcKT1wj4pP37ovXx3fb03dPCQ
fyXA8OiiDrDrlI6CZKS1J50106qUhsu40ej0L93JQjte13oIEHwDe7g+e4ZN+tik
UNS8rDvMubOGC9nmGdvWjf1GOdD+OtZFj0KxSDis9XdwVdb5g9Tyo+W5xzlTazlW
mKiig2xOKfJ33v62NEPrwPtuuRiKQ/SGwIA/fYX24dW22tWBeYLJp1bU1RoXoN/1
koDjHIJuVazSXNLRv7xYiilNDHtAMiZS8+Z4+ubt0ZEsiLWectlLm1X8rCsvqbb1
hqCu+zPtBoAR63I4kzH9erlhBi2FLWiNj7B79qzkqHsB4B4iKaMnlnbh4BnCTrzB
kTAp76teN4+0JgHDTyLkuo+D8jEDeZovW/fqpxRx4k9IRe0tZSK3nr2a6fQxa6Sg
HocJWj4KN9ZO0sQkhIZ9U1P5tf5FR6ojnOlNPIjzPu58ChzXV4jYi5Ifv0jMPY/F
i91sHCh2un5cginb7+TnUbbw2izKzbHO3gUjeWZ0bEIG1SaYssZYRH8VTm32b7nU
HEzkqWKXbAS3+prFJAC4xyLQEMuaUqjlmkFaRL7MwwTHTW77lyLB52BF9jhpHXT2
R9tB9LQ8O3IEQsUXGyCLdyTXazceQHBig5/BUhdcG0iHm4jfjD0cRDeTzyqBibUx
hkbW1DE7U8S0IQCWEfMO4eptfNLtNo/u3ioeqs+r2YMFQDpoPHjroUgHcjDe/N4t
a5HHCcOCaxqDYdcdSEzkblc+sLeJERoD8VogPlq2Gguaz41i88z8QOqapO5c9twS
CR/8TrchUtzz7M9VGQKlFNkht8nPr3zV1Yewatap7UBC4jLbQmOFcPIgWv7BFK71
wOLtn6RfMOCPG2gAPc2EPf5CFwXZEDI7WRuTYggJAHZPg4ORl0xFjZrjycS3ARkY
+kgP4I94PeuMBQ8nJLHF/3uOwEilAhpMp1L04JemZ74ery1X9LwjU8v8K6HbpDUn
Kczwy3Bt85ERaRFhQPgu/qJtp6xx2p+Nh0YDNlVL+2K43hVkyKoiSmaqQ5gIdsGI
4H0V5a0wPbXdWHhr9vBgTqA5xvLrbW/P4L17p9Q0o3P+jrUNEHo8tWGEvqX11Fsd
odRA15xcGDDAfrawRQH1PwYjXOwo9+/SC1uwgxh4VGV50tVmi9YaUD1H0H84vgZt
45hnZhpzfBgzMFrbN90Uh6ElqB4Z841JfOtYDBKxdwn4yrPon2hA5DWUrKFmp7a3
RdtwefptXYndsuDXCl+A7vSp8Xd/HlbdWyoIAVzX8YQs9RREvfS0omcZa6Mgzgbs
pEAjk+YNNrtBaFUBbG6ObccPqFZ07dffwOnoi4vI89V9f0xvgb2wQL8d7Cx5a/e5
HLCQYVu+VHDgyiftg2TnzFgRrHMK4OxEmeXAs01Nc9PUpEg+l+Ej0rUH9wffwGVW
x6e9PTacp4GCZkNsyZXqiEjPgjf6IcvhnK/je5BYTGPS9bCXblDJHvjTAIZNGdJZ
MPfxE13X3tJRP7tSuBR0hN7jASUTTtZHwghh7nIuT8vIwLVHssf0NfHH35CHOYau
Y1C11REggh68exRxYuT5sQGvni+sPy+hFhvrw5KE24C/8iAMhESP1uVOg+eBVEq7
3q+0UcxEsjTBJV/fNhudHuhepXNOMPxbY3cjauVGgsF6Ka6mq+8RZis5HyFxY68s
Hh0OTg8n12WldTRtxUiWakHoIUo26DGV+jPBouykGV+7voBIgEPrMPHhgCcXilte
IsoYl+s96coUYuKhCsF7A0NIvvvfM+7mjy8dMUFH4ZCj5ynjwEzgek7Q64QCDyhy
nPm6rLNSibE6oRDfr1SYavd/s5XXwrnRSi8FlN3PVNTQZF0+NJvd0QC9/UdBMl8E
l2/6DeslxBnWDRo5rmSy0pIhMNUM65HSOb5QZHm79BFHzd0Woh8WvxcvLEDRzMDl
ymclZ6D1JsHxFUaG4OG63pYgmS54CQ8OPVtCcBrHdCIAiPgUrkDSLah7u3ElsN4z
E+sBQYpi0vXpnklS3xS/jVgNwQI5h9qLef4Umiz6N8Sa1DMd4WU+TrGGvKj0uZLh
4AkxyzBAoYJokeE1MOFSWsxQy5HoFPIxu3YL8GqE8etpEqSqkudlqzLwn82LE7C2
FJPdU1qnVuUhlgHbDo/6SrCKg0Qz6xmNYwDoUy5Vav3RF+XZPRIt02VyKMZpgJa0
VYIO80FNxNCMxPKC/+16qj29WoLWGbBZ89PRwJbBB1MV+Cvcqd+Fk6kgKOOmesXY
Mwz17XepHPRIVbM4q76ECf3S4tC3K/FeO6DmJZFsGpj1cIlIr0aGvcuj9bEhaAm8
rmJpFzhfYtoYrtAt+H/X4SZbQ+Lq0mk9sPprzeu9L1rv7DOEc9LiYsZiWW09cEhQ
AzbQv/owQkmG+eEiz+fXE5Zr7a9gxW0tP+U+++hbUb2Yzp3J69eVB8dtnTWjPUUy
DGSxbs3sa/6VdmHZpp6Ry0VG8aMZQtke3nMe352LU3GK8Dr+EffvDlkWlsA9DOBQ
11+MMYkebTRHv0oT8wv/NdknE4cYE5vmVjGzhpnq4MZklSpD6vRp9KnuBy0hBLHP
MWQBOz/CwS0eW/iVaTqLzTXzw/zkFsPUUMRcbqZWIUZcZbH5sS6Wr5ca2UgqR97s
84F3mNxLTTTuGIj6Jv4eNlS28s8YKxAx/y7+bwGO+3mysNAxdFunLJ+BwzO4k17/
28sXK6vJbB0HFwxGhTzYATYZGsngyhgnsSiysfg75zjnZbsInGuqcG0MC03iG91x
Z/+HhEZB9BY08so42AzPL9G9J3w/wDk/uFCj4wUuo3yi+juprKc+gKU0M2MYHUms
iTTj05mUc9VL0CFEn1kKUj28QR0uswstjKwbw3H2ldCcwct8NnbMOCLiD0bEw+N9
EoaVd5zjKehkE1Q+I+hSQucWlcsC/gBxuKvOJkVpuFkhJ+KDpvdH+8GWbIYhjrnW
dUhBPAFGOGKgAVuu+zh6xhJMFsduPyyX6Kb2A1PiHBl0EHM7PCjEWUsQX6yzR0Nv
3YS+IlpqozJ2GvRw6pA1fcaj87m6chE+GUJDb5M9dQvLsp99Dv4xSsQm4C9BuIvj
FoanVSNTDi8kfboXO304uQRHLkU96fjIE/rCzHCxqoI0vX0HMvF469MkQh18wAgu
IJg9nVgbSeZGuiylHkkmKUVxbiNsCMew7PbItATcv8UNws15OkiTe9X6caYpEW8R
2rmHhipOvAkDDyQaIgfNd+bFV5WP8EDvKSvujt285nLjRHNty13lKIQJfdoHfns6
rgBP37uiL5TgPefauRkYzBXln6x+/Cq9UIc4ygaMqooT/YzLEYrIm11Oqn2rinvM
XrjVGE+PQ+HIRX5xHYYt3DnhLs1wJoQkpwAsONnvMDdBMbS/kVcrE0Mn+wz3uu6k
961QSjkHIOLLfkT4C24P/8Q5dqjbAnmIQQh37Upi1/9pqXAsmFoFNZnHMOp2KOWw
+HDb6j+qBv/6aGWoHdUMLzkKugR086zn7PW0OjWwH1qJef9Nm6pQTQ3T2KMNaKz5
a5TvsR+NZf7fQl6w+7eZ7nAu9O4zw/qYPqEfscyV78k16FezSt1PYd9sLBzEpLfM
HgQljSk/awIuDXocElVssj4/3jiZgGIJUF8jOo8D16Eht41semxEe4ndiwgKmuuk
50aRzRsmCZoiDukuzTM8Yq15K2jhjzkEqjhFFtixiV/t10Lvgg+tyDJAgpTWYRuj
8z+JipyKGCWUQD5lvo2WoISOiutzTiSjnrQIR1vWp1r2D/Ufyns4q6MGyNGpPTtS
1GKK8VeyxUAfgCuAcgw4qA3KfygwpJdsPU9w9Xz/+3m5fGC5dcHipIU/pVzeumnf
a1u7iPsRFMdROLf/x6p20LghY2ryv2XJHvosyiMiHrhOySXPQHh/wsOSRHMl9fu2
EWMZp05B53Vm16OeE3dK6PxdGaeOpfyMLYFDds0Dy8jhR8Yd/BtXLk+Jbx1MPNDA
RBs2RcdJMsQxTPbejA+AJVOGLdUAabcTaDAOZNg+a2z0A6S684jsFS7jBS5+EofF
7xl117DbJZce8TkHoR59H9B8W9IgAkIMaHc8cq/YFWAjLSHxd5GHI5BRe2lJdZGa
xn38XbuhwOhoKH7kzGJsTCo7GsfKDEj+uZShiDgKe/POPq0KKKz0WrYvD3nYsqtU
+8jKZM/4HQF2jFfdYLrBBZ+lngNvCg/esNsFLO3sIxcTu6TzCJ/agpfsH0NeunSu
1lkEvhpUlmEUphnf4LOENyYUtVMG4cKpk2TK7tT/o4I2UWWndqdrJ5uvBoQZ9wTM
Z5X+p7Nk8xAKvNK4Za/VYP4AbEpcsVvOGPqwrFKTxhENLhE6aGeGkVlNMocuhidl
Z6uBQ8RoI5umpC35QeT1TDrwZULXHTkvYihnRCS09wgBYDnWxaSl+9H4wdUiaURa
f9JqKgTpeEHk9TWIG9Vq+I04RGaUhpyZiXCt4167Q6MXIH0GA0da/Q+OXTYwmql5
v3kmV0A+Udw+vJlwPUyJ9IqR8gZVA+GK/pST32vNuBTe8ApPkGU8AM9IOERBBt9+
Z2kORnWEYru4Dx4WSzyfk5aZpfqki6xP0XiOxd2NyWnmJkPj0/IhxmXpElt61Cic
ZY6HGtEqBA9KCsiNoNdIMUsGDHUxSCnYGH/vsPMPnbkMpQhIxsdiCIjoTCDzlPKi
wCFNgAPrMQXCwXiuSbZvazMhMRzBAuU5umdw0HWEqbaccNtH80lOxQjAsjQ0ZfHD
LqDA4sm6sXJvMYMyvCFSLYTmgEtvF7o+92/QYIJqKn2EqxcC4bMStLYu21vFUd71
HwrbilGtEFoAvnxlFZ3XPM8VexfzWcR2VFajSOMJIdtDjbKP7Dzgyd9s/xsoj+Gw
pP/R0X69CPS6w0jrZ0ttCOGuBw1O6obvAwjhJGETrVNELBRpLTVITmBzUongJrhH
uBJEqDkC8xBbCiCTZesLJICmLSuL8X8NCLqRYDB1kZir3YrrXRqLRhuAsvquDWgG
HFQT3vTGBZUKv/EfRM6sYV8vb0zAaX8d2+3svcMVwdO4/+iZ8A3UhLXcZEDdh4fY
xeaGpj7qjPcNVsFaKb5wA/odtsGzVzFc8un4POAuOPfnpIN48srkJcaiGjhcmlKj
02GBRZiL1zEpf4KCBsul0jnoQDKIg4Ff5JPgxnWbFrMRaGp7qOE+ZEA6GZNN0c1Z
nrl0GR9kEECH+Pw50Xk8HSPjXGAhtRKNT6SNpRTgss+DEiOFTGmda5Hl3IbohRtt
IfrBflMZEEd1UyI0RatI3IYNPZZ3SFdOwZtg/fu0NHGFfxzTYfYvp/HK4xnG8K6w
n3ZGhaEX1XPI9h+uKhE3CRnEV8xZqKwskEoIm9QyoYApcoldc9SvVwpe3p/C10jg
LazZqL3jDDxKzAtxLKd8TAS6nUIZpZhj3Yt/UNBt2FA4zE2AsaXVLvqkpQ6ruXJ5
nE334AXfHWb0yCNoV4oi3dmKflJRSTE/mS2cG6y78+EBCsFwEEm7GLtLquXKk5fD
obFPMQVHNvH9Zk0Rtvw/ugrnkQacukP71ZV8GJoz9VvImTnwXBv6MqOJDhFhIZ9v
40UxHWUS431QhBkTBdR7au+yguMXkCuJaaBkD/mVbu2w+0RFycSiV6jhR3Yo8e26
t8mZNC5kf9dN1CMlEBIqa6bWme/oSyASnANcwFWsF8+qKF4gDRMXKZdN/ZG/m5au
kE39Sdljd6P43yk5Wh8C3p4sGHcDF6lrHaNlPH4s2g7EifZTLVELq/rud/UMl3UI
1tiiq7r+y41KmsxWRmBe4rq4wNnUIwAs/EEH7L0HIMmm4tazBjdjJFMl/UopFZFS
nhYxSByHnbXzSkpGgtbUGxW7pUs0VYczePEyR2tW0xhMI8lY9qcfegknOkta4nYO
JyiLOAfbj3II2fBbhtwJ/VxKwTmnF3n0dcyIq/nH/44H3e4ZG5A+mfgpnurcpPSQ
aTwgTflVx+QtzxLWN8/PuF5tOMwRyFlln1mqlmb1IGhANedru+Gf32WXiU/2jEIy
zj06NjqE00NhSi/EcCjUVp9fKH7pv3jEQnrNqSu+PQlup54/v7yl62zUpBBsdv4i
KfQB6AN6Z7EbpoGnLSLmahMgHEqW+soZNXgoakbfgJTPtRBSOl1Mif30rXm+Ts3g
HOpLzw6EIMIMiV+p+k+5w7tjN7OSYm5RKpNANMbhfnQB/5vt8orfrbZ5CLVCjQRo
ANbsxfDcihl4keW+0FnQpNc6dR7DicNUh1cGwdcDkogDjwxC5OLjbI+1AcoJ95OE
3to2vZVrULNn0cS6yCq5LWHLqUei17eUVYuUUDWKBZYo7Yp0a3NBhm35qjmgZuIn
HPKBAOCXDtcEPvcP69Jh/eDd2/7lL3XpLlVa0ZhHasLvwNSKcfI43Eo4ir+1METX
RtiDw9MkT2gTeZ+rgX1ui0Pau/fsbKtRB7vvBfRJDYVOXW2kpk+HbW4hNAReVGg6
Zwg9cap6Ot9z5sTnTVOYtFJJCFpCu1YZo+EOa2z5MB3zU4mTmmxdE72jN4hlceN5
fn5Po4GGLgLU/ZtvVpROdEoZ1VxbEI13l+SfmhWWywn5SldsgOUtccZPUcgXR/5l
4HlsNuZiL1Fa0PEVxgJer9heOCYMVhZ8ONec79APpXOv2VudvJv15QDeAPp5SLW0
9/IqreVGu/yF3ByhmcX1+RMGcEyv4e7Fp0DvSr8YR1070MBfD9Q2ejHkudT5W7mE
lV96JExj+pmviWEN4OQtE/6KFbQPwesRFJcodtlrha4Uhskv3Zm0rj7R7D0hqgXe
5MALpLq89yqp1mXIr11H1KeSkxBHCHcBwlWmDMFZr3HNv6FFB+oHLjIjknA0PE9B
QTe54m6+cQ0yywpNay8QEG+RvwwKi6bS/SmlGhjU62L1O26XGXUmv0/nbPBbdjsF
ExcUSDHW7iFuTjMzjCjSoSrQCatcUTqoHLVROp4tloFz2ay8GRm2rx1GpdJdu11C
KLWSciBp12joMEpqffd3ikK4XreeBgOF1yjxxSCs5HY/JImReqKXJySgKGt7ACKD
f7dghp1vF7rYYhd4OtESQxLmcaY02gulJVKmpFbFp7YqFAl5nEmroIiEDw0oCmQ6
Q3ggqmsmkpKZBeqZMXNm03cNFcIvAfQ0X+2n2/M33F8F2uIXQHG9Ek+S/0NLzx4b
z4LLUHnMlv1V5/JKodM2TTpgHdbzoS3hk+ithzUA1AkLqinbkeVzZJmXZ0dGWW8V
OJixljZCjub4gQs7t1hZnTwUZYmQ++IOjo0lMbnn5PzPWt2Z8F3K90Wu/AMClo6Y
A9s6PmVvGWC69FTNBcb0h7I+HXxUXS+a3/ctkbIgkI36gj1CFmwFQQOLnoeIKjR3
9uLSH/q0zE18zbwEKn2HrADzwG+ZttENAx8p61mYt2Hdj5um5Zdn7NkQ6Ncn/oIX
7dOJMcbt6IUD3eR1q+vXOLAanrcHPFDfnRnmSwMbxUWY3UhF9wHXF7PBef1RkEsT
uY0l1bP2AyOFS1YyXR3+jhkFe53rPb8NAu56kkGcuXVyuLjzK98ApmJb9R+tfhaL
1vIScg+sd/0EHKTkgyE63KtKwrn7FROUHOYNKR88/6cXM3ERo4tMHm/GJM+YEjtE
7f7dmkKHcGXNX1zw1gw3/PoHGWZfjhd6sg0RR3BQR4byutBrKiRJxXHnzjRHqHlu
VhExspWxbftkYqQGC79Q5aEFYYRxbnR3GCDvdZFWKwd63Le2BtWoz4F8ZwarxqMv
gU/NWg/+F/kLe+Efot7PP+RlzkOxXYpfVxamazLTHq5DJPnIiJ5kFQWFmsWoFgHx
5JaHmwT2RzUUggArJTZ2QeryNGfUemHTLVS8R0KcYx9xT4qFdrXt8+1RqlO8mimZ
/ffC75wWXRp+VmwG248XOxoY2FayBIt56bR88rgRjJyg5IJCfnqC7AQz7ywWH6dQ
MH81ppEg/nU8yXqKlhhvLcPm+AQ6mtRPorPoHxGNdBanOmpJL3BydAHvV/3Xj0Jn
cDux6mQOCBY92zVdqzUZ0vv0nBOC+kCUmBdxPklgQTOt3oDnw/AGpaBSwW8S2/FL
oMPstYHN5EajWRE38E7qZBCZo1/ZMnCeXZrT1GMefLKlgaqGzya55ggC5LxNVpTs
pq9I1mYpqEKE27S/eAXAu4Q475+ViSI1vNxGhOC3oTqKolatH4MkfeD7ZB/e1OoG
OQuNFx56AYRsALffkLPcVpsgaViNx6KcOm6V5nKJCtFSenmFrBe6S/i05/TPUIJK
6oetzf+D2oSBtmAVKBoOD5vrh09vqqiwOxlj6uhmaqGYJ0gHsO92VD+Nfk7Oo1YO
GqqOm9dREeugA1P5cq86e6akBwbhd8HyokVGQZ0+VosmO98PBQG1xmoOte2u8tc7
vr6xnlH/Scg/D8lRYZMlfjqrWcW+HZ8wz2YPX7PTqpkhckzU8bWAZwg0XzYMAvvz
Y7dVx0L1Sh4TGOay7iQLQDiHlVJ5ox7LwS+wpTliJgiPNVVWNZhGvVnE2SoQAwCZ
aozBkTEtTOf7caC13EzDZi8JmR2Cp9oAtI8mEWNL2Cmc6b85SifhM/mPP+X3flEk
giLU9xqoPc6gZEtTpiVgRqyjV7OunVTlxVTSp6uN8KGFoPVb2t41H6gElK+oMj8q
xzLXyVLvuM9/Z2z7oxdOFuq8PEQr5plrm9ccidQhUNlG/F9Thgns7DSEFEj7m55b
G5IkyRkkaG5rgeFlMk1ni8+fNjorVObColYUzUKgqkvnXsVCyRAxSuy2e2Rwdson
JdiFUc0oRmGs8f0EWHoJ1zJ3ghjc1mlNz84V9czWxvpwFQmC9gsve+ZWHRI8gnSe
T58O6tecIfCcPWhTI4Uj9Dxx4zZQzkNjKr5bicd0Q8w4uoUSSiqw4R7ykyY0Z9eW
w0l+582dYEXC2+Hhnc3y20jyjRFKMhyIQ1TBTNZQTJZZbxHq3mN01NSXpfPkHg0b
TmQc5m9Nltws/OlLA2oHyacNP0prN1AFQPRzqn3wbOQf/9/a+Zyi9pXarqrBxPSy
QaEMzU7cHNojZt8vrpdyuvlOg5vf0kdHK7wsvWciEjrTljng14coqcNn4q6253a7
8EorQfZFT5ORlabYV0LNHJSVamY+3UvjxX4VH4PbBNI5QiWZ98AEbhlBHU8Q5qwp
vpsMj+YVhjlCtUdU3kBbJc+GAB6cjjB8deY9g0LPsCSsUk4zcB3AsmZ7X8STK+bs
lpn0MJL0Cn4ykLTqyNk0RQvC8szBx3KZ69Ewgcgs/dxkWK3kJ5dRcpJ2KY0PRnJF
FOSrw3FIL6w11L7hJGQ81y76sYllQvvlBNHnfMZJV5b0Tn+HNTwV5uhfpSw6yX+t
UHIuznzoBdhSqxi79lxlWpU78ETUauFd76rsXcMX+5jXr5uiSS/7jcBUsegjVTm3
YFaoJJIwJPEu+W0uPXydKQmH8QkWbJr85a1q/O/sO81Uk3OM2g7lQmAYQFyiESE+
AG5jQZqY6GpFYZx0ANWm1o/kLjSRFFMhZKhYMOuqUVOSohuznD54TdgI+MO/gCKr
trg+EJzTg1GWzAVUqIiXpqLo5e/wKf3vD7ErGeipPD5G13gwZhNFnbrTBi4FAwYX
z/uZllAWAbpqNNhuTEZkjBGcB0F5I6/Z7iJrENUH0TbfLfpd6fUF2/fZV1FXLUUs
ppEymgu9GlI7nt2RGkFZn8STDNd38U8Ke1En1Agod0I9eXBnlh7bqSkTWFXXSCDd
r2qP5DktKZDSBy4LMG6kTuInSVkgdlOfK+UnlFMUNXYCVlSFc32LRsn7b2yfo0P/
ZRNXZK2lP8sQFwLEF0JFxPe9z1r5KF2k9e15q6+qwh5jg3r7JOxUl/2YWtx1yoAu
RhrzvBi/UvDRE7ox0slAKH8tCnxzRdPDI/ke8UpBISM2dy6EUYTdhDUtmzgVBmop
9y0PFJ1ndkBM5YTHBlrPPhCJZnYRxE8rWcQfhbn0gOBs0kzP9Wb/7Rh7I3pmGTHf
Veid6Oh8mvuq67tRT7jKOOZDIKY1zjkqlF5uKbTErMflPu0wAMEe4nqy78n3UtnC
30lIab+BsWJoFZdRvBl5TP7/WcRdgQkIAkVnJ1BwI/6dp3xYSanLKT78/JFsvcYd
qgdYqySMjaMtIjAztnskEjov6Xsf4yYBGYfHoCSjTwa+/8Xipom6wbSziPcEUA8S
P1HV1chhHNhIjzAhUkEgFzN5+CHg0eeY0t87DkR13nD52tosFuP3KCz9kBM/bt5m
iYY/YX3KuYQuIwJGaF6w1lC7PwC9nMzj4vsgthQGE5Eu4SPy3sUbyAalHBRP8Sby
ynqpyU56GRX2QcJa+JFDFDLubjVPJXRhYsb0EKenx2fdr4Q5P1UEmJ5en5/Gt+PE
UFeB1MgSe5WTfIN1yCz+iittClpBg+Iw2MGVi49eosFQ17sianQ4uauuVkL1G/P6
szFSbszGV/CasLUOp/Q2PsIsq514hBmeBMu/2VQuy5gtnMe/nn6mo+tg4FgN+DNV
UWSbOPj2vM3zRoQQ2I9cYIJ43uRn9ca06Y3GdE7ZwUOKRGpAFClygRgP+pLPB7Q+
F+K+PiL3VtNdAXk+Z0dfpD2Gqr1CAHtb8BsbGE46WwXMUgsadfln4A9k92DkK3X4
joLH5qf4J8OJmCe50RtZkECuW3uE0SES8hQyLDl7s2f8GEJAYeSrJoRgU/6y7KoC
7iyXbYgmLtxkvSbgumZ1kc2TjvymjTwQ3lhjw3maJTw0iHtlmn90YjRS7ppB5XpM
/czN4TqOC8hliOwxA+URhd9xLAffeQhK5SgGtbe5aUDmBY08KvEkc+ehkVfU3V2J
Xlej8OvjiLgmTaTQW9YXsw/kEgmh/LpAyP2zyFhJW2vxLR6efdaiZmTft3PVibaG
8SxqeNtZ+1OylVzw/TSac60GN/ZmpFC1K14+s5vE6JRqNat2KQ6Di6uYj6hX666J
tczvt5X1yh+kGKLDSgiSAGoKTs94E6A+Y7jFVWBzHHNokpZSm1NCKkVyEf26jljK
jrgoZtRS2zLg2aFd5c6sw7hK5MnQVr5PqELl2TxXCSKhtVkirnyONgxKz7zvUiMl
fR0MOCMk3oYP0gDEO/dGZEd2oYYqz1qfYW70CYU6hEZ2oE+PP+mmaJMPTE0br+P+
pZYBABSnthOFnCxJ6Umr397+km/B2k8hu8OUWSPeZMn13n4pQBRWRtd52ycQ10wd
0ESbs9Mr0IjDGmAHI7AjQ/g1D+aXuyPX3by/8H203A3CasFU+2Wh3A4/KtIp/y7k
zu9WBfOMwpfX8SkGjJVc2AEu1DMIYmdHevtUppjQLhUv/WUAaG+eHJJ0i6mnxpBj
nJVoijfffBaduhc2+Ei6wwVCsuIouJVt+DGaNmoRPBE6RrV0Evbv3NPZceqwUiwk
aqww3LV9cAQdMJ4hNZWbg1V4iyxLLiQb2fYgI0Zztkq7miUS5e38Nm5mFOXw7DIm
72EApvrk//A5TANRWKOQ06zDEUkEjf2oMm2qsRYIIP5ID3VcrcThCDhe2j4rDh8a
Vog/L7JajUnPoU666dqfdM65pl8Xr2psCTjcMLYKgZlvdPIRatBPQgMDppnEwsyY
FMujO1jWQ1x2w+6fEVEobu0BfaE70stD82+PGaMRPMsOWGHUcId3/3YF82wkuYAU
1Ll1Mlpxikg6OGCoMEQIRh8veG2gzzMOZRYwOfR1mmF5x8LtPe9xD/sOUUZCqtpP
Y+i4it7TAa7iqG3rSb9PTY8yWVox1M05Ce22gI6kd56mG5ObgcOUhxPcRYuFDDiD
0KDQU/SENmQao14JERb9DGSuV7TGvmUK41uinfRbWspXkz9WjDDod+lBh95rZcCJ
tVBpi24lNL2t82o3D7knJj+HsREhcAknXjFQFIxA7tJziKmr6MjEtM4b1+tp406r
tAdaDsPz00Zs+/Gx3D54SK3DKj3qICK5Cz6Reo00kvUqdL4Y0ILUa0jbBWWcnFTR
8tmcSWv+Y2EYbKygHZngQ01QzVIxqKePHjtP5SqG+kKRvedzAJfURCLCz2usa1o3
WIUYU/8C7IZ0gx6K9Y4X/FQ8py/p9pPIAnWiiVZppdmvW5skyGB471iRMGXrt7ni
syRF2io8vyXawAyjLjLM8Z70zGoxp0rZCydIr14JbcJDprTjwEH5gnFRKVKnfrkb
0eF/tKNBRbEJtc3dmmGcVa7TfM3j83Ux5lbPJJiF+GTRGI5y7MAM7GgNa4nZT8Ye
2Ch7P0piAl16tgNOtuGZPB1lVotIagdhrttKeKEBmmV4OrKnISvuvhFP8trsy1jp
R/VsEY0mnjs5D7CxKwV7YSgN03nP8N+WmhtrkJHQ6DO2Xaj2aEiFISNFBa9q/Bth
N/T2piBSIkrlTi0zdpKY/lD1u0pFDQKtcNUm9EjXz3o3LNx9MtHLp0zXZ+3gvpAL
6odwNZz5RCvDF5IwUmnJO+yTHYF8golHxvVDvyBX/WSK5WNImLnrwGbEJP8acpY+
oEHaroRCh83MUTuStBg0OVu9Dje/APmEPg2W0IC4lpilyWhcXj/FojNF1LNh3P6Q
/SR/jlHiFb/3bhgPH52pphUbBXi7vkynshmDobtp9U1el7KLg0n55Ozs4v989aOm
P5FCs2FhzM1qBheWxqd0RVoJYWzxWKe/oYtsgebwa/z5NlxDu53j5NeLx3KV064v
d7SZpG+y99SFQNT8yPuBG1cTsiTDLA0Z+RRPi4cWysjtbnxTtorVjW1NkmSam4qF
vO4lG4ZcTmvOOkg74SLEmHJtCUxRfYWLSsVbBAIR79Ygh7IMfC1qXQ+EC+sdxU8E
vY4bVqYdVO4gz07suzUvpqTpyNlB4u7t2GqxAko36ScOVbr3Nd38MhYJ/O7Z6vFh
Jz1+cce9YXrzDCIWzlbXp3rQejfJ0r+i0gzsu0SurA6xwTTEDfRUuqcQnRWWENrS
bxTcQ8UPJOkCviWty22MFyUfmumSm1oxqyLUKtFsm+STVb7gZCIcRcV2CXu39Bsa
x4BcyL3G3A/4sF8bsEPigjMqy6BwpkzNQMlNch2i2awjcJV305BFoM/AdrO8nFnE
oNnvHITjjFGVvOQGdn6uF2CS6JZyb4Ls3t/pRfkaD4MbX7Ex7lL/dwT9uKpAI5t/
Hfgs9Bewzb+znnuGUTafv4cdyCC5E9wp3aslkJgzTUXwfbLJEUF2SrGmp53tOcoD
ZJCt3j2++fcyi2oUhDApQVyq3YWqb2DJx+Do2qtlGpAe+maRaXvE1MemnGOi7Af8
3lokQfR7p7zwBlSfPg+Cx+WwzncrsBFMXmM4eTfb4AEmh/sk9LPwoqCMf4afabGP
6OBrFOoLJzsMcmUW5rs7vUdciqGX+o4GdCN0mpF+8ByEMg6493ny3z+EVcC/MbWj
iKg8dSqDrfxv6tDibFXQcnjcHajj0GukBgrj1ydLtQRt0keveLp6MNFQ6DQlkCXR
THRv0uLEmf7kUqRFg5UfW7kjeNG9lMG/2aRX0nHIzPUczctP9BR5pgENat3WQHMK
RWA0E0pwJnBosWvbKiILRGbkZQY5/zRG9fDzmKSqcOxVqGFtT9rsPlfFPEjO40hl
HgMUxuEoKGDG8g+C+zAo4VLeHuIcqJaDu4KG2UMQNDEQ3Nkbzbla10TUOd7Fxmzr
wM2xStfLRlOKRY7QWz/bnW1xR++QDKFnReFkGDrMcajkBTeXPOrCkgC4gwtP7S3g
bi71Ghh1uLPCOkEGsqhog4fe8bxTwvxRjO/ihmo51sC5noM5edfM0+xQzUejFptt
0jxPrIdVRBDw0qSWdznRCJau1+Q92aVrIBZwl1tIoqtrxCfQJ5A/gqAminrhJaC3
zTahOfy8gyo17AS6+ls3wDL4Q0d5hjJd7pcuxTdVtrnzy8IlybA1CbFr3US44+J1
P8civxA4qEkGlsQqEeGquqMf2SvcTNw5Qn4lago83KKwrkVLaNKZZwU7GXb/a/AQ
ENYNGHs72t9g340NwcRH8Bj78JmT+/uHm3CBUd1ZU/87K4LgvsRZTuqgYF/zsNof
P1gCjLH+hyq3XIhyhIHcKuuJBCArKQQCptEAte1Md4r2Ynt7EQ/aq2F4BVvuViCM
qxtuUEDnXqXh7vizHaZmlModrA/t9SuD6FFCJJJoOV90ekBE5kjxy0WfO/RrSF81
v72l2mhBfHVu4Udu+7G8MmZL2mOKql7liz6IEoVVhHi9XmOT+JbLlUDuksMOVOFE
7IoDuqySdi6OZ2BmE30Xs3SU76Y4ZMsvNmSysFefxI5U5BimoyZWEO0LYPuVDwk1
N89o9AmUckZo5OveLsdEgYORB6hGfOAxvd3qukALsoxHfphAQ03FkXi+Yl+OjL83
0lwQ+d0dP5VP9tvdO2fXq3rF3DkbfXDPijfB+60rg8YTGBX8vxEq31IfH2c5SCIH
eWPKg1q6oP9LMIIColRXYKqjwaDX+DDtF9rkxDr5iLdb/CfTPydEg+FRr+QMrMZz
6S1uRjFFxLtABZHnFv1cBq9FrqZZ1i6cTxhctYFYy6q10/2nxiWnMqcXMP7lXgxr
S59su6q+lM2rGn8RbxUfIoXGAVmzJVC7JFb8owmiz11BgxjeA+kDH0foByp1CvZt
lSZFfYv/lGXOWAXhtIaAGXN4AUR6gnd8C/GdLxttdYFHaVb4Chhyik5t/TIG+/vE
zGIwUxxwA13I4GuTylTENnSh1+OhX2rhBXjTIjeRJ/cOonvUUZ3ShRbCYt/osoUY
2m+3ASGq5ug43Hu+PUOcWh+DL26XWRcA3qDKdGKXfFHPSaDeTKluOVXyQhgAZ1+N
Te4Nty1q5XUQRdPCaeN1bvL13jSyFsoMWVw0yuG1quptiU070nIqD/j37/Go/DNs
5p7sPSe3CF5PuH1O3kn99j6gHtI12ZmHuhiGdZ+G4ETYQX3ceh/EE6uIZ8NDfTfw
V1VrzYk0XNTQgE1rzDUMOQUzHyplgNAzWNvaHuH+XPVEHeB3iel6ocLnrMie61mY
ToWJyEuRnNgGZHuGddSb8+muZBSmh9NKjw5pt6hh6YeakOTldgCR5oc3LFFvyLR8
o3tfVg1sQULucqprBPpzdHLJlNKzScxs+npzE1ELsoWbWgoY4tsNU+t/QgOW52jA
lfgtBboeCLLSETTyUSQFpYHlZzrJaWVnnDIO4D1E3q9+Y1wni7HCH4gro7XiE+5T
5PMgu+fbI77lfjXZRVH80hQESktaKTvqM8F75WlcHjSV/WYyS3Dbcabn0e8xr5St
9bfzncV5KdV9DeD5s4MneEJfytCHDykxmJ08zNq0qj76B74d+rkDUxOsdY905MY0
iqm43Nqhe1pyckegOpf2Fb7HDO7XHE47NoeHMyd7+nxTnk7uXQmKHU+jaDFTxPB2
SnrB59i4thYt91lcVcVvZrdPALageg79g3RGKynoLl9RRV5vNCKdEjzXFmHNki07
3jXhWOFT9CfJyTp9IwdPSKM9BtfqPrzmbMBtrJ8CW+b+vf0tEVWAAMNBG1w8e77C
+K2O1URB4wVvi5/63kPmnF4wcI5v2vxrDFxmmRy2+cCXBko4vWLbqbxO7VA1ta51
EZ9eptycHYJvt8ZeKvpp2HaXkV92iFGWrRfoqSxXcQp3FdHT1SBSimaPAMnwUX/Q
yuzzVi/5oqZP0XTsQVtN/97+PUWCknTvFEvtFs3gmY1n4Z/UW000dPLnCwcMLbki
CeAnKTWVr9mosCHdztAA72l+/mEWMuygWIJZpFmSFu5/58NC83nXFek7HwTVAppP
rvof7XMui1vuELbs/BM7wGFd7Nt6xYV+QkwtxctQkwyoFCcJPO0IMNrXZvSaheH+
ImDjWaCtw9iaFYvBT3c52Zp8zbV9LyiSk3hPoYTz76PGWw4lnHsuU671m5rjyJjj
T/9t161fcdCH7kx/tQ2+vL7IsnUXhI/ZxDymCkcJgJXnGJHecQ768Rzbh+inQjnV
lJuasoUpBC3YKTAEfIuzNtvor2LEM8uQ7P/Ej1kz6gY3rRzu/9MnGgFT9lf7TLl2
HjpY4j+lJlsXj/PF+A89cZAJc82bIvq8YkXMjesdlwya5o1TkkOYc8S7EbC/JRvM
+GnBm++yrqS1Kul3LkeTy55A3ImhKmbthypJRS6KlDpC3jsMfYdNPRi95KZiE4m0
jgdYaC24Xy+pKVh97+DbFdnDcWzDp62VzmLVUKJM8dZogUectMaIh7akmyvsAp/M
4c8TYx571JGmUKUAxCz67KYq2gyCXWG+r0kZOfGmLLJrSeYDosbBdPCDHSjbeP+L
q7vV6zA2cHtkZ35ZE23Vc9pXn/wQqW8+VtnH9i46stYv7OohYXsVq0iohbUhef3Z
z95OOTi1nMjy+2KHg5AJkZaOKvr4jvdaLLjaXc8CGxYu3OfmJgbz9ab1XynXGFky
j9vEi9c8C2DHj6iQxTinF2g+yzo8vpJAeN+N6V6nJKNr9QnpFSulkOhaRvKPuztN
+MQuleaW73RoplhpjHfdC/HT+6nf5BtPGQFWkz2+N2zBuR/nJ7dA67SWQHPhdRlR
gHMCH73wFKaekaNSEwQEEwc3JUvjC6sB5ReQ30IPw/+8HJUYINQ3qrsvr7gy7xxj
9UCu7JR6+cEgLD+coM39wXDQtAAf7kXw4Vp8J22JCR6vUjXEmGSd74dC0UKLOSZi
8tjP7sSw2Ft5aW5AqSdncxVBG8qtEx9S4/IOJ7Y9etwMYeRXrmwuMh7ggGTuKdX0
S4fkbAeLa64LxHf2IWEpz/6vlr2TDDp50gSbmP9Zc3Pb6DZ6B7+ve6IYJOFb3vQl
qfYMXlnyPli8IffkkjocUjfoaZteL9GcF9xUFxHGrXypJuUmjbD/fJn6CsZD7T+c
diCjqRr+Zdw0GaxX7HrdOZGB1YFGXnabckEIS3ckfI+Tbz5OUyAyIwpR9ma4MYJ3
hV9Jh8W8VFh7zAo1H8r9aiwUrmsXa3GfOc1gjjX87WkbCc7E39+Q9FVaEP7q5fkU
qVBFVuhu9wlD55OMUBxdTNWI46wWpHO1aq/dnCqoIYSpYVrTnzh03fF85OhrHgn4
53M6Ii0G/wHcLqK1C40m6AcqVpAv1vTknBfStCWM0G7ZMc8a+QbMOnIahq4Q1iHQ
SAHDRfUDeBQ8/4N2wSpt2DVp3v7SZC/9DdbqCWkLz0wd3UAZJwjFe1WL7u2XArPx
MvbR4EeXXguaAk4B3/kB5HPr0maKzAKY7wIOz110JdH1Z+HT82GZ9tXo90XOIxQI
jRoihQGGJ2r697WSPQm3OGMi/i91aFzjmiCcO1BMey2W05sL6Lblc0pa9lTzYOnX
QYTVhF0wRRSY/xeZZ+r98Cob+gE/geq6cvVogfCl78RLrLNBarDAzZmR3npYb47b
48VIGXJJrKVBtVqecvkKn3GBqS7qCv2ju+weqHA9M/ukn8hrOyEq/K0/X5ZaSWi9
4u6olezAL5nYcB4avrL7+4AKk8ittmgYynYsFCqs3ruQ7UaTdRo3CRfzzMK247ms
4HtJIwhXfHj3qA80EUm2+Wrfv8amcBDREVNyoYY/CpHStHjVdpg7loxyI9OfHAFY
D7WlhHsb9b3RnCSqLb0/LijQmop2cYaiju1602iH6Ax5ReI2VXDzTPqwyaM5DK4l
edxLsMhrpgQCesH5S7xGqfLmmrtvr89EnCJDmxNWmy2vo3G532LmX12fD38B2vAl
6umZOSTgzqBTmC83CY0K8UAr1AHdnAPcDj3OyCycHEkulLjtj+Qfzy9a5O6DgUJQ
k8+G02P1B3TXBhePK/mEM1qjRVvRndok0u9zBgsHNH916Y12SSwSjPUdR1HR6gUy
+aUTLu7wFI8/AuWSmukfUrho8SbrOAfoRfNablASQLVJJzXBjt2WWekSyICAzBCb
cW2b7+dB4fZrTydgZ8Tj3WLTCsO1XP6z7tUE0NqP2SK79XUxxMSBHWHoWB87hfP0
3MKfzjI5+NeeSftTWXR3nyFwyFQKXO5boA1hXqu6YSAplhodqqqtlhodKnLPM31p
rju5zpizUP81r38JeKxRiIps63ZjFbwp8kgjqUnDypeD46CK2VdXqe7n2tdLE//T
N5STjwmgWsbO83acQUekNmLUTueByil0Oxf7B9LTQFgRYkbTA7dh0dLMvLWXY8UJ
UrtdU/643A4JdvEBZYDIcKegZfOfjBOr5KosSEzimthusKMXAbkt9fMngNCvbfaP
pMAW/bHLn64Kbq+g69MJcEWaZW4vxGQ8C8+ZAIb+U/R/4afTx8iZp4b/eRxfoDYC
JT2jDo4Xr8yc/mfV/5PNBQbkIPecBjm5f/JdVPARui8AG2dFz9nuSH+wSIGWSgve
BEYmdQkLYZ3albrCwRFxvd+RxtehfoFJZKTW18nB5RAEmU7MZGY82YGl6TRLM5ON
xvzC5lF5lDmQtI7SLV5JRNG45KQG29wVsmLFKBYUmbrH/2sC6jI+3ngzORd3hh5i
kw1wpsAxXWsTrwJ4/AT2+NafoT0B76MVoChjeIB6ZJeUKewuYoJu90raPt5udCKY
+RTHMAMOAVm/NnDkgXpVJo3s8pNxWBr5c45Wku9mZUFcz2t5iQt8NqxXia5sIhuI
EpHPYSjQ0ggJy0V5OVRdMxU0eRHU0RaaRzIQ1l9fHRfsDiZ4NCD7XdmZRNyYPC93
pj3JKmMVBlCWGl8l82kS5ObjCi9OCUIibZeJz/SR+xa8yq1ZCQCnhHlM+1yscI3F
j1kkgdkMsfFVdLG595Pmak9oEx85J+70cD8SFhUjGy7ZOR1VASPvIwufxyFw2RVC
a8lo594xHNqM6eYxPNNxkw/MA70CzeUD+9oIlC2tmNgysHyJa2cId3BrcVwkK/PP
avrNk+1d5z+rDfwXlCvsjMqd0ljjUi3m24C8C9h3a0MMMhsc96rRLM/3eOLz9kS3
FBWfF8AE03YfWoJV5+mHqHhDyhXEd342s7Qjmr8zsGMJvEeJ5RgSrwaDW1DS/Rl9
rD6TE6I5TRqswsHfrWc88Od8I5enn0yX63XaAvae3QrfSfBa5O9fKr5stROkTvCG
cpq+gn9sB11bC+1j4SEefNKMRPT9esruBDvL2j2hMDAyEh/CguzzyIaRpPhSFtHE
0Fi7hSAuhjbPZnvuR83sj/DksiRXzMQvwgef57aY4+FJDKaSfzx9U1WcEHKk2diX
2u7gmWnE8ZxCDy4d6SbStIJRiF7yGsP/zjpOyJlT84G8K27EzOuRzo/d5NjXOU6T
0FOJg/z8Cql/MB8+/1urwYXjVENKZYf5cwgQJwkQeSm2mfsKArZuGBd5gv4G7aXU
3oMMx5EcQUHVwFZlClCCp7ynrR32MMelK9CH/naMiQXbmYioehS1M0eKBj08/xDD
WWO8Rlak9Ztj1kO+fMYC270rXCjkzVnWxtO5VU3X85ndjiaumj5ab0irhmmCX89u
4ZOlN874VVimcMdF2qjbOWpNSJQGv1VGEPCsf2xnN2PO6P3xXYs/YvYZr39XD02R
G56jKTmG3kayWk043W+vaQqoz0ntzHJ4/tMb8Fx2h2urj291o6SRFdt7DLwH/egD
R7FhkJd1+ZszGM1qUBrAnjGuOlbIKh+gtIbJ1UXrsSLDciZyM1pps5Yrq962NI8c
eEv61DhRS0Beojdb3/ZMXDkpSCCVOU5WkPjCTnVYnLPjNo6CouF8P9boSFxCbzB0
kLHLetwQPccdXEHCwprL9zvrSnnlKQjFlP1SFz1/4y0CnLqkUjcfBTcMOAG0Z6tA
wcG7MvjsDiOOqCFMLUc8Lq4hTNrOXBHMz8IUBsf7EjN/c1zxfTB2uwjd/eE69SKn
x+sJwwhjANDoykUny9usNQ5SlPLFjDuIr7iCfdcDur1bZ/WR7MT0uUSjIS15P316
SnjPDKYuNDwHVXysC3FlBmtqtce3Iap2tLzoMGukWysIcQTZglgJy0NTsb2RaweP
RTa6TR5mIDHtjRHIlA41AWgvgMgY7l6WM3F4OUhYoRF6ljC3wx+veZfrV+D8DZ9s
5Uq4HMjhAjt+Xs/4x192ciToPJdmQ8WbToPw9iyj2x3eUdgccV+zaknTrI9ecNfY
Q9BpkxAKwweZbayeF0oI0nJUwhLSE/5qpOuf1DcDJGvuapMO6s2K7GZ0Dj3PIy1u
wE2KhSMulsCC1hxLF1qnGc0kjIA+kFYk+b/LA1PVNW/VAIm07aZBlj7ORcWTaKeR
lIDK0XXAW3wIoEk5VBxnqlt8BnYDCdRDj5g+Nwz2+Bxg6rLp2nDULC1w4NgUtX7S
5cHSFJxnVWUfSctvKl+y6SsF0+VVgtxB5Vjbqh1s9bsx/8Up2nsxrcEGjujd7fly
dh4RXIqsGtK8GVTKaGCjRPu0SOJahtoS9rEz9sBCEyV0iy6uuyGI9NNZiUy5wU8g
A3xTibN5eQEEN8EpmkOW+UC1KX30MzR7gRVRr7NHF/QrnmmX3cZQkrTEkAfkfBaQ
YVUhBVfyPhylk4xMLyvdPsc5Ouy1+ec8LzlggjAVO5IBpgIC1QoMr3BO6rVI4lHF
bPO8Z95vWHPqfEC9jummLy807UPIXBZ1Y9izo8c0FcIkyV9EltmrmR4bCuksuAYP
FCo5Fo/2qplWn2ZUlmfrNcAxtofYY+FCpvGkTmDwMjZlbQ3ju4AjxFUasuisvOSi
gQ3nGiR2ByCltgXsYz2Ypw1II6Nd2oRKSXDlejkGkHShfE6P0SXY8vcasEl7MMUI
uwMs4Ki7hxcK/y+NqoXhFHjUJR3dkx73VMs0My4sAT14iOaJIczpuRRvfoyL9IKl
0g1dur1HsP/PaVgzE/mQ0MZv0egFk+ORPSoKMfjOwl6jDXOkFvsxvlJ7nlGRDs16
FCG1/Vj3/2h/i4XJ2OPEWvAvgTAPIF4wkCNYttOJZoOJezARSwSXQjTe38FxFwPc
H0nt2j6OpJqVHTMFwroreAb6ihaqNQjZleyYY4uYjwNEeNYd8Dh03hfEtHKxYQ7I
hgeSMGpiZR1XZbu7CSDNbwBJKNS9RvaJawoptntb/S/vMfdZci6o1FZXCNU4cd5i
d1C0uXphPCUS/3SrPebPGwPZ+ylN4J1+J9PhST57KoQFTf/JJuTvkiK0SxAXPjnN
N8wVUNz2aVNNW2OUifbB9V9U8ZbUGa97DyPJfvrddSPB8W0hjwDOknqRM6Nm7NRl
HotlZMdPULq1T8ZHvspDu6mnKFGl1WJUoGj8DywHVyuAYLChFtM4dYo+3pi+2g9p
ViUj8dwIZSQhLxkfLW/213SHSeuRX2AYT8RIq931RlxBLvyH1oLJbwGA62aRBL0S
oi4S4wRpsGsENx2YsfTp0iHghPEb5PjycoYhHxoQR0U6+7RARYNTmiXScIrUaZtI
Hlvf2px1rKbPkEzau/FzugtQIM7wOzPl0ebFOVWKIRl55AdRdQa038hD/ygyuobv
idMjmjXgGOUcNQrz7jTUgUOKD6ZeF3mkhDYWRQV6sYZprc8nW5WT5/ob0LztQyQC
kFFuH+zNvUUvRTP3dLlxzpzxU5wDA8YB+XowuX4BRD0rh9lo/nAx/6PZbZLkN9Yl
u62iQb/awz76rn2pEfT5GinJqZ1lhFx5qCIfMsWp/cTPYgO/bEAlexH/yAMUZ9+5
ypjvf6uTNoC622FbrHiHXQbZjjPkKSYBkt7uGhUvfeZMCGAtd6Fm9OAKdSfxvEKl
XPOIn2Oy+LP9stfvmb7CQHzDO7cEJONSjlzoQudAGcuUWLF3aO+VWTag/jn51yxM
GXdRlyr2bO6DSgsCWmJyQKwHwEgTXl01xjsUbLvNWMs4WuKAYJZwhU2skAhhtgWm
tYlV7QJhJ7Bshi0uemFpme7jRm2DtwoZBjIsD4L97ZzJXVxxOWnKGR7ms058K2ye
OFStwQBMkPyvYl6+0uUQ+pHaqeY3S+PjRy11GN9M+kOZqbt6YN/RY980mWvp4MDu
FPSgNzsK/70aXAktCG6i6KRy5Fk048aKEEpjdUqcUNLuZadTfN/83wa0lA5MDITv
qc+hwZJbjI5M0tjOfdptvGO7VQucNQfKA29yDhKombuHkXUZYWsbqvQdWji62+oL
s4l7y10YfcK4eAF1nVI2ezexKKxKYeSZCxUFs0EPEkeH5VTCg84otHavEFqMPY5B
OSucpz8nHnRRYcL9+kGvhloG0fUmPDkoAEIaRzWg7lBZ1eu/s8PR3fboIzvEioB/
tKbN2oJqPEJtVYzPXinVYHzKY+CO/R6p/st6WtzTFfRrUR5K4DBhAiMsHX4uMugF
msFpep/ren+v6NflGmspUU1bLzkyyypnQ0Hl/3abCPwtvNhizjB+zy+5O1GOgK/B
IZylPmqbP7Ai8Y9KC4dLtFTkusHGjMhRHOPsofPdU0ezeHTS2W5LBNmfpSEilij7
vAG8MWmroDMDqoGTrrkEjOHw2OpiVSPlrja+V8vsuI9RRKIEyZvNbzLMHkmZkK6H
2Iwwfmr53PrAb3m1+ciBVbvNMXIGnugItOrMErMtpGCZnifWByPEVsfdo/BG6JMa
nrSkgsHRB+r+cHi1tytIrKMQtM1nMa5XQx4wPHgY5qgYHw3XqXesOCK13KKiSWSs
ag3gCoRgQCs6EvymBt+zwTzBCjDyUnRZadAJ33bIunIHCv6+BijY3PVWiB2d+8Hd
X7vBtgNJy7gP+1amZXD1UVVrafoX9HGcMkFI2yA3tUrVvPd1fyRyAoEuWq14anD4
7ibdQeeY3fp/gQBRlvfmQ2l8txyHplqISVn+RsjQRbcxzjAQiMOUW97SFkpfnq7O
t4OypAWxvIqTqWn+CNCoWoS/buLnAjW0/E7qJMy2RwicMkInkqCaIhOO0FgxE1BJ
fJgapqfI6C5tGVa329Xpn013NmErGuKySrmqEBp7eEFKll166dZf8n24YTd9SglT
p8j0loEkorVn679ug0Tj/W6ZxO/h2nuqTB3gkALsCUwDmZ3XlLfzQsbBgwKmeg16
pzbWIr3WZ2Z9CKqlm5wz+LsrIpkhNrh3uHwVvZLwJ5lnQqT6yKVyhLzjRAJ8WzoY
d2fZQCUrpF8s3YmxY2M/hua051Ne4ef91ORdF6LEC7ikPbAUoZ2zBbswqIiWCnzy
L/nf7Bu/RzGdA/PeNtjGhZvNEsj3uBM7Jbf1uxKXCfEauIZwhjgPSgLOLODjVRqG
bSG+dmiKsFsgssm/EUzunxtURnxYTFUjkKPu2FzyTm+tQMslpAG8w1nhe6gIDoNH
bIASwu/idXWhoJz4xJLi/GX42eZ71cFcAoVxHCa6KaO/l7Vmult7bST5t1p+Ubma
3rI4sMiNnTbVw8QdMUOy45254HFWUaX+e8TgQD/sOXJ3SfqmiHqVtnE34XyUYYUZ
hlWeku7CYCEefaImn96puUwHjP1cc4vWVi7LSTlJwpfEP3ufPZlUn+z6ygOp1HOn
CfBOK31bavSbhrUUeXF4liqXMeW4dN1TEbNNqwrKHfgtKmuI8cIgLg1AabT0hmEg
MhYKdV+WeblIhN0wmFFp3yoRQUAcEPxuyCzySt1GJ3HaTrREPP0eSbn4dsAYvO8H
47DfgxLbrNpy1fWPR33CkBpOdiKT/Ww0sQmWuDiTiX/PdeaS9F6+Hur67Kk45rE3
uBjMmOimgU0Mzz179jGrseVZUDbvw/BBoK9B5RL2N88s5gDxGoaBwj32XSq5Xx2C
bt6Nlfs3TfGSx9UHlFgkva9IyBEGLXgD46nelIRnrOLHzkblUfxQc2xA4nM0rcHL
O9Lbs/f4TQe1M6MkYFV+77T8Yl4CAn6t2BBHFJtbPSGe37P7SCKicstLn076WFkL
S1cNbRHAgdKLDISq2/KsYNEhqHbQ2t4dGm78vvuNYw2GY2SHdQiF7DIYX3qP8tVt
KLRSjPvXqRXQtytfpLd4j79OJHZVefK8mLiL0LuWUcQVQw1cwGgnAkNedvvIQOOs
WTWkjYpz13n7pa2ZkojAuCLliwgKhFsjqhKgBAV0Dj6DX8ABPIEcsUvl1l+CWUwh
GsV1qPE3R1wgRByoa0TB46UbVHo3tLRxtfSzAOrf9fSEAVzbutgCTl7jIWf5T+0k
i+uLg2UnhD4ePAuxsP2uhHisAAxCCFOyD3g+082q8NIAQP99YMSsGSR+fEoaebYm
s5Fy4GIsk4055Hn5CFYRCX+fE5mA3tOA+Av8AoDBI7xcDWGdFV8RRmg2g9h9Lkll
s8UMEtWXPvfGYN+btTS0hveB4v+Hd46/fXkqlznrMbeT2RXYEcTXqrK2vR1GGnfR
mFMEv/cUPA4C1sv4nhc1ymAnCGH8PUsUL5yVgWXVoc3IV/pjZeF/8GS2iHAgh2HZ
x36MlfaOFiif743w7uGlEa4vG/zFd4rXR/Iw+H8xI16qS92bwfL9l4tpbVOAtUIP
bzrxp+sBecZcd2NRLue0tihhwyiGzPcD7xw+8dSUPuZjkUX+jf7VAeyEOcd/cx+U
jRC8ap32MXaNlL3GQSyvl9wN2DNv2U1vqLjSRkTO/aKwnUrHCw6dp11wIVp2h1C4
rekFxp5+B+iMFkasvvqQM7X5+V+mzTCgsRIQZHD03EHLc30MTX8VeSQgWUCmL5Vm
1IbLpzi1rNEkmyzsLk9BVOhsGbf4dUq0Hrokmij479gW7HhdZ9urlV52NUXorJMN
xiqkVJGAs3XbRKfi26ykzYXmNc+8DqbbikIsw5J8yBOeeg+FKpr/MeK7grxGv3Yk
STo4yWGpoz9Bzkkc0GEXhMHJKjZa8N5dYDnYJNfv66ZChgDGSTccppdiMeLU+Wyn
yrW58EsyqQ0Uk/jjWyc0wC5qRqTa7nzTavsUyVkmM1Cmt7UjmesIJmHHbsffHAmy
Dx3mhk9uSAMrZcpgDF0yk7iAVGEUT6+XmWAPDxoiUPBDa/umE09NM0H6wlBsB0Bk
Y7CTOjBHSWTm+8SfXnxsPqprquJX5VyK7ArtRwFRquaPDu3/kth8P1M+7KwLX20t
1oV1AwR0xmq0KuNQ1lo16Uci0SC99iBSKB7BF2eCYt2HxUyKMQaupLLu5wKqTqqa
kNwb+444w/TKn3U0BHpB2IIuhC1EqfXyl4p4aos0CCsPlQL9I6HRSxew5fyAmvJi
xa7vA3xteAW3HTSAlf8+KXDjcLuy6ueaoSwCEXQGYt3V++graVquRPlhifXCJrU/
Rh4hePgyzN7gQamzTqvqmMmgaNRQvdIzCMqvEualKPpPDRC0Z9aVlJ3tXZrk6Rum
cFyWxUfWlo5KjoXMSIBWrJ78Rgod4TIOUS3pwi6G3gc5S/Vqu9ZyjvstggeTXKeR
2/VJPVopqYgvZzRviuRDAGpdotx0jBhorBzeWcC/YlcJjDkskZj0U0Ll0o69mMDh
N2Z1JhiXh1m671PHpInVJnb678QvjMLt6cUnfhCEDUNUrwmtz4G0KrybrH83gxW/
h0ZggKjOojWwoyyK72I3u2iUBjpse5WVQv8ib0NqvQhy02oQPLhKnDgdq0Tcf0Ar
l/356tpojXf570GcGFyOgPseNgi9KzSyNmCE+p9IQ30uY6NubayZ58lfvxPQ0KFc
wmFYAa8R7sErqY9sN5cigZQDo2OXqb46cMuJOMKSskpG+PF9hYymd00GZtbh0/yg
TO8CNb3l3HQy2ETKcSsxayQYRJ93fDouVX/SJQhFwvWOnQ+t2eyo2qaIlSJONAdL
ggQP+2fTDdRpj9gn3yNPhUxMX/Y3ewskCuQY3LpDymnlka5r04fe9V+2nu1koQ1f
6SwdI5Gus5f5t4yatrUnQOjOPsSjLhHml87B8d9DzjBFhbKVpS7Dr5dopjAxq/rS
b+ECE2dGFT89XMdN2EU8gX3gWGdcYvnX0t7JpnNUouiS6AffdzpazPa/z14pYIpv
tMOVzvJD07aMTiSJAjVVkrQUpHe0kxHilwwweShtoXQst6XH30cuqOhrxPEwdxZo
7xjsdVVkvQRtwL0aODMaxUWYOr5HjDcOnGLGE6+2zUA9jleLK2AzVLq3KYnrOPGY
4Fb8cDTY1Gb8HEdd0MFdywQYtFN0BgM3T9hUr9Nr25CeDcoR/gB+XIgGpTK/VTwE
Pfl9Lb/nCCwCf8OySKdLKDXACr8ox5/jlJTqkelnv1+7eP9cv5AJlj5eXoxkga/O
4795EHESwD0GR1R3lla6WZF2/Slsio0njshd+A1f2FAVfSM2b4xmMF/DLn4klzee
kYdq1Euj/hAYomHNpVKiZX2h5pva4A6Aumnd0OmDUQAWlNXrykOeRMAKnLqb2Rq9
l3ow3l/w9WWRWEIz8Rq9wpTzQkffaRiLO68q9IFMbzC9bB2ufkNepafClgmjWYfB
MkuwhQMXOOdPur+GbW7tOAhhcPdlmaB/E8Ztu741pkH/p+VZDg23oFqlG87RkmPB
SlEqr2HADTezdGA6b6CRzHSb6+bzD23SxxaXyA7huA+ospz85pxtAAgYNrD2WQFr
H53pJ/hxoheRqJKVr0stKqDQDBR8FsQ3gws9tIknBE2oMZRCwiOk7hAr7EbThzDt
R7YBCpvlPkvWbo6KslkrnSjEWIDUjikvG78fAppaeqKBVBElU2vhbUOiBBo6i1fX
Hx/xJ3N9sAWTXN3q1Y+w6jOaVE3jnRKDTfvV6v91wauPULbEbjGK/3H1S+eZniJ/
ca0ambVNrcmy8vH+X7EXVxypDQx/ZcJQsoFkVIf9oP1A8zlpTSg6xl9CPTB1TpM/
PxtCPZ1OpxS+OtCH5pRvzuQwxz+HZz9xjeyH+8rzDuDiebUJ/Yg0B24lIbgEcD07
f+RCReJxKUfuKeBpQDvI3sU/VSr0fcN4xL70aSV8uQsppyDTO2iHASZ68uge2yBI
ATC8w3s8OLMoNTXncTYTm8emhCMk0crW00yY24rslBwUcs03ckcSVZmJ2i9Py1aD
aMzz8Z+VyFheWjpVbfyRFMwFWdLDRmEgrhWQRGjaVk+coOh0X2h8EFnKeDT4maJ+
cE0mVEY/xjMVIm4KyEptg79CBtsw5KkMo5WWF7MK58KdLc9eCnVYvNn197tL6I8b
j9TKed2Hk6D9fSRZZ0ePqcvwDQ21Y0rvwNSgQl07VhaDillHXNEL+yguVZuEjpIv
oZbc0D8ZetAAAUvB4Z5sduKxMdxUjbzKV9TR8Mnza4xdWm7qTyG25idAZx93SMwX
5ssvofS1IqE+3hL6XyXT02QqQBluRXinYuGEqmOCenKy0+FleDPNiv5OaLAMC14O
MPmPRkv5wFydCMDu/dbMosvaWn86LKzrgX+jqLW4wC/uYggfXpveZGgdDFhy6ww/
cY4okHa8yuxElSl71FFaaUl5Zn2mLADvPVgGQKibco4axE+XZC60MzMi+lKg+yIJ
0kh28HYqpHEQP5cZvSQHWNDZ1acHDg8psfnVdtRomD0nEitaqOWURJWCesxils53
L9NjS50qhl2a0wIQInuhWLHJUeoSyIFiz9ymm1Ru5rgmGIai041VvuqGd/r7Akcj
RxM6slvI5edLyiOCquFz+RWnHBhrfPrsEMap4NHyf9ZNZEsNotrjjTdVslUEXlGo
icIjdh/uStLi1ta5JwLnhN3QVqxmDyVeXucyQx8bqNYzRX844WYG7kgNjB/QsdD3
zuIEW75idx28hbu5lPaj5piWtyTItN7ftVQIbaKtQPm3AbbVwQO5Qu7HRlIlNyql
ZjCkhoOLQck48Co85dgalAC5lxWdJhMHzDin+M6Gp/fHgLN7WYRQeG+wXRG0SgSO
LNH8M3EwJM3cHi9H+iq+TBwTDCPOHoIUFkic8NqdG8AlbUqPTdTDzpDWlsELsCY9
qc+NkMTgkwadJFV2x1gzdXP1z1CJpeo0kpzEYU7ykwAcIDRyBPMdmlJtxtX3+Ago
MD3Q6mt4FH8hKXS8oiVVcUMHdts38icfGF8u3MbDb7X/UVlYeSEyIVFxAecOw+y7
zxQbCr5KmN5Li4hvsmi6sxvhjcGnRjRpKhR+OR0QdigHw0e74fUY+I6zRheZ3UYq
iN0/jQ/cKd6xjVqipyCpGPGIdCTn5CUlf8i8A/Dy+UCTYqB1Dpqnr01ZzeyZ9498
EtggtD3JbidQbxrjX+ngXZzsOSRa5ezGDdDCS69XfxdYRkwfxOkTXUhbRxo8VeR0
WF2DOinkAOIU8oo12oApBJQ2LpuDt3zcPapI/jEnbL4MT1T7jpvpZSCis6JANIZe
t+njEr4dEElqbxwFhsr/bw2uS9+qdIroBmi9vf6wFWT0zA0CtXrwECLB/jMXviNd
dcq7JHiOUrexFccRwnAHmqjZ37odL6tp7Lqit94wu1Cpenprg2qBdCm/+GN/R6X7
yDJ8gLcuQSWbO2gb2HyWf3unIN6ikCp6i/PmmofjRCpjDkwD/sRi0wZqJQBG5QH7
XU2umR5UEYPUmDz2C5RpYKArNiXkiYfGAFGHZ2mN/aocT3OBhob7pEsPfUiwTKoa
EiuUwmY+QdOX1muhx9dI0HrP5TvMYTM6v4+mr1K/S94kCLh2zfL1U9YQ+4Z92P+P
28Z8aSPsQ2qDgzYlwBGBlFXs+efiGb4U0P/Vn+8t8YWOnTjDvS5MYnGn301N4Kmx
/Wp2oVGSeehjhn4G6V29UXok1xlrJ6O3HgTA7iEakWgRRQd492xcgZJSHrHTrY7I
4bf9HcBmqvfyRdkWHumjMxSgCWrhh1+yP0ly474R1eAmv7KH76cY9xSlFLoCjNDj
nNWrdqo8yqFPlXzmfbM/6LNCKJLtjwQ6kzfZ7Do+HC8y0vB60wVBvZFp4Lt5hwE0
UPU43a/CrIWOaJJDNLrUxHLMSTvO2PYmiNXwkw6JlY9loEOZc37lrRAq3uqSl1nG
Hl+3ar/EdxCN38KBSqEP3d5XZWrcdw+A7yEt6WbrzKpL6b7ZeCDSgXMlvdjIfM6A
ithkWgjs8z9pjywJeP3Y1YZBmO4y2jQSAm9n+mLO+GRkqvPdVXUfIwww6eSFw+2z
5n7PkLf/l60u+3V7HaGWv2TcPiDkK/r0BuY+CNftVrd8q6BEJh7vC+UqaiiP2yQE
qYdRQvIB7zsyVUf81I1tddBUlgVhcT5NYBZ9qG19jAQ9RqeIXhXVcFZOSF0IegbD
BV4GR4/WKsu2BxrDn0it1WE5/gcvvwLXUNF2LPCEi09m5ZJSwk8NisU7/Yl9mxUZ
4WUGCllL31JGMu7YwUqAT6XsMvhBEe5ONvSqR/0DZrGnyUQlmjee3wTSEYtnLlm5
iBoc02XzAHgP+0rXK5IXQBUipMax5yRwMo9jcLfYY4/zlQXgow6FqIzMzOav1fCb
bTbGEM4Y5cNiBU6xO7IrJ9JmI+qhV61zJaUL3JNhfv1meIAS35V4JeTZL1qiAevA
Y4Ep+CNBGDQjCAIMLYBFLs57smdJpHkZRDN/WC2QCY3G/iWynHv9Ps9+QEPyFnFb
Y7NYu/80lhO35egxkRLVf0jTdZOlkaEkxgOguLwOdO21gEoEzekk+RaEqiIIroXI
BlebC/VL26c1Hp9+aFDClpsPZvSVgNB5tolqDUop195Zh1ckjk0msnniN6HDpPWq
T6Iy0LBpi4RNgX1l4ApXMBvy7EkWw7GTpmg3xNAV+qP3zqFufQdV8ZT2nr00rZxM
omlNhb6IMHz2v4JkbL372gAZLr7pXmZarLGq7VC3HoWyRADwrAxSFnQfpLOpnjjc
SZdY+nivShd+Nfrb0gDDvsGSjaHDsCkW3jwg5jRC9uVkT6/0/T5BuUllNYRqC4w6
R3V2vRogLLki/TWErXBR/xbaUBwAD22prA99GKXaU1A+ktBvHkO0wskY8GIjhSuy
OlCI6grF+onqUJP4boaWErTwoVEPlhLFfl+r80sbacTKLhcEVl5xeBmMwCw74VPM
F/sUbS40zXcIlLBukqytRF4s7CBio0cF1cLa6+3ugSEo9K/0E6mZ/7fefwok9Oda
C2nwXvmmdB3fnOwBrfolzpfWfyw5K5kKyvXFU+ibmbNyOeddKhDBfZFUonZMDVkN
kqWCse3V97aINF3T7iyFBHgxRLNdd75Fc+Wi/OnpvF+tO/Pv2aZTNMSzMSUI/whE
QJalcqFHt6u9lTSkk559IxG8Voa/lv5sTJOkHGgYDxCaeslVD6FmoCA0/p8DX4l3
hYbYBTZ4NgQmfGZr3PiBQawDDAu4QwTSHYwZbUGscIhhuK40t7XwOPyYPlCHOs6b
TzHj8AusGlNg7rASqgzbTFOY+CbCWWdLGKt9rSo/2I2qcF2Zq2cWC1XjAarJQ4yq
WBZXMSZCnhVxUp0Cab2GEy9JbhPsgVi5eGvg8onwSm0NqFgNofN//VdMLYDknbej
E4FJp8Wn6pioW2L/VDXlIeYBRCG6lAVeUg2spiBlM1/26lsochRkwTn0oMGQIMi4
yfVlibKmrY1D61qMhcKvBsmTxM7zEpCbqBf1FniuJfCN+h4QbWr8/zHniAbl2E47
Iojs9LkcXhuBhsqPF+oZ7FbmbhfsYxb6sHUedx31yJVZczxEIWvSsA0FcnX7KSmE
siOXbdsmAgMEn6ORJNc9RTiNeEX5VvQ5aSY8/Nveb721l2k7t9b3wChWXdDrkSx8
FXdWDzB3Q2v+JcNuzgYpnWvKTacp3sKhzhtsEWZLhIyDyA6QyYcDJIxUTtrgQFlE
mqBvNMozLOBnm2UlpM8AQNV6EUM1atSQFAHZwVdPT5hKnegb7bEHR6KNOx9OGIXE
Xc+xmbiHCkx/LAmwmVYGzAkaWoVeXf2o0nT0Vfxb/0Luc//WkMZ6o1dPHWFBvkXn
8JCIlsnmNS5+a3g8Qlj6hSaY1FFnRXJLPqZkA/tgjl7Uw/7Qp7m1CDM+0YXCusW5
YwJ5nhEv+NyHdXlb8Vf7Kho4YObxYfhRsoI11lLL2i6A4LnAf/i7OSTeB/0vCGoY
qi9OICLdMv8hyp+HWTPjOyMXrXi8RBfduG70bdwUM4Ipu60kkbjCcMDY9uA0qM99
YD8M9k/Wa2NNYNkS1I57+6PQeW5S3M5KCsJyPhXLYsP5NtUZn1wkhzGOHmtdxND+
+owrrURbfxyHdhdCmtYwVSIKvH7fdzHLDb+/Vs6XXthBMORT6nE/3/vl8gCRLd8D
xZDjUolcXCizjiTOeVf1xc6neLBHuhHBfjqACU/+eq7ZkFHP9BU+am9UWV0FRE3w
tXtTrH0lCLzksXu+IrM6GHYUSQ92vyvP5uGCKofV5HdF+pY1fU3xGc6M/dx6uaG9
0ZiEF6cgM8GnXHY3h8z/VB+f8xTErEgeVLHeYx4TkA0h7KP2+mr0tf1+MJSX2wPA
Fdvwuhi1AVZ9y+wLfwzZYT/obMkMxtcK/9UFWFkfNPJiWDmnSwEEAWGxSsOnbmob
ZwZP24SxJM1IMwoGhpDw2L4ucXxLusGWzdQk6Czx3ecAqfyARqUbFhEYdxJItKRr
4Sk0EaEGwp0+i28QG4JevYamQmTakvvzrDrTok1CuuN/6zgAfSVZ1wiN2Zb6+9T5
/pdl8CrHKgxfBChK8Ktuh7k1t8YIKPycKOuGgAhx09fJBGvB3xl1FXFj4R3VjnYU
zmWl7qvMEpPq1V/cejD8brwMvNI+THcKH2Sguq7WYIqrPBZe5LO7mzEh2WYG5f8D
l36ErIIItbqvSia2zxi6wguC6ms6K8KoIHEXGgVebBUNS03EBmCI1CmjiMuBqi12
1FamSi0QSLiGHhvavmj+1jEhscjYElymBpi7kSpmGQ/QTe4vT5nOmKi2BonjW9Ns
+l7zvQGHCc9lgzmMN+4zO4lviSopc9mYV1odStHnt4Gy9N9lpop+/mn7OS82J1mr
Mv7hikVV7HyO51tiu/YcVhUrNBdzk1daI9N7Gk2JkwBdIPUuNwGNXToUStTT/1PG
rAr6/023c2gHCiA0Q0p0Yjp9KuOrBp6TNP5uyGU/P12qeM6m0mFr22imHDZ7Y8lQ
WJafApsQfxBBhsrjx116wuJKAJlSMF8vGqra10i3Y8W5Bu4Eof5fTxKxh4Emd7se
ElkZ+vW8HeaXpXcn5VaO3UrrnF+4Aj9ZlIIcA7xSISAvZtan8daKnzauC8VUCKjR
nKb1HJcK5tiO5RInN9lJ/a3M4zsUTbaCLruyLDE/U99C88Y2EZfBF6JBgBERtV4X
QYsxjnopk8T02RUYU+DW84GdBlExGYPoDqrlImQVdAPdmCoycIwgpuOM0JPJtz+d
yd2mOQtykZ8BQPsF55zQ9+VQM3p9T1JixgUkD/gTyx7yTANmozu6pR3M4ARTmaU/
Y1Wg5cvtasKODMnHIvW/tg2NziLhMuRsMu7D12tRfE8FuvB64qkWgfITqHKvNLQy
ruPE8OV0iDEHmG621UCgfFhbRY+osNw+mUID/m3kDIITKy1n4YpTuCiUziOzsoTO
PNwK/bl7PVX1gNXA49vnW8y8NVkLujaTv3XdDt6iwCrr8va+fdJJPXTGwnpQu17K
2k6YvPES8+behavoGUZCJX2IrukW+2TtyeV/o35ARbx9JPVNp8mcmZ/HSbFdqO1l
4G/sfuz98pc0EqrG07h7pJYFJi0zZVa+wS1MV0MsvAYnsgkBU+GuOXWHVW5OI5SD
YWx2fCR6q7ZlqOwA5o1wGUHydDnKG88XnkNT3xFJBRFrGfeFn1qWhp0LGbOH+KWT
K6FRhGkY4wQ3JgEYvOeK82NOjynmXpC5PhbBfEJdFQBMAQ8B5mbld8Us3AWuKppU
PV9YkS/2iXKsHigBHmUYxDkyWW4fhI5A9PDM4u2gjUxvaKhV/iIvGDFNGi8zxmgC
wH+7PvIU78BPPNaklwz7oDyy4B56gm+DhneSi78TJJ0Z3LBmCd7hVZjcw0su0oJZ
1XjdRr5F/ys/zCPQnZfzMPiMrbyEvvD2HGl3eMMCT9D9dPCwqRNgXqYV4Z86Qg20
QGpFRAwaBykripJLVCDy6KcX2RKGOC98++NG9wsQmRQOK2CeVrdlbTXNu9wwhmas
P2STcG5Wpf2zaXh8NzFcs3Wcd0tNbYR7YkgbGcRGfAwQab7GJ1DyaWR85ywCByQe
Y3oDPMmlnu4yI8ys6rkG2I7ZBEkRNtynlQvSq5YMu5U7qRgvirhsr2F8JugKXqst
fNyoLpLLKUeHt/DO6+xXetamOZd4nTByYbQFdrbUxDVD8E4EwybCac2LDFysChxd
zGVwKX4bJC2FidpancPYgX2kUxNoSYWISFWJBKdDG3krKdgHru15sk3CscjW19yG
xCiWFI7nXTLYHTUA+Y5LCA/JFrA02TEP3HETKd6cadDZ9oOI6mW1xdvgLJl3mLcr
WafhLdIg5ouOoeX7dL2uEUWn1tz6s+8rSh7iahggvYRd0WDuDlQHHuNozrZ2hz8Z
WITP8jPEdUnTLhVBkHdzTi/qxJWTMs18/TJuWJPaEWQJNwePwQN09n34GRJ5AFGm
GHjmMiC+ZuMEwK/nqXCE7qAjFVJnfI32X3bM1Va9AqSSpxMT8TNwKZJInnPXHftZ
MfG2a3SJYF0RUEFT9zVS0U/iKTAIVX2nzik50Bz5AM4QF59Ww9tNroNgq513rDzV
og66iN3lVJ8dPKon4v2vMRksEBG8XcjCaRxG8gA17a4YdmluOGRiLHGQAfJrjQ6p
E9l9iZJVQp32G8j4hGIVI1vZQJ+Wu6eQOBZATXRiWG/IreXCLQ9bEw2dFOnP2Vnt
Kx2coyradBvwlEtvsriwjCLPRXGweOSyXAtu2tpVwBH80Y4ZANrepqCujlMz1BSz
Czeih4dbKCUc6RaZvUzqRDyJewXycfFv+37gSLBQyj6eYLPJBLpfWTPozSO/CJVU
UlHGM2dPyZtZPywoyQi6Rz0AB9h+IINfwag5xI9jPmI6HfmSpzx/6zrC/27UpEG5
P541RDiH8n7gkVU+1I6rwkzMNn5/mNF6gHI89P4yCd3kcNAYEw1jfkDkSXkX+GTA
5JV4qmQsCTB97y1NduX/OgDpchYTCG88kDRH2myRsGlGkUOy7xItyceUMMtWeptK
vweJImpiE6TYaPBuTBM3roRPbzEtn/omNaQiK+nDBCDBllHvzPbRUoMiu+FJsndd
4fVPDk5WKnUpPyJeyesELHQUQxhiW/JOTpgVMVHJZxI4/lVn13nWgj2zaW++cALT
Ip45DzlYbPe97kob1UazBSTEi4llrWvUhmaPLNQx1ltVxLvlL+4/UVIxO+gYFiZN
2C0cqK3CffQXnK1jsSB4A2n4ecdrXC7+ThKN/Gop31CxxouhBDZhqa7nqP188jNz
Ch8ln2j9h2xKNutRz9Mf2H7YD1cgLabfkaCoY9ikkcHSUFvmT7OtZN2GbMTFEQbS
aD1IDtliCkK98cSeuUoG2oxSGhtHv+LlSjWKUp8OzBUbWooPmk/52s+vYG/blnkB
ziCcbz5cSxtaVkQwGhBRK7QZGJS465M6TUvrTwIV9Jv3inN2Be0DYYd8RS+IOW5L
QCSy1VTNpSQM3YAPMz2NZOnq3g2mnlTfSw5WzJkmq2D4FjLUtLPbVKfTOVhEo2E6
KKnue/dm1owS+/UsM2mXQWwgok/OZdrMishEtKwP29n1vkJCUGqhLTgF+s+bvbcd
OY9DSX0T8PKZpq/6k9spWTbGFIxnnfP5QA+2NXN5unZlEHDfmDhBHkFgUicD0pI1
SlPNeTcc/IGzkhffPv/kkMAlzVZi0pPX3hTNGlvqbDR4PECr05KZTgtUQpaXpafr
YVwVc56eg3pyTgiwcIRnSB3RN+v8a+pRdMENkHd3hX9U/8y8Gup0fWTNGYhfSxvY
3ryzBSm2A0B9onkFWJDEmrvOQce0NuqDDMOteO/ayrCju1Yrn0GNcINRj/8/4msN
cSvCfw9dRzdiEYXXXdwQW20M98gRCSdadfxuZGTPIrJONByJhploM19IJPeCd38s
Hga0Ti2vkHxBQOSD40A3pyNCtVTDVqvhc9/YrzHJQ0SNMahnszOiE4AihabyBxQh
uRxaljf14HBMblWo0Sea/xFQ7jLam7nbty9m2KE5RjK8Luyip81hRVol0G6mDpp/
Z84N+UFIk3vjGAeQ8JPsH7vqzz4ARx0+MqmJzotxPpObjmndQLPGtenR5sEea268
REu/ms+DHrWINqJWroHZkTFiAQIUCVWTUuLYgyoHr/JNkzELGmuxISRj4k7vasMZ
jLrFu0eMr2bcXbINXuJNiIKR8Z77nlulfETdpH4hCgiH/7hoWjKiMe/dJ8St580d
acDSVXk9W0S7yN7yeOjuy7hLo3t8igHAvAhASkBcF+/FddkUX9G6B4YlFdEk4V5m
+g8s+m0sKVm5powbrLgqyt18Vqd3Y4OElJiJ8vYo0LlQ6epe2mEJYiRvyW5Ui33C
Kn+10Xoyex9mETJ0cDYwHuSBnkRtp4f5kzT6HqLOw2yAZgvNHnNwxhtxqFbD23Lp
i5NoA7w8z5Lg2/mCdo37+6eIId/DTQ4+lWUB33uO2E+wcO8FJNignMHTnO7J/eJk
JXZ3MdSt6ZDrIch5wnqV+herJ6IvwN/OUFifo8KZar9bPsaLnSOo1gnA9tIJwWq6
ord7Nob4/r7uA1LhDF89tcCxP5CUDterdo067nJGxm5uIcmIA01i3zgx9duZ2By8
keMm+gyCUdXexMo/Tcq0hkjBaDp3z7kt8KKdmenvTcXXi4uiPq5H0nno1iw3Gh+K
78tdabyS2eecG+8KWb3nJWwqhrjkof418sw0NHaq6yQEYxmDeUODXmc3W9wRWQUm
ZrafNRhDUqfbpGSQSS6Y9Q/QFdWLTknajkymiyFnJzlaMJQtCt3tOOvF4vhtOIY5
IWBXAEMsfS6l02TGLHlkr35t5yNGEZOAS5eEA/6SG7M34dUrpCKL8Mx/jNO4WpcW
PC1f51GtGb0xbZuY13k6E3Gon3aKvEJciocx3jE3W8rRUV0cgw91VS08GWbDvT6Z
h9nuEG6bDoLWxsWhrpXk0dM32m2eEJcBcvEJCR2TkItdAWEV8z0QZgtZGqBnZV6J
MJv4vSj15kqXfYaAHKaxmVV4msxuIxTxhMBGjHEMZQfmutpUQR+gnmyr1IUO+0I2
DiNQF2CvxrVYo8eXoEZf2q4QLKiTyNvED38n6GIw7uhTifitIfbbX2fUSgURTbwg
o6kmsxG+AOrmgerhoQk0RachhqcNm7ycSiS6b7kF7cadIWWxWxEUJULF8kXSSs/E
ZL1bl38Qxl8iI0RzzYRGszJWRufYZGCAhEq9HmHJfjhGqpjJF7Ri6aK7opdSPkQs
OEa8pmIcSxsUFEH62MK7KYUf2B23Qqod/o9ZvcpiLsZrXTxtVfExuKIfeLgNQz4M
zMHsVhNyxM3LdvKBhtSN6oUwG+EQqK6cHmg0A42MlR6q2RxQE97Hsr+xWIoT39+1
D/b/izKAVUQ2iA9ZzZpx8HgzTXdblGEw19AOs0SAytd8KZlxjkq3wAsCwPT8UXef
Def73vGieoWIDhwdVnwkc8K9UzFwywUHCOFKZu6NfkWKykNoYWZfGQIe9JnHHJxI
6NqGKzJX2LfV2jG9bRXsEpJQDRVIuOaFV8MhiyfmyrzsCogB3vtA0HQevhlbW0PI
2ll4DBYchpiLdelIAmGl4+SrRVsglHsJgEAPDT3krl20KlSu9UebJjXZGvzUy9wS
rOJ7Vy9fFIilird9q9ekFj1OZZQk0dhBY6CoEs20px9rmLd4AZhhfPrgDAiLdTyU
hKmcNf5Cjyo5QkTN9uerQu8pGK0pj3lkKZwJd5FqeQKadoBrZcdQrp/GU9LLSaTd
DJVnzioX6wqeiSdmkLc7Zpeek+x0rAxKxy8NY8dqVAmWwgR0N0OsUB7m0vHSmUhF
SELjzH1Ea7rYSSrij2TNI4V5e+PnQ+pYD9hgsH2V5mNwurwNWZhITlpptpgZ1fKs
FZ+aB4+O5p36VQP9ZAVz9lkbuQSs8amkvT+TqO1GMy72OqA2uLzluN2/UAn/EhT+
c5ADm5CEW5si+z0ralZ69iBfkCa5iPNH3ZHKschDPrwT2VEI+340k39IaCQXpbVF
WYfnZRM/k6WAt3aMJ+RZZXTkFd2rU3bwBwdZIMH8cDzbigo/IaOQvCF3rZM5H4Be
LKkVnBYwsRsC2Y6V+UcdX8pus0kj9LfNgmsIa6Ri1flAlMpLNFh1+WhAVkXWlghP
3xhXO+XARKTdkMEtAcBJDyghbaN9DF0z6cBlrLmGDvAcLLvux2WmzLKBjL4OC9uJ
GevyTNjYwjDDKLrzMJXIdajPGKT2POreKsALWgNKPbcPS+LNcupPRl/I8FToWvEe
YlH1Ir9Wr9j05AmPqIYMyM7rYHZb/qT46dOV91qYiFy2d2eeihFNkw7y9OobM9qd
a+upTqVwcpKq3rlkd8zJWltACjm5n7Ioz/9zHyhQw0/CZSnq2Go0JWm9IlAb5dWa
hn/pCBlcsO1wf6ZXFCCZdn2L/mP8GAqVkHfMwXI0YFfhtWpz6cZya8hCp1MRoFF5
CV5zuX3EwpIEPkLh3x89EcMB6VgFM2oW2iDjMfMio383yUnjc09Biuf4ucJIMeKI
VtqTHP+ySlALHodlOqp8Loeq346sauNl8UACqShlIXcLuB7B0XaAU1cPhwVnOL17
b2yQC1Fnogr4cnwX+REz+fZHIIh6187OgUkX31i/C4rLXUbqUaPFtXaJ84MgY35f
cSnc8eBHgnssh3U6D4HVtJTANUUIXjNZ7Q6t2VvrI+PW/e6s2s/Hp7XqwAmMW1vP
Byd9DfUGNKoxT+5d8o28j/zJy/jNNvDNX2uCRYAXdy5HMObdFf21yCQqNm0u1RLF
MIyEiDADaENAzEfdciP+lF2Mc87I2xRqNJGNlFEwIfFTQm+5kGxNS+lDDpgShWmP
PYwEuit24U3jVVJOktzNMdw3JgF+tpCl73UkTsAonH3zEta300V6UI4qd5r7yJBo
EaN+0ehrU7Hmu7kynoLSUmfyjA7x6vSbsF4waKsFd6uxy7SxNhGzn4S9h58rkin1
6rQEheaWYHlXu3wS4+/ZfzHN2rJPHTX8y1KOvU7YCEgykZOlTEazRKfeIyH3fyQE
nIduWuxI5ZfldYdF5LZr/VyxcLtXBTG9A3gsT88Rndmm91ZiGZDMYT9LWa7BmaC9
chnnLH3djQBmSS6FLdfq1O8vsXVh5QtcwxoZSUFRRUwie9HZHAr+KT1yHCoLO8XD
tY+IqIUx8QakXNI5xvJIUNOchBKx0jKw886PQAjFoNFYXu0DkHG3ZU5/UtrrPjrf
inl+ipy3898L16nQ+nm2ROyPiu1NPTfF7vH9/6hrjCg92+q1WzTg6iJWANvN2QFl
v5Y8A6ZeDwh4avQK1I7gWnhokBXz+xCbJeXjDj3FiYmt1Kw9hoStwzKZv39V1sPL
+HDOp13Z+okTbvQH0YHBEGVQ5sj02qLKNyVDcT4OIQ6E1OmRSrALqJ0arKQlgQfF
hKTSp6qJXg+x5K8CJjluVYi8vcgzJ6KTYXkHxrrlT4DKUcFhP2+L0DBg388QwNAG
ICw2vVUqouPbBxrHPo+kBjAh14UW33A++949bABBBPgBjszHDhuUbBsx/z37R9cu
ObxyQkAJ8VNz4A7CGLGHzHBFtA8WK+nWpWEvUB+fscOFWhq1zp1KV2nSGPmN2krN
0zWHtglXp0uP0gSaYyrrP6dzW5EvyL21PiSQZm9MPwKNvJ4OC3/Yij7e4m+iFg4u
fgXDQmzAzFJJfUqUdxqNRBYEB5jDkcDInkxdJ0+palAMjDBRkmmntYT4SMjbykJU
ocOYU8JcgYB5mztZJSfC8P4+psfDU3j7Hno7+xfnbqgjM33MN+iHTa24hNZcnNMa
myIiUCcbTT4vxfOouuUPph7f8i9U3AIPIbjrZg1tpaGb1/rHs6D9J7mk6V3ykxRf
nnXVfqGG5dV0I8IoYHfqDMT/EvnWhMaY+Xc5K7llVuozAXOLa4kMKLaf7kqLepx7
3VYfntaURwrZEQtqrfELi6XkE+yD8qrXe5+UeVkFxL548TI8TF+zQ/V83JDypsk5
pPdMA1UmSzDSDtkU0jsi+WAccu46QehjVxLwVgBEewdhoiOvA72m1IEqLFfM1ynV
rxFMFNh7fm5DGLoBwHl2ljC68AET6VUpyUyBn1mVA7DxEdQ5mttldiX/d1gImMSC
2kb+dVmXdWLKVOYbt8JHeDOAYuUBmJgU157SWil7oh3/iSxqjZlLNXdl9gAc8sSq
CMOt5KOE9XXoR4/BX89o0WQ/AuXnWb3YsGehsi3ldNRdSWxNAsx+4tfdezWNWjXF
zs2hCWn5ssnSzTxp+BuE44vdX6RGSXc8SpM5SOvPRPGLEW1qDG//b1jZdyhiMarq
THXwFBCrTkY9vckXTX2bvjWjLwIN6CtqGXeWoun8XMERegCkr6OzFzYr5PEAPAWc
vWgfNU0EUFWz52+d1+ycWX/dzOW9OiDcqT2I1iNUPO8kb4F6bVRhtH7z+/dJqJCS
NI+TnBaSyfCp50GtKaAGuK7z2daY6ejT5B6T14FhDBisw90fB06FiWjgddT6/JrU
6YXato8f6er9y1aQPJsCgv0CfegvXcjjD1DnbKiOYpLQd3NrII02UDkYHxhTYUw7
et4jEct5sFeneWh/HaVhumH+7BMxfEO+NQcfAyfxm0oL5u4i1fMkaQD7WoL4EcDQ
CT231A5K4L5Ej9Z3yZt8yr6WA6xHseLBDHwx+bBg388IEYBY8CuiofrHJ2j47MiK
uA/9UFbHyDXjgSvrTrfdXj8lovyGFilty3FfsOb8wY7KiegcjG+njZzAx09AL5vS
s1nCrtKY6c0xWh1cbEbiKSmW6wnOhHkVIm1+U6050SJBJhd8+IKW4d7n4RpjwCr5
Mfs9+tilibg6ofpeAwyXJPNHD6clm7tHzmqS2LCdWOu4mGwLMXHzpjUnHk21qIOM
XCJRhpKrBkjSKiyb77KrSEE3w2P0ZPyOb+1iY8TqdugSiO8TjJ6JciluXOVCPRNB
0Ox66kIFPHwq6DJVEFLIxeAUETCCHcszdhX1i9d2A9f0jTtii9WjXyVjp1GcfQTq
gpN9KO3DelUgA0Zd1chIlrlw2/De+3izjTSSpokv/mJTX52QMZQVLdWIM+Y3ZAfx
TxqMtzNkO8YjXtoGjSZLtRvCcEsnDGwaphSpgSbGQAdVOKYu977FPNV2ZMn/8IOV
XKEE7LbQGJuaNyvBQEPOD3KDvjWyiIezSeqxNdIZlJWSEFWAH051v6aS+kfJab6s
cdoxA0dkmDGHvKnW30v2jeU5ALfRjWERNMtMbvDgrlaGBnPDHMyhZ0A3w4lgC+0B
DQS+1JxxZfinBsHFBz9L1W0euNhKJ/OJRD7ifN9BOiXBV5jALtPqq7gt/TZuSaTX
r//fA2+alc2Ev8EsAiT6T/akvQzbW1xqcNXBuaQTH92XnsPYkcHvgDdFRH97Dtzl
NLMUlqbipEOVMsk/Ehkj8Z7nCIyQTh0QWCKgEaj+rQp9j9uxLc4U3aV3YOga9Z2T
9OHxdhdcOFuPfZ2dClPoB510a4H69qHKQ/inAThuSZDTiacI2X/gNI0Zm9MJd2xv
Muew/UzeMmLHMeUx9tLuy+Reuxp7HBLEUDYApSQ3ZAgMiPLvsRiW+bXNFyVO3xST
zEpCgzrGCGPcLEB208XdTHu2gtKJbaCOVJB0TVZtLOsh94KIHScNxaf4sMujNbCm
PLcbnNCp6mJffmAT8WUxZUiNpGW1Dvlyq0Lhu7aH02ibj7L2I/MTHZqnk0MdI2JA
45mqqHVV3Nf+E28z9Wz47MaEzuX6IkmoSfoJHMPIMOlZUOd7xpqIOTrxaM9VWhfQ
L+VGnvJKKrjMynjEb7ddDYpk4SnuYE4CAPdE1nHQjWS0Pf6tIMteYHGtfDYCfuqu
lzxOQAIzyRUVWyUC6YnpMjLMIQZu/SCErx5wsKIh4WkuZLWl7zQi44gmpUiKwzVH
JwaMZrNtbI4joP80KocOP9gAFtx7LquDKVQYJHMrsmGu10G6aGm8AUDPtDRNtK8K
7jU9kGGPu/gidTG0Uya2AtDs96KYp+WAIguF0Wnjo91zKmoXf53r26WkqQ0ory3u
J9r8kOIvwBYIEvWgEsajuk/f6ddfNldpsOc+Y7MIa0EL+VD6578uqOSMPnrpCop9
sXVvfC/xWn2sV04/FlfGrD77XOGkVYeWgF3o/ih8WAKVrhl05GhIB+OsHWcPH9Eo
2FGS0JMs64KO551CLn7hsQ4UOYb3KTjCzqEn8lTmiPz2D2vizvI4zU+p8iwawOaD
1B9omNL3Xog9EOQ+KMOg7MKEy19XJUIem1790bRpLvr3owOPZbnTe4/DalKRiF7v
aVfnsoy/DcmpXd2RZ5ne3IT52Ch+GyAXEV1USaO9NyojT/RQCu5zYOCFbO8zN5vv
29bR1UOFxM4QCbuYpNGWNuQqlst2ahxYumd+ImEdr6fiJEIjssU7ef29obtS6K+2
lIrAE/cT65TF/fNimsJNaY9gmXFtzDNZd27fNFx/YCCQ8BtNf6nv0zaqagB1ylc5
eEVrR36pz/WboTvtd6lSwrVURJcPTKGNyIOzOCeFnpBCE9WlZThOkq9+0jV/alJY
qrFIHcgUN76S1IPlTqAKb0mUC6A9bVYUAAOFXnckYkjfaUwJ+TyLTLPJUaFYFuD6
T3v2INcebW2n2lAtkcT1pA9KmurkMJKsBmqScNuMQ2P1Tu+xVMnULGIKRC7gAPX+
Q8Fz1V44y1CP9NNZ+l3vRiw6s7LQiwVuiSHe/9YoCzzjATD3B8/8r6nfU/HJtRBy
Gri0RMCdjQHHujYDz/obF27MxOfi70Hvd+/PLsBBAjhE3zCZkEw5si5kK52y9dp2
uqXgL8vkKyx3FiO3q3G9KScwWzMG3l/AdT+ivfbRSYP5cMu0l5xDoXED+aSWFlnH
K+mFWZbD2EtH9NMQC22Sn4ggQB4Wu8EVcUAOELNAZduwnQZlVs0up03sxJ3FYeSN
T0yip/ZemuMK0kp9GCXpwaH181kWovkHJe+nTIVh2gz0x50lIr2seAzxu7Gjd7ra
MsSHUen0iunp4T0GC0wuafsMSXeF+Bz1wdt4i13hcnra2mIT26Ll4EAUt7ICB0l8
WmAlBq8nxNYRM0Um4PDIJNFPNEEEUew4GS9+3IcanRNLTjiAbV+NSDVKB2haeMsI
9d47gJW7Mfg+l+sOTPMt3Hg+y+zOIWlL7DU0jeSfiElElXOMdWM1eostYiXl4VlC
bEtaDaHKQOE2AxElxhz1VqY7Y3TDGi/pY2WRvE8Ds6CoO6Ig5fPRZD7faOzhsDSF
0yb47GGLp117TXhs5CyaElQX395EjfLCS+8qbYENKWaI1/GlQ+MDI/adysl9vonn
BIN3SPCfQGFJeNzSrYryTypP/1Y6SaSXsCN2Zw26rglanek1abgyyZyJmmi/Ac57
5yEFEK/pWvxLWGheXarzd7+tvTfmTgToijcqaoJexF62Du7bzJlxDKJvyZM9Agrk
wg5kVW5sHEzf2GV8WRv6wllrFalBCnODdXIs+mKsdGAzO+67blN578G4UXIZkNTn
cx16qAeE7wJmt/GPTetf3edF060W3N/NC/QHfkp2t8xbCz8TBRcY0nVd84klX/6T
DWOMV6FgZE0jz3xw+TPAWDuGCnLAuzYy26wykpwdi3BnyJtQXJthcFkjK2qEaEXp
HleP7b/2j+590piSdYmeGRBYfMffPBb4vE8w2XfUbgWGaasOS19ykM3r0cu1m6tr
75nOMpb2RB3f0vayHEKb7rsyxXd9nftNPN9tGauDBhWSWMKs57t6s2viOAFQp/J+
IkpJwWeSCc1u6ijsnk9VJdIvQsBH31gyk/3R++Zd/AEqCYrLMAyCbzeaXRIbBrH5
1wFwO3wkV7o3ozvs4nAZwm4PJS0F3G4qiMhZqmApOaP/f4UQ/2UcFVe9kSUWgwev
8Y2tWWSxJCqBoI9Gq7RPEHkPy+6NSvec7Z1cA7ogWwT6yZYixUN0sPAzF+5IA/5c
jtIq8drXUEKBbIZDcJbV0BTpUd7gpr7/bXcm2pubeDuSbLRgYSKCMrXSRhnAXwwL
r1IlzoFsVSMgF4z5JuFVKK/7j67K6jT2ZdldPJtVvGKECm2Mj017SrHEhEI2X5Ny
ez5l50kH1uv2Vb36nyyiphsEDWyuEN4+G6OBU1RXXYN9sEQHUa0xtkub1UjS79to
IAeurEU38uQ0qQaJCHPJPmw1Dct72I3/5TEjyYIx22vbkI4uNtkVdK1DMIkzAkM3
Aohqik/iDf/VzJ604lwa5S1m/GJX6uj8xtXlH1Np6uFlCxuw3jc8THty/UWIfuo7
3i92mT3w/AtD9cr6sfD5M48ejCpbMf5k2YSY9oIqZ2jRJDYlndGq2Iuo5bIiesiU
/i66NaO86YTpXu55KN2na7/YxdjVqXmTEQbmiJiZUYEGs7N/tIcXNJiQHFNpzLQm
2c4J/047S/U1voq9MMY2XOYiMKSoSFHLe2f5AXgo32jIfUUi/nFgGSXL0RfjnHPz
BaWYyYB/8UTJtMsUnn4qg2EGthFrRhBLuFrgKT/1oIRvpVoxWEDOg12Zy+XYuZS8
u6N2cuJML45iK05zRvW5OWb6fx4ezNWK+LaAN0Y+1d/V8lOAwDZ2/4r/1R0gQpCd
ri9PXq6Xw8xZ7W9DpM1U8GKLcRGeK6IKD29ztSKe6yKpII7sT7NDqG6d7CTXEKot
ZZx1zDahQbnRMMdgwfMU4KyVfR62HQzSlYmbPhXLrGIJX97ba4hFox+dYbLdxTmB
0J67ipZsj4Mb3kpZ1qH6pNCSRZlN8GCNoATV05DvQkslk10H/HLT7NPcSX2unipG
vrD1qtjuPkc/HPMJty+tDVItGJwDZSmMTTYNXX+PcmjvdNDaUwkFjBXb92OKFYtR
NjOpdgThvz4MA+GLdnwCMu5DMwBS62ziPM1sCPjtzFM8datKLbqs9+LlSJzrNdpY
WRFg3Qsmnk9TW0GxBdI0Wo8ptKlI1NFieNfHQReuFknhKt8gj8Mg/ucXCr7X/WWr
9pUSxeYWQbjvyYFgildtsbNRomvhYlDmz2FHKBN1XDbgbPdcKmBypYaeH/XNP2TR
ZvK2NpS00c2yh8KtGSe+1NXcP23CIRAriGJLFJCzA8ktHHzHYxQ2TWv1B4RUreD5
s9J8GBEP/HQDb364mVaJU+4EZ0z10Kw3IEACtzqJWCTYpZvjfoih9z2cMoMVlk+L
DAhxuh0YQcARxzsbsxXwI0ORq16ANGw1AGHYU1V04oqJaHi7W02lPPJtS4su77as
TXhsRKXmAkt+9NqEOoIe+3etjCKaTnXqEIGLchQci0Vl7OzVnwPA1lRa9eF91XFo
FvhZwTVv9xhH0y7xfyFXfheVsfKhi2oaaATc8vEzkAD7C+eJMEy6QhZ7jQaLrdsY
hYjnqL9lWmqXu3KQKQ3XpBzGhCtraoVA4kXt44xeyWcYEOz4H6CoxRGYgWIGp7AH
beKBLp3PutLBtqzoUQpL3PkQYq9iUCkzQErbaDcu7cBAAhnKGcTVZBIrkr+JnBwm
LwnwdGI8VtgrpRUmGZq8L+KR3TV4eD9aeJO71wM/ZQR0NvSlQnOmTCQ5qrTSffSF
DBWGbcKqcJ6s08ciGSz+K/p2uw+/Dk8HR4oY6BDyiAmZGBk2flOUWMPuA6APo3Eq
O7knCRneiL8M7G8ABRha4tQhxvgKJZd//IrKAgXKQ1kH3v1PSCU49xKW8kXlIJkh
CDgHrfeerePp1M3DlJ+gTtOzxqUldLNU9zp1QgoirpJoOY405VaYUeCJFkY8Ew2K
PBrn2cjnQzOqqjnbp6Kj6POeixtxT6465scJPjlLPSdY+wLn+Hp9tr+6Gtb/AZhX
24yBBbKcnfpZadiLhQQy/hXjcACQMjTinaHJzPVHMemPSJCbpXR0ma+dgPn1q7T4
w0AfdwgPuYBpQ4V1eTAsgvCTW7kDPMlk+lzO/LobecbTC0sWpbrL7VAZQ1BHa7Ry
P9xyYsqa7lePCtweKtFPWNLonL5n2GOxWBhQ3ScXcz5OdEqrJE0Bl3+O+HvSmQfQ
Moe8k0/1NGpbmi00T0gP8ASXt39dSD9L4IBYGYBnHzXKaxxjJL4TwTzL7HU0FWfF
NnbQIB/KeX4eu1w6NJ/TVyHo5b1BPw1F5qvs8fedzzuna7R3Aj5Lt5AAT/V6jI4n
0Zi5MsBy2dNWxeRq4M/aDd7BpqTGdUwSu4/betXV9z4qIsMlnJZlVa4RuowhxHJA
hUqC8uNv53p+uEIBuNIHyPDuVJdx9N9L6pqTa4rNlaIeWoIJv1qGT26obZHJXc0S
mLGvH/ZRmskNVES5Uw8vnY5WWxflu33rR8r0LrRmhbgSQoN8u1Z1rwYbBnQdJIz/
sJ5qej/saqLOUXqPd97H5o3C0eEGfaSn5x+TzgvsdsGb2M+VLpTw1V8mWv/RRwGa
7z4CTrwGMN/rrpHqB9RAjg8TbW/qNUqyURsXN6YVsMRdWDzXd6aB5WRMR2dgtUZJ
Yptb+J2oeGZ7WrOZOiETXPAD+FuxkQlW6vx5pWyIPosfCA9bNcInjwjFUYJUjwTh
nTJXLmV8rvyyxKkivf7j4qUwztWZBdSC03VM7BdFxZbuxL7+mFwPjB4RuhMwKFAz
fXpAWV2HIdvat239u6t7aQuFm7rqpzrCsQXHVsh9kZoMCoLTq0KD8rX3+gfO2U38
H11aiaBzFtFilIZbI+NVhLP/T/3xK8/1sQBBAgExq5satet6YCDPzSJFujCWZuuy
LlSbkMUq5zgtQESN1b40aiiKMTE3gPX25K5CQEbklElG7d4wgBu+4igGDI5o39NA
rdVg+NuN8sDxg6K+TQQZSVhjUCd97BnDJNBN5KMHQLk4DQjWX4LiVLFn9XGnOxk1
LBxXGRWjdThVmg0nZo4bRHMz6cH3E4EhNmPSKVB3a8BHEyBPJDJ93/y2sGcNOFP+
6e9/Bqd5wLf1a/Vy+XmWvrg2MH4ms6tFbJVwGeTsckA0NGb7pvZ+u2GJpFxZ0YUJ
gfFYqEhDdC9yq8/Y9KbFV+juUSMq2zgfKF454rhKXoRPyVCLuIUsd8bKsKUKbZf9
ZNrkjN20Obm78N5OQ8FoWrp8K3bHcy135O9FxwkVRLfNRlT1zfZdNj+112PyNztp
8Y3VZehwJDEUPefMB5USNLPOjyGgUdBD2Zgbx8Y6pIjEvX+NgtXYRIfu2Y4LN3Mx
BLMS7ancu6yRFXt1II3p0qdICYSKSsPCrxtVfSH4IkltCMJ4WbTqy/+iAFP/QE2n
DvkNvSNpyFMpN2fwK81ZsBWmG5YpodD2/Um0lSWRiYRZZVpqjrtH7Erfoh5TzDUS
7raYLkhAxU1q9NuDimELyixo0a+9ac8umGmmiiGLRxwor89a7dhTOQ3u9Awp9AK3
g+GonUPSIJBH39UdAA0HfcB5X4TzinCPavCJQ+ays9dVARgx5Gs6gsa6/cHxUjEt
GTccpGUZFQ8NANKD4po6X/exlwFfE7yMpLQfxy9XjIpKvD4nKpqFnSB/SYU498bn
qYhDb2a50jg+Ol1QC9vI2gLB4IEuFvg2EdA7PGX6T8+CG9Hpo2+wyXNVRKwQh4N8
HqFh5LxHlsITUuLuE4lEfJGxHNRO7hhHT9PxBGulKLYtUJUWbrk2tV2WcMJ4SNo4
8GSe0NhAOTnJlALW/WaaUjuC5CNdd4dz/41XUUlj0rCLOUbvKmqQ3t15a41hSFSV
2l+/8JbdYjPq2Rg72NYDvQAxJGoiw/yGPRQC78QS00t5E4IVEX5LgOuGvFrqreOx
WBGDrVqsSa787s1MrSpJtrj9ZjNV98nj2/59UWPCZxguG4RFC4KXPCijJtoaxi9p
rN0mARToHEGxfyHdDlIT+ElmQkcxAc6UbjuA5XSAbKB6TLuianOQYzAAbCZMcKHq
2TqVeU+UnL8/NsBN6ZEmBM70AtEHQVeESJTgLcV0G+khSq9jH+I5e98BHw5fzhWt
6YFprmI0oYaRjfvq7V6ePtIhdpRnkQlNf7DgFPX2Nwno83rDYY7VHyiUKqeQt7zf
xXLR2Z+iiyECtn7YhEI4/RLVsWrPLNtIWVusgJ977DBWvgTGZWBWn2PVv6NAkbdd
xvpnK5qTUR+11S10FMcIx29yAOKrw80zgj+oFKaFpbURds7Zdn5NUeQp1Vt35I7L
io5PJmSnd7HMme5O9uQxqsfXHDhH9rj/M/wRhv/rrfdOUnVXGGKI8MUzEnf5gZt3
WCd1VM7FKTEyK3r+v2/6dF/0OJnIIL/1q3OoYaK64VPOgdzdsmma0FFz+JjbAwtF
+TVfRJB91QcHIscksxO8HFMha++OY0fvh9y7HIJhhKQ46/fR2LnDaMY0Bnewg7rd
9OxOSuYg0zjMPWnRd/YLc1RRE1DaeQay3hSxUJmr9iAKwa3zO+dBlFHzTrOuNiR6
h4umDF5lSw7mOyZN2rKYXFF7cfe+KUN+q38oK092HKRov1TNR3NCSMH5mmySjL/Z
rp2dQL33EdEdratvv8nrYLCNYn/eBnzFyj5cLczcj/Hvu6KjSs21caG/1PE9VIdG
2nyW9IEXle2SIPgnj2exgyDVM0ObbPc7IxBTKd3/X34O4E8IHcMEBWbe+0o+m0dM
BqQG/QllEGyCrgvDBTlGVJgOpMqmON6Xm13OcnOBz/eNdAUxlwuIkk3FC6botAXC
j69B4hs6OrbJG9ds3qYPOLO9xcNT4zgazB+PurnL8424t/Ba98SNtBTzpo//0c5K
AvgO9eb/yClkRZLYDj25z34fch8kBfvrQD8d0qfB5R2cYfR6gEl1kEinUqTgdA4t
hvZZrBBRDHPBDEyIekdvO2dkp1ZsRJiqEwEhMyVd+GsqpBIAn1qKEDdIlvO91X32
5JO3IApuWcpd8m4ekEUUzmS6uXqazKlj4gvpwotINOVDx+eQk1WlSXt+0WDdl8d3
UVBhrjI4lP/w3ZneJv5PIkP97uI/TmKssei6Tmi9ecqnGyYDI9qssK+wIWz1R89T
W7SmaRxuv28Yx3gkqfTgVRIVUXVZNx8g+HJYR3XbuYIbhqjcIwLHdREDgmBTacD9
UoY1geabKS/fJu/6Y9Dyyoa9IawqPMMJNm8PTMkv2hXpF4MoZugngq615la+enJf
yKZKaasseThLFrBSqG2AsbhgNHfi6DkNQ1oKmE+/G5+HaLu2JcyFKRjZMOQwnFAa
YmUUo/MaJaMqO8lac3/zhlL6NfoQvGJg77SSt8m8TR519xpESpiiLuCevPOiMsnz
8xLWilJ2ogNxqGeTFwV5GGVZH9SCnfGDuDqeC+6CtxdbQOG0BNO0a1RkIUpG5pen
CCWwvas3pc2zJSS6uZuQvHdk6Tb3DlTW3Z2Ef/5KTW3U1wKGtNexBx1yOrrcA5h/
0Vxz9i6w+jEsrZmehVFkghRVIgb1/Fa+ZJ54/QfJu8+1WkjzbZFSV6UkuCQwueZK
+Ky05eZUr1/WJheglmPT2kvwiz4yhJk3Zk+sI/+ShNyKNCyl1Dvk/ySGguuSfHyC
WAqD8Y/oVFAidp/E2dQzJMO2ZiI1THIAX3pL+YLya3lZNakmcn8tuLifHsxV1Tl8
WYsfnHJ3JHl8uve/JXezhx391Ecp3HDq7AuszaR7yl3pGjEQHJf261AS2aguRPsZ
6nghdgFbpjZAD+2fPnNZ5BSD6Zp2E1fm89AUoQb+9s2aojja3XN/YD5BYn9aV3vG
8+lyraxqLC6d5dyOjSQfclMSfMLJFqcoyaZEz59RsuTgac/qshgXIRy4z7WFT5U5
7IJRAg3Rb/9UbLbQkrM/y3jjezqNaJMfxi6T3RDGGGBs9WrUcP/UaxvR55KG6ilt
27fB1/7jhMqXCjimU90yDsEinCPZZ6vn36kDrHODOnvp4Du1gAS44OAGYKLC1MUa
FB6BA7st251rn6nf7PD3SLo/g9ENI9JvsA8Ln+BMx8lSUuX6GgCYPpQRVCSFplOu
QBerBUyUfGsABN7ZVR6Shgw3llcA9ng/qifis+WuAeE77ChFOv7rH01yvcLxkJ3u
2OuSG/WomNpK73dDfx1BC44G/Ja4lMvQMRczwONG4Sr5+xZ3wBNkA7UVSPmeMTRr
XN4pU2BgdxPXFPjREyD0fYHbsRrCUWuj9xGGIjaegfS+J+h1ZMDCWg69xaFShvue
zte2P/06gCrjF6fyppbzDauYl5fcJHQDjmC1Aif00Cby08s9rh83hvDWZQMuyUdi
tq/NM6jW5fu2jm8YR8l8eZe1fBM4LgjYQUrotNEo0ltWBSHEFeMXEXhwkBIj0LZ+
OHBpJdkYJ35cP7PAZuhNlARIzuTzmuR2h6ZAEZjAG+7EmWhKjM2H0J03Y7T7Phq/
bqJKGHkLjC4DlvtliqUuEQ/0lI0vagFowurCw4+vS6KYAGtUuQDybfR/jZuLeI6U
PspNbU5ElOnGAC4AP/Zc8YwuXp1n8bqBFg2g+U/1vQ8ABBDB80bNzrW4XldaVelg
h/Qxx9d6aHm3zQFsS4Iya45dfBcUQI4vRSD0iJnyEZbrZQR8nGif8Ljpe0fA4dko
TBBq/RVBLbmkOd+6dOh38rXk7didWZWoLTd7uGk74sirVu9lRbGBXfJkGFDRb8xn
JirnqhbhNico4eWO1c6DuP5gRT9Ag1m2ujg5hFZTG31OYnlTQ2AnIlYzlUrEcKf8
Els86U8oAqEiqzF4/osBpPCA0yUe+IgG8tB92FGj1ZgbaFx57t7fuwEut5ONRXa7
vvekDvP0jDNO3a9dVEUqWNNPBDB6dRoIT3RiwW+ZEhVh2bzybkUQdtglYFeEnCiC
+syf/bZYYiyPnKvV9hnUnk6xNwmndCuXqHs3VaU3mZOtQRraPmuYlunzKSppZQ4O
kRlxSeJhq9UivtHsiRcaPYFCuPF1C2POmN4xqgI+2yXPrliUTSveON7DaosNbR1q
dgk2695SysdLbRu6vubLmwtHk/mGDGdII02uZCvdXhYciaSxZDRaxnCAdFwM8FX2
iHatX6ZFLkBV8ZTOwjFL82bz+2YGyw0OlS5F2u/05sk7Y8QrxNEK+/OL00D7K2nw
SQDKIKHm/4jkxz+d4zAQTdz7KlaGtrSggOoEM01Y9/RTSj9trsyboL2QTu8qOcaT
6foNcsoZ6Sz3orRhZM0Ypg3PDc5TUsKRU/ejIUAzc4OBh/MBBelh2T7hG9C2I19e
D4esxMsf9l0+eFp9hXQfXnV71XMH4kZcKyN1GWj4IAu6J73iqGMkkMKKz23vGb8u
HEusG7YdCCAAF+bP4Ykr2hZfTvNBHDJCtsRCQFBRlfZwsGr1qcijqPp9LSc6i4E7
W2dqKwn1zOcJ76sfq4itp8aZJKgpvMCrT7mmB4LRsYWpWhsyJTPjIkOAZC0VmO2S
CTfde6nnZzq67IdOn4iagPdlUL6M7PglQxg/7WRZPEauDUKVfazzPdPdrdhYOOeh
eKhFbjr/W/eZxwy46emAgygehp0FoFLVSP5o52eeqVe1NMxoisHW+jglutstYcEA
v6oq2fya/PXpTxy1S7VUxtOV3se/4uO6EcsZCeMwDTORFoWaT81h1mAwtdzNdrZ0
AU0W/ZfDw8YbBGb0R/82+Sq/XT1QDf7GXYJX11SkwcBg6PhtrdaX+y9jNPFblwnX
WQRXHopl5AhLcKs3NAmIY1ci8da8xlrJrkP3z9hddkeTlFXuxZS2i7bWKyqJK17r
zAZEnbOVTVog9AyHMa3mdl+BqqzVR9cjdKYJWZamNOm4rc65Yc/YyYeHlhIdZ2Mx
/XQMHPStNObr1+mmiNBxHj9xOB7b9cBq1BnGuFZI7r4B8MmzHlPRaWKPvPY3irfK
FJe5u1iVMeJw8GyhsGnh+O/SYRMuNb9neqtyQJDAij83BcsQaOcHC9rnnOk3F7s3
b2KoFPsN2DrZC2LxwJ9Vw2jgALJoBq5Svu0gafP4+pCpcouTL7MYbgANUpuaRjUU
D2je0g4IetdcK7TfPjhyE0as5/6DksYD7Z68XCJY1PFUq0Gnxr8mDeIhT8iYMlt4
kqAtc0NkGRcrcG4voyGqhZztJPxzjVdituPysrUfpjKMVShQ1+562w1UpClhS7dK
hfbK7pWfK6SPiJOGjOXAvSvfDxKqKA7DakGA/XLzad3uYdx4X6fWRM15uLxgaPmj
Z92MEmCxvh9o3dMjkYVdIV84vk8TRzaPHjjDfXq6DmhG0xdXyqpngPQE+XQUm9WN
fEzYsEN5z4P7iD1wK29cRv2fSD5DSzZQWN8UVrxDs7ckHTlcZ0/LK7eW3WaIYtnn
cPD+zHFT/DtWpVFNGIbmb1JfWpP5nWsGyArgDwClLrXanj+NScmr0ifVe2IZAWrv
2ntfL6gmtGUklgBMZ+ihVyC3kOdLNz5NyhhNPaXPwy9MdZSBbJd1gVKzNH4ov1+w
KvhuFstkky0xtllqK4g1m49NjYpdnPJMklRvNMOlqBx1voSF+1RkWBwUz8ngGgm4
eIbmLb/StlmHa6K/9H/oqeSNrrCWAYORsR9WME0QLpZxwFL1TVgQB6ALfvBo7Cty
8Qg2UVnVNosifxNVJx5+0fx5vTjwDYs2ATHJTCg1licr27yIboMXQ+JdbQPVUhcZ
DjGGqZuy9lp12cXu67PRdPJjpNVgUWE9HWu3CyJ+tSSRJi6DIKxXI7VMOfEEf6jS
T81inGC10p4wqCQIx1U9ImEYEiAxtUiZu7Kg8Luv7qKSXFlylNnLXFgyiTVY6kq8
Y1osk7Kydp8OnPf+9566s6/F33k2JXiE1sTWQElK+s2gY6bA2yiV2C546hIa2qzp
Qvw//aJFPB80uPKCjFzfCn58tWW8yEyQcm1FHUhz9VEpuvr/jjcZOzv/TPHQmpFk
kcFwox3nJ90B2h0XQfgcbfjrYlT3MV+bHtPKRiEY748KICyhJiVbcplawTS3DAwO
Yu2u6PyhO7wWyERz4QM53fw65tDbeJnfXH7G22FiSF0R0km2wgz0oPqGU7prK75u
YxJvdrGnaiNyxe+3LQ9LEp8MvblCr/kgG50wZejLTh/rNjBsPTZS4rAUwUc11E9d
uySQq3ycPgrDfMATE6rsaCQRHqiuKyxaBYa07RzFuAUV438xYxDox/lhwNbrEFRu
Bu1Hq8+vMGKYaCmSj6Nox0SGVM0G7Q2ylPkqz5cHc6KqaYfBQvmtZCKuIuKyveHz
nxjGQbDHkUl6MraF9AqHFSiKf9lc5wGD7s63IpH/d0fdIeC6Ob0Y1NA+GJ30yzuG
ARG+IX/OG6g/FyCogJfFTkt2jBOQTlY7PeZQsNGk44fqPLF4dIZf3Fdnw1T6hPtK
MdUvWBNjcmAio1zagnKVULr9JUlEK2f5mnOSl8y2yMFih7A5VZOQMLeOkELobOxN
TSu3u64zowBysbREteTnJvPRZKQXFUucHzQgrAnYVc12LOSgC92SmUtuf2ArJ2GD
QfuvEyn1kT9BiZYEbX9m+rW9ybhHdTRjLCfyn9nXIiTo6QR4fXs/L2020Gvn7aoe
wazCRIKlb+YdxJUxeijBC6gZy4s+bYy0HGKI7wMtc3Sce5JRW7iL9zvnStiDtC2Q
J6l8TPdcQnnWGc6UNKq3huYWfbatR8/JK4uS/lg+q+rRusKzLG9s2MqDPV8d0K6o
7KZlofcCcE7lNH3hWoXaczyNgtIocILp+D6ydD3+sQIEQxzpccgXrVHxJ4UeQzzr
ljRGo4MH/jYsGN/pHI3N+uH7bTq67XmF9Lb3bKlicbRSVEGLKuMZXAgGkFsvUDsq
QnB7gOJi//SACqMsZnCBx9K+eam27vOHvdxvnd8YR97vJTL7UEPewY58grk5a0+U
FENvujrXKoCgHFXe5FOhIFV+AXUTxo8d6O0D5UoPpI9f+bcK3N1hLZ6XyAX7asCU
P7HqTYAv1CgQFcQOVQj/3eIqv+CSLORG5GxwGI7I25JzpvZW5bhbvv+8VsjLU4J2
J7RQIdwvEHlt/EdU29s1Cmw+/YWSojRyiWZd2jBjlnlfzjuyghy+vOVz//LjEWyB
nq9S4Btt6npQtVeIPSBRkXxFTH0wEcV9gDlc1PkvRaKe/KMzKEgW7FrIoByt0I8Q
tOEAqnNrRGwK81jU9wJIe7Z66A+w7vpaEspSbbmE2mqde4qjadd5vsB1/g7dQtfl
2EodKNvScZLNJ9RxKCbCXu6QM8sVbp5VGU45u9mKcthy0IHftfhxnCQdG1aw+uGQ
22Z+t+gEyqaM+syatdq6sK1XJF9ovkWueZbaIZykagUyPRFxlRQ9smP/L32J2YZT
d5mh71biHJWMPHSjOhfeL+UxM77RHQU7MQcU2IZDGoxaC/Z6EnsQuGpas9p0EZda
9K5xKgQYKL3bgYIF5JRGEBZ5AOxwA5UyIKbuzkK6YqwrIiPyKJgDx7tg4OeLrUlT
JlyN3qrxqpJq4OpbHjt0MrIrI/QLGIxcuVuQnSGU+/A2w+y4r0iawTiwpVnorPGy
3dOHCnFdlNyN9sfFunL5kEQmtXtVCRWuuqUW9WZMmGngFhUsjorGWnmCd+x18MlG
JUc5T4GNZ60nvKvXA6uW7sK9xb/aszo/iAKZ4MWsRtkZsqTKO8U11EMaUd5ta6Gb
4GSxxzYLVJlArj5ptmGw2o5U3FBatgIMKUzMqfjTUkJlVW9AqaDM6EbeD4a+Qf5y
K4AR5i5Zr8JNSMuZKAlW8Jj5IYuEUucqznoAyHkOeg/jfFLm/J5PsLSY+2D9dbY2
XPmlOVORcTxO2w1Z59SzKxIPMR7EQ45lzI5lwZhOdF+kL3QiHbZDlCoFztFx4T72
NBF32nJb7zLcX+UInbRkM5JglsvavjGBTHOVql653EC1ZxTlDvnwvssE/1Sg8ZRf
79XtIYnYqQ5nNpJ5b6dubNW1YtjMdhvyeh3OTSip5AJ9pbshz4S1wntNWCP1i0vb
EZDvpOkX9ZVn/gjlJSOGYDICmpQY3vWsFQ3Q2x+dcQj9/qhtEA1gY+wNJHrtTZ1Q
eD8+X0bpSk1uohPrQDaVJcK8SOuB0KpRvYg1dj11PWbCWsscuxyXggmHS5n3wNQk
v2PkOY6NCHKIRTtMcUQDt2y9LLkQGsTBEAo/N+R8J6znFFKddCmJ7p2c5K3aKIZV
s4JV+LCZqrwTol32J4ldeEtquW72PVER4PwEh31k0SOXM0Ar7tOQESHqeYSOmSN9
6z+7TtMvPs5u6v7aPY/5R7xJc+gkOq1IoOa4dVBBFGkJkpPb4u00NAI/ddgPiJjH
T7haYSFUeM+M7EHzv71YEWz4o8xLo72oNWhulkHHDWHoafoW5oOZJln5Kyyb0WN7
EBcq9LHgsyzgXJD/+6x+VPuNVFm/xYTKWHwPngl/EgPpza7kaLy9ko3hPH+BOGHW
aeMOJIR5WUHEc/WJlHNzpexsMrf0GvvW5QcZqW89Qwhaqyje1/OmH4yrshut16HR
1Yfq7Z2eZ+Ou4QAsVJLczuVLQqyuH3HgRjWNzbhQTjT4jmqRvP0DwVFwiU/P0Av5
rfqVklr1eKDKHYD5/GIKJXCuqYs3c1TNAMcLR3cDiECWj4SHfHKPQOTQKkGNq4tA
V8SK24GeW33RgXlb2qaBBK9+pzYLgdCiHrTWorjdX13NnU8MOQFA1Hm6qii6/kKF
3n6n6632YbybOmYfcNrLauRM5sU7KHNr4Ce4HOTvuWiNt+OKJyOZ0NPvangP0T0c
K/8t1SDxFMF0wQgs1cUp3cnvnztVFmMwJ6TRqFXLcn4l2aCE7FpEaiTeJ0VaZb6M
DMDAiVPGSgIIeCzpJwbXPBBagkLMMpT0X9gPM0XZxw9kXaYiFAHZqffUvoN6CqZc
7rj+J+4sBiuyyojxQZTt+EvU1R6K7lWIrZKQ5NFcRFD99Tj5QV9kekLkhqiZcEi3
w5g7CyYAVAxRLPJu0ftqRSYaPkHxhpJvMiOKzjiBuamg4LI+orNmK/HcKgvcgE/1
3Nue6lxPvBjXTqflQp2cNVPog9R5byInF6WgCabwz0Ki4D69VL6kjFBfLRShyB6B
wHClDDSzG0wzQ3LYuzxR7LZQv/Jpv1UXPHNUaKab9weWxFp/c2Vmx8MavHvEN4al
k8+dZ64fcyy3XHFTdUg5aANtMiT4MXs9Fa0ujZUP148SvfpTOBAO0rJFUlqimXN/
ty5feDafQHMCwOs1az+p46x18Z0FsK8EA6tADgQ6s+0hNpqjA8uXV7qF+dyx47ot
PKd2oVtsMo6XX+ZdokNBi+VREHraMNzAifTQVEEjfqh3ubQGXr0xt3vUia+WrnMg
YL8v06nmRIMikm6zbgeD3pd8Og/8p8NlvgZSYVtp5rLNN5farJucfVOHrjXdIuq5
C4vRRAKx5t7y7dqWUB1XVCCkPOk+C3ebNf89emnYAn5xj7QI9fqZsJlfTHzIJ6eG
BrVipAQYI31oYv4Dcq9eZjPl49Q7AaQE1KdUTU5gTYbFJU1uGSyuEei9Idom2Qlv
GxThGL0jcPyvihAPx5gyzLsXi05PxiYDz5dMkVg0+xono2DlfKOJiv4iLskaH76Z
qHSWJWNpxV+lNiLddgw/cUdUJPl23lMvbvt8dpHovVA+PwTdlzkGAXD8PGieeJ+d
+4/XKjm0UTNwDB6aXS23nw2+4nqgT2Czoc2Bc/tNMZJzoW0cLp2ncs9UeQI1NxrA
APTVRHwzvbP/YjAb5V8Joh7oUMvNCKdIMx3/GNVGhCxe/OLl5W3coQgt8u7EHtmy
6N4jSyMLtqatkGtY5k95HJMkNlxwVmOEHpXIznaB+1i0n/soBf+vDCuSkjvae24F
eVKBIZQF1Yloui2i2Hz6+NFetqyz7Byi7jtq74wM7ZQBTNAyN/LNqX+UzeRsK0IH
lK28uxpVyYH20UbI6OrXWastachCfZJgra7+n3PUn5S+4kqNWw5nwT4+JlB08Gt5
c4C7GSikF6CEsWVn63WDLk9RB71sl7EdJOqOOzg6ZYoHBLvLcy+qyybiw4BeP7Nw
DNvxH6RUAEw8phjEJdqL+iLsOdrCn/5GyWK8oRzLeMOArDkAPz0QbvMGqScBnN+y
1G7xdwFD2PSHApNvswjpHFMdKF1rGCa4Q4jHhe0qcQ6G7uuH4kt/WkZNDBvIfO6F
pyHwFzf6GJn+KFwGPI84RD5wJvDa7URtpZlVxrI8qs22CPGSyvIlQEtKzmkZfqDL
l7/UNb0DjqKBYZ2XO4H4RNj8p8Bi92nZJ7C1YxK5KwaSJZFbFeP5WrJ3CMiZ7ESA
RHCxZbXFskmqcrAfQOshOkp69/yWPFDOa1ogBFbGwRIcm11LTlcoTeQTTZm5JyDy
jFZUU+8ESvT69d93jdUl992U9ujnN2KOYId3JkxLE+ZBiBojpK9UEPM3oRPd72yI
xfnd1YAczCuPj+gIb53jkrj8HBvTjNOixQ7BWU9Cxn8bM+HirRJEXp7Uk8IIOujS
u8GtsWmIZpgU3TMrttIXtjDDesn9hilu1euFkpddy+an/JJQlXCSf7giWDAXIyAo
WwA2kZM6o0GdWP95s7isyFoizKjO3RJsldnXg/KwrMrG9IeTUiKUY+V3s12jDL44
kl70+VaRoaHH4gCU4aue+w3+a5CWBom/S0NppHS7mlcC4NYvT1eN6JhBI8/nf9Ra
290Mxe8OTqaCCdh/05Vv74s5+yIKBtNbCmPwyHffmM3DLd7vuPQjQhycBw1VMlaB
YFEtNcVtYccRuGhndCmNwxgdy9I0Czd1VfQORyjTEOWVOfAB8Pb/Tgc+l67sEEbZ
8XV9HhOMBQr9cHn0Nb5urknzgxyVcG3vcIFye7VUoApuz0aB4CRM0terw48/0q27
XizA3OMkVDYnn2kKWObH6ibGaT9crZd0CJWf1qht2CAUBavXnZ6fTZWm/SjY8OkA
T/2FahOEyM2ZtoGgdDoHOxAHCYWa38IlC+dLRs1bY0d9wuFgfKuGa7yvg2HmOYBC
bxGLv4YnxMzgiCzNkbTguYRUPpyY/pNRk2pP4/XKwPwCRVHfoXPRFbfYF0l/xrh7
JtGoXMADg0iHlOeAXm639VygbndXDsjBopXFJq4swCEkIhbfbaFE2y8gz6+cSFuZ
SH6DS9CasENA1SGfQEfqxrf4cNp8tEei81KeuVip5kdlEZVb2wvQyF8/BxUkK9p9
BQYAfrmRLUanbyb7CqfqPlcF59NKJ12k6u+/tI5rq+0mR7myhAbXrkPUAgDlShG7
HeaJrpUIQDmgZ2XMq3OfGxMWQaG74muAHYYlmqs/kO6nIDoVgULpXrFI1rhlZ9JP
UeigKkzd4yIa/RwEUDY9eNAYQFgiOIHn1B1oLmgnfjeVXMA9z8DpDj/NrML1+Sbg
ACH2BHcOSkEHDcQCkHw/qq8yp56+VQfxCSo1hy2yLY8lHqtl3Ib0KXiGaj/5JYkM
cllTr+1Hasc+dY2ifWWd90NIihsfm95rkoB0ZOmmUtmi8SwqqnJIEPIG++Qse4u7
zlaZXcjM6BaMlh3puutdXs1e6dSElDdKf13+kvZtQE0p+obErOjcI1k0qOzN8rXv
ukoxn4acMrb8COCjmsxhk53tDK8KQU67ChRnEHcNumquceb+OqUOjbwOVmocYctv
1Y1/xZfC1lFXREcnThcN/r8uZbBvJVTiLumg+rJ6Qq3eB88fHL9u7IgVpMhsusjn
+elMtP/VHj7hRAXom5ZORLZQib5MCtjyLETrKrCSfhKudRNOA3pFaUqCvWFy+30Z
+7/x9T9SCvYFJ9w7x0VL4Ih0BSeaGAi2r3ncQMVQ69oAYXkXqaPMzs0oS+N1kI2c
gabjr9EUX47sBwz+rGO9cLoX4GHp+0VbHzujrjUbF32U2ZrkuOvrhz55jqkYSS6N
S33yZ421Dx2NX2AHhIVfInzgfzRWL32NZKES6lTA8B6d1HyVjaWuQnIMd9K2A9wX
s7+xq+7EltXpAYtLyrbMmqruA4PVDWQh94gTaHPnXIMUfSPIo9f4k7SqhpoAVCiX
x/k2UwQT9I03ElMQUjb+8HEj+NyxiLfUH+kjYRuGooVR9W5DDnJ0f0vjWg6gMsvv
r1nAyvWYHBGtQn/gkpaFDpGAwKn6lcriM8fs3iIYUldOMhm4zbnQAVBP9IBfm5D8
AM+wo6fKe1CPIRmWnWxqN4N6jFlvdzgFddQKahPfxwfb9mLuVJtp42VSoRVXh4qm
K5oBu3bdTNQbRMnxrSfqMty/4kycY7WhdK799QjZyBWDGtfAs4wcQSfGVmN9kave
asqVLOBKazrrUF7433TUILPtLRKFLXUq4B9p5igmp9TYoHb28Gi5jYND4iJtKi/3
SszwOnUidbEedj15LVMR7B0R/gKUkJAVwZbMhxVXpOOgNVDJ5mU+6XWsJL5e3yWm
B8s/7FdfEzGj7StyG2IiSaVgrw1UBRexc/XCf3iTj+NBr7GTOBRKM3ETeCuOtkRE
DKyZ3x8l1zqu86Ak2P1zbpTB7FNY98MWloxB8yvkQKVEqs8eBKMbx9rcIerClpsS
moCGV5Yzks65j94EEW4pJS9MNX7ZKvebyMmekutOV/heFgoE1TYKIza32sZ3hiYc
unM4M5quksiFgyiEC2EOxmofPOvjUCHeV+JbBbe0NjJTv/8JHqNrnGY/sdaIfoGS
klZk3SQzi3aAK/NnKehMCh/VSbZT1FQ3ixiBPLfmNKih8VBNpvIYbG8Y1zCrBcsx
cH2sgW84mAzAAoDb82fUGb1PKBRh7G2k4srzpfvuU9zy8zBG1ZB4e8d8e4LNEYjK
uj1RtPvMsCGM30dCPxzxLVQhPxE6i5DH0Cz77BIBhB6CVrmPU9ROvS0jbiMSzh7B
54h/g6KrVYkRnXfZxJHEkPpfXmoeR2ALqv4cEvfl1iMYHl5k/ThL5EyuSt2Y98yz
+iJssuNHXcXZAxo21Pp1ls+EOJtTPT/nLKVB5dhHabdWUR2HgYHZuZgobt4KUZyt
clDpLYYFQk2SCSQsUlTTwVW1PJeAAc6uoqJS5Bg+q6YFiW4m/UDnvPDHkA2MtgM3
g06gVhcE8frH0VWI+TRZz+UtuCxB3mO/NNiUYkVXzduPtN7n9bR0UzSgFFcd25BG
Zzigb12olbv8KZjRQKMToxopIZmZCEPMM3F4yFpwwCGtgm2TQ3CQqmpI36Fnpk5+
bNox9L6/lK2BdKGLEWvuvrWvj+NbLVurfAOn7ZoPpBz0aHBM4zqAdm8Elti2E3ub
eWCtgWYL7OIEkEHkbUMRQUQLGpID+FS3CANNJjcZUqkECqyL21QHcLpWUSArF0qc
HOW6fiB3o8mirXONtVp9d7ntZFynfmkZG6SFSDlpg0Bvsk1dJ8APQ/y3dtBIzQQL
sU7XcuPxhEx5Q5pV3YgoL99wwvd+ctek3xT7W+ByOKEYzEMH08AdtjxafQG0VzMb
75S75va0dn0uu8SzDZsehDFUnm51Hj7jyLjZEnQetsej2dr7kY7vQk6Aq0AdWtmZ
9GI6em62Ls8+VIVZO059RqmCDCM432JEXlelM1pkef8TFRUZ7x94WDtpdLbCDVdR
mWLnmbPw7W379oDWM6SEGF6xcYrJPWr5CoIYs+nxBYvS5u4vTr98W6tLThDQN0n9
23MR/vIHsZTKAlQbPkWmErLot5nAnf1Hpodw3y28UgjfV71Gudft177efiWSDgfk
7MVf3XWe4oTXWhpZDVhLHDANe2xRF2f3bxaNKGupnDacFekW8hUKY4kyktpLGbAs
fw3q46FgkmxbKpH61k//8vTYRpx3xefZJdB7siLl9VZdNLkTuQSUX2LEbbVJPI5h
zhYNj8cNJlT8EXIfjH+RuwqpenJx/zMWbprTVZrWcLE/FWyGMjdYvcg+zmJ77P+A
arzvWIPEemtoiuVEF2kP67M01i+OD7j+HMDw1N07SRi3qezA46EADca5PjNr3+OB
QtMTryQAFG2zZUnHlwuniAv7yQDeScMaGbFEu/rWGDaA2c22PDF1iqtFUtnzRvD4
MhjSsONzl5UFUcFSyIPJ5EswatoR8M1qmGTlY2hHprGIwWDOBZr1W97hiBcEimhk
uW+bD/wsbul4dzX2xhZmdTTLGlQfcX0RBjl9l9ul/B2iz4LFVfWqMjK8htxsWSxI
1j4ftYF9rqVg0lLsAHzuvYNT1F27z9C0+0M+V8x7RfFvPBTeCl3MsOEeCKAJ+KCj
Fhg1+nKa/cbuWjOpm1qNFLNhMHYwJOLAYUZAuiUxbROy98sU8MxKmCpp19sdC/6H
ex937jHTHFTfwLyeHgRiDzbhIf9ixwUHFqdTV+tlYe0gN1UcKpxORdtkIjPhJX/b
v5Nbef6/33lo62QMVz3o66vqKHynH4Ml0qEsK8Mhq8TrCorewnznpp9cRx0fdo3n
27LTFoIYcvskLzwXMGCmzzqX95eWN9LI1FenygZTOV2lwF4VYcnCInILQB5MTtFI
bXXuxy0UMFA1rAgLzzQZIx1M/rQv2JksrAs/uWnFLxX9bZkhVzK6Z3THa73MsjKA
0C1R46PZOit9HuoT4hI2zrpv7ymys+4VQRoSkDRwAxWHIi2OcorYoiEAx6O0jugn
4MwT8+AGPGPNVxQHuHq4I8etqQaKIzqtJnzY+wBWruhRCrbctgwccQvzYRI/Ptv+
/au+aU9I2+CDJSk6DkLgZdbllbd7iS2uFD+Q83Yr2VsGkXERaWSmuIiicMbanLmK
Rn+wFiIIdOuLviJWIbcQyLFaxX8RVtCv4+1bSB98havDJrQM8rcMu7FeUS/42amN
sGHk4GazCIX4TjGMj2svaHPJikEKq5D08pVL2fMOFB0x9eFhA7iT76apKoNQvFuM
g7wkI6qFvZvvMle1V6FtnMqmP0Y1OKE7SZdcld619KQXCRwXqWSwHEzSLpcR/pGO
KyCO8WTnru3fE/cQeYkC3AV3czhsLS4OiQm/h5gMOl0OXm4TGyoh1e3tcYFsF/CW
enZT+/6c8L+uTrZWKZ1EEzzGc9/SESZpp/cdnSv1rKyFroQ2fftmuDQy4g/bzycS
S1lyxpwQzVSqpAbf33QjdVURr/7MdFs/pc5QzPcQXXzvfZChOxi5vF/3wrEoJ0N5
CMYqMOzbu+O9IqVowzo8jTmI8fKbhzHl56OPk3WfxzLj+zCnPGvOuGyxztparNZn
+NHEpUN+Ee/5IxzrWUx3wv3IIo6qZ2LK9+ZN16jK8w7L5CkyNMRX3irHcAHmG+eT
HTSR81I35VORYIwq8JdohG2DFu8dBj8fuUnX4RxhDVGEkllo0ix86+m7Mc1qPKCB
0/EceTxDWerLsfIVpeXi+qDOANnpDImSZfh7jZvSmeglqYTW2+wE0Gf2h9Ain0E8
vyFtxV5/Q+yHtQGsTwnrApXBjtjpTU8uqAK/VhpCRlTKlFTFkKLtVUdB21NOElgX
6EqkL9mgonuxhebb+3RZY+ZtFlLAzKe0d/mCZ/t5kIywVNqwu1737lXvhxaFXzuz
arJ7VwQR1VlozolPXJSDnzzHmWRorA+BUPJiuZUis57DlJ5AaNljDVjWlbazRG5o
bsIf2aySS4KtdT1EpzXijRJGpLDfP4+6xE5gYfSqz3wpfLm6tEqdGLP3nb6J7oB7
6sCd4wkaLElHRR5W2FSMuLPT/sSljefk++EvAbqbY0IoN0fEoAFGJ+pdkV3rfg/b
bHDuKFy9Ba5kVtnnQTqanl9INpbyNP/uETm2Ek3jv0SdWMNJHoxUCWZSaj8U1afh
koC/Ozrt3y3dHNh3FjTDbNUeJ2kAJO8gtSB8rmFzirmYbzqZn8bBjD63zPbTHW/n
5GFg+YOL946Ktr1FBm80EiyHbyXSU5vZDYgka7Z88b97rVjxfG3/M48r3KHn2DOD
fMG35t3WAR48Z6xta4aafIySiLREYh6XSXi1d0deazMb6BMV8Xjij6uoHvzXn7sP
BILewe6lFqlKKdOTfPnVakH7DEAcW0gOeiVf7+d6t2QQGS1FyvkzyBiXhkniN22H
u3nJ5iTNkaX0tsCinFjwOZ2AhiF9LoTM9NgihnJlaqm4R213djWgu95VLE/Fe/WE
buJWJcVEjUmYF2lPPvSSVdA5iVf/NwqtctDQy7S0oLLximymwDokMHJD7kTuySd7
Rh5aLMguRtk1uzUI1FNNUjFRzB4XKl8jxONZ5wUJqWtw1dssKYh+fcX4aJTgmffo
UWIpP3DV+tyNVyQtE7Gc/LCqQ+5rj8nck4Hz49WY2LpgORRK+Dbs9EuevASo2rKV
/dOnfLCDCdKgB1R01Di6O6BB7iU9QbhE2USocWfMKsE3h6rbvJ1dZFpiKNGraVhP
FWWVysDOW02p1VzWbKE8FCXwQmG+gw0B22fnAysA3k5rVqKlNuva+5k4+wTap9tv
KOoBrHoRpedFfgUEh0zbkHTkvjg8hucinfUVGPgzmXKogShV3V5yXTo/MfLU5Yiw
6MiFGjyr2Sxoi23/HHcVooFhjsgx0zLAPpSel9ofJglaaSL9QNvdp6AiAYQ2DNv+
vbeRWpk1VexmwnJLrW8xnbgf4sBjwfP4x85ALv/RzwiiFLPwTJbABMM6wdrqggqV
pc98M7pdzLkL401pRkAsabFgmusQk7Mpcs5q1IaDd42ks4rmsvKOZKRuJ7OVynR9
aiGPZSPj/Njdbuxi4ESv+LNmqO8nxKRG5VpqNYBZ5e2UG9SexjVuJFKRra1Krpw5
jCMdqZZHQQJYTpq2rMf8Rjc4+ozP2Ui6DQAH19fvgCf0Y+QAw+piKkpFLhG7Nukp
vcCaqz5127KmZYpRihJClSLa0ZNCwJw+htw1c4ZxKoEjJQ+oRslFVlqOxrsuXiF0
r28qU9C+4Se3t5+AGGOLZk0GpwEMe7lzsCp5sW1BtHxxiFr3txaHfyKz9wGqj28E
gcOToeln9GGe77b92WFxgEAazfHfl4n2wZZjZMzpyJwkNRdHLrcUdUH5IdkLlQP/
k63fdsoZH5dmogS1wnZf8NOamaN5PlSUBhgfTBgiLwKxHx60a1/bX/jeE0LqgKZ5
xsmzZUkut7RKCkfL2TcjLh1Fk9IpHFx+0vFD8wBRSnpwR4bK7tkfgfxF9KP9lYKn
SgBJkI0b9k9x34n9NPLKw40v+rAJ6Shm33O2ari3RzPaaM2ixL0DOj2NymdJvDLp
s9Li95Z+/FtYiUrDdxCtixnZs0XGwbNF60wGo3azHirNQoajhlx87cAOK1SSPS7i
3nSC5+qVOzf7/5vTmTYfY4Suf22Ohj91wWgiTFZRXsSHOQY3znK83e+97+rl9EVH
XO0Hky6hyhLr2HGOthuVGi8gKXU7hhWvjaG6OCC5SfkoNpknOjxL6yWT4x2StY04
ngMuN3LQrRmd9InG9RLMTiBLUpLTAgLthV2Foz3oPvf49MLSTZ7kju7Wcne7GPOH
uuW3sTpm+i5Cj8TgcQtXVT49D3Pr7ho7ZG/nUZePNnEegud7aZp/LUQ5vQwy3sUL
qUEvEvscYPrfM5hsordgy1J1U9ARNDLggyDpqUpa+YMSENJ1m1JND3PrzKMWaJmL
fcA1ZRQf/Y7ACwCrya0prmj2oSsehQXrM41htwfvWNNiJorE8YIWC7lv+4MClJ1s
zNKQcxBhsJT2i6cNnM3w123zd0dpgMeqgw0+Wr8VdM3IIJ6qarKZOCwV6/oJ9m+1
Fv+wrZU/vWK2q72A0VfoLjPXwEYyW25tC/d7hOuYSKSm1NkSoQ438y76+H0D5KhR
NVeFUd3HYGwvgBAh2LTabkQWvuLMj/R3wBHVJCDwfH0VXq/0eipxvjcLH6Gx92Zv
xoC6QjStpBW9JN7ogmFXmLoK4N8sGh6PN4Sj+V64hefJn7MJPEf5rcCnPRenC+YF
DAjqYjG74FUeLmVR3RIwohClJVFlEKY+ffmOpFStG5SONY3BNr/gXrX2bE8J9A53
9fNNaNLgZnxT74IbQNh33HMOGdCsGQTlladzbKHePi7iOji3IKF1DZzdpcOCn901
u+vPMN76DLHpnND+/RSsJVE335rV3i3cXNu+6NFQbQV0EdRL9Tp1NxyWFaCIzORh
sAsQCavFhbaKP/kwrQkOc82YC3nEstGK3MytvnGAQ6knmtY50vKPjvWBt3sLOy6v
/X1m1Urms1ZGOpo7s24U8DEbBHKQUQ8a+X5hfDffwNo/awEvfCsgnB8YCC0v2M7d
hFY4P/cTpRi2F4xiEZisVG+zQ17FtgN/yPSwOXy5J2OSU9l99+ngCXEgc1ti8bE+
G5JZ+yQfD+KawKhzzp2uMq1au8cuEYXOtnL4aTmCbIrDnJma5cL+eQS1EzkzXiRK
2DlcsutmrnirvHSsvdh3XBPFybIoObrehGjmtyDVvSmKZbvelk9BFlKm3hd13ofw
zbAJR8ZE6c9AzGQ2cjB91YH8ZhzLViB3uL2yRoRVq3fwRlFEaiRT8MU1GzCfS9M8
MuYuWTrr+sSFz05HJR3Re6kUjKCrRwjuowOcOeeEUUaw5d5Vsao0RjY8bW5dGPQW
JGpxE+ln4AxQ8PY7frnqiN8Ykmx7vTM0qcstSXc/hBN8EuhBY+3evkyMUY4+qkkm
lSd1XGB+qImOpfYdVBr0mlwe2VsjBkWDI+GSHbapByW5yKRVFsJYQ6D7GxY8y27h
jMrfvNQ2Sqngg6k4kK5MB4QoyOeMDn/uJiSxH5+QjCbZGZnnyF9/AU9B7EPXaqkK
5ywbcPYag7JAC7qi9GIuHl4Pi5UwTh8YYzTqvqBBNZONfsUd0GXUN/XC0jEuyAyj
pQ1EYmL067euugqEW6Qm+yxx32ytPTYcO4luF0kb4r3v5JECVgqkdUsCVUVQVN/L
LUt/IHUwRIa5hd+Hbo/MHYxg2utdIjIRbrpmf1Er3VQp4+mMLif7qH93Qy+gaqgJ
U+5G2/iglXKdtCRY5/2g0KGbEi+mpwitgKTaVFh/XQKYdyTvRLifAM01Tq5RjzkL
6hQ7YeUhmgHrWSCvk94HjCqF8iUDefHEbsVPgW0wCdMOSzY+KYm4mVn83XQaLIpO
Bp/6q3RCbpgmQuOnkS+5wFbctlJ1g/75bTMXF2yHywPauz3eVjonEhCF98a3B3Sz
8MykOyq/aquG8ELUNAfYQgCj3emabKg8Wq0RCC4plSxOqgzEt7kB4yCFwMonlss1
Mq81wkEu0nRcvjHm4heKW7KSBNypZqAHFL5OOw3wRkRMdvxz+QSrnksjsvfrh8tJ
ypbxIvqNTSiKZHEPFuzsWzsG72SBWdBcQ7cECHbakRqMtEkzfkxb1ItIpSF5vjRj
ew+SSbK5JW0NQROb4JJMUiBE9mQcoOQh3a/81ccpNPYWJcGe74+rG19I6sn0/F4y
78XYLdJ5vcVYNckjVVZHwoBrTsmBEhzeLfISQZrAy6ooBSlPDl2Xprul5tuGUmmv
2rYPli8WvhxQjKEK8E7YQ/cgz6gJ3B81KIEHQKRW3P0TQfjLWuAPqtfgXbTm9cdQ
87OB+TR5fWU26SH4zI+x8A1b/F7/k5J1vLYAVXK/cD4ClgLnI+Hozm1XQlQj3j06
ZsoDBUfdDRMvZZkHeVy6p8muhoxYaostVO456EDLhiS0au3b+pcWzCwuvu/bZqEo
9RGbsjoEcd2JSwot5H+kvTFZHD/9vJyMPIJqV3vrrNdvwjRs4FW5BnUxfwY4RNa6
lXEgRFLnRPzsKlBpnbnf1U91jNF4/ZciwNBExiZ+x8d3BvaGUuQpq+3PJlW4E4gC
ZbPDDwtpip2MRYofu+bUha8ysAqqKUSWO+8h0RVSlT6gDqjvznen+FULh94e557j
8q6sPp849Esxj1jiWf7e81wktBWgxz82dOPHx+06sU4E+aaokBtu4hDnbbFprKhx
49W3J7FlO7Kbibu20Fzqqa0Wy+OYCt/FvlTlNGt1Mf4K0OQMxbY8TkszxHJpkyxT
N+YkAxKhz7ybxBAuPmKaGucYMVtNJwf7kTUHyB8gZBTJQiqiFV3VPUZGW2i3E0yz
bx31X8MTF7pE5HfLfw0Q5V+gLsTBLARvRJW+64sgvq/P7Hn3XNVYlVrk3Qop8kT+
dyWLhEF5XNrZ4sWm6QVBZnbUXtbHHAQpwkvgYGbuBcDwjnATfbPrjTdMQo0+gDAX
3BtsHm1XKv7Sz1Dvn6F904D3HFN+2VDHBGd7rzvkdd+r70TLTdz3ldUnFGfg/muu
f9H6nfzUA6qVDbkpEy3zvihY3/8C1R7N9F6AODpAwRZVLqZ8O61I/KvuSFMFq5Fx
X/PTtWY+GDO2t/3EYjZii8NguX5Jx4vfysQ1Tqwf+xC4PkJS8um96gQalsfTw+OF
0JHP1Awh57RQACxsuYBfv1elCXM3WVneIMgwAfVSBA8d97qUH24kMEqUOzP1emQk
iJ27ez83V2lmTPBwiz8crJuDN2+x+vdDb1cM0VSk4PSzKfUxSmIPLsAXJmKEc1yW
t6H5r8SgahxuCl2S+jJjfkjW1MKoCu65ceB1PVF2RYAMO++9en3GZI0M8Cg7iIQd
ROX4nL9o56DMAe6NxKR4drWy5Xqsv01zcp9Ka1k5ECAMdGn5erdTAryqfMK57/9Y
6OFcOM27s8RrJJBWIyBrpCRHpbqqiEObk7puywn5mP4rbwG4pr+InqgKfLj7Mlkh
uuyLfW3Guob48PGgwgEdmcsT2jYIJ+hcWJBwEej1EkvEwM/H/DQ59m1GkfqZYI3g
6iQhiXnm033q8kdx8jsmFJhB3LhPEMByCuedtW+/7hpZ40kHy+jJLx9e/5TZ4uyJ
pvP7UdhagxrToSspPpe2oCpGKfCB+swpQqK398f1/PENBPAWQx7m8f3GCvuT2IUg
Mq+P8RSr5wzbnZgxxh+ZLK9gBxYXKar5zgf9pUTApfANmUqLo5ki9YpnafmO/0wA
l5GTJUh44x6y1tdOlf+UaWob8gZMB+iHNW1KEB6B/wqNZtwe8HG9/NbuDUHOHaNA
vzYIG8ZakxWJGuvLL8ksRHbAaGOtfUb3gT33yvMZwty/KSKJFSL6DHlB3Twl91uN
39fYxevh39ZoqBkapEzzgAUlfYi/zNVLGW0hi7met6DDEygffOF+FBT+dHi5ShS/
euAWHFDJVqXwfhp5r7qGFuuWLdsXU2+XCKQSMJ0pR2Kb2rupUWXeUC1mOj7hX7MT
ah7Qn6ZhzvFQ+iTpITNmURZ+j4Kh5oXUGtQa+lUpqg0ck3oWG8WBKFnO8Tm3WQMP
6soEUrj/fswZnZtFw09dZ5f1d+lmwqYdLy2LI0upE98HHciOlvhm3skpmLTlIedL
fjbnJ1jX69sxn6w3SpUce20+plFJh5i5g9K5j/LEW9fYRDETb7rBya+4LMs6Cgfp
qT0fMew80wQ3TAIiIOMqgxg7Kp9UjWDXYSHSoYB0qat0K2VC/I2H824SVvQru51l
8og22UYJHLFTIAILIl5q6ZBNKvt2j5PqLN7Asb/rXDgZTsPzw9y8jpF6N4uh5DJX
8/OYyVrB17M0YSiNviqcxSTFbKDCDChLPpb9iY+l/pcstbfV5W2K2o0dWw5GUmHe
8xFByXU1mLIN59b3k9wYUsCUWqbNgtDQyElcbgoJE+FrCtv5AHlCeJOZEHRq7RiG
Yjn0xne/hcxkHBemRO7CGLX9hjHMJfWgs6RZL3WZXocbvvUwnSCPiP7M9+yLdzgw
5+Sk3pWonQ+ZuWC9CvsfukqYsOkvGo9xpsO0bLOqvh7pWyW6RGbDSoKR231i4Itr
yoqYjsovGlbNUMKgEAVmhYRC1sX9YHswRm/WDXdiauz9GYMw5PwDmQNJyM3q2WSo
Vry730JRHbaib9rkU4UBp+0IUN1acFtHXLOzvwWURk0fKz9B7K9UNB/aqHD8p3bg
QIC0qgx7XduCjO7DrwIFH6RSNzImrcp6zJ5N0zc4iQhwULnTZ/Jr7xDTH0vXf9jw
wGL7Ji2guY4FfEH59PozGzTUqY4l29cBri11Vy3o2iNjXUL7783jeuYp6mcGzBuB
eHbTJ7xG2wCP140pqEadLI2TIvNNSacNdVZ8u5Tsi2PKhIhrzmpAAFjXlYCrdlaL
BxFdZUQKrmgFm6gGmMZzwSWFmQlimk2g9wNve+1lSxrggHKE6sqAr0Go1Wsv++ww
w7pqICySuqFs+OrBoOQa7L+E/jvdwJRu7TebNOk9/BWfmPk8uxkq8EmF+hEQMyaE
BJTeumjtt9BVHqth7Xi9PHcbLanWWI4tsRY4O0HJ/FeEDF1IAR2bcyGUmJSeCr+2
SCS+WTvXVQHIRs1OzzBKyRi2Ue58WtZXQjrHAb/CoDg/elB2LKNYuTAEwLN1/sMm
+9z33g8byC0ddYGwf8So/7TPlLRnSb13EGqgyYfAMkvzplW2G0BmUNh+gW+3AHzI
vZA+frSM2oql+5ZKviYfBTIuIFgZQgKl+ddTIGickkkSBs+ti6aOqy7iCkT9F4V+
yhwFzK0oLHPW2Ukm8m7WAIpeXo2wqb5mEfd292psJ2KxnMkizuKbnOUWwf0VQ1el
eQE3PyhpQfY3UswjdGbvATxex0FZd119DZwG5yH9eg3KPs6SyhF+AjvNgGGzTTq0
kvA3u3r3W6/7EJ5bTEppH5r2NfFVJ6hf256WTEWjXgw2H/3NPFzTk4TXbQlq0pxh
1g8XWUDrhuOTRswHkaNnc/DMXscEglct5E12hI528Ld7rj1nwXzW6wDilL0u73xo
Pt0y0RSlLyWJzMrG79WdB70Yqq67MfVFZ/nCntGYRs48Z5lVHgMp5jAZVdKzeNbv
kFD7xFsLHP3yv9iKFX7k4zZ78s1nU9tsRi3epG5Qd5Ebcv1zK9V0dmaiWwBUYZbW
hZlsydEdXaRgtdYY0qnxdfxWlHnr1gXhDmT13skGbljDKe53ETPlZWima75R3pgY
s+0pcC581DO57c/ymQHrUZ8uBFnDKgEoVhKv6haRr4dpo9td/lPFb1eKPzVXZEzi
TOrR61LWpMOK+eAskhrhZ6f911A3qX+/sa5GyLnYDg6foRf8oc6nQYvmS2soDWeH
Iam3xTEuXtrytef1JBllCX292HMYH7HBxkG4eAqSH95G+Rhy5TR3ecz89qJCw0Tl
6fVmTuC0IxTKq3oFNaTC2MeoRXfSLH/awxVNlVyd0XXo4LrRt3B9sqiGSnR1P7iB
7Ej/thEV7NYkRoUviU8BSJStQkBEe+LdkXlZijo3oIHxUU6rLkd13bhgBxRsPf2F
RcYhNQGq/x1JVv7F5fmB5Ygeuelt4zeSvRNNhidlakoVVC5pgnycWqlhVCbWaxO0
97p7ms6ARnuG5Y3U2J1o6fSWBdAbXDIt/kp4pW+3+K6lcUODnYJXD/JfOW49ncgE
He0rdkL2MUCsR/ygeChKnvqNhtLpmYg8EMR4/PqJUx3/CqQkx36BpR2zKBm5DabM
OHw/9LxPaN02wXSfIgXcbmTD1Nmj3GqnuFTZoyPkWYZS3rh8qMc6/EuKKizM40OM
Ua8gr7sLQW+nQVbtWv5vb7fsdd3pCMYQd5e/IYwB9qo3J85vY1KgFPWMXeocBCRE
h6tevehRgvROUMvttrGcDVYYnM3tH7dJLa3+wvUIJMggwd1ypFKU66zvaBtAhjI2
4uc/SbmCCJjVOgX0IYOGMm98/VMwMHwd0MU6rmwj95HYYxPTVCWGZED+tNe2jcFT
GY0gcQ3DtY4cuRVvLbOWCQ4mY/zay29OZuKPHsn7y2p6LN1ThU6+6hWxmyDMm95V
Ww0AnRYJ2tBPCWH6BmAB3qxsPtKj7WFKRzHbvZybkb85EURhmhFKk91+gjzklUsZ
OPZh3EnqAVkuQR1t4NXE/232U/LKwg+HaSTXyzB0iCiueJQkwrkiBhSnIX3gPbiA
HVpC0CHE9FSnMBWGTeEVEmggexgQlZeO3E3+IPaafcjL5pG3c4dvhtTPrV3ECVDN
IFDSKx9zKck+fazNJlSWgSQX+UvuetS5InPBmpM7hUdTFMq1D5UWwu9wAGfJUO4k
JraJsxCsVwaYv1NHFyFBBuKjoP0lyB7srzHXCvzcC3KmMDjK0rUla4iZ5cKggxcS
3gFB8Q+liLwEJZGvOt+BSBYh1BdqiivS2Vcoz9KKbR8yjn+e81C1xxeTC5OD3OGu
X0rcW3md+ihyXnK0L7n8xKKdBaMbGCYU5w/uIj8f8msRV4jyLK9UWt5QtAAiAzc9
TMQyG/v7ZFmfCA1OCbODYTgFmzMiHTL5BuPO5ep8PDVIfIXZ/15wzmJZNWpkXZeS
EUtQNohCNReyI4iGOZfnBgYESunKh1VfMIb9z5TsWKOvBvz0ZyOOUl7Fp9NPB7pZ
8S18FdqRUgiuuMetTeKm8ZhJ+ufGMa7ZfrLMJRIjT5b3gaV8jlWRHjBnFyobRCCJ
LA6U3x33mvBcxA1mU0KKmmU6DTTSvsMkGEp8WTT5A21ooNETFi1091XSj2oOnpF7
3BYGChv0UfDyNBdpA1oTk5KQpOBLiEfSoy+uGsU8TSalkgzelpcCJM0cZYnDtRgG
e/FyaT8vgEF3OfqVkSf9MhENYPGEoUEidYFbC7gKFzZ9eHx0eM781GAKqF2nRd1S
/qbzh7iRGYPibgBgG8ODTchwD0hb+9n0ANKEiJewQuQjERIypK/V5GwGUtg5V2DB
AT6JFcY9Ki/UUgwUproCXjNIBvwzLvfsjnH65NAwP4koBR5T31u0b+PrwrVdtz7M
2Z9f3CjrlUY2Ev3uW8KQgG65uOa4wlXadfiF2DeEEpRPVYeXgXktSQFv1zFdNTQh
BIpuWCWSt7rlD7hUwsuBgzaJYDuS86dbUxmCkLE2kn8JCUwMSkireQbBI/gOdFr4
3XqhXEtXa5gQjhKAEmKyr0da5V5J7K+0nTj4WPjRV5DCPsr3YFIvttsP7Mok2nNy
/9CyZoG/aAOVdX8JIbnM5+Mt7kLeH85BjJbnKgyHh6Pd4MalcFW0hHg/AwCyFPW+
Lmrm/hiT2cHporXXkLavIxhMHwimQM1mEOgtMsqWFpQLIZHEcVfpmtZuP8JVh3Hl
LZPFBthL+THtS+TyfNYX4U9ibAU+ukTjyB5cWWrKPkjNXGxLq41AAytAFfjdLehT
dH6TDGDlT5aZX7MEwxTLMRvuHFfq54b1yHohCm7iAV2QTeihtnKiGJ+vbVt5jKWo
fCzXbviClgajZNEiYe3b6T9v2X/rgMOFWRtQ2ulslEfuDEhx0QAlA23UpZxAc9Yv
ZfI2EM6fiYp+ndwQcL6TipWJ1N/ckZYioW1o2Ci9JKQciKwjMwHzVyXEmn8i3YZP
jToZHMMdgjarpYiaB7rH4PdGCfNtKwrgRaayJVHFrj5ym7v7Nt4lnUz85QLmczQI
p3FbILLc+pU0cutYYei7+gwGGMYDVUtzdA63BhTLBsJD/9tXrNl2/yqyfCR5tI7Z
gU4Gt+2ERrM39HB4pHlchyjByUmr/puEjyC4bpIXnyil8FcO4JQJHT32CcRGHYwQ
v1r/sf71+Dc3bSQN1IxJcF5xFirPX3rPytEq8yghEj9pXGWFiMsWBIFf4zPWZVtp
YK/ePeC9kKftwhuoUg12mR/GWq1K8/I1iKHe/wjSo/RRTPaaSFbFSN3owkBrX43L
ZABptWY6hLzg90UgJuyls5AU7hIP3d+n+wp+fXe+5GsOVvBVmlV/DesYCGhXzdhh
znLmbp+jormNTXuVQqyA2fe7v+Cf9NVQpk8TVPyVAAjCaJIp/YF5BcQPfAAYjvJv
SzWnmh0NxvSOLYiDUY/K+Lyqbi2I8v6VXRHVXvx8xIIj3sQMDEULJ5+utzYuvjvg
xgr8G4dx9Hi96HQy24jkaY3WNFjT55aXqtJU3NlWYgMh7IjowwdPjVMsm6pIx0ol
MKMPEGT7BuJBbr0oEhh6EmYPTKzglr6MXpZnWcC3YzkFaIS+zNWvhq+ur+KD8Nu+
YX5DH0Q1NqBoxz5t3JuS7zpF/0egFRs9EC2d1Yb6u4FGahw/T5n969DWdS5lX0Wq
XLWJ7Z8O93ggqFJq86AMkcLKWiOX7wdjcZhRUEiBnVJ2q/irVuqx8HiFVz00GDOU
lRCoeOkT/fTzUM7qVtvuemZOWyl6Armgut5X9v/PH9ynFXU1NQjP+Dlcoh/7z+UD
5YfceRQ9Y0bnf73qowRyJ6LK1/VC5I+QlpGfIeA/qkDVToBK+mlVwkMIO1QlzI9Z
WMym+yhs1wTP13ggg3nghKfJPDJ8UjeD5vRZhprag1VX3v7mJ/8gxFoUNyS7HpZy
NlexVZT2M5bzE2+WAN8P06UWNdCC4ssM2kiFDTubdd6WqJXnsKRhB23byr1z1e97
gb9QVxY6LzscjvKvFk61rFnyH8oCW4pvOa9PIPllu8/bDNSyfcJRwQcosNcDWVAQ
d5pnsl70DOHaeTFmeucG1+ZZzFE+51l6Tod09MxYA+AQBcO5B8pZX7vULRE7tsSd
cSCXwwrHQU2/QU5dB/Kxw+A0VJxmjJqMx+6rOQLeQjLF1RhoIQsi/c/DbgVUn67a
xzOknYaxewcVSMfsRnGTp0J71UEWMfQ8HUx8cEcklIRqizzsOOy8igybR0LBM4Z2
b9FQpMAHq5ZpnRAZpYA1inZXRgtfyFgnpC9iAZEERi7xjKJ3K4s6Y12sKrPAf/yZ
xobCNLZkZV1/wn9I8EhGNyowb4Ee8jneLfXGkZ1sq1bTzFbX89IPuI7mEP6E676k
9T9uCG7W6azwQyHxE0MkfETp1ilj+TJSWotTgsfAfaXesIlJo2fudijFrfaqR4As
QChhaxCEstOQ5HNqaccUxqr6BdyMT9FOteSxnwSzl9v5P3lo7erxQa2d0pWv5CVk
/PdbPH2zeqARXveMdga2DVroSsJDu2zTsIqg73zi+l8koKmuPHxyO3YJaUfvsueM
27qdFwLdssRcPAeumJx5mJeZJ6RW9/L4mNGfKCoUpXcPDl12T//nwPlWDPHbFDXd
moilewBbKdqFNilE402gQZW5XFaSRJHzIPKksNLj8fSJnnsV1Q3dUv8x8YlOKffv
dxOymp0Iwf5+u0TqyA/QNVF/TlDu0XjxAAEWG9PLAsha+CzofwcATg+SVikI4lIO
e+pZ+N67Q+yxCruTrUqf1s5KFi3ntbgGZALiJMjD6o/0mYzSS20h8b4kP1Z1tieT
laVZC8SlRn4GnUwgFAZ+YK1PMRCSWs83LiekhQNlcRy6IfeF0r4ZCLmkyPoYP4mL
YQNVpLT6M7MkV6tlqG6J3AWNByVZffqtpsUZ1y8x1AXhTmGw39fygpemg+tj2ONU
f0HLFkJG/GPqk7SNyE31+/IcREEisThKS7HgA1eT8oTr4PWQoEGfX+lU12E2kNCO
LQLIqQoLMdq4vBdRQUebSLtAy4pmJIoGFf41ZB97ZS5HGqBpaJWi64FZxZURzQ07
7vkJxJGSW/vf5k0cmd/EovL4cMAXJht8dE0PjA9MNSGbM4i/YnXZ/DYnsUnfFoyj
8XgwlMN0EjmaKNkb8uYsGFC6CvLVBU5sMgf/tJLSAnIBaEAuPTfXS010UVI45Guz
fmjGNfBsU0SgFp2M3d3TbV0mTTEKBtxCyJoddHZlRLNCWU6qsiLWB+QzbbCTB2WC
/F0WITZpwPM+GOlrFYyS5MlWEzWGBpHwZVofPs1ziZzNiFudMRZ2pSbWy+RFX7oa
0hEkWvigBW8zQuwKcl+xAGqGD5dZIKRaWe63C49VXAX1sRScHU73JVuj7K54VrQ2
kjvVRToGtxLITjbDcrHwkxnM046k4w2/ToQQAw1SduO1THd0U36DSmKomcG9o3ON
Ik8iPzuyXPZckwo4ldMucJVFOseAdP1U6Ag3ecBMY14u6Q8jvgZQe2KqOH0twNwX
G9A6Z/ORDYpJVGTO++FCghmN/ZMP+YI0iMmAcXGAsw0Ps8/SBDdUTzsN8LwHjxsQ
c8LXar/JMmusgP10i+NFLAKcUIOwQmyPGUXUfnUw3coh455SYFWa1nuiZrkGxYlJ
27MrJVdjr9r0b3rfkHt+eY38LxMPW53Bokl6HXNVYIXnth3BPEBD6ik7SyJEebmL
rdxccJ3h4OehdAUN/o22GtIUG6yfxk+TD4SeUcGjk0tqXdwvr3/YSUamG4ZhAHt3
TqMobWhy1c2dzNOpMPJ+VqEqtd47LjUxMxdEWyDHPF+JbxZ+NwqAsv2JITR0Crw0
0nFCxHPrdLQPvShWlVl8CzGWcd7WrXlcuD/HAVyTixcrRwdsBAtcNLg5O8VfHSqs
/rfDHD1ZfVeKQY/JcEdidfHP16wnkfoF05B0NYYeGOj402QsNeEJwY02oHViw4mk
CNxxfjmYes3+TdRWg3CmDsHzJk3DvNv/YR9rN5P83zDZ4sgyq8CgYZwcwh2VqyWq
1U/Ckxi/uTcJzkFBzg//basFGvn4PtEMRMrDd4y1se5bs+afw9ShlpTM/aivHEcp
YzcTcxuswl3/Aun/S8OHkaTK/0GfTQBq4lX3gux1/6fHs9m3AHeAB37mMBhoduVe
Y6hnzI+aCTZ4FX904WhjyrSrmpAczGtP+wGYKP5kkkFNBLkriG2plNTQMU8uUZSw
1k7HAMJAwf0d3AfeoQaPqXsf1GPKpx3133uaWBYZUw2A0nk86tM0xzdx9rlgSalh
DsZ90vivIu9iqdKVe6JZ1KxoLkrV+QkRJtTd3yXxEHgUGw/DAbJIHsJoBMdmT6dg
Hz7tmSedEsFcblN8oaNbGCQZLZSU0vuOWsYSai/l5wOiiYRlkB7mfM9c455Jtd/6
0jzccUn3Rp+i7CDjPKI/NUzBLqJ4Of/nhYyCNTnFoqz05ebtbnE2olYINF6USpgZ
47MvT/xGUfb9YKAknTmpsg9EqjyjFW9v5X4iqLnPVh9UEhBIHute8irofQijW4S8
P8EKp24Kc9D1G0Y+LhH04/3rlKwCvRzvOtcDF3DkJWH0KBFy6o+D3jzn/E2V5HGp
ti88KxR/6tovXJvCxtIQoVpPpnJFgPw/2Oleu2lAo8xMo9IZB/ig1OsNjwIJnpzx
lHRJ3yyIEcuYYwf/nPtxIGYxmWGlkjSAY/k+mUjE4FtjFhC8Aup3KV5q8IkfH6wE
R61OyOs3YnrfXwqZq6p2dXtPfnW+0vVwQpKqAk89sUVRgOG+lYUr+8zPUpvubMj/
uLYj7iwU30ZaEmJeBiARYMXRTDHIQ48omrQW+6LQMFmD7FlgJiV+lokyV/gwuzr4
RieG+VWq9FxEQjpGHpf5oXk2KqiVaBjceaTJuzGV34XQWupiarfjNY5kN5K+5LT4
lcnOElpllo9AG3hmD7Dr3qfnCWB3NH24Yo/bCer0JSMNN5y/h0MDj6NaJ4pvaZBH
m+r7tTERiSqyEJq+wUd3GTi04pgh7LvL6mcf0A0hrwPCbgII4zcBopF+/4LXoe0B
hZ4H4nma8Iqb71ckgIjAaQLW+CcvnMWuDiRkSVjtOisEW5LnSrc9hhCKbmMe22fH
Gj+i3ux+1SlkuOBLHKBNIR6QkpSFhZbk34aA36nXWWei6uhPgMgIMnPckEA/nc3P
fh6j1RA7AwY1N8/XVL3HEVhDCnmmHyA5JwtggTEH6MqlxTJoL1E5wic8saoPTKYQ
7nJczQIZkfuUdaIpHd3FBB7MscftfVP/EzlM4/uD/AxbXV9OItbeHHGKcXEAwV+9
t+qPV4R7E7825mQHOj+0VnDa0c41tOIhTP2WlqrhEPLkstBZ7fC3TxjJtkr7PS2y
170AJqNYJLZJepogFfF9YcsPQHCj8B64OrlVfa1tc+7Q3LzyOkEng0iZKvxvBW4d
HzB8sTNAinjmBQ/4CsXNWY7tvTatkhB1DD/hgpvUpiNmcFolm8r39roQxvl9Gi5k
0K/VjiMRFHERgEgEUB6Hl/rMl4Qtzn9LhWjByHOTUYRrksbEp91tke5RQ/AN5jq0
5Qt1MQXIiLBjtMRgftbbb+fegf/4AjbMPAkTimZS+JLoBBSMoTQJZsFscC/JUqwa
9ORwcc5fW29ITnjKhoOJdrKsnfiXHRjvDXa5IGX/uLet4BmVv2k4pCELzyZULmwR
QWj6PxADZ6MJQbDAGY6mQPzURIUiEkkiSDSD+9/gFXhDwncySalAbFgztZCQ/9mI
JY1X+uVeolgDOsWVw9c7h1yLEDqc606daX5fkKqFd7px2DqhUet2288h024+r2WS
wgMKo9UnjEkxlWD1mpyhr+OUUD7VTieT80tqpWNMUEn4eYtKvoqJk3pSNbtp2HF3
siDcA3NCddjCrq5M7GgAZjIcIwmVAWwQrANcO+hP7nQq4evB/hV1Lz1HGJb1ThUl
cWhvZWfESBPTVV9iY8mVyHuo5/6CHuyUK49K/uoAwcX/HzPE0vmGK36NE6/qAQ1V
iPdTEhibTseVJBubDwwfWAptljHzZA8tsCr6Jq8UvChDuDmUhZ4+t0B0vQDlfrrW
DLegJq8t4XRfZL7NdQBhJZxpIfXvoBG74LfbtWxEWRYog5RbyIo9RqhuOEtQ86Ej
jR5CQbZuvROofuZtrBJ00xAI6VQCfc5UzEI0X+6URfhAkd6jKFZSE7YiX4XemIVb
glUXvwvH5GKmj7wiSOAxrxuHJbA71hBUNEM8Bzp9xUAYeaypQvAQiOlhtpPP6KN3
5wjs4taDNFDUszOurORCjFljn45osDUnzEWkfC2nB5ZPCqjI+RnG8KM97Koxn284
KEe+fBtnlrI6SA3IIXCu4DDzKI4doA+xboKkbumUxDCFEXED8vatymkRODusWXNN
AwnBi1KjpbcclcXVPuRt2RZm+gPyjjYRGRZgXb4Txg4CDCH79qdKUwb7lQ6fuXIW
CvEDstvGSlnDAt222tVk334vEExDreZ3x2xxE1P0+5UQE2q0tJkQa/u6j3c9GiAI
Jg2q/OxrM6OLLRwXYuzDY36fEAZEwZLbuCMld8aQxj6dAivCFpeASeEUm9YnRuBz
TjI1f3gT/jtvR93Hf86SKahf7pZ9XQT2XUG2jlxvCNnwBB7xZf86GIXwirz9qxgQ
G1Ylt+VXeJnNBpGEprlD0KVVFIG4YwJh2BCraCnUiemPh9eOKDE0x+qtO9DI33zm
AeNlj8Sh0AimKMLJyYfCjBVcha9izFx+GGme5oobPWgry+tZBRaxM70xMTuL79de
6eav34LU5G0SHMVruKmcNyCDk8cRTBIh753l6Bh+BD1pl7l9Q6UtdYmiX4u8Ey6v
+tPEW5iiJzo94q08/KqFn9Y0b4LNu8rUsUwhlQd//8yM2aNv41SLpMsqzLbUJS1T
Mwq+dveVEgEEp0Nq+9EM7GtwuymF6bQUd5kv4OArKLtZnpfp8LxA9o4BGtXfUXx8
SeB5XFpLc8qD52+qnBGH3FhSck43csHcRUVU83cYMFXSdmkBEwI3bqtVufVSf49v
7Ugk6ClxVHkJKhhFuxCDZ/G6WMhzM873gYXxSj5tJxtqms7YSDWPa9kD6SC3T91m
IdSdsBwZ4NYfLiAyS5Cufuov7ZB5i3Fju+T7xxIn6ZlU3X7RDqik0PFlon2amGIb
eoBXdwFp5s5bM5Fqam0SSxpbycuhezZS8YzNeNfc1XEUAMszXIhxxR4CPIm8JhBM
TAiB759mmWQZcElsvnKCMhNHxswr007ulbAFFcfDLodobHIztuhavAhr7TzJbegk
HMB18roLfi98yqhhIELSurN3Cwpza5tYKM0Uzy23Bw3F21mWxaa9vtz7ntA1nzhP
uPLzsVU/Cscr1QGYVQTEW2inWlnOoZmf6oVYNuomJ9P/Zaj79IuPwiTlmGupCPis
lSGhy8TJbOq97ZMe1cZ1WW01YJd0VbG2nCvWaV+y7+2UechVKbzzTZ2b87yUEsS0
z4UM5In68hL+PglNTREZMpPoEV8/ek9y1BR3CT3/dEy2aEBsESus8srKuXwpVdCR
NOslzBMFdsr4wO4njE/x0QthRW+ESwtdesoCIp5KATDfPQfQ3zhIzHe3Jn7xbOtr
zGvBOYVDcrrwSeqX/sBw3AS2f+OD4jPT3PCL9jnxf19mE1Cf7EM79Xd4ytTya+DC
1rx3dOd2+osoLCup5TaaOgGyrsAbxH1u4T0zHrwfoPk9HKWNoyIEb9jpU9qRt4lE
LGEIrzKsliP+deSQrcBTLQdVMRR8joTOqyIZrPQJLbLvXKRbUdcsN3VWyk2TPWxt
bN2yKxVvlhkrbOsQdrdTVKttWLfy+FqFVKaFz9xyxFJU6O65JMpOYl9cNpsMmZsK
NQCA73zJNL5LqhoA9YCHKoCNsiyJDbIfxLKSTN6vEjvXsgcQJKN1twWa4F9JZL+H
mSQUuFov8+gQlPyuVVGWRxyIY2JX0F7fFaOHOJmIOsEvBEAwXPfwiA765HtISMiq
LXF9IouRinK9Au7dwZ/vBNORMt6/7uHxxzwVSnHxjhNpmbkaNDqgLWs60h8HOU50
ScNQlfRv9jOiVVWQs1egCJngTM2MesJfFp62yooOuV9VqeVM8vtERleSlJvc8i4q
hFpGWKseMA/V1D5WtW7xinDrDfBiLCOL2I0mRgl83cS2dKtgNUTNK094F/lQIkvP
lne0EbrEl1W3HLF0xmdsM1FnGrVQ8CiMT7EJGqgW1aVQ+EAaTtEuxhSrs1hF+Nn7
bnvtdhZUEsfmYWH5XOEwQXi3Ul738OgG5oI/HHTfCtjpw1BbeZ/Sj4P41D0JYI5T
7QXTy6Hq8JqtVIaDOU+1ejGEBrRoixGM0lH4cLqfyd6uo6v1UdUjLjVcKDJAqiDQ
3Z9bLcu71GNAM+omuItfCH3TpLyGsv0uZ3z7FTunWNJ5SOGSzpuQKa4h83uU8yXc
l2amGyDYXJkGicsQMDF2ym/jitsauPtWuA680bA1SEkGJKs1NSsf/gTAbpZoNpba
JJSN67tB5aVLTRQ/9+lcRQBHqwOomBv+Ug9Sm9aAKW4IX9eW0su8/bzVhujkuxSs
UoNYWQ0dKUUyZRK9V+W634sivyoHr06RR6VaPIxeIStm/xlxFlyUI77ExyWKcDQj
LeELb4ele3AFcKbQmvN06THGTH7lRSMEluKPCdzCejQEh+F/pEj1A99/4pcsvW5k
gGlJLXC9KXk4DT1hV1zy7v0XCTBfPFe1uEPvLRRGmt+GpGwUvXhpKBicdl1O1JVO
gxlYfozrArsCje/9E87/oR5wceJKnxGZm0uFiQ1AQTbkUWO59eU26rPx630KKjya
vsCn0kj7cpaEUQH4EkGhfXd5MGXtATAImAhInuKQ5zFlKDhr+dL4nfOxSH38o0Tu
XtO43V6B8juMyOZLDBd92RN4QqeqSHJo82tv/Cj7icvFOX82vP9MTA4EQ55Yr8lH
Fs1SicRgH3cIGivKtIHqIw08cP9r4SPyLf50XInzxdPddCqHlI24qaqzh1uXRqN5
cHZ5+Se4dVYc5OO92kyVXq7yu9QVMS+aMWopge9d8Y9skm8XSLpupiAZ1cMRVwV5
ZaaH0GDdtGELu3MZbwoLVZKWBtQbhnNmN9l2NinqfXbygy+Z6Ipv237V0AJoNTqz
wA9fzB+KihMtYWukZRkfTTlNLWYoKSvT3IGUyRKcDMgTloJSupKCWt5lsQdY84HB
BxDRKV9wKRs+QnhtZXs4tkTM28lxA8LtxiNHxgEgMfalgvH3l+QLDBiudvuKgd5l
UKoPhsqw7E33eobzvRe5GAX3cqRLr7bB5MUueBZyB1XMXQsQp0v6lWjjSh1iFaov
/8g9HLMgUteNSlrsqLJGzFnBJO/WAj2GV6cTT3cD9jLnkhOeCFF9Rumz0ip1jB5z
LJWNBeSnHLOVW2TjxVjyZeBhF9YxpundccJnVpV7Dn9Z2E9Imii5iMwjgdRvGCVO
w99+LncRjU1CZj4eJVs4SPoThSF+2voi1CpDzdkmSN8T9zcMgL/cmK7YsiFeGwbr
gMzB8+rv9YCXpSy4Jp8ZbuzX6eiC8d6Y0hjKBUDWlM4keytdA1QcUqhHkxIsmYzR
4uY28j1VZwebRbXcLxVtBCMfUXwmo57AAgnY9pb9vgGIpYgN9ga1yAL/VSA3+3Pt
WM8MOJ4pW0eExYEFVjdy7z8tRy+GKjRSqEWwZXaOxu8OrPT/vgkwnPcQRTvRM29j
aqZlNzO+D48UHI3tFCFy/MyA+JF84s9DhjgTDzL7SlTSminoDSaWLQ1GtWV9PVBc
YKgl5QphNG3Ari9X9apqKWgOLLhH8m8XGaRCvn/KLvoDDHFsd26UCwv0KF4UBo4F
mQVC/GHe/CkjtSZ/EkyEeWo2HPV5k3q0SMUNJvbVxiM//4TTXSw+nUqKhf9buBvW
trxh6zbFq4jUGmUIYi+ptGhPTiC1CFm+sS9ZaZehv9xlEh8x35vOw+U8dsOWGpI0
Qej+GQGcI8VsMK20LctqN9K2Ze4rbNhJx3vr2rWfW4m6zPqwYpWQAPX4So7lud6N
ZYp6Xfur8kjTTEJ24Xme4+ubybgyb5TJ3Ax/oKi6Y9XFsDwAy1cQoaCdYrxtQGUW
y2n8TxkNG5kp71gpQfKuW9pSSZ84oa2MM1D/NsFZLNMbNKSV1SUnjSJvgr0hFw+S
xDwCvQGh2JqqzXO/Cou41iTk6HeVsYAVypidyUPBxXgZJ8gKqdk4o6I2n63+oJ5h
SlCURLj3X2FOrMY2Wl3X1VbCyVA5YRLN6kva2tM+NmUh2jMLm9MDBoRMlBjR3QnS
nNfL6IX1h4cmPFReuGePoOrPCYM97odc6oQGTvSsPfeg+rMluYIhOsbmue5h603a
Dq5FHrm6iG644QFfkRVBuox+00Gu1JvCefiGocr6EXhNjGXLg/UvEfi6p1hHkajV
snSQZ9UG7A9yjBaeBxaAwn5O7/FuPORhYOluAq3K6GCTGJpAGShFuEEvuanje4/Z
B9OGD2rTfhJAzdeMoF35Sh8qy0IsyBLQ6B2jSORqgB0LpLwAextx77mF0V2vkDDd
08fOSBfUm5jnZXwn6rEoZoS03+lf64zX/JGPPHxq3jcr3ZMSUYGQkHYNh3iNYszd
PQylDR8m6Tu33xSmTUhUCUECxLamgv//pkO8u+0zvHET96G6ppt5y8TNZKp6+SXH
1E1dlPBZZYqVO2hQq9lmSaXut0NscY8hjRsP5DyaLuPdDegL78mlUHasiroVL/xV
qW/CAafpBQSSrxoR+rUzZ2quBs12KLf4ppxXfv6vYxf36FxIuoq5LmjM5isLSEMh
eV3ZhECAgh2C/AWd8YcJhkPklzV+hz9ibmZINaU+qop3FOnXNNjbALsp+hwUZ9Hp
6kXj1yE0l8lHgU3eox7fWyd3FwME+6KJkQQM1soAnIQurFmxti3rBzTgPay3Dumw
G8A4CsMj7Ljc7qneBfMAWUND8a3nJ7PsT+oSUm/rYz/v7URO+xzvWCCkhevPA2M5
G1Uad6k6OUgFI1Qy+mtDglY4cLb/o9NgcoiyvCXuKGd0Btm75WpdlK3e+SsJSzno
HwQH2sPExnZjK/EOjeCdAE7eGf2kig9K9rpbOIHbuWh6A38yKeaMhYB70TZ5b+B7
QTi0aeW0lfImWFWjW/dEaWOQSGxA7tZgspEB/T6zGtNXvZr9clWFdD5xafQIjU+c
CekEsIhEeXXQGbBm94d0FoYXCTAPL18FhIU9EDU7oI5vMjIeZC02dAexWZnrnv3k
qZI8WygjUaBC+hKwMUA+4PI3snsm7Gr0B+OXhxmFlhUl/EWuwwg3RzzkOea61KZJ
CuwruY+m8zALyUqAHWlFmMSlYtoe5qfWVqmL4ac/KXWh/v0W1/stoeaTV8e18MjZ
aLdQkVnc8fvc5zkCh3M2KLB6g9HFU/Z9RES8J2Iz8sYqCuw83olt/hovgDNUnYeq
m14nbzIRKV5nnhFyPFZnhEV3SWWEUon7hc3W1EgWhE2+sV9Mh39c4ULdMJXUuqVU
aVhgP+q+3aOtf9YC17AW+XaxBbTVvXGcHsKvGINMuddr0ivoELJcwk5TZr1XQ9N9
BKY34P1i5BDbPrGZY+mnyRR4yq+4n+0Wu70h9QR6XpWrTlWT6eQwrvs1nT/PIn9s
suJ0qxYVI9Oy9spFDz4uUwUmGHxTjh6FBeIYRaoQ6wZ0U3aw2bD8JCqUU/zBzX8Z
osNl7Nbge6nAtZdroevhCjh0QkVLTy91bOza32kriRgmAA/WEJAuvcB191iSOYz4
cxPR5QWAZcQBJRxGJU4fX0oJ1yBM2TEf3aOK7gyD3qhBJHb3fats0gO5ovfRuE5t
6PYxHvVYd3zB9lVG20de2PSTU+m9k0iLAZ6nBAfqX6tdvW/a+CZMP43n/gxIo5lq
krOdbf3v+72gVLoAXc6RqyHDENtnnil5JO5iCXzorvaXAHUdiA39BeBEtVgy9nxp
Tloo6mrSVKFKQTkZZOmlOo4TxHUKPieuwelCZ8sSs5Y7LPsMrx7IJV0nWPO19HFS
GytS0VICgsrQfZEVNCfxzfzHgNN7/WIhS5fYWvcRs4kczDULRuWIApGgRA2d/Sut
iyMkfpiYTyEzWeL1C32tbcLZJNEQSTGTuGj6Ckkw4462RU4qf0xVHFuZdNLMWobX
gGDH68Q0RWB4WEaW7whAW6xFlsfy/utvSMfbUouMNIYbQ1KU2jjjA5AaSSA4h55l
jsS5YRqLFIZbdMzOGef30tUIjJGjFTr13ISb/+d4yk5vTwFnEWLI8T86ITpTN0kQ
fhpmEjUzor6pW1KFnwsNWmukR5+g6PofGuzQtUyMgpWEnCtmbAM2GUJW35jeBtEi
QHSSluP80oh4JyaKRtuvTPmSb+lPWggld4uUSncQ2qdg37zTG+0C3U/Yf67zSZMR
S9Cc445Jqp51k9WiKWiLSRbpgpSPXmr68ke/vT9vzW/v2Up3I6t8szPZP9G7g/QH
JchUFEC04piPCreATd4HZHoQKavcpejflfnSr3k2iE/dpb/4bvVnLGIqbYBUFo+i
8G5ZjJxDjoKq/VAfZcGPDqqxsHJbexeQvIoTSSCxd0LqYJRQkRJISq1q98eHGFey
GhfLFUJhnjXMNiLD5SQD69hCw+I0Tm04peVFCwQiIbcUA1GdcpeEOPKy7lsU2tbB
l1OcAgatjuSSMWubfEKfCiE6ctuPhZ/UbZrxMLp+/YR6VGpkxPKSB5G9QJ71qXFc
3zQ0BB1KG/BOCiNso+VHQVCbFifWKn/Em0i+tYyx0lnqPGI8Dts+tmTMmCfNDcR5
tLMOsTCW09FJFQGtietXWKNJNf+Fh4i1raHYG5WE5xiJMofy7K4TZYp2j3ZWbayE
0r2wAS1+KgoTQVM7454kwdK3gYNANfreENqr3NTD0HgiqnZWNMpzEwUSeXhr7lqX
h9KVO1ri9KY54TIZls3xWQ3DFI5d9OYmxmjWEkuWN2AVbQoYO2GkGKnC2z2UraWI
tmmgdJQl8Pc29Exst/mrE0CEfCNFQTjcDhoiZJquYIqSsquPeMoWtDB83d9skjju
7dqgBxfeM6/h1PESjMTWSB4mH/OmYLJL0G4VmA4LRYctP8HMQ/C2kiV2SylFg2x0
MBIoEuhu/3F6NT9QOYI47bO5BzTSlFS30hOkPeBOpPsKklaBlkp6Lq1tiu20aSV6
ZuFx9OpMbL1LenUFTW/Iuu4RJ6OUdl18N1kp5ZfxmXZQW2pYSEkHfGM1L2WE4OU8
h0JRaQVAgFm7AbmZy5G10bubI7+s0c3xfjBUiKHLjcQJQqHdZiQEH41E+kVTHCZs
q9zMkYsAdz/xiFuh2HQoy6NARUtjzoASlxkeI+tTLaHSKbTyHYlit3KbFi6+JXZL
72LNhITd37tdbaZglBK+3ROTU/Rm8GqWvIWCPoar/IDEyvY6XcHD8fOn37sl7l7p
6kToV4Pw+Dx1R80TrRoUVjuJSh77+LYyh603GaxDRIE1wZG4SUoeVoDylujA+KSu
PYoxkZOlfqWPei9jyEGmEIAIOOMJVLLBR633x4fVN6+DS5UcXyzHDqdstHsyjjdP
3wf0Sk4Pzp0j3/kbWTSW991/d1Ffdbvw+Hwx1TCEmnDsKh8bwhd1M68KQNIwbieQ
jercz7i+FNUVLA35TIb82d8IFBamuLJylMcVnvsZ/3CIU+4vhLYkFBwfTzjsWE0g
IsHMh02jDcbCV0hbISxSZs7Aq+3l8zY9D8tAyDUZ9uoeF0b9fZPTTkiJfRwwKNfK
IMWQny4XvSRkbO+gdpbLpx2jahCkN+7QTxUlCS0ShTdAUnQ30ur41D3liMByyY91
wjCT9JqmmVbtjNdJxh6xAIe5ln909dj0mHXIrs5J6Xnxt/5jh6bJGuIvWYiyVRdE
3zgb4MleblltAsMTOWUzsoU8W7wIv6pGcd5lhGzEunNE7pC8JiRZTH4+3sX4vons
pFHvt5eFY8mZYQaK0MDMnmeEO4az02WTycUv3VZdR3z1H/wJtSzUrvJhhm77Zr2o
G94x/ve/Eg1RnY50rxsgTauGbM3oVRiJN5bffP3OK/sxpHqxWeUlbcNIcJHCvgMJ
CeX/fX/ksnNVBmQNxAdxIxwn8+B3wPsZNR4GKbZ6fzoxlq682BuQV9Hs3gTH7QI2
bR699Jsf4lgB+iaowRDcEFzJr2BQfS8ZbCOd7CKlWiCjSMj7wdInl0m3Hfkz/jhE
p4WW/HCMKtCn4d2t2vKGW1esu+sjVbfO6SXizSqU3K+PSOamOwEe0X9Qv5pi16sS
MmWpfd3AhmHl4XTKn+nleLJQlg5Nmv7cQZewmSBN+CMjjxd/+4imw86DPX8LnpWi
cWqadaYMypvr9J6+D54WdkElWxx3FBzJvmKzYq7cxs1RTZOuFHj1w4ioUqYymXlp
yF1Xy55i4FLrrmWKQioN9ZLrpOopLlMEE+btnbThzu8M678ivdoggS3WpowcA2Q6
CWZQdn5eRkRPYKZd/xQsM3rWO/TsGD+M2aaKituhEf3qqBtAt+Q10g1Shm2u0Jn7
uiii3+NRzhnV0VoLMeI684w7/JDbDf+tkvYmCh5oFLkUvXCGD/px+1vZuaFagi7N
+pjqr4qewQWAmV1eI5eeyABzm/GpkT9sTRA61kmb9XTXxZnBRhOecaVhCgq87/b+
lbB2CEJAWGw8v3kY/reJ5mFa/uGvEMp7XYRlH2p+wUkBcKoUT2MLXZEufgQZTXyY
SMfr5FhslPz2B+nsNA1+HqTi0PDgGbtazIxmiO/zHbTfUvKYtRW3/bSKipfwe3wz
s4MxaMYXNs/pLdGx62VmcZ268WH20JN6wkAGQbpNDDyRKZLWq8k5GpPQmvqG9FvG
epvMBiUeDHeXGJP2Kgv4pLDvbdxr9E2Vs31aKzTFDvlcG7hXYgVbxeLMck5M4GyN
mE41/3hqxfpfYYctRUmXneIK4GZ+hhVcjH6I4YVuX5zOapRtVDeZnPWuThHnC6cN
1wSxEUNZmjufTFZYuVJJDE1wKEBJQaPLTtq3NmrKti1VUjYAOMHVki3kMaFfCjo7
4m7JClSWnBbvZC8HA5Y9hrH5ElVz1pJkjxyuHLoOVjt8B6wEU5ZTMgliPLN+oyAK
ULZQeXMgI2DEC5tsA/EFvW+xsqoV7DjBOCRuWko+G4K0rVgX5GgKe+gdSN5+M37m
AKpMuVBTvgdR0+xSKG2hn8kz4Zyuo+mngJKOyucPWOEVMK9OF38VXHlh8/Z+WFNb
WKnCS2lS6Pn48gLLsFGmygcyCQ2ri7WaLqxo+gQ+Cwi8xqulGbzXvclWXpdgy3eX
jhCFikr0e9yzB8zYnACZISNa1A1Zc/UIkZSS7SKKY0eVZuycsK5avzJkyxZ4/TvN
/ObPYSc64iwI32smcfVpHjMODGCa/l1QgRznSJjU2opUry+IR7NXYMyhh5J/edzL
eMVXnoXyCqgBi9mZ7luBduPgrYIseHkYwi1eEQcaPH7q8fMxGjB9DhgT7/H8ko1j
S+U5CKnGDGlzTO3wzrwJvl0qSwv3pxZ+KRhXGj+hdWgggf3d2aG9FIRZpI8boP39
6GvaWb3d5itevkhpdL/sMbGW6Njg2gAGrbR9ez3lsAziypzZFXl51rNzUbBSnX9G
dFj+qSmHgqd3YIqBR8ylLolf1W18fJdkWGeNcxOfe3bGmOYqZsQrC5YcVtDXCm5a
/0TanVwM4LhwzJSEONcpTJKIqPOoge74Ya8cRUcS9ZOGpg/ekZKWw4FAwcpHTdWF
vv+BFZ5IWgHEYLhKqnJdwMMEKh5j3RLaHFFKivx24cEYRXQD+eCBO4V9utYmUOpk
r9p3jE2ru4wRupyw//m+MvLlqvUvNTu26hjpp8IUGJ/x85V8GFeK7GDHGlY5IUft
f2Wi7BnKUjOQ6fhH5Kq9yvmApZHDeJCEVK+U2xPBiwQ2rhoR003G2gCIczrh8IFS
XY6u/9LtbCgmP6a5Ra1HzKzhCVhSGjJ5EYEEP4siBm39zxf1dWIuLLPzf+DYmKyC
SZzL9WkFRhISW/+C9kNj3tHEK9c1ICWlPhsa8ffDDL3j4kda4wzoJ9YPUkOvyrVm
WfmP3ybc7apxUeN19L3rKrystCEt26kHWIkS8cZGm0EpmGGUtBrff5tW4DRqJodL
5kuKZw3LXWvgIGUIN8wYCyiWlUke2tT98/rykP1rDUfCZL5JnHVVvcv98h8IpiGz
6rFKk+LqIlqYkphZcnYISgon7eUgErLvUF10CXXc1glWLxPJ/SL4O+AjLRFqDIc5
akWiuGPLWz/IxnJr+I68O8Xi50JYGcDlfKnowjj7xuuZgY1usDriXBSrEY4bDv1U
xfzjVbwoGruZiBZEX7sUYfcjwJ7hYQK83eOhp7VjQxO+CIHEXNrsw+VznWt0HpB0
EyNbW5G1zGyiNjIVQs8mnxwd3Hd/DViso2Xeu+MLu0fJqvY30UmoY6hEfV8N2XIq
Zjdhp//eMDV+q/7uPu/mp8p8/zf46EapEiw7PLEASHYMlcrVpCgwE4pH8xe/bKQl
pjmJKTb444+kgxICZ7fspviguA/7cyRjvWIYQVpB2aUOGWEPDQ2izVwlqtxlRACp
Vl4KNtxFB+2UanDm01nHF74gfILFQHtYRR0PZnWfEoLd2opfpFV91Q4rFuF0UKvO
WhUJTpihQJE4M1miVYgZhNVJ1GFDJjx8TNCBc2q3YS5HLzKpMo6m7t8nINTVhq6j
5zU8d8jWRxvKhCY16iJJ+95NV39lUFfA/tlZnRphbGypcFOFOADIZaGCaY7vruZJ
I3C6Xdfr5AcBxxtrl5suiSgJiyrZ6QNextGSd4zS7yZQbvbuWGkioPEzbEZTia3+
snvpx2/TLfwyC0Bk+cYp9S4+mBQxi0OVDWihe9qCfxHQ+zP6oxVndi8RGU4LcZon
zi6GWpj4Tez8wDNzr6m4ctJncXxuwQc07eci1b4OwSlwILjUlWAlwNUykLwdYXcV
59CoZ9Qnr5trr8/5LbKsrmO4OLvjf+QgBGfbo2pGi10k5X/zQJoF3nAwVdyebq+M
dWaHigmGU8GUVEu+hPfI+ujVRP3DV1PL3pokE+Fl4ozzyF6q082WkARJwQzlzuSm
9pomSnCTAnV9vCTrZ+eqZarJ6s8nhR7f7WBbxgA5w7qMC2SR/l2ULO78J5kQXz3C
rxnN2oBQHKmGmOUyJ1FgQKZrAOD5ETe3AEPBWr4Mk4+WEbwUxbTLCwmgeSMEX3s3
xihLzi/1EqAlEZvBdcODHAFoIETbdOw5IIlEuidlf3QPqTA1mOoOfbaycPQLFKk7
hiVulMR2vv4/zhLXeXvdxMA8jik5fhvlzbDrs7dOBfnfIFyjjJEk9MJSX0Ps9Ot0
PsR21DI8+UwX8fC/EQNGZPVvGvZvAimr5TDffd/7qQqJQirUAtrL+lAqxHiPm/LN
pCx/U/If2VFgiyFhoWmVlF92X/WSamjABtiZeo+etX1EOS9mpssddstjbwBkAeGC
kZeiu2GjgjDDlKE9avljtTVgdYEqax8YlVjsmHyArdkPAEZ+IyEnlJstqj0uO8yP
PgBR8ptdvv6POCqJccYOxFNuH/TgQoN4Nu9uqDrsUvdlWDidI23Pn47DFb+L2V9O
mGAwa5fdke8gj+4EWlLxQcKZcZtltz6A768gJzKPDBlGiwC273qYMUySHcOg0cbR
1wh4X2jOUQoHPwLRRQSArRegeYYOo/NSpV1ugfkjNaLQz7xyn78OpwaBexzN5EZD
V7SnDIkr28LON2KuVoJ5NxxA13/4aDF9iZ7UXpIXwna+439hP0TPe7t8k9IA9T7F
yEYVPrV+kRuXlYynAZOwLjtcOl6QHN3xgKzoOpYqMxfddwte/MaSZ7daMUkemIQ6
0hvWnJu3rPBwT2otBq1iLkD9JloGiac7LeEGI6hdU3f1knUp/NI7RSNcIG8bPfCM
ngPzhe9MRwP+JZuUJAfgEiT56Ai1QcbpWsQioYIWnKFtu+1YegxK35uuk6ZOoZBP
qz4GkWmT/YKjpXVgkzuosFjPeYOFu1vni4Pgwj9Fk1yDFESAnSBRTxuLqDPXbZbo
5u+L0hH0hvmWrdPWRC6+wUYjwB2LxczNvGOGtWZC9wvb0kq5bxE21QivQcK6SzDh
FfWicUG6k4NfgKnT0d7+Y8pDa9IQusrApd9bSYmKDBiJy26ux+yYilEaQyJZt6E6
puJt028gV9DqUr1olBsIMp/ScRxwY3jIYRB9X7IE4+QcYOobesXy8/hCAeS0TqvV
gDJ1Rr+7DAiLQuZdCaCuzQtkqu3Ye648rKtygyrcPAvQnecRypxVjr6gs/AwaYM+
7eGt2Ky7ldBZtLjioRr0J4x063B86d9BNB5vA5tE3xqPtpKCXw69msNbpco8TSVl
IVUL8+QsCBEM/i5e+9eX0a0mlAM22bH8BhYiySLXMNl2G8DZwpXzqfxvBITjKFXV
B9gE+jsdaQYipsPU2T2uNzSz8/uaYV1RGkZo/8VLh1zvkmi21TqVv7hvOzpF5bgO
ARGPD0mG/RLq6S5CXlwoupcuRdUk6A9nkk61v7BxoY1XsefeyRA5F5CKadCAjRPZ
yp0QE3OH3sxTrIE/PYUo3UOtzCLK3WVZzboS/F1TJvQ6PnCvZHyE7wgalcV1Fbtl
6sd094vrcpSHOjzQkx+eNjUJN+kCbKocD2pISGEtjj0FLqRx1xy+CD4uG0k/oAeH
2qTBuQtzN9OoOZNnLYE/GWbi1JWEMhDaYQJu+ssUeBBIicn6qJQZ234JPHrSrDaM
kIRBwHJNqkvtiDxUB2kGODrlU3/PDA+rYjpiDX7LgxFouyjZ62yrn+g3DQPf8lju
bNhAay+lBvcf9qrslLcqdhztk38bbAKD9VNHfzs/NmCNDyb1sZvgWo2qsQg8iUy8
K1+Jpzvmbxlmc4ECgYGe+rBuC3yh2WtukC4j428mo1drUoYmr9LUXl/slWXSMdRN
9JDXOLkHd5tVgykmCeS7f4O7YUohmN5SHWjpKZoGl52RHtRoUe/FzLezf1toGc5s
gNuzOax0KqtEFqZ/pL/rc+t3WnUPbjtlFCDNA+WnLIcOC9bCZGh1dre3aFb3Rhpg
/9cu2ypuE6sBD4evMAFs5QPHL9d/qoYww4ZLQ/IRuI/BCg4sRZ9qAcrTTMEw9VUH
y1YbVHaTm1fx55ekC8WozmgDYLiLd6a5aYQKO70K96B5cAwiQgXf/OagBh8Hhhma
uZzH4OF8BFy9JRET2Q8xhIlFdT62SHKdLyVA9Pita+2Ee2w4K0MRSdXuPoStv8/I
dsB/FJ7RZP+dd19BD9zh4DbS46WO2NrJjzzSyQHBIq3sDG2Ql1ywkvX4sJEz/Txe
LcDsqsJVF69a4M52IvC0pwhNGyAWpyx6sxKjFsxBTCl0AW+En885NStWmYwAv2LK
zu35pJ4RFlBPuj57nmpU1l/GndqId/3BnxijcchqpglRuIz4Z2wkob+dK+d7fb4n
kSl2lRp8MM0g8TE2hG/WggMowyvZ5NmcYdbwirK4/cHnin+GC6sjjdvJSZGfL1j1
OLVBHqUOPgFv6sx9CvvrosOet5wyeFsa9xzjrwqQOb4AQI6g83T1cl5Og/TPP/SU
8DzxYThMtuVMATG5Gb5PgcxWddIilt/ddmVZJE3EnG2YugQlEr1yCa39UZ36hr0P
pdaqE7nJ7rS2XR95vho4IujGwI+vffZqATsDPb37ANLDZDZbTAABbUTQYAPU0x4t
wl9kXWGZNYaKIOJD2DloJbs4dogiwUoqnEMH//12tCW71q/MjBtMlKCHLTuAz0BU
eyp9wOCvAzJerfu9gmianyzXG1O1E8wPH3oWVh5Nhi9zXrM2kHXhBmcofVVUvgwk
0htvC1rg5noYjI2BSPpfBMbdaZG15e2qdg2tW/Fm6npuHywvUEqgnv1c0kgYwgkO
lz0ePf9sEa0+RhbmAN6XarOlV5fkSwQaOTVa0vjlSzenjeLcyRI7rmvSothYU+OS
4yLpKUNaU6SnAzmfFpAlPxxT1kLZiCuPSGITmmEcueW8IfI35X2PaM7LotXNpkwL
t3PmfoG7KCxo7/DgHBhqyITlVIrheG5AQTB7ORrDloOPYl/PN4Ss4591/jkZsnKD
ISkDS82PYm2UaQBxljAAljIgzZdXy9zHphF5ya/bLInLzP4lJuTQrVH/ndvpabIN
5hGp5sFAgXKohl8usWyTICCEYs5ZDCUlQO3H/porOuJ77bENXDNdHbEO/bGY8HfV
Gy3aA8hnA2P9Id9L8gcqBrNkoi0Vp4uXAEFNAzb+8mEMQULXFRs6IfJ6VkEJKrSl
UlD7oGYr7+oRuAknkYD7EWz9TdytbIqj34z3UtZ7MZTYVGJWep7ApVlhG7fhfUev
ZHE/Ic9tIIoYYK5JuNUJnN2ZewyIeAeRq9dz0/daVMqVAFhmkiOdXu4uKoeRCPW9
vxQkpL9yH1HmUUV++4SL1NM9zsPzC7w/DdAstejc8kyPofRy1gjvpqOPGQR42Lp/
/HXN8788hdxWFyVOMv944lAJHwq7wVo9WlpvGRVLFR9xZvP3rtLLm5xbjuShjNMI
h4ANtdDPrWOphk9bHKEsd0ta2BCiqoxw9nK55Y/Rbl5iGNI78MDJhIG3k7Dg9gTk
HczBfxYzArfs3JpC/e/RSSdUDaVGGXn+wAis0VpSD2y79gyfoFj4G7l0CubwMvBp
+8Au34f5F1C8jGsjbN384I4+MYwBi5Mt6u88gL5BNjGARKm6pKzFieskIb6n4Uq0
pyxNI5WtyS3PIiQZwKwl8xbnOaffC+d3++73FmZtCBdHWTALPhAbUof+rXDF3GhE
I2MGsThOure2N3/UftfPsjgfgI2+3+9i/GBgK4Yiv9gk7AkaIFUCuIOxvj64wvTv
x/I9sw0veJ24ZG5ATL8BiuUmb3rGAukcxhdFuM5pxqKxAnj8LWow5UuSVYAPiWlH
LN12EXA5ks4B/DREqNENsnvYfudIdgzngqicLuXZTjXJjBH744J/miA372/7r4nl
/GwCOtlXrwMHpTlzDzdmW2JWd7ISaoC6dvzcLHEXmip1mHHEzgurp/bEnuDkZA+D
xmq2zLKCYTNLmPg1FyWjPg2vJmw5G0dyxlNcRhvHANRHbXnUPj5dNpgOOOEwPF/H
ctU2/swhSS7inU3QsHfKDHehjWybr0M530e5FKwT3q/5h1xE/skAHuPLfkoHmyQx
9b37LaMWkj6K/J9BUg1IotPUtVfjYPOVXXjjVhvHik8=
//pragma protect end_data_block
//pragma protect digest_block
fhT43nbC8hpLpnSv0h0qyXIfAoA=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yQIUP2lw7ommBBbZEFluZ7QKjCwd/j7vbwP3xla5Z+EIIwjaEUSwSHQVi+FtqL3L
1OpyOcz6JnR6EFqXXFHt8CpiSCWKOs3ws+X6zyxu8UGfMor1OylU3WU/i2RsRUmW
Oa/w/p9b2N26vkH+1Od47PRHg+0jCmMlwDryxIn99bZcBXgOv9/pMw==
//pragma protect end_key_block
//pragma protect digest_block
bTqZix9X+VZwWP13rGYh9A/zFNc=
//pragma protect end_digest_block
//pragma protect data_block
C5fTKRytUp6ALs8YmKwopp2t2wJ3FVRdUSV1wuvaABs/QQKTvtwpQO9ywQ8sGNh3
wr8aq/c2RsbpnQrSiBUCD/G19FOLBivm8O0EE0v/+9X2nmMIsx+iFdt4kLpBJ4Ti
inb26Lsp9T34E2cJSmBdEGBiWMyDpZOnhcgfJPZxF3uPoIwzuIVaKcFtkIFNlpUw
p02Pe6sL4xFqSw1s5FcCYU9e6Q0vNPeJJno97rlK/ucQZOk38KatNJjaOubn2J1u
Ub/Qa3xU3GWY3zNLwcORHBm6uneXv1day8KXrDYjjdw94/mjHlNm9/LQdxVnO4pP
IHQJm1bUr5vzt/98/a2E83uchUM59V5QPtv9Y480b1rf5qMmoubIgwCBy8/iuJGd
p2dEOtjnC/PONs+jFuhTDPgXzsfTPTst4dg93ft2r2ugWKc8fxITIxKfwb7jlE1v
sDW8G/MEzMGMTMpfEmk/9jI+0AP7qjvvkZXG0QX2JtB9063/VIfEk93GrTVjvUy5
oipHozP2vzgpYnviIljxgTMounrN05JMM9PdRSIkQ50BjscqcFToT1olujz5eeFN
u6KnYAHQBvlJwpdSCSMF9g==
//pragma protect end_data_block
//pragma protect digest_block
sWHNO7Hu8GqQXTRJiYy6rqwgWNw=
//pragma protect end_digest_block
//pragma protect end_protected
             //vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LEg7IInfOswN9JdaevXBTkYdpZE4ET07mWqKe2CAhJZ70r2XN8lCxFqfL7gKEybW
RDXJxjTDW48JXSnTUOZdjlOiiRzu7sSrkxcdh+7A/1GSONVWxd5tpXEh9lT7mW8u
IDL63wtbb1Jrr32TR3t5Coh5TwmVCZuJHy3sSDizh8TI5sm/E4xdWg==
//pragma protect end_key_block
//pragma protect digest_block
8vH+5z9Emzs02rtPHAQQtrjGMgc=
//pragma protect end_digest_block
//pragma protect data_block
AHK8VBWBJBwX4ErGz4ZajHBkqwYTKzwJdroYrjXSqe6JDW8dgBKiM9tAg7QUiJxU
g4s1LWEndcMk49WvY6etkrhPSVIXSoUs97J0L5ANy5ykKWWIlthTlkoBFgrpRiyW
5CCaoYNPF268ePkLHRK9QlQ3CwnoxGC4WNvxUHC4zXXrZq3dG3swwfaK8k/IHXcA
CwDLjyS2YjA1y75tiVnzAzSk/l+JjkD+u+mnIMSUZ75OwCqjn4IghHeYyPgGJnRw
I9bP14frs2G2+9Zhfq0G/leGXPLBEJNRuD52FlIo4sQyyCmWPzNCRo80glJMhR12
yVWlJDW3E64y6AoiQFGvAxqQ5LuaBUk3zJqjRW3OFIIHCIrbH2grX4xCeogXLc8e
NzDLTP9Kt2YjW4T93avvEY1cLagU6CyTcEkBei2jEZoThMWbuaWEOXQcdBQ3T5US
VNKXuMV7hPzauRXYNEB2sNVH3djouyo0ycMLHQd7PBML+4LsJEoO5GPkExn3L/oG
6CCXnJArrwI5ZLY2K1nuIoOSki6A03CjtG6f1e6ZtvbX8tbyw/1knRps3ZNx03YI
D6h8YEQLZeny35xCdatoPxndzX4GiL8AZJ10KKnfJVQrvzeYk+hSs7vaFVtcw7IX
pAehN5m69Nx3QyOBjt0KlUCSZ4e94mNS/Vk/DzGkZDYd9wbq1S+X7M/+nBZmzH8l
RksY3Uq3Mz1kNu+8PN+rs7KF0X6eK1/Z8V1ESpBuNyel9ZNF7KoVvyTIXwUXK2bg
wocpCQJN5IdmWR/05T8/uDjuNlGSycGm6UjnqfKP+SWgTnfaLYeY3WTLKxVEAHEA
8/srCDbpwm+emR3qLsvj8tIC1weqCSpaW9BDarvGlECjBHTR3x93plgGiE8iZtxw
dY/QjOC76tiXtni3irCnljrMpHobOTlDdarczfmQQPCldKbTJ7IBcnGgKmsfOsgn
8EPo7E8+m/abqQuaZ1PhTL1ADJzdzBXJYuh3WK11qfnGRm/fKBXr0yLrV4y7IQ3s
IlEK8hfQPvouqbXHRfFIUlRfdgfolVXeLbhnKI2PQ16iX5wOPWXIqaXVWp4gtARG
IhSAQQlWWdrXU4NywC2A2m2ZwyUSIKGy3L6EPsktqOAw9Im6sX40Fbk3iMv3WSEs
3KtfA5RztzQ4Ut3JSwMjlzIB9iH2Bq4d9Yos2tYU4WeDKit7ofqU6b9AXL9JF6CA
PASMWIFdhkzIQa7d6chO1facPMrp9pQ2LhUnpE+TVf86EQwItotEpkxyoPM7zlCp
u6Yu0N2E9xcw06GOLII4ZHJm2TB1XzZD5pwbj5X3+3XT5snwOOvpWW845Blwwe6/
zlbDJUzF8kMuWfFogO7XXD56R3Hb8Z1aL+l3yACmgkX7oZBO6PAxalfF8HBlEb/q
IF8E9e0DdoixUZAiZOHFVBHbZjP2qGaRNYNjtECLRZGsAJP/rSpPGVCj/0QsG+x8
oxRQucVBsvI57QqGlrUHWB296p3kgdzD5pTQUwIDaxZU+zQuepWQDzalag1FA4TO
NMfBWO0q8iYkWeKgr6hhaaS1YMx4yMekC9PbV6NbVVZf+igGFVbkbAzs2QHlxgeu
iJBP177FfeD8hSvcQMirx/Dbmz0xYP1tUYsnhFAbyg+nHHd8Ck+onreRwCxNSuCj
CF2L3JlHhQgiVLm4Bj4Sd2f4QY0eLWYii4NgA5VWYl977pVmySQNVjdbkH0fytRe
nMDCAXZ89ENnd5kbZ/7dZKtrhxdc7Kxrxcf4Igv0PJXSciWouX1WKFiTFrGq5tNB
RmOEGF9Da/nip17KZB/i5K1JisysSqY1ZOWQPaD8g//En/eohBXZOIpISiKk+yXT
fKmEwfqO0DHl/QM8/bPA+rxGVjwOpQHTLMByWUDmz1sRF0GMJln8uaBgWXpH1+Jc
KSL2J95f2SOJrvX8oTIjYjYh+/HpHyeB3jI5GUs9NCyCdw44QS2x2tQvppDhAOnZ
6fE9i6KhHiHlpZ4a2SvonVqUF35yiypDTB05+zYXdnASI5DkqvRssPVsud+JwJLm
v4Mja0dpvw4mDxt/Lb4ZkFTNtU7z/K/ee+O2FLGjz41GHRyO88x+maq9M/Y00Vxy
NhZsKICZfaSnxN+2ISYdijUOAEPztB1A0RDXdlYye5I8Zivlk6y5bCoYHVnbzl0S
Ufkb0mEmNxMriN1RMfvJ1EKUmiPYKGafKD9HFu0yhBnHfjJ/yvytBYqouGVkmp4s
6Ax2IlIHTXrdLqyFM8UnptMMaoa7kwDF+pf9xs1M+fef/FbdlzDn6P6GKCYqj3VX
xpU4YNxFD/e3iUIMwJCaGcbc5XB7DEMySnaQo1GJlSk5W3QnWnbbupNFT32U4ekm
qcbYhMWv4nWe4Q+d9NHfbZ4vI4KzWj/KJTkZKn4Bm96JrMHZhm0utvEJ+J6IrLEK
YfY03wvcjbQtz83g5M9nKMbyaSB2uSnKV9trbYRcPDrNDhJn4Iz2NSntI4imo2QQ
ewpa6Xo6EnijiEIJHDyDzLUo2dLFUtNtrOE/eZdbYthDMUaJuz8EEAD6+ZQghatp
sx3ga3XhmvbhIHaI6dlKd6HauaksRpVI+PCzHrIWCxt/mcesv+Fci56E1O76gP5S
YJV88X/yfS8hHynkzg6AJ1BpX726LDob5kJ6wOqpqTQ29QuYLdjN53ZEYqMrLVQ4
gT9b1AUy9k0lR7cRyHXHzGRlogGJAjzp5oKLJQtv8Q5EGiVJQoTjk4lYc/5lZbt/
dC0TWgTZ28+kCg08qNpVhBRphcfAiT5egJe/ot09BXVpkofZwVNI5CEkMONTF5+f
P3suZA6/xNvQNj28XomFwjojc2AMe7/KUY/Q2xogodYvFmNOf+dsXFYpPVoWYk0v
K/Qc4jl9aAI9Q2dVLRfzlmDKyAxmQC7csDDKlUmxyskaTwQ6TZOL1MO6qjAZ/RjK
ZJp4lBxEPjolMVpVIUtyicoD8n8JBE6hzScatXCCRuPeHv+k7ifcIgmKdk9xpW0d
5K9xS6mYu3cCmTAG07q3T7oc9P5lEy61FrHuOfBhAqhQf9BSmRmfpmcQAt9WC1D8
6RzL+yNnoi+BOU+VuI023Ew+zQmgOD5PmWNJgB+ZXTk0j9omXUI9pSpeaLbfs+vd
Wo9EKbFU9HzCZU3eQQ0vRO8LI7qlgje4JxEr1y5UiTBokDUcbTMHueVQED4QsphR
X9+yQrKGi1z8vu5IxOafkMsTyQT8z+d1+ITDmYPmOJRSu2RC0kxJOgIwC2Rs1RJm
zMR5WnLyZQWRD9t62TDzyo7X6h3E5XATPDL/5yzRzQEXW8FodTW4bm8T+P47pXh3
jV6/MIAN4wnej87ncJm2gLkyMWA6MEVm1T4Gg3kufKFWxhvl4IGgovzLqWZaPVHL
yJHgND7Fsq1nOZDN6ZC7ViWY971/DgGYBEPbPu4r0mEvbkrXvh6Wo3U9vJ84Pwcr
PJsKF9qK2IRxKnlya/S0uWmVwduUl0uryTl2uvR+lbr44vM/k+uqP4fbvDotX//Z
MjNAF9VIITTu9QuzQ6iTZrApZ8d70T8l4jRfQxP3eDevY+7xgGgfHLjg83rmk1Z/
r8d1C+wLeOP0DwQyH6lGMbGKc6YFQM6Rm+dKZCOYQc1zxUZqG4Lv+WEl7/w4EGaq
v2YdWS9eYPpCNR6DOCBjuppJWM0v8fsDGUBuEa5pb64ODdvzFX7ccoqDag9zyd2S
FgTg8XyK4MhQXNF3xnYaHaMRJsv1zdqpGWaQsRfLMiNo2FZzEpZCu2pTrVxdoGKb
W/3PzWFz2WdtuazGyHBuNC8ANGYCrmYo5qYM0FiqahAIDSwxUrHb7lnH/3B8M1m9
+FcN7Nestf89XY6xt6AbwRIjNtYseEHjwc5F8DQPTuxJMpZehH265mHYJVQbAABX
l4Zs69C/MHhgYJo15uS6QhJMs/ITtwyUXF5V2AeCeA7n35G051/IssLfcklD8pUs
Wku2TiR9foHD6Bl84Lsk4Ga4bw6zpzyY+MT3icKK+CSS7YnOgw+BKjiZ3vr8f9/M
P2Umw46OveeLF/GjOgwyiU9pbtzejzQGYb2mgxOhB9wOcPokrWNR1cGii2fits6n
8bJ+W03uyDkx65NQ0FDbUfuyoGdVkNDWe7Tv3zgjzXWSOMsHeGWiVBIaoWYwqm8/
c837mrRe1hhKPqdSXwsAccAxvzNcL7WzxuiidqIIRHMHDGJd9I4kDlXBVd40KvYs
Wyxjj0R1PvrwHf3llvKTKAy8OBPlyEGzdmaIVMUjfICV8R1cbQs/GBbtT2pU51Rf
xAW6oj6GBKqTFMwWIAa0ewUze9nEWppCBXi9tUQG433ysI+PL3EqoAtAPEKHNkp8
Mj76Mmiod+VdFjSGikiTx3226cR34mBPIetaZv6qgBhKvTrchPfd7D9GS/82KR0h
UgwIcNu8oMCvbUzuN5TghdlMrQcLFTdhDzvRbhPu4SgyMRrlPq53KavyOWzJaP1U
FC7wfPJK1B6Mk6mHNR1oZGDS2EaRNu9M4X3GaHffX9nwgxLrW/tgHrpaQWWgWx4i
cl1S7GqUZqLZqP3OoyLz7Q12e3A/gY+xQm7IZkowd3i/a5MRmLMKyjaUsLgpeBIM
qk1yU0eLmof59qyezoNDEPDVACSDgIY4kGYphp2kOy95WAnRdtXrU/O2iUWGRPL2
uNM4+a+88qe+UfWKjDFh+sgoL2Oh8LsCDcRaQpOmdRIm9147Ez+q/Yb+kDdXQQGi
aF88VsKcQZFG+WKrBjM2fCQfxLwZYPIJlszo9q6Xd/MKFJpxo7WVDIPzY1wBIG+e
qHADr46ryeaXsV750K46G/hlA/aE53xf8XcPCLQFtZAHVWp7sP6rianbQTbaEXPi
nDnzqlJSj3nPK+WRnYopx5M2ojGEvXamvuNJKCcQccUiHyAHS1BC9zvP1ZUdKHCA
b+6IbMumRx4efcPNWtGyrJyk9CNtpcm9N4MQJfuO4kWGwNua/J5ZAC3nnIwcFl7e
qgCKWMBp/rZIwyYQK9vPbLNQ1mOxM1ovYmTt1Bx6yL7SyxwRr/U4gnBNAExFnbz2
JKnO8EstgBIvTxhdbRuLwouIwRU2vA4VVjQOgLi2YfUPb3bnNODi/sEw/W9y4UZq
CvxH1tszWgtFrsEjf1FyHM38s3VkXWfDmWdGVMMpaKuK5QRLmCa/MK2lqJJjbAer
r6Lanf/Bn6ABgunZ2loaM7xhDLUjaLojTyelX0HSUzoe0upRvIY0Bl3H4MSOk+St
3fgqDtG6bqd/f/IToETBh/T0P6+3nbCLujvwZT3hYgB+hfMGq2qdgtNHXhqSRw6r
3/Xsr5t/z0EgXt0Zv82YGUXsiKopfoNFpcfhRIxpvI0WR2LVGFycxYId7OsdvAld
NmuRTvcEkYH62JP84dmaLMwNaz4xpgrpx3hBbmE0hWm0HQSqYI0f9Pgn59zibAkb
o+l4hgiAChWJ7HNLTiqHUEF5WJhlUFojGCCvRnCOsCzVRe0HKLjVQycQPynJptkD
JMd4VFmsy4eXiQmT6BzUrXW+jwxLABAJbMWmj/5eXUmbIIhVsEbE5wap7tA5GNPo
ZYwy9FJ0lmnQ8g8oTiyKjKcnBwVDEQfaSFKPJZUmiIlKQ/ICfUYK2Cv/8W7aVND0
RAaIszYvCBMNsOwtCXChHmOjIk+3WpJN6khlKtsMIPxIJzgnM+MEhE86Rr8w7lqP
BsA3M59KD2QIkPzdIF+VxDbiKIVUqudHjimxiVY2EjrxPJ6uUJwDwSqdSEowhJZ/
400TdyftWwa8ESlK/tDZEr35p1CGnA1msTYAxzO+Tw2E8X08JUgVw2Xilfal6Aaa
k2xVVSUed1klFxN12td2yOmLYL7djn+eshBYkC/0y+f0aN0roX8NLzJDO/aDjaNp
gS3VARRDo6nrx7U3mKlBprNdUwEuXSM8WO2t85ZrpKHrlY7bNH93xrHyW8MSWEO4
v1SLox6Gg4XMKPXBbXi5buB7iN1P4vK2QiIZKQ9vuKw6vZGtGOhwMqt1Rb+p6W2f
n07AmRzwVHu96ODCKKMQXLY+imDEwBIEgO7SfA+q2cVbpkic/zvMn4XY5S6sAi28
2XsLDeHyskRpSATl2Kn+ZvlmMD0CAvfm1oHomSlTv/eoGWKhsJrmcjKTnff67Om/
61i22xfeD/bc1J4xPw3rkmQJjQYOyOI5YwT9d6x3kIxMR5Qa2qZvAtQThO54/Tb7
TvzBaU3usXLrICRmB2yGxajzyPiW0mb4u6fC89iC9+bBJ1wuzYYQXf0hIreBinHN
q/YC29DwUb9CdTrfbQnQBYieJd40cNZiz2x9FVkrfVFGKB9tMDXV/jXTak3/x50p
xJ2dL7WT/25iAV3GhS05qvbiyyPZut0e7WG6M+7grVnAYAGCmaNsWhoiHymF4drl
w/cKZY52w6/+RdaAj5rEEWgV2Wn0gPPhok2LROMVmA5rSfClsiD9wgQPMC7Eyzy1
Wf0hUbc0lKZznqKrWz2nLIjT0Fvp+qIFBpO1w3NRMo2iwqt/6uDziR/ENV5iiWK3
pXvZ0y2YjQ+JfVVZfHvYanneWtFFNg4l/FCe8mAyS6phJWnjTCPeojnmQrEPQmch
2C6Pb6pQxIoYxsepL9vBrfvqOvbR8pBZlhH80qg3aJ7YuDxMPAyHVgtE2KdZ5TCZ
9LepRaRQHOczdVFl7Oz6Th3uN4TXdg7Y6Bi7Yt3gZ4cRath5uoUdPs4KMxWP4VHx
bjSlhxPI4JVI2PHnmmJtEmyx1y3RxBus9/E70QJfhiL7Rte8HZFdnAVX1vKhLgzL
cDVVziMv5y+7eNq03H9Yv0ULaMUPGMqz6yCC9nNIQoFa+v35qdEmKmY0CeJb4Dxn
tJv2lg001bY5lQ/gltqxHwxAnNwmBMVWpS4IRlMVE0fcZNig4W4lUkkSQ6VJ40hr
QHnLxXhsdgvyfpoZ32VO/zPDl5d0ITKBi7CMwl8Yj+m1BDRzNgchvHZLglyjs1Bo
5kV5qB6niGZWcrMHZFRZu77D7yHlvrv7SaOlV3QRpPOjr0wnQsniC3i96DAJ0Q33
fr7E3er01hDpnYlAoOhgCIi/DJBaNH/YO0105/L1jgy+JTQFcNHXl9eWQPRY4gib
YULt6TpYFcF+yLEWxTzjYoAb89hZIJ1c0ffvwj37IeJGzrOPoeBVPzrviwbV8ViE
MEr0gtTAY3GhGpLqpihzIgN61R714+Go5OzdUhPC6NwSWANTRcgrCfflGFpGldpA
xprr2+m2Bz6nzj5SgnxGt2NWkDXqQY34p/IogJHsiC0jdStarEHttYsJDPBq6gnj
6zXnf0xrDql62NLHicoznQjY272jl9I12Ux1DnkX5cBDXMscZaKsvItNd7/tL8wV
580BoyjidRgBby5y4fvME9LHlAKxtbMKy14Z1pa7Ex6O/BJoaxXIvj4WSv/8RG5+
Ty6u+Xe6n94u0WJAwoj+cZuAe0vYINmqUOTc8FN6CdrqbhyhRr2QUc+ZdVEkJxqO
zOQ0FN7LVHX2WhRMeeCBvKBebpmSAX5NDgukAFk4pRK7e124z2OURoeKhbqwjoda
/8aQX7aXdIiE4qfV7PGg4Rpaoiwgg4UUhxe/cYVX+7ktrTY33QlMfctLogFXd8gt
2P6UPanKCBI4p34a27Sx2bd96gnxpxAUT0XLri5WsG09yBALFpiCI1jgDfroAslS
DUZfb1aVXpd8swYYAY75BwBz4sStOrl+cBIOYWU/MdBroh6aYUwARScjckRcbQ2b
fzL2RcZxpiESEWTVG+GiqxZezSQuymjWz0hP7itYbRuwHFygEGN48eygzXIE/COo
DcdrVkkZ9RR2bHL3tX03bfo7jtdWDG626qIg5lNbaaj2WemJBV9po+zruQ2ygM6Y
kivnycabZJf+jgIBmqbJ3LjyS6nEpNzik4xU+YEsGHpt1DF0Ne3lmwfknEa9g8RX
yM3hkfndckbqCnOJTeujyQlG+Nm2iAQ9+VHgsbFXZHUdQL8iZUxsW4cMsrJl75DZ
q5WNr2wYgSWL34JgS1BWQntmM4NvmV2Bcwb2cst3dNGcpsYN0cJH8QI1CzpUDkZE
ERdxUcUTAv821OJZuAKRmkXmrgZj2n7BlNHMJ4OE4rqKLaVF/CoC0xa/ZIn32FXx
OpnQ4J33Mk/QJrEQfPVw3wZkK2gmE/lzPMoe1Kg8uCWAUaKnvwXXSQuD9J9xC2V2
LpwGr5tS3Lm/nWMDh3OaUzSOYuG/UYKYXZNWk1bL7SYEFXA2ER3QcAoXLCgEBJkG
DvAWniYE2q4NR39/V4zmgt3UGnQBmtXdGn2peSFJv5bexm2VGauLdKLrEtcldW0X
PV/UZTMVZcAEO0ZRVSTmp2B8TEknjGZnLNWsQ/0sZX+PzHzGFPejGCK3CbA+J1G6
trOey3r+mJIAQzkkn/8dRstBpPLDluIpDb0hq1PSaq+RcK71TG3zRHyKJxk4MtKH
bM2mXHvkGR30ysF2qVTUcxuxCMxIWbqmcmr8mvD/Y30/wnmCwBYu0UvHNXY7F0h6
U+ABoI01b4jXT32uyzsW4SG/L/7HhR6hmfJNC4b9PEZPcQptsFbFheLda5rbmWO/
rU1gZcmWV9Vd71yYYPhiiT3AZ1uK2OScxEGhilBAbLpI3CRSh6NURw4toQHs43en
n1lxt3JPHz0JEArekEPVEYoFOdKVbuTvhbHDmUA0+lnMy51jVYoxB4HHBlXRKTof
+gmR0ZCzGpxE+eaXKfX9RWjlEV7RGDTiidjyc5JnrN4CX24tRLoTvBnAaYL/ZY5K
gI2Pu53IAFqsesaqzdroHiXc21MuIgR8Ay8aPDrutLP1M5bdn/IUk3R0M3alEJq1
1NzpkvHxXCAXJIxuqohth+s9jWIaEqltDhCrExtbV0pQ4ihP3I6mb2INw+U6qaiL
R7/1Whmzm40AozyQlLXWSb3G0xe9O8Pw65ecKxXmJGnWQ9sAmxRh7SWcjIxT0gYg
mCPGPuhYIYUYl1QVxCZQ6ZwygT/ocXr9+j5slJpsXAbMhqAjkg31IQPFUJFrJ0R8
oBR5IoyBc7vZ2qYHj49XAesvchllkKD1sZK/y8pLzq/9sdm2ohUq3AAaAywfdccd
rtDrp7U2eCt0Ot5jdRjkeAkNP2cV00eOLkFzyRdEu5/8UHPyYcdeXT6BDINVjp2H
yN5SGOREHRPM0tf/vFyxTTyTy8N8UwdL0YTtFqermCiGrllxbDQa7cxB/FhPgYT9
Y2U2gE4gRi+PsYluiGSOjkVThybQ6ynnB1TaY+2KH3ki8pS+Dg2DLF66FDgm+Ck+
fYvNL4fuymlFhEDUb2b7EJo5Ytwg3GjwCI3St+ufQxHQ4tJnBqYmfrpnbhNuP7b+
FM97WPr0CjnuwjVi8U+PWBgqGNKHpm1vROIc+SVRJTtrV1l94ojUXct2BXlKS6mE
eKrVNjOfsWwDuL3RYnQngR5fZgN9W446LG8/Zuwevhz2c085uVAZouLYRDbaYxy8
Er7ixxNDAE9BVExikwH1AVFEDOrAjmb18jSmePD7ld5w3dnHXa9WrPdqWv9O9ZhA
RxKb1it1GY8z1aotyFxOctQndPGrY6aKW8+YgjxTyhRFd9NoS1QBX/boUZ/+lSkS
8cNDKsfnNKDcNQ+Tx1ZB7Pv6VSN5YNUMCuFlcNgBdsNLjgYymaz8hO0mLsywIvT2
LWniGlmNOwaH4k4eYDOot5xVO/jtPu2m7ooHI6QkWCSPC2jlEkKU3Uy+CijxYNu8
19qzJW2y9KOiXM3fgbxB0VP9lejIxiBGm7mVlaKn7DjLvrnH0+n1FQA8J+iY0OXu
YmQ63YLiDbstj00qPhIthI/bB9R7ROOmEqo7GGO3AFmgtbdcovJ5O6xjVtSwCSn3
yKY87Qf5AJJdzI8kvcp/CsEmZ1yQ+UpkuWeYNt6uNhdXvff5RRW7LvALu5M8xDX8
G5FsSLRbbERIeCdTv+8YBzEzaV2zY14niLZZzr+CpvZqVhiQRmqmd1why3LDYn5T
L4yHbkYlVlsqdD2zIKJlwFfITgnKAlZgoJyLueb8c2C7Cgf3eoe1cbohTZdg9GiY
jgFfySzibbBB6GbcjIq/fueRXG19o4DnkkBQ85apYTb4taS8/yqKMBHj1rZ3SmiY
kHV9mnXWpaV8RvfNDxQOsf8VzasNfY64Lpu5e1pfOQZ7WT/K1rdoXM68T8uoqW+s
gxdtGhcn4oFbtQFQF0o17ut03y6zu84kr+xJitQ3SpTh3WWSgwW2e8U9j+NsVmU8
YhwfJ5PLD7EPJdEQHDNibtmSnGAz55E9HRqxi9GZqeUA583p5d1lrzyI/4ss/sfT
zHN9XOJZ4HN8GquxsQyTv9qkRqAch/ubQfAjnUvOYT0nqIFNl4YZaIHWXZz6aUiW
1Maq//2fY3kTVAOJ/7QMUYw84FUWgHPM9fZC1IhGVY+MvMlE07xOcfO4vOzCrvLG
V+Htf0aXrNMyMkijenK8dNV6W70QvRM+NoJUUr3BBa/kJ9YeAqgFOLWbJoih6Syv
0SmG+YSMJ4/lXjCAZ2c6CijC5pIefMI8QKWImQ+j2VllRAjQ5wANFcsgIJtDEh7a
ZeI0r0TMniMGnl9lIsi1W84BQUpDavAMYfyOlNgBLCJO5EyHSVwnAFXBqHsKMxYD
+WfcgPK8MWI33O0It6eGZSwkZxF8zhf2IuIUB2+TC3WtBxRGhDHeh9bzFJfuEPKF
GAJEa4bIkRPyt8GKkilQaT/2Pi9g0F4ddZiBJ6A380G/pWvkN5MWGxpuZnp485Uy
wQ+x8CPRioRry8ngU4tGajDcDOL+1OEdqrC1FXkhYNXDt9nnuVAILKi/TkYvsSLg
GHeqvdFr/eTRpH7ZeDivGjkGiOvrycgbZzUlvW5RUi38s4CBlk/lxRa4mS9rQEq9
02RFslBjeRgm/XXD1lxixQLV/80uX92f60av8RbCYxH6fXRyQg7WT6xzTwVojx5I
tmintD3Cm0Y0PVU80hdpwBRYPvNFRRgwd8ubZ4K8xDrpQ0/9HP7riYWeaAvhMq8Y
VXC1IpwCmxRttret7teWYsaazuQxm0qbLkdC6TWS1zyvg97mEnAkBwAByg5kHVwg
qB19FA2VEmpMHVQjsxdzWk9tD7VmKBwBNr3g0PJx15NUgdtgodLPtz64XCM6BvtL
a0LD+TWUCMLDBLPU0Qj+kkSJVoZWjr+nOq5SomP7Cs4tfUyBA/yl8ixs5i5rr1OW
2ziFTu0OzI6sCtZvK1mGSM2ETVHnfDFwtziwg3eL8KA+Lpo5Phics9gAge0WBbLF
hzKm8KCZOMI6L9vD2MPiBqjoqJf9/B8jJ7Y+mUpsVDZqMbdvVn/U9OQgx6H5iEtx
fyR0yTZExDpwqpcVjMuKrL8383EXWHaOxvO4NvcYI/6D9cym2YYLl37J2WDosYQ2
fVbPBud07CCI9Mgd5/X1qBNTbxOtj92p/sT4xnbsCuiCm/QSZVNoCuEAKh0u5VyN
yT1dJZ3SFrdBntvT31dFCORWnWVuO6k9hqpz+phzLcXZL2K2hTLJM00QtTMVUy5B
aqaJmpmqJ0ACIsrLBB4ZdL2SpgLWyFvDhoU3IXLz2Fu47ZjxEwmXyku66B29zuOU
asbGPftkXJFuHijQdXoIay/Z8XAbLbTJXxNBwvoyNZBPTc2HC0Pi25Usx+ug70j+
SuqZiAEWNgdoa+dlsS3triGEq1KlQregrN4sabCZqRKZFhzNm0h3mqak0ZraOKpv
NkxfZDxquEJYRoHJsRP8sBbkmJ31R5agenJP2J1G3Ti7NSkyQg+70hAXQog2dZ15
f2IHK9qvx2+E3vTcW3XPDxetGgWlkQJFjIZpJxPQGHKDiBFOz8Y0Hag7RXmBooGF
eV4PGqBndKYl1M5kDmo4FlyZqoGva4y3DTCANH7s5QX2xmm1H//VInxFeP2ThVZe
6j2YR68jQaS0xcVw0a13+HaY6GRrqDxCRehxe3Ztmw/gl4sIb+qpXepbDzQurfK8
4KCxRVWwnNOyV2W6vd/r8IiUM2R947r45atXNFegmEqi0FNpOEWqGQFqMW0+uViy
ZFerWdwdA590smP8tlkAfAbfhMXT+ysxMFHrmk3oxuaw5e/yfDZcnDcGZRGViRL4
JQO86zK+H+zIkc2IPMXmYoYVOEs9HgAwAR2Rzqk1BNLY0St3ZUgj2imUZ7Bhzeoc
13CbinoJW7eWMKOuNehKZv6Hbr5QDnW5t53ad/6ITTJ1JbOpQRVcK2xsQ+Z9a2UE
JCO1tibM8tL9ZHY8DW193EEW/dr7EV5pqlMtnTDA8YdBA/93dmzvqicm2M8FWk01
sBkkd2QuMA2zgKRuxs1ljcKJoUmSwfGzaXVFDPllWQHw71JrO8aK+ZO5QiyZQbbx
zYPHaiPZ0FaGi3959a/IThYKYidvNSkukoBRfBF8FLIxUIRlFtyef9MQ8uRdBIsH
9G6Z3JCiECsvhapbp6KAYYhJPac+ObbE3knFnXQCdC6m5a0Zt33Zm6DncWhPQfVs
tg07VRvfnCxrPdBbXfEhJ9nP2usRvddvyPyksTPCaKr7T6XDskbcKpOImrKAAiVz
raRhAGSWTD3N2Zdn9v8Yo4zjo2RfZ4W2Qb7MGqTYgqmFGK61eVIonC1WfTYa8+/Z
djkF2c8WHLex80udq4F1/2rXAoA7bTo0H68PFrvnWN8rWC7m9E4rrGPSwzaHV/r0
86Bp0z0nTYkjDE3kLVH3GkKF1cZsH6OKcTl6se5okcT4kmqvBcxLhct8EfLxp8UE
V3nVbwnSE5QBn2XbTGLPAmzQUOwYOTku/v0VdaRL5d2cIXR8qb52DIDoqD31u2er
gNyC9/mFYrqWxD045cdshMRwJxiSKPI1ur0YDChRB0jRwlEtPrdqETsWtA7Svqjn
TJwwtAonirUzbD/4sJQovVbBSBjD+UdvAFW8RQNUYCGo/vo2m0nHaPvCG78ipIPl
D1wYiLRIdM9PAy3IC4C9nuNGFYirK1ZF3xjkMAlT8t+/plct28Xaa2GYIf17c9Uf
ycE2/lFXlXNaqV2hW+BegLVgm9JVTUTHsQfQsfbQIhQLloeZZlYaa1zVgMQIEKA1
kHG6sbjcB1u0eZ1CpxOl7CTt6RcnDvd/89Aa1h+H5LjIz16jkleV6KOCynWOIm6q
C8FKXWp9sG0HBdi6kGUJOhh3SnPzz2RUhbi+Z6XdXJPQ6mKMuWGw67Dkx5GbfMT2
/ULE6z7jym9VQmJ3tdgNlSCUUCFzxE8W2tyKl9D+JTE6baWAQHSVgfCn4iH4Xt2R
lcE8AqRAq4K0cC08HZg/4sjxhSWK9upxpVf6hBeIrDMpccud4e8cgDNzkf+WT8oI
0ZYFCFG0zrQ615HjKZy0HCEYzH8VZUqjq8hV6ugkp7spum/Hwv7rnbscrb7z7gkJ
t9gI5JPS424WhJKGeLYEoYhbZ3mcel0lLOE2fk4bAK3kM7xfuxB8vB0nyHM7MoXM
Ml+EyDcHAXNEUismSnf3USTG9VwvwEf/64jWBwTOT4keNoRjpMLS6DB6KfUqANX2
UlbNm9Ph5sAjZyUgYBjvHCmQVDmpCWJctmK73LyjKLkSq/MOUuxRSk3yaBnvfga0
8ODDPL80Jt5zf/1qvPyAAkyAryueB6zfsX7I6SU8OZiup5cykcSptQqXPGJZj6c9
DHlENLezzi+ChXp7WgUPDsSgwqxSn/oKiNujqB6LiZQdQBT5zOSLu3EjxdD9xHYu
oS8nu4XcXw+wp+Fk2ok5QQ6s39r8HFlz216TvzRMMv4nas3x47x4Bx1tIQ1hBy0c
m+sBXskyab/0mb3zlAGkBOFN90mt8sIDOT2uhP5fnld75/zSsoeYWlbxCultRSHx
eQW/feIv160N+jUSama7noTsPk96vsXSaJdF2CEuuiwEzkn6+NTYbdhrqAwdu4Xz
pXNUUXXyFXlrkfz+FFA4v6bS4ZDwZq9JXmwU1be0qsEbvzmLfMhfgxTqzrA0LOj+
BvqNdI+otWzJSgpGbrTfDE2HNfjtj+j9HbUnY9cLd3UJ7wfS125MRFPSGnERPE9w
O8gIIyo1i5tIFakVk0vZM0oBhN8uq5m+oerLpsdL5pqwGhWdHVlPjjq3MhxIF8/Z
9luHejliIGKFpUtQgIvr6eZJSEszW+c6pimgp3zaoB9VxxZV1Pow9+b9c7PkCU6D
nIEDOdq36GybqBMyWD4e6pFnspbMzDCoh9906JD5WWt6i+QUrqxK/bTb2gn+VZyl
n4i7ElvLj1emUyE7vNoBI2EfNw/9NAJ/RB5sJamC1XBEizmhBLrTT6HyIt5HF0Xb
i2MHGy+6wAynyGWqDcvN/1qf1KOiwDqmyEhfOACZ+erkyWCs9tPXCUAmBYO7VBbR
+RCD8gf3by3BQpKnCdL3i46QAneYpqfuC451YFzG+jaxg75mSFVPqsGWvRS9bgZX
CwDoiopzCWXpZOTpOEpots0ANTxuXNRpT7nMSEF1JmbsIsrBxBLkldC+GOGab/TC
zHRfHBwxBI0j+bvC0x8M7tV8B/wtD1gdWpSH7A1KQg6k3ufrQl3M77xN/vge0n8W
UkNqZpR9VGd5SfC8PeAZ1XaBFauvaMlC7STIY+ZtgUGwLZaPPRijNQFAnQcD2q2R
lwdWSFJZPLuTyNPou2CqozNeOftJ1F5QV64vOQIVCrjpbFvGkwcK7Zm8Lid6vrU1
XFM2meAOYM83nA9oD1BQPE8c+0GHSCjEXf2opkPzMXgb5d9fNtOXcE9r0NPI2m4O
uBbSM5QWEm6Q9T6upcbufesd8mf5iv1eB/WgMtNHxI1aTOQHniOmIVFX3O12+dkp
rrIezcA4nC1LKzJpLvGPv2t7ukJSqm8qXxEdZrJT1GN83wKrAocKa1oyKjCJglqn
BqMyGp6kT//VmLG5v2bxAxPWXsr4Vry0R2I7dc6afYnmmY6ksZ12XV7K/OrmI5f8
LHQXwDkphmqq/tBPn+wze0giLey3VDSehAJX0G7L6R+jBKrXDe8loYjeCf1aIJ7k
DUoVTAlr4EEiFXRWIVoMPSWgnDkgk5Hmlo4UthWP5LyeetzUry6/4hZiCP5mkVAt
ohVUM9HikSR96Vq+m/tHnltNtIknv//HnIHRYes1aeIDzbQ//stbSaatT/Wumk3G
Abk8Qogy54/Q1fM5QnlEOsX2p8AoMANz/ET/NVxaYsnfLuKfkyoz1ZaFlgiPaFi5
KlYhDzixPlGqzC04rd4tOUxHu7cK1lUHAdNz8SakEeR4FNeVOncpmjsVCdfyKM2h
/Sf5/FqlwVjqClaa7pfnOlhASQ9KoyXFY5KsNzNoGq5IZ8AmW+ZqbfwLDKTpj+rN
x5T+E4WZpjZ4Bi436sgRrfoAZB3PPdCcYOjSUWCIAGmWNRJ793c3an42hRXed+hH
SokYz9zBZ+bk6jwNCDBXRGA5VcpyXW/gtlE5WesJfM5cGw492y4McT1/OhuLLufM
IG4unYRvW9LjY2tkvEvI52PfIvvn6rdA9rGKSjpj2oVHYBYFVz4Kz0ll4fx2jy+I
fu2B4zpjTRuvq73kzpd1GJKwNKyY81WiiCDa72t7Fg95dNTuYGq37E4vZBuiXK11
ZjjBX9tWi0xvtAilSt6HHIlQyqCJ7tw0LXmwFohlDGWKlaODaQ21vSvKVXlyfyp8
9FGR+TGJnv8OFK/BXez/iV1VC74F3NyouKLpx+2/e3eSyL4oiLPeCKrOdngTVumh
Ky0s3JXz24Pg03r0qJ9CMenThqsDPK/L1wq4l37o106wtsTELa1kwUZP0R3iKm1b
dKVQwP6Ing+q3t2iWf3uQtj+AwA00x7TXoeu8/BhEoZOKZ7rPw428vGq7cSQ2mdN
NzXCbd3pAk8UKJfqxcoX6DPmiW45eC53l83VXnirIAfawG+H39ZSRSiZ1HOwWhrk
vmOjnWXKsMdQq8GFlMg2XBqvtSC8pYD0fNeVco6YE0lvGHgAydAz+d97ISAWL0oB
PSl5CPm9AwEsBNMiEI6yQ+VjJH+gbBuo1k5Pai7MkAKF2B1dbX+OF+0GLk3hei5c
jHZ1YwtGyqTy43MaoomYmqMx3uPOb9/X0rNN+4OU+FEu1LaBHE8jk7P6whXIULXi
z0t5Uo4K+BCYOr7fCcyn6rvfy6wEeIEHgAElaEOTi/biKlKJ/vutNK/ErJ/mehFj
oe91ghTGTha9bFSZmdEiYcXqWVv5T2q2mDEIbfArw13LgjJ6Og3yxPEt+wWaZhwf
obWHSQxePVY6/vE3aBmn41a0dTwT5I4fOulyCij3uVrZVGoiv4B7GGNsYu6eWlwg
r1uSNPh1PU1mmS/Ml04iEL564+s9J5mTmWZ8ZI/rMKPXW4lHhVCjC21OszkYiPik
1rundS0Bkto1dgNRIzAKOeCJuYQuz5/GiX0JDuCVKYoWBphDUYj+6JuQQKSDGJNi
fJK/hj2BQ91Pl+BBfvWGVJik7HWlqvu87QAoBX/M/wrsPUK9JfpcZNNIoYIiCXz4
YzxeZ3NayGCgajzFQVjQfUdS42xIvoJ56K0bxP0fbsBmmxiPLrxpuKiF+KINz53e
2ClDbmDMom4OnN0/YFfOZBGX+Agx6PdJM9r1UhNx0jHmXNmdfM1J1kYT6TLDfyis
qv3nOCy4lDVFTWO8O2lgEny0qYHeVT92B58KC4BisMaD5SWHvF1JFuvab74zdxCY
j4miQZOl0nQYT99kO7Th8UWGda/xmtB4s0Ao2HLyP6Adu46KKXrgkPs7GNVrTPfV
cuPj9IIHV8Aii4XPJHDOcNqnxwZcjzzbHYuc/OR6fJvPFvFKE0N9J4RgJotNGfBg
oRyseMBICAkoYL/rcXbat4JI5/S7MbVN4Y77OImnp9cp0NRIYKD6Pp0TYQ30Ir4m
W3BZh03cQmy829ZIm0TYFUknF1Rz7FhsgosYplW6shzdp1Li1YGLciHKWDxzgOnC
CBSJeZP2MhyJxbOvGWB5JU9gIg8XhCLBcm4ava5q0ATIJ5D2AqytEMm3AoKRDC0v
mxd9L6rWU4inSyvxIB4pZKm25MjRX34IHnDOqCO7ztUFc6w1dY8CsDXg+wZLVXNe
5f4MIbMbHtTNUSUEJ7RXBFVA/twLINY3ptR8barSIY6TTJJsqtgNcBAbDSSsHpot
3TtPcYVjls8nW/oGVc2KX09M5nF7dmajRf58xgPeu3B22PnE4XpAk7l/1VRsfygm
E60ocfruFQZjhh9/Ij0AZ00WN76hNe0kb9XtJdGy0rwxPQkFIB2/d5ft3F3/PaXf
1ygLZEqV0O7JSksgPmKWX1s2MmXb1r4wfYWLtR+gza888B7rpXucE8cRVhu691It
zpYW++c12qmUBQHeJ9RrL8sc6+Uxx3TwEMWx3ks6+uyEZe78hlrQhg+cArKmsfbr
5F/DptJnpxK01PUqJjyOyFWlIEHcPsZPEBGQXUA5Jy2Bm+LVromTNMeMKTh4rtyP
YyPu4wwVCfAuXXSKf3KD+QfWBbDY95pCpvFJYifRiKmPENvBK02GXj0u8nhg3PYG
zesEmyqJcZ3hdVJUzzR5Hbp+iIXIhuyLGR/3qDSW70EbudfHcGh8v9iK2RZigyts
lEeOK9Rmx1BOvIwElt3QI+za1K2kpxlWQzd3Y60jHkJwVMZMPC6ga7AubnqH+FRY
pVykoqV9jyX7HsKlwngngYGf0Yf5lsrEM393jo0ZG2equkn+kzMNCRgwLld1v8RU
EI2Xz4sa9gcCpTm72MJzRCEB/xJFJEqrcBrHBYF4qKSZM7BYkWtlAJPpsz4SKI3j
HOHRvZlKtcnZkSpMLbUMLeWNgJTQKpWVYeq9e2G93ozvFv2mkJ1cj2A8R5iVAjBj
fy7dHTNaJhruMUb0c3iaElQ4cPJ+xtehN8Fs+HUyhT/I57huQc293MItD4C/m2V4
FuXsImJe+W7LRFyfLg+RyesXA+7StQW8KGlEwHY/XMeHMObVEzBAsiRcxpuPgN8n
F1joBT/4J9VW/mH+0c7dXG4XVKutBbRRxcLGs6sY6Y4HL0b+cdRcpvaW0684xZJ/
8l5+TzlQat4WPPV3FowVf9XGqTb71bwMOxxnTssEC0a4EzoyzivrFzsGvE++hnGb
9XD20zuHrcy4V3GtRSbgSw==
//pragma protect end_data_block
//pragma protect digest_block
ovehDt0or0BXzFcx6J14dY8u/Hs=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
