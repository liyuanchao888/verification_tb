
`ifndef GUARD_SVT_AXI_SYSTEM_MONITOR_UVM_SV
`define GUARD_SVT_AXI_SYSTEM_MONITOR_UVM_SV

typedef class svt_axi_system_monitor;
typedef class svt_axi_system_monitor_callback;
typedef class svt_axi_system_monitor_transaction_xml_callback;
typedef uvm_callbacks#(svt_axi_system_monitor,svt_axi_system_monitor_callback) svt_axi_system_monitor_callback_pool;
// =============================================================================
/**
 * This class is UVM Monitor that implements an AXI system_checker component.
 * The system monitor observes transactions across the ports of a 
 * single interconnect and performs checks between the transactions of 
 * these ports. It does not perform port level checks which are done by the 
 * checkers of each master/slave agent connected to a port. In ACE, the 
 * system monitor correlates coherent transactions and the corresponding 
 * snoop transactions to perform checks. The checks in the system monitor 
 * are geared towards checking the proper working of an interconnect DUT. 
 * The current version of the system monitor requires that cache line sizes 
 * (svt_axi_port_configuration::cache_line_size) of the various master ports are the same.
 */
class svt_axi_system_monitor extends svt_uvm_monitor;

  `uvm_register_cb(svt_axi_system_monitor, svt_axi_system_monitor_callback)
  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  /** @cond PRIVATE */
  /**
   * Port through which checker gets transactions initiated from master to IC
   */
  uvm_blocking_get_port#(svt_axi_transaction) mstr_to_ic_get_port;

  /**
   * Port through which checker gets transactions initiated from master to IC
   * These transactions are sampled from the scheduler within the Interconnect
   */
  uvm_blocking_get_port#(svt_axi_transaction) mstr_to_ic_scheduler_get_port;

  /**
   * Port through which checker gets transactions initiated from IC to slave 
   */
  uvm_blocking_get_port#(svt_axi_transaction) ic_to_slave_get_port;

  /**
   * Port through which checker gets snoop transactions initiated by interconnect 
   */
  uvm_blocking_get_port#(svt_axi_snoop_transaction) snoop_xact_get_port;
  /** @endcond */


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** @cond PRIVATE */
  /** Common features of AXI system_checker components */
  protected svt_axi_system_monitor_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_system_configuration cfg_snapshot;
  /** @endcond */


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_system_configuration cfg;

  /** A semaphore that helps to determine if add_to_active is currently blocked */ 
  local semaphore add_to_active_sema = new(1);

  /** Writer used to generate XML output for PA support. */
  local svt_xml_writer xml_writer = null;

  /** Callback that implements transaction XML generation. */
  local svt_axi_system_monitor_transaction_xml_callback system_xml_gen_cb;

  `ifdef CCI400_CHECKS_ENABLED
  // flag to avoid multiple process getting spawned to sample cci400 reset pin configuration
  local static bit cci400_cfg_updated_on_reset_done = 0;
  `endif

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `uvm_component_utils(svt_axi_system_monitor)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************


  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new monitor instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name = "svt_axi_system_monitor", uvm_component parent = null);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
  extern virtual function void build_phase (uvm_phase phase);

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   */
  extern function void connect_phase(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads that get transactions from
   * ports and monitors them. 
   */
  extern virtual task run_phase(uvm_phase phase);
  
  //----------------------------------------------------------------------------
  /** Extract Phase */
  extern function void extract_phase(uvm_phase phase);

  /**
    * Report phase
    * Reports cache vs memory consistency
    */
  extern virtual function void report_phase(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  /** @endcond */

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
   * Method that manages transactions initiated by master.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_master_to_ic(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by master and are sampled from
   * the interconnect's scheduler port.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_master_to_ic_from_ic_scheduler(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by interconnect to slave.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_ic_to_slave(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages snoop transactions initiated by interconnect.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_snoop_xact(uvm_phase phase);

  // ---------------------------------------------------------------------------
  /** Sets up exclusive access monitors */
  extern virtual function void set_exclusive_access_monitors();

 //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_xact</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_xact_cb_exec(svt_axi_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_slave_xact</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_slave_xact_cb_exec(svt_axi_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_slave_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_snoop_xact</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_snoop_xact_cb_exec(svt_axi_snoop_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_snoop_xact(svt_axi_snoop_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_axi_system_monitor_common common);

  /** Gets the system transaction corresponding to the given transaction */
  extern task get_axi_system_transaction(svt_axi_transaction xact,
                                         bit delete_post_get,
                                         output svt_axi_system_transaction sys_xact); 

  // Checks correctness of data for transactions that access multiple cache lines
  extern function void check_cross_cache_line_data_consistency(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,bit[7:0] mem_data[]);
/** @endcond */
  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
    * Called when a new transaction initiated by a master is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_master_transaction_received(svt_axi_transaction xact);

  /** 
    * Called when a new snoop transaction initiated by an interconnect is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_snoop_transaction_received(svt_axi_snoop_transaction xact);

  /** 
    * Called to override the expected snoop addresses in system transaction.
    * @param sys_xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void snoop_transaction_user_addr(svt_axi_system_transaction sys_xact);

  /** 
    * Called when a new transaction initiated by an interconnect to a slave is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_slave_transaction_received(svt_axi_transaction xact);
  
  /** 
    * Called when a new transaction initiated by a master is observed on the system 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_system_transaction_started(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);
  
  /** 
    * Called whenever system monitor tries to associate a master and slave transaction.
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association Indicates whether the xact should participate in transaction association or not.
    */
  extern virtual protected function void pre_master_slave_association(svt_axi_transaction slave_xact, output bit drop_association );

  /** 
    * Called before system monitor prints all system transactions,
    * using this callback user can remove the unmatched slave transactions present in
    * the sys_xact_assoc_queue.
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact Indicates whether sys_xact can be printed are not.
    */
  extern virtual protected function void pre_unmapped_xact_summary_report(svt_axi_system_transaction sys_xact,output bit print_xact);


   /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact  A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void pre_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual function void get_dynamic_coherent_to_snoop_xact_type_match(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts  A queue of all associated snoop transactions
    */
  extern virtual protected function void post_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

   /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void post_system_xact_association_with_snoop(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void override_slave_routing_info(svt_axi_system_transaction sys_xact);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_check_execute(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_system_check_execute(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);

 /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual protected function void interconnect_generated_dirty_data_write_detected(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual protected function void master_xact_fully_associated_to_slave_xacts(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * In some cases the attributes of master transaction are required to calculate the slave address. 
   * So this callback can be used to assign this xact to xact present in the system configuaration. <br>
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations(svt_axi_transaction xact);

  /**
    * Called after a transaction initiated by a master is received by
    * the system monitor 
    * This method issues the <i>new_master_transaction_received</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_master_transaction_received_cb_exec(svt_axi_transaction xact);

  /**
    * Called after a snoop transaction initiated by an interconnect is received by
    * the system monitor 
    * This method issues the <i>new_snoop_transaction_received</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
    extern virtual task new_snoop_transaction_received_cb_exec(svt_axi_snoop_transaction xact);

  /**
    * Called to override the expected snoop addresses in system transaction.
    * This method issues the <i>snoop_transaction_user_addr</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    * @param sys_xact A reference to the data descriptor object of interest.
    *
    */
    extern virtual task snoop_transaction_user_addr_cb_exec(svt_axi_system_transaction sys_xact);

  /**
    * Called after a transaction initiated by an interconnect to slave is received by
    * the system monitor 
    * This method issues the <i>new_slave_transaction_received</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_slave_transaction_received_cb_exec(svt_axi_transaction xact);
  
  /**
    * Called after a transaction initiated by an master is received by
    * the system monitor 
    * This method issues the <i>new_system_transaction_started</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_system_transaction_started_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);
  
  /**
    * Called before a transaction is associated to the master transaction by the system monitor
    * This method issues the <i>pre_master_slave_association</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association If 0, the transaction can be associated to master transaction. If 1 transaction should not participate in association.
    */  
  extern virtual task pre_master_slave_association_cb_exec(svt_axi_transaction slave_xact, output  bit drop_association );
 
  /**
    * Called before method print_unmapped_xact_summary in system monitor
    * This method issues the <i>pre_unmapped_xact_summary_report</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact if 1, sys_xact will be printed. If 0, sys_xact will not be printed considering that transaction is not matched
    */  
  extern virtual function void pre_unmapped_xact_summary_report_cb_exec(svt_axi_system_transaction sys_xact,output bit print_xact); 
  
  /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>pre_coherent_and_snoop_transaction_association</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact  A reference to the system transaction descriptor object of interest. 
    */

  extern virtual task pre_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual task get_dynamic_coherent_to_snoop_xact_type_match_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);

 /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_coherent_and_snoop_transaction_association</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts   A queue of snoop transactions associated with this coherent xact.
    */

  extern virtual task post_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_system_xact_association_with_snoop</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual task post_system_xact_association_with_snoop_cb_exec(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * This method issues the <i>override_slave_routing_info</i> callback using the
    * `uvm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual function void override_slave_routing_info_cb_exec(svt_axi_system_transaction sys_xact);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * This method issues the <i>pre_check_execute</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_check_execute_cb_exec(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check.
   * 
   * This method issues the <i>pre_system_check_execute</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_system_check_execute_cb_exec(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);

 /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * This method issues the
   * <i>interconnect_generated_dirty_data_write_detected</i> callback using the
   * `uvm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * This method issues the <i>master_xact_fully_associated_to_slave_xacts</i>
   * callback using the `uvm_do_callbacks macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * This method issues the <i>pre_routing_calculations</i>
   * callback using the `uvm_do_callbacks macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations_cb_exec(svt_axi_transaction xact);

  /**
    * Called before the system monitor adds a transaction to the queue.  The
    * user has the option to indicate that the original transaction must be
    * dropped and split into multiple transactions by setting
    * split_original_xact. Transactions are split at the boundary specified in
    * svt_axi_port_configuration::byte_boundary_for_master_xact_split
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
    */
  extern virtual function void pre_add_to_input_xact_queue_cb_exec(svt_axi_transaction xact, ref bit split_original_xact);

  /**
    * Called after the system monitor splits a master transaction. The transaction
    * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
    * Once split, the user can modify the split transactions through this callback
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_xacts Queue of split transactions 
    */
  extern virtual function void post_xact_split_cb_exec(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
    * Called after the system monitor splits a master transaction. The transaction
    * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
    * Once split, the user can modify the split transactions through this callback
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_xacts Queue of split transactions 
    */
  extern virtual function void post_xact_split(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
    * Called before the system monitor adds a transaction to the queue.  The
    * user has the option to indicate that the original transaction must be
    * dropped and split into multiple transactions by setting
    * split_original_xact. Transactions are split at the boundary specified in
    * svt_axi_port_configuration::byte_boundary_for_master_xact_split
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
    */
  extern virtual function void pre_add_to_input_xact_queue(svt_axi_transaction xact, ref bit split_original_xact);

  /**
   * Returns the contents of the L3 cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit  l3_read(input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                       output int index,
                                       output bit [7:0] data[],
                                       output bit is_unique,
                                       output bit is_clean,
                                       output longint age
                                      );

  /**
   * This function writes into the L3 cache via backdoor. Backdoor accesses are
   * direct accesses to the L3 cache in the VIP by the user in the testbench.
   * 
   * If the index is a positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @return 1 if the backdoor write was successful, or 0 if it was not successful.
   */
  extern virtual function bit  l3_allocate(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                  bit [7:0] data[],
                                  bit byteen[],
                                  int is_unique,
                                  int is_clean
                                 );

  /**
    * Invalidates the L3 cache line entry for a given addr. This method removes the
    * cache line from the L3 cache for the given address.
    *
    * @param addr The address that needs to be invalidated.
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit  l3_deallocate(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

  /** Clears the contents of the L3 cache.  */
  extern virtual function void l3_flush();

  /** Invalidates snoop filter for specified address 
    * @param flush_all Flushes all entries in snoop filter
    * @param addr Address which needs to be invalidated 
    * @param snoop_type of the transaction used to invalidate snoop filter entry
    */
  extern virtual task invalidate_snoop_filter(bit flush_all, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr=0, svt_axi_snoop_transaction::snoop_xact_type_enum snoop_type=svt_axi_snoop_transaction::CLEANINVALID);
  /** @endcond */

endclass

`protected
P.9^+85Y1>>UYBK&?52dR#8H<1[[442_3/_/a/99CNE6U)9XRGI>()P97F\A)BTR
PS,fHHc>,>-8L8Mg(c)c5G@LfXWC0[TPF8W8YeIGONYP95=:N=86N=8dc.P:3,f>
2A6X&,^R#@Vd;\F76\4V0f]/ZA2WZT;e:O7?]?4S?;R;.6FY\\<BA_,+9<W;KE6?
V\E<X@:VOXT>F]f.0-]]FX&\BOIZ##-OeNRO7J5>3FPV(QN76eHXSQg-U33.PeU#
\=dBcLG\07V]>N4cDdgU5IJI];C-CM@:_7X==@aXT>[a;?/5Dg.H]Z):K0XAHQ0L
.,X[a+.JY9cd?f9U_,R&<6cKARDLYUKW,,;<BU^5M872ITM3G1F4:]9;@Be0O0/4
SbY:LBI#:6BX,>,Q(T?]T0a9MZK9O>E>7KD@&\H2&]:/;?[3\V(5YDa(95A_O.G&
F,bgCK-X@^8:4-]9e++ED.RR07]]JLR+YT&[;H2Z2+T0KG1Of^S\FS(J;#2USYA)
<T2?IFU:W285[Zd6\^=-1@gY?XeT[5-.Z1_g<ID[L]<@d\INcU+1W.8,+g.5NTZ:
Y#E9R:,HC#8N(>eF=g78AY;e;OKDQ]H0+7(L4[,@/7MfO3BQ8[Gc)Je4+4M?ORdK
=+)[^DC>H0T@ZE_R4bF+\];,<c=)MA#fRO2W4].E311^Q6I-8GRDLZ7KZCA](&.E
1.g@-.CBOFV3dSHeX)RWgOL6.9TTdB;12fF9?2(=>81B]g))P@>XMFV<+@=d]&4<
\[d23beOJ29dJ4@Q9f+ZQN,T2;9]I&RCYL:<<VK)+<QUK3MM4&S11)3676FD^9WI
#_4H=F2/8aXWC3+-_-9,QCOKUF4&L,@5\RL8DI5g?G?UE$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
de3(HbGEC9dFGP5VRa[5^F=>W,+JZZG21+cf\D<R\.KaPI<bCD8D)(&YH=cMKJB#
9a.Ec;4-)KKRBY0SV-4&TgSTYgLF51+W7_>ZX5gH^21-gf:+Na(,F#KgCb&CIGb5
?2e_;7^6=M<(V&4+FZJFd\;DcNc<BG>VN,/8&cAAd)#R)-ZBZ>GfKP]J;Yf;(&)8
#cg?G&@X-#UbLI?d0Bc(XJ0b\^P^dFd/-.T\?OV(24HG9S[:V-I#Y<4^]b@<OT<A
gZC5?@Y\W(4JeG]eb5</2UIY@g/DSeYDXD4M,(3,K:0bCLEC8W.4OHc5#S^8IbVT
XB)>\/0OT7JUD#gA;;]f2?Y[KUb4bO-<7MTL8T)Y6cc3#.T3Y:.1BR[bE]1H\H?)
(#9UYH/LQ?,D\:[U7]VgQC(6ZR?Hf.:cP@F\E(-bK-TgEa-O?;Hb9[=@Jf,251_c
\UIU;CL5Pe;O_&TP_:K2F;.AG^X6,+aS&MJg8DcT>2Z3WRR[dg)^A:D-?^ZDQ#HX
UCC:6OQ>;WI8<QYEU88[f7c1V1VMeU<=.]Ad#d;Q<-NDT,+1+ecVAZOE\TFYXa]O
@V62?61+PYKb3.,<80M7c7,6F8(<SIY8f/.:#X[MVHSLGb5^^fC#:B=IXcI3Q\ff
Y>O&RYQe>Q^WGU\CKJ+KBOLXP)Me8\M=K7G;.Q?4ZTXRN5DMRJDcg4&6(Lf1_V>+
bf@J/fM/@Cfd@2X1bVJKSG^7d)H^,\->M&&96Xfg<FJ>RF0AFO9McQ/FC<eN^#GI
BOcY5YQ:4VK;GCDUX._0#/Z#bV#]2TGBW1)+aO7Nd.65;58_4KY.;B40#eQNaUSF
?e,B]WT8;gOaQa5Y@K&)X](O\R@K?O,bXN\_6aS<0#:I\D6,(UCFMfPP@+N2YXE,
#PTTf_Ff;NMUST18eFcJJ,I8)\W?B,)_CRKZTAeB[.(W@X)(>,@9\W1FMRL<M:.U
(;KZT;8EWZKfIV0,3@#D-1\\@+85-+gbe6Pf43(M#@(KPg][Z[5>[Ibee7R5@gAY
^&f;NUOP_(-E<BV0FF8ZT=78Pf7H=4aX[e-@Yc+G/+=VU(4T_=MM5-4+0KO0_CE&
]I-3G/NJS8^FX5S.0[^O/ZeB91Vb(6)F@#TJXb[LQCdW<S^6fB>>.?WEgZGQ\fR\
@5:a1B2I5>?)LR]E?d5OO]-[5BL>U#bfb(?#M0SFSM\T3FaV:,W]V-.2>-c-9Y2&
eSdI6>Z#dFdMU/6112-QT9O)<P<97YI.+-/U6XbS@7RW9A-?J>&Vbf2<&G&a&AX<
^>2=BHOU6,/2-D1(RJb5Te,gE]S(4/Def[SW0(.a6-)MgIQ(;Q?1MEFO&g.U83cI
Ag^.TC[e0:.Q:==aDIEEI\_,#BV;XV<+-.&R4e\aR&KM3Re7HXK)UUQa2AX@WBFG
CP+1C,B3O8KR.5dJd;490<,0[1W1X0++bP4A/^#_Z>8_&6eUFYU-MWT@<N7ZBg&^
;f@?/TM.Z;)7P]c42117M7d-;a<PPaYP^e?]FP))#DJZ2?IO89<FG()OBF4e=Q_2
,a24Q(-ZKT.CDD-#^OdX(^[<d3?@6M+#eCeX@><5Z?N\0-Z]A;5a?N,C][M?O5LI
#8Kcb#GS&QJ#0>J\7K^H6CBL&O<GQ#YIM]H9EW=\SG\a^5.=dY63XM3BV0c^cZ?T
#4#96XAJgWZ^-,aIZ<60e9ZOeSFHHBG=^_:J-4@CMgd>&0@0K.gM[^d,P[@eX29g
/#bQS&MJK#>4U5#@a-R8ZNC6b<(Q(.G0(E>]KbS6X?f^6\gC^O0G)5ACNVY(,4b6
RI__1=4+L/-bKU.::ZSeW3(,FR5-,XCM@@B,WUMDCD.>YX-0J+KK0I^LNO3:_d0N
;QA?=.U#(EK4.K?Q_:K@A).48ZG)&Y9W2.e\\QV3-TD7L)>I;fV[U^B_^\f,+&N#
G:@K9ZF@A8=DE3+88I:4;?ZXDWQ?&_T7L>#1:@P8Kea0Y.SO:,8Q7b=6@e<ZXS5S
JBX-<@OQPI.(,=,ZO54.GOAZI-;DI7:B^9P)&MVDH7(8+Dee_eAK9PYdY^]d&)K6
>2e>B3+.6YeYPW.G7KI4VL-?:EMVbC5I#3?EZ#=BRK4^8\+bSSEU>A@#(@V@[Be,
+3T89XIZ7_7T[&J?T:&ON^[Y&F@:<KLJ&g]d+LcCMHa^S@c,@L=J??-?6B8?]_CT
=ecQ+Fe)Y4=80,+E4TQ/LOAG6gEQ\Jc\LO@6>/PGC3_^C33XD)E-[6/KH=BB:]AO
-21VB51/<1b-V)<d6=Z0[G+Q]V.<2Q(N9K:^6KND([@C](4DFGF^9AM1U7KTcT9P
[De4c>1Ma0N=G]YT^+HP6e.I:aMX.-S3S4G:]a+X-+G+T(R1A29UT5<QCAE0-AcH
L3M.#:7aaN&B1D]0](U_&gJ(Rd+#8;)HP/#aBK?+U6Dd<H[d..-MML?O1)?NMP1#
Z^2^3)/b3d;B^LYZaSdH/<WF>>M:1IW)Gb80+c\<B@;HT-fBJ(.1QEY\YENS:f\J
\8]f#[Ie8gD+X+RGW]=P]T20-aW5Yd,5L(ST&EN_/+YY70c0_I?K)b@@a&PTRL/&
C<P,6ZT?3.BBCd(QUcQcKDZK[=4@-@&84;+U1<#c+eV,1FPWAC]@MGXIXaDR0CW@
Z?V+VT[1N=GHA^6AD+5R+V4TNWb]Q&Hc=>&3,HP+([>b@H;78-UgcSF,H>d^=MX)
YRJUZ]A;dB>OG92U28OGAU5>R@B4H2DeN&Q4B0>?Z,DX;;Kg\84H;d1JK[+)c:H9
8e\\#-Z\0:BCZU.\8-N9b8UTA=1aRHf=NS)Sc-0>:98XU8:e]H&IE7c]?,JISaF]
\NST?+R?bHG2IOS0&.gO/F]FR?IdR;_H]c0g,La0,Z<]2\(T^V9?NK+D;6R._+=2
5^gc+:-:5]I(>^9g3fY3TL;RT;?&_RM>RXG9BFaSP-V#;d/NB&_d3[Y\9Sf,>Gdg
dB\O<6IYI8SW3G21/D&B6KgI/W:,f9?+J\&:Ng3DUNXN7_U#]/./4>?L5CXg;d@R
QKc=J=><JX6[I<@].Q\:0X>ZSP<P1>D]FP9OaHARCL2KCV=?9=STVLgH:4&\:f<P
O26^)+K_#7=;4WNZg&)A=@Z4PROg&2gZO:0IY_CD\FJ@g_32RWeIceO//a49fA48
MNS-)\IZ9K3;,H>[4b7RS2EPY-)AXbPBC?FY&^V2C>Ha4PZ-4L9?c1#9JAF-=R9<
1W4g_11eX(O3JPL\^[-RCB,TQ5f5.);>5g#;FRd20<?e;Z7#eY+#P;<fO1eL^f/(
46]T@F?X1@++fA53W@IN1#0/QSSYFbXdE^)5,G5fg/2AB5#,)Y\47c;OG2_5L,Q&
&5>ZX6H[2(eO:5_6CX9=6c^W?J,Of@1;/)0KL1GJJGfM/Xd:_cFT,Q5MD),JX8.T
<7,/2EW62M=N?WF2-@[>>2L/dg[7A)^GA^<L[?IE3M1f?-gD#/WK,VQeL,WQ2dC?
M,BBYCJI54ZVSHfV2)(e[C7Q)W,ZV(X;\OQHN^fO4?DC)K38IR:EG.K1J@O\/QWJ
C?->LF<bd6W<[D[6L\#AS_74.EGTTgNQDgH>Ke_S4<M5J#]]Rd?9WXN4B?G[2M.#
N?VG/A.fabZA<gEQ&9/I2gG53bV7O7g+JD@LNd>UD39\a[FF,WB+Q[]A<aQR71eX
IH:Mf_N^KCUWQBYXN2f]FFS?1+UYQE[f:MdV@a4^0ZIT)L)2-bD7b8^JD5>)gfEe
_^Q9XDKFQd]@NH)JGEg=34[[f0HSg7DT5f^O,U:5UM^/G7ET.;A)^g?HE\M58g\_
[ZYXY??R_]8Q)XSE\=TT2<-Ef+TVU7G]X(@)I>R5.V]9<(:(JRF:ZQ=eDCCeKa>I
3+2R6R];1@:/AgOQTDNJ+I&32GA>+AJ1Zc(&SY1.a#X;J)/+_[AB+VeP57<2VMZc
ATQJ4a#H-#?eTUBFG(T3=#:\IEf;\Y@9WH@/U46)Udc9XEOY&S2f@aL05Y;F.KF2
\&_.,URP#HWgR=ZPB/eeW0D;@fO9J,KV\LA/8<dH3BMSN368d>ZF3f-e2_OW9[b3
f(cF]bg)gfMb\=Y_TcI^Af4[X4aFJgE=e;5Z=45SeOT4[<ebL^B9Zf[\MXSbd/3>
N[XT,]TI8YRe)c7/7f)<Fb=<[d#19=MR)B/<7@4U3,\5?Q@J/^I2Y?E#A<RSc-.,
JI3<1)cI@>JZfL8P2C7V<^:/JfR7:OdfHBEBY@XDBbG3;,&d3M]8^?=2J/QWQ8?]
)e^I9TNJ?U5I#XQ&T_B7OPC:G-D2WVFF[FY.V9,(<#^092(8<d_9e/VUeV6Z-cdP
C_TC&XWKK_C).GT6L+4MbP.[U84HPcEDUKB\FF^V>gX;+(-6;T/gI/.P3GL_Q9^S
BW7X^F<))#N1:\Z.1aW/;?fE#-e8b+)H3K[A3H:2C/9+X3bPVSB5fa&=M0-?]Ee;
QJ8Sb3LI7QJ028,BeA/bM:S-L.\ZH7;I2)P7.XNVID2PEX)J#5M<BGW4O?J^B(D=
-R3ZE=\RZCC18#U.F:QB4S2.S+D1=)D-a9gB4AT>;-9:dPBT2-&:#0M@_0EA,(G1
EHQG-\.KfE69)#5aZ4KBG59^R;c/@FbF@9JXI?@?YQPQ98MS;+-B9N+I1Uc-]K>X
W2+R.a:BbA_5.K.@5cB4&>#]>#BWbIEc@-N)IPW8bH,&HcIeASGcC]4IJK>UTZ#J
V+,_Q51:H+-IdSFJ\WS8IH#d)GVQTTLZKIG.;9aYB]RU\fFNQ2fQW#)0QQ>8M6fB
.M)+^1C@LdFVRJ?A67dg?_Qc)2Oc7FZ)+B8\0N(LWe9[]8?KU3W-#.f^^CG4@0L(
)&=G2)7/?.74)\SSB3Nf[Z9Pg8)-GC\)EIT=9;XT7#O7)#8L/BBU@M:30GG]NM>Z
]_:2E4/EHJg-T9R#UeSZIbc-LETF_EC.39(,g1UAUZZ<d2bXO,AH6S^4><8ObJa1
D>Rf\HRE[@X^J[UUBH.<#g+;(+;fKbM:SV&c6Q5;W/RHV\R^6W@KZIRZ9U)Q+3W[
78P+<X<437BdZ1&,WCgJ\CAZ7KJH&6RUZZef8\:O]+^]T-fRW]M5&d\2)W4QYU[=
b:8)8SNK7S.U&V5_-X+XcV\C@6N)->?A7J.9XDKfcIF63K<c/DfaN3E>LBfD?>-B
+DeDT1&40<Q&9+cRb\XMW0///-4HO_af6)gS8C,91#[8Y1VH./(>_(ER-#b@a[F#
M:[^UK4W=(;WODT]Q[]GNg?_NG/D>81eER)KI-b(QIQD)_@ZPHRGNGe5GaG)593V
MI?b[S81M1C0&&1a6+/)PaOVAQ[e_d9,C+g4K,W>Q-\#V&R/>A\Ad6N\6KQ>O+KQ
1F7TJ6#D;G&UV;?\+7HP\aVRdT8R7Q@8f1WN7ZfTRg#M+;>L^c17&:\;82].;bB0
[0A\/KcC^K?/Z9[-=MJ<10Oc=fMfLI;;@0KNF?(63Ee1&/DH:NMN:<>-B.&M35W=
I[#-71N1g,];N-)0)G7&Y0^a);E2b2b^MO(MJRLD=RPIDLOX?&?IXa;EO@+feNg8
C9W/Q3-fF[b)0OU](U[7<HAVD<W->XAXf9dGD=#E[g39+])a.O/+[=3J>7/a,V70
cJ4M^d7DHVXZ2Z<@faKPA)VOSfcLK6TF,?SH_g/:WF(:C.G410(]3(fCX<d^HcQ\
C#EccWcPVGcA?]d-5OG>7,W9eWgL>JG&..g2F+,g=:X7RVgT#1>>62BM;c^@8/5>
HEcC7GgUb#E0]Z)f^[HL]_@-1<f#Rf-U4c;cgTf,&.(4:]+]ZSg2U>WL99+L@71Q
UZbWZ3U[D](6ECEa](W^ZW3eZ?(S#OU)1QF.]8\;JO[,UdbIHcX/(UK7+1D7NQOM
.\?C3DDR\8].@<MOPZ\GbBG.\4=(&f3cae=0XcYO/;NIPeP/XY=-/2e4^3S28EdR
(#B=Ka;?<gb7B/E;LcO0K:<<F;6PPRJDA@=RgP).-f]E\:=baV.3DU.^>^UE_gIV
)-DaYLEGGDVCI0.QAF_.I1_d>H(He6S:@5C=FNd\J1HL&?SFb#8[=fG872,7acP4
YC;B4UWX8B^G[G.4@d4FfTeRUZ2UCQBD4GW@(/?O/a#g)<U\G&(ZBCDCULTXHBE;
4aUJ<5#F_HLL1KJ.R-VC+c5RM8)(:<TG.\Ida93,-@\A?WX_\gfC?3&?K(W=C6D^
>MU:S]3W]Q.DN()9VY]5YaYP0.\LVaeAA6<g>,8Q>#QAO5W\b9#d._H.2:HXSU,T
1;M]Vc#HcD[3:b]H+1GdUCGgYK:&WeYH^;=50dXR)5.-)X-ARH9_5&BD;/ZKg+:0
Q34XJIPS[?#[+B>-U#C(X=8.(>7[&@)G,cK^2g@dJY#KW)B?>2^CP+;]/+#;c3\5
7J4;9B)V+C6I?G++d\[S]W9-]WI)\>]D^fAH:@-#g&YWW^e:[WE;XMGO#2bO5:aO
:^Q3XEDSF45c@<-Y.G.-\;Ma,WR-cUd@+3V=TNDW^P>-OH8Y4>d9)?E.,Ld0#WBF
T_g3@D[c4+b\4SG]IH]-DE[?Q2Q]^La39gE5+G-e@+H1Y1NT3>DV._\P;.7IJ;9F
g9b4O_>[@WQg[d;P=)CRd,VdJBK0V66<#dV:dTP0d:2YNE+\+;\KSM/a2:3MPSf9
3D,+OF4T[VWXD>&H1K=)P?NZQT#9Ug7,9H_aOM\a7(A]&a:UTK7(\<NaYAd@2T35
c2UM<7B2+f9ZEB\16.G9/aK2;>I^ZN2<OJ#,4^5#CN8X+H5XZ^b;.<2Z6.P6F\U&
7<POaC5<+E6[D(g/49N>Vc1RCV?6XAMZ@FEK,,,7f;_@<b3Qc97M;IH=Y25I@A:R
HU3@]=RHBJdA]#SN-PRK=+Lc<[cJMOMdA[^T3<WH/,,2L;fb]fUNJN3_@F3RSYN9
WDYbK\J&]0=&aSRJN4b.LF#-d+MNIV;8U7K_^KVK??]50&_@HWS:WEST#J1#EdFb
T?25Z1&&f-Y_UD>ZYJ)QG8Q);D73+E5U:U1\I<P+5&O7b@#>Be<2#NE27+?X.=[+
b:QW96S;TDK44#bVK&a5AK8E[2L9X8E(A#Y_SLd;4I&Z[H[3S/C;UG4V-8dHG67@
gQB9MOe,+A\54?]G).4>a7<6_&0G2SSWfAE2?>e^GW@;B#gEUV:[TQ=gaCd71>4=
d:MOb&9+(J8PDR6ITRNdPQ.W5F37Z@@;KJ4/@#TRaA<KU4Z7eH(^?PZRSdO[8_Ue
S?+T9AQRTcQ>B^VN+<IPB-=UHggR?V[E46YTb,>/T6[MJTU#b,\HV0::;g.AQa0F
;U^gM7Y>J/9FId=g.V/LKZR23K3W3S^bH^FH6HOB7XF?&<4)<,YL.0S^Jc&W)LQd
CY9IMD7<7\VGeV>=BcYUWd4daG_95MEaS[)[:cW7Cb58dA\AX#>Q>gZZBVbKdDV)
K#GgO<PdFGLHaU5T:5PX:dAM(-0TM5[7]geIYWZ\^,3Zb57EASI-LH)\IH@=.R@F
XU:FS++b_Mb1J_Q+#[RWU&R1=OWX3gJLR@\IT^JCU6\JU_e)FK&d0O43HI=3FH,^
;_=d@JYEJ9BK6-JDTV?8gW:E=39R]@EYF/f>A.;TD7T9aSbC07Q(W3&b9C4d.>JD
W=dP(^DKSWRXMP9>/^J4S^B#G>WZGC7HbZf1^gUL1agF5@bSgNgb@OZgE5^@:\A1
8F4=:R(@X&/U&#Q]P#;@3:LBK=TZ[a3_7?-TJdO1T^)6K;4-<>TJYLeQBO8;cS9J
-g[FZeGY]&Te>\,5[Mc9?+-#21g@67\DYa^]KYFH)BU;^CO/c:T/I-HMQ/Y/d5?E
IEHI-9]e:LJ+S/,MV@\LPIUfHf3:D?9dI^Q@G0+[fge?Xd6a,3SbQZ<e(B>FIU=a
.a6Be9>DOJDc]2-8XD]L=g#51ZaF_A)MN8dMRa6<I]^/H2#TU9-2_^1+fI\5fIRT
(5E=a/5-\Z9S7ffOC\X5?96KTWS;/RQ0@-D9]g_XW8L6eQGJ7KSQS<Z])d+cB\6U
b29C8G_?HQKbY8ZW>[7eZY93[BR[I#b=-X5QDDS^UX8<^WWMg4DeZGf69a81Zc<Z
CCO_g[e.>+5gPQE5c^C18\g]F1?Fc1-.JS9..7EGWSD?:.OH,?_;59(fM;2I59Z<
2aOD6L#X(1F^(>LZ:&5GYc-X4bSG&dSOHBM^RHJCNc4\:#9?0HBe^Ga)5])X^/+9
b^5MBAGeA5@H>?8f/Y,.cO@>A+U<;g1e)-N)A?D]bE:2Ueeg+97GICfGAT0DB0<E
:W<dF&\9T\.b_1cT(E#SX/c2);cYPgYU]]Y,U>,6WH[[>9b+d5]bIEB)<MG(RI[Z
_HCD5SQ8U<=+PEM_C/61(+(,IFcW@V6=XEMDQagD8QOS@?W@S,^g#fO#]GcERFH.
QKX[MM@-2-E1:7&8_JgF00N>C))aN/V+TQ;A:4QG[J/<f_FEH&7dX@^LeMM:/ff#
>Qc&AC&8Y6:+.JP(2^^F/NT#@J?=;==4K&2;T8-]Egb6?BTWB;K\A0:fP3YDU)YX
7-+))@EcG^GMV2=/b\fBg3CC\ZVV_C)754?_AbU-5TF9O/N;9?EXCMHG@/E7.?ad
6@5)#]I@<g,5K,,I,X-^e9D(88<1G/WdMGYI^YVc7NZUMTKR8GE2a0DA.Y4+R7-d
X5&Hg9<GO5ZQPA[DQQf\2C=&fVZ?76IC>R,=a4+2W(/P;ORUTd#J#K:bDO#,LH^A
<>UFTcKNb<Vb)a;e8YdXQBTAd1a1fU4XFdbD^II8fdN8cSTV1;.5<,--@7[gD@1=
Wg>IACR9&^R.47W>MW4gN_HL4=0.93CD1/H1,4SDF4fG0:?P+(],[R?9&5T#\G[V
#2CENOWPH#61]L>2A^HYg2.\3Q6013+JK.LE&T[TH5]7-fc&5aF&\#0)AMV<2-G(
+BPH/M>+Yc;ASaC;>Z3GBM1JY24#S#XRQ8S#L\c7N07HcI<Q\<<JA3FS\]K6Wdg2
\NXTaE/E3>HLW,QYAEfX?@0#V-g&Aag>L()+]UL4gP6BdN<&-:H4[gfa)U/I=XDG
,LDa??=;-FJb_?7/:d2H:&FcERP<K_:G;=8\IETRb4_O9N/0+:U:/2S/SX+#LKXW
aHMH+NYKNK/8OU4dMWJf[H>Y.9TTVcQ=SJ>8-cW]26JCX0]X6P^RIeA^KbPV(c75
MF\E&&I@(8YN>W<ab-2_UO013<NA2N@JMM0CQ.&e1?46.aaEX1/Ia5EZ4:UEH>G5
P^J1A0gFecWFg@ER8^UNP=T74ECVBY.Q4V0F-R6B]_O>N4F4T-QeJS)4#WU.44EF
5CKEW_ZW<MQ=);[Ec706H1cFQ@W:--6]V;4WI<831)51R^NUI3bO&g\FF2.DSVKC
FTHdG.<Y#16#f)&XPB@P]&:Y,391;+^T.E,J(J1)MB-^C2ZBD@UIYgK<V0bbbW,g
3&a17U#=g-[I)a03&/N\Y-6>:LJ5T5AfH-2d>FUOD=)?S2<98SC>H@[^GI29FK>F
G5P][(=_3>FSa-(S.OHgc/4ADMQa8^+.S.Ha\c^C8GbbKFE6e-ef0.?0NW;ML50M
MK(HfLSSTa[43(Xb=\4@.97FgGJH]eAN,C46L[571Ae4J(aW67;):[bTaN_gUVQS
3?><7HBM<[QZT,3HE=(6GYdK)cQ;2Hd6P)D.1Fg./R0VD[gY@1X-L3JUGL]C5<Lb
RcUL2/N96Db3bMG#a2(6+8-g6/<43P?;@ULEf8LO<V&P/f+XYG:PXKTI\DT5U1C;
Y\0TTP(<9aY)\1ZO^a3;AT.d<P)^&b1:-b_f/X-?=3a5TDB^^^Q5<DWg,@DMX-d\
DDI)f@IN[;F/\4JH3/63dd)@9TAZHCDKSH+VXCOg6EL>0C,Og>;4Z[HIZUcf<860
NM8VOZ(5+,+eZV^[FTO&P]bMWbO1U;.1]>0ELE]McCXfW>_f87,e>C&e\1U87Rg#
,IDS1^/RK[U6-M=OFEM]S-R(@3HBMS8YZ7d&CWfPcMWHRY@:KJg18bR27U2a9SN/
7H[JZ@=+@5T_S&H:[_HF5A[@6V3)M8JDEX?9SV0+)&KPN/:W\\R4R(YW1(A]=d4,
:=NC6YQ9AVI7gdcUVeI^.=](NXASASWCG\WR#4?=JB3b)#O7LJM<L1VBWV24,TB4
dQV6?#+,4/X\+)9f,+&MI=9R^?<YM^YXP?]EV7O=3cFG=3FeH@L.S#1)L..@?IW[
3]]4[V[Xe?/WZ1IFTP.B=-KD2_KTU,5[Z=PP<-NHfIEcIgdB(])Z=U]1&C1?PI&7
0XS.;HAb;1H)6TV-58a/A:Sg>B,KgQJb7_M3\K)F8F_08K#3O#cRbD+?+C#9R2)/
^:0H[<3C8Yd5aP5/U6F=NOMZAQ[H6-8--4^(D-&cFPV?FNeM<R7&H+]C;>c0X0-b
O6XJ,;2A:3;+9eV8F9)@0QaD#3\(F(=+9.(P4>.>Q1c9]H\=6fI0@[;+CE0,(I;[
?O8R(+fQ@@9_9<C9>29/2M)8HcJC;/.>gD[[QH;9X+1R,V])dG;MS\EHc7D&)=6J
@I&^LB[^Ia47XfUWND<=]/E\]R:KV4&_#CH05^/AcMWQ,\&=L83YN/&XBIa;O[Xf
UJX;Rgg.fOUSGM>41)\<a.5a=e?4;E)TQZJOO(6S3+ENCU+H>Qf#[W^L;F,,)eE/
_,FUHPOCb]0\L]^]L;(ec9:&c<@2]f#N8QX38<)ZY^7?.A1Q.6;,5-HOe6f(CG0G
)f&UQMa2L?8eI@=\ae(fJ]+8I]^E&2E<a>G?c/F49P,f6^^P1e4O\[\J&>X[WN63
6(0I)Te]_=Z@AO^B=NH4\0YK?G9FPaDIdRT@DF60UP&3;_,_@8>@9A:cLGW\DR(L
9B,IPF-g^E1A:;)6T6[S(GAd1YFS/6J,,]<O\_VegD683KYVUM82+DCg+a[0gYXW
TdWHeA?[A7f>c-,(OEfOA_N4=YF3RB41g=PV1-S8/C]]0<&VHRac.Y\C.@J0<(+>
^OLWNKJKH/WY=Ye(d\g[R2Y_3?<1^AXJA:Y8aOH3MPg.+WCTg1)OZ?T<,(0E]:+^
<E3,]09HU.YJ&D7Jd7gR_+Lf;)C(R_P1Ud4d+I38]<K)+:-.8>/6166#LQ2:Y<36
Vd^WgHI[[eTe#f>8E[N1+>QJVK+9>FT<G39.HH2G0Ff;,S(M)(_-_]K/>bF9=IL.
G7BG,,N>&O(T6OW#V>/>[HF\c1NQLMH=JFg6^^af9,Z09VAaOBL;BFG4)FT4XaC4
F6B/3L=^;#b7,/2Bb;-\Y\SA6@<TBV;7KE5H3FS/?HZVN[PM@gG-XTVL#JcNGcI@
J9f4LZd&:A2cS@H.5@V2QB8KaL11Nfa:=?U)6\ScV?(\/KP)-MW6/6C@P-]3><PN
NdS:6RH@D57>@(8^T6C\@=<f=R+c&dT8OV6@0-A9P]f;P-\>A5WUQ<2G[gR,+,H-
g1VUGWTZC(QX,#V/AVCV1+58g&AB1dP8Y8?.9/Vg?_F>+8\XOKGFQ;PAU6SY7<YN
?;7+EJ/AW4&CS@HCg/bH)Wd[#=7H#(>ILB/5U<V3WQTdb+E<PNBeB_.V?PW:H3?M
c+U_ZcU?XX77QPC;LPR.4ODSae(Sbb6<2)ePeafd+2DbIRab)T)e^C8/7dE0L:-.
R-4>bI1]E;)5K1@V,(;#V]T46a[g.TW]#aXUKM,SNPR<YFKD80#9)2IIS:G>(gD/
Q_bMDT4EZ_CJ^XZ:J4M4>4)T0GOM+SU_E#g(CdH:DU3>A@8-^?L-I7Y6G?(LP9LO
75OM-I,E56DX0e&AQBV>Z)aU^3c:f7N60a[F&/6^FE>X,Y:^5)>f]YTZ/M@G:bX/
B6=E2=Z@V393.1/QUE.XcQFQ)JbG.OOOEFgH/ZQ>c[f>f\/G)_0;98)C=1?OBH[@
K?A#,,^]@,&P&46YHVdSZ>E@YQda6RKWU0XJ2<;=6))#BFV5+,Ef(X55Fa30J[ae
]XaT7,1)24O5f#gc3)7g;4A-)Uf5aR3)\SA&_P&:\E6XMMF09)Bc(?ZW.&<RBB+[
&DR:_OB9[g-)5d8>3KHW3Og6@MJ2Jb4=/2gY2OS2CagHdSfe)@JJ\(6R)L<YH2]E
Z):@;>[N=U6[T6+=7WPeQVDIL0,&8L2&[OQ3J=&-W93EWR9CC\;XNaeW.@6SK&\b
\?/)[C79>2^N41C(9H>;-/D?]/98]647]Gb(aW5b9g=O^I-HD]aQJe.WaJNeV9fc
SX.)E(E@XT+>RQ1D9Y0PJ&EEED\U?CL+D,Fc7eZeOA@<2,71/E9+I/-G=1E,F<G3
NK9S0A#e5P]7CR:-ebGeC\?GD79O^<]XT(6Og@_g@f?Z;0T?3c,(2g,J.>f)S15J
[DO;HUA^bNJK1,U_UZQWg#@R/D86P>W^e:<.AC<G=S5-])9[N,RGP&R/F19VD1&S
1<6^+9=#a7#HB^QG^L29/Tc>M0:f:B3QU[Q#Ug;4=>,3(3=J)\J8P(KbLX4[4_Vg
WGL0WR(bF3SWH^gd@FdP=<EYV7O:C0;g1>WN+M),gN/f=8MCGXg<?J0/Kf46>FA_
72GU5B1g]#V=&C:.J8Q360.cDDPD+8PMX;I_&3aYVb2aaa:,3-E_:gbF[<FY+2&T
P/T#JWPMTLEOFRZdd4E](/&@\b28f:TE=P@E&dKETZ1.FgX7Z6O=0eQO&\3?U<R6
=g2)4:S7^:#H(+=EM@L@J;+>#4SMa@8FJCZ<9JgBY[N]I14VXI,25:./MVNg\+1T
C_8<4D03]@Y)DV\;0^_C4.1_c1Zc.A;LP)XL:+Md8[-.T>=MP][:,]4&_9X9.[+H
-ZJJHJ,<I(,+K9JaZ.9B18]Z/FG&IJ^+.8)]>?+-]0/c3A9_735_S_[RY_fQOZN;
e(F,,SX\-M]<7_Y-;]RH(LaTP(ERZe71,I=6<8?)VF@FEb<-D^LeQO(]=^,XLdGA
^EV3F\G9X62@e28)P7g>1@[#3dbW8WB,fV5G><8C]eA-NS:8#Z4IEK#MFOLf_V7;
V8L]+B6gHEB-+O@2FFXON1d]P^X;Y_LZ_Q5Pf@b:&fRg77O#1^aa_P4c^(/(BBbR
c:K/U]OK>-aTP5EYCPga^S_c,)Qa^15W_7WW60eZa#eaCM(@9Y;,4]U>FdH<RWP/
.2UTDZ=MDac#NST+2/BB:S6[9BSaN2c,^(Z&SV#gVM2KCf-U;CQSFG:>X6(/+dJc
2RB[dI(^\56=X6A@b6RFC]OPWP+3ERR=W-1(RXDYF=42<C>DG;^(4_cR]7^/_J,Q
<3^?N6XF4BEI#YF]AMVTBN>@D0Y:MPRFH2\+VAfdf?_5\+HGO8K]&P:N>[d]N(:H
OAM6<C[Y=)f1.a>A).?YMLSHdO-Ja+g72E?(D?ZXFK6/9=KD>IG_&6567(Q(e/4U
V,IQB>[^?=/F7OIX+=a8>OTA9MJ\.]AKe:d#:T;5cH)DB8;>5T\]C@<EP7efK3M=
S7V0QYGL910a#R4?ECP34J\\<\,.bXdIL]de51b\]J+ZcG@[;;c?8W]C@fX95:3S
_=,)2a+4-5fE&.KY,=/f9)Ab?R63)e=Ca4RdfeaWEfM\P\5_K2Z3^MIBE(ORFWc7
EAKbgRU.OZafMc(]2MaV\XE\^3KWJX^#-CX7UAJ<8FFSVH)FEL3,RXY=]7;e8&E+
.SJPb?>OgJ]\^]4S?)IaK<8RaX^eO93<_O);X<gWF@<@ZE75cb3dUa4?QL._c8D0
+ca>PMSOeGaZ<YFY_EgW4#1S.1\?ZEMLD-(VPF_K]B8cW\.U5.I6^8_bgBW>D?7O
6W88>CSRL)Q9&eAR)E=PO=K:gI2d^f/1baG0O:491B5UaZN:AY]Oc[.40J8Z5S4)
g<,I[B7Z-]:RS+e[P=W^N,WSVA;5ESVG/1)+8;,c6@5e4?7WgDg&VGYTM0:Wa_KF
KTc-Z\>3]C-LTAUaBO\-_]N:X+[N_EV9BM(BB:4,([_31Ma)YaA1@H#AC84U?G@+
.L,c:c@[10,9+GD6ZPO:4f\;N8JN9]fEJTSRK\2Za0,A]C/JXMPEBC_]RCe2:]7)
.@FR5]/<W8e=)SC(8-S=dNWYV?g9[C,aA^C^32/&d@2X2_LS]F]#,OH3]O/I=^c[
cY62JPJJg7]=9V],3fA)0T3cbDA+R#^eAJbC0T^X;C@3g/&D>c8dRJ4:R#5V2II;
6gc3e4K]LD6eLMcYK=[6]Q02:M#(?6.SLbLgI8<+c_@5)W\U=Yf/\+I@8,d&aI<c
^eJ>XIH\]Nc\.eCg7OVW[;5.QG<9RY0L@58.gcLP#0=f9(cO]G)IM36&T3#d,^dK
;a_.gf-V:3(I;KR/+DeA&a,=B26]dJH=)D55fJg?X0RU-<&/F;4BXTM7UZC^TD[N
,.I8VBS45PAQ,MP_#N@VPB/eA(2N_P1XA1gJc@9-IU3aSJ.=?d:D/OA=<7)_CTZB
cG0UG0(\O9NFOKWZa<J>M+C;8.ZfS]1);ZdIS\QK>1SJ7_^NVTFE,,WSgG]X_2.C
Z&U#LU3c2N,)Y/^S?<#d?e23VfWBT(Y9@bN:[NF[8CPODg+b[666<P+YQ?b(D5bW
VT.&eWM?.b66S#O9YRJGT[?a(+&ec9,Qebb8OK3B?Q]0bPdB/.CG81Rf?(MPAgCO
EGg2/DLCJZWKfQ+D>XP5H1#YWZTJZO<8S>HQWUUL@_-Sfbdg_NM@_0^b,D4KJGQ6
b&;D9++gPV7d=\QKD&b@G]2TYL1NXQTWFV8-KEBa9/5097JK)b9S25A5@LGX50V3
\SXQV)&?gF6?2F\R)PQP[JX_6&WDBNc_8=OZM)\g95+[],HO1;S46J&30>.gE]AC
C@5L5;eQ\D_Y7-P)=IVK_^QL?GI;]\)>2)49^6=TRLbbM#B.(1:DNcZH(T<[>6FJ
\R\gJ<)[K<\5dGR#4_0J/?g)JZIcMF)N.^<2@C#O^:JgN>WG;D2bdII=DR=c8;U\
7HC)A>Y4?+,STS8R&d/d+f?=+N^E0-8I+Bf\d5bEcc;4GGE[b.QC@f8?M(&_G[P/
_KU^e,e-NX6NCB<V2)3^JPb-MRT)f:W6QCc)N:e#YXR^7VP6,1,QJC0-+>,T/FKc
2d3M=G22=-#Y[d+FFR^]Ef[^3Z.OV:C.?07?BE+-&c1#M@L28M5/TGaU-@]9f0gH
X_=0A;BT\13L=OUND.(K9UX(AKWW?)FX-gBGEI)D,Q@DP3NXAJQgQOf-B-V,II6X
ALYdFQ)K7R-R4KX1R1V[U>)eR=^][>fG7QJFB\<S92#CP<7?H:AFdd)+(\4b\X9R
0,7ZdL0FCSZ;>PT]b,B=7#=Kd9)^)^:M46]3(+LF94--?M2V5KI?K&2VUKa:QF5=
B4DW]\T2[=<,S;bX;/Ed@WX.b/D7G[Fgc3\A^9Ig5N4.QVM_CI5cMKJZ[DU;]Bd8
dgR@b>JP-e/E<8[N1MGaS#^[@\bAeI3c-;4:?.2RgX-9ReIB/A^e].8BNG>#984K
b)H-b6@/@3.R04P0\aPE^2NF^6:CdA6G;[1dA514O:fLa/NHbIO^0ff@K0gZGV(2
+,;eJ^cIWfc&=X5eDa-;-X6Sc&^dY\fc1XFH.^&XY19;KKEbDb-Z.W#@LBR\&=KB
RVI_02&Z,X+5Sb,L7VNbR2-FU[2e/KG>WJ0IZ?MTW[QMedN@-S++^O[T@_(/b@5^
FbY_D<GM^G&G)EG7.0e/[>S>&Ca@F^[fcOA[fCecZNI@^)D7;<A[;+ANPSSY&).E
09.\UXPRgH,9<5YM6HL?a@9)I(eMET>^M<ReC\LYL;FS?a)I5N>Q49g6D?:+-9QU
)JKS-L==+64+@dUAb1)P0;CN)0?2^@4R=NF(&69KgaS\\^#Ag(20S[M@K5A\5Z>[
IKY5MN;?5DX@USOVCcZ+T]C/H_<1T[,)&J;_e]_/&6\f.NCW87.+1,b>(W2?Q]QQ
cSW[TGY4O[7fGTP^B63N&EAd.0>T?A7FFb,0Eb@A+T8K78A/W7R1BSD]2.aRH>R3
1dUE60Vd(=-AMMd(W5F6=dYAb@a6#gY=\S9FWTQ1=3)Q/E99H,]#;_-IbAddbSA;
IC31>CNM)AYVd@0LS74#-Ue4>ed;\@<<OT08a4I#[eKS0Z?[CJ#4RMTgF-,->Zg=
TMfW8\VbP?M;bN]8JFM/&QSC4U>L^Y1dWKb-2--OLLFYB17,&5I[OZA#-S)[Sf[,
>):fPfSS8.:&.>#LG+AQ9YMa-0Kd51ZC+UE-I.4)]F-AO6>A3\D5[D;a>2GHQ0.5
,-GO:eI-Y.&F9eW(2(Y_I=WbA(1U1X8Z,KdE5K@A3\L3IGMOS#JIBcbFFU.gKF;L
GB(aZ102#^a+0DMF0-E:SdHF8a,&XG,15;[N:&.c5fB]<(FKQ/Q5a6^;,(Q8+./3
e[<Q/HHNdHGD50UP9<[Uf7/?0GMGHSOE]XbS-=G1]G[3Z&Y5CBH32\.:_ZUb)gXJ
S(9&(0G30-2f[?CMDA8Y>eTf&9X=):,TP2K#RZQ@+NYW&@b&dU)JY^/B;H;M+ISG
GL\)XGa&N@+HMH)+RA]MELG7S3?HP:YB0AZe)E5[4UNI(L\J^W@_TWR8C.4:a+e]
AV2,ZgCEX_BG/V6^=b/WU84U5g<^-M]f+Q5&2X-RC6#=+bBG_f=DQO^IN@.3>c:I
<_2]NU47NWY?#TMH6E7XHH>NPXB_O+K@/gW>VQ5,K#a?N]GU097@A+:?+aC52QL)
:-/B_<#B0<[.O5-bbP5B@61JeZ2bMYW<]2OeK:S?J;0ac2,_CYC0c2G:420?EZdD
:M^3+V(-QcZ-L@Q_JUGgVKCVM>D5&@^(HY4^aGL3EZ5BP@_cBY12T9>:5;GJF-4f
W2KVEDU[6KPd-0>0LG&@72B\1/V#4X0N[+VZaZ9>+#(#/10bGZ^1(L/bU:UA)QM0
fTM2[<,]&RQ>X+?1<]P?S7X]##5VKZ-J:;)OT16^N1F\VY]8137JUW0.5c;O-(VS
EB&R,,HEUU9dSB9EO+ZddeP,A3+;P<e#gd@+QIBgdYKVg5V)_0S<7ES5V,[7>PG?
D8^FA+K2XdX#R3aeDCI<;7g#_105-;6?,69=PdD)99:KFJf4V;\T/3JPbNPe_(f.
_^e>T3LL=URK(1b@BU/L>_8B2QCW/@VJWWVX7LG@J)4;1CH&JRU51,>L/N;g7c9W
7IeJS6\(f_]2@3LHfN@AXOa<7,0-d.[V<dFe<d/K>AF>,7(,050FA(^+83\BeVD-
2LEW\0Z@g5=,:f:I<eI-;EHbCL2RO4TF8Z;)W6)K>#^EBO&E5V\c>4]R2a#fEXQV
gPV<TJ?8Z:MU0__<50G(0_W8CCJN+;Ya7]&>8>TFfD=#)C1g=KU@Ig4\)5I.9K:R
#5FVf?1b(V#JH[<VE9BHZ=GQ1C&1-b[Y8d?G8@7Hc<IC5ZD-c=DVNI,_4X<QHdU8
2-V>&]@DD0LDGVV?K/IB.U<0>Zd0d8dRg[2=6?M;]FddLN0G>7?<d0;QZ>g#9GBE
GMJ;+d)LF(7O3DbRM07G[.1IWBO&+I4-L)D(a[I:A;5e.YH6F&18.=T\7S#@fCbU
743I.WSI^_?GNZfR=^7EN-Y?,g,[&/c.[BX2I=^^]1U.BBYXR@&;@0KGNXCg-B7Q
OT06NYJR&[];4b@9b6^SC8-5(eO=^ZQ/3T>[63JNVTW]FQ9#)WTQKYN.:G5-@.O/
H@9ZeO-F\;^U5W(GaP?28d+SWM>c\/\b][G3W3,Y2J#S1.0N&8B86;Y&#FW-eQ\O
fP+(YOMbQ];RAHGN=g9QMgO_IbFH5Ye]NR:@>4OZ558DE5U:ZL3/)IaHTY+\^O(d
F1,M#1T/U)[7^N3+9-.>G?U:0SA:1_FUVSX\2=5_[JE#/R=dRTe.=L\,DN(=bK=O
ZR=&06cXEL[?2V-eWRc&:\-+8<5KJ85dK)Y[65VJ2AT:V[F8E#CDFS<3<YCP2C#I
GWdePHbG.+fN-8Gd]VVN_]P.6:5-R5&eBQf1/Xd4@P[<,U_JGQPMgbd)2]9eQ[-R
BA&=BHNcLe3(/2P[;P3PPRH@)4E0\O-c<LLd:LdG^U?2d+^K+\\:MF1/TV@5-16\
F,QQcSA\>fc3VX/UX=c/3>F\E+I]\1]+)-R+5^f/TBUJVISQb?\]6;.bW5:/DLXE
.>/a8g5YGB@<PO3N_WgWGD8X/DaNWL;bL/4??_,a^ba]0T)S3IN;PNEPP2-b1e0/
8SI3gR[CdBA?F7cEgZ1<HZB-K,b+&e^6TZa5dcIVCF+&XOY<ge>SLR[QaUN[;^A/
PX_4T+^)dbb4/7<aJRW393LEKII\[:@S1ZV]BW2H/M=JA[9-2a#^V-+T\/Y2R\F1
d9NL\T6Q)/Ge(9/][SSA1Y\XXP^,M9?WBN[g?]^E</8#L6XY?XUNAT)HdB,^F32.
-Lc]\d20S[EDbF,H)HMgP4e,+H-K<f.;\MPa(&FO=Z7fFegXY9/18#X]:c-:.Qcc
OL)DbTA4>-\V@M8+3[PMQCD+=b:-?W7W6<aa[X=MaS3=^DO8SJH-8W0D9.FCaZY-
0dE,gALO=C4@LF<AECXL^[L_Mg>1I8=e.(G3AJ<=?J(?M.1TRD3=-11L;BJ_>EOK
M3I^T^W:OH2Q4[#V6L37eOHdM.W]Y(.2^<ef14B>J;?6=M+QWG5&?e6]OTPZA=IT
g,_KUfgaUCEYCLbKA;N3-2f;NM^^Ad,<UQMXTNH98<G2#@8Q>W_39)6cf.=(R/0Z
WS0BB/(K5d=EE8YN&:dKL,K7<IZD3A9\JaB(NA;4MH\HMD)[>>5/7(2b4CL9X?1O
P3=MJQ/1dSF7DD5:K7f9gJ<X+(]T5&OLV_BNe-N)X?A7I5K(O)F6f2VY.E54aDNH
9UIF2TcR[JF\TTG9]&7gBI&6OG1;^C3ZC^KTB(NQWAcU1F/_LZWE0Ff>Xc=>d&FU
A?2G6S+8RV(&+(_8/.6LMR)A_ddZ0C4XHQZHaE>?ae=R,][W+8SM_N<)Td881QB-
_SW3KXg.&:)B8OH_dZfRN@4HW35\-9>[QAC)gO9fDa1.[aEA]8T02aeE5a,(&3cT
FXLeSJd@f,3F3<A&:<G,bJ:SM4:K(7NHJ++8_A?XTZg(>A/;9]eHK,P.V5#LFb4&
:\0M8>R:0M^3MD^Ef0XEc+b8KDPJNCM79T7#.@E4W\WN2(YUQ2UL2SS,,P?\W_B2
eb&/Cf/3EV5B7FRf@@35TGcZ.6\(QDe8@3dV-c-ZS,R+_6)#VM<O?)EV4V-3fC;S
24g<5S3F+\.c<-@(>UYPR:+H:b@bXW/FA125Z,380WGPQ&7Be-1V@14?C:-fa>T\
&;?A2BbXKE5AH\MK8.Y6</;4HUBTMLK:1^W1.F[.<fWd)6QEf>3UgVdY:[#P4KBU
UOeIY]-J5TLI8D-Og.FO=d0J4[L:TA>bBA07@G2/0VQ#bXe]-L\WE9S<\(BXbZ7:
JQWB56]./<bW&_^+DFXXKcO6^MEXa+\CaLD]=#YNNR,fb[-&Va)#R8H^(PC1:&:-
OLUeJSG?_EY2-cH9JCLQT#SaI:#YdHFAO6G&XU4>,YGAV;O\\fbJ73bZR1ZeE;2D
<2(b=PbU<?CXFV&BdQ,fS@MZ3f;f?^9<T]4\HF[-\/dLD5f136)CHX/[g^32;Y-.
S.4]TcE,UaY#/,4ef?UMO775&^M.?N\>K\JAKD:&PC==QP#4Q0.1>deV\/3I9F#K
_f>6?)Q^4.5WW+)>TQDAHZP^8&9^:GGfW>A.]P(L=UaX#A@<TDe\L/.M:F_>UfTG
f4E[N^IM-O^+\G1Z70JKa-?Q(]OH67];(cEc902]A+IZeDTOE@Ub?(]e[9>7<NU(
+:_G5\f,cH1R_M1,:F/FI1I5L31gBZO-eX7UEIL,BT,9,bZ=AWId;C)05/RNGIM:
X@QaN;<I6d7AL]^S&f.UJW/<T3(A<(]aPH20E-a-IU^>YdgBGZ>1DS@1M-D3?Gf,
YX(7/&Fd4XMd:aZ4+Fd09^8C5FTVA;)?9PgB#44cH;dJC0^?YKCQIK#,MVM:4^K2
fTG#F,+YMDTY0,R?G6aI;.efJ1b-g6BHS7E@ZZb<MU\GB_T25bNHcaE:3.C3R,4K
Z&_TKUOcE?(N7,79X/fgbNEHSI=A_/U.>W^2B1_JEa+FOB\dI(JfYO]S;Y)MPT0S
g\U[I4,e)f\[C_MQ5AZC<Eg0Jc&ASfN].2]&5fA/dF7@A[W78W9/,Vc?ROcdLRQ0
gNBU8PF^GA^JbWR1ZKN&J?8[4)?Gc_SL/ZA;)cdP(c8;SUGD6Y)eJK::G0c?Od6(
@]^EI57ZQa6C(71Jg9-@?<eJ#)N,:I#V-:L/(?Z:3b]&.OL@P=V90da9WVKa&]C[
&c4K7DD##2#AVea#<0M4=Bf)546N;VUdII9Rg0Bb^Sbfc:DSY;@[MUM3c/4(c=/X
df>[a:/<D2HPXdAM.((X#O#DK#H1eQ#&AR;#@9JW-J:YK]VJf(gAQV47+K//VUP@
<E\)-9(41JY290aMc.V^fOD@W6OJ+09Dd3P72\8AJPV^f3e=gY[Q\aE^4@SgN)-,
T)(6I[6[ITZc8a[PaCK8e?XTUR2GG>fKS)F-:4AK,,:<JPXJaCYQ836,TI?QXaL]
.VcU_I+XL4IR@E).ZK?TFRVV3(U(eXG?\:SFL>c=)DZPW[NF_fTQF;1c])cH/<YJ
8#P0U(&FCTJA4\@HS8>]8b[L4aUd:Q:aX+-1fe^WT\7(#>[gcV)9N0=<:;b56F(J
TbUWQB,3=.59aA_MU_UPg1JJOee1GXLMSE\UP-Pb<<9OZNRV<:&K2b156&JV=Y4c
ZU_.SGVFTAa115[L.5\3\W[O^YK^J?5?Q);CRH6Vaeg\Vg<6UJ,_QJH:HUd>+XCO
I^M39^@U:X3]NSd#83+QFcO3B:@dZ4A(gW72c<L&GA@c?c+FZ=C[5T2:T_(4a5d:
GEA85>YIdb@:Y:K+/e\g+E;-5Y@[d3Pd2+VH&Y8[&R^FOF/9TUgUSR1PR^27NQeY
aH(]0]KOWV<ZE0_e9=<.cP8:Q-P(E,a7Ue2;ZFW&eU4(b#K@+FG?5c/V\[2eU\ae
MgL+R)QNKdJ0,Q:c_P]AN7+[=eM/T+:PA(3MY4&9EDKAbM1g((.##b53__J>65dP
SG?L42ca1HE1aL@(K/L26A<Tcb+8W_/,7[34:4>V(g,ZU8\EWc.FVR.(f4R:8a#b
\P#_HA;-g4IQaI8LOaL+4aG);^H2;_/)B>d_RfABPB:aNX)[/4Vf2>C^@:RdA7K+
4cDAC1@(\eOC))gVNW(dI5MOBLe_+C(,f6??O:+-6bA\6=R(KWV\UU@Y,1D+H<5W
^GQWZGYLM<.+=@3Z(<:=X>,RJW1GEbY3\O.T09=5d&e]4g(?G?C:=dOC.^Rf6c_6
+9B8,cMI-M10=LE7UQR9d8[J9V,7;;YP9VALYXR-TOXf+\/[4BM:36FR==S40X3)
DA/ELeTY>H/O&cA,E,1\E86c;EcHY]U>P])g&;?L/B_.fO(QFE@Q^c)E;O//bH7R
g:<:.[R+LH[,5W:@gJRD[@K^V,AcU]c8[X/X5(Ib#U.A#EN15U;Z@WOP/+Y;JVfa
WG(?XRZPH,Hb[12<8W@VEe99a=ICfJJ2COL;1g7e&J#;dce9U9d8DfGOHacIURAB
f_J>LX1H(-XbOX1;ZFdKZU/(=FI=&eKX><<,GICW0H^O#Z^Y.eVB[L7E2&7^BYOP
bMZ(,SNQ8VKN<D8N0cWNW[^]^ZX+IVeF;VDDSY]Y<b4-K7E=4]8cBI770L0aeTC#
;5)9<)#=9gP@Ze8:6]>ad[I3E2NEV:BDRAY?ONL?9EA@CIT]EBO_,>_fIXbTeB,D
2RX(Rc>3cZ.6W;f-g;e/cP](.GRdEKUP,58V0./FV_^M,TD6[(-?-A._)J]::V)Y
]1X#J(SAHePR+V6@0-B&c4N;JQ,KS&]US?KQ^f=PMWEZdCSW2Y.#ZJ>9b<8d9##N
/G=Y8XUSM9LIEUaJ;(@I+1=_Q4B+H0K^[cV]/GK<9aUUa<\g^P^gM+.I:^.g8U[L
?a>NV:\;,YLE:Z)U]QAHI/?@If2UQC;+Q=&)YAD[eTfO\&_feUg,JG#.YR7d##7;
\JHa4\BY#S@^_)U(gAE46Qb3Fg,ReKQ5P=E10RYPHgJ9YKbC55J/4[J>K.0K1&98
,BS,cSbSU&L=1E.FCW6gN<,g&LB5O\/E#WD/1fR,AKZR?XR_<LD@(BOTCMa:W##[
:IYc?e:S4\Jd2T7:X>UZ\P<IU,@C9(IIZ&P;/5EVbN&bZIG/eb0=f2+gW9ZIV7&N
OYF>=bZ]aBK<gY@S2(+D^fVR^F1dM8+ULR-EL5VF5[MA1A-)-J4FR)799fg&7&4>
dX,^J?CDFb^.C8U_L/B@B&+S05(aQ_U:VK6b)SK&LGEdXRNS+UX3YS>@V;?Y3d&+
LU0R1G8e]B?F^BM-NQ-9C55fD,CD;.Eb&.-T,,=[Y&]]=Y@X6:VRd>>8G1@7]3&B
=@^I(ZS1TaKP3?/OAX-G,VG/UMQ:.eB33caGBC&\#9X?54@T;SKTVP44P5Q<BVg.
-QBU-Ag?(;P50@I8A#ODc,EVL(QHa4J/2CbGPM9&b.+VJ_R5bX^ZZeSPge_BP=63
3NLdPQ;ZW6+B^Jdde9PCKcY/FcXK[UV=0NUEB/L-Fa9(eSB4PM>cY5P(O5dOe@P1
Ab35YQ,E_/T,]+,)(5D26De/&Z[\P?UJ[](d4gS5T8)4d]RV>I>LLOHOWdW7Z^BN
4?c+\)Z61AaWF[Z/K9E#.fT:O2[>@@(_ESV;eFIZH]Z5OO=^B7__FV_.FNg7[Y^,
XJ0[4+@ad5;+fUF4c9VBdK;U7V[^T5OQHZ,#QHZ+bgWOA&T)WK3QQ8bE<LbB-\B;
9OgSgNb4:A1;L24^bd2@@2?S0@9))9(@365>^)Z+,.1cNUHV+E+,b:f:>Xb,Z/NO
4IXH;Z?R;V<UVHe8aF4N9C,&TF[LBBS#>Q\[_N:7G4#EX\cS><7JM_^3+M^gE?B=
FLS?QPI)WZII).T6)M8eOZZddQ^U2+01\@6;e\BKR_6c4RGS9<N@d7Jd6P.SbN.5
XB<#SHJSa7@7\Uc2<;C;S;/c3c7feJ/2Q74B8&>=X7:8#?NEaC?1R;Bd+7?YgRV,
/CTFM[=Q^AFVT)caN6@Q+B/+D_Z&X(EY?@W_F72B\T)4c9a1/;W+T8/N7_CD1;HP
V+6_NCa.&V:d\1J#5+8Fb<acc+\YbV^F\f5Zd;-SB72aO_\&c/\10?M<@]+;ERE5
Y,18aE_9E@_g;P@ZZO>1>&SF?Ia/X?OFeS&Wae382bWVPfF^4G#;ZdbP#a#?aCOD
bRdD>]?aFL\TSLZOdHOLfK1(SJ5X0QCJ9a-FSa?[=BT4]8Z2&F?0N83P=GIOf7SZ
+Y_E0MN>^;D7\+LJ@8,^3I]1&>Aa+Q7:),QBf(@6\WGPHfX;S+G:]RO;AQ/=8P[(
@<0N?()O3-DPfe@](E]DN\V/&49L(&g;WS6fB/)e8P>O&\[X8b8GHI.>Wb84L<SC
C]#FLEZ]:Z3cOY2Ub4+HZaFE\<^)A3(H88O.3a;&<Mdf7f@#U[^U14G9Bg+^9eLg
1cB\.c[OSS#L.f^)F0P7N1@R05bUC(;6cJI8B&e@X2N+\1)fKOdHD]^=V-=.Gd\W
.[&]IDMP92<IO6M3W4LMNC+KccMBJ<D.3999&B.=Tdg)#I=HCPE?PL\Q<Q_V<&&H
9CfITW/4cK9A>N4gW+Lcd^&#UfOUb3;N6V&#e6QULEPceJA(H.[/G4D/L@[)=^WT
(:#((,2L_@@.[-87b_;?.4M.4HDTV].(5IFH=IcU0D5A/A]gfSX0M^.MLa6_TPFN
eP\A8JNaQ9NJYdEU>c:1H/aXg\BCS-XI3V72T;#T]=D?B(8/&K8EW)7dH8I1J>2e
@RCQY-MJVAQgM-:(?+=&_;1fICaOQfZ>KD+PcCT2RF]8#P<>2L/71^TS:aMZXcO[
@)V(<5d.FWgDRN)J9P\X^CPCBAB#XC/)<1J#I6IB@P_Kg=3S/_BTF#@<:f3]G+9]
&:BY0E@E;SVgN:IJg?DfJ+F=7KUZ?1/-a9_44D9g=U@S^&c-YNPXcf?(Z&)Z/,6O
V-\&NP\Y/<+?H[WW3N-@P&aZM3NGGE0)JVB;)3d9Q#^R,2d/F=X-^C6dQDOS49;(
bSD\9YNe63T@KN\<=Td2KfK+g&dOO1Ta:9Nfc#QDb@8Ge,R?)E8/f0W\2WHO)IVQ
SZ2>L\0^:9VA5VG>=X=+YWT/WK-0M]R4eE\E\.)c:BXBOTUSY437Y[0SCf7.,?fT
CK5C:-A1:>:YZ?UI8aN^J<BP2U^L0\KM:T_T?aB3;CUU7L8L0>=ZVSG)L0/c&H.>
.;:&;>YLF]<d\Q;\(=c=(4U-5:4;9F1_fdRJP2dLaC5=VVM<QS[9FQU5;f0.?PSH
1:BAK4O9#b\SHX;Q]CMEI2-9,T=Je?JU,T+OGOaM<32Sb]#0\1A.IN7.\)Eec55D
2FUaea/bWCgWeS?1-ZL1c]]LM=P3&Y6)HRTeHcD8FUK1&KKKNT3,E,]X97f>6&P\
b1[LM<FJY5NE3]KE[FW()KY]E633/fBgDQ3U8HCI25&O9:YOZ5_J63HDK?)9=g?Q
US[4KJGH&UE4QGL<C,@L&T0VH/d.KNM;6BAe9aeWd-\EKYYAL<gGP1)(bOaFM.8E
.Q;\?]e>L-&HY\8:7-?<aQ.DbB^OY79IP;)@YU9QSDKE+IG5UeD601]Ee6UF5NYT
M,BS]@^a59ScLY;]acZa@VN2K>LNJ0G?\dJ5+2\8g?74W?V9D5a,OQe+:]G&U/=(
ZMf(c=]=5WW;5d2:ZBcN@FfKQA(AU5JLg040IOFC)1C]2^R2,g:^+@\GN4cMK_;L
YPT(0.B8ETb=>Nb;Je&:YP_3X^0Mc0-^@QR+e:^E65c1?/D[cR&I7NM6/[N.Ge7f
VQS3e(U5NgS^c[f5X92Df[gC3NU8=12)\RG9YSFHGZ(ZaYF,SP@?C[f0MUO4[_(@
.[-I6]^g4BNPAXU4D](JCINI:/-#Q_FH\=JfU)/QMKC(4=^,C@]U\VTHFC&V^d:X
KW^2KM??]5GPO1#=3K\URF+bJ,T>>0HMeZ4IdV>+TJ]7WUVM4\V@N#2;e/BeJ&=A
aL_)e#&].=U#<,[CKBNT>R-KIgRc3P&2BQ8a_Ta#@8[Ke33>2.80V_I_<GbQP.5W
^+0]_ffACMe4#YM94=(,7PA^gSV/P_R3BaI2)@XT/Pb^08PbZM]0eY9@&?Cf[<d,
d<:LELfSf&8dH71)92FJ;>L26T+IRD.PU;1ZF6#7)CT=)4bULH_DKWIG6-:SR&Zf
Q]YCOV1d9+5W[e2M,XO;03_G4O9QK:Y.>Oe;\=]V,0dJ10eSeBEJ9]+eU5IZ].-Q
;1A.#^5[5^R)HADc(1DaU[dQSPEMWE4aHW.&TXFPD(Kf]45=AS_L<A,IR]/LPJ0(
HXD&dGNNMSTF@NKHM2:L[ZB&bKFJ84MU-XfN4MI7;5LTO(:LVIgBI3;:4<&DB1+T
bKEE;=:I=O4GM&3VZ3M3X74OK/0b<+5S/F9QUJb]_63)(<Zb9L<NM/(U7ed@b+2]
BQE75+09K)O8YHOQ2F6[1P(Ke2RGORe7NKg;@M_c?_#:#[AFOaF+E.OdGeK/54g^
<62XaCcLC/Kf:QU)Z-DV567aO;gQ&?6SNb.I[gN[QAQRf;,1DVOX<HHZZGXOA9+8
a]6CE_GgA/1Y(0.@I?LcFAgE0O^7CP>\;[\NQKAC<HcU/NXEOd7.WNeAbcC/XS^7
\.OYafK(8_;5,/#AW#B&BKRT?1#L?T&A?;2\fXEPb3.2L[5]E=U)U9U+.=(ZQGEf
9AFdB@5SLa(7=8U@)+XL2IEI-aR&KMA],J<dfM)4E//W5W:WYWD\\R]=Ag.UgAS.
DFC8JDFOK:-C;[8L\e#7VDTM=N(B21_MF<f>+3]cMd>OGg;I5PbQN8_Mg=_\7:XL
S(.IUOE\6^D-ZL)2>8=:b1L[\8c:R<Q(;8B?bEg:XI+[90?DZ:.[,FEb.BSM)G_U
[7[cEKOV,=L7X<P)#7d^eUfG3SB9.-FWY>PO\XQ.H-R]46;M^&M?QUSI6(:/PD&4
V=[=W88MKcQ6^NC,+eM9KJ2ZLEH/[&>HIPe#O;ARE]@UT;POQSX+6[b)?O.C=d=O
1-4F>)EYP53-)XVd?e+OAgP-W&375_/27&]gXC?Id4@1CMaQ<eVX_^F+1<^+Q@Q(
?:PBe_&G\QW^?B][56)&_O/PeT^.3S7>PE64IDT5aDLR-#e4APSJ(]ZW2[BMK]aV
;]BBBWMN#OF@-Ie=V:EJ?)c]O(LHKf-?8+K#PLBC8LW3L#KW7b,D8=Q-U8.ACd,a
.[E4J.:7VZ+JAaKR08S@&b3&^YM)(EEN7PO=M5.R_,4+M\].HMa+UO>P90[G2?dD
6D-K;cL\R[,^@IaMK7D_6&1#Z+KW(?Da8-B3D@U/K9_)BULcA>\+<BVbE9L>X238
bY(.[QXXTXBRU:/5;Y4+);U4BY;8Ad+X4QTB2fDY//:(;XbEfcSC--JX_P;Z-KGF
dY&<0,)OBQc1ZKI4M@?g<SeW8(7acRSfbI:2C[.\XS\fcESF5_AS5F4cA;/[Hd=c
M@.Z/g18NGZ+98GWg3SG<\W0YOLDY6WTVQ.c4eEeH[8NAB;0U/@[#ASaQN^W>DUR
)=@faYBS0\-L,4GE4eZ@ORO[Lg5&(^NXGBB=Eg,67Ub:(RgI,9fFCP\H4JDgAdce
FW>MbH;7FC7(8#HgE9S<\bc]M=L9+#IBIYRY1JWJD:D\Qa]S@8KCEX0Q6J=c>L5U
9dNN6+\TUb0O],]A=Z:a1EIA<L6b<IaA7AGIg2Kc&_.6W.\]JaZf9YGQK1RcUebB
1<_3J,G.[P=R<MeM4#<F(B\=9c)L_Z:\5YXIf<FUL^01E#V&c7VEg5MIT;AIZ5O+
e[dAM=P>\3KBD/&?eC#ALGMF_<#VMcA>Y?Y;F4.8eP^NF>8@V17G:SU\aQf.#P)(
Y00Tc]a4e)ea0OQg#WXe2RP[8A<=:[3J04;<XP:HV[?=B,4-#37A/CIQ[&?2S8Uc
Y9I@\A_e7A/>FC[6OS4+1D/dR-)?E@I7FFW#LB?P19EV^ea\CD?[NZg\7R:-;J;K
J62a#Y^81@:d09)bcc8F7FT#]9O=W7SQ&D11AB1b9:8M(RIZ^\JPMGLX7Q&CaMXg
b;?(^e=Y&1(I;aD;+;5dD^Z6cFD>H[@0LC[49db=ea)-5>JBgag1#RD=b9P=g81V
WV.]A3LSRe.NeC+#&dbM[2.QF4E)KcYG2[:6g@WDWI_d6XS+B\+C;a/Q]-dOGM.I
dBX_HS77OZeH;QT@CTT,D/P&YP^V-]+\_?T?R>5b[ULW/dKO,NbS/:a=Ca0^75>;
^KK5^PD\5=62Fb;<U@?ZO]Sd8JNM-9V<<1(fN&T-:87[dCGI05Q=3]9@Z=VGEV#/
Lb&5^<C>QYNOa7K#;]9-8X\7NaLYS+^6bZV0D-Q-DQ2BH8E8MVH/,G#.9I=#/_c^
JAR,OJae8ZW^_R<0WVA1-H-:2H?&bIDHZ:J,S?E3=,O6B@2QgLW9:VQ&f),&0]YQ
QXa3(NCSdeB&ETE-YE5KAS-D#N4P3UH9K8g0544J98=+9e:YV^[0ITD)aKSbKC[O
fZWeaOLH?T8G5QFN<XYQ(Y,:BgYL:M1[a>;_A0gM\6,aJNABD51/5B4OU?74=EO>
68F7OB]H^U,WJX,>cbJbegG?^M2Z_[1J69CF,eXD<QZg>;Qc#:>VHdPa5^]gbLN.
E-8:Z;0D6,#/L\fF5GDB1UcP,eI4D_a^019&6V@TB6Z=CQ>HdNT>1],V2b^3d(If
<?0AOXS_<8Nd)_O-4^TD@>KV;Y9e6KC3/XZ3CP#E\+&RSY=W(+2\CBfI[\c^30V\
FMgURFEN)REU?J?W&f.)@XK+g=K:)85QI>ELKOV&.(V8>dKE&VPVT7@7\64#BAJ.
Hd0/(gAJR<VS_//1)3Kf^8[Qd#C=CFXf->64]QSD&=)Te0aIW+DV\\6ab_=4eN69
B[I>TX]UN50+8d&DfMa-Ucc\VJ0PP26g<I<<FN@SABR2XZe+/7gJ&bdF^L8ZIA8E
Ff=(6.>+VQIK@XD8^fM>#CBCN,eQOWX2]:C]^\0c&b=#?6a(.58fJ8[X57c/,d1Q
R=7IGKT3&S;,&>GFa/PD\X^V9J+9;#Y9FO+1&YW11^&UX@f<<TaX6_DS1.8=Z-9=
:8(\:O4#C[KR94>SKE[4NK?,K7,/,L&8H/Za0HeK(YRW]0:LUY#3>Q^@12aQ11O0
U3.S<_6]XY8:egJ\P5T;\@d@RIAP85(>I)=7((<T^5#@/<>IJIReOP550]ZJcL7K
6<WZRE@).J\f0[^W2eP@L83dI2<F4dDBEgK&EZL6^4+M&K&)RBQW]_2(M)GINc3:
\?)P.K4;1D^\94GQ/Q_N^M2KR-VN&6BNeg>L5C2J?34B^EAXITK0@/0]]>L:U</[
<K6e3G:S(^;)9><d\C;5?(W7&68bJf_(9EODPNX<A,?\0TRObUNDeV.FYW405^Ad
-H]69OX-4QRJ/aMV]87/0(95b<]KV>AT#)6Q/aA>@#B<>,6dc,ES&,K,\G)Za9XS
QTP3_F,,JY22.>/9>>;[M5^B:#61dC<A8R;(Z>Pg<TF(HNXZ1LS1eA=E.ST1;)Eg
K=a907;#:^HVKM^S-]S5BIZLgB(P]CUN5b?UDFXc3MUWK\Ba&a5S5>]]BgNb5N(@
W9NaXPS#+NCfP;9b-3BF99WLI5T6\8I8>XL(3EaZ=)1<6(/L5;8K7O(OB=2+NNWJ
F#d]<W#+;,3>-QDHUc8AGLGI>_?,G-dgOHTW04H],TaG6_CbIc2Kc@0]NYVc?+g6
dHVCY3E5T,QG9J_bSQEabN3.KZ^N+9<a.XWVbTg=AK<cWI+8XSb]SM+_(^BMGcK/
+d@LLZM6?7H+?R[&I=]I.1XH/N#^Z[&b@VFPPDG^<Ked_:0QP@0?bg>fLQIZKV#O
:;?aVCF#5@dD=8HQ&S]>Wa#<9HfBcd]AEN9dC=PK97aV2.8V99a/Bc;^]]f+..;@
>8./Ia\)3fI+:RO<\[6GO,(:1_TH[Af?Z/UTRCa?(B6]F=R7[A.1>a3FFBb8fV(D
KD,acH2<I@[10#5W8?KF7TV0K^\Z.MFC7g<TZ(f]bV#,B=c7ZL@,gUTCIG4SRX-,
?1C(_L4Q9(5V:SLA;4KXR[D@@.V_T:&_SY[:G9VI50g7KW?<)EF+9CY9_cXSE0aJ
4@M#S^3c>-+a13fU[Qae3=Q4RNQAc1;_bP(fIJH:d^[BL[@2-eWF[3LWU(_#ZSRA
>.SIOTZ],/GR9+g3155.cd\b\TcAA86?8f)B7<IMMcLP\Of:.2bAeX_ELSDeVDba
g=HZaZP/?2LY57J+SBbI>NMTHc1_:e(2<]Y8eI(N#HZ1<=N@c0QIZ8^P4?dN5_O;
Y@d;N[T85(M2=_:L7Ja0NV=-IJ1@EKCKKd3#IeLAg=<&1fQgZKbCF_[c(I^^e,fJ
&3VaEGAQ3V/AELdMa_>L?]&d\:N&J1@e&=U;<QJ4)Og9@QGS-EQI8^#N<Hd;<I05
^(_O.T4NE9F1(ZKb?Y^,LTN0d1:#b0T]&KP9]<]65Q^3#/3I(^F?7bC-GUgE,7,(
^2ZA^+[31(E__;;WR8Cd-G6+<HC6ZDWG=1D4,FY9]/.XZaRfC-,LFA.F+@L&5>bb
OO6a?7b;#bIKTc_9NB.OPLCC-=O8U^C3bH,Tf3O;<P:7-0cURW3H7AQ1K#X[,Cbb
0/5e3S#Gg4=dd/M4f#J(_Y58N7N>6^9E<,Od8G-fJMF+TUT=E2K_HcHceDJ_QgX&
3B?Ia70>[&C7=F8Y:&a^eYL+P>=./OGSYYHN@_IN6S>R8cN>FTeIX[H,09L7O18R
:+9C=CSd<HLd]XdPY64^1a[2(>dUQ+cJb&O7>X-GbM2dQ:3@:WXQ94L=VeE=7QAP
<5fc&EU8XMNH^:gE6X6#,c^C4[]5O#+3:](TJ+Z5HU+Fa=+]RZK-LDf=?ZDC]B&f
Q6FbO7+(F0@[6BM-IKf(SeA54-NB?FGIaWX?WZE03@U134e^L=.c;+?JFa\e[TP:
(5YT(7aYfHK+d:da&X&TTCaM;&24[f7DBE3[GWTL2UMW=0P_,H_@3;a)bOEO3Z7V
.c,5S#MZG6#N=PPA>4=CWWL#9egH>P^6a.:0DWJ-/MK8TZG.FJIXO55ODI&c67W/
_=a)RU886]N+;U,LbFDaFYY:K?S-_T)d78Z:R_34W,?R3@8-^bX?e>GdfGZ\VcP3
<K3Q9AV\^3dSCS=1)J1-G3c8G7VCFP:SEHZ;J:HU=ET+?+K1XCJ3NJZH3DSCb,]A
BT8/a2O6E9fWFB1+4Q,eCTbg/JVSLI)<+M86ZADHA@<:7:eMI^I8.3AB\.0T0=f+
P=-+D=g7bF(<L,fAR_B+J(6AJbE?F9(2c-X.2^TLUYPQHZ^,e6-<^4-6\L025[<c
KO7.4f:cQ3gRKG\@S_K[^QP,fc(LI2Fe.([.DXODGX#\?Da4?4g_9SE2ZL)7_)?W
L^<eRFW\+;:c>=:48+dIY,\KS/>7<C2IQ+3-YTX67c;YZ<_N](.CTOEC+8F9&6=D
86?N5)M_d2/I0M3B)UMAIMQ&VW]0#?V^V.958+E7=X.Z7)=-U>\+\g4H^Z/:N_@?
/2[(V+[IEgB\Y+3?N(3DeEFGM^I4b(KCS5N3RgBL)_^7SF56.V.G?[+[GL./93&,
J/I\A,,72P:VQ&U12=<g8a2RdUX/SVM@113@(>SUOc9C&dGK/c^1eN53JSV(c4IJ
6/1fE(DK1)3IIJ)UF01a,]IA&EBT?S_Q3E+VZK=KO<)]\WU,.3a?AZ:L@CfVXSMe
MA32;JW^MaQZ<U4J[,3<cU+)7LNV^NQZ#]gc@c=Wd?b?9V\A65)OO2VO6TCV#S^O
^/=.Yc-XRQ.(eYD89Z\PJB??GIaf,>OSJBagJS<_&]P(7P7&)g5=WGKc?H.W7XYG
3g<)1D=1R;K6.d1XHBZe^<2/ZMS(OPUO3R+^(NV-cS^/BJ10S?G4^W.d<BAT)O1c
#YCRN2^#^G:b\28HE04a?QbOg-9HS8I<R^d8\7)HVV:1+0?dg^gO35[,cd(e;eF(
F?>OaL,2OR-Da=(8T=6(>S\35PGN)C9e339KVI6+WgL@\g[&WG\//X#E>cGa\PTa
TN>]]@DO-F)EN:_b#WaOUGNg_OU4[R)Z>8?,RaQX1MZG\<TcEIZb4,2g]g/aQ\Y^
MH[eI4g9?87DNe8.=]^)dg00?6]B/_.YNd.;3+/3TC3ZJ4D0)eW:5[)OC=+:AK1T
/GDJR3g?R3C1E([cE-E=fT/<-UW;aNI3DX7J>P(Je0C#(#F_^;[T\C.D]6fe<(R(
&e2T_B-4a;H)6]QGa&7DE#G@5cPFH#MH7DFQO5(;#Q,S_X:^_:H#<4<gOJ-GQ.4;
;,cT7AcR3U\e<#R6V<;b3HP42&_ZU3^(#Y.O.e6BFG:V#Ree>@5/P)MaNeL80#7.
GA.(]?Y=YB+]83YR4R/,T,#MOaU2b6cQ/0J413P4A<\RPV4BeN;eU1M3.eW9dbL9
Yg:FWXRQ=DbKbcg96#]B]&efAcEU:X/9X18E>aKbL<:/RK7.7-)0PYUZ]-B-.f9?
+S-S:_G^=c=,dN6];H8(X>\U+MeHY7Zb=G9@?_[Y3.3C9bd5FSg\5KcZONJX(=-D
+^cTSQc(d69]3P[I=\=F&Df;XW@U+3ESF-:<VZ:T<LGC0F0J;7^9H2PF(=dN3cg:
-1\UZEa-HWAAF?@D5U<8L-OHM]e4IePN6-gf4T:B7N+SGYE;Ye_d@VEKMgb^UD:[
G(::SUMH)P##a)S<0_XNTZ<PY;Z^>aEQ^F2:&=X&3#Ygf8fG#QWM^0^PM)2#.7C-
FJMH_Q[=^U3fR[O:>V+&0@[9^3+,>T.(\.C>.P]MB19QDS7G58R7^J-1-RM+?Q#[
JV6/&E+X]\FI&HG#/<)1J2,M>N)A(@eC[H=>bW^dN1@#JaNOA,eRCeJI]9:^CVW5
K:4\>OQG[SVI)OX<eDF<a79HA=1R(,P_TR+IE-QTf/XH3a(Sa0XK?)[)EMD[GKKD
e8K<TFb>-L3AF?&NOOLg-7H[^B4Oe(=#VG.c:6R>8/PPGM57ID\JGaKc)bM_g-fJ
;B2#6IcGNU[:Ad\a^dFJOIGC>?+2FN.UA\J/?(+-Wg[KBXMWEI5[)Z)CYgBDI6RG
FbVage#_?2JQ&T:fa3e#YP-4<930J4N\0I2-,C8Q1\FO(e7eHB=?8/g?1Z8I9S^#
ObKKG6BV)<VF,aR5HfCXH77UP[;4&e-.KJdWGC9>0(O<NOGdgH1&VMJGDe;TVBY;
[>L4PI5&,:?],af=5+?PG7]6]R;:.5&(S<M=Ca0UE)JST_c/<0E(D)D8ZHF_XA.&
9@ga>KV2Od52S_O+MB?>]R<RY+DDUI=\ZMP;)<CE<Ib.L>R8E]:1OI[Sg_].Qg>2
T_gRB;WH9_b:^R@48]c4>[WfJ(#=VOPZ69_>4\-f0_L>,HY[R-NJf7XZaRI,#TK9
V#E-H?-F8HU)N;2\8RY5CaRdG=NKeFbgL7=OBe&\U)S0,#7)[R[g<S5d3Z(81KZ(
,7T)3^(91MASXE.M_;73K040+@V/5beCM\HBdPdU(Pb9(N)d=98A3J-42Lc_KSa^
AMF0,H(+-VTCe,>IF8WY8UZTUC8U,#RG<0Sf<\&]F^DbEGI@-66NZ;d9-a<]^9>V
9V54DLXH3N=+Ya.4NOEM->(,UL+-:aPJ)GK@N3HFZQ6ET,SXg[EDJM?K=UgY/7/c
R:(:f)9?_YUK2QS[NR7cV#(,31@cHI7R1V<K/NS(X/g3-Q]H^We?QQ:V<U::G9V<
95a(9f#g2fFZ]7,&ST/E72WWBdP_)e,?34M3Y@g[JPNGX0_EJ8I.8],8_T_/@T?5
M?OPYFUH_a0/K8^/.,c8/:HCQ5WZV2C&9RNBE:_838a(\9MV[>B:P3;N/_MC1\C,
AVT=;QI+8)_dU^69?NBA[T#B8^R#EgUD?G&+:B&b_E8</5]c2-H0,PD+MJ[.U=X&
Kd>;6?&8NCEO1ea,ML,,5@I>8R_0<_F78C(A:_KeL;K3>?fWGT/HabW-bd&_GR>Y
NK8>ZP)0L0.R<<V,M#_d1V+(:YD4H[RHLaOPZS52V_TF-^X<FdO_H)SAV>B5Je95
S6@gV(/3Wg)7W+bR]Z-)YWLAa-KbL1-ZJ7,775@GfM5_JfQB=)^@#6VH]2cd3R7c
_ULc,9#T2L+)A\6YC>^:7XC/dHACC?U<WJ;N\Sg#21TUK(W9?d81N<<+_eR7]5#_
IE,dDPPf<KWR>PXLg4Sa/Kcb=U4#548bN\3]N]03HEeVW>KO6??]Y=7CdTS9&CVS
C4X=6LL_<?+f+[b<AP#P-RBSfQUFJE[C35^EK,Ub)9<71Q\QAgEUDd-/a^EA8\(0
^1=MKddNL5OGYEKgD42?KT-Ff/B?QeVLZ?^3Ne2KXF@S3cNI]+:H(-KB4Qa-M21-
\:SK?fcWdE@=O/T6D,60ELP;[fLGYUNDe8=BX/+T@OYJQ-[)3;,<g[O5=Bdf,BO+
RV^WfD68;>IWVbQ,B2PQ.FC.9VaQ,3eW[]2@PKdO#=OfY59MaK@RV;O<fM&:@D.\
BgHI\26FcdR:fGfbeWW90KU]B^[(TKR63aP\Jf-5:3UX_W:39-@O/1G=L.Md@0&2
4\B3CfM9]G5BaO[68GIN4XDXN7eQN^4[Ob708B]BaR[G-#-9.fU(a=,cN\BFQ7Y<
,T.IZO;IS4FdAZDf?[.0XWXMNO]OUV>3S6ERa1[+=PfZ+MD;#]Y&)YGZ./;FBf7I
g^f<\G_&H\=G;0?NGI?O;2I,&&(GQB[E\-.LHFHdO#Y>1<g(F0/RW#QF6<Tc:cUa
)Q=NP^8X#\2.5+d5[?I8_&7NG.\:1U6^f4gI]#?1(HC/REb4fDK-Z,B\].Nd+R^,
<G,T/?]G@^\@Ieb4=F86WFdJ2]-2a8GK?\eVVBA=4a79e&FIgZ^SA#B(41UUGITP
I9(dF-]9GSBY8dL/M9f48>X-[\^CbQU=caK(N?5(H<5?,Z_YJODT04fIAf-ABOcT
V9LSNSI=Z9AFgYK(4-I/WJLFfZQ1fX6C>2R(8dGS.,.be2#FGWE-XHP9::H)=Ua_
I2a9+d9)&JXQ:D6]#I\,RNYDL<;A8GNWXaD,+XJ;<EJdSW:<c02#W7Y^)-e8LBRf
?3R.:g5A1SFS;ZeM@(AfQ^?fWR2.gY;+4d/MQTS+7LQJG78.95-99X=QgYT4F9GI
cKJ3BA9R/?1g+&FS@V\cJ^bB@5=<+QT<;OTLE<O28]HKZ6Ue.X6D=-Gaf0Cc>S.^
PHXY7PS@_f2CPAcG5\d^Nb[:86/UP?B7_,W.ULX\T&XMf-T>[1c6[2VUQ-ARULZ[
ReNYZfDJadG&=9SL1DGV9G[O@]_dR#1.PB:&WP4:dX1B<D4.e01M,K3URT?BKFR0
H03aD9VDg,f5PQ[&FNM[4#fH]]D7A],O^QCQ&P,H&+P#C57FdF.C^b,,#?F&NPTC
GfWE7#]25Z.J?HYCPcJUJJL:_BGVF\R96DfA@bK5?,aN[,eWZ/9F]YZS05_f[WP;
0E6I/22,^(gGID5ONa0Kg1-[)7J-/[X7dTW9EEU4>L>AU0A:b2^>LT__C>QE#6ZP
EgTbRCaH-3N0))0L;H1gC[H&T@G(1L2YQTL<^83^LfeK#HPRJ6T5<cMQOdg&#&U^
eD3F5X4Y@L#D09A3#Y595:e9]E3^H_F)PJ-:W2g(EXPee4^0A_#CO2(a-8\;3c#_
6F4#=@)<d;edMZYcCO8=BE+O_,aa:<(WGC5F6c#PRN5\9RVV2g^^QO@4AE7E:M\W
;XM&g4Qd(5K^_(Kac][#B@,7D:S=Ia9YMZ(6e:;,6BSR94a+Yc0BfQ;e(7Vd5R3[
d1fV+^S)6\+KO>I0J;52cLTGK-fAB#HRAWSZWNFLR<T_@]B]O=^;fc\6J5\#]#-7
Uc5=H564[4:\V#O&fKOO1BB#NBYT?3^eg79(HZ29GfZFQ.@Z/5WTB/dF)5,Ffe-/
4+RYPacZUUSg,?8Wd_bP7R9M[^RYENJf0bHX@f<d:Tf1NOGE@2>U-K:6PKGNDWaU
^Y5O/^4.e&3)Qb7XgK.2Tc/W32f/f0AAH\_1?gV4.UJRXMK7S3^UKFT)66O-2P8U
]YZRXT)#(bDQ]aK)+-B5C@2_5g4F/&g9&b9aN>[>T?IRbe9:U0+];9V5N_<b-aK5
MF-]=D7ZNeR;]:M\Yf&RRS+A>Ce>F\ZB/@>U8-E-)3PYEO1)-RDfJN-.a;FXcMR8
T:K(^IaaDD_)HEYcVG[\\14_-X=:A_RM@gLU.)5AJ)g]R-/X@?N2V6>ZC(cW=HGg
VRVfL-B\&5L4=8.]M7MR&INO?=&8c<50>+g8(49O6#K8?B?,,(89[O5OK>6[#&<M
Y^O^B&N9?HMT<G<_4PeIAM^HG/K2ED8gZL;Q8Bc4Y.4V;]+MggWEV(RA^C(1gW&F
c\@Z\LYf&,@KX2L;YR+2TF;T#_B.B9TPI/]RGWSY>AVIK9VQ\G<;>41/#UE;JdOS
(bW1..ZAG;g]^Y>58VA1BPdWc>gYTO^28U-#]E)(GD,(Q:0)3B?EP[D)&TVPbcLG
1;/#:U^KBVacb292S+G0&?E\:F0O(EM9LgU\@3R_+4]6b-M=@B[Z\T.CH4A:9T:L
5.20GW?\YVCS8>c7f61O7Y7<SeW-ZTIXI@eN,([aM@:)#+Abe]WJE1HB<-^K(D4W
HW,=ZfIQcR32<QMVaS6DNFPSGAdE.QL:,VMZ\ERJL3FSN8Q\Y3c9\RUGee9g24B7
=1WBF5C_[F5GDOL?:Qb45-@NW-Ec(d?2@gN+46b5LM6(ba7aDWC:4U7,d7..WP#[
8H[SHd_5bK3[bUKd2Gd]WW^;Nd8La9(_e^,c6LLZ1)LS(U_1IVP&Y239H1R)]+4K
/B8M/]=BH5^XRTaW]#4@Z@\]]Y&^.^8W5+N\8:LC95AM+4HT)SH(eL,UZ(M64EYN
Y/#cJ(LLcJ,Z0MNW-1f/6d5gI]OGbTR&7&.X0FS7J&Y+D0MCa+?Ha6&AQ++(CEB<
@CZ#X2+WOVdJf:LBNKT3[5MPa9eEe=#YeBK(>gb[5aL<E3THX_H(]1Nf0IIc2)/8
[T<?GY=Xg8UDPK9S7AYP&H[?@<D.baQ;6+dRdcI@>TJ(Y60ANEa#DLL(ZA==OA\<
<2?+J#:1eeGbg,Bf-P192_2RVNN\BKLOS+GL0@1CC+H^T=cI3K_Tc/XQAfFK&BJ#
C1A7CMUC34KD#J_S)<:Y&6)#SHFaPMKd7HX#b;NQaf<_PbBOSQ-I@eg5_QW7ZS)f
)EB2:<ZBB4gGfeC)?-V5?]cd)KP&b(:AMb&3,4bME#CVI1CNB[(T^bA(:?)1:A]8
LR;M,)K6J_.&>gWI[g9J<K_&]BKgKA7F9644L,DEgFNVZS^#BW]/>QH,<?8;6KF&
gS/@TPf8FaYYEK3-.O<Oe.0fFL==+FIg,YL:J?/Yd,>fgN9JEUT/dI.3A<_2XY^2
+?I)EaaW6^OON_4\P&:VV2)b(\)gbG?JW#PXC7)0[:KD>=()3.dKSBQZJ:U:?20L
.>d>EKO?XaG;W=#/OL>.?>UZ]5gMHOVDDHL?]eM/536QN+6XXb@)/4ME5E5N;9J7
0e^/PNLFQFBMX[UQ,d-]W9fZ3IU++gB[dV:6_>&U.8I5KA4]-1?aK_[PKE3T+/<E
3=<a=&-V^U1>fX^Z1g3:#@JGO>(VXFf1GE&B>DcLRDK5?4<V7[3::aE3Y3^;09,X
>IeP<bG4)(S2H8M(OeNL)_M3^B;69EbG]LHO+Ea/&MeN/IBR6/U;SeGeII.NB8g)
#MA-X9N=YF)EfB=XT4<4=AGg_NLCfd;]GB;E]2#/b?S\.fU@=+G<ACQ<:JSJ1WM4
WUKeKTX+[KX7IUW5V:C/<RZY3<=DcXZ.,Vd&?7=;Z-I@_09VGUE91Q?&@HIZbXY,
469<Lf3]?S+<-E\37[Qa80C+e<;71-P:9IK&.S,IIAd0CcQ>:LZ;R<4Fg9b4WYA)
X@#<#7E>0TFfL=3S/-BAAVaRDdgf6)&P)5&6((T.&03P=b,_+MF>]eZZL#(/GP(7
+GK;9KDec:K?60Q>6.#Qd=JN4RdE>L,?/bD&.OO+,PEO>NR[]]=B7@&]8R?L2_U)
V.O+EbN]+IZE/8#P1D>W^(21JX.DYW/8#V1.0TBM#(Hd9\]4/2^\BPFI-(TePENE
,W3\MDgODJ8/YcD(PW4[-+.f6fgSW0^//;\JHP?c<XC<g^b+d,5QEW2>;-S7?C><
Df]/3/^]fIFJYT#<\Xf-c7a,Y8+Ec=P]c..g)O65T=ZS7-H6=HAaFFP?J[VbNOT/
R.L:UTaRa[bYK[YNeY)8WIbX#-3;8OIff#1EHY0E@7B0M_ab\W[8_C89@(NRBba2
O6Se/G61-[\QdEaBYM-^/[),9@?JYgJ.M-)&M51PS6^#<ggP^M0#Q#,YD;_10,2c
=C#1cXBbTAH0I6KSgL:\HM->=VIfW\S)4UaAf#MG]N,[5;LNKKfBSdV+Ub1Mb0\-
NW.F/cN.@&]X\S\^M<J:-P1,L7NgA#+F,bYa]^U]7ZOKC08(D[_X4E0:18^>87>:
XSK;56c6.Q]RJC#PTV;:g=/DDJOee=dfC.J&UP\C>[>85D&M3GRTD6T1fK&F+G7Z
7>fOE-<U[(&Y9_13#U.7&1;/@M1g074/g^L-MQ4I86S-GH/cb[;;Lb6_F>&HSfRX
D-,XdN<.+V/80Jf)U>IcVN_?2^^XII9:#+)c1GO[:]<-<4?PQ9?(717X1_c.(20-
5V315@H9Bg)M&Caab(8AcB2&=bg\,U\X(XI0MNC/2Q7.5I/;#S?13;6E4P+O6R-_
,,OV<a&)./DBC02@ab8e2Sf#eHDFV-.c8ZT8(LY1IIg)S\79OY=Yg^2J,[:)TUV0
,^b8e4T[AL6P9S:e\7Af:GC5G<gVOO]8KcQ>00ND@8QQ>fAeLS4L.)a^fAWd]>9^
5?d1-U_>)/.UV7;Qd\MX^1I-:<O\b16MX;I;dSK/:LCACL[YN0Q_?b&.3Ib6XA)J
dO9c3F:AOc#^_^Mb8O:77e3[5K8X8&ZV?<Pa_f3.&:,IS<ZG:8ZV/,ZPI?=#ae8K
_AbI-M#I)TJ[BVfQO42GWU=eOA091]PB5]/2;;/9[8[ZebG?G,#M3V/,@aGSZ.P\
D\M[:MPD+.KO_Y.6I6<4,@JWa]Z2W0\1fB=@1#9AOE^GX-_14U/)0UTETH5]/H1]
#8EL)f5B=fC-d:^QCW[1X@Y2cD7Ab2AY]Od.f_>4)HFHKL+N5#T(&c_Z;0b>PeUd
ZFeI+5bJ;LOHJfZSMfQ/[QDOV;4dD7WVZB^76B<BWM>AY>:&F>+_76ZCXW.G&9Oa
F5>[N5JL<UR]9Ibg;5W=SK9@@(fGWRd[0_BP,O62?P50_Y_)OBP5gQZCN$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_MONITOR_UVM_SV


