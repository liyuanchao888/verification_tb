
/**
 * Abstract:  This file serve as a top-level test file, which just
 * pulls in the individual tests by including them.
 */
`include "ts.base_test.sv"
`include "ts.directed_test.sv"
`include "ts.random_wr_rd_test.sv"
`include "ts.amba_pv_test.sv"
`include "ts.override_test.sv"
