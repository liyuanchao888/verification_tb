
`ifndef GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV

/**
 *  Master monitor callback class contains the callback methods called by the
 *  master monitor component.
 */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_master_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_master_monitor_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_master_monitor_callback");
`endif

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
mxJnJMxy131qGuUbB6UZCbeZHiPysuP6Cr3ANH26Om8ew99nlakT5VclxE+p5ECV
HueisRMDRcvtKQY3pCxoIIhuZXAEDmZ9UErNUE74sYTS9wl0G4L8RdYfi4YLWX9V
75vCFcCQcNE8mNOG9CxLfhKJ2imYnQBzSroP3rZhPFk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8874      )
EMgE1mqgxIg4RoRpMRSc9oX9YfWm/rDfkb2roxeQ55cGzcdtx0EyBz+sWGv0niYy
t60IS4vrsPueU0By3+7CH3ZljP4IgIJ/jII7kR4ym6WIFTkdTbWq5U03W18l5oN+
NUC3bOBJ38/AcPl/7VZH3z5d9t5qm3igAXyFfjS44uOq0hf8zca7l/SXJejpbgc9
BMaXhyoiYMrhKLdr9nRTcE6wHQrRDq/xjGkWwUHgxZ6ZSMb6KS6pjzwVImMonjJL
X3nRhVg3llLpHehpX1xlJ81h7/gVyle9D4+DmkXHfPh11ECJxb52uNujpPNgn44V
rTYd9y4CIyOTzV7zWY7OTEue2dAdghidcz2WCObyO9G9ARYZaOWFJtj1VmRd9JEM
MJ/HSLNqxrkwe12ptHyHRrzUvnTgFbY9yYgySbH+KekvZZrQhrAciEH2aKSgkrdR
C5gF5QuK1xc7pHlVeZy/QI+DmcsOPRrxu0iJx2g5d279Ex0TAqNJAhmvpScSV5w4
Pq2HvCtnx355IoUrp/zuIexoxmQyDPKqXk7i7iYEiBzEBmB+r//fcIs90vhbTAfx
l/vHyOebOqP9RR8kfj4CJXX3ifJue/NgZq0zrIgbxTnfpiGsQOtL8djbLSQJ4bEj
33SM3w+VDxWcvADthIP3bEOGSnEdImQT4zWvMqdu7ElAnlg//v+W5tbDOX36kCZI
9wAsZujWFUVP1XRWmX+bZou4MQ2ArnVpLYPL/7mtdcRBebVe+XtKtlsp2uhM+af2
bQkq0yRJANO+G22iN/xH+CrGbMDk7VnRQx7sih1m39JL3UVwgQm2+N3fxhgHpE5G
7ycFGw+r/f1tRzc20OIzv7wGKudqpK2Q8TbHzbM3MNbREvOv9D/mH40aTjLDpnFW
9hNF+spWd6E/kxihkrMP/LcEnt4Db8VnDDxl9Q/9SeVbg7lGnZtH9chuZQwFKNir
AecXtU2bR+ZS42yT37KkGAap69fBYahaPFONyVEXhveFkOVKgyJi0vJ+MtTKPa5P
fgst4BN08+0CH0LaQqKrSuh2Vv1PF7TAYeSa9XAW/+gLpiimtR799IoQ4flNJXtK
IofuiIzGCuJhTm8Wsn8VnIW67fO31gBbFazNmuIYf3MrNStXzDCX//E36RP7v5BC
snmMYO1l9z2xrAXa+K+6qoKcRdUlIeXSCU64jibuDWX2ivF2x+/g8VbhwVtYIWOL
ov68ZNfA4pG91htj1tcl1FSWafrEtb2eRCDJ9RwOZAm48HGwbWSe84/03f26XKrd
9GAmPJ6Wqp7xmyRsdg4ukN+zOwz///5vOnJ6lOS5JxkdymsuIrYWAWLXwapvkfeu
pPpZiQFplMlTZmIaXXR6ZF6hR9swb8gqJhOj+ueY6QUjZ/EBJwwGqznyF3M7XcKC
2AYkvG3AsXibU1b9iwTpSbIx2g14Ozno/PxYaAJSwaBbsyWFQWW/WmVItG0tE+lb
eK7MxPFdENQ7fY1Vk/gpn6QtanCWB2QjI/ThgoyHZK13g5gJUZqyFYQCjXB7QAjF
6oQDodT1SYxpNyjeU3H1tILyDzZHCnRR5uNQkP1zwR5ZJI83lrmqJS0UBbtCAFaq
T19LZS8k5K0LbU+Jn2Wrlj5CXGhj7o3eCUdd3Q2v5N09mjFI78QbX2dsEpNVK6ES
2sHUdyqhanhlBWqz9pSBQE8Zl23RPmjOfkE1dJK7DBRD35z2uz6Tb+AHChrZpZd0
VNfAMbACjkq4I81W7jskXe+WkXJn1UMJphSD2dyjnc+09Ov6dnMgMHuDwfvTAP2v
SujNmma066dwiDwLRwSKM/6gWGe+z154asJmcgxhuSWLN6rgpO5R9GpqiTrRWSin
KbX5E3cYLKgBEDXPyk7r0/mNY+7VGJNK+jmD33Oeqr2E7gb1CNqLhHqwIQANZ60I
+QScEpjA8m0IWoeZU3RuZU2RqNd9cY+OanVp+ytTXjFjemVhKx+tcHAX6fTd2Uj6
/dtn6YOKdEO+maFDYGo1/P2yplCDVDA6B9OIqzFVqbauhjOBEOT8WYoYhUkzEvGF
d3mbWNUvFr7pJJGkYWgL8rKd9g2hgWPvX4Ph37NMHmmCaZwyW3TC8HquSt6RHgCU
FanavH/33W2gpZgqSyl1+79jeBdupQqlUiEjsn4zljBWulmCgsirgfM9WGsR6Ic/
nG49bG+zfzmNpKXLhDEmUxRV/c722+SP7rK7mCkuPpnEnQnBDYAl750olx4LCRcB
Cra1cjGIDhHeqHNjYad0oyqAPKdN+ZWi2iWxHTILbGnaGqHtw5hPQbafxK00vq4c
ymCJsjDvhLkay/oj9UHF4cfmKd/Gev3TwhYLCIYWTxqud1kWsWDwrXLzvP4ymrFX
WDSUvzh0084149Y+RyWWJyqMkrYh80N+j0Ri8SI/I+7nQ7pvyDxdLuvTzIaeqPgW
uKcD5/ieMXKo+8GF3XYWH+q7LJQDgASGdOAd91p7eaBfLsbwEv7h7HAdHkzJ74Gu
0Dcq3l/vkUVaKDR63gn+7/d8tVcR9BqLKBE2jsry3Q1FMXD/b6yu1SBHw4h2lAKa
al3+CXFvfpPtwnrCHIbkZf0hwsIt5Go9v0nXukeB5urf2oTkN8V7wkV2Vhca4u6p
gyXVj2jJyK4aM3qlwsaNpBEEcF1xPliLso5GE4rfQSQeeMgokvBNi+0C14ufNCHt
8DVcwy+7N5TJmGW4wSX86JpGv0Bea5BydOZjlft/Y8JlBeuygLpopJLJXL/BGPO8
T8mV2dVWTBsYzfCH3TKbLFI87Y349AYz+H/TcTKYeYS6U15VAfwWfckZhjV/ICF1
mENB6jSW2bPGjqsvO/r6InK/ebslFfDLopXvtEcct5CtKtZN/dcY/lEyPFV7MVdP
wImEIM0x16yktDUyRy36dUn+ks4IkFPMLI77eFm94zAMPnl7REkdnIusau7kerf3
pwciwnpPJ2MYqbZO+PwIsw5yFj/EIUXHHqJY9PDMUoha3LGZA/knE2uqY50YOKcd
liVw7h/2hQVJEZloG3I5rPCjveFS4Fb00doDHq6JJvwfcQ9eiRlGfusWYuvqhlpK
dvo6fttdCMdFvhQ4WCH500rp9u66uTmROYhBeH4zc5biKCXIpzv2TOozkQnS/ZY3
gjzpe92zeA7lFlKrlufkEJnOEG98Q/8/kQwoMdYXMP3073kQ/Z0OwpaLz7t59DcQ
OXnTlfsB5GPmiHa6ZTCcjlYGCwulzejNGwGucoyccO3i777VGYgSHodjt/MSsEW1
r3zbPrT2kRSzz02ACuyMH/M93HM7YreJzSLHGxoGvdvx6W1vw7TmO00JsPQTGzd8
dQrgrx5MHyPhEKXZ/Y/fy/BcHBy8D9Stfz7utA1lz89soA0Qt5MmNG8FR/0tDd3R
pv4ujwPg/1LP6C1YkkUJBp4LgSegACuRKAYaZMZzOd0zDBgH35DEXO6eWBv3+BDr
yQAIS3qGFh2pjHORSqYV6EKcuPutalhBEjQ4MrJj4tIse59JoQ6/Xc+KyvB5wYov
AEVF71cMbir+anxwHs6FN6BNMDCpik2xvc33bgmtQIOkExKP8UTKh76qpRkmR7jL
Vp2vNGtWq159dQNzCh95+IkrkYO6bG2sWkSscssCHt7KqDmFxZo2I2bO1MF3NH1R
p3BPOY2K3Ey6w0vUSZm/s0YKCryHx9F+cOerChsDg0Ng/utoulq6CWD6ezepImyY
n1jJcVoJ1Xcbh0o+9GBFa//bBEql/wu8yZoZ/rxi713MU6i8YpqvUumQmtMKOnGF
hKjHy65yEnPDAPYjSz3Cs7tri8rFHmnMhowiMBv5tC3XUUjPZQfta/L3ESeS1XiU
J6gbcAyzI9/WiCrRRat/gwnsN7c2id5UyGQPeagpIF9peXerzezgpChxwjGNImdp
LKpWOHrrlG4QtI2RaJtWDFu6JzbBRu6I1c4Zjh1vV6X8YZk4tj6VSyAGg/YzKfRR
a/KUVwmJ1CqmSPQ9Xa5rqQMEVwXzVMujE5roQFHamILMUS+GeMX/OSp8Sb453mC2
p27hEQZzC6WUg5e1CpXRzFYrvbrcTnINEPdzKg70guNHr00IVeTHuJ45LpOIYSZV
f6BMudxxJX6dcv8P9bLA/WIpoely0zdhm3b4fXq7Yz8Y4kgDgobhRq01GtUQDIoW
L5TRzYHpK8B7xOj8M4pIN89yOv5aBg2/1pwiv/4DflCP3ny1H7lX/vauNoIzibWm
yQm7gzLJxsTRHglMrXEgtX9Wdth5FZ0Sma83ydd/m1wzcM8LAbDoiTlMUBPlEFIN
H/QEmcySrfMYYVRb49JjjJ2u17aHfUPar5fmfrae+lOD9hxoBvQjJO4IjQ7XP41n
gMyeC0QRjML1n04ZqSoz7s41MrxxiHJyve3Up+eZEQJn0vclRfHNF7cfymUH/5Vc
lJM+TYZpe5Oz690bNzh+oNeni2ugKZb+kLDYfUyLLI94ig3ajnOp/jWOWGm7zYix
dXf0vnViSYAgc6MFn1lETsjv5aW28OA0vSOWogVKVzHrYXYLL/+b+XVBXAhFq/09
WE/C6uRFHEvTcRwG0WsYRgjSTPNd/5ZKjyuoyot0nWYKcpKQokxDa7KhgRBLMKw5
VdyLYxMUQGkD601GEbVQfx3CQ/MQb0bCgTBnlldl1OmSYVu0fCmZ9a21wA1x/SHO
rZbC4CegD3TN773gu20eZpjHFiZZaTBNgTiAgBp/DRaSYAt3SJI9gkyfIeiXfJbo
/r52YdPAcz9klELU7O0iE4ZefItnJ/NbUYCO7n4vvM0nsNxaStr49ngwwdH5GFC8
fAvd/0TyfROaiX1QSrpP9MmIQiEUSlbFq19682JSUwh3/qT5QduLR7V9qW/ipx0Q
FIf4ukHGXLsPmbH2mGmBfSLQBz/LjGES/Vf69E+bFk+52zdtYV9Quj173MahBEWs
sdNzkBM8UTSY0kDf79O2cjjhcjxcW00uAlkebDV92jzgDh06By7LR3o3IuzReYBM
bZpSDUcIV+VYuKLrSxXKfai33zDXlNFPjvRwA7CYMpniVN6dtFnQNL73rdtjRovQ
cu8SoF2HR6t984m9gNMIZVDilE2Ue05tHS/ykenzrw9hbKocsrQQpv3vpLkwVOBN
osEuG8TtgefeM6U1yxez4bRyr5X39WShXwO4IPIJfNl8TBLUuFZPdZ25jpHBjkWe
7qY77rB+E15qtz6ziMGa5ZDyxZQFcaedkt2lwDQpkCmH2ltcCVWgPgOvpRcDWNAj
VRPJhkw5P8OPfwS5kdb7mmFA6/8R7Ym5y1lU5ljGxanDql+xFK3qCfdcuJbPvYIZ
pFRXka1Xe9o2K8k2xMUQBE95vGiSObTCajhBq2NhqYhvU7J/ddWd/gyHeehPPll0
+qc4jCJ+ky3IWW1cBwDy9xPBEaFDXbMkPQzZh4mgADnJeeoMml3j0Cstz9IARs8V
1O6igU/OddYZ2cslCq8EBPsd/XqdHFxu6VcEkKL4770BkFgNq4DiqfF/Dg2d9oY2
uT3FUDlW7WzO+zIFxnvtke+A14/1j2rtyq05LGiIOiILFfEuYHme9lvH8qFlbkp/
J2nCvXJMMNDWLPNc2SYSyP/l8bMEMHcWDJaz1+iPJ+fWFJvc21ddMsZ37Q+9HBYs
BDxPcngRAQoIurfEhy+Van23cYYwlllH/oG/AXvo2Gum5yEIKJyuN1xXqDHEIQP/
wAF/jFccGYv/VFrdUKloY+S1TCIuyilRnqIijmOp9g7MdRcySQB404b4OiBvO4JZ
qfV4C359s74t1gE6NFO2LQnc9lKIzKlv6afjnBI9WRZl8N1OJ8xht9iAdi+oNtv8
ISc63X9BbKIU/Uy9ZOzhV55Y/OYmfxLbbRs+WIX+mE2QdYA8KtRxEFUvhBw3z3k7
61Iczg2khJyyvwa09hBFCayPLyW51zamza3fqG1Jgk+o8gNiMNt/seSpskp5Ynta
vKlcE4zBMAW0MehHChmExnMFLHYjbswHLISrHct4AsajBkjPkWTu9htq2kFo9W0v
rmd0SIUrFzAChejuH0NHC9rEbrVmECdF7xuOBJSCgsWlC8pS1vpHV5AKZWlVUdDy
acZAtR0XAONH0HI0/SLlq9PCc+PdrPaeWmXI05JdTIfHp1HGex0lFDOMgDoOzKQS
MmyX6yZBC9ncmHTCthdFQ2GhBb56mr0eV8+OgzS2UlB86VgQelA5Olbl6Eqgi+af
fShysUoDT2s86pMpNyIU1lHbBxZPdi3Aztcw/d8ZwfdmeGkllXxdW9N8ZKAKGFJq
N0ct8CZagEHW+WVGPQtylDZKCbvxfZFzgbRBqeII2b/+ZW8+psJij5DnPGOKTDW6
PKELkX1XftUyuE8HzpsgQg1K1ZA5OU58EKok+LhhLg4hW9DtchHSoESOVoSMa51S
IWLv3Q+ju4NF0qt4lAGzl5UmzC9Uj5aSc2tG397RsS3ABZ9T4DLpK6nn8QOH3JR+
XOBF5F2qK/fQpHuPXLrUFjCY4jyIyltamXBnJ31unL1IXO04nvL+fHpBzV4walZJ
h1cOTAVjR93QeRSPvuoGnfw5If7tGZcb1SnF1z5eW/DOpF+citcj9+E+fRilmSJa
28Z8gI6pka67jnGB5HXOBgIfI2mi54arnk6Iy4XEeP4uKJ/kMQ0QMnuXB72AbI5z
C1L7PONJzzIIsLjsK/hwJHX09jG+oIcZq8gAlPuxvQQb2zQsFtDuHRYKOXvyFv2V
noYiRCusbbjVE7jqs7Gld/Y3rUE0or6HzlOARPz4BOuwyc4T4TavAXx81DApKPkX
CsaBJXItG8+n8zXtrirVRNhTgxIYThsWE2N0sZXbYQllkz4L0u4ETqMz9kb7+UPL
eQAFfxmu5cqZw3jcumh5i4ZdxHhubn/owB3RzhQjqvrkYCPFHtqrEQhY1NoxSVk1
H6IH8/WnAIEccVBxfYQmZGBfioh5VuZHdLmWUroXcqQhIgsuXdt5gefZ28uErT0L
OSfH7Olg8ir9THNwog9WXv7z0MbwsSW0DwtjOba7ysa7kK2mU0UgYwvtv2894EY0
MpQeywHFZUmwJllgSZgnfjFDLdx2AVM1j8FENR4sgveYNyeOi9tXbB6XMbeHnO2g
MKQ/rBVeVufAW/FfuabwUQmekRj0jxlcwba8ekGbfguqJb5iPXnWT6u7MXLXu1Ay
I+9OXICfevOgPKE0TTiUvD23pTre+cm9mZ+uhkMeAbr1Pdf5VThCqJzyICiH9Vut
93Pje0JONFRZTVI2FYeiC7CslY8ESt21yAGt5ZuZbZL9qnUrUZIzVGm8n1puO65/
n4tVD/Aosu1YvIVi7xY6YprXBHlrRYQjf23PlTmRfYYtlbuUsav0gqJyIJ/1clwA
KJ8isYjuCoZougoeAFwIV+Q6oyE0dNhcwilfP/nOVeo9+B0+zrxkqdr2sfCY7rdh
jq43sROyTCRBXmDlwEouaeLssVdd1rHdKfBHwlwq4BYdDX7lKvEZHXznmSA8QvxA
e2Jr8OZDxbENvCMBryieaUc56b4jAimph4ZSUiSIXSNIlLWQ5s/xpJ0puKQpE6wz
bnpQy6m704OG76eVvzOjaLCzcCXm0OtrgnDKEhah2mdhnd+Lue1g/HWYN0hJlzwo
L1HmvZiyghjiBJH1WmPn+qdz7rJ0czEPF5U9KctjqVYz4b8a7Kvgjww7kegLvX7/
1B9gcwGIMEmpIUPvo4YkDKoNgZzrfFRAx2jMWS5dNptBCwsvmwd4ZVBcWpQCE8aP
CseI/6NxAoXEe+UOnF00mlP42d/KDOXYotMr5khOUO6zUA/h2CwletASps3x8/qm
xthFr7fM0CyX2IoRh1FYBvzPqH4JpzE4x1BUAZ5VVA3ZdvWK++y+Ak2vpOjDibp9
Tqs5GdaCivKAOvbnR9PQ7CQI3i+5Rjwh3JtUTUbJKGw8lQrDfaAJ1kp7ozgjT5rt
1P2Gi6PWnwuhcDX/kjn2xGdqpF2G7LvLiCZtLLxfe6/7AwDkCxc6J9dVswMfWjHW
aMhNwFx1SUBWy9xPyJBmkxD4LcDbj9d2VtsSWxgtRjHMS3xhxN3niLyA94bcDf5x
q9IIMNvAz5AQnFBKgXxG81BUDHouXDpLSKAJUUyeQPbgkRBpPaigWE3z6+frfGQS
m1wlq4ce6ZAC8Y8LfZoWvrhfPEEV3biUpyO3YCpd+lq40AwqU3Hf2VICJmZTgS0r
82ROe9VlP0yCoX1kUYqOsHCUZD7sKmc3gDE06SVuULPdXB14hqXjtfpX5YUoVc+D
v0yzNsFCPPWnNEnFguToGUOxqr5xLt3+YlIPXRm0hU3qX4ClE8t//0L44jr9r59l
Cwb/THzQk9o9cXfQcgjpugQuFlKJJMGab9QKqkhJUVSS+UkgtxoqqRCjsLm55tnw
QFNswgdM/wVyZP935IfKlsISHPywjJvENYQ8lYKz0MlVHsIukOC/1W6l7lU0PBsM
LApZbiqYY6AewZXvpCDiEnD+mzfzb0gVK71ePI0dRPcD8rz8Acvil6Log8VdW5bI
qbP0Fk0u9e8LhkWYGOg0Nzd5LBwLg2FB2P8/FlOYjsdy4UPqZ1B5+4uCpXiYXiGb
yWBB4j9RnLDdZaUgTiVYYu/C+vhCmFNvV41eLLrZahK0voVrx8OijLJbjqKZOibj
ZerGrXHhXc+pyDt38M6iqov07NgExP7Xkf4039qnPORyzGL9bGdCO24gzVaRrjYW
pXD10kax9G8BJSMoyksjAD0czfvIabYGYr1OGcRS6EPGHhCyBIv9zQX/iXBhdV+O
B4DaOs2aW77n2piVLnVQv5W2RdObz2+NJYN+UN7JQejnxDZ88pdSD16g2KNJWGbI
CuZfJA0A/wYCoN0lPn7H7cWmeSa1QkxuPxstYAiP/tCYo7r8ofOLlp/HOH/an5u+
JqLBy1ssmfskjQlcF59KFynWz+rnDNCM1Y5S5xbIpawdZFe9Y6xE80ZzyPNNUpUi
AFnAhtGSZosXmnmSImEtuyfNP/wf/P+vw5BdaghpbtWI52aW7otuwn61X0QqTb9o
BRVKOsiepx8/owjv2I6i1nMp1C01qPPeDWj1O3zauW0dv6UEgECJubP2jNximxDZ
A0/rwZ9wn9CDevGnRDC8RxbW+y+c4+sBIIUGkoMjVJP+1XfwLKl0Mu2ZYFaGJ6Zj
HM2D+L39GRcG9fRMkOPd+2+qLuULO18EHfYkcgLZZ9dy4cLRB9AcburbA28XfAnL
LqguJSG/xU62SpFnNEy/WaD9Es2FqWy8wrhW3DHqJTcBte/KkZ4Ch4Sgz8yfGM5B
jPa24r6ctbxlj7ny0LnqiciX/Ar9GLH9SK3Wfu+lJBsguj2ZRS6J7Zpj/OwGZcUr
6gwCUTeOL/TfQHtlh3igPnU9vDtZEWvGQw6mPM8DOzESCyxC+OJlAQ0zyi02Xa8n
lqamoG0RTeeGhz+7jc30fQNa/UTOluNz/zol/FWdpSG00ua+nFrUmxXbEh9iwZKy
t0TT6Hf53+Hxm9xZfrJ/Qm39Vq1CqUp8niaiVg5xw66m0oxFN8dcVROsY6YwxPe+
pdawjFC4mUt9unpTm32pzWeL6Sa1840PUuND+nMl06dGwvc/ULCZ5U57p98/hNAM
sv+whv+LmPOAstO3+nACS6kN+Y6s4ucUUGzpzLbm7Chj03HkmGxa7OV+hZbQriir
Q0kbUpDUPvDovAKw72EX0cabpjn+3uCBgHXjjXyR4692hqVpD09Xs75dms7PYm5B
/Ozo+0J+lyCLCYZfVLfrPagntaywxwwM9FgPh5H8m2zX4Z3V3XQyq4ModAx4zdpj
Amtr1TSMaW3s+lIDRxyhbjmnZQNQg1TjvnI3hc6BPmjS0MAudFuQ8DMREMFTVxat
d9Gy3CP+mxPux/oXfZL7Ag+dWeuGQN2mEcZ5inJeEcLfgWqLvPT5SLIZ8Yb6YKLb
dhEaSsH37i4nAp8Up5UXoMLR9IIRJUU2Ej2HNLM6Jg0ersSee2eMBbBDpnccA7wg
tjQ9OjYzZuJiOtC75GwDfhPzz3CyOlLBOqyeVYOvFZtYnGMIZx39uMie/fn5ui8W
LEg2XNLRhcDC0SqcH74DhkdR6K3tBrjtxR28aIogKFYCfyZ8ifzcnVhjWsfuD7Cj
dqezC/5EJpS9WUSKSk7YbTTgXK7QO5GwZYzCSBkje4QoInHtqWzhoERVdnvdicIp
WKDs/fOHPDBaLSSfzyPvNN4CxWC7hlPoZgUBHNq5cO3su+Uo0Q2KmctIeU49yMLz
TQvt3Lzya6IkZeqU4V5B3swSmnD9JGK6OeTFXlYWVfX04ECl1W/bWZwmkRvgW0wY
hUxtfo8qe8ZIuRqVnK5ugmAqDrp/BsayZFppWKswLuGN6N1fagS5ThyMVum/o+Fh
VY9nazt3j1czBAikK9lor4yMdG3ou9JHtR8+ktj30NcXHnQCChUMV6sPsJOGFE5E
+kCbcWriPfHDRgz1sJuG3Rc8HB+5/gEbqSJBuPiWoWilpNAh5KVBVNxrWabHty4w
cCiiKIEbB7ek/O37VDtJU+PwWJWQbeyEBtqaWN8OsEP27EGfFCooi6hoEAez3ujB
HcBbFa9BThoRApaU6gh7fj7BV9oQV/IvwkLuVdiZ9nKfGnanYQAwZ+Ph7YqXq9Sj
dkI1ITBYC4dQ3zu3prEsTRm0FQKNMQDnk9uAXfQ9Y2CU9451S/ft0JyYHvPtEtnZ
oFoA0npw/msCwd/IzsR/Csu/t6Wz5nhNNTXXgz0dRLgqhLD1SNn8N/n93cvmCFDa
ZAYBMUTsp+85FBBq3PjCDiIOMDKxNi7My9vPyLuK5lO4Y1RrSxZ6OfEtzjXUTl8X
tbUxR1kONQ3DasEMzPMqRpeAD004sXdA1Ccac8Jk2oW7c4/PC76PKyEx4ZFhduN5
WZojQBA7Cks1qQWSTJgKgCY6IV82g1TgWCBvzfrSOglPuaftKob4kGcdACG4ff77
JKF4ooJlCauS92ob2V0YcaOSW4rzi7gjsYwdbEaidKkqVtitkKnjKmDGH1FbSvfP
aLaHSN0E21lBgQ/vQpZ0qBPAhvFmKDs71l/erdLKveWqJOY0P0cP0dlYXoXR5H8j
REh6nryH2T7PKAYjKUqKoTaVW9vy+01TEYrgWzqhbGJwtdwuV7jc8fIWacUjpLtV
xs1fDnL+2PKec5e4LrOX+Db+n15pJ56ms9Fy96O7YZw2I+n/RcdGUsZuDIeIajhv
LImeWPsgSSnNZOuK4FmJ9Zl20cSSRibZ+jY3/UWDEQoUzaanC4iFBBXwVHStWWVj
UM76pxR3HWR8cnKh/+QHNeKbCID3PzrDxw0c8KmozD017zta3poW5RWDopGktXLG
4/ycKdyEyq1kIz8kxox1g1/TXOnnkLy1pjVV5naFRzYX9FqWde1U6a100aXEtFW0
YTkom5C9xeBD0JkL0YV7bBpXxd+UsXHEEiumlLmpYvFCoBDKUFR7mcLiR/Q/J/Sr
TN5dQHQFPMCchXVNx/Ql055XFU4NLodNigwqsdmbTQbd2bZrcgAvLjnFyAR0fmc3
xpqeMA9t+fYT1qUs9dR/fJhd5g7GwpY+sDYJIriALUcT/iTioKPGh0XMcq3rFl1c
i/XjDts2fnNyA71HJOguo0STmRmoKqo3kv12iE0L53D6oTdBahczzDu91+MSG2ju
f0weMx4b/5RmASuPQpJ68HUF3UOPQal4g0OvxcYkco/ARVwfVF9zPJKXa+fiDDdE
MCPtXLNbIc6N0eSO6WK4fzhsveQzzL3sO4c3Fv3uOfb6QXBaGUugOB6myHygYkNf
BGuYqZUYU7r8U0wphi5fFRp9EvaIl7WD1WRkebnNo7qtk/vZTkKidyz70h2jsag2
`pragma protect end_protected
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
oa1MoKxbTh6RFBLCSr+Gbgf8CWJdBfJY5vGLwLEvIcZPF1Z4pSJj1FmVxFwlQ7RI
HQmZg93CdCiLj+oj1dEqbl/xTIf0Y0BDkrUpB8WoIMBrwQbKFtLzgb+MuGX0jx0r
WdkdfC8JU06ucu5zLXNRIn5lp8ZKq09bkl5ORu5ZK6s=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9276      )
clW2dzKam7N+sHo0Evy77fyXFyKZUGsETmlgZMsis2jyO0eusze8XxZ9ZhESsMb7
hy+lME1/VT7H/5gLBm9O7MVTmzNPSqx20cO/qZKh8+ENYMCN9xewe8a9oosilGeh
U4QNGYaz+ZqdbE7Hxd8ifH0FWkM6G/kvBYJhHv+l9UT858Z4rec6USF1td1zN2VJ
uU68Kz6Fb8Sp4/XJaLgBZMRiLSyLyIUJnaMES+C6YLX07FvVBqEHN/AT99Rjtt9y
OGhh+6ZduQoeR8AgqzFBjILm5jU9TNP8THG/CUH43GnhnQO8lm1wbGd5uN4nl//4
jRhIEiR0ceYDUnu2T9Sm28TkiLYORIzNgHbPCxRwqHnc10WFpKAnWGMsQXmuy2h+
M2204wbwogxd9Fc4W+VmqA/FqApumy7b/Gk1FlFYL9wS1fCWKP6+714JXi5se6Jm
JyOOghCjfSa7KoOzp185bNz/SMdrZ6S5+x0yNcH/Yf4mo3Cn+qFmxuU3tZgw9lCc
tQjh9t8kTTsg9xov3M4nbMQ7Gd+e/Vn4Vzp8YI497CM=
`pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_MONITOR_CALLBACK_UVM_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
cGjs23YBkVD/yrLxpcd0JFf1zTFe3CvmNYfSUrNRF3R6DXHzM8j5SSt1qwr90d7X
znt5kucEtDPhh6Uu+ljtLsYnDIZIHIi4QlfsxZoTO6T+0YYtl39OoPwUld4s8bt6
zBNxW2qVGIddnxgy8cUb1+V9cQtitzr8YyqGCO39JX4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9359      )
N3WiwlMDgthkJpviXUDGaKUnuhasIW3WhblI19Jt2DtKKE6c5WFlHuPsq4JewG88
qQQERngbpT1ZQ9iP5KRIQSZ1Z2ABVB72Uf5+2shXv3he2TCkiXP9EnabUDkLMBSr
`pragma protect end_protected
