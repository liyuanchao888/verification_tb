`ifndef MY_MACROS__SVH
`define MY_MACROS__SVH

`define DMA_WIDTH 64

`endif 