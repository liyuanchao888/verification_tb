
`ifndef GUARD_SVT_AXI_SYSTEM_ENV_CMD_SV
`define GUARD_SVT_AXI_SYSTEM_ENV_CMD_SV


/** @cond PRIVATE */
// =============================================================================
/**
 * <h1>AXI System Env Component with Command Interface Support</h1>
 * <hr width="75%" align="left">
 * <h2>General Description</h2>
 * <p>
 * This class implements an extension of the AXI System Env component that implements
 * the Command Interface support methods, as declared in the <b>svt_env</b> class.
 * Apart from the constructor (the <b><i>new()</i></b> method), each of the methods
 * implemented in this extension will be <i>export</i>ed as command accessible tasks.
 * These tasks will be declared in the shell file that implements the AXI System Env's
 * <i>module</i> definition (which is instantiated in the command testbench).
 * </p>
 * <p>
 * In addition to the methods described below, the following methods are
 * available in the model, as command accessible tasks:
 * </p>
 */
class svt_axi_system_env_cmd extends svt_axi_system_env;

  // ---------------------------------------------------------------------------
  // TYPE DEFINITIONS FOR THIS ENVIRONMENT
  // ---------------------------------------------------------------------------

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** @cond PRIVATE */
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * Indicates the last verbosity setting requested by the user via the
   * set_data_prop method for "verbosity". Used to enforce this verbosity on the env
   * if the env is reconfigured. A value of -1 indicates that this method
   * has not been called, and that the verbosity should therefore not be forced.
   */
  local int last_verbosity = -1;
  /** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_component_utils(svt_axi_system_env_cmd)
`elsif SVT_OVM_TECHNOLOGY
  `ovm_component_utils(svt_axi_system_env_cmd)
`endif


  //----------------------------------------------------------------------------
  /**
   * The Constructor simply calls the parent class' constructor.
   * Note that the parent class' name and inst parameters are
   * not included in the parameter list, as they aren't really known
   * at the time of model construction. These values must be set at
   * runtime via set_data_prop commands. 
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name, uvm_component parent);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name, ovm_component parent);
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run Phase
   * Raises the Default Objection to avoid testcase end due to timeout.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern task run();
`endif

  //----------------------------------------------------------------------------
  /**
   * Updates the env configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for the agents.
   * This extended method insures that if the user has used set_data_prop()
   * to force a specific verbosity that the this new verbosity is enforced
   * after the reconfiguration. This is only applicable if the env has
   * not been started. 
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ****************************************************************************
  // Command Interface Methods Implemented in this class.
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * Instructs the component to create a new data object of one of the types
   * that it supports, and store that object in a command owned reference object
   * so the command code can get/set applicable properties of that data object.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' only if the
   * <b>data_class</b> argument does not specify a supported data object type).
   * 
   * @param handle Functions as a <i>return</i> value that <i>points to</i>
   * the command owned data object.
   * 
   * @param data_class Specifies the type (class name) of the new data object
   * to be created by the transactor (must be a <i>supported</i> type.
   */
  extern virtual task new_data(output bit is_valid, output int handle, input string data_class);

  //----------------------------------------------------------------------------
  /**
   * Command Support:
   * Instructs the component that the command code is done modifying the data object
   * (config or transaction data), and that it may now be checked and utilized.
   * The result of a call to this method depends heavily on what procedures are
   * active.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to a command owned data object that is currently active).
   * 
   * @param handle Identifies the command owned data object that is ready for use.
   * 
   * @param delete_handle Indicates whether the handle should be deleted.
   */
  extern virtual task apply_data(output bit is_valid, input int handle, bit delete_handle = 1);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Retrieves the value (into the <b>prop_val</b> <i>var</i> argument) of a
   * specified public property, in the command owned data object pointed to by the
   * <b>handle</b> argument.
   *
   * <b>Note:</b> If the <i>prop_name</i> represents a sub-object, this task
   * stores a reference to that sub-object as an command owned data object, and assigns
   * the <b>prop_val</b> argument with an int that is a <i>handle</i> to that
   * sub-object. It is the user's responsibility to manage references to such
   * sub-objects.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to a command owned data object that is currently active,
   * or if the property specified by the <b>prop_name</b> argument does
   * not exist in that object, or if the property is an array but the
   * index specified by the <b>array_ix</b> argument is out of bounds).
   * 
   * @param handle Identifies the command owned data object whose property is to be
   * accessed.
   * 
   * @param prop_name Identifies the property name whose value is to be retrieved.
   * 
   * @param prop_val Functions as the <i>return</i> value (the value of the specified
   * property). <b>Note:</b> Regardless of its actual type in the data object, the
   * property value is converted to a 1Kb bit-vector. This return value must be
   * dealt with in a manner applicable to the actual property type by the command code.
   * For instance, the command code must understand the int equivalents of enumerated
   * type values in the data object.
   * 
   * @param array_ix Specifies the array element to be accessed if the property is
   * an array. This argument is <i>required</i>, but is ignored if the property is
   * not an array. If this argument is out of the array bounds in the object, an
   * error is reported.
   */
  extern virtual task get_data_prop(output bit is_valid, input int handle, string prop_name, output bit [1023:0] prop_val, input int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Assigns the value given in the <b>prop_val</b> <i>var</i> argument, to a
   * specified public property in the command owned data object pointed to by the
   * <b>handle</b> argument.
   *
   * @param is_valid Functions as a <i>return</i> value ('0' if the <b>handle</b>
   * argument does not point to an command owned data object that is currently active,
   * or if the property specified by the <b>prop_name</b> argument does
   * not exist in that object, or if the property is an array but the
   * index specified by the <b>array_ix</b> argument is out of bounds).
   * 
   * @param handle Identifies the command owned data object whose property is to be
   * accessed.
   * 
   * @param prop_name Identifies the property name whose value is to be set.
   * 
   * @param prop_val The value to assign to the specified property.
   * <b>Note:</b> Regardless of its actual type in the data object, the
   * property value is sent as a 1Kb bit-vector. This return value must be
   * specified by the command code, based on an understanding of the data object
   * property's type. For instance, the command code should supply a string for this
   * argument if the property is of type <i>string</i>. Similarly, the command should
   * supply the int equivalent of the applicable enumerated value if the
   * property type is an enum.
   * 
   * @param array_ix Specifies the array element to be accessed if the property is
   * an array. This argument is <i>required</i>, but is ignored if the property is
   * not an array. If this argument is out of the array bounds in the object, an
   * error is reported.
   */
  extern virtual task set_data_prop(output bit is_valid, input int handle, string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Start any sub-components
   */
  extern virtual task start_env();

  //----------------------------------------------------------------------------
  /**
   * Command Support: 
   * Stop any sub-components
   */
  extern virtual task stop_env();

  // ---------------------------------------------------------------------------
endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
T2SSKD]Xg?eaaS1@GL4.#HSY.Ja/e=9.ZFX&-d=1/V@SUdB#0]BL+)RBB.6O75U9
3OQ49a.ZE.J/ZCGXI::B4Z5ea+5Re:O49V\ZS8=9N_c03>\]ZK,Q@;eM2N/Q]:07
#e5H=E2[<d==52=U[B(+Rd>6[)TcJZQ8(b3_UeHPROa5b=(C;aG,CEQcC)O0=>GM
/E(KMAB=M9Q,L2K3)[.S)M+1L(:,MZ26L@N(U:YSJKdN2,CX3];LQB0+=;#R)Zg.
d68)K<=^=YZ(Y;)T>1a?4:ScH)?Z5VRGb9e9+LY0;^Rg(cC1W;[#)>_874e2UdRT
S1006^^FXV4VQ)#Y4/@GOQ7(DI+Ud+D>3W^US&VJ8JRKYWPI88=7dcCQOe;[U0)\
N4Rf_)BLbKY\)BW;-\7>#G2b?DGPJH,,\TbR>2G_;B@RU/_P(Y9RH@S9(U<2fE8+
AP<>(K]?A9(.:2FAaf,]<c+\>D1#T,PQDc&3#g\[f2T+_T:B/2Kb4#4YeI(dOYB9
##Y+.520UG(gTI0D9DC>&_E9Q[(MRb<1>_D6E.db[NfR7b=2cf0LJH^Qb;4J(7@G
dC7^Bc(T#J1OEYYGN5]9f)PZ.W,T?_YbG:T90@F+ba^LUM\&;-^5HPZ?RR](Y+N-
FN/L&a03Wf=D6+6/[6.>a74^]9Hd-U3&b5CM-9+J&N=SbR>(0&GLXc+g9:@A8P:\
@DPT10RJ3LCZF#cZ6+TJ;LH\fcf+^e?b+(5A^>O^@+:b;2ae>Y3C9,:f-Wb05gS_
)W3-LSS31_=[<Y:CQ9MCF;b]AO>JH64V+aSL1>=9(]XR^8:TegI&KNeX2<1bPQVV
cBFYc/?XfRd84T&Kg60DEK6G8dR^4J=20L(,#^)H^?MHS29D@5)DbH<2+TV=f\KN
^\B[R[Ea-:1GAEO)g-<&LfCYB]9??XEQ)c9/09S<R)P@f,d73?4;;WF8_K]Sf[VF
d7&eFb:91;FKR19>:A:R,X:9FXPM::R6?)WQ[DKHPIK;FZCPH@2NCS8SSEE>E8a.
/GCBJ:_R5E[RDETP4^fD7a1Cd(:&B7].FDP:HCN-,1\AST\8_Yc[-]@60F,fUB\]
-OAa4KK2Hc-H\@R.Y.3<-T(/Ta2GX&<bfPbbF/QD\9H&c2<8QH<VW)6?2C4g7ZZ/
g^07>A&86=TgI9P]cENXc+[E)GD98bF/[:Tgg017TX^T]?K]LSaV_7DEGef#ZU<6
6]GZ5@IBWb>,-g9OGU^LRF^Q.e07;X9,>$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
cKV4D>&Tg1]2T4eH9<SY@/8#a=-^6P[G2+#T,Q-B^b&KR9RP3DW05(@4[0U^4b[/
)ZMRB>+YIe=&d:UQ7Cb;Bf@,3_gS]4-R#454R9B-aG.eN:YEcUQR=7g?8,1P\B(,
Z)979a2&-IR3:F-^&1<5IA/.GcWOa^gU,E>[Vd.KgbbO4\+@I]MYZ?KFa^@C9,&I
6g?<\feXZKG=U_BHX\-4JE&g#fFMRJRD,[4Hg\0R]G83<6IQNZ810GN3+g3g:1H;
W<D6.1VM5P.#)d55W01eD0NI0bH<K]A5?)4>U72YeT3fJ7>Q09&O=P+\g02JaAQ8
5I#e,e()=;=2VEf.KPb4+6;^K^K6=7;[B(H/SYU/CfSTH1bDN?>Y]]Af7RR;BIBF
E51?^9+HEP#\@5ga3]BfeJ\?+<gC(FU4^Q,=2N,OS=:&:ULFc(1>I]YLEbb+E^0T
Z^]LbgE@UUMA>_X8;&YN+/&KWJO5_U4JUQ6K\Xf#Tc1BXNFbN.#,@G4cLX4WHBZJ
7g^/A=RcL:E_];5KZ:34AY#BZ+/DOT\K4K(EY@,GcKZf4ge>23.<,=^FP/RJ:Gb(
6EfdDI/;Bb88da2a2/AO6BfO8QP5c@N_&WbY)6(U/@g<OVAFF\Z2G6NGZcM47dA6
=M[#;G8]\&)-cKc?&:_(D=^c&M),/=\4c]6&d_/Y]?HLHbcWba=bE9(;E@]>>7^9
NPZbZV)Q:?e18()[(?CM>^@Z/W=B14IX/0W0G#=\1=JE,fJ]:FFfVI4]G/dZIL+J
JV-(0>:MB<=^P/9<<1a,)-F0gA80GW6MNC:fC>9JeQ#YB72@WJIZ7V7O+Z8\;5QW
b&K[N3SeFTE9A@,GDbCb]:K3c+.3IK/_]#bE^9A6.NMR204Q-QB+8\]^1P?-CaFS
/3P/D><35>JPd@cN+V.4Q5>PP+_;H:1]1AEebU,LfB42QYVa#Bg/gY].0EM[KYdR
7+O?L^-.>VG&;XY@FG(c9U_4H:Of<d9>f#++<6^(4&FP7-U237D_36Z^3M^8Rg9_
UODT6O[[_^&691VQY=^VT)S<P1?bF?PF=EM\47F^<-R],0,T@fO(-S-=(Aa^,P]H
HDL^@5Tcc:BdDM;d-X4-?9<6SKO^50eX1N&16MCcWbW@KO?VI&-X75>ATU-P4RVd
=a>IEEOLO9bZ=c(Cd#CcA,5a<NS#):GGbX(RENU;&VaDXcce0aNE5OL&d/.--:3_
FE9+>I/IGH7OERL(TBCBM4;NfB+0C)g1@V4G;O,e[0BZ.QBc&C;QIXSdW_Z;G@91
/]\O;F94SR)&ePG)8_XFZ+cgDV&LAWJQ2Q[+;EF405GJ+S.14afS[]OQ>&OLd.X:
(2E7YPFD(R6a<70GE:+R?Y-KK0JX#)-c]_Z35(O&5,V/?Q1D-]&=D2B\e8V?_eNR
2>N)U1=I+X81N@2._dZUa-IQ@U,>PU8g_dADM/23&Y+f)E;R?_L[,695Z;T7/FgA
WBgL667ORLVJ3Ag=b2TE(/>?<A<4-6Y_K:^^<<Q=Wc4B8^-;g_a2X4:M0KKe0E)d
bF]@aDN#W/P;O9[A:UANF?R;d<d+)R\<a=b]T8?gd:4R1GJ(TAQ/dg.I#6J6_d5c
-ZbMK/Z#P\13-gdDe#+JBeCd:g&<N2>IBZVKQJXOgGQGJfH(5gR-G1=:P28VG@d/
f=A<McPBLf/I=KJ]0g7C(+Aa)U]4Jd@MG0\DaOd4OSF]4,Z]Z?\gYX?5L>WB?]BY
A(MCK+^Q]OJ8H7fQaX7E6RU?^IF=b(P-cFba.N7(NW=K.R15OKZ9=3#-d65=0J\Z
2+Y&Le=:19gBKd&]=BcaMG5;g0b^a8+?JSc#GNG30Z([W@DQP-BZ&U+E<DLAXe-F
8Z(7g90IR?Jf9C1+2]:H#a.@L;8;N59+:E(;g(D./H^Vc45]DUE(JTD@dS)2O(+O
^K?17Y(CDL]Z0gQSCC_R\.7(LOZ.a;)/;K.@&/#Ge:cAC_F=YVNL\>EXNbF;WE.L
aFP(5]D,FTNW:)Qg]FBJI>U+T(f7bX.J:cdddU4KV9:#MUAb<U#>[M5(7>.>7\(8
WSC-6OXM/Q&:JgG/QHBG1;YFO)d>IY/=/FY5LcHQDEW+(R4R[_]WDVbd.N3#=_@a
4W4=(@/88[,=&Y+G[-U/_XL@.4fK#HTc@K4A2IOHaX@R3C;(5/>4U?GAa5bU46Y4
FY[JEQZ0S,:JI^(T2#W&;9H?4N>JM=:H0U.C664G<Cg1:Y>4&CCOD-c=&\WIH=?2
c/e4MQ2OCPH@@@[:N97(N#Z:VAY>)11C[F6SHUTHb[BEJ:04/5=F8_ag<]8.,2HG
NYU&),Y686\WS+a+g5]?&L-=J#:a1d&@eP]HF^E/.eIXXg>T_H+,VJBU\c9g]3Ff
CY@K,)[G\[6F-IU>+0(Ye[S9.O?LK<AT1L91)54[J@8D?g3.FAAPCTMJY2e4^GF1
>(?RK^JAPIZDP)I]K9.\<MG=K4UH6QK0PTFN)<&?/Ya8@SPL5]4L/+LV=EVY_1H;
&f+b8);8dF_I9b08HJ#AgS5&Q4VX2>/I<#,S^P0[C?3[K2BI&S+&H9RFM_Z5O)08
?T6;eDZ>)UJ8-KMb,-<0+Jfe^?+/AB.L0MRgTLY\2XD-EgXT4FJ,4R:bMG7SU)Z9
.REb)A[U(EV1)]d8Q_(Y&C#D^+EdFIYPF15bRQQ4YZS+Vc^LUD)5Z1eag48A3eI)
59]+3,BA/^0-G.+SL0U@D:#TY=G\I1QZAROO=2RO3PaHQDM.1]+VZIJRQa9cH^AU
^TaJBFcbJE/6>^O^Z6cbVNAZ\KfW9,bX7HW1(4=Q9SI/PAG3>W)OV98>(12R#a+M
=MUC8(FV@P[fJH20]\O92WT\A,a[PcEYMNK7E<<eMdSf.5LM.>-U?,)=K;I827WZ
XU^4??\5F-IMDafCPN#SPA5e=]e(;^\De69g_Q,BQca,HGLYN+I[EXBDcG=H[0+<
:ZD\I#<#2=7RV]dfRM=_ONYO5a)\DG\>+f2gW2RCN4LZTBe]G.2\a[HWO=K[/P@>
J4/g4TA;@f6#N,8(?_fNNCX;[ZPBBO#.]SK-gJV?=9K>f2Q@#bLQa:#MNd_)Pd2#
QRC,2Fa7B[_7-+I:b6cJ3f4a:W+_KIZ.U-,?;,?G\5?/&6=M@LEcMJ::<7UP<4>@
=]]N+)-)Y00D)T1BdD.)_2WTb6dJH>-^ZS0[D>I=&[)bFA=J9=@ddf?8@KAA(bZ>
FNCRf@TYdc5g5X<JY&.Na\&EgV]U:eDOdKD?&4V_N?DP#F@LJ;S3R:/;7SSef89,
I<5Y.8O.fc+d3>\f6>S@dF00eB,0P\7;9LJI9L(QfeCgA4\\4cD[+;RT2HX/6/)>
S(RKPLCHeG-TK/JgdN,>f(\)A<03HW5EJZBAbQD)@NZONL@FMc1^2Dd2:0B.3:,D
>1OYVD;&6DcMRL:4LKg\1[<[e3I8SLJ=&dD6B/#37@[9/:ZKTOH.>&98>H;,1G-+
2+?)gU8=BJ8b6L@4+;7TW]-((Lc4\3NZ@b3D5;ZB/QFV;U+.24I/ER=B;O7c/>BP
7La[JIb1/A3gI_@I2O2bMb_:XGAb_MZV[A[,:\77WEGDbDF\SFY+Hg&KXR)ZYQAN
H;B@;:_Y.Qc<(:PF9/F#7LNDc?-:_2JTGf[EEDX:J1]gbQf+d4ZId>@gFRNXU;gb
E;;H#O0X?RWgfRdRQZDD.O@US9TX6\]BM?<gW>c+&CR,2>N7.D@;08S_4/QQg3LR
=67R.U#XK]YfgR^J)RGX&M/2QBEHWVb;6SY_(S(^g>K6#7D?HN0=V+=NZU[Y,9[3
,>6<<R8RS#-B2T:.12ATbb]ScV1E:V_g6\7#bT//H>]IA7cI+eX3MHb0Z_+,aLBU
#NE9AYcQ7X&U_HQE37BF-fZdOD,([A5^T]]-@TK<L3F;7<:,6T9[P2MSZ@0WXP-]
8MFF/[CMa[Q#4MJTe80-&KRD<E^;.[^87bag<F?+]Q(9gQE\]4W/7[.KTSJaVgf;
bU3R+MYO-HGE]>WG<1#@^eJ&>2D3;\XW65@D9[TQCc1]7d_eW,[9aFY(e]HO8_a]
3G)YQ4CV-YM1WQVS74gBTNg=H,IFYab_[0SQcN0M(5^7+e9?7_g_Z#(MD3CTFRc=
e#P]R@3J[L7;c+X&PRDRg_>^RX)eb.\-.FZ?&?PG+X:XAf@W&6eMG]720K>@Ag[7
+0f[<#<N[#?8?6OSc^)Pg&+F7E9[DEYfbH2T_LFV_>1GKDCPA(N0REXIOQ1YJ@9Z
M^\#\9eJ35c/a+RYT_aD>&3IV-3QJ-?4\V5+)N7^DM5DI^Q;NOZI_D[7L1^>Y_AO
BE\=.=S&7VTJ^Ia6.3S^PG]+C)?5K4bZ^3Y@X>A+;20S_dI-LCX7W=NK3UaXMfC?
Db0gcdL:<98)ba5fL2<^9SH3B4[/c&+#B.LHf<P44.NNE]9\bB,b3>>?2Y.&2[\9
P@eLFdeO9Gd@P-MegeO\QR:RPA@@/5b_GIF/-1C0>L.9F.-L++=&(7SS)fXMOOM0
S7[^bO9d5bQ.IN6PgP<FbFQ5,]F@RX:6[51(:-T@AV=Ue-VJDdJWIGJWFee1e&=-
C-8K+<.]O<F59aH,[X8JN?7a,3&T5K@:4T:/[EV-g?DNX=R^Q72=OdW(]Q#DU)CQ
PGT[P1G#&8;g677g:>33PVG:dedUb80XC.ZS[S+SZR3UK78)Cg5CcG&=P_a8R>NS
+g<,2\6MQ;W312(QgbbH.#Z>aHKC/G?(+:aW(SXBgL^D>Bc.8aK#KH&7Ue9NN;D6
3Y6:VFPef<+F[Z@&V4I&#H2PY2F+M_KFNBZI/c;e_F8#(4aF]8\Q^/eF?,NPa5FG
dg_f<JW:]Ke0,+-9QaNc,LKU.7Ic(I5U#&+^-0XC#BU<R<-?,]c?DH3F7NaCHO?X
X#2;PKZePeQ5@,#:M[#bKDc@OR<.b=G7WNC^W>G;+35g92R>5UOd,L3Z+=A_F^:[
&a6#PbV=DOUBD_eFQH[Q-d9^BGTaa40@_X,HBX?fD^R]5E7<SZ/8;CQ?HJ?X0;H.
[3Q/BB8@JEXM#\X1f7&4&9@eA^&YHB3KN9d@@Q\/]:1P\+F,VHB@N/g.)8bNFIPY
6>(]D-0O\YQXZ/WQ@/a\K?Nb^E]@aY1KCN[P,9W(,,#L3SKIe=32Ag2#2.4_N<ga
ER(WK,3TFA1#Y^LN]/[ZG8EMYd>a_;;>STaPG2AP/#UeV>#T6bageZ7fd:FK1:><
>-OI\ZX&W_TN)&]NNHDaUU,.7[#8(J#);&_H5dS?)DU)c;:Ae0J0_2)154,c&@eJ
D[d,_^PgL;+W6)HHJ5F,VT;cM6@C.N.fR:VA&a-/#cTf)7/c2SYg[4)fUA.&1X0M
CF[X4:U3XQQ.5+_&EI4@8KaBBb.?G6-7Z:G8@b9B0=SbPSMV7UG?0ZK?;0=#bY;.
MN.@ee#L@SdXSX-gQQZEJYM2)C#;HZ:Eb9_NLRPO8DP?53:\21?HD(g#R\-/ZfY,
-Q=\4_[68b9P&_DRI:f4bW:JG#WaLY[f+0PM&I?B>^KReNQ4=]VbU.(9COI>2UV8
^Y_;I<XSQ^TZ@10HaPfO)0#?@/5HE^]QA<3KS#UQcg.cAQFVe>GDO/(+@FGa7M>C
W@A59I+8\R-:]L#?Z0T6KC&UP)#8.eQGS:_&[#]f]V@?c/&[[0Ve<R[6fH,Z/<7>
O7;cRH7D(eG5B=#[g9.M_9R^[=2@c8S(,c5\Dd3g@DVFbCW3G?LLRefIJ511#CF?
AA4-bPCOQdMH(@-.56eREA5VR>FP,YQC/GWAZ>=C1O06WINR]&?d^^gT<]Y32U<G
dBAKP2Y#FfIC?>_#fN561;ML-_LW[MA05,NP,^X1eB)_(\c,f-GePJ21BT1XJS&I
M6-W^=M@60/3_HQI+cQB,YEPTZ1:U\]2P(8O>8=N1?X8e\_eN<BO-J<8RY[4&C:f
>1<GAe+Xa37&(V)a?J(b4P1^@Q51?E_fA0N6f>-f9+c.JC0Ua_f9<e/U?CEOV<TE
UN)eeQCMaAe<RTVEKIP;Rd.B\_C@W7VIEQ,-EcAaAYg_[,+3R=DdU+2^S<1a<>NF
N+MN?D)8[307:JL)Td:\X[[KFRPK0eG_dL+]+T_V<\Ia5F\V+g3<JBf+UU,2#6[F
/XT_dZHWb<:E99&WN-f4g7_S7/^QHDR#(Y4AKO0Qc9VS4X@P2YSP^aE5?d8RdgC[
3Z#]-e9CKF^C1Z[JFa(fC:E4c_f<3=X-2S;cYPY\;/TSY#4N=>7STFBY<fX<\^3d
00#^SgEJ3RV5F8>2U0474OZ.2,=T3R>66UX^dBEbAERfJ4&7YFJ[)Of9C_ZP5Z26
NTIRV).Q.83ZFdcSCbXTW(CF6aGOcARXZYZH,N\T5/Z[H59/@@KY/IC@.8NT07DI
::,5:>7P<W(LJAQC9P_gIWAZ&A?a?5539H2aWWNa#6X3+=+-7V5.<P.,]X\E7&=X
-C?+J=dF?bWK7Z<0BQWJ47\.LZJ)F>^E3f]4@WaM>4\KH/BC7H_IaVd.Y2.T]M8+
TgfRJ5A.<.;;bFC2)F>?Uc?&:SFU?/d1@Q,QSHd8?Zd3a&]Ka-gTQUdTSQI30@=_
4>HFIA+657:Z6SV[>Ne)9D3/[1HJC(K<?f>5>18Fc_?OSK[A1?Z3AJC[8+aW,\69
]E(b,7_g=d56)M8?3D;](#VO&2/U8VMG.F6]Fd[XIZ8,M_+Ha)#@)@7b.UY6_I<\
[;2,EId(feU^OODQ&9Xb/V;F<VfDA0eeX9C<5W1Og3Sf5].=&PC^O>G>TSB+/Z86
c@D.E;[K.GX(XWSa2N0O&BEJS.EZVe>RK=_C9:J,?3f0BDVD&GcWE?.28X=c3^a[
@a-4]Z+>-8=PRFf\&@f-7>Xb<HGJ-P@(B9._eE\bLJ3I(3T^O+I<R<SS:0BD_]1)
Z]^4DbL#VCV3:N\D[I);C..D6>R#WfAJ3a39:\U7]/?+WG^3Ffb-Hf<_F&d5d_f,
e2RXg8TP?Ke8GJAC=\[;MNOZH6[A#f=TTRG3H))#@\QW/534=RV4M_R/]V<(#R&W
Q?HeDNN1>e&XGFDZ>B\]UZ36g#(d-^S3U0bgd]=@eR+=?d/AI6P,F>/ZC-ZU5,0E
8MU-g00ZUV[E;YDffI2-VdDMHV[?e=253LO94aP]ODTH417g;Q3&(T>1cH6^_SVa
TWg)/0#TEKX/LC@=D:K89gU>Ha_O1#B-eX\E:R&AL4c:KS</N]CEcb=+3R7S7LLY
,94LC&Q2]gOT9GOMSX,U5YaRfK2DI^0O^>Q)-\=B5/H<NgHVQbNX&DI_d\R=^]>N
;I8#e]HDf:S&7+IZ3^\6Wa[:B]#_4CPb#[7SM,@Q6=D)U.##b3TLZN2T,N0G>baI
2Z=O_,45H>fDZQZe.-e=/KLW2K#TPWQ9-MKb3Ig22D/J4H[1H=cFL<N\:;f+B[:T
dXG:K-/(2TJAEFNSV(LWT3W/Fb)Z267Wb2H]aR^7OKP,PLIZ781TAQ@5Y?Y]8cS,
ABPK]3V+@\):QZFS.?;]d)LIfK9WCCXbJ5aM/0LV30b35]=S\>B+Ra/(?US7c<TA
f<aE?ILeeE-I_e2]5XC^;L0V^Z@W+]_&^9F#BK57-V=175cK6]J^3KSaV5OeJ#[_
8\WPK;TcO.4.;a.=b@?e^IPPEaVaP0KF]b@G7_7GPCEI1](V5)53)c522I5:<B74
.GOCE8VQH8R2agWD&_^6)[O65g[EA.Ta>JAMJNWeO0QN?N93+.2eJQI/,>Wg_69Z
QNV\P4bRQaNNaKT>e<)S1ZTXQYOI4L1+gJRP#(aKI;)J:;A:9XQc.<5Z^P[e5=)+
:JeVF2aS]4:g+f4L0b.aYQ8A<+JX=HFd@J>_bNYV:a>Df80SI>HCHOY?D7V(-T1V
-=cL^WK-@7)6:A_-_8/9]W)V/Q/=3)IgBR8;\QKLbg(2WLcg.T1J(T8]f42a+e.d
NKF(KSPJ(+[2dNVg])R9+0-6ePJB5^:(:bB)1;g6Vc@3S;OB6\M,ZWAWf&]#?G[T
2bW1=1X/Q68_X<Q&&#1Z6J>UH].NIQFBP(f@O.\6AILcGP9bYNS1TK;,2ROf:DaO
Y<D4;4H<V#,IM5@3;>;[KHeR[4aS51^]H1I.&+?OM.VRV32K,)fIDI5BeW\/\7<:
Mbg\VF6]06&F3Nd4\63(_Y/H7\CPLR9fXNK&N(bYA3]&+fF#Q7a43#BHJH-<CT#K
:\.b[dOD.NJ3cDQPa0/+4PX<;9JMS6;QK=[[ZQegTZ^F>[Ec.4[T;M67YJ7AI/b8
CX6.O\WPf]@IWB@UdS:^3-0@af7=:bb(cG:dRI4K9+9GI.6Id3W1=]P0^CZ,N,^G
8.FPI\<-8OOWR_UAA1=VfcL/V7fE_L,9W8cZIG5IRd_g[VHJ;87@aZbJbV)8@;/-
Jc0LNI#FA7ND=BB+D]5+TIWe2</FCV([O>g@6#BY\_=G4K.N3U3LbH+^2F);H2^[
T;?Af?f?fGf&,KOKT]Q@FEJC2-5DDg1W&3BHQC<15D^\S;X#X-Af+7&9__X]-0GD
2G#/RR1]+=:>1XLc@[)ceMR]TFdF:AA[R[>2S_@/1LE#G55_V>R6g.Hb#cXRXX2+
Y-C?:Z)DGY#DC0>(LdHXde)Ha;d/)H[7S68fD4</3&K_H=IIC70d_1<cSHFN,WEP
0JU_D15ba:-Rg1dI6F@?X?;6A):XcLe[d&[J0QK?/c[K[\d_6/>g<-2()1VQ/@ON
M,SP/CR8aSTEAeg-VAcL@0OfG-ST88#]/PVgA#&K;L_5?>POU88OPCb(;D<;\2g<
5/V1Y.Z[&fA=;VX#4c=cc9RA9_e:2)UAFI)Z8KG<LdYbRFFX(_fVGK43OLB6b[?a
<E4?1I&GN2JK@WS<WD@A\dg:MY_)N79G9HDAf;dT&D<P^V^1<=/:X8=)_NCUe7/D
PUYE,bCA<Z(TO0H#Q8aWV\G=#O3Z5Y;d#RI4]gd=-[V&[K^C87V_F+eIMIe3G[aK
WE#2YB>B5b+W0^58Y(N?,7YUb(#F5(gR]@>g9bDeA?&0X-(aU]WJBRg5QFE8/4:C
&F@TIM=QA_F07Nc=P_H#)H);FNG5.^5EG620+fc/:2?FEZ?^5@#&gM&eE1]QRN:C
g.:AOCN+QCKI,bYK83e^L@QG:::JQefGH;]<caK[fV7X&a2C_(;+9I=[DT/L9BeW
,\UIOdQ#S/J;K>1YgQBB_?R[9FW.&1C,B+1YSQ;TFIQN1ebb6:)d#3QPEI]N[Q[]
NBb<LBG./DDM:^^5U80GEQ43(#QfYbTE<+IEG\5&cH;JVGHO>@?L9,R:M@bKEJEI
)<_WJ0XI[[VKL4]L7>]85bfDVRS^dRC269R95YY/[E/9&1_J(b)556/?c,P5?<&G
8=R^U6XSZJ.^:_Y7]AC2-SP^(<C<QfIJSJ&:7@SgcL<^0P6O3XC])62^#[DR\56A
+FN7)G,FP]5OLW1O84.HRJ+AE?2IP97P,RFC6HfW&MFF#Vb9F+W@CGAUUa\JFTMA
R^3]?Y:05\=PP+H<4XM>c]TIOO(HLf[Q?ZYQS:D(N)&1(=0_;@\U+ZfJ[<,V=(QW
Jg8H/&XBKAL;ggV:4J+[B._U1b76/]X&13>b6eT4HO4>A7CbVLK6<L^g1,1]);de
?F_]EJF6QZ<=//YX^@09J&-_Q:,7PV+#06d_\&#Sg(>?V,:#D0>M#ZYH8=\#\d/,
L)_;Ac?aa3+8_&+LRDP[JC>S8DK1JKaWIENGd>P62D?T(KFGMFDPV4N+.ZaPG7[=
fe;H0A:/XA\AJNS>VJ=33WP\&S<99-a7A_N9.fAOG,<<gQ:\@HCe.H(=[XQ&&-(2
;/(X4fab^5/Z96a&]G1>,ca&Y3SP#IFO=dfU5666d,W7IZI;-)^K6Z0XB^@Pc7#M
I?HD->XT,6[3gNF_Hf#80Y4]EG37R0e_]=1^X_1d1HY]W_bIfNX&G[@U,ZGQ3W2^
W+GU5=N?Y+WE,3<eDT,agYR2_W\+3HW6Z(f/J:eVd]#f6_=C4XHJN\;[87)K1b]J
F0ZV>=3T+Z^IdCK&;2ZRCCT<;^I.3/&?:bVCCA-V)b+b]:X<PB1K,g7W?+-c#IL>
PbW[P^a^#=&R(EXRSF[-bf]6):_9Bg-<?/QOON]>XP9?,029,J<2W;YGfEK68Q(4
A323g/S(@62dD.NBW\Ib3<J>R/YEDJe9STZbQ<-K].@>EH2cM&4T3JG42GL1I?SY
79]6N2cMNVg>VXF##V3,bO;:VFIfQ1Xb,4K,?@egH=>B;PM-Pca>=7K8PfE2#(_K
Pe_8F.Rge:R^1A.03C3+282Q=+R(bWe-[HcUaX/PYP4,G^\(cW2^HW[0)Cc/I@a,
5Qfc\M@\@?>QZ/8L^<a/\91INbVW-[;\/@[N0JRQ+TfZV&CLY_URg&<(&D+YXZ#V
Y=Ged(8J<I;Z?>,g:TA24,YFVS?4^6a)[Xc^[X,YB^U)TP=>CC4SDV9?@U5NYVBT
?Y4OW5aCRRVcGU3WfV:3N?VMOJM]O),.CB-U#UHP_RK#K.;N;)>,\[eAL@<DdS]]
39Sb^(gYIE@WT:>YG+##MJ2L><B\RB?WN02MU.8)7=gKbNIP1;+TAMOF/3RV+8LF
U/c.V&4g4EdZ_\M0Y9PN&Ja?V1HIB:[fH/T4Z7#6I#:cGQHX2KN:8@[g39^O[>)?
aVYJC+M:QO=-?8Sa^JbM?J+d^N6;VQT_9d,=;NSX);G)+F:ebG>N_9KP,FFG6.Y@
@7S:?I;=F=<;gJ\bIJK)O2ULU)#C#XSMO,F?8PGD4OP^V(^)<@f\QKD^:X>Qe:-S
]7[_C=YO/HO>b(ab637W=YFYA0ISHP#7a+^dZOabH^ZeHSFaJWeRRE)\@PBDMdO8
ZHU#24U@F.YYW(<->S(Pe9S,1)IRK2])WXc/-M/L,H#F2K<05F:AbAE-0_eK1F#8
cgU^D9K9RgeQ7daf3;1LN6N2&)>AgN:)gRf,UdR(A:(T&40Z:?GU(/aYFC]??^N5
Qa6R/-VbSK@4+EMc4fAE90-gFM&fK44;:5I;[;.RK&aWODA_[9=NY57LIP0=5;?3
3,UbK:-YSWT.&B.bK[Lfe#^aSC6N+-XfB3NV]^@ULOKIC6DP_eW[e=_dD[gde]<d
a;P.aIU0L3\MK2eZW5])0(\FdfF+:AH?A=?fC1UQ7;J6ZS8,NNFGM+&;Q.56>?g3
T7]FUfVU.]Gbbf]R^F-)EY/Q#3=bdI2Ye56JbbSH[^,M:VHcR:UOMV&FJ-=#6b^?
Z:M@=;BI:X0.]K^M1+5>cNa8.>He]YK8#1+EWd\\V0LC>G4[6B\.O#MFc<+_>SAb
=)#.I@4M1Nd?CKVUJHCM/=KM)Dg^g_D;gd+4#PP7[0cA]ga1>VOZ3fd5Cc14R6.3
&O6\AU2VYQ.AY57cbLN<_aRH3H,.>Z9.Y5Y1@UK9NfC@cS56P9^3<@NLUD-,/9H(
Rg^5WGTR6]/NO.W;cXA[RU](fdN43]T.#J;17Kf[Ve87S;e,afVV/\M8]fJ-)J[g
ISHQ>+^fdISF5YQ.e]Ie<9\F,MbaHKKEMUY;bND#FP#@U7e2fBV;aJ3[MXTZ.B>+
IQ[e?-XYYDYUeG2-93]N-1PCO?5gaVT-(J=LM^(.P,D95.GH-J.)(:VbWJ#?K+4^
(<[CHHb:I.>./PKL^+Rb8<0KX]9\SQ?V29E>D5R6N[U^TZ57YY\=/:^FNH7>S9aM
SGO?O?>4M#c)Cce6I05S5C]3W(P5^2><=-2-gb>4OP6QX(HM^3\_E[Od@(9>.P#6
NO_-WM,(J6aGMcJ=GU5f\NACEdQF31e^a;QMDYK1GV/bfG0[ZH\e_f>A#>1&]f)>
6Dg-/G)_WfHP@KNg.>?@d\IHYE[cc2#DBO)dY(.a+T2>,]-2/J351Xe+8:++F\F0
R3@Xb65KLHL+a8J6J>DT4ES1T-?LRD@(KcfZ^9BaF?2:ZPTVV2>W41@]B_L)^Xcc
X2TV5HW7[R1cZfE^7U;WHgDNd@LBT\gVCU<;b>;.LFAM&C;F4AS)#WIF.Pe;Q/],
,9d7,+eWVScfg)DT5+.+8Ae3X=6].M]Og]E:[.8/5A-&?:aLLg4RL_)ZHAT@C)f_
f^)gRU5+Y6-3<1)>eV+;3@)EPHR26&<:d=K-WP[1SJ7.A[HB]2/@fbN8AHMA2BJ;
B)/&a=0[-5RQbROUEWaFQM59(<N3)Mb[,VF,JBc+O5G(P5[H@5g2c&PL^,N:BK.;
FH#59SGC<eL8@V9Bd7?BC/EEG?IM>YNH]?RbY6#(.Z;3^;2QWGX.M;N0=#N.L_d&
gS9V61GBROWUH@M+&^0/8)92K7+Oa:2GJPbUHD\e1-PD6<X@-5QcR7J,PH(3cOVC
OA3D_C1;#c?_TP#G1A8X<GeYF&,K;1Ob[S.Y0S8_W83;8OWP[9NQNd7(56.3UAL[
=MB3V9=f2dX>#6?FdZ<e=GCg.F,(b,04\g7SaUWLae=S\HCFF<,;:P5NFH.2KK[J
:NW4Y3R)(Q#<eQDV/06=1_d+KUF:,F)g)9_-PP-I33IK37<8[9UE-OT\aEa,82FG
;=->Qb9aPL(dR.cQ&HSGg+#IE<-#.0c6&Z[YK/_b:0=]+_f0Yg+cU>QXQ#3]+[(6
?.d\;4RE^T:T&7/C-fEA)J)VD1J1fY=KP&)f)7SVb0\bfYUYTTDKPR67RE6>67M@
YA>#aR:>RbABG;#V&a<2510cb_X0)-f(9fABYT6;L@\c)?T+S0\AGd?TWA29&N4/
:T4O_BZ90;+bgfW@NfDT40MT+2/?bZ<f7@/fK0IIe2X1^.V0&>8=U&ZaKA(eQN/.
)&X0#]D8T@;LbK4NX8P=;D7QH&-EFK@(-<(1f/>U,RD3&QDeSNW=KYdPO5JKQQg+
=40\DRUFQZ+E]5gP8P?0e&PcTG1H-6<=4[)3ZV2XD#Z[2S.)0DY=TQ2TeCKFE?ee
E:5-Je[0=L0AGN0N,)J3R#SCWAa3BMKVA4939J1WUae06\AIV,X,5b>H?>,;2R_g
V)c&W]7GdU6Oc_bFR)VTFD7-+@\f0(0OB[<455;c>=aH[QN0Z@@d?bY&2gEXN/7M
Z,fcbCLT@7PD;)ae(,2Z@T<X5Tg.AJ2X9=aFH_I=A4)&dBB.LK<#=DWY?/LOV97N
5f454HYJ:bSY+UHF_bYD0#>fB=LK]IL#a(,NRD#O[N2P<&/3e+4&.^B(QBdD60a:
;#P46I:TI:U[^D/T8COO.A^O>eX7+ZTR3]K:d.OPXZ&B&DGeV74ZIGM7D>ZQ;[/(
J5_>\c93EQdN0YA#2908K8L,8:48T0GeT,]::<K:OS&9SOW/G=b@82XUNE0XP?FL
^f+XE\A]^a23:(,=cHK_f:X.8JIIG5L6U^dQ5)21fYXB[#\g\K.#ZI1Y07Jcf[g[
Q9bLBZgZXS&GD8OKS[N2(3>TZH1,L5_,)Z=Ud+d4LZ2J95=(7&;#_/[CU/6^<>MF
,UH&TPJP\40TLF6IFF[gB[/b5</2c9dWeUGT92<DS5DG43&L[?0.,6XYN-QK_+<,
ASbXNG#42]J+Pf<IQQ+-2Z>5(@V(_gO=52Tfa/Z\?P-N;46>bZdQ)M>OKFF-FHCg
.X(/C4)8(ET#UK1C@cb^=Q=DeE5DJ?BMV^-LKaMe4JF?108\PMNX,EXV\A)>0ZgH
4/JRHU9V/C0<Q[B[2VS-(8[.TRC5cP2B&]a-06GPGZZ>\42YT<gC,8356>:fAF3,
Vd-a:+\aH:)A_R6N>.0)W8ZMFDA)OPVZC4AF<WbO&\A2YdWQFDB<1CZ\0NGXb.W>
b7Sb&P^<QL?A68^eR2>P;R\Gf>L-DQc^1W,8\?g>5@R==@U:GMbETPTbZ=<)P?CA
DD@;]<7==^3+,Ed@A2cFV+G[D46Dc_(WN\=0_B@DEgP?[VYA8R7SWIER,M>WDLI@
)Z#,?_-::Zd<PODW6d92]5]JV\^IGe6.NO<K2?:B9)K\g@\dacKcWY?[?)Ec9-8c
T+EIfD;<S/0F:G0SdCAK#;3+P]G.G&b1\WQGSS,S7P0gR;QJQd6YWC8SU?)T]-,J
T,_^7DaE0>?aJUQQg,;:e+]_^[cf;e/LC)Z+R6<@GB,cHdf&gP<@aK6WH]3I-F;)
[1G^gI\,R,gM2Sd)Rd0=-35Yb9Zg?:5QaQRBBacE9@KNSN3]+4U3);ND(I_Bd)We
]PGR;UYW>S(9-VX(fBD,-Y6GDC.HCDOCUeG\bLY1F?AKA@c]NU/CVIF>Y^^eI&;@
#;X.gE4.P>gLKSO2:)/18C<Me?_-Of=ReJV6W[FT)ebY4(.V/7Z+/P9BG;A^PHJc
/6W/#3Z85O83YA3646UQe\BQKbHgT#4\&FY<C<404X@3LG3g,,EYM#DMO#NQUC7g
4e0&^MVN<\G^7R8X7P#-B7:OH/AE4La?0_Z3X;J#1FMQf]_e6W)H+7;XQde^f(CT
??./.\fZPg3GF1VTNL-QE:#T]OCD<\99AL&@<L1:N:CY9/ZENR_/TZFSZ-,4>Y(A
1?E<b5(,eIVL09edR,e.U#:DLVO,EHc<b)-.A#<K+Y02]J7XM9KgNH26?VP^C]U=
GW>BV#LJK7:OLITD,W).A+2ULY6AfZ#40OS;6[G)+PdLbSccDXT:F:2H=^eeAg)_
b&KUV)=UU5IJf1^b0T6c1Eb#/eK8<dNCLFDe:f9.S00R=1H9e6.de\@4XRKUS#eZ
ZU.W-gg2(a?GJ8G=3PPd@GgB(P/7P_QBAWgb/B/5H^PPN;R:IH>d2&@.MN\P4^).
_CKWFMaa^)CFeYS<K6_291X2C9]OBN+_AH(GGcGL6JL[,f8\<E>(,IQ6Aaba:DWG
gA+E9eN[?(M###9R5>.SO>[CI:0g82&6AH)]=&ZUX8faSf6]?EJ-b,V,]ISJ92/^
8-7[OeP7f+2NAG)1=EBd/M1Ncg5)(&edA4+[&XH-G)09GV\[ab(;:[/eD)a^E\bG
J)ag<W>aegKY11,YG-DR8Z_1H6gXC&VMf;^(3gGG2PFIe?X(W73;f3V^#ZJgg,N?
G&,c<;[55\&MeN\Xfa(-B@6NNfPWa_&5F>C#fa9P/.XS.EM-0@D9JNgGD:5_E.:O
/SQ/dcB9PVYFCF;TZY;2[N^30R8_C#?XPUR+S8b>G_-V@8UERZFa2]eW,/G,)/WC
RN.+J<4C?I76^=7?,[_f/?gNfTg-;BPdf1E8G;)6Cb1SJ7_7439,cW+^O?,#ST9Q
2A5gEcL(<ZdUG,^cTF9YY2dK=5#F5X<AX8-J)\cKTZ9KZ/#P;6SK_&\NQ8-e.;KU
/Q67LHWECY6WM7f:09.dVDAbL2YB_RDVA;BBf3EPK:U]9V[VPJPaR+#[YeAX1OEe
/b4_e,HA;,A4NAc6)=-X\UNRc(T(H85W#W.)^_;YA\bcPXGD-VUgC1;g?+>WNbcY
IS(2W_O0:LE^DM+1WG0D=PCD^<HW6Y(RVc6aAD;&7D[Vdg@0bJ9e,[bf:AX#JeP,
S:P7>Ka[SH]G:X@E4N&_dH#ZX-K&aPXU/Md3gfD]ce\TaX\.8Of_Y+M],F\V/TR/
5@1B;Y0C0J#?[MF;/,eJae[/C^bOINDcU#:eIZ#2?U?[>BW2f(L#6/>[CYg]f[GS
VfGA.Be.4TCSCW1GJMf90BF-T[IF+\;R\e8cE,YNM2J+5<#MUAS^0,J8a;REg8)(
b<>^H]GE4E/SSCLa8R^(F0dCa:9dHR:+@7CF[FCEE2VY:Q.EHR]&_VgRY4fWOg(0
U\2g=X3&EM;BVD_C3TEeCQM-&Eg7PM5gGVBA-\\8(QHJYK_H]RPGZeJL-A3-D;De
2=?<d4HKE>QR:6)cdJB7X^6MXe:S^PC49dSH>G(T3^XL+Y@Yg&DT>a]&7:KD.>Zf
E;HJg3aB=SX20\R)GO8g(2@a:S@b2JBc<>#,9\I7;CRf7eG,&a[f?XX&0=SUSUIg
#>>J447;(g235@\7-dHC12)?gbE&38NZ52bPc:G.M5Q=>ER22:.1H2f+R?P=JCD4
C80464AE&AD0Q2P^d-P73,d@DBX0cY/#V3S(5gWL)2eXC6MZPL+bC>[@F:00OcMH
K?4Za+cC=PaZ0,ggY\Y8:R^U2Z)KO\Y9]>TAMaKNW_VL2.>4fG.30,4+cYY)V:OI
JHNHD:a9LMW+XE0ZXF^a(F1LW#2M7GH4gILUJ9KTE0cT_VK#CQVX7ZQJ7f>J>K)+
]aZONH5Y?&X?J,M/6EA/V4\gS)CS?)eDVTE+GZ(f==gL<7Ad2]SV^GO+.CM[[f^Z
C=)a>b.Z(B2OT:Ke1VJPPMV6KUX2840,0YY>DTNF:[0KC-8HQE?JG11+.PJ6)BJE
PX7XWOG,b+@7M?\.-Fg@?[&J4A;?\:J)V[9^\135Q;#-E9)T8TdH01PHMVFSR0e[
12A5SY^3?f9WGd[&=KORNSQa.d=\K2JDd@?,[dUd@F4TB1MPKdV-(8IXe8&Xb(Q_
;W6dSa7)BD@#9?dA2.0fbX&Y^XS&\]\D;+df6K(S0aZI&8BGL#A7NRIOQJ@<TB95
N2ZZM&c@e(He7#B?H>&7DZ>SZ[>g+9ZD?(=RHJ_Qa0AeWbN@7?5d_73<GcX6^]_[
?@K:.UD,G<K(G+:KU4O-4FNGZO)&6,0(+A6NTUe8[ZN[bb2LDfQ09_Q,3D;BU_+7
HEf@R^L5,7V-;aL]#K+eF]@+\9Q:AC2&0IMATF.5-/\b56D#GA09?VYKV[aDGY4#
BeVP^=029&FUFaVY?ZOgF3\f7:e_D1MbYX2F_K3G34@^MF<0.YTcL?3VC.<cQ)@Y
Ie]gV3++Y>&7O0>,7RL5Q9)P>N+6+Y)Bg=8AD2.U<e0dONQD_GH<]\0_B)+=/VW+
L\/3eRX9>\9O]E[3a=]FZH(P@(#9))W.JXA5[;UY:(e1a0V@VABU_5&NE/WfMZ02
@/=f+8-0CD&&YPYEQ?768/KfSe@e7YZWGLDFG\C5b20I1-\bKBS2dd+Qdd2F&ZTN
/+e9AI+(b)@Q:Hgg6S_KJ=-4f/B-.cd8-g@-RbV)4-A<)VZc?_f^C71SPe5RNG.^
Z3E5g+/W3SX:LgTggQMUXC,8OGD[:-36,Q(>I[<TX=:UH4\,NKcU,A9W4TNa]KLG
+-4+BL)R\@^J5QN2PY1TN\LZSJRWF;:RVa:6A0QQZ[_HW=740g^O4SB1A\a5\&\#
U;];,^M.+QUGG>Va,-e/TQH]^<G(B5D]f__ZF]68>2I48X[D1;?D0/bDE=VX2T\S
Qg^BRCKc_+CCeeBOP#_\H7WTF^e;?&K/--I^bZa(-0Z7<1M5b<X=I+#?)G1J+bO5
:WF1&1MAY\Wd6WDbKE]A)XBMM#e>KQEfe\R1=,ZWM)72dgE#WD()1a<D@_bO<d:D
P=&.ZJKg@;]?UFJBGaP<]3D4SQOBVL<+;MT\5.g+F?IT#D4-5eZZ,(c?g.IK8,65
9,RWbBT#RWV+^O^JI<<CU@JeL5b]_a>V:2V0MW,8AJ88[ceD5P_OO&:[<;<]5fQO
]6?Ae6Y#[,X_Q@VJ=(8e>&fZ_b.B]#TNF\DT1\CU_,c7C[E7,gH\3#,?;Kb:6RgA
&-<:C\=HWN@H&/g;XM_TAK/^..]ZL8Vde#,g[3OfR=@4XWYMgJ6;3I&@VXKM##@R
g3g5VSZD-85EB#-TN@;K_;3.f_3ZGOc+L62NI&e2c)GPaXK4ST0[E(=NGbMO]UD9
Ab&M?0=O6KU?.O.6f[V?MDB&VZbB+gBQ+gMU<O?NVP9J/1A[^[]MV[TZB)a?:]PU
W].8;_cS/?T03N2c[=G>bUM90AEK?QF-eAA(KeO=Y2F4Q\/;Od[/SH/F&QX7<EDX
Y]VACaO@<ZF:<<L)<a5UF8F^PX)S_FT/<0>+R)MJY]aY7Bf]Z0RFC8U>8LG<B/=F
UEX6<OH:/)ag5GgQ[2S)DTP7.IA8^dH:0VK?\-_<++0_,d]^Ab.72O]AR^]_Wd]M
/BLR2aRUd;K/4/5GBLFc1Gc[(^71&5P[<,4\aN#&3Xd;4WJM/a+82U]AK$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_ENV_CMD_SV
