


// =============================================================================
`ifndef GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV

// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Request Order Write followed by Request Order Read
 */

class svt_chi_req_ordered_wr_followed_by_req_ordered_rd_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
emchjl51Eo0rHqwZ+0bI4mhUN+NZkVrdhyVpYJypWR4+cFy5Y+J8Fie7EjGmmDZ5
Jp6YtTnGArNApLVk/eGzkh9+cOAGhLR5RhpXuGr6CCc1tXpkMcvsYEnueyogBr05
vYfnq8wiPebRItwQWZSQXQJ/9lwx1GEuhYdDOwO9VCXJZ0M0iYrJrA==
//pragma protect end_key_block
//pragma protect digest_block
XQ27COTopVkR0g31/LSKg1YoERw=
//pragma protect end_digest_block
//pragma protect data_block
EivzCX0gGJBV2d8Eu2Kigb8orb8a1tqXKbolbWsrPJdtdjRXnfvpkB0BxXJJa/bV
+mpjB+XkSJamcAWhHR+B9deY6EDPW6KKRnFdYl4YHWwXS8qGkQxBjKwNkIHWXLHT
4OOSHdxc9bB9MMYjzOJnKFcPzL/u6PRGH4XaEqN0rpyivkouBXL5lbleCn5KS+ng
142Ue6WQi1Ih/BvCbsohKT0qFUlN1n0+NTOtnfZTv25lkWHjHa1dnAnR2yOFHWg9
/8Z8EUkhMBg2QUh+ljPkDd7eFT1LvCvEe/H31UecK2eyNSPz/7NTnARfXf6Bo0xq
nY9PTCpyGh6dOxXbm/9AwjZ0os2mbCCJy4/dhXlPeTa5hXAmaUf5Cfq8ibIShUUL
6l80yD9Qmy+tZDCo2Rp3s656AzJi+i4qum67+0k/w5w63Q1eTjr3QDGZWwNOrHne
DIssDLGOZH+g7o8hq+DWECrC7QfWzh1MDouzqRR1n79xvyWs4jbzV/8WBdAS61K9
3sSE5LbF/OBWTYWVfxMzab3MrXDkADNcc/mibkpUfAJ83orCrh337il27vtTAVeo
xSfhggWA8gyCjKzxlnFHtZLIAE4ll0sQVeyYPuf5WaaHkhMuT5WVcDHAsyFqN11a
DnT7ybHEBsPBOMNkdpv6xD7SpQ5C7vPOt+XXSkQEMzBlxqimYZ+UMvd/XHux5XrL
zuBLbIJcUP+KqY5ivwiV7ghtkG8oGNvKtx8ndV2Lc2/PPAasqBIx3nfygPrhNRtP
zleYs5MVgYvwXRD9lXXTCpeup8a0fLp3w6IBR+/YF18ItS3A80Z9m+Y2qLorm2vs
osv//id7/omtaarEK0ygTx5JOdf5jy8YJJcIQtlng/GmRk9ON2vjT9OJuR5G9ekr
rLTXXxlmgXPJXXm1T73cnB+Z/WvYRzjFIjb0Qhr1KBYk/vdCh/uCNdxUwtljWD60
1vRmpxXQleIrCnMEHWHqmWHuDIZacjWfsmmzKsjIOy0eEThGyZxuFGJZqJsU5AXm
ETaGfwWO8v49+VUMxjz96adetao8BujHEchddnXGacBKBWo9MfnarluuJFxG6AKH
vk9yG6P49uXe1Y8UxNRkeA==
//pragma protect end_data_block
//pragma protect digest_block
KID5p0OUDGizOZKtB2CCDE94nkY=
//pragma protect end_digest_block
//pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Read
 */

class svt_chi_write_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8VC8pZiQ73hWi0NOC49k1EOMP3hu+fAZFls0tVG7KbLbJf/sqF0MCZDIZx5WfmhA
sRW5JWlp9/Eiel3IhtY5oq3QBlaQvVs6n5kP07QCk7PwW2J5O2inu+kQ5Z2OpxZa
FTR9R+y01Nhy5psOJ5Bff2VJad2IAeAGvz5vrwcBQJBM361y3vDX1g==
//pragma protect end_key_block
//pragma protect digest_block
6hC0WlEq7vuU0xcmG6SOaaaQ4cI=
//pragma protect end_digest_block
//pragma protect data_block
F+V1CI/eh5yGLvflGxEqgO83wosAvaPvzA348RqKyl4SPAVX3LIqk31Vx/Hr6SFE
KqV3XPGzpQfiWmekKKSBiIubdlnS57wlEr8UMm6xilh+w+MmQ0FLb68lMkJ8k6ab
93a3bitoAJVWm0WvldWE02vbA5Ht1NUkYQbI4QiWzOlrhIhu4L/r3qVKvbpkyJYa
S8Vt9jbH6SxzrJfWVo7mrGU8SZ7h8DmSdOffqpLEO1dG0FoUK72W0T4CZenpEqE/
ItWIhK2jfJNmv9h/2hifnMg1Q0O2+95zZp2I8p2V9t30Q7YpNd36wu9bnUNfRmeL
cUpH6PsX78+Po3wqHAWVN74bMmykY++8mPUAZxtBSal70GZgKR3bDzOw/aO98yg4
KQworCaBYd/B/kKNjE6q3+aXLzACYA7jKvrXiKhnk82XeIiTmsShP6+4GuhGQ6Xq
NexR8rXMNackPA3Fq7F/sLDyTk8XsWrfxxGYHKQiN8qGpXtTDxbseaXMp8ffSWsk
1YBgmz+T2jQDvg6RmjgHvECLpTJ+lE93VuMe1Q4KuxCL8JhU/+IqDBzcGHLBS8me
xlWX+e+k5AnfCICsgzMoy5onxhVphBEvQRpH7Uns0MimUwHr0KaoYs+CMs/Dyl3c
ozkE2Eh73e9lFC0w70tjzNkpH5EjSjIMBs0wpv5hex7jvJBo7nZLOkrKEZneylEQ
HU8Tx8DwVhKVYxbmxL+XWXTEwb2lXOhY0ZBfYJ3EXnGlKuFIGEALWpKvTCrB28U2
AIw/CtBswM/6OT7z+5ObyBOqWGwksLJzo8OD6cJPqk5LBtylgaOllpmNYCnQHiP0

//pragma protect end_data_block
//pragma protect digest_block
MhP738z8XFdQjwjuOFGSAnG9qS8=
//pragma protect end_digest_block
//pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Write followed by Write
 */

class svt_chi_write_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DDT3vfIuLWgxZV+Vhu2RicU6ywMeU+fYkVmwQx3+QGuBVh2DeLKFkbtcOO0Va88b
pzvrY6qrQSX8jkJ8PmzaSyMUnt5QuiA1Lmpsa+JAS896RgGIyM/vIbhSopLKsJHG
s7u1A8e4O289XqaxlPVvsUdFvHujx6Z5lmzWTEojFHpw471CoucoAQ==
//pragma protect end_key_block
//pragma protect digest_block
fS4Vp6uSJ5qe4VjAA3/8lAwTvOc=
//pragma protect end_digest_block
//pragma protect data_block
ogHsjXx/RC76IzGXvpzmZ+tFU81P9M8oB3FOPlMXVNzDjSV7eDV2sa5JOuizto2I
exq0xMrMNLRoZfr85s/1nFREuI45T6JWLcXhlOGPHrTK9fQTO9fUqWoU9O6XJEaE
y16zjVj6J4uEzlOWEC37XD/KnflRqb9ZvIdfVC7Vi17VP7GWxr5B60YQ9Krj8Nul
okrdGUcaPExcUQvrytB6ngh96iiVMmLWJwF0DPWUv3EeWst44R71h/wYLiY/IiO4
0p292qxIug7vF5KqRJZ8Yx7VRDOttKnXNm6LxQZHfSPnsOZQLwEd5e9Mrwbrc94W
DA3D//rcT4lGT9OmrTJMqsRmV5jdfHz51uJlVHVJbMlhLEE6brCQFlBqj/KZ1OZb
DiEsL0CNe2cuUbYz2Y19JHpacNTM/jHkXjcZc4w7VF9JsALlAz5w8u3NNDe99fjp
pe7OCeNQkxgV120o1JdiH+WGRsCa9Dc6jAABr1arkFPrPV2Yi/lf4OXP9yzS5CMY
SlkRxIiWejfMEJchw4uloKap0HH7HpnzanGxI5OEYVzyiqrp2k3q1/f69M0wUHrg
GGZawD9nrNHKtOphi3mtigtPpZFFqjRpBLuCO4Miab4wk9RmkFMFZfeNyU4n1/R5
wo77VxvR9Zf0+8RHI5NqhR4TBCST+Sos8U+2H/aGeD9dsjp/LKocAYHGj4veVYU0
zf4vYrfRwUW8FlMWrO3S/1J4RJ6sXpAvMZ3vF0hsA/IIraC004Gj2LvP6pkr7RB0
3QS167YOfgl5uwByNPMx9DZKO+dPkbqIdbGH86f+fzau1FVSwvnuIQEM8OkCxk3z

//pragma protect end_data_block
//pragma protect digest_block
gaO4nc/XFYqiwN7mLSx82TLn60E=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Read
 */

class svt_chi_read_followed_by_read_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yotRlLzwHypftd2pz2tZ57vZdJsLuvIN49ruXgbqUJgDBg54wTIzHrHUJFGf/wxp
5LHC0pqdHtYFkRFBlTVc/L7MjSnAOMSjIffzM2zXyEHhwMa5asWZ84xP13aCFpSi
3Rzw1II0xsuccQBgXZ1AZHeiUIGmx1qqjFtvcOV7hAW6DxMsCP2lYg==
//pragma protect end_key_block
//pragma protect digest_block
YXpya0Mi6ydQlpv/esec2fzn+nk=
//pragma protect end_digest_block
//pragma protect data_block
BgHXHHNEBV3ePvEaLQ/55G7qwHxUtuxx8K/Arp78SKwbLeyJZA6J3O2lQJWrhL1x
YfA0VKADLl05yEqqANy4AfQWyUyfdolUSvMBnfHVZg9F0MeyJ9N7CrYyG+Tj+tci
XdQgUy10oBDW/Ga8Tx4LPpfCZZrU6fsb4RMToQDvftUxbNP3V8oqwr1homb4NR1M
aUKoYswFuUUjCrXk77GP7QDCGSGS6Ehj4Q+QdaA1yxfjlTfa71q8aM7WzC5fg6Zd
TMPB2At20zshlR9/gvcUpH6ElfP44rolYuMTN8XsH7tiWOHHwf9kidkl7keEPjOD
I3Q5iHWE2MKktK80x4WiuZojFO44BV8KVPZ4oLVRQxyzIW9fBn0/Qis6XhItk5o0
U9oivImziuahcQsXqtWFfXWZEZiEmUG58dZNOtkVdmOWJPE9WDeOjAHhXPlCtKI9
e2GuqofnBS78LL76/CuoKDlN8uIoXDjUnIErDkCF/EzmJPoht6XV09RztFEwyMVS
f7dXKixn6RCzn86zJumN3VKdMeMrzPqDFxj+abGHonwLLDDOIGNXb96azb/RiJiC
Z1g4412z6bPjjyfQNXqV4yNyOrM4ocsjwIF9EnjKJqTOqjtmAwpx49HZ7qO5fsJp
v2AoFkioU9R5T+LMvwKgwP9MefNhtezd9dbQuqXOFhXUZ8d9Wjg+kk/+ILiKEgEy
pE+5mGCmUBjfg1mn1OtimFYvOOYDwl+D/ViNpKfyIciz1hQNXmR6SACXI40cCNdh
bfnRCsqtUBO5IuM/c8uF5aZxvFDUhYFh0jMV/97QjgI=
//pragma protect end_data_block
//pragma protect digest_block
tsoNEytID+2LISuZVU1ZLbBCsiE=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Read followed by Write
 */

class svt_chi_read_followed_by_write_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TBVhJFK+kbFbutiwkb3nWIrAgO4GDIOJVolM3WmzI1ooxOxrq0/ahRzCJWvgqgeb
2qmI/r5xIwZ42r9CRk/M8JEmV4UuX+UUiYzv8VuzlGZtL2n1WWXSlck0uhtzh7Hu
VcK+3FqzdukTuctpqWIITdHbgSpbq8pcre6oggz2k6f7EzwUUdf2Ug==
//pragma protect end_key_block
//pragma protect digest_block
0AatXhbbPLZ4MPK2UgWTUy1ND3w=
//pragma protect end_digest_block
//pragma protect data_block
LhRiGwzEkFE/MLZDzFPjCeiAwaWEPcxoqmpPtPrKXW3YbifL8XAFo+cEIUkbmrQg
4NYDMzhaNpL3RffbmOikfUHUD06iThZTWK77/aocBCrFdbPcASW0p9xOq+5SsWQl
aA3MnEA6G8QAqVwQLqynSzJ7R1h0Vui+VmaUg16Ic74DYTfvdYD3OpRDiyNLVUgP
DiqOgiJ/rVHps2uJLwJkMb7QtO7UYasw32uiUkNiCBQBLHyuviNVzdpecc2G3GpI
l9wEk1MFmxj4jBf9v+iH+PdL9zc8Df2iaRi728H5ifgxjURO8kY5NShzeogxhKEj
yTobN+2bqx7tawvutN6iktVSoVTG9atqlLYrZNNIItIn4C3djCivkLaQTN6yb+tj
hgO7ZkSQHf1YSbeWk7bXAYMP6U+vD1cTUd75OQumMyPbHbMt7gm39/LTnkfzW3/K
cVIXUHXDG/u/RpdKFb2j+YefeW10isPc6Z2zwLTiX5o2RruHTj1N8EvWMCIyYwK4
zI+zF+ErfWhWtx3hI5OD+sy4wZODDeL1y2hV6TV75gZIgmj8LWq7gcg6hR6NaJl6
udfMvVDEdJbNX80CE0XYLm+V7GLn31tWueNCAnHRVOI+Wsj9F0BElWCzLoLCZO2M
vgf4OH3KCW9sT6psd86kbFPR8IHL2H5wf5V2uRwBnWQ2xA9Vg3OVZPKI8KY6SlTx
BljwG4n1/q0X1q1on16+EYBQT+rlsQd0qTvj2Qe2lVjlzUknJ5XK/LW7sBdnKk8b
6SDMIzxMfE2WRUFJ7z9DnFBCU8oMWXD/chlaO0HP1VPA5wYcPtl6st70CnMYM9+u

//pragma protect end_data_block
//pragma protect digest_block
g+NIGrPks4/E9yKIDaG8sCBLzNw=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back Order Type Transaction
 */

class svt_chi_back2back_order_type_pattern_sequence extends svt_pattern_sequence;
  extern function new(int  pttrn_seq_id = -1, int unsigned  n_times, svt_chi_transaction::order_type_enum  order_type, bit  match=1'b1);
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
S6Zgkvid2sAPUxrImQHcthO6CEf9yLGKLVNEsPjQavMByBQTGfqNcICbWFir9YUQ
0sSZ963WWpqjlrQF6W6oZAoljTQXQNeUkcNBr5gr25V1Ae4a+oIo+RvDHoaQ7Tpg
kJs0LwKSethdImi76eITnqdOkndCeT/fUv0zhfbouBgQBg/16eJ45g==
//pragma protect end_key_block
//pragma protect digest_block
3y5tuHiuVVM4AJEz2nDyKxzSQXM=
//pragma protect end_digest_block
//pragma protect data_block
FltlBZqK6U1Vq4Q0RJog64RnVTK8cUhKKOefl+aYuJQ0zckNVTM8xNgIRRAmcIMC
MA2fGxT+YqM4BcjQHhsRrrCMxl7c/rqGbl6Kkznl/fRr8Yml3CA1rLs3yE1QKNTa
LAnI2Ybgo+rXFeqp6d8Jf+3bnx62dJ2Jo7cNa77XUz9JEvOsJO60BH1STr3eb84M
VAkpPoq4BdBaut793B228wakGYUJO2I8hMYW17mrfCzFx6JWy6ZwDnFj/oqBJPMP
IYPhbjzkmoTb3L9PCYbS25XcQZiViIHrI74oUbHUxop/N5mWSWe3kARQouynRLCR
ZeiZ7hwim+c/p+17b5vF5uq//Dehl+A+DbKrm2226V5Lb2XvwLdFyOzbyT1IruBA
tQ8lph0WJWQVicTLY8McvoetOPpR5vAd0Bkdq7wgY0b2qHM/wPJjAspbQJIgPdri
EvFi3twM6U/iIrmIHAbPGmPaetxTC8jxGAi1KfTTbraANOHHHM5T3cl1O6kHr/oi
nlKQAxINAarrPK0MniDkzjAJUyiEVnE86mi9AXVZb7RYMtDaSBfYctrmVy4QblnN
djHUIGiHGQskoKyRZfLR/pN0ANAnHzweG3YXYdTWZSfG05y5gNz+p7pfA9DZipia
wnJEHLnDJwJ2jkz9oVVTqoPZjpQjWtO/jbGoCTJ8g2mCHbZrH06+a8CSSMJAS18C
C/gfCN5TISVg2Il6GKwk9QRHKRBgMseH+WcTLcTapc/hwt2hU0WY9WUGl0TSYJTK
+7tDisG8c+BKOR9DWB8qC8XXQl6cM6ogNzQHUEJbEU5J1fZPPHqxL0dPMMGFQ8QC
U4gs3sWtmMTL38b7TgAvIAAkKeqH5DbERojqc7Zr3whh9xzJUov8foSOATUNfMuJ
FXxakOFKr4UKuUK2ak1iMYck2vhM6psbIvjN5uswZBJJazA1cgtedmIYJSQZNyJC
1XzRsx1XTNEC9nrV/DX4qI0nMcfPYnM30RoDg5J3msyOQGGfVlZtIGkcuehx0q3q
LxnHBvJkqEE2KxeED8CmQ+ojpu5EvAcIc4uL7sXlf8znjlvlnBCaQ0q65BsVT75T
caITz2isAkNLvr6q7t3JtXtEXajNDvnLOTE1ymBQD/vvyBG4375L3PKdSwFgE+vj
kBO6Q1ejPb1weg30WItSldER7h4nUohlxZJve6ZkdXK50sciABHIndTA2KgRg+P3
piGXKd3OFE99W+k9drlFLd5wVLDLm7AAQiwGn3QRFXo=
//pragma protect end_data_block
//pragma protect digest_block
R66fvOZOsTHgtdviqcSN2pRKt74=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Non No-Ordering Order Write/Read followed by Non No-Ordering Order Write/Read followed by No-Ordering Read
 * with Same Address/Different-Different Address.
 *
 * i.e. '1. Request/Endpoint Order WR/RD[Same Addr]  ------->  2. Request/Endpoint Order WR/RD[Same Addr]  ------->  3. No Ordering RD[Same Addr]'
 * i.e. '1. Request/Endpoint Order WR/RD[Diff Addr]  ------->  2. Request/Endpoint Order WR/RD[Diff Addr]  ------->  3. No Ordering RD[Diff Addr]'
 */

class svt_chi_no_ordering_rd_after_two_non_no_ordering_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6rs/LFCTc9smpTY7JNmYYUhG7U9EF+7+pl0++XdWIwTCvX/JSHr47A9JjFIofcQK
OM0nSYJekjoC2y0XHGELlhz24jJCNmCbEFlMuR4NkpFmV+R3eYwz4d4DQtruhXEY
WEz4eFr22N1zbDJLUV3WwS7j5uX8/TfLW8dBcmkGiabcXu+3W805+g==
//pragma protect end_key_block
//pragma protect digest_block
syBVTQi8DbzduHei4+Sdy9TzxU4=
//pragma protect end_digest_block
//pragma protect data_block
qUqPjmugYgLkG+ZHwotnJRwLmrdXhixJ/s4wUQ5LJskP+oVtxzfK/0c5hQRuB8Lk
5ghHbNBM/5vuv2Szjcra9bAR0ImkJO1eEchjP0sEQKsArbM7eO7AIMu7dbQM2N1x
4HlzmhEtRnCXQHpv3siggeu2Hi5Su/x83ovLnrkoQxEm9OWM+tBUUFFT8Vw/WLBu
+9n2yNEdB23ncgCHMP3zgRVBt+sy52pVfq88xBkIl8raqhCE4NciGX1xAxAvEZAq
6bzYCb2ql0wNZZYdFLyMArW1oMXIqSrceYiiL85W+9wX5TjrEGpBNuKHFhdLTM31
I+YfAe05aMfFvRu2E08a91AWTYLYRLIH+OF1tjlHnFONv7O1LL4ZVAq3HqFFSs+m
2soOUdjeo5KJZmIJ/6qDTN/EGg9lNZfI+RbUAcN1slR3NNAJGyqwTQr3cwJ55Nje
NTNQIIMeyET5Wj1U3u3NK30cEk7n0nZzB1Rbbf9V6hh43qjQAxFkreuVM7g4Pc0l
rDI9zJWOOKv3mzQrX8ZG3TigSDEzuFLyHsVerpXpkppppWVRk+IMASHoe53AEnrg
DkbLGebkmz1ERvRe7IxiDACTeoEe05seMx0+ZIVYMFn+M/BhlYgG2sX8Wsfh9l/Z
eTpgJ7f26uXPmFLmYSJz0bc7ziNkN/XeBN506sx0M7/31vVJlBAn9+3sb0ur5tuc
6G7fHD7mpBdZQlhDzuLcnvejQdUEXIOqO9PDLdQk3d34ZEM7kOp6+7BsQrEsjFhf
buRz/IgvNTaJN9hAr2P6Bn4m1Urw5vWt7QfRQVw5qNv3vQ723JOsmi+4ad5aGDpT
c+4nPtKX11XvBeEiWMwEfPRLTB1HWQdts2lC7OkmHha4aU+ykujk8M4AAuRQpGhS
B7DviDGySYSwbq0MDUAegKHdgpgTuXwlQ6qKvzvA7J0vwfS6GUJksiJqXq1jsVKv
JspWg0uaILs+e64J7yBcutbsCK2azPRiKebqri+wpxonUrB5592TTvrqoEF7dNVV
B2ADV2SkSHlEdaK349vP3rCNjeZ0ArSrWkurhYo8CakRVPN4T+uw6G50jmKVlFot
I1mpiROGSsKtoZweWQUvH68iS1NNYj1q6JaE56mvlgAyRgMpoBMGxCS5yznHBitx
Mcj41pVNLhJVVQzCapfYOlK/+Lk3qxDiPPQVLS6NxkPMZEvcN9outrqGti+CgQil
tHVilS71CPgtOIdboQ7Hl3fm8MwVWFyfba6Fa14/aqw=
//pragma protect end_data_block
//pragma protect digest_block
08EBYkVuURqUT+wFr7nq2favF/Q=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * 'N' times Back2Back CHI Transactions of Same Source-ID
 */

class svt_chi_back2back_transaction_same_src_id_pattern_sequence extends svt_pattern_sequence;
  extern function new(svt_chi_node_configuration  cfg, int  pttrn_seq_id = -1, int unsigned  n_times);
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HtSHSK6AFEQUNsX78YI5zcNFvIqx6w2BgFmYXGnhEb3bR6xTI/lEy6vYQ7ekd9Ks
CAbfXJzRC9NNN6hYSWttzAT0mfom0cE6KfEu/XfNNTGME0rdOTOESMMmacGgqNIb
SQUGKxXYvP7Opiigg/ofPJcRuKwNlYE986Fcv/wbMDXOmPi+hKE/Ag==
//pragma protect end_key_block
//pragma protect digest_block
5IGji20NJtPCm0gYK5Wx/E+BQLw=
//pragma protect end_digest_block
//pragma protect data_block
WVSli8IKl7PZNUx3CNNrHDfir8oFdMxKOKoKFcfxF2ar003f1PILBLzlJUW2Ici2
pKWdKD6Oj/YsPFIhAfYdv/U1pPsp5f0gaKl1OS85u9fnGv61ZN3KMjaMP+Cwqvra
LpwN5ATgmowt4ANk8thgPitYIEOCE6DdtE7FQ0dolADqvqseYu61VNCL0Xn76hyi
LpkFQOu6W1Hr1TBQ5h7O1XUliUqCoAVJQvdfyZHjl8gqjvqh96oWIAOErLfoZsGJ
gpsx2dSzmQSqq3yGE/73fhSTsTLF0fsN4Kcq8y0qBmZII/OYIMOrgHLDAhwH652D
+abnAO7+zxESLW2LALQMomhtA0W3ofbuz9PjulYm0C4xQUBHVcY6C9OHIQbkuPbP
ZnmfiNqDKklZ8ezccTsDRAiSsxrtImnWJ3JybXv9sa45oFWL5vSvPUyAebjAOa5l
CzgPYdSC6JuY7zPbdDsF7S2xA/knn3NwplX/9Qd49eMmbz1DHo+iQ7FosCt9/iSq
6+hG9zErNR4pmsJWYe9nn3Npsc7WOabbpSZGqjgrs0PyQvLGSchTazCacnrLOYDR
d4j4dpwzZe8JzvG4osDt4eNiBH+S+xaM8yJKeCSceEw4PTHhL5tkOaxFNPD5eD9C
gKHeamh2vNp2tzHFYX6S/6AjJROgO0RLD8CzZfvQ5m/ZvkWCu+HAFnM0DBeW8fRs
1KY/yMEfrZRJUGK4ccTlkFgYSo7sGEWaAuDxfzVPE9cEtl821iCudXWmqHQhge8g
fqO/uD5dkDIMAaEFZU8EVvRiOn5omfPRNKmNso6XlBZ/JlbXalAdlYkiz4rzKAa/
5UHReArYNlpuXO10ivnzO76mdti+kyHBkXglLfubIM8xkcMpmfAePDdsS3qFWO7q
KmJOqob+VNkZhxisZ+WLNq7TNPgYv6wXsQv17Lr0J0FqAEy8gjx3EEqwNuxd4687
nRFPrhtVODBRjmcFqIV8pOl8c6XueZ39n0Djg8J8gxVKWDq424b+t5axUqYvBgPk
edhYx09ZVkYFWLWSywpSvaqAhmN7ryPILxGwM708+92xpCOQ/VBrKhOhzFYt4/oH
pWVe4+dkHTkLqz8A45rDnvbCVYtZSbuScudlIZdmI9hQlm81/ZndIkOB5W/LFJhG
ZqQlizYX42RMfTLz/SJzzKmJSsnLGNWgfn6wnYiXE54FIzXenzQ0r2VomgvGlWHq
jRBmUmm7Q84grAfOmNNzkuBMfxIcZs9buiBIPU/aj0fDTQB0ulHacwG12qVQ48dj
ih+/X140RG6KPQy+GU0tpWEImrgPkrK+SHzX+YLurKW+6KvFzIAsTvXKLxaLt8QH
HmqCS+jXZAKGuogvQ6MqXT2TXOEcXcYsLDe1z6Jlm0OJZnvZggKDiTbLGCb7G6QK
Rt0qga3OdpHowKmbzODJ+0VjDA9W8lBkbs0q46sWFPp5ArkZQvDcyu6yYjMsZi8w
n2JXSfr0eHKyuhE5aDBi7gWV/x+UmbM1kFLzPp5kAdw=
//pragma protect end_data_block
//pragma protect digest_block
Eduw8XdITP0BSwJeOHvc+w5+L4k=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * CHI-B Spec Figure 2-23::Three Read Request Order Example
 * Ordered READ#1 ---> Ordered READ#2 ---> Retry Ordered READ#2 ---> Ordered READ#3
 */

class svt_chi_three_read_request_ordering_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UxbW1k49dKmSLUGfRYTu2SnM16HffaCUM0+W6L+Od6W2wcuFBBhjjMB0TZ2eEkzc
QFmlq8cHCpUZDqoOnrMwBBeAPKjrFvckuFo0kQf1QMluiaYlcDZditKmOrrp9cNO
k08JNT7HZjeMg6hT36hbPmkSW8Rowklxdba/2yjB+ICmoQsLoafuow==
//pragma protect end_key_block
//pragma protect digest_block
wGT4JQXHfLAQk3LKf6j1kjst7VQ=
//pragma protect end_digest_block
//pragma protect data_block
4+w8DX5PNAveUYj6JyxHr8RRyVGI4FO4ZhPIFpvLJUUAcTVC/jV6qBnattp4Icxb
B+/5PmPJfbhbdtC49jTWCVzbKUYsNZnb+RTDeF0L9jJlIJc/44Y3Hl6Hr8bnDBDI
shKfBPusBS8BW5M9MrXQi6KvawLynHXJTNAhSaB0Py3b7hX1n0FewQLdgRK7Hc8h
MVFS4EcCi6DQwX0zcukCwNx+G3N0Dl/mp3Kna/wtthhQz5mNDfFL0DX0YSuS9aYb
pPoBef0nkbG8MeYd7FZxeHlsDIJTB75jZQc+pOLfxhUBkgJPxrBZQLL6WGgXgpHo
KWX+eAy1g0cy3zRanlUF5b1DrL0FF9BkAVBoaYdO2zm32ML/cd9KKKpuLG4BNanE
I5v5XXIgRVbfP7oYp5MrCUNrWvnqtOVBwKOBJJIe7oGAukoFQUQpclXpoOKfhtot
wg+qbZUe12WLKW+7ac0KM89bwzLcRIMclNEoTtvz/Jy6bnV65CGkaOM7tYC4WRqx
eBIYzHxTMyoNSVy3oN3wWfJvYEDEXJdHisYtXNz0GnWboH+2N5D6jtcOh4Cvzirj
aXJ1lL4JmLtJrR25eCo/1Mo+LGKLQZ+ENbVUd7sr6MqC1Q4jKGCkVkLqvdbGEvms
sT29gfaDs2G2mqn/N3hc6S1RWx2SsZq63SDF5AKuJKHMFcwEZYHMnxp7wWp9UsqI
drRRcfUIN3keSJa3OlTnkZeMBRL7dw9QFvwzVxY21Fi/PmnFu+XO7C7cDo2rbQ8l
oC2xr8gW2I+Pn6u5AEuKrhyLwfO+VGxplFM7AmJNiTCjuhhzzHFoAGufhTSKXPza
4bpWCQB4lkwNxALDL2cE3P/z9MG74FdEO+1yRjafdXE13nzIqsyd+xzhhO9J8V2u
unsYdXho9xwyFElRKWsuBg6hf0O0xWr8n27AHfAuZjbqpFm6THjZkJ19+KAb0dru
SvQl9/GmWF4Yfe1lxi+jOpZsn+Ulk0aOK4Z0qyDXCEprBX6g7lDd9yoMQr7jvxYp
rLLLnKbegokuOl4XVEC/ywyppko93I9wusS7syNrQu0SwhgsOYSz4e9Ibca/blFT
+Qe41aQRjEQzKJpxgJhdTJ9tP6yeYWENpPjF/87MFE1tCQfvk3RLuBMqsNi282Yk
npqLJib2E898U8n/ayRL9WMThLZe9mnKvNEva5PBvJl1qlvlHQytCqxmeHoQGUJs
sgKTaCzXUY0Ok2krgnV3jzcMwtr731LiJVbyN70X9swT9j/v+n8f2IugimZ9NEtn
veBHE0OYKXWNtxc8bSdBD2oZunb7WSGGaGOIOTFY/Do+6CXymxA/rK/aXUqxr3NN
5XXWEeURayqx7DM8k4rn2tylGqqq9opeY9PibFx6EyE4Y9OqLXym2WdgbQsDJgnP
RMLnMoa+Y/VRpNil1SphZphM4kwXp6kx+4wMsJ2gyXHn6ZYHp22/WE3AP44FkE+F
EyFrh+DTBRnUC9MrFvW+YuWtf03fFeTfbdxTHFpQWaKzIP8KkjGf+w1D29HfV7te
F+MUjwchcOE0GxKZaguwr5+am0eneTeYdAW3Fp/+sx753KdaOSsec66OoWeFuiwm
fjnuTIoU+wd0Rq+0mgXji7URcxNMEomP++dwG4GegoCzAa/JHHKrXr2bP8sVhlTJ
IVVcYNrJ6f+UlBLu1xb6rD+mvkTzt02poAaW2KrjFJ6IXFZDS/7BTXXjggi6d6ii
pgPrMNGsuYV38AtCG9vCHa3riGQI87elVqbMm+uBc5o/lSVOnYkVMKseAOINBEeJ

//pragma protect end_data_block
//pragma protect digest_block
VM3f4Ej3BGXe24fbkb2hFCPzkHc=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8kcqoLFLbsflRRZL30tjUXYDA9mm1054Fleq8G8oYPeXXPaZ3msshf/IwzLJQ6t8
3wR0lXgjjgjSnC2o7UwdCkgwyYy7DVW1Mvz6msRmz9m8jWpui9HWOWty1HfbiP3U
pUyZkloXkJPhdqLJxGd8umgsiCVHfvYlcts3/KONT1B4y0vD4gEt0A==
//pragma protect end_key_block
//pragma protect digest_block
FtvH0qfZGogtxYH07nCY1pZKD4k=
//pragma protect end_digest_block
//pragma protect data_block
3/5l2A7YwVPoAOggUfFYErbICP8Zbhi5Lx27cJWw2bCl6hwPXuci//ecpbLl9Rvk
e4ZAoQZ6cHeIWbmk95emdoWd+7ops4C/rR9GOu/CD31Kn6DZZA7qKzyRAXLmzfJZ
Gmf0+bxQ8+fFKKzCBW94AyNExRaAZ8uj/IVi4lc+qC/+6BQyxPXRXCQhsOec/ifH
TFyF2Hl6T5suUAS6tolJ0X+94RFbYrSzJidbU9aa7WIl9ubPrq4q4ng6aGUcaEZG
Mnl/71xOYAOtvT31/U1ioLfV3nZiiptsYogY8Qvs48H8kEBl8g9iosWbG+0eNhX5
WhJKCD8/6T9cmsLFMt2SajEf3b0+IqP+gC3jqy4cFIUqf/Ii5PETpCi9Ys3TcOX0
Y8VRifXdRhQlEco+zh3IXyYfO8VJj+Obfe8S4BJqtvwjODh06EeIy3cZH2Ay2OEx
670vbgvCh3wWxYU35mOfIl+tmC7Y8M0FlRi6oGJKUg+XMeKIyHIsRm6s9499K54b
p6EDHg4LIpJ0bspzgv1VNYXBeOvdXQRlfACfls1dT7hMAwMiSbeae/NxC6SySdFV
bQsDnjGqeIZL8lY6E4Nwfq0wsAa2gK/lQ8RlsA6MJNqPVysTBbcSa43TjIzIWuWa
hm80pwSCQGifEq1VB4wWd6t2PGuiakUShhMeSISbrzDAipUhTii+uiLUIXKfHTF8
S0AC/jzzbP0R8xxG9yMIew+GPlwVFFnINV5w6OjVHaypd+HQw+w8dE+gV8xOoRcJ
oul6jODMp1rqkyUxINYf49lVRxqpctjXxTSQe0vBnvwFCRdVlzcBTD+CY0ytiznc
A+zhz3WD4kdl7wlgVQf2RQGAkfZOrfcLOLuYb/Vvu6BMjSINTvtsUXxmUVhGOBQ6
t5kDV7XNIhKC6DbWaW9oBL2hBSQIcPII9F5oOJ1hIfu6gfCAcM7if6QpdyT04smc
PwO5ZMIrd2+Z46LytM3GWw==
//pragma protect end_data_block
//pragma protect digest_block
/qMTtth4Udx0V5s8ehVyhmJI+kg=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Cancelled Transaction of #1 on Retry Request ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_cancel_transaction_between_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SD8trsPHo8t5tMz9TMmxp/I3E1UqT5ipicUkqABc9dgcF+ibbK03vz8U8mzdOleF
S/AcPW2dR6tf2eVX1Tv0zn5sWjGOsfSIq6OOtkOmdP8WhF5UhgIPx26Wza3CYwq1
qg3bUEfct0DF/YVDvK/NT1JlMe0DrmVqDVaGxn9zT9ylTaQ4Ih4/KQ==
//pragma protect end_key_block
//pragma protect digest_block
c1DfbMtBSoSzXdj8Kk1QF0XRAGI=
//pragma protect end_digest_block
//pragma protect data_block
PyH32otUIU+rx4Qvmc/OW4JeNWm8WMdX6JdqKxrggMW0VTT0rd21Wecup6V/Z6B1
KFu8NMJ5syVq8of8RN8wF6UmEV34Sm8u2DMxjXaVRI4PDZCQIBK0+u0lo5QWn5wH
uSB8Bju9yi7ksm9aA7e01oDxY+2nwtfl9ZXVRDMIlu5FP8W8AiOvfjmJP6WHp8nT
ByalMWoicPi+71sjds1UZXIHA4hbhF0dnwyHDMUtDzvqaABoYa9qbt/Yl6Iijilc
I7ucXUbuvMH61nQ9sQoBe/L1+JDocJ6OU485PleH/xz7pUsu+9KG/ULgK6RgfKNa
J7H60caA7NGkskEU5wumjU62L/Jy0b9Lh/XpdlpyXqg/y6xln8l8RByTCSDIGCle
ir6CE1GERggRXcrAdIPevYgeqAzSZZ1elg7J0KwXWNT5UfeSEHhrFqGtTU6nt3q8
9Fps2MewIHRp8F6cUOVurMLV2VP/5mkzTIeyQ1j9lAwQcm+lWtj1WLE+WutRh5tT
8yiK8yEex/3V5+RSGa3cJ+Z/am3ytDpPMLbrQPkp1QLXWjKh7Sqw9j3PXDUR5fE1
kAIYSZCYZE8LRiTXcG1Xr2X6UuRWs1f10xuIQEztdM3TB6D1yJR3H/AhJVFfMjbD
vo3gqkk9N/1ST3wAgulnrpFKQ2Q1ZINomhSyuiFx/vwBNXWoh/feCaMmLZqlSNso
XA6x5G2cHydAJ2GgtDhLmhXqNrsPpHwvvkEFozZ+8lvqzBy+FkEXB/WJpqozKQwZ
DAWyVMdSykpU+KSrWtrXN0V0YxISXVv9YBl6UL6uaqPISnfmvUbyKjtgDjDcbqRd
4c4CCitPSu9gcIZQooG/qyzOd3Pw5r3BSAwsWtivn9J3bn5++773BVYYIw8/2PKq
LTH2QZgDTSsbye3s9t7wie9tIad6Yc5rsdrmOSEtvnHaRH7xfXYvjCMsqxDsx7dF
mj14el/jBAx7KCcFyp2zqIKBaSbMjvZuJRBt6DHHuvqOZtpHGWud6Qfx9EtbgfXr
eltY7KdugdC0xIijgYpGOA==
//pragma protect end_data_block
//pragma protect digest_block
EIgeBJpz23BfGoi5CIjPmO3C9Sg=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Retried Transaction of #1 with same/different TxnID of #1 ---> Any Normal CHI Transaction#2 with same TxnID of #1
 */

class svt_chi_retry_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
3tIZIfFcz8BH0Wtj6i8lA/tmD2YADZFGDgacizJFg/0wOQbGazF2hG4qFl2NQl8M
b3WSE5CpScvvaAlr7KCk3/mcaIJKoYjqL5cWDmBFXfFe+FfX6gNDcgUCQA92LTTo
hWdYEUKb8hgncginXxReoY9FrbihCNDtkEJ3REe1hu88RcgZkFHHKg==
//pragma protect end_key_block
//pragma protect digest_block
IeNwyUcvVjOhxWz01wihbSfviGk=
//pragma protect end_digest_block
//pragma protect data_block
3iw/DSpGv3rFru0zYf0F63rCEIVKxqy3o6CXonuVHp6tHGjRIs7fmin8CzaeXedg
SVpxvypCZRcTUAVZ3q5+oTZXzvTzof9g7i321lIRGYUVVWOQicxvrXHX+7g2+zy6
B93ecKHms4uEEsOzA8/mfXH9yJJYz+Cy29zI3gBfR+LU9pYmh5ImklbBDomLdjox
FpuJ4EeX1iEA2yCYdJI5ZceIgDFCgnSTfxQwf5IKlWXTGBOk4E+MEnU6v3OG5KP1
pfPOXuDkNP1Rlcm2SDgwqZSik0Kg90lLPlbR1XaOxwRXvpkHdzjnJSXw+tr+7c1N
IKd61xfCvecrO9Vmf7LMUzTJl8EK7QeL8HAU9KhGpTxNA25VJf6AXNX+d7roWlj7
tDf30BaMX2naB1tlguUKC8qnBHMrebtc9TMhgZ+y+n0i0EutCqqkF6gjNdEXkpSg
jS7SAkTvJglAseOqILjFG+9+Cb0cI1QauDzMdKgKi1LLRXUmg96cRHZbOreKkumj
cU64YRy9pLfwoRNsQ44tHWsfIzEgJSUaEziDheActE8Ql9DEe0yUD7GvWTxeUtwc
Jmd46CEeFqI7wqSPRdzi8yfqaMJI/qULTj9yRn5RPAjJnTjn744DXM1jGAM8NOrn
stQaQE2D2GpiAucV73+6Hri2vXyQpNk8qTgQ7D5+m2MpE8nxZAflERC3e2z7jNGX
caMntsCxaBXTwTFsbOUOrbnlBbcVnoSpolWeKSZot/rbvDBdZbgfo+JUHwFZluyQ
YQRpkVM6iIC/oYaZRs5GkpLTJ2JKdEaP+J2k83xPmL/e7CGdJSjmXKES3/iuA22/
4dntvacK+fuE7MDSwikl8S5moddMjQIlqjAklU60lEhHikyXd9WySKhtWPW6FtJI
XFqAq7B2Ji6/SFsb6F+Cui+kyuGjoUutVZnlot0nBQzDOQ8hPfgUc6HXu7yaPY2x

//pragma protect end_data_block
//pragma protect digest_block
GqWKW+rSKqSrki6sqoUunQPnojw=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     Any Normal CHI Transaction#1 ---> Any Normal CHI Transaction#2 with same TxnID of #1 ---> Cancelled Transaction of #1 on Retry Request
 */

class svt_chi_cancel_transaction_after_two_normal_transaction_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
r5oOdpae8ZJp9VkuLoURY7AIppy3l8sHGih0kwWWW6g2XKZpD0KD/wXSL6Rvhvn8
19x/nxpWI7veWCv4+Zio4Z9e4skK1yXA39de80UQCK8WMPApiaarMn+uXaCbNAs9
7nF2eiybolTbLqOYwd8Z+CERMxktcUIxOf0DDQZiLTPUF6GnG4HLgw==
//pragma protect end_key_block
//pragma protect digest_block
c0s5jL++f12KuBxvCWMyRyhr/XU=
//pragma protect end_digest_block
//pragma protect data_block
DRu9sTBIpETm+zKxCxV8OCr0B8ymBI0AE+NGYJaMq7MLgJ4kGvJafzJk97Mmb7we
6qO34iov00cGZ+L//GDuhbPPApdrrev8oxoTwQrPUe5F+WUAFh1OY88GWLcQaOmw
YTl/IzCUC6j8sDdZlEGkvrQZW9LypxZugSIit9Kp6a2fSYjXeYi/xH8YMUyAy3QU
unja2j09+HSG/BGji2FbSSTvCSnKeKR9tx2wj9YO0wiMWdMD/M2rq2+2yasDxykM
Fy5F1yO+KTxf7VE5RcRp/mNrSEAtM49PoSVh+qTMhwgNU9a7oB3c6Y+zaD6Xz+Vk
N5rWZdOALeShxnpa3I3/DEdutswQmQkLxD/EUjwa2sZNLghB74XW19leAOqmv/Zr
gCX/MpzChC/KD/12rIH5fiZCGZ1hTxx+IYG1j4kn11Vtb9GpY6+S5XCxZ/OUwZQM
cLm8l+z4hnG8ExIQfvyx8Od+q5PmEAJoaeJFPR37qPEX+P6zh1+acuHib/i+urfV
OFWJF005M+3zFYAJnq1YI80Uzm/Toq1C4ZwuvQj4/jI/KhFC/ny2EskZbEXAHipo
CKnFZlaMFdLEY5B53AJNJP1vrbCcIT12uW/+hjdLr2+zwF6fYNCjgB4J9ir7HvBd
ml+e/O8Ix4Jex2KyXSBuox+UUQzbzXnne28ldJ57RcktwcXIyfHhtlyDQa7rlTMn
pAizkh72+uJylMFH2bW5HHTLS6j69R/Jlwes28G5aC7lYOHHY0WxtbbtjCYuItPr
fuDkMFNLgiDelQ+H+6YE+Qd5go0fHnt4G+l0zol12Agz4ulp67E152WMBv94HEEL
w4TGw/lOoHnjNAknIMuD1Tyv6vZNKOh17HYc9TXxtNSveOgjEqJ7YhTIQr6ZSVOH
CIKCnWyYK4Ar8vOI5i6xsXNS3L3ihJXgmYNNMxXSKTMKu1vXofS+4vokmp3wGkF1
x0Juv/vuBh2ehVyMrb0A70e8AMpSiXJIs7Sz8lPMMzOb+1CRecXwdq+tzDjf7d9c
uT26OW+/kbElMCSFrVug8A==
//pragma protect end_data_block
//pragma protect digest_block
LFvKz0geEvcVyxI4yQ8JbZl9oIY=
//pragma protect end_digest_block
//pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
W22ya+CDHyzAqjETq3Kg/BUrRopkVPVh4TsDY2YWV7ps7CxkXf16VI+vdWPuzGf1
tdaYZBqa+SyPWr6sntgRahxxf0mGxkZTf0cqUKz6xatGcEAdlHzo7Rpg4BHi7BTk
qs3SWtUIFJ23gpvTnLnaU1pUx9eUNry80fSpDE6SGjr3XMMr+d9tAg==
//pragma protect end_key_block
//pragma protect digest_block
EHF6jEHYKuo+hTvhcP152hA1UKY=
//pragma protect end_digest_block
//pragma protect data_block
LKOa9ib3jAU6wzundzaAYZJsg8LUnVBgbYSLCglZmRuy2Je4HL/wGSOg8numkX5n
g2ly9kO7CwA3xHm9Ft0+g3ELkWLqdHoO2FWoHpFbBFw6VQzzueolPSxZreDudkcP
BfbR6D9UZN6alW1B2+dmIycb37Vn64Z1WXuhJdwlFVS3p59GfOyJsuZwrBt5u4Wn
luAll0AN3Hic4xtQ6W05NZ+zBd2afBBq4sPyN+5IQ+LhNg3kzRg+ABd+pyqBDdvT
33d0Z7VK3G2WPLh9BjT0kPHulckQ+lNyrE9Vc7ZsZIXiGPUE2JZK0IJwShsrOfSy
HMRbICNN6pGm9k7pOSmJp53Kcr5aua0r6aMa+EagmJepzdDU5ARyBLtmZXBSzNcQ
uev9zRGltPbFXSg/aq9no/dNCdvVn+RInUZKbV/U/w9IJN71bI/3ZpDH1/ZB3W6c
AeSdMwSokpq6ZS6Q6qYO94+rlKFBaH3o2vPvEHqaiLIqlJeNi056LW5c/6vlQ3Ru
DnEXTR/GgENVPILin3dy3HCvLkG7WwAius0zahcT8MzUN/ip8F1G15eLEeWzYkqC
R45WHkQWgsClmJ8Zt5aRMuNaNuvpNbOhjBjXJhYu0GR/tEto8853LewGzig/BKg8
9/L4uKzHDQXiI7h2mBC87/FHcQrbfXKDxW4ch3narLB6qDf+ydHgvHYupjfSsfRj
uYUs9UKu7780XCNPFR7Do0XzZ4KzwvovzLnb8fDulxqwr3xjCE4O4ZSvxykTumIH
b9Q2I8BAaeACpF8nudkmxdHskXIvDQTQhuHRelpfYZaJU+5dt2sNWk5SGIK37elv
UmJIOnL6HWbXavaA6zlgBKajIDQoq0lnSiSwZt4CybNXYe2C5QICLf44UQqGm1BI
3CIP/OfTxtm4v9zWm6QaOK3CVxUEBuf5Wvsy619gDLS4rmkn8+7tOLjvJSn+jONH
o+kS97OZWVJpD46yHJSLDAPlSrCWLP+x24ZpmV6WQkB6SpJRTIPaI8+QpE/kolki
6/Fo6wtkhpYtwmhFbPDgdHefG8HZAinXbCiEa0i2/pTGHWB3EMXRMbPrKe29jKUJ

//pragma protect end_data_block
//pragma protect digest_block
DFUYKyrOfsm6HcNjzUlNHreoPhI=
//pragma protect end_digest_block
//pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp Sync followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_sync_followed_by_retry_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
q7sffPxLKGDY17DS7lVfz/k1gIMCUIoMkH9cHsyTIJc8PK4dzeHng6favIPd4QPg
ahPJidjlnO8ecXSn47IUfKmFZL1E23LzjzkRHchS7FiTNwl/THZhtft07qNCTJ+8
uPGlYZ+W4zMcIjEqj5PEMflbqATb3R//WmPOyNjKN4jpMbgv23U3Og==
//pragma protect end_key_block
//pragma protect digest_block
7l2RBeIa673QcW7ZOy/+PVYwwoI=
//pragma protect end_digest_block
//pragma protect data_block
4pnwJHQymYDcxjiNE7lP72irV7sGPdF3E2CQhzBgCMEX9nXCBc7tiIMlgP+5neCr
5NWZTo2x+PcAG3uOPPkIDcdLek/hpDlRu35lv+98wzYzDVvd7C0vaKAak/6bDLxB
+E1rnVpY/vC2F0VzhJd+OVprl0LCnibT71a2FpGnep2B8cv2UfaGiD9gw9GVaDN7
c0aUxgSD+wKfaIe6r+4c/xegIGa/n5OKRMVUf2JDc4HrgQYqztD0mn5IwGEr7OEx
yQPPZRp6g1241NiiKtXMxuEdp+pHaxHaSBG0UHXweSTDyHx/mb32hon83IWwOXAf
8QPdn/9w+yvNOk/UuxKWUqjBxZvNoZKkR8QOlk0k5HVpn/vAu5xqEuPHTrX6s2Tp
TG/7OXjuxegS2+JnqWQACG6+xlRRb8IMBtg83Dk2BWgFmDOto37aptcSqmYPXu0A
0/uBHt0Lkb/tblG+D19GIRkhHitrpKxz/o71dXqZVegBK2QdpDrwMDt3VyddcK7g
xIBdqCKA2P/pFqaA7Ch5lYpnEVy0bBFwZkbV0PHg8a0rAQt0lvJXoa/cd9rJA4H7
lOUHYisugAoan6HheDWyTVDrFEA4T1l4oda3RDc5djrZSqER8jQdlkmWNJhgwGT7
3VbXDlhNXG3dYjq2c1ntwDAD1GashAE08cJc0Z889AjR/sdFTZOA8GuJ+X37KKEA
56+88I3JMTGTQ1+BTFD+DlPsd83+L9zCgECRBvKqzn1HxyZSFdcSojqE1JUArV0z
1J2TQ46xFLf6EiixJQLq4hqaT2U1N4MZ2fJ9PI9y37cXM7Wr8N6WJSA6EdEw980r
zyGdJPLI+XbKdphsksz34jsesZLHPXWijKx/EKn0fh0VQz6YlCywcFGYyLZjAh0b
amlq00VeimwTc73MmYYQS8vVXTuGqRdKdsHKN2TY/S2l0fDdHYsqCMcWPgE4jnIL
XoEjvL+uROHsdLGNA1ALbnKLlbQP72EsMREIAoGyqPCDoBqdwNhwWKlIlzu9kkwf
zMHetdiiETJuG7CZ8xF8OeyHr4ChBeMhNCu3Jr4wW+2XUsi8a76ZVr/bZFPn7Qgv
X41FeF6Lf0ED9w5QEhzXCwv9ZjwAWbxx5EVzZJBfATzekA1sohrIxdkYp4EXWqUC
9tRIpKP6sNVNzn+OddJCDOEKxXqn9a9MksaMJkzfDwJN9OS9bT0o7D+G923MAEn6
495q68EgvCq35wyJJ5E3tbqt4DvB6xsVzv4aTabQszmksbz/aiz2esXjdx++iOJg

//pragma protect end_data_block
//pragma protect digest_block
FSEIfZ7uOv7TinM9/DXrCuxowGM=
//pragma protect end_digest_block
//pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI outstanding followed by DVMOp TLBI followed by Retry DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_outstanding_followed_by_dvmop_tlbi_followed_by_retry_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
i9L9k/hk5Qwr7cro7iCPckL55RMwfHXZvEs+EjdHJJkBQUzDiJUv8Em9baOzRJAL
i4qdNzUB1kUFt4FOeFtS4vWkjvFipFcesfwygFs+nv4HZn3MSDD0Z+X5+TZOPtZB
sjBl7YQVqDWf/vr08y9ni8P182wO92TtI0AELPJhPTEui2YF++IoIA==
//pragma protect end_key_block
//pragma protect digest_block
kfbfE2fDBFWqZ+2k1q/YdqmjzMU=
//pragma protect end_digest_block
//pragma protect data_block
GQPGgkmjrUIUTlYuaoqd7KnQMv+25+82ln1duzVJTFsx+3/NSh8tbjXplG4hmiFa
+QLHbjwhWzT4P4MfdGfmzlxGbJbGSev4UD/gUYCt4JsqwFlxJLmnmXvf2orOIF9g
NeNBetcfyKHpjXtrqEwwXh8Dp0i7lypRd5Ki2d3pe2kGNfWdGDl+JNxjCn2bw17T
JV6cxlWSsKmb//w+3KGzTYPUWS4PXFQh0BRKUeD9ZaPq667Gdnmz9tgNm2Iu5XuN
QqhmhCykKhJF/ZjSQU8b876iId3F4OWcKRwaYiGIB9QTHSxVZXrzQU2WPjtej27n
J/mpa4sDYzlKwOu9J1E64P4oj1nb3AT5TnTy8IhoMehKSzsdXSU7jCwxjQwtV5fR
1esRhwpjhEtnssF//TMAyKsLOWvdDP6Z64RB4z7m1k+MK4rgzoe2YcQpPgh2gevm
6yf2WIQFQ+vxW4bIafaonV+6Sm6AVZlY16zVD18muj/qdbkXUYZVrmKY2pHT+iF1
9DHB+/Y5vNLvmDOG9lIBEQXqqNqq1pidzhQ7ar4cFf6VLgLMEWHXHfpzUl1SFE66
KYvPE9yDYFKhg4Y1wBiL5rWS/cd5R6LqgoMNCWjhxh1nA4kE/YxzApCsm3O+dluM
aZY5QCx7jrwPSgENwUyYR/Gdv5LXRnKc3Bf2N0X7ueQYhtTVcCze82A3hfxTJmCr
plvSGCoaiRrZtMVcBSBTjCBjDtKAwHxQ62wYBAC7mYlkPoAApkdOMB8uN9SbqAFn
10SbjsMnz/Zwt+g31H6wWrYXFzVPLE+54IXQux6zABzrCxjWUtXGzROCSBruJzR6
JIhv9k/NmNcTs3+TtJcXeCQY+8BTNy8kodVMqKTaRUBaoGT1xyn23YOUnIY4Tzxx
rg+f25HW2O5dj6LRdVwYnv5SDCOexMPd+DpAVy/ywNQwu/W9hu9/IqmrACbrIPYY
dw7xoVvHRraQKXUY9kFN6tJ8TaVTLpK1m5ZqeLgmxbmRfqGyucQ/9IjL4tRB/yID
+UY7onP0K8k4chMipyVUcu7RtgukuWJ8AxqmQe4uTbCjmBip90+PUltTN2YPZeTW
QTPyIKJ4aflxG4qEz7LaZ6bPHHms5uGIk3SKAt+yEShYtgTdAF3dE49/C6Y/lJ+v
ehSNirXVoXtJf1ZgsMR/theqQ+l/zEz5eLb9vSZfQpIRG7mgm+qpisrpsEoaY053
HYErlVS939MpBieCHjGuL6hKYQPzWjwlAZFBzMxG+cR1PauSuTfkZ4WnPwW+KS/o
pMfQyE15L+S2xz5pGgT83Cal4wzHZM5QEZsdt3rmYm3r+Ok5l9hJY298LH5bg4Ab
fFz4YBcafs2e4WUk/Sb2GQ6lh1rTzwF229QMk7YUw/OWEZVW6IBFRRjnt7oYhegi
3j+7O3howWoyicxJ/JjEmg==
//pragma protect end_data_block
//pragma protect digest_block
bcEBoxcAPX3gu/lAQZ+wkjltK5g=
//pragma protect end_digest_block
//pragma protect end_protected

/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Cfmz9QQhz8SXs8/a3Zct5jvb1c1/X/OOVhe/5zOIKTvAY7X8H0hBs6ySlRmwLGos
cAOy0fWW4c21UZ43tOLsZ6nBkwlz/XAyxTtypy6oKCiIycZg7mz6P36xQmpukuO6
pWCdxouwbIyfUblBghlHIvyDKIo+HCKYlfH/vqzk5nIdfxgG7AgjXA==
//pragma protect end_key_block
//pragma protect digest_block
fGQ8aSJRg2mJz0kpsldqIaZRWuA=
//pragma protect end_digest_block
//pragma protect data_block
UxH1PpINeqC81pXOegQ6dHpiAi6tXqrrN2YmKRV17wGMLjvmLnhmCQ31iC7WoNkt
P4LVvFxVDIYeEhcslr6z6FmWi90j9bpGZjwQJbcdyXCfZPxmbO80Hks8UAddZpI/
XhfoyYdwmRSYSGxct15xi9aQE4He2lcbWqxOJw1WTqPHIf0h7rxZyphwcU5WSxFE
WUrB0OMhwZoimIggMAIaE/b10UCNbOLVjOisNjqw37z6qhimS3cH5QK34mdDxUtA
jma94qqCxr+Zc2QbKEeewOHLZ8LiV/JG30LbQynni5BwMegsuMALLtLJCNHh9DXC
SbaJ+cGfj0IAAdck6V4rq40ko6ZNoVvCLFVe+4zz3E35Q8u4/x5YZOG4QuLVX/od
6QoQ87dm+v/JWXdU+OFGdq0twpyQoEVVJOexxNjY8jT/ZZZr1a4S4Zof/+oCSic5
6GrIoBdcx7CGgLGvdYOeOF4lmp8YSHzao5exx1ocUWGlZgRkJrfV1vRCTJPvaF3x
vrCEpx/k1MJGI5kV3lLM5BCT4xAnsTEAiPAnVupkWCp+CsZ71AZVeMXwCnAuTaoo
DtSjxElI3XwDT7v0OpQMGVRtDZLLQ8Y5lwHxOB0FzrWjc8fx7pbUI3gXe+8c80Yp
46JxvAM4x6MAY75TombU7kswPKnHkOWXN3tR/hKhCiErTi7qpJt6N32gBvIE3xDi
j2mRbpWnPRTZvzQkuC3CFhjWfh9IM4bIJXM33nnvDM9ICeigfzIJITNRoN67zD+o
WtecbNDwuqBMXJ7jtYJ+a3x//J/DJfjU/2pmyvO+7I7iMnDuA0AhOqDeEZx1JIJf
5LoPbecR+CsQAXoCPT6TM4dmFmNKQ8kxXZ2xcOoA3EV7DEeDJ/XXs3x5+Lja26Qm
hMOdLaVFiRM9zXYiSDr04uXS2T2RGSxI7eaZwfQ7HV27V6TXUio6zy9bPAzkwoR0
y2NxJAGmM3doaBiXeuTfnLzzrCazT6xEGUoSTLnlhY2+TLFxROyZ/WQZx8PSbTLC
GCnjoYOpfOgqAYdSUnWxJU2soaU5he8WaSo07Qw8y9gxpSpZxQq5QKlUXaw/xDmN
8VBuFGn8ToVYZayvqYngmSjtsBBUu3qiDN/x3ufUBVShu8geUqndoln6z6NP1I28
XHDszUUmcju5g8ehSXVkiKi76QQWzBWAwx+Vo1xZSgnBDqwyF0WhSPRpwdxypy0/
bGRZR3vF6PAyMiTjbIdozq7kDiRnyAUQ1oA+yQuum6Fsn/0jm5owhMKCTLJgQtlE
Lox/hNposv4jtFBu33mDJ9v6duimr86KyzY1vZpOMt/fMKZO3ltlFNq7hw1+bBje
kGchCEsi1Tr/8ZDxciz4yg8+7X3HD4EmutIuohRhlDIZ4ed9AqAk2gSEa77mIOJI

//pragma protect end_data_block
//pragma protect digest_block
oG0NW+l7l2RFu8WPnoMC3xwgXT4=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Retried DVMOp TLB Invalidate Transaction#1 ---> CHI DVMOp Synchronization Transaction#2 ---> Retried DVMOp Synchronization Transaction#2
 */

class svt_chi_dvmop_tlbi_transaction_followed_by_retry_dvmop_tlbi_transaction_followed_by_dvmop_sync_transaction_followed_by_retry_dvmop_sync_transaction_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
LEX9SfmHnUf67BBFflQMYzpEMsjknyopMuPU18mkSjmqGplPjym/9G9LBGft/x1M
7gz45BXE+ZVa4iFTge6k9gBiWqjOis0A5Dy64QLKHOKF77IpxoUXEZEy1zqgxi10
yC1dDZAzEaPc0ykDZmdO0pNN0IFvXgU/SvNIocZhZz+qru19ihvMVw==
//pragma protect end_key_block
//pragma protect digest_block
y9qL3HUQ/wNZeKoG4bkZ6xDZz5w=
//pragma protect end_digest_block
//pragma protect data_block
xZgnhyKwc1EYmu0KPmZ2YnMN55WVra5qRnbmVFhA9RN6h3FqmiasTA2ACcwCs3Ct
ioN3EO4dOUEx5EbFcIJ56R4Gs8RXNEfLQDvFausQuEwB7oEgHWi6cMYrf6DUk8bK
L4ye8JzU3XxZ4HdCeawfsrZY6mW9bow5HCeyT2hwM/6zyRlP1qFmeLPfxWZFy6+A
WiYxeP5DcZ8gpGn7zeLB0b5nl59FnsqSxYYgAAGH8bOxWXFL5gxGgqlTpbRjAoBb
pt4go1YdGtVXtM6YwAbw9Y9Ccbku3IWpCk2aVsMgI00CA4l9FYoTP/38WNKidSGh
O12b46OcgsVp4nly5KzARNsnkD9ffvDdYkDZaHsl+NoZCfNxinAyOKE+L7fV5dKh
9Q2tUxLqyUroBjpVCvqyN70XRm9shA2uAukWF2c8ZKjtF+yNMcafQNjv9K/+Sa/c
Zz8K9WhbGYAscdxUuzsW/N6YlOO9Oe9/e6uWr+UZl8sCpHulpPXp7Dm1K4OvVyc8
/noZZehjW5mZpxDUwlYav++keqBz5FAkWO5TwjDCCrZyAaCKZW9AWpgMVsLmLEK+
GE/+ES76OD1+SzgqUzpoBnpi6/G9bfuk4Yr1LI+Ql7ZKkE1mXb7N2chGvxnSLziU
tnTaTbikofhKuw9MxXWU2/vJ/GcNEOF6hU0NeMDhZnHVSgVLGGCKO5Pcx490v5G4
rdR8/BsBB/juLX3kYUreRr3Sm+7gQib+D7olbmX95gHRpEgpezipTL14JwP5gKSu
sP+gKraeUlsuXDFSfEyuODjxmyyVzxXGVKDTVkFeFeqORNRmnW0+woD2iD74jQ18
fG0FWARUiH9FIzSAWgt2h9q2rHIR3iRPIFKIf8x51oHwTMbDpe2z9HjF77q8x4sa
lGrZXp/YILpr/YRXsOYzyf+yzle4FoQiPyBPEhYPmXhKqb9v2d6UZAoIDqbxmmIs
+BD/9usQjC06bimrvisO3+tTNGwl+kgM8M0WqpDOJlk4ahc0iiFYrkkIyIa1vczr
xFL8Y4drLli4P/hEDSZz8d7nJY1AKNVyE175qwYZP1EdtE5moCcyzvDfkO3oWcLc
gOH1x/n+7+y50qPoXccYJqxMTusRL5OKazqYLIkDcnFWepTlg/G315uxiVYf82CC
CtsJZ3MvopL25dEIzisHHFv3806nRWz7Nl0VDrwpaI/ZEhHM6fPX9nOr87rjsNvK
j8xx2xQ3bmdLRaMRB7A2ZDq6q26N/cwgIC/W/45BJylqqjWXEseok0ubMZYr8Z4J
K9rxOQSL/Eb1gyJrYzMKYCK0xYZlPmDavNsMgEJ11L+0qHPt86uMOBMcz+Gd0GhU
a49+OGm+tXPAdwgmEPgmhox+i35oZyEM2v4hHScXjXRhL0D/vAp7uT0DRWSSt9Q9
6ALpw5noS5btQqf3l6T20Ikiv4y7bM9CV67zXp/C3/cdeBqwv6UrjOKU+CMrkPRd
ixaTrNzrfe7cgiwWCMtl8aKGRnfUEmWNcHkxWYKqNzRpRCZgBzcmoZwvXAHUrSBn
Qe9b2HQ6LgZlaImBbFD56EsSrMvrxsNZ00Cdv0ZNXBicDQp39T+0EoKaWhMczMpJ
Dr/FEerqbbJi4gMq8+XgurBt3jIASDLoEy0QdxocDBjiGZP+v3Q3B/4h8Mo9tszX
4w6sP/WS/NrtFkwMu1aeSbDMMRHmPlU/4bNDjIr8RBbHjnvnaegzqZ7gm7y50TR8
ToFC+/3+IQpFQjoaC5xmzjSM2plARnirKlJx+TDVnW4fla1VwKzw/FdpwCRAkujr
m9a6mLVm4Zrupb/FjMXLPKqozzgqSARHvSzOyR4IXbUAleZ8Jp1jA1rF5QaSN3ZY
Ki8sMBmQAYtFJ1urjDL6nJiVFcvF5NNfKwsBQi1d3hMmPcBjEaCkyodcp8+btdh6
0Mdl9BNo9wWB7pB9TfHMOLSqGB/FifS2Ap/bBi9BwVZbnu70jlbbd2lurCFUbtc7
on9L1rYAU69KqjKvzq5U4/Q2ENKPImJdO2PPG/ijq2h56wHh/Z6WYbdDWZK22Lnb
2gnlc23NRrUD1eJYzVx6cGUEbpyNaJCFJSnGPcbOPz5nI86kN8Wp/ECnwLXqNVfH

//pragma protect end_data_block
//pragma protect digest_block
iacwKIxqyCFIyGcLQxoDz8y5BCw=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI DVMOp TLB Invalidate Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_dvmop_tlbi_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UIUwyL7I/ZsBIIBfIZktGsKOEKKcRZi8BcV1eyM+Z/UY97rDTPlv0pfvgIbE27EX
LK+QFwEECsxZmfWrdyoHNPlOtjF3m8edkbytQEvOXJkh/jSikdecvwS4Np84W1i3
M9lF6dpgoyOxa/jLZVUU4EqR8jTSNFB8N5Vv+Ixpgz7g3/DVEmZ1pg==
//pragma protect end_key_block
//pragma protect digest_block
kfXbukVqLZq7x9fM3JV5+wxZgGs=
//pragma protect end_digest_block
//pragma protect data_block
0RDtqjEMtXi+LEmoPipoksTDqKkfQlgovfLOvrea1FUXGg+LmPYdweaL0rsxNFHh
1N5peDBe51EomMq+OUnnuUihIqjlR6wfBc2Cqdval/cJYErmJTMxDPDmXJgWmJJW
0ciV2ZCl4z/oowONFQm1XKFP7tKf460PmqCDvufe9ZuHorplK1OMAAnrJwwWmrrE
i4ai0Z70SPa2rQGG7QzfwrmWlzV95BmRJDAdxyPjUxpbRc9ux7mqsznsub3LLnHf
WsnwCQG+lUPGJD21a+A/AZPW/qEiSi+iD00u/bx1Z5wxPJh29iVVhug48Hg7jb6U
X8P0y0bpy8olFGddQXh/Ha3g5XPYglZFA7q5EYPG54zJajMfIbcXTbBe5aKxyRtQ
zwGGxr3hDy5BJvwdaFNzuviG+k1bBWwbJijxvRNqAgjy3jpTZc8/ND2Pm9Pv82je
52TUigY+RwE2C0twcWbn2Av2Wb8d8EUVFMzFpM3Wqw9xQUl9mCgk5Np9paZMDHIJ
+wdUAvY3LGDO6muR+O4gVE0AVHymARRvFXGRn+A7msdu+rEVn6hsbTAfLfccjhI0
I/BqyFADKV1+HFQUPpyL4x0Yk3yxgPLp9iQSQH/Ob0KuPyit8q5qOHp8/dr5DNsa
yeGs7Mjtq42jG+oe8uYU8QhlGHamOxgjsPKr1xBX8+7c1dPK9XWJenfQY6UuQL5T
scWPEC/FVV3crplqgeQKdYsKPhhZdMyT3evOW8nImqbh27jNzwoj+OLwmIyRDdW0
eCgmJpzbjMgP9ESnx/HUUUktjZyPURtPTJ2QLgpYDTUUKaiIWEU+JN4pV1IjN9Zr
C+rXeK+IkHWNFrEpmOeI9zhFsCBJO58ZWcyw6iY1OoJDmDclX7NuJlM2UVfLVwwP
z/ET82sUuXkXu/Ddw+TMo9wp8JSvrNRFssfSenBEVSGwKvy7IzsCfLkx7L2D6IJf
Po21JOviFy0mZdTnDyNrqvusyujDY7Ek0B5MmWHZXYJq6XsEFwrazTeucOPwjLlq
OvzE0lCku/Ox6DzkOyAnWwn01nvIcyJuRXR3RBeyUH3ki4QKhRa30s7RBvHYL17q
O3K5l0hn/B6Kp787UuXESlcvkc1zcgj/V+Q/bG42AaYn03USQGieW4KIH1VFMQ+g
tXdgX3rC3TRBPrHhxwfksgJVHVgJWxugsH5BPBw0nBxxETh36wf96B5M1uAZYnJ7
lzBNleWLzHFSeqJxbwOmK0P86wCrOBcCFMMY7gWGag4nZ5Bun6TUu3PiwbQcRzwN
fAp4bgUaapOHCKfllFJDHaP+pt5lHqtN/MC87fp6PeQeaZuVKq+rmZWuj87Bo5is
XkPErnx8yOPw8S2DGC+Lnau6LmnnXQ4TPWySJPl6oohECZ2WhCY06KVtpdYrHMWs
eWy/EDjY7FH9j74RPeCa2ZSqZ6U16qtpJZeFbAT+FM2ANG+X30gK8ZLxBG6+nnJU
+P+nB5KC5qPto5oCSytTNILdwASnbMmT+xwETg6c8wcP3l0nvUaKbt1vSmxOa+sA
iArKqL+XP01DSGmBjoJE2F4/uZHmijazh2gxrtwhWQclz96crNBicvTZmOZ5HYaY
yOVZ8aMYCtO1hKha1ZlQOqtUaTXSBvMygGt2VUuzUMwZfVPg0+YYfP0kvV8Bdejp
rF7NwFGQBuIIdU1EJObzaw65SUz12cM+zX0yUbMcVWl9Qq/OGIm+rzIS2/W8MUqH
t+ZKUpJeZn7BFv8A4EP07gFvdbYUhmZ/HziukYbHaQ0gi7KSqkeeiP15RIOxk+1B
J8NZrZK5Sb6jhO4rx3ilN7yr4EqZpqEb7wo5TcE0AT5w0Vw3th6XeofytBk7/m9D
5uF1s2WN3CpvUQ/OLF3xwdyAn+dID2nbaloVHpRQoRXLdJzJGyw3NQJN5FbZCTX9
IJ16t6O3ujvejgG3DEjlCJVxElOZ72rSSZetGuCTCTajng2gTB9udQPNeVL34jcJ
vJGTOSZLJKWOivFeXrsWk9Olzc3nBfsA0tEkV01dovWgRBlr4i9YzLjzz53FG6AT
W/EFYmyhQE2dGn9tFbG1xipbWn3wK0VFx+2QELbT3uapv+ei2HH9dKwd2a61jeBF
+5S85M7pAffaUQeVwA4AT0AlrHdPZmFwhZxekPA1aN1WPYgejqJrDDAo3azn6Ig3
ZfQdCnQiFFw9Oq9QYCPc0Y7CaWrRqLyEMcAiu+HlrB0Zqx+KrLONn+AAzxt7y8+j
Nbe+jbg8d4aYJoUkMmcL6eRExVfT8cuoJLVcsaUWbT9wVikIaQcqHzTfuqApZa2S
vbpAbMTA8mlr5Crym+5cFoLMfjd83JNmPY/HMqyhVJaqFfHfnsWq6TyYlvVR2wZ1
UUwLdybs3rDlTpMfoz5O15EyPbTxwAPzvtnGrSVVrNLeo/o8+e3FvcytrUN86McP
UaaTEtMNbXyGTMHdR3xmpCwlhsvub7PZRjVlPWOGD4wULqzbSIGHbdCReJ22X6Iv
MTxSRuusd2qVi1PoHDI9kW52N8/EIaQTmzRr2hGQZmWVWd/oUKSit6n1wAbMJrv2
KUxmIDaqq2dA0qIepxyojtwCHFkQBPdjYgcK7bEoyumEKeofm+i4qNZs1QJmrRMC

//pragma protect end_data_block
//pragma protect digest_block
yawS4Bvxts0yPDkcCMqYxc8LzEA=
//pragma protect end_digest_block
//pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by DVMOp SYNC Transaction followed by DVMOp SYNC Transaction followed by DVMOp TLBI Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_dvmop_sync_followed_by_dvmop_sync_followed_by_dvmop_tlbi_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RIY3XG5sfaIp6SQMVJ0SfTqByj29EM63bwhqrBuG0dOW5wpfpxdcMXtZUH7nkcj1
jKkvPaqpr+xN4xwxyNZwKIj9e49cp+rC3YAMbD9M08sQ32vD8AcXUoM9/0hJ2+mR
yjqErUTWYNle10ZRR0RUx80EzNxqrMJZD/vLSJqHrKCtxS6D0Lh6lw==
//pragma protect end_key_block
//pragma protect digest_block
lAP8Oc1F2lDjZveC+55dqBH5JNo=
//pragma protect end_digest_block
//pragma protect data_block
l+VcwUQgzbCrK8U5Oa7o7IP6MvgmpEcdoN4xpK0rnc/sYSRcCKbfSQdc97SHgEaS
NtthxJbsRy7jF4078BBgNM3/2VZ4ycG1Dep30y51R4L5h/oEmDw9ESC26y2tpHEv
W5iWWMJW+v4uP4FhrHvfqinPv7UX3Pl0XioGcMBzz+0S/x6I+I9ZPocjqcmxsO3O
zWo5auVcQHu2ZeA5tRZZAPs+fTV0sCURrRTyZbyUiyJYo2H4UsrmfgyMMakjqAXR
o/H7RQfeBNrX0oRvJUtrj5xMDizQjx5hApMI0s03Y3BbVnl1M57gfdPx7Lb2UALl
X1408eBorIAR8wb7K4vnkCnM3KWsqSoFL1Pc9cdZT+rN8tUI0gWEvHl5sQywKxhP
gCeG9r7UvLexAZu3Ay5ddXcVZG5IZkEfBT6V/J1OgdkULhq7j8UTPXmtKA0zMyas
N15qAapV1/ggdfqGSRfpskCd0S+sGwR7tGWxGj+0JgoxJR7nk7VISyUoSOVqc/iA
Bon7UldR/hRx2s3PawCff1/fpuvN3yb8zVXONYczKEIfy8dqOYKOTSFGBLlQdQt2
qjzJMwpV91fT5vKPZTGvDSzZx/a0dCpKxyAZ8eGkIKrLHOKuDxuZHI2FcBWp8Vqo
ZwvmgmLzbuRR2OVn1Ao0CeN9j6BeB2+0jdxrsetEvlTyPHVE1lB8gUuQB0FbIKZ9
ny9YyZkJGIURrLB0BtfOq4AiGypjrhFw0ysS7KabpNoysi7QZLv/KgL+TuK2KVgC
SaFKcAIiitOd8lvQt45vWlzPMOdCWhOyrdCbx5gryHi9+Tq0kvf3ZWRuTt73+Nxg
23r35psmOFDDwxtORckT5jb4mlSq7MMt2j5cYqFdZqv+epv1+gr+7SCmFYNvjb9W
mtELqpNAPXb9Qmvy5b9PZ69EQnkuwsREW0xrSvNn7uSYx/i354UikOQVgF0Tt9Ds
GcGh8jf/zUMrS+QXV7zEMo5piyvSwykxM/9UEg+Wss/mftbBQwf+FjtPh1g+WFgt
ZOLVp5n22aUPePBY+ygopv6sbRgkyqAdYrQfEEAcDTDbW4r6X+UAD5+WZCNRAhlf
CPdE6TPhhyV0kFXwyMb/rE4i5EMCPDgrmQKUqrykmFJiLt6CaVLHYsAb0HROeMXP
o75hutu8URrjpe/Pgzh1bQK+1Z0zsa5y1+qBOvQqWRzUtPgZVr7RajHpIal/pkGN
FJ2cmP3Bb6GWyxvXU2Ct1BbdmTCbsJWfRCE+bBuLDS+76xX3oAHfsxTjpOlNp3HA
kk4SlvvBD47B4qZy/c9UiyvnmbWs4vPZSxqwAS8Gp3c+7pHdX54GJ1ENUL8g/FMM
Qvd1mkVU62zrqs7FOlLYTsB980Ta78hx+lS+F2/r3woP1Yb3oVl1TuMAsxlGG48V
fRy9xguRUSvio0PxoSsBOEHR3E/3dRYgimuyzMiQ539R/X1vlMGTQz0adBOuD3SB
6+D5G9mTVCsERi8MlBp0x8fg/f0GX5rgtEWPU1OMPpUQjdq13XyNnG7XbW1Lktf7
/KnefJp2/7wlJj7FNpoZ2D5qrTC/mPcM0N0maqL1oKd7VbyLI9faUAnpFS76PQGC
BE8rKVmR9VWjH0k30sEw70FyLtuqhCzGyrukPn0x2HWn7S/Uk+V7Hurl3KarYPvN
r0zrZfK1RZzZEtwsKKeTN2SMJDmx2/73Yo3IrgGMkGuU2O4jFoDGTMejWMXuSRhg

//pragma protect end_data_block
//pragma protect digest_block
uxh/aWWWwxZIITMArOebJPDQgCY=
//pragma protect end_digest_block
//pragma protect end_protected



// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 *
 *     CHI DVMOp TLB Invalidate Transaction#1 ---> Cancelled DVMOp TLB Invalidate Transaction#1 on Retry Request ---> CHI Non DVMOp Transaction#2 with same TxnID of #1 --->
 *     CHI DVMOp Synchronization Transaction#3 ---> Cancelled DVMOp Synchronization Transaction#3 on Retry Request ---> CHI DVMOp Synchronization Transaction#4 with same TxnID of #3
 */

class svt_chi_dvmop_tlbi_followed_by_cancel_dvmop_tlbi_followed_by_non_dvmop_of_same_txnid_followed_by_dvmop_sync_followed_by_cancel_dvmop_sync_followed_by_dvmop_sync_of_same_txnid_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
eTO3bG1xDomMhCQIJaX4dhLShHrvZPjCCltQwD7a514MMcpHHY8dowaUM7ZasPsv
Fh1WjvmbNMfXcDntriMJnduNelWoPWyPjy0u3ASMIbfAiBHo16L9f8CNKLJEDQqz
mhwdYPELnXiRgX4dEOxcV40oRobNoTBTGAaPsm0xG2Aqzn40CYgkCQ==
//pragma protect end_key_block
//pragma protect digest_block
ndDabPtKdOluhm7M72Jsv8IS2lY=
//pragma protect end_digest_block
//pragma protect data_block
I4O0mHOCa0a1ld8lGVG2q+UZFOafm4ibwj06VwhGwTVsQFtN6fxruG3dLkJKfljg
vh5ZVow9Bie4IoPTwO6iqc66Zy1y0+hucCIsEvZuwKXD2BTiX3CaTDaS+B0WVS8h
2ZmrM2EwJ6AaOJ0SUJXVCud4bz8W86rfjeoFLqxX9bTpS7Dey/2FnwFWzLFjIKwI
S+NBn/3Vdfwk/b2L52zMws1XnxISVrn8y90XArmvGQzcW31kjv8+jwJhbQ/n7PTn
T2KhbHkTnfbfAahV9EMNBOhwgPIj7PYsP413VuDAQK6IkYusEGD/u1+WhOY2/z7c
5oN2gnpiUj838ImWqkMJ5GL1kiErcoAOfs72Vo8DIGo7+aPUFkb69z6D1ALY7TcV
sb95WSGAycnfQSlx8lxPjgD66bzVK5/zXx41WZsAIV62cTMTDdjKM1pZT5bZfhmW
LslCOEo0go03kFLhsZOxSysfz1u2j2yQZF/piL9u2eMgemQXTDgzBMQgpqNbnsVt
NkKbpZ7heHa5U7Z7Oq1LosXCZUGsg/UAn0cgtQzIDxnXEO9dwnA1fzvOx2BLd5UY
o+rQNUw0Bjd7MCT/xLe9Cmu9moBds5WRSPOOuvjmlLZu1XZC6i2N72qP5F4EQ5L/
pDUvOLo2R5kBDXtaLjLf/B4pUDRV5FgDt/qY4KnfvCb7+LkICLvIx/aJGnvxX+eT
dY1yjfFtMc7PTss5sG0AnCa8UGSmymyhAAQ78rSEsT36tTlJf+Z2ndlikrONkdTh
UXpEJg8KBtkw3rmex28izvjiz2Zdc/ppguBtkz8G8cHBMbghBe63hzGrYjaGIphY
WLHNGG4gKG9P1gKzmyr9yWjTjO8Ruwtkjo/smWeFrJTL4ok3KsOPamdGwqF0I7MA
CN0qjj6QOS8PM/wt5Vuz2xYh657vtiBigVCs5wwXe6pO3bLqK3587oUOHCmeccIN
OltyvENrzG9ztDToAmPUr1LZqgMH52XXaos5CS+x6YN2sJEzM8Nfm6blVpDLcLIk
WVoLUtUy5n1LS71GV96Tbkwpmj3E+GWzgQwN6ycqTTCipPblvisBehO8D8QCq3fe
VSKsLZ/zx/Knjx3qJTDKtYoxdi6M043PdF3tp3VmVORxdDwY6U7l8xHaTTjqayfp
tMuBYjdVEikXzC/5B2bQiN/TUoKfPCrr8L7ysmvWPPzL9W0V4hsM92M3B4dVeYq5
jHpMmI5S63VWQqt70oG2MdJUHiSSc5DKaFWipYqZaU45dWMmj1MnbTkXqt05kxmF
slP/9VKlTLfc//EVj+LM0YUs4AMf9rKQYNX4Te9cKaOtDFVgzQFgycJC0TIueMq1
+zu+9p0uyzOzVICDEwkJfCuyEOYF0TVdapanT36m+EndYC17KaLd2SxA/uHigfo1
dkkksr6A+y/wopdhxObQPCOTq1cOSPmNY0KHKOXU8Ll4S0SE+kNSgG8sfuxGWBlR
GoYi0Wd43weLGQEs2B5X00a5l8jG70YyYOmqVBtanrvHhXjsUhVT3R60ws69a/ny
PYQil3+yQnGXmT4Bi5hYFWm4kzj9kMIGpP53pkHGs8pttctakaiyC4auMvw5oz4r
YCgUHpuO/BTRZv2FPwU2FPthF3V+8sKF0pLkPIrztwq1EyGJqsc4qI0NaxCPBX2F
RL4tHTSitlOB6coyI0+9atqvIDsrhw/lZP79DR2Dw3wWWsXQ7PYowVEK9OWupx8I
8rnXFeGJq11CWbqsLXu8k4zwFum8aeRVf6QfUIpFWusJvgecEBvsh/Dxud1zPawb
q5RkEHNsqSIVB3FJyC7CMTHUXXGqdtnr32xL1FITk6SYqY81qh6ebKTquG0UHAej
0vt6TPgoSdQXwQG93Ra8Ch0d1TmXOtnIGbN9SQOeHMZTjYPxguRcSxndfTuVoO1M
hJLwEcbz0+I1nSqFTA09O0o4YeKi6XTCylm6DHUE+9axfAumt9rzaUQ5pWmy2iFI
QfFbfEQAtMMlWgFNwVLNKiTKs2O4fdgKYKSwE5/y2XxKoYG47QQed9wZSOxKsN32
pijzjWCB/jh4t/R3Ez6WTi0SX+qE3xkyzu+GPQTpafb6UKvoWJrqOWpyBZIOcnSy
ah7PbYuOfI5XhlX5f3DrYkD09lnirMlNltEDbQgdiNHxL0X8SIUFS0h49GfdbQnj
fSr71A8F65o+FKHeCxbBWI7gALSv0+XhWB9hlcFJKMtD3nmW/Oz21z2vR7Hh8OsL
41bYdXZH77eBVQ6vlQrTilANRL7FFCcYG9KZ2qTixU+++pLQV6FUzEvVdEPUX8Tp
ov2TMDDHRtb1iNztKY3XpC8NJPLCDm9q5fsTegdyrPCN3/jUd3qIhsSAp+/9mJwM
Wc62mXm34VwFG/EM8B2pJdhkQnMOn32SYdVUW/8nXDVZjz3cDChCrnMcGo468TRG
7rEyHB0Pm8kGRIQ17mJsgn3r7n0j6l7C1yGYBMMbd1lg9tu2ooeCJUBJNdi6xy2f
ktoLO5RCmlItOKvgmN7colkoiOG3TgI2ri/KXG7PLew=
//pragma protect end_data_block
//pragma protect digest_block
To5VVOejEjymDEVDVH/me59ay+c=
//pragma protect end_digest_block
//pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
1yLzGLmMxRnLvi1vO9EOwGqRSovVdKHf6Y6kx23VmmJqi/qIdw0iYHYl5RL4ltc7
+0h3TMnn/9jRN0M2OTkjzzRTT9KMGN6XB3tL8hZi7Loe0kzQ+AdyGisS/2aJyR5e
kb3xB58EKJC0KmMm5kSst9991TFfGEM5OSw73fZ45CbyD8AIBh8oSA==
//pragma protect end_key_block
//pragma protect digest_block
knUcc/QXEqG+oLAz6QPWTN04Yfs=
//pragma protect end_digest_block
//pragma protect data_block
OWGj99rvI2AAPinuqhl5MfNflaaydFxvn1N3lkfYTL2tVpEC0LqG34pdd6VXByah
00O4H+wAhm9J3qDfDSi3yTKoo8cWQA9ZFP1fHtmDv+NBM0yt9RS4mABLE31fsHZX
gXuYyyTS6+hQ+I935498wCiM70IOwuzqdwtFvJNV/932aY/nGIFBkGdIQQOJsbo2
1teq6VTe+ew4fjgoWYi3Kp1iO6ESnELC/8Dq6aGRjgkV2Sm4nrWKiK8RHBBICik8
yg4arHlMMZIfmUv8s8+W5iCfxP2juWx2NNLC8m4JDjtj2kfEcPdrYMdG2bR3Q7Vc
lv0W2POwLTEKAVO5SopMWfrhY/akyyln4aH1Z7NevIihrjOvBSHOWiOC7uUGJ0ts
1z1itIyivxi0PbcJPadHwtedTmAd/Z5c/rHqrAraIFx5FzBythMybtznSrsmgYua
lSK0+G3M+XHPKmYAXcEYlISnQ9trCOxoIyBqz3jAMR/G4Zf/Z9whN5i4ShAaJre/
XmEfE9ckaa3t4jEyTrboigNrD9KXcZ/6O/MhCydAxnHKdKxd5iNrBoNQhJTZZtxW
V7mJT3KyOj1nihETCmjMe/KfuX6LPtg2KYdYddjRBKrAoWQnZ9WihOpArpLvLLnM
cugCGOfds5ObpLJaG8inD9XdIKNmjnku1beP+8AQ99RMH/mHmCBv4rhl4Uatnu0z
TD86ggrGE1f+1hLXL6zLcZIpm/8VGoH5g6+UkgBv9ImCYil/XdgYwyoDN67WNkiX
hwUFoSUiesPp9c5bDakG0wkrQPGD5DSIYWmgH8bvMuKtsez6uHHRShlI0zwVhqZn
Nf8uTZSwSulwnwmlEjHl3xOFnOWJVvHFJwYaAMVYGji+e1jNy+3olDZJkCJ3sWf7
RrDSAvGefJP3eWkQ4nlH7GfgngOyu0x45C2xvYKcm8axNpj1DOTHRJ8d/DzaHfm0
1SFYw6x0iLmNQ/iEB6bavAGx7Zj46J4AADcbD7M74zd3rGftNo9G2Li08CZv+7OH
wmzVcIX7YXzeKljn8S2j59dZM2FVUg+CXuz/0lecS/1mdscUTl76WhN/iCA0jxWy
w/L02d5ELjJI8CU51f0sg3KGejoarmRJ9Y6a1Cso0EYR5V05Cb43f8AtRQqrdUya
g5Y3oNabnnkc1KPtoEo/LF9MfsGvlJ49+sEUAIs1kFtVHFYh4kLRcjTkIWRW/tN9
ShdQXBKIuYQUv4nj/feKoFny7goK51nhwNmwtKBTvDZkNwCdYGRHfPErQNsKaX6E

//pragma protect end_data_block
//pragma protect digest_block
LP4Xn+j2lC5lI4dWe4nQk4rjYdQ=
//pragma protect end_digest_block
//pragma protect end_protected


/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * DVMOp TLBI followed by CMO followed by DVMOp TLBI followed by DVMOp SYNC Transaction
 */

class svt_chi_dvmop_tlbi_followed_by_cmo_followed_by_dvmop_tlbi_followed_by_dvmop_sync_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SnAB4ddjlEGPmLMukkRAnF9AdtDo+825/YLNpy7/3xeKy7kUPSdTQ1U1cM+qO3xT
MenNr4rFRKV0xOLVipwrHy82Ckrj3BsOOwFUzkQltMgFttyUxzNPElPEWikE4QCx
b/QrTLZPtXs6+30nZaoJKaBnVhrNSGjLU8+Bt8h8F7wAWIcRHz1XUQ==
//pragma protect end_key_block
//pragma protect digest_block
H4e+fQzKTilSU7BVLLybLa3gH7M=
//pragma protect end_digest_block
//pragma protect data_block
HfR4IQWLjvJUEfFuE4FqW1iokULDCFUjbsZHE/ebnQVVpp6lTn9GVFXnPGnDkkd3
+D/SoieVFvYTvs1YD1FNVpUTEjOaWg5vHGxFJeIaGRchlQTRN95YmM2J9+yKEk6U
kRnzs8i1Tzn4LVCKdSItxZ64FM+BH8sLPzaX33e5sNq092PdvfUm9i5c5fR1myLy
i+ae0HJzeuMT2FpS7NbL5HTaZ75tKpyctbh+JcGekJmxq0j/xgUg2KXYnHrRYtAx
/oKAS8HxyE8m6f+iIpCcIjsBm8W+iITL4eLNk8BvYsIEMBTs64dUPgZeqNDN9+lC
uEpfblcT31Ut/Wyj+wyqybs85LRud0dK8e3JM7Ursbw5SkuT5yS0dQ9sNSjWk7mk
XMMAzcrFCPVm2yP+Mn/ptX5W+WVZUNStUjcPE7gc4sGcuAYUivLidsDTNQ4l/ahc
aGPc2TgE8TGoYgNL8Yp7cQ8EtIMgZ2GS+CHemYiTf1iU8eMaz2rjfvCWzXao1W0n
UdC0RsUQgUa4pfs7EO8GRuyWJnYeHCoJFqULLXKsABNJnccgkXIO6zDARmuahUhX
W8i9bpbizgvK5faXkiZiaAe8XjPql53mCIPbHhURahWKdrnf59LqsVmhmrPcFQ4a
7Y/LayTXSQ6JK1jWlVzCpQ5C+U5/+XB3WIDixXjnsW1HOgmlb/rkBjphpfcwEozx
9U7R04Bqn1/26+BAnROUShteB/j1A1UHzrSZekGPW5B50eLh675CZ2BY7HvxhKLC
wyB2EwMbRr+qs3yFyLITCf7f5ceeG7lLrr21hfzKcSZg5Ea5Vgfp9gK7Z9yfY5Ju
6tgbvEpURE1I2nFZQtvLcRiCtcdBDNltD8NJ6YqkFxnVkc85v/GtGWxUBDuocsex
9jSll3IbOBmpmiKI7b7QL4q07FjEsVYtEw5+MkoOXcvJZgVX6pTzoiBJPWmtXbR6
mYDyBOt4xcvJ0MXoqfhRWuUrkiRN0cpyqmIseK/n6A64Kz09LdbMrIDImUD5dxGu
58RZnGqwDeWviZMkEFz4sABlvZbdh7NdgX2Ly4/CaAurRYqTMJeGrZM47rrnNPuI
Tr//I+AIU5xP6ij2QPFkHjeslj3v8MAfxMih2oM7qp2YsrIhZDkA3WOWK5IqVSky
ycq0siPvMWpyyZ/b/cuvJfg2yuAcGtrPNUorxq5j1Bta0oyQNdtlSRggSffUFTCg
c3lknkO8Not6IPUYJJrr59C33taqNCHS4WANHmivHJiQyvL1FXZgoX90XUJZjFit
3xUQc71l0YAVokrYl14kNwZxBL9nFL82hSveltfIDLDjzCKNy6ybt/fVTjBNItLb
FUpc53JY8z/BBfVOJgAkiZ4zFQlkwYIPWZvOIA3WO69nk8wCXyzSmUsUfIDA1/Pv
MGd1fxBdWNf/RSRAehl9+AP3PlagEHUbmufeoltVaCah+tac7qaSVGVZqDInFpwE
ZrikciBbg4CuZUGDtg15FbSEcfdDtxPgc7hAeCovefDBBTCwsk3MUhFm39QqdQgG
FYYaXo/GHHYTZ0fRFZXnkJpWVYqKYO+skBl8qOipUrWMUrB7QB/4IxbP5gbsUhOd

//pragma protect end_data_block
//pragma protect digest_block
FIvW7xxL0NqoVUh9aDz0GCENBEk=
//pragma protect end_digest_block
//pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store
 */
class svt_chi_load_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2coj35PH8gWRlZg/cdAnNsRE/Emk11lz43lc1SToNrCPJfbby7u9HnRLLt+z2yFt
6hF+v8uWgawa3KiglZg4qLCRl85Qv9MO87DxO7ZJ4rRPkCgtgyBeyqU8J7KToqU/
AnkZTqPQ721kbuwlz4IZ00ylt9alihOn5li/RyuiK81JG9tUIGxkFA==
//pragma protect end_key_block
//pragma protect digest_block
KNQlpaMLzmYBIV13H+ROMzp8y9M=
//pragma protect end_digest_block
//pragma protect data_block
uG42+h8gmPzwu+GqsMqDVdfQVt4iXrPC5bxE1taWneFx34ehENYqX37KVrRkFjUG
6XOl+jdfjmx0T3LYD6CjdaDEkz63WzHnS8A+wDkzHDvqYx9DVOn2NMTintbRG+Ol
2MKOmQfBenQcY3fttQKEbrk/88M9nQ22yS2mn0MFWYOX+LjmwHowmUzWQaNxiQ/2
kPov5SGUaZFE0CsiAeYrWzVKutGqB4gf5etzNOkMGeYhzn0QVgCMjx1p39mgT5Q8
gMBvPShSOHNChq48MK/cwCOGBFBc7OpzBdddUCnq1IqCvkx6gxAFkmrieZG/cCdx
48LCFWCNjog0cMpsF9lUEwgNdirSvnXwf22H2Nje1VjZSwnDmiiRykewOyENa28W
gTxyXIeb588MrqKsyIMzoB8njuWE3tJ1P3yEmRPRiEZAtEfGcV9tQ9EJxbDS2R6M
uMl8TW4CTOVty0WmrwXS2HDS8kZkG+jrcmua7rOcE0x1lN9H39uE3kVj6eIN/bC0
+ZF4T+Um+pBOuNDM/1Uf1S+JuG7achXknyRbLQQwRTEPz2PUVoNBOsbvMtzSJSpH
tDM+YpBiKepAZnuuPmZnkH7LhMVtDdbo7EEbWNLJ5odJC4Y3COZSozG+/g2/i+IE
2G4S/HTgtLDOa17Q8lOuLRwS9Xv5FA618Uksddj9ooKy1Vp03NtWNihvfb4fh5ct
IyQwkY6QjoBIRzz698cBjAwxtYT+Vv+/FN842M0GRUP0FinZ7dEv1bUYeYTVh/iC
6RidVvqD9w8xkDH0wWMTLmsLOYTn4Z3a9neDL835B8GlrS4RmM7Qjtdfz3P9K/H6
eO9H229afyRor64uG4MqMIM2V0KZ63rQ+EIoT5F4z7U=
//pragma protect end_data_block
//pragma protect digest_block
rwHAdHsBPL4UNvlmgTOV68f3xQ8=
//pragma protect end_digest_block
//pragma protect end_protected


// =============================================================================
/**
 * This Class represents the following pattern sequence, which needs to be scanned within the
 * CHI Transactions.<br>
 * Load followed by Store followed by Store
 */
class svt_chi_load_followed_by_store_followed_by_store_pattern_sequence extends svt_pattern_sequence;
  extern function new();
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ubTzQyt7eUv4TgalCXX8mIi+hyke5mGVn0d3P7S1c4i+L3Z06hv23hvnk5ZNXb6o
sg4I+F9qpKtlrvQ1eH9GSPZJ/NvqE7gvi3P/TQ0c5DoV8Zzm3kuyi3U+11ccGdVS
7uWhmEgLvjV/jel1iWExFuguUH0e1djBxzjWiIkGHpDSWB7GCqa9lQ==
//pragma protect end_key_block
//pragma protect digest_block
DR4cYEW9f1nzRzY8zVQHYmBWYm8=
//pragma protect end_digest_block
//pragma protect data_block
w4O/hsy5OC5b0t7R/esDQEB2KvCNbf/hVE7+GhjbS4W0LlLiUV+1CYDTC5/Sl0oL
NJJvx71QYoBpbdFihJtd+ADHOj50/grYjWvJLEXTdqsYgjfgEm1BtgaqSBGtWW4c
L3sQS9d/xQSfhjXI5YOvkHykoVUssc2blJkpD6XRNuVVU8/4cJi2ANogrX8RWfAx
9IqAXxnSnGWm0driuQ248sdMD4XEw6MmM0oj3n0abg8i/dw9229xTv46yLj3uECT
p5PymPjU7g9Xs1f7+pZb4gDzRQgMaYS/BerZ60Fx+BmO/hp0CkSPaHNp4UqbDxEA
PESYPmAP51cwLX+ruDpJd/tgcnPl/hh/MOKlgXHS15lyDbCZo4fKfXfJUEabU0yU
D5hOcdJP0QBrtnrVhmaSY5oRMxyfgndGxS3wpqladYicJUb9PVz2usYigf+QYkFA
lc5YFTVKisf0AvMnuw/GRu5I1AOh/PAz/3gcKctT4Z/9POC+MpJ4xXvhqfaru+T2
mVfh3pw/Dv82oR3T7zuubKmQwGiFzs23Sm8LGZLxtX4uTRokWIZ1ZonMmhrJd9em
/Tv/CLgcwN+02B3p07CE41I+H52hw9olk/VdwhlecLzmiffqhsAZXNDFJoqiQeJ9
aWvF47nfIZX2qBoZdRSWCUKbsL4nk8RVsSYIjZUQpZlIFEk65itERD+nZFF86Mdx
kDo44ZzzaRzwPtyKQjRfkfcWT7GltX74Z6ed/Gf4VPbSCuqVouQaCg3kQuTDcJJk
3/YI4KnfFIZy8a3q+C7WTRlNcvU1DxMo2WH+JrYnTI362v/KXaNo9/wFHxnXN35u
IKse/O9fm+QH7hWszEtnVAuqyYHwBbe04ERDAA7d6GsNSPNnvO94iLGqiN5xjxZp
GybNX0b1VyfA3YtXmW1OiZwVj2uSMuE7nnwIigcsPO9VC0+iBmPEB8/2itx2seq1
Af1672/Vks6pZstDd8L1FlK8n6esYF+a5hpSGH62gMFfDh3UrHWiYUMNZSatAK+y
VzMNXmqVQWMmzNsnq9kGyETdBtoCIZjDy1+86KM7cTEbMX4ULK638vfRsO10DzUU

//pragma protect end_data_block
//pragma protect digest_block
U/nKAPmVdQ0sp41QnPlyHh6q530=
//pragma protect end_digest_block
//pragma protect end_protected













`endif  //GUARD_SVT_CHI_SCENARIO_PATTERN_SEQUENCE_COLLECTION_SV


