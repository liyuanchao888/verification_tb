

`ifndef GUARD_SVT_AXI_PORT_CONFIGURATION_SV
`define GUARD_SVT_AXI_PORT_CONFIGURATION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_system_configuration;
typedef class svt_axi_system_domain_item;
typedef class svt_axi_slave_addr_range;
`protected
T1^R7a^O76_HgK=D75L)M/O7H12E,.,4U<4cg#U[7NL+_60V2<OV-)SADe_e4geL
OTWXLGe&<MSH?Mc[=I&M??2CL,+K+776S\/-aBe9a#IQT-353^KNeN:F?<RJ0dBM
(OWfU4[a)W<<VcU4<LMRK./HdF5eUT9K6ReF#?\;/:,6d2Fe;\WS;>Lf:8dJFXR2
<>H[2N(Vc_d==<A_D(#2WTW:\-JMP#+<4=V1#FV2/=+7e.>,F6;OGf<KA<&_[TAA
^QJ<:W9)T?V4He/K91b9DWPW:8UCR0f3bH)1]TC99DY2SAJ0,>6[Z:W7(-=T>=P>
+>Pa4:e:U]40RVUNM4?^0J9a=:d2NQaF?>Jb0-&gBgMc9VPR^)&ZT-d.<8Nc;7I;
aVg9MEOJJW//fFR</Q70g5=KJ2KUD5>L4UMCBHOK0_#R78U-0^g.&B,Cg01_5D-W
;V=H<3:\TG47]+80@d^@,/b0?.U,AWNGX,G9RX3HNQ+IbS/4=;MC.4>DEb4afA&2
C&X.]OO=>4W6=dW4/?@UMEZ9ESQ_A[1H8f>;7QDCK=C@)KY5FN/,]\4MQE<D^a0V
KM+5-.GUON<bD?[_E(Ta@@++,#-c2]O>cHfe[WO3UU)a_X;fCMf]KC>94C;48?#J
[a6Kf]VR0bJU1&1)B_?5Pe);OT]HAd2<U(]f@(DU?.4bfLQ>V<&-I#-f9+aE]+[T
fW[9Xd5<DfNJVZeMZU;T7/)<Ng)6ES_W:PV08ALaIgg1)4]@JfDI3<T48XA9?G4;
4=?>X8I5gc]ROQ;7B[(PL,)5O^FZZ?5gTSTZLAW4(>2-3TA_fE+d&Q<ad24_:W#E
a@-J3(4_:Y_\<@bQE__.?0ZIN<-?GUM7=\,gU[XCXK&W,.76c(O7d(_^]W;4Yf5.
9@L#J;R:FT\\.$
`endprotected


/**
    Port configuration class contains configuration information which is
    applicable to individual AXI master or slave components in the system component.
    Some of the important information provided by port configuration class is:
    - Active/Passive mode of the master/slave component 
    - Enable/disable protocol checks 
    - Enable/disable port level coverage 
    - Interface type (AXI3/AXI4/AXI4 Lite/AXI_ACE) 
    - Port configuration contains the virtual interface for the port
    .

  */
class svt_axi_port_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
`ifndef __SVDOC__
`ifdef SVT_AXI_SVC_SINGLE_INTERFACE
  typedef virtual svt_axi_port_if AXI_MASTER_IF;
  typedef virtual svt_axi_port_if AXI_SLAVE_IF;
`else
  typedef virtual svt_axi_master_if AXI_MASTER_IF;
  typedef virtual svt_axi_slave_if AXI_SLAVE_IF;
`endif // __SVDOC__
  typedef virtual svt_axi_stream_if AXI_PORT_STREAM_IF;
`endif
  
  /**
    @grouphdr axi_generic_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr axi3_4_config AXI3 and AXI4 configuration parameters
    This group contains attributes which are specific to AXI3 and AXI4 protocol
    */

  /**
    @grouphdr axi3_4_timeout_config Timeout values for AXI3 and AXI4
    This group contains attributes which are used to configure timeout values for AXI3 and AXI4 signals and transactions
    */

  /**
    @grouphdr ace_config ACE configuration parameters
    This group contains attributes which are specific to ACE protocol
    */
  
   /**
    @grouphdr ace5_config ACE5 configuration parameters
    This group contains attributes which are specific to ACE5 protocol 
    ARM-EPM-033524 Version 2.0
    */

  /**
    @grouphdr axi_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  /**
    @grouphdr axi_signal_idle_value Signal idle value configuration parameters
    This group contains attributes which are used to configure idle values of signals (except "Ready" signals) when "Valid" is low.
    */

  /**
    @grouphdr default_ready Default "Ready" signal value configuration parameters
    This group contains attributes which are specific to ACE protocol
    */

  /**
    @grouphdr axi3_signal_width AXI3 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI3 signals
    */

  /**
    @grouphdr axi4_signal_width AXI4 signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 signals
    */

  /**
    @grouphdr ace_signal_width ACE signal width configuration parameters
    This group contains attributes which are used to configure signal width of ACE signals
    */

  /**
    @grouphdr axi4_stream_signal_width AXI4 Stream signal width configuration parameters
    This group contains attributes which are used to configure signal width of AXI4 Stream signals
    */

  /**
    @grouphdr master_slave_xact_association Configuration parameters required for master and slave transactions association
    This group contains attributes which are used to associate master transactions to slave transactions 
    */

  `ifdef SVT_VMM_TECHNOLOGY
  /**
    @grouphdr axi3_4_generator AXI3 and AXI4 generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for AXI3 and AXI4
    */

  /**
    @grouphdr ace_generator ACE generator configuration parameters
    This group contains attributes which are used to configure stimulus and response generators for ACE
    */
  `endif

  /**
    @grouphdr protocol_analyzer Protocol Analyzer configuration parameters
    This group contains attributes which are used to enable and disable XML file generation for Protocol Analyzer
    */

  /**
    @grouphdr axi_performance_analysis Performance Analysis configuration parameters
    This group contains attributes which are used to monitor performance of a
    system based on measurement of latencies, throughput etc. The user sets the
    performance constraints through performance analysis configuration
    parameters and the VIP reports any violations on these constraints. The time
    unit for all these parameters is the simulation time unit. Performance
    metrics that involve aggregation of values over a time period are measured
    over time intervals specified using configuration parameter
    perf_recording_interval. Measurement of other performance parameters that do
    not require aggregation of values over a time period are not affected by
    this configuration parameter. VIP reports statistics for each performance
    metric for each time interval. Each performance parameter can be enabled or
    disabled at any time.  Monitoring of a performance parameter is disabled by
    passing a value of -1 to the parameter. Passing any other value enables the
    performance parameter for measurement. If a value other than -1 is supplied,
    it will take effect at the next time interval. If the performance
    configuration parameter values are changed during simulation, the new
    configuration will need to be passed to the VIP using the #reconfigure()
    method of the top level VIP component, for eg. #reconfigure() method of AXI
    System Env will need to be called if AXI system Env is used as top level
    component.
    */

  /**
    @grouphdr axi_qvn_config AXI QVN Configuration parameters
    This group contains attributes which are used to configure QVN features in a
    system.
    */

  /**
    @grouphdr axi_tlm_generic_payload TLM Generic Payload parameters
    This group contains attributes which are used to support TLM Generic Payload feature.
    */

  /**
    @grouphdr axi_traffic_profile Traffic profile related parameters
    This group contains attributes which are used to support traffic profiles.
    */

  /**
    * Enumerated type to specify idle state of signals. 
    */
  typedef enum {
    INACTIVE_CHAN_LOW_VAL  = `SVT_AXI_INACTIVE_CHAN_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_CHAN_HIGH_VAL = `SVT_AXI_INACTIVE_CHAN_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_CHAN_PREV_VAL = `SVT_AXI_INACTIVE_CHAN_PREV_VAL,   /**< Signal is
    driven to the previous value, ie, the value that it was driven to when the
    corresponding VALID signal was asserted. */
    INACTIVE_CHAN_X_VAL    = `SVT_AXI_INACTIVE_CHAN_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_CHAN_Z_VAL    = `SVT_AXI_INACTIVE_CHAN_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_CHAN_RAND_VAL = `SVT_AXI_INACTIVE_CHAN_RAND_VAL    /**< Signal is
    driven to a random value. */
  } idle_val_enum;

  /**
    * Enumerated type to specify inactive wdata bytes of signals. 
    */
  typedef enum {
    INACTIVE_WDATA_BYTE_LOW_VAL  = `SVT_AXI_INACTIVE_WDATA_BYTE_LOW_VAL,    /**< Signal is
    driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_WDATA_BYTE_HIGH_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_HIGH_VAL,   /**< Signal is
    driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_WDATA_BYTE_X_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_X_VAL,      /**< Signal is
    driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_WDATA_BYTE_Z_VAL    = `SVT_AXI_INACTIVE_WDATA_BYTE_Z_VAL,      /**< Signal is
    driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_WDATA_BYTE_RAND_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_RAND_VAL,   /**< Signal is
    driven to a random value. */
    INACTIVE_WDATA_BYTE_UNCHANGED_VAL = `SVT_AXI_INACTIVE_WDATA_BYTE_UNCHANGED_VAL  /**<Signal is
    driven to initial value. */
  } wdata_val_enum;


  /** Enumerated types that identify the type of the AXI interface. */
  typedef enum {
    AXI3        = `SVT_AXI_INTERFACE_AXI3,
    AXI4        = `SVT_AXI_INTERFACE_AXI4,
    AXI4_LITE   = `SVT_AXI_INTERFACE_AXI4_LITE,
    AXI4_STREAM = `SVT_AXI_INTERFACE_AXI4_STREAM,
    AXI_ACE     = `SVT_AXI_INTERFACE_ACE,
    ACE_LITE    = `SVT_AXI_INTERFACE_ACE_LITE
  } axi_interface_type_enum;

  /** Enumerated types that identify the AXI interface category. */
  typedef enum {
     AXI_READ_WRITE = `SVT_AXI_READ_WRITE,
     AXI_READ_ONLY  = `SVT_AXI_READ_ONLY,
     AXI_WRITE_ONLY = `SVT_AXI_WRITE_ONLY
  } axi_interface_category_enum;

`ifdef SVT_ACE5_ENABLE

typedef enum {
  STANDARD = 0,
  BASIC = 1,
  NOT_SUPPORTED = 2 
 } mte_support_type_enum;

typedef enum {
  MPAM_9_1 = 0,
  MPAM_FALSE = 1
 } mpam_support_type_enum;

`endif
  /**
    * Enumerated typed for the port kind
    */
  typedef enum {
    AXI_MASTER = `SVT_AXI_MASTER,
    AXI_SLAVE  = `SVT_AXI_SLAVE,
    GP_MASTER = `SVT_AMBA_GP_MASTER,
    GP_SLAVE = `SVT_AMBA_GP_SLAVE
  } axi_port_kind_enum;

  /** @cond PRIVATE */
  /**
    * Enumerated type for the kind of inactivity period for throughput calculation
    */
  typedef enum {
    EXCLUDE_ALL = 0,
    EXCLUDE_BEGIN_END = 1
  } perf_inactivity_algorithm_type_enum;
  /** @endcond */

  /**
    * Enumerated type for enabling a particular version of ACE spec  
    */
  typedef enum {
     ACE_VERSION_1_0 = 0,
     ACE_VERSION_2_0 = 1
   } ace_version_enum;

  typedef enum {
    ALL_INTERFACE_TYPES = 0, /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE or ACE_LITE interface types. */
    AXI_ACE_ONLY = 1,        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to AXI_ACE interface type. */ 
    ACE_LITE_ONLY = 2        /**< svt_axi_transaction::force_xact_to_cache_line_size 
    will be applicable only for the agents that have the svt_axi_port_configuration::axi_interface_type set to ACE_LITE interface type. */ 
  } force_xact_to_cache_line_size_interface_type_enum; 

  /** @cond PRIVATE */
  /**
    * Enumerated typed for the memory kind
    */
  typedef enum {
    SV_BASED_SVT_MEM = `SVT_SV_BASED_SVT_MEM,
    C_BASED_SVT_MEM = `SVT_C_BASED_SVT_MEM
  } mem_type_enum;
  /** @endcond */

  typedef enum {
    RECOMMENDED_CACHE_LINE_STATE_CHANGE = `SVT_AXI_RECOMMENDED_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE,
    LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE = `SVT_AXI_LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE
  } axi_cache_line_state_change_type_enum;

  /**
   * Enumerated type that indicates the reordering algorithm 
   * used for ordering the transactions or responses.
   */
  typedef enum {
    ROUND_ROBIN     = `SVT_AXI_REORDERING_ROUND_ROBIN, /**< Transactions will be 
    processed in the order they are received. */
    RANDOM      = `SVT_AXI_REORDERING_RANDOM, /**< Transactions will be 
    processed in any random order, irrespective of the order they are received. */
    PRIORITIZED = `SVT_AXI_REORDERING_PRIORITIZED /**< Transactions will be
    processed in a prioritized order. The priority of a transaction is known from
    the svt_axi_transaction::reordering_priority attribute of that transaction. */
  } reordering_algorithm_enum;

  /**
   * Enumerated type that indicates how the reordering depth 
   * of transactions moves.
   * 
   * Example:
   * Consider the read data reordering depth of 2; R1, R2, R3 and R4 are the read
   * transactions to be responded. The behavior for different types reordering depth
   * is as follows:
   * - STATIC:
   *   Once both R1 and R2 are complete, then only the reordering depth moves:
   *   {R1, R2} -- to --> {R3, R4}
   * - MOVING:
   *   If any of the R1 or R2 is complete, then the reordering depth moves. Suppose
   *   that R2 is complete before R1. Then the reordering depth window moves as:
   *   {R1, R2} -- to --> {R1, R3}
   * .
   */
  typedef enum {
    STATIC         = `SVT_REORDERING_WINDOW_STATIC, /**< The reordering depth moves
    when all transactions within the current reordering depth are complete. */
    MOVING         = `SVT_REORDERING_WINDOW_MOVING /**< A new transaction is considered
    for access to send read data as part of the given reordering depth when any transaction
    within the current reordering depth is complete. */
  } reordering_window_enum;
  
 /**
  * Name of the master as used in path coverage
  * This field can also be used to specify master specific
  * slave address mapping. Refer to the documentation of
  * svt_amba_addr_mapper for more details
  */
  string source_requester_name; 

  /**
   * This queue will hold the names of all the slaves, including non-AXI slaves, 
   * to which an AXI master can communicate.
   */
   svt_amba_addr_mapper::path_cov_dest_names_enum path_cov_slave_names[$];

  /**
   * Enumerated types that tells ERROR response handling policy for AXI Master and Slave.
   */
  typedef enum {
    NO_ERROR = 0,/**< When set to NO_ERROR,vip should not report an error on receiving decerr or slverr response. */
    ERROR_ON_SLVERR = 1,/**< When set to ERROR_ON_SLVERR,vip should report an error only on receiving slverr response. */
    ERROR_ON_DECERR = 2,/**< When set to ERROR_ON_DECERR,vip should report an error only on receiving decerr response. */
    ERROR_ON_BOTH = 3 /**< When set to ERROR_ON_BOTH,vip should report an error on receiving decerr or slverr response. */
  } error_response_policy_enum;

  /**
   * Enumerated type that defines the behaviour of the VIP during reset
   */
  typedef enum { 
    EXCLUDE_UNSTARTED_XACT = `SVT_AXI_EXCLUDE_UNSTARTED_XACT, /**< Only those transactions which have gone out on the interface are ABORTED. */
    RESET_ALL_XACT = `SVT_AXI_RESET_ALL_XACT /**< All transactions which have already started along with the ones which have not yet started but are present in the internal queue are ABORTED. */
  } reset_type_enum;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enumerated type that defines the generator source for slave responses
   */
  typedef enum { 
    NO_SOURCE    = `SVT_AXI_NO_SOURCE,           /**< No internal source. This generator_type is used by master component. This specifies that no internal source should be used, and user is expected to drive the master driver input channel. */
    ATOMIC_GEN   = `SVT_AXI_ATOMIC_GEN_SOURCE,   /**< Create an atomic generator. This generator_type is used by master component. This specifies the master component to use atomic generator. */
    SCENARIO_GEN = `SVT_AXI_SCENARIO_GEN_SOURCE,  /**< Create a scenario generator. This generator_type is used by master component. This specifies the master component to use scenario generator. */
    SIMPLE_RESPONSE_GEN = `SVT_AXI_SIMPLE_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_simple_callback is automatically registered with the slave response generator. This callback generates random response. */
    MEMORY_RESPONSE_GEN = `SVT_AXI_MEMORY_RESPONSE_GEN_SOURCE, /**< This generator_type is used by slave component. When this generator_type is specified, a callback of type svt_axi_slave_response_gen_memory_callback is automatically registered with the slave response generator. This callback generates random response. In addition, this callback also reads data from slave built-in memory for read transactions, and writes data into slave built-in memory for write transactions. */
    USER_RESPONSE_GEN = `SVT_AXI_USER_RESPONSE_GEN_SOURCE /**< This generator_type is used by slave component. When this generator_type is specified, slave response callback is not automatically registered with the slave component. The user is expected to extend from svt_axi_slave_response_gen_callback, implement the generate_response callback method, and register the callback with the slave response generator. */
  } generator_type_enum;

  /**
   * Enumerated type that defines the generator source for snoop responses
   */
  typedef enum { 
    CACHE_SNOOP_RESPONSE_GEN = `SVT_AXI_CACHE_SNOOP_RESPONSE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, a callback of type #svt_axi_master_snoop_response_gen_cache_callback is automatically registered with the master component. This callback generates random snoop response based on the cache line status. */
    USER_SNOOP_RESPONSE_GEN = `SVT_AXI_USER_SNOOP_RESPONSE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, snoop response callback is not automatically registered with the master component. The user is expected to extend from #svt_axi_master_snoop_response_gen_callback, implement the generate_snoop_response callback method, and register the callback with the snoop response generator. */
  } snoop_response_generator_type_enum;

  /**
   * Enumerated type that defines the barrier transaction association approach
   */
  typedef enum { 
    RANDOM_ASSOCIATION = `SVT_AXI_RANDOM_BARRIER_XACT_ASSOCIATION, /**< This approach type is used by master component, when the #axi_interface_type is AXI_ACE. When this approach is specified, a callback of type #associate_xact_with_barrier_pair_xact() is automatically registered with the master component. This callback associates barrier transaction with normal coherent transaction in a random manner. */
    USER_DEFINED_ASSOCIATION = `SVT_AXI_USER_DEFINED_BARRIER_XACT_ASSOCIATION /**< This approach type is used by master component. When this approach is specified, the callback is not automatically registered with the master component. The user is expected to extend from
#associate_xact_with_barrier_pair_xact, implement the association of barrier transaction with normal coherent transaction */
  } barrier_association_type_enum;

  /**
   * Enumerated type that defines the generator source for DVM complete transactions
   */
  typedef enum { 
    AUTO_DVM_COMPLETE_GEN = `SVT_AXI_AUTO_DVM_COMPLETE_GEN_SOURCE, /**< This generator_type is used by master component, when the #axi_interface_type is AXI_ACE. When this generator_type is specified, master automatically generates a DVM Complete transaction, after receiving a DVM Sync transaction. The delay between reception of DVM Sync and transmission of DVM Complete is determined by random member dvm_complete_delay*/
    USER_DVM_COMPLETE_GEN = `SVT_AXI_USER_DVM_COMPLETE_GEN_SOURCE /**< This generator_type is used by master component. When this generator_type is specified, user will need implement callback method svt_axi_master_snoop_response_gen_callback::dvm_complete_gen. The user can program the delay  dvm_complete_delay in the callback method. */
  } dvm_complete_generator_type_enum;

`endif

  /**
   * Enumerated type that defines the snoop response mode during memory update transactions
   */
  typedef enum { 
    SUSPEND_SNOOP_DURING_MEM_UPDATE = 0, /**< Master suspends incoming snoop request if memory update transaction is found in the buffer, or is active at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    SUSPEND_SNOOP_DURING_MEM_UPDATE_IN_PROGRESS = 1, /**< Master suspends incoming snoop request if memory update transaction is found to be active (addres/data phase started or about to start in current clock) at the time of receiving snoop request and provides response to that snoop request only after the current ongoing memory update transaction is complete */
    RESPOND_SNOOP_DURING_MEM_UPDATE = 2, /**< Master doesn't suspend incoming snoop request even if memory update transaction is found to be active at the time of receiving snoop request. Instead it responds to the snoop request with allowed snoop response while memory update transaction is in progress.*/ 
    EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE = 3  /**< Master either suspends incoming snoop request or respond to the snoop request while memory update transaction is in progress in a random manner.*/ 
  } snoop_response_mode_during_mem_update_type_enum;

  /**
    * 
    */
  typedef enum {
    SNOOP_RESP_DATA_TRANSFER_USING_CDDATA = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_CDDATA, /**<Transfers cache data of dirty line using CDDATA channel */
    SNOOP_RESP_DATA_TRANSFER_USING_WB_WC = `SVT_AXI_SNOOP_RESP_DATA_TRANSFER_USING_WB_WC /**<Transfers cache data of dirty line using WRITEBACK or WRITECLEAN */
  } snoop_response_data_transfer_mode_enum;

  /** enum description for various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE */
  typedef enum {
    NONSHAREABLE_XACT_FULL_ADDRESS_SPACE = 0, /**<allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE = 1, /**<allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE = 2, /**<allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
    NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE = 3 /**<allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE */
  } nonshareable_xact_address_range_in_systemshareable_mode_enum;
  typedef enum {
    STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 0,
    DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 1,
    CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES = 2 
  } source_master_id_xmit_to_slaves_type_enum;

  typedef enum {
    FALSE = 0,
    ODD_PARITY_BYTE_DATA = 1,
    ODD_PARITY_BYTE_ALL = 2
  } check_type_enum;

  /**
   * Enumerated type that defines the modifiable and non modifiable cache types
   */
  typedef enum {
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK = 0,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK = 1,
    SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_DISABLE_CHECK = 2
  } master_slave_xact_association_cache_prot_check_enum;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************
`ifndef __SVDOC__
  /** Port interface */
  AXI_MASTER_IF master_if;
  AXI_SLAVE_IF slave_if;
  AXI_PORT_STREAM_IF port_stream_if;
`endif

  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to the master/slave port corresponding
    * to this port configuration. This ID must be unique across
    * all masters/slaves of the AXI system configuration to which
    * this port belongs. A master and a slave may share the same
    * port_id, but two masters or two slaves cannot share the 
    * same port_id. If not assigned by the user, it is auto
    * assigned by the VIP. 
    */ 
  int port_id;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Name of this port. This is used in transaction short display
    * to identify the instance. This is copied over from 'inst'
    * attribute.  
    */
 local string port_name;
  /** @endcond */
  /** 
    * @groupname axi_generic_config
    * A unique ID assigned to master/slave port corresponding to this port
    * configuration. This ID must be unique across all AMBA components
    * instantiated in the testbench.  This is currently applicable only when the AMBA
    * system monitor is used and is configured using a configuration plain text
    * file (as opposed to a SystemVerilog code that sets the configuration). 
    */
  int amba_system_port_id = -1;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether output signals from master/slave IFs should be
    * initialized to 0 asynchronously at 0 simulation time. 
    * - 1: Intializes output signals from master/slave IFs to 0 
    *      asynchronously at 0 simulation time.
    * - 0: Initializes output signals from master/slave IFs to Z
    *      synchronously at 0 simulation time.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit initialize_output_signals_at_start = 1'b0;

  /** 
    * @groupname axi_generic_config 
    * Specifies whether clock should be disconnected to this agent. 
    * - 1: clock will be connected to this agent from the testbench, 
    *      based on the svt_axi_system_configuration::common_clock_mode.
    * - 0: clock will not be connected to this agent from the testbench.
    *      Used to disable the agent as per the test requirement.
    * .
    * Configuration type: Static <br>
    * Default value: 0 <br>
    */ 
  bit clock_enable = 1'b1;

  /**
    * @groupname axi_generic_config
    * Handle to the system configuration object
    */
  svt_axi_system_configuration sys_cfg;

  /**
    * @groupname axi_addr_map
    * Applicable only to slave VIP
    * Address map for this slave 
    * Must be used only if the svt_axi_system_env and svt_axi_system_configuration is not used.
    * Typically used in an environment where only one slave VIP is instantiated.
    */
  svt_axi_slave_addr_range slave_addr_ranges[];

  /**
    * @groupname axi_addr_map
    * Address map that maps global address to a local address at destination
    * Typically applicable to slave components
    * Applicable only if svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper dest_addr_mappers[];

  /**
    * @groupname axi_addr_map
    * Address map that maps a local address to a global address at a source
    * Typically applicable to master components. However, it can be applicable to
    * a slave component if that is connected downstream through another interconnect/bridge to
    * components which are further downstream. Applicable only if
    * svt_axi_system_configuration::enable_complex_memory_map is set
    */
  svt_amba_addr_mapper source_addr_mappers[];

  /**
    * @groupname axi_generic_config
    * Indicates if WID must be driven for AXI4, AXI_ACE,ACE_LITE,AXI4_LITE interfaces 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit  wid_for_non_axi3_enable = 0;

  /** 
    * @groupname axi_generic_config
    * Field for updating slave memory in request order
    * When set to 1, updates slave memory in request order that is  even though response
    * is received out of order, memory will still be updated in request order at the last
    * data phase. 
    * Default value is 0.
    * Configuration type: Static
    * Applicable only to SLAVE
    */ 
    int update_memory_in_request_order = 0;

    /**
    * @groupname axi_generic_config
    * Indicates that the monitor will check that recommended number of transactions are used      in the locked sequence 
    * Configuration type: Static
    * Applicable only to MASTER 
    */

    bit check_recommended_xact_length_for_locked_sequence = 0;
   
    /**
      * @groupname axi_generic_config
      * Indicates if X/Z checks and signal stability checks must be enabled
      * These are low level checks performed every clock and have a performance overhead
      * Often, these checks are useful only during integration phase. These can be
      * switched off after integration to get better performance.
      * These checks are automatically disabled if SVT_AXI3_4_PERF_MODE is set
      */
    bit per_clock_cycle_signal_checks_enable = 1;
 

  /**
    * @groupname axi_generic_config
    * If set to svt_axi_port_configuration::RESET_ALL_XACT,all transactions which have
    * already started along with the ones which have not yet started but are
    * present in the internal queue are ABORTED.
    * If set to svt_axi_port_configuration::EXCLUDE_UNSTARTED_XACT,only those transactions
    * which have gone out on the interface will be ABORTED.
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode because in passive mode
    * or for the slave all transactions which are in the queue are already started
    */
    reset_type_enum reset_type = `SVT_AXI_RESET_TYPE;


  /**
   * @groupname axi3_4_config
   * Indicates the way VIP reports error on receiving SLVERR or DECERR read or write response.
   * If set to svt_axi_port_configuration::NO_ERROR,vip doesn't report any error on receiving decerr
   * or slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_SLVERR,vip reports error only on receiving 
   * slverr response.
   * If set to svt_axi_port_configuration::ERROR_ON_DECERR,vip reports error only on receiving 
   * decerr response.
   * If set to svt_axi_port_configuration::ERROR_ON_BOTH,vip reports error on receiving 
   * decerr or slverr response.
   * Configuration type: Static
   *
   * This is applicable to Master in both active and passive mode and to slave only in Passive mode.
   * The default enum type of error_response_policy is NO_ERROR and is user configurable.
   */
   error_response_policy_enum error_response_policy = NO_ERROR;


  /**
    * @groupname axi_generic_config
    * Indicates if VIP would use separate address spaces for each tagged attribute. This simply means that,
    * if a coherent master or interconnect or a slave attached to such system, recieves both secure and non-secure
    * transactions then both transactions will operate on completely separate address spaces and result of one transaction
    * will not be visible to the other.
    *
    * Slave for which separate secure & non-secure address space is enabled i.e. bit [0] is set to '1', it will accept both secure
    * and non-secure transactions targeted for the same address. However, while updating memory it will use tagged address i.e. 
    * address attribute, in this case security bit, will be appended to the original address as the MSB bits.
    *
    * Slave for which separate secure & non-secure address space is disabled i.e. bit [0] is set to '0' but, configured with secured
    * regions i.e. addr_attribute[0] is set to '1' in svt_axi_slave_addr_range class via task /#set_addr_range() in system configuration
    * then it will accept only secure transactions for secure regions and all transactions for non-secure regions. 
    * With this configuration slave will use orginal address while updating memory and will not use tagged address. Hence, secure and
    * non-secure transactions to the same address will affect each other, if targeted to non-secure regions. However, if it is targeted
    * to secure regions then only secure transations will be able to update memory and access for non-secure transactions will be declined as if address doesn't exist.
    *
    * Slaves can be configured with secure region by calling /#set_addr_range(<start_addr>,<end_addr>,<addres_attribute, ex: 1 [secured]>)
    *
    * [0] => represents separate address spaces for secure and non-secure attribute if set to '1'
    * [\`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:1] => RESERVED and should be set to 0
    *
    * Configuration type: Static
    * Applicable only to MASTER 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 0;
`else    
    bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0]  tagged_address_space_attributes_enable = 1;
`endif    
    
  /**
    * @groupname axi_generic_config
    * If set to '0' then Master VIP will not drive overlapped coherent transactions on Read and Write
    * channel at the same time. WRITE transactions received by the sequencer will be blocked from being
    * sent on the interface if there is another READ transaction to an overlapping address which is 
    * already in progress. The same is true if a READ transaction is received from sequencer and a WRITE
    * transaction is in progress
    * Example: ReadShared started at 1000 ns and WriteBack received from sequencer at 1200 ns when 
    *          ReadShared is still active. At this point Master VIP will block WriteBack until ReadShared
    * is finished on the Read channel.
    *
    * If set to '1' then Master VIP will drive coherent transactions on Read and Write
    * channel as it receives from the sequencer as per other coherent rules. It will not
    * block as mentioned above. 
    * Certain scenarios that involve a store on the read channel sent out
    * speculatively while a WRITEBACK/WRITECLEAN to the same cacheline is in
    * progress require that this parameter is set to 0 so that cache states
    * reflect correctly. 
    * If snoop_response_data_transfer_mode is set to
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, this parameter must be set to 1 to
    * facilitate the transfer of snoop data on the write channel without
    * getting blocked.
    *
    * Configuration type: Static
    *
    * This is applicable to only the Master in active mode 
    */
    bit allow_overlapped_read_and_write_channel_coherent_transactions = 0;    
   
   /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP can drive random snoop response for
    * WasUnique (BRRESP[4]) even if the snoop_initial_cache_line_state is in 
    * UNIQUE state.
    * If set to '0' the Master VIP must set WasUnique (BRRESP[4]) to 1 if
    * the snoop_initial_cache_line_state is UNIQUE.
    */ 
    bit allow_was_unique_zero_in_unique_state = 1; 
   
   /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * If set to '1' then Master VIP will allow burst_size to be less than
    * data_width for Atomic transaction.
    * If set to '0' then Master VIP will throw an is_valid error when burst_size 
    * is less than data_width for Atomic transaction.
    * This is only applicable for multibeat atomic transactions. 
    */
    bit allow_multibeat_atomic_transactions_to_be_less_than_data_width = 0;   
    /** @endcond */

   /**
    * @groupname axi_generic_config
    * This is applicable only when interconnect VIP is used, this is
    * applicable for all transactions. 
    * So if set to 1, then the interconnect VIP will always update dirty data into main memory 
    * if it receives dirty data from snoops corresponding to a transaction from this port
    */
    bit memory_update_for_pass_dirty_enable = 0;
 
   /**
    * @groupname axi_generic_config
    * This is applicable only when interface_type is AXI3 or AXI4
    * If set to 1 and axi_interface_type is AXI3/AXI4, system monitor will update
    * the port_configuration member axi_interface_type as ACE_LITE .
    * In addition to that system monitor will update svt_axi_transaction::xact_type as COHERENT.
    */

    bit is_downstream_coherent = 1'b0;

  /** @cond PRIVATE */
  /** Helper attribute for specifying solve order */
  local rand bit primary_props;

  /** holds total number of enabled tagged address space attributes */
  local int      num_enabled_tagged_addr_attributes = 0;

  /** Supports four state memory
   *  Default value is set as 0
   *  If set as 1 supports 4 state memory.
   */

  bit is_4state = 1'b0;
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  /** 
   * @groupname axi3_4_generator
   * The source for the stimulus that is connected to the transactor.
   *
   * Configuration type: Static
   */
  generator_type_enum generator_type = SCENARIO_GEN;

  /**
   * @groupname ace_generator
   * The source type for snoop response generation.
   *
   * Configuration type: Static
   */
  snoop_response_generator_type_enum snoop_response_generator_type = CACHE_SNOOP_RESPONSE_GEN;

  /**
   * @groupname ace_config
   * Defines how a transaction is associated with a barrier transaction pair.
   *
   * Configuration type: Static
   */
  barrier_association_type_enum barrier_association_type = RANDOM_ASSOCIATION;

  /** 
    * @groupname ace_generator
    * Defines how DVM complete transactions need to be generated.
    *
    * Configuration type: Static
    */
  dvm_complete_generator_type_enum dvm_complete_generator_type = AUTO_DVM_COMPLETE_GEN;

  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_scenarios = -1;

  /**
    * @groupname axi_generic_config
    * The number of instances that the generators should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int stop_after_n_insts = -1;

  // ACE
  /** 
    * @groupname axi_generic_config
    * The number of scenarios that the snoop_generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_scenarios = -1;

  /** 
    * @groupname axi_generic_config
    * The number of instances that the snoop generator should create for each test
    * loop.
    *
    * Configuration type: Static
    */
  int snoop_stop_after_n_insts = -1;

`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in UVM_LOW verbosity.
    */
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_HIGH verbosity.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in OVM_LOW verbosity.
    */
`else
  /**
    * @groupname axi_generic_config
    * When silent_mode is set to 1, the "Transaction started" and 
    * "Transaction ended" messages are printed in DEBUG_SEV.
    * When silent_mode is set to 0, the "Transaction started" and 
    * "Transaction ended" messages are printed in NORMAL_SEV.
    */
`endif
  bit silent_mode  = 0;

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`elsif SVT_OVM_TECHNOLOGY
  /** 
    * @groupname axi_generic_config
    * Specifies if the agent is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables sequencer, driver and 
    * monitor in the the agent. 
    * - 0: Configures component in passive mode. Enables only the monitor in the agent.
    * - Configuration type: Static
    * .
    */
`else
  /**
    * @groupname axi_generic_config
    * Specifies if the group is an active or passive component. Allowed values are:
    * - 1: Configures component in active mode. Enables driver, generator and
    * monitor in the group component. 
    * - 0: Configures component in passive mode. Enables only the monitor in the group component.
    * - Configuration type: Static
    * .
    */
`endif
  bit is_active = 1;
  
  /** @cond PRIVATE */
  /** xml_writer handle of the agent */
  svt_xml_writer xml_writer = null;
  /** @endcond */


  /** 
    * @groupname axi_generic_config
    * The AXI interface type that is being modelled. Please note that interface
    * type AXI_STREAM is not yet supported.
    * Configuration type: Static
    */
  rand axi_interface_type_enum axi_interface_type = AXI3;

  /** 
    * @groupname axi3_4_config
    * The AXI4 interface category (read-only, write-only, read-write) of this interface. 
    * Configuration type: Static
    */ 
  rand axi_interface_category_enum axi_interface_category = AXI_READ_WRITE;

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a master or a slave. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is of kind master or slave.
    */ 
  axi_port_kind_enum axi_port_kind = AXI_MASTER;

  /**
    * Specifies the impact of svt_axi_transaction::force_xact_to_cache_line_size 
    * based on the axi_interface_type. 
    * 
    * Applicable only for ACTIVE master.
    */
  force_xact_to_cache_line_size_interface_type_enum force_xact_to_cache_line_size_interface_type = ALL_INTERFACE_TYPES;

 /** 
   * @groupname ace5_config
   * Indicates supported version  of ACE specefication by AMBA AXI_ACE VIP
   * Default value of this parameter is ace_version_1_0.User need to set this parameter if they wish to
   * to use new ACE spec which is ACE spec version 2.0
   * Configuration type:static
   */
   ace_version_enum ace_version = ACE_VERSION_1_0;

/** 
   * @groupname ace5_config
   * Indicates cache stashing feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cache_stashing_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates if trace signal feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit trace_tag_enable = 0;

/** 
   * @groupname ace5_config
   * Indicates whether the trace tag value will be directly reflected in the response packet or spawned packets generated in response to the received packet.
   * when set to 1: The trace_tag value will be directly mapped to the associated response and spawned packets, irrespective of trace_tag value being 0 or 1 in the request.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 and svt_axi_port_configuration::trace_tag_enable is set to 1.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit loopback_trace_tag_enable = 0;

`ifdef SVT_ACE5_ENABLE 
/** 
   * @groupname ace5_config
   * Indicates if atomic transactions feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit atomic_transactions_enable = 0;


 /** 
   * @groupname ace5_config
   * Indicates if write_with_cmo feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit write_plus_cmo_enable = 0;
 
 /** 
   * @groupname ace5_config
   * Indicates if cmo transactions can be sent on the write channel.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit cmo_on_write_enable = 0;

 /**@groupname ace5_config
   * Specifies the number of outstanding Atomic transactions a port can support.<br>
   * This is applicable only for ACE5 ports with atomic_transactions_enable set to 1.<br>
   * The Atomic transactions include:
   * - AtomicStore
   * - AtomicLoad
   * - AtomicSwap
   * - AtomicCompare
   * .
   * MASTER:
   * If the number of outstanding atomic transactions is equal to this
   * number, the slave will refrain from initiating any new 
   * transactions until the number of outstanding write transactions
   * is less than this parameter.<br>
   * SLAVE:
   * If the number of outstanding transactions is equal to 
   * this number, the slave will not assert ARREADY/AWREADY
   * until the number of outstanding transactions becomes less
   * than this parameter. 
   * <br>
   * This parameter must be set if #num_outstanding_xact = -1.
   * This parameter must not be set if #num_outstanding_xact is not set to -1.
   * - <b>Default val:</b> -1
   * - <b>min val:</b> 1
   * - <b>max val:</b> Value defined by macro \`SVT_AXI_MAX_NUM_OUTSTANDING_XACT.
   * - <b>type:</b> Static
   * .
   */
  rand int num_outstanding_atomic_xact = 1;

 /** 
   * @groupname ace5_config
   * Indicates if Memory Partitioning and Monitoring (MPAM) feature is supported.
   * It can be set to either of two values below:
   *    enable_mpam = svt_axi_port_configuration:FALSE
   *  When set to FALSE, MPAM is not supported on the interface.
   *    enable_mpam = svt_axi_port_configuration:MPAM_9_1
   *  When set to MPAM_9_1, MPAM is supported on the interface with mpam_partid_width=9 and mpam_perfmongroup_width=1. 
   *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * - Default value:FALSE, is controlled through user re-definable macro `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM.
   * .
   */
   mpam_support_type_enum enable_mpam = `SVT_AXI_PORT_CFG_DEFAULT_ENABLE_MPAM;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Partition identifier.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_partid_width = 9;

 /** 
   * @groupname ace5_config
   * Indicates the width of MPAM Performance monitor group.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   rand int mpam_perfmongroup_width = 1;

`endif
  /**
   * @groupname ace5_config
   * If set to 1, it will enable the master component to support deallocating transactions.
   * By default, the value of this parameter is 0. This means it can not support deallocating
   * transactions and any READONCEMAKEINVALID or READONCECLEANINVALID transaction initiated
   * from this master component will be converted to READONCE transaction.
   *
   * Applicable only when svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   * and svt_axi_port_configuration::axi_interface_type is set to ACE_LITE
   * Configuration type:static
   */
   bit deallocating_xacts_enable = 0;



  /** 
   * @groupname ace5_config
   * Indicates address translation feature is supported by this port.
   * Can be set to 1 only when the compile macro SVT_ACE5_ENABLE is defined and
   * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0.
   * - Configuration type: Static
   * - Default value:0.
   * .
   */
   bit addr_translation_enable = 0; 

  /**
    * @groupname axi_generic_config
    * Indicates whether this port is a interconnect VIP port or not. User does not need to
    * configure this parameter. It is set by the VIP to reflect whether the port
    * represented by this configuration is a port of interconnect VIP or not.
    * .
    */  
  bit is_ic_port = 0;
  
 /**
   * @groupname axi_generic_config
   * Indicates if the port_monitor protocol check max_num_outstanding_xacts_check 
   * is enabled or not .The max_num_outstanding_xacts_check checks that AXI master and AXI slave 
   * are not exceeding the user configured maximum number of outstanding transactions (#num_outstanding_xact).   
   * If #num_outstanding_xact = -1 then #num_outstanding_xact will not be considered , 
   * instead #num_read_outstanding_xact and #num_write_outstanding_xact will be considered for read and write transactions respectively.
   */
  bit max_num_outstanding_xacts_check_enable =0; 
 
  /** @groupname axi_generic_config
    * Disable the association between slave read transaction and master partial write transaction.
    * This covers the specefic scenario when master partial write transaction is split into
    * slave read transaction followed by a slave write transaction by the ICN.
    * If set to 1 association between master write transaction and slave read transaction is done by the system monitor.
    * If set to 0 association between master write transaction and slave read transaction is not done by the system monitor.
    */
  bit partial_write_to_slave_read_and_write_association_enable = 0;
 
 /**
   * @groupname axi_generic_config
   * Indicates if this port is interleaved based on address to be accessed by this port
   */
  bit port_interleaving_enable =0;  
 
/** Indicates the port interleaving boundary. The value must be in form of bytes.
  * For example if interleaving szie is 64 . It means interleaving boundary os 64 bytes.
  * This port will access address locations based on interleaving size.
  * Default value is set as 64.
  * Applicable if the port_interleaving_enable is set to 1 for this port.
  */
  int port_interleaving_size = 64;

/** Indicates the group id of all the ports participating in one interleaving scheme
  * All the ports which are in the same interleave group must be configured to have same 
  * port_interleave_group_id
  * Default is set to -1 . 
  * Applicable if the port_interleaving_enable is set to 1.
  * Its value must be unique across master and slaves .All the port_ids having same port_interleaving_group_id
  * must be contigous.
  */
  int port_interleaving_group_id = -1;

/** Indcates that DVM transactions will be sent form this port of corresponding port interleaving group
  * This port will not take part in port interleaving for DVM transactions 
  * Applicable if port_interleaving_enable is set to 1.
  */
  bit dvm_sent_from_interleaved_port = 0;

/**Indicates that non coherent device traffic will be sent from this port
  * of corresponding port interleaving group.
  * This port will not take part in port interleaving for device traffic
  * as Device transaction addresses are not interleaved.
  * Applicable only when the port_interleaving_enable is set to 1.
  */ 
  bit device_xact_sent_from_interleaved_port =0;

/**  Indicates the order of this port in a port interleaving scheme.
  *  For example : If the port is 3rd in a group of 4 ports .If port_interleaving_size of the group is 512 bytes
  *  This port will have access to addresses with addr[10:9] == 3.
  *  This parameter determines which address bits to look for an interleaved port.
  *  Default value of this is set to 0 
  */
   int port_interleaving_index = 0;

  /**
   * @groupname axi_generic_config
   * Enables port inteleaving for this port for the device type xact.
   * The port configuration parameter device_xact_sent_from_interleaved_port
   * is not applicable if this bit is set to 1.
   * If this bit is set to 1, the device type transaction is interleaved like 
   * any non-dvm transaction.
   */
  bit port_interleaving_for_device_xact_enable = 0;

  /**
    * Indicates if this port  supports the setting of Poison field. <br>
    * - Default value: 0.
    * .
    */
  bit poison_enable = 1'b0;

   /** 
    * @groupname axi_generic_config
    * Indicates if the transactions on this port must be processed by the axi
    * system monitor. This configuration is applicable only to the
    * 'system_monitor' of the instance of svt_axi_system_env within which the
    * component corresponding to this port configuration is instantiated.
    * It is not used in the AMBA system monitor instantiated in an instance of
    * svt_amba_system_env (system env used when multiple AMBA protocols are
    * used)
    */ 
  bit connect_to_axi_system_monitor = 1;

  /** @cond PRIVATE */
  /**
    * @groupname axi_generic_config
    * Indicates that, if this bit is set to '1' then user needs to externally push
    * coherent and snoop master transactions and slave transactions into the port monitors. 
    * port monitor will not automatically sample it's related interface and hence will not
    * create corresponding transactions and instead will use the user provided transaction handle
    * externally pushed into the monitor.
    */ 
  bit use_external_port_monitor = 0;
  /** @endcond */

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates a tlm_generic_payload_sequencer sequencer capable
    * of generating UVM TLM Generic Payload transactions and connects the
    * master sequencer to it.  The master sequencer starts a layering sequence that gets
    * transactions from the tlm_generic_payload_sequencer, converts them to (one or more) AXI
    * transaction(s) and sends them to the driver.
    * Snoop requests are still fulfilled by the svt_axi_master_snoop_sequencer.
    * 
    * AXI transactions observed by the agent
    * are also made available as TLM GP transactions through the
    * tlm_generic_payload_observed_port in the monitor. Note that the TLM GP
    * transactions issued through the analysis port may not match one to one with GP
    * sequence items created by the tlm_generic_payload_sequencer because the
    * GP sequence items may have to be mapped
    * to multiple AXI transactions according to protocol requirements. The
    * TLM GP that is available through the tlm_generic_payload_observed_port of
    * the monitor is a direct mapping of the observed AXI transactions converted to a TLM GP.
    * No attempt is made to re-assemble a set of AXI transaction into a larger TLM GP.
    * 
    * The layering sequence that converts the TLM GP to AXI transactions is the
    * svt_axi_tlm_gp_to_axi_sequence and is available at
    * $DESIGNWAREHOME/vip/svt/amba_svt/<ver>/axi_master_agent_svt/sverilog/src/vcs/svt_axi_tlm_gp_sequence_collection.svp 
    * Transactions created by the layering sequence are of type
    * cust_svt_tlm_gp_to_axi_master_transaction. Any user constraints specific
    * to AXI must be provided in a class extended from this class.
    * 
    * In passive mode, observed AXI transactions are made available as TLM GP
    * transactions through the tlm_generic_payload_observed_port in the
    * monitor.
    */
  bit use_tlm_generic_payload = 0;

  /** 
    * @groupname axi_tlm_generic_payload
    * In active mode, creates an AMBA-PV-compatible socket that can be used to
    * connect AXI Master VIP component to an AMBA-PV master model. 
    * 
    * Enabling this functionality causes the instantiation of socket b_fwd of
    * type uvm_tlm_b_target_socket, and socket b_snoop of type
    * uvm_tlm_b_initiator_socket, in class svt_axi_master_agent.

    * Generic payload transactions received through the forward b_fwd interface
    * are executed on the tlm_generic_payload_sequencer in the agent.

    * When this option is set, the svt_axi_ace_snoop_request_to_tlm_gp_sequence
    * reactive sequence is started on the AXI VIP master snoop sequencer. Snoop
    * transaction requests received by the AXI VIP master snoop sequencer are translated to
    * equivalent tlm_generic_payload transactions with the
    * #svt_amba_pv_extension attached. The extended Generic Payload transactions
    * are then sent to the AMBA-PV master model via the backward b_snoop interface.
    * The receive response from AMBA-PV master model is then interpreted to
    * complete the snoop transaction request and executed on the AXI VIP master snoop
    * sequencer.
    * 
    * Should the AXI VIP master fulfill the snoop requests natively (i.e. the
    * default behavior when this option is not set), the snoop response sequence
    * should be restored to the default using:
    * 
    * <code>
    * uvm_config_db#(uvm_object_wrapper)::set(this, "master[0].snoop_sequencer.run_phase", "default_sequence",
    *                                         /#svt_axi_ace_master_snoop_response_sequence::type_id::/#get());
    * </code>
    * 
    * When this option is set, it implies that #use_tlm_generic_payload is also set, whether
    * it actually is or not.
    */
  bit use_pv_socket = 0;

 /** Enables the UVM REG feature of the AXI agent.  
   * Applicable only when svt_axi_port_configuration::axi_interface_type is AXI3.
   * <b>type:</b> Static 
   */
  bit uvm_reg_enable = 0;

 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables checking of wdata/tdata only on valid byte lanes based on wstrb/tstrb. 
    * In a disabled state, whole wdata/tdata as seen on the bus will be considered.
    * <b>type:</b> Dynamic 
    */
  bit check_valid_data_bytes_only_enable = 1;

  /**
    * @groupname axi3_4_timeout_config
    * A timer which is started when a transaction starts. If the transaction
    * does not complete by the set time, an error is repoted. The timer is
    * incremented by 1 every clock and is reset when the transaction ends. 
    * If set to 0, the timer is not started
    */
  int xact_inactivity_timeout = 0;

 /**
   * @groupname ace_config 
   * If this attribute is enabled it will allow snoop response data_transfer bit for
   * MAKEINVALID  transaction to be set as 1. This behaviour is permitted by protocol
   * but it is not expected snoop response for MAKEINVALID 
 */
  bit  data_transfer_for_makeinvalid_snoop_enable =0;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /** 
   * log_base_2 of \`SVT_AXI_MAX_DATA_WIDTH. 
   * Used only as a helper attribute to randomize data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_data_width;
 
  /** 
   * log_base_2 of \`SVT_AXI_ACE_SNOOP_DATA_WIDTH. 
   * Used only as a helper attribute to randomize snoop_data_width.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_snoop_data_width; 

  /** 
   * log_base_2 of \`SVT_AXI_MAX_CACHE_LINE_SIZE. 
   * Used only as a helper attribute to randomize cache_line_size.
   *
   * This parameter is not required to be set by the user.
   */
  int log_base_2_max_cache_line_size;

  /**
    * Indicates if the address range of the slave component
    * has been set
    */
  bit is_slave_addr_range_set = 0;

  /**
    * Stores the log_base_2 of the desired data_width.
    * Used only as a helper attribute to randomize data_width.
    * This parameter is first randomized and the data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_data_width;

  /**
    * Stores the log_base_2 of the desired snoop_data_width.
    * Used only as a helper attribute to randomize snoop_data_width.
    * This parameter is first randomized and the snoop_data_width
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_snoop_data_width;

  /**
    * Stores the log_base_2 of the desired cache_line_size.
    * Used only as a helper attribute to randomize cache_line_size.
    * This parameter is first randomized and the cache_line_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_cache_line_size;

  /**
    * Stores the log_base_2 of the desired atomicity_size.
    * Used only as a helper attribute to randomize atomicity_size.
    * This parameter is first randomized and the atomicity_size
    * is constrained to its power of 2 value.
    * <b>type:</b> Static
    *
    * This parameter is not required to be set by the user.
    */
  rand int log_base_2_atomicity_size;

  /** @endcond */

  /** 
    * @groupname axi3_signal_width
    * Address width of this port in bits.
    * When svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE,
    * this parameter also sets the width of signal caddr.
    *
    * NOTE: currently same address width is considered for both coherent read or write address
    *       channels and snoop address channels. So, there is no separate snoop address width
    *       parameter supported at the moment.
    * Configuration type: Static
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE 
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH;
`else    
  rand int addr_width = `SVT_AXI_MAX_ADDR_WIDTH - `SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH;
`endif   

  /** 
    * @groupname axi4_signal_width
    * Address user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int addr_user_width = `SVT_AXI_MAX_ADDR_USER_WIDTH;

  /** 
    * @groupname axi3_signal_width
    * Data width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_width = `SVT_AXI_MAX_DATA_WIDTH;

  /** 
    * @groupname axi4_signal_width
    * Data user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int data_user_width = `SVT_AXI_MAX_DATA_USER_WIDTH;
 
  /** 
    * @groupname axi4_signal_width
    * Response user width of this port in bits.
    *
    * Configuration type: Static
    */
  rand int resp_user_width = `SVT_AXI_MAX_BRESP_USER_WIDTH;

  /** 
    * @groupname ace_config
    * Cache line size in bytes for this master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int cache_line_size = `SVT_AXI_MAX_CACHE_LINE_SIZE;

  /** 
    * @groupname ace_config
    * Aligned size in bytes for the snoop corresponding to starting address.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates the size to which the snoop corresponding to the starting address
    * of a multi-cacheline access is aligned. For example, if the cacheline size
    * is 64 bytes and the coherent address of a READONCE transaction is 0x70,
    * the corresponding snoop address may be 0x40 or 0x70. If the snoop address
    * sent is 0x40, this value must be set to the same as the cacheline size which is
    * 64 bytes. If the snoop address sent is 0x70, this value can be set to 16 bytes.
    * This will help in more accurate correlation of coherent and snoop transactions.
    * The default is 0. If unchanged, the system monitor will use the cacheline size
    * for this value, assuming that all snoops are aligned to cacheline size. 
    * Configuration type: Static
    */
  rand int start_addr_snoop_aligned_size = 0;

  /** 
    * @groupname ace_config
    * Number of cache lines in the master.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int num_cache_lines = `SVT_AXI_MAX_NUM_CACHE_LINES;

  /** 
    * @groupname ace_config
    * Enables AWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default AWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit awakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Enabling this feature will allow transactions to wait to send address phase
    * until the previous transaction's datahandshake is done. This will result
    * in unexpected delays. Hence this parameters is disabled by default.
    * 
    * This parameter is applicable when 
    * svt_axi_port_configuration::axi_interface_type is set to AXI3 or AXI4.
    *
    * Configuration type: Static
    */
  rand bit prev_xact_data_handshake_ref_event_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles AWAKEUP sideband signal in the VIP during idle period of read or
    * write channel.
    * Asserts and then de-assert AWAKEUP with the range of programed number of 
    * 'awakeup_toggle_min_delay_during_idle' to 'awakeup_toggle_max_delay_during_idle'.
    * If there is no transaction observed in read or write channel, then AWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int awakeup_toggle_max_delay_during_idle = 5;


  /** 
    * @groupname ace_config
    * Enables ACWAKEUP sideband signal in the VIP when this bit is set to '1'.
    * by default ACWAKEUP signal will be '0' when this bit is enabled.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand bit acwakeup_enable = 0;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_min_delay_during_idle = 1;

  /** 
    * @groupname ace_config
    * Toggles ACWAKEUP sideband signal in the VIP during idle period of snoop channel.
    * Asserts and then de-assert ACWAKEUP with the range of programed number of 
    * 'acwakeup_toggle_min_delay_during_idle' to 'acwakeup_toggle_max_delay_during_idle'.
    * If there is no snoop transaction observed in snoop channel, then ACWAKEUP
    * will be toggled with respect to programmed number of delays. 
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Configuration type: Static
    */
  rand int acwakeup_toggle_max_delay_during_idle = 5;
  
  /** 
    * @groupname ace_signal_width
    * Snoop Data width of the cddata port in bits.
    * This parameter is applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Configuration type: Static
    */
  rand int snoop_data_width = `SVT_AXI_ACE_SNOOP_DATA_WIDTH;

  /**
    * @groupname axi3_4_config
    * Acronym for "What You See is What You Get". Applicable to the
    * svt_axi_transaction::data and svt_axi_transaction::wstrb fields of a
    * transaction. If this bit is set to 1, whatever is configured in the
    * svt_axi_transaction::data and  svt_axi_transaction::wstrb fields is
    * transmitted "as is" by the master. Also, in the transaction object
    * generated by monitor, the monitor populates the svt_axi_transaction::data
    * and  svt_axi_transaction::wstrb fields "as is", as seen on the bus. If
    * this bit is set to 0 (default), the data must be stored right-justified by
    * the user. The model will drive the data on the correct lanes.
    *
    * Refer to the documentation of svt_axi_transaction::data and 
    * svt_axi_transaction::wstrb for more details
    */
  rand bit wysiwyg_enable = 0;

  /**
    * @groupname axi3_4_config
    * Applicable when #wysiwyg_enable is set.
    * Indicates if the VIP should consider validity of wstrb in transactions
    * when #wysiwyg_enable is set. When wysiwyg_enable is set, the driver
    * checks that #wstrb is set only for valid byte lanes of each beat.  In
    * certain applications, wstrb may have to be asserted for other byte lanes
    * as well. In such applications, this bit should be set. This results in
    * the following: 
    * <br>
    * Constraints in transaction are relaxed for wstrb. wstrb
    * values will be random and may be asserted for invalid byte lanes. 
    * <br>
    * driver does not check for validity of wstrb in transaction based on valid
    * byte lanes.
    * <br>
    * Note that this will result in a non-AXI compliant behaviour, in that
    * wstrb may be asserted for invalid byte lanes based on what the user
    * programs. If this bit is set for the slave, and if the user wants memory
    * to be updated based on the transactions, the memory sequence shipped with
    * the VIP should not be used. For VMM based testbenches, the generator_type
    * should not be set to MEMORY_RESPONSE_GEN. This is because the APIs that
    * access memory are based on valid assertion of byte strobes.  The user
    * must use user-defined APIs and sequences to access memory if this bit is
    * set in the slave.
    */ 
  bit ignore_wstrb_check_for_wysiwyg_format = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal on byte count calculation in the VIP 
    * By default this configuration parameter is set to 0 to calculate the byte count using burst_size and burst_length,
    * if this parameter is set 1 then wstrb is used to calculate the byte count
    * <b>type:</b> Static
    */
  rand bit get_byte_count_from_wstrb_enable      = 0;

   /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWREGION signal in the VIP 
    * <b>type:</b> Static
    */

  rand bit awregion_enable   = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARREGION signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arregion_enable   = 0;
 
  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the AWQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit awqos_enable      = 0;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wlast_enable      = 1;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the WSTRB signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit wstrb_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the BRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit bresp_enable      = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arid_enable       = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLEN signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlen_enable   = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARSIZE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arsize_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARBURST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arburst_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARLOCK signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arlock_enable     = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARCACHE signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arcache_enable    = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARPROT signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arprot_enable     = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the ARQOS signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit arqos_enable      = 0;

  /** @cond PRIVATE */
  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RID signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rid_enable        = 1;

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RRESP signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rresp_enable      = 1;
  /** @endcond */

  /** 
    * @groupname axi4_signal_enable
    * Signifies the presence of the RLAST signal in the VIP 
    * <b>type:</b> Static
    */
  rand bit rlast_enable      = 1;

  /** 
    * @groupname axi3_4_config
    * Enables AWUSER sideband signal in the VIP. AWUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit awuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables WUSER sideband signal in the VIP. WUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit wuser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables BUSER sideband signal in the VIP. BUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit buser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables ARUSER sideband signal in the VIP. ARUSER signal can be used when
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit aruser_enable      = 0;

  /** 
    * @groupname axi3_4_config
    * Enables RUSER sideband signal in the VIP. RUSER signal can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * <b>type:</b> Static
    */
  rand bit ruser_enable      = 0;

  `ifdef SVT_AXI_QVN_ENABLE
  /** 
    * @groupname axi_qvn_config
    * Enables QVN support in the VIP. QVN signals can be used when 
    * svt_axi_port_configuration::axi_interface_type is set to
    * AXI3/AXI4/AXI4_LITE/AXI_ACE/ACE_LITE. 
    * All QVN configuration parameters comes into effect only when qvn_enable bit is set.
    * Any parameter which is declared as a bit-vector to support all Virtual Network in the
    * system, is sized by `define macro "SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK".
    *
    * If a system should support a maximum number of 5 Virtual Networks then user should
    * define SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK as 5
    * <b>type:</b> Static
    */
  rand bit qvn_enable      = 0;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Read Address channel
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_ar_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Specifies how many Virtual Network a particular master supports for Write Address channel.
    * Write Data channel must support Virtual Networks same as Write Address channel so there is
    * no need of having seperate configuration for Write Data channel.
    * <b>type:</b> Static
    */
  rand int qvn_num_virtual_network_supported_aw_chnl = 1;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Read-Address Channel.
    * It provides an array of bits each representing a Virtual Network in the system. Index of 
    * each bit denotes ID of the Virtual Network, represented by that bit.
    * If any bit of this array is set to '1' then that means Virtual Network with ID equal to
    * index of that bit, is supported by this port. If a bit in this array is set to '0' then
    * that means Virtual Network with ID equal to its index is not supported by this port.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 1 and 3 to be used for its
    *           Read-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_ar_chnl[index]) qvn_supported_virtual_network_queue_ar_chnl[index] = 0; 
    *   set '1' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_ar_chnl[1] = 1;
    *   set '1' for Virtual Network 3 =>  qvn_supported_virtual_network_queue_ar_chnl[3] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_ar_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /** 
    * @groupname axi_qvn_config
    * Lists Virtual Networks which are supported by a master/slave port for Write Address Channel.
    * This array of bits also indicate which Virtual Networks are supported by this port similar
    * to the array qvn_supported_virtual_network_queue_ar_chnl described above.
    * Initial Value:  all bits are set to '0' i.e. no Virtual Network is supported by default.
    * Example:  If a port must be configured to use Virtual Network 0 and 2 to be used for its
    *           Write-Address channel then user should configure as follows:
    *   (manual configuration without randomization)  - reset all bits to '0'
    *   foreach(qvn_supported_virtual_network_queue_aw_chnl[index]) qvn_supported_virtual_network_queue_aw_chnl[index] = 0; 
    *   set '0' for Virtual Network 1 =>  qvn_supported_virtual_network_queue_aw_chnl[1] = 1;
    *   set '1' for Virtual Network 2 =>  qvn_supported_virtual_network_queue_aw_chnl[2] = 1;
    */
  rand bit qvn_supported_virtual_network_queue_aw_chnl[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] ;

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on read address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */

   /* If a Master is not able to use a token, then after this timelimit that token will be reclaimed
    * by the slave which, granted it and Master will remove this token from its reserved token pool.
    *
    * - So, it is important to set suitable value for this parameter. If it is set too low, then
    * most tokens may expire before it could be used and hance leading to increased token request.
    *
    * - If it is set below minimum no. of cycles a master needs to use a token then all tokens will
    * expire and none could be used to issue a transaction to AXI channels.
    *
    * - On the other hand if it uses too high value, then due to under usage of token or over-request
    * of tokens by a Master, there is a possibility of accumulating large number of tokens in the
    * token-pool of that master and hence causing possible blockage to other masters.
    *
    * - If it is set to Zero then that indicates there is no timelimit for token usage i.e. once a 
    * token is acquired it will remain in the token-pool of that master until used for sending a
    * transaction.
    * .
    */
  rand int qvn_read_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write address channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_addr_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies maximum number of clock cycles (interface clock) within which a Master must use
    * all the tokens it has been granted on write data channel.
    * Port Monitor uses this parameter to assert warning if Master didn't use its granted token 
    * within this bounded time period.
    */
  rand int qvn_write_data_token_usage_timelimit[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Read Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AR_PRE_ALLOCATED_TOKEN
    * Example: if AR channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_ar_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_ar_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Pre-Allocated Token for Write Address Channel
    * An integer array is provided to hold pre_allocated token number for AR channel of
    * each corresponding Virtual Network. Index of an array element indicates for which
    * virtual network it holds pre_allocated token number.
    * Initial Value : all elements of this array is initiallized to \`SVT_AXI_QVN_MIN_NUM_AW_PRE_ALLOCATED_TOKEN
    * Example: if AW channel of Virtual Network 2 should be set to 1 then configure as
    *   qvn_num_aw_pre_allocated_token_vn[2] = 1;
    */
  rand int qvn_num_aw_pre_allocated_token_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Indicates if same AXI ID can be used between two different Virtual Network or not.
    * - If set to "0" then at any given point of time no two different Virtual Networks will
    * use same ID for transactions sent to AXI channels associated with those VNs.
    * - if set to "1" then same AXI ID can be used by two different VN without any restriction.
    * .
    *
    * NOTE: if same ID is used for AXI transactions issued to two different VN may get
    * blocked by interconnect in order to observe AXI ID ordering rule. Because of this, a
    * transaction received first will block another transaction with same ID received later,
    * even if transaction that was received first, can't make any progress.
    */
  rand int qvn_allow_id_used_in_other_vn = 0;

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on read address channel. It helps in defining how system resources will be used
    * otherwise, a master can issue large number of token requests and once granted those tokens 
    * may remain unused reserving system resources and in turn blocking other masters, if it shares 
    * same Virtual Network or if slave uses shared token for different masters.
    * 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_read_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write address channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_addr_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of granted token a master can keep unused for each virtual network
    * it supports on write data channel. 
    * NOTE: by default it is randomized within range [\`SVT_AXI_QVN_NUM_MIN_ALLOWED_UNUSED_TOKEN:\`SVT_AXI_QVN_NUM_MAX_ALLOWED_UNUSED_TOKEN]
    * 
    */
  rand int qvn_max_num_write_data_unused_token[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for read address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for read address channel.
    */
  rand int unsigned qvn_ar_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write address channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write address channel.
    */
  rand int unsigned qvn_aw_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of clock cycles (interface clock) within which slave must assert ready
    * to the master requesting token for write data channel. If slave doesn't assert ready i.e.
    * grant token to the master within this specified clock cycles then timeout will occur and
    * error will be asserted. Master driver waiting for the ready will also come out and abort
    * the transaction.
    *
    * NOTE: if this timeout value is set to '0' then timeout will be disabled and master will
    * wait forever until token request ready is asserted by slave for write data channel.
    */
  rand int unsigned qvn_w_token_request_ready_timeout_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];


  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AR channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AR channel
    */
  rand int qvn_slave_ar_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for AW channel for a particular Virtual Network
    * This means Slave has these many token resources to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Since Master is pre-allocated with certain number of token Slave will begin with 
    *       number of Tokens as specified here minus master pre_allocated_token for AW channel
    */
  rand int qvn_slave_aw_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies number of Token Slave can have for W channel for a particular Virtual Network
    * This means Slave has this many token resource to allocate to Master and can't give token
    * more than the value specified here.
    * Note: Master doesn't have any pre-allocated token for Write Data channel so, Slave will 
    *       begin with same number of Tokens as specified by this parameter.
    */
  rand int qvn_slave_w_token_size_for_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for read address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_rd_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write address channal for a VN, 
    * in accordance with slaves acceptance capability.
    * Note: This is exclusive of pre allocated token for the VN  
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_addr_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /**
    * @groupname axi_qvn_config
    * Specifies max number of outstanding token request slave can grant for write data channal for a VN, 
    * in accordance with slaves acceptance capability.
    */
   rand int unsigned qvn_slave_max_outstading_token_for_wr_data_chan_vn[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

   /**
    * @groupname axi_qvn_config
    * Mode to control the assertion of V*READYVNx signal. This allows QVN enabled Slaves to assert
    * token request grant ready signal for any Virtual Network of each channel AR, AW, W
    *
    * 0 - Assert V*READY in responce to assertion of V*VALID for token request 
    * 1 - Assert V*READY before assertion of V*VALID for token request, subjected to token availability
    */  
   rand bit qvn_slave_aw_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_assertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_assertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
  
   /*
    * @groupname axi_qvn_config
    * Mode to control the de-assertion of V*READYVNx signal. This flage is only 
    * applicable if v*ready_assertion_mode is set to ONE.
    * 0 - Keep V*READY till assertion of V*VALID.  
    * 1 - Deassert V*READY after some time if V*VALID is not asserted. 
    */  
   rand bit qvn_slave_aw_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_w_ready_deassertion_mode  [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};
   rand bit qvn_slave_ar_ready_deassertion_mode [`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1:0] = '{`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK {0}};


  `endif

  /** 
    * @groupname axi3_4_config
    * Enables optimistic flow control for Write Data channel in the VIP.  
    * The flow control of the write data channel is determined by the settings 
    * in num_outstanding_xact and num_outstanding_write_xact. Based on these 
    * settings wready is deasserted when the number of outstanding transactions
    * reach the threshold set by these parameters. This parameter controls the 
    * deassertion of wready when the threshold is reached. Since AXI allows data 
    * before address, a new transaction can start with data. When this parameter 
    * is disabled, both awready and wready are deasserted when threshold of maximum
    * outstanding transactions are reached. Note however that this will prevent data
    * of any already outstanding transactions from being continuously accepted
    * (that is with wready continuously high) and therefore can reduce throughput
    * If this parameter is set, only awready is deasserted when the threshold is reached.
    * This allows data of outstanding write transactions to be continously accepted
    * with wready maintained high continuosly. wready is deasserted only on observing
    * a new transaction which will cross the threshold. Thus, setting this configuration
    * assumes that write data before address doesn't come once the threshold for maximum
    * outstanding transactions is reached and thus keeps wready asserted. 
    * Whereas disabling this configuration assumes that write data before address might 
    * come and thus deasserts wready when number of outstanding transactions
    * reach the threshold.
    * <b>type:</b> Dynamic
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand bit wdata_optimistic_flow_control_enable = 0;
`else
  rand bit wdata_optimistic_flow_control_enable = 1;
`endif

   /** 
    * @groupname axi3_4_config
    * Passive slave memory needs to be aware of the backdoor writes to memory.
    * Setting this configuration allows passive slave memory to be updated according to
    * RDATA seen in the transaction coming from the slave. Note that the passive slave 
    * memory is updated when all read data beats have been transmitted and accepted.
    * For an EXCLUSIVE transaction memory is updated only if all beats have an EXOKAY response.
    * For a normal transaction, memory is updated only if all beats have an OKAY response.
    * <b>type:</b> Static
    */
  rand bit memory_update_for_read_xact_enable = 0;

  /**
    * @groupname axi3_signal_width
    * Indicates if separate widths are required for ID  of write channel 
    * (AWID,WID and BID) and for ID of read channel(ARID and RID).
    * If set to 1, read_chan_id_width and write_chan_id_width are used
    * for setting the widths of the ID signals of corresponding channels.
    * If set to 0, id_width is used for setting the widths of all
    * ID signals.
    * This value must be consistent across all the ports in the system.
    *
    * Configuration type: Static
    */
  rand bit use_separate_rd_wr_chan_id_width = 0;

  /**
    * @groupname axi3_signal_width
    * If port is of kind MASTER:
    * This parameter defines the ID width of the master.
    * <br>
    * If port is of kind SLAVE:
    * This parameter defines the ID width of the slave. If an
    * interconnect is present, the ID width of the slave should
    * consider the maximum ID width of the masters in the system
    * and also consider additional bits required to represent
    * each master in the system.
    * <br>
    * Valid only when use_separate_rd_wr_chan_id_width is set to 0.
    *
    * Configuration type: Static
    */
  rand int id_width  = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of ARID and RID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int read_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname axi3_signal_width
    * Represents the width of AWID, WID and BID.  
    * Valid only when use_separate_rd_wr_chan_id_width is set to 1.
    * For slaves, the same considerations given for id_width are applicable.
    *
    * Configuration type: Static
    */
  rand int write_chan_id_width = `SVT_AXI_MAX_ID_WIDTH;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with barrier transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit barrier_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_min  = 0;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for barrier transactions.
    *
    * Configuration type: Static
    */
  rand int barrier_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines whether Normal transactions IDs can overlap with DVM transactions IDs.
    *
    * Configuration type: Static
    */
  rand bit dvm_id_overlap  = 1;

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the min ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_min  = ((1<<(`SVT_AXI_MAX_ID_WIDTH/2))-1);

  /**
    * @groupname ace_config
    * If port is of kind MASTER:
    * This parameter defines the max ID value of the master for dvm transactions.
    *
    * Configuration type: Static
    */
  rand int dvm_id_max  = ((1<<(`SVT_AXI_MAX_ID_WIDTH))-1);

  /**
   * Indicates how the information regarding the source master is 
   * transmitted to the slave
   * If set to STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is static and is defined by #source_master_id_xmit_to_slaves
   * If set to DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the source master information
   * is based on the value defined in svt_axi_transaction::dynamic_source_master_id_xmit_to_slaves
   * The value in dynamic_source_master_id_xmit_to_slaves must be populated by the user
   * in a system monitor callback issued at the start of the transaction.
   * If set to CUSTOM_SOURCE_MASTER_ID_XMIT_TO_SLAVES, the user must define 
   * svt_axi_system_configuration::is_master_id_and_slave_id_correlated to indicate
   * whether ID requirements for master and slave transactions are met 
   */
  source_master_id_xmit_to_slaves_type_enum source_master_id_xmit_to_slaves_type = STATIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES;
  
 /**
   * @groupname ace5_config 
   * Indicates whether data check parity feature is enable or not.
   * If set to ODD_PARITY_BYTE_DATA, then only on data check signals odd parity algorthim is used,
   * every 8bit of data is calculated and generated singles bit of datachk parity bit.
   * If set to ODD_PARITY_BYTE_ALL, then on both data check signals and control check signals odd parity algorthim is used.  
   * By default this enum is set to FALSE, which means data check fetaure is disabled.
   */ 
  check_type_enum check_type = FALSE;



  /**
    * @groupname axi_generic_config 
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If port is of kind MASTER:
    * This parameter defines the value that the interconnect assigns when
    * routing transactions to slave for all transactions originating from this
    * master. This value is specified in some bits of AxID of the transaction
    * that is routed to slave. This value must be based on the max value that
    * can be supported based on
    * svt_axi_system_configuration::source_master_info_id_width. For example, if the
    * interconnect uses 3 bits of AxID of the outgoing slave transaction to
    * specify the source master of the transaction,
    * svt_axi_system_configuration::source_master_info_id_width must be set to 3 and
    * this value must be less than 7. For more details, please refer
    * svt_axi_system_configuration::id_based_xact_correlation_enable
    */
  bit[`SVT_AXI_MAX_ID_WIDTH-1:0] source_master_id_xmit_to_slaves;

  /**
    * @groupname axi_generic_config
    * Applicable only when
    * svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * and axi_port_kind is MASTER
    * Indicates that the ID from this master is passed through without any
    * change when the interconnect routes it to the slaves. If this is set,
    * all transactions from this master are not appended with source master
    * information when routing to slaves
   */ 
  rand bit is_source_master_id_and_dest_slave_id_same = 0;

  /**
    * @groupname axi_generic_config 
    * Applicable only when svt_axi_system_configuration::id_based_xact_correlation_enable is set
    * If this parameter is set to zero, system monitor will not do id based correlation
    * for any transactions initiated/received at this specific port, this provides the option
    * for the user to avoid or select id based correlation for specific ports 
    * default value is 1.
    */
  bit id_based_xact_correlation_enable =1'b1;

  /** 
    * @groupname axi_generic_config
    * The byte boundary at which a master transaction is split to be
    * transmitted to two different slaves. This must be defined in cases where
    * pre_add_to_input_xact_queue callback in svt_axi_system_monitor_callback
    * is used to indicate that a master transaction is split and transmitted to
    * two different slaves. This parameter defines the boundary at which a
    * transaction is split
    *
    * Configuration type: Static
    */
  rand int byte_boundary_for_master_xact_split = `SVT_AXI_MAX_BYTE_BOUNDARY_FOR_MASTER_XACT_SPLIT;

  /**
   * @groupname ace_config
   * Enables support for WriteEvict transaction
   * Configuration type: Static
   */
  rand bit writeevict_enable = 0;

  /**
   * @groupname ace_config
   * Enables AWUNIQUE signal 
   * Configuration type: Static
   */
  rand bit awunique_enable = 0;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of outstanding transactions a master/slave
    * can support.
    * num_outstanding_xact = -1 is not supported for AXI4_STREAM
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY/AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * If #num_outstanding_xact = -1 then #num_outstanding_xact will not 
    * be considered , instead #num_read_outstanding_xact and 
    * #num_write_outstanding_xact have an effect.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_outstanding_xact = 4;

  /**
    * @groupname axi3_4_config
    * Specifies the number of READ outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert ARREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_read_outstanding_xact = 4;

  /** 
    * @groupname axi3_4_config
    * Specifies the number of WRITE outstanding transactions a master/slave
    * can support.
    * <br>
    * MASTER:
    * If the number of outstanding transactions is equal to this
    * number, the master will refrain from initiating any new 
    * transactions until the number of outstanding transactions
    * is less than this parameter.
    * <br>
    * SLAVE:
    * If the number of outstanding transactions is equal to 
    * this number, the slave will not assert AWREADY
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * <br>
    * This parameter will have an effect only if #num_outstanding_xact = -1.
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
  rand int num_write_outstanding_xact = 4;

  /** 
    * @groupname ace_config
    * Specifies the number of outstanding snoop transactions a master
    * can support. Applicable when axi_interface_type == AXI_ACE.
    * If the number of outstanding snoop transactions is equal to 
    * this number, the master will not assert ACREADY 
    * until the number of outstanding transactions becomes less
    * than this parameter. 
    * - <b>min val:</b> 1
    * - <b>max val:</b> Value defined by macro SVT_AXI_MAX_NUM_OUTSTANDING_SNOOP_XACT. Default value is 10.
    * - <b>type:</b> Static
    * .
    */ 
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int num_outstanding_snoop_xact = 4;
`else
  rand int num_outstanding_snoop_xact = 16;
`endif  

  /** 
    * @groupname axi_generic_config
    * 
    * Enables a separate port/export in the slave driver
    * (delayed_response_request_export) and sequencer
    * (delayed_response_request_port) through which the user can input response
    * data in a delayed manner.  When disabled all data and response
    * information related to a transaction must be given back to the driver
    * from the sequencer in the same timestamp as it receives a transaction
    * from the monitor.  When enabled, the user has flexibility to provide
    * response and data information at a later point in time through the
    * response port in the slave driver, although parameters related to the
    * delays to be applied for driving ARREADY, AWREADY and WREADY signals need
    * to be provided in the same timestamp. 
    * Refer to the user guide for a detailed description of the usage of this
    * parameter.
    */ 
  bit enable_delayed_response_port = 0;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of exclusive access transactions.
    * <br>
    * SLAVE:
    * Indicates whether the slave supports exclusive access or not.
    * <b>type:</b> Static
    *
    */
  rand bit exclusive_access_enable = 0;
  
  /** 
    * @groupname ace_config
    * MASTER:
    * This is applicable only when svt_axi_port_configuration::exclusive_access_enable is set to 1.
    * This bit controls enabling  Exclusive Monitor for AXI and ACE Masters.
    * If it is set to '1' then exclusive monitor is enabled in ace masters cache is updated on successful exclusive transactions based on coherent response and exclusive monitor state.
    * If this is set to '0' then exclusive monitor is disabled in ace master and for exclusive transaction cache
    * is updated only based on coherent response i.e. if it is received as EXOKAY.
    * <b>type:</b> Dynamic
    */
  rand bit exclusive_monitor_enable = 1;

  /** 
    * @groupname axi3_4_config
    * MASTER:
    * Enables generation of locked access transactions.
    * <b>type:</b> Static
    *
    */
  rand bit locked_access_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of barrier transactions.
    * <b>type:</b> Static
    */
  rand bit barrier_enable = 0;

  /** 
    * @groupname ace_config
    * MASTER:
    * Enables generation of DVM transactions.
    * <b>type:</b> Static
    */
  rand bit dvm_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only for active master 
    * Enables automated generation of DVMCOMPLETE transactions
    * in response to DVM Sync Snoop transactions. 
    * When this bit is unset, it is the user's responsibility to
    * send DVMCOMPLETE transactions from the sequence in response
    * to DVM Sync snoop transactions.
    * When this bit is set, the VIP master driver will auto generate 
    * DVMCOMPLETE transaction in response to DVM Sync snoop transactions.
    * When this bit is set, any DVMCOMPLETE transaction received from the sequencer will be ignored.
    */
  rand bit auto_gen_dvm_complete_enable = 0;

  /**
    * The minimum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int min_auto_gen_dvm_complete_delay = 0;

  /**
    * The maximum delay that needs to be applied to an auto-generated
    * DVM Complete transaction before it is processed by the driver.
    * The delay is applied from the point that the DVM Sync snoop
    * transaction corresponding to the DVM COMPLETE ends. 
    */
  rand int max_auto_gen_dvm_complete_delay = `SVT_AXI_MAX_DVM_COMPLETE_DELAY;

  /**
    * If this parameter is set, when a DVM snoop sync is received, the driver
    * takes a snapshot of active transactions whose address or data have been
    * sent on the interface.  The DVMCOMPLETE on the read address channel is
    * then launched when these outstanding transactions are complete. The
    * parameter #dvm_complete_delay is not applicable if this parameter is set. 
    */
  bit launch_auto_gen_dvm_complete_on_outstanding_xact_completion = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables speculative read.
    * A speculative read is defined as a read of a cache line that a master may
    * already be holding in its cache. Consider a case when user generates a
    * coherent transaction for read of a cache line that a master already holds
    * in its cache.
    *
    * When speculative read is enabled, the master will transmit this coherent
    * transaction. Also, the master will support cache state transitions as
    * defined in second set of tables in sections 5.5.1 to 5.5.11 in ACE
    * proposal 0.27.
    *
    * When speculative read is disabled, the master will not transmit this
    * coherent transaction. In this case, the master will only support cache
    * state transitions as defined in first set of tables in sections 5.5.1 to
    * 5.5.11 in ACE proposal 0.27.
    *
    * Whether a transaction is a speculative read is indicated by read-only
    * transaction class member svt_axi_transaction::is_speculative_read.
    *
    * <b>type:</b> Dynamic
    */
  rand bit speculative_read_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    *
    * MASTER:
    * Enables restrictions in the master for support of an external
    * snoop filter.
    * <b>type:</b> Dynamic
    */
  rand bit snoop_filter_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE_LITE.
    *
    * SLAVE:
    * Checks that cache maintenance transactions received by an interconnect
    * from a master are forwarded to corresponding slaves. This check will
    * be performed only if the system monitor is enabled and correlation of
    * master and slave transactions are enabled by setting 
    * id_based_correlation_enable in svt_axi_system_configuration and the associated
    * configuration properties. 
    * <b>type:</b> Dynamic
    */
  rand bit forward_cmos_to_slaves_check_enable = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE or ACE_LITE.
    * MASTER:
    * Determines the permissible cache line state transitions in the master.
    * For each transaction type, the section 5 of the specification provides 
    * cache line state transitions for "expected (or recommended) end state", 
    * "legal end state with snoop filter" and "legal end state without snoop filter".  
    * This parameter determines which of the above state changes are to be
    * used.
    *
    * Below are the supported values:
    * - RECOMMENDED_CACHE_LINE_STATE_CHANGE: The cache line state
    * changes as given in the "expected end state" of each table is used.
    * - LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state with snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 1. The actual cache line state change can be done using
    * member svt_axi_transaction::force_to_shared_state.
    * - LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE: The cache 
    * line state changes as given in the "legal end state without snoop filter" 
    * of each table is used. To be able to use this cache line state transition,
    * the configuration member svt_axi_port_configuration::snoop_filter_enable
    * must be set to 0. The actual cache line state change can be done using
    * members svt_axi_transaction::force_to_invalid_state and
    * svt_axi_transaction::force_to_shared_state.
    * .
    *
    * <b>type:</b> Dynamic
    */
  rand axi_cache_line_state_change_type_enum cache_line_state_change_type = RECOMMENDED_CACHE_LINE_STATE_CHANGE;

  /**
   * @groupname ace_config
   * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component.
   *
   * Specifies how master will process incoming snoop request when memory update transaction is in progress.
   * if it is set to SUSPEND_SNOOP_DURING_MEM_UPDATE then master will suspend incoming snoop request and will respond
   * after current memory update transaction is complete. This is the default response mode.
   * If it is set to RESPOND_SNOOP_DURING_MEM_UPDATE then master will not suspend incoming snoop request. Instead it will
   * respond to the incoming snoop request as allowed by ACE specification.
   * If it is set to EITHER_RESPOND_OR_SUSPEND_SNOOP_DURING_MEM_UPDATE then master will randomly decide to choose between
   * either of the above two behaviour i.e. either suspend incoming snoop or respond to it.
   * 
   * Configuration type: Dynamic
   */
  rand snoop_response_mode_during_mem_update_type_enum snoop_response_mode_during_mem_update = SUSPEND_SNOOP_DURING_MEM_UPDATE;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to ACE and it is Master component
    *
    * Indicates how dirty data in cache should be transferred on receiving a snoop.
    * As per section C5.2.2 of the AXI specification, a cached master can ensure that data in a dirty cacheline
    * is available to a snoop other than MAKEINVALID in one of two ways:
    * 1. returning data when the master completes the snoop
    * 2. carrying out a memory update, using a WRITEBACK or WRITECLEAN before responding to the snoop
    * This configuration indicates which of the above two methods will be used for returning data
    * Note that if there is an outstanding WRITEUNIQUE or WRITELINEUNIQUE transaction in the
    * queue of the master, then data will be returned with the snoop transaction. This is to comply with
    * restrictions on WRITEUNIQUE and WRITELINEUNIQUE while a snoop is in progress as per section
    * C4.8.7 of the spec
    */
  rand snoop_response_data_transfer_mode_enum snoop_response_data_transfer_mode = SNOOP_RESP_DATA_TRANSFER_USING_CDDATA;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE and it is Master component
    *
    * Describes various address randomization mode for nonshareable transaction with domain type SYSTEMSHAREABLE. It indicates what
    * address range should or shouldn't be used while randomizing axi master transaction based on the different enum values listed below.
    *
    * NONSHAREABLE_XACT_FULL_ADDRESS_SPACE :: allows full address sapce to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE :: allows only address sapce outside inner, outer or nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_WITHIN_NON_SHAREABLE_ADDR_RANGE :: allows only nonshareable address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_ADDR_RANGE :: allows only address sapce outside inner or outer address range to be used for nonshareable transaciton with domain type SYSTEMSHAREABLE 
    * default value :: NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE
    */
  rand nonshareable_xact_address_range_in_systemshareable_mode_enum nonshareable_xact_address_range_in_systemshareable_mode = NONSHAREABLE_XACT_ADDR_OUTSIDE_INNER_OUTER_NON_SHAREABLE_ADDR_RANGE;

  /**
    * @groupname axi3_4_config
    * MASTER:
    * The maximum number of active exclusive transactions that will be initiated by the master.
    * SLAVE:
    * The maximum number of active exclusive access monitors supported by the slave. Attempts to
    * exceed this max number results in a failed exclusive access read response of OKAY instead of EXOKAY.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS
    * NOTE: if it is set to '0' value then there are no restrictions on maximum number of active exclusive
    * transactions. VIP will not mark any exclusive sequence as failed because of this parameter.
    * <b>type:</b> Static
    */ 
  rand int max_num_exclusive_access   = `SVT_AXI_MAX_NUM_EXCLUSIVE_ACCESS;
      
  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Number of ADDRESS bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    *
    * It can also be configured with ( -1 ) to indicate that address ranges for 
    * each exclusive monitor is defined through user specified start and end address ranges.
    * For this, user should configure start_address_ranges_for_exclusive_monitor[] and
    * end_address_ranges_for_exclusive_monitor[] arrays in system configuration.
    * A svt_axi_system_configuration::set_exclusive_monitor_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,
    *     bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr) utility method can be used for this purpose.
    *
    * NOTE: configuring with value 0 means, no address is being monitored by the 
    * corresponding exclusive monitor and hence exclusive access to different address
    * may also affect current thread.
    *
    * <b>specail value:</b> -1 indicates that num_addr_bits_used_in_exclusive_monitor and
    * num_initial_addr_bits_ignored_by_exclusive_monitor are not used. Instead address
    * ranges for exclusive monitors are defined by address_ranges_for_exclusive_monitor[] array.
    *
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ADDR_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_addr_bits_used_in_exclusive_monitor   = `SVT_AXI_MAX_ADDR_WIDTH;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * ACE Exclusive monitor will ignore number of initial address bits as
    * indicated by this configuration member.
    * Example: A coherent interconnect can divide its whole address space into
    *          multiple ranges such that each PoS Exclusive monitor checks only
    * its corresponding address range. So, if it allocates 1/2 GB address space to each
    * of the 4 PoS exclusive monitors then num_initial_addr_bits_ignored_by_exclusive_monitor
    * needs to be configured as 29 (1.5GB - 2GB ~ 31 bits).
    */
  rand int num_initial_addr_bits_ignored_by_exclusive_monitor   = 0;

  /**
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type
    * is ACE
    * INTERCONNECT:
    * Number of ID bits that need to be monitored by the exclusive monitors for 
    * current port in order to support one or more independent exclusive access
    * thread.
    * NOTE: configuring with value 0 means, no id is being monitored by the 
    * corresponding exclusive monitor and hence only single exclusive access thread
    * is supported for current port.
    *  <b> This feature is not supported yet </b>
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_ID_WIDTH-1
    * <b>type:</b> Static
    */ 
  rand int num_id_bits_used_in_exclusive_monitor     = `SVT_AXI_MAX_ID_WIDTH;

   /*
    * @groupname ace_config
    * Applicable only when svt_axi_port_configuration::axi_interface_type is ACE
    * INTERCONNECT:
    * Indicates whether Interconnect uses seperate PoS Exclusive Monitor for 
    * secured or non-secured exclusive access.
    * NOTE: configuring with value 0 means, interconnect doesn't monitor seperately
    * for secured or unsecured exclusive access.
    * <b> This feature is supported by enabling secure address space by configuring tagged_address_space_attributes_enable = 1 </b>
    * <b> User shouldn't use this configuration parameter, it is going to be deprecated </b> 0
    * <b>min val:</b> 0
    * <b>max val:</b> 1
    * <b>type:</b> Static
    */ 
  rand bit use_secured_exclusive_monitor             = 1;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will not assert error if Master sends Exclusive Store without sending Exlusive Load.
    * However, if Exclusive Store is sent from the Invalid cacheline state then VIP will still assert error since,
    * that is not a valid state to start Exclusive Store.
    * <b>type:</b> Static
    */ 
  rand bit allow_exclusive_store_without_exclusive_load = 0;

  /**
    * @groupname ace_config
    * If set to '1' then VIP will respond to very first Exclusive Store with EXOKAY response. This means that if
    * no master has performed any exclusive transaction after reset is de-asserted then the master that issues
    * exclusive store will be responded with EXOKAY or VIP will expect EXOKAY response from the coherent interconnect.
    * Note: reference point of first exclusive store is reset.
    * <b>type:</b> Static
    */ 
  rand bit allow_first_exclusive_store_to_succeed = 0;

  /**
    * @groupname ace_config
    * If set to '1' then Exclusive Monitor will get reset once Exclusive Store is successful.
    * If set to '0' then Exclusive Monitor will remain set even if Exclusive Store is successful.
    * Please Note that, VIP will still reset Exclusive Monitor for failed Exclusive Store attempt
    * regardless of the value set for this parameter.
    * <b>type:</b> Static
    */ 
  rand bit reset_exclusive_monitor_on_successful_exclusive_store = 1;

  /**
    * @groupname ace_config
    * This control register indicates different modes of error conditions uded in exclusive monitor.
    * [0] => If set to '1' implies that Snoop Error will cause an exclusive sequence to fail only if
    *        either data_transfer bit or pass_dirty bit is set to '1'. Otherwise, if snoop response
    *        indicates error bit as asserted then regardless of data_transfer bit or pass_dirty bit
    *        values exclusive sequence will fail. 
    * [31:1] => Reserved bits.
    * Default Value :: 0x00000000
    */
  rand bit[31:0] exclusive_monitor_error_control_reg = 0;

  /** 
    * @groupname ace_config
    * If shareable exclusive access needs to be supported from ace-lite port then this parameter
    * should be set to '1'. If it is set to '1' then VIP will allow READONCE or WRITEUNIQUE
    * transactions to be of exclusive type.
    * Default Value: '0' i.e. shareable exclusive access from ace-lite port is not allowed. Only
    *                non-shareable exclusive transactions as READNOSNOOP or WRITENOSNOOP are allowed.
    */
  rand bit shareable_exclusive_access_from_acelite_ports_enable = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of write transactions that can be interleaved
    * This parameter should not be greater than #num_outstanding_xact.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted write data beyond this value.
    * SLAVE: 
    * Checks that received write data is not interleaved beyond this value. 
    * An error is issued if write data is interleaved 
    * beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int write_data_interleave_depth       = `SVT_AXI_MAX_WR_INTERLEAVE_DEPTH;

  /** 
    * @groupname axi3_4_config
    * This parameter specifies the atomicity size required to check the address
    * alignment for a given transcation as per the atomicity of component.<br>
    * This parameter will not have effect if set to -1. The values specified
    * to this parameter should be power of 2, in terms of Bytes <br>
    * Default value: -1.<br>
    * Allowed values: should be power of 2, in terms of Bytes. <br>
    * For example: 8, 16, 32, 64 etc <br>
    * <b>type:</b> Static
    *
    */
  rand int atomicity_size = -1;


  /** @cond PRIVATE */
  /**
    * When set to 1, enables id reflection in AXI4_LITE mode.
    * This enables the awid, bid and rid signals. This allows
    * an AXI4-Lite slave to be used on a full AXI interface,
    * without a bridge function, in a system that guarantees that
    * the slave can only be accessed by transactions that fall
    * within the AXI4-Lite subset.
    * <b>type:</b> Static
    *
    * This parameter is not yet supported.
    */
  rand bit id_reflection_enable = 0;
  /** @endcond */

  /**
    * @groupname axi3_4_config
    * Applicable only to MASTER when axi_interface_type is 
    * AXI3/AXI4/AXI4_LITE.
    * When set to 1, accesses to the read address channel and 
    * write address channel are serialized. Thus, awvalid and
    * arvalid will never be asserted at the same time. The
    * address information driven on the write address channel
    * will have to be accepted before any address information
    * on the read address channel is driven and viceversa. 
    * When set to 0, activity on the read address channel and
    * write address channel occur in parallel.
    */
  rand bit serial_read_write_access = 0;

`ifndef SVT_EXCLUDE_VCAP
  /**
    * @groupname axi_traffic_profile 
    * Enables use of traffic profiles. This enables the use of transaction
    * generation at a higher level of abstraction.  This feature
    * is only available as part of the NOC product. Please refer to the NOC
    * user guide for details
    */
  bit use_traffic_profile = 0;

  /** 
    * @groupname axi_generic_config
    * Enables FIFO based rate control. 
    * A FIFO is modelled in the driver for read and write
    * transactions separately. A WRITE transaction can be sent
    * out if there is sufficient data in the FIFO to send out that
    * transaction. A READ transaction can be sent out if there is
    * space in the FIFO to receive the data of the READ transaction.
    * The current level of a WRITE FIFO is incremented every clock
    * based on write_fifo_fill_rate.With every data beat, the currentl level
    * is decremented based on burst_size of the transaction. The current level of a READ FIFO
    * is decremented every clock based on read_fifo_drain_rate. With every data
    * beat, the current level is incremented based on burst_size of the transaction.
    * A WRITE transaction will be sent out if the current level is greater than
    * the total number of bytes of all outstanding write transactions + the total
    * number of bytes of the current transaction. A READ transaction will be sent out
    * if the current level is less than the difference of the read_fifo_full_level and
    * the total number of bytes of all outstanding read transactions + the total number
    * of bytes of the current transaction.
    */
  rand bit use_fifo_based_rate_control = 0;

  /**
    * @groupname axi_generic_config
    * Clock period in ns. This is used to calculate the drain/fill rate in
    * bytes/cycle
    */
  real clock_period = 1;

  /** 
    * @groupname axi_generic_config
    * The drain rate in MBPS of the FIFO into which data from READ
    * transactions is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction
    */
  rand int read_fifo_drain_rate = `SVT_AXI_MAX_READ_FIFO_DRAIN_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the READ FIFO into which data from READ transactions
    * is dumped. Used by the check_current_fill_level_read_fifo 
    * method of the corresponding driver to determine if there is space
    * in the FIFO to receive data of a READ transaction.
    */
  rand int read_fifo_full_level = `SVT_AXI_MAX_READ_FIFO_FULL_LEVEL;

  /** 
    * @groupname axi_generic_config
    * The fill rate in MBPS of the FIFO from which data for WRITE 
    * transactions is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to send a WRITE transaction
    */
  rand int write_fifo_fill_rate = `SVT_AXI_MAX_WRITE_FIFO_FILL_RATE;

  /** 
    * @groupname axi_generic_config
    * The full level in bytes of the WRITE FIFO from which data for WRITE transactions
    * is taken. Used by the check_current_fill_level_write_fifo 
    * method of the corresponding driver to determine if there is enough 
    * data in the FIFO to transmit data of a WRITE transaction
    */
  rand int write_fifo_full_level = `SVT_AXI_MAX_WRITE_FIFO_FULL_LEVEL;

  /**
    * @groupname axi_generic_config
    * Determines if the READ FIFO is empty on start up
    */
  rand bit is_read_fifo_empty_on_start = 1;

  /**
    * @groupname axi_generic_config
    * Determines if the WRITE FIFO is empty on start up
    */
  rand bit is_write_fifo_empty_on_start = 1;
`endif //SVT_EXCLUDE_VCAP

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, AXI transaction phase level information is
    * printed in note verbosity.  Messages related to start & end of address,
    * data and response phases are printed.  If unset, AXI transaction phase
    * level information is printed only in debug verbosity.
    */ 
  bit display_xact_phase_messages = 0;

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding transactions
    * per AxID is limited to 1 for Non-Device and Non-DVM transactions.
    * This can be further controlled by configuration
    * svt_axi_port_configuration::single_outstanding_per_id_kind. 
    */ 
  bit single_outstanding_per_id_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set, maximum number of outstanding AXI4_STREAM transactions
    * per TDEST is limited to 1.
    */ 
  bit single_outstanding_per_tdest_enable = 0; 

  /** 
    * @groupname axi_generic_config
    * If this parameter is set to 1, all delay related parameters will be set
    * to 0. Note however, that actual delay on interface will vary based on
    * outstanding transactions.
    */ 
  rand bit zero_delay_enable = 0; 
  
  /**
    * This enumerated type controls the AxID when
    * svt_axi_port_configuration::single_outstanding_per_id_enable is set to 1.
    *
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * 'MODIFY_SAME_ID': If AxID of a new Non Device or Non DVM transaction matches
    * AxID of an active transaction, the VIP modifies the AxID such that the AxID 
    * is not overlapping with AxID of any active Non Device or Non DVM transactions.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated
    * by the user sequence. At this time, another Non Device or Non DVM with AxID = 6
    * is already in progress. In this case, VIP will check the active queue, and modify
    * the AxID of the new transaction to an un-used AxID. For example, VIP will modify 
    * the AxID of new transaction to 4, if this is not used by any active transactions.
    * 
    * If svt_axi_port_configuration::single_outstanding_per_id_kind is set to
    * ‘WAIT_FOR_COMPLETION_OF_SAME_ID': If AxID of a new Non Device or Non DVM transaction
    * matches AxID of an active Non Device or Non DVM transaction, the VIP waits till the
    * corresponding active Non Device or Non DVM transaction is complete. Only when the
    * active Non Device or Non DVM transaction is complete, VIP adds the new Non Device
    * or Non DVM transaction to the active queue. This ensures that only 1 active Non Device
    * or Non DVM transaction exists for a given AxID.
    *
    * For example, a new Non Device or Non DVM transaction with AxID = 6 is initiated by
    * the user sequence. At this time, another Non Device or Non DVM with AxID = 6 is already
    * in progress. In this case, VIP will wait for the active transaction to complete. After
    * active transaction is complete, VIP will add the new transaction with AxID = 6 to the
    * active queue.
    */
  typedef enum {
    MODIFY_SAME_ID = 0,
    WAIT_FOR_COMPLETION_OF_SAME_ID = 1
  } single_outstanding_per_id_kind_enum;

  single_outstanding_per_id_kind_enum single_outstanding_per_id_kind = WAIT_FOR_COMPLETION_OF_SAME_ID;

  /**
    * If this parameter is set, debug information is driven on the debug ports.
    * The transaction id as well as the transfer id corresponding to 
    * each beat is driven on the debug ports.
    *
    * 
    *
    * <b>type:</b> Static
    */
  bit use_debug_interface = 0; 



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checking. In a disabled state, no protocol
    * violation messages (error or warning) are issued.
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol check statistics collection. In a disabled state, statistics 
    * on checks executed are not collected. Enabling this has a run-time performance impact
    * <b>type:</b> Dynamic 
    */
  bit protocol_check_stats_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables toggle coverage.
    * Toggle Coverage gives us information on whether a bit
    * toggled from 0 to 1 and back from 1 to 0. This does not
    * indicate that every value of a multi-bit vector was seen, but
    * measures if individual bits of a multi-bit vector toggled.
    * This coverage gives information on whether a system is connected
    * properly or not.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit toggle_coverage_enable = 1;
  `else
  bit toggle_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables state coverage of signals.
    * State Coverage covers all possible states of a signal.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit state_coverage_enable = 1;
  `else
  bit state_coverage_enable = 0;
  `endif


  /** @cond PRIVATE */
  /**
    * Enables meta coverage of signals.
    * This covers second-order coverage data such as valid-ready
    * delays.
    * <br>
    * This parameter is not supported currently. The meta coverage is enabled
    * using port configuration parameter #transaction_coverage_enable.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit meta_coverage_enable = 1;
  `else
  bit meta_coverage_enable = 0;
  `endif

  /** @endcond */

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables transaction level coverage. This parameter also enables delay
    * coverage. Delay coverage is coverage on various delays between valid & ready signals.
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit transaction_coverage_enable = 1;
  `else
  bit transaction_coverage_enable = 0;
  `endif
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables protocol checks coverage. 
    * <b>type:</b> Static 
    */
  `ifdef SVT_AMBA_DEFAULT_COV_ENABLE
  bit protocol_checks_coverage_enable = 1;
  `else
  bit protocol_checks_coverage_enable = 0;
  `endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables positive or negative protocol checks coverage. 
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables signal valid check during reset when protocol_checks_enable=1. 
    * When set to '1', enables signal valid check during reset.
    * When set to '0', disables signal valid check during reset. In a disabled
    * state, no signal valid check during reset violation messages (error or warning) are issued.
    * <b>type:</b> Static 
    */
  bit signal_valid_during_reset_checks_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid. 
    * <b>type:</b> Static 
    */
  int cov_same_id_in_outstanding_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Set of multiple ID values used for matching outstanding read/write transactions for
    * covergroups trans_axi_num_outstanding_xacts_with_multiple_same_arid and 
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid. 
    * <b>type:</b> Static 
    */
  int cov_multi_same_ids[];

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching back to back write transactions for
    * covergroups trans_master_ace_lite_coherent_and_ace_snoop_response_association_with_specific_id. 
    * <b>type:</b> Static 
    */
  int cov_specific_id_in_back_to_back_xacts = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables valid_ready_dependency_coverage 
    * <b>type:</b> Static 
    */
  // When valid_ready_dependency_coverage_enable is set to '1' for IUS simulator
  // the function cov_sample_``dependency () of svt_axi_port_monitor_def_cov_util.svi
  // consumes around 10x more time. So because of this, the default value is kept 0 for the IUS simulator.
  // valid_ready_dependency covergroups as performance intensive and hence diabling them by default.
`ifndef INCA
  bit valid_ready_dependency_coverage_enable= 0;
`else 
  bit valid_ready_dependency_coverage_enable= 0;
`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wvalid deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rready deassertion for covergroup signal_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which arready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_arready_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * arready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_arready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid  need to be deasserted after
    * wready deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wvalid need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wvalid_bvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_wready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * awready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_awready_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * wready deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_wready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * rvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_rvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bready need to be deasserted after
    * bvalid deassertion for covergroup signal_master_slave_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bready_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_awvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */ 
  int cov_num_clks_awready_and_wvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * rvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_rvalid_dependency = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which awready need to be deasserted after
    * bvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_awready_and_bvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * awvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_awvalid_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * wvalid deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_wvalid_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which wready need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_wready_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which rvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_rvalid_and_bready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * awready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_awready_dependency = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * wready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_wready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * rready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_rready_dependency  = 10;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Number of clock cycles for which bvalid need to be deasserted after
    * bready deassertion for covergroup signal_slave_master_valid_ready_dependency. 
    * <b>type:</b> Static 
    */
  int cov_num_clks_bvalid_and_bready_dependency  = 10;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroups
    * trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_write_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins each for 
    * covergroups trans_axi_num_outstanding_xacts_with_same_awid and 
    * trans_axi_num_outstanding_xacts_with_same_awid
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_snoop_xacts.It should be programmed to 
    * a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_snoop_xact which
    * indicates the number of outstanding snoop transactions VIP can support.
    *
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_snoop_xact
    * <b>type:</b> Static 
    */
  int cov_bins_num_outstanding_snoop_xacts = 64;

  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates the number of bins which will be created for covergroup
    * trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid.
    * It should be programmed to a value less than or equal to configured value of 
    * svt_axi_port_configuration::num_outstanding_xact or 
    * svt_axi_port_configuration::num_read_outstanding_xact if 
    * svt_axi_port_configuration::num_outstanding_xact is set to -1 which
    * indicates the number of outstanding transactions VIP can support.
    * If user does not program this variable it will create 64 bins for 
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid 
    * <b>type:</b> Static 
    */
  int cov_bins_dvm_tlbi_num_outstanding_xacts = 64;  

  /**
    * @groupname axi_coverage_protocol_checks
    * ID value used for matching outstanding DVM TLBI transactions for
    * covergroup trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid. 
    * <b>type:</b> Static    
    */
  int cov_same_id_in_dvm_tlbi_outstanding_xacts = 0;  
  /**
    * @groupname axi_coverage_protocol_checks
    * Indicates if user wants to cover all the id_ranges of the outstanding
    * transactions. BY default , Only fixed number of outstanding transactions will be covered 
    * <b>type:</b> Static 
    */
  bit cov_num_outstanding_xacts_range_enable = 0;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awaddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and bresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and araddr signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and rresp signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_rresp_enable = 1;
    /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,rresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_rresp_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic_type,bresp signal.
    * <b>type:</b> Dynamic 
    */
  bit trans_cross_axi_atomictype_bresp_enable = 1;



  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arprot signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen, awaddr and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awaddr_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst,
    * awlen and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awlock_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst, awlen
    * and awcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awlen_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst,
    * arlen, araddr and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_araddr_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arlock signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arlock_enable = 1;

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type,atomic_xact_op_type,awsize
    * and awburst signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_comp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , atomic xact op type , awburst
    * and awsize signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_atomic_noncomp_awburst_awsize_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , bresp and
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_bresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type ,bresp
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_bresp_burst_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type , rresp 
    * and awlen signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_rresp_burst_length_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic compare transaction type
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_comp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between atomic non compare transaction type 
    * and endianness.
    * <b>type:</b> Static 
    */
 bit trans_cross_atomic_noncomp_endianness_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write transaction type , awmmussid and
    * and awmmusecsid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmusecsid_awmmussid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between write_xact_type , awmmussidv and awmmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_write_xact_type_awmmussidv_awmmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type,armmusecsid and armmusid signal.
    * <b>type:</b> Static 
    */
bit trans_cross_read_xact_type_armmusecsid_armmusid_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between read_xact_type , armmussidv
    * and armmussid signal.
    * <b>type:</b> Static 
    */
 bit trans_cross_read_xact_type_armmussidv_armmussid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_nid
    * and stash_nid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_nid_stashnid_valid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between coherent stash transaction type , stash_lpid
    * and stash_lpid_valid.
    * <b>type:</b> Static 
    */
bit trans_cross_stash_xact_type_stash_lpid_stashlpid_valid_enable = 1;

`endif

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst, arlen
    * and arcache signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arlen_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between awburst and
    * awqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_awburst_awqos_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for cross coverage between arburst and 
    * arqos signal.
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_arburst_arqos_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * bresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop, awdomain 
    * and bresp signal.
    * The EXOKAY response is permitted for WriteNoSnoop for NONSHAREABLE and SYSTEMSHAREABLE domains. 
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awsnoop_awdomain_bresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awdomain and awcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awdomain_awcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop and 
    * awbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_awbar_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * awdomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_awdomain_awbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (MEMORY_BARRIER and SYNC_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_memory_sync_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arbarrier (NORMAL_ACCESS_RESPECT_BARRIER and NORMAL_ACCESS_IGNORE_BARRIER) and 
    * ardomain signal.
    * <b>type:</b> Dynamic 
    */
  bit  trans_cross_ace_ardomain_arbarrier_respect_ignore_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks    
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arburst signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arburst_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arlen signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arlen_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arsize signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arsize_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * araddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arcache_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_coh_rresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * ardomain and arcache signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_ardomain_arcache_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop and 
    * arbar signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_arbar_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between ardvmmessage and 
    * ardvmresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_ardvmmessage_ardvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acaddr signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * acprot signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_acprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop and 
    * ace rresp signal.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_crresp_enable = 1; 

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acdvmmessages
    * and acdvmresp.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acdvmmessage_acdvmresp_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between arsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_arsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between awsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_awsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables ACE transaction level coverage group for cross coverage between acsnoop
    * initial cache line status and final cache line status.
    * <b>type:</b> Static 
    */
  bit  trans_cross_ace_acsnoop_cacheinitialstate_cachefinalstate_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_read_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level meta coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi_write_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level meta coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_meta_axi4_stream_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI4 STREAM transaction level delay coverage group for axi4 stream transfer
    * <b>type:</b> Static 
    */
  bit trans_axi4_stream_delay_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_read_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level out-of-order response coverage group for write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_ooo_write_response_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI STREAM transaction level coverage group for cross coverage
    * between stream transaction type, tid and tdest.
    * <b>type:</b> Static 
    */
  bit trans_cross_stream_xact_type_tid_tdest_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for axi outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_outstanding_xact_enable = 1;
  
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_outstanding_xact coverage group for
    * axi barrier outstanding transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_outstanding_xact_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_barrier_pair_sequence coverage group for
    * read and write barrier pair transaction
    * <b>type:</b> Static 
    */
  bit trans_ace_barrier_pair_sequence_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables AXI transaction level trans_non_barrier_xact_after_256_outstanding_barrier_xact coverage group
    * <b>type:</b> Static 
    */
  bit trans_non_barrier_xact_after_256_outstanding_barrier_xact_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_read_burst_sequence coverage group for
    * back to back read pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_read_burst_sequence_enable = 1;

 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_back_to_back_write_burst_sequence coverage group for
    * back to back write pair transaction
    * <b>type:</b> Static 
    */
  bit trans_axi_back_to_back_write_burst_sequence_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_same_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with same ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_same_id_completed_out_of_order_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_write_read_diff_id_completed_out_of_order coverage group for
    * WRITE/READ transactions with diff ID completed OOO
    * <b>type:</b> Static 
    */
  bit trans_axi_write_read_diff_id_completed_out_of_order_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width48 ,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width40,trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_tlbinvl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_tlbinvl_modes_virtaddr_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width48  ,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width40,trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_branch_predictor_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_branch_predictor_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for  trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width32,
    * trans_cross_ace_dvm_phy_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_phy_inst_cache_invl_modes_modes_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width48,
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width40,trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width32
    * trans_cross_ace_dvm_virt_inst_cache_invl_modes_virtaddr_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_virt_inst_cache_invl_modes_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_addr_range_width48,
    * trans_cross_ace_dvm_firstpart_addr_range_width40,trans_cross_ace_dvm_firstpart_addr_range_width32,
    * trans_cross_ace_dvm_firstpart_addr_range_width24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_addr_range_cov_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction  coverage group for trans_cross_ace_dvm_firstpart_secondpart_addr_range_width65,
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range56,trans_cross_ace_dvm_firstpart_secondpart_addr_range32
    * trans_cross_ace_dvm_firstpart_secondpart_addr_range24 depending on cfg.addr_width
    * <b>type:</b> Static 
    */
  bit trans_cross_ace_dvm_firstpart_secondpart_addr_range_cov_enable = 1;
  
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_state_RD_WR_burst_sequence coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_four_state_rd_wr_burst_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_four_excl_normal_sequence coverage group
    * This cover group covers specific combinations of exclusive and normal transactions
    * <b>type:</b> Static 
    */

  bit trans_axi_four_excl_normal_sequence_cov_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_lock_followed_by_excl_sequence coverage group
    * <b>type:</b> Static 
    */
  bit trans_lock_followed_by_excl_sequence_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_fixed_burst_wstrb coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_fixed_burst_wstrb_cov_enable = 1; 
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer coverage group 
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_awcache_modifiable_bit_write_unaligned_transfer_cov_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_arcache_modifiable_bit_read_unaligned_transfer_cov_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level axi_wstrb_to_signal_unaligned_start_address coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_wstrb_to_signal_unaligned_start_address_cov_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_same_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_same_arid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_read_outstanding_xact_diff_arid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_cache_modifiable_bit_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_read_outstanding_xact_diff_arid_device_cacheable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_same_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_same_awid_cache_modifiable_bit_enable = 1;
   
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_write_outstanding_xact_diff_awid_cache_modifiable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_cache_modifiable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_write_outstanding_xact_diff_awid_device_cacheable_bit_enable = 1;
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_multiple_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level
    * trans_axi_num_outstanding_xacts_with_multiple_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_multiple_same_awid_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_enable = 1;
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_arid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_same_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_same_awid_enable = 1;

 
   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_enable = 1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_axi_num_outstanding_xacts_with_diff_awid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_axi_num_outstanding_xacts_with_diff_awid_range_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_snoop_xacts coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_snoop_xacts_enable = 1;

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_same_arid_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_enable = 1;  
/**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range coverage group
    * <b>type:</b> Static 
    */

  bit trans_ace_num_outstanding_dvm_tlb_invalidate_xacts_with_diff_arid_range_enable = 1;  

   /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_arcache coverage group
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_atomictype_exclusive_arcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_axi_atomictype_exclusive_awcache  coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_axi_atomictype_exclusive_awcache_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awsnoop_awdomain_awprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_writeunique_awdomain_awprot_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables cross coverage of  transaction parameters with slave port_id for
    * the following covergroups.
    * - trans_cross_ace_awsnoop_awsize
    * - trans_cross_ace_arsnoop_arsize
    * - trans_cross_ace_awsnoop_awlen
    * - trans_cross_ace_arsnoop_arlen
    * - trans_cross_ace_awsnoop_awdomain
    * - trans_cross_ace_arsnoop_ardomain
    * - trans_cross_ace_awsnoop_awcache
    * - trans_cross_ace_arsnoop_arcache
    * - trans_cross_ace_awsnoop_awburst
    * - trans_cross_ace_arsnoop_arburst
    * - trans_cross_ace_awsnoop_bresp
    * - trans_cross_ace_arsnoop_coh_rresp
    * Basically, it covers if the transaction properties have been covered from the master to all the different slaves
    * .
    * <b>type:</b> Static 
    */
  bit cov_trans_cross_slave_port_id_enable = 0;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arsnoop_ardomain_arprot coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_readonce_ardomain_arprot_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_awprot_awbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_awprot_awbarrier_memory_sync_enable = 1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level trans_cross_ace_arprot_arbarrier_memory_sync coverage group
    * <b>type:</b> Static 
    */

  bit trans_cross_ace_arprot_arbarrier_memory_sync_enable = 1;
      
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write strobes 
    * <b>type:</b> Static 
    */  
  bit trans_cross_axi_write_strobes_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read interleaving depth
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_interleaving_depth_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for write narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_narrow_transfer_awlen_awaddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for read narror transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_narrow_transfer_arlen_araddr_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned write transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_write_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group for unaligned read transfer
    * <b>type:</b> Static 
    */
  bit trans_cross_axi_read_unaligned_transfer_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction coverage group for master_to_slave_path_access
    * <b>type:</b> Static 
    */
  bit trans_cross_master_to_slave_path_access_cov_enable = 0;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_enable = 1;  

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_coherent_and_ace_snoop_response_association
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_coherent_and_ace_snoop_response_association_enable = 1;  
 
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_specific_id_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id
    * covergroup
    * <b>type:</b> Static 
    */
  bit trans_master_ace_lite_coherent_and_ace_snoop_response_association_back_to_back_xact_with_specific_id_enable = 1;

  /** @cond PRIVATE */
   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, for non monifiable transaction cache_type 
    * and prot_type fields are compared.
    * By default this configuration parameter is set to 1 to enable cache_type and prot_type comparation,
    * if this parameter is set 0 then cache_type and prot_type comparations are dissabled
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  bit master_slave_xact_association_cache_prot_check_enable = 1;
  /** @endcond */

   /**
    * @groupname master_slave_xact_association
    * In Master Slave transaction association flow, cache_type[3:1] and prot_type fields are compared.
    * By default this configuration parameter is set to SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK
    * to enable cache_type and prot_type comparation for non modifiable transaction,
    * if this parameter is set SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_MODIFIABLE_NONMODIFIABLE_CACHE_TYPE_CHECK
    * it enables cache_type and prot_type comparation for modifiable and non modifiable transactions,
    * in master slave transaction association.
    * Note that to enable or dissable this feature, you also need to enable AXI
    * System Monitor using member #system_monitor_enable.
    * <b>type:</b> Static
    */ 
  master_slave_xact_association_cache_prot_check_enum master_slave_xact_association_cache_prot_check = SVT_AXI_MASTER_SLAVE_XACT_ASSOCIATION_NONMODIFIABLE_CHECK;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for snoop transfer
    * <b>type:</b> Static 
    */
  bit trans_axi_snoop_enable = 1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_read_with_same_id_to_different_slaves_enable = 1;
  
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_arsnoop_acsnoop 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_arsnoop_acsnoop_enable =1;
  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_enabled 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_writeevict_disabled
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_overlapping_awsnoop_acsnoop_crresp_enable =1;
 /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp 
    * <b>type:</b> Static 
    */
  bit trans_ace_concurrent_non_overlapping_awsnoop_acsnoop_crresp_enable =1;

  /**
    * @groupname axi_coverage_protocol_checks
    * Enables AXI transaction level coverage group 
    * svt_axi_port_monitor_def_cov_callback::trans_outstanding_read_with_same_id_to_different_slaves
    * <b>type:</b> Static 
    */
  bit trans_outstanding_write_with_same_id_to_different_slaves_enable = 1;
  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transactions on
    * AR, AW channel waiting for snoop response
    * <b>type:</b> Static 
    */
  bit trans_ar_aw_stalled_for_ac_channel_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after nonshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_nonshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after innershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_innershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after outershareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_outershareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction domain
    * after systemshareable barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_domain_after_systemshareable_barrier_enable = 1;

  /**
    * @groupname ace_coverage_protocol_checks
    * Enables ACE transaction level coverage group for transaction ordering
    * after barrier
    * <b>type:</b> Static 
    */
  bit trans_xact_ordering_after_barrier_enable = 1;

  /**
    * Determines if the transaction trace file generation is enabled.
    * 
    * - 1'b1 : Enable trace file generation. 
    * - 1'b0 : Disable trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_tracing = 1'b0;

   /**
    * Determines if transaction reporting is enabled.
    * 
    * - 1'b1 : Enable transaction reporting.
    * - 1'b0 : Disable transaction reporting. 
    * .
    * 
    * <b>type:</b> Static
    */
   bit enable_reporting = 1'b0;

  /**
    * Applicable only when enable_tracing or enable_reporting is set.
    * Determines if transaction data should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data in trace file generation. 
    * - 1'b0 : Disable data in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_trace_enable = 1'b0;
  
  /**
    * Applicable only when enable_tracing or enable_reporting and data_trace_enable is set.
    * Determines if transaction data_beat should be included as part of trace file
    * generation/reporting. Takes effect only if the product of 'data width in
    * bytes' and 'max burst length in AXI3 (16)' is less than or equal to 1024.
    * This restriction is imposed to avoid an overlow of characters
    * 
    * - 1'b1 : Enable data_beat in trace file generation. 
    * - 1'b0 : Disable data_beat in trace file generation.
    * .
    * 
    * <b>type:</b> Static
    */
   bit data_beat_trace_enable = 1'b0;

  /** 
    * @groupname protocol_analyzer
    * Determines if XML generation is enabled.
    * <b>type:</b> Static
    */
  bit enable_xml_gen = 0;

  /**
   * @groupname protocol_analyzer
   * Indicates whether XML generation is included for memcore operations. The resulting
   * file can be loaded in Protocol Analyzer to obtain a graphical presenation of the
   * memcore activity. Set the value to 1 to enable the memcore XML generation.
   * Set the value to 0 to disable the memcore XML generation.
   * 
   * <b>type:</b> Static
   */
  bit enable_memcore_xml_gen = 0;
 
  /**
   * Determines in which format the file should write the transaction data.
   * The enum value svt_xml_writer::XML indicates XML format, 
   * svt_xml_writer::FSDB indicates FSDB format and 
   * svt_xml_writer::BOTH indicates both XML and FSDB formats.
   */
  svt_xml_writer::format_type_enum pa_format_type ;
  
  
  // **********************************************
  // Configuration parameters for STREAM interface
  // **********************************************
  /** @cond PRIVATE */
  /** 
    * Signifies the presense of the TREADY signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tready_enable               = 1;

  /** 
    * Signifies the presense of the TKEEP signal in the VIP. 
    * <b>type:</b> Static
    * Not yet supported.
    */
  rand bit tkeep_enable                = 1;

  /** @endcond */

  /** 
    * Signifies the presense of the TSTRB signal in the VIP. 
    * <b>type:</b> Static
    * Value of tstrb is consider as 0 when tstrb_enable = 0.
    */
  rand bit tstrb_enable                = 1;

  /** 
    * Signifies the presense of the TID signal in the VIP. 
    * <b>type:</b> Static
    * Value of tid is consider as 0 when tid_enable = 0.
    */
  rand bit tid_enable                  = 1;

  /** 
    * Signifies the presense of the TDEST signal in the VIP. 
    * <b>type:</b> Static
    * Value of tdest is consider as 0 when tdest_enable = 0.
    */
  rand bit tdest_enable                = 1;

  /** 
    * Signifies the presense of the TUSER signal in the VIP. 
    * <b>type:</b> Static
    * Value of tuser is consider as 0 when tuser_enable = 0.
    */
  rand bit tuser_enable                = 1;

  /** 
    * Signifies the presense of the TDATA signal in the VIP. 
    * <b>type:</b> Static
    * Value of data is consider as 0 when tdata_enable = 0. If TDATA is not present it is required that TSTRB is not present
    */
  rand bit tdata_enable                = 1;

  /** 
    * Signifies the presense of the TLAST signal in the VIP. 
    * <b>type:</b> Static
    * All transfers are considered as individual packets when tlast_enable = 0.
    */
  rand bit tlast_enable                = 1;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDATA signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tdata_width                 = `SVT_AXI_MAX_TDATA_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    * <b>type:</b> Static
    */
  rand int tid_width                   = `SVT_AXI_MAX_TID_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TDEST signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tdest_width                 = `SVT_AXI_MAX_TDEST_WIDTH;

  /** 
    * @groupname axi4_stream_signal_width
    * Width of TUSER signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM. 
    * <b>type:</b> Static
    */
  rand int tuser_width                 = `SVT_AXI_MAX_TUSER_WIDTH;

  /** @cond PRIVATE */
  /** Setting this parameter to 1, enables the generation of a
    * byte stream type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit byte_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_aligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * continuous un-aligned type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit continuous_unaligned_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of a
    * a sparse type of data stream. 
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit sparse_stream_enable = 1;

  /** Setting this parameter to 1, enables the generation of user defined 
    * streams.
    * Applicable only when svt_axi_port_configuration::axi_interface_type 
    * is AXI4_STREAM. 
    * <b>type:</b> Static 
    */
  rand bit user_stream_enable = 1;
  /** @endcond */

  /**
    * Specifies the number of stream transactions that can be interleaved.
    * When set to 1, interleaving is not allowed.
    * MASTER: 
    * Does not interleave transmitted streams beyond this value.
    * SLAVE: 
    * Checks that received streams are not interleaved beyond this value. 
    * An error is issued if streams are interleaved beyond this value.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WR_INTERLEAVE_DEPTH
    * <b>type:</b> Static
    */ 
  rand int stream_interleave_depth       = `SVT_AXI_MAX_STREAM_INTERLEAVE_DEPTH;

  // **********************************************
  // End of Configuration parameters for STREAM interface
  // **********************************************

  /** 
    * @groupname default_ready
    * Default value of AWREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_awready = 1;

  /** 
    * @groupname default_ready
    * Default value of WREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_wready = 1; 

  /** 
    * @groupname default_ready
    * Default value of ARREADY signal. 
    * <b>type:</b> Dynamic
    */
  rand bit default_arready = 1;

   /** 
    * @groupname default_ready
    * Default value of RREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_rready = 1;

  /** 
    * @groupname default_ready
    * Default value of BREADY signal. 
    * <b>type:</b> Dynamic 
    */
  rand bit default_bready = 1;

  /**
    * @groupname default_ready
    * Default value of ACREADY signal.
    * Applicable when axi_interface_type is ACE.
    * <b>type:</b> Dynamic 
    */
  rand bit default_acready = 1;

  /**
    * @groupname default_ready
    * Default value of CRREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_crready = 1;  
 
  /**
    * @groupname default_ready
    * Default value of CDREADY signal.
    * Applicable when axi_interface_type is ACE.
    * Applicable only to SLAVE 
    * <b>type:</b> Dynamic 
    */
  rand bit default_cdready = 1;

  /**
    * @groupname default_ready
    * Default value of TREADY signal.
    * Applicable when axi_interface_type is AXI4_STREAM.
    * <b>type:</b> Dynamic 
    */
  rand bit default_tready = 0;

  /** 
    * @groupname default_ready
    * Default value of QVN VxREADY signal. 
    * <b>type:</b> Dynamic
    */
  `ifdef SVT_AXI_QVN_ENABLE
  rand bit default_qvn_ready = 1;
  `endif

  /** 
    * @groupname axi_signal_inactive_wdata_byte_value
    * When the VALID signal of the write data channel is high and wstrb is low, all
    * inactive wdata byte lane will take this value and valid wdata remains in the 
    * active byte lane.
    * <b>type:</b> Dynamic 
    */
  rand wdata_val_enum inactive_wdata_bytes_val = INACTIVE_WDATA_BYTE_UNCHANGED_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_addr_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic 
    */
  rand idle_val_enum write_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read address channel is low, all other
    * signals (except the READY signal) in that channel will take this value.
    * <b>type:</b> Dynamic 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_PREV_VAL;
`else
  rand idle_val_enum read_addr_chan_idle_val =INACTIVE_CHAN_X_VAL ;
`endif
  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the read data channel is low, all other signals 
    * (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum read_data_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * When the VALID signal of the write response channel is low, all other 
    * signals (except the READY signal) in that channel will take this value. 
    * <b>type:</b> Dynamic
    */
  rand idle_val_enum write_resp_chan_idle_val = INACTIVE_CHAN_PREV_VAL;

  /** 
    * @groupname axi_signal_idle_value
    * Enables toggling of ready signals when corresponding valid is low
    * The exact manner in which the ready signals are toggled depends on
    * the values set in svt_axi_transaction::idle_addr_ready_delay,
    * svt_axi_transaction::idle_wready_delay, svt_axi_transaction::idle_rready_delay
    * and svt_axi_transaction::idle_bready_delay
    * <b>type:</b> Static 
    */
  rand bit toggle_ready_signals_during_idle_period = 0;
 
  /** @cond PRIVATE */
  /** If this parameter is set, the master checks for any outstanding 
    * transaction with an overlapping address before sending a transaction.
    * If there is any such outstanding transaction, the master will wait
    * for it to complete before sending a transaction.
    * <b>type:</b> Static 
    *
    * This parameter is not yet supported.
    */
  rand bit addr_overlap_check_enable = 0;
  /** @endcond */

  /** 
    * @groupname axi3_4_config
    * The number of addresses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a read ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
`ifndef SVT_AMBA_ALTERNATE_DEFAULT_VALUE
  rand int read_data_reordering_depth = 1;
`else
  rand int read_data_reordering_depth = 16;
`endif

   /** 
    * @groupname axi3_4_config
    * The number of responses pending in the slave that can be 
    * reordered. A slave that processes all transactions in  
    * order has a write resp ordering depth of one.
    * This parameter’s max value is defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. 
    * The default value of this macro is 8, and is user configurable. 
    * Refer section 3.3.7 of AXI user manual for more info on System Constants.
    * <b>min val:</b> 1
    * <b>max val:</b> \`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH (Value defined by macro SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH. Default value is 8.)
    * <b>type:</b> Static 
    */
  rand int write_resp_reordering_depth = 1;

  /**
    * @groupname axi3_4_config
    * Specifies the number of beats of read data that must stay 
    * together before it can be interleaved with read data from a
    * different transaction.
    * When set to 0, interleaving is not allowed.
    * When set to 1, there is no restriction on interleaving.
    * <b>min val:</b> 0
    * <b>max val:</b> \`SVT_AXI_MAX_READ_DATA_INTERLEAVE_SIZE 
    * <b>type:</b> Static 
    */
  rand int read_data_interleave_size = 0;

  /**
   * @groupname axi3_4_config
   * Specifies how the reordering depth of transactions moves.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_window_enum reordering_window = MOVING;
      
  /**
   * @groupname axi3_4_config
   * Specifies the reordering algorithm used for reordering the 
   * transactions or responses.
   * 
   * Applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
   */
  rand reordering_algorithm_enum reordering_algorithm = ROUND_ROBIN;
  
  /** 
    * @groupname axi3_4_config
    * This parameter is added to control the reordering priority, in which svt_axi_transaction::reordering_priority 
    * value Vs reordering priority scheme.
    *
    * This member is applicable only when svt_axi_port_configuration::reordering_algorithm
    * is svt_axi_port_configuration::PRIORITIZED.
    *
    * If this bit is set to ‘1’ then transactions with svt_axi_transaction::reordering_priority highest value 
    * for this attribute will get higher priority.
    *
    * If this bit is set to ‘0’ then transactions with svt_axi_transaction::reordering_priority least value 
    * for this attribute will get higher priority.
    *
    * Default value of this bit is set to ‘0’.
    *
    * Applicable for ACTIVE SLAVE only.
    *
    * Configuration type: Static
    */
  rand bit reordering_priority_high_value = 0;

  /** 
    * @groupname axi3_4_config
    * The AXI3 protocol requires that the write response for write 
    * transactions must not be given until the clock cycle 
    * after the acceptance of the last data transfer.
    * In addition, the AXI4 protocol requires that the write response for
    * write transactions must not be given until the clock
    * cycle after address acceptance. Setting this
    * parameter to 1, enforces this second condition in AXI3
    * based systems as well. It is illegal to set this parameter to 0
    * in an AXI4 based system.
    * <b>type:</b> Static 
    */
  rand bit write_resp_wait_for_addr_accept = 1;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address to be received before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID is received.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr = 0;

  /**
    * @groupname axi3_4_config
    * Applicable only to active slave vip.
    * Waits for address handshake to be completed before driving wready.
    * Applicable to a transaction where data arrives before address.  In such a
    * scenario, if this parameter is set, wready is asserted only after the
    * corresponding AWVALID-AWREADY handshake is completed.
    * Applicable only when svt_axi_port_configuration::default_wready=0.
    */
  rand bit wready_wait_for_awaddr_handshake = 0;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This parameter is added to enable the structural dependency feature.
    * User has to set this bit to 1'b1 to enable the structural dependency feature.
    */
  
  rand bit axi_slv_channel_buffers_enable  = 0;
 
  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write data buffer.
    * The default value is set to 4096.
    * This default value considers that the AMBA AXI supports maximum burst_length of 256. Since the default value of axi_wr_addr_buffer is 16, a value of 256*16 is reasonable 
   */
  
  rand integer axi_wr_data_buffer = 4096;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Write response buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_wr_resp_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read address buffer.
    * The default value is set to 16.
    */
  
  rand integer axi_rd_addr_buffer = 16;

  /**
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * This variable configures the depth of Read response buffer.
    * The default value is set to 4096.
    */
  
  rand integer axi_rd_resp_buffer = 4096;

  /** 
    * @groupname axi3_4_config
    * Applicalbe only to slave.
    * Number of FIFO memories to be configured for this port.
    * Each FIFO memory has a specifc address and is given in
    * #fifo_mem_addresses. Needs to be used in conjunction with
    * svt_axi_slave_memory_sequence for UVM/OVM. For VMM, #generator_type must
    * be set to MEMORY_RESPONSE_GEN. If there is a FIXED type burst access
    * to one of these addresses, then data is written/read in the corresponding
    * FIFO. If there is a FIXED type burst access to an address that is not
    * configured in fifo_mem_addresses, a SLVERR response is issued.  If there
    * is a FIFO underrun when a READ is issued, a SLVERR is given as response
    * <b>type:</b> Static 
    */
  int num_fifo_mem = 0;

  /**
    * @groupname axi3_4_config
    * Addresses corresponding to each FIFO
    * The size of this array should be equal to #num_fifo_mem
    * <b>type:</b> Static 
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] fifo_mem_addresses[];
  
  /** @cond PRIVATE */
  /**
    * The AXI slave currently supports two types of memory:
    * 1. A legacy SV based memory. This is the solution by default. For more information refer to the class reference documentation of svt_mem.
    * 2. A C based memory which has more features compared to the SV based memory. For more information refer to the class reference documentation of svt_mem_core. 
    * If the memory type is set to this, the following needs to be done:
    * a. Pass/include (as elaboration options to vcs/mti/nc) “${DESIGNWARE_HOME}/vip/svt/common/latest/C/lib/${platform}/libmemserver.so"
    * b. Set LD_LIBRARY_PATH as $DESIGNWARE_HOME/vip/svt/common/latest/C/lib/$platform (or prescript file if using dw_home build)
    */
  mem_type_enum mem_type = SV_BASED_SVT_MEM;
  /** @endcond */

  /** @cond PRIVATE */
  /** 
    * Enables the internal memory of the slave.
    * Write data is written into the internal memory and read
    * data is driven based on the contents of the memory.
    *
    * <b>type:</b> Static
    *
    * This parameter is not yet supported. The slave supports built-in memory,
    * but this parameter is not currently required to enable the memory.
    */
  bit enable_mem = 1;
  /** @endcond */

  /**
    * Enables address generation based on the values configured
    * in {nonshareable_start_addr,nonshareable_end_addr},
    * {innershareable_start_addr,innershareable_start_addr} and
    * {outershareable_start_addr,outershareable_end_addr} which are set
    * through svt_axi_system_configuration::create_new_domain() and
    * svt_axi_system_configuration::set_addr_for_domain().
    * This establishes a relationship between the addresses (svt_axi_transaction::addr)
    * and domain_types(svt_axi_transaction::domain_type) generated in a transaction.
    */
  bit enable_domain_based_addr_gen = 0;

  /**
    * An array of start addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_end_addr to form an address range applicable
    * to a nonshareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_start_addr[];

  /**
    * An array of end addresses corresponding to the nonshareable
    * region of memory. Each member pairs with a corresponding
    * member of nonshareable_start_addr to form an address range applicable
    * to a nonshareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] nonshareable_end_addr[];

  /**
    * An array of start addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_end_addr to form an address range applicable
    * to a innershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the innershareable
    * region of memory. Each member pairs with a corresponding
    * member of innershareable_start_addr to form an address range applicable
    * to a innershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] innershareable_end_addr[];

  /**
    * An array of start addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_end_addr to form an address range applicable
    * to a outershareable region. 
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_start_addr[];

  /**
    * An array of end addresses corresponding to the outershareable
    * region of memory. Each member pairs with a corresponding
    * member of outershareable_start_addr to form an address range applicable
    * to a outershareable region.
    * This variable is not to be set directly by the user. It is set
    * internally by the model, when domain information is set using
    * svt_axi_system_configuration::set_addr_for_domain()
    * Applicable when interface_type is svt_axi_port_configuration::AXI_ACE
    * or svt_axi_port_configuration::ACE_LITE
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] outershareable_end_addr[];

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the protection type (as indicated by
   * svt_axi_transaction::prot_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the protection type properties recorded in the cache are set
   * for the auto-generated transaction
    */
  bit update_cache_for_prot_type = 0;

  /** Applicable only when axi_interface_type is set to AXI_ACE.  Indicates if
   * the cache must be updated with the memory attributes(as indicated by
   * svt_axi_transaction::cache_type) of the transaction that makes an entry in
   * the cache. If the VIP auto-generates a transaction for evicting an entry
   * from cache or for cleaning a cacheline before sending a cache maintenance
   * transaction, the memory attributes recorded in the cache are set for the
   * auto-generated transaction
    */
  bit update_cache_for_memory_attributes = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * the cache must be updated for WRITENOSNOOP and READNOSNOOP transactions.
    * Currently supported only if  cache_line_state_change_type is set to
    * RECOMMENDED_CACHE_LINE_STATE_CHANGE. Cache is updated only if
    * transactions are a full cacheline access. Transactions with sparse write
    * strobes are also allowed. If transactions with partial or multiple
    * cacheline accesses are received by the master driver, existing entries in
    * the cache for the corresponding address(s) will be deleted. If this bit
    * is set and svt_axi_transaction::force_xact_to_cache_line_size is set, a
    * constraint in the master transaction forces all WRITENOSNOOP and
    * READNOSNOOP to be of a full cacheline access and FIXED types bursts are
    * not allowed. The specification allows a cacheline to move from the
    * invalid state to a valid state only for a full cacheline access.
    * Therefore any backdoor access to the cache to write into non-shareable
    * region must write into all bytes of the cacheline. For a WRITENOSNOOP
    * transaction, if the cacheline is dirty and a transaction with partial
    * write strobes is received, the VIP merges dirty data from the cache and
    * the data in the transaction and transmits it. If the cacheline is clean,
    * no merging of data is performed. If the cacheline does not exist,
    * allocations are not made for a WRITENOSNOOP transaction based on section
    * C4.8.1 and Table C4-20 of the specification, since there are no cacheline
    * state transitions from an invalid state to a valid state. Hence, a
    * WRITENOSNOOP will modify cache contents only if the cache is already
    * allocated either through a READNOSNOOP or through backdoor access of
    * cache. For a READNOSNOOP transaction, if there is no entry in the cache,
    * a new cacheline is allocated only if
    * svt_axi_transaction::allocate_in_cache is set. If there is already an
    * entry in the cache, the status of the cache is updated, but the data is
    * not because this indicates a speculative read and the data in cache may
    * be the latest copy.  Cacheline state transitions for READNOSNOOP
    * transactions correspond to section C4.5.1 of the specification. 
    */
  bit update_cache_for_non_coherent_xacts = 0;

  /**
    * Applicable only when axi_interface_type is set to AXI_ACE. Indicates if
    * data must always be supplied for READONCE, READCLEAN, READSHARED,
    * READNOTSHAREDDIRTY and READUNIQUE snoop transactions on the snoop data
    * channel if the cacheline is in a valid state. If this value is set to 0, data may or may not be transferred based on randomization
    */
  bit transfer_snoop_data_always_if_valid_cacheline = 1;

    /** 
    * @groupname axi3_4_config
    * If this bit is set to ‘1’ then transactions are only eligible for "write_resp_chan_lock" only after 
    * both address phase and data phase are completed.
    *
    * If this bit is set to ‘0’ then transactions  are eligible for “write_resp_chan_lock” after
    * Address phase is completed.In here "data phase" is not considered. 
    * 
    * Default value is ‘0’.
    * This attribute is applicable only to the READ data and WRITE resp transactions processed by ACTIVE Slave.
    *
    * ** Note, Eligible transaction are given the “write_resp_chan_lock” according to the “reordering algorithm”.
    */
  bit write_resp_wait_for_data_accept = 0;

  /** @cond PRIVATE */
`ifdef SVT_VMM_TECHNOLOGY
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals spcified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * <b>type:</b> Dynamic
    */
`else
  /**
    * @groupname axi_performance_analysis 
    * The interval based on which performance parameters are monitored and
    * reported. The simulation time is divided into time intervals specified by this
    * parameter and performance parameters are monitored and reported based on
    * these. Typically, this interval affects measurement of performance
    * parameters that require aggregation of values across several transactions
    * such as the average latency for a transaction to complete. The unit for
    * this parameter is the same as the simulation time unit.
    * When set to 0, the total simulation time is not divided into time intervals.
    * For example, consider that this parameter is set to 1000 and that the
    * simulation time unit is 1ns. Then, all performance metrics that require
    * aggregation will be measured separately for each 1000 ns. Also, min and max
    * performance parameters will be reported separately for each time interval.
    * If this parameter is changed dynamically, the new value will take effect
    * only after the current time interval elapses.
    * <br>
    * When set to -1, svt_axi_port_perf_status::start_performance_monitoring() and
    * svt_axi_port_perf_status::stop_performance_monitoring() needs to be used to
    * indicate the start and stop events for the performance monitoring. If the
    * start and stop events are not indicated, the performance monitoring will not 
    * be enabled. If the stop event is not indicated after issuing a start event,
    * the port monitor stops the performance monitoring in the extract phase.
    * Note that any constraint checks will be performed only during the monitoring period.
    * <b>type:</b> Dynamic
    */
`endif  
  real perf_recording_interval = 0;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a write
    * transaction to complete. The duration is measured as the time when the
    * the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    */
  real perf_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a write transaction to
    * complete. The duration is measured as the time when the the transaction
    * is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a write
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_write_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed duration for a read
    * transaction to complete. The duration is measured as the time when the the
    * transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum duration for a read transaction to
    * complete. The duration is measured as the time when the the transaction is
    * started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is more than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_max_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected average duration for a read
    * transaction. The average is calculated over a time interval specified by
    * perf_recording_interval. A violation is reported if the computed average
    * duration is less than this parameter. The duration is measured as the time
    * when the the transaction is started to the time when transaction ends.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_avg_min_read_xact_latency = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for read
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected throughput for write
    * transfers in a given time interval. The throughput is measured as 
    * (number of bytes transferred in an interval)/(duration of interval).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a throughput
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_throughput = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for read
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_read_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the maximum allowed bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_max_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis 
    * Performance constraint on the minimum expected bandwidth for write
    * transfers in a given time interval. The bandwidth is measured as 
    * (number of bytes transferred in an interval)/(latency).
    * The interval is specified in perf_recording_interval.
    * The unit for this is Bytes/Timescale Unit. For example, if a bandwidth
    * of 100 MB/s is to be configured and the timescale is 1ns/1ps, it translates
    * to (100 * 10^6) bytes per 10^9 ns and so this needs to be configured to 0.1.
    * A value of -1 indicates that no performance monitoring is done.
    * <b>type:</b> Dynamic 
    * When #perf_recording_interval is set to -1, check related to this constraint is
    * performed only while the performance monitoring is active.
    */
  real perf_min_write_bandwidth = -1;

  /**
    * @groupname axi_performance_analysis
    * Indicates if periods of transaction inactivity (ie, periods when no
    * transaction is active) must be excluded from the calculation of
    * throughput.  The throughput is measured as (number of bytes transferred
    * in an interval)/(duration of interval). If this bit is set, inactive
    * periods will be deducted from the duration of the interval
    */
  bit perf_exclude_inactive_periods_for_throughput = 0;
  
  /**
    * @groupname axi_performance_analysis
    * Indicates how the transaction inactivity (ie, periods when no
    * transaction is active) must be estimated for the calculation of
    * throughput.  
    * Applicable only when svt_axi_port_configuration::
    * perf_exclude_inactive_periods_for_throughput is set to 1. 
    * EXCLUDE_ALL: Excludes all the inactivity. This is the default value. 
    * EXCLUDE_BEGIN_END: Excludes the inactivity only from time 0 to start of first 
    * transaction, and from end of last transaction to end of simulation. 
    */
  perf_inactivity_algorithm_type_enum perf_inactivity_algorithm_type = EXCLUDE_ALL;
  /** @endcond */

`ifdef SVT_ACE5_ENABLE
   /**
     * @groupname ace5_config
     *  It can be set to either of three values below:
     *  mte_support_type =svt_axi_port_configuration:STANDARD.
     *  When set to the above value memory tagging is supported on the interface, all tag operation types are supported
     *	mte_support_type = svt_axi_port_configuration:BASIC.
     *  When set to the above value memory tagging is supported on the interface at a basic level, a limited range of tag operations are supported. 
     *	mte_support_type = svt_axi_port_configuration:FALSE.
     *  When set to NOT_SUPPORTED , memory tagging is not supported on the interface
     *  Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
     */
  mte_support_type_enum mte_support_type = NOT_SUPPORTED;

 /**
   * @groupname ace5_config
   * Bcomp signal
   * Only applicable when SVT_ACE5_ENABLE macro is defined and svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0
   */
  bit bcomp_signal_enable; 
`endif

`ifdef SVT_ACE5_ENABLE
 /**
    * @groupname ace5_config
    * Enables unique id identifier feature for write and read address and response channels
    * <b>type:</b> Static
    * Only applicable when SVT_ACE5_ENABLE macro is defined and 
    * svt_axi_port_configuration::ace_version is set to ACE_VERSION_2_0 or higher
    *
    * This functionality is not supported yet.
    */
   bit unique_id_enable  = 0; 

 /**
   * @groupname ace5_config
   * Enables Read Data Chunking feature support in master and slave. 
   * <b>type:</b> Static
   * Only applicable when SVT_ACE5_ENABLE macro is defined. 
   * Not yet implemented.
   */
  bit rdata_chunking_enable = 0;

   /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunknum signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunknum_width                   = `SVT_AXI_MAX_CHUNK_NUM_WIDTH;

  /** 
    * @groupname ace5_config 
    * It is used to set width of the rchunkstrb signal. Applicable when
    * <b>type:</b> Static
    * Not yet implemented.
    */
  rand int rchunkstrb_width                   = `SVT_AXI_MAX_CHUNK_STROBE_WIDTH;
`endif

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /*   pre_randomize does the following
   *   1) Calculates number of tagged address attributes set to '1'
   */
  extern function void pre_randomize ();

`protected
HZEgE5dd4PGd0Z@QKLeF<XG_@5Hf>9)PPQfH<NdF728;La3]<Tc]1)BNH2fJ:PU(
\d(MIgKKbZM:=fN/-WK[1?32Hcd9U8E.^)JH^)8N3<)NgQ(16KY]-0D?L+O1\MJC
#I3H7g/H2X&^V\>BN;17GVYO7@(L5JAM;$
`endprotected


`ifdef SVT_ACE5_ENABLE
/** 
 * Returns 1 if bcomp response is applicable on this port else returns 0
 */
 extern function bit is_bcomp_response_valid();   
`endif

`ifdef SVT_VMM_TECHNOLOGY
/** @cond PRIVATE */
  /** 
    * @groupname axi_generic_config
    * The source for the stimulus that is connected to the transactor.
    * This member is not used.
    * Configuration type: Static
    */
  generator_type_enum snoop_generator_type = SCENARIO_GEN;
/** @endcond */
`endif

//vcs_vip_protect
`protected
Jf8eP:(:L/\F6J@A.gJJYJ?=H9deCGD>Z,N<9N5)bM8b,0?POXYX3(Q6,BPX5c2/
Ca\FCVRZG<W,b+1/LA+aDU[R@L/7RB.TEW_,04KF+45;AC(U.7)RS\UF(c6b5KRD
=eO&>/#Q?T(ac/5#e]5JC8Z15B3P[b>^IF8)3eec\SY5O;5bB?FSANfE3MAJ3fg;
0+Pe,D0b<_7AS[133H0Zf-X,,8-7\<)C(91\ACT6:U1f8GTQb@1^&_Ug;03/e\gd
&a]&B<Vb2C]9NdLJ5U7H^L/VP;/4U0Z@E0<J(X\9b2:f@2G1f5;JS8B[R-G8.(<C
(d7_?GaRR[]D.9D\1-(2JCb/fJSa]L=@.^;GbS]26ITJa[_XNZ>aK]Y9M+C2E,c5
+S8)b[H#5&-4X1PbJ9D2W<>QJ#T+N9AaCbNG+]5cZ^OUVW1&-CgPS#/]AF+T.NC)
A4J:A,AE0K6XBA463T\?S&1PO.OA2-G:dZ5(c25N3fE,[A@S(>@&#)M54.A9G/.P
CAS1S.4C,=A8=NB72If&[-NA^WJ))[+J?YIH?WB.KXP86+@+c-\]cHF+c]=DGS?D
g9aa<,M71.:4P>)?a>8K+>=F06ccL)@bTW_>>e:g@JS]I5/=BAdZ?,VX1@Ndd-X,
M:FV16dGM:X#3QJcTS0:FVcEaQd(>W^REOTP11174NNR<,R<:g)C9FA>(A&e<&G(
/ae)Z@#>>O0]C@J^c4^e@g_(+?/:,2g9[H,KE5I\U8cW]=Db_(G;\C(LH9Pd93Y.
]K6F5PK47R7J^Z#<aCW]0/TaLLa6JKg?E2b,U&)U:cR[[KBXfH^.XRHEOeNWD9C]
+)Z37<SI^;C<CUWPJBB5R]1:#8/9T5A&X.[D-A[F@-UZ4Q<>+.RKO4:5&Q@[aIKS
<PPM#EDdLeZB&9S^LP=;;1</B\0d,-P=>G/cV7-4d.d2DF^GbDUU:,V.UG]J?(KL
^?=A>5U+,H/;BQI:97K\MX,faQ=DW)^C6ef2Rg.C6)d\GGK\&d.93<cdePM]4gU8
.99ed#O8bCJS=YI<eFB5f5+,;#;IRa7/QBVQ5W9-1K+6QMBA@[9?4P2Q2=<KJ,57
X96LW<C9Z[I3fg:cE5]dV]3B+X8ZI9>D.RA:^^W_[W;+--M4[?6]VV@AJO(:HEYG
WDS+411ZDEcR-Xb2N\d?NS,3X_C3-]M.Wc90-,R\cMIGX1f4V\0gL.2@4NFFK+Q-
X&0IUPC[OW_PSa-bZ3Hb<CYb?[:LG+ZKDCDVKLH)JY,,CZD&3:1dF3(=cPN\2#35
e/>F-?[_V(,:+-O#G&YccPT6C4VPT^J[+[)Bf?PK7SFa[f))K,[^(N(]:dR30FA<
)2-G_TWV7G+bE6(CaeMF>,e=URX7S,#=A6U#Pge^@IfLdBVB#;K9e2cac_8RCP:K
^G3+L/DZ/Vd&A\)0S-3./S)bID[VW&cU^E?Oc0;J9L]bYUF=K4,<)H]2@/YSZ+fP
K]33KT+<eDO&QB</@Tf7H);+(7@eQd:\(=AI]>6UF+E_V,XXQM23HD+?O=8VH?F=
.TE(>>[=-Zc5J@ETU:2R9Ue/8+N-;AWE))O>4X722-I>+GE:F6SF#+dI3C10)[6F
XEb<]d1[b-=M0PQ>8e@_\9/4GQY:HQgYB,W#3c5YJPW<\YDR&1>K<R5QNLfRI7XC
0#-F@N@0TV]EeZ^8(\F&OJI>M9HBTP7e0JJ]8.dX1J6F5ZY\S0H_[MI5WOU,BX##
d63e@SGA_YU8HCaA;e3eG.0-a[TS\e2(BCJ^cUXFEMEC7W[=22.ZK@2GeJ)H]TGJ
<L3PH[]d#HBS_NW2CCT2X^>aG=MKDMIXR0A^/f_HS\N(CI-7JWE8J&OAUU,S7RQ;
.cOK_\KdL<G(G@NQ+]],/Q;ZEU/TXAG_Q9=;X7+@-4f,K92Sb3V&2H+MFd27OWNb
Y#E\Y]<#GE=f,0f\CKH4OEF:A-GC9c]SQZ<R(#:J]HJBK_Q\@;3e-7XRZ)3X,1.J
UCZS7RUW\AR5XBJ0+WG;5b_NL::JL+e4HFe=Z6-5O7+YHK<I5gZ?bIL[T[\XYDNO
Ld>4a<6aXg>;8,R4>73\T=0YRFePQDcE]9YW:g9R_--_XeJ[6Z2Z3/DKfeLcMIB:
\N^+NB#1OHPdR]d@b2Z+gF@.LJ+<ZLV[MMS[V4gRDb28O_f^)HJ?@c#FL0=cCHAN
+A61LR)M)BUfE+FE?=U/eUg@+B6H.;PYR9<;=AfO8&Q2JNAaUSQ\I1-/-M7e<aK[
^/ZEKfUUf<OM@LGT@@(JV[LEP0/X:NfQ.UA5WE^I;1b5N6,Y>@G5QWO6;;]+E-bI
-:BU8[DH=(gFRf85Af1&NQ9g][gZ=NXI_5?_TL@V@NFOGa\H6OA)\>S.=efDg5E(
f\5<cH=c(_e5N0PH;]M2JHcG62IZ.f3O^3KKQR>/5;15^^X/FVgb@G=?cTD_Jg(]
fcUQMRaH6d@I#/DJ_Q-^TbPUNFEJF8Y0fRN1&)LNJ/6fK83J9DfbEQ]]eB)62KS;
_[?a,c]?L9:,2J(Y804YA9I5WX+@@1ST3-(I^,geRfZJ?d^\EJK&G9SL6gX;RC\P
)[RE#1YJ&RGN[8S@O6VCb.4XG3CA^Z0=1b@]63;7)B\5aG==S9M(BA;fX]\7&.<E
&2@B[aEe^&[,[fgB4\b>X&F7O5<]>VK7@/.fbJW]BXL>3[)Lc,^L9+#N5T#N#&O^
XdU^eX0\T1a#V)0YG4([94M)FWf:NWGU8DN1gYSV5H0@8eJA_T]LJDK1V@-b8;GH
]>VEM\EJWP)D6\L<-<7?4A^-P<G7RS0H)#0=1DM:LP_NVVP(EAF4H\TYEC15(I48
1-_G_^gQLF<Uf)(D9=U&N0ZPY,Ra:ML?[2FN_+(VY.TTHH&6Q=Y092-7EJR(O9EU
3L4170H.V.B=JWRRSP-#Ycb]H@,ZR9JEOR;]ZS6?9WZO5IT8Tc:V-)OCSeZ85fZZ
S3@?7b#?I>WX,89IC>1aLVS.?K=dUTGNBA6RAN)-&PaXC-^EI(US;gZD;:ETR&Tc
O-,5M&KZJJgGG=d>9=VJe-Og_g6)FPOG<20_8PC&8IeU/3-1b;GS;96f#V@//SL2
?600bcgU)@aKXfO6VI,D@1<NZeV@)ENJb3IU)O7G1;\X1J>;.9G^-9\57<+OL4_b
B&Q#V\D35]REf4_Z7<VD+0ZDKM&NTLYXMLF]@=E:cR\CGJ?PUb]AK7>YPXL0)#P&
^D@-(+f_2Vc9(DW1QC#4H3O4WWW:D(_O;2:1f?<9;RIW9c9bHfX#FZX0532;/S[A
,2f4I1JI@XI9@EE2Oa#(^gHF7Pg4)DH4H0PgAB&]fZIgJ3\/GGI4Nc\B2]UQ7Xe.
Z479BAI-UQX,:BX(-)A>;0aggFLeaMOG9_W-5>]a+;@^eP@4..Q?D?X^#d):_7N=
(G(cUN#2d/9-\8#@E-Jg0H-f6D1L;_>I2NXQJ2B&PY0-]&YFQ/3G-^]H;#)4?=9R
eERd&5PJ_gOI3:>FEU6fG.H4A^QB3D?AR<EV)5?W#2<71-aA09H<eB7d&6d,,#?J
eT>a8Dd8=Xb9E-XWB>Mc;UXcKgU&6[UX\/&aF#38R#X.877KEC7AYVf&&01XEGH2
AG8WF20dSU\&f[b^=6CcVCE-b5.Y<ZLP7A0&b3UO5McQUH;+,?PBR0G\F/b(9b])
9F7ZP_FagCAC+c:8;3?6;W9:]=A#\KF]MO<OB\.-]9Fg:f;^FTeNeKL556VPI:YT
Y42GC6[[aV)6ae8f-PE/#YJWO86/^9H/#6a(e[U0I[_f[c/FEaSea<MX\OPVJDT7
Y1,5/G@:\A0dH8HS,E.X@Cf?9_0f&+V##82/#-I,W=/@Ze4U2BS#aMYc&]H8S@Jc
5+@CL)]fPI7]\I>_V/<D^TH8=UO1gD.V#PcJ<RMC=J^B9,G#LWQXb+GcG7TbV5&,
YH=g&P)23I?@(Pa9,/AP[E#@fTYWYA;LcBA6S14OVYQD.]XS8Vf@S)5O>Qc]2#R,
DL:T.J+gY\(?0@,4E/VUP@_@)M8<9DY))4S042BG8Wb-\Z^2f&Va2TbW1a<3>bTE
;aEPcd@;WTVDWLZKe3Md,SP7N)CQUNUFQO+MJ.e<gI,K9L[61@/Y,@CTGDDc/#b6
=ER&ZM>CSS?GfJfJ54eB4@JfVf#)MFCCbD=I=\0SO4ZMB8c>TKQbO^ZFbFJ,\KCM
SNe#(RLd#M^Y]e&.cPE+G^+_8O01&YNE2VQ@D:I_3:\I?U1,@HM-K1#1YC@^_aH2
OQ9^IO2X,Db3/GfU@_8c55c(VV9f(>0X@0)U1E?3=E<8X&E4S#_X=:_b+#-gR@=.
+>KeGe6(J6:4E#XYSQ+:T+fPO)Q.P(-W57_XR<L<UP,Y+[#4ROB3)VK=TVa8fU6&
5DgC6J23EN?.f#_WaRG;=W:/)P[Q[GHQ6(SJ?M11L-#MV?HKa[;8Fd,5S:]&<,[(
:J+>UVD[bd_Sd4B41W(KcAg=B@Ja0@9P.V_3<.2a.JK/H_>CA-)<WLA4>[FOe_a9
4=5Bf6#c1&T/U)XK)IR5ECN:#Y>,_D/4:VQ730fTGTMOLE5DSZKZ3]\O<EYg[GB3
XeS5_CXb>L/[6W_R77:VV=)8Z3dgF_a]E.R;CPeCFDbg^ZI/D6.&61KZIV5DV@<<
gQ\?[->Bc&ZWONS6B#9P#NA<[+)K&IT#RZM]H<+GO6UbO<NbE6+c74#<84af9a]H
W>(gX@X+IfL8ddPgD/QKE0Ce=/;;+TLad4NQEZVVOYW)e:X>LWI25;FE#VbRYY(?
b-4/dPAd5?bJ8OW7fc5]>O)9aeYBdWIR4ge.,Z5PD;Y,)4VFg#TLB[M/58VH/H&0
9#>Xe13^74V\RKQZ6NI=PS1SO-dgG4^J6c^Yc[_,0Cg[II<KR8Hb&:XMZ)>61eDJ
MADS7^4[]GKOI/GUWVRAJ=CNCe\@?IQ8WF.6II]8eY)]d_LKL8HE^/[3F35Z<]0#
VKXIe9Sfg^:/J0Z4X(dH@2aBU40:Y8UPbC0\f+Z@FBP]6]YeV]48.XJ6VZY1MZ15
6>+M1T&?=2@>9UUga@#YH]LTKH7[PaJ5dR+)6HcM@EG=HYgN]5U-/W^,K3+O\]8S
_aC/\(eY9+]@<V-<X7TF[KM:.,^>S6X7AJW\AdH?&A9JQCe=SO0Z^e,+M2Sbe0)_
?WWNF&4LR:DMBV5)dC.+R,X)CCR.BcENR<?1fCF+QN#IYG?=[:TP_C=W/>af2L5+
M\@<##c&&?=fKg[;e#fIV.4DHAKFE00,85)1gd5QZ3<fNX?6,P5.)dZAYR8AAT+L
#)[]KR:We6P\LGTC&/(aO6>/VB71R/],_.UeN\K,^Xf^&Y=EQ:+?\8Q9[1Z3KY(K
aKc._(]#K&E8cM_7Y1g])SdNO27?]]CLZ1Y>G55K_2I5^YeB7O&&WMQXQ]1?1L^W
IJM)11A+?:@#X(gMe,0/AB#8B;_eI&eU8,,1&766X\8,dIULRFG1aVZd_5)ZLM_T
KVY2(DNe8I2#J4<:)bK-3SJR(M@]0D&8Je\I@J_44:(MUDZHNa0EAZ^SEP:^IWQV
W4J5D#GI9fRM9a0XU2-a;6;#)-T&N=]@QAE5O,>Z_A4<S.CbXf,GeV@-\\4B_D1>
9T3MTX]WR#\A5>4GL.7L1CQQ(VSg),e7PW>,g^\P(,cc9e4a#]cW<\Q8)UD^21=?
9J4@=ONR+IUY4:Cd\1f;6C6H]Y(FFBa34=/>0^;?+XYNHcg0dGI&AQLBe>YC,;&7
K<7T97fSSWMJU]@7@V4I+5A&7(90R<1:X1_DeL#dGH9?/fbS]7HAK.10DL;/d)64
.JNEZRLT<OGL>BL?Le(K2aR^.PFO+MM<MG(GP:d&M+/DRXKQSDFYa)EK5(^RU5H9
UE:O^]1cd-)]aL^b#3?+@Pdc0DfY:<Pa&9)bFE@a#UL@1X:\\1BOX0ge=EI_NE.U
(UbVN[J\4;?Ag:0FY>HGeH),,/69CB<?J\+73002.L]9((B85WWaAF7KW0RQ<V@K
??24>@T>-IgI?afef,1O^N><>Dg3?eMCW\AP15I:f/bc>BJ,=?&a]HE\-[E1KL:Y
O/VAD?6S,BIG159F#_WJ.&YB#[(ONNb924SA9:gS&14=4OUM\>?aL71gK1&_0N<R
RI(LcR-Mb/Od]Q#=;3KP1Q+0-Fg5C_b0:;e.55;<eZ8BXWUI93=UTg1dKcQJJ<Bc
1f7QNI<;N#-ZRe]Z?LRBbB:J8U?67^0Z\@YZ(B(g-31)K(R\M=(K,d,&&:N7B@fI
;_e7SK=@65([g8Oc]H^aVA5ZIDa6M@1=ZX+G#C.2-Z0MDW[]+V1@]WV(5IHLc2c9
H6N@6WW[gFC.70/,RKXE;P(>dY)@>W]e5JGc<DYe-<?@++,=BLE@8C5MW73WKJ(T
\g=cV#P>W3_,L?TVQB(I256Q&_/6MG,YZ,)X?-FXTfAQANcd?J86.@CO6;&TD)S_
7Z4C/&3XM[C1\71#)JM+gb/^X&RgeDFRTHKNZAK7cDV^ZT-Pga+,TM>Kd@.SL<;L
U08\;/UY[?/Gg=1-eP;FZPX48(;BLcfWEI;Ub&@(MGfLJUICL^;<FA.H0bC1/f_6
,3@4<g0(RYRQd(H][PMBd\)L]1;>)V[ZWV0.1S;abT><E9[E3&aaV?<fA49^c]2I
5Ja<S@(2:];I-YLOaWR.P,51T7?Ad^4Cd6Q(O2+e71cSIHGFeH+L(Q/g4S6^[3E3
JMf1(M0WIN,G.0S:46>1:TW.HS,d4(/^>6Va4V7]X:9eg4.(f.0KAO0B=HA>\<P;
>^._bB)[K-<IJ(_=\N99g(_N4PF-EEd1Q1[Q_M++MUa.FADZX_IK;01gF4aUSU=F
X.ReDSd[UDBMbE[.6-S7Hd2\Y_H0((2#?7E74UC&O):__ebB<MHX&:&-cD-e[52B
4+>Qf.YLT?_TI9:WDe[ZF4=YE8P.JJ/AQ0f/LgT3a9/caOH(2[QFJRMXEHZ_IAfQ
GM9HeA:9@+ORYacDAZfNOS>PP:Q/>I++>E0>:3YQXZ_^LUA=ILA26>WDG^ST(Y&&
O/9E:NX6Tf)MP&#0>JA0Y?=CAS0TLSONNRPZ+,JFP,OU+c.90\.RHJ^=IEE<[:](
UN_R7,>O-75PDa:60:1WI,H1cS7]PP-Ab>RCM69UK9P1Z,A/V?3-?@PKTE#B&Xd2
9=BdM]d@,cH-^ABQ6>W6)=F9>,A(bT+8:PVf?IH?0C9PSCcE1TSOC(NK>6+NI(9a
3LdbaHSEbW;A4G.#KTQXK#+NEH(a+fKI\82;,7#5MfNI7gED__4K]GVb;d\-B/B1
+710,3T9B#4;NEEJHZS;e#JMF=_ZgQ8H-(H_aH?C/ZaI44#0V/7EY=B;#/g37-,Q
&7JYF7\OO[/#+g_)[.M3RM)c,WO+S.8U52=PXCC#/-#Q;a/BC2^(WP\J0ZfP<[g4
2LNgC=gEP1.[Df4fER<=EFED#fa]LP&;Of=3/3Tg[DeTg@:1_)P=G8gYQD?;dB.9
<.3G/3&H#[V]E2UR,&dDY9^,+V\AE]\OKffVS?E^R<Ob,:9.MJI5.7NDH3=J>HYQ
@EQ[NcLL[.2@-AL;EC/9-C1L5aPW#\2LI)HGgB9fb\cfURG1<PcZAE:^:+SSA,a7
V\HUX-JQ1;c#\E^M-)U0QW4c)]?<RNY(c\3LGIKLS:Y&:23N;.[gHDVbW/#2,U>K
PI90)LDb@S6L9-M;g,O05JFU[Fa;=Ce?Q,VVWE;[cceP&)?;_\FH=,HN6G<BdQa0
f?+0:ec7+I_E@8=H;?25;3,A\T-8B8H-e8(c>a#_CaC;F2:Da\P=++,+:P#;Cg>B
XQY&E>]Ze2/C]dX+Z47f0f^7aUN]H5:4AH<8>H>:X-HTH-5f,2Y;&Lc>dQZbMSU8
2#XAA-4A+c9S(VCQd6/b<X^#EU\EaG;Rc/2bS08=:)3?CNCEEH#(&f/9.7I2E@C;
^[QF?/4aYHJ/Q@I@U?f8(EF1Ff5GK&7I..Ra4^]Qa7PDE[/7;G+bCKOT>AE_YV\d
B(a/Y\86PS@5Q.E\cefRECb8Pb.=a)OPZ1,EL_[RG@28N_9b922Bf6,PFd0_Y@VH
aO;7dJOPDfXR=HRG:D,A<G>-5ZV9c+2(f5NK92@XR-.OA<e-e?ALGEbEc2CX95f7
T2VG:g<,ID#5HdI2??2O?H?+U8O1+OT3[dK@LHg@CH+D9J06XL(PD46PPA+UECG[
7a=(g-22AB/CFK3B8&_;Of11TF1\ZRM3a@.[#]0g?_7_IC@ZPLdE7,-=K[KW&KNF
C0&RaaS#V)VNG411U-,ST(;#=M,C\CG+QJaU[O>L6OT2VDLKHNa?)5:&)@O\1MDZ
<ZTV5bdSI7=#,N7R8beZ?T3:II1ee;G^LEHEPQ/>6GU=@T&=R0M=0]UMRV3KZa77
4+5?LIa]cf=?UG#&X#9A4]\ZX>=N96a<T0A5=,1;2.G>EN)9G/OLY&4+C?5gPF5f
](DA,JH?R]D6&?(KPC//&c@UG35Z8P55UUW-8,4HQLcYS@1dVMT6VR.B/9RX5Ef5
T(KP,;DEBd&PO(3==UEYT][NPF>EK/VM.,Y8]&RUWd#fUeK7.^_@WCFaAR>)1,eb
IDS&Jg97gT<EZHE1\46g1.Xa(&B0/@Ndcg-Z+QYe_4#O^ZZd&J)CK<[D7(9L4_Z4
>@7Q(BPZ_BEXB]9V/,Jg@eY=3.Q/0HdT7&1gWcbTH#/S98&g_[]KGOf2VOV#WSC,
-:b>7GG2=6f/C(bf3^MO&-@1HNOB):7\[H2]9:SgX^.<Y>RCO-gN[&,D/\ZIB?5F
?_SMUO3Va1X&gT_(ORA5ZF)TLfF;aGJC6@17.9BD615(c,fOQ^BN+\gB-08?Ze2[
&AId<[OV^SR4.bR@0D>J7C[6HOMR[726K.Ub,7DC\#DFF5&eYgJQ(,TXG)MI((,<
>IK[UDfJ9\65Yg73X<6^LO:19b-R0fNbI<^1P]P<gU^]QT#IF;IDg?50\]g;J;>H
_&NUEgS_AT)bBX>#0_SZ1J\;E&+1eYG,G\Wa#52IMPTe^FX4\:Bdb#f62?.>M#5V
73=L/B<\=RYeK,<7C;#\SbFGbDVWTUYJ4_ba4:c<B:;DbCXJfZ&b::1JG;HSJ4/M
GR,X5K,67EG0VK71DeC2:+?Q1&:Q-\=GAeVFB<3cSH1T4e^L+&c<N>NTf^:HYI>b
ARN@N)ILWJI8OE58&34X\@]g^Q9aPS.Pf_M8B]44&;d2[W9X<GQ9]6^TD,dG;I^D
6aE>fN3S,7R2GSML\g9cQ];P1DV@ESN[8&6II.^O)P)0]10La@\\fd\]K[2&>8AI
@cT.dH(@_F#57]K6)P<X89e[\/7Y;Z@N/EQQ<5F4Eb:0gPV9\376H:K9VNTg<.J9
IN8^/&G+RcIeOB<DK4\a?W7J:fMOAT/DIM\P.[.VMa+O#\J/J3L2&2X0aNCR]77R
NU_HBbIW7MXe7Y>&G[e(RHHNIHRb[O]1D<@+bLeP3bYG2W7XLVI]4F\(Q-ASF:.^
56;MM/DZ\)KR1<PP[?A-\C>R]?B39X8U2JP<:gHd\_N;#PP7[;OYPRX>/OdNT<H>
=BOD@D]Q<&,^Cg)J3a&Ee97[d?54]BK^Iaa(I;#e]/CDR8g1f=SEUKQ=#B6bCW/&
aBE^e&8K27c]@F#_Y,R[6d9[a7?B__V?:@?]\+a5G?NQ\IBYV>b81:H4g=&gF^Ie
OB.D;IaQ^/W(W635bAG8]Ma@W7A?Y[K-g===H6J^04V60ZE>HI[O/=&#NGI[;-f1
TgZF=d1]e(f;NcfVD7LeO^C_OIR;9H)KX9=_7;>QYS#.ad3Md:9RHRTI;g^CVZ4\
+:]BQ=A,WF(A]+E]WZ&6bT,UCW=>c;24WBEW:7BU-dQ.NW-\1Xb2D84[1.#&7OQ-
W82LO67/A-2H5M<P6U1CMA;XG,)&2#)RF/e8&V5X;MIJF;7B9SdJ;06P^b9VB=BO
B_B1Od8;YKdI<3K<^4/PDW-X:1)S.FQ+E-OW484W7]f13@\/;QEUI5TT3\?@FL2#
GTEMGfVd9NgaeK(3G2J(I_f=,OeYZNJ.Db7fVAS^aN^TV9:G?JK[.S#^5R.aX/^5
EfNO@TH(I_;g7U_ID?LFKe_RH(47V\,2OD,<8Y410@:TEBAHec=fc:J1=F_EY=MH
53Gd61=a7?cf95Z.Y_SGeI]+HF/\PW^5#4?7e]D,)LJN_Bd3SXR7a[5J[,+1C>UC
2LFMa/:X_-UY:C.WcS)<0:6:c9XJXRH<T[gKB@:42HZMES[/(E]8PK9(LH;N3UF4
<GIP;U>eN-a,a/A#6&ZU793&HTG[1-YR12+2C,.S/7XUA2L9MP:daNK;M6>]<N+a
#F@CD03O7Z2WZa/AFd6.CO[<\6\;()X6egX2R.#T6X6IGa&2G&T#K(UTcZNg2D><
008A=ZTAC54/F7CMYO/?5BTg01XN[XY5[bFc4)<(O37a<ZIC\&a/0cW(WQ-Rg>ON
^10(AU1Ac7KQ.)8+L[\I4=E;>gL#d(RZ67#b+ea.Q_03f3(6EL]-T9+Hc09UG3R-
^I5/GeAV(W@6?V;_&44LF0AIF#8H9()2JDcb;Mb.),Sb<IR4dJg(NXaP.H[dGQ#X
6MVM^?UQ]3dBgLQUHHbT,X[I9GUJF_XO_S9K,E^Q?Df:U@DCgWR&36Z3;P@37Z@g
3A+_9=2P+ZfX7R#:)<eL,(=WgTVW[/bNM^CGc>,,4ec/VZ7E/=/;+?A-^;BX5OQ7
&J@CT&=ZWg:cXD-(_6H/_(M?X/IIE1(@4ZbNb;/&P1SHO3+Y0<+6F^eTH.g>#3B\
-_E1B,SZ+#?e:K/5#a>^=eQNT\HED<=gc0_<9G+V>V6,5cgPbQTF#YM8gZ;QAVf\
cP6Pg?)/f#54NJd9E(Ic]6?>D9EOf\07)RPb,>?B&E66HCR#L;c?:5>[gA7RfK\3
WU0UYN53aY,&\ULAf=D]65cB#N]/LD(_ZT]<FF\X[=GY_QP_\J))6bLGPOgA/JN:
5;cd^9\#_6;-QN@U#(L5NM(L66T53OZ8E;=^+TLT<85+XMFfA:G,OB4b9?J&N#>e
E1b)HbJcO-.W2==G(JXf=AKR42:H[K-UBeeDNSV=ZHIc25WFJ/K[)Ma]8I1])503
6eU+DP[R)_0.Z+g5MS48Y44b/(BbYRPN&:08<BTLD(2]W2&5MJUYBe>:KWG/[#,c
&/ZUd3^(XX-6^R#\bHYaa,R-dD(O.K3/aIT1Z6SX-L<9MLF>@M3SOW[F95Q[;2L@
2^NOE-]=Od0?ONHR[1<EB.N5DfM3)45#0S@#Q6e7LQVb-aCHESH,KF.I9HO62d-^
+8R?IAEHD015[INea2c_3JSNYgF0<)6KGLL<;VEZV??,^c8E7-=/R629JR<.dPMX
Z@JF4dPFRcL3XR/e8Lg-dA3GI^.ZC<#VSd+#g@_g)E:<D/\,O(4#P:;fP\<)(PCK
9:-PFT[fP==I0-I(g#Z9CQf#2<4I#7ee_6,LIZa>SGP]dd(0;<b[bDbbBDaa=):U
b72eY,V(,S6)S6=:/e^3D6=>-P8a+<2R);PV)Q[[De5H4.:F24-_3DBE-KgVD4d^
4D3Vb#0H]@STIXEPEL:/)eWM;_?#XRKAaL,TA^]@)dE8]=agQ9JR3T?F>BK903#L
eQRF\CJF64=M.146fF<b1Mc]X+[M&PaeZBSKWXZI33N6IDEHa9bM4g+8FW8_NfLA
77S>(B)4/ZH<X-.eII?&.Kc-/DJ+9eeN2MN.U#Pa[GLNc.NJXIT[+6^)f-/Ng3RO
OZ>,d5a#Z&,S^[Ee)Q=2d7A?B\6Y;7ca+FVZ3QWU#b:ZgPb?N1=dVMgdTD0U4_-Q
KZ(e<2K-)JV<&6@2-_eDN15faCLO2FJMdJQ]A>aJ_dJHd53)]CLY.JXSE=[]9<IW
ZDBZ8d;R)c;^G]]QY7F7-F-9;gEBD#0=\;5;B\e_U7YIGgUO_eCVB+GH=d3GCXIO
?@(cJTeV^gUM(5bbMS\<(6BHIHLdCWNRXQFJXGN&@UgJ9>U)4\DSG2W1#2.01R?L
Se?)=(d^EW>3a?0,WAL.A-R\M]NC>W361=JeOZ3<-9B=4&bRWZZ-I9fLZcNO^@8P
QN3=AQG#F\gVZ_F@(3T[W2VQGDBILg4<KTEHdg1)+3[D&ZF>0d0T,)c2[PAXB[A[
7A:KbO#K:1.</UM])4B<<KWS<L=#FWWd5K+JR6))D7CDdGb)g32@Af7XH0.9@CJ,
6&UC)^VgX[?YZP##1,U+EJ5J=Dc]eRR5:B?5ITcI;@HRaGgG>c^2F3@+9B#_ZGFO
SP<A5^4_L5EEF&<INZN&[Mb>M+Y0@>B\1X#B.BB-;C/^AI\(EU4#U#7#g[7_>.;<
61,6L:9I-ONdff-V;&Z9&>Pa(TV7W4D-W9NMLK]?H8JL^GKK4@NLB?6502/>ffNM
MRKQOMA/M9;e^<HXA4a1VRK7.D,8TAI+FZ-@0.-&b6X2K43bd/H68F.g?A4<=4/0
HCfF9e(6Rg&Cg>QZV<W9PV\_W:AL,62;N\#D&G2+V-GAUYM2)B\7g:EL;^eY>59X
?]cEW=/UfDQSBKcED/5#\ID]2P5C3P#@QZgWW#CSUBB/J<78a@.+XXZcM<3-3=VG
?G(&DO1,/=6b=GKEH/g/NL-_e;_-7@XTGbGWb,F:,1<3DI.aa7:?2S;[aG9,,^S;
T#(\O@5QF9f):V,&LBVEd6(J])K_H2VD2L4e8T-)9TdXfGPP/B[E8);/R#E,7:b1
7VUXCV>?cESGF6T^>bUW>c103U#^YfFYg(+3E8Ra_5)54?.A)51E]e+0-+MdEB)9
Zea.JX\-4TLFgQU[PV3B?\]1FF?aA=aO\_/S&Q-:H_A2dY=g9TGYV4fXFC>(9PTX
Sd42(SgKTF;,@M;0dIYF?/NFLf3[EX<EBYSc<D+Bd=NDVI3KCT)Mdf/F2,5C5YPU
T-G?P-WTFM.Xd/GXb=g622=)7aH)ADR[3JK;/W4#QZ-Y<K0\<JcAQNgDF,<]+]Q_
,TE#0LJ\S;9aC8\XW/a?]GP^dTQ8?E)JG7W;K29cHF-U#^4-J:W,9\afIRM#VCX]
4LWK_^<g3&.?24/YU4:0M+UD99AR]Ngb;J15OKET-/Y19)cTIVbSc1IYI67a#M.4
4Fa.VYXGBe#HH(3).#+5g5=a@d#6.@N?gW;2&Geg2O/\7-GK9,e5]]\=6eQK.^@N
<2?MJd2&Rf,AbV6EF8O9UG;W@2X=abb/]Oe@eTV=A6DIVf\YBG8+;RQ+3J[P[33e
713V=?VR=(HA&=Ab5G?QINe_bXa+_T^F?0OAS2)2BY2AObaYb0DO?<_&deGdQJET
X8/>#dVG]2)Q_+W2?/a/_c4C\=B]X[H)C1J\E2eDS;.9ZMK3.fL;QYF>5IKSLL>O
fQ(-QQ;@--SOQH9AUXV,./Db-#KN.d7,5UV=]/0(<&>2)[HU[^&],RT.=)]2NWd[
T3F+99R.aaP4(N<f]O4aX3e9O8Q:X&1,cc;AfPfHAO1OK^.VKP8ZX3+E3Ja2:XMe
7>;G,<8>:/^YLaR,.YI/=WC:58PF.DVGGDb3+d13K7M8_1X=>?:CKZe9Dad3.-ce
0I#+04R4/_7TYc/6JK=&eIf@F_f,^Na9J/g2]HU\[,/&a.4^b7aN];U[--\57V9S
<U],A,9P?M#BHAe><c[S0:d9W#7CYI[AL/KQ1EaY[a2+O+I6KOX5#6=HKXbF=;M)
ENT=F8NXG_Ge8B,:;G85BdJCgXe5^Y706cWd\<b?N;>Z&Y\d2cK3(fWLT8@eO9^3
.>4B2UU50#fI6N;+1?QS@NQG(7IUW[5fYTF/I?(>7TeC_^C^ZS;/;Kad@9\M7LLV
5f801AI2c@:.c7(,71UZ&Qe0SL\GNWeM4NB<.L)A_W/?_(XZ)\H_>f(L+7ZZc>DA
bCU^;XAVF;#X.OLFRA23TB35Q0c7_2D\OHW5Ke]e/;K66EE[1=G^YO6+7a+&JeS,
@NP2_>KR^GF>dR/3eJZAY=FM?1Q&/3Y/^/?T7:9Y;<GeREIAdGU6DaG\V.TS:1+g
:VD)(^Z/32/B4NKRYCf.:#N=U^(2EcKGZYZ\O2gafa9/eKDQ:d^-7JT&HX?M4a27
X[DU.U><,Z>_G69eTb@DL;bJ)G_.M0;FaH,>K0cEIL9=@3@O_IL/_e08>;cB^71P
]G92QI2>N8M_)#NO9_g;8:1e?f_a;#_3U01HXD^RPNOcbIY3VLR\5ZXCJL)Nb_3>
XdXT<fe5gg6QQH>HSgWH]5GUYSI(A7-)g(FF=;X__S<^Wd:J+0?EF,4FPW87&U\_
1b5EO^NF#@EOY6WGP/OfH>8YU5_.^;.[OK1IS=QWfg[&(3C=>\dDP8d]3Y-F=bbF
Z&=U<ZS7.5IeSN[Ug\27&LZZ:FM+S4\-1C<?=9T]Y78X6@3>,-6eXP:O8KVd3JE-
#)HRM7Z7d-Ye=SJ3XXE8-]MP>68IDV54Y3[,)D;^+C43UEDV6g:>V?>FDK\Mfc8#
]\XFN5&1AXFV75.Y>cG7a-9K5#3f5Q<f^O,?O5(CX_PMK<:gIJ,eT2@4f-DPE4M9
>dQ96ag7GMb1NK>R4GRA/EQ=4TD73.XDQRH>Jg9D/\E6VNCeJ(Xg1DPeHWOd+fcc
6.(K?4@GKLE;gf@K<^LX8)YPJB9gG+OX?c:\]J,+;-Uf(I,4a_G<<JB.;L6[75/c
4DC;V=@[_#UT/#X9S6AZC-)b_bJ]-(-2.-/_HB\/6;f^Z_+02(8.UK)a?X0;/F)S
JH9c:3OfEJ<A-8SO;.#3gS:CFM4?4MJ7_0M+/B8(JR4c>O-7YA-\a7e5CF)M64>\
>\:TO^6cO.RN]XZMZ1VJbS]W6aHUIZQA>\dEFW&59&-I3[YP8Q)540.0IXS3ZCMf
\,B.efP0b9XKE>#RV/;]Q6]\DC/006/FR(EQHXOO8_dKL]5526XgEQb;\:Y9JL_e
UI7[dL3e/]#:.-AVYDf4/Q7BQ;>ZLG(?bf(Y3)U?4.H),B;><D<L+ZW,(dfOQ&-S
UdI5>c;Z&OKSff5Y&9+0c^d45G&gD/:GN3\.8D:=/PPM+98cU,UPB=(1SKScG=6.
_7g#V=.9bQYbWd4J<=,WJ&B2Td4=bc\T:=a7G)e1^?TU_Ya;+&5-43+=(d0>8I+8
-::2V9Q90.?dSATT0EY5^a@R]=ZbU01WHK(0OY6BVO:7eI._)<RQ([&eF<-gf^1>
@gHcK=b#?1E]JII#bLa/<H:UFA51D-0Xf_5bDVQMN+;)01+;P]O0&SF4@IX0+Z#Q
C>JN=5.\R=Oa;1<9#bDG][LG?DC/:+50V+S[[RcJZ&HY]W\)\E5ITY@-G],>g19(
B2+2fa[@COQ(-OH:;_]fP:OLg64f0PQS2K5KQ(4-H7_N^70\&gABb<GTI9\>50]f
<NRA/=0@45E77WPB)N;.9H\AKf7bPY/M-@:H\CUW@#BU/R7[UA05PZYM:LMZLIQ>
-1bXE#R#;POE8209+8dO(:3\<<dZSY>LdV9I<,N<7OeMOX60IZU[b_:F1fg,bO@F
RbTGSC#.W0e)0Nc7;+-AFQ;<,=N.^Q3>R9@d)T?b_7DBFUSX5/[BI-A+#>?#8gIN
^ZYdC&Z3FF1ag?::-/._0RIV_?_0Q]@O#gWbV3S?WAQCNI2F<Oe]b&PO5#;.AA2P
2/=W-@=+/(>JdG5W\K<cA</\-J,.85d@<J\S1Y1?#]KOX\f]RLK[\>85BDe9^DU6
.YUAY_,AEJ#FS[G+WLBJDARfD5P\2O2I8@<Cb34S0L2EbSB^Y:[BCHebEKI2K2^]
&,6MbG\P@a>_R/SG;HC5KYbg9^f][M67STdP84&2+gP](?fRM6CB5[]/LC/dGGDX
^Vf/g#<,/?BV?^]?,P_]&.b./\LbV(c(#)Mf+0fa=3BJ[-H.dIdLQ6O[Jg/cc:ON
QF4,MN<5fD6U8Y7;AWV-/>.:U=(=<b-U>G\A12K)FH[^\88QE@@Me@I)Z-9M?+Qf
(U-D:_J-aOE4IfP&PTQeJD>.P1\W[&O)eAY\>\;;3@Z^#2KBYE[#HB]Z#XWRIUCQ
[^K\a2b25=4FFQ8Kd[&T3e1GJGIQ.,)2bQ20U#X/GUN)7+?Cc);_&TH-C<G0;2Y4
:S0b^967TaZ@D-GV?B6P-0_V2<]FgfW1R3QbV#396O0;E^a5a248.]ZXY/7g:5EM
\)JMIIHbEd+A@?M5E<_+H?X>(-3e_98;U#>C<[]H:&&;Mce:F5JSVc#=&Y81&[bX
SII-396;\<M--HL2EG?D(&a8>B+IGLZ#.;A1_;WF.?W7BgEFG:=V<UK\P.T,d^b6
eEA=K2+_P=ae6O(,X^V#XU_2U5J9O0Lg24aS5YUJ=@0V.WX65C&F)AY?\aK4I\T3
)?E4B3-IC5:S-VS28&f^4,a6g7R&7Ja11T#9LO\>?U;AKF-X+9:PXSUCQd><6;O@
MVgHYO?AO:B7dF-^HMV8;H-VE=PW8VZD#:VDIA&U-OSQ=IX8#D:/f#.#e(>T()Q0
b,TBYQ(()\)=D/B6N9W&eFU3R(2WHbLdUea#+PVaBRR@FG>=Ig-)E=72,g8YfO-0
6/X&EA[9,.&/CeZ_+VG-bV.@VH7U)SV?BPMXHSQUA?LWQPB<XCf#g:#T.\aCM.(H
8-C-YVO<=&a<=NfC8VTFg:E2D5OU0]P#R+7KB/6U@KX3?O^7d_;0,\fUM3B0:Y[[
CQW5CcHZRN:+\J>)f)MM\UdeXf[Q6b)3)ARIgN(^:>b):L+P_LEIZGMLXK=R<?\Q
;UPf07NIX7M13M^b_J?8]+675;Pg,W4_I.df&=K]c^@;=JWXW+(?3?LV2d(N?QG]
RI5S\/;<?Jc9e.5d/PA8Z5e6fTf>gOEL03C+)/R1&WZFe#Da:;Bda;MOYc/6bG.8
,0LOBMaMB+8W\9>9;UDJ<-P#2_9CDH<-=U<JQ<<KYOW/M;/11T2cZ^P.C25KJ:D]
ScV+6KVZY=2S)+A&d7+0Ae[MW2JZ9?UVFg+4&C^5OFeGB4,+4AGC&2?]-A1\BK>4
+7/<M(\2+bM64We-QN-eP3b^S@5ZT12&2A;@K<7SX_#NG72VH14)YQFW?)HWQ;gE
ZY]Y]]gTE.Y?[:K4&KK>M)^gBQ[VRC#27RRE^9\0JI[(B]7:aa:B:@KgHM8=G#(T
1Sb3.O7)ZA:c]K/M(GQ&I+:+LEVb\BT@=]gK#UN,94&X<VOOQ.1^OP]c=-Wb)0GX
cYY=<BPGE+A=2XA..4U1VNJ9@<Id&V60cd;2ELRUN@93>00U>\dEc_W<+a:_X<YQ
d0<&L#TLd+e_]X+_5;f2R>88(D/?RKZd)8d<,PN7C4A^Q9&<eM:A?PI2?AbYPHV#
P8EWD-6TC\8R#T_Q-4QCDgP:VKbX:2P+J\BEGQLLAAV(_]RbRdZ7,G<O/Z-]1g2B
;BP2GO,BEKP6CWBBc4@@6;ED.8I0d#5a9GGNC<4b(:_f81Q@9VB=-ZBXICWIaI<?
=PcTa+O&HFKD9H[DYL2ac56RKY<M0?G[+TEILbD64QaA]NE\?a(GF-Gc75@82#KP
:N()ZTCW?5Y+UG8#-E<faY@V4FS:a>bOV/#Q@T.D8^L0KE#/S<?HZ:Bb#R=R.[QR
9_)SI/,ALJSd>#Z?6B-cHd&cZ@95S(\@&WL]W-<3E^MF8KJ3;=U+II(E5+NBBaAM
D?=8.Ua:HIS6a@@@2RH>9Nc57SfB[QLVV?0[5JbJ5&^4e12[:]5_)F9-gR66B\Bg
:(/);Fd(\[-J,MFXg<Q\F2^CEd,[GaB#,X)DCNI(?\b<EQY05e-81L:1UDYXF14K
IFX4=L;K:2Xa]>2bB,\KTF+;^]W(\Y>:LDINZ+,fBQcYVTd<Z@2J2ecMG1_=WIITV$
`endprotected

      `protected
dVd#QU&4gLU+/^L8e]0bWW5fJZY.JPZWD^2?KN.HFTUKc;3eNBB]+)#>HHUGMADS
0Z8+JH#EX(B#GGPP<&QOG25f6$
`endprotected

      //vcs_vip_protect
      `protected
95\9Af&XXFH@FK8DX+eZ#eR:ZZ^<;M.31dM#[Af;E-XLNd^3/(]+((I9_GL4-9I^
BMZ7I:1I0V:I3\I7f]g19LfRYP9Sa7UdT^b.N#>)@Q</,.62W8RF[LCdT6Z8S7bG
_U=;&53.AM=;W2Z0^FU>6Q+ZX5UV^DM:eV,T<GHaUE#Ic/)&TMJPOF98OHYTH\>C
&FRYOgbN#8582fXDcYUZ#-F=U0/AM7XF4@7DIS5,:72Ic_B02cIMZB51YWS@eg,\
CFB4PQ^]e&@G]VeMG/)&(gUHQdfIFX4Y<1F87Q+@^fd3^]38&4f^NQ>UN+Hg1#KK
Sgc1)U:QG>?&=0V(T.OYV9H&20AF4[OC3f(aBV\XQ8OA^N=(J4S8Y./6>WUb;PgY
gP6eC5<cG.MfLG<[\1S@8/cg;;;;#(g?HUWV_^I7QLZ&4VdJSS=OHQ&M-YYBN5)&
J6+AI5S#f0V1+gI6UNQH@]QX/aV2JFPeb4.5C1UT6?-,III#,:ZD(=Fc)eU2JJ@2
FUL0f1-K?O[9Z+6+DG?.E6VIN=(PA]D\-M&,=4dPS?7FO@X;TYAS9\cARXHc7FI.
B):G(-VX[N&6Q8\gC&H]VeR(FgTH1,;,&O)\\B,385\D3;.S&AQ-\Pcb;V8N1DL<
7N<5+=VcB5/M<+G02WMf\gYb-HP83R1aKHX1Md@ffIUD.f>KJafJ(2<,4f)2Q6RZ
aLe-0/9+L)6+6dQ0deWI-NRg3JE>URQ;P+UDBFI6V0]3;<>EbASIZ):(QE@+<Kad
PY?W2]O))[0WT@;9cX1&ABM?N+8ffIfeB]KX(5I23LdO5BU>?[U8O[bKI-G/P9VL
g;92-SP,ZQK0=>\X8BK^44f[M8M1J+^.NeOF(8dd>23\_]]U7T_J=>#92C[VI7g/
F2LgRM[[P/;@P[>c939=Od11L/.Z_BgF:T@Q#?aFV=cCU=,bX-G0/+3dL.7fKWKd
<I=)H6eTZ&3Ja,KJXH,B4^&JFUfSEB,XKYM&4HK@<YSK^J&R2b\gF<3LISG^V#(Y
;3Mf4UI8?a\>YHdX8A9?d0dN#cPO_C6eYN)7/EIb0/:F18;d=,NI4.,JZ#0dHAQ7
2G:8YWP3d#,ZLAXdUXZ[1AGc2:9K[0,PU8fA_C;2aULKHB-XL2gI03:VK_OLWX3H
>\L#eX&A>[>XQ0)ZUFVR=ENVB67eB\5OVVbF_aKE+8)Z)598g>G1=J3+M8M-Ne_\
FL;-:[6P9_NS#Y=^U4&K)C>&IeB0V?Q(Y#M8ZVID-(/CTA1BX.;@H4C=BVFGH-NT
BXGKPZJ^W^C(T2WE+X/-@g^?GR:K:=R482PC6>6>T+3IO_ONQAY153F^G._f3_(/
CBTF\FbMdd:FU1gN7=cCDL<b?#\=#eG-#T<NC-8YB_X1&fH9L8#BWY#-7&2g#cCe
2,]Y^R&0S+&/RIE\,TCZ),6aTgGE(eHF_^HYO-B@@8F5]E2]OE==Jc/Q2/TXW&Z>
S9=CPI]>HbXGVSI+<,^Y2_7^W?26DYcIVO[cc(#9WSK2T_(ENL-EZYS)2DW,UG;:
6II&Y;).2AedW&G,E@JT[./0XabHZLQ=YGH4?EedBOGTXYYUIc_\XD@S+#f1DCDa
J6]=>Sf?MF#00<P)bGP0GTROGFdFc#04bGQK8=N;A:\e[d>?(MS;GV>IMD<1C>6<
fTa6eBWQ6Q]D:R+5-]];:W7ZC08P>aXGPIVZ&?1>bAAf=^S#CgG8UfVN8N#>e:5#
9Z^WfVc5JC[S>?00e]RE0fd+U]E?:[7:8\;SMNR@:HJ]NP^#gcV:P8-3BG8C6?We
::EQ89+PY:Re&J\L\>Y27(///VNE>dPE5Z=U9A(U]55[[0+NM)[ZM=];UG]@VWeS
--A>d1P^S.HWZ7Q:eTK508(eA.I2TEgg+1PG;@/H=HUZIZOK=4Te.;U[LGAg-CH^
FO=GP^;23VH04D=9F1T#IYM9I?IWH7BOJFR@cfg9E#b/<5WGV\=W9Q:bQ/g1/\1-
WUfI.g\XQD;7)8.1/E8<Od.W/WZ+MLK4\WOd):BLTCHL[ggZU-LR&+F+L^.9b0#g
-,2HXZ(P#;DN;,>ZM^Kag-J]gc?WZSSH:c/J_5Oc00:ZK)KT/R<-0bHP@J1Id9<6
Ed1:V+8@IB3S5/a3)C2AI_9^/e<;1K/SO-eaE8a=0ee3&^73UGC/#)HPJ$
`endprotected

      `protected
ZN\4V>KZG35>f_4<Y3:RWSXDB(DC<gFdJ8eGfC4(f9P4ME>D[TfQ))D3O?NC3)93
SXAC;K\:aM\5YXS0DZZ8WaXD6$
`endprotected

      //vcs_vip_protect
      `protected
[Hd<ZAIfZ=U&c9b6@94e)K1HRU_+(TcG\^:-^9:=IE4Y@7/N7C0a)(Q4U@#@A<CI
M?H3EJWX)Y,G]P8\GIU:Z[WKA13^ZXV9Ac>T_5-.@,63>5QPB?:-b42F7IUWGe-f
0;<L3@5CeHY<G1&GDM2L7FJgEPU[_5^Vb81\X0LM&9(VH]UI[Sb?MZJ/U:L0(?^W
K8H4C+.WT&e#V(0<b&0cUKON0I@Nfd[[<UcC94Xe<R1-@65::1#-1aD7YQf()Y.g
Uc1(R,V]I^:93FWJ(1gPS6NAM6&/++,&gQI>,?<P-<cJ3=L#--fcPZI&I4U.1@;P
aLAY4G?Bc=I=YB/&K;#:@dV]P.MSd2#GIAbH)9#TH<8EfL)>;@T9_<T+eHa&5_X@
>A<X4M-R;G@-HUL@(O&6CEDTYAbgTUbD@::J0+:DgFGEP/4_f-L6IGFGWZN#<dE0
]Ebebb2)fc,SDK17(VNeEgV6#3?O+dg<Xg8,#)Ve0IC^GSCCL&I@T^-HKd1(51X?
=?7(?-=?);EcC^:UG5NGbVE_ee9X[R:#&]BJX#Ra#75\#TVL+Y6JcI@?.D84[33d
e^QW<UVSMbd1XR+Q1M\b;Qc:/M_gbLSBB[ebK,\AW7d6ZJ6ZGaeALS_Y./<APXOV
6R;/\HZaZ5GGZd)YHBBb(K:6R:b0XO2R)&f\-DKBT+-+e+VQLa;COg=?DX@<8I.;
DKIC^T;;//AJ#V3WHM&B-D/K+@aP+GLEXQ)_\+2=:7>?GGHV:(AUcV7HUb-2aV)D
eSARfZ6LBgf^Z>SIb-=[[^U>/&2d26.^3>:[a4Wa7?R(4+7]Wb7ZY02GNA\eJ=..
JHPSJ..O@=[Pf+]<?-IV9Y/Y=(=Dc8WC+O:IQD/B1LL?(&#>/NPYGE]=dS;VPC\C
RgV^U(.:c]>S0NZ_M4S3T],)@:R>\0^.FCaZVf/f2:TC@[2N(+=0E2RZ)/^5g<MD
589HLNS7+9&OE0?Td8]SZ@M/+A=0(DbH[O8<UPa/?L7N-7;M6/1TeF6Z?DcY&,&\
7^DACOTg;=.YF/X@:XBPaUWWYI>04JLH@fg/#YUXRI.:+cFFOB7bWfK+MfaXPcQ-
0<)G_Y)TD?(1,Z)L-2<_((?Ye?cbVeD@-DPBGN5D2a<,\1dCb[U:LK9H\D=OA3?Y
NKIAIC_)8M<QK(]d<eA7&cId>W1GK.<PF2IQ//8CfA]@B1A8_Z15g+@EFJNX7>28
@Z?@)[#HOE_eG3g>5QY309BX:^e>U(?98OJLD_--[O)KdY[P@JSYQf4G6U#\6Q;[
X]+TEaGXJa8[Y3:1,OH2.&[IWe0aA&Te\B+)N+ZfYY,abdE@Z#[P9d)THE:Lc336
DT/<#E1JeIJ=#:E=MM#(BG6dReHc,F01&7V_Y:CP&I@--020YA)UQ3@DgcB55XT4
N2,0LJ/NFL:0(B1T.8D9+#JWI00ZTNcJVW-\N^I>6c?C^_&B@BF=@[>cC#B@0,__
EMM#T15_IJJF@gZ-F[bP_NTIdC@5Wg&S/]9Id2@dUV-QDZ[JX-204,YXDK6fN@A6
+)bO>^Q4_.7Ve+LFbNWa\E+;+2,@,C>a)PA;c#E/OG&>Q//O)(3QKL#P7=-SZL:L
LaNN=QNe8E&EI-9-5<MA;Pc1:Ad]S-3#b4P/gW_8YWcE?(WH@VZL]:_ETcW6^:<]
<:4,W&dG[ae\VCL.?:cC)T;2aGRS:7/T=RK2.]IQ41_QPEb>M5f^=d5&T>^fZSDR
,U<0,BXHB0,dI^/)2N[6TCACF6dT;?d?Bc8D(ZOUJ(,,]X(/O4+REE\KcaLe(1d_
G;22@M+(-2cd+0B2XOD(6L.>S/L4HABc7Sd1BWTVPRO>(P;<.U_g^NcdT?1=\4LH
F)<[@XC(U&3\B=>U,]?a[?0>0GP?(E#J8;TgP7R6@Q8e5LW,V+)8QNNF_H:(eHLE
+@3,H=V#]EZS<PT;bFT<Cf0<Q[,aI=__:3?aR-M5ReTI:cE>c5VAIaEBeESg8;<e
KO:[I78K5@-UbG>OS/,><UO6+(\#eM8@P1GA1gQ5&,ZL=eUT3#U0>Fb+3>,?J_E>
S\cL2f(1[P.7&E=TS+KB#,,>DS.]ZMYAZWKYV,c&H?^V)Fg17_V3C/M0UCd:2)>Z
3_?4N27<(Pd?7YU3OfMfa;5L>OC=02K<#FAUWFA\^473M&19]UH\;66BV@+8eG]W
=AIUGQZ_GJCGabLg/dOGdAU,5ZVX0AHHSE;7=MX?4A2PcRO:M]F)GIcX6:R1;a^+
@9V;e4I:)LYc2d,Bb_23B68O5gJ04-Q)+b(CMG4a1S;6AF6)Z(+f+@GECCD?N5Vc
cbe-A6I>;Y;EHa[f2O6U[&@LQ#e[7W&-c)]&Nbb0eE<U/WURU)Z#=Xe?OG3ga[@\
U=>DZ+<4f92\(3?f0Y?\M;H2(U4UZB=5OO&,EKBHdfeWXT@2cg-+P5cd\X_&9b.<
6D/C]MUT<WV8Q6A2AR<5#39P3+dG^&07L^2Y.OHK7C;(eNSC8cL(H,&\F+:1T.[:
6aWUPFAZ@LUM.DIb5PO=>f(-f9.M=/a,.J:Q?cM2(L4<KPWX/,TP7\+TUdA9(DG.
)QI=dJVV1COC?b9H+P2HQP[AT&C:S^E.ad(O-3<P0bD9C:PCU5>P^NQMgA_X:6Y?
YFXg5e)ORcNd318:AKFR\_d+(A28^\?>O)8PA2+26[f#OP;Z&85U;F:.Z#dV1H#5
>E=\W5M1\<-]BdUg,/9(&?eW1];OO[P::b1C4a;7LM;YgNT;O7?7bAJ3Ea+Y4+Ab
)MN\]1Be[E;:UD98FO-C0^5S3+2C#ENTWJgS0Hc@e<[/1.g,ZcecNDHf\2,8@_dg
C]X9f(f;dFYBB(1EWG><K/]]deOXdBcM>g3KLRS.WeM]G0-=II4c11AN\LLN_,d;
.fQZ5E]]1+RYa/a4?=gEa_NC?R[D_,BEXBRS,),cMBfMAQ0d=+A]V+L/AeU0@Kb/
VXNKYB.Y_4XfYY?PJ[B)EFc)L3@BF>^)KUUMQ,OIUde_0g=,C=f0H.5II+AZEW=A
2:2<A/fI@YB9X>G(feFD<daUV]W0NH5IBEGa9_eP1YU=Q1<bUBYWIOPBDEb2JE6<
bAVd<e=:>S,40K_N2QbOfX.I>E6VXG2f#d?Y,((HBa@)(5<;KCf-0WMXCOeLCHB[
1>4L5gcC/Xf_:Q8B)KT9>2H:@0?J4b^/_D6H&^d7?(O)^]aaeF2^eYDDUbHK+-1N
eC2T,G+aOZbYCf66]VOA:;V9\]a;gV8SN#K<K?Ia(Yc]4,M-\PNUNQ7L21<:F4W=
^9MM<^(WUE8:FVF<-AN5[cH)RXR9R.c6V8C8T(2>SC&[Q/\0g]I.+KcE_LXDf2BT
-3R9F-27LQAUR13\T2LU0c5_-cK?F&JK-9&YaZ8&faTQLB?G4K[#5&KXD\Z_\>J6
0O4I[-<#[\U9cf_SPG?TfN_,EL:5EJ,)PecE)R+1:0>K3bFG^Ob?=#)C4@E>1+6/
3W0)6&L+5N]dT&Qa3=:1GBfAJ3<\M.]NTRAA<TcPdQ[@E,gY+7de[0W2I4:f\X+I
/_HAc=3_=VUPeGGR9.cN:0]=QAVODG0\S9g2:F=2R=;.eK^cU9OVD\UALA_#M4Ma
30G=)JDO.U69:E,/7HZ+.L.4AYD)bJ00K?-4Q<8Sda:fG(IENV8+\/3Q_eHC&HZI
<-4TB1d2-W3SZ1+.Lg[H(&:1Cd;W)1U;aQ^AQ=VSMRY04G<_W.(_NLV?d?<4(LWe
8[c03KYXR(,c2G63Ocdc3Fa@UIYc-bZB6f4S@3DE[WF#-MbEe8JMPZ5?/e2OYBcT
daP\:aBTS5NeG\gNJ4Y9[EYQCVKV;FbIOXG(51T:9_VP#:[OJUA]U5(;dF_,\V-G
RF8V+>f3W\^\5CcK]7=\E4Q2UeKIKF-;#)ER8NJW@_KI<?-WdM1a&Q://,\24&-b
A,\Zg#7N):_Fg\WVg4aJ,97G[A>@V?J^d2CA:E&V-B=OV;@5N]GV0OXdCZeHM]+7
dVAA7,CL@aQfP@H-(2SGV)I5bET=IW#[:12VK+@KH8#aNTG,(L>2URa+.bLVg4H^
-B,Ef1O+?U.bc3J0cDc@<]V+g#D=+R\OG&M#31[O(.9)/c?fY8]T)XK8gQ2VGCI;
9?-0?C<bgQ?J?B;R?\)]3S3_S49_OQ_\fF[V\+D-GeE](LTgW]UY;61b&SX4PB5V
K3Ce+_0]#?3]#6R_>#1PJS?;>;UCH[R[W)/f5W=_LKI9-R:cL)F]#U-#Ld]BSY0F
658Q_09VCEL8SMg+GMAN7&6>a[18_g[/EB@4B75FIgB]/bHabN1G(@._&3gc,EPU
=4+B&6^Q^)ZT#,P.(CS&4a5W^+7-_]aJ];BIM3JEED1aFgVV0O7BG;Q?F9=dVGKL
W0HI0OS=K,Y+0MHU<3STR@>)\Y)#cK5)8Oa+-Ud@T,d5b/37)56W:\5a&TD;.XAX
/C)),ARd[?LC3=XaC6d<W3?PC07e)bP0##,JVJ^^RET)5e[#L=&_b_c<HBeUC&+B
\^@AIHWE4KR<7Y&^fWK4=)5/;[#;G]e:efAMbE-fE,9Y>.8<G:1XB9\+B5=6(G<X
(e-&(6NGD3V<4f.NU?DbBWeMTRV0>NUQ87g8eQ??\2^8gC4DfQJ2THXK7<_2NCP-
?689EG?5;,B7;^fOeH^NM;(((3)NHMQ/gFaVDFKOY;#:7+:aa>Y2&]W))L><fJP5
SbJgeX6Q(_[P]e3BFR+R/TIEL)_J/=3&TLcO,+N)=d>785Ab)JSNB/+X6@cc#&KP
>9B2#W;-5]OC]Y=]ZZN1Q=IU;d:X#_X1HeXB-E.gHT2LK2^KLa#]4;PaVI__R3P@
SZR/67FSJJU[C?Y<&+,W9]=#)62GGRf2]CK6bQ:--B9.?AXf:,cT+Q<I47B+Lb3K
D9WP.27-0)-G5Zb2IWD?A[3_^,&^>2&/6HYL^^.b//T3,fd1)AEQ?:6LDUC@8ML)
#-b>de.FXK[[c-Y4OgS[-Z>+:H+9Wbd2W@&F7\<+QJR5)UY]NY/(8fPRL6:(5#09
YQE^N_^=ZU.FM[H#IKaa?UA][=(E?8AP7/KOKO)F0ag@]][Sd5?/X/_08cC7F-PX
J?c<&.;Z<-cg[Pb]Y2U?eec-,Sb(U+fY:F8YN1P=)=>;43R;RWf4J)S(G=6Ag5H]
0XDY^Zd2\&G&MgAA_<OZ]Ma7J3/_62EL^@:DAQ#O_AOR.F5(C,?RMQVWWB:^2V\B
&QY(Ic;>:UJ>FLV_c0YQ,(T;:RC&Qa)L5;MP\V5WBMaH-9cDNBP-_;bW98b]D@7T
g84C<4(;.85;LVZV](gDZ>UH;Zf^<Y7A1[=L^E-bB7;+#3OaLD^AW?(-Y0RDNfR;
F>aYC,P0F9920+:XYK^a^XA+YB9U1)4bD<N:TDBTdN=O:>JcPX5g:4Q@W7H]#FX&
TOMObTXSR1HN]d[&X&cNS@7_:bO_^Q/F^:-@PZ]^U__R?Dc.&3(LJ<SGX\b25eO=
>1[c&g;Y60MKC7&OG>E8f+Kc5U)g;gZ^4P[N;Z@<Lg\R=_0&0XBM8AQ<I>M8;+Da
BYX0BX_LfT@GEX6)7a/D]);+B^9&>PBdPWGTW3_4:Fa>QQD]Ka#0RHL/#_E8-fS?
0X&d;1D5g1>1fd69e38@N?X/SNUD>,&3@U.d1WD)fVV._XH91YM)0SI/2((_03/I
TNK=)GQTPgYLULVBJQK=O+a:CdVO3WU;4WMNLZbALd_=Vf]:Y)SL5_ZQfLJg_J@S
33)GU@TUfY-f3I&PX=[\GSf2?,XF4O#^Gd#@S&b5SfaQQ5P1W._U)CA[I3Q=T2U:
Q6OVe/UId<FN1G+a,WdA:)H10FCYT;gM?EPc_-c^Ce/6O0Kc&N(25f[V]I1#[):L
=IgaXDOcg;gW8MFa-A346R5CcTB>b(LO[.5Y#N532&6Q,@H+bHW-c(+d7&YHB)\^
M_?G)0FQ^H)0X44VU_\1@Y_<a<FQ>8^EE0IIEI921+BZ]?./J+R>8\)7\NFW.B9e
UNF5:@_d]X;LcC#EOf5I3<B->SM+3#bgDF:,9;P\+.[YB?^Eca?U3fb7X?1DSLcF
W/KHW,XV@=X^X8V-f^:/RdcKKHG],S0-6gX]#R>^f6@/HR@4)&4fU\&cXgS;2,YO
bQDed6FLVK/QB6C<)c.(?BYLMIX@1(&V.7QM:WP4+LF0Hd<SFK,)-/KI5gS.4_<@
-HU8>cZLB;Q1J6#7c?FDYFBa62M6OQ;RaN]1<GM:=GUaY^71KgG6/QUJZ3=a9JM0
^.7;<DY,:CU4CCH]A+;<d1JdVgbb(J?NTM/I<#2aA,UAV0_(WfH9#IHN:^25=cSL
\-:F8HF^J5J:Z&RB_ZB;B;3^b3U9g\\VbES#&/a0CVBeK[Q#UT8Zfe4cgQb/)9bK
D<J=/W[P3NfHV371WANMLZ1gP\4H[YNKH&01BIb7ZZPRT#MGP]<T2QB=Mb;Z8V_=
#K1:-?V1ZWO^,1-E?YQDHQPe,I.6Z45D5#O288dHe=f=,V]Pa7C,LfU3<cG.QPGG
8FOFF[45[1]N<;0OW#cFVgFF=T25<X,dDZY=9R>[C52Z=XF:]-8I(/5:I-9C;V3M
+[9TgL;-8_@,R&\0HQ::bP5OE17d]3BOCV@OPWe5-2g8&cDN+JEKYe?>RRC6K1DI
J#OE@(MJ\dX>0S\L7Y+3?CZ)(,H@>R,MRB]_5YP+X\\4dTCEN\?cY.e.L=82R\K5
]H7^5G;GG\FYLaOB\G1&3KcWN;ES?7+DFG3+dC(7_L[L1bdBA-)gH6/@E7Qc_?&b
eATD&+X^K:?4#N>?^Ec>D-ZQKJfEZ-[,dJ.]ScOO(a._RG^@J_Ld+H^E6?\d1O^>
^B&P,U8+A5:0-D-64S1cX-d,4\LDLaG&RVW:S</ZN/HI+TATbO]UC2D5KH]3#3X?
OCP-Bf,N&e<eOA]S8W0b=GNgJdT(F6R-M#IYW]>3<NXW\D0]_cZ+ecbFA&B3>DfP
S5=W]F^H.+Za9We5@cTN0KMbf3\F2Q;\RM_JIa7(??6&89/2H1ZCZTeQ)Y9LH_B_
I+2C5LP2MTLJV#MBb#VMG2<?Vf:MA_.\QS?(<OKUR;AZY4U[(-WYMbL4F(?__?UY
b=WTVXWRQ6BYe]L:GTTD3#V.)V^@)#]R\-Q)Tc=)Ba>1#4f0[+^FQM+0P@f&F0N,
#9acIgCZ(]N)c1b8ZDNR2aK3GcQJE>;[^fJ>J6#32;?=#U?8g16LE_LHWN0;.d9b
4)OeMFUfCPI.CWRR,B-]L_09GaV7>-@-OAG(,SN^TOY3.3T2SBcHWKb-93<WWMb[
EQ)520NDW2L9L]290=Ob25^O6a?LZ?UW3.cFAUg61&&DHG[UYG6cZ0/?X_#HVU?+
Cb\NOJgD5S62X>M,:;;a-;aQd,5-(=GZ9TD^.EAUCNIBX3-)XcZRdXQI,:XYJB_&
1Z[[S1)J/^O;fQ1\DbU+RG]5M,,@22K9IG;+E]>Ka26QRYXC.NbF1C2_)b2Da+U@
U)#BN9:BCQ^SdA:EaUPV+(XZ7&I?)JI1Y<DeGV0bcK9652C[(RBAH7;:84]L15d2
(?BC,S8]Vd,EM]9G7YL_S[9=1@[2PJ@U3_FOEKaIC,]AK#AdbWa;II#]GaaDJg?a
aSa:W5\23&OF]M_J.cZSY8QIEL0MCFSL;4b:>=A(d=[<e/P]XUF4d0[+O5/8&d[=
eF#0a\;5.NT:)<?;_Y\Wa7.#@f8S-RM4<_31M8=6>Ef9H3CBPbZQ.LB=?88^K:Gf
-K3IT5B?)aEWXb)QY>-Y.?FA<<-SK=f97_(e(.M)&g0QD2d7?JY?3M\Qb=YBI&[S
:T8SF826CNfS+3+aUe/VODW0+JGXJ@U4E2Eb;9aS\<J5.;_G+9Z#&62=V]BF+0I#
=USe6TGI)=;&XEf&2ZIG9OM39;>d_/V6<HFQ7M8Be&UX#L+fV=^R&3_T&7Z>6E0<
KR_e)9>=JL-6T7B@BMa^]+(Q?.X@KRFaN;S;@+d8=/f@AQR4GG(23H?3#6U^)=_1
0A]c]MO4bH]UU8B&Z_;=:I)\/1K?L<(fO5MEZE4A&:AdB/]Z#H;CGb^1/JD-+cIB
D^2ZWY]L,ND+H_E^=RJ0Va+J6gL>U/XAdZ]D1>=Vc]4>dS9>@b/R:g>_;^XBCeH6
K;NK(c)97E:O(Z5?bPY];V(E7Lf6M>L\+X(++51+4H(M63;,YEOO0KIG>DE4RFB=
-/VJ62&1Y#&M?1[,)X@4>c&YKWgdS8\SW^d4O+<IW)KV5Z]U=F4Q5B@(WDE^/\17
/Rf(#EX_EKLHWdQ<.R3+VAK,:PFXW6H(6X,D>XW[9J4g2(18T9LcRIRQ;Q]gH_(U
DM(#TMY^^1BI;K3M4Pf-bOT1V\V5UUCCQe@Cb@P[N7+L>1B-\1&(KNC<]PbUL&P=
]+(,)])0[+:D:]DJ#b/&0I+#V7\F<XU/Z/^YS2CD6;C6B4(&6:A;76)D-77cO4M_
UO67#&V;R1ZKgagIc:O;R9S@I69(IdD>7NdUbC(C4-)_?<Lb&KPdB^@(&O1V/gZ7
VF4B>3-HPM9=(J]B8gYg_c]S2W=UZ[.]GfT52:3#U9RU29V_;6#4O]WC;HcY_9^:
[S87Qb,P;<EHD0:B_5DSH2=Z26XS(FV6Vf#@Tc^NXg+X^3V9EZFWP?LL&EbgQ3BW
]f:D1)\6=VF5J0G52#bES#B#TVUM=_[3/a&KUd0eM,H@=QV8]X&GL<7B,;g3PV]G
bfMI+8T65\_;e=7#=g+C_I]:d@a79[?L5=(Jg++,.aD4;<WRWd+F:a?(F[Q((?d\
f6RX]H[dPM25Lc#UJ/P.:O[e[.ZC/\WE[NA&TU>;,.G@[?&0>bGN>>.JbEIE#AV&
)2Y5Gf+Ng(.e0Q>F=L5c/E.5g4(L5_eD3T7K=S6])ZB6:T:XW_YeHa)5a=caeG\[
XeGDU:?Q31X;1;GP6B5]M3EO0,OKRC5+++3>P)3c4S;+ES:I?E::5=CM07/H+^6K
9Xae,eMFL?(=A/AE&VW/d8be9+g^a_-_,d:C_07Z&dN_V,7X2J6GVL31P8LDHTC#
,_(FUa-;&[e2(e8a#f55KJIJN2N^+-/)VIIM9E,8)P4gZTEB?-Cd]L&QCOMO5e_>
5X2E.^U?&N>H[cEgbfa@H<]C^CM@/RW8R<+SEQbB9cBSA/M?SE1A910ZeRafc@BW
H/Xe\4^FK0>cd<QA&0JbP8K^N<@&_Y;USYHWP?EEM/YO-T/LGVL>XaOa(;0ZA><Q
9)5A#+KBF,.MI#H^M^2d^=W-+\GAg8#DE+BF/QR_L=(Ed.TaI(OcW3OGT8.XD=HG
30NRWSJ5GN9@4X/K6f^K4]3\5a4.R_:0M-PICAf8Za383-DI:cF8e?4a)=]Pe;#0
3&]A-UcCUYOeaS,>g)&ecX1MXERG=NC>E&dT7Sb&SCVPJKa[?BE_X7H?03aZHF.T
R:/fJM1Q9S2/e+^Ga0C?^MaWB)YU?S^1AdRNR;;Q^VF4gYLO.5[H>+JI0L;<?+WH
\X]bQF\4R5fX7U[U<4W@>.=2T=6FC?-<8DMg-gAJ>.L^Ofc2(PILPIUCF&,Eb&fB
BX50eS(E\#RE;PFKLI46#]K<&(d&acMCET:8N>e9S1:KB):cT]08JF67&aga>H5&
R2TV^?M2<8]IW01eZI,fL[):G0IG__38EB2X-X#+AS7N;#SR(YZOP#_^H&<P)<M5
.ZXV(:A;HP[e[6Q8@\e,FHTb7cMVdR9:](GK.D#M;O.X9T5OQ6AeFYg-,8LTfERZ
?/gES#O=,120V<ILCa=OLY-FU5XCJ&BZb@BGC<abJ:(fPFHD=9#](<@N5d,M-((T
A?-Y52Of_^X1[LK4L-fde\YM.S53AX##-D-NCRW)YT5Ef:3][[P018EAP&?7fA&\
Bb//J=7=S?XCA8<8a=RQFbUF#B+d^KQXf9E=<-\MW-Ke3&d?#F)X:K(g,c2J0E/M
0C74bg15SU48dEZ?Y77#T11@SR+c-)-.QR344PFQTCS,&S;(Z6#O1MM)X_([/=QW
eHG[&_OM\RF]P_CI\K&3HWP:)C-MP>b8B@R8^R05HYQ]\(D+]N:=-73:W:+LR_DO
@1:F0?)\S&:VED85FgQbaOc;7[@(^[X4X40D]>e1]<U^bde3/ZXAN1ZOEDa1fPVN
5(5>N\L202Z64\J&MZE7P(#gL]=(VQJSLf.>S<T9g0FXZ[0ZJ[>O#7N9d7SGK:eO
2DgBNXY(Q_TUb.W35-2Q8fNVIIa(4;dA1R\e3R<5:(/G9[JeBd)--L]_&1XZeWLd
-.JQI(M;-M)_F@>U7+Tc_2/,WHA[KW]N:A4GT)#=D\Z6>g(4T5bQeQI;,+(eAWL7
Kg^,78L/:,9F)eYb1S@T^a9.L=ZDd>,GbMGN-TAMb+/Y4[EQ6JRLGV=9#7X7>5T)
BV6.F^56dJ-=Z_fYMQCA?aTY3@0K]OKJS53T);;]VJg;]7>(YaTGY],?D]BT0LMR
;gdd&TE+]=[XU.7>-XY[[<5X/2UMFd/GNc?&V\LX>e&F&1-6E@P)MBM\.+(=EXcF
VN.V3DgXYFU+50<0W@]G;LPX4N@T^F>HB18-e_OW@b__KdLMI+#e_ZQAI]X[LBD8
;+<\4/AE>@#8H/cd:)L.XA7g<Wd<90VC2.d>U(DaYa8A&>9];UO3b;K;EJ/MXE^^
4D@Q+.7V/V6O]ScQC[_E/6LJV-JT0<F(eF;g8._,J(_B,eHT(IL1Ef\<V^7>\/H&
7:4fF=?ZJF.c(Na;D<:SQ+7._U2FK<73>:d\2EM4((^J\&QJ/M)BD==1Qg;N]dEV
GGb0P,AdQOO1L4e8+>0F\49XVM3F0eT-1AE+;Ybf/QgI\;>__@D#SdNd:T+-4)::
:3N,b?UTeP,Yf5AbN:6@Z<F,\4^DS?CdgL213e?K);7,\a;/@X-GD#b-1?4@c?c2
BP5QYZIf+MI<4Q>2Q_Y@QaISVGL59AeV6+CF@:<FQ)_+RIUOU(6dSZ3JCCM9>NdJ
2F-23Nc/WS0:#91U>fLXYU=gFcL7.:46.L^A]ZD+D91g<XEf5T6e((/\#=H>Q/+F
eQ8MJ2,=c>6EUWYf>&:@AEM5UQ84KXY,NS#d1&X3AXfKQ);>dSTR-)eNA4<:AC.A
F5VE;DNOcFYMT+U7EdE1?#,#64ICEF2FcIRLRg/7?NE>0S94_XWVJ^[ROO>-PKU?
g-0K.SB@1McLX1()7&SL0UD87d,0#CSe=G&(g(VH4XI@]L<0cdE<+</&Udg9Z9.-
CcK\\;,Z7gYb[2,9G\VOG8G1?eb\ZR3-YFPKIeeCT:L.5ZNKO+EJ8<4#Ic9c<M.b
;\c1(3..=_cEPeW^PZ/bANIQaE(9d(.F5NN_1M^5V)JQN[M.&54L&20\eX[gD8&J
cQ,5cOe^F)f)I1I1Q9I(]6>bDba8XVCf,A,P/W5>U26JE\Jb)OHPGZU,Bb-b8.4P
6a&I-A+7AH\L8E-0QJ,(Xe7PYPJD6KeQK#:P:-1O7JYE+f5TL;]GY.Y7a=MAZD(G
_:,@[O7[?64(O1IZ\A9+X;,QOQ.D(PBO9L=OP<X(SX,We1,]DMbAI2:#C,L3a9>G
GF6X&/M&>d?9J^[)fZJf^Y3)\Z8)4[[+4@M?@@Qd41BZ^5IKB6ZG._Y1MbPc#g3]
>S?8[BPB4ZKfM40Zab47YR_NQ@>]<+<CM9FRdPK@dRdEHCAYGHd/gP>G7c0-_=6\
SZT/<4/:_B&8WDBPK.@WD.VJAIefF81:Z>TUL2MWV(194=.5gI[Y)V<0fd0994(M
GGEQ5B6QUT\cA41DP5c;J79(M(e/G5O,AU9R[#\TG84,MAaAQQ2EP7WT\)O&01._
(+F71K(<A2P1&N-@=W\#GE1R]9)I@U+NXd(I6S+1R@EF/SI0\8GIc>bV,c7]OD-Z
1[e0b0,-GfJdce#5B<#:_DbA7P+Q\V+a>I<+b[I]8Ne5KHaVd/N8RD?3:6#ad]JG
JZEeW7-cE(/],Y.&O-b]egZ^9<H==W&0#7?):e@M9.>(GC42_)&JD.M&L-XH;E>J
IS]]M&(7U7(DY2c;ZeW?8)((e>]9BCT4L4(<5S18CNg2-1cX:-+??87^7BH66L5-
PfXJ:-W)>WZSO:6YYMN=-b.;WCN#cDASM)g&HT=HEZ^=HL2B;<OS/;FKO3IaL[@R
N1VYeJ#63I<YZ+9;3a:M^7dJKc+f^19::VJJeSA=(+(6G(eD)Od2/YV2Z:5>MaL6
PB5-+:1NV=]:f3>ALZN0+L8Fag7J,@]_^eePU_JVTXEQ3#\[JO^(4NA4C-DB.=#^
g]Ra1a2;gNf\IXTLE-4@cGA(V/6W(-EKXMR/e#U)9IJ7^Qeb=f=5Z<0FMGO)6>>>
6M,fDeA5P]G=H&9]WG@@GFKU]?GPeIK-.7gP?0c&ANcBWVAPZ7OS&cNJ2N2NLa_&
aJdVb8Oa6OH-I_MW5:;]0-_A=dfPQ)?T1\2Pa<F4\=VL_6ZQKSa?:&B<\2#3_3R[
]XYIYUH@MFXb#[d[+E<TRdcB#NdCTLb_]H3VXQ758f2(4<.NDQ2c(aXc@&e<B6bX
:MaO]Y<S9_JYRE4LKZ;S9=?.KAcddJIc@W^6&U1D4N8c-@^459AWa<fNe15:f]LT
S4-dN:?d7Z=/#,b#4[#/^Q7KV8/.GG[&NYA,;:VK-)CGMQ5V,^9(a7[:9<XI]PD8
W=S<.Xf9NaO<E<Q69OSSRfGJ=0-U1LFZWf,cV-=7F:VM:C@<AZ=f)2Oca[d[I<4<
,A&A])7P?\3:LN;abT98d[CT7[:7?K?U_(SGb<)3>CS&A7A&URMBE__<4)_7WIU^
fI-X7=3NWE(P#CWX+XfX=_58Z]-PFe5c-&P<a9VO9]I/75?<LP50XC1\O9R)N@<e
RBV05L.[0::O<aZBP,U9NW(.,eK<OL#1Q(A<M_DWNC/UTfOVSe&U(L+__bY<#M0N
CKEaYQ.><JZ(HCP(:96=A^T\/;I?:?U3/R7=1H3<gTJNGUg276)/.445[/I&.T.:
.O9edg:g)10</&.(_SfIG=A1G:O=fRJIOU(H2RC1\BY9DF3:DcY&+8G5M+WUcd)F
:J]5O1FUKQ.M,DVG:^&/BE.+NWg-Ef@<6g+6X32UVB_JE[\d7DI?0G^S?DY_I_>D
gN.FeXOPQ<a/c;14[D)Fa/TfKKN45\-JW.Z-Dga5-KZ6J#8d./9#?HVc,Z18MS1b
II?^)4\&9@D/:ANF3JX-34b3^:-^T#>&O[e0BBfF08_#=>Ac;Q_FAE5_9V<HbME;
YS7)T@,,aA9f&fTQ(aLK2QI\W>#C_cSdgLHULe[G-GTHO_P#aAbNWGROS)Ff?f^R
H^L&N6QP@b,4c7PcH+ZC>BJ=I#BUeMC7&0B9(#VB>M>3GVc7=KD)W<RH0&7@G89X
@.eOF=[=9[)Y[8f?31?be-Q5I_R0cH?Cg=M:CE:<g[M^W?<#YVL:FN#D6XcM74Y:
\>4Q3@g.Z,3M;>G#-\(4UF>Aa73VC<)FNd,5X1./]&(F?>?gWd.+@&/-IT.^Z:b2
UA+(O?Z)P^Lf5^)KJQE7H[777D>7I+:;^2g=?W0Q:Q^.9U76^8PK>)[#Z#6B50Ib
@U-LIGJg6d#dG<U,f>MeSf>\\I5]U2BC4:A[SZd+B#eA)e7K-OCSQfH8F4bMETZ8
R+5g70V:[:.)WHU(aNcO>>_K.F88@EG=:+J_MN;YeDVdM(\\W)U6B2)W3@.+M#JH
^+O@EY#XNM)3Y1NT6_3-(R:,G66eTY,.ZI?\[VcGb1+.=(S+BCE\Ie.L20UEa)PB
=Y\CTTWMC)\aP2ICK\W11^2@GO7Kd^IS7M?(^[N&D6#CTee/SU,gS]KaAeERDP,]
-Se,X[G?,=TDTaY9C)eE7VPU,Y[:_C^X07MRJ>cQGD2/)=AcR6:LP-e3[/EMPJ12
XZ]&WZNB\Yc7A[8c+^d/P&=G1FSYb+I+WUg1/==U-f;QF0@F-.+fb/F]+BDZb.AN
A]WOb^2:=#+B##W?C//SPK[OK6HIV(0I+-dCJQ(9F@)eedbfc\<.G=0/C<]IL2N9
TUSeD)X^/1)fUC=ATLac2QNMY,c#MQa^JS;)=a3-08PNT&-.KUZZV1[ONF>AVg,)
>5cICT53#;3PR<Mdg+^>09JVg5:2g&8OTb@+7bbE:)QMF0J@ccDd2I+a:U5E[cRS
@JIf,L^OHLbM/->d88c0Y<ANEK2[#5829L4fCU_=FYbC#c6]5R(0YaXfT]0C,PR^
KP/K^:4Md6C0VO-Qg]L6AZeD;f.3[:P-:/M^[cBJ35,HGH@YDQFb;_1#K6NESg?;
ICVIDOWBJ>E9Z^(WD&/Z;B]:F\7ZRCdEaQAKA]Q-[QAAA^P+=3KeL7,a@Zf>cOg;
>d^e-L,1&dZF4c_8GHM67d4VZ>G0FUWfX3D7?aH8QaZL#J3>T>>P/]Ud[2P1C<0K
+S/gbO]DX@RTd4d#R+3#\8b4<QZSWK\##HXW0@O12G1fJf^KTVXe<SY4d5L#DTY\
M@[3BCfcVU.OAN@bQ=6]\d.0M&53<]f9;)_eW+[S04J#b]YI/BJ/eO.Dg8\[8F1Q
\dQ;,f.8DPQ&)/KY)=V^101VOH+geI_H17#X1Z^L[Q4=^1Y,ACVK<6@5=cMTSe;&
bd(^,<NTS3f\?OT>^C_@OED2X:+,PQ#0J)94=&\eD/NI:f4/3JD[06fLa3U+UB.F
29>9/MRF<A(UA=QWVE5LWe;3\Y/eYN(bHS>3NfGY_>P\S-5F4eY7cJeRA3>aMXB:
0[eRM[=dUd92(\S,W2MdAI/A]+geQG24M#/0aCe;?->V#=b&2Vd&GU,D5E9)OCVL
6AL9LD_?ee9#bHOMX,8WFBG2gD#Ng(CbcT_VWaTTObJ\cJ,AeNWRaE3g\_\V<+CW
a\,1[:Ug)[KId=XCd9>G[PN?3Y?b&_IKW\6@1:]2V4f3JP6QFd[,0Y9]a=^#<fXB
X1QP5Zf1V93@+U\_0f;WC]5+GT+S=PLK#)5M7#[B7]E8(ZQNVW@Qf4DF0V),7=?G
c]Rd7[3NCe5+P1#?\KP])@);ca.)3g4R/YBB]\/<8_Jfe\65)P8R@dM]d;e16(?S
PL@D?4^9HIKBDb(B&8L#XCA/2d[2EN:e&Bbce7&b=(QE.F,BEd9MY>&?1(=^QVTJ
V9OdJ<7LKYRJ0H@H.N@G?B@LTD2,X5+BZ706&=J:L\#O8,Id/K8?=?CN[4]7@gKQ
X=[S/QKegOTT-=DT&]:Q]Ba7Z^B5R#N^RD&]fJ,GKDAg-L-TEJ723]=DT0+M?-U1
+(203\SZ8^JZ45BH6FUc;M9\>W5=[Q\6P#E_LL8-?:1K0:0Uc9\[T0K-a/c3N#_#
WCD[c>#bO(2ZLcV65CS;P)[da-G0MJACD<9309]JfCaZ4)L=P^cCYP._)[3;>.[/
XI1]117JD.:M:C.G4g5f^4H-JICLKe/H)aI-MF4O<4]WE;.IeEB:@eT4FfCe#4CP
D@(2MdE3&1WE+Q\/1N3P6+BLXRLaJce[>Z)E5,E;.f1CZV<[,?EeX,5_1BD]@KO;
YQ:(Y?:O5db2;XU>b8]T0=R+>bW6,:_B.^PNCSfFTM#W4>JcHgPH63+-ORES8HgP
f0[(OM+1DR;Za(^[KUVZJ>WcdHgK52WN\->ILQ=gfL@e8aW^@a8=4^HN:Y8eMec)
0.5.>/A.TLbM3G3&Y<7eSEE<.&:MMQIc[]GO=Ma=99P=d+e;>2D0Q^E4/:[:FE/Y
]PUdgB05_eT7eWE9H2fLEB<#SZ8G<WZg6M[K)6C1924B7Y-&Og3-ZGe6DPB[1T@I
\^><Xb2;DPQ0ED&5E/)I>:YOa-b8c0FSTYb7HMf3>+\eL<.RK.DO>c>Aa37f-8DX
K7PA)R(XW9aDNIg:,#8JaW5gW2Sa\5aA78a)GCE/KK89/#YK,#]-PNT0.NKZ_+fG
f62@/:#1b,)E4geCVDV/W7;a,&67P3RGO@7^;>.6JfQ8?=XB&a4L(bFIB;XIb5,H
=cdRd6dB.]b0S,MF]X56#)W/POfS4d;W2]Td^U4Z[OVbD\6_B7K],e7-Qd&X#,TB
IM7e#]L=S/[gF_@&?7PMXV(bg;4>;f2#EIc:IUX_GA(CDER2bg.3U/T0HcX(;W?>
PEK:F-+[U=f8,2+<?2DZPKNMVPK>c(?:fT1C#9BeDV+<Lc?N\aC1-5;53H3:Lf8C
XYJcO5gS=M;90DD.bMb^fXPe^V:5)EQ)TdGJCL37Nc;.Td/bA>d/I8YDI_L_N\.>
\d[:;+ZZ@Rgb0MD\PfN,31OJK0cEe^HQY=SVN[#N=D4+Cfe[1d+X(\5FN4]Gde^)
E/E^VU1+<Vb9f=?eGddK93/P#F@^JZ/5UP4-;#C\[PdRYKAWF_R_Udg@LT7.1@GO
T#9.HY&PgOQJ7Oa2CK#/;0+:XCHgI,aL0E3^Ud;PCcf?+ea61bPff;aV1&@a-1YZ
@FT5D,&8<5d-3>1GM>N:6,:8/B+DZ>Ib>FCK<VcEY(.W0PT\2#caZ/^8e8RYCHX.
4fJIT_HLM[3dI&?7df1:G#2037L/>KA/@68\H[&O9//Ie3Xf@<3e,,<T4;^<QcI3
a=0HB_W#9Q&KNZRVN+>>dIA>+0JaAX,DV?-M2f@eDOT-?Ebb1]+AB/(Lc4YFBB1N
b1F7QI=5F9N=YKMD+?,A]=;NNB,S(X\/[R>YFH57I#:K#9)]6ENUBf8^#JA.<MEd
@XcO>28=Y.5.G9^MbQL(>UYYYIbQ=99\a6K-5[Q>F,BNUN:5c(c;KXHa\IW:\=VU
/>4.2Idda)3X8FHQG>7]07Wc##X=W?O;R^(=C9\cPR6+\3=FfX&Ic0e8<S^2(2OY
H6bD]-O6\/4,c.]fZ&^eBN=4;MYZ^M7eNbdG]fb]TI4EZ:=KSf[La;5B>:@JU8>A
-;2/+S/6(b95@6ePW(=TJ8HXH;A5@-7[DG:+/bRK5;^=77g(_5Xg<gb>UH12ZO4d
)/[1cV_(FC(G>@-91PZXgCR\WP>[/4H6N#<F,?K0GUdM#3(dW6=40a8+[R[fT]V5
<,1>Q[R>?5KA2.4BfRd[V64THQO=:4P^Y@5+;HO/XYT#_EDZUQ8)::R6)^]:cHGR
)^^^e>_+2W\X:14P2TFUYMP.)]P16Q[HF6L?f>&;.(X\CKMQB0S]9<EJaRBX8>A0
OGKSGZPX)5O9UP-KM7=(N10+GWUQ6=H=W23fG>U/fdf#JA?+;K>,f4-D--N7&S(#
([7P&bV^)H:5dLZd6\1M-3MFX_#b[4Z.TUZK:#1RU/ZD71R7e9CQ0KH0UARX3RES
(QfDJ^g0S_>gQO#[(CHJ(DIVf,V4=DaAR70QLPRfF:eGKJ[HWQ[LTM4G)/DQQgY1
\32A8SR1#&#7PB(60[\?aQ]\SI/@KAPQ>gJ[:5HBdB^aY\a+-MMf/.T.62cgS^cJ
1AUF8<]F3Q8&a2MY#M=M]IBe2cb:A?c:G7N>-,>VQ?5,,>e-O^d74#]E:dR)3g;S
1eE[,]14_5886SX+VfZNLO&=Ld<d\\S(PLL.YM^-aF>@&<YT(&0?L6KScOJQ?(3>
\6ZdIG>SY/W(.T60U5:RDFX:-<Cd4U,623G;X]a=c<PdL>Sd)?&Jg:+Q5E-1/I5<
K4^,SLQ2aC5HU^OGTT3@;3S6G=>R9K.&cLHK:JQbMa>RAPFZ\+:dS:..7<:/1@=@
8?gBE/b^,;;5M6@&e5&OI;EUF.NR\b)38D-4GE-.g<C79]J;@M0,ZM>).>0e&1TY
<G63Q=?4f#T2P>FXe[@_@#?c9A.7X@:HVPSB;JY#S0KWZg=]0S:7b;];8QcH_I5U
O&:;XNI+>6gg)OZ:aPQ-/]9f66@]I;cXM__O2ARYX>OX]:4S76c]#+;?)=H\U.31
Q/^BU&OLBY8C(J/Z1aP&=T7-E7<OY.85.6;4eNL5G/6RL[]?L7]/LC.AdZ;:3If+
e?B(?d99:],_DLZK2S]/E)YaHI>]^CRAY0L&,(=UB[3@#B.CHX2ZBRe?[DJO58fG
);dc^gf3W1[MJ?L-G<ID\e3GAMES9aL;8e/T(Y.YG6O+Hc/9cX[@3TIH)-E(+R[^
]B=[Ed,<7d20X5g7MDU_V<D@VEbPAC4\0,-W1?_3&BM];U;=G@Sd;>V[fUDW\R&M
Y\\D,L,VI-C)L#dU#BD.@O,cIP(];JfG7OSSX\:2<8ZRELb1I<5Lb?P6bAWG^>(D
G/HbATV^+HAU_,I&B7D/FQBPRcYGB.ba>@cW@-YO]>?V/N-/V/YfBe7>Q,FI_Pg=
RUIGJHeZV(XL-P,P+B^Y^;+4RC&g(AC;QgNG1]]REJOI2Uae?29-3fV(DF[^R\@O
/ZLV&b:F]WDFQ;@Aa@H2-6G^fYf=4SBT0CSFDO[d-<a;29VDDG-.L9d-If11/JBL
fGWgQ7KIJWFOU0^F,;RJMb\I4,-N.ESHU8VC>Y0af2^,1VXNI@#?3Me6gdd>?[17
ce4fDI^:\0OaKE0Rd5b-.Q^QU#e\1[(B]93NHE9FL,ITe?VUHMAc,LcV4P7B@-c;
Wb][&P92E:J02]AYBUBFF6D5aYL0YNM2VMW<:[UeERCR]Q1JZ&N82UC?f=#gV8fP
H\&-Oa]FWG=7-O5,O)G@I_Z;4T)UZXW)J<QVUVgKZ3T^QS-Q(U.2EXe:eRR1g6/\
.4H^JgeN8@3#?>E.8DT<0SSL-]P0WdDeUBMW?U/^^:H>1A(#P5;QMc#2-K?=><d(
gDP6T[T0dF=5]7[Z_b/KYY1.#-7LJd7Q3gH]C+.U8^NdNf9P0QN&02TYGg=cU\@M
8aRP9cSEQc71U?cO21dQC-L.feEN;Zg)<QF?\NfIH^MB=3GM/)5)CD,0=#U/[Xg:
8KBdA6EON9ROeD2ZgHe[A4POX^1X,C;,)XE6Zc6V&f5I3bMJYTc]Ee5B<V>1:&PP
O/-^#_B;JdI757Sd[f15VZHFdfXT26N:#@.R;T@baPPXdAeOFGa^-EO[/g8CT42R
4ZXc&bNA?)MIUWF5Nc_e<6^N^]8JCT9J:/AE?7;/TDf(40RW^A]0N8V+.(+->gK5
@J9NA<-fS)PHJ+4I<\--HJg<7e@_+_-AFEJ46P-Sd..=865VdTR5[#)4?A5@SYDL
1B-Oc[7P]C93X:ZC-8.?,-[F;H+ZI;SK-1HdO=YK;^X;/[EO@ARSD\W&>88I4AFZ
VP0?>Mf_+>.O537>CJ(J6N7-VMWNMd2ZNVANRIYWW6AY[=>aPIVXSW(YM<VO=.E:
?f39e/KM,O-9B,(8E3Z[LTF+=4]9bDSRGg2_fJ;D)?:P.-IXb<7-7V)6:5Lg5TL5
Cd^MCPbM01f&7WQ8c;Z+)/BP/2O:f+8fT&XN+,TO\IAX?W=TS>J,9&3R+#[c.@-@
+7=-6ZZAR6,84>CNdJe:DARB#&YGb7GJE/I>?NKNE8C<@EQX7OPRf+D,7Cc=,==/
Y3].VUZM-T_BN27,=RUQ4L[9e05J\Z[P?X\;>GAbAX@L6P8_9\1Ld7[b+?)W(\JA
/AH31_&#QPN<>BT][)Y0^D)<+4V5FO>T@.1R&(P0<:?H;>#)feSbORfS=<5_YUX3
_N.2;Uc=B)C5+D@<>E>e[,R&M).IA\TCS)(\2R[K\9BMgE@&QK,ReOaTXATR.@PE
NU2RQ],HP^WGXfgGV#-QbYcNP+D8&XX.Q?dS/9U<PU-=(<@eYLT(,&aPd@Uf5)U/
bXJ]YT#8AXQZf0dT?O&7P_B@>@M@9(4S6bX/5a<gL4<(2U<2,9/(==J5^L)1\-2I
@W_X5K0<1MZHEgg>.L=.d[;)Z460^A7dVF))4g@3Cc:W)M6fEV@3+Gf;X[1O\/]&
S]GJZK]SSZ74__D@TJ=E+.V51a)^^1CJWG43N/.^#)dG((FYeVB6T2#D3:H?TfE#
;=_@I#N-]Ba<4YePePLg@&/@Le=C<_Y)dY3U\BEfA4U-20<YCY5SOQ@:36[c<0Hg
0)X?\VgFD5C?]?L+F+7QRZNCHT/EH@ICbeC)57])+O_b)/ETB,649T(.g?:W.Zf[
W&;g2IB2:TVBN./\HL34DAY?0]7F5#;H2Ud=:D(O\/HQ/@Na=eJ=;^HB38>?H#D0
9fQ]ZHaFM:+[=OH<BJZC\Y@UB;\4cB\EJX?L8]9QCDTB?+>@Tg\#c=b=0ICV4R48
Of#K]U5D]M#S][R=d7A6N>1,#1&;a>?dPZ2#.?G7aFgWeKI?)[92)W[&6:,K3?9[
8eTfNc.1LVH\cW3aV0e1B]<S@K@KS)ePVEY(]=cB_aEYOQ<X+-a;SO:::=L3KM31
7TUT8ON+U;</TG^6H>W^#HI:5&=[2D<=WRQW&c2K?Q4[+0abcD\&+V3L2=bW+cVM
DSZ21Z9Z=VIaO=VK]NIMCX,^CDNZ2@U3?d=38fOWRMBBe</L@GK2^9JHHWY]ZCfc
N;P:S6L5_6J0eZFc)Ab2d<7aWN6ZgLfc83HT?6E[1f0](aD3&b?#d.cA(6^7dB@6
I>VG21b7fQ311_:V8f;AW4O@.7)/@ddX,1I8M/.b>=OYg2BK^SNI,WK?P?2Z<7XH
SF4<5]475TRfGO6:fcF\/E()Vec+P_>#3JX0IQ4_>?51@8bY_X78Cc+D@c#/+E3]
3.@6V)S?N<?KbfS5S2>#.6eR8.+M@7U3OZdNHRXI;2Kc-&)8/Z&.O,ESb6&(BN#[
6X4^bU&H9=367?g&:&>Mg+C1VOKQN2?8?X;\1C_.89b/-::DALBb&2YLYF-)4W<W
gEaMG-?^=\Q2#6YQcJ:3e#G)@2-J9KM01JWJ]JG)Ig2AeSf@F_c-B<V\(FBfBX.+
+RGY=e@SDge#O&J6M(e;J/=)@>fL[NE8U##+f];cW3\G^6-7]0<Qf#aT[I:[B[g?
[,#/Y[[eT-0[EdM7ePTR7G>bJ1CJ3-\\\]@b@5TCXGXAB_=fd7cZ4XHP99U#X2-/
=27AHA8g_FRE^8-.O08P&)JBYYXD724S=50QKEFTL9;+REHQU/@7D)ceQSDI+L7d
1Pb?#R9//CP64#NI8A]\C(9=bUcP@f0+6C?^SH/cZ9S]?HHY6\V1:7RebTX(RO/6
\XK.8/\]/O-KdR4aEJ;)?>9Xf//gJ7,BEI,@1J,S@9P;^D=JCNgJ6:I\8M#_.+8g
PJgLFG\YMUff&^KIE\?fL.OO_e3ab,5gc>dO#5Q9;/U@KLUZ;95B:cL)K3=eU\bZ
d9dP3::BeSU:CF04\Yf8;HI^#5?1:2]Y@+3>)GQ)2eC_b+Y2]c;^d\EOg&CJ[^V7
:/]VN1_[.FLJW>T\A^,Z=Q5.,O_?(0^\W^Z,DX,5F:O(@B/4Q(YS7A^CNFM<O6<T
UMdKJX[gdc]0V,e^Q_>R+N-=c=NYZ\1d?@?a2<P:9VZGGD4RBQZRO^.TRJ;+_PI;
dS&6P?JaJ8.X?Oa^]#<8fX?72K&R7;KUGSB[9G3#)^E:KgK=7IP3Ye_DH>3I8a#0
JFb7EG](YdZccaf0O2:,MgPS_G5A&CC<=X3=?V@-4T@V-2;PO-0,O//7Pe6_Sg8C
GGCVRC33<cfY4fEM>-5\.FCR2)d4/F)MG9F;9OU#+=dCQWb#&96H;?@/P8c9N+KJ
Vg,S9cJV61AC1Oac0#ed.;(QW2.bLgFPcY1ARd8\\Ra/;#;Nc]T(G6TO4QR&37XI
V1J7XS3)S3QXNPY3[1Pb5F1M<caX24=VXAXT3c0J?VCE?N:GQ\UAbD[@^HTE(fSV
/eI9WZEC;9W\2/@.=S?CN]:XT.dTWJDTPAC&H>_VeeEUDMMGN]8Z0T5&,DS3+>L#
L]TS?eDU[9YCgH#H?XXQHL4#OJ3-3?Rb-QDSS/0a@JQdP_[Z1U(D8T@AT-Rb6OH=
OLDC(X9_1O&KP;PM4U4[UDB^^AMWY@bP7fg<@H,O?_HZ6MLX<bSBTKB)MW66DIDa
5<X1@5:4STQA46/BKL/gE_Y8]TYJV/XfT([.d27?=JO;797ID_?2YHQ6J]&?N\G?
4VR-B4d0<4_PT0(/(d7H=V2g>Occ)IcgYdIR)\S8-Y,QU-<82a2,WMV4(#HGBADb
2J\H&\>=U]9>\:W&?@;ODHBKgD0M-SX/KQ#(ZJTX=^4+;;YbI]^5-63?e(<=IaYG
G#A>41V0)>-80;[C8_++L)B[[)HWP<ffd6gKF)7R/VEgdZYK1WBAM]W1dWUaBO4Z
9O8e^Y,GCBb#UQ6#_NP24BfXII-X,g\eg#4Z+VFH0D415R25R4Ia\;O(YPBXReGM
@W#U2\ILKKMK\gO.^BAO]3Y7\B<@B5Da0R2[4d?0@IJUB>+WcPLS?SG:e.A5CPJW
IY;f3#D_ea6L+f\eWUY:8]<1bTIM)NSe#<[DcRXe(#U<cP]Z;,H12I#I94>Q\LPT
5Q2c.]5)?>+#.LC2OaEO8MSU,SO[+ZD&BZ.5)0M(6>R/B_<)U=0c6LC2T_RV4V6H
;/gH[NBTKPU<?&>cMcL@FL7X44=Z_I0Z6_[M^<H-L4^1f;T]KA\KH\HdQ-=.]G0E
(G<J)N#A65XWF_f<M:#F(57.P(.bQbg<eBVOYZb0a#M=J^O+F&0P.OQJ0d^5I)X#
7GK<ZG1;RG#g4&Mb.TX]9J&JgEaB<R?_]\e_C6#F.d4G[@09GF?VZ221A<\V6Z?J
C1L]8+cFY,VFHA2gee(Oe:YU\eAR#-[TFO?LIce65:,^dHKD6P+F[VN=M9<c@2cO
Dde+GJ=>#KJ]3T8KI@M4Ob33-F0GRVRR?CdY/5VE2_A/F:2)AJRCaR?QaZ?SP)@(
W67W3fDF9cT\/JXAA_J;J2\</H(DN+:dG,9?;;57/([b@NB@IYUCcP#g1GCJ(65C
7:,.c&M0Z0GaVCF0[YBOC^[&f\A+I5/BQdM?a=4:LAAeQV:Zc)2UQcM:/4d#SPPN
[R,M=eXLG=JWVTPb_gdEZ5<a;bQS)>F:;IcFO6T5dcL<2+GR.]IO.Lf)F[Z<YS^?
]4=H8)F<HOL2Sg3HMQE>[&K#)M#C.b&T&e/bCedV,+JQ3;[?EU-cMaVZ7CYCL:9;
GJ=@VMNSJ99WA9H?eE?)P/c\>FC\FFKFVbV2F[fYe/edQDNKRV;J0:SASY97feW,
</L,+J5<EASd,-K409;)\:Oa_e:(<9[<4:)778R,[R1@DE0N[U97#\]dMLD)<+#f
>P05:ZgN-4JD,>e8/L)^LLN4bRBafdP@@&KC@Vb30+1^JgaIZW&SQ;&:_ML4D@g7
/H[A7VVUa&:80eR@O.P3^SS(XS=:O#34NBaX-7FO@B-66Cf9,g_@E6&S)JZW&_]]
5Jb4e)NZZGKe#&892F&fHaK+5>VKZ+5E4>;Y1\9MgI\]Ac45#^.GCT5X_XQS.)>U
=+NP1G4F5LE(?f:[QN\3=7UQb2KA]U/B9JJCV&?J5d@U1gC.&e\^X.7<;1B+Ma#3
F<(JcJ?-6bUT2dN_+/,e9DBPg;M8.eTdd\ZO8?N7L..OM3,:9bf&H>G3V:c:5<b1
YT)#KT=#@)3X4>79<(SDBf&Z.+gcOVK=K9+0De34(bRQ6^<6WX=3=MZ\2E@C[_]/
))RJS87g+G<HLFe2QHP<W3FdQSbUE?4G<J.DURB4[9?#I[KFET^H63Ead4<FSeNK
YJ<,7Q@0=PW>E+)Qf5/g4e_OFP@A<RE:(AH1R<CdVI8)KWPX:G,D31XC;WAEfS0P
BJGaN\N4(AG.101ea)/.;;=\g;146NRLZ7b<@-4&#NKEXX:#d4TW.>T:/@E[O.8b
TKScI,?Kc)&E_(d7[;BH:33/5A?S;.#UEMX=G4aG;VYbL.U_KJX[8:0CdAA/3Dd;
eeL.5<H-IW+gLE<a>>6\?ONAg4XG]-XaSSA4=R[/;J(NGVUGK2=dN581J?)(ZR+G
g..0#K@9QdXCK54b@63A6/RCP7DSd,I#3I/7J8@Z<&4@?KaD=g3IQ.a]9D]S>OW.
[6@+PAc)g.dU)/R>;BVNJfA1a<74#1dP)SU@aV//PPAJ-PP63-GMKM0VKN@9fcH)
4\6\>\g):1&.GM[V9?ETN^EIfU@ZY9W];cK_5Z@\b?PUDGWcBTKCCEC:VWEPa\ae
_:5\_TSLM>].<Z6e:(1aR2;HKMD+I@)@;X0=b+BaL+&<9=OA)#B=B.:eRJ_UcX+e
X33Xc0X)K7,:+Z_?fV@22:^1YJ^c\G[F@&e4/R(42LQb]3,@;I.dJ@I7>EAg)<Ug
5b+0YAg[T7ad;\G;;OD)bJ@OKEfXIK2#g0K6L_XG))=HI;<-/0dR17cKKF45d)F_
b[E_U:\ZbLbW75;2<Lf?dP;VZH6#ZG8<E=^YI@6Og+\gUT8<Y1APfOQ>^^OCb26M
N:\6:G+J.K-g]^RFKZNY7aYSa-=,B;2^Kff7aG?O>[;TSQdCe4UBd\0YKS;?[TBH
:BW_B<?92-D[[ObfPV\R8IJf.[<g[6@1A)TL+F;DTV/^c;g)<#PQ4BDEV4GL7#eO
XQ86][E+?5K3d9H\&7a=_c)^R4DL>KDKY^dS=&Q>)++6(7/-,/>9</V1BV693#+e
^L[D2d72+MZOgFN)Yeg]4RL>08-P@BDP\\1SY/:)+B;<&_DDNM[X]@\[(]8XQKT;
>7FG0(;(g>#=)gK)[e8_///WgF0?T=-MMA0b;HECTXJ,P#YY1bBI[JWPHKIcT^<7
HG+8ZNYUbBNGJ1JGQ)1]FE8O[YP#&&XYe&HE28Jd068MV(eK94/7C]\?DFfcK>MR
A(O:@]7Mf+TA\1+D+^/LII:<BAOXg1<,U<79O1)EDVCAK2F0PK)P/+U7#3QGN^9S
YOU]>=G.\:_\-;@2FW9&:7dRHF@N4]6RL4]LTJWUYg7C@Vd+;D@H^6:E]EUQ.=V/
QNV<(FFJNC]UOK,JN5CW),:OeH8/?M?8=@Kc,5,R:@-N&?e6f?C&+b?ceZKHb^>>
2.Kg6caZa3I(,d+7797U//,3c-6_7gd^F9[f0G0G<c0G75.9Z,0fXQ^OZA4JCa^A
aS:edV=AeH,.?<g&F32_\YgK,GBD9[TV[1gI[75caBHDD,T<WQM@;Q[TXL^>98;3
:4J[M4+bT3#7g@0KR1Y9ZQRb?Y++Y@VR9SE/EQ?b4,M?4AQ[>&J2&N]7\g^43?K&
SFB#C9)Y[638B]IXWZ>+VJ,/b+ETgg92UJbN6,#MaB#UTVRb0__:B8J=UGE6)(BH
g3;[S<OYC#a/UO[K:Z)Z.gg-<?gBIS4fb_JFPE+3e)\FD[2ENc0X:Z8_\)I[LS@&
)6e@8QdbXA/T]52(g(JWD;[Q(DZS]_Xcc_aUb>7-f.44/71&dC)+^2S(d50T3FW8
7/_2X4Bc1>/aF\ANLN8MCdL@OW&LODPbW]WJgWK0b0\gV<K(VcPBV^HLX5[a4<g7
d_dMMAf?cgL#&e>BW>VW3B1&4/;8d>CAe].ZI:3&)2QHg[D)2DB#,,AY<GEH84CD
K22ZG,+T0AUR^Fa:_)INfg:E3\;,E(/(fLO,CGB<7K&25ZHb0U79fX;e;CS:JRC2
=V5)Ig61BZ#(;QZAB5VV5XVfFDI^>+f,RFX.L^@a0b)@XJ6,^DM_BC.29L739)6c
e)<-]O:SaA8f27a,?dgeG66^KI3fG)\E)IENF+Zc2V0449:LZ:g79I/IcMP>R^g/
=2,P)BD(K2S2L2/Tc1N;0)1[:?2;XU3Q>_H?SX><V,>MHBc>MHdF5@6.<8^@:TJ&
&efS7aP++<b9J?.B;UGT@Ec8?1Ld[3bX/#3(f>B9aB(?K)#f(gYac;_V]]K,O1<H
40\]DOXP,Kf]g#@de7926(8/&?e59<;gZKOS>KEN5PEI\_V6CP@Y]=.#KZZMd6I;
[YD+]T./GX0e4Ga0=R_a&XIE:96>d)I(PcDRZ0C#:RLMT_&V-PU.#[6c0U:L<S^W
A5C\7N>O](\OF.+dEYK^QEH/Q)D,Sa30LSa?e^:6LSURec_Ae=bX9JI>S8Z)USRT
8Ec@3cbVbF<V2-S5?2MELP^dEMGV:5M:JVHDOd_B.[Y)KgaF8[=MA9e/QfGegc10
EUa<?WL?7]&Y17?JZ)?BC_RVR,3BO+6.BcZL;]LPXF&[fAG6_4aGCMK)=G9eRF;B
,_28G5YX\Hf<7V&AaE(FPVA.HA5[J]bLbE6eKLFB[&bTS@/ZABTHZJ^0)W^H(L0Y
=5E<FagGAIWO=M(73(/0<cU<M/]fdfE/QX>NFaEYe,]88<EU]@UEW\=_X[@J2GQJ
&L]/]M[H.f3Nc0c_C@IPg&LMKMCFLC+0_NJeI5;YC[4c+>N?EO/:[Y-8SY6(.JLT
<MUfF8L_69.YJFddBEKZCL=PI5\E0,-X;K0+MM;3U-PEbC+R4(8):D+H[\X.[=?U
JP#f1/#].c/fUU]3<J_20T9>7R?8U(g4F9gIL49e&^]L2)/EHc?8HdUg:HfcVg/B
<U\>3((Kf/2MOZ4H5?<7A2=PV2<U1e4MK\KgLE(D,()UR@7>,#VCaAY+91FWDOLJ
9N;6G?.H;&Z\,N4Q<c]ZU:4^ESZg9N@T27G+?9)Z7RGE3HO[[LHSeX)GgHBa2].R
SGce.O(<K-7XG#++F4FDPUS;[TWeVAW:Q+_;FY0F?\@cc@V>G@)Og-I&+;He,1gX
#VIPA1:Z&Ye5QPSH7:XgIgF<#D67aEBS<0DgD?g,M0:a:7?HaMZ01MCD];N-AG5G
c[69F@0N?B:FLY>/=X8XfA\C..7]<D>^B^gP?fY1;73G1V&2)ag[VA.EK85G1A[T
Xg@N))f9Hd37(6B;Q#A)VIUV_CQ@gN&TSQ>M_79+WHScVS.#BdaUZN>MH,=NBEbH
K#BB\&HB+JGdF?&>,[#ab]N&6>(JaCMO5#F2g9N9</=O+:Ne?2N016/8G>@0-/_3
X+0=HRb\];Z)7c5f3AcVN@a,bL_S,3K:\MC)U(K>N<@4._?C\7SdT#TL&A7MZZPP
3O/bZK):FX)TTRW5@=WTa#_4[J549@,?,+c_-\cK:IB:W-4b0/WPM8J1[6_(aKMN
W&ZQ#=C9Y?33:U+0YO)]78/I,aYYJ\Nc4bI=,_NMG=D=]dV;Q[+#]DZD.A+/NF6b
T0/-)Q.VB2U3)/b>>?ZU=,.<<ZKZP2_UI>KE9@/5M.d@Q<g2A.4Kc/ZSc=/G_M<-
=AFBA)QRI):/:LJ=LN8=DIVOQ,@Z-AV5XAT([YdQ7Z8f2.=R.&B:TVR-W,8.M887
Cf7W#^f0\61KDLI-J.e<^Y#c:eQ[M(C]?[:;&F>G?MKd&bI&EDd>6<0P2Q7K<G\N
-DSgP<WXZ]f@bG7Z8:9])RJSDX\/cOLNSVVZ0BbGH2YKU5WY(dW15ca+F;@e.2#U
Q\IR2&YJ]\_XUOPF4Y[&@?I-\-CEJ.d<5)5=M=U_[aOV?^,AF)OM\O\Z:12;+-SN
_9(-U,P/-<:]R>NO@/ACS=DA]67#d>IJGaUPCJV?,Xa)=UK_S(=e&,8Z3SKRPKL-
2eWV@N85X;6dgOLObOQ/:UJSOEJTNH0_X7E>T,9,I[K@GV18]4^>^XHOU6R2V0a?
c;-[3T>VO\3b/TfS9Lb&IdJ=T@<F0^]-+=B0Q\AW.f4\DY/#7cfDW]:7/JC3128L
G6VfD;.e&e6LFH(=<.>TQV-gL<D@&?_<I]3C\)JUdO;?_RgFF&YaN2Y]TFM_dBbF
Ef,V8#+24MXfCB3S:a5E#LENg;E,M.B/ZVKSJGAENXHQ:F_X&g)0\AB?[WcT;bGa
4Z]E42LIDfZaAONGCI@&AC)cT_1KE4\5.0@3cbQ;]YL[JXD)a>@^ePQ5&@D1[)8>
0O85LUXAT2AYX\=NZ-]MSI[1AB9?ERNY.4)=.0&XT]#&FM-E&MO)MWJY9bQG:DcJ
R[fbJP9:O#QVJ<N[M^SO-eB#N^RVTSe9_Z7d9QC<8HJS7)/;[[K^@RLXF(/NG#QE
WZL_;-J=7_](TgK[T24QJGHQ0DJQSA+)7/]&JX^=+W+P.SLNH6QAg)+#=Q=8GSTF
<DB+UfaIb#6?Q#Z4GHg6A)&V::LM9Q(0-[U\9,);;8<Qe^UL47+fU,)YaR.Y7LCX
T.H=b5,GKYTfUDF,N2V,,/LWNU7C6WROLTF)[f)BbY5ZZ6SJ2c4<b.0SM>\eQHgY
:<13+HCWgeLCOY1Z4UT>,5Q]Re9/\W#@Og:Wd?CeLJ2B/)^Ra.9KZ.GLR4P:0BJG
/QTR@?=TT4U#f)9&d+W@B]FA6PeG?e:,RG\1V<7WHD#MM(M;6@e62;T/G&?=>H)\
\]&&,1S/Rc.+d>=&g?Y\g0XHMQ:__/GQ^E<XYO<94R\]agS6SeJU.&1@Md8.cf<G
PUESB)V@bA]H5Qba&#g8+5gPC2g>MN2YKF[RW-^KP(dbT^_ee]D5a@^SY9INLfL1
f./D;Oe381U<:L5Zd^C-d=Q;GW2NP7+40S?M1+Q9S76/ZSSbBP8FeBUeF5b()0e-
WT1a<Q0J=A\TS3d[?14(A?LeS3SI)Cf2964N+ae4D6+>657H0);(LA7a?J6<eUR]
7O?6U(Z(/CGDI?U#8O8&MU:A<.CgP-^9UQ/-eD:6M<?9@P1cE0.)^GM/gK#6JVT0
e\gE0-DE&KF5egY(UM:]2f>E_c98WCKETea)MH6I.EP34G9GB#\U5CTIdTI,FBS)
4S3a^K[ZI1<\MdNZ)A+S:[TaGVO=(5>TDB:];;#JSOe@2;K,,>e43G>e<:HbM.Q4
gQXAG[SCf2c(C<7.dS9D)C@KU<,+g,Y4U_^+>DbH9^FU[D?beHg17[-5QeCgK#^U
]SX3Ld77ENMXH8f&D;:ePd1<B[Qg8ed;U.JG:5O\]JC8PRN,MMc9@B?Cb\/#X\d4
5>(URQ&cX-[CCN43.YZRCH?/dKF#4Z?0@f6IV<8IG-1&E/IG)8gQ3,Cc^cA&UN9V
CA267N<KF_dP7&@bRY;,LLS+J;X-QR/2A9WKJfS<174DX[EG-.CG[[/;\[d^6?)V
:Pe5;2D[Ad):@g9=/DT_R=:[R9C#[V]08#c_2LB>gL;]&F@2V,3gBC<>[ffC.)Y(
[9ZYKJg(B]739JQ/LO#Q,2]>3OXfHNB@O/0RbLE8&QO>P+:^17.+)-6HK\D\/8QE
5EZQ9:EDJL+L&gA1KH])3bW<0#])42J/[.O1)CEc=ISB[MW+U.W51\dE6;(AIQ^;
(&5O#CbSIPMR7):<CJNB/eefJ(?8116?(MB<))XX-,M6]>Pbd\ePV-4g)]\3M&W#
QLBVCV^\?dN0#XAg5^_01Lb@>@MPcWSQN\<DYV08\VL0ENQ-;MM.e60K:;C-g)>D
TeDUZ>4?EP:U(#HM2RC/V40AG_?=;)+LCTXbS5N^VAK2He9-;C>_dJGJYL=_+RV(
LMZU(VdaQD5J8#MQ>>6TZNb9c/9C5,8U,@Q(8];F4+2,UGBUbcB)(E73NO./dS>D
JJ#QfL?bTE^#VYKTECT.,AOM/<;UOHc9N^K/-R7^Q;)S>X//RZIDI2@LT=H;b.OT
X\9DKCKbKL6DKMfIQ#>:^A>d[g1X#@B;b.138[-1WC.G4/@eA_TXWR@IOb21@I@X
gN(2bWQ:SX&B+[ATY@P?^>_+WP+J=Sb@fPX>73^e]8&]gXc,La;X8[4I,T3dOU,H
DT)G[4?3<>3>M57J72Z[,2^Z=]),QTK/FF=FU+4:?cW4DB]PeFd7O=#MZ93&G>MN
B=AI&,S/8>c\U>CB[?A9E.c?KQK-7?[aNb4d;dI+Y,bXaFVY/0]6#?g^CJJ4Mf,X
SW?NFF4:aM]d#^[aBS?X:[3/Tf25.F3cL7f2W+:J,dB;)/3[4U:BUEYO_7@T<g#D
P12?,0521YI&).a:__\M?>E8>9]e#ENIJ3J9)C2F.?6Q:Je99\)]T@1Y?PM<0N.N
]#AWKODWCFEL\_7F-@&XL/NDRdSZ\:4L0F[4^67)PQHg<N6L7EK18_W-A7X</<fH
a+>J+5PB3X^I\22^0,IQ5FMR<g.98bbJYS)7U2#J5(BQFX;G#FUYW&^-)bLZ^+QS
3Y5V15QM@(_/_a&8QO54?Mg8BR-?Uf00fXMf>=P1V(5)@PGO/Y(D7T-^I.)<+/8Z
BC,bNR@^E>#>eaAGcNOI1TWDeR8,6F@C-6Cd:EG3>ZAGZc/:7a1OF3c&O2E-CMJ>
;/5dd:)>\XQ,Nc,RE3L[;J?f4Z1KS9\/Y[DA/e;+:2B;+F>FC8>]FFaY@0>I#Q1+
P.58H>Z9@a.O2=K_?5TY,<X&A/;P&Z]dOa5JB@G5/ZeFR@2[;++@@]XBZ[?aFHWf
S52)4@QYVg^94YN.,)gRe92W9S.f+:1X=)eE\IWHa_X[T8EX^d.]M;e1],Z<AJ,T
g8DdV#TU>D7#/+OL9Vfe86=MR,BZeAG)e<BdS-3/UA.B>I]##)-FI4:\D.M;cCFG
4)[8Nb-cYYJ0V60>N=V)AZ?N,MJD[RR^b;7IXBJM80;B;#EcU:D\ZXHf7becPDc-
.?4Q9Q^0])&7^;HS=dR(WQgVLPH;-;c1)3f8>W+[8R6KXQ:[7b;_dSK/3HefQD<&
BF1P@EQM,#)PJ,MH#(eUGf5LO0fW55cJ-0]c-EM\H/g?NWR=-W=G1E>-df0]/g2C
Q8bWcGPX9.S.PEcfKBagWW&;U2>GTf;^;]Rb/?.XL;OC@CC2cgT.8&X.+^+F4Z37
]QY;)(ccKC<c2dFY(C\NIOE5:E]IHDKb5PdTD40JS@Lb5PHJ,)<8;bC^g(V5W&UR
C^#e7(5T]839b(fK[RB05.KRXf^B>1Y2\+PEIC+d0CZVPJ?\FcZJ&+HS66=2BeN4
0=I[Wd^^G>\,dJaQKYJ@8,5DV2?J<^(+HG-GHJZU=Fa^LYeUH2edU<<\WXb#9_gM
?;3XDDSUY.a:4WRJg,S3gBEM\&YX(D3?7AfARGgMfK=/4?feAC[OYY8;[CM+Qcg?
0,K;4ca.=RV)FXI#07Q6OacAH)VQ8ECa)-:Z.M>a+2;YHD8?X-]@(dEF6-?EURT2
T8:/I@@3(FW(WHffMKN29X&4WEXfAebWE9#S9PUcVFeZIc]DONZ=d-@QHF6M5<L8
]8[W/1(Y4a-^)]Y#?@.AZOgA7#W1F^+ZP,6dNb@N3aU)GHST@OT:Rfd\gGKdHCI6
XWWgY6J[F.\NXDa3?P7f0J_AM^ORFS\H+O_RLX(K^fTUdaYB]G4b<5M5,T_a;>RQ
IVXCY(XK2Z,@J8O85VSUWLZS_84=gA5I6dGB8cbEK2)QN;I-UJ)8M,RdO[\QQ/U-
E;,/_H6ZYZ/b7cS&7]Y&@PQ6f6&cBAEcJe4ASA2K5X94AgSa\(F71OF+>40cZ,]G
E]I]-9IQd]@QQR=O@K5]QC5&VN-cLE0<@@d7?<#eeFLWCT?S9T<fbBCOR^[gO+O;
>8Sb&J+/=0-/R2I]T5XNU?N&3df/FgV8A5.:BR^2MQd/(?+YeCfJGPO6RK\R6),<
_ZB.<Of7.T/54;b[D\H/4:e?gWF(B1Ve@M087.6^OPCB(]>^JK6cJW\W>C5^Z=4L
bUMW/_3XcYaARJJPN&Ig6Ag_dbVI:5XS>XC>GUNH]e_7^G8c55O9-L798(_;bYbG
e27O;,7RfDQY,ggYfc(X<CF#3M9+O+^PXa]cT/_TaAU=.Y@8DFV(O,-a3D6LJ:10
0JCW_Z,1>LB)/PA-g.?A)_Mg).VP]/+e/A)K22^6H8ARL><<bC\OA23J6I7E<64H
@804Bae-GVQ6gKPf<U.(4FXS2=4H&bI5NU?Fd,AFRZ7.<03?U,cb^/;QZ4^K-9gV
N+L]M;D-.(>T(I#IW)+aR_=,=7D\9cSS?eaK_0;-eUFTaF00KH8@>&[gd/BX58=;
](eZY&M9/L13U#Qc=I[6M)L)XBYg/5:B?C(EJG3]6J8bYd:+5KO&7\;)D0]^(GOO
>Fc&4T5[,aN=SR80(DC,G&96S<bAICI1ZD;0N\4^Ycc(#@-CXX,P3[;V]f7X(T[W
5[(;]O74(<2:6Bea94;2#cPa]a>YW+@#08gaTdg)Y6#2E)PgJVMH,<J/,HB]Y&JI
<[O+K1?PfCUB=@.&W8>XdS:[NMI=,?XD6:VG>O:gOZ/D?@K)MG,>5@VJ@MBgJGQ\
3^1aCOA>A)?YJ@>XR/S=J#6Sd=N[9Sc8A1_a3Be^.Od=bNS+IUQ<A4.,EUA>I0?J
M]E+?KI2.V4^[&MP0&UD&TN8Q3]ZWN,,E[de(ENQeZ(2HNVbY16MGc,)_9a6Ga0.
_bYMF+U3.F@c@/C\ZF?=75P&E^1Jb-:>RP0Ddfe2]=D)b:F9.2c8(aOMP<XcSK)A
=Y;f,PV/AF85G9@2?>4B=3E^Sg^]3Q:Wc2c;;)2C-^O-?4Og#2bYP==b@H&8/IT;
BTaLAX#Ibe&)Kb&M@(.PW=0,(>YK1N6O/f^0/L(#fR-TS6&b9]>(b_CDf98c](U0
M\5I:5PFL5-fF5O6UB414f4NL4@T?+Xb3J4S>ILdf^TF+[PeQJ28cZFE:@;4RQ71
;EfOFGB#=EKZ#K])U5?Oc4L,LIf&X-6f0Ig#&4&Y?+<2?&NFUf8[cENdT,F?Q5I@
OGb\=VDOSM-)87Rga3;LWZF7MaOFfeXQZ<Y&][7&.cV&T(DbeO=YL\)-OTAV4fE1
Vf/MD/2DgQ;eb+?U5FXYGN10&ZCg>-2Ke9X<IU@5LZ:36b^>;G3f0K1HJ@&Y\EE5
9Y1(LIX/BATbHZ\B3I=\Vg4ZJ\TCcaQbZ#AL>FMI^g4AERJ;(]BX#OIdCE3=cT;1
V]GH5a=?EeL-0I^caBM0KFgY99^5D-[V[1-5;,F_beQ)?Y\292^EEd2NZ[;<24,d
B);QOA](OG2@b65/7f2F0BgUU(>GGDeV9V1D3NNC@caD^A\<1YBcPZ73?SW&_49:
KPf9?09#:FWFZ4E8OcK@8:2b8>g65VI?<J?]Ag#\Qe)[<d6FZ5EbPVWYcTE+UU3G
8@58@GLEFS6/(;8Rf\:K#/+6_>):<@ORVG2a\E[YR,]cUV+#1T\(bFWZcH,AY/=M
)A(BX.M;Hc=\=[8g8Ka2F@U8@@-G_RI+HS(^G40eU/PbYGVA:KUR6:07;AKS=\Q&
G40a]G0O?,C00:C5F2V]9b&F7eUD?1Z3M0M4ag4b?L9bYe4;PSAW\f<-.ORIWM2?
T4@7>MW@T+&7e)UU2,(Gc^_0ABMUEX[4^3L?[1IPPZR)W@T@BgL4[-LGdP&IN-CL
RaOab8LE8<(8R.16bE7U89OB2Rd5\(T#/B\eTg7-.DOfA#&\dXD@:W<Z:OFP(HTS
X7G(g>/<Z+TM55.SV#d)/#aaJ2BNO5f;9WWb:65A11H?Gd9RZI\IcTR6?befc7F-
N0[N8d]R7M8Q0YCW>KFbUVS[&>#]@#CET=Db\3O7feY]0-^BKXXV56I.;d1f4#Vf
^R#5f&G]NZc<VQea3K;Yf=A:OI9-,P6Eb2//-I1BRg.O<>Z>e5VNL=gI=2Q07ZbT
?V#<,RRJ7GV\\0=X:8Z2eZXNKW5;E\=.3bY2HH:W0cPBQf0JT2W<U412GOc>?LV#
7_Y_8L5WU3[>=MAMHTGd@V+UKadJ2ef6?/U<HFCR:Q,4d5YC4.BPZdY&5,,32bZK
d3.3EO.]&N0<?]R(98G^X>CK^FH((M7-XdM1;N[Y-S<CV6E8>^X99&<PGH?OKK4L
X1II2CW)cQ]P?>:g0<6\7d.30cM#UNbZaR6b6dBZ(ZOb42-OeV[/Ca^Ce4@@2fGQ
1/W]((;8-5F/ITS40,,0I28SH0GFORTXE]#U\XM:=M5OOU?4N=Y[gA;/NG=E(7/c
#GVVae90JaWS9B@ZfR?>80dSS^CWM8F4[.154ZdH+Ib))([U:J6+9CIf5YUc(N?c
>MRKMaLO#-CT9/-T_EVNYN_CeP.,9<,C(T&E9OIIcC&-d=<JSP#Wd5\SJ/(;R+=W
.R9BIOged(BfK-?X03(V8Z:ZRY8gJX4/(URLW,.aOC/>1a2ES63#PW[3/E4):b0?
Z6^T&9<>J>1&1d0C0B1cJ=#--27G9BXRN)F>@.88868FN-^bSGW&57NL=eMS2H9>
^A[c@49,4\LT,H>4g^7RD=2AF7P]R7:E#/M_38IXOPGf(;D@)=]KUD.GBA,WMAV4
3UM<\4LG8?GF_R=GYZ3UdDTMg1RJ:=LVdgQa>b^9+(HA[fF1bJ0G?Lb5?e,C:DBb
PX+M(HZ?f8157Y2HX#E<C9a-PYS@R^W)F19AWG.DfHK?K/U@J/a8VT46-WP:::b6
?TFYW#5gA\(\GJH>II/Ge1#[K0#;(5)#M=\Y(]Ca^KAS8J2M7\C/YIWG>?=^XL>>
7=6=7e<3+/d^DYK-KNX+_0K/@3fN:gSH5a=fT3\]O#^dYGd6Y18[J-c:<6CS9STa
1PeRUMe<T84#S2R1<2>/\9R]VW>4ca3W75/5-gT)I,OBR\A3g.PL;(Ng<\DIA/d(
IZIVQN&N/TfTG5[N(c+KPa;G>.;DId)C-5\_aSQ7R)U&_dQW\9NL=7?#Y#,776=D
B,9]Q<7RXgZ5MTO(U_HeWIU/.L(^accRaX73VKYf^]DU2=F_XPG>MDFZW>TV=4ef
7&NB:^cBbR0.>b+(0-gSL8gd9>_@-DMYUXJ\cCeQgO(W/e6gXY57N#.AD\N;?eg+
f(dM&)8gE0Kd>:_XNE<G;&c=\XMK/)c)Cg,(;&.H8cE1X10X7a])f25VR-0AeR95
Ge^XE]7M=ER<A^4D7>M]VXTB2-DQT^5_2e+O=:\Lc;C@JdE\V3;TH5eYVH._gPZV
DN50MJ@B2F\?H#XY93eAT8/(JR@?f\]FFU4F?f+.Wg>XdAF9;1H]7WF=L6BJY<TL
-8;=F3@ab/]Mgb2TRH\3.UP88Lf/(J>K7a+DWdd]0-_0#K5FO(aH3T./F_I^HM,-
^a0/C1V&+f6R7f@C@LXVA:YOIZ0\-W&^&2QDbM#<O/5G;&OOVc^fe5>\;&HD^VM(
b)VITTA#B9?.I75)3:d1VM&0U(QD/,9UO]4aO]^-GP@?@H17[>GI:)^,@)-ZA6aO
&9W82F^-1-dJCP7(NL71^6K6)LVFMLaVc>1A+BEgb;,5)U6=@5(/c&Nb5TF9K1-E
MNT#,FNbd56a;O.dPTK;B1_Ib9.+NZ>:R#DQF>3?/a^KK5(JA<+8JY.S1IPa>447
4+>JH)-5f;&2OKHgZHDSeH<1?MR_B#gGAN/AFfZ6-bH6Q]c@EDdX)?[1-ZNAQb(M
9?X@P=.SgfUVQIc=GagOHMS#?1daC/9SZb2+(GB(S6(O.:I7XBRP)LdI_I;HZ^(/
fLX3K-+ND1E(6VF(W^AO<&&g?P^X3=-fBHd<ec\TD8KG0:M#1MQG20@@W.fFEJ_g
degB:&Fb]EaZ)/Cd??KBNV3/QK+\KFF\NDQ4F(\,\Q[BN?PFL\<_&d^[I1>J]B#&
O6.WJHG([=I3X0c>C8L_A_H:c7X8_P)c=8_OB+ZC0<H?_]O5_E-ZL:J_5ZbF><cN
-(@C?>g/#@<;J]>]?KNG<7+QaEMb>e/YF]Wb;^2G?U=d(VWb1QEOe]/]-+H]2/_Y
YAPT;>UU8I0.)Ce7^L+]FQ:JY]&QB@M#)bYDN:b[Le<NBPa.EWAdER\MIeYN5/P[
^9:g[<?6^J^eO=R.3^]MO?cSJBb&MUd=I=TH:IFV+NB)GE=>O9=>H=:X^1]1T#Vg
GWXU^fY,F=W.&(Nc3cNYZfGXYSLg3S3QO_F@KFM[S2]]0_Qf#1RL;=GPZZP64E//
59Y0;]bMYIA:5M0014A30)@+?D<TDPELS3eR[P+3e)RC.,g?Q6RHF=K2\O=SJE[S
e+#XfBfU@]E(LAATa(RaJ>XZL>VU)9RV^/+LU2aJccK<2<0A(_geQ0g6,4BS-V;@
Ga-gd24C]OHSRg(E)6R/A\D,8]eLbEK73;U2-(0+6#@RV/FTb/3BUL4dIP^_9AL@
PC+O[HZ-7;[5N3V,__0J:H6M;?2P[,0+FI<Gd_[C;@b.&_D^GC]_EP+Pf^M5)6@/
\bXW+_g-(++WV874WA<N[=&&.^D\H54bR^DD11,:O62LEZ+,JEDG1&d4-RGA.7RA
]:]_M?_435O/2=UNe9V-;&Q#8T3);>9<HB]IeWRER@A?O4fZIO=6e;4S#@/T(Jf)
&gbWG=PBdUMG[D-<M45S[\g^=fD1#SJfV@dOJ1<aT2]KWf)Q2;?WG.:.]^d2AK)D
P31SU6]N]FeH-3cU])c25G]6N?P2L@>=+PSL^+M;E0g-1G+A;eg=/Uf=,eQ-bK4B
4^NEOOaRS(GZ4-BTFK>@-ABO6Q;KWK;H_a[C0IQ1ObZ>1B8Q;AQe[=1&\^K[@7HR
DX]4JC\3KQ[;P?#O-FeBPCQ.Ua&LAS^,(;\KeH,JS71ccFgdP?RE6)W=CX5Y0RI4
c.#cK[^\UH7MB^fRfD#_4[=O-(M1\H/Y1T_UK^6.U4HQ^DKR,:OA+YcfG7<N-P8H
b5a]VL:Tbe]9:?Sf=:T8KAA;Qa5-cAK^FUE^+gS5VD:JMOU2VJaCO.==.X/0G0UD
-W4GFaJa?-TJe(0V]N<FKQA;5$
`endprotected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new configuration instance, passing the appropriate
   * argument values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_axi_port_configuration", AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`else
`svt_vmm_data_new(svt_axi_port_configuration)
  extern function new (vmm_log log = null,AXI_MASTER_IF master_if=null, AXI_SLAVE_IF slave_if=null, AXI_PORT_STREAM_IF port_stream_if=null);
`endif

  // ***************************************************************************
  //   SVT shorthand macros
  // ***************************************************************************
 `svt_data_member_begin(svt_axi_port_configuration)
       `svt_field_object(                      sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(slave_addr_ranges       ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(dest_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(source_addr_mappers,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_string(source_requester_name, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_queue_enum(svt_amba_addr_mapper::path_cov_dest_names_enum,path_cov_slave_names,`SVT_ALL_ON)
 `svt_data_member_end(svt_axi_port_configuration)

 
                
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /**
   * Assigns a master interface to this configuration.
   *
   * @param master_if Interface for the AXI Port
   */
  extern function void set_master_if(AXI_MASTER_IF master_if);

  /**
   * Assigns a slave interface to this configuration.
   *
   * @param slave_if Interface for the AXI Port
   */
  extern function void set_slave_if(AXI_SLAVE_IF slave_if);

  /**
   * Assigns a port stream interface to this configuration.
   *
   * @param port_stream_if Interface for the AXI Port stream
   */
  extern function void set_port_stream_if(AXI_PORT_STREAM_IF port_stream_if);

  /** @cond PRIVATE */
  /**
    * Updates domain related information for this port. Relates the address
    * range given by start_addr and end_addr to the domain_type in domain_item
    * This function is not expected to be used by the user. It is called
    * internally by the model when svt_axi_system_configuration::set_addr_for_domain
    * is used
    * @param domain_item The domain item corresponding to the addresses given 
    * @param start_addr  The start_addr of the address range corresponding to this domain item
    * @param end_addr    The end_addr of the address range corresponding to this domain item
    */
  extern function void update_domain(svt_axi_system_domain_item domain_item,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr,bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr);
  /** @endcond */

  /**
    * Gets the shareability domain of the address specified.
    * Returns 1 if a shareability domain could be found, else returns 0
    * @param addr The address whose shareability domain is to be got.
    * @param domain_type The returned shareability domain type
    */
  extern function bit get_shareablity_domain_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,output int domain_type); 

  /**
    * Sets the address map of this slave component. This method can be called
    * multiple times to set multiple address ranges for a slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * @param start_addr The start address of this address range
    * @param end_addr The end address of this address range
    */
  extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);
  //extern function void set_addr_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] end_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH:0] addr_attribute={1'b1,{`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH{1'b0}}} );

  /**
    * Returns 1 if the given address is in the address range(s) configured for this slave.
    * This method must be used only if svt_axi_system_env and svt_axi_system_configuration are not used
    * Typically used in an environment where only one slave VIP is instantiated.
    * Note that, "addr" provided through argument should be untagged address i.e. address which doesn't
    *      have any address tag attributes appended at MSB.
    * @param addr Address
    */
  extern function bit is_slave_addr_in_range(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attribute=0);

  //----------------------------------------------------------------------------
  /**
   * Method to turn static config param randomization on/off as a block.
   */
  extern virtual function int static_rand_mode(bit on_off);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);
 // ---------------------------------------------------------------------------
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  //----------------------------------------------------------------------------
  // Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode ( bit on_off);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * Does basic validation of the object contents.
    */
  extern virtual function bit do_is_valid ( bit silent = 1,int kind = RELEVANT);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern do_allocate_pattern();
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the AXI SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AXI SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum value for range check done do_is_valid().
   * The max value will either be the MAX macro value or parameter value if 
   * paramterized interface is used.
   */
  extern virtual function int get_max_val(string width_name = "empty");

  // ---------------------------------------------------------------------------
  /** returns total number of address attribute tags which are enabled by setting to '1' */
  extern virtual function int get_num_enabled_tagged_addr_attributes ( );

  // ---------------------------------------------------------------------------
  /** returns address prefixed with attribute tags for corresponding address region as MSB address bits */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr, bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_tag);

  // ---------------------------------------------------------------------------
  /** if tagged address is passed then it returns only the address part corresponding to the configured addr_width
    * removing any address tag attributes appended at the MSB bits of the input address value 
    */
  extern virtual function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  // ---------------------------------------------------------------------------
  /** If indipendent secured and non-secured address space support is enabled then it compares two address
    * attributes and returns '1' if both are identical. Otherwise, if indipendent secured/non-secure address
    * space support is not enabled then it always returns '1'.
    */
  extern virtual function bit is_same_addr_attribute(bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib1,bit[`SVT_AXI_ADDR_TAG_ATTRIBUTES_WIDTH-1:0] addr_attrib2);

  // ---------------------------------------------------------------------------
  /** Need to enable enable_tracing and data_trace_enable */
  extern virtual function svt_pattern allocate_debug_feature_pattern();

  // ---------------------------------------------------------------------------
  /** returns ID width based on port configuration and user requirement.
    * If read and write channel ID widths are same then it just returns common 'id_width'
    * Otherwise, it returns read channel or write channel id_width if rd_wr_type is
    * set to '0' or '1' respectively.
    * If rd_wr_type is set to "-1" then by default it returns minimum of read and write
    * channel id width. If use_min_width == 0 then it return maximum of read and write
    * channel id width.
    */
  extern virtual function int get_id_width(int rd_wr_type=-1, bit use_min_width=1);
  
  /** This method returns 1 when corresponding slave port is same as path_cove_dest_names_enum  name 
    * and is_register_addr_space for particular slave port is programmed as 1
    */
  extern virtual function bit is_register_addr_space(svt_axi_system_configuration sys_cfg, svt_amba_addr_mapper::path_cov_dest_names_enum name);

  extern virtual function void set_cfg_for_rd_or_wr_only(int mode = 0);
   
  extern virtual function void set_port_name(string port_name_);
  
  extern virtual function string get_port_name();

  /** Method to wait for next negative edge of internal common clock */
  extern virtual task wait_for_negedge_clock(int mode = 0);
  
  /** This method returns axi_interface_type as ACE_LITE if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set axi_interface_type will not be changed.
    */
  extern function axi_interface_type_enum get_axi_interface_type();

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_port_configuration)
`endif   

endclass

// -----------------------------------------------------------------------------

/**
Utility method definition for the svt_axi_port_configuration class

*/
`protected
5?Rd][f4@4AL[@c]DU?Lg9C0P-KIW?U0AK-(Ob@B2CT).K6D.YT9.)Ta,FA9A)RS
;R;9e:OEUA3RP9/3>3M#4F/5<a/5bPUe.Wb185L@Q:ZLANJ??/0d.fW+A?=U?N;8
6OR-GLQAPL8-c;\FKa\a2TZ;ZC>)c.CU4>HbHO;gUE;-HgOZMVSLJ/XQ-V@)@;LW
.#fRCJ6OVE9/:O9GDB\cbPTQQXQDAB40K0=C[#J09M]U.V3(&+TU9R4\_(6d4]<W
c0Lbd3,aF679S30#81<>:@_=5SUFAegZ6W=S]A^d;/+=][K39P-=YbHHPWR0[_9f
d@W@P,<D;K-ca?50<gWEa7BdWLRXI.]/PT_5EdcCE2??(HYNI:4FcX\^/J9gDU7f
TQgK/QN8PJ7G,5&T=;)^\085W\^?1JW:<&QGUTWBLgK^SU+BV.C+8]89gYUa1CT,
LV]eJ(ZH8=HL)BJQS-GOEM@AQ]6NBYI>^RDd(4JfLd2R#2/ONcegf->J.T3,C_=C
.DA:#WY(DeV9])=c:0ZL=cB[ag><-GL_180RDYBa?0e9daW]</0ID)815Z[MT=E4
5]d+N[[<+:(O^LRPD6ORPa;CBb>EKSd-L9K1X[#0#IE5H\F0G;AZ0BM]558LZ1JU
c-KG)5+^3)PTLP94PD9I@+XOa?S+#5-[c-Vf/P7f@<UL)J&F?Rf(IS>J1dP]L=b3
PQOb:+;2^3gPYTU#M4UYIc(+aU7G82Pb\SP):-A9<>L/-4bA725VUaOI8.eTV0-e
BEJ3DA)OTQ0U/9\14X286DG[5[Ga)/3+OL&0fIc]aT&aYBdQF/HO[e7+N5f5]UT2
dSC:G[bXS3.,@_HQX@(9L#-^P2/@S>B99Mf7@L(-LZ/,c0/\1R[YGRMZ_7d<GJg6
\W8VM0AE8[\PN/-S71d]4;7/D/+Z()A[aG>W>?S3N0=7g[c@;LX<;L3fLG&_c09O
IC(>A;_afP(90;YA6\A=/\P9N,g,Kb#cPb0@g@Hf/aK90DDAA9P;6EQA])X3+<<<
WF?BS3PNTB)+[a\fU.0A?Q8c[XK.e=YDETN_=JSW:gg6FN[<?0),)],7=gHfWYEe
>-QG.2QWH;>RZ9>I&:=C2XHNC_M(;^W1VCWeO>Z.)XTEVd/)b3(PC[X+3LU\+N)(
K<T3<XA[T_^&>QWC.D8#/KeT^+Ee+6\2a+SbI5QH5K^a&;[^^US=EL/aPX;F:>.+
Dc)P&bA)D:a7A1-<a5+#YL?.,bd2ND5c::KdYK/QHRMPBAVQOM7aCdF:-7XEYE.(
&,eU_afVZ4cA(>@Sg_PO:b,LG-1FUM7Pd,edRc762A3ZI<=aW=Y>ZEKA)7P\V,?c
@;V<.60Wg#8G6);9<TXE=5K[J+V_WAVf1DB&>6b[?B93#+U[4CfJS.5@UeKBa./&
@4J^SddUU9aWMTG,0Z+QJ6T==aeC\.C.W/+8-C_<.EZ7=6V5-G7;PKOR^daf]8RE
/F;N9dQB=UFGbS_c?#URQR.QeF(EG(N]aSJ;Z(/1bYM2<R1R]O-)Z2IU)(7T.fGC
e=JeGG]0#)<H(B(;_db(@/7?#;[A3DX[S+M^#G2I+&7,Q^EIdW[/cF]RfW;.dc5>
7Z/<M/03O;(dH[4eG[X)BJ]/Fc9M9A;AZ2^ER0=Q3e(02XYQB4B]TICI76@\&&b:
\aZ4)7)CHCP#9Ue)VRa-WKa((aZ-2M6L;&OD@DW#5HSW=/S;RLJL/gQFR,)9AGM0
C[9I#)4WOdOVbU)[XNNe&^1D#SWe0OKF^+++JM4ad7E^&9OR]5TP)K7-G,1YY\G<
dE+,a7Y_G8b&8)gI1>FVLfIP]3BIQ#dWVCg9(-RA\@Y,YX7W]AFGQg7Y^9[V-OKM
BE6[C3G2@QM5VI6AC#O4W58HO)&I5<3^H+aF52+<,>:fU(aAMB/eLJ4J_1Y(]a0#
QW6I&JB7M9W>6MJ#c9@ad-\XS9cHFV1d<KEOF4TZBbWLM)+\OSH<1C?N+:->OF6I
2L,MI4CVa>(.C)NA\Q:Q-QLAgdMJ7FJ2C\@^GRV;Xf[X_,.^YYMI2M&?dWd>TS=I
X>,.SS>6[gR00QUTB(dfN6,[ZcW)-RYQN=8L<ZaOK<YF-T@Ia>(8[ATZe<\@-:S#
\Q\.G)]^RbLAO2J]X?B99g]ZMLfD5f@7&DAA;U=,_K0b@J4GXR:=</:,HLFG5<@Z
6)T;F3P?3UaFP2a9)7.>:OTe2+NYRGJ,ON7gb\HW9U-#3SM[#\d^7+O[0R9D&1HP
4OZYD0F\665<M2/./LJN^3d#7(4FLI#_4C>OU]/)GM+f#\7Y?/E95^>JF;_NA6BA
X7=Eb4AJ@T+@&.F&DK<DYg3WJ-77+>FAMHW;]AMMZf=I[97J;D+eI:9\GLI[6dIC
gFZJF?gVZ.@]9]&@?Q2IN+dHOEcVOW@Q86C:^D6FNFbAeY)^8,C(DMQ(^.]TDaXT
G+/aH9K[gcCB+SE@dU6Vb-E_+ea6>-Q2.T;Kb6,RQM^HMKE_3V=-_S[J5:F5(PUG
_#38P488a2E&2WQUD)U(P<A#BGM<K\GZ3L7+8WEgM^4@K62dP<8+SgcZ\<RQ7)FX
7B>:UBZ0&Oa9F;B^Kb@_U+R9F^bI[K&-\+6,9c@P>))H7EB^9F>=e5/Q?WYfP37d
W>;4ZRBec>#S7d4[,VV>QK:RW;)a91^AC,=dK>1TD@\O+dJa;;\5>7H91=_.gFIe
e(^#RK?M<NCGME[I>E_0+61@UU<@CA^I9)]a2.7eOb5JE8>844:R&WUgYa(U41;[
0aL.(/Oa17@gL(b2QJY1JE6;,/d3ILa=fLURO3XPSEB9JL5[\_I.)@_aT@X./c,:
c+@BUK(PG441(.4ZI<2@aSfYg<HWO73NZ<WZ1/3U?JNC\L^EZP6:_JLOWIWGb(#?
8]CaD)@2.TCBXW_RcAYP:U]#EB8X-0NBS);6YC+CPg:[&\SS/Vf\;_?^4?172NN(
aJc8.LDRH>BG@YUY-\5<#3;LHUBA\ORX/ER,OWa84<7B54GP^O-Sa_IISb^P5YT)
L5(,VHe:4.+TRfeFYDUC(N@7Jf7DbcDf4,ICDfGIE)2.f_COAbIR<fS,B;N0Dd3Y
fI=SCIJ=I2)=LRWR1Uf<HJB:08#5+\6KgH;2Z4<LR;X:4e>LBf2SG+OZ6HZ5@Nea
;(Y@VV,C6:?_NGRB+EM+VEJ9F,SS+0@_bVgG05TC_@)D:eUaF=#bHA14Q#3I)@28
9RF^IPPG).\=8^-459Kc0DSPW;S5e6_[dOW5^LPTHg&XGg(GP)YaWWNU.21cXcbW
\R<F9gU.7e+[eRVB#IdG#@1ATO3-JG0V<b3d/MNaSK[VBR9,Re;S_FadCBVVU9?(
,NEENL)+N_TB_5+VNO<:83d]GfVd9:g<M-Yc0=LP;LgZ,S@8@;DD)9_L.@0K3M#f
6Q^f2FU0d^\89\/IDWfJ&71M(V92DcPA@+8K;_(##<Z_dZ+(IGL)CQD()&5EJU]K
LU=C1NCFPQ@OD?EV](-8U::B=\V,\EeS,O(c\I:P8]g/EID]6X\U<LfYb#aH23WZ
I5&B-?X4@VD6PaRff89I1>MCL^<:B;K99cA_)X2]H\20cM.MU7c;8Ie@=Vd.<8B7
Y]]PeT<4gZ)+2URWG0)RK/1BY)0<,CZ)/O-3ESC[F1CF^B+>gJ)6B01#.B4]UVV#
UBY&CY5&,\>4dP@C]g[O2<EZAL@A&7M#\EX9#K#@a#.(ISFN0-(ZR>[PN#+:5^TO
E.<K3,O(LdTO3>(VfaHI6020U@Z&5a^e\a)6\WOCe-&+dLcC9MB>#IG#9HE</J@&
)J?(UY8EFTM)Df2d2Q1W0XeG88NGfDWbL5M(DIP5][?.TOZIHOTBM.+Y)^DOGGK0
G)1gAR36X&4Q,AZDHOcXdB6eEVG2)8&a#UW\aPf/4#>cB2b<H:S@7g&[]M[;YDJZ
;4A=.>MIaLGV,?gI4aRgQ/M1/O87#U5ef/&.NU^aFPY&WGIRdHJ-,W_O4K2Jd@)1
93SG\)WMaZ6/?4A7A5UV=bU)GPPU59O4ZE#&=D6@P7dO;2d,5aMP9=Ng[_5/d5CY
-:(CAMNX_L7VdMb4aYPU.=Ba_TbaH8T]70R-WO7GCN&R\aAO;VA44>K=RZI6/TU8
:>&:aFG49-2#&RBCC2\\GF\O<Rb#O;8S]?1:Z8J?3DKO&7e[\Z]V.+:G&;FaOHM?
,72QdKE&dNP9b4;FB?8-3RGXaeeM(2IV9J=_14D6BJN=<c2ZMPH6>/H^?[1TCS6L
C00KDdT#R9VZN:&A<WXAd_2)32fe,TeJ^3<65Bb.,U\]R.X2C(GMCAREP;/3:ab@
XGSNSZD7VT?aDg+eB[cN/T>T5T/C5;HA:PD0:^:E1Z1<<ZY/OKVA]2R#&G7KWBW0
ICeUS;Oe>QP1^QUdA8)1LTfReE,1^c[EgS4/[3,Ld?T)3\CT9=]QON0AC=JG>Hg>
GN-EV/ZgWK)Z85^5,LfY<\?#VQf]D6dR>8(<5ca6=e3M5Fb-/abRXR,b+fGM##Cg
aCZ\RVBWe<dO[=JcUKZ8F5)@(2N2XVIL4_8\@.Y<8J3P^3U>V6,_@,]cRAV&A+Pb
@12]J/VcN.]P7UINgM8K+g<d(bT2G5bT0-eAS7I,eb1T3W1[^[4]V/+/2[\]6[-.
Q,#]+_\Z[gG1)W;ZMFJ,DI9^\<5JK&1XHECBfZNaIb/gWd4Xc6O+FY+/I$
`endprotected


// -----------------------------------------------------------------------------
`ifdef SVT_ACE5_ENABLE
function bit svt_axi_port_configuration::is_bcomp_response_valid();
   if(bcomp_signal_enable ==1)
     is_bcomp_response_valid =1;
   else
     is_bcomp_response_valid =0;  
endfunction
`endif
// ----------------------------------------------------------------------------

//vcs_vip_protect
`protected
HZ3Sda-NONVg/YK?W3eI0VXI@,\\D&CHGc#_J4bI\^JFW[E+N&fB2(4I@?>GW_,6
9K=RQ;,J/EeCf#gQ_?@V)9@+WPM=JH3;X;A8KM2gC1;=\Ua/McQCO?fVdY3=T]9R
^0B^3(1dX1FD-C;:>JG(C;3BPaUZ-e_?/R[+K2JX5ECW;.WV37+aN5gQ64ZJ\OfO
,:XcKB/4L/ggd6_PK4O/_&YINZ9-EO._c:]+;/bA818O37V]ag]<##BX2E)LR\VC
c+9QE9=+Y^fNUa7[>Z94]>W&UYWP1>dgb#+>^V;+[/3.,SJ9FJ34g4^,_PfOBB^.
318A9b-#f;Y\::X+48)_TJ@?-C^gWQDbCLT+Y3BVEDI801QM4V44PJB8I3fX>YWe
RA#FYfAN^/79&,?8ZFL[G_6WZgQ=3(2;1XY6a&afQ-C/QG<aUF;Fd.[>C-=W.DNI
c1_C44;b99^0cc-B3>]9&8-NV\XeE-g[A1RF)B0S9T5<&Dd14QcOZ7V3MO2aJ/TX
>D8:=3f@;,5XLQ0R[c^B^ecNd)T8d_Ge(R95A_gPAKg:d?b56]O_)ET^#(F]#_Vf
K?L\?P+;I>J6EX/[CI)^Y2;;1bZf@PBRI<;7TQP]=cJf\IA1?IfK;T>0c-4D;_eK
@]YOI&c@EUc7=>WV@BGgX8N+BWMKSP#G/6G#3X_1M/DKKOJH^9X.#Z+2<Ab<HI]D
M\Q/@A(VXTHC]3Y@A0^0RJDU>eRLF<?#64dA[Xc^U52X5YYMUf37D&W#<HDYV<_<
C_.eRLW@C(e8QE2c&57a]/_6aI/8H0(N.-?(/9YZ\FII4+XaFI>VgDA>;eX07@57
<,W^f89_N<K=;L)INUT)HBGD)#,94A89aG-NF..+Q8#^-J-98c+^4ePDgM](WAXK
K13=G=;T<K^CWcf<V]g5QZ[BE^M/cd8NfZfM]R@+@8eLK\>&H&;fK.c56>eY#@?P
++13eHeK9.;1_<c6>1fFT=#G8.JCeE2feQbL8+KQ-L])HE_+e0Z7feX8R#<BX0X)
T#>Of4#)]W=^1RA/;?UV6N,Y.R8;cY&EE);DTGfaa.V.O\fM;03T1a&CSV69?V55
1a2A7E;[MYLdP6;=3I5^g&FJQQ+;;9X#-4WbaVaS(T8J8ZY&<d1W7g?aI:PbV/\0
HG)W[gIGK;8@LTe?X_&<@76-a?#-aK.3]._LU\EE->L2[>U6R@>#]9T:3UOMZ;.O
+6TN02LSW?D][F+Rd_FWaK0KC=d9(8Y9&?=X;/.PDR^T1P)=&Yf,Pf143G4fLL9D
^+^=].Jd.eb3TbOZV?a]6bBLF-=[E,Cg.3Q_R]eM);4ZIY(dMB.QY[\?:.5d]YC+
/[cSdf1e)VE(bNg@.(R]^65(B[Df79I-1M/g6T(Q:OZd+IaU@DUA-<;8.P=b7C>X
_V<MJ4Pd>>D\EGV,(64.BRTDGI+J[_/:RaJ;Eb^S09=e7gC>10gSZKea8HgZJMXG
-XF[YB0I\+-ggKc,278R].V28Q@(a://K>:^USC1.0d]:_GdRS/TB0I6>)C.B.1Y
\.9H.DA42CbgIc,7c^8g@8b?44GF>#I>4C&\@9X0X,IONL&5/3bL>89\-^EYggb^
cGQ=OW0b2(M-Q_<:X6C+UG5MT2+&GS-C8A70=RR,bI,ESD:T,aLd]g.PRCgT9]U4
b@XUO28b2cVW^0/1]\=C=,MP(W?W2>;;/3M_A8;aa1cJVB)XM(XJV+Gb#F1aBZE3
EZ-G]Gb3V?7XaZ+UM4>19R_L;_Q6#98C=E&V#0C.E>[2&T#W0APV1+U_<47^W;CN
<&dP?bLQW1f2a#(fTBe:M-7&1>0fOb<X3fRVUW[I\XL-[[1L9IGEAe.XQ[]3CDAU
SJ1\.6T3\7GQO8[cON>D>J/bYNI_.4K]e@:2gL,@XCUHcYbHc4YY?GP\YG,aM\QN
DGc+]g<5:gbMZZXEK1>6O&a;#)dcY#314dD3=IB301b3g1faH].]=T8O2@T(c\&-
1[Y)bb\WE.NN83NZ]_;d6#[Ad4:MeO_dcUEfC7I,KdL;c57GRD2(),[d>(I.HQ&<
B7NcVP9/#G<O[aKU<U\))P>=G9<\<:6e\:&a5UN.g\L^2=?ZX1/(c.)5D0BFBV.:
>8fOe?ER>4&:Id&bGAd&\EIL07QS]]#Y#bBE.1M5Y6.a>+8+GKHO[&LQJ+Gce7I)
KNg&X,0SL1H9gM^dOK0U==K=L6cWFe::([WATXeQ_ECf#7#>/)0Sd+2.LUEdE@1?
WPdC6??A],I;Le&e,b6,dS=_RZFXH=Qa+\EOF_2\LKF.NC(2_)^#S<aC0[g^Qc(\
^AfAPBK:CL&A@3^;H;/Q<_DJ)b&:3/0/:I7ASb8NQ[;BAX,FI+J=3EKTNY#1\I^0
[P?S\0>6NVaHNPf@V]^H+IZ7Gg2;I,dBaY>S:@aPJ5YSeX:P5RLN_\G9M;Y5E24A
<DA\>GfF/f/dU@.WbXIFfdGdfd,()Z9\4-#aZJg^4],;gV@]JP>b#?V/1?fBLR([
[bcHQge^D<X(QYMb\C7I+Ra3aGZS<[>QY6BG;XRVd]4eP-9^KSL&@U4Y\V2(8TQ=
1Y47Sd.LMY>:\T)<ZXHLJ1G)8gA@&;CZICIE7ffT37fSN,]:TNa=7T/=JW2a?M68
7;^e4YM=NW.?2OVYJSF,0SX-05bTRcGK1#OX,QL9G,a4/DaUQRg8FC(9O>LWFG,/
bJ3Ne:QgNONUC,aLH_BTf0MN7U#aXL3fEEe86/@g7?.4YaD#0cd0-Ra)2Ee3P_F_
VPW&LAEfM]0QE?D3Q=/6aE8G]7RUfX.67L?5)1dNX3GcL5N,gb[,H8#_@U8(R:7.
9EUA[+M&S_\,;(cMY4HKfR,3Ufg(SEAM;4(fOUOAWbMPe0T=>(QU0aR@U8EZF,DA
8/\8aSVb0gb;KVW;_&2QPUST9dP/^^2EWAX]Z=bc\[9J=62V;RD/(JbeJ7/>GNEY
Q<2(DdIb.f#I.R7QA?TMd@0G8@LT@4.]Bf3>]G1IgSWZ1)14cQ\SZX\UL)M/W\IE
B?7fV,OHZ8d_3YPd;\-RVg7d>DFM48CNbe..TT-Z&\gbX4]VgcD(_Kg1HI49,37Z
e-[;T&<QI.U,L41B&2Rd.Xe7#@U8JWJ;<EQbYI&<YbH:>?.DGXEAO>=a#OY(K1?e
LJP-3Ac8JDD7@+V&0U5M:/&9_Q2bRDaLe[96fS(;gA9=<T87B/KG5BXND9g.J6&D
>DbD+f2bYLQV\OG2K,_+(V<GZW+[b0_d0N7aN&OZ7O6@(E[V)]0PPK=C2#9-7U<5
dg4@<-J^PMBK:G/:#LI+g###Ze&S_\:CcIHf.Da]IZgbJI3^TOaN+->c=L.2C[U@
GSb_1HGScP+:.:8KS+Sf1FI0ZX51H:E3^;a25BXMR1ICI,H\<S&4Yf\N9#CZ4+7C
L,Bc--DN#ZG(e#^]Y:04-E0\OKe@)eC-+]d@,2-N(2;We@[9Aac;DPJfO6d,U4)R
cf(2:R5U(d3JHK/gFA].\@IMA1[Sd[6F()X7H:>aL>MbT:]7;dJ93M(I#3Lf#+WA
&AU#KP2:3[M1U:LV?6c.]4EAB6V8K^DfF<Sg5GeI/1gDJ;09)XX\aN/FeXfTW2(@
Q4R=7T-e[,K;8KdH:M.I.7Jb)\40M&aT=-M^W^7_b-X1L+cORGR.J]Y6GD6b#6OY
H=+eMLcOU4Na;4VG6>NYb=E6Wb\cC0-K08.dOU(7KUEd>/4ARI+N4<&,/:NNEWT6
V5,e<N]ONOeSMLfOeb8.e3PIdF8JZc8&QR/H[9VV+7,_S1-\)ER(f&JZ6gVMF7J8
=F.\F4JdR=JE1BV4QeMFKgFc+,&EG<Ug\LS-5CQPE&?\#[bFY;A>W#6?/KAG+Va0
YZa>LScIP1,a6L_7&W[e;cgCX[48&5ccORH]?E4KTGdb,WWN]ENO?L2W[3KY05d8
SIQ9TM9-ZNUE.DX3A@IP.MIf5]MK,J8<S?/>d4F\VI0a:03Q1SR,MDM<DK\QT78M
:K9/QLUFEOP>dOXP79P#>O9fPF.Z6IF8I66V1+96U<V[ASN[ENM(^SJMEI<@H#==
GP]9H(bL2;RH,]HI(B)JKZ+9S-]K[dbQ6L-\ML+0RK2f72T#V/1T)#>RbAY.8SUU
(SD/\g)2/.7?NJU/8O7&,L);AYNXU_>#6fD?bEc52&e:Q98.\X&-J,(1fT<AJ[@e
AQ)M:JId,[f(2>4#Y/;WIb<LR1@#8G\G5\OM4FE)W+<-V,+CT^?/fRXN49d.)#00
T:UM5RD3KAWd9Z8.R(\UaZW96FQ(CJ528C<1)?U-H-\O7_BKTQ=Q04_aW?0EcT-V
4bA)7aZHHe;6G+e6d-4Vbe[UOUA;^4QZ@aD72XP:H__g.76RA3f/)d6GD.(PQ0Y6
[06SRUN>a2]=II.,RUeD_?_#Y:@V\4H_^Ee)]V3AE)Kf.9KD-dXQH1Q#UD?>=3BX
>H.>f\\4C7Q?IdY]Wa,GX1EW(_[<>AROdX>#GU1Vb+A@1=cC:I)2bS&MD0#(1?,<
U75V-:a0bLLC4K?H/da(ae[[@4Q-a_D^Fa@e=\FXMU2P0;ON0PI^+d]Vbc=][F7Q
(:GdT:8f/De8Y7[=^?/(Ng/N5#Jd(1a7.b;_VB;EAP-\I;K4=7K[dMT8>MfUWR6^
PDP(F+<?&b.FIFJH7_(0-Q?G0M?FX)>CgKbYd:N1J\,>[/MPOceJG,AR788-;;dN
#/99TCMa2,MQe-[H5MD/b9LK>R79cYSVIZAC<I526@#Z[BOM591FFeDE[\+Jc5H8
c3E,ZRB?8]UWFbbQ1&>OY([agTHFEN-bC_R0E9.6-V[&VB\J2c94B5GBJ@e>PEX?
HeXI9f5.+4DDgS<ceZ]K#egZ[<e;5:2]U:V\1^cQ2ZDLa(E9<]F,#9=_F;).g(<W
LOI+-]>Mcf[f\F39\^]1/ceIZ5&D]S,GE):5ZVTD+=IV?1TSQHTgRL1]^9)R-=&+
VEWA+@DA,KYL\=CFLV>3<ba3a5F^(]KT)\FKbB0a6OK&.&]UeB<0B&f6^3#aG&R\
0PR_>[eE=8T_cPbP7g,LZ1#OKg)XGeN6)5O#-JL3ED/;CUEfE#UP;[A>A;^8&PP3
J^<3Ya3G64^.JF?eBbO7cb4Re+->FLB[HA55\/E[EF@@_NV&E4L]B6S.3S/<X#M1
\O-#bT=@H92#&386G@2_:d?d4.f8]UQ)4.O9VCAR8@4G2C>;Y3)+VJ<H<JAbZT5V
YK#bQAX=C^><D)9T&VWIZQ/)cFVK@gO<8CG)N\L1=2M0YeHR+.<,9g^=#3]P;]53
:<W66E6;:Z4G4]#?Y.B8VDIZdI]1g4UQA.;JS97<<R&4B4CTd3e/eRc#NIB_VVg2
ZaPNg&.^Gg=(=7,1c^:CTE-fE=OK@I2DWOP0()U9,BND>:R4[-WRM&c?eZ/5(]Y\
P,64(IB60a0QEUWZdF2#7(V]_3HQ\?G&XMSU.f<g,A[22?.d+MUD>X:SKa3/S.eO
B#M?\7N^>d9_K.N.YHO_c(Y5UFgPX<BdT#@MC@a\.XZ,Ygaf73SOe?Ff.][PY383
ePDF>VDBF)4I?3ebPIf?a&\UI\0B)?KBL_W3A:9ODAc>1e:Wg/1#W@[+D<2fa6/a
fS1#:c>]H2X-);>e45K54.89^\f\R9YR.TDeV.,?Z6G_Gc=HLN=>[dP)QfgN74PU
7(Z^YX:(.c[7DEO5Ae^?<3gAB^c2PJ&-ROc>OA1Z?.2)(QY-b\/bTVgG5d@e?I+d
Y5J9J4YV.A\)C.C40e4HF]Kc<34[f)I#1Yf7_0SSffIWU@&V0[Rf]J8U]@3]_:@4
H6MR1V@S08X0RU\Y(A78V@3A9f\VBU_-3D17SR;b@H1bH=CEZ(38V5H^cc8=Ud,d
<gQMB]fBdb:S(bF?MP&,gS]ME>.O<6ScH.?fH&T)6.])^=:K;0QSLcHf(H.=FM]J
V3e:f(>C]PcOBL>:g\CB<-KD4MQ\8C0#BfWe?/Q\43(-d]5PW#3g^e)GL@HQ<#Yb
G7AGWaIMT<7\AZIcF<J[3;(K)#caKT@P.R]M<JP75S<,MUARMPC3Aeb9_Ld@P9D?
d-g77M@_1bU#F0/U3Y.M(9VV-=C9g10fHbAcEI(G(I7c@3MB5QJ;@=e1<dYZ3][_
9d,Qd55_1;-M49SN19;\>NVJH0=Ye,N]0Q0+0]ffK)g&#SI1fY:_;JJAV_3&Hd,O
IU54aI95L(A)gQ7S,&-8>#0H1_CNW;2QL@S7Z>J&]<XNX<AGNcI+-(J-=b=<DKX=
-QYM@fL6[07fU)L_#?TBQZ\/02IDSO;RBAa8cP6bS/CSY-PD#K2P&.A2JS9.eYO1
VLI?=@,.[_6#BI.<8/AdeVdT]NR94PTWWC<+=O:C8A,9D-Af05&eASNaW^1X1@W=
BH+(\]/OQ21/>#CAECVdF[e]LN[Lc[/Z7?L#G,M5_[_LHW\#dTDE=6_@GQZ7QZ+5
]P&)B@-2JM4/=cXBQFe8#4E,@S^H[1O)fJ<1Ua&\[C[@cgM]6IOf649YPLBV-PZ0
H(f;g.E3=EYf.;dI._S=,JWXJedE3PP8b,Q?B()Rc-;3f>]O1S>aW>=#P1;c5T6)
<28PDX195/?8K-KPPT#7,W2QL)&/b@f2J\bed0[&BaK5ZcNTGB9270RA07[P-VX\
(M=NS-GH_HED)P.(QIA4-7ZT[_XNfYFF[M_7M25SGY8;JI\O#QR8dgU(8TE8d[H0
8:?FHCWTCXaN&fSCC,WeB8[cF7a-/:_TH<UPf3T3,MZX=g=AWQS1Q1O4BX92CRaF
,Z:W)Wc<++B.KZ9?Y6QP2A.O=C)Bd1U))>YE14M25<S-FP+;EWYPD86)BFOeG@10
04B/JS]M0U[_Ta8a-V_69M2?+PKg66A^H3#Ag-6dV6^D5O_S[5B?/U&He+d@Ga5T
ce)>-a?T.AKW_K#6KAP/AFQG[QOed?e-JE0@C34-c.OO^P9]EZP_8]?gK-;eEIEO
7bP5]Ma\004>0gDT/Q#I_3Fb6aAcOVDW&cWQM_-)Y9d:_@L3Sb&I;:326f911,B8
].#,TO3eT;UF+\)@>QW7#KVAC06Qf-bD[7Eg-O7O=CM?WJY@1M((1SeR8I.U>gFF
V97dE9K.I+V=bC8:#K.5f6OM@47/E-3@UOA#T6+PH,ed/a]E[=>[PP<YS^3([)TH
H2,AV>g5C(G?54_9B=_VNW++BYA@LE-J/=YCf)SZP_I;Y4^XS15\PdP4?f481BZ6
TD:IZf)fA/-/>N\gHINZ1HX4JHP9[\fcE^\ASd181YD3S\88[CaT+_a4H&L[)^EG
6@Z4\O?>4FB@2)F-IJ^,VYWDa0HI?NNCEdTC>.[KDP@+OgG?[NUI]X/_N,3&?4gU
K/2?(@JBRIOM9\aQ=M(@0cWN/6N3]KcZ]?N,BeP+/+B(&?X/9KR:J;UZdO>Y]AYD
Q2I1THHM[SIF.<TVVOaVUgCPS6AMTJMM#XfA2^/80DHS1VMZ9IC1^+ZG]KMg&-TK
?)[:MCX8f?gV4HP9E7E+0>R4J84/Bc5=He&?B\NC\-WT2d(<A>Db@ECgL--ZM(G,
\J>X<>GM?6>715I=-R\b7Y+(cO>aF>6E1Y&f>IMYG02+Z1A7XegLJP>7fL^JSe9[
-0+TH\BbLRMcb0>=HeCV<U_G,_Y3>TdD5PNe#ca.5\cPSCd=R)-LB598>@H^a?Q>
&I?+.XRcBQ0F?3a;eM/_4)E#(/=:C-WZ8O)S;1-dAUOP:dN;X?[>9&:N7TM<E8?_
QK6BESE?5.PWTg2E891e@&TbO@d=#>^F3M,Zc/?bHRVQPdeJ@edS3S-2@)VZQb9:
9I_Q02g7]CY@TG1LZ-XaBdMQE3Xd+ZM2Ab;WI6#IgIIY?#V.\73VaU4)[gD#>W3Q
+3Y6#2_#I+/(A4OT^(e0EST@8e<,PQ[B\a_eAJ@6KDN7>_)Rg;0FIE3aG3(NF7CJ
S^20@/^^C&HcLH@](bULC+^3JOS/AV>-/L;]GS]P<1aK5aEGM;ce#d9I7JH1L+f1
+VbN3K]@/2JX&+V<N]824]dMBYO6\0/-G>b#0Y5M<-38HPRQK^_W5B/KMaH_0YG3
/V._B5Y=c<FX71()]&N2ZQ=L4U7(&7-L7?>-f1K+)VP/)Y#<Z_@YN]f^X4(0V\^:
FGE]@aL_8(?B[SGKHeJ7C9WETIKPaCWAMMY;f_V>Ke9-ABVg#9gA/+\2,^(/AIEZ
4e#AWNANN2#Z@YE)/M_;ZYZ8MFY-&9eWFX\LIMBG>[eCX+gS5@WF&=&60eSZgg?(
eBD)7>N;UZK&ALIPG=?cV&(^\6[2V-[PD3/?[@P&B1Sga-[P,g=7gMPc+^7:N2\P
7Eed)??G__QE5#=>0d([5c2A.K;abATDQ8g<,A:1DT?E8B0_NdC_A@#a+O_Zf;GJ
S-[aAI7[EcgJ6XG6&[CEV<4BKX0NX<9@[He73HV5VWP1fT@eA960J;Db5P[NNI_M
FC,_6<GSb_Y05G3YAXO--7.=5E/WL:D]<RdSaJ5H+]fHU:=#Q7S4=+)d58&:Z_]b
B(O33OVT3B^EYYdHD@,[<IZ3b9=U^_(^GD,fDQ^[^22?7F4U[:,4TN/NSZ=)Me-I
F5fHa-+<#F<NRIL&/;9ZQR#O;CHEK9@fKX^cP_MZNA8fTc0gHT+F_N?@B-a8FH:,
(\CTZ#^W7NGNITf37LN+XEFO7;eXQ01gT2S0Vcf4-_dc_3U3dZSDAU_[cP,1,4@&
MW\9##MR\_Kc73XdAf8X;gb/(L3b:6QHdJ)3c@HWZ]d^7Ra24[+/fV9dQXCB\7&0
RLZ^/KO0O30Z+,+(PD[7E)^Q]BZ:g.a:WT?eTN>DL7TBV?C0^Y2\aESa35G@#W0R
b4Y\-3V-/>)4g(]8X3BW+^W[VG]F]O0APNcB0HP3:BS3V82^TXcdU7KS(]/3T(6d
TR0Qaf2g-]=b,2-?#C6U]ST84IB9P0V/B9GVP9P/(8T6Ff2XfV6^:f11#f+[3F(P
]gDQOBb0U2^GcXGG6d>@B]6Kb06f-IQ_<dTEWG[eKW5a1G]Y=>9X)b3bF:Fd0dQU
+M-__/bZ)3R>4;,,Z00[\F:E&IfY896)#eC[A1T,edcPAFP[WVQ_#g&2SHc;H6#B
JMPREU&00#(cT^HL2RC570V=)Q5-7QcJ\S7KGHNQM&:D?Y]fc7,1-:+RReOYHF/7
ZKN.@BR(>6U1a<=Q=KGgO#T?>X[X@DALKB1S3DS.8IGDU=+U;KVBC^UB=3/S6[f?
Vff-E9^J@/=+M6>ROFZ4:=8d[4?:</\ECBGe;UY;#)A-7g^e&\FL?CJI<NEZ+1af
9fR@4@/5K.,WP]ADDA(XQ-]QKD;<T65FA=ba9O#34K^S^F+XKZ9JZHe2Vg@AVSKH
Kc\aeD/Z)1IZ8(W#M-(cdO9&]a[KN(Z;,<XUHDD2@NZf6.O?E\5--bL,Xa,SW:[+
BXb7F=FZCMQ\]1J30HXPUI^LWc;/A7H9ZH80:&a<UQWQ0JI2D6?T\eXJI]BV/<([
^W(K/eAeF(57UMJ)]GH@EXFX@8dA=L6.c.X:ATbd:9Y)4-d#3E/K&ICE]Je;MM\A
Ff&[KP5ZHCa>fd[e/\3D<0N:8W\#X:8A&<TCY/#M)g)fG@\YNP0TB@2TDSCKFg70
gb)#TGP_5OLFA1aZM24S5FXSJ-KOfDD3=^X&UH_Rc:[6>cS&6-9=/Jg8Lf-C/JQ:
=g]FaMCS4aD@YTM..(B-H6Q_fW#?A[UU6NS?=B.WCCM^@=L=H+ZH_<+X(a/b:?_:
HGI85+RFM4QC/X6FC]Z>&P>2F]U?GcS^<>@J@NKgeg#.:892+Uf=:F..1Z5Q6ZCW
E57Mf:0.VD3QIfAN+/Q0]#89b3_2DV>,^.3>[==5G-U]U@-F>&Tc2S@7/1Id)P(c
1M+aZ7GHc8gTD]>-UR5JdIA#e2f^BTbC\@Y9J4@U6@L-NGcDb_9fO14T]b2D(;LK
CJPO4?bNBEF^fe6#M<+V>0U5dYKAGLBO).Ic5G(M;TX(^KNUHR8MDg]#Y[;3+?F)
BIaFMTT]>1HI(aUKW/)AFdFDaTUU>#RPKCG(1>8c,R92HGY?7T^(Z+c)TfN6Hg:7
b@>5O.0UUYTA43L@C+PEV0T,6=A9]_e:4&_3VIG1Z954BT1DT9R+YV6[8H.Y^;UR
L2;8+ZAU>?YAU5H0a=.@9]KZZ8EYGSce6Q3;,/>A0&:6]>BZ_WS&9-EYH91KL[5W
T>P73Y:KX6Z3/._[a,-K#SDg\HO5Ka=T26)8JE[G#Q1_PKOH7,F@NTaMF6\01dcN
62QDgA#4E7Ka7Lf9\JaBL(S\O:@a0]/A.Wf:)XGC(OL&Rc3W81X9WBI[LS]=0M;b
FQeZD))H_O(64Q,^5d]E^d4>5#MIG=I?KY2d=gIe5Y>5XdW#(4G&RdWBbI<f^5&0
f6)gOa=fW[F+QYcZW6YA9NQg?RW-<_Ede/@Ie<6VTeXbb#&CP^9PBQ_6.^PQEK2g
Q]eRG/J8d>H,KL58_eFAYEZ-1;=(>;.#VL#?7#48[4(W25_XKRBL1:[SBa@>@G4[
WW?g4Ug.a.VHTW0]Le6.e[I6>Df)Y(X1bT5L5>K<bZ#_]GJ(EP.I?^DNL]L_<5D3
/P>4BI=2>T=[3GDR5.c+-]]E-U0(W+V@3#df8I2?I9eK0XJMO?_=6^.8,#=:Kg_/
=dd:;_WJU9W)HDeQZ97,GUP=:?5+,DS^7C;&UeDHNO:CD:cd#e^XIVH[,??U?\fe
148BA^8cQ1C=@A;fFT)S-LEXDI?aDKWa0eIB9=N9&IB<-UKK1a/L;2GL>()]e_db
ZXF\_T.fH@Q.E--4J\<a[?/@1^e0dUY>]-9U&D#gffA1CFJ;QT:40SeP+f^-M8ZM
/KKYg,=1UbZ+V,+[gAT\@P-O@K48\D6d-d7EgQ/a:4@XI;3D9BR&DU+_;IUWPZ1C
>&B_f>-WPC9[BY<?2\Fd=AZOVdI/KdORI7@eE6G(YAaWXQg1]F[7>cR-eAW@1BT#
\@+/[3J3NC&)<.>66FD?,+a(]e>8HJMfS/YaW#Z5Y,b-:590810dC@@1HD2R(QX3
_W7TeC4U-CDMd(SU>\9COUM2EcdIOE5Z?ZG_bN9/^>2M&IDgBTEdQc_U&T9PBQ,@
7J#^P[=TX\,7]BUG,E>:C-9PA__S0b-@WF@2OT@^a8I3gf03&GR3Z,6CMU^@=I]J
WdR:-a-ZJ9W&V5?:HJ?0I#QQ[;c:@5DGVPDA9@WQ-G3VEKD=@0W(b@a:JdaHT5Wg
)UCcK5&?0d_;&E2&6gB6B1GRRIgLS+3P6E?:7b4+0\?_&)H(N0=BB2O+^/]9&SC9
06KD^aU<YI05ccE8_]_G7_-@.:12RSD9:T#(/gV[S>DO^/1:g7HKJLV2&ZVFEA#g
>Z;9..N>?^P5FCALNN6R5,#U>d#N2<7BR6PDP(:-a<,S@Nc,@-+;AAO6J&YN)U=T
gS3eF<J5K<fI(O2)#cM2AQG)M4[:f@V[L<83=O+;(P+O/\bG04.A2M<6eJKb-A3U
JJ9QIN-Z2^cJM-F,P@;33WS&L4-U;M/CIeYNNHD+dL>XQ1[g3RSN6B-RMf?VS66(
</c#U4E)Y[#[FZ/84)ZgMg^88U2YORV_0UH6]^eIfcSZ@c)H;ZffSeW>[M+:e-DO
BPELAG4[?85PVE7=,/-ZK1bNCI[,+F7K0<5FV(A[93@SQ=_f46SIdN[G:)adN-b@
>E;752CGcWfgfXP3BIaJON7Vc2+9R^_66]6-,Z;U.EZ;D:M//LP)+TK1g4V\;CT1
7D#DT0DgaCPPZ950(Z.bUe;;dXe<^P3D1PDMH(\\1^Hbb@]QD,3P3d[A6Y+N:K_>
M=(C>UP?J?[A(?#_V8<7I<I/g8[&2^P2U9XLX\dPY\I_X<W-Q<RK;NKLT66f/L(M
P(-W3cWC0-bDb\Y?X8W@PG0B]9-<YEW<)Jb4W^gJIBQ;eK5U0bODW^99J57?+GB,
O:Q\>ZC6S\\[M<2=_FR:G.b602]KOf@[[W^McX428_c[5>E?.Z.6AX25TSWDAG0f
T?+@L;S+[X[JdZ2@<ZR&][I2UD<V2KF]09&<Y42d\BI^74QW7VLVJR=fE&/IPWT#
7G@0@UCd2A\b@-c;_.TW01:C+<:e32WK@QDN[#]@g&[^2d8IL4#^)bR]+D[;ZMc_
O^cOJ7#d>.5ZPSK0RdQI=E=]VF_EL4D\gGP#US&V6=\9GKbgVebZOb957##);>=P
f1A^E^.c(g^7>D6?WCAb6TGBLT^\dVTFaQTFJ6Gf_=OZcOSSb.G2,Z?bZ0<f<FV4
XVAMQdC,:UMN>fIA[(\5QXV@)a+&cK63<;LK2[2f=WA=_\V95[MTBYY5:P12;EHf
X./W/c+BHIU_1M@VO##DMK(=?UU?aM2+&+cWYJ\\YMc]R+dY6SN>:>S.#)XRY_?1
5,,7WcVf(;a0gD]+5@P/,6SG7;PIH/9aQ,<=.<N.>)d8fJCFA7L[d;2:0<ff@YC[
DC\A\?OK#]4^8I;J]aP^SQb?EQMg)YRaX]ZQge5FE]A]e_P8>@E=DX/&+,.e=6EW
&DeIe5,fUL(SNNfPf=TdV.bF42.3]&6#(JCHfWLU,S/0I6eH9g[KIHA,5KQ&ffb(
bSe:HGTg9,./MDZI)[VG,I,.?OE?J7eT\LO1F=>VW-\XZ5eAX3.>?S)9-:LePOFS
Rg]5H8]_]?PM:+EB>N6WCSOfJc2D+^-NWN?[N886<;T:18Af(:e(:&1[#dE\K-QG
LV8S&,g:UE;+2-VF/IG24)XQ4_/AV==5<gZ((7eR:ea_E0(5XHC<:A>Ab]1:bCLH
A2\6W).6\J]S/M3OF&f97=R.#PM\deIV,Pc0RDf):C5Cd^S]]Z_-,,<:Xb<]RR^&
#]B@5TGb:4JdOF8@&Ecd3W<7)TT/eUS2NV#(>9C_F6aG5^1N(A_CW:BP[gEMWEHS
QZcL/;b.ZH/IdYQIEIbB^ee0@/7cRU2;G\_4)V./AGg7A_XNR_V@fRA6<H@O.93c
Mg@Z^2HLS3J_d^W)H+AEYH[PT1)S6cf>XB]7PYEQ=f@6cH]]4[Q(I7FbLZ&;fS\I
(-Eg_JE-K=NN2R0<fA(?X_dLOZ8,EKeNP^.LR)Ja)TLH6Z(-.F1+QKA[6D_=RY<Q
A.]6KAD^.SM^NeK^K4ULS.;A_U5XR?Te,gSK.3ba#MM[H9f;^-1+3^-&AAI62_c3
<VBfU<@GafMWJ/YC/=V3^HdH3=dX]D,^(1TU5:]<b(0,#cVJ)BdC1?3eCb39Udfg
\E>R2TAB,Z7EgK_28DcKJ?7:UE5e48GI2AeA:]8;:/<-P5UVVS_IU71(6)S<9NP0
5)FM<E/[<aZKD=M.>_g4F(b==Uf,R&aF54H/Y/?HSM]NT70O4dPSW82eAXK91YAH
]7f1JV5_.<LKa0de21IGaCWHIPKdL9R6V<J?G=L,P21/c==4bH^:a,\NLQ,NQ^1S
-b_NCY;&/WKB,>+EYXdTS3)CW>H>6TaWV_1EUY^]d,6+LKa#0O>-Tc#O_FOR>Ef]
SKGcEWf)g/L_P\(\T(XD#T)3V/9FI3M>OaCMY<g4L2>7#LWGT=96<P7GF&<11cg@
#9)R#KDT4K6:[fXX@/cA(^PXEd=6?OI>2-c)#6?87/c^a#N8&I6(??\1f9KY#)T;
=,=NXaR_F_OA<MJM+G_HT][MQe[a2H67a?b-g3cT5V&A-@d>=)N8O_F881?.EDRZ
\5TLgObZ[RPX=UOP=cceQ<KI1d4,-&)N@<cQLd/GJJ8I4\+f727<YeJc/I]>NFX-
fX_X<ET1:cg)QE<WaT=Ke1O0BR_;Mb8ZDgCN_J&IHaVI^;D8^AMP1-@W0e-8E]1J
I+F=LM1gF[CHR6^e54J+?QTKFYD=eK2,<Q)8HV5K=Z3^^28X<NT^4\>382#A[ET&
O;TId^C^YaQ6,K6c2=OL]XOS9ZcME1VZ.g0EH893D&KeJ&;>VV)#<D6@T@#Lg[<T
.NIH)&O:,?;3Wa=+GUD/5Y&R\/,e;K5Qf.CW=WO7K46M56:A[N7T_9APY)bYLZUE
(5W[W,X.BBPZ78L?/dQf#/IS]H:A^>F838AgNI10FSXFJaW]E:[_\1;3MG[I1:Q9
X)S?KA[WQRQ1K-9UN@PeId\dOeZG)E_OGf,8F^a;O@6F?29:[MV(43#JMc;<+PR3
1FI@S]dL6L=VD77Z=g[64P\]g@K>gQ;PL-FQ>2\W1[,UJ]:D:..]RIb5Z@F7ASe?
6_ZS;JFZg8;Yg#Ea]Y7/S74HF;>5S9Y0==BX9R./[4dKTBK=>,.K3REg74<MaM.9
U8-eFbBF(Xd/QB:<+c)&+>,^I>#3-[NJ/S_53f+#R6VA[)?I\J<5SL+(4[<G3:X/
/<Qc<3;/?K3Dc?,I,Z\@3<2S@ffAO]L2<J,HLQSNY]EPV-_2I;3Bcec>D#-L9D8a
.HAB36E_MT-8:C7MO_1:>IB5V9bS/gPZV]UfDSPf\OWV<LB\EK(/.;WaZ9d?E3C^
^=6cK6M;3YUEe>K^[[;M8DS<_Y1-8+5K)KRM_1eD.-R[LD3Ocg0g9bbT:QKJ5L)e
@T?Z@0I)GU;V>,1M3=^_\MVX0>#0g+U6NW.3/X)JOdVC=&13ac_:]:e>RKc645a)
-Q)9@0_fXWLe;Q[=U+)>BfYVcAf+<;=EbBT[&M3^[_40_Z)259F7//<E>XJeAEf&
eb[VCX]1EA\EHEI\)J0a49b-(7J-Qe2U2gVGWLU)eZW)+O9cd4K>-=aDZFI92@(C
:XEM;Q7.4BNWC^9WEN4_2>3ecbGaMGV:M8W;S8J/@6=7NTGEb.8:eL_.6OgBGIO@
(eC-_[>.#K;T)U-;[3AM<P?2)<YPS\,:[?BUW,:;B+[V.O.(O@:6&QFaDD3M<gH6
M:f+[WY91c12J^-?FS_M58?ICGa3QgcI&C0_,-AH22ScQ^-F>N>G6#8=K\6^?\-,
A;@RRbDF86]PU&dSB&,KAZ-LQ0F3.ZB_)Z0EaKY1KBb.&-)43S76I8a\ZdL#VCgZ
A>55A+6I+HAS8<Q8JdTVFFbL+W9>T^b)e2aVBE7UJV]/L+4,)/HegY-bN29_b6#@
YFYJ-D7<UaNN-,WI-e0a+deTBSe.D>3+8>,Y8,,.SJO(N><ML1KL?_^4_dB:9_5=
SEY+,8We09>5<]:KH]Df\IA19#J,1D9f(+FJTQ;7IBJK,F4^VCQD,U3@bRNdO.8;
g-fE#PA_GC9]2-&S+^((@eB=2(-40&dXTR8I9:C@L5bP3?7fdV]&S(L9TJg]JaQ^
SeB\_5K5EYegDQRg#CMJGJQ(YN06O.[N9fJF\6F3=FJ1W]1cDWgDMF1Q+<a21Z@?
P3U/cT83_:)&)GB>eP3#WW2:,f[aBF0YNEVRS1OPIT;LX\AYFKX(M#&<UbPf?+cd
CXF+/U5YDGP^Z]bc=bSQ;MF+aP;eD)U;.f,A+,.<QM;cdL^<XNU,DeVE7bd8E/:1
KZ@F]AA\Y=1.D&>AY\aTRV2^d5Y<^[KO.f]e3T9EKQf-HW_JL#:^>#)ETD56Q^+[
(Q9M.YW39=&L^fVYd0]fKZ1#/F>_8->7H0,J-1?ZgJ/SPZ>.gaHM)GB7Ub,a[#_W
[<4OM0,QT6a5g^P/RVQJ/Z#;gOf?RfLDfDI#KH,b;H:@0&9W5>O==[/RP2g.@AHC
:(P)NgP+5W4SK\+f0V;_&AZc#>Fb[F0YUfRa+AE)fH/R+CFdXW2gHcJDJIaF^6a]
/RF+HH^fYS&@@6]?SV/KDN];^VM0GD;_86NU0X5Z5F>NO2^HOCBV=8<&Q53M6aQ#
)OAS8N+[5G1a^_bHX,F:Z-22KR;eW9KV#GL0/8:D_;?b5G6fU#cW]YeOSM+BJ83<
&,,>8F-=K9UIF?QNgO6FgIITdEM?9G;]Z5<:<VACI4MA4]KXQB&MZHC1U32Ia1Hb
I.K..9.-4Z5ALgOYc4-U=N+c>X1W_[AbAASI:/(PEWbd3ZP4ELR^\93ZZ7Gfg2./
BFN2-A)65[E_=]UN-d>8&K8=NJRFQ0C+e?2egf^)Zf+NAF_1?E93TbVCaQX3[eI4
<0U4];DC1d.Rf;8SL<JTa.1W][=ObA42GA86BCVA1)S\4?.TR3B3&&.KW;VCKD0c
975E\54C8K>9X#0AAa]EOXcJ1^:Z+cJ32L13>(A:=eCSaWHB^;YR-2K0R8Xb@_C?
0e8T;Jba3gc\H7ZWP5WBU_C(^68L>5/_R]X0@KKcK;6INb>6a[&dC#)0Ef8/K=U&
NfK;H;04US3YAW4PB51\),cAKQ,5R]GY[W2LMOZT=?cN?8/.gY/DK-Q/&)?)#HRU
P.Q@;ad#9>8F#cEg(BN>&AOV3;38bVHXG4GJ3.c>=H2Y.7=a75XHH_IL^bL7.c-Q
-YWI_9Q.EB^_T6U?)We;54CQ7,)EPNEgJFP,S)cM\#V41-cW^.aS,C,T,@4-SH0]
f5A\.=,<g[/dRZ;2+W6TSRUQPZOWS->C@F?4cOJVUQ/7D6C8&@Bbf8gHdGDcF7<9
J,65]R&5@PC#HVM8?X77Lg.))BR8I(4_c(YP\8@+4IKR;ZS2bLLEPI+<=@_>Xe/T
&W/^LR6IH:HERdeY-VCN9L\E#Y;.+8<J/\G2N]P,M5f,eZ6(1)];NCSHA6+(Lb\b
7L@^M?&+OBTb]Fa#4X\aV(Q9:=4e3#@^9DYMDTdHX>G@[g7QdPc>R(QNVQ04^Z=F
&OZCU3WM:+^?Fd[eg&5ZIJ;J6@_WPLKL96OP@HTJYN#GN7^=WIg8Ka8#fN,cK8DS
R4,58Cdf/ZfESCH>JV+O&fcVH=J&da^2-0I&68Ob;.?5?g1<.ZSd?]BQ3f[7,D:<
DTIJ>f-f3G1CCO\6XTYF?:[g_L^\V@Pd[<I0S\OZ5P?S@0AgP^37322/Q5?(0Y6C
=_8NS8a5:4EX9T:GK,F]afH-IN3[]8EDeHg/aT73F+/1-c[T;95_XQBXNQFI4P@f
#^4Dc@COg,=\^2Q/QB7bB<KSH+dCXYdA#V6\V0gfI;=\LP=B,53M=;T0KEW4N65H
gU-F6f;9JQKg-E9&Ze=+GKO_.a&1S9=e^^e=F_4fgJP\:/KHAG6NfX@)4;OVCD,/
VLfC28TN44>]Q>a]G<.-OLc,N&F+@<2B?@PK1PU90=;E/.#.+XX#+d.:O)+-M5VO
>MLd=OW1e8M4LWS2DGSEB5Y8S[[9b0C9IJEM;^?WL)J8F&S,]>D85G0W0F+.b,5,
)VST2ZIP@ASaUXbV3+3]ST.-XNGP2+f3UW)PC[V?J;1L-=d\IdUOdLTIfF0<UT=8
+K3dF9.YP<N#YZB28?56^\:]2HC7U>4\#J2,DeI\\C3A/gEaD?V9M7P&=4/&S.08
/Ud9P3RZ:,e,MI5;Db-#Za1OefYFb59dDgYJ-]J]C4,aJTMEFE,/4O.H.&&^>-B:
Q:E=L)^6#/4f:1_0^VI^Vf9Xe8@_DGR&.E5P)=G#@g6eL#e2g4HLU8+_4Q02W<I\
Ub3KO_g_8LWW<5XCTJD?X77==;]2_02fcV&R[\V63C5>#/Id>,2KZ,J7\,69MAMY
@&F\e5:RJP)ZH?>ED41(#RM-4^=,4?N-F@geBI?>bcL]:4(OUdgDHL&X2>?Y.PYL
:;aTY2eV6F=F(A6K8>O0V[2?\IL2Bc2NZD?GbCf/fg3aO?2M3>@@NR)S:3BS4X&.
CUN>,-JPIM1ZQAQVA+2YaeAN#(F6KY6@I/CO(#fGfZc72GeQ4c4?S2.TW1N13fST
g>A[=#COO,dB.]9;)<A[).8<D,5SQI_D<W]#Wg^TeQf<GB)7G]d\LfA>g\T81,0-
:2dZI7]^FP2YX+J;c.E+C/ME\CUFZTN.aC\>3F#Xf]aR1/XMNMF+;U4ZZ3XJa1SM
9B6>M)e=X;fUL._K9XC4:gRf?>:AQcA&fL4+a#Xd/9+O,T?6\[P<DD4.GZ#HAZRR
R&9J>S3CVM5&NM>EHF)UfCd&<SO^gBM:Y3FK6IW8-L2_\dW^0P4-4D[b]f:a7W9F
;3F+?5>cAB5N#gBUB-@HZ&EYDUc^gFH5ZE3ER\P@FW\Y?:T_N383c^f3&5U.7/B;
E4IJUGU4ELeQG\^4.786c8&3G:g-\fb1^MI90\#)UP59H571LRf1()H_OJB?Z3fV
Q#e,:;\A396=<a-I+bA\8LSFWFcBQM:O4WJC?Jd0778CeZFF6AaOPZY.HM6H<^<V
]VHXeWAV2\>Fg]SaLD+>W8-bF,S/)&BX:38QLHCURI^b\7W4Yg4<DD+L7dG@:0^?
8QF(O,Y\_FFNS;=g[-<O6;INA=IT&0BZ<QY#]CF^?58abc\LK&0>7+YUP+Va]AZb
_MLY8Pb3H,TVIDP^VHQg8TN--Ve9(RXd29S33TNU?Q+SV#<cN3bN+Q0Dd]4\@HA(
Ae;K1WN]X9+/>SU3B&be<GaXb9VUdd#3);T6OZ9??-S7Be]9TLL:9STdWEVdIH=T
CE3fL\Uf[98BN&SM@\9XM@Rg)Td.G6DD_HK3bT[W)MXL@/^1O>OCBS#:G4-(I+B0
^T&LDSgD:0>2L-Q:M\\K1c1IcF<Xb+84g_Y[97@YcPN9S(K,EV<K9f+b2]]L\f&X
/(1_0]_gIfX\#XeJXS?Q]5aIQ^eN<fdeRQ#6HD8G<AO+]=be;1XFcPMa)=D6C_KM
7Y.H1DAB?fHC3:fDec5)fV7J1fg@H0b7]Y2F-V1D<L=f;Q8?-W?]b7BQa>DGA/Pf
f.d@;8aH79#OA/O8b,GSe+-Z(g47VaO[FY&IU>GN7CCg:7>-KJ\=T)G\a.G_A0_D
R,:9>gN2A:bF.M=N92R5C#X:.T97NCY?G#0)CI_2>DTb=fP5,->:6a8;+HAU[=98
@Gb3a=.1bTOAeJ\_c17.,5AVgXFHWVBeOD3ZY3<PdI:8FNVadW?BU5(,C1.,0[-]
2<4^0U)JF:L7>T&eKBG4OK&[\cT4PUR/3FQDIeQJ/QgTU:U2Y8ZKHef.VU:I-9?2
;46f]LJP[gW\LcD9=Ta8A7?aQKKaS,#X7MNgHIGE#T+:FW:4IZKW>7R)DgMT_KK8
+4:-M:T)>#4#FQ(=?QBLg,:(EAU?IZFB6ba+d#GY+L@R3(9CYg4S0=)OJ:ER^S12
^5;DQW3U:)HP:/&VV4SF2cZ0U#dLQF].63K,)@T:5<V+1d<=:7L/GAB(R(,:#-&I
NJeEV@T?M?4Pe,F>:CC&RN4gO[CK>;VS8TLK<&,)L[;2ZHb&J8Lg>Cb(QH=4:&Hf
_8U8&M3R#[U@BKECa6?P^GHW13K7Y-P8ZT75#9WXd9J@9AF.R&;V+Qa-Y.=abL=6
a80)DE7E:05-5]A]eM+6G(;c1f3MB3Qg^PfZV30eSC8;eA3HU0ecP[GV(L^>,(&)
[O#)YM4Y3+25^@2.DD0+Y7=;J7P#0[Wg7[1^9EP4Id;C_,+LDJaT58>NfWaRN2(+
D@+d<>2:U7ReQ4WGB8c^=):(8fFV0YGeEaX&+adJA(B1PM@-TNgL,6OR#4I-d@M7
:7B29Q?[RF]YNAO]Md0]-dMR?Y9-7=Pe<eDJ<O5g^3XCGeCR;@T(2:(H;G)U;7;(
HU:&,5=1NT]Q;WA,]d_).3#,7OIQZL0K\R@^[W-AGe&^N9T>XXU>7RF5UAfWIDC]
=1_E.=@3KTT>,HY&Ja6WQFeJ.a,WD&PYN;AHE9Q0J+1Q(X>GeFEG#NeA:7f_d[FJ
_9(YL8Yf?&/f2eO/4@[?ENg&C)02KLVJQ#^8\b8D3<FRF>CK^#&e)Ce)&@9OR^>&
]FT?2CRG1^bM<6H934b[->9EG]XI4FN=L?Lc?JLXY[?b@CZ\V_E6M3aQE6\E#>Zg
fc;=WJRGVf6Bg.e&>:YbBMV1A-Bf)WO?PL4b>KEf_#0>TcaIIK_HYD(@=:cXR8+=
61^HOG_d6CI#6G\/GLMa#@P[eV,FY1+0;T-bVOQUH&:Jbb0e6[I(=94_K@+KEN5J
fOM4[SRC#A9G38J=^JBbH[LO2S)&O1_2W=M9Y7CV1gM\I_d]LfFD,YU\d@9QB)E[
DZ70M>gb8.@50&@#[+VLCf3SDF&3R32G:T]9MPfU5)\<[&(K(Ob3N?L:[M4W5AD1
3T0CQ;Vf@.4[><I[UY?@[J]IgL0eKKPeEBL:5DVNT)XLW)g_<PF&Q,gK6QB=g)Kc
U[,ZKD,+BNEJGXJR-/CWQgeP<LF5-VOf,GK8OR7?Pbb2C/6#N[,[L0BLbR2[7g&M
a-+GRb65I9M6YP&)(/TO->4G\-Y#PPJLRIBDDY]SP70KPEZ//\a3f<UFS]Y-\fgG
[8?].ZbAL<6VLdM1FA2g0C?A2#X[T@-G:SLYHR<)UH(#FbI=2Q@&25?a1^eS>>ZO
4UJGX2DXRLE9<.T\?_9]W(_Z:&,DU@NObXTg28OE:&RH;Y;,]7+MY<RdPP7C1:RD
/aI)Y_&X&88Q_;QYGVe4,ZAO00;EOa-/d(G-VTY)95NVU\DH:_-W?QS41V1ONd.C
+\Q5G1<DI3a;S&c0?P?:ABNXJ@7b+ZMC.0M]]?cUaT>-9[]UC9FfH7#^R1)f<K^g
QC5,3&LeI7SL1.MD6-31C.&8<GgGE_4O;8L@&:>,PID/X.H+c6;^Jdb]2?7H0>6U
G-0KgM],=B/R94S7@ZZJJJ?)V;_<Na;[M6H38;DE@-B<H.RG21Id(/,B&IA0B0cQ
JIG\]-=3ObM/A^D9LL:OWUb:94@a=?2R8_&KBZB#/E)8fP7E;7;U(T;Igc6BDWZB
6?&.g)JM#)QFb3C<+<#fMUA]&6P]W&?R@faZ^S)E2BV.dMF<A2Z,,,US4QZgf^M.
H1bU,=:7<T#3(:TA6?<dHa)7e,GHC6cK2=VW:BK.BeH552Vd[[,X1)g<2Y[c\965
CHO,92L.S4^WO9EgROJ>a9^[,D(PM6Q5:AZACFW1ag^Q?><MZ0e\H&_c-M[c>-5T
)LLHV2J:34T+Z5,K\MB4MTF#.8VGJT=<L+=3VGc,5Na33Y,8LSL2a^KDW:S.@aef
7IX>UL,I[U.KQa5>=.BG+Q-RZ4W:UL>HX_g)92^dS&IXefX@TUT?^4MQYb<7E:RC
\c>dA<Da62K=N)-L\K)Q^-EB6#APTTbGR.M6>XG-5T&#:HH5KM9aGe/LEM3e326&
/gAa+F)SOQFB1Hc5+[,+W-[TaNC7X3K@S3)\\\(a+8-5SfW9JZ22UXAg6(1&(7:c
,4/AC2V/W3YAOBGX>N+++2-+E#Ea:FE@4gELYBfD,<a_4TdKZf1C&Q6:dL[,MXVg
PX9./GVRY=D:BD+Ge./NQ<>0<=a(2-_g8dZGcAIMD9ffSI#G)CE?LIU61?+XabM^
][cAJ-D^[J4LCL7IOaE4L>)1OFDH,1KLQUX:>g/4>;FMR;<&ARR=FO3R7.9BOcV_
.6(8d_BKa8#:)AdTa\5a@A=J\;5-9g]QXHY6_<1BWVIdLBU@2IIHNNBR-.Y=eJ+&
?7:4#Ze2>7g_;GF0E]D0;#64E10;7X:-&ggN[\DBYU9;_fARRYN/7e3Y:&G6;BHC
DQ8d#HN@ObJ\.Q[V1IZggR+/g91U[-6_S?8I-6e4UJ2e2TP,M.E3I\RK4A1C<(XU
4U)@3aVI-N2<\>a&LUdaI<@0727LKMW9ITQEfgW]R?g+.\WH?e>LP_85E^^HA[K+
S0=XCRB&ebNE5eNQ=I.;#\ST0;07<&>.\T?\JW[]HfELHR+OWB=b\:5#LEN0)?@@
=UEfaI?B<CRN0&>C3WU6IWO)-,(50&#ADa,NDH^MR2JacaT6NJUUNUGe1AcMad(<
6L-@GLdALUD2=#FIP3YH14RA01I4O1T4W.;e[2>_0Z7]^B)>.M)^V(#@M4H?2V33
4XUSZZ=6?1(+\5<FPTId(FVZJ/fDHQ0\@29C3f:-g->C.0MGHfME.6)(R[MHU&P]
=34JdgQDRJ7G71R7.b[:<ZS,1#W7+33?/PUW#SCY0#QRKcdMW>4a8FUe_@DeXYO_
T&/3(XL745O1cPROgbdG\^gB5H;;(T?g<OD5RaP-CILAT8M.CJ,(>LVE3U7_GL/9
9:B=5SLLWg&Y(U]H3:2?L:DEV<W)\B<N6#8I1RO55KKGS<KcgMdMTX522?M\;\AZ
?8]-E(]7>B\_Z0b+MSg5#(-RF:.6;5;\MXA=aO_ZcUAd1J0cHa,SQ.:Aa^Q^.GO9
Q#;#2@bR;6W>;VO0F;4IPN_9MHK#[AYXR=gfHK(RaKR(a93-#4f7&?;&VF&9cL+=
J6gT3\;5c525&>8TA.8gDHbd.J(QEUUNQ8B=8ABV/dV2V4@_.A;H53WcIaXeM)HL
IIB?C;ZH.TKH:LTcY2fAQNT&_^@J>+@1X0Y8.Sc?^a#e=Fc+52(C<@5Zf?<<@RN^
JMaa?^GB+B#TL^b0W[&/E^MgMVAY^P;\YK:I2&I#S<H8<E;)+g.F)NB+-O#^78W_
PFWcS<P]YbTLgDZ_3T=/@BBV2]+9Y_C;V(T&?0DH6K]@RKI]5(<R&ORBFZY+Ec]F
IU9E)5WWHXYAHa2VSB3B#?O;QfEQF?QOFbHJGDQK&g3U1e+QU;&(EY<7WdP^UM/:
3g3(=/aH_F<FRZD3f-2#La7YOGZ8.YG<b/LZ_T-Q3-U<1,Zbc)R[Z.&EagV+:SNY
QDGbRI0CRAKBGA8FJ2T6@5R8J-31ZOMM+&<6IIA/c6)GA;HSSB09Z]<3MD.31IcM
8&g\O5I05>_M>WdA8+&FO2Z[)1YD(bO^0VgeO/(UJZLM?Z[<.IDMA,?B58U3K-K8
Ec52U^Q2@aMARaI.feYF1;F1F:RE^PdT9dfFFa]Fc<.D<LPC12.QLTAE7:NZ7(;.
YC&eWX]9<HS)5H20Q7TcL[F6V5314H-@g58fgTK)8gST\g#V(3+]GJW7fNLYX^/]
S6K-d\c_W^YSOGC]T&V6GfgF7^/#65]R>C0YAD3RY1RgK6\c/HN::0d8<LTbR[\V
:RW0H#\6M[fQEd-43YaZgA/MPcK@>-Sb/?B@B?C#[dA0YQCI\DYSIe;QFaRJ=/.8
2,g9+4L^g28FJS]WBPXCQNd2XD#V2N8D4-VG02CgZ;^M?J<RP+>XfZ\)J;S#RX6D
:6K[X(&@ZK0bWGb))Z-?BgfZ?I#:N#E8_\MW\[@aFbaJ)W_F.U9&&ad63/;Y:?d8
>L]GV#\[QM.<W8FGQI\IC2JKZ<-CT\ggMHRJGG>gT\+0OOX=#aNY@C::,86-<H]a
0>)O,]=&2g],TZeH#T.f^2)-R7^?b/36S/S.J68?(;<@@^4#^];Ab@be2fM2]/52
?KO.C=JOgc<EMV8OG-TWWD4A@),Q7L\g]7[.\G:D:YH(5]fOH=.L/a@\7\4LLO9[
LdaE6_U\^MH:_e1L;a,g#SKGNg=B[P126E1QL5.fPL)U\gTIVg2-KS8A,;&??S/N
J@0:Q:-E>9BR9#442\+S.1;)gD[NJaMEE^^5SE4G.RS]WVUL;6@_^XL#Edg=O6K<
\J)=g(ZAd?ZWJ9G02KOD^P-XVUN.)8#aHV)J-b+Kb(@AHT#A9FKeHU:0=T_5a6N@
TUWT9>bbWL7\I2g:1_G^A[C96M,Qb<[YNgY(9Hf.;G7J<bWH]/(Y86+?QD&/g-&V
N>6cYU&]Z0H6=a_TaQ5d7.@V\&)8,2J)?YH?,PLeT9cf2ZNY@_T;H/@J:UX^9+g+
gIQO&-C?Q_(W/F@^:\.(>\g(7]0;C+DV@]J:1]bB1+GgLMLB\8;?;IA:?b8I8)^4
@SR]gM3d2Ub1BAYVeJ7_Q(3DaH&fX[&:<BeSS[7[T.(T626T@f)cWM]H>LPc@d[)
W(]5Z(aLV4;I]EH7e6O>+Q9KKCBC46c0_#gI8.a6&7;L7L97NO3cg6b&21R-d#]S
Z:_N9CNVCaF^#-6Q+VX;>[c=gCd-\[:,Cfd+_?OgC.+:d-:ZG,,@N:588-fO;PP&
2O8L1N_,3Y7_LbI,(DU+0]DW7/A).1AN#PBV7;g[38T2J@,4]C;-fX57\b>U),a/
/01^]]J)HD[8cdIc:/?9-dfaD3]XO^dW+/_QbU^=_71e?0_+EJQ4ZHF7HBQf>&:W
cXRGcJIINPZMNfILL>SYdSJE)-2+2//BQE,:@<f^C#<g3E<16NLNDc8bJ,+R/-WR
YBXbF7c&/&R\I31Le12;1G6YW#(^AF09VEa>+,^e.AMe18FNK\2XPb3N-QQF[^Ra
>L-V+D::7T1W0ZIQg)?ID_=I\Sa#CH-F(Jg.+^=JS59R<;e=a2a;.OHM#?4CDWKA
0FdAYDIPO(@cWaBK=;]0T>_WN@XIa-_<e7FQSNF3E9g7B2I5V1?<J:>HIS:\<^-C
-d[#c:<K@1_7Y[8P1M\MMf.,/(T>D#8D0F>;XYY3XZfFI\]A?FE>)c.VU##MCa,2
)A:81H=C4CYIZPIWY8_M>@S#c=,H=bPLb=I3:875O3M?N0H?.X4QD<4+G>T=P]W@
4S2NgQRW8-+c:WT5b(QRH7+,O<=Q?N4#_OO^8P)\5GQ^U>+:HMfDL/_HVc0&WVDg
=LG^7IVfP?5B<7SYB^+7/&@J\0d_GXD34HXHAd+N)Ne56EC0IB]D7PbN(F)Ie/6N
&-UgY\Zd50[Ng#H0\f[&@eM_WIga,X\U0E\APf6;PeW46,WDW)?fFbFRG.;gOOa2
XcfL4\@)XXdcUUIbI.X2\d=0O<T7JHA7))CP9<L;A1=ZZd<9Q5d5Y6)SS+>;A^WV
J;6bHUFRX9Wd8?61?=CNLW)4Q\f8THM.BO5HH;W=8_PA8HNe;)1Z&a\.L)Vg[83O
cCXcL9-2://1UBQ_dN#9c<eK_#[;61b:MC1gGETEFSM.M<B_;Qb4:d51#)EI/g9@
.L]..3]e6?EWbO56X?HE5DP21H;g?+S1F5XCL]4Lc8G(g+NOHI(,TN^=:5C8ZV=0
8@&3:EMP5+;gXeO,J1>NMD8&68NT<9U3JLKeD65)+V/B?gK8(KV3^DZ[R2?@YP)A
R3+cfUcfIf,KKA_VKNgLQL\UD+^=>).5Z#Sc.L5Xca?9JV\cA<Z8-6d0LPW,\FS@
N4C:[NKcUB0P[^1G2c12D/E#YN0+&Pb[CLFWF.=2P/U)5<3#9dS.FZ.ZO[:XJg>\
JN,R#:.JHRL:e?9@d.QPC0=BfLNY#Yb,LBJ7+<_>IFF(JW_Hb3.IcY.dKDgTHDG>
>,N>+_g+d5b4d[E)KW36F6JPN6a3<Vg.\KWgW4FS7[A>MJI1&Rd55T76\#FO;\SI
H)8&&8VW4:#.U+/6O.XZcb>RMT&#/4\,HfQX3A8c/CSa<P&HF5WC0;#4\T2C_4=?
?)e]c,XQfgL(DaBGfCUgf(;EEfPDQeLbM)1M@d/4Ue05#B)4VY_7b4XNaNA<#AYI
Uf+7ce^IE)4\+Z@C\J,HK1KbHYY(0e0(B^Y#dYNJaeBM.>Te,=#T4I>FF\[eA6CC
9+9B>(F\Rb]AKYQc#L/&J3B._H0Xg7b]86->-Q^G@]\CVKOaGbGZ18ba@JV4VR[Z
RV6c@9ggQg>JR2?PLeF>-6B;IS3]d@WZY><3Ag6QY:+HYGA;^;I=A/AC2fd^14Qf
GFaR@d.YNKE(g/9&Dc&4KN8eK1KN+#0gPd1CMS;Z-S71BI9_a/f?G.A^K,WXf-?_
Re58a)g3(LHOCY:<O#V)C33e+.>MEe47S8FE[e;ZHOW^<fNb/eFa;:@B:V2W8CFM
NY.O@f.ZI..]#dZ>0AUbXHg;FGTPg6R;GOS92UM4eVV^be1GY8@6;M^97GKJU((9
:&>5HF9N?)Ob35L=<dc]OIKPUXA^<>370@,3CgD#1Of_D)f-Y[TgV8GV]E&#N)Uc
CQ+Y?_>P7)bL1;O\),>G(f/JeRJUa941H.X//249]#@8f.X4P9SE)B1NWZ<^>-G^
:+/Je00_I=]#IC,_O^NACD?BG+5?KLMK,8fRV082g@1P0\V+E@)b\67KGPfJB&@A
F1#G,8WNfIT;+,DdKS@<QUD7Sc3UC?DTY\B)30>QOMfC7BQ=2Y[#^B8>,NI^>dE\
+W.UYW,/BVa,G46a,a,3(O())Le]ABZLfVP=+E.OZbQUe5Z9FGb)_W,#9OD50A77
/X(]HB,b]__a9>Q&TDVCOT8&<0Z[AZ1J51@SX+KSG]eC87dCS-Ad@T0PFG@6ePMd
EQ&:U(\J#EQc6)F))Zb9_gNfH#?&:[62C3>?d>38IW]aY6<c/WKP48DS9&@HS8f+
d&?6YcCac6d69>8Z^2=(QQ.C(VAcT7DBH-2YYCKSFZJa/Yfe9<\<QL\c+QX>P.&J
^VT]N[IQBPUMA+^6PANd>AHd:UB&&f9_@(P:R?1b(//638@BJPL\3N2-0(7I3PD6
S^]BV9f@\]XD66fN#-XT4KJ:N+&MGPUI24JQKWC#6L9/B^8eC,IK1eVTNb&^X4L8
?U\Dfb/N79GCA^c2-#b_324;0.VY;YcWH>-(+BR/6ZPfTB5EDf^5#GXCJJ)Q(&.U
cL7@+fb<DEN&Y_;O,ZeLc7OF42I]YVWCSI,;fA[.d7T\gPIZN(:a>&X6e&_0>E&b
I0\3Yg:6#G#H,#QJU[/H<EXLggXL<ND>_((g@cP@JWX6X:2R]BLXY3LDO/,C,DZT
6W^Q9/QIOQ7PW2Y4<3)9[<#?Dc/_X:T-2\)YT(K&Y^P4H&K>--,.PSK.JfQ<8/W\
ZXHb<](+M\R^?QE30PRX+71OKc;W<6G?V?+NLH.E?2X73B;@OL9#IeU9XgLK(5;2
Z]I>6M#==G)[AT]c.?Fa/9]\aE[VDbWK2dg=FdS,eS_NfYU+ARCg0R;STDJPa<M9
-&Q-LF450[>92H(YCMU2cZZQc\\Tg4?[AUU=DYAS<E&/251L93[J:EaKS=QWTRHY
/J2VMKC[[XgTH(E+/7KGSS(YTDY[EUgH0cMA[:cbE/X^G#3(?9B/922\VS-,8cd2
F@dWLdB4YT&6L81UH[ggE#gP;2N#d2/ZFR1#3)L>WcQe\GS-aK/>D?5+PT3PX(d(
gT=DDNGS1W/EW;dcBM\&Yf1QWOU#VUWbJ+9SL18+Q?;5[E+2c2+;G-G^)_b_7VFY
b9R.-(H;F4LB_0--R8\YL&/Y?)JC.Z)ZN3a5a<b(5ZH@1Z4McBFTC-6GdH<R-dY>
73FWJ:N9T?P2c5^@d/Fcac<XBaJedTb6aV-6\/U;^L>I/5G24gURgWWZ:P9R4ND6
ObYAcAVcCRLPL[#_=L?]eF?88beH,>R([5b^30O=Nc=aI<S(1>@7(,b0@G+@.I@2
]a<J)P&-WdMG0LJT[9g7_>GQ=UFM/f<>U=CAb1ODOG@d/OaEO5;FE.,#+/R]F&R^
LVE4aS@4YC>f2A:=E[XO3AMcOPY4U^7/&WRV@2PX(LYPXWf_&[E:I+ORIS=H<.2&
0QaXRT9gVK@4ACf3A^/<-eY=1A-]#?I+KKSPNZ+/L-GF,eD&FZ#0@1R(VX@C59U3
G1eW1J0ZEeXbW./\CV9RAdc7VP7f\.dK[[=CF;?PN?D..06NdNeKS&GQ,SS.53F/
2Z;NX]gMOJ;GeDKfHN@WQW11KT-<Ug/@_JMS6)eg&f=2Ca8F3.GE?Id<X6/<G-WT
8gZ#TB:Zg=[0(VIGeYa2gd(M&=+fgVL/5DDL74>11=YPd7B8E_[R,c8Kd?7=3>c8
N[Nde9/W=I/[&VDXX[;)]0SCf[d+N(/eF.E1LR^9/(6:N5^^MUeY@K;=TZ?_1f&8
]=]f_;(1F\^dN/eVabDIU_D7bZ:(Y]fP5+4LVBZR59GTN7Na.UAR3?aSL8]P^KFL
^V+KK?&R529S4,6;YJdcaK#(/2M6067SC;[QYSSVOPB#7fO820X:N,+XXONN;+_f
;4RRHTaEM]Y\SG>A#U83T5L>D8N7c3>C8O:(3.G1a(WK39c;^eeM+dfBB.75I8HB
SO#aV9B]^)1M_3(8dP@[(^RIGXW=N-JK&WM:aT3DAQI/Q#O#-FeX:gXYW])&.aUW
.-0K<EI5/H:[A[+8,DD//Ha^1gO]O3g;H@f=bYE[=:FX\,]E.=12Z2LL,5ZT&J/A
>ZETeP7CY1CHMHW2,W)(HR/bKQ1TBAgCGd83[B+S\.])WPF)bYL1[97+5K/6gE->
BG(>_I^=_JC[;<#4_fK+K,X(.WV8CB;1N7TZ?.L1Gb_f(?\^.3?5f(G0LN=/7CP8
S4aKSdR]\\\]D=Hb;(K9]7U3gT+;3-)TTMS4[7(_MGH>#OCT4&2?OD8/N]>@O;W#
>QG=eI\O0c8.MCLAONZHdUZe46RGYRb,X8f])0bQ0=2TJ1R4Jb5[UHGR.^QbN:6<
B5;JOJ,.P=+.,8J_7C:eMYC4cWI1Gfg7:SeF]CY<Y#&>9\S;\^+N>dO>#QCK]T_Y
E\<T]6SPg.=J344Q[6GQB9R)\E[G.d#UY9:^CG9&_LQg8H;+g:K#SO[72N@TQ[C=
R0[?+NIQC5d?5(A#)BHVM)T_.X-:YgFA=Nf=G12C)Zbg--6E8PWBTYbOeC#I1]J8
TNEX3)X@5X;fCZ#B]f/[0-2d?@6HQ@42S#e9N4fWeY/DAb\698c.?EE\aVQ[S,R]
SBF12g^B(eP[AbFUUcB]U&/O,/[#=J4g8)/BV34A+Y)&IM<T<<4AZ<^NOe_2?M-S
F.OUJKI?DAANSP2X,<(DK(g&4Ja/-Z]@FQ.\\TIG/4Y_U]N2JUQXL6@QH-M)7@-Q
P?_LbX.L/\Z0;TY<;5#e(6c#EXU.KS3F=^K(84((\dcJ<gH2LS[HX:F+=Df?HOfP
P,T,=ZV3<,-1+H6Tg9ZW-W^<;d<[JN\83cY)0dP#[32V8]IMA2W/R19-a3&=B3^d
+d5#LRd:b(B:A[&S6)Ta]-,:X+VJS,4T:D8&>eUMY]:Q=R3)JegfGN.8X_.NfgaT
(EN=_#bY<23d<b^KCO3W1U<;D#<B4#91?@;8ZGb)DERC]Og5GE.#Ka@HZ.7##27Y
&J97T]>9NDJ1I,d:FTH^d8PBP,/[dGYZeF^D=I=VMegK<f-(a4B,b,W&<?ZF)9(6
)G2S?_N_c.EDaddSee@U:N61g^eK2EXPKC;e?BV90.\A4B&@K321\NE9g4TR?:PY
4T^#@VNbUDXY_O_R\90VSZ49)b9g;Q470696+RU1^[(cK>,g8\aU<<1Mg3e60LQe
IG,5Y)VVA-eZ\]6])?3&LX2JTO4750Z(e_?\Hd<.#62#Y^g\_/a)#[DET/4.^(]J
6=K>R6)BQ2^9K#J@TPNC(/JdH9]D-C(<CbF@B)?]T=L_(J;MT?10Vd+<U>>=F2WZ
Z=-?Q<LF6K;(:e[#B@5<:-/X6VXM<=T^Z@GM9NI<LeVV//=OS\I1:JO-OFUE+H3D
GE^CfMGO3=<V<?H>Eg:FAQgfH#:BK8AbK8ag1-82WAA4]<>-F]_3cOC&M4Q&(b[W
QN-8CQQe9f+NS0@V5U_2#8-2]?Q@Ad@-;ce1X\RT.>K1YSVHU92)[AI6d3^5e8JN
I^;SgDa1Sd^OdDBJ#dW/e)X?&LC;8bdOKQ#_PYT=B<C>e8@-LgJO\0.2-g2J-,9:
>Y/>AD)K\A_)+eeBeV;[GSB3(;1ZgdZ6KZX&2+.a=[g27\_1C/4cG&]UDEYR_&_O
1_N7CKSF4:gKfP<1dL^>0+c3XdR2CP(G(08D8VCIA<>RUV0aO)b<\=1[^4((9SGW
TT-=e/U5A<_c,71dc19+UM6B[9Z&C-OI8Id9fS5K5KF-#U[M9N.FFb/T:(R,;]58
KD)>2@K1C<XJ>a>[SDI&6)4WfIDER1]U[S^HG22O>#91a]JRE((Yfa\^2FB?GaM9
=DJdP1\Z72+S<&;#Y\@bXPfP+TLgPXH(ISD<A[CK]\;X]eB]a-.2X+;3UF0EF^K-
LX8@E3<H1X(:8X62Le[4DWR_>QV9Y5J5#GB)eGDbN>VZB1XT-@dPSIZ2_DZ00J61
C>9--a_/M5G^KK_]RVSF7;P0ZA^:WVO0?L/W9Zb.eV9fF2^S7I_11#f9B+/LfGPA
d_:W1/;SE\L&d:c<49aG]dKE,-8IUQ^_KfNP,/@SWN2[/YRU6D\?SYGc4/5WER:/
aUM#TT3CH33fOUeJ-gcXS=/<c#Rb/c]f(8SG9J?,U,[VF&72b0W+?7#fU;B\4(P0
ZY)N>ODSTK,BS]QP(JTFE[8@<U8_/W&#;]PBdO.HOHKeW0F1(U:4.3)VUK=><#:2
f(15cdT&B+E?A-UMKORF_E<2J7TGZL<>4]^Ff_8;+>IZIKX3,S\QEBN(cVE_ND@-
Q)V]I7[GNc.#LCSIP@#3;D&F/>:L-5,)IF(WaULP.N9+Z,T)]=:eeON,D2GbWefS
X?X7+GLQ.Y9M^#A6S2N/CQ?8VI4CAL2]D)#eN^Q\D5OY8a8AfX9=DTLE;YHg=Q-O
J7;LA@<J2+&I7A=I/#K2<OcHg;FC@Yc(VcJ7(XWBF]<D7e;LRNU<aB5SZLQ2e2LU
W-=(5[BG/eM.@g)BE4=@g5D_RN/J_4Jg@cbL84a7NP6dGNQX]O=[e(EJ&RS((D(M
C\3:7/,KeO@V4,X/-RI731LH2IWK-W_MNI0gd.bV_2[#/a:W,>_gN<AFGVY;OCN=
12WgX;A<MUWH2)RR/S:9I5UGM+;\HDRX3NQ23F9RM9E[UE8OP5SH<N]?.f#9]Y.>
bLfc[.A<]F>7Kd[dFg+(5\HdO]:UELb/1T#W0(9HaKZ4dG)Y5SJT[)+D_R@0d.CW
AX8Z4A@M\MAH1\7+OAf2fYcW^EaO27@8/)&\Q4_J.f3IL<+dd=L=d:,\XNcB2,#.
6?O>M27VaaNa::9CXW-01.^eG)WHIF/dRF-HFBR-S5gQF]/V5BfD(]>::#>aaUO)
/6^CN[Nc9UagG^&U)?)a;T7F:RPK/ee]fcd#>37dB1XT]#3&IY@5Y[LG7eDFa0JF
(>V\@ePAE3_WV+AA5Q.+KXM-+6,DU0.gQL)D;S@g[73UCdgGMGdP/D??J/^==(B/
Ad0:F.3A#=IKD3XO\PE.0aG]PAeZ794SG:.=>SV/B9NfG_\Qg8:/._#?M5R&D<.J
1T=fG(KeOPc_+)Y1PQ8^Xb\C1Y/aMLd/AS0d)gg5/FLg88LDOJWP,Q#aFM\Z,-A&
#J#7c,&Egg@Ue\+2d5E-f\\[SacC)?NJ]YDDe&\HB+3,F6PN732T@@,42&)5KN<O
WCI:\Q44dFGD<RH,XNVLU>V&AZ:PF=Q;\Qd?.MZ4004fKN(83T<^KYN@&N]bOY+-
P)(VRDbTK[G[K>)XDE_E7-CeQ>;/S3dQD?a^3GP)B--b)eU04SZ1Of9HKDSY@085
&QIVM@f\aAT=a,CLE.3SeEZ;7H1.V\(<V>E0c[faM5-N5aF&T]W2MRgBMd(]5@H6
(@?8&;-Da.FaZDL;4S&FdW;OBK?B9KF_eHeXKWS+),?6/gTA-=3U8-d:QN<aAK0D
X:c<d)G]Z<?Q62>-4TA/YFc7GHaWPYV7JU?XH^J4J.FbK3eFFdfPXdR7\(WcV=,\
3QX8-P6E\1-F(9VbFVD]1FQ]17a=P4^>3SWd@WgZV3>Q]+UO808YX,]fWYB0:(A/
Vg1e(3?47^0,>eQa[fG^;ZbEg9\1FPJ1B2OcaGV^5-f4EGNc+fPZ8M^(?^\)>=3O
P\FT-</XMBbI&b(X]_?1Gf\Oe[()3KD\E8fBX:,[XcOD<O/<E4GRA\80d;H<NKM,
fCI0C::R]]Z,[5QggHJ<ZKc@]O8]2(+JN82G5\#.FD>Qc/)@A3015.[_^JEc,3Jb
:@B9C1a5WDTXRK;.EP@NdE))4R+0Ne=bOSc>>gfda&:4,/#278W)DcK_>YUOAXb2
_U+LW:LZFEQTe6&G4I5/_bN@eeRdW940cVG,WU6\3G)g6INa3?_fA8-AR/&1W^ZU
AJU<^.fBIVZ/eYbWD;N\GY.=0TfIJK/CI1YU1X@>/NQL9AZ#Ee)]A6KQ>=:B=57D
1Q/0DE5(]XLQVF7(<;3_;Qe,6PbI]E9-^BC8,g>,]A:(^P>)]P4bYB)#,C=,4^\0
86SD&@dM_-a9A6K:-8.=TdAgS.S]E,A:;9IYcET781<[9ZAcQ:FO+[+a@4b46TS+
2@HgTcPU#:D/3(&TN++F4\gLL;^K\JG1G<.O-aTM]D@8S;.\-A^2PCPXLAJCSYUa
8BW^#MVF.J)Nb^bOcQ?T)W],K,9,PXcHE5Ia?3B82M6.0#U;@?]d36KDZ9Z6669<
]7Nb.]B9U\,FA3+71U6::KB15?E#J&43=0d&KVHP2#6+)LDVJaW.c/eR.[d?D4/]
g(VP0B@NN1G@f?9]a5;H:,)PBU[3BZ<<HW@8cc&Jc6=+e=LNPT:AW6\[Tf0-B/:(
bd]=C<T@HDN3Ha86S=O9:D/M[b:4N3:HZ5?JU(d:2R&A0RLSe>\_OX8_BM]caLI2
<(&+?A]9H[VdfbeZJ8d<V:aY)EN.2B(Z/=2CD]EY;11\UEKG,-7SA\O#(WOHSTLY
S3cB/#X8/;EFM0H1:ANIR+1-ZFc&BcH739\>)6NALB4BDXD^aWW<4(.,f:M93dc_
[bO)1TO_b-W#?,_NIggW_\@+2RWFfJJ+0Z8A&0ZD1G?Yc4P0V:F#/=6QDUaC(0;Q
WI4g7gTdO]Dg\PWYI]^XI?B&=(BIHJFDB3LX./N-:_@M[HKB@-b:6-0DM5&fW\E^
UGCHO.MX\5-D8_KW<U9O.DSRcgXgK@N:UB#IC6bW;J6\EcDa/A/_577[J=LEcFc[
S:#2\])F.A#78Af<.T9,J)8O.JP+2e<6A_8H3:6c5)T>_[@_]b5&P&IVQ.T14CgA
O@[&L@L<Y4->25<]0\:]KC/^_N1@Ma;6f^]0<8@5Be))W5FIT2NQ>-WA[d.<6MIU
.6-MVS][b4R/eIKHQC+],d)CAaQTIGNJJ)aK,:<I?2)P6bQFJ[^INY9(JF,<F7IN
M.]C;SNV,V@@G&9-+^U>fJWA=&&e\+BV)H#UM0d#L95II,A&EF3.S9/CMcMA0eH@
G/X_ZVO86]Y09,Xe\\0A(S#;Wc:C2^#_?3e..U>Y07a?]Q:2eH<1bZOO2_3.\1FS
6K?>?B-<.[+c]DNVHbbY(;Z<?/>c^e.cbA:D=/32D:DRAcK>_6fNT-LX;)N0STGJ
b0I]DGWEd=9>+f[3>S&d9b93\)T.Jg@-=/B;F1]S:e>U>O:F]\?Q:AIU7a45;C^5
Z;V^?[fLO<#TfF@]GPAS?W+9-M&QFB(HL3XQV5E?2S))@COL@TOM=P3WTQ](ARO\
0b\8fA\0bTX-UJJ0f/NPBTCB6Y;@5S)bIKc_OI0Vg:-T&GFL^4<eO<^XNg=K.EO6
C9b:NV.WV#T_IdIA3&4ETTIM>(OY9++]KYJDAL+TT@=MSb\?P(eV1J-EU=1TFJKN
B(@aPZ.:K)MZ8X)((]HAR/K^,aG=7be1CBEFWA)7Z_gM&)VBURCUP1)=NDL,f_)#
1>UeGEX6eOBI@4BLc.YOd#H8TCL2[D#c5F,K;(7/_O@Gf6N5g3R+BDA)MVUVRULK
R>LUUcAeB:ODe&X=USX_@UH:X9LWHHaa&8DYc.#NNH#YB>SbQf&MX58GdQC?WJLf
0L:#;7\R/L(+HH>VE5<_=Y\8E\D?[Q?9X3F(&c5)c=G32P_A::U)]1@Q6@FKY\GB
cY6S5?VW&cAH[N+9^C7JL,WW6RfOVJU4HdV=/#,/XDLgCg7).]37-GEMH3ZX-5e[
a&GK+ZOYb0464\e<IJTb4K,90b/UMOe7&4LH8@@+f8D0EQ=N:OQRI=e=B>BS93a0
6J;Y#RTRT9:S\X(Lc_\&,FFXab6.[Ig6O,?g_G.ZDATJ5+.6.62(11,#70F9:_0U
&W4NQB_J95>c(Tb^e)L7a5#;MaH\\=)LcZ_TIFS)>P,6Q+UT+gFMaT^HIFD4]=I2
@-=/3.gXOHH58IK5KA-\?_]93bdLOb<T93/b2=7?LW^5c^[dBF,R/L),>]&Z/;KN
C&b#6\ML#.=R@T2Y/Z92Ke:=C2#eM(;F4V&]]&#<GF9:MP=():5>a=a55\I?Z@HH
M7f9HXeNKJD4C(2gTF>Ra<&99Q_Kgc./;A-PYf?=DO\6dH+B@Dc,AHa&a&[g_)2)
C)FSd(]QLQIaB-D7[d(HJQIQY#0BTVJ^C?C[DD\HL<\cS-_[b@FE8ge]P(3bIRJd
V(egRH&eX-I?]/7O<F:E:6=cD1Kg^P9YaPG7&RMDPfb.KGeA<&]XS)4g4#H3Yb4=
FXTV;#67]:;WZ&3_M?42+C12Q4RV#Z@Hb[:gWbTUID8UbA7dLW<1eN+8B^9V,:J9
VOYF3cH0H33SK@740HMg4P-34X@#ZZ:Y8\aVOM:O6,,+\.A/,;)B\Xc)A(85_]?K
PFDC).X-ALP=@&HE/1W3JOcIPKgb(YUf73/G&,3;^O;J:GS3R^T.W7P?KTIROK:0
.C^\YFPbI[H):18TI_Qc=TX0EV#YWNUME8(dCI\+-)AM/DO9aKP7+MIF(LP^/GUX
=EHI<#RbY9M=7-W/?4./OJL3=98;U)LP/XT/N@9bD::/\YEC&YAZ7.5g/->bDCfW
X7;:66)+B0PQ/<CIU-P.TNVK]G)JIg-FbWZF3,>#Bd];1NK::HY25L?H3d93b8aL
\Z+T?)ITVd(ONMH>cKgYQ@](@LfJW..8A/+:Zc9cE_g<O#fe:GP62Tb,-&@8f-#&
U(/DXCAJQ@0B[Z0Cg.,O528=EUg4QH(Q[7YZTNf5CZI;&W;ENaH+&McKV@<<0d2d
#.C7L@Y>-RP\I8,H^Xbg>?<J\:;GS?4K-]S#B()+Nb;Y\:T_>JCXO^^(Hb\MFd.c
Q3\M_4PYIFc[cR#V&Ed(1)UCg_,9C;;ZOG5QI-[>aWF^V(bH3L#W:5CYM=4)fGUC
KQ>+b07]^ZF20E#5[L)9AT5,Pb+@<V<C5HLWQ=18]KSAT5\477TGgVOI7-_8g8YY
D(Na=b>3d(3>G6.D8590OWc9N;9B060)/^)>]614\WDGK\C,aJ[@5E4dBW3dL-dJ
gfACg-5+/GRMeG9IZ?KM\7OW?W^TX10SL/LX1d]V4G#D<&;&ZVeR@?_fS<Pb0/0c
>Z8G2@;/eJ#8/V\XM_D=_g]2TJ+-C+b##=^Y-G(/#Pc2f)2CDUgF9<J:?LUWeGEa
_T2+=TN;X^=Q#5B[OSTA<)e#NO05>XVN7Y6@HMCER^IIVLKQAW42>?>B(M=<H52T
8IAKW6VJZI5+O(L[c)W,_+[HaI,[TBN\@E1HHCHX[RQ<9T9)5C8cCIYHEd.ed?gO
/::d@#GQ=BK;1b<[2R)KQV_Q;g2X):-WECDNc7B+^R:9/44a3e8:\M7Ng0&<Q:A=
3AH_;Te3f7eb,)4\R(EY\8(/(0+g[bKT9c6A,Cg^V.[9A909-QCdGC-bB_1\(QVN
-QV(J]IdM&bTWLAdQ#gE1)N::W9XA1U3-b=U-Q,^PD-F3H;72_LL;c,5\JF&aYTD
Rg&G=1-L5ESB@5dBdX;UK5R@[1B6G7CRBWZ;?Q?2-We[YY>NR-(_N>430/B+HKd@
Oc3=1XD\I&_C(/cAe=]N^EbWe\FI=Kd7ZSTI5Gg76eaS+PdZMOd)Z@Cag;-W5A::
AUHW?)27?QH\^Y)\K0D4;..C.M-bCGHNER=J,^Od2dUN&4e1MSG_Y=&7VgO0@H/U
/Cf+L@54cQNX?0-HgdG/D6F?RGPf@4AGHaLdE\A6]@Ng,+LA[&IS@9DO.Q,Qa&A.
C)K7\e;J9L0G?;;,BGYS184OU;GA@ba0.#bK(4AM9,;K(FA#8DX<\G,A.4BbC>cZ
(^IcJS(bLVUfK.9G2e]I#2A+PX84XST4AJWbPdRBHg=c0,9gbg86SgDB=c<dZ4aH
9SJ78]4eYB/[WL.Y8A^dD)(^XO0K.^&R1F]DR4d&X@5Df^Df6\9/_Z^O4g)J-R:H
b14=@eE[N<Z3g@X2-1RQ/,cAH9<KI2gaXP,MWNS:9@;,VCT,aLK++fbY6KV)ECCT
BKS71Ba:\897?+CC_(2_M7GHRcdXQ2cWC[c.:#J+I<>\;c_85U]BD2=M)UQ(P14P
<:)G&Y^EX][RX]K:6.SGgUaLX<J-O7g&MG(Bae4V:e#Z9IHK_I0H5b>FFUE]9HVc
\0/A@N>..PdXPB0U9(I:-;dG5Y4;HL/eQ1QCCC\4&S,XHQ1BAK/L>6;0eZf_D-_T
8LE,\EJ#AK+7fbaU=CX,43U\+R.f)f4+(740+_DFUDL)efNW6()&>bT.SU,804X,
_6-:J]ZNX0-e]=V2O1:_(_7)<PU_N<Jgb#^6dB0I(W(^MVT5.[SK5.>cb>=.\./&
2d0J[+A&=;RKe/XO;N<D>OQffV\[:C9U)LgGWC+@/[T&=O):4>6BCU4LN&UQ:-bT
G+e3+NI,&WC4,QVcaT]+a+AcA^fEcgA_5e:V,GQ_TfPVBKHY6^UfUfSZd[SU^DaC
1UZ\^TWW+2_gK@NTN48DT/:deB+;1A:1>XGfM_U=DfDQJY.&eXYBeg90H:EGHNJF
B@W\F1GB0cKc2GK:1gGfCdYMFG5,&3dOc\.5U0,Z]7J<Z#1Ef#a:UCL.N^YNOD+&
70?8:M5R_O=0[:];D==PaB]AQJYO3J[08BN?K=T6A(49b[7EE#68G/aLWR4J?;?8
<8SGX+2G@V6]f<YSa@Pb<I>C=1Z^d>Ga0d^U?d:QTO/KM,9X[N-1,)Q:U.Q0)\\Q
\,T);]Qf?JL9D,7TRCTQ.Tg4[)VgSUXXV3V[ee1ae]c>GIb5gd^.OR;aI(NJK/@6
#=8;HU)=J\Y,fcGbX,12F3=DQG?aaS]KER7@OT&?cAbG/OWfVgN?+,C+b1U(5c0d
PS+FdVQ/\7R1ISR@HRASN)#^\NP-959fG>#V_P>[F=<TbfJ\b59JdL.GZX6R&DMR
&Y9]Q:O4WNHg24\_T(MWU2Z]K=eWU-66XPF#10E6Y3PQHIef>U,FTHee\Ia@d+37
#1HW9+OY(HZ-c#BUWAG-4O49PgKKfS.T8SDJZ.-7bJ.DO25a+TV_-gKTHTgE=XXd
8T@)6A,4,)e_E6e,9Q3NUT.FZd+5WDHR,;E1]<<DgOW(4>+G1QTJ>TG9.@M6<]<_
<TOe,LD53OJSJ,38^#DJPc#(c.GfY4?[)B<[Rg#C>_+X&1G4aA,&g=,M^2UE=<>9
(/Gg6J=V5IY++WbOJe\b#IL.1?)S5@?aeNXV6[5@S(9R^P=[>Z6MQ7KQAg(1L:#^
(KNS,,C@X;#=2bS0N(@EQ&PR&@E&SP1S76=AeR^WH2gP1f;QIAg_9L_ON)GY?>@;
7bLaHf?SgB7-AYaF&6^LYDUDGZ]g8:gN0[ee^H<N(6T>(Z_DT-)GWaU@XS[S]g5Z
\SV&bLIP1CAMRV^&DO1?)\]A67eB[KH)[+^Be9\)W5Z;:-<X&5]XTIF3AS\)a)g)
KF?.E9.a8H#+:Q=X>;X4XC+CH7]Y/<7a?JMDWdC>4I.KYc;OWGN5/),eV.]E85?c
;>Y2Hcb2VW@1&\d74Zd7DPcO^7P?2),;Xd>DHDCA)UF:M:-8bTbffC[&O/Vad-(5
LVUaX<c)&YK>2+PI[64RNgFP.XUQFS&:T3.URg10dYM@B[3e,396?(f9/\Z\,T^]
:1WGaN]9#WFA^WcW-K]ID6RL0ee-&C,2R9FYY;,d>_3/VJX)A^H&EMR&;0Q_ZFY)
RZQP9F(O4WXD]3>=\<?YI:F8NM093._I0ad@c?X7T]ZDUU^4SVJ?O]27eK)4)d?/
QOA]Y6ASEOAS0U8J_+N2ba;#YIL\YEG;ITLE4VFg&#Ucf+Z]]_8)-RHUVA-P5-ec
?e)#-+(5=A?[,P.)HZ;Z;#87QXV4&D-bMVB.V0OD?=CH9P3O<?V?dTb3Y3TIefb5
De;;HYg:5#J_2HZ3Y/]V;P,gN#Tc[3ae1_S:C-D7]GZ+NYI.I7eRG[GU[Y(^:46H
;(\M.3S)_\b7&DCQ).Z0OJ[N;VT_g0:_V@(\?P5G+2#H(&4RZ[NddL&2-V:7I=&I
PB6C?T\,J-VCQRJ:4<aL1LQ9MQ]T@O1=L;c]TZA4NXe5ZWHdZcC_QSI?6/J5dE[9
@.6FEUO-e]f)#OK0P(TX[VN3=ZHRLUD,Zg30L[bB=Rc31)Y-c;G(.e]09&VUBF7#
5F/:>>\F^UY;D=OGZ0,\55@dWab4OLefCGSd_]J8]MZMCXb=5[3;58:/WggHI6S5
\f0fdO09I\DAUY=Ug7BSJ6eGX==K83PC9EE6NFVAgd8G,;Lf,9^7=;BL:aAdY^?>
TCWDT9KSO)Be530)2Z;S(>1G)._f-#?=G:6-)ba7:.0WO;OMN[bA\4?>)DG+9NES
35HY9Rdaad6S:&YZPa??fZ+E4b_)ca>B8W)=U1.QSW(B+OC=DN<N<5JB9NfWR>4T
\]PeW2CfN<eS,-1>c9;\=C.U=:.C<RPY7c.NS@PaF\2B)a\#F#&GGd)+R+5>a=KH
,&9f5@.Cd,(/E59S68^4W[JM_S.16A+L,2+G8/O,+4SY@OZaVTN=ad@]Z4d>5.8b
W&48)YZc?#e/HfdbPDK=,L(PQSYU^[BE-K&?^+YEQJ/5Bc<=TdJ\_U]):Z4K\9_]
aCbPLY([F_XB?5R;8X?Q[IC<6KGd<)RZg?@TX1B8,7;?=1.\GeSC)4fDN-gHc)5G
?&5)>2?X5=f6Nfg;ET:0e7#GLE2M[YH>95V2PL8J>Q5^]AT]b@\e;+3E_7Z[BV?a
69?,X96=8B(b(SI6<c2^,]Tf6D3T,BSPEW\JVK,>4=O1+:WNIe,>dBEY\)F0W,?e
PVRbgf[7bL_0g[aK;9[-DPDZ1#L9bZ<:G#@1KX[+Gf/S(c(I/aQX0Ff]FQCUL9T)
A;QDWRJ.XVDWbB5FFIOR=;FAa?I=CR[,0;P+::9J6:FY?+gD#K36H<eF^+HQ;;UH
>UIWGWE.c<OZ_P[(42-1#L]029A(M.BJ@?67-E-GT#KN2Wd1c<776?G2S?:NNL=5
@Z>EM#cV6eDQ,5BC^)a33<?<7/H70CgU)F_ST&<>Cd+5+#P;9.DXO0N?L^_[X=cU
+JK0@+G.Je4+^(^cS1BQRYb]YXASDP=b5d3DPA)+YD]Y.ICIf5cb3N@)RF=06=P,
MZ@;[;bT8C&f/Y_gEgV&98+3DZW5F\a>0fgLgZJG8I.:D+_FfBLg90.=CZM,7YJ-
WV1)#WOES<D6g=<PMM4bW]F2(_Ig)/BIK-^JF:gd#;C;XA9:V(B/3FGf@fd0E0g)
\\Z.C8Ta)^8[cf@4:Z9FI-Ze,[<YgWYJ97K\//e^^c:Q\\M(>A8:3.&>C&BPdK9D
[K1Y8SOE2V2V)>@KTSW>G_)-CJ8aabV6)bLN,]O:R+,PaR1R4>^HB5.a;/U3Bbd5
O;V:FA4WAE&6OdM1<d0.CQXIJ&V\1MCd=K8DC=\d3A-]4XYOZAI?^^5bZ__C7>GF
f4M.YaOfU_Z>fG\TMZ8TTGCNC0/D,[7:-HH9XgNS#+LM0YICg[V,7V+eKD<2&_4(
Y<bbUY\QE;f3O[H1+<@aON.59ZdT1eQ:_<C[5&OUf[+=T^YA283B6(=\RLAC2P\/
5C_0GcY>^NGU^OD+g&(:_T+KN.BY>[,B]@0UPE]Yf_L63W-V@g>DgcGf[;1_HP&P
MG&1I[)>UMMgM7LS>1:;EDAA6SHgRCHYfJ;=R)^_[.(J1>J8((CTX=/R.52G@ccC
/A?>gTRHcFF[-39QX=;[F^Y4b0J9OPZE/AAT-dNI,Q^1TF)<VF62)gB<<E0H#Rg\
V\Q</&)gE:dT0+caB]c];9.+B52_]54TbR<0,+d26Ta.&.Y:L3O]bf>_&]EJc8Z/
VEZYQ#&?bM8TQ4X>;4\,fKf#@][F3-d-;=LQQ\e]ZZ)<-)^#ZaL#Q1>1PLHV0&QG
geY[Z1AJ_9--?S\419@H_._P4-3/bHSO(_7SMRP_^E2#3egKW-=4ZAa(b^-:<3WJ
&CO[<[#S>@+72Vd>I0VW977[9HCX-cWbV,BE,DaI1V>>_61>FM.74D,5c/YQ34\4
(V0P.g(:H>c(8>^.3HYRWEG[P8-CI=TYCe]LI<PAY<dX\RE<?^EZX;W3&4<RNLSV
HTE@g>N+1#U+e2cP)]&dOAU[#N-KGRc=TA0SL1;T@bPD^LZ<WS[,9KM9-=IP,2fY
c-K42_?@(:]Z;a2H.+[\N1_1.fQ6+FR;=AJJ3A1#S(_\_5X#S@#0==V0:<0cW=e&
3DS:].c5)9g]4PeecO0-geU9_A<KHaGR3J_+I67WF\IH_M>d/AO3X2V@U2&G&7+W
AQ+JYC1PS]Uf[@;R.ZIGX\c9b2Y2eK9+ON2KX=&@][9L[(SUQMS-(KJ-=<#YJBdB
\8Y#>RbHEQFFNJ7V#ZLc\+aB0aZM[SE_-<bMFNC]]C#G<[&QZ5?@79&cPe530:La
6bV\Gg&#JE)=6]PG_/WL5\d?Kf[;>6gcT5+\>NdET\@SO44?<>79ddaIdVT[L,9D
,c&gA2>[UGC/X[HR\Z\)>O-Of5Z-&N>^\I=^f3G^g3a2T_(&B#:VF.\#VKE:0I0P
7F(S35\E-ZIM7@PL>7HeXJ=4N[&c.@fC<ITXWP;N-^6MQg[gG<SJM<@,K9=3MA?Z
WKXXS:aOO-<X5T7@]2^B#OH)DL&A>Z^3MG-J6fP98S?DVf1I,c^77D8F/XgGUENP
9(?LNRNRMf,?fdd3>3Y)M4.Q,4F^bU2U^MYWO/ME^HQ),H-5aCCbVBYH?e[A0K1H
G^+Cf<XQ;Z[^JXI[,:[RZWQQC:XWD69=/FdcR6AWeQB^ZMU4e7)CUQ-#;d@G>>S]
[#5/;T7Y+dD7_WQDVH4]&PY^3f@Pc5dE?,.2QE)?AdedPPFNe[P-.fW9Q[452aK/
EaO+U)Y\>g2;23dfCdX6,<^=c;)98<-G-d#HD_);=U&Y8>a8>.ScY,NM>>RF:-c/
Q\;6\C7,HE1>0V_,6JSA@OIJ83a&gG>0^.[9,SAG7a/c=CdgB)I29\?5J^#_X=d\
(6O]<5N\2L@27DND@^?PK0ScYg;E+cX3[ZJ,,ARQdAWMgL[6&:N_Lb6AL3?Y5^=B
5;V:QEc),Og\&2BIB7-I_BAFe>]P(TBF3A3@[2e9\)XMBZ2;1ULg-W1bBA/1WMVQ
ZU13WIYD<8,MOB@)5\0d@[VT#[9#2Q?;BVE?,QAK0LC-W^XEYB5A)[0UO_aB7D)-
b<GU-J+#18G9eQ.:^8RN6aJJF?(L_=b98>LQYDSLLCK.4_+Z#T1cI3AZG2GBXB[5
<]#>[(Oa;W<Q/]1NJD=IP-][Y)5>@@[9@I4Z@U]gVDLN&QZNN+gI<GN<)e4L+B+L
gOEfXOc\RS?e[N:gC8g]D0F^)MRg/=H=FZ]&[JR,e5(A8#)cfdX(-Sg?]GKJgW\P
4Z0Q_1G]3-G^0U\_RaaOPME8]<AQ\&4/@3P-;7+WT[Ld#Q9I1dY84G[)R[cEA-P-
3I_d=SQKGZR)8cTFd-dc=af02\bO.^)O.T?Z#:)BN(C1=IRGcV2PDXF=^+[5b&.8
d/@A?M6FU4:c48=ZF6.,PG_U8_=&a@?,cUL198-9:3cD4WSHYN[-_P&[B463fQ0[
V/3Q&/a3]=AS]M@eI4_[9&D4:-JHXVP:RK/<&(2KD3)YEaD5@4PE@IFF)II+5.@g
DbDc8@;dR;ZP)6/TISBYBT09/-E;S)4CYeaBT(fJNVb@PF7H/V//1#B1ZBOfM-BI
I(;c#8?6]8PdF8ZcQY;S<F-P-<00.G&F4>ZbNP\XC.IdONE3@9?YKMT7BafY_gU-
ZKFc29PVe/+LPfE/8VgWIG/SBQ6@50=JEIe)R>^70Ia&CX8d6M&[/VAO;CR.MT<1
==)a6YI_LXZb,?dA/I-,F]OC0;YHZ@P7-E/E.033+)2@OWAFY8WIBIc=&N6A3.L+
060MFAUI^3:[Ud2Y\cW1XCBJ+0G^G=.Q7G<8.?CdP1H6-ZYC+]=\A8MWO:9(Ig:[
+f060,?)#)b>@ZgQB#cY1M2FB4,IO#@8.BY110_JR\146IJC^f2OBRI><5>(AFZ=
@@X>OJ6NV\#=8WE\gIDR&0(&3_TXVMYC7FOYNM@_L+7gfI^b>MUZ9.e<ZB/H,SC)
O\,;3MXJBcfS#H?RDBgEJb3+3^?(KS?FB#CJO3GTEPGa_bK-@0NOaa70QZ-2:^(_
H^TgGZB2VL+=Y(If++\=Y?2-QLO_a636Y90_.[0)61?ZBZ40]cd^1c=4RPK==(17
Re1eVd<+K7fWP[<;,;bZ,YK=10GMd9+08Q8)+DR]81>=FXKUEHe30WgcYPOVV&5@
4^Z70e9Kf8RB+#Y;]&31?3T2fM:PZRcO@(:&M3FF4,VC@dXU)XKM4B0P9GM#K&b=
-7=@QZ-N1]LPY@3X26TS]fNY#aZaAQ^(N9W8<B7O?..^9/@#g9:NEUH7S31N:N-0
9J\Y<MAL?(VVfF^gX8O>:S3DSS-,,aa4AW,OE)VbF;N+7UTTF6\a8S-e(;ZQ/6.,
=1Z]-B-<f+V/9A&QUF=YDRQ8JXJfD.eL<dV0VGS^>RJ;@LEcG=61+a0:g:+1P7@M
dN6=)N.fd>ED\<IgD&.JLgeF<_F4BR8@KL0X5FV>I10_-+RAECJPYQV#+E\UAe#^
bIR07Z_14(E>6PLE#f:Y.^b.LB?Rc\Q/2-VG8.Q@KB=A.>SIcH8eTSWA;YYBZ7/B
TT>\d7K2GZ8N_I=<S=+LLCSfEdLAVfTR0^LG^BUS4D>J./JSFH&c5X4=?Y[BCBVd
bZ,RW/K\=3D]a]CRfLdUEYOU\X#L>VN\Z8I8gf[[CRgPV<0<^<c7;7@1&D3>5:_D
]6?@O5>)g\Fd6GTdE9[?C99eH#C5#NCEdGYQeYLG6IE_Z8CYKA0c:.g0=DY)?GEd
UI_T70&7g=UHN;G/#_U@49(bDY^IFH,cH4?.1N_5P7V,L]dEHaDA6^P[@]RVa)6C
);X6R9G)&cRAeL&5-f00Fb?;DFAF@8-DJ+5^-C&Q3#[+H]MZ@+-)@b[0LPO6M4d\
[(3Z<BVT-\&@D@IW6@fg8\Y5]-/:X[Q&#CTEN)cXFWY+WRUHb>.S8]3?.#G\E5SJ
a_QOfC^)VO6Y?4;&dA@N[G7X5L4F;L.6JfYRMc/e,G^TP/9Tg9_44-_L[Td64)\<
N1&fTL57[d@-;AN7I1+XTU6H)4ETTd+[O>AOR^3T+JS:+6C^UVX+VZ,N76G9b^JH
X9:BA]HV_0gHXJ;WCXLAS_,MK/6NAI(ORfA)J^5:f&]b79e9F3gDbBB@-\+Xf/NO
TWHZ-J2J#8MG4b==ESKF1MLf1IT\19[Id:Ca^XHY:&RY>U]Ka#K(OU(=1aLEH0O+
eXAPfDf(cOE\1M[JdX,Ff)ZL=SZF#7GY@(Cb:3b\>ZEfNQ/eG:N@3JWP3+g1]563
60+X58Ff5M-5a@M#e-2C#A5RbL47HVaR??V.QCGfMC/D=;IW.J82\C>X)[8P.,7^
2f7:+.XABcF-CBT,IVJ^f[K7>aBOaVEVFd&Vg1UB&1Xf5Jb^9_X-B5SYESXN@/5c
.XM:[0YMQS:dI#(6O9GZBA,TXASKI<Gga,)@@B^3E5LWcK5aN_4D[J<LUVEQ,3df
fJY1<I\+\X6VTd001ZV2KM]^cU1=TObN.Z:92d9N8;.gX4Q.(Ad/3K7,SbdQf[,]
1=JCG-1WXbV[cICVHLV<c\N_K^-+RWT?MYBN.N./4#4PAQ<5XA3;9,R46Za[.K_+
fL(KH0--LNUd/.>)Q_.ACSLA-b(KHN(c+J/8a7-L12+:?^UB]J@9H&=gY;c:P[\Z
LKM,BAfJ4+0/>Z(HW94GQEVDC]Z<_a<10H:>?59U-PWBL9.T2NgB[Q2)#5A-3B\c
)O9FHXB6EbXQ#@]&K&=/TYa7)0</aG9H53VO7F@cBE,/Of^DTd2=:9O4CdB<F\5E
P?(>TK<cg9bJK_J0E4a5#ZR&V@/IP1UU3GLKFBGNfdY,9AZ5RCPZX;H?O@/54,#A
c#;R:[>gSSILP@2f)AKL1W\ES(2.R]#Hc<=4=eH7LfVM5M,M_-TYO[K;A(Cd7&81
TZ?C/:;_FN3L=&KTF\O6JC6Qg.BeH:CYU;Fd3_UK&9Wbb&.S\KH,0&&;S/LTd0=f
/0?VF90>0:[P<BF>(GU3gCZGLZQZXMYW(2J2d;[3AA&ed/DaUd,R<#IMXF1f<eSZ
@=ARI1T\T.>@&bEF67bAI?fBSJ0Z+5e#T3b/DJ(UX>I>DNdNYXO0RUQ#6@BLK>fF
PX_BWIf9L#/JcIfF:Ga,gD4Jc35D?Wa3WgW83W+DMdf&6RZd]Q_S>F_S\5S&Y6-)
ee,J@7<]Qg,\L1WZf&:W\eQ7XOLAeZTf-@SeVH4_J[3]e]6@LICM[4c2:e&;0e?V
FA0:BP:^Z@5SCa]4NFOI7)J#fR,b8YHK8FGWf);A@?G(Xb7L(O2BAg^U5M3NgBQ2
G,[:-ff)[aZ[[g\U@F9JYc/]K2?[HXDU=KbWYCb2S7ZWXgVdbcV,[a530#AdHAJC
2D3Y,9>1:#B=5V><9@-&gJF>4P;5RA4((V>>XX-XZZ^QgA7I,=(HUM^4B>;-:&(T
8Z5Q(W_1SV1Z;Q^?A&;5EFE=IAU;.b3-OOIVPgSUa;]D,5L,+@&6L&5:?X9A1JAX
Kf/I3T8J4C&D>\ETH:A6[]-:C&RM66.(M7V;b_M2OF+I<+UXVC>gTT#G/SNMS<g8
Wg4S+EF(YRAVcX]59EGPK0C3S,@-<+/Z6/b0DM^IbG6:/B^SaF[UOeUZE2Z]RDCb
J:eV>,d8=#6AJ5.RP(D,G9V&BQ,/fITAY6VE0eP:+HQ;NU3A8DVdFcJ;Y1V)^_U4
(c-SW^Y+H>,N^9ZA(TQT7-TYRC+<U@E9K].[Z84#JeAUESH+C,7LZe)\>0IPDb1:
^1OXFgX,JfI\M_2/IW81?B(VQ&-?GG3LK&TeLMe59Q<VIQ&-Pa;E).?#/?(7AWHV
J1a>ag?.WbE;fV<=aI6G7CA(@]\ecY?KVNT11C<<-W0ACMfPERe\LAScXMKbW:7K
01YdN>1O4\:fT.5T-Ke\XM#E]1Y6#W>,,-5B2_W7C?QB0gPf@0Q4P5c>JSP\JgcG
TJbR[1;A>EF,2L93NJ=UdM>F+,>FPe\eEPTbZ>+VcDX-[9X]0BCU=;]X\XK3?a>L
=2-V19CdMS+La6g(O^\Mg((YU>#IYKe5Gg?V]a&>5326aJaA7-/R>?,6:H4\2XSZ
aSb#PZMcUe3[>gH+A\-^BUU=XSJB&54Y1<_Z8?UWe+Jd_fEN+HN]g&9VI/G]O9GA
;>S>@_GZIe>OYbJFCQH7R/)F4Yg&LQ;.;6@OX@/#&:)6VS//>5-N=6QZMS<0HHc]
d-AFVcNa[]O38G6Z_e7(N]S>cOWJgIOHd?/R]U1[Z(=;eY]5ZF]:1:L5MA]TbP;J
(3V^<P,B]9a1-7)b7FEXeVaDT,Q4c1>L;\Fd7BN4W.S5)cUDE#O(>PH5_:\O?If=
=TMd)CCdC]85UAAFIV=^B]?(UKb7_BXL<X8\2JY=^E7N/^@T3^KA1,[&/<]=O6b=
a?(AYO6a91XY=7/W);)U\W6@C^TD[6=(?3BU0.>aWgT#XUcHa+L^9+EOBMT59f[/
4/b163=I;5HMEc#Q548bUXIe8D@ZMf4Y_?H>ca<Qd1[Q^AUTQ\bU(\9(ZS2g#R/X
&:?EecLdTbXY\FNG&8T>\YdL&QERPA:<?FgI)W(cUTIXE6&6\0D&T5[d.4YO7>A)
#C]b@MS&K+TXD4efDYD[C&KJDUV?[c(1SdJB<M;9f;<6fH2JW-[2HB>A\0M9Z>(Q
IE]:b,9O?D&,.JRFQP[TI:e\AW]gdH\@4N:g@;HF4g(0(\17J\?GG2C,eaHHP9)>
&_V^5W8+@LgbA4BdIBSD.WU3_HBG&SaA5?3</PWb7bG/TeA?@WS,YJYg:E75a/.G
?X@X]7E>WZ^ZANb;9O0PL3baa62/Z#3)g@S[[LM:_Y<MS/5;?_:P;EZQ]&DY[J6T
T1O,0eU<[<CKaYUKM1C199GA,94-)[]=ECY[;8_#-4MUKD7;U:;D1F4,fHB)9RK(
Z8XdbcVQUQ1@beCRdVGWT;a28W9S1C-V<I<B&CfIBRa3]7<B0(WOD@W?<@g_>2-+
+De>Pb:b>ZKWLcQ?<>]H5&+[#gY1bgNS/Nb2DV:b9IPZgIB-LIBC7f:445&ZNFV0
G>1/\cW5G=ZSdF?-=D,D\=3Rd/a-H_=16P9_XgNEb1CR&2P[bXBaYF37A4059C:B
4>G<aHKO)g//\R4aJFFB_G:f;5]IT?SHPgX.9e<DEg(G>)WNST_BY\5KPJH\>LKb
CXIZF)&+;g?3+YB?V7ZVI=TEX(1;?CBFAT.KD5TI;Y<\]V:;LCXK5^c+1IVa<e\;
RGJM6JT05e,^^V\9>OgT?BW-@E>Z1#](IFGCDdG&<P7O2N)PQ/^QG0fPE^b\_J[J
,0DCT#3.cb1bAbE1bE#S+:@[TeN\\4O_=d_cM?IEJ3P7dAM1XH;>g)H\c3Y0-\00
B(Ug_VdD;.Dd;45Z)8Y(/IWQYB9U13abPSTMG@\ffc0[[_g23Z86EQ,.Ta<ZC;e5
47>bc\PYXYe5K@E)NXQA[PN/2[>\3J34bEY/Lc6E;).=A\SZ&e)K@Fa<]IZJ>)-.
QU\f5.D^>,bdE?I/Q;+Q8P,D^NV.YQQGM6(9Y:[J(b9Q5+<b4.U,?27\#7->5:e0
60FPV9XZ28(&B,8NR(+0&V-Pa^E6I5g0X<@VWReNTW?;_A;C^XMbD>>C691-0^Df
]G;V6Q\)N+1D._&NeJFMXW6ZQV(AVGNMTIE4JRY:1EE-3M^#NSNDYAU<&59@T3(6
.WL(C36a.e_9C?C2Q2UTCQ-#-71Uc5041\N.L9W5PY==U3IT0W)f5J9XH@=B87.P
>]ZVL4GV7UYUBMK\A&<4[DUS4K?0-#WaB9d25cT/8,BY70@Fdd/Y>1#274e0>WNA
B?:O[3D4S0FAd.T;>5V=ZdIX9fc?T^;3L@7A?7<TCH1b)C#:7@\LIU1d5?>A#8?V
J5\&8OWQ4R@Lf=1E;H7>^c6bWaR)U52f:_=3ADg<9ac]M;,:@:4SVBPdDP5N8X@=
^M:Ad8]R1()926?@B-#S/=\X2FTg-G)<5/VT25N(CQ81TX3Zc(8--&\b1U.@]d.2
c1>W2JP=N7GbVOW+5,?(-4?+[ZUGd3AG4cK>\>_GdI8a/T=?^;MEFEg)(5IZWCXN
0-N9_<Y@I]+2R+ffed]W?/+Qg+95e^&ZO)[T7=+T@YW/22cD5H:@gYV^KB-]X&[#
(3WbdL,Aa&-0V4bSWWV6aFDS3_b]R44DT2U@EcNQWW39M63dM)HOJ46[56W6&;bM
&IdNP-DA;,fYGbM&_M-,\X7T[HT>_7M8bfc#SR_cXT)3I(/#P[+]MM6RE1D5SABN
VPH3G>]EM0Z.D<fe>d/J@NA_45c8MMM0g2U;RR4<7XFJI5]C??2+MPP8ef&ScVJ(
_XPE,Q(0WP:3f9-H5YaLcTfdDMaSS[A:8@eFZ0b8/UgdObc+Z4R^5/eMbCa^NfPN
(EZP4SJ@aR0<&7Uc.S&/^@4^[HA@dd@,?A/fB42#HVbOcJ4AI1>Xc6FTG^/F392?
BgPgf0[T[?EC.a.STCfgTY^&@)2V8)MI,;,?GCXYL].<DW\#RKVG1=X&#:@]]e;J
Kb@dePOgb27(WS<1,MDK[&9NX4AC]O(2Jg@\GcAf-1(:SMXIO=+fN([F(;eX._73
N0d(#2L=P6;b_bFLc<X_H_K3B]/@Y36--=>XMfMG/,C#bF;3)[><(B&X+H,,=4gW
1E]+eWIgDaT+FdBcgE1MMY<#\SLZ9:+>8_GC@6;&S3,bU(B1,7dCc,U8871><#3I
_B4F,dVgDYd<[,:B^,#1W3K;K]54/_WBYa?BO/Y?:\T5R3E<KP=P/#]UO2b@+_T_
F5IJ,]FXOX05_WM88P:f<+Kc;g-0?9XR:M=QJJNaI6T_9.6;:UF1e>X<DQHU^JOR
WFePS8B(c8=]WS/eg];cb<Ba>)HP-d_S1QFS@CWRMZN#3:Ed[#48LUgJH>(O1OMg
@8>HYH;N?3,_WfI:2]6+P)f&gP^AQ>+.44FETBZAd(W2_K+g\SfZT#ZQa<@^F.3e
(SUZe^YJ0/6K[bJ4],]c[;M^?5VJU,I&bb6FV(4C588OYcH/F4(LCSL#J:HVSF9K
72,e,@D(g)E-S2^FVFb?0ceMVDSQ&(NT1\DJ+a[7O9^eR&?4b-;,Z:IRCR1>-V)M
@TMEMB?_N&C0Y&Y(dCZAZ3<NT#I]0;bD/.8gG#N@g+0P87:d:6X@3.M4FINZ)X[>
IgIaH[@B[Hg)Q]BB1K^CBF=(H5a(23L06Za->&61T)G<0MKEX_M=<(.McF5\ZAT&
/\Z^S/K6T2d7[]6@4ba,eUWWH#XOHOY<e>,e\dZ_>HJ=X]IB67NEf61=6V388(Lc
Ud5U)/Y)YE^_CJ,DbaKR53J(;-&7cMV7L6U_G,3?4<3M9\<_EPd48@T5Fb<(F=ZT
097QK#(fGS<Q;ZEdX;\C^N90-?I1PC[AO&FRVWfD7R7DMI+IY:R.W9M#/_.@1/,,
WS+]Z45>YEX<?[)IH=8_Ca[I3fH^e_-D)^HUZ8+:3[Ge(9gR[dRcWCG]]@V:^<@>
FDcJ5Wag--;XAaD>HV]cOT,;F]dDNgeFL07.@3QP=.g,=7a@C,Z=;aP1&\TPFU4L
=H1]L=]B)a^@EAOW+_5C6-ENG7&Je0EL:)S@)?:J-EV):1MJ]aH/+(6[4e&<<O(&
J20.d0W:H=YFDWM;K_LXPQdJZB=\YJ0-X?O1[3^W-EaF0^V;,&dIJAWJf#g@F9,=
c<?YId(1bBOQ=NDA6LS=S=]a1<>1.9\AIc0<gD?-,FOF3Mf:dBTCN&6RHONJ(VJ^
Y@T^D+D<7QW9<CT]4,&2U27DZ^DSN-PHE,IEd]=YLf6P;1-N4:D\WG>MF+S>^>BA
_.82Y7,6\c(b]@DLDT^LM++7X@HHN32NI4EcD]ML2OcK=B?2:Z_8,fC9c8f(<LM[
B-H]#fPgK-9PU?TC\aXV#>MV7=4Z/4E-/@VeFL[f#JM>,C=E0KdI&3EN(.d#Y5SO
2-+3IbGD:B;L@@@gQ=e=C-V4MGQMQ+2F_3<fUJ#-JB<Y;&XHc.SL,@0[@F;,9g2W
efZUIM92^5M^X>GK.Of6d7^0A@^#WC[a:A_I@.U,7V(2]LG0J7.a^>CBef@3,+5Y
<(53K4WJX4OEC\0YFRHVbGGBBdg4;D;TVdITN02JD:[J.8Y<[XdF4-O?VXU^8-?A
0PF6O4<[3feL_?Od)2-&BdZ5OBP7S9.\0<[a_86V=E.49V#J:=8)N52@9Z/8?FON
&cV_fZf8X1,\?#YQV5NH8a;KGR:>#?-e0;LBFf?f5e[J1Y;QQaR[?1OY+J3N_:>V
U]g7U[<AG[:/c@M8dC(c69L<38T^19b[EC[Y=PdCH+[/BM[/:g?,N1LGA@K96&a@
_2GB1FBZ,Id04T]KVIQ2dg54L-P0J7,PfMV?1EaT-S82N(X)7WL\9[Ve?POa]49P
_]c;D-:F>8@<M\47-H9O]1YP5J]V#[U(\Ff8L2b?BfY=)E^dHS=F>^<U4;g_FH1U
F^G>;Q6\/;C7<-6QLb=X@>K0dRNY,J-aFCPI\JER&U3D-9de8@]#>.IAc61Q\gJT
d6g((0O,Sf2XF0?\GL+N8.E4P@S&/?fW&APA[GWe<_55[]A9SD3fNc7S1[+BY];S
BUK\106=_?bOF#/;E6/?LcTf8+eH\C1X7E7LFD>6(fH3A[Xa#>Q2cJ,@:A6SO;[B
>;Oa+a^fY7EVT=6bHQfJU]aR.>PI/>8C3g3,10XTN]5;O9O.-WZF:7\dP<=:;61f
B6eD3Z^U:5I]g;\-WPK)#Y+KUQa[S:>(B5?71gd?/-0UK0PCXM>ddMGe[;e8-)F0
-C^O-CUFgGGd?B[E^SVVa_PIHM;)/L;@[X,]D/8/[VWN^eA\_;ePD8^;Z9QE/.Sd
@QQE]KMW+?5>HSTS/U/f54DF=\L6QXAa/O0UVAX<6]f^>e349GD/OdEU-IU;4R/?
U8+:D2DJ\7-?+,1/1D)#9O1f[]7J<VHKXD.#5Wa+>F[KHY0UKEb]),Q,RIE\T)SQ
S\]CE@1g^<AVESGG9TeC0:D;[7.U/-FN.Xg/^e2.P(WQU.5XDKQ+1,,]0[EVM@S_
Ae?OXP13<A/EV9>CY+)f:A?;f6]d;_/?3^WX)I3+KNda]8:Ob0883<_JF3JcTHMD
[AV4LT^LYN@5^H5dH=:T?2TZZ@4&)g^5CAM?X;D26e]F#Wf_,AWG(ge=cUW&ZCE?
\dD?bf4Sf8g1,L1&D/6-a=OYBM4[-Ld)TE<WZAg6=COZ@Xg5];P^,e7NI2#ced==
?)0]@3PQJ?0LCFMERASCB.#//BUQVH>P43QYGNG2O,T)#9F2Z5S^;7?2EH.0YLE1
7/f-bS0KO4I&Y3fAV-);\A\\&We2Ef>^Pbe_@KO29V98VGAMTCaU:,&:g6],Xb7:
KM=KLA:[GK+e@];PQZ.AC0Nd/>4gCYb@;:&&M]e\/?[G.#J7U-33-QD_f9+]^->(
dLA_BfCdW>D/T:dYa,EK>fM71^M4KR9-A-C-XEZV8KAee&:\g9a8>(^UR2g89+G#
^5Sb:#1fN)PEDN3K+_aC_[+L3)<MHL:OX7cG/=K?+b.U][AD7]S>LEY@,\@f/1,F
4\=(AaS2QWCSCWW5KKV>?Fb=@?bDH[VKU?LJ)H/K^R:_N8#I29L\S7,UOK/JbW7f
JaUEBCUe:S<f(;M6V7XVK(RHg9G@H^BW^(@Y5?--7fQLfT7cEQEbL)3<=QOe=+;]
,bRCNYAeM-Egb7<UR-/4]H?>3L(K#F<X-F45,&+H]D@>0,.e2:Ab+HWX1.g[,LE&
S?0=^6YU=XOQJ^QJS[J[OZd@J[SWV/BgWP)JSGPc=Z9XV[_cf9T=)@MYI)9,N>+K
Q5ObLfZIV>Db4;Q<>c6G-R9K18[\?0_e8>4,A;gS5PX>LP[)d1&\0-+-6Y8@N>H>
+P;,6fY+?-2X(5SJged,9R\W:Sd(9)V9V2]R9?Vd.,<U6U\Y]Ye>RQ+7EPFMO(&Q
-Ra<&A>0P(<Qf>#LDY2)gFe?]:MBb0MS9;^OX>5#N/^1)A02ADXL0=P6G)@+fg[4
J+cDMLfV3:eCJW>1=Z;S+CGX/)I>&N,BET1NQSRL;(U5+W3EEbBWJ-J=.BZ6W+:_
(4D@=NXTaG@<@UCH2-#f[J5+P&LFU6\Z(I3AYT,ZKVH;<@2f]?U\PX=GX@AO7&G6
E3DU^Ga1;cUTYY8JD\^@VbYAXG#+)BZ-&F,)]M+8>^ARUIN[C.R86A\1O6Y@?[.=
CP7@[=<S,<:(=H2^TI.F#5b&>JP&E=5K=D4IdD>:C]59eNT_#f=N3@fI-^\;3>a&
K0cC42UF3c_B(#)U[YQIDYM4T#:dU\:28S6Z<_:(@WGY0-<.^gbY?8&5Q4.^J2f[
U5]@8CA>T3^4d>@-E[DFQ&>-/7S6MCD1\g?#LaJf:VQMXR)EUQH:a.7g66,a)-O@
?W&3^?YFG,JX<M8-\,RY8\^GHZ:^T2L.>&e@C4fC;CBE8RZ&E.be^L04VgFSeZ:^
#Mg]-181\aRSa>ca,RfaW>8cGcGbS)CZA5PN6&D0eE)-]_W_gVFC7-6[);OM:Q,W
[EJODLDGJI=C/f1M3V?F[IBKF,2O#T<0Y+<b>:7./Tc3V?e.8<f[BcOV_P((2R7Z
DL:F.FI;)&37IZDG.](OV5ZA+SACTW&ccS_aFI?eHIW_81U=cHBQV4U26(D4Wb,A
C_Z8K)5(^KB<PB1KQZ>C)C.5DVP_<9Sg1UB:Uf-770f_f,-NX_A0+=XfOOZY\Z@0
SRVUO-N]bHZV\_daT@I3O<TI5GT&/<J,#NAXL-E3GQR^/]GR#d;;A[25V:/[P3S1
GOZ-F>F[OBeEQ:\Y4^c0,?(4.SF<N2VT1.:gZ3XF)1gNQS5EE(D0M_,=U8^6[?9W
=IFLC:,K\#b<N7Xe9adde\2dFHW=2)]g4LIT[=E<&:D+^_fbH>eAM+#@G50Db[.D
TT/5E5X^QMd;A3(CRHXCc7TO9.FaV:])FF[9fTZ@;YPX>0=Y]AK@cQU:.?R-3ZQ@
Y4;&]IQ,VZ@B7KDC6fE^DcHcL=Q4_\,N>D]6N==e-Kgd@V,,a1]Nf<6/T-0&Qbe>
8_6a1g#(O55,2N]D+I(<KfSaa[AVa5Pb[J2D0<5;T+JC0B_fVB-e#8aM@8TDBVMe
KGHMP:?-/Hc9+L1fN/863faM-ISN,;56@a47G=NPX<>AKKWZa1Q)1++0#YO+gH=J
,.,.#(DEDOF[_COWV]2YNB-=2E\bHFXKTO>+8A5?Fe3Re?AKDNM,Y4\>(ITd4e\-
.bU8GXEX3=-X.D19#UJCX<K_9VTOaRIC)AY&5)^TD#Hb^JTL+Ue/^PC#adQ&Yg8N
7ODa=gd[G;1^0[,6HX-G0g,S5/Ff&bBN30#Y20g3^=I<dB2O)XHLG^DRDd/H_I64
W2\9fL:E;K-(4W;M)Y(AN1a80BZf[Y8C?-<1,<Q0<5W&d<A4-I1@&>O#EFe4=()a
9Ufg8YOMN8^Y1fC(CU)YU+^&?g-fJ/IL_#;3:eZ(aa(e0^OGKfP36X^6eIIC[]J+
MR[9/8Y.WY+VZBQf[I[;_9?a=ZU4L7fe4IA^A[9ee?eV9^+8ZVSR.f7;5SW-?(:g
&NX4<LB-2MUWWfK]9/Bd?.4AY4ZcVR-:,2Q6EgDA>G/@,[+R+3VS0:F(>JYNIgI=
^bV17DVO.R>JGd+YeHD^@;cH-0E;9MH.eY/2ePg:\90I6.-5+Mee4/??D](TQPY[
beK..8W+#Ia&8#(380]L/.Me056OZ6M)Y,<#O>F5LFF8U+_2Q8R0R^FNN94C^4G)
\2.JM7gQb\0M.5,^#d5J?7G6ba<32#H?K2.;1@gP#/fg?9:-13BERHYS+UFHZ#CR
d((fc1_AA@bYE<V9bd[8Q5^)dI9T9W,^dXX1=4aC4Neb,(.a>S<NR/fACc;RVN3c
5?8I@(J4#1FS0Ac8^F\GE7DIO_3N)_IDf;Z/FZc#B6=(UQ]aM3>C1\1+ag#UXC@6
?E)&ES[JIRFg?7X]8<-M>^L^b9dMVU34GG08=O@H<aSD\7TdC1a0-YaZb&6e9KIg
9=0gDe>\YV5V2]M:e/W_DMN9@Uc1Eb-Da093Kb;PXbDMc?J;b=7EDcZ<G&+G:)2-
.J7]JA@I@>e-7KgUYaO2=Q\I[Q)<6NfKLSe7/^)X?I)g9e)-(Af78+[0=^F5bJ58
fKN-X=fMRX4S5dE9K&XeT323KR7_LLG6&g<\V<F=,T\c3_cag:C/5Tf@0aJU^RG#
J#FQ3JU6O?J^=2DU,2LCWF4C2LVd3[O(U373&(FR[DNeOC+8a_SW7?:._DQJWK[Y
1PJK):AbATSV5:W&D+RZL3>O@^/:/AOef1]2^,<UaDJ>Jb,-DGZC51+P5Wg^26A-
]9V=59K^T^<9R]?^BgJ>1.f&#6,LB7Z5,1;)Q]T<8bG>]7C<=Z;?fXbH+?4K=cf1
/LL1#_^gOI#WJ=(XXVI7LUfUH1/K4Z^EcfDKB4fdgPVfOaa.ZR\BfK_G_5J#<^E_
C<\OFf(<1X02QV+O>:##26.[@#R>L)G>4ZE;QGQ-bUZWNgEFQbERO(3H91g>DNAg
\:2E-YKAQ0&Q,T?6(RH,4,bF6fb,c859OUY3)JD0GeFb<O\K279V8CP]FI/F1S_R
LD.AK,PeaA@&@;V,I&X]E#8-bQJN#CT;\3FDb8c:ST@Q3)/7@eG9\R)DOGZ23[8e
&c\Z\dJRb>X@g^O^T.NC.EAD)\7EW(?>Wg<XZYO3#HS+PWQLWXR)eZ^URB5\V6g3
S@Z5C8_&OSWJ[XRUgeI[f#0</A/P7DX031A/3@9IQZ<_9fB1Fgc-fTZ@FHIPV:Z@
NBf:T2C6/DA<DH@F==3U:G91VV&)&WFTUa@JOT^)&>X#?_PSae9:d^I\\g9V&N&B
Hd0dRJHH)(3VNN+T1g:M\+fDXOKGbTf(OY1cRQG#G8IgFX49,9Ma6Dfg=;D9R[@K
4a829.ef>GE^&RHaAMg0A;,0@:S=f_G:].2?R1KQ6F0GC,B1S<S-P=bgR.8XY@c2
\C]K.<,1K?SYEJNaPARTF>:#WI./,S_D^8E9\YAP^eOLOR1L:SO573ZF8JQe^A>V
+E;BYeUXU:./_-1(T=J0Eg6.8[K]..V;NK4c,Jb\@&K)AB)&+?I(#OHH>K42.,B;
G^>W=VWIc^bIP,=5J/Z4WQ5D;@N]F>9T7NHL)=,@2c50DUEdD9MYVG-IF53PM_Z=
+aV-6.1JHOf1@HAVgbA8b,M+;G5EQfDYZX51dD?1,?8G)PR0>@H2Y1P69Hf/LK_;
fZe7Oe<CJ1#W1=)Y4U?T7\UJ/>8SDc6?R/-+2SWMVK>TK,39]g)E/+VTM-6PT/\/
g;A5\\=-LXL?=HS0=4fMY&BDgVUMTg3X3F[CMJ&NbI;@2]Qbd(_CT6gLg7[XbOW]
VWU>32#GG@feSEaWFM;dgVNGEV=805W=U]8N&-2L5g7AAV.7S5O&-ANL5:#4)&a7
,RQLd3RV:RKBfg&(LY,Jd&fgGGLTR<7K&EcbL_G^Q5(G]/_;@VeWWE1FR5)HKLGV
=7JfgYI#HO_UHN4YKgEYF>0^3+V,g<R^M@K\LcOd93RHP=Z2&U=R.W^7>2b4@eIA
=6&DL^Y,8#1(E&\7W12c,bSU>9>7.I[DeBWTgQ@1QeXVg/88Gb1[UI1>aT2R@Wc+
b+-Z+=fM:9B0L4BD[H2:G(2&^bYA0@7\9N]MJCcO9RaXNg45<VVYY&7aL<EbVA>-
Ia@abfHG&\;8/KbOUGfIcG7WA3KX?3,d13W[Xc,2+L/Oa#SB,I7_FNGUf\:\K[[;
M9QP[_]]TJL[O])O2YbW;?]19#SJ/?X;.LdANBVNIgF79G5dcZTVbJ1W[DAeH1U-
8(Yc3g@B(T\ZL7)@3C9I(<PfEI6b>;?BA0)._.:4D,//J1SW[C2M5ZfR5BAd:8EA
NJJ8TDAab=<&cAgZHCRA]UKENR@^a:SHgdgXYBW\J);WYcES=H>UFV52g2J2[cgY
X2_Da>\HRUQ8;1L<1JINf461-N8K._2BTY2@PF)C;O\#X]HeT5B@8JB]dfZ#<@HS
^CNA^@a\CJD4@Q@YO:C8&\@ZH>a0db3cc/41CJ=Wf;B7)R2P7GW7VM.;9Ef&H2MZ
LL.fTIQ:\+_KVU^P.I0SNMVFNU_GRc^6EX;C:O8I/Ec6fQagS[H[+63KTfZ]-^IQ
+9.9/ON/+UVR=V3:MR0F]).^7ZRW/I>P##4FW#PSAX_CA)VBFJDC1-JNg7NFS#3K
LC]X9c=2A6,;@Id+Na/>0;M[FOMgb,XTHc]<?&C9?Y5,Z\;6,N79[2(@#Fc6d:3L
]AD\(^f32P/(8<WB.-bLV(;eUS69E/dbJZ<,A>KET94V6AQ_Tc&8.0cgX\RJ@PCA
H8;([.#[FXPL?>()N;IA)[Ca[>\bBTUb;PbD]b]d;9M<G_g/WU8eT?&W6.H.#W7V
HD2.O1[_4^^V>]+F/@27<HdIF@eAF/2GdO1HA=KH(gRcNB5+]RORLf3BNcC_T<4+
\/_PW4Z_([G-HL#PRK77JX(0aAZ[]2H;-JCE#C:1,1CZQ#N.32^^O7Lg6^VfFDK,
-YUH4Ed49AW]>D/P7Cc36_eKgW^@@X;fNPTQ;_/OPf@7&)(L4BA^&758Z(d)aU@c
>-D3._#A@TSKSJ7[)70a6E8Og?FO=9:[CO[6&@B/O>#2e_W;79KD94]g[Q/OT4M8
S(:UK+_Y0PW:3D<]8Q_K/B,E-/T53c5E.AT@(T8;64[-cU,AI1#LVWKS[X3b44a3
^?bGTXU,-#cJNXd0B/Hcf#5RgL7G&5HRdSKdTaPMYE8RW#P)<_-Z;,=KD8;9b:=W
.RA#U^,7>7eBWPN^Q6LC)9G=(gLA&D5g3.@NHg^+W)X4XN0.T:Z0c<.N>=c)0=K4
>Z0eS7VG=:GQT[B2Q-7_d08QNd)B@AB/EPBJO?bR(VQg@XQI1RI[HP3_RCVU(cIY
T7D5(W#g+9WA6+)=K+0UM?FS@\J;..-B7KZP]?^R^O54LcIA/O[b::MGI8=Y2U7[
T#?ZRAe\E)R5;e5<A)UL:._[CTY[f9cf4=.2G/0:(bM3#e;f_CYT4cgcJ^PI1NU9
;-4(Na6[\.eD;0;e]HQ09c:>>W81\E5c=4#8N0<AP6\P78J9<WPJ9LOTV4]URPb,
Q(BP<JC#TNQ^=(QVMLJWWJQ_#J6UPA&<Q^TZ:d(_CgJNbS7e0N-HVQPa-MC7N5Y?
d\8F7g>N:X=.QF;0AXCfLF@/)SA9.fM)@6Z5K;5]H>a-cI553B5D3U+Ke375]QF8
<0)=UW7&:]TLE+8)EOY=aF?)8UR6dB<>dE>?_7=#VcO1P[[8,&B=F/.^:[>6Ob1R
PM/b24@/F\KdDc3Y#P_d=@[&Z@PJL+OPQT6fg2P\bQ+P)#]W?PEN\X04b/Z.-f)U
]G_V-fdSa\)^LCX;Qd/@]Vf+4XLG7</:;@IBCca1:4>C[X:P#Y:4?H[,\NYZ1]]&
.J=W3B2]((+0=?gE9@8b#>>A:UAZO<[=NII8^;]fET0SDB-#WE&)8GUL;,TLd6T0
D98.CgZ^))(a=,Xab#b3QeB,ZEbaU1^cM6=ZK=S1N9H6-@#-NdRV[9,5M]#eeF@P
)KE\db<F[D<&^(2;UgXDV6I:7LO6f-BcXLCA7MML^Eb&IdIJ_#VF6Kg>XJV>baI#
@PA&LS=BMf]CPeS=fNB]e+0CK858g:60:K=f87dS(@.N(Mf_Z<3.Z;\eK<2:J^)Q
NT<4+BD-F21QKT7^c-#GQ\,;gg9:Z0:A,1-76IAEe(]KRD[e98bA6(TK(OQ+<A)[
&KXON@17LRSB_.:Yc+-PHZfe,2Q?HbN/^b<<Q<0#^b.O[]K3Q(DSd0Ga=/IQ:JCD
M:NE[P-Z?5=7g]/_9>0d(Y@M:)\B^6d@\g=(:;g9;fQ^7I2+:JE+(\NA5HRf6->&
.<[dYX]e#&(cRL?#BdcgcP/^b,2)R8d,P4gD<LBIQ1[OK,GI]IG]-=&KUG<,EX_U
I2-9U<L5JFGOB=UDV(-OY9?7PS6Z7<#Jc.D;5W2YW>PZ+\^+.:.&+/7fL7>4EAgB
^-LO+2R_L:;2&5FRZ(/aI)>D2]#AO,;.9eUaHgd2?<]&C7[@:_ZFPK#E>&Y+?H)A
V-a4JK9K50,eN2eZ8Z/A_Q]W:4bA68J[YNWWAU0&3b[AFJMG;OL9V@EPO]QM(DJA
I_^5A@e_4X)g.UW0#]]<^LdGE6OX5?=16/Z#1(,3=]JKI(\/9cb2??>8T>V:6d<6
bCW7HUV)2.K19Q?SYE:JQe4JZT6DL\)g)7LZ/;[B1TQ#A4)bcY(QaCY/B/9b3&/?
LPW4d8=>^PH1b52Q7OHIL4/5Ya1;.HI1J24BL[V:]aO5<4c0BeQ)/9U>?&SF]HL>
X]S9C8F(IY:BQJK,S3b\Q_9I=^6I3/X:C@L3L+I4_.=EbSG;IJL#A2R08_A(7AB7
H_acKH)+B0VKKcLD=-TYXB;+1).UGWU=+\FB,]^-;aeA\GeBg8N&#WVAA9>^#KT5
&4ZZD[VNJ.-\#0A0cO41;d+;6f].E4J+0WI;Ue;RHdR=BaOPP)N&G##=J>^fcMTW
-2bM<.:BAf#-FUW2C4\SaeJ_S8<SB+1)YbI/N]@22276+7R0&Z#3;]JSMP0E-W?+
8/g&6DC-SgWb1_A6+CXZLdU2.@gE+Q]N914.D\XHMJ5P&\d9LWT@XQ?ZYZ\XQT3^
Z]G/.3\U@8+8)36&^#JE-MJTQZ2\Y-c[-VV3^PG,D+OaXJaFB6>SFRN+e/D;Df?H
/UK+8/=:(eV^L(XA+0IAHRe<8g6]ReaF80@+]]9bRAQ\16U5RQF2I^),[+Aa3),X
D:/e^MSOW(N:US74STdg.YQde:g4/X)=AKKeKe+AIggG6,]bS6U^C#H#HM#2X9d>
;JGE:\<Y4eTe\93@)3QBFE1ENcM-IH;f_W[cfXQ=IC2KEQA+>PS2,;TGM&#KZRH^
60Z8/e\;b+_];>Z,Ub2/5YM3E6M5:6/>F3/XBY0M>S9\-_b&4;AS^UY:&)[YAA5O
@c+g^ON0-@>2E?&:2RGgZ?9P&OD;4/.8)5eTaAcN[UT04SD)/RFcGWYH>>0AISG:
b@-dS4I4A=fSI#X4aCN19^b-K556WYB=[9aG3,P#?>e3-9+JL3?]=&-)OD=F9-KU
YN7-4G[TGW9>YSW+946BU8D;Y&#(=7]QWc/^D@G/O0ID4aE><95<L#I367SZ])GE
QY&Qg6bKS-Oa,;IO[bA,88Be=\=OS807b&O/QIac13^4HF]4e0acP#:#4O04#6W8
E-]MUVSfeJV]7@Ke+F-_/,bI=S+N,:-N)S]^ZG1,_N0?76VS&CN8^:PZ8[abgbO#
NA99^NI@J=Cc_8<_b.Q=]E3Q7UgABI(\/OF98^7@+dD#]b:<:([/5<MQ)/AYdOP8
7[DYTD4<<])S.f.PfEI[U\;]L?0QJ5JA\ID0[)a;d7&O(8]a?E^_+/F>Ed\^@X7d
=c(Q:YdR;.-M[E^Y>A7NX-0><=.S7=_U#7:gN],Wd6F0S2O1Z\VR=C_BLKI:@+/4
4XHS<R1Y1E)/0^UD#8P39BAY><9I@5C.CRUK^IbN5cFFL3JKR[5f&T>\HVA0R\RU
53]1YYTUbSV3()P405/-G&I9PB0LID>:]b1cGdfcPO6:Nf4E]M8]H?b(\(aeIEIb
_)dX2Vee3/C](L\bPd-d.deN]f]DEPbHH-.-4aVR1<<1;C-\2=T-)-gQ/[SXcJRY
2&5a9=AIA9;NZ,,VM)P33IMT(Q?cNRR#=IZI2RE:0WE^38eC<c#)8<LWP5I13F/b
8@W_<8LDKd#7gRHc3g,dY].JF(K<@FP#O10FE&Z]V(;H90H<R,)\GZIOJNKDa2XA
-;1ETd-NUVaC_,5WMe^a;;I)9Pd::V)g1HOc)AV_aLVDB.JcY#-dg=SBVUf[f8VC
TI=fA7:<a]:?[FVJ9U>B8#&a0PX?6AUSaT+XG_>:JFLg^??ZZ8&eX0+N;OcY<G2R
-A/1&^(=ZdM(MH^#4WUUGA7@C&,^>85I-X&5=S_G+<T0_\0>BRM0W_f1>GgR?Z\2
d\<Bd;U<ZfEYB^+_\V[gJOg/@B8VG.Y)O53+(W,0HaMGT9P3MES:RL6@,U;(W3&<
,T#bZZ+(+8F@TSRW,?+K&d6B7eHCb8\J8]_4X7c,Td38.1;20<JU-2G8]3U[e9S9
[ObDRfA0QM;dEH24/&>RFDW08U4#/cWOK-SM@GJUHT?5(cD&FW5A_:QfRPIdHK^0
M>=<^7QW-?3U^ZWN4]8XA][J2E\Bbb0[,O\26-2F>#J74bU]GC7HgIHf<4&QH&DX
6;#M.=9&HVFR:)9Kb>\@9HSVb&R(MdWfgS9Z4MdQ70&_G+PN\I6bB8?\&Sg/;:Q>
+fNA9Hf4Lb-L:QAE<W^UTQR52M.XPM41TfKEC,\XS/D_H4=SNaSI3/]bY/,GLUVI
L0BG,4N2PF3FV7aA16Y[R/-48AYJ[d7gX?97aMf2SV)RXSZHV.9X-9:0g5&7cL6A
Z)KWJ\D=9-J_RgTbQdNM-]ADK^R>.)T<\,?39&U,#eS1V6@^_-gXP2,\F.cSAW\W
6V#ODWH(]eQW9C2P+49#_6N8CK9RUOG;S+CFM0W#>.=-UfH\P)1Me+KR=L:Yc12>
W@dXa.HJ?>[_e=PTTO(U7Z/^KVL;b@9b4].dBGWCd+]bDNX4f2BR]Wc+0<RMGMH#
,@ffKBTdfcdGM\#dbeUGPbM?/S7HZ(@cB#b>QZ@XgDY&A1b=Z7&,[<A,VD;NBSIL
O=M\.5X5OUXY9QR\@)2TZZR3][=f]BR2W17_3,SP#+<gF2&LCRF8G740M#.ge\c)
6P8c>E1:Q\6A?]L,\)[cK<B.0F9S47g2IHW</S;/N._9d&.4/SX[K]YCPe=Y:e)Q
B_fJAf6AXU4I1Od>HY^V2_:/1;?gEUdB^,X>2fH=?AVLgY.[4>6;:+]eH@fRR05Y
/-NU,>gZ4b[[I3BD:&@A],<.#?Dc33YAS^XbH9f\I&N3O.cL\,1MZJ3G@KA0a[_M
([c)46B=D(Yc#fC[W/:7,\6XA@Q\FG.Y-04N7e1ZY\QM&Q)?,/=Ra<;_DM=Vd^IU
J@5(&UL&JW6^(4M2@\/KRY3@Pa(X8#UWfU5VPgN?-=Z6JMCDa_E#Q4TM?TV2C5g3
/?N/gA>1bU+8@Vc=,b?Dc;-+U5AFI3>QBM:K^M]/1\[d9MgY:@7G-]NP=](DB1<[
-c0NP4PAI]2=U--]ZT2[CD.e6(JHRVCdfZ-A5FYI3=H7CB02I3B_Qe#I8eJ7S/QB
L,WLP]^Y0&T7^(aPYB#)VA\V2LZ34#O_bSS0XbCg.T32AZMNW4PG/G=QKZeI8<4e
O-^D?X>&\MLL2Rfd24P3/f#4:93?/3e5Cb69^B1[Ug8YUIO29@Z_FTBXXESZ_d+V
?H>2V)4YUIJ+AHHNL:4)80:J9]LM4ZZDeY[O/gVM_<JO33-c1AO]_c#X\cQ,;IRV
64@IOP+F;Bba(6T-/<Ac@IOQ[157([C:7K;\L^ZgdXM:3I43,c/dX@/PI-<?G@SV
:BT6f9N3V7:Eb:FJ:D:MM2b+B\eX_cf1SE)+LV:b>0[46UL,1Z>5PQN)[C:HCS._
f&/cZDIM;4TJRCCab46gK<\_81,Bd5T;@fYD?<)FE2(5VE#6RS=O_&OME##KZC\8
5)#.I]I-<c:DMW-MG?6_@()NV2F\=X43(ZV8JO7I#]ZL<8OVI-GQ7fDW#\C04);?
;/N9QHQg?7>-c(&E-Iaf0b/\[<94_@U3b_3fC?R+F<&c&5WbBVD#[Z0B/_\OfJb&
-NW^gQPRKBZXRF0UKIZ52[5e>A\CI_gW>e4+;VW=c/D,Ea#FT6f);:^H9e]?DZ,[
.ZN7<1>#gf.FUdIgc;006Q89C6QfL=23E>2JM::_VKc5&7<>_4)WKSddKQ?SZ#[]
9[H2V^d_EHTIJU6&eVRYXBbRb>\bgD3Q)..cJc4QG88SW>3,[PcZ[06HY+Ed]/Q+
/7AR?1-dFLWT;7?V\N?<H1gaDT[<Ta1/JP.A#@&dc<[2Cb,M&\HaYH2O@YV9<b]5
;#Tf,RDO<^E21>\RR&0&5/\0J8P?&gN]_]FO&fH4LQ>HJQ[>X[V?-[Z14R#3cWM\
(R&BW?K@,c876-NDK:W;H<H7gOLL0J)eN.ADD.-8CNJ^BF7gU^Y87<fSeK6&T.N4
@9PB1N7f2Z1(d8;B^85F=H_#@:&\:T_EGOb4e13\E4Gg89^^U47;AVV^N)e1:S1F
<)Z+DGQJ.U0DIFUAEb<WR@9[#Z(EA-/J8\E=@?2Ac52c=S?e[fZ?McB;X)bRZ:#E
0,,5ZWHO-R)61gZZO(WScM7fOYEG@&aD#RJ98=:QE]M=H;g#2acQRdUJ^c:NgXFA
ID28]eb;CPYQ^Te2KGO6S?W+[#T4,\6\47->ALfVfU5LV2VBUJaKS]>)2ZFI/P]-
3XC.CHM]5JAA^3fYfP\\X>RT0]21:Z[6O6f[TS-.a=<Y@C+^_6YXdW-B7bD&Ne<?
F2JcN56V^JA\5Y(R9]J-fN3V>G&[+U<@240ZQ)cf?Rd7>.W3WR:L,?\FMd2P0a#B
a@[YS91PRGCH9627S[>F3?NYC,fC?&U1R=:\[IA,LP=@\0&<P1)GF]D/gIZ>+<67
P=e>6H7W^KGc_3&QPPN+TF>VR#]6VAa:WC(8HX4c8^0SI2_,F6eP.d>=2HOg&I^;
f2MeN912[M7G01D,O.47IeK4@]RdJMFcW.X/Tf[I](P#=\?.cF^(#?>gRECB+P6:
Z.H_c-&e0HcAO)D^Od\g)2TLQIHR<F6EHWYb;a2DJ[V?Z;.)V5Re/Q72e?,:B3-@
RQ;AT8/@R)/-G\8N]fR]S8CF;2,[3+,D.c?B\UGKD#BH3d=5VgV\A(Qf&^OZYaE(
6RIb8O_A0gN\C>R6@+(6:Pe#-Ja\6>SX+_C-QLb1IdSdL;N(^V2.3>FIE,ER\UX<
SNFW>2S:[J1YAGB3C_-1#V)a@PU7]7DBf397UEb]37MPU^T7:PCG/dB>4gcBD0=N
&@SWY?@KQ]M/5J(3#e_L44(DGJ1U+0.aU_#(e#5aWN/fYdLCM>B0,d##@L6eED6X
&D3T^-@Td<D,:=R4;;EHM6P]?S,3IUMUF]0MO.5E[4HUW#Y[T>)K2/W4KL6<^A8e
^aP_T5debW39N\cR4XK&BMGH&_>P+@A6QP9:Y7>QJ1a.6)(R-[)M6g/T+ZO+BR5]
:.f9c9Agd4&4)E1)Re_RH3NT10?_cEa_&fV\D^d1>]g3Z.H+V=89a;,3&XSb2XN4
a7F#8]aKZ@bG+5fb6\IS81+g;H2./]\VeCe#=+I6Be>PO9_LcHE3>PQ<FGaE+4AT
&>EV:U2W-AVUGZ.T5f.T+[BVM88c0dZDQ:CbQ.Rb4aRbL2a&5PaYe(0a@Bb;c618
R83+27K/0+P._b.Z9K[ACKB=fUGGRd\TW#T1R.=-dbSZDSd;:?NgbB6S@c_I_ZH_
9HJ\WPNbLVZ_)7aY?0ZUWS)&<8f4<S=+K9P^eI6)Qe^FQS_7OPZC3QdFZ0c+9^TB
3=6S#1<\e#eH.ZC7:bI^B=N4PU[N5H/;[<;d@+e-;WbOBB4VQ[HA22eDCF@H.BF1
gNJ3?.F5JKHR&JB@He>,88XK)/L-OE.XXI9?ZS:=ZAAA7F5,EZLAGa9U)=?&f_6P
f:A<H>bGXfE)IHg<f695-L\9Zc?]Ud)ZQ)TB:6PF4K3=eH9)<_PDH3=-SfVUNW&c
[/_:?2JQg.+VEA7c&5?].OQQ_9N^,H]627X(IXEVNfF1a[/.G<R6V^)I^MYW.?BM
JM,/EI]Z1?FL:V?C\I8E^#IC),eZW+BVd:A8#[H=F.=.-T6c-F8+33c@PR+RB4^(
P4OBP0Zgb55,DAU_(>A.F&W[.Xe;?N1/I_R1M336>YVO<W\D]@^c>(#V6-b2,&\L
>?F:Q1ZZKZ=CcMeU-D4))+0B#Mc#;_#+@Zd.33.0PF.-1FE#1Hd1&=;YT5M#8Pg7
&_ZQS=_R1ZL-fgHfXLC_-C7a7#I]&\1@.H(NS^6>b1V_MMVOGH[M\6I:;&/5\+8V
CO2b7.XbYc4J/agcXU\+[5AAHA?ge?P)BFNQPH#&/8JX6>+5\5O<7bMD]BWOW.&6
XU2\925NJV@=+5BVU.\6>PNM,-5L<c<Pd.-_&6_4@V+Nf9EG7XTgJ-C-O\X4g7YK
=c#_ZgN]gcHWEF-(V8e6AFV;YY\HJ(f=d,VEN5WP\R(5K?e_^HdOEccLE.:,3?03
AE4V;aI@7G-5a2/.C2ITX_CO(R?dH9cHe<AWf#MdTab0=MDAYf,Y^T,8ZD^#c>9E
gF7(DM>L7&=HRO8\0A@\[2Db1)H^T07^(=,N8S(BLO1&OcQ&(<<eDfB_^TG?VHF5
HXX4XSJ;e&H-YZMaQ<T^FR\f#V?:-aV9(WgNf0-G<^GggN_,84PQ9&d4FRJ+P+g;
OV(-#X-]^c(>&U?ebZ=#D#8WQGDZXfO=@JEGQ6+?7\)H&?c+^UaZO:W-1.R(bZ(+
@?P<[Oa<IHHF:LaEO)6]0cda)A,eB-fe&,7&a\MSB1GMKcgLX^>@+&d8<_N#>8,;
?OYV<FHSA8f=&M<O/d-]eU&@8S]GY:=+#0,D=ZY;@M@A>0c25<A5)OXWY-H?e-FS
:-C-LY;\NEe;@NbH-Pba-.cU3S()2+BGPWBAKZN=[_/FA\MD;#,__BSRaBd]K)/T
<V#T-<e^D/95.@^,7Z)0D>9I<\+B5;CA[B7LUO]RSG]^;K\ZVGg+&\fe.(K,#_P0
dY^\4a^V3NC_CHX]Y;]29C0RIZET1SUNW8W1OP5aUXNX:T5@1XB)_93gA<[6(SH(
WTTETdYDb8WY_[+Pa+1_.?WNcJPR^FC?XH#TgR+0Z7M]:7Y,#HNCR=c/ZTI=d06O
/1#K#cd<cJ(]<0NaGdPLVf,O[(bG]9YUKA1R0,dEe@>U<.d>,YCK.#G\R2^U^/BN
@4G?d1;<:??<L4d.B44O);?^@1a-1LWQ)K_](_fDdTg3MK:1(LH2>DdP+>,US3A0
9&CC.MY&/&>AV0a2X&I&HN87V8)C1ed591D96g22K_.<=N,38WaOHQU<1g4-Rg_J
-7-1efGGK[HSA;:28-?,&c@Ia0_Oa\Z)=4#7g<g+)R==BI=,E6[,G0_Na0,_X97:
/^/ES&CP>+7V=EB8A,bDI5?U\B/e[fL9d<],48;.DKU9#TCdTP0VE)<\U_DCf[A:
)LD1CXG+>H_1fK?\,P+SR<(+L2/.EGH=3RZIC0X#ISLMfeg5#a:>XQYQH=8KVR7^
c-I^C+LA:bcF:4U_XL;W.:L=:I:Xb@f?:Uf79LE(C4A(<+0/(ATYgg.>NZKBJ]+Y
2fR7FI3cU,]ESO(Y?SMYNVE89^a;&A9?d(fe<^DNUg2(Obd3O#;QS(T&63>^(Z6N
_.IN5fP-egdWDVD<b2&4<]N)TCEV_.SbAVWd#QG;(:]V0@F<<?_RW/_fcQ#bJO_O
ES80B-13ELVV4D;;W[7ORH26XD?Xe(OggIPg7-g^EQ5L;;3,><=9T2TB_.+2g8B>
[7#-H2?g2;9/M=U@X-RW)\MKUJ6ETbTCS#/0YdRK37.<NOI]1A_>gY/S-^U80W8Z
G6>7]]OGX<)HQ>1@FU&X+PaCAMI9LeS#,BGM6-KMI<^TAXYP=M)#e,3J\G6g/\g/
T-]\fePgWfC+0JKCXYPD-00XPXE53a.Uf&Z6Eg\K/Ze@#=1(_c=Y-Dd_IA8GGZ?[
B:]9B^aOF+gJb<L6___O4@Pe>b=g&I4S4OL\POM#(KU/[LfTM346YU?KW/H1Y/B^
;T@GFXI8;1\JQ9S(/_H.Z7GN7<e#^:@V&,296g<().U0G@YSQ\;b7LZ.-C9?bf1C
1J@A_20f?XIY&FZ;OcVEH]#TZE/4_cB9#&,GSM6gTdg<PNWcA@+gI]O(VJHZfDJa
1(+J#+:U1E[SOGYV>A7VDLW]W<O.UL(9P@F:\85+-^CI5bX.L[];8V&-).,PTP=1
&4L^6>@X[](/N&Q&PUD6^gdQJ&Q4[?eMaFL=ZQ;.AN?c)-9Q_4A87/XT/XAaS3X8
KSVN/c9B+HPE&1c9Md2==/B\1D_+A5HbC>Z5)W[O^.0QF&SC_TZ2,Lc?a55R</CM
HEL^5+_:[A^VT)\Q5J0)^)g@_35aPK)R@SJ[4NT[0-Kb4C7W8bT<HB/Y>(B/dIOG
Rc/J4B(?R&DJ]@B88VV&YA&-S=7OL^V58G27M#a(,C)K3RAeGE34;E86JP6Jb=G7
cYT=WH.@IDbO5+=a?(=X)]50HV7_1gV@VOf:<9)J^PDBO2:O@B[[0;We2H&=MY(?
L2MN9D,ZOf6?J7>d],PMKK:]XWN0JU[PRRUU0aI-d3e?eXf+cf;OB)8Z14YDA4<c
\cEOH1.UVKeD>C7EW(NXO?9YBQ_X,D9I2dCU9MPEEY?L8OZc??ZF5W/+3_fOV9.f
NMEBg:0;T>@MdJU:0H([]>(V<-VRRH6CR=EK/Zc;-9,[_9(gdSKLJ<7F<>LSD2B[
<A;1M+2^B2M+ad4;;H4aNRQ/,;@Fa:(CeJA2QW1TLV:>dH(eQ9G\>--;W-Y33)ca
UEaK9N)IKddK<MFK54-5eWAN)BA@FgS:JAW14MWW1V>0_Rd5#gDT1dMS7B?=4@D=
3OfeL)]F@3P.W)WWbf\)-e#@f#O#T?F9W_U(E&Q=[H5IB2#_;V#f:F^?D.3O4^.N
R7;\U0E8Cde0dN<57fJ5ISS,63_W3U]=C(5=)NG>,TY=PJ)GZW>P+YGe/=?W6UQa
_=V(eK1G)A:a#/++WI26+H?/WUHZD2eLNO#]08,BGOKS(ZVHB@)c280R8_>QZgEH
H2ZF63RSGFD0QcQ?RVZeRI)b]V]#E,1:0>4C=KdLY+05LN/J^#VZ(?1W]P^@4^?I
N]CcLPIA>K>?DP/?/;gc/K(4d2dfT\D9fUM/A,(@7U^B_^T#a=4OHAIXcId,5RN_
.)P^SBD3cc=dgf#3;8ZV4#@4Fc8#F>KFT)>\BWdT,P)></FT8OG5GD;O=(Na1C<A
<2XCARP.d7[cHIf_L^OL<eIeJVaO,H(gW1V[[&f?YgM611E91WU_)4Kg],:HYBeR
N/@Z0UNX-N)5F/0](CTFF+<3U:ZAe@;RO7TG,K@eaT=1E];NDHadS3EfLb_PI_H<
J.].\,a2;0:I=ZRBHDSGK,CdL[\cJMHV04<?KVZK9#BbLO#g8-QZM&)FaKEVB2-,
:;0JE-A1UdL6^VX@g)L_PL[):YD.7C&&M8V?[c6..4(NNMD8.5_U4&.6AJ@b&193
WMSS@_XZ);73DR)Q#MVgP-&d?]gf((,1><-fXeK&ge1gQ(99TaW1Y3\^&1UW;#DN
VUW\0VgKA]/IO2IJMQS.-]XMeIH0(UZ2SBf[2e&5GX#e,563d1P.L;\6B10fY=#9
3OS4Y+dNALYf(LEF/&&+S831+2F(L_Ag(/>/3(X:-ANY-bSFa<+A2._/0,6/Q0_B
RJc+T9Z\,cKH?+d1;0.TUe>L<D79;&)K8;Z0IR>(#K@I84N26=cCa8F.JW6EZ4:-
AV[P.(HKM<4a@CY?8M4Xd;C^;be13-OT:103^#F11H9RPXVd8O]4^JUgB3Ib3:5N
d)R._?;3Rf9M8#4c(fSFfO(WS_HK_\DN2,CLaG9^ef8E99JX3ZJ/@+(6CAL+3<J0
8RITWac]Q@BGL@;O+ONFUAF;,^<?GE-CB,@(]/4[W>4;&UOTDeZ+2959OBX#//^d
AfJ]4^G-c.#E(KAF8Kf??XY4d)1(]4:24>1X4];CJBdD,-5:dG?FR4_N<H3V^<>?
a,&7=SRL^;9/JfE,E1@f1f?-5ZbWbaRQH=.&-R-D,FP]4DI4N=d-V0e0TR+^P-4S
V4>(0S#_Y2<-5GaQ.Zb[Fg/=4FX_VB0&?gE)UXac8I;VKV(e09(E5W(44WI;?3-1
+19,,K9@I8P73RHPQF0a3(GMegF0:_H&;=ASPZ7C7-;7OBb=BXS3Y>cT:P-=bd6Z
I3KITIMUYeRPYBE>gOE,-:ZQH)>PN@F_@DCCL7#cS#]VNfH7OW9-S=2:-)OJ36g3
E<Nf7]a#UB3>GB7^d;.X]A=]_5Z3BVdTd#-7OVd+7?(ce9gR[5.ERQ)V+2>+Z4FJ
fQBP?T>-[9J=47-6dC#9a6baV0]DcAYGYB(eYHGL.6^G/-H)\6b8g^IH>@+16-.[
.:RXRbGd.,:=&;A9E/MRUB_F_+O#=W7XF/-JXXJVN8:4_&ed[\Af7dgU,#UQ^I52
?<GZ2H-WJ#R^.;Vc^&\CCG0eZ[[gMJF7@MA=&-E,[.BYJK3-V.HaZB=(;XOK.ea)
fL]V0PGQ:MH1<HU.LK:JGCB-7d[;,b&R6+QC)d+VK<#g6WNBALD@<A:1^<fbJ&Jd
b@6VD[3G[.YVC:U:HNABMEE@^[JHe^U[AJE0Z9O00a@LRX]Z\c_86JG>2^IL:/)&
4/6\(-@H_^H<FM3A\^[0B#-JU)Gf8T->C#F-A&/bQ:_(4][_1FM/bF_@\cU/F,;e
VP(7R5>#9P3[[&?^0g\S;9YLU-4MI9eXg09g[f&UC+X.d3XYb[D7PQ01f8eZ:Wf;
]<SZBER9Y]HU9=;,]@9VO.BdP2F02NTJ@J^,YJT@]HT0QE723TTTDHJG\H+?eXR+
_(#7]NY6PT\E>3f5APc322M]3EQF+)A&M1N-GH/.8,,U4--Bd]1)^EcN]S7HR=K=
+ZML,G2)6?R_GDYJMXg93)D]YYf3)dU^eS=J9T9SAef-6#cb#FDUN<K)c:J;,ZOM
,,TP0&)IET)O.[#=>E>KZP-0WUWH[2SF]84&,bT-I-V;:cg5(SbY#I(7ZSQMY>&?
:1_1Xa]RKK_Q:V+85?S(5:Z&;LJd,B]],fR)gDBRR/TI_[5+J1Z^(NJ]4@@DSAd?
JE:1&CJ_If)W6g4AD-[)<69aO8c]AH.YLVC#VB+b]0.gSGL2)4EF^Y]R=R(.g,AY
a/.g(9+1>,8)UJg7/5,@C/eg724:3a&<M?fK9,_Mgd&[AS4<>;WEFNUGEcb:[ZL8
I&;:5PRScW<b98UZCW?:H2Q5a].;4I_7fI.9MDMH=c[WEV1AM1B1_9;eI/Q&?61P
JcgZK7G/C[&3R:J^d]]SIRE=JT#)DEE1-b:/DKge4]B_RXR1-fSc)S<K4(G_]2<D
gSZ^)Ed&PDU;@PZ1Y.P/])b<L7b<G6UIE/0Hc#S]X&2f6O:>(3P2<Y2HJ<55GLK3
UBCN0MPB7KWH(fJ7g_^&R5Q&)d?.UKWDQ328PggXfD@\^@4^:;VK72DdN+G8^QIU
TgL#FYYC\,T<(ALgV#>-5,/HA?d:<06^KD/_VT3],V2fbE\eaH86<;45TDQH2)eb
4G4dObOV6?ceV)=\86JXG(cZ2EQ7IBFOUQVR2H;@aebVIVH=3J]Z]g_GL@N]GIX.
^K/-\^_?R9L)@:_O+.^E;RW+0-BXNA:/Xg<A0#W@:F?RJM2V<5(b8M>2ORAY_UA3
P]QLQGg0=^XKTM6Qec.&G:I19_H.>8ITba8/VNZd\Hg[WG[3PFV.,ca:&Ge<0a]/
AIE@HgLJWO.#T0;5aaB1=fM9CM(63LPM--&\+R?YRLX))B&KL&3Zef/]Z-)Y.F?.
,])B9GcAQZ/T#PL25S4EO5JDYMbeKJg=1gaYJd-;>R.YLBRE?1D(]JKV4b=AY\ZZ
M09fH,c,D?BQV]TBIYBW<1X6]c3\H7EE(2U1P\WbFHOaAA_.N(RKJ&ZQ8#XTYOX+
b]&SL:&3\I-2K_d<JdN2RW,<QR.?/?b7G4)<6ZXG9EfMP/Ra=S[f82UbXC(KSQXf
XZ.CG0Z&9@]EfNbRb\1^23J?]5>:&Z5gV4H/H&2CO-g)UEcYZ0CQeea[ag3P?@TF
^A<]:3aa&@G2VaM;E_+8N<a4ZDSF08^1QcbYGO#IF+89dc2B[,@,EQ1W0dE,@/&M
TR?40Cf++0/ce;-#E4IZ#gQ^I?4:F/3UVC,V>[/ac(c>V?8@a]KP^;)B29dL21B[
_AWe[L_1>GKFBGfGd^Y[FJR34M<S7N@M.a5b/&.4S0.(,8R(.YEOUI</Sg&RK+8<
Hgb?A2(O-F()@Q]+,^SNf7)WIEdT-/e/0AA[KgP\,H(_B8MbSK2F9:H7/+&7#AeU
I(78-92Z]1G:XW)G2F)#XKEC<N=M&L<>&c^WJ1IU;Ubc/.9JH9MYJOFK73ZE:2<Q
9OA^EJX/4BV-2D4,a+2&[gLCb551V=aOL5V>g<WEYBN8/#gT_G#WZ)?+[6]??D(U
8B6S<eHNXIY6T0PLOC3R>OT4e)/XM@WYa@&.f)SU\JEdW@VTIK\C274Z^94FPFU/
eWcH?9GBH7D[1QYI3e>5V895=:EcBLT]McQ;JHVJ.@_U;?T7HWKaeWM-3?b<(/I<
fZ3JN6@1X_#P8];H6R7?H1:gV;5B.B5++D#14e#6FYO(KN)C185I_^ND(6+YIWOE
1aeIXB<#2e_0ES(//KYM]JPedFM+NOALFE9A__V[<.gXKaaB;W.<;ZMeURHJ2M96
D^F5_7\(;gU>Af.5,+T)S9F?1:)&G6E\cGZ(@IBN<DGMV-(=M/2W;9#g>,#\aYT;
F#0e;(JabICb7FbQ(&dG??Y8_?LG4>N<OG,_MXFP^QJ^D/b7a?UE&T+G3AH0J2=_
ABLE(C^\_/4BCVe,/\)VRLQG1K+5DBc#3)\EKCH.RS2RRZC<Z9SXKHY9Ec]^2,A7
f:/g8&Ag=HZJdJ)F7+YdPSA;6M_aFYGT7&BWRBW.;1G?TM:LVU5P[[&fC1CIX@V^
>0UO?dAJ(OWcHQPXf00YE>CC(Z#\C\\.4IQC0aW;3bXOB8Z(eA],6,]#X[W5+Rfa
/9#Fe[XB5E&_bP4:-CYIOUD^G8Hf,>2R<_)S@NL.(Y>;QZ0\a/MQA&[).AVcBgd?
9[1Ia#W:/_Vd-_;Jb<]^BNC@&bI;a/RU+aLF_ZPA=>g[4DI3+S9c2^4T)2)N-OU[
+^-f[W&&^.f=Y>BP2aSd#(S>2_O#:9[23KG=O_^=7LMdH0BfHX=BZ\:O8,f\cb5#
cM/-0/4[+F(E8)dGf/-ZAPIN^-Rf/COXKc9C-K1TS=\X&Q6FM&3;X673EA3^KA;W
QgH4PL>)Xbd[R&KQ><K6F5H)NeSE#_1gPTUXcD:CF.:63QCXLPd@:503=_<ELU:-
^M:WId8L#A8_@bCDQ)E+NU7A8)<=HafR[^S_8,a3a-4<+C4SL;_>TT(=_ge,A;8/
VG[+#3QZ[H-SJSM>7b/=.aDZU>cdd-P:=O\WXP;-_I\(5+B2R5dGgd>@L-)PgVX6
e(G<N.2QEW#VJ;&Q^<ba;IA^FPW:HI(58ETF?Af]cdPf4Jf>gC^\?WDZ=f[[0eR&
g-D=(^Y5f@5D\=_FFB.(CI=G;A.C9BCKI6L+VU=P5Cg<Pb^fF[1>):0@[H\6V_c-
+5O[R:Xf)W,[F<9OET[IGd]H3=D^;>(?1=bYSUO)NL]TLHLZgLF@WZY4H#/_d?.-
]XVUTFD=-@?R_&Ke<1bE#fOe;4bgH49@@856#0V:RJ&2?YEI8HUC/2<N>O[/HdJ^
TKS&:LI_W>eOTO/&9bPIV0F4ZH>fYERR0LGP.]bEC,d,K1-cE\eV0ZF]T+HB]UUI
\DM4]cM7V[,4H&W/4Hc5QP_)LPK4@7=K0^(Q0L3A][)HZ79c4RbQW20.OHMC;.X>
4B)P4L.6REM6-U.WCRS1.e21-SNPUQ[RDU9)W,1R0.=H8M4IE#&4C?<:&T/e_9W>
\JU\DF?J/@]00.48gMfS,aYabK>D7O1OaTIJ7^,R#M5NBABWC0_>]RW@YWZM,TRH
>4XSKAR2W2+KcO(F_Y1S>G3K89Z2IZQ@HPa1K6-[Ig@U>.[7ZXI<4W1JFBIFF:b+
8?g]@:=5S[B&\U-LQ6IJ[A>^^Ia+O20gK7=Cd3I7OV)QLT5Z(&4;>aC(1R(R1)4L
<C8@^DE,@PLcZP1f-^+N,-@\f3XWW5##1^W1fEH8D8-(#)+bc6V,L9G[>fP4>X;2
UcU3ZB<2I(Q:6<>NW5MM8^T>[7#G-PUO\TZZcSe<.+b58]YO+:K_O4IaQD,:[675
Q)cJ2K:4M#I&bFUbR>/_@HR=GQ\H[EBSZ0g[SLZ9SUO8&e99A>+JKT[QeJZAd#;/
>5A-82H;)RMbJ72N6.+]bLbXYDLSa:EfOM9:GJgNR>R?f?fDg]6/f/1@X6&&?67^
Uf.@Bb1XI>gJ77=WXST?N?E1;H()6aHZ:VBIdcO]:DE2&SP\3PITY[PKB+Z18H@+
_f97aM^;[8CU[WBNN^H=HO8T=+0)-6@HWf1\d+bMG&D:T@b9Ja>gQ?(?7Z=+(\aA
F/E?.V&01;WOYZA5>Hf6?EHEc.>[X5=9VEXV5=:&LfK,L<KAKPSf3H#]RE@??_?V
E>B[_JGe^EbX[,Pc6^AC[2b^dG5=2bD\;(TAZ5,EQF.+&d4L<Y,YOgR-fM]WfR_X
>c/:f[Q>O)&JY#PaWHZ+G4g7&0FC27_K#)59?Yd^Wd8Z;\3a+V2LZE^E7UQV72c)
Q-VDIL>Kd),J.T(7#6fZ]K7<fXB;653=Y2R+cK_WCW/B>:KM)ad([K06#R3/:\bN
.E\V4L6;T48&H>FPAX35AD6;e7=]#4;KRJ:WNRPG2IM:-QLR+a=GdbXCcg1.]U@N
:#BL43&Yc9eK1VgQ4:2F?_\Uf<J]HWLU[J:#MYAR6/#b1FF\>CBC-\6BZW/DYU9,
EJ=b(KW>@RWA,86LO5g(gbJRS4W^W0;EbX4:P]>[fB@_:F)YX?bGgW_dL?52#E-(
].I5d1BcE96dbC]KScc9E>deK,f&EJ]:&5F&;d0VFK>&)-HL?>>FQUL+df/LM^3Z
+J]@AUP8f3EV2I2P1:XGT<1G_41+(3e05E&TgFaNaR:B=MFd>6_7H2^=JgIAPT1U
T9U3+-F2dE)a&[SK7=9?A:/=5160L0-/B#QZBQ9HNfD0,g9,)K@IV)fM;KYc@[Q(
P_7WBcXPD01b,_[+(d90^\E37M5&IM7+Aa#d._3K:bP&D\bAF;WFJd0D::+GD&[2
0@=ea3e6CF1I5>Q(WCPd32A:e#9[3B5:[bTc(DSP-UFA8[N7VV5e;<&JBL^:2b1f
;[g.b63aKQ@FaKRbf:R?0#dU[;SKWcUL:=N.88_>DWW+5]\N<WfJC=f)>.c&<Y)<
f6+b0QNUZL+,b<-KL0BbKS>a8Gc@;E_PAEPI73eO6gE1fd<,RME^G)SB2PS)6b77
.b9YS0^W@++dcPg6Z;A/fdC(.=QO1(<T7H(G]KF7,L]M?R<:#3[<A-DUd-.a[M.+
X6KUQA7KBB_/L+/<PY^/_6#I-R\+&)_F>F;1W8-A9Pcg4F>;NebM&9YT-9^+1MJP
cc)QJ:/ZOKF+MLX=e;T,a[dcb7=d()_:f&6d\^b<?g\420E&HOX4e.G_eU#PG\gK
&-OL85-aQUV9bG.6^;6C@gIb3.ZC_34:\SFeW_Ne&@_EGE=@[5J3JI+R?G8N]_Nc
O>fPB:ddQD(T@-6FLTeITfXKKA.@@Q?;K[7-GHf5U.09Ib,E1Y]<_QMI=X(XbG18
[KWZHB\><(ZEf.48L<;&@Hbc2H;;8XbTQ5Q5Ae6S4?eG;X-,<TBUc8ZS0=g_T[]C
G]PV32WgA)(NP[,3\^(X8<&S=f60\E-,/V\O7XY@=d#0D;eL204(]e;]C47-6OMe
9O>.G>&74R\PYbEES;PD;Yc<VL0PV)FHT1GZ(1Bg-UHS2OUgfVY+@)TVXTBXW6B?
3(>QNd#,PK8\GT)VfOXPPU_U/Q&:CB&\6\W5a(5<g:VX2cY:24-/4/X9C;5UY8-/
0Z.==OK:87)_9>:H2WB9d8g_[W1R,HF3N<2W2,JBYGH7a\c-eL]4N6FAB^BEMP-H
VD(GbI_#Sd[E8.8BcRQ5BI9:>e(QCM164VHPd@Q\W<#bYSRDOX#X4Df6_87^.#GG
4g>Y,f2KbHJ\#3dI.(^1/6[V<)BK;BaYa^L?+5RR3&gcW0F\)c/K[9O9^4SNG)e=
YFIW;,RE;YP(0Kd5b-?8SW<b_1/#g58:=>Q]I(VFS9.GB7S7gUaE0?1KD]RG^_?I
-L&NX1^73^T.GX<V)^_aL/PcDNBZ3Y2+XK6?HNWN18]+AOSADG8Z?E7(<9TMGCa)
.WYd9DJ]YAXA8]D1Z/1]LR5F6EJ1:7]3XFTTZJ-LBDD\G[KfG)g.gWE^O<eYTf\#
If/MOeG,__fV8,0H@SPS9SEYW33N5GTXGg[)1LbQFT:F,b^a;3MdNQfO]Q(3-VSP
F55ZWaA)OLe+&+c7\+P2f.D;/@1EO>TZTX4=&[/SE9AZCH=46)P6(NPZFg;bec_Z
K06>Q@\Te4-T4cXcVfMgC7RK=/T#EX@&KNRaWS7M7MZV\[\4E/]/SgM)4MZeZ;VO
ON-BK\(\=HYFTYH\I,42H[5-UCaBD[d<]5Gg?UgI\4W@^:aR.#BaI28]XI<0__:b
S:R)e:2-))M:]CW\S[EdDT:LYGL^Cf@bJ9TXK?IJaN>9[\M4746)M)C_\dK@C-bD
N8^-FE]J81)c/Z6Q:9&55)0>7(&gQ</&+g?52[O+6I<gBacXHY6AHB<\D4KP.5G2
KbM0GPddO>E:3HD#\daN-;EDO<_\#e[?;FVU2?&:LS&R)O6eHJQbT5/5f^Ve;b3A
Q#R<:CR14+Te^5](<d,6/?Q&c].@4\6^C>X@76F?DT5(L7-[b\BA-NS2E+c3S3)<
L2F#97_S&W:6D/1^=ZMIUb6B.MF8L2D62CeL(?gZ>U60\,;R>Y:(_M<R+([49<-W
).SC)XM#S1Z4<FA+I=8BC/H68+FbRIWED;\NVJD&W[=:,]eJd2K&Z][PO=LEV#\6
+,=bU^/1XJPIP@U^CGG6RX6M2CYRaZ^=]2J)^:58Gf=Sc(\fgPa_>Lf?UKCJbU[B
J^P[19dfHf4Yb&2B[FBB=7SCfNLP)]PbV+E4A&;eT;>3L:g=QH2V<Lf1_N_fJS\T
F3g49I3gYUO.-cdRJ=Qe01Ib<Q5bfI@^3CP-AF/3A_fDR)U&4fW?10NBO\]&3/Hf
XU=(]]VXV.,7\S:YVUA9KB?.?6,XP4cA)(bgeIOb670L<CXYTD#[A8MGUFT/6HI.
7cGe2dORK[.gd3.LBEKDJU)32_@V0d/40_L3P8f:R(gM_9I-F1.G#,F73-W>6g&C
LF2S8L5Y<)Je@O&3G5)[-J-]bY0eW=1FGUSF7b/]#][_bNDX2,;U+(QK9c4=cgEM
GH5<=:Xe:Hd-7=GFc+E,I/fS9:/NLANLM&L]6Y3d>>6g?e5>aPD9CG),UG5RgOGg
H\2Q?/6\]<L,X9WQa?N7BPD6OL5ZR=8RY6dCbZD@GNf?K=_+RW0cU3NZ<)P+L@(J
EKS0+f1CP1,KVLFBP440aMX]gJLGSG,C+=d\UcF=3<Cb,_Zg?Z/bBMDB]b]AGCKZ
Ad?1)2d@QgO>V_gR]PfNK\aJ?,]f^6B[7]Q]1.S@GMT)0:?GSRU<K9],G#&)beRe
Yg#IE=4589;QE];#d2OX[3LP1;dEZ6I1G,b::-T@61ZQFLJA,IR&965L#VPgUG8e
Q_U/d\V[U^^L3XQE+.V(7V@edAf#(GG8HGN&@;25WWOGK0DM4dYc-88JCgFgP7Ud
@V:=,(Jc?9?TMgTgXN8(XMP=/FNJL(C=,V;TY^TI=>4E5T3B=aU,?-DE5e5#K[DV
0^bI)G#DI_>eA=@T]NDfJK^OUIT2aVZH7]]g=HL+8N8)LV-6.0(1R]4N=bORe5NB
D-J8+U.-.X6Pd/==f#2FG/40>?^D.IS03f-P^^(A(]eW@ZE?:.DT?DX#Dg<e=R;D
YefPDc5Cg[7.9FfLQQ10>ADF+:JT9MHRO)SKLABKHJPCZ>FM1\9LF&X4><\KLFKL
DS77#LTO]&c-LGHPR;Cb;L@1?6.@d]Je7VN@=VVZ><2Q>OWKB]C?3I_C5?/W)9I(
U?OSCZ6Q_8,]PTI97MH;]4&?EH6NZEXAP.A-GSe,HI4_\^BO^g,FP94APfe[I(PQ
J5-7fD,02O-+(C3V2UTCM&[IHYDcZ_bA@/FD<&CEE)VR0TG^@W;P[NcB<32I@XPC
UKDFcZZ[_UW=cF\7XI]RBY+;QHfG]?L)6[[C=4PU2J(AA><aQ\AFP[_LIL7M_7MJ
6_D0c-bT]1F6,<7JN]^Ma&62/)cQLH^&=aSJD,YS0^(+/D15B3_JO,HM#L+HBaD@
@4B;:GbGYOYH-,=G8?NVd5Z4T1a/(bA_^:OUU2S2TU-b[dSDKWb58#2(;fKW.:F6
(<?e^4XLGPXQMQggJKBM<@)aQ8bR4CG9G?8OMHWS(A>Uf7)W5@(g)7/YWJ6NO[L?
108)B9W#9?&XFX,-^]d@fg,?&Jd3VT&752U3S9TK^9ZMD9FPXb-Be]]^&>eXBeTE
bbcGZd[cfd,:#dU?H8EVT+5_<=;<d\_SLf]P7HFQP<<d9)4L3^ST[ICO:-#AQ9)2
E_3Q/g)/c>VQM)13DDQe2CZBd1ZQ&PN\4(c2+(_,&+(OF]XH7H6)edV6WO.c-#X<
+048)WS02;K[PL-YO+JEHFa,]+EdcgeKGQBAJGD2X[NF^_J[1R5YI3JB(<0P2EVA
A6^^dc\<L.KBK/Kbf>Q\J-_&G.L69e+_W[d)Q]DPT\71Z.NANgP-C[^BD#L#88eF
M1d9JY/)=)U7KFI?@74M&(\YY#NA-e:D\V#-@F-XA4[12b#1QRZZU5Pa,.b2X8/2
QdaD:?>3P_9fC_>4Bd&E<R8R4-QHHYVXJf>DFF_eN2DJS)+W-)&_]3CIZYTaWcdL
^M.F0Y7,J30-;-^,ZCS7?UWN[U,(XISd:J+VO9Q4/_[]7]aFJSD)WfJES1TU_8:L
&>@S1S.FE104M@@^G];SW<G=bZ,b:@7&dK-,W7AH(&D\=dd8Qed0(9=Z6/R.M#9H
[.OC;<#[O\XHJ&[;9]QHO;J9@_cA4ZK#\5#GG<KJQU)dBZ@TW(=[4/a8)5-A4K/;
&:-NCD\^;J&KHB8R?44^E@+>_OAf\08VP1V0(@ZEKa9=Kf1<0JP.d)Ab3PYFWVfS
S<bJW3ZZ[31_R./PN[(XR-B-ZdcL<U1#.Pg1?ES+g3,]/a1MSf2PI6=/^O0K(+R?
RGg-\NL9Q<?^=4Y:C;U7O[6R)O+<S]eC\59<I9_9SP9.9Y(?1C<>3?,:,<;SUORQ
F7ID5a&b&;38Q/6^?R]SZM=BEQ[^=#N(BW\Y/F2>+4TcU(=F=>S3C27^IM1;DR#I
.N3_7&IH1./(RQ8aK-AF@\11)F7W]cZ@\d?.:AM^Q&&KdKgJDaMB]7O1MFAPEA(F
+QU,NWdZ0<Le=U<BV4N1=#eW6W.FJ4#>fWN7E&4^D8S5^[TP/-M70]X[eZ8_F4c1
4SD>1XU\&ZDS\C<C,V(d371/#_-@eYQ);+/,[>b#^[E#@VJH(d(FXV?_3]BcIga+
PbK:19-e5<[&PGK@,H^;O)3-?\4L-:>&5<4&B&gC3Re[L+=[XK@R8EcUb2WM#fJ<
,3S9#?>F9=8ePRG<2^:[gd9#8VX1QA-,(08Ue2>JJe+<CVR9US?g9a,:_4&^,]F&
?6DVP?IY<MBJ=c)^#ea[Q(c0b@=a(_>ZR(1XUa]Vb>7@@>ZT/\=+[2,V-_J_c2P)
fLF1&;JVM,4G5FB8D#R54K\a;J<5+,8DHKaE,Q][g8bX?O9e\XaU8B>(^HM96[.V
eWD6f-WNMJXc@PZ2S_/Q^A0@WVTFK:U1<F.-#GP_E-C?0K1U76.7N;a;G2>U<RAX
-f+MLIW5_D:a:IW#EaUeQ6SQ.dG9BD\/CX=2SQ5@F(+4@g5g?3L/ZGIB9?[7&5eJ
0,AZSK.@QaT&Ib/;&5MMNO_8;K&=OK\JE90XU5R)#^>_gYE[)#5UK:cGd[V=bGGV
EPPM<f^-&:S[@@a<W@VYNX\M8U.)YR\_PaUa/I+4GYX1B8C+KP@I=(8+:@5:2=QK
_7@],=e0+e^KP3YRHV_NL@;+^OcbB[LUc,IAcCG6+M#+0R\/Va@BF&)RZ.QH@0<U
b?=3(ND1e48?23^0&2HAbLET-L43A<JL]B0J-fH;A^;0SZMc4#:I]_<fI12>(A9X
@8NK,A#=e]8eAdB=EV5BYT6<aXYHZY0<FAU;)+a5/^3-8B,<B6S6FPR5DBZD7E3K
NYMfO/\FI7:^&8W>GY;;_Q=GIHPHP:5RdK;442e&>]P8FGP:AI/X?MEA+>=fe5Se
XM[=5a.R\^;=QJARZ(cLRAHZ^AfDfXTI&RJ^NPGJ9.^J]a4gQ;+@@Y?L.)b_<_b-
N-2W>QCE\L:bR//8Q\QYY)g.PV=gV]JGV./FBaY2KA_@a2S\1Y8AeNK?[I_Ge]>O
W4+FK9M4G5ce8LL]9#]N/dHRdS<1ZQKGWZ//V^Bd>-L4@bKAM>>5]Ug&A2]+TRX[
gc)=ZMTd,@776Z(Ue=3Q<bC7[F2LFN7>:Ja75KfE=@WKcI-2A\+5Na;PRL/9U(^S
Y9-4>3Z=9G99K9ee#6Q\#X_O1e]NRP7K\6,5[+@\8Le?-MgYX.D0/3dRMSWD9VOU
;0<F/IZA^0W1](S#2,9,2Q5>DB\&5fV-RVbMXFZPXT-\gU14FaJ>ZY=e[PCT-&(C
DIeZH,e.C>PI0-F4dd5W&LW<N<Q)WL\;ENg=2Q0BOddMPSee&T:>IQPgZ/TfeGDL
0\(c<5#YOTAR=M>c_dUHaVN5:T(c]FV<IZ9(K,/A0-af;Y\KgabWE)5&W_2RK0Bb
+][611S:]cb&H5?1X?]SB)=H)]Q<4>9/5/FX48(dOQEQEaf::);W+RJ@?VI@3<K6
.?8DWHB)&e8_CASgBJ[3\R;9LE<RJ@b23,WKdGY([KCV-#DJ_FE419BDaBZbfH,G
CMM&H9Z36ebOMD-9MHDb2:=LU3d5L^GA>:Z^HDCd/@T8F[S(a?Q8<92<0T_+e_T0
KH,QYfeT+gdf]S/R9U_Y#Pf#TZ7&45YfD4^.UO:JNP0b:2R:.bP0Ac0&?AB&.@8P
KC,YaZ=3I]IH+B6=EVK;SeN?NWENXdJDb].5<:W?N]IgU/J24#6^7E0Cb6;4RLJD
B8-fe)LXN5^e/e+;a&f<FXI6,5bH?f8Jc:+ODJ:]6JC_P:@e+]<IPEYSK9?[ZABK
G/Z;-#2E@UR-MO\9YG<OS2@5b\bCZ6V57_eC#V)We0-dFG@G81PEgJ]>fZM7]a>/
g=<J>Bb,OA4MHA\W:4,(N9K/1KaP1^,_E]NA&(ace3U#VKT#YE9ca#b4BMO0e2cV
^ggEW<ZX(U^+>&MNe^Kf2DK?fF>gU2Ce(a6#?>d,AO8&UV#a<]6V><<C9(3_,,V3
dN+,N&O^^=[;Y+LTeGXWP<D2d+SMa6cRH&3Q/G?SLJ.fC^T>2=KON2(Lg/)[5S&C
eMHK]E(7C4Be/D>.X]<T14)_4[_<fM\)a0+dRXEZa0F<HKF)3^YAK)be]1DgPUY=
W\f(Nb)8c-MV7EdBKVPF_-aaCcb05TC-U:gZD:[-Z5=dc+]2cWTfYARX<\8@I@ZR
Z=G4IME3>0F:?\&[1DQ2^Gc40\X<C.]2SW8<?5L0XGQOe+O.Ke3)S=@N.<(?U+^:
5@5X=8b_STeOaXG#\2LTM]J_c_[?P:4R>I<E^Y7Fa<OgY0W(O?TRD&>?bF.5fA=4
#Fc89([((.YfD&LEE++@\)MRXcK8@5>43Y<:Va<XZR/-C?+A1:S/1]0[gDLbV<N(
1ae_cO68]K13FICRF\@\?(T&?))8+_X,c</9LDK;>8KYB=fARQfU=a^F\#)HeM/S
[)5_KLAV@26-PNfJbe@YSB>46V4GdO#@#AQVc^V#K4YY[3bU8>#TGD]B4;<IULY3
=27LCa)40<A+@V[NSZ2G0ZT)VBZB3K_(+^I8,UNb^DdK_@^0S2[H6?RUJR-fb>2.
dgRaB4>cTL]7+A^_f4LIOH-#^64b=0G&P8GaUgE)5HDLDcCW(856)IIK;IWU,J7(
8c6ZgZ0#+([d,Y?JfAY/RD_F)J\FUWcFLDRU?ZRF?TCA?Q+GYHR>L>f/AP-PU:76
f^0_&b-/fD87C^N;A6bY#<(/3cZSEN6KIZc/W:\4_&^FG+cBMgdbQ7O&4MQH#XOT
-LTS?fJe-X_10+<U)5A_BB]MST,+D4C]@O6U4^F=cP7Q.5OX#],&#G.VYUF.QMY.
4]&WgV8H2AKNc83Tf+=<>_)D7\L4;6DTg]\#_7^-]bPJXK9f;3A4Hg+;+f&ROEGc
:]e@.O1Q3[[C,Y:4eL5<MGKBeOHD^3GM2=ZP1.\B?5K35C:W>6L2[(XWV04E1A+_
]Se3?8]eEWZ0]T0d&EKF2_TMT2bcb<#cY7YGaX@9E1-J8AO?;@CNCO3G7c:S)OK9
D25^9V<[E_31Fg8\<W#ND#&KPJ]7;I=)DS,f=Rd.dc(TUQ<2R7WJ\\1a:[182Wc-
d#?T_&cVGE0&J01@aA8EMY>Qd@W+eZ_Fg\ERb(ER&PL=P_+g,S&:=K+dYSBXQMSg
U(>VYf&b55M@W<..?Rg;a6SK@\)TQV[]MFY781?10RB6+b5#5P80)3\JV)-edLDD
37@L3Qg^@YR;;G,A@UBEO<10ZD]bAg-Sb[]AE]BNO0Q]K0DS^?6,&Gf3PJaf&&2A
SL_BK#TKD;NVDOH=0PVbA\YFb,/T\gb:H5TP^0G[#5F4B-Ia@M?15DX@V#W9>[:E
LE<^ReVfeZXPO)&9_MUd+#)ccUCb2;_=J1FX?FaDW4e7e(AD@YC?]:-QXOCf+g#:
#TQK#M.3<FUGFP)OU48@\V[Z3<@;.aU]1<#SV-J6W43U[4B(6>J&S,XZPUgXR@[Y
7(D-M98\bP&9N;2)H.N/?eYgcMHT0]Ndab?SSDUFA[;VdaD)+&;DeIW07X-&C,1[
IDMDRbHZ,e)d5(/_L0_^A4MJW/e/H#Y9[>;>UcLZ8EZ&EH,Cab6-EAdM9+HA\C5_
K;FAP:DM>9&:@>B9R(JJPN(A-,:E&):[P64W)g+a?SaLdJM+5c-K=/M38:1U]A=.
EZUE:.G+]N=OW?Z&SD(FP=]ZKB2ZFL/<,Q6K5+OeSQ>fd>C7+&(>aMNG1[;aB9XL
-ESF^)=MD?E)PG+KV8]QWW)eQGKQe,Nad(YZ4_R6@:f8cF^.g?\RAQ.NM[aOIT9Q
fSe\OCaO3Ig-W3[7)07aM#,(THEf^]OfHGX]G1fQ&DQfJH&+Ce:F#7JaF#0)c)Cc
S:45Q/+WS=/L<S>KPXP@=fT(Z+G-[NaQ6FFA+GK@FB#1dH[FFV4@CW1(e0N^-b4J
b<H>;-04A1B^J6>;)@0Z8b0202]GWCIOJ,^3P7G?F7aL)O8^abKC)4NGJFT3^Qe0
Z(b3UE3>d&7DN+FU+:Fe<K[dL<V9IXD30fGXCV1\\V6UaZf3DHd1[aWQ52EYZ38X
3UYc7KKVaXT+>/QIT)dB/O?M/K>>:0^[9NNaLd,(80DI:=+D1_(4X)g9KE@HC>7(
,KPB\U3M&);+O:W))65J0Xggdd/a=O@LU9#WgYB3WC^_2YCRc5g4H_]QCO7.V>/X
KTX9)=\;;\g0Wc>c(I]T#ZFR?;LZR_H\&.ADYL@@ZgS9Q3cA.3:#aPK^5X64&4;V
U4I^>DG#=:KUVOS,\G]^75-)JJ2b]b&1POZ&\.VE:4CG_#&>Fb&J6-C^M[cT:1)N
g]8X(KR<.R26IH:\XbYc,WBP9M?66b3X=),KMVJ-+8D4U_8=\&ff;YLeNG_>N0;&
US8Zg3B1Wa&0.=[bP#N\AN+b4819g/;aaZEM9H>Y6b>?T+g\Z4SEKJ01Lg]NJ1S\
SZHAg6HO6WW2K4M73RP&ZAG:&TM>KG+U-+UUeU#NSC^9Ra?gZeAHa6^@STX_Z#a&
f#9PS5X-F^1W1+G+X9A);I-@+IL.eP+dNg)Ya:TQDcc1O>.BA7KH&#\SG37fOJ3<
L.@YZb0(&\;[4\@/?5e;0>J_9#9AET?M\M#L1/I)<:YX1W=BK45ZfI9Gd,8)BE:J
N@XPH+:AJf-6]_.g2/B_#2<>>=I]17H^XJPQK]]Z#W3eO@I<S;^1=gIR=G(SG5YR
<a(3@PR;V(fZ?V4,4bgWHBHL\X:CQ4AKK?Z<:;=PD34Z.=A[N9C#)MEVT_#_E3OJ
bfMeJD9=bI/N)@MW7;6APM:aX_-cGU[HH1,DN@3<f_@/bB?)7EXT@=./d\\K+dG+
8LK?T8#FfF+5?5WZNH&KOQ>b)F6)N-2AP+/9F>+28W4Rb_ADL0M)d^7\MGF69C@c
cF<GN)23Se#=dNa^WOX7XfUP.<0C^-R5Z[90W:K24E7eYgXbJL/gU:ON3Db8LVG]
f(71F.bI>L;JJZ&O>/&&Q^PTE,;U&e8Sf,2KVNSOYR\@G-QVGc:)CZV3]U3B5(UD
A#_e#2ceX;LV5KEHcZTPTa_4]KfU;HH\H\_+E;a,P,;8cFEST:\85VV]K9;PR&[O
K#PZ[QL46A(0OR8_OTK?M&=DR5[-Z^e7A18;08..\S6O9fIZ1a&<NVL5,gMCS-B]
PH0B@H3D7E1K6B4<_3@eMGc^WMKMSWVJ;:UQ5R9-8,6<QLH2?+9eCM);M_TE2Z>J
C;6R2,5=eQ?0X@#.5+K>?);fL<&-#6\E+\^5;TD2SGe+O(+aDc[@]6D1>0aP9b:B
H&2)5gf8dG(])GfF0C58-;L2<^6#7HYFXWCKTP(QI#_2b0M2T^J&abI0]M#&f1Ra
D>bfdGV6bYR1V>C4WB)B1YIG@_FRbB5T]FHW=bGQV4(:HSD7)IJG.C\I.?U:#03;
Zc:N0&a,\L69c7XZdO&41CgMWa>1L#._U#bUBfKHG@9\-W9e1PJ^]M6)cea1L&LU
QfSD:JSYP_2V9#;Eg@C=)Z+HZe#\]B[Sbf[eYKM[K&Va/^O#gOIYeHH>-D1XO(bM
_E\HC-)[I5aRe.[@.?=SEV1)MCV7@M)3d^.f&9^KV/,5gBBc:MPL<VC1_5AMK7L6
/@IN1&C=Q[3OH,DO-IaYZ0IL73Q?QJ+STG9PeD/:Z-7<]Qc/OFbb#;\^EZ;O#(/W
2D/74a-N5<c5[[VH4;PbGV^=e<FC]9-Y<+5K21&c^AQ;C\KGZW9baS^D^3-^4ZB<
DCF(232-f9.P_@7.:c#-S=^?W:<7PL<P[W\cfdP>2)H:?AL2SHSY>[Q0FNF8ZP96
)W/5Fe7F)EgG>IQ3.)[.-.Z[]4\]H?.^P1O[;(6-B.U>Y0_+C(N^b#A9-Z&fVSa+
V5;?Y/CK<db(f.fbJB)aL0WAE;@aZ]F<7Y\O,e\W.+]6]_UK?O@dSY4&,2-TB1S7
EE@3Qe=//WDJPcPB();b]R_6A0bX7\>V71V6g:^&/gEXL:,2c)4:MaB703DC0;dd
Bg4DBC=EV[#0Y-\g52cB8d;_aO56&\[M_#fg^ABZ8=eReOWC61&/2M_4N_E-L+eC
WD>1_WWg/(O_>a;&G-/2;XIPgQRT5B>I)U8]-8H58)?^.dHe)3V2MH9g\F#g/XPN
BX2I<]W:@7g0U]aQT8RZ@e])d+;E92(9-c>V@GZ)@TGVF#/1SPHb)<H5FYEMMBeg
d..YWGa5UT^[I+POW,#YN3&^T1aBd?(-0]TL;+?feVO@&VK-aE@7fVBT@^)&CXg[
^W+0^UeLLVQ3?AdcfDVfd]XRYU??+[JPdfbP]LE:),(KYEdFg1O08a1?SP593[Sb
NC1OeUQP9(JL9]U]=F;J67[B>_L27&LE6T+5=G(5W_FJVYa+dacK.eY;^g3CP<D[
]ZT+eIVFE_XWc41GL6#V_C_(3&O#E5]&L_YPX-KKA(N=.)=?S2=.:C43d(6#8UYd
V),YK+cPa8Y/;716O0>Bg.YY\SY-If-SX47OEK&aNK,Y4MLH<;H8FGf586?1)RAD
\)0T[/f#Y\@OeWdC:<>,H9/J)=:#ZGdXTQKH=XXU-UH;W<Z0=XLLJLR[K1UM/M<C
;B=YX1,@DF:EN(9?gU-8:ddU_D@9T^e?bK)I:BX&)F3ICfA@XR\eST@JEI@?U+T>
a&e8;/e[eZ;0A>+EDK)1KWaR=,,-.6G/S_dbY_/.;Y;)g-INa,DYR)LbW2&0FL)Y
OQE>QaG=&7P:(@[7#O^>?.5,(MYH2949HdJT.K#[GB=,U^6Ff,XO(C/JOUXP3GT9
9^Q[DE?RF4_-:1d+:ZAg-?^3cPPC&CMXC8ZN9DL(5/TEa:N(gPOQ#NJKT2=c4.fS
(KRDU7aTYU6@DRSEg@(1JMM9CABOMW.Z9#^\U2b5c+/#E?2+N.<SbMf(7(gX>T16
X-0.5fG);,566AS,e>#Bd^P3=W_<_L[V2gIX6QS5MW+=QVSU\&#Xb>-4,ORMQFAT
eW#-,JR5Q5<fbX8:16eK]\d-BLM>OVJ+@V/cg\L5V^I2/XEEYI43FL7=/PJ2@-QT
)3T<gJKBWN)L08.3&V/JTS5G)eL/#Y:?QECB04CHEDV[=]P:4P\:O:AGg=@-Y,cJ
O_1F/2U]VE9FdeC)P@EOT,TTU98eS55d?2A,2#E(CJ6],LO/V=(RK.O^.XKEOU78
7Z3IO+&L+\15A(7FT-.@8V5T7-[;?@4>UW?(Q3W0E/;=Z0aDRT]K?XNP]JZV@FbV
VDdffKVB3fLZCPZ3G2,;;]=&[4-3dM4+]WbK)7)-68W46Q3\d\#F3^AY0JQXdO?_
6F?/6C[6<d+I#H62^9aMVR;U4ZY1(4G\U1X\a)AJMER;RJ.aCW5Xg\NNeC))[e4M
(LP]<I3?)\D1HD?MR5?dIZ7I@MEV1&#;([.4+Ee@X<-e>E8cFLN&62M^Z(aWK4eY
:NT&#^f-EDYA=-[,>f-G&/S8UR,K.)3e\WZS29VN4\b(OUeC7bOLJS)Q@,3R9RP=
eFGEZ3[2F2>@Eg&@9ae[6d>K7EOL@Y@eff^SI@ES[^_d7RAb^<V0BN671WYYJU/P
<&46U@6d,HOZZX7RG:Y[_5#U92[:5HK.W>^V6&W[>fM/=YVc5+?FL@KS1a-Ce\a8
[_Yd5<ZCV9++fG>K9)+IWe]UE<3CUS2d0<X:)ggW(93Q_c+eLg+LTd-<MHS_ZPL/
A\IVQVBA@UZ3&UF2g=O9bOc:)9-IGH2A=Rb^)H63:@-8(]Za+)SM@ZGbNT2ad\0W
H_XbNc\N?<P>5TH\[S#CHHXB(EFY-cfedFE,L0B<X_#&BNBM3;[3E4&Wa@9@/N0H
BSLZfg<_D9CXf+:_-?7NPO.==-YCLR&^UWX\:fg)\T7ed08WcG=W3S@-C,)f=Q&H
\.CK8IG7Ha>GGWN?L[T>.5+NDPfZV2C)0PNE8NK<JP<TH7f1WS(&c]CG8U;D44dY
W:JI/b09F^X29Nc-^]e:I11Y-4X)V<+g?,&Y=43Q1@-1g=_9:R@A8T7;-Z0aASbd
3aCZdCHQ@?:V3V.?8?+Hc0.bP5f[^c>DE1bBfMU;Qf1,,fCET+XS2J?ZY[?:+ZBU
O-_6<W+JgRW[8S,RHI45[X,Jg=F1KJ1<b)W0,Q-.5+-IHF],OC,[bZ34Rc@e[K1J
;O9bV7SOFgdf(.PFIG@/.K--SS3?O5]F:;E//#:5Z9<R\S.>&4R^dTOIED(#^U0E
dQDQ+2a]]CHGP,3U8e0>)=CPVbee40=D,5cL(_[XU2WG4@]eLZT:LC^\XPcHTF;M
:C9Vd3CP)=H78S?,)Xg-Xg9;ab3bZYSAc&fdR7FX/f>a?57)-@SPCSDe^V\0\@Oa
45Tc2da9DfBfTCe>67(0D;9[cB&dPdF@4L_@#aI.W+AM,2b^aU7/@fL,E=8I+bP+
_BFB@:F<N7M+ZFF/8)B-J1.//f>WK.&e)adWO<_cX7YV+W/BTGeQbG6c7c:,ZN6=
e5[O-Nd8fS6G[)RG72<AHBOQI\#M<\9bQbEQRF4ZXFU.A]M__B4/U6SWJ\DHTMCJ
?a?:#@(+,eTC16]bER\MKPX:28:>&KQ<4FH\(;(^)>R1H)b-.CDD#^G\BX@M<Sg1
\JfgQ_G2H>),EeD_a6HEG+/5f?7WQTZ@RSd7X5+VD+Laa6H_fO>3#+DV\PQ58S=0
L)gFR?)EI?Y,=S<He1DA2?/R7\]-I=@;\4PL7,#E3/8;E5eGa@9=W;7)&a15ZZ<U
d1@>gdW(K^EA,_Q6>V#Z2_-Y[4fB.VT6=2Y3A<eWQC#Q<;b&X<&551eP^Z\IM?]_
K2f@WV9U/AYW?<A5<RYOWAaQ]60=P34O)S;_JQ:JG=<M5W\^5(@=g-I]0,^gCa_X
ed>2^@+0]N]48UCHY+fc1dERbKCO+</65)9^THROOS^777HQ@S;B;BU9QB[f8=41
J.=aH.+/34BU64.796IS.:G:BMVdZH03VZ4Y2KeH3d<IO#JVJeDN1J6/.D;@eECN
UE3bYbcJXJ(#dA;6#\a+[B1H<26WbX5\SJBBG44KGJQN-fP.EAd&/#;,LLB;DH4.
Of=8;R:<7W]TY4QbEA)K09#=7bA:<Nb,ga5eJ=[?GPMF>Q@&JT&DH^J4:TM5>T>H
H7KRDbb<g1AH1LN&AK[8d76#WOLBF_)2@KK+/5-BO)L2)))Qf2,R,GAb875>Ja4c
6WMDa_=L;H_0II[=M_8/Y>QMH=L;X=XW8Gb1?,LYc<I<X8Za4D7W0fT:(79Gb<.U
?R5YO3C:>gBTQXZeA?V\_bMda.ZN;9K5^(^[Qe=cJD^/d(&ZP<Z,:6fBEaCfMG6\
]LY3eC63NU=3[>faG@[PD4P#CUCMgL-9LM>ffEVA53HQTK@(RBO-T]4?e:2&Of-;
]G.92#L#T9gX:#UP8K[3#_Y^\&&LB:NU9P4_QJL,RLL^1UZ37LWHCC797\.J:HE\
0HXCCK>F^:+8^2dS8;1aMg&DIJUAFFEK,>L.D0DXJK7,/21<B+KfcXcQ?++=O8JD
&JGVERKe1P930-dY64Ef)D[cWG]M_dEbS1J0@@W/2P=R^5@e8]#9a5]fg;8DADf8
,;CWc1:&da81].9QM#;&)N8792&7CAJdZZ=<GbM08YZVE:(NGcQU2WI9B9d&?K>9
I>/01S<fCO<T8+-/RV419\bYcU0@Q_?LO?HK3@fC0N+N,C5CDFdb4-0JOeVWKa7L
VN400&TPNORfIM+JW[79aHSeZ;T)I#+S?aPc2[QE2d/ZMTB(Lb-P7WaKCb[Lb7@C
Q2HP#8dJB??4+DFY2+aYPe\<SUL8EQP[O,@BOBDIdKSYQ3T61F\-]dQ^3(g4@)P;
1aFfJ#ac2aYQ:\?WfX-0,68Q-J\KJ-3?M#Qe7&TK4#^+W7.5>)PaT;0649^QTPD+
2B1;.Kd9_5[V5d900/\ZB?D-P5-#/OT3W^a6M76:BDQD#C(gF9H0QP2IN^R.;/^\
H7WXf+:1AZFWJ9XL2XON@b1+L_@]E9?;LN<S2\&KL]SPA-,E0<)G@(#<5OZ(-+d<
>)?S#BB4Dd+/dID\KI<SgI9fCO1-=\^L0_]I.511_DEf.8PO].E[Qe-H?7Y^M7P:
XP7#fYHSE84.;QPLBQWDUJW95VO3]CFFI<9#Df4@P29A5:8U-24G_H;(aYA+Y@FP
G<FK]=;WX<[>5e+2KY>\gEGI6TW_RPPCR5\<Q?X;;R<YS,88_)?F;0gcg<R#&KT2
68&f5,^8T[<N<UcT+cU:C&S0Uc-/;1]F;@5AY6C8FM,4aLZQ@NZI:R-G2^[N1WR+
#,@>AH51OP7^>&7-;S)-C9VBJaNJd#2<+@F^(@T\7a<?-<)&2LaRV49@Y_/?G#bQ
:W?gaHd\G\5^F]aLW?U+KQUJS=5.)^;fKGgfF]KDA),)ML).HQ;[CKc><,O1]<G0
c]2?]KN?@b]Md+2@Va7K7T]J_e_Ue2;9VEd.AJ23G0:gT5#ND86OX)S5]\J.1Ebd
(B9DBGGa9U\8IX&8a3TXB+>?]O#^LBD6R,OA[S976cB[a/V_F8/N61><DX]2bW3(
H2,6K?8K,_?95594[;eOa40^^,?[L(_XQ0X#S&>=aAQ8^>;dC\1Aa^bIK@=:^][,
CAKM4XI0d;fMDeD+KIK.FO#<\==9>fNE6W4M?4&;=AOGFF=dU0,Q/g&9RCFJ7Q<Z
F;H;8@&@2.a0SPc)fCN<U.+\#[0WgS/&LX_P?g)-@N=H171Gf^.\):[4\8aV#<?U
P_E]7(F]KF91EJ:/6M?17QfSdD8,JWfZ1DX=2ScWAFQ;JDDa2+9#GS-Sf&:&#?c)
;20g0WF_MWA\4QE\-CWPb;8K\3+>2(CYWLQ8H4E;(DD4O;4+FZJ0RMc;^K5#=ae.
_XL,Bd-<X^TV88E4.;>0,#P=/?J(8ZY<YcM76#KfbN7Xb=egFd;T:<)>8I;B_W<F
(,B6<<;4DU/8deT(;ABf:ZFYL,Q(4WRA.79C3^-J^AUPR3VdDO?<(<F4eB9/P]?a
:&E4)>_?eg6OQ0f&?8WdeV5^AOC[D2_3XX-V5F]X),cFP1KDLgWcc=D0IM3HM#(;
GOZ7e:JGD3\dZP[EPg(]HE\F>5:FMP&&D&Z0bV9\VcZYL>gfJdaH_5#Y#TZ<S_8I
fIJ4@abbAb:Pf/]LP@cAV<>4.^R05NBcbf1I5XZMWCKUB0UKBaY5^=:MaZKD+ff_
>3Z#>fY]DQ)<>0RN9JT[S<(7#G,Y6g-3JX0CJIK2\PEM-^:\A^c@=85IN-/,7aL0
>Kde0EedEEICA/DKY,5\gVTE)6@MVF3JU-O8_(b?cQNK[(\^ZBDE:gL0B1RPB3Pd
>2/;0)@=<-?Bd9Qdaa]6+T)1CZb.Y.^<HBPLe[?.>PADGD(;Q&C^0OX2\?5KEObS
Z=3b4PL-6Uda<eC_08c\+_ZILeY)B&H77.((^^<c8D@?/a8:KQ>,I1/&OZ=U@U3H
HdNHWAZcD3VP(LGGEL]6J8(,g#B:0N_M7]_Z60OU-1+(.K)=D;a^U)#]b<X+/4DX
3SK&,S+(EC^2H4.8))JYE5eR=AAA0M#WK?IQX;?Z2(8K99@RJ3a>TM7/N0EG?S9g
1N#)>K\356@2b=H-):@gC66SQ.#I6_\0,4C.XNU+IGcA_2BW3G>F7Y6A#H:G&U>d
[ULLBO?ZO)NF[XbUL:KMVHUY;Y8B2;SU@8/X7].e(CX;XS:^0F,/LWXZ6<e>RL1O
VGF1F_>CP/eO91T6T8Rb65:.(?NaFNe@4((#YY[.8CV<f)fR5d>[@[S4DZCNI,=Y
USO#/>eTRd^;,47NHa@J4GO]:DIP8-NLWfY?^E/NfQ&M38;,=G7EJO5.PPf.P]T1
E_=eUT4Z@Zc+YQB0e8:33L8-K^4U(V&.1NOF<e0,/M9)4OYZJ1GOL8dW+X_8,T8L
)-F?]5De)EM&3(H:U<gPa#\M/E,N<RfK=G9ZY7T;L:XeH<(7(eXd[2XfcI9/KbO/
_E\Z0NA&JE+AcTDA1F,VeaT,fb[8?E7AEAI5dN.Z\+(7OVG>VDZ6\Pb;Q/2G+G:H
0J7)6]Y;R<E#N._XW;/BW+,[?FIF35YX3:fXMJ0-,3a3I#-Y4WT#;O&&T^AS7:^0
7YK]2F)MCF(WO4@XCU3DGN-FAEET4gR.SE:XUZ7V9<3P#)=baZ)_X620&@5HfXgR
Zdg)4?(9>@C>?8B>F[3CCOXH>-0168>M.)a&PZ)&O3c8C7YJg=8R0cFe]N9_B+WT
S8,G48MB(O1@,-<Y5DXdM>1V)5W@2OC(S>F:/UeEc=9af[c3)WTa1AS]6):D>VA)
A63Pc1=O\^((J0B29cA52B=]IO>&a4)E0D+M/b[E77BVZ9RM7)65b/(>YHB@VX\:
1V-?X_Rb<<DOC(J;f(;PcC&gEC4(T/7X42)G<P.?,ed?ScXS(1KD@])03#[.PZId
>>>gM1>/&2A<AfJc<8LM)Xd31a=WQB@Y;+2D1^[+<R[FQYdIX.-+WXSXJ@H,VO;a
URE[OgJ]d\R2EO)0F/03e0#Y7a&G-,RY068Md\J/Z]QO=]L=,4_>V;#T-V67@XOA
Y@5B&,BJg8ERZO#J480eaK>3]^GQ[_(;YP_.Bb(A5L0QC&1da<9(8Y39B5PP+E:[
@J+OKWAFPVI<BO3U7BLcYaY[3MER+QPJb#8g4L(S0[]-TfAT)>9WdfV?S+eLG[=]
:UYX5ZL2,X9:Jc9-d]Z/c9#<C0@Ha0;A^[bQFUaG6L5YH0=X=&@0EU.Wb(JE29<A
7T,8Vb17T#fQ+U<V)cY3?[fd6T8?885H)E0fZE+-.-]gZU+6aP4W#2X:A]ZW2>)#
Y.LQH;_&,-:I<^/;BV-Od==;8=S)ETJL=7IOeU2X:f2VeI).P:Z<EW/RJMQQSX#T
315,BZC1\F(.KK[<dM)4OBNfPU)/ZWT+eXX)\FCg]#gTL?SK.b)MO]H1G=aHL2gf
DQa0H,8Ef<(R:ED9]U>7K5NaBLYE@DBRNJ13GKK&C;),bEg+Z70[2,3gS8\N#SAJ
ERC&VP<e21?Q<c++/01&8fWU_B9VWMb4_V5#Ze&A8=/SO\.WAF;,RSGTg5]X/b\W
]ZfY9UDBb_W^SgFU^FJ&-K5+FQ;Ff,N9.g=[0[;:db/6/33__L1#J&#b)^1TASUY
?#>a<9@Q70]7\BF)X1E)-gCdJ)H_Q;:N7Kd)fO>OZ2?#2Q@+=,/IW,@O]/Fad&=c
6\J<37aAE^Jb.\TC2A<]DVgD>2\\8/]PL?,1+/Rc<^/_W#P=8RNN@+6_\87#7IKR
5d]K^E#GF72H5ZR[g;5+d[DVJ\SeB<K0agV@(M._0KaLQea]&[NM>]BC9;@,(]-<
PJ;=N.7+dfGBIGdE8CQPH-R@(3eS)U1GJ6PZ]H^S)V3HM[I:Xaa7LFSUSA4]9^P;
8FgCdM/=F;3@A[]cd2e(MS-c>[Zg0N^^V:[gBd8)S2cf+<-e,OHSUV=(DYAW1XdK
;FS/K=JBAa]-(NdNeb31,P93L9W_UV\PE(169=?5NYQJa:DG=7UO,),S\aPKC:.T
:,2W^\>9QLA\J2494\VWE8GRd4UB&@E=@R?]^(,X6AIgI.SNLG@ddg,W@W,/7)MK
4QQX9[^M&Tf8HcK.L#\\1).Ff1:&BFRABI\4NdWEG&cM2YEV,1UIWgGEAJ/\MJBU
LH)PDIOcbW2]ZE0TbUUR?^IA:_eLYZY]9B13(N\HE:87cRCRfU?>4dPEV@P)LEIC
;[7<X?6CdSef\BMT?&&P,US]>dL9MM.WfVV)E[YA/dC2)X[NC,,aOOOAf5HFG_Te
TCW;_NFIeH-B2M2KO,8]-CMEMbW\&(#D6I0Z32@?6_Y+L6&CK;DgCYIa,L,1]GE=
&EeXDSGg:7.I77:L5-M&S?,AFB@)PcW0gT[[9MDQ31Y[ASLBM+E,_1O2,J;2-OVL
X@0JVUJW5<K+C(/3gK#SFO]#<\E)TgU+,:H--eV/WV2G1\3P_4NeU7PDgNJL2>B6
_F(>@<U30Ha1g,S1+]7aI-;d^<I@:XF>J4[R@+7bTZ@Yc3A(^18eUJg(>^0XGa=6
=d/JR9AF9>(F76NKI46(2X>B;9XTXI)(8W0:.N>[8A]c^QP_gdZOA&MNGE,IPY@.
)@V;SPEZ20S/A4E/DgID&(+/0\M6/_b_K-N#gKW[_:DY<X&d/[6N/JbO[TMRLKOF
#)XD?:,:QbPJAX77d6JZ<Y>Ka(:>4g\e)54+]c.3DRXX<]CXeXL,R-3NBSWW98V-
K#<XC0egdP?g.JZ;>FB(b=eBR#@HC(RB-V(RPH;XZ0<F;aWK-H9>;&CK>-5V1_XA
(F2/RN3-<bg.N/RVG(I?0^#g-TSM8[VEX1f-2&f=#P,7MEV5cZ@>UaGGCQ9c+5(<
5)8TWCY>;LQDQ<fT4NB\Z6LEL<&FT#7J/[b2VNN5cgUPb#YVIMG=:YT(+OX]MTKO
=5N]8^_FOGRdT69E6:1Lc9_,9XJD/21<I63D2P54V0CA3510.cY_Z=8RX+R^)?d\
Q>-1/J;DV@)MKPf;L(9,gdN3ROXa@T(#@/[P8673bfC<:,d\eW+B_LT60BAYRXNV
/WF;>B1&)Nfcb\+bG1U<LbUK8<.&P10eRR6U:^@8?7;W6G_1;C,>WG>\8_ZHW#KZ
E(V:WW4<BOcQAS48,Sb[W)K(da>AX1WeQ(&4A_Dc,-8E-JKcO9;5UdT[;EQ.DEca
3cZ&d9-&9O>YW#H0<d9OLQNbP.HW9WOW0_F30C68N,,TM:ET>T_/)[<N5WGXP;\5
SbIXd?^K<GTJ4>SU<X/b;,a)_Q2L^KPRFC@N7AJFeQZL#(>X>COcC[34/DFZ@<\I
RPLA5JV=1G@dNIM,6J&X\;?/?K]<Jd<+NHX:=HOR;EER.^]Mg,1aQ3\X9g^0b-+S
W4R^AfN(7dJ8f)+JIS+0c6OO_MCEB]:b;_YE]+62M(IIca;C\f_8cTHRd;QT0##8
CWM.3f24[Lg@9B_^I95YJ^ENW1PYV)GGFe:/8/P3@L0cQeb6KD+2CL8\NaP7#.7O
1/2fP;N5a7RDS./)E_\86^J6ObOU^@IST5>CSa#:?^F=R@5a=9IN1N9,DAFTD&IQ
>a2A-)Z7\GS3B<<S4,W,?>d+:d&;4>VB=Vf5Wf?J^Kg(?a0W1gf59Pda\==:E6I^
_PR)^bO@7;+3T4Y5X2(S^T#gZ@W9,Y_d_Eb2<^W=V/c[I@Zf[JDCA.PaQ<DdL-.6
g[TQS56b<N82)/)JEP&?#IG^F=^3H@PC1/-J9/fF,;LBB??(/\PX-/Q)4OOPN@aP
JS4,f>].:M(7<.U86WB<(PK4O38B?J#DJ44e25]\9X?@=g=QeI-b=;Mg0Z:4(L29
-b@4c,],&+W((g,EVUZ:8^[9/69Y=19Z@>R7.6Bg&7/4B_ZVgb7T?SAW=&>0ACK5
R4#gC;]C#)16F)EV0:9cebCWJ9f@)=GJB_&3JY8Z(,dZ&7NA]CN5(;VNHVfJT134
/#/b_YIT=0fBB7\IVHf[I5HI(Q969)Z3?EG9^LPVNSG+TM>GN4L\\8E:[33&F)1[
H9TB0BRJWXLZ:TfP;U89ELMTA_PG.C?UeQQE58(S/NaEE9f\#9(=SO8IO9V-:&M:
PR_<X[)a#gKL;FN]H:?@QLH7-CWJ=c[^U;_UTDM,71U0dET7GbbbKE?gEWgWdFAI
a6#],@Q#Z1R/_F^=I7)&R/1Pfa5F06MJ>T@68gDP)cfQ1DY/B>:RZU/;]\)TgB.f
<KVJP^C69.>YCCL[4<H=f7eH,0XC4Z)eK,R4^S+CS;+WTS/gf-3<ZJb47@?HNfE@
S+GdZXcf24R_R=V(VDT:BCV:#S/&Q>=2(FSR:N80&OGced?1-U7KTGcF5L5EdaS<
bf24b=L&?N^;.MK_PC/c1bL2HR(c_2_Y9/U@&MDZ0f/+?gL4\E4eKZQG9g^<[Y;B
.7XdgN;@A3M&I@aPE.dJ6/^STd3]_+V_.2?_EC;.N8&2a4RNJ6T4Z1AIJ49?7D98
EdZ)GgNZ#J-=[6PJ41S/4IEDV?]4#+H)EW).J^,<-@f@a-C?NcdgZb8MLJB_FUT-
Q3TK(G.L?284+W>EP#Ra()1#<U)[ERY=Y,e23(9e7YFa2#_+V/c>D^+7:FfV2a;N
dX2J@?Q-LJQO>e=e2-O_DKcPcPSM16(->(]]_97<.\7GD65.FU,IW=c\9e3HI@+f
eA8?V[2E2T:&W.V2@JAf1D9E\.[YU>W&B@P[_Dbb]Ad6+H-F0&]9TCF+8OW@-&8E
()TeKfWGB2#[F?(f(_(]EX_+G)@G>-L&KFOD@P@f1MTX25DAYX1O+cU91I5L)f]R
4I&>3?L&f/#KG]N/TCXQ4KA:gQ39^#<g9^]EHEQc(d465BH^-fb)fZ)+AN340G)b
KU7^WOBW1#FAg=dS-)U[f.3;/eNb\1[/DZ34[^;HFS^;4Y[;Ge1@\,S&#VTZ-OC1
_M=;?81a/@6Y_:Df@;/_&]M.4)7==1AeEcPB,U]QUS^ZVX=P=Mg5XJV1I=TYQCa_
UH\P^FS.)-M_0D6R.\1P\Q2<28#WaUGTCSY_D0VJ0\e:PS?9bM5gP,\WA2JP4X_(
Y(L=e9/H(Z#4ZN.<3M36-K5@9M+M;WP8EG\PEc?>^V#W@P08LZW+2[VgLf.S:fU0
SAU1[F\gXCGM6Q\WYIU[&5HD_1;>7+&e0b9<S;XK98Ze.,^BV=Y9AK3X>RZ)95^f
EAZ->Y:b7U<X92L0<]d77>=K;=IC1)7L(>b,CQY:A8IU,):III@)C_L^)A1e>[R)
K;9Z5J[4X38_PY>XGT^58[HQE(E<?8;21-bg1C8dH1b_A?R56<NZgUU1>(6&@)Te
d1XLM;Z)f:06D#B9ANK84Y68=M&@d\JE^^@NM4;-D9#.0cX#^Z(#UU1NUYa.M)GW
FT?e72L#NCB2_3Q)Rb3]e8Q:B80eP):GG4[[R_#L&HVEHa+:O..eQ>b(MH#-._YV
:??;840+SeP]1bO9_C.4?aEEL04^L//-=&VG8JSYCcSD[,FO^.aVCAN/XV7>B5d)
g9]Z/T?D\O;J+T^_bY(@;WA[I-K@d#FT<Y+P_f\7UGQH.Q0ZB,:Id_e+=IcGb.QZ
/R=cUV909aVg:,Z&4ZaV?gO)/B]PF,aI]=OA\a:T(5P?&NT[/?cBb\bfGbFP^0_V
],D+^=+:RDZ-+LX0gEc7>3K\g.5ETR\PcTWOT<-\E&:925I(SW8fB([I#1[28A&[
>DF6Ef0[Q214R=M?8\M&-d1;?C5,]=?J;O0F)O@Raf.L_NDN-J\.G=c)c.>4FJV1
/fJ(8G)XNeX^/MaKg53/R/0ICeIfE2_80Ie8SY1JM4:+64Q(#R<XbI:3bFIY4O=9
eU3e]<WY;BX:4dSAGK1]YGS._f2&:fVff1C;S)QW=XbZeZ&LHb-e0DbJ)A-+A>8d
D7A[^SK07&[,>]-?O1JZ3P]d82DGW7)/X]W8@e-L8SRdWC-g1:bTMG3Ve7bd02U5
X7(5cg&T6Ia@<9.HcRP;ZFYQPZL,dK4/<6H;OPe2Z@J76C+a2b??PXQ;JHE^X5GD
Y=Hc+GO?9(_QIP_V^VI]-THYZ[D#.^D-(6.d(]#FIEf:+S_4I-e90ZI7\[f>d+bg
7MaXaeCgK-cJ7)<,[8SG_S@6Fc=f-ERYQ+0E/Z]3AI>[A?C6bQ?]7c>ab2+3/0(W
MRB<5UI@SMP:f^J(-4D.ReR5P^RUR8;]d==#^E0JA8[_XG>NVa->61Q]bgY(OMET
K_b,H,]d]#/Z1L9gC>4S2cP&5:T-V(83DJCMDKeV+TG7GV0GOI[RW>c6HS#RFVU7
.WdYLN8\#-LZc_FY(\YdVc0]O_I?;6M(7b.5=,-gC(KSK#ZI;E)]>cAPU>SP/SaA
BGA+TaJ]K=@TYbGO@\])\e2AK39O7T2KLY?0gbRR23=,aV)WQ?e:;GQc;HQ6Kc]E
HKK:G=[\e9+TF3L#P]ZPFBU:e8&@@8<YU@9,V.PTXRGZM/(5QL4HcV;.=J^C^=65
d.=G8C];PJ3>3C2S>Y>Za_VV=<@P5AV_MQJd.L,7YFcICCTK@@;]LRF4=[^(C;dP
6E4a=/E[dY?G?=V^O5cbELg0fI<NfQ2I[HU2\gPgFOW:dc:&<BDA^E7,b(7b91Da
_(aXE4OV1R4G:HFN?M9NH[b6:^?.DJPJKPD:G\7G87+e?735=P\)ZB_[.M_7f50)
J/d./^(=.Y0>a??Tb&\cSH8.c?UcH)bDX?\B(SgGT#U&a<<Y=1#NbSB_>Aa1(W/M
#.W/1N,g22fJUN,^MJRLU\64[b(T9fb/+1#&^LI<IE)Z@d(T-3V?31<(d[f7Q0NH
LBQ]K9bR1RNZdFf\+[:EdRb&BAQKd(AaKf]FC#=KR1FDV.D>P_NATVM0+Y(7UP,A
(5;I.HH+TSAf2Z7?8Z,+?=2G1Oe@X1WP08?7aV_J;K[J[\cY])QaT9A=L2EGG]04
.W\>LDMaK,cQ,fLCU5Z\P3B2;8Ffd\MYeA]CLCeMb7cP4.M^B__ZdAK/gK>&f-g+
&\IFf?#7e39WQ0#._FY_Z-S#:NR[Cb336eCIe?U0M0aSG64]#59KX.Z7=]G3@5Jf
Da4H:.g175@M2bd1@MFMOdZBX@L@&K/59Q/ZBM7EFT;D1f.6_+?&6_U@9,?.g(ON
T[C.MSg&\)CF+N()VeOC8_<dUW]58gGPJ<aESWBY;RR#:]U_DKXRMb.GN:I13SQS
dX62Ee]39ZYS7ZPC<gRcFc#X#QP,4<M3];b6gYO1L:/^J2SCYN_aD@2IXJJ0L1P0
f=:##OWWF6P@>-Z^&41N&KN^?>N[?a+P4&_fVC#C#T-/@YWbBcE=3Xb4f>]32=<J
\.gSgg<KXL/<@X)^T-LFJ>0(E6BTXWX6MI-3Q,)_Q[Y]&Pd-T3-\K#[,A.eAH\9B
XUI37_2N@96_.]Ad_VS9(6[f8DPV4)EcUHG2(:[Q;I@K44<_9b.)-==\>R,&(:-a
]^-&YD^DAN/7<X06_#H_-DV0O:e^H?N,JS/H_BC/V80;CV&>[7R?f;N>OMSZFP2E
?Y^#b?@bLd076>0WL.0FL;DgN.W@Z?,1g2[Z+(3c]E)71(?I_Z\M6LD^F0:5.cga
JJSA^0]^@B^dK=H3T(&0,d;N;GFFWNe-EEdZ,d^Ig9?dQ5bQCKL^GV9)3:PHDX&M
GCd?adN5Bee>1a:Hf-I;EOMY\CA@@2;F@+#S_6XAQ2Wa5^.)#gPHeYI]5F^H_c9#
cLFAd6f]O;E&eVW[_LgWYC\Q7KW5?ZffG1&7DC.Z^)7VVI6bQ<7:6P?Y6XM=CDGQ
K(bRac,d>D5Q@EQP[-@U3GSI;=b[REbS:O,HMCK+-&Mg070.,?A,UA(Q\L^K\]/+
dB8WYFUbH.\8QZe.SR1Sb#MZ#_/JI\=XEJ//b&_.Z;\CO?H1]:(X@<.3FMaQ1P48
H+-Y[:0)5ge4dLcG]>O1BHYZQQ8HR)KFGbB@d>7@=[dWY\Oe>gEL7),d+],)0_S#
8Ya<OWG_IFHD7[9B0@5^cXM\bZL(0[GVN1UH4.?HQH^GQRWSUPQP[c,K\a,K;F]O
8MR1Zc&D^7(J<&+0XP7@cP6T?:6ARDIEP=A-WK67E5HBT2P4XWMZ->MXa7ZWJ_D2
69UNT2:E.OBWZ/#/;Tf19@H2)f1UN^M;>dD0^@05:6O79/^g_ZBd;_Ka4c(LD7OZ
CJ@;)ae<9CS=ag,7A1f)MgLVD:9#,8LU8W,f2(G4=/FM4DIQBRM?)X](QE5]fEdf
ZBMU?(?ZMJ:g&=cOIJFS.XA8:;f=(9PaIgOX/5fY:1d8]VG<VZZN&T7;CYee4.g+
TRM8FM:T7bBcV^:bbC08Jda(N;^J/XfY0QMPV1df6]1(WWM.K02HW-,Y18G<NeC>
PNgR&BXG9fS+:YB18,).8X^RYc_)408MQS3\EU@VE6/O>J<1]0J@.5]Y[+]A.Q_4
M]f)c(6A-8KXY2?6cRWQ&^P008g6HYH&O:D,9@FVLMI597DY<Z8QJZ]cM]E<1[V[
cA[1#:8[048/C/Zd;H:LbbN[a+ZJ/BIUT=Ga+7e-HHG?,Ka?X[,3eL2#d.#-cM06
5aaG15S+3(&+FI7;S(5M6=A(V&-]E&,1I#_2ZK<.XT6^[AA[D4G_49AKVW3,?,Z^
aE@3S0bZWV].U0QD>4[bV72EB?45Fd2V10adL8V<TYaU8\I43V,M+T,#:#-SJ,/1
>#P?[[ZGVa^=ZN+.Y+P8W?Wc;\gWO,[3Ib&#aZU-.V_QDG4(P2P##g<Q^)1U,2ce
2fA#V:-ZKPE4R:)1I3L7F46d<L-=029W\M^LQ\@C:Q)_Y9X3aZW>89YT4)cM<d3Z
?Q7,c>AWLT7#R5;ac-eC,:W[9Jb<VKFM?4cI0@N-TJIA)gA\M67N-M-9Q&J6eAaN
(-+>4@U8XL##H?[_V^,(R1Fe[NN8#CUEA2=38#>aZ:2dW8eQZ<4/0\AEPK.IBYLH
<_E[]KgB4+52JNIIXZJH8OK@HZR3FTLC0b_H2EP&P&:VNXK/(Jc;#]cEL7[:eF4H
,eYB,B-0)g/5:E\0\7W]2YTbJJOD&B/MR)FR=g82b:/O;gN@#/Jd.>C(C3I/F1Ta
2E/3OAXGYR-]8D754HJ_#HQ6I,HX+6+H1[.+ZXRW2L#E]H,7V;0DSBBCGe&G@ef9
@-[2+C<-cZe<gAJAUOe1;GOIDY-VJ4H7Bgf1GU]C2JAZQ]+\70X?OP9AM;LE4NTJ
N.<.#e8,VH);I&1<Ob+g:dW;BLU(NC:8DZZKS;C=B(>+DKDP^&bE,6D#\;SCB(+Q
;6/LH&cJ,RH^3)E<VJ@OHHKRCd;X_9U^bcE9_&&N):Z(6E2HP,RNa?gbT5KX:U&C
O,PfX(\:;Y_QaE-gJ;5O1Q@7O/838F8Dd6U@UV>/6<QagTV8YE9;+TCgf(R6]ZBg
95gJJ8#dP.f1ZOcK.])A5cb@\ccF@<1G^/4@KUWPDJU=?>#UL,F:]fV/AFF6+XI_
0F=2Rd0EI;5WX:;KC_Ua0U]DD/.;e))#YRa#4+4.7cP^I8JfTHTH9e/<FOgOUE3I
?3c0)ZTD^;6A=WcXf7P3E_PE1XZ+JQT<DJ,=5:e=(5UK_5Ug(2F9;b(^KUVgfV;Z
XXRa,<,PNbBWM9aYab.5]BabOK^[ZC,_/:>_D^^E1Y_.6P3A(;TFDeCJ()ZGXe?=
LOIXFdcJDW_8ddQf\a)W(J7HA@5LPX=70cAIG:H<.<I8a9Y6271fKIcbDDE/K?J=
)e[O^4O,K6>AT=ZcK;]YYZcYc0SKeP-7+L.2UMHfF3\[O^1Dfg+_._>Xc:#B1bf/
K0Kb_?B3d9H^IG3?0Wf>GI=P-V2f&F_?I[YY]4f\V6KNPWM1cd366K+2[1&AU>a?
VVWf/?1>&cdLNPHS+Rb\AX]DM7MfKNM_RR\)QcUOOKd#^#Z+P/=Tg(_=IF;)\8?_
R=.KFO1_c18b0EB2(Z4#F<]]AEEKb-)^L53f_fO#-/N<5D_+5DeU=<4+LgZ[Z@H;
IgJ>\#;WKMV+3Xe\4fF14=GZTbT8&_^-052S7XWR;/C3&Oa^,<Y>GTM;E_EE_Q?L
TPeNgC)Cd?[8(G9gP8&]2aJYfCKd9>NFD0+1;4a?G2G0;MB;>?IJH^@Z5Z=XM>&W
3D3QS7]e)(Y#T]2:)_d)@TcK,)efd;5_0aI?Rf=Tc9:8?790..9]8Af;XJ^\]0I(
FKY?QC@=)X=.b-Z;)RLa,I&e_+;97GVX76c02]X;0#1F?E4Ce5JI?.[+5&5.7&[X
D(=eg4bD?O:N#^>5gga6\(+46Q0QEcCW:NeT+I;CJ-]^7UeFP;T?4SDL^6H[PG[#
GSRLgRMP1V])Q41+,ZdReFU^]cgc:>VI8?=QR\bA)&R.-8Y=Xg-,4>GfZYddcD2(
+V;OWY&_2^AW7@Y^Fe@>U/+0,bUgI:WO[+O@28Z9)a8]2IfD>PE+8VV\J&Y2E(d4
:-E#=KfE6b@?WgPTY_G?(R#>,);Ma-:^M)R,0f^\=#F8OYI8_MD,F=QKW9QAF)&3
BC^.X?TEDf;FgYaIR2;;91bF6e(?<MbN[Z\YBVRC<)VPQ0T#N4VOfR469/]@d4-C
>/UXb6AMU#=Ed#g6,NP?)0=6NN>d?M,J;e/3UEGW@MaE1M9_5X4<Q8N_SP]76Y0&
#Q5gSHE+DZVI[-OTYX([#/LH).)].W7:JeICdLQ(MJ:-+<e4;-#g(P@SGBVE9Uf4
:MGV?G&d<\8S-BH(g7dNcT0)JECZ)XZAd.96Sdc]4&&:IN?WB-B]OR0D7TdCDZRd
JC/L4W92FJ.IgANYJ_DNU^FV@0#AYO_]5K;16R5Ob@A3]3S3:6K4N=U<abc5ANL@
&D@WAOB5)6IB4&beT^>=+RZQZ&9_P^YQ6HOQ(eBedB/I&W.Z:--aG?O,bUWYe[a.
,b+b485MS3#HFYaP87-P1+;BJ&86UN,DQI8<1+6bWKM-L>?EFVcIUG((^B;9F<F^
R:I#UQ0W)^:bDMR4Rf#>>_\cYV;7T5]Z=/WYAT0d_A2W/?)MRd-(L?5G\G.O4)c:
;JSK+Q(JM-AeF5ZY:RBC<AG[J(PdBe+>TN)\[H+&HB9L4XO3UWaSSVL)S(9.JYS.
VT8A^QB69d[/Xad;5N>.Pf\N)&QXN92H@]YdK7@1@]4+fPa<T#)F@N;AfJ#d_6_6
bL=OTPcgUR;IbBU(G#@V#1_-:HNRJM_,+1PYI3gTTS3<(]ZGaI]J<X0Y-(HGTGNL
M1QRQC,U.eMG1aWZ/(B_SD&[RHC:3eL(\S&[9]Hg9>L14ST>DQ=3:DZ>e:[FGAAF
SE+IINf.78<U7,6PT3EL-SX+0IYQ,FLMT1d.+gWfQ2&-3gC[daMTe:Y8<MLTU;LW
D^;=7J)M2FdgO@gedO4HJB\\V?L4@A5WM>BOHU?#d^VX9W29Ig]B4P4PX903XI:0
S^gb;aTEeQ(NPbAF9<E^HL=ef5?d5<4S=gDIb2^Z:C53ec1QAGFDVL2\g:(;_Pa;
,/?[3KG5E6dK7;Q2QgL0DdYJY:)7<N2^00#9MQ;f+cNP^-0&?BY72[,f[d6f<TD1
2E.QQJA+WS#>dd^35Jd0]]ZEc0GJGdJ_84RU0;V.(MZP).[GA@[ST<&:^?PDM=f:
2NMYUUR0<J:?Qc>-UL.V2JZ+TSgI?4-1N?Ja&A/f5^[bJ/aa0>-_R^FHQLXMf?+:
YU(bYR979Ef/B/=#X8F9\/@7?EM7(??2I58gJ.2@HNNc_@=+:=N]@I@GV#X=WB6V
c.RG&#\Q@;RdS=3:KIRCHBS#f87)Q;O;K9;ZYD;<Rf60M@E^PgCNNIJD448)EaKW
R/\8=0[e49&5?QF1GGYaK7S09?=\@L4<f5L0NC=5bX(1K>H^6A;SeOSAD9<CIP\[
g:DRSV6O@#89f5aeaO8ZICB@ebLRHd=GF3&0XC6d01e3-48>2E/>=:)5O1R-1gM4
9O.0B64OS9^T,bK@dc@FR^I9/f9Nad:;FW+dRGfDKO&P])#@>eN&ee.0\Q^(Y(A^
_:gF9[7e&FEN]0X-.GG@=Q[)C_=VM0762F\Bg&PH=<9-P5cJBI._)N,&^NX=A5)D
=C9+(;C^g97TV1H>O,0G8P,^EINa[O0OMJFWHa\UL?U)HMM3V2EJ4(?C?BJ?C<7<
]H>P8[^N?b=QS@EUQf[&<,]?5V-.(]@HS/B/#P-@O4F1\SDP@O\22(9.VQ0fVUHO
0BDL\S[E8:bc;UT2F^E63ZIZ=/d#_P/HB=Je9P.WV;>W^,@T>X>9:O5)Z<0c8H5&
<U)CL;0T+0@LPDT_6PT6?S1D,aW>18fQ0g,;]a@D6cTGAZ.?2c,D+BaVS@b&HZ=>
/220eb#K3:dH.,+01F/SR.a<cc;PB>:4G]V/RJ/J^+N@UeMX(.0OTEVD[a<5@8+6
g8Gc04ZT[JR2a;AaZL4;f\3MTT.BbK58))#EdK6S>XeP#?LK)4</X^df+3=-;@5f
d6WQE-AEcW9@<,(7AH,86MG<Se5NB5\731N^N&V=:?(f;LZQWGH;D0J3dSPG-X^:
4FW2+V-c+9:)6E)f4[)RD;X#SJOF\/)e)cG^4M=(f/@QC:^?E[YEb8#5Q<0<4]3^
Y<[O&#>1(<gZ9bPMW;1OVI43?6cHCBPA-@Rdga>f[8^6^,V76_L\b[)LeR@(aa2U
G=W->__/IA2R2UZ&b,OUG9Y=Z;(PWP3Q_e;SCG722N21,I@LQ]T:CJcF\Id&BQCb
_+XJM.H0PA,d:O3E.6Q9?8N9FZB#?)b=GUZ)g.J#=cI3EeY&TCS/G]04[F+9-()4
TY,8^;gZ&_;f1:26Z5Q=Aa[V9#;HQTe_J^A6K0NQ&B(8C61O=Z#&&P=BB\J6-1Sb
,QL_0bFU1AX0W_EA-[)-,QMXJ11,I94-K-=58=JZGITYVZF^N;f2D-#d4KYR:?g4
CcH88dKT2>\I9-e8fEC:C2I>d(M_LEc1UR]L(A-^M5U:^bg+13ES2J4[42Q<d^C?
fEf>WMALS?A3A7Q[A4J]R]dOdU;\XAO-^_9UZLLf-P@MZb\d;BT3TQJNecSQUL,K
)D@^[^Sda2d[(EILaR@(de()MG5+]HAGAGY@5A3S8)W=<VNNAUYOD1g+(a1@9<a#
;>+;7S?/.bbJF6e=fYIW?7NJX]LB)QPQ3:8Kb3-1=F.V=d)c>5^PK>&[IV,QCQ?C
[4;&N_,1RQ2Dc=d#SQQ#Oaf9UKDOJDBdAaZb-ZQDJG=(6WJfN;98+3/.&=a=+A(H
3#AIEV]6X#=M-I)230T]<U3[a^E;[ZUVTOVDN..eZeNPWgagI1[;5<>8TTQY:F.B
@7T+KPaSb\)T((^Df6f^&+OT<_CF<H]A_ME97)8TDf81)d]JMJC087#AgVYOM<db
R/@0PN_I__c?EGO/Z/=[>L/N8J;UPeM/<5UQZNXGH^,A(N.LGbFba16UK&20dD]6
\147g7BcZCY,,&I0EMT]61=d1afBR4F[SGO#Eg^25=EGJDZB)_X+g_KgP@0INTID
)6W8,8K/L/U8>Ue<[]0R]_+&+6^?R>>B,]0:N?S,(NUR]fR=@ZBb=J[_9:YQdW;8
IR:X)8OY.TVEAd:eE8+eQ(gWYM&J+>QIKNKQE9_=]V[0Sf4dG=GafE-(N5]?[4Qf
SaP;-HeaGM3W_T>Abb]P#>UKYWX863bK9[/9CV&c509?<@K]B<(28a]F.DG8UgVS
T+=OGQ3O?]fW<+Y1Bb99e/6GYf@G-6HX99/A@5):M_E#.42-f&gB,5P=RWXgC(F@
K#>BY(a>++T+HMIcZN#MTYI7<NDJ=eOa,]B\C@WIcREMS@?OQdFBZP\&V.K^WfFC
_FV/)]f9G1?T<E.IDJ;H?@U44IGT6U:#5[,[FeT:Rd9.&403^\#JTc1,1Q/K-AT8
=I6TCW=If(_W5)U/Q+-gD.ZE/#a+YGXcMX]II/5:L5(4JcG(7MbE9d+V]OB)SUBU
A5#YU:^1c>D3c[NY\PX;=T3=U\fFf]_QE?_6)H_a^X+SF9/1:7LTH40#A[^?XG05
B;(EQ:XV-SI?5#S6_Q<1/aE+,X7=b(H_3U)6=9#2H06:17IcMDV<adf,E8&CGE8)
JM9KX];:)9c#JJH>0UXQ0>+gCKB6ZT+.8,b\E_D((^&WNZF(c4J\=Q>N&3;@91T;
PfJJ?bfTFE7^V5NWHL@3g@ZeA[SH<L&g1A+Y>H)=0YN6fCX#A=;G\L+@g(-ML_-6
6ARR_7^>)@^2+JH4GD)06\.+YdM\6fHP4d8WaG3SHdIe7NZe#U2WJ0=,F>4I>AWc
A7K/N]OL-F2U0Z<Y>eR]E6M>0a]a&?54L\.WIR11FLIU+E\gA]0-\;JXfaJ@V;LC
4M[>,#PL,8fO;AS=CA[29a0J:>99R]^^?,@->&CVF5Jf+QJGSdbdV&3T#?HM^0Xd
3\:XTW0O4)CV[J1cV>[CT(T&:cTV:RG#[HZ5A&^G=4N.Y15EC6.2)QRT=95KV4W<
bcP=aQ0LQL3)711gYUZ521^I(Ge=AN<5M].RH8>a(&M1SF[O?71XG;U,c3OBJIOe
KI+WJJ#b<FaA]S@2P6.HDfOWM4+]\dEX1.LVb<^AWPF[>J,ISd1)<&a91fPSaP/S
5+dE&04^Q_]PF/;fZF9-<N6_g1=:1PdY/T1YdIPCZD\>U+7<?c.M<@0@/,=gH58c
gXdMa3=<.KeVUg.=Y-(1^3(KZ?=?a5S0]Xc[T:GG&(?1[aTC5KDbVY-IO2SN)Wg8
R/R.2YWM9?/TA<X^33RI^Rf<./P\d(&NGd&D2MHQ>3=]XILNG/R+/9Y@W^02W\3a
6,.1_/I7GRd<ZPKUM+Z=<]X5@#GGCd5AEL9-fNF3)f<=7f>A[e_gaAI,[P>HX0MA
#V<;Y)-fJT+NR&6\#6c,M^M[=O=(>F>gV7H+CLEI[:L66.?G<2^2,#R1WZJb:M.c
GLEJMd:MV?WQH[=eXF&75D\>.+ZAW#D^98V0H[YIW?He+gFOI<YB(?Pd-CJR[Y]W
01JZ=U-LfeH(;(YVL&#F:W?Y8(&<DeO#WF24Z.S1;d4A\WG=4.g.QJRN9IJTJ,Yf
B;(^H2M)]Ufe^M-8PU\/]QObVB^43-a>18D@S475GfJDPD7POAa7?L4bQ<Z;dQ-5
:ML#_ADN@L8W=R3LN0^L9.L]QR18-I?>&BL_=@f+9=1SRB9+3R:cV@XNX]R\7XTR
:I(a)3\7#WNb6KM4T&g1VKMPedCaQ10=(F5fE/dT720/WI,34L[G[9=C_&eOcZEF
?+#]AZd+df-70W6](/LQQW#8#(45QH?O=4PFI297LRI1\A[K++Z\7FI9O]Y8IbAa
0:A7L3+QYJ?-REE(d_NWOad0IbJ\/R0@68EBKQKU+1a)<63J</:K=F4F6FU<YY+)
I(:@U+T@W&RLH>beW2TBHZ64[.cU3WJ^#1O:c#:2-0;5;G,N&E:1OeJ-A[(:WK5H
H#<&X=Ue9+PP<<Xc?M_M&QL8OGC6GC\]2]GKR?J^QBVQGMa9LJ7?)BZ8O0>7.VDK
R8LLV=&+If\ANSG4c4T@9;F&>YEC&)NI?cg30GXA^DJcXBfV[3ARc.(IHR30D6L<
)d32a<L#<>E1??H8fOf#gcEM#&GbE&T##RePPK9GS4S4Q(BCbY^8)gWTWPFQ_Fd8
2C@@A@bf@.NYOK,dTXgL:.W\4^Y1W.UI]\.KF/-6G_e)X[/fA0CC&J+<(MWR@YQA
gB:U/]YS2:.7;&-V_Q8cH)T9aAKUVU)L_1TMSGGUCV5BYD#)PWJMDU@[P&-@02?<
>a6f0S)&CMMC&691(WSW1)L=<ETTN\I/?6,(bdX1^>NH2eR=HTRC^3GWKMKd;.Z)
;b;E_]V\[7+,(G3#<f5bTgLO]BIf;^U?GBOS)Xa/30bg>N_46]cadf=a;^UD3SeW
P02\aTW1,Q^GB8+NUH9gdGC?W5?KR97d8JMgf=^Y-+.UOaa)R6[DH=F/gCdGDBU@
6daT:AVPgD@[ISW:1Dd77GN+NLX_QBU^D-f&0K2a5-.])U06H;LJ)DV1R7fD(2>E
a<Z=[-ZWEQTY(VOe2@JJJ#J&J@c]Nd<H-SWLDMW5g?YV+(LY-]I2d=I#UgJ8b:c1
C1R,Cg7b;-7Pg7PBH0eT0^1Z\?S3E3(9W/(Y\,)CK\_G?P_NH+D#5D0gO^&.J(:Y
87D:=3TYL0+MUF]W#)g>P-#R?@B7XPA31b(VOX/Qd^]3I;ASUVI0[R=a.c7F>]HG
M6D]/eIe-3ddBW@O)0>G[Q9-=(fcUc4R01?Sgd>/:b+QB]=]@V5\IR@RF=Uf&][<
bDO4eRR-<,/,JLRY3)YJ9(a)>OeB<H_B=1^_HSgBe8;#LKI=-XfHDEQUbT.CT4=R
gLfNHM]&YUa#7;TO-J^&gd_+Y(Re?[VN+:<=2-^XBQZLEe,dK^SL@2,:0O^HICOO
G<W].?HLcc^6XEWUX/a]1WC@C8].Ka&AAQUb;_/T45bZZMANbd&E8A[J6e-VI<#Q
JLdLI]5_B0#;T/f?\;5C<7M-bfR)7E3@cA^.aWaKc@Y9=ee,_)U__9C,L5N&KG7b
4)b43O,ZUgWc1#bX>R?g7S,L().7,=2&[^DG.CP>O1BdP29).,LB5</O]G;^-L8#
^6VM7OLCc5.CXDMMTCF11aJa#,d)E.RL1+#Q>;E<-?<+f<(WfU#2^SHWE.c3LD(K
g?[@dUGL<71Y&@6S607ZRJEMe6T=@g\YbOV@(NW)FRQ>6V2VcF9=A6[;9>gLC3JV
G2;-Rc5,4>#4197]LZRa:).Z6G>DJ^7(F[3/GMJ[\e^^)M^=GE1cF);_KXf)Z;-(
=R&1LeWBZN4\RVOBf[c)Ge:ZI<DL]bOLFT?BOKO,P0d(fT]Y?M[X82d:\OA)OANG
Q;_=GK<Td&Mc60Ea(5<8,B^:?]#11[ONbgaX@8_4CNOD2#X_Y-54.P>gG^NRFC2g
79HZ124,MX7aBJDJ3/gUfJ#bD61F<<5E=QLO/B6Y?XI(GWQD<0S+U_YV?Y]Ma?1S
4-J#<;Z9YR@Q=DdMc9OM.a^0M@J&/U+Gc-;LfDP>OGUa/fLMY.^=c:51VYHZ0/=A
\Lg/:;Zg+>AI?.N^@P<@ESbKSSJAXg0_D:KF2>[Z&EgV&f482I-M,UH)&FTd<+<#
49FI_8E<;6CAZDVf1KYH,WIfD?g-A\C\^D]&(>)d3.fZ>@SOLLTPWLfG<-ZEbB:/
?1RC_)2]NbXFAZZ]Ae7T6>A0EbEAH=Jb::ETRB:ADA<>2Fb,0BcK0>&cW9b(F4R_
gO1VRaKVc.::_&;:EEXE#[7>SBO:^/ELS9.NDRU55e#?I5--cU/ARA#UZ^5\^WA9
6=98]@ADZ_Y>6]H2#(Bf>_Ja253I[)KX\X-ZLaQeaXe004Bg;W6gLC2<E/F#TdHJ
>6SFWOZ\>I42[_>X0<<=10:7DJC11@,EMfZ[N/(I+dM\^Yc<<1-.);_DRAS9eN74
;H=M1P\XIUa1OE;AWSbH96dDVV_>cW(<C[.d:N61\f]3&Y.Xbc:)2BLaaBW(I+G4
d\2@B\SdMM\8cdJQ+3R\Je@?=VYI@>1dB&-]F,JP26WCEZBFgI)bH]M.Te[gX-IF
I;I.U3AFGE;&06e2gE2\F]L+^?W\bZI?Ab2V;95RKc&&^_#8HXcG&,0agE09]]W-
9Y7;O,9\S&D7HB\VKa5N&[I/b9K@NCNT/6VUCVI]@)\[LG=/AE.+2-HCK>AcT7W4
&?>,6Z3@46[eYVbCUQ53g@Z(J0S;YQ^)X+-.(/1TE[1+=R7f8,>1&d<OQ^\gV)N#
QEI/7NHB,\YM-S729e7PY/JS#dfE(;87]Te;.fW/6R7P;C86_4@OZ0TP#866M=Gf
1:MfPR:K^Y.HOW,A2(#9dTG?Z\9HTSI6De=63<aS5_Q7[01RZ<52f4=(#NB=VeR<
#EETbH6b3GQ^BE^@.NTD6N6#O\^L#J-c<f5Y185JLd,SCZW\>L7#VJ=SG0F?QE@3
RJ^U96U,a+D.)0/C)#D[eCFD&eeUUdS>YZeN&;NQA>G,Q7<2^UY?BM4WRE,8a?@F
LRJC11?;e?V6#;/N(bPg;9&fFD39RUM.YII(K_G2:H8Z^D4<B9[07g+;MS+M&V=I
GEO6g(TR@#3T(28&_9Y.NJbX280=[VgZES4WObPOb=beK@d8L9;fA:Y7F-8dOT@C
O2M]HgQND_b;M_YEeB0O=[/BIZ#_Xd598KHE;SWf:#G(0M-2CGANSf.Y<_)+8[(:
JP7J9H3f3_SX6?O7P9X&O2RA?Y]WO@#L-9PEV-@-=(5U?<e9D\,SdQC&QaE[2Tc9
GL7L0:0aSV?M_?48TVU+DYA](A8^Jg_]+EKc6&21f^C7Pg+7a<a?[4P=6cPGbd.8
PK>4BJBSbD/+@7K:g#&\0G/;_;e2dX:?)UPf?KUId1&@f_W.,[]ZL+a+(?\][>HE
(6dL&2A)HA0^@VZ]aQg<:/WObb6K582#J-)1(&dYPY3WGYDW?QYPGJ)9+YDG:Y9T
<H#77)+],+f>bOFbgAJ.O&)8GM>e_Ma=34BdD(OS>dd\NQ[E_+)X?8X52@;OPJ<;
5MIRWYc#](]M4LR)0HN^VLf_G/E4d&:OFPP#bIeb,1Kb^c66A)&0/Vbf7XP(N&UB
#[I_2I&ROKRZN4QB4ObNFXOE/F835bGF:Y,H^2gI(SQ5M0DF+7?H1WUKI6D0Y;d2
;4DJ?=E-/XSO+6F>XfC?gJ<]]OXN^Z/T+MUe9,+O4eUZG1USacQa6,8E/8(V\^#c
]-J)9GdO\(^KKUXMd0:K-c?N8X1AASd:>&:CF-(IYb77)NOE1Y\c9N#Q#,)5b)d>
US&R4W0FJ?(G(eg^<\3<B<B63<]-1P]cb0XN(-#GOK7I^BcBRV\Yb^bD2<6QeD?]
H.&S=XQP1+K^c>Bc:He+SU,ETd+,#EaRYC(E?_#0dcX-e4XD1#9M8;UITZA+gKGe
,Dd<32M6O2Sg#=d[D5b<Ffc^U2(N-2U7WE,f.N0M^3#BScL8b@F?=.F&>fJ8&EEO
cBWFQF8VBEMDQXP@S@5b[WCa&\=](aG\^Oa(B[T@VZYXZ33eU-H42?O&.LC]TFe=
SB+]OJeZ@d.YY<-=:_F5&-&bLV-52TWaT7R8YdW?/^2bJ9F#Zf<1>Cd=>_4@S+SR
S<b62E.#0;5I.TAD+?>0^^7;+bUIefWGD1[C=P7?,-ecVc=FN85W;Wfc/G3C@OeE
@J5CWaQ#SOS]+:P+4(_QAH[I,GAC\8G)f3V(4X@6:OB]I91Z.(U2(PF0C#<@XBLb
27_1GBP\W:^?XPV)&5CgGQIfg-:SAIZC\/cOR77aWU1SS2>2KBW1cK7RfUcbO/,.
@ZZ3X&0HFNb[PB(>c4Xa,HJG15R>dM4Yb_767??YOX<\-L0a\4BJBc,?T87?B3NF
/1P;7e1\Q38?:T[CIJ<OUB(+0=NFXW<E73=I63LIe23a=7g(<_J/JCTI>&.e^;1L
(TB:7DDc+^/TCU7FYE+;D81;f(3T4O\<PG#E,G,eC.;([Q\1e^?g6a#b?aT=3R5T
47+dE:d>ESPI^DA/,Bg2/?f&]<C_c.7A6/P1XQV-:&JaLW;_(Q3A6DcN+[8PHYWM
1[VA2M,[+)=4360:E#XcGgR?;:(Ae/4J[MMX9UUMLSQM&N\IRgGB#a#b+ZNO3QWd
M1N2;8(J7U2[<g/eg3(YYUA.^0dXFLTOLGTOG:/\:;,W-SD1ce3dbOWGT;]aDH@g
S8bEgUVK(X7UA[00C(W0>O#bFISC2M,LGINTGCWCQ\7<);;++3OHBae,>Id_11KS
(4]R97]OT=[Fb0:\P3:b]BUKQV5dI/[F@aGW)a/g[PK0G2MK6d@@9ED+;,1\.-/9
KSaRe>HK7R3)H,_;78dSDY+/#aK&g1Db1A)(a#D##8N:8d94GBG/dIY/<b(THb+V
-/b)[f0X(I3c.?ZdX)Qd3PI]LTZM#<+F@L6[f?+:d(0\6cGa.P.I9\Zc?\&BKeGC
fJbcOb<EbO1\fHLNBa8#9,.#E#YTOaBH0OQ-YCQLg)GX+J)XUc6\^_0a.SDMd=43
LRTUX1?X,LPY>KC^\S]&FGJOb^W=YDR:QZ[UK&g+JFA7:T13/O]@fbBQ8H6;KJaO
94Y7QR4I#R69d.S-2^6L1&+b,b1+JYUNE4R.9#\[A+LB#XUMQ_gEV2IT8=F6A>DS
Xc3[TGR7+0eZC#-SM@Jbf3Z43RT/</F[7?3,e)\>@F6T:eK7UT;;<c)X=@PVYOAW
P@/\W_0+-2=U[[UfGPZ&\#CU^E8YND:Aa9DLO:O\fbI[5^1MNcKeQZA6XY=QDR(R
aceKAFA72Ee/:/R_@N3@+=e\CGWV2&(_6Qa&a3/aK>A,&gH;.NV/S6g5RF<fCH:1
WU:E=AA@^XI(VE[:Lfe:ST;ZT#caG7ObX47a[D^<IG[b5^6H&8Y\.8cWJL.BYgPK
d@608WOe7ZcSZI7R2Q4SW&^=.VVCXYRA^6fQR506S)_a4L3TJ0_4,MgS=g5M9+JY
9fR^3XfM^RT\U)\BVL:ABVXPUNaBA<<E]dLBJ.]W+RbK/gJ<V\I7dOL=NA8;7>Z6
FA(,fXX@4#._b@84ZVR4.>,0GXWPV:c<Q)&,KL=4W_B&]FUOAbG6SU;Q,<8]/9I7
;-(]P3FL[1K?HTY=WK3>H#[W#Vc7bPcceSL-c,cW)ea];\0->CHgKNPCNWdNW07;
]S0;UH/4CQ,=F3fEY-f>?PG6EJ+WP/G-HU.bN#dHO[\f/OG#UH]UVB(DBEGfE\3A
c@FXI\#=FY<&XUHZ&4Q5::CZ#K#?7@4?,MA?#He:Wa0\##XXfQ2.^I#L);;Bc)^.
bACeI_^fV?Of3a-JH:Q,e-1XHKZ1Z?:3[X4@-5Ta/OC2RO(0,,4B1?0YBX+EO@8b
;A^NeA,MgEE0;HBZ\,b1Y1[@@?A:-@Vga9=,]?<dL]TX)JXg-P7ZIad_2K4^25M=
/?F/T(8.QHA&/PO#c2N-X9BQHUdYLS]M=<P/+,K>=Hf^dI==,64@.Yb8d0><9\,W
Y7ECR4T<dYQEbC/:FcFUYF<e>,CKRVU?:4U_XOA3HfUC0_,RaaKCJ=aR-[VT_?VZ
S(D/#b8\0^F9(@@5QJX\Z.0QMg0_5b9&M,+S0>&8]ePW=V^0=-:]1dODXd>O)[6:
;@K?c:/<D=\F<)a8:-2T::fbLd=C=++](3T29U4SWFXS[F]DA)Fg2GP.5>::K-#F
Y@bB006?IMX6.1-0Y;OOg/>A?a(D<X-:d<=D\dQK--)7#+KHSG/]A(H_X<^;3U__
)TM0W&XB72>_H)>FX:/6Q2Vf5Z\W2(f1P(:#1F;B(1fD)=7-e:=JcQG\0\\IP(cG
<4gL0?FRPEVJBMfb(,Q2[fd;&eD&N:TYdN(:K&?T8_g5Uc>SAQ:KL_0Y-_HGS&1F
I,Lf(WdE.9U9NAP_daWf8UcgSR,Z(-E.1Ab6g@M#U5D1P7K[S&e6T&?71CCC-M@#
;,ZR;AXA=eP\6EgO-VB-WYL^K34U5#3H5aIOPGXICg^1IHS73/1.TKN;11\NH8\<
&LPQC&2\<b;U9JH=Z1BI1,e##VN]aQ/GV6K:]2;#1feBH9Dc@NRRd5FPU^fC[,LM
8=F9)6fb&_X?2P0AL[2LMgLNM3];@gaWf;-VC#0e@+e29MP1gN.@,U+KbH9,DLS]
WSGUZe-^4/L<.F0KdH@[9C[0\>P/GC&(g7)>+VI(3U?SBb7)[f:e11[-JGQ8:0X=
cffEXNOC;W=:NYXAFF6I>3U9C;D:0D91[BO]BTD&:G^@6.b7@?Q-@HBBT+)Ed-Mc
,FUV[DF0dfY4.\YF9;2:a-bM-Q@e2#4M>.UG2,_FQ2G5S(DN2K#END@GJe5>;a=Z
RL@W0=4.4c.C9NYR]I?Y6--/HOJ/)f:OK#R))8(<OJcF&H=R]NdN,[]5BS^OCT>B
AaT5+O\#(D=\Y+B2::[]cQ2f_J5BCG9T7C:6;M;OLeG7)9B^0EKD3cGa=I;]H>e5
X<Ra#3T?Zb+b=ZSc+[?1.LU,:e-VaR+C/+GZg6^1:U(0#A32dB;Z^9J5<PVb)[N.
O2gD;Y^7X7(W#E\3@3/:+.Q/X@26L0BPROd,9B4b#&G4f0f:2?f16^?c&(ZQPCdF
WJ=HFY^DOT230V/VD\1b[HBdD-c,8g?Q\[GVbXTS9]=Id]_Bb5d>FTdF.AXBFSZW
X#/O;cc&9O7SM#IVXZ5NGE/G-3F1V3O5SE#9N3\H9[c@891OB0Ka6T3-AP2I>cFN
&:3B?MIa>CBUPN39[fcF\g1baVXU@R;LF/WH9AFe3V>-46I:\I_eSOG@:W.-V.K+
8dNJ]8<F/bfOcS+JV]7SKH>V<IMA_5=;&7VL<RGL^1WQW1+f0gXHHRKW#\BR[0g?
D\>#73P&d@-/>2I@9fg#(WT@YS(]LFMI_7T2VF4>\>(cC>TBGSW7OIM..XPKO30[
=U.cNX&gdcD&N#S,[6G;RLKUF/:ZY5&ga:]/UEB1C]=WZaWCGR<)+KT6CK7cGf^K
\;)5;SS+<WJ@?\eV5Wd#:d=a4[\Y5N&+#T4&XeZZZS-]YY[,,9O;0QPV]NWEE>U^
YbQOST&F#D_]JMMAQ/H/(,d7/1OJ6H(A27)KVFdM<AZ2I,D3[T1A^.Z?=BP\1:2_
gG,].[X3\\<ag1,76+=Z?([JV,0A,O9,1B-?4f2F1T1N<7+O/Ya(-aVL([De8HZ,
B2gC2,PM_e349P2T^)0.R1+-<+:1+;GBIF2C[L8W/4_/_#QPf7]bQ45G_<1,_RLB
?-S+fAcMOd;XcTC=G.W4NJ,GC:>GgI+1&W3##7R8P^W<87Y8g#UM._>&T05^.>1B
bPSg4]ZeA;\Q&2PC^Ab[IWSEbWQJW09+^3H]D1=>ad?2L?fPL_.fcD+=gbX96?62
S(T1&K0FQe6?/^EO^>X#-4?,P3)-<:O(T=Z>JSD<_1,Z+Xd&]7O;WbV7:XETIaOZ
4b:5)bJ/dT6ERAGMTKW9XE78fP<+_<IKASD7H05fRF,<8e3]H6/a=JM-&dVIOISW
DRO;I[9W)_XZX@T2XbM<WdA[/.@O&\6O>aLFCJK\bJ3fg#S<X)]:PA8E=f^dRacS
65L<aD/<.d7:]9[\-5=JU/EP_PE<H)HO^E#N0#+-&/UD\5XdgU159UD&?fZ\IM>Q
MJPMd/ER&^8@D@RI]gcHG;d6LZ448_Y8T0b\K:FK47UIIGZ9b;#XFTD(?b0)TB07
\d;IPAM)fY6C(^2WZ0UW6N3T8Ndc\Z]bKN3=(W(C&R)=+)>G>-<KcZIZd&U&^>TP
/VVV]g,g?Y<@Q_)+SV??M^R/PX:>,/6@9X\JB;<000LOE;3f.FPD2eRI&ZHJ5IU;
gIb[&/.VXF&;_?T2Gb>9(.dC..eSX^/XIN64HN7MJZNd#:KEGY^E82J5&Y&CK?7C
d<e)9_VC#B(cLD+6C_Jf>KfOZ)[X[d2_JE/61B[DCGT4+A.#&bE)XVdN+BQ/QX71
@F^#b_N:KNG/1(Q8/Q9O>aeCNe@J#0AV?5(;CCHO^\VcBQ77CIH7=cg:LK8+#YbN
=(_e9&a/\0TUV>+(W8P_1CK,]fC+fA0A)d0VR2>eM<YER)@W<.V]Ja.R]fMQ]TF]
>6V7XL?=g<\DcI&=)@>fZLTQIH_#ZH^9B#/CVFe62;\YWH62DV16L\6\gbR03VP9
1a4\GK76Z=M,Ed:OcG>dC]S[g/WV7Ud0/RK:]N:]#daMMMR00)#GLWAaP-FVI(/(
=>Vf);Jc8B+J]AYLY]d)?CY4Ea<URODd(Oe;]#D0fcJ:Ke,W.8??H_Ua/NN2F>I3
b^:Q5J5U;()H+0BQ::AgSFcXDXF5ZEWIKg+7J&\G.LdDGITcfbZ^N1O5RA[C#9=]
W?cQ=>2VP\\P5H8KHP:5:FPfPGE,:/W7&M+V=]:E,)cg\,d^02d#=GTZ159fY]SK
B234aZEe#]fF^eKS-LEX5)FCUPT0VLa__I_;XK@<J@VeSABQ\X&,&E@YCQX<XfE&
g<cM;&IX4cd1(?f^bOWC8G2OG4Y.MR6Pc4B/@^E)<:.75LA@6@H+Z#c);H8a3[G_
?(<7NE+eK1UFXbB]1eR2LHC<CcMOg,@X.5D:\<?7D8M,Y)10[3&M:0fN_2S[V-Jg
/)dE_dHULcQ,]Pd_G/7MKFK(^C[VN-f@\/gR5@>4&_,7SIX_WZMFW?7@KO4UZ:G,
P22e,JfC,7ML^cYQ35N?=;([Dc73X88.D#<.TfGMTT#NVHg61&H\\>=g6P0LVH:V
L82WOfK1Ze;EaLI<e@Nb+Aa?TIbX@3P/e[daJET=GRMCgP/]GX]4<R9g5T(U;XT@
8V0Gf_R#M;e/,b>?M[M8O;>Cc>H4g,W^5Mc-6(<SM4D/OOHE<[]0&17YRQVT/4BR
RP_;1:L-T18HXe;f4WUPH2]\3_dS(cd/;VGL3e[--KLbB<O.VLVWHS:U+Ye46WAQ
6Y0-/\R86JA=#R@\b<&(>L3R_-bVY_f/;[)EUb/MM98T+XcCW_,UaJ:.@,BC&/R<
g]V<KN.]S9R,Z,?L(fR51-]-(7;#[_V0CQ#WZX_XUR.^[_R,#8--LfZ9XV5:g4]b
TMe69I3b7Q>bAIb.7YaHKAbG^N6&cHP#,/<F9g,1>^KbcE(cL55SHR14Oa(1KEJ@
-]_>D_5^fF/>5.2JQ1NYS&GUO-N_B8&3QO<R)JJ-HN=HI.>.d1MC4f(AE92^3387
_</Z)O2/=V425XFb]_HbT;U@L&-J3GBAQOZ[]O8JL#Z0-c=IJ7b?G>&1\N6\HY+[
-^[:?2@>4LGO&>KEO-?LDIaZT^dLTS/0FPRb1FQKVMZ(B[&,N(TZeObQ.gO9CYM<
0fc=W6#S@[Q.VF3E4cN:e49c\.L_U=R_TQBDX<CBBQ1=:AP.#7KFL@K&)XMc(b1?
Z@J1LDP)X81,,e:=<^99bTVTIJC7]0-2IU,ec0[/IR)bXKZ4_QJM+HO>9:A7Te__
K]=;UGTTd)Z^c=3PW0Lc=AP7IP.XP3,TXT;Dg^0LMU[[8=J>Q@fG\QI0^HWMGQ^#
IB=YJ;T[:8@,&+W]JW;3#N8,]gB8:cAd>VQYeFfR/X2\Be,-[-B<PeH+Y@L)SUad
YfOM6fCH/>\+S,S1=F=@FPB2(f>G87<^NL=782\g+,P:4Ug,J-;9ZI8BcZdAQJ/6
ALF<S]DQ>GHA/Yafg:E:d07JgCY4OabX2-^MM-f-RA9_I4UQC.dJ.V?b]eSW;@Qg
XI/-Bf53X4(=1T3fW5)1C#/3>DH/aP\ZOQJV,B[+PSWF[)F)>UY7D<+1+-#^9<+A
Fegg8S],28Xf1?SS6OH?)=,3>acJ.:+e@0N\>W2FX_\MGLC=A0)dA7GTe)fEMeMX
-SJXX?2e5I88JL3aNJE&f2-3A.8<-UW:FS22[8G(1767dNDWJ8L^@XJ>=d>>U_+D
a>QbX_YHKPIF]^;?>#LO=,LDAFB=R62PXOU#[L]TZY^+10V_WF4^H^d0=O9FR_ED
)c^];61U^O(K[?REIZ\g>/XW)JQ=:^99b]OO\;E?<.3da^F#SI_dV:O#/aVIG#K,
e#)gX5E,D2DT,U6_,_faQ_H<]W(Zf&X+3L9[fX(=OXN(5SH)DON)SJ:EbXY[[:4c
HW7>)^9_;Pg5Xg>eRR+)<RLO7A&XRU(OS^=JYV7QC7f&WP:9cGg]^)ZdQVYD-Pb?
(a?)+Kb\Y?7a7c\0\faL;/^-<0>?VbT4;>>#SPJI3JK/70]c5]Y_6Jd>J<<3b_4g
2])M+:YNS1U^@?9#0Uc31TAagF\.1TCK0R5XeJSB,f+WC4O3]YK6>=-=[:TVKM>Q
\TCeeb8,fQUCdD-,X..=T2;f)E&VL-(2PG914X=b_PRM0,A\C4eK+GL0I@_X,;R4
XfBPGc5Q+g&S#R:NMG2,O-<&?6,O3cY+g6X\OS,16:Y6W#7S_.8]V)-dI:Qa01]L
S0]dAQeX)UR?K>5V\db0KW&_N;+Q()RE\.?>N7.@E(TUD\EPKY&K_WBX[))D7>O=
CJ\8CYg0A?AT_d]UW9,@Y/<27ZGBOTNf,AV:>W9^c)MR6/R4K\JS(4_@[@VK<FCR
M_Y67&H\0#2YO/aBXH:YDN@\FQ03T068+ERfBd\VG[K,Ie)cV?&DKY>[ZFHa\B?^
ePLK-G;VcfF2T:O1TV,2;#<FC+Q#WY)1S@a)X:_U)X\\N&RB<EbD:AE+WM9<bgM2
D36Ea)Y,_(WVd4)3](LaJfFT+PJQWaS90#+79KJ[\U0FURM(KJ#)3:U&VdLN4K0M
][VB+I4LCeTMeXF&McR;dHdFJWON<QQ=9I<L+H6f7U9,)Y/CEL_^I[0S@-,L@0_?
Pg?0HHF_M]_KR)>=SV\gY?<F[/J-1P5ee+@F<P,S[)@Z20P=ZaEJZ4W17BW9E6]G
fW:MAUg-7Dg.+^EZbY+]eZLE+/:C8V)J\+5H\DSLedTZ=UDd#Zd@fe^.7./\^0\_
9V>FHDR,36>4a7.<1B/LD&(4Tc=9-TBcaYTdK)E.4;QU,,REd,]<@d.0QU7)d>gR
.de<G6>N<fCOR5==:O4\\ZT-H,_9afFIQ1LaX#VJHNKYg3P1bESdHg,-VXJ_5\)D
=,^A-L-a-M#6[YQS7/R=RR=JD<.>)cPEOe;?G@9F0?LCJOJPW-;;d4Q(6=gCaY7O
37_1Zb5)9=C.^[(A:BGfgHO^ADQR,&12OX,:F3HJH(#9/ZAObg\_c\\+DEReY@P/
R+KW2fI/YPCYe_b9=gGA9AHR@(_BZ/=P7;Ba>@WPK1_R6?.J8K,N4a?2T((&H6EG
Zc+&Q2L)XGQ/N/#TPcHELD&CcDMORPA#BQ?_7(+N8#_?\eDM,JT4[(fH,Ng<@/a-
c6aY+X?d2LaeSf@-0F\M937M+:,/QTSI-+6.3H?db.USA;A[:RaH(HC:1JgRAX(P
WV+QF2LL&aYQ7)f2RV\-.TW.+&I(LU66RLgA/dY(5H\CBKJbX-S:a7MVM:[F4BB;
7.g.a4]WL9?(HffSa##\WFYL8ORU&C9,GBO)0W.#<,86_6@D_J3d=P@0gVQ3C1ZY
-d:@T06H5cJ]X(&@?b8[Q/6SGA:[B-1TG8?I7#JX7[6->gQ6(ZB]0+a4DaWObY3)
Y9RIXGIX3b6+[gFEOMAT^Ra5]3WLZ/UH0aC6.CLU5[:&07Oe(O8R62NfX6(NT<83
EcEDRS]CX3VaHSe<LC&:g=)?c_87MANQ+0Q#D>OeC\]/W7Y/3^VfXE]F)?;C8B^:
60JP@52;E\\SGJV;VMTPebS87Pd\OB=,CRJJ8G@\fb8&>34&JJCb5)(G=[,A_L4J
+M^XSNO_.D(5+e)F_[3X3c\.853bM(f(O5a>>]#)KX.[]EX8a1)C.\T]]1I0]aWL
cPM1OWadZ=@,+1>T;gJaELaD<@RGY:OO[XK_Ma\Z^>Y8(3IFd0JLA#T.[bUW[+A=
1c\;E9QgM>NJ(<2e2+LbP7\K2PM#(EFGOT)U,JfKMA,RO[];L9LO,=N_O<?^:?M&
&+b##cCIT0FG4/=\f5@N.EGUU<gKW\b[6VY39^ZPV9N<g2=<=.S<JBNW@>c(X4E;
3\>7_GcW(b3+#EH(LOVZdMbA.MbG?QP[F5TB3.g&^cfENGgH5_4-347TM?]c]QcI
/_80^>0(>F:]S)a]N863(2A=:dd\ZZ]]10-&7#\U6?V#\gREEUf>.=E7FL:bEA/6
O:(?e.S5F[e5QTU=dUFNE9Xa/6fY+@L41g.#WX<O<J<b[VZ)[K<\Tc\Z7L:_e_LW
D;-HVAFR8^JZ8.ON1V@N(=._2FGPB<&\-4^[PZ7,B5a];X<RWIQ_Q;7O/;K2@D;b
fIbF^7Fg;)H)4&bgb[.V:]-EA0eNGX>?ODQK<0F77V2=PI=7M^K))5P=J=a15?@T
;4aBC\ENF+TeV46e4<W:8@,G&0L7Sb8VZ9FgPe<DI8O4_Xd>M2^Dc/O;?&IV?)_Z
DD_EFZ>XH;3#ORQ_YMgf>0N.+fg[4@6-,3BH-8Ua,GXRGONc3FHBYb;^4a<&2\<a
E63Ke+RAB&+ST(H^6>K^\)Q4;eb(e34SfJ^48bUg9+X0RETa:.OC@1+>O\>LF5\Q
(WN>U;VNZ0MN1YL7E/O]Ug>]H59:aO\8:#R1W5g\8d4KJ13-)@19ef\H6HSQ-J-b
_?1+S&[f-/N]M#@<fIbC21=+gTe=/?OG3ZRO5]gJ,SSddV48V,=.,NJ=,<6d5NS@
B,JNde>1BPL;M2ea/2X].Rf2g]Z)QM-EG0<3VgZB86)b95<WEeGP_e[Md5[g#Paa
)E3CEH3A?#ZYLd5B:V]&@IEK<=Z\#<NY2=0V48B_<F6FFT;Tgg;)?)Se4\W7a>&I
f:?@\\+J53J?AF?5#9SOON3=)([XZF8d&MCGc@EAdKb68@S5V\Hb\e&O^8Za7V3-
GOa(3>:<VOI.JN3F?^#GX2\QS??I+B\,-b#H8G&_71cD<5+L)NIWY)-1XS2C\Vb7
STUH0gK7dBgK2\=B4S[(,3<8>Z6B6:7[;3g7BHHQIH.TS&(]MX&UC:8SMe.3U+.]
V]&@?E5N0H@(W2Igf&HO9BS\g-6:R<O4\P-@-MUA45PK011Z@c2@E&EILNBW0EY3
aT.]=RVPV<(53/&b,DS\UO,&;Z+M_YW;AAc7)ZXcM.E4D&7+PF[JC]7OGK15e48T
#4fd4Z+F.#\H@H-RFbKKfJ\C\A01)PT8R@@2V9fJD^5QU<YUB\(P1G17LS[cfISM
HUBEdeFV75[BUN[V?/S=9_);.e:W^?cCQS:G-g,TFC,7Yd;e<GPN^\8MgQbb-cJB
e]d&J<2K7[B#)KA?SH,YT90H2fV\8f:aLf&-EM^8LBM6YNg30A#9]QF5g=g=eeR>
7UK-6\32](W)QYHR/\.B?_TXP/fe-c77-6cY&+:)ZH,Ze?)&;)0D:e_S@C1:fb&d
OB2>9S&,^f,aFGYUfVIT:IOAJ4>=6d4#a]]Z5<a[,d@BWdac=G@@,98750H8B[)U
W/c_?O,N\-5]dI[eYN[7Y<K6f,a=H7C1TaN>K6gZLaPbWW9][g+5BKee50d]cQ>S
YGN#=f==22)SRF^=9aZbF,bZH3:]bVF[REZ[LD+[1-PMWEFWF<>,_5OLd35/gVK4
Vd-fUWF81?F6dT?[]e1JI5&7?21_#Y\AC#E12,?F1_+gRIY)@YP4?8c:BZ9=/\@N
[f<=WT06bS1CS)WN<+Bd5S99gPGLGA+KV17UEWE#YC,@HeU:FE[IE[c4O\F8IF#-
)eV19-48A@9#>YDRL9X:g4O\0SZeGDRS4K9^=T^EgY3)<:3<L>1G4_@\UB_:FH0g
6J(R__#/T8ddSO6a[G&A\-,AXGN.Q<UXQ5=F&TM4@<-<Z-?Ha;AE/.Q+VTV@-X@?
2<AWMdbR6W&-]@_gaBf7./8E)XFHH\SQaPBYF?>8Nc)=bW@c:3Uaa;DfV13AZ8>/
X1Xg\3)25=X509C#,&aRE@5[++Z=ZM:RDP?S?R,A;4(A+08Qa6Lf,1fHDO59\g2=
,7;]JMdZ_Z+fM=8)fJZ&XQVPg?J#71VD7ac5^C&;ZY^H1d6>\@_0JZHfI_E44N8#
SX7?dRN4b?c^5263?Y:/?bR:0RJgT&6VK([5?[KXb]Af]5dTJMb5VKVOJ+71A9b:
FQ8,RJEd6CYRB,K.L8E7E_)2F=N/M?J:GI+.Y/,5RR_;0Q1T[1#AJ/IQ76NVM,<9
gVP5>9.T5LP<(d@.Ic+<YBQg0^9M@7BS2cE(g+a09cFFdcVN;U2L]Y)?f#[#A1<4
T.K&/Z30-LQX3c#V)=R,9)0eU(dDK=[64-eSDQB7<=U,=47eA<Kb8#NJ]bG=@f&E
\SU7bT?YMHR4c;K(G_]1Mg8RC1-IgR7T&LJ^>AI2W<H/S?[ZGG7U.A7)4_,<E\T]
.K/NTU93O7Q#IAWa\@G\1[<.+<d#g]_Zef>,>8ULRC#Y;S>YgRVae&8T&T=I]+K2
X1.<M:DXTLUFO=e/FaP37V.QdPb[F\KLMA)=3B>B53bZOc.b?FI6W5]a\XTYU)]C
SD8&aW,<R>::E_[F?R3GLA5)QU\Y4>^.XeEJP<R8]gDRAH.G]YHcRE9R(c3d^I5]
E4b00D9:87YUD_UAQ/QMMbE35+G(Vg@Q;Z4(,[4O[;R0A?<+.<I4:MJ8J_F-;b4a
^^ag8[d7Cf66dZMW]FQ.AdC;]@?_QJVI?1DVT9E4W9-fN1ZS?\?-9CC>^eI)aW2Z
3&J5R\BYD)3K+.795O_1DO2SILN_W\>DF1B\:P22DG?[dSdP)1JT3Q2A(G2NaOGX
6K/CKaR#<H/GOE@1>(Q/aIG;Q[S4)c/#?_T1LFS7>+0dZB8+KVd:B:IS3(Lc)Ta0
ZVPaCIg?=71_IAZ?5c=G(QBE01H]\)3Lc\ZA?bM:Bd(a9.?=[JW_6Cb?Z,1RYQ\-
Icb41<CD18e<VGA9e?4d3YZ4+&Q06OJA7ZW[2)S=)=SFFa7?Kg9#&Q@4Y8G+dgN[
2](_@7#7b>._C/-+]:/&1DOc7\GgXU3HP1HXJdR(Q(cVGSG<M<2#1&e]F-^5,g[M
4SaZ2^5V\GFZ>g&T@S[CdK@QJ+V(IPP0:PIVLIL7cG#ZSF,FLIc]+-=^G;9[1/Y)
D@SZPW\@d:JdJ5S,5;McP.JP8?A\09g_KMA/5N(OaQK<_IU/T6JbgG+QH1UUE<7Z
M(Ua8+g_WSH?LX(_]@ZDL+MdWEbIg?0GD\?d)2J.^Ec..Q)VK72Z4#-7)J=@OR+R
=VWS:>P#W3AKg.XN&Td/W];QZb&T-NNX3])V5G@A.c?dEP/Z/^CS+[g<g7f\G<7:
/[9E/QJ8g3,<BVKe[C.+\RML\5f-5H[5<?B-NBD@D#AGXO<2(&1_?.X)&7-@Z>)d
:AAWQb:-G^6FG#TO8R2N(T3T=TJC[c##PYg4aS:O#]d81+:Y(ceL&MfMI(7Mgf)@
aZMJB./64&?&F3C=MXcE(>A=:>G:&aL1&=aCBG4Lf_/>1B5bHMKIbZ9E/Ye0QZRG
A;N+g0-:?=SF5-1+:O00HKC5b)/&SEUMT?8NW\<FUF1L8=eP(d\0P?J6K_CWHK1.
Y,3Y5^ZQ[R((,ZB(@5DX2,YW^D<5YX(W>;6JfP07]N;/3O,@/Nfe#bI1&@4c4<YJ
]9SE#@IZ9H#/QVe6<?5S/N,bSP60g7Z4XUOYA?[aIU\O)g)+IH1QP4DDW[=BcM_V
D<BE+<<5P@USD,dT<O^0:W?<&4Ka/ZVC5.<GKM_G=ObI1.H26[XQXM1:TZN7JgD<
e[OY6?GVcA&5^Yc1>c=-\.:W,ReSDI@2PW-N^4RAXZHA^HB#?\6ZYR_d)R3KYaGf
=[M0FXc<=&79E8AKG(Rb\A&WEg4gW@D2]I[Ff4NZ&K&9W^B_E;39_9Wed15AP5/V
]P.P6Ib5.1<03?a6-I:F@?;AUb_\,;,-CK.D/^#XeE(bJ,[ZF7#70KEZ96:KIX0;
P7.2DUX0LQSg(K0O>3;D@aK<N0A2/E@Y[\KReAJGB7N-TA-CIHZ+31&7:=G4/50Q
X=HLCEd,<F@TZa6DJI]1Ag1=BXB-_;a7]DaG42KU+_1;d-R==(b-4A53YHD?6ND^
B#:UZCW(\7RHfG@G<D-[F:(@,VUXK<a8S)MGUY19]gTRYHY]693PcF\86..BV;<<
8S+U+Y,<[e)X]a>3L5#HK3c((Ed,4@TR4?6QGQBREP;R08JI[+C6(B28g27X[1HR
X<:7A7](YZYUgLJa_MESFP,QdP-KC4M\)b@G#U,<DAWW6;O5VSQY,a->\80)@T=K
[N5bK?A>FX.R3.gL0<Ob+4SMU>UF1YI?H#@TBMTd4ZMW++.ZRN<CDX=5DK.O\712
6XAUZHX:Mc-1L+5B85;99PXC;=F..FY&S)W:P,>5Q5a)E8#Y\N/aE@;L^@c]5E9=
GF9)U)L/HFVgRFNGaZ6.f^<E8WYQ13Ie#4UD)dB[<>&J;TPZD@Vb8gJ27/>Y&D1d
TF+Id/YCIUE_XQ8a^XHBF4;+-d=0BAT=[_9;I3B.^@P[Pf:I)M/f6+0N?;2Aa64X
16SN@.Vff7df4^/7LL/XR5f5:?IAW@VKW.B&CPF^-F+VN#28LbK2J#BJ([T1KGA#
64D?Ue^BPf2>=@A6B0>/LfPaUV=)++IgJYTP62-X<=cD#<,^97b-Y9=-dfCUZ0\O
1Ef47fU0?AT#H=5GbK1V#5B^Nb;_R\T)>B[AX.eLc0DLOU)Z_K7[+d^>3P-M2ZT\
/a9E.aZ1R/87O2bW5(D(W(e(,P_)DH1R7>80V(QR^,d7;OfgG:WZAR99NQ)U-T#1
IeYVA?JB8T4V^1=@RIbfS=]@+<9F8NI6@e\:(A==g;;D652AZU<C9UYJJTAdZS+?
ZBOdAA,cgTd,bB6eS?D&V3)5H-W#?CR)g5gOD+#7,Sb-VZ<\J@0E[/KT3bM3L6Z^
(R8JD03g>\9fQ9DM/WXeeB\S)a]QU<;cEe6SZeR)\IZO_28TG5#GHE([M3PAJK2]
)]A4SG0Ba9Kb.96634[UG,D\/f&]^QEIQ^FdLRVW[@@=3(?.E+(;X[[W6_RP93^@
U?,5gF=)#74B+IDVYd(D]/\I8WX=W;UG[;)/,V.c5eS8I9XdfN7C+.^)-&E6A8NS
NBN@&CAOSAGNG\I0;6a-X&A:8V\BbTAQUZ#>1PQc77(KQOK#?6a\#J78\8JQ,ZPN
3@O)e9LJ>I8a4L6L)0HER4X#[KIW_?gJBKN3L]-A;0E2e,[X6VD#/bgVbPXFTBb-
((#YM>AEHP](?cWJXR3ZC1011TY?d[&+cMFQbYbPU1G,4Q0&KLfTFg?b;14),GX2
]Zf0.F/<K.4.S=X\NJ=ZC&IT\O]IB4C+W7(&c^;0caY/X]NF(HQ6:@CGKaA_K]b>
(MR9e>bKf,;_CE1QNP;H[<BMVcTZg[V596V^eSEQYR,A70#Q3I1Y#O/Lf_H]..?;
J??#3?IJ^]DcT.<OS>-GC.Fg14F@>Q^7?Nbe+;[+7_QaS]LdMDI.0W.&@22dV4@R
+LEXH7<c[0_e>[L.C#QIcG0Wg<M_J>--?aLd+D9(@HAQC2Y_IYd\(W,+PgED.S\S
RL8JO\YJD->5?-K)U&CQ?BRM+K)/1/C+H(-NW7IG(L?+H<bMQOR1J,Z9P1Ac]<,?
B#-Lf:f&K-gd@W<&)(04]I^>T?FJ6GcGX65MZ;P9+e4G]74W_ED.)<]95;8K^bga
C:;/Z9,)>ODJ#MNP+R7<[L8A\Gb0Y959GAI<)KCHgH-aQ]^Z<1V7=C.Zf_4ScCKe
-9FV^f<<Pe4\aZ;dQMG7BN?SB+^HWH+#<SJReM#+BFRA^1JZYF6N64cYYH?ZJ==M
Lg\RT0fL;EO<<C#R+U\S7?H^([>8W#@<a:IND48:0E#AZ?Wa@1NB7d?]#g/Mb1XE
:FSI3TS#5>L.<WPIF)&:8,+0>L;#DOPCb)&DW</,?;.T@?bW?g3>YI0e;ZN;3]T.
#54.J9:P2__F]5e/R8Df(e8>1?HbLFX:QOB0=>S1O@+QaPP.(21;dV;e]\U^P#4P
cHd@6W-LQTCWFL1I/M.S;U,bf,7.U0Q6])T9@\g&X:eQ/F5a6).GJU,XFg(CC=V1
>-,MFD63;0DF@EZDVef]Td>Z:?Wg21Q4Ib<-609C8gR-=Kf57EUGCES(1[G):O(9
WXF@?_cad.8-eG;Z-Z3PdN.dT./0U:X1279K?/OKAATaX?f;&7(X(YRS5Y@(QZ@-
961;d-D7SGgSeIeJF3?XT9MP4B,QW^1PK\39CU<a2GC>b;a1.Wb9G8caI299f&b9
I)M2&e-cNOI@g_@V,Ib-O/dQ#PX7;E/D_,JcY?gW?13f8V<J.O6V7MLOI=NO<,dR
M#f&@F/[TfF;^Te7XWYDC=Q]:B\d8eGAF)4YT+/).,;5]2?Q_>28,aRBaKR5C:cb
=OSR35,PXD36XC^CPbKeLUb8Z(\1SAQ,5>J.8IcaT]1gV)C,Y5@_5HZ7V:dMR^eP
cgbA\G^<?<UGe39R[E8PY-REZ7(K7BGA]_8+:\V>,EbO1e:JL^^\5aCJ<2L2BUHT
W0,:P>Hg6UcLO=DY\ZG(e[UWJRL_Jfb[(+W,I;0:^2X_.^=1NVRV\5bHDM40M1\c
gHdeK8X?//@0^O()Y=:H9V[K>;1JA&=SJXB]DZd[F7/2]Oc[5UA[eO(.QT6J7:[J
C3).TH4=dHWWEG:9#F5c_AI-R4Aa&?+IDLB1Xa@H912_-_#(FDJ\60a5H(T7(PW4
KcWPe9df@ffM?cS4;b4U[b)U8<_O,#FEZcJ)&<5CY8Pd,7O@d&[fRV<JGR_BP/99
2A:OCS?3X9^HbO0_9X36)&U^.#Ma@3f2(f774f/(+BF3+U[E_baQc>(bJc,O:P.6
EOC\.BT5RV[fX/5d&f1dU^NDXRFP:V#O3LLYF2O;,3VQ7=J1fHC^_8M0U;YNZVLQ
R(F=QHg&K]gO>)<;[,We&,4468MAGT2&7TBXOD&XP.3QDR&EX6K@JWUW2PG(LQEb
Sa+YVB)Kd[X/CJ.;3Z9W)M)8D?E:Z.bEdOS/PPMJf_ZXLIS=V[d,[]M9Vd>]L6_:
1Y>c2gFBOK;?<UZ,_?3gSeYQcaZR)g>UUcQE?EQVg_X@V8BO=LR9URW8fRW1VD_Y
S&)RQ<TO+f\T#/KJBW);K1g,e,T1OWG@U:gE;WF4WYEY9X-][;8Mb]T?]XV)O<PZ
^V^5;5=Pg&UIA)c92V0;BT?AC[\JPFf?&Kf;XPCMW0&-[UbJYec<])YH7YPed([&
L6I@fC4<BOZ71@^(#C3/MH?@gW?\I1^H\eII@bP-->ZHK8NQDW&7-Lab^R66I6(S
d1,IHZT134)U?Q=bU&MA((,R_IP?WSRBUNY\SQ4OBU+C^5g8?1YH:/^.+P=^Q2H3
)WZP?&W\[MD/[&DW>HXWT#dGa#UN@YKXbXF6Cg_c1eT=#O(D2cW7P:HfUX)Ye:>E
8+?T?.Kc-?1IEPgX7QSK#3+35.UQ0BJB-Y5NL1[+IAV]baQ>cWF54)Y>>ZgdM#3a
XZKR\@BDfOP@(;SMf#g=8:/XGC8e9_)DEdNQ9d]PTG)=ZfdJWQ=/b,0]NeS@7LME
NAWT._SVZ?WVZe8=\\fCAMDBA^F3a/cA<1>29DeVcWTZXX9-U<9/;])bHcYcL<JF
,g=D=^#30W,PP1-egRE(F>M#4Yf#K?fD2R7:eTB;Yd](?6A(Ua(;eRA^#Z#I,a-0
\Q3gBO0_(V^d=9&PeJ[1@b?C<8?+_95(3N(QC+DXCbXTIC/?]08;/NBK[WCd=:g#
RfNeAO+0RILDAKWdIQg[D==)g.1g=1F\)[W2AZXSH?.\aT#_=R(a1D-:[@NP@UM=
L)SX^SV4V)5d6];](fNCLX6;BQ(E0U6[AVM6^7FedbbMf-?#(WR5L,7_WQ(F#[H]
^O#WcdPXY9;7E^&->>T1VXJ^>fgL.D,bD@4^PVbN^6SH6W/.Q<U6=A;eGM(Hb-E4
V2][6VI&[EF0CCWJ1,),d?O910?3^8f\^A&XWbZ8R2?#Rc>O0_;BKV6LG;)ZOGf9
,6\eJE-EW)GC[#UGZb>XaZaa&7PC>48MV16?9(>4c<A>Y(S<<^\7[2[cR]E0+44M
Y[2KA>:-8DB2YaK+<QND61\;FJ).59555+H<NFZGg/#W-06MFgTZPB=04a1Ve4LP
1=OENdS0</aO1dPW^?S@?Q;^53cYE/(D=T6TZMA#)29OY(5VT_^9Dbd/RV<\\BK3
^>b]Lf2MVdC\=-6E@++YVE#T&\L&),)R,bd(@NFCUB6K(2_g/QH0BE<<-QT;7-bB
aP#g2F30A#3V:DC[,IfXEaSPF\NAAHVbJ?TO.e]([6XcOT][1WNIG-#2HN8VAZ3Y
<0,/^YS9@WZAG7LO24:[D<g0>O2JQ3CC3OH5gOSW-dAYPF\a/)L+ZBM8M8Ba>AA2
ZD#O8;&:DZ9O43e1OP59O1#OY.6f8f54EV+L2YJH?E&TIVAC<aLNd>_./IR+PRg/
W9QeY\e;S5PANg;^G5N0.5]US6>2fd1e:]_Y,GbIK(:^^FZB^:[/@SOG,b9&Q&4?
AILSLUB>Yd(e,WQ&UUC3CAYD):;^H7(Z38V>0M_aE+]d+\[B5)cMa[2;_-)HY^A&
<:@<2UM<RUM0P5C<g2-+c@TQ=g,>(^.UNZa6LUa+(-Z/X8fbI][bTd]\9)2>=8=3
I_Y?a)2)@+Rf&_5[d_(K/&O0HQ=E/2cAeE_;9&O;Af+SUO@<Z]AQ4J#aM6>?-LZ/
=E7H@<cfd)R8NMME=:+U=fU.]WQ#&0S0X=4\A.ETZ<8>Xg<;AY3dAcHDKV&?JE1U
4c1?c[:_]9#^0cC]JDeZ/g/Vb5gT]P3GI:37b?ZR;U;./M1d9,a:(TDKHXZ4<#<]
3.HJc8eaTcc?P7FJZCd>XgS4;0OgH,ge6<_J\+UM+A:7:+75A2c(Y@<a=W4Q/AW0
<F2d6Y^Eg9ZSaQTHIA\Ed)gG^>E.PQ(=USWg6K_-6a@dTC=[)JR+UOF<VLE9caHQ
[=HUf:U_.FB)JP]g)O\SN?Y07EIXdU:,9S)KC0_YL(<><2=dZYWQZ><,]H8^b3L/
5\FMdFBSI><bOa>@.5?<F<TQa/^B5LbM6GCG?P=4-@#GVfOW:>[cCSe>=X97,4WI
G@.Qc4Z<7Xa?DR/:O2G6S3V)]O]8TB_(ea:NK7J3_c?5TFBX.GP:W-78,^FbUEdd
7E=0X(?W3,6;f);[&6.11^Fbe+&&<>b&Q]@.&P&QTSKJ/1QBf(g#321]D1[e1?B0
QIb(/,X=VG;G/_-[YCALWXPC1;1WJ@ZEFSK_YW_>AFD0MY-U>R1QT)[;FLC^EF@?
b174]gT2JbPQ(S+#aRB;DVcV_/(R;K,BD6@?2-UUG\H]IN>ec3&5D?a_Ag[6&-(X
/:7-=#S14558BMZb]aa=MFaTX@X3=D7S<+>WDYH=&V#[OIZ4OSJ1.@3.]&c@b1YO
LA.@gf8]07Q2N:>VAMGBO4-BN?5YFE+<g4HXEP(5e^4JG9[Ld0AeOW1XB)Ba,NVW
S,9(e6bM_8a2+U_@bVd36XH_Y;<=1<;KMM<RS:7ZA9H/V((7DfCCADTG^T9HX0d2
#=Ca.dY+M_QR-ZVV-L--VREaJTAMD1AG]AAMc_SS@D<?/[G#4G6(W=Xa:WCZZE8T
PG<20eWEH[8SQf(,A<HCF@IZL#f\QY/HQZf?,1\\=TN#8(;Le4/X,#\G;C+IfGT:
AH.1MAed\O+XH8(,-T\<94,-VOa+a-<?;^IaD(R-0GFPfS-faEc6QLU@?\/S:ETB
?:f>_O-eCDN;]5,5HGZO9a>(LXJ]\,5BV,4OeO=_J<G.DTXJR\791TTG=C=&C,>0
X2R:B@[ODG6e4:__ZRC+IdG43HPC7B6DIgRYFf_.LFdOLJH/dD=CWV6F\dG+5H1)
V[43()^UXM+G/R47gb48-MKf\_-DH^C\<HRYa]1d>2Z_7=>_EJ+W\)Y@FHG_AIDF
(\/Y49[1MD(;#UP-7S.#&+Ff[]7IU\d463:W?ZNFB1XCNR.4G&+8599.acI.>3VD
N2]8265ZP=f2;]<=gX\[KLDeY?1DT5M;S4FB.\@8;RYfZCRX;fZX<X/EL_/(VP90
2aA@]Kf<XW=3c@),f)4>9@7&1O+E3,6C69BC=0c5NP(.CfKb]/\<):0JUf5=DV]3
g992[O]M\^.I>50Ycf6b-X15><]<UQMd20DI/[#J3g=:P[.AUG+&g=dR@4K:#7F;
0FU\XCQBdE[F^)gJOY-NCJJVI\/EM,@d.#K]\cFMCDc35:?W-_d(<^_F0\N0CQ-8
/<-Kd>[bRa@WCac][H887e4@8_TX4296QTT/a+0LJM_HgEaH8MRFS,GE--cVP8KQ
4(1X\@9R.1UMYge-F9K3YbWGDH:-_3EXL<GY/eg#cd;#0=?X54A3E^:Y\>^I+Y.^
K.4JVC1\:QPa<Y^LW(I@])E2WZ)D(CUZgVL=6H9feC;./G\]+a8Q1-4DJCG0D-D8
2&<LN@(6Jg^#IL[5Z<UG_[4dGA7AQY3>^_L+KVf#3@U2RRfBQb2F.FUUZ=CJFF?9
,JW9cCX]e5.e:F]UXLVZa@-#Wb.<E6eH6QbbQb#Oc0&0Nb?Gc/VO?R31A,\0ab>6
T&F+Z7BCg8-HF)=C.:9P&N@+PI[N_;:ea_)0IVMf@,X<;EBcNa30,(K04g>59]OE
ZO<+cS(;.EJS3U_9\W4/eOK02Bc<XgaND^X/a9&>(GRZUY[aNND.[>R#W^^2f.D1
^>;L^Ha&4JOg43KGSCfKQU,VXbb2A\3(E8@.6RY,B^=I5T3]STA]VO_0XeIOQ,S#
CM0fE,H2^3DR@UH]HWVO5eL<:;)2NfSYW)\cV+EGPH3(MTRefOFLKfS3Q@aIRAEA
Z,-Q?74?WZ]#H3,H=^D)M-MLD7B]^^ORH6Sf\[ZS\=gM01B=\:dHL\IBT8PD3)+I
N61_OgP5UC3P>)b/V,Pc#T96K0JfTF;e_WOFAI/6CYC^Q<_:1gWM=@3)I&SHC9./
+aKH/.?X\L=F21#39?bc[@13:Da29.GL.NC^dDdL@/V=e#e@f-I<3+Z1UEQ<JC-<
GIR#bHNSK)@]R-K8eTLe(F9=QY[PeU4BAf7?1;NV<9HA<-aU]Y:8B:@[^5+,K1S+
YU:?NT[#PQ>2ff[+YK1OL49;N]8UWeWJUW=K>;<>S;]0=B(VFaA5:835VUVA^e61
V>Z/)W6KHH^8X>MGRa&QYKf(FYVW47OU?b=(><\DAVgZecYWW+Z5DAc9gR]B5VM6
;fI?7]E.+2b(3f.I6\FK4;VcKZFGY_YX=QcG=V(dL6(/5&e4MN7-N?&DaXe=D#2C
IfgJ?KT\\YA,^4EfV,5U_aaOT^fK6_Z/Rc^gSe_A,.;R<B9<K##Q9#4\dVWSSQU=
G5J_JA[XY6JW2IZA#OGCO(IRf?dWI>9G]]K;@N\DV0(C0E03(:BM??fNL4SUMM><
,+_C)<?Z@dVV)7[aOY1?P_>20;ECZB_Pa;M1b,OW#Cab@\Xd.O(;RA^16^DY>/a@
:3RD_4dfZI(TaYG81_J\NSI8S\X@&IQ,F7)BAM#(8.]0;e9U78=UZ=R58eFC#^g2
,G6)#);7.O3WaU5(@@cd9J7Ab(WRI?72D>=7P4R];T,8/Uc4ZbF#2,,KHOLPVL)Y
<^O.-)(bCE/ON(L3_=84OPTIA\3HZX9S2L3COgIIE-XD1-H>3BcdHCRZQZ,V/._7
P<R3RDU#KfFY3N&<FVLKdI>5gCH/BWQP79<0a3BJ4621\c4)A(+[ae&JTW=^@M)A
F_R#K&3^M\+C<eBeVZDagV,Xa\2>WH_ZB8-f(dTGBV>1gDc7b8V0CG>\N8ePG?BK
EfcQ&M8A1Ud_<>XFJJHF-PU+e;fHHM72&??)Q)9><)U5KU:dSSc.ZG/=(O63HCU7
^SV0[RLI4_\TLS3,3Y@0[GP32,dU(R=EZ>D1LP2A95TGOOCB=V=)-^0E][8fPeXN
F,SK<.REQ_#e7&=7L^9I71IZ\<F:]ET4_4WHgcG=2b>6ODK)C1/_9g\AF(g:@DXb
gFY-b0>]K.B:=HYX(bU3=7d3L?H2_>P@8e.fHG3;O+J+/O4c:(C;bc-_.cdCB>34
]bO[.1/2L]F?F;@1#GbL7=4+D=T+V]=.2M4GGI7526A.1dODCR,60NI#GZd3&BDZ
E8<E26U-6]T9H(CYTOXFXE<<#9RX83O^IGdadX];NW+GJ6.,##c0C_X8UX(B[B:.
9603M6ca(;=Je=:7I36X@6/5UPRR1;5@L87,85bUZaM12P#M57DK,\IL6M2>Zd);
A\20<4;>IaILBLf)0Z^.E@_O4\4bBE5JZ&?0a4Sd3R/C1J0:SQ=9Rg+e7KRWFDX&
E5\:[#+79&L5R-f0=&124Sc(9VGeH49U?U=BcUNR9JS\S<^d\L5c/Q@fAb<KK#Q?
;,\GQ7f>D,#RJF0gTAec_bLd1P4T;M7YBW/1#aS0?gee6)WL2d(4eAW;afGcc0]f
4R6Je]W=^9T0_f\)a3KZ,F@D\AKEaKLMG52)3E9fb3[O_^cd)c6__>[TQI5dcVgB
LF+4RJ,??+PUCG/)Ia:32^f\=U+c4ObJK2_4RKge9E>Fe_Ld.cBJ&-5IeTMMe3)(
8V7TQN+BgWZ_7d6D[E.;<1UaOWT9=8(>c09R[<Za<UN7bGJdYB25:GW0gbPN<G0a
1OF_BRJ^:E\FPST,)PI^X755Ca)6EQIDRHT[g?K7865Z@R5G;IMgW6+)1+fd@TK=
H@(Yd_e.]\E;TYQbGeBA@9De\PW;<NQ8H]_C]G3#VN.)2-ecYb7;9RTF-#SDD(6Z
OR&WV.9(Jb0;HcV0^eJb)(3+\gR^Pd,](GTbE??f:8JN>;V04,THe+)aFA0]2LIS
VD15;3I^e/9B+?JYaUc,gDNQL_T.Je4gNU@L<P35fA\CCV\):K9GfS@eQa2@,EPR
51=1dNWBSeRFDPXMV?#)USED/;7(,6EY5+R3K1NHCPXTB=;M&eO,cW3FY^35QE:H
5g>+N\P?Xff4CeN8<BDZ-##I4/0^<\&51QZLDE(+BR@(O.4U[ZeaD_GEZU/7gGKF
YR-f9JI8ZCg)E(;HB+=C/S=3?bL\UKTeDDOSAT&aS&dVaJ@,4&6M3-R(1.6U+FZM
M.7S#\A26=U[DU?YL&/<F[aDK5#7;MD&]\DQ^A@.HE4c4U>+?:VG^X1CXgHIEH\2
[b^-0>E,-WJ;OI@,U)eFCa,,B)?9RIgW[;VMM&.W:/a5P^\;JSR.6&]9DR+OAbW4
ST21V.8b;.F.ZePe-1E>Sf_V->]EO9#R1_eR?;B#QADRcJCS#8gK2;>.KEfVg]K<
g,_3e:SQ-bD;H@eI3V4^F3)MO7PgE^C#HFU6C;]KGRYVQ_a/B/+ce2GQEA0c_eBL
Z]FHP2+R:UU@&?XLKX@R_4g<RbX7C6Sg08:IWS[Bf<##^T8&6D\W53)P/O[KC+@K
E_MR=bD-.1F3@V32/Z40/<>G2_H<YF(B0=;:TL>;9Rf@B.bCT)DV]S3QR+8eQ=O2
[4&&E;0Ab)5?W/:F,T-3\QSGbY(c7:4.]gDR>AJ,W7b=&?TP/^CU_K,[;&EV)Bda
6OA/TZ=FC)5U^)&VG\d9dVQD@\QO-=Pc5>Q01T]18()-\W.P_D<ZLaKa\._6c733
=PYQUe\KW;5I#W_>VB1?P?+g+W+06&geVYC8)K6(HSe+ZC9ZaSPIPb7_A97fg(6+
;#SDC0(H/H8+I>(&]9:gJ9>QGD-DE-30CX.ETPbDM[JU^65QK8Ba^Y:ILZW4c2Q_
,QAP4G5SSJK@Q^f]OeGF<5CC.WQ_-dVU8dH>64)02X6Z@Ya,ORJU/F[cGL@NM40L
?29(+GI[Ja_)d@8gceE]V;HZEO>?Wf.DeY,cP;O-I@,<c>,A^b^7M474U4,AHD0-
Y]9EL0&/<aUZ-3)D=:cWbb-7Me0AAR):TEF&Q(>K2[,Y_7/c(^W=aEZ_]ST1=NMV
WGJM,f2LMa6HY;D>8U_#H5:^ETL7eTOZ&dD5E,H4O>EO267EE3T<+b?L;BMUcZ/9
<2)D5;M)J@/)(5Pa&(e#MZGQN,:c229UMF9,;fCdQR4a:.##/KM+=bX?3/=EKKN@
@&6HD_I8@c03TIJ3S3K4;cV8LW(>adY1PBaIe;#PG^;BNB>I_[.61IM5CK<I3>?M
?J>FUIB]W+;;(&8RPe@Jg9f[,,8M7<K;FO2K)L[8_1cWKJVUFL@=.X7R7/#CG<9A
UOT0e/+3O]KE,FA_TSg2_XfR^#<>\X;6P<)I&gLbY[\R3Y^1g#XX2,?68:QRJ@9d
6Z3+g=7G]:+>Y]RP.\ZOD&/UZ<;&>YW2PRSRVaf5>L#VG)8)N=1(-(9D/,FS(KL@
OXdQH2T@L9_IU4)[&S:6SeI:52]Pa<M&R3@NdA57GY_GdXb4RaWVEBTK+7Od9C)9
bD-[fcP>P_6>;],20<=^=CB+_V^K<5].D6Z5T,R?=8:R-K=E8JcI=F8,N_K(HL=9
-,f)[G^JIB+0_-L5;&5dX[NK8<g4;\])(2PFRB>@;&@g-KC^=g5>b5_=N)LEKPgg
;b77CZ>7=M/b@1fEeCbMJAZ821J;d)DU;?K3baD]^[ZC02<f^L[VaeA\HeF8gPF/
WcR@T#_G1Y;N\RP&Z[L>gM:^GA-A^e#>]B8^;B7[>fG\,&JWMeeJW6XTATT<.V5[
SC>C)c1Y@:Z@[WBad/eTgeADG&A^;RfgR_?>:-8NU.d])Y7^?:Y^.U5JEN=]S-#2
:/&.@RC\1TY(a7=CRQJ2_S.,522&N)-D\8;+K[#UKIC)8I:fV.Z#66N426IBBJNe
#/KA>FYM]]_2?RJ1Ud<VQ\X30@RO>@I+H=ZNC.&H[gUb&#:\9&WGFG9LHd9GD3L.
2K==,^=C,A.a?;4;f;3>XJL4..=@4dc3fFZ7Ue9N1@8^WaTDBfe7ENS_GeD>V#KS
UE+/O/V&eQP.M#WefA@T^)BI788;KQcKCH9H5)5MQONcKGCd_7>P?/CCUL8&YB/L
,<N)MbP2+]:4)J(06CLA^D[g2ZG-Z]gP-7ZQA@I]?=H+E)C&W=ZQV):J?670AI-T
3;PXdG+9X/g1#<@QMYV8()bX;eJdCXAG?3NTXU:@R^]#AMffV7aQA^@EN1f+XP6@
gF566?6PgD@AVUKCd-faA.-P1(;O/P=U,A[8.Ye_VKH:+LJRXJ&)0/:9W#(Yg5_f
4WHK,;eQ4YME521SYJ1DE7eRg\fG@G3eD=eUN5Q8#[/cFF=bg<bB,BHFU(-FaND,
-R0B;E-J4>eF;VOQcaQc45PW:FV<^=aKR=g:cJaKFQQ7-A7_HR1#c^g0^+]](FM_
P:M2T2X\KBb<bK4N9C?IgE]1<N26WfIYHC^&+<,K1O1U5fc3[Q>/P::#.[;F_U8L
N.>R-I(#5f-C2>?8X(>2S0#92AIO(XAVf<-@5-fRAd4Y114_Y[&fWD-Db:Ec3:&)
Qd70#P:Y)=A6OR;B_S&B,(R_]\IT3:8TU3/IfbZ6_\RK>Z57C65gWd)FJ][9aJ;K
&I<\;;U@;3()F^gZA[K]ZEY2_gG.7ZBU)TJ6TO[d[L<@Q)g4?/4UMbAVOaf_D=g[
68)2-.2HCMFT;5F(A::[P57:dLZXAe:F&d?4WL#JCZ+WaaGH?RT75W;DE,0D.bE3
_CWJD4I^B<V&@3,BgVO63_2bJSISY.@G-&B&HXe()85bb&)\@[A:_>CS6T.V16>C
T?ZfLaHBJV70c?V>9M18bFZgO[L^#B<+.f)=2bO#3-1U0QM,AVP\dZU_#^,S#F+.
065TF.L-)RVYESe;9ENFFYP@>ePb-HRYDRIg^aVGf4<ZQaD9#<<b2LBW\>T=NRg)
NE7.0,ZH\RQW?+HACCC&P2#=ff&EcVUaVf5@&4_4=O=CD+DJ;7Y]RXZ;,5ScN@VD
RfRHEO@4RO3BFb:VY?&#NVFbF\K79I#U><c=b#eQ]1Z?@e1_@(A=4.LO)X00]H:f
QUAE]9a2SQNJ9;WdD0Qd6BV<JXe5X+#:d=;GCTUHZUG2_J7<@S-(#I]bO6SPG.#)
1e.>ZFDY5#P^(Z+a=Qd-AU8E)0JYWEb)OVKKVC)Ea06,He1fU27?1/6(F?(=eF)J
:aN?D(N(WbKDF6eAI4XAA_M;QE&/N8G)aK>g4d>FfM+WXX[H[L0c67>C7H.P=KIf
>F:)5<T=/LfD7EB0=[Z[3\&<0>]6R,^]YGU9,ZX8(+F+QgPL:2M0aO;2b=U[M2PY
T7Ye.-cC79V+BC6acRFTO<eI5Ac?7OEb+&#)6M_Z/.c@\@5]>4:I?]aA@=bcEbI1
J+?;ODTAL6ggH#.KRJgcJ9]BY^?8#(I[b0FgbX2@H?Bf;RV36F^b-30AGLDRf>6b
@OUgNe)#:&F\Y;-0]f?_e+),/eY-;EN,_^?,?2CRJE]MJV,(DP2QY236H?LSR9(S
OUEDa+_(H)^1\^,VC:?JUfHdKBf)2GTB]W]@\S[)1?H4@G^:KZ]bbS4V]C<eEJ=.
LJ^BI5+3]WB2XH)JUM8<1^D^aT#GA3R)ee_N28gDU#d,8?fQfDMa9IM\R7YcHZd&
U\fI;_E2&N-1M73Z20]fNBZba?Q=,TG?D/5/=aacP-B#\8TA[[/-fXGK21,=QN66
f@S9GaP,>P_DP3Va6cC9Hd/L<)&b]5\4&73Ra8NeMR_cdS+M>O.&>)TZ,O)d-+]:
ZaSAQ,C38EBGg/1SFE1J3DRQb5])>?ZBJW2CAD--@d;6/F2:NR:JXS2#dce^Db[Y
ce6cC#bd/d/=Tf1YBN<JEY?c;dT[/#)I\Ye@2Z@0AW^_[GP&K^c+AQPC@4-)W9JD
/F<f+Y]5/^DZWSXCf#4,81T6SIA9T36?^BbN/:[SeL>L8J5NH7/.5G-MX8U/VIVI
=BB;Y+U<M>b.ZaNY[MZ)<2Xf=8@MVdWJ@[0-_HBQ_C>;Y&Z/;P.JI2CIJJ7=&A0W
3,.f63CcZ@-0(@#W-,b/LT_ad:)MDDYS1f):^MK;.S;fgL::V,4,MLW>AVT3B+.O
R&,I5F:P&55+6Sf=0#g-YX#<W(c6+3gQ;5-P.GA0CWXc#IYOe2#9JKe=cPbSN_/8
fN.=995#L8/F69_5VYNTRKQJF58C#(=H7+6&bKT]Q1,3gA1&0]T5[cbDJRL(EU=N
,]AXCVS_GP[6f_1a5)9&_-NTXO<V+/LZ#;XcPDCGb7cg+>EX7<C.DeZ<I3RA/cd)
0[Mb5;M.H4ZW_ZcfZ]FE16FNLXW_JCIc=4+aL+aM\W[EeK@QRJAO7[57;WE,cO1Z
KRQJ4?XPK6AQ;b,gGYSB8@cPMJ.8.J^F6V@F0C0<U1aGG7#):Ybc39G8<JaDbb1I
bP:D=?bLQS=+?:ZU&#^.feS/(K1gJB;8gbTRE6KJOD??(=F(b?,&GLD4>PT]K<(f
;/S;)4[094OT5U=0:D<FRL9,2N;cc159YDEF^.5a7_,+D5X&RRAFPSC2EL8;UA<?
^dX3Y.bM:(Fe10@L8XZIBX><_gD;,Jf7:F.(X7eJU-eXJHD6f+,HN7ZEMd<:+>H?
Ma0DJ-OC&UY>&O\<4Y?bD6,R3XfK)?(f+K&0-A<YdMPg&CNGOR-@S^N>+fRC_F2_
L4S>DT.S(Uc@;De,aYAWf@D7HF9MF?W)ZBeK=Y_&Oc-)@_d[La7S/L5V5;#(=W=Q
YD;#2#6VBS6517f?POXUY0XJ=[A,)4-N_3@ZBgeJ,&?P:5NE.@+Nd?N0f47Qc5P+
45EY.5d:<(9-V78_N+F])e\.U.?BgS9N=gFJ);=Kcc,S9M4f]a8E6@<aF-H6<#=H
[A5AQXU]UFPeT1db#(<BR4G5WYT/EJ#.@d(S_K,ZF2+UEXM)WJ]J<CDHF6[.bCLc
cEF9WH0<b6&W4>B\.>E7gWH7],(.BG-HG@FaT.Nae9\#f&<_fD>YU51:eK>)]STe
P9Yd2[e,;LYf.O]LUc\Ib838A-8\7c[eD06/0da\#IDG@^,3:@7O_FFGf8+(4&5d
G4+XP^;,RIWf#J\?gFFTW=B;E(a\]dFX+)abH]P.R7BC?cdLX#K(2W;&WHV&36d4
2>[geGOCWR)S(&f)0RKL9MMC5/dE/N<+<WILg+Z[V6eJ[J_)(e>]+d^c_ZXbdO4-
=NBSD=TCfY\ICATOFJ7e-,PW.fWE4CBQR#^(3.PIN@@eJE];-4C;G)]L4RN-c-S/
UCY\R#UCMB<aLIJ0<Y?&N,RFS=+#e:US6gC]5TM6bJQY3&YV?W?]9dRCELaa+V<+
U(fdY))Q;Q0>.#BY/K@NFba6gUg#V5(e/bF1AHab\T.E3:a-@Kd[bW0.9T0V3J#C
DEQ6/2WUO_5_?ID8(R.__:;((+be7)2,_&Oc&;0D\(Y.bP[bQ2F94Ha8B(S7V?@d
0V:/fL43R)TW-6dgfgW-P7<QL.:/<J@AV8/f,AA\]T4]5:/fLU@SKLITc:_1FA=O
aW_08]d4FbaCJMS<+VA^M^H(J[cNG]^aA[Rg))9(NgNJ>N<d.9Of6P71CgN+<#&(
K2QH]gVVcPaV^1CGFELJM36_+3bfM>G,M]X=NOH@1\AM_.;3#K<WA:<5<Yc(7^G+
I@gD5Yd(0:4(=6\]^f+JaN.[IK6M,GH?[KK@#cS=2]IG&/#C4-B_aeX/dBP:e5/S
2.145YJgLKB/[2D#)3J;^bfUVCTU#8.8P[Q^7URSK#bcPQO7Eb-Q/FS?;@;EB9B:
eVG>eFb@N_[fQLK9>N.EQ?H6D,VO@/7=HKX^5@-gU<D/UZLD6M3L+RY?JZGY[#CB
e7<Me>T3S&fgF9L_UV7F@W1CKQQ@9bGB@Z9;74<=2\U+@4b8UO^<VNQc\M_U.BNa
>?VPAPgAE,8Yf73M)HEO8YBS;)Y0K\7dRMg#><aTE:/&LcP6#bg[D4Y>.LFJ;5&g
;AaVH//;a]RCgD?7Sc3EKHbV_.AJE@cF^+g=5dI;7)RT</IR+]-)Q/X5(VRR0;)6
6YLG<@OGe?5D7??Q&>/e:KLPQ:egdNQ[#@UR&YX:T:=6c]2e_8CSD>.8<Z9>CN&D
BSIgBN&G?:.bR?@a_(\A#Pbf@C?_QdKYf]]4)KcM0NV3Z9U)SMDa>g9?Z2IEO)+G
e0+aC4CO^=AVIKE]@[P?7N_<bW[/U/+Y];C0.0T<CXWN,@5F:QSYO_20XA,G(/<d
W>,_[Y9IR>8V+EEU;EE2ABYKV[c^7_c;a5<3F@^9_Sg:OGGdM?P_Lc]+R2P7B<W&
_9VbHC(Nd.Z^cLH+60e]+fc1Pc>(4&2A2XcJM1=8cJ;Q1T=f:3BX6H)B\]^WC^_H
)YE9Ecb\<B.,BP&aGg6UA:gC)/H4R?&&Z/M=[MABSJfO)aH7;]9=UcJSG@cLJJ#E
POWZ6]I:Z5S/0)^U4Ucg[a+]/?e4(QP7BVe.F)7_A88/:93TXG#.YB4gFUXOUSP,
N]XQb@fOf;S+&/VR?Z7S8<6CHNGSQ58:WM(e;LeYf+]0BC3(_C1S4R,Ja)\a&e;X
^<L?b=-)LT9]MVcCY.,\>-<7.e:G2adC@f+VTCL.^K\;395K.,a+bZL@Q?YQ5Z4a
A<c[11gY)9cKRWBW-_PLMWKLCD/PRQ/F/=QP>:.PZ?,MQ0Ce_-[0,]eFcF1a4>,e
:AR#dP^(8(1UW+PB86<L#F60.?IW;/gXP\XK@6KLAdF5e42\6Xa.7SH,V@?1]YQR
=63dKQ/+\BM#51PfD)e+_a:P5RN#_D_d(73c>EW=_-Z#<25L-9X@5Wf:GJVV0C1&
[Qc1#_7+6]-Y5OZ&)?J>R@d16W-S24,8>VBI\0?e+\EF+#]&^E)0,\;47D@)@B>g
9f6\VL,Zg;[#(FMK<fOIeQB83Z0gIY4=9[M,N:)=-d+X/JS\e0^KER[?W,7MC;eI
Tg>MB)b(/],2Z=H))33:A8SgggLW6DPZ<edXbI>gc=&Z4JRHT9U?[/US67JT,8.1
De>Y4<J<SB2^>0W?I7;;0U4Y<b]WKL24GJI:8:b5U5;+SAV)12Hc-.(<0_3D+RHO
&8c8OVeeMCBSI:baF:[8WF((FPPMDCe#C(=aBU?DTC,gJ@TWBMJ[QMS>UgLIDA(5
P^FRS&XS6JE;9CS?C;b4a;SU]ER41C168NFOXK.aW&W^7\?[52a#47=O(F?/\;UG
bI_FH+1&OK=b)fD#UFPX#P-cPHCJ&@?THa@\a(PA1b3H+[aY#P[UGd>7aBX3c@_9
NG^6d^E,,gFUeaY)ggWG<=W/gN;M(:aW78XM9LC9:0>-fe?]Pe_>)Ue+[V1;<d[8
<\N[T9L#WT_0DG5/P;:/ZOWIC5K#LXT\75K,Z5\3X&RAD@&/DCVea9]Hg^P(:J_=
[U2a@WHO&H3#6c,QgLW?E#Ufc?RS9c&>-c.ULPTM]HX\SF]3HW4[39]#J7LK6^(c
\)cfRQ6IUd1/.GDf2a50H:aIB]T4+[^5TSA8aG7DDc^L<.c[I7fY&VH2+RBOb:6B
<XL;605YQ-WW0SU\7DUa6eRA+2_PgV^00<.)]EBRNc&Q@dYY9]f.RQT8H1?OK4EN
2HI?\)@MARHgKDI2NNGPG01a+=aDSLeW,NV)73>cTFPS5g5;a>[GBX>S@cU<fFO^
C@^+</>aL\(:JQ&GRBfKTbM<\EXZ9+541S0T:14X;96aCOE>[JXEE7G8<E7&@.ET
(#Z:0KVGZ02G;&GZL4P&=??gJaA@9(eIX.SO>gGJI_bL)^ZK0e+)IEF^55.-S^I)
H3J0W))BS+MSXI0;_9&6cQX9c)Ig9/ec97WI[e3<UObFVMVP#)b33UES,_ID/=JB
CE/;\KSJ3d#a,LWeUc3[@fAIEB7Y??/21(D03DK=K.U9f4cf<\J&4G#11=3d,aC:
&H1D]<CVC9/>[CPB5FCO;^[:@JMD4&8eGV^Ga+)GHN38<DTa9O;9T3SJ^=HO@af0
0HGIDf1D^W3<G-\B7C9)+#Ua&<+-4H=&Z4dfbDX@J.>#74[bfd+^#H4X1eDG(N2g
D&gXV&N3:?O&BdZ6YE8U/?3bZVg6R,Y6UP1MY\CVZXKH9(_]L<</>d5?[ON\/NTF
/EG1PdaC(/.a6I-7-V/UA09BP5M(Z4_,=3EOf^[T-DTf0ID[]0?&g9&.Zd<1/)D3
X53_P,8OP--9]8.RF0R?[GUW)I(01Z2aVGYINDcYcCIYS)9U-<)f0+N4E?,(fLMK
Z@^d7WcDA>5HFeOX4a.)/N7d3[<;6T^V<NT[e2T,eBg/53ME:_(]F:PGZ@ZfEf1D
e9Dfb?PaX@5M1.W+9:Ug>-U@E_-N1J)TJ+]:XT9@BVGa(TWg9>1J3U=A:W2,A9X/
3=E]3Y-T4J@3A[0>d7WeH?3OS(1A+]([U_e;R3DcA-8[K]_:^:AT)\UMQMB6-MXg
OR9P>aS>04>3P>CPXFLQ,>.NG#A]^@HL[KdEU[d97-OFLc.Q@g,)-?HP3V-7c[MY
PQe5_7DO5):;]<V)MNb>W;/[AHVGZE3^P_UJ[6Sd[NUP,eZ84_ZXc7.bXD]UcLTT
T3@^QVWG(@H(<3-g/,IH:Q8E9fA4_8A:VHS53=8::APFb/9W[G5I)29FWIMGP+_U
N;e/JHcM/JE7X&9/8IC-51C#d:GT0]YNbCcVa\/f4@L&:b?L[&&B+(F//8SR,8BH
#3e&YOgV-_8GKWK7D6,e3I</gR4CS8PMQ;-GOHMGPNL[O[bA-cUV>&G,HRP9H]KB
/b2Ca,CK<6YdO#(V<3,DT?9b<e6H,N)=\+?Ra^YJ2Z5V^P)+)_LNP?#NE>D@ZL^Y
R)E1[-5-E]Y#>9].H^Z;J+gC3MX4O0&KI3CTdAX2)f15OG8WLG^>O0\,R4?[>Rb,
N;9,RAf8Q&=MbV(Q2KQDKbX.aY4BLM9eLU0+L+KLW<W14P_KRPT4W,0PVf9N<(>\
XEW4)9H^V3;K2M4=X5J0X95ecZAa(L&C\DQ0VbJI>DD+6&BRBb,WA[A<OX<]A[R:
Sg<\_:J@+a-_V&7&bNHE9GcALa?)ES56F)0/UW@dQF#0:#JAfGTRINW/eF65+^DF
21+9HU&EP=A4D9/3gf[WZf478][T4&c\B(a9SK=PN_9L=4WKE>CZ&,WAgV(YdTZ^
+L/fe:R]<.Dg.D>;0EQ^=+X<AA-OTA@..N9#>UZGW;<5K(0H)Nd/O:b58(K&-A/=
V89[e8I_=S;9cA@G6=]?f@)IZcHcI9&aV7)>Cf&-A#O)@B>7F__<JB-@FPBEe:&V
Sc^KX;<2=C0+Ib<(OM9J]:Dg0.O?[d+Y00ZP8DRYI5.b6WD:JVJ[T8WEUT(^2DU4
&@XXBFH01@95+C&KHP.T>Y/eO)GN&8ZYN/O?DZ3O:TCH4d\QbL[?FJMJ1^\&H5FR
4&N(]<A-9E9fAQR<2]<(HVWgWW+80-I)./0g</g:&RT6KLc7_S&0WB+TZ;QgP44+
bK1fLe5O#ROR0T1g0(\9Sb>32_3N\7g=HR:TcLTf4TUCKQ-6N<^D19(KZFAS-5B:
H;#ca^cHea/._L?OADI3RcdF7aMKZ08YcZ5/^aKP6B>()144LSBZ)A0Y<^893=:>
McGKWe6I5b6CBR;>>+NX+1L69e-;Vc7)>AbcC/V,CE,4IU4@G]LcA1LUR\Z=.5fA
b;O3UDVZeVg.Rb9Z^>N^#E0-AO7C_MTM>+D_7aY?<UaGTWP_::V,?]<a?LPRHZd,
85W?AZCgG2,-L4.a1YB6[&cE7S?cH5:JB9gaCVUVIYZ&?-a8_U7B^>eS(@&)Y>1I
92<.:W6ZcDY:Z:RA.L:8Cfc@IVBJCH&WN]0IB-#Z0ESQ+Q(7UL[^)3Pa[aX(_]V\
--0OUg(:N(=0WP]?YL7Z-C)W;ROYC#bg=81(NAK5-aQ:>a741[H.AOO-bDfU&^KA
F,7/AZL./EAP(E@)bLWV&,6__4ROE7PNO,6U[94LOGJGCbNbJe^;6g/^<U#JVaG#
+GR91[N_]e+J/4/_0NE,IW23&Je7F[G[=K^:EQQ,1TM;D469&-=e=X#cX+L\72O)
;UIc##6XB@-N:Z:L;<NTW5&LgGY;=]6X0T2WD;8R@db@DC+K4^E+_2A?;JL)d/#_
W,)&U7)POCb3d:XWA4(d:+C^e_EC=@O8-U6.D.])IK)ZQ/aOYRZ4f///JfY;MAQO
P?3-_IM>MP2a-=);+cC+4+YM,5JF#D/d]a<#E&JO2-[AR=^GARAH/;UT6Q5U9F\2
aX73;81++A-YO^&X=^FV].9Y=1S0BQP6CR\3(@MP](BCV/?N.ZE1S.865Mg9AAK-
4-JM9?b5P#XJFdTbgMGA6AY7W1IK<Ka.fR?UK@P.WTcWRTAY-VeK)JA+<EDVVQ8I
W[I?K_gC3afQK>EZGRP)#OCDdJ0(eT.D)eXPF^)(?_R:W&QH+UR5Z.8W/?UL(I(e
.Y9WP5W;BC1;(VgUfb/]G6NKO[(VXO>>5#d,\;.+3MQHG_.8.e4-N&K/d])N_c_7
/R3H98&J&=@H6F)g=R:d16+9?Zb(&ZQS#]bbY^]WN+Ye41Z.,CXO62W>R=+5OQ:@
WUP,fAP)BcfBE:6,JQ@f@I/]:a6OEM><\M;&JY.H<KYCc:d=Xbc:;]SHQCeQA66@
c+]\OO=gA6[JR:>S#A38_S<FgbeGD\_<S51S.^,WF;^EUKc_0Z#(8;?9X/Y)ISI=
JcDW5=6BaHVXVW7S5B[5CH\c,-]G;X;7DHO9&B9eZNd+g#,cFBA9#fMFLW2];=ZS
+a)bD>c9?B@TEREIAS0XfRO-eQD=]ZXO2Q4HMJ^ZU=/MK-#&cH,OYNUdZ#5CHQ2X
#PD+FC8Y?]NQ9Z6^.4P8J,DW:72ROQFcd5K80M1.V,9QQ;#c?GgZ_c>cB;\>;;WP
/K@=D,c>0Cb&W=_EH[:Z3C8N->G5VbF<e@4.\=cgc_ad4[g.<aG18UP>>=S6S,1R
_A8aZL9F[OQTecA3V&TBT)g79TVgCE^.O@?6TRW43NRC;8+.,K)AC6VB-A+P2Qa[
Q=ZEYZBJ30B+F4gAW++EF^,PBH>V5cge_EXIFHSWb5,dLSR^\8eP:caIf&5^+GJT
8<]V9_^R;GH.PeEDO7TNOQ4c\--0a+2>8>#;;M+U_31CB8@LdD@I@W>+Y\-eFZaP
b3O=1?Z@+C&8[O)/30KQROZ8cCFa:;K[Qe#/:=1VJ0])38RKXO8N&1O<AbUaBX79
O]dJ704&>Cb/4#S[8L6+c,6<WZa^?:9HA_81;^dFGf,PBM5]FaWT\)RZg3Xc,5-;
Ke;3(a6+2P=Y?cR(gT,2H+HL/(ZUV9Xa:+=CR\-GF(]+Y7-2Eg0>5NQAC-BC5\TF
:W7OR&>SP0JF78L3#5CGg0<0c=E5,F09KFG>S-WH)YN8f3-N&6>5O,XAPXS3IJg1
eOPEVKb^QJ(+K2DQPO+]FXTC\5NUS/^0S(2Y/Q>,43HG).S#TDCT2KJ#YAB#(UP7
W0XC^C.)&C#ZM-C#MLKWaP8\f6UgBUO++]gKW;&.U^],U?E)V^Ba::A3Q]f?#)E4
:>CMFJeaOQ(^T2VXg1cHQ6=UST6VQ_>DF\d]L4<S?0)Ce@4,2(=J@Q?<0DPRQLYC
V/W?dEQGLBDdGb@[6(&:HdBAO93Sa\,W/6A,HR37)H[BNU^]8NRS;,Eb_P/O98DL
XOI-Wae;W9BZY>AHUJPZ+VO&L0YEM6Z3Y70CPG)[,HVO7@)08<a1HUK=-K<1HD?W
8&#0_&BK)#A)0+&>2D#;dcL(fCZ@5a&),0=6M]LHe-UK#)7ID>P4OIO.;9/M-fbI
);(MR0<c&IbUcUBeOefP#91<3<e7@bS.H[bf6LOJ[4](_CaXd&X.NcTf5H/4W_DL
H_<MZ8:(X=-KRR(2CA&X,->:>>/XT=^7#+<+V84IS(-HM0.3H6f/Q)15XE9cFcMF
-GdEP1530)7E3[L2/],/S>7=HWH/EEHMUDA[297Z-C_)D3aY])JePT#BU&_:2>eB
2NfA,^dTd[H_F5K;H-G@W)3S6?c\OK+;I.URJcf<X>:C^@@08JD;B@D#OYD.R.J@
T7J&IgB6Cgc@c70deBg1<GAf2T8.M^AdYO\F[Sf-e1@_H;HbY4DM?RRJ\V6OIW=9
Z?YWRg+c>ZgcEL2H#C_(Zb1^3/SFaD3.@\]cXBGR=A,/.c>Yb5_+.D#<agR1&O=3
PcN9P\_Pc/MZ\M.P5bSgI0&\V)KJMeD=R)?K/7#9SMb\b.ID+>JWF]\IgQ+aAY80
cRS?_=<(MP^^bJ#6f:UX\QE13e[P480fCZ_OJ&b9AG>PKfI0/?)VcB:+US_.VbT>
f-4bX+FAT1U-KDY&I>]E;\Q>[/[&2^432IMUdTP8^O5?JIT<6)&La2Z7(>,\f774
VUc6GBRV^bEcU:IPDd^LJ(3A\S=K16fRdYOXbZ354^L\@Y663N?WMBSXBZ=5JH@U
RMA&:g:T@<PaE0Qg.GL;5V/IbU:D,PSO.&Z8_\S#\_90O_,e][0B+]8eRC>d5Q&\
J(=>,\7D:Z(<L<+Y8JK.I)J#SP07TMFG)>PC0HW-L&F<fHH;8XGe/Q9?&,^@EJHB
M1?2/g3,6CgWEHE\>Q;X1PTB((e8I=9VRKRg0(3L.ECP[1/;UeQDZ@<KKH=RQ[Q8
X<Wc+8N=><b,R#1B_C>>=I#<CFTS8KEHH2acXRF<1?1PQ#V7DY5EZ2#HERLM)b0M
cG?7_;RVQ^);M[MdZASEdZcDTR0[X[4Xa,JG1[C@^AIL05gR.C3:/J8-BK6g^R>E
X&@+B,b[IS3)da9GOIH[+bU[2#UZ6Q-GV2,G+T9T5GOgCb^VRWAZHG7(C6LS[FL=
@E+WGG?_;f#cD]@])CV.0+S=)Z<N-\.BNaF2(L.W9U3D[C+eVLU=3ES,P#[c=@Ug
-:+G=N@+,>Ca4eff.W4\027JF?Z#8eX3?WTgR2T7U,#BQE9[MOL^S]e]T8-UcAQ3
\DL9)^865_P&/XNIFVP;+WYK;#S@>YA/6WJXTUW#I4X4Z?LH1&fd.3>?KOT#Ze]1
0JY_RQL<Y[DP\P[LSL53M?_A45,A:F/VDQ6&8J[08:?2T.62:;4@WHZc?CW3QBA:
:M++O=PHT1=-9^Q[3?00]H=BaD&WX2&25SD2Q/J3HH#U^)(,]-QG4C#]8I8?M0]+
>6e@Z?Q#K-_5LS)ER1VS+=TL<416=T+])S0e8G[-/0Y]6=N^S8:G[-#HdeaY1IYL
Q;VF,HY?gWW2(2IO_S.KJ9F2)V2Q9_R#MF;.#,=;O:9E#3(.fIHcBBU-FCN?=^R#
^R)a24Z^J78fFA^_P9cOD3;-IIR2TL?1E3A7Y>/2Ic4SIFc.E0)I:^S(VM^gRYYN
CD@YM[AN6@^fWUD:b&G?>MGa26SeIB:5GMb];/=<^TT^&D-@Y-V<6&WPCV7#FP3Z
5[-fa?:XTFK)&K?_bI5Ua6[^BD]>CVScaKPXY.(#2Y:.SG212=<C>BbaLWgHMFE<
VV(@@W&_L,#<dc.N2))dEM8e[e(,S?c@DS>E/Q_U.F+O@A#XU:-=_T@#N_V?_\1D
PE\WQTGAE=.;?#3[C,#aGZAQ=#aK2LOJ:CYE/B_2?(OcGfV8+BdFD1G9A1G=<Gd&
]5_M<RF+FY<,R^AA]?++<#1?e,;[a&IW;RGSJ7=\/bNCF7a<(^F^7#<JWTXT]IVW
;=VI8?MQ@QaC;222)70Z6If3Z0FF^?FT9d=[E7TX^+LdeBU>d@#OaCZ;G5C<Q/QH
a-EQe5@1W/AH/7N;,RP1&W21_Z#SX/1ZVRNcbc?Gg,A_WV1c<T5<dXM>_=4V;6@2
aTCV;8S65aG;@]\dY/3GVDSK&I@LFSUY,[53F)SJB^:b7I96YGX>d+/CO>&JR?2\
cW/ceS^<1aNXb/Bg[b/RJ)G6Q\K5Vg58K\-[\0X@:dFU[_SGWCP+DI,]WQP@[WDS
XbLf8<C5YFX#6dS.MZea#OQF/V-.a:PHY_aUBV+R^&L/(C]\..PVSSUW9Z6&?=Z6
fR5A3Ud(.FJKU637KOaf7@/S.VFY[U278&/.;D4)dKYW:[>_]BNe[5CJ9:Q2\<A/
F>U10Z/:Aa1(U&LcX>2_[[FZ4O6JXccKH9Sb/gU:,TI9O_;5@TDE?g/)I+Z(=HM0
a-?,_5[X?22f3gCT2N<[98R^8[[V>3WdO<(DE4AIMc\g:PK;YV1aGJG>B;bWM^\&
Y\3;YT@+@a^D^4Ib7BU,FS?2V_2ORWTDNgDM)_=eH>K4c-:a8^&;)Me0CP_O@@U_
MbOHTdR&I-?XK#_Z)VfFK.PJ9;VMDH9:LH+2R1^6DCZe/=&SRb[<]DQbQUA:6=e2
VdPg0H]#UVV4UHG(4GASaPOY]NNEU]WAAS@5X<eZ@7BI6N,W2;Z-9NOfRH&;@0gc
;4E?e+E<=aL7\97KJ:30[B^J7LG-_N<A5HN3bV_MF/]I1HF8JUE@Q\R\9&5QL.6Q
550+IOL94gI;OF[:/c76;H?Pg?U\c-#9#7:9>[cJJa^0VOEC3W.V2gE5+[f#G>g-
_UD<@,cHD&YFf(^fXL?\VafE=>]N-b0,.PT7U/7P:1Kg/2:OUJGK6=SHCH:?(W5U
#)\0V(.,e<;8.M,9ge=(28N_OVW4dFcG;Y;(KD#KHPcf;9&1ZJMN(.b\L+/gX45(
[B>N+PB(+GRKDGV?CZT.I<^1M++/D?YA^=bKEIWHJ2/aK4KNN@C=;<F=.V,=0SD+
[VIeaP4O_TM).d&d,@-NY^7;0R@5Wd=gGb,=L&-[cX5J0)F;T.IJKZ_\:=beM7__
\?<NdB0P43d/DNN63T4;&eVD@FDZ?=UNW,HU2cEZK)T;cIGWCV<3O?H#C^VBc=87
L1OJJI950[/gQ;AGU):9fb<FfE(,[Yec37XO#/#We7>P=K4]PZ&LH:=QZOIX3YEQ
PVR&9:Z\]WCQ.a<;(4Y=86KYVW5:,S>3<IFL&^3c>AG^Mg,feMHOG&M5;AYG)/[N
eP6+0g[ZBgNXA<JH[=#>;I<8gI83T<MG\Q@UFLP[F+@W@gMV3=?XO>JQX\=,8,]f
<EeLXH3a=YQ8.#[^E+e[J(+MN#;c@X2]4Q;?L#BTHbK;QC=S.Jd=.T;FcFL9CW&W
-a?_5>OBFG77\<a)HKe1GMb=&GQ,>3H[]K8>U.H9SMFG4,Y(8KYD1LgRdM2=S8d?
83J)gC-(2@_&KRJ?:KM^RZ]O\L.+]\<NB@c2@@f[VI&fW/<]V@&KT=4,PEAO7Me?
=a?3O-HfM=\^>W=F9f(fEZBS/CYR)<=(GC.],E,RCLS_[+2=>@#L,\7CJ(gS_b<N
E0&:+1SWF_<b;\7.T#>YG^\\+3WOINV<(LR3S+Y7\MU\X+8?06471UPMFU]8+U)H
\ffP3E&5)<E<^)S?NH[05<&gSH0g3<aR=QJH]33e3E2L.cQ&1_7(,F\D3Z-e)UUd
>,GAFdL=A_QGZ:9Q7QY_U[)SS47eY@Ec2[9P02988&8MW_8X9A4e6V=FEABZ;CSZ
f3T/LB7KCY6>R]4ddO@Y0e?YHEO&TSHJ(3_a0QUTKg:A:^7&Z:+,HFRV8f_F@.-8
8<>=C0.)FYRbS;];4fY/VN8)T6G(^[Mb(FK/E27;SF.<G#_ZA7+H\[/RVU)-8<<W
1V5c#L4caQ57=>NaaHG2I-]7IgfD).QREP47D<Ef>gPJ<HP;2N=X,:BDDL>Z3Zbe
H(eK8,&BE54c;&CTU-,D1J2]4F?M<DQSH<_6CM=0F-^Vf28f#1?f.BK/D8L0GgN<
Nc#d+H0.RC:a+\?eb14JM@aK0c([S\+daW+?A@9K_5/1[eK36Z_HMefOAFNTT,Cf
9c3Z(JX6N,e^MS/B2D53&6(@R[)8VF]J#XV.b;7gf:Z>JGHEC4STIW9Y@cYKGXBb
T:DG;>IK4;3WL?J]8c0dK\HV](_H6CPAK]MXc6?Da+:3D&DH_D.<e/2U0fF^N3F1
F:A[.SA/YCd:-0J;c<,)E&C1.].O\J2<LVF/Q^0&U/E]W=Y6CQ?.GEEHHM9P7?&^
ZOdTfZY==Dcb.2Q+/4AXMO\QZgKGERA1N1E@FWagU;=Y?EKST:F&,Z)IGU.dN(9+
7)-99W+:0eK-42U<93DZYV-b;T3+Fae0JFOg)/eJ>W1d8U&/XQ@(1f(#M^FVeZ9W
1Sd8:@Td6820d&OKCdIP<EBH@Z0g9,K5#[IB@80@WK,48T:1?4P]G]DD(/SQTLc-
d0c#[g4J&QI-FfQF8Z#-A)8.U_F^=SM;_f2(Y?JMS-0BY.4G0>cTO-M1#8(J?>AG
X)IN=\X7bL\GO:IcWFC,3.#EJM8[CA\.YC(IHPd.^aFZ7>d]WMJ16CJ4<Pe@8c<6
_G;1AP8&T@D_ZJ=3M)G9]>?cOPP3QW4.,d0(ATf5-4E-OG_>Z/]b^&,N_3Q#fc^;
W:[]YGb?a-LP1Lc-Qd:[;e4O7(0cKT[bQ<D,eZ6cf8OU[W+FQU/Jc8T48a:YNN10
A\]dD?X9=0VD+X(DSK6OJX[&.HUX_6N2e^K\MV]a_#.A-FCdZX1F1@Q8I^01gDS?
B(V5O;e@I1V39ce;&ZdbGQ<\/8=[F.4Cb_)+fX@=[I]?d].>AR8INN]X8+NS^5,+
L9Ve>_M)3.7)d#R,fg=T)ZCKL+FV)Ec(W+?:?4N[g4fB868)_aVf7dOQ^C5C;XWX
->cd)\<@5@JA4K(?DVRY0UCI\?85KWg5;_;2@9^A,a&LNO#U?V0c38MT?N:-#Ue\
:&TO,\DS3f\(/N5@R:J>VP,L>;;+8UfXM4V=9H3N1EbTg[S@UPfKfg;N_E=ZXa&5
CSZ78a?25+?aS?2>].8eTTM;>.)V+=f.3&R7g#JYK:b4IVPX^,4MRMFU&Q^e=aH;
KW=V^U6f@2^^fW-;N&:9b@^F8Uc[UI&aJbb=]T2C=K-,(g:5_E(JQ5GbJ392YGT9
#QG2;QF^BaUYI<a)309714V?a>f+:=3_W2_6,Hg?P(e?:+>bQ.RfU2YC1HH6.F]K
P.\K6X0W7LfcbS-#LCMTcUS#>IVXXOP[EXBP4KJ,DLJ=W2U#QS<9K3+Af\?dWPE>
HIbKT2.ER[9FgR#Cg+6a-\C>e\aGAWRGQ/<P+L]QVSd?YM#0Kf3b9Ef2Q0MXKPWG
3dF4(3&/=E,+d7)#Rf[8+9;RE/^6+>CgEb;-S.XN&M?3)1C[#;B@9SX?d<DK<@+c
4^NXa\aB+4L]J;@30D<8\-QP;2dRDQCUPCgf.Sa2A+[UeR8TfDED4:GD:._JK-75
gAe(d(+#+K?.G,RC7WQ:N3DA+9#E;\?fa1EM_b=>Q5-g.RJ(?XE)0<eE\aRdG:f1
W&VMgaO.a2VVN=SIb:S?7UF(TG6SDc6gRe;_&RY9K=BZ9ZSE3E_+&P#D,E9=AQ/P
9=[,_GZZOHUCF8cZ2MKPTJ5fBB(/^cITG2TFP0Qbc/GWS)P29fC+7gUM_-(_,3V3
RL].^JJDV_dWS0CBd#MF[_A+PCU?>6_gb_MHHe.TC0&,H/4S2)=_U\Nf,RWZd>Z]
RXDQ,R.-fVT_:-+VE)HFNN^[N]+0+EC6K7g52@<>b\7<(5IRQ7/BfBLM2Y]K2MZF
[)\d]aB^/-JQcD3fY,;B,+g_Z?4^c+O9;@,A]P[(PE><\+Bbd?5b>>6[IDFd8#W(
NJPD6Q@?I6eNc^?,Jfc2D_2b+<4fMR+-\E#1V@H#^fY<SRWAaG36<1E^Gb?GeeW>
1>4^HMT-JMA\7^_MH11IZ//R^D4c\Nb3QbO_Had1)d,KI5S?T/K)H-&QMXVXF7-]
C>AAN[N/A2SV2-gE8=@3(27a.EGWcA4C^O=R(+ebS0V6-:_YTR5]G=_7=GM3_?Y/
#7J^Ra8_]G<:1^cEJ[8X-fb/,g-]/?cPeHBNJTWK&HAD\:7KET6758[(#<=S8J_B
c3TD1XXU7^]A1BT?+87.(a\^9B<4X:7Fb02DT05?[@Z\/_Ga5a4Z;aF+A:Z)NOC&
cU@55M@bQ@T9X>\1\W>VIDSE[afbM6:?+DH,4:a0<;]FdM8KY;N-?f]D_UJGEYG.
OX&YRJ@PE3./KO2b2M=3E&KSHSETTgI36(XZRb7U>?TgCC@9XQ5&JZP_LG4#^,[8
>(E5-S\a<[(_X^JX+>6LUIP_SR&_0^I>N#EPc;#V#S6=4<_=I)Nb-?(aTA2>T?))
P>E]d>#OSYI;3L\]WRATJ8+S1S.BU^d)HSc<B8[J]_Jb[a9NOMQXA^.^I]@P>9,E
;Q84Y744Ce-Zd(]-C144;dW<K0U#QBQ@eE]JBL.F_O>6JZ04BBEY=)@8RO1TPH>N
M04)#_#=M+)6a:[-A0#B9aBcf#(,eCPJE0IgdcdHL0-<bNdG_]VIPT=1^>gF1<6g
8.fZ[/_O?R,<ec-1@OcW)LF2ELfSM1F5g#BR.&65D/0EeT\U=[-<cW]F0FQAKeI^
W&33IMO?CY0IH\:\?_Je,a9JZD.H)@G;VN4?aY6F0c280L#a2Qa257RUa6VS5PT0
[gXgL9eN9Y:38-&JZNPJG2/IVGLUQgR[VSB)+Mfe;;3G^/9g8TIA#G(389eZ?/L3
-_BAXL9L)8c(1ZAB\F.Bd5OM;(/07fE&-bB&C..^Z8I,6Gd[F(BOg>Uc[/\,TN/^
^1Yb@(/06IYNFH+:.M9NeETW/L5BRD..X_FWb0F0N6Kb:a6+<EN:.+O=8WUH<_3S
KIEb2&?)9?6O50A:TUE5RF/@<4@=NS&T5eQFeV&3<D_=NYOaRLCRY;6_B0BR_3Y&
9A7P8/\E3<EPCZ2O3XEb>VF-b4\f&bW^=IH\2_,2DP#KCM/;_@LIBMEE-K529]H\
/C,C58WG;+A2R1bG#;&<?60Q5?T:2ZB]6B=,84<:1PYc4]:^a05)@FbZ7bSIHNDb
8Kf:>WW,+c4@cI_DZ1PIVH3d^C8Q)f1EOHc+84cbLQ,TG_20Jb0#HKA_3eE?X-db
G.<<VEYPa[a(P?0F+R[/51]QL(5UE&><.g#.WKK[g?YIe-;N7M1g]1[NPY9aH&6M
KGZ))&+^@>Xf=R(UI<f?A_6>fF7TW-2-,(37O_G#3^-8;HKG<[LZCP4E6E+gZL18
\B]CDb[CYZe7U.W#D<Na[T/W@+]6Q-B#-/gOa24W:2/e@eN<#=.ZFBMI05&+MY8,
E.6U#UF][f&E,(&ec9[;<K0B27L)0\a(?37T(N-V=@@B3@-C)f0C;XSXV<K+;T^K
?.QU/9,BKeIHP4N^g>b0B:a16P/d97I5^fL-UC#>Jf?5\1W]7WV:D5L_gbZR3GgN
;XOG6W6EP6SXRQOEUHgP+,XM/^;E+#.006g-V<=<cPOYW=G2>f//LCYR=\e1CgL]
F+9;[U._L34G&9+N-?7(Zg=g7R:#^Cd3\V+H<_VZJ(9ZW#E)Ha6VM;GE@X(MVHdA
@K@g[0fKQ7_1/@K?OH/4X007_E_LJ46,8/BJg539?\@?>[cU<CT\#Q4YVd<;W#8&
Ie)GXBM(DeeBZf530U1A+UFd.JR26>QK[TKW+^dXTN,\5FNKa8;W[IH6Lc^S2P7b
E:\9@:[Y(B(H0e>+M;@R;9[3_BPD.HcCdL_VT\gBg]F=XZKB(N-ZcKBc24dN7?\E
6M188=TV/1>_;c51QG0&>S.<cU^IK&?O20X(.e?4BT<3C[HF?P@EJ#,+<+>&@a\E
cEW1d/.->6E>fX&?5M9&UJ&5:7O4\#C^[XD-NfEeOPGDUWBa&0d5O#-a#Q4X6.[Q
QZOVg?31Zb&JZC4g_#.===L2_C5P=7],D[SRZcI6;fgHGa]=cD,3(Y<Hd+0+_H^)
T/0:]:]JDY6.+g0]^<PI0HAGN?+B]dRLgM^W,?RbLY(#&L\b\N_-Cg/dP4Y#6P]>
fLHM3DD6GG,TEN+749aD7fIGMP\cPARD&)ST7@ZW6b<b.6O?.V4Q?U(\e&&J5^#A
^TN_D0K+M:P<F2+535+>W^BV:?IH905@QNZUVQS<fFB:]b(0DU@AXICDX(3;,]?a
?Y52@TSGJ)(.=9&&1A)CcVb2AE;cEf(EWDJJ0^D.^Z[Dg3(/NMQ7TZ)UbP5]d0);
dSD9B:D]TTgVeDO+U1TbP3XebNaY^,(I9Y&EGH:XBc7K7R9ag0..G74RTNO[Jc>9
=AGQZTLe+)UTg>(<)G49]4XcHG-7,5F_U?.R&^1UDSD397g-\<2.W=Ub-)9^T>KZ
\NVAd^HENKDdD3WbGG?WG2IACX5/FCU^?N0BMS65c]P3\eEKaIeaKJ-(fgAF<B=f
Kf.6X_:@,G6)HOGAU:2HR+@/-#?-.:^b?U+La0YYHB==036&\._4W64Pd>\(0F,K
ALE?/RY6g=UPFT2/Y.d><0+<KT[LbX\eVLfc?.,db+V;2;S,AF_B8L/7&L97WP&a
:X_7=9:=LEf\OOC&4b>@0ZN4;X[_McPId7XeP.>GY-#FX2RbX&(/+GD<8ZbCc3fa
QOM3J^5;a#@7K(4/KafO@cd(cbHc07B[aFBc-GGI&^#X6Q52WCY&#f47.D:LU>K6
U8O@0ZZH1KYf.-<TDSC.P;6&SD#IUZ6E?KIXa5-[)V<e?IHG6RT?f;>23e/UU\V7
dYKTeZDX-g3g<TBP1T]bX+_BQ<7#F_efO@1OW,UMb4_&Cd60S>cXf:bGUID.OW)6
:6d-D=4TK)KZ2<O1U@D\A<:a=AfbYNZ)WB)B?+QMa.VK-#a7;Q(f,7ZGYbA90.?D
3?(BI\#J)b^FPO>_XY/85.Ha]]N[Z.R[0+V(0F^F#(fP@8#IA>J(1AKa31XOQ^91
VJ@C\-D=#O\-A.@Z#=ZIcM:]I=g]GF\P<GOF#f_+aZ1Ee8:5M/<3;V.E(Hfc-A(7
B.:-Z14#HO[JHd_SCaNAT#/FTRSO#5?)C+KFLPE]M2#37&J>L9S[b]//Xc1=e@]<
W4&A2GXAV7TE./8.1g>G/FH2-OR(NBICa1_ggY(QecVZCRHMNFE4fN1^^fccIRL[
:&3X]S6H&O6A:9I)D_Mbg_11(8M7C0TWN,B9\0S^_>X95DMg7McGR@AIfKg?55.&
6==W1<W>-4VB^P)5HdH1YYSQ:fBLTI(A9f^R7OV&Y)I(=,HIGA8GER()FLI1f<T5
@<.@+f;N2e:O=B1[WLZ9G0WBN8V_&2E6#]_&YHg=GET3,^[TRBdXHgG[4Yb3&YK2
:VMSE-;Jd;5NF,]I.87Z=WSEN_Z38LMY-:ELHS-YJ^]YN#[ZRHK_M)6SHBUM0JM+
-:H6)0]&+NHIK[L&:67)=Q#YSLXdL/MFfZIV?487O383OW&3Xb06.ZHga2;EU<^F
0G/(0+)?/F2SNF@/aVec;1#ABSWOdH8#BWZ<7Rfbgd83\GgLS9EOUZU4W3Ke_F+U
gQ34>RPC,]_B0\#b2>56G<M=_JG9;gT3<b>JUA?gQSHe^>I7#+e0^]XRK,JKS>;_
QeO-#4YJ76T3U>T=DC+cTE9AHV.aBbZQgGX<gI9,?ZC=MXKRb<VJ4M]ZUSfQE,a9
<CZX/2/\U;;OGGNI/[NRQcW??WKSZS-5[@RT/>9HCS]&>ScAU3<^+QadW\=)A8WP
K,dBEVI:Ja=7X36YM6_&>cK\6:8,7eb+GCCB2&+&&Lg=DIREX6:_&T:gU4CR.Sc>
I4X()N]T7([\K:,AdKd>ABOUK:K>K(XREY2<0I3[HO4T;H6C_N4-fU<[RN7:;/=Z
+=Q27==0OHH)R\/US?d#KT)L&BSQ1IZ-a;8QGUB\3dCPW6?3fGSW[(XE@[:bP9b<
,>D+(9_QSLaXF5)5+>C/2L]K,fN7Q)bTJa=?LdAb<Y6)O@H:bdbHG#IcgOSL5>RW
Q#BFO+Z7VL=K^F[9MW47>CH)C,B9c^R;DIbbLT_4P363ge0d@>E<UO+?WK_L@?PK
]8C^F:,dQA)3F&-,51AWRY#B@J&8Q8@.HNC[>,X=I&aQB_<;O]JDO?28QH5X6WSf
E#GUS^UZM+Qg==SS^)gSZK)@8,7HL&V_)(Ncb04\,#J??A6/QT\J0F:^X9K/=YJ#
#f&)<7e=303]F8N:IR@P;V^4;^MYBQb8(c2Y:R(.,XC6D?DS+XV/+TZS?3Q6E]0+
K)ZL>M\RQeWWUcH;C:=CLT&_2Ra4]T7[JH,E])-G?VBL_X=_V0A<6IYQ5]g=?W(5
G<T<0H5aAHJ(DEfP<DIAF_-Kb/MJ)5INJI]G)/02OXXUMR[M>aNM#R_e4Ee4>Ze3
fG7bDYV()0Y((TZQ:25-G@e[+e&EP3CG.-A)e@+&[9AR>K[25.DdcGSMSM]XF:[=
TU[KWdb+UWEQK&-d&SYead&;R;<E7b<LFC6b?2eM5VW]GgCQN(LLDH8TdLDK6>BT
IWDg[c9#;&S,fLG\<;Td;&VG1:>W.8\[@4Z[59W<5XY73baAA4Hda)]O_f(VLXL&
7E65bP62+ORPN.dNN\U#;f&L;<#DeK:;#]@T?K;B8a:[RCU8KL(\CI0f2?W&I?>@
HG;UY-[^:7-3E8G#O.<-0ZS(K#Da0S1RHI>>,(V48:JS]-/173^PW,QA.g8>F#g;
d8/T;cXT5(&>[AF]N,4VB+]QUgM13M8GN,K;+I00P@8YGWe/KS([U3KC]UPB)9gO
2/Q3c<^#RX_WF&?a6,/<QDBO[;-89NGadWW4UYaVB+420.V848eK&?SG+94-69WL
a9G2+f&/.;8b\:MN;_=;&>UZ:XYAV+FH)JN7GN@aBZ^J2d6.R=(?.;/T=fX#QY&Y
ZUD/Q>OPdP<Wg,+>8IK.N+U]+[/4=d[>]/JF@HK_6,3X:Q;0]8X-2)Da&A-b?:5e
6bB(G8_:c#4?MPP&GVB=OV8IEOVU6\IY[ZM\5b9?-7[dCBL5f_O>Jd4=T2TF,AT0
&3K7C64KQV<U3GBFcB-V^W(#_?fa7dY]:,SM49>XMF3HF9NYc927Q[bgRKKWR+ef
,G(8WFcJB(MJ>IA2EH<L4-7Q\4O_cWgZ2dJI4Xe<MU+,TJ[=.LEX4I8f]2#O6F8(
F&6I4&/PVZL(MER]C3L5:gRE8MF/fccM3T/cHQW#?Y79KZbI<9:OHDP6PWDf2][,
V[Z\4&\3F#,[^KDC/]<2V\UN,><W64&>0/1b^4.5RW)dNGLP8]>9_IJ3Z;9;A&4?
a)N8/>a20L<bGMY3bLZ,T)_eeSQBIBP\W-S(>77If8Xb\(EZ2cK[+/ZA1,UI><Me
BOTD_GbOXeE.MLI4]1.0D.ZFZU&@c?eC9TF[W.V41\GJ_9B1<7T(Z4WgV&6@,>Qg
1cG5aW+W&8^H<3>C003R]/?<^d8B2A(GO7D>)H5[.+UE5\Q>L@I=60Z3P0Z9NNc6
56[M^c@7OaA@#T?]8Pa0X/;RPFNP-C2;QPPS4S1]U(fP=<Z#L]5=QRP46ge+^&K7
Z</_?KWE;W2LV<[2Z4U-3c3g9_,M:3]K<#UL_^Mc(P,CT+)C.Idd39Z+Pd,(#VF/
.YV:dQ34D]3V64C>4;g0WL?8>U]^(5PPK,3Z\W:C90Z,&9f3D=J/8AN=D96LDc/U
+92TIVE;>.Z\K@&g(J;\LI<Z\BWRJ9]+VU(IV@63<HEY0J/6TB&GINgb2]P5SSLM
6b;JK6V5B\7MBeD6.ZTdQc,bDW]-U0c7ZA1?]I_VE>YR&E\C_BEV#JUL^_RD99=g
H_^Q_g9@MQK(0eTa1\837(5MFNX\1(=;3,?Ff>gK15>^gS\5e9VEJF#)#c\Q+?ad
cZ\+BKHKV/YM:Zb)MN(_>;d1Jab&]95+S?a[cDL_C.S,>7aSa36D^S[S6ENW<<>:
E6T\Mc/cf(V?T?c#0HM3I-Q3/&D^+g2^:EOF+09_@+ABU3/\B[=X0BILQ^bg_8Q]
bTEW@ZNB7E4P[)aEA7a8@E]+.NN#?8T^/C^dK:]>U#b)#UV^I)4_A;WY-E&9U1[b
Xb4\_H-Z?:A(DK2>@?O\2+I4a&cSF>c?V^.9;K1V\TG]O(g:Q>/K6<M=X2)#^DR6
JLXZ6L&(ZOKX&7QER\fU/@F2Yb,08ZbLWI?a\M)cdF>U6)7@aV=acFGNT-&3+WHW
SP9&EAG+J27?;0<(R;THKNfQ=0PO[G52[,g^:U:W9DV.N7[9<8QO+eXH^278eVb6
SK:GDg#7TJ1\IURD=#]VL12D5L;Z(;6?\Y17_,_#6)0D&fX>I?Ocb/a\0=NZR;(<
8LV4TG</QT&WQ(\(Y?)1UTKf_(E8e;Q_0YNL#&89-^/P44>#/?AUWU[J7P+dc<X/
H)[=M+P-Sg=FbSRB@e)..e;?[=S^2VB.<6>OV@dbF7RPLGE=-7;/KBS=T.5X;6V9
H,HG<9cI6F7J@+];cUIX;IB375,:ASR/&1gKD.1=@Sae0:F2L#g3MJe#VZ6/X4C-
DI9d2Pe8RMP+@@0ZAe-4KQ?>11+-K.c^<6-+HVD_0^_X7dIF;2HcCbXND@[DJUL]
(.,a[#Ic#=F=>>@?b,4/_,IFG_O4_RT.OM.)MG>34T]@Z7?>XDRXPH]N6V]LBf5)
M#><><eea9eX(#UO:Q.>1],&11R;8dQ<N05.[0\bAEHVM3;bN.X9G>[@&3X^\,FS
WH1X)/1_6ID8._agfS]I7<Z4JIa6/c:9TBDc/7YT\/4^EMdD7,2NT),NR::1-_E6
B9FUgX,Y-9Feb@),MS+D.bDY@UA^;5:1IE;;H&VYgFW1)Z[eGUg(_;^B1RY&.FB4
==?+a?Y@WK]7(D_PALMZBU:A(g.VCPaUeROO0\c>\#fY,T.H9&54.5b2Oa19-&K]
;G#P1C5g]<+LCeD4J#=4K8P_9b6FFbVeLJM@DdY;:=Hd5=YP7e@(a7F>D25BVHg_
CR-6X\+2LFZ/:6GO^G&U\#=PPBZe?DV3R9@2HGWDW_Sa4CaG;(IZ6P5@?.M_2R>-
&=a2F1@6M1>+\6,(P?QWN9[7+/F^-<ff,bC&8SMP4eN,(-KE8fK,CKB^=T]#e[1a
JE.X\b6GWKK&1?gY6O\W:M&].g<,-Pa==SZ660<9U,&7C+g,(Q>.f^@0?CMUI5g&
_-:XT;8#XFUUV6[KJdUG-JdM#R;?,;YFTQ,\bQ<7K6;3Y\bUCXJ4NbM>V=Q[P7A#
faCGQGZMQN9;G1KX@,85EFHQ,)cEA37)9L[W]/WW-Y7.8Z5<GX15\#L]2,G&JT&V
Z\5]6IT[/.cUJK&c.WC4#e.T-N4CaI/C8=CRDMB98CT&/L,^BV2;Nd#PKG/?Ng_/
X5R73^1GGGH@P@[2;ceY6bb-9J+AMXYcL>1#M/JAg<2I+IQ(ZF;;7;+MQ@H\J,Q,
RBDP&E0S=;VfVd94LQ>a.2P:@[BC#9+^6ead0S?4NGFeO=A69E.JWA(;Q.(e56[P
XY1<H_SPeVb:.+e8XOL(>JF<K8;JdH:9NZOg^6ACKg[4&YAX#)O/NBN(7NRW/?A:
bRfPF19ZcZ=313W4?PL&^K(-F9,@#>#9:Q:ce7K,ZO(ab)PHY[>c)G^/c[CO7d&G
FdR.7+^e>WJLNP6X@FR]eKB&?4UU03X0KH5&6b37J-RH&ZD[6Cd/25dS\9X[gUD/
#479MIMJMPaCGHf]I/8]A/5JXWQF9NKSFf4?]X)E0Ef3FV:AT<bV76-#,UZ7NI48
EGg;b)^-#ECB_GRJE-c#EBH\[fT:.==HWgDFPPKV_Mc3[d[G].VUVb:O8@Kc:cB/
#CN:;#(VJ-@15G1\GQeL((EPKHQ1@FgR)Z:W78g1ZK82)OHTVI\GS75fb8+I7\1H
fG=[:N?b1W;ARJKXSg.(@S8K,PMW_?TdI6(CFg3^P3CDe@=I4MHKc<We],d&__8d
XKW=H>JK>7PeDIRTO>c),ESUS^f3G#:#Q(g\F\UL.O]^bT3>A:;DQ(L(2?>Ec[7G
EYFacDQ6+R<3/,gRL<J_fRFcK[E_@++#S@L?\,SdU<de6O-LOH\H(WA\>cQO[GV)
dJG?Q:@LRgadgRZ[SR1Z4^D^M#G/N/b3Z0LcTf;JX\ULDTdR1KJB7C8,SD_,(<#O
4E8E,G@0/DLcHKQ68cEReI8G05;U>@+&2a4#S;QA^d^[2K/cdf?Qc/>G#e/MdTH#
>AO9W.A52U)fEU2_F:=<A4f)SDa2.Q@9Td@?8QK,)?G4KT/aR<)9^+@a#(ePH@+W
Aa/]I5_b74e\T;JB],VU\L^V3gFTe.R=3a42N1aG@V-.<caY&5V:(9HOH]B\QBgT
=S:UIDPB\H^IGZ#A2O(bfWIH,/^\.4&TX6e2C1NUHV7&Xc<S>eKO.XMUMATIHH?;
A<2I4WE1\aP7;aVP8Dga<@Xdf]V0.+K,>R_^=1dU7Dc;15<S?KcN&eQE<X)WY,6;
YCfbM@b-1=;/9,3T-BB(=ZYC6?N1RTWEOUAIdE\<^@-2Q50acabN_&eHLE8GMY/5
&?@K1>3&HJEOOSTFN-4A::K#Vd3-gSC8d>VQ:G<G+=6fbZdF+E8eE-=L,],41:Jc
@=b_D.94CBITE^^NH;7,-bYS\dM\<[GefS,-(EZ_RBTSEL>[1<<D_GB#0e;gY7W9
6PZ5-b;C>-4V[4=TB3BNRWZ^0;75O-^GQgd8_^JC@5YIRDGg+8Bc=]Z;7]C531X+
1]_P>RZaVX<M5;BZ,]Q8PT&_;+_H-_4XY._7+-2:8G;-/VK8(&[9/BVT#(X6HL,7
@^5B&E(C>A8PYaR[Yb9@CSc-dWDJNFGVD\Nd-,KC,20/dgZ9>:T9a@ZII_C\JS4[
=#c?I-3\)7,O^5N6Xg2;6e#_P/7&84A]V-1\WXGb(+DH6<],:2=9BC,;B6=fD:V7
FUQ)Lc6:ROZZcHec-L5[_^]N+I=[W+AS[QNNUYcD(1V>4dO<c_3_3;(\FL.8a69Q
+#]B:UTE)=8>b6gb#R-c),63F]_gION\4a/-g(WZ7?+L0B>Acb4fTAI,&FG?8(H]
VI[5><YVe;S5g.N?WXW@(1^;.])77cQCT:VI30:F+MQ9(WEXWYNVZ>]CC]8^0D4,
5IOb0f6Ce/_0&YPICe^#;<3F7eI[TYa5CI2;[2N_)3a#B127BZ5Q0+<FO>FN-2f+
#6#C@&8A]0,DTIO6:^_8a(6\be9,\8[-.ZVKcA57R_b?g03@Og63.P+Sa[\M=_M<
/7?UN;bE_gVd:,XE?Z_?X2@C;f-G;ZBW)0LS-_5\N7GVK[0TK1.9F7_+gY;_A6EM
[:G/\@]\3.bI?,CG)SF(_;3:b-D>77=ATN1(DG++B;72KH07H5(R=1A,I,-?UdX)
?6.<ZUB]E=<F.b[-PHCVAG_6LPR,d?-9P&]397\94E&Lbf)AM[Z.]XX[X<F_M^d\
/d/f?DaR/KA)LG\CIXY?ZHTIV^5B;8D8&Ab^PS1M;ADD+B99fJY9d;EKW2EgPX=9
fD4/f,.F2^VPJU)@ISE7AK=YC9A[.(8\,3NHg)IMRE,_327\T3/I&_,/1^O)c0-/
_T[aLbE5YXdYV4-44@61=WZP8NUKVDD5(,5&:SB7]cM>@Z+>?>aJ]O/G;]Xb<+WZ
X]3+0UB^;L&JC5fIP8IeI^8>/;_HH<f212N6.HU^+(+):eRb>@KRO_A2TR4ZVe?e
8agGYUAaZ5H.&Xb(GVJ\##RT,c5T/daKKEf7[<WI&NgFA0TAMNO;E:<&CT_FVF2H
-fK](P8YR6(B1NH/_KQ2A5e;H[[bJY^THd7?bEVKg[5:g93]\6A)\XS3:?MS+1)3
QQ#N)UfZg?NY-E6ZL4I0\U/1+2eJS43Ed094S6g5\#.?G_1We<^[+,.KFf-Zb3dZ
gVU\[8ML7A)/W9CCQM>[7.MCNcg\FG-1.](#Hfc\/^N>FXUc?(fDXUfa2AfdNMbR
E,+=>.ea+I7g[FRL\1OLT_9DZD.0gafVM=QEJ0UR9fB[.-05HS1O#RBdH7U>6eHg
CQU0O19:1SOGMOIF(&g#bPd\#.@]2_\0V6G/:G\;<e@F^(O\ODG8a)#/I5XCI>P]
-:SXfJTR-H[J)(1D9ZYg9ZPMLD&(R[6;MID04^2:72I?[D3I=B&J8>0#Q@6[&Z#B
.Z)-Z,V5@&[#\D]H-&/)Xd=5.K\Rb=1<2#:CTGIJ-9Mf3AE8MC)^&-)aN9P#e#>&
F2DD5+DFI\ac<2_MC9/g^aIZB,Zb7_OYD+D77L-?cfT?8[??d4(-QUY-5VK<7)Db
#D4H@V>F<W,MdBVd>OI89L\7+WPH:c<N_YfBG^3X?5]N:=_H<RL;Cf4_&BJWAe<f
L=_f@E]KXd=+,AK?#:2PdS,5/1OWC->G7,[4_,HPMOTVH/V>5<@Y^<bB;78;;S.O
VCB\6,Za3PUca,S/@=AeVS_L0A=McOU^KC5@<&L_;a/K#3PEM34WWbJ#cZ1HY-I8
aKW8JXA2Y5?__S:d/V@(4]+>Ic.>B78@+<gOGfY=>_c,F7Wd+7EIM^add>1C-5Y9
R()eEJJfc[O<QJ966LYcI=+.:6RTD_:PG7_Z9DA6=YbP<0FEc8-X/e/&2F#,(TUb
059W]f+K2E/3[6L:)aUJ]gA,C1fcT)Acf8[BB[<O:_3V;aD84[GS@S[R7ZKY89C:
;Mg;2[SHc&4AS8^[4;8JTP<RPPSJ<1B=EM>=Wa@?ZF9P)0g-;g\?5.bg<FeWYB#[
@=F&ZLY(9\HKZ5;^72JL4^VWXQ;E/:(\e<_A=JKaC1]eGC)U>7B3O)=F#?;HO@O6
5QDTL2bT\b43a[.0cd<873KF-/X/9-]gW&1c@Z:U.bE@T;8H]O^>b)GBFEAe+2?e
FfWG0Zd^2JMADK\,dI_Z#Q#@1:da2@_b>^?FIDgT_aLF<(K#LA:LV_O+JA\.<71Q
b(4f96-#&c2_a<AZYHc8I5F)-6Z<U:LT@@96P\WNfg28<&7U(\_fc?C90O/ST=U-
=d3gd3&e+A0Q)E,W<L+^ROZ7dTMZF]#AJ;JWV:Q9We@WPXBKBb6PXCOb^I<76)7-
.0Za@^6^-0AW?._7SKLDPYXCG:\NZYAHHV-A/ZA-+QTBSZ9[gG2(fJ-D0HX1D]<4
f3MdNUc=3c>4g;MZ;).[aE9,EUKV#MN7NT@cSMHLND^#L]V3K\I4RF@+^^[]:,c,
ZGGbd@NHHd6HN>[d(aFULJ?EUXZfK4#RaFfO/MD@U2>cOIA7:\<4LD;YTZWD[[MW
Z[9<T0d://4I#2f)QH23I(+&Yg4AT;?<K:^AUd(_G;W#PcEY^M>#F-A4T2a9)ETb
WBE#^:VYa>>@f>A[F?R-HG7f(_JC\JO?6EQECLMBG([RZ.0DP=A(eWc(.\X^S)7\
NW?GZd/PC2>YD&P3<_T8a08IeHfC^N_#/c]Sbc\_DccRL[\L#UR4ADFB=;LA>XQY
YH&<0>W/::.[+Zd2G>10=)4CPf9NCfRLF60Z4I2FXNg?Y+,I3.)0:ZL7)?TR:fNB
B3D-<cJR9A)C(&CeG^1_+T)74e@\Vg@FWZ0)\+Za))EHW8#?dJQ+K(9PB2WW2Re1
dUQb@<3QTBQ1IYe4MIf5SW):=FZ<YWME8JTTa5VbgOVY<>@7A=L(&8+BUF.66W]P
0<.CB.<@M.-^Q7.d>EA-C0&7d?6+[a/G;Of)b3Y,1[dcSQUS&=aE,b0?O:W2YK(/
Q4f[][)[ME20JIP8LbVb0g9IZ4C,+Q69A0SG[VaFb]IB,R-7+L=Zea8ZH7[X,3Lc
9g)YeMJV?A_Q^]TKGJ)KXX65_G\A&52F1g/dH;H\N;EK@b;K&_##P4J;4AZTK1)M
_@CRYP4_RK5+US<@/V[K_?PbRf\JC[=QW^P;E:8EH4SdP3P:f#N8ST4S,<..N>GI
K^792-E<,J=cC(E[@&8F-T1RW:,C5@=_K6IFDF2Y6(()BEceaV7IV?RWDSF-S?2>
aZUYH-EK<615_8<LafTeLOac>ePK3ML5(bNLNRE[26SGN,.XZX?.X.f?HJ+^J_(^
HSJ_+\86I(COA&>IU\6<<.6XO2M1J;d](=D2?AYA]\?>f<]0)-HF4aaHeaSIf>Q^
TGM,<(U8M@/>\_(13cIac+E2?e-D[60b[E[;+^?[f\IAG.-<DH)@fZPY.UV]+.S.
DR\B<KQ#:[^SMG5K^.b)24NU0RYOeWUR=f)3c<TPLfV1#&/?KPUg;5d6PH?\4A\[
>T@#T90>g]Q6Ag&#3fM70VCVaII5\8A>VKCKL,Sg?4f42XHQUB:@D=ZNP9e9;X/_
;)McK7JK@?AGb8-.?.>)3e/R+M=+^]?B;N8)3^2F4U7;V3)]ZE+[&AL6c,\Z&3>+
V..DV8&M7_5V\L(]H[@?O>c>1;c)bcCaK/?U:\ZE@8]?#JM.I,6f(V+_9NOBg_RF
bHIW5>/1>a()Ocb@FQ,B@N=_)&&aIU1OQ,e,5PDIMVQ8XOK)9Y:]<QGL1O@#HRMM
/76&8GYU0J<WG9C:/fcWP]2c)+.X?a&bT<KY/C\fDK^N5b/,BZEU[\6#HBF[UD8V
AI96.SNR@&:OHG)9@Y6c1TMf@S+.OHe[L/GH2II>5.)?6aZ;1W?CTZ9)U^8^UEg#
[bMF/+9CL[Q-26,cT4QZNTAQ[VQ;6\\@N[g^/T8a?@d2Z3JM174dC[N#,fgP1P6E
L+]X+56OR0[V8I#;++E0OI?U_I4<C(;I:^78/47B,=[5<+aVL=26=.L[(44S3b?d
\U3;&O1Pb[T#Yf23a#RDdJdLSY2B[-A^]OZ&O?.0>]>cU;9&@5A@0a6+.QBWF]1;
S0);L]^-^eMXA4N=_EO7fI=JC4S1;?8VRAVdDLdfK5-0,L?2,.b+A6K.XL7TSaJP
_X[&JU)+^CC62^ZLObJ-<@^e7fU70G2\\gMKPaG<3ZT=XZS>A6(bM^5c3BMfSTF(
e7O.SIKdFDZRKI<Z;3c1ZY,BZ;Y4[#FEGE?K3(W)Xd.g./_Ff@?bIeJ3I>>YV1IR
&Off9b45c:/)^2C?OdA&#36ALH>N_+U[ZW/@7+.L_,SKc)6L]SaO]Gb?:FGWV?bD
\<H,\5;L;LVN]aYU^/(-H>^/ZE=4>3A@_P/99ZNgD/MWWgNDBP_L[C\J=fSU_N:I
;BbTXV>JbA]_&g714HIZJ(VNMY35dN30X[-/O8b/L>2-:?77Xc868VI+L4QOL1.[
PX.5S,e_JMTK<8ZgK<a(<FOW&bKJ9@@01RK?=:&-_W<H@-9BP.RP/XHFG(+E\]6e
5/GJO)ADV6f/&8_L7#0;U;<KF\JD9#);3BKf#F#K]D0SEMI)XOV8\B9RKc)UJAC5
9MU^+(\,V;X?=JdYagXCb.-):AEc2Jc4QHd>?.e=ALY(IbUF]IW42\?BCK^e:@&U
9F)@2K/-c4K7SYg?(0R@\J<;d5SFTCKTf;R6_&R01KTB6_E1f?,a+Jc/X_I>9f;1
O88UO+gCI6I(SLPB.]&R<=g8AU4\U9X@0e-DVVGO.]+Ya5,XEJd-LJI)0Fg<&SRS
LP6EYUW2]EJKV>8eYT]Ha6J\/7+UMY#d-N[/&]SE3@c]b\4FA#deH=RYS(KE1Z_F
[BN)KF7g^(g=dD[0SMKVAe[CXKDF9\0.aLec@3ZY1J_5T)J471YKg#WFIQ-BD5af
A6#62EG;C=/B9-#Y&;P(U?Qa&<:1ULfT@/5FE,-UPMK?7[S=dPA)H26;YP1FEV+4
B-2>)4]@eI;3f\Bg90(;A+SX^P.#?FJ_E=60&Z&D[bbT;.3.CXK6)&26M;Na6g>Q
OO?HGNf@O-#+[^/:\@CQS3.,a7bFUbZ=#QI1[fHdK,+#:@c]U3cb-SM[KS0@-]gI
-8C&54=&#IWO;bAP@C]C9eQNb:+_6S61OMF<O.GE].A=\:g^dQQ2M[We@OWcf7<8
^Qg(cNgXC.:bN4fXNRFPfGdeLUf,(8e33G#X6gPbKGY&RGOcb:,5e<e,AUA?Te?_
?W):@=@.8L:d2Z7M&ddg+P0)3--W.N_e_A=<_=4e/aZENI/QDVZN/FZER8NDVXEV
[VST(_fN_-2:FQ=(dBUR@4LED)HCA[Y7)#J__0G?,gZ+Q)>+d_.D77c;LMOQ2J8M
_:;BWeGQg#4E7PJM&G3Q:&Q4AN0.:U-;;-35[[P9>ge]@&gIIULbI?L6a@AY0H/P
Z8_NJ]7DFIPGBPJOS5aO=dVYI6N;H]MR6JQ#4QO>+e\f?/A;9HS(()B@dN\Z@7^:
BFDJ?:9&2f-_QH1OU<7SJVU9_NS?4L]Z>_<5Xb9B1,aZg:P4IDD3S@c,FJ:V&0C?
NgAaJ)3bX:?\#+F=YcfEHZIQ\[KA5=&.0WLE<4#QGC7U03X[&8BRLW=^N\5b#N7^
)<b_I0;/3cHQ(R9>)DI_111W;gXaM-#8Kg0@3RK&;;OgS<]EgN>T>NYa#bJA7XF&
K=)+c89O19^a&WQ.SFVSWLDZZ7E5eF.J?#9dZUE48R4;/],-?;92c)CFXeAd=;DQ
),S3:GB#G30d=?;O/aOK[66gD&#BcH,7I\AVFR>T]]_3\23_BJ15+/N2Sg5L#>Y#
WZc3P-00(LXb2X+_1dZH/8bM?SO@U(VICgA/1deH4:21D46@5YJ3bAAZ<W;.L9JN
ZXJD+1[Tf[b2[MOf;6K,-P4M>RW,6Td:BIaW+F2=NY9@I-R@FXY2Q6YD<S.M0V<=
0Y/7\+gQK[YE9LEPcY[QOVLS?cdc/79&#F7]^EYC1)d-BJK^G.2E2=eB>C&QAW9I
VT^>afC[E^@Kg&6K7JS(feWEN04YcIN4A+f0fd.B=Q8-8CcdCL/G(P<[dc4g@e(?
R]C=ecING01GdY.OeQRW8c5#MTfQgVEHTIg4JeT20d[XCR[f_^:g0-K_KA_V.E?<
_19aEH1U_RMW)YbdMf4c5B<e91@A=P-_e71AW/.;B15YUV_<-<)9#f,QY_&gPYV1
dJ>,&DA<f+]Nd^>^CR\S71a?SZ#_(Zead-WL_@=FINQb:6g[PC-\1LKN(5EbE(8b
E\?JI8]0LQ#UZO:F]OZ^^4>07HRH52J.2<<85-#Sf./D:4Y@_9\R)B<aa+W&JNE@
@e3H18JK,&&6+TDC474\W@;#[_a)Y>F^POfTJ<:=gT@M+C.g9-NZ[7#Y]\]063KD
75&4;=,D,M.Y&&=DE=&>T2Q1BT-329&=X9/GgKNAUR+5H._eR)LNV]BS6E+HSfeK
0FdUdL&XGMaYV(#59@)^cA1?H2QgJe8(R+[D3259\[5B:_.MM4gOQC;+4535VI.2
S(3@;Q^K>1X_TE1ZA)+@D/[F;ONSJg.F1(a]cRL^\\56\1,L3;0ADXa.gZAI)c?a
Hc/eEHaCJbUA.a?,CUMF<??TBfA&/+P7@Z?4c(L+[]1>-C7E:FB5Jg?:TaI_G,0+
E?Q7/?aHX]gX_3e<8IL#T[C?^)A,V8C.ZGa\D7-R_2,Z3=EYXYJH/1Z07>FTKO9E
?e9_&?3M]ZgX:<2<f<3Kb_;,()@VN0RLDSZ/fUO0LLR-Rfd?AD_gZ@7d;^19_C)9
Z>]6YP?VFGCKeTY_f[R)LMVd1AcS&:M>UN&;Od(\=G-f@1_>T>?FLX._DdOa#UfC
Q]^\SC]gWETJ:2L\+4WR<;cG/YTZF1L[bF+_4[X\Cg1e0ReX=:5WL^DeW/I=S(),
3ZLEB^g#+,A2KAdRP;:7[XJ7K0J@^)b(dI=L#9,I3M98M+P&P+Y;3@N?8.(dE:8>
N_S=MPBOUB-0HFc>G(/O,F<Y\/_HF819Z@X3^25\VS&?<K)\K9,UCD6:N5Ff/>RN
E?ZJG)GSGILY;b7c(DRg,WF[8a^.6KG#:#DSJT8-EeL:e42MP0SM&DdXIQa-SVDE
d.GJ,&fY_,\;TY<Y?8&\6H>FYU-\9?G\WWdP&SKDaeZIT[S4U7^#VgT8O=Y)CaM?
2K/HbH[5)Q7X6=BaCb_eMF]7(6U8:2LcW/ZNCH7a(+Pdcb>?478#LAbEeaL[;,U:
f.a\OE-aZBFPaO=BFZf5bLIK(^I\N0UO82Q+g/;=dTC=.96KFYIQP+M\1Vc=B+EB
#2K^UI23.3.(e6U9[g;5HL45\]eJ(/fD4&g?5IQY5W-#+D#A9M?]\G]^3aIgUF1_
:[./&FbV\cZT9fPc.W2N+.C<837Z;dWR=UP1>9<PUPN/#V<7GC-5PZ?SdX/RF9)@
;fa/NLT)KMN2dWEQGdf(0PJf._LXTMNQ5XQY^cEZQ-C&2@)79#)]CS+8JH5OH(>(
c4LCaX?T0gc(I]#1SeZ0Xbbb28YODYGb:,1cG])MR;ca(e,-9;RPG>JZ?;DG.P8S
_>R2d[S8Ue=_0/@M1a,e.V[+[M3I[8(2c(/M&#69Qc7BC5=02UYHSGGS+-RXc89K
F>ABggRQVWQW81=aIUL[d+?]93[)=NP/-:1Leg.06GH1GT-W/+V_^\@&OM@9T+BT
=f=:)&Sb;>=8H<,VA]?;#Ncd1N6YZ5X-6e@]PNIDVAH2EH@^^8#9=3E.c\5^,3+.
geZ@65HR:N,CA=B0,+:SY>L[J\C@Ma1+0];@A5LVNg8VE1(95).@1@0U(f2YX<K,
MT26)JCJ[QA(f_-XK;)J@5]2VO..1EdANTL/:;cK#FTBF1P<2ScEFfVIGQN?:B88
:M^4[TB0>F;9SAaOI[c4^<,T<L[>4:5gAZRXC0WYcT5U>7>aOKe<d0/fG_.^F36_
7QHF&g:V^fJRGg[0=]..3(1,-QQME991=DLU=H1D4,J[bY\P)<^\;#-^g#QE]eQK
3L8^ZC/\gYS81a.?E]?I4&T#LWQI^1MITQLGf,,?(:A16bZQ]WJ_C8XF2L=Pg9G6
-HR01U1XR[WU@B,M]6AUCM.C+gf5__^e;,7N[]T/fEI[GC:84;4b?:4N8LTg6)PN
fGQJbf&R\3YO6>/UMR4:a82HFC5a^fW_)W0S]Db1A_@7;6gdCDd)Yb?0EbHX90Uf
+K&]cf=N/@PI7F,.0OB;97)/e<I.gW&MW2@Dd;9TZ(4>IT)(SG5b6M(LJ+e?g?@G
D&6S_QZP#P39I=3WHe4.4e.3O?7.6f9ZgV\-/,G]Mg7^GA]f3;_e?-RHWYKd0ULP
7cDGac2,X2gF)e)&FX-Xgc+c1AC(/42P^-<S-@GD0g2^?L3X3E)3#F,RB^TZG/V.
7HZc@(@J1^B[^_d/FU^S5K3QD9T#ADQ69ITX:LCcaTEUNO2(6,LV[daUM>a:f)(<
-DI[\-[N0)d;@11fZASA/]/D80GR[g<1B5D(Xc)OHS47+.XB6N).a^8;A7efe/V:
YO_,1ReScMbEH)IAD3edCL9E.Yc?5:/D(NDT^Lf4S;9Y+UfRRf]TMTfJZ?GFC9/=
S./\/@SQNe6HT^2\8)#^SG<9>E9dFA&1YT/LVd)E^b@@62-@Z[=9-T_9WEaGBFB#
0.+>gX[P>ag[U1/WXE,Dg=]X]Z1L91I04HK21)R-Bg0B?^NG]]BE^H)21)EA^f?.
_/^7_>)gV]b,IVf]@#d@@aYV160FR0f+K&G-6a2^B^@^af;I=<R5P_gUKH&fMCK.
,358d<^0.6#3Mg\Q+P8G_G-G@ULf6,:<47/:V2N7J,8Fd],59a2KX?56F+.8N)\@
@?B7+AH)SeJ9MDX=6[L.(-_C2_KU5<(&Nc3KN=LUB5a0@IRD;:^A:EC9,@RJ?\E_
6B)BG4L#OfF>/U3/\+?G?0;f8gGJcZ#R(95g2P<g+ce/BKK7Z[bTXOEI:N5)N&.e
B<Aeb0\I,B)?cX5@0N&\H.MeZ(N.NJ0f)X?W#JFOEGWHB\4XBED7WTJ@&6(5V1<8
446>d(T3YO:DAG056179RO29QXNBJRJPIFGH54bU6+]bO.1/SO/2a5I^B(2QV><X
F3dYV(c9V6Jf-_><IFXHT)AgSC9DdYSQPe\RQ:B_A(@+L9A_&c:R()]eO/.+(g+T
3^,3c3W6QM)U@WQP7+TTDK=8F_O/FSfL([<SB:AOeD8a(\K<#-\^dUb0L^^<JO-&
-gLcgEO-PM:#NH93.;eTDfc:a]\_]Xa,;0NDI<Y<bV3#0=>/ZDY?-Z4K^MT7OHXf
C\[/L9V[>[^WT4#^DF@EX7FXM68>//bB,NGd1P5fY-VJe:P&-4ISF^,Q#FZ>QY_/
=b/2d;dLYWP4L]^)bLZ)f)?bWaB@-8gYR74A>b/H&<0#QPXRNF#=Ef.+2UOHYaCC
<VI71d=IQEXFI/TYM5(_gYW.f(Q1Q,&G.JW.Y4dU7RB;SVJR@VGeP7A_KG1]^@F7
6ZC._b)-B79BAC&4#TJ6WAS0cFdA+1+?:L;.;49D,B8cgaX>(0;)3E4I6]##)?U=
UH^^@c<EP??8Rd4MK.0YRNX/)&F)d,43J4GDX8IBO5++LY+Q7g=D_F(gAcMbgGLE
E,c&6]DC]5]KH#C.=.)cZZE&N_90QD;PJEPA;&(+:9-LL:5[Q_3a1ZQMSDUFCDe;
P-\bW8C;^VWTT6WX_H2\7EJLA&gH5;749:JV+^.a8H0cQ&CVEYT&d046#/DI0^_-
f8)3M0TL.eO0\G6N6Q(+QN1YC?,&7W7U.Y&b1,(5S9;]05-e9f\#gc(6abL==/3K
&I]bB:[fJ15AW/3^EgG=1,H<-^_Ue?7C2QBcW;;LN]W6Z/HUbA?#3c5W/D(dN6WU
;WO2A;e\]Y?=;<9H57U75I6)fPeQeABY^F,4:/>2eE1d(+(_Lc5&E9?GL#2\(fK&
(U)<Bg)<R1ZZ17Zg&L9=8;Y>01/b.]ed:YbW,=a(JGb?<_^\E&OgPea1@f#/31H:
.]PWC(2FYIeNN+&>C&A;-c>PU-9T>T^#^LeT[IK7<2b<_#0)V&:NPVQ_W+7+4f15
FC7?Q^72M:9Z4CeG[d4++\E>56GE.H-QEfD@FG9DS][R\aPO0?:975GN]TQXE+<g
YV-=W482?F=12[NE.J-cNW.?OGdI9G35)aG;Rc6K1^_KD[Y/OcYf/3XaR\36L13M
>(<cZLY.X^\;G,Z\3J=c5OV>\BGZR>TJZPA__>)YOaaCUXf/8K0SS>I9=XQGe6H=
aSY.;9)7SRe,b8QP-Z90<A9b5U=-ZQ@4/29R,Uc3CL-bIBd-@]cZT8Oe8^C6Aeac
Y\^SY=YT20XS_LS?PPgG.\GEb>W.,67f+c4U6CFGeOELW3_g+65O=3T?#FI2_<RC
HGfC-VYL#^cbaXPYHWKM<Z28:\D-317(>[YR@;NaBF.Zd@1J7eWT8FT/PTCR9#P/
38[Q6)Ic3^5Sf//\&80FG71J58D(NR]BOLa\ERXGZ/gb>GR3>OTL/XL<A#5cEgc^
X5LX18:GYK7;N:P6-8G8T18#EV4:?d:?87gaA/>J5CBPI&)N@Ea4VP]<U_;#2b/=
c=:AMe]1V_VWBJC.e)N^[QB>4_KK\+N2#^Ge8US2a</7:1Y79[J7VGZOaP^dV4O(
[I-<,CL)J,<,>^6@ZR-3;=^\)9&&fIDU#gC06\SWUf(#KZ9PcFU@XbPKB9CTO<1M
^K1gdRC,J=;2;DTH@gJ3Y7;H\2e4\b8X)@XVYdOG_:DC\.(0WFf)62.B_J#0-dEd
HbIgAGNUaDTP-D6=dVML@5dS1[ZH[bKOOHEOc6XK2G6^6/U-5bOP:+ZBOTCH^Q<d
FVO@-HDQb__N5.G<XbRFS2Y.=f2GF,TWdb,N\eeR[H>ETCUSdR]XMZZ&6>QG<d_&
L.VdI#]]44H+D?6LJR1V^N=XB=)=?>B//@YTTO>-TY6)8+Z#P.B^\G,0cSe[_aUd
=[.bOF1LNJeDJZPIaM+UCYM(bdD(:XXZ_eW7YG3gDV6Jb6^WF78:U9,d0:_<^],7
7SYA\_-.X8Z+B8\/^>0M\IU5Y[K/A1P;Ffc^2.IYg7GF)(dPO;I3SR3ERBO_6:Zd
PN4]5M^_CK8/gZPeXNfR))fOBWK&b7fNgcbG[PDSQ8<2cZ-1_S0G\cQS5eA?;dU_
MN53(a)Z0^9a(YDOHR:d>X-&]Q8<]V?cHBGefY)B?/I,?dNOLec]^3V46CIeKCO-
<Z1EN8FO=PX^eCM\3#LEI08TTVY3^d-V5,&>c^U<gHb5/T6MN94@P8([E(W6CZ1Y
PF.#5_?#6AIL@3A=b<=:dQJNWY@?+_JY(T=B9N71CNVQ;1=E>b&RI7La[BVU8L\]
N<G]c8Gb5(0^@c9H8MI;MD:P.DHSDWA#D3\LQ5?W<]J_D;)T1a#P=M-C]860?\Rb
fW@L^R/,FcT5.UH[GJQW;(DD-J;[^bS#]VP;Jf-D[QLHJ/f63DE:7M?D4ULdTccV
QNX>1(/R8](_6GNBcB.R_Q]]54[&&Z6K;Y8@0T;@K[JVT/_ZU4_=6(+NK.[^/df5
I[e(=0g/\?ePS:5Z_O\VXgJZAV#aYa6P5XXK>XZ,fB)HRPWQ1eb+\GYa82QT2Iab
OM[UT8F,[L7e;096+-e4FcT\]DTD(B/D&G=fXC^SE.b8C<A0T9/,M5c.0b-90U5I
.TYP\KdW:Y(.>J)Z-Y>cc+JO<ZV;&3G26J;dPf@@JT5+S\gRL=EP+@@#33Y#F,WZ
6#OdU+IV4G>IVI8?W:dRED2#0Y)]/UYQ_.)H9(RA@VH,AEP+E+2@BH9H:6SMR670
@(F#_ce]Id;F/CFA^aB\+C&C#AL)B?1+Xc[#L&Z>\]THf<(?cN=]gb>DPE9Y3TGI
\2LOWNG+Q_<P]&]eBdRYLEJVa8VV;I36]H&<<g-:Nd\08<dKPSMUcVI#(gSdM49M
20XCP.4Y]f<=5ZVY1.B@@/Y)+9?db);4N>=K<[:A(/2K,Z9=:3<&6Gg?a):cJCRV
RY53(?)<S5EOeVMA+4gG\U-(_?,-Wb)@X/aXO;0IcANZcZA8Fb4@_e]].-.O0:[;
H\07J+(</fJ103cP;dW#39d,KSbFM:UY8K63Z#KL,W2Y[E?\?1^_10;@)7UH-b,b
(4C0dS>5,G&Y#_JOP-=D.5WF3JKQ;dd/H3[;Y0(&FBN?[IV<FA(.a21D4(EZa2A=
Q@20FU_fZ81ZZNQ[gHdS-2H=XSQ06O]eUU5-c(#c_;2XQcPHF_BE3g=UHRN\bV>J
aU9_XZFg1(]N:MK9MT^^aB\HXZK&;#Y7)SG#OKE:;L\YB78/(c/-1U5H[EAR--U]
bc2=g[[1]G)KY)&FF>GKU42_A^@K43^>Qe/&Ca?C:Y7bgA<63fT/O121Y=e\NX/[
7?ZdWQ#5MP?E>;0(6/D[/MR-3/LX0Z-1F?6RdWbe&U@-0UAUN_@PcAI+DU\?:a(P
&TfJb.#\,P\UJe51QBF@GX57CSJVFS=-NDYWXUb\]H48P&(K]-S&)aQH_P#9Z2];
M>aDV.^3?^D?#NASCQ.]3B8@M7Ac)IV?:#e2SEa35ID0Rc+dXTMI\3F@E2O?d00V
f:N7Pd4UB6USA3,]^#YfLTQ5J:\fXLGg+C(;A_9e(5,\5;T8-^f69#PBIWDb?De=
@GfgUI(7T+?=-)A4_W;[PC,b080Z@N9VAXc0GHd</>&?YdQ1&2K,]JROKC9L8[B7
9YY>EQ-WQ#_C4V,U?X[(:ZTN(EJ@a<Qa2Z4<>73JAW;SV-;NT/bQB2UJA;28RN04
c\XQZeM2_R0NeLH74=#g#Y69#6_>LL#P?91#]@SEB8RJ,6:GC@+c-@&,681#FV<D
N2e0_.V-GI,ZYb&ZQ586-fddfUHCN[#]<gXXddaUC@eY@WaV_]D1UHMM;e#>YaV0
?(AGZ&=LALH[-JW4F,7a;@#I+KVI\H9QMbV&Ae,>0HN[F_C1W7Vba,)TdDGTcEc^
V88f@^dbG(+/,O6SXbK(1#])T.9faKdJR>O7afBR&JS-C.2QPVX/=8GQ#Vg&/,TS
X\d3cBCU\9G_0+[9/cQD<(<KVbY&/_V_AGUV#P)H61U?LW#?QF,^H<M2#+@[5S;f
:15^ZUY&a/d<85Z+<(L0Ub5\,K,/G?5fIZA17c,ENOWER](9-_d<RQF04TP/-F&+
F+LE?^@+5PAL3,fAXM@HQ=0N1=g4];N1g:EJOOFDFVIc?OCe>HEHNc)SP9cNg(..
/_8(9E61(7B#+2A>]9M3[?B@VK/8c6fW\HU9&//RPaL8LCd\O>G?0E@X]AId#c)7
:X8ZFQRSFX2X6\e4)e9d,:c\@gC,L0DET,#^&b,_>D,MO0(@V_7.5GZPODKaGd0&
UMM(BWbB6CA0JIJ=9?4?Ve5e2]^T3)D1<ATVe+]?H[65E_d\A2(&1DCb8eKB#TDP
YM612)C?3G)\MMQf7>HgDbgN[B1FUGL4&@Z7PG<E>6HWPN3^..WFG;C?f</B5e<R
PXZ.WGfYa:@4N0F]5e)E[D<M_8O5)ZN^JE1WA625e1J8)/:I)3^?f24?41d6^Z?\
7C34UEI4HHKVA[KC8gaZNXTaBBQ6EP+[fBY3bCE\\K5P#YcXW7G?98b;f=_-Ac@J
,:d&g+2-gHHB_,)QST-B9-ecC:dH+:#PF/7VAe]TB4.bW6e5#,E<U#P,]\[b#2gJ
)UEa&<&>/@Y>4DGBI4BAFXPK?Y#_@,P3S3RS>.4PO&Q04+LW3:K>N6U7.XE,g-HJ
N\<Ha2>3gZDAf3>c?3a5ZUAX6_8DB).#4TPSQGIT;VbD\K>^6GUSZ2NKH->+&6CO
#;60V^;9Vd]YEAML=7CG;VB,^(;V0[,X462?KP+87IC)&51-H:KAM=?Wf>>,fL-5
U.PSV1^BcY7>Y)@;17DCMc.5J86(GL@6\M\;23WST^ZFD&)7-CBd5cN/IL4QE6YH
T0B/XIX#MC;5?2]5ZZR#a9AVFa<+e?J][L+B:U,C+LD<IPX>Z.bJf#?a@&0MPD-^
H?D(9H[[V_FAMZE<fC,-a2+ec_J^P7f+eE,_\3^KI9:;[W>MQF[.ABZVEB8gMEVU
4dM..d@N35OW@@JF.0^Xb)Bd+Fa\L^0RQ6SNEYN6MLd+5-(WE++\//f9U70QNdPc
3H?43a?aN0V00@2_UY\6W<D#PAZ0>SF[aWAb:AaQYH<5Y7D-LH_(,G][J6-P?PMZ
PRVL]86TT9(K[R_9@-\F>cb0<:KCF.]Z/5-@4BK,10\6&#Y_f[\aKYf3PAEV0D8:
TTQ<SF<]Wc:[;gI?N1I0V77=6O^Q(\RM2L-d;V--BB,:N#:>.gV;F\g<[ZE?c?YQ
-0Q]&K#J7Y0EZdef)c9AR\\)83BR.b5+U>,-(,+BSL6)<VU:f8HBHg=FTS2TRg.d
-=8.V\L0Q-LJ:3=4,A=L7a5DZMG>9B325XM#O1@\eX^Z./V?J^K[>F5Y.:^c11#T
0&fZ1=E5e[YecZ5W>#O85\QD[ENX8#g.>E1O6@f+F>+)V.6C_37.PY\-01c3,GZD
TE1[F95DQ)V5E(.gWFOb(D,)BY/V2\)8<-)NF#cdc)Vb+bIdQa51,,6PQ??=\4cI
<b=M]V-@WdbG,47FXIfHK>#PZ?)9E0.J4LW>+7[f?S0Dg-MY,Z2RU64,dIYH)B2K
aWO\FZRaE-^I26<:PN,RT=9-H7]IgfZ3R5:U.(Y5.Dg9KR@J_09aXQJ=M^H4P0F<
f-?3:e8H=LH0:HPE5_YMHOM694e=MTQNC5S@>7R4B^>\:8V75I,X;Q:_#O_^aM@/
S5688PBBEf6OG/.6Q3NJPeKb;a^G8R]bB7)Rd_>=Mf\:&KED,W&++D:X:IDJaFTA
D8>)+gX@SGVNT0\gYR1g9\X26]f[T?#[g<Zb8IfX8Kcc;#aRGDY5,=_aO2<5b6I<
&@C[(W&Q:2/RR3+27E9C[.2G[+2\#eXK:STf=0^\VNIA[8Z/:4f@cSfd\F)YY,</
:IQbJ)=Z;Z4OH4X+-,UO/TPBYIDG<.81K@X<=YBf;g[9Y>^&P/14UHP45XBA\V:K
^3SZ/,T6cI3U2R?<N=J9ZE_I/:AT7N;g@RP/65(C40661XgJ\@DNKQ2[5>OH7[aB
_cD/OT..F=bOgW/BW8RZgGG[5Z<?_S+KU=AZ.X29fL\-#[DDdW-KgC;d[g_f]3YF
[TZ<<]TI<d65##c^494H;GTER^5aZ5KO:ggabGAY7X#fG)V009Dg:Yd>X&Y/CY8F
>+7dPc4\#(RW0<DWBWKJ5K6Q+IV+PX[\A\gK\Pb70//g.WgHgFIKXJ_K\1,104P&
B#X;a68(QCLGE<WcXMD173<,1BWYW,:C-C[]\X)F1/9@TV&T]5::U5302g8bI26K
>bB:;S@@O:bS?+HaZ@:X>)^0>01-0O4(J?M9,EdPSHL42/WG=]^gBKL))c@E@X:[
b35QI?[a=WS)-+/3G:XO.9ET(<#YP0WZ:8;f\D3VSTdEf9XI>#.[-]ER+3TQM+C,
0[<>87N3<(S?BeC<ZN0#K]BL\ZSUXG/&,N-/BU-:=6A6.d:R2^-TN(I<:FRLQJ)@
Wg<W;E+VMLJ4S.@/_=Rd_P\5LO3R<9]:GI:CO/I8FU-eC3^E/9)H^PD-Wf_(HfTY
04M^;K6?/:&Y.90-N55:-\<L+Pb9)<Tb83P#KKP?K/;(dVS[^\A8<A9d]4RT_0H&
3(2->bEFDG#g-JRH&B56B8.UH3-MZ1XcK9FaVbO(?(>cQDf-<4QU4K:\Ke-+2d<+
:7f2//T]b)-O\:(67[WE7^8E6ZC0]Z>HKK04fMbH,fDSCI7,RXKdAY5be>@JfX==
5Ie1JJ75eNWDF\Z5SE9IGG-4fZ]QY1CRf7^gXS2BRGZ._#OgG-S[C8d8DPROKJg<
1MG/+1G>X0g8Oc)F[-]Lbb;VBO,<H8B)G/+XNQTX+R32d8_P&_C0+\VBOME7B<Q0
2=8CfW62efYCC#8JfWKfLU,6>eOOGX\0[R0D<\;Fe]JSP/-ALPMX[A3@I)R][YE?
fWC;(_2d7ZZ6;YB,/7\BSLeUKL9H2dK51)Y7I_-<:\H7O&:eR<6=?#WQ9T6)eM]W
/>OCI)A<N?XP1A5)_G+>NE9F#:P,Z-gK3Z-BG\GCc:95b:8HeY@BG9,5(g(6>E=B
NEA5<cbB+_RG&;_C-)VMJ;??)+ES:7\1bACf)430_OHJ?&e&U(_B/0Od7OB;C[K6
-ZV&GB?+ML+?0S9)ST<NUSW(.-M]APA791WP_9[c\2DQ6U/6=PYZfgIWbg#:2H\^
TI3?J@IQ,8\YJeY&_NRM8B9GN]P#JVX-[POR+DeR@+DTG#)2SVHc5bff<0(7Kf)/
H7P03MM=0eS]dEL@-GB9LF=Jf37aGW@EM^R5PZX/NX97F@?C)7^Z+=)<.2F05.Q<
aJ45.?3Q:da3>&>C^#?SGXZ\\0AR<5<<)SgX[RBYK>=)T&8&),1#>76MAEL>_/DN
bg_@bd522-INCN\D//-T@ZaUa7K,G=5PQR=7-Dg?dJ>MC;G(<L=M5RMGGZC7<eCH
eJ5-XDg)JTPHTA/cWZc<=+ffJC2/AMcO^.^0GZYUU;M#+=A:I\N\L.2D>O>L]>9a
51.Y;J+8&db)g;_ASK4?D1X_70MQRX4^<cX0g8&Y.cMW<B(J.3^X&W\LB0<HNF^_
Hg>7Z)Z-EFP]gO::5K/YaD(dL?=UJVf,HG@AgfS(47ZTUbS0;8VF856>NN]7Ca?C
<^22P-dLM_0WVdNZX-e.@SWO\@:/C743cS0)D/BU8\ZY34ALBMA8N/W9f^[O<7/W
\MX0aIS<(g[\A<((e22Ae8<H</015ELQ7?./J(dF8dVC[E237]ZBH^90<UW+9R)E
[65PL>+;fYDGAL?a^GY\H4[JO@:-a)N0c<EK]-YN@.cQJea<]7HQaRAA_T&\5NHQ
[Ob;MC7?B=ZL\5(bR7A(Q;C]aaO#(Md((Z2eATO4];)XA&\@4gW#3d)&[HXVE^BP
9g0K<a[9AF4@_BZXOX+VZIH0.a1X)..,TMRe,GK2@@RUGR[.,aB=N,RJ\4Y8K\/2
X-V92fEcKd])Nfg:#.9+]X)3aR?eFNLLN3KNS_:AC,=/Ob2N<;8\\YB&N_))<(R+
KN45FJOG\#a/5W)RUAK\NHL63B2QYM3e?OTP4aU?4^+7F=-S>6\KV5WX:C@,Ha:8
KM1]>Pd?]95_bVF.=.;8ZG#7//?dED\G^0b_+UEOLZAQY;,:WOD/G_VUZIEN,LVf
4RSHNfLI_=L2dY^cE:1:PEd99dW\:5:.L&D-bLN1Og1TdO@_U>_4[O58GA2Pd=6&
_O1bWS8F-d/(Y/V6cB1,^RcLdF>DVL],af_bU.[Q<XP:L^]D#OO:7HL-_3USa_f#
@.,Eg,]AG)QH;20PJaBCT=8C/<dA[g=)SW1W+R0<Q<1JV_\7EN>HFL<PJ30JA,eW
R@Wa+BJIS)L#><MTG7>P-dZ90A#TH/&-J;G\=S>6Ed]&PD.Y[b2:J3P)[T\=P7NV
_F.4X\+H@Xb(0,5I]QUa@2P^\/P>V_/3cF^VKJB7HZOJZ1](\7f7QdW4</J_-JQ3
VQ0S=c#Yg#R,MZXC]>-N5O]E?dF<NQ_>e/#E#CgZ=JJLC_0W<)-YdM5Q#R]fLbUV
9_YB5eTE56:K,5/PNGN1D6C7/+f\:-NEA=0N(A;N_Gg^/37F:@f7WFEMEUWMM_FO
@1@@4gHNa[E,OCZ=g)(&J73:3eV/\Ec95c-dH::4RJfF4K9&/0H&?E?VRXCdX\g[
,8/33T7;JXMI;G:3Ug^-dKQ0Xf(I)+Z0aKf@6d?Qg&GBRDMd^U9QXga8VdBXIWUU
RZ];\HQWe^FXWVY[P:BYC>gTVEH:52d0V?DK,=(Q5AT(VdH:LETGHU2LgUXNGIHc
P+2?XF[JFBTW>]4JW1N-;M1TeEbQ.EW&TJ[A7A.,?=.FW.?\TUS^4QJH8D300#fT
W\BLSbINfBB&^C[>&#IL#L;84=[C7/W8MGEf1<b+6>UN+#0NJ;)82Ib[Ad?6I&8d
@e19@OY,WHYcNQWX];?8KdXY]<^f/AU/Jb-K6-O-WIe_W&R30XMF@WZ8><M_WV(Z
?4-9L_PL=HM>2B]]4.?#=1T\GTF8B:1[JfD,5f.&Ub[TEC<5g6J7RO=P?JI:;LWa
\6)fM8S.d&aEB_aG6X]IRaRZZV:bI6c;c^d\ZUZUFaNS3_P0?25T)f(8d\#]f<0A
FN1U#6SX#-f<Z/gWFE_#Ia@#ZFfcd9^aBdVMMG<S;+:OAB^#Ad-fK(feLI,+N5WP
=;[#,R#3@G8d,_E./<7(ISa9[TV,YZ^=:SQDQ(?D6+eT_5Y.-EEZB+6,gg:KOY;W
+\,.If1J/,6]U=egFQRF\V(N.G/(g>0VS23CA4GL]UQaO@/S,g8ARb(IPH&7P04]
6MFS3/OaQ)TFgWdCJ\Z9&>Z;4f9V4YgJMCb:.)@>92A#Y\R_+MU3M/be>,&@\6T&
G\f-[W\E]^M0TG9+4Z?YNVFODLa3geV3B]6OfD&@NN6K.<C]F0.MWAYFNK<_9EK>
#V/:=KB-X3C#H5fJ7eW8.)1Z(U1=Z(4/bCM54L^7fRT5RR?\#0fJHRg(VL-9QLRd
Ye<Qd^=b_Z4&bfL6HL\EAB]1IXG-&#V20Y1c?4H#O]F]0BK5_(:3]B<OK^_gAO>B
>XeFP#CW@^E=F+Q\Cb@VCg]<S2=<PF,gId+/c/gN3@@@&Z.Ic]H.QaE>T2@-C8Me
^Q4I4afO&a0P<]3dDcVa60f;(DO9:<9SH^=V/<1&GHYQRY/:e;]/=EV5(7Vf<VNU
T+f[Q4&:eDGJCD&3.:)aI^Ff;8]#/0&:;=0>E0]#/b8GDOHQ5).C7Q1\^;a-ebP5
1PR1OY9KUBc(MeJ9d>)=.T&W4H^DHCWef4S82)^-?4#2T)EM<T8.WREH_[]fE),I
dgH[W]X2_@TBQ<BNOc,5GP<\Q054YA6@6Yb^G;2=-<_5WJ[Y:14HC>cg>H^U&VMA
X_AR&:6P=/^_)b:C^04?(]5G=cFe8&MOK^4Ffb\d[BY,PU&94cb^T&4CZ[\RJYe=
N.[fJdVg,;?^a3fS-GV_L.UU^/HNU8_;RI#2aB6Q>VcKYbQ\M#/D\I@&U:Q?.HN6
0>MI\+,Y7ZK/Y6:&fF;D2YAVIO)#<YI8IB4VJP+;WF32E_EF9^-cUcd,AIM#;=eJ
W[5-]B[?<TNDJ_T.gB(^,D#2<H?:UV<DZXQ8;E_JYR=6[FYR61UH(3EJ36A[2M7@
ENfgDbgLe+J\Y)3L)-cU)A,=d-E?[?9,_MXM;ZI_5O^0N67IUL[K)[TU/OT7ZRCT
9WLcU+N5OMfW-<NQ?+T3E/eCTYUTe9gU[K>)6:eED.7cY;Z.@?6N9;E+7+C35EIN
\<2-I3S]ZYa_N#f<V733U\:.F)F9+]OX6gRO;9RMU8?Q39TaDGHP(9BI[#CR+T\Y
BW]4>6QVDEKSK?:Z:ABNXg^KDGH<W5O(B93#&IggN3V7^ALf>=(eRRS&HRRb5.PZ
:-7BFe(;gU,Waa-_-[dH8V&]MZ9W/H?6f_A&1^WcOPX8V(?>9LKS<,E..YH/@1\/
G]=+G+VaK77+ECBD?1a4</VZGX<F(;g_.G(7[#AR-/L-QVW(RH?9gPS3FNfOI8=K
>)C0&@?:J4OE7M]F^DF[4A:2;N0>ZMZ:P1J230)<6>2LR=]d9U\\ba<ZHCGeM:VT
POJ2cLTMb.WUa#^Zd:M8ag0Jb82FBe(D0]7G-+Y3Dd1.0gbASL++=Hg-e-H/^]1N
d#ZNS8=THVgFB7M.:d#75,30I2#_fdFJ]YGZ9\21BN\HX[OQ8SQeP=VMdU;g#31;
:e<Z9Y64)W@0(646Z;@L&@,]YEYFe3,<0BB(,39@[._XK,:0B8F_GZ2T[1S<Oe>X
ffXaERB#I.HQaK6G)5X(#<YQ+^K(QfV_@ATV=>\G.D:W<#8]B(@/VG-5S[ZITB+W
AP(YK>5--fA\e8/&1]beHAPG=<:Kb)A7TaX<^XAF^c^_(D@Y5\K8D@,H8d32[JOb
E]B37OBGS,a19X]-cD/S=1fCOd]P3b1gYZFARLM/39O#8=CS@U\XN+WYA<L?g2Gd
^KK5XU@M/-@c\(3LfHgXBLZ:UgI.9:Y;be/)-?25T9.IY)TWRR?;S0KWcIU5/Q,1
DgGBB:(cb\@H=88#?[:fLT<K:FD3@]3==C;5=FPD.NTbB^(eHKL,\Vb2).QLTFXf
^L-;OOZfd-M?-68F4fK6T?6QX,S#I5QA&OYO:>KfX,^cf^BD:=]G_X@>7&IaGV#<
^d4J+f4K1]4<(F6[0:L8XfWD5[81[KO>4A-8@R>9]&=A>-P1&>d>\Gg_)HP/C:/0
B&_C_V<</ga6/<W2E:QYbK]B.KDLU58JacU^PV=b,dHC02=I)MPC/)768]J=XRU]
MK3EX1NNI5+SB3UP:MVdAdNE@4SVH7#6#PGK8b@Q+XZJ4(.9=C=.?BEN=H+U47;S
6a[:eJM0Y^KKEfb-Ig+Y:^5AQO^1F3S3^b)fcR(5d[cIf+.KW5L#^d.dHT/3:I)V
gNX-=/M9K\a#/L4MADE90\@3\8K07JeeLLP5c&MBH=Y)B0]G>,/Ddc<dH50=\.c,
[DP?fU:7.Tg9Ue9?N.IW]b.J22<21CNE&d,\YQGZ>/d#&7Nd4-HOL:T?HR:gg[fK
;WL3VQLR@W89R(B1V7=4<T-?aH[KU5=2M9M(+WFSL63W:#T6&&Le&L;HBd-c[V@K
&M(,IcNG4ZHWd&GH,E1E0)F0eU(Y19D;=6R4\Z9b=^BfZ_,-:VDb2fDSQQTH/OHe
D7=_V7Z,+W;RTL.I7UUO)93I2#1WGLBS40V+&G(+=J)7U:7LDf?1FWO9]&?W,DGN
@3ef_ME3MJU-e#]e>SC/PU<6;8>-g^.C2@E,VIU4-)O7#aQ=^N49Z#J6D\FT/2QO
[+QWLP:aH8e,M;7E&;+B<WZ^S=N#IXaQ-X@#AN61(8fROEACb/>aAbKRgd)S4If(
(\G,I^1JTA(1:BZD8g0SVJ3KXZX;3ab#U]DZNHS6<&Ae7>(1(;N:cQ+Db<1+GZSI
:Jaa9?1.<a&bKGK2NTJM2f6d&d@=N<:,9)XBgCI\\N_EUKR9MM#I:_;EK.H86>&C
97<@Y]MC==/70R>K-G6Xf-E+WC#0\5S)O=&-@>C>AOFQ3f9[K]E42NCJ4DR)4[BP
U435J,8WK2L;X=JKZ&FGUM9.Re2?UF@G--d1/MQ:SK>&cHEAcW\.0Mg8&[:6/&D.
.3HKI#\25RN^QVTW2Y-Rb;>@>++F[\]_@b0ZC\.KH:Fc\[WSMN/I(5a)L1LePgfA
NN&129:B6&aFA.ZAU>7#5JC/@,5A#1\N<)IBa_N:><X@08Z_e_+O?ON.#Wf;#6K=
]:RX3-Af95OF].<TW]TeI)g8b6#KdHKX/.>Df??Td_6^0TbeD0_XZV#?aITS1+L&
7,ITc]=RE@d/^P(#)R8D3ZH9KcaGO]^9T,B@INZ=AJcf95R6U[1NAV3MMLKMR99_
-(T.LN7C@))@;U7eEMWHKV<aWWg?>\<7I3G.O#/<]3)_;Mf(04;YWBWRJcE9]VcA
J]CC4eT4=?He0&>@B7SE<RHFLU_V;FNFa,2G9ZO7QLL=^D.d#Y@<,B3(=_KAcX@^
V6\&c?<I9.2)DC[H6e3H7[H(,UCXA@:N.=..EV/UV;;Na\NZU\S->Ea8;0BYB3SZ
,E7V:&^]GNZ;-B.:\.;?<NF9[+,PZcA:YFa[Ce0H<c>J1<YEePO8\c?d?CLRI98d
g8L:GR;S?93bA&2BGaOXU<8TL>:;,0d:g#=Ig,OA_R;2EUGW\X(M;\4M#M4B[DUB
gJ;gQd_1fM&D?-5X]?cMYG/b5ZA,_f[(5MF?Y&?eDO/WPY0IHEaKH07dNJ#WMCd0
X38Y]SR0\VSIA7.dQa=[Af0efD9C&[]RDW:7-R#GSXRYb/OJ-Q4YBa.CG)Z#-E]2
TbU<^V5f1J@KEOB6_Z,G.52BH_WX;<B/:OQ:W;f9HFCD6RYH+JZ+FG^+2EY]=76W
bN>UPXVTY8gSNgMU.X-)SGc4PB)\<+D4K)=fP9]YN[XEW_2T?MM?67;KRT+/K:GB
&b-1K.^d.AZS1^M:[E9,=F1-g?26CE)O0@H6Ea4G4TG[]GF3YGN5\gQ90cL+f&a1
TEYFBJW<./,S\P0(cS8ZGDY<GIJGU<[fI;@ae9/gO2L-X?=.MUa/[X]VLeOJR0g:
[P(9@egRXZ9[@9JMTUECD#_YGA@FACeI+(/P_91Y7?aP,BO=0LUF#c@4:3OGNQOF
1g#@4-39Wa#D,WZK+/Z54Z+/\Z)_g0UYQ2>=)FLPAc?30UF/0<YIHc=8[O5\>).4
LQ8JFIRR[WJg4Pf##A8:2I;SK@b(PND8f7=FMYCIE(c.IR6UgB\R=ZLRSTIFZTOc
7:]J\.(1HeK2GIK/Q1(2eTDI>e&VSW^M11-7>_&Tb=?<5T@NLQ4<c2DUXDc4]Z@;
BBfC:O\cN@G2+:==acAdRdJ0N?DCC(6U@[g23YM0IV7JZ>&,T3B9YYI+8+8DfZfS
e3f3da17JbgXSR;?W=L/@PefZRT[-J)dFLY@T6@\[C.9aB?J:<1LcET0/I6:?OWc
P[a@0Jc\,L3J^GI.ASRFM-_89B^Ka675JPDb?=a/aQE_L2BADY-YGT=ZIWCeV(.<
-/af<4ADD_1RSUD]eT/DZ(9B,K4ge>,:;?M7=S^_?#a4T&2/_K7cEa)F&G4>g&\A
2=g=-E76O3KF-DJaUPP1f-YZEZU,d?+b3P30/NJCJca-ILF/JLO<>7U(C2P-3CJN
^X4WMME.,E?a<e@2&+=,YRGF7J=@UX_g3g]cS:A9c+M/_cTd9+eX(2@WEVTOL1<2
75BD\T^RdcN?6(=1GbISJPSVD3\eV9EddV[R\1XcWd&T_>[]=\\@88d[PGAIAZUc
?deD^P1J;a;HR(&.f?b\BHWIUCKRN2SR]P<0GeFd6D?\ZS<9AC<adgb&>.@09JcX
c(eeZA-fY-4IFW4PV?^\E6cR>g/(#WC2Q7SE_)>/aV7g9XaM.>^Bd+R5^d1D:dQf
,M.1ZCbe+,B??7UBfgJ/+?bO.^[-9B5a_;\D8Y=f/L^S<R<FE,J,FTQ@1=SCLKKO
101=c8b7dSBW&ZV4W#bg((@g]#Yf1eCXZ8A</WYS+1>J8+/A7FR1H]CP2;D/>G>(
Q2Xg&1R<3B^<KaX<cOI[<ec(SO8/PL9#_0<;[MAP5BS,->Vg7\^M,1L8Z[_.-OE;
2E0.+/=C.?PXGEOGC[N,>YY3Db/N5-\ZY1@cCaV0+FP@/N-U^+-C0F)U)#>Ve6D)
8=@Dd/V1GZfWX0DW5]b^e>JaB_Q9X?@<F[B14#.Nd=AT]7KF@d6b+N@a2,0A3+.-
ZC</R9N2BH@P][#>O#._1<(E7W],P<274B6?D[6:YQ.5DB;@@NCE[&TPa>?VgGa?
ZNZCe4dWdAfBH81DV8&,7H-Z/D-fI=\CEP]T<V#>E0&]_P0#YPH>aJ&?GSGKK,AC
_P./=S:9D^]@Mf^BA#AHYQb5Ba+fYCec&ZH=GMN@Y?gR1MK,4#B8/<gaFWCAYfaS
#,4WVg/.2O@YG_0>3b;;F\MB^34V(]VYNAV7LgO9\,R-LN&W(PL^J63?@e^9.K9E
D2E8WQ[YD-#X//OB0GTS]R18&E8dUbKIS/N&D[3;NM^KdI[4NWaJTdO-d(CE?P;d
[E0]>S_1CJF9Xg^5MdK>CZaOX:-QWE_19.BJHF]WG914U[>O:8:Y0?O)N[4,CKJJ
ZNK@e5:E\76Ud#QN:AE,YP=DJH8.>Q9;8>DO=1XeBQ9F4c?8[IDFY@e3+)IS0DQ(
?##W8cD8N]8MUO[S0>T<T/a1BS\C.4TQA(=OO_#@dE3&5V>2QgYM2+REJ6BE+XF[
Yc3&03@P-5E2R_P(FBcS5+dbHE>Cc#MKe6J[;G]1KWA]>\gI^=VG&5+cKfaMHIDD
E<Bg].E@)(Tf/UM&a&#ZA,3.PS??=RT:/5L^XeHbPC3J/=cU<5]YT[HYf#dURO4,
1dDO@3QY>:?K>/EZW8=b)_fJfaVb7N<)XDb]V57-e:@BW#c2QK84BU4-<H92==1C
6TODF4Pg6,CQ[Y]ddKCK3B&JIJ]YSZO7:\B+^#<U9A;\&3(TD0II68IS@XN2\ERd
HL_bbT5]@UIXQ9E9ef#9)8QYc=O8A9cG-M=A^A;a14355QI+9Pd=Z:f,[C0/L7bM
QUb8<E>^F<-#SLX>ZXcA5a._8K>>&,LBT>2-F[[D1eE:M\\J=N@MGd[7\&a3QLL<
8<eN;(.VS2.C^bB@JRB,ESN68aR8(BZdQ?].0Z-6_XNU?,6#cGAI/2JG)9Pf5+&>
39N8We0SSdISK2+g@G91H^2PLeQN;3OSBZ<,)44@[(+Ac&LaTcMG.)[&(#7];I)A
J&829/7[RTcdNe<^52^>NGPe0Z#]SW_&J@Q2.a4[EW=E=S@TA1C?,B1LV=KQ(DXJ
W)OS;6B87RIcg+.4G;&[RX)]Qa4/2/H=H]76UW>C),-SNU^.^Yf-O>S(_E=(BKK7
>]_O(-.5D\#\=cd&?;I8:-\TWeRMGXP^L86c/)0H@(#:^J,3aY8e:7\;P/?<MLL_
/,4M\IW8HL3?@#VMQ<7YE/^18ZDPf,&Bf)W:157=^6BBgd.8Z;+-ed(;9@MOgJKb
5KZ[)YWWa:c#V1@[-:_cL4b?LeXLOMeA)IB/OQ_Q.RH<1&X4\HE@LCPG<SCVLEMQ
KARYYYe-@cT6_CD0<dRF:K(0LI.cB6NP3F05;6V6g1Bb[^X+c?5b-K><f1VGBSRU
>VBM5[g]aXSZ2^CIWLS+=5O3?FZ._EfM4:2bOXVY1NSB-B2AW4gT@If5R)5,7_(O
O&5>5P9E];58\)W4#WaG-</eYTK)?@:DgQ:)\\48SZd#d>A)M1H(U0/SDX>JURE?
eF=g)+6:/#6S^9SG]^dJ5G6Z9V[6Z<]\>aU-UKgEMDZ58D,MW-eH=M3_M\VgX;Z=
.Q;&[gS^F8:WKc>?A8XFTG4H^acgcDUW\+2BP<ERCF)+UL<(SAc7Cc&ZT6:b:=>S
S,)/7F=@TUe3-.\gOLFI7aS1[--b6=<+I<2G57./6MWYFbK_O&8QTA:E(?1_R^eL
9FS@g<X&J\NOf8&7+@BZ0\11HV:3^f9P3e5^cY+g.#T>.I77R^cC+O+BIQ[@+<8.
KJ9L8E5Y,O4#VOf-/E75fT,c&:)<Y),+D:+2CW6E#ZAV32O/M@;4Y68D-9GUA-WL
C,^31RBI<.QccJD8\7XBg3fAC15U(M<Uc973^\e:6&&LI,#fT,YbGNc;IB84?4@5
>]1D&7Z^G,dMC#6dZS3>2)7f)O@],71FRSNB4G)=22D)FKA\OF317@7=NaP\eW3a
RNB#36-C5a#D5(bEL(D<QE6_gN?aZ0Y7,VR<ba-2PH#?@@B-J(EB4Qd&SF<_#1/F
HU?Y+93U^FK)c^=7ZA[TfbZ41:Tf>I1[gfDDS3,WFfSLH<96:5740&F2\UWV^1\H
;/=Q?JX96;6(DK,<<c+CKU#e<TKf2[L6;\VW[B4Ag9^N+c[?((8V)J.8:O><Z_.a
\\0_:5&.Vd2QNPOE7:aV@,4EfPAF#4:aBfWK:,TIUE.L#^eVG^9:cbM<gdTIF1C>
aD=+2MMMDW#-<HQF:\CdV6<VG7-UP7ZYFIb/QY16PWD81,IBV:gMT@UMCMG=U8T0
#YIS]>[>910C\]g0HO>(+[,HZacRSQMc\<2GRca:T>f_)EYbS/=8Ig6\WP]U:.OT
36TQD>42<[#(/)O:HIE?:;d&63>,X<C0^P1fN87+c,D8_>)<d(J6QQ/Z9]c:71AN
.;9D=^6@\N/^)91:61J:0d6O7bHWH@LA/T]GXX0WM.A/N6<9AaHMNVV#9D+JJV:)
\SL;6WK1:X+M19P[CD,C=-R1c8K.ZWTNUX#.EQX^67-K#-M:<^=;3Acc1e\YU)0P
cR;7W>Q/)\/Q&^,UTe-5SB/@T1;_HY/M_VLG8;Pe(?E?1g.-G\(FG4eF^;)WQ[&K
SAIY/\-(V#2SN9R6<DIf>1)fNIFPA+f2gIeL+M6<3[0MA;+VB[g-.9)Qa[AU3\13
3@BDB:Q=;(<QB?T?Y,ad:-\XcTQTG8)>XQ+./D=I3@gYYZB?/6M;LZXTYS&gP[WV
a/06?XXJ1fP4ZW10AXFCJ#0GTKMN(=(cW18OX4MOVJ;LF;HR9(U2O\=D?U1c]@4b
C:/40:;g4@>KgB?.O,PR/H&C_=Y;aTaTSBCf7^#T6FQL:(;<JLK;O//bY0HHbM7H
<R99/U^\SZb7C&Qg.-?b[EM[(ATY.b&9F<O>^L5S:AOLGUB0R>PFdK1Dd_CU8JaF
/JSDG+2+;WMfI:UIQ+1JHP3A/Md6Qdcd9f@27c<(HVA&>1\e)\9:M@E,W_.)3[gT
g#F298d9e@=)+^aI1U+8HcIMJ=NPJZ5L&8eg#1RcFI]dVI5a3WWSZ<cS1,\VG?.^
US#\1fgGPA.H(#X]ABG12SY@<]>>=UYeeFOf0&KU]@Gd;H;Y0R5L8[9\7,d.;VFZ
M0,/YCRO4KX9#=9a2]Sc]5B.=Z[<6GK3&=(_bHVBI\O=R?B-WX8)4+&1X(WKWF7V
cX#:(=0E79T:dCd:][NSF3G[&?A\5TT]<A?Q&]bJ2)J6,aWda@a_+(,-642K[[IC
]DC2]T@D\[94)5cFDZ&6AM>H+1&D.K]2;KeO&edL46JIEUY<(<fNUO#WCHCY.>57
f>HD=3C,RQ]RHAU<EUFJ^)fU1]6MI+&UE-TZRC/E9g.QD?,8cg_1PY@EA@C7Z2+]
(X>1Va)L<_gZ[_BK][\2.SSF33Y5ANFa/QaJHU-8C-K&dU)GF/8=_W]2D^>8Vg>_
@K]abY9bJ[Jb+NXAAP+E]R<J<VfA[XP8cPJEf8aQ6Kd890dZ6F]X@cHE[&H6FKTY
eNHb>[Hdf]B\e^c?B:ES(N,)\U6E,LYUf/,])F;b+4J9B3N?27S,N0F3(T5+MJ[_
OBWB@J5[NYR0eP5aL0WRW1\4)-c70W=JbZa45QHT71EMDfSVY9gG)CgG>;Uf]>(^
[2(Nc:4B<6e:Z?@T9^:Z@-Z@Nb<3Pc^&Q59P19122:2Y@,NIfdMKcd82]^]#HCX(
/#S[7Pd#.)3aO/36^VMeZY/]#Z;V9b[HS,,@B+R>e]D<b5=#0U,Y,/A1+TBE;3g(
KX=AF?=V3AL46#)5#_(BOeJ2TQ<(LT&B\.RPc++.93HIYDb;A+WID(7_(N^CX,#>
_&-c[9Z[A2XTL7-A0fOeb.DSbG.X>&=SARMM42<LBPP7BTUd16GDJ@f,OL&M7JL^
AV]XK>&J2SE0#c<\UW7S@PfD5Y@2LP&HAM_DD4@O:Bc-@0^f<3fC1)ZW@K<PGNAa
]KQX7T,?J[AZO\(2Gd-[?8GXUF@)dFS-O6LRG8@gd^.S\1;OI,d,YIgS>/.JRf1D
Q3JY3^;(eND/X2,D.K5)JBAC8DF_N.YQZFD1Q&I];6(?J_L:EUEIf7I)/;[]>(U6
)Q>F3eGVOZ@H^OWB8NUJ_;:CbQGEGE-2WK1=^SdNM&M,_aTJFC.CAMV>GW@F/M]6
=33IE_F/C-IYVXc_ZO9e1\Mb3STBKDYG[<7Se@P[PD]^OUIGZb:IX07b-AEU_aEB
e9BDWG(TP2XV<@8M?JDgeG4JR)A6H21_+^SSc,P\S\459OWAE&f\GGg]6852cY#S
(CKK4=;5[fZ5/M9)BLK)V#\^1d:GLI-)801HG@?VI@H#IE+^d;[^1gBQOZS&.g_Y
K)SF_9>1dJ6HKCAc&CB\SY^INN(fMD(5;.LV+BgPg)M-dY@0eP.5-\gc_5\N@J(f
5(2@TP2X]/:M6\<-Z&/#VFMI,/,3gO2BIRL.@+(J7DS1ZU7NC&K&fN23OLgFa:Jc
4OSCB?(@;#P9BdEd\XN]#b<g@:cMQ9V,IFPKNRN:-H]S3#>ZcNBGdQSO4^^WF#eK
PQ)Ra,M,6][cbT_AD4K>YX@C[WW6IVG5.Sac)(QB]TZD^9]f#EBU&#_BS=S,Q<6d
1N:TP+\D(<@FOL_S.GIF>63a>P5d+G<GE#BNJ>#D8X4bN:9<.:]N4NDP[RIcCKQ/
.(gPEHD#f6[Fd8:O[1eCJB;N/Nf594,D?.a9)A@5+Q<,XL@T40b7<Wd0eF95PLYb
WGD5TD>[cQ+\N-@;I.C<;+BD8I<T70b[bMVCK\-g.<Ndg\_40^NC[,YZd)Xe)=^a
M&c\aEDY6#.aYb>[EY.6MIMdRK1H3QEe(4gTB.</cF5EMdFUZRU(dcaRKS5W5eOU
<)C22WMO[WBM-G#M23e4>1+VI>1gg@HY0N6CHNbP=@M5G=BT_6d-HWTc?Z(DFc(;
ELbU,5>#HQ2-A&A<eF)6>[[G)8-Z;X,&F7Zb7I^.9^T);PTG&,6VAYf2@M#9g7?-
(7.K+54G.IdJSQ/8B;1J7T6F8eg1;#eM+G+VJ\;F[;U+;Z_K^Z:]>2ED(g62&QQ?
9Ja@/3R-,KRY>L[TO_\86X\99F0[\4\HT-(I(353H.a@bD-bZ:QCKR8\:=GgV3X>
U2FVI+Z\MLFCIJH8;0VD),=6QZU?-,RGC2RP8S-2S;LfF2>JUbeM4WK@G-6SRGM#
2<NXOEC6A\DKUA<7G:EeQdG[g+)@B?2SNLT;[^Qe\=78^CH82GUePa<aZ3ZIg]\N
;8<9A4,>])c?XALK9GFGb&@^P]c\-7N,RTA.>Z7<Z1_dTNMN=LC:cM]#9Y^&<6H/
GG3Q2IB&HG)9bAGD2-_d-eYVK:A,?UHY\E_L[2B6Z32SX5b?Nc<L>T3e=^bc+^fc
#.\d-U]WYH[N/6Vff-]Z\R(9a\-0L1ZK&\bPU^fXACQWY);(9?K&FFY67NEJ5>9@
DQL+b(Y[)\3f,@Yg^\&OV+S:;/VT6JDV5L:U[7cX_U#4S7+BYQXZ6Z/dR,;7FOT2
(\_KdLS;<U><[05A,:d/1\L195Z4++&S.]P#6:<+P^c/UU\d(6=);6;XQ,V,47V<
>>=B,bQ>AO5e_fe\(FK&7TeH>RO^LA&44IC^YGNQHX^UA:SE+\+b_TURM@MY03V<
#:HOM]a6=,Vab1EV2M,@aB<;[W/>G;P6D\+N8]G@7E\T8^6IYO)RY[]e#6&+<C2Q
>fb1,U;/P=B4:[53=c,MD]A,(?B-U]ZU_Tc-\[P<>5d/3aB&&X.)ETGZ2D@Y)Y:C
b&]bD+S<<6C.0=fdJ]FVGaQF/L3>b_Sc4f)/gYQOa4GfZ9B3(PO;+82[+Z0dSX2U
@EQ-c_\P@8c^M0QG&&=)d3Zge@??O8XV#NHHg[H8O^/44.NEcYN\@N69]/A/8L5:
@.;I1H7@X6V8UL1)FSaE#eT5N(;&X(;D(6[G#2:4WgOIf<[b6^3_+Q3(8;N3)-6P
f7\c95__K\PZC>,gB8\V1JM:adaee-B@0&/E7fFZa;BC)Z13H?D3,TIK&9YObR;/
.>gab<3,AYJD(CbEa]HgWZTK,3\eW2,]#\X>(7:.N;:JP(Nef9aD)OP1213P9TT:
)>gD\9d#3ZK9AZd-aBMZ8bbX\2@W&X>&_][=Z<bU5J6-,UaGL10OT@-]aQ]W6CN&
\=FTY)22MXEA0=</&WZ^T>QU1gLgY4:WJS;g_TR#LZ-5U/_K7[d(80/(A,]<S5:4
-5]1&F@Z10VYZN6XNd/M@C=CR/bR1VNCR6?LSRJ[YgWXG6\</(?=6^)YK?L3B=a,
YgTb>XU<[Q;>IC6+GEPJ[+@UbQI[3&:U;X^<(bN4+[7ZJ,aQKf^UF91<ccD2ea>5
V8:^-d(U-\H]gc\=CSfF8SbX(:X-dWdKYb>I].b,E=88G:&IX+f.?<:@d;T5^[5B
GW:28KX,fHe0HKIEDABK<E^#IF+AcKM_O?f_Z10Vg&3/-J0fNSIU;<]Z\QJ@Cg@G
\.AV4)3;cKCe:3-3/dAJ+JD#7FfXF9MWK]SLT+IQ0,:C8d)9M)G\H<7BRKT_,F4V
-&GVMW(+3+gFH5bTL8>T>&?N(aC<](.&0R47-<]g5>.KO&dTQ[W#BA+.XAQGc5/L
#_Pb@8@F<c39;.5,aQ5>8T2cT.JWS4\;)Y=^RaW(JB^<]:0_(H.<RK,)+KZA7@D:
)=E\(U:7,OG>U6?Ybc5;[G-?M;dK)a>@=6,K0&7PGf^ETXDQ]^;8B_0<dW(fM:[L
JFU\[?.RD9XP2R3NK2ZcL0F-R<R6Q.XJR/c;M9MOZWeHP,+[<^YGYG<fNLP>&0aK
5?55))Xc#:4DK@MB9MK-:;eM5XSZZCg<aX@VQ@^F_Y]=4F[B==9K@<]RY:BC72#\
&)ERQ+N#Ped:UK14[5+BT]97>-[[QNDeB/6\eSVbcaaU9A9D--XSA-.Fcg>)g>ac
_\#S5g)S:CMLZX5;J3eeI-P:RIQ&36-/2Q3F)H2g^>BZFfIEBb/@GC2_>Vd<X2@H
J3409:XP0YX)7WZ#<eZJf/?cM;N:SEI^dO/FbDS9K?PRI9f5AH+?APRAGc1&Sb/=
D#OSTG@;T=I,C0@VV&R<GR3gGD91LJ,FJ<76OH5ZD;QG)9bSf,Y;/edVe5G]X94U
T?5FW^]H]K>:d)L)4W^Z3<WDaSK5D_ECBO+QTG,X/O[g[(#(]-@A+_,JG@)^DBKT
bWd?g8E8X\<@Z4Y\;0R#D\A833PT&=?aRID<cT24+YP^@C=NX_5[]K9SFcQW[bdU
U_7.VKH#U0<<YD13Yd;<^.OE[FaaILgR-dZA:g[?cg:eNOB)bVC7T?4H3dOV;Q,;
G#Ab&eHRL+=?(bK;4PC/+?7HB(IUCY+,=6AgHNUX(.b;JWcNB#]W[ZBK]<f]HJ57
aQ\&LSEM<K>+BV[)KI^H;PC://PCF0#-IA#FPeBDODbQ-Kgf3E7Eb0LVHQcMI<:^
A[D>V2>d>[5QIR8:5-#fJ4N.+;Ec<?TL?<:C\5ad9:KaY:ZT5HCD>b&?N)RFHZT_
J&G@=.BN>)XFQWQaJW2eMZ06RC+[Yc9\d34EN2H;0N(MA=Y^96:@+^C5_8HEdcf\
(4(EBFePAPbX(3e>3>B&,@e(5/U_7bAY7BO/Z(12<gYQe^(d.FUMR14E>SQ0&.P[
(ALS=@CMD0<D(V=I@GLNPX\?DaQHA21NAKFF:;\GQfF.5_TT<cC+E\ZK=1:/6T,\
&AX+RaAJ:)DAeOH3TT&89,8cQ]#^M56;):&IB:Z1.LZIVXbGM+RbV.IbSV5MbGL;
3V/RVD\J?9<VOG:(R8.,M3DZ;)31T?])7(/0LTKI;Q@_:N>Z.6UF+MX.\(?U=V7L
GU\c(cdeS&7cM^HS<]cFDXG?&d#c/E39\)IIB3JQ/faT+J&^DeK/fR_e-#7OL2&(
H&E>;I20Xf/Z-86?9_8#5c5D6gKf5_C3aN:-HXfa?#8,bGIEGXgfcAXK3H99^bFQ
L(J?N[T^eU4<@GCVTD9,,d;YY3;#.\<W6E-c8>K;OP1980@HHC;=3EV0EZ\b,[Fb
415OXF]7-@DaL5a/ILgATS/bU@;b9,be.#4Z:>]dM&QJ6G:HH2C&J)9DPR&[CUbT
EDTD_]g-,Tg-D/f@Y>N\[,>&I#:HZg>FN+R01168@/d];<QB26L^Z(b.80eD&:S>
)?BNaHXRe>)S;INC_UIEXfWBYL2Y]d@-=QAU2]Z3\:(SFMfXL_gfH^?]ZS.5W6@?
,(.WV-W0V:&^I2<Ea1=4HKcZZ9c5Sa.R,.LTe-aBH3D?\c[L27C5?NYE(_Z-Td,8
OCT7+K[?DL^E9^\UE.K3)]7Yaf.gQ<):T>O\Y<X>>&1GZA_MNF@HJ0e58(0Afb\.
TFHDMg#<5R04.-41HW//877A(J0=<<(#Q<L=M3ZJ0)8cad>BSO4=DbP=\:S&84?@
Yg_g#c^T4>GL:NB&+eK^2.MU02=JN-HeIAGgU>GIX/NbO7gc;E)cW1\BEdJeT9WQ
V)14g^g;S#cO77I&6S5V9DEEL./.UPRPNR0CDb3AXX8<]1cBW;d0YL>=Y,1_QO:3
<K&H81B(N+=<E>TcbSg_[AK+7R;2B)U]>5)8DBGL8PdN>.2Kd\D5&H-SY/ZY[#QK
.8(N/+>QOQRO:I<[I97P(8?/-4N;BS.PCa+)Ed<RJ,7U;f+fEZ]Vf6HC9AQ>Z]>L
-+R=C@b/5C(HcIG9WF0?Q:d,4CP):>IYHLDWM]e,J;_,V\NeNN;6-90]>V9b2YSV
-K)eS(37=RHaGd?R/Kc_bf\Ff9)#bEWEW_&0]019E-I20R3]Ze9[E<P1-(CF#QHP
1U&(]eFeOHGW]Ra_g#^Zg2(Y>FaY<a)3N03]5<O8-BX^fSaL9aYT/I+NYFG[CN.O
FeTBY(PV;X(1gL)2gd#e0gS<Y+0QI(Q#RH0I>.(1,a0-R.5EXeW1U:;ZAM8_OFXT
?b,/6>Bc?dZf(MJ0f>(D_YRGG)6Wf<cX5aGKY1C)d7K,[JQUGUVe)bGW)7eRDCVG
-TKb7a7a89eG1E\B+>fFX=(g)87GgA,BY,VO+5bB+V79c5XeZMXRILESZ]4M0R8^
^:-+JY.12L86\&T^A/EI6QbN,UMU51861IF5X8=FBD8G8H(0aeQZbS/^URJ@OBA]
@e8GZZIHN5_)6MLg7-9OE1;&+WG9LV8F#@cRCAQWaF1(F#,D#>dgGQGN:RSfECFS
LM__-\^9[eTV+:X]NPdaC((8CN/N&5>Hg>7B7DOFS>AHATEY45PD?:P&N(>B_X>&
E_dP&S9gE,S_7OWdH5UJRKNZW?>EALc0;58c+]A,\.<[9MbN+/eQ@&Z9QHDNX+_T
QM[KZVGP;:111=Y:e>,_R&.<Q0O)d52O/(W8SbJ6([;]Nc9HO5dU)LVVSM3XS>5&
12;TC/PJIG55cN,c&/4TE[</L@JP6Jf,RJ)fB9B/A0aJb/dW)N+]WQ@706b-40XC
Y8f,DYL\).^0>;.?T[[:GD6@D^07fJd)ARK@P:4(0>&7cYega5^1L)RSIR-c@5Ve
3a#AMTE3/03f.750ceNNFd0\HW4WNQZ)[cV9RVM7TgI-C#@aBX5a;B5>=,Z@SFF;
6VN2KH)4Yb_f)ZTK&FW+.JCFSW3P&<a\KfO/2bIYJL#6<D<QY_?LXV2)=c[#XcC=
S+]f0O^\f3#,-&+XAEc89F:GWg7P;/>C7ddI\,;WK/-7@:M;4BdT6K-+/4-cN,,F
NL)Z]H&I(2E/YL7G5K-g[dM=6,IaO5-C611R2+Ma_,Y.8IY:]U78e[g)H_1(0_4L
e6F?>ecaL@/f_-aAe9;HN@9,G#G70fZLGW_Z^]R/@8(U)1;g>4?FH^Je9,NJBYFS
R6)USVKSG7A#M+aa0FAg/UOYT[-GHVFgd]_eWSP:[\1K3G9\^P.,a@c]G5B3<19_
/1ID)Z?-R0:VXQf/AcF:3V-BZYM/B1IXI-&5AA]g8YgBPbeTdJ1,P(L7fTC0L0U6
;K&5)Z;1/2R[He?.@5L,@=db=#&(NQB90IN[6c05B5;,].:6@PT+Hc8d8-Ub.ETJ
5bU;K;74agL]P-LSW5bQ\ZOWg.MF@)4AND[&aWdKLP0b&D>5)^D0bZOP=:S;fV_8
aLSLPX3#8:QO:/I0@H\R3._OCMLJ_YJHPVD/V8aQ1-_gNd.FOMdCC<BX>NF0a>8.
T&C)[/X\^cGCIbC7dG?S&1Nb++H5&N33+PG/RaY3IAdTV8L.]+UHF0:68I;QCQ[:
@1#RXD;5=ZLSISgKKJ=/_Y9B_8-IDDU,g(=CcV.-C>1Jf>fG1YcG6:]PM]d+efNJ
-1/UBZ-A-_WE/AG+T=G=F\bE89?TSHZ)=^OZC\;B/]W1G79fOE)LY;Pd/F(_b.C&
gN[WIDEe+87[0?Y9G)XK>I)0Xd#1@^4PY.UH(/Y:Z286)9N:M3UXP,MI(ecIb5YI
3QWLU#OgZBYC7^;,&BKB-3f]&[E78M#AVZ+2Hg\]SZ#(N8>753SD4VZEG:@AJ<H1
7&b:)Ze;;Z/9]@CP\eKOXAgCJKELF/BgSDZ)AV/9361(\2T;G8K_9/X(GLE(aa2[
EgLQ-e-/NNPGV=eX7961VMGN9]L2XN46.-f<W+N2#-:bb_R4GPdF^KOYf8TMcTCf
a?[=^-7;6Bb4PML\]Nd/gLa);c/2:DfNSYM24CbU8Rf5EB@AJQ,fb=MII1#3_PeB
6aZ,SBJ.gQ.5;+^O\#]:GYJ?4-VA3g)A&;Of8BJ>9CfIO=c4fJ-Gdc:4#9M.G^a_
^+(60?17V16U)HZ)_N81EN?KI.X;KF(MZfXI/R7]DNBZgF^@;b(?Z8I9F^3LN^QA
W^@:[XaAbCW)?WcDgIMFGU(>UC9(O>bT5c/^RDDb];E1N^.\YS+R^X1_WX5S0Tc,
MEAB_OZ]IB8#f7H<g1@ZMA,9QKDCLH,3X-.S3LZ+M.L-04VV_7/[.6f<VB6AB17U
aXbB5d3KW02>BYFH)D4[<,BE-ScF#YePHLOeJO]=g^-d=X\54GUZGFG2?S2Bf\)M
.JH]]2e8=E5F#M+7=&BZ>c.WH;X;MBR1DZI93+f.g&e=UW.SQJX4-H0C_938R_TN
6YI<(-8M.YK^gaPO#Y18BJP@L-.Y+GQ8#PDZ;]B16^;fg-=&TC_//4Kf+eLeP6=f
;\8I(4<?Q63>U[TZ0B#-L>_XABMQeP>G^/IT#6eE/\Z[BFg04DCY89<W>2+2PF)+
=G,d[<(@EA+YW9dS6c\8GQ/EOW^7Y.B2@gH_f[V(+INYe4#M<[151B4&JP>9)gN4
TIaf;Z@FDD1>Y6Y>MC?_,JI29WM=_D>)(^^WTBGN3KB>E\W<;>-c))-DP/-a3V\L
(.PRKdd0X)H>,A+A;:<I3G1f6YS=\:eGWacI^bS1OS;V9;aKaG/&&4a3Pf/f\K+1
U7K=22=^+G<D+gP\&;fBQ\#=QU+NBM/>&1cXe,W5B/PRdR+O(--<\<2?=Rg(K3bH
@O;QF[J,3XfL08:bJ-B7U=9LS>(cT9^dP:TNH5J88c9MaY29cP.BfccL,-\Ma[PR
0Y_=f2]ZSa07dY\_=>):NH9]8cV]J<YeYVBDHK.bHYd)+EZ?0T4HfI(BBUa/dC#=
.^KMHV9?[]9T6IP:2LL1;5X\cT10WW^4@#a?YS=(aebY\/0@\Ie)?d6dfPDCU2MH
&CIfGI?_J7CQ[7IHQ9W67aXc&D/^,_UK-)eC92CP,d2bNO8TDa;Gg>K_\MgROd_N
M2U@9\8ed]Y-+Eac[.a#.NL:TZ(>a\d<4K38Rf^b2=M0=KHHaIND4I<fCg=7@W/1
a;ZO_V2c3J5&\A\OaO<T)8IO36JG4e92e(_9_#b&=aX.HQ.;XVI/QS(9b._ASX8(
g0X53:+e=;g1C=:.:T?aY)FF5Z@S8+J;H/VD>V+fT&FcfQ_[N7WWXG,KOSID4W3N
0XQT.^VZG<1W2<I#U3_g;?S,7F_3V/NGUG1X3H>LgLN83J,^X8FKT0+8BI9f-TT0
1__A8((,5S]]=)VWVVKF+BTaHXYY2+A0EYQ<Q-9_S6#M?8RB2+;+@6AB;+4/PR&C
:T#U^0d1Rf[+FD6@9J;OFC5Y42\^TQKLHN?HaZA&SEdHdU+=>B)ZM=ScU0YB5XOB
19&71g8Aa7Pg.L-2XM-.=KBD;0;g0TCb49d)76[&8^_:=77U0.@Q_@OIL5AX><SP
ODX^bRb@RMJgHe2eRb,?ML8N(cER,]J+@8)Q:0VSH#7=eBL<Q54A4_4HAR/I?]MS
NW&-XQARZH:W073W1#2KPYgB0SKDVD;1FF__U^G3fU>25Z(LeLCbTM=B>,D^BdXa
gYQU6P2[+_6O^#6,F.;GJ2:7YI,E(BF<^OB<_P;044,>FKTDT#5X-SMNZ\(KGT>8
NR&f[d-51\TWP-><JF?4&<L9fe&45?8AD&WaT&:XVb#VebFF:?&WM(Bbb>G>^.TL
^F72H0f_FeBP^]Rd8SL@RJZUBSX)Y)343cF7aSGX56M9]GG4.+_8ab^TRCJL/=XF
\(1MLNC/8^dJ7^>+3QJ,J-\&1@dZ(^_LF.X?#>a0[WZC+CI[3T-(^^e?.1N^g?a-
_>-55c)-,\bO5GVPbK(L(Kf[E.]Tg)2N]OGH&DMSF[F6GA36UR0^@F@:FL5Vg6VF
9Q_\5^2;BO[EN>_/JW(/I9=]ORMUH[2;P32@Q;c3ce.1NXdfM&@ef[f^<#f<LPL+
8L:UaO>>#a#=dNNYd#3PL+@F1S2/IT&#1LBOYEdI1VF([\;U5g=UaO[EK[SI]#B-
?f@,7ERfI3]+)Ea^RfRIWMR2JMXWMZd8bg[AZ_9_JaYU2]Q+DU2b)H_]G^D.](d6
9KdOO-d]G_7A)^b@&G-42JVfM3cH:FZEI+:aA(=2<f3;TDC9F4/)F]>3ID#ZXV9D
KRMY/Fg(C.=:Ab&J4G&D<(7?U-R;2##U=-(G(BJA3V[/^#Z5f8DG5O8A.XBcY9<C
;TG/Q=bI_5,8A4&;_QHL.),ga<R.P>&DP]IPEUEG8gUKfF[BKRJB,JC)N.)I,L?;
eb0a3#]Ac_OTU<eLED6+YE0HN[IF?E6&J075;TF>PCC0JIC&WO/A.E2390(A?bM0
[@P(.>IKQ+I_Kg5+JT@YHVLRB9[M2F&@9;C),g:^bFW-eS;C=aC+8MAY7)I]6McS
#(68Ba^Y.LK/^gUgE&N3PW]BC7TXTV6b7+IKL3Te&J7.-=gY#=A4E7K#KZ.=PRGX
aNW)N82MaVI-)YCS^9f(2:7-_T6ERL_NE8W85D&>.=0[;@4J8a^AL.H5;,PBfH+3
8M-He\9[>f597X4>dP3?^0JJ@.S@@\.=GL,)#6/Z]9@PO/WaL7U^f=MY@4K#/D<(
:,H:)=(Ha00>6F+7G26_6POYC;\]DbKfI0E50WDdf&@O=NW9K6\QWYJ?7&-R]Z1J
FC=H2ZFAT#-(I.:PFW2,VS?U@9L/D:]a#L6:bbD88.]2a9#WaI3+G5eB,M[50=WV
>89]IU&INM)Z:1PF,DP?<U]]YK]I&@\V&,8VCW_Y-)K2BS;39>CS?LSNYBL(B7X_
0_T._e,JK9I3:<6ESJ\Id5CZ(Rc_Teb5W[63W+HF69\VdV6\gc1/(+)]G,T1b8d(
KM/C[<66>e>+T+a3X)<(61L,IQ9-PO/0&9U4\:@bN5TMH0WQX,(d33c#NBe6>dJ(
3_IY26McdMcG=>-37NT346E.(Q6UA=[#H[?/IZe1.[Y)d.(c/955b5R(B1D.8X^=
:f7DKeNEd@1][G)MCS?d3D76L?Mf63#YfO&:D4&]W\f3KJBZY].\IW1Rfd24B<gN
QEbS4]V@QeYR3H8(I9?[.dX;EE#1LceeDT^38ALZR()XD[dIV1?YIZ:K@eMF;^G:
T)-fT#e@2^NA\IL)&G-f_#)-)+:0[_R1,>]@^d0_EARLf;W5-O7TZY0XdFC?<N+2
U5)a#7;VGOB)/d64BSMK8PcC56:,1g#;N@F:M(Y=-G^4[J1&2CbV6.dR5cg.P7WC
>0;1??=P\E8M/(DcK:C.044PR:69Z#:&,(VUJCP4Yc)U\6bL_J>J\3QN(WZ_DVY_
UC,Cb)_A]<D#5)(&DA)O\<?#);(H)c-4(4Sc6[MUP3L]eafO1T2J5dIa>a5(#+fW
9;afd62;+/NK_+@3g;&DdaEE\;eG+SOdP5;@^LX2d94UR1)E1JRdT=[DNVB)4?W.
Z+.b/.cgP,aAXe5]9)d[]P7@gP46g1V>::P@^<2[dGMbKG@<74Z\_+0>/J1/^_5d
M^UK:96Z<9d>(M2\[Ec8LZJV2D61SMTC.@Eg11d(GB96BUZLHP?7^K>]#\^(Q4G_
O,^L.1,WZaa[L#eZP-Y@KK-Z_H1-X8cE>&/^6Jg,,,(X=\;]/[GP6B_T-DGCZ-d[
MIN\>;N#J]SRZ<.&7=7@?LKSA^2F.RJN:7UH#D)bbf^5DIX.I;WaAAf][/@JcZLE
G<\@>FB]D=./1KbDWX;=.1e+bY)^)e(C61N-AM0PgeV64/4^ff(g-[>O8TbY;E7^
0<,#\9?9g<XB[Ka57gNB+PO[LTd=7?/+9TV?=<7d0C+VKDRXXS.1LWZ\]PD2d&87
_DcI,YU1SG;3L(C3IF6B=C@D#QY>SS\)=E\bV->/bga6\W?da06eB30?)IA4C/L9
2CS/;^MUYIP.7-KD+F8Xc3?NY#@-Nd5)O?P=X^2N=X>Y:]JO3e,+5Ga\b>32E&[Z
F&bX-K9SI:Z\6c-gDH7dBZTY<LB6/_GAg)CT(W@]db1g;+U__,;ZXL>0&A09IeMG
Y<9R:_45eL\6(_Uf1fF-@A#;bSbS0N3P2O\^,74O,KJKJDX+D@6:+a&O9C\:Y+WG
;)CTPFcaZ_6LKX]e;YWD]dU1N8#>7L#XcFNU-ZVF=K,[HKHd\f]B06L>3[+#R>1B
Ib<dc(\J74&H-YdLbHa1MTeVf=T/GCdYOZfbTJ4K[A#-#df5;4Z&UK4eS3BO5]K?
M15E1/)3eL1-1./_LLG[:YDbJMa/V(e4],E_a^U^(aAW:Y9Sa]eS?P)G&6DOM6G?
3KSEgDJ=L,7,1QVYf/N=^J3cDQ^G(<bKUH+E^g\1cK18NSM@?6P]=3A2[=F^YE1T
[:bQ:O3-(36699T,Of-UcgDa8I9>P-#UUc2dPMaI,N<3M0SU[VPNS8B&3Zc/.8S+
M252SW8<aMR_4U#B80W.LXgK8(/U:g_?EFYJVa8K5RcggVb?LI+g)3f\WUV(&FJ1
A2/ZA8;7]]Uc+>C125NV?G\NH.:O\6IZ=\@KU+;&E\(SO?\6?^D)1IF;0L#2)+\4
.;N[(MX(H#(VI4&P(ZCZfag?W)L2@UU3bAV.4F5L/da?6Y+[[5GAcW;Z@_b\1E.I
#R7=3,IP98b(Ta(]49_P4V0A\GWD/#R\Zf>=[^gA#f&7[1_AAdUZ.BM^P[GEe2__
8G@.64[HfHIK^2.fII,R+^;NXZb:Z/<Q)J4Ha=U^@H3abNW1[W-N51;4X(NGY2JG
TOB#4EKKV2Ngd,5Fg(=HW&@Z)73A\cZ)A=(M3QHWTCR3;+#DIM25GDEFD#:YOYVF
@&/1EHM:=/9PF?L7eDd[--ENS7]Y_Re(>ZV0W-Z/Sg-4,H+]9-8bGY@=57P#CM@U
1MA30VVg-PaXPK^E4(SdS?VgCLDG#5V?E0;)^K2fZ9<C>\RB[#e4QQX=PadF)77[
0VU1e_X;4;FgDUTB3WL^><ZLD:O@.N/a<@PELb^M8J-N=@D^8MQCE)TX]^=B99-5
ERH7P0FQ;BbI[CZ<L#UHY>H#+@T8[c[>.=R9HYWSd]gbQ8Z5#De4f=LR7M+(]EZ5
]X(gG,7K-&F-E()TXS<^P8UAF-)4Ke+X[JTM&PMR:@DP],.fQ4BfBV1]O3ACaCZ2
6gAg=>9V<K4;S:(>N\0aM#ZX_TL:B3<G[U+#G8\6AaZB#75M:1F342E4eN0CaH+b
??XeWeZRcg]BPSfOF@U0B1[Q[:V&.IW474_9a3<Z2XaB([28#^2dO]f=JI/OL:P+
NZYY3V8;^@@^]IR=CV@)J3Jc7)^U;WNF6-9?NZGd7(B^g?EG9ARB8QQYG7_8,23E
aJ:;dOX\2>68D:)D([P-+.53+AD<EVOD]LKH6(T_4\dECId[ETWGV\=<9g7a@-(5
\6DJ75@XAZQX.>[MQ.>2(NDXL8)#KdH8-,U_^eS+4Qe=100+S,Rb&\/6)=AG7/US
</L=UA)L,b/1-&PCP5HX0F;7gT(O+fY+dCM@(Vb-0ceLP7f&1;a1G0X[W=NX234R
g(Q60XXag,7P\(:#LPXJ)_.\_]>NOVe0cBbTP;[/@SI^Rc[Cd9?C7R,g:_BR]^@/
5&U6-D?Vd5fS<;(3A_&4,fVEXRKZ+;(TH0YQ9<KCWgg2T3I7Q;1\O<I3MBf;ES/K
US6:M3cOed8RC10F>FD?PRB@P>dgd+JYCW<c8&g8Y,?<SU-^KE7L>;P+T;F(D==b
Z6@eV7F.W.1R\c2?F@KHJVLAJAS,d+_M+SYNE6Y/Ag85e>\1D3b/1J:CQT\I-,f,
13cHbdc)NJ8DSZF51(D0UHQSUABB^@g9E4-bL,3^W_ZQB:-TEfaeA#B:^Wg(X;@W
c:L.3WP^AIRU@X:&1bcJ[I&+9;>@N3\d4O<(dK2)^NC0-.H/GJ7F>N.D=-9@,,WA
@R3/=1c@#/I_SB-K(2YSc_6(Gd;04(Of&P7,09bKVB\LNH9QSMbgCcbgK=>)(=40
Ie]M.Q#+J+A?,YgT7Mef19cfgf@S=:1c^/IcA)N1@9@.GH/YTYJN2,eUZ\5Y#C96
&I?+CP:WFKS=6.5QUF[/BB?9b4aWGPX]FR.D)>]S54Wf3(dWY9UF#&?VT?4V3dH;
f&K7PcWUSNa/TH[)F-O^>N85I,]OeQe9:6L+7IJb3<b:#)BaH:g0D\FUf_K8d5_+
#H\B<K9TA+_5>S7Ng>^F@1>g84KQHX-Te;5AdSDPY,e,@S_;,TNH29W-X=.f0_>+
&2G2c/D,<R.Z3C(Q-_=1gM9d^IAb6[6.Z##PJ#aA_HFB:Y_@c;5Y&Eca4[9TEWaR
/D:1K>aS7LR;]QC^:T2;TD@H\ZA+[E=&RdCP2EIddP4?8KMfQa/)Vc01,L1Mf,42
XAFYO/OZ4eGf>1=-[/RWb&[>\Y=T9J561TXZH:N<\ZI#K]aaC.Qb63&b_M@:cCH)
-d?RAKFH0=3C_-N#:V[CWI)K#,I.L=(0DeP9HJ@/&,8BGd+Q.4E<PA&(^C[2I1I-
DCe?UBM.<6PKDWWLWZdfb&\UG;MT3W26R;EPgU=GgLOYa8[_5-&BE>.)]7;S+NdY
g,XG6BW+fH>E>R<]a_VAXE0caVbW]V3C#Q-[(H17V>5AdQ<^\8)H)9dH\QK;T>P2
:,37#]XMO=F]H2JGA\8cR;-9EG:>fF2aL?fX=YF(TSAI3M(>23#A8<0ICX8c7?MP
6/LYM&T?@/3CR1aE#[8[=bS?(c.d=W@#3K?YI_c8@eB\:2T6#A.)#:YWM39H;GQ?
XZM&?9.MY(D+?J/\e8TU&Fb@Q&=f1QPg@a&__e5Jff8aQY@3/L[;T\O@LD0=H#9_
FN642N7&1,8bM(eXFBTU/70W#\>X;29B3f0g6H]e\-Ocb8e:3eE.\G.-Z\Z]Z6SW
.2RC,@e+^(F]4S#N#G#0.Q15dC#-1?IWf4NRM0F5G)b8SY:^(OCC[P0,4&bN39;B
E/dM?9BYRFY:N#>V&:K8@KA=e?IT[[PIf8YW0P;<f2W0Z?:0IK3Ya(#FW=ZWPCeE
^-5RU/7#&3UbO<N^(3Jf_[72=c0K&Q,A&X^;TRe_@#94BU&RaSM>_XQRV/c0K-N.
J6d[MA2,L\M-S3^KT_G2#a?Lb=WWagZ/1_8Q[F^ZFMNg;gSCF:]bg?W>U4+OB&?C
6.N+?9]V+O48NS3^(]d;_3]H1MVc5fW#aYe9JRUGV-IQgZgE:4B.GM>Yf80C^7.#
9HRZcLZHY5AP;5@YZ7_TLRT2K=F:OSAf&0BbC3GDfZ4E;(?D_fY?09@9.6NDc)f3
JbeF?Oa.PGd5GML0#/F-D2NHRJ(X3S8fNB_3ZKJE^A3PX4]3(R[[77dM&^W?DXN3
QZ_G(TR8)]OO>SHP4&)W.Hg]NE2^O?;SdW>4,CGLHJ]2XXVeS.aL(]U9\J./)1U8
Q&^/LeJ2EQWegY>8H7(7fZ,TM1f^CM?F365DW3&(Y#&65>gAMGbIAaXVA,Y5&f2,
BEG?FbBLeSI4LOA.9@[.KBf;Z+,H6Y9;TEC-<[f#[N[)STKLQVd-4CT[L:f5_0L_
U,P<_TE(XcP:e_)\D/(Wb;JRN9,5V_EJ8DJ71O\JLVb^[_9cbX71+\\XR#a+K)9,
22JPG/.W^aN]8DRcd6]XbAZd]DgU#V0CCG=LVC2SXcJ:IGQ&Z]18DJaQ3?F[Lad[
UJ#UD06SW9A[S1(Ad8Wg,OU<TI7?M028b<KYb1.#&W-;:P7&-VM]?9@ZA:Ke43<J
N(&+\N_4LF-BSOSM.];;#fQN^D9[=R1)W</ScX(.=<.W7?W<XH+UCFU1M9SA=Me<
_Y#T[2=_IOP(@E:H^IU>RMc@53>Q\d4,b<C3C>4&1HY3;-<0YeE_/3(81T72gd/d
dZ<B7eMV@PUZ)89)B=L1@9=C9eKP=_f:O+T-:PU?8?1S8VZ7LYN=1\07Rb<P^XYc
SaF4[ea>6/N/+;HL&58LS9df.8@VM6])TcSfH7U;+7LR,TAR:SD5J)5M?#Z(9CK#
?JQX:6H)V8S5U4W-IFA2T;STCS.edZa/:0-YUU1HTAc3(#]K=,X6F+,(0-eW&/J4
\YJdS/E]<;d=\0NGF/@D:C<-be08=c@WS.7?7B)B=dS.Pc\4+]4cF-:?TM+MdO]g
)[\#AS;_(NQ^\IZQb/3X0A)R)Z0A:R-+^IQD-@NEJ)IS(_\#^\DIg(-G9H-1d8FX
]>\b,4QCZ+>G7C>5eDf_2YH5.aR]-X+@9X.ARadORFCg(a)F1K?TV&_T@>/?;,Z9
@7c3Ug^_cbEa]1313.RBS&X?;GC@1,ZN;NSe^BS:(:=ZOPSGH6Ig<71W<9/PVUgZ
BT&IeKBfM+6:7[>e6O=>[#6U[W9PMLN+^O>H94&7>R>6>J2,9I\,U0BA\I<^UN\[
HV<O^,1P+_0FQ[Se0&IG+F@TXOYM3.Wf2Ec1<#F;LbI?-:RH;MS/GRZ?&9[dHC;>
IMIDK)0:>VR)-(TC:9DZeD<=#59=T0.\8E-JY\Q@>(PX&^[G?1]9Zc,-[gV@)5SE
SE>/([3bI36ZZ)1M9Ka+X&<d=-VeK-@)).?MHcCAJ9Bc+N7N/]TIa.V\fXYXG&;<
<2K4fH;4Q/gO\Yf?44c^-T4\g:Y)9APT@)0-XC\WO,(V(\S0g9YOL#\,PG\143P>
Xc<V8ILVAfL<e4V<dP]Db6d^bF_FW.;d57EV6+Kc&=#SSUSc^>CUAP\RQT9(?]L@
PYag8_QIQ>a9HcHF/6906CE,BgG#fD-U5CYTEJfNHE^a?YFa>X23_OBN.G5e6c\R
KNC,?5F?/^ad7DTW9Xb.c>9MG?Sg.,YMRbAKE[N/0G]RV_&)16)7/=[Z:=eJ52[A
0/LD^4>(NFYbFWD6gNUZc=5JeOS6R-K_c7b1ba01B@F[7fAec9^bIEa\b^XNJS1;
UYW/@eMSMWYMZ?8UMOEXac3ZB@(&(9(,/?0][\1-9:^P:[MMLaF<&:8Fb)>)J6[J
GVHT3D&V4(D/&<3b_1Z3M@PDc.QfD=JTHabVIEP#O;ZFL^E?OBMGc:TLE>(+VfN+
^BEaca=eM5W(\P0]TM4\PRN3gYQZ8)7[M,RN/eC-0b0(L3A>^FS(ged<XZ@BU.Q7
[[ET1F>5><HPZe]1^^T[0_-d-YY_6CN@;+SDU^K/7A+cL.aWV,cA[1LF#A2R_c0N
=Jc2\>H+9Vf)J-5DKT_/UZVZ5_J<Ye)GO4PecD>JU6KU;:.;)^3^23bcHU@WDdWU
>O.\,aV5#0.YL,RHO(?LN4H^V5bW-fBd_D\QH^JEVI7aFa?<=]/VB>e+T9@4X[>?
Qg2IR?g2SXa&A+52V]?(A=LJ-J[T\Q^@/R=RRPW_>JZ-/.R67SWVF\RZ>\7=:3ZH
2^N\CU4Z5#48MM#(cU3FMfH./aH[82&M,D,;SfIgAAf,[PRPHE@;F9B<YRdB#=WU
c.GITH,80>S>dK_)0^=W1+-H:U_;A?(HMcD]:B+A[:7EH75)eN5F_BgDbNQ#5:3K
B&3A.1A]fGbH_S<CXb]cb+A_QO-bY/?I<5U:9I>)#M3E&J-?U04f>Gg5GW#UKeE8
ADB;;R9KHD_5GK?HO,4\]V+6cLQX(&2TC6eBCAHD:GN;#]2&VTed3@^Ae&&gMT.;
d9@^FP0gX,f9dR4=1D9,K1OTHCVL5CRDS38//2RRM0#SO77H4^b[e86@:(7(;BB2
b6]XHc@e5=2Ic<<(D)-HMPbA7DHNI52/\ag#cW]RRYO86U2Y>XZNMgYG7@bJZ]UU
-@.S<#>\6+(d\&&3X>5\=X+Z0?b7/]YXdV]NE:Y,BNeI+_G,7f?&U&:)3:X365(_
d+e]?IM[SP74Z8,\VPVVOB)[9ET\VGT2;/aY7G>1AK_L_4^R7S-6e0=0(DU_#&P&
)J/_-IfO50b=K]GE=/dEd6->]I<g/\9fFX\QL7HM6K4F?^cUJ^#Z]7#]=.=VfTT=
2cb4HQM3Ge>?BK3)LKfa);.4J7>G#=EYA[Q=U\#-_@U9.]3.AX3JX948GT0Eg<3f
2V<CJa+@\ZY:6IWJb3JQecZ=MKb,&cRNPGWFZ(P;<=-9bF(cZGE_?A;Be);8FZH;
+WP-\PcB<:O.H([C/O;()D0K_=a\\<]GIT&?#TgU#LCF;+2;@)K[>2X^?[E7NTJf
LK#VB,?.-8g:KBBCa\CU-H)?XB)XE0<d;O7\eL263bE;2(=V(&12A,?&(L&W_:B9
-6/MbbcO25>L_0G3;6-SAT<KKdf)M_1]BFD)Z+Y?e808+M;VMS^V>eG:E51eLRR8
TC3]a3^S8Y]/R8(UQ&/3^Q?gE3;dVV=)105Z3-V21=Ja?K&bF&bU41\/=6Pg331R
^.0d(L;)NKbGBgBQ.)L,,-BC&6TOXVV)S==ggCT.8IXeV?6IdX2&-6AZ@GJ-:5aD
9c_F69_7>)4C1@AgL\[H[LJD6QJ67G)@eCJP3B7MLJ5-C[2_XKd4,Eb?<H^=fL4]
Y52LdAAHK2KBO>7BU7OAVR3XK[>]4aCScU9WecXbHN,fRNQLL](Df@PD;FW+f6YQ
WTN.#>Q3g96<O0^D7LC9(@XZ/aS?BaU-3TQM#HbINM(4PQYP>C3gE7Id3c0-MLTX
fV2;+HgU:C+&T1#1YA2SZ(H+\\RH-A]:F.@HUE-::=b4X(L&4G9fD_CJ3<,CC3X:
ZE[H?7<F&6E-cgWVL^1JD3e+V<R_)_N]WN])>4Y#T)aQC([)J-^D934aWW@CW.b:
R>fa#,>R,N?VEA+RV4.4&PJ4PM:;]=R/N@]UcD[O5NO7#;WBKC&#@=CF8+a;SMa^
6N24d7g#>f7&2-cdUDH+a<]PDCC4aa.C7DBc\^CO((d?S,,B/+I,;c-^EH3UYa7M
Ke/S73[[I-Wc<Q]S@=fBI,,-RXTDB25Q:+7b<XLL>Jc5\UOA53WVac1@6Xec4QYO
:OD1-\#G)OGGYXZacZP4-,BD/[Y<D>.;X#JOF>6;7M<)ZE6_fKK3fEX[-=c:RYEY
E7J(G.ZO&C2PRgPFdB5M88C_6/?-fT6^FQQ?Uf420EM+C=41]DgXJa^Y7TZdf0@\
M-gKAFOfgDS&Y???X.UA3-O;\A2\.aSEf9cR8JF.V#;@&,I.;7UX6]Y6aVPE:gQK
1X-R608TOCS4YK<7>VO3\0=-);=QV:-CfT&/<&2A5J]gdc,JC+)W#6F#=a:efg61
:73_\I5DDZ7ORPIcM[JK(Z,<Y-+^ON>0b3)WM)3.Qa6;9^FR5O(dS>^d\2NB4H=5
<=\,+S,JH(b45_\8]<4SWNY22cUVH^G<^DWI_?YA0?-UHd44-88X]BWBD<<,G=7?
a6)SQf[R1C/-G(O)1-V[GI0[>LK&?K9LU,A1(\5A5,HZG()ZcBR1AL>O&<fVSDE2
CQ0A#H=@\)@+,5U4?e@:^Jg\E\F25fF2SM)_T(MSWPXSRF>WgC)HGY3g].c@g&+f
_AV7XKUJVI-UUd0@cde]YCU#;c>9fd:=@g9EZRM_.QXS]a8Sg=2AQN09UfP-JaZ5
(/QIAB,IR]\-S+@<f=S:g]FQC5EK;NW]U54FX7#eg\+:K.b[#+PGcWCO#J\SV8f?
YX@=Dg&W>0.8P?L?,/92X)-R,C:&fVbA23IZRM.(P?(KDZZ^J&ZV;M+2FSG;Q?+;
L4>HFeAZM=gRCC\+5:-HgDc9.S^1]=5f=c-S^\T^LK>b@.MGW/U8[CcPXfZNgW^C
fECNQXMZ9,EG4L+Y?KUMF_d5;<>_1[d\+SZOHH59#:MZC<WQ>K+Z6-9J[KJ@<K16
5K9OYW8:<K1FK@:8599AP>,g9Se.K26M9H5-;78^b];=.c=CU>^\P59MNZZZ/DcV
98J=d[E&[)aBKP\IQO3:NJ;4bDP[-\4XEF+1_[Q.K2c2A;b_^QS2SK#JV.1O-R67
[\E+LZLf#bCXR^EC8847_M,367>CgLB7CVHR4;+S,\(X,?ML3(eGEd;O;@[R7=GX
7d]>bJJ?\M>fV:/VG()^9P/7cMT4MJ2\._V=C1L,__K9X8S5FaLHbD?^9M=,d>ND
J@SW#^DE6P]W3?E6I,PU-67<4B/U>e9^RLK)BfWO-FOZR_/W\aI9VSDg&4986&Lf
M4+P[Q0RfX;=J8gM;[,RaC4J_-(WS.1P_E^IJ\G<B2b87#6IIA[A.SWe/<VUO2;+
7P@9OOK3Kce;?/=V4_].VNO)[X+:&;RY+e]QPC1NH7b]J8UH]J_CV)Q_BR;\W7#g
a+I<J3FM=S7(<VT@B_I[gfWbd5b>WL/Q^UAP\;F/JX:.ID5B,QO2(&;FHL@7-I2a
G52g7d@2SJg@f\(L6^RJDHgMI+2eK7X?J/BaI,.gWZ]R@Xg_WW0CBSN.11CQ.fS^
47L<11ZNAgI4UeK[6UYX,H-Z9:Ee14fd\@C6+NL?H\G5):]>VPJaGZJDY^GTHK5(
fHYWV8bSQfg@/E:b,T>HaXX&YSDd3(930O,AELL,d5/K&E,E]MMR4/,B2#VWg\d\
@79d-L&746X:[QQ^UDYA1G_]FH/SG38;Fg0Z:MNb7X_<)G/RS_2ZN;/>#3)2KDeG
HT\J;Jc,T6degKMYGACe,B:Fgb,Wd3b_5<I])GCZDK/TET64U/.X8.0_7)9:CC=A
0?9<\,4E)I+ZZIYI1+a^aKZOR[J2JPS.E19CSG:VG]&.0BdaLdd1RIF)e1>F5#1_
^&9PA]>@(0LX\M:BAL3<<[/\K05ZDQaB-H-_dKRN^(C4D,819Z.K#P]-F-<Y],T1
WUCKPT<0MZ+[>51W4_AT40+,X&^DGC\Z??T8Q<0[5NS/W\]KdE+2W;&UQ67J@(b]
.5I>FfNH)OOAH[-PQ0e1^\__^W<9f:8&EB+[XW/PP.IJ#4#B>R1B+aH2TV_,XH1R
d\2YD[/MR(5EAUZH2-6aNSDD@Y/a[H305CV_]9e0V5MV91A@J\_3DKJgZQM7+A(d
A=c,P?P\.CBdAJB(&SKU30W7L8+NQ98gB580+5CKdV0;N_CaY?]LMgZ-16EWH6\&
QY(B1PN>OR+V4ea:dY5L1?;[c8U2UUE[[M]4dD>I,-1O@1\?QTIS.]C72/MF(ZR(
,gH_1SFV0YO8?_ASD,g#HEUEGNE-&[aTIfS[#cA:.)9IOb,L3MP[\\=#DEPXeP/Q
&0UIP9I[WQ)d<gaITJ[7L8GN3eMbZ4\IYUYCKYZ0KI=#[d,eH8V\;&95Vff,8&4=
E>@Z?FLI4_Z@.)PMG,=ef4Y@2VZgK7#9R&F-98NFPT]M4MJ:^:EA2CdGL9A+DGB/
704K0]=f@O<;+6M[Q<fgB?CI>VgY\V(DQ)_PBMg1\5[&NPRFUIV[gPfXJ\ZOGD-)
PVNQBY^ZHIJ5b_IQIFV=:[\D1ZOC^V,gLIc9g:A,Wg(a<-_I<_[#cISNO&_O(1TA
BG?fe3G08\W)3+2Vg\Y?NOKVBL>=N7ASSbH08E]G,R_ORNWUc4T3^.J#^GG?-GaZ
R0Jbb?Bc^R2A;VXc[e87R/1[./UD@DGPcEH\f[(7^QZ/N-bYBb3MZ2JVJUTQQM5A
#8+UR.L@,GCbA8aCa9[MSCa(>+7Y13d0LK.dUMQO[47+,VR:bBV#S?4S>\\G16&X
ZS9MabRPT_,;UDN^1f8G2>L/:,N^>&FZUA7GP/LPLDGKLB[6/.8SSg2e#_g]N<:_
X&+379W([/H,J.EdVZYfTQEW5+27WcZ1&4TE?#)3aK1(#H@DT-5YLK&\#a73?#f8
C<O:-#HL1DFBP<f&S:b]LH8E=CME[&+GX46MN@f7G+E\P-9AP0MB^EG>8?6^2GBU
LJVGA8dH<D1F]=+7]-4>@Na9K?HZgd:;5eET#_6J75A9e0IHMR<9UU)ZV.f=FM+U
K,eEM(?959eN^[6?CPE=W/<+ULCTYF-bJCJG,\MQXS.+_5I-=7+92@)59ON=K+N_
?.;U.RJ,70c8(C[WO>_)=J_02@N1P0\\2^Ra..CYR0g;4YV9J9fOD<ZWF8Ec,#,9
7He18/KVV\NgBfD8J@fg)b0]ES_E4IKGA#FZN4W.d0XEVPZOcWZ_GSV3/+9:SXFB
KU7c<Re@8<9N9OYYggV0+1aEQ[L-E^/U&b57^-(JJ\.&(ePIY1DYBSa(BO7=1F\W
8+b>14AJ(^-fEVFK9Z;QO[dEJW-BM9G0O>>\U@[MAa#L6:TM?,K\@>A)^)aMb#&4
7E5KZ32]ad[)Nb14O8ZR)bY)I.I\290=]MaQK7W[0<+W_-UW-Gc)00S=^E?GC&>J
Nd?@ZH,<LN-N<N5:bId#9Xe3Z-O>c:=ANf7RM04X:@FD?EY35(NbK6Z97]=2^8Q<
1b3P&;.15Uc>=ZTF6TEZPE.R@GYEMB7G)b(S[c/>?YZ\_Bg^PU.(1X@3b#gc?P@D
XHJL]29-QBgW5RN-];D<>SI6VdJG;d.J#R=gZD_L02]1?5^e.XVBM4.+>dG>7P.8
=fbW9Q:)G)B2.DD&1B?A4Y=gI4]b+JV&?KOOEdF93_NN6LYecY?.&SF@4=GB>P\b
5BdSbL#6(2TGIM;AX0fM_)&L88FGNB^GLL:]HBBQfJ?,B>7ER9fgY@@B-A>\+3V+
G7>.9DM;K86>0D<]EOX34=^bI8OTQ69cFI@Hf=Pd2>YNDLD5DbE39(/b@KUE^cNP
QH)+N>MWG(6Oa]75Rbb7^2a):U;e/2A(S[IA0a<H&65BW.A7M[=?dfe^K0@[7M=S
/:IYFfQgY.#JHWS_W5S;>=F5[,Gcc=EcRWI[&C)8g&::)13?W73(I?EO;;9&fGYf
6SKYM5YOU=f9YF#RMUP?g4F@03WO@QDW<:29:4fEY5P,bZT7KWGfCG0K1M#7\ZAF
/Ta>LN2\=Hd(@6L/R#@-/@PJ/;Df4Z-F,Oae.JFT75GRN#7?)3RM(CUDIL=9d]Z.
WW&A9eJMQb0EC<#)RVA15-5NY]HFd9=L44CNB)Re&6>4WN1XCDUZ1b_3]d6d;X;+
TMO-^TDg8@P&1f6;2RK)HS69:>\;PIf1b<:Y_?9=VfTXV0KMV&KG]]-1RLM8b+)[
W.^L8c3\YU2U]62J0N5JSRFUXOBWT5=E_?@?_C5]S7e8g<NOW5RTK)/;;34&3PJ9
TIO0LX,S.RN8+G2#MdD1LV].W=,(7dHaYBV8NfEN<#1Zc?SLS2ZFI/6C6IXBS7d#
.6B\I&bcK_Z+V^>4<3c/6W#3OA;TB2X<MZ5dEc)W1&_[c_(cUQK[H+-OSE/@ZR:e
<J6Y.^P5#X@2(K;W9B0)-Z<]C)_K.>^Q/[1OHF\J[NQ-eX+#c?(-50SI:V)W_<BQ
\?;-6;3@9ZU4?4[.\=9b3:_^c>9#>aD7;\^YRF1V.T<MDFGa36>6HQW=#^.1_2FR
ABQPcKb1S_GWYBR<7#f.]+,4/D0#0K)G3;_7^)0Z_+QL0UBXID2OECKOUId\19)P
V,XK^<f;R0KGTFT&-?S(&KQLNN@&TJcgM<6\bTB8<CGMJ)ac[^TYM+G\L4AAK?\I
6/VS)FYXK2J9C\bb6aFETU68193,,cN0/BV2&&3]3(^bE0:P#Y.0c>XT6:Q?cI7E
&8a42fR:c0(eE.#0ZM[WNcQX(\AdC,[T5]QDGDbZdL>d.I4R7XbS_CM443#;e[EM
G0M9=L+1a.X.^GV+Kf39P3<13&cbfS1acG2CSDX)79C+NUL5Q2Se^faHRd;XG):U
/?-Q08;AFZE@gDF8&JA1OMZ,M\[S31-P>;6NeH#N3;L,UI9U)P>NYSc9PGH&RaJP
G@5Z,b7&>&OcKW.f45G/4370G4W\T+3?JOLOLRMe<7(E8Ua?4-]:#P6NO(;K/[cN
3]Xa5;?E2XIX:7-YZG/X5G\-1f?/@0\EUbFJ@+=7Y@)0>C&eULIT3#@RY^Cf33]P
D1._R#FNX6]eJOUH)B5=A3R/4WHOU)<+_UGHf^.L;_Q^VVY@NU\2FXR[+=Y>\HdI
<D-K&=)6Lcb4bPPWG2=Y>NNV=U-Vc&+;Ba;50]U@[MdgW@CK]P.RPgX)0;Q]\KLW
DEX[ZG<MLg6UEDH_T985V<adQ4S,(7>[XAM@Q.^9\a@;[7EW>.U+c0GH+#K^&J<c
(8JGE=eL,fL1N3fEaD4@VJ@b_><[?C6W;UNW]<;J]@1NVF,]eR\(c7&0f@)L3?4&
#(AT_S^QEJ+G3a;Nd9]EU,6c:6=Z>.^/\4/E,HDZSWeIf,+JT2_>87f(G);;=K.e
93,L9T<I;[509F#\E[d0V?dY[AHP5RF218X])I\TV_UN@TSBKaXTH)g[B^V.8G56
+8-2\GI_Y\=[Q<E3S1b1cA;?62bJ(X<UeHB6;R@Cd<<#]/V,BF^^9D1AD)F=2bfU
P-/\2GN\W\ETZMX1Wf?bX?_;0#,KV08Y8JdO?5Z&-I^I,@3K?SQec/@E3NaPR:KP
2J).9ac+K[AB<6X,Xc3SM_<1-]<):HH,<JA[[e0Y.(RDa9+P573R\a+VW1bMXFP/
S/NPI,1;C,fZ(7]M<_[DE&H<+C)SH+NZ):4.MYe8aS8D@UdJ8:I0CEUK0PU_J#D[
cHg0gO4+Gb1B5O?c)Z_ZeDVXc@Lg>S-OY;CRH1M+S34Z,I:I-M],^:OTG,K9/[?&
P_R7//&7+>,6Z1Z0SWF:CSL/a#[cd&/>5Jg]@M]35fKUQ\Cb#D:OaY&)HYS=4d6L
DSG[#8&W44ITT6>0GZda9NMBV;@;/5;.YbUI/BR@/<L-W]F^R7]77GK5_2d2D:#7
^(BO92XId^14d1>--K;B^<FQdb):_YW?cM+d<>QYdI8]2c:WJL@[a@F0F&_5UC23
U=QX<?DBLeH]d>N1>F63D00Y2XQ@R3X(5/58=^<7\><3(X1KebA<,&f&\XDFI9AI
3SE^70gL?2OU8SM1@Wg;5W(\RHJ.MZSL53Lee=4QLV(g5QL5M+(fXGcXW#7O66&f
e2<VS,H\2[?X])YTJ:X\-Id3IOBR[T(c[eC3_M?GG]SXWgM_]_-Na0NT,/4H.KXg
>>AeQ,8;:B+XaW6A+U^2M8+,R3Z>;(_0>&SERd,T16U/?K6U38b>b]4#_?PGF<J8
_HE\//-Rec#DeRfaDffZT/M5>02Z9dE&+.375)E=/6=](LdPc[L6>TTc,X^[SAIe
4P4WQ7FGWR&[\3FFDO5BS[U=b8S1(W8OWQe#JV;=PPK_2?JQ6;SE21RCX^A=Z65\
(29+FTfSHc;HN>E#NIDUMNg^UgWT=N7EF(?PEU-X:A6<?G:1U?eZI2B\&:6,+Ofb
]6YRffa\?(<>_c/PE[)cB25)PUL1\>-(eAHH9HC_LW]^/<I&&gSD<aF37DP&?ZJM
YIX0/\5C9TB4[W?<[G;#=]-<Sda4#OZaL0._H,e@=_3@]ZP0Pef4U??FNGNNYN/d
a;,&,^-5(_2XJAI&,5KAfZ]F-D-/1cESa@f]^F)8^;9&XWgQfSSQW3e>V-+.-_AK
JD.N/OSZF,B&<W4T8TB&aB=5X8Sdf\^35\PWcEQPP.T;)<IR[T7XWDb\7?Od><[8
EULHKJEP5gB/EE;?VM1PQ0HCg#6[4I=O>d@99Ge-1@VHXG6..F<@PGe=HAT7U<56
SPEdQc^/W6<GXXG]F()<c\H0I+Z;//6+\^63,J_,D]=TO9DJ1Oa.\=/93B2^WE=e
D:;;K96A0R_Rd@.]G2.fK<(,/B&O.B,[Y7@VLbD5.YZGF)]Ha+DdQGSfXZ8Fc:54
aJ9:<McXLU<X/W4XM]0(7a3[#;:.2]EAX,BQ6TLBEDL;J[?#[IgO3W27H.(?\G(=
NXTKeeJJ8;V_HT+&6BC[0-YcG&/.b0NLYNZ1[371L3NTCD+SNe_9RbM,KZ_I&WWY
[H6a3QFXZBXg,],La5Za7/Bd6;e6&2TPE=]4@1a_XaEb4E#dSK)aPPf#dY\F]]RK
?0.KO]YQYC\X(XO)N0N79W=NJP-A@45^]_9Z,afc1&T11b9L7HVRR&Z+FU+T=1Y.
@f&GH7V6N0ECJ(>8.=#-#>Gc3T(Q-)e/c#R2RYTVKcOCP;K&O8&bZ7/[1Oa-^c[E
ELERc=V504D>D@9>T9Ke3UD:A[(cR#ZE>d@696NYeBTc9<0D\A[G&^c]^=+R7.L&
3,DZK#^FUQb:ARZC6ZZ1c\;CUF8:@[a^OP9g\=-<TE47>#8VQ)C6_X0FgTH@]U;E
#B25@K@0fHa12gQN\GS)//X)a-27?<e.UP8X(3KMdc^@g=gR((.\)Gf;W/g-G;)0
0/[OO)2EMINefFK8gJaF.,GeKa0+2M4L891Q6))WefBPL?N(6B\]&;/eIcR9D<gA
57&)(NX2Z,B(,<GP.^JOc(Te45N2D-YJW/OZ\G5XR)f@;&fHGM>42WX6@@+70eZg
3dF3dd)C(Uc[I+a6P^H[c8=VDQ8^U_1(/R>2[)&2;f?e8W;4ZP:UFL\FY+fBbCd?
&6<&9Q@2F_FL.XR:)/Je=Rb:H,:L^gSL2deB[[2J:>C#QK;a9R=c645V1EEX/?5&
\Q#CBCH4>a:QR4KO:C<+EC9-Ybc8A3FZd^_5^-Y;N;&ISQ2X6]43:a-]eYS5dNU(
cDYPI;f@>aX?@P##OQ<?BI&-4;=A^-.W#NecE9I7-.)I_#I?bJIg8GU_Ee7+MS8W
^gH)-7PBB=(b>f1(-&/,L-&ZM-)<2N6W_(6,W?H&KXJ:KO5X#O4ZHAY4_T9g=?VQ
SXa(DZ9KAcce_O._MQE)]F4Z^5UU6g.3-Z+be7+C5V<AfWBgc/8QRfE_a/7IMK>c
dX7^SE1J.3D4U]b#d)R>EAA?HE8=KX7G?W?^eLb2CU<RYd[g=/M2\.P_JP[48:X>
J4)ab8f<PM-@X&</SL1;Q:Y)XLT\P96+/+aS\.L/KK<>/R@d<beYb<XS4+DJ8J=A
?BfDMA<3IO4Md/I+bB#,LNA6a#Ca;0F2[?S/VB53DT9eCJA0B2@+:)IC?;7O]3;S
Z[VKS39CS)@K<0(I)PG9CB?MZMZ;L-bNC]OX,>[?5##EA+AVA7)M=b:I:;1c_W@/
?3BP5g0Z_1OEYA4TO72<d_.X=W+Rg9VdRgTd\B:B9HR=+fLP@?&+=a&fNAF/b[(7
gM=,IV=GI[R:daDUUbeHFcV=d-)QEX7@b8AGH>?4]@_A:,6g+,FVL@+V,4Fe<<7Z
ZfPY87=71fb83-V=1.M,E1;>C\(SBPP4CaH>5M9W>J<S2=\DIRe)5N)5QBW\6gL2
DLb/^Q);#M^GE5<T^_#0S+&VL[\WJY\@]62T+&f?-(@UZTbXG._,aN64D^]FaV+U
-aWGSc^:8L(R&F[dG)B2W^Z<VYSAN#WP)cgPUPgH<BKF17fM&J@eLVQ5gANbY9RL
VA7O^4cWdKD7S_=Tg&SYb2GW)5?5&B,^)&]MCW)b5Og8/C7E#P.@fEf&>@GCe6V6
GYadX+V_-/T8ACJb=)]U_Y?3:g+B+bO]BXB3f-<)O9J=_&b..)&\CQdCFOI8TeZW
-P#R1U>C5#FI8A.JTI<c4]5;e[0H2aeS^PYT^TZ(=,8f/R/6F[[aI8c0?:_/];8Z
G0f_PGeH)e_9E25X4LXaL_L_DYaAS;_L7a#0JgJC,6A<C0MBe[cTS>[\O--B_2WQ
_X]Q(V0T>_;S,^P@3CT9-3/VC)WG=VGR+#=G(b,2.PP+cB].^HB4MC]+US#HdBg]
CeN2[/bN8A+@V[Q-T+ATFSB1WMT3(F,cTb7OB9a2XYc^J+MBS+L0\R8\aW74Y/Ka
[?PX1=O0SQ5Ra^-C5.JG7],8\?J3O#;cW9G<JF4VS>)GS.<+,0N#MACOf0\R-^_+
>-[D?WEM<LSK/NWccLI[g4A2\F]M#e,Y<?T7?BAF:7+b=+b,06MB/.7NcgBaL[(5
NI#.0J^MMDIA72d/&ZJ,M:WeDGTU/>6dTWe7BbUTP@,G09agg>[+.VN&V^fOBb5Y
9bMc+KEI<&4a=KA,5B&-3DDU^Q5[ZT6A)[/+c3MWI,1>ggTfLFW@@XYUBT+M&b6S
0,dO(Mb2Jf,US^JY\I&_+EV=J^DRX;[?E#+>]N\U?QCG+<G[RfOUbgJ@4Zc9gHDW
b+UdgdMGYRVBb5(1MX+Fge:>AB/PL72dK2^PL\;AaS,L2[&5Fd1B#>d&)Z_4]2V.
7&H#FD/[5gZD?KfFeI)<CPQW-PAS^1<==+bWGPQ#@>,_bFd9Yf)-/;?g+D7MfIA0
^?3e(1c;?\&)X?#?[-UD/]JLU:S&>F:1&57B5=-e0-Ld@+@L+PdgZ=cF5,ACYbPC
<^Fd)3<2Ac-KTAe+=&BaEZVKPU+7\V1IA=M6#[.9e4D;U@ZbQLC6P0FE]XZGBH]g
S_Q;Q9A\[M-^D[2>]X<:)?Z7>R]/0[c&X7JDaY-.cT)JNCM<2YBZ84V\f30)JM/2
dNA8\D.VP;:WOP@AC]WWYI+_[CGP1K(bO1Ge?fd:\PB[)UFYZJOHe[(@6:X^S\bN
M[@?S2RP;V:U<RZ+J#LCFe+J1A8/V&1Z3-255:NXAY0:c[ONb44K[&2V5AHaZ:ZS
K14\-.WU_E7TRQ<V40&\N(CM?4F\3gBNSOCAdTDa<0.a_/R-R=E)VO;>Vb;[V>>?
E6Z\I]+_-MXGA@fF].IdR@SfNa9>AFD#<bIC+WUGRFa<T.DRU;R7d<,HLdNK4dBA
,7YEHS.3QHc[T1g60O.XXc5]^OFU??1Z+(A0eP&&a-T50>0@Y:OG(IfFc42e+UY+
C^1@\?KJ6HYAC>A3.T94O-28g<.6b#NTFDHD:98c(UGWZ<_(N56HbeQaKB0D7A:/
P8+5STgd23-KF]>X1Q8FL)G/;RLN@HHV.d>E)#V)=4BgUJ5PA8QF?bE7P(b\35?f
#3c]KV+bFaeE2JID1(\2]dBTP&YN,:TBaEPPT+HbOZ,/SK#:YM#+UG/EN2DYB/=<
cE9)2;0]M3(HE>_Q.=J+dJ<Xac0O)[C5ffWP)fKaeCN14dCIO)4bQI6Z+I<AX(-<
]^/8MQ#@M#^YJSMc[BG+_/f-bM\24XKPBda3OV[cPN=]QS;@YW#W]AD>&#K1A\@4
L-+YI&07IL1b@1AZL]9RPF8?G3,QEVHY4bU<?K0OXJGScA\83R5Y5JZQ\:@eDa[=
60U+JH:bc85MHaWPD35_C<NA3=6H[67[ZC[L5B?Wb^e/VbM6N/[>K/T_AZS8OBZ)
AZ06-;74@5V&?b\7WgN;CY#AO#\UV;@Og=_.5ODB>)cg@P:U4Y,Q_MN1^E>;b<0\
9VL=;YUB0-.KedeVI._\&9_#9&J,F&e:5&JFF7N/8_Z>;DI[c#R&O\VCV=?G_6T(
>5YC3/S--8E)SPMd<^_CF&,b5V_-)8>5We4^^&(?JL,D#/B@UagMD[T[AQIZSI(Z
OS-L559D,>C.NJ#P8UeK7//bBR+>D14N>fD3fU]7dN=0-SGK_gE#eV]\,+=RL34[
N/Q66^?M@9K23-5318aTD:/(=5A6D95>dJ<eKg_H)3^+B?Q(_dfG54(8:>Z\[^/Z
4RM9OR^V8/_\ZNeI5L8/55365]Ce2RbJbEU9[VB.TPKAQcT&B;EQZFR3)N4Y@<Ba
Ud&]XQL.,/<IAf86d?eI,9L/>H:&MWMN90(2VBEaX]C=6P[&6ELO1I+<CY;-cKGT
\3:\V.DC@;]D\^J/#(0/#b5A]0Pc8JIZMGZ5WUD^PcgW:4-^8bEON9?eQKdV:Q0M
J[:[/<+/BL@1bQZ>6HI2]^NM:+>6HD);c49?QO0A<_g&)^N2Qg.+S?5<M3-[Q+[G
3cY2=[^YJ-]0DURUS3/4C,\7]C5.4f7PSa/AR;gR->R^0@_41RB+@G7QH([DJ8-P
\OBA@D>]FDKOX/Z-_Ha?:3E<SSR\e9@cY4J(3eD]3QMSVc[M)Q_dOfIYGTECLV.?
NJTQ=OV6D<e>-a+(Ac9b_-e.b0(5D5[QU)?E=))&g6f[2O8A\/cgBO1Waf1fB=/R
.&L;/gVb&Ff0A512b)J1/(@[OYTC=JeDV.MCg-[a933])83HR.F]Ng00d9=R0#S@
#U50&SdX/R2&(;A^Lg=SX3FfC27;T]I,eZdQg0gP)9;MWa_f[gC;M5/cDA+)2[[B
A\_D;M2B@@)&CS9L95J:JDL[,,C/8Eg+(2<WMdfaedVd/#UL9GP6cWbVPRYYP=W1
RW:CU#9CBH==#=F-U;,\9J)EJ]N_dH#4f8::5X5G;\><T>cTQD\XEb[UZQ?C\<.f
YB[<RgP80JG&CP7-@G94C.]>+I&SdJ\.B:bfe4B3]0cW;D(\B^KTRPXS=<U\V-+>
Z>UN0L0V@?:c)JJ)9Q7<a@Y)f(6:0ddS=<.EaFYHd_dQ-(fX_<=E/I9Q1C/B5BNK
99VOOVL(VY)BIK69&@c,ME^XLT6&HP50TMAY#ZN(G4I>Q1HCPfMMb89[N,-^+.2(
4O;TS7R#N9;KN=S:8_Rgb)QZ?8TSA6LAM]KB^/CN)LYGfR[-);RL=1G&Qg7WRBdN
Q^@QAE>7Fd)SEZ-aZSc&;^b5QG_eJ,(6H]8=/),2a_I\RN^:1+8T+00:/,EEe0P3
4II>6VAZD:5,O,S,#CP5591UHNBgG#8M^+0\<?FBfSfOW]:7@.S?S4(E;-_J,,/b
Z(?#Z-b0+Rf0@1gaHT]Q0[\)+22Z@,V#X/gDYE]?>]YeO(FT_-X6H@G7<gPMOU60
>6c1e4]Xg&^7B1[dQSd.(RX?+O];&OdM\_FX[9=IEbJ<Ce#/\b88W4SN;C:W=cBJ
8V^cTcM\UY[,Gb(<?UE&UNe,#+/FHOCYc4g9^AP>-2P;?9<;1BSLbdBCLMJGbgYe
Hd)2b_Q_+0F3MI\.H])b5-.OVa),I/C7O/1XdD?:9JL7MXHO#W6D),9<2:F#E50I
2gXA^>A,:_IKFe4a66PRJO.XLHSLE,>>7QYd3\^R,#><.9YAO)^2Kf_:G6]4KM;N
8>bebe>#gM?72P\6T27Oa+_&>adX8#HJHUW^S\&b&ReM?C@SM0N_-a(&,bBA[,<J
HQQ@_;FF>[?_.0./DYQ)(6b:)Ka1K<743f.;F;I;Hb.7)Xg&@]1.3?0GV6.=N]TN
V\+JVEE?DF)N\ZHK3^HcUa;c2OG1[IOA7NbLKP8/O1?NcDd_eY=LGA>+P=YdU/+K
6?;a^Z5b^#@E^OQ-,D<ACg=A4O<cT6b2Y,Hdb)8HJfIG::f?EOCf>,T0cdYR.68<
:0[]BQ:VQ:T+ZEG+\/G;X?^?62-M6b8a55d;6RWPG8?;=/CD8Ka=N-6(?cAU76R,
=063X78J@7HC+.C^+ZK/NSPBg1,Q]_N^(1TB/<2:AVL2R#WC&1152Id(/=ARTM5M
RRT-157W>\97+U+AIO-?T;(L/;15TcXAVOS:Fee[U8]T>Q^@P?9?:Z7E]<6X?dJB
430dJ<ZGCcY3]#G\_<(SIFfI-gRXK/(7SfDEXIDV])SecITI3KFLC^Be(dT:6,\)
Y;C7a]+T_e1eTMRb)8^(fA,DFS3TaU;3)_;&FHEZ^=0D7X37M(bOXgIS5-,e1X8d
Nd9E]I[<Y=2WRXa^VQFS+,1YB2>=[A0bU-#6(D;NSHYe<Z4NST+24+<JcI7)IXcV
7(Y4gW)8c][gY#,S#9,D0-30eY0HNBU/A04Y]0+Z;EC^7ZM?[:#(?_;+;9C-J59_
1gGA+]6RFd&.6C8\9>bgZ;E?[X6O0?:_:OTaaSfW/6-DBac-)?62g.c#O=;f&U)A
W<[>7GMI(:c97g@7Dad(NS-FHH64eKVWV>R0eF.2eEO8=.9;&:APY_1)31OO>I><
@,?,X[#&;/Z-L@W=A.\11@1FTZSX;??^LX;BN./3G>S(-.W/;L\EQ.(BL>)ag;Bf
\CVbaIbCP\M5E>QW#[.OM@+(a<2SRd;b8.UL2Z;VL=d_@X/BcbDDFROcD0dgTYXA
/3HVU>EWd^\fBYC<D/;[726J6W;PV3.3\=W8FH/\Q-]dH#.[GA[EGfO63AD><6).
eKETIV^(ID^#)EU<M)H5(FJPA?8;6MEU_K;gPX)B05=]J&DXfG8=:1?6_2BT]V,Y
VJF0d1_D?8eeGCJSaMH]7-.Z5,ZKb#:Y0_O-0;I.,gC^LgAg=Hd3D]F;:-_W=R<&
:YGb[XJ]<SU;CV>Wca9V5a/<[(@(]Sb_^E9LPM5YeR5@Gd^[68^@\W#PB+D0GU^-
J[>FBLZ)Kb=ID^2Yf[#:J:UI[0+H#I4)[(]Mc&Q^1c.:/Ha.H3\;.:I]HY9Of6HV
@S[WJ1LY;W0g?+ba[b5L9^ZV=U1CCFVXR4<[e)<4=>CH#-A4;aaOC0DP?B[,[&JD
C1&QL44.;6MQVG/Y=]fa,WJ0eT<@44ANZCf:eO=FM-eC^4&AND=<KYb/C_GXXDY<
BR\GE..KR19(ce/:gV/>.O<aH4&D5A#.:JRJ3Hg4a5B>.K=<-:dZL<-dY0P[K,_(
0J^cHcZUADab&YNE,FZQU76U)U2A\;aM0J1UB#2?NIFCJNN;EbR65U\\:E0NNO)a
32/7)7W@?6EWKP754MGAg.c@VT.[FGDR44A,Fe(2gf&ZX+;<YF_X/UHBA75()DB>
5/@Pc01&cC_/^eF)0N+cMVdI(Td837NR;L9#E.3UP[@0)+dEc,=e/9)RL&dcF,=.
M5fTE/MQ8LGGFX]09fe&MAUEZWc^E1J8NWSVM2geg;\1CJ<HZ[&VQ58KKCV;gH&G
g;D3H\)5?^Q>9]RA]3eM/10O&EUVf;H?g;L4(gN?];\B3Y3KPEQ[(\I>)8U&24=P
.0-)[aLFUD)1Hf1eJCT)^G+d.73e&/-QbDL7&&L##>7NQ(,T29c.S4=I^0;Q&ZDT
./G0I9e<PB<;G;&;eZ822R[+b\c6RUEH8;a)>=:J1M9D=@5LaXO@J.1E?JF0>d&d
]K-=>/;[Z?7\eD3/2UT]-6dU9Dg=b##/BCBe/.M5,19TOJG\E]97?19+1LQR7Y&a
:>:2.1,CMDYWC2C3+X(-Pc)TG/4^<C)LFW3<=4V(@@O>3J,/)W0YF;WNI,2CH>2O
Zf1&@MD&IY7;KR)_@CGO<5TX\fG/(6C.?0A7egNcV-&?-XF7=f(&eCPY4D]&D/QV
ID8bN\^FA8SfJD/GT2;3T)^5>Q;VgP;,E<agHP2W\=54K?Pe?bGgMgeTX?KF+Hed
V#f&9dUaH9I26]#HN4I;1?FY,M@eWLa1g,Og^H\KPP(0,5BMR/YCZM_5C_?P^b3.
d#TE&NUcS;A[BFEIXBIHF/#Vab&/VRgBJ=AS[B[79CH;gTUOK&=cNGXI]<Ud5R,H
X1BRL+H73.bFDQ^&Cf#,AQWbKdXVdgJ^QPD1(3;d_EQXO,Y8P9Z(Y>N&(+bQ>>LT
fOgB6HKbIE]NQ)(BJdV=390MR5BO\30HcRZa3Yd+#22H]6-OSB8@S_dUSN]4N#K)
).c1H5cE/5;f?16/f#3A6[eQ-=eEQH4aP]2#[TBFLO?)-Q0T&g^2B3PDV71G/d^f
N9^I3O_<Q/TP.E;?RC9(/F]L@_D.a>L@cPYD[RZ:,2,^-Pc_GSN7/N<2@=9E<[(W
1/dR2HHTKe^S,-d#>RP?/I;,1e1YESJgU&ICJf-HP.Z7/NQaYDN.G:.HWG>U#H\W
6M>)USUGG_I]J5agJMP9V/)?&NO6J8#f8=d5Q5Q3:)b9X^T#<V(IDW>55#N^Z\1>
H2^MO18E>Z>M.Q\QF?3)=5VG4BdWUBRB#]6g9,6)/:c@_<QaM#@=f&c8,\JN8K_H
)c)C=H>W[[:X;T&+1HX<W984EB1b[6TTCO\;FJaPEgJOO5<a.&#:A^NRL.H];T:b
FKSJ<1BOe;3KMe9-RgKE=dC^EI>@?0.D;Z=^Ra@>,U<--_^OGP8N(50Gc:?f0/FU
:S>ZH/-7;T_51]geVV8-a6[[_Adc5>eD1NV:<feaAJ2/WH,^?&OHN-7U1&2>.Q((
?0;gEe?,8TJJ[?FR/BX9T_=.U#=g1;cK@@MG<RDIG5I#[@1TS&I-WV8UT8a<F.cF
R^g>7MU84J-O&[Z.3/,=U[83E3>BFOTGH:-fQe&B.3&T_39^J3)7(I[c,=BUGQ5B
d_/3V50,]J)D;aQ;<6QN&9U_b1RPb>XWB])AD8IB#T./8;,<1O8MOf=+H5Q>,]/-
)+^FW)_5O6e+ZJcU,ag1dJH29XPHM3J(F+eLZ)610MRVRD]&,26CI-H;=e9ISa)/
]<HJg^7/W>8;[LGbKPPeP0JZRBE&g9P.IOX^?WF;##H5PBfM)@ND?RNJg1&Q.:ff
(U.VCQXZJ6S?gI:^#]gc5-18QJ]/ee:eY6C?I@;_^=NdgeIS_?cdXO>93OL>WO+c
0Y;7@V2P-d9C.:_8c>AaRg4UAFfC5Y\6W89()8;cXGRQNMTWL_cO>JOfaL)O(AI_
3.d[<)GW[]c>EE,<#E>G;]K_>R@0bV(bWN[RE8P:U33C^/V#\+D,FcP_P2S(F.MZ
Ee(7W#)N^+JC[0Kf);PHTUdJ[+;Je24UJM>TNeJZR?\cH\c+edYVS8,[Q6?;fDFX
-;SZH?b7(gWM@0;67PLE4VeX,#&[ed4#F@\dVVBL0/.G:-?-,4QJ-KOd.+W]Ug5e
=E.HFb,d]\U]<3I7Q8F0J@M_f6&M_1\43RWEN9Q7\2GLIX.6.OaC<4>@cS9b>UgE
]#@I\Q9/8b2BQJ;77B,<GgQ\c5cVV,PINIJ\N3Q2F,?/IK)fGVRa\60285PNK^>H
T@1^3cW-^dN#8GVU1H75K/Z&gBN0U._<RcO5.IZ;\Y20WZgKYQK4=\X@^DaMG<L^
ag8.7b#)5/R9]+,?bM--O0SD-HALI6Qg1#JGSF,+9g99DXG][@cFIdE5ZNSQ/.O;
ef\J=J1Vc@D/T@.E)Z/b_&FaCaQ^PeC,VFdJ0e=VGM56f:S\fCZX2VD7QFVM>[b^
(EM5O?.(d9B0b#[==EW=8cVUe@S)#,3HIQG,Rb<]BN\.48]_CT?cG.e,WIg,,W(X
g)2?NY>#G.24EGJUA73NW^ND.?N5)W;6KA]g^cG+dH-VfS=N)Gg0[/e5G]25T?J_
I:cZN1@;2X,G47#.\Nd45(+/6XI#4L2C\SF+R<@)bVQ4c_<V(MEe-Bg4A+(U.K:5
9N=0dL1M[PBJ5TUCb<4?^U:7D]0#Z&F^DN]MGC9ZPd>DM55R./#fJ_f_?AcI9DO0
,c4XM4RdfM=YVJ9(W7RCQeKIOM[,Nd9c8;=Pb8<(TO@+]-\#+LRT<Z.@/8O[Qf;L
eac1)CL&KZ,eG^cN^OHK=C4+\LdKX5]K;Fd]^5&5b4WWF,-c4&X=[f-VM.A_4\S9
+;M?KR+F/:W)7.S4?JAG\4Od421]D@,J\/@5_8)9dSdSB.T6=T-D;:\\f@RJea]V
RPf^eJNK@Dg6bJF@=/9d\4[S9KQOO\gaC[bK]-@1P8V1g#A.P\SJZO@7;59&(5@Q
K83HF22V.GA]\&O#W5Led?_\YW<C1V61(=+V)(gJVW0)Z4]d@@,->S)\?D3,g&0A
[FfT3AbWTT]1N#-V,Y@_O[,A\e+d^ZRTeYgW)(RN,-1#)7#^9)<?U\g\<?fQ2a[g
IH2A^M6G\K2]D@E@ff14JULY16eRS.K,RAB0UHaU(,+3R\S2@JEe4P--08&FdO;J
Bc8#U^;TH[W<,C=YXXcWFeRIR&D)P=[\9Ye/ZK.#c9QG>UB:O8.2Q53B8(G4c9)+
DY=9b5Z#/=ZB3=THB<NI-=H^?(VI2b;;46J)T+VC-82:5\G-<A#)\UY\4\Ug8#.9
Me65B,S057c_7DbU7Fc)K(]8N\-56eU,a]a^:QY9Ed.GPI:PQ([7:S(J[[(QPF>A
Z8UZXC;-9K:d#?A(.&c4Jb/;6IO^^g<^COV3IAJf8G82NNU@C(gT_?C=8PaTKP;8
S-M:^X4(Z:Kc&H+<83Z^KUV.#;ATgKVf?]Yb]a<-\K6EE@AYX:3][LQKPI;Z9+VM
a&@XU7d3G_B\,cG4>AGFA3]TDGT>:9_-fT)FFZJ>[8?\O]-b8eLDX>fSQ/adT6>G
YPH18bPNCJ7)L5g>VWbJ4J+;]^(PbF6H0L?\EeIIL1-f/FMYRcX.b9+Gc+30L:<>
g-c)PDJ,<F5JNKOFfd5.PM1XcQ1(&K]BJaGa<#3bg\(_,8B2O9U&Q=N\2-Bd7.M+
MCXJGBHI#PLV;UdQ:)1TOTc>?gZ98R0MNBW5N3;eO3=RBK3FWEcU):(H2g:G1M9e
(E_RU=>&>H+1F_C-Q<9I8)HILbKc(a]O4gPLO@-5/0Rb1b9=fd2E-[--.bV9^+)7
^XgBN5XNIcQLL#\-e,J,B#:<ML,T03D82G8PDc-7(LMVC,dD5[LdCEGH,dA,C]00
D4cF4BVO:2QZ2f-PG2RgA6g,K(6fYXGb4S/Z^+];=C\J3=Y2O+:2T,(6,RALDSL;
N?[NcgYcB:-OH1.A3X^#VT1+(ffCHcbTN\?RNCA]ffJ8T4Y1gH_M=LFbF4<;[g(7
:TD9=>DbPd6YA2AcXU4\-[NF,WSOU?KQ^6#0Gb,E7<ZWB#,G>T.e^GbBT\#G#)NT
EL<?@\9T4:@gN]G;PYb@.8S7JJODY^E,?GVR-[2Y;[J:B-HT9(^(5..^L0G7e@/B
6L(R1]J.DK_;DS^N):DdNZO57b;\U+13TPW.9^dBgbO_1g4J23P)[[FGF?aGa2\P
IG7SaD1:d#2g(7J=Q9d#\be/:Tb/3C&;5N;T_99Z,;:[GP?^<]&X[>^U8fBc9<?U
566^N>^V;dH4<ULgEX1I+1:QP4A^2Z=+:b^7#2<IbI@6E8[1R5XNPQ(E.&#686f>
J)))\b=JZ0U2]Z;E)][Y)H79_HU=J=5^G,)D5/g9@@[TMT(JcJfdWcLT\e-M<?b9
,;ILT69,#4W937P#fI>M:Tc5>,5g?K^O]D;AM-AVf\A<\f&.9K)U4)\:+5)H=g#T
F<70a;?;EHIV+VZcVebXOK2Q#7M[:MT,W:eHb)df)Y2@>NDA=SZ(3ZL-5)?TaTP(
,^fZJ>8C]BNce:;3(TG.:>EeA90Z_TZ@A#&X60f?3B3<AD,?TC]HH&+C]Z]N2fb;
.ST<KM4aXG(P:-g[&P&#9:#TJ@<&O\<POPQg:BF\.Ob[LJF?4SWD#1F]D_U3FTBc
ZPZcE<Q[g=EN/0SO>)\N4AWc1?fRKTaHW(d]dS3K5X-bE0g^)<;6[F\EFE3.\^7?
?;<@SMf(/)P,Z)b)PDR,aT;]Hb:bD9JWHXPY&CN=VGF&8X-7B/=2Z(5eG[WM,A4b
,UGA9Q>)M#B3;4?R#P)g&QI=?I8ZFBgb7Y6,.G.4afW0H,9b8B[J8#IG0/X8>32W
MZI)^F;#OGW>c8T18a>2F8BA95e=+.YY]7SfdQab@+X;[A)+-[K:\/S&6F=>6TRD
\:,03B>2]1?dfX4E,N/6Ed1J+?B7A8f3gf](<A=^&STT?6L\53dMBfQHR[g+:6QX
.fHS?DPK#eQCRYd1;<P/cRB9#H3272)L7ddRag.Lf7R,Sf@D]_NAHdW10:[babV1
:.D]3F;44OM,@9BBR70Z6QfO?:4C+33Ze>06U6.SEW3H#8RKg:J[NLRg<+C\67B3
=^-S)KJJN^51?CFY#<LFS:8[e+_B,8)4=)=)[058#PV^=7Y&6BEVRX7[MP-[M\#E
1.](7I]EA5DOE;>J8O1,#bTe-:DPJ7aV(WCX\3FgF:A@.?+N1\:g4^X#P(=7eE+J
),&JKBXA##L.9JP897fZA41\O8P[+NPH[I4@13\R]EY?b8S6e?/N=,#S2:VEAcJK
;+]FN62_\;MZO2V-AT2adE+VLQ#<\(+T#fQ8X4&87DTS\2T;MKDU#KG4HF:YX-]:
GQ]AdZV0785Y?#5.8^eD3WS\WKdFC[,SV[R6]^a3G?PV;685&H>YC>AU)5c_[8ZH
)fKBDZ3M/RBPW.3BQ-<IOR]AfKJS)c)V8A0^aaSV=C:TD65bE5DPPRVg<P&0Bd65
V\/1Y_XZ=2(,^BZaffZ0B]EK]cCb56C3[#2@TfK1YVGUH2L+NR3MU2b#42EDJ;gF
:63\-G0)8gETMD#+Zf/b7K[YdO,B)V.P4U/#1+3<;#2Cfg>cd_7I@a0;9@/;L;dE
JEY<X9M?T(HaRBg7U=(&;,TJ.Q3B0-NSdd9^HcT@BO>97ObZ7\6_9S,N7.-6WJ?g
9,N&DEK<[e4&B18\GUMDFZIb:/@8YIKMIRLWg<,/4,,T^6ac1-Q.U5X-6]V\@F@#
&RKb\M(G>0P;.WFd9;R<9@f\EaR;(0]X8K>/]F?0KZ)_O2-P?OaSgZQA>AFN(-/g
SK]N?NAbN4gJ2<P8a,3O^e3L7Z/LWgF,fHVF)c4>;DHfWd<Ge=WFRT7\@&(H&YQg
T7N)bVQH5B;E=Yf1La5JB=<UaBQ[KJ\TH#g(A\P_04aY\&11N,4g<>B_3..f;9_R
5V-D5dRd.a6G<RJHRabX8C3aGJe4c_.gHJH)N_7:eZB5:,F@;CdY3e<+f\GSS61#
5M3fdG4,#?WK.BVcPZBB..f55NI8WWZ4c>S.\3CWN>eM/^YQeZS00M,366@]PSPQ
5-(S&W^K)<g7c\E)&PUg(?1P0:8V9eTO(Z(F&FQQ#Mb.MDCR2ZRZ0,DN@;,PHH^W
^eec5.MCY,T3/.OCEX49I5-@ZD9E&cJJHA]G6-Y)M1Ge3F_)+c+I\ZJa&_O_R:NA
X36Z)HTWEeN<K.dGda7JFK,[4cL0<GP3+f7g(+TCPXeaCI&JAK;ZH]9>GIZ:YCO+
#]4\X&X_:S0H\TXHF7^2&(OeYW1]W2?1HS6@#0gBL-&9@X-1YP>HAOKE5GPQ22RW
=NRW_9-Jac(3^)35gB2Se))JZ_Q)GWaZWED#XMN4+/Y1A<AY#Ea@d_Jf4J5e:fHX
_(d5ZLL-Za3cYSf2P.DL8TF4Y=?N;Uc1TCAc3+<FHY37g,eTSfQ3XK0^^P->3.=9
B>S&&344L#)8Q@JY3;RH9BcUR,]DSSADTPRMA>0aZ\=Y72R^9)2=R>9SPQ\<9&]4
c82?^Z\.^;f__#L@Y)8+?78^DZE<Z^(#]^eMddT+gbNGK)8Ud?ZN+>HN=d0gVM:]
K?b[]eMMNUTb^9\a[TM]&ae@(&]IXQa4VY&8LeF],-&E)P4.2T]SD3V@TbS?I,,E
LX4gBV17I<[O@T?X=YW,R5Q:78P9\cg.:256aa8Z;]F7>[A?OXD=[[&+8WO]VSKY
RgZ1WOEZ+7ffV5aaAPV]5K([OeICV5YPJ+=WW9V@H<FR@\c=#BVcZN)5J@cQ_5&B
EQH0>7I8\FCb-ZAJ\HB>^)4(SU5dY4#GY>TZ@DLQe>aA-DcU.[?C7QAG9=&LMfG:
e-A[HPGF-]_&7>ZV,X??)5IB&_IHf?J&PO&&?,JW_0UUYfFF\LaEU,ESA2)_TVT3
XQE>2=Nd0aJ7;(ZVbJ:=,MS2K6YP.;6J^SQd58Gf#A]0fI-(S-FRaO#2)=@;,X2X
L_YVND8)M>.CE.2H?0@5YG^Q[0bfD9^Veg?1?g:@7Q_c?AOHA5ffd4)E9;2SZ4[L
PHfX+JX=<T7cYIb==Md:<0W9L+:NVF)S-JX.WMPbeTR7DE+UG-4/3/,4[C7fKM..
GY?M?KJ5UP@eR4Xf_WXIA7=/K.AcOA^dI/AQ4d0PaCZPa-&eCSLF&<85877V,Jfc
95fN)LYZ.g?\B2=BC08&7(cXKA7SfGPe_&CBJ6QQ:>WVUdaTPg90VG0(F^L=1NL8
@Jad9V6&NJEWPdIW3Nc<8UT84_+RdPa8Za/@@V3aV]6:0^e=eDO\a8#fDVb7B_bM
(:-b7+67[BZ5/:#0N4O,f\EgXF.;TICI&&VDcL@H.W\_PXg26D6BU+dRY+]2MRT\
;BA_Y45^9P^-PbS_X_M;/6;WL;;<VHdCH&(78H:ZW)_I#UXK9OAK-F&]WMY8)SMZ
R6DIRJV=VQg.MF?&<4e?B+L4+5<g0abf+ZA.66D?X+,FO_?:GUEX:@8,)3G+_.\g
(Z;YgRc(JE/dN+f\1FDAK4VLT,E&-b)JLP-)0BO54+dfH>BHGbEG)\U8^;3\cW6)
68L0_#Z_M/X@cOU2TW6Z6)RG-HR4_@[0JI)#26=D?1X;CQa#7K(U]EGA<QD]:Nc^
XI-LTag0RCL\I+ERgf0@Y.E]@^CWR[8^<QHT]b?MGgNJELMQ@RORb@GR[;,[HG2Y
Vd4HCY0)MVBVOVF/O1?=VaSOge9JgYJI&#5OfFA]0L\<:_?S?@?VFCOY8\ZDW^YM
_ENJ;c\3O6_.^Q:IV?J&Q[3S(W+MHY:[X57@7-;28E^LIfb3X<b]5de]Ne_M^AbQ
VAOXZ/2e;IR7:+Q0L<1?,Uc9g(4OT(4:F2-)MPC8aE;#Ad#)KS?b^HeMESNRdd>P
\D[<_]8;gT7DT:.RV99E3X2cZ_MReCI)QR;H.dE&K+VI)JY.:FG?a@C)W6VN9/+B
&9GPe@4MT5HdA1<dg5-[84(dFN]&_&+2g0:Ka8FeC-B-,dKA.g,dPWddc)W\S9U7
7<QO8AQBAJ7ZLD7F<?cLIe;ONP9KaQbAF)68HB>9/We?O@;]5L#fWU0>AR)bd:S5
Z_=]Z]A4Y)HGC]U#5<YI,\^_8;0ZET#^-ZEdEX&2>Z51?GOBfYAN0#4d_Q:0XeM[
(K\WSSFT4e1]K(G19H0aQ1,#;H[>bQGU&dJ9WMHQST_@9QWIR;<IJJ@)0]71Y(6T
b_8G-IaW,?)A;KMa6dK[Q.J0>07S-QfaQ8,1,_LI.?O?9cPG=7&(8WXK+gaMXb^D
@a4N#)#8+gQ@7bHJ6(a?ML.c.0;UIKULd-#=H;UJ6WJa51P(,[YKW7<J.FNLW>X2
L9cFCaZ#da^[CI;2W7.;;=SI-B(P[:+;G<I?+2g>geWMM4KC8M,cFd3<7>C<+J4L
+.6:&O/H<#,+DR0QD=57_7-<PW2Z>d6[3?E\@e<@D+e;RbK-?H)ZAEbMPf,<,P79
E6=6KAeD/(A.WP</Q_e)L&X8K)]+b#^_-JUg4]M>YM5CKV5\#(WZ=AR(T7DbQYRO
?)CUQ-48<?gTU5=(<S-#@LbB(@(\4R3cI#-F]<DbA0?6&<V?XJKC7TR-PLPKbQ6)
BSSI+Z.1ZWN=#N\&@AACHL=.;g5B-1L;E(\FNMI;LK)J+H\2Ca_9)gfQf7?[=#3c
?g5[TNG6:f0?C\,;:<gbOUIT8ScL9OK>c>7AC)/MaKLQ.cUGG5EHBO2<\^LD2,[3
5a<T8:TJ]J;ZTa7234)E<+e:H\&;F_NSLbH>FQdACc:2ITP-KF(G-0.I8)S&.>S2
<@AW+=>G>H?+O=c>V?PT8S7a\_UB1:^f0g17YG2SO>QP9+[-A1X8NP^K3<JCVJ@&
f5N_C/AfdD(-VN.9bF;PG^Ha&5<^EbL85BECX17&?/.<\@@</Kg\.OK:.&59PZSS
d;3<Y^&INCT0D@gcN0d>Yaf5cAg(M:]9,O9X;gEK]+2cEX?#0/@?,b8\fDIF[20>
1,&NfFZa[#892W]JDFS(/)U:@\-J>gA&S0ZV:ORD^IO3CDcf?.7[GW.P;?Ae;YY0
H+Y0NK9bY3_e(B3,P+84Q)#7J<9:P]dZTUeefVLG&MfQN1\,JJ.4<@>L:]J.3]D9
O0e-.I:?fWa(5EDVCDNe=597+MA#4@Z93O(0#TB+SBEZ8OBKMS@V#6V.(H7PZMg>
[@9,@_c212FY8I7fI<TALad,&G1_<1:713/SCRgS<d><Q,&fEH[)UV.F>SWE@UKd
]QZXUeZR],+7;B73c+/+fXSI?O7A6<b[^T8:YX695.R(e?=7_G[,P4YV(+4^5?4V
^W\b8Y_5_(VER@&:J<g[Se+7&JR@][[>6,#W)HbF#g<VM.>WLC6Da+3b/9<)eXDB
bE4167]=(aTRFcM.))Z:T:E)W8S-]5bg9XD<<9C\ID2#?5ff_)UAGCINJb#VPBU1
<H:X(2-7FIJM+YL3WD<2<=FffaYUPLCU^I(IQ=JcH@?K7VYFbZ6_ENJ&_.^0VbVT
@D]?_d\7I=8?F1N79],_Oc\9Ne-_T&)VZS4;+YUKC;3X_L5c4]EIM.L&M6(IeF=.
W@8SNaJ_TKPNT[7@&]#ZA,dW8cU4AUH]Hg]R9.)ZJb5cLd+c6c[W<+XAJIBGVFX@
aJFaV6cZdDe?XJ83dVKA9QJ@E4D<a/Fa,^XU?3.P<=IQWN][J]/+Ma?^>/:[[5<+
CPE55;dVK,GA,CO=@76#88S712;)bTfdR#cCT:fFFF)7UU])VZfEHXINV.^YFYWg
b,U9[gLdR9?M\<U>:AKB.Ne@3YVf3JcJTg[48f600fgW>L+&-AQa_cZ,A\GH73^4
C=Vf@-=S>QTU1T72#PKCe)G720.@0g>^]MXa9#Jc4eEX[;2A-V9^Af..7Y?6c@>6
)7?N,\,S,GY11.7TJU5D1D(;e<4QZ,=R03KA#N+bLbH.?\=AH#2W9GN0R85f_15b
;c4X1^IXY8ec-b>&EFb(VN,3A2#WNML),RDW=UcYgV5VCXbgTe-bQB<Sc74(+&EI
QWH\aE95@dE>\[6I040ZY=5PDGNQe:E@#AT-^\;.ad@]CbU5BO7YYT<]9Occ?BKb
D4W89Q>K0AM92,_NE;A<IW=f<>BV[TMdU&c2>R==b\;3;^/O4S?/DP6.Fa#B)<b1
;6PWW.9b9P6=35PGJ;,C6JE@63F__LZ^4?8A#@J/(aLR;E;/+BGBMa8c=8Q#/-_H
X+#2]XfPCY6[4C<LQ7Y\VT&.aJ3b<@E<MSZ^2,+f(b:3?V>OY\D,SM2+[8]0fE23
ML950]?K/3:A@>()b6M@;TfL+YF0/_(FS(4Ja0Y2GY^POH_c)J0O&(B63Ff_-/.U
5G:N>[+YVHF\LD?MO^5B>)NNUN7VZML:aN=bf[6W356B.),77D;9,3R_X5^gSC8M
/X94-W1U?.fSF2<8H_UYba\1?B?4W\fb^8M\9&O410XQ)IR&0.S6)=[Zb4ed@5Vf
I#:GZ[G61HAJ]);1RZDTcH3+;5+_;ZD6)PS#\K@YH)c2]ZDMHXdT:2^#c@48JR<;
ObK/EGbX4cgH,I#/H.(JK[(56+#-L0(+AaIa#2&BcE5#<@G?3(X/KW5H0&VaGH5R
U-V&R3@/\@^65#=1H[b7#<.Q0P91_8cfCFa._ae+e8[#/OH+@a9/:2f,/C)FT&CR
g+4c/G6WgF9c;gVJgD]GIKfP#]LQBE^ZAa[E</#;6CaK>)WE1PKgXB<6F/#AK29L
HDWf<^9eXC7cJ6:#d<:9M?Mf7:EMEIKT9WHHEM.ZbPRCMWJUH>7VGdJ0AKE&E-.e
-W2NQ^-IeJPU5LD_cgYNQ]d@YF@)SE1aMQNf>[7U_DdBJ:=)J>A)V&<7J9RfbF6<
+KOa<MO3=HZJJ]8:_3)2(,GKV;]V6+93eT5ff38](XgO^=L.Z2KRf<]bK_)KaQEX
dV+[W;BfN,AE@X0T[8#)PYe)?HR3^&)K_U>OD#\1.JZ/.MAbSLbX=WF5)477TMWc
L=,GO<ZRcJ?:RJN3KA@/3TUc+S5BeC[DgT04_aab<2OM\P._NeeIc@-ZV^#53)C>
c;YFYRF8d26>K=8GCB2>R,F/4O)X-0Ed#5dC;,Cd-[^#L;;A&aJ.?AI)@MR[>I_W
N3O1+C[#[6VHLN;KFN8@=KV>,<_,SXG4a)6Z3?=Id5Q6=OBUERJf@7bICA;dGUH#
G&>TV@U^<2:OZFFPF50Qfb]Z)fYg6>L@_eaVaS.cT6H2+V@>B0(g&?_8WAd3AY(S
L?R9N<OZga7=@]gUG,16DT0\<gAeI;(<0:\W2JBUd[27a@T2cQcUYRHSUb(c5[=2
.&4<SF/Z>;/-GRTT?8?g9>X10-NH<c8U1E)QFZM>U<I(/a?9O_5EZGa3K)2K[KFP
EK)?(E#5#f8gcP)DWDA:OHK9F<#RFOfTOXKM#V\QHQMWUH/#T]e7E2UQHGO?<S4B
Z[<X+G=?2J3;8^:R]B7?M(1#U56.N:OR1F0b(A\ULLSUGGJbL/N:Uc#d+^Qf^Fb)
e.)Z)BeA0g;2C5b_1e50?b>)/IJ2;d3[1(c/M5(GbOE?>\J300P2Nb-7H+b2P(.C
M5Z:9_P@UV(/I(6V[]aUNA5VK,[4D4/A5Ceg8(gUEKNO=T5;G7GSBONFUdF-1R-=
()g?UAS5g/^(/YAU0DQPF#MM:gYNP#X..aAGVA#A^4bSOeFUOeDeQDRUCA0+:Z<#
\Zd2-f33<b[GY@dG9(>3S/?ZdCC=#B,;DKg\0O\HU.93+ZC<09NAP12FgOXb@?f0
c0cCJ>66@DQ..\OR95K(H&FV/XKP2B2CEB1L=S_[/.WSE)cUITPN8DGJKNX(0AQ4
<9f:HgOPe-INb1a98=cfF>.,][KaF@ec,A8PbbYMA&@eNc.IE.FbK=NV09aW^,S8
@E^2C#fXH_TVJED\Oc;?Y^>N=\V+.C34I4NaK=B8NJ3<Ig&:@>3,X,JWVL5<AM+0
ULDUJN@BPc.]FM(+g]BEQ6+QPVW<2Y[Y30<W]R11Z1Ug:(5HM3H,d)[[YY58FB3+
b0L(C;05b4SC[B7^ge\IZ3D<HYa3L@OLUKCZ\D:JN[64SC@Df4Y_A[R2bWP&H>^1
MM8YH]5H:\cf@END&I1d?6.)G[8W4ecA7@;3#LG((+,aW(2/EZ_5a0P\8A<AF)8c
LMEURQ6G8)M7A=_[C@@S,DL;Vd9R#2@7(&KRV=6;/@F35\(2\[R,;U)?9@:WVJ.T
:d?-745UZgB/Y/a4+4@\L/8@YD,bf6H<GeEZHSTa.IMG3agR4PdYc;6aeQ78(X/#
dZ&<De_RQISKV;ce9[4[OQ5.E7ZD;O[I6/cf[W&S1>7M\aMXg8E#@V8Y9SS:#1e,
bc9XbW3\;7#721b>-/VEA/]]I<>N_R\#=Ng&5DG7(fA)8_dY,PA,e]d2.PaWYJP5
-c6J/DQT>M2C0_3W6BJ?.HAcVG?QRc.]V;96g,Ca(UP=04E)R/Pf;5K^<C+(P6.d
RW<=8AMU,10:(.7^5GPVN4XKXXaZe&G0R0LB9@Bf;&c6DbJRZW/G+@H<UGXfO=J#
1],8NSQ76[YD4](J,V@O_62(H[42c=[JR^9WMP0&5D:KFbZFMKeM8]5bF12[VeY&
^D;K)T2TW-0??8,HQ(f>)3K(0LLEbQ@E_KQKMI9JZ=Sd_AW/aG9g;YW\4,bF:R.d
.aM8#H2d?,c1g^<J]R9c2A/P2;M#UDD5YEJP+5IJV)8aDE?-bIa.A1I642-_b[cQ
3.@^0@K??^_6.>I8.dD[^GI6C3GS6;@-8cXZU8:K;\<&OS^FJL,>2:,F7NRZ;Ce0
K5bBdI8NJJUeY@Zb^)A4=7/[L_^G[=MDCTHMQ=#b:c(54RS17fMH/_+TVZa97cf_
-2.1?YaA:fAQeacfJ4AEPPEH#P#B<YUcfKfM.7FgH,GYECXK1e?)de_X?+:LbVF^
RX=Kf+>+@)RcSFP3K]3MLfdH^JHQNS8+Zc2bgeDC)B;8P[EI@<+O,=\,+536\Cc@
5Q;?,Bfd?b<(J23-49BZZ^R7E-9[Fe#eW-8KI88[?TI6^LX7U]RdA7[SMPFNbd^>
VYWA9eN306[\9292P@EENEe?#c/RKA<\?C;BgN[O3JZ@aQ,PC-S^?R<5188,G1L^
=e+&M^7U,HETX:^\gN_Hd08OH6LY.N,@fRZ?F^FB+/YGGI/KA2O]gD7=c[O41PG.
S#3IPHY)<cc\I7H==26EG]..EdF(-Z;=BR7WH.d+]9T<AZE:(A>(_M+X_Q^ZWOS-
E[Kg:??KbUYN5e#7.0bWY(d&=6=^&ND]G>(WL#YP=,KJ>^0+6g/PH4V_,.(7&/VU
B.]Ag&10gWadKO)-VXW4.bJ_cb\49=PCL1VdOL6R#bWQ]8DdgPH>SeXYa)NXA^.G
^JC6XVaSe,_N][W)PLO/dBLM<B=PRMaX;8)MBc8U_7-fZF4NKC7KaNSEc@beC)3C
1;7#A;7.\J6NTVSOgCeVT^L3fO(Z/1RJgC7_@;S]#JgFYLBX+;WS@a/EaZ043_6J
QQ]9A:U31cR+1KH;.b2:7X#C&cCXdV,FH^M78[f;gGOV]JY9>eIUeUd1+c2CNKM&
TE[SZLM9T..&aR9^FXDS>WVTX19WET6)<>/Hg=BY^9:7fRQDF=O9[AQaeAZ:2gZO
;2L]2\SOd6SSA\VC(XE&@X(#\2^\#MIEH1fT;[?dg(J1V:]aD&]7]OVK7GSUG:M>
3I_=_^KC7I\:::3&BJ#344:Y9?Ged]?EZO4,UZJ-^F?\Q.cd.1d\f0D#WJY6EFcW
VF#4T5>_d2g@>P0[6bKOV_3D(>QGI0?PR[7ZIT]bLCa\R3BWNH<JgD.cF5,/bbIY
QgZfR>dPFJUNW1g^;(g7GJPb+ZEW@?P:S^4N<15#8J-QZJeC>,1/)3N]YDX<5He4
ULDW7BaHb-V>ZOa#MVbO,/N.88C(TR\6/\c8+;_Y-7_c8FQ0+\1P#RFY133KG>Td
,IC,&;PGBbe\NB+[0^>R;/=C]?8INXdY+/>a8^ML\?A.&[_c)\bc1#P,#3YU8L<@
aJ.[J:L(^?)9+GH\Q(>&F8JMEde=RDNR/<T.<\4&=3T(;J]&X&3^<A)C&@<CN(AT
\ESI;g?AIE?UBTFMPYA<PA:0RS:2W\8@-(SB2;=CWccJ7(IFB]N3Z^fadE\-DeWW
c.Gc7TMFPD.;>8Dc)SE?7@F24\T;d=&RB+21>YNfLG9U>eg>QRW\U^YA]8b+>?./
T6OW@F&BFI?@]3=(J872M><S<.c+1X0;P-@Fc&&(1TY;&W94SbbM0E0R&Q60J8d]
\.2bN#L\M\TgRRQ[M[S.ZT/?eS4e#.;e5\6,b/@[6:6^fg1NY#WGN4#8T#+4NJ,R
.T<E2&X3V;WeZJO[^bJIabQDM?_[gB-;YBJZ<B&E\aZ4Y7VC]b_KREIYPaXAJaNE
\/5.NF::,g-<N;WN]Jff9K,OCLB1CbW4Sa#OCeLA8C;5WE3\].N<?>3DLM-HKZ;D
.#UL_CM3.2_3I-b<SYZ7#=b/D.GVY^-/#U58If.I6,(0^WPE97_6(NaE29LbA6L.
=@0C3KO6GZ:T-.^EZ(V242([V?_^9c]UA]G?U&N_O5TcXZfOb[WJ>L)P]2568;bE
@AJ]]](R^VXLGggL#R;)LBNXb+E<6UX31,D7bP.6_GYC((O.Q-^SNX#FHc7]MgJf
SB71)^Hc^e\SOZ[#WMJbAB-Jd,bVB,ATS<FEEJB(IH,?DL#K?7IO(:S2],eaBeY:
cPIB9H4+ATOJKYD)=9SN)@Cb&L03dIG1NdIC@17b+O=\5S^SDZWBcc\1FdZ92TWc
,D37fN,58fSf7Kd^T>_#b]MeUFQPYG].IE=HMaWC2ca)]fb<bJ_[_a?Aag,C5/38
K\4++@[._aJ\46XJ&W8G,/WKB[@&aaT;_(>FJaD94WYU.CbZC?_d4),7)+.9@N0Z
3VfVQ3O80C^O>D6(eM:.-324[1fa-RN,PKOSI#_3g2PC@>b8T]J\CaFP,-BZ=#?@
M98WF5C0L;=A]a9WG1W;-B(VcZHO;@V@;bX>B@0b@aE.HM[CBYg_).5g<D8;=X)J
a8f<FB3YDgR\Md+DP+,.&ac5)5G[1QT\YfE788VEC3fe#g;cd3NV+2_cZV>U0G6g
I>]=_.AdO&-?3T;FBV<(g6[^@+4ZCWHB5R3Q2-H[K)RP-^R>gf4(_]5?e&d>P5O?
JE]Ue]ET-->>A]Re)5I]5T[N=(eTZ@^QBTf^6VX=-Cf?=T2(5)WE)=#7H?e(?]-)
2H/EULZMLQ#UQUHFX?Q^@dYTQ=(#7?J;2;YI=HV?,O,N6eZO[X.cHa(99MH@@9)/
NGJAUIe1::31b)LT6bLT5[1]#QII-8T>VQI#K,YZF]20/W,J=--\/f5IcSPEB_=_
K0?31YX^[fOC5<g7>7/T^ZRVWc_0STRK62KMb>&&fGaK/B1P_AB.a:2B(a/?E+;2
YP+^VD:E+GX\55,b[?>fVf:ZC_NZE).L[A6E1,1@@=(&&L/27g<4V2N+EV^88>eA
&,F\bd#:TSQ]]M>_L,.A.I,;WF)\Hf-YMe45GaN\(LSYYY&J?04OAS8f58A?ceaD
E4IcO8MUf]&8-XZZ/YXH:+_g5UB)_;,[JQT56/LQI\ST,_>IYY/\T.[@NC#)56WZ
0O+]R,L&f/Zb]-cZ^Xadf]e86V]JSOA/>gA;;.<)\,6O=?D=_F@dLC/1O0;?c@FP
1D.]ICMFF)X8X4>YM:_^^R<W8OedBG5F<7c/3B,\W]@+^-/AA5UXHH2dE?2<d&R/
Rc1&NQFD)#6QP03RGO4T1^)9C^776,P:.B10#RU<c,8I.X9-#dNVFC(98366RGG/
=?F[F,POF_YU(fSF[L=7OCQBM><,-^Y?+FCBCJg;a06#/J72O>(AETC4EPe,=SYX
F16;4ReY1)CaZa>PP@[2:V],H:CFVUC^VHb<4).].)Ad29]BbZH1;5DWAIVQcVL,
(G0P]5V/L\E--NJT-fIM;1UGD[TJ=;@A832SQO3K[6AM-b@bIDUL@UdUNe9;0G=U
>O>:2,5Sab(UdXVG0[@EB8e;PLN8]ea^[77#S4,[SV2<XgXf(:FUg^(J0<W&K5CP
<d0XW>@gB_D8>,;5I@E_6L5cgO)-S:@P5).QMG/fM^CF]1D:D,M;dLW>ePFg.c85
U\\LB9H1]5G-XT6<gRN<GfeSRIO3VL;T@:1^bI&5ffP=,CNd#B+c>DS3T,)[a=GE
[f.UBZ-[g1Y94?;GYLBDT-=UA)=T(8H-=M.9Zf^NFJ&c>;QbbQITd,],FTbZZ5B_
\2>fS38S7g50SEFD&.RZ#fC\5\I&,1(,QP4)LB\??&C[BDH8d/1^KJC8DHR;(N;g
4<W,]?O(MG4[PF9OCO.R<9CY\EEY94d6aQ)bd[>9d\?bYO=VbWJ2c4_5Z,@0C?;Z
.<_1AR(MR6V^^GBF]ES.-Y1-b5@)P4]\Bc0SV(a7CQPW;S?Y@8O_>>#/81YcGPZ/
]#[+5c??2/g<d]0]GgXg9gC<Y[@L7T2fLQF,7.<8D]<^0[D4WE=KJHa=AP#X]+DS
IQEf)_Sba@ObfS_DZ_;TaY?P<[.R]YA#4[E8V=MBA8IC;>R3F6ea8Y)@Xf+dW/&3
T72?6^46WG^fZZLa(UQ37-#+?_HBbC&KGTa6:PLP8dd0,dVDb/6,eD\NJ1QbDADd
2@42^S0<4MPR&>+Q>OdZBH,T@53VII5\5NM;(eV?))<TNF>=F=L=EP1bQG8Xe(U=
9)GY_=\5/[5]_H0Qb=A&8Sc]=4FGBE5CbM/&).J\e3^2>_\P5D8/3S,?QC7cI.6F
EgH^>HcFb69b_OUCbT\WEL/8G<,,S<=_]U=C.UF._:_-f(3ANNQ#9=c[8B108E1T
f#E1,FbTW+5Lf(]JL.HEa81&834;NE,P)@JCJ#Tb#ZU6Y:cK3H[FZ?N.J#+2U,7B
<J9T3&>;1:e=]TP6?:,-+7;TF?U54G[U:V)5DI>1>d@(BAfT._G+J.1#5ZHGGJR[
N^Gg:#605We0C\,2=J5.<ZPWQ]1+EPA2gB,2?<Ob:D)9SN^\daSTW3[<Z0XfN@f@
K09.)[dB+;V=C]T<ME15[>O.H18>)BZ2-#D,]]Bb)<B8GYc,X-S>@KLMaM]S.)M6
((_F9<d8/57;LHVd-0#(8QT-]T>Q;bPKYP:@403&DBO#O/DF+>gJA<(+3J2==_47
de@#+3]5ZF_gcS:4EHYYT)2ES1Dd?<N_6:B^=Q,2?90CL?216@N0OIHSb,>DaI)F
N4b)5>AX5#IWdCWcaLdW1>8<&aN42:T_E2a/PZ,MCeKObEDe()#)[3EIBOe(BHb<
YgW4CO]@-g#bUX<GdfSegEB\Je<Z4]O&e/g8_6F[VeR+aV=TTG0QSR^M5R5A8I+(
X6aS<0XW<1X=H#CB.LF0O5QYcacV;26Oe2Rd;X,BLDP+@a=Re,-VZ2G4_>AF9&4e
78>387X?0:b161>XO)LF.#Sg\PaSSQ^8,L0?FDM-OP?U3K[E(9L4@X@dZ59ZZVG?
\94]LJ=79[;)BK=,)bg5&P4fg.dGLZXb;CF[7\A<8@9Q@KfI?3,O7a[\/V.Z<,7,
PU5T.&2)+#@fg3T1QNP]+5=KY5aF>[=]Ye;84AK\VF4^&N:1+aK1P(9_J[906:.X
90P/cUNOGT?TeK8+DTQC,d1-&B<;L--367Ya^D4AdT?G9>;<<2NBSZNE1J[HV6^0
V@O:C):&XKHf=;b,g1+GPQOSaHD8(H^bM.)MOODRU>F#:GSDf:\a(g&FKQH#3X6J
JWf)dJYT^.d)cOEK<4C?YGd(F<g/@+B;d4SHd1.FHLJL/8Lg&:97_5]T-PeD.@3^
>\ZY]7J[FLeW;C)@JIP2aWK^0S?&#EC3Y(FG9P.>TF9g\WU4UI#Fc<9DEI48^d:_
X4-@dWg^H76E<\=7C-Q4+.<Nb]H9B81BW)B+2@DJRUYJVNc>D<C#E5E>..3\eB]E
@;GR)XFXV\QQ(0-^>H<_:<F5#^-?7&\+>UBFa;?(G1Z^7f_2)E.]/?/Q^7g01>QZ
>[J(^P_Ac@]0^gCK7[G:DLY0dG.I1PM/W#Y_ee\PQ0,S#C5WKSD;NJ.7T(8_(X\.
V08FBV9<ZMLW0We6Z\)Of>MU-+O9@K>--M17M>cTe^=Xd.V:2NO6H@L8b;P)7OGO
Ace(IMV9\4;VEH_15)9:NLLdH9Vd4>USb=\O=#YS3161Ie+\9769.e>eCO)=dQI<
=N&-R8gLWR2gH;G>ZMggc1\?bN?5_&c1B?Caad6Ub?cLK\^Z_EL&UIIA[EUWgE37
X-K?W/:HX_S+;WVT?DY&-ZR>Y4R1YWON=B>>gDe<E,SPZW64fbD2Z6GP2a,4<L>F
5;MH.<_9IgNV(?5T)C<B-N.-J_C6N-e/,-LQL+QRe,2?C+B#^2USQ6)1RG[cWa#7
AV^TAST0<0;_ID4M\TW__OKP+_IAXG4T8><Q:/_Wc1+F^cf.20/[d4)^GcXVAR]c
#RK\f2UYgV]c05M&V,.3BB2CCCFPIAd-.bI2W;67XIffUY@I.?AWI+_^cK=,W&R<
<^FeaZb6e_,\9Mge+-b4-0W23N1O@&1R:b15=c;HZF4B/ZN-EM?;F)[_T_3]A+V+
OcbL2^5@@#\,X32G+aXI5@4V]BaX=&:O&Z,\g_C_2TWNN=#7(Jc7AVBXg@B^YBe-
[<dWabQN)+98YREWLg+JUc..ZM59ZY(OGd0<DBU0G1R3Wf855IJ33.ZG]N:3a)D#
Z-TF-P?b#=;YDR;,Z,Q]8.6Ae457_,,)9#\b1]T;VW@aRCB2(]W-.02._0,MggOX
A6&PAT-92a8b2<:GO;IS/NWR]756E^3aTc&ebNT>ONJ5&XN9]F^ZHOS[)12H3fH;
>TA8]@0AdQPRd=Z<X)VSW(ICS;QZa8P1)HY87EX&IEI_;E\0S[3W;:RI>T8fF_ZD
E46<(U\CcM=K3MVV6P.7g4J<D[#Z0OQda_FDL=c7YJGQU>-R>K5FY/JPXfc<^fBC
P/I>A)\IJ@G9;MfVGU__X]6<=HKX/QL=4L\.Y<0.fR4EOOSACb)OG?Dc1E901eHH
O_ML8U-C_?7g#9H:YgS5f/\6:DRHNXP^^a:[Y1C6(]I<-QQ\1G\L84S74YD=-]\_
OM;0fa#^d81L^Y^Wec]7c9Y>,O;:-#gULCEQ4dS&,Z#Qg?,X94]&b0-a&[bY<f29
bX4WJCU),ZCK:^C+X(N<EdVTFF#=^@:7M>I=e/DB;aB250\[BFAbg#]<P_O@X+;Y
I7OO).W2Q?R4^,4f@g_MJV>=&[(ND26=agI,\JU)fdA.#00)EQ1b#8D70aH92)&2
e&\(/IJ(WVed.5<+S[;1#?/OIebRZIGZ-F3:.dVP@42WeJ.2-f5d/.aH=)N(ZP@.
CC4D)6;;.X<)C8FU7[X139L_Ma786:CYIG0?.TZP2PL52TRO>7HMI3T(I:K+RNN/
+..[OI5&cUF\^G@F).MBL121TRQ^4+2TG&4)1\JMJSABfUX_8NII^?68=;.DV5eZ
-^8M6[,Q>:MR_&9R\<B^&YC[\#.-/T9(I0(2d<<V22G:;&SL5d-.EWaa8dX>YggK
_\1/<@,ZFRI^QZM2>OA_8a0?0]B&9/L;^0e0W];X62IS<3&OBD\fU;<;71HeAYS7
CA-e:.+@LGH:=b/?5d0K9:8dDSE]M>#^gI-]FCZ@:#I/5eP6-FB,G41&gUSW.Xa=
V]S]I;&00\;,E0.TD^T8dcS::+4\<PWV_0G+?6LGJ3)F=MN#)<BMGe[7RMI=cQdg
TFMX&#HM&N-]]X2W76b,Q]T>Y&/F8EK5[Uf1dZ+694&0P6F9Q)ZEHC:BL>_R9Z91
,DKZg.NI9CF>^TPN;c8d;[(Xg&\O];_a,W[d^LcXY@V87RgU=E;CI0dL;aP4RVgd
S50OcEFdSbaAKJE)@U2^Cc^&0P:L7[X5Bf@fLL-NV_JK(=Ac>fM^F6TKB2Q_9Z\5
)TXRFF#dEQQDMFR:@/Me=3+3:cWY@bQ\7[7Hd0L(5;F#UVHbKgH.]f?H6([b.4O+
]VD(aPa?+1Q<_:@6^MOU;b&a+XFK^-B&.8dSdN/0RTcG^XD>-J.19P>2R27)Rcg4
.0;5:;UA?P1a=LXEB(>LOCCAAQgLfT/6,3BZ()&_C1[-4X[f@f7Of.>WSR\0&9<A
#-,UG).TgX@.^ITT6S_?M>d>8[-^X(bb0Z)+4>/AV5Tf2g34Q[Z+3\Y1]\0NO2Q:
?::F;(;DN-Y36&+R[ZQG7e1_/(#DJg8gYbRG?N<Zb5.39W2ba62d9D\8c?I/72,0
M0GK0^\PTG_6Z5OER+TFO\#4dX6L(2eQ,M[(.c>4CJDNePYV&K=NT(VD6LX3;TKO
JG0K3O\?O2U3a=_E@LO3,9::U=.)UGaf4@\X7T8I&d[7bPQON485R62IWF@5e(9O
_1Ob=P/<9S,?D>@8[8#511dPaZ+</-EJG6>Zb.[N<W@P8f+=L3800]EXc&O&S.Q]
bAO((bG#B1;I<#Wd1C>O3T4BZ6?+;VLS)S,9J=VP&;(JC6^>/-dL2=#Tbg-Q+#.:
=?+aLPO8)2;dK45(5+JL#2(D5Z4?1I+@ZC.NGW50\#O(DR[NB_U^_cUI>Ig5I=C>
=HY.)^XYe[B.9R7P:cVg4IX71FT2)GSJfSR(59OSWY:]=H(N-4EdP\/V1LS@bV3(
X2CcMg&;:4WT3PO);O/=/1ZMHOb]/?7_ZTDC(Zb#6EJ)YQU9IgZOd:ZS<6XQBLW/
80Pd1N=&S0P/;6a?I#fZ@;R?])6gg#BIF\2USQ_DU[bZC82;L0gR]PLPfUYUSCTH
02H4@RA^Y^_)W)SPDF6JDK?[_9=U/X?6V#MW<6VcBB.@/^>X3(/ed#NKDBV,H6BX
)HFGPI;XXI[/eFT>ge3Q0aJFW/U]/6RLC//7;XP4?fb0Ef8VOa^A:]1\]H-8Tg:L
R+JI<&2U4PeMf_7FASX</;K)?J_ZSWOd7fa[[HU_Y3BY/+6GZU7SV:4fR=[deZ_T
P@WS[[8dKeCPHb&F:C4.P2_Z44CEM7?V59]Jd.05ZQ4YHE+R34ILa_],H(3f,WBK
IQd@YNB0daJ=[9Vf4;I>fg0.]1,[cTMAW8RHOP4Qd\b-1A3N;-54e:aIJJK\)8S^
g3P<NOZ&aaI5IG)L](d2ZX?.G@6MgMb\9[X5<2=_QP0=7S(g33bR/P(H-SH)X<Z\
#g4UC,DNSg0(T=,I>Q.@ENWOd?I\8XU+^)1)ZU=-7D.=T>8O-.[/cM)-(-]/^97f
X7VDMHV7I1_)Za0VgQ\Rd;D+d)2(TG&#dN_IN3:R5b>,]>Xg>Tf(>-AC5>([A2Ya
E)TNZ;]L:Va)=O;bZY>V)7,eA4eV25@^+B3Nf8?YV5=;f&F(9bdAaM_fFN^cC4-e
V221U50EH2We1Y/agD#:,O=d0b?V8Y0bf47K9dOK\HAPDe):0281;QAR:<S]W([T
O<b/D:33<4C0dUV^&&.DF@=-K1#]d-;96,-O)6EgSR4J3C=S\bCCaU+C8CXY.#,c
1(=YCL[+g9a#_73d[M_I?F#JJ+)BSDRNeT4[>e9fZ41)\4f7<UgOPT:;T0W[d_#)
Qa2Ec:GcH)8[5BN55#Pe:FSE^TJZV:.6-=;C3IaB(#cfSVe]@TUCK]I@A5V:FIWN
gTKUFCSBa)_9]\Q:?caF5W]/:.2e:g7dP3A-(#/L>&M=2e.8&09T&d=eZQM@)U&Q
89FL&818Q)M=1#4,O\9fO2=fN,J\K4X[a[6,4(?H^^R;ZgGG_<;=F?:M]_RN1Y=Z
Y9;.Z-6AUDTH7f^HZgV0I5]9J#Q:aSc6-V<SH)K_ZTf4bDNPQ0:(FaQ^2,@e3[^7
R0CD^>.7E,8Pf08<//2SF)7X,_9D6\MZ6?RXc=]c9[9bMEg1>?A&c)G2RN?C]^?O
6f2&]MO2-TgTM5W0)a=[V:HSJegNF&-cZaM4Kc+S#d+IZd3+;/#83/)&_/_.\7G\
3:X5Z-H,,IAB]G^0Z#Y8Z5=3E#GLA=7cf,1J#P85&Hf82CT?d,Y/LOW(57_C0aZ5
A3Ja_#0e7:9G+X;XfFJ=/_<:_R6:GKA&(AC>cK[fEUf\gP5e2O3a.I7NN#g=B?HQ
a)N=NI]OMc_d^S^WdKS^5.?+0=2^[]Y],F9)TfJZb1DG3A&^I]H1T5_[aH),5^_2
)W3F.A-SaO/.8]Ga7XcF[8]1/agM^OH/H5?PG3XOA1]@G:VNSOT7C+cH:[caQ9//
/HYXeA5;.FP<K0J<BM+I@_AVITUZI29;B4V-b-c#O5^cFAY\Y#PR=S@00NA\I9HQ
.\eQ28Rd4NKJfcT58X;O<@J?XHB\V45]5_]c^V>?4W6ZFeX09LbeI?.S]++EV;@U
S/(>EBHd5[BA<3gNVV+BW8H1bKDAM_;?>.7B\(gE7A+V(PfN?Be_4M9<5-@R.fO1
_)SD&dIL<2>R&LLW5Q0),/RPE77,DcK1\b>4BS@5(+/P375(EM,^(R0+41:#M6K=
CQ&9JF]_\^<(g,2X57/-US2b-_3IA5dH9JOHUW.T+5Y[8X.RGPH[d6:De[^OC[G-
/0N._ISG1)QOPRWECQRedFJ8I_5THBEf0L.+Y2aCH-?f@[TI)9F?b(YgLP)BJ<Ic
L[PJd(T=9SIBP8W7Q2<;-H-3X81SF=.]:XcbL,D:_aTGf[[@]_>+A@U/:)1eb?BZ
YQGZ,VeZ^Ef_C8@T2dd;/JY&J7RTV-=Ve4N.fSP)<E7>S[^6N9K#^:(F@<A[L2#5
J3@TMPH-EWTWK>=IEVF6ZGRf]-B:4Y.0CP]ODNY5@UP)K[+K+K+bN_DI\-Q0=1E_
R89.g11C[^=5Z->D[;aebeM]+P5>V@RcDB?->g5(PJ-H^PYZCMQ1>))_.:]GRb:F
-PX,:Z87<cLO4?g)-SAJ=R-+Qb(/Q2)/BT2_Nf<EO:C-d5;g?RdL9G[N;.:G&aG5
Fac,_,MJ?R88]@J-(&^C/VBf-g;RN?P#WK5[G[R/eb&^]-(2cb63eRgMU\(JR2XC
L.Z0d@I9N^f-:8M_;?I3)J7[R9;BNAZAVbM?WgY8.U-B-BBQ[[@4C=EPB1OHb9g4
E<ER8R(e;[@QPP#?e1[dc6d+7^41DN,DI#@@.3#^fCS,(01@Xc:,<@#b6GXZ^S.M
eW5O>BFU]96)HO;#11dT>5Y0B-D=Z6,_D]T14RT8bb=HEC]LGXKc0aR/];8^J1ab
Y]HCT=dQ\\D/)a,-]/?.\OTY_CL61eM>9c?0L:d6B?FNNSQZ&.4#S?gRLUcae#C&
GH:9-;5N;VacO?;9RO3Ec:5A1##_#)ed#51;^5+<XUf3,LL6R:4.ET;O(8QcMD>D
Y?Uc[5#O50@[XNT\YR<PPXGX/HAd0?;C824GRX+@L7BPDa-gA73)I?7N#\GaGH,,
#U.Ga)26>>2\D\4YC1O(O^-L.U2.J_fA1HD[HAF->MTJXfXBE@L:E]TSXS+OGc8D
[DL/[3D(BZ0BBJC95F3e,X^KMS#8@9bM):55VDE;(CM:-)D8DRA#U;JDZX.-<^EO
K-J1,J[2>,feVKAR#Y0YIE]1OJ]-OF1+UbPBERQ]8d:&4]g[dEK)&IL@T9^b:eJ>
fe92Z?],9E9N,7B&[G<_gb]@I\8?7UDHLK6f+ge+CRJMf6D>HL[V.S_,A3,B(d2_
F6((4GYSa3geIEKFA5c)aH_6E)3/2CXa4YKAe9QJ3f.FIfPYb)4[DK+_g\<X6SY9
#9WV6I9Z7AA#D5_;Y5AOV^U3/C4Odba3>a&(H2W9U,K:Abb5>O)-,fF+4+._921O
W3=+X.D)_VG#_15X]:R8aEH#F]A^T7LXS^[^&G[cd2GDO#cTA<a6BFV<&c20#MDZ
+HfRIcC,./@#WQ<[:YGM4CTXW@ef:9^;\ZNQDdP=\[5=Z0/OU6/>48(U:.WPK7&D
)\Z=DT2L-6c1L]BY^[ceNbIb-[Be#CC4\d#?TRR+=ZRe@J+1;Y=R,QO/IL]M.L^O
JA68LV^;>)5bH8GZ#g]RZB2b?N?WJ1[DZQ#@d-Qa>(,#=E=KX<O,TJ(cZ-R&+S?&
:B41;_Od_EPW\71GgU4(ML&eBLD)HWF/99Z)-AE<:.Q[1:@6^R:.HdeHH2&(D[PX
E-N&E+;f9GR/4]<VLF^NH+_P0L@O@NL]S[;T65g#ZfRCU\ZI#P/.AaWf2R(L)EK[
.PNP9a1R>9T_OKE<Q#;Ea6D_E6e8T>e_;(Ycga-M[>G]@RL#3MP17<9F-^CDC0H\
N]V_I=>&d#,6&<fL@^4;ReN2a7SMGK&U-IIP&:K[/+2eFR4KW7_PIBb3RW-+CUFA
_bF5=#QW;]Pb:Q_\13f4LRJQI_\QA_SL7aJF82[CT7MJc)geVfB\fC:P\^We(QTK
3CcAD--GE?CXZW/@9MNK827[HBgC&J=;O#-[K[9>fdCXA^L60Y1XWF9e9BQ.<eS0
f1/3A[4)L@P@U3fffTMT\CHXJJ#YdL6BgF25RING/]#@HZSLN=)T+;D-/[AcHNgR
K:-MIZYeG-5e\g3O-ad6S-\C^.E/,RCPR34X@GHUY&&9XYE)B7-GX:Da(J#gSC[^
g[Y1La^8aZ(WIgV[?7bN1R^:OD;4AUST4X]Y4_/1d^QePgQD..H)f;WQ>[JD&C4U
bPOeVLe=XO.&\VVZBbb\N\1NO^6fc9Ta<T)M1Y20Y+#[\L,9;)00T9/b:/AK1_e-
U/<_W_A6_8Z9U<3?3UW5)5HDW?/-+c#\HN2F26=W?M8AZ:23\H<C>]IPUT3&)EJZ
BH;3OC-#-]THX6gF,&>G.Q(]4?:Z2eCcb#0fZX;O:1I9<(\P23^ESbRJcPNaP8?X
-:4V^T)84LW<10e#3=WIR.<.6:a]2]A#ede3I8^,,B6E#07Me1E;>UY].\g@dDb1
TD62MadF#/;QK0@#b#9LKf?F]L8=_B)DI^C#\?GT,fGg]1[Ic15.[e)fACS6TPD8
=P]]c;:Q5XL_gM5G0V_X4:@S5ICb<3D+eQ=1Z8K:I-RHOC.H3U[7[C95-A#F=I?<
QX>Z3ONXW&31c6OJ;-5<AH8dcEGDdK<GbA;;F=+G5,NI0VWgG^ED6<].V?5K6f]Z
]3_,J7VK.R>M62@<UE.ZAN_IGYXIWAL[8A)W^Q2BQR;WYV3\E@d(.1J1-\+^MQ[>
a5PUH?V:]ee^)?P-H/8d5/F,0cIRV.@174?X[_Nd86dc\JPa)/df7Q/_c&J]?da7
TNeI=F^PDF0L2[OB=S.a>Wf7/aUBBef\0OXaf4(LH5/+_&#Qb,ge<f>1P2&Ie=4]
NX^P;M4>#\f/ee0WMK@8QE-+0aGXZ?2&#aJ;8;Tg0:&.bDP#8F_Z(/Eg)RK/-7K9
5BQXW^e>B:8.02&QIM.5Fb(4:Ofc_4QDF)WY)S5:NO9E<7:-bfTG&gA5<aA#e+?I
L@Pe_OYI=TfLM2ZHZF7)1BMg+Z-[K[fMZH2NW/](?LMBEF-M@F-T6M3==5F5TcPg
_V5(LDG20OQ(?W-U8g[F-D9WGgR9?4SOY&HW+^f>?6C>&[#Z_&b(:U]).KBWfO9f
ODP2:a/Z;<a0S&>1TQN^g0fIX9@G-b0?D(HW3FN#=LM3bfe^c>R(@&K/;E3J48&S
&<3MN(d@5gc7)>6,f:?f2RQ5PN:,_+EQ(HDZ_TD/@]9T0(R?Te?B+>dBQ&2&X_EI
eBPZ.;4R.^6E(=a;[]:/+c8Oc6)QO^[?a+8>(.aNAbDJF,A^UO-K0ZJ,NQ9_8^H.
^HEV/fe/OG/TW(0X.WbF,EEZ8N+PWdS]GV8J=0g=?6Af/AX&2I?QXVB\gW,<LRD#
E(9#CC8NVPYf0,Y)&e8[T@W9.^-_@f#7;UTbFP(YUR+;],U9/HO.&?a>[9d1Q-&c
)dNFRH_R/&+NF439fc21c<dNH2E.Y<D.b^3[4?;cYE>QgfeVQ=L.QKd:dCef^6=N
[7XdS9[,4+=^U?,f9a:eF?E1YVZDb5_,)\+X1ZNUAK,NHR>?P/XZFD=ZX[R9fN17
SYb3cS?cARDR>4/HM<J&W1-LPO>?V.YfY>(bX@::,_@EfI<]#g=1H&GRc[/fIO1C
\\X7O]VZ?9RdV-d3)a.&O.)7McFTf&UHW_4E\0JYf]eY\8LdN^>VNS2aegH_UQ_1
01gG-WC>11TRCgYFTDO\CbX[7=^Q^?GcE&,,+^SNX)#TTf=DV5._=I-6>9JUAc[9
^d.2cb4V=LSRROHP/3,_6S,F(dG?F@3\Z#K(:3<7>X0)W9S5WERLA+I0:PZ4Z<Qf
0d@8)cD>9/a]240YgTbIQG#B1LGaN3\SJXU5c4e^3;OPd[E#T[.CK#7)EL9Ra?8#
IWf_L)N3XE:^QQYDV&JSJ:g4JH6^>&dKXR>.OI@+EN@B?.1)-<dR=f;)9NdMcI^>
_RO41-,7:7CUdFEU@(cg[K)CS?5WM>a@,0KG[2.J\N8gHA\b5T\]f?K,LZ,Tb+XL
G+:V4PQ;.;;e1V(.V:^LX>DD-<E-dGW;F-)EbCWQ)BL&=WP5(9_D3?+D\gV)@AHb
d.X4GU)Sg7P0_@SeF-:dRfAM_e2,S2)GQH8bY(IYc&f#0Q/_.DWNXU\d&5_@<CBL
DK(H>A7[=V^G\_g1,;f,U@8e2:d?3YdJWC#2_-]+[cX;9aNE)DN<94(&O@W-?C#+
[53\OL]RJV2PcO@96L#H&94NO@];#5\6X2\]\Z^][9A/ReA<]JUC(FQ@(-8J[X\K
P99VA64XR^2U7)YT=(f.c],\#WaU[HO#:;1b1CK(&2BMbP:^YSH(eLSYUPNQ)8\4
K>b>J0,FJDR8066[PZG/26??(e4>b5W?B:>-UHaV]^W=Y0@ZgR6+Qb0N?2)2bWU5
^31f(^Z-TE9R<SGSPPc:6eG2dagBD<>f&M?3D@BMSAV^e19V]QCLON_1\Q:e078;
?7[4fR&5dTOVT#7W+BKAL>NTGaVfXQW1e_F;3R)HSR;,BS#cDB-V<8,(8d&^JIB]
&?&e)\Sg-951HaCH\(b:/O^bT<J\B)50ddN8>=WFZBR5G7W>eFG4GDf+BQ2bab^>
MbfJNN(W[MeG]J6X7,MF]?O(]EO[=H/a#=X7^OURYD3WX0[UX02e0]2?\=8+1Y^P
;YM26(UL(5^O+Z0eAH)PDD[F]9A5@1-#F>BgWGXe[?86F:,<8WFY-YQM^IW<A_W3
gC-,TPGO.c-&._O-6X450bE;4a\X(<VefY3M.&,\9W8P4T6d@7dCRU-:]PKaUZ+A
:d/d/SadaYJZR2&b&fQd[ITJAFVZ;BE^E7e<[f:(E,SVP\MGZZ,[5,TO;1]ILBcM
W?4R-bTUEY^=_#5O(G^(gfZST?,-(F4BbP^=8CRI7TSSFc=(VC\(X^],D1:^KS9J
3LC:E/7gf#aKJ^XfX.O,g&&,KE7O5-IDUbcIE9>Q.WMAS[Q>\LUfXLa?MIG1E=g>
Y(MRI:Q;\]WYW9800UX<:FS0[YT]c?H5YFN+[-XgDT=TYdX?,&6YH_,6TD>(.C;T
D92S/7ZQU:dK7KQfQK-V@I/]4A.N5[>-Sb^&Dd@/R[JQC;@-Y2fX8PM\+<f^(_@#
0,+gOP.5T?;.T7)L.M2H\BEI=7S8W@;?M9edc3#&g)>[NU>.;^H;7(LTKC<g8AL\
3)ebEF8_E9eJ-e9BT>_>Q-RV@WJE.AA+5^7T06)60B]SEJ7;BE2T#F](]5#9/L85
V_E44e3::,VX-AP8N65=BTGc,/6X,a)RH5Z0JP]+/f&PVd&-4?M9_XO8N<U,WW\Q
)aeG)TY[)gFVURVEb?&AdH(7R+3N6/]CX>A<d_HSU)bdHAbUV/c<6UJagIO7&]+4
9W?d]99:\K5_cb#K@,O9E:HPMY1f2F+d3/O^5E,,2EaCYb/PN)I+WgC4<gd3Y.?g
64W0Wf2dGO_ZS[gOcU.PUIC0D:A)E[eQRfZ9I:,d6MFO&8M:_JR?\SJ(#=e4&K2,
QNRCY-0Y\Y:^R>[3Kg>I&Aeb0ZPb_5,I0XK0WC)&]KUXSY=@CZgAf[a0M_7CeYLJ
:K-:[GEfC4#<g-a)&\]G8:aSLJVK3LNbfUV1;/]<>-<eeOTGa_SaCY,7E23R_9:+
Td^dX1b<2WT8,OY\b2\N^bf3_fa^1eUQ3HVS.(,DEWSZ_/K3bW-@>V^a9O)&O^#]
[P[6H>\;DO]=,LXQM+VWPbCPRGLgXeLEE;HZ999#0:2_4gbTe[C_gI5T[TL<6;BB
M-c=B6XL?1195RYUG&>/GIX[;IZLG9-&#RI:@g7[a-WM<@5CW)/=EHe]R,HMXD6;
RYd2?6<=:^a>;L8]_??<AWTgg3/8fRGcH-;TM[@cL3YOQgT#)/]\DK/=?5\3HcY[
&2e7]10LV#X\6E/^]AN;Y1EWY_gFf^,(aHN(Q(]F704(M1JIH<6?;E7IcRYF1fZN
DaYLT-=gSU2KM7IPKW:a;)[/(E.:F18O#:Q6RN>DbUeIL8GR)7@-VAHS15U>DPgP
-fK;9G;XOVWWCbc0/WTU5gG;I#9/[((gW=_R1BQeNR.ZNZM426-c?3EBE61<BU._
6Z.ObcC3X//F;;QE0dd:39&KFPIM9IF(cUfI+caO&GZ7T=a#),IdI74Mbc:B&JK]
:V44/9,\IId(K#Q+eW6[2#-UBSaF^-;;>0&0ab>H6JW2@(.&-+[6D[YKe1?eNOGS
^;CBRXT7N\c;EZ_16JZ@XaU:T3aAY[NN443FJ7#Z0?UP\4\NG/JI2Q6cU5C-XB[\
AA.:GV<(P5<cB6U1:Ve@FY6RKW=gB#NbT.O+A7]c2487FNN.CVL3P2Sb9EQ?:REI
,@A(^.@-;LC)A.e-8J]Y_W.NW^c.PAMBA#L46_aQPXS9Qe_O:ad:8FTIU:2Vg,DD
3<LN++VY==+RBDfQeT#-Z[83gR<b8eAW@E.VdKI4gb&8>Ae0:aGA76?+[N;/DL1a
C-C]2X@+0D[=#>4f6I80bTQ]FWL=,_MUNHgN@<Aa\\HdDOG\IB;KG]PdKKZ:7LD#
81/4_(g1:50Y-ZY+D[+ND-JgCJQ7K>:Y;2,X2Ve7&L2Ya#,AZ,>4d2Y<BP)<+\56
=gJ0]b^W-QG<2>&dI/aEXedE>44^6R_+aD.)IdBC(.a:5V4>7>KCVK.AcP5+3L53
WZ5<#Q77eI2\gY>W23I(,M&A1)+a3Q0?=)Bb?N;5TA_e1@2B8?f/082#-Y3,QUbI
4];JDCC#b(e?Fd.9g<BaH?SZ(4BKMZ?LP/5EVWMg8cZ1<K:d6UFH\_3]X4^V6(Rg
Pa2P5:UPZ(O<LS<]RW4cMR:-0AZ.=KUK7/gATU3][g[(Zb5T]Gg\;9.P00NG=XT=
<<SPC3^;GI@NVDMeQc9B64GdD75/2&6+<?=(UTV1/FRO]6MX^P#V.Z9-/GR6;eKW
X&-.G07X0(YK6QX8;-3^,B:8XY<4P770Ua&BeDeJ,06ge,>P1R</JU^[R(=[]OEf
::Q&:RB_._CJGFZ:JgT]]J2[[=)fLS6=_1Z,ZLJK:f5Q[dEb@:9A_EP9@dA,&2CE
YX>,3?WWEY)]PJ#X2_(L#7:Igd#+QG<cT;X-_7[-0]4,:7.I&Veb>7eSK_J+@QZ.
MTCb(gg\IN3T9UOScM>[0^Y^:(BMF=gK94&QAb22\CHS63J+LM)E@K^D#CDXX&I+
JQ[34MN3L;f37(G[Z=D9\9I[UBUY?OL?LO+A<Y.0_J1YKRc..H^=QIFM[e?=N1;O
=@B[_Z?,cY=7d-Xf?aOVQT=(R3/=+6VcgA[N](MLIP,+fdA7LDZ1B@TISb/0W>]<
dEZG+O2J<]O>)1LKaDRA?1f.JBIC#90?22Rc+g0=1H5EMG(dZB]?LL5],,AIDFVY
)UeMVRdK::X3TM36?KI;^9KL>4d?(aOT+ALX&5e?-EUfeaB:OdU0T+QVJE=eEb^5
:5UUD=cNZWCW2SIQ3(HGG7IG,&X7Tf3Q.H&VVD/EdEZV<]7bXYD^<QP;926;F+19
:]_U3(1OW=/eCX;>;3g-OR4-/@CU^4[?Pf&GF3T+TUI#L@XNMV]8U2K9WaN80W\7
?IY@a#PI/]B/TFb5=R37=cf^f8&gUb_Z?;42,=5;eIA;L.-e\^eDePD[W)9XQFR\
CTL^P1fIGYPW(H+RLbI#;#;N>FGf<1L#-+XK_ATH2HO3,1E;=g270>-8(K32W/\e
D;YFD^<PM-L6c/A.8Y]EX@L:1]QT:<\()1ESNQ;T.0(^./E.MB&T?&XY(3Q@PF-T
bU_]/8P]?^6aHOHZ91L.8;SV8DOV56._O#e+6#H?e.04g@3]g:\:9;JP@#bLF-FY
fNT3RIP(/YK_(M0GF&9L:-WB_VN;^(,H3JZUWJW233B.eA_Z-7K=6OCY3A+>KLY-
Y5G#27b:9ABcA3_0Y8;M0NG-.LbXBKE[A2F7c+\F6O6Z/ccZ)dK8-1/L)M0H@#6<
Ig6c5;4a5d+9gC18)EDMY2a)c;b#S.UT5Q[6^Y1TR=8^I=gEa?&B4V=SK9AE1Z+?
bg&\5&Jc[bB=_ZGJY&3U)<EII6^HCX^&1Y5+P7Ce7D_[S70a.0[V0bbQ2G6Z]T#=
#V9M]c+FEPX\H_0=UVgb4YZ3bH2K&,3)UQF=OG?]_d9DCZG0MAMfYV&D&=.FI.CW
fHZYePOQ0HHBg+?Q5V2;6H57C#I9TV2C-2)RM@M94SRc07Y?F/T@I]KDcINSDK-(
]a=\XNF6<7a:XO^5dK6c]CZ(gZ?F6M5.6ZOXF\+</X4dR=ECSN;)SbB=3X(f]FJ]
T,^T@O9/B2A_A.=eQbQ02TaGUG)>8TKV/9<fM:B(?)X;V5G6W(W).FB.N.BTJ-YT
C4J]1NHGVR+KWW6f[.PO@09#Ta0Z^HA3?;&6bJ^?#(7TD_Mga4XQ1SdfS)TdZ+HC
X&W?=>99dY:bB#SMe[(W2,;=2C&gJ6(0Y7MRQ@/SAe?1V3P1VFd7XS&b.aQV9SND
c(9IL+PH?aT#?ad[.:DR((@+H\]G1bXbH^6_YOg/9_H.>fQHE25A\FcHI&)>7cac
4)KAMSaVcU)C-&(W.]+X;e,Q]6W+d0>-=-?2WI,/KSLD9bW8@Q6S#c?F^Mf^6_5.
[e&(A1.d>b+NU94g7-&-=YCXe)1S_a>[1_/>H;8>>dU;PTYT[W);G2_2?H7S>+=1
.-U\5_g5W8,9^+\PZWNONg+c8Y81;=gF;RJ_-S./9IR-L:H[^FBDVB;Yc1HG=0#.
-E:.GF-g;J+:+cM<gN9ge3PG/)Bg#^QA-Y47>XF?OJA+GQN?PZ>8R\JaHBH@^G6/
,F+[Oe]TD]Yd77PG7fgX3+1B8=Pd<6DVV\V3\9HK2UJ/XZ()S<b>g:&[04M<gMbO
#7gaO]Y\07-aU8N-I\W;P+RG-8bNR7GAD;R1YH5;PJY]b#K/94F:Bg/(7g+&a.6Q
H_TY&<?TBA;/Y^EXe3/5+CV)OB@)AGNX<e4S9RPeNSbM=&f=H-.N+K]^U-#2H8WT
cX5bAV&8^98U(JGbSW;3Ja\g.#,QV<QA?&C=+9bXX#HJB371(4TJ\KKb,:H6O@9D
2??:?9Z_8[,H<3K^(dQH/W2@JX,d(P;MCXGd=&7LU/Z#_Hc_Q\YD9e8J;^(RR=9c
^KM9LCfE8N.B>E\-357DS(HZ^N=]_FG-9+7O2DI=.@>4Oce5L7^V=W2OP4UWX.;B
Hf]U1M@#DRAPCK/<:NA4NP@ReF7(A.PS-a;6FLGO@MGPeI32?A;T(13\WL6O1f^_
#)3)A7-UZGDOJLT47WY:C1bE#;D[6_#:d12N+-U6B/0dCW.S](0BEWc2LHAA;9X\
e?fPePECAVP)B,cOVFU^49#Kf[<&Zf:f,5YE?-/DRXZ;HHX^O.[cdU2c57+^be18
-J(W<fM]b8^\E@C12>g^OCLG777#>g1M[4HQ05U8;H&=dW=9DO91E51&I3,101aO
P]^#cFJ#/BA^f-QA>X_dCC>eFAIba-HY5IU5FQV;g^7L35=T1+e^+9[=f7=EE@f(
UUAT#45\]>3(cW:R8I-Ee5RQ-3fP7XYN[dZB,0G751>YKYR=QH)@J2;=fP<R0JbT
P9[?:2@PHJf2L(d16?YFVDf#_.c=MA\2fP9LdHC3-#bQ]32d][[HRa#\P=Y9&^dY
],JbCg7fffV]:H=a>;_^eb5c;FcKK?BDJ.B&a&RQ10(ZG)68B,WQJgd4)<Vc\Z.5
^2RTMbEP+B]Z=&;(.)9TLN\d/JU5@HN2MFF<GKD8FT0^5+3g&1BYG;1,6\H[)+6\
U7LfcI.=&b\QPJ@16L/K6_FBSeNLd@>495=EfT=6M2?K-@.;W96fM_Pc9^(;S:cY
d6W<C2O<>,,9<Z/>>KEg,O(eRBM4I#NYPM+5eZ4KJC-VE+D6F[\/LF#1DNg4Zbg9
?f,/SV/-L207;S9^7.cLKDE8H<HHdJcTab#^8+PU^+WDGY/[I3_f0UE[^JA&A.)]
4+-<aIVQ>bfe:QS&HC<NKE0&>R1=#&8gJ_1[,&^_W[6F^\]X7\94X=].Ig^6ZQR9
g+I20b@QB0W/-C5_]c-Ib04PCK<[eN/3,T8GD8HCA:/f90YR\_N?#MeQ64/<_g1^
MNT0;HdH9MZ/D?RV:B;[45-+5H6aDUY2Y###J251??Ic=:=6^CDeG984aF/W:6K6
+Q/(L,+PX>Ua60fLVP08_TR-AV/BVC\:QR1QSBXRf+&a(@^:eOd3&O^->ZWOPT4Q
9@52Tgdf\b7&3+#739Q.W7A>MEf52dK37?T1DXGG0aS)\.UJYSW,CA[\<;BJ:eAI
HQ@db5]f>6E#]DZdOMITHHQ5LXE^[f7;OZ<.R<XX##M]H.^V^3M?gJ,)FCf7]Q(6
D\HXW[a0R^8<g1a5)=WX,[(9eaFE_cCF@D.<5J+e:^W5Fc>bg0ZDV(H[#\8.YBV.
QA^dJUfTE->5C\XgN[^9V[Q<U;RfRGBIK(&efI0cMQ2FKI@-.A[(DDLG&ZF4FSBN
#FM)QW4,&-PQ?>XE&?>WgQ\)eIb6)(Z]4I>/+@+PJP=0]b\\7cSR-HAE7FK\8D0E
GbLW:S28Q.5K;_CHY5Q\CRdJ@KHB&/KH#>Ef4;=^e:[?ZQc;NZ^:\QaIK62M+4I,
BBA/5LE[,V8=#3\6b)fQ=MZOCW[.TcBMPLP2a15Z#D;KbIZ&Ud&_I#gbc&^e@)S4
7R.cLbD?I?W\2W(>#_0]OYe/6]d6cd@HdE/Q3Z49g\Re@,#5,3^;;N?G#1S_.cFC
KDS(5PY:RS2[IHS.P.SYG@I/5>O1-3F^bc7>9_ca5?13_:EC@>T#QX+McS+.?@&0
[YBV<(.)Y^BS1P7YM>(+V8BB5VCMb,4Od=#USNBT?CC#,6I2;J-^WJ@bRE6UbI9^
J@(9#79bcAH#f/L_0S_7FKSA9++E_)J6GgVEAU?fP7HY&ET+)DD:dZ)5J/bL1WK0
>7RSEN4JZf-)a\L4baZc3;M??P4S12^CAB1GP;F2bMb@aFE.Y>I=3f=9a0)+F-;P
W6b1DUeD=5K0XebGDJI)eLZ7E&_/AcL2EgG2VT,AVe/>CJ&-#Z+WX=HEV#O1\&8>
C1WQ7V8MB^VFVgAU2#+eBSM/FNW&=?gf_4RZBK=B(XgS.-Xf&SH?&O:I()0:9RZb
[JA=JO6<0FB0<;(?F65E&RZ4MCDO4?1>,gAW14b3I#]V)\+fFQ,:D3[Pb6A#4.LI
,fGMC6HL?GQ#3@I>.8]I::V=N29^\bR3L1aD?\7TEXC]GG2&9(LcM0\&G;VLO+@7
NO[5ae5NbR/A:RZ^PFZM2;U?^CE>@U?.:OI(B,0]3;<<fC9JK(1ffZ5U=TC^7aQ4
R@#RLDJON>QM)P7/f@Z1P#WZNeWP\&+0,Me?+[PMA.EMGXJFf4UX68J[BTc\Z#<Y
e&[Q5TI&bEAL8B<I6(g2W_3\C\[Pd7B72XL;4?U0QFa=>Y8+Sd/EM54]MW7@5e7&
141FKe;Q&85#6^EB4-gA#-cFZTM_/ZCY353QBF=X1a1g4Q6dcCAKd5W9a6I-(US8
2P[c+;a=gY^PV_JWR=Z4YKIMFNFC4d0P6TQ]@NDJ>WaCFc_F[NKC&0g,<#.4J;Q1
>.I]]01;VaA.8FDVO?3dU)PUIb_;Z,d5>J3bd\S?;Cd,T#\>G3X)TLPb\:)g<UEE
ATeNJWXC;,22B9:)C8T6gX<g6d82E:>4(aT6KadAFXLI.C[WU]bK/K0LI=<?.\fL
d@0E3cG(04Gb+f8G(91f3+aG+cc>VO0^2H_N+bfIa(XG+>2PI[#JG2NcZHK24.,3
2]QH1#JO/bGN<gbg4P#CZY>DKBWUB<\eL]K,HKaTN(GBO9C:_X9Q96@HRf<TA\fG
,N#Jg;0KU1KV4MdDP4VRg0N.L.J7WaZT)IC&@60KBLPgVd)&)9gE2=<HMWA1+>bI
:62M/.Ld8\:^,TGCD-N[OPH_R)1^?aLXH+6e+(.CbH4BNU5,Pbeg=P^>-(9A?=(Y
4N],9(1M[)Ze\2+D;6c7?17Y_Y,_\,;+8f?U/^GG@5V]_OR/V3H;JKe_B.?MP]0D
=O=/&Mf]5&1F&c+2Jfd:#[RY7KVS4ab?G(b?/^FUV?PIQ-Z^_FaHOg,I:c6[S^7Y
5WIL)EXQ-,3NH/SG5M#:>:2/_N67,<HZdUR+-MB,I2g0RcVLLQPg68M+XY.Y?MB^
NH&0MQ./#dIN8P1YV;[Ea2P:.+0SOLN(IQg=&PWJaT?0E<2,F@#X6-<A#SGAgK/P
NdX[_c#D&2V&)UF>\R&,X<(PP<b4d(O22JV=NQS>9[.[JAG4Ng&R^9QR4dG2/?DU
-)L65;F_3-af0@C1RgO<>W#Zd4Y\?_ZVDAEb6VZ02Z>^-dD5PTV><H(BL^c_-K=K
X6\HGTNB3E0.BI[6CHN3-R51OP;GYR82(B.ZYaCXDQ^QGDRUPWGV-LLG2)?PeFHH
Q[P57Q@4E&?@9G[HWD52:AIZeeJMI>Z--f<S(8+D5cOAIJ;B?6+K(0^fE8@b?5ES
cAVNfS_@cYYAIPb4fCU?CR-K@K:8Bgb+2@\gXWbFC&(_;0b<8@8WGP@JBG.P:I]-
:S]5dUOBKf9Fg73/4=IK9Q\;\#T+;:Sg6^DPP6+L#9XNUHM@\N/eV;RdV;6Y-L_Q
fB>CRF510^?+RE]?a-HY>U4H9df.B?>F.bL0>,,[Bb:E-EXY[/YcI66W\7Ra.E4\
TH^]CNCWT6^K,1L\<(;PVV7XJ:Q7D9^>\6>O9KSFF&;,Z3+FEg<K^S&W??YJe-MP
=B<6YV&9>21E5GYC\A@2-=Mc3c@NN@C5AP7Z\2PJB]B9E-4b(6W]>OK3[\UPQ;9:
@_@d=L7Abe>4:&+#GUQ7#UM)Wd-CCE;aJ[SN&Odf]eV,g>C42fJ&.M/R/^]7Z_Oc
)?/Y5;OD5^Q-<B+2KT=29H-/+:_T(T#VG5K->)LA4U1_7aS?Z/.TG^ccTUZV]3EQ
/d3HYW^T=HY0>]a1U&B5B-^882Z=;MX,P/=_d/PS-U#1N\2CWT<af?J[aM>ecZP_
b=FI?OP]B4YW)e[&R2?;\>(EY^(Y:R^@#H=[;62QW,I001JD,S:_UNFfJ7Cc2CL,
H<Q3JZ;_.eE]6J-OG)PZ3_M-.6QB/8F/+5\PZFbG)A__SaC568Zfe:=5(JS#3&45
J6?UX&FT3Qc.WYTG^HL33).]-2:JTGER5E1M>Xa]1?2c2@b#7^-Ie>DQA+,B4@U-
H^W6-dDGUGFIUJ]R=NbNgWSf+9Q9?(K4,C4+bcUV[fVZE<efE4.UY),J6)KQ3FY_
#]a=/@M+4f<G-E>>cSP)TaP)Q3PGLRXJ=DW=f7)7ad[UPA68>FTN.(DTT(Hfb(8>
914EO:.QO@[[(2Lf:M[JZVCJ9,(-e77Tcg<5=bK=LV@LW8Z.C/E.P.(DY#BU6SFJ
BHD4YQO03DX[KB9R=>#bX:OaAcG_#2>b\LD;E.@V8IU6AFL9deIC.YJ6Gf30^<UO
8Daa21&UO2[]M\;(=ZT6ggD+WCLXRbXbCa(84;ad_[,8U\K,@c\=BeHZaf]\1C)>
5@IDMdT:a3I^>Z20L5A1RI7TFG3c?>N-,2>G+e#@=aVFLWc:@QP0a4=Qc.YJ#8/e
GE#N:\XCNc/<6/K<6U5:KSR&YC,2d_;bFS&:RM64Q_Z-BA>_LZ#-=6W_WB0DVQ2M
;g4YHg:P#e6TQ7_c?NN/LU>-K9FdX010fQ)L\7XQH#1Xf[>8d[e2Y/7-1O=6<=K=
;N]CIN97:^c-L>JZJ<)_S^MI<G&O9f>V:6/F+8)=c\N0TZ:AVW>>.)a(MG\8SffK
[W@]8(TNP:?:dY^:V)OeMZa=G#O.:_6AJ2PBEK^NN:-FM3ZSC=A7/FL0E3\C<(5&
\X@.(JKVb(f/UHGQ:L,bJ&^8V(/H0\M?gMAcYJTTZ)=B01C-;)[@0WG=G<X.?;>H
4^.;VY[_4bM./,QQ-BWKeJR/,739BS;f]d([bHK\ZcDDD/fO>/^fb\J?f;LI5d2_
H/L?a>S>=_GPMSQ;<]e2bNVd86VfGdZKELd+^b_:a?K_SYMQMaaV;V[UFccK_4b)
&#4?76DSGa=VbC@U<XQZc3NA]LR]Rb@)\GX=VQe_-6]eW8^V?M36.P6EOgP?W[MI
UEceKO1^P4JEAN@XS<@Gc6W#=GG#Z#;IHAb)F&9Z)K_5C1YG[+AK-N0WbgD[bD</
:J<^BDS6N:gEV_I@JXP/A0EPOdB/OG4,U1:045O^a-=,BER:^3?/FB=OXO_,D94+
]A@GM-^A4IQG[Ic26#KJKg?0/[VN5&[2ZTJ)WG<B@8)RBfS_HFS1e+MdB-6(C.S6
;F1:KbGb:#091Ye<Od,aV)WN0VW#bWE/K6NYE5e9=<\9M=<f;g=cXK#e3J+U\Lg3
]3\2fYD9B].#Z.49K/?3,RTG8cdP0H)EQf_<b8WL0P)g>3PU_5,YHURNJ]0F@8(N
bf8R5+VDT]<gW3Hb[/V#TUR0T9BZ?EXaA9R)0Za#SJ3:(G\DM(7\DgE-Y4YgaSJ8
8+3ZJT98)923Sa6)(\-C^JFD&B^)RHFEP58EC]&eX[Y>4ATWWc/9f+L\B3#fW\S&
CHNF1f=3)._2Y<U-FL0/HR4;e^7-ebReB4I6;NK\=ORJVYEBA#T;SJ(@gIOWE7?>
S\MQ@J.&KOR(Rc&D<YEDf\&WSCDZ&C6_cDg-c.S7@T+[M_/1#d\(NB2UC:=,^^.J
L0WOFfg(a[A[L\W+YW7E@WP]fYU^a<TOE]T^OECEE=XO]Qf,@L.2PM1,efWFL8>I
RBaX+P0I;2S?c+\13S^/a[MMST@T6-(/ER5ee7-E:aWO.F7;=/6;TT>VJ:e7O4L0
dc7\O?;G/FVZW^c+5N?Ic2VZ(7]\.6gJ6b1C3aC/5cd&.f\C[RY]GCMg#]>P-->T
LQfC&:DV;FK&F/X0(:\2>S\)L??SgA15BQ646a/S=;O8B:R9QX=R=G(9aJ/;HJSZ
FdY5bP=7#a?LPcLU,Y]d?3fY5&Y^MF:9?8;(>a[G6?+:SIVDEA&3K0K/dO-:W)e^
OL2&GETb#]D(3&d:O;3?Z[dAT@&&e<9/8L?J-1Y;LMZgRE7BM,+R,(FI>IEFA2=B
d1=g-7K&Sec@\#2<V-.8cK=I0DQaQA#@CN<=D)([Fag2:?1U,O4<V)b,_a^/#D3Z
RJU&e?.L8gH<=43[_R=T+OZe8WXL>ZS<#&KJ[.eOP.,:_>KNXR(WBf]O^_Z6bPZ?
abAJ+2^]Pc.5?QEeJD&:G1d1F/8?[6_b(;EdR0c;+LMd]&]\&=3_#gC<O@5Sfd2?
]+P0=FR<79[^(.QI[;eTHAagZ_HMBSB?8]d9:B6((V_CB6Y>283EJY6UQ+4:1&Ge
YQ&_d,CMKcB@>G263:PTd)N(-=<fVX8;9dIO-d<E:6fG+5.7/T;OFU.BF1dYK0dD
B_2076ON)?ZSZNge+FM5A4aBd6DLEcRDXD1:10LR8:d@6:+?[CDLS>99;F82>>,R
@ebc0LU(&G2eC32dfI5gKXZRf_YNAZ)8Z2Y,?M.352W(U;^OY,+(8W9[=^KKOG#9
2>RN.f5MdFQ\C_4R+7ZZOHOY-22adE&V6V@.1FYdI<e#,93J/5I1(Z8MB<3-9#51
c8O;YaKedMPFaNP#ABWe=N>6URY7W-8[#L9_WGcQ[L,@;-\Oc-9JP;R=(GDZ\_=?
F(Ld))633GI@;Gf+5IW05R#I^?;dG8J82/U1PKAZ?ce_d1eHMZV^>GHECQ6<e(,R
W<W_P5+/]R71#QP6CP=F19WQ@;DQXfb4VZ0Sc_#5.KRYH@]7@?:Q4>@,4LR_JM&X
R?APcLQ3I;;NP97YaWX1D?L,@Y2dQ5dJfHaB9L^c1SU4;UQ;Ed#)T>b>d?C^:+[6
I(X1&+C2\:RG/R33;6-21R2S1<Z88AgUX^]9^W^-W+CHS,=Nb/KaJZQ?6Q1I;26:
.@Ua<NX0T5==F9FS5=SH7dKWVe?cC]SDf>GM&ND@T1(VJRb+A+J:@?E&F=XF]1eE
Xg.^H:((gOgM#;QDcc_1E[68fSIN#L&1D<75AK9YUa^WOH&D&XGe5\T.V#OH5RO^
BdTBG:Q;5Ig+P?4Z?dO&bfFeZZf4=f52Ob20NDHMHH4&Z28<QCF?Jf.[&NIE+dE+
76E>@Q+UO>_8-D?9,RT_W8Z(0N80EK)S>.IHfBB]8)W<@EdMX3C:T:R=;JD]?f.8
D(X?TH[Ha;EE>SFKKA102>YQ5I^RX+R.7d^+)GFAM8gF/&Jd<&R?/PF<U#J(b[M9
K])9#F6V=-HQI5)JEZL&<MPKY1DE5ZJI,F)3;D3MbYXXN<&GX+T^egY=.SZ<@BA-
:_8O=97XSTS55XfOVSP.<PMOK/A-O/HOA-S6\KJX7N?##f_^W.NV0>;LS+\_:P(Y
aeZ+<^O1E10Q>2PA4CRE0?bIL>g@>BSeREe4d-eM/<@H57.gG=MN+[1[4I^C-_Ta
Y7&;)L54UEW9cP5Hg,a;CeL2R28;=0OW&E_EKEO=?(bFM:g2Y#dY^=0K4N=/e_IA
KP[?/BY1VdHHPRb2T+]M0#O,^EMQRK_#TL\UdJGIUJM^^SddG\aTKT1&,(dU>=6Q
YS,0:g8T?cCF.L6VE=>H>UFWP4F]2W&1T0@;-/L&<B?G^.?M8E:.L\b(G^EQSN.I
fIF\Z6<;/)\9cB:12P;09,&a#bW2+:4b_D^_e<<3XaS<P\[2,(4CEOD[AVRLY:/O
Ma3da?;/[C[)YD\\YM8dG0Y@22QIYRe+.Z,f71GE3=4ZE040[[4YG#=Wd[,JWFVW
-=V?0W0R(Y=1(c@-BCM/7P7Gf_N@3)L0>7WD0#QCI,7P.f<d:c-4OCMOU4WdZ?Nc
+GC)T>fF[WB1HG]E^)0Q3KW#Q6;7GeB=1+.77#eB-b)VN4Y,d99H8Z?fdA](MbGW
]S_9J.G_-=ZMOD\+<@bA#AU@36bSKFD9+?ETKNCCZdY=W^+:Z>?+gS+.:NNZg1(f
N4E45RI)7Qg&/1;/7W,;;_W9#E7@+eV>_CFAQ52PY,?da6<5Z8Uc.S^7\:+EfRP<
H\1XR]VZ>]G51/V]S/-.TbL3g&O2XacLC9S]RAd/>I+fH[JbT_3N2MXYa_KfAC>]
16@.U.M9/M7EOFAUfYSK;J\Ab+F]-.DUa0:-E7:P?EG^+G)379P34ZUgN#?OQ8A:
K<^e(:-Z@<.E7&&C_Q?<I/c30]0O0R181?[D/Bd.P+<@5d1OW=f/C?+0\=UE=)1,
FBd2TM4LcdQF[eQ:<0QCP-g_]WB=PV</?I&eJJ(<X>(Ba?U:;VHD\<P1M0X_DFb5
:Y4_</P4CUX,aO[2ZK[&fOI63[DE?2&Z#]6HDW4J))3J70U-):VG8D0eIEDR?0P]
\^b&^YJZ13LUCVY5ZJ4=;ce(9A+77@@.cQLaJ1]a9a0\VQPf-2>SRRJUVOVJOUJ1
)3_d-<P@I;U25]X][3>)7,c6C+KJ804g,T=5W2ZI_N]Q2:X;FH\K/7c5WF-=^Q:[
R3ZG[3-:C@XX][g4bFE1Y#ReL/aRH,#W\3+6X<12]=-Z0e3+aZ.GJGQBF;Z]GgeQ
K5;)C]E1.;eZ^1N;@R-f9]SE&IgS\_Xf_c(51M5:MaN5L&bEZCM+;9PEIfO(e@?b
/Y_,e2RQDK8/aX28>VL92f-N+__@::57\^0O8?/a.<7?[&<@.=WADNJ3<dN3]Q\b
YQ.VbFU2C76(OZ_S:V]AgO40DX,4\G+ZWO#&FW@RM&??JP+Z.C;4H.,JJ<+cAaYW
I]0A6ccc51?TVP\94aYYRE)>9(7R4]f+cEBL6A>7,KA02[@0JO9=g;,P8f48aG40
dg-c7UOf1]/ZXNg^N9G4TefPDg0MIZIeL)QX&:gL8gQB:A:c2B/TbF(,Jb=8XQ5.
^M+\AXSf+F)4>[CZ##PMaZ945N+M?_SQNbf_eB4Q\g=&Pb.R9H4#>188T@b/G=Tb
YWGeNaHOVJ8a2V>4Y#&&35WbI8GO+PeQZ)#[D9Fd(C84f)BP2,TPA8a3WVFUR5/8
)Cgf#[?=50N2Q+:=HD77C(e]4SOd=^U>G6R3/FZD<)JA?_DgSBF#2PTQaV3@=,<Y
?TO9\Qc2C=YDB5NH#J&G[:J9Ie0;SO.K>JMfNN_DN6KH7G3;f.9.Vf.)PG(.KU.-
3e3,XB:7V6&R/7LMR@DEW:9-[JI/8JESe75NQYHR)YF^TM+6Xc-UK)OKJW+W;USC
T@@THf<8I)0NA9KA;P@T2f\C4];X=>](Z(]e2I;0)-:6,e;[)C_<2Fc/ZeJK5Ue@
Yd-07T@N\&AEL8GSNX]U[(I.4T(3Q[?&;X_C;H#fCb1aZSefDaW14.50UGMIRYd#
K/[7@#DKcJPA#Ka#O_4NaNVLG2fgWT2afHM=PAIVM749\,1@VE94f2+g;&2-ZZ;U
38SGd^P1[^+b3ebdeM_OVI844.G?,9+F\8_VQ^,/Q;OOG,X6DP=DZOf(DG<V<Y,H
TU-GU4-@-N2#-/E1P6[LQY.[7+>9gR-/>_b3<Vb8:914)EDEF4-=1cIBEJ[RF_aG
GKRc.X3:I\^f:b5?HB4H4RF>MPE0,\V:L/&M,56LP3SJ41=K0=?e9G3F(?JSES_>
ge4dPA;GVgD<QOf#GHE:+Oc0G_Yf#-7XFUdP<)47bD3_;fTSHf+.0I>L-AY@(bM>
^gHefG^?GE/WMVf<YD);0)&&&Z@L#3S;^PXa-OW&>FfPJ8cRE:cT:I@;f3(3)6WV
g;4bg8&d)^QRae_bYY][;+>S^_aIAG<.g>&]<>_22?cVI]-e^2^=PJ(e+LP+O^.W
VUc=aMGb4<g=^Df=_^<e0=5N.I>P_dYb\5RM6EHW#fT<<c:g4A_-(AJ,-@N3B0WT
bG(?@e6TT:YgHK[OW/29JG\eXXL?TW/]CK7U4KYf4+/Jd=OJ:18Ag,(1JA]e.(8R
D7\FH2LY&02&1,LPN<((1PTX0\YI8g90;E09.NKRB\02K3geS1M5b?e.[34,IUR:
dWO2LIXaM?dEf?)]Xc]0PbSW2=eeTIX1;(bN5<7D]N<.e,2.#)C),NA(N6UF9W,M
RM)4L3;;/\O/g0^DVSAg4Qc_]L8_VM[PbA@>KV=RKM=[RQ+f]SMOS?HI:[AZ#,Mg
J(X->(V6A4^KVNAc\?Ua>5#D.8RV/&<F]f9I+56L=3)a6_HIUX>7DJVH7W0@HA&2
5c\K78I50/e;@P)S9[YUE:cY902Zf1BRF4:/:fDR9P_E[=C.N:8I/ffYN@fD.R17
_7ZfIM)#LP^0ASH;g(Q/MU5.K&T4ga9gM^MeSZ6&=7aNgb/G)DgBQQUaZ^SII96Z
<F_I9b7(8O-XV.e8YV/C<@56><ZBgd75+CaT[b?S?Y9[N8Ca[IggF(EYU+ZG9XJ3
dB=W2RF_M+BR<cE_(0F/YJ&Y]@02H&<g)c70+BSMV-L/94:Z[N@29H9Z7VO/TYFB
gE_:KE#SfeB6<EcSA&fXfJ&#@=Ub+KS(][Oe2#&RVYZGW9d78gU@0P.8<)U^M;M@
6IXM#d=b,)d4J9g3)GGB<4)\eF(Z3832O@MQU,-V3C-fg&9b@#_[)?98/#:+(M[_
&b/D/cCPP+O3[NZ@]=_aOI2ff;bc#T_ZRY]G4=ZK^Eg?-K:G9ecG=IND[g0U2,:E
5HK&3[IWU3BbU5B:^.Kd+T#5,B2GC#L0P;E8^?2++Sg;d0gFXPa6YF2FSW4#Q9g^
8S)_5OfP^gI0LfFZ:;7;CACg<egK;Ea<FL2?H4U6:.Q9495NB.cN@)CI?d-=\4LH
d1Ag2./A8T/HZ7R-\&4PdRI8RfZ2V15+TC\T>;d-dH5B.M49>HIA,K50>GKZ)f12
J7fS=>aQ\,=T#J8UI&_6CDCY\KH(g[eOCZ/1\[O(>-YJN;#c\UVPgMcd50L15V5[
/RTR1ef)gYU6ddL:6?5+;DK,8;J:Z36Y1,f<bM0@RCF6d=4;(,OLab&&#Wg07gD5
)-;35K@>M<<6.[@G_PE4VA@eTOG;Z;FHgc2N](;4^(b84GCe&Y\g9R>]F8dRfJaf
:c<5.YOg1Wge^TAN#&+TaEdKWY7M(P7LB3HBQ]fKX](Tf\,d]I&^[.Q0XTgT^UaW
R7HU&0R@9><S0>:EA^D72AD/aIa0U5XQg:<^05a>g8JH=#(dPSE=E5;/+P7PJbg9
]_FF-X331B)H+K>fAX8&HH?V3/L@5U_f-;0W<I5>W2fEg,555OL<^05H7-1OD.A8
&EFQ^;RUD#:fS1RIOFJ2\TUegL#+<S\5-]NfSRKJC.PR/gL]Fg>/<(&]0M?HUC-,
MY]:Z7Qg7T28?A-SYQ/G/c_a.4TA#0Db47Z1Rd,1X)0M>#e)O\QRfZ=48U@:9,53
L,).I)4BAa5438MNa1C&5aYNDI+-6T(78V/Sf-e\)KRCXf;P.K]Z+D+\XW@b2ER:
LYHKG+:b[1C52/)B>WT.CJH-XN?aYaD_30YdAPd2BQKb/=8@@D04_YO7K5Qa#?16
-0MDH;0[<Z=2D@,[)245^^??]/A\]/=KZL@0Td?(5aL,^NJOS=8a&cBF?@N&^#9g
Id^J.AAC<<e@a,DF=V51N9L)bbUfZ[N\#5;.f;E9e-.8cG2ZGEOZgO>CWDX:;?>2
+b(VGQ1E-).gW#QNa9d&RD#YZdL+N,2Fc[0UUDB]E4P/OVKO-,6[T,X<KeY\T9b[
92,MWf+5?C^=1=F1&JANI6#feEEaJI-T2Y/]TY8+>EIN/U[X\?&cP4V_Rg:4ZG>f
Q=\dM_]K\Yf2N:/,MQ2Q]NA6AC]R;CM-\0gCLCL9bEG]F1L_D0#CabN4>B;DI8Y9
M;^,_Cb>b5>C.MGMgP,GOAD^RI&X\E2UT0eI,&b^@-YP1V<[KEXX&L.=L:A04(@F
,UB^M[QB)1\.Q+\IfaJZG.+3\Q&XDCfV#e=7J:3bfAH49O#,9-?67Z&FCT7K&2EF
#-UdCZ,JN]<LKD1CYC\ef-(_6)&-)UaVe7G)\a]d5ZSTe0C@K.YYa24Yg^VY,-D_
=MUU)I(83Ce4.fa_g-4\H[^8T@U8K>@O@/D,&U(Y9<L3L[QT@NP2P<9<.Q0WL(ag
P&#/4cd04cf415.gd)UGTOSV>E(75(QcLcA_Y[5OXI6^(((3\7+LF2g]WIVaV[30
-)=L.6e0;eO/06\\GZ4,^E6bQ+LU/>:;\16+EXXcIVC?,#ba/d)a=F13^@/QUME8
6Q07+0Z0+EVbS=KfQ)CHe;Q[R7<1=-X[VPA:EH1ff@,[QBaf-bW/S5X@##3B5=N(
8:4-O-EfSKR8T5HXUK0WEGWB(8UMagae7#5=+7GG+G<fCc7ZdB;]97F63>g_9JF[
D3S;R+32)>cc,Rf+&IU:b>O22FQN8eb1NVQT\5:+FHN^I2)(Z1>9OGZY8U2T?84(
VgET;&5WNQ;:0BXgU/GX#7BgNXc;]9TP8a<-S18:X7K[\U9?bIa?[89\7Q4<cD>D
f/6)(1YZ9bAbcUe\]\<5>O(L\HXW#;U4)3A_,YR<Fd(U0=0RURN(Sa0=6DD6S&8_
cd&]E6Kf=52gECT@@<?5TB(<TV#M?ZH(XN\b-g5C<W][SJ::dP4\LSNd7TgdAD?Q
/=:4Y-2ACK,f7O5Z,A#EMML+93c8(GJS+9^V_4(E]B(]YYXH3LUXcR,B3F+W:]16
RB=/#P4ZVPfL:I3RJ#?fIYK74]6c\W6bL]89f.-f\Nd&gaM)OEg;CK]bBELIK->]
f7?D2/++D(CT42P.>T5b+:PI0MZ91d)[ZV-J,>=Vccg4XYgTSAX]P1060a,+>YaI
e]6NB16d2&.fVb90-O=NfDBd2_)cbg5D6F,\PITPc(AWC)A9J^,I<-.@Pfc65C.a
68-[ZV/60e/fgJ/]LC2gFabW_.7g;5Kf8e;MYW6;<NJ)P/Y3c<1d&L96g;ZGIYGD
fEB^B&M==,&@9+D;9FTDOZbT^378K00@W6eG?0M&IE^N@3RYc=fb^aO_+9,++C41
W7;:g,4gB<4<R=89?->T?)1=SP]DfN/J47&.K<=0JP6W^B<Y;MI0[P;O,DGde31Z
#Y3^(^W[fGFVPPaDDSb6R=53d)e&gQ-52[0-KR6.<SdQ,;Ea;K:BgI9/b3&9TB]2
a5XL9J.L.Z6eFE<Y.eXcFGI[^1c::@><2Ng4T]d/>7J:CPDDH6=&&P<B^J69CBe+
Q?R.LgCAL4H@I?([e[0-FCc6E^ROM?/3/=WCMHUCX@e,&Q<K=XaO+YY/a[H4c.CE
Y#OZ,BZGZ3T[g9dBTMMUJf9-bVBWfZI_EgN<8ScKK)CA)]S(J;MU3,NH];_W(:7T
Z((=dYa4=HKR^EQ[7\(f;:g_6^a\7&&QdPG6^K3V=T__+F=MJD1,.CW1KH6;@1^W
STcSGD3IMP_G&E+60YY65A#RPQ35Nd>R;W2T:HV19B_=bL3E,80)d:\:FeQ9?T[A
f,G_d)4?GYH4.5_<RFX+NEXLDKJ1O16LI88#SP_=C:<Eb+8Q+7UfEDVH5-=CR=T4
GKL?J,O29^]4GP];b(1cOJ2;d[1O9AHBF6A=Q)b#Q81-5#:GG9,1IXV_Q9V@^V@0
0c7&Ec:S6XRgL-ed@TW_:C;H\U><8dI0^d3gB^aVTJZ<YOW4(0,6ADfIa#a^V(A\
XT8KG,-OQJ<c+T1bRbK0@@IeP_VgN:3G)RXA?_bg@)[+J(eK,&aCgfIV1bQ]SO]U
L)D3bGI<=_VJ08FR@#:c/dIO/FYP4D#<KLJ@^/U?8a=Hf?9]YdEX^XC]EP\6)=5K
edSJHL>7EH<D.?#11>65V+I3=4E(I,:R?QF0<GeQ8;fRPG\N-,\;GIB].3C\=#0>
9K.(WBYD48AC.T:e;>V&;\;M@+[YM[#QNWe_>gBS5J:S>LfMC.NKb^&Q@TGYG_&M
5LT1UCV)4]K4aLY\dER^eV[eD)Sc0N:W863B/-D4e0LNF5J2g&cEe2a9BbG4U@,K
aC-G+HCV:e3e6eYBA4Z[OPb\/AD@ZIJS[]aa,?;Je8E9F04,56@e5b0S8]Kd=E/(
I(N+dM9\W/;M/O[\\O]BC&GQU^T)IVd?L7e/]9.a)-)1;-;IgDSW[NMF;4]AD9:.
X21/4/E+eBW87:+N.C;_Kf+8(7&7_YT(5Xd:/6=+:E_aL<5@_4_;05^;S<;HbIA4
+BA11g(DEgN/79<fWe&[.^YL,<.?1DYS+d:(b/CJA(fK\B\/N\Y5+9&TWPa-LU-<
J>NM@O@cfW-bI(K6Gff7)ZK4HMEET,\dN5:7]65bB)1,&O.GZH<39<;^9VLJ;9a4
dPJ24#b?WcYHJO7GGLR+G@-GHJ#g8Q:cN^e1IB7XAQ<Rd^d6)[L@4O=1;JV,=6dc
=DA#&fZ</6S42@NBTG4b2/N2;KabW./@Y/c_44I<+]V#R7aN;EV(^GR+&8CfbQ5_
>H;.B<N21;I4_HX#_;a7)dS;L2EAEM7KX/F\FdT@VO:Z,<e/[7d?J(?:2P31N^He
.W<QFQ2/G_^RIASC_N@]MBU1BQQ_CX)c_55X+T7?[U2>\3V9Cc<9HIU)YFJ3,9KM
)^KeNe2.)W33NA<_=&JXMge-B:X6H:eLLGG;TTLFW7VOYI)LO++GIa7(P>TYXgO#
,K:6B16.I[A)G\V\&?2FL9_=9C.++4f:Q;=TI]99VO&RRE:MKa7<JT)RO]Qc\IEU
<-9-dd]^Y<fa\Ag6SF4K)fJ?PCa,C33b:_Ze&7f#Ie:65N\+8+.OT^98#1XZJXdX
X@+PLA003EgR\T5.eH@U89349GPfDD?:<YEgDSGTQJ7@&WY5=gBOD>cC:Bc;.-5R
ZU73I,6OYI->g]fALQE3]Z(,/<Z/,?@]e_0XCcF=QP+7D+JKD?YE>ZACU]BIc:X^
ZDF6.U#4?Xg8Z+/[T8>RA]ZO(81.Lc3fDMX-Q#REFg-SA)[J(7,35]+#JEL<4)@,
WcN)0T1M_H[85gI@[0@:]S1.,E;^+JEI>L[2DZB2bPZc^5Y=IUDG/=Z7:P(1aAG1
4/).cJ5XbP9VdQa1\8PX62[#P&CXe<+U0&>=7..LG]6<PS6Z0#M-0d(Y;(dFUM;a
BS.FPN[KWLd0Ia\5OF4:N9g.OC<H>3C1UM93ca(@UBO0)XaTWcREF^8bCZN5BU<:
O=TFWXdAI?dO/TA8G+IWGVHYHVU)Z=R>0LG[#<cW2](FG9,e(&UK>B/>(]Z5SLT>
)ZQ=BY22>@#.,c#EC@AQ3L@XW5:B1WG/Mf&3cOSKB475=SbKb53F5RZf=W&>8\d4
@9FD1VEDYbE,PgAF\e+-,#D5]C8732#2\a:]b#=c8R5gC[1SV:WE?,N46#:ZWd9\
+UeR?7L4B6aZf9-B++F55SG=:T89\(?S=S=VHUgGfKJ1G&JN=&-^W].U7_BCPO[L
1SDOD2]/5OX59D]K7LOYf1J#V0F:CRQbF?4e=)W,(b#0IFfOU#[c.H?M5eWOD1A[
GDIR/b&^@Y?_D&SagTRg0?g^,QH04.+KMaQK4S7P]VP#&:3Pc8-6db[OA3F.+U<,
I^)N>UO)U1XaE[J51D.^8+JHUcRZI=Dg<VKC2IV73dFCbN88Kc5XC>bfU5)/A6]F
U(I[U;:\#D^Rg0:@bJBgU-YAT)@Z3Z>SfeV<39-(G];,5/Z.eSOI,R9;IMgdc/3a
b5@LWO&.QEVR7OCKI&8gX-EF/T:ZS+J[4ZP8f1=33^b(^?SBVAb^LT>BBY1EWW@8
U]bPQF-[=V_=Ve,P9[f;)H/?4QK/_fF7dCbO9fc#J?2dK<NI39bHP#</]8aD^P4<
>RKV5W@3B#NCR=PRH9@g^O78]d]6AY;G-cRJ1#ba[3J-K]a6G2aG)0.2@[H+EIB?
5.1Ld0[K7RSN5R7QGbf1PCWZ+QGWFCF(]TC^ZA)3MB#(#Y6,b3[[&e_#H4Ya(87P
7aC#F:LAeU1PYa_,6M#]H/B4]HE=a6,TY/R4EcK.A<&LCL\L&I@QVT_V#A?9U.&U
[^?c+[@_J_0,O)B2OC,b45?LY81Y)@R,@S/[(@OKL7,N.9-J[HN+B?5)S=34S^OH
G26Wb[Ea?_?)-C_b^<e(&5ea)@E>L6^A6C;1K2cIU#X?@/RRcG#:#2+]E5c[/O4B
Ne+6#E/2>>eg1OR(XQNf;<4[,\,B,U.JV)XWI6eYW9KX.1QPHVaAf,8QW(-&cfQW
RDB8\8U_&R/CU2_=YfHU13CL?5OQK[R?a[DX4b,(VN+\65J8O<\>L1>7\9RbFONK
4.O2f[IaTX3d3N#1ZC?<5LY2G\:8#._f48c.[UA#@H_I#_J6fUMHf@DDefUcO+R]
1eO^_L8CKAQ]2d-CBW>ZCd#d,6>#@K;dFcB<7.f7;?2Xe_e8<6OJZED7X\?3KXf4
W?ZHc7U<H.+e8R)HNDD1\4_BM5+.ED[9&AL^ZQPFP?]fWWQe(>=],La2X8U5COEN
L)fHHQ>;@;=2WeEFCcL6V_gF3-LNB64V<LCPFN5(X9+g]#N3]2&2<SEDg<fHSJb#
8TdMO8H=HO(<eE9g][.Zb9I4NGFQEUf/08g/9THC]@4#1OH/(,KHf.Kg.#?ZD+E<
bbO<1-EE.69C_C)=dXKS1^5KT:2RbII\)#Y)d:;7EFA9=Z34,c;7R2VBN2O4WF1Q
85JQNb2=>&AK1J[JSY&#g[#WB#Z3PecN1\4gZeaIZ\=6;U<+K;b]a,Nd\15fXMDL
)1[5R-QJe&@/=dZeKD=4b=S.c)G7=P5#_g+2[fPf/?McQNT5M5[7U#bb/.SB5M=e
d<c0JE3:=?fe12]N(RR_9.2gLTSEWWFMZ@F1:7)CP6cH,9>2QO^]XJZ\Fg0SfN4W
6WJ,WBU?=I::L[(@WLO72E:SHGCg:.aYD2PbQ3.<JPc:(BZ6A+HY)HCQ;=(H@M9E
47I?2YIZ2+]@DaI84e_.R=e4&c+JBHg1aM^RYf-C8:H<[=:#1e]O26+Q]aV^f.?2
/F@4<ScJH8b-J/J.E=@Z^f8@XS+_R#J;\5>X2dg7(;\UCF32C=V975W=<KY?g?d.
46H>KDW=;0,@c#8T.6gL^RO+d-D,8_#CfAN+6ZOLc<WQWMM16gd7L:-I@0_PW2CS
ba247</_=2#f)5^aU^R70?(4/F/f4I-Vf0L]]a1_I:@UVH6?LHRbOa[6S<IF01M:
@C6eHUD28I1#c39Ad#R=3H6+UZ3YYRE07dS^>)B<^C;>EY4Qe=C[NKW<]\REV=X/
EgSe8]5NX23AK<IR&0QH5LEcOH6gU9S(YfV)-/HJKA=4-:dO=^(-d,G^:(eC_ZFU
e?^I).)#?H@ff9]NTFHVXd7S8C[7KgTQ29JeTBEB:Na?UNLWg:3+N1aCa8YHJH&]
X=P]PfgM^<Y^PQa&7WEFUR,VYfQ8a,cLO68V)9:b9,8N(]Mf;Bg6K19Z;fEF(@__
=Pb+T[7cEJ/5E]3E<d>V=.<PD,,^#1>,DD^E),:5EW7CS63=GJIfSM1^M#fDeUL@
de4?aBQd]XfX,=87/>V9S3bAH_-9+P^;aVd@50M:2KA=6GFRL\,E349;eU@gS/0Q
Z_>1U5NgA4S\(<VVGaDM6g=UZ,@_7RKE/,[]@9X-d#.=-]B6=bP\76JT&&[UOAfI
&5?O1ZXc&>/&5#_LCQ#V5CfUgU7dV6E/D_E]@^1J62J>V+g_\3gEe:0a(&ZJbI.U
:]_[\(N59Da\aFRVT_O27U)225TZ;abef51#>E,>@);H=;CbXH,)9[QE&H-8(PgM
22Ne4?#O\Y>3?6/^EBG9ZAVe6^BQY1E(TfT.R@-R9/JU7)>L5^AGH>0@5_GBN4+?
0]TSB>=O@I0WbN-;b5+Z?9N=5WQQf.OC?3d:Y.9aQcL:0e>/8/\MV6Q,M(Q\505a
:QW#cP@L^PI:19@\<S9(KZ1b3]3f./J,02_.NbRR?^ZJEDge]BD);)e<.b)M4Z:B
V<@bB8e_\fI?BgLOeEc?.I=AbKBagY[TY2H<aI?U1,ZZcFaO.IN?B+(aPfT1CJFM
\TW6GQD0#?Y7Q?e(<_[@>#Ac-He>OaG=A_Cf]g,dGc+#5ZBXIY2DYM8)X6N^Y>&K
-],J/^.;6-F[+=#<5e,_7)WY-5V8_Z9a]1#g\[EM-_CK>F_2399dRP^e8_,;LZO/
T/.NR8dc6_1_6aQ;gWIN<P=Z3-35aD-OY-Z>Db>]e^gMKa3YTT\@9+-Q(JI4@92U
e_dT,0&T\LTY5.F\^/(5JL-fYc-JDcNJ0dIAF&d]IMR@.>gLH4B32cMg,HEN?GK6
eF8_DY^3<W525B=+gHNN,aQKg)b,b1N^K/^)C15S/[EB\e#F2PXc1WgCV3]FM8@?
&(_TFA\>W3I,3cIbbJ)IGO6_(5^P<Lb=:=OJDVa1Y_,dCZIH=02EA<Hea+0<P\_O
]IHB/<.cWT^7?/dRb1HMVA_S;Y>B\e,f+<DT+NCB/;)WK/D@.ZBf)eEL=^Dd09Be
2c7LB-8W;&YHD8RIb8ZaE4ONGP:.VW+,I4A@3\#@ZJ;AP?(ET<0gI?E19<K:LcD0
W)7Xb+9UQHHe#c\LcVUc3/BMZI96#(b\NVKPb73ee@423W2B:1:Q]FKf64S5AaFL
^D^WeEUWf59^4XNPdKPZe;C.5_3VY/EQdHR4.18/X+FU&V8:ZeZVWD9;&3N,4B?Y
17_c]fZI)Ba>V(OGg(<#\b]&.dK@#PE\21gF)LgGPX]fPeJ:I::J5:9XfUa-Vd++
WQgMJHG4;g,RTGb\+gI+JE,HS4#\[8fA+N\,#T=\bB3)\e#=J:2NNFeLg7:7YBgZ
D11CGf<a43>;I8(?<DKD_P0J::=Ff#/I.<A=NN-YL)XI)D#7;LaT>eJ;:V\6QRRK
Da>aIS+GTJf\-E;C9>.FF3NNU)H9_0;9-R7L.8BNV4=X>;,A?f@/)R6^U89J\/Qe
fENG:/_><?I069@JL9>PQAgKgW+;9=ESE?SeJV#XP?&KJIUVK=[R4_I4?LG&[8L\
)KRZLLY=LY5YK#L1/bCJD9&8D,-#:7gG<(9G.(_I75L<LUAe-IT8f@b/f9-G&N:4
P[?U\[aNITWTA/?+>C(<&5dM07Jb)+PBe?Te1g\1?Q-(D,M4[ba_5/H-fZ+A:,6e
VA50QXFfKA&LTPBT0BBV<AC6=f&-Q&,.07G;NO_()^ZV7B.VH;:,<acQ7E=NeIdd
\DT49=-&6S<Yg+3BF5GHgNS39J-\c-B>]Q]gP/bF+?D8<YNbRD6b9>WX>&0-fUfe
7MRKB4)N:=R@(/Q0-MGKO0K-=L<-?AF:9eN2Sc9X]H5H;fD-_::01\\=N)J;1=eX
fPO/YK;PG=1_&5I.::5XeBT??U655^U(#U&d#C;ARGE3ADA/;DN\L>A/_N1L-S?-
XEI3abR9H4WQBedBA<DZgd/B.31ERdN\I8^/TI+OLX)dc8S;]?NM;4FfKS;1_^e/
Ec1_9F@98Wb<Ic\Y0Q<8d#=VJZRF(T1XfU]BAfAC,,HV5M?CM@OL[/2?R(B[W9X@
XUBCNK(@:0+E96OV#:-GRGRS.=PNC4)::;^:;c/^8#Y-dXATYN0H/P,U8;UA+3cL
G+C,WML3F^EHG@g;:;eXJK^&/#0IbWY;X:g41)38DIgWgL?ce)W6Sdd[20EOd4D1
)G#/U^d0<INLf,;UB5K]>8<g:7Z[EDB[W./YE/JeG)_\aB;I1QXCad:SB&+,SPeS
I+JdIKX)0,=G#UP/_cRV9<E7+34#f5&:8YCe5=ZT?a5AVd4O@S.N6bUQFPTfC\D\
GLNB8N@4cKIK/K?YM)N\BNeQAgaDfFdCfEId4bP9^<@[E,AA:ge@TN/?f/RcUaVS
=:N,OJLXD>2K/8dSP8dV[)?6(74QN#-Q/XI\:J8;HA65?@Mcb-#b7U[+=;E@>b(H
-:a[KTQ35.M-UHg\fWaJg3XX#FP]+;5K<_ICFXY;O[5EH8<UBf0:cMQ@X#_\BDPB
c(E)f7HS/X+KZVER+c<-aY[QSKP/ZI,+HPf0X]b-A_9YK1KXV+Z+^S7/YE1;G+1f
#g_NMd>=Q8P\L#AAdEWGSK3e:b\GU;CK[gVT2.P1gG^2\?QL-CaZU4VDW[A(00EV
SOXT-P[g+<YLUH3.4<gD?CAF,eVYDNL<GFP@GEO9?UZXe;NE#)[2d@F74/Z6)ZP&
a]B>0E(P\0XB8Cg;_+0e.I>JPHaW4Z01(A9D@NJ)=^\LZV9K&9:F8eNKb0ZBUbSe
fSCPB@+LJ+6a.0d7e0243d\#bTL;A9CWB0953:f,&0OeMcUR(]6&F7X<BNRMT-/Y
Q7.+/>cbQ>bM>31S\P7^FQ9-1Q\1c8UFB[O60?9eU+0Pba9d\f0HSGWf#_P[U.N-
6,UXEJ]M>f?/3@fPLV6Z_a2AS>J\aCB/SGB[RV/#^3T8c3e/XNU@e5gG;B4:AY;,
=^204-&U,TZBF2/?/,)(:9P\-(L&DDe,-V0cPBRJ[D0H?L/e5N&2@dPFM\c)gMGg
/:6L(VAX\3RbN#/2\E;a4\X+B9MQF&7[N1XC+0]dL8?gg.-26>D0WCZY8:;D9S?1
H9/CHBbGUfR4a1..,fK?>[Q\CZH6_::I<7M+[Q)UUQbPcIG8.d05W;O4@Mf\g-FU
ab8G9:;K5[+E98L+03GfP4_;-8QST3H^fed-S]C48:7JfY[+[#fMM:JV2P6@Id5b
8Z;;CRcUE-Z0N4TX2>g#b6EB0ERL\a=?EBJ>LQ1XW3(UL-PVB2V@Bf2P2#DQE]6)
QSJ@#KG8FKWcPXbI.-;\dV(:IXW0@1g&5T3D_&Md@6T9\[0FSGNX/,TX36Q+XTA^
B@CX5;O8#eW]XU&L]W-HLL&ba^8733fGb=bCdO=dcdWb86=/HHS27/V?^4.&STbU
&:)a;2N5d)e.OH]d=\EEZg3;AUV\-G#4CT,^.TG0+P&.CWY@gHNJTEZF[G>5ZFT;
@QD(g_@(R@U@X;?EI]6,1Sg(Y=_7ZXXK9[g72?(\F1EI7.d;1HB2[;N/O@M>6JHW
Z\Q7dX?M[8T6)?bBQS,5XgDePg4Q9]ME2D;7JeBT]QS3/EeJ<?/3YeE@IUS2NDI1
[P>J^Q5N,(XZ=G?B5I:X+eT?,0WSa553bKR6/+-Z-D5F+GG@:^R=?[a<U]S;@YXD
K>Y;-2]Y^QY9Wf6&E<HQ;FPTTeX9)8UU=B0ZZ<)PV;;Z.F@[1BYPNH3C0.(GLC/]
/=g^CPf1]9=E3Y=U^AZ1D[g,;VLK2+g6EHId1Eb0.VRP@+SR?&^:b40<.#^@:RZe
;d-PNU@07^NNRE/GMdP&@\I]-I[@N@L</P?ET1WQa3F(4_+?56Nb=f)G6H@=T=KF
A[2gPOET5.=fO^K(Fg5EM@NgHDe3=7S2>Pe_+WdVb8S<ARbZ/MT48L1^fJHR&cKM
1R-N6WbHKbS.e5#<\)>K#E+\,g[=Z8CQ+,CSTM(Z:PN@?g5gDQfY>g42X5#<@81)
Ja(SO6@6@SE7dDV6a1^;4_^O7[D:3bb.O8;R,K-1?RN@\SOV:6GQINEEW0=7<?Ag
0gDeGHSOAC2f]ZI9+]I/X=_]5Ta).b17_OCU9SE,ac#ROO/DMb.,WgH;0B=X5J@O
b#C,OBdIIHV3WKHLZMGV_:A_WfeQ5Yb4;B(b?L711:4TdZ2]FeLIF?D]LWg<?T)3
bU/)=J6@P#3RA.2DfNgSWD-Y@0EQNg/J3[4K@QU=fPGNWE9b9ZSKKLOPIag/O)-?
?bP[S/4LKT&0L8[]Geea>2>96\MPA(L,(WPV1-&>.F\4,-<;)<=\FePa5]_g=0?.
XDMO03eDXS+A:9ScFc7^S6W1O)0QgISM(f//d4#]d+a,EBUHFb6fOCIB(?)\a\ZO
9g7e@8]F6GeC]PcSQD.^K5D;6e6agJ]&2Q+.)b@f.5YYgRd<,S&V5b8]ZWWN?eBc
/NMB+AB:4aPLAcX\WZ-.I6-TQQ7<,028c<(cT588a=X.4H7E[M&?EgfFEA-Nfg,R
UBI4X]NJ;6OVXO(e9UFb?1U);Q^XR<IG-5(=[Z(1VB0;?&1LK[E,9&MJ[EKDS7EE
?(]@;fYB\OZb],<KT0QV:)&YReT,M]+&I^[\XVE=1M??+N[3e,7^;)c0aA8@.:T8
(CJe\:Y-0:Y&MNM/ECeUcMW;W@)a&6]R4X^bBYOcH#?;BW[2]5_#)g+T6JH<=@cA
]&#gY)RW/8AbK]PgI])f35g.TA0eV7JZP]861VCLaWZddDK[Me1MgS;XcM.Y3,4&
?J>SK=,N)DZcdH[>&D;fCO(g)9NbZ3+S/d^3K^2\X^J<P)R6[<H1:U5&-,H/1PDb
fTLV7V=+U4LBLWe4O9BQ,\GY,/=^7EQf.f<bAL._5EU7V_Qg&GK4QPc@6cRG?bd-
T0_[b.)/YFF60Z(&3SU+Q20QaQTBB4N]R)L,F>aHdANbA=Z<PL09V\Z_)3Dg77AZ
G(EbbLYS##@edS)4/gQb8)Z0U:-LO8OYIPQ74)]B7D&JDUaNA[Ug4g.UAgVb6]ga
0\H_A)<V-B;U3=d+#Z.R?9cb7UVY9XDJB(/aTa\b<LNAeZ[,OaE8ZMVW55?.#6SU
gM[BH\Q^=4AE<2UDXEWI/TZX(gEDJ4>[;&4TUU\BgE_+0-gU-(NYAI4P7Xf?P<Md
-9J,0=YS1X>JC6?TKOg:@\U59DeQb.A[A-^N#bY^B0Ng;?.UWTXH>d+[dUQ3LPTa
3?2)B\dP4E_IfL-Q[L3^1ZAUfG3DXB0OUb6R.ZQd^NfT#X35T+N0?Ef4ISZ.C(7d
VVf?\YcFVc&QHJM5E##R8)?)TL<bL8&[4&b,9K(ff6-+M&[8aE@>NO.LWS(O4/[,
I(fS_>1_9/af:602T>@V8_F8Y+AB6),=2d0=>1)IXgTL,EPG=F^6K;NW=)WA@-<S
200D2aJC(bbLN3>e#HbP]X<5EG#&_2SN67?c&fR):CaG.;Xf&#ZQ#6HS;7J/DMVa
\X,0YUELK\DLCJ?\ec\bSTL(7K5GQ_16K.;AJ:e1YKK,/CLd^TI#.P-M6ScLbVNb
YI_D6;AbMA6TcCW+0Z9P/P4@KV9SSG.f+@RVcCM93L)G4\Bg5(LL-H#@/@7@@\G(
ZUT63#W4?)7A@^7#C-Re#Da#bHKd0;E/:VCX\PF,6]L.=.Gg2B=a+9B3[-c_a..B
,MMe;&T7d46A?cPcE2<71AcW\_YN<4-[YA[(cL8I8TBQNT-]cO)E])=,6e94]8]0
6BR^/S:Z^2N-:@b:8ScLR_2[=e9+CbgBPg#<X1VX\A4W[\AGVL)\2Fc;?NTJ^9O8
)BLZ=SP:g:+#F_-:/K5^R3::5BKd7QL@;47fZe9XeM<7Zf>K4K:\?7TdNA0fKH_7
H?+/V1H>E]2G_,Q(4=RV8^@P)W9.=N]TPF9O?=PM)+^F^N=RRSFQE38@-e8E^Z,D
/,aPKB:S:FZ=(#AK)8d4^),4IMRLW+Z^LI&R;XQeWF^^-IX?dDB2E/YS.<H<.5g-
7X,1&SO\[>.V#bKQ^dN>3ga=2.B^d86[/A@FUCW&MW)&31E^7P;gVaQ#@<4Q@-B2
GU?GU9IgH,9?cWKLV.Hb1\O:a91,KVbZZ/JV[<Z;T(Z)0I)D+8JXB:SD3XIXE6DT
=&Xf6ZB(<_UMU>5G_\MKEfVLVX;D4eNP(A&_bO<JM&eHP@>&L=c]b,TB&7O86IQ-
\=?Xf2Z0MGA0BNOS(Y1A@\;b)4A5_X[L)&d5+B0-EF1?J1(FS24RMD(-ZJ<aX\M5
16E\87I@QUEK<\PDKAY;K[-R:5>52R3F:U40e6/bdBZCBK]A[V9c9)?,eAHXFILM
0-XV9,F4:[g&W]<A57@T&;9X^-K>69S\\ccOEQ&72/a>AUDc1@PMPD@EcGEO5<bb
U>?/EV<LX61;bDa14FBCE/-LSeB4^W1Gg:C<Ha@RJ\_5NbGRCaZKJ[S;@\:-D4fb
3DO_;QT;?GCB^I:6T,eINOK7K^b,6GMdbVdD/9+XRJ?.BCLa2#1Pg)+R)X<<HZLd
X/NIO4@]9a0JeXcFE=.+be35R.O_#5>:=E=K>K_ZE:^6C[H2aQSG8f7V/5Q@#3\W
7M=HLNX@E\E9ZO7R,^DgTe0XL8_V<WAPH5f-:NSOXfQSc=^Z/>;^>+GNZ(C&>aQ;
UO^3BQ@(N/J18KFd1TeR&\V<Sa/SMLga9#@Ae=6JK30g:ILJ^+SdH.Xf\63U)?BG
9,=(EOQ@]Qf:(fYfLO#TXS&)VU&g?2PYg2:>Q([+C5ZJ_.4d^/f+>,[Z_7bOf+PP
G>OZ&8]_+#f^S^QYO.F[@HUg-R+(+#UF^9&&gEa:bXfJESGSUQ<7HW+BOfbYZ/HO
>M&I=Q\H3)f4eGM>BF;_Q;0Q9bCJ8RQL_/YYISgCF[ETUQ9DcOI@KI5ARb.aU7\K
^6g1dO2X9XV]+F@g5Z-@XES-<TMAS36RT+=9>\V[>#I9>1/A6g=UHAdS;-W?CR[T
:YHBSA0PM8DVUFRf1M]Mb_KX4;TaH8f(7.@E;S&QW(]GQNM;]@]Y>.Hd&FW<fG_6
2?#W0&/cE=0Te6SU=NS63-G+fA,.:K1#]]&1WSJG;]F4cH.37&W>R,\3Z,53T>Y5
M<Y;+d0?K5;NL++A:;XMV+YUUVe>MTGf]U9Be2-?#:b]^Q,Fg(3H@46S?-gZG<^9
S-7e62<VA@<#+>E1VcZQ7\Oe5ZPGdI56]7H9[O>K+42g]:U5?,12W9;<L,4M]7UM
&CY7\EJ(7HT+:7KgO14c2+(S,=f/J\D+5.5D[7&@=#c:J][bO0^g,4,+=)T=G#fX
JAS,KQJ)&Nd+3eKHIDg87>f#9Q+PI:B3XfA8gg]M^gd624dFP(cW(?Ef;2ZeP6HI
a,KJ8URL;Z7;5([#DM68\_[d7cRB+0)(-YIa_K289;&^&ET162X.fDdeIcH1=R^^
IH9358K-#M;VdMVa@YRP8^Yd+WP98PaPD1I9G/PcgWXH>Z,98AfJ#L;dQeKD)AF\
)0bH]_A?SC+9=O^a)NG^cT+3;4C;KK_(#7OVf&V17L.:,H5:2\FLa9EU[ZJgKFZf
C]G/V\=]H:A.OQLdPMW<QI+J2OVBY#-eg&#=d\dZ(Vg:L/:4WX4X_HHE0JJ2g=@,
2c,9EH)edG](dBNAD;ABLJb)-0P&V93BZ_@KLV.@=:)UK17.D>&>N<XKH>NRBIJc
a.D_K=Hb_-&1S?SEVFI62-0/dPIAE=]M?&W=4Y7#6.QI/)H.:^VSFC2=GUR\(bgP
(H>>PM,.WKZ#g1O_N1?;P^f<,R70DGJ2K\(K5H9U#(_GL<I><:R)CX50YDS5;37O
cT#-a+M&/eD?;_G/1#RN>QfJQ?O)=J&HGE^?E#BTge92(LI]EX\A37c2DO4V)D3]
[b_I:N7fL379NJ:6E(<CL8BHT9Z-]T6b7afU=&1>O9&SFL9AB(@PWgJ.ZGA?QEL1
adXPE;+JgG(>,b;(=4_X^fg/=gAc^R]fgIdO]+Ra_/bY1&,-]HGP_M(SZ^M@>6#c
QP0XW(eYTabE^>:[_/;B-d4JY[aggN2B4>O?)IURb4>F=@>O-3f&(CT8L]2cJ8P(
bR[QcK34g0IMMFWPNO>L6[NF#T&W<^<<V[XZI999&7GP--GWP?XbC9#48G9Z;<PX
14[g@c4?)bQe:[Y]QTXY_@^L:@>5K>BJ6Og6(Qg</.RH4dFG5aYPbHF1=^A:^dB:
R/3>+^&#T+6,0;)f+e[b&S;58=N)>K9=)66DcHSL&-NSaA?G3+@VHQ?dG>^/)3@W
8f4IP<;H6.0YH]H,)-0KfGQYVe>K6C>9dJ0KA&:/gI@+76]8,eRCg^Ta<bV:3[D+
9DfDd)[U?(&-828A.T9+VWT/9@BK^_gZ)K#27_1X.^UZ;,f\,e9.BG77X;0c+-J8
?KP.DdI]3]@2S^=gB:H/c-/)deWX-EY3:YfVRA3ge<S_:A&P4A[_/A1^e#M+LU<[
U[68W(2&FDN[fM/ZW],OL1MJI2&T;USea]cE0da65)9LGD)JP3C\;OK0<0O6+^MH
UMHDaU3eSQ?N_P]TDD-TcIM>-g1W^,;&5PZVRKZ@4RN^.]\<ZB^M=G[)&(2PKP2J
[+MS-DV@0]0cW2Z(/E)]JaG\a]aSED+OcM+8[F>02,da[3I#-;#E,?+bVUabfSSf
7)ad,(9EPPC=(.:1f[UXAc:)4A4W(7JEH2L&2[D_YMe7AMH7,^_.<[RH9JK=G7G-
B5SWNWAT?^;J)?NAge[JINBe(R1291Te?DWG\VW#?5)&.O08dH?=(O=&:IbI?_+Q
L@BT#?C4MfQaLRfM=Bf-JF8+K]9H)deG9N4JF+5(0@R,4_5U1\CW3_XBY5FTcNZS
TN+SIeX3f>#[fL>8?LTXWPc\8.M.P\\6<3NG8=Af780(e-I_4&>#e6<RK@R>BZ#<
F^NX#NN#9MQdSEL&)JPS?R,\AS\P].ZR>5fcfGg&-J6/R(C=()=NBb17_G])DUHR
03cTZ=/S6SD4>T+6WC[T<YM/VFa\[/LeT#acUN\A+]XJ@6ZEa[]/CTc^:DAV4G+L
9:PHM0,@d&5M0.RTfg2#>=9\Q3.B@W0c[40=a\USJ,I(>C9)CERZgLfb.g3Z_Lf,
WYMDLE=_SR[JRDV]:VZ0T2PA,ag7>7M39-\]^7(C72Gab&f1N(TQJ@e5;fB?,+\:
8:42U84W/OeUQ&cZe:#5Q3g-QW^8ecFf)1YdIVTXD9J(OI;&_,Ff=ZA(4WL40/J=
cWa_=TI4MY0Uf@7;FLQ2,KLHBD\5LW;VJ5e4aB+?+\56YcZ+d@((Xf#:DDK/E]IH
EWf?/NYd5O,aTZYSZ0Ae.^2S.,5><8;OEd-EIF,^+-M_IaBRH[NS3AF_+FG#Zb<0
RVU+D]QaD#6[]/UMeCH8-S6E4K8)?IM.#[W=&Y5F63.S@8BS&<\/UTfLMaS2K_Y2
C@;D&#-2aYEbac]A/082K,5+<,SWQB8OW2K4AU5E^IdF,0B+R7XJ<@86d=?]3=?4
N)D#;WG<C7Q:T@=P2N,IC.4>C:c.0RN/dF]7-K0J9eY[Y]E@W^?2BJ3],D76Zf^f
D]&HGacP)KDLSBZRUAU5S6Va1Z^KTYMB:,B&[RSOW/>X>8fX),;85E.E\,@QSb/R
R0Y??e.4(#&[b+U:RE>9aBU<=^NQ&B>[]De_ARG8LIcIE;8TP65WB5IXaa^e10d5
0[@QaNHd3^W<RLKJ.J@9-QJd[G]U2M^-&T096\TH+C3U)/e:?d/)YE]SKEMU]3]3
<dRVd/&//X4gC[XdZK=S1/>I:C3.#V6<1:SJ7c[ZR[B5IDA4F_LN?Q,JeW5fM(R#
SHZ)&0V:A]I,7KD6B1MK=C+Tb0fMLSEc^:9V6bFM<eRI/PA0P=)2ZA/31=?I[HP&
I;&P8VcgS2b?GP0[bZZfK/f_IS[870d;H_fGPAF&7MWCE<NQKBIgfRW&[Xc(\0U]
O?;6<<O=9K-e2H)5=dU\M6E_>L/9OZDf#fg/DOG8Y<S>g)9C3+RN8cO(6a7^QI,c
<QHB^edR-GQ(09gTR(b)]E<&fITXN6M>2Y#D06:,#,<0@22PQOU-?U;W<[-CV8e.
U>#Hg0UE&eZJNFF#@Wf>M.P_1\1=O>gNQ1ORP4\ZV_4WYBGEQ]DaIK\?cfT+A>B-
?9KR&K9N7e/8>>1@1R6@K+])G@X6(SEVZ9V+?D5YURC2<=bW@2;3X[.0UNJ8LgLa
9>X+d_cE/37QIc6\=<Ec@_.H0B5b<J774be,DUVC#^Cg.\)gB#U9&Wb5882UA-3;
,ec-Z,FG?IQQBPE3ZP-Y#18D=7)fa;,c]8^WDR6cg4]:8E,f<OFG&O+@3VXS<;Y@
aE2+].ZQV&-1c.9IfgPD?I-0:H_OLcV#,A@Q-Z75L\55?8N&8SbAaI>ReO@VS1>M
cJ>2Cc7\Q^,LG96f6>>8][)&L<6LYKH?)XQ35Kf1L#/aUL[N/7[SL:Q)3..PcT[1
Xd;a9JDQgdfBa/#0f8Fb\YGZA(,GGC-4J4RdVf_<J+HY72=2JXe^gGOcS9L=_P17
@EAEbG?G&VL,LW0S[6;M;M=2=H><_22@OQGZHHIQDO5WZ(1MW3)+T1>>U^ZSYdYY
g@&JNW<N9NWJFOc=GQ>V:3,().M7OUR,B_eD.HAD,)D/W7d^SCH_5fCT:N>TWULc
BT^T[)/b0]8YffCBGJ57+0W#YC\2&4#T/+?UWECOJ?0]@fHg/JG25R_#YZAb]+1S
gT=AfC8KLR:VIUH)HJ-:fR)W>c(A>,8U]F5@X>)5g6102f0-][e8;Q>6=:G?\JIR
K\FdadU3P=PHWP6MVQASP]PBFc:5LK]BA/U-62dOE2K+&Re:JgJ2aPQ-_8>A]>,G
+c)b1I,L1=:;RYe25cJ3SN0D6\@/9GUIG2/?V;3O#U,1EUaBWJP._f@862UGe^//
GR?a5S6:<f3W).IZ9A_B;-QB-1=SN;:;JN3=GD\A-DbH/Z1]B-X6+(W8E.G9C-e.
bKT@ff_0EPS5YRR(e7a8cOFK4Q.^@E9Ya-DTXdEG&:U2V04<+g5PI[>Te8C\ZJP=
M_I0eLC\)ebX72BXV5Z=>Kd&4PN[71U5TMR\#A6H[YA\-L3:\/E2NAcVW5D0O)?/
?OdG)c73B>(bOBf3D53PbeHT/L1RCF8K.297S/^cX,?>;gJZ>^7XG1#9U86\NNbH
fY;MNDPT4Q]C=;^>Ve1_W6A:IG/#O:d/Cc]OLH23afD1_5U;,1A9]KTBLJIN(+GQ
N;\1;b?eVD3<I5b=O<f1f>9JM;NdUV5::3Gb)<0WR\8Yd+]A=;T[dV_?cT4FJ^W\
=;AD<[(NeE@TOB5]&F\BXbZ,93]\1&#df3SgGDfCK:fdEc8RS;VQ[GQZJW_DX+AS
^6E4YU8f(2#E6eeTLHEZC@K/;>-I8<O@^M=&/M+A+g#NW:Fa7?c;0#O9UD6D[BAS
O=e3;_LX^c93.bJ8gcN1Q899+E:7^T>;DMeN^8IG03g&EW_)YC7[]Gb/]d\NV<d]
8CCTd]WJ,C4NK&/(4HR_D;U:]EDO&W?R:71?6e/FNf7ZAYJARfDQ_a.[#3[&4Y&c
ecM3MQCT;;-a8EHXF=KZ\IS@KWZIFUBRbQgFcea0E[g5U7M_X-^JI#T0X.ec,PKJ
WE[?3,OM929VQHPIET:WJ(<DY;g_G>32/.)Y_Rg]IDWU7&WJ8M;.a?D:J\@fI>\)
ZS(D#9M^2g.YI@G/O=d25LYM&TVY^\EYAH#(a]ccd6YNP]Y[@:S&EPJZEPV;;4KR
:]_#@(fD69>?Cg/-b5eC?L7@5G@O]gg144)2<]RgIdKd=df(O&C9+Ea_D0;b5KZ^
O;;.KC;V/e+,<VbH+g-()-/5])>)5eBe],Pe,B;,2)EJ@g#O2^\MU_6\A)TT_)EE
^8>dY9<];6a-KQ(=YdJUJe+\SNCYL-)^E;b>-]cKDU-ESDT6D-T-_=_cLcf]MSWR
L:?4ASAK08f4d0O&Z7@+NJZHa4?d57XMD84AFeNBd#,J39UZ=ZC;#_;],TOM8BZ,
CfO84K0KZH>QUU3/73)Q3DQW[FcSX87ZdT:A28HNKf@-[6Y&5VL043VC=06Q5?WF
^W;^VF><6dg9H#GNWPfb8gF),f^/dT(]>O,fcbC]\O0/6?4BeXXA=ecV2WefRH.,
)_F(48][G\FGIL>b/XSJHd#TPAHC84&,eX9Z^MXc#b)(b<(-UbQ1;bBB7-RDO2X^
H9DH>E9MQK>(<c(U/_dV/;c>;75c\HFOKW[L7.Rg-0A\[^R>@DE0R6BH&,,?6NRb
1fb8#>60\8T725:&bR^+XNb./@EB^<RP9Q#@f=;JYdTP+=]T0N&Tb1J\VPG[W<0P
T=0WW\5+Lcb3SXKJ=5,BN9<5aWQXY\ELGbg>cPZfd55?#X>I?6A&.\CG[G8&XS]>
-Y8C,O:CG1H),f0WQPQ6O0=F-P\Ig1RG?MQH820E^Xa(>Z4bSOD@TZ7L6<QS&@1,
O09e,]7eJ;KVgeMM<4c@gARA,:L@^#M[\>0,ASaFKX(DYS^UcH]DbOL=);dL>B89
TW/TS@T30A^IO#A#=g_X/I&A[b6I#eg)N]:+O^VF>,8):L:9aOL<]\KABH0MONH#
eHA;5T5,LWD;17OC#MaC/6)T<J:=gAJbR@L6<Ye?BdD/^.>_0@dDed^PANcPMGAF
^],/[J8X+RVNY<D/X/a.VXQf)7JgGD:bR>TRX63ggSP53fL)BJT2/b&>\AGC0f.L
^N^[XI.)Ra->/4VB<ZDZ#.JEa5d5EH=@VTCHg(/4N\-ACb8cP32L=g9#&KfbNbfL
cW)BW5U[+\gg5:TIA]1g(:X<]4-5^[O[,J5]X54f42Z7f:fDTGNSaF.4<,J=B>\K
CJ_YEFTB9L/2CMW(aGW\HEPP?UCeU.L3g5)9D.&,(ZL55Z^:>NQ\@]H6G,7,YC:\
,H=Uc\bH<RIVP.JD_b6UJ.<Ld<=0XLKER5.O-YG.LQ13g)5W63Qd/A<PIL_(?BF1
EWHH9#gIVaG]@5GP0WfT0CJ-G&Q&f#O^;M^>@I8S7f+C8RD/E/R.^O+&VDJ^.OQW
_-.R8Y)AbY9Y?=d52abNDM+B4@[BSYUNR6(J?8KV=/Ea2@Xa\(ZB<Y7[^BF/B(@]
_M1F/e(/:d(4;#@Ef(8#d=>4.dO@&^&0XG-4#5V,I6HCaJ.-^/HacdL=gAVU1PYC
3X<BB;2\[dS)K-M4:c>b&NP2=5)+36;391S1U+bS)OIV.Za]?^_.?SIfWZ&PR<OM
I7c94)+8,)/;5YL)OT3];f73H?fY=gTg,#=Dg+dSec7-f)C-/#>08DT^Kf&@SX)]
g=5O3e\#P50bBX^(Kg9+dO/FP]:F]@>:-fYA9_01gE.5-8W0Q#EKA;E1ZN=LOT;=
9H2OD3_N[S<fOS-J13F-U>dQW,31DMH^8Q=:1;eUZG54>=__>Ab;5Q;#;fMGQfYL
/S.-=bDbDR<K,JSI6KJ89,;3:+,8=9S5THM->BD84MP[NU==P-O/G0fAIEG6JJ@<
gVb-cI)(Ff(6)=\ZB&.POYU,O^e83HYN>;98XGMA4TL6P13NES+:/?PD)F8F2QP)
7FJdI6dA^V5U90-H?761a8=.)gBQ_>>K,VO)^>?_^P&ad8X^[_+)9.WL=9,-/4PZ
&8-^FT?D91P)Te,>UJE3<cWK?#ag\,](E6a@E=bRR]L8._.^OAfW0S7c3)XY9YXK
+3UKcBg^c5-O1E]\P=N>?Ta,_M.bP7CN]bOX;?cdD/b<S.CVO2<<;6>]<;AE;gY:
A3\XBY)c_=1=V1:G3]XB_W<><Z.&T#BN39ff5EB__N(#[9gT>c+,5G1YU+?@V@fB
6WgMf<)]_HJ06G8TPEUBPN+18LYNYb;bIR;YI_-&,+3\>c,BETP7\>a\FHbX@c7A
E+Pbd;4()<?H<JIMEee;:87@GW.95E]0fOUERW:BRXF4B-OW9<YE^U@-U^8&?A;C
D,AMH-Y:fBJ[W^1@a?V=,QUG@?:<^L1130>;/I;,dYE^eD,\W]TF9YW/M4K#(@H)
g<#3END\-NP.1+I8Yc3,@5?K(cYP8O?4VRT6)NMX@=G]/^^F7GaSC0UG[.ec[QF1
G,\AX\]WC:>VgK>cMXD.7\e97a9@L\7e]@;.FD/gVA_YF&]FC;@fH)ZJ5M7FM[Md
XA(;33#PB&P&UABZV?/CS:85a@[TQ?aWKd26V7#)P1Ae+e2.D)R(8GGBQ-_a.eFG
^MJ-7JgS_U=e9dU-\)SQ#:?QfTR8)U4TYXOaQ(JZ^G4A5?O.9&RNNWC]gABb]Mf?
E25Le).\fY\W[1dX&,;&>WYU>TV]TLLE:fT3<6a)1NKD^fJgJeU\:),fXA2E.2)]
@53?L:@,+^Y1@/eJPVLG;95JaD;+(0N4;1_[8_RL;ag[V2[7F?I)QB?6QYYRb3H[
9>FO=Y_E5S/aV>K<0LaY=@21-8^Y]E4W^D7?]\7VF_Jd0Mc/2URARLX6I7M>>\_T
EI:7O].=_cb)#P/X+bcS8][8TM]I:e15QY;SOW7=3]-E.UVL[)@/4N=N[X\g3TGf
.)Q@3)DS@eQ5cZEc64?<=UXOL?@RAFHd/c@Pd5E6@eJP#FPCI;F(RMEgTU5J3N#a
<89\[W=1Q[+VQI2U7LFP&];f<:-OADCM(P.PbZ3H<LM[8I)UR3-dB4,/HI<P06N[
GM(/E419K(3TFW6JA5C/=Nb;5DGdD9YYEAFdA5;&A8_W\GEgN.B?C]a+E=1@S/Y.
])?e(5<+V//<a(CEa8,=c:\IQY.[?+^M3TY-[]7VHg_^a-OaC2gY7D?+<G?]Q#G3
LF+:]+3Z_7UH:10RH<G6/f<HJ9dQ:6gU:)@>O.EMY-N1;e?F\8C,Q&;?AO?^A<S[
7\)aAC9D-UEPA4<CGb)USVIc5>CQ97L-?I0&9ANg(@01Qd)?[6ANVC0]V7;8>91J
WX?0HRRDLG&_D,K;HMG1<9[g6\)A=Z6_Y/L.9],eS1\DV=X-(&c3gBLc[W3++Ha=
Z8]3VM\FC:f23SL)KJ(WDa/;R^@]3JbGB3NDMO5@K>2B>8-/3#cS=;b7?IFgUa0V
80T2SFIXH1R_KcI[NYBf88a0/]DIWfN?HUK8Yc&?#_CT1fbO[PfPKF8,)2=Q?/gZ
+C[=I^fVAZ2<J4d^J=^N)8BAI=9dH(bSFa;JQZ&a+-bd[f6#&@JS.f3(IRO:D2(Q
EQ78b>P/I-+G5a09Y179?O#Y8c=I=K9;EVU?a\&M&D4_,B.RUU-g(FUP3K#1^[<C
=F1\P6)BYFea(D,a?DYb/@.WG=EB+8U-,9HLV/\Q:Oc)XNP4Q;BeSRS5K-ZP6^U)
8R^2A@-_3gS:R)41CMND;Acg\[7.O1?,Z_DP28[5f\/URaP-)9^HgY^5bYAMgOUc
]Y_aUT<_N58DE4#P>\4NE88I@(#G\MeF&\Y4,6U1Ue-);>:CT,=WH-_^I0H5:X:W
6&EYD:Jd.CF>,6c=]]g&VH=<cR19b1/B)(OM6^3U,c6>EOAHL4_LJ]1;dDIW@5b:
>Y+:MV9QFa64WYS4U).ZgG9d)U2+=Ue\6P)K>f;>,KcKL)@7c)eJ)Q3.;cAf:eHL
dL8;NO&64g(C5EH3cS3#<EADe-0a=+/5DYc-?4/JQ7?)dKN.UTHU&FeV0W@N<R0:
C_8X\NRL.KZa^Q351#1<^2D4+#=M\Zf^0eU2Z,Jg[<7<G_VA&7W97LMaP/)37N?G
7a_A+]ESZ[ZU@)M+#Vg8T\dOPK,:FHT(4I.N-,8J?]/]1^]48(2\]HIX>[)90EFf
Y5XW-Z5?S);YBYF:1]J9CS.@dHYBA<_cCBIZ&f8/>YU4Y#N8IN?cM=Q=4(U8OMGf
?ISW6T7Q+]6H[VPL-W5=O3^PRBF1J43UV1NLgBXB<#3;,Dfc8(EJ)AD9;H2YV=35
9)YK0Hb\<4:E9-18Dg(/T/D\PgWUeO):KZc3MeO&7_O/=f<JZ?@7/(G_eYKRe,.9
9K.3@Oc^K#MF@/0^(:c<49#gRF;YY]gfN.=^6_eK;8K2ZBICJcR#CAb+bU)>KU7D
f0NZ4.[?75EM]e=@;2>U9]@UB4>\-&/[.C3E<=RMdcIUE6Z,3@bP7+e.Qd&LGK]B
5(@/G.?Q[:@Y<GAXG_X[19a>T<Y/g7-8@>)X1FJ7g^Xf]B;DY4]MBP].PF^S)(I7
e,574:NZGB)FOI^8.C]LV1+TA2YbD=eA1--cR&6\XZN\f)PQ179E1L)-Z=U.MQZ@
S/aK-OK0X\&8Kb@+.YD>P0eSS<Cc<@3,?CLDG;)/->E.KC(&F:/WW2?,>2b^,ZVQ
.aB/:-?K=EJgY+358YId2dTOFM;24M@5eDIeR7ff5Da>I1ZA8Q\3I?<0,c26)b]D
?29-94Z#:Q/)#Z?IG<1_-<48NDK7ab<c.[K78@TJ]+CI@HZ+e,6g+KJcaXTBSYYg
3FH.fGMbb]LYT:[f0<_]MFB)<99=,=-7c7TB63Aa5(QIDF@_Y)O()H=2PdX(AYR^
+L.JD(H)NbZ@H-gR)D(;_&&fA4NKA=+8_WDRE^VEE2g#2TT>KYd1)C8(.-4+.7W=
4KN46T<#-#&D+C>&fSaX696-]O6#UJfBVHLdaI9+7eF[gM/6ESa>MQDPSQdQRNZ+
@B-QC<e,^\A\#22-K+J.#G)FdRIDfg83:G5^V<OC.d\PX4N[9#U/(U8--.:WE7JX
LO,JO?J[S>7W40Dd^dJX]0;N<;20YUU=-g:PZ5NW8O@C++Hf[;d:,RD,>^6(E]+L
J<\EDW29:1ZM1[@^ca\DQeOM@C=_1=W67e,7U1PKKgcUL@0>((aT4<M;;Rd4A7Lb
(CKDCMeD\)>;\Q-QU46P4-5M4Gd,14OdY?+CKZ#e)eJ(\6#S;-<;LfNC=LDeN[.;
)&e,XRY51cW&g-SN?T]./9)W?[4/HTAFVM0Ke+H>-]E=g.G;)EI]IXGAIQ#,A3&d
0.RIc7@Q,/G]RE&V[WA6&^g4;WYA5U<b-_B?,H_]\KT]:U0\6V4[MCI\(_-):bA7
>23E[E^4).8a9?RK^OZE;P[78Q7f1VUYVdb8APBJ(RU;OV3R)TR_5<ZHe)3[9(<C
dM.#>PT(1]>\/;UZG46<2IEMN\=a7S+1F+3@OE5^MGPf/J)C@:RaaT47UVN@3Q;d
[#]@]QgF(VcS02cDd)(V2_(UM=<2]XCJd/eYB+dR[BK4b.NB<P)(;@3Y[:7LMeJB
;U(T-d8C\0YX0^=I0#64KFAG.2Q0^5a.WE^WG:(^R/5PPaYU.\]:P-&:0)6>4Gd7
b[eR[&d13S#(CLaB-F(XQR+bKK(d+]]Q^Z(GH]a<2K84+)AMIf;,&Nd[9[W)2[[a
=9040Z-1a0Z)B:WKdbOI;[^#Ea3V10UNDagQ1Y-3)H>@X?58DD<+I8#-WacTE6@T
E5.(YSH5V\a53e_#b9#8:d,;W6(Ie78=(C.X)JcEH)<AIUga^7,g#J)L_bf.+>B\
W3+GGFcJDfSf^=G#bEa<J1DMWMF?M),eID?UedS:XD6=(5Z+4?+9efUYI6D;Hd>:
:a+,OKecVM=bSZdMQ2E;G-_bXJ]\A.@@5AL(HK\;1+VJ:&K-Z5?(HK<(3,=D1YW-
21&D]^V8dC_HTR)[;8=7X2fEO^K/PVX/@EDN]U&1Wa<eCf^gBg_HfEXGQ0@a[#2g
&aX9f_GJ[X\O.(ZFHJ#9:Y9WNU8I=939c_T<Z<g>TEbI=O_4-+ZJUP-38,;3K795
I^1/cN-<SgPK(T-UW(d8?5dF7C98OWN_Zd0X6[6Aa#:&_,fFZ277fe?[C10eW68.
?f^a]OH8LK(fZ\EP1TGYb63P2fF#D(_M7@F-:31g1e8BX3.>)L<+>12X3VTMOP03
c-[&X.HQ2+])HEL^&02:6.?Y=4>T0Nb(J,9d7:=A]d>:J/@)5@=cPAZb9;f/8B>d
EE-[B\<_+e(a@KANTJ-fE4^ea^MU7LcV4bQF\PO<EVd/MV+NW&RTGK)=[@>=a7;,
+V)RR>HCTVJGdKED1@@N&#b1M:Ha?C?KWbcVLPAHSZ+Wc9.Nc.KQ)2LIc0;G:<Jg
7CfYQ<6--@#e3UNRNKbU=G3dD<FM83e[BAdf)b&P:9PI(;>4NE<4PXA=,WENS-f\
gJZ5GB7[Rd/<b7S./SM3#B2JDIHJgY6-=8>EF)Ja96dC\g]MG=Db0).^?WCS>_Z#
AS5P.2.PRWP50.U9BGEBK9E>VNc)[D\,6>1;^]bPV^Y2W^N8ZR?#2b#HNFCL;Zb6
PBI-BBRM:<^>LJIU4:MaN3d&&^D+06ZBM&<6GMYaY=P0NPTCeQd:gfW<@@0.KP5H
F3?c&>==]dA)<588TfRM:0NXS-cef?^G2\[fJWITBOB>=)61dMT)F64/ZCPbKgHZ
\\Q+La9H#<:^;<TDb[0KgPe:.N^WAYFe,?]S[O#:E>&>0INc\4[A-B(.KY1.V_e[
1D2HP.71Cd0)>&8b4:P\-1Eg(]F8U5bF?P2]HXNNO98gC=CUH]O9WO[P4;#(&L79
O-ac.IX.WSMYgRRE@ZO:??J>>2P]a;WHF6>:AWS4Xa<;1G[-K/1U;Q2/FK_8>H;V
eI\-fGIHVZZYX#f>]0223#8=MDUB(=Y75AZXHYC</8C0\D>+24S-F)d9Ca]JfA6T
[0(bH:S04bO,-@E\6G[;WK55eVC>3Sf-d=CeMQeBBXMJE3D<)gGd/K4cOU^:)95K
THAIJS9^=0fL5c[?#)+VG=d/@-<1.JFGQZGXdXO#;L.J8+^^8\,RCF(+AT[<JX]V
K>7>7XU6GTFY5P+KfP&6;U1SF-.cQ8/(afd^0]e4Y\?8^M5#6_IB]LLP,FL6Y?6W
/F:9Eg/cd_+E@g5Bb^RYd#,,EC56g,+XU3e2WOWLT-N39da^/-3VcIIV9V(CT9B@
LIWgf@V9#U&e]&YBJEf.fX?N(A.CEH#a7BM&#BI0+[^WFC3&:IZ:B<H4cOfb8U3c
OKTY>F?TQWLD2.g.:VWIPDfLVR?OE(,-BbWT[#OcJ(J(,HXQN;^G/#.]^;N2dT#G
dTa7?6.P#5<Y^\fKGM9FNC9R(bdSJ@O.7WW^5G#SVZ5SFb6d@WG^.)>J+)R\aVf(
@)I5WcB,L+_b?f,RD:;YFC(6cY3V[e)7E;+<:ROPQQ;0d)6?BAU]S8eT<E_#M2.\
&5O:L^Za9;+>_RDd=>T?dFf<^ADcOFM&02LT&^4T1=eQaKUH\DAMVS#@fU@EF^>+
,e=bRO<:[^eR>BF4NM^0aWT5Z7f)Q18dB9E(+b0]SIHBK<\RZedL@VN95Udc/#D1
F5++LV+/OdG3(dXc.O34(1B.&Y#)2^e+V]Y_eTX6@S]fU_g46T=e&3_;VTI,Xf;)
2>-aL7geY?R3d<=RNE_J-Fd=R?_?O6X;S;U7)YYF@f_?6N8_QBSRZ47#SOUSDa70
N0_5[d>OCRM32QNa_LZO\f^T#2af[Bce9JL:g^DOWX?dLgcaWAKT]JE1_HQC:Z]#
4FORReMVQ)&V8VGT:O<3Jf_E&N_IC+8/8S]^5X#\7#=-b0UfAI\<YTS,JCIDHBUX
FMX+UdO_\S^R/BbbAbbELZ<0=G[J39?PKJB.)LEGB35<Dg5_/V=Tg(1TBFE1I^-d
I2CTR@8/#A\I/S>F(1B@M()F@L&4QC?1[eBKN857A+TPJ;=UM-]e#?-7B[ZJ#[7d
gA<GL;cKKc,7V@LKPRb;W1:cD3X9:]cN3@Fcb?/F_G.dP[c3JQ\Q8_6>>bdXf?O5
RTZBAbY3O>K[9dX(dbKg+@X7LWN)78,?g2]AVR1RFG41K8@GU9EKg1>11U9SCA68
I9]CGOIdVLAGHY0K(0RD/PaR.8eHgT\C4g;8WFYg6)0B,X4+L+>:5^\SV.W5f8G(
8abaOYO3D,1_E(4ZU5-V^,aKP&)SYD1@/3E]d]H]f32=]DD3F(,@&cA@-H0CcUNZ
dE#<bKS\G1&\]P.F(6GIRc6HX77@;U720/WJ&0d05]Ze#L6Kd=6TU@Y#)A>A.23L
a4@W<(GX.C6_-S6>_9G>2bCN3^&aNIM]e-VBaB=JTcH0LdYE(EIG#)=8NYBga3BD
+X:PT.Ydcd=F<RBc0S0R7TATQS,48Z9@H5&[#+eA4]6g<7.^g6.BUSF+G)JAe,Ac
_;97eP,R<0.QgT,(.>bD.2E:1).3JKD&VM5,=PT+7\fX9(DK_W[QM-UYg\N=e9]_
Ic6d__/L@^@SB>:[;9\,?C@RCL6=E+cKE2CYCfXV/2ILB8>AaB+0cWZW\N726V>.
X/IX/D;:14dHaQFdA5BI,W?[2(E].<\)a3^WO8HZOeK221<.?@SAHB&6C5<_54L]
#D4F,P_\DIJ;]3bK3AP)[\b3MOM;7-VgA+eHBR^J4P)IK-_;.9R4KK_FGY(>-D34
CQB);2O@-c;fb1CK35F#BD09\9OBWYEH3;D,&Xg#eO\XT7&TNc>,@;eOBI>H0\,K
H3(4#XZS<;)N8F80T.Z9CGJ1?2^@>^ZAJ?S6e=QJO>PKb5G=L0[O[+R)L;7Ua3?O
GV[b\Y_<<f2XJS[aL(a&HG,ER:Y-E=SICH)H>X1]g.DUD[)?N^8:MYW./,BX^&&S
[Z>>Ie2d_:Sgb6?XOH/UNM[(6<Y8Y>\?2P&<9P#WAW_&MFG43N80?-FJU_Fd0KEI
WTZ+70H(=b]GPK69NFF1UC(^,;\:K1:-a,,ggIHUa[UFG0EfM=C[OOP;f73FeD2K
P,,b::PO>;g^97(;cY]UV+BYL_4]KQ?3+](BZ_=E,P:L.CdZdaU@=+:/NacLKge-
51)6GO58+^^R:WMO4#-\]b:O[J3Q0]CI&XHH3#N0:Y+Y0XBN>PIJ<)M/c@_EEC-9
Dg]UITMYNCFd<LDUgVXV(,]2c;>M2N[f:(Xg=>DQ428d:KRP4YH@I.MWJMLN5@CX
WcFYGFd[[fG0U,2UNQgYO-_+N[<N+\YNaeS.CQGV2>B<B(4[3,Y5ZS91])@)DI8=
X(Z,&c?Z.8JPeC4=E9-H?W;b)RI&S1#9WGD&3Q-X0bYcZG-)(fe,@Ya@</,/Q]Z1
3M4N0TgEV=PQSR]1S6=J[d_V>A_C^\6A]P?WK92KWKXfWLeCPJ,e\3(;T7@0D]T\
e,#D](ML+S([2#QS&X3->(KN,ePW?^A4<31-VDC511gI#0d#M3+9#4(0YS?E:9=.
1B(b5O.+LMM:b6;G2;QXc\5+5E-9Td/GdL&>ca?RI\J/gLURP0^#NTQ^6b,@ON2A
__[b\FNSHR=Z+H-CE[J-FZ\7G@VCP\BT\3VEU4=34,@<C+P?6F];53)?^#XFYJ7C
+R>;UKP&QdgdR@6S)fTM@0?41\CUc@\^\Z?SPFA(95H(QDY8e49RITYPEe@+(I7F
-FZ]OY:DH^4E9)D2<X[?gE_2CV#2HU@LP,MSYAIT07H[Q&JeJGGRZ^Z8T:gE]eLK
[dKGV/FCARUD6(Z]/N9+J^7>N^TY2FggVf8TA0R4.SF7/JXGJ5>MGSPVdIVP3Y)H
+UD,2C+]dG2(DbZ@N>1U3PY\AT:a4T,9#Tb<VQ:Z>43DeG0A1PbGcVd1<Keb7DJ/
)]Lc;_UdTbH:[b-JL[+:.SYJ8H.W(LGN]X_-0/GKP5P2d&VfN&QO7(1#Jed/A,gC
4B^YV/X,e4++TVZ.aId6T<^Ge-1VSbQC4RPE&]13BB_=+_e/#/TPfSXC\:-Xf]A,
f&bA/8N<8OFL-8B)^-\IM1WeDRM2PF;b&\HB9R6FZL8M1()VDaRb[444_Z^/EY<3
5SUK45KJL=)IU69K>\)MZI3N87T-^6#F-=()?-?A8#.<U,+6^NeMB?F97e7NeS>A
<E/cLFdf#/J0P;\0V3(H>SP[TD9KAKc[F&AFc9aU\CY^R&L:8eL1eR\MR](/@N+:
Y?03@^>^+<-XGfZ_edKG/dZM3U=-P6KU8EWO9@6[gM5>Q.T;.\S/_-PcV/91X@O(
][A(R+Q_G\]EN1+/0DEH#X+R1671^Fd,+EI<;3TgYMK0e7feUYD;B^gecKDU8,\0
-a<RZVb.eeY/aS:;J@)P4/J5V.cP_:a+aM,dSG;J\2L/b?SV=R<X<.bNZZ[)WEAF
;^]9]B>S1#XKKYH9_DBR,+\b;.;aZ@Y+NA\7F,[0-AG7V2I#c<UIN=[g&dXI6G4C
#>N#54Eg?2\)(IW5=?=T).1Q.Y=KY,d,gVU+&(O9IG?NEeMCI2BX:_5QfGI4XN^+
/6W&M4A>\g(JOCHMD,ef6#O[ISWEG65#4OD47WZ=a(.ZdQHU#R2W#?<b>TNSSe?>
JX[1?/YZN)6\3I].X25U/c2L3CKRCT(c^96F@e?bRFQ&Q6]G:BRacHC8=T@#_NL)
\#Z,\-R_]F:7\1A.-GA,QfQ<PX]f+YB:RXPa)2XSFf7=G^aD<2/AaF^7Y#.Z3JWH
S<@JY^YSVA;^M22@TP=32-61@KNY6,EFP:d2&TF2JH-PP5C^.MEYJ3E239(J5E@]
M^^H[Q)O6HU+Tc^,QI&JO@FCV?#Z94a>LfJd/E=IUD]G]cJ?+ZSWVEVV+I8P@HOO
5_]ZW9C^P)bNXDIe\D0c)OS>LV_Nc&>IN;>RK.U_BJ5Oa:?/3:@:L?:1[V)<#VQ+
5>[]?ad5C6MK9?N8U3JALZS>1H5\&8<=1]3V;++<a9I[YK1)[7]X?D3=5d?dUUEH
X8&F:ZcX9ZERWL-b>/dCFLC/[]I[1)#0QE8QKgef[7WC>d9d0<BS\f&C<RaZZMIf
KFXgV+L\dVG7eP>f^3V_B\(7X^S_::,K.X-V0Db5L&a^EK6O_Za7@-L2HQd;U_Pe
)^KaHf0_O(^b-B5SgaCOc</,[KI56G(/cQY.a>g2?gA9C.2VHF;b,b:JN@)W)0XB
^W40EMKY2Pc\6c4K/3TQTJI0fPgRH;:FAKQ)bM?)K\_,DeD1E1@SM5@HR91O?R<<
E&:0@Mc-8SLDJ1L<E;=cP5(^baLUQf@Kg;U(A>LW-JS4IYL7b[[_a<#F>>\:J<3X
91@bU0?g_T6M2Ac9(-8eb@P7=5X<HZdE[RETfYdJccX]-_Z#;ZAZZTQA7)fKGaM5
;-@TD6_V3OR)4Z#HW2a;Sf<^P&cA3NaH=>91/<Q?SYD,T<04Macg,5UWB\M\bDI\
BffcHEPP@Y:<C^O=B\d<]O\YG9X3IFPST2Z#a)B;a4dLN\C=4,Kg@9H=W\NT1V:5
X5\>MJYZJE=f1^Y^/7S(\;d89O@4&d7&.SLH?AT(#,_H9.NXdb_<Xg:&2U.W0R#f
YT://;KJ]GdX1S-?9T(78-CD4IU(<dBBAM3D_2=-I=AdA/]bHFA#_T-SBb[@:38+
W_HH\c]?0FSUMaD&0,/RXNO[W3I&<\WLR/g+1ZZ@EZ?S(b_X\?L3U=XKdW==<#H(
aF@DX48U:dg5&:Y5E5C=:^M]CUW@[K\:9c[<gYHBW0,9/)]&_2P,KEd)1fgH=1M(
bcgY+-eB<&0YR;5?RT7Mb;I)RS0NR)NL=0NM2I/3:71C[;E&N62b/5Ee8eH5M[7P
(=aJ^J^=ZBMWFT@@M0,+QW_.?L.648>?JDfEL(MgdZ^[a314cH1=ga@O[(e/FBdD
?W3KTP,_,_?Z6;TB9]DL[0U5=Yf)0:d#Hb(-5?g^=bDNL<,,\a2?&99[NA]8UYQ9
4b.&_=<UTe<3A.?:aNN449\MK1A9Y0VQ-Y:OKV_IU1DfaScG/7\^\DNfA&I@XMgW
gIX2?/LG14f.-Z2U&>f7U,MM\f.D^.MT=L7AU8;[8]6Vf+,U4fLdZN7)cNJOeX&G
#&E3)fIJfDU?SK+a1^b#d]ZE/-&[Wg^8.3K\U5M^?Pg/&J+9-fg]F^U^2?)UaKBF
0H/KGa5S)1U-ZGcT[2S2<0?I8(/[bOI1PY]Z8>^U>IcB^YRc+TS^F\PD^4T3W@M_
[4X/:TY6a01cfJ>S,f-ETG=LKAW@FVgJ>]QOc<MU&LX#_[1CK^0=MLU8=ADTCaYX
RC0:)L7>FS,+NQE)H_I<>BH1C]0E@1):FCY)O[B?b1Ucefd3O]=?O=^E4(,=eP@A
X&3gD_(&QRO^1[A-.1GR:-IWF/:.Tb3HIPJLg+^5Xc/GN(:&RfF[10f2dR5T5^Mc
TEV5(Zg?:3;+6]YB?,6b:Y_N^Z>-cQD+L>?7N[@P;]cd4GN^L,9IMb,Z5WJA0A[a
LEdHgDHV7<)J/327I2g;ZEOW^A.U8QdKe.-f]2M-[/?a51dXSGHTVb4dX[IM3+#J
#YfHEg0X07eTHec]=OCBPRa2U,LO?cQUCU8T-.):=C5Y29QB/d(fM3Z8)F#FSKDG
[3Fe-]XO9Mde/-9;R3YQ;Z<3DT3CMQ;GCaC#6X.(6\48a:efVA[X8d8?EO#5LGJ&
]OF<SCc]gcKH).\6I6DA_4eXHA:P0A-?)d#gR77)dA7,@=<Q0E)3/OUO+EKUJJWc
7Z_4_1gC9-90LT4KT7,@c28[gfG8eZDa9a19N7#1Jg<M?M[FH)IUUDJg>)+>]K[;
:IRSO0K8aX&.L/e0(E2T#.b_e;(b?A(YHA\HKGDaAJ54+8IZ=ZC0^K/JPGDLCAGc
IS1cM#Df)>0+N1]E6OH0O?1cg@=F#N2b.LA9LC90RJD7?d+O<L73c2D7AaLSF=JM
e/@]f^L7YH3ZYLRMD)GM@.TT3:2LHL:0_-=bOGVSbEH0[L(Oa213J,=eL4;HW#KZ
D&IO4=gR>9#b#IFR6?;XS7JP>&^N=(]<N.:)Da]/-4QF2\9Y]6&]EYBU8ZPWYOH=
\PD:cSPH54//P5111e&CYbXc/TDD2]aK(87XRH)?g_9=?eagaMe9,&9RWJAQ6WUc
(H:eUL/Ug^#0[^3#+KVFTa#(2DZ60c(,?gDfG[RKd5,Y7S+0f6Q.G6T1<)Q.D\;,
L.9\U(TZU+.B>+(_.)5BF+gP_&]3g7=ZY2I,D=<#dV3H(P0deUI8\.FgL,;DR2b2
V97@C0^@7=O-J)\<4+3(^FH,2G/RI[UWD2Z_a>79\fY3dH1Tf&,NI1QD&;7=c99J
WZ9:TbJUGPTUAEC:f2@[LgDG;#AY:T=B@YWZe]^f;PC&]8Z4@779[2_.V=cX.cca
0QG2BZPX3PBENS1S#ULWHcaOT/Z7eEeaX(J-.OYeA\7\MAAWI#7MK.dOY<AQF4<\
e=[K4U(POKB1Z&4LeHOca?88Fc)#A,2\9N/(dT/6W:B&S?G\PC9Y_;7OYfegf35c
R4-JAb?9ED5+;fH:5A,LIeQJJbIHLU#Y.F[(<3.XdZ(,:0)?-dI,=]GI+O(7YMBZ
#7ORB@-)Q>DH>K[GbX^2<:6d=R>>fIC<-\6BCUP3Z>G]&[+=Ee/A74<V6Z_aP<,R
@0=gGZV^YE2)DL6^(=gCbCLe7V-UCbME?8&@.@RPC[=Z].2<=?WAEYKPfVC4Q-Q:
Q<^Q;#9>2M=Hc1P88NHQN[S>bPZ^>:8]M/,.GSXg/H:92&?\_g<BXKCBE(LN5>W6
2-bA?V.C7)ZR#Q_/S+Q^X+31=.gAe-cRA+CV?ZMC5@F:GKaOXQIX]ceP&XeOV>3#
OO@J]H[ILOBa?H#FOZ)[VA2QL:@X4:\TVW(PdO&>9H4/4_gaV?&U1\9b)D6H3-gD
7fC+B)9d1.c[,VU6Z&&\HPS5ZCY_VL>]K/US1B#G3NZH?T.Y?_LeHVW9G<E^H&bd
5J_7I>J:-GJI/?a2_5:^>4BAPG[D_f9K40CY:G[>6e#G<Ga1L1Z\f9[],E,D0R+#
LcN+&<WO0,1[g?EAO3BQ1[)Vf)bKffg&,-+GL3K.H8<bEC&N8F&HARb]TZ#G6gY.
S1Q?[6OO33N/:1Y[ZI4EfacAGAd/56F1)7TI:?-2\UYE19G6=Y,Z[?A?C&?#.W<D
IT0?gH9F5090)K_9J>=5]ZY[bQ]ET)=(cB:TXb9[CJJM3PfFP9Y,:Q0c:<YZL9^[
.:1<]7.;7?VPg\WdUP4(BAHS/+93MY<TBX2OQTMU6FRaM[/VCA20N[,(>B2Bc1&Q
-I>91<7gg([[..?KSCU7;\3D9OM:)0d<>NZLfcaIIIJD-P2eJ^[]>3H\dSZd#&g^
KcCVGIMVCbIC^SUU,-(NP^^QSGMSMMPXL@cT\#[,CEH+?eXVcZ),Ag;.Z>3bfdgR
f\IaPJACH4#VDILNO/_8:d;S9gL6d?BN]1\Q#JT[]_H1cFL2]DS6\@gA5?PG#7[L
e:,eEaaU)gcKGJ9R+CQ.a7I@91SOcSQ-2bMF9+-Z\J)JI?UKH88]D43C#b8II^9J
I+_99E]7Ec]L(1?4=H#G)E6X,_&MB:2IEOXFY&(JAAD\EdE[Y1^/W/,R(/L;&5Y-
-51fI<<SV;KFG/ebC2P5B/:gUVC<<c5e.&#G>@YPNUVN,/CRE-d^:4WG]BP+RU81
ZefIG<(_6TRLB6\<@^bePc9NgBA-JJG0J@#9<B4f;/DcQg<IA=BMM[N]c,b5U=gP
-H8+R5eCY.(B+87-Yf<bP9ZR9cZ_1f,K]c->VK&3REPP=E,E]&/(U&W)-d/)_4B<
36:HU6&H#;[,:>Le1B40K8FaMUFB]2)dWKJ/73/\cRM4I6-W@UMXE.;bU^>M&2)U
OH]/,^R:D+SI5N+\)X\?M745_gT?J7fVf@=OJ=UJYb;,1&f[SfRK;+N9(N6#[^bA
-W6G@5VMZB-[2&_#A8f,Ff54/L=H1VP3ACgOFY8W+?\OMZaIbFKI^>7PQC?D_5JK
7TSZRQJ&\9\RGea)@?&>YG48bB9a=)=EHd+RP:F9aUQ#WGa+<3cDLBVY0=SRJ8+/
[gW+E>0K(PDC-Me@Q97[8PaS70>F&9G:Q-:DQEO>K@G<e>GI1M-=PKDX6M=WTQ>)
dc;I6AX5#?&Q-APUA4;dF:F7S/eRT[S<8@3C?,41^Ic4/dS@f5K0OJ#OKZ>f60E0
8BJ(eRR:P]ZfHfQS9#HPB_.7_FN_?HY8[28OWFJ2e5A/5]/3]<K\Q@YR5PAU69^7
57QG_O\e7[NJcPX^U=bK:@Y5R;TOAKHR]0P?V#@-<D4D<UHcYD_M;3A-7d\\,L=2
c=0<5UC;DN,XQOE^SE:fMI4T3bZGEUQ..VFX@Y,1O^1XC&1=[\O32,[/LS+:0R;\
3+[#C3HZd>2KH-/.IdQ1MbFKNHPR=1]A8D_P#<\NH/T987L=?AKB8)N8A5[Q.5;H
?6[03c/[<(Fd,K(VTZ8OaU8f]-<PBALBETY-U<D,0&&8@-L2#P2Fb.f1NGKE)0/-
4fa6IJ(6WbTU]gD3M2Hb7;H\_c.c)(:PNF5BK_U@,:HY:_)^>5#MK(G8S>5TXO^U
KU.VFU_^a+5]KdNSPFRT4;97?8I&?447a/JP0efd[SW[N-THZ7TQI+H_aFLPLNUT
[\/0=Z18@WGR3KRa8^P:2@CaD>F,c16E.?,-a25+4C58#40]?aSG?/#<O__KBcB2
K26SOOG[MYQXHUFM93C(J)_fW:VU71;5/VcSP1EcGeaXC/A0d:gg@cfUW3(9VF?3
UPe&1Q&.aX0^RdQ.NL[Sd,0X(,^/&Z4Ce]X\YgB#95GJEE^C8#c:DD[4?GVWMHa?
PJ&OR:Pa92;@[f;@&I&KHMRW\Z]BCbQ;HIZF/NFZ6_<:4^/YG=2f<G]DY7GHV.F5
64XRbQ3Yg,H&X<E#92@88+fcT>RIW<_4Bd1R53Mb]a5:R^SgDN]AN/Z1##G/3Z(1
+.OR)^)^24g=>\KHd7EWNJI6J-8-1]6Hb9SPJ;_C^/c@eS//(YbDQBI/YYe=+SA+
KK]^OK5LOJ#gG1WGK]EcO[6=Z.]1^884<GPfA&e09Y/H+AcRSEA_[O]@:J28/c5E
6RS\5FL#UJ/)^]2,@bSQ6P#/1;.AR;I0fTC4S;_b?;O.e1/CL--C7P6.ODJ7ZZPE
a6(#Z;,B(@fSIS;@WZYB_K?RYfa[&9O7Y:PYH&Y&]C/BDeT\(.\f=90S)JEBK<K]
_\dT#[#V:^&<\I.7^:VI>A7K&?7@eKMac:\@C^bZZeN+NR:fGX26BaJCcX-W?>A#
SCfH;+cP?fED+=]3IYY@4W8=F>Ka^RFXCK3.:O0AN1^LY+a-MN9NB1>7-d\&]4AE
&F@5Z#Z.\E+e;:-TD:1Q.E@/17.Dc6[?]0@@LIg-4:fRIY.KeXMGbGEH[8a6/4&/
86a>\5:J5DTIQ.J=XR_]4I6+TQXGLKKS@c08#W+H7dIdIF?f^L1GL<8I]#?23>;C
e>(&O<fcY-(@bM/Y8]0^d3Y1VKAV1AD=3X.65G<JL9^MO@G[6U.V-[7CJ<CAC;f:
V&?cD6]Y/1U8<R5D2EG^Z1.UM24M(:5+J8[JH&d8(_8ETaAPJJSIG+d,:83CgE,0
A9]]^@LH^.05\@[&b[S88^Q;9:/a6adX>;HD/-3B[XT2Df)3<b\0W;)0AU^9gW/[
@dW2DV6H_Q=55,eMB.?/c>5?]-QfMUgN02@A@J,]^KDYb_71-gW0]^:[7-FAJ:fV
&:=4[AROJbO.,P<>XC4/2Gc<VD9_H&3^^@^_&_PCKPfEK(Y1(84D78f]8R2K-7eG
LB:?)4H^(?)X0YB;&YUO#H:^X+C/BPQ(H#X,fMYMf0A7X@@e/HS(@R9WJ>^VKK7E
AL_9cI]V,T?#?;e&QTE-1&:ad&T2WdXKV^:<DdG3X+UB)S^7Ka?E+[3F1TGWe73O
/48S@4;JJc7f?ZARUBDRY#U8\D(O@]6[/PgPd+Rd)gD;K>/UW:8//F+01bPFA(8Q
H1LRB;_?]CQZB1TUVJdL&<9@&R1YK@d4\)-WgP,5E4VW[(UDWJODEPXIe-<1V&5M
K-8V33[ebZK9#;?.(E<5#PK;\HTNL1X<NPPA9EE+?RDC(O0\J1:Z<LMc1A5eIGe]
7[)1)&K@81KIBBXB>?6+(^V+F@XCB#WC;0HF_AW1#P7?VQ8[B5@.1EK+gF=GN2:C
&IQI8QT4.eIK?@2PS@UPeBfIY6M6VX^E@Td6HH&B@ccM)?[U-+4QWb0_e(4N8bAd
6;WY.),C;F#]AGG.2ZWO]K(@KXT[(DZb^EM&[NCa+C1#ZaBb+.Z2T_c;0:I-0P>Z
?/B6dYH1D>Q\=f#D9@)HVZc-8H>f00[YMN;9?80af:;RQI=;5@f17;;NFXOF)]9V
W<gG]dV](M,_F_-2>D6gLDcAG+B[QWGV&WCZ9PVM]8G^J0,[0Z(g1WWg)O:GD.b>
c::Y0d0ePYc0(AE,]J?VE7-FUO\LOE,_(>NU//>;N&N8R010WC)>Q\M-NGfQ:N;Q
Q0SM\<-XNFBOIcT.E#W53.+BSf;M6d,3#Y_bNV1N/G)/&2K=OW,V)Xd&1BCf6V+2
+2P23+62[=bR9Ng7QSR0Q^55XZWNS]X.#[JPB^F0QCg?f)W137aD@&N0X818[WZ)
XdG1K7WJSM92>@A2INRD8K1R<<O(-I+F)K50^TG94b4VHQ7AaYWFfOKA5VZH?&Q^
VFQ6+4<L0/[?0FgGGV_6)U@S3B>Pg04]OD[MFg6Xb=6Q5Q;#/e>E#VGfK82A;e)K
38DL[efI2d#ZX(cKT[?c996E+WUG@..(6GTf4<J@ceeI0fD[EUR++^0U]+I4E<Vg
ZZ)OUR5D@AT_)7K6/\87e@4D>a+>Xa,GDTGJTHGdD..<0D8TLDD;S9g@:efb.=^4
=4IB89EIY&G>=O=ZE/CV>ReG&7R0<0<V),)]65D=XY^LJOc;eFF+YQ1;fG>/Y40;
?1Ze6&S4Z88DaD-&9)1Ab_,0M#7R>^^ML#@_<c\Y\3bA+)<_-b7a0)bU21JJH5,<
A.J-=G4Q<N9Sc>?&:E?aTI<dNUZ<FXdTKP/;5L8XD-Y[F0QMJ/,B634O:>IH#[[C
D+D;]7[C@#_YH^cO2e,].X5GL5:91c1C;Y6a<IYMfS??E@.S?;CdYZIS;>1RNg[N
?-N9]A.1Id<dIWTW^<8D1V308B8aE?fa>e7C=PE[R;HR8/-;8XSZFM>62&#,][^;
,S+EE4(:7c;_H7KLY=8=J(M@E27<XgE0QDB5ac[>FY:B?1?7_bK9S(]H/dTbJ9&\
@(3M.X8TA<JP17^7OOP,\OA2:9eI-R#c=3M7CHZJ(Ub10.dDCeAHC^ANNSg+Y\M0
N-NQ#<0/(eEb2gB1^_a/G<2Eb)L<@LSf+a?B_&.-FEeB7(a6Q>L_2feDJ=[GU+\G
OMT+4d7CgOR=^BK0CO?+Oa0B?6e90LEU[7dL,;dLQ-:bdO9WcPQN2X:5M&K=D<SE
U^YAPNUcI3Z@9RW-:5IHS:B02PZ:3YfB7(Ng5_@eD;,+?A^b).#63I&bZ9:D770a
\I01P#J0@B0LYJT8HZZSG>Q[O#]6b0DF3URce0.\S_DBL5FD]Jf,8DD.AAZPG<+0
WLB8\dZb_BaQecM6e.548e1UK\I>M9B>6CM_1\4dZU9-9KH_G.-N,8J;@PcRKF5^
1aFYYA591Z-&[8,7=7VBNa]H2;6Vb>4P-PBda][cI0[DcZ,a/,.Bd@a5&;Pd5M:X
M>FD)R.URH8\g&^-9T#WO9=19_)5&2)2OMfgW5>U208YIeV1PB]S1XQ0=]Q;3Q=V
:PI.)VN:NKC].RD(&3.P2&Q\D04FUC=O,]C#=e>O80YRfeT(I/eM9&KW8c/.)WLI
GgK&#^3_/6M(/U.:eaI@X0[[F4:/IbcNY\5=LZ/PaG#QR:MN]ZUS-N/c(;<WV?86
7;He6)W8.eM&Tf3f_)e:WQ3dL3J+>R6#SBgL]N1B)VYGT<-\+T3&G]2)b?PF@A9R
<Lb7?c_-eP>#c43ZFJfM.P2HfB\A[9DB9JN92gF^BE2[;f+dLK]P4-,DI8_,ReY;
A/c@C&P=63FcTfOc+ff7+&77;T/f-D?3F(U+4FFSY31Z2fYE8g]2T.G1TNRF5NB6
I463b1I.V9VYS:<.N[:SI+R-4PLeIX_XT@#+9A+efg,-[:2;:6C9eY=ZHd4HE4B(
6#Pg_^#N6gWLZN>6;PTN4:9SXDD)T^)PG=^Ob0XIGH?E(b5Z)4d&(N;J?+:bXF]2
YVVQ6Re_DAg0(ZSc22:EZ@5#NS9?c[_K+=5DVA2K(F6/12?]<NOfE8EaH++IEcRM
9Wb71<R6KJ9)[?3a9L/RS;9:+OJ.V\8J#SM4^f3-dV6(\AY6cB7<2Y^MKKA2@.2&
:B17O\]LOYcCc1CS-B](.2Mg(&Nc2<B&Hc<1\QH;O&I#6J8[3G3#0:MddL>_B<ZO
DM]D-X/T\KSfP(Y?+G^G&8J&PW04T<FNP/bTJRCTV1&AL8@:ONH6Z<ba1/);<BCJ
DQ^W.ML+PQQa7GbT_e_TQ,9C>0Y/VDb1#@H_WJ&8XVAE&,@;6]Z6]4P0S;A=F3+P
CA(P.QRf<@V_HB=3P#6MT\6<gNP<I,[&&=PV3Q,I-[CI@2P.I+@K5(I=#a\W&cD2
WELC6_DVLd].;>5@67Q?MOP2.E?<^/O-05S]+@\5XN/\9[#d&5Z89./,6M^=b:/I
>T:5=G2_C[IfcOcDRHa<]B+A+?A81c/A-6c_eb_Y-=_QK6N87aRL@B]+?D1AdQDO
A1T+Y_DL6@<4)NM(-E;51Ta-C=JWFRC?DLNH<c2BRE0dP5c:YEUW1/e^&IHfWJ,P
_Z>=6&O]YgP:9G?^UH#5&_8Tdc4QBe[)M@+G3Ed]DA,6?bDQAUBBKOHHg_D0HIB;
CcbZMb>PBeB9]bcHC=DD66X8H\1)WM9<@A=-NQNT:-P:@0(,.[SXPVIb]95Q:LXR
JK,,V4e&(OM>YMNd(fDIfF>CY:HC&K?2]>X0Lf:M?DM>^0P)>RE6_>9=CS+c5?Ee
=<2SaX4XLI62gT.(d:LB]/:.NPYeRcI--Q6_eT1fbIT7DfE(7Y(+H?e@J[58M]\(
TI(QUN<;:)BP:IcE<5HcQC-#>K06SYN#9#LY]Jfe(KUNAa4X1W<TaR>K>>0O2dKf
2HJ]A\\bI8W[UMTXH&TgPT+G;]:N=S_SP@4C7aOcfNaNbT_gNK[&\MAU:NYfZY=<
,,a9Y>4Nf7-bQ6&Z?RI92+OT9I+T;N/0T3BI6ETeR<:=HK=3Cb(/c//d@;Y6=^f4
-EU:T4YU[.Ee9CY05^+D6).d3e?#=g:9eBE^J1W?<e0^&(39[/=1HQ_Yf-f=MV5g
=TWRF6HNgfW8F=9Egd_S3_?#MUH9LW/eA\?EeA5\[435e_Kb@Z+>gVEf8AH3&)R_
X;FHbRT=g40R.YfST&<9JJ:D,;QF1;6X17=F@gVM=]1WJ9GE)?ZD_RPK<M^:4\PQ
B:R0;,P2gX94fAF27T=e&c_>#OT4U/O1MFgADR,[=QLeEL;@YTgO99SNJ@JE?Ve3
L.R#J6V)RE(HX,Na,<4.a,_6?#7d:,adD475Y\AM@>E-e+J]3W^BFCGR?(Mf^<N+
0SgTdQ+>^?WP;gOWONe@.bd15<^^J7.NB:AdH/^eFIXGZ?B[Y0d)=UPST<1-6XPC
S/A:O44QK<O>2DSY7QEd+d<6SVcY;3R986fL1.9F[3.#JNa/MJSQ1-M-C,?(B8=b
X:U5V,ELfN1\MeF\.-75_a+7@[gaC+O67XX<U^P3K5EeV)e,5Ze@#d.^LL<a#TK8
PNI0e)PQD^aD@e^F?:]A#LgR0VT#X]0<UNZRLKVEE&K)57C&\bWKfMV)TIO2D0NO
)V#:(bS4X-&7\::2KCWA)11/F@S6=JO#Af#b;.\_JF7a3?VaGE4C>1)>d<=a-0<.
a/bQJ.c9J-3gYV3ET-f<6G#a@EOd?LJ/H;(>SfE#dS])\U0XNgT0\0];TNGNRNNa
OAJR<77PceBTcL3WHEHZNAX)M2EAdg6092RBLJfF?\81DV-);7UH\ZbLBg)5gQ+Y
]9<a118J(d@_3=(.@OW#GaOO2WA@CF?e0DPDU7R>O3Sa3O]Ig1d?EC0XP2+[RO[:
b8/c#ML&eK>3.=0]KR,+a8K#7IZGTMfFX#\0U;5R3,g-B:LZ9fE+Ef@AGdJZaU(7
>I[V<V[>/,:ee7H5AIcg8CO\CNERBWG9KF<BW[E[V1@F)&>?O^^IRN\SACH2g5_[
Zc62H?/2E0X.?]#f3B2)JFLSLaCTTOM>DXION;fQeU:S/POSfB3<4=+9:3C35O2I
;?2bL=]_N_<UU^-0CBcF;.gZ[Ye4H/0QQQ8CB>VS)\0_0L]bf5\<4L9:,.[8SdJ_
&ESH\)CLZBI>-?V+8fFP,NK.^=8KT>B&dXH+gKT0ea93)AUe?FG(=O-LD+:-E&)9
CdNG?fF-\9a4X7SWO,Hg7,+8J2T308HVSa3gU-W]GL_A-]V/f&bBNT^/9XbW\;WE
JL3_8U[0#2&;<5[<N2c;QT8(YX^B)ZR\Eg+e,=&9:RE5c<;7VOc8M@OOP/71J=c^
DJ]=B;@R+6#X89Y,[T5HO[T@Q,4H2FTZVVI.YF_c-Q,Y#F/7IU[I.S9]BJ<TP.:f
O9\]8@@((W323bMK26ZeIbPWR;R>^I5bP\IYdI[.Y<Lff)5ZVW8XgE86/T/]JM,_
3f87UHHX0J=U)5V(g)Ad7[a,MVeE#PLHYfbPGUK+ZA9c<N?44/OC=KBeCLGD/@We
Q;I-YT;Df=SI9@GRXR,_T\:U->.&67.=S52:^K66K@aZ\3@BBcAB+199A=<G+2Kd
>Y^6-4E(66-J9+U)YTZ61HA<(:UY.;4_CcDOU.9F86QI20>U&]ZM.)[f+I[4Peb,
XCA\[(5G),4YW)@EB1EJAE)7U1GUFU/,?=/Vd9KeOQ-INYaH(Y8]\Q1Z4?-W):dN
4,;eaZ&(J>2^?8LVX+JGb+S.39AGE/71TR>\,NSB->#);ZeX>+&^^+d3,f:URZ^@
bGQT,ZRFb.4W>3RY)5F;]>f<L1[ded4RNA)g2[.X4U:M,5(_0g@/(-=<[^0<@QK5
BKdT-_caX(_NP,?+HDEJ8_=Uea\X<4X#?MRJUA9_d0eUgFJ1U6^Rb^5^N7&\&H/W
Z8f+:a<JdT;963a^A232+]3TIb@g+ARdGYRS:Y.N#).AM3.A.HU@ea?)0YJ9,]G?
MYE0]WV<X:gZae\415(^B>cdMPNB/0=#?U[\ggUHH_HE#<BPQWU05BcCg3>7J1O)
^QNAd:PR1XO-f>]_g&4ML-C8;(6&4c4C@@W,5O<GH<8:7F^_NI:#H8IPJQE)e:W&
JNAG^35c_)6d/D3Zc+6M.X-Y.7@CXN9:R(0&W_5(^RFMEMPZVeHd#PKK&/G\b4TQ
g64X+[c:L[Yf7(b\H2KFU-?14UA,56#Q2adfQ1(#([S[C.,;[J\BDA)e/IZLPfQ=
XNZ<AMe;6RNV@gK<<]7dXZE(Xa4FW[BHX8(c:]\TV+V^R7Y_R=VeZeO+F^)&J6FM
E4#f(FV/[IVC=E;0d?T3B\f3Gc_F;^(T<6dE09038Z3Q&f.YeK=<;)>L,e@-JH?8
1ITK3_4,HAe#(BEK3K0E71[;K(a<<=6D)V#(-9@;e7G8UWE1TgfW5?^;HB2J<T(d
&.e<g2K6dDc)#SX3YKI+?d,@5DW)8>AcB4&BGP&W,.H:CT;HAUM]YIWU)9#]AWCd
dZC9RPCT+O(DU1dR&fA>eN5S_-b2dPW)dW&)5NM[KOaPbM>1R@5Z=-60/=QU,+L\
^+6R>>X^d[BSQU>eV&[F7>^<(OUccC:O-_L7/eR2W+Q>VJ#\LGI-CCDc-Z\M/Y3X
Z/;DIdD,Y4:Bg_A^IT,ZI&Mg\c(T\S1UELa5+>#CAY)caeH@DP]c\S)YZMXgP6fP
a]&,R0+_J6I-PZ#_\c.;HO_^2&U]gC5BSaD1JH96B\:a<fA?]Y2PY8^WLHHGH^O7
3K#,79:5^S^Af=M.ZWdMI_P\?3#JfMACR>G^_J6YS&S8D4K#4^W?EAKPaC=I.>e.
5+5EI16R4+))+\/\YIXN6c6S2GdI]7&N&H2:F4J_-S_8;W^H=bDX+YaA];TM2J5]
6QEf=g,IBO3_#10X\06]T)+M379)bGAI9YU_:8ZeJ<=E(8QT>L1;CE?3a]FD5XZT
#dY,9^N>0#>:F\>+O68dPTJN^EcXVVaV:F^&N+(XU3\[TbP)ea?^geX)@+)f>(2D
EfAeX.4J_+UWZ0bM.+4MJ2P7@LY5-b.OS5V[Q<De;bK?VMc\2?^CXV-Hf#BX=83d
(\B_#7KG3[C)@<ZF6af@LP)-VR-?5P=L+aT-+eWGL84D<G2;XJ+1XX.HNE]EG]E#
.;84K+^aJ;-XV)=g_&b).,4?KZEI+KQP4QI<Q+3J+/I:S[I:H&f:D+8d+G>1R:C^
bH.@P.S.&#37?g7ZA4SPR\Q0;K,\:#g<A9O\28/MZT8d\4@d>,/+O0>.=(AA2E[<
)a)c<eRQ3B<(gGg977:?YWTOI9Z4/ES4F5N63R-5IY9f]4>AF)2U02C=-4/bUYLA
JfcXC=W]U<\6&7S5RegMX]R&R7#d@HRJ#/RM2::?Re7Nf>RAW?UJV<8&f3J\Y\X?
&9JXRWCAZYaVg+3dWTWIc=4:>:b/)>H<R@L/>4Qd9cY=P#FT8PYeD^23UXX^bHCF
&DG4g7WS61Q(bd0HQKQW^@>JE-c)R^AbW4A_Gb=>/58eI;>4R)WCDK6K5IKLe+AL
G^Od.06(084T-bg_?X5?9>SV)B[Y0Y88K\+CWM:5c-9)5:J\&?H<,NOE1UU@2MP]
#13(,INE/H-NW-V2=FUP@TWJG2G,bW&1(R[VW2TB9(A7>_[g-Zf9O_e+9N@SV>VA
SRaY<0D91E-O8EZ[2:/,Ob7e4S\=0Tcc:.U^a_U5#?cN<b+b=;)MP:#G+O@OVDW_
^P=;1Y657:ARR#[0K4;;=<eO-KXdMS=]Ja.E,R\3\\gOAZ?4[2MXdcE\PE6=\0KW
\(]VaScAY/1V8ec#R2SJ5.&8fF]E^Q<Z&.3Le_,fKN7,bUAL;^F5,9L4K]g[7+d\
N4[[[DMGb_).R#]W4>=c11Fg2^NU,a)V4W--JB@3;)M=BF:]K?d1^+(N>.HS3[.6
CJeR+]Q74,I=Y?(:CbDG[6)T5<454f+d4<O#@-35P-TCI4SDfWO9);+FE94?Pe(=
6.6<DLUU8/0M>4^@O:5g#&K\:e3<5I)g<:Z=1#cQCS&9Q,69YN?N8+Q-I-a,L^g9
AFa[g5;IWO(O#@5RHZG:OBb9+RPX1T,JACG)DI8ZY1VHd.YE===7#U\Q5S>+/,JJ
gEB&J]\N^:P]S^T\a=@a84GZ6Y1EH_-AL9S,G#^Z,GfGbN6&[De]JGNBV@(I?TEM
(^LNHG8T2M3[@G(d\1H1>6-?D,0];OcO^]UUd=W:@HKX4+8a2HQZT\9/T-KRbA3Q
CAce68LB;N(+F74PcVJ53Jgg?&++&@+06RL]RX8XU/H)OINg?F()cTIcg?;[>[K,
@J[=e[7J;N9#Q+R,Q0VaeIb0M8#F+Y1C.OIY^BgSZO#<92_@D]^-C:e5X:.9)P&Z
@ddda(AeU.MI3VO0OdG8GN.A.-b=I,E0KSSG2d@ENZ4T6??W.1+XYJVELQIH83#d
9WOG?8R;#_O&e^ebe]>?ZHIER@/8Xd=W9HCS27KQ63gY];F94-4[X91]gdRNSeNb
.O,6WL9QFQ@N92K0PD^#8PI>HLBKBCf<OQC(Z1&DaU9AY=TF33cJ@C8BI+,,SJ/I
L/Y/e13_+?,+QXaF+GXVXPVYgQg=31D-)&.,U=X,K0ZH^9KEC^V09>JY^HH\FVEE
@(^X&_5fU(-W-EdQ0]e:H^W&5JAaOLUSZ\a5+;X^[#Rc^8=X<QPET?4?a?d9>U3D
;H(AYLG3M6JZb0I>[LE@3RLJAUZYHZgAgE(6dVE:/-X&CE-5KZ[&4V7/KZZ4cg#D
1MbLIDZ^;V9LH2[90EE=+Q)g>XH7?8,635[G-b)O:IT1KYM]a>SfL;(Z)-@YgBH9
X=Q<2ZZ^HM@>J]ZU?<CZ?#P1,4GA<REF6U[9;dX?TD=XWQ,H>OeaZgL6VC0&YQ[f
&BD?N>:4\:fWQ^,GJOa.A(LEI;eUf<gHe96CR1+71M08MLgF:<SL.2JC)QTbDA]Z
aeOXN2:&?;@/,MQd\G5g_&2a9UL;<TZ<24cR4a6=V_2-@(\Wf;ca/[XQaV197W@I
eH]CJ]+^Z=EI<<Ze(V4V4/1@aCg#=b5&1(>C1UO7/Z4a_)bKXH(5WY3C+WCC+/V2
SC(THK<&WA+_-+X26>gTRD7A>PGc;.+90B?LLB(0B1J_^_OC/-QS+/aQX7VZK8e\
F.&(0:T/C#OaaOgIBAWV9^,0#+M[-;>PL>[aCcA/c_<+,H7Y)Q@,\C/5\8f8^.b-
K@KUC,AN9Hf1]B;H-cSg\XALf3?Q)(D.TcCD7X(KW[g-Dc15MMS=XI3DA_da5:^[
c[0W]^3KS9eUX&.FbgM1P_>@9egSOC78>AZ17<O7F,R4BKdfZJAKH41Wa1-c(5_:
X>(6M=5V]>d,W95[Q<Le<?TYe-c#E=#U(G\Q7AVBKD32KBQfec#1,QFN82&XebBR
EDPEA?BQ)ZUGB)YDQGJZe+^fZcK#57U-;_^A):aKP4T9f_?ZQ4#X1f+KR@:9f+?S
]dX\KINO:8#3[Dd[J.LD15K;&b+d[.KO:/\e>J>)MI[P[0;;N8dg[3g3aU-J0[<,
-W)OLfRae<F92TPR:-<U^/GEVQ__a:VOb[)>c)ad]LG&FV2P5N&)^&4I85A9,KR2
WH@U/;ON+eeH=&E;3RXd+cN7E_93W78V7E^da<#Ab\5QA[G^[-ERb4WL->W>/7M;
821&E^#V?2+0325;PN)KYFc)+A7AN8^XX0?U1=#2-38,H71a3UA9O,XEX@E1M75M
9b_.VRAD#]bN/?1S=(^d0:-F7CBW-L,cd^OKaNEe<7+A&1F?19cbe4>\TSQ8:7>e
S;YN)3I8M=D&0@\Hc&L^D^8a(aA([+M[9Y.6NYE+aUHNYDJ#T3,^?),\+&4O8Ue=
V^&+(V+#3DA^:A+NQcW05D7AFFZ]g#YI)NWET@NEAT2d@4aEfD/?f28aKO)/4@a;
+9#,K5@-?MENDNY#/.eR4AR-FLW24/]MJ/Q&]2fO]N]8O0=0\,JCdT&9MR5-0g;0
/M-_>_Y1-[SO\.9ObJ#D0+4L.GC7C^[I3]2bJK^A\;a4<gUR85dee]5/5@?N1GO3
9;e+a4\W8Db8Qf+(b-K#)XcN6COF^g,GR?7-9_KeG7&_/e7?bP8ZCf(OP>(5b[gG
2/X2KQ5P.CW9;Z.>e9g4(.YaG4IT4dN;e_#K>BgbZ[BbZERF>.)GFF\\E(DDH3G)
H+OT7V]<L:#Y:;IJH7:AY79]M;X+gFD^P7=,eETM_]0GC(&A0?HBP[f\5R?K#(5U
c146AB2Ie6>0^A4SE2DM_J:8AS4&SN;.VQL]SWcbK18]WMg5RTS@KfD5W\,<9PA>
G_]HL#/3fd=&X:I._4XC3=bLODfMB4VD=P6+6S2VaOR3<d76.g3Be+OF\+O_1?R[
,CPb?UV[R;+GK6XG8BggVab15U<RJ9JJb7B?:;BLN)P1H439acXAeBPNC_BC/@P,
3[.#FdaEcQdP0@K8Aee2[]UQda;.#EGb^>O:P\H<JG=aTWPLYV#K[538gE6d5LXd
OMKSd;E?-;YgHIc^GK.a(./@OE:N(Df13+E:bHeO@QTBd+f1U)GW&[2QK<<RI/R&
M)62X.QL_F\9cM5@#.e[ZaGM)X<Dc/Y7@TeAAc[1a_g8^2F1d)?6G(OD.@^-B.;d
]<7SY:[af:c>cGgP.4f(Z+YJ]eS3C\R5[1KJ-71/Q84,[Y^)\B2aNB-,-bX[]YT]
:=Z:1UdgOB?:G4e@.UHD/?5I5@<5HTLQ;:]Le?F>];YFHU>@63cVC].<^f7:VXPG
0e,gP@eVRJ//f=<G68d#LLfQ.ea@FS=<d5#CD7cNcZ#\YED.TWXe;)JCNJA2(:4T
CSB5RB9SXbRL+KEd6eb^X,N+D/M>LJ-CG)EO&YA]Q]_UfP/J0XULeUNJ3+P2;DQb
KK<I[A^&R7.L782=EV>Q:.;]OKX2\CbB;C4?_U<Vb9N[R#5QZD6=MQ+:#[HZB.O]
cZD5CE6:.eTMDOgB;RO.>c,f1@b892X54W(4Y0:ddK-\e]NgOS/ZH=GX=O.>FH?Q
-+YEBSVSPNdLRCN98(g;ZL8.YSHQ=]7M@cW)6EF=@1C2P1fNE,b.LQ\0F=.(U,A]
R7,HDD@832BKd>90b6>_:NLFfB#ReIF>GQL0_?D1I+[5XARg2Dd>BbI9+gG/<^A.
SJW/MC?@&gHXOVEX/9_@[UR2TNE70#@LQDZ;2U_#eSYKWD[#GXLK42I5,VXM=0M:
NP/3G,OPR32XQb0+XTc2QfKRfVI?K_+4R6d-:?4/M<-C_Z0PFa\d[#G8AL)fR^9D
@/8&]La2fSL:5O.8Fgd9IOZSbfI2=<5G:LGK-aL</I)22<:?@HEC8UH]NS..KTZ>
MXMCW7UceXGQTYTR>BX;?6(:a^JdEEf1O=1:#O4D/W^2a(E7cWdZRZCU2cc64(eF
NDgS8Q,_F_)4&<::C<_BCTeM^#LRGF;B=Bg1g-EWPT8fOAXJG-H_c=]SY&WaZgN:
E<&/X:[<5+Z&<ae.^B-V8bK97??4_a8A3.SMA+4b[]L:6e\d>&bEIGFF/-.M5B&V
0SIAZcAD_D.N]&L<^)_UY>_d--:UH]MS<Z?>RHOfaNL1KDc1b,WV.(\WR;^LL@SL
Bb4c[b(M71XK&V>@LB#P;KBdKC+\P08\-6XV]=(VAP-FSaPCHO/#UBCY)8,UN&Q/
,Se4a>-3AYW:/^KYAA7&8W61D;Q3QQ@,eR9X1ND:EJTVcBS^MPf./&^9V#,M:7-f
5e4f#c:C;0DMY\ac[5KTU7Z_0:[c/e:Gag=KERad9^UUH[CBf36QE#7c3+cceVM2
7Jc(D?XJJHYe#P[^P[3+bFX^b>&D=V,EU)#X)<?NUI<BVTTg/SXHPSTEPBL(55;e
e<X(VX;KC[[)V-0RGG5>O-,@ASF(,^]O/\d=QO_<GSSV.OYEc+dc\(R[BW&IeXKW
^11.IS)E7YA=,(KK+JHWRTUGC^f;N(/Z4:;CK.0I5Kd#T=QXM2VKBTMUb8+X&NT+
cb2YB8T_7BD<P6]&R)UI]J[BO+4W(c3(7>AA[HR6MJ^Ic;e,17N/R6GQ3BXE&I0>
=cA@>L28(JD=KWVgWRW_a8X9U\:OVT>&G47R76>D4Qc]BR=4@/J_E_=LACUC-(/6
dOCe\)0aDOYTgHG:RTPd2CIG[=GG>PVPC+XNOU22K_Q;3LC,I>:,8M>:MV8OX]FB
gW97U(1(#5^Q5c4Z#8_McPLd?[85)b@AG0d;BW\9YWOd3P;c9Y4YOXe8YUB>GXI/
?+^NCJ:>WB]9H64X^BFX#]5Nd^XbK2)bX055N]bE[UXC?>gLR\,SHY.(O3]EMMQJ
15DU;Tc;\R==cH1Hd43Te]&f8QTb^^--cN:aXYCbLfMEY)g[>HGW)a3#<(V>E?a3
BNYDJX23Rb<<=#^-c;7K#,\b0dC#E8LGYa@GXP4.cMXGYNa#->f?QMW_/,Kd)_@O
1&<4KAL4HHT3&:+e>fZ9Vc7U;A1?/M,[\8b#:>N.[fC(V6AFcBT4#(RcSHMeX(83
OF#E>Q@CVL)>:B>J0W#+Sc9VK>9RWPVF#=GFJH6e(Ag:E;-4g99H[2D@f[Y7<e0K
9(M;XGS/)UXFZ[QKdFM6\:K];<=X_I>+<6R^@@DQM7AL@6,A&TXSg@EJ[^BSeK78
>Yc)>f4/3_eeW5_VLIM:7/8C8U&QXfe-PZAENCIKA\(.N/IK[UbD72Yf]BVI0+?b
2&2G4]K6f,580+FCb],;[fQ2bDO(P#?VU\H@Df-O(B=1g].-gQMaW[SB\F[SK-/+
9Jf;);UDBIWSJ>C(PHXRK^/4g[?^EOV[d,MPf[G-0g/_[Q#7P&e&>AWYc<A>L9/,
2Ng;bVOMUPSTaTLObG_0/<aIFcP_?GZVfEX?/B:93T^A@K)[EI&0_Vg/6@aP<4IM
A]+=K5GJ2L9O7QOF(9Kg[]CJWXdW56bLdb(]+5f[F^DKO>+_D2d=(cQZ<[\f-FXG
eccJW3fWe-e?LbDR2AX@9AS#S]U>Q@Hd]-Ke_G]I2Z3D@AJ(Z[6.ZT-=XINX+]Q8
3B6GVBgU5F?=f_2dI.>3dMUBH_)f[dK-&[&J8/d.T.a&\e\(L/4@WGb?YTX/Df;J
=>(,]F91TS.]LF&4,Gb,,GReUaF=O)c-cKcT6R_7R5PW2VG:RYFD@[#RVO]YVS&b
d]f<<8?YM/I6d:4?4K<6bRTQKgTDOH@A7O]O5?5UBAUO+=,^F;JG3B9XfKQ:Y>#V
3f6D&E?Refb8P\aeg#CKBDY]TTQU6QEH9#.]5?a^I.:C#QN)\dGTf/0:,=/9>TIe
HE+@U7ef4K,W<CA1#UDZNH\9BP<c-9TYY-Ce]6fPOQ9DJJ)38_P#Z4SQ5X9J59QI
OM=1c7g?]+6&Zae?(9f_BI@g]WNa:A,RKeIL@Z5(G>N@>-OX852d=c\H8U>LdeCU
UV#7MRA>QfB9]Q1;E:.AM.e[Ed5D6\B?ZFU^eY?R1Qc;)IH^;P6N_8&WaeMe0S/g
dNAdB@:(LH9g;Nf]<8(6fYP/6NE]U);0QLc__V3G>.)e5(3-P=(;+?a,J-cM6eNI
7,=?[g1H^>/<2^9/)f<)N;a<=&@I23:aBG[H,BT7fW0/8gHO:R;1</70cG.2.QT-
J/>R1;1d4YCVU-CJb3>1L_JV.B\=I1?_U<RPcPQ\2(@IUdGR222,@aNIN,QG[L):
/GX?f&6ZX;aGQg[>F2667J.W3&1YJaP@#EI>_=ATM@X^_=U)Ad=1D30#7&2M9FKE
ZGN>GaL>_0AM]8Vee]<N7,U1LL@K\6=S#g,LK=g422:IXF5GZYd&74&&GT38?I-0
6,4QGY:MU[2S#LP;]?+dPQd]E1,YP6]Xf_MOfXO6-XO:@<DeP>:9X_Kegf;^=.\e
b_cEB5Cg1NH,BHI#g\7X_#d0PH^MK,K+@eC[-6(?LFIS6<USVKg]d7^B(\C&:d??
^#R\/KK-H68I3]@:O5\<Ae;HIWV8FD;J8d6QJY2A06?TSE1(.FCAIQ=:C6e4/.\?
D/,IF/3ce,)80#&M78IZOZ-@LI2_c;TY[AX^Gebc?]L-];bFLV?)8a)2H3ZgR<M=
:40e5[BVSPOT2BO[1:05Fc0-E3QC,.1?C8B8c7^-(fN79E;UdWJ1ZJ3;8Da_63<P
6L_I:5^.;Tcf+]Y_#_S\?.S\+OS@F/c[358QdOgVM62;3R/WC[_H9:dO)-e\fQbO
=>Tc(Y+ac7N+eE?cW05?[RO+>_8K\HKeD2c3b>F1@BELGg=G,<c\HfLKUU&X0f]L
Z^)GS/IGKK^Z-ID<9-3:d_J:EGD3-BIgQU>/gDb)\P[8SaA#:\)U2[[AC&FX[ZUK
UU,D/LNcCI\+J#)c]GW)T2@U5N:QR(PSD_(b5_(8fGLM\8\^3.@50?e7(_^\S&KI
;A-H4:+P8_bYY:8ff[>e&>QfL>6):6OYf=;3EE?FF02&fS/15b&NN-Z6+N]]N=Sg
I2(TV=68(ccUPPb9TVM3eJ)aG,]NL7e^L2V2RI+TP9eGfV[H7?8BWHgKN(11?4f=
fOT-M&-UgX(eJG>^MM+.J<7#R(&\C_+O<R[JOSd32^4@6K)4P,V^@FQZ:Y,&X?DH
;9960HY0\@/IHeQ0/VZc,M+6@B@RY/SY8&2:FJC?SP1@?ZBaWL_H=A=0);;(=?E(
J8E+^^N]18Q#+1#2CNQg(A1c5:@e6YHV4B>AHXZEW.-IPbd7[:F__5]-1P#[Ag7_
&7\DH&.UG)b[fPQgK)f.>e_-7_[d]AIDbXP][IV7PK-NQ[LR;,#+\0Hd<eN3c4BH
a(;#//)EBESCQOB[de=\9UYR9DP<^?<(V._QS5L3VG//#<S)4CLWS)+J(@MU4EZI
3LK.>_/E-K/]b;RD6@3UEF&L[dBTT7g>K:[;1A#H,#^_0&UM#V4-BRK1e0N0,O./
N=b/G76G.Q,VIWgC@#=#KG04=X0U9A^LcP#9<;X.a_f578J)&A0]86-HcgcKa0g8
U(/RDbWZb3I7D[Q([6M.@&ZLLLNaLHTU4U<c67>H4Ld<5U:1eH4Xc:9YT&L38O^6
J^^Q0/=^L1>dA<c(L#Z(g5I0E+TRNE6_;DTS>93&5c<[HA\HJ3I,Y&BTUR#XE;(Q
THfXDRHI]QYZ<aFQ@0c).]6NV6<D(FYgPVMEC2-UBO3b7c4,)@(NM18UCI[G:f<d
bGPGd9V&VaG)JBYZ,geO,TJ-CF&0A+O0eTR^&WfGf>C#Og)5CSPKdbWPI@:?]87,
;/>-&-e]FaBQI68SQ-EG9T8bdIdG>FHD(^Ld>.?RWT<\cRW812EIX?XS?#>J)R2=
g+cSe7N2KA<,OH::e.P1>:FD<XS-N,94e#1]7-@]g[:&)GZFQaKS4L<b[MH)b/]K
bD/9[;0M:DKK<PXB]SD>R<eK-:BV#X(S?,b<10_LC50,O)XQBUDD9e;ZI6.],O+&
0WJK<B6C1e99:IX_a4BYU_AYH;TYfU#XF>@)@/OYLX>TC^(.JASf^#dLX0Y.I[:R
\0VV7e[5/bIA=\B/ZDC7N[)(C_;+NL?OP+_Yc,/;R@0-FGg#9)S4dL@NBYD?:=dI
1IWTD5XEe?_[+:ESK91F:TISUdZV/f5cA[:768Db+?4\:]LD6/+-??:7(2M:0-c,
?\LUW4;GfVRa@8K_H@W[H,[;6:Ge1N=?P:,.;8A(CU4R3f4=@>W];+W.<a-[^Z/O
8(O,93U8HY7#79-MP7-=4bG5>@#9O.fJ4F&?2IfV8=9J;H=H;5.\#393H,U5-2@\
JeT#9R)POe/#PdXX-RU?@7/VW9?eN_K^HIb-K5G[\+.eGZeO9G+9.:\?9ZcS4-?X
c/7NAKNB@6MXR+;C31P=_BD6[XZZSUC?Ig30fRd5ea?J9f:4GaJG#)g=bWJBH^;D
/IG[S(N6];.0]RL)_8@c3OfPW9+;C1ZTE\>+8?9Q3faFBdIZ\[YIf.:^MM&<Q_ZS
Obd@DaUVM,YF>G@N#DKPZe>]EWJZ9FJO4QW:f9>P5>;^=,/N59AD:.2@gKS)1dCD
NZ7@T2O/-ZG&IE=>Z91:]U,0[V[G4ISc&9]HNWZUgHaW\]_eWK<g:2G.;gVDVDQ,
C)HULZP-ZU8UFEBSe_+5Mb#3NZFc3bfMa4[EJadSg=G8ARKRf;\CM<81L0UMDJP2
^3718-C.;<f<C?.Qd:R,0S3/=2?\P3\@gA[bQbdO4V/4ZdVc[EWX@>_D\<d?8F4L
faeS:ZdAX@XH;.?1&_0IFY+&A7U;2Q9^gQM?Z1>FB,4^(Q-J8SEa.]B9RF=d-HG1
HXB?OZRZ]VVIZb[1UH0#,8+gE)5/]E85JG8ae>JA[b7FZ)S_>gZ[>SBbP(OL51J+
/d0aB0I/YYNWeMCHdYe[M1(.e\R2(,.f#SXC]#^SSCfY(UVc[_EJ3A.LEPK>G.f\
1LOZCOWf/P-d.Kd59-c4W#NJIYU,?0)0(HHVbEb=3O@Q7R^G^b5S7.@=-Ca#>DA7
MVEV:d5#,\=eVd8;gV+KYTL\WVAE98c0bCDc7N-a]DR:C;)-)NT2WUfQI0fW()A;
8U(4?;)U&4.UORDeG;c\YHZMXE^AL16>#\@a_4QNZ4&cacc1La9D0ba6IR:,7,1B
)C/_LD2E@cKGZHAT3f#g1[_3TJCYDA1TJ8\67D=@MW@&;QNG5ZN07dQMK,RbT+bc
f?5cC/]=\7b^K0<:Z@d79.F<6PQL=fM:[UC+BY3f<W]R1[)H/&gc6g;Q36g1;7YP
:5B-V,E-K3&]K)6\8:P2Eg?EeY.A&MFWGJ@)^-WC#Y0T@]c/)e:6UTDHc<?DGW4K
)cA?C@:&N2TBOUdg4=KZ7Z]D;Ea6H3HD)bJMZ8X>Zf_TJMd#52=VJcELU[bFBJ@f
.PgE:a^&KfUa<+DLJfA#RJ\gd.]HZ3\#:-^>MZQ/<ND-)RDEP1YZ9S;O40:A+\3G
3g0/WSY3\21\JE9^F47DV5ecJ-5LTQH8e)WdQU_bWB6X.d.2UR-JL@8UJSQYbfQ5
2_I:5XYJ5=MK<7,f-Q9P<@>IMTB98eM)\Q<NCW67]#6_XHOMP[=^-Sda=NDU\cLK
60I^\E>Y;3/VB&9<MTPI[9[IN<##S_=aEbN99bC.W@Q;=[EeOd.R32EPW(K;#)(K
I^be-]\7+A/#S&4Q,YdU)(7I6cPgdU+J?)3a^VV].Q-+<U0>\CW4VC;MXX4VGZ8H
;TT\V[T]5;=V#VGeQ=d66=dTU\Z[,f8@\;5>;MT(g^V_Mf:?-23+G>-gTe6J]NXH
KH@-BSY(H#>##V8TS1FHQ#Ce;@c7Z8ZLXBN&?8_)8fS<J]:CV1F/OU#B?S_ULMgK
[eK1)GQX(aP;?4/V[]H9<L,?=ZHKB23,+YY323KS=a:,fJ)GF^W&QbW,8EfCFc+b
J6eTg2P[b3<UM3NHSEU_2#bE67bKUS&/C8XH,b=9\9>+@[C)D?8OID#US))Lg(Nf
c+&9C[HUO>a)E@\]D/=1H[Q,94[VDfFV&G]KSII&a<A9LX51Re9WA[fd2(F#&EWb
Z6e:Q_^1]a=-B^D_=]>M?11B/DOc&f+.0c9J_U^A>94EM&-+=06+5T.WCD#O2YG/
^+)>CF-9-U3RJNQ)0+cefbgFECF-7V-&_UU&bJ=5G6=?PNL#Z>LEb/FG[..ZLe;/
\N(H2/9;2Mg5XKP00TUPBVdPKN7J64:>8<H#>;3.YK)<PAc.]#YMP08TUUG,2L8Y
,KdOfbKX^NbaE7]T203<E#5)B8;I<_/]-9.HgFO:L@;dYSPTgGGfU-PGCM1aRHfG
>+J@a6E)Ec[g(BfBRGUgE@bF:I9,MLc;Fg.O+Y,E@?N8-g^+5X#RTY#dCT^GJ4Aa
GQ#>TU]^L=XUMN>OT[d//RMT9]5)6[^=GgPUB[<UWDRYPMWM_V\4CN83[>&K?66e
&^L)IYdac0#@I>bC)/B&@UAP1KO\CE14==;fa(8QK=M9VXAG#f6a.0;:>bIgVXLL
Z\=6,HHIeA>JN?NIFg+:882231<dF=FMI7E:;9#^Le0@\^,933[NcV(/&C-&_M.7
:)/-a-)0I(323]X\T_CN+02SOX?Qb-&?a?2d#R7NC/SKMY,X11cWT#9^P=Z>L+3#
)\0H]]S>QLC)SO:(_AD.4M^3fI4Q#WFX?4g)f=7I;Se6UCYNfI@>4DCMOP5Pb=7/
F/UI+7>\F[6SG?W9:A7/Q_.8[0Y-5TT#MS\.P3d^V<\R&(<4GC):WZWWB-]C0C8P
d#g]Z(P,4C^G2,Kc\,VE1,J\SCc>G>5Ng7RI6(P6#?HG01efRMG,)R)aDZ-&99.5
2cE5K\Z<?Me#>+faD-F@[OP,_XVSAf\ALW+GO1.XK2eAT:C;&eD7Z3T60Z^_M)=d
(;U,38=eO6@]5\_/EXYc0:-J/-DNL(14Hb;PEQ#LB\NOVA^5.#KRG93QJ[H&B5F7
XfGe_LXN5E;gMfNTCLBUGRbbMYVeQJTX=2P8.aeOVJ[QS5OFY[g=EKHR2<FY3Ifg
Be\FHF0W[d2]BHC6P2B9XTJ>2c:W7L=8fW4\AK>Vb7->++X@2\NB;[E;4C0H9/P#
cf_R[[Ie.A#;+AXe5E/4)^/8<[G/Y_3QOY+(fI#V>g<X.RMBKR8dgBc5@EZ\&BF[
,.DY/(<>]X?VJ2_8:P7a\Z[,f7dKH\=2+Q:<A0_9D(,/J_?<6\]BM^AKTL7BJ4f1
6F2cbeW.V;[Sd1A3FG,YV79c8C4+ET1JKbSFYX8A2,\=d_HPc@.<G/)15&L]J;Lg
;gQ\EgFG,8c;LAJK#c=fY-(3,ecIJE_W^]>aC@aSHa7Q/X9TBZ@K8R=eMD<0=Pb0
LYb(bXPZY7g8?\5TZfc[-=a:PZV7RB_L&_&4S6EVQFJK[gKFDa[S-aM_cRH85>5_
BgA@f=Uc?+H,O7UW4O<I3_SM\FBH\95HF0&&TB2Jc1Z_6=UWNcOW9aeY+I0AM05Z
7?&0g+a30dQ:)cYTgG,<&BQcC9ZI_1MY,I2\:Z=Yf.aVY_?M(A,O2bCdREKYXHIa
DRM\,)^AT[fDT8d=6&7COcaCZM_.-Md(&BF481@E4JB=22WDKPX:cJHH1R-4]-f-
5OfI(3Z4670gKT?.XUZbE@f4UAI.7e)RR@ZIDgcIC]VHL[2(G,eHFY6L]RD5H^G-
V:3/:<9N7Q+Ode&>^=2C,9Cd]He>J9Me:=A2@4ZWKW3&PSON.Sfaf?[-@c#V<Y0)
b8D,,Qc84@XB8<CP9?TJR3dF0F4_-JfP#/:AdMD-2:O\(?P_W]7P-IPKDed@F-,E
87AS0-OQ(4J_OO+Sge47bSb\DFddgGIdK#DGg1g4B43/P:]35S-(d:-)K-MQ]O_;
5TQJ-f8:,?)I<bB=D\DKVDY4)ZN#_GCB^^5;.D)J=Iea\U5-W582bJ0Q8S:3M\)[
3=3eKe?BV5:ZV_T#cf2gfU^b/;@.KR9-PGPFBS;WWP@M[:F]?D<NQ+.RdfFLAQ<G
b36_0cNY4EEQBL_FC7[?J?dIBM3DB/JP-cN[1f,RA4Fd\LATO.7GLaTd-GUZ\5;L
W+Sa<I+AQT?QO8T]TH[Kb;4;;geI2&Ua\YgN-gB6G>D&\]T]cQ1?-ZgXQGaDBLX]
C@W.4d_;05NeVY^L=I=bA56<AO6E5(B_g#A#&9JUeMZ]V6?&5NYbA1?2\9-dcNQ3
6W)GR@@(IQ53HE\M6H0=/e0eJeHV_ef)>98U1RFc]6H+f,712E&fG74=Q?Q_K?((
8Z[UP&R#TDP.L,Y/aP&5Y05,NTe5gU80Y@]RZO0\+4eMIFQ-CLc/?K9VHRKOX9YK
YRE_]AfD2\J@S3b7&Dg<AO3Z;3aKg(b>Qg_;9e1#g(;:/WM^6D+9Fa_B)&>7IVgG
gM.XON[AF,:E8:Ha_JUBP6]LG^0a?L[8F3#XQX_aC,1YUZP&@PF]F,IPG)dXa[L=
#gf59SZccTb>#G54;ZAgKJG<NO98#K]EgP1@#H>[Q,3D5MZ8APU3>>CIGbL<_LW:
;UQ6ZeA27:81F>801E=PXcDbBP^:Q2RO:C:62;_8Z7a3I7[@1#/Lf_FDD_c=E./V
10ZccL0)GZ8([?61NTT<,dH>#SS.H8_.&HGeg.4H+.SgYGY;TaXCJ>,[Q5H8f)[&
F<QM+7>S>/-\(4?#]L<;-\9RR[Ie0c0B<AeK,:5B2O4WeZ&Q_?,DCAc.S&193=2=
#/g0B=:cZX6014a7=&&;c+eB#cR=K1;8\eR=ZNO9A;,57OcY(dbV]/PQI3:_TX?=
NU<8//4fO(6gRL4.&IUc>?gKe\F0ZLBQL0S,:g4b&_6\Q5ZPR@G3Yb#CHXHP[Kc+
JQ+5g^@3e/Xf#a>0N<B,@dP2Y@>?\\O<dY]..fVW,-c8:NKRB3;45_8e9JS?Z0LI
H-+Y1)E[?BBa5P@OcG4Ucf>bRFfK?9Ib0DC#AgI#[S_#:9-bbd62cUY92K7#N=T&
F)d7a4U/Z=2^fW#6US;=KL-b9FgPI4IE2S/>_]f4#330V?RY=<-a+J=,D=f5NI;^
9Q);9+]J>\TE)[<A>EK_TV[^ZC,Mb_2M5WORI2,gMOaQGQ(DTOZ03?3QVNEHS86;
W_G/TN/Q-\MFT;R8TcN8g?<H&fdF<D6V]LE[R1QLdX4a??_0-:&I:XG]<NM&2c@5
FeDL@CB]gUbeFaKgXVcPO+P7/0L=ZKET81.^&P9Ud\Z&QDHVB(ZSZPVeJF51:@GX
UbZ<9ZK+K5<2V2+gOX08b(D]TNKKDQLCcQJ;E8)b8A&F-QLFB)V?2X7EfX9T.CU[
MB[A2H6)M#:_[ACLM><Re1RJF)?S9Q7aK8+bW3EEbA-(.B-(1+7/&;#.>BQD9P0E
b8&=(W0N:]d>87bNPbe-6-OUcLe]OFcA<.J,>ENNNX-0GK(f2[DMY)DEK,d@#Eea
H@1?QN8=cSM5I2/Y)(,d64O<VNK-R[Pc(SW^D1DeG7DJ&beT3FKT6d=bG;EG(H)X
g1\?A55[M1>[E<gW=]3J96YRA5(>K/52ceMYc8,LTQ(F0g<OETR+(8MZeLJ+XMbR
\E5;H6/]EAg.\ERP=(a9=2P/a@,Kc-YTdPUW]D_;QaER>MHa5WK,+PfWaU/Wd,(H
&LUUJf0UEBDY>W8XJ24XG(2X:8#M8D,--e(M4T83[BFL1>]A/VgR)0HQf38LM,=H
IDL9^,d.18?d2.T;0]fMXO.A&0\\9;1):_7887<RMY_8)Zf/(J6b5SfB6Jd31e&G
\IOGC?C,4A&JWK]_A8RFF3.,6=M6055IKPID+X+/\&b\6==)/1W\PCT#<B+ScR>Z
,VRQaG.GOUBg:I2J9+1g5N+1S#[FIK/9&7.ccdP.^P:NcUP,a-ST1E3eUEMA6\b0
_<f(G/e=27-XUUK.E,UN7VBQNF#LGOXKNL#dGK^Pg+ED>)g>W2#b8=+WC:MaL:c6
_0>=Q1Zd+Pf9)[+S+R-bVCB[CCc1BZX&,Q9aV5S-WOQ3?R(9F>1^-#^YJgN(0KOc
SU6HYL=<PfNLacB7]0=W;[Va[][0))0//_e4E7ggg(+9P9I?TJc8e/_=V6/2@HZO
=U5_82)XS)\U35b0@@+ZcdRO-;KD6abR&0S=9>];-IUCGS;fA8:cZ0Q<V^,;H9Uc
\YU8a:+\R7,\Pc:DIC>C.<d;8N+2VZH,^M+,4M@.C#I1],K1N#_/fVYQ&HY4=].D
b7^7g+7HAe<Wb)^SDe:TBX?.3?\fMbg)c#Ca,#fLdAA^V3UNggD/RUS;=RS0f19?
IGPXa7cU0g<=[\XP[[;MT\HPA^bFaIXG5]R7cBdM<5+<2P>-]:^.f>?WR(gL-5IG
FM3b#<(d]CZN.,5C>O<eZ3;:QU_=G-CC_MV\G^\aXSI?UdV=-K.f-+>IV6O(L</9
I5NDI\\e:+.bV0.(?A3:2@aH@CD^MHXMR,3fQc-fGA@eG2gAdd:4_-&?>-gD<d@U
+0QA:gAMFDaAL2,.N^8<7;9?bN:30b@CC)Q>eZ3_OPG+(Xd7cN=>;_>LI@7aK#AJ
JAdT:=HC>a,cR0+C792MO[^aH?+G2O0.QKd]92a:S[C.f6aPJ.+?PbMVaZD@72CT
+2b)A1&D3RNW6@bN_(:0@D#c-b;_Z5F,g0O637Uc[FOU^[0[bgT@U)FB,91.c_#&
#^OZ?SL]Kg)&fdO=f&KVK/5QLO1N&JWSN8IA>##GWFIO4/Y#,UR59F5ZS3)66e6c
O]V8->^+COZRWB(LCGO=9KcS1-=d60&W+V#NS)2F1)LV9OUF-Y@6+XF\gcKWMIL<
D<fZY@\MQbV)[gf;(MM4J;;RW1VU8Ca(?1M/OJ3AME^IKI549ZS0MF7DdYWT@gBa
KUYa[P^F:^O1K1FNU19\HWDKZ)Ad85/LLVMWf&BF\=)4/7ZR[FQ1Da0Y.6>7>SB#
H&e]<M_2B5#\HRV:Q3?0g9JSD86P>NP>\/IJd-]7^,ATMYJ\^BI:M:[_/ON[@4)O
:LKdHO[fC@#CDFG/2+D@3bRGN189URTLC@)IP@W:I3.+Z3#W4FV)\RT7cM>L0\f+
6X<>2^D6_be26Q/B+FKdX3Y3/F3\R,fG<Vf0bC?R7MV/+a>G-B^-N\9_VQ;72C?=
0EE&N>_ga.a\81gAGX<9M3[7IOd3/T]#KU/E)4]fc2e[,=Vf71fFNUOTSERfZD)P
B[A07dca+X@)+:/VJUJ<Df:-H62X8gN(d?2E)0(gL?+5]X9J]:U_9eC0\KU+LB8Y
T=d^&)5#&I3NHJ12J57>=WJAI.NfI]MBVIR4?E?];&KLC3TSTJ]8BIBL\;34C6]E
C]M<_JG)@S#<-dcc[6^-8#6Qab@R7J1OOg1#TGHU48G-@bQC6Mad30;fC,M2+CFX
&Y5.L02I7PYM0@I5P<aU8&RR\gQ,MTN?=O>2Q9OAL2FQPcbPQM^@#HSVYKV<a\g#
O1<LRJc=EBgGUSXM/Y.(]>,C<>FOb5Q5e9_Ua_6-)H76/H9?:I405?:dTALZf&eW
[Z?Za#&&J108ec2T8YUF]T[A&=5S2M?U0I]<Ac?-UEY?JV.>ZN(<O9#^2ZC\+DI\
DMKT3BV@)(NO(A>Z9A)-OO7S1Z<I?4#K/,Q;LaG4N5XL0+SAC/@a/JK@YV9AK=cg
KUR@=7NU/eNJ)@=\gQIXAZ<U(0)<K=71F7_a&WZ4V7YY-P&+/c]P7Vf&-E<JC8<0
8b+58Q]=dIFKGJ_Gd#d0gA27#S&=@49f6H))XIH=)PCY?V/GU)#5K\QPa9F9,[GM
a9FPA0cgg3e;Y^7Z(f-@7aTQV&gV-[]]0e(HD\\BX][fP<\MN.&9eIbI]R]V-/\0
E00QMHcM&V2Hc4fd+YO:P\Ec7=KUf#cC#AccH9Y@.GW1g.bH=[VP>7/@>BL,bJG8
YFXV5RZO09)#Ue)J:b7e_2A3c,^7)Ub5DLF9;3_(8OK<A+?L?^T4?Ib[V@]OT/ZG
R[X(GK4VPN+.Ec;F8_f1eEUT/L8a@eU1f)90C/=CL-]&G4cQJR7K:0N#.;K]>9WX
4H3[CJ[)aNa?69eTHN;<[^]e2aKJ;=d=^H3X=:?7<]a\?:>\OG<Z0PQC^0RD.d\=
^I:d:80E0)UB0X1<LH^?5AQ6cVH,aAe.RPR0]E/8K[^f3E;B[;5<;]],?b4b/Xf+
;>2[1K2;4FM);W9#[dSD#8B3Y16-]@WA198S[7(QJV?eE3C<0#_#Mc6D+T:ad#6U
&R)CG6@Y=:2be\K)W1C1W+7\B@gAURK7N=.ZgP#<TRI(09O,6>7LZ@ZEF5-QRSbb
.GE;W+H^cI5EJ/VRdTa;AU:2[7_L=F_CL(MSBY6:><9O2U5;()><XGfbWL=2(A6P
BLHS4W]6_?g#bL;]@&ZNI8aCY9G^L7P/)409RX<_&C;0P33?:L[Kbd/;H[KA3Y@1
4ON6KX[X;XdFJ\TXe=FX=VM,+X1S50Q)C+-X[\DR5^86(.E,]]bFV,KN^3=LJe7-
23R[LQ5fHRPbO\8:>EVP^P;<AT-X;^(>6FK#<Y7CVNgR6<F=H[1B-Ab)R4;g]fOR
]TFTAGD+2[2ILZf1G<A,V-BfD_&UX9SU5D#3.3AD216QK[ecU.(V:#@DQ7.;Ga=;
V<4-:?Ff,<7,1Z&\AcG?eX6,TZW.L(g9+M+>M46^gZbQ6K8&-P0YgRSc=4+AMO.)
0:\U?M7X^8Y+;c(E5;,eJ^.Q:#cfU4R123Z_7EgAM]>Y^307J=LMMSRBR<KAMW[;
1@:98U[WSa&GG?Q,G3TT)9FF>6e3.a<]?8:^=9MGOX0ZPHaUU.4=&dQV^722G6##
aL7+7EBRQ5?#6&Yg&D6UAdYgEc-O1+Rb>cD0W-ZN:N<572gBRS8+HLVHTFE?WYQa
\MV1[cU7\2a&P;)d9BOAVLN7/e?=P&fNBNL5>0]7]R^O[JHY2f/V7LL#IF,&O1D>
QW5BS8<B,eFe9T2.V?ZEM97OG\:D#U2;Q\)JJ:=VcQOHFfbX@FNA@_C\P;[cQM=d
P^.K.T-2Z12,EZNDLQ>8L)1Y<P6TFS43TeZ]K\=KZ[/1SJFOePa5WKY1K8A0(WC^
+dF<B6)fVW\.LJO/GJ_)]6fG2<W<M0e9-<H0:.8[KYFeH;X?^S\M0&G4g]g/Q8?D
(>3>W_?EUY5.9A<BcTBHGY?&T6+91PU]AENa)YS7RWW?&XZJPCHfb#=(?38YbeRg
a_UFMf,Mf7gY1RRVgB.5QJZQNOT/F[#QS..<F9AL7I6bDMH7bL_.2@5^EEd<X-,[
]JbXY)4X4IWQ,VQ>fV2.&6-f\PCJN68Ofdg3.8A.YPP/+[N&:31PS\V4TcGBK:XH
=:/J0=2^MLgN_.?X&<;RDQX,R[#2EEO7BX>IA-Cb=I.U,fIXR?Wg_NG[Q=NZ(0A:
ef3KYCA,X+ea&A@4<)=\+-ZJYH#d,O5=L/C>L\,K0ZB)H?#;SFeC_^1;D[T+YZA1
/fL]S5^YTKGaW:L<^VF&OFc]+#_A60(\,S+I/:<2]c#B@K6-Z2?6WgHaG_B)GQ9A
I>fc@@0\Ef>,YaNVXaERLG?P_eXQ,e\GTAGC/CB(-ZCI?Z,:=5@XbD9SN[WbJ,)B
6Nff4F6M-.ZG&=BEQMF<Z&beE[_^<EJ:S+Y;:=/0)>ggII(NcJ,UQLfQGS>d)TR)
W&,&^H[L)/[Yf&GZa2MQNZEWLN)5C@2RFQVXM6Q\FKPZ(<WdE]ZU8@GIg6JeT4Y]
=\YJB1KT](-K5Q6J2aa^>/XZ4eI=B&1QCY]Db?(\YKSaDNUMY[U/N_T?)0c[B-.[
Yg<+KU0PGJR_KC:E9178OE7BU:+[\N?0?UQ[;8)g]3V[0aY8@FaW,G3<J6fFGU/&
,F7<c)gD^5KV:V+K]QaO-UF,WII_HZ[^N-afSO^1EEWVUZ7RE[-/cMHLROV_FBX\
=&B2_0P3CfM7e\2#CBfY]g,Y<G<WfHC?ccSW,.<[f8&6EDC1MOVdFX;TgY1[THEJ
U#;S(,G<d@HfeKU8-Y],9ALc::)AfNNV-f1c=2bO=_E_S7&]aUKYRL?&16d?X_H,
\9Q9-B][Z1\([_^>+;WOF+_@XKf/+VL_fUC5L/;G1[;<7H01#Ca0^.-NRBE#:LH0
+f@2f,V8_bJ=U172&IWfb<dL(WTP(T(Da>;.df_EU]O^^\4P/;+S6Cg7&+-+0\(V
P)UYRN)OLA@MF6)J(H#c6b(e8=^U^,gK&)Z15>Z/T)F5O4XC01MW1YR:<[G-1#=)
HGFC>DOcY)5@>MV:]N6MAAZX6AgBHga-;:?WBGQE\KJRIdb^T=4WFG^&E[J.e@3<
?f6NaN2N?)G-M]fTgN),B/fFG[;+BLUC17eZ7]5R.Eg2caB]FRZ&8Z<@KSCKJ?25
C9_c7S]AS1&5ZR^a,G_3_?V<VTG+?-Z)]5@b&\I&XA-=de0]PHde@Q44_)D^;A2I
KEQ+5:bX,aBF(=5)3LQ<A-44ga1CEQA=:7F&>\4@2<SW<@_>3?aAFf08?TS7U#f(
FL#.5]3AM-2He>M6Q[B4\:HS>Hb>7#3\,.2HG8=4[b0&f.ZK]S>(2?L/Fd681M)e
.ZD:T7:#,Gc6@2I<\^)&#Nd6Q:#DVQ@G9c<Ib(]<>C6;>JVD7J&6dXLb/PLa0,(d
[&IHCHYR=^3Rb,[8?X\0#V?P8(#f-:CbfTa.C(E/ZHYRM/]3S+3?BRA##K5d4I+O
g=67ZI+81PPV]JN2:/(c@=?\8S5.8?7>Y68Me7;V\4FeUMYBg_SaU-b.0&LU_6F\
_+[0(?P?dTV&<WD4O>+=fB57_+P:aHZ3fEgCK&E:R8/94d?B,?=NG0_2C/5@fS&a
JG8cdbSS&O]UdEF[1f?@=d1X\f>0dgAL8bOA4=@D1:KAM-Yc/#@HO1fZ>X;6Ab:_
7?@#(>Q1e\VSC;?R,I7B]Y]E<\Ea\&BSaA<O&QW#&a0AYEXU6/=.e#]7X[(0L-?P
b&158_GaCOY8a2UD#(aUZfRQCg9S=YHSCHbDAa(YMSfIDIHeB\Z<:(XJ3T8R(D&_
8TM8gG]eP4;0;KIT(^A=;4S[)C>aXbY\6Z=QW\(1MaKHgZ514O^\>[:BKeY^//Zf
,I96,O10KLKG/5WN;TJ1FG>Y>MS1LO,DdMW_[\W:3eMP55<I]84[_H>/^1B_^Y>D
.gfUH:PMUJ=9ZLd;QNSA)0]R7EZ4734,2S]:II]fI.C&f<bbH]M>8V<cdXee,M&F
)#_FA_e14HFO]DX=E9(CD3J.-7W,5]]C/4N,FOO[;;\C763F]beGGM>F5VZ<_-))
?bf&Lb[]M#&T;d;gYU-&0ObP:_IZ;&_[Hb_Ag-PPM(062UA,Z(+;?MHUg)GTPISc
4R(LUJ_626De?QFDb:cI+IL05;92S.AI65bCI4bI2gY&Med7X6g-94Y@&@>7bJ,,
gCI0XS8+/-N0/D?@K9I-(Nb[=HM4[b4fc,1]0GY4F+V/W.;S[#MT,QY-gg/ZWa:)
PaDR=^JFED4+G:d3PXgW>L#9K&0a,7=S3C#7d=.D(\6;7TJUX_G5&NC(.c,LY[/_
P#?Yd4bQR>N<gJd\HFCHL:0]a?^E(+YLgV@->8TM=^7-gbZAf-\TOIHE<@cY>.O<
.Q>+0UDb))D=e>5ZX?)(I07/80D3Be_82U0dWI3@D:(P;V8JC/-7adY]ReWb@7Eg
S?.g5Ibb9BFV+2D[0ED4Y\#,S@7=]dQ6e(1-O..SV0B50DQA[/U/5_A<fgI?9P/W
Dba3N6Vd7F-+6=2R\eOUU153IH:\gG8Z=0Le81dQ<NS5K]H4eG>2D;8:RNOfXTML
:>10VgWKfZb&,:W#aJ\AHPJ=HT_bX=a,O/I?fLZc-&+O[RSN[NDX01Z_9G8;Q9]b
5<5(&LgPCb9O6O-7QTS[/IcO4HDQ9.[2O@TM\;>@GgbR>J-RPI5YG4WN\KTA<@L0
N&C0dDIMe+E9W0+?KV=TVN?a:-^[E#<0&^Q_Q#a3K,)ddYU-UX42f[b?bW/31EXI
=ZLZe3>2Z;aMX:f_EF1#b9:bg3X[J?ce88XY5KfWLdgETHXU^TGa69PK3bg-=aQ&
\f9?LAV<]e8(<>#T7OA/cM^J\G=KD:L&HB9EG:Wb:18BaWAC4^LP#R0\H@F(;I/W
8d7QQ_:E;RK[e.f_^UM^W;K46@R.)KfSEPKG^UBK\_O#9+.BE]aO-0+IWSc?Yb#\
a&a7f^W(\9V6;SL-.>SC]Y]ZRIL.E_SAJ/8IdARHR\IR[&M,KTVG[[^+SM0@6T+6
7,HU9U3S[SgRd]DL15X-46ReQH+]CUI=LNK#B)G^AL_\Y0UNde9C7]6aCALY@K(D
X_\2#GVMPE3\0/.b-@4.[f#Z(&OS-E7K9WV4VGX9X3ZH0;45#cUHc,(MbAO7e1;B
J?cI=a,IIbA?J-A]I:MN7N3UAHZf7TbIcYB\^NgDJ/XQHCX-@P\DSfN@Z_7+O;8N
=X07bL\ABd39K]\a<L#WLL,?8Y3e4e19\[N(NG1UA/?EM]9N1\T6c9N2-<5XTaI)
aVY=ZV5K;1gFQD6dc,6&)?.B>-)7I-]JMcQ2?Eb;-[:U3GX8TF<:ZL9(7TI41//\
&(0U=D44QA?B\E<A#RJfUHZ@B+?eM59a&(eKf-J4-6@LRA^;@18_O/:SP\&\TDD\
88[)]aC&+b\+F0\>2<>NdcYBNH&1T.#A3eZWY.[T/SK3/2TM3>EV]D+M-C=ZCKAN
.;7=QH0Q13O;e[.cG#fCfS?788D)@g1eV>/RHf3@=3:48\6gaCHU5EF0U&J=,O/P
:c7\A,PT&J@@69<7-:CS191cP<K;D^).2cHI+7XaFa]55@]9@>TJV4V#2IXSBN_X
@1]O@#EEg[3^I1,R@XE,[S#We[E&>6J7.)<N)9bMNg&&^PIRaS:RBIg_&ff[@)RD
T)dGb-_Q:Z_\,W\-CaY\#(JG#5:=@3/8S4O7F:N-MEXc^JG9)4BYaVU(84V:#135
6&_Y:OY(g==I;EE[)0EVYTHP)\6W)D2e4]AD-:FTE8bKAL#Y=31?f?.Wb\)-@EQW
H]a[J.YVgI]=/5L>?8Nb;_)ZL0G,&g?b<]O&BO^U=aXXUNXRK15):<>=HgR:)4D1
OOB_E/(=Pb<aV-O<RB@?4LT0+?3HgEJ<XfF-[_O73XH>A:A(^YY-FFGK&#8d;B=9
gE1=3>aGX.TO/=140CaT.@+L42&_@\WPUaY\;.Le<X-IDP:I9@F18CM;V9WfRQT2
O/b0P^IZ9V0W4<CVWSAJW9QTW[S5=5.2Y/5c>AK)2(L65OAJN39S1?3&YMK-2,^:
8df::;>gM)[d<IB9\6YFc0W-K-U:g7<]F@Xc/abU/^F:N]@4M8DT,?dYcfR+W9;&
I_@MQ4b9F&-WN0F00T-KHF+Q0JBNUcIZR1N0>c8\ZL_<P1H^0EeQQFd8CE@BYc,&
JDMXV=ZK]EOP9^/,FVB>3D/GLUKMdDJaX6U\(J7g2F(cega#M_(Oe(_=_:?+7EH[
TL-B>=HL4V?+6EYcK=G+)=ZFe1I#cZ2#]d(/BSa:M)2;J>#WcMV]7b^:Z-bR8B):
5a(?S/D7GL3(W5DMR,<JgL0CP)#J10Z-WO?N[[WUBfbC;5gXcTB1O1#d.(#9\993
\?53H;>2,f.f]/#V0GgX^J70d;WQ53f\GM+Qb7?cI5+,C.;IM=0TA]Q@^VL+R\U?
K]XYUf(=E3>34Yb3Gg?/?=,/4>[D:_9W<]C,g])>/1M;dfFAF^74ZEa?X=T:TN74
])6Ue:+RKV[;31OKM\MMRFX)_Z@6XOJ1A=?E&>SfA.O-Sd[1<+O#CZa[NDV#3;Lg
W-H[U,8ZKScRFNKIEK3Jf)@QQ6;CP1DKE/B]fE,:R1PfI.fZM@gIf)8P9a3_:_V^
=.M.<^((#]P<-3Ba;C9N5J1GOe&U&gJ.LAC8S#B,(7TPX^de1=XaN#G_KU[^V/.]
&:QV3b,M=J]QUSKNFES6.BdV>:6cIOINV0XePZF_T@feA5PO=CE6?O0F281\bR51
&XBgM1IT980;VTLP?#]Lc^E:S<=L@X09E3N=@/;0>,V;70,<H#@S+.5^O:c&aWP_
6@2^K=^[48&36P-<BX]6S16^0/K#&F-#D#4c>3[MdE@V()MZA+M<G?[He?DU+IdO
9A3)J]K_@=T]D_<5GKdAY3:#KEdR-O4KY<TXR-^E9/14MPTX_&S84d-X]/1b7DR[
.[DeK8SSNXc:WKA(F^(=QX-MTSJ@7BGg4B_RNHE#c[VM5W<_JAG<T5M#-P57(UD\
/a=Xb2KLG9HX\.cgCXdMT>Adg+,BIP13^bI\ca8g#[CD54XM3WEPM>(@@Q39_&I)
J2OBE;[YP2d&/)R/b\PgdeD0[d0+L+B&XbY<-_W]?W,,R7>Hd9\BF/9NMG<MS7U7
2PR2,T^(W]/aVH_OI1\QY\&]FCSaIU>F>#>_;6gP4[Z208IcXcY)FFPa\SS(R879
<S0#dX(#R_495UEXH@CQJOQ)^)aF&,6.+\JT^T^PL:SF^JdcP08eR<VNgR6YQU5E
2Id)&Q7d7>?WDUGKfBV<F[5]B@fEdcgc\YV._LHYYHT)]&LGgd#ZG2_a#F,.15AW
fe/B4VZNL6Y<c79G)@4CV51050f/]4/8&1O9Q#7eOJZ)-D)+AFLg23/5>]EeON,L
J)I5gZG5]+cP\A:4>TI:43(dN3QX,/35JBWgTf_.+C1XGg:#;4Jb7FI6NX8Ae^&B
MG_?MfdB?:#4EMdC,#LQ8M5dXdYdHGdO8X+Fb8^gg0DCRFbD^Vag2LGUa.+fgW/X
)H6OBS1CK4[:Rb(:P)JdC?1&IRKYSF?S3QPR8UXUL?@L+-JYPd+FM5O8DQcU;WF9
WRQQINb\R]W.X4X96Q3Y4)]K(9P=ELG0_]FINI,/eH1?\@LHY:O-SF2-/<Qf1DP6
M,g7B&aFXUQ;UK,DMIR,(,8Z3eEY^KN;RL?e3:+F\d[&Kg3K;9[MFQ#WY;C-4<BT
XQN#Z#<QYD(1^:X/6-&O6f1D,]UJ=^5Z0V8-aR:abM3\ILPY8C(,.b^BS?KSGTd+
GTOd;_BaEF6T,TffYFTSD:\_3,ESZQ==O.JT(Oc)UF?IF4[gPNBN6:\AHLaUQOY?
4S.-L1^L3+19_(H3OdW@1\O.WT.T68-Ae)D/KA^G5Qd(/LQ6fGd2#@8LP0RYJ_U7
R..\GdRY@F6V@JaA6,IJ)cWR\XR@W>6H5IX4X9,_DA/;QA,e.af+DOO]b1QDBI?a
FP=4\dAW3bG8PB5Z\IUa7;7JY+\Z9+FGe3>=Z(3N[2HTRE]W]0=dEFCRagO:UL#J
(60\A-L(SAXd6+XJS_K7gDb.Q\TPEOb_O?YRV>)+M]JX.V@FVK>&68a[NMC7#?gX
P/C@1(##G<ST:9&-#Q#Hb]dN@;+F3?bf-=^5b<@?87C-N<dg>dHYR_;M9XH8-3bQ
8/W[G9Q#@K?MZf-I?Na[A#RZHYPP9R/Q.Q6_9KM=-fI=M0OYI4F<NZ^c[7M,(e_8
@ET<=DV);c).,eDHO_:_,3f;2_+XY@-K=GX\JRPTC=J5X&1GB)b)M-257Y2,QMFV
K9H<0f28:469_eWX1N:V7C6+_JG(C@a&QV657><FCAFaEMS#Y?KO&F/:TdeF]>)D
/@EE8aVa([DZSAL:_)?;3,K[6@JU+eNXADO.YcR]RO97F0D59UgH1]<:3dQNLcMO
T^RO[L[g#]d]1WOR1@F+Z[d9H1PC/<VPQ^PJ#e21;d_fYWN^Xe>[7&[Z;#/6<7J:
PP1UP0-<#IT?M;TLaQ#N(Jf,ZJ2NVR=NF,L,SK/+MT]gZ1O;U(;ES0MD9XPHL6-O
?HQEGC=/Y9Oe91d=C9bMR@FO,?X4F+#_F6]6N#[52PN.)_VGH2B\+1YZL>a>@f=S
DZQ2?:cCWFW@0VN;dP;_ASQY5/[R9bD;dDUX?6M,0#DO;RbFQK64dgZ+/08Q)[W^
\\.,f8>K06\,O-KCUAcA]_B1Ze,?[/PXAXXOP1W8^VO1SYYS97QcGd,QR6e;90AT
HQ_K4M#fC^5dWW[H/cW[0MOHOe1IeN7-+5IcJH/MIFCD[^X1PHV&d4^9)&HcRfQA
BH)F]V4#?SAO/[VJ0A_KM51W9:Q:^.Hd8;&M@\gZ()I7E=Z_/5bV1dbVOEG(0^NZ
OC#VC>U/^d#B[BD1_bBZH3DeP=c_BI.953T]OGNLVXL:#QdR?3WPF&ARe/If]&__
],)OS=32\=b76bOf2M(E[RHISfU1Q<1e-M9QE[5^J731KLf:)B6F/30(K2NaU<WO
V^LNVK4R^0cBF<<d9X.QeTQf_C.^eOQPXT\V?N03DK5/_O=J/Y4HXE-=F:[Cd<[&
NLGJUEe8&L4SB#AR]RD&M)WNd>L_XQY7E-^0]:=/F4Lb<YZ(O;?D_/<P/LW7bbcf
\aFJcP^4S.2YbN,HK[2H2Ib_>8,]2NZ4]c:;Ef[#SO#9eA7gA;(,-R@I@1D\Q(#/
WOJT+>g?^N/O[E)SN\^E9WcdMJD3NQ;^QQB.#@g@#M34L92=7,NNCUWSVGf95>9Z
28G9YARTPf)Mefg2L8@SW+1,&\QIgM]T,a/M;1#TPa.HfBX2:SY?EU:Ca[c30/(L
,2QK?+af&3V4BJPRH9]N(3IA5a8V0b2X5#AZYAQ1D@4HAN,(RQMZeFPe&^U)g^fC
81(U&U;]?a]\5&=Be@UMLZNRNKaZ9<6[+0?a.DEVDd9fM3cLMM-c\N^8g56P67e^
+CQMTDT7JARGRgM>24d-5A?^W?5>Sa[\d2&XK#g6Wd4.@ePP>XQVdOLX1+,Z-Q+V
0(3\(NQN39d[,,2QP65YeV3<aQVP6JUd4IgD6g/Z=HAI#WHW2)9[&ZZb:6)VLY8f
=ZbVDX9U262_9FY5Af8I&#;.=>Nd=+cX(?,@WQC^IUQg@4QL3)B@QAKG?+bg)T-/
S>E-=TAU^S@)E]fAR?88UPN96)^8F0>DRH0Z3X&d)U<?fde,WXR3TV]>DLJ:=?R8
+MCODHV/M@4F058P3.H[eL-52b;,5&gEa5O?<1<+,1[FN5Y/>AR/Z\GO^QegWT5(
LC9L,1(.99,gEQD;fY;(a^\IDE7YXFfUY#)UZZOdW/f4/aLGF5V7?-XSG8WGc_Q?
Z4GM,+]BDF5UNP,4)dL<<TU@a30\K9M^=02^#6+K9DNR7Q31cZd=].Gd@dW#Z>+\
1WKH#B^];]S[HRUK\^b56B(;I_0(WH9FZ#:gV/#>DF>A88KZAd7:PUB1SBC0VYTP
9O4gNd2>VJ(<J1(.gESag4/(c],B-PVT#9M#<A]Gd\,8TD=eD.];dQJ7W[JLe->e
.F-O-52cFF2Rf69=+X&KJ:25>+,[YeB5d;QZJY.[@d#W)(WPBT)Va@bJ,YLAG1?(
3W&4Ib7<+2a)5AGSVUe^GJ+8ETOP+0cU1;R:Gd^Z]f@=<P-)e5fJcDY@86;c2,fc
N+_^HY\dF8X/PGY(#V-SPAK18Ce)/AP+M)a4^0X;PR)GPdF&,0V#OFSBS2[c>ON[
]R1C.MW8D#4Cde55:33E5=Z)8-dfZBSO6EC]gCg+9^c#7Qdc2@1ebREV.V]T6[EE
=+HdMc4]/8ER7-2@&Q.Sd;+6/]7MdMZ=SWPb\,ZM7Yg79W.6IN,.BX76U/=L_W6C
;[<P9N<A\R3Fc8c1cgb_SY2:aU^BU=f<cDZb+c7ZbS[6LTQ\,NA>L]&2I1Tc/P18
KI6^XM=;0G\W+OFP_a0R=c=c_f?-Y=LdRWXb7>2EDg3:@PNL6&]_0)(_5aALLAa:
UAUTbRRJPf:cd8)W\d#VJ?/[[B,G>X3OZS4@:=0UWNOPGC-J0aIYO502Q,#C3C&R
>EE<Aa=]8N0PNU2REA8P]BV1M7GN1>O3:L5S?(fG8;7#dV7/:a\[9afbVH08cbR1
K/7c]f14_OH/bXd;?9f//8^b1.(\MT7eZ-(#a<QITQI?)K0=,Z?F/;O@gBLAMW]&
?OQgOQF/K7^d\Ea92I&^61:3gID[GZGQI,;fCf4^04E,c+R,)G6)0,^[\-2gO&#E
QLXcP.:G>(A:,I1CM9F?T5CI-[;VMTZG1I+[ER8GM4d?P8f]KF,?H9eea^H)0+06
P,S/Qd<ROOBE(B,T;Y&^JZ\7F^a+&#T.,fJ.H7/bSVM[d+,4S^RMb>35KCX_g>P>
JFe6CH39-W2-bB^8[(.PK3,aU]Y;(-aA54bb\gET-VD_YFO28bf-1_E7UU+]Vc+7
LWW:e)9LD6IBBW;G660?:e-9:H\(gT,>1?<bNYgCd>02Y9XJ#<5S8KA2c@2Z75XY
KB>d/G:5_FY.+OL?[0G,@Z@B&UXc3JR5:c>;U00H[07A),O+d+S?aG;:C.ET&fg<
GAW[74>T\Q&<ggM+Q-]Qe@1YIY5@1/_(BP-_QR98AFI4d#5):_[FI\c8]B=O((KX
I\K0R1YI[-C?;GcXIb;^J\;E/Xg_NXeg3D_HRF)B6=J@c&7G&YaD4_D^XTI]_\HD
PK44BFb8aXRY8WU7>:J[E]W3M5/_Z?@d#UE.R.==6T/LCgCA\]<=4?E,49/Z?(5T
;U=ad]DAX_Y=\Ga>fM&W9@EV(d2ZQKN>\BMcRe6D#Vb.MA<IN^6=L:b?I0G#9c+[
(H8+,NIW691=PH^T2J7/1)FQfQP3CX3@_,B5+RB<4_>P=dPFR<&&2(QOGc=H[aE)
ZfWYd<VK,X(<G^A^(8fgTCK;)]:eIL4WT)5U?[@4S-]LW_5YRM7BBMV4)eIYZ5\C
^LCU,4:1:?+1Z:F@#L2DcY[Q[:-)T-M\G2#4L76GGd^3[8))YXE=5K,_fE:OFANG
J2EC?V5D52,</HE5IM1L-_;@P6OA4\e59]e@T2WA]T).XN+dV?>??PX[75?ZLA6C
\H9eaQTEXS7cJWS@b./,+.Y@DSgcAd9:K\^P=J+Y\95cJALSP-.P3[N];gAN:;?8
5Z4,HFLB#:820K^K;WHc8S3753f8KQ26T[,0>7MX2K/^XgEEW0(8c)18#a<^14>H
TI7C)fID,>g(@8-eb/:QJM6g&<?2Kf\LK?7(BL.3.X:HMPgGC6>:(VZ72:R_B4.e
1S4B>9/4\T-4<VHV<3MHF5b.Y4RXZXM;2MQ=U5T6&X)aA^4^bPVV>G<^4LSQZ8#J
.Y6N4#77]-\OF_,.D/&V9]C>6)@1S][./43R\K31&>LGH(KVaf@?(=c)U,#F[.0H
YVGGU46;^Mg@ALcb[G6W57Mcc1/fgCP3=K6f95eTC,;4fZR1eZ7\GT_[-RO6TNR>
YT29<=]U8_=?#I)UH_dW:_+8TYA6EECb7\=^OH3)HLd:K=Gc4@8Z,25O752-ad-<
\^8Q)7VW>D6=PPSL2H=XV4+DaSU.6,F0DA-2YY5./GYHG_J2FW4A>.8L,^1AZM1/
TZOYQVNQaggUFCD^WW.1?13D<N;5@HG00GC7P^^)K(aJIZ/eYY1]4[2JUQQ(G6IB
OS0ST,T\=/S=ORPICbX7>>ZW[C)]2:M@c^bUO^FK3C5W+c(9^&0&^WV]F,5<0VDf
8f+F[7[<U[;E19Qcddb:TCeCL/T?g3b]88T=G,&3A)Y+_[GJ>aG<46.7fZJ0-(J/
@@\4H4>9NI(@L_6e,T?AVZ)@A0_6(@))4:7Y:&#S^^.12A6&)UF)-R6SG&24UIZI
5D)Z\E2+]/GGE[VUUSOUV#.T,P6U&P+T]>S0HQ^JIRVO>U6,a(D5/VU<8R?_V:+V
/;Q:W1<.BH)bgE&F58=-DU_+N;2QW^R=_AYbJ3A9KD1bg3De:&(YM(MBI;f;NIH#
VO9]6,aCTceBCX,(6DMLTH6Y0]9;:ALF[M+ETWPY\09Ta-b32(WAO]D7RM,,SLQH
FGCbX(\#<&9D=/DR1I[E0@gQbeRP_TA.7bQGVI51cXc4QO_UaYX7G<IAcAO]^9C:
&Q_=Y6.KS?]1TOO5>_[HF91G9B@/JUDf4g;F0fM-\_82U_a0;1#S9P.dgON?f?d1
<D/QI^&Q>@T>_79?2)JMY[>ggEIJ1SW^Zf\6QN.;.10\Y,P6[(.V2-84Q_9&)C06
W=1JK;\1&V;cZ[a;Wa<:YIQKFb[XP294HCQTG><TQ-R[9g#a,b?OA.[9fL)0A<XK
6>ABQAQ9WfeO;TT>f>Cd2_9f7g++?I+\I[Cafe#.L(^TRM^>_S254GfR.VZ&UH2V
&(@MJ6&-@RODU>dEJ+9:JF/U#aTJSgdQ:?3LB<JK>^CWB<@.#+91<]=T#IIVeG,C
OH@JJI+b9I-P<Z88I)8[J\+9FW3TKR1?^-<Lb)G^a]-FM7J#)Ib:SZAf(D_<eDGE
VTP[^dEc)4U8Xd0C@C;C?L=UY\9M/??QbXOZ2BK]KL[(aT2@5ILPZ5^V-;eEe:f_
0-TNIGNfZ^VHD5?AVQHL8;+P5:UI+9O,0,&bK>Q03.f/G3:\DAO@)Y]NMc5gM>-g
)?L(&\.-#e:\.C1HX6;TB(/;cVFBa#S^-4](2W6fR[QF6E<&STgX#daK=N5AMb<<
Y_]>Q.5QF-N1]W]KOR]#Q-BA_T-cDg_.]4#Y;P^,9731N8d,b.^Q>.fUOQ6?/eHf
YeXBMS7We4^E/WDPR+9,?+V125[2+K3,QJbY&#JTdNg>BNSNTKFc0.EePO>M/=QO
WY6@bCaEP6J?8(.Uf4P,17B>8J9ED#:1GCP)#(;>-7)&PXHHPLY9Z7RT;7IBW0]I
?.BJYDN;aJUY.F/(E6b^dW[O990\KPL8.?2MM?C4F[>GbN8Y8fQ#DUKRI@?3S-C?
P\A8\\JVN)KS8e1>GBE[:&=D&bPB^9RGR+-LAF=:R1<LY=3<(/.OM+I^gZDSU7.5
]d4C#KI?,MUf-+8#O]Lag>WS:<aO.9049)B.3=Md.-;Ea/3EAQ/bX5BdC\AB)E(2
,geP5^_RYXCUO?:-a=[BTH,VcG?E\X4<CNa^&=S8Y:9XAZL</_(PRF^GOSUYE>Md
U48BUCZ#V?;E:\cOI[P)HHV8XS8NGd1F&HZUV//?06I8#J;4U]B>H[d;J\R_-:aW
@R0a8/6cV\^eD_.ZE?GP<_-ADLeeGcJOg^f,L6X60S,<fKIg7]U^e?S4/SOH[0g.
2F2ZR>.-VJf&;A+7eg^d+e)b@1?C<+4_)#g71EOMKY?TLCf9K_^b_V8cDU1_I4(L
W\:J#OX.Ka62ED>0bEUae<##;.WP/<cJ3@.WEJ-DQD+3/6Q6[=[a#BdQ&--(/2S5
fW]80,#9Vb[0TB_-JJTAP)3WR/cBMSW@T&ZeYV19>-_CLA#_(2XXGK-U6>^4O:(?
-OIN#/aFd48<R+fceaBUa-M^.)6G0bYSR0Y.gP/<X^gV1b;36e)BF35RJ[:\=Na?
Hb1_B@#V,3_;cGVYaE+YNQ+^N.^=8J#CG[+POK\HPX10T]2IW^32AQVVUDF<Y+6_
LR6JXFGO;AV3<Rg8<W@F2#g\F]T:)d;dd_H=]B6H\E8C<P[/gRd68HbfJYCc=R)(
[)3,FPNA)WZ=J@KT4:YPFQ,K1<d(..S;U>R:T\SDTWEFV8/^-71d,QC1MYIa6QbO
VP&2O[N=(E4)D++Y?KDTD]UKM&^a3fg2MM()3,&)eE8/2>9>NH;^^]H>\I\c&9g9
d7IUPSg7=-8-L3AD&KgN^g/DF,B(/L8c(/e8O4LJZ,R]]E73(OFZgQ?gSP4[8V(_
F,d+<0-I&08,B/BV+UZ4)OKM&;#c=J09O@dO_a3QeWaeJP5WDU6Z@YNN_eJI&=^X
]([PMY=&I+LCa:9<_d;gcR,O3==/^(0b#]bVCVJAS65S)B2b>bW^d+I,0_V1P8MR
gXT7ZR#UAHZEK>A@_,,U_W&ER5c95/g)LI15dD=/+_R(O;C1Q:O[RKGg1-JObS\#
P\6d:&g:Jf>@FU6E=_-_0/;)Lc8+^(D2?_OBD97CaN0K/T?&2SS=F6=IHXe<BeC.
?^&f+U\)fR_)1CUO?/X7T[F5b+6PR./d</-4-SWV&._(0KNeRdKJE1>7N):5_GgM
?=B9eEf@Ba^)5L55f[Y(69d5FG,IgWN3KaHT<eV?=gZ/K.YfZ9Z0gFN6@R]]g6]9
S,)1dU^.f;0IdVdCgHRQDJ4?SKQ64a>\HU/Ee<<R42(dbDO@beA#/_2=-W<TU:Z1
cVbP=V-G0MX\>_3GD(&TSdGOC\8IFWHGR,4AE8^E3^@cK<AdO3G>IB]U)B/2;^-C
2IJ^T82#H0;>.^fYIE7A,T;9]gLNCST,-P6GT&FXR-4KHfUKQaZ&V8H5EQ[.Oa)c
^F#G:LE>C87;5HL<e#-d->,dT&WE+RVR7b8cZ^0>,CQI\LWA6C]>W&XKUa4F[3d5
E+3GP7M-1KBM6#8f:+DZa@SPEHX2+D>10Ga_QM?GB0#BU^:JV]Z9&C1#DZDVEA9V
^FOAZ;7G@];FN2Qb?.6S,fQA(?;ZCT73C\O.7T1c3/.,JY]be?U?0Y9HCdbXa;X5
PJ>JT]/C9/)K7JN>6fYR?3=>dfP)WW?F79b4cV<b.Q3:<62R[<g:69:YeYTg;O3A
XLC9ONc;VJK423E^1X;M8aUNJ6:H_O1#SbA1.TZAFdQW4gGK?cc[Z:V+Pd<eJ^VA
;fWZ3Ie@+L?O<\<RJ14,dFb/=K(2WKZZd/9UNV7f<,1A4TB?,eb:gaP0V<GEdfOC
.c+<>SXDQBDf>D8Z6c+O7CF]5<CB^1PDUK-&[g+^B6CM9>RY]fS6dY&LW6>bV/^8
JK9V2\a4?C3?G1OeF6>f833TdD#bNJMe/a5X?JT>Ba(.AQ=?LJ(\W;X^;G1[)a.H
.,\YZ7:;XfX709-WAdN0)-M,7(N=g6b9.&@6=+[+_>\_@P87YI6&KIE9a7I_EDGP
Sd)f#T<G(&MVLSM]D#UN7,88YOed-I<KS&^/M3PgI7b3+f^gcKgIagTQD0B,,8.?
YWNPQZ?<IT-YeZKO)YGUUF&-TO?,U,YIIgKcJPQA7W_75b-C[/=6UQ+SOc\e@G57
dO7O[I:_b,g20&GW6c.)S@T;^@;YGe1cFH3LL7LUF?.AD/C0,O.QbC&<.GOMP?ID
d/4&eO1V(/eZR?X4a5Ode+\fa,g0;S:AG.Z)PSQP599g<<X3e,@P-48Zg9:OcZ[U
1>:_)(A6f^DQVP)aR0TY5&<6@FH9QZL/K2>Q9eYK.bb(gd:^Qa#IEeARJ6M3E9C^
:6?CgS(d:[bK[.9:\8@Q=;Y3RgEfaJc#@+>P-A<daE:BFRe0/,(BLB,R,^R4Y^Gc
UJO4Q(RE5RN#<4C?7@G.4UW,P9e<[9CP.S+)>bWY.3=+?2f32Ufb5?d\fd(9W[QG
,(\I#0K1<MCSeUaA]]YfM7]3bKKQ>N@]82?9cI/_#dTJP)\\ZB@N7gP4:^_TH[ZX
B,F@OE38202agYIE5^<c.RD?cJD7[cU/dYX-dF_,8CDNHPQTEb6&LJ+A;70AJEQd
:=FCR<+CYKY9I5M&16(427F@/O3_6M<>&=D4V#20+EcO#1Eac;e6+_?M,K84Q@90
V0EB@2VO.g;<MU6AAQE77<_X=4(<JdYeg^I[]EVfA^f5I6M7QNcRY/a?WHDDO\;.
3O-L[BMR,7RO5.#-D^M&ea=Ob5L._8Pg#g&T,ARF9+&c38(Mg/<FQd.QA7Y^;FdV
f8\ZfW5g(.H/<=&LK#4g]Id7>Y7FE:Pg;HB4KN(/3VZ/,8W(XfT#YSQYFXLWL1W3
XG/Md9,a]MACfHb4>=.D@6WIS6[gb>)ZFOC]C9+.BM.bCO5RV5QDIe=/W,Q5[KEP
N_S:,\FJX4,-E@NIYAMUK,#^T5G>V?[gXe:.RSDRU0768AJ9AZE\+\/X>.8(<e-B
,5@DbE0#15B+N)YJU)AW:(;(3Z0M^2ENWO#D\YVYG@N)[,PCWF<d@DPHM#e?&f-3
=Tb5UI3DYG13MS_\\G^C=-41EPDD7>;E;K53,MAdTOB0,[<g,^K=e?3\ZBF9CJ-8
eb(CQ+2OCOINIKRMCb^K^=&7F(N\<@=?+CV.;HM5e6(HeQIXS4C./@@ff/_?EB,c
.\E+a@HebD9L643g(FXI8,T;BB_CQVG>gF0<Fd<YW>d3NDf7dZF#eV3M7,YKQFZK
I2g_]<86@7,-NNVVARFC??dCH.,L8b-0]?_[,CS2,W:V+&:IS3/#DaZ@X,A5[8ZW
<4d-5TU<(55#4O]10FZ\^ILP(H9Jf8C_Y:c_4Rbb@SaJ:Y4eMFMV=[a;;-4R&-1C
;bCeL>4P<AZD79:WGAaOZ+8?3Y\SXG4_;0>-_9N;DV&Q_B@GCe^N;V#:25_e5Ta7
eZ;[.@,M.f[7W1(eOL)Y]RV(M[E67OA)VD5GQ=01JZ,\VRa(@N:A<4PWLL<adYLf
2Kb><W+FL6R:)WS<faWV#]aRX2(-FDI7Z>)3.^]@AR,#DXNFX(?A=6IHdDB.WeO,
Z2D+YS5b-a&=AI[8XL:3_-I[#?4.B\UH8Jg+JT=OYYa06A<6T@cU?50]9J<=/9B#
@a>55_Q&E8cR7ecI=f2M/5CFB6_Fe3.OI_[U-ND7DQLOA;QQUGBZRW7Kc92F.;=-
E,T\SM0X&:6Kf.&G-TA^aFL9#-@P3P&TZ8N^#d?B)4HeXJC]&RM\X,7CS]+\3.3W
Hc2#cCH>=S2X?fJ8S+aPO8Z0Z+BIX@EbB2R3[1W)FKaD@(Q8M>JQAgV(BRVJ:A0Q
OJ]@\Xe4Y))]5fb2D@<:ZK(cg9E\@2O6O/(D#J#&5g])Q>R?Qb0d^.N-^BYH#1QJ
c,_N_(dA:4aB/c=b\g-+d],L[Y,?e;V0TU:ZK57HIWO/M)?e7[ZJ[HB5:N0J[Xg\
QG?I-8XJ;=UIZFJD1LA1Q?[eOHc:.RF;JC?N[42?AbOV=&UbN[NBL)EW;#MG#GL-
OEZ8+B(NDZ>+1;DTVC+T_c>Qd7?:UCC+?FP+A5cMg6BUCD3WV?]LW36DSNAX5QQ7
c^XR1Pffc2(@(SD)W10bSFW5e9B5(9b?)&[.4B(-g11CfM+7:6H^b4N<Y1)d[<f\
KL^CX:8FF_(A5:<JX[LA9;P3W.:Z#;BaG]2[;T?&e8QO[IE/YO@?C_I_fG:C/SN4
X86LHGXOcXF(#AH,CQ&_C]W?VP7>#UXKV^A).KD:K>]JN:]/2I15cP9RMS[ZRO9L
EFbE6R.TP1NJWO(;-<<7VCY2Oac^D6CBB+)5fRL[@G=-ON2eW5HT4X/[3T^+?QS\
E89c5)a29[gH<1e:/1(SaHf89HQ8&>_1TXES/I2Ca38>aPJ_a3AeO.&T0#B8gG1\
B5AMYTWW4,?S?QE&R9J.7RK341:Hg]87R,6/LR7MFb9=_J3a00Gc9D<M_J8a1SC,
,K9E;-O5XP;gHcA,D^>5PQL4eR/],MAbeeW[(Fd#_G<ZfbXfBgQ<-<5@G]5HBBB:
LY1?H96G;J_)[0@?Z3<T#DF\K5M>SEW;cPIDW#X&XAC>ST,:97eSBbV3-U=SW?DL
OL05MF#BcD0M]G7=07,TfBUEU>a>+ZHaKCSV10V)YAAaW_U4a#ab(Fd?d_3<N9Te
.IfTe-\.\P\-bd+JaZGgCG&FfLQ5IL1E5_dD)X+c\,7:]E=AXc)Z8UeL&22DD/E4
V:I?9>RC,=8MC?88T?>g:O]3(WAH3#A+8_W^GRda33G=M#MU>1HObHeV)YI-c[O#
Y8@?-7>;@&H2MWa_U:#GS?&MQ:&fDd&NEb8bY/PC3RA1SF+A_A_,1,,)G@d<e7H-
]YXBA58<4/8\0A&-5-VgK0bCBH4dYJMSF8c13c)0E2U5Q[A;)K9DF,MKg?fW8=TQ
/2F:69LX(H_K?FJAODOW4R26DE8M1>+]bDD@BLZNA+Yc#)O8FINCROWZ.IFS04,b
+APLT<R_7cf]4HS>WOFc<(MXbWA-CIM_P_cC[X#d4:LS(WeYXH8O10,3/f=:RN.3
=.Pb+=R9_NZ8_T)I<Y9[WNaf:ceXZPMAQTEWbNB+?J>&a#6@g6PbP-+7<:CNG&bf
)A@Rd7T&-QEXXFeO[_^f=4a->P1aaNd?8dLC.BN0F)O8=F_<,g8<3gWX7;MH1JQ@
@8V-J04V-ZPVWFW,-^=7\>JHSE<(KF)N<D8MWUJeSceSS]?/Z3/Q_B[)C)=c47H5
B-PL0BdLFRb9VTZ#66aO]ZK-O?I7U<3cbJ[L82J_X3BGfQ[+8/..O&?>0@S-/A_T
SRUe\^fa+S+PR^.,6X5aP=/=dYOHA?0U:Yf\>?<_UAG>-;Q-F\&?SW&T870S^867
YL4+:.>UeOHGPFba:TQd1P)J97,cBdJ,[=.b=[;NZ&XHTFA(X.\56#?eb8P76>CS
MZ+3Ld5(afP7EDfBB,#B\eP-\Rc+:8G(]Z;4\Z#+YeF64>?2EF:A:VSKFD^D0K]W
^X8@a3(_D+eV.&XKNHJX+A<5,g(M:R<@8MCZ8-H2RU>X2<-2L:fgc]c_(,TAMB@I
Fbf@>TURFIBJ6[4A;\I3L6VL2=E3.bfQcaW8-cfD-9ZNf.+_\E^^<JI8e<4Jgc.3
Idgc7/LW@;SN.0.g6(>ff^R_<G-\f&_d)]1CcGX[YQVGNDKc2d_K=CMQ\&&?PgWK
NN4VC-5df7ZcSXH-@?R@K(cBZP^ZUbYPd\eKMSY-^eL;C#:;^>+:70SI=TP+BS8R
YGE=0=5F;G=,[SU3_<-e:_4ZKS5YN@^@5LCe-T.bR=P,7e11/5dN+/2T#X.:#5RS
R\Z#>ZMagLO5QP:0P5QY3LJ0@Q9@a_0DBK0T4<CH/\3-<Q.2/9b,cXdZ=UJ3cfF:
V0H6WGS/JLO?=(g_a+PHH5I;122HOZ>fe7aU+[]_03,g7a0X<8bf^BWc@&5\]VdO
X<Z,?geEV#&5a487d@5;..JX1fJcC.4AG,F6TOOg(X^V,TebdU3X6M?E04KH:SK8
:WZL<CZb2/?b,FX<=Y1e#].?G2b:0-<];PJLUS)0F.DV:(Q3Q1YfY(#=WRg0_bY9
:7W@4W-A(gGB8[LM\UAW?@.DE_@NdA_LTJ46\VOPQUK[1FF.W<_K=YG#&BLSBY00
;5)2:Rb(A2]M:K@MRCD?_=E^WYL2VRVU>>O1_)d4.5V-J[bf6\F0R/Q)[19YPad2
\I2NaK\>#NKcGIX8,VKCdG[HSQ3UZHHcDT^aHEQ1EBfI\ZP>8JN@<EHQ[C86),JX
OP<SAM<[@[)4CLGg2dNG590;3W(V,ZdLIdP;?6/bNZ(LL>NI-/baFaY84R4I(_/X
ZbY&PI^S=-/S<PEC0&0D37CTTb+2UdLJ73;=8ZeC8FWM+AA^&Q+>M3\PH-Sab9T6
UAQ;-(,@SE@M7;YE?((Q#RB.;<BN<Z..;Y9([?I87##[1^MU4F3UBCeT/8&KcRK.
VX&-g5fJ(#ER,88aAVadE.@M@bN\f)VNH5[E91b=Za_FYL-:&Z\JW:K#g0Y#8-Ua
[\AE4gc\U>1U+I15Q2dNf3MZ<99C-b5a)36TP3#@-9ZUWFeePL;e@?5?+T])1IY+
^(]6]GS61:^M]KVA;TTJ)P=U8KLMGE7=HZ\2ZZEa\0T>-/d9W49WN]gK0IK=)ML5
P1;<#@6=4Z/8[8@UKPdWXYf\4RD,S@MRQ.8f.0]JGL1NC83PYf8-B.9:P@Nd\#g>
AE6Qa/OcSZbU@NaG.5S\,f_E+(2M]0@7/0Z]eO;2\-(8C9=7#6OYF>VESD798MF>
7[Tee8TL^0MGV0CWRMd:cd#;,(gM[IAGJ9-QUQ)8A/)KQf/NWb@Ha2^U;^FG=45c
JF_2R]>-0;e][ZJb(_@?N:7AQg<TJ6VLURA(\LCM(:&.MR3^>S8JS5e[H:E5V27@
:?#D6A935G<S].>>2N/+.5OE8JR[,G5]7@_3;Rd[<fQWPA]E6U0.8B@Ee:GTOE>,
T:b_L]7(8E2RM@H#ON66;fA[G2@7GgM-?]03:6(2SX<W5XS8Va4>O[C7Xa[P+GUR
V]M0N7_95(MJ588f\G4])EA9?_B4NS)D.;I9c4F6)VfWK)P]aaYY>bd<I>DU\9P]
L8<<S4Db8[7g3Kdc_L>GGA0[<Y?W4:>^d1@[GZWc3f[WVf)86C5?fGd363@[+H=O
-T>/[/9;/Mf=FG]?:E0/I-[1KgO&Q?#1FOC@?=d(RD+A^dK;O).4Ed4H8gT87Y=,
).cUCL0c8fKD0S#Q8ERPCfJbYbTW0dL9F:-@/44=/4;[6^U66dJIL=O&FLQ0JBJ(
KKU=]ZF[dIDNC1UE;7WF/QX9MJa(XM?)f-1&Q9&]DC<R\\]U./>c9[8+>Tf-eO.\
K^G[R03QN=daO#:b_OJ[>e6W5G@a1L0>M5&=(YR&d@Q-efa#=@EedG=^TO<NF<;+
XITO2a@Yg,CIBf/\1>Y6NLdMQ<Vf,J?FNTXdf3?Q=OKKJ-DKY@g_B[^1HWDUDA9?
-YE3G^10\;D-^M08=RMHedFS4>L[VZV9O(/K&NMH#F:5.J>f-<Q;dF>1]a+B\&>6
0\=B.;XXE/ENZ>0H1PU7=?U?@]96=NOc@Z2deX].4Rg?-873&9b4K:YN+3,a:@CW
F(REM9]7AZ,&U3W,A1R7cQE;M;@/T24d2+-_55E1/;gG=.ROHE2I#O[[_bHVA#XT
YN@EI3F=LXaFO^5RS:/@G-+&(Ce_P&g=>I,:EA@VA-2#^D+;T,X342.?PR1;_JYV
ZPH]ST82Q=Ff_K2NX,-=WCMdbfMXH[;6>^c,MEC?4#8:?5BBVcWCaf@KD#bdCKZe
JYTH2K5Y[YIE3^E)Q:^g&FT7N772@b24U:B>#-H]]f_T6WG[],D;_XO>Y5TN>7&B
I+IN6a7,e;>Z.57[)SMbZ3A-=)24a3?.]JcbHb\:N/ONS53HdaJc(3ZRgcfYW7f@
0LWYA@/eab<\V1N+fBFA);-G^QRKe>#JRXW5+gg+QHOLA3:HW8/;ARQ5J]WBMM/[
+4+Z,V3ABWL_^CDaH&8E.A[eOAV+=XK.^;d,Rf^-EF/0Lb160eMK\9?L+1@E#US0
@UK1:F05A#NPNZX:Q7NKGJE3QYLD72(BK_N&G=BW@39PUTK<Cg;?<X@UR:.f,,D#
JXSHW[3&]<UU+ZgaO9G5TJI^Re<c@X\+Ib;YCZbBRO3WWgD1E&9[H^_6J,L&/,C1
fQZ<)/GbW,?baH,@6G^F:8e@09XGJ];TVdV4-44ZGdNUe7G)ccF@/P]:\)#GAgBM
MTIH,)_U-2,@]I(LZH>Jg)24XO.W-c-9/Aa]^8gd[d]9/O2=][#EO0?\DNC?>P\#
a\@Y4Q/B=PYH>KLYHL?G2I+fF[Ea(9M#8SKMc/G+3eJHgZQa1.^T1[Y;c[:CXM-X
U([LcbX]D/V72V;A@5?8N@R#&8B3#7D>(f1>9&N4U/::V9e-FR#CRU_7[I5=>GJf
9^2(9Y_bQAeT)3X(>2P.UF;L(#Me[5FPP&Ld#\LTI+&>J.2/I\RSc-\1YT>CHQD8
UZ8U)aeP.=8FNZSJ,J=gWIJ)CEaRI+46)21+-.\;GJN+N/Lg8^:=MQNBa6FX[Z7#
0e@M6F/9)R7-4N7f)&+7WHab(S^B5S)6=?e(SUBCJ/Bb4LQ)b:,#5Hf<XP7]B.DQ
H^-)LUAR4MV[33Q3F4L)[-MXY(B9X9+=+BX=26WCM9-+GXT@>9d_8[T(dGffffA]
7,A&CS]UCBZ4.4PZ5G_F7(I//LFVY4_b>f1eK:C<)TYR7Z#Xe6f-O(Vb28T+O.W5
P3X9N&+c<@;1_+6JU2[/_>8F?3FY9PB4]M2M65NB2#GMVOW=0[E,#T<\/N^g\QT/
VG/2.Df7#?(4C-6/&C0:?=N]AV.?PU;-6>Z47MHF&W^\EQS?3H54Y,YE+(@FN94)
O:b<3)>K\7aI,Ua1>C0fU,f>=YMNf//DKKdXMNV-FM]?YfdZ:1XL4/Y^_/M5N6U,
W6R,V53H>&I1Ma@&g,?6-?cAC82)@Ab3U#5aMNFX;cW.P&#cM_\S4AeeD&LC<d3-
Y[g9aMT18Y(,GPDbF#]f;FQI6L\LZddcKc76b.7NPa=AFg)RAgWT.Ca8O0>M[c6E
V,6S&@SKaG8XD;+G/c#KJ51@^,-9[5Cbd,gf;UBRF&QWR9B5?J;@E)_:@)QI+3ea
C?L?JXJ[d7/D^I]CVP/5K^dP-4.T]:.RPC;N[gf7Q3AOT&L,P_a=5f:d(YR66=65
A[B>51=+A2P/2X<9RHH.:VdJ&JVRe:DK8F5ZM;EJ=bOD(=Ld1e&F>.e>Q-&Ia/PB
H31?d\A7C_QT-YJ,VX0:SSL1CdOUOX)T=RM)IN^5:1_]TDeK8/&S/&)/#V=AN.bd
f7Oe-Y)]QD>0I91A3+\)IMEb/CfKZN<+7K/RP5FOe#ZL8VW@.RDO<#a+>Z=24#H(
89G1D+A=1VO05,7H<YC00VWOH/@X94P0>;P-??e=2d],U8;\[,bBXZI(fNgK:#[R
bTQA\3R>N/47?)f#^,43<2CbfJ_1DUAX6gYCS[5:RdG)FX/MCQ]dFE=>9N]JFb_@
2A=+@I>T(K8[+(1@Y81Vg],QLET4Z;:[B8J>D34&P@&?CYNc/.Pfb(K)6A@8.<B2
N:--^#.VVCd[=DG<9HC+;ZF+#1#eO@@Zcf@,GcAZL3S(8Q]+-OH5N(+8Td.>QP&Y
:&;NZ/ZZU)[=c20CVWWG116e:=7?CC=R>fCEC:G7[5#6O-d5Q3KBP7:<==L@_=PS
IR\bYdWG_EJb[Za=>\9ceX+II/1>4cA)V4cFHFJR^DKJP<\\aV=<&CR.d:E-4W]/
;C_-6PW0\#[cVZ.HDPC7R]&[MG_Jbc2fFI)^XO36b_3NSd=<V_dL(\&P_[XI#:UT
a1-a.-PYYAX_R3MU]2JSc08LcMR;f-:DfWXDQKf:VU-E3B98(d;[](D87LV?3bNI
=J^O??&DD56&c^+4PI:Y7?&OIa&S6g7KIYTUETUW@#W_VcK_HGTZ[57aB&bQ-.X=
Rd88+,fHO0/<cB.ZU6.4^@P+F-7f[(P1OQZg72:aFfCP(0X09Y4Cb?EMC+L_,,Fb
[f(NXRG5/Rf;1,D01=K]5TaZ<RRD<=&D]]@]03Z;cCf])g@S&N^<P7:[T\D_LJK1
cKTVE&6I@>QT0VT0-gC?D7)]:5Z\IG1f_Tf9U#KCM0H7ATc68Q)f(F]2&QX5^.7a
<6fQa^CCgFA=eJV52==N9S?Vb64+F9#/\0#F@e-V<Q]ga73B9KQFcfWbWB6.MHK:
ZgIN(E:NUTFH)NgfZHa,[;8MbX4K_gAN)a[?[W6MSJCJ:9+,VIS&;A)DNdHfZ(]H
(K(HZZ&ZWCFUYWeI4KJ;J-fX/BedL?L?:a.;H8(;eB:GMLUeF.6F,]?Y2c5f?5Ae
SGc8UWN.C\&_AMZ)#E>PZ;+c]1G0g]GeR;9TZ#X6aE&S^]WP?R^4FW#X64N?NR&H
;ALI==2f1SE1=>)D?Kf.4O9WO5J=UXDe;c8/e=POAaG_e=_g+GEB3__@c7Sc1T[7
CUP&5<CLA[-,(M:DEb>)a:f\.d1#Nf^1A<VA,K&#.^3&F&g_[+>WJde=T80@2#6E
\,5G5,YL5(9c??R>g4\<d-85K1BONQC+LPT_D\4cIX5;OA<9REG]fQU:8/=H]2KR
AL8R<@K<@+E\D+TSDJ<_#A/9T@^7g[;<gF<?.DKfU#C)JHefN[=,&G8=:?S9&^KD
6D#(bGLD>2#g.S\PU[R\NBDQ,&5CC:QR,-V^35H:g68>F\VD,fL+e8cV/.>D^N-)
2PA1B99dNS[Y0^_:@gN6c8U3^:[:L].+_:FRb(&ee77(]fZBS2D)cHa\Y8W1KWYb
6T?_HaSKb0)X,R&JP((L/0N.K^IB^\]#E,K;80b8aD3GaZ,G]CPSf+]S(BOO(\:W
<FSG.^e7]9\WB>]:&D,;.<HFg_KSQ\Z=D]?0N4>fAQ5;@1G,D.ca09f?O#^?aZ:(
.7VRMd\EVQa=:C^aHg6S4I&A4GONFDPdfUA?\WUU^Z&TWER[O31&A?R:2F8dPFUc
[IYWE@TA(fA7=TaIT@KR&XPD@e98OdE.6&dS9/XN]2?7g/&B=L3>-e\>I/X0VX-E
9dYWP2YW^fE#2;WNTK^A,RceEc9T@<WJ.dQ<1gA9JP4N8,D-@_:=BdR+)?SLQ2;g
.][XC+Q^bQ89FM63[?/,=PVL_HdX=9#[Ja6&-OV+;U1Jg7Q>c,dbXb6//^I6CMC>
7U<R<3C,FPeAXF<.MXJb^5EA/7\1[17aDdYdE[0TTYWSMWPXM8(FMg>9HZF7V4O^
f]a(F^HMOXN9e^6F>RK3ad=,E[^.gL9b?D(_U-fYVaML_+:fc7C[XBHNHfUe<SE8
03B/bFY;ZPYeXYA/JaD43+ZM#eMZSJA567ZaeDg=EP?NQPN(77G0A.J\UX/f/-[S
AJ48d/VfFWDJBZ>[K=R1aGTJ5:c.+5KEeF?a(UUeA6<&+4O8338/R[aDRf]TC[9H
:dFfCGW1f&70R9Ya,#>.g0T6:;9K3/#dOF&]C9;b?IC4P/;\;>c>21>6?UFDa4CS
=\JGP5ZDd1#b]+cW:31W80IIC=)0L];JA>2^Jf=06#(T_7TNdNR^?Tb2+0)@,c2H
@76V:Q=T_S_4P55aQWNUB^Q.-\O_CQ#<RCTfc?NU./.-^A8Qcd@KeRV<cJ-O<5a6
NF\?-P)KFOF9G:YcXgSb.@M;L.V((gX^5+Cb1C-S0BO^+-UbK0A1Ndf&aa<?-D8C
VCRbA:^Z=IXSX@=,g;HJG4D->+eC.RG#3gI0XVC[(>)C<Lb)1#g:,FRJ5SIWM@cf
U90H@#WON8W2I]CK#H5>^_7Z[::g_K\bZIP(Z4,>&dJN:EXd);4@GX?FAN?-\PKJ
0QO)>>T\H_J5OVE<c>^Z/c(FV(cGBR#++H/2<\6^>C]\R^9X?)2&Aa=#<UO<6V4R
KMX:HYR::9B,I=4N?KTNY[#@.6_]F:5W_dgYE+@M+HJKecWO+)KT?+QLW_&S7WD0
g6?S#11H4.CG/,G_^3_B9/WMCF9G=ga=HSB5[WKAB3-HF0V?aeLXBde-4MQ3.VST
,gL6WQLe2?ca3P7/8P0\372)PV1CMf7CINGb?ILVGW6Q;TPJ_,#[\-]UNL_,&K_I
<0OR3Y8?@/SU&IRCMK<eMcIdR0@B5V22H8f>,RROD8FO0;CR#[T+W3S6N<16>IWb
O;NQK43WF]I3>=Zb4E34<Y;=T.PF,)V/#M)S_DC1,/=H2>OC;DH?4#8^U]afBM9T
I,4MQcQ/:YSEecF7LeV63(\81gM>EDdO,VDSL]D#+3DMW+,WQMV&ZFMfXU<F-)F:
<2KU/LS]KN6Q392O43>.#f2?\46W^@S&@f(BYZaEM2;.YX2XXCIc>RT(gY4f:C)d
SDc7.T=A)K&UJ:YdDVF>,SXC;WQRSW-5O1[O..>SL76&C[7;P<afFFXKM2FYYTD@
UL>[4DUg5WAcWKa3JEY1-7fO#Sade]C;dX^W/_+Y3Q8C?&TQC^TfZCM8bWQBY)0+
>X^3^48Bd;YQUJ+ON8F>@T_#^=NFBZM1_gT7J2R^A]T1^A9/U4Y&,?,63AVJK,&4
b]JD@^B5I5\T=/_P/0L]<@CY@]T(=a,P?169^c?-K=RY9IKBSa=I?G#c[W<PE@>P
B#VdRH4W4B93^aZ6L_Fd6(\fa1ZLYUfg-ZW1F]1D=;JZ_/E1+E+=80@b<>]QY^I#
G;_K0]00=[SDMSNE,Ua4]?G+5^H&.@OZ:_B4b[[B?1(BEPg,=QY+_;+UJJB;.R,.
^BIQ#_URfRHOEd<GdM,=,GF43<PLV3WF[g&4YXfGDA9UIa>^A\Dc7Rc5ZME44(RM
BBW_/d_9?[QLYA_5F42)fJeIb)S-B)Y),+1LCQ-c]Z+G2HA2f#E,:#3TC93eS01@
):IQdXH85A<,_TW>>LMOWHS,/:\1II&]^W??c=?/)WMGD6\Y_YH+C]R#-@.YA@Tf
dU:.M<MD_AB?E@ENPY)g/O3b5DE#X]K]M<01;M6W>Z4]UG1DGH<:\JZ<bM;#A0Xb
9[U]C:gO:5J4U#N?M5gMD=UW.#M5(bPeRBA:dWY-,BB3cMUX&5dH(/^,)M_gW-:6
=Z@C<VPI0^[CH+<KF6eI+DF16L9>1_a2@R34_F(]6#W<HeMK:98&B4@9#A7^J8V9
&JMBA1-X.8/9\G=)RAOKNVbK@&X)[W82094?)cP?W=KX/L;U#B]O6dRdN]d-H)<W
B-9IB7;F-_H+JfWI=EAI2S.5F,-NW^F&IW8:[>F0Qbc(T\Z/@58E?8Q_gS1A-+G@
1LQY;Q@cY8J@+KTZ7Y\:D>?;Z5#^ee#0C03EG2@.d-_f69,F-UV;f>d^M&(.1c0F
]H=;05^aM;,AZgEMfQ,/0)KU==E^X5.=6[+[dX^D=9BBRA./U93X@8M2bU9S[)b1
NKD.RBO:,0a/-Xe68+H/WJ5a[RZYEcX#_g8<gXeQ6HeTSX@&5M0NGT7[-KSVc[G1
@_]:&#)Y/QQDB9aWHHBE]LROMAW1#6d)^M&Z,eP5_K(1UT@I><;:9c2=EN9=9Ff:
\9Z?[R6G&K_WGT2X(?F]VC2(CA:>E]OLbKVBAQXFY5Y/#b4c;J]bHOTY(F<7KFA4
.MW5M<;73UB9f;^9I.#aI9G8]T,V8^E,dB7LS-,-\/^C5^J;SC\;UHLW(=AYZ):J
,5[F]d]EVG0XcaT,f[00Z721/GS0cL@7ad/G&?bS:G1V4;aSXPZ58&P;<Y]c2J?0
aYJ)RYIRa+0.D>DU^]H6G1B-(aW(>:c92<B9X0?\3PeQ4<8NJC3MN8g3PXU#=M7=
L70=MT9WEUc3gJGMUI]-S56\#;1796dD/0XA[bfRUcTLDTOL6fE\+.[U58BXS&I[
\512O(-_RTCLgOI7KO5CJBM=/:[Y=9?#gW&5H:(WCOe.^WZ1f]ZQc,=3C,I6W5e^
TR7_cYAEMDZKZEXaSIN)3GdJ3YJ9WASFVXVT;V2>U_Cg95Z9\=aJQf96-^S=gQ1(
>.3bW5Dg6c4B#AMg3/_&(O+:U_b^PSZ?aa<bHZHC+4\Vd+#/1L:G+gBLIV^HI?X]
ORdF;W,;O7M/N#Qe86Z7N;J+AWTQCB,D2VNPK.>d97M.5NgJSO#=+1&TP=63e8Ga
D_DS?ULPFGeNW79ISg[8YT==b@R\@/Ba&RB(1A/Rd(+S/eN0fP5,+8#14Y?gN&[X
IW&0\Qc9WJDfNJBOD.LF.B2-_;Q./JH=9=TZ+@EI0&OM(2VbB3>?^[cZdYLB;,fQ
L8VK(IYQS_T<^161#aMC=+07]-,<8:Q90+(IIWFIb?6.5ZIdOa:X3Z.gMPH9EfGV
[KCFREc(=Oc0Z/XKd@]cHT;_-6N,1e6/3N,aVIK-GHR81^6N[VW<&__EU]G)EHdS
4:0e>dCO8C[5W+XTdadZ>eK//ECHRUA/bd)IPL//7A\&CB?]-.D>[-[2Db\PLYMM
+<R&+JY(/O:bQY#1JQA#DEG@_C_9)O_ODdU\RA[:6=2E,8\J^^(JOI+R+]?4f#D@
8d7BF3_-?.9@\2Y/TW.DVD,SO#X5+DAEEH?>fX2\C1^e24d:S37NQ;3]&X61U=DZ
B.<72OFgG+Q@&a@17AH&6ULd]_-g;f6cIGQ><Q2#80cE5WDDQ;</fGO-1R7;G7bE
&GI93F<-@[E&#G9QLE_-+9MX,S6a<gI5VN90T9?1#OG=a_FX3Y_YF</#;)?T(+7,
4-N\-?IP)VZI2_NPE;3TCJNZBabR(6dP>PL(-5[ebSB;IPFQM3I6VUf?ZD4EDRBP
eTfHVERT7;[_g/1Cg7)fXL48Qc/Ua+)84Q0+>\5C^IJCbf#/BD)cRMgAR=FVH7?-
,0dV&?R^L+942:_23Q>IQ)+NLAdEZL,,SWBf?LEALU/THX@OG:ZdV[YM+Q^QEO-2
DZ?UKJVT36E06_HS>fZI_a\G=(;6=B/,d,_-Nc(MJKP)1>bb+?YbZ[)HQL[;,DAd
f>[]CCF.^B,eBb_d8Y@#b@SK5aL<#A#8((D0b?<d(DXK]&eO1Z(37X_9U\MNf=8J
STCKH;M_f6VDV<US.H;-LVdOF5T7)I@?d7_HIYIW@JdgAYZDP<JG0Y2&#:fD-EU/
N<^F/\3.QDZ&/&K&]K&Ze3L)(WCbE4V692-P)2g2TCS@ZV?9=L36J7dA6f?@4TA>
>g@L44b:_dY6c2^fI@#bB(5JDP-1UL\>\ZFb)0.2Dg?[E2a>YM26JC;OYEa3EVZ1
56J<9WH)Vg;\X5_4.d17S\2:9\),[,E@J>7S\Z:V<MVPJFA-_fR-N\75f./S<L(^
X/e4bN^0(YW-MWW5B).GR1F&SV&/L,U=dW9L>P1&CYGE@NR50U1-fS5WRS0]69e<
)L8^c75LGZ7IWaXM)ESW9?>5DJ3d?3VeBg[)4^.W\S#I&&]MDcaI<=RNP^@@#CgJ
QDG#.De,.,_5N1b;T6R.^d\#+/<&VdLUPCJN_gI/MVZ;Z>?1;Z@])7bc/OI5R_e;
8KRO6BVZXCQ(N1G0@/eA=W-[-696SY(XMGP)e85WTf,aOZFYfL<K[g5:DXK5>]_N
e#BX7MDMDAT60F=PK-6c_NG[SgJ#TTgIWW1ES#@G?8.c3>1ffcFOSNU6#CgQH^0K
#TH;fILAK\[/D<8K0NcZ.QEHSQ+IDML6M;1W8P^MNcGWT>=K?,#1(.<_M8Of.U\P
?g56D&6\aVM>?2EYH/]N:aV68RA#M[][c3OYcY3SMSVM,?M<.MYUI5N#]Q63DUJS
HgLc-QOYd1EQSX-]>6&g^I^:Ka-9Ef[fG#\,X\f>6T212@IMgP1Ff4O6?^7E1CQT
fIdCO-/DGfL=b\)TEAOZ=Y@g[cGT#R5Z[ZD1#A0>cI2;F;Ae.d<dT#aA>9J<B<#1
CV[FefTQZC/OP#[1PZK[,KOUTB><;]WNWG4G&54)Ua/M+@XFHaW^<A3PH8JLO\99
O.5<WR&e<XKVA_M0^&Vb.e.Z@.f;0dS>SgG^6c)#1XA>SZ49M]2?0=V[bWKWIcbF
g>V]g&4]=G9NZ)C+_Ce@+-aYWK+.B->?5DFKBH(#PM+=\N0D9O3Ie-;(aE5CA9Y[
:@MF(JB8ZZ.c5\Q)9fK\]=1UEUKGfF=:6baLN(W,6AG3;:^E#c2(^UW,7CO.N&2R
54g=3Q0A;:XeFD,]=4B@GX=b7(VX<Bg-EFQL5AW--(3L30ED,=,K<L&._;OF_N<;
HIQ-4+XG1?=YU5T(CC<,eJJ(<=)=e,(AVO(:0A,.ZH\:M8/2P+ZC^.^8\g5ORPZd
EX9I2>3]HMZ12Z[M&Mb4(A8]3_VN=K6N;O<Gg<LOf>,b1:e&9;)-6L5B>>M^N4IB
/Ff9&]9BA]FC2Q>)0e66?<F2.A)5,PF-#<CYXB\]\TPe9+=.3[PH-VOGbb-]fZ;>
7Z9K]KfXTAHeS+._Q6?cd#S&:&W-VZFeL9;bT&dDM_0I^Q#b#4]FL4f>L^SbIH5O
VS_1aCRSI7]>M#d12;cP?5GBE6L8I?[GJ\[VMCedgaPB>0Lg9#\_9A8X4VG#20J1
1?T_;<[7_CQ5ecORg<gKdRPe:(DB2UbgC6YG=](SG&bM7Q30f)AHGTaOc2C?d,FM
UA8:I4,#Lf7;,CQ8-cTYaYW\H@E#a3F26YGYVb6.RO>5NZ]3O^LfDcMb+.g?8KPA
N+YGC((d<(2F.91,7X4?#FD]dN/^Ef+5D<-^@7VZB7?+HS5WQRM1D#R)ZJDaSR?e
6K:+@ZZM:a5Bb<^+;VT#52OL2\?43D563XKa^,_Sfda9#18;P+YDD+g8SYZ]eFbV
IIAL_GKUY#,d5[O0P1_8V;>aaWP47DBGH+BLAS_/:_d\XP7TUWPR_B9DcLHaTF0R
5b/Ob44D^@B.))9/]V_6+1bW3NU1.NEa?f0eQFaMTQ7A4RTgG;Y086-(fX-QE-2&
=FQ>,[:ZQ]IDR,DT#>G5)S,,9[-20bT(\5973IM/?VPBLe;9MRd89K5U._D=@Y@U
6ER:P8#8F\YA;,P&BaT93L)QP<MNJb-LAEcF:HJ?3Wc+TSK>_Q=S1@;fX,97FQYB
XIc.9]?HJE>40d8=WPF.P,&W-<HAZcQN&R88^;gVWYJEd_I^]Vd>/NY/C]HW1.F@
+E81):eD?B4Z,>#<1UK2Q@.\3D=BgG.=J#1NV,QKeG]1GUBbg;b>ZU2e9c3:TG)2
&ZXg(d)XX?KgQ)=X9La2<5?:9W.UV>NHZQ.I(FLY/6F5\\Ze(/B2SRZ_(.P5c<Y1
H?0O0>LV3#RB44I7S1U.Z3T80fA225@.)E>LbQ</J:DO4^BMcP.U#(W-H3Ob3f^]
SWZ\TP-QIO^)?/;N;J:92PLO.f&7H#WJ9edMVIH9gF0WS]FBBPeNM=Y-fS1[Q^GG
BR5&.&:T+/.?H.OY;85b)PYNDJ^ZY?C9PGHRP=I&E:A19SR2MR/->UY.f-LVGS9.
^c@B<YL06F>]X.gX+-V6?=9N(O&WBYL\>]W(49G=ZbVR_7QcCgXPO#=-3]KB_ERT
fWd5WILaZbES(IM/1GJ2S#ba/AB0TI\V;a/6R#(5^AY:KdKTMeDcHYUdFeYRRVZ[
KGGK0VFW4Rd27(Te=1+_DJ)M?IYDEe+Q]M5M[E)ZP1]-?T_^S>(Ie@?Z##0SMBf(
1^W(4^TFX+U)AZL.&JJM>?QZ>C=,&Q<HdVE.gLO8LWO/CH13@P0S?]G?>R;eF5^&
X_JfeJ&[#<]OTUS2HLRILE\++bJT)OdHW[eF#FJf7?bRPG_+<F=K0bA[-L>2QM#0
E@Y]c[2(#g6#^5,>;&gAL@9cWLL6U]-62#YG^X5;(<=3\E/SVZ><7E)3H8U-2IAO
;;LY=b#6C[((db+Wd-f/cTPH7#MTd7fU3<7d-<8I-OQHL]E2@-];&,C9]Aa_a60f
0QZ@Q0F3R&NBc3TRPPR_RN=M]=LROIJTQOO5f]bB5-7HV-0+K=9[2a]G4.QCfO1^
BDMY=[DLE#Bd0T4S=2Z_GNTgYI^f1OK?D-Ob5S>EUZ+H((L)>WO)&Rd>ccf8B&U^
fEKR73[QcCc?,BYRE7[[7(K[1FB&8I#,3^1fS@g_7M&IIbEB,U(N7NC[<FIG:ZVS
=G&2,e>+57&B8gFc<GL?D.@V@[2>ea((:2DZ#<=.36bebL=\6BC)=0Y#<PId=Mb3
<=,^7)ZFX[@S;O]I7DR3ZR.ND=[FVb0U0U2+B=Y8J_Q98;QS0O)K/1W15AYZQ<Kg
EQ.eHcS_V96gB&(aJf=e.F5NL_<+9,>;G0=_B_;]F<AJ]F5[A,->CM>,f>M5>QD=
CN[+I0:MRf91H\,Z?/WPWVX@BP@F(=2>--0.Vb@+1]SCT4e[dFT[GZ.M#F@(,I.\
agU533CBP/I9HO,QQ9,(5cIe3V994gSN@+\Z)028M6L+1[8P\MBGUUccBL1A)D@X
VKN3)KB=>IN2P:8O+^OL]HU/(<6H?ZQ]M+2L42aCfg@]+EDC?(145GEBCJ6\6d]D
EgDR3OLXO/DCK<<D3Z8VTL;?/7684[GF6AZ#fVb9d2,]7\bZ=<e,X=LeA>(C>bfa
0IU93GX;06,BG0PSDIb,PBY7c,SNd>Y6V?AVL0XcFfD2cdbZZ4;>T2W,^N0<d:<,
5dILa,?SCAfPd4^\Yd+4EC.[^)Od9)<TLYGJK<\@G]-CDN0+T\O,L96gJ4A0B]A\
5/+UCbK_^3XTETa;\/Re.cT>[H0Q34<_#f&a5c7J<:[FN1?f.2D>6I^#28HU5]5I
DX0dGZ=+)gdV7K43X3,HLSCU;[3edO&PMGO_6A_KDc+;\ac=d<,FH&V)d#GcWQ9<
<RVX/.aN45A=,JBL7,L&;cP&R6]6Lda;Qb@SaFgNW&#dg?T^UF&>GYE#5#DS242H
&_)?9)Og#4#Q:_\7XZ^.VS6U5aH<(Vd70]>9KM,(B_HX:R#E4^.B#ND3Zd_ZA^]]
d.f1AKOKQ=:eFS/>Y69P\F)dTA[D.]^?KJQaf+GT;63cIXLOfDKfM1XABa^e?H#R
9?.QdfQa>HU,A;c8c@EAVJL39\KF(bV?,_99[5@G8gQBXTBSYS-V<49US7^+PBJL
5G.4,X?+#EYQA8=(6,>._1J+G-C0bO[:>.1[c/4L:9CBbeBe=eFT[a&ZR+fMHGT+
NfP0[D4Q)aNG:bbT9&NZE3Pdc>58D=4.e]WO#-#H&<d_GUW65H]3TUHb;9ZFCSdL
?E<G>3TESOJa;[V&+?O\IG]UGX)P\6aYSafN,32,,5S;K67U5U,0)I_T87Y<8^Mg
fgA0YfA4(J]JE-EPX0gG6Z^YOe=G0M8bEbWV(\WE4GWA72A\L=1I4\#eE@;7F4\^
Ng&5@IU0WQUGOd>7H,DX[(5QJ8K-_\AVIA,==EI4JX.ZaO]Re;QH.BR8GO<g\O.S
0fR2PE_QCSP6MLN#aF1^E>2&c)+;@_\/c_-d.?1N9Y4WC+Ia[O>L0@e6=^3=_R86
+7C2K=E>U#0eM^CVX:[OZ-1-,<_bS.__N]_[7L]_Z)04bZ4e];D9]bH.f1O5=&.4
Z5#6>#CID?&g#GZ_D?\=da.2F==36+-1K_JN.@<2XI;)XI9K?5RfgSeD_80C?H0D
YH&.9C\C#4(:;>-+fSCMZ@JW(E/Xd&]2:>B:+HWf-b0/a0NAYUQ1R\cd)?9[_ZE6
+X5f5=E0DC,9](Ue_CP-&CED)aSgb4A:]UGB7;6SJNb.Cg>E<K?0E-/>VP=DO&(9
R^-L7(E8LMRP7N^1Q1Cg]/@e7U6])+10fBLc@XA9B^eGIJ2Y\:e>dFgGU>L90Qgc
X&36:LV4?8TT,4U/F^#Ig#aW.PMT@>.8?V;PX2DZ?HITe6:4B6SOHU_+/HE@AKO8
]BQ3+22>(F&3KIDK;eF<7MQ7<H4g@)USb\Vb1M4Jf;0LbF5R18+&-fW7@7]UQO29
<Q6;\3#?3G\F2K=VLEOLEC]LE7\_()\@[fc=TdGQfYERL./L2SdL437[J0F>NJ8H
.ad6_A2JN2.&2<;bOd3=2YVQ>gI..VAbfE-/<DJcT7/:W._>7-9@a7[N=-#XdF,J
.IECgb?836VSSbFa3T0++V10d#Xa32JN&FE,?dWZ?6cNO?A:HcPTf10X<,]c@6V8
&Q?MD[A^9/4Z]__/36Zef_\[U5ZK_#fOO56.ED2@eBaVb#AcJ^6#LY0IPg_WY?\c
SO.d\I6F\0eF(_^4YE6Mg\S022/F(4c<b9+0)Xa;_K\M1=BOUa2b<O2Y#D/EJHVJ
:<;TLA0&24Z&eL.52gQPNg&f7H86?Qd8I\cAJ7^U8fgW5c;.+gG\bQ5P\^/e79KJ
<]=Z@3.0?eT.[=\6+=;THZMR1cFcb69.Hcg>R086/(gYb9NGUDf3YcM=+RIK4;VS
^PD^M3PbV_g+2a[D9LTK2PCOU<G6H?/5-QG\?HBP8RG\2P#BdJ+Z,b05V\<_:?^2
UY&FS/FSJ\2.E#&W9f,?_)13.;HI9\Y7#:3Xa65B6YPU.4eQJa;KedW.=O0LE]Ne
?Q14_@2?L7e(GgI=dHQLG_&REJKfB3AJa[M6W@SIJH<]@Pe]3?2Gcb[ZWLBHV,EU
_g>=\JMN8U(+#\+L=e4S/C8[(Fe>6OFL\dFDWH>-\H8B8(>T)P/+3NRF_@I(7eee
D)g)DPPD&A+8b9R4G7S-2WRR^d5N@0FY\Z]1<I,cR>XI7,=fYX,WO@N\Q7_#S91A
;)NS;L^\2(EV.8A9E\@=RM19,Z;?@=O&g;BEOZ28<97/:d,KN:&1@1FgUQD/02Ke
aT8L<dd0JF?\3__N=V]7._BL(R69Vg)eM\?:N>GJ5OS2)I&]O1SF1,VJec04P.UZ
\be1)/PaH1>gcSM/e_61E6(--.-)O&Z<,b:efYCP@5);7_a[XLJ;L_@&W,].OPT3
9&P[50?+23BRW?4LZM8MGd(^OX^Z)WQe)-J@bT8+9d>-)3)0F[]VI54\e7fJMAIM
=,#-+36,<;@,IO<N0Mb2R)V45MQGZG,B#1BBKWCg>PT<HZ7@J63#;L?5T3:\a9/2
O;KG>#>7f=>PDPe_36#X9GFAcV59XR3e1e/Ob^=?OR#KdEY+]=QL(>eWdad<#H4V
8edZLQY]V3AaV3JO29PO=ANCLNCP0ES0YJ(CF3RS2,I^fGD0@=&>U,E(fRca,=,f
UZA9#&0E>G^AQgY5(R[JG\S3g_RTZO)+dUDE,S7@+cU=[KPJ3f7e<)O[<U2?AYHC
OWMS;6(EDZ3bf.E4e_gIQ4[/\L/Of61NL.GH2;>AK@Q,T]PUYABEe>GO2UbGeF36
UT.C)DAO\EUG\+#eeJXf,H?:EIAa-8L]ZVa4(V9;W[L2@eNRQD7&0]_TdbU2Jd0U
XB#QRb>[#].;bO6[\)/GC:<2_)++?82ODf?I2F2?\4g5^H9.GXC=?aX?>H1S/XQc
.1\SHcN][Ca&?HdZ(:_R.=[^AAPU]H2ZKfR2-71Z=&B8WEM.@OL6MLG\RcL>]TUE
<fBQNCFF]V-O-@aP[+YXI@\a;N.a>U4(/+51(BZEMZgLR;8dQ,=\:15S2ZP,T/Yf
^LDQFe)fIfcO.4\c?FN7g,7(@?L)ROZ5(1fSg;>()H2QBL9&GXf54#(8UR(WagKg
I?>1IBdeJ/+.C7,1XST97Nd4e(.a1,.Zf0Z</B8ffa[/[QIbgRA>Nc+.L>O7MAO5
A?(.CX/:aIKc(-)=BfLI;=,Bd:^Y.(1N2O7)<DeJg?77Ug+/6f-0Z.L^O,)F=TP^
_/7(2,5V73D07b=d];W;\LNf--[^E\/>U<8AH+G;N?Vd<[^QQfR3K11[N(3PRd7)
2ZF7H,AbR)IYgP(bT52-Z2/RP,KLWg&,AB7)-3IBKRHVfIWMfOefB@Y7a0)&,6RE
1eP^BSLP3\/d0XE511(#:7EKb<XOJOL#4K/X)a05bSQQYLMEA)&5d4Ae[61L_VIN
@C8&9cPWU/C1TSDB<AQaF,=.-/7;=[eZ55d5,W<dI>Y2bPV;;W4])PRUSB6O@<E<
O]03\@BLCL/e&LO&C^XO(8MN4Uc9QOKd&H-V.+<>\:H/=^>3][#WH><gfZ&J]?c4
(MNL--H.B/Kf>gG\3^[WIcR?0(=B1;UWJ[c>dPg=NAVZ_E0(M5=#6Y&M,B@=AP^#
eCP08F?JHPcUC6UIT>:)[&6?75eSOI4O8,7)O,FE=QU=HdE8(QKMBef:]=)R#6c\
+S3LUDH;\@P)g4a3RO6O1=4<RW9fU@G8?VYJM:\?K?1aG]&45I0--FK4RL[?7^]E
K1O>5\>:.-M[f23NG8Zgg>EYf]1:^c<+]6.X19DR>/YYNOB/@L=?4P^WE#K)0f=8
?[eLV)CO50^?50L[-4DJ?@EJ9L\N@ffY/Ec;60II/Ca>MFTA)DbNIQa#/.,f.3)]
7(ZN>AWQ@,BE<#E.U&C9&@8.bES(G<>OV9I<@+QeP;7c[E1ggWd;+Z]I-f_7RG5+
DVR3X(>@g>a?+VcQFPPdX^1:b1-?8[>AQ@^,Y\[)feOAVB9E0#55#>Rc;C:,SZ/A
U.T(.^-)F(b]E?6N66ALIJ=PW2L;IA_egX<UPAf#@>T88DKgU+0f2.1.&)-A=LA4
XA[e5XY-IgW4^ULNaSCgHWWC_WB:-,f&HE;.f#fTFKBOXS.92Z&A\>2X]:dYFV(R
:K&AE;&Z5SD/XS@#Y38M:?HcBJ1VW&\54FeaAdRZf@+aQVfT?[B/UK.H7@,?.8^A
3aCP2]Ef<#MV9/OeJD0PDF6]L88dc7_bRfd\5Q_>:[EHTg=>=)P7LOL@V+6^+\:S
bf^,__@PUBK(XDM/WR>G.5\5(9f^QDB11GH?8KbbIRG00R0Q6=@:Mg_V1@@QP.K-
N24<DV3]RBS3G>EO-#[fK<F4]4]/4)JCC2GKAP#X9fZ,T6b?LSQM^LF\_2?F753H
X;X)&2#/=R@Bf9gVQY(b9GOFVaJKGaeFMI&32H-C?dH:d-0T4LD\5ZA]M9VCX?GX
/CA,?JOK59G]ZRW[M9YMZ9d1H2R<Te,@YLcWK-LYSCZFCHZ?D6:6Sf>QdV(;1:Hf
SH>DK])W.(5Y.X1)L]NFdN0BC[J;]4I.X;RJIf;P0@T.^C.\.E1)f4U.PKG2b6@3
#FB^<8P[LR[<\L;DENX8<XPT[g(^&dQE^+I1J[);MDS^>e8HV0@/d5Q+_>O=Rb5K
10aTJ,UBC]GTL;N/=4@0KGJ\=[M>DIaUYa90\GCLR\6KB_(C2D5U:&VW.UR9(P>7
6:;[d[c8CI^:47QNBNgKb:-T=EYM+;2A-DDBMKF+,22<E4<))gK2Z(Z=fdYY8X>U
6V[3;fY)A=]VP_de(_=#/>:O0@:1=aWfAE2)S6bX:)<,e2g2@W8-R^UH09CFd;6f
KTd?)b^\a7SD\1&fL+)c<\g6P=#[O):>a):0,b,N[7_R:#Mf+gZ0Pf[?R2.4;Q5T
6G3VAQ/S,Fb5MH[1G-;AS7FC\Ka1<3H-EHg7YMQ];B]B0B:>[&72L-0I;-0Y)<8F
#8XDRA2&dQBSJJ&YE6^-=?W&I@TXZ<HSPeDRNe:D\QQfGbT;G8>L8GW#,E\8PLS=
L>;U_Z0cL]Z[bU=:eG^=GPT_Y.IQFG0bX/^Gg(\L4>,=@SR6:3AbA^PVWbUQ]6N2
A.;1XbVAMSY7Yea_Z:@J2,V>PE4A1g[==7(,_V<95X/73J;JPRf:-R@6:\[7f=4O
+EY.b()#IJ^Z]H\:U6RGgYQ<aZS)d5(H,L;V5HJ@[&J@ZL[4gff#2=K?US3<RBEM
0QY1D[+McgG)WOe=+)WaL>6D]9.(c,/D?7U&HceJ9;,Cf5.;:MT\ETN[=:db94<.
>8_8#4bOZIJO/#eff#9S3NZ+X.Ac#PUR]b#b&8@>@<\9f3.RK/4PP+P^\g[LELGP
U6f7<SV#O78&37:]1T?9RG6W>X@XP72SRCR1U:/^bcF)2S95_):_)[5UeaU7^VW=
OLR4(fC&(PE/8<EESKNQS&FN?gbG8_K_?>1S;^IPbZQ8]4@SD[cKG@SNaV)QIX<V
BR-B,)KT]ET5;J0R^OW9@J9b\N[^DEbHYZ_R8)(Y:PR=[DX?/(IcQ0A31D7OQ7&I
e<PfU/M?eEG=I,bZ7J60;X(e,_<1U2SBZM=bB4.XE#>9=[M_-S=?\\\f2^ITY@^=
Ge]KC3F<BQW6FFGT+,,fc]a0f_L,S#=0=DTAIce8aU,.7S&&O,b\SDcT3RgJd9<=
[J&4Q&I0[JU^N&3NE@8T,X+EM733[&]B(DP;aA##BEIJ=X0H2S+L;-<7US&O\Q5A
+21N\2.=4=NHaZa80636Iae,IV#PE#cg=.A]7Q9^]:45XZ2&N2<J#ZJQ_;\a<#_L
]M5D^]=Y=6gVf.S)2A4K58)TI@\795_NN?-+)WGUK7RHa1ZG\e]=e,2]5,O>T#@^
2ZNZTKLdSgY)=aGT[K@)W(;[0@S(./8SN(G&@/cFBIag(U;0M>M@YULFP(GKX(::
K/G(dC5G.;UX.<^FEKOe_ZL&:@C<R?F(KLcG7d&H_#P.B_-K;UMJ7DJ/P7-;)0+a
b,#Y7_&f/#\M>R?G?NLE43&><;:9X79eJbF3=/W@S@T@4F[U51&D@FBbZ<McZI8]
8,E0#b@Y-..:D4]?)7gF[9FB6b+^_KRgYS?aKZST/+6@70_9Zgg&.?;_gYN64V_+
ZVdYOY42O,d98a=@8V/P>d;_31+b)c,0H?a8[1==,=2Wb&/BZ,D_7DKL])/CW=cQ
?4PY];XEfeMbNJN^ccK?EZeV3-C,84DCdA3=#.C\X0WGO9EfAUbY<UM=2CQL3?SS
:F27F_@>Q9gA&F9fY;S&-/OH&K/P283b]05[+96T3-0YPPQ?DcWSHK6/#6aX4@?B
=1NNbC(1L-aH8L8VBIgHf>62:&1.DPZ)M:(&_-SZVA:QD[:B6&D(9KOAfbPKF5?8
d(6A&92B]8.(NdXR8Z[S;#.J1Bb_L&Q#TPdc/R8U0)K._Q_cBN<H;+VE-CJaX3D9
&9KaHO@&02C2;FU3cH,4YL]SQ4::^7.d],(d0VC&.2A:U(5V\_3-YD\d,G7KL1A9
N@Q\K>WdaZ5=H8_9f55SLZ30Lff8\1;12,BKM\.]6(c:\P/P/IXbX^d/c4A)[4?_
3T_?S9fE\<D7.=eK4#LQa(dB?R,/ZAN:]Kf=6=OOW;fFfY;0JI4U@GJeY(B>>+9Z
T#KX[MgDX#N^Ee/,R398-R.Y[eCId&CDRTS?(GY(L<CRMN=+2A)K05&<,CNZT9>7
K&W5KS7VR1LQ_R\PGMT\A+Q^VIN54e2BA79KZ/0_R7OeX]/#Gg>;-c(N_cBH4C-)
S64_ORNOK@U^MS1H0fDS6V(&L1<F^YN,TG=]AF>CU/LE4NfIa1TYXE4GBe)cN>;D
/7J>T=PG2]]ZF+8G@=Se8UEc/2NRfL\D^5.e.8:e+:fbRZ)O-@a2<4<R]XUX5D0&
4&OR;W1[bK8MHY<8)a:OSIM9:2H122b<42]6-#?7@6H[UXF9b<EI@Uc1L)J7,V(5
0<SAU^#R)#YM.2X<d<X-D1eKFR&ARM4+QT225Q+D7K^CY#+A3OGLSE3+OfYQKR&@
:9dB83XTF-35IK)e30N99,T[DJHM@\VXST7TQ?GZNW[8cUc8+<a6>W\X96XU6gPc
@34PFd#8BFG;6XZ?_N(fEAQXPX:;I;gG&=JGdE^N9CfTM[3U>XTI+0\NaTa&cWOe
8QU2H;545VHbJO23NYGE<a>H3#FL<)[=F8fH?[c=ATT<TA(M;/U,<>7Y>AS\&EFR
@DAHJ.?:ce_6RM5Ic\AT=^04&AC4I@72O^+&ED\)^K(GH#/dg.JT@V7:6a;0a/UK
D;A.0f-H9?ZI_PQEV)IM,<9@VZ/QM9cKc3b]b>N+6@?>>>5E<NbXCZd>7c-?,ZeH
]@-#_3GVd16c8>@FL8RcNTR9E0aQ)_UII<U\>JY9<f+BC.E0Dab=cc-c+gG^7QA;
16RdLO7[eD:DEZKd#(.H;/Q_;\g(+HV/L<(eR2C@2UG<79#>_\3AgS2@XD7)eB\a
CCW]6FUNB;;)(JCb[Q^>.LBN_C8?VcHQD9?7&0d98gZCf9E192X&<>B62;=c9GX[
,Cf=&U&7I]7V,#?PZ=c?L]?=A,Na/:FAH29V@30FI/c_-HZ&N3-8J=;e\Ke<ICP/
X/[1>D<7J]eZP)DW(.cg62074BGR[R.:>;<@KYJJXH_QMRN6J-&bJ]C8+S4CU990
#FZC7bEKHORC+8EUEJQW:d<\(f>32SLRf600SI)g3S(&Ec,=R)D6#(YF]ZP6-C,T
>CAc8af3gQEd(KO\4_Y86=cV^@d(U>,aJA>XLQ6H;>[2]HWd+_+E@=4B7M)SRdR)
EQD/_[8K-TJ(C??CUaa8Tcg]d)-B@+T<egPf4VJQ260SaWVYC,P0YIA47]7Sc9J]
E?J^-HcS\PS#P].)0PW@b@,e2/a=-3D>4c]bP10EFQS>UCX,R0>N_(^(TEK\-Q;g
<eH_(N4RgC:H,4=]S]TCM9[IA,W1LZT?DgUM,E^[(K37SdbXE44@3c4H=GQ]-g99
Y3Hfe@\SMdFFKO-R]b@2PZD^XY[+3EgTg4c<&^g)J?g+,8I]F_LTVD_(RITM:.B^
0@NDH>M-\\Z)EYYDGf(PKJ;MQ#aO769<-/[R65U2&X67-Q<4Vgg(Yc&-UKUdOHDF
<H,dQEg_?N&eS-=AYGIDV#3MFM-7@J2K?O3/U(-b.fg9IMR^YeE<4>,NEBd0.VYQ
[G0=cIW]-eaJ=4GEG60I0RgCZHT(4L7_T9U)9>)48(QECdX7_9?#\=HE0,E560J&
]ae^J^b9)FXf0<S-\1O<QfTcMDeW1.gB0AB5bZ53HL9_4;UEKBf>@RfQL/&cgZ0C
9S=PM<T8U)K]/f=caAL40]WHE;2@3Z=KOHT[5^028P><_241KB(GV0+b,U-eW(WH
@:,HF6+g(PD96.[?(5REfOWA2?,@C7O4_)C#JA//\QeF,MMgM:2E[7Q1-)@ILOKM
/2L:Pe\R]U.cHR,RX6.3gGTJ5I\2QS24Z35\5X=\H&NP2V)4F8U.@>EYZL,AMH_F
dW5cE3AM=<f?>IVXT)I1.0T#+<5b7MBU64/OT@(4V<\9@0I7]HXLD0RfO)(^T/BH
<_A33A(H@aE<C1E+U;VE5G\MMIH^PS3BQ3+=R(C5@^#^_SR\X4[3/][H?TAX370F
Q9gKM&1Qg,_]A)R/c)L>FF;d2>b6;Q]=<YN)Z4K]22N;_@6HgbDT66P&91CW6=6Q
(&P:BXb)M9RRBg^HUP+;Y>_6484U3Q:-@_NDe)U4Z&d^S(D.&XYYeLG3c&&+5WB=
^D]K^D&8&c(0-dGO05;XIaTRDYAO/d95_N0G8dNFaYTc<W_,L8.3(DT]P6U,+&M1
&]3/(TdJ2)2+?;VU0R]GS^7-.agGXdQeZ1fQ4W8O4.MggeR^SJF7(GHI3J?GGLOH
<BDN:L0IdIN8\fRR#5@PS/D69fMa:OV\;K5dU?b(8=[/XFPd)MBEZ]32C&=S\@E\
N134A[?#C?DIA[3a8aP=,N^@GDZRX4a8:LFM?>EL7@2c1K>M19Wa]LLH4dAX]d,;
N+c28(&Je?4_)8S/#\X<12BM8V(LC_R3;Z;4BFbJa79Y7=43LET(V[fH3/#eS9@I
NHH]D74_bHP+b#L5.>Xg9Gf@J.G1FC(<R)7\::M>_:[>)5;])M.@A0XGFKT+[[^Z
W._CN8P<ZCGA;,=LY[H[OT5+P;/E[:8I6GVW/Jd\BN7eeg5&LJYA#49(35TeXK#(
E&B\9G?>LGSD[M_G[4ILEgFXTS4+_H96A>&^(U:#49L7(LfZVYZC>cP=8g=(4b&:
R9R-=a59BXSNFT\FE#,HUS28D)dbM5Z_=X6(>#UENW516PO;,/Q/PFQKF^/\B6TY
&>HMYJ\WS9#X/@__fX63-+eF(W/K/1W71,cXIX]B]R0:7HQ8OOR1D<RR7.N,B0+g
H1JZM6JR?cX^^3Y8K#^&G(af[<+)g;:?DS^1:^\PB&+L.[]:,XP]f]aB0JN@R6[1
8[>P&V_JCHOEdCT7Z<-)Q<4bL(>XL--,UR6gUa^6Z-^E.CHT?,VF@_;?QZFQ#<Q[
@\O1F,fJ;;/eSO&&e+TR>Xc\aRLEGPBYOG/,T<ARbZeP4+bY:AQc7PI+3:2b&EUc
+I+6IXKJB-:SVPBIXCULQU8D6/NDa;6BU3Hd^UXEKSF-TbW=V70@_D6R7H]9=faN
\M@ab8YgZ5A6Q4Z3O+\fB?DC@^2)OI_XZU>H??edc6Q.8c<&[gT703,N3RgA&J1(
[E]=\?g1aNe<_R0);aPc)(SSP>geeRN=AM3f;UZ7d4&d-OU2)T+57f&]WH1YC?cG
Z-<(I58DP+K>VIR-<XF;;V7FJ#XKKb#(-X.#W[B?aQ9+=B#U3C8^^/>+?Ng+/JYf
S0]4eR68S#eN4OMF5XR^7I0&F[?_fd,;6S1-[B>b29;RXOR-V)I?Y+3;-F[gPT0D
\1B>fKceZBT\J03QCL47VbK4O_XaE48?WB:?S@JN?FX^XYT,B+U>IYU8c#KPK&W&
+JN\8c^f96Y0QS>TO>aJ(6VO[C8U&Q@2bZJbfRPEB:4_ATBM@2#b?L.:Fg2Y]-#_
MdM&8BFXFXQc?Ec:==d</Of.Pg?2:D^D/-V\A#I:9:1=:=&Af1ZG5-M3A:+\(..O
EF4Vd>6JN9b_>8,W@/?_<6L\1<+La]R,20,[JM-Dd6_E\.\:\RBF[6FJW^WGObU@
f[4W?;W)A=IZ?V?+A6B8#)#Bd9d8F#3aT@AcTF</;J8MfRHMb#d&UDP@H&^?MV4B
;L2+T+DDHeJ.?<-YU8IRAAN3dNO:dcS<_F-+PRb&@Q_<&ZE(XU26W(><4.63gb9b
S\XYSZd#a1F.F^-E8fW-<J1,S289XNO=A8X#OX(PJ(T8,.S\c;Af,;@9V^,2GZE;
/K\;:S6:A>GgNe[1a_c:D1&#CdI5(3g&7:/P+1ZA5REMX,_01cb;CR9d9(+&eR3g
UPYe\K)QWB4]GGdXV?P\NTNU-KYOB(E<,]?(P#S5;Q)P)&2LC/:(/.,Y>_JDbYSX
S<g?eCQb8b/J8Ked[.R5>\BbdA^A@(]BTa^GQF@IH1@F2c_0@e6=LZYgaefO1\E,
^RbX4JQ[@U81DJZ.(W3&ae/-Pc8A+FIVDL+F<N\Uc\IV97VOXGIHNQ^/#5KWOCFA
]):\GPXOWNY?2(H4AKXT#D5R4Ne(SS:0^&[JP^T@89WR@NRNc\AfAaVM_-T\aFWd
/PWIF0<Z:dL/H32:HJR(QOIGf47DRV5-_bgDgY9fX0(Q&4&e\2[48a.?HOW[(U67
^TH64&HA>M@HSKa7gV,1=(4MVT(4:O;\J@F(O56XYXF3@/X0YCaE3DJ#(+G3X?PW
SFdQg)P9])=A?@\cgJcK?NH/dFA75SJ:3BfW/^XLT\R#Vd4/V081f;/BY(7OVKK[
f[=D+TegWf:SZ(UKB5bKb6:P<^2JN_e/OF.NBE(LGR(24(</?I56]:B8G59V_:@V
3YaNd[FO(C\+_MRMG:K:&BQ-FD;VFQWWFZId7[Q8.VIF:+W;O;.HG-S&\S9C#(dD
@VO6T\A7Eb^g[QLIeI-,45/Tg?U8YEg\A?SeP>RJA:HJQDA6cBS_bg7YVE;.6S@N
BW7M#J,9I;XgFOKNZ1f78V4/0Y[G#IG=UUP3(f+3(PHY/8UaUY9:[6dLKEZV@2Y2
UU2+RA5XO;FYfU0c598TNeH=NTb.2:d@[ME^dc4AH.&(J07,),N9,A,>-(YRb+M.
dddE:<CW5NW42Y/0ZT&LJ;U,Ue2N6f,,K4K4;ZG2-BT@1ELb@DCUIF,;_+6)&S@d
,d0&>E<F0GK=?&VZ>YQ9:2W,=V&DLYeYJ=FF[[g^+>UB2<>[N0)W(Cc,M;GKJ=CV
I<R5ZSg+LV;e:F8ZB[a13^X[7^18::4UY8D<f_c.J#+e01ZFR&?#dH?NJ,SKRafH
=2.[_GX8QWZd39ZC?RXDME?R)O7L^gYJ97^d^/Q\L\[I]_:DMd_;&^W3ZY3F(Z[^
JVMg[R\X=SR:gQIS-F3;Y.F/NGU8QcFZf[J<<1>U;X_@+Zc0c9gLK:2\_SP<CE&e
AcBU?>Za&YAF4aU2eL&OQ7)5>U2PUAM5Z>>[/CV;?J)d]C4A0,P/aDVH]dJgdLWZ
1&)X3=WB:YUT^bQE0NVc7c.5B)1K4.c;bKYBD<:M/WKfL#/Kf(=<BbTWJ^))Ff:0
AJaZJY.5bIVc&5,_(>YY84R#?+e/1Dc?S2#CaAR:.]>#e?FD.NI\?T(VN:=OUc=<
&YTG/B[38[]G>-)V#4RXc;#[+657d@00f=QSb&#2M0JQ;&_Z#G1W1[dKg9_)Vfc?
(0TZ1_L<@4C+==ZA0ZB>\KYF+/L#(cg5,0J@YH>-VbCe<7T^#9IWE3>[87(d-7(\
IDEE7eDcM4KA5aC:[A;\WVT#23LLTY:^MFSE7G[bK6Hb3UAa.fOO1@.NCQO-ggY8
^f^gA.J5C.XXb/@5@5c(_;4.Ga381e:SZf1-IH9G7V;A+.:.SZ;b;/c@V_[?:T=S
1dJR4N^TdG\G._#eW)0[L7<.BF71GSB2AI&aH+AF5LFa>6f=;0)Ud?4Rd7(,=FSZ
.\f4(QTJ9I:g82E/B4be7YL:<^=Yb8^gNH]P[A^:E5>D#ETHWN4>a=g(T6UHS&+J
PO0P?eX_FUPUaJ>Z3,:0QLXMgRBWeSNJYI=./^b=ge5.E/ZD.E]F+d4H?PW<B,@#
@a/e-L.-g78Qe[0OL\U--PPDF1,SJ,Pee?GD)\+EC?#7C,aY,cc#/QHa:bROQ2H3
JcHE>(/0T]L8]9/Gb4W:ZJ7K)dUKF2P4^a6(bNFCY1(,LEC@4^=J_FW\A;ED40-:
ddIY9>C&&16.-F0^KQI<2FdP2#1C>+7+Ba&@d\VIb+35TO(Ta==U-67-AEc;B[U\
18O@Z):+,8G,J.^FZR\b9B119Udg1NbFD@XA.T6)(&dK2K.g<U8&T6[e=TZ@/<)Y
8SR?eK(/>;#7\C\TVY/N>EM>VaMS#MF?^)Ufg;[_c-\I#ZF_<bWWPY(Y)YeD7R(J
a&8[AABJI@A042W5Y-bbDKbP.(0T0^([RG]=YJE/P8.R0>QTVV:.aSKc:X@dW;Zb
Fb_TZ,EP.bC)YOIJ_/HAd4HO+#3Fb.OZI0RF#gb92:R.A2<X1f.CB;g5DP2WCec_
K29X1[-NF-U1CB]J=;YLNg)C_&W<f_D+QWY=SWZd08Yb\TCSO?ce:PHCHNR0_>:N
7]c3JN<^?YKD/9ED:g.7YYC.C#SOJSb@CZEG?T)7c6gX8K<ZC+MZ8gWXC\Na3H\G
+.D\K;W/;fBAUB=Fd=VSGV6:?OIcIgDG[fZ4SFge6d-c8bT)2&P&+g2)+]ZWU7\G
SMH@_-^fMJ(.H&0=TBR=N4R@O:(HJC03ZHB10_:^X;^F_&=:Va8J^\?XDFDa:8g#
N)R<We7,NYL:<b.?#gB@YcbcKfCdNeZgfTNF9@:OUgd7b:b[gK.J4#2):&;T?7L2
\N80,.&&C(LO<cT1V?N<J3RKcW7Ab35DZ^egYc-WR>51b=O=UaQD0\:&V^dN(Dac
&/S,//&a_4D.SbL;R=L]-O)MD,5L&Gbd#S6/?=[aME^M?9N33<7U<1f;<gG30MUQ
,;\ZB>X:<7e2f(XJ20L3.-B(U&c9_=B6f,#I=]ZLLV4CC4]f^fBe8[Z^:&GVf^]E
fYJab3@#6&]1XRLB-aLD:8bFafeVYF>,Y@S6Z/\JaP#^[a.XLU+R1D8e??/UBP[_
K-<6/E.7ed7f7MdDZ+Q\d^&I9#?\IOT40E6@<(-Yb>=5AbPF7M+QGY_LQY\64N@/
>NV8++0C7R\5TA6.9ATR.YPgI7I^@M[@KF:X^B3JUc\5\U)ZV7f;P,g#KWdg&TK0
Q.6O62a_N]=[477L^40K?LA7(Y6MKc4J20JDSeA_=-A6[U(MTU#3M=4YOc]]899C
+L52\@J\3D[-1LLU1F=UID5+YL4a:CH\aQc7M0^8,d\HT;]8-XfSeU/9[9@cg6V.
9T>@?1>UW3H1EV0VPD&bVba/V4:[_R2^EJDACgR2^a2>;gX>1G&fT=[PaIf=DG]F
3ON/WZ@8a,0L-(BV[1)0Ea1=(N44:,W;G+V:.0W67@7#\N=LR+X0,^QJM\P9aH;K
7-)8WN5+D;b,=Q@ZJPTQb154R7V>O?2-?.4TBFBZSQN?7P4@JK&76>ZQR7I\3d3d
UPBb\+D2DU/.WQ&#0ZW;I@11,fQU[MU?EB_.1\67JCPT\(7VHAX_Qca4)KH]#&>[
.B1TH]AL.M>[b(^FOYRfC\@7K](60YS81&59Z]?0N1IA7C9Q358^JRbG=d:K6ca#
6E]U;4A/[V3J2gTT#e0FT(=6:Q<1Dd3/BM3dX>CDSY7Nac=>=AdfR0@);]_6@+@&
bG]XK-aEgYT&D?Q5&N3^MfL/,[>\b&LP748:3_e:C2#4EM[K^_LKT8@Z26<1XVZd
3-UV9;47\OO)^]]f?b9=.#0:\4V3#_[^b8XZQ6KW41#K+G2,M721gU<-TF17UVFe
d0H(Jc5TIc42MBCWcWZ;^]0GY8<)F.#MBA.Y3Z@)VM\;HHB[)_+4Qf)DA11_c=#<
[EgZUHXB^HXVe9d4CF51NVPgG\Vb=H@<.>Ge&SfW]^J:NeB3R^W_C_\1Y;\b5f?=
KeG+:)&7)B+dCE8K6bFU=1cL)KGW\c9LcTZ/K;>cUTNA&J;Ha@c1>)CR,bFg,B^H
=g[S?17bXZ>W1N_5eO3DBb;[4=.b^c0,8e]4HRg:\(82U0H=E/V<9QdFOCDbO5<X
;-a99WeL-]^U<B<LZ#-;,J/F-(8Y<.KFU_K@fY/C4BcWW0=28P+(Ebb5T>OH7R.d
NUgZQb#W6H::6U.[Fe9=P)W,b_Y&2LA8&S#/N_TJ]#YDM1C(f0IQeMY,QE&[,U0B
W]c_,79BMcAXJ#KL/06<,WaWEG?C@6e]cVdJ@F\&(]XOT>B784VeJ#9afN;QS\a(
[1)B?Y]LA0Je92P5=,XCaeO,WE99BO=:f1Zd9KK9XN:V4QE933+-T#B/U8[T<YS+
M=39_AJOV#Ma7>Y#UaAYBa6aN:FgUXd:G/Ce0c5&[^^FG3#gQJQJbFP5>:>\]RMK
,V7g3aX&H,^fVHb6[=ddc:?)^?:Y8H&Z(-T4.\R09GPP0VgX4U57GfSWEOdZG>1:
CDW1&FW8W<^W1F1L(3X1(d>4ObO@-H8&Z2>T,N.V;6&_C5JSG;&X-1Cgb<IDRA<=
7fJGA/c+QCEHJB/2^>7TdL;52-&bdFWQC[0ZI1VA&S(7[Hc4W(/TXK+:2?;^8/V]
EG-@5-D)F:g39NM\EQ:AVI6f1ML/:5XP1&(E6>@@LV4Oe:Y74gb:\K5&N8L_Q_(]
bWUF_LSW08F+-?RgbUP]bX)SHY00&]C<1B])_V,.YaeZbZO-TaFO\.\@&VWK9LQA
>K(?IN4LaT;^-8-NZedg+:La3g>46^]TF^TOB@Y4BWJ5(M(3>f#7HZM0[@+A[3+V
MEP(JD>1XNPXB9(<:Y^;P^[VOKT<da[fO)<Oe+O87c,fa4Q_SbED&^7Z3Wb--Q,>
@-4M(H[_2HH?+CWQS6g\S?-V.6QKG@N]3a23bUgUV_;@4DD8a3UVEQc^8?IZS@Kf
f;I6?5Z>/C.D4<K(dgN.dC^E]PNLEVJ=XC.[?2299AJ8X_-GIYEdV8fa#UH#QCGg
b&>&F_C1P\BIT<IYEUAGO-L<5HBSU5:a,-[d?c#QTXZ#-:&DF5YdCC[_:][c<2/b
\/1g\@<#WcGRTZV3f6T#RCETYaY&Q5MFb)3(0ZfEKMN@9[U,.PeTgOg^fBNO&VPO
/AW?T_ZW-];a+8,aLHO;b9NKO=7@7R,fU<Eg1L?#:1KG6BRE,_1BR6;d8XedB9(0
6310^0e3].I^>=e=Uc80Cg3a73f_FH0+:]3AZ>WG/]7/g&BUaI>>?,W2O\^Q.4#;
4G9C,fMH1(7D3E+>X<->?]@dZbT(QUGTJdcR<XS13Q&MF7TB-(ZW;NA3Z:C?OgP.
3WKfU@0@.K]-9L7=[(^P@IK5J/XI6WCGfM6JRQgd1F=@90KO^YOXg,&Ad@HSVc;-
KJ82LL<ddg[H,V&2a(;I/J5L/K<W8&QaY)QLX+a1O.dE.W?6^g5N3_47[FT[RLU7
>TY7Yf#E7f@8/b8^8.P+ZPJIW6H0fbG:BR>V1_&^VcI=Vd;0-Xa/;LW:Nc#I(N@&
b(R)_+_&dZT;SZaVf0BYa)^+d>X;Ff&Ncb=WGY>2:;44R5<[BfECCb^T7+C4V,DP
H0JT^GGgD8;>]/eXgV)S/=VW&BM?1a,SBQKPYZ6THW(I4WKP42eQY=P<dKB>9N5N
DZWA_HI/_@8gKOF/I-WMZ@\U<^S+1[L?0a.;a0?NaL-+_)PYc)=JL&B@<KUFNE4J
GWE_YY8:3AWG16eJ_M]EJJJ]c]2,_[X[ML;)Udb5efe)DK0H]gU,V-WM<H-_\@aQ
65e4H=SXS3GQVL+?MOVN5/>Q^7cQM40Q;cdXDH]Mce-[>OVcCe]Of\d<L,@^E0M9
&TQI96G:?:5SaXg7;0\>IQf\HJDIBQ>cDS+Za]4g;?4WDXLUKKCW<IG1_7(#8@Y1
JNT>-dOC1U8#R9IKb4JgcZg12:aa^aXd\7aOO,D:\=((e@9/,e)6I9L5^PZ&D51P
U)F=[1=EdF+P3CWEgZFDDPcE5d(dg-=PIGF?#Ce?D<T-a]=-H223b:,\\T9_bB=.
8gEeP?JPFg,.457[717-ND&V&@X;>)fe5dLebEEY4#8(f2S9A9,TYfM[^I,TV1AI
X&O/7FFQ]]SK\VO;\:\2Q]3MN6W9RX_a0=b-5MgFBSVUXV51YR>fO])N><Z]J?.:
2#[P2?:^8,^PJD]3>;(_cB5L/O0SHb+5COfge(FOW<A[D>,817OTZWaY8f3fRRRD
YF1K;XX6JC68V;&6a?)2QG^)MG5b6EZ3#UN=P+I/[dfU(-CCY7=V672>TI<S;O1a
g))SHO@FR<XG68a\dFMDb(MGR^)#AgX56SLVbB=0AR.D=_Z60SHDIKSbBJfA2QG]
8,_6<3#2Ja&Z(3;U6\]U:6bK[]I-GNXfg5)Gd,LIfcE0H,fOHV[08E1_OUYaMV_D
6CDcO?\5.V@QU<(1(_=M>cM0Og6cOXG3_(ZTaeFN#80eNWC-VQ7G5@9AU(9<FGFD
c6c_M<g94P,g34Xb6=;1^-gY>I1V[,e@0L,(64fR(WYB<?c5Y[N,,PKPdE:EYO_O
YY3B=]WU?g+)@.4gcfE3VU:.BHeZgZ1Ad;8/d2&V]aVYHS@XF5(GB#g>^XBg<K5D
]dHR=ML6Iff5F4Y?U=d,e4BJLHfLPYa:2d>6dWYM#:.0R-TL(W&CXOLKFZ_8+E[S
Y@-.U@RSb2gBb,bb_/9cZ]4d+CX\Bd=DDf4N0\<BZ+ONQe\P1S/MX3K;+6I\G=<C
@Y^1?B0FL=>2H1?NSXc=L([a(6dXTL.H7T82_fG7:[4+?>A[C4>W9@(<0O#Z8G&f
VbB/gCcSNL-d]Y,@QW,K]WCeYX0b8;)^P,K9)88)KTD:GQ50,>[O05d>\/=JZ:99
GX)/DNOW\f&=^a;J]Wb?+).=E]GbO6K.]<UE+HQ[1DJg):bf#8-L=TDFGWP6fO^P
7fA/-0KXQPVP&1?GG^L<<<QUVB0_#aN)GO_<&6KC14MTP\,,FD>#g<4@3_XJ?dGR
(a4e2A022S5OF_9;^O0-X2R/GCYXd<2C0gLf;(dB7H;41aQHHFJOU0F3>aEZ8+[V
cR#eF,D&HdTZC)O]>T9S3T-Z+JgN^N3G3L7O81;aMb#e90C)+41N#ZP_T9S79c7a
782R)FZ-T(.T):43/)DYU1Of=R9C&Z<.bUTR.D^IJdYK<cJ6+/_#8X5gJ-8FNQ2C
?5RPR=US?8(>bJE>5R;;fFCLHV\<g_FaHe-0+7:?SF9@&LX7D3Bfa-.)^.+T&3DW
^F]0g&TG=gX)Q?>9bT]QG6e+dL#^)_aO7I=T?AFI;KO[ffH;;D==B;A=Y3b?H?Qf
Wg^F:3;R.WF0,UaM77=6H0LMRO,5H2Y3XC^N=M>eR#98Q^H5NBK-A43L9.IPb^FX
BN7<M_KG65Q-bZ<\&?dR+H2E8G.-]A7_Z1IT@2A6+-P-9=OLIK[&1UTS+8H?9fEN
g9_V3D+WW-BfFP4W0QFX[dI6bA@aB4Z\I>c(cYB]I^<2ge@^370X[RR))/Jd?M45
4@d;M&\W_)EF,@R&BF9P&2MQ1=bT_>BH>O(#(89^OVc8S&<XXe;SL_\+91WASGVb
V4f\XDC;NJMA+2TO8X2](TM5S7_[<,M+J,gE,c,cA^2Q\7VL)bf=>4a;cYXQ/8fS
H;UIW34V&fJNV5RL9DEgNf?EF)U\bGLE?KA\8V_6(Vd;cOPRQO.?5FLDdeP3PaCN
Jf^#CgCg7XDBdZe,S--ZP=<9NBaJKN.D[5AaZY/^1EaB29STO,bL:;DHZ1JY;4a6
S)b,YADP&6>8gWF^&UAR5@I[\KN^3B,SXa;.V(d6>?(cbb=(PQ6\)UJS8-S/QQDe
+_UdMOg6C1YBEB(CK_&QS&?:c-X?LC\X6,EA3/036KRK18OKPe7)H+a>@U9:(_.3
<-/85TRK-TKd1Q12@P&8-Fa)?YbTaP20V&S^8gIcM-:U\<4)^VR.DU-0K-)d^E?,
b)@fW.)Z;Pd=S@>>9Q.-1,T[+/=G8E-&gg/#cU6TTcU]fad/X)&\CH1S/.T??B7D
-2VeF462P3_)LTS^U_AM[-fV9YJ.>c^FQ3QbSbQ?<=>JXSA>3COfYAM-bb=Hg>ZZ
?eJ)e-^-IPafY^K#:fPAeAA<2V]:6?P8)@&^RBK)K_-V_2:RF1,b-ReQPXBb;8,G
4BJ1,+&22CeL59f;SDg,@QP64=;dTVd/:d.Q&e:33=S)@cF-V^V-(\N:&&9P&<g.
;1[@XQ6gKM37Zg])6-gA)aSecg:#_[(J2V#01AA0b2C4S+=7&\FVF]a427-eK>4?
QCL]5Fd3J6^5@8e]b)[NP_Od]F7GAQW,P7[?6I2N)],,,.YXB],=Ra\\1?7Q@;:Z
.D;CeJcg>^+NK]8@5JCaAQZL#;D2I:UIL#HV72\M+aE4UU>;64GJ7D0+TP;^Qb=+
65BQINa4^AM3.4bZeg3Q6N2^a/9c58HQ:EJb5A>aHfbb[Y?JH^<5X>GObBAX/I&J
@U(;VYNZF:egD;.J8A.gVR6[O)K^Gf4W<?\HA8Pd\Y1Y++d5IEHc7RB?cQ5c,,6K
ARM@Y+fDgJg9IRG]OW36UCK]#=A:E\1;FV<U@<7T?=E;1cTQ\)b])YC9I;La?3W4
UT\Ff1dL\Ga_L;8fD,KNMdTRNXBT:;6W,?e3Q53\:?JKEOD1/J4b_/UYPd)DW:8f
NfbfDB=]1&Bb>W,:WcZ__d7@9W+-a:Nb:]f7e7TN6Uc/3[)1aZ.]c[A@/&=Z<Oa<
e7YAJY]1V0MCTIOX8#4fBCe:]RWQ_M:762<2I@>U@c4O2&#X/Z5@YFO[LC92OMRX
1@#;(A:\K>D)D;?+ISbBJ6bBDSL299a/X_G]\W?MH5M?BDb63E<>F&fRXZWKH2Of
AaQARWNef/;gXK#?JE8bF+3-OcTDa5&2>#bDa=>@b2#IVg.48?;4@8L5_U^H<b5V
37aDKE?aJ45C.U@bc.Gf?EWODW)82PX2^c#^O9+>9W-@X?\Lb5Xc^#Y(?eF2>Q80
BDR\#_+/\)&?RJ/+a[5N(9M>[1cX/B\?LU#43?R#_U)Sd3Ned(YZ^-[cQZT4;7fJ
A6BRCPNeJ^5ADMM,C,8\SDM#75/=_O4N?:Z1e@cb7IWc+c6:7E;^BZ&2[&=X6GE3
XaEVPCfQ2.-GU?Cgfd[+^05GFJ3F]cJ:7eI9RR1-^BQU/Q&PVG?gEFe9@M8:6FE>
06UKG;B?#8OCS/[NIL6@W897>U1.X[_2M2cT>f@AdgJ#c]AFRWMUb[4HVEN0gf9Y
^&.N#N,W^];<]QY4J(:;ZH8eE\b0<J53c9?W=A:gcF5@+dI,_cSP@f\6M7-a#<S=
-3QeJL66K3&&>)DG#;BTMRgB[9R[QFNbQCRV4R;?YRB)@0A1(Qad];ecab^23NN/
?09XO=AD>_;RIXJ@-OaZbU3G@(6bc#,b_89f^d1V85SQ68Kd/E^;]#1/MSbaF_0&
E=>GgWSHK,?VcGIC]2IZG9C]&HMY7R/P3I,,Mg^TE;dRH?B-),JBQ9EWT]Cfb3Y2
2OI9P(5R,T6@)Hf-aa5-a)?;7,3ce3:#2DA9F9G@Vfa2_##0/E?2+(d():=WbFa-
[^<fRb:>Q<XLG4Q7S#d(FNT/C@HG7cL16TIM&/;,J1@=01fB__FE#HKR9+__IgTe
\,2\a&>Ue5.R@S5+HSbTE5&M9EUY2JJeS&_ONd=IV0NP;P(C_RCa6@3cV]fYX,Ae
WXB&<Gb)aU?b<FbN3a8R2Yf)Z,..)/b:cCA[W)2cgf2e)O6.7ZH./ZeRf:3ObY,6
\;^C?S8g^b.1-Qf_#[S3S/ecgf8BI]91FI:Z=KPT@NJ0,RAHOK,#Ce1042Sg73TF
?AS7QH]6cXV5:W\P5_=Q#Vd@6D9@X[.35G/@__W4H/;.Rc>0EBN,b-ZLY,:<VQ2&
dbQ_IN&FA(#Ka.dR^@10Y,T7P:Wd21XMSfcM(^0;ZQ0K9ge1O^-Jb[]L\c?<PKfZ
ee4D#/=8^NJ<JJ&2<MIE#M6Z>D7B+c[7eP^[0,#)K;\:AHJ,&-CC&&E=K,\^=XO=
3?BI;AJ4G<#5F(6J[,LIGJfF]24c<&S],OJRIR-5BQ?5ML5))X]+FE+bKWV5)+;b
;_db58_/#Ic)a84?J_KCWTV:1J6S:-X?/K7[LZM;:/9[OOCKYZS]1LV1_.bWI@30
TW-V@G631WNWAF,,/\Pc=T(ID56IS,FA^B&M-BU&=4R)f5ad+VdH&Md1#&K)8U?#
YMU?R@>K^//57+(Q4UHIF]N+O&Ja10T3K071F)55V0YB^W)#8X.SY.#Bf;1H3(AV
>RB.a:R6Zb5TKZ#CX<cK3OY/dS5[aVRa5.O&YMIGD&8>;B50YaNE33.,fSB/TdR+
1I5C._dD4D#A@Q-GcBS36@3#NP+)Z#f\8EAS?/45F.3:.K[G8-R;;@Mde]CT/c\Y
).9E_\.NJa4#F>2D)#5..R&F#P(V:4gcB\_1?6[^D^>+DJJa>cNG6T9\IBWZW6V2
]ZH?RdI7b=@f#(.2R<NTB#BIICSBZ]W\/OZA7<b[Z?WT[H87(f#=JNZPEa_XYN8Q
#HCTCfAg@ZVS6/CK&S+KTZ7JMJZPdW2GF^ORIN0I45M/>Y(;4VU3JKA7,.L]_])9
ddEBIWP99@\f18INU8G(V)I/O\&ICALP80&L9)]Of/HAf.6_QHZ-de@QGXYMBF-?
39FRN.6&HKV]DV)/:=@8<LD7TN6Z3>1\_C(fgPaCFbI>^=8R:RZW)_;]UOECabV>
P@:g43OSfRP:Qb7W;[Z<dQ1M^0@3WM3@9\97fYC9+Z]aTTXI+)LYI0MJf=c4U@7P
=GH><QDPPG.A1G&Nf@7gYGIHCD&0&)+8.A?Y8(VIcb>;<W,d5FgM9e@ZWfK[=aa)
O+?X-/MRaKQ:=2#V=<ZROaFc@;Ad/S+?C<77ROL.@FJ0VXT7#NCSY>6NRa5<-7Q@
565\OcUCK\VNc#B=L@CA1Gf][-;0REfGYR.Y:cNUSKU9IZ+[_G]Lf,.IV+:ZZ]7R
[S3GcSRXb<)55D^DN;_M3V(I+Q4BaVd^E@5);]>++<#/+42c,M9;8K)#aP@E06Y_
\_/GF#>/C)9T35;NR#Ib7::b9ZA-W+S)-V;MFV\Z-.M(?:WOZSbL&]9A0^[e?FaW
A4J+]PGXg4;+BPJZ)\e<eaQ5;IdU/DOa:.eXCG_a6XYH)RW)BUg3RJP/T.c<F\6R
B?d>>HgL/;H:;4cf)@IJBJ+64ZTE-T/8XOb&=L)3ccOMI-c9,K@f_>[QNCM:75.(
Bcb;f8[]@\+5@C_1NK6II&\:4_F##b)_B;?B[gJ#\CeO_KR1CfP63W6X7\RCX=F-
NVUI[V^Oa4UJIFe=U+J/+b+H8fBe5NF/I?BPR<4O^LJZ7GN\PSe([NeEc2f4)F2\
dJCb0T(,(P@XSb+-<E&;N[eYNCE;W1@a\cEZWX(3RTJ\+9&XBFRAPWeFFaM0TSOA
)3KBd._[[7X4R?17S[19;B3c.YD+_9(:IY\K:Z9O^c[KM:D\cI#HN8PR(gcPH^I_
U(S@19^/H#WKHKfU7KR1QH;0C:7ZP_fH/L>+LZ#cO(TC9ETMaZ&)G[=SLEL=#2Da
T@A0gA4UA@:/=OBg/e..]e+7J>WQf?V?&dN(N,<YLAS[0cLC:\H03aYG/J:7)K(U
f3J]H?MMf4DP)>1P>?#;1Y7B<P7Y=2D[>7>0J1S(a#AT2ZC43.:I:QXa=_-/cG4Y
9d)[6TV_\)SWZQ\R@S6NOGO#]4M.MBZ2;1fX;(P=);f9XI48dPD6CeV@A.C=-2&H
(3abP2I3Y#QI?\,^QPVcG9-HGg\ZEG;?<eDJ9>OIMH6(YEX9&&:[)dAU<f=;_G+f
F9UR,b9_EX,H:FJ21/_PCKMFGeM6E^G)<O+DS96/4H1gVJIJ,IYcV_+M.fdXbPST
X&;B;aK(=M[b+ARcI(bB(<94@0M^9^I<KVT&?@W,bd8N5fag63&OK6Zfac9I#?_V
X<Mb+PH;52F?P-G7\>Y<XY0E)(#Sa7B,9Ad5N/=c;b+gD_;1_E6^fNHH\>FO_-\W
SGD87[W6HVHHY1P<0=VRFYUc6&K^970>d+d2P>c&g@O8>6+8-W[K@D=OS,)>UU._
^2-UTBeU5[#\6bgMI?OUW4)FcL_=[4e5eNdS8O)>4d<.HXHB.L[F;IQ>HL5\J8d8
8?)24=K3;=W4Cge>A8&Te?;/D\9-0PM<=5B8e0<bA\24,7Z:?R7a9Y19=OTd=J_@
^#M,TeaZ9K_,6.,2IY23>#E,15((K<SLFBb78JHH7F(9P7OZQ6>VG4G2;O.bV7b^
dRDCJg1c#.b5fOZ]&QeQe(?KEGF[c,EQQJF+OdQbF.4WB1/V&7(FOP,Qg+=J@=JB
X\#I,LPS@S]Cce>3M4>&g)YPd7O_RX[#Z7b\=LN6)<92PJC89QCP\F?;VFI:DG/7
bagc/(.e_GLR4CRQ^+OUDD9fJ][IULF?,c4752)Wf)V]a.4YbYLKM:gV_L+LP>]U
:]^J:b>K],J,QeG1JIL4^TAg3JfG)0>CIXa))S8B.^^Q4:2GN_&(]NGP2//C&FO^
VPS]:F>#8TB+:3DQ\eF(+#O]9PH:7<@c3)I=#-=Bf/BAgeS?[0=(]X0:?Y@V,I)L
YX=MP3=+R<Tf^@+(.DbTH3#cYF1f1a?8;+I\]UP.\T5QQ1-@O:7\,f&b6ZG,)-10
TLC<cN,@9]D58@W-J-T+AUQMdV4^SQ0d;]+PDS-;^dWQ>HBOT8:S^JS_6T7?1[RO
AIEbP/>A877/W>ab2(TNTe\Fb.#=Y-KTVPgXS7,6TNY+2G@dYH2;P_0YAYF0,\)>
SdWd>I::8T6B573aB&Mba<-f.^[9?MG]=_(70f+TA1\Z6aOc:<9M]APP(7.T98?R
CIa1IX1G\KgVO8ZV^07+W3/N1Bc)0R4#]Q(/#]6YW=92cggG(Ee,X\dg8WA-V_^,
BMf:f]Q/eD<bDS&H/#0<S=T_Xb8g<[bRL2V\57TSA&TE^3F#-gG1A_g&V@WHLeH6
,/_I,dHEQXd7YQNb]Y5\CT];bUcHZ9;WBQSNRg/\M4bZ9CQaR,C@^6X?,>,c-.T+
Ce/(XMF^GAYX@,bLEYUY;FfFg\V(,[R7eef>A^.T^NGA4CWU70G>[AW<.,53]_,e
]&_f0De1;BR_R7NQQ>gAbDR/e@B4FPf:/Y+F/>IG]\5L9TELRg?U+3d:;<eYc\5+
RAHDG#\?-O<7?4@@K2E/Sc^T[DS3Y]5]/MRB6b;(V#RdI9AO]FU6#c1D(H]LERd?
3[WJB8:Z;>4=/OT</J2;DgO<aaXR,fQ[G7#L_T3M+4:V.G4b):L&V/W\),XRF/>T
W9]OfK=,eS]@9a?^V#Q,fAL6&33dS1NJ(7,=O@OHIYH(N<,9]I7BGbBW?P(U\_J0
eAbc4&Y+;bb3N[<\.-#B.\O>YGIf3e0@Y&?NP/QWKRb&#_]g=+6R;fe7>LScOS@c
UbN+RLaP;a)4)S8)gB2fZ:)7,Hdfd-7_V<,._9d@3AW:P/;ITM9@d58;IB(O.O44
^(+]8g#.TOVLM7I[&J]S;&&+@)3[;7&ba8&6ET^B^Tb?BJELXD2,9KD/bT^,MWQA
^5,2LdZ7f(G.[[GA#T=[^8:GF[Lc56#DWAOeB/@2HKC1(EL&0c;^DFIgP3JVSK^@
N,.g&7\2W3671ddOO-JCZH7,PXKg.&XLQdcgM@J)9+S5R7\;_dY3/8?aLLNDF)OD
7:F]aJ7Of>@Z(:aH8^d:C]IY#YX-T[1RE.33B]W+8dcQY]OME=S1H_&d7F11b<;]
3Ic4TB(_BU(YSOAd2-7+d-0F82.K461=2ZAVQAfQW;EO7+3Z6K@K_3<A.)X1Z1R=
KFK4f02R\O0c/]DH(.,U#DN:;G5A)C-5S>c6<6GM:g6&=/H.7[W8/@L7cK:9\G[[
.LG7J7DZ1cT/Ab4VX/,g+53bIPg5OR36KN<UH)+,J9Id0[#dUJ:7.R7<RYG+ZQU-
O/Q6J<3f3.>bL[M=^e5NPKDaeH1a#VUN]78T(>?Y9a6#<cR+BRGagOf;[4.=<aSN
4ZQ@F8W?\CcI^e&3ORZ0.EM&WCS3/:AJRXaNT9I^:ZAD^XS:O/fG>e8/X:agL&DW
WF=;RRe2S\b\SL&L7D]IJ)^(>9\<B4XAYB0>MV+E^9DS4cNC#B;TECe1=eV7Re&6
Y:.,:UL82<9VPHWC&9Bb[e_?We5dL9?&F^Lfdf1L2addHUMfT\O[,UHcL7)(0HK_
SV945.G5c1g?QS?fYgOa]QR6d3C9bOM/KUFf-3Fd-8UE\0HJAfJ5f2Q0bF[?KeDc
3TZBABT+A^G]P9CJUY>=^<bR+N&LG4-;dRW11.<<?IN63Ic=,R9?F6De,,FPEKVH
YL2[LY7\[>ZWOE)<,(2^&PSNXNe^E;78YSQE^,Z[FHM5?N?K<4Z?&bE76<]66/7&
#fF?X=7,:d@0ZD2VG-dLc3[M&SFYJ-Z+=]3B.7fM0PM;902PYR74Fa/.5f]ecAQ5
[UX+5SfG_edGHA23O2\IO[J5VNO77T0bbbge#U63M9?PP7&A=#&\J;#e:D[QCUWQ
dcdbWR,V7&9/(;-S)gI[DHITd7<E)2_JW8?.e#\>[)SMX@:#K.RcCFJ1#6;2Wb7d
U0FD7,OaK)D]>2L5JDM2=b2_\:<cfQd-AgJML8=#FV)96_HcWM.(UF(&(RDWaC1e
T3GDQ\/S9F6G>c-0O-\@YYO3@bN1I54^^5ZgC+)R,>&E]8YM8\ZM,Le6N:fUcV&_
Tc^:80c;B.&bTP2HF#0f<@\WN[&YTE^2Tb]9a6&B@X.[3#O?HVS1@;F@b9<?4?,Y
G.=#&3>:YGL,?(AT0.f-AS-9^8[fUTBIFTf:0-V_>T)Yb3O9GT@6>F,A.(+/<JXc
I_-3BBgG]H-DUCZ#.X6[5E.]Y=/OM/F)gZ5N[LebaeYX_Z9=b5:\H&[a]CSfJg-A
[-YYK_b/]=[W1GPBRWb[?JP2;?3CO<0T:D2(CG3D5aID#8&=]?MK3ZN.)2OdKfO\
=/>DHb7H;#;VE]<LPP)BXY[CKCM4O9fcWBK\]CLf-V(c1YS]\G/PKQEYGB3aIK<B
Y&gLbQD6a/NE]K@PB^:(1C:^H?Q_=VE3361S(V^J#>TIB]@+K^)0Z?Z]4>3=bTK]
O0H,P6^V?L,c4#@ZE39OLaF5GUP64@>Pc6=b.?:R?4A^^YM5GE5=9dX3;N7PSH\D
4bCB^^?K8c:]f^F<+J;I]Xa&6H2]R_gg:b)D=WXV#=(6-f2>,,E?)Y@fEY-PUT0B
dG:&,_JJ_g-),Pe1E6[>&@_#,6UX,b)Oc5J@A5./Vd/b8d@<VZ:E7G<f0\BJW:#c
AeL8/gVXRN^9D.N;^f]-Z+1dJCdP:09ebg0>>PW.TSM6;M1RCH6-&QK7W:PO2Z9>
^V@,(=ZCI.P2A[8U;)_KSQNOQGEO[M?T4_fGS]GT,[W8P;Tf./V7,gM?69)?U?VQ
@=(2Sc[<A-/6d6KIcK<]KFX,(E@ETfGd<2-Ogb5N:.W3E4JE7F6.ff[2RS8+G2Ba
EIe7A(1R@?6:-J8PMc2]R(K6V<(OAbTOZ0/=NFSg8_A2LMaARAF^Q:GN?W6H0<1#
8&f;-1/_JA[AY=]9UeW.H\PYA/@^>Yc=Y#F)dV]Sg/b8_ADYd/PJ80=E_/PNQ90<
DCa+RN9IbC9OeC>-V:H/\a6aYa]d-.37?BDT.-/Y##@2d(ec/6&g=0.<V,cGD35d
3LC_F?]Q>NG<+;Z]Z.F->U@H,@DUaWJKZ[IcbA.7EN;D4]^L07Y/UQZ)&+aH4\Ue
CX7[?-A<UEFUO4cd4>+Tf0AD659&2fXSIbAg4)18g-[//:XB4<BF^eLA=9(.I/J)
R[f-=I:L]#IYF]P09aLdJ6>^F&[/HG@PK^\NG\(fK>:_BV-bb17cSQ-Y&d,f.g.U
VWM-f&-B[I]L35->5L-8+D(^IbW9L7^#GKHYFaOOJHU/5;S=.IRcMfC.E7I\3W,&
;baY1</7V[d@?K>0/9cYH+L8P]Fe_&(X.6AF6V2Y0N(VC6E4R,fE,J,8d,bb_V#A
;/bc+?-W7)<X1^C)&FUR0ILPL,4^]]KUH0/O3d>]=5#>#/4LR7^;XY430c]1)9b?
g4b0cZ&EO:=+,)c77?d+HODWXa;?1BUFVF)/ddCa-eIKOPA=0X#,4.@eYGNIFL,c
AbM?/[HGS<]IK+JKEC:A(-6-A6efd^RP\d75,031<eU@XCX#M6<\KM(KC-4G:S/A
+AeQ50D1g_VI0Mb).Ec3<K0B(V=&3;Y.]9/[K0e?P&,.XKJ5)-g&6];/VH\S:2.B
a<^#OKeV3C3TeBLO0K7JGM4>3UM\B6F</K5Tac./O_<L6VQcZ@2?CE;FK2A?Q(d-
bYTGOD):(J;6[U4=d43>JN:4O>aGBXfA+XDB02KLF(UH&/&KaQOaSS/4Z#V6VEHK
994_B5EZXJ\[BSGe0TDY@,<H0DOJMX-[UH:Wg6f;P0B@bM8EFQ33CDR&4F40[WO1
&BZ^>-):dD0?)J:)=XZ]-WU^\_.CAUZ]62bY)TN8V\PYGUE>W>/(3R#/7SgFeR+]
<-&dMQ;GS)Q:fa2EbWb<O<JK=H\:P5Q:V5>d<OAK+)dOaaO1YK>_1K#G>R@G;bC+
;?]C_II9,B44B986U)JRfcLfAIB=VPfAM]f^I9H\YQcG8?A8UcESU<Ce@YD(A^/;
_P@K&2HO6@/TXD:J31@2MaJ(2c>_Xa)8D[bfAf>aH+DM=_8,f[R0C?DB]XBHJGY-
.^.]dPU<#e<f=2I3V^?-g4)]4LaTBU3;CeMJB8[Y2[FBegZa=0c[59E0,NMHS)=Y
U<7b7X\I+DCH<H3H&@2CJPJNFMB9W/G#8^CYPO39W]K^6;Y3U.-T#?eBLUF,OM35
9VJ]ZD6)A=J[Y=Q2g5,aZd>?4-HU[MA.dZR>CRg<LOE4U,[Q@HP=.@bU&O2[1]#2
fDV?S]\\Y)WS,=J?Rf+KXX+d^UBEO58Ed5g4#WR<g3;WOfKSLP?CEfd.J>@F1LXO
(STaS5H+STO\(DZQf(/WX[IcFYA6.4eM(-2a5LdaVBRa>W#OcZ4>F^NO]9BdE(,-
-AeQ?YOddd?K=Kg8AKE&L;ZWa.3c?IUe6]JcXbRL^._3c=RN[TQeFg:eS6Uc&dHE
@DRgHd@DQ(;4SeK\+]PUP830I4Z)bFZW3^2(\?>JGd8PSYN71^#95Y[T8H]7VKXP
,?+FLJWJ.f4\579bCa^12_S^;HFOB?675T)YK@KH4/8R8WY.NUYNO/KD/IgTHB-)
Q9ggO4QUga,fbe>K+891Y6#f[cOGUGRJJE+52&1b78E7O\N;U9TdI39-e>H.VD_H
QL:UD1+e97[?->F.L86=gE^0\U@8_>f;e;5OO8?g-,28K-O\,Xbc1B8YeJ&\;RLU
<(7S.N89RPc/e]V0aB^92RR4EEH_KA,N3FL.G#G4V8C\NX0U+b/4L288WdX@DZSG
#R_5DRG-A].,^EQ;AbaVZ16RPcF,?GO@Nb#^./S]SLU3C#:fF;=Y/ZXSX.2D1WfU
@#Kg_1]&Pc:g\IAD;V/#8cYSZ((057=WKgMET9eFZGT7c(G\Z1WXLa>RHVVaVbR2
ag^E]^#^3J;B)2+);JZ^3JMT?WcJaR(bRfEP&B:IOKHT:\_WXA(\98Q+RVO?1_8]
&^D1C8f2U;44B?ITSS]N-WR_0aWU[@(O/Z2@-^[?(&NX<g/)6P<0SgQK543@ND5X
39?O&@LHQ?#7.H-HP@)R?Q]])&3QU)U&7e#W)]4M/5:),gEL/A#R=P#8X=d42_#Y
,F8V]TZTQVMF/C(@M9S(]IdN#.TRXJfTe3)EI:4&EePUM0JORFU,4+.7CCZ#eMQ^
\V?/4BcWG2M6de72,(dQQ(\G(g,/K.Z^8?a0)6Z?_W_,6LM7ZQDT@ZeS4DLSG\&/
FW4@M9:=^S.eAb+,UO95P#3=Y#UNeP^>)=552G72cG[?+a9g[dE7UTR-^,/]=#bS
dXd@aASMBfK>GT7c?GcN@@1#]8]TFDL<Sdg^R7X7X4.55O>fDP,6+d3J6_>1U3F3
fS18Fd58<6dN4P0D8cf)F\+K;_5:+F,(aPA<S9GTA<#H(b8bR\b^e;M)44NY.ZaP
-\:_LK1H0EgRLHM>UAc0cE>Xb2AgBUTX/?Z9/\00g>3f#E@5+OJAbg0WbQ;/^3,;
c:?7^-K;1\GQbJD8(0X:Pb^e>TV?)/L]>_L<8^+<)J>W<18A(W:ZI6d;a8.;69+e
O>,XbVM#?O^814/F&35O;@)M.:JD/8X_^4=<f>B-T949+9b6RX9SL==/G.>Vd3S@
;>KeLIJ28eM^BdJW_]R\Ug#4Qdb5]>3G=_K4J6FE^K;E^A<]F<3DNb_B#-ND#\+8
bYI2GY@(OJe\&OIIGc^:W9f,]c[;Ze<S)[#5^X=O^MO#<._AJ[M;>E/N8L-d?A0M
ecN:UO#b?&[6]_,e17fE;E@8L^R&J)JRNR@L(D;P>@GL.DCD;bY.(-:UF>Y0CPF8
;3>F9DYf8_X+VK,-cRZA+debO.WgWC+JG(ebBQ/cG\b_SNB0VWBN6VEDAH38?M@/
U2)X33;1E9e(FL/ZMAQeI+ZA9G)=\I&U>F/\5AA>+V_J.9#.?JWS^10P(=<60UEH
E\:LG\[2DO5V=-QCY5KVRUB_3</1U(6TOd9_,J9Ug[_40US?4f-aG-YM)8)ID4N;
1RZ1O=g6,:K#S=WegO;\]B4cQC^0(WHVPTgZGbFYY4K;Y2S[6&V3I4F#,HUg,-?\
OS?:E:0[7G>:aHJU\5Xg,X5e@H=JdA^d-_NSTcAe:DPR&\&;0/P5.#aB7+&5(=/;
(2TNH^Z;NT095GFg@dKTL99d_OA5?FRWaUNFX@0BK:bT9&OEfR/cBC@H)_X2Z=KT
6VZT]I:]=MM->6>><8W5KBV,,1PZ\S3E.\>.)]L9_?>(ZQFMCELX/cY74=.4]1QC
e[dYeb9MN._D>_IfQJB)@W-_K?TPQ)F9;MA(ZYCd2Q\[R;?\GJZ7?[d.-5HCKeW,
e?:_D71#ZTBMgXV=SGJXcgc0a@84Q+R<0@SYL7)1KZ_:7TJ:20a>E7RUYg5(MNME
da@>8gT]+^7e5APK0PT3@SMS:O0O:JIdK>IROKIM)=Rd)(3>3(_M36g@L2<EXT[G
2_Vf/4R^31U@MK6XBQA&[S@=)=18FWgB:51IY(GefgeA5c>OQ13+A5;MBT2X4eDN
2ZASLB,,)&?99705]XB]J9>LQ6Y&Z<V<U77eJ3;>eH@aC<Y6HUM(VVN4PXXPJYO7
gJ)g<CdG8a26CW@?Q._geg\73#(c#SJA5Bf;1[W,_H(U8_1+;0QF6d=FWNd1.O<1
8MLc2WGfWbfF,]XK_SK6[\V6WBO1@>29\>95f@4=CT@Zc-.cY<AKGf^,-SLD^ZX\
;gSdYBKKTN]e35_a04TRX;>CgTP(ac6#123S6.+>3B0<1E68g3HC4(=.I(D,364D
H\<)ZAd\M=V0^09/ST];Pge9CZTU1X.^64:&eOFK[CJ2=?6(P?VgBIR]D(T>[A41
#S^6DH64d6H;GM/(X.\7-3T+<5K06Cf6HL_6cb5.Le#)5HaI+Ub:JB#U>AE(:F\B
1be^RF,3Y0Tg-;HMc>4I:]7,YaM&/V(+U&ggN8#UKC.Ye>28E1IR;299<>EMSB_+
MT<eH+&I:E1=OB6gc;)X4^Y\JVIgSJ5gNQ><SO#I_)\gI&Ib9W)_=(ESd(3(_0Eg
([VD#2cfgJ/5EEf(\BEDO<bKR9K)S#NNe@E=,_JK[>/A4-e-<>Lb8[O.@:AaW834
>:_/fJ/IG&B+/a43WQZX-4VfPEL@&@QX8+N)N9]QP?FWd(g]R[O:AO25G?/?M=@b
3e;@+Za6RB6<aG^0aRNBObL&LR6&5HT==e>_gPd?R<(^3+##E.#G6Rc2-4.G/H-<
Qe]9L7C;)L19e@SO]:CfGAR,NN:^a()^QUL/#e>:ZS/5./Q0<;(OOF8C(OCSK.gA
bG8/23HK<5a=[AMQJZNFI/+]dbHOG(P@W_B-M5DWCe=XSDZLKe#?3S3g-Sd1U<,E
4BJXSGfO#1eU[)VD2:^,Lc.fBd2<^FO)2(3C6WOR#,6IFPf\1U?0DJ^#?f,fbZ7;
c,Xg=BG)e3BO7YA:eB,WHL9a&d1A)E]/R4NQXebNNCYD7S_H,=^7OE1A7BOU)B>A
3>54JEU+_;-1a@,P;.@/WW&Ra933S>>-(Rd<AYTH4aI&NZ:3#eMB52O#aT)8(5/C
D?K[_NN+d=^IbL?#<9[CS.=8@1?/DAIGP3e]PfV+;4E+7M@.K]/FP/E8YXE:O#SV
EVZJAWID>:UP>0CfML&H0/AOLF-#-.D777V4DMOLTMW+2HWI:&5>2A)^DB5SH:KA
(1b?S;C0U>X65L4Z/Z&aQ@^5]<L<1G#....2?)7Zc2da4S@b205IXggP3O,[)I=3
d4.QaJ:#57C8?/JXZ:-.K3afcZK08GG^-CB-VLNLLV>,A9c\d,,A3UJ2XBg;=XJ+
#<Z&/_7J7FG][]45I+\3_=@^ZE_.aC][PCV4)^A[,]4(N\CK>14&gdLZR.0+@X;S
/&0,#d3:)I_9UgS(NU-4/K]1VPacBYgDS1;]W.f&a0WfC?1G/VE@_/7BdAd#=M,0
?)^.B?<<>dZ;WROOe<-aJ5UJ\L5U^5WB#+-UPJ_A)eJJCR2/dO_(a7DQ^Z516FM<
,\2)C1gVC0QbT#/BS2KV_L(1V1HRE9-J:UE_G0ZgUI4([7IS,9/g1gO<96D5<b/L
16gH@LR@(<<<Za,?/c\R;35>&PDWG\J)R40e/77N[=^D?V@G,TN?/QCMO;Va=/.L
^fL=84Rb0WT1<TR<fe779TYO>T,=U?d^eb#-ZA?c?AS<LKgPAN?TQC3Q)d/9cGEU
LE6/O8L3E_&(TUEaN_7gM)Fc]&&BL?+A#M^T.D0OZ4_bQN)+Z(CJb?dMA=O^U@ZF
ISYE(Xb/I3#I[127a1;A9GDb[KFL77Q7+b2,P3U6.JfJZ(_(bMQB:bU<Q2bGC7/0
EM,7^Y:_7T\U&R(f3X&[d(_eA5B.F]f&WT2KH]FM6__H2,N7M^0E36-A[9&^Ve\(
3Lg;6bF4?=HE2d\@5WS_dF1cDYdeE?.@TX&^/RSLG9+/4dOR@G\_6QRH,KDE96I#
+01L9[1d3ZBW:S-,bDU24K&&[D)g[;4/aYXBK80AFDT:R2I5TN[CLd>Mf(BeZfQ>
fc;.AOG5GFXgc<dfI-_[2>ZDQURa7\B.,+HWCSN4a-B0^]T]f<(4/<6)aN/;7g2[
JM3)c<#Nd+&47L]+D)BFF?)XQ/J7#O4B+Y)Z1HPEdT)?N6X3g)4H4\?DV-Og/:G,
aD<<\X]ML,;A]PM7DWX?[86^V@VONXKJ[TXNKcZ[H_9ff_RRJTS@9FN.C60-QfV^
fMX>;E9A/aX)gg:BY4f5DW9U=#_Oc:J][[W5=BYIM#(T8\KB^5457f-G<W0FJa3N
b?A#D?-c.7LGKcPS.NZT2TF,@>KUJNSXX#^c<ZPC(WFB&]8g.3D73=4dgO5a/E<H
D;>CPfd]&a63XF\(2]9V[Y)(dD/NK7Y.>W<LPIZ3#TVcT1SF8U&(=J<-1-E<ZP.W
P<]2^2JRJa06<9Gf.>a&40bW926?@V#PgE#/AaU-g-0-.Xe@@0?MM/31O3f5F2fH
QVW2Y@J0OceHO6GJN#b9]:S8RL2;QFX0LQ(\\I(M^W:)gD\\;f,=)VTRS\ae0<Y?
3bH1Fd/fPKSV#/<G-QU[ZPbHNB4DM4ga@7S@69f5Fe_&NVCa=/35CFM_?/.>X1a4
U4;SY&#aLY]_b&.@WHA[78K.;=R\af]f3GU[YGf0eYG&dWZPeJ?d-KZE3DLU7Z.I
(6_4\Dg096#URMZ<]?VG=H3_,LBV.g(DB@F.RAe@b9@G@+8aVcOS7[QI.:;(TAg8
AF_OS0J9#A7Y;Qa&5bg)IGbdS7fXUWZNB.3>BSI_5M#E?U]8]JfM-</IN\ce[bAT
&SF[_JAM/3I4XB5fab^L^Wb89M5dBCK91PIC-E+GX5->JJFZ._\H=4H[;5IT5IBW
4TE?+K0If^2SRH1(_9@g2T8&ceW1G-KaDI,g[OWgLAa@IBH/MC9YSAT^@.D3#UBC
1^/YHM;]^D)&PMU]EJ#_W-4?K<2Ud?&N]UWR8:gA;6Q9VFC7RfeeE,7Y[cg:WIAA
HO::3H](6,a1fY@-1#5CD(BIO3-Q,A)^Ce)S3=_9eV=/e<AITDS][c=OQ]]B6O0e
;faYBf+I9&M::]GXDA\CDYF6:U8YHOK=[/3VD7YE8V)SSX;<WB:A_\Z#V4Ad-1)+
:RCeT4-f.F6\D[/1.3EZdR/,X/aKS)W(0P=CXec1bYTO^dae@U2&>[)N(I4bTb#\
;A2J-<JK]CN6,QUD?I@8AY8QbYH)6bMaJ=JVSQ82QC/J?7_ZI?Ea>Cc52E9f\2<;
_XL7N>;Nf>cOK(e08D15/9Td[<&7_B[B(<)d2a_BM,[,Q1dH_C(\D3#(R[GgOf7e
&;f#;9ba-\\2S4DKSd5R:d&7Z(#[<)X\JMMUQ:3BVgR->UaB52GfUOSE7?467J+f
I=(<Z3G36]T2e29fO\Z3\0&3,,YH(WKYG:D]3V/I\3WLTBb,FR#[UYX]IJ405?-X
1eOb(_e&?<SU0:9:+P\?2CF@D+X_G6./fP>JEA4EAOe5.5_2],EA+2@I+e:?ADB:
R&OHC,0+WNK<dSXQ-Z5)4J=Ia)d3F:cR[Gd8\be]6fg4ZaN;Y9SYR.gQ3M(X(Vc5
MJ[=\M(/I8deU#BcV&S1M9/V:fN7F[8S=K1Y_bA>gJ9Ibaa24,5&/ZJ_B.UZ#d5T
Y2FS-.])fK41/R]Qaf;Z#\\6e,#PXM^S)=)(^23G66dd\J3/Ze?-:;DaLR<>0:[.
_TKLW8Ec8A@FU;Aba7:Jd56EQRK9b3Y1^)_85.Y?CeCH+;9&+S_#?)C:,5;8N6:1
dC6Q9]6_.I8\PMD2[Pd:JF9E_WL]R9BWA91PVRDD==6e<Q[>FH60Cd^e;?C5b_EC
A8I3EAIeDR^IQ)81dJ,@>]OL/85C;E2bcIGW4abV_M14_L,HO5@8HBF+I@&cT=Df
OCNCP2:U;AD0+TaLGaV1T>JW>e8b^D9,9eNPa5H,&f/3>6@#Y=.?Z1RN&Ad/\8=,
QEbU:DS:U)OC0[K]#_(B>CMI)/2&7]VIUJ]M-5AJ&FZK-6M-?@,Q+Y_5a&6LT]+\
RKIGB==EZ#8QdEg]8YS5806C[X:1Y_Wbc.]/U?DPLX\7[U&.(Y;NHE/>,bC-M];c
]b_bM@6PE9U:>(->JJQ.ZX2GU&/QQ.fO0#WJN:?&NK>P@W48:JZ7.8L?9ea(YUSD
dNQ>\Q?7]Z+3c<AJ2]75ZSXgAeD+#8TZQXB4g7:<K=cf(#7_2,2<[WSVQ&.P2=,A
VD&R29^D(0I9/QcD2g<AgCEAOgWAb^I562,0LG&]Y(8g;X=c0/(ZOd@2.^QLVUOe
R:G:KNK=X4\>KEF:c1R(ObD<3F&#BLI4IcaW1SJP:7Q1DGI&8Lf^IZB\g5@2HV4P
K<;_N<dV1O#)13U2?Xb&/=Z57LRG3>K?#R:?8M#;.8>bWJ4N&>04QWH2^\MQ+/Nb
DfP\_T3\?X#PAJd>RY,0.gb\W\_,X-a?H5U>&5+a:GEM(9I4^5EMTIH\P0H]ZJOI
;Y7IST?LJQ-C2R8aJd5;WB,e)^R@A9>RE=,,K\OaK)WIT7>Mb^NAG9N687cFS2T3
g5Q]\f4U+UO8E>:M#[7=6)(.IeF8:.aT(.K2ZE+E/+K:Q3g<eLL0DI\;Y_CbUK6L
K?PX?F[\\FYC378Y,;]QMgI=3b0HY>RHN)SAAZdd;;<e-F/QfMBHDUQae(#V2C&^
1?[7B;GQ5Z;bGX9e2;UBWZ4.JPPN9=BHS>MX](;8g^H5/A:1O8]>&4g[H:AQ/2?/
/7I7BS/_-TEEb3]dD+F6;1D2[0^X@:2Le2.HGS=a,H36Y7cgA)ND#)>bK5;]E[0R
RT[bG4DL?&@H>g_B63A/a/S8ccA=7W>?Re1:b5HT#UcRRg>bC[X]RY[?Od]4^6D/
3[1J3\,0)-Mb=]AbK_TU3fJ)-8M1GL0M=RWN]E;/fc(6CaVddA9\\Mb:Yd=TR:06
f^5.1J,,>5^09J._V7_^ac2Y1=RN,ZDO/&=_BK^dEDSYDI-\U_?DK)-H]de+c#;e
MF0@EB+;T2aVd,^078&RaR@)SH<P0eT=L^RN6<>WNC5R,>bWX+<50V/V1&[1&,,J
FaG025X;^#.;<J@<RMNPJLO,2^,)f&RJ+&413-LD&N\aY_4VEdL.Ngcf9,Q?J9?c
89>]gC+T;][GSPTI9,KYc:S48<OHX@@.^FPR6X2_21-Q3d9TdcHf7M\Ve_Lf(dXB
3ZD4JSaIWZfX.K;N,?[)\GGSV4EBKOc0]?/@+F?b7CMb)N+0L]BIFObHNbd]+L9>
Ld-6&Y\<DP+&6a<C2,MF<ZFgd?6(K#C)6LRJ4+bM<aDA#GN\b.AaQdC7e9OQLcNB
ODT0RIdSJVK9PGXfNABD3\>dN>==YZL?)J;R\a0IML@gL=_.:@@CD:aXdQ]PVUeH
Z\Nc_QF#f;(5DS_;\^b&A4cREYM#5VAA[YFPF:PP;C[,E\@fW0:KE86,Y83.&M\=
=H@-YN;fe^K_=B[HS/dZ2dAANEfM=#?S-J1,L(f+O;S#3-:O6OH5a((3&?G4MEX8
&/N?FENO8ZT\FW2S?)K80R?:#HE-f3c7Z.40,LRC(:3&_f)+fY2NV-::V1OgE-3a
2A(Yb8>[TRW9A4dFU08gegGYcWE.6GO+9_G#20A\Nb(cH@ODZ^UU3:gRVA=@55PB
&:^>bU]Z5Xa695f^-Z<U[O/4N[F_?bS3)[Q?[g_5)_[[U2aUQN>3aU9@dZ-#K\\\
AMAPUb9IM2[eeH/bM4B,GB2493B>5a_A/G\9G6J)LLX-fCH:5=1cF,1B#3]<<44X
g=[D#bYF,c_Ng=K=6N/P^,0^#^5-DOSN9[LMa;/]W]S^+FTWG_N4O;68YK3FH3&Q
=Af-c+MdVG[d.A/(D=<,(aZ,d)3@QF9,X-<GY[TCTW/MC#>][dNNZUB<TI/U(_XQ
M?TM=BXLN6G9T:5^&>U4X]aI^7W#KR)]:YU?adC>FK4LTAXPJFbMb]+@MF==THMZ
-aMfJHe]dX:ZSED(#FU09d3CK)fAg3H4]R2>?Cc/E34QBRRFPCGYCRdS;O5TCQ.?
3XNT)1BbL5;4O<^6D.FQH-b.&471EEX1U1Q@Q).P)]GHE4C=f23acM:N@R<8FX2g
WXGP,YT)VV8(9ID/YK7ZTBT#e>\fKNBU<NB[(G\JW4F#3ZNV60?._8d+9RA9c0;Z
:Se)MG,VZDD_)?2IGc.JYJ\A8@gN]]#aBD96<QdFS>f7,=#,ga@E/[9gACM1H&L-
6Y#>3C;JTAY5^E\K:,[;BObaZ&H<Yb.#Aaf:Z28)&g8/800OJfYO(<#ROOY>NCV[
+7UGg@;_W&-SWBa(0FOV69ILRd5;;Y4&E+HPcE60Mg^gE(^DBg2B+E)gI=XNS1BG
fJ9(N)[g(K;GW+WBDGdEO=X4_f[F3.OAMJW3PH,7+NT3>(BRdO\>CbO2PgL4VT,d
E(JJYe\?g5AZP+)J^,?BF>KV?9T:AP>292D:AdH23/E=<:,N#@TfF;]=eDeFGCD.
<7C]/S,IRWD7K>AR:P#C,G=g+D6Q70A-I_GG<dJ#2)/fbP8QB-\B:JSH?(;G?dUU
?)H^W,GO>J^E[E3FDW-7.fDP4^39S=<IYB2W<N.^,Y,=EMKdNVQMSXgJbHOEJ3eF
;2UP(48LV-K9C-Y2EMDTZ4]TaaWd,#&5L0a0ULU)X6Ib#cYK5ER;.>0)/fW:cI+B
7N[+LaETA]4(TWJ?Hcc[EIOGQ(AJ@fX6cB/,N.1dP>9U&:GF?M.46]]H@eWa(;I,
/fXK_UTR^VB_&)FF\a&(#CBG8M4F>&6(_]BH.54g<K\8X)E0da.W(&AZNcWXPE])
F9[)3U.K=7>:-X/WR0Rc#-84QTKF>SSE@fdL0d^MU2d6W)4E1::-21HM.1:/;G&U
/9GA\5I-OeCB+[0c1X239WI6;I_D55F0R@9D1UGN#a5,(?RL3Y+gAJ8S2&CJ/Y3[
WCZC7_gcM4T(D=5<GLg)+[aM\F;M51J>bb^3C:>20/8Gg6;;#E)7#>JS,0IB5(9#
2E09cN#f@9JBB&<&S(NcOKcZM:&_84V4=aLJZZ1gR\86f]5-9)I-QaV^HY+3FF<(
_&K-/[]RVCZN29M1TBe+W-0:92-OaC41W[DV(OLW?_](5;79gNdY[@AJUd20]gN[
RG&?HXVRMEY:?[Dc@dN>L8@@)5/:<5_?22RH]VXCeeEdQ)O)K?V_2V7Q5W5La_]X
?Qc0J[)]R9&)dX]I8;fa,/GegM;/Ea,/SgS7>J.(P?_0=b+;2UEDO^-NEFQK5D0S
7U:@AU[^+A)Z?\8S:?3MZd84]Ae8<:W9b?Fb3Qb<32O4E]FYeK&e[8HWE8.598KL
EGXgL=I/Z+96b/c0L0+J]=^2QBa@F^UR:#;?41&beH4T7gBdV8V=VRP,13Q&B7;8
AGQ@V@E;35+O4>BW,43<a)TQP.(=W;N>N50&E\+?]<8cD6V^DAW/f@K;;^\)&Z[#
0H=fV.3g6;WL2-IdK3IAJGJ?K5dGZ#8P&ZG#B&-<-fc2_6TV:)1FXN1^FS?J33LD
7R2X+#Q>+A6FMbC-_Y41)dL-\HMeQ_VV:UO92_L1D,E9c5Dfa/B]5b(U(g)J6Z/.
/)[dNAF>Wd[=:G@ecG5F1ZdC369AAKVg#I\d-QLI)^1BP2bGYf7;W/;2<FEXCP0I
U(U=M.O+6PK(>)9E_7R2EMA(0P;,7_9H4^IK/bO&Q\aca\(7d.ddI6Bf_)GgVGc-
CbA2<+bZCcP^Oa:7</[JW?b8PCRREGG88OgXGGU8TA3)DER_M<7,a?,Y)f7V4O:_
W1MCTOf3^YZg5ASQ28QMY@TIH#HI7b0/78a/TT<0Taa)&N;.La=^QD)b_3@DR5)Y
?X6?+.J2OZE9)fLDeQV\Ug[AO>CQ\6W0&dO@fW=6(@9g[9;Wd(^(9Q_XHZ-E^7X0
EAM.GLKKK\68G+BWNR4c0+Xa5^+NIa5)Eb8=7=DZ=(.]ZA.L^SELCJS#eRPe:G.T
b.E58,QGP+0EUeF+V#>3N;08043BZ4P)#If<Y.NB.:Z:,5>S+8JfA[RZ?6\\Z,R\
7CQ?A&CV8fA,LH^#R.Y\^[CA4?E[(7AedI,S);@T^>5BdbWWY\4^,#?CS6F\,2Y-
BHY_6=c)Q4b)?Qd-Vf3<:D=U];(BC2ZC:G<[@+NCF6.G@3D_&-I_KdEWPWfYcIc6
+3VU+M@.D<Z+3//NX=,5cCgPPJH>5&F9OF/8]G#8&7(;;0OOMVf:SPgL:75Da5(=
e7MKaU(P2I7)/GTbF0IE/H/K,67EMe?7e,D@29D/IeE>,O5=a<TW@;OJJE8NJP7H
IeVGO1=[=S.R_L5g/L[3gf9Z-^T@]d=HN1M4PJ2673M:EJ,&Hb0G>,V-_OU13::B
B.G#GZGGg_^[)3CaJIC@KbBf0ZL;O#aVQaKCd)S8W#.Ed4,(f]:E=PIX2HY-+YaH
D4dGLXM6K@VAb]GDOB.\&U]1FSXFA+/Z)5),[XSX^HP95D4eAEVNS++9=d9Q?31F
8gcRL0bRQ68e3[K/Mc7d\2CU?[d>:#^T#)&P\[#Y<E;B)02>2O6>XN;[7W\C4Zc5
[W\Ze(F^M@_S]M[Y+0cC\g^:MW#X(a7]gJWM8C?BZF;ARdU(PX9gQe=,_26XZ-]I
(6AN,SI9a8#?af3E.Q5?MB<3)+86^cR]J[Ye7:/UX8^SP]aLT792<g.C?_R8)P\R
g.OB#@g9;N&NE26HaK^AbJVBf-FSOAB_HS<4-dWMG963>M,HFG_]3-]M6Y;=V3#W
a6P4+E#J<GDbb)CD7=,82H-D^>;Q^(VN3UMK9dQGbbM?XMVdX:Y(:#L=c0^S8FSd
G?2]2W1Q>;3Pbd&#D3:ZO)QWGV^]8f:E6a6]fY&7U#L_Jd7+VSf:^<dG5,WXHaM?
de5K14?^VcM+IM0URK]5TLc&4#_[b4QBeF0//L&=-f:9eJFX2D#BQ.N3H0X)^@T)
B](=<)c5AIT572=2^>:M[KN6a=:&^GU:DZ=M#W^CG+OC]>f/TB.Aa^IUaAO+aX-T
9EWQVZN)D,^Z0N_2EN^dK9g4PN4Z7>#>aQPZ]PUO5_.C;@W89+2GeP0E0>VP8LOW
:]Z:/Eg_f=0OGH77J[&dE5)XS;;^&f?03;,>4M#W)N+R<_F6UMLf[RcLXQ9C-;cO
T<cCFD-@a0\11/H-PdIWM08@Xfa<\_F/gRbBQROCP]6WA#6H^_D=\d.X^];^JZ+H
O<7Be;.O7a#0)RHM[Z+C5T))YdX[ZGHY@(<X>;26@@_[RYO>;CYBTWNAWV3DG>5B
eJ@&#5YETW]++#[3GJ#B,Q;FU6AWU^aOWC-IU]AaAW#)0_FB+W?#4Y=G6&R\O[Y+
\f?_P?;dI[b=DEeI:]?/)NEG:K//?QH632/0?0<G,d&eSDF]c,5FPKU\M>?79B-)
;S&XfCc\P4OJN&1Wbf9F4=9Gda2XN)eC2VH1S4<8?Pc[4&K(ZJZ1G?HVYQA#5]<<
C^)GggeB[a>cJL]baPLg65]<ZEIJ?/LGGARLeHd\ZAcMbNI&GA#CKLL4GI8&T,3V
K:OgUPOGGB^[]T]H=],NXR]T>?2SYVa0,U8J6>NW843_\]e@U5W7d;X9\IO-D;L^
>M-bN9VFKX_3W&G:LSIUWB-T6aFJC(2M^TMc)QJ6#JSM;,^NcGL(@6^&,E@,#7S-
8[Yb&=NMMKd@;+#5dZ/-2F0-,KJ+(VMJ)-.Z6;UFG1(/20IU58f?NW(K\H)V=>;Z
@#[3\#:QLD=3[DOc&(5(9:F]A5&)UEF>#0#Qe9VI-Tdb>SDg8>/-JDA>4UJ]-GD5
-.Aaf([SLKNT]:EB[&U/?aYWg?B.ZU@ee0ARA[L#Z&WFeP\f<2CBa65H=^OJ?W;O
M,b&Z(LNXH=Z5\aE,LO.2[O.97Jd@B2<M/)0gIIWEeERbY+C/J>gH&NL1\[Hb)]:
GH@F3^+RV@XCY+7KRTQPF2.eUM14S/P,SK/-7#.Z++/BE;8,d1?;34LL/,D^1;P\
J1fH1^;He1(;]D;M)NWDDb\DGG@Qcc1NE\(+0NVG_M\N+9:dH[1FQaN-\_Ie3@ZW
?5/7d>/3IDBP:MW\AgP)<M;8QTc9Hd@JY9O-]Z.2H>^>#eJ_EcJZ?6TIM[U,>(.R
8L]MEd^GR27fR&TK)\g2CY2A<;GCH=OW_bP^b.dGKD\e(ef8Y2Fbf3)8MAf_U9fJ
9@2]C(4L0UJ=-d-[7LKW+6^N#OTE<OFTS@(<H)8Z:)<_<R];3^QWEK.?LO_VDB27
X.Hf9:<;VeW[GI#4JE3fGP2Z?aW?MXgL1.QY;Za>GY?gPc7P^>G+UQ^0Q&.Xg<,)
JT:/)gWF:[[]QSBTRUeS/NR7bOZ0+1.^QH@[T?-a#X1&LGZ6<?09F\ZU&1K?U.Q8
\++E9LU3?,3b[:7W)K70a(.-(cRb+U\=8aEKI7deAO<0,:R6/+^TE<RB/8RW5P8A
eDXc3B,>L.O];S38e1E-[GM?I=U<Y,469+4G]_\-#N+2#]&cC=2KdeKDYB_6<F;>
852f2PC5G,N^fe-Jb,RIS0A/;D2FPbE0KL-X?,#EJdT;\?1/:)dgD.6K?+T<0Oa=
\[M6)?]QHC]\M5275/[aA,[-M+)V91\@NCLZd26a18+dH(eU)1T3L4J8R[fO65K(
fJFHAVM/[@IG[O2:YY#f^?Y)]SBU8>.#g39.Z7J2)YAdXMYMX2;33A+&0CSB_\R2
3Q7S#)M+f9;1R&a1FM5aEHIe9E;D2VQ/c@@_bX0R_cf,\UMf\X(S(6\Zd[73C;2;
?=IOgQdT[:Z7T5?0A_dBCgTe\^2V>&CP^eB#[PcY=b1Yg-5,YM7B2(9d,YFgMPG>
F+RT4d@L)g2SKW\WO7e)c^9AdZCR44Y&GQ0,c?>3E3FYWOUS[eT0f7ILF-_L5-Pf
CfaN9E1WM5(]aCcGfRaN]bN1&I[VB@>5<JIOX1XA4H/CVERDQ,;c0XA8\O+Z&D02
-DJ\]@AfY6#_@SSC:JN@.E>5H1.P<U8eWg2U><4(7P4]=.TCZ;]dc;[<<NTGCLK2
K#0c:T;)?Z#(5b#<WHER2aS25JeQ+cW><UXZ(0R_#[=UJc(5U3c0CLb_Kfc_7--&
fLF6b3?1fZ9WGK/]Xg.OO-)-3OR&W[b4RGR_:HVLV>IBP</J@Xe(eDC4;7\JT^&U
F3WM<e@b4(F8(JD\3UbRBT-c:07,#;VHdI\8:I)6^Qdb+DbMU#J@_RD2ab^_O7;Q
+M9CaY2L83c]_ULb:MF[VZ565,&#[\IcCM<(;MF81:;L0L@2f7).e4cC.W+MQ@OP
T:5N:eI9E0+-8JCL:)bfDQX@C5;#M#T]ULe]A,UVaYQL>dg2QZFK@Kf2a_&-+B]:
eH^6dR->]gE5F&V;_5K4CPXR;5Bc@b[FfOQ?FfX,WFb&O:J@NZ&P<D-W+L[W>/D0
R7aa2aL+<RR47V(57:aBIKY+#J=9B(-Y)R82FL&+,Ne/0291GfR)4(A@&+dWg_>F
N/4c@LBIQ>LS)&b)1X4-5M3O9_MX0.RC#UaRM1@4dVg]GH,NebI#5L2JOfO=._8>
bd=//B7(=X^K910Ad<4E_#I\,0[)8A[86/VK7^(<+e;f8Oaf\0.O.?A,X@FSYB2N
4F7FQ9TV8S>cF>5ZJR=?.ScE<\BPWQ7S@SB,]CC/Y_>QN;825C.C[J;F.E_IQ453
)ZP187OJQLYg8GO[a9)9bQ>>F.9_3^N[>69)^=6c]aM.21.4>F9C_C;M;\SeBQ#E
@W^XV#:4LP3B\7+N_5E5;B_QLHS3H(E??aY\g-\,NZfO/H0cY,gTb@f(+HI9>a<M
(OT6&>>2a)P@5:Z8;,\#1FX:a:&?^(K#\a#O=0UJE].+3g)/&T5<M&OfX9.d@=fa
f:7&^2JQ_K6ZR2?.Wd\;TNd&G);Q(EF(/>9(>Q(#g&<N>\<RR4W<3-(.@DNIZ5,[
gHdG;5DJR>O[U3]cS?F;<PZ22T2#\PUEEK^J@H-gW9A_M]9>ODEGa&b8?gaAaWRX
].K/]fCP>FBZ?473EG[?/WVI^4@K4O;2HMR0GY;]Y[C[N,^.D3_FDa:+3[04C5?F
3Z\?Z35?g4:Q5:cFg,P^7GJ((<Y[E)bARf26R+WM=1AJ,)I5K,GT[-I4\g2gMS^P
@8=_AB]:&3&G-Q6LUXIO8Y=9^^PEJK;&dY?:(NNP,5f\1N)RAg25.Sd9P96W[XNQ
&>J;F_g]&\J3d8QfT;]48&F]7^68NSS/QI]6aC:Ic57JT,f?FF(Mc82BE0BfbU;R
?A>KTH63CCfJM4gd?KW()S<VMWC_ZO9(Y?2[@fVS:JZd<X)DKf5VE+d_f8aBbKX:
2S,3S.48dSU4N_BcN;CW_+R,D@Z/=03.AN]19NEHGaNbg<5dJ/1.c8eQU<Y;A2ID
BN&#V#YZ[S1R+DLT.eF+g-OQ@69>57.-R3Qaa[1@7d9;f76_ZM;+gZd6<SU))=N-
ZgXO(gZdX2e>P@[gDdV8UQTcVY2O):DEO5^65@PA;>fXE7L^Xg=/,I@<1?/ERcML
OSP4_#2X2VONL,UdIL(0H6/79dcX#L[WR]AAbbI>DM<\T=BQ_<NMJD.QO)\2W1ED
g)HS++X/da@Q8RR?W\R04g==6_O]WG#QS\.N&Q24K2/RJeU,4e+CfU#g-H>?&X=5
L_J(2I-+]^NZYbS(L>SMPE;VEa_CY6BT^d:?+)I3BFbZbQ/V7\5B5;GX--H,gbG.
14Z)3Y.##7NL[E#BOPPfK/3/]5fXQNKccT)1S1SM]7I)4?)/T1]7X0:Z[&DNe4?Q
>70T-e_=/5/V?=TG>\]ZOOf7CA>64B^-5g^QcSf_SN79H(S;NHg5Ee???-4S6aEF
S)H)6AN1N-R+VVaa3J;C&-1_]/3cPgV&IA2Y=d&)[G0Bba#4<-9<S0D=SFTNY,Z_
=PU1EK:8:#FPW\.SQ/&4fK,>9NJ2N:Xa1KL8=J#Y=G<[QGGB:D:P6Q,R4?PT9F&G
72=c^8-._]+;g^c>R-Le,7EeUQ9YQ/GdaJ:L.->.LS;fcJA\;1C0bT=:I3b0]Yf6
<SVbb]dLMFRYN?gK<f73S8H#D#L2MeC^=(PT5SPfab];?^;DNC>5V(O8_W/gM95+
]XHc+K)LPV,OP6/dfE67TYZHB08Z,J[>OYV+E(#8OONS]4UP+&0S\6XX.Ge=411@
=PIHD^4,15XdN)bW:(8759/^<2SGAfJBf8M#GS=J^/+MNHRWb>](2(WU,CII/]aE
]_(?RNccV?_(BT^0dU,CBL:c,4,R1ReG880O>]-dP?O&A5MAAfZAcJX;&Q9eYc(#
PL(JdBT^PSN0IEN@2QF&B8c97N&-(\b.O>81527NV@4PJaZ86<;3\e5VG+S>fJ2L
F.FWV9[T]Q#CBKRGBT=4:Pe)DX_(O[G0^7Gf,]ZQL>cED;+J;aGG>B&QOYW+Yg50
FR#aYJT5BbNUf@/3f)/V93c,S/YNIcY_L190g,8@;dQFO96#Y#?;-Z7fMIJZ.6C)
:.5d4@+VEY/Ba^9@UeIU8Ha,[GJX&\fPVICX&YO>;UL[0#<NVC[@?5>U,4fE#P]7
+ba>Q-U,Sc#/G-M@/4&FSd#g=O06(SA576Y4)=T#U4<\?Fc@PA(R<0/<HRZGYL>]
Q[JdIS_V78Y_QQU-/CZ8e>;<X9eZUWC?XSKP3:[N7;(#VCZfY/QB<C=7HU4;#&@&
F@]MXX=;QO]BR]aKAAYD)8]-L&)5UV?TN</1)GI16NL_Y\:T&/]+IRY^8CS0d7+4
^?cLM^QC7GEa3LcF/OP(-BV;[f+?>7(9W5gCWaA[COaBN6>GX1Oc^&G[06^ET=9L
1#Z36a][LT(LPI^A_F[KH[Id.:-f2JAC]_4T<BU@,T#2+JK;G2M+D<9UKgTKgY_@
SWY(bSg7,6Y?MQENNcQRYEaAF=U<-;e\aFY01^bI?S8PP5M)Z\BKa[,HDUA)OCN5
Y-F\X]=_.DGTXdY([)HT6+6f]c7P-C)40G;D8)(Rd^MaNg+5(g#]TeV8b8;Y0Pa8
[O55#5eX:eDJ350N<>67,1#45TIe/S7OO33.738.Q6R=e84;L^ULZQUe;e18__90
HRF\e#?WW#>;>,LZ.8RYg/5>.;C.>B<G+7SI+@DQedTeU19:C_f0#^OA&GW[YbJS
J,&aLS14g:6gg]W-_HQ,g9KV_^Ef@N<EdM9\COP_G6eFC2:B#>0/^VOQKK9@[0DT
9dW#:c1g;ITW]gJKba9[[+7]?K^306e,f&O.d99\gU26D^P)HcVUN[5J?8ca5LJS
1K8dT[[3YF2JBYE=8d.g#OLe:;B0OgQV;+I7KWg)dM4)M-a@@9?WO42CGWCZ<@M?
XE2e7RK@/.1#Q0#HA-M3b:^.4g96>)0FXaB-7e-]099a_K30YFU>T+/e@AF(C<D2
f;PT-ZL=6HgMQ.;L@5@SabQ^TIK^-FCgJPY#P2D5,BH[+I)^L;,08L4f^#Y60X?7
_J_KH&>g&-Y__c](2>FVHF;S9I&0]OL2IT=ZW]XC/6(FIQW_++fLZ=\RX0,5:b>P
McUD7c;+,Ba4R8I<V]E\>5Rf^KO2;TY5&\Da=K&C/KYRCHUP#-X;0^U3.V\4ZK9c
O=5<WW7&@.5RJY_8U(#.@(<3:3T&[c1?^4]F;Id3:?HW@59.<BK[fQPGc4>@^#^7
@2YR9>3.R#?0;YG\94Z-b]+4.;6O9Y>0I.)(,PF/@@\[N#_>Z.I,4>=EV@d7^-L2
P^-6N3)194THH]>8LPLC#7P;=XG>c5I3@e]9>:I9Yd3E?8&DO&bWSSE[>XWIJ,8d
:-59\WZ@Y=O-9&d)IYHRMd3?I4S>Za/?<,;;K9V_+4#BM4=#+V9CVYK,@b>cDbE5
3Ve;/IC6G]T.46D=^1/b9?X^R-HWC8HS(e;A\U_O&\Kb9dHU<,,M<F&39==M>VJ>
@JdQdFH4W_0:J6@DU5?E).#&GB+A]AXW/c<e0A(4FN)]&/f^DDJ[77a=cIg]dF+9
I=;R(:bBL=:(T;BVOEc.R(]]U[KB]Y4d8J4ND+.3(FDWf1Lb]E,JJa6>F0-V3&7[
dH+d;b]0,=XPB4+KX]Z<B.0CQb<B)ZV+6<J-Y<?a][If\>#)gDMWcbVRVX2=d(_G
.C:F=#ER-?RX\(I_Td,=T.8aUG,-6fG.(NZf?YIa/bL<PG7_=B4DP2&U-AMGfCMH
8/RW(P52W7T)X]B7Z<04d#ZW?GJ.O@J3]NDDX@EO@gI,0bQ0V?,8?&N:>=^0f88d
:VC[S;1J2^:==T^=d)Egc6fC3Ig^:bQ,6]6;^e;=#P/<LW43d?<>Q=5@K]aZd\b>
-,8].8U.C;O=aR=X/,Ib?K4^gc.XELV?ZA/gFAe6RH\:X(MJ#)OfXAed69LDZ;&e
U4K)C,SK-)@NMR+d2D&\\XH7P>^aYRM7CdY08TIKED&Da>_a7@H=JG0b62<NY@AW
f7QK<P/gJfN9BDT9Eb.Y+c))ga)[?^Q^CF1&+]WOSY;2LE_6X0b]0Z-^Z\g8K<gS
YgW973;>^eW,R13Y>/X8d#6;0JV,RA+)_4?-fEP;+#G&c#]X58/-B2.e@1c)6N#1
Y=a8f2?B@CPU+Y5,[Y[PE?YK-6&)L\_;8X]SS\&S_&DTV.E(+P/d.#VKfFJF<_aH
>G5cgd#-VeVb(9WdYZJ6dQ>5X(FdT>g47:c=U[.a:ODUa<1TUdT&a.aNP)K[V:QH
_B(SGa77aF^669+V5,d.U5;N51K+QN4)7c2WW2;ad<6(X3g3M/;aZA^d9gPfWSCI
Pda\M^JMU7(58N9VG,_PIROYV1DgbeRZ8)bC.YTQE63?JKSO>1><La(.95:0Y1EK
T5&;&YWW_NV+)V\dH4V+<f/g-9[W;a8f;>:^[GTLc)ZG-JC6dU+I52DFPW?0BR_f
,QOCgUEa+PJ0FP8+EeQg-?)bIOC:-cOH5@;RQ199N8\^CL@,2NIfb9(HLN3W@(;W
JD3.L\aVf>)I(5cGH4NE20>f+AP?LAY>c_^N0>f9.:Rb2^\@K-H;,[H#;XJOY&GW
Q,3YQV)6:^VJ>3L\=X/6_?09,>T64_];7?I2c[@aT-YJDIO9RCe,S<fI,I5F&7X8
10HV_a.4fH86G4(1b=#=-Q_LZ]>@Y?7[OF3d6LLY;-b0aJ<Ma/DR+ZbW\MSJ6?f8
_E-Q\+SBZ<TBI^UI@>P9^[K)LCHc(O#]8aL_H5ZV?A4dC5_;0fAM3/aI)]R8S.-=
)GE2N,M5+)\DE-P;AFZ-b+gJT)#S/)A1Q)+5V:;NLM+7FeA,:D3.E,T1:V=J6OVV
aa9TT9+EGK-:d19,=eLR#CGTBVc+05@A/a3Y[R(g.e>-]WdDEU<P:[74R)9SVKF:
.gAK6Z_G1#E8Z7eSJDf3Ae))dd=Agfg?Pa@fG>OS7)N(PT=MdL2LZEKgQGA+eU@H
<cbEHg1/,\7XO5H7\;:Gf1],Yb:6)L:Z0C0[/3G[&VW.)3PSR946+-bXF>f;0[_/
I^&4/WU#/=(U)S4@fY0SQ^Z\+OeE;g]cdQ+48&Rfb+]Q:EaTOaZHD=]WKD1:4@Oa
OR2>B33R5V#T8KDNA/&^ZIL8W2PD6-K_Z[L?DKb2P,8VEb,HR1\CSgBYO#Q<.F:d
HZ:>LHfd=_9Re;P257ceM6.ESVGEBD<QSg,<#6TQ(X29f1[N_c20/g_U:g.^IC,W
HN7+UH=)X9J6I\,B3cQ.?<9c?&5][V4<Q7YDRH8D&6US:TV[>]\95CB2[G=>^Rg9
IU(5SXZ+:fgFdR<dVYg?GaYIa60WWFeOP2cI4XF>WG&N7bIE4U)+4H+2]LM6e?^C
Z:V=\ZU2M>JC+Re@P1WO0EB\V0DePF73>>GF(1K>^RbT+4V:gWe_=2ZPP+IFL8,L
&]&A[d,+)H8>J8>\a,8/fZ/YSbbX5a1AW<TK;Ce/(_W<A5&K4WZ.S(Q+0Kf_V5H9
+(d)/#fC^9^5C\&A/0e=7d=^J0Wg/596R);@JgJ<.5W(I+E&W^):1PTJ.2F;?S02
N2B\dI4:[^bT-f+>]#HAV=)&G=A21dB83MX0c/_T5K_2(6gaO3<DA)UXAf951a5R
I,)B-DW@S/RSJ+gF\H;-]3#dI=2eYN->7AR,CG>9Z3(#5f1JCU.2,AE,0=E5,>4T
2,E1UQUa00NX1C2&IYV?f.>dRCWPPSX3K;9MN5e:]_KUXYCEgU[WF(U5=V?\T_YM
;dd?B?KG.#QI(4I;c=\K29W\JIQZ;GS9<632^g4;F6:FagOWZP3J_(L0>+&1,&Zg
//(?MVdgN.5ZOA6(4A)c.P0@,;3--aO>KI.@J#CW(RDaI0>OE(/?)2Z5HPb@f[L?
Ba&)SJQE1(B6M3121\TUW)Z8TCDME:&^)gZ0A&TBeS2d7eJfJ]F#3f#?&&97<N1b
UYRB64=,.g3Lf0(/.-#,R4H:K#CT#DJ-0J^:,#Ig58+)7P+Q5SBg_Q51H4&C9-=d
7/d[MI(@c-18^^N+g@\@@)9DSE11Re:EK4(84/B+LWNe5XPQ1MST8H?^:1C#CF&b
bcH122&MS,CDNS7A[Z@W23:88W8JN?SW\6D0B-M.Za>SS&gXDT2&7XNNIQ.6E^@2
\A];2fDZ50A^.2H>=R-RZHgM(X\,Zb_B6aZVRf8^E7d2VY-A/5YDe;L&L2NO[[4-
a[B;0@5NSDU@Df3SZQ5]A-5G\bKOI#?<Q/KFRgWQa&Q93S55c]&VX9XTM)4Z[0I]
,NVWQ=0N70D4dG0a2.8@B34D[,A&#c)@_]Q(PGXdL&BCDdS&F+aOOd=;_O.8U[Wc
AM&X.Y6L/>[b01)ODCRW<F3c^9cDSU.D/]INbKL>+XA;Xg=d[c34gC_W;-MaK=QG
K2Yb0#=KH@fI@AL)V.^JgdbD98P@\->[0RWG.-Dg[0daOVB&^TH((Z9U3GJ2?7MI
OZ/Kf<C6++QR=/DJ&d-X4\I]]]N[QAeVAAT&\B=CNYMf7N^L:W;HZ@WS&4\=c2UV
GgfQ<RKBL-O0b@?C3GKVEC3?M_S+8;54NSV?VUO9@YVDaWE[)47#W_813>fT-B]?
#Y;]0/@Ze3KAW?X0ERWP9+dPUJ#PK,gC:+c[e<b:C)Uc<@N2W<1Ibb0IKMdD\b1M
f4NE63W[5+PE,&/A\NcX]]TEb)?9?QU.[8S&6T(499NNE-NOFB6NbD)03eJB?W:F
7[0O)Qe3fN1&Y<C[13dWO?O]4b3QD;=XB\DDD8K3fK466>S+Y1;I911dYO&&aPW0
PC7CaLCNIQbI+ce-0]PMC8\2KITD-0&6+P^^B[B@N8HY9D3-D4]D<Xb?d:B?&2ZU
]]S#TT(J?Q.f0-e4_O.V88D0<#L&K+?d@RRE-d-Hg(G<F7SIOGL\8cKdBFZd8F)3
Q9?U1ROX18-II4B^1BGDF,W<)<PLO+4d9EGIB<_4Z__aFWLY6;XO-MGX<0G[39E0
=.Ug_NQ;T&CT_4Z&fS[0M>M)R>Hd^,\ac[L@dKE8XKKDM,@_YcVD(BJV2\CV.49^
(fP4eBD2UPgQF5O4YRE1EP^#8Z;Za).&VYa_(J:065<,&G1@.^;&X1I&9/-296@/
^DSUE2UcPTC,>2SN0>A^CIA\>1B<FHYIVD/&Fc3V==f<XF372LN6HEb&6?d1H/<\
4697\&aeBg],QW#X>>QOZI)3EYNTB4g.GS=Gfa0#82/VZA(<S>N0T:[YbVG_HTQ=
-&62@_+#&ASNgcd6a.N_-#WcBBMRIPAX;W^K\D,e5R=BWSV#:d5T;\A+?:3]NCMZ
QbLJ8SPF>H74GAJ5OaBY7KMB92\.5A<&\:b.:E-c\fH)BJW.,f+1^c<X_2YPS)UP
c06Me:FVe8>\:J_+#XZ,1Q.#X@5IX(Q(1I,b\<BG-=P6MPD<>40>WAfS]OV+?KeI
K8HXD1RHfLc8<>HIP@NB.W<_bceD(T89]]1@-7EeH]ZA_&P6OJ=I@a_76,fcU=Y3
-^D-0I\?3D316KUdWH:g#=eW@K&S7S^CfJM>XcBbZ_e[S=.4:f@@+\XI_]>4/5L.
1dUXe[ACPeYW.D91JF(f8>?77XT)J.6-<2J>-N+f5<PbM7_=4BHJK0TUT0T@80AD
UT&YHAULGQd332[:))=A@@F4/^eEY1;EJWFa&8D8f6VUEQW,)3]-gRRB@<J?6[eH
Hg\)b9aS5g9[C[?@BJ8Cac,HRRQ\SD\7]R6M0-5I6F7ae,a.RT7CWFT@71OcC>^c
O&V7bUg8gX<4KdJY/)T6d8B[^0X\Ga^)9RYA_,^KdI1\WID42VF-,HQ]=:&RS[#+
Db0MKf._QT0ODEEgJbN?SPWGO[b&aYaF4,b(8=E95[(:>BCN+56LV5QVTGT9I9Ca
DBLeGA&Q4HV(_:0^W,-/C5da4K+SX0&7AMLJW_ND8;g/[H:Ae[G?3&#H0<febD=_
[=OQ<\J&L[(a(_Y/7c._(+T[&F9LJ48cD,b\_[(_4NVHUQ;b95OAKPfg&AF^P^7N
b_aCbf#CHT[;P7,T,/XCK+Hc^0:]HeK0eZHWMR3B?8eBFc+0],fUa-Ea<&<?)COM
02??0D-<,&0QUc[@F:C42@H&4+,f+M1U_=#D;]ZK==XV6Na^bC7@.O&LRFZgf.=#
,gbD(ZM9caeO:IAIQ<@S?KcF,P0FFY^:/P4L4bXHAF:+]/-=WPaUP]CU=Y18[SG?
B5Ye\Y=4RB9bR(/5fJf1/OGXA8-G9U+_I_Ee3G-3D>KQ-Y[?D.aKZ^fTCT1[,>a3
M=/W./+VZA9K#,CSQYa^#35[Z6@a8^Y7g0@UHIL3>?c6[)3.1SH98/?AaOG(VUN:
cE6ZL-aCFdT)IR/CIK0_gS_Q3&7d>e>=K3G;aXH.]cO6:1NffVaX_.5M1HY+VcbK
&(E7NDFbKQ8KD^ZRPP0N/,bSBf3=L<DRMHHR\)fNZU[:,SXHOTBG^Y:20\&6>B9V
(PVTQcL/Ag&5gd7&Q,&BNXP?UT)5A?/>ZUL?9W6^K5W.>X/FQCR@>7(IL;K)_J;b
_0.?dLI(Qb9&)[1(NgJD],><2?JegF@3>2NL#,C.DC._K@bE;.N5U#,[_<f.WZGT
R-UbXN.PS@5B_g6U38L.)^FbD)GXAd38f()<>D@0/B+))57O@f.abY8G^W?fc]#I
ZG0gQU]=[L1YV4_\I1242XF-WW:=#<+0LLOIIS+a403M[3F#)KNX5c-.C+PAPFO#
BV)NO68_HAe0;MeC&JIXG[INF3AE2JEb#B&71]^O344Y<G6\,7-G?Ob7@6Ke=,KZ
KA81:01^:R[Va#D_<LXYI0G[V#05)G^Y<>#O=P+SJ#PQN]ge/XO1;S(LVCSPN#;G
@fUb))JaY=NF5<0(Z=54-W>+=ZNQMY?0S[M/EQZQ>1:d+=5cFARa-?R3..+?gCD,
[.fe4TT&H;\@VfBI;<b]Ke<f5DU;U&.7+\LP8WU<);9YS-2)6-RK;IZGN;3\Q7KH
[gTD8KNDLa\I0&:]V\?N2>SUIXb#(/[/GfW#Q;V<1+F^PAGVRL23D?1_bI(FDg77
&.3[BNWdcVF->KIaPDVL)?0FAF)KJ0G9cET&;T/S4?<UL7\6N4ff=g85)8?L.HSF
]\:b,PGX@[g,-WfFMA4d@aC5S.KD@@/S([:50HT7+_G[SRD<]8KDL[MLT_#U_0?I
TK+9<7\a-1VV[Keg\3OfD_;TPg9eFYbT,LYRfRdQb2+,eSIg]SLE#E_-;@=X1&8c
>)BFY&STYC^--dT?K>-#1A&::_TCY0R:KNgfHS4U+Q^0/+PMA6L@Zd,035cFc>TS
7H>TE+[71YfR0L:S2B>ZNP3]LD-SSC;XMCI^XIR&55N58;0&PJ,._[Df@6Y#?Y@E
?6cC.dHU4?:16D3F>.E-Da_#>WD.)Y<S_0Z@<fGa;0]AR#\@(H28M/X6?5GH./7S
eRWHJZ>FQGPZ=K/agH]-#7J18M+:UKeP?T)FYAAI=D)GE^U:1/KOO(c]2^2=URRH
L>#A>C3e9+e(2\ROMcRKFR3G8@[D.0QKB[J[f]RAD&_F(/72gDJJL1e,WP>GW+aW
a/Y+IeJ-cU^U6H@[/bEG6WZ:e)###81#3OS=cSJ3Z[WGSC3eQNe7?VdC;4V^>cU)
L3Q7\5K4@+1BB@_?)KA(8?;4MMLYN^89SM2cMQ;];^,#Ef)U[deUR@F2N?OMBd02
6DQ6;@(g),2gG>8N6ZH2(.H808S)(;g]_e_3;C6.g1^KTeZ4c?N(]C_>41WBa5_?
R>@F[DEYHLe<,cT/.b(XBRLHgZI-\-MLMKf2\NS#_KUMPJN4dgBL)YJTO1E13)IK
dRU2WK]WRHSJHL3b+1:BK6\bg@C]W]Y29QM5dcBU2YFY7UK@\&OB7,H-SG/O^#J,
(UMa)PR,]7S.67_E\P=5WL?-F-SZ??4a+/YB=-H28f=-DC\)4[N.9EP,E9P8P1T1
Af3+6PSUQ,CL8DYdBR:8>+1_3YFRM^8SbS>>K6=[+eK]GTRg^S6gS,]P@77QgHeE
R>CNe8G-+7gbf:A/V\9C;a(f6X)bfO]?Y=I+>0<PD><3JNO6:Zg(RaO.H7CP7<GO
aCf\E64.(dE<#^<;Y-L#ZC-+#WAM1TRW#8X17>2bJS<Ob(IMH6YcZeCAB218_91>
P^T(#CK\,U^QeJR95O\Sd(:B8EDZO8Q7B.cE(6Qf=Z,>E>1HQBGa25Q8UX#V]JWF
[K)^;F9<P28T;7B]fQ^@JZ2FA/K>UF2&0_9+8):=)/LV^^L[dMM7O+-+2A;7-0D.
bb^,-EZE/_0/J027U?fB5<7)b#7U]P1ebMN58;-+Z-GE08]&W0QXA+P@#M^ILb/<
TI,/C<R=+Tc2a:=FO_^9]J8<H^Xb<LPT_ZFOHc9g,O4:^Z+Q+J2>OVI2YHN<:eLV
c,1(=20dPQeca9_]/,g5,YL\59B5;c]4R=95=)X8-c]P-Bg3G7.U5b9EQD6/?<XK
5eU(+UIB5fXg&:MbQT0BBZI7(fW-?Gc3EA/.MR)Q<ON\N8d,(Af7;Wf/Ub#g]J<5
0T:\8=^eXfH,O+YZGc59df[d6AG<@DKCDQ7IQ_d])KVQ]X[6+7X0L4-64fc@-86a
]+;cF2V=dJYR20)A3dg,O56cP@]A@9f,,CKF6PL0VR=&G@H@6gLDF[dC<LD:UNIN
?cBgT@>R2&7C=-QIQdI>CF-SeNPDgVA[,+eI47C8O9)+B]+C.:IQ+eD^YXdQU(Fe
<7:+E4I]KXR7W7M/DecCdY.F?&+7[dE_X@CUfc-cO2/S4VQ\X3VNZ6L.H;DcL[UA
CSe0Q\:3V4UJg^Kd](+-FLFK@_/FNX)TS2>WBFK_R/NP,7E^Z[@cM@<ADH0N+3FJ
>CIWUW_)E(2HX[aUc@TUc=(I7aZL3ZM/XQ+/ZU4JMgW:UENAVF3KMbK\]b0gWK3a
PD@J@I,QJc5J@:ZBX(D.,K<.f/Y.:\ceISQ7c]cHSR>Zc><=03L5+<c.\QNB.Dd3
8][A_W)W/7EHHd?9MP[/B>0TL0;KW7.(.QF?L(eKX\860a,@>9/WfH67?bXZ0:8/
&<CXN[T@/&/+M\^:<Rg2NJPJ-DCV&EU3G^@ZVY8B,#U,/WaZ.1\T->\4)CU\2-#4
\fR&JdLT#1VK)HTURCYO/(\IVJ[_M?IcW=4T2ed\f>-CQ12,@L=Y>?S]fFY&:L?=
+O+QY-Mgag#ND1)C-VN=1DfDYIZ)PV])VV]1Hf:b6TcEcN(H<L<64[+?J[8aO[g(
0_eR/a=_Y[QVEIYB(_UN#.:&V\97U91622[_<-N3J;UZbF+Fc&6HZQ,0K_I6-CJ9
fa=37QOd@S:IYUPL>^KK64,AWf:7B=.53RQJZO_?YD=M:8#F302LW7<cU:#bW(]E
NQMfT]P><bZH[TK3SgG4&SXa+^VU4?3WU)_6(3^A[W029BGDD>RX0SB+KTK@N=+=
c,ZV@FNWf:Q[S#A05,G,N.Q1=5[#PL#NULNL<)UN7aXd#AE<(a_(M2dF>H@A6/8W
HcBBE88XTZ2P4K>-=R^)LgaB/IGI^0g=V=cAUXA7WPEARAb])L8MB):-_)MCfbgI
L78b_?gVGLTb>-RcVOP\6BR:9:gH5g]M&[6^c#6:G#EPGCX9I5T1Lg3eN([(-2QQ
SZ#Wg5X;N9\TV?L_gMNW5/3KK4Y12@fF[g4a\e+4LA18PS+,XZ1EQ9;aK1>JLZ8D
a0bKWV\c1CBEN.U;>#_-MO:YdaN)I>R-d>)4VID6G(4369Ha?>;W18.#JGPf@35J
c\=QK;f^?EOb-5N4E]/<GY[QFL+]I&#8,-1SE4S,YD0J)f>L^TAPT@PTe6>\_]A<
E-S]W].>)]U8_^a(/PTX.]+)N&Pe\6_G<_/b+74GbE#^=YGNK3XXD&4OQePU\Y-?
fFT[.O(;95O#)Oe.Kb;0bV#3.>Y@7#-;bL@N.IW1#?X2FdbV4F75+XQE<^72d_Vc
[EA<]Q+WgLB8JT2Z&6#XCF_\bA.D(VJLJL8KQdQ(N/3XFVReTa;Z/(f>/a6HQOT^
_fY.2FO7OI?86O68.X9/AZ=F#7b)WQH:S^dD>NN7JE+XT2B@]I^f(+Q45HUC/.0(
EH,-^fB71:.F&/HF;f8P3BJ\f\eZELX5)W92GK/d6b_?9AL)2g>eNK@?Y(>B?MS-
K0M])KAg8@KUccF?c(fBY;XVBPd.6AfTRU.G;W9JZXBKDa6G)c3D50UGKd2ER]^G
Sa<_e@H2eY(CB?&?S/f@O=7:5b/7<7b7OO\4EgWII2d4C<#8:VUNIO6D=2^YFK<B
?T_WDNN_,6=EaX8M;8)[16KPTgF9T#?=X8T;=c1H1B=+LgXFKM<M0N][U6<K2G=-
:B7JKC?S/J9fQTQ)V)Bf?]NL=A@cOP].]T-2<KZKeEN\1b9,Db[<0[HK?Wad+:]1
R+N/O/J7DGIFJ]bH4#02/7^R?TdTScQS--[g63DTIAd4/@;)=C=9KVW0SeKL>@98
PN1VKcT5>^5_)aM6M4R<9ac=P&Dfe6Hf7758T-2X?V3eHJ\87V0NM/?Z+RbT0\W2
K4.IMBYX.H4Uc?2)4dKA&Ic4Nc_HN:e6:@IN:dT:F-QH(QZ[HBPU7E<985YHe,A&
CHW^42JF4^Ke9-/.ceBEM855V=95L[f3L11eAHP#<KTbL9E_#P48R_:R&EB^QDAa
c[4cU@gE(X5_fT//BJ;3V6NKI9MC3C?[VD=GO=&cNR-JRZ/.Q0)]GO(3V#@.)]8b
T74[C#ML^;c9IbcV[bBgWKa+1[g2E_S0Ne19X\d(-eLKf9E-I-Yb(3-LF50>HMQ\
:5;A[EVJD)[EU_5(CCPPU)Kge5^\<I[HIE.aXMe1:BXL2C#.]gY\-@_1#D<e#VH5
E1[L2XF4=IR(HGIP6Rf3#MM3=UbNEIFcU&d+ebZKBT86@?WGT]_eI0e9WTS<=]J8
_J9<+T4QY=9121RD)eS>@)X-9,\U:Y(\,B-#HIU]@01aUI,XF/BW79LA&\A;T:e>
PJb43A;_-T<GQ=PO7G8(4K)HD//gM[(af>=e&/-;;O9F/fVHbQK>6>XgW21\MPBA
\-]K_M(7Y-T0M3K0E8bQ=OD921b+c\]I5-aV_TY1A1\8><G.eY/7a)Y_^-WHQ8X=
[O::Cb;1TPbT4bTJaUH:)f0CSO9DJFBf:P1<ac7^af/S+@Y9B]OYMaZ\1D.CbPHX
D<cP].8W-^S-HW,ff6cSMHS=U^PR@DJEMJ:4\F\&-?cGVRgb_3SV8]d[8FMg:H7)
9A=BbRfSZc503Y.IfD3Df[;4PJBUH@f;(+[7Ue=KcPgMVXM-f:CNB=75[PP807,.
/^R=RF[4+Z(a8_XEL<[Ia4O]CH3#+HB1FSS[90DgCEdZJYQ[)&UeKe#8B,Q0bb((
\UW_X>A9\UDQ>],N]VB5FM,71aQKdR6Xd+C)a/+\=<-,^F55Bg7cWA77R16B/PF]
.5ILeBb0a0gZ&PPf2Z2d0&26+N)RXI_0).\JR&_B;UP>[UXFFSaY/Y3adY9L@ICB
YBHI20Q5gY:WBFZ((?aWdW4L,S2_ISQEa14]MZ#>K]H=Sc>1.@O@(&8bRf[83f5P
_P1e<)R.\>(gD)ESL>9J)3U:gWRe5=cg0b>2RTH3\Va5SUgH^-ICS.^-(J@<2]#3
6[8N:&F=#Dd2BR1VW_UfCQgIeE+6[NO@^6[PB#WUE\5XTAD=NUcK\2R7XG@6>eB<
N3Z4;]<F>3J-&+^d4X=f_8a9>8LETGANI19E0OQP]bXJ+(3Kb,a)<)HeM7P),[EA
H6IY>+-27bSRZFO9I_/@>R5#8bA4FZ#e1+<9D?NMN)IX#7I#K7;DN28b[3c[9#ZL
K]L=X.g[d#;:5VQ]7U5?Ve7C-bZ.cK^6#gV0cc9P8YOAP[Se\>1NFH8[<D?;d6+9
O]R830+?\YD74GbSS?AB8DDJ.2]8X#I>fa8-;fLGDDCQJ5VRR#d\MJ&/QCEWdEb=
PZ1</8g1K6AJ,W#=;FG(&BWa>7.YE=6OWE.Y=AcAPP>QW_:8MWeH_:\,#.4ag]6/
NI(Y[NRDWFSTgb8d[)N;V.:7+B)<:aN2QcWMaOHQDJ,XH.\I<6#0fdYM4:I02U3a
-[()/7fK-N]-dJOb\?YV^N71BBT^3N+?_fbO+-UfedGX\1/ffTFN>;eEP#41cU:G
7dYA4VN_L0A)O1fI9A>\;+AQEJQ02CP)=g):>ZMHZc=2aC+Ud]OK;F-G#Hd@RTc_
8:2RBD<4N2Y9S;a/YJBfIT&FJd]?>PS[\H60Z-YRd-cY_Z8ZNGI7g_CS(5=Og3M=
UM\?DU-Je<D?J-(Yb8H#;aRG--T0F,8C&dQdE<6-EdAQ.<N]50K#[dN0e?Q-aHW,
01JIXG6NFL3O(=))HJ:8bT7#F+668N3Y4QgCb^.Z>Qc>B34=)<2\A?g89V:6LRNA
=NS1Q(Mce\6C\+D@JNX+X4CIKf+f@M1HRHIg+G>U?H^:\[)X&FV_O^OcD?R)&H3J
A;-;1ESc:7LYJ4H0c\RW,#J<f#=+((cN_eM42=88I/f<>1V4]#BR/_6c+c=IC<B1
;Z&JHEKgG)#ET\M9+)g@<b8I_J&ASH.OQ;R(@9&.c0&R705O>g?_2OGPF?7-WK>9
\_-M3;W))&+AaB0RD6=PB/aD3b8KU>5B\7O^T?f8/N-\?5OLcE3(de]F>S9RdHLX
@;:]IN\O]S<b#C48LH[Q8(4W1])?LfJ9#);PXG+UI0+Og,e[\94Y\GSgPJf\/(4,
XXeDF>7]59&K/XEGYD1KIK3\G^L_9f,fYH;95cU3@ANFEC3c7RWP\2U6VEbW)Ld0
7,3-V#-4?C<E=1&9&(&EI85G]5II=b\]_TN3]SI/=E5,PU&0#)6UAX9,?e_KEX^R
<L9<e#[9ZDP54Fa0=ecC&LV9L+H]GAcHZN0LcFaL(-O\[[,_4I>_bb&@:<A1^B;[
\\Q;Lc3d,Z3JeG.0DQ?0@c+9N;c4]Wa^PJ?;OPRe\;9F-E]2,/1&ZKO=IK4?b8CR
9X>X6R3R2F6aVQg4KV8)9S&S[;DKD@;W&.3N1DNN2\TQ#LKG898g-?/=57]CQ7fK
=S_=eH#d<W,?54?e5[0ERc\T&C;>cJ,aWYUa<ZS:()<O3CG,YNK9/L=@XQPOW?aW
)g9U/44?0>?@7\M)M]60?6_51X<6^fH8G2M2BZ3bQe]U<MVdWQdDWg@WE:GI@#0g
H7+e7GDHg:8bcc)UD\R1gRLA1O934I6:95;E:SQXSGB0dOe/B.-DO1EECLTC&G;+
?GCd?4b,Fgd4e,7MX=Y6Z=HO?C:82IC)#K>)5GFI8L(c1UPL2^3D\Qe,_ZRAY^cd
;gJA,d^W9L<OU[(5cX+MP(_I)4V/d2fK&=cB.ccSNUYbY8@>HUU<BEb0aSVS=_\L
<-)F<0))39^gEW<MC?eN=^MJ&]+CF0aYI2eO6(Y(_CV(C)6@#Z]V8+eHZITDB#0A
7MKK]gRB2DcC._&Y?W;K-1YD7_+)9\O,b,V2H6(b7WG.]9,/e+6\,>WJ.+Y,FIOZ
^WW>bAVHY>PGSfDZ:[+K;)EH>>4HD4KK#EQ()3WW?RR=BW83Ibc;RJ\eH#0A)A3)
L;\X4NO/MOGP\<1AC?I,\Y:>;c.;161(M9.UKFIH3.ARL(]A2e3=LPFFR\P(Q1WS
KJW=9GLL^=J13AG_a-L<4g2Mb:Sb1e4&C&]:g8+3[;F)XA#-bb7RQY,?O5<&C8ZK
@7XXeCb^.]fSWX+VW/^gbF]QE6YJfE5K#0=E<=JHcW6.CZHd_WLVa&E6AKU[ZeeE
IC\@8/L.)6a>^Q#F_ZP3eOZ/M#E4-D:ZHV_R@ZS9[QZOSV;Z^g.7EC/QJ2PUW)LY
N1?KQO]O-?#SIKdKZP9b:=ULaLK8X@B,C#-839://=(2;H4:[-,[7=Ac2F]J?.K8
K5e_?IGb\)fOg_DUcf047F/f4aVC#V0M2T[+@DHCMY/e?X8/&P;\;@@JCX1<J:8<
;cP@YH_&d354<Z;G)_:2W?(edY:=H&,VGKSCE9=,,3aeNL^cF75<f1Q+R4c29J2P
IeYgDI_?_.&[Xa8;ADfTP;NTGC^N3LA\[c8G#0dW/H@>;@F4FFHD9]7PUf;.?\F^
^W,PX(F^O_)f(>7W;\9-+Lg-Q9:FKd(a9d=c+CbQ1T-ACg9<I[))NHCPW,b,14Y[
3+L9E6B7SBg>MS:)UJLD7JYV[^HLK?J.:;.L/bB/626UHR\bRSg&;P@IJ@P4[V9g
1e=,Wdf[?\d:Xd<f\_Gaf/Q,]=/9C>4SSCfEEdeL>LS3\RB0;2QY\;V8J>G[E51]
YP5V+eZa^][)461CB+4gFPFW97@d<CHW0;ZU@G:24OKIR;B6:].f2fdX&.)_#E^2
&EMC[;7,L7#\Zc2KUAf8,&5VR+9YZY20Y&YP_1FaN0W+<Z<OF@ZN,BM2e-Q]L>&8
8I24C^69MCFKBZBJTF1E6GH+,O0&4QP1(?NJRW/S()FRH_Y2KXLHa\?SE]WXHJcV
O<cIDOG<WC&NWIB-26L?YNgI7_^S9E1I,b<=>6T:DEVMDE8UGNd_M_\MBX#Q8a\;
:8+AYQf5d;VY40G=3J_2NaB&Q\<d)5ba.B[G/PRcNA1@.J8CWGC]UBa:8LH(Ng=e
TOJMdd-[^#g5_J#;LT1:1#HBf[:U<P/7WcU4S@@ASGFAMNJF_&O&@X&.89?=>&YI
(XScN\VaV\3NNZ7Y:[RBW/HBY8O<5[gDc8.-72J.cPNQJIaeM<@#A,W-SDY[>\3F
0T-GJ,OJP(6:?SY)CY-eZ^KGADZeA_Z9,_C4\D;789^A@<ZGY_W?U-=,KCN=3SB+
]??]/5=?5#9+2De&eRXT0-X@5QP^M?J_c44[8/[V9BCa6d&S-9Q+g/>T9@/a.U>5
A@.Z-S#C.130:^BCTG6U:SBe\1aTVM9/>:e.02BPeL&TI=-J4..I,DC^^JN]b?d+
cR((f(39e41/87.FV[aFPWcX^[(S5(DU=31UW-f^0D\]7Ob8S9/6WZV=[R0-:SR9
,FKLS/?R.)[PZb7Q_8E001A^]1R8&Y.PH,X-)>+6R:OHFc2T;8#()\EMA<Z+W6K_
YZ:L8:2T1>X3/1a2S#a)ZQU+;VDS(_0@f=D][9f\.X41,)McVQEF:?1Z)34BOP0[
84f#,Nd_YQN1d-cKE6eAZ4]G@X@LZc+[TT77^Le#eZ@/0#H(4UdZ@N:2Nd0L5J>_
MJ(P=N>PY\BQRS+HgEI&_Z4,C_Y)ZK&@?:@;C\2/=5Jb_R:F&94/YH5RSDOJG&d]
:Z#J#-HM@3JV&H_d_<-:X5d<(6..2KK7\.eM.Rg]:JKH(\/2:S.J,=3P,bI1dD7e
W7Z<Ga@878_SCZ/V4CXCL398MYcQKALH0MccP]_[g7FJaS/?(/aR[-RM;D.]G=Yb
(YKQ..PLP<S^WR2+Jc^::X#/,_D8];)ag-P8VJ7IE+/Y(>V:W<WQ/BP\>Y48\HF.
#TW+G2]JNO,MJ)I<M8EDQQ,4_5:^PQHdCe?RcCBDS=Y&;3eUc3NcIL9763Zg)\^F
afEJ?X[(&\(JJ>_?EPQ146C<\LAbG]?Y+bKdeYe[Z+(U>b;Dd.MG1RIQR>S9L#d(
H.(ZDMTJ;(W-P66/g:,4bHD_L;dbF1c7/[00W[E9d&8ONIC5OaKXXIW97I7-^/I6
a[]2BD[,4,X2bV778fWUTZ?B)8O3B<e_\^T:CHG3(OH4b5fG=@M-8;)R\6ATfG8;
TE(>]K(\:,=f#Tc(d1E-<RdRR0/f2O;UQ_E1IT8>Z>@QP=d_F\](fXOP@60F\;.X
VdW9/;>I8]Y4A,AXPQ>\4X7Ca-O-4cEFZLX+:XD3_P7Z.5_TUEA6Oa_aQ_GfBELS
aH\I<NP(U\^9D=4)>.^1WF898M9(5Q10ALWV/>IZ[O:@C7@I[.3A:5.(D<&0D3Xg
\T2Qf<LFB6U6+YAdf5Za4K9Re:?d9/OJ.[[_4UY@QdY#5aE#R^+UI3P95I^2:ead
=/X3b,b0-<UCfD6>?/3Acf1W:fC;.TUA]dK6aW2AA/F5a00=NJOL>XIL_\A<2FZ5
\@,;dLP-XQ9)QcZ),X/-O(7TV8\X9[+#DLX\5@9X&e:4#5[Od3TV&fDc>5:O<4H,
I@=ObZd_c6>R/G/7gZ;fV2g8dDZN&?Qg=0OP5FE7Fc\b)VUR5-:J<=^c4AJ86[3/
Wb[?+c[a&d5ON)D(VRH+X#YWO6,\0]\I3Uc]A+eF8,aKA>;HfH4f.14BFBA]?M7]
(G58e[3+T7cVSO5)cL&#_N_75V_(S>BE1[]QH&a5>=-RE&S<U)WR;L-]IV4)9cN(
:UMNeASL&UA.B_-,@)H)Eg5Yc8552HZFK\ZX,L.(/<3g3eL.@W+:_UWN7MCHJg?6
\SK5+.?VNJ0(2H3<,Q@[)WYT+2O5_TE^##6<T&W<Ad::RN4-VR\(Y<]8;>8e>&7f
:?B7Lb.@R3J]#XA-)(Ng/_>f))J]d-#RFO@6SReEK8Vb3_7eP5G\cV&[;^P,>XVI
C?/b?MF?-^P;0E7bf=R\89.=Y/8,V_CG)d]R3-@IQHE.-TS\cMP?,L(Z&CF)[A>d
18<24d91S40)Y8JU((:gRL\Z]eM[B++a)CWB_K0>NY]d&>G.:HSX;5Hf66.MDJS\
WEI(K-C2SdNHT@ZTEg^J&H;-;7#CUGV&b^)<9FRJ_=f)R&.NeVK/&3P\_##^(K:.
/&gPfQ<7S-.NAP=/+YB6#Ha=]6-=,-P:KZ@)BD9cBfN2;fKX839OZ.A2;#=KOEBK
WI1K\PR6+>:._:E>6<I5+QdN43MG@<=4e+0b=S5?OL0JX&Jc^WTX]U@d,@<SBZT#
-X,E;3S@27L&FZ,T.@9@;d@KJM[^0_JVE-7[??gf>RB-]OZ7cI2e-?GDe8_@:Q1g
Z]9P._d^XdOc)CO?\PDT:d>C<.E=VSHV.95:M8>(eMOH\/W8bd?GPODL&(-WNWCA
.Hd181Q=VF4Q;\WO:C#T.EbH(CeE.OFKd/.FOAI&;+&6<2+ag?KdML,BBBP8cIHN
_I\9?+O)X8^&.WZBbY.7J<V&U3-fHf0\/cF[ARC29\9?\H62_M&3IV<.XMRJUN3K
()^GGEY0\P(VYJ]EU]0R83\AYf@EQ8WGGcDY65WL@>gW?G1/N[[^.K7eJYK\fd.d
R4gVW(c<>;^7/WZH[OKaObK--EW+Ne1W9BLY2cD25g.<&PQMS5PB\Y>F0TLg2Ig>
g4PE?\P9,9S2L)=NU&:\cfb+g;[d=e1<<JO^OOMO<HDeF2&1c_/B+2R6RK<X=L>/
8=2c,F=;GOM)FbDHH]0,_4[[/cS1:c,@AYE+Gb&_;NP+6(W+5,:G>e>-cY7MX0(2
12N=CgbB)6I+]a3Z)DSL,daIbN#?W=Eab=J#-1^S\H-,9C)OIS>ATHgWUeX\YYTT
fgU1[gJ)>0e;7;N22QL]La+/gK+M8a^9g\U9ga(Kc5aQ-G5KAI:+FXS9(cFf:L\:
20P_>@DXOBT4PP#5ANcCBQO@11G3O[2C)gA<P=OUN6GT<V\6&W+,#+aX<.AV99R)
E6+9>B<LeZEE544a-cW^X0>RVY>BQD+5g=,\gY1Nd+_Qe<CC51VJ_D<F.,+R8>.J
DCASf<8:C#6)P/fZbL=U[G6H2)Q<J9[:K[OD+gA-MXGLI::R;QZD684OA@XV(RO3
Y13EVL11?\1,&T57XP\:-d]MIaQ6[-.4[D:L?L9&b5+75J1]EP#,C2T)>TP6@a#H
?[V@^MP&S.#\OMf:WZ5VeZc:6-OL&9:eST8F5#bYW:]+S4YY-PE4#R[]T/)VFg0P
CeTO+]=O^[&_BH.-S11@\fTQYV_PBH]g]+@4db=fFL3QBfTeYA(WR6QfI1@4Y9NC
N+76^1&5DJH^<Rf.c1gKR?9X#)@TdY[2#OJY&=@51#_N?[JBM\Z?:9EHa)9[+&8@
:-7D1VX<,/,5@>R/-#5SD533_1MA\PaNCA8,ef&_IaQSF@SG_(B#J\O-W<EK@M.H
<(H^1G-eP>c9S)CbI8AJXf3Y0?01?3P<YV,^2VE/0(=N6S1&RR-^]X+.b[[=Z2gC
,bB_2CMcbJIZ9\;EE4I^K+YZPIPICSZ0[H_N8Q1gcO?19C;ASA#dMXY6#=TgA.?1
LfX)+BN&\?_Fbb<IC3De0(Vb+<1?e:&C2]8DI^(BC0Cae/#XeHF3##M@-WT&5@64
:WQ]Cf+1Lf=,Y&98WaQ#BAV_1bfK,6E=\XbXbfVBMWQJ+FM#2R1#ZB-H739fAXON
KaOC9NdDB-b??:HQ-OY_I;3\99/eVfHe-,N:OS[H_]=/XPgYgcY/GA,aHMYX@^)_
EAMad,EO&<7ZAG2,&c=0@.5PB;;L\dXbQ>CKa>_4N_EW;V3(#R\RMLU(P_d(<af?
T]CHb2WGE73Q@QPc41X(2/2QG\Y5X)XPb\G<W4LI&/CX@)[.K:B_aC+@WW[U2Tc1
6)X>>?8([.4YQa0-)-D48Q)e61Z1_I:CL3+6AZKgAIFSY&?).Gg[.EJ.R=^g)II\
f&WNb_JHH3M)Bd4MM^R67N08=6D;>N&.?_N:V^-bMM)^^8>>beBES#(N58OIfX?I
+bg/^Y^_+\E3I(KR@<XOX=EMNJgR>:GcORa(IAG]9K44XRB,HV&UPAGSMLZ1EC7O
NFLV9L.X9#F?bH,P<C@8M(B;TAPG[+75J=17WSR&5_LPbWOOg;?g74S<F9V]&fEA
-e>2W^T\5MALAeBY\NTSdO-#42N^?:-4X)/+=1ffC)H5_SgXe]E=gASBQJJGd1D_
Sd@+GA)76a)Y0]fJ(:,,8#I70f]AKac5be]Wc/G.g[#+XHQG&Ec:8Ib^H0GgU[0@
G_#,QX7Nd@M?eL[>VT;65<Q_L<Cb:W>Ld=Pb.eWM^6b(DA2D0e3:4e\X;__FNdCF
3KUM>]Z<b@f=RCT3X=GK,MHCIOL=eGKQgc?DBAL8=A_Jg9;S2WOaSO^(-YX[/JfZ
(.Qd3A?V7BQQ4QA1)f:]bYRQ9/0-0<4)P@@D\\4C?E<>+3?3++?H]E6)H\NbFQg]
F+gb(MJd5A]5H@_fd?RWgD<W0bFG[2d\^X0Q6?.71TD0XWKS?^Z>cZH6VIWR71^]
Q]>]Eg>O3<>2T+<U?eFbHF.:SAfO^<Ha>,H;K6HYX;V#9FS=1H4XROC/(/_&A;?^
KO?gH.LgH@g\0f/]OEc34b;)A848Ua?,]>EMTbLS_?3DQYY#J41B5\DIO7JKSObN
Qb()@1LZWMB_b5,dI.PSDLW3AQ8deebAUeZ<Sd@<)-J:Mc?f,B=/ZOY6])RC_]I_
N13L/LA(9&=2QI6(TggN5MX7Jda&=b]IAdT[EO9A.a.ca[;e&IT&gE@+BRJ])I^S
@0[?H#-&T4dYUBKE4/CG;/FWAN.Rb^Q4WU<^c\DB&aB^<CbA:.T<.CR\dO#_/4c&
T>8d(Y80<MT:06N0,O#<4S]AMJE_>HQ:B6_,+V=[A&<157Y\S+JX_VL]=LOQ/I:_
/ObYR4_YO5a_M0Bc=L[WEJ@[1cRJJ><=)5J17QK[UT)ROJU[0P=:V93&:J^T[gTb
FLX#=@f(6XB,FeINJGb(X3C(>?Qc-(S><X)V(]=a1QN++<3NV29)3=8D8MV&D6X)
d+2;<=0A1?PF8Yg)T\NEN[/bNg4KN7X5e.2I>EYDf>gZHW@Q;9aFOLQH_>5\.UgZ
HK(J6b3WNZBQ7E&=(E,_YAR,[EUFf2K/M.)9.&4dKT()_L]eM9&.KW.CSW?Z>/-\
82_L1)NTSY<[B_:B^b4B98LQa=W/KMa6Y-=g&gdKP4@X,aUQN=68DXXdVSC9=@;(
)#g1I,+AcI<&[A7F_(F_2?_)^2e&5&L<I^QN,<3)WIKQZdO_>YW5Z5X1I0M.bFH0
/gITF[R^OI(cRNV(Yg:4g4Ig__@V>OgU54]?eCPd=a0JA(34-C(O5GE\bTEXf00@
fT?LRXbX1UU5A(fMO]4e2d719A:e[O5W5ZBKH4f7&3a(.?K>.#R-2Eg-ZQNF2c66
K7MQdE@HOYZf0dJ[Q3CTWcPa020<4I&T0^PGd=7fcG@/&KeP@HOQ)Bc5S/142-=/
)Z)ENNNRdK@dcDU&:8ge:0Ac7X#OUR)QK>LaIRdLTLQ>4Me2KY9TV,8T?<,;&[7=
e.T55c.C<?F9QL(;g,]T>)D7Z]e_0b9]II\>Ce3U\OL4[ReV?Q0ECA&]-6GWI&2+
8V(Ue@[BX<=V164IES+J6[,1_&)S+)LU=0XT08+ESP,V.80^8CIJC^)?2;,VW)e7
+>OEO/0Y&HaI+^9;3FCC1:0-5/@(6WTXHIYaQ>T;e,7a:>V?aQQc41-DUOcN;-;#
PU\G:WOGE/57I,&e1W,?=+RK1TGJ3H_\I\O=BY0KeX=?FEM]<H?FbUW3A?3WEa+g
IXS]K#OQD[Gb_@bE7LCMMV)K1gYZGUFJN)1+e<6=DaRdK&+C7A1G^4KI=(APXb1<
d477D1]\??2U:0?3<=Z7O4@EU.F)ZX^?=&#@\4L474,O)FAO:Q0\>QW<-OD0I7@@
IW;NIX;XN.O03S+)NEFQM=(7]RZNN65GJIU<N05;BH>^IVgZ>YES;ccOI_QHBNG8
HddEGCU5PJRLeRLX7YIB<H]+8@LCKA>GA/7Td7-)W?:^5LV:B_9HSgMX<=4\SA.]
8<EdVg?B:?0HFH]I&;FA^4gAfT=_6:[8M9O64_cDY[R;N>C2@_8&egT)A&P]&TO?
VVS8If;-9Rgg]O44&f7JKKOQb,=L5-,da(@_KU+#L4Ye^,P92T79)[2P8LJ#NRB\
T5RMDB7S:c1[Y[L(L0gMCD^J,93F77HE6f..ZM/@W#77>W35NH(M4+d&D1MCXE6A
4Q<7MF9(&7UVB;+a8a_^HI4:d6SA9\JA.^[BACF5L;DIB?<Af.8)bL)LO^f]-J(g
7[0/_/2WdWYfE;<85JRgPV+AZ.9&>V3:/:J>.^)Dg?K]?f9NbTf[)]TND@FVR.-C
?8,?fO/?17\?46W]VN^CM@50\L\6IT5-K..[?_=S>-,C\E><Na7;HT(M4EYJ5P@)
W;)2MXT_B<R6/R9S#b<B\FEBWgGTH[AJg@;R=ZMFV11P5JL;EF5+B6DP@M?bXg>,
D2O21)XXUA>;1D;d6D?LBCY=DQ:BK0?\KLROUX;&S5_Z??#BfPXO=DHeVE[_.+8G
,<KOb(?)(J6&H29UUDb[fgEPb3FM;^R[.O8,EMB[3<9NWeT?fDdgCCMDS6ca0S^6
,B0O2J4aTf)OK1f_OG+5g(9bTYDMdJN06:H+a=XLb(EG7T5+BeU3XD39L+We8QDG
(<;D#?Y8>E),8dR,GTT,d,:a;E+#X3WEZYPWY_&Y4D6X,c0#Ie6P,RF@._QOIP^#
A&0XD6+8R-H?\,6U\g;#aH--.4aZdc/TPN\LedJ-DPB&?&)_:fC(JS[AaQOA=?1X
aQ=\W8Y^)7_VSX&W=)g<^TVVCNM1W\)&b(_@N[d0ZS]g[E_BI2)77C,(UK)g.b^2
2TJD0VB?=44+gTO?ULdE)>\cSXF.YO6MF+VaVHTK;T_A>\.NZK,5.&6H#AC&CV&G
V?S?:]UV(ACad[_#?-\&@IOC9P6-g.S<<-Ab-&?G>Z7FJR5\-LVE:HQ2P<N6,)P-
eH&WL)XE(KGB^0c-8@6-=E82W;HGY,QbaN<\fNYDYZQOdC1@OB+7LU0UH\(?OC1<
;VeSdTM=0K1=J-_(g5,4GE&/D54eM(OH4[P-eg^6^#32_c;GJ#6DC5;IAXc:TS@6
JE4DL)Wf)&e:O2f[^AV\=->I\JS?PB75EX6ZT@R3TG;JHUaNI<+)gcMZ]eMUfSL0
9V()+N3cGGc9[2c@C:a1+ZPQRGCYO1UE9/XaV:KCJe3WOV?<TW,QFZaT[_ES8JVY
\g7CF8VMLFG+(e80/U?f,V]CEC\G)QgfE7=?\(;/+^ITc.05[1@;9c49EJBe2C5f
ZL/I\BRWX5ee3,6[9WO?Q;&>5F8fF9SVaN][<fg=JBe#8))E6V;Zc1EG2?SF#?a&
a^WFF.;PX-8GE2RNFPPJ<Fb(5\#;bN8IeU\FYgVa(J5EMON,U_A8[Td?(\dSI_Te
b0U0).KTA@dOP[Z+S[@-Eb9F,aLE,O6M:/P0-C)CLe5fecbN3]973YRM<#d6Q7gL
c_gV+9V?-^1;UP=N32==>Og4=^==bU;1T4HKS+&OI)L_0LZ_GV9DRd#EUW3KL@La
/_K]JDD^Pc2@,882Jd1<O/19E4)^>@2<bJIP.S=OdFN+HGP@W0K6#&Q][^,KA=HS
0X9O>P-]?6(E4<YgMJAS\/SB,R]W<XIBQMfbG3ERZ>0GHS#43>W,]E42N]X&4I8d
A\X/eOK;_HNDg1R&C>JQ0SBfKd+,3AP63KT-YLK4??5PA@7(5SFNRAKd6GU^=D+P
\-AeN_UFcO/_Z5(K#A5;K>B^:FXBK+#BER?96YTeD&bXH)_:&_8U_0>NX1Fe3-N>
:(e&HdNPbYKJLG:1A](N>H1--;5,E0A._L_TKdU5Ved<C;Ae?,:P+]U\F=De.Hec
8TL:HEJN@V3KSc:W&V:<56&VQ+.#/4]TC>d:DVY>Y0IAXLWW+V>Z3-P\Yg2PL.OW
:cUGS[G+Y@/)2K+AA_O/K&[1F)06/^_C.cHIg(((aG:0\UeWIN8LOGV^Re[0)b#g
DKc?FZJ@XR.S_f06#T<_6YTdgb)XX4^_=ZQe#3QdE+b[31b.Cc)8)WJ9A-U261=;
BFe5afVdK>=0VMZF3Y9\9]U2b&]2X6.EJ=[MHH([8C]S[55]Z.O\IJC0]W)U8P.-
7FD>4[XR6=K?K.f_7/T&:aK+)PT7EWQ&-G8]Q24.b68_=]V7<e&EDceAVA4O6\e7
44c#c+=VLY^Ve1NfW)=J60<G<UC5XJ0,[d572J]gE)II\TOIYU1:d_&-:e2g,0;5
,?AgXJG7]@B27#&YU<W.HWeIXL@+J+D=X1:\g\VNEdFQN>(NW_g1_,-#5U,IWgWD
NR--K(N.[4(H(@C.3D1PQ:@L-5e>Q98VX454LB1OHK#5P/+GE,:NT.AD65N3&?;?
b7PCR_@UL(W=bZR5K@(K#XIa0TW/X=41/8PI(X(J9ATLVgJH;GABLD8R;=U_X:XW
F>dU:D6+Q>/XIW&PH7.<W__Sca<;NRM\a9#=?2@CK#dU)8g,F2?f&[0aLM1H;891
ZC5=eFY:@M+2Ae)-69@eM?0D]793I=89:.0C=O]b)>B_?fT71JdX:LJ-A34HHY81
JE</aT1ZOM#3527QZ5&J5&g,@].JN95a6>2OBH87g?SdN5^_30HC^Oc-+DW]BCb<
ZJ6WOQ7-0-(DLe(f+S<3B^YQWZ.[0;CO0eKSfDf4@\C)6d[?@IR=Q;/BUX_DG07+
YW6Ff6Z.?e^,WS,S6CQ#)X#+DcU)B\@P4[5UO\J<,1_c<b,D;1R:-Q=gcE,K3G0.
?LX14C34GR@LObC/Z:FZa7+#&E_c5?H]79\M&Y>S&@.;e(bgNd_;PSdBN87Cdd1?
.[T:&J]P[\0Y((,2+,bSgXdL@,GeP[<D/C93R/0I9/edc1:RbG\L9e7.5Sf56g:-
FQJ58D#CZIVVg>[FE25;/QU&1LN(JL6e/M@D0fUY&]#Bf=:SbB)(3W/TAcZ5f^8<
E2IURL=Tb;8#?GPe?.Y[UJ&f1UO7G+JG8bV/04S3#]0HIP))V9YY\<S\Rge.T=cD
_7(Ac2462DG-53GMb1H-;fJNC_\AOEZ4,)#1baBMVKHF&OJL>TXJ_S(R<bOe]gFZ
R]DR+?2>:III9AR7eJ^,<J1AdDXcMCH(3XU.CfEGFXU)A\)T>HXJIG+5S:gVOfIP
/9Rd#)b;?fX2HFUQR6b.R-_eL]7Q9R_BS];5aPeQ6C-Z?C=8O@0dUR;([NJXT5[.
:Z,Ba1cW?X.Hf^DC4J1[-D:S/2B0.G<.d6#EVgO+=P6KFDdD4E:00[W.^/+SB<N/
/RH<e\1M(d&b8/,2.BOe1C-.,<(WQV4K#TGI3K_RfDH=Y1,ObdJ>06cD82bXX)2E
eAdJR1092[HMdEQ(c^F]Q^CWW@S&F8#c#c3(_cE2Qc9;IGD0U(N?/H&N;X.-(gIY
JaNe+c]N)1P&#-KS-.<)[QA:J)GdUZ@a(WZAZ)T:#HE3cWFH<ZOK1E#;=PVKOKLI
c-^LH(ZVe@]=gG=_(+:5CYNNM8C/8?ULP--68_5:8983-3c.J&NcBZYbJ7MJ^HP[
E(>R>>(-=A@0LF:B]#@W\fF?9)3MF@H_FC)69Ve><gVd(KYOP+I.Hc&[U7f9Z&P<
e(AX-XI.f^]b]\;XSBLFQ1@:[)_R;#R[J.XTcWe,FbNS&FI57C3B)b=UP/OTAL]2
Ifb_WW9>>WBF>OT.&:6ZBd86+cW-_/9G2dg]eSHW9.\V]^+#WZ)04/NQ^B0YZSMa
e>I^1A[ERA6+BIVS4GN9g+e0:T,Qc\5fIXc?0(aU9[IDUY8;L=4E-R;HJ7BGER)-
3A<1\;ED+W9F=FFP4aP(S[UGFd)2X?.Z[IMUYM:XMJXU;?7[B19QXd83XAXZNI1O
?,(C31NS#>FF]eN#@1OT-c,=TBQ/FXK>)KZ0SJg:\7;=DTJf[0YS(KC-9<V^;47#
^B3Oc^UaOR6e=E_EGOE+K4B2DB;f/.I:)?E_cBC/Dg6HC/e@Y_JG>^BdL2NZefae
5ZeM&F6[gL;)YQ5FFFK:dU1:B\d+]<J13-XeEN4ZPY=QgP/HFQ(cCA[-f/NRR#@^
F/R(TV.eU97E>.X6][88gL\M<0.L<fFed?H>(8;];J4<^Rc6O[ZT,>JdSM=f533P
,17G\)_=R7:I?]]df:cZaC2NP(:E>C[8cP(-)#[84&cI3+\#\;NIZY/0<fHC)LDT
.-#)cGC>63)1?OJ61&Ie@9fY35D;#SVdWZ7/]AQ\EES7G\4#\LVXVU)ff1A[Yg:d
<7N1331TW@P7SO0UeO(_0)T&<f6D^BSYeVZ]+KT;#?-=+:A;]87U<JD2FP<>TZCE
RUDQWB9IK86)9TC9P6VOQC=\J_:f=fJW8#cA;N0HC3Da2KOXI>52@Vd#(IER?733
>W_<ITP5@9^;7RDMU5b+U8Cf1^N)Y3>BIUN(a_?g[CbG=0_V33X99-WODV8?L_[R
-aHNR8=?Z&[?L/@+GX.<LTV_QM6CPU/4[3C5LOA6?_<MX_Lc3_#28GO1Q?[JA0(;
9D6=:.UOFa5R(aPU0e=^[g[VZbB\31=[TCa3Y\Z5(W8e10WS#-=f\2Zg#c=F&^2#
A7Eb#TO=+G&;R@HP3a()P>DbASf\7#D5Ee_-E_Ld><D0ga870T?Kf73eQN)<)T?U
<P<3d=Z/0SFYDGH[ZMfC1+SJXP6Hc.&;PSN36:f<Vbe/G?Q=T0@91E2a4(UcQ5a&
IX:XBVPO(;de7)a2KJfRIK.\V:E:2++G_1NL1_>.1UPR943?/7\1MIHL/U:3<-<:
0V)W)LEC]&K;F;L.L5#Y-W&/2CJ854:X.WLgeFb1K.@\[^K/4FYU2[Tb^BU^Q(Q[
7_Z>D;)T;W0I>ZgI_>aK#bDO00O:.=4Q+2KL2[ZGAUK>+c+eN]HJRBQKYR+HM-<3
/c\<4IT\H]/=abZOLCa\RC3VQK]O0Z4&16[gYIZQ3&E@?)6)KZ=/L6+78<E&Ye33
gf_O[PJ#La/#Id_-ED(0X6e/J)O.ef[F^Ra\#3L4e/\XMY1)P>5;4fZZL7Ue3?/4
c4\F7E-:B[,^Ka4],,)Z;1@)d/ALO)KC+ZI0g7:W[3/BBV8G>EF_dIJNH.3GH0E3
WSMAC:[MQ0-,X+91D8ABLIa:I]4AERNT?9W+c/24W1H<:df8S]cMG\.)M12IN[D>
@L-^a:CFWOb#(g?3V^+B@Q1HN,]O]+d,gFg_+)d+,?N=>@)f_NWe[C+J&bEG1S1O
,C-]^Ob7aJ-cfMe,;OgK;#RY^X)^A31(0d<[?/[N>4UQgY8\7[P.ZEASPb;g^Q2\
TJd#W^#b]?PD[TNQ^fGAZ1.BJAffYfe0_)JcOg,-[2A+J1aO:9d8ecLURgE+>SQL
OObG-QNWf9&C9DX1-66]UfS9/U)N;;10T4T40QHLB:b49<g&(/+I)<,7b79IC=3S
[aJ4JLN7U&6.?0;R)IEII:O\A&U5XXf@4S=A[^c@H)C#=9I+=KWeZ=[0a<X@#.E1
Z)fA#N]>b1JE>T9a11eBedN5?C)A-ZMPX1=AaE=/G1X3GI(;dNZ2,&e2^;ML?_dK
d;5)A;W(TH47P104//Fc/2^<.LgR]+ZQdHAFINES>>_@@@6>[]W+3B>MVNB1eddS
Qa[e?6.+JJ9^aYgE8Jg.b:DK+55RXDF/QBOEG(b/T/#:0=G0EdEdRBE7_/R:cYSW
Fd(NO>,MHF3.N&I5RN-DdD@A[;J#D>.=&:>X1SP#0R#5H^J_bGe7BY:7U[&fALN8
-AVKLg(SdZgRR?233IW-DDC/WMU,5=bY>g3CA2/?I[HPK)g+T(J;fA,P>d(85C-D
W:e->dA;(QF&DXW@YAC4U=Yb@6M#:2J3:QPME),]\Z.&8)G/((&W?6e5WG1T]\9X
&.OS2[>b&-ca46[>J<V1CL#-O?Dcf9I71CI4L7-^^K9H3=Qg[5T<#<+6HgF/BIMP
(5GB>^cgHQS<fQH,g[gg5SEQEP@SP(G=+0>L(NVT^H?Xd5?[=J0G()_YJ>0Tb]2S
fgN3dWKc)&@-YI:fVN,e\LbD>8Y@3)]BV1T(A/L0QI>ITQBX]U-BVEAc7VQLZZWN
33PDAOE5?#SD9d0-&YMG)O/^18WM[0IC-IZ5B&<3OPX06(NJ2J?FbTEM@#)ZWG]<
:GEc\E+g#\?\_ZM?g3Sbb5LB68(\2F#<K-@6-&^GVa6E<PX/)+5\F:T<a,(_1bJ]
9?V&A0)VOD8DKNUe&UA<Nc3Sd3O([G\7[]L]gAXU43+gYF=:L)@8f=e(])a-#+C(
S-BHd,6J,4]e7XW?H;NQc&4;RLPIP-H(JeDPZT1aEV.(K04>,N]&W[2g3RKSGHH>
..#TZXU\8QgY?_R,a@&Z6BD0H7be)B/DH2>WAb(HO?JQ6P_\c6J4K1--L&6WO=,0
S9Ud#YLK3a_7O^a_6\b=I+2BVLB^LFH+3W#MG;AMf-LRUZ2K_LVFg2>0Ob6XZY3C
13gK+_IVY<,/((ITNb=]J(BdKfVdc=2#c>@aDINSZ5YD&@A<RWC24:6DObc@&W4>
@OR/.PYf@H[dgDf--e+\AED.DL0^c\I.6UQOD4:811=XB7>gV?0U.dC8PUKVa]1<
OLS4:((R<7D0)#eS=9.1E)[Tbc1+;G20bJTLS.Z9DX_FafQEB+N]TBfX7V=]I_M?
L&:]S:X>GSU9XQ+HMUdM+5,8UP&[NH^.;DaS4\L].QfY_CQP@#AEU[aF\IB-0Y#J
Yff0T#E4A-Q>=aC7L+.@Cc9f/.)e1W_<f.CH.DNH:HMdT#Wd4Wd5gcKVDcP[aLNJ
ZSV[P:E-@=fUI@F00SU2)AP9KGOc)H+BO1B15Fd6O6=C-/eIG1F\JM5[>;Ig-M_8
#ZZ[/+?(+<TB,W>R\4,f,c1BO0D_0dZDLE-FX)HZ4/04G5;G(++>I9If6RIYFO6F
UQ<_=[a\]b;Gb\F:B/5d#1e4cYF-9C[W?&W0_USL:A>52J,.KPdUCIQfF/(TB+A;
UJ)-):;\b3BFLa;eGa7Ig,bI#c-=;L\cY_ISKC)70W0QHW,(<X304#AR.gCV/?R@
\c?6:;U=3)-1V26=0Y[;AFSQ0]0/>6V_>0Z9&:2^M111:0[=G8D:Cd.GH7SDO5^e
G?BgA_8OTKTe54AE6\S<P0_N@BdR8R?TgY)H<U^R-V<M=Q=@B8D/[\[.XTW+V+Hd
Q3O1(Ff3QG_HR0+b(N[KU8aF)f1K73C17;PS\f:>RQf5B6aCb(]cWJGO8J,(HZ8W
M]8.<K8.GgM9E_VABXg)[DCG@AASg<VL9TMb1\9YYU3T\^N@VFad\X(a8dbd,LcH
bS9e0fF5eBCbN>RcP0AY]EEXR88/1E8YHJb:)H-<-G[XGIc@5?2&BJ>.QY3SZ\Kf
aAb=JH243U]O=_;0<4R\aQ0;CP]L\].WfTL@0e^\IW,E>B^[>95^O9;2\G@e,K]0
)D@Ag5?IMaIS#7aKZQMQZQKg>RA@0_:9CDAbUSaYOfY5(AIf<JM1:;@U;;(a+#F-
^5ffYE-9LID6MeM#\QN<NGL->WB2\?&b[C?LNVJBWVBXMW3D.F+MQCdfcbIe[B&O
I_FHfJQCg=O,[Y<Aa9XS77\WK/-_OK^LKPP0RDU:]\Pb\d_94MX^^.NAfI,9KF7E
a7P0\G3-U?T]Y1S6^R9CG69>#D;2FfdMV,Q;^eUEE)P].7I>.K6P9KLDDeRKB)W2
.O#HU6B4R^&\MY/_:TgQ7F7H4\<VgO]_KO0VGJH=b-f4I((MYEJ)HdeV@eBG_#+g
=0^R4OH?Fc8J6gG)AG@C1V(b?2fddU<,QeW=Q7;_JLQWaR\=+SeR#(a8&4_#M#8#
BDdB(B42WNVd)Sc\E_M(8HIE6FXK(KQ86]^JEZ;aCdQg)b^YE2_2/[=<5OaMS3]4
JRX-5/]RGY[M2:E1fL->E-#7L]27=+E\FHVJ&cB9-F>&G8.eM//-e+KY^LXFPXZ,
/f&6?<^07a<6S5O&]>5<V6SSJEW?eT)<.f(1RWU-;VF1@c@_DTd0Z9:M:Yf>,I&G
:.A#P^[O=^cI)dXTe7&Pb5M(gPRCfURFHdNIYV>D7aEa]Cab+9/>/]YR-+UW2KEK
BbYf_6De#/^3HI..MXX;5\>P6>Q1LSfBT[GD_a?]-QMI0^]bgM^QBePF:TLQOSU@
Z8@/(Nd:2M[)(9IGCY^;98H0PeAe?K83(fb2SVe#IHdOG4(8+M,N9KE&QBF0fA#I
LPO_W-^^@83P]fc3==FMa7<_R]B#BQT+b.a_gH<N[TMS<8@f+Fd=X3.=>f@@7S-K
TXE,_L#[GN1(c&:,#_ZSg8gV1WW-_4++J(5&,CaK0Q.3L2g4O.Q^8,.\TU34R37@
.MCLb8BLXF&aZdfaR&UeA/HKVO,1g&Cb@d]QK^f<gQA=DgG;TYNOa;0eFA+3J_6#
(T2B/PB_R0+.W_F&CDbB&PFE.ZK([\^)V+?CPCeEZ?8>@7PZ;3DQaK#]4(D>20#2
d>Ede0+_/e,KOU+aEeNdJ1],A?3ZVC2@N^/YSY//Yb2+.=9#II2W./Qa&cgBO),C
;=1f82#Sb.<(&IWb2Z5Q6UafYJ,YSJQ,FROeEdAL^CL#7,g@>#HL0eF1DB&,UOM2
M3f/N,7U\E>WF4_J>QQ^-De^,,./EJc@+1JQLM0V6[R7a^_QT.:D:8\6c,=Xd+-g
dO852?JNA)B2-2b+120OINDF-B,K46/S_:b=TT4T^AL0b([B1fAIB\/9;-QLO\(W
.IN2&23TdfBN5J\2)Q5>KUebc.S7B..+?]C4=W]F@I-.)8OXM=eUW+6-=+;PD=KK
J:e\K[&g]50/;O<\&U@G62/ZZ_C1H2g3.)-M4LU?:0,TV&Id80&/XCQFT7eGeCIR
@X8+5Ua#?QOI9M85DM:&</BH/:_Q+Ygb,gT(3-MM12,9\5VWce?0.8-bSOfR<S3e
WW3bWc,@-4U+^e&93__E5?bM]-]BZeNNF-aVNO)N6K#H9dcTZ;feS^[1E)75J?VR
eZ=&39R]ZK(CJIJ:N6T6abObKFb0ZF85gR+])0aRR9E:&:gCL]3cd(]47\gf<I.T
XY=]f>_V^8^Y58FM.KIT-G@&MbA=N91+:aSR-AJ\U&70U^91GPMSJRSA4VEE[g4?
:UW31d)N?WdJ0;9DUCQZf2XE#:RgE1Q2d^d57^_P^1G(HcTIE<HWU.&-Uc8H_g_I
4)00A1c63S^];56LE9:#7ILd;CS9PX-6(BEO-ZC^9XIYVCdLc]\/WIRL&S+1#1K5
]d:<]C)\6f)(a^UUT9/dQMGI6AT2@X0gPA70^J:=UgKO,edS@>FG<AXZ0CLfc&gP
5))Eca8?2e=W)8Uf3Ea9KK+Qc@aKN\Cf&R5fU;Jag@5:Q.A96/<K)gG12O160L8W
=L]&YF/0BC^2_YTI>:a)@LQ)Q]?-A5e1^27P]:V:c4ZGfT?>f1a:a5)1?1?Z^Y<G
_=cf>PbBZAE[Yg;I:FR.86ZNFHccD8GA+?]b)+;Q\/@6XW/e4RH;R#-XK2:\1+.A
-TP(LE?)b&YE5#15/Cff<K8#U@FH.-[[JUU2K]8Tc)W#>P==?)D1_E.f[JF;(Ua8
,;>Y[RSILg/)b3EBG18c9JZ/#f><0HJ5Gf22R/23TZM.:+d_6e_]J6A;^I1^.E84
<KgG3I\+&9IHPPNb1[QC,gX;c(73#IbM&.3\IFW)^#c97<NfJUKQ_^N^4e3::K.C
;0JM#GJZ.R,g\9Q&&]+gg?3^R2?7Xeg?F5>J;M\2a9)7CUPR^=ISYO;ZMb&PU#KD
.MbacTU#\I/[V&XQ9G^Nc&c1_>,LA=KPJ3N(fO#XPg6b6R6_>OXa4E>RV2;Aa(;J
GV2Le5NI]O75f,[UXWc\&2X=MX4FG_3X?IQ#1=NR9)I#P2S7aW6-TTCG1_2T4>KR
eICXVDff5KU=GLPa(1;P6);_30DJ[L[#4OBKS5Fb=>ASENQ2S?&ac/b?=2c^<&.X
[HO]V^Y5?d);@gg\N_+@R2>IK3fe?]aA1YPJW)a=:]PK7Y1&/eMI53K0B(4,Y3G5
7++A0=4aM#>BT>DN.\TGTR#9>Z?7GbbAYJZDKeM,V)X16VQ@X7UI0I@[/[eOC<bJ
41fRd=/QeZ4;UIUI#NPWOG)2L\[GS?MK\,N&CYC2)XBb]TC9>QO7N#HSA5M-b;3-
T5J<44?B(J+L:@;^3S521TcL]bc@;98eF,_5AJ^R&HQWV^(MVSN4\24a0\YeX\D>
C7b481LTO><GJAP4?d9\S@aWMJKY,B,6TV52aYQPU@,cUDAH2W=8g&6(ZYYA93F5
LWHRdB+B64UTZFO:YA4#=]Fc+f?,5d^.bF7,;Q[>?@+\W<]/B7Y&:5./P=JI/+dd
5)5E^.bIY>b/fI@#/&b5W,<GYa8]WM@a@G?cELAO=1>W(XYLfNG&Ice\R6[]<;GL
WR81gRMECY<@E7E)de4@:N>,=,]65Pgg:88,Fd^Lg[eV[>:/Y)9:GB+J?;-)1RUM
((Ke[.8Uc&885?=#4\KV0f/APE]O/+7K-,(^Va]eMd&V4)=Ab4AUf5XS/^77/G:G
K7U>_3Y]0FH)JYGbAR(ZP_V9SBLdda.Gc963==PS^1/)VY<9:U/S4:N13O9I3,\(
,]C/I]V9d+N&^VA(#PPC=MY>S.;0YgO0B2C2K_VC8D.=NX\?IgC<89g#VIP+?b\X
PD^H;Ua-[8LB/G\2#gDOeYa&eM=KX>+-eKb&8?/ZG^149<S>N+fTOMV(G>9BEg\7
#<(JCXZ7-V4FH^]:A+-#&I_-#e3=TJL1AGbfOdPSLM7<)I>SEN20RV3M9DUPZ/OS
-e-E>Q+);RJM=1@11G]68?J^:TZ2BG@I@f1LYfN4=/fYgg=F/+CGMXM-Qb[d@g3;
VPC;6)[O3dOaNdP;e_7I4#Ha+74ITE486G]SC_+#Df,bfA4+aH4deG?<4KH0O8,2
ZffaU];,G@[cZ]IYR?__(3CV=0O+RRZR]LU6E0]V1;dW2eX;CNLNNNVC^-H-TbH=
>d,a=g8Ve_KZ3[Q4Z5D-BISaNF7YY779QFI=JUScTPQT=^>]GM[+\^A&K5cX-ERP
\J+R[L;?F54Q7H&RU(5A19G/g4C5C]/?-T=+ATNTN#9fJ7@@A95/J55cR+9>a72g
MQBNE:bIG6Z?c<e^U#;W@CVB#)2ZRK-M23--WT/>c?[31@A/03KgG?H9D32D9dYL
cJ2Rf:NAUT4/B-)&U[8B>b\ETf+-XXXd@fB2:#/]03K1WP)Q80/cUeD@b7eS[:d_
OMFLIV@B;T3E_;C@VF4BEe?@4N&68=K0?=.:;6HHWJSYcRT47gJ])>b4-F/Hb58L
#;PB1U1]44MO5M^82S,>7;.)ZB]7L4472/C_^M1E2/MV74&X+eZV69JDb7TWC7e7
:._Q/GU3\TdT5a0KZA]8I&7.L?1B)gT)?[fSSN=_e<]/W<5T0C,TG^OJZf:L:6)c
1HV,WION\<LY/MO@O819f94c]6[\0H#/U_E1Q&4,aX_^=VG]P;G/RHV>10d<N3.6
_acP)GS?<^R^:^(D#F1d25Bed;-R#A?#7a3IFDHP&2N\_[+>O^PfD.6a6#,4Z(<H
#;8_b#OSGb#5X;(:6ZD[N+TG.C)QC0679(Z_]YS-cB>+.36\Da[\H<MS^5UbR0(N
TTEaSMAeT\NLc4/IGVb0/;,ea5<ZX?=^]=SL\]1a6KAFNMS45>DTCN^b4VG./Ke;
1/b7F?<S6BZK[5gO@MSZ4/+#\e0/8&\d)Fb#S02DJ])VU48d0J;-CBZ(?VE]a7F/
2bc&Z,_<(F.K<HTM,I<O/Y36#VR6DKA\].K#JfQUZeg<>O[\D]3PEE?gc]/c-d:b
C0H1N3;]g_fF2C@W@V@2T6-gW\\bZ@<4I_fZWG4FU)?B[DVMZ/XGQEBGHZ)R\b]N
<f_cGOf>ELC/ReRW5/#:]-+@MKK(VH+=;]=9;,0J6\T:<.DPJVcZZ).U\KZ#3XJ(
OG5D8VJM8EUAVe]BFfP_=Yd7#KST42Od0Z>:U&D&eZ0VUcb[[F#dVFI@03f3ZL<9
MbPJ>4Z:I=Qb[#R8BMIGNP.c\6I=5Ag_<R@2?f,CNN,:\((Z3I79W4LA/[f<)+E(
^DTeLCX&[f-Ie@\KEGMR6^6MXa+ZX#=gI@gN>d,\@\0Hb#,+BWWOK]J\=&>U4Y2J
eFU7eNI;7U_E[gXP0JEE,A@^eR<FBL@<3:N4^<)4,^Me(FWFX^DDX>QU<(_F>0/A
S3\39^7&dWU;2(NG->:[-U4I:ELX1[E\\]\<SR93W?G7cC6bGW6T2Y=_AXK^A3_L
)OfR-MQ(Z8[2d]Se5\D/ZOb>&Q8UK5?3+;)W7Oe.\V6CeO3--4]G9H;?T&)@KJHL
K00H+8JTO>.>HDMC49K/aB17VJT(9:SR[G]DX7aU[L^QMCe.QHC/G1SRF#1O\9EZ
X&EJGLW5M@R/4a^d<-[./C9b:e#6@3Y2^GU6C#I[6dPX)KfU-70OQ74(F_JM3IGH
3\YQ_5)bgdX)F=57N)AbU>A1]8U(/3T\6(PT5XbT=W;ZB_661^R9ddUcXTDFa[6+
Q\XD7L5f2G]]=5,J9>fJcfXC3]^cgYSP;DWVf-N&ebX(@3d<HZ17VP;A@S#W/[O&
8O/YB\DQcU^_B3B::Ig3<>R?;A@?&M7&Zb,@M=Rd/:X-LfZ0\^f.]>B:N..VQ<f/
K+\6--Z-/b,?>\4d9GP.E<[RedeI0EN@<ad<=:R(f6Y2E]Q)AP6/+ZD)\3HJXH-@
.MW7GK0E6#F>3T@9)C,4MLV-;+b,(+4)YHc=S9-RQf6:L8-[:+M]fR@L;7#CfB2c
M_OS,&ZZ6N;S+.5B[5b<X?0X&_W#Ub\_Z4/Q^4d^+M-\XV[a=^,X;Q1U^[O5#aL7
TP30=UG+5J/GT=C.-R9GQVNA[#HU+;&U-R_[JTa87A8MaFEV8\/>GLYFYQg?7?K&
9,D5db;cE-6gaDZ:0.A@7=K6?=eXg,Q;_/?PJFPOWL)P8VFZ0VB5,gS#1GS#55a)
9(F6HD2S9=Ua]Ec@7U]9aS80-N;]d>.C#F\4E5J]]5G:K[O4XWgDaYEW)a/bJS#W
U)-+bO8\HO/bC2EccEP#@,a)TZU2ZK@,T9J00L<V1E&8^8NVgDIMN?=.)-K3KJbC
Z\]K^fR(;XUF5BKb>[LdRA2;;@_PHI<[I#8)ac-PEMI>8ZRFB3_?)+:K:>+I0HdP
OZfa^MIP>\+?@.eOL45W1<M^T^&2Y)I0IaC<,\]G\g8#_OK.0Y69V@0TYT)9c7/b
@:>B=RbfKTMf?8Y:M2baS:bIOdMIYceDEg1YFZN@)]L9.&&)4PAMAe.=K=BR3VO(
]C\DB#)R<Gf2S^;HC)E_c_MC8>Z)IIL:3Ha(W+f:/Q9F:ZbN0aD18Kf2AdIFJ?T=
4(8^c0.)L9\d1871B4VF2:SQ1)[g?4_0LM0Y0Z=PIWT8WL<7YZ_g^Y\UR^c_8-9Z
\TN@5,29+W,_IK\GRWb)#:+;F2X]ZH5g3IB&K]6D]HOD)>QR9HMb<)M8&ZH@#^H<
HE,RO4?]>H@(_dMM&CbUb.==<+3(fL_R:e,QI/9=E0&<)^F@+8?a=NP]1;=6.7F6
^LV32#?(L(VP-_K0Z#;\)64^^CgHC?eKMEW#_+XEA[=J;AI;+)?[^8041O#NYZ3d
+4[PSC3<#TPe:8H?PMG02)405Y[1CZ=A#0A8D2\:A]:f9:BF<B\7SC>B^geW7TA(
;C0_[J^ULa8@B^X@3G>QA9HJ[9#3,f9ba,QK+H?df;^[:]5=1U4FfZ4N2b7=(UEe
bU-AA3\3Ag1T?F>SY+F\B)UYOIWHG5IOM-0,J0:[PER=bV-2F_@1bc3&e_QCSKV7
FfF;5X1#].1;Dd_(gLMT4R_BMIDBB>/IUS+6/S[@CG=SM)baJV3K?H2//;I\8RT0
8#dO:OS:(<6U[S]SA:WNK04e<eH/c7Bb6BYL\\L;6^ZU0X]ZLR>&_Ke-1H.[318&
5g<EFE;7,:48&1(-,CPe[LB[(9)ZLDM38;8K[I:G0Reb;+\-;ZI6b:K);[&\33Y\
H6=1<b38Z]:f[N2QA3K3R/aX.2X)H.XJNb2&UNF+W(?B#ffQ,O>IDQZG[B7e/5cM
QVHXL7=FE5G0O&T.&5DR/a3);>V(<\W5OgQ+5:+^8T=_cKgNNd=aQ-R4\&J=-fYF
?g3IQ-aN(+8a0WOZ5HHH,+feL7C1N,S<YaD9Q1=G2LJZE2G;KP;bFP)[O2YTL--d
-9Q8#cb^^?_7WXV>2=6E\,,^)KLPfa9F5(e5/ZX0Y&Ld3e.a)#L,LH6A+9PG&Z41
+LK3CdI15f@\Y[C2CH^af0V4T#2JK8S2F&^FKZ61/R&;1<PJBaK<2(:=[VV,@FaE
NYXDAcGE.\W/ZgN&UDdVGR9(4@c<+A9KRL?8/6RL>W5_Z\Zf<EZUbE[->O5GRb/K
d3+T=)aNTB[H/f_\]U59>^+]QTb1-O;Rf?IU=F-6=/Y<3cCcP8GRTXF+.;Q6U;Tc
c7?<-=GQ>YND7O9H;ePB,\_<Z2>+66<=Q;B.B[5:7VXb2+PZVVdF9c1a7E/Z17,e
YACZFQ:?&3Wc,V-Ld:UI#VGIR5ME@I>LR,Y#YJA/)a]Xg<L,bW6&Xcd-C[dZ;?O#
CFL+3T<K.NfaY:&Jd#&7>1<1LG9E@fGDD-1QP8XV9B&W<\c_#F8FCS+P9>_L=NT:
1O&<A_,(^MIOGFHF.1ge&&)T?VPE?;?)[Xg@J1ZEC[L)Agb_0?Q50Q-OQA:XQF7E
F;-(GFKWIL1N^@H-TIKJg+DO:N^,T&VA)P.STUQ8-6GXTZWJ5+K?-:P+M9&NME7;
SE=UJM5X^>78JZW[KPc9(0U\#^VL7fCbV_J3bQGZb)@a(g\6\1BP79)&XB1&J.3]
_<TRDd__M5=f5Re@YX>-;)MT7;JLRJKJ,B)/G[Z\9Q\+[F(5Z,X;+C/?1JeWC)3O
V#]N97VJLB-Aa2SBaHJ(]]FN_R;Mf)E/IAXbU9:B;/NSZF2QLO(bY)BOe[)RWd8S
=1?O(fOeWBTIe2<7J?@?4;.TDR@O<JMNM2HGHd\@S8a&e>#1V-CcR7+UdGbJe:(E
-W#)</]ITL7YN^M>S6--R?YcGc7]cPI>&#2fgUbAIY&:f?U_g93\J4,+KI=<U-&X
a1NdC3^1QWa[bM?-.)@NJ.)_,NB:Z>D=QRdbCN@)\:6K\(\Le\Yd<CNe,H-(#29:
74b=.[M#HPfgd#[a<BR+1<I(B:G6U1MA#XPA1RZE4g<IFKJ+NBg>W#30++041_@c
9c:7@A3HDc@D,Ue@5\PgL;CO(5LTUY.WGGa-AEL9a2/aHQA9#M]2LVXRL_A>\QBM
f@a?W-AYKO#T.MQL\;WA2gLVIE&3e1F3H?U@NQAZf3#TAWLJ)S2=_D]8TQT&V:[(
EPO+ed0Y5H5I@[G:()TTD2G-I=d7]4G(_VFZf^g.-M_Oc_XQ22ZdZ\f?]Xg?-\B?
@X_ZgWPX-?OTb)9eLD(<UV[VY?c,SUMD[@-+_+6Y;O6\X2A;LCg&F6cTNGX0#\/Q
VL(/JF@-8BSZUXD_-b]LeY.5QSCFd0E?/MC>T<ES)M@/U=22g1,HI5W&1ES+^9J0
4ebAd0/TUc<GE]<O5CB#YNE(RYPC0SHfI@SI@[2Yf\6]-V-RKM3dIWYB3TKe3EHZ
81bD/geY-bSKdI0ZY3BS\Q\<WLbM8,fW9<:b^eeHA,bYBgA6(L/C2&(B.F6DgRd5
H4Me]5W6EIJV+_N[9Pf[dEP)gJd/F-K>.92]DaJ5f@32@6H-ZI4/[URcW@EW7VG-
8ZLUf^62LJB#RY(AG1T7Fg@:B_M6U;0L4\XB#cC2E&2cFd1+/^UfM:BXR80DE6SY
7J]2_bQOe-JP=d_<DT<Q[ReHF,_\P;SU(e+J#9?DDWD03(R>@fK3#SM>[08a/HD9
UN;=1X<8;)QN/TZD6=Ge36/9;#HX6,d2bGUE=:1>XPJ&6G#14CLdXM1Q+KQ7D#aB
H6BU@]R.14(T0N^b-C\I4@VfOCN:DCQNE&.c).P>/>RMfYT@GV4fNL7A]C<POW-4
:35Cfc\:Fe;5<JK0&f?TL2+D(GMf#Kf\?LIYQ40L7c44-JJ>:cCKb2e+I,gf\_7#
;LB)]@aY0\]LD+TF@.a)O4AUK05;eBISd2)bAV;XL\<f]]JM1[RSBgJ:6Q\(UK94
X1E<;K9NEQQJQ;50A-__cddP)TWTWFMK]AZ)cBIS>@,C/C#U(J8@0LN5VJZg_T:2
5\]/4^52DR->?4BD_bOW@A2PXD]W/HLCD:T,ZIS]a53gO9YTJC]C3(e#[@df[B@d
C+d)cd((UUc2bbfBbY,a6G+D\WH74+&_10>T8W;>Wb0=d>22+A)aHgWHV#TXQ=Fc
dV&JdXG/P/1D-L>,35DbRJc5U25Yb7>c?]Q<e>4#cA;g^7QVF2D^6@F[HSZ\1SVP
(dUWOJWM3GKUD&=LZISI#X>/-@D.6NQeJ(?8JY>RTTH=@^OSQ>@@N27&=VLQ\D6P
26XH+AVZ+@@:U_d3VD>Bc9<ZZ^+)C9a_[7/WZ3L(#GA^5a;2A.X41D;33&2^#MCZ
A9)JSb?fUOBU?a8);<#XG;G?9K-d8^L@DP,,9;.8H\(fL6PV#FK(3Q&Z>H?<UD61
EFON,7W_1#2G.]A6W\>HU.T8W&]2&Kg)US^YBH_HgGfN+@(=2UOL;U#KJ<9Mc;ZN
6<I]7T(@BN=Y-H^S#D/;=NCg]JYD[Hd<Jad6#eD9@\EPDBP)?WD.aJ+9VC=6(1)c
a6&U5IWe0N&YS]b/5?LZY-B_d0b[gLJH=Tf2\B;M&N[/HQ@6;c1(#e<VHeIID)]F
1.5S/IR634H0PM(.d&)Y#b-X/:I?Bd[N#BRJZ<7C+51ARJ?+]=>+U7N_?)4ID<6I
Xe^#^[#6T_6K&1F=YW^0#>DcUKf/e_8HVIa&[cI2G7L,5D(D^6)ZT-N[D6Y+:]H/
#2H9fE=K1JU69Cb\[(cS8./R.Qgb\O6A-_3KC=,Z=UDeC_8MDA4>VE?EUD0,gA0Y
QcTT]fMfg0>=Q_(AE@cEe1K,>GGS4O&_<E[ETfVPS#gH]cEMUS]OH44OLf_4UZS\
P7Z9a3L7(K4M9(YA?;MDX5@gIV1QY-R)6[B_:YUDP2AB0UIOAX4&^/U)&\a6G]=c
-R;VW2f_-+:G1B7a/1KH4-JJD4RIXe4_)XDXXPWTUgD3U7+AS/&8g5b].T0(ZY1@
cWV;d)F3BLY[R@Y7f-YN\M5Ic4a+U>99dDZ=,./_PE2(b&>aYf=VK1P1\B89FGQb
TFI4ZHg(eJ83Ka:H&2g1K8D4,,@&g^ZC4FA3L)KZ8@F+KR6fIa>dAAQ(D[Ge1W6U
IMZ52c&d2JKgS^25TL,LA)\e+^_UB)A3JBW<WbRZeZV.L4Mf.P5_H:K;\MH5e#(M
3+G(,<A:H,bN]Xa9^^d7NK]EKR=YV]c(<#P39S4We:H8Z;J-_0fDGV],KL<#T_R&
&a16TYTOg/];RSO0TXP^;XB?/C4R-3?--\V\K[>8EV/)J&^g;TcdHZaC^cLJ+f[W
:Gc^]0YbBA^aH+gNB(])7BVIF?da@(3><9f\CHZGEe]cc8F>R&_?1DX17W?G.+1T
fDT)QHcBc&-Dg8:cB)YCW_7OIN:FHA\^@,A:/)42U@G0B?Q.4H?+QSg:>e_V<KG+
2EF&Z9WL0E=gG\a=?KJ_)M[EVUIEX^/FFd-(\Q^JU+_cFRH2-B4T,d,I]RZG=+b-
Fc4bA#[GJ>9gXI)\a3]D1#<cI+IN]=cW8cLPPR=EYEaS#<:>N&(M5Pd;XgX6+,:#
B08K]e;:[]OVWH4IBI>gZ7Q?RS]\/538E_FOdPfK2d^MfI90Y+?\#2PZ><aUe?<S
E8/OJ]HJ5:gW+^.N4F<8d2/2SVPJ3UDL>1?aZT^_J>Q;W9\XJ]);QgT(aRKK&CC7
>NaY^JTL@XEZJ<E^aICc@GgR&F8BSML/1cDe\3B]/AO\YD>f;Z54?7Td.PT_5bRE
VRd9CZ88>H2cNAU4/@c[_g7c\DAEC)4.1M/_OMAAFBNd9Y.<:7NIIKd]8Oe_e8L7
bG=PD5&)1VK&c@:QC[Y+A4aYb_Z>F8c+,-b>U4,Eee()I,-0ACYJg-G,A<Y.0J1H
YY8Q?Z,dCNIB0)EFc=^B>K?::04f4W)/IQB@_8,(-A3J+;UHM2M+(dO1,,Xd:OR:
34@gJcc@;R_ObPQ;gB5--I-<V3U275N#YXg9b6K#^=X,-<OADTd3WMN&/ULf)^Gb
.eRJdacMA\XEQY0,I(D/Z9QaG+RZC(1UaQ2gf(]11b31>_THBW1YNfP&KcU0<I2X
90/K?1-]CJMH3>5aMC=4UFUV7^<L2WfYf3QZ_9EJHZ^@X+Q4\Y+V/6[,70.62Fb9
D?N/89<.QR;()_6RM)B\(HROM..W3f:D4?QEU3:3ATSZOH@9PEZ_bFOT=OfLFB\R
/>FPLYfU\gf&aNL\-QAO2#0UA&:0cL/3F=)&XU-8:]<RR7[8;+D#-]M&WfD9(A]g
3f;^S-SX38QBI9R+A&>+2T+#DM7M8K\BJ3dd[UE5QBNSDQ=&<NPN?8<CbE>>AK,5
bbK@0D:(;@5R<Cg8dAc&0.1<MQXWU/[YU(\bg,gM<2UHS@&bHQE@HW?5e+GHg=+]
JO4)J?JOI-ZZ5U.4?PWa6e@V>MLZ:d+1Ke5_SFW0JD/^\d<=ZF)7E^bF77T&IQZg
YX,AbWI0cOfgc6BKgUM3f_d3SZO,9:NSe(M3R)I]//Pe?R1?]5\4a9+gG@=J#9W]
K;e>G-)B8f:)[[5W[6a[ZI^I&>W0_#;W_@QDYOVdI?>2L;@2)8OPZAebHQ8T1d2;
DGYA;e3N@83Z=@a\+fIc/&=[L.:A/@HE9cN7(?8<[]U-2cH2J3<_\VXC1D^32f4&
LXUe,F/#=X\V_3:g:,32f6d9NFLJ3OK0&MLBbLcXCY5PV@\6(WN]PK2WI1S=&9@7
^J,Q0C]]7ECgWP5dDQ90-T98+>I?>#6)V>02NK&Af/ZQY2>)N:O&JOM?FH7OWS<A
ag+P3R9O-,Z:Wa]gU^Efc/@)Y)[Zc/[E^DE.P^faH(8KH_Ld>6ZV>c,eH5H,H2<C
W,Zc5C_>ZBaHC@N_b(WOWVga\ZfPMgIgE\LE6K^M5aHR\J&A01O=d+@^?-d<FH:I
d@U=X15S_K4F>6f+0EX23,61>/gPT\gL[<>SSSV4Z//\b3QB6+gH+dCZ(RdF(b4J
0+)7FaYSZFIg>6V^RBVGe8[\E&7U2\9+3S-E_QU@S]-?+D>H?)V>V.TC&d1CR;P6
d2>+eaC=fNK[B50(GQ7_^]9M(P0B:c)Ndd^_=413V2NcS#32.]WXYKUE[7CMK?N5
Q:(dG4FO]-aa-[G8ND:06B8YId(a;OAIcXUX8R:P+B8ZY2Od,OZ:#[Uc9aTDO5OR
NY55]N#9OC-PfQL:1^f^CdKD15BZCZK]_#T8S41L:ZX5/&]P=7^2/6M78XEV#N6#
A2g;I76F:D9D<MbGT<\NX7W=9(B&::;R(3#e[]I7SAPKQ_ZU4<VS/VY8S1U@JWOP
V&ZJ5X2?AN)ZHg4&W[;.L3C?g-.U3WQI#J;HEGOLa2MTDFDP#V2DWd<9KJ#?)/d1
3:bI[HfJWECJa5?#bA(&R50KcP>BXS9/PWcWEgDS;\?C]R93:8Z7C,V0b7>Y6T3e
PUFUS1?);;-;4RV(,>ZS2P-c#c_))gfb\@d:\YPTT&Ug7?bW.LN&GD6)88:XI4KQ
]8HE.g-+?5O3NQeb.C&2@Fg;?KO#@+aE,/PW7:F?A7^e-&JIE<5:aEWU)JNC1Ca4
VV]<C.EBQOae4EDWG,P:dc[#NAWfFcPP+_DPCH]Q](8Y;eA9f9Oea:H@^:e:H]KG
EH-Y+>+>d//eg]bZ@50(gILY_I6I/+:.T\dD1^bIX7)3,=?0\f6Nb^SBCDAeQO_7
Z0NZH+.YaD?,fND2ZaO@BgfLV>;Lf7K\+NKY/_Sc49/H:60<e.R,S49H6aL4[KN<
f\\MD9JUW2URX-3S6/6TOU&S6<CDV(\VKJdVD@J<NfTPbU@Ug_FOOM]NYXBb7A:P
/7)>?5d^P1:R&R^=8Y/HE>aF1Y,,>H5JbL].Og8YRK[dMf=^5B#UEF03g?2M6BPA
,)a7E<OC@<,.L/D70URa^4?/Tc+\W32I:P9\?E^+XJd@6=6(7bV?<8d,VFMXT\OL
deM,N+68?&CD6&&H1-F0<0EY>>5-SHSE\afPQ^DGMc?[N+UEB)DJg4>-BFU),Z/X
=GM#ARcB6Z>A&GEXdP,Pb/73J:3133e-Wc_ebfOU[/GTgbYF6EH@L_SST5#/f&2N
&f218HYR)P5.0JL[_:a^HfZRL@@-@dNFJGE\(ZPPa.M^\_cYAPXf_M]e83N3,P[@
1<@W:C.JMGH^bYJ;=03/VD@8MaOSOc^7f3XdFZ(R=JONO0Se0&/>++&K1UDRAd)T
27XK.+QfO#<[\LG-P+&f8H83N7:J\7->Ed;^>6;GAE8=9YK3_HM+b]IZP5T?PbQG
M(<aJ]SJIME85;#E?c.^47Z#0PQ@OV5\4G+aZZ_CX7\;(^R>VHT4Z22Ob=[R362_
UN@ZH=S1\P[c?&-<O-3_K5e:e;^WQ?#FU59U5,T8?<E]7Dc-3SA]f,B,=]ZU3J9V
414Z]DP,6A/Y]OQfEJK,O6\OZd)JJ<N-B0M/+.<DG#^6TK^F1>6=Q@POY1R;?:g2
:4EZOeRX8W)NS,Va\D2):/ABe:7XbbeeGEZH[FRM[/d5OH7ZMB&O?K;=(R@Wd9A&
=VM<-ZOR#b)&52.QH?6SF7@<&B>Fc#fG7a+:W)gI?5A(11=NQG:02b7Qe/]3OZVR
4=@[?YQ9/;^e4O:BEOX\IfJbGFcA;d-6>W>&D(BYM7_MP_-&L_OASMZc\2Je^YN@
P=95<]E-:M,/2MZM9-H<?97^RWBSQ3(].[cG\XW2NafU<DYI;?7,@<URbgCQ@L?^
RUOA385:I7WGfA>]K^[Nd0?#M1eG5\WI+.E^ZO;_61RJV/3Oe+Y4V0>Z[.g:ag=B
a)<2A3PLSO+&S2Jgb<IISB<-aMT06\B-\DKN(?-(Q&H+_gd+;e<@80\@5_>IX>34
+=4PeY8?eC#Y:+J:Z\fE/4#\9AYGAF)/NM_R8SXg#NPD=A[F>?0/:>;&7V97_^:4
beaSE,Y,G&PKbf_7_;\,X:MK:=VaXfad/UC?]4-g+^ZO(E.[.)>6/g;U7B-+f,C9
4)Ca[_.T=&]?3X:Ef5S=[c9B4)g+_&.Se20W&U-\L]3-.2?0VQFg?bfTHd_EB/08
]UB+0QMd]S0<<fKQaDJcN\74.TLS2QE&O>7V@3ACg4T&:UJaR,\;e4PI2#Y/65Y5
#-?Vb1d8N^Jg8\W5bX/#.fdWcLGcZ&J@BOI^3H&ZYLGGO>+SfX.17BW^T-a[@3I5
K6&dS?9C:CZ#W^I[YOUULA6=(9c)RJ_C^MAN39aL,CCKE6WI(R]K;0+gUD)..P,#
;+>P.0J>QN&+78JA0^^6IKH]W@XQ]c#S:X8HY7[/24Jb1:P/gUU0LXaUO9J[-/4d
#\^ZB9Kc?8FAKJQI<I=@28V>&SBN6OL>KX]4+/>PY.VA76/)=.E)L@RLO\e0F)ga
e_:O0)]D5cZVF02AL\]?1D8ddPUB<TT-H;5E1O\79NO3[[XI/9V+-/[1.,S((B1&
X#O)>N@>XRE7\/1354C_+H4_[Y6bCSCGa4W?0)TQAKNa4SKR<>?Q34YaI2DAQL2Q
U>FIVc@/SGXY\^X:1:[:-b.);49DRe-9Z^(FFcI2gZT<D[)9\QDR;ZGPaO.4B[_>
D28(Xe4(6V_UY-G9_P7V1(U2D57.03c?TeJ=.bQI(eV726946L8LWC&(D;ScC(3d
J1d4?<6ESEIOW?]KL8STU:ARa0Qgg,@cd4@eZ#Q96.&KV;VUX@>2WIFIS59P\^S)
a.7LGe)N?4B(\^aAS[/(12D38Z;.3EI1R&QG54KU2C)5e]LR7=Q-g-JPd.J<(C3+
Zf5g3c=GKG&\0^VKfaRbEHK-ddKD=M_agfA#a\g=T?2KJY==TN764@>eIJHdO@UQ
EERV7CPL;H0:A@Ag2Ya/VZ:>M+HPD8U5X.\PR;OAI_+RS6,ddR/EK71)F?cg61KF
JM/@(41N5PQaEP-I.CH#gJKIEM7OY<1?J;_(f8W&+>.P&]5\ae^,Eb&67T.:Fd?H
J6I1\2MVK(N-bQ@2Hd2Q>\59MMc9[11^a^/R^GW6da-bc&MUZ=/ZYT8g,&TTeb]=
f<#]\V79:O1\T);)O6Y??V:a7@I]S59gS4Ze_@aV/F?^1@U:QUKBGe#-PVPK4:)-
]NQZ._Z8-9YKR404/]H/fd,/R2bdE8C#YP7R?7-eUX(A6[MQfX/AcPV.+DP7NL6A
@CQ5XK->N#[;22eWH^2d8&@;a4:+.8F?8X3RBcY[X[SA-f0W[C1I>1RG0Nd)/K+8
,[A=L)(7IS/&U=ZII^[7Md4Z?e4)T\(=X:-8RLg\YB)[&Y)-L)YLb\O:eF\M8)GI
d@-;]aD^;^c8@(P?T92PMHRZa6[OP[3EggO@APZEQ_YE/K9HV/@9dWee^9e_,S5:
6>D5T_e7@\(R6)Cg=-Q4:Z<gQ-+;TT85Gb[+U7A/IU9R-TYdGaA&g;MFcB)O-X\9
EOC?#bMS,)5T.d\b6US4L5X:PWDX?C.<&_QEHK0BJdZQNH8cYKH&UZPA]DP<fLf4
?@DV+B+N6\UV>0R7I3RBQYF,GA5;YTe7#D;b/]GX[<R<1J,9cY?[2)K<.YDQTZDA
-RS;[]E?<a0DeD+^Y)da@-#a=fIBb[G#1:d4)E)]@)CQg9[\.QEWKPHYTJX>2.DW
eUfW2GM#++@7:>/4[5I06)g\.>;FXN2gF1\ICD]X1BK7PD:I>Y]F-<DHH)N9&W8E
.U+WQC#2_PWa8^D]G094139:S#3aHT<c,2DTcIbMM##cS\M&(4U;_\-IdE8GO=>?
.<dUPXRVf3afcE6fER,5Fa&)f=?9C.1_7a\Lf=R8[4D7c(-,(MX,bCP:M&--7#./
//=N9I])GWaZO)5>?-^X:ZW;g#YgLg3&TS;Q2&D:AfNUUP2;-:=B]g67Je@cU<W]
2=F^X2VBU7/6G@5E,&4J/M2S8[>:fLf3+WXe5490AL2EH8SfXBC+Re@FaSMcMWBW
\L?\S)LVM=eMeT-Wa_7eH-VER@=YUCeCF/c,bTX?4=)([UCSRU\SYD>SCR0K6SEW
^RE3AMCX@<JP\Wf2dGbO;:8UDbZ9KBR9PBeC3(A@I]O/UA/LM3/RIHJF^V/fR;fF
]aF#+g4RLLfCJR2e^]M3)2_90I08V0g5Z[:bZP4[:2>=?&TR>I1LaKdU[MSJNZUI
O8^6O]MKCD&fWK#EEdJf9Z/7)[FL,8KXTT^^@Ld7EcT;Ug46D5UCcgd.>2Md>Y6;
2&<\4[PZ0J8<gGU5L]I2E&M+:Wd)dc\[1cFGHb,ZX?(9QDD9RO#gF88.@bRA5Ka>
-T6V9;A#<cPLIIgK?3ARc6Z))2R)d_)ZRRDOd963gXSgO]Q:O+&F1:K9J5QZYT@\
][079H8d9LSaQU:2;LHJ]>\I)15f)LB8K\VA[VFB04.PV2L/.ETR/B^5)?EKWWVF
IE(\FRd@B;FGK9XfTLO__F^K)4IRN+e_T6d#M;Xd)W8MR#++;XN/0K[6@,.4_VXO
Bb9Z6Y5\XT6f]GHYA2?cQdGT9=F:THS8e/7\^gW-gV?GG3A-U,UN9H8+H,J-cKZ.
<KMIYbLUUeCd.C7?BQ6._f@3OC;9W.CQKLNR6aRPGGV@^bQ^\6=AR(e\CQ?_W<Z.
K<dCa8V&DG_+V]T\Ua<9P1?U,7Y#@JG-,=#Q5T)&__-b[Z<>3YOM=\7@)J_-I#]8
57[&@1<[?S6c#?1RCbI6&BZ#ef1aSX46S)(f\QOdBcg,g+2db6H=L+TK?H0@(Z?>
C6,H<5aI5\R;F0[+^TGY.Wf+E(.+gb/UQ7gTRL<,9<D5A<N4[4&RAQ?Ya@d.JH8g
7#4b/WUDYF>P+^ZC^be]&]3.f85I_X?0,e/Kg_R-bDIKG7dNgbZbV9ccMZ+.eQc.
K7e;LFM?@:>U-Z@Jb?EWe9\^aC3_IJ\Q?YGg_U?6K=[<e)Db8e0)8;S=OQ@b?U=b
VF<9Xd<d=6cI9A&MF<<fS^;Z0eA^f^f=N&aM1M;B]N.]7>^@^^[[C?adCDFR4Tf\
PH&+O)E0\0CPM<g:809d^7O-LR0A2RKFO4^MK,L-EKWC:eI:XQ.=:Pbe8F@VUZGM
UaV_FB+g2=A0U0Vb&b6Sc/gT+(_>OMc\E:1fU00;fQZ5737L1S,V8<\c2K+.JA<)
cZ[\S?##&]4fa&^EdD]5IQX:((6>L.[9(H&1IR[8(_@;7eCDRP#5L+3Xb@Q;;XV(
AP2g&FbDB)I9Z/V]@d/^X+.ISO[J9NT_ff,2S,.E_#.[WKK3\B42UR]>?e1MXX.2
a6EcdK8,[IKIA&6/.DDe&.\NaBQZ5DSe9D3#=QBf4^P.<V)0?]aSW:ZAg\799@M-
Ue+Y1Sg7/)5KA6a9YF#@?A.gA57J6e#D+b7WXX[R[ND77U/HDL^dCBA4@?>6OgfY
]cH,KHJ,f<ML-=Ra9PNIQSeMb-M.]]-=_)C754\SNAY9Q@aY^R[R2bDc)765FM@c
b9\MX(61Gea=PH9SL;?2H,FA@3Z=;a+X(a1:@^49T12=EH=&I/IQ/W;6,Y+>f)^G
\?K3[BVGe)YOH,JX>\WB##-3FK^K.NDcH@N;Zg8_d^27./4^YSQ(PBb2eC4<8MZ@
db:2#[6>>9M^PXL/J8)00dKP<OEW=aJd(<;T1=5[WAH)dTZg=+;f0Tccec=V;ZYa
-;X/;W7aeCH)C:A_YS54OJR?>]V@H.Df[aaW@9R9ab@dZ^=E7I+Ha5K7<\f7P?_N
>7\O,#g/@)YFW;P^<1(g=6;U.)gT,/<6,U/2;1fH45/X7-1BN1Ef8H6L&Ba8YL4)
RKS-WGDDBS>aF6N97J,BR^Kf@ZeY7PZE/.LE,HW)[/&Fa(O8V-G4>\(^JOK+4BT>
308#=\-0??fVP8;OIeZ0<^4X&E8gHFR:b2)Lf.2H2(aP,.b]VdDO\)-G=dM?[5>2
WR1[=0;<V=b2D[R>>Q0KU5OW(367&W[B7CN)6NI6<T,5[QcT+D1V1?(Se^]F.H0#
R7VQ8C32O=K\JX\=^1E+a(QDLC9RZ[Q@J@DH1&+/A<7R9@DVYQSB[cWVXMPX/J)V
FPMd1K6NSFVb@acf6RF[D00\-/DQP,MWZ@]M4dTAPEJJ=e,F/\[B84+C/)H8HBQ/
O7KMEBVX>_9WU-aT]:8ETF[C3efUQYT?[ZF)EWY1LS^EI+OR&I<K7bGP&_3VSNcF
J.H#f0,[b-+,S;9+2^8IU9D1VVT\L>=P_>]@e@V=D6/^Z]IHd+,+E2f3A\#0^1WJ
SJD4c8/SQ-M.T8U6XPf-:Rg@Z.8@H+16>6MC74ISJ&Fe_4ZIFU()6DBIMEXaF@72
]>;&>dUg=(?I+YEb3SF/OKL<2&UcXcVKgJ?FeSN/#,.43MM[T8KH45:[>OG(.4=#
B[-G)_:GUcMTR+WM5HO2QCM<N<M,HK4ead<+<Q]0a.,[&]aP>JJZFMbFW96VL38b
K?RW^<131P;P6TGFZ6&gBRX6+aMH/RgO1)]LP/aM\SK00c;#?][[9U8J(.0O:bg@
EeS#9\LDMA1IET+I31aRVd(_[@KU_X=-XaVBaL\Y]W&,67^Y[=8V=KLMGN70F-V1
@P[K[+Q=_-g\d5/b9E-cQCXKI:MA-N.WV^8+]Q+\\6IaYcEMLH2R7-UM.SJ^M1,G
A9X>ER>(S)M=/=UK7Da0[7#BYAG.,Z@a&0W6.E?NE].M02RN7S2Z(3<,aE6+;2Wc
#P^R)C3b_[L?=L/5Pd\3.H#,(E<IIeZec-QR+b>[&)(HP,7]D7NEN[eIR02_\J_G
G&D53)&fC_N<AaG&d9c8Y;>Qe]Q\FB7&0KH-0[g#agX>eP7Cf9+F@P_gUH^2C@PO
LfTQUS/VfQU)8)SHRa+#:::e1\\5V0E^K18:;A-FeKUF;27F]V\M#=f08/N=CK6N
EJ]W<_3ZRG>;0N@CU5FaY,Y@dQ_5GC#TTHJOONC>fg.VUJM^PDJ5R#FA(M5Q))K:
5U^[9C4=P(F^+_UEXZ,W/?#D_A9/[@J6Xa4:I,;PR[Dc^6LC\6<]&bf<7L[^/9\@
@TJ];UI7Q1Q#HCFHD?PE>g^:<)E]K,+fQZ1RY_G>62HJJHa,\C(PWZV<)8TSBB&X
I8AaK2=Xa#WV?XB#\4VRe@QX6.JU11V:O)bL>_/HGUR#3,LQW04/5f3F,bL^-13f
dG=5+P=.\cSHReV1a/ZafeF_e9<JWV=JOeTKS=;U5.GW,gJ[9OL0C?X+fPfAK,d[
P4_\UV-3\bSAYbKVHR:M,##B@76:5U):VDX)5HIIcH^((5W+V<9YI_A=[O(2P.,W
d\MgL(6QJ)1RHVTOZ5e.\42?3>gLd,]I.eNKC8;&;;@7Dde5WL4)a24+g;>P5GHO
ASI#,b.-SWM]#Z;97/5:b@aL]C(85W2BLbW0EX#fNaPE6JY0>b,CVSL47)PG0@68
_\8?;\-D[Gd-V-7NI&ZEK\gYRRK?9UH7ENKW&^P96eFSMbK;PJe=7QEeIBWS,1aX
(LSQeYAgDS4eU\[S@SUY,cQMH]]K.@\#V6Ma,HbT);,(J)?3[I[\e:g,(P<e#HaN
?cQW()_67-K>f6eW>GO3K4&>+ESDB:e+M/-Q_E(.-KC?=d=/L&N.FbfX1ef;D/TP
61,QX2&9Rg>]3:+UI-RD:eR]OEYa#[bL<SMEB3_TN654M7_HNUHJ:5c9UcRGADJV
4#]d1)ga;/>@gYb3XDZ8;1X8))[21(:ce-6AGb]Y/.e20G-3P=Z\^,]RJ[e[d4gT
SbZg@Eee)O(4dd[Z:Y=]&ffLZ[-PO[U\cY22U(J>RSaID\DYPb/IB32V9SM(J4Ug
;@Kd/]Ea&_[72@07/JN4A=9\3[C?>=D>LFY3^PP7?-bKT9]51J;SXCY,\<aF&FD,
W.Y^(c1^W-6=^>^;-a?I3S_7d9=(4@]#0X>[J1V-1L=c;cV&GJ3JK/UWETDI@d;D
1;SWFfK<_H\Na5U__eNX#.&C88LD1[.>&G(::[@/Q&ND@7g\Lg5S5f+8/2O^1E^E
YM:EUX8a#)0NV:NWbAB0-Pc/YZQ1:2QK-82&YJ3S4+5e#2KbWTc1U>MdR@11RRgf
9d>KM-LZ/OS,_dD25BB3YSYb4(1,PMKaP8S)/1\USP5d7NM:<8_M_RPCFOJV3cTT
Pg82+U=QZ@5EWI2GD\P=>L33bG1a#[F#KP0F4]X3>e;aQ2JK]?-?fX,#3X^EHa8;
F&G\78V>aW0D5V^@1[I8EH;7WdH7(1&aTJ5_8O^G+g,V6S+e#]24T[,8Zg>-]T?F
e0Ue8JM-4/67#1bRS5OVVbLCaI@4FX/Y5EX[MWOS5<d05fUaC;IaQ2Sc4Bb>#T(^
J>b0VVP.C7ge[LTcGZbXP&1-JQ->AgNag&6XD_A_[S?R#FOTQZfOcSdYD88(&[\-
JC:UH.2>b=V&9M\WSg(3R<ZKaZXS1)UJ?Q;2YW(4C2856g4R#c2=:F53Nf56,R2=
DAc[bafgd5DcbN+11XEDeY3J)c7:1:>C_/8LG30fPQd?E[9<cE>_Q?[-dX061^.]
A<:G@VSfRNX8F[EQbJTJe[AT3A>585XdP5QD6RaLZ^4TL9CCBd_L\;7EaZS4+1g)
R9@#,2,P5@80^O8OZJ7=BcdaHX[,Jc+OR;2c+^ZVgE1#7]/FU4(SF6F/I,YPT:Df
,g\2UDdN2T\+8g03__Z@?\NXYM0E/EDKG@41f1\5B?3N[^-D_Ef2?3P:()<&DH=f
^(M8g8Q]HRca:,300d0Z0_FKF?G]\2\#AP.NdS2PV:8#aB(g,H6WXU2NI6cF7+TU
/2MJY5K3a^<Z.,E7OE@Gf?g>K<B2PN)HO0-FH^LWSID=c[[CW\8Wc(4]ZB40gPKc
.3Z-&@e5bSF(F]0I898;e;AR[bFWI8@+_0Z34(6RfB)+4_g6=5JLcC+NdX\7E;S5
dX(O]U//;VJW>X&7O>G5Z]4G1GRGVY>17GR8LaK4RJ=LQa9LD/5Y99E30D.d+\87
3F).?XN90#1LK;ZKF_MbZ/b/&5\V+7E4fab9aCV2MMF\/8ZD)f5Ia[2dX/-A(;VX
U^6JXc81e&a15f<(CCS7:>T4#6C\LVA0Se41:B/1FX-V3g&g,+HMEV\HG#+4BA07
J10&:Y/X)6#gT4,=GC6@MRZ;]A=TV5(<\(U4G=4N.#)0W/U#4[]94-0dN/XC[7M0
U;8:Z^M/T+V0[WM-Nd9:<:>7\81/]^=G-;.L;3CG39@#=QD9#Q,_U86X.FeT3TN;
Q=).e0dF4_&A[N#5N\EUEa,4HF34cG\1TN&O.4?_<QS4>47?MZ)2WIT42fBKDeaS
_SPP7:b)G_A,=#^I@b[1DMd.]Z8D40910:8RTWK4KZ73+QD\P<)6EKcSSAX6_6F)
c&Y6aW+8PBf3UZ?fL;/^R89Z]NgAYPPD=<g1^]O805D0ccQB=_X?A-9Vf&Z@5K7/
\U(N76[G;b+e:Y@T2:X_DgB^R5T2-MCa7GdMNNcI5@[T0(<H5bM6>T_@O[(_0YIg
YB(;XF=RZ,EgJKMDFCAK_K6D;R;e:abf&c;HRRga0Z_;&/ERCQ8PBN3d=>I#[]bU
C3YL.C&#Y81g9\T(5-1f>A>6<g3#K:;gN;.Uc7De5B][5G?bcd#TM(7]bV:2a4[>
g6UE/01gd^@9+b69;APDbcL+/VeJAN:aR3>QCB94:[6@=)R@P=C\eO-[/d+?eP]^
&]2YAA?cE2-BYS(RfEcUXIf>Ic9&&d3BV=+XCU+<SHNZ&\/:/B/7&gP[>)AFeH06
RA;DWbP6\RF@gSa3)D?_.(Y?,-Q<:OLG?V?FI_@(XNc.=_dDUbSDO[>R99Wd37Ae
XP)@8#7JN:>R5@T_OTb>9UNb8bG=<<HVI=T<S8IE,SWU-gU&\AD?=Y@2U:MR@[8K
WcJJZcC-_(B1(0G#?\Z(I:IIOOeJ22Bg?RL>eY>>QWc7@I=U-.gbHO?-FP&fE]05
<J[#0ICa/Q<J88bB5W#P[BE(7;d6L0]=_7,d&0fg.HMKJdfV;d6+f)Q]>2>a<48e
gD+7eFaZD#)5+_C>TeB_OeY48]&Ee0c5-ebdN>@4H@F+/2=:H)9_5:;BC[8D^ER^
YS[>XYD8]#cb,?NC=KOD-dJ-HB]&7Xg7=Q0gTID\Q=B;O^fb+YYVEg9S^UH=86)G
;7NZfRWW0F7<Wg5f5CB?L_BPf_H?P+-04)d&S7]LNO_=UEGg@0BdZRNgH/LFMY1W
0U6W>a52;QZ.J<#<fdYI:]<69XGPEg8GE]Q0Pd52)HA+K)c(W&+M?6L]]?XXfGH(
\T?A=(ARD+C:UKG@>=0A^dSW]2)\c(B98H]#A=IK;^?8d6.RAXEg(8U4Y83bM-cG
O>gYR<^CNPJ#-AKAN8cXDI-/M1^O[.(2_3KUbO7Be@._)XX;TLHIbL=1dLd5NE?f
Uc1S/-WQ<9@Kb.7a=f2<04DQC9f,gP5/,O@2O7#8Q=f)L.V^\<_SV)LYfMXBYc@R
?UWF_;<9#TUfVWeHD4+\MbJ&);;O)1G@PK#WJIRSd7V[+9aC=FGN\;;?N(3E6?PO
LM1);1D)99=@_ZZA1I7a,eA2X19:GD?,<#LJ,8YXZMTU6FM\JNE/:4L]-@gIY<Y+
ZD[?(Q>QE98G^<UEDSA.432TVaaFfEB2LF7E.?Z4I_,aK3SD/<Y>Me_GT7QMcaB]
b[^gNZ_7[OT#b#KZ>631OBK?W==,=&&E2_8ee,=I?>g(UU#5]MC?a&2]GRd-3fSA
7<fLOFXb(4YdK-><gHG5?X-,XT2dHUf-^)I.Na:])a^[2P/OV48#9X\c?4&,Sc7J
L#f/#Rd[AGA)I,&[b.VFY0>+39L=4[PfcQ9)a-(gfY\5g+OZc@g4VVDN]aL0[W3Q
JCB1\<].?053O6,,-KXY;)e@_M,>9Ha_.,[:gOeI(5-4<RTH&cB+:[4R\+9^800F
:7ZVDP\P+/9^6#KTX9U](0^O(,#WI>TKS.8GF[,b;G&WBAab#Ac5b,IG@W3/ZYS6
#_d^aE=g7]KM).-?QWX6:[6V_)+bdG@=;@JCJ&A9[D^&Y(a^CZ,)YZ<W3WY>#TJX
E+85QEcD[7f_ET@&7H[4=(-7-A9>EDLW<<&UIROS7(0>+e3L?=?&J5A^\BcdU:[M
bTTX)=W5e^S;Z;T+152-PNOG6^T+1F,NgDMY)@MW3K(3,#LLU:[UCR9R_M8YD22,
b[T@/SI/6R78WL]T;[E-==L?9TOdZA\DXB6[5=?J<O2,-RYE<?>=T_K61(,TH^TL
2P116M\CPcK617/4e4F>fe[V>-AIf469@./U04+fb?Y+W/J(dE69d-L2DO/FA0QF
3(2_TAMU>F_VcgP.5/^)G1Hg7UD#=S7H:F>N<92LTJ(P_WGB[4UfJLf2D);.7WY>
E1507LMLe7g02gJ=Q+]X:_P,GTG6\5:Dd\45fgG0JY7)/1>;5HO#0A8,9]P2473Z
E&2TcbWQfTD?VbdZJ)NXaM&7HE[2VbKMUU.PG><;-4Va8F6f#Rg0JOeJ_,SEGX8f
J?^7X\_DC_Z^=?Vd2_c9J,W5WAc,MZ?;7M;/8UMV<B-LAEAa;(&^FUL=/:;b,3Z0
U.#W1UKQNIBDUc?RV3U-20NSR0+0.][@E^OF-SYf)PO2H[M<5T2@fW;);1c6,(&N
\ccK6]\T66SG<V[f2Cc5<Y?XR<M?IKY^Z5.aFK-VX3?I(7\b1XFa5EZDYD_B6M?7
1=AdS:PJaOF@2;COC#(];d).d?1cFB[-RBPdURE@<ZEDcIM<fTSLG.&QAE/);#g6
LAf8E)<_HbB9W]C/V<SVA?IPgWdL6^_@]S@3-EP_<Y.UU\:Y=IdA5M\GQO17fH#N
1HA,84?J2<>gG\G:DNO9N=9G\,:EQ3>bdB2ef<Z_K86YCZfYeA?adFNY/<g7Y+2V
?R5I3:X6a3_8A2GLO:O3UQYKV2\He,Q?2[0VD:5#(V)/a5J+C:1BBDg_9b,e:cP<
8J=-L-GI9-.F>E3H?\a,(53U+(O;0^#8IZW(RV0&4=O(USO_6A88H4Rag>)VfI;H
,L>5WFacE9;TD6&bVP_S<Q8LB5@OU>N+GC+DcVI)5BX=._+\>faZ=K(SRK-f+b6X
X7Z7,R-XY-Ud=R5J.B]g:U]S#DMVf4RZB:,A>5gPfC^\R^@29]9\c/XO,4#gVW_>
SDUG0KQHE4RCT?8d#B:W_=_:,SHdZN<V#RPH0PbFIG\,&Qg,G;KI@L1Jf,Kf#;Y6
3Pc\EI4B.RcG<:FeGF2V)_0.Qe1EDZaKB)7aQb@NG;&]cZO3K>59Y\HH(2bVVPTZ
38L7EPJ##T]0I&&&;BeFEW:eb&,_e244+(>=OcTNET,ZR4N1-O21#A_@/&Z;2L\J
F41FZ7ECAT_Ogf3G,X^NJ53&>@D(@P83VJ/XYJaWV.+d)Y^eREQb+P,gIfa1#Q5b
T2PeIFBO&GP,)EX8gf30bg65E>KM=egcK[bb7?9.+WFQ06K=P^\UPW.M0c.P:/,0
cLH>GXUW:/7;KGFIN4f:>4\PI8X1fT+eVHbTPW1O:DFB<]QML(/AWDBAR&S?\Z#R
?L1P<\)?6Jf[?K:SZVL/V,U,<]bM;6C](N,T&)c]=B#\_EMTDdN_f86Fe<RF).F<
L</3>VXX5DA3PB>=Q[<:ZF;J:AG^aMB<B81Qb,A@eI.0EPRS=gO:OVbOB8H\IU>O
f+8C^P9_F:,-1)g5836R=O64:Q[^G8A#GV.LBK>KH08(Y(=,6_YZ6Zf;\A_ZTLd:
XLag,Q@EQR/C[GaF97H#T,_>L3NJea1SY0#aIR4_F7,#1E_)G4cb:cN[PeOIF(HC
5O.T-Tg6W6QU36UT@HZX&@RU(R+CZEEU#/I41O_;bAFP0H0YG#cUV.W<E><N4#V0
c,]G<H;7gGY^34;fdEI=ZDYe2^?_8b8?36a5FW;,;ec&C-0)1\_.Y84?MdW&[aDP
;Z7?CbGJ,a3.HaHS(^M,4VWeQ/E7dD6:7@QX8=QBeS?KQGW,>94eSR9MXXV#V=PT
F\e4@JCQN@_]U01.J6RRLK<;IE>2(LKC<LR.cF+)\RL[MM5Ma?.XK0VN)c(FDRVJ
FRESRK#YQIK=9_9OCE)0QGV5FE]aF?Y###5H\&O=:]C0#)^>XL?JY#Q0d:682e2b
]?V69b4BFJ=;ZH&N?Xe67&(-LGfc&=;=32I5D<]E0,G1KM:0PBDW1-,V<3.9-(6N
8L0f55X56MeKPS.H#P1OJ@ZYBQ3L+b\BK8>YJCa?)P3P,RFF(fSWdDRW;1A/dD>A
_^ID+[@X5R<T@);IJ]T5?_N.;;O8Sbg@[L?<HG&SC8_<O^T@O&>c1M^SBFU8:?)O
V3c<;9SP/;N1+H?aeA6gf)\I,EB.:TQRI;1-d^7A(,g2M=K),_T]CZKW?:=dM,^&
37d;8gIXUH,U[\8/_HA0&&cH<g:D&WN>K.3:UD+b7E3:CELJ)7R908,TWd(&e-OV
BXF4e_O(]=7Q:dLSJZX:FHEd9I5BX=G^.BZ^FA0D6IHZ@26<]OP)>5B[b<Y<2:#<
<>3&2^\W/(^HUA,X+?:H]5S#A8#6aI,:R3PXJ#/F/>V#eS#2VYH<F=eZ[C3(TcfD
e.PT\0363E7Bd9<ZSJ#)Yc1D8N=F?BJ\0,F79cKLU:M-b]E4bS;4@=5-SW3]+.[:
>+KC=Tf2:=(KJQJW\[L4KF_ZE,CHHNFCA9I6Nc>J7C^[667I8\X.LVZ5UX;Q[:-\
R-dHaP6Y1VBT_&SA1^5]Z,/f656L+^KQggfLZHeSO76PI;d3>QCC1>9b:&BL:Bg4
Q#)[WROXRCKf=;L5e5a70>4L,CZ=6Qg,MN^^<#FU+DG1[-3L;ABMg-Afa+IO_D(V
PJ?0QT31db=T;5)E^TQM2^8@X>+3#9<_645@<H/H5UJ&5CS]-QWbT7[])IBFEBDO
WX<4S>[;=:7bBCXb=C2FOI?P<K:g_](e7IXGeF+9PEKc919bQ(Oc6MX78_H+.T=.
A<>W48P&UZ=O^WIg.CW?H^@?A780JN#g./7?(S.>Ka9Xfe=-d86?X<DSDfY]BVVF
O34M?._/G7PDHBada+<B:T&,\:[RVEdF9d4+74eeE3[B@QA?6LTI&I:J&;.&9NXT
<AK?cH/:C(gZ9^BJ[/_MSbM7=6]CLLfB&HLGGET</S^-E2J,W;KKD\bJ8#f=e#50
EAGW9SE9&,#[G;&-R+N2NH&;cX?[cOf3&+YB0ccUGHQ.VI\:aQOW_FS\?Jd2\[KM
K:JREbB8b2+-]/.I2,3V&>e=/5;R]HXL5X&WA>9P;ALb<?PZ),(W]L7HIbW&9V=S
[6WSe=1V?\E\DQ7e6PUE-CKV-X_/?@W:&;4<YZ[c.0>dcCAS>c?H/RM4_V(4#PbC
_3V^EE&H8,X1>5Y.&TWS6OUACJa05Jf.f.80g=1>g<b.a[]3GIV_NdUZ7V00G@NZ
YT6cSF.KT.[IH8R@#)[3G8)W\Zf-+O:eF6VQ[V[<Ka[A+#g197g+:g9S7@(7J7BS
C#d7fEWHIa;Z#+S)M=#_-e84:\?UI><AN.e)H8XZRgYH=;[RA.=K5(:(<(]X75YM
3S.YgA/[?(C1ADVL>1cQ?C/AULNPE4+9:d8GJeO5^AF7LG6DFY9(eK=3U?\D9@N2
LK87dYK\YIVHVWFD12[TM>08FEN_LTTg2Nfb6W4HRQS?>XfP\L_g_AQg,7D+S^f@
08P)8cGbG;e\<7dTBK,YZ/7g.X48[E5=7gS3ZPDZgTOLdE+[#eVE-5AAU\?R3.?H
PP,;SYM3>^&OXS,JYO06@-S0++\V1DV(T<5gKDR-=&ROO<ZVOOCS5MH5V6_=@\/7
BDLbLRfSgD@UY?VWA;\18F=8L??S<;<P_=@TF\,\QJ;?dI_6P^UI[eQ1^NP&\T1W
b/3:AId>N-2421S.8U,Y7B+)&T[ZFK4CN,]N0/R+2CMYG2gDTG_#VC[.XO5HB7<X
7<FH?KVQ4+NH>TZ^acVNY]+U)QT>]g/_K\005MR,/eA41E_ZD+74=Y0EEN\ST(J9
Xg4S=(\bM?(=9Xdd]6,EfKORZA;aP^IV=RC\1IVEJAPbFEdAYYBPJKR&K\.I<9Q/
ggQ.;<7eLSP6^TfH4BaU<(F2NNHPaR6Da^XX3WWNfUeLdWg_7V.P+\5R;PZ28DW]
/FUd)gVQG5/gCBgDaCe4-W:-I+217]]J6HZK^<KXd7,P?Q@f\B6S7cWVaF(VEEb@
^RUJ400cfP.[NP>>?AJ?XP5J4fgd\1CYZCC\63:89-W,-M&.CT/bg#7^<1RgDc5C
0gN](7@HL[=aE^2YHP@KWeVVT\/?R6.#=1P;SGERP2;G,>#,G&^3?/YLf,7RDE5<
L1d9@ZI]VR.?eRM-P3gTFWWWPYW)7&[Dd/.B3EdZEW#^5MU[]\>A9=VcD/JHK(=;
Se#WQL^,50)c>P0UJR_U3AT5+]:.2\9E)A_M9.FRLQFF)0].V6YU@G(\P1d<7aAJ
P0#UN2G:c?Z,7511M;OTg6J#f5O\Bg:F]#Qc=?bZ<S^@bXLebJd8Ob48,B/MU01_
22LYSD6H76[2HZJ)bILY\F?-/FUXb,+dage,?M1KWXb;=@gGa@7d\.Pc_HZB_VP?
UF3c&?f2W@?TMc>Hb,(N.Mac/3K[eZSGFOYR>T/#Ab,.EQ(_>3::KVdTORdE&BF5
H?e9[]/G,FfQb#@[,&(LMNeIH@ZK#\4&^BE>-;gPBV/_PRRZ@V\C:R&G[)XU9W@N
d(>E_e;eVVPR9[Q5VRS^TJDW0\)B,W3:FO&Y;3=IOZW0.YAZfb(49d;Bad[@0TJ/
8)g</GCQ5S+Y/9]Jc3NUR-Jd]IbV06/S&Uce3_ZX8+fIW?0VJ)ISZR(_8VOeOWac
YMF8];^7H(/@6d8B:@+^eE39JW?_UCO5,B^T&5a]>>D82R_WMVQL,4NNcQORF:XJ
174RV7XcWE7>FIU+UAW/)R.(OeSTb5:APZcN^4M,;Nb:HY(L/HAXQUWaf4A2HS#+
;#9O\\<:(>JL,VYJ\EbBMcYY,Tb+:&_5SQL&YO4]<IF1C;2EJL5^T<FbUBeFC7\\
W?+#-CJFd7KW-N;<1,fe>fcU#?gT0[5<J2b4(0YdI+N46F=)8#BagTE8]WC_bU)+
UGIEfJNAaVPR;d>B-9T,Q&9/a974_OOKVV?OGK^_bd1=:LfF(NCT9J=]Z>89W>WD
0Af<Pa>C#F:&MT\)S\US((N[;LI3\c;YKGeZfD:RZZ=a\=AS&S_#&M<1&>cE0ZDS
A0O4Y&MW+TZ3+B@EAIF[\C(QU<7@+)#@4]\X.KEC&gC9BG_-,J?3P/TQAVf(ZEE?
4.VcW=]9Jfd<,B#S11@QeaCR-3K<3KL&^Y+Gb-d]+?C@Qeb;5F_W\Rc:NHU=8DVX
:=T:H@_P4C^WegKaKFE[AG.LF@<R=KMGWd((Y?(OAfAG;e,7E0=^fNIV<4d+7Z6Q
N;1PRY?0RIA?OHYDV.X@QA&:R(&6_F#e;db>&Eg@F2]G<FN<fZ8\6UR6gZCQT4:=
2GJ4O+TIOTV1<YE,<VX-QLRdUD7@,Z^b-EYG(5#J?W^.<,.e?X?aZT6Jba1>Q[[(
JQR8A]D0X^7ZT<V,e>M7?7)gK/OZf1a3OJEEOH[GS3GKBWN0]F/ae8<]N7fH11E4
+4[/1&&:EP>X,Ac))(#d_ZcSUVA7E[8^XE^GL=#2d)LebRGRVZ(d8e+;eO2G_B[N
.3Q[Q]f3=3XRL54MUHZLL+=W8FVcS>c7T\..(D\\dPTb5RgJ:;2fR):1fSScQ4Ta
1a=/DdR/&LRSdaN>YW8_9^eBJU_@S\_PD:>_a9Q/FVa_U#K9(5F4,NEb8JRM;8>A
egS_Rc/c8aZCFRb+CZ,Y9]fL@0^O(V@?/AN]G;AFT)4c=CPS/b>#0NOA:aDJ_IV_
52G(D[NG]>B6GTacf4T0+3VKRY]+^QVV)@>RKH2QKTAZ;g,K>ON2LS;4HC41g.^e
edD:<ITA+4Y_B1VD>#2gLA2D8UAFI5S;07aFA]IMd7GYgRA\D@_N[bK>Y_0?J-RV
&PgaD+E#>A;32-G]Eb1K=:0,)^B8?99_G;H_T0G:B,Ue[<UR4^?3@dDZ5+RY4LC?
aQ)b\;3Y>BC2?QWG=&dW-^d??F.>_eO]:ZEd71M[>C?:bT]0[24&KZB.eN5N,-Td
K3PU+7@?&;V6(_D\OAOgRJ#H6&dIag6A:.,[6?Z(]3#_FdbAMSV,YZ#82XV;BMVa
.A/^S=+b3&8@ZPV(5\+Eg8TV:A(Q(1]WDIf.DFb:J?-;CD6JVR7(ZT3@Q7EfTF)f
7;9W7PEcKNDJD23=]<15U,_AGG\=R],R0+GT6/f738Q10@+L-eRQ==[H_=A)A4@4
VK4@.K?eN2I9&P48-+QJ>G<d7N>@.eUU.=b\-4T^+J,/_FSS3UB1NI05dH)-^cH3
c.EZ,QeO/VP_[M?;KUL2EVPVSGD_1-G.>f0a;P;9ca438<Aac8D>+?YIOV(&&J=9
AD[T;X/BE.+@;H;a>N3[)+_;FDE@eO-]b1GZ;G&\1gYac9RDCOdeaR,V4+T]8O,J
.FW88IbeG)/<JJ(?187^)/.Q6f7:g8TLQ;#OVD9]JWe3[-UILYdg9K>TR(?<AN\R
bP.9=Q=Y<U/8O]T)(<O098>1cM/<:fNCBB=:>:3.E)XFG0d(_UA#e(GI33:4KPRQ
3-XbSV#TM-/N<gF<R0@,BZR0.MGR,UEb@LS?J.6)IZU>S6,[MO^e<9H[9[&-AH(3
0&SIf(f2a??<2KN2#gLe<-17FeN@3H2)R4.1155O(S#1@<6<Wd,13@_J)17&UMc8
f3/R7_QaEX&TWa=Z\]\L87S3b.FQ^TSW^F:M-EBfLXCFg/g87GFWL;He/#0&M[<V
U]4bgU99OcB>:4]7HI)gJU1L>T5e(U<(G+_MXLEH-U0D))5.bLT>U,@96]f>&>#@
c2(^9T\^9M8YVGgHe3Q_\L&P6EI-5+3>10dWR?<_M.G@cNKegAHZ(Q\A(FVg#QU)
+>eCa=.NL<FO9O9P6/5A-4_f[JC8^=^+Mc^_8]Q3BBB)M#WUC5M&c\T_W\D+_IHZ
.\NGQJ^/;_QN0?95@K[X:PFG@K21/I^8/M\AQYcef08PL21)[BW[R3=BcIYDP:CR
2M#S::TJN1]:P;3XEQf.-E<;e+F7(2P+/Dc:UXc(Vfd;D_EGO<dS\g^SFMP-JgH>
d23(F:<IbJ)BCZV/3ZA<e3L[35Ea1c>.],>_E&5_5H#9R,14A(O+;DQd>XZO].YE
1+N.FYXb1C+GJ4Lc[=\L2Z[UOR-fJ6)WCJ0[aQ,8/F+;\L01FI[1bfNdLeQ6KB(D
FDNNVW/gOZ-H7PDGY0K-=BIRb7+L-;3eUP]a]O6&>_Ie:IK].29<2=/T#a1T\=KD
P<_Q4/K)_Y\T=MaP-[,B<82Fg1XdOaX/^_MQA0fKWR.Zd8\MU&3X;5Laa(d,>O:f
12U84HV392#P?<dF/]=X=>VA_0:B0;d^fG41c[#O0SY<W5WKAB2(18GL2(6c^gYF
LCU^N,OSe]GfM0M-PC83?<T&.7WT3.X#[1_[J[+dT)I)).f?C.:IbIeC97.c-UTg
BEPdO^S0)ZJ&c@_\\_b4U-;MP3^]5;>UB3_9Q[._8X;]0S5AK5GI<-Z+<bJ#DROY
;#Z6=TNe[@X76edNCAZf_+5S#_?-1c_D-R,]STa/,AKL]MK6BS+6@,/_<[=-WH^F
36Q,>\c/?[Tf7<9?;4](9(3EbA6HYYHRP0LYLA2G6FDQ@55[93Pd=gL1F5C=SIT+
G3b2NOM5SZgF>4&Rc;O?Yd1@Fa9N:V1HYL=b8OWfG.#<#+W/X\7H@2O;,BAa^<.K
IXO,9_JgUK#8;I3[M+>?VUe\Taf0B^]baGdeQLE]9G9VNA(6>ZU.=B=:+CQ1DMYA
>URLBbK[aIIf9X>^bUcD7F[gJbZVFDGQHcdK1\dI.@Ea?R8:(fJY(>.JN(:=(-(/
[,]EC[B#=:egY_C)aZ37F30(KW.MZ&W=V4L/O3)c[a\CQRa?03@5+\8U7+1c.OZE
5_((F_-C796/P@XFb6),CHNE,5c6a>3W_TBNL+BHSMTe16I31/0a35]Cb8#&)9&;
eXY8C7EZg>R6JR><W/;8a^b#^[A\@2::3]?ce_HdO_a7EL7:J;,ACaJE]]/+>Bd8
f>>99)A[TPa#T<9=VDT(.ILFQTW,(W7X^4<L([)B&A&J;Xg3#<XE\(E):SQXd9ZA
.4_]N5P/-QQK1JI;JecFUf^Wf.F3d[PNX,CcTG+W/S8LLSEMNIf-3[]4=AS5B_Gf
2b9RPY_F5&GGGDV+[(A/Oa.S&V-,<1M1fa733#8E,GSQK\M<:@R@TLF1cG5LEdE6
g,71B27C8L,X.S33:8S<W3B<)D(Uce3-^-OA<&6M=JJ>0HXI0dOCT.RTA&XY]/gF
>=F7#.\17g]8CJ&C/)G-.&;]BdJaUO0_J620/<BB.eA5^EQaEW66)CF)\ZEcSVM@
]W.,fSF)-LS8S)&f0?YOI&#3g<ag3UV0OQMLI]e)\&C#)8GFcXc1(e_,AW8N__T<
8=+M^;;Z_\O43<g@fMV^+F+fa.?_40C/,,U8T>XO<NUG74#g0[YVMLJT>D[Yf._Q
W?#/fH]91YTX:W/>&R((;D8fUT-P+>5VOFdWbFD=IQJH00\C>XaGa,.d/_[A<WOR
Ee?Q5cCFIQ:HOc=c8T1dQ-K47e>LG:IR\e9K&:)FA&R[2(G9C;g=@N/BGRUU+^Je
F&Z>>0c6RAd&c-?=VK?WR4XF5T=]W0gX+B57ECP=Y=N5Z8HIKe_bYKg>a[(XRF9^
YIgR#456X=@Mdd&-WbFP..HAN7HdR)_TJ7/<cEOM,6I68gQ-_/_1:a2F\&RgQLH9
1=^DG:V9W?G)78@M87a)22Z-g6L;e?;>07_=3DPafVWcEBSSQYU>VLJgMW8(2Q\-
UA5TT\Q#[\^VA]HOf+V5.^+V@D?(Z5ZW.[c7D](3B)fCDZKL16N5@+?0+=9U=BU3
WI68?Oe?+6cT_<,+2K99W)1:EdJ<gJSU5GO8f&)OQeb::]18M5a(@2HO_X8ENY=]
4J+1<LM6W]776B(?N_X1RTED6X-N\Ca31,A789eS1Xf)TJ,4,A]45XHG0P=R9,2D
\AAef,E7>BL=VR[7WL_622?EWQEf5-X.==-(d>.Lg^>[?/b5C3\GdW?<7\=KCE].
&D;XJbNQM/\#3--:\]0IZ^>_<_-6J3:e#7-8)agBXT13CaXN;[_;G_:_=;#)QKZ<
[/eI2\5>&M[@/@_S[_1M0MdQQL^5&e\AYZ#I&&6>Ne-J3cZe9Ce><NI33&NKJ+ZL
#@-=_#3DbcaDPRH-&Y-<\BU&MM;(Q1W5gAe@5;>YW8];=/]>QS.))ObDHP/EG]B#
BYO[]If575gQ.U^b.&P.M3&OV8[.O[R50)]HU_g^_>/<DS:O+:KDDe[P]?]R/L(b
JYZ17USGN_HL6:?cW6LROe?fD\7=d:LG1.);UNWUD[)9If\0aA))LWaPbSS&-COV
<G>.SMW<TQgT:2@4_ASFVA?&?V0^C\(]J9e3f5K:W4<UdX3MM/;QDE@52];O1?GR
64.M4bBC6-#KN^?;#[d4PBYFgfSfI_=WHI;[?>L[E2KObTC;Z0=EcW_<bWH7,T/2
5->3d2;_ac#QJ#YW@27=TP,H-,<:4:Z6Y<<TdJ>H1QaX_@@82?^G+;Q?CX)2A\O5
3P_+;)[4c:IB1a6JX^)agJ5;_@9I?&H)0]D&;[5IRGOg@^2gHVX7Df+.\/4@LZRN
+[(3PE9[+aRRSTA(8F/@5NPH_aG#Gg-2:)R7E?cQLQ/@\X(:O=/d_>AO&:02bD/[
L@/e50\4G^de5_-Z@UPU>2JHe]-=?c-6J5dO;37?1Me&I#d48=8QJ=0AUBHB=5I,
DbYM\9>Z\X>DFT(]G/F&BeT<7WIZYN\CKP[Ff[\,]Cg/2P,8&-+>E1YEYgWb4@J<
#1bA/7C-8#\J)P(f]-de?J;YcSF?6Z]VG>GP:,/-DSe<DRJ]<=JfGa;^EPH+Ee(L
<A99)FfE)=UJ8LP8<W-YA2I-8[Sb=7>E)05V[T]?;,WcCQH2^1LGNYU?&AWV23De
\H=2Q<.;b?WU@OP]9)Hd1W=>3JL9.]&L[;CP+/IF=K,@46:^SM8(+T5R446.DVb:
4?a+WU5XSBZI_#/Id.7eRE7cc<X]fMG\GJ(c.BE<M88OZ\SHPZ\=Nf(W,MJ,CDaH
BBdC@WgODd]RP]=GU<;4;AHO,\A>5egK5McM^dC)S/9]XZA25VV\C]DARQ28(:Y]
BNc:J,edYATcGO++efXL<F>dPL?6>ZfdCYT4Q==#acgS+Wf5J?@ERTJb72UR2:A6
#&D,^?f64I?S(#PV+I:M>e>+5C1:+(a3N(]CM&.GCYObX)BS>+5aZY5ID(8B(]5+
4W6.^3dgC#7@Ka@.5XMOMCRG=cKA3YLLB1M.]5]Xg3cd.-)c6V6=</^@^691,ID;
4UAE;[;C:_C.S]dXX[6QKf1YS_J#VK>SYIO8d9QCacaWOGX->14XTJNceHXR\1bD
JdW..RBF=<1WcAJHN2;QXL4PD-fRa3Ge,T6bS4T+We8f+?bIG2R(0WBf-WC/WEYY
6f/B2CV9(X#MVFPbK-b,<KH/GeE=D;[+ZfFfd.@307.g7OG3DOF;-ZJ</SP1F)ZG
F)[g/>f5T^(CZ3@a\V_EP;1EYcJB86=+(Ka:_Ra&H&F?7.a6=A,F8)aXUR-ES,?D
4a7Z.6bfO-/LNYf#&:X]Z=G,2DBPW>1(F#L..?9H9CE_Z66#K<B#&g7;J2MSb@;I
B:JAZD0QBFNe5@bU]a:5S2R6P<6BE0(>8[fHIVV=G@<,>+CR)A30)3Q(,7d-6dc^
Y.Ob/S+9JeN/26Ifc_<#aXXXVBa@C5G8?/Tad_fE:7?8;YD\H#VR>&CD[\..>V4A
].U.@(ec^aME>,3(G+@#2[P5^HY7f)K9=g9a;1U+JB)OWKZ)ZUJcFA90B]T8)I9J
a8:bXY9d[2?O27U[@S<(&FMa4Oe\K2L<84.N]W@8?Q/W^J#JN+;7SBF4#Ub9MWOP
0g839X@eQ.e<)1c1Mb?K;X=\(SM?JSaX<9c[T<EECbERQ^#37PWb[RZ+0a]URY;L
X:ade?1McZLS<bf>Yg>KRP)dM8a9D5C[C(L/&+Vg@512;6_00=CIK>CN.eb+<3-7
a[B+CRD=H+29QL9==PA#R012Jb+I&[IVQD@\0;BVQ&6;.Z4O2?-&bZ-6J#2=]F4Y
A\bB&_Q]3e43EGC:9aUV)+eIV>-1E1930P+dUCG^.30G.0+b:egF=IeNTV0G(P1G
,S9R?CLeeY772;D.K2T8-/W;/I)KfA\C_8=c9RA9>+KY-Qb[C<Y:f/@3/0gU2)D+
AYO;ZS@HA^<R,JLeZB+(RgGMDAf-N.HCO#UDe;XE)\.@]:4QR-(_?XYO8faV(IE9
X8?/7e,B>J3,K7ISAC0?dO-ZC<&<T#)[NT1P(\R)9YZNE?NKc1=AAB\],Q6.Ea/O
YHV^OeZCG#Q_6O?0K^?2&DW1<0]Ob^C_?eMTY0&TR,G3@<CXX1H@#fcgYT\TRR.E
+ccSL?\\LbW7&TSXK3;D7@IS6DAKI+/2+LHaTD1R2>?I@B>e19QMHI1PaJ7)L+b2
,:JSSKK=We15M)@d3^Ma6f4<JU-05CAfVa:6(#O9BW8CYC+eR==PgYac.5(XeGXW
,EG3F;.U]1U_70XeL4/Y^^)#<^.GeL0\WPKcC=b;ZD:.3LE+7N5f@K[6R?KgVOWN
O5d[CQ(^NVJ7(S?L6e/_GXV33\,05e>1CcQWN63R4VgI2>QCWRgcK-;=Z?+(XWYO
?/#Yb[SOJC=#gXQ9cU84=JN20Y;,)K[;JQE3._?-)bSDcUQgAd0>3^dd9/B[+J^2
4+Q&ee9W;LG??F5?&T0]:Tgge#/UKHQT#+HS600U<F&6)6)\91)M<ZJdCf;4YGXd
(3cSGE=>\bGe=TUf(J?UJFJ7V+g6>+Q6GK_N,V1O:Q(ZO)Z&BNX2N89aQTGOb(?F
F;6?&5A4b66bW#-PDF7P]1SE4])(JcK=E3XQ)R;<b-<e\/BZ@HeLB\\6\-BPZ3\e
MSHQ&(gMCRDN2R;KU^17@J(FB.d9GF6+^8>H33gX\UP0F45L&-IZM#,KIF\g]P:[
<&3S_TZ4=,d@U[;6-3U>&WX>/41P1/H\Y-+\NG]=2dQTP@=LJD8E@DLcDEgR[_1Y
>TOOa8+G47\6)MS?[C#+W0_PMeBSD+VR^IeZdS4WDI,5#Db><40>(FOTS(1EP>.X
7Qf?5HEP\cd\U?I@Y_(E:F3.bA5^P6eb-R)DfXce<g)&Q#N3dSE7PZVK)&cX?;>?
:<9W/-2K#AGX]g6ZT(DeQFU;:a65F+[UDYY0SG@K+;]>Wd^9S0W,JE@(/QKg&I,;
?#ZD/J5f9]Y@VQ&@DH#/K;]gO-@L<&I;V[U\7=d23@D=CWbGA7@2O.IH+@6_\Rb6
9#A]bKY_?\XW8X6L;DN/.>UPLd9H_@EEG,7WC1cWW0ATNOH&3(7W0CQMPOCN,=/G
R4N(BHaWS1LMYc9+MZa<M]#U9PU[>L):be&+38JccS,K(5>FK;b)+RJ7A>PQM_8T
Q:(&3cF-W:c;Z)Q5SW3&K0>PYHgH7fa0g,V?J?Z_]0P]5)F99PO)GLH7Z1<ESG?3
A\gfX/,@E;-<X(NJXJ1eGDO=&,eX7LJb_.Hb9F;fL.L9I(3R[KG.H>Og:&:BUSQG
XF9HM[50fL\b,7UeVQeY]8bQLMGI/#Sc(_<L5P65G4KVEW4c-9V-QU@]1LB7SF^g
EbT1ZBHb=5\Gd3Y:N#ECVO5d\XO+7P4>K+YfdQ<2OR@4dMfbGH^=KSZa8g@C)4QJ
#?/BII?f#?ZK,XDA_W^fMTLTbJBVb/8A-a#W>G9M]/C5K+R?=7b;fdf(R5Bd\IA3
&1EBa7YP\Z@2:M:X(T8<(@GMW75Y)UUTfWM9X1H-YW#_LG3QJ;EVaeY\31c/2USE
d;DD.#WV6?C?JP]6T)O#EfPc9]cR,(H]^4+MeU6cB:&P-HRDb@fEA\L>>5.cSG(9
R5)B4-dWR]J&2H0cQT/F>bA(Z(04#5-3GVH?HHA.dL<?C@g+??UE24[KK&^W+]6=
:Y+I_QM[D])g.S)T)@4_;948&2,(4^KBA4ZNV^b0HMQ#&[Y^I&BSEL#d_R9G.(,I
3Y54^O(We83^HDV+&2FD8.cTfNQO&&RK7a1DG6\:([30fY_OV@6RXW#P]6U7<XJ8
NF=>e/QESLa6+I&H4A_U)W\:0a-BFLY(/3[D_).(,ZY(9S/A:+,?CP6gY7=@^W@/
/#eMZDAD1+B&?.KI=MV03c:cf&+L,VX4M.Y@)//TC>:YA+Dbb1?#VB]P]7JRY>N]
]_C[PE^_MQMCW+RD7JZ_WKX-PI=gS4Z&):F#[0=G.\A(,H^E^5K_V/]6XLQ]bJ9:
#O?5J(RG;KfPQA=H?YYD7B/bU&_a/de9bXUTQQ#,E>RaEEF9d=O;EPDXAdSIVK63
f^E1.fN?L.K\GXU@.<_DG)bV1(66&d:B:aNaX]>HI>9Qbf\SV?3^T/6EOc=TED^;
]f^/P3\b)(7SE.7Z.M;9?[ZX)N#DJCMQ)JcW/Re+Ea,e^8N10WgR^GJ6fU_b:X,_
:_1L5[OPU\I6B(7DdE&V-?>KP:gG6Hc2Te?e]8+;TWbJY>.5a\C^CHV+Z-(ZdM=T
7^aMTX>P5V6\;a0feV875(gcD0A;SfJ\C;7D8#OG3?<<c>[<;ALZ?AA=7.>OZ3OL
D]-U7c&/.WQ\2&M/6?a^a+-FF-JW:QP2\B]b./G^Z]bY6,863Q#8S;d7_-ceMaSc
b4K+_]2II9OZ(5,B;&#d,Ib:ON?QPSg[C00SPVDE+\/5WQUD9QS0+\RR\OdAG==,
D59^DR/S_J>YS=WI\ZULHU5#4[V&BD>PeH1G?1(=V[\.1N1Te@(\a5Y[P0L&)cQ,
;(3@3e&[RK?O9@]M?F123PUObR5E39MR1N1?;@K9\,g3L+=-HU5/e+ED(A\gQc_<
(>FR&;af\I\T6R_e)U)HH+La>\2UJAE^]Bg_GM>P;P.4GFNcSB:WGIKJ=O(,ONQ(
FIe3B@-V,f75+BY),A;cBC;7QL4?4U8#A[Xc.G.5+dPd0N0gI8G#=E7PMc0LCR65
Bf,f.]?WfHLD&>N<#]eE&N0;)T1/JD\+78&=4H-:CPS<Lg.X)_B19(8=#^429#N?
L_TZ;Z<LFHS0Me.X<M]10<c9SGd;7>O/:7R;=<L2J)?F1@T^ZVELda0=:L0E?ZUd
ED7?7Q?baETU3B=T+14_#02-)LZ?+^AVR5/YFD1cWM(#IdfY+H>L=X;SRB_E27Qd
L(>2?RS42^6T[<?15[bBOX3:NH@\&4-c)ed2>#S5742VN]PZR8M#_NTH[</HLRM(
G(fcf:(<]HISg:gKWKbM,UV1K3#U5K:EN^EK9V99;6UY;A?^)1H-ORN@+1-AAS=N
<f#B+\+YP7Nf#2HF8O^>Qf(6R?(G/NU,QbES^_P=E.a=P],4=D-:U\^)U2IL<c=1
Ye]\e&f+#_(=LBP-S3@BcETTVJ09;>#F4V>K@L-FO,L@)9\>,L.B#,/aD14QN#5a
\BYYW6F(<f\=1+OOT#g#IJ.4<1XD[2JF5Ma[_3+d_(_e=>92ZVO4_>aN>P#.L[:_
1_5T1N6B8Z9_N<86TefgJ,K4(R\Q?cKHW&^e@7E(F362:2:9[75>^5b@_KA_I6FA
aN7Ya+515]a5OGB?d3VT1eG29098b@R^FOP&Xa>\:B;f#_5:c#P\JB/_CQPM6c,E
^#P@1e.80M)@WSb0:WS@Ee@O_]25Y#VB].&Ee:B<LJb31f9bFXY7abda^&Y6+JC6
+Y5K18D:/>RH+X=(O&gQ1VL@=_4,CgdNK(>Ga6O4)SF1_?@/dRPH]+Pg#0:0[cG:
GFGALOG)1+H(=S9a\\LV)]aLG@^VT[GF72L#=70GPeUE.DOBK@g\+MM)6=bIJ-+N
+I8[914XJ\LW^H?FQKX,N-f>AG\Id6VJ(.+RZL.HL8)f=BI5BM,=[a9/0;0H9?eM
@6X\-OCBLRMGf4_NH2,?MDdWY?CGPK_gWV6H[]<8M2[PG5;?dORaI(W;eR#/2X7=
[Y--4@#G:7^XI(bM^^a(,V/D#NZR:gaeR]HEA;VF8U#.W92R;A>O28IEH3&;U4S@
I-6KQ=g])HCgf+:G\c7(@_<MNSFWY-a\[R=L<XOM8a(TIA.SgDT6,^4)6I7ObMZ+
c9??9_I-&Fb7P?);&T5ZRA7Sa14PdKf)UU/[H,;b+ZXG6?P3^QBOXX3(6\;P8QI^
?,1]5>CU?8?3c?M2,AP.0Q<5:FIKPc:I#A0)ce7P\MZOJE55)9V\6Q>NCI[RV<X&
(\J@SQZe4AR1Q7:2Qba0RB\4<7E^L[-<G[.8LN,<LQD]fBP\)B>B\JQ@^aTDBV]Y
W8HD-V]?6X:bT@RaENaba\X1+/6&F,;QUC=Ud9X.cC93?P)#e/B,V2Je7U(Z5\4.
VSG?CZK40gA_cHAb;;fX82#V27]adNFePXFF0/)1cd>2cKF?cX7A821)NA0MJ56:
<L,:N82<2AJ_LR\b6XaW9;:LGGV>:gV\H3)[gfMV\\+Y+;G]I1M10UdQf:F8Q/FF
ID:b<TX.XLfDHW@8ddf3:ODQ5R@bE=D=R3;1D3Z/d-)D=_R83YYXL_(g:EfHF2KS
DY5/+[\KH-AADFgR4J(3G@471MMfY0ab[<8_JV+<SFT:8gDW6<gRIf:X4/O4b47]
9#0a+N(c+R7Q&4GS-;,S;B#=)6,UEcT:5]Fg=OeU=MVPZcB]#XYRXfWPI0R&6?V-
HGVIK4CI?c(<ZSLATOD^gM=-#L?P-:7<JN#)5WeAK&:0G:#+WI7(7\V34aJ5-@@H
B2K^=,HR^/OBU6L_1SAY:#V1Sd-)=VTIE:T,e7HC=9Wc9F\,d615T>QfLMd?)0EJ
VX]dM^2@L.)R_UEM#XFA@7&<PAU^_.P+:]P[[RX(dRM2A+5GS>2WWTdb4[+#WF:]
X+T#P;U-\),TGHO+Va/bSa4QTC-N2cD4V5UED+-L+ZO\MDcAI5L+)FU9X(1KHYH&
M5O3c\b_aXe(?W,84AT;\8-^G\eHf.#R=/S/S3A6I@e<>+N-]PQ?^1]X\;MGb-NR
#aQ.[TO.O^&S\I\BXcK.Q6U\D:-fP.BaMB+77-M_):YdK22GRgW\1Paf&P]b@TU@
[[\?D;&5L7#BWN^1dH6;?f\@PfA8O7LE<>OdK05_=dZ_?^OHW=[TUX\NI.8[4N)d
L+3^W<>YH1\DO(P(\TZ)]e&>.Ve;TT>N?F/,RWd6FCV\A_[86cQLeAS_5DVfa\?X
9^(a_-?6XT1Y-C(X@7DBM9OEe<fN=ZW=#6+=BdG@MGN:?YQFGD7(3CH)60U:8M_?
KZ7cN,aALc.gARMd3[4ZH:N-WP0TbUa5@,O5T>WdH4cgV03W#(e<M-g1RP,f:W4W
MGBR,OI8#8<.7^IJYdSP;c.He>\He^PaeSV/0\@8F]=;5bN.Y<,JT&TcVI/X,QRV
QdBY>IAGX.8g5;@F21Y4Z:3MH>4N3Jg\71B7ZA)>c5]M7g,fZ-ZSE?1\8d>6-AG0
f.3@Tb4:CB4]YOgW-#V1;5V36&\J72Q=?dZ&YLLT7J#c=;B[([;4-AM#QG:3FKRB
QVK:E&Sd@\IQ=G5SZ^.D)H;F-GJVBSOfTGJH4<ISIF@eW:LEYPT??5G6O4DQfN-F
DU)8B@JeDRVGQ.A7.,J2@Se/eL1E#;),D#PHPHQV:JPJ_#XBVJ\=HgA9WLCCP)?W
^Nd5>8NW1MSPKNGP_9CGG]9BaYO-cWZ9Gf#[/9/3\PM^W&V,GUX(P,TbQQIL55>H
[]T:L\B<:HH[L43,10fIU?_1^VaC[&3#DOKO2gSJ;LKHFMA;F-WT&WVA42B(/@:_
/8.b7cCE63<YL+=[&=@,<(X(O6g]Tf:#(M&IfabD^3(H:[RU?Rb=>:4g0GVL7Nc-
D_Z?G\Q[9B(=6[,:ZAIdBY8Y30Qc^O<BWJ:U<7Gf_Xe+TN:XeMD6X2;9N1CKCF4(
,Q13=cPa#HJFPPEI96VMV99,Q#,Z[aN,<Ae\.O@\[PW43eA=BKJLA\A&XAFfYZb;
GEQ0[NS4^E>>,WF(g&<0=LP83Pcga<\#KJ,,HO>NWUJ_3BFOYN3H;+T;<EIG.L@.
EK80\MC,IZCYKW9\(&<0)J.>?4CL#D.Ka:Q9^TP?1CX=?aKTRDSTV6<Q[\8.VZ0=
_.g4dNK#YL]gO;]c=MM=W)=Cf=,CdV=g^f:]6C-4DHg3ABA3^-KVB7R4.TY^QM(#
/g^f,<Se)fC8)V:5c.Q?eDZ>+5d+Z4RI-O=BgZ?#:?2/)C_@0[,4gJ/S9B^60SY(
PX[2dB7@8ST_OF=O2X]8D_5X>T?_d<0UHD7:OX/+RABFb[MaI\;[),7O-/&O1+:+
T\Q?:HZ1Z^d9FVZf[G9SM;)E7QU(>&JTW#UHJ:;4),d@,YEJXEB<B+:Ef5HAKf#4
,c/Kf^-^&20C_fJ@adM<eWSc]7W61QFKS_a9AKUERF+Mb:Z6X<N2VX9J-^>7EBC1
LOC;fG\cL]gD4#S_>dRW)6SCE,HeNSQ&\.AGg1QZ=/V&[RcA-.NNg60)@047_<WB
RA/KRXOX5g6J]WF+1OeD.0_QZb40&McD-,g4Y37EYCe<?+V6fd<MXH;@+JLU@L[a
gc\+EbU0WZ@[E01V0]6a6<-FY,3MKdc+gE4@C&P.GNVYaQ+,]PH;KP&cM;;&O[^,
8;[3\0-0<\Z].W/f::YB?)(C.<QAVXBOWK8QG:8[L,SE+UJ&3DLd1)N/^14K2:Ac
O_ESf2UG?g(GLC,0g23)I>cSPg<R&gG,-gLMF>TY/Ig=T>62,2^?FN8:c#JdM2Tb
9IF@K0-QR@Z0\g#Lg[/N1=dacGU0)=R+BJ:gR:(4/d^1dD(=d#\JgUaNBOZZH9>H
F?Ff@&^^X00_REQI]=GQdCg+WUMf:LXA)</\;.9X;V8bU(=,T&9[H=9AN[a6)4OM
g8><dc2@0P&gD2;5N\\ATIRJePK2\-@F>5fF)CUF33YY=g2=1OQ]-8d].RaK]?CU
D@G7>(DIAWa[3=K\R1\/d;3GXAXQM>LM]b(SE#.+W<4V78\Z-@N2g.GL(YeG2HFJ
>&^f4X=8L5\7&.GICV&7WK][S;?Z&M;^P6,9ZPL&VX;O=@8L6?GU(f\H3ZPZ=F5)
U6<9Gae/>d3&T)+YL@?G__cgT-^)#gOZOT]>1eO7caaTF=1>8]Z(J_XZDOO2.3bb
/L4ZO71CW]Q>KAfLKTa21TKB_?_9cM8UJ@A-S03aM1GK3^D;DOJ:V?0,&.PK:bGg
[eU;O45^Ab##eMQf)L,bPT^[P;M(&e(IG-a0/-d5aS8(226G,]B@XD::CN0DW0V2
3dWH]S.[03SWW<SW\AG6NKe>Q[d@CQ\UM6\PVP4Od99THgOA6QHE&_K)NdSXMCM1
[9\f/:Fbc)[f<-@D4dZ=Q3@b0#60c&TH<(bJQ=8f8gWPf/gA4>RBX0LDX/YM\/#;
W4U7W(0&IE?CfPMcS\9>&Wb/>=,LK+\U/NK:2+2/Q=>#=J.NaVQQ>-7TKD.D#DJ-
<+Ra/UQe[7M;^I3RU\/dC485A?(12fNR;:41W;X^cD:UJbF+E-VWF.-2a_[+^.Z-
^LVDbg>b,4(6-3MM08?BT8eY>EO,WgDNA=I<F\/)G0:C3b\(Q,eE\5-I>V:)NK#U
(gG8:<I/)@A-&F4#<MeX(W^OgNMAM65aF:P3f[/24;a+M#Sb::gTRZ8WAX&aM>=J
ee4[ePNQFegY)9<IO?HHI0\U1HZ&Vb=5Q3Eeaa^[\77+XE]?0[d<PO-QBGA_A41B
=(bb8,G-PM100HF>-#:<[I;f-570&J.U+QEdWM]#Kg<>=3.\S>Ca,dGOf5?d>K)a
X&:M]<]Sc^g.J=#\&2\CQ?^:A4BKIU-#M47L7AQ=KbEJ06fA98Qg4gO:(S<I]/HQ
(I;N(.NJ(ZW,g;QWgXf=OG[:;.B<).P.7738CfHFfP9Z#HdO(a)K9dgO[5CE]M9Q
O+N@D]U7KK2:Z]N2+\B.QKaJ+5(;;/1J<.]2X(]\J#gbMDa02eKE]6>6:@a>cA&T
-L#]+\bf0=IZ_Q&UK:]=Bd)a>NQBNgKO;M<;:2<=KGAZK&,U,)M_+^)+42G6Y;ZK
9fUYTQFUGb1^KVWO+e<Z.&-9Q.ML)S8YTOeeeYD^..g0911/RQV=I<@ADF^cM=I,
9<9/]I_RX5<9=Fd_<+U/(7XYCcHM]VVcT[E?/66N525+71:^#5(@1=;EPE)88/g4
C?9F;Rg)C)V>>ELW^MOZ+B6@W\#C8R-V;_eK:69F>U/<1<(XEV1M(3;\1[4.cJ91
Dg&eM0>0GSWH]_dJ<P/+LEK]RX9MTW@;WXP(.\M:,2N)E_0_JC(9C#&7Oe6R;De#
SIb>WPgK<fPcIUQ)a9B0&18PKOgfC_L0-SI>HK(B(fSOR/M9b=Z;a]C.KcM@F(A+
;1^2RV74L.g2.]DP#/JDU4._]][ZGH^+D@L18U@\C@b@)bX54Y20]8S\?WFMI[+V
OBC<=Y)T[:eY3[N2gQ<[?]\1Y]g&)O=T@W551d77K#ES1Ye;<GdIJ(9_-6(8E..Z
b4(86975eWP:].E.U&GBB/(c&:eSN[:@<S(.E9>6&3[KUO<ZD8BRL.bIeO)-9V.,
DY=N?ENPWY:-JfU#a:PN3_F2Z+-5XR;f[BaY8fXgbTFZAf3c3LcTQGUS3=0#R[AR
EbOX>XD^^^>COTU/J5Z&?b16,K#Eb>&K^R-Pc+EEa1IFZ26S<Ca40#Ld)01+C]Ba
AP4;bGZ>;KFg<:P;?&adMDeg9]Ea637SU&M[?,,=,6=OVT6E=P(\9X#=ZE_4XA5U
TPFTd,^5IF\9JBb-^ZY@FL3>8AHIHce@I?1CI;\&fTTC^GRELJB)23FPT=gA0=R^
RH]P&I74\]Kf6-&][4cJ+Mbf2V>TZ0\?BUJaIbF3d:=2?4R5.]2S=EF,EAFD7CT[
FOK>-HC(a@7,_8B5:;>1,X)KaXHN3YVafd+#faE2?=D#O,If[Q\R_>HTBbe#;&<@
G8J.X8c\Z\bE=c[MB8_-D/[UaMJL]QW#8)5?=O0H<8HZLZF6=MFP7L/5IK9Y6,S^
=IRADP,R\PR/daF\FV\7=RD9OM9fOZ;aRLSQ(>1FI)+X1;P,.gFa8?Y6<cQKK3EH
Wf/d7aQ\OD[c#K3BZ3#b992?YOHgB1A21Lb(fd7]6+-S1W8CJ(N_KD7UQ2WQR;#&
GTC7-6X:JL6;3_#)I0M=AW?ZNXVUEE#/]Q=5dIa:5.VBD4):N4O\:dc@MAe(TW#4
[U\S+fd:SKBWOT(?J7,Y:_Yc=H:ECIJ\;VVUC+SJ3QX5,TZ&GGPX1I&)+a,7a+EE
D]N<\B3#VgQ_T66VWWGQGH2U975W??+\,M7604,5(Z]FL-ZMRbcWBNL6gMZ:GD[X
fPaHLNBg^eaN\J.Q(^_aU0(L2#R]/3GFSeEDXdIT4^a74?DT8BI&_3b0PXdaXT/0
CQ<QVS&,ceJ788MW/8H2T09<#MEg@Ba0KI1P.A.^-\e3WN/?DAg8<;DI1/6N8@^C
HMM\BXMW?WV0?QgXA((,AQJ/QW665L#<\aSaO90OO;C@^Z1IS3X9YG@0N4LAW-CN
S5<[XLLcZ71?8a9bN;17?84J_;XGSX:.N7C0e:+.fVb_DUVB,2L(LXKUN9J0e\UD
EGM#6WZ91;XY1CgT]_U/CcKD_@=K^TKQ=g6],4PcBY=X4N&@Z80-UJL@eaILC:gW
=XTdd:FG5Y@MJ1O3#^-GM(V,SOb7N].TV8KeR/D>I#:A2>PT-R1ff=8c7S:C2^O&
TD(TNA\X3HM+(5&G/aZ2.HK08@W^]0/RR^LKUYUY1LJQUE7O&DRTQR]8gEAaL-46
--62ZaS/<(.;d0gcdX?3>&:=??GAW?BLcR49RFT?)-[;.ICC89[a+G8UPHZdJTQ/
L-;b@+ca/TcX?IgB[RTZ:V=B\73FN_4=cJ5>F1fB0Q0D4O?8QNVc\(.\9B#Y:eFQ
,,Q1>.7P8HET?IdUVO57\Zb&cQG-&X#+,EF_]7BQD>eTM)+2.,M9e8#E7[<[2bZ,
^&ZDYD4M;A<4[2AF@N=[J-?a,^/9HYGdX5Q4IZJ_#0Eg)K,bc]2.A],4P_WZ48Q7
/;8EDUS0a/GJfFLPf/JC9OSe\bELF\RF?O+gJ#\/V;R]WdNYScYW,6DA:.JFSJV1
?+NF;9AfY&;,dc-HGA9\YbLf?BH_#]Sa=568a?P>JG00CM^6=4^SK((Eg4.d.cU#
0=Z@6a>SEbN_gGLVE1PX-:4/V=Z,V/&<[\bYA#K676SCNIHLOB9V6<=UW]LMR+7?
YA(fS0:CM9<0;ad8B3>dfSO0gFJD@&L=ZdT_J:bVC#Sd<H1ODCFF216.Oe?Dg][f
4a:-c&7fL#R#4VM;D]VMVTb24@_ef&>,Ic56g(E9Md#ARWE2N8J2fc]O+Zg1.0@f
gWA(eb(JKBf),JWN#fXLPECX.DF3:J?6g5Lccf((PW2e^P]V^?8[H^#&.IK6Y.-T
N(,M83K3Rb=]?VVLOYS83(?4]+[6(#E^SYB<UU73-9O.N^6;[4>0?]52F:NLP(UK
P0U,(cSY0HV+4\[2O]bKCG-L0UDA)77gW,a2RagPN&J^O8(ePW2>A=cZKS,)XVY8
aXL_d04DL,_.8@6=d]F_1Vc)W#>(4fFf9GaXF1W)&)HaC1F^&eR0FcgfddcI<g#^
#Z6WG)GHDU]&,[0Z.H##fB8b\:)Ia:TVCP,T?38KDSb\3KYSe,M2TWD-:F4\a,_3
ZU58\b=F-^/ea76-EZ>b0V[(T:@@H>.5GNRGO/&/F1N_8&4EfSd.@7,?XBWKcXEC
9,AO=D2S1>=^/;dLbbVUC4>Z7EYLaH@A)H;O/(Y<FgK@2+7ZBYII)6UE3[).He>.
+BB_eGFcLVJ0&#?,]XP(X>a2A#]]=:#IG0H_&PDBS#)N_IA=_R?/_fO?gN<62=6)
@H0:Ce+-Y_WS4W=)L/JNIM0DO]IA>8-R<HaSPb7g(P,(=eAH_QAb3I91Z8f(;(AT
<8e(3NU<3P?d47IeIMA<+f9:=B+Ib^]N[f6g,Ug8X:NW0c@T/;HHWJX)=]A(,/LE
bO(Y/EI;(19d1?#(fM0H3cQfb8eF)C/-]_]Wa\g4E]TaA+GKDK+I7L4;cGRH1fQ3
,10&T?]/2MX]M<H/,&J_NMJa:DCgR[,8SFbZ<aUFfag>\7^F.JcCcC+37QVN&dC?
\2fdUFcN6OFJE3_GR]]9I34-CN,AAf#?HNY?(g:KY0J&Baf49?M7YUXZH[Ee+\VO
JI?D,F4YHA=J0TYXRVAEH,e;ZTBVJ/d/cg;PJYBHYID^<LEgGCPc7b7c@T5[H6,-
I(>E]eL].2MR<RW_]QPJ3#PB0+0,))EMY4Y,.4Y7G-]^]OW0PBaQgXMe_82P#:HO
60e2SE=@ZUBFbB(,PARDa#+=9gb0cU@2]8&9_7>:M--4&YT-7\D/bLba:ad,0bc3
)Z40C;Q)Q+5@.N#]@1-PAHT9+V_3+<5),6:C<8JML=Q:\S\(15GeY4>&+)0f_LX,
8V]P12f(2gUVA:fR<I#dGTF85\_>XU^?<IXGX\@7N?U3C)VWSJGLYNO]N8]2g7e;
cY]RM@#f#P[D.@3,3]5.WH_46-fCC6A;HE^/1J05JT1e4N4_aAY[BIW:a\Y/ET]H
.=7/Rg>8XL:5KaW:fJ2[V9.];M5EHKT.XDA0g6Jb\H93B0a\97UcI(^E2^LPQX@B
>G7XG7PY4+a15ILW5G@[cUOScdE+&7LV\;T:PH3+75FdY+;_<cF.FQa5_5-=\Cdb
(52\5OD22.EFBDTcO:4X=d7^_KeKU@[Q^Q/77C#_0C_EJRSIPL:ML=D/R,<bR,F2
]]fJ#M4C?X]<UD_E+0e8D=KSRSgG]/=1EfWagR0H@YM:2:#S/bQO9@SHbVJEc,0(
\87D,QEaD[;XTJH0VBQ<^R?WfRC9dd?&R]d/WfYX8OPI8].4DfJ6FS___WbVGFO#
,6K;&S+K&L>bSR(5JB16EG:S5?M1Nf@I9L0&>MQXQHAIJf0B7H.XR@]<:f=e<Y]Z
+Q?:H@7^_OU+6#)7;g>P0R,b6?)785<5T51BMd1=+=09W3@+6LecP6S6/R31Rg_b
UXFHXW/G/Qca;e[TRQ=TOX:S&H+\IO_=0>bCTCR8,-b03E8H2=,7-XYb0S6AE0A\
Yc:T^F)8KWIZ\5bda8:E0@X(9a.\@LA[QO&3EPL9D:/)f@,0d;AC\?DW:VIR\7bH
ZH_CcYc,378Tba[G-WWWF7GWR:QQ#ND<bN.J/0d9O=+Cg-M2d3-EC^\?[D@,X5VV
-YbRLBAgPKge&1OT\dUYUg,?e#gT;GM\+7I+V)4&M?ca813NUaSgC/J4H+=IPDHR
9=G]_I8b_^DUg+U;9^@3FX-F[cTL@1aLL2Z##g2cU7Y#@=MYc,B#CO;#+=>N1dM)
]IH)=R7Z(DR]=T>]QdO^&gVD8JYf6O?JCfC<5W2=K9ae&EHb#,OKJAY]&eCETF6P
@W\e+10BC.4EQ/KDOgQFdG:g2#L6T+cA9E17N_;O.\M##9G\_]ETf+7U&V#<+53Q
dNJae64<aL#2Y.(fe&FK_?d);44g8#EX)(S@CL\-T2NE,LeW7#DR=,O,gM,Qc8Q[
>J1[3V9U\98@(#ZX,b3<Ua(Q:?F1@+3LGX&7c&g?(d7CT>;5eN3,RUVRFR7RM;S[
FbP_&0Z2@:-fN]]ISHNCE9ZDNLLU,CSA4KgP)?07<UR<G+X1;(RJJ1@@XK3>^VQd
BX9V?++8(&^G_Ab_8cg.;?#GN_WBWAI0.FD#SEDENc11;(3)SgC.:UAF@5Ua6.,7
:^R#V,ESgO(97eYd_SNQ@fYH,P348\bQXdg75Z96a>\IPCEK_U,;#Xc1I-d3YQd/
@A4P.,2(-HLX#Fd>e-9b4S5BHY6?O:7RVX6C5G8@_Ga9X4L&,,-C8I_4A:P.-M#R
Z]CW9ceAU[B&V(5)NLCNK_9E6K#>30f]W7HfDb1@g[8X_9[FRWN-b\?4//6D]Sff
4[-^ZJ6#faKXTADD.-F;UR3Q2_.9INJ_F69=BebZ#X@C@6TaKbZOQ@8#.e^5;Adc
PG#abf3g0_&D5fa<9bg3JH\YdLUK5)M/@B,)TUI44N(,V(I[5+e[U??UXF=VSK/9
<E6EFKT2FV\O@9(TC4JSYGW&/:JYb/TVNQZAgQ-_e)YeI/C./a&,H:IOA8.#F6Ue
d_S8Ib8-7>EW9]_3g)W7M\-+P?cMWGC=.fZB2RF\JIAFG7BKMC=[@g[f\^?S@AF9
AVfRHA92.c[Ld.>HXPK+J?53GO(44E3?YH@Re.f;c3SO]dD-V;4+S@ZB@)ZT9X46
,OPG12JB-O0#LJ(a78OL89E.CKZec>L^V2I1-PWdb.cb^>P5Qg(PG3+5]<Rba+S&
THeO>#F7f.DRaO91QO7-^_@J1eIWP6L#VWLJROD@Og;Gc&-[a#^bW2)049S#Ea7/
I>\3Y4f_86a)?0UYBXfIPaHA^Jg/<Z(3[4IQ,6P?>W@^Bb,RS(VO@ICWb,QZ55Ub
3cO+AN0/.-@:E)[A_95<EBeP9&M(A[RR/L4[LAeDfe(>fJYbM+Z/EF\Md7,f?1J3
MT(C9Q<KH:BE6Je4E.VXTf:ZZPPAF,)&XgSa3LH.5#KFf47]+G?_YYa;01f+UY8S
Q,./L,=6^09EDZZXH>(5J58Y,ZRbb@<e;Cd>YO1URC\<-/):Be&V)2Cc_KV0-U&d
cWI](1Cg.6a0KW4\QC;e2TY3UHb2ceea[OK;fIK#Re(A^8?;?;):_5?H@PY((Nb\
;UC]R_F5Xb&2.,MFELI3MQ6\E0G/D^<Z=I?#>2>>M9=CgLJ2Q8.a;<\VKVBB@g=b
Oe\O9\gU:>Q6T3IJ>,^]Ic9VURNB=:_]^A1H7FPX6UYV5MJ;QHbP5UR_8X>6?M3;
L[F4IIWJQS<b6^a=>/Yb6]\<E2D?ccF@bH>WTK\EQ<U2ac61aB=KJ&&#XV53fTFN
ABQ)A9X:bW^=)KDO,/b-gSG/HZZQ@1G?V3UCUNKQF#b4F9;.e9MO)HcNdB+UX[e<
IJc(MQNQeQCQ2X_MXOI)9D>DUGU.86ZY3A1&5L/E>e_A6R_WGIG##G6<@W@2\E5V
[bTDZ<U.a^WE45,Mf<e?3IS&#3WVZQ9AD?4]E(=aWdCP9/8KEf6cga&g1b9&=B@U
.+aG6RT1AZ0Y[.I04GZ@1FC17[35V-Z^,,(&TgfS_Q#XENL^f&MJFZQ79ID1H1M\
a-D>2J<YY:CRK\]Q>,RGHM;5O7dT^,0Z1X@dNR8DfH-^Y5JP&9)+G:fM0<PeIN0(
<WL.SC:3LaY4@f6e2BEbd=JCI(ba]<E=We&ZN+GE-)N69&C6YA=YB.Q)_/;OP6+Y
0GN2Gb_TRg><d71T8d,.H-AXQ.g8eGfd<KRe<:6.E]>C(@IHf^8NbPbMM_[;=[:>
UWf,</_N>9(_<1@URI5&f=GB+TC\)S__:f2X7Q6d^8RPeUIdd2g-\4<K5#S?/L4I
:#CT4I)FIF/W1M@./O]=]U&T1+24>FJR4K<OCX2Y.O).Y;S1+aMg,X_LYa=7d10:
KB(<P\]6BaK3BXAP73I?N.,_XaP6/e?[Ne8PTB1-25_\SXRE4/;bWbB/FJCd[Ud^
]g_ZXF/T.a5_T=baQ=5@4&eHaW7@6GPC7VPABJW1Kd4]T]QR)Q\I=WN@17?3.3&1
Ib3f.8e6PK238V8YR7P(DG?]J,[a.ILL?8H..DWD=02BL?^^[1._MLQO,3PRD;E@
S<QX-cPEca9&AAIbY506R0=O^<,AFc+6AQTU[<4\:eE/C=^[Q@F>,EF0^GgJ0N7#
5Uc@(Y.M,]<AVUO45C&(KD=1b.&dI11@>()FX;)LSB]@O<X3.VFVb7Z\DUU@82KS
U#JMVa\gMZAR\1:PTUINMPa8Y<_,[9c2M@4Ff/++2UU]BdL>f48fVaeKOD-)+f/S
LGf4aQId,W9Y5-\DU[JLg4cTC>9e:HX--4)cQE6?&ORE#0b_PHN<5faE.[G]BcW^
<DEN:090(BH],1:EgOXVP:]E;FEV2A(Ab([V&9HZ7G7M.^_P[Cdc1,6_@7YE]JCA
+Y[0gPOad[UfOHFLIWMe<5<dD&a6<:TM]a&-WT<YMfcPZ:VS#]P<[/^&HXa>U]9E
e:,/6Q;S=,ESbF\2THVJ4-IJB6TD72&5d#FJ=G.f>?42Q@5;1fOTg327T1a[K9NR
)F-.#&>F3U5S7^2_CPKAIE1_cNSAV^D[)2)e?KWTHZ@<D3>FNMH/B2Q\bD7bR0Za
TA+]P_FN2O,JB&8_RJMaL3PM8/Y).K1PA)R&;/b/#J;0-0GBF>YRO.eEN<:&;2A2
SGQ<30g?>04BISKO0XR^N@:[dL4LAB-N;DKJ#fUC[JWA<77_T=<0]06S;Y.Lb[XN
86.4O5(L,ENA2,Kd;3ME2fW?aTP7BWO?D@]+30BeGH+1g1cCE56B8V.R&L\AOIdY
6V(LAUb1A0=II(H+\DTg2-Db8MT.0:##bL/Z:6&W;XU75+D[NN8KH.N9BcJK<R_G
ZT(53SUHECQ8AR/(;fZ)IVQ8]T<^_((IM/Q2;VYdB^;A3U_(g;\KBPggE_EA]Sa(
QeQ+Og1_#7?aFWC01^H=OR6<=A8@DL:_E5,:S+,abRVf74<_W9;3H[Z5#8_TG4AD
F(F;M_LTZa(Xa?Id;:b0W5;AVI?]2<FVS:CZg8?2(X&?S[JQ.<+V7/.W)RP/+,PZ
E]/9eC\?#I=^)5/:+\B5E?=c+M9c+U\gc9Y\_PCC]HL+MBfV?2)UQ127BI))\d[;
27;KFf4bX+#+daI-b04E9?8VI33LIPK#\];;.GKY#WNUW;d,[R=WXJW,U6b?>MX\
)M;YWe38c/9N7WdV78\I;(/RQ[TdLV)XNAV\d\S,;e\Z/45NL)Q6a0#FU?N,7I]Z
DaOEI&=Q3:)c5O_2^UZ<WR;(6bVM3&;:E<c<3.7:H7Da(B8>N#b)YaH01bB2&)/C
gPJ&S,9gf8MDJBfN60EIHaS?_>>gfa<d1H-RbVI9\L.\YS0FRO_dI(K/Td;/)e4T
8He4ZXfK;L[<@_/1W[BT4BS:O_[cS&V^N:.dVA;gA1X,)<AQbb-)JaH9b#03N@4[
IQ3)9,>7dI,H^L,@@M103X<QX7?7J?a^GREJCMJO)H_0@O/>ILX9]e^.AebXMSW.
R4GJMU;<F656IRO[ZKf4gJ3[Q]:/L)ZN/a.ROHO0T.YN&OfYDZ4VdQ?HdR-OJgBF
E+C1\L@[bI91BcHE6J_D5EHPDS/G9#DOI>AO8aa2ZC<]<5J]KMV8E[dQ3;?&PRg]
CCBDC0WAT9Md30QM^Pbf]=(&Q9Z6IfU#SD:_7(f^Rb?dFB#cU:=EIG<e[0e(8gM^
7SVA,9KNf@@<3F+,5IALG((bWWN[)N)Z=B:8FRKP>FG?Lf/;^:B-ANZ/R6JN8C;L
)5=-]WVPA(:6,Gd#@K=37]bgV<(#P=M&+E+)7]_26E-:2a0CNUd_O+IcVC_^ZQQX
:(GDV8a\P:YOaFaKafYf,Q:^@KU40_1YYIdaPG__EFF?>/:#K<bD>#PEcJU:)I=4
?1aa#4LYP]/4SC062,3/=f0O.I_#PaLDG1fZZ19._ge^_bT9HEa+eTdD(_<0G_T?
DaGHb+CaI_&A.e;g-05K:H(IfI<AMf&e=bPMcbgP..d4^A_[XKSXTd382&>:ZbCI
NUM+96cQNg_/?Q67(\RVTg]>5@EMPa-NAae99NM/+12,7L,,^&)@V^.bXN7IRKU1
_MB)1.WaSQ#O-#DR-6(ULU\Q[1#4./#_3c)X4R4g8B5W58:QZ]+9OND8AgV4;#aZ
_J>PaW4>eG6@Nc60I8UF<K^&:72/M)PK@.T=(XCb7OXOBGadAO:^1YCJU6NVaL>)
bF(OM-gg01W[@cQUbFScQRIYOCLXJ.1cA.]J#Q,W@W[gM)))T#dO_,AA+Vaf7-ad
;GG>Z_(-R_R;R[^+U7RHQDCEACg.G?YcNZ;[W>:-?#IPb&)KI>N0VLOTU,QW6X.#
T8bI8TO5a#S=)DWeFB?/7VL7-8:B)O(Ca;aML/VfV.D+E.DC)RNHa6A>f)]#?2//
^U_SPG7e@V1,)LTQVZ[=&;dB]ZJF2IUHX7ZcY5DUSY0Y2A(]73<=WM+-8=bXG+\3
C7e53A+9E;S1MSHf[FZ#cH:W.QJ#,+\94#E+C#TF=-4^9eBVYRQeE9#)ZgA=MGg(
_EHS(;=WS65VFM(OCS1O-P/;LK#6CTM)/K;SdJbA9bN)0bI9eUBY>RFE-+-dBY=U
d2c\fPO/R;:0M7_RW[3/^?1[J9/9F7g^3Y,N)<K:Fa4?;RZ(0Fd^c<MJ6f5T9a1[
;;ZaeAc321Z1LZQ+EfD;ADR0C7EL#)YD26Z74#Ud(\T/CK_X>d?AV#,:@7ZJ6E^-
Gc3-#Q8+XY[Va&X9,GJ_),W169GcAFL71=PFX<,3Q#&d^cgU)-0]JJ3)Z.<D)2V@
DH^G5R=N.1]^L6EGJ7?0XZ(7NWJSF;[N+F64;e&7WL@ggD[RD[>QdbBE2c^((PeD
/=^F58W4D[a/DUI6B,2;P6gS8NJS;,U,KZ=+CbV[\H1-+Y;H\-55(QIXN,ZNJ:T3
,3ZHMG_dNQ),f1<2_,9Oe]4ObUbGGZ1KP86eX?TPO0TeAP3bO@MI.D^<W[dW[]c1
63b6=Z&d\YD\^GG1Q+MIT.XGR]=F-VBe/<6g.7dVV7+P]f:H7B?DfRdBHRN&UO[=
MS[dP5Lc9L+_[:=9Sf@/II>05cdT[0c6/DGX&=AL_=QFDBVcEBHT^LGRG\Bc3=9(
KgJH,1/OO550>3X)3KdK\cd&HN()M:baSV@[I,IKLN9=U)LTEGWGbN/^VL70O[40
H95bX&Ca3/C,4=<a)3f+,WC6::6UJB/(,]XGO@dATd#QK0#].W\2YFLQ/F2/^7g_
7_Kdd12GB<J2)7a3LF#R3MWeJ--ZAd4E50)-&=/aN:L/3,1SU&f4UHM^-eHE8-[&
MT0DG^WQ_2+/g.=PfJ2#ASU;.ETZM+2X1^=HYY#)SM?<DPe7gAaTUfFO8A._V01D
QX1dIJH#AI_XQ?eWB]O&c#-cI(TMOPXA:)-UBFR\&0NM)S]X20cA&3>2.?BG(f-/
,C<8AR0[GZAPd;@MGOM?aLN5&V&2C0>5I55#TM>[Y,-<eI<U@KE_UJ>2KSG/;G7.
VPYcF+ILF<XA6I+K0P6@Y^]J;F)CW?W]K0.bD+-d++,GZD1TSR5.)HcL?TB.NLeW
/#_1SH;\g9Tf?aUA6Qe:CA.?@^>#-LHP@TV3U?9TD-WVdf:F-QO4GF-:6:2+/75d
-_#PT.\VD,>c-KJ4Vf:VQ<b4=fe,9Abg3;d5d+If5a^+7L0F]93#c43FI]SPIgPK
,(6Q:g>@>Q4ZI<)O.G#+&MGZYI)c>e1_WU^:>8fXG9#<L_((J9BKTaEH[AT2e<L6
#0gabd>9KZ3)MBMb3\#V/+C&RI9Ee9GICb&2.<(GZ#35-#.KW^I?R;XUX75d_KM:
ADCg)\#EQF4gN(Ed^-G?[4A780@GL+;2]N9A3.N4Y[J;=P<:HMb3PgC2a?g_D^fO
IA0]Z,.Ge3=dH?U(HQJHE68795\D12/b:IP1U,H<IQfGe:+[Q(/<Wg<]8U>0C[ZY
E3eHNS;=gHY0<cA)<16^RJ]TCZJT@E]GB-]NZ_Lgdg-H)CW_^\+6+6D0.f[#^fUR
\53VHH]5b&fV[T2G\dE&eK4bR9BaIP/4IZ2,DC?&/AV4S:)W[>EObM^JQSQJVF6[
3A-fG>dCESLYV?-.5MD=+2EREg==d>5:]1(M4_P>fXc\>O[,/,UG2II\J=9,WLB<
^70I[fBBa.=c<RKV+7HeP4T1@Oc@T9&CQgP@XH9AS9WN:##=J0RB.]>#0L:U,7;4
RH0(0&1?7,ea@EO<^I2;YcgZDZ\;O2<7I^f;K#7Cg<TBWY<Ue:\:a[+cC=_OS_PC
HVXBP>LKR5CVg]V+V\b7;G?1LeQ0[H<S]UcIT[1<P&0#WP&ZLEZW)UT5I#/W3f2Q
Q;;6;C.CSH1IMKH)HLMf27?YUZEQ@BHf@$
`endprotected

             `protected
UUbV=U.OKOO>6K67_+-9V;1dLP1@FO0KP0GbMN?f^\049g+Ug3+(+)/FLa2KW3ET
be?SXf3+OMA0R_]CKPL90.6&MO>d9&(_>HfV#8aacM6^D/gNbf#=ET/E&ZC7d8P>
0c2Q4XZ&+)b00$
`endprotected

             //vcs_vip_protect
             `protected
XTFK5L#_LZ_ESbBZ(a7I+d-BV0AgS@+-8^e8O@/T&,@+4>FNWSUH1(PT?,HaCLDf
#E/[Z/OL__#?DTL:+E)g?>^MC3UI=-/^/=/5@YC5H>&FW(R^-B.?RGXG+PaZOWR8
a&c0I/e\#[;C_>M@2KbW@4?GL?(BDAFI24W5f]BO2A2C7=0Q[OIC)-MQ:C>G?]],
/A8WB_Q@21U.<=1B3[6#e=A7-Z4F8[1N)?KLN1:EeY-?8AU7Ld70.@DgXGK3K+gR
X3AbIPN+8G3O1^7-X37@;.X2J=Z-g(\(-c-UD/.W]3/a9WBf(I1A&7[,PW4DD?S;
.6NYY3QS2J#aGBCK8A#c8f\>&M^Cg:1]+WPC@^GG6MNd+Ne:f2[:)2.YNEb@[N/e
(2L]O5-?;TWM@3E+M\00+1LcID^7d(R08I0Y/G1P[1f-N&1+3O>#/@)H>5\])Z@H
IL6^L)_c:ObM;W-=1RBX_VZ?2182-IH/=>W;O?_ZE=]3]I21ab?LIT7<5,:L?X?^
U\\__0Yd)<JI1AFcYfeCYba/[2_-aN=CFN?R(dQ+bU6Re^3U1T[HL[VgE(8c6dGT
0f[9O>1=H6MC_61O<;X6eeF3Z+BT@UAZT#]N.V;B)_b=_<_;\:/1LReK0J..GO47
7(F)5CDSb1(-FSTA2[\1_XX6Q6I45.+S1&9c6]/2QI4,+J;D:XNVWWVfCCf0de[8
geR(@e)d47F:GZFbH+OX6._D;f:aXf>HM/FCY1\]X3gAg121Q:_;GJSe9(V;eAAU
&RZIfD9>&CWU.VGDJDf20L#V,HTV&3WWb5BU^KeH@X8050#b==dT<R211@a603]K
Dg9@Q^,HSMQF2;XX:E_M#5PG=-;3??YL>V==FE9U^dO&:&O2J^;?eKDUDJA(_:I:
YJE34UQc-520L-Y.);c@;RNeCV[JT,9gb:Lc@:T-DK/9e-S248V,&@TO0N5CW)#J
.-:52MKE/_;)FRK2#Q]HLe8O;@dBSI@^#99-3Eg_6#NgEb?KZD<&5F-?2@g2L/T=
Q1b=:=5^N+Z,C+2fZ]fC<N5.&c#Y;9555A0c5-QUY4ScQcP-?/[+SX(.g0,0eEe[
.O,=:cXCgR?c]S2&)Tg2.&Zc:Fd9WdVDQHJV5W93+_RSO-5++;&&F>,0HZ4aa5>(
Z#VSGcT_CO,/K?.7aW4E#:,^C-3b2gLdKO32]S7b7VE-Vb2#6SfW2.RY^;SH-75I
fSV>AKG&DM6+TI5&WM621Ea90VSV2;<2QD:W7/gU[NI=(_#Y[Y)^]NDe^e5LceD;
=L3Y^6(=#<MB?5.f_g\dd?0WKYI<fD3&2)7LN^;#@Vfcg?/eeNf[?)/6-GXSY:\S
#<A>gP7>&f&KdXKF\dYXB#R2]S)\64QB--6W=aC^I6RV;ZGXA&LZ&,ba[U=b+U.5
^LEd05;7LA>/Tb@(CZ&0GBAQ1.GYOH^I08Z<8FFe&O4a0H?8e_F43)U\OEPE@&c1
>QTUEI;(B>&Bd6+_B=.4DS:8V@U\_]HB64FM+)O8Ia+HF>[2\aP]@9;NgfH(E]I/
_)5=aW+d8[aCV[b?9O:]11e4@26AWcJTgSGXK;??14<D_#/GTF/CHf>gc[5P6-.4
#K\N<VHQSDVRY]45UECBW)WbE3/g.5/S\0Y:KS1\EU0^[CDf)eLYWg\]8VaE&H\=
6;UfeF)6S[H/Z1BF3Ve/[_F5=@G(WYe3V]LY<YXY8g=Jfa0AD5)36d_87+V<@ORb
fQIC89RY9c]G?OUB_+Xgb>Z[aA8U[]J-:/HWH/=7WL9-MFe+9E6Ue]8@BL<]fLKS
GSFg(aKBCP?,-1bY;(=J^IdNVC;6GUdX9/.gP=G>5G,d;KIbEb]U0><21TV_+egL
DeWNH[7-TU[=&71Jc=/3[?@?_]+NA[<PPd^/,##a<d^+ZX5;]:JB-#?E&]Z;1UMI
H;(5,3RAO,K3]G05QSgbJELQ?+bVeD8?cUgZ1ff-9.edP@V<[-^HBR.,faKe;\9:
W]#>2I(:UHL6]48(9e]0fNU,P6&0>6B,#UHPFY]1BM8HI1S&5Z?#PKO):KTY.ZF?
c?P)[c8[MebJ2>G>F3Z1K];MUd<P39:M)NbOaW5bLX8-4c:SC(Y-M2WZ#(W6GX)D
3QF?dT[.^)]/1<B8X;&@;V\17.fNbV7B1PU84bJ1.:\KF[f[#(Ef-f5IWV+1NPg+
5PSMSTg2dZOcL;c_\@EOY[Y33UTCR,K1L?^dda.-#@>XJBE-U&B+YC./4a,2TIGT
db-.e&9@AD2[_QP]+/?FVg.U@^5?[Q2;eZOQF=gfLa8MM92E7#7)]W9<-UN.Y4#<
B[7QF,M6TAeEdee\<^<V?8L608_5I,ABb4QaD.71CZ0)K^U9:[7PDOWK_F&>R5/\
gDH<_U^IFS^I&:N7Ee,]U/YU,K?N1><5U3OTI/f2XK@1Fg&G.?I&3OgF9)C8gP<[
9?gUA_C^FNVO[8O^><W+B]?CDfUV,_M@AbDQS5DA6]Ag&.::N[-C:9G:)gOSCY<.
=c@:JCaMgeDYBZX0f=Y@BDR3Z.DYO1[&62B.d3/0)b+c+^00aaKS6If9N+7]#06a
HXC-[fbe9HRaKR8G[8Z(/_=B_1L75>8KS6#S>9NPR9:)98Y^V<845-1:ABbc0Q\\
92@W<M8aFDVN=C=.8JCR].B=F&(&W<H\1+W,G5A;?AT])\]KOR2G_N6SM^9XDXPN
2.Y\L6f1;a;KLS<D]YB7>V1)B;_Ze:G,Y9.?38O&RN:f2X[Q3ER^e]6a9:Z(6Lb:
7Z&-F\e9LTX\03XF=W429I#5G(:D-MNUSg+LG,)C>11,f&8.>L/QV=78/;)(Q8TB
A@Y,2LO^Pf<3F<U0G\K=<_TeHLLMH=HQDUJZ+eeGPdQW=g;DH3EVRIO(gL/C0-Ce
KDO7]+OL@N?H_-XXRLW:Z5S+J/]HA3e82ND(=;F)2M0d31;?7AFI@Q8L&/dFDV;V
SIKC1TU?&OGL/J(#4b9M;6D-6]G>JC82-W[42J;Z6L>(XU_T)>(ZL<J+SR544Y>D
V6a8<9\KB>&gDM/^EABXV:9L]#DZ@7]]-S8g0.>8O-0b=5S4\3Z,.V#+?3JQa@;V
0V9@SACJ+)P[J8=fK-7f#2/#-W2f7,=@BI<?9NBF/U/\+,OH4;HPbV2)13?X?O7Z
d#d.Z\cBH\/GXYOC5R8G(MS=[]-cE\]0(#ZSc#UWfB8:OScWGA[JaN0WS=HN5TL]
:=;#SAFT^I[&L56MG:706=VD8=-I7W,G_]2f+G7#6LHP&H/&T3.J=+DO_D=b.:e\
@+??K@(4,/L6#eY^[1)f3U;aCZ#4_Pf><>)B3=E+T[CLERf=8K341dO-G8)b]#[B
^F;S8O/(24SG=XMQSNZV[.fbCI#Wc=CX8dPd[EbgHNBKKM9).S:Dd8K-0XLLCG02
\K^bHNDDLB2X3WTfKZ]N50XWFH>YL::UX5X:.b<18IIY8\DIY+:-/&#,IZ:9R&9X
Ed]7gTc722E8-IEVQJe^J?\>+J/VbWQeYPY2@J1)Q>:+S3S74\0_U1)T8:VE/[YB
c4GUGNedQ3+./UN^P:TBCL3Zca_@>A:A,:PH.QYRS0,baL0)GWDJ&C2./Pe&ge;(
7U781I7\Ea^Z&fH+A<J\_ME2RVKNIABAQA[I+]KZ17^<.ND(g1AO<:=PU()-B9N3
J/8c&=Nec\)NVL.b_eD8FH2<EV/6I86,[?gg[<0Kf5[:ED+B280D+=VeNPb9Fd&f
3Ha&O(777&16LE]/C+Q,gb(FE7F>Q4\_?)JC>de-cOBYO-fCZGO8?XRA.g6_;=+T
e<d&(S?P3(Z>US@g7Xbg3&8^0T0AN?,\XW]FYCCb3)8_>#0T9dPX15HU(QgB1BN2
V2L9@/.:ME.A9S<9DFOBU@g3T3@)>=<-.fcA3@^,Z0;/_T=.Y0QD30A1#I?H5+CC
#(QABO6M3Je;aFeX#PT\QIB)JPFGQ]:KUACPZGg8dO>cS=efACN5:4RXJ.:4+3Z0
-3?3<cX_X7=bHTEaK5:TO7&/OC/8>J+e:OFeT-#Y-@0U?TNC&PW,ga[P]Q3?;=0/
.fK0SaC,Oa9(8OcDe3JWG&5gRN?;e>P<4dBXA[:Z;&S/b0HY>DA@c@gJ8XK[;dA#
dHIO<VZHJ3&WK63INgVY6.+((+>5E5ffIY/<K<6RF9?9I1bA+>>Ka8]\^?SHK@KJ
#bD7gE@e>FdW;-</5K\9-<bOW]+[SDe09[a?+4T95VHDb;#^,D<Q;e_8aNI^d:N@
d@gdQ[S]F;#9/U6_[-LX__]7X>=;+GOX?SDUeR&Q3>#b:)YE)QZdeBb_[3<a5/P<
&.Ta2.>,C6E9P(5;bL\Q.7=I_9^:<3EMSSJ?))UR34JOGT,f[2Z.<+OA.eV;a^5>
HCA#._>_#:\)W+LQAI?d@):882?^ZI)[P#T()VW]2A>2[<_Q2DV?g+X(b8@XSN+1
ATRGQA8?ENc=6U0FgS6B-&D2#U=f(Q?[ZYXG58K5Cg1UVBQ6LSP+UdYf9.1N(_Ed
G(0[,B@g@-/SYFeb\XW/JOY11AWL7[9@+LP#RSPDYO=M-TA@+2cC97UK8b^L;O_)
D8J#FF1LKHW4.:D^T];)Q8QbOM5L?:R50I\PJa^99O;d3REU)CLB=cdcT72PTeE]
D3FM;7SD?1@cI@39fDY#78/1(W_0RNS.IOZ6T+P7B4JZC^a:7M><CICDf2P20aA^
#:aHDIS.ggT4(MK6H<TK[X_+8Y<\<4T>U]e;#.>2.NT+g8/.=AEGX=;a;U>H)FPK
2NT]TO0N6Q-YY2NEBSU-:^JX4GS#62#D6CDK(EP.@HX:_:1AUdIEP7_@RM22HG?,
1<V1?T3QbU0&>3VX/YP\&9^4=B8S@gQMR)4B81L3\<R_.Y)_T.>Y_?J.2b#@LaNT
f4+2_T,3E[Q3S+3R^M@3?=ac;+b7R^Qb/RI.;W]1AN#c=.IFQ@SaU/d]K.D7LX54
?NT^8J2f?,+S94\c,Z#6T^#;cg\?IY#-SA6E#+@2JT8@BJ)QPK/EDL7S9JY[MID+
:&NFGC5JP60C4Za6B=d.Q?]g9(>:-FXJ>+(8;17b057>Z(Y@<K]AR(_YKgRW9:N]
K?1\a6O[[UA#Q6NM04eD.&e47FG1[DfgBW<67P&MBU:9L7&TD3gBZaD_7@R\@bG#
7DEb<9Q>HK?GbJ>==X\8^/7V)JW=,,CMe:U()<fRL4O+[FKD9I5U8g.gG1eb=_G5
YRW0XY_ALQ:KUK#?7>2O_L6>/S:M&KY_2CI8#3&T<A59A;N9GWNZJ<BH<&MG0)B_
.AB_(_@P_8NHUBc6XfS<e/DT^^]EG_43=_>;^F3S0:EZ;OD7caGI^BJ?8=_P>J6?
\e_4,W6(;9T:O0\]PPc_?S[cQXa:-=7dfg[Q@P2WbVGL8\ebJdSW4d?N?I,9UKY2
&c^RT#[J[#HdAX<3T.eB_A[d;EUbL#6UW-L)>66Q8AHZYD>W[KTN>A^A(HKF#5Q3
X@eP;FI9:]FJ_GZQ[,.1BUOS;e]QFgAXPT)U(1BdIaAQ,WOY-<<.eNL_\WQ>^4]F
#Q]XG\-cWB0/(A,>7:A6)]=(XUZ4FL6?>C0?N]AEZYMK.+E\WO#UdS:[0]&.)5[Y
G>\(M^?T[K>C;e=J_d/XS.N.MVU)6RO4e];.<5>/LU;Lf0IGf;N6Ib.#[bg5VX19
K?_N;H^]TG&\>[DdWV3_)(3Z6:O,N)(_-W-/aK(L4L.3\THW/JGOb]:dCVd^fQRB
bU>f(K-T?M7Y)?PB#.EdeIT^A#T=+NdJ<(Y#W^IV(00C=\AgLf@)<0/<ZbN5F08e
PJd.H/-NG;DDT?O\Gad6fVUfGQM9C3gVZCfP<-\IF398fbLRc?Vbc83\]bDC#eVb
2TO^#(LES&2G,\8YA]aZ9]8LOSdPcE,-,:cF1Z53NILYZ=ALBXS5,]3fPHW,9GR1
\ce<<4BPV2SPE2IMV42V;E&5VA]Sg\_Q[b@_FG>)-WA2>R130aK7b1HK?B8GHe&F
:(<3<DFO]SW5UdHL_<+NY=,a4_O3(F\U3aVIR0;\O\bTebU/]G4_UcOC^eIK2X66
M;.Tcea:XbF;6aTGg4IY4X>9e@4&eVNC4_JW?77)WURV-5+A-)(P8g<Y<]AbV78-
,NP-Gc.4HLYc:>;-B=#=NSWd<XO+;L@Z/:KVFaMK#=cB(,1N&^_KTNXfN0Vb4N@^
M>=/C?,@8_EG2+GGgf8-P8aB]fCf?Q=;]SRS;?7--[:,TAfD105H#(?6,42TXSY:
S>P=5(H7d:\(Bf13A]UR:^E,3H-R<.a0fQFUF(RCcLSDFAI(#MY#J?c,>X;C:C]E
WWJba7cfH<=VP,X=7&C#:2=5/_327M..6X&0<Q4O=A;/^g\H/>FBbV@F(#)d3LC\
/O[87d(85c>0VP-Y757@cAH?Kb9[2O/(QHg)V43ODB93.:f;L.9ATCaX(9L8[.gT
)V58@L5=ZOA3_e#8&P3DJOYMX?WI(aL[W<b#DBYTXg>12g4fYYcM1He6c2PZ@)D7
CK&E+QRbfVWeb)AR@fHJfbAI?14PbbNOKB6SYT8V:LAQ>/>P1dH[FE(B]WBF[?UI
=a1J^O:C+ZU+1EK/f-ETgI?dd)3:g8YKb_USKDR9d^LBcICg,)<aXA2DcRaA^GO4
E7e5Qb^9KGA,DR_]GBEZCf@g[\-<e+IE^c_:SF92L:T_BJ5->Tc;#;_KN64+bAEB
W=;=4VUFY.VW3([O9M[\E]67A+8VHKH/A;13UY9:g1M(dTL&N@5ZCVRCS^?bO,EB
R+?6A18D:_E?)+LH5BYWAIfJU\&TVf2UCIJN.bZad/T[8SY_3TU_A@U_fDUY]IT<
0S)_1W]WI):,?FFbLC1V-4Id[G2dC,CQdL5dcADGL11#+8/YBcGFI=Q+(.aPT>/,
U\,1#RO\^G9;AAE2F[VX9[@-#7d420&YA9T#ZUK,LgQ3Z4&BZc3cJUP,.MVGUZ#1
8R:_f]XY03f9SYE+gV&W<?63#.Rd.6:_H>(AXB_ZEX&&V8<@Y3S<0JUK>\12e>Sd
W-B3]TI[5MQ.L8dK9DgT96:F_2D9N)4_3HY[.C<UFW_#:#4/68bKb+KQWWc/MfdM
-[0+O4@,+gWgRS.MX6C\Ibc]Fg^B+g,5e_EHcV@G;A<MG:5b46>@,9UZFfgUQZ@d
7/CYIU56GN.C+U8;<#.1]T3V\<<T+?_28XMF^Q/^Fc-@GQ&NPXdZDL>/<B)^[Y[W
^AbaAg><KbI<=AdFU.I7cSZ&4cVcT8ST.OVbb<^,Q7X[?UaU>H[&Z?HACdH.VJ.Y
Y8L8A=V&?N:1IHQY7-R=\.3>KH#]T&U;4=(<;]L-8+@a.#^,Yb=?F(=FVJS2]01?
YYPPDaN(>S?P[dS<Lc]IN=@E(SEbEFA3DdMOa5I.QD0>7W+T.Ga=CK\70FW=A^2A
>E<VN#=\+OcE/\I\A)f9f)3>F)F]_TO-K?_-+0RY+#c>3(,B@:VC@I<D1gPTN<be
VFI-P13S=e5G2F0IL8&1Hd,.c+3M/S(eVe7O0e=MdOEF.b/Y(E72;?>eQEgAFM:Q
HBMPK:)DY4&0#5J;Cf8)Tb0>@#XK==7NgV8=:?\Z,::V5bW8.6:M35c_U#\OHD,0
c3L\L>O]Xd1EY(RWS_ZXAFT/7Z:1R-?FGe.\O-R&451P[@@a;6B2_6DRX7G/I8_N
VY5g;D0FG>7[)L3I1<BN?Vd)aZ;]+=OG5EZ&W]#;U=@S^>OU>)9N1Me\>Ag:?\6C
HPcE(699D1-T0B@U?TAYO_)@T9)0Dd?-R&S(^S,)D>QS[HC5C)g]H5g;+/8e/7Xc
3;b2,c4c.FD-EV,ab7gD\^KP<[KP\HB<R7bPY>G5XScHPgF-fR5Mg(g80gKYSbL3
BFgeXUST]4[.;AI1S@4E]#-ET:cX<&e9O&5gQ(8:db5R,^=d&+&Z^Tb#-G81IG(W
P93cA#6WJ:RfYPbUP04.2JNI/0W8@EW3N-PX\La]E5G6HU@-ZKQILSeX/)=R3CHU
^ZS0L<]CX=YcReINY^YZ4S#M/T?5UGB/DdaN[\\#5=Z@b5b)P[.W=M70J9Ja(6)W
:FFX4@@QWKB_\].;<Aa^C#3H(9d).\?78c3)P_)N[K<,6/J]VPZa]E]3f?G[<SSJ
<UZR0QJ3cIP#[78N7]Be,>[WQGNR_4<Xf>E4P#IAA=8R4?_bV+94,R72/W5@:Y^f
9.6FV+BS?AK?(c+WgbE&SdFg-g8f;T^V;;IK8HMC_XB^]+b-eBC++U\QEc4LZMKO
1#]7,faUNg2R1LV3;H9C?b3DaG8Y5UKRGJ(@RZ.KAMGPQ2D#;/MJgS91>JedbBMZ
+OEVAH#C&HL?E^f,gXSWg6JUXb=I.7.aFQBC^.@F#cW/)Z2836VIc;]GAI6HRG0)
A[S9[]/@,H?2aC@/<@&X0N(>,F47.MBT)P3@9QX-J8O;NC\WYZJGgcAa#S??_AbZ
LXGDN@LZb2MN^V,GKU+DS_RS<)B70T44F]P@aY(cU29/>Df4Z<.CD14IIO82CGG;
ZLgX\)UKg<.ePMQF+:Y=d1]1eOIKC^f8:3;<QA#_RFBJaW,E3RW;TcLNC=a-X&>?
be0U1Wab8g7dAgQ]QP8]&J>d3g)0G_g<-(6F4gdTY@F?#gA,@9eVQ3T,OOL&]H7X
V]3I[PHW7K/O(=6(Je-KFLUK9=a_[/(K3/ZC98HGHJI#5):N.f<ggFg^b(2@.a&a
3(HB(CVC8Q+\P[T<QZ(8N7@7eYbeaR=42EL,[:RAC&<^dbBPBFUa_XM8bd4#^HR_
1a0TFCW1J3-?W<8,2cSKf<-^2([#,RG;Y4\JZ:cWD9Q_BTO,K(_7Z]M)=U>FEN4-
7))Ua)_<U4TPC)U:R<_Y2C(2T>J):-26&MW-Y@QNO&9<(_@]6Ub=eB>8Dg<KQagA
:BO1;N7/gUcW/XU12NgV]1\VfTD@0TR+(6M)XY,C^P/^L83KQTUMIMdLBAU3B1E<
0>Y#B.5daZa?X\JW,+GG:^\6>:/YH[/;L7;_9KVbgB_[2aHaGba>eK]P[HN-J-_Q
C_2WDV3R7706=2[5/21_e.#-+C0OM>#@,+&C9PfK]LA:F]E?6R-=d3DJ;d#VQ.(U
gL]<6&^#f]5_fV]SOBIZ)9X(g5,LER#X-,aV3ZTcf9ZEfU9IbUKRG]]8I_AMCPaH
P&b]V0_ZJ7N)YK]1QJAfRTDN&6fZ)XfOEL7XGC+U]=X44<44bL0&^#OfQ.,>dG0]
87=UW_7d;:5[R5dGeQ,[F+\X-8f>-EI:6(;IX?/Pa(3]O\^NdP>+N/\@^I083YH,
:^N1/?#a\G8f]=HAW_4GQ;0EI\?18O9RN.AZ0KXO@06BX+F&e0NTN6.QF;V^#@eX
eTfWTFYG,=6.DG-5I(2Ac,&eBRgNS5Z3Z)3R;,3RI#6C0BNBG=RXDOEdE_a>(NG-
JKYF]BaGK29>&A=ZN49C=J6agOHVdT\GW7^<9PH.3<\OOeKEFA&@4a]e&,++3X=9
X\>\IegfR??LIP@XPa)OBRF)Cd@:eBP^>+5B;L#AV>WR(G6Q?59.8^bV>V3XF#;=
.+Z=)ef@Z]QAg1DHU(?X#^_cX\LcAd,^EG7T+5fTL[V&X;/cA,019=A;TO:dOJg(
0f[e8[8g-6N^cOW];cH7/E&O,?T2e49/HbK9CY:5VFKIeL@(MXRC+5LW2a5.(H5b
I47LgdJ+(8<LeFe-.]_O[eNGJ1XA)/b5K&L&RbR=KYH>2BL0EC@2&dP_a3Yd?,fO
e\]OI#[PZ-c0AR/&Q+\?+3;Eb3-^gTS/>^^b6H&(&]QUVcS&H(DV>4L#N[0+):FV
&dH.g]+[WSLYE)]N84Of1V77RS/eGPV^f;HFMbc_^gN^/Y::-^;GTM_TC(O[-Z^O
(O?6R>E&T)UE,T2BNLgT:A2JeI(GCTO0YE&:V5NXc(^#M(N)R0BNf&Ja>^06?TZc
-X7K@(e1JI^R4g-O8&F?XA4]-1;5K_aC+bQ6&K?O@f2R@QA^MSL]Ca/OX3K0>P5X
#(//NM[8MEN]@<+].5e,Sdf#Y_g.d&VFdg1d?[;Ca;A@c1cg,2bd;\,QP(d:WC+D
1P^?L51DEg=>?RBH8JK0\97&3CEGO_41:X-0N#faf5<;Q#72eQ)QB<M[GL(0L(1g
gdHT5^.Z[G000d-f/BIR2Wc0>QBJ78f;P24LN4:YH89WI<C.f@gN>(U]W[c77PL,
X#/RO;^R>[)(e/,cT[30KQ>,dLM\b7+<WdI2,1?f+:EHM1RL#4&TLLH5_,(<U3Y5
P4I-\S8UCc@\XJ-E6\<72LWfNLBG]>]&_#?f&Ld+Q,<:WM-Z(d7D65-;/KFM[aXS
Q@1#^Geab;d&WPTV&88L.R>12G\(F^(4b\-+RL#BJf/+MIE2L?B=fX?ZLQ_P>-X7
IR1@Y><(.NbDYf.B2DLD(BV/-bF\7\#TeNa0S^G3a5=)?;.gAb65FQ:NS>^c7?>Z
_E]e8DeF=GfQ>TcGTOOR7#EX=d2AbH+6.,?4Z].0GHHR[;d6S)ALHC=[H0Z#Z5>/
-VV3R3934@;K85+2:6Jf].M-3_VZ-O46)&.44(:6=(2-->+8a_CAbgT(C.O(MI3@
]DgR)Xd-4OI6bDH>9+3f1,6N0]QH<fMTgCe?UR_U^I1I,UL(@@?/2OLY(/0B)PQT
)LGE9_aSbT,bZ]/47I[1>KD-DBGB?.WbI]bD51+2FJ1+..3[,9b+ZBTZZLYI1>Hb
;^4GM6bCa2E,7Ge2-D)d<@DD0f@Wg]TW>WHY.-F+/cF@>)c2A+IE:e@TAB,C7HS3
PY@/_]V3#e//>PFHQ0;I0STEbRAP(3E)>=1/[TDF4T>4\>eQJ();I00(4D>F][0V
BN8RO.\Tb>f8c>(7S;^fR=]N4Z^M[?7O#8Ia6,-Y/K&\3?D1<F=3cd/JR5g&ZD,d
\E<@69G2+C=V:1dF>U8MQ]]c+c]&gK2W(1T<(,5.:@H[3VVaIK52UIdQ#]Y]f.<=
_b=2g.36eM/NOIRg(=T#D6=>D/Z_08T7PBID__b0OJ8.[I.Y#NN#PI;^>8+)R-Gc
DdO#ABOK_<)\We8ULV+MBfG>2A4Z)<>K;7<6aY=;G;dLFHS4T+3gHceb40H1\CL)
GdZ,R]_RZfeY4NJN.1UJ,I=2+3&SWCb4Q+-e,8Efd[b(bE4P[K8XY_dH1]a597VZ
dIaeWUbY@MH[(8M6?_SJ52K-\3a@TT2d3F_5-I&:;U+fM)DWXO<M_)[7UB4))6fG
EX7Z7)bIM]^>19Wgd2+Q&H;^_8b,_J[LAg:Q/dO&8>858-9N>+AN5A,45(e2+IQb
Z6cccEe<]e/<LJ&]=.M<8S4XL#Ac\G?_]T)aTaUV13V6RF0.HUH=<JIK^]7aW4&+
6-JVKI[92_Xa7eF?5D6b#MCU7W:_5E5@TW0@cCSY_013=S<48MU]3[BO&cb-,EL-
J8&2A_W5[])TcC&HK3H;YSG1J.MAM^BbVf@,eRM]MdGYS=^XUN,0X7L,N7JK2WSZ
&929K<0TgOb=.51G<>9f\@.EJK#>bQB??5#b[01E_H>WD2X;Z\1\K(TQ^.Q_K@QD
O.A?)+E16PM/;-6C.<GGW&\8Ka0E)EHV70F\@C07KK1)[SG6BMXdAG+N02+[:3>G
)V_-.gWW1MYOP7E[F7Z1?1]N0XM39/+6DFZA1T<=R_ddBFcBUJbJ)SRg,eM,#QbQ
<FP4]GDd&=_c:WS3\bZVX_ePQ_7D3MR7S8&3;?TASPVM/Z_d?>,=MSKH>/H:EMDQ
Z(4(V5MAJVTT?.=CBa(5W\48DND:4#X:Y97IeCf^OJTZKZ_-L#fM[OdUVF/fHgC.
GT[d-6&L^I]5-,1>4@-IH2b+ZZc=CFITde1^b3N+N270Z2eQY(OS<O-9FU03K2[R
^^RKT_-L-+HaVc.-WDP[=:-9^53e=63bG@-,aRM^Ug;3K[7Qf&I>9X+(VgINKSDX
(GBVR4_f+^>+@[&C(LFV@:caRTVJ56<U(X_.IW._^<T=fcf-E1PfaWT3fbK[\A,)
Md/.P;>O#83NCYNLU\JT/T1VRPW#+DB0^JZ_3+2GQ0-YTSMCLS,^A);XMA_+1WaO
ab=]=(BP00G/bF)#:8Da2/:M[TOH36Wc.O#8-N^EGM@LcL8f\QO=2c?<&+G5ae50
T-I5F5LDg8_+=JF[gBC<cO:^2<b)?N,aUJV?H<dC?8P;8P_.OU1:Q?TE#97Q]D0F
N_L).Z)3RYU5FWDN6J\gWAa+6#JJ48Y2Q=;CU\=W5,O9R[#^WEQ8aADW>dL.P<Hd
5gLX\SITGZRNb\Qd0-(aYR,4,A_C)=Ka]T&1TJ(S/,fM2g[RZ?5I^@1>b:B,DYAQ
WfT26,M\T6Lc8#C1PQDE/,,5g=8GU.d0CG98IgL\<3e&P/1c.OAD\:M\9BdSJG)7
-6GJNf/TG7U[AMY_R.)ePHOWSNN>?[#A<0Q5:eJe3,37)D0S&R0.50A8:-0bRB>,
H,?fb[W?f#?@JN<ORNed3L;F-ZA63LP=^DT\956^H#S.<E/(JgFA=SDCZ5(E6Yg1
OR,K]<4N_e)>XR+:)-FST>Z]]AT]<(.9/BU91S(LY[HIYJff_)>5YNBSKU.YLIf4
baYc>EW\TY5QW0d>7JOCAdK6H?IFA(Y2Ygd0gWaQ:)YWeJ?.ZE:MSV3TCL.M5CJ,
IeS+XC+=L1SEa36GHLF@7g:H/Cc,@cPF7-:[cf[8G5OEfJHeB/^fSD7CQG=MFWI/
+gFZ.YM9;&)&^Q:/&O]D0S6-^PM.FW7Cb#;N1T.^Y6d^.L8G@fZ,SbT64]4?\JRI
5Se&_4Q,2eDCP]M_DHa.EKMNdZBCC9BQCL8XaKJ3<g@?0_3T=[IcY2H:7&(GAbcA
7KV(\9Z8OZfLffea(,N8G>\DPX>dUHL:@SP2J5PU9&J3Q3PKZAX9VVgJ,07)I]c7
I(2GV\Q]0\b5DeP07Dd12Xg;]QJ3VYNDEU+E.&&?-W&]PU2GRRZUO+\;a<\W93V/
SOI\&1EQDOM[G9=LW<VHBYDb)S<>7T7K<?=HK/+.I3<ZB=D[72/5J5M;\;I<b12<
],TUN9W3D(4beI4V&UVB+18fU1M;(O7e7-YZDO[_YaBX1,MM84LRXg?3.15_)LJ:
TN/W1/B=15[QRfD\II>ZbT3FX;_O644\I()db;V9PW5O_/aO47YYR4(C<F[_7d:0
J:?HE;-gDXI<)Ug[L>N\9W(>1Eb(Y[]Ia.5_M=;>PReQ=2PU:U:G^TTL#I\PUV^L
ER\:47Y:aL<:=(TIIMPf@=bXA\aXb/K5=M=+d#CK/[WR-:&^[,Y[MF_C3.,L;L_#
R/QPZL1\LS:?.6O75G^GR2XJ9325.7[fa-Pf&ULJJ5?\e.ZOGR,bTBCd9g5[,1W,
IZJL0+;=Q&)3eVVQBZYBCSbQ06P@?1NDTWeS04c/Sc>:D+<PWY+VO0D4f[E:/,5F
K(&g5I?CPfCfQHI70g^]1Tc.64f-=(\XIIBB?3]Hb#V;g->(Z:aXXR)>KE?,Z>;Q
R=HE#cQfN2bb+(]X=SBI5+4NCS3<-J6=?Y0#8-:f=U+Y#]<(a96OK<M/53aQ&GJG
U(Hg834MGHY-]ONIMC:VaEZd0RfT1SI6UWOe<MG_B2724&+bVd787abY?Vf_OVM@
,KSfGa1Gc3.Z>Vc/54.(&_C]6X@Q#1+S3XGb5T2e54#C-a_Vf#(BT6.0^c<<UXJ#
fQEf6dZ0L&gIBN=XU:_bceXff<,8W9V;PW/AA:2HGJ]FMO@d#+:_Te,LB):18<gH
a>I/&+\4ZXZB?A@U_H_bV2RU_[-9cb\E33d8_2U=1@/-=6UV>\ZN9]G&#,M0c,c/
Zg?(.@))4b&Q:PS9-]44.aPQS(-9]>Q\YOcM<\a@C+7][<NAB5IJ;R-Z2Jd-B3S3
^e596@dPFXYE)XS8)5D/(/K1QJ(_]\K:6JJ1FJU/<.Ub.R#>6:eYMW2Gd+V7-F,)
c@/a6Q#6#7Qa4S/)dTPP1R7_>VWPLD>3LVC1HFLW^/<@d3&PUb<.cTVXHD-(4S=/
(BPTE8fV@2cPNEH8CM2gN,)01PDO5[CE9X+(@YVK6K5ad53g.f,dBEE/E)1dVOK4
LEF+]/BXZ(C485C.;/PS5Rb&.A\Ad[GAEe@8AR-Vb]5Te0cV&X>GDKK4WNRQI>)C
R[^B0A,K1L7.fT7DgY<]eV?IZ.(_\QR3SKd\K=aF\\PJ_WJ#F3+TKN-XK#OGfdQS
OgEdG6OWe.^S^7P\<M_NZA?\9Q#4Wa#HeZb9N[8/:Kd<91-/WcR>STca9S9CC_3M
KYe7EK@2F\&X[&I3D)YF0XVX#cJeES2P-U?XWKN&Z+6_-KfZ0g#NWW3H/@aAH_G9
5X#D2f=PH>;R9S+O4,UO/9J4cG1^3J8Gg&g7<0.QZOJ^=\[#D@PX3a\B=4@/@PUR
6JQT@7dFUI<JO.4.#e]F-1X/(c<MB#QD5?-a@3(DcFR6C1bI&HSM-4T+B=H<)b[\
N=Sgd]3bOS8,^V/JY+EIQYI4I.,\#fQVETD^09BY3),AB/RM8a\0]?5R?R4=R[?=
/0c&QD:&^He(;e)#Sa)FXI6=KEaeN_3H:Y0Ud?)J_+gg#GQX@\U?[B&I/+&.:Y4)
FBG,ERb5,Q?W/7=a;J2MX)8X;Hd.#Z4()30#OAVa>18ELE80ZSbN[\#NR)VeHG4F
LY6F.Bf(9)</5OZ9QU-[-M<PPPYE8D^7;,>)GE]5)KH:@_M7V_/9\]0+Ncd&ePI,
,dX8[B&VV3gK;4P]La57:K1(NYACO8ccgdE31/W7)6eDg&Ee2[dERC+=f4#NQTQe
g#f3JI>XU#[WJT2d.Q<O1EaR0W@;9KgHPL^D^:ad:,UGb@L[IP?d:f#VS>e@Y:Ga
/MP/:2:.8M#0d\eGS[fa_aga-c2eB;YEeHWQU\7+8#AQZ;a4aH[M,=@O-6X[C&U]
SJ3O-ddB=?T-ZWHS7X]#D-&9Z_R@OKKW95D2/_Xd4K,=O@6/CZM0-EZ+6]WJ^V-e
B@RQ<Q,^4Q1Vf(1XWCG/cDfaB89.\?2]a-4M[6\PMbK#01fa84,HbJ7EZ#1_)^M&
4H[KHT??(S27E&;7I[,JG2YCGb]#_2=]40,82I7;1a_F8:1T,Fb3VY=f8GZI:8M3
EfU(d09(&c#8fH^O&XHL\&,;ED^&G:D.g4BfK,P1QV)->daR2/N4b.J\M/5.R2I#
Yd/B+6Gf3YF5YI]K@DMaU23M6L<7=?N5+gHJ<>V@FP^89N&35S)TTK<B=Hf:g2][
0H)YGE#b(Vg#<K&-ae9FN^>VH.D9cda)5Uce-.KcbIX:FB@ULG5cM9cDM3E[FbE;
J=DdMX>9T:;YMQX;^fVc_SZXZa5B;99U1Gd+Z?Q]J[YePB?=,eb\KJ07<?IN4&e4
R<UF94TQGF)d225.1g^_&?:J9c#:HB[SY\]V2PY9X&N623]BWRfZ;T_48GcZ-<6e
;G;@@LVTb.J>?9V+e-HR#4+@;YXQ90DV;L,50;X#0:]<Pg]OA\5=3Xd:e[Y#M5N0
DX>Ec\_Q;YD_ZGASDN@=-/Q_^IEcgeDZN636G2/bJFKDPbS7E9d>;IZ:ME(]:?5_
:04dL,g]dJ5YEOK5-:,T_M+</-QR([423R-8Z^-egaX-)00<dE=TIA@;I]g]:_cT
BP_G3OANRH[KD9EH04TAHD3e3^0.OG>/A-4G>>U<YNb_RBRXO0<.,2<dSYU8WF+]
Uc\8^O>gbKfT]\SL>>]8+5&,C)<e2T3XMQ93\P:/7=J>R]XL5V(/G8FCd5^FDJf^
_WXF6:HYV8D](KD;-.\I(WTK6,Va(.(VY3)\]W:]S3:@)<-S(NE#J&1-.MZW=K5W
B8S:XFZ:+P88</153gMUN<:A\V4P+UTM3g0YMBTC^\XV^LQI5/#)JL92-Kd]U?H;
dB<I1)]eZAB]MDYI<Ceg;NUd)g)&dZC_>GZXS(ERd9B=LM)(N<Ad2&]BA+9C7feO
4/Y7f-9C\P^)@a2BL^Z;4GQacPg.W5.7N>:]X6#/UFPY_X;EgfQ=AG->6OK+7&Y8
3VR,b#=-0(L-OT#FGEF4@g_N?)2]gKFg_-Z]M-##//V,U6#RVb[#@E4/[Gc06Z+W
X\)B.8787O:>+I(P11_L?FYJ,4dW@;aJcDC3CSG<<F]B@Y.6C)TX6Z(TT5e,AD5,
?(DPa[P,5N4(XI6b2Hb&3JMX;PM,&S+5/f75P0[fLU1a,c+H;?,M2b<g9?9[;SL[
Xc1:bCCVf^THUH3+MY1P=7PL:B+KFeN1R;Q]NE0[)5+@(.W[-SJM86DSRGI)\eYa
(+-7@40QK.W9<4^9B>B<UZJ2N.MYH=2f]Tf:;[T-#>[[9Ha:eQW1JH4aUEe&HcU4
#YY8CTbCI)N:G^2MG[\0)48?5ZMbW6H_HIGSH\B8F,dZ,IFC,:\c^XL9<-P,KbT-
_L/N@SY-_>+(]:UeL(S3,[^?9>2Z5<4692)P#B7-Q8IE)Q6VA/A0eBW);>CO?=RB
9[,JE&B,UKN#)0M+e._@+Q95OU-#GPKA@We0M8d5c4;P6D5&C7OU#,49RYJDQZMc
B]:G7bEYH9\BS&HR.OKC\V8)JCRYFE0,2Y0&;X-FQ>f2^>-3cE@b&X3L:,BW(cdF
LME5MPPcWe)>fK6@4)_@e^T2</RPSSe6NHf2B6^H7,22;Z]Y[GW>aJB6]11gGF51
Q?2Mgf:+^CA)g?:W(O#0a-R#/fI;/NKOd1R_^4Sc1K-aIN@AS5_>6@+QX4#eYO2M
MKS9L.477/Y@M@J[T7^P=Teg&_4BE-,T:cTL/LIU@BTc=U<;2O:&@&W3VOa2Wbb3
1b+AJ0#^]3J,PM-F]Efdf#dEWG@b,:A1DM]@H>M5-&96SEBV_]XTXX8FL]Q=G?E@
N0HLKC6Y)#83+-NfF.N;WGUM/6?:/-:V3[:dK6cU3LX9;UagPLW6?bRUd11.Rb&O
;M7F11[&Z\Vd6Q#C]EIF-f5FfgZgd^EJ>g4.:25OGB>RX:9EC1MbaS0Fb1_+YXRB
eG)NEd4Jd\Q?+SfJ]VR</MG4R\/?OW#fM5??)a=SA6ED2L/O68AG9X?,61d5W/<<
K<#,>WI));PD-1M+VID60\8ZY?BS:,f+4(2V>=S0[0Z7+E+JAYE<K9=MT(?\Q^YG
==M)2ON7T6;E?7^]8A_#^3Hf27?JGI]fYg-1;3((TXG+]NNI;Q:a3b9@>W2Q>-X_
6RK_8BMLd(8QZPZfI&#SMJ#:X]Q[BODJ:@M2LCW&g67Nd[4NYaXDd/9,I/4\ADO=
)ZUA<ede1IYP3SL#O@d[:8O;I[4,1)aBB5^._fBK;YG.,C:MG(.NRbPb[K0P<KV5
:SK9>gGFQKQ,[Re(U0S&g]He:S3B9Y,:K,22330b<LD&b)a=NX33Y]@e)RaOP73A
Q&NKZ??LR#[U[(GJ]8=,2LI,a-=aKN<XE96R0E?c\0T&[d]aJL0V7^&.X5L8b-#6
_FHMV,3(B,3Q8=c:B8[dT(L>HDYR71X4+7IY:(L_HYM8cG/SGO>4-=f_8+g.5>VN
/W-.1D==>LJUIc0NPB>D;&KRV[CP1T70Qe+T8VfUS:Uc0=L3abOaL\FK^HBJ5:ge
fWcYZ(Yd>G:RY.X,J<<c.U18IIK29-K.^(]C/EL[>[VG&Fd936+8XRH/X0VL0?5Q
U_4f6Vg+M,]1R3A[Y/U3_7Y4B^3&6;#H4L/,86.<\RV))[QE7IK#XBd@cGI=<Z2]
(,4S@[\-3T)\C9,D=F]9B,KIPL@2(TCa/>CN0Q4f-JI5I+O@N.cGbR_MU<W4XV,g
F3D[WKKMWOPWddMSVf-/a?d<7I#5JJ#?6SdZ.D^&Y4[g]AK^7F?:K.TX:C,\ZEcQ
F:L;K3B<f@e<9_0:c?E7:d[QUPc19:7J5.0)?8:PG=d2fgZ84/#=<)#RRJPAW;CU
8FEbS^F:<Z[H6_X1MJQQC?83F]A_[QH5X;DTPL-TTg2bQScOW,;dfX-D4OM#R4Q.
SgV>^M];dEVH+$
`endprotected


`endif
