//`ifndef A_WIDTH
//    `define A_WIDTH 32
//`endif
//`ifndef D_WIDTH
//    `define D_WIDTH 32
//`endif
`ifndef NO_OF_SLAVES
    `define NO_OF_SLAVES 8
`endif


// ******************** Global Parameters ******************
// Please change the A_WIDTH & D_WIDTH with the respective width
// of address and data bus
parameter A_WIDTH = 8;     // Address bus width
parameter D_WIDTH = 128;     // Data bus width


