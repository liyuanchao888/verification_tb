
`ifndef GUARD_SVT_AXI_CACHE_SV
`define GUARD_SVT_AXI_CACHE_SV

`include "svt_axi_common_defines.svi"

`ifndef DESIGNWARE_INCDIR
  `include "svt_data.sv"
`endif

/** Add some customized logic to copy the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COPY \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COPY) begin \
    svt_axi_cache_copy_hook(this.__vmm_rhs); \
  end \
`endif

/** Add some customized logic to compare the actual memory elements */
`define SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE \
`ifdef SVT_UVM_TECHNOLOGY \
`elsif SVT_OVM_TECHNOLOGY \
`else \
  if (do_what == DO_COMPARE) begin \
    if (!svt_axi_cache_compare_hook(this.__vmm_rhs, this.__vmm_image)) begin \
      this.__vmm_status = 0; \
    end \
  end \
`endif

//`define _SVT_AXI_CACHE_DEBUG \
    //`ifdef SVT_AXI_TEMP_CACHE_DEBUG \
        //`svt_amba_debug(cache_name,$sformatf \
    //`endif
// ======================================================================
/**
 * This class is used to model a single cache. 
 *
 * Internally, the cache is modeled with a sparse array of svt_axi_cache_line objects,
 * each of which represents a full cache line.
 */
class svt_axi_cache extends `SVT_DATA_TYPE;

  /**
   * Convenience typedef for address properties
   */
  typedef bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;
  
  /**
   * Convenience typedef for data properties
   */

  typedef bit [7:0] data_t;

  /**
    * Enum to represent the different cache structures
    * DIRECT_MAPPED: An entry corresponding to a main memory address
    * is stored in a cache line with a unique index. For example,
    * consider an 8 KB cache where the cache line size is 16 bytes
    * and there are 512 such lines. Then addresses 0, 8K, 16K, 24K etc
    * are always mapped to index 0 of the cache and so on.
    * FULLY_ASSOCIATIVE: In such a cache structure, a given main
    * memory address can be stored in a cache line with any index. 
    * TWO_WAY_ASSOCIATIVE: An entry corresponding to a main memory
    * address can be stored in any one of two cache line indices.
    * For example, consider an 8 KB cache where the cache line size
    * is 16 bytes and there are 512 such lines. These 512 lines are
    * divided into 256 sets with "2 ways" for each set. So any given
    * main memory address can be stored in only a unique set, but within
    * this set, it can be stored in one of the two ways. 
    * NOTE: Currently only FULLY_ASSOCIATIVE is supported 
    */
  typedef enum {
    FULLY_ASSOCIATIVE   = `SVT_CACHE_FULLY_ASSOCIATIVE,
    DIRECT_MAPPED       = `SVT_CACHE_DIRECT_MAPPED,
    TWO_WAY_ASSOCIATIVE = `SVT_CACHE_TWO_WAY_ASSOCIATIVE
  } cache_structure_enum;

  /** @cond PRIVATE */
  /** 
    * The minimum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_start_addr;

  /** 
    * The maximum address in the shared region of memory
    * that the component where this cache resides in will access
    */ 
  addr_t shared_end_addr;

  /** 
    * The width of each cache line in bits
    */
  int cache_line_size = 32;

  /**
    * The number of cache lines in this cache
    * The cache_line_width*num_cache_lines defaults to a 1 KB cache memory
    */
  int num_cache_lines = 256;


  /**
    * Flag to indicate CHI ICN Full-Slave mode. Set when CHI Interconnect is
    * used in Full-Slave mode.
    * Default value is 0.
    */
  bit is_chi_icn_full_slave = 0;

  /**
   * Indicates whether the cache supports storing poison fields
   */
  local bit poison_enable;

  /**
   * Indicates whether the cache supports storing data_check(parity) fields
   */
  local bit data_check_enable;

  /**
   * Poison granularity: number of data bytes corresponding to a poison bit
   */
  local int num_bytes_per_poison_bit = 8;
  
  /**
    * The structure of the cache
    */
  cache_structure_enum cache_structure = FULLY_ASSOCIATIVE;

  /**
   * Indicates whether the cache supports storing Tag value
   */
  local bit tag_enable;

  /**
   * Indicates whether the cache supports partial cache states: UCE, UDP
   */
  local bit partial_cache_states_enable =0;
  /** @endcond */

/** @cond PRIVATE */


  /**
   * Sparse array of svt_axi_cache_line objects, used to model the physical
   * storage of this cache.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  local svt_axi_cache_line cache_lines [addr_t];

  /**
    * Array of addresses mapped to each index of the cache.
    * Whenever a cache line is updated, this is also updated to
    * reflect the updated contents and may be used by the various
    * cache access methods depending on the structure of the cache 
    */
  local addr_t addr_mapped_to_indices [int];

  /**
   * Sparse array used to store the number of reservations for 
   * addresses for which cache lines are reserved.
   *
   * The array is to be indexed only by an expression that evaluates to an 
   * address within the bounds of the maximum number of cache lines in the cache.
   */
  //local bit reserved_cache_lines [addr_t];
  local int reserved_cache_lines [addr_t];

  /**
    * Array of addresses mapped to a reserved index of the cache.
    */
  local addr_t addr_mapped_to_reserved_indices [int];

  /** 
    * log_base_2 of cache_line_size used for aligning
    * addresses
    */
  local int log_base_2_cache_line_size = 2;

  /**
    * Semaphore to regulate cache access. Components using this
    * cache model can use this to first get the semaphore before
    * accessing the cache. This is useful when multiple processes
    * are accessing the same cache. 
    */
  semaphore cache_access_sema;
  
  /**
    * PA writer handle which is used to write the cache data inside
    * FSDB. The data will written out only into FSDB and not for XML.
    * This means the handle is instanciated only when FSDB is enabled.
    */
  svt_xml_writer pa_writer;

  /**
    * Transaction UID
    * To support cache operation to transaction relationship 
    */
  string transaction_uid;

  /**
    * Transaction type
    * To support cache operation to transaction relationship 
    */
  string transaction_type = "";

`ifdef SVT_VMM_TECHNOLOGY
  /** Shared log object if user does not pass log object */
  local static vmm_log shared_log = new ( "svt_axi_cache", "class" );
`endif
  
  local int dbg_indx;
  local string cache_name = "";
/** @endcond */

`ifdef SVT_UVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`elsif SVT_OVM_TECHNOLOGY
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param name Intance name for this memory object
   * 
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
  extern function new(string name = "svt_transaction_inst",
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`else
  // --------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new instance of this class.
   *
   * When this object is created, the cache is assigned an instance name, 
   * cache line size, number of cache lines, the cache structure and 
   * the minimum and maximum shared address.  
   *
   * @param log The log object.
   *
   * @param suite_name Name of the suite in which the memory is used.
   * 
   * @param cache_line_size The width of each cache line in bits.
   * 
   * @param num_cache_lines The number of cache lines in this cache.
   * 
   * @param cache_structure The structure of this cache.
   * 
   * @param shared_start_addr The minimum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   * 
   * @param shared_end_addr The maximum address in the shared region of memory
   *        that will be accessed by the component where this cache resides in.
   *        
   * @param is_chi_icn_full_slave (Optional) Applicable only in case of CHI
   * ICN Full Slave mode where it is passed as 1. Default value is 0.
   */
`ifndef __SVDOC__
`svt_vmm_data_new(svt_axi_cache)
`endif
   extern function new(vmm_log log = null,
                      string suite_name = "",
                      int cache_line_size = 32,
                      int num_cache_lines = 256,
                      cache_structure_enum cache_structure = FULLY_ASSOCIATIVE,
                      addr_t shared_start_addr = 0, 
                      addr_t shared_end_addr = ((1<<`SVT_AXI_MAX_ADDR_WIDTH)-1),
                      bit is_chi_icn_full_slave = 0);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
`ifndef __SVDOC__
  `svt_data_member_begin(svt_axi_cache)
    `SVT_AXI_CACHE_SHORTHAND_CUST_COPY
    `SVT_AXI_CACHE_SHORTHAND_CUST_COMPARE
  `svt_data_member_end(svt_axi_cache)
`endif

  // ---------------------------------------------------------------------------
  
  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   * 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given index.
   * If the index does not exist this function returns 0, else it returns 1.
   *
   * @param index The index of the cache line to be read.
   *
   * @param addr Assigned with the address stored in the given index. Please
   * note that if the address specified is unaligned to cache line size, an
   * aligned address is computed internally, before doing the operation.
   *
   * @param data Assigned with the data stored in the given index.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line at the given index is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line at the given index is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line at given index.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given index
   * has an entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_index(input int index,
                                            output addr_t addr, 
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   *
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0 );

  // ---------------------------------------------------------------------------
  /**
   * Returns the contents of the cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param dirty_byte_flag Returns dirty flag associated with each byte in the
   * cache line associated with the given address. '1' indicates data byte is dirty
   * '0' indicates data byte id clean
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is off
   * 
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit read_line_by_addr(
                                            input addr_t addr, 
                                            output int index,
                                            output bit [7:0] data[],
                                            output bit       dirty_byte_flag[],
                                            output bit is_unique,
                                            output bit is_clean,
                                            output longint age, 
                                            input bit record_to_fsdb = 0);
  // ---------------------------------------------------------------------------
  /**
   * Writes cache line information into a cache line.  If the index is a
   * positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param retain_reservation (Optional) ensure that no existing reservation
   * which was made for some other transaction is deleted. The cache keeps
   * track of the number of reservations on each address. If this bit is 0,
   * with each write, the number of reservations on the given address is
   * decremented by 1. If there is only one reservation on this address, this
   * write will result in all reservations being deleted. If this bit is 1, no
   * reservations are decremented or deleted.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the write was successful, or 0 if it was not successful.
   */
   extern virtual function bit write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit retain_reservation = 0,
                                     bit record_to_fsdb = 1
                               );
  // ---------------------------------------------------------------------------
  /**
   * This function writes into the cache via backdoor. Backdoor accesses are
   * direct accesses to the cache in the VIP by the user in the testbench. For
   * example, if users want to preload the cache from the testbench, this
   * function must be used. This function does not delete any existing
   * reservation made to this address by some other transaction. Reservations
   * may have been made by the master VIP for transactions to the same address
   * as what  is requested in the backdoor write. Using this function for
   * backdoor writes (as opposed to using the write() function) makes sure that
   * those reservations are not deleted.
   * 
   * If the index is a positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param index The index to which the cache line information needs to be
   * written. The range of index is between 0 to
   * (svt_axi_port_configuration::num_cache_lines - 1).
   * 
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param age (Optional) The age to be stored in the cache line. If not passed, the
   * age information is not changed/updated. Typically, current simulation clock
   * cycle can be specified as the age.
   *
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   *
   * @return 1 if the backdoor write was successful, or 0 if it was not successful.
   */
   extern virtual function bit backdoor_write(
                                     int index, 
                                     addr_t addr = 0,
                                     bit [7:0] data[],
                                     bit byteen[],
                                     int is_unique = -1,
                                     int is_clean = -1,
                                     longint age = -1,
                                     bit record_to_fsdb = 1
                               );
   
  // ---------------------------------------------------------------------------
  /**
   * Gets the index of a cache line corresponding to the given address
   * If there is no corresponding entry returns -1.
   *
   * @param addr The address whose index is required. 
   *
   * @return Returns the index corresponding to the given address. If
   * there is no such entry, returns -1.
   */
  extern virtual function int get_index_for_addr(
                                            input addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the address stored in the cache line at given index. 
   * If there is no corresponding entry returns -1.
   *
   * @param index The index of the cache line
   *
   * @param addr Assigned with the address stored at given index. 
   *
   * @return Returns 1 if there is a cache line at given index, else
   * returns 0. 
   */
  extern virtual function bit get_addr_at_index( input int index, 
                                            output addr_t addr 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Returns the index corresponding to the least recently used cache line 
   * between the given set of indices. The least recently used cache line
   * is the cache line with the least age. 
   * @param low_index The first index at which the operation is to be done
   * @param high_index The last index at which the operation is to be done.
   * @param is_not_reserved Indicates that the entry returned should not be
   * a reserved index.
   * @return Returns the index corresponding to the least recently 
   * used cache line
   */
  extern virtual function int get_least_recently_used(
                                int low_index,
                                int high_index,
                                bit is_not_reserved = 1
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry for a given addr. This method removes the
    * cache line from the cache for the given address.
    *
    * @param addr The address that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_addr(
                                addr_t addr,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
    * Invalidates the cache line entry at the given index. This method removes the
    * cache line from the cache for the given index.
    *
    * @param index The index that needs to be invalidated.
    *
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit invalidate_index(
                                int index,
                                bit record_to_fsdb = 1 
                              );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address.
    * Reserves the given index of the cache for future use. The get_any_index
    * function takes into account the reserved indices as well so that a user
    * is always given an index that is neither currently in use nor reserved
    * for future use. When a cache line is written into an index, the corresponding 
    * index is deleted from the set of reserved indices (if present).
    *
    * @param index The index that needs to be reserved.
    *
    * @return Returns 1 if the operation is successful, else returns 0.
    */
  extern virtual function bit reserve_index(
                                int index,
                                addr_t addr
                              );
  // ---------------------------------------------------------------------------
  /**
    * Gets the reserved index for the given addr.
    * @param addr Address for which the index needs to be found
    * @return Returns the index.
    */
  extern virtual function int get_reserved_index(addr_t addr);
  // ---------------------------------------------------------------------------
  /**
    * Deletes all reservations made in this cache for future updates in cache.
    */
  extern function void delete_reservations();
  // ---------------------------------------------------------------------------
  /**
    * Delete or decrement reserved_cache_lines corresponding to address
    */
  extern function int delete_reservation_for_addr(addr_t addr);
   
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_unique The shared status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * A value of -1 indicates that the current status need not be changed.
   * @param is_clean The clean status to which the cache line associated
   * with the addres needs to be updated. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   * A value of -1 indicates that the current status need not be changed.
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_status(
                                addr_t addr, 
                                int is_unique,
                                int is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the status of the Tag held in the cache line for the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param is_invalid This specifies if the Tag is held in the cache line. 
   * A value of 1 indicates that the corresponding cache line should not contain Tags and the Tag state
   * must be considered Invalid
   * A value of 0 indicates that the corresponding cache line contains Tags
   * @param is_clean Specifies the state of the Tag held in the cache line. 
   * A value of 1 indicates that  the Tag is held in clean state. 
   * A value of 0 indicates that  the Tag is held in dirty state. 
   * . 
   * @param record_to_fsdb Indicates to record the cache operation into
   *        FSDB for debugging. Default is on
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit update_tag_status(
                                addr_t addr, 
                                bit is_invalid,
                                bit is_clean,
                                bit record_to_fsdb = 1
                           );
  // ---------------------------------------------------------------------------
  /**
   * Gets the status of the cache line for the given address
   *
   * @param addr The address whose status is required.
   *
   * @param is_unique The shared status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is not shared 
   * with other caches 
   * A value of 0 indicates that  the corresponding cache line is shared 
   * with other caches 
   * @param is_clean The clean status of the cache line associated
   * with the address. 
   * A value of 1 indicates that  the corresponding cache line is updated
   * relative to main memory. 
   * A value of 0 indicates that  the corresponding cache line is not 
   * updated with respect to main memory. 
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
   extern virtual function bit get_status(
                                addr_t addr, 
                                output bit is_unique,
                                output bit is_clean
                           );
  // ---------------------------------------------------------------------------
  /**
   * Updates the age of the cache line associated with the given address
   *
   * @param addr The address that needs to be updated.
   *
   * @param age  The age to which the associated cache line is to be updated.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit update_age(
                                addr_t addr,
                                longint age
                              );
  // ---------------------------------------------------------------------------
  /**
   * Gets the age of the cache line associated with the given address
   *
   * @param addr The address whose age is required.
   *
   * @param age  Assigned with the age associated with the cache line of the address.
   *
   * @return Returns 1 if the operation is successful, that is, there
   * is a corresponding entry in cache, otherwise returns 0.
   */
  extern virtual function bit get_age(
                                addr_t addr, 
                                output longint age
                              );
  // ---------------------------------------------------------------------------
  /**
    * Sets the protection type of this address.
    * For is_privileged, is_secure and is_instruction arguments, a value of -1 indicates that the existing value
    * should not be modified. Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address that needs to be updated.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_prot_type( addr_t addr,
                                     int is_privileged = -1,
                                     int is_secure = -1,
                                     int is_instruction = -1,
                                     bit record_to_fsdb = 1 );

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the protection type of this cache line.
    * Definitions of priveleged, secure and instruction access
    * are as per AXI definitions for access permissions of AxPROT signal.
    * @param addr The address whose information needs to be retreived.
    * @param is_privileged Indicates if the address corresponding to this line is privileged
    * @param is_secure Indicates if the address corresponding to this line is secure
    * @param is_instruction Indicates if the address corresponding to this line is an instruction
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_prot_type(addr_t addr,
                                     output bit is_privileged,
                                     output bit is_secure,
                                     output bit is_instruction);

  // ---------------------------------------------------------------------------
  /**
    * Sets the memory attribute of this address 
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address that needs to be updated.
    * @param cache_type Memory attribute of this cache line
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_cache_type(addr_t addr, 
                                     bit[3:0] cache_type, 
                                     bit record_to_fsdb = 1);
  // --------------------------------------------------------------------
  /**
    * Gets the memory attribute of this cache line.
    * Definition of memory attribute is as per AXI definition of memory attribute for AxCACHE signalling.
    * @param addr The address whose information needs to be retreived.
    * @param cache_type Returns the memory attribute of this cache line
    *
    * @return Returns 1 if the operation is successful, that is, there
    * is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_cache_type(addr_t addr, output bit[3:0] cache_type);

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
lvRN4QYaXQlEEcoNxHI//PNt6PfmfxCeRnDWI2MjLhDDyT0b4YpNs7Na97ge16ex
4eMgPzxuowTB/h6wizhnd9bq6FyYwRjEQWY76w3BgFbOUroljWfMun3xXQDpM8SH
c5MznOq3h81pY5j8co5K7xZ0zPBqzHw3DZfvZn5OfIA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 802       )
sJR4WMr7hMBl2ZEEWhPh6oXvl2tKktJhYDEl44/mSMrLRcB/DpuHf0ue14CfLZ6c
NOGdMb96nzxkxtuOYNqd9ETRw9Aiwc2qup3ILOxy+QIzzJlvemZOwZweCUq4c7yx
y8nhqFRJKunU/R+pROoHfue44ZJ0tU3WvoOyB2Lwap7Jds7Dnb4IrQczwTS29572
Wn/9lryB5Ru4kGAR3VEhiGhYPdqmQGlqFy1asTr80aIchp2YGNKVOTLLndPWG0zr
nr1d7Xfn2he9zHF9Mnus9mcWPKcabtAD+S5HDQ+DGfvkSgosNCbcIXewjk8FTwwX
NJnq1Qp1c+AV4G8u/1V3LtP2JFSuikn6TQS0OrtVxLCrjir5y3A50W8OOLVTvD2p
GL2pDzNV0DoEJXk4MsIKASirxSf1DSJKJB/bscSq+zIS0Ub7oX0SygsoKsyeSddf
zTNg4BjVOhjX4otwO60+xgKfi2beDwKqQ30Es74jtulMBj/QTuKR9f4Tq4j2dRol
tID3qPZyUrHk7/71fZSziXzb3L2z4ElLBNNR+DCyPqUXn9IiLAzEJ0GXJOyd1SBG
4KPldkn2uYn27YyXU4bH69+qwZ8hR7xpaL01VRHLXiJNDrOOUaspzZa3weUW2qZC
twrePIIm0duEvo30TjHPw/JuTMRRn7BdAqqpKRaC8CLW4TPwJewlq2FFu2ZYaPgO
C2bq18uVdVePpfyilnUHwxnHnz5B3qCplh4rb+KK4I4vT5Kq65FICefJyyYirO4X
ocbKkBQv8AlweE3ICelPHHdU0wiFBtzYL5uHqaUJ7ocWbrgiRXbHFlv/kgPjt1AS
qixOesaUUhqmDcJU9jvrEvIfm6a1DjeEY70l1nmt+gJZVpUX0YJBshWF/L+ktWeU
LG8udDaBNTfThUrEmBDOLjhd9FNYWxLhjRAv9itMEYxCyW/HHDH8YorGrEpVXJCq
yI4slpKm/+bRkECgvf0d3gQSBTqCchRVSszeqNDLA8gsCYQC42ovirh+9kRZr5i9
B1B4aEAvE5kmgg3DQzJxexviI5UT0R2cN0UR7+twehrmINwdBgvAITsjufJaSrkj
`pragma protect end_protected

  // ---------------------------------------------------------------------------
  /**
    * Sets the Tag field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address that needs to be updated.
    * @param tag Tag settings corresponding to the address.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags must be invalidated from the cacheline correpsonding to this address.
    * If is_invalid is set to 1, tag, tag_update and is_clean values passed to the API will be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state must be set to clean, and 
    * when set to 0, indicates that Tag state must be set to dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing Tags
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_tag( addr_t addr,
                               bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               bit tag_update[],
                               bit is_invalid,
                               bit is_clean,
                               bit record_to_fsdb = 1);
  
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the Tag filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store Tag settings.
    * This method must be called only when the cacheline corresponding to this address exists in the cache.
    * @param addr The address whose information needs to be retreived.
    * @param tag Tag setting corresponding to this cacheline.
    * @param tag_update TagUpdate settings to indicate which entries in the 'tag' array are valid.
    * @param is_invalid Tag State setting, which when set indicates that Tags are not present in the cacheline, and the Tag state is Invalid.
    * If is_invalid is set to 1, tag, tag_update and is_clean values returned by the API must be ignored.
    * @param is_clean Tag State setting, which when set to 1 indicates that Tag state is clean, 
    * and when set to 0, indicates that Tag state is dirty. 
    * This setting is applicable only when is_invalid is set to zero.
    * @param tag_str Tag setting corresponding to this cacheline as string.
    * 
    * @return Returns 1 if the operation is successful, that is, storing Tags 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_tag( addr_t addr,
                               output bit[(`SVT_AXI_NUM_BITS_IN_TAG-1):0] tag[],
                               output bit tag_update[],
                               output bit is_invalid,
                               output bit is_clean,
                               output string tag_str); 


  
  // ---------------------------------------------------------------------------
  /**
    * API to get poison_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_poison_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * API to get tag_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_tag_enabled();

  // ---------------------------------------------------------------------------
  /**
    * API to get partial_cache_states_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_partial_cache_states_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the poison field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address that needs to be updated.
    * @param poison poison settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing poison
   *  is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_poison( addr_t addr,
                                  bit poison[],
                                  bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the poison filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store poison settings.
    * @param addr The address whose information needs to be retreived.
    * @param poison Poison setting corresponding to this address.
    * @param poison_str Poison setting corresponding to this address as string.
    * 
    *
    * @return Returns 1 if the operation is successful, that is, storing poison 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_poison( addr_t addr,
                                  output bit poison[],
                                  output string poison_str);

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DGCqdgSubLbdXyp7JzCp9Qy4VBaRcqXI7VUKvDMHXu3w4nKuVYLOe9TZ3Vw1/3Lr
RUb94C69+CfEeJ2dtLtaN3iEufUT1ezlteucecTDyj3WBLcKn4mlhuMGy0Vb9bhh
/yeOZnW6wKTdQnn/cMTs9pMcLcEM0krxAtVXuE78TeE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1217      )
WsL48NZDm2/G5BBWAf4AxSzn9tWw3wEQcWyPBRSqrgU9v0iWtvrLxqCKO98ziXhk
KXlwljxCH5NHljeu9H1a008OnUH26lR8GeoypGmdEJ/Hz6KMgAyQHb6y3rVI5p0f
qHC3eAN99ux4S3LQlckdQZVxwUjhCPknlKq+Bg90W+CYmGIJ9qu6+nqM9jK71A6g
AayGg6nxRV3RpsEaycTARCHua/y90vUrM4uS3YDwsfGQLiqqajY4YquEQgMa7wes
4oPZ+9bW1nX+HYNCm56CqEFAZZgnFBcG7UBFbYdopZJrnBGAFFsHvUvlJNlgiWY4
SLalAYucFzGgmyVXJGRu5AZAY4L5xvZYLbQE/bcrpiqopgCNkr0ZsGhsfdbELlGr
IApGnj+dDyYv8NzwjpFvQebMJugLTS1XJbCgyFmQKOV1iWvVz8fpexDS8ncb9FDK
qyTu8n1JDiIt8QXRkaX9H0mwHQ4SKY/m7vI6giyhqQBLg1C04q1TLjiw4yQbkJQc
IbpN0l6bIPOGTBcucNBeZP5OxWKiPpwxcgy8D6JI9Hk=
`pragma protect end_protected
  
  // ---------------------------------------------------------------------------
  /**
    * API to get data_check_enable flag of the cache. Must be used after build phase.
    */
  extern function bit is_data_check_enabled();
  
  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address that needs to be updated.
    * @param data_check data_check settings corresponding to the address.
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit set_data_check( addr_t addr,
                                      bit data_check[],
                                      bit record_to_fsdb = 1);

  // ---------------------------------------------------------------------------
  /**
    * Sets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * 
    * @param record_to_fsdb Indicates to record the cache operation into
    *        FSDB for debugging. Default is on
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit set_data_check_passed( addr_t addr,
                                             bit data_check_passed[],
                                             bit record_to_fsdb = 1);
  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check filed corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings.
    * @param addr The address whose information needs to be retreived.
    * @param data_check Data_check setting corresponding to this address.
    * @param data_check Data_check setting corresponding to this address as string.
    *
    * @return Returns 1 if the operation is successful, that is, storing data_check 
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    */
  extern function bit get_data_check( addr_t addr,
                                      output bit data_check[],
                                      output string data_check_str);

  
  // ---------------------------------------------------------------------------
  /**
    * Gets the data_check_passed field corresponding to this address. Must be used after build phase.
    * Valid only when cache is enabled to store data_check settings. 
    * @param addr The address that needs to be updated.
    * @param data_check_passed data_check_passed settings corresponding to the address.
    *        For each of the data bytes and corresponding data_check value, 
    *        this field indicates whether the parity check has passed or not.
    * @param data_check_passed_str data_check_passed settings corresponding to the address as string.   
    * @return Returns 1 if the operation is successful, that is, storing data_check
    * is enabled and there is a corresponding entry in cache, otherwise returns 0.
    * 
    */
  extern function bit get_data_check_passed( addr_t addr,
                                             output bit data_check_passed[],
                                             output string data_check_passed_str);

  // ---------------------------------------------------------------------------
  /**
   * This method allows the user to get an index in the cache which may either
   * be allocated for a cache line, or not allocated. If user specifies the
   * values of arguments is_unique and is_clean as -1, then an index is returned
   * where no cache line has been allocated. If user specifies the values of
   * arguments is_unique and is_clean as 0 or 1, index is returned where a cache
   * line is allocated, and the cache line state is as specified. The returned
   * index is between values specified by low_index and high_index.
   *
   * @param is_unique The shared status of the cache line which needs to be 
   * retreived.
   * A value of 1 indicates that  the cache line must not be shared 
   * with other caches. 
   * A value of 0 indicates that the cache line could be shared. 
   * A value of -1 indicates that the shared status of the cache line could 
   * be in any state.
   *
   * @param is_clean The clean status of the cache line that needs to be
   * retreived. 
   * A value of 1 indicates that the cache line must be updated
   * relative to main memory. 
   * A value of 0 indicates that the cache line must not be
   * updated with respect to main memory. 
   * A value of -1 indicates that the clean status of the cache line could 
   * be in any state.
   * 
   * @param low_index The first index at which the operation is to be done. 
   *
   * @param high_index The last index at which the operation is to be done. 
   *
   * @return Returns a positive integer if the operation is successful, 
   * that is, a cache line satisfying the requirements is found, 
   * otherwise returns -1.
   */
  extern virtual function int get_any_index(
                                int is_unique,
                                int is_clean,
                                int low_index,
                                int high_index        
                              );
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /**
    * Loads the cache based on the contents of the file.
    * Each line of the file represents a cache line.
    * Each line should have the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file.
    *
    * @return Returns 1 if the cache was successfully loaded, else returns 0.
    */
  extern virtual function bit load_cache(string filename);
  // ---------------------------------------------------------------------------
  /**
    * Dumps the contents of the into a file.
    * Each line of the file represents a cache line.
    * Each line has the following format:
    * <index> <addr> <data> <shared status> <clean status> <age> 
    *
    * @param filename The full path to the file into which the contents of the
    * cache are to be dumped.
    *
    * @return Returns 1 if the cache was successfully saved, else returns 0.
    */
  extern virtual function bit save_cache(string filename);

  /** @endcond */
  // ---------------------------------------------------------------------------
  /** 
   * Get matched tagged address of cache lines with is_unique, is_clean settings
   * @param is_unique is_unique setting that is required to match for the cache lines.
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param is_clean is_clean setting that is required to match for the cache lines
   * - When set to a value >= 1: considered as 1
   * - When set to a value <= -1: considered as don't care
   * .
   * @param matched_tagged_addr queue of tagged addresses with matched is_uquie, is_clean settings
   * @return Returns 1 if there are any cache lines found with matching input arguments
   */
  extern virtual function bit get_tagged_addresses_for_matched_cache_state(input int is_unique,
                                                                           input int is_clean,
                                                                           output    addr_t matched_tagged_addr[$]);
  
  // ---------------------------------------------------------------------------
  /**
   * Clears the contents of the cache.
   */
  extern virtual function void invalidate_all();

  // ---------------------------------------------------------------------------
  /**
   * Returns the class name for the object.
   */
  extern virtual function string get_mcd_class_name();

  // ---------------------------------------------------------------------------
  /**
   * Returns the cacheline stored in the specified address. 
   * If there is no such cacheline a null is returned
   */
  extern virtual function svt_axi_cache_line get_cache_line(addr_t addr);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM display routine to display the memory contents */
  extern virtual function void do_print(uvm_printer printer);

  /** Extend the UVM copy routine to compare the memory contents */
  extern virtual function void do_copy(uvm_object  rhs);

  /** Extend the UVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM display routine to display the memory contents */
  extern virtual function void do_print(ovm_printer printer);

  /** Extend the OVM copy routine to compare the memory contents */
  extern virtual function void do_copy(ovm_object  rhs);

  /** Extend the OVM compare routine to compare the memory contents */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);

`else
  // ---------------------------------------------------------------------------
  /** Override the default VMM allocate implementation */
  extern virtual function vmm_data do_allocate();

  // ---------------------------------------------------------------------------
  /** Enable the VMM compare hook method */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated 'copy'
   * routine.
   * 
   * @param to Destination class for teh copy operation
   */
  extern function void svt_axi_cache_copy_hook(vmm_data to = null);

  // ---------------------------------------------------------------------------
  /**
   * Hook called by the VMM shorthand macro after performing the automated
   * 'compare' routine.
   *
   * @param to vmm_data object to be compared against.
   * 
   * @param diff String indicating the differences between this and to.
   */
  extern virtual function bit svt_axi_cache_compare_hook(vmm_data to, output string diff);

  // ---------------------------------------------------------------------------
  /**
   * Hook called after the automated display routine finishes.  This is extended by
   * this class to format a display of the memory contents.
   *
   * @param prefix Prefix appended to the display
   */
  extern virtual function string svt_shorthand_psdisplay_hook(string prefix);
`endif

  /** Added to support the svt_shorthand_psdisplay method */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);

  /** Added t support the svt_shorthand_psdisplay_method*/
  extern virtual function svt_pattern allocate_pattern();
 
  /** @cond PRIVATE */
  /** Gets the address aligned to cache line size */
  extern function addr_t get_aligned_addr(addr_t addr);
  /** @endcond */
  
  //----------------------------------------------------------------------------
  /**
   * Sets the 'pa_writer' required for writing the cache data into FSDB.
   * Also this function records the meta data required for cache visualization
   * in Protocol Analyzer. 
   *
   * @param pa_writer handle to 'SVT_XML_WRITER'
   */
   extern function void set_pa_writer(svt_xml_writer pa_writer);

  //----------------------------------------------------------------------------
  /**
   * Sets the transaction uid for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_uid(string uid);
  
  //----------------------------------------------------------------------------
  /**
   * Sets the transaction type for cache operation
   * To support cache operation to transaction relationship 
   */
   extern function void set_transaction_type(string xact_type);

  //----------------------------------------------------------------------------
   /** Indicates if the cache line is in partial dirty state 
   *  @param addr Input address
   *  @param is_aligned_addr Indicates if the input address passed is already aligned to cache line size 
   */
  extern virtual function bit is_partial_dirty_line(input addr_t addr, input bit is_aligned_addr = 1);

  //--------------------------------------------------------------------------------
   /** Indicates if the cache line is in empty state
    * This API will return a value 1, when the cache line is in UCE state  i.e. both when is_unique and is_clean are set to 1
    * but none of the data bytes are valid.
    * @param addr Input address
    */
  extern function bit is_line_empty(input addr_t addr);
// ======================================================================
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
l9LwRBOUUkxgp/3lhNoAD15BEpPjnLddVnpxdkayiCQL6RjStTpx1PGG5ldvurfO
K1BcqFGsS3+JeKd85n+k3+gtmOdP/PnXck6pOmR/NdN5H8JNfcfxWWP6xw2uq/z0
9fG/8YD6kHox2vQhG3UabyzRqTXht0FNZ4yDcUXPRRQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4193      )
tgwR1KBkrVVo6e4Xp/GFV2rTAxl5D/aEOFW8y5gZKsAKTcRgfGARqKsFw+5Y18Do
H52Sh/tsWMcurxh6Es6uDOw/JRCUdDR7yMjkOn9KCDa1k/X1mJLV7OSjNXzMpe4B
IBRvZJ3Pb0Fj64ozxqmfMCmM6Y9RIs6d7oJZ6wrvAunbgJiC5JzS9ppzSxl/F1CD
S522JSIflmx3aTrEzZTzJX1bTHh0alsIsDuw1OeR/r0NRT7dEvpgNJnfumPVZlwk
Msc1p0Px7e6oqqbeZES987nV1ApZ2YrWvzdcL7D/f4EW1kILPZg5lNEp8N8iwVGl
ihhC8nOP2x/QXf6AmuaNVAGJQpvf5884X3w5yqQ/hDaQbrD1MfKwX5ZLtjjw5Ekf
5aBpHWV1DVNCvq/axBTaLhUKwIuAOtMgV9GQcuhjeVEhXsWONeIRWbhR0B4CnUEt
/2ApbBv4q6RGrzEzS/NZs4VAcGl5I88ItoLds2p9bj0FOwtoB5piAOMdApA+F3qJ
cdNULzn9h7gcAyRsZ/ZvrTN8/sLfYEfwBWQaImy+pNLGtG9n4ClW6lGbQ7ea2mFf
fltiToI/Gx2NSCeA+FLNJqnFvz0APGEkBqtIKaIZUPl0TgNmMw9AJSibNGtkAEfP
BfFNr2Uv3j5tUuDj40I+5QvfGqRoGiT0X7lzBsOgdT0gd3kYV6RLnoofTb98gRpy
z/jGO4Qeq4tlXZfrZy+OoIEw70m5ndCZDaZpO5R03ybQei9P8CcAg9UnLEV0/Zcv
LW4VL1bxB/Lru/nGyrki9VTojEX8ZaCJZCfXmFOytAJJTrkzqDmYNgdXvYfvf72z
ej4fEifliIf9UbzUY/PRO0oeELSwV8ElLsP/hNemkLJkK1Smtnmvj1F6uH2/H535
BRF+d8b8YzejrhfJyI4IoN9TnD8fbUAUQGmxI7aO4lrtihCJto6oAazKpLPVozUv
ut2YXBVIpUxS/MGmZwX9lZlv4z/c67chskYJ5Nk0RnBdtLL95guQfdRbIjcEYgzD
Y0yKnD/+VIyD767aCqPYVvYB0nO/3xVKSmzysGihAmTKFOCceFn28kT3iW7YvMmz
6ZBgpulbhkANbhMIyNLHYth4rYJeCkSaP9oDJZG6Qt9AKDqYrbnmlL+d0MmDJcUg
E5fJbK+4mAhwJJWUoF3xZohEFhObp3WIv9pURyTnmnZpJagASHWcRhjb2IlNKVL+
/m1Yot1bwraTL7IRA+0DYKRNDPBDwfnXhq618hMd/sLGFHrAw3f+praX+bQThP8M
VAwUWEv2l6MaahdBWuAd3jixodIu1lh7fkaSAUX2KFMsW/6q8Om640IryyUMwfoe
GBPOj3jHdK/EH2Xyv8k9yOO8AsNgjv3X+mNhE2SKXKtRrY+O3w4+JtGRlJ6ziI3E
8+g++OuLElxhpwrMBZvBWyniT3LlCNgJpenacGGonvDUvKiN217rVJt5Qskg2AzU
XEx+4xXg1Pq5qhsAyJbx7m2k04tOH7yyTuAGlQj4RF/UWYgdRFTaxvB8sHIFLm/3
0XEf5BUco6iZOmMTh1dPFEitKlbjp2tgxuFIhbENRorxo6KWJvgOVkyTOt+Jfdga
OymwwA58nztzfB+O276IOqtByH0cZOclCt+ybd+ZUOdxXO6XGLWTpHZh0j103InR
Q7rIns6P2Ot8k1KinDxMLWtFbER8f6bg2FVvjxjXemamGdGIz8G3VuNSzBBcedUT
2zaDNd+UayNFKE4qDkvmwwJg3uXE9g3zRgh5AlAkHztppeqkPG0YwETn5lpDf1h2
UqF8y2NotfCUIGflP53HSqILJmdCeXp7Bo2RvVeJPsfD2pcyVnHCJksLXpfLGj9U
EMUx8kh2Z/fMhzQ6t3dBFgW4cYrVmQq/1lvoWV6DBJS/QgQBVZllBygK0FSuE+cM
nLtuVK8W+Yf2FBGEnw92DeQxOynRit08McAKSL5cqACUxJjvty8jS7Yi10otgKgo
tOGCe44gECBDfxcqdSfd9ASnizGAguk8rofl88c7Laa3Rdy0ZWdhdQWTqyZpjBEs
ZecCkFLmzDoNPpF2HLSJ1iO0iHyWilKZstDtMhkCEIToNP9OTIq/OT1yXvIm3uCK
zE6eTcf/+jI44HqVkRLOep2CxpjWkR0Ya5PhBSUQeQx0e4/1vt4fM2JawRkW1pxY
s6pG2ZpBQOcb6h18v3wXE89SlH6ZjzCQjvpMMattEQpqVZwxCxg+76xPj5GbF/AV
1XtllmUx2/cSgrqMNVvup5Fv6rKRCEAlRs1/OEZMbltK3oLngWSE1/msvaw57UAO
lUPNmYM5u0tklpjjS1n74YxZTElEcfAYQpBWflXB59DJ9I858897NnjnBRGfDK0w
3awctIRr3c3EBP1vRlgsktIZQEoYpidtD6ijOVtXv8ATF8Q4Gku9bn2anjzJXbFL
ETcxPohOy8V5wL2fpZxmLcLRLolWTe9kt4ojeNeEogLQBzlcCaCpQbiw64aVl/y+
8i/jnWJivaUc0Bnt4xkTeQwjH8YSEoSD9munoRYe9/gD/nK9aUjaTlK2lTICWZII
cooQu18cBlv4n2Cs/0LZJbFkFNLag/qGVXi3WQShD6oncmGskL1ClcJvyn2hgvrp
+BPSinwDQ7SDgGdDFzf8uCKmBrkiUxgld15HADvaHBLMXTxCs6+JoNPqfKQa/JgS
imStP39fJ37dqyho8UgrO9WrQaO3IgLi5ym3RyQLAPJ5YgSBDzsQTMEr4ZbgOxMi
AlpGDBhsoGyuTNaPSz8/+w7sYGON87pE/Ib3n+a3mpknD8GnolvRL/rxv31qnRHU
T3akclQePva0wa8EHQGS/JXXIRsSB+mWyPkLg81Fw130cvQUZwTjbLVsF7nmAR0G
l0Ylst75GFKMgJw2WpIqRzSaFllubG0EwqcVDAwAQQax8J7hcNz41CbrGJo6OJ3V
RkqkoW8FF2YzTQBrJkOhdc+PGL7wGgISmgqJOx4qk+qfINOs5OH8FuZRq1P4ssng
uoDNGC44ic+rXJQgWH2EOKdNv4WZBRFh0Rz4QKk3bP4nZSQLSms49efIHs89o8jW
aaEeTSspMk+EZ8Y/InXvvJE1hmB439/sZRKTRcF2Wtox1dvI4hh26CuFPdHMiuO/
OjH8H+IioH0lqvyR9VWvdRrYh7xMvUt0EXwKPo8bu1wZvOzmCcy5Yf1RK6i/yIZL
TQXGGtacPwzErzqiDrSA62ovsaEY/UDwG4uTDxQFHPu4APYwyRR9TIwoMrMUTkD3
F4t278+K8a8j6gMHueUoXRI1Kv0/Sc3m1Yk4qOQ6oBGuoXPpEdyQDHSfaisglWpU
QhQf6ful5dpU8DAEuGqebyp6yinsWZomfyS9avSO0gobUWvRbv+XvzLyQzCpKB6V
hNvPLiLPV416WWJfbRV8rwkq9FE97l9/4c2xKU6WXbbC8thm0wuQ6HT7rHtBRp6p
QcLLaRIKaRpyywrYXjqTWanvdmdQ2PogZKsevLcuLUIV2y8NGCmNBTJ9i5cwa/2L
cxozsRPY3MLCk1oYsYgJjzh89bPynoH6dVhsmwgME6dfv+yK2tqn+24e7zpTGl/v
RZ+gNKQiuR66oxMHMC0enJWcoAyfa7KO41XwajnVlIGyxBfkQOxjYFlJWgSzkcrI
ANjw3XExo9RDJAMm9eKSPhvU9VlPr1dcxvKPQC326PdKRPsZbQW6smHfS+xLzXJx
IAnu9ioFmERLs2GkcDuzsZwUY9mxn2TshM6MXflSnohw6Mfv1sERbDCVGOC4YkSS
9HFDhZ/tcP/4q/cGIeFaQEKkPBP29sy5SXHy0H5WvCXQYxRHs+o4gPMPq72rALLt
bekqhXom9GyWON7bmKw8yoS3x0AODKrZ+QdMHv0yD4CF0eXV+Qj4E03u1mwZq5RS
SKhaPZNOdUAZca+tn/yXP1rsQl+4KhtWvCRK9pTAd3BgIF/Fh5W7CRjm8gqhdyAv
CI4yaZlqapyR1ee1wug4Tg==
`pragma protect end_protected

// ----------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GcZDujq5ryL12Kwr/erumOhh4i4ui7V6hdRrWnzpUNY2di5XMv8Xfy5X6eW8ynQa
ACMMWMic8ekprWN276sH0dcJcHVnPpJ55uMtGS8PFbXEwF+E+4u9EhXBJYi5jgrZ
G3zSdezGBcrZ20d2CtCHatHPqUcLUxODBzJGujV7FtQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4424      )
9MHujof7GcfzjPjRuo5mgXKIEapLm8kgf1UnyBbXt7YxEZRW/Gi3chsj41oP0/vv
M7X1pozoodKi+Nw4iwUQsGpIaAimmleNf1J6p2WNNqWm9OhxHVDfD8z1bLAs89lN
Q4sv/CzeCbcqJJpQ3rkNVnqJYgYIX+WnVmiGhnVcOaHjvspSaj2///raILZvkPlB
jRfajTjF7lHdKgySWvWz3x/TEsZ1BqV64ERdU5Q8sKZDIzeGUBuC8IAPvF9GGzs/
/sjJW0PhozNxQdWlbsr7XMJB3sPX+hZJ3Ebujwx3D74d8W0djAFE3CW8mhZNLtp6
`pragma protect end_protected

`ifdef SVT_UVM_TECHNOLOGY
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
li5r4BZUwwR4LWErwompnoLkF3KOSckllm3sEXLA6U6YrwHNt/Q264GMEmi/PRvc
pkB53Oe2bqnCQsCYBsAd5gZjXm5o1WcwCzqYzsFt6karAudDFWPlhso2trW3c7Id
WCy5luEbDNe0c2zU7MrlsRpLRUfKpp2eMrH0csjjU5c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6633      )
xVhREfIF7y3BjGc8pZtgolnST9GtPft7OrnYLuMDtJLJlUm3e2+gKYSmazfMNuH/
4xG8/j5gKl2v6JBouJUm/lxUIbln0N9kxm/BxOB/jKn2RXMPYxBfCjqJjJ1Hlk/S
eBUY6pckbpIYtprHU4DVbWEgb1nGluR/ucZK1edod+bxJOmaUKYC4jfRy3kizPDk
mBkLnXej17a3oS/PYuJWRaxRYXSf+t75cm+yOrMRlEA8CYgkBM1SQcezvcYsqXzb
mPmnS4N+jGJC9KPcOU4DcD5QWCWJvhlasBVv5rhiC6AXr3quMv000pp1BJtm+pXN
U8DBEsni0HHvfAmFxEBmY1VPaITiKQB/nN2wKTAskj6Uxz9ZhfgtLPoR8SLe7q79
Ol+AzvRiVI/kE/gScmbCQ3Z0wVVeKFuv7GvKSA1fVYJ4nN1+MxANGyesoYfu9JE7
u5ERGyuYZmkq9du1/5Vrh6vcTDwYvyRt8JsGcHkZZqEb8MAcuQizz04BAKC+H3ls
eIYHIidxxeGuN61JggsZpVbHRtpxtQ5CIcvTzwt/1JfmzIEdQKs220lXEWfznFab
CWkwVmYW1Rr3Yq3dP+2Mu05/8TYnGitI8MAj4N3sfpMIJ6Q3AG8yCbyy4ZYQ/280
lsDcWfvPilrZzLm0YtCGgFtgLzJ2chqgRhGr3YOeJWTTBDYKG9NxZMCCE5zxL/GE
5tPihKTnx2x/pV1az1A0AYm6tCYo05QzQIJX6W54ei7OV2XXil+RWOJx3mBM+/b2
e0UcWG44nUm1EbwpKDy4XNJojFG2bNGwc4/VVQXmEhAsSEPReP2BOfwdelmxpXiP
r1PLD5LO8XTyFycfPo8XThOME9T4PkgXFkcI4BaS/+P+xLpKUXGN3bYW6E8bTsyg
Arhxed2MG8UoB3wfgjFtWeaWuXyXk9EXGdUMDGMGufq4VLj9YGM3myCkf6aRoPB0
1Icr5/KESXfU+c5N6QAQJ9wQ3xCVoE++jT4KYT0kaML//BggQMTXaeD+AAyBs1nX
RbPhwC3V5e0EWYiIcJPv8S6y3tRA7qC5ljn9n5/lwl9udgnT7yUr+hTB8kJRdm6a
9VHkgIf7T9524BZMk8i+5sakxmJatTdnMU33+yRJtkkfxDWgol8mQG2tJPELw7Y1
+/U6Qjd5GXu2mHuO+VfQdGwyORmrVZD0+AB8JBmkG0ULtBU3VnFSsjEMlkLVfZ/y
l3q5N7XuLE/uHhPRYEXEon914ww4iEFlKoEZVrchr/P//8cvn86lhtXnr/dC//QS
Jochy9gSx3WMsr/xWx8o+Mn2u/DMeaI/5vM6/ewVpQgF82OOOCNXotsv+ffR+Cvp
Is1QB8Pnqg5qGj52N+FRNBEhBpvmeHTTsK1C9wimsn6oYbRMrUdFkC0nIEd73/X1
qJ9Ghz4vZf7Q3s8hhkmskTa/F60ak/WA7lAgSqXgVJ8UqE0+RK/WgaCwel7rWZJJ
AvThYUfx5XaANrKK5L7pRPCjEaszM7Rv1VM1r47PespXbIX9W/1tkJ1y/u7SH4PE
TgVU622amKQ/P2ZffFGZUO1P6yAZi3kAn5BPZjYRJII2Y74JQ0iwjd3T02v63R+w
8z/hR6mFGecPNtrtYdHx+DP00FRkutOb0RUMMl+QeUnhxzObNsxd6XC98pnishLg
rUuvvUwgXOrn1iQ9vRy2tXnsuQfyHdkY+NLjym0IYGWF9NEjW9Jz+3CL0JzP9MM6
a4Kd04fTDwXs3VKYCDUXIkg7CNRNm28/I6uOFKy/8JIkY0u9zr8Sv3xgrnpar8PU
KuTZrEROCbP7f6nPxcAvAgaZZpn8mGsUgAcFn+z6/6ovOJ7W6phZe6TqJAZ+Abpx
SGGreenQwt9HSZKjJoz2RgECWNk5MzLw0wpcK0n4giCUVwOnEnKpXTBJe2MNxz0N
vN4oSFGM2V0xphfkOtK0ry7LiU0jNO5cRnRwKril1/4LE4enR7bzRsjwNmT79zC8
zyIOaf+fdfGrGhBTBAQBUXPC/z36Cr/n5gUO41LLD/i6NbdEZj88sRnzjT6SsMs1
bZJ043HzOG1dwnSX8d1VEHBDxVgvq1qzI4MJbCvIXJE95LOKJr9zmgQHXOSF5OpM
NZs9pSJk82ux//2zxTKH4cwE8sgZo11p/O2JgDV5UGyrcJLZWyKdL36LMQ+dBGLr
RMWiachfBOuQJxlRtq8AwmuHvGfSYB/MabHHUI+3CB3aCqI3D9SBFYjgwD8OedbM
/RW9DqSJFJugC85ftQPleUHdHbOdds+5+0EQMOmxsjyVjdKP3e5p6TNMO4zXCKYj
msKUXJ5/STgH738hlAhOzRpJNbNkJmz0sC2P2KOpmt/3w9gUVOIHLbTd5S9PffMf
kAJEQeJyhZO06Ugx/51kWVDeR3AtDZ7QnKc/iR0bE84HMpJ43kb4bp0NOR7Cxk3u
z40oBnlEi34OPJ4MmByGOI8f6V8iGG/c129YaayIneqdvJDqrV3SR3B82x3WTgpj
ZnF2gmKKpX0HOwKsTmBYK3TW2NLIBiDmPo8YlrPE6sclHk3NkEOu4+PaGbQofu5A
nV3PNH52iMR7dYlPnfl+A69j55ISGC7CdYtlp0O9iSa+7r7O9jxi/zTCvgZNJ3MQ
dlPFqZ/UeMqExIlr3PlhBw3qob8mfwUay5C0o1FtNhNi6jsfXbNXuwZXUe3ml1kE
Fmi2us8AOdXrsyraW/AmUT2M4N/v3I/qrG6OeC7FMZryTlATAJodI8FCkqRvMHqh
HeKG/+asPhA/BwPJw9FNO+37Rlwnfj3tweH3HTv6c2v/PLgvgUznUaJ2LA6M7cDx
ZIRCnxMKSgrN2b4/F8P1ElAymSLKr3ep7nyoMZ/w8OGFdA2NkV9c4TocUg6wO+xq
m9jPJ+P1vEHDTedyWWmQyuB3vyzpN4/l8+NrwZgivfzHS9fafWAvlNj//AQJIJJj
qHm1f2t9rNSv0qlCEJjQwg==
`pragma protect end_protected    
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ijZbQxRW2viZoEjl1+CwcGZyJOMd5DtqnAY8I+0lk3KIHtO7J88wu+uKNFJZRIG0
8dSI5rR4ZAaB3+e1tOiwX6r6t3ocaMs/bVjlzEtkg0m2AYMRGoJYrCY8Pr/yVR2z
cvTfvpUwiy3PTSfTK3/nwEqrXo6WSktXydihyEvwI+E=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6849      )
Hzp10FCaUfiVQTQgGAVUjtq4qgL+ZxWGzWRGqp+YRv57/qjCN4IFGYo88jMVyu0p
vmXy8BbJ/+8pHOR5NW4zrkIte3hW6ubOA+V1I3hGGDaHGN0e1s7Nspgy58onP834
0/Hpvvh1x5TzRW011zQqjryE94v9lROATmC7SFKKz/m7Dw+z0J8pHdPQ/v7tMYv+
Yx6LqXIkBinrylFBiyc1N2d/NchaFtPIdsQwYnIIRpGBcNyRciZGYvYOroDyPQw9
m2oEhNF4OChsjOnf+7MaFl7ZMtSE9VybMH8d5sb2neM=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ISg+CZHrBlulHp+oXbB8A7WDUfVlZc+BBoGsPJwb8RlpSPu2byGsqVcn50mmErYI
c7EC0U+X3hhVWMg0ysWS82z9xa2T21nqWWx/8Li9UkSXwTktsnGifAElYaq8t3yd
ErZJqIfw97Eb/Ei7HAA79cYRpc1ibdxK0mOQHcgVa0o=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7345      )
XkxNJoqh4rgaQrmixYxbDU8YqP83dz6vVCWikUvkjXGtUA1HFyKf7iw2+jYZvoJx
wHPoJHb4OQERPrLTwYFSmesjb3z3hqA66Y+I1SYE6NWR5g6c4Xlm8+zTusHhEDv4
EieWuvtD57Ao+rnuSJd0yLp2nFIUhBf5fnsUkqq/BHEN550tos3StsRE4Z29b5zL
4HBDWYUPK7FRWCBjJuEpNljosbKI9jhgGpTkH82LpHbba266RB7piuib8CKcGzR/
n6vfgj20PJOq+jfLGUBWw59tOyN3bMql6Tz1LH8ccyW6tzKsjY+Ppq2luBSRU/y6
K8XTIW+bqPKsk1kBIm75K72h0YQufnz52ypKdkttw/F950vc/0kCOo720214PC1r
EWo2WQz8NCE51yURATU+gZ1yiCgGEs8yr5J1DiO63+YhTpPto1zL7Fg2OSx6LFLL
4QGILMBjUzWKjKinj6zCUmAnlHbH+OPcxwYRCyeEFfX1xkHCxgMAc8e8cbOIMBTW
3Lh21VvWlYuCbrpcQfMxbSvZU2+7KYhGRT0MvxpIF3UmWCS7vjRIlRA6rHwttNnM
cA+0HRhlr5KOdSxTP97WR8dIwfleVH8U0o1e/Wf5cb7XAdEK+wDEHvh1kwFBpDEx
9TgL8F2/lJ8NIHFxOTPkhjWLSxZ0Ot5WyfoJkppg+Dc=
`pragma protect end_protected    

`elsif SVT_OVM_TECHNOLOGY
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IiiS/oN3UQe9UXxASxfEpts+iJmNGbpA8JqdqeYpTyzIw/qjK6No75dFgbM/UZ1H
J3rNfSEyqnfdUouP6cBIdHXMMr5MzdtjA4dDVqBuZBBq5PhcG+E/0jKI0Z7ESghS
ekM5TvZ2BVHDALz9aGaav707Mct1APh+IfuR2FGqhD8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 9979      )
Cq4AZC2LjtjE5NqewobDCmb60huPzvMCKjSVyLaPsG2guKQmuI5ZDG9V0AH/JhSe
h/zlbpsRE8IjN8JIgazRHBqctvRKhG90oh/Zd4d70EjTmh96Z5vnvJBWeTsqV+bi
PDKdNgJFepQRc1XRZZPGF+G/gIqTsShdRpxGmrhn0LiwwnFq6FQmR21OhnAhcuuq
KzhZ1YZsM3JxZ4JpG+MaQdPhxz/1PDeRSL9wv0U9vyTn4K+Jx9iUJm53UFQV19AD
VHh2MHuyq3nynh8+LRtFQuGUliz8x5bE8cTnSADsVd9QGz+sb8mIKnGq2mA4hL13
+LLADSY5t50emp5tLKsGVA0qX8XYEP5VypRNcncCOZ/U6EjH7D7+YFTEKhjGCUcV
3NWhv15uDtfX687eXnkuhoLO9O8AhfG92TmuF7/WKnwcnEPdAT9UHM+vjirqL7Bc
lEMvPa9pNdGt18jRsEeLT5IJcBl+FWT4JHnKgFTiMIb8M9+5ALtrEDrzOvAuFlGP
Tnmcjzb4y756hM9CRwISf6LSdK8lyAksI70n/FIJORXSCxFPRwrUSqvxYPEaI2lA
WDELZqI58Urctmf9gxRp5KofcrrvtUQ5P9wLfqXjwHUxylbYufjvpNMj703T+l/J
vnK9qJy7lJwC6JFdhmL5UNhs2bG3fKErLpR9xMD5H21ZSuUXJlSWmKh4oXWqiuB8
NNB4iKveY2zJ+dcuQ1F+hVEfE4lWjSIUZaPYaZ+U4Vt6G4xFaERqIRKZV2itVI0/
v4AfpKCC+RFKSSPnF28rnVroyjKQUu6NyzLZKWlCOV2hbJ5lirFEup7udb+uHQ7m
pGmyvgRZVY4H/tvK0vis/q8lk01RatSZ/3c6HXSd59zvWj7SmIG8wj5XBdTlSaxy
WRug8szgHGNBi29WH2ekE3jO3xL/IM4mXTEOeAb2p8lYlbZy2J4UB02D7tD04Gc0
SAVjiLlAFmWyXLuW7RASbssNzS/J/iLZjdxTJIKMrRa3NclLG2DtYfx/3MN00G3c
b6lgDaKc7xMpPcrfHCGVtFS1kZtGGFzpplXn8ByPoSYZmLmQ4qmD1owuua6J4ciY
iGmWpLzDwgT0lEj08YOrYddyteFojjr1pmupNikEOEUN33tawzhz6oKt4v+BFs9b
puauecGfkNWRbnVifNjjZsdB7B3K0BF+hcLYoyGToAmOOj0gcwNioMlncWzgIVoz
6I5DxwNji1nVaD3HkZP0jd8PRiLSDZWHbvAjbjcOJ/HhSybumeoe3iMdpoK/Ijne
+SLruCmAYSrD/80XiOrjMq36+HjJ4Jku87NUowHcrOF8evA9qAOPP4g1G92R3uIu
AdyVHVYc5RvO6umzVllEDrfCNv/InnxehnUYZfVsEU1AMvb8UI/GHBJTwo4grySc
B2Q3UlMDj39xaqym8Bj+BEOoJ+yR1h2yfQ2xJVbqLa9ieMUho1dhv0Bt4UVCJ55F
aGBfO5pURKietXkI6YWDAQDMxgH4m/x/b3pte9YDg6ji/diO5eI2snORiTfQBYBJ
LIKT2UOcHIB3TmjHdEG3gRlEABhBi1mFtdFM/oU/UTk5mA2R++xRunEUY2mSfPti
WQIb+KiFgOZTL3XIKefFbGP0F8B1BSBc7s3YUbjAKx1qLSUSTEMEVOW10LD6pLo7
Q92SszWWSRPMWgI/HcdngLZAL2sL4HeyfXA1iK8PNibwIId4EJ2OkRliUMLKLRGA
vMbOovU1KNMEHL+tLkXZvHMad0mnF9huJE+23pVSzkd+gm68GZQhxvFcahwF6kgI
Ivf98jCAaGxnXJh3VuiTQKl14OFTWUYDy2gk15LGVWFo8jHaPLObVChTiz1oYyvD
3iQVi71d9bSoGQaHEgIx+oYU7zFWH5bhEqvZTHoLlNScpr9q0rmFjHN7qKcFAxuk
1/0vnyq27gKSq6rWEWRHsLzEegPHmOKRbxW5qKS1JG+LDuWHYtw8Au4/gUJKOwVc
SSU6sAqIwGM008zBb8EElU2dfzecIcPbkZkNw7ErvWeVrtqdUxeACuPzL9uiuTXg
cOOp0D0P4D2t3ero5jHx8BCTOyXRPpeil9IJiBPbH0mTbnlE3yJ55usHySuCnQyX
uaCzTY3o+Vt+JPGS6lVnnoHMZHFFcVD7bAalF2ojdYTzHbNcf2nug9HpbgaHrBEX
0TLTvzRo6zsFqhIbu4qJC3WOhjHS0IvamfrzjioJn3D3H5V7ihjgdim8B0Sx43XG
bMmK5NSG2d5NsahfnPNiNwtV9tvi4Au3Qfce+wvdLxnA11gsJLbYzxSQBJr4xhq5
hdF0X+7LzUm+EfOrq2vagQJTpXTZ3OkHCqtdEI7ApTmLrXuQn2f15njiKcVKaXZ5
xqop4iqUxpIYxDIbhMSCZbEAhz1n2lOe9CKRxJWXcAv0zztfmzDFPEekt7onhhb1
ahJvSAn2k16tVwYz7I6v4R3jDVT65RfHfHpck1Gw8tlViRZ3ET5wFXELV9QppE+d
2O9dbbjx0r4lsoRlvSfecN57me2XGNfj2zHd+CS6LsZnGLyY3ypSH7DULUkBgxWB
JhZ4KMiXPQuBJDqI8fUBaRx8ZyyEnhqh8DTe+KtG+IUuFXyu5jIhai8elAJa6wsi
KC4XWOZgtpGbKGo15jyyc2O7aKUj4Oo93q93cqp8KKcHIhiy+ir/tQhZVzXtN15M
6+RSh+XWsR+vAWI+S9b3Vjw2236uXDJOibV6ueKSNgjTv9/sdCdV4OassLKlvJ1N
M99dtPEAsdCoteH+aSSnGbg6hjtpcMvZLohx4lzqqdLfgd+dSWn32LRbs1g9Sa3M
ToOHcEJKqaKyXiFtppy3Qv0n9yg/kjts5bNTva1tb3ydh3w5v4YK+4RKJtB0wjhJ
W4YuAVsDOq5/8f9yJRY2comFQIeRUjjhkoWXxs7jRhOEVRul/DIGfTWQi6KRjdPo
1r4vvZ5NV0uK3gU5vxLO352SJlGUVAqtBNbVCHJ1ZsOJXKSGFkaQvl5saH5RbyVq
k7mUlskuZlk2hvRZdWZBvH5m34zUoKmJf6g7dOfIPhfne8TL9OqlW3RkQighJ+tf
qf3yHt8vvQaLWreRtQhXoMcDZ4TCHlNWRXRnolJt0ulizuNUGyCCfhvESrC31zIk
iBiZfQBNB2HVuQuz4637sNMcbSVTmaXa3qoRP8Hdc0h27N2dmcNJozAn7TC9bU/U
ZvQt9I81u27bZ8dDKBtJu68REV7tl72/e5Ec2s2y/K043c6Mff9JpcXvZNpOQ/pp
lUkqawB6JgwpftCWkmZJdtBJVW13UF/RdKhLD2WSdg4De9wYPHUG74ZUtSPivIQD
+yGWvIQb/R86ZqpNAnnvqTEXBT+2EqExqrIhrP4Knp6NUKW8kAOi21HyMCHwX9SL
q0XYfhqAnDZXQB2qtzxDEOuTKa+K/QH4b1paj5S21V9wh6LNSb3fILjs/la9VS1d
+DAuDYXUpN/C2XXbiYo9S8QUmMEEJCEDA8nPnq/JZkcxEXWxxVtz6wsABOpusf4+
`pragma protect end_protected

`else
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RPRi2G5l1HfJx3jM5UTbPCHnFSDj4FY3jxqksCMZKPNTQyEMdVqeme2dERFUHgSX
8BPaPyn88tcpxw4qX/AIkDnOOgpXPOgKLugy8rqOYtKCWx39aH05UtODPA1MQ1Rg
/aixbVC2AIV/aoDWbVu2Lg71jZc2FQCjgtHUak7zKgI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 15152     )
YG8Z6dzn/pGnlw6RtSErJjKzUOtYoUbZYIK3Yat/cgjStDGNed6Gbu1ZtkjmVC7I
Zo4ofVMG9Qqo4Q2g+hWyUv3vuRbL2YVCdwzCOsp4cHtPlwK9tAz7pRJ0S0HNK+hE
PtXtSWgl5AyKwUjytOTtdEcl45RkPelU+vzNDR9yvufhQt+mXYX9UUKdchcr5w27
WhW5ZvGKtNOS/ttHjwSbml9fRQq5XZIJYh0kbxWSn1abjis6gF11nFuKhOWzJatG
hOEOxp6vWYWUsd8L9005e0Z+0vs7usi5RecDkJYghOEfghse/g8QEeRf937YwHj1
R++2o1R9T8VOt/2CadRQQnqpAohGixoqWGHqKO+h2XiRykjeFqpCqRO8jQz4Gr/a
oWZZ0SC8kO74CRR1yfr7gt5v9WHDyWSUAOYHWsNFiSjS3gaHZRQjYuPNcqwQek5M
xh9/kRkchecxyXdK+FrEr7WggPSl6bgVQNY1pMgtN3snt9R9gd3mzKaNeg+PeDN3
sK+qqs6NZiSldRetgUgWRqj0H7/kEsrrIQ6JvslXqbHUnm2lQT8s+DAQYO0yqTt0
K+cwjcTzzCGizjQEL+xeZ1bb9m0/567hzkm7CdgAskRqTaEQnppn9bGq0pWJEhHy
z0SOmY7ODjXVszz5DufRzsAJc9kGJimLp5G+PbI+SiFf7PAnxKTbXjZ0+mWOrEz/
QVZYYKgi+PZTwajatNW4OyWp17rMcggStvqkBCyrKO3M5HpxQgHNeEffPNepK29V
sWZ1v7wtZUmEi3tTIfp49waGTpTTpkR5Na2oV3JOxz8tV6dfooD1oHVL/edyJ/eT
5LetT0GuzrO72F+qXp87w8YXCdAroF+HOQpZkPwND7/V+HQDF6Dia+IjDF62YXHc
wSphug6X0wYKtd0yW+Jl53VQJgeAgBu5QNSDXhNCpyzvAjGPYTku4V1G8lAGB/lQ
oCk0JRyXuUakIqAoleveoRNWMeq0bKHrSB8vRYkilWG60/CMF/G+wzXhA9bbqkTc
Mvzg1qB/7ClxpdxWZcUMUmFHEW3ytaoBsTpPeL9SP8AjlraCv2xvXZM2LrE/QAIY
JTc90lc6ErhMZOC3LnETEL38qYqCKgyJ0Mue7GL2Z7Tqu3sw8r/hTjv0RAaHtUJP
0ocvSiX1xCDpVrS3OsjZYbBW12SePJy8775h+5cWzSO63LMXOiaEbtUAkscchW70
Q9C/TcLJnQSUKtilb9owRrpkW8RtK3hosYNyEff1RGH6xuP6INXIZV4lDxByqu7E
HLP0RZc1ltxD+Y1eJU35EuHGRTVI7X1qLzOQlauVMO9usc2M3syUU1iXgl8u5tnb
RyLWNheDnyhL6nIlmuGlR3gvBqYVEBX+CW4xIhZQalfcQogUI8G6JtgdkLdLMFAt
Fq8H1j6tRHtmitPZUeFcNOvB1LF6xrypiCkQm1A/plKGtZLdIkEv+YbI3kARQzh+
rjoqs1dKI0VRhalDPkV0CWfhO0LUAsq///IZJBKyD6eh5juLdKD/PiMcIIzZWj2L
WVskvhbTetIXbXJfwcRVyHeWzRn5Lhrl93bPyA1be33f5egvSAxEcjHEpx+pXv/c
MMF+A94JpunBliwWXJmjEWO6nohFRPz5u/SwsgTbB7aGEqQ/u5+s3z1TBEkcDDqR
HiyfYnsTvwul7ztp+AHK+k5D8zlQd7ENbMpfrLrCAQPuzTZzIkhAfBFd/FQHTpvP
/EeUl82wp3J1N2cMC1qsAXDe0axY+rh3QS3dUSYSWE+cTnAgtOTa/fIjafhOzN4/
cBPJ+zhweO9Hv1AufcVWl+DaHyWmkNQM5Vaer1TdegKPLBj2rEQMEtmzEdcnWIFF
CpBWMpBqp9lb2OxT4GTdAQFP/y2n76Tyu52ga+uhgSpesisDBY0hJkFFSy55OwWh
z6LGAzQYNzajz4FijGP5DzRAgFWxUnwFpMi1UCeyz5etm4bYwYCy2QMkdhR1N9nj
vryWE/e4hbNCNbZdKUpw8CeJF8RDN5pFeLw1sSxPTH/X6/ZbHkGpVW5RXqQj8a66
dQWPGYLB4+pvGu5ZEORUKFNLCZxu6k5Dvvgh/MKAQY/+QFW+eTtcQ3/K0F6CI7uJ
FtTYbBdIQqvwOA3tzSXyUyDIlvDVN/P4TuXtA6WpzG0Dk7WkLj35TF7+PC9tG2zQ
Fn1v4GR5yrq/ZeLWUEBJUrDia5ZV9LTEboV08lhB1xYxVRvbJ5WBdU8p+IAvJXnn
KRLjNYKaeVTHCGCu2Nbj/GRE3HpB0VB58FJOBO5Oz91Qf3xN9ddDM1PV7hliHGMV
8p6jVwC6G/JCcJu68xFPJKAc2B0mpJGvjyIFztkhh2EgEBrILgV9LObGtSNZaEOk
B9faPU1GQNMvtQe2c1MC8TgGJ60oaiqu6OF7bP96vmaBqrBZ3jdaI4YLZAN4ozfu
WjhgPVmoAaxv5yORnvtu+xU1LsxkXU++PnFTOz1UqoWE/lOkaz284eBcdVVhCKhr
Wz0Rrk2/Gczqa39ZqqkFKGCb+DQVsCUIBNfhYWRE1N124HkxtDGQJ1hK8e/COJOX
JOGEBl3PycYDQ8+7sInpOsmS7bUyc0ZRKcLk4DwFE7LOHTgjOFW+cKrlkClxSfzs
hU5ZizMj2PKJQFCYNd+ews454VNT84J5g1zPm+rv07LE4z7pon3n0gIYO/BNQRl6
8sYdZzrjRgeuommeKR8OOaXL5RMQT3T1zsLHKrbdEzJnBfvpSLRRsQ4nlxSuFr/A
qPnrUnckjN1SClF1mc33IBycKEAGmzvm6L8hIkGnSD33amjKgbPMwJOxIt4VqGji
lTYvkxvUtA7HbCNS3MqY0gRA3p42EdBJGDu+Njg+Hv7k3GCnD44zDdEfyh1rO+w5
N674bnxJHL+n21Z6Lj8JuK/g7/WYDPrebQkXhZAf3O2Ee/7iT76KMx1dRTtBARux
OabGPlE7csg+N3YPFscuIitU44eAXIMXdOyMAX9CDRjbkBjC94nNPT06MnRnz93q
wMt8g2uTGre1YlLMM8vrS1yFrfHJzvS9UyAuGt95d/g9ByibGJ3JswcH5kk0A9oN
i91buVqw/rUg1/zLsb7GKTcVwyJKqGCxr0v6gWQIyyX/0VUzy8mA+FAU8MRqpWjV
QiV9xEtE213mb2jzwdDlCbxcRzAs+1HD9Z11x527tzSbQxLL+7wLoM9VIh4WFpTR
dbssQQxZAOnmlxv2R0kVsSPODh6W0tnHQmymPmjkgLtFhKFlDt/1bu9abztUPO+j
nnKAoUbuTIZVhiT7ihRZgmixGIuM5URmIfluk/rQ7uQF/PrXjj0koOoG0+U3sT7C
7KeNrg0JWJVuS+oMdRJPbq8Zo+MTY03fq2Ya+c6hLbSsQLXknqNTXyd8jzC4rF7s
ZKzK0F5JA6CC0rXSol1UJtptQ5w3CKGwRWX+qRfE1t7uwvk/Vvwb8T9JbvJRBBtM
rhej/aZsQogJJst0kceOnoGHooN42TWS0YKNep04GM15tyySacUnVngF7NcRn2No
l16XK1yX9/Inj8fEbGxv6m1N5ZSjpeYU+oWgbU7AXjeC27kiM1tm2AWlzNW2I1dJ
XYTdXj5FnquCa8USCCcmvkaZDrPZKSgyJsmlmp3kMGEMuLzQ0p5/XN8g7XxahGtZ
5qH/zoZPQTLL1VIZxqG3s7KfPW9AOHquwCNCGGNWPgjh37aJHNd+HNVsUgoavVx8
RYh4mS2rrZcioTlZKr1uERIAPimMqKELuhucpmFOy8IZEmmjQlA963qzwuhni6Ii
6j0LmGmnzlauUFbLiiQKbA7UbS4HyxFy2g40VXDV+aruoq2mybPSGW48Ib9k/XcD
8n0l+0egPo8I2LCklcR6cUVlhDThJBCB1q4bOFt3DlkaoKDWtbiGOqBezHX8vj6p
KoDvJNeJySrjmopBym9mpm7/nWzFfrH3m1c3CAl6oBwfuNfdMx4LRblZjw523bOI
1RJmkvvY1OCeiC8m/hzVjbvCXGUwDRt1DMOR4QzyZgtrn3sDKXn1wbIqRCmKAG9W
VvhSECh0B7Px2g/46yxHaBzX8cYS9kE6MtmnmPcw7IF2qlanZcQcxVKqiKD8Pei1
9McxNpRfd+sPY/jn9hwqzXJW8EtPZZR7C+w9AtTV6RyW35DJRYl9x6o0PPyQFxSX
Ud+Ddv+uKAXjEc/ufEPBrohyVceUv18gPgaZSfhueTPIdc4GhD2Es1kbzxdy22ZP
ew+w7afJipHQEMS5AlhA9JHF//pK0Z4aBgsiUp7QVLflGseZTqkMz6dvWqxbjOoi
cW/LAWxzscjbZlqrJWuo7F3JIZRnQAdmNT3zIqMW+NY1qa4j21YmtI0MBzjpu8C6
h1/ns8ihYemuZlXKRa/TiZPxatYBskvgF+eracW4IQU3kqi3JwZWorr+UWg5Y+cJ
LJUovQZHMEwbu/jwdFcRLQZynCWKkMobkXVbVWY4NxAj42PpC7COoZUtcJ3kk7IA
n/bWW9/SbxjhN3ADdumz3E/j8j6t4+v6r4oE6bbkzTNKI5CCAHh4PPlCVjN68mJs
nrYTd/RfRaZmExGUfbxHtov4D5ZX3a1dIonpLKLJSHyRYwRgiIUJeIMLHCFeJTai
78Cx4Ogv9TSvrmCAJCErv8jKs80Je3scF08MLfk/6KQE+VBeN2FXJe5yTgfSprGR
pEHLvLgnqKc5+q86/cGD/g+wjQpWXcVNzNfgDbje2xkyGkvhJTszp8sK2b7FM9xH
YFhWZSB2O8ltZRYew27cC46vKk4irZV0T1WqhGGPsD5kH99g2oFxhJqZ4OcH02QS
Z+ZnnlaABlKcesIMGNxlGZocJjTyKEB3MSUjSv5PT/tJNIDj9wp5r/ExV6M2YYhT
J7dPMj58G6HzeEGcvR2w5i5+j/OlGQUppl9t4s4kxAhlfoI4TiImcWoLae6cYpE2
GoWJzN45kAT88Cm/fhRNfwdmp7R+WiItI/ZNXn79+8FGSmrBH/prPaNmm1y9IwhF
9BKq7/jOEq0u1g1u7hZitu6RpWgj3Wueiy+QNbk3Ac4ojFxa+5GQBodJ6zT/bPpA
ZVVS/I0QS0SkkPMR7g96mKUtKBT2+P11vHcO7lkGEKnDpbDJ5VZopsm95HJSgyaI
DGt9lsWdwgoPNeY3fi/k5CbXHpYM23s7eCtkIdpsNxwPeQ7yphv+ImvF1chSeaOq
hd1Y7jCtysP0uA7JZfoZUspFBgSPFgTHtiZgl5TUSt3q4UdGu9hT/ofAzgDGw1M+
i9mzpgZklYIRR0CeOTl7dUf3S0THEZPOWu0Z9IakxABLyWnY+7T3AQm+klre2qli
cyJ6bmnbonPK+XWBrAPjluz0SxZVATdIofAvny08q+yY7ZPg560RIuPqxQuOZspm
586ox0Wz7ZE/DByxJoSHStmyTFgMrwpbxojkr7JybWzaahemf686Newntl1wxFok
Eb1Ow2CoOzCg/1u0fQ/a3+Bqhos25wwoMCZdjGJsM9IrwqAokVE7cFb1phr2WZ22
1aIwHV6sFTfsXQc5pmVd5i2Vt5+M4kCC++LKAzFVoAhuddm3yiZlAMSreqgiJOtn
wTlD/WvWlIgYx3J2PBgpCUZ9jTAvamxvCU1LsseGeNPZQxQRNXRaSS3TQ000rBYX
29nmcMO3UjOH2O4D+O1UX2XDvh6bnZCeyJojtMi8eBeTeoSo2jM8iSuuq4ayXgtG
zuLkv7PwPzDa+TW8zYe2TOXf0nBsHgKoO4MqY+RiNTDmyapv280I5AaspXnriRL5
JmfYMFU5PolWIU3S4EU4uWJrDSC+hsMW88AOvvhmCHkldTcnpqCPgvSLoLBuLFeQ
D9HKqGpBlwxZeI+WhXSr8N0Xd/8MwIJAvYyXRkTBJVLylmVFdetBknTMd94IZ09O
1WbgN79N75wIr8bD6F1sr5PEN82VpFGHIdceH+MwC2mKWMZYOrsuKRQ3wj2QPCNU
VhY1CB1F00aunsFcCkDxomQicOctHxaH3doFxchOpp1drZASaSJCKR9HATBtMieD
t5z39RMA7nXiFWxCpwo1wPjnNM+LEzb9TyUCVGRnepGlD/YWxrz4tfj5qRLYgau5
TJjEq/ZnFtENvKho/DUqqHsfEimXCim5bMVZ1H+I4bRetfZHN7W5yXme4+yoIg/P
sbar21/D9iBGMpY0YGsI03N2NY91UsCWgVQgU8kVSv+6lxhm6GPi4DR8YdwbpWhq
2jjQ1FwMa9QFyOKu5/yHfGmxQOshKp9NK1djE1Y6RuAwVtDM77kW5OQF+Ya6aoZw
TYl10IsD7lRHKAz3viW5uNOSHxT7pn/mMlY5l+yBqy5nXyBhBcHnEqwX9Iu7t8Bc
8PfZnCwq1UmOGDF1Fb6ofc2eOYrpPDFX4SGY2IqZkMmDino5bk23Sx7uvDV/inRP
ZepDvTlGXTJpL4uUalUHDy9jT1m7fY4+SDpZh169f6r5nn0/TjBBoXZTbzpaWdHd
90WOqmw2huVdI8+KY8os+m774jIyTB0YXvcuK4sWIc5/PXOvsCq9NM2+BEKr8KOu
3sG2aoVdUltojEa9kmfUxLNEoBq7+oZvaj/8anM24wgUF8a/BZcBR6/7IqL7rthP
ryNQU59SEm67Jumf75PLfMWdJpXD/65Vo0s+s3pugHMAKU7ZYDYbWOgaqZZAv0DG
YEBbQBTtJzvME2wrdpCvLdfm21OzODcStTMYKf2Qm0by+9rXpvGjZus31CckxHVz
nSCCcJbpkGS6+R9E8vrw83qHrLd2afbktVa00QafsB6u/yxWKDLZPuFGCVe51HTh
cy+GKSlPo9aaYzZ9DclI8NI5t/+iJ7zUBSgJOREd7Zi4QyqxcrQP4PVMniG0sjfn
eFOxvDBQqxqIHlzg4sfdYf1c52NWljYBN13VWN3MG7PQbeMYOnOZysvVcs5JgC6i
`pragma protect end_protected
`endif

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
d4z6yqEBTOfjy0UULvxCjEXIvUCdD2FrTiXH0vmyp8XAU/5lXRDI2wCP1Msi3BNY
QpRhNa2eHETUGLHAs8CF8MWVr2/j+4HFJg+eezvqxXrT6tSAc7RDbcQr8cfRd9rp
77s7kLVPssPJJdv+ZDAhtii+AQLRXkjOCu/ixPhBGZk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 104599    )
NZibmWU+RdZ4oOg3Oof0ud3Df2bngXxA+B2FDxbF6z9Wpv2EfM7s56ZvKsOYJPex
dAr95Io1qzYIfXNFX+nBtnjccN7P59nN7AuSOfmJVQkDzfjS6aWfN0mrNWL8oi9V
TSPdDWq2koq4pkudSkd3SWnSzAo5N5pHrmazxtGymcN0ehu3nECIO6yztPngPUh6
yC/KgTwc66ldJ5iYYYactPmHcq01b67Y1EJe13FK/7uvxTMm+Iiw4nohbWhb5Mv1
dZlY+CJhkeOcuhP6YvmwsVFSLuUIMJxXIVdErI5Fbhdu05pIYMuFlJ9x2jTRhlHU
xzaWJMRB5kr/HehwizZAIYskCM3EgMLyYeuG3nHwzCsFqwWzFWZDYfwQVGws+pX9
9oe+QsET2KYTiiuD4lliaXm4JYz92Sulvs7kZ3UFrmNUQ/9Plxyk2XvyMfCYQvQv
3xQ4bxuLV7Pv4xBGfaHPGS1pZTjb1FIBp7k8E8Amt9LG4GAgPPMPyNCERnEJWyxD
pF9GYbt1TcsaefD8wgSRWTgMl1QeumHJNyiCnUQ7CHHs7N8X2asaCW7E/g8VtQFo
kA+99GIkg5rrt9IT5DExJsklOktqya3hG7Iu9wQDJR2yRBqHg0pYcSspRy2+hRTe
QlqCAaxXS9r7kQh8LR63bGpgWmj+dHN6f88ZSSrb2VKz0jLEoaKAE7iauWtH5owf
b74jggj/kcuSql1UFqh//HfSFaUZ0Cjo4TKGOmuZTXOmpOo7RksLerIcxJmaLjSq
3I3wkwCzYta55XEJ9o9LgH159ofVkIJtY55r3p8k2J8VJejCBW8rw20amIBNxdaA
BEDyaGuqhizOSoUCwT6namnGLKwEHBCEzK4GLp1JzvH2DgTQ2y5GcQNwpcYKFaRf
7RDccq0aKllnEo18GMq56e9gKaXPY2lR/3uy37uVphoK9eVBf1Q5XXoI+an4qEMR
kGtAnTjrfomFtsIbnaMcflI5/+ZJ5aj0srn8iaCxBnpAxwFFuMMFgUxKzYyrY2LW
xqtUT+PW71Es9x0aK1nUmI7zpz2I7FLll734x8fSsjOY14TUhYFgWsJgLe8CrFd3
Tw/8EbG42Ks0pkVufFBNhDRr9S6nbzxYVjAl29zBz7Zt+qDxz5n26SsxICS0qdVq
U3jHdqdw5YStiEYXh90FBFbZuRSj9MikLpVJb2QI92XlD/TyvzqSmDLXDO5BRl3y
vnBfum2h5NzmdN2f/inOGikMyJZ/XNQryCnZigATR71UPXSJq5vQuo/5QXEK18VZ
bVu6mb63348gEihWQyd/nOqbIC7WkuwTiVQg1Iu6gFSlo6deC6B/bLW4UDywW6b4
Xx+LgD7M6WcTM3iUWOcp9btC6EvfJXqsNc0Pgd3EG8wGdzNXRgu2El8GyBbDCZof
u5OFT3hQcxn0GxiYzyilr2AMnbuwfgavGQRSuWao06xFtXxP1+oIrQW2HuXr5IJp
VOSYErLwdkYWJDZIuq/a+odf/Izj3JTWVKdCSzdOx3rU/0GMlDJoL2wfx+SYbU9z
vrX3/mZKQlNPSDBjHAm/deOrx1uKxCJ24ezCPn28tZTFbqehhBLSU/PG2qJiPT+w
69IgFOQChhhEp7HX7G8vgRXTp8WXx3FAUyvo+kkvfE3wpaHU5s1Ism6aWSY2OkiC
zMvbNh9ToBoWzwGNsbCTJSoQSjiOpLwzm+WpGzxlQXg9EXQGTMAY+MjDT8ZbqWKL
udWWHBQYn5eWpzglIcotxQrt+gCvCMIoa2P+D3D+6+eWr6VXi1t6yVQ92wvW4YY8
dJeFs0rnDyoq2d2/djDfinT+pMfsi44viSEaQdGKy4acqtEjdq4zZtOPlfUoXN8+
yqoIYGVKxl2ss6BICwAhk8oVr1iIBby0sdDNEMTQ6Hymt6mJkoLNQgUC6VJknksV
/POSFr+WR0uHiRRIdQvDdzcGVHa0C/4+EFXvB8iYaCHIL1jSh73G/lRVGbgzN9lL
3g76y9EF/XpI2Zo4a1XrQ4jdtvfL922Z5Q6KB9f1DPyEgzLFqadIyeD1nA+mMc9z
4OHiPocQ7C9HBQf8qg8ykcRDvTM9ycALeXkWrmRiifyIFgMdf3KYOSwWxd1z1a9O
Ky8glmwh+TkUK2XeBloP24h25BY0LKSYFj/mrG7qUOWjEubPN54a64f0ZPdfkZNV
7He/NkHVqOs+tiPdM7KA3OXu5IrnI/9+BC0RRf8Coma5fTwZP1uNXckFPCsrn7lp
Li57dyBmTWnzbKlAO/HUcDh0DXdp/8keGbWNAcQbPN5PDD6iNQ94xyWepLUPj78n
I1Q4B9NUT/TLXZIcK6+M2/UiUsvNL42NKCfF4UTe8GpMQYP0SxBYQt9zOjjK8U1I
fWqCEyW3JH8H/mKXUjABZtc6i86hgbJQ2+jwSsEy8YOJ/L6LVV5sdkOxrTh2Xx8H
Ziuee0/CLMExtX0gcBdmroqKuU9oO4i8wZeBDKTEA0Vf2uVR/JH7AjnFKGfM2yDP
w15QkF1623WaHJTYdvwGwPNEDmbh5mxEtU0gXnwg/nlLWOTW1ObKoz26mIiYnko4
vjm2lDEPrixP5EdkAt0j0Fm6u7GYy6vNtfAMs1YSkYbsEo3m/xEMxU869qFA79rS
E/QXOSMdQqS7hwWbLhF5fFftJLv1fKmdUbC609XpAJnRlpNfce2THxvATJori7PD
r+LhkFEgvAFqjtuKJCdXjFRgm19loDVoGkXrQlr9cJMUJ29H1B6d8dzjRkwyK0w0
+7xpj1CLPV2abxLlRkVUFqp4kuUKjA7aNdZksili34mwBpdVFeGTWCK8R/EitsG4
ZcKG4sfP0MxPXBwLUwRo5E5IJ07mKtJ+I56lSEBAgb6deqL9UWAlAZdgTJ88iQXR
eYy7IPLCrSqNRbfZkIRL87xhBdd/Y0qwlZQkH7Hmqy9FGECCWdk8O+hwq3GY6jD7
GWIeyF3r6U7tcZBhLdgh86dGDHvEpqDw0/E3VX2qhTsQ2ogCkcA2a9yA292YdtlX
/+wchfXlLvVZajWviWMS40pUrDzPmjV9c0ff4gGOScfWuzkTEDAeUZWkDzSI8a8z
3si9ul4kKMCGHpjXjla9UL1pjn7X7QgNFBJHEsY46VzV1QuTl2Pg86Z5IvfrRBMd
0Py5qH5MkhVfLDUB9ZfoxuV6hzjz/x9Jl9ZI+DSqr47+s+bAX7yIwPV0tls3wzcW
t1EOmxz/ZJq4L/sbCN0W+0GDNzLtErgBH5RCP61MS745FCpfTn3dJM1wxGdOaRWy
C7KA5pi4xyRGGon1Aiq7j+B3PW7V2NAUY/yPT39V7L7cYrSVIvKzJea2t2VvKZt0
Mmj2nJhE964Fee9YCxG+RpdaR34QqPujU86Zp24ymBDjlnUtLMln6zj+uZKAEU1k
sbXKV1I5LxnenGL6ftEOa89QH4piXxm3NxwijTpVVQv325THzvpweMukcfBJuLkE
xkws8yCVOi6oYq2hXqDwreqlnvlD5mRFsG/WRdMeEHHRXFpNpBj2smzfAMUC5Vzi
mxPk3ctwUUAN38tFE1htdwxhf+EvxJXLSKDYmYPsa+rOuRTqlSz6dUVb+mHSTpX8
HPW8oD5wWYp+aCc/SRq4vsQ9qBwEnGpUH68WMlcLrJpics2a+E+6fw69/Ypqcw6s
eoOlYBnnUKQ8vobrxD/ar6RdGh1MhvSXqErDJUSIlU3bTOrW119EFoIpJNwrxc8W
PX+MGaHROWHGR7oERAa6daVEsCDGdf6Wh5mNXO5gXru5LHs/APFncJcq9stgpvnz
W13ba0QRxr+Zrv8JOt+VcQShhf/v0MCYqoBuka/36HywixNR4uRye19oRVVctiCc
GtCYpkm7robu/FDVPGwNuQ18HicMuPejI956LwXGVk1BcCHjcfbDT/bZOjobW8EN
FVmaDHgxysfWCjKl92tPPZPTgTUnf6iUAwjEoRKUf1gDBeRGw3hmXVFriDDuOsCi
B+5ucX8uYNcEsUG+OF8gGSkXPB2N/ybYfEHYvLvuz8GEGRDRs2eersmzEDC4I0Xb
LhROs0LgkVgc5DBDPDSKfArOX3e7sHZf0qe3ghx585JxKHbfhmaQMxLvOGVCcXs3
JgH+q1wmQMpulALXi8cfL48vhvZTSd3Qj+BOafOcN+P466RozuZdT/cA9yk5w9Ew
KJhy9UlMkywDE9VXfdOVwriT32qYpo56KW8LD3p52o8StsNc8rhCIO2gOos/nFtX
hZ+TravnpR8Vj2NI9/ulPH2O0G+kg8eMTMnW7UC1+n1Z8cEqaxOOGFXDm0LLML0f
q0+uWhnQVb/lQc65NtUe06/zC+hSD+tYiOoG15p0fsKDYt8YjWppxYfduxoaJtnu
SQ90FugvhC1NcnFecIK0Cj5ZW7PO8lc2RG8yXLhlPIKTz35uM+8guXuF/iqOQMc5
9u/qEpx0JwoqUcRtVqCi1SN1SejcbPGjGimCz+YrYrBDx13K0vkq4+2YiQnvm5ER
LvzXFFt4BtBwWk3rbutc/VOzMAyj7E18Uw287Fgcfa6wHuNFH2STYHwgsAiL30wZ
jhwrWLp2s6IBjTppTZvOB1TYB7Oy+v9mpJgIZKI0qi15wyVSjAlIbWGi2Uit5YBv
eMItQrbmE8GhUtbkPv+Oky7+kDC8c3K9wLdPxC0HHeDiGoDz7NKFDRNwgvK8r6dX
1+DHfY+lc000Y3eIwyxISkgkqCorm2LS8b4YrYCo1LTkWXJSOD3HYVafaAhhO8Ey
xbRhWriA/V+cnO4UDh0tAsd3UH3nknbS/k6uIlMAnssZ+yzrycEY1IiMFgr+db9Z
PhU0EevknGHBUyrC3DYS6qc8EhtYfv0/KUD2V1qrwKwNX837bqzBibdVyfyXpGR5
oIJH7MiMZQdexeFd/mmDsX1pMzK/rxmQuQd0Rx6dN5EIS4rcBWXa//cGlFzIdSYf
LBwIA6v6+Rx8GaOhmI08SFTuNmWcLIbi3aGET6bi8FRjY5bDymCAvmfzsN0U9VDp
dbo/YRiq4smZ2p0fqlt/cl5T0kWjXlETp/NOpy+E6gWp53UhibwAEq0aQkUIQTyL
hcnhlMpixDwymQUm59n0fXG/IGaDYdgoAdM15KDjBd4rQqShP0MXHc3Id2ApTCIj
YSv4ugwWwXexdk8ACFeNxt4yljvrk1q2kirMcgiQ/7geaANZp0YClu0zirpc66o2
+4Yjy5CtPkEFQ/Mrc1YoVykXRtY9PeB9SrmVstFeftLAXqeAMaldr7fqpaE4fIxJ
jw+MRU3IJWOUX/yBnPNDGv5kbYgaCRHUGx6BPyaDA2GhloiMSiiN0diNLOqZ2iCW
v0V2KcyL0X+Nm+KYMiMPHov/zXUKruh/kX32HgYlIrguacai4iqRG59kRxiCYST2
vwvGmPyV8zGW+q/ELcI0HwNej7FAmP4FeAtx+c223u9K9Y3WdShe7P9+Cn+S6k8b
WQG1IGm+cXIDyAWe5TAXL+IkjXwPP9gzcfxBjz6zR96y5mXDOD3SSqpoE38Vs9XS
sh2ZVGLopBYczcm4ESLmIwsj84rp5qw7ZprH56/JxtDBvYR81Zw4U0c8gd8S+1OQ
JhQKgkLjPtt3MKxZrHF6EqcZbU1opytXJJlKIDLkiD0CRQxK/N1H+NwT6OTuxWaR
5wOmcaw/M9d6y+V7eJM8SkRS7S+cCH5ulPsiicm+/KT8f4y0XSYG3+AXDOVfJWY1
bXD+n1ieBJZgrmjsLrX6FI9lU3yTA2vZkD0BQE5+LcAlIaT7TZFrvKHqE2FvoVzB
RDGvVyt9bopDNns8QpcvbLWZIqDKQxSw84f5S1zb7iad0oL48FzmLVqzvHpyiRWa
kSJ7FG0wrSqkAf6mJQUoniAHMIRNMRXuYtqWfDjtrXO/hdw5nlcNxzXUTWJEt6K6
9ELLuINbRfcKP3cCM4ER8WQDwa9JJkcgXbeuPTRt9Q62DqVNfUQ2w3bv/wuVRj/w
g40SqQwvFuoHrcSgxRztzYIl+lq8eJr4KH9t/xPDHe8ieVe4RX1iNgexhaq07H7h
y+zPeMMgeWOmgNSCasBERQv78UzrNCxzBZk6TYsL/nWXwYZf0nyp1oG5KTq/VE0e
Ksj5jCqg8e8giXZocDHG5+JFOTABEm53BTv46jZFaYRYa10UZwM2fR6I/2WEcomN
qsc6v4EPjiwxRLMvYtrMGJjyvPAans8QjL3hUt0xhSlOq7xpfiSMg2qv6VktfGMo
C8nTR1MiPYXWBNeHvI8PRqRE00Uo3M3E24TqDD3pMKW9Rmt7G1iCtzh4wUaarVMQ
atP602cFmDWffL5rs9h+L2IHntv6RiqMHm6DpJyJPSpPpuhHW26rpPI+APSsCDED
ix/p8UedDC1ZSv+Q+ugfDYXlwlQ+gD5Du5vzrJC3SQaR2zSg39PRlf4QNXpwOcsB
YnyA1Is1c7yzchRixWEL3iLY6/bhN0xdYAxs932cMUBCYdEA/Sc1rzkqlAmwkanD
hXRPAYk4+rxAGwcKhydNtxoGRZViP5Brc30CiTAWo9OJ/EnEetQXbYAjxgu0fDE9
MAZjfAK5fL9iQz3r4WHGMKvxDd7SuZiGRdw1YtpbGIN46NhnoVokFDBE0SR3WrwO
wqrtoUtdcjOXk5fQpJHi6bCjoeh74m4xVTf3CbQEEUm6j+5crc6WRbe2Z84h97Ug
A0cnW7EMOER9kW8YpAABNKsa7wOOtNziJITVF8AwerjT/38f/CzemrE+iv20bYRG
cQzIzKk4kzrNfjpIYdyx33L1EPluKwyYzgqQ+pZIRJJUjf14RthDT284Zl64I5jg
aFDRwskwbgiSsU1tRIjsPljsqqneJXrC0Q+ltsWwJFGPpjBDeDxjCDowgiQhioiV
QBhN7Q4BuGnZIWb/aEPXEohghbjKN12m9+Y2w6blQYU3lHHMWnmODjjchFo0uLBQ
ZJRzqIR0RmS2nrT9uwNxhX9tH1p/+YqeOllDMHWDPskS1SrnvPB890CStqdyPThB
vUBiABcCzeozoSVibUo9tlp55M4PidhqKlYI+mXvZDPUCB/lRJbFsSPas+dltI1Z
ZiiWK2SApKqlAGVmKGYcq6kQ47FIWGeqCwksTsbLecOJ0yHVIbFIV32RW2hJIMI7
FmyyQ+Ny4O48H8sJd+wDkC3ZiWTM21+Ik65/pxHElT0bISmiFeR4FHgGq9vgGSmO
frYLe8NHNMw/yYJ8yCxCSkUjE53CNNubxWSkzXRTXFQ0GnYzXN5kAfLi+nZdUnGy
LscrS3Iln1nQVtjYA2cn/tOWI2WtBF/iSXOUnUI6FCsnY4nRwZcK3GXUoErfHbXd
Np6VdlPf+Yp4jX5c6keCH46K6hDHhwC673bc+RVqoLaigGhJpzEGw9+Zp+O3ChD/
fwBXbSOAws50lxFbbtK7TQJRAkD9JmWg0zwMGQO1sWl6EzUw8ch/nMg/v/5Nx+bL
ADSCYl6HUANPZ9wuJl50f7J9itxLp1bPKkVvERbLODpoLAYImjmjV2Cmnf4zR10Y
367JXpslbLk3JUBvS/HqUq5WpM0/wSs/xNt5c1aUK+m6jNIUT/aHqjUquW+WRXD4
OlRi+FbL/0HQyf8bkDOMbIiPzq7N+Gfa+ZWtQWF3VIKsDRG6M1eK9UA/nwYh1l4/
929vX30FDPTB5+dJMq+lkebCExFhMBS92g7dFmdhOUasDljW8wFcXWuJCoPW9ZeB
DHQeIpv6EWsM3NKL608+fuKK7U3+5byHSuL4v4/ICUKc1hPj/KeVKAF1sB9QebuU
NdxBlSscBIqPHWTFHi8vic6lBy7BKCU8YyRB1/XopuNjNv6irbycRE1O4XsWOm0O
gQGD/Q77xLTKKQdgz8t6zS7+mXo9Zl9mXQMcaNx3KehFeIJ/VZipaFxAc7SVje6t
oAwTanPExT9TYHG4CnSRbPwedvEhdB98Mss/gb/Rotn0AmQNi3zIjAh7dRr3C/1C
rBDhvOSOn1/X5hqMYDLjL7xuT/5+qXzZLenZhP9iAGigTwauU1sHcUYL+5GMcMii
W9KyEyX30hhjhd6KKKiOr5E9TjEaEe6FfG0vecWzcptVIRe9P3Y5QRLbi0HhhIhP
diZdwdjhA79R73OHrkV1iPpkoHFATsU64FWxLmkSNxXdkkE+iIf7UmXjDMpspbQB
1BPiBMR6fx5MMNWUfKF1BUfjGPTpS73MOO8eAy733KVdksPayhlxy8921ghvQTdr
ZqpaBdXBmAzq1P0TKQ5CFaVOGPT1eBTuH4DFOejSjWkoToHT/t2w9yfKDbJrrKbn
5iSuoGuBvS005yT6zFUYrJ8bZeUyfbsmQZkb/mZTrZfT3/nxj210S5nLwVoLgyMU
meRAqAPXoJ0D9hYSqr1cw7cAJefxbrbYth7nPOPAuLbAbQb+M+mJoNcHljfBxyOq
opfu6Cxh3jsH1VeMoSHvFUNHd7qFroeWmjGIGJFWGamIkObre3Hv6gsEaxYr+PKe
0VVfbTZzjeaCtL4VdP/bROuqMTS1SHSx+unBfDjF58c3GRds4cux5DefHKHpi42U
zzbA7mEHqz0fUZCSXFN4uJiiQTx2zLD/zeToELeblbSA3cTx689FCQK6TCmgWphu
XJLc9omd2Wd7ZRNVwk9Ft/eWC+qcfFDct3mYX8zbxxRuMC8QqJACEuvcRwX45Ot/
2DXzNztx++V4NXzIUt3toHiKfD7Q7LZK6I2BVZWE217R7DjbrBy7O53651xEG2pQ
Lau4bMPUy3/l/qhrS5t+Ah/+atkiTsuetcOpzvulVuTeWrtJ2qWnPn6CiNEMoeF0
hq0367rm1g2eUvBDQDQi8XtvyyuQ4fY5zVekNhPKHA/88nmmMWmZmcc5TM4E6h/o
iELORMVXRWa36nUPEEzF9o1I+zLRrFRr46SrhYTDm3twzPtaAKDX193OrIxZ1Dox
HsAcZiNBwwnGvk9qn2Kzx73fy7Z5xNKFncKM1Vx/Oilh/Tl0XBPFzedw9SusSXXb
n2rCJFDXojzV/8rrAqmLPeoc4V/9a9m1FQwCDt+cpE6MDFijSNLhyFLLUM9cQvtV
XntCDKg3uQPmYJrZjXs649I+WZYxZPRVKKiwmENAP3patE2l3Clknkg9fubwkaJM
UX3R+t9X2fD34zkOxqZB9/y/xnMSWrqNdi7z81jIr+sdAZRlBA2QnfJUjDacRz6H
JqCcZunD/cmaQAtryeJ7bMTxBLW1dlxzBrOvaZn5457V318UxF87qpV5wa2KdMAr
VoetZkjXG2njYOX6/29QMdtDl76w1QTYQFLPJQq1KdXmLdntfywrvTV1sE90Bl61
32ZntbKSTag3MGnm9y51gZp6pI+2iRZuib69RdpW8Tlm3ODmHq6Kh+q6rbVBtRyX
wjPESAcDGrhrwK0pg0kYCxluQbzz5jLsfgCmneMoMELSM1vhVc/qBrqlrtDeZcYe
4YyQvzKCixHxcvKe1FFSkHJG2a4PuJYKvr/+NnAOhSVlZ2hAF30vcxhsdFk6h9UR
/FRPeixpMDd+/5BpvUbiJ70aCvr7vPA5ValWIKsiQoPIN216agnqI81VjvBan9NF
xuAuzx+gzdzGdBZpnn9RZqFZ4RdJUFf2gIRebL5Iz0VGqNg3Bt/bHc4jEGiGW7jS
YFjgAPRRYtK+Ao460HsEInqQa5H4jXeQWW7vBb32IVBOYsRdcL10i4EqpDds44/Q
Dy5mTXQLcZCKSWqztFnl3thzc/D/FLz+bS0Ob+yaC1cM1bwsSdAwx+t0LS9GRmNl
n+w7LDqvo2WWMeIiHUDmnSsm6jqx3eQcIfUf/O8SjyraOSgNA0WslEWtz+QuhvHe
aM1GNEzfZrH6tbPERFX39SaMtuW58oE+nPoCpR70gO5WYXzPa+PV6vgjgsF04Tpx
A/eLDakEBo71snZjIXzjHBEdZxKD77RTcxdYyPl0QX4qjrZ+Tm7ZxsFB2lu195nd
xyYvy39yMLvXa2mxytaMGHxSkGXxBqS8j4myUYJtfbwFBGKtYQaAMMv4cWREHa8X
x9Up6rT38Py1h7eGSjOuQDjhT27kapP6bLsPs9Xbu3c1rAdCdnlokGL0+VKU5G2O
tAXrHb5yFChG45wV4Crngo89Sx1EoU8pdcwSz6KF8aBaO2wMtf35wZfW8oLo8XMQ
DUxWTaLnwFMhm4HPeSak7j7ZQM3+p3uuimS1cKt0dhLmgv2ShAvHkF6ZMfTddx8J
Qz5dyEA3g14Lksfk9CPd6eblYw+Y8tdIKTVdMrOcijngcJ946XUw24vpeKJufmZZ
7p6kbfKtvC0PZDp3n9DJxWbVoLsq+zmKjJWBB44o8QKx+kwKy/gFK8B1sm3H7Liy
/YRCosXvcBp92VawIC8mQvO4nfRsovffwJxnGv22wTaHZbsxYmjvbftgLVpIYedf
hEJrw4Hn1Wrw3EYA82Oww2OuvuDJnEJGwQ0H6DtP4xitsOxioRWjIhmucnr0Ar4z
n1tOHmT1XzkynvTxbwF68E+BdrfX9tibt/lDXsCTvhrcvydVOmFi7lLSb2TdVRvq
d53FZsI55hth3MCQl48MkJDHIcHCNPlp9u4CmLLP9DxJDPLW6LJD4ftrBHxCADx4
0Ky8k4WGo0FeBhTFmqaD3YULAkd6sLl6tOu5WXF4PSFfiQMZOV1jG3/V/eb3a33V
P0JVTV9wNOnaFRMEdTGV7UMbKL2zGIDBLF2E8iaswspq5oHZ2+975Xhx7aslJThd
gPFfsI6UAQ+0enMXCmlewi8Wbz+yxuMlFCj+XnboAXbovIik4YkccHHPpsWzyZK2
oGwnLMWWmLEnW9tuwUhTmZhI+uqqZlpDWAfL7Ewm2J9jXS0O8j8mTsDZYnQR2Kxh
AeBCJYuahpHuj33kNsY/HqZND2fcZofCB3Sm3ksnseUwK5cn0uoNIgy9I1jvZnkh
uuGyxeF1TAH5vxYHNabVTpvguZHHdQGKZRI6C29LL9/0D7hI0LXANWdqaBJTAZ2p
ArDbcq/Z3CiZn8WIW07QKyIcSCZCse/Dw6qggCRcz5KJO3cPrZB2CQkdvW17+lLS
UoUIbusJRv9nl62wT2Wqgh7gf52yCntIggevgztswYjASLtVF+EUhYy3DP1v3oxl
DipFZDm3HAtr/UQj7YiZ1PaDq3HIVXeNAA+byxPW7P0QmwA8DftlaB4HH2dnU+pU
tsfC9UJ7I/3ppvP06SGiedJa3Wt/uOUP+tH9wXuz85iMxWphWXWLlg9Wg98jBJ6n
+ZpkSQn9TkUMcVeXTvhgjt6Q9C9X0BKdB/Ui2DAiT3Cb+PemNwYXJRXYN3e4ELk2
NzYf1RiD90mfOlYyqDo/nRkDOciAGedAj84EGih5kqVfmrUmXBhUS4VKISCkWme0
5HdqGD+a2Jj5B5plcnj4CChB+5+mHLnm6VHuNzBh4YyPTkSC8InTtxnjl/IYS4ta
gPovGIIHxPZGaf+/dWVdcC0ZfRW8iARPB8cYsVKd4E3SKx/bPwItrzCRhOvo82Ha
JzwsM0gOn1yYzMVj2yiHwhlLvKsqJ1y+L7FKniGbmWuk2M26WW5fDOSWpfMWNegf
TSaiCHogKrH9a6PDPdPO9SmmwBRnHS6MLhtptKv0kRvTJAj+0zCYN5DzdwHwQqxu
WlHauWr8BpTpLPsYYF0IPOjSWiCoFqwDEfo1AwXuvAkz7zqt5AEncF78NsKUGiII
eg5A+geVQuYGTzj/igGutMjWf2do2ILC7kNtmopLo8nvwh8g6+tL60ipTm4MfcA6
/umJeIPHB7tNzL0miVZanVi/lYYKYkCBWLnuVq+mLB0JkTkG/AaYeiZt+wD6JEnk
zhuYS4OBWLlAHs+ta9LB7d81w3b7XORaZBcyF26TzJwaR7R8WI/m1Ev2sejzMhAZ
1uzFz0515Ez+VOfFECFgzO67zD7+tkLD9whwTMiUcdQZuzriRraZL0ordPmFBOQl
mNc0XpeRbC/5y+meaF+15KtNXznaBG8dw+K4klaUePenZ5GykPXOodVe2BCre1/F
YbOnelXZzugAChbz++5SIQz2Zv0QTtV2gU/YaWag5qMAIDvkN7Fg0zwLgH8Ta0yw
RMV6bV/PYQZ1LEg4QJ8blaPswW7JYTfENv59LFGDJmZo7xjZ3iLNnFjYGw9GeguF
tSkN4N4Yq7Qpq3yw4L5cNCviFByNuP4TUZX1RuJAJ+Dt2un2sMkP0RdSbg5pSeYx
UpfFnY05XOyrwWl8T6bdOzJe+bCnRwVOvGUktZGX+BcDiP0A4v3y+gbtdiW9hCs4
6rLM8uvIO+ZjNtseWiIg6mVg0KqFg58FMnzRluhlgkMGS9TPHM3SxLrHoP/tcMQ4
oiecSMABbYs7phEwedc3t6rQ0wOjQlTr6wlo9bdgHLhr/5glhJ7V3fJ6JOQ8dRWC
05kW083Hq3n6Nl7IbflGAZyMOqNpB2zHIZ91xmcSg2WDCAufyGr0TPOZX7MaO0JH
8jFwvJBRNGqNaQo+cG34E256GarM9lKlm7tSibpirpum4Glsi/DEkrUTAK1I81S5
O++Q7T+TYz+InvVP74UltdyHqdHQblxDnirb5s9Gd8kyDx3mACbCgZlSdQFs303X
EG2OBkDfbQ+66aT6g94O4x91k3ZkRR+7q2B24Ln9xqevvJLcblT4fx67G1PUOqoL
KFZeCl7mJJo6ev+2gBSTnfE6apbaS5V7l32+b96ZRGNM/2zMuPAEVY90M+sN9I6m
nHEItNK67dpIsgrMeVWCdnpQ2dM7s+oUO5Mhb5EP/j0TGpSBtW2iagsJrxo82zbq
16RyzBdhVPvsIsMerHrJklglWLXOX5O4M0fxby9hJ4X2ESKOsM6ng5MVkLHuSzxw
Gpt0NocTvi19hpXHjrcER/nYcaMoRZ6CpwyeDp1u8pvoyRBExwsh6vjjxz5c2aSg
kHBNdhzKZEXEprs6mvjXhg9WZZrGZYSum3jAfm5oj/h7sO8ODoKXE49p5GwD3slX
mL7A/p5t5lw3nonnyJKe+J0aEVDpnB8CgBIkiDPItzSMAFuIK9mGSgnLX7ylNtmM
k3QdQlaaiY6TS1IK1qBV2VEhVW6uuDo84vXhtMt5+oM4D8SVzAkt3Gn406Kyu662
fM8Uo4XC5Lk0/uwiIaxiLAE3UX2sx12UJIZQ8FP8r8OiDJ6NM6CoTkJQ3OnnWWai
yFhPbp5oKjMU9epObim7EVcGomNgnpzrdo3R1wA7RbxHHVKT6AvwEez8zgxXAEfo
L32C05Ovg+b3eTsMWbujJ7SOhXfvOJH+gAuBgDv/PVgT6TM73flT9MPIOMs7RNvj
kqIAVu9REpW8DH3xZBuvV90k/9kiJoNTd4wVvxAD/W6Drui/l/Fq6eUWN5d3Ag9E
XrLpsBBn6MO1JsGlMY+5DQNIKWaJ/FvTp6c5nCQZkfzxk3S8pyR6HlGut9Qfa56O
IqVKbAWCqHVnES4Wap4dlyz2ftVUkxMeSRSXxsJpQVkZwPI/XBJvxLQ/s7E13IzR
6we0xLX7jH3Cg2wP1OBHHKo3TDr0q9CIzp2oTy8HSv4aG/Ha2OHZQkbHBum5TB5t
fC9J2RZdJppMVmTKerHTn16oPk7OtXGBO+hdwHsTLUvOjWFHuxNRjbNrf55ex5hJ
Bt9phRSs8G/oq0ZEaZMak57MSU4xcOw3EW9HjAnUuKjtcRo+XfqW9ZbTI1rNKSks
Fs54q+a7YO8npBFBrqZaR+3NgKRk4nhjo4ejJp9PwKG0VXflZVz8L6nU8dJNQlJJ
AU1RMBz43BfSHHQ4gZmstGfwpqFDINkKYQtS7T1P92ijE8Jcx+0qk0GM4/k6CTYe
7I7yN6/gn0Za295l1kw/y0TI0nVhFhsoqvQgE0LaZdz19g4dtAYkB1kD+wNg6oRk
L74eyFVlF2KRp4WqtIJKr1uBN5f3phhs06M/y3nbmNuBclvOYlhCozfb6vuHD9P8
pZPwZ6V/iHM8WIOMn8QlTKALwTQ2xxPejCGasfsAoS4T+Ww6Mr20Qg4W4Xm7l1r+
Q83erDZc+MuauEqVcw3WVRhp5qQPVf3QPdUxGSCdB9Kvkps2dnVlN9a/s26tvhkz
9kDdyoQgp9zTUmp/HwsUnu4FxsjQ0bIZxuGuftRH8cx8Xi4x5L0yQ8kYBpr3ywCZ
19mHP7FAdFpZJRF/k1z6SMhKelBafFiNZH5vcEw9fL4KxzHkCb2wiKuVf7XfWMWR
0c/YUnj2q5JDt3b4PUlmhwP+ZXcj+z98fjNOF9YYS5ANf8lc0aTDCUhqdAaXvYlC
dIpAsDAb1/077+VOs3bg7IINiQA+c6zx2Kf4cdylg6v/+9Yf2JRaIf5T6jFmE73y
GISa4h6smoWX5DjYc29dmLIEF61/rLw275HTxga8YBTmX1GybC3nrVVuZ6i+PMlW
ZDh1SWci+W1Ste4Mn21oh7zIV+scYM+SMAwTIPxBlM4g3NcwZFPuByBuy8hTp250
4KTWv+1vpiaeq3g8H3UyOLNIs+OajQ70XKYsyAcqohl873kXQydqaFVp63HckbJG
qjkmOkYUmuFWxGEiBdRC7GBhellBkR1Q7GtCAcl2F5aJlzxyPlS/G4JY0mNjrRJq
a1uvFhjsPe7sVzEOxmaWKO74vi1CKcsDlCKbPzm2BDjexruEFp0as+C82FWGFZ9W
C1E6kvHUCusyW6RmZrl4tY1coViz7bbX76oQz3fmXkrN9G0da7ghsEMjhAQn10Kr
Sk3JIH09+LTLqF+KsDNLJREtTFEW5QGsZUebnYd4R6YWTq1BhB5sE/JO6N1VSQZc
WJchOpgJNF/Z0kKrGFHIpOy7qpCiBFVLdMieVgIRNGuQsRBarhrlxTYTOJg4peO3
EXBJQqkRgLJP6YTrCr5k+0bhvwbOu1jX73Oxs5uIEOZQbW+dtvZ31kPWoR8xv1cH
EHtr5UUhzGwhMbgU3pjSBoRAZyXEzNNfSAxGiPngLFaAl7oPAmi75g2LigbPjWxd
2WGBRGXSrqzTjyz0IplFEUZ2n8G/hhThBJmxVkWJf1A6sbdiA95cwHN+fXFlNQLK
7JO6EWM4Uk9yDW9o5PGY8M3Cl4DAJL5pTctIagCQdX962tv0ifzyNYVK3xRlFe2P
KejeLf9C+ZFKZ/c/5RRGqKjbEiuNMKM2YKB2IZFqgykPgBod70ssrSyD58ib6C3b
jSnavShraBuFSewaxNFM09graT+Nlr9rtsJ/7Jqz1TW0mnoDn4fRv9SpzD+7c0yP
PXQP5gdp2KY4x+IVHYJkEDCpG5j0RrK/vEmoG1fn64zmAfSGp25ExuTSOfnkbSAj
kqNLzOv/rSycoPdXo/cxOhZsAyk9GtKEzfLl7TPtUIKz+BYSZYNeJQxgwTpZUs76
rykbQwQxH40Qzq7flfiSktMstu67jHEQ902q5afm5gwJsm21+M+LrJXdyBgJ+E9o
20RImSZlznOVDqwwVaq4070H79yFY3wCBK023NQGF+L/Wcks/PNcY6cktW7I7C9H
sEAC+jlfxgVMUCM+8zoOYTkMMKBJ8pi+5qrIVlBSf/mvPd/f2xIGBv+DVMLeraJ/
PY1f5Ev5z/wpq+3Fw8UkYdnhr0nvdE7OxfGQdxlteenZgqnOHRTUG4I+drvFQh4o
kCI01be6f2xAuLSzW8Xgzu2aHxgK3HnbRB9wIaOsoEzf1WHaoLz1QqClgKNs9W07
95XwxnlzHWEszQ32m6qNyfdaqCluW9Et6R0wX2FmTkez7r/X1Qv1tY1qIrjZI5lw
wJ1xKQ6zpdxnEqB2J5S5pksFMwVIR9/cnoKsMe1R2C94OLdGgYM1a9jo9O9irqeW
dbnsUgU3ZpxT6roCsGDdMYfMcM+Hw6jym/got+1u2f18rf3k7YUfHgemhNhlTYuh
Qixvf3JxEOPjyeLBzJZmPmxr0ZdnbcQgPzi9WZwh6T5GkG0amVdAVTZA9HhPIGyS
DI7Rb0NIpwlZrFqaqBp24UelK5inVGIcOCyuYobl+tX9T0KPYAuXLl+khfQkI/Dx
eZFwtGXf0tc6+oasok/u2CM6UR6kJ3ze1kpSgG0Tke+dHFPV2SWdt9cdDAfLbs5d
jkIvhOnbGGCuFLDCNMmb6E3erB7040raUT65r2OMy0D7VJ/tYlVtPc1iO+/LQSTh
TjoAv9mM5NqjtGy85dIQ/x1Y83sgnE6W7Y913BIuB/ddYLZ/Li7Gye3BO680/gIr
1O1ya1i9PmiUYZP7XcrOHUVHvfesD14Zsm9sek1NBcDMJqQahdvC16H6NikLZ7Xr
7vLul9jmD1Ur+sx40+FW2y+ifIAb0eFBKB1mtEwr4EkedicR3927IS7dnnP7v0+T
7xAtTbk1RhuRSILo8c9mqJ0p5z5Ia7vKHpUpg5FwvOVD/zDbgQLQrfkNaDejnKMd
URfJMTj6LJ8OchbymuDEuYbiQrx0euGNrIxXP9beLdpdPZk9Tv2zP+RaNrmDITJf
j8/z1tfdKUarqoE13WPzsV0e4br5U9IJJpJqdGiGdiSHLV8B2EvZe/PXbj69lrmL
WIq9QXk2R7ax/bnHhqk7h9gzKdQmiPVy4BHyItfSptNAqkJfShQ4a0+VB2lFURPS
VvxiT7n1kVUbZfWw3ht7AqNy6WkTVu5IlgXpwipMrYZoBirXZebGmeWs047Uvvb8
QhY4IAOwreQwk5zZNcFbRLSfek3x6FpX/ybwksObU5noy3XYulUIcyfNFaqptdwd
FHb30VunZgbqPFIVOHtdcWEW9Q+CdQML/OZow3I6PDQ+FLaIFBNynvkMXANu1dJa
TAAAgfbffWtuT9FijodHsda649AEuYOt/VsEgAi9PseQvz7jfK4xofbUFAJ/zh7N
YKBSjl2FiQNN9bvnGsQGTJ3cO/JLZFaJLdlsrGBnKQoik110bUx2nOd9FmabVRJc
7fimSS0GxsZQEAiRUv0L8fqGhk1z4p/Wz+NPLWgydDJHM8tGpvrKsofylFr2LvZR
fHXZsvy3Ac3b2/hSI+vjxMErXCU3uqg6KtAhtRBMlOFFvrswRqaWhwtE55Q7dPvJ
6dUhp6YVQVdlusyuB+GmKkX0jtoPLFAkiqcI6+pPiAzK39KzFKscwkFafIDHQRo8
9lH6eIFQqpwugFBLxYkpaQo8tH5o2u4iIW6QhsFFq7QJYpsrwNIMcfCwYNXgLyR/
9j6UNPbyZtRqu0IU3m90JJO7gV7sjDic3LEsOeqpV4Kj3wLmevPlUjCJB/JBSMzi
7hHuUiqQix5JasN4QphLh0mtujUtxJB8+RIzsAgqf+GURJZ3uprsetcuKeVKBhjq
n/nJIl3eSnZYYoJV0ku8FbUX4kuxzvzF7l3cRh5rAsaAzxkT71Q1ch29jdqQ3zXC
RkWHUBwEncRTNteCQDft2+nN+vpNmwv5BknGhwrp/Gpz4wMGzaEwuONK+G63G9kf
cKpovbiDj2LbUrPhBWzTAIPIlD3DAYdqpx2ypHkESIYlja7eR7sRk5dqWY4IgV/6
5giZi/svrAdArnLolB6Xf0ax2j/KxDmjiwHNBHfaVp/5ygEzeKmfiQtCd6xryY+C
WYnAsK78P/H0wyYi0U1dmnzfg74R+3Stxmqgecww7R4QQpX7NmnlOWdE7mfkIQW+
EoFCyN+VQEFJIKLIqupRqux8DP7knP5PG+0K+z3z2eewd6i7hCfVifSIZYLcmgR0
NGayLDYt07I12Gsn/BFldbxMFivqbBQZOrdxx23T1I5AW3FWhy6ZkCUsCqlbjzjU
kuUeXshY2XGzbN86JN49ZDcQFi7AyVzBhnMQAgUa+oG7JU91MdpIvi6sY8KQzw2L
qw7WMy/y0SxI28lvZUHbEOSaIO8JDgDV9kZ8nSDB+l47uNlSCjFGNPKgpC8I7zXL
JW+UaG8TMiVj5NHZQ+Ta7PHw4gH8z0lOxeOYJzxl7VnhDwWE5Y/Jfh9Ro9GrjBqa
1RTacu7++loAFc8+7NEZlb6VYQ3L5IvqdeXJFACtda6zlZHcbGOTIgoNG5OReEu5
WBuABv+YHvRv8UTvh4DVE4NeLXrxAFCvY8BqSvMvXaL5dLj5phB+xDF6elPYeVUs
E1JVsnY6eM8eMr5K5inGoMP7B3R6jfga63NBpkK1pOdSR/+ZrPiDNnrMy8ubyc3L
yrQXcUL2/XWdJxM1aHqiykRi85VZrQ+AOPRitQXKm+QCha1PGiQrqTd6oMFvByNd
IdLP6jclyVUpFOIg38U9oiYkkFaEQuddGTvOvcHSc+qcNW70DmEyKllcOtDpkUwr
fuxwd6nBpKaD686+L/rAqeCeKRcBXe1S0fns0HmRK244XGl+LeQCD0j7pO2ndmvQ
7W5GrV1XzDhk9iA1tnsTfBaga5GBoxv4KsdLcDHe76FfUVoqaj9c15iEnaXb+qNy
caPun6fjhmjzy/NFbzjo5+257K9SuB8Njc5s7ozpMGWK+zG3iGkuiYtErD4Jt7zx
7N1Moxd8vftiF8a924xSO8kshkymOfGZ2JrspExq9ZUqiv7zp6X48LKmz1JdbZok
ITjfzjVG2RFGJ7gRedmxwvpJBL2a2EUxKqprWl0htpjflR54hAjnFLWpxnLvCHkz
RvH31a69t7pgPAZuPP0lhuWFWya14pNXvgJ+EYw39YIBae69qrf1XNpCiGZ5hAZF
sMNFqYMwlD95fSwfOneQ3VSJvzWAEsg1RTYms/QRIc0Vw5al/vVY2YpM1Z2XVbFY
61b+7+7xxOq/svVCX2wTK23/U439KnVSS9S82peYdgFsBy3IcCS0JFvjVDZPKlba
/U2neITOmenMUvuFMOzRqEgBw7ez+Qjnid48aFT5mcXZ0YNxA6JsAZs+yjTYk64B
WnwPHOwmM0/817y0+8/VPWE5+jOiVE11jAXakV3UR6hnQTysWKObb59yHVCqZAyd
004amqnDIwcAhKkLcJWHW/8Zu50CesBwUj+/Ba413dmrBsu5sU8QPEi/B8lqbVkI
omBcQVNjegP0UF+T5cW0hBDYFd55hGiJGivUy9f77VllGrAyukLF1+tFdvr9+0Az
bBvdtU/36KN3dYdOoUfimo+DNk7HhBGxE8tV0h0SJxFBD/dmalikcyCjOFnun6kP
nBXbaRqZE8Ps4ySEOC1rZnpwSox92rBO4bxCouiYXppqgeIcSf5f656wcZ9Xoj8V
jBkQPmce3dMWRIOTOwbP06Bxul0qVpG1BKnvY5IE/jWMb9RGQwJcBYCT01uMF+xB
BhCS25JBzeroT8v5s9obXuC5dAQuc5nUYAQ4dXSgfyTOQXMp4K5UQ6nQaSwhull3
RWqJrPmV6ea85ifL4SWNe/Dy9Knnv4xF4ptAm1Xp2K9hw5ai8pBZggAHx1qFcByb
00n0HMzlKMML6TEQt/8sGDLqbsiskYJnhvCoQiUyaJQQ6d9IJtVSaiwPCpFG2BG3
JtdEQoE+L66qndQBKstc10YvwQvP+qHoJT51/mjumyH3qP6HYgnOcl5wNlWyY7+c
oK6m8V2LkP4OQ9nQDbIB3VtwLUHHawTE57tp3EEZ+wHxe4oAu5JXuhnuY+jEawcO
MnyeNmcHDgNV9v/3l5oyt/7gsYeqxtOCenLJb5t/ckwDjNPlXbWMv59C4KoBkVli
Tdml3m+XI00XRPdlK4O34inwTSP95ZOCXUVxY/z10rl5beS1s3+erw8KUf10Ffgt
efpdfe37V+eDhS8zTG8nELY6ePo02dkGxBUsQcRVwGLt86nuUOcvc86fJU7hnmMi
Hd0SNS8wX7ZNhoAgH5Kbagh3RdvhARvhLo3PS7t/ECSqbP+evwMxeFq1L18eB8WI
o/8OgeSAvd4N2Fi7T0kpmK+cEPzom3hAj9oRPYcRC2z0IsQduY584+4Ylo+1a6lD
HSsGu5F37NrjmtO+ohvlY9MsjCXF9g1ENh97dEaSEXUbA29rhPoyOYYg1MxLHQhq
MKtb09cXT7Z4K+6cW4jXLsBkfWJeNok7qhJ2RKyrqWenf9g2JK7xSzLIbPyLoFnJ
EeOZkcMb8J7QvxrObCaMbuNc0bIa70sA4k67BZN0HcGQ5mbZRL2UJJak2xxaz+85
WodWBfWBm8SluBZikzdpszRZSNHuuNky6PEDIcpukhOC8+iohAHvj1sOoPVEDuDt
cW/I+CIwTxGp3bBflLn78jqXbL+ll6whyCftC55X6vekorfN7tAFwsO5zhk+22D0
j2a7lw+qJ5dvrd1G14uh4roEbddgPsvYrS9xSrk2QZb7HErB+mjYKX040Cg/YGTp
OSb7F3edlr1e2Cl3ltFheWBPwRAfEy8UnjJBJ4EDuWGeQ8eeHxM3/1NrfPVGUjfX
vU0d/EBDOLaUDspoqww/xxZmIC+UhHNM+eNv3KDIHEIsNQ7KlJyfspaW04OXQGvK
2dvGcSGEaVFXhQhEG/G9WddrMeWiugdrjLzrkkq5wboxLB4JpQLQfLcr3U/5yPDi
jxNr91ri60ojLxMnvSeK8ApUKC345lmTaZNVvFnQsc1VMCmzefjDB9dtdxn6LVix
TgNsV/Qz/Hfy/BL8Syo81wsRUUMJ3rWFmwcOUF9omJ6cQ11GS8CHG9Mg2iYi4jmT
Ea2Maj/xh7a8U/R+DAxwcbR3jS29GIQvJTPOOueDme+jOYZvLPuyk6mI3wR5kIgX
g+UNwJphIHgWHNR0RbnJ9faYgAG2Ne8KpzhnbxGC41GB/mFrbRnU5EG1YoxZgzzE
uL4TQwoVGYzsHQe2Mi4/Jrs4HBYQm3NjsA/pwaYN5lB8f9w52K9+mlIXEJgsszHY
Xi0+kQdbLjJOTLHHl6hOoaWvLeYOLr5gsUnKag1502SSaT3BYdBrgkffvZvnJWx7
1S92Vg7BoFFXqNHI9WcAuXbDw0y0fBa32ndvj189jSbwJPbXHIAl2ECej0EUm/Cb
tD6eNa4qAQDu3mTKansVNNEqXhyktWASVqYckMk8BBgQPu5umagwQt0r88U6o5la
YxFWZWH2SuC4pHbxRmpQtst0HXyK/g/cMax7inK+e4M0auOe6m4SoOPuiq32qgNC
o0GVexoFQh2z24LUBeeID9AOgAl/Nq9wZ8vc37B5FPiU4fLkOM5a9ruoz/oVFng1
kWQx/eWKm5/Um4u+NU0/UTx1tc8S2keXzZtU3PEKgyNT9rcunBa5XN7n0wfAgxLO
VJ7jeQgTDXwES63zBl1tzLaxc4cVOWC2km8/o+n+aCRtaowbkXj1NSNWe+l8VsHn
j5FWnrXrPn30h1ppPuXpVjnFT9VXBwR4PdzQZIA1EJdDTSFkUiWZyI14Qwws6VkL
2o8O2d4biOsIoQIxORveB/JNPrQAqpaV7J9xHCzGMXlrtPxCJFBRrOFCRU0xu3GA
2R7GxjNgZO4+mDfwSBLDltE3Omx7+lSQgNvNclBPGsAbfFAtsUUZ9/yKx/cDUJdC
JXRVPhkvR/CwZtpghaa3pFv+zOjbj4aLwf0bMPTrkPx9nvC3KKHO6JcJ+ycFfZbN
tOzdup3H8OmOKF+DipOzrJ3Ala/r7svt0zUsj+EgZD7bp3O2uDRbE2RfPE8NJfTX
YWLiT6VEUg2D+5r7MtX38mB21kBd7G4sIf0jdK6o+zcN+iI9vPk8kU/lKayRyOgw
kBeEvnpUKZkg4YPPBbQKwiLxV40f0yHGYYul7gCRCDp3/1DZWoaNZ9T2GSL7KUfd
5iEy6LJIisC5oBOdJuHAzyBE5cAPwcktC6KC6pwY41WIMT9jEnw6O6tn2UskcBBi
Z/nkFe1I70BHUY3jccHVzolBRjgEBSWc9JoK7NsQowrxk6M4uc64NPszjqjdFutj
1aMDjkQ4H266IzqmyAaRKuE6xjM7X2fOvDfJPsf2s3SK6vaklQfiMDPkBU1snI3S
30TczUk+z2OnlSdUgCUAaPMg39I9cFFNwtqaBgvVTXvYzobVJJFdiHiXbu+ZhK4D
T/DoUIMGM+bzDMcfRV089CBS1JKuIB8Sumy3NwPtaHCXyFH378fJVzfzCg655Yuv
Xxd062cichBJNc1HE3cm+O/iYD68MNd7Gbt6pyvXo/YopACRGZbNKaC54XHPg74X
/QDUjxOKcCO4qXhF5Pe0AowJCe0lNxqkC+hQfZQOc6XWSg9qBSLHJUZx9QoQ590M
KzeKRYeykuLo+QMtfrw5FfCDaPEPE1kwrJBKQiAg59bu9Z4/WiQYPsGXQ/EXjtGT
wSFW7zWVRay0Fqs+Br3RYr3b57CYjm/31h2W6Fvj8JrKFj+Zi94pIYNPKBG0cEpk
EpHVHKtZnC4iX2XuKtOpP3r8FiWkwF/Hx8DVptRUJdhTqoJpFotCt7XyyrA+MG9n
r2m1EUIwZTCjw+tDzxuZabud7XF+oJjHGiw8Wq1TRH7emvQAD/6Co29F3NenaMnO
JyBZ7qAa000bxdPyp0nCTLxatoaW/tyPhkeRUNCuH6iXBEY7E1YyMTvmakzGgXgP
0OoN4EAF04UWe8DnmE1pTzVPtjeQRL/VjpH2fCY75qr5FzvcwK69MQpwG3AwDX2u
C8YEZAMZ+aRrvrSZJDRXchg5dmrn52nX22hr26UUxK4pCrcT1XqqmLcPbVx1vs3P
aKXyIYjijrJl3lhiihL6SZylLPgMtKm8aeZusTiBITUCY/3+ietKxzxuJPb/ZcM6
e6j70w1yARiXzZ6B3+ay1YxXljiY4Yqrp4dhGkqgoUCxiW+HfnTnjqVnfENII3+7
i5Kue9IbjjLDrKjZsugJLn+Ya9X+6sAmzmzfPxgnYM+OWW+hSg/7SkjuD7mhJm8G
L4VMNF3H3jX5aXGT7U1dmjrIrmNVifOyUp2mQZ3/p3N7VtJ63zmQ0guhDmfWpCyC
2mNA14VjQjMrAmidg66VqVbUvpu5GJIkY7fM74gl9OtEKBpsAbwJ/IEvlXKE0DSi
UplA2CFcDBc9r0qLrMd/j1nqIwXHhF5KqMfqp10fjdQ2VfY8Y6rWPmad+wMmaqiy
GRLOD+5axp0kwGoMWDpFWC+jtEhU8jWPM39sUkbHozzx5CW7uLrjOfwakZwwjJjN
XD4ivmSe6QITdQ+Hv95bUQSOk5N4lUW+0FtaU28uRVl18aH1P9eTjOpte8ym1oqT
NkCWeFbhUu1sbkiOkDnuKXO1N7Szcn+12tB/O0r1i/CVUTIYr8ksXgR1onrE22hY
2vQdMykdPCjVMged80oSyLQzDTBOcJ5mf0BGADM1BUGltTOwG0nL+TpMVcm3Zqxq
9aqrJ1dCA0CX0fEAROXEc/lt2NL+rh/7PI3erfd8CduHVG/IxEjVIPulYcARxCYt
lDf/Jb9JybGq2btmVXAd6zSac3wmYnSmZ/4U6xJHJ8JnjO9erF4cQvwp5U7owU7U
zVNLXp46dQH2uwKdRrx4UEYt9/YyCm9NC1W6bG+TU8a9q7eilvRC5HDjacDmrFg+
eZ6kE5ZwjCFTygBr6RcNc37aP92qX1myhfxXa//LL8hbgma/14pRAChnCzKcIX/b
uO7aoZXTGKGcD61xPi0QgQRmK4AfMVH1/3C6urmpFLCylLFhXIDJq72gzOBGCtHL
p4Ah/IgTG1J8l1kmyyEiVOMeU09+6iw4FwUQADdyE0zwFLQNMestRz1vl7cijHOX
xmkm8siz7iLl5BYnYtSICuSD0ndhv9B2MTXyD65KM49tFR2PO0ayh4T3pHqr6wVB
bNDk8SCczp/ynIrsL3Pj1GhdDN0ZASGSKXxKxd76zLBKtIgnTbdfZZsQP0vZrzGJ
fTv4N5pGAMTcHZ5S88kfjqskFr2gF0J55QNP41W7AuDwUTEKUUY/8vQsgXnY1nm2
8wBut5ksR+n54oF461CVLhYyHIl6oWtCs9yxfG/HMHYDgAAEGVp1VHL8HtqOlrJs
t8VDEaWpOV5WsOsFhTa2adVMGg0OfMlvmBtiVsanociLu9VtbmpLCIj7fAgrNpcR
Ezd4zMywKH5cuK01EGlC37ga4fDwkOJ47MjwxjVxL9PjHiQizE48IVV9Zm+/hN2T
yBgJsC3Yca1dQn1jeqCniVUXP4f3gRAqfbQpqwauWOpBxEFJJZmB0vwfTJY/QsMI
Ubo+Sb3IseJtXHvPJIAqSCy74f+zt9P6K9SgBwbkH6rhYb5OK6VMaqA2vKA8qZE9
kmJmsShPGL4Yw+cWlD+EsKvSirv1GSubbCxppZp+XT7Dp19c0L3JaVoWRW6E66Em
UnCrvNvwfmMjqooeH3pTyfwMl2ZS1M9cfxBl8Pe6dNzyfukLvKCm0S22SgsKn4Sw
tySl61NiPnFNC5hZzAM/1hh+pF1hk5M62kUtvV2dHFFgk09vreyZywzvAWPVbYcK
GGpuTf0r+tJCsgflMj+0Kh6d/dVJ1r/LhJNFrGzzBbkXUngf7zb53uNTIVMGqr2w
QdsV2ubPoBH3wlUSV/7uBG6PtFl1DD8SNxRh/cgobW6gw5C/XmyAQHkYngF66AIA
4X4S3ORm8HthagZRux5wrKtKCOZ2VIZXZLvvTiY5bnNZUlnhPYAJhVXUr8wLpgQC
ku5NMqnAWKno/JA/cdyVZJEak8TkKoAuuRP7WLBA5tPgBtv5TSCN1GraCJ3XFNJv
D1l+ZMgcYhUYVLkPK4l+6I7ADvxIPzUc8dsFBvdn7tNMAlp2DlDNcerr0Dx06p/x
bdNqlU8phzEseFIZgDujvUfwThXEuWKuL55YmDklUUGqmeRyK5giGhEHXmEX3x8a
Jy9PcQEjpGvso+ieS/JTKheoNHHHm8Ma8jYPD8+FLnppif8i716i5RLj/AyarL/a
7PmaB/n4hl+rxubnr5zOXIUcAgVD4Iom3K6YP0xrihpGR12mtF9WVtXCOjxGi0Fv
TMK0BwlBoTP5fWVbGIfj6IJftfQNm4cGTjj3N2Ulld57BBfe2dqqL+sC0YnqlIDE
5NMGrmDmLZtz1WUuIxcZAOkAA/qMNLS5mnmzzMAQQw8cDkPtMnRbVgHLUQ7JqJhH
nHoP+7Rd0dGUpzQeAErE4mycbIZ6ETYHHdm/cuJoTZ44iS1ecXpgUG2gwT/SpXkE
1YVdFj7sfNYL2gVsUL3unwLW3TNvkuBVQkS3eRh2ld9xHEvmsnREQ8JOVgSS6Anx
nd3o11O6DItjsK72r2jO1vd4ewtsAm/4LiB7lh1ggot2h33Q35bEGAOWUx2KPH8G
UlrcjDgBI/Q1YUc198blHmMDr5VmKPnPFGCh31JeVfATtUxvW0RjqOxGNeL3PC6l
IRWLeUg5S9FKbr29p9tXyptOUJugyavxGL9gIl/uJWIFEf6un4gCos9ncV0calNT
d/0tXWwvhmnROBrULBvdVZh5saDQM7TySQ3SP775mkMzyyiwTrmHlfgarHW2G5yG
LBZss5kSD6RfjeQYy5evglK7KyjVbRZWvyGWxBnz6Mzp4yONZFLtKMoy2gS9yapx
DwluWpiwO9ULxhp9YT7AQEFMKvldpw2hZCiP54Y/e9TdvBWy513/STrm8a1TYQwA
AulqNFGcLTxqS35yib/9ktTLkOFNpRlAKGQkaNRLbbyrUs14F9YP+jxyXmgtQBgL
+FQhHl3/SWvFx10NUIgaDTBocUi+UFPmuxq6JZuzo1zPBpg05zQOIKPcJyT76yPV
gLfpu9q1z8wGJqSyVcHdc0Zj/B/IiD2VWY2pKJTc6ZI8jDzjkrfVgyBwIfN4fM4D
QG8uqchnlkAXV5bnxGr9Q99u3J/kSfAlDAK/OEIXIAWOvpIQ1zsEBZcpOzeotsGp
MNOHHGnm10bGG9FB0xjRcmC/nazT51iMnDq8LRGjrT7fjoqiau2jWDpTDTVnc6KC
od+cO3D30rSssSDlZQruefJKBQ3x9t4CKSIfOZWAX9pk6G3YWvT/w63BEg5YNgcD
uJLP6dlOJ6LbcnCTO5rNIkMYAy09nfRx8fYsYFJbR2L1iqMMio12FWB+6aSpI4nJ
1ALUL4iHVEwciMmGd2zg7MSaQXLVRXh7Mt9zw0k9jyPgJPsli/wtOj9pzjR/bPUM
4JSyKJXhKiQ7cSJU30eqoISSXHusRVgnYhwDBLX7xBogaKXQsPoYgFEkqVvPqI93
pPSiW+t5p0H4pgh4yaAmkcVpUeHHqkqZLgRf2rEdqoVX21Q3fJYl7AmdeILhmazn
iPVdC/U0ZcLE0u3wXKSsoi6OWQNT9MGN9Li88YG11//lw/dPrVKBRJQoIW8X+lGY
7DO56RTpzc6x2OJC6ymZa+1SuhpxpCj50ozdvOa1iZwXQUeeghXEssCMLcc0wpUe
I5CaNIZmwni8/P1OP+JWLv35nqABZ0W+10bkjNUGJMzxh/pszx4Wpd3fCrhh1Or6
oOdfzPVyLrnh2IiSkLy8jIwfXL/tlO+ejw1Xk7TKyWbXIZrTuvoxx+UloaD8Rihu
ACT5dZpzuZvamHMIccoDtuQ2iXSiydOLdSMVBB3mOLp5TL3LP6o0hztljDd/9+EW
NdOsKXi7PhUlH/9Jdjk+PJOlSIAa5YRt2f6Lu3VA7eE4DDG1k+aotU+6u+ySFwJ/
XcAy3lZf14+8LrjvQNeusG0IWMT3JAvCPc4LMiEyO9vnHRZXwztJLvSUDp4YIRVG
vMZYMJ+jQq8jplptBC+NC9PcSzl1xdIohVzUffyTsseDBfsHmt1bh/eZA06Cwgzk
LtHHYfLGkYvWQzrLMkRd3vm7GZFanrKPMyQChepD579yasfb7klHyvTwrQ6jB+PR
Pkb+B1eBpIWctOxlQKbaPQtB9aZW5xCj69/8y8BsGUHvvWNHyU87SjdS/0BNmU0R
+A2ZFBKf3YZ0NVlMfgKVxtJkKmx42zslQx/ccTpeH80eMM9F1RiGyXyAvacGpmKU
BeeakCdWmcAhwl0Pchb2a0tRLa7YgR0Z3PiTb9p94qn1DFGIOXJJMByjJ9IcLkRV
QqOuWFQe3yuW3fi3fn2CYNJAWEQagtx46Wgiauovvyi0CaiJsn+dbZwuwOgIhylF
c3Uw6vumhnKHQVU+StZNWEv3wgEWN6CZ4Z7dcRYmg26xhGhnrnbBIe/9q1Y61RPx
exh6p74r4QctL0gWoTvIbU32j9Bpa094+KcTQf0zV+oQmQvWV9ha7SN0/IDv4+hG
PZ9vsnOx5QX5BrUXKIO1krwWS+mLROs5iM0M40Gfhw3GW41O0vnIaSCOYueA9oZj
MyK8qiy/DH8jel87UPVcP5EkEWPKd7Z2S6B+0/WhsaONpDALCYgmzwwWLAVt9j0F
nAtiZjwAsjNIP9j8mn3xIYRJVayTcmakCGp1Q1Uh1WStQAXPmt3Tii2lJQloNt4T
74FY/UtsVzvEYj+efNxuf7Cg3haxHsOdW5UMArMKqiFT+JfTP9glDnwUmK1Qc3RK
FetnNG2kja7dHhZj/yUGcPHrW58lxkIgdo7fihzvaBy/7lqOIkGaY04t5MjZwPpN
kGnEocuLWdVNTivSkHBe2HhfbfB+1QSgT4R8HE/TjkF8BYnOcZ1IcCUXUh3HGN6z
tofAPBhuU+HE+nwmk+wobl96j4vHR23csux99tkI7zHdTNh/TJGQUL33EWmuwOnA
1i+p0GpLAI1R+N8/fjpJEKn3nrFOd2ZcdpMdgraE1GuyPztr9GcXUQdYAuTCccRA
4FAb0Y1iY9z3j6E7WEjQS3XHcguzYKGhWFG++HORl6J6rJz6vtLSOCQAHMP76eY9
h6Lsn+l6Ifx9+5JkNq7JV25K/WoIJdR4ib+cIrg72+Hk7TVecksHK9mOhvgJL8Cy
rnoenNOEQytPj6J+JhnFMwb6aVlOoL2/mT/jkNkqNEyVwpvin++prkJcaGFjPwWP
7cyDiOJRGB9b+c1PPx9dzBJwBMRsEGtDWtFiDorCno2XSJ629S+i+3BKZCD9v9G4
/MX+asfvi8m5C6juvhmw9CLLxAQ+UyRH9brnTN++f5V2O9gkc9gSMZPU5U7X/OeZ
mMpG/+ihJjQWFlFwduY5cIoeKor0fsSf/Fl4ZlwXr+M4jO9Jfqt8ldvYlDzyQc8n
QT24u1w3R/aEOZ/+yQo0te5X+Z0/8ReVSiRWQAyJJr5EtaMj/TegNyzd3vK4q9Eh
5AkMFP45fCFGrnFC0SYogMhSP/rVIdfg0j59gf7s52CQUCySZRX+TWW996vbP0OT
k4Oooqo/3QkMqRJH2XcRD+uU6+gdt59CJ+jYfa646fJDkB96lTascxYdNouuGgOZ
2qywNZJMSb8NysMryiB54Bl+OlfJQbUE7F3ue9TbsK9kGjWu+S+mZTuiDIRs3iWb
N4qvsZESm5G3CAHa0R4y0tyaf5/ewEHTlqKUypVAns4wPc7+4OT5EtBn5tnJiYoW
DWR+7r3f7PTSbcWgqezriMYreU9bxZnpJYR7cgrwjqJfSgQ9UB4Xlki7qYk/yhWv
pXn33qF+QFu0+KaCOpctNLpRsQyZIWPeSjCTM1eTwFNUG3pohyfcNS8NLEjtBQgz
tDZjNBwOEcEgl+iX9u1x4UEysTKN+5m+cdF3RPX5i1tHOVjtXekeAX8JbK3HbBLd
7yN1xirQYUn3A+JFl0J6c97k6/NUoteOTKcso0YRPAkaAuYlgZIILQ6ODBanwldI
ACD5NJzpli1/LrKJco8pBdir3SL3m8PyUmtUBVHuwHdLKSxGbfGb5VPX+6zquufH
mb/qlMbvn01kUPiuj33ovGVamw2iRt9h6zznCAPPyxrEraqVj+3dN5+qrCh7IQ3Z
tAvu5M+WzxmFBbuy6FZHBDg0SIXJIBnts/FeL7cDrWj+CUCETBbjsQZkg7g0H13V
wn2ovqVodYZx/vaJ2NcLn8rU+RRBvkPh1COERVvp+XmixYA/d+iXNKWQGPDQNuRi
tgQ/+c1p0zyFoP1F7YKEgZWQPo9tW1gaOdVYx49N1WGZw2ur2W/oyIqJdozI5XJb
pNiBm4Yjg6UdBQI9fQiXe2syRkUOsRSs4svSVeoBr8WhR5xLHkBZw0TMwarMUcrV
4hnaE/FWPlybYfCFZN9WOslAZ7UxvUyTeGbM3103nmDzDCyOSRi0wi6msqzG+r3R
1TS2/wxjM0TuQZwsQjpN1GwYxXF7yS3AR86tOEPcQGbnVA4Z7E+SP+08uVN1eair
gtY2fp8a174T1WBK+4h/sdlb3LIhHwHzc+T5BRJMqFDW2WncvW//r8QL1V1RObmi
CNZhMUHitisScozayYM+myUtdyyoknfe+1q6wIZvkI9ySdojTXJfjg5GKQApQ63H
PLNWYx6xc0brHxNzECiLSBSxJZS7e2jHYAnf5+YlEod4skRLltZiulj3bwkUiMvv
dfIJzciEjmtHzk+LzI5EqYo/klZOkQomdJ6lQWHDI3J9HMlfxDlbykJkBX6PJ9BB
JPCVAaCVne/B+Ncu+WZ3zu5dsgOMMxPjUUyRphPOmK0+QhrPYAWBXStsxx0QSb5+
entiwc8+CJS3wzLNEJz7B6TbBZ4tslyxp1HpFrtp1M+3oAgAVDt97/NfUtWtACpB
28KhiDW01gW3cs5gybjo4XfjQwQMQYWIbrGyabBHt4GY+hYnxDIu9uAKbzs1qeIP
1kU2nQf22dBIEWhY8+Xub7OllEccVMdUGzoXAJLXcJMdmGnfbhwDfDZNRuwst3N+
gi3MNnwtQPgoqTbDwlnRNAhNWeLB5+Rhw7OO67rYDzEeN4C+x/0G5BDqO3QNOUy/
JP00vMZSRuHa3eoZksBSvyWJZlY/ENjqOkgFlCzcEjbnur1489VDUwZtf9J+u5cq
plgWdgiNYkk1DT/0LBbVZZGXqrTYa8PoCDdq49fL4NplK+G1Sz5z1JbCxV1QjopA
VLfJHdQJ3IKAhuiSogRTG2bNAkw49e4+tjmotk8oYwRqOhLEEYV6rToBmo1TU2aU
BExeXftH6O4Yy/bQtSeoYuputjwrv/Xep3vM6hw7SX1HSNRzd+waqJq4eKKfnDXG
1bEI8qI+aUitsHXNZA8ZmoeNPNWaZYumLs265kuOyVLAPT8HVt2ulasM9boiM5no
p3Moy2MnVSYIiwQgU8mc4b1NDfwo20dcYEraOd9PKBbl+6pWl/FrpAT+XB2nnCbH
2DTrosgvQSyuKYY68GywtJ0mhiOJ5UBdKyHaBbrSkySLOEQ2BtFIzCLebAyQStZV
2OuxseDU4ekNmPXW1/ET0Vv4k8/VFj7HybUwT9/smEJ8tgIqjOsvm1VnwIyKXlLm
UalPidxHlqFj3tHNQPjuZptr2AQpoEQjqBbsqoEZKCptTkpn4G3oNIqD5x7ULKKU
fYtO9F9jPGDleFIg3AbYT6zHd78VnNTeu7jhYhq03SxAzBOgthQULZraVhTRIFER
8VOWAdy26ibMTecoMEx9x+sQ0kDxbufpuWfhBvtEXZCxPEeJXCqVKbwhOiptScn9
DioAlpUpHf4IvdavdhfznTeHXA29qnFFVXVkiSgi0azLH7pSkKqSdTqdR2SQwK4H
IbDyjbH7qzQyAi4CKS8gsXtgvKWbReskT9CWLtmYOVoFUF6AB7C4zB4f6L2P6XtZ
0O0VGrP8hjifieT3gzk/o94/gqFGMVu6b4jfuucj2askEr3MBnvMcfR3Sa58prD9
BMmNIS8dS7y4rcK0ut/Ms53cfz/ztaspZkOpo/sH9ELMEcI2Jxk8mYRGSNnNJDJW
0DTIu9xXtcgVYdAYCyTY8YMSQwuyveMAe7rbJb9j9W0nV1LAt/0IyqksfZSQbVu8
J2SK4NW2iF38Jj3bT4UT1q9SbkjJhcK7mpcPTmFI+RpEQpGKfi/rZ1LFF62e5+kK
PHIj4gHZLRWKw4NW/NehQzQTPqj5zCp1BbaaL/qnmq0tX3kfp5Ir9w7Wj0Sa+kRR
BEFfC21YZQhi/s7hN8G1NQ9rlLIiKCvcvNaVGsamCUEUlFGHKGevo2McXuBBr54K
MtPYACspq4wyh+2pp/ZprPTFF1ynlJRzkUd41h053r9qNzmVOQkCUMZC3Ncqe3PQ
lc6AYupz3No6OgpTWdg9OHZgDCZ798SB1ZyXV3K7u9dQ8S9fai57LsmzGQdtxf67
0vVCAqKDDYbnaIl0p1gKbvk9bIFc5splspZ1kyTnsALiMH3KVj+rFob+60BLMeCM
MKiQ1TS1s3izXmD9lZ3PL9OKtubgV5JM9gcIuwq3G3Fv3UtRSF7p8AeMgMyPRyHf
I/Il7tQY8yntLODRVUUtxJK20XCHfGZkR5pFrBpKcc85gqJG2i6OSpg39b0dBqxn
eHLxCSAlKoRLtDJMBR/KphWNgLedbgDFKwFtzHavrOPUfeokBExknLT1NTmOgkz8
7fr5ybEPLTf8uS9UBFX8TFs5CtAEx5xDYlrz8+ecByF+ZPtloRsKpBP2vtwnqjfu
NwUHS2/fYV3tVS9xMs93x6gxGiLYj010gko/G6xHiuPKg51f/bmgdwMnx4gc6vsa
tMo8KMVUPZ1PG+5c7XlItr9dNuPaotDdWdad62Ka5UeB9vt+wV4HSfAU/mFkSW/v
ibRHTZJJN3IgN4rWkkmQGOGE8hm1kiRrH5ar0yheWVyhCQmh2ye46rx+Xke2qU9F
3bMeDLsnMeKOIg+8SLwzX3WsvX8BXiVJCaCud9BE8G2BMMQkSRJzaZy313KFQIRT
stU2V00WCva4l14tODrYP5Va65K4xjS2V5bepm8I86E9N1UelFWduD1QSN4KCdcl
FkFij8DMfYzrd/zTIQuiuCGgAfYcA3vuNmI2g+c6TzKSEymtVz4lbiOoFyFhYz9B
n7hhFYy1mYEoxmoiHE1MJQoXZByrKQxrww1LAKT5ijHY3eJD9uwr4ql9IW9vfUr7
TeASoniQNPVr6/X/eLH9RAGAN1TEM2cVT97YqM/mnZtagMnIAwWoDIE7MJCN/zhG
u8Onhw0bLKwgRBBiovhpApdmJ9DFlqe5v4Kb4XKBCXlcUHNYCbxtLtnCoavddCGV
lwKr7eoTIfMGnfAZfhzn4/a2R7DXhPBVJwcKXNWX+Ly4/IH1x0VBO02MM160YCP0
k+tYPxUmBeZr2zWOQZH3RdocxYOdjfxfopNe+zUzkUMLStUX0Ol3Gnlvea7NDYuf
5bsyt2BHGL7ihuSNmwhjSqAkVfeG7ZfvJPQCGPlTBkn66UtGGpGBDyGe6WEU35gp
9mMvdkmTsnND2zSulWuXiKnQfION0fq6xCPEQFjRxofZHPb+yoVaCgJr4Bjs1EJd
WqrDUAYEbbfjJfp1Jj6VmVMx9EHBUW4wPR9b3y/bAI+5JzbAvq01liCnN3LTq0+m
ex2O9cer/y5ISGW9/1ps2UQUDl8wAdIyWVJqG3Rc1QRzZERt6w2AxaimxfWXUmeP
z58BYedldvllBgc3RQmikuGblvCtoj7ENNWd+vaNMf1LcWziSzAhOvQcr4espNRX
gpOmDQXI4M4Eqwk2MyqtAs+7MOQBPjsoiqQAE1G+gZaJK0oiguSZNrDjIsUx4/Zl
4m2VHSSV9SN+j9xIfUECE/qtS0z85erFQLFk2HCrMGAuhLtVADQ/PaNvr0b3vnRI
Q1yjC3mIhpWldnRh7FX5TAXCvIlLgByJVgqMoNKC0Iyf9n0arwznyocc67FLhVsD
y2tI/Zbejx+mWF5k2wfZMfAEi7WOUzkQboBSPyove8GOJz7huRsV62FgslK2LMBn
nCd/OBBtrrBuc3Z5Un2CLcT754TFe7Fm8mexWGjjUH0afmdw6Ep2lRkoVJdpQgl3
vnMP52skLtqf+IGU4vCpwQK5k2vl8P6svQiw40cxQo3NM2rhJL8MX5tjJsrUQQkt
cjEZGJGMeMXSxImCroge0H2QWePH3L2orlZKHiUGH0e955mzcyV4GJJGXbzqzv9G
0NwrPCQ40RKml5wL/44Yx3RAg9ONRhqbn8+vMWw06F2MTNF9onaGtuVX58j6xpwo
/ksm8TggPogccgQKrFAtPifzYppJrRSMpWXdK5UE3C4z1PlSMaHkRZy8yYJDQgMx
t5rS30vtweqJ3OI8lBURpvUxJ6kja4zP8s/aK1TstlFSwkNfKGnY1SQtuyzso7Cs
lvpkCd/CS2FjfBU+U384Q0p/kBl6f1hjwASG9DjPrBhhyyr4kfWgMfYBo5kMEyVp
HPDjJga9Z8Djou69JoPwq/pWSoKZlc0lA6ApSN1cZZH4UHrL6nuLpfvw8UwaFWdR
BxhDCHbcAPFFEHCYzvgV7rVKyrQYD4UMUHhotpqfKG6/b+gkF4jTsE1XiDApLbtq
hvcMM+q70tHrbx6QzAqvwsMVTBNnGzW3/HWYVEqtbkdjtfzfmURDrqSC5JUehgc5
OqkvhelFYXgOxBw1+RaMSVeFx682OSL0B/uNwDILhYBAWit3Thdr+M/kf1yfFw64
kD1poqSi19f/v515gFgCLB+ZTA3Lq3RhA5BoX2F7paj7Z++BqXLjW9IZIPVgtC0t
KmWRz3ZCjTEfl8EVz7dz0uRagHHf0isvtOnMHTtgaQDSxwYcqSeFQFSFwxHwOYSr
3Rgm0XPFlSV7zJOvCeBzVPw2SqxRzrueEA3B1A0aaOEUriwKCvnRSe6jijhW8BEd
RtLM6pGH7j+LH2uM3TYsWCw5PWLCMzOj/bs0mTcDLHB8wy8MqkM2B1EREJypaqV2
V65czZvDb2L2ms3SKZeNNWY6BuFyeyP9GEP7Q/Ob3GFk7gcQ28x2AIXPOw+hKP2i
0Ycxxs2Wlq8ghUn0XlxlTY4J6F6TEuNwML44CzPvHucQI4EmtBkRBTsEmOQgJoUp
7BWCGZI+tsuTD2U9jvPPmZ8IQNmk36RXd8ZQlOCdDViTeisCFcQXDA3koHvDWDmm
MjNtMdT3iRtlTuFn2tYAWrfnPeQKJNW6kMw/kbU5CbIrUpzxq7sg+vAQ7owN/n2N
4I/AWyomXzDSDwosW1KzCP+HAs3zPwxBbXXcC56XxilQ8ZyWhGH67T/LKKyVXEZf
lWiAsr25uL7hCg3ETvwAX18NV9KmDb/wDna42E8Xg/lc33jYaGUQItfnLXDiARAx
dUHQVHN9BgcHqJrUp2Xvhm8Oxnz1wLE4VwNqOEld93BFCj24ycN+sHKGFTRBRVgF
x+nFfBqfzMtrl70cziYbNTfoHJhcUjrP+MLKJWuqEDQwOzU/IORJ6WHnfUVup+Tf
Mn9NbrOffKNZAo3F0XrDE4sbejCSEGvrXjSoZsyTMrDz0Q0O89c3JQz3dKXH5yEJ
DeBfMfXgTtXjvOPxDEtVqdZmdLWvsK/lSUaJ/qhqaL+dSK/QQNP3UAPmizq6/4i5
5/g4NAp3rwWyC/zseGJRfKc7cMXym35QelAOOcYuLcq2Tn0DIhSll8xn6U+dp/CK
g5RmtU0ryquVn8f2rWrF7sYcN5LRRigkTcCmcp71vA2MoKbdkSAiboqolBUHV1kf
UmgNmFpgdM5Mn+VUatJspDwacJufRQtxaDOA81cXH3FmbE1kqC6dBob+tLoYrrvG
7Ac3ide1EoUnQoVsgU/4UHua23LGv7ud4bZon5gaNAspJpHlYhQbJWPEh+/0eHcw
doOLfeYSdXbafJXdLcX2X6N2Sa7sec+LOAp2jqP394+6LjO8WaJpNpFAiPI7piox
GR59t8KwvPpEd7hMz1IywyHVGVa53rmQYDeHRrxPNgntWvrscxW6pzpW8TuMjMOH
UXR+rBErhQcjCYAreVOlmWgGI+LgJZ0hMoTEvM0d4JpwciWmC+GETz4B39VWnGpD
mNEnpzSWhP+9t199yCWWynF3jq7Ek2B+WZq3M2r4Vlld9rnv5Gtwg37uCBfl/n13
URjLmzX9PRMvS0QrXR0AmHJg+WSeFLTTReMe5nLXIl00roIXvAcEZx24J0tw1OdD
1RvkNOuOtAn3kkkRw0V13SCOq2DRDl/pU6Tiob0VT468dxf60qWFGixJ2EH+rr7a
DqbX8RCQqesfUNtPTXMLoCgj2OGmN1cQerMvvHdM3aAINPLr5TqO3y4eb1qkc7Qc
qSbpGf2bxqm3XqDONcX5tkVWlLbbhfR26lTc5/1qawxDTe+EJzO09mKg6whK5BVY
8RVIQoixTKUIXJa5yl8qFB8pPApxRqNhQTOLPVwoKpNB9rJH2t20mFpABPzQPRNN
y+bjbXMyQfO4/N0ygIRR/M2CpQ7Nj9iomQ5VkQbIe54bUNuVzNkOM3k7C0OPXXpM
Xir8ZF3X1z8EBTdVkZyff+8yoGKMf/tD44Ck6g3jcZf/SZdWIodA0X98xD/b1LR8
I4P5K3cwax2mYvC3n+wKj5/ibyNq4g+7s6uP7oibfc8Kc5bzsau8Ypv+UQWXQ7N2
IV87P7zcUeTYUiRWVt3egE/H2jr+aLdiLwx3ipU50RmnnLCdnVrp02HlR1IeU3Jv
ltN/KcDSTkZr3JxwgBE7ItxCQ+pnZJhOVCbui6gHTJKuyIMrmtQYJUFuVerBEjh4
FKcU7ujTDAKRqhK0RgFe7aP0976mTSaTvSC22xdueR7QwqChcbt2QwhPsSBi4sAb
7S8XS9ZUj+Z3N8H4x/uwh5Xe7BMwldNkBUxOy/X/hb/efzjdO9ob/uOc0KTzQM+2
SO10d0022vBSXCD8lGo0nUu+C7omiyGH3pQ/v8wybtIttWSoYM95faNgs3QEa9m4
zVNCXZznCk1lxxXN1uJRG6Dugc6bTajBCdugOv94H6WcZYiUc8k3ma9g5cfP7B1r
VIvJ8b0J5gBOwMX/UurlAaDd2vU+E+KR/MWMO2GaUpzjtqVnKRyCfmvJwKH2JyXR
DEAKBe7fD8QTY7+nI10njUMyhfeHT6ADT6Byr2I5P7x3mDoctIQjQ0se2Jzw7E/W
1yYmNwFbY2USbdOhwPw+quRT+6csrd7jGqkSw+wYXJL4kHkz77BQ7+jCkprlj9et
H9/ZW+9Wdu1hfGRHn6edzZLcKRUHSum9hfN/gI71KasrpyH0BNz44rZDP595ds65
sksjl/cJEC6Jq056s2W9yeTCA3TWUXvI8QIH8oboxvFZ3bhf75kAN3I8DnKoCyy5
mlFUo01BGuXyneaZBPPqLovfdXXxmEbMCoSQD3xEf4B+u6+pHrs17wuU4xe7VMWU
FDMhQmk153Of6FRO8PiDMPkVUq7HOPkB9BS59tIFmYS1zuucTgPl3YbZbNGhdocZ
xyToRXQ7bfK/XESU5/ye6TteXYQoXyFdCmCPZ+utuD9VREDhIThTbvqNKtoPrA9F
sGH6tpfT1K9uJejJLzqRIyuuf8ViwYLd84FFZ53OYilzXTrNBgqPM8sYQxEad7tO
e7DcVowfB5A9IRxtAaiBzqFQZivbyulFx/Va7nKJQ6A2tkkUNZCbzefIM9tTwFsD
cfFbTyN+hEe5/702aJ7GK5nPoX16YQ6yRFYnU5Cs2Z+JoWSNQiD5kFjcuOa3tzvW
fv07wVeoeEnIGAW2Z0PlD0QdUitEKIyoJ6/aFywbtX6LFGYdI1UxuAVVEZ6PlIGJ
cAX3wShTitMlRQ5B0fDixAxXhw8OQysB0GbUAbctqS9o7ewufQHrbtBY6Cui0Vuv
WDnG0AkPe58/ruNdDbFZJYjdLFQQYcyQkco0Rd+IneazGCyElvfFR6Ejjzeb6iE0
kJAkBK+B6mqaA78JerJ+WfczhCz8hrAM24P0UJoV3kfuHQcIh2taNDE9zCFpl/zD
cFT7SY8xnL2DRREahqgAjlpikbJ/cSgl/L1sX1aCQHSIa60NVzqOzWVZzCTlIBFa
brrB4HCtSCU+BvF4TQ654o4ALf7SCUVcPR5t4hpW8jyqDxJunvUNSx0JTpm6f4ZC
8ilalIAgRD1SqBO1KKkgSDDbp8CsQS2IOQoLQtk2Xg/DNmWLy6bJ8+2EZYF/rxvd
320n+Nl9Dt+HgcYTsQYKmL/A4i1SRMOyvogFwmKiCZsBaiU/ZgihNyBd/ejFGENu
/FLNeCfwdGn0//gQdDApyFwYDgEHbyzCOh8xySaBrQoX+vMPtdIEtuc/bQ0CB9rq
L4lHVAM2itdQJyp9/fyUD7NVe0D5gJdyCXaB0odCcOPgfLJ2FfFLWf1azAZl93Ar
Dc0qFxYV6izFIhCQi59jBtSwEW+3a9yoaxYTS0/UIxFSM6fchsAqfnCjFPVK/4/8
geexCryswfA1EImMtr7e51Xg3ZVK2JpDeCYNxeQ/4U5ZVL5flQy1PSaljzTNJM1z
diCW+QYgbWx+/GgR3fXFftQaLn6cGka4l2oTkZ59bCKuwRZAGxERe6rZN8iMfUvx
WNVtemLoECgT6tpbiNnIFfN5lfljg91JvD/NxLefgpjfMeJVHT75rfqwqkjR8Acw
wgoQkhmZmcaz9kn6Ea9LMNKFifTI0+kOS8sgXexSAwRL5ezjnP8fNCm1APrQr/hy
xMQZn5ggkxLMxrNI0yhnggPtGFRqIA7C3MzZc/Wv+oltrFnfSXFxMKN4xWbAeQPJ
qHFE5ak1NWWuPx40nk7rcZhSlcJ1r1XhP8A7y/1oZmoZxklFBh2/kScAKpQzOGaz
gZZ/Hwu5CFyMyh1525ssKYOXpSD2zDAGwsDuYWsh08DKWqE+aoBbmusdhnyg/U88
NwwLEXM7gPPpygtTegAXRh9l5p8oac423Or68otUJTCL/r45aqFmBHZjqyKISkF8
82upyS2MZ69BoxZH0xxn83ajnUcMns6hVoqtxYKTCpTVf33g9GL0pIY+8jGbrkZ/
fzjlz+/ZatQaT+8/ALyrwRbZrDj4xjp6Freo/eubgLYy+tCQrz32lXj4zW7W6FKd
64VqKN9emC8BVDx4YoTCdggdlyXjyICvF9yW2Qlwhh4Bm/3aMKCQih4M3LKLDfIR
JlrkP4JDvSdLm8+0j4T1/jZO/F5E/up5hRGTM2riNFNe9pkWT0u+LsUzspnHJU1b
DTfxR/oBpiiiycN2QUt3xoB6m9jPwT9E3OkEubOS8gqcUoqbXXE7FxwJ+B2e5SKV
bM9GAP1d5TF0kOCWWlap/fQnpKVeotltv/8VcrdJ/nvKcqoiz8f3V6vaCowz/CvK
R0NQxvqZsr1VtKqdadcxOP+nd0Ncm/ZSPG/s9L+CcNfrD/KVJtJAIExf6nW3g+2+
4wsBdDbYyyGw5vS+4CWDLren1bY4EAIqOakUc5cVVSAnTS6uLMzA4HUElm8sW+XR
y/deTMUYxjhlcVYjLBkgcluwT9IBG/Ct9+nssRf5UO4u7ZbcVOH6Ui4NSN3c6pQb
43F9D97ZBU5uudJtBMJuvDDfXpRmn8/e2YdOc9juUgMS9xzTIjUQ1GsjrFBdNPbp
kdIfvDI4P2GxjyeHh9SkAj3OsIYXvvRfzY0ZqyDVC/jj/vTzd1ukQzdGzn6E4baZ
GoKE9IMr9jVzRExgR1oVQpX+mzEFmJpXevZ+3VmyilPY6fxCaFIlrRjjJlMHfsEY
RwSD+AYDFX+yN2K9y1xCIvBz/QcgiMnrHOeP7QS6ctBr9mRxqByeSdHoYzhN3H2R
7Ca9k+vOi6WNwyt+NTNpfAxxyPP2P1wLhW+I+KGm3Pft5dbOqkrQQ9JJ24w8Bnl9
6xSJf45ZExiYs3FOA+cdRAPiRJMx7i6zvFbUR3AsWVP8TwcSbtyWyNTep0Y8Z+ph
oaZ+vV5Qz/2WdaiOrGqjDuqsXVyKNtXEIU0be5KlkDEeyNL33WzMKFanf1V6+Alq
AHZdclD1efcenxJ4buKh5Xqiksy7lp13ds/x6Xs8LfimZWz9QPfw/djLeONwn6K5
ol/mTYD2wzULsdh4YXUNB+bQ0naAHeeFT8xDPga80HXnhmsTK++vvbCgqQXQkszo
vYKhlQVwjh73O1kDCy2NITgQKDM+1qpGAn/nOFfG/WryPkAmS4SFOQliKWaKgQ3O
5aTF8YyY4Gki2gfQgjgd8PS+6Kq65Jf05InPhz++3jaaho3Y/JRmPE7Mjc5luBgz
FlrlWvjChjx97utQSLPEu/J54ZbHxXggk1zf5rBDo42eVwg9XC0ffDY9NhnDggIf
K+i/PTOu3skkzTn97ggt+KIqRCriVTaizT5W62nnWtUhyBpSrM1uMj+lUhXiyz6c
OTA1WH4ZeS+vSGkrK4fRLc600XS7yHhBy97Mk2vpn21Ano9wq2dVQQv1wAvYsywd
AssqXfQpWLHNulPZ+CpXYh1JxRMaEiey/Oe54krvnVOYyAtDGlVzPp5VUz46nZzD
QK6hi133ouRezOrxBo+D+UIyVTI9ewadE4KM7k2yhhj1hMRMYY8Do04mL2uHGQUh
aEQMG7n5OIvwLHugKLvbkiYc2A6SF3h12qq3TvytHWqVFIx2sZUU0KUL6rTPO+z4
T5nzk7Oic2ZlZNfK6ankxqRqD04f3PAs9MyjFVeaIWoPOc0p3JQq9PIl3JDqT70m
UHprIGEWsoFESvTgp6gBmI1dPEUhaMrmrh/xguJJp5hLS6u/HcHrIj2jFI4CUjKm
NoNX4lo1NI4mRv2i8HrF/kUEpEhJnJLj3tLTM73bmjvv41bazAyz8/FfE/JAhOyi
PNFOGvgrOLmIYvB1rL1tiJTzSLi09hCho7wAyhFEOyv3vAq4f1CzJNrJudtlpBPg
7foz/ud1s3JEyX3+NV9kan+ZALRT5E7wUZPmcwFBuyOPM2gdiUn+6E0lscfu6Ndr
vKTzLxUK0MLkVnF6ySy2KkBLslErOuVH494fVTULQGal7W3MS3ur914yfMaRZuzY
0xAPSdstGtcHWU0if0so3rlLIa2YtYHZ3lozf+stzR3ViEQqygkOdDRnq+vOgk5g
3+F5/SJGh0JE7mqCH2XK+ASJvbeFpqPdxAmbrX6imfiILQZlpYJ3+6yjUz2ULVsO
kscz9uqKJCHH40ADXEkRKN+ePNg0JT2rEpwKf1Z3eqh0Rr3uemcW0+tcw8mPX1WL
Q5A5L+AileF76x5dnHB9vOkxp22xqNS1qtFpmBN9xFkneotD4aMLkdgjB4LWFDqe
sdWmk6fmwMuuUwhQFfy0wOxmsQPG2gLr2acC/DMgfqVNr2mnbSWJ+kMQwnrdqNi/
Lo4+8WcXBRSthsBPzSktytW//fi1yawsGpaMO0jVtmcDh3bHmOlDMWI8R/qeNOdP
H+fhGueKJAa2drCLtqXrmgRfGz1jsGOlAoP2ZoRLSbAlpwNnxK89d3unUTCTmOEO
A999dgdKCnQVPr0pcZnVobL3WmlJs4AP8U8zRFeGcwOZVuP/269oHhiPEdYRz1xB
G+RyATr+mLuwvLB6TJltfso4WkA9p6PN7zzFPRykEZpVWqxZzTGuuuUjYTTR++qw
oNgliIvPZHf5fnX1wxb+/tOVtycMXHMh11sZObCJcheA61gezMFQcdzNaMpWyw5e
rHINItclZBlGo/yAAT1214FpOo92zK0+5mRFe/u+ymZXzpKOjEwh6HgFY+Fxxv8c
v5LpfeH3qqocTf+Mk957ow6XYbQ9DCnbHeVxfZG64RKPXemWFa9LDbkqrt56F2Vd
6xkTmRQsblfuf9OZZTfcctU9LioJH8hTUho3xxXaVWPNJuxWbUifyG7qaJ0nMo4w
XQ3cWQnpcUmIX2a+qA2P89T83m82dWjifxXnpaES3YbSdYHTXicCRCzCNNhTqjxa
8HpSVcRT3JLhHXkdvd+mKRETFwWMYfhsdiIp4pdRLRIRHeG9PjzLa95E9wWl54O8
s79kGr+U+dkwD5SF48rJz+4KVu31mTFqSv+uxzkxMvDYyWA9Y0PBAjOM7VEM/rMo
IalesC+c7w7WGTIxPCYbATssxQnOijlaKr1ZrCKMHXEdVhyenOmpjfADnHM12bVd
AwAVge3Ln8G04TXXuGdMruGmi4PFMS55DkPcZf5g4RqWr3H0SeeH82XgFV67ZG7T
m1rV/BRPwZADEiihURStWRpqawOmJh/uH3mec2we/LRYFtiE1YooMSHDSUU2KZWk
eVthfkXhZOKYHDMllked/XDC5YzL9VEy4lk/dzDzoOlgmnJk0+/MLBM820foHRp7
aVd8bBGqegjeCiZj1uB1XLlYi0BkzcEy5JZxEJ2smrKnnzTy35JciHkW+oPk8zxg
Umg5iuSxXH2UF1Tf1RAmDvgAFeGd8doq5a/AZjx5pWrjGXEoSQG/u86i8DRnoBkv
C4hGgM8S0eVBpIeCwtRSvgRLD6KLE6pLb3uAjK0qjXueDZ+8NVjH5EcOgl/9x6Zc
bGTES3K5Ti2kAEUup6DpBLqL0U3Y9rQN/AyHOGnofCY2UmQ6Gt9wW9gbC1GLUve8
VFY0UpinOqzxzY1KnyVuzU4s4Fuqbpk197J9P1LdGyP3W+IMtTx4oU1LndH1wjuD
WQv/gU0lDQzBkjCtTPdCeWBDj+1adIQ0UkHNICAGALr5rplU0YmGXIA6Ii5dNC/U
+b3uASad8TdyVWYmSnz9sJl87hB2c1hINitr+NdDHL+4c+ZoEM4TPWBoGpTqCdMy
p8okydstebtg2FBbDGirkwxr3IQTzExgXfct+yLtquHWDWUdQM1M9CW0URv9isw2
PYwqlnGXD+20A8sgAISWtN/sf3WtnE/GEPGYyQ8IIsn5Bli7usgFIkmg9FGXStm2
4X5z5FSnMMnLqIj7exm61PM3/XKNmbkkeNKBTBRRSHEPfqIhRQ9pbEA+G66inca1
8wrFXowO/tZCJK+hDFdAXaoMtOn+d3WkQe2Fe81gqmpROp4VyocHvh3dWIsZpa4W
doVd1Xnxf1Td+b5arSn3XW9Dfeq+KFZvUEImc8As6hwyiwrpegP736zBt5qGFcOk
4fPhTvl0Pihx0JNFgqz+Jl6FatcV9PmsS3USmELeiEYv9IyBsZw1tvzsq06hFWFV
VVkalJTIAGqvg6ZHcEx62bHCWEPnnwda6QfSnPgWoCT8x/aNl5Jw8nDah9oULu85
ZVrG0cnaFE2mKrb4jbVDJfqztiJwysS4bXxEnfhI62Lgk+YFbGhgRp3ZEpNuRVtw
pjLnMThV+iY8AJAPsky0ToVwEIn1JFK3p3ZL5SuJiZoBPEt9B5SnNgUPsapeJzhI
LxGOTho0bQteH2ALUiPcUWm1FktsT+AtRrRbpExYzkOWkiYOMWYETkaVz7HJEhOT
AYfh94P79BSXWlx7WQ/MXRc6M6bHxXB9X6NRumCR+9aUs3j4NOCMaakA54NzMNer
LS7DbcMQqCcKwPywQMqZsaexHU9NY6oV8lxMjuMRUjhtassF6xwUguOCuR8AkOMW
/IGROpIBa/vNxOxIJ9zAwuzJJtJDNr0wyALaviAi3xijaL98/zNTb7gOm81GtHF2
JYqRYjqYyARIwznUmxen8ph1AYOKvw7/K1qf7aPlymH+KrK1Xtbw8jh73Ge0PK8/
B7EGVShCgUgZ//+j0TnCGs4QCKq5LZB2MqlCl2hKdDXgyBEeAB8c49N/Y68wxU8j
Pltl9c1ouvgMJnAs5hZF47LGiZs8g3Cdt1YSio+c2DdeMMb9jwKJXGkeRp/970cJ
I5Zdw8Um2xIid/LS3FDLl3xu+zDpEeTx0i59GnY/Xp0lm3abh8ryj0FURYAo9NTJ
G23zBnwZpDPcOmaUuXtmvRDYqL0Ai9S0QTVEZZqz7722vPNfQhK19Lm22oTKN7zn
2Uyu2aFHc43Jw/pVO5wZVvSbBc9+v4oEnSepOWwGHuKpnk7b7UwPKoirx4DT3kD4
prqwTe9AdsRSmbyGowWTpvsB3vLhvIOCc6KgL1SkA/PhA3CiOduGcFqwtj7n96Xf
hb1xT7BL04ZCNfzUyfv1DrCw2BjHv6BpyHoIuVEIhhLh1rR/78Rgd0QkhMhMX1N8
3ReMR805bssqzyB4l6TzfTniRSc3JHds4gUQ9Ve+2va5RpP32pyeX76B46In3pTp
VaV5LawuWVysCCzddX17lZPYkVuSu+mIiVlLxXWr4f3ajbRgWJ8FrbmMkhsrK/fz
GeizYoc2DgnnaGSTtMlyVQuLocZq70A+jILqgI/QRqGHATJH5AibWjs0+pZms7lL
dknBXRBxXtSavG/OnQtW8PDnSsDm77MJS+QkcczEahuiHZdj+198ka1JX4Wv9vQT
e5eCylK/3nv5D0KLR+7EmXOF5pMbuUvMaXJMIQ0GVBV55hD/NUJP2pFcWNNJC+ey
8MlCznpA+4/Gc1TXCj34ql3O4elkj/vSD3SLdW0AHWmV4r2O8RZzs/kgPu/fEve4
LOJuay1QXayVYPjCNmZrP5GSmDudYg3gQ4Ct/AxKJ7Bt+Sc/HumqML2hxreeLVqQ
JJw0PukxfvxaLiQLRER0P0Yfz/E17uGC/Ce6WKA3gVVxZp8nD7Jp+p3OJT1G1wwG
kUlgSkcA5woKECd2/pOnGs7I2ct6/h9NHO0d+jPMKN5LSN9FcyF5CyX/tr18sXs2
TBCEPqMhhpHKxy0a53diFsDq/0bkbA2wJueXVU+Bbym9Ix42OqX1kVgF5e+jjhQl
IjkbHcYZKAVtKLynina6r70Z8eegmYa9dXnj7RkT3FAW+GGuy0kX2e2j2V2VUk3U
pysGLzK6K9ZAgSZHSesHFtESU8MSJtKFHnjAReuJYp/z/fzIGWa98/3KM1LJrSQS
i9m4be5og40Qi4qEImCWG1ChhK0XrWSh3f1Nyi6izGzYj2jupYXhlnjdDw+WJfUi
zcaLQOm4/RR4rFJbD9VTOLooWyl3m2IPcjVV0a69Oa5mUJKL74t40Koksyp2LsvN
ikr/d5jQybfm7AY2kIicBjkYBtTZTk29fPZWdpmWD9UcnexgHpEstzgXdb3c5jmS
ZXqUMwq+2Wz8JvrCwdSCJBj7y3fLif6NW2eJhuv84EvHpFvp9QfkXfJd/kz3ZMBc
BiybrGuKJzSvg/g4YjSk5sR3Z9UeFlbkhxr3ISYpqGKo/bRgGzwUBquy58cuJwhM
q/f8b6ugrc6kZsi9tbhcgoEXvFpT9v6mgVf5oVcSawDbrtWMkx/tW5bTG/jnldLP
Xmkqt8Vnb7rYmIv8XhrcNvfY0mLWdmPtWg4NqrkPvdFE91fhFwCn14VZN5uxG5z1
hrbpHBaL3SN9hTaZNBCJ+dSTu8uKEc7CIdF4kiLNtfpR5naiGLMJDe9be+n6USwZ
C/i9ieEmJV+sCZaF5dK4aRIslo4OkEP86CqmZk+SPkPEQPcZBLNCZ+/HJmhTi4ou
hI/j39DU7VYqs4boh9LwDH1qlv5EmIDFxVlGHoYlnZzW+xFtH+t4UEsJA1nrEkVB
ibEDab4CsyGX7U7V2G3FASbnFcU8VMTkGElnBkwZjwKsS8CXlF2bU0JpYPVgjvmG
c9tVwrDqaljfE/dnTLF3ClNSTDhK0MScKBjI2+WGG+9ZC79h+VEMBZiNAT2WKY0U
ly+ZZNySTjh/cs787Qh17M40szalUZbKzqzhmHWR7Ec14ZTP4fWk5Gt9J+jlCudj
cbY+d1uiWO5hs9FGHp4COnaGY0dLbITS8oVmt4ATgz32Gk4cu2LBokpAG/OCE75+
spNndKToTZZ5Sef2Tj7DU6xmo3r7NZHTtsBtClBiMpmQBvkZpLtsdS4/GRVkRHvL
b4uE/b1cjpYFlZzDaF1LnWAT9Z/4dijNA5a/bDRqszbzN2PEdiiyIjxOwtsIqVJz
Bq2UazBTwL9cpapxwpxKx5gh/aBYu7HpWZ7gaXjAZ8fmiOABqRT67XYrN69c+nGk
/JJD9/OpMOTe8hzXiWlIS7Vg3VUWgE4m+5iN2vp7X8IJo/gycbC2RrJk+p0FJ6Ef
NjPn3Fe+gU0Ivx037Zi+tAPzFTm9wkE1LGFoIBCnq1oQxj9dSz72pFp4xHFjGhhT
piwRZGIMgdJtb0GBfE/Gt1/6ctmnkr1i+heQu3Sdw6ReCIsyM4CW6SFnsNYsE8oq
C55r5QbXa4n36q4g13z9E5NRT03HCvymdzY5votrhzNmNiBhheaNFPoLg7ix+6Re
rmOqBh+ftoX68fZtVrkGZjUn79i1/eaJ7SSIEHfxxq6om0uTurV8L9/eLnRatUZO
X1nhLMDfy5QqAFwp3tjUc/cYunSotCKexGa02unheuCjwZwoM5WYVu05dlXA5S8a
xaXCdp1ikyh/4p7TTgCXD3/+MmebsA/mSvwUc5zjNmJexuPN6ZSVVppD+eo0VHVF
kQVt5PPWN/ztnyZo5n139h1KXbfL5xG2KS8rRZbP0izX97tb5wK1iEqjHQKBlclI
h/uvk6GkbuRA0jFovfVnJFO4E+Amcbi2pm2uJDVW88wtBicRlhZC9HZQEs4tyqlN
zv8QhN38V37Ihc1XU0iffuKS+EXjHAshYpTQdPfyHR7X/wJZPIQg/AGj0WR2Jwsh
cPtIcANXsuaNh+1mqev6QadhYlsVIyWBo56Otxw3eoEQstspGpqGmWepWjxKPQ+C
gj/970I/QC1ZCHZNi/QYBQhegby7misy56LqWm8LmYWJAfWuyzULVL3oP8tkyXCF
OQuRiQqR14pb/ZGo9C19KxYUfEbJtotI+MNtPEA9F03orPvYhiBnU+f4Gh8RzCRQ
bR64D7TY5WxAXBYOk6rCccdSLDmCBZ/iIXGH8djtsbwhoCi9IbBXgTk28gFpgffv
nfbtQsknYheoNWfuONlBV7Osmd+sO35sCIays/7ElUAxvfMnSEDOoxkR3+4287t9
UjQNfLhCeFfeckBxzfyYcsf4wdGs30oBX206O8zykVR+nLO/mrqsualA3K1ulexR
APCeheI3PXs6ikG7qTuQXveIu5wqT1YVt1fncDjsMOZVXgus6ZZat8G9JulLJ8bk
YP+2/rg0cEvIUw3hkj1vIaYVghWBMPQ0/P079ulfQ/2G7kKPrwXsKtp7qDTUgjOZ
n8lJ6OnyZc7nnhE1g03AD24iawmdZKJ7S9mzjO7cjwH9NNQqjGVlf6/+HF7gkMf1
N0dUA1+9bcND7luW27+DwvXgizbpsXXl8MyfRexqFGW3mTruETyMLb/6xYZ3/+OD
yQ/dK+XeVVQXYfckH6e+F2x/3ytKkOWEiJL5+nlH7sY000ABcDzNMiEHSg9O2jpp
Sng/bKG4OG/GDzAFHf6QepopZ6PGii7uSzBcWbFmL+Q1lzkUU0ruTlZbv+L82cXd
QPQKTVzkjLMxo0Yut47J1FrjzdneIADSVet5fpIPFIkM+cTguKCVXnyP76ZnjVc1
bjBBrUWUaThYN1YU/igEbjS3w2TOzAya8sl8M43RfZoGRAfKBkrIXKTIQWYevwOL
RlE6nd8c/i1KoOKhfeMOvVLIaYOOimTourXu4GznjtEOLEhO/lrvlP6PZzut3RYD
D4QO4r/uDZ8ksi7NQcA0Q2WIGPnJum1cIHz/faLr/D6HAxD64gH/G7KfFXVe4QLK
qMcxviEtj2nHTy/2ODs6O3zpZRvH98WrbcdRBuvekJFUReBmcxQBaXWEwlcwVVXD
dtwgrK8a46IOd5q7FEBJGix3zFmgneQuwq01sok6E4JR0rGUFV6jgP/9tjOZAyHr
15VYE7eX0XvENSV5UKLrzV1IzconBvOKN/SELKhl1oqA5KGL47UFDeLmxa0RrqEn
+siLAgktpVsmMPFRIrP2oJpxaVyfLVO991b42OKGhgd2wnp/Jvr1cykiRzv6Tnw+
VcWWdHkEQdw0Q7WiJ99TNCTVOEwE+tP3+9rmG9wBIh09qBJNcT3BC7NGfMxGZiXb
2lBCMoY5qdrvo1olwa30G9NAjw4ou0fyetz4PnpmmwROqWhEtiYpISQ/WlZwyzEA
xyMKHSjRKCEhNvBsfF3RqEQVFK7/ikwL5oN0kK3UceeiFND4XTnFPjmSO5y6QV0L
/jqwf+o5heQSKeYRYhPRv212BBaJFolyvV1b3IizXaOLzdGfNncyfelS1vGvPjOU
nRWWI+xHh22JdEdNqaJPPDKNuqcU9TwLUPpEw/AllUtynVbrTBThCImRPua0IIHc
DYPnsyWMaV7TH8PT808K9qsJwT2Iviby4Dc3FV16PVlGZ4zau/uludaLSx2NVpht
Z6TtYrjJlQmICInUBZEFgdNlOBHBGLOPRA7Gv7pl5DFhcCCjjpXx54iL0HNVIBsj
mSVyT+GHch2xlwJ9ZPsCfRXqGL8oaN5W56BBIG2fddUglNlfql6tQEZlD+jTPDZv
qxUh3yU0hX8yc81FjBuqXffcOvJRu0TrGnvZpXQHGFDK2cprRUEPLC3b1pNIIMmc
TNkLweha4YWaEybGyKXbzBSn+v2ah06RzLatf2/tOSJf7hqiVtUzPBfvH7/d6kal
LtA52s4Sfc0m2bCR7OUav8h2G2aq3AhNwHfOUGj+IiYalO8LfB81dRIn717LIdvu
xBsRBEOmdsivI/81XNjcw+5nHjxhq4c4JigrOPcgSwkjsM8mW5MmXSY6D7H4v2jH
2M8V0T3A6r15kmFr5iJ+693vC95MpYqf235X0dRcuap2No5l+MhpoXWeTUlMzdLM
RT0zgWFQC5qlKnBsdFrJ8Szfr0uBQuUhvxhojmtZsYO/gEYhyzAEXI+JPNH3YITB
o8Bp4NSzkmRvyXixFBqFUtK08AR0eXvawxyaep3oUUoqC0jFdOPLw8Wu6/iNBM0r
FYuEHRqtP3s36dyMKW2Sy2ZqWOiqnsGMh5jEflSfVz8R01+79a5S+Sjr2P2hk4ap
VaN3Q3I9VhcXR0PR58qDUx5fBeGCnV80LsEiIpIX9/C7Q76NlmoKmOhgPWxrDe9G
05F/2D2jifSZNDYdzkOVwB7ZR/BFfoH9M6viXdD9uQE9tBzjRHYTjfMfDnooMYQW
Rtz7XQScLwLZ1K9tr1Fn2NfJUKIVIGrHohzDnLt/cEsXWloUlBcb58Sb6njjH/tu
6UGQ286kO5ygWtfRziJ27JhdwPOwZBi3a8E7MSszsQFmn93Sqc6p9kv14G2Qmuf1
8Y1W/pa3wS97tVzEsnZGlKVXaqqji5Wy/C0sDViD1cQoYIRxfE51nqtnySYYHegb
+muJD/iZA5UHOjdxLKK+fWDFkuW249hnZpwp9pP6HXrUqUU9fJyaVbdHdgSb8hQf
9+1rVE0tW4oUTLpHX6u7T6YDvQ/ZBPHIUg1pQ9EOxAz8HdPuhjxaoA5xTnJteX3+
xaCwRE+aMm1yIN8SmNgoir6sKbRDSECqkxVnzsxf9D/icKmba3NPz5l40EuhGoMv
qzlIO7amgoynhsx4lVcHOiPiWfeJpH4n9NJsPfZiL2EgZzG5vS0pwZtJ4D2FN4ft
23NCd9NkBKvePZrXT/dPbFO6QmnFjgnjd1FrT5YMXgAyY43224NbQYk/3zm2/Iwf
Z1svSQppWs0cAjblFG/EF7JwvWPpZuMGKv5iOKt0NOJzf6UKdho4iSlX249ZcZJ/
9agI8Qj+QyJfKWFn9C7I1Odcb4J6k77NiFM73QPSL8VMYJw5opVWanwf4w0SgM+D
B9YLoE6yQ64PHC9rS6i/mkNWAee5bHKJvI0yQUDWR6IOOy1XeDX0LN2HC/yLzGqt
BfZwd0LI6Q3Jk6rtvaeBWdoaiNKaxe/hgT1acerrGHS3V3zyn/25UKDAYXOhOo+/
Ics++l7Vfw1TllGd/miXLyUZ4KtuLJc4AsEphxIlnXm2Xsy1TGyRtYk1Q1BWzACO
/k/zfp3ZCoTSBA1V9NGBb17yX19NxpXuDI1b6gdH32s+LNNGG528jRbN6iI4zCHL
qNOTAFhnS/mHv6wvaMUbqJPHj0YIekjTWjUc7tso0hqvSynoL6hAfaOgUwkfyyCO
cWglHYGXTIqQtTYHt9MAafCVvctRsTs5s+05zxCNXayuAxDxQlxa5JoySUzlujnX
VT5mfK/Q//NUD5vZaKfAwJumzjiZ9RWlF56paG7MaPFWEIlwfqVHR7gHGkS5z0Qb
6Govt068SoxLC8omCLGlw0n9InUEMZe2tBVb12tTUXeIo0OxeNgBOhKOcMWtJAFs
6KyZ+06nZxBLjHBGoPCtDZnEtyaMb1+ZTeWmw4pzOjMla/qLenLmnX1zFKGttOBa
L4OyU9k/bN3fKsCwayTLxvIVWjMpldOywqPMIRubEE3d7+y9URuR/L4gNFtLlDxk
i/NFzSSXDnatV8fh/Jp1VqqmhrM59U6w/9IZzwnlLvBNxFHJWi45vtq842+WuUSR
FmzIDLITbSOIqpKpdowPhWpMx+ZIt/1tvmd05ZwVCLo851Xy25gsch1U8zJf/Om5
3ud9ZNu8nj7wW3dqVVI6pJm9luCi+0N8vtcsJC2Rz6PUHHs+QlKkMCDvuiUsZnms
UKt1isxTmwaAVnLxUoSFhFKgJn81Gczr2lfUEunDByOiubJZEJ+WJgCkeNgpuiDZ
PNlxCrNonCbg2oKXfECne2dykPXIJuSsEl8AjyiFYTv4oB9eH3nOjzOkCsKyNApm
Oe5upgRSMnUMQjjKrsayLSU2mQbRJXP/LvqU1O7SOy8nsL5v201tNX8JKJ4QVaYb
kvEYAFn+948S5netVIN3D3ctAS8FO9BPAWIOEme27FaQd5/Y3Z5o5CVY3ce7LabV
KS345Qzo9ktaD16dcCD/Sjv74B/ylpb3pT+QICRk0mmUzHvvS3iKJ9RsmSqgWeY3
dTLsC3fGy4BXmGM8VHdHUt/zcYPAxVFWCAU5iWdRbhuT38cT3bWxXyBydFocLTId
GiJHBDRarcR4VyLL2rCdq7HuYf1W30O5aAcNwvIeX1VFk4yZz0qOAyUT70XeqAjA
WN3fwXTDVdGgl6eQnw7kkunrbIcAL3JMG65jnSozu8KCwB3JNBFg0nm/wWLvk6Rn
14IrwLZd4NYoy/dNAGzsF86YmzGJiypsdZYE2qYP5ACN6IshzJ0grIHbuWmDmI8Z
4ygSJSwnVEI8dDZF6P7QlYvLrFOC9mpavYx+Or6o+RlwtrKI479Fz0yJ9UnHLKSd
fWpgiZJroLAEhdl3l59YLmRk1l2cFdRN+4l3s5zLIh2etpPVwFJsQFLOWpXtTAD0
68NbV1EFPuJgfwLzzJQVzvEL88zJpRC1v+8amNJcqJRMuE+KGUBAuAEhcIdixNoB
3K0fOOk2MWI45Je48G8XI8rkFvq6T6TNtU5B3DuK5Be7PwkM4wsyBANdaBJ/BLNf
y6iX7FcdpS6zzrXNlXFx3JHDNUYShyJvJv4U6CE7/PONS893TR+gpuedHEeA1Isp
oSHxJMM5JooMuI9pyjyOzYqgA8YcR5AfPHnSSRD4BfmwScTAWMu6kWIfxt6aQCBY
n9aONd5xAg9YG2UcGTr0nWKkpcIlvGKq17avHKBX503cZ/gMb2zcQKrJLjwZOKzy
6JQsfPisJyBO0h3pAjml/0UGjzaUX2D32/0tETofooua/Z/AItj98cygeSyEbLFc
6wEYafgg5IoBHovuJkEncNmKBW6fZiTGMGBhplcUdCaCN+GugOhMHqs2ZRcHWNu7
FJeN8BVDKPzimO7ESF6+qekmoKFu0ZYI1fHI767OShN0ASLf32q2umdGScVJ0Iej
keUh34h2JZN6hvYVw8R2clghSEZU+Fv/zlCtdoi+2MX1Swf5Y1Q53qdqew37SFPC
U35KIZOHngbSF5lgJcqo7XNf0nyZ1V0EbL7au0n9+c3LwXylkkmtI026rMDtf46I
AEuNnVqsEQ55zeSJ53/GoQSjgeLH8llGUv4BvTj0SIPCOK5fbWOC0/omIogqMMc7
aYMw1rS0HBwKqOHO/9gCf/J3c1b9nyIp1+4LLuc5lVKOyYasOKnzIduWUxfScDE1
8xMrOS+B5U/ZAx+6OIAVt0+Dty9PQBBwWTrpVZVoM+RqydtHm6Cb+1MX1PkA4aRR
Cq5VQeHSOjtUamlhXL0++6op6CVlc98S93xzHGhQofKpUnQHpMNzBrxFMXPnDk3Q
4yBCOFTR97J7aP+1eXz/fySRy+dZqGtnHb6dhd8yuW0Hg1WUlRISR8Dk6u9I7R5j
tQs787A73/JyeyyEFoSqRBl1dwljaHmohuu5R4BEKQogYT2V31QyJACyOrRPY/FW
1YuY9mii+RBQTs0tejAumFqVpmUXsVDohSPnghJO/sC2WQ1D6TKY+PyS8PW/1geG
W8bt9aqzqqHKDwcXSyGxy1bDo3ev55iqd6q6E5vo705a7dUgkXBBvVzzxwTHnoCM
ZKWvnO+Vdia99HwYhbHnrmik3YyYLBwfh4K34MSTx2nmXheokmpqJwl+WN0YQezR
uz0emH0nRnGGP9HOJV4kYon9XpIc6hz3UEZbAdWbqNJzT1G3xUM3K6OQV4VLlU33
XZBwEooaynWLZb0a0sybjpnDVOXjGl7xZHsLltMZko64fG2lBwqyWGtnvYnnTNfr
uRfr70tmNe2eH+7Ghz6BwxxW7Pe4RvHuQQgR2vaEsVWNimDNVuYNFVEbdLzykcwu
WyLuQUhqCeAVvSJLY4LUSkqVj38DLbJVxl+dFLTAadqNEUUQkXNFrFf+g29qwdcu
UctnDh4GkrDMf0woFhD2k0ZvU2XR7AFbUsARyZbGtEsGSmXoUy5daEVSW+Sm2PoG
QyTfZgHex2S1tRuwFIzSsxsJPWZ7aXD7+4j1B85tsipeKNH6CckldraI65HHid1g
1fogUPZzBxgp+gx5ve0ProzwPfvAiZ3TDtE3CT3dE4TDT7ZWq1zhHTt6RrbglVi8
MX+PstHK1090VbeCj5B1KPMg+eaDcZh38eiOlzs8mL56wAl/34g5HwEY715BVw03
2FOgLFALLvZP2wf3Wfd4RQJ5QNWyegf+HOMjE5mDmVb78VF2vPLeWzWseJ8vZDE0
Gv+rvBNByQNzASP+FV8hju57ms2l7gBRrS3Of/EVcCpwqTrx5ptWBUO3c9TQacQI
DWVJMS9ZGgKXrDWM5iW/zjvcpkeOVULuIcCyoPvaVYtkjq1e4A/C/02c83mKGEmP
Zpn1uuge77dCRukishhg66zL9FU8l9cSwZNfd29mhxVr9Ye4DGLbqnG8MBK1iBky
wB6DXBsVNh0WWqCrzeSptu9c26/PH1UCogodjp4GuWmMJdv4MyUQvvHyRbKk3ONo
9yT6VLLBkrFxNkcb45oqyicB6aDbO28W1wiwLFE7Zz5t5R0ePCziwhyObClXDHNC
O/vsEyaQv2WNboqqohKbP3HGZ/cFofwXoomnpdEIlHzjNLay3AppGR56cGKeSLqB
iwWvk1zN+GZoMXCN7h8Dz/Q1xrvlRQDaqkGyPxVKpxRlPsH7t/GrTwFsjdn+gKwi
7XJ50+hxUMuCLGeJefBXLKjdE+yyesS/5OnUx6W2KYxSMnB894Fb29JGee09yLRJ
GJB5+5ZnPYnumOnePLCZxk3Va8xZNfnYLcRelB291EAWhMBA2CCRnWCm0gb3Rcbd
X2prm2JNAgO6ueRNKuq1M692oIMx/OQjl4dj2poZrs19XxeLcIFPsCpFqJhKdMP6
scJY59GGudhnMewrjyG0p3/w7oWGST5qc7HQJU7yZCL/yLieuCXETqVPt1eLQ0Vw
SLjmelj5RROk6ccrOMivXfM3natCSmsmMe0sot94nLgJ3eQH8D3NvDVDVsoQOXX5
l8zq68t2J3mtOXuCR72C0BQgvUmlgRdgM3CybfH7QNKWv7jIJbverrHJNiMY1jaA
1/1akBb7VK6cm/seQ/aWMLTrnNM5LZr7oemQYLK7IE/pl4TyOnYBuK3N7S+kmsbt
P0Ej1eYgtWbdDB6wd+ooB+frzytv0ZneTzLLjmsZ7Vaqqnynf9e1G3CpoqK1YVOd
FDjqjhxNosKf6QUPIpsVQajCLv/LdgR8asFM4FEG7AvRcvIb3gZ+ijH1fI/6Iqhw
p66EJo2LTGhR1tJHeSRULFtWD/ZhZh+yVP+NG0qR4vI7nQvOvBv6N+CIEj7ElmTq
gXHt8deFjsCZBC7LyiADN9XM5MCUUE/TBPYwhVOzYtxpTg+ElRDgwYOQ0Kt66YJB
FUIsJHqFWs1LD8K2mse918H+/qLmF2ymLfEDbK0K53q9Jc7DIl8kvpZ9+IsbS10H
ifuYdwfif2cN7NiID/bLLY03c3H+cOwBIaRUv/do42wkyqlCYaSP3oKP0z3xScJJ
XgVv8xgG+bh0KbYcRv6vCQShrgaf6IsxWDIzivRh7j7YQcGuikvEgeG8X/APMioE
lEXOqDZGSkyzih2joRix8x6kWryNz2oCyznMwnjxK0l+row0n4PovTsgXi06zckh
GaA2CVDTTXaC7yxxMbXv6o5QsqZe/VgJHHdmG/VEIjYRRAUHDxlDEnD+lZW+tTR0
dYo7ah1xGA1qo6oIUofKOsyUmp86Fk0dE3j84b0QFTOLdnv+mJoat2yJL+w7+fmL
9J2PEDDVRT3kjglqfYkgEpaIlfJSeKb7eESY2d8OzLXMPXmvvIE9HuHQtgrYu2uP
q45X3sAOsKILLDRXHUw1E4x6oJMJ+pZkzM+7tkn9UmYrlXPpvGhxlbsxYjbTajyz
mnVGvokJYDJDdhmi+8bQMaVN784PHoZlr0ZPoEInzLnHHddCKUg8Hn5e63nNycYd
gNnl5jZjIc0ApvbDym/+oNt7BJIlz2MjMW+6takpmg1VvvELucEEsnCl8LIkkUsy
wpND1YbvhglrglCacdHBo645JsGVTY8j//5v7mlXpzg7rs8LopO7ni8QXEpI0EXH
rEcUgLiFs3ykK+dgyYwg7KjOw4YuNltVWProoGGMlBXYehRKB8Syfzgrt2zgxJOX
24pxrTZLCrqn4EOza3v0tuOM0ZIfW0Dd9EOlpQAQEBsE8wL53o9scI4aF0TDvhN2
oTcVQkWdxGUmpYVmmX583TuBwdr/OBmJi8jM15CtPrSMPrcj/dSoQnGFsVbdDhh7
ArKycma9qfPh2l73IOwAv/FzpfsWcCCQJs/nXNkF40BcDd3xmwFgzdorH8vO2pKM
YIeZiWU2preu9rWyH4lBkdrYTJuc9TnirZulxbZOzd8aBQv7qQbtA8I4IiHbF0lf
ItdE08P4Wgxbw7r81reCEbB8+xesCyJVjjI3Wg2gx4z2PfNxVDZZFC271Tx9K2Ae
ljZMvMyFPC5KITShSWT93vLXHc1bVx6mhWXd5x5suz+PkrKKFgbUgxLLzjVYaP7o
32JuaIQojBUf6URUcPrCEP99mBIIaVYRfsDd1XSFsUQct08PVMFc/nhScdCpkq5U
srXRPFXVnfXDo1CSEd8EfyVEXSDLzt7pf0tTDJbbpDdbbIxF/Szs3OmO5X+vZlmB
tnhlnK86FGOzgywgntJtfkRkGtf6CNo2PWoADUXGdqibVwWH+aWyxoh5wdi0Fl/T
cEQcnePPsTMtvRgqwxt4CiyAQ6coKDtyL+zBXZX9nkmOjWK0fttRBVlkRIcMa4HO
TjqWsbUm4hTNg+eviHVdxkXKQ12fZTCjfyeG3WAUhogj1tGajw28r+99Ueg7hjAD
ZaCtiIdC6u7dvQALTL5fZHROJRtycuFAK45j9DX7kB9cLdqZ2/WMeW/fhFhlUz8n
o5MPFQ/FUWF2PQfi+fFmK1+iAUVPqZ+0J0LR7etYL8fVmSP20DW1czNSWbbHsQ/H
ru5+H713csHOtBZMw9BcHnDnqDYl9H1VZWYJtrLCHb0wZE3uOGw7LTaaVLoIseV8
YBgNUC9e5elW6JNYzSjZ61UGuLxfb6mHeS7EZ9oea6ecfYgT9vDlLf8o3SaS3NhL
FV5CiUP132jx+hAHQSbSXfOldMNtNRCw9IQjzdj3Gkw28Amp4utL9Rgmi5ddAoeh
vvw0sgjfo2J2vN7rs19Me3hYom2MUhHSrDDEGU7z6MnnoQID0Fxd/xHwpYTJBzLv
mRmfCU4yX78N7EJDPi1thO7h3UEW39zJ8th+yhnhC0mP2r4aqJywLRq+e1bqWCzD
LgkOWHLGBO3t2mZi4CSOrnSEFtt/ty8JkNiy3O/0fhHqKiIXnlLpL7ocZSHg7e2w
BelYCJoxkwztjRx8WQmp+1rasPVlY+cFzXWGyvK3NZvaTN3DTogito5WmI2+eGpK
FnmIkQh1uw7+JSxIqWJusfHM5vIx9mJLhU2AQ/8FSRU0HRv/wz0Asoy1Bh19Gogd
K3dyvBO4maOSS87PG5t3buf3R1yaPAludvJlQkDcnhsIXp+JaJ2Pc2r1J58iR01Z
2Gkax3ZYjcN4blLGzaG74ClJsC+r9it4vkVvZCmxlf8SuXcVjKDhXyNiwmkeZuLt
2V/qUN1bEd8GZGIWu5LZLf+CPqrY5v4u3H3qeYjFnwFErV5otxNwh7i1r0D8R47g
58hPqkq/ahSXffozCYQr4U7Qxd2KhrRulcaUp5/fpNns6Jo9aTbP1I7njT4lU7lg
82HfAyZAhBRalZlOWr9W/kQ9AzF7Fg7PFVhLC1z6kQNmUxg6A9AfmClE60dd9Dse
XQnmcPd9RmGMFrYtdguG2U0Og7Pa0KWFsQ7iquryIyBxe/uBxJRo7JTdJ2mZzp+t
A6mknjhyYt31cH7vVo3mbqcuWW5W6vw+ZZ1kPXZnV8ZbMSWGbfG1k42Na4wqOf4a
IjyNQaSUJ7JXTHscGHQM2VbwwTLJpVCoLuSyrL22lsdgsaAImEuNo1uqgVS3HCee
P4b6g0vKN8JIsw/CaMRC9fswNyjn6WWsolcRqiU7tk6+1CMiNC5cCWBq/41Y+0u/
UXGXEHZmx/Y5vecdcnwg77ewG0J6vaiO6yB/jmc4FYBd9q4YuK7L9WHbW8iIs/6p
SDgSKmYA9DuPKm4rE/kuLuHGs0l28uiwWPXlCDpfKoylRH3GNXySVFhFP8LtWfhY
6BdWvKsSbrZQoi+GTztRS9zEM4Sn9dgzWpYz4p61RuAuxypuy+qPq30EonsPlgHM
uZD5UoG+nI9nqwdLRVw2fHQEYgpDchJMjNZJmvZQItv3Ri1T51bK7+IE9+wU5nAe
wAKeDOW3FANfjwr4hjmFO9JxQGwFojyWKxkW3sZjD6SSEw17f9lU3GNGWkfpzXya
cxqgBbIzGI6dtkLvrtsxF/rcm+Wtjk38CLcuxEXnYRdg8e2fuHxleyWsa6luFldq
qCctNgf5FHSP+nQMjwUxtugNmpneo3qzTs0k2gPhRAv5kDIhIK8KmtbymWAujesp
EFu8/usJxgUCQ8JU6gh/bcD3gBt7b8vFNACqvUz5BDg3Haer8TpOtqOyHn0MYHcd
72oQaRQp36QZSow3B/ja8p7Tg9DzC4KhqZkSYQXi6++tPF4MUbrV62QrnSqROzEi
8ajLrkKPxtZC2BMsMDfhCmLm3FeVRuLME+8UgBBr4ufqq4LVP5TX1XYpTDZqnxPU
UNENS/xBckqdIzK10nB7jmqNENUdXYIgzLimqOCxPp/Rg/MBHOhO6ZVls6PXpKXJ
H8FmlbNoVCSqojlEaOMjZOpWx3J+YlfiI8s849kPJBKvdLTtRCjfBNbHzGsmcc55
wovdTvknHZeKCw8XtbV8iQGzK7b+wkEJcyxUC7fSQv1NBNnohS+E8EO1S318H7Zy
Dn7eB9CKAyeCjyjIflHoi7P3sRX++quPgXlitO4YEQcIQE1elmUHrV6hbA6E3oC7
/KyyUkMNIjcV/BgmEazI1uV851sGf/mg9LzDYbXTrg6fFhsrEWHRbXHOtI8OAbFM
n7omO15gJ9bAdFqgGYeLMsLbXqHZ8pWUkLf500BWDZReItdxvD4OpSM7GlxPyb9s
zFK5epInIkWwzOcUK6lAj/U4cYS6jSCLEYZ+ni4wTbq2yCMGMUhtTk3zzsIYvrF0
tnPw2y35Va/8gjTs8uu4I9XFETBAgWyTfYP11S9oqD/McN+17SfipplngH5Vh9kM
Lsiy9EGRg76Vqb1rcy7g8ZYdDuD70qqoCeW2KIsOC+D9fR7tyVyweHFNQfnc8Axa
FjoWs009FpC1S58+wS8xwekhq2y/u442PBiYibKThxLANZIVzIoRgpz9yA0M9W8N
zbrJObTJogogWo+pHMNSFQZTL0/zgnY06VjwKrbzeWWCmdXhGWs1aA5MnjQKdD0k
natbblwuBD5enYDCPxVIPWc1B48zIun3KV9yaCKnsSgzdY1nShIg8tb73BMab8P5
rl4jKpTrNvh77S1FLiM1EU93lMfiqWu3gq2IC5l3mPfPrpxCf2uAuF6RB0YPRsXL
rns5VkRDdaMvbZbjGUa76lfmNpsOYFiGkE1smviQJEHG3N2lFxMLsGQukJbGFgF4
auTmm0z3zl3jpgWIYtMYoZZmWhKVIYsLGeBkRmnZfMPnTXUwc5DBjmFTkuIcJytu
SrxJLvwx5qnb0USUwt0qtuc0w2Y0UIkEweU51zPC3t0qN9HxW3EKEOvINqL0yGcA
w+I/ULihi+guFNtr7GIVhil8heHHT6TfdeRlbcCMMeL7eYaRvcO5JZP2YaL118TS
/r+BAAHaGl1NBeYuLl5Cih6hCrzUGq9AuqkeBGZNjl685eR3FyWlF2W7Xw+SI6V7
tlK1H3WwPhRNT45b9pypTv8Vn9Cjig4Gj2faApernXuxDMydfQB8FXDBK61I1ZsM
7lQFqYmQtO+/49RkEqtagXlOnVLgf9q6OZU5S5rT89v1hdPh3or2g8PKReMWGn2N
TgVm+k7jkaFga8zRQS4T3Gxj9JJRmI5hoKQOB+ldCGx3gaJAWo1wB3WCdABHM49f
5VF17Zt1vdJygRH17b0AaxcmG/uZd5ZQAvc4xOSTUPeD+m+2AktkyvzJgbO6FwWE
MPwyFFS/HDWXZ3TAoevDUHGeh6BXNsA6fDrjZRB7WDrRY5AP/tHXWAp6pYK0laRU
TtKKb4FnWcmXmLj9DKx3CbOYm9Vj/+EPrZAsYext2Ut3GoZ58aoiVADJIoi1OW17
1Vy20hKheASjozcb4tR1ygkS7cVZp2juJQO+cQSmsut6qq9hPw+OwUDY9Wye96Ax
AYuFCJnG+sPbGwq1aHSnG93rcGl5eBI49rGgekLqSZMnQDdxTMnpF+go8CtAtd1O
ksinLDGqZOoIkghz/whWF7KWqCe31v+oeC66cnpqDw9UQbOferg4LWBZib0lu5OU
AhxnHDX0jNFXcSOVi2J8OesmhQCasFAsEBOV72LFfJ6R+9rUUCOAnrZO/zOVdMDu
BR9BrGgdvsoDwP7qwY3M+TC76MeP+ATy4MXbqulxYZUW5qWUklVV2KMZUfFvOxBp
hP2c1as8aVgybCwci0E88ABDMnz+3Rm0rsbpB8FfOnt7HOWOkGEatIngDh6gPFe8
MgMElBtandO7vtEj+g865IhJwdyFFHdMl5AXmId1fworgC8tJWYIrSHi9cEPcR65
CzDifDgMPprfqrYMxISQhLYbUtvPx/10kKQhlucp15j+5ZpOHJ2Dd1vu9uGYFJcv
nAmsJRpRAJ7SlD6ypCfjnYo11KcY3lELQMzy5JzPLPdbPdW/z55pRaiQ32WgfDWB
hZ5es62cDtPuq1mhyZCyRBJ58UsTK9XOzpgNflsoc8f9JVsN1DHreaRViL103y4e
2sMjjfdPLFA1cQ74MhimWE58h3o6dyUzILy+6h21b7xiL2b9ESYoiRqLLrEgcOcG
E9KHzHjv0GRBeeTwe5x/MkqXqDOX5R0MZ0c70koaF9kWpTG45AzfUjq8rFP7Ubhd
+nPw0PwxA33htkJJVCIo4aQ/n/t+3pe/h4MdM0FJFxy2aAufMh20xHfEdIA9/1Q9
ExpSMmkyAtR/20KpHnJ3mlHM1lXX1UZoH0GrlPthB96id2sXk07BTbFOVVIuj+oJ
oqDy2g3MrBYvh4kEB6JZ3T8YrZryj5AaFQj5PVp2hfhWl3ccnkLNiIE5tk60BDBK
hTGcY4B9ybVwpPDYV4mnNsIxLOAahzHetex5zgiA9cYbgLfs3lJ9RzSfULykSazm
C+a/NFNMB+QsIFB+HZjAV/viZIgwXTX5x3MARxyR//B74TRn99/9B/d6kHDnl2YQ
2+xW7IqWBJRPEVH8ed5kwaod5QDv7JTC85tBkxn7gXdSSoavj0EJtvF7MlivFgV+
g04FOdZ6hhbJ4m3LUJ0WZsPsZVLCwEXBgPHY5dXZZOEQLqEB+PDPvMjuubAArnv9
ECQEq+YLygFE+LxuIyLnh2Q8+VhsnA8xj7xKmIo+4bQlK2nqE31VQoLIEJDJx0tS
uZHJuSFrPIaA2O6ecYBI+j+Xf0nVCMcZy9yNyY2l0CPGR4/iGraoY0YXSYh5MTtk
3VDBXxfYMAM4d9c7l/KA0pzjBHJz/nWe2SDfD9OQoJI+aeScK2Smbc8sgXq0V9/p
YCtkC6zVzJmox5iSId8Y9ysQvyrgivRjoHUlqqeFqMEIEHtA4o6pP4dx2CzsaqN7
oQesVwdJcG42qGiCh8jQoIy6p/tC6Qd8Cv+N7hH3gHy9QJogtIKilBeesB3Xiz0m
Kpt1wfGKh43zBCl95XApX8ehPKxl3cA0CM1ZA3+4a9t7c2ptwt6M1w6irFQGzBNQ
fN4mEAR8W+BMy2AlK9fGYyUAdkt0hmTohRPUe/GS4Vb9gpj8jf04xPt6gyaby+aR
2ThqVyPlIRxsAanjXknrKuDHS2BrRFmzjsfeWswtdo7nrb9NeFSdUXskNGfhIvzJ
ApfMvti8jz37Flsz16CrzRdlWYHMmqZHuqTiVJJEZGjabqhpHLHUxcfM0WAUlOTA
YgfHGJv263+UI2RxI6QadMaxeV7XMWQkcBTBQeFLlGEc0tW2AGUNM13Gta4LVps3
+/FFuWlsqQ1q7diy4vau3TtiZy4Sq7cPUZ8xyrk9RCiHjixp/edtGds+sC58h6Bl
FkY1H9E+g6TaOqHtTsRjT8+xFCVQCmU4HbiiKhqLmM4RlI0Zyj6VQOm9WNJbCW+k
WuWNDpXd8qoYdh/MhlmNIyH+M9o1WxKXXU1/cehYXQn9iTgAHraYrw3yyJWwKOqM
UbUz6eyjUx8o5DFEW7sYECUXkLhqUbTHnPxjUqsU4Re5TLpsIl2XLiP+MXnv/4b5
ihlSIIxq20v8Jn+NOk/YzqFpOy6uMX7PzEAO3sz09MXIG/TiVs2y1jy+CBbrpbyX
Nf0rXlLdvjAQ73qB2ukDxbO7Ag0MS8Ted+xrZA9/PJVzS12xgI2qSXR3Z69Z89Gs
bAv6SMhD9QHkg7ZtkqbyPuRVjmSObrw8mBxOBla+HnxejWOyZiMR76IYAb4aZxtC
pjA8O6n+BaEyAMox2R+30AabNLpZkWUCsN/B3bmrrhO0AxdWT8okBlW6Z1YiSdt7
udvbIM6EeZmb8G0CmIDcMyrCXva1oM6ZST2G3dT+ycba5LDbCsGBwDFUoF5yUbjG
d0FnO6oJL+4+V/9+l3felD5KbcI4BNV6G+E/24jsqtclpgcmtpzVowlBtzU87tiZ
LkL+bOPxxm4IFgm2HWbKuWzcaWPEumdXXrUHJPAW1yPlOEoLfqiH+U84bHgSIsei
xspZkuN2entwH54ugGzsFYslMz7Pc+kg5mo76SHZiR0uq7NsFEnc8pDnCo+hypKS
ezsgzhZ3neYduzgR88eZPQlFoxkDzMbmZPP070uCXriazJeJ/Lim6/iIE+mfR3KO
BrYRTmiNp3Xb6TGkZb+qdjDVuX2PsOY0OjzuiHav430eOwlI8SBHvAZ2FtmXP7nQ
uKcC2sqgCh9Nt3gbn1fE0DGc5hL0dD6CUmmX84nCNo3pKVa2BOmegwDcPWeltMKC
iZgNB5pMSidj2cq1Cr5sUJFLOX3b+q8pQDO1sUIzjzphbbMTaELxlNnDggaTqfc1
K71WSAp8xBLIzWd572YT6A8QA9fWVLNFucx2B/vcRw4npNklFDVD4u1gTNLNb1BN
7U7KqYgUSEIMWu5NxLrFNWDH+7rKvULpX0H8qbRAox+w2YpEIe9mw8CXcA7Ine+/
ce2BUNyN9OaMAWiwcYA28ZWlAO1AfCttvvxAiRrVJkSiT4hlf5Ri57gtGPT/Lrkx
at4PHuc9pntTGklUcQo4E+xyKW230z66cFh7oAOWAmVzvWCrkOTUmT4ydP9GMxLo
u6HDl/gtwdX4EwjV33bGAAr2v0FeVc0/3TMNEsb6l7ZKUD8ZfAnO3OUpL6t54TC3
JO50bkGg9gmTVVrmLkd6Bn8Q1rdk4ImOHdDErJu02/bqzbpfQbTVDT/d8sizYrZC
0yfX4geIQIoZgwf3GxMMMlNxbr0InsQGHOLtvVXDW7FgkHTkO8Sw7MyDDlaSNPXX
50E3MH0K2+/T/SvRkIpscQKynJ0gVVnHgiZm3BPwGfTbcSz60iqu6N2vYsYurK9i
vXqpF9ghipcO4eiYhsSexedl5GwDybrxMfSCOtMA2Y1mhpZGPAnO1i3O9y6V06C8
hIqcUA3pVJMYvCQRBn1xqiw16pTxITWOgo1JzfTa6KuS5TnpiRee4JUNrt+wtIZs
OK1YRoh1B3CZsaP+C+ffh98Hu0zrW5f8UIs2GjK8Q/rdFM9sxkwU4ukUcQA6CRo8
NmoDldC+S9+wgdaMQTpzsQLsA+vhgxAQtimsAlTqqB1523M3Gag1uY+CPm/B8S+C
V59urykKn95fJoES4Mf+4pwG/vWRr3qknjpLlaldCELGrmv1coXXbhjcfW+Gegh3
7eXZ8TJEhDMCoTmeNnOPQQhmiYJfEaB/aS1xoAf2jE3g8JPov8dKO0X7UUSXYPME
61Wc/EJemRcYl1swraCInNJzigDdB7LNHJ95yhF/l43CNy6ut8tmxS7FHJS8vm1f
uW1woDbD86/V7NqMadtegy5vGGbZ1YKql47Z335Fr0bnGh/4PMLMVHhg8x1pRxap
xwMD1j3eZ5VW8lAw6floNtykvVHQA8Df/99m9i0/nRN3GtImPeu4aeKKm6zwSP4D
vI6ipIoxYx1g8iARZ5Do4Wg8Frtg7YJ1EEIQGFs6lUjz7cYaAaaGwyfyx0gbTI7W
RaVQX0OawAu4BT6110f6YUUIVdSvtvTvpujhAlxFpT5b+TvCdoRvKL+V4HKIPoN1
spSeIxyD0UInW2nPTmxCnLEjtaSjjtKY3WgMh8baIVp/NyhQLqtpeKkXZwpWD71g
HgnmWAShKPSsZweJVs0ztP1UMnP8oDbEFJGGTqR0so1GB1G/LOJNt2uNlmMjWpx8
mNxf2Ibi9Zts8TEN6wY20SkEF8Be5v0q1wgi6wbNL1nmMlxQE2b6dx0PJP4cezun
W+GgXxF9q4miZjFs5/u8/iGNP6jtzp5U1zyNdOwoEV2pU15HUVTQXrSCesVTlqgZ
zZgpQ/WmpfxdWeLU8NbRmHjJ/xo9yatTDNt/qng8mDWcyZXpuV6a/fBE906It69+
XHiG1+z+h4Vu9hEAVZ1kUCQOixx0DNaT/nGQghbWIwrsgtMKxjSNd9JU2YVSaOTJ
y/9/r+6v93432Ax5wAnpAy4lB+97tP1aM5P6PeNRdPAhgQVKYQ39r3ZrNocmu1y2
aygj5punrwi7YmWdxCHNrsjJi6tOhw8WnYpQaX3wQvFOSLg88rfMawTrxdOVQV62
7l/88KZGJ0vB7rGKseS3V6fHnnJMlE3mxDB8uQoWgSsleUYPFUndu0ot1P/zE5Pk
uneEP/Zxigz9ahyUPD9UKeWilYTZfjzaRq4F4pfXQ3hdIGXwLfcAEWPR4iIdUUzm
ASg2Ts3a+2FeO1DQ+lDiStVTAuCzJhtzO79QWum8P/ztH5Y0/x99OvR0jJJpsYgQ
n3dIql18f+Yifn/wmMShgZCJ9i37UmejAunAxsCACPaBYOJY5sexVbMoAi9VDGH7
Cx1SjK0igsFoi7HuDGd3Nau5tMN2BppkdHp4vV6a1Pi/KO+Lm8GoR2Hs+9+el1Cf
kMweXU0NOklw+i11oYUk+Ex/p6fGIYGKAmgB0Cj9xcCRfBtIwLAA9/zfEBKg3JL3
po2vQoTBdz4OfgZePgGfIkaJlHwCNGXsBg7/cMSopzP+dEYzX/X5o0dLhXmD5oGW
tjWHHnCHXdV4oqpIYxyzDLxYGL/RodVyuzZWixHclimbJ2h6FMYu3ofEGxWmvF3p
r6uafiu3QFWP6ln2nZKpUGYPva8cyRCNzlSEIU/r4JML6oXg2nWY7duImodI3EK6
DqXb1ekYxAg8tXKtU3JM3/qvu/H+3rfzp+OJD/qH9LbCM+1lOshKNLbyDiiemhNb
1cRNLgk6TSmfh2ia8GPGs6VAF0wd+njwD3h9KRcrfaHkV/dphdkAeytWOjgKAKFt
AzQvzKyUayyNH2xjS6icj8HGMeph5vausXEhXrchvLH3uiOenb+W9xiWPNlNIFOx
T3ZwGs+bW85Lz6qDBbP0zywJkhimuWievUk9O/KcXqadwZ/nGBQdxUzNd2AkgtuD
C6WTq+kHSEcb5AhGu8EGV5hTmGlLOqitRvGGC2noHeedj2lr+RTnqJd+DXC8HPCT
jjRvY7CYfV1SL53lh1NcoS3cCsqyl8NvshcnD4JanzIO/E84wxoPx/0o/4IsC/Dv
bMGHslZ0gxeUOehx9qXXdk/2b5aK2k1vdU7gvBq30xmP+PheEIag+7JLtqCngSkr
CaQ/RrTBsfEkRUO7j65foqO1hcntKuAE5OErK2vo4FNKlOLFDz41O8YbTwacH9IT
cC9272uVOnbS5K7DHwq3uFsKFjGmFyULEaziotBCSZ7PdysloWk1NAIuivVU2pQQ
9LI8yjSA2CduBnXUT0ztniRjiDytuj9ZXe2Stm924ypIi2TaAca/7rfvppreH0yO
XtmInYHXLSXgkglPnWUUu9TZ3yszXjkcML+NJxXtEmCM2KjYobIW5nSMnlupcvLq
3avLtH0tB6fI/E+eBRPAG4FbbjNITQ+8Y45gGjGAV/rQfTLXYDIbOXLFUL8Y8DL/
2zR1+gIJ1FUh5GxXYm6GZz3xwxeyb7UidBMqqsS24zJREsUNq7q+bRdPLllNL6nX
K6qP43UxdTX/rNP2krDeYGUR7w2jfrBRVjPwZ2K0IjBLuDoqjASDxd71KbvgJ7en
xTT9u+aCwiXK0UQ2i+urN4Amj2kb6pKIeVp+TY6rBsTDmgwSx+MVdG88nj0O4naY
wX/uUXt6uQ76h5Q20LVh3uZ4iQin19PK9R4ryrNOpg6BGBH3wmELSQ4ySXu3v/gm
6+3evMXg+J/y1vBllwRYKWStA4/cVOabSEEoNo+veAdpZFhUW7QHLAoyEpWS15z9
E0ICaqEPZhobnQOnTa3iAXsxicqvEVA7jvV59GNy935yLb9blsNXg4fqDi5W0dWt
b6AgTZ3mhCw6z1GlIfZAeMXFFSOsQV6Zg2UUeuP9hXfeeK1Ub4KDR5R/VyK9HYW2
wmSXP5pjjun9zKO/2EBF3k/Zwwn9Dz31+loVaPfa3wypOLtzd8h/BRwK41sHqjtR
Xhuk8107Px9K0fuQKBlZ2lRfaDzKjAmErq11+5qC7NGZzxIG9XkPgL0DrG2ptlEN
Wyrn+lGDfLyBQniSBit3NVjoeeTHx6Q2quOuf9gIlKGP2Bq1pgybqfCrnPnr5sjc
tp4XSML3lhfsuDF+7GUppgb58ns9bchRJ1G6TCd+7Mc4kMShaYaId5ZLslTxiixe
qY0sAG4Mtv/4yLrZxlg+IY71uzdCdMLUF7iByX/h8Cj5QYPDHXsPmDM1JMSXmRt/
Y/vV3uUcN0UK+3ItF5u0xzxEQaUJtJVGycM6XnjyizMQcXg1Ennk81GjasY/SaAF
fEXQZ5mgfVN5BMjPQ/WzFg03BMWTfu0t0x1QeHot30oUqYO+JWNibnkotSdb75tw
x5m55ly/yhiNAW75X2eY8bIEZsNAxLpHV7lxddCcwrSBygfbWU2SFA23a9K/4pLv
JiamLNRCmpciqANg0lmnA1/mmnLnGtFx2OasxxuJ/JIjErbcU8HaneyrKp6lFN56
aVHUvLKFSqJLxWKdCp6Ao3j5Kyer8hulxSMo22+Ibg+MUfMHzHJLwjvJegX4QbOE
akdcAhS4GRIiBaSgnrBOb/4EuyRMa4ycVU1dKDjsJyf9IypV2to7wwPiZgmQ6TnV
+dJQSifW7/N57+PVG/3H1hDgY4lp++el325iHO/oQ3pl7VogjKcBdU7eSHGhHL6g
qw3QkIDQJMUqNT02+yulz+x0m/mlN1K3tZVsurFBkCYwPXIbkfKXAP06cgecyt0+
5XuNjYmmsoCc81+Euza22m++I+o4uXN5lcMYhnYyY+WK8/Vivn5sLsJjPSh/ICOg
YGw5KHmJ6cfTG7uQkn+QN2OU9i2ogkXd7HacODZsEMZKnXZUjK+15OqJVt48x/bL
SNB+i/6R/oOTNOVb1iwBKIHHakklxtjYnd5SqRi3ocZHZ6lBy3Y4khuJO5bexYU8
hSLxq/KMO8PSpcOQBju2rmCkdwTwxhiXm2rSArlhQInwJrhRSGn7uqmXkWzoDKBj
C1rexl7nRAprCOEmBYZ0c5kYTkmdkNTXSsZrY13yI/9OcN33v2SzlOon7b5YeM2k
327jiSHFxS90zdp+rGACQ0pONm4+sw5D12p/wTSZzFUgSrSQsctlVkL5rPBpHJQ0
0YchX6oRx3VlwnDjjUOtGd1Pe8KUsbrM6opbetWocPEZBkUW4On1iuL+IYlM5Xbe
vH0daVTgfvVa7ew7R67QVi94ozef3BqK6DfBDKegjps5YBu/rxGsJlIOKO/MN8Uq
vRp2RnqO/BYREq+PgBEMFCKKWsChd0bDAqceAJnJOm9VC2Qq6z5M2LIHRvNUzYJ1
+3I1jPPMr+Tv5omXStq+tzIkdMYx7hl6evyWoi1d5hMpaNcJvzlTBUILtEK2MyKj
f7agIA8zch9r2i+SJ0jb83OuVdG0334csV0l71NoqVSKdVi+gGTGAEHgAaWPPCuA
kWKqyKytJCg3ZEyocN+9tUJI94opQlmfyCG1sEcmTVNozVBCG92MtGObO5v9vJgf
jQUQqsmbL05DcTsWd0+/GBvXPR71LwnT4okL1Z9ir7i4H5jdQMgTLu0xh3zyqpmt
gL/CxS1Xx9n20xAoGdnlq5LZ01ebi1MKLipzaxckXeeWOCzBJKkmmkd/ZoNQx7xe
Bdgmmo8n2OkTFc0sDcA2AkWXlHznzE7VX0hQUBwVRXiFC0GnxM41tV58uJgZPiOl
R+oqgzOCynuby4BzhdLkAvh6kfT1tNoT9W+PnluRKM7ZhFtKt+I9xSCalEhjduJl
ACfjWx+jQ7BWWbxROjzbJnA3rKMUknayVj51JHmEmXJ7mJIhexS0IjNBDwuxDn3z
0bHGK33wS10yZFIDE13iz1fEbCzJBUO2/0FJMgYrR2na8ArpPMV9Ow7ffJzUyROm
sD9j5UsNKFc8XOCi7yTkU+oR8ft58i+Ps21F4T0kEe6X9lpVoLuMyMYk+9KHF6Zr
wjX0IItrfXl685EdsLDCwUyv6BrFjeUN6QUNf6V/XhUSdO/7yM/5jcd+xnU2DMKu
e+9i+jn2rV71sS12PQHyppWrt/kZ+o8WPjz5pURUliLvxukBRNFQa6DIQVKWRwCn
REcRam4MGtczV4nBTtCsdjgBXqNkBhDMXARp3F9Y07UcoJAGCvoikqGyHLDJk5Bc
tWXpcpDqHMgI7mt48eSZFmop7U/ZDTMXgZnjQ59/so6MDlmdXhKh4k+51Ov8t37L
zgvEurE2JoYZeGn1dOyvDVHk2IX7NQCAYyE5/MkFbsT+SzZGzV5zdpPrcRIRcBxw
OC0RLLGk1LRZ9oX2R7teN0nr6LJdFp4fOod7xn3U/OzAfZcWVsNipc0nraj8+1Qh
upc2s9/xW91yOW+NMNhfVmnLsoltunL+2uX+3r8jDV9Sdwsf3V702fd33mg8wice
gWvFfZHLYvMY48eokDyn8E7kzRGh4QI9C7O/wCl55/FkzhKTfgueeniMH0oG2UDb
3071/GmUrENRFhShuhjtV1KNr1qLZ2zntsO3M+aUdLvR6cGMkm/gfnP6hj5cwU4a
1c8wf9B1KnnP42roPtBIlmHT449ZF0jRMnEvyRPDsNQIIgFWT7Oql8BP/Em3GyX3
8cVVsD/dd57SU2/UzjqZUKQ3lXjMtL1xbhaYm+C9kxIhFaEb83lOTvTyJ4uqVjrK
PrRztV0UJqkbgRLmOrhDSF/zq4Qjji0qvZh6HbZrPwi3n+/DQY5CfzamN2TkkLrl
72Zu+GBv8NsG+6lK89HX/qRRyjDgKixGFk9DUIA3Kh1eyDWUsAIW5AnvilknMTpz
0gdwP9I1E12+fUCxJya1NqwtyncWGiZOmi1jtsZHTTGEoIEBcAt56W6gT8isXZl8
xoMQmAJUj/Wfq28Qnpsvys17z6nC7WWc7U9/XiB32/88c7N/3rCQZiTZWjGs6qc+
JtgYwUroS7DC/BSXReMiYNIz6tkbdIHaJMAWPwHa0zK48W0GnzM9Us0itzuIu0Fa
d1X3f2sD3BXB1HWVuxg+JEHo6YHHOhGaJq9gnxN2BvqmNJq8s6AijnCqqW/X4oqJ
yj5JUjgOQOLx1Fx++4f4T8X01Ssyo+J9Vuzfg2lKoViQZfeAhxAyn1qM+SqrHYla
d4U7MfMNQYhFnbuBs2LCci7iTXN5Y7Y1GrQ4KlqRt4znsJ8uxNs6LCMipqDwkWlj
OJtnxStC2luhDk+4Da3MAtgwY07CIxXBv9Fh6EeZxQ56HlNxaY/WLclxdPf7ctuK
KXo7HmqXH7pRpeAjxF69KxWjoBu3O1fxP+ZYbFBg5e3JCeX5ppF+5m9i6oEQrHMb
IO/8gSDPlDKokWW/irCi9lsKIKqMX89UajBLbZ442PIhSzRhhA3MPYTWa93mxQMe
1T6uqjVUIAYL3tZgF7PCcQ7hlwZrO1W6SiN98xB5p/5kkQgrx4KFCT9BNvgGU6cU
9mXHDTA1hA2bOC9wUu0YthE+q4hunSfybbD6Y3HWmJhaxI42Mjv1T9ui0tzbHdje
mT0utPCmXntghH/V5I4p93UXECd58TgA81Jh+MRkvXLJSkULt9TdI1es7aG2Tph1
x0HjuRF8wOLQK+Oy7vj2bKarpl7aLz1XIeGzwNXpuTo2E/v6KGbRZNXVubs+w3Bd
mdaZqM8royBpQcxHK+j1DwsUboJXQRCxyvu6PCPjHrAtpIg7CST5NM8q3UMNEa8C
T0oFkTOtwMUtW6lBHyrXiWkTuuil/sJOFU+WBuQ3FlpwWkcSSrTwuDl7rBYRm4hr
GhAEd+9Sl/an3NzU+VuctZKmXmUJ2bfp93ZdENx/dOB+INTsnrHS0OSzX57Li3Sz
6CbjlCnvA08fGoYIsw4e/MPlLuWy05Fik0QB2NIF7k/6zarJ4EW5y/AbA4JxgrxP
HuzSF1fKPWIn7VKj+ieMMt3n+RnI2KrK3AE1y4WIypwEcTmc3HeJ4aJu37Oa5uKE
n0nBUJKx4k6fkC8IYNtvAMs5CPTAED16z5yEX9dazNPuzLbl7Wwmp1bSGRgNGA99
A4DKAxVxv1lG6XludnApSZ+vGbUxQeABdLaIhmw2azgoRRf9Lv5RbNa4PRaFfG2Q
/VvY5bdW68y7Cfb3C8OPrnVfaI2/sdfhxeqygVPKpNBmFumlx4nE1dbKV6edvFXT
76na6sgnE3hBIpkAsYQaU3ixxXk6ZJuIZxUhdHj3OJsEpbozq9ny5pNdpZu953Zw
n13DH+7CyaH/+QDIGuWShuHPohsZJpdPkfLjxMYLD5fOrH8H0GjT8i3ZmDY/ZqUM
NrOHRxvtXP2XU/Q2pd3p2VPXBsxCrYa4tg8y7beQirwtIC0uWmq5zKRf3uvwIUaX
6ezyig98h4gvOCqkX98Q3qbfAyT3v34wrmqgOKbbSUI1LNiOAuO4K/e852abHY37
x+AdJgPCegvsdVu3Hlorij2aaVKBBOzid140XhiCY3Mr3u3pvevlErbGxaqKDmw6
gMzwW8mWoZ03FF1GkwgUj06Wxb5BH6wqvrXl1zz7hDtdefNpvDUUmYNAXYkvtfHw
mdUJYvnWiuKsPumXuHEEKthylXaAFbwpBvxW5YqICjRTxwEi17Ml0gXv2ASRNw3o
qI1vQP1iNSHzYVdfPzTQFe/b86mJLswv2NV38E8jcyiLtjn647YNYLwT3OkYKALg
yuMTKLFCad672CUQk78UMD1EYdnWkRRGqTCzuy1hd0ZGA/hT4w8mdvQ5WHZvFMep
TE/UXRDYgti6XlcCpQkN6xM7d8X5jrN7pRp8k6YLx2SMD0Mcu7GYEVZuZGJwXIvH
DR+Kzlq7TxJjE1/lvamyxAiCdLsQnaJuyOrzkfPSj3ZU4IKh/q5eNVnLQ7hCZAEW
7cvPhilEOoPpRV7+sgLcfRqhTjaSGXn4DTIgR0txe4IZ194ZBsJjVLlft9iyooMW
mvUS31FDe9zzcbZe6cxnCSJHS/tFmfInxliwdxBYGGeFdllBrAXJF0uU6FNrUfdW
aX3McVdag415uQcvF1/pZXQwVw+i81N5pOAOevWRtqMb7K5wTJ8C6bW71rT+cFJF
/iecAGwoB8DZdzBVUHH2K+9JfEYIGBaeKjoxqDkXcqtCas78lm78bOmzipuUz5cP
ohLkhs+xEZvY8dQORPxnhM94Scc5bb+n0koAt+CSOLanSJt4G6ScTrlW4huKqcvR
cpv0sNjJKvuTrHZqM2Mk99YeDse7HZoDC4ve2k13bADkFl4cKIn6Q68e2hGFiurq
H27FYCa3gfwqv+b9i9UBI0+ZJRKe15n9N+PBGU6xSf8B+A8G2abkckUfpSctlkN9
rBGcFGjADMIXdJuOFO3xaR5VKRsvdjpuWscJK4H1ZmkPp3XSu94sSCDGfTkIx/tJ
clqTuc3xCgLYlX7E17L6RRE8naCdukUg5+epsHdejRrsENqDnrS9hxIm4HVuSmOi
pz8is9ft/tLOVWD7JfVzDj97BrQB0MCShvi3wd8uY7bgYAM/25Hcqwe/Vj4FYGHJ
1J0WXHEaQdOqWto9os7lZTQXRCih2K6edts5exNJcu3xQ6ExIkkfNMRus4maK9LS
yxlewUsNDb3IYveM77cffMNpA/FO4JBadq4KUjQgPjbHpqCUkzQ1+VGm6PLpDObt
X5ZOVjxXBRVLnRuhddHmOAfxTHfFJl63zMfEmfDmEfaMDaDH0c5dJpYYg2ip/Wd6
eq65SI6Bbdjaru3LvaXuRGbpQoSw2Hbjdv74TsK5D6Kfkd52jKkntHYIeHfPLgOq
YtPSrw2OYHz1/CRkB2rI1SicRF3ekjhGuWku3nkzgCZuivfx+pXkBHfHeekBhKaW
xRlLlV2zZtnq9ElkUOL+pZHclLYDR/GZvcp67UigX/+u6L/Ozbtmo7XI7FrgJ+cS
eUWtzI1qTBglyc9fzH9yl2qFpE5O8S3tadTWopEwVnUj3i9TfOp9zAYs8oZaqZIy
G9Grkcd5R4bbZ5R0HdNlS70Ht8fA4xhUmRbo6DTR1/C/mzvoFTEt2gF9M53Xpqbr
rpjujzQkUtVIZ5PRVdShnVhQShYsi+EzGFf0XOqrcRGl1hvEmfQTdGYv6WsTKIEp
z8j6w6dtz+Yex9rUWnS8aX5xfiExEl2aL/MJMa6j2P7V++VQYFa8kQFqPae7xdxz
p9a/4nd5SxOdZJS9WnKkCw5ReZrINoPM738OLNGnC17d1isFCkuZ0ht5d5b377Oi
KONDR2oWyCLwZjSdqrRjbK245jtVT7I4pCxWYdRYM5NM9IzAnI6B6+PO7rQ25vy0
vL2kl9IBXItp13OU/Q/C53O1A9nAE9KrO2yoBNxvmKcIDcqdIoXczW+h0FWnrCpY
nVmbV7VFM5y4xsL4QKwzWhpPkHV/JVQwW1XSMhS/Asohewk6S4u5jJe6MORrXTkM
vGfDyqc9f2eP3+XGdMXN+hqPa+kxahh5x7oDNOd8Fz0IpsyUn8flMnV1xzoTScxj
usbSWB/qZeoXeIOner5Rq2iwCTQtDaix2x6zW2YSQdk7GlsA+TVRzNeNuq0sDkSy
DBbOSfj3b5ysTZEaiBp6Ns2UzKEGNN6SvzYu+Ac6Pf8C22480zypPJWlOIw3Q8i+
GtShJTnzEPK/cXRk4OxrPi/jI0CUXlngAxUKakrorTWaxlRnNdV4Yp92qpyueoVh
PEGz5boT4T41Ck97qmmCIa6LMFEgvgGIjMVAsj/zRo+DxmweAtFvXGSL5O0QT/qY
W7/jdNtZrBDqUaiCo6ECJvMsaZpWGy0FIZaz/pvyxx6AuAiCKJ+OdYmZVDhzBLgD
VfGH9MO/nSkdVykWHx3P1ZNNBdVTL+RUUupSMplQw0jeTPBVwt/4PUrUg87S+43d
cdrCxADzw9XFDKwoksNdM8Ajg8su/S1jC48EwRttbO3fni5N6ajG2AzMVi4xtTnP
LlR7xptYIf8dmSsGoxEWxVrowsED9lRiKhdVb7ZkAFssct6rRySnCXIeMkYL8rvd
ENVZAmpCPG/yoAe/Auek59d0SbgH2Y14QGNYVLb5WFJxHk8DRic1LOmE/t0MMCQG
po16pMV9u6eR21Jz6eTTKTOa7f9hTB6OpG9pbfl0zStvSiGbUidBbzS0GXthwCDP
vje1FkYzaNhwzA84VkE8mmcdmoq9FC9G5UG5e9Sv7EF134bS8PAXsFoqHqU4rtKN
WnJvX9q/BCPbHXJzrX6fv3WKr14z+R03e4hmPxyml9aVq7GXrb6y/hBZPp69mjxj
Bho9PgzUSBaOvYlw0yDKc6tpBRJYKHpdupmD6GtoY6VeW8rYld4sXoWvy4trmSet
H/4BJJi7pRTuSQcd/xSwIgrA2RpvJqpe3L/FmaJ7PP6+awPioFh5O0RosHhqU51C
RcM7h2iI1OFqtF/hhpQ/Rs/KNLVgKN5UEYfxcNojQHK+a6yoBO2MWUXlN+lsQS0h
2BRou1PaWjOZkcx48OF4Bs3y9Iaokvckc3ULVlFhgy/VT8BOjmaWI1FmvRYg9GSV
7T+hm4TbL3O31hFahT7yUjhqWMQEqheNa2fwOtkFWA1i8oVUoujtq5rlMekaoKTj
ExpB1g1cTo2I3VoSRu+MELPICyl1E+QwqI/c2iNTTtmvWZSLk7wMYicMhrDNxFmj
cy2C4tGXeRBdd+AWjLtblYnemojxL4ub1tWdGeK0qUSZ77QLNPMgEOoHCK0MZqax
U8EVG3krol0YYw2lhlWn4TgXJmidgeWhF8tzFWhC4ysdKPmzsR7tO/o+lpg4OATd
eAysXOZWI4v2YC4pfS/dDGBUrbNi+0W/h7+9z0HXdhhh0fL67Rt00pzWGrOv6RGf
amE4UrN+8AVQen4y2JrPGiE2GtlurinL/QNJPlnPHWI/w3OfK+n6TsyaN7oaqyCP
zMudTRmN9hIWtz93uhq9uvWjbGDu1x7nfAaPUZIl4kBtycmCzG2erRcmcHz4mDiM
QFNGTWo2hdylhurPBh9Xtk3qTcL2XFYNEZF+kSMlhV6baBE1Wne3zmdJMewtgDmq
YOv1b8ta6RQbZQgX73Y376HS9hyvu6g6AZDIXtwh5gk9ETI5gbU7e3H6qSnsVh61
lk1r+spzEhWtn3ZPc7RH9FJiao954v3MyQCd5Dls1hndK15PffBW2yCYHQC6GLVB
fShE3dVe+R+JYIVqgJBrRgN0wLbYwGdmHemwqrqSH6cL78mV4gunF91lJ6OM0Twx
UST9ANSm8Ikj32LC17kp23IpZqar8LPQZP4DOUsNHbtCXYycOAWB3gMpY3gfx5mE
jmDqm1FKSF5L4+cArZKP+jYycO1ILfKIe6ux+ZS+v7t11HLA5Gf0Wlbede1HJWVV
KbRNIHUrB20qrO56RezNklZXo0c/XHBnyFyHU+2sWkwHH6Vzaj1ITJJqkUF//qOa
BzOgTG0gBr2I5aFE5y+ujYcDo+8W2rwFemX+sRWWVtnq8plnFqCIilQOkyqXVGaY
Lyngcxr7OwNRoTYq/r/Q38HKdCWi4FRXnEVO4FUjwIstwHAKXZ5PRsJvCccXXpF6
wEv+IeU3blGWJRNAkUfCKtcIhSlUKqf/beHrhjYXBl9iz4yaYv0L4Vyf5fks0Z6f
UwV7Pu7qhBdUYG+dIRUiEAYQTokqFgUsnDPdHAyPrPVxxpihxKSB29Kms3huNqYW
vVWl3HaJu7QdXcGJh/FKGG8KNl1uPTdKZ2cE4BH4HwH314uSZ2ENtOFN4HpM5rI0
lMtNwYyyHfouDvPFbXVoQnRTt1dppckFjBIlYNu2gjldWwT2Sl5xHh6pfTgsJzPU
Ns1BFmI8ljEdx7UVh/SDJyka3P9X8Oi/YbUcZdUqEusshKNO0/D4JzMucK1Uc2Vl
YnMgiLcPOLws3ep2s7z24nDIgpzqhbWky0HtNKVYa1DUOcr9/kfI+MusWIH2IS/5
idhvQf1d3eAbhZv5TUGS4i/PlYvXcK37zr3omI6uKk9qVn5w+AvHH931ROnyrGzt
PFBDeFknoVAHnaKRrByYJsKruX3WOuVfvVuGbrYr2B9rOSht76vEqpmNxel9jL1i
4U3ljapJOESU2SQJdLYg3Kie0N3KANc+MpXlXEZUOvFklz6Q1Krj6j1cB7Znmqhn
tv63lDmdoXQwt5abM5WgLeXCxX9aFsvu6ho3MXkKXxPI+2MO8ZyVyBtyp0vW5C22
CwzxjW5sSLOgPfAaxZysx6RUX+551zc9ZQLQA3qr/tm63rNL3pkgdKdjW155gBzw
o2aWU6va6mqS6yUB2/EjFMTyYvam7MEKJIWfYKIjj66avrA5MM27z8YopT8v8hms
nRv0DSvMBaJS3GGELlzNv5ZUzqnFRoZTKM9fSK4F3LV2gbej9MKGv9nUIsK7+6BD
CShk72QgodwspGj4V9U7fukGhzyPTer+2LfEuIQf873kTTeJ7/JCoYpknGBxHJNK
xngvvho/63u5+PAMkoWYy9/KKAqetmfOn74poo74EltphWPOGPuZWcrjHoqE07HB
uvQJealKDKFuK+AI6yQFVLbqBwh9L/FPc9ICMqT7p8F7mmAQz4Su/wVVNvPQBAMO
qtJeQUFvwo+2JeXjjnei2aX9NYAf0ZIkuzagvbFHClzNrtNeNKNSvkfuMnVrq1uS
VRZq5VakjYPoPSWtjmSH+zkmGwFbcbsN4yCHjax2UMAZTZsyqiplTBBn4qkvaSkB
+fwMuEZHKdVgnKC1G/FphtLTcZO5wx23cQ3DQdvFZ7iTMAh3ZgnA/glAWcZXgaRG
C8OSgkaC4e7SvhaLRXYEmvNmcaQ2Nc0sAmhL6kfNvSJOzcOPdrMix7vAgJJGOekL
AfEZY+a6wfqWW0uBtfnKE3d8xyZsw3elyx8hJ8F2Gqy0toIUrTl0BEcPcHyyUHcR
xKT/USDx8/Dr6WjKe6VZREl7gGw0YiT9apukwgwvcHOUXl7hE0WWTNp2801AHJOP
unpMGb8myPWsWsbshKfs2XLRcXt8ba88MDJ/q4fCL0fo9XVlz8GEni3Za8ZuuWzW
gEMQd3PxnyXLITJYuVmxSoZD32HoPFIF3dlpHZLIqUFJRpYANLLOfDkQEXccIduk
/uYlzzzWN7Ff1NdVwuhP2M/2nWPznwQ0rWfOHIeU1u0Q7h/8m1JjVoa8KaJ9oEHK
w9v8sgVJIKqvySSDRGkdoRzh4QB1qgPsFJ6sLtwjab70ntrincABCelm2+plb1lO
7TjeNOgGUCenY5WmVE60Pixr0bzaK4LAtwoL5ySkU3z0/K8xePG0AKuC9Ch3RmZz
nf1dnMAQ2CzhRSenwKZaakbYlIqlYwkAUcK0BI6mQ4Tgu3fdBD9XIRt2hazHQD6i
y6mOs8hHlZN62OuTQ7zkHucu/191HcFdb1kmm1ilRVUNc9IcbnMnLdrS3GJ7X2mM
8+J8G+PlwsGMewZKj1K/kKTcg1HQTB/0RG+I7ImSK+jCY13iC1CfYssSQUTMOJnb
062w/jDsd3Y/knMDPvfwqGeP85f0ZMyo5G60O5+5jSm889Z0sDiy25osnhHlvP28
Z+Ydd1JLBSiDJ2emGCIb3UINKQ28ky4SDU4rtoCn00/pxV+0f8rqknjjmZf1SFYD
rs57E0pTEZSwuxFgQSL6XiS8rvoi6Joqc12Wgd9g3rXXh5XuGuyjRUQUuqyl/Q7O
+KQv7XFfiKcCdLHVhCz/HyBO9DU/SAMdQB+jKAhgOKNhwj6eFGFzNpJdYBrrITL4
qAic7qcdEdLFqHBcT9tqiNQybdDybzMUBGumpUji6RuOngWPr1jaoK+Eu7korlgy
y38Y7W1Buq2qp6VLcmtizaYF8fI7fj3NSqtu5KXkvwIi0utku0w1tpicFnG8LVuC
Nd8uaO21x2r19A9nv+3jMW1/qSOh/qgPCvv516SQkUz/m1YaiXRVk7aa0DA1QrVV
+0+yrRIvA+5zX7X7iyEBRLHRbXtvQ3XtYrbnuW2VXMkDKCZ1L8La/sJEfWPhwCM2
HyhO9rRK0AQe83DtZjd1otZfLMulZjaKSbcaPk5w3RT9bLY2hVFngeYh2JEJXUtX
IS3EYPMSk762xU1mmQDZia9TQEuPX3QdV0kypPNa8DgHArnBxcFPyIF9TgFp2OwH
LZh2AouSgN62+ca29Yi+7AknXml5iRLVvXeu1gCT2e2C2SI8Cv4Z11dmxzQIvDjr
5/uNEHCAVj+InQ9kr2z18ZMVmqzh8tiXvsa4GX8qjoAwlPcVI71HiEnS1IaJ0NK/
H2cQU3GaMT3qaqALHnCr8oVj7xXS9Pa31y9yNZpH9sQzbhbzz4GURiSft9pcbo6t
jGzg4HlxinUXYi5kL6uCvSvIIYbqju9MoqcgoW6mL14h239DQm1rtHyy2wEv4bTB
fd7JroVBBQA6weobxC8S0BymkPKyNgdJHVd9xgPm7H6C5veXxr4RrsearUrRJiEd
GUD0rw3Cs6GtEbtMT86fVIrnyrpILaQdVA4XeAlV/zoJaZpeU89PWmV84NWrFZIu
+wH4m4vMU1QrVTaUT242l4VqU5PeO5HL6P58jWOJ+uXhUACTXUQqWvNmWSTEdC0x
wfAneESeOEz9ojPD4eRjA+BIuGfxd+D/lOQJZclnovdci/R62l/acSB8vQnr1kyz
eT4PeF8/NcVRHqT8lsbXQBAfqJ5oZ5SlNmdEKCFNuoI2rrsqiG8MCtnKujrtIHpj
YUdHUXgh2KU+z7eZsN5bXTJVfJaY5wXsbhrPRq3M9eXcKV9/Op8umgIahQIFvBYm
g1VtT9MPni1wzRnjNvhzUQHdeBGrXLqsbHm5Mcb6IZy0+aiP+lLCWNEEdb+5WmcP
/1I8O8VA1VW7PHxlNzf/EKpYUPCeSZJuYaMSeLBsWgM3CBkfaX9cN/xqZFD9GB4u
YPu7u+xgzC7q3wLhjfSX1Pqt1wojbExw0ZktF8MWuH3smDIpR130kSA787sYNyAh
H1dkbJr/+BDSw4GZ/qWRwsC5CkA6pZTFL7ubNrom7GmUJ0reoH62AcLNpdcnCrZU
YUNmI8m9HQ6xYVuf57Gpt++MfbPJOi0MzIPC2t8eMUtvUXJUHWJnOwYGj2UyAGIU
JaWuD3fpmmF4r7SvH+9bghFnGU+ELXU1IOErx+gZJEWUGujgLhJL1cjlBClvsa3s
FZFnSTbhAxtzfLi5m1V9aH6uvEnaD57g8G+GU14FXi+BU2nQDewnHWpWTXU52gHp
jEwnpMUQm3PTnLV30wU9jOFq+DOSkDgH6tQ/BV5/Otk4N4J9Ja+1bgSnDcTJ4mQG
VJZbEtJZ/DQiSudAlmqbzW83WbHx+Yc8cKRelWhRp5VRdtmpaNRLLvSuj/b/P3nX
FQD33lA1+5adYWnEp57olUJKAhxb+/RViWPKK25abiyeikfxiuUEcXm1imJ1DFzn
cw6E3+4T5VDO3CjO6nW1Kz+PBIKi7hyS5HiM21y9Vck3nSMcyLXN7T3+Si2DPMwV
LW9sRen6djgdCrc9A2YfdxBmWGkbKQybS6OUAJWo9gjmOdjXh4spVn2UIrpNVnAf
2XXBFKbfxRPIMWGvjnulT+lFKbGCGA2oAkWgUD0gamcdhbz4eyW7YkO+IZcj6HhP
PREhf4LnE04F8h+7bp0s9aFrtkaMKdBsvTLTa1+0oqWNp4MlltRKvm8Ii5wQm6a2
lkWInUHhprJyqvO6xeDgNVC9m3l56GKrdSMpnGLbZm6besDPYwHYxESWXbpnG6KV
VRzEmWz5Qws3Ho9u7OV2qHHXR40ky9KVbBQrnZYbnSElk9kfDmt8mTzCcPDdEX8B
x2hUf85E3yvieN1yZd83kJuQmuOEImRj0eJkIJDw7JdIlk1rpPg1TNtWYEEEY4I9
EMzdf44yGGUSSOTACclOzpMeAvLKTFOP6CrBektYd4IvfVi+WejILziwCi5aajmh
DgTOxSkEDrkKE7uylTvHfK4PKtxHPnVi+XC4uB2mzll0NHQiler19gNNQDOF8CIE
Tn16X9fPce6qjhhCiSlTeHhNSev/uGiA7AjrBPulUce3DHgieW8/VDKXM+41dfJJ
M9gXnnOdW+XJE2o648ChjCpU3cyzZpYbkcnsBk7Z8QPt1n0Ze1XCLFTSwMgL3abN
czSx6ci2grLt61iy+GSpNGF1kejQGbflXP5C/Anr5KkdUcUAgi0P2MCP/KY3NetO
jCCnXH0GFbMpKtScqxE3RVHd0xaD9fAuuNaPo1ypU2HgZhMoS8+ROo9jzsrOe9Am
Ql/OUMLm3RXlXvMogmwQExR138qjjBHoU6iT663dAbdzLXQA/FK5HM3D+23OvzIz
n05ynX6Q4PmW6Fqt16YVibgFUsbcO/3BXrOnfr39IxxbxYopz2SyUpdNGjjO2H+E
OdZN+RvqintQkKsUMvEMsNi5kWX28/KfHovJFJa8a8ACCQjOT1FzxwDSKCVAxsLQ
LHkIifRiLa5x3ZVYfvFeLuwKrjURGA9kINOVXpWTU0blKIjLrWSjcomROJoT0mSB
zW9RWw8bObb0vdGrWl2lVjPtt5ernPynJllhL+0fbyyfNsuZpbzEiTVTgg8bB1If
YDuFa5HAdv2L9Q3+Pr2oOEvDOoORb7yCz/mgDE6AnjhH6Dkh5uN+bCsiKNYfEYPT
ZmMfnOW7/eCqO3vKl0H8gmeqIF98F/IE+/5YuVllYni8OsCZhxOxOIKbSWNqgtFy
2vkQXepJmsJOrx40y0/tQfGGsDmrpeUTNxFh5yzmaT0rqQDxtkM3RLFceq6BMW2v
JlDSiROUx9+E6aShttlg+NZNSF3Yej0+OjtUN0JreuAzwrZoE2ww/E2OsVGlxYJD
7jmnSpohLP5602htAUZ4maSYmzwX2FrEDTJPH/mWKXOiErooKOwFM3ZnjEvfuDMp
5jegQ45MTGpvsx/RLxe9fRQmFxN2U08jDxU48ZCh6kbV1FsSNQXCs6K0rWNdDvfd
2+2xFT01HAEJ5llu3ejFK9WvWbHJMRk8GSIjTBx4Y/fi94ei/d97Sbd/F592wh/R
lT+RR7pMN6h803BoFxvjmiNvoqIBQuVdOv8VhY9Kte46HTLzIxjhhhWWDEGBITmD
e6YU6qvDKuJuOhv9GaoxTSIpu6nfgTrWwnJSLiXBavywzAqhh8ODC6PJ2hvz/fNP
vqQmn4XcOMRBpyFeDfmji/wVHeKF5H9FSV5mwiniSMtEDXEAGrwvagIA04S+6IK1
w8b6LR60REZo5rvZvIeDGnk3F1qZARQJ7mZ98f9cpUtDbtiVZk4zXskeieAcg3DZ
HeE6UUlM5FPwkpPEmQ4S+xRqRn2o/RXf7/Ng5C5XV7QcqY6IxUFa3oTUKT1gLXDv
3/pM4boWhjnb4FM1pwep4RRW1s741SZe7clCX3WfnSeqb4g8Q1mrpNr/c/a+n13U
Bx8mbZPIx7XM9ofGTJC1v5aBvj85HRiCMCvkfHiWmGPe9YCYyaeEEWqnLROLETZS
/YDqF4fpfMkFQp4ab5tjHVnVVUT4O2j/FZ/avcGO8S5aFSSBw7ibpjJsXZBYU2Iy
mAXx6qw0QEApqd3xwa545oqtmAcpIjIukCqqnWTI/jKzcrVjhek/vPN+kInktxez
ta9MpUoUVfeHj9GsOaM4f7T+f6YeKrgYHmMHoswP/1OSzRHvuZUTbOb0XMqmE8U2
L+pYk3PcQXwcUmiEIMytLgzGGpOwFKOAfY6i02IW3oBvCT1i2gLJ0B2pSLX9JhAw
usJBiXHqzBgWdZOgz7R0QZ4pgicHeUWtgEwg8PwMEpD0+cnAVSIRfcc27TcjHwNk
0hVdRo2t492izId9v5Soh0a9wbNvR7yH1/DVElhYcyxl6fjZ6eETwbyYl87mx2tS
2kI8s1xNRZb5mK5kV0rJQhwFge1W+uXm/6knT6zb81he1wCSzf5vTo7EBhjB+K6f
DK/alLzAcOHuSt54nLf4ROZxbcQV9uQxnQUkGnsMNmc+iu/OitbRoewbcMwLBVgc
RxyAmbosifrKfHorp87DnzoSlx+Ddn3huqnmVFJhuPSR/93fjGiSwmrHk4DLvBaT
0uAQro5Dh0+57losvpfeTN8CgAvMAYxL559d+qOBd3bE9FnV+Cm1twL0meKQ3Dbb
r+bqajth9op3+obntajcDRrUuYVW0+F2vrMUEfqqZocMbRPqhNSxZTEIxnzUQXUK
IPFJA5pWUoRIUQW6JXZS/vul1wBMmzrkOpFAbyYhMU0/tBTjxD4CadG8ydf6ruFl
+sdPpEAfpSfjV396XByl1RdpbYCv4ahePlp5GILLGtLFLTwf8qdUfU7R4XNJG8sU
7QUVzo2ITLZ9xJ3K8IkS3yv7DgLHr8U85phiXc9DothbaaUi80AedT6rIicrUVeH
8QLOZSxAsdq1e1ZgoNgrYQhLL0CYtI3+XXF5MImhkbylRfICDewaeikXGl5HmIxr
GWEr4DP3BM2f1zR8lTIaD9JqN6TF5+XvOn55J/RUdpuDGA8Zqe5LeoiciaWBAJp2
qb4bSQqnUzo0aBpheEXcKlJkbDzPQajRm5u9A8c58e7+y4TrNA/O3iI7MTTaPFPI
T8nsnrCSrd5uJ9A2REKHlxebr20JIPldTUb1Qz0v9GmL/FsmCJPrvd6xyDYWN6k6
w7mfuWiIhsTDE74PsXam0BCwbGrshf8YERfLQR9Rqv9C3HLAX6Lbe3atiupMPezB
9wNFcqr/IAeWbeMWUCfKpttqNmPfQQeqHtoYEDC+kzF9QSKtYgPLa1SOZZISz+DC
9VwASv4SwSUcmP/fh935MyIebO4O6RM56gSkKr6SRfl7hYOJXGbIGMr0QK9iMipJ
H6QSgw+g8nvZFDKAUT013IdPXpRmVjyD2X/ZNWtwhwyC1DOEmGEnVrL1CMhEEZJ8
xy+HWxp5+m6JGkjKfjkAYLFyM32eGNa9vUCRmT8QRP0yWq0MrBWTjokg91pEXChm
U5OY2U/4VgZ8c5nN6L+OiPjV9MTsnl7LNXc09d6wQaCw4XoJ4PBgL6peYLliq0wN
+utCFADTANnVipapTMOnFrrvDfzde8iuW9hp+xxNTFXqGUr1KoheA59wehtEzwuO
4cIlOpin+/TmSnOARSceTEr32OqcMPu93d+wS4FfF0sU4NhixcVAv3g87cdY5Pol
REtlCjVv+UQtoX8zefNzMIlsew8ORSVaFdqfyNLrvniFZXe6DgXu+iu85i5j8wte
1e2b7FphQBT/z0X0PDlKhUWPQUI2fK7NUgdTonbwz5D+14aLBW9kUIb0sRSkpGVZ
kG3I5RpwFp2jWpaXexa/U4tAKo9vWKZbJ6KxqZGc9ghhI+RCWoajUcfsXieXzTVk
IDA3DXh2GksA+AY/AFLK2srx2OxZYA5VcuwcyebvjfDMc7y4mvdIWRNBdo4GbKzP
8HKCPFLDjqb6YPLVzy9sJdku/O8Lf10201buXziqGNph9UdyMq/+EQ54+J+GOnOL
ZPcqJ0lNiCsc0fmXfmxT+9xnNzoLQI17w0yX4WZZMxBTzQ5VYPfjdHfG3HncCasC
0tLabyLFpHv2+xhk1Vh3o9VaEAr250xaGpAbyKaVFsgmWyAJDJvVpKjqmPNO+Up2
ruvyI3AucLWB8ls36V3S/xml92Gh7bS/hEeadHGt68+kCN123cF7A22+xMXZoPYd
TY1apQVWTskLtPG8+NVahSjB+L3aY/06llT/9lsCm1bCxDR/Xkbq2I6oVzG2dIiz
0FzDsRc+MiPD2HdMfKQsYEh+1VMLbbrOwkmbDYGXiAfpZdKqHKVXpTeQG5+7xAql
Cf5BZQtM1R89pOl7su58TCXR/zIKxAcKzcghibCEs8gFeCR2yLpXjCJ8QMjtN6k7
Y3q2oWLeH3F8mfPyXNGwnKhGp2G9Yd7C4zvFzUqiH+ybcLTkWaVDBRghNOgZQ+ga
IWW5J7BLeynOc1fh4OXcUDlcvz+aLIVTMCpDpajcjcndghoJqpvXc1+I026WFFAH
s+OegO0cd9Fb6EJVNmuWpRQCAV+RlNlHaYsO4uqXz+m4jliPH6hNmoUvyjE7NvLF
ChJ3Ko8OLX5/1YqWOrr68rwGSy7QaoV1QjBMyQtPzNVJfvpBMDgUTkUmYYtmm0+8
eaYm2/KyS4Ic/mmKmZw+CkW344AyRyMRmbZy8RJyHmURjflsQg66yNuQghkeiT8I
RX8cgH4g9+qH3PJIBCdYi1hhBjB/0OC8+FSkkjuDD+2KrtJV76e6Z2tsCxAuvD2J
fNeBoLDjiVw1gvkfwWAR8tgEUk3tZuNCGRCleHhgl8zKtNsCVZQnA/U1rKPR41u7
3Q78CILLO17ridZmn+I2vwJAGcyKNX5E5yBHJHTDdy6+kPxPmfKdB9w/DaPOMcP9
l7T3pdTrBWqK1vozrBy72l9q1lXpncaV9UUbYN8mYKy0g3XgkYQULCJeSDON0jBV
mxqV/DLjx9Eju5cFpKHSFZHnVdbQMkuGIaFFo1OI0iIMyakkhqKBfHbStAcG+q0m
5ynLaQOyFRyjy9OIDxXedubAk2VUwv3Pl8xMs4zv1dd6KMZ9XiuyjqmvWZK5fciz
0lHWlkwhA2kardCe6vkTPk8LIQJIHTF0bVsw9rbPzK01Cwl4N9pzL9gxhjsAi4/x
p5fnAmVRbdHXOufYAA+5ZmzvlaHQxv+QTDRRc7l/urCfQxQfxS4krZ6JUkt4v6tT
8XQ4QxBTTjOn5egiNItTAcxyBIIdEHEvXGy39s3foCz5KW7+xqywiUl/oxNtGusg
tAqSCYw8cxT8qKYlk4uA7xr8gJXLZzVDR4qYapK+5Im/bk+n+O5DvNpfsdnY1fnM
Dr3Gs5lsEYHNVh8D7xVOb9a9XqSyiV4hozWgOG6Gn/DT9H5V7yXWbOi4aez5Be8J
wcWl4e3SvCyD4TLAHyuVwZ6YBVHG5eEmAqDTd6nyoTfhKIh0gmZ3NnpjcUQDutWR
udjwi9bbTQKuVJQBtzeTPT2q20uyIR1c27KEvMQCjBdYyhxqFgtoOOqnM0FMDnQM
Dl39917FTaqK9nZEw26n60cEDiMHx9oT6QOwjI9RY0WHKGcLd6bEjWpYaGqoP+x4
DxbFFeuMbCHG9xL7Y2cXLKCmQaM7VkKlbfBH/dihanzjgAVXfSxX8hbuibrXavdF
TwGyFsI3yVDe+oZka/XOCy1zValB22cPGjdthAMG3BMUdryWE/gJwBSUQj8uneMq
+RKoHzChi2kXbSljqy1dyYds4jPjsIUTY3HUNSj/URrCUu2377ASIttvSby24P/U
asWG5cvN12xzn3hHzP8V/Iv4KgZRjFpNqkXz5Z/F7HUH9276QJ3a4ZheOjJk91bf
hq1M3xbLWQZn+8gGLB8a2IsuOPgVjJbU3cPcmlEP+OEsgJ8F0nXrZbYR5W8NKAci
Fg3X779PpqidwURDfaupw+rg6kQbe7TDisuVFzzanMAzQt5AOITGRrXfX5Fc1VFc
FDctMRhBv3Tpd/tGnpq9nDlEu9l8sFC6eWzNBqAI6PbVnggJ+mCV68fAVEQZC04q
fRBw2H4NTgdqDHmoiWb2KCNZKrFQ/1x9oOLgtS0F3gSiRkvBkwyx3WtDUR9OGRg+
NLcYagpW3EoQ+mm/IKxEeGiwshTEVXYeadodSnFSQk68Yzqyp1qsWaujgqDLZ84i
SwF7HNcPAVm7zUjdnDIEX2W9+dPeXGD9Qr9MIxd8noGHb+xkp9r5E5FdrLj6x0qr
elsQY2BUZVbsP51aWJrxlUJRlW4ITW4TyQ8kcmYPpnW0paBC0Pt8lF19HDE7yFN/
79PcedB2155oHI1pbl/KP4tBcf/7dlySXezRYFjUmqNuaL3GJk+uLAxdh2530LZS
zPOQhwOXT48qEx1493d1kMbdM0ifQB6fYcRjz95+rf+kYGlYg2J4rR5Pz7DLMdgT
IpXOMSBxQ1/t/46BT0CprHdNEG/C/NFteeH3EYhc2pyPZvg+fsnWING2JT/KXmoN
6xiyZ/JJJikXjhryFYIgd1U0Ajvf6m3yV+dFnOUi9RB7Ut906fXY+V0SUQeZjLk4
JpNEk1BaZP1uP5m1YavFjKHe4ygXgSfJwxD3X9Z19FuEWVzbpJt9YT9nj96dSm+u
d2kVfH1oOKWET6WOegs0/Pdf2pnNfnCj855xBvFlKltkyZdJz8VCqHcPUdQEsc5y
IHZfH/ooi3HakEnuoDDYmhjuCm2iZbfAJpacxBJBr/vif+rH46/hMugY6pHIUXih
fPO8KfZbU3FeDYA+rZR0v805V4UICLq7zO7wUtn08cZUYdMpQu1/H/SrycF7v/a6
FeN3KIlsQVZDDX2vzIIm210aXvWShJwkWP1/8QlFhaFq9Wyqhz73AcS8ZVDDVieN
vQNBnbe0ShDHxjwtq0oREq7gbjKIhTeydJ4buJULj4Q0l8WoRcq3ekHPLne6vW2b
yVjRJ0RsnBQf1ciyN1eQi67jtvEHSqcWBS6nxeGwqnARaulGtiS9KDfI+AdMjHUy
kNZAF+brzbQLS7bjqnCT6va0MxWEe/J6/yCx7ZrLImwSP3jydBwhpVd9B/6k3/GR
QNWKy9kg3eI5AgRqnMFrRUaOGwGw2lSGAAgudo6VeT1kXWMgvqEEOeREbjvgDkSF
52u1E89C1Rcm5m03EOeM1xoLRveGveNOI+3sX4EXOyTQ85oI78M72y4xjDR2eYuo
tujj8ne11LeSU7xUzr3GSIO9ILr6PI1at2Bh1uZ6vjdkp4jdhroe1dZnKr2lzIYn
yN4Z3am4IdAxCuIsQ77Cnqwq8azs7KO/X5PMsq4aQca14aSwQnJncaKp9P0S7tqx
SeJvm+qY8dnOOrZrqenJE8tjYhHzoLp8JJWvR13xJzfmlY6VImSNCPjOlTPxEsAM
/vu29oA+wRSv8kpYJ/pQUDvNwgZYPCYLOrQqXuFA5QhgFQqQh2z3Zm5v9Qvh/Hil
fosXUNt/0lP6B3qWd28QA24pHLzSdcSMU/p0Vx5g1friLqWFAehJiF5r4JTdUo6D
P8aUk1Of3ELzva+kTaqNRya7A9QhqqvekPeggzLJtz4JQyZegGsk9S1iKcZ82wwO
hweNTDBPsLmyuzZIZne4CIBgP/hyURQqEUMuw6a4DpKgKYb4RZa3STXidnz4v7Df
WKk1y01ySX3ULik3GHfmt7BaPHnDSIVs0uPnrKOjb+4ME4e4Xhxw+RghaUqKCFYr
paxNJMOqGLj+eJMlvzjmlHICAtoQElF4j4ZMlPG7RVAOEdCbdCQzZDrUXwSLr5fB
2spAbRXYSoIoU67KgykbuVRfpGULAkaBsYgOfbEMg9rinrm5wEMe+083dXnah1So
RM+TOlLx7y6iCVJpvZ43CaQq6cTGCjY1Br9lH7VMkH2W57Iesc2UUZUSIBNMT4MO
tF8+A9kttRNwaveKhl6FtL5XIY5fquombDnq6/738Bg4/3pHkmGqLKx3wQXDCYNT
nujnVpQjBwu8k5ogabq6NHAFU7FjOJCl0NtmjH8HMxUBQY1C2NuHDU/isi05kkVY
KPstFvlk1qullzs0hEUzBpoO6OF4DmAIw1ffv8ES16oSVEgMzbtVi+I9374bSr9Y
HPW/pBuyybwb5u9BKGUIVXA9PFTskO8KTUp9joVtSbgrlu/rONOlI+kKzCK2Awo5
XVnbqFzAP446CH338e9Yiv6P3VcMaFqnzFNKPUaDxPGBMdVFLTR6wj9NOIQYyq0o
K4OgALhkh2pz9NQtbBKwojF/KrZkU0QDalMML25qg9e8W7C7Ffe8FsQ/cdhYnwL1
pqNjhsG9Zq4ZKsFo0KRfb1YvgYRJSp71SkqeVbhzTck2t57ZYWuXqbzOzbWZpWO0
IPu3NUMIWJ27yT3aSMTQST5pSx4K+aEoOsS0qvfr1glR+bTePAHxy/X1AiSgTlAV
ssp5px51swOkRXbDnj5r6YbiKckLJ0NZjU7VZmao4inFskZBT3jyNLhA/z4G7tAd
uSP9820v3+vcAos6rTY1aopFVgyC0gekDAslvVPhjPFCfuCIMwhsuTk1BuHGRUbr
Ns9Qim4G0tyPsulKF2zBBPPSw9BOUJhCWiMgxmXIo6O6+ms/Wc3pMu9jRIX8Eu62
rKdS4/sjAerP6mR9Ngixf1Pa/z8ACI1cFLw/AY2YFXoUZykywrAwzIYY/I+6mRd/
aWmkQLUlFFuRbo3SO2CmodgQH/d1vnLMNhC6vyE2bH7E9DIP+xys+bdziKDk7Igf
7mbVWzA3J8nkB2WoWvOnz+feF8+Hk90DrIj2dJ3BE/VmZhDyCQ015+p+F/nxuDdV
x/thjdvP83U+vdnCDQ/f2QeNuRLRz6wcJEELOXjF0QkD1AGPs13cSd3rqwd63zfm
Qk4hIn6PsNEtquuEJwzBnkEq5Hg+vE8y7RVUgsQCyl3NVIJEU96FM9wl4XP5D+OR
GU/U029l4UuFZx3D7KVUC4vslDnqi84ay3mLu1AXggiSWZZE5B/iKpeX+OZC+3WO
LioWMJ81G7atXU8siVD1waxMLd7+gqQYwXjf5moZck8RUURcw333wAIyBxOaKRZc
fdegQaf6o2/xFf4mu4B+2lceji8ACKRsL6l3vAwok1rGrUkQBD0DZoK6rj2/0OQu
Ya5RMNYVPVBlgLlfO2EKHhVjabx44vvIHF3k56oPpb0EnQkBasuU3Cp8ctxjbDVb
SbRV3QhmGtsfxGCQXLX3dR8H9QpV6Bz6XyX+5eErGiUllvReG2Qau5SFSrk0nIrW
/35AZcBlxhT+6cL+Lw0QcL8B3n9cGxlXXMTthiTtx3imanwePJgIAwz0icn7ghxI
mdcEL/ztt9D6Mr9EWRZUu8CsBx1486MUQwBw4eNKt1YtjVHPjx4e91vBoF7xJAU4
zYeXfS3MveZZlZdMDpQRnhgFTwapzIQ2MArpY3Gw84v1U6afd2KoAUckCJvMxFno
vq+wC2zR+Txqk265TLwWPHoKMuJaI1OwUWy4tl7BGWVX11War2sSIRrvYeF+F7JQ
C2wlvw2IiXheq/Oblcl9IrLB+0riq0/8QYAye3SX2y9iqb7ElYRptMlFEQ7xA5mB
gAghTpjtsLZNdJjnTXRFbfEbPCX9/fU0v4RyVwFrPbTcdQOp1jRSmi7VWUeozJJh
WClKv1gNVr+5sNMkByehWEab2dWsvt8Bl86i9AySlCyJPIBcdi7MzmKTGmb3NwAN
Z59YUpgRZoFEU5TdrpWCxKvmbcFAtMn1JixnGIgerlP+0s3D2Aug44Q1uuLHWeM8
Z9IanFH7xLYB7XrM2bkwBE0GNpancPUmp9rvlYn2+kHNzHLxfM5uo9PoT14ymk75
gGaTmgWddzhkWULvUZzuyCqwOgcqo3qJGZvxwG7mHwhbeQ/i1xo8uw1sTa45OPg1
JEzHbPIfKjefzoKHCqzjVA1cC3Z2bAmjm7iwr14YMjqjiiXKlI4umsspnO+W6YIc
TH9kcJyLcWE1sDhYvRMhV7Ezp6pblbZ5WsRSFiGOo8YKQSJCoQyU13/QiTb8jkLb
gJmFP10PJrcSbOWiShxGNBQtY+Sh04aOxEJv245f3J+JYB/O6WhEzMOkksYrLzcz
68xd6Mudf4UXR6oO6gQVVekX3cfTX8XjqMSv6MjpQaR7iej+K/XR+YRxIl+yzGmz
08MylEI3JTtAtJWY2rITDi9IRKJcKEmk7uEqWjM2QBJv98AjNt/AdanhijiZ+UBv
7iMTn1uhcDmkWEItGiCmTIR5In4lSNRhJcx3bpymgbyKkYFE9XJzhoZxDzvGgr3A
+zks07myScSmkiEd6BuBGzljdDQ+AX3ojYBZaPB5hewzykFAbSFEgy7wl6cODlVm
AWlFMoVTKG3xtwKZCsd+c4xTsxiOMnOtJebMXXXx7V9yD6O+Wr/7MaZAEoV41hPc
6JUZcvCfQBjYmQRM4AjNKDWp9IFk8np4jpujKp2JBlXJ/sxphhGzNx9olkx9mOrI
+4WestzVXJyhd9MUKqUrH/OzyL7N7kel33HUW9geYElP5Yfqm3IYZ7cLK9WLnRPY
io7kuC/xO9diJu6Clj7NLDGDDqZ+uyNE5azKkowsccSjHm5iSCkybL6u6XE1qxWK
p4cXI1Z3ssmga69Sg3uA3nn5Gc+iT9UfeYe//GHP9PcGiDnVKCOoEdDGcS/iE920
CZabkwLKOBnMEOeEfqP4vqSKq19Am+vW3RuSlB+HPSWYsocZeISfREj01uehnoyL
XnV0ijMEktPxGJ9xf+9WSuT94z6dJgu/fFeKZYez3lFrBo5eNLBzBvF456k6n+0N
X84Wdz2FwDHW/3l1Fnq4dRlChULNUvtamTKamja2xULaSmbGfkcWO3YzNI5UQDvw
4ynBvRMRQ7uJbXmWUQA2sbDrCHAX0lHb4ecqZOxb5mUcnva6qOwBEoXxI2KfKbSS
WfhLVF0UIxM45/YEHwuXVjM2HIs2uqCoQp4gVseX5NfMUg7RN4Obz1KR37HtgycA
fdKsoa00SVi6BX00duV7MXHqadVjs3NwCetP/bpwldj3VbEizH7kln7ygLPmVKh+
tbX88tu7TRGyQCv30H6zPyuhvFjbDVmWWRlAClZ9kBBjJlVz7Ws2nlU2N8oTjcjq
FzorGYqivaMhHYZxYps3QUp8quzhbFsNXD6ADoJzgKEULt0xthA/VoIlFoHtmX1z
k8DFF9+gTMfPsHif5CaUAT5f31BY2xX1TUDzafMyRqUAKD14vShYFs/s1g3qdNO6
8QYFN2pd07TA9AshIdCjedn6d/kxyu3cZILtMFFUBIbMx8kfwuTNKhm8Dy1XLVbM
qXMqcYEyn+05K+UGPuj9eqQ34wNNM6Ewl8yDnDKvfdN2bYPPyn0vXXjM0lhNrmbO
ILI/ZECQSE/R9FtIQWll9PHKsR2OOPkTcjaKx48q9ISPv9jHfDD1/05ll+uhKLYz
FMKkyfJUnVJ4oOjwRwEVzMD8ZrPW9OIAv6E4cLTlVX0a9/ImhtCcYaYR2lxBiQ3f
ONzMJeFJkuf+zWTx1V/QJMsbtdQ1tnYWmH/govpV0QtZuAkIEtdMIfhVcX9bGso0
VBIkaIHyOXzYnN61TzCmSf6Inz/viSfEe4+AfrfdaFzEcH6G/dQUw7dvoJIQQ/J3
vvOkVjRHmRZzG5v7BBs7LWzVg97y3i14yrPVjTKno7p+QYxvMc9k3g7jS95HploT
601qS23P7LwSwLHBhSSsB9pJoyGEHZ+ZLmIkO3OQFP/2wGn/SRLWnV8WOZlBxQxf
gpK1KgYooBrq5jLxg/MWRxfTFrvFhfB6fXVGFWL5I1Dse2TXCX5V2fn4Xtksbo9w
+aCHJguw60Vv0jm3C9sPXf39bQEPG5T61Fjd6c/ATuLErDPz3wsmhCBBu2eM+Jyz
7nm22uGgd+dwVrGCNgN3PkY1kBTEv6Z7hrToBMmyzFA/rEsr1mUGW3P+YdaTxsJT
nuIyDHnZN/e/Wv2uN8XF8/GyRQGPCj2yAO8AOJFP6gk8fOwQYKJejvW3REazwaLY
FoR/eI+eCJDQnKWOfVVEB9hAkf28F97zmqyXAfStkA4rELlE/Wlmb/i/rBNc7TdX
CM7AcnDkd0md3XuhRH0GeVmyjWoTzSshqyg0rOHSe1Mv9Ne/X7sNO9CWI5DmAsxr
vRqE466c+fHnJwjOUzBKS5odMyMXIwBJx8RKlnHXAmQKle2TG1TmvQlU2lFNAeX7
tUzLw6J8F5erWtPQGnaZ3fI/bnKe9jIoUDbdGbfcmys4j5PtVyPqU6Muf2RSmpZN
evdiD81XUHVEtSZ7zFTDtQXJa9MZ8Ou8w4sP8zol3l6JP3kAO/eevcs2bx3Xtjip
vGI0PeVc1MPdYRyBvvYH6zK3zCpNl/YCsn+3WpdmtENqDQUC44ksZZdtM2dyrVg/
MWAfLuJ1YVbdvVmtoGCu8OOOUuW76ZrDMcfQ+EuDyBG9Mn7tDA0TEPNJrAfM6kEe
M4FJK0z1cCh9JTjiPGJvPk5QMYGmjjdxiEdnN5UIctjeV2MulEabhBOxW8qZVwNP
zZ7cH9vWLTYGd+/1cP3KBU6YSbWMjgKJwMiCwG3/yvf5aztsrcqGgXxMdmlS04zI
yXU44ipS93oGQD+/MQ/MgO6rS4LJ2d/s4Et2TLG8KdVBua+W1a0jS2zJVWocMGYU
Lg1CADS7Y08fSAZ9oXjxlz8eA1K6YcVKohE0mJYuNJn3juB3/pTiiLADPruwub3x
dw0YxybiwqwcYuUYOpYjqN0CSByvLJf/+godv1G14fW9apkqcCL/MkUNQ/G31eeh
PQY357mxCNyHl/ZYw62ODkSC4JDCP5fRVGR96O5MMx7bghnLNtlIkCgdwi0nmRqF
WthdkawvtXXk0PEqi425+6W3wb7mMJc/9Uy7zmPsca9uGeoS0gKiVEMQ0+NuASGL
MYP6bEMKDhmp67Mla+FUzd8dyDLi7a0nMlWqCCrN0orHl8zxeX0/+fzHAgyK1Lmx
V9/bbPnCk+lsVX8bRM++q15ZX1kseBf3QqEKGHEZiF0KwMqZbPdj/F2LqIzzpEZs
MEQ48xHTde9kVonmPHLJARGvLf3qa8Uvo2XeOKAHNdNq40iNAinlM3VT7Pa7qeer
WgpAKXgzP8CznC5ltHsliLj6w6gbztuJNURZoA+BY0i7KgJHQ1TJRi3cZB5Fl6Yy
0DY38Vs5aLlt3yl76HAY5aq4zHYvGBE+gnRRVJuMV8jG8Vik60OoQqUJ9CfXbdGf
yzAR9JTMYGP4fxzip5r1XmD9kvhGCHp6unyZraQWZqIww4R6cUQ1TdGfgLAkqFNw
pW1Yp0lKFv5lo1op2Gzvyl6CLi/6jxfZ5Wc5Z+hc7aynuL/88cRcf6aMlFc2nwGv
uURbeDmf7uMyAYtd+u5IsZaroVvU1n2u8GSyojWkIfucO7NxmEkXpnVj9erPLjAV
ZpZVx0VkeaYuMduHG54EP7yznkNHhx8ul5J/jCiCPxnwI0PclZ55KtkhgpxqETc0
VnungB4vJoPmO5JSP8ggVJMyP3gwO/gzCZu+W5EacEV77R1fhA5Rig8vKnz0CUvR
Bm/hh5wOAMADbosTumYROHtJMYZqQj92z+uYAcggg4Ve64BdroNFkrRcUPx71Y4c
kanNjLMl/f534aTer70q3bxCyredPBbamnrPac1B4ppUS0XF5BfWsvFWFJxMYvaQ
mTni9nhXScaUfj6u0inInN0XtyLhTearzuut21ww39dutfVrOuQL/sGxTS+dG6aD
1l538BDl1wAqJUFwwdMC3iv3aDqfmMhHj9gDPWW0VcyfZWJG3VEWQksF4xltf6Bp
p4B5IItnZJJ1Y7GsRbxyaUECxIrch364l4hII8BOSjdyXqTFyF5lf/ta0ehOjlo0
es1ZDfVcVXCJARkkys8W3it1eMGwucb4duWaC06+DUIjEU6degavlMX53pNy6C7P
BTvOLOY0JaaJCL5GAFI3F48wgIPzdHV2FQmL1JUjj58EUo227PzmlxPocm2/Ic3/
Pfve4djjnDaG/42gQbXvusc4BgV1MK9zcONZUAikHfe4fa2VR3RkvRzedIduCkty
nXM/JIz3GoaWGfwUXuNX/4LCU7V+ot5pRxwXnRvVGjt8CAXVYn/6Tyv7XkXZVYb8
J0zvc/F3dPm14GkREOpfFcMmf9YRl5IC55rGuV0D1homsUVpKTBIIcxi4cigorqa
EkfvDVQ4UbQRNyKCWjSGT1/w+5ehQ5X6TWUoIdZrQxyIALkuXvpXkqHqzQkYQTI3
vSmh/3fP2tlE/fLfVb0an9EBR8QFvdxTLQJOnC0WNZD15deB59EfFkl475xpz2YT
bSRR7bU1inaCm3xlwCfqOrc7mT4BSH+mJyKXKpueul3rFzvkkunWwa028V55NbMC
Ia4wzRew/YoIC/hsx1mR9/bt3/Lm75APba4/aE2ffCG0mJpTVbQKq3rzPvUzt+W1
y3ikiArD4BRcpzv80wldpt1PBVsRrJalKNum7sMchzxFen8fbwwX+2KsxOJhmU1S
bAwqQ8X706nhm+gcgr9AZyzBxKXreaRIWKqMPwOwf+kU73p+IU0fNwjUi1NhjArk
kigGpr2Qy9kUXuSf8TB8rhaJOon/k9PTy4upykF40/bW+p0yDID8uUKyha4nKxcS
nrB01fyERE3FLNzI9i5ZwKwdvs6NS81tohRB+7XamnIroaD5OFX0jWKyZ3l6LEJA
M/Up2ksZxcfzthIgbZmfGI7+DoVs8cEb7MoqzRgp5g3mJ5pOkGDBvsavBpczIAIt
vLaOpxkAWKpfySqBpQrz9C7NT7zt0rIqKwcVELrC/H/+EMoKXlUgix4N0mtWbjd3
ByixEK4R4mtwoFt4EcApbi+nYw/nCpqHcJfRd5D4u9gvaxJ0yurBU2XUfkqjzou1
+ogqtzNQBJikN4ul3jmGdG7X/3jl66whAfoa/Ge7I9xzZ4023qug9G4quy0nlGP8
0/LKm+pzE/gp/BplyH9Ww94vCdkQbhCHvjwebU/V8GiGZ70UipwnxHm9uxYTKMm6
daNhDPFdGXXdH9DF6hxj+DX9MfvdDIlp6DU3uKTQtB6mJptcwCw00E35ZnUAfoHz
4tb6lGnGJ4Cal5THDBGG1W/G/h+T6D8lbpEoL4cz7RMdfL8OMELaXsbHCYPEUKxr
GX9YUDCJWxPoBcLCyTtf0X8voCetG6Osfu8TKso5FKp2W7CV7R+AVxH/I/MmzKDR
B50T8a3FXmsoyJO5q7hodpm8gO1EcOlFylE2ALGrrfOX103lHU/bdOOu9HbtaJZx
y2JSguEF7SUHeudSbmbOZ3Vxx78XxGmZptzmAsjWI/lcGhLssWM2xHSGxSwdZgOH
e5665fRqL8eBaUbuUO/CQKEkZhlGN/DoQSVT0looyl6jb7nVUVntba/Ssao4tTBv
aXBcli+h+tiNVChLSe9Abwon+/9m9K5m6Oc+kJJrLQQCAcPpSdNQZpwEajD9+2Yt
G47MiPMizgOp9ZqiFtfwvYaLLdvTLAU2XoTc3pUb2plpwYZjaptHbFLyFoeaJwVx
pbixeePWKVjAG7lZjeVpyRi7SkdIWv0udoNoLND3xu9mtfv97szBJyx6d2mwsE5p
XVCgcFh9d0ZeAAE/SZk9tvT/uFq+9RoRxqdKa7ExlWQwluvPgk+SNTWrDaWUK0kH
Lg/pp9rcEp4aibMHLrE4BQ6MANy0gn+TI7tZ7KbzsgBVjj+NZahd+oOlk4oGhUCZ
5EAxLPW/I3LJyVo6YPJWJZxHidENT/xmPyE9k0e2rPH1VDFUh9ck1ufzMOEnTzzn
nSTLBVEG8AiuXbRarIbjKEoXtD5ErnXPGhafm5/OcWcDt5r97udrxXiYuQ8CoL9p
ARfnRlT3oOhnUlL3jNQFPCIS0WQFXekdfWERGk7nLVbnpW7R25q/LtjMZmzrH9fT
nudYJanNqqW/52q8z6CMZuAPkTs2j6/pCAP2d3wKvTgritKt+F1qgMZ2NXOU2RRu
aNZIidHhevlT180INspPwvh3LUNWEZZrHfb++POvHMrYZtr5SHQDUxJcB5/BJHYV
CGcVW5XgB5/Bb00+jPlq1nDv/eQTuY/++QfF1zfgGC5Ml3S++5yBBVjgtoMlsIQz
8MjS7SyIbPn3PzkTBaNrowIM1B6hkjDnpjnI4MPAMgXlMFNkfetqtOcFbBvkWudB
aPUmd6qHcydyG2kDuiQY9rQ/Xw0UY9z7DBUzWQommGuMzVX7E9qiE74cPueP/h0t
q5TG7pi0vFDXhK20DSafGf0HmDVykJJTtdE08hR0FFjHxhAT9oQl6Q0JLeXqVxrB
NkbipROyt+35L7yq95U9c/Jesb1OGvtILTgej3iQo97+DfI6/KUVBDpqJE/j7p5T
dnmkI5fbSPmYgmKdmLBXYYB6shym0AAPvXo9l6+c740An4tnRmrZGwUZU7wwDkyk
ED9YslEysSgKGP59K0osKudXus3bgRp2d2zd6HTeMIrdYsx2mZVkWzb+pp521S1m
tbyGE4rxHC8jCynzkyJHLouuAqm2gzG+sW+KyzulTPvIku2Jl0rtPjyy6zuJRajt
k0bIhILHxpoAfPQ/sNoa7TBpKO0Wv48mRK64hlFT+1ZaL34ps6WX5HNA+yJMqecS
FAJMyiQ8jsZdsZOsXMvQLjMFxy+rw6fUBLsbzuvNWwCj95tV6A+WKhOmJq/Whj5M
FcpFtpyy3vqsSEkidKWS02xeGWgFklqFUoeZ8tak/zyMT6di4r8dBDFrpuq5Hn6X
kylrS3XK/KcfWKuSDPog3cXyxYJe3et8OkdHTSC2mazMme81Isg8/qip1/7AEhum
b+Smhu752cREIujHCxhv17SAanvvcv/3AdTCJTGCbHqPN6+N8CiRtHIKQAA6ak+8
PB/tNLxWRviQoL6TeQZmCElzAtes45y3pHMmAwhvFWvgHsDBd0pLxBEgRGC8wycr
N5QYr40s6beKNSSubm6ZT7l8TKa/+mcAkgB+6zOJ2al4InfuALA04NImnaspiJV+
rraK9vqOnYJumm106lF4w+hB4GNlP4d172gyMRsRWWbqH+rYEORBokp/hVJWOToF
AUwmLU8eWcBGAZBZ+u8NTLDP1DDGSRjNXkycGFia8voOGuooBGw+ixH0iANF1ju+
C8CbU0XKnBm19o7yAoMJCq+zSESvXH7DCPYzs0vDxisvKlWuwFYXzBSWoYotN9ms
eCpRyE15io/W6tkPodafwQ5MAoujBjBpVQuoyjn+wVsE/QQRl3MpAVTWhJAvknyp
C0C25VF5Qcto9kRc69Gvkr+3RExr/YsiCg87tVWvazF04RvbP49C3dSvYEHXJhPM
8XX9J2KOiaTyc5TwezeyTj9VyUBZTmhMOCaTivN6gxsiSwC3kgggqehB0HuPvlJf
0Le0/CXGrUhW/RlnQdNSOX1UM89z5EUQUomv4cKb+2v0e2r+hcuLpAPmHJEqHBze
FEqM1n+l+kLDh4LUd7h5D6rBlFdtQjMaUODjOJ0eBESwvpKk88VLzC+C+3lKWx5W
DL7FcPymhkdG7FgRmqJxjO0vlb3yqqG7bODlQx9sjgmnZP9OtWZLYcHoi2oafh6h
56vne0PL5LA67QWc7IlPpehba1GS3v4QoA1JOE+oSSAdOP2tlafmIlfteJXRasXH
Cep03oOIKpvIF1zJsDt3I7Znxw+jk98SHnSD3YuvUezxL7Zdrw22yD5Wr+iXihw/
3kdn+8jzVrlgK29llOn4IjGcLBR7SNaPv8O0fLBxxQvlUF8+4NFITnefhB4ZNJFT
O183evp2y/OFjF1fMah9XOr3xysdwAdFI1zZMPuYVmV9CsUt2zB+OUGlztIQrgJC
d7fpgWe434DbYdPy18sfVt/mEsXJdt0CmGexVGmE/wcSd/epBvCwjtkBIE+9SZE7
hj+L0FOuvO2QjVs8gMsy6jCL/gV186kHz3+RwQ+dbHVuh8QzvGglgrRHfm05DH40
JD40z9uSMJz8D2g6X6gWkkX/05jDuY+2d1TajRRtrr1x/kkWMqCmsg+rez0Z4GSb
MV9B/Y/oha0UUagmpz1UeZogu29kUYl+uS/I4rS6LZledcHh9dJjEgXuymyMBcWd
QgWX5vIpKSxx9CFLk/WLpb3iyO+O5jtfDaIEHmMq2aRyuNfNoe3AOkJExWTWmYtZ
WMk2XFbxbYBCm9iPTAjU13nYszaWgI3T78b+sFPmWb7rXz3U8Hw0T4xFijwoufjF
I0zjdYOuY7G6c0zGuMTVYdljSOiwFgRiAsdw7YXebCY+HvO0xoenWri8CwEpb90v
usIUW60Fvq/2lyCEQ2eFu1ijatSQKGnJCFF3gX8NsbWd8f7kVys0YuCd2KFvd531
Wq0sK9iIrf3KfkoaUsmedVKA7K3IFbKYl9zYlWM2Q0pXF0Z9oEAql0By5XDXzFNl
1RvcNcxe+NxwkmA7h4XpF8dvJrilwaBxtoTFSxZliJWwnxUM4kvJo6y07nWDfEzN
WQj2geJeQxxcIXWLr9Y4yt3TeN87eS/8C3nBCY1uH4BAbxFCQSogO3Su+echA7wD
ElDwEd56OiIzz6Nh7d2FIX3WhUpJFj1X4eFTBao8PNxODmMNPg12+AbJCdT4SaGE
D0ICY7V0W2qVwwVCH0Xhs9hxYIZ7El/AO8CbK4pPlceHUw2KvWYAoa39dTsp+IZv
g35ZzFdyHXPPL5uAUo+cadgXX3d/BkT+h0hMtUYSkN9rzRG+fSioOLX+LfzpfHh3
jHQI5ZRno4HYP83i8T5tOSmvKv+BcGqh3fBD46w+UPyGJU0NWXhT2pWdw5OOk01G
Tfu21pqReao12NDDsEsAOHQ2wwB6whC+jl3uX+Nr07Gg6Ibl3lXNWboHyEZv4sht
cEppW42QHdO5I1xkSP1HRmqnWs53lEMJ1jN4wtKN37VzIKq5092JvdYpb9lrmtFz
xxeovi89GrqVOQaBzF38Qry3GdgRmFPowGUbLCsFD+FwfEGbRKPcvbOLFVcwnmC4
/BbNvxc87VGbWnn+UtDPvl22ZOcXesqJcZN4sIkCvKTa3H2Xb8tumn4h0hegA89l
q8vTmIJEQNyHSVaDfqOwqW11KiXBQnF4jpthScE8rt2EH6lZKaVG/boYFxnesIpr
T+nu3R+D4lw5e32pSDfwJMayaKCKczcvjLKhP53SNEWzyY98R8eviRQrhk+RSh40
V4oPVO3nJE1s+DqmQp0j7sqQX9hGjXidVcBfUNTGRCwXzC3yshkYL8u9zCilhFBK
gHwQQxgN6zReYGtA0yuQpsV65pwBxDHu+8L7EJkH844ahmjqhm9uLqjGmWQ9NydM
GevcNzi+VW2D02HEeWh3KCSRoY4X9rvMwEjV1a3yK1hIabdiKm2zvurc0WSNwqi3
P3urvcBsggCXF36+oUUbGhEO0W+Idietg5hfJfflM26phBRIbtIlIlFSVLd/dstv
fBJKuJD0fdVGvrfz3ZCVTr3Lv6QpwI5OIHnLZLJIpO0mBrOAXe1HgQ3gJygw+mUA
ZdwLGf1K67jSiESbfSZmhLRIYOMLA12MTezN15+eQ0Rp/NrZdwYYD2sM4gypUwKf
N5kRngGhJtF2zjcl6CyVM/RA0H+ssDFynmYmEmXlpjlgFsmuy+Yj4cHhBIvx7C1I
v+fUPcF5o+xjPPMhAk8l5utvIWmkDtmm4Ah7cAKUgDMvyaZb8ddqIjoFAxu1+ZTb
M10h4xJf8JgfUBrXyctn1YsfbHg7tvscvMuouhiZu8e7zQp29uyjzrCtuwr/aTpF
IKQoCBhzapFOEYSBLJmpOiC9PiZyRKAhOv55RHLsqtrfHWuNsKCxdPZ95Ziy7VrT
VXTepr7FjuvMB65LaqB3+hhSQdb4ceLLpStrkEL8ayS0e549wZComLb91KQQcOHb
4yjzS5qXoDXRZm90YpesXU8K8pEa5CPHs9FZQ+AeVphxYu2QT13enG8UvJnjL79/
rRPsuZ5L/hfUD8TL+AqDtOrBgpH81rFOr7KpzmYcj0ewPLpir1/xT9oBP8nACQga
mJsU/m2ho7Q6FKYiWMNK6eGtUo349ESKLw/S8GSwdPzO8arUOOyUf10pCeWzZ/pU
f08+9wdAlZCS4kS8JC0pcyjoBOz8OWvei3YXgHrTj2/LYKyE607lMAgWhLOj1B9+
9vmZEnfKuVWI7H4cQ+mh5syfwOkd223958qJ3sz8FkXBdPGYbXJR/ETwcDX2ByBg
ZJzcvlHOrFd6h6513oDdPKmBvg/wdog+9UoakAB44Op85jeODNHnyAUkpOjSs80Y
FwVupjoiQT9XFQ8xduCAy+EzJRzvVdGyqdzGvMxMM3FExZ4YMyJacb978uYy9YHA
gnr4YQFAMQUcIsiiCu1Cy9w6uwsvR6zB6+WSdRvJTXaYaSnIOui7mFopsN4bxIyz
g/+5/ch296pr+O/sMThLINiFFTg8wfOpgZTrn6OYdyVmTBpOthqzJ5NERo1c1wjw
3pQ1968FUdCH7/rYqAEnXW6IlREZHBOC9Ueo5qFjgW7sYMxn6uxa4+sMI1Wqy/Lj
KaNJijDouFPWZrHpnv4xn4gSzgNLMOq/l/4CnrVfWh3LuePR7ff1IV4uif+UiedB
IRVyoFKzjFs9Sfi8Wdk8oZQWKSB0Wt81YP7gUDE2enXNg1b5jPLBP1luGRKPG0Qf
IeDFHI8Gu/P/A77GLQiCUbbzRXV/Cs2yHMP/2ac9UVhGqDMkpn5r+EoEGixwGyW5
/Ss0uoyoCPSY5GQdFkI+SMAOTOj1JDD2GLkpcI8Lx9N78cN03R+vsvjxCRgKShS7
FcIWE2Ksa9izkZ0GMMb8Hwa/FxoMTFUQ8mEwtcslQHpW1JjMIVtlFci5q5+hXFLU
MzCQHWZpLOFyk69uTHCg7UwPCUwYtkrQtitCJt9mY9/OK6kOBV1bLRCFE7DVqM0v
z5u4ghKCen4ZgzNAafWiryVlWi4irjBLf8c6b7rRBzOAhJgo6FIKs7TLKYWUwKee
U4AeSKQrbNLQy+LuZl2lQuR6B9ESUd0bHsZL8Hb98OTgWE0fozmshEljcyJ5o7sn
fmdBKhjiJDugzdtWRju9C5gQPaaT7dpCODlg+dbbkoFqOmv0HsyxdeQb30uCYiIv
npwBP1aCgbL976CIai4+ARt75RKzXi6S4V9ZbFuwWFE+pZ/j96dB4XD9DCLyWhf1
4tEZ0RcnO9t/h/9UaWd4w+ANSs3rotpbal12bopVtVSBZh5JHfq4fsd+q13d3lVE
FTRmm54hPYdv6fKuQFiMBbL6Qk4fuHN5RGrGOLgP2+mMbKyklJOQxBOPKOJHm6Xr
OPWkosCujWmm+K2mhXfYr1S+z/+7Ds1+W3nyLEVWGFNzcwRGJ10GLhz6FIof6wac
gajUao4HmMVt00z1pUklLFi/L3esF51y7CHz7zfklHzqYxjmTehE/qGVA19ZTmfK
eVfkcFzKz2NKqTBJVY+YBGm0DDohcvsQu38M/1NnqLUCmYN2+PpOdfH76mHKffS2
+kBEQPI4K/6n+cGXMR13HzAMBjHWZI6EMINUrwlv/wDGPgR4CSIMBT5mT0XcnaDm
ffkeu6e9ksZUA1BDeNvERWLxIlbK6AIVd9VsBhfw2lYyeinhL3VouNGtwaYw/zJm
LYW/CVhQokPs+2wryMVZlfbdbhBn7LgOJ1Ax4/Ln3T9LOGJxKnrzY6K1E7lN1vB8
Z9gQWOAHal+tFjZCQBPAuI42V2e9aU3AmQ9XxX8ZCG2OjfKPHSvpUfYw0A7PQsjc
HTXMLR0XFaWia/k9waZ1UXsWN8b94+9jANXt9xMraEL+p3H8yen0uqNcEk9VxWLq
ud+eOYE+EvnD7yR5IxhwliVUmiENvP3GuMjGMaPDk+c005u4Sbt5YEY+wVOZKoHT
tM4AG+10eOLBCXAcgXBgMhOBDRNWvOd7kmXFYVmgnC9ZFANyMRwvYqN/VONR1Xq4
wcpIl/+mY/GkvBr39ATEdd5KJx2GCefKThtnVwQsUjxpxC2AyQvm5zf/PwnLVjkS
tqMZyVZzYtcmQ8lrMYr6YqcP5l8se6TDbE6jH+1Sn2lo9mR474khnpJ+vNaHdNyW
81lnE/z0paVwUIBqOQgWZytrjKgB7TDC9sGOLTULIHtdYMw52QtwD+oOB0gePcR9
uMpjwvNPylUoWNWY79Yp7lwC8lm1tmgRGVoxzHYWA48svGCb86ptSZmJk/tyXU7G
JHQd+fJpto+Um4B8kEhlIi0/ur1jOMBU2RHIkAErU1GQgZQ9eK5/8zraWYE1Cmop
zY76jij4MxJlo8Y954s5c4/18drbi5ewXhHTIkFlUDjZjxOo/oBrxV0+aoVBDMNp
RQYJCmffLKT9wJZtoKE3CqMom0jqkWUHnZhYU1yQxV3ht0bbABAoEP0e4P56edGd
/xf3RxF1wwYEpj6ihoNZiR1GtTsyn1Pl+xYuNoRUGxe8aq9D+J222ky4GgTxJm3r
p29TOiK4P0+mGKyoPAKASPkTznFN+Iqfn6XIU1dR1ssG73/ncicqPu6y7qFUwrpf
fbafJaakEZTbV8L2cb6ehDkOYpp8Hg4JzEt8TV18PHg/udx/IIMJi4naoOSHifqm
T0pJllCpzO5gei5BXFnzy8KDrC2OtVEpOK4smefE7mzesXHrOjzetq0u/ViUQlgi
49G6pTo+WN0TAaWMAafFzRLCGUtcAth4mAduhxERPagtyU2b48QsMyuodpH0p4/I
Aa/jWQYyT6iz8hJAoWKh7bt768GdEWFAtY03+q1mRAxyVyIoy0Y/D+yqvS5bD2r4
IBzm+kFDeRRNWEK76Jp973o4V9oMIeJFkWUyLeNraDaVFzZwzWyQQaMrcUTzbokb
minH/uMO20hT6TO1DcwJuFBPoFvlMAZmgaYlCf5N5oOQi+Abl1+3nAOkZlhdWcg9
VaTWlhicqSYMC4qqZLq/v1YBhutjTSV3r/oFda6MayUvON6wsmbbzkSwU/odtZSY
Pa+bgobw9Mb/tyxTg63dELpytmcAX2rwRC/uz/1uJsxT8YCgyWmS520REChkkFBA
5qMzgGeE/qpEJJKzLZT3NWohHHuOvOBLvcGPmeJdiK7yvDAfmhqvY1tkDmXOpXwo
UQuosmpxKP/YSMxgVveIuWWoowEvrEJcvKV5Ej2YUd4QQyLy+zkr+plnwe6r/n77
3417aWmKDZt1MvDVnDEuC+vcOMoZEeMajFp5RZ3qdiciNvEWe1p/lepbsaURxSuG
2KioPyv9e/u0TqvEIetO9WveK/lr1PoDQxkeYC+BBDaTqfi2q9vhFmO4lfmWIw2y
4IIDmZlMGtO1WdZi62dTeSAZBS1hcBXW2uNVc+Xhe1L9/rL2EzPwjHAMrywnPL9T
KFrMtrUoJf3DwH5Phy5MtO351Xr+vuKvNvaJXccCJ/FTinMP1jyNPLdpqfzHYTnA
oUQSoMgtONONdJ+baWu5PbdR2tL7Djw0Y+Z8PnMbA4VEV4/F8gWYVKYjBUx6j9Ud
3cyWGyVyfqs3Eege+sB1Davz1chxJjiQAXPjhh/FnFPnQkjEuyy2D8sQAYe4KQY1
N9ImuINrtiYu2Zy9sjzr6q673jBwWZIFUh842I+rAC7sLPbF/3zttSM3WMeGayoP
rxHxg32d6xa4xtzdSGX4fr9uSfOrv4a7Jxm51KiyEuO0fIvaiinAY/zePcB7wgUm
Iz4/ZfebYtHCyXbujcZa84lyitIHEuB4UoiR3vPfJYf91+FKz+S2Y7g74/d6CWx+
Yk8Af1yw4tgaJ0PVfV2fvdgbJDAdH+OheRTYcUTMUwBGclUdMx160Fen/ym9jxJh
Cq4gZKk0o5WozqYO2a6MwBtTRHq0Zoqt//i6mG0+57xw1W8UjofWFSrpp7kTq2Sy
1n2nZbhzbsR6wTeQgXae9FtBrPt6PRL+IWKlF1/d2vTODL8AUuQmfUWt0pSkLleD
cMm7LvU7t5+qbMoUkMhhajT+fcnlc2OOjZKf3AIbEVeJ5NU9wY1uOjCmyaVEi975
W7ypOck4LC8k318rrrBqk776Au66Q89/H8TuJJs3GAKnet/av1mpO34Qjfkv1lzK
d/al1tNB3O1he2CQBfQAl/I09ZVET6M7CJVQeXwjDDhgyT6pjOTlBHiTfFY3EkYL
fvpYfC69biw1tSSa0pKoNdhecF4w+Dj8Acbg3qCRN/iIG2rDaLS2Kuowp3j4Etk0
ukksPoD6pZqWlmKaXj1xU3+qDwKD9DUg2KvA6svv40LZkrIie/7VRmajcgJ9P5hI
n1EflJlUvdwokquj0ewPvQaA+6O+3ee8iQyxbHb7lQv2DiE2VtB12QTySOOzdUPb
ItUJS5s2pNhTCNA2w014eIelGftSXwoXn6o771vqvbr8V1fnmH6NwkHAh0NKgiC+
q4dBX2IvVPCDq8WBLfPrzOa5yzbzsFGcvQDWnbEHACp0P3mvpsufOzKJ8AOwXbJA
gt7UUZdMx/ELVSL700XPYCCNu8Q88TeAgCylRDTvhOmg6NCRXB/oKgyXkD+N90I3
ToY0Ke8KAThfbgI8Ru/UEoYN2jP0AfaKbMQuB56OPb6KE9g7wO5CRgtyj2K2uE7O
PMdnFbak6EK0UiyEbaeYUdUP0lCO4fTzOW2LC/rPLAvBpHnu0bxzWJ1CWvZG3/5z
Pqe+qvyOkNeOqauhim/BN48IjSNNedObRHTnmKjqJndIld4gR7vz2WXVwbV+DPCW
wtKr3+Z846BOzxstEjnBy4o4jZfj36IBxfusIEuW/PP29Pd6ZY79UfXq/pmzoSMa
JjBCfuLysnicrkirufyp1Yj4ILrkDKmAOM8idvcLzC4Zm2RF+yaniA7ms9mAAenz
BUqEoFm+C35KHJ2msbTvxMXuMprMwcD5/L1kTsScRw8yBpCHyel1vgb0xLNVY4mX
65KXdN+bdqNiXka1DtgAJ0CKCYp9GGZ6SB77AVZgxb5MzPw/cDRWDknppyYwaBdo
k8JdIZu/LFmafIgwG4I3zJ0fxWEGZY4n5Gz31nh5etCRWLEgjFQ2aXgvP5f9djhq
ks/R2FVVRYyRUlkOuY5Y3q9KEfSuF3zM0PdayxopYAWNZxrxZukxomy7RbRqBY0+
g8uyzURVy7X9TRAiK59AwE5ovurL0rlpPFKaHOiFr3RU25Nj9jrODv2tuy42TT9Z
MgaVdH6rbwXxkHuT+hCvs+YvPcvILIxwrb7NudVQGMbbSZX5gVlEnhUfu/smMWru
tEGVneMNwVKdIYcpjs/nAspQn8kmIlKzEAzsd4tiMppsrksfyzx4kyKODF9F0ZHd
d38RTzI5MqYb5Yt5/Vtt0mppVEoKJmoxKm9rQ9sR5SEmGdoOsIES3jpkrJgLDk5Z
XnZhdxeCYavRqAtNsfgy9lTAvEwf5NHjli5/+mCiBrkIUurukGKuuiWBmiOut8wv
4gqFhzMJAL+k2IDeXOpHSYbjwKtRoJUenjM0xSFXGYxoGvIzZytgxAlXbYjXYhXD
r3kNC9zsGLzzIfwxL+yTlY6+7gDQR4NjrJFEqNrHXC3TUpvyA2bGoTF8rub45obN
n89qjTHsiteTv96xZ92zXV7v78wwJ9xzQw8zwYjaNzeYFPkpFWVHoIfVJ1HLCxdU
GqdL5fwtt6W2uEbK5b5B3rKp70/QuLFCqYnjeTuHGpdUSAwl1P30KqTcqFAm6VIp
CDr31YROV7Fl/4XqZ8wy2+SwTTStD4Gxy1JDyzwvpB4O9QASzZmTYXLMF/uThIMk
Z6S2XMA1co5BFJCh+D48Bfl9DKFZDm0I3tAa/2a6AhbWsl73GxLjXV7aAs0KVf6e
MdmUEO707cUbZ4oJMlscHhJtGzQDeygH/0F+xNxDFOOLw16qaD5E4FyLGINjmHTP
F3/M168LWuhQk5x1bpDgMe0Cd01yRPhRLzlBPRoIWSzHJhw/ZGeBHZbXfxqGqUf4
6GTbJ3qT8R6us1Y7xDQcOSeC3yAmq2FQdbxM71fxAulS8gkSASLOBmOR7og76tZM
y4BOfPnENe4yM25146Dibiofh4aJpLZTEYjMUX8Qrjy3ujHZSjbfiycbB1GSCdvt
D6SvpoaY64cus2jQu4VgaYVdtihdUj9LoFoeGupV7kKsfx/OzWP1PA520SC250dx
T8uByPXspnP3kFFiyMYjkbSB7igrFxrB3qsC7/1e3Z0cUMTcqC+mAk9hQXGZqI5I
FKi3fbVH6A1DI8UBjlmwyuirF9jg7DZACd/rzqCxawdmKRV9tlUjTWUo7eEUCa05
l/S81crNqDv7YQyCBSfsTnPxUhydkMNm5xoKCVqdBEdaJs/IdfSt6T/T77tzrvC7
q96hN44zjwFOGdJaX7EfUaqkXv7Slcvp8HwFy4eKYNfLYdD9W0SrfQ4oUaGAxlTU
Gvj4JlMVmGaqvUpUfKuemFXOtiFgXerXYPksKZrMCHs1cccivr9MnkonoyB2GRiK
njpCtNdno+hkf0yx7zimUsuWmfXAf8tJ57r31gDmgEO8fYwpyz05de1HfA8Sqc/K
gcs9lHa2siIr2sqo8XNDGAFy99ggu/KeO8WwjvUIURqUTUR5fZ8LgEd7CJGOcq99
ZXzSFPCqPQZqjQC6SjCyxU0fSKk03BAa1KUEF0lv8UyaVW9ufW/YV84hPH5HfGZD
KwHLEFyLvScVnLvkqgLmpNWsXHSTBjwo94ot4je81FpjmfI+raqArrPOuZwZNnb7
B9p/sdTWJOas44A5CPJl3B7Il1JKo+iSQ6u5G/RrLPJ2qWO3+sRpXNK8JCIz7UFg
xhO1vEQBi8h3U0JR54v0RixVvsRGD70sbN/y/4HumilB0Cp5vL2p86ryuWTCRS86
6cV/4QEdNoO3lbaEICgXHisUZNYkVsT7tFuzx5QNIYrY2GLvAK1YucmDJwaeH9PE
R/5NfayKm51TiiHpwUzKuFjsFN0/LHbf5GWJpy9+HkoeKIdcRuRnYsA/02hivA/k
+QapWHftT+ieBJGxFG0G+UpoIxzvtWmRExQXvzbxLGNcfnEiJrGa2UYJJgZ2vwHp
ejvFsmpJwbHGmvtg6u5GQsmWtsqQbV4bGq0t4vz6tt1Z0awBp9MYEE8dHA6Yc0cB
i104+QoO3U/qGYFG/jRVIC5NDKYxhWco8Ym2iW3cT74GTUAHBSAHLiOAAlVGZWON
fbbq7zChlFD9eMa01B1oqrIcLH8i4wW/sywNUMlLM5+B4T3F7hf1lfNbv6dsKkUv
5WmcDyuEf3fbQUASAjoVEHGgUcBwGv0MHmgFP3Z1Codnyd2Z9F99iGy6bOTNTdYR
ILWm9JtTopdpzQx5Ly0PV0q149AwqEWuzqeWuSGHUDo+fp15uKj5sZl22sU3hbaL
G6vClAROdU/tFZOovzheWgXJXw8gYSrMqg84eGghw8Gp1DxovGA2cCzbIVnerN1l
TFWMxakYu9IwjAkB7h/KiUB2zj73CO5ARbOQQ2+YJVqbTE3sD2sJq0qM9fTauQt+
YlHKxvjaqCNq0ipO0iQj+77TzxTVFPT9GciHoSK3XLzkkWPoY8aJTsVvnO3Uj80G
hCto52paV4Op87bPWqh+1+JPgGcmgaoIRfyckbqcp6wNRrWOcIbVJsi42pjK1n84
lieKnsv1PYOOskgWoIMhhDCADhWGVhirb6LqFdxDGwpAjqQWTz5bLbVVzAZMhNQ0
UfPn9zioXsexkjb03b/WN+685Pl+FMYxpSETZek5HwyrOB5tV0a1H8RjiU0MPr7D
ketuVls4L02RtB83+Rd4OXEcs+/aJnitlmqN+pPZzmTYc/o2jUqOqeU1Ox8OjVeN
PKYR8Sr77c2ZEdxINkdCWnMbuNUPKTmMnVrQbItAD/VaqaaHw+k9r92cPiLtx04q
ZATPWCTb2mv75P6xzoep9pRwW1QARLS6AtNpdlo7MzqyCoxYLmnwGnd0gd59HM/s
G7rqJ6rOinJ+p4+IVQ+/04TPNCaSkcqolphG+WZuhRdJajWJ0OW13ldpomOK6Hqy
LoXDVkNAmCymj/fBKPP80YEuX3PM2KZvVyQbkjstnjkBek9PoNym2at8WjM+Hdkp
hkeDSbqEEf8hLrF6MdmvF4+gW6TbaO/bzelwoN6/1zb6fpWU32naVIyhkq7BTjrr
PkEE9efBq3rSyxqAjDMf6I3ZKBuapg/qy9EPfnM3dlaY9/AB5mfnegg8zgAAyJGn
Dhim+3C2Kz5eozVRuoMb23qgAjxjE363K69T49+EAttjFX/40wxprASqGsxUtk+K
38rFCU6vldZ4/wj9jxEe70eNbmvxuEFWaYUyfQM+vVbAznSKcOR+rRbuhHsmfwIc
Dhe5ZhWbIWpDBugII+HKjW0dTYs67tauWvdaTSgkqBKcGcWuowmlI7pGV3AEgggZ
NpcgJSb4uTruxYMj9uHq85TLgtV5DikaXRZSGHJ/QBlrhnFv9HFyV7JKRl4btYKL
9k5JMPBKL3l1NCVooyhLxo/kfvwEGSifQk2yk1rhtJ4UeB4ZP6lEDz92OE00TG0u
iGMxwqugxJkhYzJGc2KVZhleI2B71WNZ6V11huQ4O5JCd23/fcNTyrPyktb1I7hW
U+W7mYBZExUdfgBMt6ZYOH5767WS4ZiCtL52m8YORSWqS2DgTSHzJ3HMrPWa/UL+
ac0mfIow8Vs4el5Vdk3Y0jGQkw5KAqSltotNzgZrq6g4xg7bAgIg2TTHxNqmCEFI
T70Mi4NJzCfD77upWDCQZBIP+K1zYPNYI/bntOCT2fo2bNZ0LtdoDdyHkwNOPvsy
76p6HULvVmi39TjxBhOafoEAR8JJk7BUjVbKVGlabadLiuzAWXA1gyu81wipOJoh
yZiAYwia804XYeZhiFqsGgwu2QDRZTOutknJO27FTzDoOBstgD4UaeoUSeteoQf1
7HG50BWYmWZISg2SpXYKxAVyeizzWjgI32tMnE0+j/mA9pAkt9LunupKBdNmfmHh
v9a9x+sJ+GdjRmBObDggp0KouPB9nZw0wIHHDXlt53fUP1PSOSpiIoyzq/9NuIVT
TenZePnueci37BlKhHlufLtEFTmxbyizjN3OxUQ4EaEP5TimbObPH+DqZjBJjty2
LRe7C19vCLWhmiGB+BZutfAWsMYmeqOwL/IYHnoY1+fodAyT3QxlSS5pQgne2hTt
Qs6LxAVZie2oOCSUfdPPNIPfZBhSQ5Zq7eeR9b+EWyqq7lrVFE29WQwFebj9OlWW
lw0g4lsrI5t/0zN/MvxLehSwXtpfn3o0OOaV3fknyrZ/4ZKKWCj/wvb98jR54l6b
ecpBicj3IldSsFOLr+F1ZSzK55qyZPxEmd5Pue9VmAdA23qKvDm1st7lL2a760Lp
8ufSUTp/lqpuVE9dn1rdHekpMpG2f8Sk8x7+KRlSUomdlNGuHUPHKx0wVEm2MnXV
b3hM1sU3MN/u5G/ffRrV9Ee4PUml7zrn56JZ3W86FI6AEBxBH2M8LqU8WHKqwlbM
fQH41Rx/xO34ifU3eQSE9qpdPH8xHKrbS57KUxesLhwnyRGh218pLDV+vrLIDKp+
peEsCQGJCmmMRruvBBtEgm6OO8+zOGpd6z0/PIGFhxr7J7nGOGONIhclwrV/aqP/
qF9fDZ23/5X39zM10oTgEO/WDY3fcf43bKJ/vEqBA6nVNRudBM9omS3zvuejABz8
c42AEYVvMVa/tlrwyyaCx7PcuWieybj30OV8MmhLjS9Jm86nliI6HZSOPdhIzSa6
u+tsrEB7WlFPboeggvOf9eiZTbOtNzZB5usDUG2txTuuHTAmQ/D+O/G6NAn8Qjyo
adjq7tJlCjMn1t9VrBoJBfCxehskejhlmcMTsLyCh5XQOO0hwj8iyZ5c45lLOKFH
vgRlSRCn6zA4c9GnwiVU9XPWcQtntgoNXo3dF1ZPs50zlCyLgLhHoxrxOC3BJ4HG
9YKcGojbxC2aLCeB0WLzPaVLzi/BMo1Ibi6heiVhDxkUmgRjTjUsrXGCIANASwAh
1iPu0kCq8p9IIq9/h+49iYIbLI4uj/3SfBwiA4E1pSMrRuy5Cn3MZx0tLd2Mq+Gk
tZ2ZGWpz3PB+JvjbQ59QGqTfEstn/t082R5jZwfvOS9a1x+72X5U70ZwhHmgdPXH
6k8Y2EdwVlwGi2QYxp82x4vKxAt/9HRVUd2pFwAyNarR8nqBOwejRI3YKepiqlNo
daVN2FfVAU3JEc7mVOmuYlaDjEbPqP96jhUCuWESn41+FlE4Y9j+a2ajYJU3N/jZ
2XY1kKcTiWD43KKqShF8rqYLSNEA9AadXMb9QHSmGU8ti+eiYGoZZiJfzcNJ0T9K
qCWr7qwX9DkAlUjoJskJW7YLK2SV3O7N+YP7JDJp/HkzRaz26v3T0FKZcWycbnOk
ZTJ2u9O4Jonz4g3XkQuRn8opyXJIhbGdvBzwOz0TOLbC/92DKlhTdCS8yFXi9mZ4
Adl3Nm9b6ysqo9+3gLH/AtGlUFyk4HiO8isC0IbeyXhTFCdWyVkE8R63Mpaz+KHM
/6WC+V/951Atdh9WCT8w0uLC7szI+o2OZlT03hRHo8aVPS7zHpdb72SkiN6kD//t
aD63HJ5AcWgGMsUjxAvj0jTSMO4wY9GMwj4oygm8BH5Uo74Rvkx82ed44qgOE/4e
9oGCcuU3P+hHCfZhMsiQ0dD4aCEwqGz+oQfrCyGZhkG0js0pJvsDSteNtS/d3B3n
7Qgq6SyIWETMZ6N57l3BwO2ZeIGz8GOEDTspW8+96odcoRC8Md7EQSoZ3Qx99gGb
TQebPM1/ua5kFgk1WPXCzAH9kKZ/KMGvtYGgbTWl41TSxFmvftflhYeUFSdp/Lk9
Tq1JUablDPIJzsdcKZ8tMl4GlYiQfalCSRE65ENPDWav3IqTP6XyMhZBnvdcxIbi
7JBI2WbOcH0h/pB2SJY7qgAZuuEopYX4ar4xNKOdHyb+QfptnGjJ6AWwZ87wN22H
7opytZN8SgXBW8EvU6FF4AgjcRxYImrS9j+qU32fa4YWB6kuWbHqWqjrRtmiNBRu
HS7N0vQM9g//c6Zs1M44CAWbYRS4AUeVFnkVrdUUqkpVWKElfz7yEdNA/n7vLE2K
6OiHn+5Je40Tb9SmoK7xPBeuZDT7DT3gGEaYcvlrAvTJ6dpS5oYFYhQ5PXlIrsbV
4mZt6g3zED3LyJaOk5KN6SMNsQOLkBAHga3xXU92pyPtLLG5HZn8HsPXdxYk8tJC
duKpMYZ+J75X/0dVmbjm4H87v+TuDhS7vkzSRZLy21TSJ5dWhnaqYAZa6YsTRbJi
uPRlHErF1TGSiYJZiNCGE/GB8u9B4dZStZNtfHAChFpU45bPwbmEmi6xt6aEv0kp
31p9oUamg69JOEhHhSW7tO/cQnJ0wYPGjKx8uJNp/xyxj1nsZT0njpBwTooRoVG9
x9lCaKkcSiHEJciLte6UrCigdCfXTymlnPyxiBAq251UehKsTFPgtTheNvrkIiyX
5fdvOwfN8Np3JKeay4CwUaRqW7xqXBUsTCm4F5+VvfvuNYFU64sXC3qOKRKL0Sgb
jZYShUfKDbjPmDlxRP5cosDPtzXWxs7HH8rihA319jyop7x18lvNmVDYZhHy4Kj9
KhcSryiwWx5CWJ3bvEhCGFtF6jWtzth1SjWxtiFNqgv1BZCe/MG8TyT8E3lM6LxE
cYoLXMgWUBBCGrs3hP9pVxlMA5gl/REBHuE4HA+PgJKn5vHISZWpobg/21j596AL
6xxkOrl33BRqV0enCgCSWxT6RaJL0YTJ3ItD4st2K0dCEDXjazpCKxnH7mhJNHUc
rhMy2T6kkkYC59dHaMgkJyTCy9uFXkmXkPWlM3VTwXhdeo9oriHTFElW6e9YEkrL
e+hdvZaFooxTuI/HyQjasRWug0FPW/gWBD8WkAbxjuP64nRXr0kqmaX074qayl9a
lOtKkdS8lSNpy36r2vuGuw8yRBmMnlvp3FZYbTKlgEZe+Ucslggun76HgkvyF1wU
HUdx0DnS6SttuZg77Ha4Oqq26iJDX2RIJF3CbkzfjjmU89+6+nYTFAjc/GnQBx70
0ZSOCORjdp86EEZfYNiWmuTXlFi8ooYZSAymf6TPefbOO47/PWgVEGpuraNmxbXk
JNUACWLLp+bTueretp4Zyf/FmLVOq98cQSpZASE40rMSOE+EYdHjtRfdVxV6gFOl
BziLQTA0zh6JRiGSIp9hMBSqoeGXMNuidiIrSSSikNoLQTo0R1iwi54Wwrn1X6hC
mfi0nx1eOAN86TSc3v55o2qbmAhE1M+Y1bQw71bFFKfbNfgrq6MgxlRjFF/+yzxI
9+mI4FxAvtVNvsLSP5L7eqJ8EYkAJbM9zHKWuIi4Na3M92zlbvL4xLruAwMN7Gv3
BLXCemeItsbB5D1gnT5I/E8eCGoaapg0Ymin8uuyXK8i7A5qLwenOj7j/oz1zDkx
V1oyG7Gd4up8Br4jLmziIDMMeKA6Q8KoOIb6/mKyxphbr8RLd4dXtIc4NxUQMiDG
EiChkAg+tq/diDApmh5X1WNKLrjRrUTPz4NaXqOPKdserQ31RibPBnUjEdMgwqm1
jJOfMG5XMvtUBnlUutojNAi7gzCj+oGj2RpZYj4q/XnCzU7lBA+Yjb3ahv/QuJ9x
LGnEtIum7+8yRDf2wWohkHJH45PtkRc7SZa9nt429ZD5ulFMO0zv/Z/Gg8ommRVO
2NJUgqMg4Xa/IUOH6HH63qJhki1VN6f3fkAXOyvbCYJFrXgxp7dBjBJ3FYq+DSOk
9pTQBe4xC/wJFzL/USPVJ7Sliy3+TtpoCLGkzbWPZg+itoU3XTMvOP8P2Q13yWFi
gz/AJTw2G8Vs0w8KHOHoIqtHTt4qYeKm4AcPxqs1QaXr6yBijfUGrP5htor/S1n7
YwIrdL1iiq0rbmEOGUdrzLJuMTDRHpjHgO5sOHhHnp/i7rK2i8K4V/n87rThP+bD
31t5ULWFDUiELNPGO3OFcCIMAffuNntgn8IZYyx8wmCH4a1QR+n/cCfYRUyhEvsp
8iHEHtpaa4ICEOLZNBMl/1Z6TqvMEuF5tF1Y75YKiKYzqsvb7Y361T/f7JiqjDzH
aVzktOIzhd7/5fckdODCpniL4qV4zqDVT8wGrx1svcF9dlVfqitOocF/uiijYBvT
Uu2UbiTbPsnbAhsMZhTejGh4KhbsevA7uVrBIQZatMy9hHhUul4hh6mucPXNE2hk
ulySwbytaNvJumpTbDc41MEvv1JJZUvlGT2V2xNpxhMIDOLOPR8lT0mROcsb5LHB
0NGr4XbnEyYxYIEjyfglHXlmAw8GUsw8+/wjrp1pvsIcL5Pd+ORd7ePmIzHbnUl/
TF4EPnf1pe6ezGXwbUIqYdCRoKQlQJeS+9LT/fxatGLWyKYXd7eptcrOqwDJM54i
djPwkMcC7U5VgXvwSkpqheyd+EaNwiVIG5bgpN0vDDinieudIg/xI1QVouRAqqOf
qKPa+BPtaxtWBaT4zCjbRTVyWzN/WsnPJlWAgxN+MRjrXnA0Z4QSr2G0+h00/O2V
paGIAFKxwkI0J15boDXt0DC20zf+KV8Kb3tBWaB0aJmw/1zkJFqMgUCcRMjFa4a0
i1JNGcrl7aldME3POn0b3lNg3v1M+KPWIXzIrVKyvm4ZtqAZr0KqiunAoo0xpxYo
C8WG8x+8rSjXgebn+cipV/Q+0DsYH2TcYprRqk+z7ebG7oEBqkyAb1HjeIYKQiV3
POEt21r8Vr8fS4O8G7wkNCuAzAghxw9e1qOHkJwlpe1knA9X8aAxVx99BCUzaOzB
Gmwm/kSqbSe0dC4n0X3txar8AR/9+jbHRgI/IWTEJrLvNDRZdrotTeXmeWKBRihe
HEZ/pafh2F9ftiGKTBwmQ515YNWrOQW+u3wrwOE1NzKWWvplzwk0rPKS5MoMZh1I
ILoIPhj/dbZVGbVzsuj7yroC1W0B/EMLOT7CcacgHWRDFOnaZJyt5EdWg/1fPOPV
nMoU3DIp+QyZN74WekMGBAliwq/XeFMkdrgA+93+OVqy8V881YMN5XJQs7Z5zoOk
fV3AGXNP1z43EHcxgf310vmFXXsdrkg6be++vrSu8dCn8bH9dphKDd+JC6i6UfXx
k6uNSDSw0A32Z60Joz8Th33aHayw1D9R5gvJIi7FIrGWOAtFNi3CAPs+0WbQL+GB
30x/oHp6kiUYROqV599gHg5vd7llBtx6crRQa5TQDHYb6lrTvk0mkEiRbkOx9hFX
FzbiAGyGl2YVhyL8p/ohxs7xNi3Nv7zOpEppJ7/hrrN9jph4dXMd9UJkOo1e7UPn
VDpq8OLSrortpjo8moymSl9rR+Pr1RUJQk5LxYeejJHBm4VpUEBXBek+yZFufxi3
uGYP8peS2r9q/yR3jaUd36bEDSD/Dpr+QskdjoEtg1rXsqrhEiSmhtwNMuw8TMn1
XzdiWwAAT92w0MP+gQ/g0qN1WcApWSZLwE6QMpUVywsFu+5X00ftUHuHEQmynmg3
V6kh/cvLDnT06Zhaeuo7Cx2c4BLXItODAPle2A4MCuosgJJSvLtQ3GDnbwRGgDY4
EJmTs9Kwp9MmbJZs7/Swg2C+PVrmVdXwI39ASFDPKJl5sBaEsETrVWubUUsd5Oxg
zrZrRpMhnOyI4T8pmuZJ7XvOKkfkoOhnfnboJVmyi+WJGjFnSCTfz9a1VzKy5Hv/
4/UhL7JTJNxjTAVh5gr46L5BqXWkGCJBW/HGBhv6N0iAQVySdK8khFFchxmlu4Ix
zwINk9hlayed/M9hEM3s+osJrExHdOg3RlokzGet2QgAK3LjhEa32z4LdLmPnR8m
FYrMnpNl089iVKVhLQbbrVRDAYO4BXclkVGVZyL8KqvGC/GpoyCK7dQ+7fbjYkHX
Ez9mHzJDQxfLPrRGauM1euG4oryCh5bdqktXOzthFVsuJXolt4AS4JzAMpfeiyn8
l2/E+Ot0eL8gzeO2D0NJ8J1yleBt3l8jB+/bnIyDh7VXkzi52lb2jqXR9RNiSNGe
6ly3d0bdtfYci9SFtgFfiTB1MNn2GXe3X44mP8w3sUm753wOXORqRbtRvh+CT7ox
FDSCLup5Uj6Wz2PI3c42aJl08bZQEQ7BL2UND4hV3ZqqGasXi7guvYClfpB/FKqh
om1bZ4nxwjNqe0xyn0XdRG6UokuaXp3O8ITLY90P4zTQmYb4mNgVsC62g3XxuT4a
oD+Ow0J+XpvhpfEDoDg+/oNfimu6J3+TK89vGc0dr1BLmq8z0qYAf++IA3qUnl9e
gv0/GwUzAPvpA4o5BZsHCk8N31wb1cIJpABQWRxFKYNQmVA6sjwx5lBHk6K05pv8
ZoylWizrV8hWAnRoQa2JEtRSMN2hbt2benR/qwLlZvAo1FDGHA5J1gD1of1v9Oq0
wLO4GzwHi/sxpCjIqYsI/RfKBS22BfGVwe9mwG2r9JbhaSk/l7RnBy+aDqbivWGb
11r7cnzmqYX+UgAURJVDgsWq8/ON1dh/9p5FVarrtIo7DxQW52SIZ23SUeUfVTZo
cPKyrM5j1OMqyv3YBp0+ANSM0tdcTj0CaTYJhIQ43QLgesbVQtCYc8FtJzqB2F5Q
xivz9zvBQWnQg5/MZylRMQBLaipJzA5zKwPOeOXKV3DFQZa6k2VOqRP+p+oQdKdk
9RR68flA0iQCvuDtg7X9/uHBjnopQ5hKOHQAespX+KaW1uSSDH4rtQek5gDFrZQl
fL7agY5B6dNpb9Fu07xXJhiLHDQwLBzakgICtC99eMOCGOh8gJt8Xbog6ygf8L8a
2ZMBr7hMKql/8Ski4/KD2wO0RK1rWHsj06obiDginZtcNdnDMlmbwK1MqxIPziRM
+HcGXO5qy5Xp6cikeHAZCSsQP4JatveOxjjQXXXx2+Hb+LqlrCQInYGMCnn7Z6K6
0bpQIhNGgPBK+AEtNJVz+BRhoZY13XtEpSYWqI/hS210Thg3NI8b7ZKDXHbHboad
4UiNRC3UAPHBLlnF0a5jhcJY2u1ppT8W5Ale6v0Whuurs6ocBk/hH+u6j3xOOPKB
UygOF2PkH2DHBaIeEsp/NnHputjtEhlbh0tYiz25DO179L7OMxyw29T5b6eMToYB
NKG6lJlbfWChifRyjzYS4JL5TIAYx+orbX4sUk75/0x6pSihUtelHHNKKjh8fkgL
VMs2RsHYvEMkEz86/6EOS1e2rziJq8Ml1KnMMTnnBHw0nXeGu4R8NUFNgyKs5Wrh
hjHPe+lRWyVtt974GMdQcKUPiyPTnOr3FXmSm9ZOqMGRMVJIRmluDso81vf4r8Uz
sMapFyTxsa4J8aQgjATWVB6GBeokOP/8vbUtjTiFe1ecAP+I1MJOjq0wdTBNc5QK
1umqnoYTb6fTSkGQtuBmcq4CsGTUmOQKDAcnLt9XrUqObHIZfy4i44lnZa4TvQlZ
zt5yzSkf5Dbj7FBllGM0+yVPP9IPcSZIIQgddB1BUxQY2eWUXpmJyYHSpTYld9AO
Gg0wi+WQJQV2n0WjXPQqtyQmwsDmcFnrpMl97R7yp24eS8F2CiogOjr079nxPMxF
trxblKlDGUtjJ5SAbiQpnBHasD+l6+wrXZc5z8azyD9+EAAnvlW9Ft6BuHIG6ZS/
gusSvPa+vlx5vQURuiANFshsQtMhky2haCAGKZ/ZdEQ6NbsIs+dmD3c/i1xy4he0
4Ko4r01uy6YeiQTF37yCQm2WIWINDYvxDaQKGpejvxqU4olWejDQ23icshxPHJam
OrEchjk0jGLKqHCGHdqc5qgQqnBLJJqwzwBt7Hpxfy/z311cmy/1Dkc4/w5B5anf
oQ4rHuplsqJxKDraoUBsmn400xvApeDhlf9Rc/71u+yFai0j+SNqG2OwW8DISL3J
SGQ3xPksc5x7pbQOfAuw/4azjC8E+XExe0lrUoe4v+dtMILlAXhvYad7nVmAx+Yb
D1c1x/AiF0kksxuTkwLO/Sbiqn1Sqagw7r9TrLiFWCimiT7znx+4xb9/PkKLmfYQ
T4TmXE4ngnqhc2GH+RSMqtNiagYfWQmBSgpSonRI7q1SKzxyMEk4snDb+IJgn3/A
r2l8qTTjq/Gvp/b4cyzHDDeVG7fqUv3a8alL8FnX7wZJoTkU+pJqDCzqcmiRq0X/
wP9BF9K+SpPmUeilsJVVsS3idIL87tFQgtmL25cNmtB4bwtkf1JZfEobdb3W3uBZ
6bh5F3EXuq5bXo2Rcc57N6I+Cnz0REgCtyJLypU/cKjI59Yz4Gm4PfDcwOlKCEW9
5nv1Gw5lDjnHwu11V4UXjen/cwOVCVNzP6rAgxv9e+NiaZwmNCRUFtqpnk3qbAUr
JS/Lz/c1bhSUgNmsnkyjr8Mdu5HEbJ5/43K3xpfbkZseFR3OsU8Fg4aB7drhsrSX
ZBA6FC3rcA3ZuoN9FZhbc6OIZYiwe9bfCUuLPH2ef7ImPN3wAm4Ap/51318WDvYJ
KXtrNEV39+w4WwVKBqbH0a8iH7OSYC2ixrpKakhjCED3iqXPfeDdjyxlJdHiCovm
677u1mtusKOWEhP2wGEqgC6r/kQzOwMNdNgurZghQnxcecw/qira32Y+PDqGlISr
Ox+3KnyTcGJJ+OxTaZybhrSsD9FEmUTkpAxGgnobKFrORliWn8bQAXVNkfX3f661
J9LVuzmy2YDni8kjd3YqO3zOM3qGX6tcgdQeN1bk8gPDslCgvYlLKINEVMSiYjtc
7qLRdOSZYEpD5XoOBaRFhVfBVzmwDbHZHTfMFaYCwT0mqes4VJW1luISZFNJseWR
xSo9rXvp1zqzXM/XNh+G5OcoYhu4UHXA6p2kjNCDNwsGhwLeay5BvJprP+JGGxvZ
JvKP8GuZruuCYjwlgcLbrauuPK/WPKJfDdoU0+S7IrsNikXsRR8YUpyGiHQBnqkm
UiPbJSIROuJ8SMhH1UoyCffh7mPINdjf4a1F7JmKyJYApqdpbtaxfuxCvqx1Z7Fv
recdC7jtTpOH2PSN6yrWsv/OAdBzJ2la9knC2nOzk/otKb/exh7rIDBvVS9BKXds
KjvLVt69qi4mVVk5brsU+zH4zuCHPBjhTQzeeAX3kEmGOfnhYGDgn0v1JwJZTF8a
+7yV6w8GZweJPUXjiMROfMZok8Jcoq65LB+xV2NNwaPw9Iu3heggf2eQgXMGu0hx
RGXK8Ic679uROJErwLqjEa2P83KgT/AbVmaLk3N4mXT03P1j91P2LFByDdjATZTd
GRSwU1Y4WR4h8LefPPpIjZLK4l3gDlmavP/ImztUHKTQL93pBhKer+f6EjQvkw9n
yWRwWK4I+S60Th6GiM5gX8WPpv6p3J/5TItaw8rghODxjgnBEYoGwGlLSlNi/MyZ
W3ntQJd+FsbWoUicy+YLaa2gTzrrC31r3c/Z9fhkikJ7QtOfq1u/FTSqitJhHgn6
GZomD+xXCcU/0K3DK5sLHSca5faUNKsfl0IKlTsMaNjXJA9dI/rzmMpZf11F2qI3
o7GpD9cErd8kA5I9teFR8jsqq/KEY58sf+B8gvzgEP9YJhXmrHDrvKXq6ElbNKPe
0BMAfHQpbLWxJevnkywFYOdXJWyTMWsbcjj5k4pJlDHEXmAj8lsi4d4bBcXBgyz9
f5JTf/Vj8MuqAz6uh9xG+PL7y7PC3GPQg+dFWbeS/EZyfVkipCyJLG2ZMzawVYC5
mg4xGR5qHDq3DCReDrE6Ed9OjlHuQvwLEYadw/wXRtXz2irfYL5/T2zE8SXupL/g
Wp4a2FJDHhCAPMgTn3xn8p0vhDTonnVnPDovdpuG7bWZ7Z8ijl4gIxZjnGwC9Ne1
j01u7ab/vN00NemSvA26TiEWpZn3AH2fVI6h5h12sNdO5FdpD9IYHpJAW9Fo2pqQ
xQB0rARWc8gOp0+k9PapdQqBRw/M9EdXYjS98g5DDU+S10NW417TH3Ore475a55B
DjjKnZYqHcQ+uLEEsxFQjw1CBxn8WNsfGXm1v6/jwXN0ITxKHFKkyU9ZN7zApHjC
7UBDM2VUefu+/DiOFGOIQfNtOvom18BZIL8MdT9m9onOLBobIJ9q9VsbSTRpih3C
WV3Pnll+4o6lSdU3gK5JP7c1LezJy9SZNFTTl2Mcu/weguV/+xGRTJNTSz3gkPrb
lyv6+i4Oq9ZybyQ17JiSkalRQV2nDv0C6zrIsx4iUrRBn2iMpWo9iLBAw8YnKxtk
3j3FisPkCo1dBxKPc+IPUbPBabmFr5D8hNbDLovrBjhQfof5atAUyE1RHzaqlWha
AsoCjb17EzE17qd6ddG+0n0+oSbvSsy18dcScJGXA7zzTKE5ubiBCPVpgM0/CyRX
ZrMekaBqogEMyCXUfNBuwyKT6k/n/DbImwSfCVmZoNju+GcKKdctXxTE5p20LDJt
Gh5e50kUAEkMT3ly5zqMmFrUE6/Y9enZWzGzI1aocwL2tnMBGacvDIuWLhOB/aI0
/VhPgDwlRQ8XmfryxYauP01dZ0OiNDPmvGj9cZn74GyHftyfoxGw/1jvhYYwZy6c
SaKxOqgn21WZG8xLqYQXUzhu90lK0oSJ15LvV8taHVHUmxysnHyzHOPbjJGOh6yt
ndpmHcRRp8bIwjSWvBNDDfdYoTPXEhQ7LlorkdBS+C6HvWrE+Xm/icD1Eq/h77tc
DXru37Rmk8ysvrR8QirwbO22vJWOQunXUY5Fo9IVmKjCMi6UVBmu3pu0+AA6HQaF
cDAIB2rvEuLWojX5h5Uo0gy6o8l3FxP7A9z/8qv+AAe8cXCMvYj7qGltwWfujD93
QPEVoXLkXU2KAsl5Gb7AVIJSXeMoiTuAJ+DrKWBjuwUgLtsRoQyQyAoKgnxCeGNo
+FBpSWWgBLkpfIWsxvXAxJ3bftsNs1GNd9b3yjd11SoVfN7EPcMHdxEKOS9UeAvs
57dmxM/V/bHe1in4c9wEpIzmXJco+X3XvqZtpsmNsaowcg10gVszkRs3or9MoCF7
qM75oStQCC6mbZfrVc+niVl6B5IgYXEXZRnUGsYtTcBCWkUozgNm7biJmioEwGo8
IYyG1XlK1Psuhvs90A53CzZkc/CVjrHUDWJh7N/WdiW6OxkuLoc6yDE2eT3ai1wT
O3ft2TZz1Yen6nDTEH2qO7D7yBMm883Zynply0ppR6U1Qx8/Tbk/ebemxFeRySxz
auqfAOoPg9cTtDxm1m7w1Ek98OasKoLVVisjvhqSO9iGyLHT/yccTJdV1/uNZ1C1
b48q+v9NMMQaGDkJ/2+ZnaPmBCJalELvHAlWxIk3jr2CP6tAP1mRl24IrdNwcnUK
Z267uspKESQnL4sKrbhBcL7x4/CDqq3qByyFAjmT/SPyWOMVwYlJu7KdLQ41eXTR
bTjaAtd801qMB8bbho40knvLxLryb/lJIM+oMgMP5IK0bKvAeNtS40B7fINEc5JW
3izMcBHj+QswM6YeCgD17+V7nv6+vF1+RTowTx6wBPBbgpbP+UmM43oWJD0mYj+e
fcVnI8i5pnNpxn+t9vCxha+m5AVv26hfQ3uSNIx62yQRPhTNtj3GNOdeqFPRDypa
+4ewPZGq0gqUHeiAYdnb6c8mlGR63dnbjuRElQM8kwpC912G/8NyFcyitpHM4H68
sTmZAZ+IiNpdBFuQyicsNcWRZZrx6Va7Go3i2GM9okfY3VqOikjqbsSulKHS6NiD
crPfSmgykJ/6EwUXG0/i07y16V/dHGzX7RFuKHldLarcE49ecUgyBYi3Mxv4ADUm
Bryc+DDxHJvBsHPDjJ1a2oeK8LqrMQsULywc1OJTSFWLpDrkNh7wDripa8Lsodo8
0r7+4r81Q2QeVcx5gyX2LctNAs2RIVlo6AqB0c5Jv2Lxd8eszclo9ZlxNLdxO0gU
6CLFthEzOx7n52bA8t9tykB9Zzmw532aMIpK+ZJefQBz0/ouculSUMKyzBIOq/fN
hrfeIW9Z1VMQcOdioG4I3xyDeKjQZqPxbQ9HqAIG/+zYKiS2vKWwhN5R3WSzqUs/
hNN6zNUIVVnUG8FhtwL14ABr4vtZi7Les2iOFNqhYJM1Cb7Km9MplnXF/z/H5WMt
HY+X2u/uG3d9473OF0XlL6zWdvg7iwAKnnKxLyzm0C/P04VWoLUur4zVynAmBCMe
hx5fFngf2IPS2DvMdChd7DXqVB+SYYvwxL09M0m9+2tKhNGIsE81UWZSuX1VUVid
h1VsslThyHvE3DcB7sB3y3RQythFylAr/q9FqT5UkzojnaMYLpS8VvElDyu3gKwY
RRShmAo5Un+SlsoiC1XMHo0SgKix5QNmArsFQ9fS19qq00WjtJPRGSMtwai67DHI
a0PBdNT81ZAYEMWKN5JeVId098NU1+sf9O+NtlDBwv++OqcFDizb7g8AL/z2OWFm
cV3QXepPNwbdR4HTHjFJv0npOA4zpAfMwq54yiWvg6SF04R37OCmm+Il53A17Fy/
H3vnzf7okbiXXv9YI/XxlyHUVqwNcj17a6fglvWL3byzmTqhYRaeGMN1gs7yOure
6xqz6Dr1oFuWaMa3iwBjcqsGQoR6V5j0z6nB+tBi8dnMTdhRiKeF2H8P7rFMlWbw
QNXKyCR111SsensXuE2heLmfPBRGwI9LLk2LnltKABi27cgBuLAJhQpNN8dDy9Ye
SlbhKkfFNMBI3a0nIaIRCUDOWyBMLTyVWZ5ROpZoyfHSdlpYoWWzss1XOLZfXH5R
JCrzF0pw2udzjjEHGqi98pypqwBuIEZ7NwXgM9+3EdDDSr7P4opYK8YaUqa03az5
Xx4Udx38sHr6OCLtyDPgzvu1LL3r6LJ94TxVYhVSrMFhXz2gdAAyqSLxK7OMZRCA
gKvo038zZDDbDgZYWE882jQI5LGKa03EBK3dELhd39kOsgfyWQnOj/i5FatWMhVu
oO50SHG7snpf832XiUqtYcbyLEZK5MGLdg978fPPAZldnfev66YX/jYj8UQOI0QO
2S4JOF3ejnP7qVA8lE1NbcMbflRasc34PgwaHRVsf4TVwjHnMswqWCweCmNa7M35
w6LQRcu64R5MRiKgpgJsrdqNXiy8AEsMW4WGhAoaBM34BdQ3Na6i2qBGBMGJ97av
YxL0/XEw7wI4N5t5AybSwN96f6U+hezXQ6i/Fn6NH0ZvaJF8UIEFV+k7v4cEXeBN
C3uKstbvjs9NrvvV7ERWEW4ox87ciSIwEVoe0gZyWCV0Q/fHBvqlxLDYTqjg0MSG
q6PGwqeY86km+s1YEgQxOscKsq/9271VBw34SdRtZrykLy/cVKCZ7C5oN2aIpTFX
dAiMflqHB4Q4Apnmu2iTiHF/6nngC9tdDMUQT1E1frCabbrMZIfpebwSWkNcH+zt
RP8bhcZ7YiG8PKlL5N2y6yVPV9z+OV2C2pBQwIYhJSwP3YRsxl2O4H2uSAxfkd1o
pII0h4xwZE/mVXad1oJJwo4b2yLmQjuB2xBwbwLhwuItY8UFH+vSCmPqbhAEL5Ef
gtbkHfUO29qda5z8HkjDCGh35RlRUI701tD9V271eBwSmxaSWrxgKPckh4GzCjEt
6St4UvkH20SWSp8dhnfsUNuquuNra2vhyzuk4qn50s4fWTFyPkYdvtS34H4thv57
kY3tfXkWwzzTLu7IjMQH3f00zX9+7MdOc60HdrNIR7J6g63M7V0mUH29xk51uH71
rWGIDIbszMoNL1m6dxBTptE6sLIuUGX6bPFZrXtJ9+IOod9ufrsAjYZ2ZVvotKqz
Nf+D6cagN6Ke5RV3hrYLbdYJhilav0Lc6Flw3U6jjK/OVic77QyDMZjbraVQEUCE
SJPOTJ7jpgifwAY7LxCbYpp79JNOsF9pMxNswN5FDYNNwxSBjZ3Hh8gBAIjsZUxo
X1YUbf/MKB2I7FQf4h0bqDlIFdXmfjSk+Aoi+mtx8q1IJ+sbCKW1moF1iUCx0ikf
6nj/rxG3gShQZmiZ1VOpemDoXCBgUlS2HxE9ZV0ryD5TDmG1oXxOoP1h2omHhhTO
wHs+gI6VzogWs1hl/q2W7lqtfRglk+TgmsRiUSr28Dc0vGcB0PMW0LLjBWOpcIc/
owb1dpcUyB352mG9ci2GBZwe8oafjAHMJgfHWITMdHdbmrZjdqhwJPiZ0lBatR3m
oWCAygHTLTIZbtNUqoUlggfdLbaCwCb7QuoRICWvsSY=
`pragma protect end_protected

`endif // GUARD_SVT_AXI_CACHE_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
O5QPwCs1GTNUKkltg2vk7WpSTB83H87/H1dnXUFqsSW5nHJheH6ogo+vz9oSvhly
/pYhDI5Qqyl3yOSJHeTuGH38Yu4Z42toxAxy5Y9HrgxxG+kIj5J9D08FJL0JIMEl
mMfXvXPkwn1l3slVRXWlV3G9W1ZFV0lqTKtOObXS6Y8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 104682    )
XO3EDXrjTukVhVhEXa/raAUGLx7oKW8fwPJg6zNJFIJ/p79OHPcbeCjSCa8u7xeF
TPQH+QjadzDGR74/PkzSSWr5VqZPVUL7pyHbYnBDZIk+JS5CkDzEKXeKhgoIYce3
`pragma protect end_protected
