

`ifndef GUARD_SVT_AXI_BASE_MASTER_COMMON_SV
`define GUARD_SVT_AXI_BASE_MASTER_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
 
`include "svt_axi_defines.svi"

// Note:
// Throughout this file, the term 'driver' is used to refer to the active
// component on this port.  For UVM this object is extended from uvm_driver.
// For VMM this object is extended from vmm_xactor.

//vcs_lic_vip_protect
  `protected
X1RNWaR\&_SUP6XS(aNUbECaa6FJJB)<RYP<aaRWEXO;RWQdX(PK,(/d7OgH]:Dd
5SA61(._fa)KV6:9-gF.Sfa[GZXaS+.N^F07a^D9R2,#(dCI&39S8Z#cP<0U56#I
\\=Z?2E00caY:0FW(&=T#4AAG?<UDU1.1a+L+6,V6_W2[:c1H^fZ9#\@:_J8RX8<
,V-LdNgBRR,>W06=;>K:T0?7VbDA._\:7+&@<TN/TQ=aT6[)7MQ5[>4JbJB[<#F]
dB_RcUBR5/bW>d5(FN+;79Df(g59cBO+1f\+c5V&2Rg-&#4gAaTEGHXOUC(K;F:[
-BE0HQc^JQ5.4?NHVc)/aK[OQSeOZ@#>R9)OTaR<S&M;#LI/L]QFWS:Ja9/2bR,=
?+0COc46ZEEOCcaGW>Z:#P99+#9IJ:TFC0:AT&K=,G\>J\MGJGgY_-6<@7^=7+--
9Z=X5WMd]FCOBYA2be:_E\TFOV:+KU=3NeP#J^1TW-fV\_\98-G_NZTU;[9Q/VG#
-&20=[6g93AC_NT&&^U&8b8O-)#PHQ#;\;,>5ANcS;.6eXTL-5^L8<=[E.6[AG8B
Rf3?5)O/Z:_8FN@c)+?HF6(FZ]9T\VVG(Wdb.bX0_ec#FUA(YQ.8N7\BGf4J7+Nc
C.C\/0<YTgQ5X8[)1.L__Q^;+F__[9a?dO0F2I]L\1aRCDO00SSB[IgP?Q/c=P)>
V+efgP3)?g-3[fL-T<dWICRYVE?0bfYWT@R4BW:689I_fUfVUDO6HG9RUbUPY46C
.1=.-LY=#<,ZG6&:b9-,-bZL0OaRKEP/#S,<\&&3HX9X&MAI[bLV#.DTB\A=WWNT
YeG.I==TS2DFUT+-.P^47[73=F3EfUc;(.#a-?Y;;bX\SdU3MUa\A[SA[&G5Z(bB
4AMXR6G=-aQIRV-/W)\1=X;>WALA44WMbID44+A8G@TF;FP01,[M:b8(eC;ddP9+
6bM<J\682U6_+<ICBaA80@M]bWJe.ZB)MAEJfbIV.C#323IRDa?>QAfWO,dSAT9=
F41UgDf830PIDa-FP^;:R_dG,)/3Q;OX#O02H3Q0<G#c8#K2UXA=RdI+_T]0F&fD
ZP=#6YNK;9A^+NMc=3A?Qd/5N2CB/NOa5XV#0V&#\RY8C>P#JD6d3b_D/K:<788W
+N+:UfZC;?e:G2##D#//]Zb(-Q?G@SNQ3gL?)#PPE75,DbL;1AD#(\NV]KHI1S5J
IdT=V=;28SN7:XTE)C9N<NH:aFD4CW8(PZ8g+3GLS:8>>PU__f)e/c8X?A/P_@UP
G3<NY42976_Ad8Sgd\G<DFD)7b4.QA>/02#^\0SWN+C>S-Y4DMQBAHb99bDO\Ug?
adQI6?;PO]bILX-H>W6Q)H^27A[Y,57BHdSE8/)N=9Q)(,<LdN^HQVUO/7@PF->:
+\Pe&G=QF^H9(>f?1YXU#,/91\PR97\TQ)2OJdDNCQB=MaE^bL:Z/40\MEV+F_XS
V;c5UABCEFHUFF^?,01<1<IE#RB0#WK&e@2=WR/7gUeQS5;a\^<^#5g\&DQOJ-=[
e[f3KWB?6<-NK3=-dMe=3Xg981RI=,f4H2gCVN_d9e[?03ZVdKbK4D\b(7H7HGYX
f>OXO8H)eb3QM^4=8RK5F&OO]48-Q:4/Z4&TIFfURBd55[L&,^-8MFUQ84gJM;KK
@6^5aPSVb_ScK3H>J@VAK^;cN[a.b=F?V1OOQNLXAJHR9P2XD>DTRBAY6e-V>14J
&_bbI+.=:C#9e58\]\5MS9cB;1&<+\gC/JK^8L>g^da+59>fb#3F7+F=GWFPBEGN
LA?^0#;[\.9FQ#A+#S>g:9c</[ZVcdK2GYN0He97B5S3+7Wac_a@WbM3WD?+B57<
DfeXPUb_7F6QF?[HW/Vb:FQg4Z)PDOI(CHZA+2B55\,S/UVSNU+Z1NgAC8>F<4:4
1CRe(+>?M7Cf3SR:0:_RcQfU?H.H_<c,OZ7,Q>S#J7>_(>N@=J:KBNK+R9fd^EG]
V._5^&gL/7@F_R_8\N>d/9bb=>M];e&35?0,22;BWA;APK4W[VF@@^AR>97;53BI
E+VbT=]+DG(/a5>:W8[Sf?4d+R9e#;[aUS7?]35YR(=U2b/BJ2.A6.ZL8T[22c50
QCb_K:G2./(,R\_\cMd\H1>N>EG&g72TO3=T2D:b4;([^>a5R_2K+T1P[Yg)J4Kb
)g_>VEMeR9V8SV1Qb6.VHRQ5CRbNEC@(Z?(^Q08@SYE&5ISZX,a).NVb&DHUDBR,
4B/fHgSBQMH1,_X1,A.CJ,(WHQT?XT>[abM;OS?EQGJJUFgV(SJBAPfE.Ebc+1E[
SQOE:c8XC&4O7BV;3(F#X_(8X&ZP?4X</IKVSAU^IQBeO<f6G&-AeR;&A-1[38,G
T8GU@UVS+.[V.9N3a20NX5F@)-T[Wa]d9a1^aZMR)b[f:)\4/&:f8-^0OK/2J,Cg
@DZ267E(OK7VH4W_gb1<H](IB(-c\+LfKE[YaUM=?JKMYMLE9BM&F@HAO6;(Vc/M
d?e:M7](DW:gQ<P55I#FSXC.;T/;W(D.45RPCK67cgY)ce#38;MN_(E?Lb3,X=D3
\+1+[,Ud)^b[GAL)LfH[aeS@][Tg^IM=1d_\<MWSS+.[OFR1UC\5WA4D:=UQ(F=+
_gDJO[c:5BA2Z&C(-9+4D)[>Z:AUB:+A)FR;67125fOAEV,#&fdM-_4_Wfc8O\80
K53g?d+cJ/CKb/5Y@aKQUE3.g0<)Ma(IJgI)_B/#U;G@6V3-DQIeHR7gD2&d34JC
:/T\09COPFAYcYdLCGUc)7/^A)F=aBRabg:0)L+WFg8VU4\WaDBZV6EMafQ4F?fb
SQ/DV(C>2>@1/?/1cR<9?RM7FYIS;P&1;YFS?;1,/#<]Z94\Y&?D)KS/S<#:0BJS
#01H2@&AXc]6)JS_D<eN/49a]HA2A+Q-e::(1(>^=YL4[A_//MFEFX6Q:M^Yf,CL
/eSWeJ&,5533<@SQJ@Md/;4JT0LG>fPD-<JUST&@a1X-9&M<W@U8bB1)KMEAb65G
G2:HC:=\5G6ASJ@Y&7BWa&DQOP:4SbND.3+?0GCR._<AcfPPaTBW)Y)@L@^F;[M/
cg7EebVQg;7_H<.1f)bb^IN,=Bee&95Be&Z[@g/^2Z\4K0_P,S;JIU97W:J5<W_M
a3Qc:ed]15[]=b1D&eGA9DA[L[)dX;,,gaa^JX@DeEL(X#@,A3<Q#Zg14H2DU.[T
RbY9H(5@QW[ag]KfUeR-:.6AfFV.4e9PF(XWLG::@;5/\Y8;,K=-<L\O8;,[@4BL
+L3M>]ZB@VMLX@RbTZ5fRV5\7G/fSRcKCgHMeI3(V3ReWJC&#Ag\:)^8\.S;VfK2
(K1.ceC5U^.CDCQT\Z:e+aI+dV^2NBPUYfU#,6TJJ2I74\](T(;NO(666UMJ](JH
66R_L#N65R.G/+KDG.QeTEXAXKdDdGVB]D@LE/5ZIfKG=)U7SZga5b3,BN8=H>D[
:O+Va7V01e\HNIG/fEPK</PGH+GDMY@TGYFLeL(=[3gRMNCdG^e)+NM_7M)@030>
^b>5T-IX:YVdE6@P?204^V4Nc6GDSS^@EJ/3_2@+?1cVY[QeZ8Ug]N3>X/R:Ide2
PGL\TLNb_C^EVJRc9J;WGL5<R2]=d4Y-+B1X7.C=_g?EI1]F4[[@^M^N+NDMHP?a
e?3Q68Db;RZVGG<gK\I_g9&0RQ?7W=O5UY_Z.IOEcg44Y=4R)_5E:P5&b=CZ#JP1
7+-Qg[O5_,CJ<gT=G9TMQ<BaT:8a?^RSe+:82,:OPNOPcY\KeXZ0e-X17#/4U8PW
<1AV2^>RW9Rcd^(BR>+5GbIJ=.O(dSYJ?Q.Vf?fc7J=M]U-AKD)_IaY\Z(Z]BW>/
E(a2ERS7NKOGNU+-KFZUg7[@KS#c8)3XW^=^M]OUB:[&Mb93ICU1CD4<e,3:V;#/
a[YKeg2EGQJ+OA@SGY-LUE1M0W8W67@fe&P_12X1?M3FKfca.c2BGPK;b,;=^1b9
YHY^9V>)(T5:7a_;[CY7)0=T49R;?\4FLeSUd@R^;[K&J]aIH:d2F8Af6&&R1dFK
Y7>XbD)S6Tfd^Z+0b/ce>_NH1-&>J40.Z4T\20X)OYc..95Z[PG8DB:)5I@6EZSR
[.:fX<V)F6>DTGb=X2DSMaI.@g(<@6.F+PdQb1Dc8&75<fg,YaE^37P6ZMU6).D?
X#P(LZ?Ug>:5[<C;G\VW]BXZe#P3??,PH@.4GfQ3&;3;.RA(IHGgY?Z3OU)P#]IF
:3>UPG:J[4A4SccMKa]F/=H_8ZeHOTZ(_;:3UPNUW[CR.0F77>(6KN@+ILLQZS]\
+8VDfcWK;&1Y/Ya(C,OeF2>CCaX<<U8_:6ZV>;N1S8(=<W&)(L9-<U/^O>)^5B#2
dXQDLZba1#TG(K+@CZHD9;SV@L/(FU^cB4K[Y;O^9?fJRBW([R;=#EZF/d[Og6B4
1QC:\JH]>EQYDe_HIX7Z:d2&)OgZK+;YAg#<\5Y.^GKOIKe+7LNN=]9HC-9e485&
(#I_JWBO@?\e>NA9e,)0:[?PA>J.+YM&I[\1B.:9A-\;0Y&?S><G7-?0\\c?Sg^f
L;WI.L.[,)_I#aF8;)7?CWUXN+PJ9dGDP\ebUX@d<2>e&fbJ:7E-C_e73bH9.cKN
JT2)^N\DDJ0E)OaYbD_W_5G:UE2@:.][QaJ)-JB/C1N;/.4O?):_1;=[Rg&e(RdP
(=ZOfN/Lc;9[-Qg3-NYfg\b]Xc-[)E^>::M_8C;5<.WYQ/;@)X>]@CHP+#:_VU-\
EV#Wa60MT[LUe:MBId+_1RFeY3gDLITg_:?HYRLFHO;<?IQaMe+#4>,^3O..NK0\
L:(JVY:@Y.8T=+QS9.RN\<1YK\SGb9NR]BMZX<L7@8@06?EK7&K^cLeLVFLd.\-[
L;DNA=\\=L:N/A,W)@,c&?KRSgd##f_X==IaX/c^ab(]T>QWBW5Xg4,UU]H&FAQd
Cac?QM6&#,CdbXP1LU_Df_0.V:Nb6Y/J&d[4HQ]&8W=+aTOcb7H\Z<6gD;;0F>ZI
XQ(=fQK)<O:XB(2\IeG-10,:Ma_09Q^J(\I/#=2>E6]MDVBD8^7\6(1W1M,KRYQ<
9dFaTe9dA8IH?fGV1c2bZ+[T=J9TDNC6Lb9USTJ^B3)438)I[8fE7S0P?T7Q<4YU
49<a?=BH2MCdNMQYOa]4A1<T&\LM#O<W>YP(=R->M<)NI6f?^g.#HAcI5J2fL<@S
K##9-b8BU\]C]R1FZL#06J31KS9Q4^QAXXZ7PCSL:GSG;N580eKQgO+:LcXg&e^V
#=W]9U9@R#^d&Gg_I=AI8a[\SbPG=-J;JE_#X,25EBPQ?1gX9<gFTQIa7O&A<-cf
U86+-T)7Wa9VU&VI;>@HZdK],f:T:^1H=.48OK#-_R,4OIgK=c.6SV=/eXSB(Q1,
:]Vc@GHa2/V:@Ua)JB#EE<3^7OQ-F^]=WK5O/Y,cJd>I>gFC6G\(;,>a#ga:,;#_
DF[SCVF.67f#^7e&0Sb-eIeHQ0=^9VVJ??F]<4#=BT<[7]B;>b>Be2K2ef+8YYJ1
ZN^E]4^\8(^=&4/J_FOK_,S5KaUM5L7>QQ3[WU,[c3F;Q^)e\0>7453TcN:R]WYD
A7GK+3S=MNE.>D0,&4b;LC0N50PYLcO5RANKZd9,0NELI(@A0<2)0>TB-5>X\g^(
9\\[#9dHKU4fgY\C#gLX<R7Eb&H_O-HF?W)B(TI9I/.2ZQc_;LEV2D\LfC>@F]BQ
N,8/FX<^M04=/2VOGC,KQOB:ZBKRDN]8_LXBd3Gd\&g@8#GWE>@]W0BP)NKIf(U6
6AZ6g#ADC.[^:\?WSK@47VTY5./2;cM]>5RX.2HRZ2:QTgY1JceZ3X/ebbI/]@0;
WX1D+._L@bJb^N79f3<PO.#T&.NH)>1.8[VHK24fNS#a[H,UXW,RN;\0<GY:R:4,
HP=X@WDIC-^[S^=Y44T1F5;Y>HC5Ibb8e3Db.?=.(/GFPZ:Q,T>:;@,#N=LbJ05,
[1aP;ZMWS&M&=<-fRG,#2d7AKHUeYEH^BAY(=0f+-c)X8DKGQ9c@Q[P&9&LV_VVV
1(D(5@C2/+bN55;9_JaDVE>_PMc];0C\eb-H7XB\F3;&P+gHf:ZF@1fa2TE.:HP?
0SM=^X-36gBF/1+/9Z+[9=d<Hg=]Z8OFaHB;VfG/\[#6-O=ON[^eA4I(J)OVQf]C
D9DCP?4c==TDe_B>Gb]YTA&8g<S3U@)ReT#d@9ZGZG^f/YV<OfI]>Q;Wg+&5.eKC
>_I:L2dL.LRN(PHf/LX9RSL2C,;g@+HEF/3:?67N_.c>W:V0<U4ME4HQ.[GI<(_Z
dDRG1Z6f[,&SH2@AG)5U4de:aF>[.;(EV<]8(@OEOIJ+.>FeMY:YfgL;^QCN5B#4
3,+cS2]6:L+HMf0<;1cdD4EQ?^,7^^]_67R[Rg(\9G5<XE>J;Q2E0UVUCO,V^^I:
/KJe^IR^ZM]d,bG;B<3LGZYf(<\T&FD#3)4aSZaR)DZA;X7&V064EfO+d=cKbVJN
>TK-\3C-G\4^EIJ&>gE1d.dHS\.eC=K)Ib[G&gKR@TN?1WDH;b?E?-@WMP&1\4de
H2B_\GL+Ja/85.:<.N>ARPD0ZN/EDG;,<:U7AfVcQUMA;)+FH2AI=J;<,73V2f\D
@#UGWM13]L^I@OE;#;c<8<gaL;NXKKEE8B36>3N/>eU@M<G--06(0dBgP?eO75Kf
G)&R[;>O4aOQ7)<=>KV&#W.D.5YS?7-TaG7EHSd;G5V>G3)c1-dbN@d@YP5@L.(8
VT5V?M9#)AaMWb3e36_;W&UIdXV[;6VAEZO@Q+66GaJ7&EQN<Ea92Ad4W1cIIZcb
bN@6@X>,QFXc7R_dScP;94NA=P9CWPV?2DEb;>]eMQ[FJFeR;2?892I#f)5C=4&U
GWV]47XDQ;I8<;IH;Wb\4b&gVTARWc]+[F_3YH3ZQHd[IY>0[+eSEC?W;=^_3#<[
cTZW>AGWUPU^1<:I2UE0Gd)QeC1f#d\#CeMMB]^TCSFR&.)PeFCV2TAB[c1#<NgM
JBP;,PPO,aDX_eZXV^>Jf]QOM:d4760)40I:VgE?:6CWKR^D;#,/<76Re+3U<P&d
dI7g@FcR0K@4J9Y(1-ID)DB0CFD^1e][;)(ZSFPF#AACI[?YV<2Z0P/Wg?YPV/.D
f6A><S)g=6.eL-DVQ<OY:>[Yf0RK35-9eQd0M5,.I;D+,(8R^)VW,X/_WS[eW3;5
29GK8WcIOB4Y6aY@02D4>Q#df2aOCYfJf4_/_&K1R<T4,ZcU<T(bABf.9./Ng4Hg
N_342BRc</0W1b4V)(D175@K[]\0:\B;5X/(VIJOD@M02)^d5@;-?Gd9eJN34_>I
]FDS)[SK,+RSS073fd[/Jb-#]A:8F8/)^(5c7I3U-5V/,D3];[_N@?JW[DaB>;M-
#(7:,cAVfR,@1873K9g#B2_]MGZ8NM]GQC]Dga?CB4U5&RR46TDD?MRPA;cUVXTS
MCS)&ScG,/4>Q/^N;\7X#JDb<5?D?0.J7SYc=b9NO6;gIe:J1#-K:Ka-\(QL_AOD
=Ca,>Y>MP^WB\Lf:/Vc7OgOGTBFKK@Z5\aW5=F_0+KF#f+XPS+=)VR0Ia:JR31,;
f1QS8^0@N]JKKV<L9A2MMEENI-/:0N[SgS9A@_#;H>?32_1)U3[O<g&YZ,>>LAIK
@KF/BO=&dU<(7a8f4VEUWNO]^+GW1gMA#@GZ^-9I1TcL-PX<)F:A/caRRM+Kd+J1
@E^cYF4NW7+0+4Ofbf_5Z>,03J<f]?@+D./[VaHB>](+._.&Q_+>Id#&O=WZeA#d
&3>@2^&>[bY,?_8XfB3dGMKA6;OE@4/3G)7C)&e;T5H2;T?J\&SUUYC)_CDbJT@Q
4Q5AP3d+Qa>-A/)J^+-A=-LMOGS7+F\UD=GINU7G/daO<K#G4VVAAZWKK#e+d2_U
0B[cE->,9aOC8Ib.QEP\&Yg^&RKCO+:NS@7,67R1)>FK_0&7(V0TcfVMX+^W/+2E
fVI]J8Z(Q(UFfW^_:d_a8BVP5U79<c>a<C/c-.VQHJVV:0P?L/A9P(/H8#6_bF51
AH<5bfG.Kae=/FI-T2:HXOZ[Z^bF#G#KEc_2RP1FX,XKV.Wd7PJ87.U,WCeVQ7ZF
dN/\I09N]N&egGgFY_6_991/3XRMG[^(X7,_=e(Xd]JBaE15/_.F/Hdg\G;IgWCW
&/0MZ]GOa_1^dUDFAGf<c3>ZeNN=b-S.^W3F7^b[SN_;JdNN7;bD,,>b36N47:OB
PagM@K16[P)0@E^=HC-5)e7,6>e@.-/5=\;K@Vb_T@dGCcTOG/K0Q);2T#7\6dCO
:5[EE/[KQ^UJ5;:\ZPT,^A7)4-FOT.KUWaf)/R/F.M9d\\WD.U))8.be#;d5(EB/
@UA_#QMHI^6aFfM03WDA6c_V(EO&H7EUTQg3)WJ60dNL5V:@_gI(N,#d)SH-IgN5
;I-gGB&]],XHTB)\J83Dc)(KNa&.f6Q&0XQD\>b4Jd40]e4W2K+c1_dT/]_L4(@+
MIf8.EWB#N[DL,?b--aP5;CT8,7>g]SdAE<S.DNJ@B;+VdN1c<Z.fYWF8E5DM9TJ
09IL(;@N\-8AQc-#2WL4W@_N)81e_T-VH1J[G5C<dJ^@8:7&Ieg,G&,V+&R3N/g[
SS&7-DS;[N7f^?aQg>9;60#-=3<-UN@0+O=dUE@U@4#],L.O0,-FZ3#CR@KT859e
,6C\&a5HF:VgSI#,,@XV;YM&8O=O?f5SR&GFGTZSa;<Y0-2;9JaWL:VG3QE:VF^I
IF9_TY4G(X[ECJ[WI43.P3<4dW/PQB18P_c7M1=[E;\3HL)(YRT._BD[56bXC@<A
2HYANZfU_&LCW)VCa5aSVS7>PMVD^=b>@SKG8N(d;KMC#YL>DP-9+>\\9^AV[FFX
,U8bB];CdJ;YPR]CP6>V:601S&:1_:B[_<LD4N+C<X[PY:B1=d(F24&P\-H&;A26
]L4X-RO347W7EBbU)95<0M]N:>.J-LDDVXV77CfOA,+MTPB>?7)=NPF-9;gF?,<+
ED?_;D9]e:^[TO=++XINe(4X[(<=aXBZgT@L=;:bb/8C8)JO;<e-7(<V\=1),@UY
79??26::c&+D7\QL6f+BNE6R+NHc8#_+9f6WHJARH2#.S3#a\eZ:SYWYBXYGY;XP
U88EdAIVcf1(,7RI?#D.X^?O?.:F7+c[8L1COHPag;HW9JcL),D?+D_^USGKM<):
caA6?F_U5FT@.=M]3O_W&^\Q_?cMcgH)J0C(/?>G>;6;&@Pd><NUV;[A,=cIc?Y(
H>6C_>3>Z=.@e]#Hb&F(]T=]:[_)e?He#4(d\>]g(TdH:P4H_]4b9=cJP\gA;9/D
#DTOaRVG:P))HOeCGMT3@48gE-31OMRY&1]gL<\Xf@<MZCLF_>)@:1DE\[HRVL<D
abS,bQ2eZ393/-CR>^J)2EJ\4[7?d7O1EXL<\dVS[eaIUFXg-gc@S\Cd]TeSTT;G
c49;-U;^RXBT^aN(g3V9gR+5229WgAS+(#9Z:<;JC:QG87H)@_E35QB0[-HM>UgT
/WDGKTBHEee4NP7N:U4DSZUM;cNP[-XV6;\2R]a_fWCT/4KLEIKc6aTMcHAeH6Gg
>ZTaG7.1eEK#U8=\[CT1W\LG]U)Yf2#@\\gPK5D,79:O]]:_@D-I]6CML^dWCOcF
EHL<@;LTe@)^DC8e2.aJ3ad)>^LR82Q/P+#J&E[\\Q[:1C\BYVU3=KW^CAM/GYNS
WEDL<W,C9D110#EVg]>fQW?[+a,[_YM)8Y##IB^&/E+<c-NY.^G?Lb[(HOSd\&8f
_Eg?Q+U1M^,[E=;#2@M;/U2L4TH_L+C)[@MZ)->Z5W;1ZKC6(ODU?&94g<OQO^:?
b,+M3M+/6K[aDM:61@^/,FET:cL\BJ669-Se[M<NAD?3]MaSbPdU\-TJKQ:JRB/H
]?B,bOZY>DKKP&9)/=5V?@LF)d#H)J>f#?;bF\F69VWJ6&SEgOgI33&\R]#=;aeb
1M_ZC3K>R_0AVYeBBU3]\U@E_0ZFO)8OSPHG(?6&1[Xf.NCPUH[=Ta5>8b/Y>@08
9?\3^dYB7MSe&AMM<-bJD5/Gf4b,E=fgN?3g18+YK&YU7]F#6SQ_88C#4NH_XU\A
gP)=Zd?d:_[T@K)B3.(a-@DefB..[Mg8,d@[03]UXO]IF\ZEPWU7c-84\_29F/S4
IG^L=+/]TZNU<dCA:O.\A=F8b0LWCMSO7a^RUbV3ac&H;1=b.Q^D1W\eIM>FXMf2
R?9I0b@1BPVDe)45Q3N;;,2&/4dL9/c@GP3B>CE>cG^HI3^f=D2\ceY7OIDET?FB
K1LE:\+4Yf>F^a..NXBeZ.NU&WdZT>J9#&27YUL&XCJA:a:9^ZRFS/9>Q)J.ZeMC
RQa]I69>VPY+/d4YG#9/UT=K[)17fLGbRcR^/fC7B0eE(;CA4C>O2OFL57U,//C6
:1CcZeM4^GgM<.VVRA?1A&TJT6\&S(#R.69^H=5^&d\7e=FO#P)@1P5VVWF(MM7b
g<\FHI(.:2I3C6WWU3[W@>Xf6T(&_XST&PU4C[)MAdY9A6]UddC><+4gU7(RUb^N
8K)G?.:GQD6(g=)-b..H4CEIgY=_[]S(fY0^#INTXcZYE0A6QB<S[R/B74+QGQb.
:KRHU4(28NG&1#U.]?PJ^31FZL]/D5<;cOMCQ?9[H[f<EB00Vg6L@+L=.>[3aO-D
?(;gfA3XBWCMR?55T2RZ+]A;QdFG4C;+)a8R3>)R&:S@HE08cQ@0)L8,DDPBL2^_
dgD4QbdS)\Z;.#dL_8NO()b^Y1^\W_;S5OKNBc_./W_D#M1We+bB(e]2Ya3SG8M1
U=P2[Y.[f-bSQY-N(H<D=YGV4P80)4Ig5>[ZKYK@)R8M^#Ld,6ML&42X>>PaE;<1
B:##bTI?+EV<>Y52aC:3T;g2GS=K5ORaHVB27FQ)e),1_V?\Y<L\+)343(ICU2b8
5S[YbgQC:Y=\Gc1fbVEA@BJF//UE<[OfSa#^?SE>Hb=[,HCbBB/0dMIL^CB>@:EF
dN/_D;Lbf-/))RAHFN;#]E]1-9_D22@IOdH>b?<cd[):\E29X/V_b-T<8F>VI9EE
#]YDC&#a-NS@RZFf-84JDH?B)N2UE_,=(FG0=S+^JHLY@gI]7FJXM=Z.2_6;Z-Dc
C9/2HLR_H6U\APEAN27]I)?bL;9:gg^-84d\J&?,WR@_=fce5/fQ,M<U#&MU^US5
/NeGLaCe8)b#I328<HF]:[BbQ<Z0G?J5\/X8fgCUd:J;Nb,ZP@JYW+@M^]g_T/bN
V#7_;),H.^IL_4CMF+bXFOaY=[Q#C,+Y=ZP=TS,(DS,>-)X_Z89@W[eNT#&Z,LJ5
7^bW2ZH.C5=7S1CVK^=RWGI,gG3>#I[.a@:P_FL3bPT)9:\gF@[9(-B1Dg[Z5LZ^
^:I1\0>;@I]/UI;UeW4S(Y\)OHK]Y(;6S5ZC;PET-]BO1BTK-\D1PJ^4bMcRX;56
c=V5436>,dI&dYSEOZ4<8R[M5UKP-fB:>V[HeSgAeQA3cf4/K,<YBcc:=a;Q?@P.
XX@T?A&8bM-55MeRQ<CCR.<>5GfJLM71&LS)XHeegEdV^5gQ(#gfLB>^;2EN]:3@
/3\b;62J)_d+Ba+8LE//#bZfU=I=L^W4E+fFBS<2g=V@,;bC#SBLUJAT^70:Q&(N
KDA9\PN8ZJ<&17,Q?b@V[KE#H.d5J4]4EZVHbaD@=Gd@Nc:[ZXX)[/&^UVZ]M(0X
\/N1Y^3<FRJFLB3-E9L7JKX./C5QdSPK9FXOI_MQ?B&3LDOe0.cES8MZZARaA7(P
Y,MY?@SI9IAXe8g7?0L?5aDI81;a&#=eYQ<I=1A:a1CDR[BZ.L=CVd,5D]&&3IeJ
ZS-3N^Ef2V72#Y<4FSCZ+BgWR=>14=KeUQ3<1fCUC/#d6K3O3?AJ)L/8X@NK>XPT
M0GE@V_)GA3T??gYPN>[2^W/K4N<B=Z+:(VN0\\_.Z;N^Hf]UKTDJbNQ+_GRIa[g
AG_ZL1C4F)Y.7f0b21)A?_HLN-0_-EL+&[_,&<e4S53HOF/d_:61#MTJbGa/GOUT
ANP)dg@BXgA^f7PZ7[fUaB9fV[b27#YB@HRN2HV<EEH,BP(M2gJ#UA\9J,e[CEX4
]/?:[Y?@Q.<T.fZ=f8DP\76TQMQ(+1fL&cF#XR84\TE\L(/96;?gV+TUZ,J/Z,Fa
L,8B_DUTE2:(^&PS\],e+[ERI2X.P//)c#)=:b>UA((ZaT9S[4=C(J>0AX(H.7)9
@;bGT7BU#YePc<_E3GU?X[/SRZ0)ICa1IHNJ2F]\<;5-g2ZJP?4\c<CCW;98ZS7\
(&Aaa<Q^6[;@.3JJfUNRXK9HIN],RF41J@g.]1&B7WIaA<JJ;BJT+T:eZ9fFEDO0
9BgL/8T+M+ZVA&XON\#;fE8,GddQ<(3QS5VH[G0E-V_>,Na9<FDWa9+LZ1Q<-UM>
aV.G\7D-V^RE>5=[UD]-DA879/FO/XG3UB7Bc9L)QXFV7P@SN?O5+^C6]AJcL6&B
0:DH>I1/AKAfc+_)V[cC)2gUgZ@=eT=8aM6,:(+S+c=:3=R/dKf1S?B76<O4aZU,
Na]^X]TJO/_LC@/g[&4>&fH[d-g#[7N>d3)YI^TWf&@CO,BE?;7HP0Z&&fO&bFb[
>TdL9Zd>VDOR+KVbM#c))LML]gBH5E?M_\\1YN0bf0_<[34b6O+JIdd87E)7Qb8C
911_/4c5QR=6+g1eX8S(8HRGC;+K/(+X^YP(80QI.eYXIJ@RQ0@TfGdEcR?JgWD_
1F/)(#9,;?Y0ObI@23^DgADQeaCO0+#=./GV>fE4S9,fR)Nb/^>UT0(HVRXg/cB3
EZ#D.E16K6Ac&1P6MJ<GQ+ZX<8+Md>=<Z-3fMdL/T5#@g7/R_67PNgGO8D,3P#4[
&#d,.E[f9ATVcT1A-18>eKN2KdAb63RNU);IdW,Ea_>,(Y9XQCbS)=LdV6GdX4/?
ZgNK7ef[)8eaA&.HEdNRLTg-Tce[+>WK+:&EKYRLO2e4L-EG][?e.4/YT1;M8FGb
GA(GJ(<Q<PgX4(;<JTKc9-a@&YH(FUSA7XPB\XEO^H:cU=7faY&eaPcg^?FQ2a2,
G]a\XgbY1/.dQ[7H:-X)<(=D.S0C<.&Ra)96YaL\aCD&3]+Vc+g;PEK?NF73L9e)
SXeHaH4MNc;@4>UggC\I-,B6V^2^X.A4+Z94#fHD\eeQ3PUJFOXXP.YbKH)#ag]V
OBI0Tf5e9G,SHafb/TG:HZWO7>8\C;<T:JD:H6_/5=H^>6e(c(ENH=S-;VbM\-?:
:9SUM<Z7X;3VbA?3O^+VBUG+Bd9dA<#W0+4O>36_)K4Tdc9&GLdGCFd[f5;cW>.<
Y()H+cOKJf31,;gCHXS5>6WLZ:L)B/[/<.^EIVI2<3KGQedAMK+^BQXZ9KIUc]B-
XPKOUMT/37F,)U^A#+.1GeJ-Pd\9e3gQ]AW+9)Qb,N,fWDJ)72>U1L:G7R8OIIPR
UDeJCR[X:gYMG_ZgC-F:67cQ1>@Le#cNP.(VYbe\C@WT58N8eC:g::&,cS?N-Cf0
A:G?cW=:VI\5;e2&B;_(>7]Me+g&MJ3JZ0Q+&/3Q-?E^GgOQDFB9LeU<7QBK=RSM
V,:)R/\UeUE([><4X;aZVI^eVGG-E9\cE7CCR1WG-W&]E+Z>\[?d^&Ua8+dB<Z1T
ASDXCLg^OBd^fH9A/S5&M_ZM:0F5N0JA=S>5c4XQecN7VC&.&(1SC>60(2PA>#:]
D:N49X7E=@&W\U?f1S3D@;^V?[8eZAJ4U.]E/H[[?cI.GHW#ZR&T2CC]E<CZ88cR
WLW=5D;c(92):BdG-5/;GU@#P/R8TD<5C,_T7UHYdZJ&_7BUdSRS,ccSgV7#;^4b
Hg3I.UHB;41WNV@bS&H^MW.59Y/JF)Z:&IRRO89SGHE6+WSY^W+VM9[Z\1=1?K-d
WF;cTTA+R#a;WcO(LeB:ERB8eg=+AX(dY]8U5=LR\TfcJ@<SV+R>N1W3T?XRc)[K
8&=6-75De5Yg2D;R5QCf9\7<8F[0[=4OSF+Ve9fC0+,<,5T1a(7c1dR^5HDAaS@S
aZ47M+Zab^.)bPNRUEKSY>a/JHKS@=QI@eK=A3>\7JM;EIacAKX;GgFg\@]\/4QM
PNP<K)(F\=;=LHePP)BHWR\R<<7Y=-^ZS20JY]@RJF,VR;XMe:a4RK(P.)J2SFII
@EaH_V;P1g+8geg_ga2UXRE]\;2WZ8ac]P:F3-V#)I[7]bgVU9[6,;I@M4ILID-#
g<O^a9JCKa]_[DaEM\3ISPF)R<-RKbG#U[R=4f\O2bX&MRGFQDEeFSTCcL.dX(C3
-,I9=9@2f20PD(PX&SZ4IPDLT@J.V<<_E+abfCC59[^RFU>6;?EFPNT-EgA_4aMT
+^&UUPEU1_+HSP<^UEd>g[&63AVd(a?DU0gG^Y]QacOKg6L&MD3Z]V^=>HFE84,S
^X)-LQ1DNWNM.Q@&ee@g0UIFW&]fD)<cWQO1d:/_:#4R>4B6&><;a>8,b;_/M<CN
L6T21M/[S3f-NC8XO6BedQJUW_H/K\WJQPVE5C->Q2T4L?eeV/^acF(7ZEgHDcAg
@#g(YVRda+;=+J:):KX[^DNJ3/>FIO>&WEaK@9,HR>F.5/==)S#F+_K)9SWJdaK;
MTf8ZK[7)?&1fc_8WbGeK]M2S]CgI1[&1)?0O:81LM8PKNT2[,>/_)gQ^bN.RX>^
d5AU(G:LMRZP-Cg51a:E+=@>A0@@)4?8@D?8+]L.:.Zf_Y0cZPJ8_]cBG&5J2[6.
BdL=H1N=FR5Cc9]H=\cK:eO7d6_3NB\^;VA>BfFbC7A+,)OGAW[O87K^g>?[;NA0
];A>SIQc_@fMc9[4[2gA,@65)CZ;]OM9QW]Waf=caM^Vc=#V&NZ35Kg0=NIO]9UM
=]cK&I1W:5>_^9/)C=gXOYAdMC9P]f\SV)+=#2#Y)_CD-<-3=/fdbKJcb,Xa#G>G
cCG]9b[5_;=,&LBJ5IbJ,>/=L(5:U,6Jf[/@[FLZ=dRCgL+6,dFMYB0.F.33\9d=
GEc[:I-]8K9,^e\.3PV2OE^cL?g1L2K286e@RO3J>cR1CKY_CG/Q2a?M4R=.8P^F
_UT3FgW;VMHfK[@\f,,D[Y(7LL?U.7P((>09\40^=(E^N1TH\1()U1<TBO((g]M:
]6;EOI9M--_>_JWI1O;(Hd#-JaQ7<[DGA6X;J/28d4,D,bZ\N027W\8)5F9X?P<\
(e7;86(aZQO&JR<IX[N]f\c/@6(G]2X5RcGZ14g72GPI\6NcS_\Fe4T^OfECEcL2
c,3T3_CPceffMVdBTR.f68:_TUc,HWc0(4B2(@Qa:K_VgL_ZV;PM?J>6^Zb[dEV/
A+fP\e?8U0],[=E/4BB(LOQOQFI,O_dF=_3OdA2eW7DTXEbcO,.X+e8YKEG+377^
0Y8\YVY9W-JA4E80Pa51E-3VH/[9(I3g0/IB?0.;(/+Kf5<MOgG2JQS2EV_7=>]S
Ub,F50.;?IJ]B+2#L9fK,g/6SYK-1Q0O3X/K-Z3;0XIe4_0U9Oc^DY]-&I:::;/7
6HO9JP?,5-3#CYeTJYV821+JfBNE^Ifb-9eSDB6^;LUMHc;C;GOMX;1cIFI23P:.
YV\_d#=O8LB3L2IDL:;ES?-,PA#EBJV8>b/)B<>29P)YQ-Hb/4Sf[2TLUX#VZ_?9
?XEZQWGSN?-gYYaZ)R-=).4F:eRD76;UHPaG\40fV8K^H.>S?)^B5:P49O&eb]3,
gI)3GcW>@V3Je5?=VENI<2AMRV6KQAB)T(&<8U:#9g6S?-N1(&V&TOgAU?FLVR_D
NY=LHKHN3ff=67M+^)+BR0cL>>=6LLCd4:8];94D8JA8)1AH69)B>WB,2CccL-#)
U.Z=+.CaWU7TGd,\-U1c=>TVfVCcF9&WF1Ugg[K&,GbgW^fVFAO+1a:()-bJNe_Y
;Ua4I:,=AgY#.@Y[ad^cIRVPb]=BG>J\9WXbK:C#aFY=+.\XSXF-:Ha;#U(T@<DK
9d;?11cb>Aa/Z+FLGDe_]3(V(Z(@S/0g_=?eL:LJQ@<+FfEDR#^fN_\U5C82[YS+
N+)+MBQ\EFCZ]U>WBdFaTb4,=7QP8-[2#-E<C-8=T/BbR=51[Z=OTGC].cLXI]KA
5:6&7N5I@/8RBK3.&TJY0Y9JeB.7@.4_2RQ3-YLcHO6D[,a.25]&E]EeS#_+/HZH
O6A)d;E6]HN^g0L.Q54JI9F:D(;+fODUdc#7?Q=QX#S[&(,U.\cA1c&C13A8a4/U
6+5CYe81B691?;7<g38PMP6B3#5a?]9NO,4-=_gV??6M6G-\;eGPY4JGJQb=gWKK
AXZCS[4<;d@g^?GgLENLQ08G?Hc.<2KVfFGDI>SOU?89/I^B^TGF0<;O^IIQ3<Y7
;e&B42N\)51@3+_;bW&V2F]3473_@WP68#[\YP:B1#T(0V7NHC8dY29+/aIRfS5Q
8O\fQI5MDQ87WX8?FKTMHXTMOgS1AC/Tb1Q\-eBd<a[#dcKS\a9S?#0,\N(SC]CJ
WED3FU[3C,DJJLN]3=eYEH)YK+V_Z]EY,C-FQ/ZRRV.QX6S&M6d9IBMW:8/PO99#
0;f\W4^K28FKU<6dK@4?JRB4:R=?-e0c(gTZ;(VT>Ic;g(,\&UH+H,-[ddV)6g;,
a_cG[T(BY>a7ce0\Scg6>P<Nag@.YW_;JJG/C=4ZR?J;E$
`endprotected
  


/** @cond PRIVATE */
typedef class svt_axi_checker;
typedef class svt_axi_port_monitor;
typedef class svt_axi_master;
// Utility data-type used to capture QVN Token related activities
typedef class qvn_token_pool;
`ifndef SVT_AXI_DISABLE_SYSTEM_ENV_ACCESS_FROM_AGENT
`ifndef SVT_VMM_TECHNOLOGY
typedef class svt_axi_system_env;
typedef class svt_axi_master_agent;
typedef class svt_axi_ic_master_agent;
`else
typedef class svt_axi_system_group;
typedef class svt_axi_master_group;
typedef class svt_axi_ic_master_group;
`endif
`endif

`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_base_master_common#(type DRIVER_MP = virtual `SVT_AXI_SLAVE_IF.`SVT_AXI_IC_MASTER_MODPORT,
                             type MONITOR_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport,
                             type DEBUG_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_debug_modport
                             ) extends svt_axi_common;
`else
class svt_axi_base_master_common#(type DRIVER_MP = virtual `SVT_AXI_SLAVE_IF.`SVT_AXI_IC_MASTER_MODPORT,
                             type MONITOR_MP = virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport
                             ) extends svt_axi_common;
`endif
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AXI interface */
   typedef virtual svt_axi_stream_if.svt_axi_stream_master_modport STREAM_DRIVER_MP;
   typedef virtual svt_axi_stream_if.svt_axi_stream_monitor_modport STREAM_MONITOR_MP;
   typedef virtual svt_axi_master_if.svt_axi_master_async_modport AXI_MASTER_IF_ASYNC_MP;
   
  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_axi_port_monitor axi_port_monitor;

  svt_axi_cache axi_cache;

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Master VIP modport */
  protected DRIVER_MP driver_mp;
  protected MONITOR_MP monitor_mp;
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
  protected DEBUG_MP debug_mp;
`endif
  protected STREAM_DRIVER_MP stream_driver_mp;
  protected STREAM_MONITOR_MP stream_monitor_mp;
  protected AXI_MASTER_IF_ASYNC_MP axi_master_async_mp;

  // ****************************************************************************
  // protected Data Properties
  // ****************************************************************************
`ifndef SVT_AXI_DISABLE_SYSTEM_ENV_ACCESS_FROM_AGENT
`ifdef SVT_VMM_TECHNOLOGY
  protected svt_axi_system_group system_env; 
`else
  protected svt_axi_system_env system_env;
`endif
`endif

  // NC gives this error for these declarations (not currently supported)
  // Associative array uses an element data type that is not currently supported [SystemVerilog]
`ifndef INCA
  /** Associative array of the send_read_addr process indexed by
    * the transaction handle */ 
  protected process send_read_addr_proc_q [`SVT_AXI_MASTER_TRANSACTION_TYPE];

  /** Associative array of the receive_read_data process indexed by
    * the transaction handle */ 
  protected process receive_read_data_proc_q [`SVT_AXI_MASTER_TRANSACTION_TYPE];

  /** Associative array of the send_write_addr process indexed by
    * the transaction handle */ 
  protected process send_write_addr_proc_q [`SVT_AXI_MASTER_TRANSACTION_TYPE];

  /** Associative array of the send_write_data process indexed by
    * the transaction handle */ 
  protected process send_write_data_proc_q [`SVT_AXI_MASTER_TRANSACTION_TYPE];

  /** Associative array of the receive_write_resp process indexed by
    * the transaction handle */ 
  protected process receive_write_resp_proc_q[`SVT_AXI_MASTER_TRANSACTION_TYPE];
  /** Associative array of the send_data_stream process indexed by
    * the transaction handle */
  protected  process send_data_stream_proc_q[`SVT_AXI_MASTER_TRANSACTION_TYPE];
`endif

`ifdef SVT_UVM_TECHNOLOGY
 /** Handle to the UVM Master driver */
`elsif SVT_OVM_TECHNOLOGY
 /** Handle to the OVM Master driver */
`else
 /** Handle to the VMM Master transactor */
`endif
  protected svt_axi_master driver;

  /** Internal queue of pending trying to be active transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE pending_active_xact_queue[$];

  /** Internal queue of active transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE active_xact_queue[$];

  /** Internal queue of locked transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE locked_xact_queue[$];

  /** Internal queue of transactions taken from channel or
      auto-generated by VIP, but not yet added to active queue*/
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE current_xact_queue[$];

  /** Internal queue to buffer the incomming read transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE read_xact_buffer[$];

  /** Internal queue of buffer the incomming write transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE write_xact_buffer[$];

  /** Internal queue of buffer the VIP generated WRITEBACK Transaction from
   * CLEANSHARED or CLEANSHAREDPERSIST or CLEANINVALID transactions */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE writeback_xact_buffer[$];

  /** Mask to get valid bytes of read data */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] curr_read_data_mask;

   /** Mask to get valid bytes of read poison */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] curr_read_poison_mask;

 /** Current owner of the read address channel */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE read_addr_chan_owner;

  /** The last transaction which was the owner of the read address channel */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE last_read_addr_chan_owner;

  /** Current owner of the common address channel (when enabled)*/
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE serial_addr_chan_owner;

  /** Current owner of the read address channel */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE write_addr_chan_owner;

  /** Current owner of the read address channel */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE write_data_chan_owner;

  /** Variable that stores the read transaction count */
  protected int read_xact_count = 0;

  /** Variable that stores the stream transaction count */
  protected int stream_xact_count = 0;

  /** Internal clock count from rvalid to rready.*/
  protected int rvalid_to_rready_delay;
  
  /** Internal clock count from bvalid to bready.*/
  protected int bvalid_to_bready_delay;

  /** Variable that stores the write transaction count */
  protected int write_xact_count = `SVT_AXI_WRITE_XACT_COUNT_BASE;

  /** Variable stores the number of active xact count */
  //protected integer active_xact_count = 0;

  /** Variable stores the number of active read xact count */
  protected integer active_read_xact_count = 0;

  /** Variable stores the number of active write xact count */
  protected integer active_write_xact_count = 0;

  /** log_base_2 of data width in bytes */
  protected int log_base_2_data_width_in_bytes;

  /** log_base_2 of cache_line_size */
  protected int log_base_2_cache_line_size;

  /** data width in bytes */
  protected int data_width_in_bytes;

  /** data mask used for sampling data based on data width*/
  protected bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] sample_data_mask;

   /** data mask used for sampling data based on data width*/
  protected bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] sample_poison_mask;

 /** data mask used for sampling data based on data user width*/
  protected bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] sample_data_user_mask;

  /** mask used for sampling ID based on id_width*/
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_id_mask;

  /** mask used for sampling RID based on read_chan_id_width */
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_read_id_mask;

  /** mask used for sampling BID based on read_chan_id_width */
  protected bit[`SVT_AXI_MAX_ID_WIDTH-1:0] sample_write_id_mask;

  /** mask used for sampling addr based on resp_user_width*/
  protected bit[`SVT_AXI_MAX_BRESP_USER_WIDTH-1:0] sample_resp_user_mask;

  /** mask used for sampling addr based on snoop_addr_width*/
  protected bit[`SVT_AXI_ACE_SNOOP_ADDR_WIDTH-1:0] sample_snoopaddr_mask;
  
  /** this flag is set when reset is asserted synchronous or asynchronously*/
  protected bit dynamic_reset_flag = 0;

  /** Variable that flags if DVM Operation has been done before
    * issueing DVM Sync
    */
  protected bit dvm_operation_done = 0;
  
  /**
    * Variable that flags if DVM Complete has been received before
    * issueing DVM Sync
    */
  protected bit dvm_sync_complete_done = 1;

  /** The cycle in which last crready was driven high*/
  protected int last_dvmsync_crready_cycle = 0;

  /** Variable that stores the DVM Sync transaction count (received) */
  protected int sync_xact_count = 0;

  /** stores count of auto-generate transactions */
  protected int auto_xact_count = -1;

  /** Object used for randomizing a transaction to drive random values during idle*/ 
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE idle_val_rand_factory;

  /** Transaction currently being processed in add_to_master_current_queue */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE add_to_master_curr_xact;
  
  /** Sampled delay from ACVALID to ACREADY */
  protected int acvalid_to_acready_delay = 0;

  /** Variable that stores the ACWAKEUP assertion transaction count */
  int awakeup_read_deassert_count=0;

  /** Variable that stores the ACWAKEUP assertion transaction count */
  int awakeup_write_deassert_count=0;

  /** Variable that stores the ACWAKEUP assertion transaction count */
  int awakeup_toggle_assert=0;

  /** This bit stores that, AWAKEUP assertion details when ARVALID is asserted */
  bit arwakeup=0;
  
  /** This bit stores that, AWAKEUP assertion details when AWVALID is asserted */
  bit awwakeup=0;
  
  /** This bit stores that, AWAKEUP assertion details when WVALID is asserted */
  bit wwakeup=0;
  
  /** this flag is set when ACWAKEUP is asserted for read address*/
  bit active_read_addr_chan_drive=0;

  /** this flag is set when ACWAKEUP is asserted for write address */
  bit active_write_addr_chan_drive=0;

  /** this flag is set when ACWAKEUP is asserted for write data*/
  bit active_write_data_chan_drive=0;

  /** this flag is set when ACWAKEUP is asserted for data before address transaction*/
  bit data_before_addr=0;
  /** This flag is set when new trasaction is marked with highest priority*/
  bit priority_to_new_xact = 0;  

  // ****************************************************************************
  // SEMAPHORES
  // ****************************************************************************
  /** 
    * Semaphore that controls access to the active xact queue. 
    * Any access to the active_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_xact_queue_sema;
  
  /**
    * Semaphore that controls access to the current queue
    */
  protected semaphore master_current_queue_sema;

  /**
    * Semaphore that controls access to logic that drives rready when
    * the default value of rready is 1. Look for comments in 
    * the task drive_rready for a detailed description
    */
  protected semaphore rready_sema;

  /**
    * Semaphore that controls access to logic that drives bready when
    * the default value of bready is 1. Look for comments in 
    * the task drive_bready for a detailed description
    */
  protected semaphore bready_sema;

  `ifdef SVT_AXI_QVN_ENABLE
  /**
    * Mailbox of "`SVT_AXI_MASTER_TRANSACTION_TYPE" data-type
    */
  typedef mailbox #(`SVT_AXI_MASTER_TRANSACTION_TYPE) axi_master_transaction_mailbox;

  /**
    * For issuing a transaction driver will typically spawn process threads of
    * send_read_address, send_write_address, send_write_data. Each of this 
    * process will require at least one token to be available in order to proceed
    * with each transfer. So, these processes need to inform "qvn_process_token_request"
    * each time it is spawned off. For this purpose, each of these will pass
    * received "axi_master_transaction" (xact) to "qvn_process_token_request" through 
    * respective mailboxes.
    *
    * "send_read_address" will use following mailbox to send xact handle to "qvn_process_token_request"
    */
  protected axi_master_transaction_mailbox qvn_read_addr_token_req_mailbox;

  /**
    * "send_write_address" will use following mailbox to send xact handle to "qvn_process_token_request"
    */
  protected axi_master_transaction_mailbox qvn_write_addr_token_req_mailbox;
  
  /**
    * "send_write_data" will use following mailbox to send xact handle to "qvn_process_token_request"
    */
  protected axi_master_transaction_mailbox qvn_write_data_token_req_mailbox;

  /**
    * Each master needs at least one QVN Token to be available for a particular Virtual Network
    * in order to make a transfer to an Axi Channel targeted to same VN. For this purpose, each
    * master needs to keep track of each Token it has requested, granted, when it was granted,
    * tokens that remain unused and remove a token when it has been used to make a transfer.
    * It also contains semaphore for getting token statistics and requesting a token consuming time.
    *
    * Following QVN Token object queue (one for each Virtual Network) is used for Read Address Channel
    */
  protected qvn_token_pool qvn_read_addr_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Address Channel
    */
  protected qvn_token_pool qvn_write_addr_token_pool_of_vn[int];

  /**
    * Following QVN Token object queue (one for each Virtual Network) is used for Write Data Channel
    */
  protected qvn_token_pool qvn_write_data_token_pool_of_vn[int];
  `endif

  //vcs_lic_vip_protect
    `protected
UD<b^DVEO2&)M<WT,,FaEA+<XS:5[_5;QZ[:J;-VJ7^Y2J+;XBO)+(:gAW=F4OUI
77W9Pe&DK[E:DecSZg6JD-b?Q7=JDP>c:Je32]Q1.##g1)(8PQ+W/e4(&ee=Y?_K
-3,e@feWV.;EK#IQ10-X6<R9#.Oe4)GZg@40Lf:cb(+8D(UJ&D565NYac((5_OTX
UWDF[Q^=8:HKJEaSFQ/])gH2d1<c5SI8+)f<<9\f=DM.Q,P/22P]0Y&I6S&CZX?W
0HPHG5]Z_G:7Nc6<CX?VUF\?;D/cG12gTgM6eJbZP4I119>5J#fN,NH]?G927UcZ
5E3CIK9J.aZ8@gd>e^P8I]ReOS\MaV?@g2DH0\be_[WeUK3cT)7aYPQP(:2G6GUL
[R?Q<K)OdEV(LEM)<c_dK@TT64>FF7(.;dNZ,?^P_fO[dP_g#23?2e?9AaWZ2P1H
QMda2O:5.ZT-@/f=(&_5e@V,>dGNRZC425LDV1\BYeWDGML2DD:PZXL/NXGX(dW1
c>JOS&@:Z&1@f[YUE?CdL25[M^DB:(FJ[/R#CaE<fY2#P<@25N/=WM;&aGeJ=W_)
LabA6(G,=7@#6D8GG5ZH]7?_8Xd@(L/+g/2,JgWD9#,75-ON)6U0,3@,d^eMI4.R
8NCKD#OME;(VQ<.G9K.A?]ZUf;)[.;;R\^B[S.dV.3MC>C>^>.\[HP7e++d8cG8V
77edYI,D8&e-Mc))1eG<d?T;b517<Q\Wb+;9Z6ABLZf6C7Ve7JFOCI/CHKc,LV5<
g5>W6Y;_<cdV^QEdM6.ff[DeH1^6Z.6f<,(@[9f;A],3cL&R]>^Mdd3>a;b;c,Ve
R>cQS/ZPAa,Q8I4,@\OA+7@^6AW2TgAf^JL<Te94;,295g=]fV_?c,aM,d95>e]-
2W9CA8aT)K/AF==d6f-//7HZN-DAKFQ)[;f&\-L@YK)L?VI3H?Y3??a\9]DLBSQ<
5M&YQ(QEa:Q:]<a^d4U?6B-cAI^-[4?H8I:C6HdR]9PJ7\3fOCAU8=XcaT=LY&BF
0UbVB9)2KF?0&BS;g1+E+T[,8.7]B8Pd-[O0WXK5&#(=@&a4>6^Y,ER2S7J/P:LJ
/(Z6>,(3fWG<NUKFgfaLY=).d^/g^4;8e22UZ++6VB\:\?O2PGLR&WDL>:GX=]\;
MK23>;<;_LA7+af_X)-^CCf,&d)R+Y/&<?,;FDS3BV/D-?f6<FF<_D)9Gb0&-@14
f7XZf\,KEK,6=>OJ9Y#?>#4b>B@[f?bMda/ZO^8/eCI,M;T@ZI=J5Z0+4g6OJ9+S
7:K1H0S&f</[58OO>^\5><M2[Z1[I:(c_9B/W[<B/0913fe.Qfe?3P].4LZ_)Gg5
9JAb4IC;gdC#M,2CeM9/^[2D=+(U/U.MT2SfUK9RKXK#@gDaC;:2W>8PVWFQOfe&
R\SV(;bH]-SR515[0<B+L=^=_W#K=J&gH^^9<@SJZg/VM-^-gB9=^dB>U5U\?38T
a==&@e^Y->c;ZDFMPIH?2WK\Q)RF/aH<V/SFMZb<&<F]RLO2&G5f2>84BTZ#S7+-
&,+g^f_T4[,W#SP@E_ZS<M@/eg?6+_\2\WB+QX+IR@WeN22NJ#cAQ@YaD4:T_I3#
/c@TKJNMA\>L9#C?F1+:Cb?b45c>bB<Hc2KSS3OS:OXeH$
`endprotected

  
  /** 
    * Triggered after sampling at every block.
    * The event provides a syncronization mechanism for all
    * the processes that are spawned for each transaction.
    * Basically, waiting upon this event ensure that all signals
    * for a clock edge has been sampled.
    */
  protected event is_sampled;

  /** Triggered after any transaction ends */
  protected event transaction_ended;

  /** An event that is triggered every time a valid is asserted or a handshake
    * takes place.
    */
  protected event bus_activity;

  /** Variable that stores the auto-generated transaction count */
  protected int auto_generated_xacts_count = 0;

  /** Variable that stores the dropped coherent transaction count */
  protected int dropped_coherent_xacts_count = 0;

  // ****************************************************************************
  // TIMERS
  // ****************************************************************************
  /** Timer used to track arready assertion */
  svt_timer arvalid_arready_timer;

  /** Timer used to track awready assertion */
  svt_timer awvalid_awready_timer;

  /** Timer used to track wready assertion */
  svt_timer wvalid_wready_timer;

  /** Timer used to track tready assertion */
  svt_timer tvalid_tready_timer;

  /** Timer  queue to store timer handles used to track dvm complete on read channel for dvm sync received on snoop channel */
  svt_timer dvm_complete_timer_queue[$];

`ifdef SVT_AXI_QVN_ENABLE 
  /** Every time a Master requests a Token it waits for corresponding ready signal to be
    * asserted by associated slave, indicating a Token being granted to that Master. 
    * Since Master can't proceed with a transfer without having a token so, a delay in
    * granting a token i.e. assertion of corresponding ready signal may increase system
    * latency. For this reason, a Token request must be granted by associated slave within
    * a bounded time - configured in port configuration :: qvn_ar_token_request_ready_timeout_for_vn
    * If a token request is not granted withing this specified time (in clock cycles)
    * a timer used for each Virtual Network for Read Address, Write Address and Write Data Channel
    * fires up and asserts error. 
    */
    
  /** Timer used to track qvn read address channel token request grant ready assertion */
  svt_timer read_addr_token_ready_timer[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /** Timer used to track qvn write address channel token request grant ready assertion */
  svt_timer write_addr_token_ready_timer[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];

  /** Timer used to track qvn write data channel token request grant ready assertion */
  svt_timer write_data_token_ready_timer[`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK];
`endif

  // ****************************************************************************
  //                        SNOOP PROCESSING RELATED MEMBERS 
  // ****************************************************************************
  /** Variable that stores the snoop transaction count */
  protected int snoop_xact_count = 0;

  /** Snoop transaction that is not yet in queue */
  protected svt_axi_master_snoop_transaction snoop_xact_not_in_queue;

  /** Internal queue of active snoop transactions */
  protected svt_axi_master_snoop_transaction active_snoop_xact_queue[$];

  /** 
    * Semaphore that controls access to the active xact queue. 
    * Any access to the active_xact_queue should be via this
    * semaphore. This is because there are multiple processes
    * accessing the queue and it is neccessary to have this kind
    * of access control to ensure consistent behaviour
    */
  protected semaphore active_snoop_xact_queue_sema;

  //vcs_lic_vip_protect
    `protected
0d258#_IO97XSS=]:AL-4Y3+:56(@F8:FFgN(cO<\B6-e12dIBQQ1(R<+V+_3[[&
@-M/T9(c)Z3JSI:7De^67K#c/.?E6N28E]PeMeaXLJ4SG2+=^++11YSBNL+&=VR]
RS.JCQD<S4WY3^A>a(4/ZUSBI@90Q?V2E^E,XW^1NU;B.0>/&,\U3)?+,:AG6P\N
]8KO<46ZeWaY_E[F][#aI3RJ:<12c:@M,LO\&>\56T^W]?H73WK+cH2E)(RK0ga,
DD2@a&4E3bZAZ<+SSQQFab#[SE)BBU6S^?J::2V8(bLLd0EY?J,WEf_9Y6HQY)U(
Y@)8X[.22GW(=RPgF0dIHKFG3gD2TQC;Kb4/Q4g>DUC:dd.eGSE7;RgQN6OI1&ML
;O\TSbV/;de-G&33QdE7/T80P]LRCW+af]/.Q@RD5SUb,IWPWBX)]=6&[a]WJU5Y
ZFPg8SF,43CQB#U7C4:Y_=VZ[KQ0)V9,,/D#1De#:g\f6B9JN_&g5f0(8Y_D8S9O
MNM\7J95D(PG_FSS.W)XR)OQ/JIEc>RK;$
`endprotected


  /** Transaction that holds ownership of snoop data channel */
  protected svt_axi_master_snoop_transaction snoop_data_chan_owner;

  /** Transaction that holds ownership of snoop response channel */
  protected svt_axi_master_snoop_transaction snoop_resp_chan_owner;

  /** Current owner for driving WACK*/
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE wack_owner;

  /** Current owner for driving RACK*/
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE rack_owner;

  // NC gives this error for these declarations (not currently supported)
  // Associative array uses an element data type that is not currently supported [SystemVerilog]
`ifndef INCA
  /** Associative array of the send_write_addr process indexed by
    * the transaction handle */ 
  protected process receive_snoop_addr_proc_q [svt_axi_master_snoop_transaction];

  /** Associative array of the send_write_data process indexed by
    * the transaction handle */ 
  protected process send_snoop_data_proc_q [svt_axi_master_snoop_transaction];

  /** Associative array of the receive_write_resp process indexed by
    * the transaction handle */ 
  protected process send_snoop_resp_proc_q[svt_axi_master_snoop_transaction];
`endif

  /** Event that indicates that the receive_snoop_addr process has kicked off */
  protected event ev_snoop_addr_started;

  /** Event that indicates that the send_snoop_data process has kicked off */
  protected event ev_snoop_data_started;

  /** Event that indicates that the send_snoop_resp process has kicked off */
  protected event ev_snoop_resp_started;

  /** Event that indicates that dvm complete has arrived on snoop channel for dvm sync on read channel */
  protected event ev_snoop_dvm_complete_received;

  /** Event that indicates that dvm complete has arrived on read channel for dvm sync on snoop channel */
  protected event ev_dvm_complete_received;

  /** Reference to the object corresponding to the last sample of ACVALID */ 
  protected svt_axi_master_snoop_transaction curr_snoop_addr_xact;

  /**
    * Semaphore that controls access to logic that drives acready when
    * the default value of acready is 1. Look for comments in 
    * the task drive_acready for a detailed description
    */
  protected semaphore acready_sema;

  /** Master exclusive monitor that monitors the snoop transactions corresponding to store transaction from other masters */  
  protected bit excl_mon [*];

  /** Flag to avoid same exclusive transaction getting processed again */
  protected bit excl_xact_processed [svt_axi_transaction];

  /** Semaphore that controls access to master excluisve monitor */
  protected semaphore excl_mon_sem;
  
  /** Semaphore that controls the processing of coherent exclusive transaction one at a time */
  protected semaphore excl_access_sem;


  /** Array to hold outstanding barrier pair transactions */
  svt_axi_barrier_pair_transaction barrier_pair_xact[$];

  /**
    * Snoop transaction that has not yet been added to queue. This
    * happens when the received snoop address matches an outstanding
    * WRITEBACK/WRITECLEAN/EVICT. The snoop is not sent out to the user
    * until the WRITEBACK/WRITECLEAN/EVICT is complete.
    */
  protected svt_axi_master_snoop_transaction suspended_snoop_xacts[$];

  protected int num_pending_dvm_completes = 0;

  //**************** AXI4 STREAM RELATED MEMBERS ******************
  protected svt_axi_transaction data_stream_owner;
  // ****************************************************************************


  // ****************************************************************************
  // Local MEMBERS
  // ****************************************************************************
  protected bit suspend_arvalid = 0;
  protected bit suspend_awvalid = 0;
  protected bit suspend_wvalid  = 0;
  protected bit suspend_bready  = 0;
  protected bit suspend_rready  = 0;

  /** Master Transaction */
  protected `SVT_AXI_MASTER_TRANSACTION_TYPE global_parity_xact;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter, svt_axi_master driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter OVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter, svt_axi_master driver);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_axi_master xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** 
    * Adds the transaction to the internal queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task add_to_master_active(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Adds the transaction to an internal queue of transactions
    * got from channel, but not yet added to queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task add_to_master_current_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Adds the transaction to an internal queue of transactions
    * got from channel, but not yet added to queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    * Checks for ongoing snoop before adding. Internally calls add_to_master_current_queue
    */
  extern virtual task add_to_master_current_queue_post_snoop_check(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Adds the transaction to an internal queue of transactions
    * got from channel, when current transaction ID is matching with
    * active_xact_queue transaction ID.
    */
  extern virtual function bit  add_xact_with_same_id_to_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  unused_ids_by_active_master_transaction);

  /** 
    * Adds the transaction to read_xact_buffer or write_xact_buffer 
    * depending on whether its a read or write transaction. 
    */
  extern virtual task add_to_master_buffer(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  /** 
    * Adds the transaction to the active queue. 
    * Blocks when the  number of outstanding transactions is
    * the configured max. value.
    */
  extern virtual task load_active_from_master_buffer ();


  /**Checks for exclusive read transaction and pushes the transaction into exclusive read queue */
  extern virtual function void check_exclusive_read_transactions(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**Checks for exclusive write transaction and compares the transaction from exclusive read queue */
  extern virtual function void check_exclusive_write_transactions(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  
  /** Starts the processes of a transaction based on xact_type */
  extern virtual task start_transaction_process(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Removes transaction xact from the internal queue.  */
  extern virtual task remove_from_active(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit silent=0);

  /** Removes transaction xact from internal queue of xacts got from channel but not added to active queue.  */
  extern virtual task remove_from_master_current_queue(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives read address channel signals */
  extern virtual task send_read_addr(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Receives read data for a transaction */
  extern virtual task receive_read_data(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Receives read data for a transaction */
  extern virtual task receive_read_chunk_data(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives write address channel signals. */
  extern virtual task send_write_addr(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives write data channel signals */
  extern virtual task send_write_data(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Receives write response channel signals. */
  extern virtual task receive_write_resp(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to the read address channel for this transactions*/
  extern virtual task get_read_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Waits for previous write transaction last data beat handshake*/
  extern virtual task wait_for_prev_last_write_data_handshake(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Waits for previous read transaction last data beat handshake*/
  extern virtual task wait_for_prev_last_read_data_handshake(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to the write address channel for this transactions*/
  extern virtual task get_write_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to the address channel (merged) for this transactions*/
  extern virtual task get_serial_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to the write data channel for this transactions*/
  extern virtual task get_write_data_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Releases lock of read adress channel. Decides which transaction should
    * be the next owner of the read address channel.
    */
  extern virtual task release_read_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** 
    * Releases lock of write adress channel. Decides which transaction should
    * be the next owner of the write address channel.
    */
  extern virtual task release_write_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** 
    * Releases lock of adress channel (merged). Decides which transaction should
    * be the next owner of the address channel.
    */
  extern virtual task release_serial_addr_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** 
    * Releases lock of write data channel. Decides which transaction should
    * be the next owner of the write data channel.
    */
  extern virtual task release_write_data_chan_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /**
    * Returns the number of beats based on the current
    * interleave and the the random_interleave_array
    */
  extern virtual function int get_number_of_transfers(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, int curr_intrlv);

  /*
   * Waits until bvalid with the id of this transaction is received
   */
  extern virtual task wait_for_bresp(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /*
   * Tracks bresp timeout for a write transaction 
   */
  extern virtual task track_wdata_bresp_timeout(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /*
   * Waits for the assertion of rvalid and associates it with a
   * transaction
   */
  extern virtual task wait_for_rvalid(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Waits for rdata */
  extern virtual task wait_for_rdata(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /*
   * Returns the number of outstanding transactions
   */
  extern virtual function int get_number_of_outstanding_master_transactions(bit silent = 1, output `SVT_AXI_MASTER_TRANSACTION_TYPE actvQ[$]);

  /** Returns the number of auto-generated transactions. */
  extern virtual function int get_number_auto_generated_xacts();

  /** Returns the number of dropped coherent transactions. */
  extern virtual function int get_number_dropped_coherent_xacts();

  /** Updates the ace counters for auto-generated and dropped coherent transactions. */
  extern virtual function void update_ace_counters(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /* Checks if current transaction is allowed to proceed based on ID overlap rule with outstanding transactions */
  extern virtual task check_id_overlap_rule_and_wait_if_not_allowed(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Returns the number of READ transcations that have started  and in 
    * active queue
    */
  extern virtual function int get_num_started_read_xacts();
  
 /** 
    * Returns the number of WRITE transcations that have started  and in 
    * active queue
    */
  extern virtual function int get_num_started_write_xacts();

`ifdef SVT_ACE5_ENABLE
 /** 
    * Returns the number of WRITE transcations that have started  and in 
    * active queue
    */
  extern virtual function int get_num_started_atomic_xacts ();
`endif

  /*
   * Returns the delay to be executed by the address channel 
   */
  extern virtual function int get_addr_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);
  
  /*
   * Returns the delay to be executed by the address channel 
   */
  extern virtual function int get_dvm_addr_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Timer for DVM Complete for DVM Sync received on read/snoop channel */
  extern virtual task track_snoop_dvm_complete_timeout(`SVT_AXI_MASTER_TRANSACTION_TYPE xact); 
  /*
   * Returns the delay to be executed by the data channel.
   */
  extern virtual function int get_write_data_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, int addr_event_cycle);

  /*
   * Returns the delay to be executed by the data stream channel.
   */
  extern virtual function int get_data_stream_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, int addr_event_cycle);

  /** Advances clock by #num_clocks */
  extern virtual task advance_clock(int num_clocks);

  /** Steps one clock*/
  extern virtual task step_monitor_clock();

  /** Drives the read address channel signals on the physical pins */
  extern virtual task drive_read_addr_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the read address channel signals on the physical pins */
  extern virtual task drive_read_addr_chan_signals_without_awakeup(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Deasserts read address channel signals*/
  extern virtual task deassert_read_addr_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** Waits until arready is received */
  extern virtual task wait_for_arready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the write address channel signals on the physical pins */
  extern virtual task drive_write_addr_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the write address channel signals on the physical pins */
  extern virtual task drive_write_addr_chan_signals_without_awakeup(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Assign the addr awakeup assertion cycle to transaction*/
  extern virtual task addr_wakeup_assertion(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the awakeup signal during idle time period of addr channel */
  extern virtual task toggle_awakeup_signals_during_idle_channel( );

  /** Deasserts write address channel signals*/
  extern virtual task deassert_write_addr_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** Waits until awready is received */
  extern virtual task wait_for_awready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the write data channel signals on the physical pins */
  extern virtual task drive_write_data_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the write data channel signals on the physical pins */
  extern virtual task drive_write_data_chan_signals_without_awakeup(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Deasserts write data channel signals*/
  extern virtual task deassert_write_data_chan_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** Waits until wready is received */
  extern virtual task wait_for_wready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit output_timed_out_);

  /** Waits until bready is received */
  extern virtual task drive_bready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Toggles RREADY signal when the read data channel is IDLE */
  extern virtual task toggle_bready_during_idle(svt_axi_transaction xact, output bit is_valid_accepted);

  /** Waits until rready is received */
  extern virtual task drive_rready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Wait for suspended signal from being driven. 
    * Before the driver attempts to drive these signals, it will check if it has been suspended. 
    * If so, it will wait until the suspended signal has been resumed with a call to resume_signal. 
    * This is supported only for valid and ready signals. 
    * It is supported for ready signals only when the corresponding default is low.
    */
  extern virtual task wait_for_suspend_signal_resume(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, string signal_name="");

  /** Toggles RREADY signal when the read data channel is IDLE */
  extern virtual task toggle_rready_during_idle(svt_axi_transaction xact, int curr_beat, output bit is_valid_accepted);

  /** Drives the read data channel debug ports on the physical pins */
  extern virtual task drive_read_data_chan_debug_port(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Drives the write resp channel debug ports on the physical pins */
  extern virtual task drive_write_resp_chan_debug_port(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Sets internal variables used by this class based on the config */
  extern virtual function void set_internal_variables(svt_axi_port_configuration cfg);

  /** Samples signals from the physical pins and does signal level checks */
  extern virtual task sample();

  /** Samples the reset signal */
  extern virtual task sample_reset();
 /**samples initial reset async*/
  extern virtual task sample_reset_async();
  extern virtual function void detect_initial_reset();
  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Initializes master I/F output signals to 0 at 0 simulation time */
  extern virtual task async_init_signals();

  /** Drive default values for master signals during asynchronous reset **/
  extern virtual task default_signal_values_async_reset(); 

  /** Initializes signals */
  extern virtual task initialize_signals();

  /** Drive the idle values after initial reset */
  extern virtual task drive_idle_val_initial_reset();

  /** Waits until any transaction ends */
  extern virtual task wait_for_any_transaction_ended();

  /** Sets the configuration */
  extern virtual function void set_cfg(svt_axi_port_configuration cfg);

  /** Waits until a valid or handshake takes place on any channel*/
  extern virtual task wait_for_bus_activity();

  /** Checks if the handle given matches any of those of the active transactions. */
  extern virtual function void check_xact_handle(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Utility function to construct timers */
  extern virtual function void create_timers();

  /** Creates dynamic arrays of non-rand variables of xact based
    * on burst_length. This is done in the driver because here 
    * we can ensure that the arrays are created 
    * whether a transction is randomized or not
    */
  extern virtual function void safe_set_burst_dimensions(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Creates the transaction inactivity timer
    */
  extern virtual function svt_timer create_xact_inactivity_timer();

  /**
    * Returns 1 if the specified error_kind is there in transaction, else returns 0 
    */
  extern virtual function bit has_axi_exception(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, svt_axi_transaction_exception::error_kind_enum error_kind); 

  /**
    * Drive invalid values to signals in case an exception is injected 
    */
//  extern virtual function void drive_axi_exception(svt_axi_master_transaction xact, svt_axi_transaction_exception::error_kind_enum error_kind);  

  // ---------------------------------------------------------------------------
  // LOCKED XACT PROCESSING RELATED METHODS 
  // ---------------------------------------------------------------------------
  /** Detects a new locked sequeunce */
  extern virtual task is_new_locked_sequence(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_new_sequence);

  /** Checks if the received transaction is part of the current locked sequence if any */
  extern virtual task is_xact_in_current_locked_sequence(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_in_current_locked_seq);

  /** Checks if the received transaction is a valid locked sequeunce transaction */
  extern virtual task is_valid_locked_sequence_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_valid_xact);


  // ---------------------------------------------------------------------------
  // SNOOP PROCESSING RELATED METHODS 
  // ---------------------------------------------------------------------------
  /** Adds a new snoop transaction to the queue */
  extern virtual task add_to_master_snoop_active(svt_axi_master_snoop_transaction xact);

  /** Removes a snoop transaction from the queue */
  extern virtual task remove_snoop_xact_from_active(svt_axi_master_snoop_transaction xact);

  /** Receives snoop address */
  extern virtual task receive_snoop_addr(svt_axi_master_snoop_transaction xact);

  /** Sends snoop data */
  extern virtual task send_snoop_data(svt_axi_master_snoop_transaction xact);

  /** Sends snoop response */
  extern virtual task send_snoop_resp(svt_axi_master_snoop_transaction xact);

  /** Drives the ACREADY signal based on the delay */ 
  extern virtual task drive_acready(svt_axi_master_snoop_transaction xact, output bit wait_for_acready_end);

  /** Gets the delay associated with snoop data transfer */
  extern virtual function integer get_snoop_data_delay(svt_axi_master_snoop_transaction xact);

  /** Drives the snoop data channel signals */
  extern virtual task drive_snoop_data_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Waits for the CDREADY signal */
  extern virtual task wait_for_cdready(svt_axi_master_snoop_transaction xact);

  /** Deasserts the snoop data channel signals */
  extern virtual task deassert_snoop_data_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Gets access to the snoop data channel for a transaction */
  extern virtual task get_snoop_data_chan_lock(svt_axi_master_snoop_transaction xact);

  /** Assigns ownership of snoop data channel to a transaction */
  extern virtual task release_snoop_data_chan_lock(svt_axi_master_snoop_transaction xact = null);

  /** Gets the delay associated with snoop response transfer */
  extern virtual function integer get_snoop_resp_delay(svt_axi_master_snoop_transaction xact);

  /** Drives the snoop response channel signals */
  extern virtual task drive_snoop_resp_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Waits for the CRREADY signal */
  extern virtual task wait_for_crready(svt_axi_master_snoop_transaction xact);

  /** Deasserts the snoop response channel signals */
  extern virtual task deassert_snoop_resp_chan_signals(svt_axi_master_snoop_transaction xact);

  /** Gets access to the snoop response channel for a transaction */
  extern virtual task get_snoop_resp_chan_lock(svt_axi_master_snoop_transaction xact);

  /** Assigns ownership of snoop response channel to a transaction */
  extern virtual task release_snoop_resp_chan_lock(svt_axi_master_snoop_transaction xact = null);

  /** Samples snoop address channel and assigns values to snoop transaction object */
  extern virtual task process_snoop_addr_channel(ref int acvalid_to_acready_delay, output svt_axi_master_snoop_transaction new_snoop_xact);

  /** 
    * Waits for a new snoop transaction. The monitor uses this task to get a 
    * handle to the new snoop transaction.
    */ 
  extern virtual task wait_for_acvalid(output svt_axi_master_snoop_transaction xact);

  /**
    * Tracks suspended snoop xacts and triggers events when they are ready
    * to be added to the queue
    */
  extern virtual task track_suspended_snoop_xacts();

  /** Gets access to drive WACK*/
  extern virtual task get_wack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Gets access to drive RACK*/
  extern virtual task get_rack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Releases lock of WACK. Decides which transaction should
    * be the next owner to drive WACK.
    */
  extern virtual task release_wack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** 
    * Releases lock of RACK. Decides which transaction should
    * be the next owner to drive RACK.
    */
  extern virtual task release_rack_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  /** Drives debug port signals for snoop data channel */
  extern virtual task drive_snoop_data_chan_debug_port(svt_axi_master_snoop_transaction xact);

  /** Drives debug port signals for snoop response channel */
  extern virtual task drive_snoop_resp_chan_debug_port(svt_axi_master_snoop_transaction xact);
  
  /** Drives debug port signals for snoop address channel */
  extern virtual task drive_snoop_addr_chan_debug_port(svt_axi_master_snoop_transaction xact);

  /** Checks coherent transaction. If data is available in cache it is retreived */ 
  extern virtual task process_coherent_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Reserves an index in cache for allocation of this transaction */ 
  extern virtual task reserve_cache_allocation(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output `SVT_AXI_MASTER_TRANSACTION_TYPE lru_xact);

  /** Writes data into cache */
  extern virtual task write_into_cache(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual function void get_end_cache_state_and_data(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,
                                                    output bit update_cache,
                                                    output bit update_only_status,
                                                    output int is_unique,
                                                    output int is_clean,
                                                    output bit use_cache_write_data
                                                  );

  /** Assigns initial_snoop_cache_line_state based on cache state */
  extern virtual task assign_snoop_xact_cache_line_state(svt_axi_master_snoop_transaction snoop_xact, string kind);

  /** Assigns initial and final cache line states in xact based on cache state */
  extern virtual task assign_coh_xact_cache_line_state(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, string kind);

  /** 
    * Updates the cache based on snoop response assigned by user after 
    * receiving a snoop transaction from the input channel 
    */
  extern virtual task post_snoop_cache_update(svt_axi_master_snoop_transaction snoop_xact);

  /** Waits for post_snoop_cache_update() method to complete if any activity
    * is observed on the SNOOP channel */
  extern virtual task is_post_snoop_cache_update_done(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit check_outstanding_queue= 0);  

  /** Does the necessary processing to end a transaction */
  extern virtual task end_transaction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit is_removed=0);

  /** returns the delay for RACK signal */
  extern virtual function int get_rack_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** returns the delay for WACK signal */
  extern virtual function int get_wack_delay(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Checks if a transaction can be given the lock from the
    * perspective of a barrier
    */
  extern virtual function void check_chan_lock_for_barrier(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit give_lock);

  /**
    * Checks if a transaction can be given the lock from the
    * perspective of transaction ID
    * 
    */
  extern virtual function void check_chan_lock_for_xact_id(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit give_lock);

  /*
   * Checks if a transaction can be given the lock from the
   * perspective of cache maintenance transactions
   */
  extern virtual function void check_addr_chan_lock_for_cache_maintenance (
                         `SVT_AXI_MASTER_TRANSACTION_TYPE xact, 
                         bit check_cache_maintenance,
                         bit check_memory_update,
                         ref bit cache_maintenance_in_progress,
                         ref bit memory_update_in_progress
                       );

  /** Checks that a transaction can be given the lock taking requirements 
    * for snoop filter into consideration */
  extern virtual function void check_read_addr_chan_lock_for_snoop_filter(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, ref bit snoop_filter_give_lock);

  /** Checks if there is a snoop to the same cache line addressed by xact */
  extern virtual function svt_axi_master_snoop_transaction check_snoop_to_same_cache_line(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);
  
  /** Gets the handle of a snoop transaction to the same address as that of a WRITEUNIQUE or WRITELINEUNIQUE transaction */
  extern virtual function svt_axi_master_snoop_transaction get_snoop_to_same_addr_during_wu_wlu(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** Checks if there is a resp to the same cache line addressed by xact */
  extern virtual function `SVT_AXI_MASTER_TRANSACTION_TYPE check_resp_to_same_cache_line(svt_axi_master_snoop_transaction xact, output bit is_resp_to_same_cache_line);

  extern virtual task drive_wack(logic val);

  extern virtual task drive_rack(logic val);

  extern virtual task perform_cache_update(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_rack_and_update_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_wack_and_update_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_read_addr_chan_coherent_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task deassert_read_addr_chan_coherent_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task drive_write_addr_chan_coherent_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task deassert_write_addr_chan_coherent_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task process_ace_reset();

  extern virtual task pre_process_coherent_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,
                                                ref `SVT_AXI_MASTER_TRANSACTION_TYPE memory_update_xact,
                                                ref bit drop_barrier);

  extern virtual task wait_for_write_xacts_to_same_cache_line(svt_axi_master_snoop_transaction new_snoop_xact);

  extern virtual task wait_for_xacts_to_same_cache_line_to_end(`SVT_AXI_MASTER_TRANSACTION_TYPE xact,output bit is_xact_outstanding);

  extern virtual task get_coherent_write_to_same_cache_line(svt_axi_master_snoop_transaction snoop_xact,output `SVT_AXI_MASTER_TRANSACTION_TYPE coh_write_to_same_cache_line);

  extern virtual task trigger_new_snoop_addr_chan_activity_event(svt_axi_master_snoop_transaction snoop_xact);

  extern virtual task wait_for_cache_update_post_curr_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit is_snoop_to_same_cache_line);

  extern virtual task check_chan_lock_for_outstanding_snoop(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, output bit b_has_outstanding_snoop);

  extern virtual task update_current_snoop_xact_handle(svt_axi_master_snoop_transaction snoop_xact);

  extern virtual task check_for_writeunique_writelineunique_restriction(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  extern virtual task include_dirty_data_into_xact(svt_axi_cache axi_cache, `SVT_AXI_MASTER_TRANSACTION_TYPE parent_xact, `SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit original_txn=0);

  // send de-allocating transaction (CLEANINVALID) when cacheline doesn't get updated due to error response
  extern virtual task check_and_remove_cacheline_from_snoop_filter(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  //**************** AXI4 STREAM RELATED METHODS ******************
  // Main task that controls transmit of data stream
  extern virtual task send_data_stream(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  // Gets the data stream lock for this transaction.
  extern virtual task get_data_stream_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  // Releases access to data stream lock and assigns it to a new transaction
  extern virtual task release_data_stream_lock(`SVT_AXI_MASTER_TRANSACTION_TYPE xact = null);

  // Waits for tready to be asserted
  extern virtual task wait_for_tready(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  // Drives data stream signals
  extern virtual task drive_data_stream_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  // Assigns default values to data stream signals
  extern task deassert_data_stream_signals(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  `ifdef SVT_AXI_QVN_ENABLE
  //
  // Method to drive token request signals for corresponding AXI channels - Read Address, Write Address and Write Data.
  // It also uses address channel names appended with QOS to drive only QOS signals for respective token request when 
  // it wants to upgrade QOS value waiting for token request grant from slave.
  // Depending on the channel_name == "READ_ADDR" or "WRITE_ADDR" this method will use either VAWVALIDVNx or VARVALIDVNx
  // and corresponding QOS signal i.e. VAWQOSVNx or VARQOSVNx
  // if channel_name == "WRITE_DATA" then VWVALIDVNx signal will be driven.
  // if channel_name == "READ_ADDR_QOS" or "WRITE_ADDR_QOS" this method will drive either VAWQOSVNx or VARQOSVNx signal 
  // only, in order to upgrade QOS values.
  // Virtual Network ID (vnet_id) passed to this method will determine which *VNx" signal will be used i.e. if vnet_id=2
  // then "*VN2" signals will be used. It uses axi_master_cb clocking block of svt_axi_master_if interface.
  // It is the responsibility of the caller to pass correct channel name and transaction handle to request token on correct
  // channel and pass correct QOS value. In order to re-use this method to de-assert token request signals, it should have 
  // another argument "bit valid" which will be used to driver valid signals for requesting token. While requesting token 
  // caller will pass valid=1 and to de-assert caller will pass valid=0"
  //
  // Drive QVN signals for respective AXI Channels - Read-Address, Write-Address, Write-Data
  //
  extern task qvn_drive_token_request_signals(int vnet_id, int qos_value, string channel_str, bit valid=1'b1);

  // Once master has driven token request it waits for the request to be granted by slave. When slave asserts ready for corresponding token request to the respective channel that marks the end of token request. At this point master will either de-assert valid signals for that token request or drive another token request without inserting any delay.

  // Drive QVN signals for respective AXI Channels - Read-Address, Write-Address, Write-Data
  extern task qvn_deassert_token_request_signals(int vnet_id, string channel_str);

  //
  // Once master has driven token request, it waits for the request to be granted by slave. When slave asserts ready for 
  // corresponding token request to the respective channel that marks the end of token request. For this purpose, master 
  // uses following method to sample token request ready signal driven by slave.
  // Depending on channel name passed through "channel_str" and Virtual Network number passed through "vnet_id" it chooses
  // which signal it needs to drive. It uses axi_master_cb clocking block of svt_axi_master_if interface.
  // Channels supported:: "READ_ADDR" => Read Address channel, "WRITE_ADDR" => Write Address channel, "WRITE_DATA" => Write Data Channel
  // Example: if vnet_id = 2 and channel_str = "WRITE_DATA" then it will sample "driver_mp.axi_master_cb.vwreadyvn2"
  //
  // Samples QVN Ready signal for a Virtual Network for respective AXI Channels - Read-Address, Write-Address, Write-Data and returns sampled signal value.
  //
  extern function bit qvn_sample_token_request_ready(int vnet_id, string channel_str);

  //
  // Requests for new Token in specified channel for the Virtual Network to which current Transaction is issued.
  // While driving token request, it passes QOS value from qvn_qos_value_queue of current transaction based on the
  // token request number passed to this method. If the request is made first time for the current transaction, based
  // on the token request number, then it also tries to upgrade QOS value it has already driven as per the transaction
  // configuration of qvn_qos_upgrade_delay_queue and qvn_qos_upgrade_value_queue. 
  // For QOS upgrade it uses qvn_qos_upgrade_delay queue to determine when to upgrade QOS value. So, after driving QVN
  // token request it samples corresponding token request ready signal (asserted by slave). If it is asserted then it
  // returns from the task by de-asserting token request valid signal marking end of token request.
  // If ready signal is de-asserted then it keeps waiting and for each clock cycle of the axi_master_cb clocking block
  // it tracks how many cycles it has been waiting. If it waited for first entry of the qvn_qos_upgrade_delay_queue then
  // master will upgrade its QOS value keeping track of which delay value it has used. If it so happens that master is
  // still waiting for token request grant and it reaches next QOS upgrade delay specified, then at that time it will 
  // use next entry i.e. qvn_qos_upgrade_value_queue[1] to upgrade QOS again and this process will repeat until token 
  // request is granted by slave or number of QOS upgrade reaches to qvn_num_qos_upgrade value, whichever is earlier.
  //   Since, multiple processes will call this method in their own order so, it makes use of single-key semaphore of
  // the token-pool of same virtual network for which request is being made. Based on the channel READ_ADDR, WRITE_ADDR
  // or WRITE_DATA and virtual network id of current transaction, it chooses which token pool to use.
  //
  // if a master shares same Virtual Network with another one or if slave uses shared token for different masters then
  // there is a possibility that, a master can issue multiple token requests and once granted those tokens remain unused
  // reserving system resources and in turn blocking other masters. To avoid this, it checks if Maximum number of Unused Token
  // reached configured number of maximum limit. In that case, it waits until number of unused token goes below the maximum limit.
  // This protects a system from one master reserving large number of resources in one time.
  //
  extern task qvn_request_token(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, string channel_str, int token_req_number=0);

  //
  // This task is primarily responsible for managing issuance of token request based on the transaction handle information 
  // sent by processes - send_read_address, send_write_address and send_write_data. Once it is launched by the master driver
  // at the beginning of simulation it remains alive for rest of the simulation as a non-blocking free-running thread.
  //    At first, it checks if QVN is enabled for this master. If not enabled then it terminates the task without doing anything 
  // further. If QVN is enabled then first, it initiallizes token-pool of each supported Virtual Network in each AXI Channel 
  // (AR, AW, W) with configured value of pre-allocated token number of respective channels (qvn_num_ar_pre_allocated_token_vn, 
  // qvn_num_aw_pre_allocated_token_vn, qvn_num_w_pre_allocated_token_vn).
  //    Then it spawns of three parallel non-blocking threads to take care of token requests for read-address, write-address and
  // write-data channel. Each thread is free-running and gets blocked by axi_master_transaction mailbox of respective channel.
  // So, at the start of each thread it checks if any transaction handle is available in its mailbox. It waits if mailbox is empty.
  // If a transaction is available in the mailbox then it pops out that handle and checks number of token available in that
  // channel for the Virtual Network the transaction was issued to. 
  //    If it finds that no token is available and no token request has been set in the transaction then for address channel it 
  // forces 1 token to be requested. For Data channel it checks how many token is required to make full data transfer for that 
  // transaction. If number of available token and number of token request set in the received transaction is less than the number
  // of token is required then it forces additional tokens to be requested to make up that difference.
  //    However, if number of available token and number of token request set in the transaction is equal to or more than required
  // token then it simply requests as per the token request number set in the transaction for address or data channel.
  //    NOTE: since write data channel requires token for each beat of data transfer, send_write_data process passes transaction handle
  // to this method via write_data_mailbox multiple times for each transfer. "qvn_num_data_token_request" set in transaction handle
  // is considered to send token request only for the first data-beat. For subsequent data-beat transfer this method only checks if
  // sufficient tokens are available or not. If not available only then it requests for new token. For first data-beat, even if
  // more tokens are available, it goes ahead and requests token as set in transaction handle.
  //    Since these processes request token in different order, discreetly one at a time or multiple requests together, these requests
  // are controlled by token_request semaphore of each virtual network token pool of corresponding channel. So, even if multiple
  // token request threads are spawned-off these are blocked by the above sempahore and only one token request gets access to the
  // bus for that virtual network of the corresponding channel. Once this request is complete one among other pending token request
  // gets unblocked and starts driving token request on the bus.
  //
  extern virtual task qvn_process_token_request();

  //
  // Each process that performs a transfer on Axi Read Address, Write Address or Write Data channel, needs at least one token for each
  // transfer. So, send_read_addr, send_write_addr and send_write_data each of this method needs to wait for at least one token to be
  // available for respective channel and the virtual network to which it intends to send current transaction. For this purpose, this 
  // method provides a common implementation for above three tasks to wait for token before proceeding with a transfer.
  //    It needs argument "enable" which indicates QVN feature is enabled for this master and current transaction is not of BARRIER type
  // If enabled then it needs to checks for token availability but, before that, it passes current transaction handle to 
  // "qvn_process_token_request" task so that, number of token requests in current transaction are driven to respective VN and axi channel
  // or in case of non-availability of token, required number of token requests can be carried out. Corresponding mailbox handle passed
  // through "mbox" argument is used for this purpose.
  // After this, it checks available token number through corresponding qvn token pool passed through 'token' argument. If token is
  // available it proceeds otherwise waits until a token is available by checking it through 'token' handle at every clock cycle. Once a
  // token is available it stops a corresponding timer which was started before each of the above task started to wait for token availability
  // i.e. called "qvn_wait_for_token" and terminates indicating a transfer on current chanel and virtual network can proceed.
  //
  extern virtual task qvn_wait_for_token(bit enable, axi_master_transaction_mailbox mbox, `SVT_AXI_MASTER_TRANSACTION_TYPE xact, qvn_token_pool token, svt_timer timer);
  `endif

  /**
    * This method is used to get list of all IDs which are currently under use by outstanding transactions. However, user
    * can choose the type of outstanding transactions this method should consider while extracting ID of active transactions.
    * "mode" and "rw_type" arguments should be used for this purpose.
    *
    * It returns '1' if total number of unique IDs currently used by active transactions, is less than all possible ID that can
    * be used by an AXI transaction. This helps in determining whether randomizing ID field of a new transaction which should
    * not be part of the all the IDs currently in use, is possible or not.
    * 
    * @param mode Type of outstanding transactions this method should consider while extracting ID of active transactions.
    *             Currently it supports following modes (defined as string) ::
    *               - "non_dvm_non_barrier" => all transactions which are neither DVM nor Barrier  (default)
    *               - "non_dvm"             => all transactions which are not DVM 
    *               - "non_barrier"         => all transactions which are not Barrier 
    *               - "dvm"                 => all transactions which are of DVM type 
    *               - "barrier"             => all transactions which are of Barrier type
    *               - "dvm_barrier"         => all transactions which are either DVM or Barrier type
    *               - Note: if "rw_type" is set to '0' then only read channel transactions will be considered for non-dvm
    *                       and non-barrier type
    *               .
    * 
    * @param rw_type Indicates which channel id width should be considered.
    *               - ' 0 ' => only read channel id width and transactions should be used
    *               - ' 1 ' => only write channel id width and transactions should be used
    *               - '-1 ' => common or either of read or write channel id width and transactions are used
    *               .
    * 
    * @param use_min_width If set to '1', minimum of read and write channel id width should be used otherwise maximum.
    *               This is applicable only if "rw_type == -1" i.e. no particular channel id width is specified.
    * 
    * @param silent Suppresses debug messages from this method if set to '1'
    */
  extern virtual function bit get_ids_used_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_dvm_non_barrier", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);
  extern virtual function bit get_ids_unused_by_active_master_transactions(output bit[`SVT_AXI_MAX_ID_WIDTH-1:0] id_list[$], input string mode="non_device_or_non_dvm", input int rw_type=-1, input bit use_min_width=1, input bit silent=1);

  /**
    * This method is used to update current transaction handle (argument xact) with overlapped transactions which are
    * accessing same cacheline and have not completed i.e. currently active.
    *
    * @param xact Indicates current transaction handle that needs to be updated with overlapped transaction
    *
    */
  extern virtual task set_overlapped_xacts(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /**
    * Method that auto generates DVM complete transactions
    *
    * @ param snoop_xact Handle to the DVM SYNC transaction for which DVM complete must be generated
    * @ param phase UVM phase from which this task is called
    */
`ifdef SVT_VMM_TECHNOLOGY
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact);
`else
  extern virtual task send_auto_gen_dvm_complete(svt_axi_master_snoop_transaction snoop_xact, svt_phase phase);
`endif
 
  /** Returns if all Snoop DVM COMPLETEs are received for coherent DVM Sync sent */
  extern virtual function bit is_dvm_snoop_sync_complete_done();

  /** Wait for conditions for DVM */
  extern virtual task check_and_wait_for_dvm_complete_conditions(svt_axi_transaction xact);

  /** checks if reset asserted and then aborts transaction */
  extern virtual task check_reset_and_abort_xact(`SVT_AXI_MASTER_TRANSACTION_TYPE xact, bit give_seq_resp=1, bit check_unstarted=1, bit wait_for_reset=0);

  /** waits for transaction which has been blocked by other transactions more than `SVT_AXI_NUM_BLOCKED_XACTS_ALLOWED number of times.
    * It wait for those blocked transaction to finish. This will avoid starvation of some type of transactions and will provide
    * more fair chance to all the transactions to proceed
    */
  extern virtual task wait_for_severly_blocked_transactions_to_make_progress(`SVT_AXI_MASTER_TRANSACTION_TYPE xact=null);

  /** waits until VIP is out of reset */
  extern virtual task wait_for_out_of_reset(int mode = 0);

  /** waits until VIP is in reset */
  extern virtual task wait_for_reset(int mode = 0);

  /**
    * If an incoming snoop changes cacheline state, we need to reevaluate if a memory update transaction
    * can be sent out. This task does that
    */
  extern virtual task check_pre_xact_start_conditions_for_mem_update_xacts(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** task to provide sequence item processed response from the driver to the sequencer */
  extern virtual task sequencer_put_response(`SVT_AXI_MASTER_TRANSACTION_TYPE xact);

  /** 
    * Suspends signal from being driven based on signal_name value. 
    * That is, the signal will be driven low and will wait for a call to resume_signal 
    * before it is driven high.
    * Following are supported values for signal_name
    * - awvalid     - suspend the signal awvalid 
    * - wvalid      - suspend the signal wvalid 
    * - bready      - suspend the signal bready 
    * - arvalid     - suspend the signal arvalid  
    * - rready      - suspend the signal rready 
    * - all_signals - suspend awvalid, wvalid, bready, arvalid, rready signals   
    * .
    */
  extern virtual task suspend_signal(string signal_name = "");

  /** 
    * Resumes signal after being suspended based on signal_name value. 
    * That is, the suspended signal will be resumed back and respective signals  
    * will be driven high.
    * Following are supported values for signal_name
    * - awvalid     - resume the signal awvalid 
    * - wvalid      - resume the signal wvalid 
    * - bready      - resume the signal bready 
    * - arvalid     - resume the signal arvalid  
    * - rready      - resume the signal rready 
    * - all_signals - resume awvalid, wvalid, bready, arvalid, rready signals   
    * .
    */
  extern virtual task resume_signal(string signal_name = "");

  /** task to sample parity check signals and calculate respective signal parity values for parity check comparision */
  extern virtual task sample_and_check_parity_check_signal();

  //***************************************************************
`ifndef SVT_AXI_DISABLE_SYSTEM_ENV_ACCESS_FROM_AGENT
  extern virtual function void set_system_env();
`endif

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
HV:UI:U^AHdG\R\-\e7N=RA5IMJ4_KB^1_0#0VbSXXdVXfRcbKVG6)9\.+6&KO_C
ZJ))?5XP&>.8?Q=#)b+=?6PK8Dd632]F_4Yg\)0,I5\KJE<VM73VS9GP(b1?1BPV
f0b<.52W?AJGbXLIGKE(-2(Yf98/ZH8eNA4VWf)0[-TDXQ?IV+>1_-&V\[F72g:A
R(?U6>WM?;cL9M^8N@[LXJ.a<H18JMdY:(<e9\[8D9P<ZT3]LHYA=3]cSe1Nb>Y1
<0C+3;^E0gQ,\<Z>SR0;A1RO[a4D8B&;Ug;<8Idge?&F>)1CII9O53\aDF[=4;aI
a1#:_4YIH6JVgDH6@J<3@S<XF4ReV[3GE?0@#3[_fJ<cN/YV43R>B:cFfgLA>c93
9W?:#eCCGI]+HB8?dLG6&0/A6cWMdX3fJ#@LNI/G>;@-@Acd3S4;WN^(WWPKU[=#
a0f7/?FcC7#O)gKGMd+H>M.6:N:3&AJ\XV1A-?VC>9&E&VS>Lcdd_7BE1P^[V(L/
7),.:F=\NZ95A6,WIOI,1VP#d7CR9f:,]4;Bf2Idd4OfGTO1(..6G6CC08KG:QV+
^]T/Q3dN]dQH0YSfXIcR5B?BF\E>KVBPe)HZN36LCA[DCF<b>eFFV&[;X54/<K:c
>Q)T@f_#P#(LD^>aJP(((ZXF6gU_(.OVFI9IJ\K]3FHW[b30\c-K5].;7MZTR[=,
Cb;ZN)H.W]f&IFC0(63EB-@UcSa]g9R(/gg?D><+TdS1d5fMZPGG_#+@#=I;B&.<
aWONC5XN--^6#0V(T&Ng))(eH7/0Z^]2)CE+@fg15gK5JYb[a&9]=&XE3K+MFN2c
B3K#:>c9N047]fTRSUX6N;WFa,12])?gd/HaD;b++a.Z#b-1:X3^T3[<#QT<MPSQ
()QK_NHFgZ9_+H8I18<FAZ(BNKFG/#=g8)5T+Ad3R&H&3[OS7TL3D=EVLV:SKC;S
4+NETV/g]@M7A9;O,Ra5D0BBGNB:Y9V\OZc:be]9PCOA8?E#UZGf;BfaUG(<W?_(
[BGUXYNOIUTWO7V;,A6fd/V[8(/V&B0COODJ0gW[FDZYPY3C_)-<^-L.Rcb8/,Xe
O.7D?;KY(Hd(c4&=8@Y61I5GVOWaU12N.@)NK<C7^X9H)7AC^TZHNW82P&bL9ZaP
S1NJHQT_WV^WE[DJT2V8-FG,/CfE=-JS^Q;<NQH[&Mc\)QM_-K(Q3@9;-#C20\9W
[6L=]b:O#S6^<W<=)YV+[IL<(L3BVOe7AN6@J/4QJ,,^P22WSM=8a).f=>O)TL4C
JPO/U[:O(DXE=+a^/WXZH5aWFPJadd5>SRQ=^?(VA@7f1E?=?IN_W#d?2+78OT.4
38X)YLAAO;=I@PY0d61]H7I=X.R)f;O=)cAN/^adGMeb;<V46[J]26Z<_F6^>b=T
,P_U9(DS)A&IR5R\5&Z.fO]M.fe4XJCB=aGPIX\+aS,FS7X>QP[13I2G;@-YFCf;
MJ-&2&A+B5\d\5?-6=6fMX?KNU#c\=P5g^#69?4cJ2EJc>H<?B<3Q3UPDHH7&GX5
;8(]P(4E^V_Y=d]XD1g&5ZW]LfaUN(_]Cf[30ZE2,T#1X?L^IH/+d(GeNd[AOCZR
(=?RC<a4U+^c29JQgDWd[)ZDAcG<<0NBRSeL>E50SYU@HU&\ZC6Sb17MEQLKD7Z)
P\)WQ1H)Be2Wd7-G9+DD8/\=6fZAC0]2N^:Ue>I\Y]/LNbFd^dTB?M.S82U[f8Da
OISYVTU/5e-6J+U[;c6G^[MAPN#f:O<)[ePdF0\.CgDSC##+;#b8.8#NU1A&Q(I5
e4SK17O,^A?9c^I]T,3W?R/OE?65;aeNSRG-<:-3DGERc1^QaV-S9g^FD4VCUA5)
PT.L@;?_@E6CVdAg<[(0H_PNb^g+&UX6=02\XdeV7[5UR[-QL,N@44<c@:8?32#E
AE2;M0,)B53bXDc:@X.gIUY1/aAFWP#6,.C(\X_e6S9.&[]9QY/-0<aGP#?;2W0D
ZMA@cOPT;?K]cGRO2@_LHR<[O]OQ)ccgF:A#Cg#@I_3R[#O/X3VSeUD/G>QKB46d
[Y;JGS<2BfG)_7>W3Ab06f_;)FU=^EE_WfQ(;8RAE#eYb/f2>@+KKQ]bbWXJGA<c
[]E,VDb3E)(eC-K;\5S5ZGQ3/W#H93ZE:U-Q].U4090e86^=358PI?(1cK\-Y[d2
=61FWV:L@I[c:9T-df)CNX[/bG1SL-OC>8/57^?CaFFW6<Q/;KHT-W344PMdMQ<>
SB#..F)&>QZgT8O?-^_,ZCW^1A8J84,/^g:ER06bge=;M4631DB3]>:AP>Fc#PBI
[>;0#5W8,6+<JK.OKMYO&P,(gH55:IYeFX-#<+_3N^&^US,5ZcH(5b(E:?6\LfPW
:ZV<GTSTPU<X/>#(2NA>>6K9S0gHMeQK8C4Uc6bAV3F<FafAFAT3^(e8KN4VJU>c
QYOBZ7]Z5-:6/2)T)&^L&>;IU8Lc7.[#Z83/G<Q,bK#9[3:F6[]E@G;/d?CX>J#e
C4.JA_O0&^5.Pa)2;>UMCb4#RR_@S):[OfADc0+2E;.1I:P8^1VQC[c8O_.:=#F(
99FO&/135Ac8QT;04\bcA-,)6/?f4d1PDQG-Z81X^#(6:;5O=GDY4QA7LHN4=,6D
:-0gIMF(4]6]O#?JB3eT/gNWb;8Y63C9P0/7W6FC7]=D@Da?:9/Q7DFYH=WO.eWY
XaBY?E3EH9Oge(T<:fAdSVbDO<]I87)B8KC_V-3NFaX<JTXD1W?LLS)D_NdO3<NG
C0[P-GbH=f]2a+,e?c0^a#9_b\K3_14\L95;E8W+FR&,QJNB?F)+8LEPZdL4?gEU
#K:ZG65WKH&AN[C>,JA75^IC@O+_55e(CM?D\EDC9?,RQTPf^X+6[P>]-\-0<cGB
R<+46O+351#0ZA.;NZg9I@(5=-5-OC.-b^AF.TJ?5S&8M<PB0Ga1>DUWaad5]Sb2
(1S;X7(ZCMR@:23H/e>XJQBAX2YPS7<0I(-S=2;G5;D.:<_4E_]^G[Ib#d9JAX&L
62cg(5A/5-_FQ;PS[W9=2BAQa0BLCA<P>Ldc\QM,Y-2BMP4,^<APG=-U>BO-a^eJ
?1&>>Gee,\.8L.[QH-16,#>:]6ZG5-K8B3PJDe6<1.,G]DQ>U-VZ/\]e2HH;,,\:
U+0X6BQgHM@1((]>]UU.J-cVaPJP1FcXZG9BZH8G#K,:=T]+6\^PN:/G\N202R^g
2N8\.3[NTB>=T?&S,?^G-E@bKS?S<KU@bJHeSMJ(GgT/F56>b3:B7HMA#24=@BI)
b+R/HN>5K=6U.X,@0CCdU.af420cS#@Y6T[<(Z-Te0<GM0G^<d#4XGV91-_Aaca>
X#4^A<2c#E_LF9A.P5f/cQ)cH_CeKcX;[/EJVg[@=7@8gYOLUN^.2.Jf3RG;H3#3
P)X==3CX953]S+Z_)Yg.F]7[7?dgF(]AT/[\7b.IOcR5UQ/^J\P[6bLH6;cLT#^S
P9(B<NcWb;W@[IYC&NA[:Q1]3A[O/&,O1?\;2cNgaB]3).g,N/gK^Fa]aK/[.e@T
eg3OfT#:e;/YI@/M,IJ?8-+(d:aT@fLLN95?3S6Gf53ORT^F=c.Q=D@Z4[^&V[+[
DgZ_8bU7Jd2KCfB,G-33PTI.N9[AX]IW#)Y+1dG0_ffO/?KMCF+MBBB;O>1&/>Z3
^-7B7;O:Kc@H_Z9+BaE7]NSI[9G:K2L_P4^RgD-J4E=J5aCA]RcZ7<4X>(U==D8T
9K#_\>PRbP61+)7,_3RBEfM(G=;U6V.5;,W-__)+Y5d_\IBg:X=KPK(QcDC1,C[,
M-C(?.X4g\J#XT?<\G)+GO8a#K?f\&a5MQ57?MKDNDD_#?6;0G6L<&>PC=90D2NG
Ca@:+#T2#gU,Z1C?L-NOH].AQ;eOEH(>9eV70<].G]U[]HYQA]P/0_YR<^.WD;J(
\YBe7S99_D;)DR>L^CQCgFD=5a7\;X>WL(.VFX-@a_&a8[L/XRR1.]4Dc?c=R9d0
CEXOcg2C?_EBO/S^;HUW8LW57?Zg@5AX^WgN0.:/)7ZXIK==D^RVFQLg(7+@Y4R=
@D@\_gDMZO((Z=:C)\_NJ6gTVa:1Z#9bJ@AIF)ePVT&5@OIF2_]@01/(-Z_#N9R,
0[ZNK22()^XY2?A2ZVXXf7=R0FLc)]W#QdQSbbcF<E4WVc3,T5)\ZfF;@)&b950)
I:5IK/F/R)1^B1X5.-f-P#DRF4I]UA\/FV1e1e(/F5Y)U0d:PD^?3>_Z2GgJ6Af2
;UD(+N89gdT(<)Vde/Y9O\(PKdFYFJSN>F^,.OR\TDF+)8;SLW0A1XX5&7GCRAgQ
/d_L?YXWK=[KWD-R[[8J(\We[;PJE3B;LddGRH.c@X4d\KTF\K1Y=4eL>.L-2EVU
YAO@PJ6VBN9&/.3S?]f?dQ]#3JNF3=BM\]0C])aa+^NEU(2Y.54.bK17)8_(Y3;@
-<;5D?^cS1-eQ>.d)W-Q&U<UQd4)X24,F&dTL7N^GfMLGAaE/M-WAK+[1dD<23S1
91Bc0P.J)65b&:R&8?ZL1dcLTM.ZNa1OK[B.1J)>,#<<M,VQ7[^3>8&2Gc=>D77F
_A@:35fH:Y5=g^?>M,9df^R1^Y]3QSD<;+I:)#BN4aLKB\W^3gIdZ-LYPa23&-L4
)3[G2ac5O(K]FcO<D[#_:cV=OZK7]R[bXLBX2M#Z<KHdc6=cg=W/;Z1.4MP4];C8
>aT<OMZI@W;]Z<H)4^YTG^8UOMV.^-g4R65-C)_R&ZEIP4a\M_RcPce^^@fX]aJ/
JLVYYZ(/#9>ZP48F[)7BU[C5XS50.E[dcN^69fFH8[EPbTZ9N&];7b]Y.KHIO6;e
2C^>2a\PN3L86[b18]SR@MQ+:?4BT5b0;GIbKb6\839Kc0g7Q<#6a);\96A>I>(K
=.5826\JY>,=-<HF+9[:,7.RMbEcH#)C/1QbYTSEc?&SNTMZNg;CUfJaCW3-ID.=
W]<2T=@;6eD/7@1@b7-5V2fA.DDa4-eZEWB,QAL6+Af:4C7CG8.[YC#eOL:+D3:K
NU8[@O:QCCB9>TNST;,f)1c\eD3A^WA#<2D>CP?QDG<dc53A:ZXK8]MP1d;&T>C4
_KHY]&5;]5C<0>Uc9bI&5TKB;2E8_Ma3,?BY?:UOH9d?2ZK:<,HE3GZGICI#DTYd
;Q1;9X)\]4,f/N=]^F:^DQJT.<P1@5FbVHTLPcVDdS</)2J;cP&BN<Mb(&b)M=?8
-5NC7ULCN:@Q-2>R#B,^,.2JWB0-0BQ-/Oc7-#E97@;e.^D-E47O;K07VMM(?<Za
6KgS8;#g_<CLJ9Qe\OW^g67X(?-]@@51+/.ARR--=@;NTb:D,@a.??_J7PSZb;^&
9:I.):AK\WWEf0TQ?gDM-e)f1G<g6YT5Wa=_,X7GEefRM3;-\1]:RD\:,P)0@,9?
e\\8G5+_6R<\VW[LR#a7XUgfFFgOP&dX&Z7G_^G8=9.0XQ3GZE^]6gM@EBc+3;K9
_&68TWR==g5;4D1P1HP9)JDQ^@fA15b0gLD0JC^b4>H83MGe^.1VP?g(J_.gE6:P
F6ZdM-bEbfccbUMW]_P(LcW>DY67/g-YSM3aU[#Af3V4?YN-a\b>]23AU,M2^0aI
NXN<RL-8\b=#2+PMK9E4+L,T3MKZ7CBST37R15K1VC^Sbd@T>6PPWO8GO\CL_?F_
Y<NLKSX/@+7NLO[&FXCT]_-VB.ZH+CP>63>PO^FKU7Y8LL1LIf<FVA-::?0f.9d)
cd&Id[K4Q8,@]Hc71HZRb4@:W)WC_W3\EZ+Ncc8b+-.:O?7>#W=[1dI9O8=D8ZGK
Q@Y)8AEe2TcbXd4:<I(f35J0?P;a225A&04FTV:OQ9=BTB.5gO+]R]B.BM0/E27H
JD56_^82fb=NYGBCGQ1WeO5_B=(GD\,8dC#KHNIcaYg[_c6f>H/Ma@.J2Y60f/EO
Pa;H,-M=gW>&)@U71JACgSd+\5XHU8+4<d8[(bgb)7T[D$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
dYd.(O58cYeD0UL?Z?=-T);O40Z6=/XGDcYTadAK=?E;^)b?#FAF0(RA0C&U2G&(
+(AADDQ8<M+aLOMI)=78&]&?F27I4U^7];VE9d46:/A1V=@1?8Rc\@0&2gV#d)BW
,42.F]dG-JYZLe,YV/@adJLN5N=MBU@Kf9&-bXLcV<TGL30]3)Y@D?a[V?@G]Pg]
]3Z#b\8?42J0\bSOdO-Z=,G^f=GH?-(I)_[/I0:,I3=&2D6W])B=+WSGIUMSaZG1
>C:&Kf38>[McR/D]CU2cJ67X/aQ@VR.FaDFH<U5,gf&^Q0/OfZME_6);,<]=_-_<
HX@D.).6Nab<90/^L..O.+@LCa>P#/N-(2e(8gU2.:C+^7V(P\#3],e#E>3^1;a)
V9@]#-b0P3(N>P<^QW]TX6efc[GQ&TDI1Nf6;5,Q:3Qe@1_7(1FK@DbcZ/Ca#3KE
bfQ<NfA81I(W[ZSY/D3PF(HY;\-47aA@Y<))?Z[M;+R=W;QR#a=UZfR=N;UIN&7_
3;Z;:SV.ER9(cAPBS?ASF7NA?=<7[c;HC57]D?LaLRKUJ6V^5/R1+ZfAD1\5Q?H:
XROH#(2IJ4QHY;IMT##]?JN)3EZ(K>X#>MT6.F2(#,E.+4fg+M_QA4\_fJ&b99X=
Z,ce9:B<_bg(1^;]A^DO+JK)BTM-Q0J.Ac8Bd1D[4J/,R/=6M.d9H4-bc59TTRIV
B98fL1[>?Og@.3>#&0G8G:@aGWa4\2eKe6X3LR/Hc?Mb(W.b47f)eXOA:89P]S,V
e/G&&R)6U?&aR;LO@^U<4_(]CT52J^61_.#E=OUA[\\/RL5R8e\V.^1?C;85:>@,
@Ig3XWOg458.45c8.?,_NG78<7Y7TdSPbc>GCX-<0VYEJS9<7bP\4AC+46+U;<C@
EfNY8B,a1cLaJQcN@2[J@a0TIJF=YEL3++L<773)<],5MWPL,OVS5Z1RB,7H1?aA
#UKK+0.J/2f:2^@3+V1J-a,ND&\XAN+4(VKHU?==aPP=N<;HOMIN45Z]V,(@G)&a
]0Wd#_4O23dVJ-5],+RG)KaLHH0BK:,g_^(0P?I4b28fB[.SdHd6bW+#(UCJbNJ-
H&eYGDC1]VQ#ScK&9KRBB3=gFCE02_LOV5/>GFF,T6W\2d4KH(Ca],MJF2bHTfHe
gC,OUWbQO74ZKT;W]K0.7^XKe++/)/H-J@HO97R-W-K9;MX>KFPI-RQC&/HNBH-=
M@AGgABI+X]-)L9##G2JfI^_L5P3)bPQL+88E0VbXX[>4VCR&11;MXT#=e=I?&RA
;dFcF?abI&5eATAAU.dd-[<)WfFC+#f\&\G]gP-D9YNDWUC=(V,dM:1YEM<Kc@JA
[+H@@/^D>Q>A,;DPF,g#D\E2B.aIa6C=71M#0S</VB^cE]@4fK[7>L=Ldgd@-U(M
M]@dA03=@?,[>D2<+S1OJY2BdH_^=L8).FX/#-^Z)[/;f&H?(84TPcc:a1cAU55P
faB(.3CfB-A?7SGKMSQ\JBNJ5e5=I72C>4<76L)TX1GKfcD3dO)O4SXGH<6+>DQ5
/Y)\]O(fHca7776<QE33AMN\JQ5870d/-7BY?^aNY9>;I)-?1=:dWgV-R#8V60Gd
+9U.U<U@[ACd,Z5bQ#GQ@#Ocb):>V?REW&:M8^,J]DFW,aWD;>FA>=T5\;)H56:T
L/48]gBGEb4PR?PQ8[TWJFXK4C1CF58(B_Ue-S3/C:=H@aTd08;A(LYHA@W@dU<@
adY^Q\EXP\759+-SES.#4KBM7Rf,&-]A.J.7;BcQg84TCSeND_&9WSH3HEVE(5Hd
PP1<WO66=;OT.\Ja9.14F/UT)H^M;eFLTK41a/\54VH_ebUgD(:TTA86BXN6WF-4
RX]H\4gUH\25U#Z+BON\YE>KafK;aXBX#()FXdMANTAS-G0F1J,WHYLG#((:TE.I
/[cIU9UU:FWORa52T0eUZd,(RZ0217C;9]c/:E5JFRb06/-ZdXHb&RGS7\47f1G1
<I/HS7,&=]=XCX]_NKHR.-,PdM=[3[g]P4X5[48WZ-GR26V8VF+b2[-PDG:[(+ER
WTcfR[@d2@#KIH9IFOB_VFIP6,D/2gW&/[MSVZO)U:dGG#3RJJVV3]WH:cgUSFC=
F/[B-;Wg:/1@NLLfR.H>dgEFLOI@1OQ:.GHE6S9JN8ZJ?5&<7Z.8>H=>\O/K>]de
;<8W:&&X[3;8@?,[,ac52O/<7,;dV.cN4@)ARV?1cbfOO9g67MW,@e2.Y-Ue>E_-
[)2;5/@UHf#:YQE[ZDV.de69>VN,dAW^dId;W;Wg.?^ebFeD8G[@Cd89cd?7&^@3
2#_+&,aOYgGKZ,=EKL7-bKH;d.G>bJ_bga642U<H?2<.Y<^FAPWXaYcRSSNJ2]@W
=A:Q<5^&P(:IU6cMU\c.F:3A_V7PU+;[?\(17+VdC89/VF.PeUBWQ0GR=VP,T4/e
::K)0A&7]21Gg@C\1X#<M&X]J\.]Y5+<5bLZ8A\PAZKGR68&4\VJ5d-.Z>:(MQNf
>/+1GZP-dOaFU;)MbJJd4PVH:QDGQRM+fR.(1g_51UKSU05]#REAgN[H[+^^FX7V
()Ja#HNS_[#@82Ae^Z^NL/O7-:&eRLA5&&M,F1<L+NJVUaR+:BK1bC4S2SV1bcSF
JC=.G=P-6B,Y6DC3^.T.Y2)O?>3VBKS.=M:F#dBgL0/R^H:-V_<5_6<26SM&<A&X
_V#PG+)6eG[.DQ-&H_S?C(3OVY7)^LLA(R<(767gBEKJI_(24a,EERU=^^e]A,RZ
4K^OZ^7_2Jd;&A09A/:5(9O5>gW:MFHTbS8.,.a0L?)RV9b.BSFDVY=T:J2Mg=^B
K?-L>M]1<A[DA@I(Q<NbER)__#>gTL4^HA-VfRec>egba<=[gS[&P]/57FG585IN
)J7E[W]_LP]KZ9D,-cebc&]R+J93K?=H8>9=#QaTL0=TEA:?JY;B5/A1&M13P.EY
+3_&d1^:HEK]d(27E2?)TGP&Qb=AD]Jf.d1_K/K(>Z^16W,J.=/Og2,5HWCb3#0T
ZSJBU2+WODb:K>JV;+5+Tb\@(XG)gNO=,gS#GAI714(Rga_#]4AB@U<XZ&=KSD>+
(HPgfRR@^D64QESTg_IX?JU?aV,]M596\a_K;Q--bfIAZe@#d,HWZEF7V0NG5/NM
LTJA=?fEJECb(M@L.-=6eR3JcDf=1<[&2UZ.-<bE;2[D+f8T]c>@1RV_CGFRGYTR
fPG-ZSd5SPf\=,)7YE_Q;b,fd<:KQ1R_B.FbE5F+G].6Uf-d;+5&0c338SX1\8/+
C.5+0YMQb<\I<.RLS8S3F?3Y4MF3g8KK^6,A)V1bF^)\&e761H:CQeYAeOWLAKI+
;G[>6BT)(+NUP@0f(:E4JDKW#/VU:UA5\YYY?c22[DQKYabba1Fe0b)MK7If:AF.
M&BE)K2Ef<N3<c5[7b4E7f<MIH.O(05._5]PYf#9MLMN]/>?CTbQc0S^KCcdS3TE
\D1)M5cAEKBH#Cf0<ge_OfBceMP=^<X^-c83YWR9?MbD(6SCU77D8H9ABa3A2OgV
:9LLH.1_KARS#P50\XZS,0Gf#g6PUWB:g[:-37FbRNd-E89Y<N@N[N2D7g^eXGH.
Q_,X^DMKPfQ=dQ^1ZB@L\AbK@##QKD0C(08bO#AV<NTZd7-e4fJT8YU-\Q7aSP=<
AfVHUeI07HFY.^ZV\bJQC/NBe@IQ;)P/cRfacYQI@4(ZFHOZ9XXL>JNZ2[G__6IE
X(?RfG2eXHaUI3^YG3L3#U&+gOAVCf9-RS@75ZQO(M?>BU@@D2@/()=\>OPMfG]f
[[ZcZEd4#fg-/S;fBV/0&FK,aHB)6I3G_3>ACHD9=FS0<0WO^GX:KSKFE=:._T?/
X_ML:3R(HM/2D,>F&WgeZ8^g=]bCH4O6DQ\H)b[=\Y\eGL44.?#L?X)_cX#.GB#[
Y_O_)7-?HPVF3]<GPB\0;X0,&OWK/V,gUaL;0]GBJ3TK7=O\@41g-3L\729:X+a4
3WIKII>[P\=adcY2)RD5e[N+Z.+:2gU0[Xg#<LHf9X6dTH\V@9W:D[:2]T>B^b_a
A.-W6X#2^4VXgLB?fe=<<>SJdQf^W26:BFE/6fFBPY>X-R7M608=3T\e=V9UCdc>
]-YH0E#R+Je55_PAeU=_1^CG^X,XM/S>K)4d:?RQ;GWYE)H#[]Pa8\6/>V-eE3:5
Q_;aINQ]W\MbIBB[)aF)+F,?=a<KI#b)dE[2TA]UIE-Wea.];_9A/W&#^#\HCY_@
LHWW^4JT1G<C3;I_./]aSN0#?e/\MYdS_6Cb1&#gI&a#-)>3>IZ.EVVK)GWL_NT7
L2LGBQGMJIW=)5/H^;GPaVPNPcc#]BcI6_gfM[U2.+(03[W,dSf[0HKgJUFG<fJL
8>U^:_(g9:dMH0MV4b#IR7K9N#aAR-IQPKT+UJJC=JK^PU;WdKY.#>15(Y0=,M4U
cX&PBQdF#IRK):CF3(Z1S5g]Sa2_W<TBV+6[NP18bGGYQ7=)7P=T6SDR1TKP+#7Q
f5UdHA0+f=O?,1/<.B9fcZ\<AZa4NJ1GD6Y1/dJ:IbE9O\>I0;^\bP>V4;ZV&;7#
J(d#C<:=5\?(P2Ed6/UVQ&?,UY6=-HR6XJY5X0O#f9LH/cV^ba9_2#c_K@Ad7dbH
d;S#Q\5_N;Q-^TT;,1RO6/AE8FX+Zf:H1&1?0?=M3&?M[MGd+=1Ac,PZYcO(B<#<
Q5We[7H/e;G7L,(U6=[7TN4,-cUV-EZ9W1QDG&Eb]?/RJ&(Z7IEY.d]=7+E>eb_5
(=:N>c\P9B03b?H+C48?,8YXM]KREF2)cc4Lg=7ZSF)bKA10>JQX8E]A1:0Bb?B5
UJF\2[WF9d\TEaeB_S(d<dU)@<#/HF^-G]L)-EC1+M^ZXT-F,9?5NJX-8]F2\#&H
(C(d4EK5;+FH)3_#2YYCWGg46X5:a]6(N;VOg\,cLa24&F-TMH]^+IB3B@d43e,W
)>D^H@4:)f5A1d<SH@&5e5ZHMLO+A;\6Ie&=bMdLUE1gJG?e<R:R53KW42fT:..g
POC/d(:Z)K5EH.Q4->H]-4)5(5K8AU@17fEY7^8BD/>8?,&+L2\7bbD:>U-U4-ff
7<VUcdKGKWL+a#7Hb<G5GZgJIUQ9Y)1e-RR4Z0)\D?N(2CXJ,>[DI2PTJV4L5U;R
YW257<EJ#JEN1(RO7=;J^U+HcK-A@KVd\AZ:1]0OcP:a6>dE[64PAUF84H\<KR(X
G6BQZ)g]a+f+g?D?MN-MfYPg=FA_eWH4CEAMa?#?U;^W/SPII@^JCVa9Pe\D9H:7
^Y0D(=0AbG71\12d;T:Y;2.>/M1=ggT2M4U4gQ86M6KUI#XYB4M[T75T9?]bW?#S
OOa59_f1?TVOZ>DZ6Q-UE4;&\6X_<W5^4M_IR_c^SNT7.S>U9I,TF3VC?2b#?778
>\>Qc6\V7)gE#WTOa^_@=f&)U\IX[0VL#(XNbdSH;f\TFPQT=ICX6G3&?\+4A/8@
T5I6I3C<N9:d:RX(g2S#H_A:55T<&91e[4\)1&Z[\AFW.)5-.LJ9KdCC.\EGFd0-
(KNG#SFOa#TQN4Ka@Ta[40,XOV6?OB?1f@W#-g0(Y4OJ<e3J&N0@6a>TB,bUcOT@
6.@#5IDJMgR)-E]5)fYRY.J9[G9N<N3Q55V9d=DB-R62#B<XE-5?8A9)7EgG5G?T
EeP5M[P.QC01gN-W-6XT]7]_e,1EH?/;/OW_4Y._g2_,\-f\R7YG4WJc5AT+4gPK
Te4DCQKG=JSP87K)8W>FgV8W3fRgW/]&#D>T)XEF#<>Fg]X)G][IL?KXW>gfG)Qc
H(df7G3GXA8gWQU2/RBDc:X9#T]H.g8a_J909+_92&e1KLTE(b@^1AaR6_@=d?,b
?,+H0PZZ0KDaI+JIN<WZ].F\=(aK/MdSLAY>f^gb(U&A3KQG?:ddY-:61(K;791[
3YQUEU&B:/R=,42F\\=A1C#-QC0^9F?#G]N:@e]eZ;4Qg5W2P]eC6DA3SXW-a/[^
Z)BMfc.cE>(f1Q-Y_[QX?R>Z4(>(Tg/ASbOUQY#P1T=HG/XcHeJX6Ic\WI_c7^7T
dgI(:Qe[c9..3YWD#>@\_W&.[L/PF3B;58)Y]SO6:TJ<BeO[70?4+cbQP\.7RbF.
#&f=gFR?5TP13;Oe#X4/E:S>_SeDC#^,_eCGB;@K_X39)V#fQ[_B9D.Ua6EeY,QQ
6Tf;@fJ>5S:]^[4/:XA4BT;+BC)X1eVYAFZMJFG/SE62PA>aa1b.<?edRQWJ_Z#<
dV]RKY)e=9Q+]gFSC]X:Q+dO4DgZBH--bZ5;?;N2E4Bce-<ZeX;V82PW0M9e&=@S
YR^I>5g:ON.e=gHDBP/a=-53K8NQ?(1bddL:X-:\YQaVY7bV+6N]E&K1[7NW.G\D
fRKPDPVV5?18:cEVUE.EG5WJ0/TbV52eTd@(>KZ#&I6]CHSEa28[11?@Y]T39AVW
1:-feAfe<49:OZB-7IK#@Dcg8f#)VVLBWdWYUY<72:N/)OEW4fYFcVa4)BDaPFaP
RcIDZ-L<P>a9F4@:#0b29>9S-,b-Z#aKcBc+ZNY(\6A5P7,eC2)BaVcM,<4&;g7A
2S;gbS^5LK#dcf+c#^<MGNf/Z[U^ZYaHWP,R?dL/G)@I7^La--IG(_ceG9^Wa#fJ
gKF040PL76IM]Xe^bOf2cG7<80_(GWIFGESaB@,CEfNX1F],6J5)2O62I4)<gAPZ
FK/A[8H4RdO#Z6RL1D4>.5FN>f+/@5a:1_NO>,0)CE08=#ZQS/ECJ-/9P&dP4SU9
K0G1J\U.9U6EU<ATA/#9Mg)_6WD#8M+IMLZd+UV]_MD&K;KP5+@=?eK325MRP(4K
.-:6LPJVA@&9Z6LZ?E0_7DM4<1>f<b9&fS#?J5FAa?V3d5gd23X[PVbRKK_I^V@.
R[,8R=Z9N9;c>4HY><D8)+7[:;TAd1^2faT?;)Q>)MIP9c\?MS1P.\?QC#VdF;(d
EAf7&;:1,AH/W<GeV0#gCZCQE@NN9Q4BL,B^#85ER)ND)6TGI6N5C5FN?G[-\#?4
=;D/3((E0We/A=6F=(URAgN6FK\X.bIdR]4LHL^>GeOM6+/61(E\(9M<GKb7UMND
;=R2/,DN[9ONEd(JeOW?E-KYca-2&\0/U@41JLD?4(>.N3(gIJLJb0.0T9F-D@@+
^ZM?d1(E(Q+<C-X&N/;3BBX+J@JNE#E_UMUZRVZA5)_^f?1/)1/A?c\[XNeMg2E?
,ZWT@+Cb)NP]\01HK9)?O/E<T,-.2JXEU(aEAXSQc?c69G@5OAb-<<Fd2I+B^UQZ
g3Nb?Haec,)/B^Jg#T992AGE\4-NK-RWKc1P.VZ.<>R[1b9EU9c_VXBW6Z3aEU3Q
;B3=L_>P,5gdKaOWB-ZJeFXg+#37=,TgBY[HQ>-BYFL>=c3_Fg9MKVV7#_DIUTf]
g)2EPGDJ?2bE]cJI(#6LeE^RW+ULM3,\]AfR1E8e7gg@/HE?8dB[I;LH#[Y.W;BC
fGQCN,gPNId;g>X)g=,EQ^;G4Hg7Y-7MOUeE;CeI3J,Bb)&FYTUKBRC8D:7?V5TI
F)U\[3=]T##c7[-]\f:4JM(@#6<BHG[&g(Re)NUCG^;1gJ@Gcd:TPM]3VN=\NB)3
_</:N-.E0+VTYECe;TXU>0+-)]MfF8f4[\dT+5Q#<.@:d#Ac952fZOVC,NE/][aK
)Z>H+6dX<.M@D1+)J@-SF[:EB3OH4ZUBB0L\\/,0c3>AF@;.@3&-+^EIQA])T<T_
P<M:Ue4+SD;FgQcP]6)1=2AP(@TY6dK@#DM&YEB,R4,PM;X5Y<MR1:gg]P5URf11
409aHQgCA7Zb_GHa]M9b[Q=Ve/[_GP+&XN1=Uf^6UJ-U,B^KW:NL?W<83\IWbRaW
;E&6OcUPHDX@Wf6.XY/IW^7SPd42C4&+#eK_W8gN,F<MME0RTT8EP(eBS8@UZf(]
;@UULM)Q#X_67AT=fPC@CRYV(\,;/^;=f.6>=ZF(NDBJf/8g4R6c4+0#]5A^DSdN
\GJ_Zc@/5Sc=]4/gUYb.^>[+<D=+ZP23X)J^,/<JHZ0EA&_<R>CU2\4)0PfI]W39
4W2QbD9B[Zf\cWa1C?C&<<aS(XVC&7433gL4NV1dM57A6K1]SLW=edBDd\01YgS]
5=12_)=:]_<^=81-eUNTX@Q@<8b(:6-#]TTLY1N)L[LU3CcOB.((#E)3T1Ud?XbN
0dWE6FDa+2P_Og-NL=(JXJ&,f468N<T+@#+\36O[8TY37:L^Se2:(M#_UL[R6eDG
U@2^IdT(J&0W5F]C?d?NIS6V]J-P3+8F-XH_CbbZJG+bF6@V]9N20RXD\N.+N9J2
eYbQ\WON633VT)7H6CgDUL^JEPC#Z>;-[PS#\LT#G0Pg=VdJY^-T)RF#b#:<LG4^
#/OC7UdYEQCNK^e9X^4J/g?(J.c-Bd(Gg1T.cd8[1G6>d]JQL&++GMU\:1fU6B5I
Zf,Mf/5?10bWbQ0Y^I969^Mf?<F,gIBFE&IRY&SRLA]K@2\,(?OLa7PPXOP+F/bN
+:ZD6M.7:<?I5;-OYQIHB;B5EIgfN];3[;#<1[?K5M8VOd8:9(a8#Md\.B7J^H:Q
:L(1eMfT=7)MB]3;TD6(A)X:aA(b,?,(.Q3H1Q3IbE)UEB49Ue)[g)-@g5C7WM6f
-4/-b.WPYE0O[;]WR2:@0_8P)..H,+)4NG[#0_G16EVQ55?K@1L2)cd^I71NSf^(
=6B?;6gK<>UV^5X,YVSg:B(Y<aNfDBW[RSQJJ:6CR\_Z^V^d:?GA@A?BdcSUDgLd
b_HB]-V)ZNAJc6)<JYZ-DWe@YG[Q2M#4CF#b/RReG8C_c8:d67@Z\4.>2N@?e;UV
52_>=N4MMbDGaB0Hd75^[CR_c;&0<FBPOg2;@YHTJa0B6J;K8Rd+L=1@TJPM9-R[
&;gIbaZNdc>5Y5PRG(YN<B4e@^4JP7-4F=dPHN+?aPT#a#B(g5JY]NDRBbHKfK#P
V9GBcX,>BC4BR8-E.4,;^Q]:D?;1a-g;?_Se36>eK#C4Z:;,O/NM+5Q]Y/9.)H).
2Z0Z-&D[O1==V@8RJPVGXF]Y^69S4](8aQ?@N;7KY;^Z/@IOK4]Q2NX;MJ,<T7Z/
=<S#C;V)+dRX<(cA0JD@AS5]WJ_;GES@C70CTNPC.(H.^5Q)e__Z_U,&+HC9B_FX
ebUM[HaeOQA8b>H0QO.S,9ec3)3K2Z7-^-9^f[.O)f<<4:f8)2QB1XB@89X91H#U
4]?2+TgOA]B1gR](_9bAOER,@e?E-FN&[edJ/+>25@,?;g5D#B^=YX_g8,.b0OED
CY(H9@bM;a3K.>4bW1NB)A=:F?KE@E/5bQ4Kd=_@P32=#dM<+F.c9V33.[37g<AO
.XZC85T\8.c:EI&S547W+,8d44UM5=;Ddf28J(ZT:#b]9+Og)5E,9F+cfIL58&ZE
69ZdF)D&[#A/?^^ARgGILZd@00B,#\60ce<e46/0#)-V=:W6,XIefgY,g-V;&CB9
X>;QN7Bf-#b/e#Y#^,aIMcL.2T^P?J]H629U8,55)/=Ob=0=H0g0TU&),(ZUA1Q&
HP;+GOJCT[&W:Z1[=+@1dBIW-NP(U6NLDZ0M_RFZF7C27,ISb<>e?Q16/bG[\(bY
I_2bAK5.;:B;1e2^BB)CKWV[f5(?dbECM&N5bAObcDYRdAZa]Z+&1RF<L9Oe^F[,
MfP)g?_YA0@4cUd6A@_&1))KbKVP/6=^7ePB0WBfgf84;V>^6D=NK&(Y=cEB>4BL
/XMeac0OD-S:f)OFTYM)UY:6@FJW&GR]9#_cWI,)8:4J/;>ZA)Y@NdgK_Z&A.&]:
-3#GEO]:FJfUaE3#I9,P,VC44C&VC([gad(;C\a-Wc.aR^CL9N9Z-BJ<bf:(=cYN
GF>5#-,)BcOd;@f5:QR0=f>M#f0)IMDF20ML[Ae3P<D\2V(AfadO=>0P:Y(BJc&b
E5dCGCRF-ULe7?T?g:,U;KTRP;ZB#eN:?VN51FfHQX5CA4E=+1]?/HfEJ[Cf-ZTK
DEE7)H.SHTB\fY+d))AeS:a]^D0dG+J0>9+3d#5/X+NeKDK(MLa)eF74YDSJS^E(
f]3CQKdOZFZP\QJ9-J7gQ2FZ6)R=9OZY[3V9;:G<<a.f4#2>?Y_fD2ZVd[[A_2Nb
&aY@.2=_W)E-)VgUaQfMU#]Y_[a3H/gPbTT:cGKgIBT#W7.?52)RP&/\M-Y&cF,N
)W80,1PH0H[0cL+b;:,&F;QC]R3S\(?/[2M66D#gBFQ=3:_3fQPb<#1^N7OF]\[D
W&YL(c<TIOJXE@G[83R_:)GM;_@P]9agTR[XL(;WQI;gQ:71V\#+)V/L45J)L=&I
/C=WDHKagH?ZbO+2W.Y+Z/29]@3K[TNSc)2:-XZ[3V>Lcb^#b1S_-SaYIBf)HP<0
9(RH-7XR#X:=X2;)?Y+3O_(cBH+WW>EXY\F]f(2LJ0eMQ[SMC2;g0AUEdLV0&02]
34e9Bca+26.a,VEJO9-_SS)6Sf;;2=QCTXb>,22=ST&C?OLY;O,BS1EF6JE(0G1-
^2(NVVSVab_IAA,b1B1SRGEB?J[,\E8.MV\[HY6OOCHYPW(6F5R^A+71RB6^W@_<
C4SBcQ7Pf58Q>H0605fT4R.-2Cb/:U,(YI_:g.UAb);G&)QZ]AAd=c1D1;7_c@W4
M]0KT2]6ZeSM2Oc>ecVH/3gf5SBI,8Rc@GU<5>@Tg,&OB1I[#Y,[(\[[>D_MC<CE
YG8,?LB<AJ0J:@g/c;CXH.d62:WRZ6U,G+AM42E^AOY>L>5MS)LBNZQ_IA>eE1;e
7GHeY;8Y_:HQ\YKYeXRR1+b2M;TS:N;O07(EO@-aUGA/BLY+9&gbE_F/2a_WXBb-
BGD@<]aP#0B3D8-FV_B:=9O&QFdcLOH.R[05X78>H86b[>JWf57dYZ@R1:,<K846
,Ke1HW)NFV7DQC[RI#1;+<&(EUI=a[QZ_6.C_:T/a[ZK3YWJC&OEa>WZR,O?bZ0A
+cO7&2ODA/ID7feUIDNKXdNXTVb8;_:YJ-><@\&LeW.G=P9<E5H.<Q:7(C5A[C0^
4/YQ4BRFUY&WA+U>>S-P47GTA)8NHI)XN?ZI1Ib\K2S-<O;332ZJQU.Lfc<</^;[
Y:dQ\9Wc]d4Q1MdZ@Hg5=@2[XZ#0@M1I/=#JXA\<W6Q.;-8UN(MS8>aC-:0Q<aTI
/J1X@:e,<GC3-R]R1&X6E=]&\E(_-\Xf/8<HYVR:J?WFgg-.Y/>58#A,=3CM?B>N
MWJW#WBK_K3N)\/_EB-M(AE]fZ=F(gZ54G[EUgH#,@FccR#g7_J/cgJSa;^\O,Ob
>7Y\+7e\K]:>F(VQW:V^.8];]EX.\#=7W:MPQ2VQ5XSFDLU)1X3bS+E:HJbI?(=?
WbG>AK)];AOFNQ&H(&?01QS]eA@JS).>c]7NV\1XJD+@TXKC_a4+X>4&]1Q:QZ7:
8IXD,G(E(2UX+)bA8Q^f=81O0X,RdHC(a\e^IR+3P?8ID3]@b95WI]]M6:2CYPV4
]]O]L_fU^_fcK84(?/D@IVJ>WD@a)Z,G5_73(<4#61E,I;R\3LQ]C_4<b:^U9VL[
C(]Z9;JWfK3R/g22BedP1.E1fR)8=?7_L>6^#,(62^[-UVPLIaK4.MI05Hg5#667
gFB_1M0-<fZ;A-^f:)\OQf_1aLBF?\1?G>g8N\C]BaNJge@O2=&6^1/+-#&M;J;F
b7Bb9LL02&e?>e\92?6&F_LWC1Q91?9Td;E0;Fa&?gcA5,f@RQ;]S^e?^9])>YB#
FL)+]IQ+APCJC3)-@;Lfe21?3:+AI9W5AaFP(?Z9<GM;UZW9QW+U.YSYI6;77WW8
cO^Q1D(]C\-gQ?dZgXXDNI0D__VG8UE\6;PXPCf5ROZ[XR>XW28)Q18@L&QF,eeX
:HX?0C2\C+7U;#&BFTZ7RJ9PbN0K9]PVO?5]X5[cO244D#W_BYPBKgRHG//fB1_g
5RGEM;J/:+6.6?]>;N,D>IKQbMB7AGB5U-b7G</R7+2R:.eBC7DEY)+Nc.C#)K5R
W]ef+R-]g@GEbF4S[gD:.?3WfSW]V1Y2HT,&^f)0F66Y\1Q9.@U6<FDQE3HK-,#Q
F,R&b?;=Rf25C(TY7F6PB<c?P2R1/NAEJVAP?52GK&@>7e^19Hb0+e-R_[>7A1FB
)QX)d_2](_@_/UcfJX>+7WHA6.6=(e.T.J-7?6d)+]IF(<_09ZAL_4]E1V7SRcOP
X>9L.B[#U@J+NRaQNfA3Ne/SEa819=GXI\Q4;JMK&J.#6\PDUY9P-0-B=W#?c9?N
3f&<U+5^Kf]VW;XCTHAS.d13(dHE0-=?Z5O#\]SOZ)C7_7QB>c=>;bUHdbPO2CKH
NfI]T+/,H>EPb&?F[[6HA]H2;^3DZGYOa;:UVXP3efUP??V3[N@T8=B2LBe<Ue/0
C0YF;9bH?ba^NIRPN:PIdDcdE=WGN8=H.G@c(D7A&ZTG(7(JDH3K[7XdYJOd:XQ.
6fRY(fd&9)7N][RA/b9-ZYR,NOY2HH_2M23HID/M90cH8Q4YY2WKDa93A<KDAJ\_
[@P#X#PVT.=<;?<I5HUT4S26P@O6f\[:MGBX)J4C<=U[;00V1KcS6E,E\]+5Z-/b
ZZ::P9EI?70NQc?.dF#g;gcRf);)gEOGeZQK3N:eUB.RcH-]I;IWC5_7d<e6P^RY
WH&74-_V5HXaXE.c/#V>N/a9>Z&H4DWNeD+_Q+?NX-9PM4-.3Z.K>JCWb1R:D:L0
-&>5O[.FS.gO=GRK7:,OH=cFM6/L/A]U6)5gB32Bg5R#XX^ENMM1a^bd5Tg:+<7=
LH3R99VG=C&4eY3N9Q,PgJVfXDR6aFYBJI?;/HI[[b?5U6a99,KH\:L+96F,?Hd\
OF6((Gc8gMHJSKZ#,-[bD6E,gHQ.@SYS:HQF)(b#b,CV&80@]1+6<7;MA5SXe?#G
#_\7+VRP0HNdH2;>+bM(+/-6;feZ^ONYY8I2O=;Eg2KO)28D:7(TK;SUeeY]<:Y6
W<L11RC.^1B8_SbG2Gc9aN@eR3g4T\B&[#(Q,:XS_Z:Y>g=;Fc6741,97](Ld3[=
)eF2^7.SbfX2-H7[#?)L72GO(IA#&WbBM09XO24XN=GB;+3UG^cYC)BGJO\);(HL
A37\ZW<KE1UX1A/OJS\_6d2ZRC;4?IW+aG#X32P.0LAd>WBaWb2P/W5;?;7-+a5M
\-TSN]ObC,Eb2F:aDXBX7-63eOI_#IC8Hg>=B>5O9J@SPRgg3A7>1JVeM[B0a&ff
5Q14@V6)]gTVA6-,87B@71dA(;P&[=>T0&2^O3[Ke<:.?<OGL6fHWTfA7,S@7;.>
29K6ZTI](H2RK:<7g;#B+C9+;T3O:;eAS+^3-4ea^.1GF[fHU.C7WL\ZP?f7Y4?H
G4(N]ISTeH>#cU2S0N9KYFGGPc=\1]ccULbW^CZ=1>GD2T>Hg;Y:4_4fbQ^Z])<_
..f6Z-_0C=AbOO&./GGgLAe/<3C8_b5]>:20RJ1:WD2f#HdRR4E1BJ6JIQc@XPN4
U#cEJ#9Ma/T1a(g19D?[,#RgMO>V2#2^1]7PF4#B5/T&P/V@U481A-]VP3U)O_,J
W3:Ng#?MeX<L\B.fL4eR[3L&FPF1ZYc_41;@UZV2M49WZV/6Pa4U0KSa)<ULJ45R
5/VI&CMB\B9[6cBPC?(;_@9)A+A0&(]ISK#-FS@E)\JGLV#>9g@c8RVA8g:7O9ZI
Be)CGJR36fe>H^6<b^\Tc@<AZfUWI[Re(J-84]4(>ZE)=P7O1.MDOUWg(UW(0+Z9
NQ\A:G#]V:W3,2Se#K6H]KT<A74#R\df68ZJTWWFf//8ER.ae<[.Mg2:\R+6N<gD
Ia-E+]#@XPQ=OHcgWV4=Kdc:bB^7Me&9]M<dMb73;=]HJFN)AD(3ZR22>[@3+]7+
Aab.-+8-WU,_2?9RcR7-35&].=\Hg^5N,dX>;/#[b>X-Y(T6L0A1Z03XSM=d)WO[
DO=;V787-)]Lbd1/TA^M5L[N8.\5CE7Nc]WR3.FLbTF/HF,9G-8E-fZcZe6GWa9(
\_9B+1N/#\R6_d@8<]eN>J-_,W6VM[WdP_FW.063M/Hd/Y<@gFKMdJ>IJ<VJS<P@
_f,a/,T)+P403:1M9DOTeFC\>4O4K#C-3SL-<0J&V\;cTA@\;P3eIC4VdH4+2GNA
F=TN#GB??4\CMLe+XJd#NV/)G-4f)U8>JgKKWK<f=I@_I,[Jd1M##/gJA-T_F0TM
&WK6ef2T3Z74^G5bQA\Z\LN]Z(H0^fGLSO=19&a?AH+N;>EOafH[bF)7550.,7Md
D;M-.\>T7cG#--Q(J[VAdMM#KdgE<?efFfaGUR&,922/QQ2_?TSL_CPLI@T<5f4D
I?_7H?/F_\99X4>4:g=.]AK8;7GLMINO]#<4LE3(MT/98#2Ae\7M18_9Y\L??Q&L
]D>..7==)03=^&;Nb]07\=RH@7UP3AfP9Z@,a;Z(C#9:aYADD5E?H@8X.WV/_)f?
.Y.fV=2QMJ12B/8R:,LUId9\LVfK#b[X<,GIUa6G4JRCQ3I&@?SD;O&fEY5?5-[G
W;(E^I1aY?,e[cYBU<<c4-OG2a#VA#(N8L6&;9#I51S?MU,QT4Y8+bVCQ(WYTX7CU$
`endprotected

`protected
N=FONXK@52d;eE/Sa(F_efX):eAgAZDR)2^S/^=T7]-+6#0X8),(7)a?[,a]Kb#M
D8X<D&346-fT-APN]EC?U:X)2$
`endprotected

//vcs_lic_vip_protect
  `protected
\X-]9U91_Uf6.7MKBcAd@YgQ5_.-:/GfWEJ_0;EW^#3FNGReRAR\&(,E<gg_5dW]
f=@&9(?e\S_;e276EA7:;c3(gN5=g^MTH1Q7B)gF.=4\&;,fEXQ+DaNQ@CX&_N;-
fN5bfPP-K6E9U(1ZO23UB[#<WI\,/R(:_B;g?;B8<:Dg]<(<O.A;d9N+Pg)0-/bQ
=TTCN:S2/-]f33^^:NQ:Uc-_Ua+5=5VKX_>AE6gO]9c^W\,F83&3_:&EUI3&#.A<
OHc.^&Q8ZBE?,(HZf\&0[H4e,fF6F.B_I7V6J@:O_ZCQ3NS)Xf&-6SSA-9JdeZX+
QG_+YeK5fUcE,+Hb]H&I]Z?+-ZS.g]HGa5HI+0;2fbQ<2G?)7AMHGNI:8.?RE,_(
cR?f<S\&a83+V_N)A+;)b>IUfd=T,Z-IV?.&X#41D-VEZ6(JLQ3)f3/R-)R#F9]d
PT:<IN\g3XMaCM__3JF8#fCHY7d)QUd=6>caV/N96H0(eX^C2Da#RdCcR@_eMJTN
d,WPXOVGOBU+G^H;J0^@A.H&+\C#A^:FOB8Xd#7#/ANI0<+.UA;(e(EZMa.<-5D_
^.5^S396c\HO[N)a^OZR#_9Ee)9RU2>:37E<DHcDD]B:,_J@]G.?02R0834&<:HH
SbKF+;dc&CUM\ADT-Hd5;9Bceb6)3f3Of>c>)GNTPK?)XUbeN?GgK[-@(7BI0EBX
TWHJGZ11MLe6)dK(-0b#DHGO=[7ZE-cb;LRX3U9^4A)^1I&WDPN<0Qb3VWb\+Oc,
>&52CaV;PS26J;>D;3WaNd_JQbHASJ#]8RdFD96(3XNPeNE_TB8L]^4DfE:MdYMc
4c1?_4C)JG-E)\^,fE#?[0)gd#:LO=&>R3DVHGC.gf-1,=P7ZHF)f(]-S4IMKH:B
=fKdKUgV+aae-Q7<1)e0ZRWWgLT^d)+4,W(Q>@NY@5E6_CEU=98+_D2)IO2Rb5]_
;D5?14>/;O_,XJ=DD1WeJ2R&?X5\U4Wd1QXfRB.:&]V4(S<gHeI,J&M0FA:.T;g+
BSGA:MBCG=MEa(S_aF,SR;LbfYAR;K;/?IJ\N8;T?</PEF08AgZ>YEVH&NS=)N;:
4#4Jd&+\C0R7<1-.9[g2.HJJca_CK.:IHGc>)ISA/XUR1-?@]IIT-U6,_=0IaZU@
OdL1X7aGRH)-F5cNd(F^Y2a/62d=GVfg0_IgI^G4F&2DM,?5APE9PPJ)aK;[AZMQ
JCfVW5+(04Tf[<A#W+fW/S2>JMeL]D0G^;WS)GSB=,J.;0Ob^&W0QIA@A1O5gbQ2
E?7dVG67KBaPN^4&G+#FOZX/Q]F.e6&G+JB:&9#N?B8HS-SAX\_2:5?SG:b7b(J:
O-=6K[H=NT=-aNUdQc_WXU>UVR;V_DaC8c1PQaP1]-\)Mae;2d#NP_Q>5[C9.c3H
O(4<T4PB,feO2HEB;L39TYHUHc0Ve+Qd+=_.3YdXf4aX(P=b3S=OJF3[,=&Ke^GK
K2a4Q#8b6:I\\\Q9)G@D1O?3fAG2O[ERb<H(f]S9DD\Hc=B3,Mc&b4X+&EHdD>=Y
Nd4&bZG_;B?(D#7C+[@U6EOI.T=(5e(d=^X+Ie/3Z5^e_baW,34F7b1aF7B.^E^d
8(7?JT+4]OMZ8.]Bd)69c[4&^N1V[P?K)^O1YTLOZ;,D.<TX3U=LDaS,_D,^OI^a
()eg<?/DMS52#/\IJ)&eQK[K>AfX^OCZJ+K6QIP&Z81fK=73]g(Fdf>&]U)NbLZ,
#S2)MZ;+F_25V(>.(L_d21X]g3S[dM^G-@)CN4<W?gQ-?)e:9D3#DCO^g;gT,f)L
Q_/R(SOFR)b].XV()3CVBD?)ZS:K(R9BJRJL<8X[X;Jbf7bNPMRZ13J/L44I\_H6
^[:II^FV<0)Q>JU4b+@Y-^4N:NKN]QP]@<?NDD=1(YCQA(QCEG+FfRa5Z.J0cH\<
;NTEP37-_B487]+[ZDFGcP_58^)RGUX[@O0[Hd&=ODJH>Fb)]aNFE-ESb.QY-]UL
X:A&cGId\OQG+Z)W\B;\dN4agHdM.HN_KS2MG-Dg@PPQXKZ^g0^GKL.Y=c5&L=FA
QUF+HCfT^J#6@XZbDg)Wa.1QM^CV-=\CP](D?9]I]a2--?9?bFHTW&4Tf@daHS?R
>Z+7\>I[F4fg^D,X1Sc6FJSgCK9G;VE[P12F,H40fREWEcSfe,8DbbGGCEIFHg+)
6>-d]6#(EAL@,^dP2Z(,KG^b7Z[JA2ge_L,g)ZE-J8#TebZ?E1(=b23HG[;/0(2B
:;_0Ocg6_Tf:Q:J:gRW[K3+CFWZVdP2L)(Sec2OX);?X7]1Ic-AM0e3(FO268a^Y
Gd1MP;<Z?eHM-O+]&:8_+;(Q/5I8V\VU08&BUCGLE;F\.FbLZ5.)_=7[bLfRK#?Z
C9ZC::-e=PI:/C+#^\TZWP3;?fZH_FD>=/KOS(]&Y6V9,cd>:OWT4fY?IW#]LF\@
Ld+Ja,;:FWMJSNC4Wf2#PFC:P.6XI<U,9-#Z>_M(2[_ZWSX1.2,ea&2b:a@,e_ZG
?LQSX.,MSD-4N,Oa,GI=1<Z4:XBM_WW=8ME;RPG3c#NfA1/C187ZCH&:?H285XJ?
HN)<E\)7(PfE0?Gb>A>SDY4T@5+WgU6A+7X;;c4(XEc7AT5#BK?XESV(M2S(1QR,
.Q#L4=<-=1Q2J0@>\SDJHD3Oeea&<f&HK2<U/X@6)]B5+/_@@L(4T^)e]T)1#I8&
\WI/>:L4AN9A8:d0YPG/bFL#bX07<c0OKWW2763II51QI2bGGYb>J(Oc2dD#,C&)
5&):)G0Ke2N#OTF74WV3FJ[Z4a]A01PWaeGW,^TCY1.,2\);>)5(#WG)QJWKQL)S
FAUFd2>eMSY[\[fPLD[GOb)?aC7-e#Wb>#Rf)<9K,+R3\U1_LF,[/-_>dSR^ZD,X
=[HK]5#:T4b71^[?JJ@9_gP,=>ROMQJbg>.JQc;2:,?[]11IRA;ba\+#O1?-(gEG
<97R-:12J#KaK:#IUU[KE+,Oge0.4U-&NZaX@5ccNa]BL&6E#>8MY.O=fc)VQ3?F
bYQSYSH554GBO2J-6:DVC##-J9FO4]=F@#5_EXU3^Eb18g348CK8NV]Q6dO\JILB
/?//LJPDA_[=e<?XRfPdWV9X3)aM@BR]=)@Q@d)HQBP2&Q4RWT5=T\RK8ML:fdN\
A/-B)A.)B8+3)5CP<Ff,-C\.MJSQ0[JbTWQ2HBcS)RA\/ZOS-(-&FE0V?bb#8a8S
g#05C[YBBJ#=eGXIF>D3Z-4:f<ReA<1fU,RB2Y8Y;C2N@NPFGZ&[].K[A>&,8;&<
/d#4W05RK]f<BL8J;V#08EHX>LC2/b/34=8UXEJ4E4D4<1<3/GEcgeTY),1<Pb;.
62SJIC/T,b(1U[I8DO:J63f<K.d(J:+LY(G-B,]=^+<JN\@QU62R4UFY6\?V?MZ#
4/E.?aDbY,6ZO4HY:S=?KV4[FNI3d^Z+H6Ea3W73O.]#\g5VU-,@+R8(N/6F-JGZ
5IIH>c4Wg=-V4>fE>/-;WXa8d[,E\dK2(S6QLK.SdL&.F+5ZNCW,3T?Nd]-POX_>
,d-?+9]47LGT&JKH1I^aK15RT[LPK9@<D4#\:=_8JcF)MRcTVF+ST]_ZE)_ODGfB
>c3KP?c?gU4[_[?5I<2/8KEG?2RPD]P7L_ZZcD1fc#<R)9fNG[-EH.D@T\X+4UgJ
S8YF\+B5\+QLWMJZK0FL55/]D[:1YC^JSfAW0RDGOY=<d8TTE+fG:3T<b)+52IG4
EEZ7d4]8U4b27f,L+4TSX75dgdHZD=P#CMHc#+0:BL3X>GEX.?YKgOJ#-Q<-Q=eI
MV]A1W4MOFe[67OC[M1,3I&6(9I-.R0e4PYM-/Y-Wbd.7I+&[):f?A@ERN5Mf56f
2c<f./?<ZA.ABX(OG<H8V+E2e7Ic9^@MYWS_22IaKB0-c?:X8#XH5H.0A?HOTCYN
R.O[9fQL1D#_3aT_,<8L-W1c.TDC9RXGS86-Tegf7;5>#L=S.7XUX7X[\RFHGAJ9
eK0?0FKVIK079EJ2\60PSW+Q]P5GgTSG/SQ3+Q+U7^4#)S@,V>g^SID4Va@/_0Z4
=f6Y0U1]AEO_TX:&H&@KZ0<1]c,V9bY7I789.V:VWb>TM)CX;1=;:IJ3VMW6]^;E
:_L[N6&/Zb?+@WH0F=7NaY]SQF_OMH3U)K5DD^):VL5E&EE:E.M5H<EW]&=U]\+f
Y&]f67dY]7fbNMeGO0MF\B&(Nb+UTVIK?U,^[DT,>@I/c<QW7UV@A7[WW6#U9E)]
+d3gZ4=EaUQ4[=a/4F260#+P<0cS(N+T7[VF;bV^+d@QB28]_Q:F@/abW[6^da)P
MTZ^>DR1[A4FOb42c<#_>(Xc99b#(/6WDVb]/>(/SW>9I/A6IRaM?GM=)5Mgc6d<
IOJF_.EVdT/A2I6LI68:-TYDdA4VZ5d#E^YOUW-B^Fdg04J7ZDeWYA5ZWJTee1_6
.gUYSDI\POQ</][0#/Y#WM_a<VBLfP>T^-AQFJA+g@0V2X?#^6XgSUP>1ZREL];B
KEZ5#6^Q+RHcccg>]4K>#QQZ.P-LD9\cTR6:<>KA[23J_0d8N.gPWUTGHO8Z[5]C
EP7<D0/)<NI:F;JP\DE/7E1:BgZ]VESE>Z)&-9X4_f^WR(IY1<C<ZgT8X2H/a9(C
fIcJ/Bf>CNH9b?H^824dRf,;19]NN?<&gU4[Q8fW?-\H3Q?LVfbI0D]I^HHKPMCD
HL^B9=ANaHKC3.,)N=S;I,0AW_9;;A?=a+WYJ(EOHZ>.XZ(ZALG(]E8FOOBD3RR\
fM9@#RN4Y(>PeeSE]8g@NEV5SIGG-=>&2]&<Zc8KNc7JK(eZ]0[S\XPBWNE(]>R7
M?6JFV<R.]@(BfXWQ>B;I\FOOaeUB8a)bNGYb8QA/9WR[KNEYJ9FN7&BD,<ZZIb^
^c(aX8HHY1+/82FNKB7g9aY&OT0eLC5QQfNF@<+CPSECe4gZYASMUR]KKBfG1GY[
./eFTB.Uca;M-BcS3g25J/^]S>:03?b>TQ;N[R.d1@fUB]=TIV5,N6Y(.B#1TBF0
9+ZPa[KUBU_USISb@IAMRY42@<3(I#=<;CF#7C^Pfa@]e7(NV/De&aM_H0ZP2RCa
]0a7#=RWPCOH\Ad6TWOT:(K)HfT8d5514HPJ0X]aIGbg/7P=3@2[6DZ<a]dKfK;P
f0OH_;VRcEOb\EKO0,4^?<:OG<cC,N<DcQXXO_ZWc&9#1c1[GK9T>3W3Z6c:)(D)
ged;O@Ef8BUI\gMV^BZ)/R2T_@H5,Xb0WZc>D9V6,T7#PP@@)WfES072^5L1K.DG
]]W>&51Ha<@a#=(/HLJ27Xg.T_Z1A;f&V6d#W7]]JR/&DHa>f<&PXgc7b:]EZP?C
.X1=N)e_05M:fS@Q?IF)=5E5]I6Z14(cTQ/,QKW5BT;)I2&DBV>&K6@e^f3YgNF;
/8KPf)Z6W?d^VG3BUS8CD]NL4Zc/G/\D7P@=9WeLVS/IWD9-:29@B9I0DWX@19_9
2XHSQ>)UDI?8,?L54Hc=Pg(^c&]><D\Q+[;PAc:e<,AT&f)&[83LVSEQe81B[DN;
[VY5JVC7]7g33[QJ^,c3>?WFd0@]RT\W8Bc0>e/Kc;fMX+g=6IL0MIc.QZ4EU..N
,H(I>]AGcOF[[UJ@>3=.B/Ig1J^);&,I(=c7HZ5J8T>2J6bbe@##/a&SKMOK:/_C
CHR=CeD;,CJ3IX=&E[[U]H?-\)I&g)_&0:#]TOF2^MCD]5<C1^S1YCTLUHTA]W\9
b\03J114&>0.d\9eO/42P^2]b830:Xa4J]S_-Z=dOa7fX8XfSPg]I\8>SCL)SMC(
57_d_=TG(>SM[Q^fLWY(1Pe+:c;.&R,P,4ed?H/cJ:,KJ+5XMb;G)N2\DIVA<HPT
TW\8ME\IKXU>?[XeMISOF8KWU<MM.R9]6@dA<,JU2M^J_7G/2UXQe/9XGS-QJJ40
E5T+Le(?V<fHOZ9YeXM\J1,)EL#^Cc:,@SU>1QVddE@3C;)B0:9.,G8FTD1\,V^7
X]:PEI;6W0SK6Pe0M&cXE\1QB/G5@6<?b9(^:aP[2^?J2+\-c1[5;)S6dVfAH#^(
?EP@_[R+?_VG(NYPN8NXbK3K,W2DXG\La5;MASN4<+AQ3ESM^M,##J;>KcZ^H80+
&B]&f4BC>cUb<b01H^I8Z&7[FXTRDE#dX.EeEP&JaX)Q2>9YM3EJ-dcM-BAB]AN8
Ee)g<P&JZ@(gZQ+W[@+DL6Z?T>H7B,/[54NKXRR>:bLQW[V?OC:&_0;)2#9gc^OA
LWQO9cd_E]fW<TX&()(G;@M=d-+J\]^(_8V_X.c[3>>R<c=5G#,OeKUGQ,(T-P.J
?MQRA#YJ[+6Z&0Be:\\::8[^CLQG-8]HT8Df-SH3OPBI3HC#:]ER4O,ML+[UBRg@
462TWQ>:EOQ/>_OY@]DBVbVRG_dK2??V.BB-UP,?1B2g8@T(C3?#04I)Z:-X=eI4
-^K<:5C-R6H<(4.L-?2;KI9N;9<eXab]b?@Q@@LF:R]0UB3-BGE?GTU0MNTRad.H
L74&#EYd4;)K^G\G22QLB0=+4[A]CcJYX=D<OdWT&09O@QX)?g;CH2-7f9?7=;8-
fbG9Ed<6DPT1,[I@gQ-X-VbWeXGbQ>OdI>\D.#U:O>;ST^N,62M3K)@(ZZ)=ZJ&-
ST?>K/<D178QNdS1B0,N/-GTI<#4g<HJNC3Ec0<&e>(QWLNa@7GAW?YLdQ&()gRL
5gX5L]=XW\-GW=R)^[8EX#G#G,[,,CGea4=cO.5OM;a770bS[>X#OAc9X5dO1e1E
CEP;?TJA<Xef<,[+>feDV/D2YdA5--c&C>8bR?^0V5AZAM_-A9X[Zd;P47DB;g9O
d+9+6UUVf)&^I>6HXB-eMG2d@/^9Bb-4]NJ\##R^J@;>A,7[g/_+YH801T8eH9@4
Xe>IZ4\93OW@@74@?aVNU9DU?GN&;O.Zc8HGZ=G+g73>L,/0S0[eQC<T5HUAW?)#
Ug6c:0HB&L)EW=0U;AB<7.GFd4g(g/IF+TCd^3?7_MeP:DO]\?cdA#CSdf))L.5<
LGJ#06cGB;MUZ-&Wfc:B;NB?0_a7E36)]Ye5g9cY>fE2VU_W=]XK_B&9V]&-BP)[
SeW/]1(.@:>+SR6H/\=#G&=-=NP3UJ2+47(7X3cUC><dI9DJ+eTWXQJ\R]L\MU4^
MH\+L54BMc0T0.3f?7/6ZVG9989]eZRVS9E3:#B?N+^15BcF9)gZD7Jadb83>JBX
V,T#BMBa?Rf<E\\NM:TE(4B0NZTc?XfJgW3K55McV^P?d#/eOBVR)=NDISB@-c:+
d/@(e,/3]f4X/7[d[.c@:CN+7N6.IF(.CU@^0;D8+QgZU::VH8a@b;Y(WI^1C.ZO
9K?IT^T-XI4S9aFC1OH@2VZ+//;MU\0L<\EaQ+3RJSRY#UbbN.66DGF00ecLWEVN
P4CWg?7Q>]RYd66#]02U63LK,d?([BDF&&#K1+?Y<8&PeXa)UU9E]^E9&c(4SNa1
A-YB6Ib+P0ee@@3c=</,#H5WeN^88;N14=;,Ff@X0@ELSQ1]C>QAe3U/REAI8f,8
DWK165YP+f554GJe@DUdC)<A>E/1N(,32B&<>Rd11bddL0[0BH=[0G5G;+:84_N0
LBW>d,1eZ-H\29([?8V2MIHVC4<AW6(R0/aO_]2f8+d?2a37W2Wb847Y6;&g)-QR
W=Qg>\8#8C7-fOTV@?7c4&9-JA69DNS;4a[^2V(Y5NTT\UUSJTdb)=8(QJH@IS3T
QISeJFBW[#ddM;e30=/#DJ^73+.Zf]XW[I>eOJ.B[-Q6M8?LCUK/Ya-J).cg+0O1
G\?[KN.22APQG&-Bf(#A6be1/_-ZQX:I?>Pd9IAXW+C[<Re:C,?eR5E]+U>2X&SV
eRO]0-a(g>]9Gb1VPYZVY\=L+FbRJYc_H-6NgWM2_3VJ_4NB^&-aI6WJCWI#OV1T
TT?+#LBIFEP3X+]5Xd/+2[T;@&CeF]CXB=Z^NQ@N-TBg9QD>D1;4QNf6R/>/0WWJ
aTW.G\>DbIO+PU8&7<(BQ>DXQXc)KfEYAYW+g\Z,4FZ4,P\:_IWF7S6Hg]1/#FIO
&5@BgaeK8MAH\;.@+SE<56TSQbc<^]<=TP/>T_Y.e]EQ]U:a06@F/Acc/+P80-W?
T.dA^QDUcc+;dO=TBDedVA1,6\_a3)eX\d1F#-[KRMeI1g^UVe4T5D)G08E(V+78
NPc4A^@A</5F7[15ORYHFB&6&fEe@G6_+NR9NBC.ZI58a7[Dg/7MaGYKJK7.8aU&
Z]ZV/[))3K9+V7feZH)J8J>.[cL,b8N#Da-3f-MGaF:GG<]ENcATIJ:,<ag-c];)
PCV[fC-54g(A^8MU=LJJS02._d@dKZZTLIa)(P/:&@RVTd&QWa/T:KZ<cD6;(>J4
ZGAXF7S/<5c7)M/9E1fP]Y;[L:a(\]M+F^;;dgaCabf/Ba[X9A3d(T=97NbMc\c-
gb>BeT86NIAJBA;GM=P5f2LUAd5FQ/@c,YYQKYBg/AV]6aH[<<0R4d)#)5]M0:^\
F7E-ZeMVc9B1cM;ZQWA-[Q>E_91Jf36Q,aNNM]D_1UVFOG/45\VY2@ISDgAD6>&C
>PF8O:2Q:S@M1T:C=C2D:IRG]6.L9M5?eA&U[.2U#,=3Z9\<R<.D&g/)Fa)1:>Ec
>S8(gBZgaWQB,KGW7X]Sg/L5I^\+KO2F<?[FMF6^92e]+IEd?(IOA,^6YI<427=7
cQcO)SE1QA]+S&U=6>dJ&6LMFafI<]([C@CdQ84[XC)7fFX5RZ(F:X0@S7QWLN#W
aK#Na/W,b[>T#=4S+3QNb2+;bA3+Q:4Z.EeJEDGF<T?73ETdZX1WB\[RQFQ<:e/B
cYR,&@f:ORYcb0>@#XBOM5[G@\@&I.5f49)gU/FFL,bR;_5GG:U;d(+9+S=8Lb:V
dDM:PeI>7_V[:.aV-(dT:J(H/W>?LE]Ef0K56b&/Q^&&=dMWCFKRPBL/->B2;T<&
eSfc)_\&2:@M8QLcgYMdV)8AVe8^G,__c+S<2@XALBPU,B_1f>AGe\U,:<:eAMZL
dAR&?@;^LG;e#828Eg;.egg8.W/G@-ZVdIZV&IYLH]F;a;YV[QZ(DE^D,LIa<XgY
]0K5AHgNGaL<(BFcO,<#?K.,4EB+\g_=RN]53JR6OP4JF4;gf^9P]\/S7T[E,+db
N^K25H)ZKfc[_T+./^FQR3A8+BgY-5g/]]RL(.>Pf6H0MdRHI>8:]G/WgD:GU<2.
+Ac^4G@X)?FSQU+f[dUM<a\^4WbZTVS:H18Yd6OMI5GD(JGP<8=:N]/M3I<.0+T6
ZS=/Z/&8A\_J>MXY?ZG5RY@Le@)CEgKRGI&DcPf>)VaafD[>)F^,C5b;SR:K2FSC
gb^NR@E=.7#+M;\AUB<._Z)gUg3fWb?=,;#FP=/.#;O8:QO\#3E<:1O[[O7cPM+K
5&?DFLea7KAQ.Ya8#aG2V[:VHf4C/BMX?E50Kd)/ZB_Q([_N-@3@fXLT?3A8b=#Y
GY,PSLW<E3\)M2ADFGTg&X)Y48I0ID7&[\QfU53S@77ZJ1XfF.IaB?\L)aGITa\>
)#:\7Y\G>;f#,-@TcG/0fQQA<f#P0CHeJB7NZRGDZ,a@=V4g):]g6M9=-Z\0KS?P
b;]5UE+\^e+2I(2Z24d_@_>&cJ0P[0/R2e@/JE)6Cf;YbWJD=[T\1H:R9+;fR(];
+7=XFD/e<9N8;&6.>5K7M.K?J<9&aU4PE2_=>6f-)U9dN/&GW(fO^H#cNKBSCbTK
Z4,X-=a\5\A@S3Ie:b^RN#N)^^Y.#AX<7D0J6d491WdEcPgRd->d)S&YLeeOM&/R
9WF&d4&=<fZPaDU<c<&1NKIVQZ^J18gB.J+-3>.5DJb8P8V8g(N4a3aJ_9gb/[,?
/S3-f-G#GZYHZ?E/^W;V^PD]01X_TSY;]CTE?#HV7Ja)XTG>B4T&@V-B:Se3(E&,
bY51B9<DHb\/YQ27EV#W\(X)OS@_g=^7[ZEH^=9L;&32JG+7H?RPfMQ@g;(\-D^K
V4SH\U;[&A;J8Q4,.O)9H76].d_7]4cV6YbQBOSbQRCGe6\OFUFPXR2LZ-[VDB[P
_8C;37U)V-Yg\fF+@X1R-2+\>fB<>E)&-HgU8bV8U]LL.BfXB@d^cKU5.=H1)888
?2f;<\L;]E)H1FIG<YAJd[\A-eaN#=\^<c4-S5V?@J5cU.RGcI(=LV0,F#SV37^V
.eLEL+?C5(.I?#H5FXO4./NbXNRd^2&6&[FZaXCEE7M-/>5VC&3<a/EGXLS9>=U&
YN;V+V\SK#&cEec>KMDEP3>7H\MQO_8UfdU>.9+FNdM-VQX\Jf7?@a-Y<+]MKR[6
[cP/A;SZc(=]O.YVbJ@ZJKAF[@9,0&61ccMIGC3\W?31+eT5D0N(_NV9E\cXIe3B
N-a)2&1Cc74.(Jc=XZc@Wb2OM?EJ[FRbbM5Hb0I1d7R]U&<S)bMSM:+@ZZa^ZdB=
K=C.bXBJY_\AZMW@0S2<K2L/7Y,Y0\Xeb\@XQedD3M2IDBC#/XHGVE?XbT5V@6A[
PD4H@B.RV3[5CV_^#EfR8\AgQe0D.L_ZS7O1?gVIbMWSBOdUL7HCIT,29BXZLFFL
DXDD6K:B\M[-fd0Q5g0AR/6eF9I92>#(2<H1&RULR:.SQU:JfN=&6@gW_EJ[9>-9
;/2[]2/N1;;^5ZL[XXHE(4UR#db-Kf2JBIg_Ye_;^R+B4ICL(H62=(X[@.^a=ecZ
(16dH9a]@8[Z]A>\OIVW<Rf)CK_;9<Y2ebJ#])=R\O0)FAfEaD1(A?7.?2H]?I3&
g@E^Jf0GDX.g:/9[;\O]7dc<MT^M2GD<D4MC;YREMBB)Z4]B@[fO7WSO[?XP)Zge
S_.1=_QC[IcZa:2JJH@T<+-FX==,WJB9@IJI9L;<JU7H+OW3f[,J:(9MPOPXbeLQ
];\V8R]:(_bS26,R)K\L6NCcb&]+VVWeb>W1.K06PT.X,_U,+7e?YH:#@5OZ(DIX
bML\&Ra8dC_WDFbG#.de:^W):@6Xe;fdB4E0dZDM28GSE[SeB_JVf?[KRcVg9a1N
/a.I,C4H^R>,\D<FeL0;5&>LP?J1R6-4D45VJ^__GIW&V<(GPXJFJ>APNOSXJ#6W
=6[5[?cf+aYZ5=Q[dM=8^fOWFb>,BAdWc#TX_:EXF^=:PB7GRgUM[R.cU,8:e;+7
VQ]C0R.+:HCE@7+C?2a0+cbcf@cZb1:I?+H67XBR6<\EL(=MgX7_=_696f3DWUW;
H>aGE)Xf[+H9TR][/W@#705P<:)/:b?[FZ3c3Hbe^Gd,ML/\Ja6A,1=dYdQ]gCc;
OCMfRbWebN?6&H_EL;d1@^RKM/d,,A8=FXW4?NV,7=f.[Zb\;L4I:Va,=UOD<I9S
\7V4R\IZW:KQ.;#Se&Xa/3+W0F4A3573#5B79]aQTKX@,I[Y6T_A+U=MC:6ODCC3
cD9-)FT#(V-KL(MLa^_?Ae-(Ne@0?>:TO#6>R(8W49+H_5N@A9,)6[;W4-WBGd,Q
a<HfO7#0cX0=b)ZG+F72XX>E+PY)2_fe40U6bE41T3/&H_BF_D;V;E-bcG@)3AU\
Sa[8&+0D[/^a^[\Xc\b4J-^D(>)+DOS:cLdFZZ.P,D[aBXA03AYXaVI?R-+)S>9O
dCWJU=[5#ZHH)OD[a:eAXK(H4W2RLdS^-R6EEeN(=?0P4V\^+57\9/a]cWH6R51V
9Y-d_K79a=DY;PL9HYb/d.Z)6K?XgMJ+M/2^V57M).QRGYdTJ9<9_;G?V;WFG0.,
4aV?O4>5I--)8A8XHS:1fH2cAQa5OKg-].JRJ(PE-e4JG>[T6f/N>ZJ?4F7J1R3X
0W^9^K;:38?E,2TE>cAfPe&e@/@b#^QaKGA&S//cF1279A5CRg2RDWU>.\/c+?#\
cg0VEN6EBf2E6\-#=c^AY0#5S#eV#Q^0?QRNWKD>)_((X;AN05I^Y(XR?X^<f>[T
PcDU)Kf,O6ZK1baaIPKb+K[[&682^U/]FK<dQ2fQf8Q5Wgg\_QXTgT]@1L02M8.e
;_9:)_)=fHf>LWNFBe2\Oee1\(X.>Ab774]7653=U4XgW^#_FYK;EPA16Y.be;cL
bc+d7^(a4bf61>H^eg]PZD/-b.:PVF2+XIB^7dJ+Z<eQ,U90&\-5^<6K/HaN7YT9
T@J>9b>;/?A6;d;gRKIC#DC@HdCg#[beDGKd(aF?B,[-YFBM,CeM;@YFKC8eF6Q2
J3+[[fBaD0bB??-MSa&=_c2X;@+-88#[0]b_:Y(D3TTVJ.#^fQ/WdDDgI2FIb/R+
Oa2^K+Q)B&6M,&:LRL\E30>]T8;-bFY==5A2g<MSGId0/Od07F0R\d5?TDe:9Re2
+/3JC=8#7NfFR):V](Y(@26:\Kf@BIFL4]8I\Pb;bT;9+^68WK@WbTP:?LECf0X8
]96)b9eO\OE=dE]:KGb3PP<+-0YS6,aSgLPVAP34:ZJIaE-GB;7PNYXNA:E)S?A9
SeWcG1[9HP4V32<Z,E>B7)HfC.(5g?ag./(,6g>^,#\6Cb-05\+RT]41dKBDHM4f
LMcYZZ+CU0V.1<?Ra/,X:JSAa7HPfE.QTMX60&GSa=6WgI04@Q@aK6=@eU.Q91Ic
5baRdAa#@f)(6H-<C4X8Gf8N:-EQ-F8R1[6_K--,a/2:[f:Qb#\E^7.]I6caS]]8
S<ba<B.Y(D=EK.)RZb.6T-K[7c_E&K1(#FQEBBBDF&g6XT=9fFFbP(BcX]):O-9d
Yd2OC)@/9-:5I4_E,a+]#<[I#^O94//:7O\Mb+GF)@&5Dg796_@=VVZcN;Df7[X-
(?@g-Dg1JH@(LGERGZ4HGYLd;7fgR6U#EDNMQCSdLD>_?^Z:2G>&MKO(3YVJ72IW
;72CCG?[=dB72RPV5e=N?-P>#W?YI;eO7&DJaA=QKWgf[-a/06f=<,B[10\\,7P_
YE?cC]:AK32LOEUc1HL/0gCR?MP(ZA/#6<<@-W>AU3U:+#;a_(e<e>KObF_UR(Re
f+N+CO;^/0Q3c/?B/_)22?R,,0.5[O6(D,1A>ZXA1]24.MRTWNQ[a@L]3UH-(/^Q
.2#La7(If&f1eG2-XAC+IVZ.a4VIAG)F6f1CE8\O3@\\RGLg?McUH&MgGDaa?FFB
:bbW@^YOK7)(\U_8O@@RUaT\\[^KYNR[4Z/J.b\FJed6?D)_[9//Yd16(1/AX;D2
[.ZG2fTJIH<))6J#40fQcLab+^X-;SQ_>;0Hf#)U=BdI7&)-0a_]5H&7FEOf)4/0
7C9KQ8ag06R3YS1Fd_FR.GR1,6fCeM,CeBZRU7RD#+VHTK8\8(e9Gc)9c;<YUIZ-
-a2bIQ(C;?BKHOS6;1(<QU7/e1EPJ.g3]9KH4Y.^J[XM0G8S<HBE8(L_RYH33]-V
)f<[bI+/4]6-7WBS9b8Fc0D75),@SN@L<?Z;Gd=[(44W91);<@W>7CgHLOd?/MBV
.0bMM<FB1AHf^D,4JN7C+NRBZcM81(HbY9#7?M+(FS6ZC4SV+](6@.&8MW#V,A9R
+NL-]K5?IRHWJDY8V+B\:,,IYZ\D1NE8&#>W>V7dfKL2KO[;SL,Z8e6IQ#EDD[BO
68#8efUe0/^;0dP^[U#&&96\\4W3<V^@=;&L:bS\1;G8I?^6YK(]2=UZ2)8-FKS/
4-ZS6eC)=#CDT/L9P\E_.A+^(Dc[]/P?[16-AeZJF,SI^:?RN4&HXW5QYf-/<,24
XO>W4D@+^7/IHgEJ,TPRSg;/IQ3F:2a_P;04B]JS[N5BX+FJ0AHYKeEc8E_.PK.I
6DXOUFRL+)2)H<HL?bB(Ug2G6)UX<_Y@&<-)^&>9\\8NfWU4bBf71g\M.?:(b\:1
Ua4<R5MQfJS/4GO/;bVfJ+WLJJIOeG9BeX0gY24)84KI0:_O4Hd]4<?ZEDWaZ0;K
g(+LEFT7D(C.\<LTaTH/7fV+_^\N7?W>Rg9&AGMfZ6/37KFT32f4MX8/QN&V<[Cb
74G<4@ZQY)dbd+eg^0dVFRB0d&@R[^5GMK:Ag2OP?Wb8BSU[X?F-cSAbe&+GP(V_
[R?b2QWa_-S/WCaS8ZJ0YGb1D6eB?U:=WcEHE,OC@V9Y<\9>U&BbKca]fecH-Y9)
SF(3NQO9,8Kc>E)K3C?b7cA6)ZI_OKcCBQV0UVaE2WC78Z0PMDE[P?+W2G939IN<
4RPcU+>\M>U#;MO]#<R_N#SPC&b]\fX\ADXP4]I)7bRdS96N[\L1ZGTM8Vd?M=GU
4>C9<YV_BaH.Y8QM^^W:&HfK?[dZE+/DAQ;fL=Y(<I6.];8cd]c8+XH2f)4;FaWf
3AbNGX43HH67A:ER#_AHL]\FXMUK6F7RENU8F?+7_ADaS6V5P(GdMJ?B09N76+M/
bV#<=8&3>b@[45F3?fNaX2[YB=GR7^B:88#O67Q>aAB>^YT+5(9EVSA)LS6;#.4)
4fD)P)0_HX23a[&@IDJ;.TO1E[c0T(OIJ2S[UeR^9)4YXgK8@/4A0[VgN>UT-Y-d
)C]ELB9gIg5Z<Y6@1NT59GVJO(ZN3T3,=LQ?@9@P+A:RWC9+IRX;2(CU.=:W:a:.
A__=-DEJIaH/RGNZ@R;M-Q52fED8[-KE3TR>dM=EBg+dVS+,.UK7Q,_3[2I/1;^T
,42&DPJTDBgZa#HJYa[F?MTGc2O^EYZ1-963?><g^G47R@3CEOC>I;[O-7c;(<#a
K9?B]7^.KA?6SK-YH+_IZMX)M_0-@Ia4Ogb;&2((\.M.:4B2G=ZEQ&>=()4a+^_c
DN+e,RbTK.4)Jg8R1-JXR5,8KA0BfDU@[&>9bIO-bR(7-Q4[T=Gd?-MO<IfN7W)g
?OMKB:1D7Y-ec6<OEOBB4)]T-fDP+T/N&2bW(JV25W,8O=)>dLT754SAZFTPK&W\
[6QD5fA,P=8_gH9W3(#GH2,.0-K0dHZOM@f&WB^O1dP0\1X;M)LU;IP_+LdUfZE8
3Bff33\<F.I-,ef3C/P2Q-\0@TbQYgf&0@<M0YEWd4Ugbd?/9_Y.:__(HOO;ANbD
3aAP=]HH91/^^B,#5\=g-1#Q[0FN_J-2ZG?I=Q7OU>E/Q1^=>5)E+;+R\^YT2;T7
ZDMU?L4G_1]&38,U=_c^#S[/3ES]3#,FVWJaS#ObRQ=K6[2F4/(e:?\91YV?CN=C
7UUgQD17YCPaOgV=f]=N0bXQeKE-YV^PT)CJY0[YJ?KURWD/Qb:Z6HV\X\MPC.2E
Z,^P+XQBQFP[W5GI&dRL[YY)N1&-c[a_FM;#C>RGD4a?RQ#=UfbY;.=1.Z:H6O@4
M(cM.f];RJB8eDM,C7S>FSAIR2RHV,-^>V->::b3ADA\QSDY?4b6a_)Q]XY^C>,<
d5-7&2a/dR9XgF-cZE.PPJFB/JE_HAAG[&#OL]H/EUDYUA4H@6H2K]@=>I(cOLNF
<-6_JD1bL7cgB74_/WO\/BJO2?ZF.:P1-DfOUU=O=CF033]14R;VTL@>#7SK.OYV
4JWWZ_A/a=PePF?ePHN3_.:E\3Y.^fS3>N4ZA=TQ<5FZ?QIKLgK:]6I_)eN&[Q)d
aUW8d,D#X/^I5LOJ1dL-##5&+&S<bSR_>:W\U)Q[#3PHC.?_P5bUOT45ffVDef]@
]2G4+X5TFNL5b2CQfDV[1_4CT41g?(A5JKdO^HXDSJDJg.OZQ(-cf[;c48,]G:<9
;BU?;B5D4O33QX>;YI8()W2>KAHB.Y35fF^FYeD,A^Q71-ETEZ\_J?6^ZaBZ_8S>
Z#KVVZRU+A@]2bQ;@;1<+I#-=gLAI<&X<NG@JE<]ZfA_+I3b;/U4;9K^5SSXd9X0
@,e73S&f[#2(1&RIVd@L;0Y3M-39<6/UN?(eZb6(AX1WD1GEL<GA+QgMZ5+Q/]0K
:T<&HHH_Rb./M@b3DGVDQ/IbNDFdMQ?eY/e@Q]D=f=;0)G8C@VPPMP&3a6?,H,bO
5T.gUS)f;A;2ScdU.^^D2<A(WcL@6PWFdJ&S-5.^beVgO](OCTXb?D@^c5c1#Z&W
G==?L-Fb4T;c)II3bG++8+CT+F#LQfAN\-1e7>/Y\aL5S1Ye<NQ1NF7VU)HXW<QT
:M1#Z)8TY,JUZM<Wc-1]L>X;FdG#1Jc)&O9C08&T7D)1M;b8J/bb@(Md-F-B3U?/
8<9(cJE+V(\H19_e)LAO,@IZQUe#?RDKeRbI_GK>QLG9dLLS^,aUf0)=N8XWL4KK
-08T\fH/T2,d>XbUL4I6(f)WQ^G;c.5eTOV.;[-_H[db,[:2YUJ7NbNK@3N1>3Fe
\AgE&eeY^K<CY+),WT?_Qgd)L3C@D6cZ;2/^7C0gZK5(=HeTJd:F\XaBg.NHDH1_
K_1-\V7-]e/J&a_:G=5914#7[<XKbT0eNU41XW@BP7YZd#RL8?b:,=TAM,YMEEfK
C<28Q4f6AU9O:8Bg^P>dYRgBUI-TOU=9KQ[KNYPQRIVBTYc?OEAM(.WfGS_(XS>N
IeJ07_/.bV#ZL18-,33A]+O?X06W_4=K?QG8(-(6cUSG&.cb@GJ9_&(AL3G:M_9-
7K80N=BDT<#+d#T2SN^4(@I;YegaYCUcT3<(fRE,JJ7XV>&Q<UDa^Z8D1\EX.#3J
IDc.ZJARUP+aO.^Z7:_HU?aF?(f+2cRRH?Ec5N)GdL+[,L@9d?>BSeda/&0aCG>2
]ZEDA#NXd:_a_Q3,e>>g&?[+19H^GG]Fd>S;?,>47.B:^bFcE5_&TK:UgH);A_G7
>QE)+:c2e\Y^]3b2-YSHIJ2BB32OZMgOJ76d/0X/]P]P;N,baYG5I:SHVJBLK8O9
<N+,8),?N2g5b7MI<<;6OW?R+F5cbY]&\:I188d6UD(^(Q]Ta^5bMV[d&6dLVE+C
E+^LX,NPJO8>T=LaB6K)EVW;P>&CX>A,SQF=R5P:be#1[\Z:N#B-04HCB.K_FFG>
ca]8DV:,2XC?;f-QV@^,Dg_FYgWPWb<5<eMcXO56?;8P???-5#CT4R:W.PP#3TLW
])7M9WKQ\[HOe;6TMc@I3CgD@0&aJ@#\NXfe9c^Bc(I+9FeFBQ--QA2J7^R=H=1K
feZ#,6?&fP>Q(1M&c[A).HF.9&3G&Y+(ER:g+8WZGR?E-AU&\,U)Tfe7=/@_-2+]
2)cY#@&J@0NZYJ@<;-e#>9/&>+>#0H\+NG(+L#R=Vd:X+A[5N4=W7XDbQBP0SG[&
NQUEI6=[MaaaTT-BgI?^8Vb.(^c3(gX3:#GIXWL<_,B8D+4HT/T,M&I8^bO,W\7>
YB&RN3bTbCcFGYA^/ce@-6G:E@]c)SJM.QC4-JQ)<>(#?9.G,TO.M8NFg<D/2A&Q
_@WK2CZ;^HL8G9a?U2Q,>g^B9G9J/I\+Na2[YE;dOGfWTCP2+:97L9cJ]TALP;?9
9=>VC/UId7^/6S-1@dG46@SAI3+^OE4Y\ZA]SWYZJ(3,(Gg]U\K\OHJ-8S/8#IBA
?Wb2V@0bDG^1<CKCDF9-RHb,))ab7/&N>AJ_-TI_@R4]9NKEd,CS30\G;Ee/L>JT
Z@2];TQ.L;E753Q:2)6?0LW3ON6+YQHW.T\D8D]BUG<C8Z?1FUV^Dc]d/\@4&0L#
bJ9761f0P<W2ER-,7K=&YF._S9RS;a)YJ+be0GaIaMcVW@P=QZ47WY1cE[V/GKea
[4R,@7A)WHYIT(S_T4eVAZL=YMC.=BV>?GNH(Jf3WIQ.G]E[9]cG9(R_ODDdEZ/a
bCb1W,X(ZH@=Q&=SA24-Z/J:FCX4C5A8dMC^3\8f6c\b5K]c7fb.Y;P0@ZFOTX^c
N6Cg_\C8QM67Y+(\aA]CXM\][UALYQ4bH/7JKNE@fWEK_4GZFV=Se_;S\CE32I73
)^+9MdS+dbTJVNDQWBN^#WM7AXWg<f+bB#8gD5,-[MH/M&F,0+E?VG[T60+EVU-D
0NKP;K^RAc0#bQDW+=[P0[XTTP0Y/PaQB:=397]0;^.Kd/0a[<MdVQ5[0HW?ZTQL
LU>1R_9d?0^DSB>?_e>=.7:)RDGAA#;\b3<gD>_L;:Rg4OP8(g]=e?YCe@INK[N+
;I_CF4H[09^[I&b6&1^#KULe<V(3RcEJe@.dN5VfWB8)e;:NW1c]Wc2[cLca#&,Q
>e?3_e7+CX^fW-@ZAbZ&A[&X6TX&gM;B]2U<c9]X;9fW:LfP:NX?C&S^eE^QV4#d
<BgbONAQNP9b5CQ6:g3WCA>QXGSK]:=(S@@RbR5]N3CU[LP5-&1b8\>NBHf8L-&U
9G.W(0)O@b4IVf9W3Lb3c\EYY^H2_P\IFEQQ\O?/@RBN-L_OU;;Y3?:]USbL^QK&
2,.GAYI@gP[V4;;1D=[Z&KL&fV<LdR3?^YD56b#J7C-a+:;LRb&V\&-Zed35dd&6
IIfJ;=]167;QLO>)T:V=U],7#6fT_gKS[(KD8=LK(#INO:M0Y.\I4XTE5EU9W.:V
UBIeE#;Y0_SZdgWRcb^ZbfJ.I2U[HdTaE;#RR?b\J@>.GTfdI\>2[8Ya2K\ZNUB?
SePT,;38.4Y--I(dZMX^;).3WR)-:LY2I6[N_RBQ_V<O.afR=^=3cA1TR2ZWTRUW
CCRL:fEgE[M2409fa>b4/A;(AR:d5GcHVFP\D7,\4NEOKYEA:3N,8gQF)@0T>F_J
Y#_44,@\E9c)bF]>?CKJc2F&#@cKB7S,NNUEX/Y0UY#HV+D&X/\,d39K]LDd]8HF
>Y)BGf8JgaW)N5&5fPeB8O>CSVcTaTC65a5IV8e#5.77X^ULS/d>aCYMb/]@V^X_
(\AV3[<a>cR+)B]N4\M#N/E>[;NN5<gOE5B^JU;R+L&_a&PgO.D,Rf6CKC2A7bD,
fX:b5gENW,Feg?SMV6;#P7N[=#)10#8&MGH.PNc<5OBcAR;S8Sg(N0NB3185_XZR
BM;A.:d/d<ZMLU2<K8N7]X&>G3B7WW3J@3=ce4+17M&f41cNK1[Z6eKcaK2aUFG2
OLL4-O[?55TDM:d:<<NX>]DKg2U8NBEE;#/R7K.6FP5\Q(7K+C@(bVgc<[)7/,8g
-TY)SI,D>?9XL+61;^eCTWeDe9/@7+]_7.LN\Q-c3RN(Q=?a/G<QX:V/WDT+c&,;
083,Q0LYPf]-8aF:PFU(--a>K5K_CQDR9-0Rb>U)]XXTScEW&ee_5V(LEZW45#.G
\Y]QY9B0dgZAGLc+M9#/0:O&\KV_#8^P5/dH9V_18A[#)],3G68V4LX7-O5J5@f&
KR#GYHSfdLJM,B_I<d3g(a4I@A/3-#2/9GV/c;GNNUE,/KBW^:>F>F\]JXFg[A45
^f4&//^NC>NbNRP3V@^Ue5JbX48H2VSP0PTZ1-PU<Z)9H>:MMG=KFI;FgU/DQ.Ob
]=R&46749a-(0.WRXYReYcHLg1CFZ7(15Y/J@T3M./dQP3_50b-SK[6O\Ee47<ZM
JTbg&cBdRUJHM=Z^52LL&gY-bZRZe;G)J21HQf9DbIJY<V63,f\f&HPBDN0c^C3&
0eUeLGOe6XQ_VBO1F]e6\aQ#,bW29]&1UG3NcN]KEeD^,9aJ_SK+G7L8[7?BIc+6
MDg9eI\=L3cb7?^SCFOgD6/_-(B>HN?2QI.ITH<F^2.H>P3cAT=[Q&\1K8?WN+#<
9c+aEXO2)8(6=T2BYE5cB:fVZ]TJNSZHPLEBbA;\VWX4C\]=[1@TfEXUXB.VM6a&
XJ1[D#H^PF;=e8A@H:,MH;A>;B^RN(78C:1E<6ccg_U\YgUZ\)#9D]09DE7P,ce(
5_6>K?C44bf28&g0W5Xa57N@aX7Y+Ub-<XAE@S\e#:A#gEG:&1bR\:4gHZbFKVJU
SFSf2O^[&TO25#61^HC9#c6dQ[;8]HO_<ZWQNY_#;\U,d9900LEVB,Yd>g^<_&5<
(6&;4fS^5(9([;S92J_PTV1C7KX\B0)</408a2;SMFN]NQ#G6K;HLBGL_aG]76ET
Sf#]\QW_XdFU8=X8YT#eIbEYGN:=Y&df7H)EFa(1VJH.V>W?FEV64d>>XUFVL?Fe
E\/I&5JJ[e=g9ET3P)=GK6?gA[-6E</FKZVUDQ(?bb9+gU#]J1fRBUKcb4[aN<GQ
HG^^C9FU+?_Fe/<-6,,1+T?g4$
`endprotected

`protected
JC).L44GbONdCFB@K5:W[X0)Xb=^TZYb>8X#(.SO>c2OFaR3VccV/)bB+K/T/;^[
2&)^OJ3XNM3d.$
`endprotected

//vcs_lic_vip_protect
  `protected
5J,-?gOgIc0Pfa_;4IYICUO?)L^[CL(UQeK[KQ^Q&E3d,,)DZ:,77(4JO>U;/_Ab
dO:@,NO8/?VR_0Y:N5E1[FRZ[PVD9]H5+@g-\OI/)<&MGM7>3=1#eII[76W-?R>O
ZA6SK#-D]N:#eMPf4?B16e-D?(Cc[e5<M6OGVAJO#T[bH[KML@4EF7,&&&QKB9.F
JFZ0/5HcO66dGNQFG3=7A.Z@AUP,B;D-C=0B@(O@KK>9)UH]M_#F?-K,67eIEd^#
)f^2US9(]c2agVe/a]+3VMMMUNbe>E/1gIYZT(2;gZT4_+YNMW,RK.5WAWC4dN6P
5,8f:YO#Q)@DHXd#IE\.QI(D&(SaR[Ja#g4W).[J<U9GG,>1FY\Tb6+EN?N7dNDW
#f_2RN,7bgeGCQ/Q6L#@+c:CP_cZ.c)d_eOK>],^.f1)+Q^2:+:6K?2SZVN]\Q/[
CM+CV0]1K:IVT98FQ93HZ^SZW)7WX5ZaRO?><>OJ9=UF&.MRL5U/9^)Gd[W(MAf7
8G]PZ9aWR^JN<d=0gOF&0_GZA9fE(3JPA)X+5K^R:&422++?9[SVaGB8\)4L)BC6
a<=Ec<HP\O+4CKON=0_cH6YJ^CSM>G:BQJR#0]).@[ZdG?N,&9Yc]-BTDaM983bg
F=WD20J6;GYYbYdDa\NBZ?7JDAeEEGF/O[dT?)YYJF:Qf3A9N:K:0OAX2ZAVd1^b
V7.3]JABZ#cCgK/b2^^He\UeR]^E^S#;I9\HJ4fLVbAIL.FW?8[G=J>_f6^ad2H4
7;B4,b+]9QDUV30XHT;b^0+dU@AC7H^aAaV38Ga-OS0HO/H]PI2KfG7<DZWTSBfK
XKd?4+S8]f2T4P\:RD2bPUDaJ?1J-LR6)LM&=6Cg[<WO;D#fSb:&VM00K+(Z_bf=
X09)6Kd[5V=D,OC#?@J_?BME&EN<4TDI=93Ld8&G7\6^QD4&\&T3,).1C<S]A1,-
UG0<?FO10-,>_IGcC^AG04(R3f-aL#UYJ+R\S\MB3gQEV4C)E.5=_Q@Z)H=)4^gV
G[3AeT]QD&cHX<_#9d>,][-A13)\Z^\2-7S?4>@Qf\CEf#XaWAM+=.B&[5LQ/BR2
RG@Y\bVN^,<gN60HDZ?A9((<b1Z8X&DQLL42WIeLA1LT6dT7cEUHG3&YdSJTHA6S
>@D]P-4LSNQW+FK9C^g_>84gBCJ1d]TbG@;IB3EZPRe<4GBb6N-1JFaC=C&4SK5/
KD;;E6K\Jb[;:dM704MUOH735&1VY;K]D,g6[(Xa]UFR#(?Acf_dB#cN_aF]^KJ-
Pb&1<+\(U7P&LYXOR<AfDTA[G)Cf?\U?3G:W3K.FXN5,7H)00HQ6^;4U&3#91QOF
U6B+@?<5&fe(UTP@^e[HVV2;f]/Q(8DL.+RL&,g0&[2TM/L/Z&IJBZHCT^&20=cM
bXXT+0UTU5bLSA5#QY3X=W\BFQOIXfgI2>XgeR0C>dTIQ^X=a][3>Y._<1DVX7XX
J2RM>Z5&,BA)ZX<0.Ha>HJ8D^WCO9.9LR38UXg<[BM^LU\QFObZAZMgT#S0_@KS,
>Dbb5KR1Q@=b]Y#M#N_HE,JEH@d>-B_X20,LZ@X[^35P]f4gKAIUbSWP>DA,8G3I
(,+T1Xg]CEO02L]Y/>=_L/9OWEeCP(8_T03Z061&0\NYZE^YR3agQ6<Y\Q&C,BZB
2_#3g2;UPW1:YSK&ZVXf4Tg4\cVcXC[\?6N#_<./BNA,CYbe-ZCVfY7>=-#AO\-B
dE:fMN-W>gF\9Y699O;bX9.f\;#KZK7;cQ9ZLS;B\#NFd5;\<0YK2IQ0TDf]a9Y,
--]:2I85H95>>KR+#gJ+f?:cI=E[c]PM3U,UdW?XaLZ+BAW9<5(#06C8-&/3\K3D
Mfd.BbIAId#/LRI(^f+HOVX>cQIG21^;GK<E:C5:b3a4U#Vcg38eH83T3fZeB8S)
[.+1]^6e+IafQ=YPNZK[3?4O(Gb@;e9a?\M,9,7A>\ZRI72a_OD3JUEOgJ7=+@-]
KA_-MPD-#O:Sd#<+=;gDHNGHf)d1b(Y9=YG]W9RGX,6J\88N>0P_WONdAT:7Y=]G
3FZR:KA8&;K)>67Y\MI&WZMW^C9:H=A&8L58R0U0a7<&;NHa0ISKB5&;&LEU.17+
TGQEHS\R5LT[a;Id5<FR.H^JB=:_(W8<aBSUe&4NBScT&I0JW/SG,KAQ#XKb61)\
#1IBa^30F902<I]^IJ/B25LU9Ze1&-G;53<25<OMECTVFB)_V0<G+Na89=F#C;_)
-f^N\V<1P<4BMK6X3b88&?f<(SVYB,A=5aQ8@48D)NM]GMDf#8J.N[:1,-F6]D-9
/SEYbK6,IRcKMMS9(bZOL<@Q1<)Z0Z<7U2,YX]\/Q_,3=5/XCWM-=7V3[HAB.Bg1
7aYR?/)\G3/?7]ZS]6W^fG4PIHc@^3SCSW[;1WVVIa>G)AK_<D0^cZd\.-V:XK)&
],\UM3SZ@^BZ[aSX-=fNY]0Y6BZ?Z>UDX0SbHG_O8e/DJ@0V^,#>R2?J\MO)[>E1
g9^IZ>5,HGNd,eS6aDQ[^VZ>T(S=<GFc=9TK/CU#A]b#O1Pd+NcB<0_H.HQ@gdRR
<ZVVbGKf4+QaMC>]8.60;4#Q-L+#NcFJ2I;]/Ca4V8-_HP/0T4DcFdDIB69a_?[F
NQ:LBS=[/SV/cNBS,b]#W-=90dcIf-4T?G_[gQJ;fAg<?(PcDbdV4\MgVb=)Z2R#
I;.1:)X:d9b9>gWV4PIMI?0MMDJWJ[D;030HXJ?JVNLZUcPGD>M5N7Kf23)[;XKN
J(-?X57876e78BZ2;E5TL(Q.;1Jc\)6Ab_bMC/2Nb)L.cL@R5e(P/;JIMGbIE4>0
EeP>N?4,RO(AQT^Q@&1:4g_+)g<ObA./b8HJ_33:8ePQ3:D<2.8f]GHW07#d>,,W
X9[7E[RTSR+KbW1;YZcS;>X^Y+(4WYPIT](GVYAV8?UF)G[WD1GW3dA<AGZM#5C2
Ab.BV[M)5Z1CJ]1DZ16ebF33&9De:A,<H+,e1,=(eg]3\>S=3Z)J8\W>U25+J4SP
R>.S1^JNA]^=Ka@?S6VQ,b0-=DVD_LWK?N@FNSU.7X/=C+B9^#TOEN<\fC\-+f-L
/;3J>X0^BY?aDe<M[K^=1KP@?R3A0)@Gg(c\D41T9N>H=J004^]@4P;bg^]6ZZ\0
c#,M&3E#S?),4G5\/8+1_^g;G^(Z_YZHUHU?fIP8F_f[97FT,6@/._?Y1^F>;U6U
HV>S)OF>(cWUX9O;X7eG-gD9;?#;c50;S\b4\aUaGQ92+GIf.FCLUc+3)dd<WEJ0
M[3@6e?&,aS<DANGVM]ZT7Tc=LE0W>M-9-=aPDOG5eDZ2R)&cB^?,<O9ZY;6G#FO
5Mb@TFH0A)_cYg@+/S>-,:/+faa.YbPT55[5Z/83RL@&cRec1cc(M.SDZ).<bNHE
eH0[U9<TL.K1V3)c&;.00EG_04g<^g3EN[Z<WF<a?eV?UZ8)(6MFD^A2B6fA#-B=
d1gGJ-O.^HV5<;efU0L)C>:9<8O^[AebHZE_fL0Z3+7FGY>F=^@]Xb7P?fO-SP)0
Zgd1><:IUg4?CX]2f]XMF5(bJ=MB[GLB-cVaR+7N0?aC(UG2eD5+#2TJIV;)]N)a
9U,YC0.N7US79&/fR9V3-6+RPI9;?2^eI_UJR4&X@(aXF0c7a7701SVU,^NU,98-
^.__B6U1M)32>H9@]>V&W8gHO1_Y/>_DgYRQ-fb]Db5U=F.+#D7Ob);aId:E.4[=
=?XceG7PS>ZP=]<,4UQ>fgeH^_af<9O;Xe&A>OO,H81BLJVFSWU-dcHZ+9(4Z4N_
<S3ME^XU=2KIEZL&aU3^aZ?9ASP+,BG>GW]\=AWW.+)Q[?+-(LgUP9Tg:YWXebJF
K@ac1([F=af:08>5e?[2U<JOJ/:)@SMH=)ZA+_Yc]cR,A+F_<gB@b6e\,)=ZBZ0P
.1OVWL0:-Xa<LcBcGUb[[NHgVGIbfU(P3O#HQX:=]-TM0(S:XF+dBU>K[[Z&:fPL
G-ISfI\>^c@40UYR^5.2Oc.H;c138U0(IO?>+5Y7IN8[5J@/daT6f[f)NN98RV#Z
fb/f[cVR\T4T1aLNda+B5@QFF:N5;cX5e.M29SbX;O6?2bOYZ7@4(ZL<6@2P/L+R
UYgDYK&I8MeG^bFb(JK?M)(LA&\AXG44-V8Q5:@7E[,[<L#QEY6]W]IJN<e=OWYF
11>I\I3&D)1;O[LdgLLPaW_@9_G&<0=Cb;N5<[B0,c)I8Q]),ZJC)Z-d[4:8]JKP
^YENW(3IJ@M#SC=fGcLU2#2L),aN/e&OC[+B&JG8W?0-P0V;:N)V9f.D4JSO-,dG
S:H)Y&);Wc_Q?6N=FB]33^8bV]b4,\ga_X1LI59fPE0IK>^c[3GHMLLRYX,9[QJ2
gQX);LX4HV8T))MaAM=W.B1_aQ(E/OEA3e?;NQO0dDW0B-W-6/eTdSbG&TQd27/-
G2LTSXWY1UF\dEO47L\YI3G,&#e)8_3A7Y8RL@ZaGSJ\-QWgREO0eIB[NAaMAS@X
HBTbTI+B.:-WWYY.C.d)BKgg6g2Y))6+MW3Og)_.[#BP(<[W<3N>+\H;F[XdLF(e
a@V3b,C9:=9H<&DLU?_[RH91\Z=Q<A3<#WO[\bM=G0G?/S\FF-P7aT83B],#e12e
)Q:9<d^OH,>3O89ZR0ab;I.<CL\:<Y.=/Z=6E2>>208?ffY]g/cOOWbNHcd94I?9
7dbJZ[>IT2(MUTT@7Z.9-+dP>J12N(>d&YUC^2b3[R.0H^_4X&&WA+3^>UZJ:=ZE
cZ]Y.LXV9Od8(<O45W;J7PVPaC\A@[CfI=/Q[2VKYFc/;Qf57T?&L31beV/.d(Ig
K#?8f>?)OfWC9-e\C:@Z0(,g0F[E#C=)Je[:[B7f]Pg&@XFSTQ#KE[bSQV?VE^I.
97SbUK5QGbQJU9:,@5N2d0#X>6MWKR3()T05.RgM0WbI@?^Nc@&L1LUe<-&,6-KY
fd]KDb\3RALfNAEbIF+H0fOYN0U<&J&F4f6,fK7\[TZH@VZ5cOM7AeUP+e57_(KW
b()),),]R3dLg_(\],HX3;6X9&;FD^G9S7EIN1Q+Y)<9<5c)GF6;[0?LZRMVWcP/
H-:QBfV(7M5PYN8K;^HJ/8X0d^-X@#c>]Qg>Oa=I4-)fS6SR-NgEg/75FYO9#B5P
FWb-A-WQJ1/2A5(8>;?#W0.>R#I<(ea(RUDG<P9(NBe)-([5<ZY6#eE?:2f.5G#E
K4R#6@+A=8NTQRRK?gL>)PJ2;c30EB/,B,<G2V?KaTGX7CH1I&M>LE\DW?KX&7KL
@IfR?BL1c(;BJT3S#H\H14N.)B/@J@->YR5,,XaQ&4+fWf(YSEVO2G+b:_P&[GI3
ULL2/>a2(-Mbg>+gGTL#<7C;.A@)cMeJYIYS@d_dN<1JTgfc)K:V.^5X]/eYLAC.
DY:FQ(6>=3[a8bB\S1LANN:X>gK<UF0VV?^Z(&6cTA157,JV#Y0UgXJb)Ea4]77;
+M,YM-OPfG#,,T8A#NcZ8PG2O1We+UZ[>7e8WZQ@/6M#N#UT>E0,/?K?++SUAC6I
9f@ICP&HUgT)<GeMN=M-/LZ:RUT55.._K7#>5cR&KM@(=(KKGe(.-R=7U6C=DBEH
IE^6.d^QTS8<W0WTSb+_VVKV3Cg7gKRGXC^a4P1GE9DB+82[ebfKG:J/MNBSSVg=
RddMKeEgMX9U.@V6DPFKF:G5R79N.&QgGaIRWDCDa+cFfBW/ddXT7de\(ecD73AR
&6I]H/)(ND=17<:GLMdaF_c8gVFK,QD[R5Q6^5\?V73<UM9B;-aQa];Ddg-]JRB-
-cd?/#EaOcBPCHOg]=CLf1+abgcac,B6SHC,QMZ7TH=\BRV(C[V0Z4PWF>fJMH>Z
PXDEdD@HbM+6ZSe4SS#-_Q9<?Dc([7?3&(Q5?I8-O=TP:eZ,W4U<S:+Ce]1g;Z+[
]7G_3e+eccF_]6+ZZCfG7CNW93Q^:?JUc.dPUF>9[fF<+,-D[,-AX,(4:F.EQOU]
EAZ:??c0Te5AdIeaSd=@>24.S0-PRW7bI^PfF8W001NM_<UF+9J[X?<+S)1J:Ce@
RE4+e[_-B8^342O9L)MeFSWU[1[^/N8ICHXR7HK03XVNQ+5/a0RE6G>C4(V:9XNf
a1O(U]b6[<Y<RSeT;KAURIP)GPS0fB60.,.UR,I)UaJdeO@EV>9HI7^&U2:7#G<_
A>9B6AS1)TZ\?5(1bX,/)X]IE<<7bQS1+IV@CEIe[Ub5K9\>HBDR\7D<3c7)#U(f
#b[Z9?&>O\F[L_1.f]JEV4dZc5WC&[7LBbBC/ZW^\06T@K;JD>N;=-=@8bE).VH4
LUgHT0<^&S1F2aSF0,9QZ9@K9W0dB1HG)<V:WHXPNZ)9L.#F\4G(@d.<4JOd&g[^
A-/8aALV,C_O7.[#AI0g@=.H?FGDg&e=4afX[_>I7/LAIJ&:()\32D/TDC7e.8F)
M,Yb)fC>CJ,BS[dgWL<(_AXYUJ,>Sa)&[[c9<IPD#_ZBb>.IODdRF>Ke/,32+e._
K,;LH1=:G(BPb>fF8ZTMJ/MK-^;AP>0gaX=UU&T-)eZ@J/ZCZ;4QPHUV;]&L?4>f
C+CfaRI[Va31eEd7^8:ZM[,4NC,+Gg:78MMA>.A_1NF-I3P&L<K&[SJN(d_=NFNQ
-D:OH\,EEe4f_E#7e.gVQ=\e2DUP:D[_B@AV#H0_ED8QTQ;;DM9Z_cMb&ND@V&D0
12N+RNOHL<XFMRfg3b0(b43c/E<3TRD7QUUaW(HNKF_N0+,-E88>].3X?-U6CIIM
R(7P[H4JD\UI1QN@=UR+744N3bA@PebZFWZ;d@L6=+bM\2CPE?41FIY:JfI-GYa+
-0@#MHcc,3Z+ddZO7>G\.e(FFRR_;RH]DT:K.BMLe-+;71d14G,L/7ECPd2VUO7A
;4&D4YDVW5-.W]4U@UC?7CXVGTMY=KF/fA94ZY?DH+.Md4O\51ffWJ2cUK4<F(U+
Z<49d8=CIgUG(b9DPN=9@1Y)19a7H:M&@PX&.dL?;\+E.,8@HAcVQ^LX03^+)G(7
XOJWRRT11?#.7#=f;AB.1R]fR)R=fJ4MA@^++M]c)f=:.QeS12./,05NbPG4;+P3
UYT>67I?I^^;Zg3:bE6_++_bZK,)8-ZZX7d+e3[[8#\:5LMC00:4[>[8]9MgI#=A
+G56;#),=T^F2GeKROfaVFbVM<;6?=gE3;JTMFa(U,]@3#W<=9d\d\PW1g&[)@H:
5e0-I_NTAY9@E5GOfS;E;TZK?_]8M=,F3M1T8A;5FFU(RDHbXQNRKJ>J9JU>C]^<
:W;0C(NJ;ca8K-Z41(=U:21NW<\[]]C7UJ\<;<=<1RUN6,b7FdaDB=<J>b.f9:;V
9:7I#WD4a_;3gaP&]dVc7U]d=3[=TQbVIXN1T8YDJLT#c#dFN?,Dd0^X54)e>d4Y
:D,910?S_8H16-2^[<D.UGgMZ8C[<W1&M^0@2OUK,g?10/b2UFQBAR7E;U-A/dPL
WcgTA)=5d,G:?/R+4:^cb+abPDY:(^/3M1eG[MeL0=\R/EENEL&WE<P7^F:RNC2K
b.<aJF<D.OJ&GM@NOCJPL^.TE6-4@U835gML;I#1D1V9+Qe-N--)LAcBFIU1;O-D
NCB#KJHZSM(3,8.7)@)g_#FV]-SXaI#ZaNE&XME2]MM-).2-6I_;,ZXI_6&VZ/\=
1N<4+KSTb/:XfP\cIT>[O)Cd5\&G-#HB<,029>?f/Q^acA71DH0[f?VbS;\a\FMT
R@[/5c>]5.([2N3-J4cNP@3-):+=Z_CX(#aDD^XE.DB37MHQd?gV9(:[>ZD_<W[)
:&+7V2_gBG:9I-A^H1U:+7UI1W5_6b\-+-4?+?EOW2S#M-_@S_3^W@>J1DC//.;e
YF.2K706]7fK]5L<dH)MIg5T(12M87Y#@Fg2?Xbc7=?/-^^4A8e4Dd#AA,aaC):4
QC@E;Z]K\)_Q+@C-OHc?,-\9@?]PS61X8bB80\e=/]G?1XIR9UF2-]YEU75CCDD8
=IRZMMLND@@+fU/SBQ</??42EHB<f.,3.1H937f]H89H6CF2L=D4d72\1=Wb3S@(
H:P3&aV)c3+S8+U(L_=&_#-S,[CKNgIFJ3PcC16<L5a1[(eA)V=]^_\#XBa6\0RZ
fEQA/ADOM0)>B=TUQ#G(41]?3/;NSgXVK^L_?a/f]VT];E@U+Y14+&a?=YYbY_U)
1#8IP;;C,.<L^=-GO35QPaK6Df93XN16dW8<+J?+55a[<:S:e.5U]M(:N65)<[bN
Z6FILd<R1E8G.=8LBEWNL>4&H:A.M9aF[F1FN^\-N<3K3&7=NP?g8UO(W1fg-8H2
.VH:+fBW\^e\[FNYD/\^M-Lb@9=O<gO<3^T.1V-[C&ZWfdYID)OV(#,>[?(GbMQg
8-#4WeV3U<JabICM3NdFW_+C/+,YTJ3Af#I/2GE6XE@VV63f6#-;/YA)Ge#9IgV^
XJ:3&#e_>-C1R&Z:VL-)&0XVd28KYM_YUTSF6(,_#K[U77B3Eb5ZRA#GHUI^\J,(
G\]bGX[CG)XC?>^-\d^M,>WSL#BG^<^Ie_R\SF#WeAZ536RJ]2@2=TWJ,_<G_<Zg
_CH-GBEC<^P123X^a:0,;TfYNPYGX@Q+GA()?20+Y&N/TE8PQbV4&2HW[A#_deKR
bG-I90Y0?/^7Z5(OePA7geZJPf5);?QY3,MPDTT=<e1Y:S_DQeVAE:V-@eI6U/(N
9H[_^Ff]fJ7U(G9V4/2NLOW0R:OUEQSA0&-E-&N&4SUWScPQZQ=,JR1TE39G5>9E
Vf^&\XOVNQAIXe-:HJ5EW@6e],,FZS>d:.4>;I<)dCZZ\OCS=H?[CcJF);YOH>+<
,4@ea?XN8Y-Z[WE=H>4-M##W@VM3R9>T#7??-U3W>e&?BfdL+GZ\F(LMf:0\S1PS
8c,1Lb9>#2]e/3cS-E0<=a.b0P]?DH[cec4]BY6][PbcLIRbL1\95U:Q^&10O]MC
LUf]c&M8V:_d0cY=YNd2+4@CH=?Z/P@7V^=;_D^/(&@22d-8a0gW)>\P)Hd8)3D1
Z36]<dO@aRH4.-dg6<>Lg?V[V]WHXKWZC8bS>4I<@^2V645.?8);QT@f@D:.5BQO
QMXN27T=LWUM+6OdKZ>&\Obf&?879PNP2RA7d]_CAAX-F3@8ZA53#6T3C&aIK.\B
F&R6.(Y^F/O3J-d3IJ-,Y;SYH^f)[>=XaE:cA>(4aLFa,ZU9LR,0egXgN/.c1#1b
T:@:_.V>DcbH&QUJ0\eJSWd\T#A_g_]dCLe9]RJZIeA<(H8GSZ2-dPR/fFVc1L/+
g]GKYM:[Q=]LF/cEBLf(8=M,5H=J/6L>.#^N#AG+HU;K:e:_B1L<\;N-HHZ)M8;:
=TXB=R2UDP5N=X\D7I0)DC&GU[#C[2MATJW]NFVdfF0/HC:&L_PAL4A4AF]P1OE-
4\YV^PLCL[0P+3MVC3IcNa;NK3[[(X.#4GU-<HIW)NQe&CEH9+dPaH][c<<1d]H6
(RU&(/=efMK?U]bcH0CAf4=T3ZTY[HEc>gA,\K?N)a0Ic29-]fA:\;.]<W-)B@#<
T-4SET?YZ^aM@?8Je+bB3)LbZZ2K8^QUZ6QN#)NP,HPAR)CY,M2<9OD1-1:QW>4)
[J/3C^0-82b>7J\+ZAC]:bXZZ[_Y>(:92->ZKQJTZ2^ZQ4S=QQe,U?FOcG][,H:-
RR]F6e;X&<O73C<SPa4/XCXBSSI:IXR4S(G79[#=J[X3JI->Gd8+O(FI@(((=15I
6:L.#)<Pc?\b8MSZBB_aNJ+:0K>R;UD4bO)>X]8WQEX[>R1XEGW;F9DC2D-P_CZc
<g\#26CdQ7_Q]:X:,__N&CAaF1Of(\/Qe9M)GPFG.N7Z(g>#@+O]/=.-]YN3G\HL
&EIOF9c8&2MW@9&KaJ7BLHEd8[:U\#EcC2DT1[GD6BC#V5_^GXb80:+[)0<)OfD#
0?2UTHH[6OGa[ML(0-2\))dF9;M4O9P4PLA7N:DaX1OM:?81fAB4?[fQG&BYC@&>
RC@,6c>Y:XX,c8(;=^J(62GM/bVS7?I:LV:([/@ERKf0fMARcF\F@SbZQ+d@0:W]
EPO-;PH8eGD5OYTKL?Fd[S#XVb&O5dB@=?19aYZ<cXLC=Nbf;PQ&#BG)D?G[SKIL
LB:9Ne_K;a<0geKXO0X.egH0S-)9^-)g=[@C@C17],>DLP-.I4PWBVJ:KDQ4e(0?
(UfFQX\+;QU0W^W-UHgDg7UafU\FQYgVcGf:;6-gO1FY5BSG:)Ig57DKBNDNV1)b
0B26TO=8+Z&EaFJb4Ka>V#fMc[fFQ=,,Za6@4QA;a8a]N)ZRM2gP:A=EV^GfA@NE
X<X<SYVVZ@LY3f5UXWQ.QZ&AFA^/:AZW=e:+?).KfU6R&,N7DGROU_^,P)KIG5AF
?a1Q^V(VcF(?<SRO2Q1X2FSDNAFLSdB/BM;6(L3HPN=?4JG=<]/;[)&>X;8\UK]^
V4YaQ=J7DUE2DO1MTEN:f=AR2@5eggQ;T[ebb-0Oe1+c2@H.1R--;RG-+/6cTRCU
;]-C:KW@c;Z)/YA+7;OPL5_ZCcT8D.\6O[JJHEG7:][XVAI_Z>P1=G3J_4<a5H;O
W6EDWIDeW?&HVgFELP291R8BgGPRN6/?QT6B+1[8#eU+OQMc6/C#:3XQeN&\-FX[
,UXO&_DEU?X98R.2SCK_1[.::.F_1MReJe1c2W83F<1Y6S(_3]8R\]_cC..VZGTS
\/>QMN:Yc_]dHaKR&@.:)__-AK&.@S?HFGH-Fc/YeJ<F.ggQBZdB]25,f_Rda#2>
BUSK#a15JVMJ[_<b]M]0fN-M#XOe+0NQU(b69#W)Ng/U[8[T3C<(D4.;b_57D;+M
<O=;dA7HF_PAS/#K<c5R&AJ,)Jb=\^aXCVDL_#YG97L#e0X2eBBc3(TGXA=C\eF,
[?VDSWJ--7g<&4F7^]gPS?\(UDQ9eV477ZB[fJ347FB4Ee.IOa>7WSJ79A?.0XMb
P&VH<b]:fYS&DTF\73B-<XIEPXb5<)58SLDA/&g^DL@K4g4HDa5)T0P.T_2P7B^c
K;H&FTC]:6A^3._X3_>?U7R?:-6I^gXUE^)dKI/?.>e[A92>RWWSEcQ#(DN51@U8
LH\;0YRN\:B.f0M2[&gUJB1.E.Y4c_K1e24/HSHKS>?>5AdBBg]&b3Y>0bA(g/aY
G-X.^N[B[6TD2L2Y<3G/ZZ=:,PE9cWbE/8([+3)X1#-W[W_aA.K9=P/P+H;1\&Rf
g+6<L0-2X/IQ+>=;[/V:EEW_#X03b_9JM-;?R:+6gLYgBL[C@2IA6.P@ES?1.#Y1
gaR()aL2b4X@Y\-^-Z?/YT#A>\;IW+Z]=/eU-10gM,<T/+SPg,bGJPP0&aRDgV:f
WT@_UR^2fZOL2N&e-PTH=AT2.8\L^3Ufa^e@T#eeXg+N[X@6+da<J)L+<JV]?g,G
Gf=;]Ug7Ed1Zb._&PSM][DJ81<XbD/e^b2dIAgIPDgZ/EeF>WU8D/#KH^DN&BJd9
?WW]L:(FU#G=T<eY)EO-cURZ@bYAPcgCE\JR;C1)?-.4WDfRfg&(MbFYJ7/X2#XR
F?E0f&Q:1KKA](YMH((.cRH;0OKV@6gKYM/E-OF@a3U.FE-]1)505H:?XIVfE7ZC
?/IO0(2Cc=:fUgOWFI+B]Pb@>JTeW]Y7=-0:J]KTfa(X]?EO1@SE9A^GSXZK=<0;
B<84@9;Q^cK2<:Q\F]3:b<1>3C33]]H_G<XUXc+1I(6?D=d:L,gdUWfX=.GHPeDS
0##.</HO+(@F[C>/@C&FHDZUH)#Y,_\6A8CDY#N]FXOf0dU^(O8KFZRS3fJD7?eM
E6&EdKR#Q8JIMX?_&Tg<5cSOGVe;NJ.DbM(O&b6L@F?;/FbQ@@4=#G9Y3G33XX18
?51]\1]CI()gY_IG&6)g&L@,OaQ<Ee9=3/DgS^3#A+FG5O&Qb8/]OB[D7LDeRK9K
](b44_8)S+,GL]FEO\1YKIZd73^MWURFGe)dZ[:QPgGd&;g2631Q\cU[XY3LefUL
T5:36630NR-[W0&]:<.=.fQ.HNUJU(3P^Gc)9.AD<\D&B34WF9d?_5V?(T4V:YYH
=7@a#+#)@;D;+KgAB&B<V>:,1JaYfTb#GB-LXP9Af.MLPMa37]I(->)BCbZ6/a,K
P3ZH8(+\gd#PJWe8b?Q#HWVQ/QA-F.MF=#9E\#&)QA0QROTLgfUbM?GaeAVZM>+X
11FA,8E4.QB=JT#Q9IM@f#VMaO6.XT7&STF_L<?<IV9015)KVBNV8b_F,b\)/LC8
T2,3EK15GYILXdNX9=SO7CZT]c6MO)-C+/K0V&ggJ([0HJ]PFJGa84=:dGSQgd[P
U^J&O[99TU<3U)(d&7Uf3e#VB-N#=+/VXG=4\AUF;]7]/O+F65bcdVb>BV3bVM\0S$
`endprotected

`protected
4FG\gK?HKL0;FJ.0f3J8(L.I3GH[I2L(:TaUNgX.Pab1fM)Q(P@_/)7-8ZBOP)eT
5#U0DVA55d9\9TR6M,AK8R.I6$
`endprotected

//vcs_lic_vip_protect
  `protected
dYF]P7_-B<JPJ)6?.0/=(2V=FS-)cQW81WIQ8=JO&)4.e4bSQ>U83(V)8a]0P6e^
EBDBf-Z(OTK];Q#&=LP7H3\Q::c93P-6)c90=(1A+fCW+_WI-CEL,aR4^;_AgF9K
EIE:JWX[_7D0L-[/MgdgKSZ7<KdJ,.[fF2MR:a.Rg64c].2.W#-&A<1A2:@KMb-N
FV-cWda)36CFeR&GU8D7Q)ddAb4XOTA0#[D,<C5Y74=Y.Tb;2UK/#/J=>X.-TBL,
XN-N>E=eSV/B6TK[\#J;a:2cEd5Ka1O.fHeVUX5dI#fD&F6bZ\)1.(#4HEKAFI00
K?G7:W(SeSAA?U.S>TW)FZHJMb]]5RB?3gB=K=)MKP,NLM7d=d_NXV,L_G6SVG_D
R]C#L_?J]2bWPK6>3FERW0U53IJFA>EYG>TBU^V-QFBA-S_.^A&Y9\QN3X>aEZF-
9H->=e4VgFOK^SDW;SPS.73_1I)ATgQEc9FJd7@E7&2=d,CM0].(,MW>,&4Ca(SI
7J9UaM]7R-@MeML^;SI4TWa)WcSQ:g.KPB(fC@6]E.VP5<1[[1D)8[R+\ff9e]aJ
A]b_LN0;_:DA^);<^>O;535?@)aLN0Hd5Q\_XLeY;]P@406Q9UF]=g^b^XIfV2+^
&(<]EUA4)E[N)(<;aQ4T&X@QOg?e)10c]:b\X7&?+K,QRO@(2J6._TU8gT];==IG
:WTT#bM=^YE-;(V@:a,HOY,g+,.>M,(dQgK]LMG19/2cU=U_?R;=TH)9G8#>-ZC?
(=4/0.LAL2>;^HD?PSfK4]Ic_FQT?E<2FNR0?c7J#P]gMR(@Wa4(KUeY72a,0FaK
:?ZgKd6SHB:4>0HO4fQ++E3Z3#W<?ST:JH\XP;b4N:2NF<V^_MODf&<?7WOg0RWa
59SEJMM#)<X^A1#1Z9gaEG9[>C.CAUS?W2f-6Ted(C,PS=0S4V5)8R;c;g@)EfY\
D@1XY-VR,7+[-0-IZ#LP4+:ECF-I].Xc7G-7F2HR+PHF.X&Cb^\S-_>_+fX6U[S]
R77JGYTTJW;D^-X[#?:SLIVegNg+\6\6<17=W8cD+Qe^Q7@[EQTCIa36QY#5Qc3^
)_?>5;1#e9ga@FX99S.ScWa.BZ]W6V1ZgD]4fTF^0a2b;S]C.bZ_U(-JNKR->6Rf
aXR1\APE:BHbO8.8g0M&L]3U^,+,Y&[D@A9;>4P5AbL2?S-e1YV=7I-8L2+\W6OV
>QRJN-8AGNK3E+8PIc#f44IDVBN&7eFZ=FaR:?ZC:U8=I6,FW_:_H96O?\S#7S9K
LOT>1e8K[P,0eH).LC^]C&Vg,U2KV&?)X\O7fT8Z1bT0aW,E.EHd#I#HW8^(aG1)
/SKY-@>#8.gN:P?N92Uc[6G#A8dUKQY2+<HYG3:\BK(<K;5-YCJ<e[FDUHK[07H.
RT.6CA_3_J?XGEV0GY64DKQFD1[W37+28I]TE5e2R-,67#b/D[JV1JZG-88<,G2<
ZY=IYE2g;0-4cE82@eG\7R<K@9EJ?+QY?0dO):OgZ(E;6#]eF5U.(R+@G?I=gcZ<
H[K]@-5TUdT<[RWfJ_5@V8X9AQ8a+=Wd<HOMb.5aeObA)PA49D><L0NSFgS1[[/9
/)4)BAG1YNgg?T_2P3Pgc+PLAA<cGDY[c=GF682fFB7+5N&),7ZHc3\&b1X,=0:8
=SKB#93=cL(C-99X72F=:ICC(a4O@;f7YgR#_71Ge8V&8.3gYC;&F]43;&3CWUZ=
3Z>.C]FEB[;5b6>NW2ZN7L2<B=ZKN8783GGAY&ceR6;MD0P?L=P/;JG8g\,CHE)V
M#FL(=TDdWINPHMCG\44=B/MOECX4X\B^F]O]b5AH#[?f6]M.K.NT_#WXMPWW:IR
FJ2K:F3e_.@\_QTWXcWGPd&1E2UDdN#XQ]FLSb7c[+g[aJ8UaXf#I7\DfU72dOXQ
:NBY&9aOHb621APIY,ZY/.WALPHCMc4:=^MBM;]YPTc.18_C];Y,TeB4#II==d?L
-b(fQ;9M&EM5YKRdf^VPd^I8_1<>R<<>MI^0((FR+/cbO&FTZAc44YBeNP//^.E1
#?BX+TP?HMMJV?TGLS/?[5N=@a6Sg@I<;d:Lc0LSOeA[gC7Y/.2M;J@Rf]^V(V],
NMT_5V^R05bG;=HeY@R8,?+?aLCM6B_]dHeSS/g1c&#R_)(]G<=G_YJ<U<(+ceZN
g:GJO^+fTgf)+Og5WeWVBIT\DCJ;a<N__4eJG(9X-N?EOV0\[E\N=+?,.g7TB;9[
2MeDLX\Y9Ta@9IMN7=P7]E:,<BN:9CL#<[[I/@ea(4M9(K;AC(9]4FfXK8CaZY\3
LK[LW,f01>X1bL)D^I4@;EU6=eHM@..[EHF?7:94(\>L_=R)\<.836<aJNdW9MB[
L6c2d4[:S6Y_ge)4LXBS9.Za3gIafBGcXG5[V<K(Q^BTYUNT4.C8KNOAIRaEeg2A
J[>K<@bX?3]?J(dE&3L(#DV>#W[973_W;$
`endprotected

//vcs_lic_vip_protect
  `protected
MXV<;@f?Q/F2aC=T&&=W6&H/BNB[OBdHdB\>[J+:T?J2IX<9_?3K)(=I[Y>]3H?=
_@gHJ1Bd_EC</([Z,=fE=FB.03#6MJZ1(L?AVPN8AMHLf7?Z8)6d[Q>AVM)\6B:N
X&K[_+cGK&(;Z,^]-LN1#N^_KSL2C]<.RZG7C79#?=c<>6&Z\,,0[#4bg&>:KK?B
bMNa7DT2?a?YS[?E;98-J)QOUd<;LW@a++18-S6.MD81=LSF#K:H84R=3SM_\T<)
(45PL1)F9c)N.Z?28QE#\WcaQF=+?FLb:5cae59TgJ0_KKSMK5=DGdVg:.GZ]IZ-
#,K4cD;/.dJFCKaOB1AYAc>cZ+JbEV+T_aPF-OScA/De?.)@?b>gDGeF#gf6_LKH
,,dNQWBCd_Jc9)b_###8VfE:^)<JfI>A1Yf?0F\FZb2&,/2dFAFb47[)_LQ3-HQM
d,9A0-YPcBH^<,FL_+7@.f9PaR2P-U6KFf96716]86XGK;1_/)P#<Sg>^KA_DbT_
e:>DRa:XV,F\]WaP5a\QMg)F(>XI]-)/V-RXb-/M>32D<<(@BM[dKBA,0U-bGUf0
bQL6Y3I&1WIF+U-@4<g;edB8MG4E7db<-a_UKVM#F_7:A@UQCEVbIcdX;6Re(OIN
g\Z[ZWV>+9P.d0Je7)EM>[e=gHR@#^\#^?+fJ^+e9N.4c8gY^;IDB#5;E_T&c_=5
R=Z;1+8U#ZKB;>HC)K8#V,/<A>O:5+>A</1WK27)[)58(OK01=-[bM&VF)_,SUPU
0]9B2O5\15.e>GBa[4JN#eTABad^@X]a7<(NA5E.W;a>#U.(gA2GO55=Ug#UORRf
?4+bM)JV:J>Ne.dX#1SQMI500:d>eJNN_\26W0a<Ve:GGObLVX=&VHS1g++V[2AN
01eL&9SdN-QR#9LQMD.aMQ+(67RCB>0eJB7:/@d06JI+\HKI^9bL9ON1CXae#5TR
/F/La4)1)XeY@-(&8d.&TCMRX6>4LB6MF@F4#9ILUZ3D\#36d]^<HU;]4@OeS.46
D9QLXQ9_gWeN7?CAZ@gNSdQS4&5#JF=fcN]Jg++6_^),B.9:\Y5R=#48V1H8H.C2
PD)1d^L7Q<JKS43g[9WX;>]:(g;f?fSNEDad_c84LI4&U+d]8&&c6YYZ([)OS,@_
E:<0FG5XT@QVKgDGQH/a[IU,.GXW=4/f>0[M8><@+T?4G:MBQ&ZPP/42S;bf86gd
AXYN6GM([JK\QWc<L[f_5ZLg+4,U(3caU@b_#(#J:b(Pg..C+eYD:5+TR/8)=.F0
dUc8?&UYM:8)X5GS>=TS[fIQ(XUfP>gRW@DfR9GfZLG\,?[J?9,OBPCcF+^^P6Z1
cPO@ADA67NcDONT&/29,V3YR^+3U97_O#0PdaDY/.#\[]6:\4OF@ESQ:0SNQ51=6
A,;K+Ob6aR75SSO[b>XT0.6GDb;_>E^Hb<DeD?LH?]=^gDTF)U/)E89K42-c^@3<
./Y:G91aT3#RG_Y78#,=<Q;L^=K+2dD,1?)MM1AdFT]D?0A(1/8)Df^/KB8,WfXb
Sa;7.I&]T10?B&8:5[9R&RU>[0<OfX.M9$
`endprotected

`protected
:F0,L&=73&WG_7;I,JR.7Eb4HP^.b[cAb;TW_04-HFI\N/<d&:IX,)=DN#_-Je;(
Z>,eOU(+7UE:aK1C+XO_GYb46$
`endprotected

//vcs_lic_vip_protect
  `protected
&aNS#](2<N>EE>2Q5DOCDF\ON^TTV(&(5Cb_RH_1VG>HfE#9F4Xa,(4ed3NMLM-A
Y2R:cH=)6G)[4DBNe4#-LS;P7N88#.0;UJf>)N,UcV0#Y4@Q[C:NbCc9KSC]NX2#
?8#3;;+G&H>9fAfPD;g_M[[;:4T4B[7R7XET7.VY9-:I[FI0,4bcZ+0^_=FHBUbI
7-HS1O?eC(YZ8bZ0U4R&NJ5AY@S^Q\#LC<F6@:G=013cAAd046Db;Y,+=Q@=Z/3^
[gLRS87C#8D\JN.Y]<IKY\4;b]C64fg^?U/UIcFU6QJ)a?TB1dH[,=a6-H3A.8PU
R&efBNAM<PZP^(C71S77#[@8:TAZafLA[^2)?HQ0&GUB+^?8g,(PB>ERCUK.8,\d
f8a60FWb)>[BFZbXHRESS(Eg2W^dc;H5_5ec6W.e5K33XIH.T##M&O6J&XA/g&b=
I[g(,^L]L)c?6,#5C:KVYfa?OR>X5f)f+d,^bLGK34>PV6e[=3aR?.RA/M82N3Ef
1dN2\Ab7Q\ZH=YCV.XR4?YaK:PGQOdR-99dUTMDG]X=/(YI&+J4aTS0TbLcRCZ[a
G3@U7_]XXa,@)BdR8O5N8C34_9XY.\10X<4&6bUP4KGJ_ZAD]&#SPX\?7,4b@[]1
a\W5aK#OJDK:I]]aA5XWGP0Q:,G?,CeIX&,VB?d/F>>g4;1H3)?DP;4X1K9WL;E6
gM&2.0;=URQdO.d=2S4I0B#_2-g,Ic5P,9beBaL)CY:Bf.PLW@8FIeb=;(]_[W/=
?J6UR?IZ/3N8L]D4ZW7^_+[RJ;DA_>USJS5dOJ2IMU;(OW>N9_WFD:Q7QYCOOdSY
24=W&XZ(e(:QMI.CD53<Xa,K9S;/=P5N=QP/UV@7J;O)aGM#1IO@()]:aJE6CJ?4
EPH]&5W1Wb?49.V?(SE[Z7DXA[Z0)KL6&ME16Q>S9d@X&J=-EUSQ1b1BIZ#_>+>d
fA1\JPRB@T4N+eV_34IH_6I<90ZdW7gIf7KB2eab[Y.?4eK]T_Tg?Fa/3)b7##SR
<G.QT.>WE@7@_KO^c-ZcN1[#[M9=+LZ5DOL)5C[9g@@GF(H12a4]&2:faP2\,A8^
gU4VN<?_M,E+2<eIMAMW7<]Q<H=E(&]5Z&g--cHT5^aHHd\Qa[BFS65ZWL22D<UJ
e<541[T6W\Zg?=,bYPS<BS+EIGYK]R&T1<+DQ?:g7D&A=P_A=K1gN?XVT1Na8Y]+
a?VUB8=S<F4eS?M)Xa=5?1b,+VZ<KYaBL5QJ/5&LT^+@Cf-,,I(8A&bGM]6LWdT>
b+;+QKRT[UGK/[OM/(_;3/5LIb&+(7g>#=SdF8VD?>\MMV@,7e_BN3Q7,7;N@Cb?
>OYfA;dUJCFS0UAT=_<<7>49a(EN7YgVEe2Z7@[g,#H/@L8g+FB:R-e#M(f.MOHL
YbXgR+<&V0OTaH-,\V8_D[9\Z;@a]6I6.IYcE\0,>R;f_=fe-XK)(cEKZ1A:7a-F
^_ZFJ.406D6B:;HE][gFL;(BT:7X_C5#=-g>)+9K@eNOD_@:U1J+I_Te[Ef)QN<=
@b#_6^R^X,(0(faaF>._U7F<RHY)EW#N-[&E?J-d.]GS,3##9C-4b2D.I75W_B(M
Q_SL(H[(HXO;J:7V7I7[&P7EPH(H<KU4^>FCLd39@?6d\0]SFDCH,B9=YT@BAHP[
:bbc\@4AXB@P7#K[ZcJ3^FUR)62-/V=9472H+)[BA^++AKKYYeC<LF9MHO6/;LeQ
<AGKe&RS#S5XcPVIM,:69c7IbL(QZ+A6Q;)-KL^&bLQ-_TJ^HP@)(WY3A+f4_J_c
W(3E17c[Bb56U4CYR-5eFCH)O.XCN+WabGOJ,EB6B/4OT2OJL]\FD@Cd7aTbLAM_
:<HV8+D.5KHQRIYFE+C9VcOe<3F7JVJS29>EH)N(?N6Kc>4D<dM:QSfVUHY]4#5F
K[PCLR<^ca1I5R5f,^>2RH?g=CcI5IQKHIc9=@)@S:_2Ig#6G01cR:A1]#&F[[MN
VIX?.Mg_\YJ-Ka[=9dCR[HWd109c?S4-1H1J9[PABb)?B3LQC^C4JA6(7=6K]AU.
J]EI@-8B33b>GKZJgcPI_XHNf8LZ])KR31FH@?T4^WI1_(V8dZ=II<27]&1-SP[a
;##5LcXV,14/W#Y_d_bd9b,^H8MU]:7QF-KO&c\]F2bBMCAC0YW60bJAR9/US6BQ
I1d[KBO(DYX&U+0.:^f,ZBfTT,DVQaJR82NG^2gN@NK_J9MU5IT<\V/A3g)Y)&2-
PaY/6I_/8OfSc)OM[2C/U,DXTbIbW5(GC6;K:8<ZS@_fNI8Q,;dGdaeN)]K:V4B]
OH.ga&eZfK.bW8J>[((c.LEaG,^:N42-I[C67,6a8J[R&2UT=;5L=1_P0<<)gcJ_
e3HZ5[5MBg3Z+A,.>[^T?+SJ8Y#aYWAT,]A7Z<9FPJ+Sc?3FU18@,?6TfS&6:Qf0
=6RG23a]0_:gX_89-?Ie0EP=M.K)&.O2V>@+W+e55+T/)_9#+EUPc].8.&NU_65Z
@81GJdK70N:;QbI_a\/AV9GX\:ZI/HdR@I1cPQQLN&U]2#ge_.@B#Ea@R6Ygf+KV
(KVTYAf1LF:25SE+<IWe=4XK/V/9eV59QB,S?JFN/(6DZa19MG,WF>+7VRb,S^>d
WfP0166N66?A3(TG29_(TaEW,d4VU<SBd)5;#&DXS-F9RV&@61a:/9?2Cb26U34#
VV[GS\&N^W2IOHcR<dLBe)#3(HeB[bBB:e]?##93/G(C740/4,9KOW?_O)gb<&RJ
Z[XR6^V+eJ^P@\#T_85WL#&]@ff5)\@>;&UIM5\(d@(Q?c-IM6>_RH)b>N.H]\(1
?BO+b((DFIBF73>+):\e0VZ+KEe[6^KHb-R:eGKTN_g5D[+^R/A<1\>d/J>[G#0\
GX[V#a5Mf[ZL^d[g-@A?fZaKG@JECY2W/>I.aJVR.HT>9eb/S;BYQ9@>)JS^2dX=
@QXVFd3#:^-/WKW8,VZ6HVEZEWe:\f;(D2J?JS?LD3EUe?(;CI.SJXI/Oa6ZL\J>
[TN@9B(^K)fYN:5JS@/dD^RMFUH85Y,57B[gR<VP3@1DLPc[Rg<YKF19JeIb(E+g
?31.;WbbX^A6XL,Vc)UBCA>,S7BI(WY313aI,858OMb1;/eG3bR.&7Z9,c_MV4,^
P1f[;8\Qf51;AIFDDS63(fYK.TK@[0>KFAVO<b0^dF4\UIN6[Md\1g<TH&a.]5Fg
=AQM@GTT]3d(#F6N(=LaV]E=AeV^;9QEU8.:=cZR=D#3<W+CCZ3)SCe)5^C]):eX
^caANS:g>K^\.#D&7a73LN,_T[8YSGNd78c1<)eVK;;cK>a#IFU=&6QJ[AXN+[R:
c,A8#HF\dI==7^aV_L,IW;K\J?2QL7Mf=):Q6J100e#(03DP4/^^0Ub[9bbH-LPC
[Z(?<-K=3B4eBD=::7]^KJ5Cd1Mg=K:-IYb]K^[1V+S23;JN@3#LMNcgUD/,b(4R
_PP=e6E@(P+M;EJfQXQ8)[@271VM[bT]YeC2Ob7>WQ<#5B,=@WOSFUadRNcBJGeB
999NKdPUF4I4Dc+^XAd5/(43g#U<^Tf&BA@X)U8[SV?NAB21#C_0)),C?>L&>2_X
eSLZF5/<b^HOHFS?9dLLZ@9]:L/a4>PVP,047Ffgab2N@Bc\5UAdJFe1b?PH(10Q
W-X2UeEG_,OG]fbAHO)SONXMFX8gO0\&,H5\-OLU=/]RVU&X#O,FFe(-ecS_=4^g
=C1PdN#5</X],Y]&VFF;:P&0agR>P4))P:2CNT>K0^HHH:):OWg5cH&4A2A^ebdH
2eG[<;=DI:>#MH:))gMWN[UVQXY>^+RI/8/\1NCO:ZWKZ:3V\3E[1#^ZYD5@_FdJ
Q>684?GLF#_dWRe.6b1L3WRDb(PPfB<5^8076&RAC-b(;0g]&FKQ?DATC;/]8d)#
-LK:S4?U4D,HUSX(^^C?9e3D])A:Q3Y1&<Y(Ga\#[P3]&@.JQS.?;:_3P:P8)YP]
-7/^4JOC4O<1-b.aeQ,71BD,#O9#VQY;a<2g1AK5TF?f#38#,4D8Y7g2/0CD];Z[
Mg/JC3E48>\SeD8:->9Z\N=]WcKc&LBJ0>1KE?#B\N2>3]Zd8D(2DQVXC)53_b[B
P308e@.I6<[BJ\;WN6J/P\A:(EB8e99M7DRLTG_[(Vc_?XBX]bd51H0,<FN=QX[F
7R@]UU+K6+30.\AQ1<VX3G:IA<gX^XBc]G;P2eGKD94YBWFQE#4;=NMfJD2]g)Z9
H,2Zeg+g@;E];>+R-+;.fE_C1_PVL)3FGWDfcKM\Wa]M1)9?VZDTGQR4Td]YA^Q^
,RTWOMIBBAM1//0R9,8ab4)AS)@IWFMABA1e<IgAK/7\GZ-eE_O/[N74X,+cLE6Q
:YO<aEY]K^a9-SaYf2C-geA,,(7-G:G/ZBZA[97SK&FT=?P1L-PS4W4Ze^GW66]]
?:N.D[VU]?ZPM5W#&5<&L7S2=<\,81e]R?5/SYL2.S_/OeYNSL9&UQeCZcc2#8<1
=:54IBDEW3Ug?)XWP6VZ:4G^<+;S.cU.[TK3@XAWADULKg4#]H.#6IB/^?;MM0fO
K9Y175K#G/L\F^1.&LDMd,[WOV886\_SD\3I)X8(9V.f76EU#d:7<GWc+5-CN\^=
)9SCTABI52C>TFLM:OFQ1]@)Ba0J:YD728;<ba:4/3]=^4D=B@0.^7HM=5U2TYOX
g\7;BYeOP-/2f+T^L5/C84eVT_dcD,.6S,C+?YU():TUc0KJ4S>0.QM+:AI<5+J(
(Kc02&@YF)HAC7Xf6,7[)R;[48H\E]Af=Q:OU05aS@IA,LM7QK4J21AIB]-<\#BD
PCJVJIWZEJ/PMQ3[c-7BF]+7.E+-:BN^eP(+]KVWRgbeSD>P/4YKVJc_a2:?B8AX
a9A[TA6_LSM53>=#^6<1(G16N+V_6.7Z8YaBVGBVb)dg8_;HaCa0(G/7AZC79@TY
7-Rb0e,+)_Q-N.g#e\Q^:R:377TZZ9Z6_P:O/M\XOg/Ad9;=J7=0bAQP<[REF_Ia
M,8(V2dSG(.O1;e0PB39?3JFB6Pe1?/N)&5]K(B](&MA>O;+]WU80aWE<SU3H58D
^e3M6Q083NR)W#TA.GUDVGGR)QI./LGOH7e.3#W8F_d;,NY,)\ES6YK)O1=]c/6W
==YB_a-4(/PbaJYb&Sb;?,dED)&Se/fEN1AFI&3E+RR^WH07,MaVZF\#R?DW^Eg3
XDXfTbdPcXd>g<T4UQedYZ?T+ad_MXA]aFD#,(;9e@#(Q>=OSR0gH?Y[;96</(W7
:B7O9;O?8Lad#1YR<)P>G:R8&:V5M=Qg?D(:M#bcSQB3>1?Z?F6H^@^0IIM233@I
_&+ZPKWb]@7Se?GML/e98A(T1b>Gc4UL-F?I6A;>]@^G\CRN13BYH[2(=:eM_=:D
.]=CY52O)Ge^+.FfS9bH:R@2NSFg9+>49[&C(;52SGf;][\^RQ3OK9LH^:0#d+#F
0H-L#QW^U.TS21cJGE8PH]Q&2RQ?bb8/S+0NWRRU@=fg9V@TZeE+@FSK)6065Yef
:,ZH<dWC]D5R^W_0aR^C/a#g[d:GJ.ZT)RS3e8b?H5A+>VG:cF:e__(6ab@K:KZ8
Z/=Z>0?I#>>IM\OEN3;+GI\V)Yf&0[V^OOdQ)bc422@6KSS?^#ePNEY1)aE4H/aP
:^&ce&-0/A_>692L=7eBgYc8,N28Me5aS/.b60(QgKeI<0\JQW5,B)f^O60W@Y[g
DIU.4CMKfCPE:Wegd=KNLZX\1FD3/MQcAC\bAX9/AT#HQ8aOLTeQ_SJX[JP9ELbK
b<)f-1;M&..-:XRdg&&L4&4;]fG8T,L@0DE7MQdXB6f1A.,>V?-gFH^3C_ZdRQFD
I9^adL#2P48M-<c]1>>97=-/AUSD.3;C7.[DXaKbd_e.)bHCFB?S5QRRc6,UFN@J
=&&_N&@CG5^C+U779YQRA)<3CV3a)7@Ba^#@BB-a_ZMI0Hg>@\)f(XM,<3@D)#\c
>==U=aZgJ@Y/=::RdDX32KWdX0/TaPWE+.=AZ&RQ5Z,b9#a1Z;Rb40-cN)NQ-<IL
Z;_T1?2cGe<5ZSS4&dd9@^]VY4K2SFgFNdJd(;HU)aTJZcN626ZH.T?.M9TNSN0O
g6Y._K32UBYF0?TBf6g0Ba+BT[:5EA&7f2JWO]G=N;Pe@(egQTeeR(/(8[H/TN/(
YUT.c2#2@Q:9]S@_LFR0H2M-I9@FLf#0X,?-K\I5IRF6U86cb((ZbV4b#/-)DNTO
;Q=.Q@BHB]EZSE#>MU@D((^eGSV5F?LQ9.;HCUg[8I6556YdRIe#60(2]<PZF;<g
[>dcMT.JF@V#)?9]d8?FU8^0dLb=(]DI=AfAWe,EEQfC8_Z0+e:_^GR+7,B[6g:?
4AaJ7-+ITc?O/-Ya2^gC3_>d(XWfc;CSBd<#c&.cOHg=&@32<RJW]eVE[QP5_cNV
0@:LGJZE7M-(2<#4,a3(5SL>CUD]g)-(CUR&9:KGT<bKb@&;TG=VM_;cUQ4?Gda\
R+b@E.A:V].J6@b,14]Ca0IYKX)d0e&N9>(4TO,=Ld_WaGTK\Z]:]A[.-gS4>9S3
SXS_0N5+D+0D^caZ5+]FCTXd7I04Z0e48/+ZC];5.)^PgRCD5S=1NMcaS1U&Y0eT
TIAJS),_c6Y;Id89d-V@HRYTV.FS-Z.bG;YF4+XeCQ6CNG:/.N6:L+2\J80GA?0_
,Y=cXT>-+#U:2Gf],@T@;X3N_-S6/8gJ13@aC?BC@f#C0[9Cc,9;^>+edN)N;O(@
GV+8b(\[H+=6BUg3D5)cAMf0F<5[]1EHL+gR(--GBT;/]RM+]O:NR[[]\+b?G7cT
LZQ8/559Wg1e3Y&^;X7<@gKF47V:+Y;ET&+,^Z\^KUC33EgGOg\G)OUa3)&(X/JS
Tb)?L0[MH\&_,.R\M>PID,302\=8QG2bR(FC#_43Z,UdN(&R=BC/Q+33;+V<W6g;
(#:QM&[(>A-OCN5P/]6XZ,I2Y0a_(AP7=:PW9LVV&0AaK+W>;S<fFW?@8\3E<<.d
8c^,4X7H:]OTR.;YGS?LHF1Db-=]H/KB:7R]\+Z)8IUcH5^^9ZC:Q#6&9=5K)QT5
6])LMbM?/3=3_fL5H+0)I(f?):QO&d#]ZR#_CWWHLOCUf-OM]3MXTK7MEYE2YaL@
X#66@TW^M\@W779c2R.?/,RFK)<U3O^?6e)I(VZ?67Ef2H\&]@#/2[>fHB<QP9R?
&XP[d9S/9E&EaIWUBgFT\?g7P4)I)Zg^^8;_J#4>J<VRa6D?#&Q:=ZZRW0=E,NGF
Z>JZV(bI=68#13aZ2#OS]CMRL]dd34&4+eA&C=8;6IM&cH4CVT;Tg;+eH<d,9[O-
O?+VQcbJFY)U@NOT\7f/+(D]g,W-e0^6NFDg7ac,Dg;a[RR+_D6K-\dCME37V<Z;
3M_?b,>.C.;XE9N,<,VddaC<Td4I4KY+3ICSL@+YUR2G>ZAI+SM9DUIH^Xef]4AI
7CP>?4[),5F#:V#<+RDc0&,NZ,U0<,PM3(\=Q<AC<5.W<b8V17>1WG#eP?S7dU^2
PH]B03-=N+gXUg)M=Y@KC?dC:U)bC+25D^=gKe.GSG4R1V5W;HPGJ5#:8McgfC22
7C7M8&F)?@GY.62V]Y6e6\2KACUF+,1bUR9cg7J#?4&E[>7K=+\eZ+&UTE?K5.OE
e:XNg6N2e4DU-8CVQ.YA5#Og2dQ+KO(I)[KcUg,Q;EcCK))>:X>(8I[P5T=R3A.]
DW;(Q<UHgL:KF2X\U8R?Q0bV:5H1@8=3T9Qc+1-+B,XRY=@L^f;1<_<#(,AA31B&
:f<?ZF-+CaVH0AGJ&W.dDE1X.a:]de8ePfQDYTPeKH2_YCSgRVUMUN;Vg)eEPH_V
8^_J&QUR-cIeJ_L?bQc+D03caBBJ@<XWG)P&_5)dNW-A?II1>WQc/OTA5[-O0U,U
Tb2.#4LH=QO4Ka5H=DgH#ECRRg8WL-I8)(-.a3-d_]+(=N3&O^LGFMBD4VD#N4U:
P)ULU;S7ZTR1B1d/=Fa=Fd0,<-8.7+dbQC+GU@G9Hd1dT=3D8J0/T9)H.gP\a<Ca
F<Z)?4U_<,HbZIR&DSN:-T.#,a@9[DE#EZFGF1P[UGFC\#e^GHD-GXaU>bBKLFD3
XN?7&FCdgbHc5T79_I5gJ&VW6.\1Za8SU,KZ+27a71TP15VY@GC:&^eP:3D@bYg>
=I&#U_87WL1^(WN7b[]&61OBUYDX4eGV?I\aa(>9T=+L#JDYU7M3CL2);46U(?7/
B248_Y9\T1JWb4FS/Sc3-3-?Ra\A\2I_V_PFIC8[@YE8=]R@3g&S,IWaU[@:^:dY
TYA0Bc6KbOQ7BM6#HMEE&?OS>GA)Y:-HRa]7+/YRa+6OGJ[=IZY#gO/_Q+5GXX>\
WFF].<:2A<@cA@+4^W]12FK27OB()]QHfY.)JPa@eG=?-8LbUW3e5KL.eGKR/&Pd
EKN3f+:#K3XN1U8g7bQ:OU>ZZ(&ba>M\08\/77B=.0,aI;I:@H+4H>?LW.Y&c_67
7_MZDY;:6VbX&:<(,c.2ET;Q9B3N1#)dO,DPPFFU8,BW)BZS2R:6NXUG2&)YT,HX
Q<X+LOW^?Y_2VJF/^_TZ(VCR@U/X^M\T_c50)-IM._Y9:/UDdI,cVRLd>R)1eC8H
^e9+3O\I,fZeGQ:-g=M:&Z/UV@7,]g=208ZJ<e-XR\/G)VP^&J(M+EW&DI;==[bW
-=,SQ71GP]/9cgTeWF.:UE5,1URNO\MH<2X2TAZ_)&a&EW1V:f5DNT/49XI#ODcR
PY\#D@6bKFZ5I[PK=-UOJRUP>/\;CWG<LLC>V,5.<L7J2_PTQ50QY1Ea0;)WNYFJ
/N]I:a9XcHU]K0e;@6+ca4-95:#70B)We.A&D_96(2?YT=I[gOH/LB2N0H=F0C+\
H7.=I\AZT..ZJ_GCCME,e]6aE10IW\[HaZ4\U(((aRXT)12^N6?8\4AR>gVQ+L\[
2X-(AF(5;8GcQCBE&C029N?F6\8QgNLgW8#\>eD@4K-MZOGO.]cR-]?METD\RgP)
)=JXU0[>f-;Gb0?5524//JQ?3bQ+?-YbN5PW[RMc(D2RU\T[ScPW,^V?-7)C&Fd6
g,Ze=1NNXb7a6;<WNK;P#\=)cf2BXD>f.8]G,Z>P[a^Y4cdMdEFU+(_MUSC\Y57^
@.:,MESM+1f:cZT,&57CgM;0\L>H]FVX@:::g]9ICR#J.LH1cg^HB)EL#>Od?Z<9
9UVMdUWbP\&AQX??aZ^HWY5YdFYBBJ1FcBg8a3=M9/=]/OV,D?__AOB.+2;[<+<a
=^:2NXOV+I;SGRS0c\f.T06,JHLI+3\ZUZeQ9(U/Q/<6BG^#f_173,RUHYD\9XEU
R_d0fN8/+46GSdV[GCg_UE7c40U;ba/?9-d).I//e._56GefA;fE4fUXLPeA7T\5
VA5bMI0Lb1F:I^NHMI8f^@G61;La8MA2@<2_XJeg->X5D$
`endprotected

`protected
]+Y.[O,()[P(cV[_D_:#JbO-MTTcUF5.XB@UAfeY7?_GOeP=C08U6)LTW>CeX5=L
^N;;]&&/QSILWBWPIc^]M\9HCFd8HV25;$
`endprotected

//vcs_lic_vip_protect
  `protected
9X?QTeS]?cP\#(_ZTY6c,DObV(/W>aM;WLbULJ0+?.R53bT(J9+^((b;=@RIS:./
@R)-A5dBA.@EaF09]+0Y-e7S#NKA+b9;WRHSK/F;.-[)8M>&S?1J&X)<<Pb0@69g
QEH\C;12(b]V&7d:R2<4aC]_UDC2#>7aQ(J\FTWKMN9eGG=-[+FR<<>:GXK@:K__
TW:32MMf/F#INCVXgYSb\1=#QJV^&f4=3deC5KG4KW&cC#^a-1/[c2_295cE<#g+
DX4Z,a1B?-?=G#_8/0/)P(<R3^]E=(DONL75@U:EgZ?J+dJL7P,95[?c-?6dbKC?
NH<>@HdD<4-UIL9Q.6P0C&81ZOH^WA8567F:gGYf<[DPE^?Z&9&U,]CXU[7>&S#@
caA9X=VRfcdNST\]M>]-;FFT[D71a0MAY_SI?^f7F7]H=(D2MLa1D;&L1e3FW&OX
^?Z4cT:;?7(#=1PVS/I:eD]1GAc,XLI;b_a5:PY6RO4F8Xd]>..B+Q?,#>Of;&7<
HOH1WC(Y4YU@VNKcD+)NZR)=MIVO&(+&(Y_/.W)e0T[G])M_]_=,_>0XZV53LVH<
6D_#C)[3Bd?&Q-<<>I&B?2CVY&a9KRE;?0^3]#E0b)N/b=1P.bdC30H&EO3FB[@1
GY1^@PEc>PQJf?JLWZ4#@Y;<>f.@2]_442fMI+A6YVM4F(.>05<@ZT]W@e?PF8L,
O>&GHCP4J_76P<2DV.HR?DcF,^YD?&GR5G)b<Fa[CM-]O#-WZNRK[U:+/>&XAb?Q
?220K7,,YK@gZ<B1HHS-E/J=JB9TL7Z7[dJdaeXYDXZU;PPI/XL]6M)1D<_<V0DR
Mg.@]ZKH8\3ZV;e/E^^XL<@UA@)7O\FI<QU[L/H=2fcZ^2O:=4;S,412[);-LcDf
SXZSKg1]M>.2PFHL+?/5(?2;eU:Gg(]ST/?Y^WCgSd;R;R(d:GE>d\B:I?D06WUd
c;=6,(c0aY-+ZW,AWXfV.J8f5WC3(9MRYgW>V[L=.,BMM+<[ecX+L5#23HRD@Jb7
6>a_U^KTDR@-_-Q++g6d^#;Q,L-L@(bC\NdPGPWbIS16L@O,UZ6bNedTO2+e?JB/
=G^4E6GObNR[5fc5(Y6cFBE=]NW&2O)95VC6XLK4=Y>gAeR9U@O&6aGd@]@ee8KQ
T/C>NXJIgA=ONUA.UK^/d7VQR=6.A3TB7P227(L6_1#O/DFMH<_)?3T)ea?KLFC?
_AG?&f0M>Y?6(NNQB,\_P74AI&5PS<0]EJf3Pb#CX@2)2L]cSdUeQ_L;@YP5+>EF
E#YR@&cZ:acC(T@4:^?Z414Z-TgA5C]BG2@>LeQ.R5ba,A0T3+];V<BSKe>G+g,5
)U.#K07R@(H)4AM(5OJAeb[:@A.0+PRY7P^.Ug0ce,<SW0F]cYL,HbaG\NF)O05]
VZcA2)7\PU;ZHG>c9,Of,_JMPc&AMJIGd>ZV;?X04;7U2eeAS6]L?dA@Nc2VegPW
RAJ.ZJY:QY]LO2F#010&NZ-EI_KN0.VE+UURN[Y0#gA3LP=QD>80[5b>STHA=<78
@5dR9>255V2a&OE3C5/AFUBQ?1/TZ0@5gY7e&_94gO/Y\4Qb(8OLf<V>4H/9FAV2
)E7QI3Y.K2bFMV&:C4,eL]Va)#g?O&,W,M(,<cU4A#04eSRd[=1ec55:[#):_THZ
I20(X;#53fX,.IA5f085X\2EIdfI04[V2V1eP5I\7L46gV=8g=J+:_U3:^TK)R]<
Y23C@COf[T_W)\+0X&&Q5;Ldaa7&?X1S?/2=(aUHGMGZgA]4&&gO3-L\RYa)_0P?
:J_0A3XM<H8FWUbG#4c2O0C(>-&(M[H&2XN7Xa/)E>9843-:NB9gbJ^HY\JQPaHC
c8]DKFaJNT(fXW5FfCfD=7;\Sa;SH5@FP]BO).?0H;55^a+6AYX.[1NYO(-@/EQ8
E7;>2/N9#:O<@-&O]2a82_gfJHQKee\aDag?bNgaC5_<gf:J3?ZbaQaE+7WUCPGg
If&fC::T3\736(A5JcQ8bW>CV+#7Z0\:e+UHa-ME,+_]d;MWG)RFJ=eZG;CV/QRf
f)fZGKOK)6Q_F.:B8YF7Y.WfQTNJ9/.aA3OY<ZbD@(9CQBb=V;H<UP/0QS7;0dW4
5c=KU210Gb=QK6#&7RfMaP8KIBQ(EO&N9YW_JZ/7>&ZbJ,?7)7)RbH(U\K=.RQDF
3M54;eTE#PQ5JK#5\?#a-^;=+Jf0XBH90LX1H;1KEcW6I,>?26X<b9E5aHe:eLga
)Da9B.H(Z)0\\0T,/)D&MJG8C1&GCDG+H[HL.OUK0af5eaOc;@[5II4J>D\]Q];a
XS1ZgS.06PK5J;,5c]3ac<gcTP+7YEf)?SYB._]0)<a5#c=,#&6LU11U+,ML&KY7
F51,2A<.LE9cbP0O.]e31<dUT,@XM.DG?B78f/(K/P4]Ad944FD0;+6,R_3&fJ>-
O(eVb.V#LLJ]=V36\b3UJ::ad<NQ5FCceOS/BcK:<Db;?QT=.\YUB;-J&:4,(3ab
+.Q>#DBOeFQ(OHQY8[66=RO^6/)]eZ7S7T(>DY2#=bH0)4I180#8YYJ,BY7SQ?]e
)Z6=(3S0DX^0d<#;[W=H3,^0G8[6LF_.dgZ<UP05CI)W>cJbS3f,CM2].BV&5@R(
5<)7NOP]_PT0eBIMI</;b\Q].XV+<E2>6DV/TfFM/<:U:J5#&,/:be7WF_MS/[A\
?A3LK#\\1GLNf:RE#ZF:S6KLe&__(;8(^\;)<#XAf(^fWfAE)DUY??UBDZ7Gg;2]
A/7-]>V_D]3V[Oc[X^_+dZed/bD;aFd;<>@9[XJ/U6\VTX^2W<@&JO6^4/4+5bS+
3HEPgc>W(YJe@3UPJcV&BPU<Rge?T0GLH7-YL5dEb=Q8/2-&@0Z[@C(;,5W>B-7]
,^1/0g3]/&bFWC:]>7295)SeKZ1[>cK@;:bJ/g0U)XV3UH0T2d3<4f?]2\=8FH@C
WeT5XY<+1cc/S#:H&767KO<\I0aR8_Q:g<2]EeIb:&>age:NG)e2>C_e@QTF1I\?
cEX]DGG-g&Q1Q\I?+P^>X4+Sf=Jc2A4ADW[9F09T1@\CF]>.\J=^Y/@C0H8?e2Y-
B>5/c<X2CY3eA08:-M;&;?0TF7)7W&U+PBf=QJf<K^1aO?L4E>DA@YfX2[R+0?#B
=U/4)NfPQcT3X?LU:7aTOX?>>Y)M9MCN=FAX;J(BHIH_?KY&DR[/@51V=TBUQd-E
W9)V[ZF-3IYV/fWGJMR=[GC5>A:d<gG5S@6C^0TC(fg4Y(?(QZ7A-H&F4fL0@Y\.
JEGWRVF[Q^T..RLGP@aNHURA7;QY3XOG?e+JXPY_0@@YObQXeO<?O6>NTIDD?.W4
HN?YOI<f5Xc,SN(1HI[[PWI^&ZBX]CY2<#&P\KNBZ:<Nd_JG5[#ZK13XC[COZK9g
cFH4a?&ZL-@MXcD(,>A>9<=7^.d=]2T2XBJ):fC4(#R1>PWdORS\aCHL5#.VV0Yc
2<E/[Tg)FIc2Ff8[XN3VP3&O_YQXIb(]HI7?L?CEH3</;+2Z(]dO7Qb]))S]TBM+
a,UU;4b78Jf0FCF)FP:K/M(G^[.c\\=>fKZ[@CWS9G]APP_NJ@O#.\.N@2\(MQM4
6&)^5N2KLWf:^7CH_6Q@I&TAEXJWF0P#S8T).FFEFQ918/c](UCBTd]VbQ6NY?1)
.&Cd3>R,C0bYX):+4#\J3\F\6fN@(0cM)FURKD;Q/bXf92]C1<?^C)R^\1\Oc6W8
3(-f2.3W[KPJ<W>FW0F(Ib&Iaf3L@a1B4WZf:6U7,([aOJcG+c1aSK-Y0Z>N=>Z.
KD<X(43>F\Z.S\X9,8F(>K_G[e1)Z:U2+e@,@,d=P4.b[^Hf(HI(#@T9ARcVIWW^
4Y7=)Z6>\<#H+W^H@:,&61EEFB=c:J7V@NTVB8@V3UUCO]ISc4dbGPeBbPI>BaXN
:=X:MfDCKPGZ@&_Ta,NT^L<Y5.TCGM4G=]4cX^R-]WgFdCZR;W<(1R>QKVV)g[fE
Z8RC^-8<C;#F2DOJ2/K-R:&HMb2D((CU&GBF,FaLQ.DVTCWefC7-RYfBS3@a/VWL
@SHN1_DOcUXMd8ACJ9LVfS?eLf#./V4[aDRf.5T3)1CCBcU_:?BMX/>=_P<KZe4U
7c_SD\&QD]Hb^aC+A/\<34MY3QGPc-dIW=J_2:Z=?)O0W7PZW>068S97F42I]aS?
bG#T,?C]NBS5_/Z;Y,UH=-cA0Z<@@ceL0=\V6)#1?DceBUF5[b&&L3Ac3I.g2#X2
=3_S?QYA,K5gW2[=]Zb?6MaU]+H6=[3?.X[fBS,cQ.9N-L(;=ab(3S@CV(WLa&O>
@)#dY/)TV6]4V6L^_AXHRZ22Db<BL&bO_@FcV@J+0WgA]/OZ35-eId8A(c3WEg;1
e6,,2fWEDK(#a)/7NKKPP62^b&Q2=I9FR=0&L^bVYZ:UV0DAf^c1de15L;(c;PN@
P]83N+5UcGF3/:).^9&MJ42.Xa@M;?)+6?#0T<>Y8D3@WA5a4T?BX.f-^[MFgHZ[
N1&Q7O.2?VYO-QVef+Q>9e_)AEF)de;<F//B>IQ#dEMgU_2-+=K>1YF6_KBQ]>VL
#OIJ4?=+?L<C;d-WYA=1Gf1D\/0cE0NaW2B9+&C8\[S]E^I6ABb\d8TG;74ga?QA
FS:M^RH6Z;I.WG_5EI)GH[N^NXKO@9,[1H6ad1Hcc?_:N[X0cd_38e8b2Qb.T4<9
OT[R/gWGK69Xf(?C72Ye_B(-#5H^2SYB4=0cg)9UC[KYW/-:5+WD_QNP>FL9=bMf
3cS^..>YWV/B)-P]YJSIb9GN\_W3Z.aM;P(g+Sdc-1VU8K4#:U8][3;20C.^L=N.
Q-ccc,,(2^=62gW4)4YI+(>(/BSC^5_&C?ea6=JMA3Sbbde;9GEA#3:>).,eY),N
<,91_&UTW_@[8+.GQ;7G0TB&>,Aca2b?AYK2YFEK?Q3Z8KI[)cT9fN&L0;E;_AU@
1N[Q#G0S?>GP-QD9.@2\45NWWZ1EILcSgc?MIGW]9-DJ85[g0/fO;>eQ>E;#<3b(
cY?e6>(W:C&N&7\(4Y8_[OQSV_TG-8Z2MG2e_=ZL:C-;7bS,;78;..ge.;7ga&Z/
b-JRWJZSMIN]FWI?gA[)NE]aC;I&egLT1@I,XK+d,<fd:Oa[8Jc8G(RREeLY[MX>
eA<N\4FH&c03B>A07DETUQ(VbdF.-H5W5(ODg9@:@9W9#LUeN1D_5R2,U_+3YDag
C:C=;ULH/W-LGMG^Ub#WQZa8fQ?S];#E3MU,^WaMFB3A#;Dd-R:Z)31U/[[VO75U
1+H/-+63>&3AR\^ZfCN:CA<cg6]A/5]/8a75EP8BfOZCc-MQVaU1@A/?TK58@R(>
4I&YGK5:7.XQK#,+5<gZ=;aDARVWR723SP[F+]=gLb@0fV?AZMCBT0)Q>Y,UPT_1
d>VRb2bU@3aCbH?IAeLL>(8-[R=\[S1Y#T&T5,Ta2[PE;UVV)_3[T-B.>#A?F9aQ
X[DFgHf-PI67fLD_EUUK(;/)DPU2I3?JVNd01dTXb:AUKX.ACU(TNV3?K#./S<T=
+IH(201\,SbJFD1,c,3SA241Q^_dd+86Z6E]B,0)O1_FS:8cW>3(=FF\:J;d+9F[
?<0G8ScQ3?AR9WI/,QLFba?9EJeJQZJQ3VWeWHMX_<8YT:Kg1fPWPT)WIa\@,<3S
#+KRLe=+[,(RG;K&^LPGSXO2:-Q,>fNGe.O)bH#O(#;GSCegJVTH<@B<_Ef8H<3Q
G]PC&2-:A,A#?b.7D?_8X@]Y?aC30?KGUZ(([eaA:PMZPTKWUZ,+.F.[b[Q3/@0c
CM=UP<?HFa\T6E:.&/8:)a=^XSeE/U/Y8]?;>1#+6@PF#f.)\<<-P?V.M..IcM#T
>#[1^NSTKFEMM1=EP[TZB0MZ6OG2FNR]=DZ^G?=5//\X5GN38>3G<2Pfec86_1G2
7:YW9ZeFYJ)bONCaLVS_ZFXE7#d1d-87eH1[E6a:SD4aVZPT<08YB1,.\MP;7V\_
23Q-8BF-@PXABO-1FE(@LcGF2WYO78OYX[:CaE)c4]P6[F@CU0.YB\X95;c6N/&3
<E.C41WF)&CRHSPI9#VMP^-_]?U.?8,Ce7MdY9/F(AVA3SSNLS9G>(85B8b\4.\d
:X.0M]7:Sg2J#RfRPL29O(J@?dZK6)K/1S&Ag:.Y=_OJRfCZ>WN;\?EgAL&7fI&T
H<[a6J+c&WRY-YdS(]65^[0D&Q&O<--FFa.P7TBMf3L+.SUEb.G5P_),L1R(QMMT
5H//[/7@LB_T^;Nf]B=36c:+RaVT6_Q8fL^NH5?8AFC\.8bdC^OdW6ePNL=J7gcA
HW0gJ2#+?M0;/B;bHUC>W/)<I7B.:]QVg.b;@\SM<9,<b8WY/PFZD,&Z^fDUe,8S
;cfCE.P:2+dcI:XUc\U)J1THT?A<5C2Y\D+^47&\UTX/+R.EF)I:)K0O,CU1KI^^
<T9T[F,=eBcCWa>K2g1J])J3))#ACc8U()9DEE?4MITL83c7KDe>7fd#./7>W:YU
66<Ad>8ESL:04F\W\KHJ6;\P85R@@8#M_dR&&.3UW@RUFB)cS@NYAWe^I]APG54B
?>+c=QBQWHU9;@2;>NcS1(gQ]@WPR8L<FRS8]=g9GBae[+QEHP.a<_aD1OL0++2F
O@^.NFb,=PSI38GC\SX<[cfD=9A\JB\^.35J>7&JcL(K\_?;OM2IVFZCOA\C?Vb\
Q_J>^)^beV)VRU)XP(EE@D7f=R#>&=W-><//WEB>__ZT7)ERef,P54Q7B@dg9^)(
(.a1:9+6e:e6.bdP.L<CW[:W-8a7.X0\^-@2W#][L(Y1J@#2O)d/)WEf]V(B?W^D
70VO):f+2b9\U493>BDPNc18QYC648f0E37]P0g60H80QJa.=:BQVd#,DW>6\?WJ
b1.NS.T77FNLMaKU/If3Pe@^?<+XeNFGYS(QS@H3f0b:f(QeGOCK99TcWf]@2c+d
&H<YU:[.MKd1/FQO=gB5\40<E)Hg1EObbGcNMQFZ9#I#S)?4f-ZE5:?0eF(4)FK.
dI+83fR^M2;JL6+C9:6cGQW#/:>PX#?N-PJ.@,DJ)5^H8-YYKFZgYa#U^,TO+:T(
6\gKHIJ3KAL57g,JPW.RPW;K:+@EGAgVROI,=O4W]7@M8=5dZOC;A=2(H(=#:;NF
8W@30H5P:_7F=RFN#g2UGFG<GS8;=(;Y_PPDXPPgZGL-O\5WL[__F.Q_#?1^ed&;
fC[YS#3QHD@3UIeH[PTg7MdW;I_=G3PE)I256cU2@(IT/70?gTR3@5XBbIeKN2b3
d?UW[\1J37/,@IReV@;8?[>-.5[KI[+JK643Z7Z;._M>]>64.CLKE#_N=5baT\>O
6;2\eM0d]<+FQX&Z0-AQK#)Ag-711#D313.#[&A<DQK6RZB>X^Yc\YbTE_^J3WHg
I=U@JbA##?5XZ8ZN<VUEC\P>/A62f7E3/>OZWX;_FN?,.SWLD>7BPLaIC-0(K?HF
=(E#33:Df.,&LA[a=J5Q1^.?7][)ZH<82L@N)XWU>g;<:>Vg/&SMA<fR95FTH+U1
Y&>OdG.L7Nb^FLTKU+&\+>_D[FbU[AK&Y&][]cU.3\9,OY=2RH[M-/HA#M#gf,NX
dS^4P4KY[7LXK4PD:f93SeX)dYgS4[eP;Mc89/\SZS1(CKd^e?1S,\bQ)e&bF-4A
VA#Z]APUX.IS1M4fd^>A[f27[=4RNLJQQUA\^]EWGbAY1&2Af3Hd,VSE,S_?D#UF
_LBLc87a6Y=A2=F5)+N\;XaaA3#OYR12P)>,#]UW\^Xb#6@O+G<=2-X-^g:CT.F1
3VL6;-\>7]6&@b@QU2WN+J_-:=BG[E9D91^Pc&S@>WW2=M9a+EcG_7a-BUP_;dPI
P-7UE?:4I([\AODWa4YM+?CHf+654_>6(EP&@M5\ggHUIJ-B_2-ZA=aZ5O</b@3c
M5eLc8aB.^/-#I<P6A]Yggd+7)dZ?F4IG]5A=:6K.<6M5++e&L14]JQNVE?K3eQ)
^9^[7UXRI;P+K:.f1gM&([N\.4IJ@]Ye_[<VKg/YE&A/<C>FPW]bL4VJK6e#+X+2
7T\W-4;M@;N<YJG],AeR_:M5+6ROb-c,&JO<\6N(B?fNTW\U9[(0EK/?#NWU&)T4
CA4N[P)#6J^1.60:>+;IVW5ebdI+S<]FY6=]-XMcYEITMCS25.M-/0^NUX0DWP;,
^#dHM^cU6PT1bF^46(\R9R;?2C[7AX2W6NTfX2ePaFccJX2XeOB&SZF4?+8ZEQf0
8P[aY<Oa4[2K,_2ObB)GfMJT2COR[/19:eNf?>afG?PQ&Za\OQV2eM(:eX8W8LH1
]9UQV[eI<MF8]9XL?/D[T:TPeL(EN;V#V0f=BN+2Wb/>;aWfa]_RbA0/IOM.GLQa
A7=/,Q61_HI]U^6?=H+dM(ad#-VGR]IB72^D//0,.IcV&,C+DNEJ0XcSV>NVSVS1
b+?GV>bKbJYILB[\+/?[d)//e.2T3+SIV#,JP<)ec&O/Y.@FI:eVK>7U=U@b&+;f
Y_&cP_#,^5?7Yd#G;:O5S[B-G7.2?Q>9.]S<>C[d_\?VOA4f#09CdZg(@2KgK.W+
T+?9LN2CV<A],C;O8d0R>SfYON61>MO&dQE-gEb\FM_F.AeGIJAM#AVTJZ9b@Vd+
;QAba9.Fb@/@&)Z;H=N,5.E1gM^Q^8FA1gOfP@@040;gV+/&J7=^0LO2]F2Be3#)
C]M-?RL4X5=^>8eg>VfgJ&P.UNI3,+^AeQ0BYD+aQ=<Uc]??\G\XK6S=H-)00C\V
89OR>bgK2RS;9TIJ(XT:dI\E[YQ-#MTET#f0.ZU=S-1//gE_=c^.,Kd/B;=<KUTG
B9c_978^)FbWEKVZZ+N(RSF^XWDP;7,;TMDU2@\AMXUd/=TfG(5++;4JAPKP^d4-
Kc\A5P[CV_Ma7b]Z0H@]BZO)-=g;f8=M4C=#.b(7SgG\N3XLf587@SA8=LFc)6.V
P1>,<,2-;_MSPBf-_M)g[>O,^[EgR8aBbQ0N3=)=V[>(P/T^+fKH0S?Y80I72H^V
E;#=>b_cQbCQ:^?f--=B.[RP[WS3Y<^A:,G;VHS8DG6ZY,/fgIL<CPfRH;8LIYT.
=;7\S28J:G=U7cg__=EW0V.:3L:gF=eZd)^\QN0HJO\0Q]AV[8^YM(2H]3;E#8CO
6_a]2CC1DOSE8KJ:.56F_]<,E^+6dYSE6N7&dPF(]bE)YO9AO3F\M/+@3X(_b.1f
De8)QK)d=)M+&3@5,B)B<Z_]ff=[GH8L7d6,L0+W&.T.O4LHLY:aBPQ=[Q>g9EV+
DMe/TLOI^3TM,OU7#RQbaG?M6)gTRII^S62E(c.YPLH[9+a4\Y1eLZ(T)aA02CJW
CO<dI[b<XX8c-DSVG@U8W9T.M(O_a>ZJ];QE>b=0XANJYFJ]Y+41e&X,f:U/6+8O
bfN)6&;MRS28IX#,02QU)0bKda);S-MZ3cZbd;W8d;,:a\]:-2FfOG<e_:7L(Xb:
@eU)+>WBg065ZV^XIS--C<9b=U7862YbBP-aYP3K?\7)dVb;EWREA_YAB#4\>V#L
OPbJQX97?0<dJ1=eQ^_gD-1;d8GQ]J7M28^ba;Wdf#;d:AP?JZ1=_aGb9EOII,g>
[<DG5@I84bSaA2=9=F\d+VZO_RX:.3+?Y-2V.8-]]AF2K0?&@9S#eTVCWcB,+ME7
;G^AeK.AFE<V7S+#d:Cc\Qe3Z/M,?^[6FM<81;MK3/U=T:=?ce7[B4K4SA79:.f8
2_T4(G?KS8+<L=Y?TS:P]:ZR[+MBgS:^4Oa).(ZBK@Q1JP]^;?:G@G^KND=bU#+:
<-3L<W</]<:\UX7GQ0/^=e1Lc\K^B45#LO+AHU0ZC.;)QUdBE)I0?@1b-EHMP]Ab
c(42A-\&6J1#28<b(eGQ?e4QI^gc/HI/6<S,Q)O/ATHZ.f32SS;W5?_22<<f:44F
OF;70:E>3)@JR,BN02<G@8(ZC0(ZSMF7a@VL<UNf7\@=L>LJL50:3Y8YaO5OFLZ^
]XKQc/d:7/HN]()U]I\))A><N_fNF)Y1E;)KY\;AdbK,(\Y:GRT:29/RE-56aU(?
0D(<gbb#(7X6M]ZKF(bN9E#8d&OH&UE.K5G32.5@>S4f^VN).M8#[#,NYT3FSFI#
Ob5=#)@X-JD\>?BBKJM)Af&d_O(BUEfOE&.+X[1E;9V_-SM@-7XcD8b:B@,MMa#U
=@C\a]W2JMd(,?,+IRDD_3:=JN3aaJD_bG2_OX7b<HG)=DM^KJ&;0YHS9JIM2728
C8@TFC^@^DXH]7&_6FX=L>Q-Qa\LZ+PXN:B&1V)?O/FbJLgBUI+?NOaUSK6#IUG&
+KU0/P;cg3)C3QH?Q<f38-4DMdN@TSd8bXMdJ?3W1QXgT/C2SX3^VCd>;Td.S1J2
^ST=@a[D[0Zd)RC:KGU.deZD4OST\GPd]IM[L<.TLQ)-W?JfJJ]2.,TWcL3&XG[W
([J=R]gQf:S6W\#dY&M9(KO)M=TbSGDN+F7;7N>#17R?eC?;TM^UWg2_,6?6[KYg
WaF-?4I]fSd([ERDX[=S47BV=N59D)D0BdgWcW<>T;&1M0P7Y9>>OVeU=<a46MP[
J,&?IaWgFO@GPG.]Pf0=D:Y.Pd]2^eQPY-E-N1>gPe1LR^K?/CLc0V?CBIL-[_3A
Q&8IA[A,WO-f0DZdKWBBH^+M()4,^HNfRPJc::P0M:e=7H/Q0S4?2:5M9-I\Y^3=
:\,SN6Q\.a0J_MQa;a@1E_)V[e;D3II@\MFTeJE)c(OSV<We6#Q&6?Nbd=)J]=V4
e\G#N3c+ED&=&8)Nc@Q+G2->V7#Odge+L(d8XXE#QZELR]@F=.(JLY@+.<8QbCfV
H1MdN8+(KTZ_7U<P;c.E_8>;.AV9IGT2IgBRGaJIR&cTM-cC\<Agg2Y2V29GZF#:
ZXE/6_I<929I1cJ7aKaVJB3K6UG>]X<H4;_;86Z/0;0F,8;fN4+DXI((Ec@5Y?DS
EO_2(W+c;6WHMEc.=H6DKQ?N\@>7CK1OXg\(#[=K6.XZR=81A\T&2FBW,A/=WG4=
NHM9;WGJN3PUZ.[Ra+^@E:\DZbZ]3WTU[&]2AE#HfXP0-TBJMQ5&@#A]@+818_N<
(<B1.8D\[/9?4=(YG-c2):2#JGbI7a8HR:(/<.Z_N]2f(+0M(4][@]Y2RKSgR)f3
a@07R+/G))1)CDB^-ddf_94<0WLaX+W/8R2b<&:6UaE4@0dI,=?:9f5N=<L1b+NR
.;OM2:0@29@\A0QHa^2;PVNa\YE8T&C59a2]@_;KM2(Y[e7ggOCZTUF@8.8>O19U
@V<g9+1Q?;Ac^]g@cP;M?ec[W?6?+\@=9D8>G2^.+0\eMbI^AB[5>,P&M#FNF9.?
;EP[a.9IMOO:?\Qg/5@PXP8K;5Cc&=J_+V6S#,6TBJ,AL]O9cM5&@1S&Z8CEO2;\
1bIR:7X,Gef<I>bF;aQWDCPM:e2agXCFY-W^4+E.,FEBNW=@WL2RM?[[0a0Pf([W
=aIU,RX_K).K_YaK-)c)EHaXG^;GHB\?Y?@2O]V3OOY/,#7>TQdN(@M0)N<f[C9+
.f)NMQ25UTd(;a]6X6TV6-N_VDMSW_Rdg&?C@f&GQP^]K(gVMcN=Gf:GLF_^S\=.
UR-eKf;MbB\6<T5;7dOW3gZ43RH[V37?WgSP;7)+P8@gGRZKU;SE7V1IIP&^^2:7
fN0/T?gQ+:6SI9c_G\<?^2+R._\#:24c</H&)Yf8V:6eT9>(2[.QBc<K.dIU-4f-
)0&#ELG5Z/5A.aU.V)AO2LaR/UQ]aUFY^4HaU\8K\6Z@9a=,B15>MfYJT41-/LJZ
R5U14=VR\OL#?AY85KBD8=KHX0bRX>3Q)9P4;].aXg9;Y)(^ULC^f&#L9]g2E+d<
,-]@5gNRR,11D>68_N7E//ZYBNP87b6M:?_7SA,ML&?/(E7EZ-8Rc,>9aNWUc]L5
518@6&\eI02LO9M1XA#3Z332<H:42c9M=BJ6;9J92X]>?AP0DQ.b+bL&7cMR+CGg
cD0\U(a94I:?E9/>Hg\eYI]d1Q0R^R-J>3SM=6=ZL5-;_?[I?<S@T?RUT1c0c)?4
fPa#:[#>5[L-G[:V(_BH0:[W^89JbP#D0FgFGJeKgI.02#_?^XfO<#CTf8^P#V]-
P-A-U>#&G&OX1CJ+cQNb4SS^b@;7V@ggU74;2M_Fc1&P^a\f3VD_eHQ9E^&XKP19
K0X??4G.CX<]bCN@_Db>DD9Q<Rd7_>-ae#1:Xg@f/c5]\gfc;M&;<fK(P661b:CY
USV\C)ZHLXRHTEH4L(1ISZ&a,N+LS^+:<QEN116CO9\Y]cM<@<F+eRac:ab\^;V\
N:,UgF;=?SX>eDc^ZS]:X=M&JJW\(B?&4B0U+UAVe7H0VJ1VZ>9TQP.^\HM\[30.
;gXA(8&>)70Q7U[L879_F37;Z^@),PJ]J95AHVW>S\O):@X-g8c&3D&1)0eAK;W9
eUWd:SNdHD)+N>/S2IV>J&LJgYg:VKNSQ7P:8a4+@^(GR0=K5=B8?86,0/HY.7^5
U<<fea8>D?gP^+:VZ1_:E1=bEPFV0V-K&1\IO4J0#eG17bG9HH]Ta-N,Y,Vc=T)B
\9Y.(ZKJ;9+\:.UK47WSg,45,^4;a(0=(B.c&W,TU[;RX=31YKQ#J<Y-I5#:_60,
P@eY4V6FBW/?Lgc8R2B6fF18<U+7Z?12R@+FA7^E_[;W8.MR@SFaK/^a]VIb);B#
O@+WTKZVc4A,3R_=)T)7K#]0geRO\UJ050NTZUD;5Hd(\PV&C?dYDA:;E1@5+(^U
M64[_+1:PVe1-d2\=6/7YF<[5(>;H-F>+LgZ;H1&<3@8-#@9VQM6gE@36ZS,@/Db
(6g6dYe>48U8:0K;;U8=eBN]UEU<VVY#dLLgS(OOMU]M0CeH=bGG(/7@R^:3eJ/N
62E1YcJ]D)+AD;#AKf@f(H8+JU?T+c6W+&_4ZeL7e:\Wf+d+L]JR-T1KRXeQf@/X
IF&91cJ1?Q5?5[A@.XXJY-V8^.^-9DP>./,6<WAD:>g4\/P0K@g.7402@@Zb_]3,
aCeI3cEDAa3CIeaLgDECSNGQJ(.-[X4c(TOW>40293V+4E+[6aDeE&S^,\3@@QQX
f>M<:(Fb@+Z2,PYG(MRH)RYd9#>?R-ZgbK1)7[9<=/T/F1SNI#0NC\Zf#33dfC=Y
_Gb7gYd5NBHa^^BQNK]:.1FgOSA38e5NVU>:?H,Wab07W8]H\c^Y785^^6SVSAUQ
W13BYd?>D78\JCCY5IKLZ4]IbU4[3(B\EL>^Q+-FPH<DYSbD5@FY\&c)+#9NaOb;
)a\?XeAIdV9,aU+,DagG=^cCY_L/fF0);KR#b7[&4JR/X;4_f(2X?4bV^Y3]-)DH
?/@G^L<1Q0a><20QH#0EeT?Q/PWd&;=9I)7MRH.TH.O/;d80,)?SB:CKcX)NW7-W
Q&Y#Z:JWfZD.M0&\T:/GLF2_B7RMNJW#e(4Z99U]MOaeU/T(LG^e-)OdMZfSA<L=
E=VMBA<DRCBCR_\U7ZD1.c_?afN3HR8g^B9^A<d\M@/A;Qa9Oe3_KZZ+gT;M^@<J
?++UOKX#;[7^/RPRH^@eT;7F1ED0BRJ05N>?>Pe3DXNW[.PZa>cVI9?=0PGUR=4b
AL0aC[R:F&WFIeCQ7-dI[7R0CT<=RY]0e/aXY5KP<@CN.41;?]7,c>^e+,Y.#38H
>PI?1agfBF7:]Wf\]0DEZ^eeSNUC[JT64[efG004MA4DUFDZ(^KY-KDC2ER;,Y9A
2FD2NR;D.Re66BH,gZbK29HFgZfT/PS;V9J19&T?9+FbbgO.d-RDSSH)]]TfU:Dg
aeg^dAN,AQ7(SK3:_bA9;bY>&_;BD6a]KD]+MZ(KK\-SeG;80=a-J1O=<ILAZ\;O
egb+S+0BJ0Z6Z@Q9-_&3bd-D]#W@T3SZ9)&:6MQ)dd/NfE.M])f6VAQQQc4OC?/.
;cNMHH.0&L,MCd4/FIQ^?:88D>SB)LRFf-f#eIe&4JBILVJ+OLf<<?<(IQ@M&,5K
U8cHHJ#@#LSCW?Y6Q/,,Zg6MaB?(.eM_N2/L7/\OVDGQL:>[d24)6^F0C@+bE;Y.
>dJ,-0AJe:)1c7+a1,1&6?\1+=GQYD#[Xf25^@R/aG^?[^QG-;;H#QT3>0fV(P\Y
8)BgS7-UUbPK5fKe@?J4=8]-e\TU:7ZbfHG;7b=a2Z2+Z<#d-4Q8SN2O+Z\gW>_@
(,NHP;/GbVf;U;e[59TR#EW)4LBVCHH@/T@0D,>-7(G4AE3/H_=4;e10a@^ZR0;X
?ac6^-Kb@0<Gg<=</PJ)E;._b8,aS9fLe.)gP>OHO&QL#-2aA81X1XXc&a67aF+3
b#3#(L^:D>QVTVG-=F#VRK\?)Ee&1K\4TVFJcgd(>a6>ed(.BD1Y2O6gZ<]F-VcS
&J<.T3:G-(_\edFX[/A;D>,568g^LfT3(LDLWYZdU3+gSC_Q]W?VH+9-a+/Y0.S9
a>=AU+,SCa)+Q+U_[J9f)F3R8_e;T9\#Lea#K2C/I@9D^(TC\1106P1AdL&e=Z[F
G613c@(,LR>.A,370b#4KLPbVc(8]He&g3N;M>&SA4T27J(^,/M?c/3f,0+[=ZHX
A8>_-6^L<P[KPe=62Q<@>@?LBYJ_Kd2:T>=F#O@=@cXUW417IP^J-)7H9WaR;4M1
a^K,e5(_DEfT8^TGd4d.BJ9?@HJTQ&63]L)/T]6R3:eG^:RY&B4,P65.=M:\\fb(
6VLf)2PDQMAU&P0JNSf<VCa;4-/V+X/@U9S)O1DLDQ3c>VO+J8X.,=8?-PECQ4=,
eb3PH@((?V6Gc<C(]g4:Lb0.[4&9G,_):;WS1^L,-83]::TL5Y1QQf&X2O.6bC)=
#UMU#1CIDLXG@1V9J#1dU.Ff&PZQPO]<TW^:Q/A@U30H2X+Q/V[+<@#c<WfWFPbg
@4Y7Gde,?MUH/N-FE(_J):N]fUORbQ;\VVR1G2.J.O\(FeX)S+HSN:cZC]0XP&/b
HW@5c&G[=_28I(7dND]HMe+F][.&.Nf+(R4V2#O)JO36;#QE=d?V=_78;X:fGV6H
=O9Sfg33UU8(8:_8H#)/O4>Y(-]a:JZgdH1/AJ)TW>VWX,3LG+:J&4.N(W4+/?:Q
P69[RPDIF2#[Q(K+7(W=L+/gZ?HYURCIX]+8]+PVX:AR:a31:PLHF01ZY/-Z>EY;
38Z,R0YT:f<Me([1Va]PM8Q^[Q5MD8cMQFD]H5Q_O/\&VX.fF1L9cR9QUL=\0Ag5
C0@Od32YFfQSZ.a9XUSAW<8-Y0ICIeZD[]B@Ne8dQE=R>(fI>+)FZ^;FC2Wc[7L:
R4C]3)fM1Z#3,TK:9a50YGP=5ga219CAAL)fOfdT.1)VND?N@3\H;O&8>Eg(Nb>V
_S@#Xg&I8_Pb1-,?J1#LAN>:XRD=5_e5?0,RYfO&XJA)8b9II?f+RFe3T.L)1DZS
=]+,L.\;<]610=WO:XO-/Y:=V=4XbQGQG103SId?^D9T.6=(K4N@K+>@5&B+R[ZK
=;ZM?G>B:f9:48US8M&f.^V+c?D^7^I^?SZY,9\JgcJT<U[PLL,)EE5SK^bSBROF
1ZcgVbRPEIE]6EJ^H?_O)aQB<()];2R\fAT;S6OUNIMY0R20EPce;5-FOM5C.ZeU
O;1)M)G.]9:;ND7-JN:^.[>:JBCg9?J4M8KBC6/RR[H\5^158MWDVND]I-64V5^H
]\<DVafcK\C.dS_3@JCFA7R7X/WR,e(K(=E)S+\fEHaPCTgHVV^1/K&LB_XbbCd<
80G=LO]KN<249(M29X<If+\g_J0a+))#(_Af]@/^NOT^GGCZaM26@C>]QS+QAY8V
#XS6>Y51Z\B/^Z7]A_d;V8=g:@BKJ0^8Tg+^NceedcF+GS+Q43+9M>c9TN:TQa#,
-P)7>dW-\7SM+S0TKAQY)>BW-BN5FVB8X1bIJ<X&d(<0I:dcH665MY[@5f]a)EDO
KcVP05_4K]&6)Y/_(WE<?\LRGPe3MFZE>e]7VQ?I/eLV(fYLd4]WOMX,>-=JJP[7
1b+]^SaJ=&4IdN9S8e-/RKVAID5L4A#UTd>NMG=,:<:3[QE9>=PJL<5QB@_DCV0?
QKNR;N6/]&9]d4>.N?>@JeN[Q1E#7/ePN^]-NC(],C(8UCT]N:I:P0/g@T_PO9O>
4APFR4I.E]c5gOVAK6#EDO11S0I?bUV0b7ceLU((IOe-)1_+6SMM&aTS>.d=63=:
1OJU=#LM9-gUbCIUX+PDOd;0EgcZ9ZZ?J/:L/[&0/PQJ3EJ5>YTe,]e6I\fKQV/B
:@M^&f=S:1W9L7Fd&P)T,G:BE)_(K?HA[>0T+gPfJ]3<]C6&&1(C0BU86P0gK7^\
ZAWKA_\eCS3g:YV/eddPc0d\;McG6Y+fDL1bdg+S=]I>9+?0+?XA(U#KJ3/^)c)E
O->Q,.A;?]&GXRK+DEMA?:[9:KZM\]E_eS&IE@P1G8QBND@=+(&R_;F4b>1@_e<M
=.O^f6I1Zf)#cT>\J+JOA9O-VSe8Ged?]g24SN,aD;,OaBMF]=.#S/TfDLGR<Uf5
^)/-2RT/Fa_FL7N,G&@[e+LT+aU-AQeYI:_3HK3gY)[R/1V43.VTGbPWC+5IXQ_T
88+RFO/9P&fF;TH.-f+5H@&a73S1SPQd(T^]@_>RSIXSQSa32>&f=(#IY/e<&M7g
3ffGA7F+[bR>Z-7aPN>&\>00VH=8MBZ2e>CHI&da;f>DPGPG(NV&:\Gf6VfZ3fg;
A\d:+:\[MA/N6&[RA-d76VVP6(+R\_<B3QU1bZ(+8LdGNOGL7:/N5S&KS],Uf_S/
.+]gc]7D=OQ8WfJ9H.0LfXH\KU7+L(0JGPaJ[Q@9:OQ08TTJ)gb3)(C9V[_1@B0,
>4-?>WM9=)@66Q).?S6e?]D:LNO,2N1_R@_S&D[)K@H/7)6M;e)ZA\>^c:)3FdAP
_R5DGHSf&5:0?JI@3ZQB_1.Q>/JP5-)H-.PVE?#Bdd8@4CV?>3#]<&P6;H0a[5B8
@A=#17P;/HR+13L]U-CNCeRXQ0VZGSJUgGPYO86K8E>9I;FePPcIY1g+?=,7K5?[
gH>F&M:gTX,bX?\XSbO)E],aGK6<OK^G8W]1,#LP>a9Abde;[6<\(L+V&7EAQA=>
ObcCLSg;(R>B>?Ba5=^8-<(ORG@.(JfHZUX3NQ3^J#:1;)c=4LCf.J0T)cd,?N08
P?)&c&MZXE:,P_Uf4,I;IUO495(K<_9^(F#bb<[I3MQ,fBe_F>K<eT1XITgZgPJV
Z]G9eCXHM@eN>bTN:4XNQ&.LX,NZ\aU4\<DUN^b#+MHQ&AN:Q43&.7TSK3Ob\>:M
ge&4]]H];..[L/[#Z[#&VMU,LS4LVWDL60#?ZAQ1.#&,FP5^^FQTTV2f-NdO+Bd;
Y?feZDC]2]#YESJQ:-R5[N;R.?#YH1DM;&X4AHK1cD0GRf5(9+/g#JEH<M1@Q+WE
RX47\;]#TeA6-+N\G0_b#ZK=+X4_03Cb;c7V(++5@0Q?[VP287P,Ma0K<8+Y7V^O
T;a(\3GAcNQU?HOBC;JCGUER+NL5gc)Y>M^-JIGXQX8G+#C^;4)<6aEU/F[&S508
G-ZLRSgZgQ>D)=?3N-@_Mf147JJg,0+f/4WB^FRH6&V.,4A3eM<QWW):Nc;(Y0]I
TD<&M]:dP-@TeRV7PD)Z_/:-TW>gQ;0;>4Q+IPZ08M>3#7,3JD-I27E>MK.,c>CG
7]fX5eJ80NTN)8^X7F\HO#J(P?-/C5Q2R.;DU#Z+0U?C51c^fMG?4;KV2BCY/Q[V
Xa(F)B-#+EA_5&TQ4[f[U74PR.V?SJ4KQ3aR5_6VG+/MME<YL06I\CYd4_Y2B^Yc
(IJ/)8OIL<?/#,\(\IX3dYgNXSI&84/6]fMVP5?+W_QJY.AJ/-1\I#DMd<#,MPRY
35b\P^&G>4,VK1EZcT8?b&=NLA#Cg5ED,:?NQKW3b\7FaJ@BE,MDF[3gVfeFXP@[
OY=K[6MUUSd_Y(48KVa&O^2e_#S]f/P\A3EH.I#^:bU\(PXg0[Y-cI:F3a<HH,<e
d&:cP?AAH#3ONX6W(eQ-Wc2:5BZ]a&P3E7N(,Xb2PL(RK[f.;76H<Zg:aT+;G16@
=2SN:J&(9_^B96\;NY?=Z7IOE<HYM;UL.C7A_:T((C3.URI>6YK@#G7<U38_NIK[
:R?]IEccW_^ZNU<?:4M1SL7b;9e;I:F;c2,a6Y:986OWa&bBSQ1_LVWPK[Qf/]<C
V8+Z#@7EO?QRX92OO&O2P0:W#ef_3TH3^e:9X2JZG>CIGS=4AV1]_M@,d_K:3JA0
eMXDS1f+=QH:1T7@N-I2f\gA<=<dB^8[\MG5[FRC#R<,a-#aZ&<EHbA]H]4CEaMF
ZQNRFG+/O.#R0,#VbdJ#bP5aYaTHIf&T^>Y+a2SNYGa^]3?>)MJ^.G=->K\C7+?D
Y-0/U<1[e]UG,R0-P;g:(_7\a&^UW)DVWP)ESIH;Q9HXUVfSG&L??:0JNNLPOH<.
=+B:fJ[d&=+RV+<@=_T4V8/.Xa#7?W:#&>e+Q>7KSbN)66;UZdJNag>9K#I=1C2(
CPH@Y-edPQ_gc0YD]GK]C(/K#)T;F@9UIJ3NVTAGGC<HCFC)g-2Y[BBW,+F.Y;27
87:W\/BJO(b6fWF(:e9P+P92ce8UP<+#>&ZV5)D/V,XW_4_5Sc^CO2J;bbT1(^;(
)-e9W_5U+U2)0/EO4]7ZW<VE,VD&c1CF@3UJ,6CH9X.c(&c<XCea.67H7]cb=WfY
RMF.g#2E9LQ4EPf.aE?RRB?+5/AM57UE5-9_UMJ#MX=W8B(<N-;9K-G4SR0(Q[X<
N?QC]Pf19U<0JUW:QaC3:R6+9^Qda77d^?Kb20a(K4OTQ]L\SaB73RcIc4EXZ[.b
Y2fR8N[M@eQJLa>KZO3e+0D[F10a>BD#2Ed^;0(Z1g]MQJ,;-F?.^H+=Xagbb(#(
0HGgFJ=I\3J\>?J8E@M9:FVAF3^^bZX/Y(b^b?YBY>37/AUe0<ZT+cc:dRRZPG#^
Sg]\K+(97-J;O81DR8=BgU6X=U2B1NX&YTZJ3;02PCQQ5]DE;aR?GDODddTJ_Ebb
6cMeLCBOb2S-[XS7><YSOZ<_JH+]3@&,0:SQ>PB):9U?/BR_FR[8P5#S#)fBFIbO
79MYP#WF-#_YIec<7dFRTN:I8g2[-?ETYLAF+#_1]cF2c4KDXL^DMC(M;67+WbJT
HcW7YZ\8JH86B\(JU#Fd6A9@X<X;P5/]X#+QCOK0CXQGRA@=c,GT1\O#RfR7SW3D
^Xba(&F,U7F0\--ReT;PO9.1ON9NK>f^2+S0U9K?^VHMDNTAMJHT^.+4_N74V4bO
MDA@ZP5=VJ:<9C^D[Oa^9F]C68;Ff_P=<.T;YNU-K:M0c&?A&g1=FSOL&6/7-PT@
-,QP0X;PFTX^WDN((+TbcE/8\8/N=FE^?/\KZ&H33V<V:c#2(S)DZ&Y_/.-WR::V
38C:\)O\]V9EM&RbWXa+(fMAReE+#_)H1463:H_5L?(T:IUIOE2H.g_[XIX]VXH:
1ZJ-R2P2De.cB3(WfCSH/dG1CH_.[?Lf5eK=MP6#L>BbLc8RQ8/_d1JUO>..4ZP@
-Y@C[552Yf.C45:2.Q[CRAF\6F8O::=]dW8R/^YbO-R^+Pd0<)/\W#?2dOY0fHRW
]JN)5)-9?ee-4?(c^^^HUM8:bbf,09TDT:Zc6bg&U/]2&U4c4I?1_MQ(LDMI#dSW
>c&#JV/B4,SN8)I,Tb32LBG>RdDAM+GE2C1YbKYL8eJ,+3]ITOVHHC09Y2Yd>aT1
60/EUN-b>9/-(_ZY=\OS:@Z>.MaSQ4f<&Qa,gb=12UQ0@69#V79f]]QX\BRcg1\]
f9X?8-I.aC(MJ+2GMdU(&LF/N=REfP(P:9ER<Xd<V1/P\QJ@@A_.8D+6XY,=aD#D
HB,UU-SPeV7;Y\e0B;Ug/Cgc,T#65LY(fgbV_G62_.K;DNU_4&E5e]OD^OY5M:[Q
-39LZCK<X\?_DD7Kc&<Xf:a\JA+_)VNa>LfQ<YZ=2X9/D9F@JN-NO2&;RY7CB[PZ
dX>Y^_,_C2[F_59FA=\\+?(a/@bPG2(3gJI5P3XY9d[:H:AKabWg8));,Y/UNR3V
ZQKB^CYc1B]D9Re]d1N^P,;],;QF8H9E=[,e(GL(>VU(4eHH?D56/SO6b@YDEb\^
Je?R@.WEFCEFYT?N@D5UTQ^G2=?7c[F^0O\DHW(I3IAITc90]bV+VgZ;^D#@bfH2
YB7D.>&Q?C49bR(;KYD.E3&F0BP/^=gYc/G7Y\(Q5P35YVDM3g/+70B6-MX](<c,
eB4#bE0(S1#UNBc0Z(LO0QVWfII_7cSKP[YPVKeYGYA8Ye&H?IF5HVHZXCY)bLCP
Lb>[5G?7-)A\]N59,@9T?K@GeJX#+eXS0eB^4E0QVeb#a/;cC,9.V07F=<2[>=8U
_M7DO@&8C.a_D\?9f_(gW0,LS6QZCVQRYBCPb)UWYRYCJJJRPe.Q4W03684[4FUV
2c.6bTPG9;G=(1.Hc?bG,gH;cF8:&)S<SceOO1f)?DMdFVG8+)76)Z;4^Nf78I^X
,e)f0+3@P8N]MVZA5Z<9FM5[JJ2HQ;BUM3RHGS(J7+=f?<\/TA-<fKd;^+(Id^[T
+ZEXPQC=M3eI1fdG3EZJeP/[.R.FXB8;\6=N]\[+2/-(e=51gS/ZBg9A^0QgNDA1
2@d#(MN^Y<>a]BWCO#22Kc;04+@X0]>.g/CEX31W+LOg.]+MOcALL]>+SYXa#RHT
JcYTMZ(IeZC:7DBd.F4Eac#5d[aGVg4Bf.N.(OD>QE<]#TR0T;O)VR^a^=>Q9)=6
DbbRE4G6M<::.a@]G4=4T/7f;\ECO;O^Xc?/2W(U,5QLXAb0FTNdAC[FBgY,IT\[
)?:e#KWLK<7]<7=W20&YTa2;.4g.aA5E#<OG^VRaA)aQd\^/IPTP84D@Zd5[2b80
L8,?dTZTGX\[UZ2?L>]eZ<B2#8?S1MN(0_)d)4a_3_X3Id[]?+V?MV8Ed/U<VOV#
3.Jb8(Ue4)<YC68L&@R6@;A0]@9<QB+OX;SC;U<&:c9gCES.a//S>]_#4F?bNROc
PAQ4NKD@-(<#D)N4AX+KdPd0OVb--]AeXEX,Jb9fB4.;F/T2X@/F\Y#BN=8]2\?:
cW/XTcYCC8)+XX4Q4AKIZ2,U>C;WggZ<a>\RE@T[OJ<G4P+6#0YDd<d-KC#0X8Tf
F=CJ_gUY(8?^Ha?YI7N6&3R7?g=4?#9+G2.8R5eYBY[G70MF._cT@TdARN-dCd13
ZA@QOJS4<<<?bA_Rc)K2F]M1cW_K3/a4Q:,OW9DUc0(8VDGR=S.G4(-W6Z8a,-f<
[f4HdPd:Hb(0X4FQ.dLZ)QSL2&7f@<LYV2OZL8ZVd]9QNF0.DN3Ug5RIg>c,X?P1
T@(OJ60TSZQ=?F[3^OJ6_40,2QgA3O]Gg>DWO,]P4dHRcR2W)N0?[3]cK-1YN>Ug
DS_XOYW]=S0OMcMXb@@dL/S]362?C_Y+e7.8VaZA8,,1#1\JeM+LHCDFUR0G);8g
F^6bUKBQ2(O93)P:WX/fY-aX:G9F3a+RZ&21A^UL6F2TML).L8[,H,JF8=cJaC)W
9B<[J_c\H)FL7968c_Y]4;\.b6E:T^[D/H:c<a4/\>R[R)ZA<YJ5[M=Ad-V4Xe/J
FHY;VbW)2J<?G^f@\B8B>8&J\b?60:W^1Q)[ZH5VdDH\aN;D.OT5]e\YGaX_g4_:
?23@1^<^-E1OcSef2FM7ZCAUgdW?bfG>NEH00(,(1<3K^-6-9<2YZE1EO^:^[>MH
RJ2gP5S[=>DZ>J=.c>X6bHREM[@96[FQI.3S@eL&^)a(Z@;#/b;]8K>3NC8#Z6C\
HB<1fP[bBCbQ<a<\]1Y3<J2Q3\JDg)?PSB(eEG[YOSG]BIYGF\G4aX1Z.G:b^I>>
=G,-5I]TBa>N:5eW]4-8^_X=0.Z_[89U]MSE2+5aWaE)\&U5III-E#\_0dcc]J_;
-+?0+J03]gX2PBRc-bTH?#f^6^OP(,egJ3TR<g^)6Cca6CSB>30QSg-IFRH2=M_+
QQTK?QbX;9E-V]R,0G&gPT1QC7:I1(NTK&-5b>1LcP:(T;OCS5-7d@@85[<#<#<#
3U[PG9CUT7=4WU=<eL)8V_O@Hca/D<Qg3L5@H9dU+=W.,C#3SR(Y,><B:W,gTI(5
6e2SG2W5/AI2#U[:Z#\b=g72b5cMN6da??>g1MQ>/dF1N#b5]DdE)MJ_c:aV^1:Q
YZI_aN20^HULERMXQQ83[]\_^0b<EI\JK7d_aW(Uca7H(@RVT)4B,GFDUB\),VN7
XJ7^^LVQLD<Z(+cC\5B->U7^(J4YQ3bHJaeF.SK>RSH-P,<+-eObBg#5Og,7++3[
J.)FT&<?Xf35RAH]JEG\T^R:&+4O=LGLAGd,)f]VD3\9JLZ<+[(e<]N>N/Y=4[##
Zab:OCC=BePZTSB(B-\=\GW),Rf2c\WB,#S(/I4LQ67H(]DZ_CKRWZ>I,8A+M2WI
^Qd9/RJ=J@=dT69QL;UQX=Ig;LY@^]R[&U]6P0/g.BQ.K_4Z[T/VK),/_D/SLM?C
U,4fS;8<1F,]g&MW,fdO\OddbKdQ5L.1BA>.P>7CXB(3d&XaFB/\VV7NG<C[3b;C
e=)KGd=e=)4W7aUXZCAK\W0b8@8a:P1dXa;eOQ<_gCgFIHNeBe;;#@Q,[KJRKdgS
g/I_>46,;;Ta=OB^ZEX+-GU:TBT<-[:L8LQ+6^]ePSf],6R0Eb87CT]@,9bZI+);
4^H;FTWO<4ENA:E<FR1:36BVAf7)3H64C0)H&@S=)BH;EGS3&OSH_9ACBU_X//^4
K3Fc_;V?b4VH7Rf9,]Cc.E_R<b@U>c9eN_&9J43BQT>O:bdUSNBX]RO#(#&=)aJ1
+>+bIcA[0\e9>[]34JT/L_:S@=Q9.2D1AAeVXbbV;>CNd,GdW7.\T>Xc2g^JI9CD
FT9df6G@QR]#OG;GH:YDF^f1FHYBAdI)+d==MHeIC[&V+)\J<<M2^egV\AW9W-R2
5POOY4F.)X<(H7@098WBN<WW]O+eeF74X6K9Q6TV/G,?QYUS=VZ<5b0FV&]XNI:9
T-g6&?3Ca#g_A](5VJe[?MW9=c9SN8CYJM_5+6+Ud]>G-=7WTY+.CBC>f)f;Z.S8
E&ZMVMEO6CHC5<PXcN.::+QZKgg:G25=bJ78Dc[@JI^c;cA:-5gL3:(Vg;SVEB.@
).?,8/80(Ggf8ML9e?X7K#ZB55ZKN;G]^QPDE,XP4TYT]W+b.78[d(O&^,#P-7LJ
/Cc4(DV6Td=F23gCN_@71#Fd\7RIg8B0BUPYOP3^1T>cMIa^AL#-CJD-O[V65K:Z
e7?JI8TI6TbU1V\K_I5K#A]AYSSAS8]&T2P]g[A5:AbTGR,&P90-8.?F6;IPH)9T
+_8NL+J,O,:#;9.;VFD((U=7^^;]gI7@<LK<B?N2cRVK81V@_Ab2B>eXXXJJ_\74
HM47b8KW?\O6+-D;cdg(,,a>6XfMKVT+eF4^/IM]f,KW7+&A>d+)\Ld6,RU.dEDS
YJ8F=17R+A/XWb=&ZcUTL3SL<;8AB9I[0LXT5L0@bPA\WE]1Ba1>PNH3e9ZMS/WL
B-8Lf-b,Z\&gZU/8\b6cOD]QI@eP#@S1O#9QTIEHH2eH.b.cENOXGUYHQ0G&@?EL
W_;^L]8E/8#,ZA[]4D7]2F<d3UV(8YR(=;eHY1d/3DR]+;#/74ZR1F-g79-IUZ-B
g;\@,g:UO82E^\@cU<]RU50UMTHA6E54:4a_KM8;).E5ZN[4f\F5cCB[LKL;Z[Gd
TCJ@&G^MP9,EL3\ABf_0ME_)Y(\beI^)QYV;e,@+\P.:L;@D76X.0RIg[NAFbCZ>
1Xa\G/JVgZ.+Q?#0+>P5DFC=,1P\@7E7:<MdNRd14&,dUT\-C],c&GV8bD/5Zb8[
cG/Z&g1I>[H:d1a;M3^4;ZWY2TR4119>0(;G/[LMa17H<?UO38Ue^49\R-0[,.e+
fUf2?JR<S8Mf0LfNCCg(A<VDV@aN2[,@3M\#(RA3Odd:NZeY,I7Ybc/8+4C=0PY,
Z_7<Z[FG<H^cGL@^(W4?_7PLQH1WI/(1K+W/aKEAQ7Z9(Tc-&=A6WY#Q^[H+7Id-
U,Bb&&_Q]V2V8]=QcO17[c3:GN.C,8.\,:G:=0H,\]X2V_27W/eZ^N.Wg+8S>+0-
0JA,dLcYG0\K=L,9F2d-IfSJV.LWO</&U:SaBG-B5G#egA.=9A^8;(?)E4eEeBb=
#9HINWWA@Y2)5O6-UOS^IZ7Yb;b=S67)g:.0)3>FNX0c=6&HG98\-:X-;6C3d1fO
BE<Y\/)JA5FfFGRR=WQ7;X^+MIR38^VNZg>P2/,cMH3-1LLQ\R[Ya>HbTaJ4&eO.
X]DJT(&CH0\)1Ba:c2b2R-UCT^/L4?NCPE8bG.8G37+GPP6HO&XVL)aJP7=d[d1P
,TJ(\#F>L,9bdVgGG)(URCFZ]J&TgWcH.f8<FCb@-Td]?))-VC>>PaU04_2WaXME
B-f(eI6RIGQIL\^W?LB<E0GR/fYf@L/7_]_BA:.:U^8_MX_MF5BY1:#U7CXR2L_#
I]^XUM?<Lc.@MN-4fK8#3D\Z2QC],GPAEFS_dQ,[7:88FP>>QZSE2[;[7LI^_R6f
^0AE^#K4YFXX/=A#^>0=9,C_@Z<HD7IfB9TAB(//R(=^aaCJBMd79e\K-6F[Fgc8
&ea5LV:8.ODK\M]ZbAJN2<A?<^=WX_Bf<J0S6FDE8P2JBe;>b7fWLSF=ReXdV-ba
&F#Uacg<>D23BM/)VV@/cWS?#35_T)QF75?DKJQOUR+,XO/\.aNA.;2Q1U\VEK??
CGaZTP&Z&F_G3DdLb1Y_0S5A2F7L5UYaD:&T7(G5):RIO[(8:A3I1VG[#[M\B>QJ
,b7:]XR[W,B[801b0c-_d@Tb5fIBY,c3S<7bS+0J+N1P6WCBdcBMV3^BN@^If6cG
EHTIaT&b:5=JX3CK#c4IB]FR[dH<;(U/aB<Ic]8gbZG]4<Je?,Kg\O[#OGe7L:XO
:P1cIbLe<JWHK-@AG_8TQT^#87]c9V:.27+a\_8fN+C(,1cG]I7<\4>[BN=/PZAG
?_cS[@<7I@OR\@ZMM73K]3)=?M]M#GH.?\3(]-.a4<TPGdLH/1^NP-1Y+5(-R_#=
Q]-H8bE/WIH@J5G9SJPD3HC2X_DUJTG,7/(]a/-\4/SZ\WW1Z-UDNDP;BS;ZJVZ5
0g=,4TZ01AHS;0A0F56/?3CV_19fWXMH)L?)_B.b;1OHa[</XKBa;,c536\91Qc6
2A37=UM+6QV1,Oa?3QKMRBV4<Q=O6b2_9??cTGg>@CFWMJ)7K^7^&XV]#0,[DBBV
?I^g\]:dX^WP6=.c(eJZ)H>[c=)Fa:K/KZ3-SLSP\SR;B9e?K;DfF85?A^A_>+.G
U5caV^V7gYFX?Z&;d2&ICB@ccXF:?Q9][ZDP09XCZO^0S80-.Z5:=-bF3U1JY+4+
&>?/?MM4U[F9c/:\KaT+eE#Q9I5SWZ?5N4D9&4=<[)bA:ZN@b_Z@_H3U&);36AXB
Y;1]E7\)C.N:6\0//B=d7D.agb_MX_TL^=bX#^gXaQ([GBg_.UT[]&6]H+5TI/M0
@::YRCDN?B6<+UfZ1N5aUGW56QN01D3&1=8OAB_@aI<(S:M_X5.DFG:AdR5?(/B9
Jb3g^WIRP_Uc]<gW5+:Y.MP&,MM4FMaGV3?,P(MA<dH)G02M_:aNG=[UTe+G/G)S
.2)3]eBa8cUb)P\[c0EBD9K/XXC2C+W4ECB^A^V.BJ;.NdVWFSSR6cS>PAN;;3#d
HQ/eIHOIeA.c6:K:&5-I2QN>#V8^LO4>U=8=N\\/40ON1SS+S-.Q+Va,7f6b@dAJ
4g4g?b]G&=(HALa:72MHaLA5U?c5T&FXe9NV,L]_6:Mfa@C2f?\\/7W3a[@@6N=E
0::T<Nf\>a48KB]?-NV(g0BUb/9aOCD1N0M:4A[)6SQ34B_8bGVM;29P9_VQe#M<
a[4<DPfc#HD7]2\4b1<gKW6BaNFd,OM?L^FJ&W::J[_&ZY/g+#bfe0gVT,7^c(\&
7&X#5^H4D1U7-9@\:ND7JP<)XQK9B-81N_),cU1)/3QUZ.7D25KLRR0F1BR7JZ)H
1K7T3U)\0)]SKH9@,4N&gDA^^+?+b4f+/#RSK1H2eV20>,\2aUMKD#G_TNV&27;H
/T[/b+KgR[/V^4?0MgHQO?PNQ-H7TV>4&IN.YbL\-GXXeRI0BB_MK&RY[F&f43da
Ad;\Sae>1R.WB2=f/^)PRB-(&R(Q0WGYI@9-(S5]:8,NKdU)e+Jd,>?Nc&^]Mc83
3CKV&_(XH-5DWP->A()O6T8C\IEe](#bI/E4a,@+Gf(R1KR?@IYS>/Id12O9552W
:ILN,[=/((&eR#7b>5P2V1,8UCOK(<CSO0RZ7AHcQd8Z?.dLU7KE3g.CcUUA3>MO
PNCeLUHHfCg3)L&+EeX+;>B+aYK&JI+PK1@1NL_1ZaVGA,-0ESfFB:Qg6MRY#Q#?
&L,#>9g7W_2-CAAN\9;X3a+0]b)@/#DW6U.0=F@(IPO7=H;?Hf,:2)bFWOdTC@T;
]WOG+=.Y@T-Y4A>ScOIJe[SRRB,<.]@#]T9?Y09\6B\LGSFCE:-V03O/;WU\QZ<N
0bADGPUZPgA7ZC\c<0a,+4=VMDJ_.=#,a_I[d_Tb;.C]T^6+W>6HCa_.eZJ1C7\+
O#R4@JGA;\(JQ:?FO=-MC4GA/,TZgdPb7P_:JPLaZQ/R(e@/(+#3J@+:e8Y^&[;8
X@[D32/IJ-dB>/^4G=5PJNC5aMRb7/4L)6NV/A83S\N7f+S>cC=1_/=[,<;TeN,P
<Lg[88<4&(#:K1(=?Y\eF)R;Na@aDc3^>E4^^N3,BK;G@F/3MGHZY0Va9d(6HQPT
)P_8&&/?:Qb7L::.RWA=O;YCG=6++C[R^-0XT=V-,6,C>)+.12g:>XMY;.,V&P\[
XRZQZ3\TQf<c@BW,&6@N+AW2)YcA]FH3]A6>eOER#,O1\OdLK\M\#=N[EM7Q2c;J
-e_e7L(B>a&7.U>^gV,_M_T,&U#OXKYc+=.5OA0K1_PYJfGL7c1JLAN-U;4.c6,0
#gC<3GS(29KV7JA1#89eX_]^fP(Z536#;TG;W7DS3d;[/,7(>5O4SKd7^48+\U:?
4:d=:21ONF.]/^bTWEX&.11=YI?Y&1.ZV&1\WfKI@?]>?IF+<;bLWIL8::=^5@A#
DO/b9E1P0#EEP=92</P;5U\\6_7b3fPVcI=d-Y:.dTe\T[\(=/^+T/DIeg;]dN(U
^NFO5P+Tc^Nf,O5bcPJ[&F=.\83D0P8F-UAe+2e^U=6DJ00AT:YRV_VR^W1[64F)
]UV>ZRG9OT[?PD;aWfLeIV?dF+Ifb(aRa>^4Z>0c&1YXg[J&+46AK<P_&>a08WRX
W5)@d:[NBLH>BG]0e&1PcIA?>5</dLOK\6]g-&=W<2W5_]T1QZ6ECKKO3>YZ;)X[
<&edZFdUW@2D(g(9)Y^=aIL4a7c:gKVV)R..-B,#U,OKF1@N?HO&g]M9A@=4gL/W
[Q2H^PTSbF\QK)7eAfSQ1IG0cYTf#O^,=FbWO&L\25>P3B_d\6;)?fe/AZG[Q0)A
W^;CK+?KNVEg0_]DgM3<_3+#T([2bM)I7Q,QTf@O;ZLf@;BD-XN-Y<;=-G9P7@1]
\@J7HVg=&C^S-\LDeR90LJE7c_NU8Ng4Ac6Lcf-<--4XH?94CVZT7IC2(N5>C.HS
&UAf^-FV9FI-=GCe=J7-2&dXc/Iddc>MbOIIC6(Bb/@LQL1G\Y4K?^eC2;]<=EEI
AC\/A5N,/<KD7g>dKI45CHQ@eRZW1=EBc2NQV9I[bX4gTZ5K=Na4fL19e:>0R]W<
BTUUMG_CC>(6D4:RABUN\O+P-E:-C-CS^TBU<?Kb7H18LQgQCf@^>HZ:(OQD(NeA
(,&g/J72P7)D<GZ(O.Y.TB]#6GK/N./;XDGO_-+9NGc^]Q70/Dd:Lg[-fdX6:dX<
[9>UA@H/T0R&?SaY):7GM@<.JDONOR2F9DT[][32TP0.E6Rg=A5_EDIIOOJUMP2K
@Z@&/9>ASEF@WX0C^N4@ZQ0;Re2M^K#,9.fb-MUYPb+=L::Y/@,g;0(]K./40<DM
[R4Z[G.D:D=S#Yc<P8:1:#--SK.Ig\I5_]RI[/@P0=D1G(GDa#-H.7(,bIQbQ5JT
e,D(=]46>gFRN]42QKc7RGDZ5N\Vb4\X@>;X[E^GKGUQ)8fB7-RdP/TNPLcV_CIG
+VC=9]A-5(B+XAEOVR]+FUcIS@IMK-NB_E(QZ,b8@::b7f,efaR5)>&?(I4(IHA,
dM3GIYCRZf@gV\<Q-[=d,;D#<H,/-UU\MVR5J/[Pg@cLM_5AI7,.(46;=U/)Ce1<
,7c@GMI:S\0#N^G5,)Y>TNeH_1cTDgR(bBETQ7_^b_7U6B14?]NGX>0UV/J#:>d4
]3X_6#A#7BEI=WS[&8@\0d,>T]5.>K;&&RB2OD=G0>]O\aQK?\U>T6&/YEH\]cK)
-4J#+P]J7GMNS1gB0IOFIH3]0K/K/JI-V][^Wd)7cZE=.D_,TMfWLKIdfM7QK.Q=
E.UF)VP7R]f+3^a=>[JU.M?NV;Ac:_:OFWC9P]d8bOXNTf+c7Z^6P5H029OG<IV>
C)_P&-H_CA<LBG,f^9]A-2=4JPc3V,2Yd7T?4e3[H?gaCLM9OKb<VdG:K#/HUTLZ
0X[b2;\@]B(7<(]&IATXdc:1D.&ab\U#MfeJE1[dIX3/aUH7S3FE6f5)200F-P,Y
.#/1MYaUW([W7/L:EeH7B,KLAa>@]FG#g]De-:HFO0_;L5=<C\(#@aFH5fPE-g&5
@0Y7XKKG4U<Pd59V:]<U.+)]PNVbFTacT..:A5C.^G?2,W7e8^5L_Da+F8U1_;^d
A[C,;8L/C\ZC5Ze;gdGZ2N#]17+CVZ],HG7#1_.CC[8J.Kb3FcLKg5YcbeLFD.^4
[3^eb?+X+gaeIX,]B=BAK?><;U:V9#JU[GICSJgH///1HX(HXJ&[N7TCE,U[K^AZ
Hc+IJWT_[D09[WgFGE@CUB?OU?1THB&/=4ZU9]0V,EVgPXg2.7=GQ-)KAWa+d,)E
Re0,OC\47TLD2.4\#X(8BF6)ZNAW,)J]MWHZDc]J7aWQ74;a]gRH\</HfO3;=:71
M\PEbTT9N\#CHgACcaP.GPE)9<CfWf\,ZQTHU]VE^/@Z3gJ2Zg>&A7Gd(:T.:W7+
6WRO)/WSAS?/T-9N51cHaAI<4Pb,UP\D]_DV+38dVZY\(aI?2=ND/U^bDP(5WZN1
EY<@(0]RO+Kf@TXZf)/0cO6aa>Z?(Tg\MaVS.^)@=Z\V16U_GdM,VD;D5X+[bATL
WbR.5@&[RK,,0.6S><13[de]TLb2Ze,g&(US\/3>[)J,]e=>S_db.3d99GEOJILC
R+?e=NY6XBZDTX3\6dRXJ(D8\F((9&Bg#Z#4).d_cgeMVCX[#_8).N0BO^_d1dX7
;=1[013-)NW)ISL#QAQQ_5EJ3?/=U?RYReVRW@F9?#UPNe7NZg1FE)<[eQTcC)],
)EZ-f[1MN4RJA7\Zc>T(I\.dB>\?(DW=<EgENZNe#dJTWTNQ-dfO26f:#:D-J<P;
>3gA104L2TC&DW-<&WVCG8a]L[N;9eIFDIUL(K_OW2Y\7TSWSMM:gJUQYHI:4(J7
6TZZe7[a\8a?Vb4.:^c^ZdB^JbVZEd6<Y<^N&L.KcGUI=-DQffH641WM43BU08:H
&5d0:b5?Q(7]Q9/2&)4CSae:KW(7O-8=8M^dLFA:U4g-<MTcP<X406Y0=>f_I9)_
TP8>JI1?(af(KB+6Ta_Z;=2fORM>Jg]cLSAePP2RG\cMU_L#6LJE8:&d,G+PMa,0
_0HUc^7caK#c&2BaP=dLXARbg^#;GSd>N6cPB6&BHP2S;eKeIVV9QIAR)5>>LX-3
^dOW#MZcdb9OW8Sc+]e7b4B]IXH_T#6-8GEQ@WXaKJSB;d)LGPC=YY\D(@2)dR.P
ZJ9S[BfVTKBX5>N,=F[gC[dITO=#bN0U1WT7&_\6RffPE;?16Z-KE[DP#)6NO];:
K2@Y).[>ZXA:O)O<0K^C[eGfPdTLCaYF(a4aUd8L>N]:Gg+(;JKfQMJ8JXGgKgYE
Fc)Q[TKQA_IDH>/aW]T[D3c]IVCHE\R<IcZ,-VF>SI\7ANI\E1)abK609WbbB6RU
COU>4OT;9RX?D-eT83JHK,/PcIK<Lb8-RL3LcG0D.@gAIE8](A?#G7-WSSWXB57W
fJ(RQ4:#WRVf-=<ZQRH+IbDg:=^LBD2db73gY8U)PO?#X?O\,]GTYFO#K\\2H^=f
_=^=_O>56?F@E98;EFg8Y63UKHC/DYT\9G1de-TCNfIV\3Q[EM:7=/R@@4,UZK9C
R83.f0T?XK2&\>.0[a/L:bd]8F86.CWV&@7H1QEU#8gCTM(P34U^N?WI_[&/R@=6
GLOP,FKSJ_Q@^=/cA_T5AGfE4>5aW-d^4@XWFE,VL+8Nd+4]OB_I#.M?+F1&f3_a
?2dCVRYVH<Q>R;c5>E&\1._d<g\.edFb>_10_EFWLfC/#FJ]=SD#H3J+[aF^SN^Q
CKQZ/FJ2,A8/8dC643Aa75VO[A_:6]#_fRI;AT@gT#XY?CLA,Z#YP^7[bREI(b7?
#CHJbR9T7fee,6b/B+.+e=[;E;?6^b?Gd.TACGI^fg+H9O=H&C2M?K:+J;)-)I0\
Q]5a]@E&gT7@:/VG+<e2/>43U11CagKbD@(d2DXcVJ^YU=,>e7?6D.&Z(1)/_=#X
56@c+(,C)I&,>W>eg=E@];[3bF6K)P2:8(#fT?=Qd&DM=2La.P-E)-0=WaCWQ(4(
::F?)d=,+V_\JUX\fO_[^^CcbYAd-+R7L_MbU[,=3gMD]VS?>;<SLZ<H6)YHPDZB
<[IRVG>,GO[Kd6^6SbU?K#QF8<ZQ_J@RB\N=@be.N=DEXf?O]F3LIL((Ub[4S>Z)
J7OZdeK2aI<F88f_CVT=Ya>6.fX[:c_IR?KYZZ3)ENBgP_NQ9f>T,1<0.eWDER[+
H:f(-KSc)IG++OX3#2DIW<+[dN7?XNN],(7U7B7RK.QW<59H(QU^RUFP&[9,/bWg
1:7T7<Dg,/R<OZ9UC)O1[cbU<1I\Q&T/>(Nb::[#.\A2#EfX]KKFa,HCYfecO#G+
PBDK=d?6(?(_aD22@GX?:8TDaWbD>JLATd1Y+RY&4Z9gfBTQ+-ZMB,:)8L7.RZA.
9L+d2?6dMN^6a^33KBbbS);Ie\=9OFKCfD2ZNO?UE_T_A[^QI^CY?b\Y9XA-G(Q3
8X]1YA1^-_@+AF;DaN3g/@CIY8F77+2_L+N7[.I>XD@<f9=]#P#RdH:,8gN76J,g
F4]&3g6]K7U&IJf,_CM=NaI]=ZCJ3P6SDNb.R8e2g94K)c#QB/2CLCAA]UK_cRW?
PT;?=54FW(DQ(/f2O0I#^#@SA0dWCI5#&R+QH6M[\IR3gT9&J_M<H+/<T8>VKHB&
K]HGQeXaSZO3+L7DbZWHRV4H&UM6=.eG6a2AE1C5;CC2KceMe0ED71P;Af\;R[Wf
&5IT?aP_@)2=-.UJ8Y\W]CL?cf+(a&4L9Z0)WMQU,#N^2[dEV-Pc68DO<e9aBVQF
TT;5/R-R@dNH.a92<=CH\ML?E=K6W9+#D?Z4^YJ2BB8bGO[f+B&93LVWN_18TS:G
2[Ja690A:b+cb-:@:K(F<MOe.b52gF1[O@?985@4GZ3e(BCX&OO[L6<e/G3dQOC8
]d8K_W9Vbe_@&[If)12QTOC+KPDU>P/CB-M0)PH6Eb],_E#>TN1[K/)W-Y4Q3+aa
B#V7:<,SG/[L=P0He0a.;@C#JJ287PQW<<_#Je<.SU=504X<&Ed1cfIXR;2N.)AM
.VZTU>86E(HZ6;BdNPYY/B@(E8I(19>WcgBEG[E4b?aAEc)[6&OT:.X7?+HK]H5(
UJC0c_>53EQdcEf[bYC37@TIR[BX#T)ec=4=1V=Pd:J2YAT+3VJ<M.MZL7e=:IM&
c3:#,a<b[J:Ag;&CG39O_c)O&=@N8Qb]T]>aA2;BQ;M;2#9](\2VXZ32KU9QE4Wc
GT/c=.LWS?+?I\&e?VU[JH[JAWd435fa0JDZ2QBBXJL>8)2D[&U;7K]7V[-OADL>
&/D5BM_R\,/PdG<+]D[B:4<)#PG(J.X_0/3VHLPCY]M=PW,[QV\#0CAe.cT78/J7
@YZY0CMH[:dMDH[<Gc<XHdc35,Z)I7V_&g>,HCF5.3.E:0=EgK0:RMI[LcC)]IZD
U#UM[996&2PFG&VGJHS^M3@.N9?bDONA[]WIS4U.4)^>-=793g2gFM)I+0R;\+gP
XScV&5][E&57T:O).B@>ZHCQP<SF&](OT(;:;[15PSgcAOHbZLf<Z]11QBPc4dSY
e=BY3?R3?]S,EaBGJ0cd4CY,T1?O+LJ?+B<4g/aPL]OD<01YZeI34KMW23EV;DMM
^0M5N.&2K6EVRV1eY4MF-19[Mg(UTYGSG2+c?JBA:Se([54_UN(G,B5^3RHV2#;3
GIG7T&NY;1&N]W[1?D>1<I?M(Naf?2X,Wd^2dN[;8,S2;V]BeaMUd7^LLbSZ+I-K
C?YaR[5@&D,<C/Z#@0#@#NYR=CgL1\CX./:6T;\/]-GS;S9T?OAA]<S09M](3+GT
d^XGYc_]WK6QG>U^&0-P5M?8[A&3HLf8D7N>YLOT=Z2Y7RE&^5fF0_[G_VE0]64Y
I8E5?PD=;6CXdFAbSP@D7B-N4L+ZAe2Z:fBbHK.G3A+7QLA\Y>NIYY\NE:Wg>@DN
/XdFGE<G7-&)(012bHGHbNEBW0g_4KA^EAJ9_&N:57\fgSSS9ge+ZX00E8Y=Q2VF
@XXHGZ,56Mf?TY@MUVU2B;4?JXE6Q#+E?3M7.:T[(/GK9)?R4K-VF\]M3^/MH,Y:
<XA0ZHO=TN>g>KF(0XQBa;MJNc\gJH1::U436Td&/G(-0^EA3?_(^JgQ)U>V)Ld&
+V16PJR9@DRbSL=GdZ)GLPVH1T_Lb.EdNA:POge[b9>]D,cKOZJb^9UCR#4W^+I]
8RMAa&A6=T\1O8^:Yd:5TJ[?4>^ZT;:f9FP^S)OT+1aF5a>Xd[SB)<W&DDAa:-U5
44?]OD4SKTa5QA4YYSZX<.T=WS4fM,AHF_\S>Z[KbFOLX?3+XFXAR()+0M-G_[73
-9)A(SL#3L8B][K]d/8NOB0#.c?#C_]25I1T;HO\R[0CGccDQ1PP)>eP3dV\9FcV
e8>e7@IRKDM1e[7QcMA7c#e#&4:M?FGWS/e1J7AW4;Y236-cRK^?R_OS-KG.+>d#
ROEOK(\>>AQ[L#,Qg(Fcd6C+#HMGY^Q52&_Uf=<#.8;&F4Z#-S1]6W387X9XGB-\
BW3D4T(g_].OLMb_D.>_Q:1?M<;V718L0_<YULG9F\+8,S9aL\=I(a3-gD,Y8)_;
BI9N9BBSfPGO79-9Pc>B_--^HRa3]N53OV,.)0C-4UJ-TU62\HHETbJc,QB=FW7Z
34_M1/a-9DF?E8<0.2FLF_N:5P:@N^\+a;N]?Qe]@L_31#b\V+_DX7cE1X47CD:f
9EV?JG+<Y(RgS@dD0M8D4X@>WF/4];C;WE^:CNNYRC;cV+D\9696U/(Ee1^IY5E1
496]02SOb:SY34DTFI,TT,U0-\cH+A@[(?:.#VT749-Y0P-eb4;1]HgcUA]feR+b
.6P]=GT8c?S<XD4X:6)JHdHG5OW=P=8ENa-X;5dJ^,f@AIf4?99[[7B3#3[GGD>c
LW@,HML<+OP,1N,S\gF[E=E8O<aOR_UOAfZW<DU-7S,4FRLX@,]=Y;->RN[Y^O7W
2BR]?0D8]>[0EM3]JEd]dM_/IWR19>?#;UQ9RCaT2=_dDKa+(6g)2.B7QHL1;&>J
7_#I+P/);;#c;&f4;4EYWMY1-FSLdJ+MH?Lb<.DO:V0.V.EV8e-&1E#UF#Y>Z3?B
HDg,3&bY783GN^fO2O&bBN).X=f[2(g-+[QW+V,]KG4-&\MZR3T;FG6OJ9C83.Na
NL?PGU)ZL]W-PS?@9&R#2d,0f,ON8LUc-PPL6^U2M60Yc#Z/d2M>C(3gQX-04d;D
:Q1<5_aG+c<BZM?d+YDc2_2B_:\<Q,5Bb>5)^6TY<GeOB1cO=fH+a_8ebgd?=>8T
\_IHV85N4+-I1Z\5VbXYWA>X4OJ#e2AU&T[a+e(^CT>P\MWdFY.T+7=;I:VZ=IIb
4cR&J2c,6(1Ng8K,F3LQ-N>Z>DdJ>=dF4PdI24M<AbWYgF?:_AU.a^I(G2##D5I5
=+=,bQI-?K?TS]F+d^^_A(_]4XF_K<]/[Y5AaI-/V5-R/XH&+QA.(;TVd/0Y1^aA
6V&;^O:=+7CJa+Q+C1V[gF&f/@6C#fCZRP#./QYU(R;4#421#e1+(D+&ceAg2V3T
e4RK.P9_OX]IYKba^VEDKIX,@QG=FIK\9:TD:6:VD76OSIVZ#dN#JegD,6WVM1[=
O;M&S,EH-7MY/.ZI0E5f=-[B?D1R7&e<5f;[QY1cT).F3g=^S;Xa_>M,C^TA7;<<
cL4RbgPC_DR&O:P&,eD.BA==_eH08@0g4[.F>cSJB\[f?:(6SR^=<06/[K5<.Cc_
W+@LN#)63(3;]SaF)=,H^II&LL/2MK2,dV-G^QGX#[KCBHHMI+AYd+:+YF7,d[DI
(6V9XA5dX#/VW9XTX\HbBNRI&8VY>@I[<Q@>LZf9^Q>+ICX9LcC3d;FFK\]H_IU;
,O5[0F_eRR<B-YE77Ab6F#EcHO?GFG>;PWX;TVab2@F<\Q-]#HEgUSK.#QB-^dbF
2K,f.a-fUSF66AW-_bdYKM(_=RR@e--\K7K->c?R29eY9T-Ad55R#b)N8)Q<BP39
W[f:He,[U5H:+N#SDMT3ABdNI3+1).P;#J:4C9+2_OHG56D;ATA\A^NA&#Y@&RD^
Q3+9S]:A<d15&GSg1?c^a8?P<G615&1QMHFaFQP@O5M_THCMd?/ONHV3(5.8d&C(
E&:#SND==DTe&VBHB5@5B.P3\4Ua54O[]AO1JTG4S\>CB_O&YV)&QV&f;<ARcS5_
>4S^fe&MfA<[TVCFI63e<)+Xc?b_AH=BL]1&]X6JGcgY#JFHPB8<6=Kc=MGU13Z.
/g2R&TZ9/A[0U^-[B@e[+bG_LM>U\H&#9_,M=&WD=e(&D--Q4H)Q>N>g746aNG3)
T^GKb-:-&[C&&eHG5TM+3U01Y9&M\:0O#I+JUB.6E>-f>Tb:faLJV#A2a69IGR17
0e3D7:U=?4ffO/W6DFEJ.00_cZ7>?18>CZ::^>9cS[<,PCcc^/e&N_49#4\C6AM[
#>K-CV7G?24AI,+;,1d&&cTeGgeJE?LDC2FSQ8C_A-,5N1QE5Idf8gU/<>&BBQbR
XY06\Z_eS?SOBWQBB@86#LD=>>Cd5[)\eL&C]fJ32-EDa8:]_W-F5ALMM7?BDMEL
5).dY?<,-A@C1;Z1e0S/(g>J;?=-.f=KM]N(;).]B+#):/05Jf8ZM.RE)V:b-^1T
aIM,fZ^..Ta4VdR<O7eA1I(E;Wf#?K6:76,Z=[c8P>T9BPUQKA\Q[6aCaT:Vc:NZ
(6dF6FfIVXF>V5,6R#MX@EZM]&QN39_T[QYg;SHP@c56cV3?WXZ3#=aR_.g<g&;C
b+@(9?SP@b@cN4fRD[M.2M;f6S(5<&g5Cf4YD-bEN8R<&.a+aNA+<#2G8>?Y;]+I
bVgf\H(X8Z96bOG>[(>E^:WE34R_XLPNM0NA174A,&.F>KK40F\Ob@+/[_]8,THO
3NZ46ONFRK#\\?Z.VO2RD/EOHHFg@UT/_d(L_/?.\#>/B465=cZLD3MLQ]3/b4eZ
H3fEO[@S<3PM,41?[._DCa<MTeeXbVIcc=G:XR1?dFQ)N5\1QPI\>QW]U#7SOJ1f
.2,[6VU?Z-THQE<3_.IAU/WP<;+<?&@3WaASCIeKd9C,21Y_(5WNU9GRA&eY\8g(
/8^^)dTT_3K6R,.^@\H-)6FK^D_dNAK^;Y=_LA\A9SGM,BKKKW/LdNH>0)Ig333@
DgGG4\fL3>c5.#LTgZ^U[LR].5)Z#NFC)B5I,e[+cQd-LV<JYTFN2)8=<1e+TbKI
dV:(f^PU,6WaMW57VcE(Q1_.[=6FG4Ifb<0N)UW&?G96UcNd@gbPd7IB9E+DB(]B
-Z_WM]I/e0W2C6,[\CN)I:ID5U30c1[]0\eIT\C3RRPOA@?bS:L_K8U03gNc=>P&
B8[Y=?.4KHQ5X@N:,>Sf?S4?I#B)3Ee5[T+[g23^P0.0-D<;(3gCB+@NFBW&L[4U
M?52M7#/[d^a]#0B;9fS(P43X]^^a3\Z[ROS&]b)Y3[+&GA@g;;DYJTX&&;HXNK=
]<FIAN()fP_#[RDD:bf7c<S,Q(KGU&7[X)\)^.;3<?=Q04BMH-bB++BfS?JN=;@L
<S[SW^PQD.Rf_Z76N5V]N>XKJcV;V)e=@e]@SI:Gdc_=/_^C7a]P[<,L_CaMMQT,
?ZaP/L;S^&I#86:@/eJES6DSbS<[-A]Fb.^;AgFgT<P\9fBgC^?MQ8]?.-T#I>\d
NEWagPcL,1<KJ7+^39)A;D[Bb#ARVe;-=KYZ]/41^VRDCU[g7(Ab5CWE<&V=XS_&
)#9>/K:0[b2>D=:R&Zc0ebCEMVd]GX9-@6gCZAL,?aY=>f)CLOOd[?\64-BS.1YH
#QYHN3RSX9gAAF&(V0,HVC6</g)+.8DN/Z3bdEE6T#.+e=WP[K+#B7<E9^f6R13g
V45+6&4?^G8.>MJ+QF7SLfebdQ)3JeE+3NfAC).OM+QZaG&AC4JZOF7YU:]=)6^]
AS>^aA3+UY12KdZfbf/b(-RDcf+L,DEACfIY9I[6;J^8.6DRa-Q,K,EC5F<CS+B?
De;L[+[#8[?((O-6;HU>XfMK>\W95FE?KC=E+9KJJSaHPeJ)&cT^Rc=O<^@7I8/g
[C3AER.=\cS1@+C,Og]cU<(/U;gN]ZK?H184F\_[5DKYD)O]O=B#A_\1FN<-14?e
)_^fXXcM7ZHfPUX6HbJUG:T9;IDY=a6ag@GR;BN1IL+Q[K8NN1\bF44S;JUf8RO4
GP&OgT=.0_Y9;I\O3K;+DM]6?KKKCO9fa8@@WdUfJ6=B=>5Y,:,(DMeSS?(bF[DC
cYX>OGcSCd.FUI+QQ\TBgI[XCAT#</ag5aJ8K?/K]1NWBOP=7-R4Q0:V+PC[[G^N
R<>U>JT(V6PaFMCS2L;+IRBCNPF4S_-UZ8/NZXQUUYR0HN>LCIRaa3K_5b4:]Kg/
/Q+F67-_O=24G+6KCBST5^/)faV]+7&dD-WaMDPcZJG7E2-;G(#Y>,/(Y=V=QOL,
BFbRaN,T#&8N]V4FY]O]SUH),Af8L;8AGV)KJ1g([&EWZ>.M5d/T;:?Da<X,a.c_
3UP>G[8@\]fEZ=9OebD-8MA4W#)W),64J^3,/C6A@2]>R46:PJEE1AW8g(-LMO;^
AP:#)I9Ng,Q<@^R]a?2ZgPObOJOJ8QZe1dJ;HcR9@/VeM>:Q:-:4V0D]JP(3S9IC
X5eOaI_0/3==O4BObIdg8dMQUb]Oc60[.H-0G&+R8=#B#6S:#_C+Z&8?-5/#LP^3
E#;JWBRFVfW:SIR>X7&J4H2KEcL[I2PT\:1ZLfe\IdD3@>/07\T,;TR8G3@@L4cE
T)89Pdc?e7V@8=NV/dQN>632GZ^a5?:G.R\,.D[<I,cUX>79I2g:<d.SAb6N8LcF
fKPC[OSdb(2;HRe5SVcK-JJO+I/5b4525=@F=;S<D:Qg/O-OX47N\;Y2#^578f>>
Qe3K-S3aR6/^:KKELE[)?U)dP94D\eP=ND60UB9bSVT4c<acGI3b8,db5LZZeO(I
W243,#Fc1SN5I+=aT3A6M.,KRI=U2,M\GW[1La63RY3Ze.<g)/gBb^RGReJ8LdS:
TBNX?W46QI,_C;=E]3bK<HJf-M5L_cR+;49+NNZK:,Kc]bEQ]Q+&/0)Q(QGAY&Ke
JMa:^&;7VW87;\PGY#8NSG=e/(.;+&(3EZ[KU=Z,VFI>bWB5dDf:22?QG5GDcMUR
TIQN]/g+LE\S-H-6&&.N&-R^;H@]]3??b\^&9+^EV<4LMJ4EHdAEPZLWOEF+P2ZU
b)[Pe+S3G0:&_0eb]X^4E0D4\K@OAF)\,g&W@,KDUI?GA6?@)EP?0Gc3ATN+:9DI
3e^34SQZOc0g;S2^f,O_2UL8^N@)@R5P:BN>KLFI5C@NFB<MWb-gD#N/(]2R+gP3
5C5IPX)M7d<DaG(]0<M>Y2@7g6WZIQ=J>0Ug__A<75EegTe[XIA8#L)A<e_U.gf#
d9bX<T&dGX;gI@#VK.g+32K04;@M([?/XHABN9H\XR[8Gc7c\@OB,a,C9M/@bgP&
9Y1?XPe)?_9_@:,&>#,VVeSdTa6\6(2PTfD&#Q2g0[fTYD:UD3HV23.aOGDd&9-:
-#]^3@9e932Nb@L<I^.2:QK7/O-a@MfMCb5H#]F3MOGVQ\72Ta<(X#4e1daTIC#T
SfcDJ7DAd3OVO,>0X<+NdQ@#O9&d>AQ1d+U5Id[[)M.L.X0J0YBa&=_A/)VgW+L1
d82F0XMaITBEKKg>VN?;BHV9-d1T]J62RL[:09.J?[&-Fc,=/O9T)ST/dT6CS7cd
]O6X4OeLaRQAZ==V_03=/518+#A[,/10OT>eZ/DRI5JC:(eP2JL5IX^^Z\>U=Y4K
,^MaBZTA]=0d?0#0T.,dTP6/X&bUa9E0P5c^3c(JcXc?DJ@8,GSHYRL+M(2WTG_1
HNXX/Z\ZI<MTL^T[RAfE[#acH[HgJ.B9I=eY1bDOb^\+?a<B3b?_NN?bfcVF5XL1
QfcP162aNN+QPCKBfQE(U5)18-f6DLJN-OEV)f,05-RCDef>@.(4bBF94[I>\+F2
ZVaTfIKHYMbMI3LEIFTKAEAF_E#XQ_T2@fH,J-Sb;2H_9KS8Y.d03:Y=d(f,;gcT
?KQ_-EB_K+eRI8;.Fg,AA4VVgV5_5I_Hb=,aZ\IC&M_,)60#@9,?;ObKfFe(f<_c
(UIO,A5bc.8SQG/L3g_eF6Y<HGY&FbbPABGQ9fL1.Z&Wge7:9cI>OQ(/#OR/c<2a
RTYVT=]3SMA_6bM0S_^<+@M3:;6S&@BNM=3+<J:Z3M5KXK\gc?,aY+)AHMBZ1;HV
CLW1db1=9.B^GP^-[fDcH>7;.&;F>T;MCWe?d?T[_?AS,_MYJRGOT?_-ZN><MAME
KNV?CK=,(g>V#Db.+g8,-[+_C](4N6>##BHc/)0eO+Q@^Y_9fC=bL^R1Y:WCA>5.
AC)2gdcMQg=]V[,.&a\&XPR7]DYeKY/6/fTGB(g(N\1_#[a-bU,RR)YJA]BSI<e3
+dAOQ1>NVRV.VHe1,68@COKU^2c./(:Q0F,;>P^eGYL]HW72YODbJ4fe&2K4dB9B
.>S&=HNZAaFg1_#?FB)^:++4AH#=:H19Y[GZ-S51\O(WRYK6<_e]DLVIS,)3[=N.
G[\(F?RHEbRc1e<)VbWL6E?7[6:<&b]Ta@2MXTQL<MDA7UT8N@5<^YLS=[HL=\\S
U[Vf#O+]5.+)R<g6@D(78+50P.SE#=G+NeBR6KB(MI78DDGTZZ9LE^E_V^MU9MR-
22]6DDC20J]]=G1FSP)c_3)>@E7R@HA3JG#?<^a?5g&5a3UUGHeZUA]0JbX8FY^A
IReFOfJMV_YS1#P>G2ac#ODAJK(\1a/9)<M<Ug<IQ;AJ=5\:E2TI?>M/(O^cKWKG
^W)MX8YV9_\Q:#/\9U-\LU+5.C:F0LAUPV&O]#;(SA=DVDIUHA3;abWQg<)5KKCD
YV\AHN-Qe?EEIC40+)VLE<92AF/&dZ+M)Pc,3T_K98\_RH^KbKQVB_S>]P\aCA/d
BGAA0b]H9\;O+04?<XF)EL8W@e9LHc19IRQdc2=^<XH\+0fXZOOAL)RV60SP+MaT
G3]UY7V)f^FP9^7Cbdb<)RW06L4c=UU7>HI?UQ4?8VYH,fW[3A+)E=[,C50;\19Y
+.Pd3SH3<MXfaSEe;:9_.g(A761X+VADOD?-Y^<+O[3N(H[dYN661;L;TKF]79N/
&7/8FL1/,VZeVDKGZdbBMW<XL,GR@KDUR>P=I6JIU^S&-\4KdQT@/NTGD_T+>\U>
:^dOU6\3D7]TM.gg2:54B_-1>+#EY^g,DQ:<1@9LL=OfNJ_Y:g6>X3BSEKWIMc50
29YEf1UNCW@8C:.]6_7cAPggF@?MQEc+I2SAWb),7,Ab?O9I3>6c[AL9KVaD4I#/
Z6QBOS6JV)A>^:&YO:0aW<DgH]..51:+T.fS2G@L;]_NZFB+PF)GA,J3M(L4b,1>
LUHG,Gg]^R-\/U\N7cBY8JV4fgaVB(.CHN3^B&[N^--M[bU4-GIf/N,ZWV1EH[8B
;72Nf.4&2ZQ+f)(La^d]BYO8<H@BI6Q<12<<ZQBWUD,V0NR2g,>N,1:.T^G4O-;E
BIYU,dG^B1GSG\QUda+C(.cSEG,.?JQ2g=#V+/&@1@\=NQMUW#WT/VD9GQA536JD
SN/[_-aJ<54BVa\dS;c>B4P/+beLM1].YJ+CFDD=[G11=[XWQcP01Vc](#e1c)W+
gV^QJD3NE[-QA^/ON\^TJ^LRNE-8)38I#&#L:;aC9.R(c6H+970P3\>EOed.6,Y@
YR_FX4X&+#P8AG]Ig=S3<UNOJ(?/ZNOcHTd?bBaU2BI=JPNYJR#./eC2/O47:5\3
-cAaHFRKTGQ-SGAW-CQ6a0DB5V.FAa?\O?Xce3<H21F9&Pd\];HE,#UTVWZ?@FQ4
+6Bbd-5@<5#BYU]GB85L]bAK]1F37>+1A7QD?_9@U(OF9621H[QZe7[bFW\Wd]98
cSDG&5<5TPH2aXVE?GF==,54H:@>dcD+He+?N1@@.A_S#XE?8U2#D&VDA:0;.3Hc
@EC5efdA.3&4F;,ES].Dd0L?8&R.1@WJ>#:,5\ffFZ[<T-PB1bJJWCHG]IYU]4/a
5>a_:bOJXbCLC9TN_;15ecaD6bLJd<W4FUU>P&ZI_bPF+1cYQOD^&I2PfI@^77)N
DC&eC3/@866fGg78X(J&YCE/[g3TFO.=g44223UU1XB3&>UC<9T5G82]>LVOZV[M
g,7g#c8/=G]0(8H.8a0>81gUWG[-].CZ\a)&Xc06LC>QER]]9JPgI(:3J23g04C1
B_f]K=I?UK>LM8EE^]RZLeYZN)[3F+4:(DSg^=H=3Y^3YeT&GV:H7#PJ4@N01:\+
GZgf:Q:gae5:CV9=/gH=f9@_/SWf&K&L>fN=?(:8&@4XU(V.N@aREaT/GTSQ&B:_
GWD5#=\_4&@f-X#Eb#)[;.gZ4M.FK/aXTMd(/BW++(,(EF<@[3SIV_?b&)7(H6))
JQD-X83VY==O(HH9NP(S5\A-DbELe(cEJA0fc5Vc)U-RD^3VZQbT]\;WM:&VY;_Y
)I6X_@eV8=N1;2QAE.aH>332(Z8A/.-CN.0f,fFU?J(C9:RVY^&W4XNbL3F@R^9L
)6C_0(+gX=FcHPD\/^/7)Pd,YD->D&4/G<Z^3GX188g)GHb[[8#F788XL^I+?_4T
ENL=?Z-3IAY)RJ\+T1RA.L5,PfY-KedKfN)#1<,]OOFHY<Q>PZH3d#)I<DD4)^9[
R0RX?/gF+C^[R\FXVR/-Q.PAON/FO@[c.8,YLWMdIBDG/+cOKW.QV4Y&L++BS@FN
M0SB.L3g+#,[d&X^;YBeZ2KIg.Fg/4IQ^BDI#\5XC8Vc9FM_(WJCda</4S[/>[X#
\.Jf6a?.<)WU&3>#a4\\FU<TA5T&^X=2-N&E5GA?Z:?;)@1A.F-4;:2TEfOQ>AZB
GUY^&>#^+[ATA2R0c3O9;(:B/FAf0ZK3QaFFMT?fDQ62Q7@+;NI,F@BV[DHV?63U
L[B5(/NZ-Db]^fA42[#/\eM4GQXDXI5>A,_eJZ,bB&a_^9\EL+23g6LTT&_:.BD9
-YJX7b01BgR6D&>Ga(61+(SDO&3Z,AFEU&B)]_#?^])WcEW/YdXR::]C<^RWe?4B
eeb1+6gISb:6e-SEf]O:P9+]49HC,T5PgF6Ee[]B,=6,a:EM<:b9)CHbT;VZR1>4
+P+CW##<5Z8#K]b48?+;<c?&CIg>8fW_Q/+4VdZ.bXERCOd)ZR/-SBYRMLLH.C&Y
f04FL/#b1WCBJ7W;QO+CPWU-N#T8fGWSI(=f?Y4S=E858EOJ4>.:0MLU?g32@+Z3
AW5eV^N_8c.WcV?BDC<eNR#C]7UJ(7.(XO9Zd+fSZ5:[(M71F9L?<\5Q[-#OGUT9
b9c3ES]aMXb^[7Qg(,=>J:Y?15YJ8g?f+MOI(.9cFR4+41C452Hb?bc^bN@\O=BL
^^DEVNXGM11>2PQ&5>b)38bcLQ1CDIY#@:,A;K3-6^ggD(DID)WB(<7U^-Dd_Ga>
A+OCH_6@?PF<Y[J1Z[Pe65IS#3-GSY2<HQ^Z3gQPGD/^KAZB16Ed:VG>cTb6)3OJ
:?+;aQb[bc[)J4ZcDbTBFCIge(7HaTU[XTZHN955^a[#&8d-B&WG29b]I#,RJ4T.
@Y5FD7ea_T9J0KL)?Z,<N+W0^LDRb9/L4)FAD6,&B+>\NUbDNVcEBRLaaA>/NU/&
/VUeF]Za3b6@;DIRK/[NWb\ec>\00?J1KMHc>EEbWLJV(Ja_8S#RA)MH]TB.1@#S
,&=WCN,&f(Y#N;YLO-L9XC67(&QgB_A(:JE<adg-D1;/O_DN&J:LMYGeWfXWG/E<
/8;5L0g<]Mf,]Q5(A+fS5,bJF((0_U.gY3:VA9BAP:HJ.HUC1.7,6[NL9#)gX;N7
cWB9_XCCAeB:^0)T\9HEFIb<W5g]Y_1YH:5YH5N@7PJ<>=BE1Zg,>O4<.e&eY-HN
TRZ_FSO<IK?e4DT_e92;57](P=Xc,JQ_Xc[]YaEfL6_=F])Ie^?O>K<U[;4ObLJ>
A^Vb?N=0FR#7(]LWEE9eQ)aRG6]_<YeQ.Q=VdPS&O^X2.MC?I&^N2HK&9+\d,XQ\
NbQgdCfC2EM2K<F\a=fTZ/AO?gZX<9[WIIb[4eW;b2R#;c:g@-bE0QYb@G-BM)?<
dM+5YA_H+YedMSJ?RV;5)8IBd(3NM&5&9F-\fe<IB[2CgI,.WP^RUbVTU/Hc4@K&
HgCY]ePd:WR;GBQ4d>OZFY++=bW5)cbeZB;Ybc7XB(HgT(0:#9#2?[^^Gcc_XCA(
G_AH&gV@:UT_P8)gE[3=-(+^3N9F@SJ,;.VLHLXDILI\<:7ZADcC_?b901KH0eHa
,ISH_2Bg]-\FR,F1NDK,H)0[-/6#EcD?+0JTS@aXZed](2S#JKX;?De?e6QNCf_X
.YW319SbP=DD1:/[F[[@UZ.XR55BS(T00HN5H/S6(U]-F_-N[W;([2Z4:;:P5f)K
A[Hgb6@<#D\B4=V>S=)c;eV4&a2-<-=-fBC=<I9?75E0]>9^_=)ATG;Cc[c\&e@U
c;BId)?NK5R<O.F:,VCK)??5SHag]g75<MU&&X.I9>-,_H3J.,J0cJ,D9V/3K.X7
LI@>1fOA#E:H,__c<RS4/L,A=RJOPVXVI#Cf2OR4Z^\)0R;<0UUcS6HU5NO61Ig&
4R[9++E3U>Z;UPe.F@#WAY(Eg_A0#RC3(gV(1W.,<gONKZP?/#9[0U[?.2e>&&?K
>aQSOEM5<-)TE3AT6W\-D>b8S&e#07AaNeG^cDcQ+?#fEEJ,(K(:DJBS)5MK9.]X
A<TJ+);+@AGL>^,cc-/:RAI3NWc:#BeHQ_Q1;#NUD.J:&UDRcQ;:&(3S[/Y4c<_]
6\T5/\K,RKVLTHS.ATK77]XAHRcG9UfJ4Z915>7@?W2>,VP45L84GCTL:(=?.60N
_AA^.;=872]?+V-91.K[c:SOWMd_=H>O&a:A55D2#ae:50,61?)^b-AZ;[2],dK_
6<+5E+04]X78dSG.MT6ADaY.;2<<<O\/_K7+\Y3,[b;HUCJ+PK@RO4#-H76U>6Eb
@_64P30W#g>[A-8//>:R9:D(<C^?5FHU6MB1T25=,?0?eD9LQZE231B>>J:;G1L9
eZ1A2-.(agR28,HeN]c7]0E-K7bYS_9\3DX0)_RF\/0LY4e:X&4F:M4Teb<WX^@S
B5ab.W,9[)??==;0gD>f:NTOTeW+YfH8ScQDaL@CbV9LG^4DKDI[QYMf2Ne9Ye?7
],7F:3#+/\+<.)b;5/GFgZ;adED[D&RJ+-gT<&BReX@F960M=-[&?HCR_,#20bUN
TU[E2LJE\0+4+IS^Q80J/cCd4FbLT^_UI.13ePdX<,5_/#(-aac&EUfgW8:1A0<;
6bWTg^S^FF-XG^@SNT1eECaVS3cGC8PD7H];6Z8/bKgVLPeV<19ED;8]a,J2&I,b
c7V&0VRd9&B#V6]8CT8HZ8HD+B^2&[PDV5#E&9,b&HVX7X[65L_.fS/2e-HCTCTg
cXYHZAMe)K5)]=&#,E0W^RN,/T9DW#^A>[2cS?@BJ@g<=F,0?R:)E617Z0L9]]T0
#HJgXR/X:I00)DV;E7_:@VA2(a<0QE7/BZ,4-GR39;++/@0G&Lf<_F9Y\DWAKZ2b
8H74-#7_/[Nd#J>Z<R5.a67FFc+9F3d]DTfAHFKR1Y-d42L13dMN25ETg[H.;62&
F]b.\c5_<:\V=)Q<O\a0R85dIK^L9[+=9D&aV2S?bHH+[4@TS^-^c/HGTbR-7_1Q
6,J7\a-81R?C.99X;8NJbRV]f[HVScDgfSc\g=Q.K>)?]SaHI+\+:f2#aY0@ZS2:
N#+Xe<9Q>/K?L.QR(U]#P#]F4,+BU?QP]MI_)3a6-O4bIE:\U)V>G;fGU-M6W[+,
OPf1WJ)+V&FQ?L5KgGQa96^PB1]AN<BL@R1R8XXNgV8\X)RUb\_4]7@<4IF=FHU1
ZZPg@N#aB<6g/-b881RBg+@^ZWZCaZ:-BICH\SU86aZ:/53K/-=J#cWUGAOR:J=H
?-.)eY>,C<f/Q#&_26.CRG=62c[bFV5,86DO0@<M014096)ASUN\NG-9GBP_).;2
UH\C4M^9g<If8#/+G2FXOdDINX.P:SBV@?ga1:#>+,U6PO>+.V&):@#51TUVH.\8
ZfLY-\JPO?U2R9VHgYDF]@2Pa[Z:L)GDH]Pcd/+aZfK_YeW@aLe,TS[cLIRQ_EHK
Y1<C.ZUXI5cD;JCR>R3G^EXS5G+D>M(DH.ODV_H+:c_#a95-P-1-MGB,@5ZG_Ug(
9G[O?Z^,.7PQ\.00(]]FC?P7\FH,_,\Ka/TH4=8WZLH3W:N__I<RJaMYdD@ZgKVV
DSJdNXN01?O?.RJZ)Y<;YN>DG;:8@d/)@K5(3eb^7QK?g//T5,#\Jc/a=eTTBLC:
W3GdBc2?^0,TeK?7MQ2U=LZfA:25e0Y=O;L1X:H6a45M5O7+#&:F-H9Q&8V_X^<>
]VM[/WX^Sg,1Nd5.,ASPe?CQ>WJ4;P#_C0]T:1+G:1AUJ6(BV/,2FL:_^;<G(+5@
R0Y3_KO=Cg6Q/Ef0^PTI:>#cNWg.H(GOe=<#d.A0\?_VN(IAGaUGaFZG?8daSU<^
=<W[ULFab^284H/ZDTfV^^S@&e)M.H?QH8HBX#d_C1fPfSc#S-ggGHPJDSb<1K7E
&O_4D>&0F4:g(#]9L8@_F3D7:LNGT)?_F].P]^TMbf(FIX>/O7PT?.O]:6U)H\2V
9RVW?&bC&1PYX:c)EMDTf6P(E]W&LX+T:?61Hb:WKRINdB>Q6,VBdB;MaIcW@1S/
?1DB_4]]@Pe&F-Yc)7X72-bfc&X]#YeW1&=93@I.E.5):LM4)b[8+F@+I4@Ia?d4
]D7N4[8-\,W@]<4P+1Wa#\S^E223d(MHf4O.8;eN^L#_^;^WWY5Z2QM?NYLOa(^E
5):UM/f&G0=/#FBM.\RTfe^V:daN<.Q)E7.AK7b=#;gY/MR>:1-=:DL#Q#a:)G:#
SO\N[:EaOC9eCHO6^PMF8E.6.,aAJ6@W1[bUCf?&UO-,8KI_<WU,33SH&HE=(8\)
SeZJZQbKfeMGKLd#BJe+1@,dU;.A^CCE+X@5Y7>UFOFcHfaPM-7fB9&f?C/g@:Ud
K&^K&.N>\BX2>2c4aGB)8-QQ]6.MVC#fYgcUdf\DEB#2ET&5;UM_=TYa0+](9)^5
L9b#/6:5L6^N<V.13\\]R^D6Y+e.ZQ(aCGKK+]KFLSP:bC84;0aF7:>Zaf7H\K(<
1dRcXPfQ=R@W73+_YbE6FTUETg?,FPGa[;@BHfgaHdGD+>8_a]6D,H,#b6:S.^@U
:FJ#Xe@VJ7]54VE[IP2;B5-Q@-I<X=Bd(_\0ZK6:f7eB+L<6XZ.U4JHd^+1e[0>&
g^7+<SQD>^V_PQIa45>M:+(L/E1@L1X1,C1Q>P/f,GJ^#SFG@b0;7>6C-9W[eeDd
<3:>Qc-/S\b;LB8#(dS\X:-;.]Og,);M//,3S+/6fQAZf+=NW5;(=K[^0YOgG@DU
=:e4:60aD#da27/0/J^KU@3gCHHa8-F3MSM8E36e2.K0@_5DeUH\VR]9bg#?W@)T
X2a1Z\;M:TD3+d(NBEa/0Y2V6R.20[]O:#1F0L^(R@a1LJFYd+AB#d#28BMS9Mga
E1cAI:CcHa6N,]>#f\^]AMT?YQB2@D&+?b8@SbQW_@C5X(g?eTa;&QB&F#^_Q,8?
ALTC?V]87[Y+&8_5LcPQ>&.Qb],UV)OBVH?LC?.R;3R]c]@S-T<LQ<HJE>B7c+3#
IR7P>?RQQ0)6c<76YbBW8#b-/RUB\Z.@7RKgG0Ladf+DSfTIfP=bFST6=VJ-bEEQ
GNO>/QgJ=/SCF&)2g?7\>)483\86cW/;@f96=/^:,=98TS45g/8bTHMbB?P/^,^X
1EJBgR;Pe6]87SZ[MW+O;cV/W-3,D/JJK\0;[@OeJc2PBMeXdbGIeYI4&OgK[F-F
JAB>2\\R@DZ5cV2VM>G74DKS0&bBAKR-G\(e\/U@;X0BTK,1(eD=?4d>R.R6:#&a
b(C\F^2[[f(Uf2QbE?2\bD<KT/P?9ac(g.+I?DS?Y&;P9g6BZV.:B4G:H\PUI),?
Z=02ND:A&V<X#6M\6b(D1#30+5/RB,E-@3@B?9d&UU7\SL348X7XKade@DKKJ:[8
E2eD>KHO7b][U/D#V>^gM(>1L[:UV^T-YCe3>Q,3ZRGBJ\DG^2S_]^K/0cLK=M[O
0D=W5AYUV@C+O<dZ_I+3^e@[(OYA&0WKDV2D/CaOB8.UJQ_-4?C?L+C4Ta<YSbA6
ULZZe/<<B#\XZ@)00>#:XSY2NR+bY1#9KBSS>9.H3G5G:XSD-4??U04?S>;EEQd=
CD]^;NWRa?HFGG:9&K;(bP+NYEg#PE6A1g;6T#F@Wc_MJ/5[7=fMAJR7Z\T.(6=Q
d1:2CGD,EN7E_aAN^\WBYFbB1,Q?dP>\@>Dea?K&^g9Ec68V/UEY&b@OVEENRgO?
/e(fGVJ4-.a9V/ZKIc2(L]KA+>dYCNcV(KL.\RMJQ5F2g+Vg3UD+/()8)^0&dIBO
>Sf.c2e+@WFA6H87V>&,S>KU;1/AeaZU^Y_0b(.]V?1Jf#S32ZbQ,-2,,Le-RQe5
^M>2XMP^M)PagNZ8gWZES>V.0KK&D/D<,QF(@T2I:>CJ7?)5)JROWWW9@K8J.RPK
RVE8<&7/J)PdW5(cNaL]HO1SD,aT#N0BOeAB(ggcDYUQ&VQ9A;?Db<PaA<-6NBAD
CM^d^S^LNO&LU6.<:aZW3I,+_\WVPe9J+b;M7<;ITdW#3HUWHJ\-3-RHN9Q#CQ);
Z42)D,Ree7^9<O8;;]D3N1@aO_^SAa0:LYb39Jdf9Nd>:QNUV,1LK)R6-4/JS+7.
:R,+=PK)&4090eb+UNI]\5UddFV&3C52_gMJBUd5)63,;Y=&C832eHYVGKZOb&AY
:?R19I0.PQ(NHAIEDG;Jd1Wd4XBTH_?R8+00<ZJX:Oe&Gd^])cea8>])+C/a#N23
C(FVJ9NNNgN2e+)N)?>X3I,DeSVdc#.OW/Y>@98N_4L?gA[D:5aO8&]L-0SfM.;R
ffZ;4b3>]e6)(5A=./+)/DX8c.2(Z;QPGRc62AXZ(+MU^:Yfd)4&3fC[2/IP3^[J
Vd?YZN&<,SaX(=-#R1D94;)M6N5b/DT8YT]E=+EaBRbQ7CTg9/W)>T/;6#0CI/NF
MWVQ<7U)F2S/e_269]94DDP9X-P(T_DEXQE[4,:c:\1:6(Me5E:=37a)(R(7,1HC
=:CPX2X(_=(5NITH8?<R_WV:TFUS/H\45FaH&4/1]2()]J3_TCQ:g/KfYfgccKDO
QYQIY^N9).:aL,>R6&)WI&)B=UR]b8T&b3+P1W?VdO_c:a0g)W9BMe()G-6cc8\V
?O53MH<_;\KJ(;]N2WL(Xc9gR9[(LF/P.Z,9G>XK9T@,9@g[SNLK9Xe1=VD1)aFA
8VU;&YM#M)bI^(+)<WFCg6bEeRC_HcW40[SGK?P@W,E1?^Z1EN+4@AR#K1VB)8W+
=W3aRKX\)U\ZgZb1aGUO2c]&a6fD=K-d#V@>,:G1_NTQF&ge;JF;TE^c+?^3ffFT
---27Q1#/9,I7#_U6PEN/D-;SWIB65\OH-K(c7bDZ,7KT46L)D57DfW27[g+#:->
=Z/CJUGP^UL)cA.2]34CgT<SVQ7Y56=M+b,aegJ;_P\dK9Ta57\F63F\(FBHTP,E
McLX>E)Q?KbNOGT8VO.=1<>WEFKRZWeF#8J&[KQQ3,+Ne2fX>(6+0W,;K&=[##XY
f@X5.ZaX.@<5<+57M^^UUXX^UR7A?YYg]K6O2>BLNVHTe9dR51](_HF[G,+68A).
S4^&(X@7YFJ&FX,\g)H_:Q>1gND,DYYLG&4-a;49J<7?/I8f/,;U/HMgM.GZQf(c
JRFJ+66QW6[f#UWd3/21f#K9[K14e18&.UV5NF7SA93>BOQ(^N+VGHB73&&UNGCN
J.+,f+,F0L&Aa+IP/^H95X^Le@O\AV?>gLMYd_1MEL8:fg[?,fFa&O1H1b5A=]g(
#&MUFP;?f1GN4Hf,d+/F6d;5Hb\)EI9dV.ggc2031\52Lc.(V2OT;;ZGA_=[.0Q]
[E><71OAXgC4&gYR^eJ38;fc<#QLS66HR(U\;\KgH(VFdbJM_=FdVN\YZARN/gEO
;:0902#:P&Nf?#2)EY8=D3IP1Q&D<W]BPYFZE&_^IE]1#b)RI^2M#BODAU519[;Y
X9-</[TV2JF59[-F@?RU_P4Gf:L)]T.Pfb]RH/=)([,c4=W\M>O-_6@7)Y-D5^R-
Y,M4gUO_YVbBY;9\MHVV[&FdE5EZ+)9W4LC&,#EC=_K\.PA7fIU?A^KD55dG\?<H
eJ?c\^6[_]/9]>_H<8g&eR,T/\N?=_3+:2SMNc9J:<W07eWaOLG)?2ZHPY1?Z<R5
RXCY[4[^29LMU3P?.5QFLbD6Z,f8F@dN9^)eJG\B#Nd/V,4COPDP&aA(E?N)Ue)K
OFDK@b?11dZ(bXG;V;TR<+eKfaa;@TE2]f>]9ea:0GE23[]1:cd9=&fK)J]f;J;Y
Q7G=>^_cPb:YN4N2beR^XD:T.Lg9Sc0)X?7M2@6RUDYMM2f69H1ZXT7F>V<C6=.R
NSDf;]bOUI3;;R8][97NBPB][_ZYGHLJ<D_c5FHQVB>],g>:97:A?<:MBAS4g?SG
=H2fb4,N.RJR]H(_L92F49MOI1aJE>e<]YJSTL._(fS_W-LZZb2XP:gDN]]&UaV&
1CbEb->)@63N6AB4IN6AJJU?8=OW@0@VUW+OGLN?BEcSTEXbg=N;K-^=FKQ0c:[_
0ebP97?1CBKe6Taa.<CWR8#/]E]DKVbEg;f\]S&cTG9+?#&(]d,-ISB]^2HLFdOM
)7YUD9:cP2S:V;.YGH>R1Z?>e@1Q>dD4^I#QB_>/J2fbFR@BJXB-H9GBS+F@g)C]
8\^=AfgKP\K6@g)XUMdOC7WM^NI5W=AZb53@bebGX>N4PNL@8g&J)_SEMWS?aBYU
:,b7YFfKJ3UGQ,>KA3R=8LN_@L:d5NeJ:_I+)W9)W-Hbf[d/8>1]U+gO.:cJE7;D
a9>_f8P[R;Q_KV9260G(@AeeT4&-[[dSQ2<IgRQ+###T57?#;J1U0,>C2W873/D)
SNYLE#8P0>;ECV<J#L@0XWKeRLFPHS18fNe3-IC=8#/GbLT]<WB]30U^Bf,\/KG;
,-,e+YSDMBOd:#WZ9VH3MJS7C7Ad_0N7);bR2OZX[_(DMeQ)K]W7[;@3FJP,B7&=
D0d6f-S25.TG9M_Y]U.U;6ce?OXF13TY?L5g/C34Q?gG<,M]YR98&F,MgBK4=X&;
9E?ITPcHIH(4,.5T8J9)Q;e3@&84OJ79gGFGU/M?D0&,S30JE]VIe#c.U@F4&W,/
Ia@NF>6+fE<bfSUgaO\MW4AF,E^<KVLJ[a#NTUCMdUZ=]CQ:L6eB&f+++dZK^G:1
B>5T0BAC\W3I87&P_N,/DPC]G0(821(PC9F\?)VEQLgYa:0La_MROC2J,Y0HO.[f
^I6]ZgIG:780.:CH-U&;e1R\=O\-VZ+\YN&/WTdDQB,BV)[2.F.B5<MF0NWT/cDR
=\Yb,8K7JVEX&EDT(ED_ddD<-ZJU-+F\+EaIJ>Z@0d=8&;+5W,-5PM?E6,?;)]c;
CUZZcV[5>)dP=[[T(NC7=15K;>]8S8=Vg36.0-L0[I[TF:aZDDX++NB/<E#\]]g^
EW:1#H\^-eV>R<g><Hc@_FT\.DLN-#AFY)3eBVTc]AVUL,P.]f16#DDKER>XcB4C
FX?fK1)K)I:@a]F15Z@-d8X5K]B75-0TFLZ,V3=)C?Re>OUZ,L#:C9B(1a@SMg/I
1>=fDAQ)V?T2.X1MS[;O+(ZX=9\d8cE4_2gaGe(CMfWDdQV9KTB>6RbMIZYYI<WB
8JM^KGOfT?>J>70#P5X\)V[.B]XDMO@G@&9+DL:SA9425G>PV8d/Q?G/)IJe9dD9
La@^/IG7H<V>2G?UMe:IQMU=P5J[+/J@)L\&EJfO4f-J)CY59]?A6H<O1M)-OUR:
4<A^.&>89cL?C3=:#g-LA(/fM\cM4LDFTBAbT/ZOP>#RCIBg<I#U1<62?1(HZEG.
&Q2;Ab@)KA#NU.+0=KDSNEI>+Kee401VZ04KI)KMg?Yf1dH5)PG>SbNLJ#\,#/D^
BbK@6NS<E?#2P_/-0HM0&c\AHDOIe3g0/_KE1)TVBVVG_S&VRQ3;[O])2_]?J[Ue
MUH1IY+SJKe#f7G<C++6+PQ#J&b1;+#+:(&^J#X/JK?D]BH.bA&07-E3H\a_L&4c
NH5/AIgX@B6f7L=I;<5CJFMK<H6Xb45-WFa4bYZb5-8+OHbKAO(/U=9_(cF7g9:V
a7JaV8\;bEDc?\,FY,dY<^Y6H49M0=cfW?:GQ^@MIRA5>=(#U0ZZT(,)e,IKFA8g
@5AU?ZR)Q9_/6-+?3_1d;ERJ+?4F0WVXJ?7Yg&QaWM#3=/M_dYVP0V5bX0\LaTYa
ONA?a)(ODfJ3dY,9J;bVccQ4,,(2XgA>a^<A\;@W9]_L;3\\7H7FJaAE2W4PDP&Z
WL_GdO+R/MUZP?\Wa)DDe\A/8#d6;H;3:3AT/XN4I@XC;H0H99e[7aa(1Q>?RH=&
/Z4&G+TSYa=Q[44g]T_b[ZbLYEHXT3UK#gC2@fTdW@34UCSgcY7VQAI79W\=&9?Y
\_-U8ALQXbS#^\[_2Y@Og#3UOQSLS04H0HMGeRcN862OXWVd:_I^bW/-e0@ARQ7[
4YP2P+]FVD&:1GUbNe_7D#,#NU-,D\1a&\dE\=3+3MVeD4a&UY_0@dE;T\U>cKW>
b.6+\#c&R2QKV/KY:I]BPIZdR#1G.Be:^E;T7N\3WJQ&1O3(9cE&&.(+/[bTNGGf
ZQ54_Hb0V-2JCgN@e+^IP_<a1cC\IB6U@Kfb0[BL/\bKA2@[[&)7=;P\7V&ZCGZ?
T8L=ga)^-=#JQ=)C8,)\KO)=QH^,/,8&dB@fCa17:^)Y&CQR?g486&_-T0CbcV>Q
L4?GP;_,;/7DgGSF(B@dVIFFc=C,<)T?5.0g3VOP\d;YC<_O)\BY_1THd]=VH.]c
1Y[]9):8<?+YW4R+YR>SU3VEX(O:@3ESOGTDZ\8Be@0Z0@N#Nb]/S/Y_gcA+#XXb
8cPA.=45Ve;,R/(5fHREOI)/0,KBd\KSa?;G1+3@0)L)(93J8/E92&+.M/J+>6Y5
V5YK+6\EXHRZ1BJ5\]]C-US1&#KX(OE@OYZbWA@g6QcdHJY@W_g^(]bfI+[fa\W[
2MY]a=#,WbK?ZYb>:/YK/V&eKML@>,X=^.Dg/_;H5+U&,I]7>@6,_b&/)3&S2S6;
(5;f:[(R_5S4=6)Z9[#L4RYHXaI8KIf[b-))FdXH&@^[13G+;J^ZcUE]d_=:/0F(
5C8GW6dF3f7Z,9_&9@?fJL<]0DL=4NOc?eMNO#\dFG,d=5MPKMA.FBY35e\X4T_G
;]bbOHX2]7@RMUAbHd_d?.^NFAU@&-+D;Md2cR-W8gYFbc)9Q#e03gR,ARC^c-OF
gd7a-=1&ZOF4L37V)eL_?X<1JIA@YMD;U[gPUK0P510[:ISUb:_C3I#Y;Wf,A-6I
SENIP<I9?I33D4@D_V]VOaQX=Z;HbXHD5eLd)RZ34HA7&:?E63C+L3e;&d9A;FaI
_D7=g:2M>FC_e\IDX.\3D]U0\D^,3+<I]c34CPE1S9<XSKZ+P4T-I[IF7>gaO0=&
0QA(e50T[5REW6N#0cXQ_L-\F)F,dJd#@N:5:POcf\8_b^.Hbd,7MT:V\64:gMeU
>@@2S)S:4BS+&e]B8U0-0+HG#abS2;;E&-g8Jg?0DG[M52b>:&19c6SSI=89deJ\
Z,H3^RN6K.+=\@=A\CMJ<Z=g-HIU_2d]288.S@6E]5O9XQ,IXV0UWS<U9;cDg@d_
Q@-eL?:[.SCbO+X2(N?:+g&A=U./5.A:ARB1.6U557\dWKc0\&e;G->D^RU,1_bI
M_AO8-,#U>bN;F3.b[UD_PY.-\@8K-F-HOYX\A9.Kf&1dB9&G=MBd^B6fMCLM_bP
,FdQCXA1Q\cfN\0)A/(D:b-1T.Y>P_.6VH18XNcYB8Z:<fe>);4+K[(b0RTER-E3
ZT]#&X<>B4#Pf?VXKU_7TN2G9c):A9&3Q/W#6[@+?MdK/CfFU]g,QIFZ?KQ5O^X&
GKK;FH5U+E6,AU).81Ld_ZQ/Z]_4dU8MLE+4JST[Q@GKMECG#1+3A^PCM]^^.X_T
F7KFUeT#-@4.>,62bIC&OMcPc&f0OC[Qfg?K5)a.A:3,_H5X(V+c\/XWRcCdN#c+
=V,RbQYW6-HII)R^/aT6[\&WdWbdR\\e;1dLXPE2U8WBC5NUb/^1\>dC0?FQ[(8U
)0JLRU>2c(5d-ZZPGK;-^<QMR-IeWd\C^@7T\.Z215&RL/&YS==(8b/K34<g8(Eb
8?@65ZfI>dH?MC_,-gU<8.5BDbLe@82\&PN=LX5W)DEANL3bKF4_II59;<3SYR6>
L:?P5bW,AN5+T=5)+5.RS7+RRDdY,I]EL=RWE8gb8T>C+fM)A[R/_8:UcUaXSL8_
4cfcT4KNZcS33I?_1R1Y(f.8;J(d5LbdBI3d-8UP=O?f+^f49gO9R/DG3E6RE2?7
]Z+g\1JA#TCE+_X@:gcW:JQ6C+>EPgZEZc+daI26445Og>5Rad3)OEN+LSS?>>K.
BaE:?/HX\&a^8Y?F/1.IF=S\c@SQ6+Ff=AMYRH+T#CF?A&+:BJ[+?^IH]A#dbUN[
6U\X96:YU/-ggO@E3V4U0YF)dMIUa<+Z.d8:Qa?US\\E(^&SYB^EZG],J-Zc(,f7
87JA&=DNA&.6)U#04RA<73L;A[I2(JI:9\SY01@faS.?ET&WFebfECPJ-:V_FK^C
LfWMG;7L.,M2,#^9\\RGd>5CBEaCMT<G]E]MM-AV^T9=X[R2]dE=AC?U?R<9;E<a
&HbVfE)YgZ-#3P6)OH]G2JaK^(bVH-^VO>EO=]EBdQQ]aGH/8\Y/R5A[0U=5@G>^
,((L:OP3g(b4R&>L\M+:HA/<(Vb)Ab-#0DLU.[D>a&R2a6a6P7V8d?E>;2=;Q:AT
R.T+8C#f@GR\HG01821d151M.gT,1=KW<V&+DBed<=6)2ER@/:EF=gC=eKMf1E5b
#Y;2]7\;S>AYVd7Z0:9:Ae.A-b=K:cF\K;_[ZGEJT2KZQ>(a]660>YHQH3J5]>P^
K=aaa?Z,?EH9,c\>+530^ebG@4T_I8+W)\H7.]VT2+>;BfRKd4FV+ZfG>2\/?6YP
d2,CXfPS=W(RT+\88PeCBV5<)J4^&HY\CCI1+B[./BZW,G:cZNTDD_7,OVZB2U)C
9A9E?T?A(FJOLF-Sg)OJ,aQF6^VE\[I:7/-K4ZZ.8,T_IYWK4L[Z?aH_+M=W,ZWM
K6MD?7XWBcIa.3+NT>+d.M@Lf.4B5ENF:\A2,P]UDMaaK+:YXH=fURI=\AGE0EAH
Z9K1-8Q&LOEdLK7J4K-5+a\)Y[b[FIM?<+TYSXPTTd+Z@TUN1PGK3/g43-@OD83N
1UAZBG(GNa26J[B7a8URXcET0E?;4NOQ&3IOQI?0Xa@N8I+4e<240TS+T5-EXU[C
eYU-K1(>J:W,)W[.UC7cU+LMGX=ZK=de^WF?793bc=LQ5/Z(]S868)[1\SDZb>a3
Ne^EPbAgcd)=6a39.&TZUc@.e8Y<.V?=N3d<&YVX^G09/,H]ZTY^VMBFRbU^&#0(
+X).g2SE0K)9[(A07/MFPWNJP4ggf>:1:<.9A\(:S2=V0dZ;8HOf8Kfa9W5QSO\H
B+8D\UKF;ID/1fWa]759ga472P=,f+BN-[HN/2EYRPSIR#7?JJT=U>Cd;CcC:FE<
Z2)bWI/4423[f]gY-J+SO)5P6<^Y5N;-N5^2V#;HNV7\RX21#e4d<^@CSDS=]YVM
-EZHW<cQACWXVJ<]e8HHa:G5Q2X+dD8=7Maf+J:ReDXgL+98d@<=9KG9(.96CI05
NPQW/J[D-cC7T:0e9f2T/)4c[Q[PdTC3JR(Cc\e_@M@WX+ND@]eA=Y?cb=TVJNJ^
gX;II;KGdOJD::^SO9E)36I,(]OFN>Q=VV5_<f(5P3NTg3LbAYP?1AHF69)dH(T\
0\P60#]C)\-6AeMdFe&JD0Tf)CFIX)\Fa2&=0\11OgN#G(@8a58EC4D16b;#dFFQ
1<YPId91O:d>S2CQUBJRM5S7WQ0Q7aFOCH[8Z#W;VGERNc.VJC:RQU?FcYXAUb7@
I(.(\bVYcc2>JINLJL@L6f1F2+Z)ee9T\Jg>;LS8K1JT>5Y0?8NcT[]-/0@6Z9c^
8ZUS<ZC81b_L2E,\V01;#a]6IDG<Q4I)4GgLT0c_1I#>[E960fL:c#2TIg;,_?>M
dNCZ2Dc=[:#.X_^Q^+/N2J-48c.A>8=gf-Z,AU6]<^5cb6Q[6&I7[>2eW^@#.+6Q
6.g8>9;5NE=B@3#S?]J3BVD9L[ZK(Dd=2ObW3/#B,?9-,TWCR093+d[/;=Yg0>gQ
#Y[&d99F72-dIDZX9)OWWCWVJ6J,?Gf^aP3)BGE5==JAE83]_>T_IDPKDTNW1QDH
GIC&aN<Q0;WgN0OZaNT?3HJV0[0<;8>(F^@Y+\6-9:=43FX00>5#;2Wg0Hb5U.&C
:+Ef,[C/UAd&PB;?P#RY)^e][SM&RARGQDH@TFU9Z8cRP.-^cI,N&.R:L0M+e?#S
bb[#Y)7f669^XA,U2]BeAN=@PCG/\7>NeOE<+62.:1HYIX=[HS6cU?OAQ9KZGJH>
/Pb1NN3R9TZ[@)Q^&-8V>Tg+JL;K=2745)V_6VceZK32f(QdBa,27S?OY=OM>V.G
A=.cE[R:Mb6>H3\)RV/-Z7HR/?ERC()OJV,;=I37=-^WE8)5RD>GBf][;P[,B+\_
5>FHY\^bbdgLcS#M[ZHdMcX2a,VF=)@e0fXXe3;_2;#/S)U+RfYa40XPBE,]:58;
bYc>>91(#K6VUZ:PNf)+E;Ye0GQ:[;NN)\&:?a.Z213VGggVQ&HVZYZbF06B0,<I
S>P&Tg)_20-S+VHCf]6.LXf((RGH#U&5eWHCHLYV[VA1\H5(HV3+2J:eOLMB=fHA
>Bb?0Z,b>OB<YAa<b5Q7R(+Z,,P)-^f-^8=?-\JZ>ZKIG6MSJGI7(c(g9Y],T7NV
LRaa=VTLdK#T_XA.<2@_;;S4J0\SB&J>082&JeEMLI98_OJagF[fQ3M[KaQ:K)PH
UH&O@XDQ(_N<D0C#Z9@G\Ue<]]/g05b@^d)e8Lg7H=&@5E\Z<P&V;gCMB9d\Y>A(
@5.&Z4YBZ8[d/I0[Z/L<\KB>7U7=14eEQ-QZ#P_NB4.(C&YbfHN6JGLB);1b-B/-
Z5ON^6S=YI[e^5(U+EfA#SGYY9#+/;5-F_)XJO]9(C+C+HOW).GOY<f3?#T9TYSA
L54:M2SUP+8I;f_PdLM=df_4YZd<YDYM?/<6IfJJNO)/V>5KggeVVPf+&EHL\U@N
>@+BV8C&>c?eHYIZEKc=;,P<H5^#I7):_C6E6>WZbYM(8F7)eY-34bL[QC?V3ASe
cQLXU+9/C:-fUO9Q_2H,aOQXP/.\4;c2.9:=2\3bY9H)e0dfe+BTd1A^)P^PIIFW
)PdJJ6STdBK^/?8SO[5F7_#253LLe#L<4\-E.<WeETgK0,F+e0gJR\_N+d2+IT1f
O1fPTGF3&N+gP?DZgeSe#L+Tc.5F=U/a8(H3WM1-cMEW8O7[T;6]eg<(]V3G=XY0
UK)H(/f^V=2P]X,WP^X@;44afU5N&S>HYO6ZTM[NbFM_O[c&+OO^OBe.1J7A:4]K
FG)3.Mb),.(b?gOA0Y92039f0,,];E@R^bCT5[#b+=@/&IY;gGSXHXHQA0R/<:f-
GWWE/)8)PILVa-3f[@FQ<ID7CW.EKaN?6=K1]HDP/>E4c1,HBFT:FD<S\YFW^M;3
YX:L9YE?H@;<6f]U<WLPE5Y1K+,,1Ha(;A,YJX7-P52acCRCYFI+9SaOOJ_)0\#/
6g;2M9cF01>1.LPb3aX#=/ZgYKfbN,2&:FQH(MUU:YgRFN18Da5\O&f?-EeZ6YOV
+g5SGHQ9M;5[1[O@5?R8/;-Q6g754.f:A24J\,.8)1QVJ)T\R;A-XP(YDP-JgR7g
c&K>]Zg;YXQJ\g1L14\AUU.AZG]R#,YJ0K9_(_9[WAM+/L51d?DUAfO.D[857S)I
Y>S33]SY4P5A+^c)e+[J.R,Q,\=?06PMId,=/fFL:FP7HKEb59Y.,dW3a#ZANF/]
R^9QV.UOKYc@)EdSM2CcfIbaSUdM)\I9CggA^e^3dH<0&BH)DAI;.3W]V9:AALS5
UCU0H0.-+U<DNM120f@G>55Z0BUYDO+TND-IN+0bOU79R5M7Q6WO>LWX@<?8=UVN
<+,W&05g&19ba6,F.cdH1#_IBga_C^D8VC@J=6U\M>U]3XO0J@Z+MQcGOS#UW32,
Ye+.ac^J3?9\.)EdX;IYLXR);T[VETA[_#Q;-.VN4Q8=J;c#1&KZ/D,HZ[d#(5Wf
c1A8J[SH[cCL[GM#A1E=Be\9E@=OF\NH\fF=dTQ+.PdNeM\#cP-Y-+MR73N[F@fF
9dV:,ORFUB)7[P,b>cV66QY0>^-2C4IL.+OeOQg:f,e9c_=c<,6\N@Y7BK7CJ]O_
)Q>Wc3&ZK1B9&g(+RgY?O[]N/C.&YX[Q#OL9g__[WMKdMfEc77.Z[?9F5,d4LQ(b
WL]g?c@Wc^?]cgeg);Y]^.\2XQ8/=e89<RS]fBO(4bf1L3\:fXVRE8fT9>gJYU9g
0/L343ET?bDS;L?T5[P-.-ce1[H[(;5FZV8?>a+JOUH3V(\-=a,?,>8edIP_d-(G
5T=CUG9RcZ2bGL>1ff0Ba1R)SS4e.cJUAdSaH^H^+T,S=W&=BN180-2&Fa?+RHH;
d>OR56YaBVWTG3NSM>;KN1P9H6,GQ4Z<I[[:R=NQ7MfB:PR.,VaN5,Q_KVN+[K7a
T86/eJ8bG6(c/L@69&-82\GCKR6DS)1c_I/Ne&FH16?C,DV8L9I+@F_bVVRIL?^S
O-cB>,E>9F#(<J>0H37N>P>1GJ<MLRW;\WC\IDBHZI<?G_5<-U^(@2(7NYfSdC?F
DOFQK[/,+#XO3Q=#-.^0=aLf12D;JF6TcI[221#B^]B)/F(Y-E^)?LLE>V5bZN0D
B.@<VI_fRHOP/[;e3>3N2.+(R5IWYMSND(AW=J?P0[N+=29QG:RD35K#1Q=_Q?]#
X/-:3<IfB_Dd]=cLFD86?2cL>I6@HYRfKY.\/.(&c<.7CP-gUM<Fd@O54F+?EXO+
JWfcedfQ:+\bB7:^1?5Oe8R4fUZ?f?UHNGG<W>L<f?-MXcR<7c-RSY?eHRB1HEN)
:WW4/931(;K5\#^>K+UTD[_>/[O8gKb-2L?4EE^4B0\-\Z8b<GW2f-#=]>^]GWJD
#-cgI8_EM_RDdbMRWY,U\8Ke0B@<F;R>7a/E>8F7TP3NaL-TG+0g-YY0F4)4]5dQ
OC+Q.Gb0?<(L)Z,eF[2Wg_NIOZL,1-JQBOcOd&T1CH6W=,\AT;C6b;JWdMC2c+-P
K/?bEK5/<&fgF9)SYWO@L@0@C1J:LT2#JWLK8+Ga>;#T0/9UFZ)LF@d^575)5b\)
HUIe_4J>CS=gB;=<<ZGXRdMZ@S&-2RBZ3SBZf>7Y)HB@5)^]]ARbUfOTVVAK=VF.
_II:CGG98X9Wa+5DVMdN7cVJSMf7XI9cQ>5&9d4F):+0WBFGM5])][dY\?V#C&K>
L\^L[T#8OF9f0KJ-.QIf3ZgOK?5L7[G1Sf)N</]WaRdWa/[;YHU=-N>.6BV6,2,3
H<_,&GX:(CSD.2@ZK6HF]TNM0F9PS(9@[?8:TE:[[N;6L>UTAPdMa)-Z,/\aD;SF
/FbZea\W_c-;@^0[=IM)304=c)52P.D=)0Uc<4c1JT@:Cg0/2[?DG4]A@Qg8PSa1
H:Q#>G@G=RPA3ZP[48-g#<&T;<7<L)c+PF62OJfW6L:&)AX##fCL<8=RMT\&-&K6
7dd+33U\#fJ)+E/:];OB)8GKCI4W)Z=d##IRINGNeRRQ5>^+8@N=7O59eX2<(QbO
E1=>PU&=)V;LYH:;LFF,CRXe189@fSe]\T4Y0E9d=bCO.gMGB7E,DI/,CFB>]6_O
3S(F^d^EBVdC_>CC]<+L<7^dZ=C/608(_TP76ZV\<UR6G.@Q;HYA0(#+J<_V2SIU
8AZHCF;4N8#4VHaJ3XJ0QAINAAKY4NT(GP&KW(\G:GUG_,UaP>CF^FE_[cWdGBX\
@g)-;8AOMf?P522)P][6XaFA_.CFa\Y^?VK-N(L_MgBLC6;Q8;ccZQg?>I4C^S:b
6N8[_Ie?#W.@KH2-0]?]Y>GLO?[-a,QR^[S_5W;.eaf68C9/dEE757f.,WD&Z]-4
dId(Q)8eWMd[MA^PQF#60X1&CFM-B/?>2]QSI,3<RgS7UKPXIE)>?JU4V-I9d@Q8
NJ8;P2E1=6N0-8OI+#:<3W+=d?:a]G]TVT]0MA29dWQ-5(B^?)LeOKYGKR..ZId?
TO\27ed8O/,;f6a^ERN;e;G_TeX[[&#/L]:>\1&fg[c4#K]/:f+4[>fTYGN(J7)R
7+<.,H_,<GSF3]L+cEOSI>?,J<N_EK:-NXMOP:C62PBM&eSEbF#?B14;VYKMTCS@
HWZZd(V3,Ve\),_.f\[4a]-R1BRR3:C1V&E?-LQ_Za4:XJ\8YSBH9>2YZW;7<;OP
6GHN;BJ\0cWEN9\N;B9E<dSL8^g95<(1+MR(eJd@O]JKE/MJSXBPaKQ?)00I.Ga0
>BgO,=d33V(6-aOe9a3Q5P3LY57-AgSeY<NZ]+T81JZe6@Z#,ZC832-^af5MY?&^
4T:\SIJDfA9H^5&((dGCV(UYKG./dIbd/LcZF_,;GAadM9)a_5)(/W1H31#G90:c
G#>>L1dd(+;BT-\Y)N7,>B>L@:e(-PZA3#EED\A./PaY3Macg.6Vg],91X.dJ(DR
W9:)^d6c.K4M=R@9DXII6efbM=B4V+P>/]1.M):#d/[CXLQaS+(0H&?SC9ZQXd7E
GH\/+>HI<7++)\-MFSbeR>\ccLXT6/)G?U\QcZVg32=VDQQSH6E5bR#+<Q.VN3Q-
>ID>&c,3W0-/\8>=^g5f.fV@+BbQ9Q3:63B5C7<:T7+36S:;U&[QNQFLgO)>gWBZ
M=XW1RgB6_IZ/c@#A+^.,[Lc4S3[LXdLA0V[46&8KOAMYL:/Zcd;R[HQ,F\1e+^a
H<d:LWU<U2\WFdTCb1(^QWc2@4Re.Z0T?/R&.PB4f[-\g9-:dIK,aBDf+JE&Pf2[
60JUf>eR4NA(026?4/#-JdR7X0E47@1c\IMg<>:MaIB[\/Z6L>Q51ad51B)KcTL=
_^V/A/d)-b8#=@TJ6;QB0CAO>GagFMJO/@BW[#Xa67-L+_)b:L^-+XQ-D:aBH-2c
&:P#T409cQ)f3/RZ^Xeea0g\63.Z\@N\,-YH?T)[c;7-+V?WC/2QTRd50gX;Y8BC
JCDbaNAS?^_->ELH(9,.(.a2XdEF\\_B]DCRZR]U^;.e+4P7VIH4_Je?IU8;e?M=
EbY&LYFGH::SgIKXX?#9:\1)[+>Id_f6[7)E/gMKf-RS+g>K4-g?74)E-bb6LX-(
P,H-R&(2GDIEQD,#GA7).W#S1\<A;G8\-eU.ed1B=4+EN-d&b3P^2[W]+JQ)@[Cg
=bZQL_7R[77>[K3g96HM/Oa.(4@:bW:41>^-_3:M):>dE3_DbX^OG07@D\16BR04
_YfdRN>D1A/>&CG7^E)9J[c(HE0gVLFVV@P]V^2(.JIV&ZX=H32XE,;I5@Cbc/-Z
_K?c2g,?C<e45b69]?gU&;A]/eXO-Qg#f-fcM@YGR]d4YA/?ZUGN/O1TQ:[LGY&B
ZZP:U2^\8D7KEeXg^U.X6]6HH#fTYdEDU)HH&>:)bX)+]G4\,dJYaG]@F82:E>8.
-30f,R5CP^=-Mf+9CTR[+H)4Wc?B&CVa<;QHceK90F#ELATATALRAJ[STb\L7g.M
U3gO:Wf;C>QRNQ96VZ3H<RVH4O4R^5JX-G,N2,?9KHe?a11LECed_^+-dU+L@]=c
bW&Q-UXM:A?_><PQ6RI)cKQA>RXaDEAFQOXZ.AWC0^U?1819feL_5d[R0&a?27,H
:LX)/<_(]e=62ELb?FXdC@abaQ#IZ@@KN9>2V<8-DH?^()=Ta4(gbAbGWT^c-:Z-
8\7WEE7\QW-e67J,V)L_J=&]H-H(6)L.<-\WT5GG4:gS(/75>6IJXWDP33D5238T
==8C9&T5@eH5R::A1\26)/fE^^R?\RXUdIDABCSW]/[g?V[8a./J(;\6,BfRZOP<
):SG^f6@d=8a>2MO.N9]_ISbff:H8G?2JOgC/]@b&8QWWSNX9fR>+CNe(6f>Z+Pg
Mc#9L1##f]Y7geegHW3HY3L^D11G7=c[:c=@E#/GVITd:IN=9HF(=)MV-.=S[P<)
(M8=T4M=QEF:IQ>2WLW@[AeWeH@cHNKD(#eOB-c_3?>W)YD:Z&WNbOWNP>3aY&I5
WUcG\\:([OcU+]9:5AQ?ANM.WB_@1I(=7@8e-V6&Z?#4HYeUe0b>bWNOL^:c-aQ#
GCH0I?AQFQUYY_)2NO^WZa^b3:]N:I65_842ZRH38R#_;aS5P-,af4U@N87@YQ/f
#S(;a1B3cFdecab\a34]Z0HX7;d0/aQ[?EL7X1G_H&JP?HZXM#]-S+9(P,1P4M6K
XS-4L(2geb0a-&8Dc_:Sd_ab5,(8OJ7(31JSd3&8KFB[BS)A35.VaP-K;9WIO?PK
6Z_GY#G&<VD&.M1SBg2?PK/bL?-FZC:H@f:cKMM,f8T7/_Fd3g38BQLX.E.8Y2f-
P3W7gLRd(f0BL5)V(+;R@0^+8,=2Z^MJY;D<.S=\+3_?gbRPCHX3>ZLb;.V&fC8#
2CYCCP?V8G;Ea>Ca:^OI2M:#AL114];fbKA4B7R7A:cAVC2YO#P;VEX)#OOb#;fZ
0\7P@fO<D>YZ/]UKFBMJaHe:G(eJ30-V/;=fP/\6[f^I6d&[#5bF0b]3/1d:_Cg,
Z1TX56b=NUFB)+A05&#=/DR0&00M?C:8RZbaL=0&c,dP?da+=3[=Ic;31G69=N>R
b+8.[((_e#R12_L]X>,GBQb5bA\gA9Xf33e<W^_V=Y>0E5bI\dZP\1)B&DF.a4bA
7d_bbg,BX)2H275#Ebg29cV)^0aIA=AeeCDELF1;Cc)SOTW+D<5CC+XBFUGV^<0G
BC>5E.N\>_Og6J1XcQUI?/J^/I([EJdEfU)[\B3LG^^UT;QW@geAMUF^,MHJd1PO
WN00Se;2;P/OGYTV9&+[4@F&^B.C;b-334C22YFA_Q.+6UX].gaS91PSc5MI77H,
S,U8+6G+Z6cYD=MF0I+9Y1=>9Cd7QUQdA8OdNTVTIK??dM])W3@g_TLT&TYUF^\&
FB2e=3#IgE#-I>2W(BN0GP,:>26ITD,&.D&_Ng-][aK37Ne-5;1,>,A3Z_C+D\)-
]6W4YfO_OA=fg&E-W@@#;CU_c(SMKU:=V8N8QZ[UM5T:42RFJ[-;NAV?<eM@>W0Q
#:=/)(Z.CJe?>2BTBAP2M.LEHb=P)B_25_+gWU[XTQP&GfRd9D1=_-\#1O=28><8
U_T^dERF0a,:H:f9-4X_+ea996:6\df6&:,DYKB)=:(W?\G5.CA:C&f9S+5UA8\f
OI)700,QXF):MSaKZ^\]:XQ4.ObGbUDB@4+>gB&ATQWE?)1DfLLU=[?c.-4\CeK^
5,)LDe>C@_4&53N4bXW:5\FXg833SYR7K<]X[aa>V#&^7<83^BU/c2>3JIA[0Z>N
1C[X27WDWgZa/.;63PF#R>S^FP1J/E@e#ZN4U2L9,/1&aV2Wd@,85UT&RNR>E]4,
baQYY<W6bUS>g#3b6+7=ccIbbbT?K7,NL,(^O;5@aUa/bFCUR+)H\<97OJM?Q#=g
FJ#&e9EC<>QC+MYTRcJHdc&;AZ9F6G]B<^E>EbM>(IYF#=bAX,VQNIAVQULWbYZI
GACOUgT:I)7gO:V>SH?D&G:fO#4[0^V?_dY_&<<R)D&)AE3JObDHcIDNc<?[IZfX
bGL-4FdS@H\SBY8)Tb,CQXIKDL_2OP#)@X27Z9Ka-1gT\I@(WdAWYg8ML4H,C]3D
/O)I&@ME2#RKSKQ_Tb3N9-H,G\@:<\KFV&(0J)[L1N7Qg0LBXTYOa(f\b0U?1O.1
-G:>&&+Vf;O\WeEOgJJG3IUbaALGRO/[a#4_A=&-B:Z6QEb1,&_2&-^\gb\;V3K9
#bWTSE_JXUf<I2fF=g-(]BD5E>V<a_-2HI5CL0WdC5.\>MJ_D3I.eO1_e-,5703g
4A:.(84We@4BC@:I8FJD0+RC?XHKeBf(P6-<I.1)d@_Ve]I_R:Z/eA=9Rf:@B5Oe
eX05)aLI(IYa1T26XWJA>Y-5OS_Z3IF8&gg6]ZW+d0#?7Y#0OM9,fW5>;>+1a6f(
T^7Z)32&B\dCGdGe_?&W(OEB^>a(/e\Lc25_0]\6e[H5aAJ]0=fgYVS#[5,BMJ.:
<a]Z1HbW5OaMJFTY?,70SM1-SESgRQT:^_5e;d35PQ<HZ\<Q9+4g9e]6c\[&e#VT
L?8P>0Yb-,CICJN?(N[#O45)Z).3?-3IU71A?\bM#;C0CKB7NVW8FB8\N&0@/JU[
T0H#X5V^-H_DU4-Y994K___g)Z>MZUL;V#a@FGS#-^.13;2gLYa5QX/Ndd9L1g\P
B4EQGWX(;)PE7N9J/NJb;\G-bITgc<2-.1gK<=.8aEZORVeV(a[2]5g35>L6AA;D
0cAK0=8A.[2S@K[OE@-HTc<G+#]c1,Ve#WNbd_M?.=a8SRBM8L&V:/L8L;C-A-/7
g-+:ZYIW(0CcYSgVPI&-e4K39]<U-08/Oa_B?1UN;4)DeD/G8X/&M6;EeXg)CG^4
CVFP4\a1GIP8#.\;fK6b)0\V2VaNQGa,c<EIE3@A6(EUBWgaKPD=JKTFNO2<[GJ_
Sdc5,6LG?Ee1ZC]><dS8-=PH?@MO8]E\YBeKYPSe[f+[_7C<3d4,f,8XR/:/<9>?
7TSYYZg_O[AKV3V91[.O.6>e.4K]^&LGYOJG()/WZFLM[g6b^?[@()X[@A1>Q0T?
6g,C)Af0.eC&2gYeE.:#DS1a9HD?UH(71:F4;A[Pe.KNE^WT)&W1\g4)bT\IIH93
/]YFT9,:ED(D+]0ecM>SS^O[RN(SK;1^]Z[+=ISKTX;=HT6LgY1A],;ZNNH1cP\<
b(dHc((3EZ)6Y:MOI\4QFV?b#[?F074FTc(A+RU]>F_DC_>T53g,\T9fW;X<.e\&
6B5GO4TVcG\e237Z_#-^9aU0(cN&H2MEP>BD[+D\]AIEO\CQWR1M+@c7BO@IK><K
2Wa8L3I2AW>;F-,=KEDIK-)N&aEW:,RE+GV2@EM:K2KdM9@PG8&U;A,^+WC4H0cX
ZTOA4Y/aD=D_,dF]7/J2H:+b))/Sc8Q:Q.P=GfbZYK44/g<)&Da=Mg)R-HRgNNXM
f+3DfTVMJ6+^ELIgFGPOGP94Q.[gBgSP1I:c_0WFK>WXN[Q2-IFcH4cH9JK5#TI?
/>8XG39,]3H>=2N3Q^Xgd+#]4ReN?I;B_>3U?X?dg;K?&;<11_6LND=TM9A.7;S.
1B+0J\D\QSSC[G9Zc?YY484PF:]++0F^WG:74D[PGOGC?8?M0Ve[ZINa,Cg;M@]3
Nb>YfA.eNF6[6X5S7/JJQQc2:f?QO^,O_,UC7\Y9g;\fLTAV8W8Z&;HDMgHD-9V#
TfW]/3fKZ>9#d2;@&E46c7UR<e.&UODAQ+4/#S[>;a\;3H]H>,5]APb#MZ00YPQ[
ZH\;]MG#HURVP.W)T309\]5.4Kd.BU,c_a99\=a<5;-_dZ_3cQ8e-e7J.=\6[?_b
#+EG>7NBKONG<\QBX_XW9:gW-ERTgUa38:1SgdE;+)3GO#Obg=HL)Lc<U#=.T1+8
e]N\b;^GUC>c0X@[6ab9;\SUPU1VDA@Ea@,F19HZa\K4T0GZ6OHEc\dbHP&d^OQ4
#2(54gK1;#II)IUaPEW)Q/<4);+-#FdX@Dg)dTB2daV)#BV\?ZLA@Y+(\/Y5[ILa
B:Q:W;R/#:>X9:Ud+;Q2D41(fHZ189183FS=XNH^/+[,X)E18ELJ4VVTV,e?geVR
.IY?B^Ag,NWY_D(1HFR6MKI:cc@^?3POf]9)3F.JK<&Y9I4TMNUAJF.O>Na2C2D+
af-SW..C[,CV2SDU\3G;TX@C+J?+PF70C4/5+M(@&Z5>07YBeGR(ObY+F5c;F\g\
e]W1HJ<#FBH2&c@_Vgb=9YG_:Z0<:A#-@f5O((eVBAVc^56V_-X8(;9M63WIX#>J
;1DI]a,bUe@O@b3.(b5R<[SE-872SE,NID.d]cS\?[\[_2NIQ>-P>N)_EPBdc2X>
;\eB#QYF8AgA=FMJ:2T25,<,2gH>ECGFEVCXI8/HN):d6SMSMY@PNcMO7@<OR+B)
O3EFMEK_@c,b#L;GB#KBRB3FNHgb[49E.(;AeD<+T6+RU\V:\]gJMZdYN+S>+bQU
;5f?&T?1E-^(+,1&85e=,&OEf8_&6=fT5PM=8P9f86Fdc<Y,YRbAEIG\;f6#EI^=
8[W/::2c(MaE14-C5Q4(5F9g5S#Ag5b[G]7fZHXLX2G-=R).61C^<2^9b64&ef(6
3Z4ZO2OMg&R=Nec2I2_;a9aYG0V17\c85<8(Kb4fK.7IeDX:ZZ-a83YD?aO>I/F0
07MGNO7,:0^ZTS@YF9@>2f_G[#QIXFQ/0SBD6#aVN)GVQ^7<dY@2IT^Lg#FNNeGQ
DA-@A3LIE@H<9H+a4(G=FMHcX1FKI[&WA(E]GE7T@E0HD6<6]T\#b.2S@P2:\gd:
7X-f,(NXbFN1;Q6dZHb:P1.-,e90X8@gQD6(A<M2?)d;IbK]UHNZ8RYU79dIF&&b
SYUca\05KGB]L^-4VTc-0KB:(IFf,Ke0+2(bXCaZ)H+B.e,a3#bQaS0#AE-SI4/X
?.98gebD/N.)Y&RTC0#8\aXeJfC3IfL#b:I+^EbO+9f<Sb;b>JJQ^]-/cgV:---S
ZM.EA;A:SMFHG:4ZO(Q-K/3?S(6=GDKWF]1@O7W6RcaSI3b9]E<7HL,V:ceLOgR?
G<=DaS3d)2CD\;2JFB?aGLOK7LC,EU4:gV[54)EcH]G0e=QV3:QL&LR23Z#L0e5;
GK+H-7a=WU:XX1QIH<<8RN2-Ie>[(?YFNMOQ8U@()=0LW9OVR87F9dXTG.@(=NeD
Uf=&GFL=(]&1e4-U=<aCSa-JA_MCDeC(D6YA4&dIK_Bg.&7eMGYV:3TO>_K>SJ?T
[aX/d=^;4A<:X)GIJ8\GQM:K)0]41SVcLag@TD/N-UMFPMSa>.)3RL/Ef.[Ia_S\
CH;8ZN8=3,Q,1K2D<JMZ(?ICH;NeG@HVG#&21e40&[-Q814.8W._,^O-4aG[Bf(=
]/fPUZGGLBM9/;b=52W+;:W:2aNcA(@QJ4A[e@O]G-d0EP/X#,:>EXVABC6YWZ;L
]DT=^DI\>\@,f;[TI-cNNM):.N>Ub_<_E-8;9bV=ZK;_6)>MVK&@&aF[_g;A30<5
b+@<e=,R>0>[b+gHAbT2?IQI&AVO2<_KEeaUa5)b6#?9E:3VTb/ALaaO,<[4B1FX
9;0/8-]FMFX41E_/VfR9(debQ<@d3eM_IM/LSJ-H3_H:2G<,]QE6&[MWI,g9,.?8
<?dK3UObO3dZ/(H^/IP^;7YgG=DRC9V/EK=dd+f)Z5^IJ30\TG@_#JFZI4JK5_]<
FK8@O.2cG-=E/U,>8)LPRaG^A1N9B<8V&g12(NWLT<P_C[Z)Ug_^K_V2XKOH+#9#
S=,78@,Y[JE33CZVQWUL=9Q1?CJ&<>eZ)__]&/e/RJVW\C[]ML-W4R9=eX&eV^83
If,P4OUf/--:YEca>#3>E0W,XaNE7/DR:C+A96PL+VHE[Y5&H:(]Y-V#cZR[d-bM
d]f#Y7[7J33b</;?cMJ3fYL#PCC+D0Ie1JE:VD3.F2(B[O44.MGMMEOf&U3K?c1T
5-;C=?fUd5]ZXg)58dXNC^ZXK&+?T2L,OKf\3d&-DB&=FaW6#K=:;VLP^-]B<eJd
Oe\d_&93fO,Z9c99&NF>.9L4)UU[9V45A_eS_bZ):;<F23XF8:9AaUcY(==N=W9[
fce:]V,e^LS\?S4(QB6D_(;&07-Vb=O>dBTYgDS7FAE9+Q0=(@]YXa44XN[>I.D+
faXS<]Fa6>=T/L(bT.[5dFQN)@_)7gPd#Q5eS/HS6Y4.\HW0e-VI:A(X@W1[K[bJ
bU96QG;IK&dHYCYU#J,<#Eg^OVK_@+RFFdW^,YJeEM_V:&Ede3e=W8H712Oe1PJT
d],DHW_Z-(g7?bGM=8dIe7MMK=]=O5aQ[G79Ga&CMPAB,::S9SN@K:NcDLfH@4Eg
3GbP4]0IK)A7=d^\ZE_2^YGSZW2:RTI/RN360&ROXQ<[,-5ASF2C(D:[Y^=F>3G9
R=C=0U;Q\;]aF//;6_8&;f?e>LFdHa>Kcc95ZXe-(8.;JUYDG-(ORUF5DB7<>199
\UVT)(AgH::4dU&BG\#2@g//7#;P@Pb>c@^M>9R[=C]2B)?+7P8I(TXMaZ^:dfR?
#;]:HIRRE=8JV#R6@;3DR@4&F8ZWQ;]L7fEP6>;;bF3D[)8C)g6ZQ9g2IV6PNYRV
E8+3\YeUQ1A/RLV9,V,T/AY9W\0U4[@Pd3HJbH[ZXEUb3#ZRSOBRR,=-cOZFe>[Q
;SG8W]F?\F)-=K]ZUcQ;f+[MP,[.94V.@gNO@QNAc:?T2PH?aR+#RB79O:UCC:3X
#\Ib+1==:X5QCS:DUUM-#/TRc@>:TJ=#<UO=+:IVSW;7gPSOYeY,9/KXY5]FXXH&
6Pf/8N37=X^TJCF4=8BH;Ia,/b-OFb;&RXf??acS=Z:CEU3,bb.YeS)c<75(2bQ<
)fa)R4VeBaOH(SNPQ3C\B59V,P3Tc@<f6<Y:OH1DKK.=e>RCb(?T+@;S=3/<?a-]
B/+2K+:QXH2,5+[AHUNCXOBW:/H(/X4R?[X(2&:f7+R4G&=;bTU[1(E?N4&-6U]J
A4XZ84A:Q#QX(AT\P1].G:4(@^:Y1f3cVNV&<#Xcb\DEF:IJ6-_8H8ZEf/3,T<0e
BCLe0:?MJM\3[,L[#I7SR@G=CZ&]P:6-[GJK5aaZM>J=I6^g5^RVR:.cT<N7-5S9
S:bE17E,<9BJZ,R9.Z]EM.;Rb8L;XX\.CJOUbX0bZ[DJ/YF/B)PD&6<0_7-)SS)4
LE-N]]NHNP^+6]c<f/Uc?2<JI3Y3Ug]5[:,Qa_KX?&YMb-?^<5WDXA&0(+O(F6\H
/caGF/bR<>VVTM6b[ER).J.];WFb?M@IP5/-6A[L=f-/b^LCWNN])U8.-0X6)8Ug
Hc6-DeC1gd9=WP4HJGaEE(XIaAC]CS1BKCGA^8)dY<&U@FWK]f=Jc,5^IXd6_KX6
W:06HgTa;cQWHU#Y4,5g&aJ2f>KO=GgPcN6gEHGDDbIe78Lgfe4:A[T_+3S=#&=S
EG?WLLg73WDA&.e,aK2&JZ]F^>9;L#]1_,_Db_LAI]aNPeFR)&E&903@RU.L2<GS
HM72--<d1T;P(BP9?bN=LZ,EQ/YEEcE[VLIF@;R^O+ZN,d<e>;b>Vg5I4/7LY3[d
/Pg^ObMD+K[Y)@4;C9)bXd<J90c,P;+FW+0+K(UPKA+#D2O_9;(P;F/0^>O&N62&
Vf?HY9dCU^?R\MbT.^M0[a9d,5Z1[(/6/+6Y7NP&e+_@5.<Z]_3ZRJ/Z[.22T(T^
SORCT-1KSKefLOSIda]ZbTMBdNKd[_D9F>HVI^Ge.1fSE^0WE77JK#,;a0(KHQLT
@?.dSf+F/-:PEfWVaHD9MfcNB:1DRTPH(.-)+:3BAfEVP8BH^XVIN>@f^[4#;[1O
Y4Z.\X3@O\PbPE\)TS3\KNV2bJ0eU8Z]40Z2gT(ER9-DcUV)RWc.=AR3/+HS:;N8
8).P)DC5FD8OQ#:E)MXS/a=H8gdHgON&,C\2&#-8OKdD/YHYQ(@0cZ3T9C:/,0V9
&,S)cP6).0DV@-eI[ZaGQ7[6:XbH:/86@T8_>K-2RS4#f2?I?1C4O]/.?@RYc&;E
B))=<4TTFRSE^U^UK+4Q?.-LP7&X+5Cf(W&/dd()\e)<^LS\gQZ/3L2FR2J]NMf]
ZRFYdgY3+O^@>gLZ7g;W)fQ54HZP@C8TC6CHJ=HQ)2JAdOQS65)VMc(9,[#S]WcG
<J=9B>VA2C?75_NN<&>5#FRB(C;X2Le#36/<NbE+[aI^:M7+Yg>S#&7__81e3JVd
7cG?UX2XG-?F^-?^.;(B_^?L-H&J&EI4Y5[=;B217&UP42?9fc.P:?8e98eO,E^&
@\37Q6L0DOKI;\3d>01/ISN/)20/P7[UC]XB]8O-QYb2&gMS-9TA.5(L+1/WS-G5
[a=7Y?3++e#3N^ZYHO7gF-#8W,33&(1>8;2?H#@F6H.O/QN1^UVOFDW>G?9fe>G:
0PK/:I)P@U:aMBI;#<,5ECg)O8@BU6K2X3_G,POJ,IHR(DEdLHSZgDcUBIg2:TU?
U+dI<d?3O@YR&AfeQdeg&=Y/T+E/:6VdaY(<IbZM<\N3?Pb)?4&Z(M6H/aOc_8?_
;0@RgN4)ab;XLX&)f6]?T#gN]&J3]GK[YCH\4;#(?L/UM0^9HfPVGS5ceF]P:&0]
5>5f?T@,\2\c=6SEg<L]cca=:JERYM0Kca;R/2&#_<_.DHK6+BGb+bNUWN)\[?&;
U,KBCB=3M.3.OgbK55K;AC(/KI4_9da5RcT<e_3/6].#b5LKN861.3GKO^_f#:H^
]L7G^Y7[#/.3GL&J7&=-e#<JQBIAc\[&eCa=I>gU8QZaMETNN^.M^G[.@^U;5+J6
/]1bgHZ,F#J_:].6-]\[N[4\8#^EC:4>PGNA5P]#W8a+@VMT2,9?@c</3d6LcYB#
#(gR/OM#EB_UR;0/e;B?/;U-B(?dE1C165Z/T\A<;I5gaV44Y@ca-7,QA_OTAHHT
KG0@/OOJV6<<[UTHbNZa+7e:I3(gWFMAXXWRb2gNVGA@SQ,^GE=S.6=Q6F@_3(XB
eG]@4-DBUHOO@<@7#U3U9E[;(=)^IdCZ09MJ[#:a?bASC?J5<B0?c[Zd[]S-MOe3
EN6]SaSYeLS730c=H1L+^TU],SZR:&[:2f)dD#LJ8J>Qg>^=><GC:^HK^d&dH6=[
59HZ5<;9(+SY=B(cW8\<B#OG+,5fQ+\;?7;4CV8/2F>\X+Ub7UN0#N@,PeCZ[(gb
A8</DTM.ZdIId&HKT&\[0OV-;,O]EKLPM3W/^,@B=D?U9]\Se#^L7E>K^;/H3GEW
,CH[d?CJ+MZ1V945)8#BVC3=?X.=:GQDfY(+L-06A>C&1^2H7P^7+0A71\TYH0f1
[<QRc#X&2gQQ_Iec\/LCYdCH?+HV)-(/ADZ^f/D7@,YXSA@,(430JaN7UF1KZ9XL
@@0bd5bMD,V^0>Le.Z>@X)1f>g)S1Tb+Q/XRCG+@(:#a5Pa#(W/,<>?g]@&/99<a
)H]H6Y-#1:\<[_b.fc[^G2a:cR6XA,1cPYe94/JaL(CEV@-:fRUa6D.7d6JH2J:Z
]\dG82DRc[,dZE];fg(E<V1)1c\e\CJ9/Fg&)Gf\XNZ6XgB2DV]=^9<(@@=Q8QPP
Y#EH;8:SNF:72D4CA(WBb8Q>MW]ZR&&R(IM#1#YU(c#4fC)^TV#W=W5g^?g;XBQe
K^(E])1?66-XY>^,93Lg&bUKO0REPXY+<:B34/?FZ]=gATN#gfHQ3\N5,A98HTZN
/J9)=DO=aXLa2_LPHc.8_KHfL[MXB].6.PD7M5:??K14:VM?TXGV.5RE@K0fT<2\
2C#^(dTU8RL.aZ+2;T)^\gYa2,[CH=QJII;_#HI7_0D38aT,#_U^JZ43NL2>@.RV
\R<_#,2f6F#3=2^;f7ZTBZSdA]LQ/755)NF[0WY@9\FOAaBfJFG1&E]Qb3:73c?E
C7QY^F[V@8NZ]1f#.dR8;\WC.@5/Z+;>?8&V2ZGa]9B43Q+\GDf3872Z_J-_Q&Dc
3&g5b6G:[NSY)bSPB@.=Q-LG7a6?OR\<+4?gZ&D&R]DF\bQ/8aT8\=M[LQ[MgX^?
<BLY_L&f@I#)e#M8T>KW+/KgG[7]I7-&&LZcDD5@Z)GASGK;BWPb.]]?0.FG9#1<
5B;KJ[;-6[(;U_+1->((:[XbXe54YDLZR,P24Bf4/>;36A+ae>PTL?HELg.WK,ZE
]<&68=S8R>&M)9cBOY=7CLJ@_#1KQ8R3[M<.;eM8ZZND2Z)NC=BG[@eQ2If?ZHMN
X_1LP7G__5D7IAJd_0N<A3=,[4E.Pd#.HGC;2X@PE:>b-VWB,_S(0P]4CR.+IDQ\
,gHTgD6[f=feabI+eATDF?#137>ae,30<=+AWKPS6Ff8,Q2UeDJA8?bP7JJT<#FB
f[e0g]R?/;HE.[)GE+c;R/NF=Gd3e0VEG05UK268(:9;[3fb)4@]Q)9KSa=V)?3P
IP^TDPVQ?@A60OcVR&]gO,?(8=)WB5QXGY=O>B\.34+3[30#0K,(bGgTFe[3Me>0
aSXe:?:9BI?PX.Mb(3?c&XJOL]MeSN.;e2@e7D_4-#PNB001X9=#PIA1_>5GWTVK
H,MU@U-.K.H/Y/-ADJSKc6HS0@WDDO)[:TGDR(XD;/=:S29aUW^M&..V95(@:OZH
PdK+=X:JeFd8ff#P4.M#EAG8>HC6&)J\,CY)-#ID:<A6NL_:^;(/.+R_eYc[<CBG
)MP)/-K[EZV7KV+7[)-g@A9^e-_]&]OU?(&AUT:IG3g6(^;OW47I7SHV#ZDg3\IW
#g;3b,+dbI)+P^6]L/Z5=f\6(M1NHA1]U;+=/02L)@M_,d@P@fFJ;?eYVZ_/NR0>
[c.g:MDI&I0Y/U>(T4U[CR/0^A#,B^I-N9g&#GY1RM09Ta(=3,?P]\HGa5e2^>#@
#V&N7?JN.c5U:9X-5)289;\DH5@S\)f[PH>Ieb[ITGM^?\WI]<:OT6e3FIE7-T,>
RgM-C>634&=YgJ+9EBfdB/AbY&5SF.N:+E?MfJbY4DgU-#dVFTQDI(L7[GPX9eT,
(b]QX810.P28?#VeP-<7OV\SV=b77G.8=d@6U9Z>FBN9,(_[IPF+0-3Nf>KF;\A-
P_=E]9K+B\<A;O6gWR+X1>IgP>4HH1de)Id_<2f^5S[#>O?/+HbM>=#0daJ@EJYV
X#1B^]52YW;OI=)Oc^cJB82\_AE95SLP8fV,de;5@ES9AS-L>YdM8RBLT/6W@,<)
Q+BE\5?9AE=#08fER(Y\a>8FC&/\>UK9S?X=>#eS;AcT\JOSfa.K?1<M)H]Z#,HA
NK13K\?(I9WC36I\MfL>8<WMA2,M\JT6c=Dd:YbXK.S&g?/C&V/T]./ef3E7dE<a
FH#KdBGE#>K;2)C),&X6=CcfLa)@3b=e-K4#BD@R#/A.H]Wg:+I;ObGGE(#<-9BV
8+PU(NO,6?GMQEWSZ#]+[EMYc8@X8X&ZLg110-a:8JI4Q4X^JS1QZ+A0eJA[,J1V
XAOXGY=^HEVIRSCeKD5,]JOUeN3#D-QT47/C5JD38,gC8Z,<+A8S\D<ACVfU&G_c
HCX&R(<RVd)^_Ef>K(WcV#+)IQe\bL52e8@;O>=)]5V[DGEd6WB8>.U#V&W+T)I]
dQ\##1M1)XPX_-^dU1UaW:\cT+/VNb75AO]f<K>O64Ad4Wa6&?DQ6J3L=DLW_&WS
b[45=YR.ac8R=>=C#YG^]4AGFCR+gOCU4^M0H>)DQ1<bUE#2\(HP#c<B,E#(G884
\aALQH]gTS8)S\12g]:dU77R#QX#6fQR@JIZ3_:Fa1?S5bKN?b5Y7AA:#&VEC+a9
5b^KMM72OLaSWN-X\@RWKKNJ^BE)@)W[g7U#DF/U]a?I)Z4XN4D.=T1[A@AJ2(Z4
J<=;+I-7Fc)^AA0Z&1M/f1Z?f>e]:_1I7SJZUUQ^AT8cBgff-3TC.K;?XG.U-I.>
V)gUI.]DE+V[M[C@;NaY<f=Z+,/>2da/;+UX?RUBGdFU@?gL):WcQ@WCd-(MaF6.
S>VfDLf)#KN\.UO:1;?WV;8R0_I67U^5Y?^f_F#5XY(^.ScTHP_\&9D(8^RaM[9(
9XdUI]&E=VMDAQIMW679>]HZ+PTOM,LQ]G=_)\f7e@4[cXC?,.K.J@W#CM,68aPE
-W:OgG76a-CWP@K&4CT<S(_5-,29@UA@LD;(HOBf^?e[NJHcGUBI@EdSB-.<YES>
Vbgg006FUQ0#O1\<KAY166K2Rd1S]ScVLIV<,N#]W:B4@AH?#4L1\Z\O)]H5O42K
Oa.L]Y0)S[:([WD4c#WQ=;3#+.eDb]^)W]9HJ@D_-O&Fa?gebS[6>JX#Z_+_SAXZ
F?N1>T:01YYYcVY(M-V.8W.:2FcF,[.T(;/=H?G3CP410@24>L8<195d^[YB01SN
]g8g64>\8>:U=5)8G[K^H9LO90M_)5bK7XgL8WAeQ,YZ<#ecNcMZ^#@OMR]33M,[
Z6)&@A=#fN9fM[4D8#+:-Pc(1Z,&LQ_GEWKNgT/T^#TVS[K:2#8.&L\_(#?K=-KU
6[L4(^DC/1S\L-X-<e#J\&NdURT-2SN/)dKXNOO,ELaT/-)IB4)>H_X7ec=-?]c&
@4.Re3T[+)].1&]\1ZEWL;(YGZ2Xa91J-4<\M,A4ZEbU:-BE2:d;Wb6YBUa#5&=g
e:D\4?K>U-(g6C,Z7U2fQb@0DOFd]ZLg,(f.I.8X7]=#J(XTc@1MCZ@1ZgaJeSIa
DV[/@#TFZf8[G^IbSHTKLaZ5Ya&&()5?ID7dGXIU[ATfA^^#-S#/<[7GMEPO7c&Z
5e=XXG>aeC0(S4@=&bQZAaaP/]1.8,71GDJ3Ud+6XH?U21M>D)7B?8eS<HG)L3M1
:C=VUCKX7X&Q:aMBQb3-c17g;@0&NL#C;SM&;W-4/0UJfDLcbMI5R>UP?XO8+8BR
?Y7fD>7Se=8cCXZ?\+f38C>:SK=Y_HHDM^aJ)V@WKUY\XQIOA[3(,EeX@CbDA9[>
([Z[6WH(2K;;G_GcKY1F-&be0Z^,IO@#4f=PO\?eVP,.^Cb.\CQ]MHDB4UV/F7FU
D]:_Ga.RCff+814HU)K,g9,:XYD.Y^W^ZB3V<?(29MHHcD]4OH[CfW5Ab)^<12;B
4d8cA0R:#3..NSM,0S\dLW^#AAPP.&&-DP2J7.aef1KKa2;5([c4b0;>Va75HB0#
,(_XWP5/b=MggFf6d4NeS[]7FSH#36Gb3PN,?HdAM[M8R>1\^CZM#C[e2;LOgMZa
(4.@S4\(XJF35B>J(F8L0S7N@NS2E=#.[\8a5N298A[P^EHX9\FWCSAdZFRdadW7
6N;TW?,/[_]Z_2MX^B<G;#Kbf3C=USE,(1SH>9_1RZe<>#AaYXCFZD];)e^aJB<J
#EC3>R+H<V/1\SI1d#0Je0Q8)<#5K=JgJ(LWK3(Y+-8H3O.&T4HDc>)gZ_J3a/2C
JWXAcCaI+eE=#^@T\e,S2SZWY#8PF@;^dQQDOd@cL_;HLV3E-a,2d?BK97-<?>N@
H2M#L)/]Na:EU-E9AV6eb38..=+Q#-\a=f5P((Tc=8[)\M&M(JZcOJ4TW&UJ:1HA
C+C[W;5F^WN0a12IQRNQD]?G(RVF]1,X29g:YS[]\&@><ab40KM]/1;<>+H+2E&A
YN)\gG5T#DN86,>_I6,/7,4SNC=((Fe?C\GZ5)GZ)0MeOSW7b?A=E6X>WF?D#2Y@
1Q4MdHFU(>Ib6LE(V,gIdWa\abE=?aU-+58Z<6^#Z?\d@TM&EY,>[B#YQ^Q?S#2a
ZGEKEB@J(P0+M6^YCF\D2XTVSH+:>I45ZB/bB+6&=3U8<,7ab[EH@?V@&]FNagED
@LYE)8M]D4K#EV#>NE;22:H_/5XRPPe&GDU?BJW9W3^c:6?H:34?VY&<eA+bCG>>
-bHGW60-\RG.-9a)V)1E414a:JP+QaV5MDMJ\23I#_U2S)3@]?)DPC;d,M;#F9aT
da=E8WO.TCFcFe?>8<9HJ#e6IT=LOC63S)R/=T57&-dbbN)M^)4I4A+[Ge=G;EP+
++Ab3L(9BIg2V0G+[bg/Me8^(6[5#-7M4.;8C=f(+)QbH@B?+/UQX9TISNTV,BTR
?FA^ET;Ob9@CWf5:(6=<-6;Ue7B>GT;?:+8=GJW=27&[&Z,Y81[GPF>HaQNET1X6
aP]-,(.^Z>]V?a5gR9QSQ\/V#(7ARAEdea;d?/TSS2.D7f4,-#LNTXH)OAG?\VL[
g<[W;_d)WA[He;6-NB3d65TR+N7Y.R6KadTI+MRQcM&:QGB1cMg[YPU.R#AXC:4Q
T-)9ODTTR)3&U(8/=g_W3,R9C5c[5IOQG:E((VBV_G:7N8@/^YA](PRD7e1]NW0(
8.W;^5\,03Ba-:&U/PVRQO40FWF?=fcOfH7N[6Z_&ZQP4N]?^b=71Y>??BTLJV\g
5EW.H1+(6;H]>gE>]?fSO&a9#(ET7/Vb4C_U_TI8S/K]VRZ?X/=GR]8fK_0A3ASF
d>U_e&EV#4D(Vgb/RQb4H5MAU(TRbMX7P:J_80T+SdK&N2#=@6.bbL&66.SbZ[56
DVZ@,B=?Agg+H.>8C>SJX:;2H4F^1&21U(0a;T)g5?eK[JMTfBS()/[K6&;_,bgA
UQSgQ_)fDLVaO\c9^U#2_6::#-a50G(M6/D[4U<T(c(S^JV^Q>Mf&Qc3J&,0[/;:
.#00b+?AOZB2BLS\T2J74^MDNeA:^4:+)#_>OJ;a6FOdE#9]LU6QJ&EMV7T#I[de
Da9Fg6>;[,Y\N3Bd[I1GK3_W5eMc<TMIYV;H:L4e-M,<+UP-->1<:\7ID=TQfSCR
DgPOH@05</\LM#DL,^BgP<BLQ/cFF\6J::>+IMcUFRKFYU0gQQ59,;6O>I[\e0>X
3FU+\6EH.YJN?IW<>f>5XYN>I_eMH=g=A-c^_5NZ&,_aY2RcCFVR8@@KZGW/KXC=
RR/<;MNaY<4/],_../[+GVY[aHOdZfXA(b83:cU3MTMIaMgO)OcQI])F9]/ZeL33
B8-a-FV.&[;@4>RV<9B&,FMP[KQ07P_J#D.9#DC:N@[)V<.P;;fJA6f0^UEA45ba
N^Z+g;I)gPKM<:=40Dc(DKd4KfT115K^QST0)I9?&43.Z^=989ZGW#DVX0/_ZSG/
HM;eX\]Wb[0JgCP7f1)c;HZ(aaW9K->]Za>\F6H[N[[;+040]eVT;5Q3=f;a;9-/
M#AaaL,IUcJW7TTIS\P#HSc-c.WHe&<Nb2<4gDgOUY,+Y_bJELL97bT]-+J3<U7c
O+feJdO&56-\E2g?@A))ZV_cCWU^753H@bV08<BM)VfH<CB)ICG_(H<:-5.O),PL
^/@S&]U@UC-@fFO14G011L?D<gQOf<92J/QO#?,(X?9KWC6NbO2e5f_1aX4J8Lc?
]MgF:T#d\_^5+a]U^E-PA?edV:Og4Q]EDZ;Ie@MH:HX8FGJg<d<AT:[>M.5\c?X/
UN;AKb5aB<Y_-O:U3B85JDQ9OfF=Q8HTe<\K<JdD)fD=Z8PfX\\,<bZ(THM_3cOJ
CTFI8#EG7eb/76a0Q-EDEC9TW0]4K<I++5V98Q+La20>\AA9/AW.g;X;.UMF[S8Z
/]KO1L8-f/BB&ME9)dX4NE0(.Qd9?ABHT3J]K56/WDTgBHPc6I.Lf6TQ/]9=g=+)
MN<8.NaE(0&6<SEHEUL]ESJ;_T):a<]>.S^J9.TG04=TJ.>aM2SBRNK.c2eA88QR
3B5GPFO#SJ^E_4I@/fCXQdfd]YWV9OfIKcONgfS^fRLGNaBgQH1M<TVefE6IfRdQ
B#A20+dXLN=S9&+;BM8Nb(VZ,gJ0K05-SQ,SYPdW?Pc8K.+#;3(/,:4]T[3e3>0f
:&2+7Z4Z0d<TM,4DJMFV0GTQLgX-/fI<(;e8[7]Kc3WWLP^cQ^JT(^R9:^/]DDGb
:FE7A.6cS6g]26-,C4XKd^W=YU0J6bMRKe.:ec?BXK)F^O6D4?:4.)2IHI62O,3.
EF_MQG[F(9M7-3EMO2J]4<b[)ND:Yf6-JEZG9W<2W;;Q5KB6;_Ab(E9,Y3DYU47?
QgNgd(#gD8YLR]P;#[M^daBO.eWHg]ZaX&OL9<A&f<eAT&EG[Uf8>6aI6-ffYK/,
JOE=B7CfK#PKBJ_,-5Oa]51?.DA#,XV3A=V),BW#@F#_>9<_WGMFQRWdd(\=^/H=
3QS@e=TYf&K@dCH@C/aCX#)bAUfTK]ZG?_&+I+CA5=XY^>?9WReU7f&89#4R:B](
T]bK<J@U^(71^HX(OURX@L.L5cO:cM8,S65>Pb^T8cCc-S<K:BOX9H<P&>XYW@OA
1a21/=XaJFb@F[/>Yfe+22S1G=HZaF8BP.EOd5;),,TLc+)D1:@[+Ef)TN5K[A1;
a8DDA#g^[UOe0?:FQd2[P)#d>DPYCcFa&=QZ/DRFBS&4R&&W31+V?A.J(Q?UQ+RJ
ELQS:B>EG\?F,Bf6GE:RW(:-#V:O?YQOeG[<)&/U,\?f&Fb\@7^(6.G8cg?VaRYF
=+7SM=:X-d8?F&2+-[>J9KB.aJfZKB&QVc:K;K8SHHV-^bd@6eef;Q&HUI1N4SK3
/7U.17cfIcc@K_gJ7YE]N:G9g3?7XgFfK4eI8JPJ>?DF/Z6:8e3X1T@T(gDKDF\/
YPa?S\2F&B\R]YT8M7JWNHRA;SS8\@4=C4V^DNMHfTWe9LZ4I5-G?A/YVbbAH7[\
YA;_K[+84Q>NEJ1gS0X/(>/GP?0Q.^6bO4C3N,0QM]A#W@6Ng#O_/e+^Z,2X0a=C
.)9FD[(c.bXRT;BA.?MWE5E=AY++6Of-@34;R4_QS##<VCcf(^9DU8G<M#6^0PdI
@Te8a[3GVIa\NCPDK=XEQIW7<82DU6F3[T(>>c\@WCg>FfZLa>)F#\<6?g(dEb?7
J&(^TT>RAK^W-Q=fHJQAW>.(7e8S(e_=3_SgOA=HfBdZ,>@&RA\2U>:.,\8OH:#S
@=DW9QY=+AMOaCQ<7Qb.fUUgXP,-gA49^S0g[L(ZEQ_KdI@Vf)18D;>f>cVAKNGY
LOK+ReR_BKTf8DHRCPe#;VK&C+f1&1[dg?+I5OU#X+8#_@]UXCW?XfJ8&L4ZcM.4
45E5WVcG8327#(aO]@5M6gMRWd&-F_ESI4,)#;e]\cb__K.6A@WS-\0g=YY^a)T0
/5E4NP2]/EM-T>d/,>L=16[-g[g\@YCc[6D+7d9P\+X,Z2&:<?)O2@YOd3R/G?<&
0.PL(/^PCM\[]<:\1J.S#Kf,W7JcTa:T\KC>:CN;5TS/E6cW97N8FN@A94<0b8DN
+D]A<G#G2SE-CXA03)@?;L7H]dHC/0=3bBERJ55L>e0ZZ5C:<[d4#AVCB?BF^_SM
ZOD?SR\BH>AW,R#HJe#IF8?e,B&,1fNMBJ>,Lc(1NOV_<H.cL(;G0:1\aUba,.#.
VUB+Z<LD7Q:/U<:^bPBQOHS[;4W=A(a/d,T8+]@;V0&7&ZA.BD^d_:ZGBaffHC5_
90N52S9G(^PRZ,3MA5VC6aNR:[+[a>RJ+L#_FA+I65+L^F4I4E4T8aNGN+QDOP=I
f^-3BWE7^Q6Hd4=BdT@R#<RcC5UbOC@]G409c?Z&8[fcX^7.afV];b<B/;B/?a;g
9WNLXQcZ>gMOf:KcHUD1,_6F6F^@JL&SCJQHKWI,^RLX2/<P24g6YcN6_+OTfYY1
9<c,gNYY;f5V[Q8\?6A1Ze0,EL-,,C5PLUcGX)@PI>N=0a,D\Z7J-<,:aSS_S:)D
E:F\<W/3RK5dA]HU\Q->M:-H_-58ZBCd<a\0bWLb1dcPI>a)X>4/QcG]@)>I]U,#
DI?2TP(e:F:ZEDBD,H=W(9IWJ,1R9[)R^;S()(_-QQbG/#IR)44dP&02^D)2UZ&K
+60R#6XE)/U.g+_>F9dVEV2_K.ZaW16\_9]\)_M8PN29eI:\PO.9IM1a@bbRSZ?O
2LQ5KD)),;D[:-HSE4:_EZO^.I:/#1=3\I+:eJ+GgV.&Agf&MU[NHYdTM)R[J.(6
EMgA>V7I=7OPJc<=D4cf<[I/<[7-:JCeE>J75JgfI>M[7=Na#6IP=1Za4/eGaJCf
Z)IY:6SM9b2g<4d4)G^0905=R-b\-2>W1.bWXEF3RR4PU/)3cHTJDN&.Va-U^+T-
;Y.1C6(O2&N&1Q>Z/aM9cY>]B<DE=U5df3SP/TV51dA]0Z6;N58IL^F^Y6:##.HQ
;dMZ7G/eTA_>\_=a]aK8_.N\Ec6E))K4QSM9>86R>1U)\)D&>73Y73277J6IFE5>
Nf#C\fB/U+aGRGDC?K-ga8D=,<[U>#WGcg,VWW)e<,N\A.9UT<PPDJIQb8VJUNC&
5eG:Vd]K-.,L5a><._KAZU?X8(bN&cX2QJbb].9P)#<ODM3+[CO:G,/.1AfI]e/\
\aWWgQ;:7aS2e=H[U#HT\:WE/-Qc<EaAMI(CS6].^CUP&1\9Y.F/V085S@H.ffd9
N.W\SAO46R^?1MS?8.K;bH7/46G,K1bWJ9N#K1f-6<JRLf0:?3EB(L1EY+-#.GUN
M7dF>[G7^0<3^9b8]:GP2(65MIGc^Pd0S)a[>LSEf^0H>[O,BXd_.4\Pa7=X;PFH
.3Z[Z83)4FKQNeQA>-<L@@3GgXFGI&MZ(;#Q+ITK:FcJTaIS)Z6,I1ZT+MC#VY,@
aXbAM-QHLKTUeB[H>NWgPc+TQI]6)cB0]2[N6N,VBT:95^I)\C^,]c#8Na12[3-E
>2W>6@A&0+A1W.GX5QcbXT=W/AFQg?T0SE8J#A:LW@af<JK&La/Z&3[N\cT(LYDE
5e8N88\/H6N]Y9:B:4GYD7F<G=eDYc)gV8E4(@@1CR5&W+43(H<T<#2]V0#b[PC,
BZ7AZGLW5E@e=44YW0a3.>-^6YdHKICL0(DE(5JW@&eC:-7e8Y-561VR^SN6W5IU
MK,3e#^JMN//FTfdKcZ@@=--;9KM5P2+L@\YSV/C3(@4&6fMKV.Z<BLc@Mg3L-)F
-DR2D9T<g-H[H-ZC2f[&&5E.=ZZ?-\gI03+?g?5?4R\fVR;;DdX11(.<\<f_bDQL
RG\#E(6V[OQI5(R,)bQ5,WS?@G9.YH7a_@3=ffd^^WR?3DB7c>B#acQB:<Q5BfO8
Qa#-->K[JE,.:SMgZN[KN@(>/E<CdT/Y5^H#>79_>NNRW<.D7L=g(P10G4?5PE/F
2S:B0R/IHS\&[bX)/9/@\:LD3@:Hd)B\CV]Z)b1J8XQYL,f7[d;(/Y?Y)TVQg);9
YF_DI4f5Q\D>^gVfg&9:)TU(2/3gfU5X5UR,#(-RTf^DJ#ZH?I5)OX>QCNY[9QcU
\&CKJbcOY92[9AKDUEL_)J4IU#^RX2RCdS-:H3b1>G:KU[+I&OUTM<GTVL&geVOR
?>ZM]3->e?T;>:NK=VZ2O+H8J7^_EccFfRDNgeK@B1,BDPaF2]&]6RbM=#T^/GBN
4TC.DZc.=PA8#8WV+M#3[7&WKTU8^fE&F)1bXRPP;c4D5,U8>KCVE]Tg=W8Rd0Y?
(63)#\/W<@3(#^.GJPeQ;P9L=1RS&VNV_#D.<T3P&c8&<f>Z9&\WEB8\014BMc(?
>KV/^BeW&A1Z??V03e[[;-\E>DZ?DD=#,S&f[AKG<PL_P&f6Gd<WEG9[&WR6JM<V
JF,4\a154Xf_9A\?YQbTCOA0_,NE^76Q-/_5IR,+Q_KaKK].-eEDadM>.V4DFF[9
G@1P4&R-VfHQgQ52:0C>[SU=UDXg?>B;_.-L6EWeA_GP\?D3gL24TXHAFdGYaT-M
&Z8B7>A49T8:09I/cGd:7A+LGE@&:_C7dB+F[ZY347]aW,V2[03O=U=HJRKTZ0(-
\G.B,LK5AUA0.G9B>A3#1-fBQ;.>U)Y(fUAJ[O[GF]eb#ag3S[2H+NI-dggbd\C?
2?cRcfV;.U1(2[g1>fMBB2HFf/P;GE&14\?Ldeada[O\3+Z4_,W>&gB1NBT<c#f+
18?&E&g@^QAXLMSYL^IM>J/GQ<L,O]D2NZ^AZ,X0>##7aYG[8e#V/?-++eQQR48c
UF5:,U)C?<A.V4PR;.cR_KPRLbEZ@=4b)=1.+EMFTPMEHR.;<.LKXF)/c=>KO\F&
C0BS6JG@?4-1>XQ:QFbM)1V/)ZL(f5eSaA5-VPIc^b<7cV2UQ_HEKS8g,.,;VTF#
+1A8I?](=MW0)\2IP.JU)(,>GH-02ANTXFYaTcT^/=g>;&=&,EF_]HCc04a.07[@
ALBX.2(>>>]gJ4\_LM9/D>>XOS9fK8O526A8AMWC\#LN(ZRJ[-2^<b,#D>;:R5)B
A-:8._O99;<H\TC2[HCX#2EaWN(RIWbEFP:5dO96>]La>9EAcYf/XBQ=?BB+<9<)
D9c1Ob-8OL^>&9F>6=N<Q)R;U&-2K>CAT6\<C=N0R;W29Y:ZgMU?S2.W&Ydg\<Z@
;;UZLRM@7c[3.7MI=&QcF^P10Rb8^)J-45TeabK^+I7(EBRK=_/gM:U=[g6CILXO
?#@S0:(AgbBZ2,GXUeM10H\/U8b5P:3KON7b,1AV72Cd<eHMCT4ZKP&]_&9LC5.H
=UWS(Fa;EQL,<9N2_XeWQ])<R&QK-OYc9;b;9C:50>_,#406K;VXTG:A>_CK]R9G
eX]-./KIX5<U[W&6IS4U1GdYaf?PV&F.e,K(VYJ2)2-VcRT_-^PW>\ZDGK;;ce_,
A7f,]_eNBM7[eCdOA@KFM4a8gE6S3,dMEJRV1O;g?J:Ia0,)#-dBN<7a<E0.2RK(
BGdE(I?cWST&C+3,.JZ>4fd_J8;20e1C-PKP9_eO,HGTH?J@(T;2&\2D@DZ[F4N@
-UUI?^f,#-d\FQ97:[)cH<:,T3e-@?+:/BOK23RYQ-=E(WN3HJ&PGXDe.S>=K+dg
L=S?#&[e:OZV1H[4ZQEE]ePJE5\JAg:M<:36,e-I/OfVW<<NCbD6]UX2[9[?G=9?
^eYAPPP#JH9D61B5d1T;SG>:);R:F@Ed&H4.EF.JA)S2SBQ1Q4H==+^Q&eM:(&#[
(1c1-dD,@J&2_6JdIXEIJ<H_D(OF.,Be7AM]_Y-B0-9\19,J7J>c)_?OK@-ZAN5T
R-/Z(a;9B^1ba]5Jg/^SJ@0fA+9V.IO/,X^CM;2WR&4Offf]Hec]17Pa@L;FW=+P
#aW&aW+&4dU8AQ(9-c?JaT8?:-9;WC7>N37:?JG0(,7M@K?Z+8+ZeJ;M?3:;UQS_
I;#@5;-9b,OTb3;TB;)J_2?9Td9>)PT&fe3FPTAeB]ggW@JK8KDPbdV_[21+C3S>
?I:Q0.07a>RN4dJ\BG#H,eI3Zg;_]?c?UMWef;82aM;#C=LH?Q?U8C?]fD;PDVV4
I,T[^Kb;Z^I5+QD_9GBG2_L.UeH^+(eVSK/M0RDOF^LF9[bOag-4X@)@ScH5JW/R
Ka2JYD3(cZ\T\WMZ7#\[a@8);<QOSgE+@)-5c,:L6F&:A/5/0dG[>F@dCg_f)(3Q
#QBFOW@5?G@Z23COC>9BZ+EGY+>EY.T-7gGA+CD(Se&ZAASF21TFH?B5KcP8-:<E
SVbc>RC9DIZ1d8U.[CU08K\_F,BW+\FRVa3?BL)S^/ZW0e=W=Fd5OEWe^F0gg)e9
U?f=WD3De_?T2US/Lbbd=e.2-^.SPL\/cfRaER=0b,I>]U.;Le<eK[QgVN;0Cf9D
+(gQW6IKQ_<M[L95:)@?8V==-7FHQ2HNde:PJ++Ideb67V/ec0bM<6=A+gaEfb9M
\2A[c&L.UN76[==1(Db@.bIA_-dG<Ygc^9eOIMXRR3PR-8TO0VQ\Xc;?TE(Sa)]A
WGDV-^XB\Gd1eB7BX5QVFf;4-OH#HN8e.]4X#c-8PVe2NX+DHWQ+a909\.gf8G0g
bOEEgB0J3,aebI4ST7^RbB/&96>?79CQFg+^C?RcWQW:(9Y2S9cG1.=<H85X>6]F
9)OZ2gV6<W/J5_D[TRffWf7&S=F=K>=\7P)J>..ET.1BZTEb7>b<#K&2f[H/V>PL
S,Q34AAfNMW[59/.#d,;PS75bT\OC;Z2T4;Q7Oe4(Je\ZB+HY1gO6/1e4;ZVN8GE
#41gSWL.5@+,XXCP#51+#=f2:4#T-B3U#J&VFE@Z0O8>Q=2Oc#B3dNG\+:]6eD&F
O#T&^Xa-3?_N@B>\E+bZc;6@B;ScaUXQ\aKX=e-DaI)OMaTI46_;E-g8XB]8dQ\/
H-[SW#G];^+L(L>BbRaX/G=R9cc9cHHC/KfI)IIfaI3=#<<9&;b::L^RQ@I#d]Z3
&S9YcNdg0P3].TLQK,C@47<)M<@7S86P6Jf)bEL4LSPIP^Md&fUL]CR3H@g4SED_
@e]M2/F]F9,1O34[cHbdb/O7^GEXGd>J1>\J&0LKd?9Z8d.XV<,EV-gGC@QP@1]3
TR-<S6#H;&VfISFPIP&[NNc@<40JK35bV]N3.WNgIKdafYP1N]T5)MJ/DOH@2ZCS
2ZQ0SA]:3;Q\5Ng\]00(WVW+OVUX2+TV_G<8GY:-&\W;@W&e([W79-fPHFNeZ7YS
;c;\/f/]MX;=Z9LMY44:(GM(@eX9IY</bG+^La_RgeYJBKB8S&>7Bb:MfEc6HB]]
Q9NR0G?).8(g-)9OV=c>gRXZg,4W.W^b]>gY)Y]L/&T-AE(:GBSW--VO&=/X0<>Y
g_^+]:^b0#A+T4Pe\3S2^Zg\Q6KOZ+RS-VK>0/-7F<P5bV.D(IOZSMDO8-aWU>2L
.aKf#4O-EfAD,0#IgDPD-K(W/FbDf9..+gSEXG=K<DP9J.F9;C;WbfbGK0^a2H\a
VRI8ER_&ON<7+F#92DKI=2J]@_;)5[LgI)F7IYR427C;.C#S,X1-aXI8cNd&&ObI
2dD0Qg]NOFX;d[&7A9?YgN_@N\/=SQ\#5;]W0Z.ZF:A?c,C6CN,4JR?H:?W_ALD]
0,?IWAa.;[39IJ./EbSG_,c^K@][H+:c]Z&__^JIVL4JR?7b)K^;XXb@P<GMI^#a
J)[HT3APWQV>7)QBU6?)Ke(^fF>Y9;MdMAF22cBR?Ea7,[S\=]JNaOa:2Z]\=NE#
6HC[[g9,U4[MCU)CT:Jc@_,(M,S8>3T,)=OK:BeXH+#;K+cV2PDDf#\1=Q,]FF<R
)]V3V2,D0E\=E#WC.6WBX2[/?;1H7Q3S(U/7;-K-3W6YX>U_)-g(X0Z/[O;IAW^4
S,_\[R(4DDfL\4PIOF)MB\fC)_249RD5c.<N1dRg79fgA^40/6./4]L_#4,S\I?U
J9MDG[-(8Qfe7e924#c\DA9J0OgCMMa<L\SB>Wc<7XVb6=#T_G8I;B?^MbQ\SfTT
LW2+Zbg45;6-f[(H+-Zd^e3MKRbQ+\4&WNU/_V@^N@SM+=#\93)7187&:^e16-d=
:-PMF^6MWb>:<d4M](7WHg&Q0?81F_:=5eX,CE]GA;]K?DIN:W?K1Zg0X;WMYNM^
)5,gV[O9&D,,FT#LNKQLQA&7E/9C/]@ZY4H;^>QRVXfc7J#IEe[Q2I0CHY-T,WS5
?=<>@C-)e/OX^EMK8M26,VB&:-CTQ_5dg>GMcAD)Zf^2HFgT;Y43?Y<DZW@FDCR[
30,?42S9BWPB^NDW_Y?76]X.,M.bVU-Z>/WK,HMPLS>d8dfK(T:+,L7\@_EM0(?V
&6GLM_CUcK5)bU69\^\bb[RHd@F@AgPRJ>Ag>X6^T/MdFSX6Y=;IH6K4X0BdRW:@
,W^L?L88Xda^6I2QHAV6NFKEg^@/.3A+P?WY\)DBeJBMOg]gC[g\:MT5N58ZQKg,
B9\0R-JCd]6XPcTMg^KfeMZFM9#21<KJM7+2?e^g1I.cJ6;a,@0,(OHB3bf4Zb?_
]B;9>R)HO2#U-f^]f=>+QEA\^9IS:Z8d4@:+<0W5c/Ga>HK@=M&3\5Rba=?/73C0
)CfVe;P_IMc2HM)ZL+W+ARBd)_YH]79L[>gB@,c?M1aI?,FdT_B7?SfH5Y&G;OV/
R_Nb[U/dM1ZP>J;Ab.fMHKc_8Wd#a+/V=O+J2b1(aT#/GBVEH1L;XIG).fN0gOVa
SCY^/]+DVPEX2,<F71R2X4g0+\VL?a[,[,0LKY\e6,(X#PL2+QJ2-VO&Z+3UVc[^
Z#>0ab?S>Oc\Ye3G)2)T.#(#,ZG:YHY?4RYG21c0MX7)2B\;_#8+9cb@@S-O,aH[
PAL[EJbNb1F7XKbWJ;MccQBCVJ3g5fTRX=VOFB:3d6J_/P]8.?gT)&ESDa+f9F@Q
E](57F:a/8MCW_NOU;]aS2#WE5@f93MTR0CV;B?:Y8<0<)dD#XPD[4Y@3_Oa=.;c
.gg;+/GOZ/>,8_b\Wg8?0L3(0SQUR)f=YEU5bYUdDJg_P/>J_^Hb-43\>&TEEDM@
Z#-a(,/1TMBQ8aPS/YYg)dZLDM[I4T8EKVe+P]8G?^c.@c-P,>,I=;67B89?cB<A
f-=5Q6G>ECC?d^>25Z;@_(:E3OR8X[6CGX2a38\70Yg6\(E:O^#cW)/DG6<GSBMC
=HB@^M\Fgg=Y&=XN,+HM(=O@=>bK)>-+C+A\-4<,HM+1HU4BS#ITVHd+E^Gd=50K
]G37d7]@&UJ^([M3]\BfYS_a?EZ=B76gJ<QNWL^_Ob>;d9T;/P)f-D\X3>=L>ZbK
6/5;@]V:ELRPSR<b4IHAA9\+eX2M?Z8?#9&f\FK?Ae6HW=:,K_fK#g-0NXd46#:Z
_II;E3ZAbSZ)1F6IATWPUeZ@@G3\SggM:5;EGZ+@K[L2+L(MBH)GIdK5_\.N)[#f
=C<f>S831bR-L,.M,M;WOB&&?T+E[#:56-E>-QCJW\-b&YNc33G#.EVH;a<J#gLQ
CV^Q_<cT@MMTGQEOBT2-P<7gRLWC,[N&L0SL\efX;aICXSCR[F)?OgOTf4LR8c;^
g@SFYRK4@M)F;_(ZW+-DQP=E)AdfQ&,D<N#SCIFADQ>X?]-QS31[JNN#W^C/E?QL
>dc(;S]N[\-7KTgV6Z@D=5-]H^YO@>T(54.K4bMA_FY>1C1(3cN5f:gU2_eZd3NF
c&2ba@b>/NY_CeF6@;#;O\8fcf24#R=Jd5TR6SVc[H+/XLgSB2QDe5E6O4;>Wa_I
\,^&fSEI]82JR?IRS(QL<d?O?1f?eZGZPKDTF>a5\=bfg)Je9T64-:eQY-3=^W#3
&gFPffP4,+>I,VYS-:D7QJ>YQHW3BE-0TS/-ZVWKgF+6A_P\KPWH=RCcJPgfeffH
(I2Cg)B6:K/J>gg/77GYF07MM&Ka[=TLMTISVS38GQ)LIC+S@UAU;,28bAGW+\Hg
OC/5Q?N346&XP+H9Mfd4+4]@_IEF.4(]9F/4E\EKgX;>S[NQO;5bgK<g<&OE-Pg8
b]PK5)1Lc&dFWA+NR>14XI@QALe4BLV[>OfSe^9bS]b>^+[=(<:ACG\G:c2H.Xgf
3F-6A)+,767-UP@IgR:\.()BREfY+H(4bJ;<F4_NZT7,9K@?C>;;A].,,(,G4=F]
WYC,]TJJbVBV]D].9^e^XG<UE7dQ/;\XL8a@2HG@f#T+OHIE;\:JeX\ZZJR)aW7_
L@Pf/.g@D:f;PYI[X/O3aeQ&X=U\&B,HJM7gcZ&(;64ZUf,ca9[C7de^^#a+&WP_
,8CD>0@L)d5JVMAU(:WNGLR^A54c#+4#)3UA-Y5,b9BD&6/+)Zf.RBL0b-]PT<9@
50WJRQ,55#-73DZ1WG2^&F:7.0B#@L&3M4aHB?LHA&d@aHK_92b&&4Z-GA(AR0B,
M/=;,eZ.&@+9#TAZTV\9>=.@E6/__ZE&a0)(8K7=N^-I3b4QbI@YD6^;LOTUbbcT
)ECUT_D2^@8feREGEbKD8&;03DB4YbSE^&&Md+=]U;d[B1+\&YM\7:>LCZ&L8G9>
R6)Ic?\_MS:g74_+]?^\FT+&]</;K-XN[_=[73;ZaC<Y9-bXg3;([WWf)&?KR<E?
L7_(0ec2fU,X\M?QTbRB+-K8(YQZGIDZ_8GYBFA5P36eP:>Z6UEc9,ROKPCXHK5b
@0L1E3RNfC\ee(]6/cSa[KOd9.;(1(VF&Y?e.e7P)f?ANT#HdcG4g[3139PNTLW,
63:?.\e);H9.Cc56:b0DE,+OOLX]Q9?1egVK?TXT37K7e8XVg(KP(X;:<L193=LV
:KbA<]KeHD#NQI6.g_3+g)KAb1=77dEG1:9=]Z(<;ZDMRH>4c2&WaCC77S_MW3ZS
0B+@B-,LJ;>+T@2DcA;2-\E/7C^fPG\A;]=\=B_2.fUGDc-;F(4(e.c60b\TSQ(V
<_(&Ge_a,94D8-=9BT2HJN;IgL:_gY=VX7XDG8dGY\N6fTHT(?33BaJC0<9MWY\T
)YF\#da^g:)e/-YUM;BJPIE5>ZG90>0<Sc=fJ6R75HFNVY,+aR6NK,\7LEXCbd0/
;2fbG^]\R1Qf^<M7G;Sb<P-K<HI1:QX>;RcdM#6bQE7ZWLH)/UE^:X0E]fU35(]H
-F^,gDD02FMe2gLeEUGK06f&2Q\_cAIfZRZN.LP)K^=7f;YQI:5b8=f;:(IA\K3?
XY1d&D0XYO51JXL9>;gE^3/#_8WT,d,>R+>->B=fIMLM_acQ4ICWc07;:Q[fPWLJ
1ZM5N)N[Y43R>EgAC6ONO+]F6eN/,F@2ZXS8\8OfaU=.GFVQgfcDY/144F.L,XOf
IS@VTJLK+?8>43V)ZdZQ4PDKgUM#Q=K?&d[#W:+)0E,AC>N=09eM8&J24:@9DFB<
FBB\B[GF12V239_&2]+IO4O&[[FcaQS_^S0e4YGLKPDLa\?Q4W4P1AC)]U0Ic_BL
_C<b#N=.6LgO@=J]1D:aFDW>J<H]U>AACcK3O^)?N96M\cP<f?CbCNJ<JKZY>OZ9
BgagBU@eHJK8@>ZLaCQXO#DJES#7W=G3_F45283&U3==Cf#46W67fY4]J0-\RRGg
[g60<J4+fY>R;3)?[B#8/6fE/RXf9QATWWWW457^Gb4O(V7)>Z_X^f>eP3B#447;
GHa\T_Xf<@M?PE1F.gE@c/&&;aPc@3\=?DFDG.F/A>g]6#TH2@V-DP#eHM?/UL0D
^65Ya-(TRX\fGL82Z3XP:4I4gWR,,);HdKbeF646Z#;bfaV7;fdQCK].\]SI2]8.
G+DZ)PLR.-(6A#X]B[)EG&AN\GRC65H[D+aK?<8f]Y1\_ANeX=H,>/3@9;R>LUe.
cObDG;5ED0@eL+UY=_?[-/&Zge^7L]K8LDfB9U+K0IZ:/KCOZS4&ZK(VLTFLLH6b
7,dKJZQb+KdTTY,)Ka]TJgcIE\K^K-:PCE<a4@>:5L22O=-dOTcb<QA=X1JgL>,I
^(XK&:7_<2S^4ad<=KJMK&EBIEaB+/)T2B.e24<2BIR(1MX(.(EYE_549M-L>/49
5)a(>A2NAab;@&Y0G17=N:Y6HaAYVYIU@.&YCD58/1RZBAW,Af&>WEDedQU>H,g/
E4Dc6(-)eUFF5[gWFdGMN:b]TYD>)E3bN3U13C=aU,]\3[TE]J,\9.5Z464a99SS
TT@CK/7[g^[@Zb\DOJAVU<Ifa&GHMN\SEbG=SBV7;dg(eFEXc\)8/U@Q:Y#&>&B:
JfT[8Y^:\;I<0J+SW;-R)eCKbL@9VD,;<eHIKd^RHFNA5dE0eT-e?MN]g>JY3^:b
-+PY-LaS+HL)2E[D/:ag6#T+\M9561_N;B3XXBf##V<SN_>-DZFCTf=-&22..<Z<
6Z\9>\&Z+a/Rd&a=&_.,/H0NF9_)Le625gfN->(>7P#M7N)X=+M+2OERK440=@&G
O95RY\R5#,4)aB3D8#8MLQ?YUWR?NO:]56EQ\QWeV0?7Me1[W,_@#B+I]g>QPM1&
4W&/]G>^b2DdF#748f^g]IX+AHK#,(dX2.-:7AQQa=UW:V[^K>/DKT83[=FFK2Sb
S@4RXbC#;(Z_?3J;Z]0AY90EP47#dNCY7d1.,3:0;7PMTf;B4+<b23B;9CI?A.[7
@)N^HN/Y@7Eb6dAV8UO-KK:Je/_IJU?0RJPOE/B?6Ub[,9)F/L@@=T)X?#4#FDO3
7JV<<<:1S\J3X+D(HbeJFa-NcL2GL=2M_dGT.^-;DD0T8fF)b_MdDM)dB^>1Y][I
OLGC&HZL[NZ_C[VeFYdJ^[eM_O#M(?+gT,HL\:.?M7Bf=BZbS/af\R#&9Z6VE2fL
:I3&,9;N\LV3VY6K[TTGd9cL=T]-)-#;:fe+7YQINEWN)MD@2;)>RET[62IUY9FK
N]6Y\F>T_^[3=>H/cVQE:[N.1IgW6B-WN,8RF>Sac=]]AeYb3F>2<HW-MP5HSD10
6:]Q.8D\dZeBDDD0S5GRHd.;)W1YH:<aWg1PC[1-\XY62=,FADKHKF-c;]FUY>B7
O+X.,WV([^RF;_YD3#E:8?bAK1VNgL8N&f5&9QQD?eZ56b=644WD+^>?ZIDB7CTR
fKIZ-7Ee/_0[^4FH=M3?M.DX\=D<;\MGVa;FYIO#[<[6dY3.0<\X>Rc3\J/:(8\[
IK\:=P=BI\9M]4)_.9T_.&JXf-&(#J)A-UE<@<N#))d:PB6e>_#HQ)4;_,HSG5H>
=0)-)Hb>>>GCLf(^BLdJfAR;:&>:Qb5@E?bJ=1SBfY-L;QG&H:6(E-[aCa4E6WdV
;6CHgC6eX\)A_\[JQY[gC@TR3.]eD-g<F#8d8AJL/TYK]T0?M-LPS.R;Pf^:ELR[
VOIJ/008a.FOA1^4#KE?:XJb5MS,d_8GU^M9DGT#WebD(F\R>9\AcB[4&W7/II1O
VgT\?aTH0)RU_J_<5LG:^6&:/ZF1XFEW,:fIW:(^^[c_gdBO]=P#AO-WfL_9g+9S
fK;eHGO]XD>9X#+U.&Aa_9Oa2B[g[cSC<<2=4HX.+KSL@UOVd+[L/5L;;6@QZfO>
f,-<bfK#K7AF,?>@R0B&;QcH[fH3\Z_O;e5a9YWJ#COEfd\4c@GG1;bf^:,^Q#)f
:dA&4,3]HPf)3H-b(2Y>.1;gK5ZfZ(fV?HZ-@73K(f2TD;VB>Z3Kb>IZ<?OEJWHY
e+-9NLdFZ,9[18c5;[R0]A-TF:^Q[[4bH/,QKH6P:T1K;,2e81f4&3TH5d;CVBHg
FLb^#.K0..U<1R3LABP9+gLF4N_3F8#DQF/Bg>V6IXCW(V<d63_/f6@#;HBPeA<;
_017T@]@T5<],CKbF9&65d<T0-^RT5,53fVT.>D#CJE6-[6PI-dV[(MN9LNFL[M=
JB?Cf3:47:MK0Y?3#)IAabPY?+A5J4N2N6>?,:1<)b@:d^\+cG/L)63Nb.W#.CQT
a#(c6HP)a5@b#N#VK>&UM-2,[fgHC5d@C@M8ASV/?dgVYCPXVB9;Y\d\f5YV@02V
;JTE8:AZ/e0;LKG/FeYN#@;Y#,;&eRF7Wc+7_Af)(@T#.3<7R@BFPDXX)-XQgX64
&K6fWf2#&L>48HS^Q=aKVN5V)M<&2QSdVSOYMQ@96<T-Y&->=>E9ZA>1N8Yd[W6F
@QHb?T0eg=Z^dBV[9>BMLZd)Wce;>V^6&c^>S+O@3e:?(,F@T-S,JbEIPEX>DAY+
FEGO&)TK,>X(gCK.6B:+(eU0>?M)HcL\3__;XdNI8b1^0<6(=M#&]PBdd,JE.RF(
=g\I)Y4=^HX5;g:\+OI=4@@fba=\U5>-&&&8bJ#@K-Q.^=#\)KcaO/(6?IFA39f2
CW])SL(d#UfTKUg]RZ\df9d(H+NUF))TdYSf]U<V.T(e34G3#5>?X7D,Ua06J#.a
;ZD;LL4K-54AFaeU+B#-HTe]YRdO^8Z7^0Tca8YLU@JGRBV+aE?XU?Z4Fb:cf,,W
_UCSNX99J(#CLB4NM)-MDdB4BUGCBbRN/W1&dX(&3/+IA^V<QKe:>3H>RZJgRH-b
\+LaWI,X0eQ=R3aYJ=e-,J6?#VIV9)(;;N)K+f4C74SH2;>K&SN+FMRf_d[ROGQb
W2f\Y=0<7g+L]C0=PD.(cQ8Q1]?W2+KZd)R66GJRI,(WV/B3RgBdf2X6#5P-U^?J
[+KbK7T#4<D5-4gMg(J:K^\_.a[?EdLRCBa3=Id\L6YUJ&IW^.?PX>.3.dc\fgY\
G+MId)0g:H3Y;a)JGWPd>]cP41;cFP7&[424]C^1G]#H\&[Ge-77bPH^0_E+4-YG
Z;B/I^?\@VBTYGSa.F9KV,[ZE:TB1I4^g6GJ&Td+ZS&5WI>_VK]8fQ<ZQ@aR:I<I
H0.<J-77@1E0[887)Lg5:.S]LKB<41S\2RRF#g:[@QI[W2205I[cd8[dSMPfYS[D
B,3ZVN=Y>f4bR8@_OQYNYTaZ6>4.\a53OM\^/E<9/#Ja,D)6FMDP4YNW^QCC;LB@
R\<7(/N/-:NH.D(,90(;3[G+QSBc9C^B<\g9&@7;Wc/M\V=FIWZYD2?#>-J?OKd-
8UQ0;BZKU.EG/>OH9YLE@,V)NDU<B2STd/f]P9E4YNUe)RcUMGTRL@6@?A\(>=)a
&\A]5)TZXA=7U]^5A.IL@G1]+?8-1VYfSS)(V_4A+P>^gE/^2ec#g>(0J1(8^Y;V
371g1,=HPCTfeTEDE>V:7ZG]RFeAFR=LX7S=@QYJ3J9,G?,L=KEg=73^1Ja[HWT#
^RD^+QVOV#Bf^,WL(d.<d04O-Va3g15,>\Xa[M)0YHKa@EM2-49bND+;Rg,TJD87
]7?&)ONYY?QG=QT&=C9.QJ39>/M.C?\XK),dG7\L8[Vf/R30><(C[NgLcJd;\:UC
_gS>b5T^]6]]O.4D_?S@2-_U75X7,4,0Z1^WS)deCG)X_2=Fa#Gg]KGAa^]VZ>)A
K1a9Y4O&I/BH6^;+GA.\91f/E+3HT=UM).IYe:eMO.1^ZXJ](E)1#fQDC78N_Fc_
@:L^5&D^ad2e+@6DC]57=+dNNgKEbVMgVAUac/--\[-9J[5#NP#U^Z>KY2cU)JR)
;02.Z-,K3LH593\^XXA#C?B36Aa(JO5&\VSLEAQ0[Z0)XH^N3Sa6Y@Gd;^36/2LM
K0OU/a+0g3E2FG+ZMUaZacT#&R_U;Q6TaZ=KWIUH3BgS;,OZ)D-8^Vg,N.5=I)?E
QQCRDeP_9R7L8MN-\K@gB_:T5.30EB4F<H[Z-0e?/G?D^Q0(AW)?F#+H\0C^8#Ob
7LU@V5#:<=Y?OS\SbE<-7UG#/KTcE+-H/)_dK0gF7bC7>OBQ]JDC6?:0c#-Y29=7
E+3902QH+F]F)]bfNR\(fX^,[E#PU31AUbB^fE_aH&MS4L@(F#2&&aJWS;=gdgb3
)a<](MgQ[BI))U#>3WO:\\T)>L&Pa1]\9YFC_A5dZ12#LX2G)+V8JWbO1.7g^c>Z
.?YI14&#bTe?Kb-@L&VBXgVNO5:AZ+<5V]dAgZS.?C/P-0_)N#M]\&4.g2K,O7XW
Ng>RFIY2+4NZQ??[Z)D&@#@#G7CBXZ94[V0fF#;Q5P_#&Redcba]3Y&)FB+1P8YB
38N]3ZV1P/Aa3_N>5:fE0Cec&3dS.d;-]X]@:[KL3aPP)\0BW&&L(J+?f<eD4QW4
><4I[^8dSF05#-UP2OdCWDfU,0YC4MONGW57_\gg[8#.c^3IYAOfXUEVObMKQ3Q6
7NA+__WH2,fAIR(&]#e3f0A#8A-\1;435fYVXVf;HI]@@/\DHcL+#gd8M?#&Ig?W
4EFONcg_ND:DRLPFJ/Me=W7YY4f<A&S]AJUFPJ08Y<Q=A]6KS?.6O>R:>L>&E@^Z
XOAN2>4IX^H/a-^3&VMEVE^+.60f=fRK;Y/A[K^BVfQFHXOV-Qc]WKI\RFSZ(+)W
1A=W97Wg.be]VE?2?M&YKQ],A0eD5@<69-dSLB?UN[@-6>MSXcBG-K76eP@P^K3=
7a/)(b-K-1Y2aT\U\6De/Id]gQG55L&-FgW^be4gT2B)(UdE7V24[3ea+T1,TI&3
g6:J;O\GI&\2X&dW+;df)AgK@XRALaRD@W.XU@NAANRL[+0NFJO=BPYbS[Y62L,C
dUJTfR?R(U>48U]_FO1]\ccQbT;eS?aM45>81Cfg?AD#/PO=LcRI8,>CJ6bLg)<.
cb:,KJ6g<fWBE0eM<dJ13R]Y,@D.^_T<;C3XV-^bL/V[c##[>#c@2Z2ZG?&=d(YI
7^DOT-J-G+2Z[9P.W]F&d1\U04/.?.<,)3IWO?DgXbC9_][/5,EaONN7BVWV)-U_
\:RH)&QP<gLb:\6G1a1cL_DF)W(4NT4_24CK4:2bc<E)W76Cd@VB)Td0]?W5b-(E
QeE2=9b3Ce45IHGF,=;G.Nf=gW)V@@984]UEK&9)0FMAZNWK3_)LM>=^4N<L4G\#
HU<03UOb?<)#9PCf^3WAEc^#W.L/#0N54B?[?B0.F9\29bTP9S>fYCDfNLg9c=UD
fUbeWE]=>/[QaV0BC>LGR6e(Ce^F.D8(\agIG[P;JHb87LBMZ0@@<CRWIC3cO._T
^CMW)26a_a:=6VWAE,E-XLLe]:b6G,.^f=O5N#S_CZN@DQFf7NWMA,S0J)6W_53D
bLD)=2VTVa<.<Fg0<^5=3<-N,X^_7C?&TAJ&S1,/6cJ0fSOHX)0AOfb>GXe,M/g-
fcRB??,J?07JZSZ_C4b0dS.Yg?P_1D<>I0,YgW<6O5?IJ3\G4(a(gJ7?(?VZOD@O
M)c]3IB?#<TH+;:;]R#@-:YU-/9eaLT\:&U-[CUAU1U@RTGU1++I8.8d;VBJY+GB
RYcO>FEZXNaWJK71/JK34=L@c=5dFN;^@14A@9\;4I(c#-#,ZW#cR7@ICR=e1SP\
)J3:S2bWCSb?e:aMZ2cM0F4Y3LfL-\ARdR7(e0I=g,V@WWYaM;Xa2A,V=:(J&cW4
?6@dP(_If4PK3TK_Y3gNE-cQ-;&<8F+NOH1)bUNNIJUFXFS&<e)X;J=FZcPOF.UZ
9[629QTW<GdI@#/52E0/M)?1F0ID[R\gUfZ1-ROTBKgW:GaRcZY-c<7G58@F_Q5@
D78@gQM)f\F/T;dF3@QWaK&e.=A/X[5?M5#M(U+D5aIBSV&J]-+JN+?a&=REdcf;
HNYM1^V20<)ceN(PV?-T?ZPH??UDcLK7./3/A?8@UH.Q85NW<f5d6TFM:Q68#\]+
c>B0Y&8PJ=0&e+@e:aL9-&TY#I5,1,CO^_4Y(VK,K.eYVggHO1FSRf&A#Df@E5e9
Q&>O8G8;9C1)RL6[N1-V#Oc9Y=^IOKJE]#C2X&^8:?+KG(]D(6D1<G?]]O4V3:5Y
7=]<+aQfFG?L&,94V@fe9dUeHKf3JIP_:9:G)\/KWPW_aT^K4GA^/9,fE8?@fFP3
fGV-5:RDXZ2eF;/HF6;/83I^WT?]_bHW2N>XBHB1W77W,R+#)&_PZ-a1Yd:aQJ(N
DS]Y]M,VRP4P8fJY.C;M05GX,LI7b6cR[ENOPY)[,Ie\E;Z__>R:2:K6/gcT/;db
aCNC<96NX5_@2A8L7B+Z9F;/[\8V)VFF8L#(YEV?O&a[[0R,:LW^Hb]9;486V(1_
Z5)(3+PbE/d)?:L<3P6PAASZHO>dWUBTPUJ,b#=f8B=6_+09b3e;E:a?()fbP&>S
SY.MLQEFJ-7F++_=T8OBKD63:4_=2R6<7)=HS&]?CM\M\7<#,SJN0F8E40c:e;_?
F^D98c-H[7H4De4cEUVCML:M82-bdEX@.1a@];ON,dVLP6=N8XVA2F=I:98Y<\F0
SSE.9OW-[>=b.7R8WG+Ifg=M(3&Y\a,aJ\+Y#C.(VObTHT6UWUP&;Ye\:>14S]6,
X4CZNPG&eS)3#I[(#7PP)-(H;[-a[\G/3#S7e0CD?:Ff7ZF64OYCNVG8N=^J[\[3
631(NXCH77dQ#J?<\WW27:GCT7XO<M:XU/?9ZOX>:\.XeA/<K\57C(?b^PfC809X
08)PFM&MePg68^:O6#H-Mf@]64-M;0^3X6d3aTeZ?G_I,V4]:?QB/S?>U1SGKbMC
ff=]7=eNgD)SF6d(^E;I&58XT7Vd265HG4P<1U([LR:aHO,+W8f@7]B(QL?1CVVe
R.2gT[Ke2gEdd:X81TOX,YN:,RU\-778Y631VaEX;0N0/OPO(Ef:/1K4PX32K,&.
G/+BFTTdN0P&1^3VA52P,D16fZVCWZ@D9&XR^?TF/(D-]QREO2FM()W/gg5.f,I[
LZ717^E^X?d.60[F_E\dCOS7N4/PWDQ;We-71AI:LL\DR[AF3Q#adEMMWQ7,((\@
&3&;6<E+DZ.M;ef&G.Q,=3ZS?8=S0F?6N+?VgCM.E5.F8?J6ZZB8]4-eQN96#FHS
FB8BKe;.ZI)IF4,@F<^MV]R?QA11O6W35D1\:PDQG20-6-b??=/V(e.d,(@AP_:[
;H#Ie#V1U?>cSc:;?TNP1+DXJ89S5VcOX?#5LQR?=JDN;4QS@FTGgWg>ReSR:gFR
[J;7&D-P,?Rb51P:+,4.bgYL0Z8Y,<D\^6&VC49+aO=^#F/3W]PC.]K6-3-\dFYL
M-+<_2b6.MA@&c3cYN17W7,S\UbA3DCG2OaX]3A[;aZ=8L23J/??a_2(KTH<@&<<
5W)Z+T>(A80PWB_bPPRUaQ_N.1G.M+aDf82H=3c5>E<9)GV]efP7[_C<+:MAN?JL
^X>2=c:_dTS=SP^9:Ea9U5Wc(V1R+EX@?6:c8&O^>#gf0FFFW.e(<bY05Kd_G]H+
2^AL_W2N74+4OAV70]F)0e5C18Mg(\Kf]3G-=9ZK=6_B.Cef&81B+VYM2\M_.TY4
H73A/(U_/#99d8^fEX<^;ME\WL<V@c9beZ@J8A\_UN(cfeSGS_0ON?f=Y_TN6UGK
5e5+R3&2K7.A>X90ICd.6O?,IM8#Q>+X9V_MKH&BU[WEXOCLM0WZQ7Ze+DKe2U=B
Pg8GC/2e[/Va<^+LF,TcX6;()9FeVD9X?UN?T#c@^UM]TO]-Kf?f^_c;#AGBNCCQ
Lf4c2,3BK-7=f2=.YBCg0Y:PC_?_OY<-.)(CBW0)fUK4fgZS_SLT:TWS=J79,X9f
1E/4@;\Z_gf3J#)f9d3V(D(5N-/-&)ND7F&;.,La/)YLN<D;\V^EUbgEIJ;DOGNa
,K8]YBMGL>0?H/aIQ-Z0c1==F&A<5QZAcg^b2bYU,]C)gcRa7d4QGY3H#2K&:^I#
)79U<;IbBYbPSe1fa\9W,XD@RWA4EH_=b;PB/13<Y34IP:,CK&JZEP4+20OQ9JN.
_a/5A_+;F:O:A7&Y^H19dS^7[:gKgL(Qd]PQ&/c2f<:2V8Z4>IFWbL0@3-B<3CS/
AQcd:D1YA)aD6X,];XBP-/f7>&C^MNSB/7XJRdI<\3fE((4YaaI19](OXDJ_>OD5
,fD#BG)90YeR:K7I&f1Y?C/AY3IXcX9Be.#KPPK/E2PWV,#,JK0UNGAI__K60.FJ
RH[aQ.I.,#@-)P8/8=15J88g\IeW]@J_Va(Q83LIaPQ8.6_1J)L>=[WFg<<O?((@
(C<f;L(E2TI5D2S8JAM0A:Ieg.8GZ9>S(XR0@Q@Ve-D]0C2HM4M>CSYXQb.<C@>;
8Tcg+KYSZ7OX<@YPY[C]AJ9ZfI[a0gF]a?2RC5BQe),D<N^5?YLE5(&B#QUFbT2?
eS&_.8X:LQ,R^&S,F#a?0U;Ec<.9YTdVIC^ZHJdT794e4>_M?VdH/2@O2+4<-X67
3^CCM3E1X&-LN/1]+I:YdL3H/R(.U5V0Df29b^+ZU[0?WF<)^BCSJg+Yc+a_,BX>
N1V;NCZ\W&[3.85=&.O-BH5@fX:g@05^AWV)1:_R1a+@0W?=C8-R_=[JN)?d?G@I
WN(X4dU2E;bC1&6MA=]/8Ief[3Q7Y+Y=<9.G_W9@gWN;FDRN/TW0a=DW2F>TS49e
,23RR[#POLSAZK,-(Y;,36\T^+H=KXgR[(XaWWg_<K7&\T;#RQTSYV3N;a7R^;I]
8R>PQ/5ddH^aD?A:QB6[aW?I[8RH&#gg=#8^GcN,6TBUCM^gWEV1,;(gS@4c73Z#
=Y&eOE_/e,,GbJ[UED38LW1U_X6QUW&YVaN>+R]E6NG2e.YbXd_R3F.I,^>1FQO4
CJP[[E#@6\+Mb>.TWNGKEP>\69O63YR<#Z_S50.cPC<4@EEFG?0D#:_Q6^ACbA>(
4L.I/c3;7+<H]aeIX?5P9J:gOG2;-fM/Ya5O>[D+(I_B=MB=>@e9WE(C66S85QS#
:.=I+AKH9DGbRD,]9]/]M&)<=N:),EQPd3/b:>1_Qd^-[6&>J#cTALX<C9Y&KKcX
Y7=4EL9N;5gKJ5#&f@#-F?.O5Ab/9H?M:B.?.;P:PX=/DWGZ._?R^HBH;T_Xa>4R
PcGe08L2?/CX[1UMCg/N3]B)SW[3:<FCE]0dUEPTSEZF@.(5Q:;(-8ccJ,<R(&Hb
W0g>^H>Lf:+;TNe/eI3IRT@-W&0]IF[-MadHPfO4a5Y)EQ5IDDCe<Kb_a\VJ65Jg
0Qd08U(&ZB09,Y#CJ>6,(d=@g1Y6]1aJ))5<?LFG5Q[O715\aWL<98;67GXR?ORO
L0cc;>VdI7D45Hc&RcUU5)D#IbA_0>4d98HZ5O/-RGRWXUL0PMIB?f4gZ;dY-g?/
M8A.Q6M(U#f[bI+FP5<\HdGR(_Wf]9WY5I[J#HcR83^A@L)a9_[e]:&f?5U#aH&R
#e6d)+^_J\>I<F0AX3;@)E(QgH#:9<64>N]g+gSPaWXJOTX38USUTM[#9.S,dG6[
PKH?&A+=I+bNeG[+gdUXHPRfdb;VVE4P)+9P@(.Kb:OZ1RI;(^]:?PU.K><@)XeG
7cA+d2W?1-V[gBddO+75RVY>ZB[UG-7#a<VF^dDPEQ?YbPIEB9,#I2\\?YCX:--[
e9^E3815\U#H+.0M&Q-[U]YR\aV9..F6<+^3D3I1.P_)/-J2REZRc;[47?/9JAd>
GP21A?HW2=>&ZU7]Z?P)gM@eB#f1H:=Q+>&Z;2@BR=7>^)&,dE:V[<eHCMA]b(I-
9T.3]AO;WGS<_JB]0<a=7=_SIBP7=aF2__-C13WHK@DNODeO\OdXRf/IBD\2NJGc
9]E?BKb0;bA-QB;5?&,IbKLfBDBTN,]W@>-6M40W+63F&L;@]g#baFU_>If)>ef[
Cb.FbIW3Z,7ENV&/,MBP]5#H=4HTOTK6SKW616YGZC2c]@-N#^01;&SNXOE_Jd55
<=]U7\3g6HeQ(+DIVZUJAbdM,]d2GDEGWX-S[L:SO++_3YcS)\\VYVPD\MIJ[f#,
K3AM&W,fRCbUWT^Y;aU2.<1GQ]APS@PEEZ1HYXe3R(GRJFc3N3A5NO6IEM@O2L)X
2)Ngb&]<&.d4(&WLW-]gga86-Vd0X_Y4A50//(^[\Ecg4B:;I==W9E@BV>-3D[O;
.#=N7_0eQS\JSWVa)g]XF]f<#:I:c)ZR;J&UAcXVFZ&0ZVTb9P4;]ZW\Uc[KPFY6
Y-a;Z<-O,-FcYUI;&/C7G4@:X-_S43T#3T1eLXH4\8IJ5/-/&._e6S9G,PU+eI@<
^J=f_0U:G6@)R]G#N)Qa.@]IIFRcM0LIR.#L10#,]F=3E]57XPG=0W77,IWX8ALX
\KR:L48H@3;0U@X5dJf/2,7)YCP/6[@U[cV7RU[1&3ZOAZ4H#\X[\PW@G_]cAag@
F[9.218O+[8,+4W:PM46?,0A^SP0bfEY[EP_d.+7CTL=2ZLS<Qf)gZ/N8G?C0VQZ
=aA@X(^Z_>fJQfWQ3,07,&G-.^Y7GO:.IfB+fe7bV57[1N9U;L.B#SM.G[CA\#Y4
P.3>WN;I,N(@&Qa7.(R[M_JI]ea[;f+[D.8XF>(VO^MI+VQUW((P9Z1:(Pg[06&@
?Y@1OOU,,EaL0S[aG3[[68)e9OR-OIC]c;GL74@]#8d3N_VVLG&7@_;LA+(E_f@:
+5[8c7V4W39BO,T6;V5b1O)O&205gCbGSgW.T;XI0_fALJ5CWfVFNe6/,^e&/@-@
[W)c1dC3PcD5B\@<\6)DH?Ac<6/@BL/[FE/&RIE1DO@=F+?8+B?B?1S4@[/ES;TF
>[2_7+9-\A+c.GIEe-K.)6#-Q;LONE+K;gB<+MM3(_]&H1gVN@I<[<3_(aKU(C_7
CYX6CAN26dJD2(5]:DDdD:X1N?R37VKWf=4R?I@/;5X<@HD+MbdK3gNOYc,+eN&[
O4\RAUKb4B[cY>YU]LK\fG[PLd#9?@]RAA2X4ECY3H44]7,1>V[J:75N549]A]S)
cU?Ffg[&&3E7I58#;,(NKdc.GEgM8H4DGXK24E88_2EF,Y9J_@6Lg>McM)3\)a?X
R=ZSbAS5O582_JRS32V[7R&KQ(0.OR&A3.MRDf8+7RBD]Ve_LYLSfW\+c=aZ_f3a
5L(KEC6cAAM?Hf80+MT9Re\[\O^6)5]P/\P))VNEBGd(cU&5QQgDSaOD=EM-)YF)
,506TB>aK\4+a:/8ae.WZ>Be^:B.bV4(K\+S,aUF.bAPR\:IG59XFGIE<)LUga.S
#WKCX\WeEACQ>IR+]f29RO90U<7#[PY=Z:f8dQcE982KcdZ8LgQe5_[F3>;a8U7@
Q77(9T)(^ALVBLM432PPC<.Y_47B]9N;S;1dB4)&;&(2YXT.^)9eWA,QC(KcEEJ_
]?<F1cRMgEBFeRRVf+be3LKgC>&BV1(dCZA+D?Z[cY4H)B-VIE^D8Q2E5M<-U#AZ
RJ1&>TJ91cXN7/F[GaUME&d\)d,UTGIM+DXe[[9[YL-Ed&/T>,60J]+Y&P7\7A0>
dZ+P.]:WIU4S>/>H7W;F/F[&1<:567ET^=d1YJcT5f@a/-I.3)[EUZ]_0N8G[9(B
,\WZ4dN3g^H)L<J,8O<,MRL8E6<e)430.SJV.;L]2C?fJSF.HdG\Z-4f+JCMS403
Y9UM(fFY2g&9ST0OZ4KRS?E)3NM6<0aI3;XSN:<V,[C^DfX:6g98N&:/F41ZID85
.A/0Xf0faM[7bWb)&^[A3[KB(c=8]6->4XdMQaV-/<aT>^VeO&&g_+@cRC^)W8)J
Ka17KEQU?,X6?>Z(ReWSE?Y_7H@Z-X(J?]Q9KUbAVQCe>][^.U\U[IF]7,#9g-6\
):@cVWZ0_B&b;fX][96T>3;54\RR@P<-7cR5\Re7F>(:A)HOR:IBY/3[@ZF9C^,3
3/c>=Ab4ZOW3[ASZAOGYE)1SAf+IQRX<cB-E.dCQ@3@WZW53/S#e\7C]+JeGcaSb
1\(Ha^SMV_Z1J?9OW.e^Z:0H=8c7.6X#=9M)R3C>S^.J597ADZ,Zc26JB24>W(\P
TD6fI)28c6.@]:CV4=5I.8R0)\JUg/[</7,DE]Le,G3e3>dT\]@S>WbN9>W0[.M)
ZZ^BgJ<;=F7M&+B=R<JK@JEWYRdVPJ^_K+L:\b_0D@\UUNd5OYdScQF0BYMS.V05
XJX<9@1d].4^(Y8#;)T;WYSd(CK;@Nf57>ALd<O>L?SLA,8QOQ^EWc::TZ4SIYLE
57;PQ/?-JT_.abO3TR.S@f,.^+JA(5(<79L^LKXD#>YY0\)>VEM9N.XP81G&)?gG
N.1W.ggG&JeJ0-H[>V2Scd,8a.@Z81Q)SCN<E.(.1.0E_::&bKWWV7bMP3BY<E:K
Q/)K]aH)F;aNG(B;Md?Pe23b]<B&d25[:+9)(8=8TMfPTNMW1GUJV]g.@+?0,Q3W
F8+a^NECPD<OFa64E(^HXafg#.H]2eUZ/YEYF7a^15.2Z2-3@I1P(DBNbb\OP5DX
JYYHeLH/^-)>RQ5/,<S56NIgH\[VI3IGDN>DH&?gG^cS9d+0MZ\?DRZ&RA2e&;NP
KV)b5^\.9,;I&>W)1fRQ]eeM-e.F=IC<_/O.@@U@NNPV0=;e1G1FN/[7dGNPJB>L
d<YOUXU:ECLBH4ZgJ[aMb1.(7AIDB)>W9bY[XPI3cgR+Y/#OdNc;b<CY2ZK>\R+;
N<@be5)Nc3&(IMBWOHaGDVGD?MBg,WG[A[S\.Q6PAdRZ^Y2;c=VM>^J/#XY?P>+7
OK,_R^(\d.\6WKK)5fF8AE7GD-&L0gTG+>JZP>3:aIF6+@I\Q_XC3<[^7R73#?V)
^.;HAb+9f4ONLJXgDTWPEWa+HU&(57K7_C:6IV7S47\ORJ.V)fF38eGbD,&C4X=9
_5e_Rd7TKCd:L[\;0S06e5;D/^O/5B8Z0ZIdS@=J337DD<-A@ARB\2.FUdZ6N6:[
3a.gBZfa&U^_EdFGcO[K=-NT]G2a=^T&fACc0fFU7cHJ?G9DZ)B<++;/[0IB5I-X
gQE:,\/^1#NC/IKa:6;ZX@P-B_A&M<^\JN/>VFS8OW+)S0L=.99?cQ]60D4H5F\O
0??J[4K7(#.N=8P>P^<V\_R-GO0g+d_OPOY[+_]0d^aXJTCVIAGW^\2)2dcbedUE
a2A:M,PJ<M,IH7?]GF[.?EO0+BI2,578QT)b/ME)7-W3EYH4&8e4XXJEW;CW61.M
cOg)^TEb,2)[++EH=23.8ST.TA4#9UQ8)PO9GTP?[eT1/\Rf716L<d&UAKO&HTP;
JV,NA/XgXR=Y[eYW0e;U.#,ITI<&Z1CAL>a5f1=DH_I#=fa^W^EKL)FF>BGCfeM[
)e^.#8I_GXBE]e^,UILRG=Cc=_2GA[=J]>9Z8fLOUH&#7&&Dc)XJPS9^N-cU/&B8
S,f#,SF_^<EOQa>#5JSZ0[JS=993N+A837Q)=2>K-TA(>.(E0:(>KOW/L6(6JcCU
0;C=@3OB,RIX6TN<RYPIgZ9a6?.4LRH/O[M[V:9+ZJ.X>E;))^ZfdQ7aI^WYQ?QE
\WT9^CT#;+1#<F>S0<Z<77/3&EQa2DU1@.GF+a6W,DY<D3@@S(:M?[OQ5d@V;\UO
6aGe.(VZ7W+7VN>EC-\gc?7W@;EeBDC@JHZ21B1.]@gD>G#TZ[0bC<b<g_f<@e>2
IC><#DQfBT#daeN&K[[),VfK+394N:GcUQ1<C9LDVG7=E0P;^@:eCLXG_G67+K_:
-H6+7)E#TQ-7[_6<X^2^2<?K6XA3P@9>48YNKOLWW50,-)>YSGR4YJ[BVM0c+Y+3
LF4eH/.N69[6=?f[MdDX&K4db-2[&e+S_6.NZ-b>NBB8#eg:O&gYc)M4E6K2]6DF
baaecD.XFQQGe.b,\:=)ScN]QO\7S=RdPH:C-,b0)PeH@_8/NE\UZ1I+6V?)49GP
/8e8T#7^EMXaEV##bD7I?ZEKG/\a[(M45M3G0798K_bYHFLEX,5FJ1.,JTDTeO&)
cC\EfC,;ES]=-fTSQHc;ZW=Z?]F9C<?1cY_N/eF+WX:b90G+&2O;4<PdEL0LT=bX
,@AM5AKN@eB6)Rc/0_QWM&=IFC\UDE4DF<a8/E60W0H;7P#ZTaN+7bIW.C:f,d5/
O-0HJKd:IRFKUa8EX+Q+6e/W^P:+D-NXGY/RZ:60-=].#UX4X8Tf+U>dD0XR;Q;E
d/-PAfV+Z@7>)2\XF9H>eZHC+6gCMG<Ce40:7IM?^SV(/]R-291g@<TRB+;QCFcb
/HK^cO7Xg\-aVf,_/?WK/>^dd8/SO;FEX4WK2M3a.S-PX7BX=ZAJ?>_]+/SUYQKa
EG2J:N]&Oa@NcP0Bef)@&O:=<_N+=Kf>5I:XJE=M2[FBDA.::E<2a9QY+P)?fFWe
7DV/Ma\YEJ;F?E<OCYLf:2f9V-?XQ7S<44?2^(9CX[F+.B4&7WD0ABAK@LA8=f#X
;E@-aF9.,K;cST]@N_Ud2^cA>bBXTObQ9G18<YfLdC7bAZF9W6#N;JU6M^GfcZc>
LD6LdJUB?8861:<fN8[Q<UDB^^OF&][JNb,MaOgJETGZF.R<O,I-c/J>bN\.-VIW
_?A;F5@X:g^(B/G-NDFFdT2:V[+T^;NCfO)@O=G;CF(d-aKB5R<V)?cVF(CGIH1\
bI^)a)<(KI_X8,/N4W22T]+2C>-I1.D.]V.QUQN@O34I_bGMO2#CHb90\K>QM.5M
#=#2-N\>[Rfac\YFVLfJME9XTafSEPCWA#L5@+H+@;GK@00.6561dV/I7^<)S+^\
^a:b\,B(gA3W2G@DAP:B6Tg=D;4A2ce()d4EKc]YdL7M<^JRW4@J,VM0_bW#(1Ud
HEV&1XTZ76XG7R-QZI<?K:H2G>>>WN2K]T2WdOB,AeBE\\C>C.d3I)U2FT>g^ZKU
2KeJ96K:5cf7C<Z9K\A;dX-gZC].>94SRg\-8d]b8.c^N+OPZF61/bYXS<+HMI#a
LCO3G^^__210]&JS])e>-N(--_EB/\IE?gKXJd.aPH_4\0_01\fWfX;NXB,?W?#^
6XdM2b[>9/I3K@_e7V=GCf[:a0I\,&<1d75EN>TFSS[FB)7_K^T<e@F6(D=JR01H
YGfJ1_E]RS90;):<_c(>_0FF8f0)/I,_9#=bRY7D#<Bc:V(ORAFc5SWX]NQU]/_<
S-?\\.VZ)dc\>7,X@?HUK]YP4.O5_L=,&/4^&7?QWbJ,dNZbVOEb5/);e^](WdA1
0Z?H(MG:Y@5>5a[N4U=Hd^59>&6HBI)J+&c+8Bd?MYH3Z+bV:0fIR&L[D/,cPA.;
:08eN;?0\F(;]f)>/OOda2)c<.#&_B.f&)]RaS?)VPI5HYNWYWbKOLD);]N0TeQU
3M]4eXJ@;]Q1\a+7/I)1@]=3ddWK/6FZ_=IE7\R7^-YfEN2GdfHHF[]Q=b3)CYfH
XCC(<@:D(N?5W[]2.b(-df;YB]d-\E^[IJTR-\K=,JH&4F]]UMMN#O8aOU,]DeS.
F-]MHgeOGW5]((H[R-(662^@;?d)T?]]<-JC@4\1,Z.dbY#&P-:b5T9TK=D7/MaJ
[5(IP(RNU._:V)Oc>eWMH5XHDO90CH3F.F)ZL[T7MZHJ;9[K->?_7I,N&YI&UB[1
1+L2V,2<e(WXf8]dOCN;P#,f082(RB1P99VFJ8c03G+3XUD^([:TZ-=F6)H&TM&8
f8=b)+3KOGHFedgYbP-=P_.=UI@Q<2VPW=7fLVAQ<eC#13b>7I9LLC-_DFIQ->DV
A+EbM\V/E:gC/N7/QTA6g>T/1GKa0(KS]aD2;[XV]0/?f_/SF]1./^)CF8\URJ0_
#64#2F6TN#/T7AbZX4(WE(GFQ=H6WC#WFAB=M3O#e\6M&P)X9(@7R556fLOJIb)2
IH?HK=]6_NA[fAcE;Ia&G91eKRb7CA4Q?^=Of7X3eB.7LYV+,C[=GEHXAB/J#03_
[<HU^@c/[@=A/14N--W5J-=TEID))g\Ia-]Na)[#GU.I@Z>L;b21,:Y?9[)^:#&b
)1e5YOR+6Q/)M+[2ICT]TgZ056G4&Z7-L^N8/VOegX2MLaII^D:/J(Kad.:U.\Yd
V=5<TJa]/==^5Y9V?6PdB>C;9OG]6bd[_f&(:<WQ^LT<@,,57^OTBc@Fc(8e&7D8
@NUV,ZSd)J,SN&&8>\M2IK7,GcLR+EVbKDHK<S^H#SKM6eX/<T-.C#[VfX4Zc_c)
C,@7?V/3F8C_/c.H@:H4GaT,S@P(/TV0RK27;SV]@Y9b\#4;DV,(d8?\36WSDfMJ
;2Q=08^\(T6A<VK[U&/&dWg5^D5e\OLS1XDYM5)\ZOLV#,._V+E]E1ag2a=_00BR
.6J.(:dQ,RKbe=Ac+BY3R&Y4>TH;d<VHCCbMJO7_8WfFA4B/LA=9fL^9FX[XG:6I
7B6T.[9f;^^.V)PHc7#N]ZRC9WJ6a,;H55KJU<<C/f7Z;:a=CJQLS6R@Y&Xf.b:/
<R4@f[V-Y\]UTXg;]FXLR<7D3^3?;NKBP=?be/4XH]3TXY0B>3>-HFAdC\]R92]R
_3E-8S?HBUa_05,?]>I-DH#3AF=@X7I:\H2<4B;XS#@;\/0S9b9[7IERUB7bAIB^
)()(YT&EHX\GId8S8?R6Lc;)c-H4R_1I1=/Ba@X;L46E,C@]XXZgg8(M/&.)5_Wf
BP@^4?9Y&;D5_#7O/a>YOId\G_NR&/Vc8V3<f7?d4IYLYW#1.S>+;.?3)G2R?FX+
^>Q;X\C<_M@dL9HU.PgNLE-O/X7-D519Lc,4Fee?Jce3+PB>E>b+\J4I]Z_UM,XW
Z4@(2.(DV:G=&?,M)&ZAa;2gSFeC78bS0c[3BeW&B8d\\>cK\6XO8D^d]QJcV(#R
9cA8\F_EZHYd4JNY^<Kc/7OJ?Ae[+a?X1W>N2J2[b?:UIWUfI\A,W/(^f9N-,F[d
)=1;gU1[1:9:E09-J<8N&7Q8L&\a)ZAgYH?CF5_=f,.,U#NSVSZ(W;1adDVb3fCK
[(7^YfffK=8476aU.aFA2X0f?)8g4:Y]Sb>JG]3dPWTR3:WM2U_@VIRV7I.V/-J2
9A6U9^Y<7V=#UE<^=]9d(1Ba3N57A<;/Kf@1N#?T=\[fG8GY,V?>@-,4\3,8ATcH
]A.a\=BB^P[0J+HG196L.+DJZQ&B=4I;P_.M1>&DZa/H@HVO_DX>X,&K):V=AOcU
J/5B=Ke#_#:A9a[,9Y1cN#KcbC@-feMKc^6W(<GQ#Y=[SLbQUYU=/,0=Sa456ONM
0WN=[\SW4BW^gZP\WL/e9LC3>,3WF#PDc?G+U1-^H#)>HP;24W[G/a4aZ0gFG8<B
5AS5Bb;>BE^9.aX8KA.L4.<PCR?C.IQb?_W[8fG/O-HX++CP-A&M_^N3[9UJ:D#K
ZS=A\,U>T3#]\05#S-\G]N6Ecf;^EHH-Q7S)dZfF]\^9_:4+PXE@9M\gP0;NOUf:
85=J6#2JN>O/d]/^^&;QG6P4SZ>c]784(6,Nc]S+KN>f9SRcR4c^)^dU5NY@e;(f
Hg)Oc,\,_&)/GeceEVQR8I#FCQQ<5Y:(e[7X^G(<K.=F?dJMFga==59E-MfP3=Lb
K6[g;=7NgC@Z,7UM&LH2EfZUW;FIB,DL)W,]FFHV)PC[(PHGU1C.)#[E4K&YaLIF
+T=MP#bQXFc]WJIVWe52FE:.P8eOF2381@V2-IR=G+b<N9cRXC2OY64?2W3ca^-S
@)?eec57MW&&<C:P90_>d5,^&Ua3>g6X;cG]b/X5U]9+QFY604K36?=O5^LJ]GW3
XgW^4:SCc,XL\,WeLHZe3/M/&,=]6H(>cfc40V#,L@3?,],61,\MA]g>@5:4J]GN
6;[#fF>^0JQ76\&A2M+-)fQROgAf0.g@Z:2JK-NZ79YEQ?K8LNfA9NB@CT]eA#PW
=b)JUc?0a5NdPQ9aO3eP@F_WXI+R\O0?XSZ==EQE6YA.AFWNTJg#0YX@:F:2/6a4
KPH0eb&QO5KUFTV0T:@V7A--/),f:>1H9)bK)F[T=\Of4.dEfP#1d??P\]V&a&:9
d2^U[X9SUHH(6Y4CHKgY3R->R+A0OWbdTWV>/UBV5fC;+9f9+@FKO@8&RF?8E)OE
F32OK,#L,N0O3fA/aASX\gOg941cA]Td<&94Ed,5+QYJRML)WcL<:XScFD_>5eB+
8W\MLc>PL/&bG)VD[EV)D+[-)BLO,N69VaIZ]E9.0QH_4:A[43I]OD\EO[e=C9,\
O=PC[^DV,DZL,S.1[Y>>UTPDfBZ;;#P1Y;B-)cHbF47bFX?N870Q<A:+10<#EZ87
0T/6S8<-:7MJ@CN[_V0:\A&LafO./=<YOa6@[WG\HAM_fS/^\+,GT.#U((2\0A9\
@#D(>K51CQ?P@_cP2Ca:@,C;C=LE,A3R,GIDBW.88AdKUZ3,L&BbSRCT4aJ8G,3H
SI:&Rc7dEE&eN[b#eLKGa-fG7aaH#R/FJ7fD]@Mb-DXXRX3\3+.c5F#8A<cd#gZ_
>g5,JAe9_9^4L49_(JNU2_A7BQ9RTG697_CX;MX[;9X]fKA<5SfJK7[/V9a-JZ8I
\>CM;2Fd5Pf<EO;&)/_PK:-)X2:1=48\5ZKbR6+aAMO-f@M2&B@V,ZgEM&aXW<cO
WO(&6VBRI@N;B-)WMGILOH8[S>XFaeb_BN,5?+cMa2\.ELO\>\16Y=H\=>(2@bdS
,<F2;/dS0,XdEARQBg:^AMUgG(5)<;g&BKK[:_6/F]+XU&_Y2Xc8K6_&T)cPF5-g
AO0QA+0e]HW-61Ge+47gJ:+<?1Q97/=M4ccbbYR2[V?\[gJa8,N>W5cWOV05AB8&
F4<S##AHF4;?_)IaOEV77Ab.78c.Q:LBUJ>4>11^QY=7=44OBc_.d<5JT-77d_\V
b&=eG5^TGXfSHP(#?GW>&JND&DaIHXE&T0KVM?KX=&MgW1[6g_M_TNa?=A<e&AXM
NSAW5F<^D,M)FWX.fVUFbH82)G@1-+;O/)FN4SG:T03W<2D1UHRL9&b),5QK^)+X
@c5Y_S<5J]P1XICc(Y4<ce1T/)JI2@;EI=O^A0,;4AVaA3]5K0D@eD,-D58NBF.d
6=#>\Ye,DQ-@-Y7HP?fF^9/43^42J^[5#/>a,B^dPD-c/-g@1?)8dG&fU@PT//:Q
RJR;85WRV7b,NL+<S+[<T]HbC)T,,NX=YSg99RN6^56@^@d(YF=G&a2G(cVCc3F/
J-4[?A?(,?])T\06g9#,Xd[J?H-A5Hc9XFUcS,:B,D9/NOI9>T6F\^:J4FB\<._Z
.R@/GN&_cT]6/I8a-ZT86Ze]RDC0&cE96^@5C8^\LUN3]/bdNQ>f-Q(P6,T#^\FK
+26SLKb^[-E&&Y13OWdXWM.gR6]IG/K7;_1WE_6)<CJb7Wb^Tf]9fZ(gb3HCBJc)
Wg_7cQ#f7WF,=B(RNL?C?C9g]g#&ZB0LNDP\/Z7=QH&2c(0<]/8BFd2g7Lb^[X7X
J.K&[bbZMKP/.5\Y6f96+=HR16):VaA\c#?7Zc8VfGMDSP5O6<9/)_RNU_N<e088
.B^(e2H\+e+d/>QP1A[9/[cS,J]3-E-=8+SgC&.G/[Y@V4:7]ZeDIX>S9;LJ^.7G
@HZOGdVPIAQ.Z3QffLGb/=O@f061>VYPUX#Ob7&M4/H)O.-/Q:bdHD44SAA1(E2Y
ZT@C5MS+M+Ze&<5&ee>Y->dNf:8dG<&@QY51gU^SegPRU_B3]>Lcac+A:2=O_c2Y
M6D=HGK(SLH7O_G<<7)J4S(;6&?C#D]?3J_3aAFMKcL/->5c\@2OEcT@3>J6UBG2
[+,^ZBW5,6LYK3@,GMKZJ<dN1:J7M4R.^A&77c.1/81I;C<;8D?61f67[0IM@>WD
WVA=LG?A_ddT6)<=])3gaYJ;e/,GPZQ-K8.TRIaF]6XGL3-fW-TVTWUafT<I_XA(
RfCSU@1SK7W;dJA..0/Bf:9f6c&8Z-0,HCS&UM2gIc08.M[dXR0[K=):BZF^Rf=)
EDb,BC90:PP0eH<)Y[2V=S.Y@86BJGLMFKV]fQ(J2C-:HI(>HPBY\Q:)AbTb2JB\
geX[6T5JU.=1S368ARY#++\4-_Wa?2DafKO]A;UI,OX4g&#4\96K?e2JBX<&?O)D
Va\95aIY6M#G@aCS6ZSXc>:)Z6cD>631KFa9eY7\.\?H;;_<7d5B_f#[Z1=/dWHZ
J8+aM5Uc(d9.Q]b&S>]4GRVL)YU&Z/Ca;H_3fK/JQ^a0g87b_&Je;-dY4VFJ,Oa\
46:QF<Z_f:LN.(De-8UHf1+R?6LHb3Xa5AZS(TfMA<(aQ/V^3I(,YO=dDR.#/NPb
(\=C7g0(G:]DJN^P82](38<B=@c7Y+,EYV)&>VS)P0,_209W;?e8/D;3HP]5QRE-
WV8506fYUPHPSABbY(3?.2&_SPRN(V[bG&J/P]J(O]b.R#b0R(O5b]b9>Zf3[5Qb
&D2L0^F7;:YbL[4_fC9Hgae8(#F#]YeU4B^[-(_5.c,(Z9:<Z#;3)DCT(7Q^X^@T
N+HP&@S[P\bG+5K=,Q<7fIF=,(;g#H+dXMfS6CPU+N;;=<L\<gLXDN-VBVNEaE,Z
GV]1VF)?Z;LR\\FQP/<A7fOW(3F49eGKQ==BKOP^FXQ5Oc7QWGRVU:B[6\b]f)d:
L9[+2<AIB2g39-O4<A/ZWC-bc77G(5gYT:W=ZX>VRcaFBOW>ZK7;UL>?6@.Wc9>N
E2Bd^a@T[=U5WH0JEQHc.&Ee:<g.e\,W:HV72;2b.S2C^_8L.QBYZK5\OM=>bT<E
/D[LaXK^SBa-R:6\_UQ1d.NJR+:+dQ3@@KP+93I,,[9RA-<5PBR>&(M&9WY_P>S;
L)bf69.WP3#b8&VFKLgJ@Te\GA4B;[2@9g(QNDZ<3JM=_IF6<:SHZ.A\-6<E8.]C
\9&1F1OU[&U;.ZE>GP93/3.7UE_bU>A2:aEB4Yf7+E&>+&[ZbK<83>Z7>0UG^LH^
_ESX;^.+EX;?&e?1,]#P9;J7<M+A,ZdFZS)-,U-aGUD15+.O,=AZ(a/(gb4Q6@K#
PO>K,9M;bOKTg?FDDeUNfG8R@D\0ZE:IYTe8=W-3N\7H_aEP7[TO(]S<.c^33T5T
e7R2RST(Xe3Agb#V)DS:@CR2]_c&YbD#46ZR24(/QTZCUANXK#(L=GR5FUA5[>g9
4@M>18<+#fH/caD>1CGLUD))bKB3WQG,HX^P1U75&Z8_3aVN=^F:OHK@cJ(]_Y/Y
N1N7H=BUN)G&(I8MUS,=>f^4I0&7-BV-Z^SE.H:5LFRE.V5a7DY[(MW55J4>U)S_
\G8NFHZ\,,b^Y=8O>)^[CgJ&c+Q&#5?Ja4ddAS.N/SA9#MbDe/,CfG]<ASFT25)S
+GbEU<<AW?.;e#,Z[@bdWSa\\;YD(H6HGFP@HT1F\RN9F8a7>IO]_B/b7Dag?aK^
G[g#;4G#[_OdL>OHBQG<5U7Le/f#&\&gLdWJ-15.EK3<Zf<-MFSMAUSFE\RNNK;:
L<Y3JK3dKgeWWLI/Ccga[D_;_TK\U5S_V._)/O9G=0@8B.D\2HLL:fE<=WZW3]?A
Y^Xg0)#NNVXeW3Zc&Ab69)@bb9->H[EMgL)?KIAWBC/,.g/F<;_NA5+;^C7S9P8/
5?K=;Y-LA25[S=Ae94S_WF.)0Wc]1BDTR+_H-6MZ)I/O8[MMgCK<<Dg8P1bR^H[.
J,0KH#+@2-5aPI:^MF<G\)U/4]G9QdXDf4gVHTUZdF79\PUfUCB5(,6IG.75fAA9
Ae)0b?W&FRS(.RLJBP<@S#F,Y/,N)MHZf7NZ\7&=cQ]4;#=56aEQRHRZ&PD,-PYG
@6WSP5(I3Q?aBFLZR1ec?Rd44A,HT)1EGYSOg+\51IDSK=41>aY;S[+,^T3eaWN/
HZ_[@NG829Xg>c/LDFg08P3#RSa/AAFIL[03>\P247egBAcID1d,S6RE1Cdb0NG8
7Og=E]WY_[0NKJI7EOO>3NNUe+cg<7b#c52f2FQGEe=IBJ@LB\;\LfO&#g<I)P&X
NTD#3X3J7T6T=NK=B?C+2[.6TB[+,MZ&3W]W2_W[_@S3cEN^/.+K+3UVO.HR<aaC
Hc5N#7c4.S+((&A8BY(>H(UX1QF&HR0eAb+<D6@:4J>SCBbaS9_>D&f4S7<?DfDK
#[Z]WJ]SgREgNUY);<^Q9JQePd];X@VS51]N+E5MBW<R,,@f=a?@7:ZZM.aKe47U
WOA7T)>.MQRIR\_[.0bAc6=]9N+BYZIe[_AFDP6M8T6@<aLM1]V=e3CW2TGZR@E?
;Z1?CI24VS.=PC-NV8<C0KNTU4.\/&5^c51<cFHG@W4(+(0LBEH3.Wa>d5W&7PcA
G8?_eKFE0cL7,gN9gOXJ;YXe>61MfW,K]33V:?PUM/:TNG206>]V;cUY\O-3(P>,
81>FX>ISD&A]\[RQ\,C)+_)N,.&2WOMQ23MIb:QO)3L4cC+?B7_7OXa(:JXQEX>f
T1//cZ:/E^O^8N?0Y85>S=7Z-(g,/OK78@ZX9LDLAPR_e>2ZcRU;3Jc5U[I5=(>b
+d(M.SL4dS65Cg.@:WP)B^G_O^)PF6\UA@?[bSKIJ_FQ=\:PV;>XSJ<]<O32EMA=
g;MIeN7J.GT<M_5)=@#/<:++N/RHO,Ud],fX?dQ(X2cF1Bac:^0DA.e2OZ647]J:
0Y0QD?[4L\#:<Q&1BU)>C#6^063^\^g0F)IT(IV5ED>3<I?J9ADUJQ,D&7K<aG6d
AC)VT^?.S-WG\R,::X5<bC_a\N+3G[cTU=F=f(bD6LbZWJ>+P+?I4906+,J,>OR(
P-]4](B\4>2:-#d&1?T/LbZ(c.D-)H:+Q@75CbHX>Wb?T3@<E+Dd1Y@YB4JWfG-^
@,RQQ#8.X)IB^:KU)-R801T=^e.99)bGJe<91BEO7KUe<fLCV.J\,O7Xdg4;047&
;Qb)NQ([E@aV&IbC<^EGZ00(;V2H7NLb?,;U4E&9[:Mab96YJ^bA=CQSGK83TN]C
ggT@.]+\PeY2&4[D=^_,=<J\RV]\gR[FNW^86Q1<J:\a?QKZJ2+,H)O[:4&Cb32?
_5B9L^])<Xb>X)6\53f/NaXC^.a=<fQJKDLQ3-GG4dK7]9+>La2-JbF]HbID1a^4
=9[4g+L4A?DXN_V.R&19.BJ,I\;B:7W\Ne^^\9F/U[?84^_@eW_K6)P:]+gS?Gb-
Dbg68.YUF9MTRH/W=7dHQVP0Kff>+EW\3U(I=&:B#SZ4Ne#c#X:LWX^e/K9VUfdX
;R7WdW+DS02Y\@G_:f0SIFO.Hg/NW(C@BI3<]Dfd_8fL_g<&(dB(GABPfIHKQ0QL
T28#9e07@3LX(4Tg,aWW.5SSafF^g#F4=-,Y(V6e8R2fI3TK3b:B9;^3S(e5Se6c
?cTOT]?XKcG\0eY5F1RM>/<M4-dBJSf59L-&a2=&LfEA9Q64?Y+V@R()OGCLZ1>8
&H[N@RY^H?6WB/]&H#YOL.2G9IbD#N.\^61:_LUEYUc[D\F)DLFZa[K8W);?(2GK
-4X8]e;3WcP)2OPXER5P-IQ^-Y(gdNSO+54]eVL=L;X)=Y-F0d/feg9>+a;BVP81
4))>.3FL.1-77E_P;2<IK/K278K&0@8bfgLc18^WbR47VA=FTJLY+g:TA7dRY)8-
PNc0FXa3BKBZJ220EL?)52;feI3TE\X^F0YI?+<WLaIVgH;I8.bH]2T_#]RFFQI2
=T34J+M,X2O/XCO[0<TQ?K,&#)S0fR/1EL.Q4+FLP3.[JPeFFcP8BWKeS)K4GP?&
Ef?R3;cG.UBBTbD9B7XA,4\&=AJVa_;44&\L@RO?]5;SL3e2I>0?(]ZE567HFf3H
gV]U6G38>8GceMcB<<K->-PD^F@Ogb[0Kc12f[<[)IJDeC_#e5FUZgD2[N][Q7M#
(V2gL<SaGODGK08V8?286;MP4Z6Y;MV2]]4YXPfD\:EU3R2)F>L-BBdK/TKO929]
Sf[)0U^gY,2D1.RLJAX@Q]+:&e^eXX/)aY66_EPYRN:ARedgDAXJ)AKe[6(?L_(@
-56&=f[gIdW4#\/8ZWYLUY&LWT+R99>NB;:Q_<@:[^_0f?Tab3S^]A]3)KOQJJ^^
K6ND]#?K1F>5U?FSS&05U]W49>(]+5((]4+##9A(>#@>d/]CR:=c.9I9L0X>QT7=
.U8X-e[VE.P9aQce+VCAJ>L>A])B[S>:X+>_9P4TUK6e+<8-)YWK/I4Y?@9(Ma,b
8\HIa/+[>B>U]4b-6=G]7NaT@)?JFb/E]a4Z8BV.]I@V6+0OQZ6MQ93CZA;@PF0N
2FB3JM39]OR3c;278P]?7VOT/LMIZ01BC(,eN74-BO?YA@;e2>;VR,,[VHE0eb95
ZG3D-^)TUH9RH&U-IH&5V3Z-+dYfYbOfPKH5?AP?:6P]7KQKR2E^#2I^@SIQ7KSM
GNV&S]^^4725C+J,7&Bd-?YZA#.S1AA?>GP4T^T>L:=K?OR5R(bQZF-&5@@-@5d3
S0c)RG3O_IQ^#JSfNW0\/59X?e9AeDPZT^fXd74/NEX,R3:7>-DKKUJg_XI;Q\#+
gRK#Dc/QaUQ\FSa<e(9Ff;Ze_6bN;+-9V^?E=U>g-M02DEeRUQP9^aC?96&R]&a7
J,BY&DT-L+QS;G^OZBFB,5O?F]<=8/IONVJ?b]90]8E6#VE^+V?WYMT-5OZ1+Id:
eb\XCFECBd.:]PFY151eTPN4\df=5eJgDc<_g8G7A5]H(1GUE-^cd1eHL51eeQ3=
?F3KL\S@dP#eH0B,+YRNW^+6?X3GGA/#PfLdRNgUKY9bd&A<d/VgDSe<VVa.A5WB
TNA68<4V]La<<;\^\G_@I_Z3LK+X2U#d^^D@c?]553LL@@CB;N:-E)7fY:5(<PJS
PPbU=&LG5W=9Mg:#PW3g4+SRR=db2(@<aW;S@#H/1H81=2PE1UGd6/0=c;5);>?/
.I=PC_eY.F02PdE=IH-T\=?Q9G):F,?2CC/fUgg=ODK#3I;GF-W/0?AB>)FF#[FC
X5X,:eaW(F(T-C=51DP9JY@B\SHcWINZ>gP>P#[Ud#&f0MMM7b9_>&6M/E;GI+28
JGBZ=0YJa?9:I&]4JR+SWPEdCU5H=R;C6.^77/KE5a=E<bWO^P@BfK[_\Y].b+MC
)=1IZ:8;V:5EH3PP4S;#_EG6X,9.Lc\ZV11W3H>cM=5D-8]^_Zc//,Z@L\_J5/W6
34U2<,&b<MN0J34)7?18)dd_;EYS-IV0.TY672[VH,X4^&#aO<895N=e@^QNVa:E
U41)SZ@+cBd@Z8g69HYG+>_ab#+QI&+9P#H\KP9>KbUM44=RJb-JPO(PXB09BIRG
c/4bdHTgUTDgH@R5;>V2+g\d#MQECZ7+Mbb/bQ0QdD&9TMN1N6--O8a2cF;Q\G^.
0T=^5#c2V&^&aJ;3A=(&=5Z:F_:C\DY_M+_e2K3;(/@S,SFA8=[(:6)IIUa/GBG#
GXZRO:<?)WNO\>B(e((PP&Wb@PE)6g@-I97<__M)^c^GB(UCeSOQa&NR]P55,E&X
/K,T1gHTR_-eRI7J,bZd;3gB/gLWbGHQ\N29IDgcFC?>_=f),3Og<X@[#=XV@VS/
B\dfO458>ePUJ[:2@/LT&FIa<(c@&[:F-IRXO79U1D^FXDA(O0Hfe-?2WLS?S5aE
M0[IgbUU?+D22KAg)\KgCH3QgB>3g:@cL9XP9R.)==5<[;[#ZL[cYD-H=JSe_cM8
DX7DP0LggC;QK@JHD9XC#JYAV-=H[E3>UaE=#5O22P>WRf\B,Q;\VF)K?_7QIWT]
XHFU,V:M_<aV,YbX<c+3(E<AE.MH^R+Y-Z.Y?O@QF94+FYf6eJg35+G][[6YZ8O0
S[fP1AP4^K:7DTSIW\:^;H?dN=P:T5[gV_gbB6YEGU_)db-R)<4cBa?MF8)bdB04
/<9?CL:D-AbJ[V<F9[D)+Y+d_AgB)Ba1:)a<OR^M[XL[WYGV41cUIM?&QO<+VSR7
-6[4A[M@P46D8=[H(WdLg3>737c6+:WARSIV][3:T5MU\[3f(<]E\WL2CO)52865
[>&_g09CUKca3)=&>O[-Yc&8O,C,(JDMKVTP>#I4^;2ZLS87:N^HJ3RI+RH9/2Lf
2cWIYbeOZ4P4.DYafOZ,.&NQ?KgK0H=b=077+[VcD\+CN4J_T1GbfSZI,)Y@E##9
X3PTf=D9f_&I/5LZ5<Za<O6&cK5)3N2+V+CC3X4W?cg+&J,LIB<D^>(M_<Jg8P#O
cDB1^&CUTI92.)N4BS=f.W=W=_DGTQ=69F4BY9]3?MWYJMI#A?e?^EWX0N<<WVA7
W:FG([RL\cF76=?fT-Z\D6I8JQ4^O&D@4F](C@?3Q4QA7C@bK@_PPUEcFBaR&bg<
)-9[DJ76Y5_(64?>c8)ZR]10:=06,=KLYTEF:bR\HZ&USZ/)JPX/H/,DbCe9+/7O
feCLH=\,::#87<+D<(g_fXKUg9dgBCOK+>8#ReLH<U[[))[F+1R-d.0DV\N##93A
H7bWK8?XWBPDJ6/.e@8e7282;Ka8;S&[;<2>Q[gWB5#AXd,O?S]6H[:/610_Udb7
?=,#ATJM^D?(+]WBefCME?30_^B+0?#.^:6[FQ6YgIRQ&Ya_Z163[MNIW]7eEJP3
O1L/-QS]MSF&b8e;I/];1O[M[FIV2Ve(d=Ya1;P][g)Y#d@bK23@&F+V\_91B3[C
-#9M#HgNOMK:V(^[GBH-TBB[[QaLGWLI6/H\W30Y.ce,#9;873+^a/W/ICg@ZRcQ
\G6U<W=FR)[a->HGObd&MTG.Ef1>N[?;Ve;:.f.WFOdDF9LOBSgYS[+X3RN8)W^6
D+c9,0->V(S[PPd7eP7-<Y6H+e^M=NMC?+Pg]39N+4H)#SKN7,SgHMR.gBIGPeGR
^_=W6>PZO8O^NU?VX0,WT.&,R-U6C=f5^eV3EDKbJ</?b:9?4Pd&:DV0)D>T1&0N
eRN&]RARI.\0GDD_CRP,A^<;;:V?LQ4@:GK4(6QD7HKb1[COd37:JLU/Y5+)c9/_
SK:;dcaHMCd9W\<1EV1NU9d1AMQ]/#^0>1e7^JP9)B8C0-5;:-N.Na3.H(R(f0WC
,&[UfL.]RQ4&gWK2M1/RM4=#?8Y^@-OUWdS&(O1_/4XfSTdb.TW_TUYJHDP)66LZ
ZVWSTKK1N]g\._PYT7P?)8#QDRA)[SAN4aA6gIC9cG4J.,XL>L&JN,1N4OP01^:e
W3QLDPQZ#6X2V,e5QDeHVac;?6V=O]]I#9__?S55V;-Ld<MLEdIUb>U#)WV5ARUT
;Q1dVPb73MLbbZO,VYgG),E6&@)dUGP[@EVB](b+31df3Sd.6aEZ)AW?]W4L_#)3
Cce;W5W0H8g@6Z@<;19O09T:T<d.RJ=YN7=;c6=M@\A/4I<_]\]D^G/Y/#32eYc^
=1L(_f\\>H^\S;dN#cXE&D-AgEMAPJG6@Qe6f9?>;;Sa1#?PO9/EWAO#U\\6A-Sf
XO#S/<8f[Ae[QSJH@D(eA=_Z;OI4.@>DVa8/T1eSM9^>&[E]5[7BfA-Bd-+@EP<G
<OSgTX:=8A@_3U:d&D3Y]^f461A6)aT2#QLL?,Tg)0XUe)KCM.0+,D#a,U(:Q\B-
VP=Q&g[FGB4R5K,.YLN+W>A2\WIbD>68SN2&H2]#bL#XI_T?I>\.>8+OXBWSDbMI
LG^5f]>M<\c+_DH?^[;7^X^OE)\UH9f4^,HQaI2G584;_NR6P\5FN=#=(Rg.DI08
3Z\2]4A,@?N9EU6RF&V=N&O8K&dOYOC1Lf:D(J56<bX>FU?Z7<&[(O^IR^cCgX4c
Pgf]0-S+F>P2U^/TaVFM.R@KS1^+cTZ?PSL2FWE]4ZgX2(G./.PdEHK/61,HO<OA
KSUKbH2GEJ.Z?BXG@aP(P(_eWbJUN_M/7F\R18SM37I1_UWb8822[cfB_5\b]2C>
/^@&LW/?3ge9>FN?PWaQ=gTOU]g3C6F8LQLXW-P=+GUM;C.FUbXI.\E9NCN@25c0
[\BUK7T6:/84=VX[QZJ-N=)_.:D#PC3YP<LdUY:#9Zd/bDMF@4\f(Y[5=/U&4X1W
GK]94c3RC30^<5N-@M&ZSK3P+0IE(3V8U=d#5<T8)VVJJ(RcO_W5c02e/=ZV/4?Q
T<PQMT;CW76P6\OK)MLT&#S7B2]R)[LN^c-^Eb?>M0Q/C7TR>X.Y&S(H3SCF;HIc
N)0KN2fTKQe#02#=a37>H-E=@[LZ6O(40RW3)W3g]UMZD@6K+08[c/8Qc7[5B45f
,O\;(f@c,>;J]\Z-CLbR1GSC2[5H&6I^dF2Sd9fdbW^ZZ9[@A5eTLY:9Tf:cF?fR
-IBO/PDXBQDf0@@MY>b&VYMc9WJd4PDS34XC,Z<eDO?BK)LEJ^?[a<Y0f/04-I^X
a^MMeGFNBcXU6WJc<XgHMcL(]a@\[(EJe@&2A>BQK8SL1ddU(#5LXS25\c:(BIcd
SR<CUSNeD^&@.e07-D)JD@Z_dB9b0aTBe5+.eCWIL.dM^/4d1Z7&GEL<)UbFV:&2
5R1;g(S(NQf3:^\a);Td;A,W8P#e);:(#aE+U(.[#[a+^V7T#KQ/,I5bQSdQ2.^J
Cf\g>/WL[[bKd.3#=XBU\IVP\&gc)gLc4,149@\3EF^EB\fLDFFHgD3UJe64D)RU
[?Md.R\F_,5cF7ZODHc/@^<=KW;AS2U-XSC^[-]@.,QEIVV/YF?V8_DA&SUeTQ90
:I]cV-WB2O+8NJ8.Y-JP8/e;,-)[BP[9g.UGU5/-<L1VWM[=5,0f4298]<1(ZDQd
M9L.W#2@?^OD=_QR_Ic4f&a-@\YQTJ0P+9S8)0KTd+:HGZ[,UKUBb]eb:P_N/[d_
1T@7<EJee26F^LJKfKd25OC4A//@,#JI1PbJ29#;RfgY58cP=]A2//1,I5H8V[6-
dZO(2G8-TK2HM>U>E1XI6F:,e^K#&64X0LP53##.&O(E;97eR(aPJ?fdLEb)6&8A
5,gPE#e6ROR8d2DAEDI=:7=&&O=S>\EYfcX7_8-S>AD/&9/9\^AOaB9;<Q;&J@-S
)adAR^5C,LZ5[2MT;Q&1)N)AWHK0)Wgbd\++eH3X+?(aXQLPZ]9;)AfeJDIV/,E+
WYR&RR/M<XV:0U7I//,#VXXUD3@^MH+f8>F44g#=af@WLI.PbW&)NZ)eF46e+JSF
WL53VO)#W,:D_BQ9_B0V<JMf&:g@UA2@eQ^B_T(,_16e@TLU4X),HSJE4]55][4O
Q(87R>UP^FT+YJ7+\Q\;E\d)JA\C+HKRE800ZdTK2a^HC)H93UL&bDWNLT]gO\bU
[W9I&[#:BA_2a.50.<-IP/6I2(A_dTUFYMEYa.7+KPRWAUSTJ[/:H>OZCR,1[3I^
V=O1N(Y9MKC>eSKM[Qb6dN.65MGP[47/cVP9?KAZGd:4\U<:NXa&S8\eQ](ONS0H
IW^VdZ^gPT;6SfS+V>Pb+M3_C4df,7.=c^aP^BZU>HR,OEE:#^E12TW#[P)e3K\:
Bg3JA/Z-G;/A\DKfYY#7Iga2)(DgPYKR2;]Y_1DEEg@)\G6S@B]TG=81#Zb7g1,,
HJ2=XE/]dFCJ1(-g9,BP?c]SSAV>XL\Xd5CeGdAO,d[6N8V)R1Q]3>71B.9K>.G8
BXa[6O;GcYWWSXG7fW39J#-PJ::@f.HcB?ROS[:RG1+:d7Fg:45L=55\Pe,1R[VF
g,P72&R?<Z]<;N57HSXHd@\^gJO52&g@dX&N>:H<YRRY<]WTf@#2M.O4(Xc10F&?
gC7\]#WU?UfC7>^3Z35_WY0W2&@9#TJSEU.<7OS7/H9g/.0CP-UPP(QPBTXEU/Z?
#aPR&XPU)d8T]+B@YA)=:P>YPB-\2Ab0.;=(8=IcCEdMF&DF8:_:C(Y-TTC;EIfc
1KdQ\2Cg8S]]7Fb@F\226,P,;VAY\BH(d4;3EE1dXe>BZO-aKJR[XMEgH13b=;cg
U90(=d,F:7YBST\&6]F<?DY>U;/+[\PA([W)\Z5IY]b<VbZSL5cZV[_GSQ0-ZC)7
E[X[(1IDYK:CG5)e0cR4Vg)H)\F#b/8QA5J807b0&USOQ/Ld=/MO&8d7A82g<22:
)K@JQA<B^IR#cT3I(>R7d:a__g#b0&TQU-6(L12d[@+QX/&MG_&K-,b,E>M)YWEJ
(>Q,a>If-?Q=TM8EHVR&W/TbXCK[,8bd)ZedM/B(@4E+[K2_b4.&Y1+[QY2+X\M5
E7G-^SVYTKK?ZYFSa:OK>34e\f+RgLgB\[>6a.CJB5,X/UX)&)c>4TL4R-BXCHB.
eV+3;VNA+NCJUGYGcBTK.6.5.:-6,KGTHIT(W=M5T,g4&678-=@F&S(:70&(K8;Q
-^YgOBZ[)d6/4-#\P1MQ>44DY,4@3BSIB^SS6<0++\+HcLQ\8Rb(dAP0d[P:.g[e
CA@1NfRHg^R:QG&HfP/b6^E6-PV]_.]J)[,Oa.A&WPEB-0OH206/@Uaaa:9@7,A8
1S022(XEFH_@3cD/B+73\_O[1_cM,=.@,W8[5S[TT.6a#(fSOCfAFgU8K,+)S#Oa
(JUUZ^@90V3aP:(M4U,-MC8:NP3(PI.?E#6@0IZFBG2aQf\>eWf\U^)N4@B^D<J>
7MITYgM,&3K)Ydg+[JB9#@\6D>:ZASbF\QOM_J]8/[)DUJL@NaYMBWCG>5(9#^3:
8G(1g6D#E)VKJWCCLFg<fXAWR4H-U2Uf7ZbOM2]DO^6WYY7.Da+&fJSF>:26B86/
Pa^U3.SA(@BGA2/QBgUUNP+Gdf9VL&3S@@;],Cb]75Tb4#6E@g/K@IBQQa10VQeP
XYW0C(HLA3]18RNYX7-G>4+?2JL6SP^Vea__b6&4E075]0\e9:cQP?04EeYg-LNN
-bfHSSa,.8fC.L+],D+ea15,BI>T2P2f8HQKcQ9P7SR(^4/g4:=&CF)TcJ^MaH<H
UI^<+FF:I(_2^e#3B(7ME_W?D4:Z+B<@Qf@^?^Rg^8IfX_FSJ<Ce8<<_UJ10CgOA
a8.3+Pe7+Y^SFSZKIKF_Y.gWY&HA6KGFDW-[?;&eWD74-97IY^G^EEa)&#,KRfa/
[F,(TMbbI;39.^L&V;&WTQ1FW3-/T&<MecM+b[T5##Q]U,BR)>]7^F]+W6c76+e2
f.a#U@3WS&T.]2AT<8;:d?M3HRR\H_BYgS\H+XeKK_>J=Y)5-0AHCN2G:@/AeY;:
7#,C).+VYgf.SWNf8W]F_2+3IU2#bB4AJG];/N&_0:.>;+8&S)B(cD>D1GG@7Ad-
W4D27ALB3J;DEc(4CdWf80.\/,AC:^]aXDM@We<0,A<S,;NW?#H.NCMga^^/\;5Z
-8M,c)II[JD;1PEW(VJ081PdX1E=L>?RH6N((0[[d&MBcb\&1,bcD<.UQ0gH595Y
Cb_@&=f+^b[d6/<e[CTX;)CL(&BBL^9H@&FCY7=Z,,CA5bSI><(3&1cUY>;GF_aZ
O^g?^J_S:K)We6E)@)P2B)0:+K6<VR>R83d)6(J._QXA-@eCg-aKa?NTaOWV_#76
?C>45IM.,e25dVZ.1CQCLR6Nc\(cC?f4;FA?K;(6\BM0S1bd7U8EAPV]dB&G[K]D
#B.gW[YHa&HegfY2#eF-\P.f:Tf3X&[19S3UFW:[Oe=X3Y@AB4g58Z\d1BdIM.E7
/[0D:@S^HZ(3bLTW(a^FXXG]1:NYC3BML(-#T+?ZMN6L@e&cUQ\CF=VUZ1P2Z@M(
57J-G8;BEB(9PP:2.Z.(KCK&+0H/;0D+45MANR@\e<9gJR8=dFJ8>X7H<8GA.#c4
33.3BXD+.H\e-gaTNFTD.\eW>XO.V<<cG#V,M:K:1WS>ce_BQQ#UaG6TI#_<FTB;
F^?Ue2/1I/(10-BD\./GS_f]4)9RD3a9[F)6-ZgH54Q)P>;),<Vd10._&JOO\I1N
SYL\+0MW;5e;\b(L>;TBT(IWO:W)O5/0NZ8IF)[>140e?,M(JV<>]YD\1R[=&UCL
Qf:b94GYafbN5/1W5f<a?bZe&eUM7g9QJ2,\T,=;=AGQLT(+Wa\#//.?3fVA2Ee+
O@V#]:??XRg.H1S4H&Uc4fI=)D7/?CQ/CWA\/R9+T,]0aKQ&F9A[FCc0VC#FR(/#
fXMJ1=M]a6/_.^/EBV/<G29:HUCYKUD-M\7b>>,B@79B)O:ObH?Q+V5d4[Kg6Q9I
ce=P\GaXB19UaH:VCBQA38/CJg4IIN&6#RC:]2]GN-2dZ6>g\)DEG(_XIZ35_GVK
,/EA&L_MK&1Q:0;<878+DM=O#@1+=AeU-7,O\NQL_O98;R?=.=^Id#gC?32-^J:=
8EV[<0P_a=Se5f.^,Y)-]Ua4Ee;B;SbQMfcX8<=^0R,E<YNcQ6#4#19<RB6fNI,<
-GX<&K5XQe6[6VX,M/F7#Pb2]E[?LG+TeN<7N@=ZF_SgBbP8:d5@L.VSa8E,PPHL
_]1LE(VC6L]/3Ka[Z)d&G\1EMRY)G]5+:ag?#Ub?YIe_=7]-MX2]A&A)Sd]5\gbT
d&EP.=agO-2<P.d,E?\1>cdMG5OP=P16)b+dZO68OIF-c9_0bX-TNT.P^S3ETaB:
&C@gQ/-63E@H+Ub>;AU^38R>K/MLcK+Y?2YUL5bYg#2IHS2JfY.\+>I&3K#db>9M
V50YON);7eH\>>482YP&0K4d56:SX>;4Mfg8+Y?@-U=VcK&7Ba/LO@K4dGRI1<.E
(-,d31B?1]X&fVa4Q?OHB#7JGC;dTJ4ZX\-5\N6EXBLQB9QE4M@=fR(GHN7KRBXe
NP2d9RB-H8_e(a1GGdKJd6,RV<eKCYA.WJDSg+d&c>Ha],NbK-Lb7\&NRLJLSXVE
OHXdO-@E4egX=\E4:S(SDF8@47NM&gDfgbBK\,A-fLQ2g:3cUU>V6#BaD\c7aEL=
Z]I:gQaMI^O.c]:,>dI\_NU#[HDB#ZCW7I+5_H;U5H17>4Ra;N/)6;#e04#),5?H
H1+Ee^Lc,X8[>/RT<7]M1^]LU_:XA.K4387DDeJH\:L\LC?:9FaC&T101GGW>=#b
.9:db=8&:;8U^P>fS&PIP<dZI<QHOfG1f?K@&KJV7P4_6>bVgCH1<4+\cX?88M=a
&6]VHPC1(CQ7S:f?<]X^aLVbKL>+&.7H/>bHg739H7b9YT.]_S:aQ&CF\/Y&(]6>
;YZ=N1P72\,J,E344;[KW0E+&DA#0]dYT&8Y10>&f1=;BbgY5?L\1bLJ=S7ZcO<F
OB#BEc+cgCG^.WdQ?VaX3WNVR?@(QPT72e;d/ac[BZ]eS88I8I2.:D7-4QWcU>CO
/9FPNf_[5B-?:)G[OM&f[W_e5U/A8K_BIH?Sd9Ie-3AX,H:cWB)DZ2VSZ?=G#8S5
N;c]\J=^(1LWXdL/;MVBeN>>J#^_\K?4]Z@5YUcF>SYDM+Z<A7P7/>^99OLLH__A
NFAB,C=3?&0]4Ldg4?_GLXb:g@,#O[9P6AQ#ZPLN:.e7W4H<I123f_HcZBMQIa.W
G<C[:b)D/NfGD=1De>:a#].6&baKB+7\2MYE+c]@Z8+Y,4ME<SAWa5R&ZcI4=U5U
T9UbTK&#He[822XJ/DM[F[XV73+BEM[MFR5>P.=\]UKG0?89YI(T<e^]3Nea)].<
?<ET#S7/K,fU?:bbgc4.?9dV+UaD3W53Sb/@[2@gU_bQ>E2(C(;CA2eeZO<I:Ja#
;H4>H^=A8R4e/.-X,W+OF3PeGF\2=-ZKf1.T\ZS&3>PQ]#3Cg,PA3;54d>HUU>?L
RXE-]e9#f3>,^^LR.HZ;a1_[+<E^BQ<8KNFH;ag1-)H5UP:505YS+;,KT-Ve]X?9
+fW2@+(8b,TH:Q2R20]RASC3B/)fE#3EU3fMJ.Ma&A6<c^L]gH]>f5M<f_CB[e=7
=];Ogc_23\,K)&9OffM9H&JO<<2]<\K+<gA7fRGMdV=NGWRe3=2>>BGdaLDIdXc5
QM:HBE.a,:eLHcL8W1GP^^S75eY81W/O2)(\,W=H[O@1(0a@X^gXOM<3f<20_G\.
)_;/N,3=VaJQYP^V2/^-C?-GKNJ;-fJT4HRCe9eeS?/G_S>QVSM4[IA0&;d8gVL=
Y/@QZfQM6-_N^Ig9Oaf3MFFfB1H0XHG11N_AeO)K>Q3UYU9g/fgc3E[JU1VR7,;B
1)H+f?&E=gK7RTJ<@bVHZ_&?Ic0U_2?D:D53AVHIS?a,L2@S+8&cbM,X/S/>9X43
86F9G;#LW^P0;R(ZQ&eV&[GBcU/VX1SVf]a-;RY28.8N>6BaH_GJ4<M[?fAOCM]b
QbV4,E23a3H[D05cLRDW&[d=O@[ZRQ\bZCF^RP.gJ#>VC[1,0RG85&G81)8-]M>5
.NXYLbGWL@=&aV?C@cD;Nb3O+S;<OD_:JYQOFZS+B@JfH3;ZJ0GbX#gNCN127d2N
>]c<9[e0.1SM(bcV0I>X79;8SKVU)^BI@/YfTW(?G)3Q[&,?:HYQ\RcBf0AT45=+
&;(a(_)=DfW?:/ScHPQUVPZ<Z#RC-WZL70>;+Ad5+=EAMAA_)BE>#[JEQe]J#f8,
aY9C&cg574-IEKb1GB;4)b_UV\E);;f@X;;/<^0@G?f0Z0T7c4b^4;-4\DO2]&K/
ID2Q6476WGK&ec5BRccc]-9c8b4O:L4Ob)V_3,a8;@IUgX=BF.)^0=A2N9YF;e(V
?3UP@MMgJ84eR/HIdeV4e7J#+O3B5c)W83<==I2SW&-=?-4>dD/Q60d))bJ?;R@B
.K:DK[C8NZR_(6[J6XXM6Lc0[gSE4OFA>#;YY]MeDcQ5(>Y_^;,a8b9]WDFdRQ6e
>B@>Z@a]1[9R/0<ed8S\Z?]b,B);:=b;[#EVI]/M69=QTZgF3T:CO<B9\V6#1742
EA2#7;JTH_\C.f?<FDP:Qb:6QUPY5VGGS@74-OeB-O)Z_A83CbeeC<H-Y2D>@#B>
?1G9>1BVRWf]#G.K.,@GUV?,4V7G:FDQKH6UK)Kg5@eYc1IHf=P935dP\^/>F&AZ
8+.=;c5)__5Z+L,G^B[Z<(IZ]a_^1EPDLKK0PN5ID-LcLIGFKG,FBNQZ[[\9U:\c
0:[/<>[58eZg)@fSRMW0BW+I52^UL;R;f1&<9eJ+._f/f(/OHQ5>cK\7H7aHc.O/
>\KRCSfRcK5C?8BeIg>fHe)eD(E?g\4\0(M6^CK^>G))&:5&T\^]VR[/EAX-<ZH1
>9Q=@6g8=d,Pb,+,bNPd=8Z6B3K-]/(:PV5&6;\bLJY&ABRMdPM[^(M#9g;MDb2C
f)@KC#3>CM7dS,N0JQ/A6\+I1;_<41X#7a=KO0RUU30#6B(\E2]/?d(?fO^bOB\:
S2&W3F)+D?\O3EfW.);48FQA<F3\#^,b,9L5H50_a(E,B1A-7AFE&W@UN=(DZF/M
:,YEC.Yc2]8;Ha;1ZM+5,]b@B];1,QR6N[T6eMYc52\:HegURC_D>BQV<6;N/(aL
EHdH)-df,+=L9g:^?+3XAAeS4c]1-7J(/I:U5I77=dKL/G;MbH#L-_#/I^6U0NFg
M^@f?:M9B2>5#KOd4F+@VXCL:Rg>M/gQ_B2)c1c3I\P.OfI6&d\>O_gY(@UN5#=V
3DYJ^.65T/>5;1>15N\,TVR\I0HTeI_:RV.2S1ANTM;MeHT:Y.KN=e+65GU5QK4H
#c(gK\A@VIRbc30(J=MM,2db3Td[GS=W+@N.,LZW;P-JX#8I;b:7-K_&5K3.<=KO
#<33McZ/@PWdO1\-ZGSb;40&#LN(>EN73WEZAX/UQg5JVfPZ_(?]W21Q#+aKDX0(
M)U4HKJ;^#gB2&7YfdEJ(\R07:6=04=F]BNbNBY2NG-3__JLV<2MaO&5+c1CN0GJ
FOYCU-T1D)EK?RL(QZ/,J9D.Tc[H0Xd(4P4ZQ\HQcB_PW,,/.MC?dROM/=^7Z#(-
IcZd(@I_._)G5#e?_eDcF5)f3P9P3[cR>JTEAX[CafGH@.a7AP-;=;^R\JU(N[)A
,SH_DNa+IYSIe^<EZV<<U#Q-[aS]SdP6@,OREMI:-<=U[ed#2,&-)NVNc2@_DR4K
,C\1VKK&(7=M3HK4&TS&SfQ&SOf@AJ>T+(-.];F]1=S__be(a.7J>[f7:7#S+WZC
H?CPHfEc/\HH:4C.CCH>--UVO50[B]c0RP[+H]&8YF[TRPV?]WAEU?&U88QPf@NC
cE<\O7F/42,A)LW1cW=V_\T@?#3ebWK8^;^B;X03@2N^,564/42Yg=[eZ\OV9eJM
XHTT.0RN;V.+]FOUGO1+.,fO2OR/J=PX;\ed;Ma)3N:+@I@67[#,FY[N8XKQ(_9T
?TJ=(88T4X?T>O9BO)9C6AHOK<N\GMX/24-BRVFY;eBY7#\=J4&g0\,DS-Pce[L/
KSf3P\4/f)OK\,0_Y]G1e>GO,^30a8KMW?9F-=F5E@</_Ld):)DFO^f;)HXc&JFH
aDgLH6?UX5=Le/0>OT3g\.0]H@;QXdXEW#ALIb+d<d[4V:IGMb)_8_SWGff5I/d<
SS_+R=f_3?0d6XA?_TY84aed6\@3+d[:^]S/BAP)G2=?MY=<Q;aZM,D:\g6\HZV_
g(RYLFFIQ4;I^_RLEf2ZZdP(/9JfX_X\Pc1a7K)TTQRCM&K/QHRUK@HG,S<2eIQV
NQ\\H2?X8.3:P>bM&^HCYL:SAQ_RYUEeYC/Y,-YB+WU-)HdEKGf=6d@:?OeIUNX6
2#3@89EaV^/R#fQ+,C8KLGHgOTK9TP/-Ka66)MIEc?)WX0eP.FK)b_K/-_b)]YNJ
3[V(g34<PLC4CJ6D8OIY)/V)9:c?=RE1adE24@>_MgdJSU4S+7GM/<@6VUg63=-V
TS1eFBU1Z<?N+K_<:?E9)N_@MOAcF\6,D:P->6&V6UUH>W(U?+BRJF0@5KcYV&\R
c0F6K-\W;H4[.f<X)PZ5Ia3IXe<K@/-c=;Q14:[ac1Z7QMgKES)9R4[If<+R(Q[,
4P4dVQ57GNe#+,-.XIFCL#FfYVIQ]0C9AcFT<WC+Kd9=c8\^G0&3@3_SM8QN0(UB
O.Dc7[RP[C;OA1AGPPGd=a/J:Q<\E2/gVBN4<Id4-\87(GXF@[MM8ZY[W@]]0g&:
AG510EK/EK1BHHLFe;N5F@XNG8Kd6+GXgH]-=M8+:IDVZ=LY0FEEac)BO\-=B++\
@MROGC;Z(3Y)aVKKRdUa?8=G(XKU18#NU>@H#=@:V,H&/XK[Gb]](aVFR.beZ;(V
gQLK##AXg634\d1bB_;AT\e&FJB:K5MbJ5O?[+=g4a)1@bQ\b&7SWE)7MfXGEO0e
bPCLIP&aUeLBMFQae>//J+CW@:+BOg#5A&HBH);[F9EQIC&+<YTe])e]U_ZSO[L=
?eIQ=Y6;VI92R7M11JWELXYa984cZ<9O-F=8S1.ZU@AMEH@cR>AH8=f,C0^3\gK0
WD99ON0NJ]A.39Bb8&PTHB;O3-4[1Eeg.&Gc3:^#D\<4cR8W]Y4^HfU_.OW.2C<U
05/&:YLEMCU:H59&8\-0YG^)Cabg_fD^1WW3IH43gU+1QSV&ADT@+5<JOS.:BZIa
X&bJd\f[Fe-2LcIaWc.;7Lc^H^99FDJ4(Hd-WXZ4HMG=Z[X+MI\X:KO?cR1HF[8/
7)_W\&+3QXA/1PI-d4@S5=G]X(IPJF/KQ_FUR+^=&Y\6JU0+Rd^9Y(/RRR=5dRY#
gBWa;dZWK\@Ig&8Ce;3S4Bdfbf7N=S9Z?ecSCbP)eK)F;CUeR7G\(O:g;Y1&0Y5Q
(Yc2GM:?6RZ^[6NP^B@\fg?2R2[PKK\4[6GE[d&-;&AG+XS+R:_8EFXK-,4)=J5?
HEQ&Ic>g+NLN-#U(ab1SVD,>)2GC)4RG>B3caJ4D<UYJ+SgQ&6=e(LYQ14>GW>:/
MUWf4Ib]#<N<6D,fA>bL0bg[V0d-6;XbNeKS4I1QF^Y;g=>&D(>PO.b&3T)RUT+.
JO3A+;G?c[JPXW<+<OQ.XDAIG[:)KI<;3(Y,&]d:AI,NLZ?fM9KBFYf^G+eaRCPV
5aM)8_9N(R6I_MbD1J@0(CR(b-\K:f57aH/fDHYc\H-f,MR-;2BID0RR/(3R?f2Q
6AI_\08f_\bcDYYBcETD,73e&FK(3/WG+STLILb5KF(c:6982X,&VCSDE^C?cW(I
6Wc9YEaWEd6J04,;26#gB9V_;.6;-<cKf&8=7Z7#7gRL53c3dQ)S+6FEA4V1V919
H)Of8T2&<^Vb<MXf&N19WW8gSY8CbP7Rc-.CDNAYbAJZ?=>2&6<;a0(,\70[DOLN
EJARbB@O;_Q[A7K.]2U69#G>8+[\f^?_HWX:=cNU]?B7H=FI:W,?=&/#W:DV18]^
[B0Ie8c6+]ZTZ)659EKMZXaK;3B].Qd>O.G0G&Ad4DGCCS/=]XK-5^DeF:JeN8/:
39GADQX1-BL==XT.6-V05[\>DG(:G]8I/dJ)@-8?@_CJRA[&FA)g99(91H9P0_SX
<&KJ\#R&MfFVaZLPDb^H454]KH6)4e2OT<01FLb_-61U@WB,cRgQ;/cd7?FPbD.?
?ZPY;DL,J9U#<DAK;T-aYUA?I9VYT8BO6R4(,7/L6<I35O;a#cfMOPUH4FE0aEe+
HN#Z-E@-X7,8[@]E05DQCMFL\C_1&X)V]S\VO>W+SNC[\R?_K61>9/J5D4b=JBE3
][Q-B9b/@?+\.LY_Seb1fX-gRgA=\-?2V3BH:Dd5D[]V_8^JeE6_DT_IA&eeU25-
JF@6MLa_STZ&FX]#cS<.a@f+0E+Ld-(+K2#A>JTc:71S3PC7aeVR.e<ZM&2)cOFd
<#U-)M1C#c(_B3I#f\GdRRH@c[,8[>GQd)Fc>E5(THS>(gKCOd33c>1/+FE\Z<bN
1D,gF2A>9T/<^_a-/C@S3.Eb.L.>HU=fe9I29LS^8Zg[#JHbZTNa=)Ja,aOe>g(Y
6,;LH>+;W5DT(#efa11.&=FUD0Ig2BJ-US=/fF6I5G-d9:GG0\7eM&MHd45TM^[U
MZ_EB&UY#8[Q>]:I2NK/PLfd)FbE1?BE,32^B<1ARcI.QH[->^cJ(T1/QaD<;K(J
>gaLeVbR]ZKDPN?V#=.&d>=;QKZUHVa2.bOC3#>X0PBQgRPIgQ&)2gB+Q6eLRf5Y
(8.:BBL+3Z+3)_482A54VUe3g)=Yb7ZCQ?.cR@H^W_5CHWDNPS67IbLP>I15(gH4
#2W1I<?D.=;.ALZ3c=RBL+L(W^?Kc2LNG)=YL(X\8fJ:I\b9E@93?&d2FW6.QF>6
,&Q-XDJFI@PLJMTcLMO&M@P]ICRJ9CBRI.b&fd@,)M<CBTEZaHP57UOS6>[0M4^4
R-W3&?5?2=N2Y\T(dM]<4D4caG;XRX?VH/&_JfCKD7W6G;^0a6#?6YWg7g)TgU#O
A8M2a1]1\3J@45L-=THaS3O.feZQ85#?()DZ)\d^YS@F(YB?<e0.+HcWE&_XYf<@
g&XO+ICH52W]<2\g;=@]PB[7bXg;A:H;>P+);#>cGY1TZcT_?L(2OMdCOQ:b.[BI
CG:ag7L^5:Q^QU=?a7aX3FV#1dDP#.gA9-08Z>-/-d84^S):<:4E4g]G1.c]VcAg
97eU..T]OC(\O\@aL+f\KHZSN3gVaFZ/1\(^R/U)MCYFEF3;cM^)X.(@MQ<dS\d(
\5YgA=QCGZC<P.DSBIC6_&DX:f-\YbM(YNbL5F;G?Z._=D@7WXg;+B9R3Hc&,X+-
De+YOdf>fD^?[N,0>e;BB)R58=f[P=\9cWa:d#AY6d\c(3bRQG@V6J_3GRU\U(6(
O(2J:Z7f[GWN80U?cYK/&]Bd/efRBQO>dUbU,?,0=SZO(RO.JL(^Z;dK=(V1.YFR
=__?YOPd9E;ecL7Q.ES=UH,b:>7-I+M1;ANH(:0&g7GK<LFaN+H;fd0I7Y_R_BB=
],g1?O6?MBN8Z8U&[ISg()WOO)_NL?Q6K<<D)?JKM^[FfQUZ>(/Oa1cIb\MG[8c_
YC5JcbbE2A]TZO]?ECGH+3+=_:J@V0QN.K1VQ.:d@QX@4Z)MQ/a4KU/&f(_\3g,S
0aE9_N4MG4BJ7^9].Qa8E2@;O[]PMgTa:B@gD8<55f\#V;U-ceUCO#_ZZe+JgUR?
IMR6&ROcFd^1Mf.2G5SD0K;BH6&H5KT_@8[d=+M;.H=<;6QHDbCT&K8?WT\F?L8V
1FOb[76@CKMZ-W^?Q1LI)]JaB8(7aI?&cgA)<HL5,V(a]QQ_;)c2B@fOJFUPGOI+
5TIAac^[_AYC@4EU,c<=GbTc+U@/@,]?=EeI<M/0&&YPTP)6OD28@VD[E?.GZ\BW
-6)#ZKYEK:X]NY0_9/OV_VL[8FJ]g[^E)ETH1=O)efNZQGTR8.,(;TdJb0N/\<IG
PV?9X6J#G^.J)>EK)#92S4^V]F4./8Ie6VIUF9XfU^]/\IAcOX22>?0M^=gV>F+Z
>EcT?=-^PIB9KHf9<-@Q2:X+,GY]1E]T-HNK68YOP&.I@7IUdS(9R(V]1U^@&HWJ
IFGU2C^4A1.,SL9-aPfBG\20#IRTC3TCJ^_3//3^[<c>a\\]@G):8QcYOVK?6Sg:
MN-f&.S,EQe-X[g6)/HZ\?)&GYN_e\==Ne0abf.e4g:WCA/5?b+(5YgZ[Qf2\B)=
^]Z\QeTPS\@>Y5\C9aT@E1A>g;>KcTZf2CDML-.JS75WQ:c2P[R.14)IN/R;KA]0
T1LN;J^b&(@R9@K=:9543S.HaQ]8W7,TFgF1eg,dM47_&BKX;58I9EPO>D50cOFO
^0=a-#&6877NJ/@@9C.Y040[.b9]CW6&6Gb6Re13e/Fc0S:1^XK.BR^/eD>-JI[W
>TE,MF8L:aA;:d]MRZ8B6@E^a3T>F[9A53SX=(AQFLDc?^#V>B3G,S)+2;=S6^(R
+3GMX11UXE/[b2Gb7J@[3Q/J#eDFbWC=02I0^;TMH;)H8.#.?H[2ga05+[\4F]dP
S,_G9,)Fc#P.NR6AY_07MRFdaPL5,86(>cZO:cB/OG_A8&b8)&FG9B^0\TQ8V]JM
4EPZSS\HfK+IdR(^OBaDcB+8B9:T\cW.YF_#.2]=T(T#+4<eVE6=>c^XP75,B\,-
HJ;,T+RD8I5H+CC,J)G-(PAXKTP9MSZ<,5XGAV(Kf,Ig4J>07,JY_.)[&](7e8VA
Mf.LD6BXSKTCP1J)]-2HaD\]cHS9ZbDg<H\OG7DPC/4]2:DM4]FKa>WE2g6)^V@V
OOHXedFWTZ^]g4a?1dN1(Ng.9DI^?=fLQRL9/#cJDQ)^6SW(D=H=N?NXFI,,A+BB
S50_5W-\IQX\a^^;DITJBgU108&eQKJ[B1C0g-XAc3;+KDX,B+5ATU\aGUQ:+0;&
Q3D2JEaWKKMYcIUgRD&fDZNIV5X;H^E6=N6BE/NQ\TZU)9DE5K4HY&:SE;\ggKe-
L+)K6T1a]a[&9W4(&-X#.P6DffLefb\P7C&[0b/PDL>97JZ;QHK_(a-1;9:ZQR]@
]6PK,(RgY<TaTVaUZJZU1a,8C3KWfbH/c(cb##CHEZ21LYb#8<[,93Mf0[6DFRZQ
.JKB(MVG^9WA4^8_K@#cI@#?SYeI6Ne(_d9JEBc1MV)9KEaC&REZ1))E6+Yb8LEZ
0&U;bQMGQ9QXaORLKGFA>VdHW5E@S],G/0fI/A00JHH_K9=L_G7,L4#)=CgaM\1G
#eFJ>Y3H?]9Q,Ab#a,Ta(+WYXUAY.;89S=aL2aIIS2gDYOYI6<95#QBF[H257.21
K_[B5B)dP6Q5T(KZY:)<.G8b9WaO/S;RfQ/HX#Q+(gG@)Oc65@S>NDf^A<NBd.BU
FeK/3[d05<YH.&G>;LO3dcDFaYLg?/JY1W1+^_(2E4EK587/dJfNc&4MPb+:8-.<
4Z3A-)4N=7,Ga;K=ISW^EC6@^IJVV8BN)I^947=c3#-V3_,GF:AUAC(=)G-Vg1f\
.b7\T4V:gI6eVFbQ]/[YcI&HAdUPIS/^93A8+5LCTX_\_5NS7Q0:@=LeXa0JY0K0
d,IJ0PV7IfIA2?DQ,e#&NEfBDGVH^-L0-4E)cD1OWXeKg&UD=O)dEK=J0.dT/NB5
CMfa16gS+_DadX>P>:>Z,::;4W.N12U1G-DEG0,<f6[JRCIX&fEU5XK#E8,?(&Q/
T&>CXI<SfX)Ed4N[&K6Z79515@F)bA,/R2>21][_b8?2Qc(L56STJ2Ea&2<[\FG1
a_La,JD?/>04K=_eUa6.C1AW+B/-BQ;I#E=7UZUX?.,;6&3R;O4:c=N)IBW\f_@.
VUOg@8(1.X?_6FL+ZU..cb\eD1>4F5aHK7(_bc1QgYb4AfQ#8bA]KIG8[\X[:+Aa
RHf-8:YRbM)\a9VZ7KNE?-NK8c-=FY/SE,L57(&d2Z_D[LY,a50\LfZ][&?>6O5^
NWZ7c8ZT+XE>a?8]@PD-KNKB@B+)Y0Z+@b;.?fbd4,Cf2.>+;f_H<]d2_eYL,EK5
Sg,H1]X\Z.#-Y<H_N5,7YcE\eQ^16+gaMJ[+Z,E[?S]#fI(\#:]^LLR^W2VR45<d
L7WOAD(;9\^];JZaS(5@&M:81eBA>eO?#)VKL\7Ve7+W=IU2BTZY(]Kb6;/#XYR?
+N1CaE#KY59Z[?[;]fLdK-^aCKL>IF&>U__):;QYH91M=PWMY5]=0J7QEU<T]^4V
P)6[Z0LAO0Q/KVH]:aPVC1B5A0UT.8>RJA?C[TOEA=<\We8H<Y+)L[Z;M2M5cNM;
VWFBFGG[BfX.5T=;-DVE^+Sac9Z<BR/#A[&5f/ZV,#3XMe/[\<M^YX\EH+CO[MfD
\EeBdP4XXX?6Ye,DK/A3<0YWJaQIZ<+7>73=bg7G8+b3FJ_a^UN6>1J3-J:V3.L<
(#_KE=2;<HX6a7M8FF9gc/<59<07]&.&8daAb.;7c2^SF8c#J/WD37\W9GSN37>+
/LYR?a#_BBCA9WG1VG@F:7>d[E)?[,X+#>+TReV[6bcNe/Pc+WJ&0\?8(9Y;AG,,
5f\,Q&X9][]=MaE8/eC#4QBOWD<7Q-?5[YIb0d.JTWBeH5<XL+X-9cZYGKNSZC>:
+.-C48F3:5FLH8aXEY&TEH[?+CY,WeM[DQ[0RL4W7=R31^=1RJI2\L?ScF=3^2@Y
?cYc86LNSKb)f=NJb?;L\?4<#BPP(g0EdYdW2(?g2LYHD5U-bH[RB8+Xb4RZJ?:[
=:@b;bLN-CPbcd,&bKD8)<-Z)9FVg2d4f3SIJ^JZ9Qd:Gd^Z7DA]b5d6BFJ;a.++
;\0J4Me:YG_Q9&VM_VRS#7DV-Ag74_X^A?dgGXH\0O)a;D@8;cX?-2YMa6F/M1)Z
2^:@&)]JMH[F-)GUa1X?;YI^&>8Ae8[4c5>]aaadIMM3?(VS.f//OI@bZU+)[f1H
R]XU]bdN8;gfA1g=aL]E>#?IIF?[-YDM0@Q(1K)#L.2Y5>.WVA;JPgG#A]E;S.J:
Xg^ZJ8#LTNK(),\:aG<;f^HF8(@)7fHO;22Hd\2IKa<73=S<a=Hc0:@JJ6:JfW@T
/16=M&LGTPL=1;HU-H(2\cCT+#\58V\G37BL-#W]WB5>CZE_W,ZBTQ_3MYM?Zc.7
W\H?g7?V[P4&d75\#IF.@>PQH6/b)5+S-dD>ZF8KBHOY-_1MKdG_UeTIe)RW4Q20
/]_-9SMR8/1EWM6d5_&)=JHDGRQUQ#RBI\/a:6<D-UP9RK2e;b,A]AQXXL7F&9D&
3f]^I&JF\D<;U9d?9FTY+RbTD^1#1N;P^DJ@<GAJZ/H\#?C=NG[6G=HSBTeDQ-,]
b7eZP>:O\a[ac\68E8K_)N8O>Kg._N1PdZ#Efg088#CE\^#W#\QGc5F4;YFX??8+
Ea@c_U8T8[f[LW\?X-9VJHJO4-@2efAKW;/H.S1U..L:6gP5G9fD[Q^_T)HR7#DU
/OYAJG8aHfPP&Y&KMVS<KDWd6V@]D7-\P6>V6>[>J4BR-eGKA7d+8.4C3(Z?;Y6]
dNbGO43e@e\Lb=M+5dH>_1_f0]G;G)GV+[LX+(0N(4-bcOF.]aS(N0XSI^\SY,&B
IDcQ#.-_Z-Vd<K^d=g/(R]SU1WI4Ue4XFOUdAG;^I^B-DD?g,(B#a:PW_MRXgOCC
WHI)->H3Rd/2Y2,\4FgeVf.c-I>0APgZ0H/d9M2C->\^RP(cDAUc:Bd8P\Cf+=T@
WC<;SJ&?9#<G91SIV=^##.4Zc3b=4\-&7W+R@[EEeR#-A\f2Q74/-+,3YT1VTI7P
FX?0cLLRZ@:&Ge0OMZ\:(]-W1\Z=N0W-NH#E;>?ZQ1dF@1G4\A9C6(/3_?2()=6&
2@a2--6=g[T2_+g3YGMW<JR)0VX^GT;(CcS5^PZ-]X/U3?E0#gYG2&KFU/I-fge:
J]+?b7fF1]<:K5BfT0TDK<=\T?1N7VILF\)UA(Z+LRM5a^&g6XWB<,\W]TU?/e]\
GJ:@,;,_O^gFVL(cJNNX.U184fSHgKP=bX2cM7_@FTB;F7<J_L?9NQYCUNJ0a,gB
;f^KRAb4IG/0.8JH2^)R>LS)&RE44ZNQXeNZFB+KDg_L(J[=#Y=XVR^QfFQAO1L#
^-/F@S?RH(N/&7_N4HQ^HKVTTOCQ&.47VeN\Za^^ge)+d;DGb.Wg5M,cPf89@-5B
Q[aZg2K_bT3J8NeUb2?S6G+;),_P?.1XEb0+D0Q((OK.UQZ\[e6(;a/#QP,:bBK_
QcbF^>NAOV(+DU1+=Y[0@]3R-UDB+PK_N,?C#XX&ed<ZZW_[DDX:A0>-c&O1W.65
g^B,(eWZ/?0a@^cE2G2])F(9b2SfS#C,-fN8=)5T<^)87AQgFde\M>g.KP#,]eaS
QBcT(93TV(S]b5CD_XKXTO9dcIBSP2?8cF4]\<eTI=LafM#<M_.A:MHFR<g)J&#Q
0M#;)K.J1abUI=ab0^&:\X=be_PCe^2ADFY;de:P59K-WF\[f[,Z]@TVKd>F>e^d
XeANb^b6SG<,A_abT=Y#GE.-BJ&&^9D5:?&@>eH)O]AC>EZ<)[Q>WI[/0Ue#T>Z1
7H8U#g27Ra7T-23f:JH2VRGEO<fJ@J/=6_Cfd,PVL93\K_LAKc><ZQ3?ZgWR@9B9
Q+U>=OMX7N&KWJ>/1&_4\1\=TL,OJU^16W1b<.U0fOGQF95[E]GS:e5ZPQ2-).V)
BR:c,VQVW[5@Fc5DG^&EU/)E)aPQ_bGJ&>#?0c22SZ3Af28Ee3S&5dWIf)Se+,<C
c5_aW0O-:-4;M&\EGe/16Vc29>+V1aM91Kd?f&SS&Z+RT\W,9(9ePW[VT:]/N,=-
<I_],)^+KOWJ)Y?,E35W@]6F^<9CX>&[R>)E/P#Z;,e,)4#&\XB^8#\Z)HA_a;/=
Jdd>JWU-9(BU=CaV<FQ];T8F#V:aP75Z;CgIO?6QW>4b=^_C@C&R^]VRMe:9AG?:
S/+-+<bJ[[_bSdM-B>0SKGUQY9EY6cLa0Y1NTZQ@L2\8;9Y1>V2S/9-)3MP,(P:Y
:_^af8#<aT9JTCBJ11R+@CU54SaUd@P,[bQ[U6<&2cRY).6/d9.W&:deXVd9Bf_O
SQ0\=UP==+-P9>U=3.II.Ld6Z<DLcC<@L[Q3@3Z]Gce5XE74<_Mdb:SJ4(V)6>0<
5IBN[<@YcDN#b9IfV[PGJ\Z@=3PUY2/OaN&gCQcU1bK7;HQe2.]2DA#?#OS.JE5f
+K1K(@e5DS_2>@BfgNVBH;EUU55?A1#C-_>R^3;/baMQ+ECM6cd+E3CUWSbZJ@KO
@,+?F4ca>dd1M@Fe7C.L\</3I(^&S#;^#a?CR3-)C^Y1FWDZ3aOK(G\2.@8;;<N]
F=Cc1OAZ;-D?,ID-eVP-(AQX8Ce?>5Y);O]cFeU<D>79;gJ:WEgGag&70TgME@)U
b+Vb9S7)NRI1^G+CIdNA^<Za:d8-0QO[J:RX>\>:aVcVXSV1DWa=4a0VJ:UV9-JS
@GUS5LR9<UCR,7Ie(U:ZU5E?X(R#(.0>4_-?->5(J,\fYK8QR#Y4a3f#1G_^_/7N
e#Q(ZOEfgLIL5:Y/[DF@]X2&Jg[+3ZgU>F6(NNZbN?&=gL7B>Z?M\1GAEWcD/<RV
.R&ST7HD1f#O,dD]JLfI/2F_(UWDZ<^(f[@[@^Pg5=VD887\HP^Y?V&H^J\2NJDS
4E9:6g&Q-:FX[E/N5CD6#0b]D_A_cPX?B9JIT6R3aN[ULJJ&:FdeFEa<XJ];e^dW
P01=,TP:\<SBVB]d>>Q7BT9@<=ITV<@(ZJK(7=)NaH>J&.;.Z6&M<OJ2Q?)_.,.@
8&dXcM/1:XN_MI1T7bZdFU#eE_4e59HC)\K=Xc0<fQ?KdbCOQ]GF#U>OOgRf27G3
-JC&F;RO2Q0=\XYDATb(ecU8\ES:<N)9F(G[1AYf(KH>?SE:e88UZ9>M)_7dfP7W
67,E)08JB&DSUOZG_1XJ?.(=(0.5,MPHADOY)D<9G2AfV\M+9&f9^[7#ZKEG)c26
RG&Q9cROAHK)XLb4D\2262T1&++#4M#R1.dS,/Q+QF_F_U8B/)[9\/@KY3>Td.2(
EQH/09TX<+HCf)e<F&<)^NPcWX;W,/.[M_FL[c8]FI6RfQT/3Qaf\46OZ<?KIe:g
4CXcMg;_[UJXJ/IU_IQ\(@(Z(<Q.fCX&gf10aG]8b/;C5&OE=\1ceQ(DM_/4Q5T#
QbW++eHC5085fc2#6+,GVaUa,WRADOcGc2E7U2.DW@d5J8K5T(@U)(J^a\/2U0@,
5-_?T+I4<Kg@13Y8f15@a,6@[D4=V@OUb5:;?PYd#F/Vf[T0D7SD;g=;9=TNd1QX
4XAN;C]@-YAR=()>#]--bKa7K\78Jc@K=Da=L_a)P^FH:AV-9E6EUN&VL;dX)Z^A
e#fL,.DOddP#Z)Q:^&1b?=gNU]4L,)V1S&:.EE1)N/<S8H@@aCQ?YXI2L.>G][+g
.A^T<<gMNNLUN_>@eBBL-Cb_<QeC^4.MDZ2^JT>IE3(gF=#0_Id)8LX]LNSQ/bI2
4P6TCeKfSf1EA:OV@eZA4]A,4D@[Q[Zf7BXI?.=/Q3@_TC6P??B(TN4Y?daKcS?a
M.:LaN:7-#dW]?=RaL83FNK4]9@PL&S(D]U]8:OZ^ALD:e1.)8SQSW/18@W.2cW?
f3134e^&VRe-ET5-dOMA^d_#IR7T>.2HGIcTS6OBSEKNIdJCb1R@/T_=P2dO+50G
E3Y)3C9f(7#Y[GPXJ/7&18_DbYEF>eY^T3GKT0?d#N\4Uf25HgI+-eX8LU+GF8I]
F;;@+2]B+GKABSME<M\[4G2a2eY:_MB;Y;YBH49W^Q/M6bU+__gFNX>ZLE,[@YfB
3JA(3)fg2S&+H=cD#H\B>?PK8gKEO92V4)6BN-@.3WE.fE71L>X/a;5GbDLbF9MV
@:2F0K9BMWV8d>EGa<@6QJ?YN;c5SFcPee>JALMUH/6^?5aXcff@]OR)53F^9f\(
U,e6^4bES,(Za^^&@O;aJfa>f:8]T;_Z_JgXS_O#]#FRW]3WCC2cd>?S=]Ta)=UA
21A)A:6-#9)c0eBO^Gb2/X(+5&Ke7R0I8bTX<E4\JU^?.5V=3;<:ZB[,UT>^FE]U
/Hc7#D#_&[AA47fgPY2^PH[L2M?3.O;RGTDM)XUN<J,^(B+H?F=@\WfeKg0fA\HP
_RcLI<]\]f2B--07&[J2c)-Y_.@U2+N8Pf0E7Sf\W=BSB4M&Qe.[[Yg\05\OZT-D
FaNJ86V5/aFD>;7EeR)4Kd@R-2+H-/bb2/4.(9RDWbd-,RII629>4TXZdeW^O..]
W@Z[]3ODWIC\N5QW;.f]322I[?0Y;+TT2V^+2O.HEE=D=F>#JZ]=.5[SYK:AN>E/
5Q(ef76;Tb__4W#0aSb->cQ<KOFZ^)7d9CRY[Z&9JK_N9)QG;fQ\c@Jb8QR-VPCe
9_-IN^IK\g)Ce[A9B^U^_XJXD)KN@^LR3487&X)FHBRZG]gCWPf:aCU=MCY.U5.+
K^#9O-=f)&#\<V/Sgf;H6,e,Jf,B/He>IT&CKL=AZJGV+X?cg1:dI5dgd_J>C=Z9
=;S[@Ve;HLP[_e6GZE=_;C,5RO[+&KU:K\21:;43D=1NPPJ:[bC=]\<G;^0bg,DL
]3RJ8DaH8Ya0N)0P3FcU,f3AJRY1??ZVQHQ\H>dCL-+:gQCCD/F.bG(TD7gG\EGf
Pf(=.1A&@X(3^O^:7b=UgWP[T<&ZMd1G:f2A-&=B,aQ(XaM9bPFb.IL-QQ@?(__,
-]R]&I<(IC9NS?Tf_+T^]LO)B;=HL+f.K3Y-]YfJP<:@+9&9_9H1+DNT2-M8.S4>
=eV@GTV2,<T+#fd2?SW:>RSIZX5LA:7?9JZBe::1b15RbTNOd#43YSfUYLPO@:)V
MAFP[A6.Z\_Gdb4cSP6NF2cgAH1,.6^9\+ggW-)Ccab>_LN;e>g5C[V=QBfG@Qc]
7^A+N]GWJLURZ>GO+]@^SWeb0X??&?eP<_dV^CO:3bA/:Lc#/MS4V;LW#)R4O^AO
gC4a54K]9=Fe/+<B=@E=:EUbf20=F);fcUFT;eQHe3#A@/]9?aRWFbADbJ.g9[P(
#3??P3&Ue>XKMbI;YaG(E&cU/ZOJ.CG-W@WEM_Y2\PgdC]UP.fRBb<04.HQ4,Ye^
5_GTZ#?K12/\gOG:6W1\FN6G[R-bEZ>DK_@fQa5E?c1H86T>a+ZJXC5W+BM],J3g
eV1<.<G)C/><N?D:M\7=FCZe]<QI42RE.,Pc<2]H]\:/G0#F(Ed<LR>DC++(F)KW
c?/32M\@GGCT])S_Y\EOb=GLKG(M7^;Pa=H]3PE&gX.AVDW>\.SN+N+D@2Q23W2N
6BeE0L>V-0f;I=Y:WP\55Xf0)W09S=3UN>2?d[Hg,AeE.9g6Zg>30RYS@_8)CY=2
>.=R5.4SROS@1gCZ7O]L9MNV)2OaLS)g>/W8MVa24F+K;:T?YY7g^-#I(W2[R1[1
V#,=F&/d6)<J?@Z=51]TgC298\OBcf)f^,UA):.a^Ue31L#X[VJ)6?]T^>POgR4W
N;3/^YQ<OE6;fR9^4E/NCZYM\5YV:HUAdAF3-T<3-)c4Hc@.<,:23&-C[A(?Wa0)
Z5GJGHZab<D)(?Y/NYZP.Nc7:)\XPW>@cWGCYe(Wa4=^)P601H_c:9LcO7:2;AGF
B^Of8S=Q7I<VVE0DYbW_+bT@J]\2Z@?)g@>D^H80BMJ3QR.#,IR02O=@ZC^-<Y/[
C@J[[J>1Y/bd<YZd@bPFN4=#J]&UFIG4-dDVK.(c^01Y0dEY?407AQNe7JG1N]UV
M?Y\CQ@b)CIFF3AIT4WfXf05]c6b,.63I0@IKH(=3JcR.4XceKMZ:RMC=BZb5c82
D\0A00HLec.<NT7IY=I#3\CacUD<&YRf#QJ#THXM+9Wc)<S4RMI43PG3[a?&T[W/
66#?9;CG(==OfK[a412TUad(+\W44)QJ2WSH6@BP-W813D_d_Tc:J^TX/cX?IeSZ
J;BLO/.G&RMP@K(D0:Md&2THd/FbRaJbeY^RF36cD<P]JcG?T;gKY9<O\f]OTbO@
<39JSa:4be(8[@3/5,Zf[cb23\cOT-)[eH+CX@_AO3^V^b3-fOd;;a@^TNSC1)P+
a5]PAQNVFOQRVg9dLg?LDb/Pgd.I3[5Sa,c^&=DW[(4^eU^>L?[-80C0G>S5LcZN
)LOR24.T_EB>[a8&;#XRBLUR2NWE/Xdg^Gb-<^#ccWD_9d>^gFI1_d@FK3fU?NfF
BNDJ?\QL-MD+G2&QUCHg/KLL@#,ABI+baQ_NE@9Z5BO]7IJ;Y,f2RK_J/-,@NVK<
86cCaHb62M6^;_DZ4CT81V^W/=)]]c1dTS??#CCPQJ@;VR9T#,O43e(>W5L#3LH0
K&&c_f@F30b/,L0-Wf@.\QYACFA\<S>9M2YXIEScYe30O+W:&M/d1_#22UHFO,4Y
agg??bRPeS.H^FSYBAFFb\Q7.[4\e<:La+A]>QS4-S<)3<eAHe0DI>a,9&V.d</F
UV0&E_PR.CLC.b&>-MP<<7DG?^/?)N/(3\LSaL(CLA9a+TSF?7I)RY/a0)S10=Sa
&9#4E3bD,N/dOcRb2fIgg88<]S<cG]NXBbSO?O0XO9)N;DY5XC9)OQBYW<d>dLc=
H4)bX2UIPEE682aCRd57Je3Y.GYdLf<e[#Kc-W@99LZY6DVWR;9V7HU\;D1CVRW@
/\4aO#5=HROS?04bJU.H>@D[e;IC^Y(7#1M=>D>bc&8]3[_\[a6;90/1:^R+?H4@
^8;_7>PBX0d7V/BB]0.a=PHNJV-KW6&e(941#P37\)-H)5,[Q81;N2O_1f.J]UT_
.cZg1?4^b0QO5]<<f.L70;>0f)O_D.K54EgbJ/)8WAU;]D4;C0J6K;K&,W1.DAWc
)#W<S9>612^.(WRINb5^Z99f9N8GbP@HDWc#TJd+I51+\XM_L=>;=/1;H/P4Z2de
d&KK(8c-df<+2/KX+4V^YS1ARaDfK6W.,C,2gVPdXg^f.DKHeM6D\]d1>O;.)?gD
egC0.^d8J7T.SI;)E4I-=[d@05@MZ[=NJPaCA\a+\b?X#=]ILJ3FOg3>4OEAM)Ye
fdBD7&-\dgWc@X-4cL=WMJS0RC50G(74[1PK]1VZP2X;Y0-7g4bN6S=QNAN(Z#MG
NB:6fYT80gJ,)#f^BWTcV\WB]PH8IcJ8S,QYLgN[@3PGe7BI(]@aV@BR<bWPUC4d
-35MAV]2FDP),^;F)S3,]@Q,6D2EH>Y3R?NBU>0;1>3)1DR.Q#M_.MOOgOZfRa;(
C?Z(3#BL@:bOe_._e>BQ?fQKd+.W-<Ud&O9M4(@#FL0?;aWAV<SA9J_MF?:\/bV#
8,Sa-VWE-D;5&]\?AaK9Ff<IgNWXE+2SOc6ZK,QAa88Y^IE:S?@V#P,L51Hf3&,[
0/W]UdEVHJZ[IY<7XA<-\I<EBP+>2U^0MdYI06\8+G7>FOV[Q3HNg-_#[.<PPd9N
g4N2cR@=#6?-G&L/V_e-O++6TZ]O++BNc?RF+K]U]/_Gb/[HR=J#.dL4\6).f;.d
?)N-bg-J\eJ++[^ffbQ?]P3N<^AQ1M/f>-#W6&99U,Qc(Qg5/(c:Y4<<QPc<?U3(
cg/VZ;<+I+aRM&,:26]>W\Cg??&/EG-ffW3_<be<Ld#e8687bFeUN5A<&OMa<J&A
\d&8/.LdN0Gc?B[#;a8,08R<.#1ZVHC(QId)S0_70,2LGHAF7Ha)N3X4DZM^6,(?
Y#7)d@d4U#-LI_A@K7)7:X/[GXVF>B>V,[>+3>aFW&0Y4J\U?1FJ5G#cVD.Web7Y
&Bc4Z(YQ:.R^;V?(<g>2GJd\NQ\[R)J2MDLbTXXLIB95Z#7#LN2Z9=YH;MRYV3PT
E+U3)0RJ3+BHVH>TcTEG6U9_b]?fOB7]8H6VW)3R903[PF5L<VaL_/g9OG-:9LUb
(_>cT(Z_HTBN<J&>PB38+&.0,-^DD2@;e=LK\e=)-O\3E+<eM5D(.LX?^[Tg8^T@
-EFZ[ZCc06H<4X\C<Yb8)L=d&_a^Dbd^?#<Af@Dg;g8P\dS/&=RaNfKGKg)/Ta_R
K,^65&):ML77(-S[&A7<_dS6H:Z7QXOU_XeNfNSTQ>]R7Y9EXG.O(1/Y],:V1\1M
@R9?2aRPRILUdId)N]:\>agf.@@0If0_cA:<&b_cbU=e#(:dVcFIVHMAYL?Zd.D\
8ZRPcc.b=HAR9Q7Hg<_UGbQ(AJWBc=-.Jg+M,JUTD:/fWA(d:.,WK>Q\@>Z=FUY_
DPM-R\e.4CZXA5d?efF?M&?.S9D-M)b#]eac8CKA=BW#5D^&8&P763d(eJ(feKCU
;&XSO&?X#+8X#fJ+7,EbF?ZN0@K\dgD)UKY<8,U@eCI6<4U0>PX.\d6;cKMAaH10
U:SdARf,G@R9GOK7>e3TMaZ(+cN7XMUN#\[A7K-#GX<IWQESAMeB[<YA&H;<44->
IXd]&T0-M636_<4XBO_VEQR01<b)U94C><[D07(9.+4=g8(a\#IZ#6DQ>T+g)5b_
E@Ve\@:If](8C=PVC2V#DYT4QN77>L6@fR@/ZfY;e28.d@#bYYE1=S@A1Cc9H?7A
cNCL9FVQdFJ&Fa>2)=F[4JO^]Q;9\0#2U1N8JAUUB0;6/P(7LHQ1\&DXL.1LZ/=d
8B#g3&7WQMa#2;67])REXT+[UKVHJ@&L.7))-<W;c=>7F^V_<G0eLJ6L,_5ML3e\
LHJIcbJPIZC=.TfQI48P-N2XLJ_J783&B27D#LYQ_@fd>JV-=Ma:999>WD^RCEQP
W_/#fdU_A^;VGEKUc_CHJ4J(:A_G-<,d9S5\9<@^f?>cNb&_d\#FGSO?BK3U#6>^
-e_#1@E#Q,QSU8\TB-8R,C/dOK.UWX+.ENP[4_0,44PcE9)Q2C-22F_d@Sb#VdeP
Y3YPA&f<=1eQA&Q2D+2=R;N;d,KOJ?=bJDRUD<EU(I[cHcG+5:D-B95_dK^8A93.
XF02F1VPAae=2?gE[3MYJG7NaL83XR?3fd0?2+.Fa(.O90;YICF05YJ[HQ1)gW6H
_Z.0Z]S]-3]dD]D+IQ7FPcAR7e@&59-UB<]-V7)#6(G@OZLa6L<V6:GJ>2RbJPd8
PD=,2&.eb,3/&cG)FZA[3L3L>?SfIEg(V2A<4g^(\bBU:O+_21JMDMKD1ARRcf)C
N0(NZPEC/@JIcS.BX7(404-,Y(9P4G45,BV_RA)#8c)T5I)/(TNVeP8<0eUM@X9>
M-L3g)^Y+>]S\>#R,eWNH7X_XRdSZ70+&?,\6;\bf7&TM8-C=U,?K^O2ER.gMJT-
[Oa76[fN^&&I8>8NGP@4Y<4SUY:VL+YI=[NOHfQ@1-68BSVdIN(?ZR4?=cHI=6/+
=QHW)^0Q@?KEE)FTNHJ\6^WAYDN]2U<-/.=I+BGQ?OA8]QZ_WDZX\QB?MQW-dO<e
QDE[93X>P(?8U^CV5/TI26Db#aNBd;1e7Wg4U&KB#(2Dc(:1BeMddBY6)H-H04IR
RXV1GSL^4?QN2&A_J#1c[XHS9fUD9<J[:VcAcNcC0aP/TQRgA-PUWP@/7UIdS1([
EgILa#0Y>LY6/P/D6L4a/Q#)?WeJZ2[/OSR?IgK[(]aIQV<FMNE^L>Sb=E_66/J-
GPFWdT\]S1^AQ,>+0CW?+?NZ_1;>OCg(<X[bCO[(bE3gZ4F=GFe:Eaee=JO9+BI^
C:a6/@_HF_6f55d^2@X?.&(N-R<dP?Q5/eWTJQW^]e\0WV@R6X]R=2QXFfLE]AC9
WdI::Z(QVe=:9(^6,/7HYAL#J4O,bc^5=Q.LVb#)bH=I8+gJE(O5QE?b-Z,SPDcU
5R<fPNW:[Q<JS\B<RJ37#AaX03gbRD1F,A8():Lc6I)b08b?-9LO&=>\20>gfd:8
YDdac96HNN8b0E,>5#7X^^ISf?:2,W=4f&RM(eH_,I;9PU@7KJb(?XNSc1cVBfdU
G80Fca[gG0RV/KJEQgQD0?;RQGH=Q,QAW:+-SEWSBCG&-3ZS?6>(4RLG-e#D-5Bd
TK8FT1\@c_b<VQYJ&,H6&3_ffLD-K,]\2=D46bf.3&SH;b7ZD?B-.^&&#A(\--f/
X>_CZK=A7B@^.[KO)ZFYLfd2X?^99F=_E.0<GUDGd/,HS2R[#E;Ya@L7L0VOW[SU
K8\6HMNH69:9_9)gH+<M8WP[KSdd1.&H=8e+I]6Z6\<GOZ8\V^-OHJV&VSC\VXN(
J[D(Pa58<LB;H:3gF=P<8E@^O7SE8:>[8,99)/0@&U6K.E90EA\-(A8GPQVgYP]F
93fbcRdJeQ)NLP@fIb4.bBf46Q44>_?C<OJ?RXZX7B.Q(^2)RaTdWMPFLS_?I@MS
1L2LD/AWC1C_U,?_,)X2.;8aK??X7c&?]Ja[\U[(FED6X+f>(N#1c()6]#NUE2VZ
;Q8Z9fBQM>g#]7aV3H_aS-Y>-+I/AL4@2>L0>TS5&cO)8RPAcAa+7:_BX7SOZ)Jf
DD+@GN[f?Hg-ZKDNG?e6&aEV.9S/#>J(72\7W-SR?YJ:gTG06C_5#+0GN&J8cG?S
WI0U>W9<2O-M4L19];SN):CR&gFX\[a7fe\CXXaa;H>#JF^)1bNa?#O1,7GL^/10
4a?-_2KAG[9-KgGSe0gH<4C3D>3)3=;cI08adP[#_0>?YU..[O_B7+GGVe/&U[CC
.X\9-d(&]B-X&9+7D-7DG&ZaUM;\_DCNK]6X+b.CZ/N[e7WHJ,(gIT=eWG-/CNc9
He&b7I;IMD5.13#9U;9d@=EC+d<e/NMKIJ,DfOMSHAD/>)=g5D:8-4\LDJ<5TTga
:7351K6]/F-9#Z3R6=VYNa+IXUQeT4O>^?AcX9+UCEgg5a,[=b&835YS1]3\[VH>
bYgN/32CCSCZ?LINW<87Laf>U<eKX8>HAG?;WX8Qg:Q8<OLPbRb&AZ==Q>,M.C&3
Le[#LO:8<#bgae\IfR95O&5\YL/>:<D=##_&:VLJ<bf@SPABCLeX<(,F82QQ5IZb
D(IHf+dAF_<+4e-7g;TVUa)_IHEWJc<KbQ&aJQ2GGR1H1]DGAFA.cZbWgXK)XcC/
AQUZM+5Y<E[B4=DWL62Ef?F?D_+IR>0JcBKX3G&eW^XNXbCe57F^f(K/O4]6#OJ/
,GHeQ[2#7f0AC]#P&ZN@M\HObM4M[9=9F3?g2>:,<)+a=F(\NAFFdT/^?1-g_:JI
c+JA_CfS:;UF,\8MFe=K8,9O9fDX+E6Z[fN#:WeQO:L,IO6gDQ/<4/+b-Z8E:01T
VQR.2@Y(2#CB=;A-D0ET;Dc-)J_Hf[VX=RCY[[dbDXTTdX&:cF=L]=_D7(M,ZLb3
JT:HZ/X?X]=SXNU;&^UTcg=T97,1e@O4(TVXdJXH<e)WA5K[BaB/QCc8bcFEP;W#
W@bG6dS8SB\gA:IL1RgR0D62L\4Ke3;3dcT9TY#>5(948\Y6T6QQV?0(,=S:QR4Q
R,[([>W4N2_[+H-EAe);3E\UaU>^f=_[,EKA0-EL)=6fG8f1S_UF#/BPeIVJTWd&
JaO3eU6.e:WXD.Vd2/:/7U=^&OT3MSOd>\DT5IgRRN/T3CZ9WX@IeZ@8IR<PUIDe
dPECBNdJ,1Z0LB/IgG<1V<HK8bL=UY4)\55c6I9^^B=IICI@aL4H70gbbO#+f9(#
F2R\[<-:OP&?DE9C\4;W#+I;2L5]J&(Z[;DA=[A@Z11W,SH/KYP4-P(e7fP:E2\T
9^NSN<SNL?@Q;ZHN#3+2K_CVWWGFE=HL@>CbX0Q1<YMO/3FT.)A4b:+()86CN@5V
YeeY+/RXc=R.^P:IJX3H@_RGfWd^:fNK\M_:NV@F\Ng4BJ<KS7>=:]S.V?QZC]HE
AE@0/A5G5-b:W2>Z&19GRb3QfcbYSSOd91Oa>P\H(TB^7-\>5CY)Ad7R8FaH8.=3
Q&aa@Fe,B3#-];)Y8G0SV1W\S^4E][e5BZ5^W>S>\ENc+/_b/<@M9K420?4BTe/M
V8>^MfRK6>a.O(bHL&&5cRDU9CJG8;L[_FaZbcP/R<_99;JS&/[FR8I5&,3\:S1T
X5geBABW<ZWO5C#?/L@Vg^N7L.f3[E988+d^]J9DZ4EP7.&[.5I#J7S5e4P&[@c&
U^Z+W\[L33TUV<>Cfd#0LfR\aD&<F)I;UBgUTOUd.F;Ge(a.bK43]V,Ob1A5R90Q
QFL_?]8PBN@E6d192+.&_-UIgG^UVRU\^^3WU1^D/A&XgE5W;1[K@g))F10S<abR
cY5;J3I.\RS9:cV=&]K><9G6C&GJ_]J_Q&Z?]>L1O8/ABRSN_&D@XR&AY^/f\X-Q
CP@2CV_M^.\0;U6):4M+&WU?_WG//#>@AebQfa:65bN3XWCJ^C&F0dBGfFE[5[HK
;H2Bb<4:S^1<NP_@.)cZQa2[YYZ6FRK5Q],=^RCW^C]Y<,M_6a;MbMF//cV\WY5:
Y(3S80+bEL(b>W7>eM)98N].Y-XKOXF4CKEK<7BU;aXG6:NKDD]AAUXRWeGA6b<(
=IL>cMG0;U\LVg+RHHde\2DY5)N[E(&a)b:FJRSKCg,)N4W5bC@^=/aZ75RGY)?K
Z^00EG:HYRA:]Y.8FD4W0R4N[XWR=\)\.,@J?R4[5G-[Jf>5/Y&;P.>]_ORW:P19
+8Q_J[NbUX/OK7@\(52E&@O^@OTC87a@?D]I-#a-:R1E2OV\-@DdaRB=T5EC<[PZ
gNTNK6LY20/>>.U4)M#W8BKTZKN3BXfI,>?Rc6#NCR((3cIY[^PHa+69QJDTd5U[
<B_]gZ56_6RfS<L\T+\K(4FJJccJ(<SPI,4JGe::gVe5?b<[JT&9?g<8+ZLbaRD=
5_Z;8U]6@4F20Fc3J_6ZPW&TG:9<]]N>Zd-K19@(R?UaI&<<b8RdYH^]A:KHT)CA
,<X1N2;G/S=782(DMV^F5.6HIJ,?PQEWM0GafU8.d6^7PM#/IeI4W?D+F0CHC3^^
UQb_TMe.ZRIQYL7?:A3_[;#W0Ya-fK3_f20+HZ@1dbS@[;C8Df-SF5f90aDAVX[?
1VH]QCdG]1OR@0S]U:--,S-C?^#;20Y2<:PNUL,_W9R5aF]N72X&URVNcK0_&]>#
63LSUDOg6;7B)&Eb0YIa=f@Y#(1G@dT/gC)SJdTe>:>IYM1I5\=dc:/[W(c0E_D6
PY3b4e,b?2N1LWL1@<#GHO<5W(5=FAW52_gSSEIOcIV5R0LX:UcFg:QY#(-_Y4KO
U8/V)+[XWNBV5OF-[GK_]L=.C,+Q4C<@4VS\9LAATNPH[<IG1,N\KZDeX0)C,+4&
8<IGE9V2>bLMf>?a)WDC>.OT46/F]@M<.9AL3Tg3AK_2D>GEc0SH=QD+dGX\1Z52
R&LYGF20=#KM\N@F:4L6.W6<67-UHZe_4&<6c7ZV(^A9ETZD8<SScIA])&[[;P+=
WE6b,I7)Z\ZdKM(6]1:[1\BO4^VZ]CL24[Ad/cPU+^:<2ZT0#V0T^_7AJf]2gO+8
GPPU#AKI/6.H<=[6PV2A4LcMMX<HQ1<36Ne(/;Rb\Y7=MN8&,YDS&))P&8R-;@c<
c/VI0;WJUIAM?HU5SRB9SKDA@-7SS@:UKMQ(Za(1TMJU@7DXfZ9=Y[TYCCT,_Fc:
d(Def>++(X,75RCCP/]6d-U6K3O,ZMRVa(7#1_A&Z+D;S>H89.:])#>aJ>P[3R+R
1&c9KEMTT@(e9N5]0F[#(R-7I]D6Qb?=@Kbc0=0@N:PN?X+N2bgd>Y?4c]EJ,Y^:
A36PcIZ]MWZD[,c.+Dg=CB_QA\7^HLA_(KU84X5EQd+LcZJ&YECD_Oa1.4Y4A598
fVEAb6<?Md;8IU+98Ne5;\.RA=6DcD#MHCO\H2dQbFbB@c>QO;4T(CHPa;<gK2Xe
a9P(2[gfc/P9L7NR6//LdKN&>=9gB9O/0I6LQR=;Ae#\G#+Sd2:VGD=[W)[(M=#W
Y)&[2c68?ff#O9R6F6b#AfP:NBcB0-f\:?(O2/@T@(Y.(DXOYa[JA3Gf7KT]<\[&
:D4TK_RM5M75Zf-WU3#2fAK_<1KF:O_2VGGSF:S@2N7;?TGcWTDfga4:=b(O#@+,
W[Q9X[E@4:QR-2[aHKQ^+,NP0IX.Hc#WfR.Kc(X[NLQe(+LLAaS).WWNOO-;F;;&
YIX6;FT_4a.E_>5&efcGf)dE==4J2IaTF>ANc5RDJ\MTdKHUY+9-2?LO,F2d,QTI
J-\A;FZQ-R(c^]d7dF>W8FF\):F&E?T50\^Ra5><&YF-BaTE0Z]X8STBb3TWQ9I3
\ZF75Z\).Pc0Cg9HO-K9V/X,<ZFfcZ91X)MH:352J@UZ,Z]bfIb,\D>A?V6__(a_
gXQ,>OBITBcRA?6PT=8R-/8[6SBW@e)Zbc=1>De3+:-fO9KKG0VC8B&MW/]YK&c2
H-I+G5P,P,7P)NZY,6-6DSI\6[>18F6Bf7EP)Rd/C:2OG0)-T?QgD5_3K0KOS+IR
0::H(>=31[a^Be5O^E-Leb^0F0g3SV5HO3.(Ze.?&I@,<,:L1)V^-+/G;>NX5(-,
>T[_Y8?6Xa2D\ZO:VTdf8IK;;:_CeS\3eeZB^#IY\[8,<DDOV9QMg7\4>7b3Z^TK
fOcB;G:5?c0Qb-FVNN_cV(SBWGN2g-D^->ZXTbI4TKHW<RCG_cPIZ3AU&U_Pb@<\
Aa1(PQ;K7e_JT8VM)]fCM.Z?[=[/.S>(XH0+M,eT55<M::WFHQA]0QWH]UE\F?X,
L-8e5J74\dN;&MgWgV#IQ)5=;]6B6af,eAMDRg)+[GPJS(FQ7,Tc@]D3SS9F+)\X
2dBI:EP\FPXgfA>:fYK1]DTAFag1Od,]632&L#..1_dSILBB@d91D<(IM0#:YcXU
&Vg\/=TT\?BC5.@B0:X[=IZR5O)E-T=C8<@KcPSd,TgQ\?#QYCAXZE3Va6ZW8#8B
@aS2^cK^I^3+.NHIc9V3d)Z5S3M\IL/R/<S.:00>(W4/K.SD9(Cd=JQQP2/-AYR/
_CW;L(]@->/GFQ8>H[,dT+\LfZ;F[EbYDgfSeBR6<B>4N[:AfX..BW/7=+f@:]TU
6?HO40RO4=aD8AXTg/+0/1D46/Z@KfFGH=VFbQ:?APTN#dOV)[]P?#\#L2./X\HV
bL#^J]>9RRNV\88L^++/ZG/7HHgGGB-:,_4/#[O(2-[@AWS4OXS^<d/RNKLF6G59
D-E7^+KK.\8e[(FH]e/V/#4_[/G+DbN5_D(3@c&A?T[g86>.d&cXL@CDHV;6XFM2
[+Q?+R//EMeO16+DI^Q3]B)ZEC.6c@((+7WSfD[^LZN-Y9X^_]2/[6I[+KROWgb;
f<g.Z:4)0_7Y(.-e?8_ba:LUPc:GFDKWbDb<&C_D6[Ba^JfOeGAI_]J69A2dPK(2
&B1C=f>Z#MR4[eXI:)>dH5@><^NH;&dJ7X54]eZF?92N5BFFOb[eHb=7./02Nf>K
C]aACJ#5RGL7-@L7.IeF:#M1JQY=U0IGI1JHQJ2OA]-;aUT?ZDO>c6-UQ1B#f11T
43;P3cZeL=d^fC(C2KK-GO6S&O,TM-[Zb=B1C3A[V3Hb/S?V0GXXD0U=[@>]0Q==
()Q#6)]CTU0EK44A)KUAF8JN;:KZVN.4)\VU9)K3T7eX]W;LAgBDVE^^I)PHCBH#
I@18,P,U.eKO<8PF>4\V;<_aM)^M4W+bC>@?B<5@gJS)_WTJgV0.[GBEWL.dc.IJ
<RMH)S8H/g_1THN_0Y=E<gg8?d(SN8SX/ZP:E@4;069:Q8ZRFA,8A8ABS^M^6:KO
:A3KT0E55&T_#U;H\0,HCS<2J2/eCCLcG&^e73PfL[C_L>KIO-bUQSPW/+94XEfe
LQ<F&F\b?T-(HJO@YV2X(&&H)E?HJ<N&a5+1CM^T6C=OdJDMa6#VIcgJ50_TL50F
4:\S(e-QK@WN#A8O[C=T\;J@IA7H=,Gf0+ACJ&(^0XNC4f@NW+LZ>(9QIA3D]fMD
\&3=;IRP0>fd6)+Ug2#L:1XM0;Oab9REH9]&D8ae]f:W^J^4a8=]I<dJ?&&>_a:I
@>4G>G&;dH.RAVeSHT+HcUX78;1V&UIL#-OW/^DV(SVb3QfI1L)96\bfBG9)M3c8
<80?3eX:,g7[;DTf[^e1-P)eX&.=(=_R++b4eB1YL4,d-a,;.I]EKZL7.F+Ac;g9
fg/?>YUU#=^<;2ZAV(?.0P&J5/+DKK.S)a8/bR?^->_T_3[6&R.)42F7HG]8[>-9
R&SeEC:QdO.fM5KJ[RVJA#JGb(/,E;Z5O;)MW3g[JCJY,IV4_/@bc(QF=[DOTc9a
XKYW]&^C@O(?6>ZQIfd#T/J@JB+JUOD+)AGHWKJYdHf53=?(YbG3.;_S&:YCa-c<
@>^1S<^DWe27#V5V8g4a3E-M0(fLOLRd&KACfB4.546#Z/?N?+-JT<2H?fX9ONM>
FS#ED=_-DMKNZS>\EZBMfd&Y)SHC1]2IXT4]0XY2T[a]HB,Q9V)0J^9YL;9SdM1H
4A>[/(P25g9KGZ-@&VHCZY12(T&?)fVOQR<E/H^TQGX6dY,9=XBcG9_&c#S(_eD_
F<D59TPZ+K59V2/^T,2\3c2ed/H=JLY0gED:<:-ODJ?GM0,,cf8MR;3<JWY@&,>+
_Q2BGE8I]dM.4O.H,];d)JcIX<Zc[7R12P&K50=+UE>XV[S#WfNd^^5B\APb9f>g
AR+g_WXOQ8_;&9b4./M?=FVQ5D2-=R4HF6OCHIDVeb0:@Ud3XFQYcG]2J.6\g3_J
T/ec.NfA-;Ua#F7(G1@_b8\:+X-QQ9c+/e#,/^bYa@/)V_:V+MHQe.3cc&:=_e:.
NNa5&1YbY1=cK#f]KZDFW5BQT3,d.TH/.E,VH(,B6\T(Yc6fA2IF]&7+e6ST.Q>L
HZ8P:-E?N?X[,?^6,;FW7\5R&-;M+NObd&_gLY(1IVEa4=V4>10GYCQYDfNY)aBa
F[0]9A\[PN1FYaL9c@bGTNc<dZfagVB1Q47#I6-P^UCFUbC)JfHJ&BQUDbKFL#K3
ZAL/9_REH_TZDbN>0>d=SJZUJccUT<89G//RQ>P.;E91=e;bedCfI0bS^R>=c3B;
FaL_e#6W6>-1B-RS>8?64;TBP<@GG1[.gK+H8(Q2(4H#17Xeb[RCHb>Q[L;]HIIS
GTKD&_C2-H,DXC3L-@+4X+T?9^Cb==A8_#X0G-Q707_7(\MCDYVZ0>JR;@7WW@V^
>(Sb1a.U]@Ob:S^6AEQ0(M3IE6#ZG24513-?=NZP:JL(]&WP9:ba<RZV6J1=We,g
)GaD.IFG?PIM^\aJH#D33>g7E28IY?G^8@VWMYJB##])<\8[0LPg.bc=H=_/AU9E
<W[\=H.[@ZZ?SD3W50-]=SG,-T6/E28ZMY9bMVWef(aIUf(LDQXG-7f\\,(&I\J_
O@/<[53UXNA;)6<>J5=#B&N-.3J]+#E[eLC<I\C=#S-6HW[TK]30)]E8)4aO=T66
1Xf<A_25LO41f?S&/\fKEOXFM^?9H,5U^A#+TGQP.?,O17d)NUQdVM]16f#5\B(f
Ec2c?cXTX-.\Y2DTa^;SgA/GU1b74g1T4)\9@54N;^4-;dc<e3;TP3.H<U].eL/^
@.)fDWQESWeea,F#K3=M@UQ;HEe)g==&eZAe8-cAI9WDK=;C2#\TXD3^CYKQfDSN
^TW1#NaL/1M883bO>1RVT850b+LY2_4VMS]C=JSN<)bF7H4+^M7Y4OL6C52)Jc_7
X2#>SQRW(2>b4\f[a?<0Z9=?M_X=T-PFV;&#SF&fM.gHbfJC8e?C>=#=4[,O<;(O
JE;855E84b:4f)]L.?O@/8+_0]+Aa<f;ZVZ<f1#:NP_J54=Y.F\&^=aKHSI=MJ9P
Z2RNGDALA)2-7[_CQ)S5\.>bB+9OMBf1@R8CQ&K4]P#Sg8F7:>#:gdJT+^0Gg0^=
DD:^3c8WGSJO2aJT>0bBgR(^F5H9^)[M;9/1^^b+<9@_<PD9.T,P^W\T7F3g=6#]
HMSADW&aS4Jb8Y^7Z?0-Zc]Q,,,TU8MN=JU#-\d5)=a2-E>M)JaNRY,+Y4e]@FN_
)FZG63>&GMKIT@c@]31D]708[:,&L;]J/((<D@.dTaGE\.g]DAOB7/<>EZZ2,+#Q
TQ?RgC(Z>^bc9/X0=J5CTQ(B^Y>U7+.5DS_&g@_P>3JV>]MG5:BH@NA+BT,&Y?&F
/HB12_P:F8:cU\FWA,9<3Eef,4.J;A\IfTL4_71OAVVfD8L@0Zb[gbHE8T]O+@B-
Ng\>d>Rge,&#[Y,g>Pe;PVZZ/?VT0X(,NeQ\52:I=KDW45-HD_G.W[SA,VQ8,J1+
T]HR6&C0(LPRG_egKVKd^AEQ/R6bAJN-&76FRN^4L,K:E<\Y3L(:fR7K.a(]/VN+
=KF+M&>F/O[)HP4-X]R.GO6-K]8aeB],:41dJ<I.B@0>1;,_d/J.N6CHM=3(g8B1
[1CMDfSFKK,/LDc-RDHIEIfc14[QIJOOD-_LDF=J&>;N__g\IRL,;V1bY;7B=OCZ
PW(HMB7aHY?K.;<@Ff<B/JZ>)#ScREg1><BJ_V4V/U4TbF@^2S)=4G2D7=^e=Qe4
,PM;g(@0DJ@ET#+CC__N&@Z3)^](83R1_A91K[K_JU=\9:=0>WeY0#T20SA]-LKN
aC^W>D]G/-ZSVJ(Q_MZF:R9^X[S>X4^96Q7&/9>/\b09feEdTJZ1W#A1\PYefBCE
d[EbYN4aUZNd9X=YZ-#<VZAC_WES&Y8(\Q5;cI648[HXCf-I,08>:6OX__U0Y[]B
b0bO6@(N=TE^ca&+B9>DfP;NTbRPc+5BL;]0MZV&B]#,D>_G,a.\\]N7N.85?&Od
+#UG6B^W;a4:/^_@GQB?5G=QAP)ZM,(;6C??aI4L,9-,XEV-WTX5[-LC=Q)YeF\>
JY,LU3ZgBO4(5XXg3F2@^+-MSXJa\b<L&Y,&e5U[0PB>d]9V8c-_5(C>\&^&)2\F
cPf3]]Q>T?:-U:O?ZS#PKWKR30^DD2De^3Vg4=0?R7&b-LB(5UQ]S9Fe&Q\+)MSM
C+6:d3P)JHA=3W&)5K(f,P9EVK:Y,@D\_BF_V^UZ:6F+K&(46A6AYQJKICMC.T/a
<&S+O)gH2TPUc\U=V@L>TF9JU-AG/CY4VWcVDH0>8&LZ?26KJ&fa,Fd61G@\F:TE
[ISP(\9BE9GL.;-KOM1fUe,U@aRQAWfO21<7?^5&(]3bEIBUIP2BY.fMMDFe[J4?
4KfBWF>[]T9cFFJCK2Q@=ZP[]1IcW;c>5IXfFRLfD+[9E\\D)H;0W7gCER4GB/^.
6^TL(8H]>OIYQJV;YfZ?^BVL2S0IdX\TBd;+/Rac&8OP?f:_?M6T\eML?Gg03c&D
<61F2>ZNT3HQIN.#&gZe6)8&MW#)V?8N6RK?ccK,=bZA2_J0[]Y#cc?W+3OO,363
.<B]@3J;=?ggW&BLTS#dQRFJ/PL/]:?GgYPD9(U#@&PDgSb_NW[+W3VMfT)F;I.+
N_(.HK+.-(e4-N-L6<bC3[4gU:=Ud6YJ5fXBP9Bfc,&Lgd7f\=b,()V?/bCBLZ).
BU,A0DM4?PQaL:f\gCH[WWK]gM#b?5DC2B/ZScZdK/J\<@E5N_&a.cXdbZR8X62>
XVb>FBW^.#Z+>,M3Ye@-ZRdc&4VX=CF3[2gD/LT[c^>6Pa(8R8ULKP_AAA5)4K[+
XT.R?0L<\Xee/+?/VE[DIC?YUMcgc<B5\LSIADW>IIg=SCL&1]]H94+,4ac<(4@J
YNVf]P4Md0Rdg)d4Zc<WO31OP_V@OW4QH25,A@DJNP1\2].@b&SU@JbH;=K(#UR^
)T5(:].K/E(:dZ@>49M5deA>.)NIDI\FbSeEU?5A[I/70^Y>@.LAWT=;:]<B->Ge
(OYX\08BAb9bfU>JK/5#efKaXMVO@7U/W>T8Y^EY?OY2?<ZI3PKZC9<-1(O-.6d&
?&9HdMYb@S28FfN3gf\Nb@49:Bd&OLKQ6XXCb\37&&GLLJ][?(;/&ATd[#T115P?
Zb7GK\9gd@,6GH_-7(G-@[QG[:ONW_,VN@e3dRC^O+CP;&N<FYd_7#Q[^HaCV2K3
K(V3&:58S1fY3+1D8X\D?9Ma:]3]M57R0^.FVOJH@^-X@S60BA9aJ-e)6/G+=;8[
=.LS2,]Y8(/A.93G;?-])/0)\158b)TC7M?e5D:(Gd=MQ5f<VYEdBE9XBPK;F#e6
U.S#/;d?b53GN?37V;/LEF6d]Fb9\(CC[,EQSGC6Od:\MCH)FJW3#3:+R0PZ:J@a
V0HY.QST/GHWIM[K6V+#C)cO5c_<T5\.)AZ7.7bO1B-74+TYN-/SW:9&PZU#9OT1
Eb8(&5EI50#YIbRFD-=^4=ZP>e1B94M#U):S9&M04A>3P.NYM@I:U,f_FYQ&)M1g
)2170]M,3RMEaLC..&T.7(8EBe@0LeM6:\5M3S^.:Z>4V40X5KLYVb4bJU6g>b^2
8+Ce>2QRfZ(gcdNQ_bP6UVAC/@[a5aQA+><T#\NVO7b&g<)=Z/e\C;QG3B6VL=cH
>f:?9\=X564-]PO&\UL:7-&M4G4K-_4V;6T6]T>UA/L/().C)32aDC<U.f=[I6F@
]Z[6,_XQE69THe23MR)\HPU2ZZ208W,?3eEVeH6;Z^Ma^D(0c6#B/WLQ.;<-_IYP
<\2QD9SO_#-3AFHPLec?Y+SRa5;\,fU+3c96ZM84EMD2X<IQ,cJU#8,K_/Sg-].@
27JA^4fOb-;LW=b)I6X+_MbX7EeBP?4QCQ#&]]MHZVB+d6VaS/(d61Y>44D3\2-a
@:V\7II3acYBA8D,RY[fa0OPN6_)GW8FQ,JRZ9LY5<?2G[98ZBSA=VVN)]\ZE#b<
8ZR97_L&S3^)BJ-c<_07-/L70/gE60K?=B,1eb27Z9L_)SCW(/?eW4EeV4^2e8(c
I79eQ><2#AeMV1U<?A,e]I@T6-a//#^C?Q[4V>OT\EPVMA<K13&1G>X_gg_?52)&
^(#a;D,\S3)@dT._1Q>M.?:L)-@/_X+3(2).L,I^<0_#=fF0D0[ed]V7R3K>,2(M
64NYcY.NJ846&^L>M4EDdSN?&fA7b&GW=UF&fPYbcQ-.E00[:467R+4DV?RXLe8J
f+d29;7IH-fD81RF:ZbQ3LTHf+TXX:d58cYcUSK\?=df^H7?5_N?483M()2;:+#)
>D0).cY&=L=K\-f]6R]D4T)=e/O=V_56?[a/>-HHT1_aD8^//a#N9Pg^L3S7^R6?
M:>HK4#6\N:3eR.7]7=9d@;,].#153_C2-NSLLTDX)-E32XfCIJQX7P/6aL)\Tg4
O((\AEQ#T([VZ8f]R.REJL/^8c&I8T9^;c(YgK@Q38cZ>1^R>.T8RG(eZbZ3f3X9
^R=Y\Q1IB>X.b#1a7@?Ld<3,/:;g<U_L6C,THH\S<eJ1Z4I7QDf7R_?_&LQP1W=<
43Rab25^@Oc6+?72.QTY104/E7bcQ>=Cg</)?DcX?Dd=XBZC1NJK1c)Z8^8CJ51(
_fN39Pe_QdN6Z:U0:0I?6O_HbV(C]P<1H\Y:<M)(0;FMS2X-BfY>Bd8F<a9WX9UO
@E?f,a\EJ<Aa\>>BaP:b<ER(]IeEYA)RW9T#V-NSJ<N#)8-6)8.\22d7+Q1.gWCE
f>SHQc@J6]gTDN3\aR&R>cJ&F&3Y/8d_R8DXVUQN3S55Tf[QRRK29QH.>b+^R.)[
g.N:C.)6KUF(.gD,.C0BLGgJgg;f)fLc^BeY4f19@0H&L+TG/>7+M/(D8PP[#a4:
5FBJ_(gc?=fJR07B>+KOP+Jb#ZQ2HQXZdHE<.f@1V#)EAd=WAQN##g2c&bU_FTK1
]+dWHMa8@abR@)CIgg9K(,.[05<Y>5<).@[[bQ0/,GK.f7I<E84O\PNgF.:^5<N1
]Mde9TO^H#4PHNAXO#Wa6:C9QSYe53T/;1gG(-21_ad/)NK0VgMUTaS#JB2+gYW#
1T&;?=V6Pf@?D#4?\(gc9)dME1eB52a6/5NM,c4fO-;6&7:Ha=N0ZIV#fYWg9TaG
df]:/:aZHT4<N,G0AL;[U9bdG9#(9K&&[g,Z:J;S/4.W+=,UW^R(]Q@f62-#B@ZF
&486CMA5HKRMBGF2CF0N>9T<^;#fMQJPf/NKg.IIAA@>,H^6XPRUPf&MX.9J<cHX
;\0JQ)Y2U+6\P@f<[?\Cg0M\&S/Gb3LQBCH3L_P4;W6QT-OF3TXTUaeKcK:&.g[G
+b]M[1N>SD?VCX+MB]0\C6;JFU:VBa6_W&-:Y?N1/;ca)(<S\I5AT3SV/86<OK^Q
-0@Z\;68ab/,;HMIDY7DLC+g3O9KdeR/XeQaeS2XbK#52SM6cY?8J/5aM_>6<<43
BCe^D[>@C/X:dg]V[7I53Z3DS7R4?d56)PI@af.TTM,eI_VJBBDP/cYCTIS?IX-B
=@E?#g23DPC3gU#@XE0QH9GbaFO@-c0b3Y3(Y?M__@0T91^41:^R07&C_WS+20\C
bHBQNbD-CQMMX=F0TN61-+4\[&S?6fS#WU&\C?S]/5B>XfgPN(&J3I0K<bH?BUWB
5ES7<D]e1JId(16/LOGR7YJBBN&K6b\7Mg6/#SH7BO4eT0=)bUJAP1EV4A#M81(Y
J3#V@AR(@/MH644E5Od8;b17bQMBTN1Dc&+H(1]66I4S2),+&AW/5e-;B.YdabIS
?/_&FDGYT2L2D(O_+5Pe;(#>+9MTDYW2\X2.=HGf,fMX3b5FXPZM2]F.0)>W;3F;
)CX@be8(^0(afK/eZ=.S=?&M:\PYTFE4cVce0<+H3.^+C);d>0[6e/NKN:JP;O.T
F2@cTKca>T6?T<&3?D^.]FNMgSLRG2@N_S;a3&+GR\gQbL=e151,E&OICIaX+#XI
8g3?]f&\O?K1FU2VJE-KXYEOd^Zg7K_S5e8U?3//2Dedb1V4>.7Y>4FNK;=ODD>/
\M^gb4,HI^Ja;KeM<11aeN@ZN\JDRb_@Caad44RCKJF)eBPKe_8-c:Y^(&(\UL1-
F-1(54fFQX+46<_[9=5.GG=4UVPNQRYM/fS\Se)g_#GMF]L[QSRBcAHXY=G)eEcg
^NBTW+E,46UX,BBf^/SWeE8CGMO:)8Q5^1)5NM6Y6Fd<0-P_C^Wdb(95Q&be:IP,
gJ^W@H2@7#(<:UM;+QSd@5>1G#^FIF)T5-bX&=fg0]5=(T\@dK?&C;=/<A]e>:=6
2U^eUQfFaN\c)9.S)f4XHF/&O7d<DcN+U6eH[?+Z=SP6,M-J)#gOYWA=/6X1N5bX
#I9V.0c^:GA7J^8T@S&00)APEW4bfb.[AR:9EQOEX9a=XKLd#F99dCO1#8,GOI>>
])=fbV@eO]3&e+?7:CK@,R3LQ(K=D1g,NO&IEVL?<67N)=CS7WV(\]W<Nf@5CTcH
eMgBF<99<&D&+<Q?aA_?ZTCR4eBY=.0_^ASa=Rb@@Mf@CFS4>Y]8)GX4B3IBaTf.
-E[FY#]5-O7TVbD&FOE156SDRcD2d)45S@TINRE=-cN>KC_DLa\[\UN:C9\0?W;Y
SgPL./e4KdJb+5^./=4X?);RRD:X<&4,OZTg4,0=T5X>eO^Z_3]2.AVKVZN)QXf:
Ha8K@L,&>;c1/)M5[XU/7YOZ:+R_QI(N0B&HG<MbQD8VZ[+Be]a)A1I76JA,eA7S
Fc>6-SWU.g9(SV^5I0-5AH[E@\\(/\045Q\YK\Gc]\2#=OaLIAE9(La^3R_:PS(=
[M/3=]N5P0bBBe&(#>T,Y)U6eF,I5/a#\HdbS1dBR[7)c,_3QA]]@-2/H7?VV/7b
GN5:ePZAB7.7@9I:08;JNFA8-Z=A?8=0PYK5\G,2;C61.8Z+XREff[>+@F2bMQ/1
+I<g]f1]f5HdBPZRWR/IFg475?gM0^.7EO\<I2geE4&eIX<>6^Na61_K78[\.cT+
FI188,P_c3AfaIWQ7BaQ+=WO0;.WO_>/?04fA;^R\KdSP>Td,]#^8a5-/3XGQ:^(
&GM^_:E3+\S<^bQ?_K4F?/<A(:([<PH3FTNST^E8X3>O^8F.f7af_+Pb+B>129E7
R(6/6.)R;O-N6,4bTO2N>VC-#bbM?12JP;?N1T90c?W9B@>+LXU\CJMf<;3K,DTb
C96ePJB86Fe[J2C<,U0[@Z5E,aZ_D+,V.Q[-P,;0A098C:A=-AES#MA_5HeJ)FJO
U6JE7<GJ,(AUYZQbCM;JZ0>24L\.2V)I-N0I^IBX=8S<XR._<YUNB2>S5b#9Fe51
7dX;>Y&28PP<UWbR_2bZT@2Z]a^N7@Tgd#b&9>J+Q1&=\RC^/X-:?+;(LN,8.B:b
SA[R;)FEY++c<=5Q(3HcDDV/#M>2Z5K9f<Q<7-A_5db;:TK:Rb?P/2dS[6-ER.fI
]6Q/Ag+U-FI=3K&XS82;CG_=+_XZ2EP2.6<<b7e63\KL]XQ^9=gS/2c;8KWQ6f-P
@dRC-LOG]\W0ce9,C:cF#QMFM3?V+g9D-d5QbHA(O?]M;:)>KUd++R.aT4SI/BPX
;efg<PK)B\gc=V/P0UMgC2gJ_.e)bP<)WIKH)9eg4D:6O(fH)/eGS1[gX00R]D#3
4B2UZBTURc/cT=^TGDb?0=fGWN;HNb3cX##DYI-T9N4dD)S_#]GB<K8C&]f>I[M#
5T9K5C\DKR(E0c^5I=dA/>6<3>B=]J1-0^&3f.,INWSf;,Q@(9C<Q^&@A,d64#Qg
E0f:PP8_]C&fgM,bg541Q8Gb)3X?H].EW[)@XMNFVBV\EgKN[8W__##8O5XT7HBf
626(O)RV#<1)&+S--+cV^]2VDL#6e=V8E]>aab(/:Ea63O1R@@X8fGGZ0FN;DbgY
fW\->X\YIbY6g:T+.\+MZWEHL[IF;I,GS(X_W8;KB:43^VVaU#Z+#U@68U^@+V7G
L@DOQ5f^e1&STX]]]56AW)C4F7e<fM(T+Qd<&:\?CFRg[M45Zcf12-0)6ZZVK=>d
0IK14VKKaCTWH4[8VIdcSDR=6Z2WZb?.6)IS&fad:9\#96bN\[I0>O-YRX#/e#AT
FTdcB]JFgZ)c#[)2OKEA[6Q^fYYUMT)2>O)\H0JgF?+V:>HI^@C+):0P,eb0BK2Z
VDfPaeeQ;f3KQE+P9EH35/SKS/Cg9?:[?Q1.R84YT#gTM>Ub6;<Z5d.DO9U#8BI_
)F@K&Z<1+]]e](#+_R,1M@HBP4eS.(GTUDZ^9T>cD0U=[LY]6T4fT0-#/+0@EY28
7>?A8Y=W^X?G]3a19[WR;1+)S<S1XHLSD8D+:EaI]_O0+3G/,+[9fb]DYQE._H.S
5[gW5AA)AC9N1;5eZ[YBa8C+eKf[R7?=BG.4V<>-cM.<ae@,Z>&;7?\HV@A3fBD&
L@VI-ZM_Ac6MNH/4;dXS]JAJ@+cLH.N6SGN+=/>#.QLBdW-F.RCACf@McB6G62NJ
f:=J@4[A#2.c=PJfTdT2\d<&C]8?XRHd:\#&ef4J1,_?af0,;JcXg8.)7XBgbaY\
d#6:X#,bb][,Ia&C\0gD3[0A&JEL7L<RE_I>[\+=\I@+L85J&1R[#/=&YM9Q3GAK
EB(Kc;A6923GW/RCF0DB84;-=_G<[b-bSVR;&(HZ53BeDY^[E7T@XC#7U@0A-5\S
^gRJ-9.S&EUaSAC<9UGP?[=RL5CJ2N,HBcK,0WdTNP,9ROgWKS(5OZB/43^O2^6_
0dTO@cBC^+JgR4R9OH<-CG]GX^6c3bX\+#.,603&f.d,APD))0_IE.=dGX_eS4=Q
IVLgS,-.dS/1CL5eeSRg94OCa;O2((;<4D7Y[c8&WSa&+RfOAdAHTE?DH..P:SJa
=[QQ[]NIg:KES\20L-H/Yd.AaKIE&=1A>P()JGcL0IRD0KeM0L-CgQHU:HR<&gE0
gc1N@3S,&B07;-O&O7:b67Z]U?5-A?5NV6#f;FNIPR;@f[;W+cW.<87V4]&a\/AE
RYfI9Z(0]FP48BTNZ>f=Q^OYaA,15<P;M0RL)-J&7e#.bQ;YV92gYODF1I8/=+d&
;@4.V_P<6?Y#TW@Tb;N;&Kaf6LWGTa#PbGU0gDHVZ970^&fSV(Z^&QL\G-[6(9+D
NL]_Ve[cLU)gJ2Y(URHM9</T6;cZK#dMP#?QSbe60YW+N(XIWDH:>2LO2aUgb.,3
RJU.J,1>3D/+Hb&Ee.[[+TC.=URN(\D6Sc;AMA[ZM;T7J\[&I7?Q._g6gR=0aEOS
T2S8,gO^NDd+a-S&FHUNO(.H^HDJc6AO+J7K6@F7YI-@XC^55K2dZF4g=PAA=M.G
KdLZSKNeIb_5ZO,61EMZ<W^U/>P(7//f;[BPW]KWJ)ONWTgD-RL9,D]J;;4^eRFf
<@28Fb0SJbbccd67PQT)f_WL-/4(:-P\F4AT+b=dS8?X<R>H\3LL1]+NF&c;O#6V
TS3Lf)W\FD&NH7&+a.B]Ue1IOX7,b)IP1WYWIf]#YT(&=S@)bZX@_g&&#3#>&@fS
V<(]=BL(+(CNET#Z704]ID#dPQ@[H\^HeWdR)PG[JY)06>9=ZWa7HEVNI22=WDgV
#/9#<Zd).c;>7GJRL)CL03WB=3_3YDY2OW_=@8a+I6(^5&QCI&6I8R6K>^gB+814
/\(P<aeUHdF^48PO)>N1gIB_LGFf9LMdDT77,7)Y5C-=&9c+W;dS<9-\HH;RQSKC
#D::gcNQ,=adC5TQXY3f7FF?RZ]8L?HI,gDB#GgGaX4N]H2bFB4Z0O-+OR(K&A>O
RO3g.9^>PB/H(U7<(DC,,BHgH+\/.UO:UVd8G?UQ4a\-96(@VeAfFIUICf]V,deJ
bN7CM.\39)C(<NFVREG?G,6ROSDcM:SFY3L[)RF:<[2_c)S+aPOWLdY_ESN<f/&4
;LR[Vb&XIA[JWG>WJ^1R#.c8M[1_G_=+VIe?<(aBDgeb[H<RI3IJ4-@6+=YR?TZP
QQCKgDUYCaRD;RB)bCA]J)=QE.OAYCcI0QNY:;E?L(86E\UbAa;FaL#g5O](,S:>
P[]O_7U8[E@S?fKBdE.HEJR\SB59;6;3)-.K0,;K2dC7+X6II4GJfZ(/]_8:UFN[
NI(V8K],AG,D#Y_/(UX8LKLK@\N?1F5NU(UCgF=FAcC_3?Z1RNW6@fXNO2SY.?Ua
IM=7^BS3<fPL,IST8R@8Q\E&TQT4KQ)J6UTECB4e=QH3,MG1?a#_G@HHOffT#ZHE
P3_#@_W<O@D7EE1S>;[5W=6_c5E,WJ3fU8]P?,EPB8_[Ca(bQE/CQ+1gIdN+-N:F
]W:-/FRZFGC6JA_YV9:b>Z,+B<877FOP[H]5\Y0(cSAe/@:JKNH\\QMP?9VXSDR1
OXRR6K<MI0WOXLCG]\NCW<K+1.7;+]Y5BHUC#(gZTDH8TeKGTgN7Z(;4\3J/?a4;
=SXJ-V,?64WH[62[aDR^ZQ+/BQ9:SeJT9(7,B_2&@--gA\7AS/>M79G@d)NaM2Z4
L+C\08NbLP(\Ig^V&D@,aD-9U.bCIXH#9X(Je8I4gX9YN.VLgc>XY>]\QH.@VHbY
IB9?6=gQ:)Sa8BK=[FD0b)[]SKg4cXEAF+[d?H4Q?cWf>&^bUH0R#?d=;d()aL_d
Y#+8/f<++\3M-[BX2c=<IRJ=;Dc8;\fb]NHKdCgO>B-B-K,:NccCK#\]:?B1@CLY
#7A:@J7M4&agc)VgA&@-cWQ->5a0?aD\[Z)^I:8?&+<[FG5BfXeT]1&?>E#R@.2[
];0G/A7aB9S3NGQPZKB&#,0RIIE,XP5d(fUH0^]#a8]8eFEd=MKJ+13dK,?6W0CF
7(F.#.daKHIPC&2T/:a@JJeSfF7;aC2(KA\a97c#(\eN,E[bMKZ;KU_Q+_NE^4UL
I9S+E9WL7K=[W1).<RBd/2B.ON2J0PPI+IW5T6(gGA:L\^QLEEb?W,NLdN-GOI(;
8eb2W[SLN?MJUcPR6e0-5MZ)WT7-4=QI:];&P3QHUdJ50\B]T0EVOJ.a\[U2#M[&
6_7+Xg<16&;e_T^079;3@P6=bHb<3QH0K8VM&1/=O_e#R;6LN7DfaH&N:=2cU6&?
ZNeIWGZ(UQV61[V0>(XH7(3D4Q2]gUcE3JPEd4QJc42HH?/c?f75(]G:9-942EgR
bQE]EPQF\C[BN^f\:Z\32N._WWg@SfZg+N#=aOGGKW8385c]:fY-99e4LSR<^OUW
J5FJ>2B?61@1HAW4)LJ9>A;XEeb-FC&79M;VQg\2UZAW@@DC9+gVaDO8fI]XX(bc
Ad<\O+OLCW)>85)0g2.@X:+Ca20K-X:/.(3VMSJgg4Z8)[,0LVLGNPK7UG&;<AYX
f5<5TRO>JC(d3;/);MbS_8#d:M@JT=YGY3&P<+P\R[8K0-]^)Q[#N2.+?cWN(<Q:
WWCeBbSVg8<aQTAVMYFB.BHI7>=U3XeM3]/&_[eDGC[c<\,&6B/F7a>16g,.=P;J
QXeW)R:?Xc2F_G52#(I4\L^74_:;fL-:@+GY7Eb([bg.<D>Uf9X/31<4?GLN:#2F
K]U9^g&&&)W<:RHadU@]/)TWf^73c4QH98&[O-S<7Bc.T@1c-RR/?2Z=5LMOe[(L
8#Tb6bQ@_\10,)MV/KNeef&MI#:a-c);-H&4L@.c#:X[f9-(gH?=U,P]^(GH1Va,
HDYBMUQ>&.@4)dVba.NF6Ng6[^1WRgZJTJG_(T=OUJH05\#548A,J9)g]B-f2491
/8O-2M:6Z>;\\[eLQ5J@&93?4^PU(_RIW<)#\((##PJ1(HDcD#MR;#U3\/O+>M];
CJ=&JU90I=6cD5SA\C7g>5;gMKfXFWXc^Y7/A:-/N-=>+/f:H>[RK]?#FeCN.#ND
XDS2(0A@4AFENHE)Z7g=,EDPT8A@gN[ge?e70&W9O2a[Rc2C1BQC/W(Z#OG2-Df,
]<DM)&)6VA59B^P[50)[Ib[\]G=WK\_+@f9K=^(.gVYVaCMP\a.FB8]3g)?c@5Jd
K;DV7M&6FV3+FOFK:ZeW?1L5Zb3Sa]d5ZRJ--T\g2]M>,Ff9]T#(OI;5Z5]W=HWJ
&929?;B0a;S]9W@J_K-I</F@&H_7<ScTaSgJ5:NSKPbZ,/UNJCJC7He70-/<>.UW
.(/YGf42.7S#[CDNfQV8[NffPRQaJ&V<+/)]Ig[\76SO>TKf>24.))Q-@=IM>BKY
SHWIaL8gK2Aa/5,,\[6<dee#AA6?5SC/AI00d.?9I=19<UfbdcE(?B6MYKT<J[X/
L3&=\e/K1VK5I12C.>5]VF3\&C4SE^dVXT+OY&H?TFb^;CW;;E(g3K71g#U:b<MV
X>B1WG3KeaQ?Gfe^aM^BQ,gTSC\:b4A;O1J>HZJf9F\,YOf\Y25G>GSV<0O8XO#b
gCF,3Kf6\^1I21JGL64Z-)/3;+#P4C]1T9H-MEaI(Y&Z2(;WH[QSJ:GbXg^?g3QB
_;8Eb2(0,PZ7VM..^/gS(bZ;gNP+8;[:<TEc\)\H6f=?a+I[:665,X75APN#0-e8
T0]GI^PAJJ^0C?.CLD2X4W:+&UJUQV)J((a]9;3V>9_7:DUY_Z#D]I5OSBL)0b3/
]/a8VK\6D>OcQAT:G6LO8#:;:<@62G-G[/G-JS+GQ@B+RS71JJ<2D51>.CAdfY2X
#TXYc?<d^G,c7V>YTcB5=L+]1:+OM:@S.V:)=U>.VMFRDV8?BbA2dX.@X;^W_<d+
:dLO=Lc?3ce2(XaJY(YcCJE?&<:/95Za2YAOAK^b48+)^b6O:3+T0E(ZJ_>3=#F0
;CgM?CGX&#)?dgO+g-RGK13@CQ1fE;8]d@^?dY7AK5\S9,c\9ZL[ZPagXX?/c)+X
AGa-fM;\Y&:XNf)Fd+S98e-NJ;88_,aU2G=H3?FHg>dA^R&4_ZB^K&#,A,[O(XT,
X:]]64g=?WW<SUB/Q-6,UMK;0<7;6/a.?Fg(0(1(0#RU<IaH.HT5_RB84cR^_GBH
Gb/W+K\?P2dcc-W3OYB0b,A8G1\37VeNFd+W\\14-Zae(B#>4V3:_AQGUR94H+C<
b.NPQF.NHBG@_e@?K8)Zg+OYY1BCeOCN.2-H.dPLe(.bIeN?N[-T?3@(=Z^fBR\c
Q/SMG:ZDVb7ZC_)89B,>=3&)IIQ:Re>7G?.<[WVFgebdL1Y3X30/K+99E(]H]^A;
7cY?:H0K+/ICUP_f1Eb5aOYa/NYROUVMGf,UBgc+7N+TRN4Pc(B&Z@M,[0MO7VgO
OB)PFB^8?A9BD8Y=EGEF.?cZ2[M:JCFS7R\&/W)LM7:.(eA)Xf1>#M]eJW]YRV>I
>8)9cggN3)72EU2.F-N168Od,-9#?/G1NdOT99.?GB2H6TgBZ7LHBGd\bL6N\Z;U
Q+)7Y]d<=PEPYEb89@)D>T)59[#0ba>@TX^9:CJ=Y#F7eZ+b1,+:,S/[\TCe,QA;
Z)3X@Q_)g)4d(<MAGTfX69=W480N0X[fE)VBX[/c[ISb\B&=>IE+6LS#QC,ccI#<
DfWHL=fN-d7e]E<;=bf8I04RM2a[-N@T\=bBS&.98\PU:gO]4I)2HAC<<+1Cc<AX
5DR3&1615(C;;;L;20:OR9?[\S3M29(Y_/U)Mg[3.D\-S3(OV@L4d+_;a44ZgVH9
@XU]THPg)e//=O4HO_YGEHJ;U)/HWdR7B+g]/#B>F]K?J#gZWF])8<[QPgHg/]6J
O\OW,YNC3ZG>B_I8:OA/WOdPL.(cV#2M0S8+\-YUN+\(LUYE<@QOX3\N20He1S35
@CQ5Ld/)N6H504YJ]6e<B[_^I>BAI4DM0]^YJOQCdG?G>[T(&([aL<_Ca/O3d7;K
X@(XN4.GIf]R&4E\7.e0M\f,QK;<1ab2V:[T:>7ND(V&.U=A]gHDdQ?)?WePD7M>
[3SXabaS]W;#R8:IOF,)+K)D8D_618\YFb=6()2.DNef2Qe7bW6FbPc4+UKWV/EB
#ERTC<?cWV_KgVV16OP7FS:)+V3SD?CV1E\SM8#?F>D1YN#AgN9g;[#Ae^;2,GZ6
EbF8,2,PfdNYgGA&&]7Q]GV8@-2=+dg2T3gf\:4P5TcdGc7.1TJT1\(FANK&/.^O
.29AR.2/BcUAD\Zc;I]LAQL7\U>_2RTDg(e8PE]2J^^<^eWA[EE]IU\]8J]#)0KZ
V[-/=g.S])XW&DEAZ:[C3U>cTDa#BJ)U7H1dZFOe5HR\aHZ:^_I[@[L06(c^I9-J
SWcA8GEX?D4aXS@H@U7OXA=c(W?O4GBZE;7_O4,/1ZI5eK.fA3@RMIR^eOY.DNL]
dDW7@O?1W2K2JVX1YcQQR#aV,b7RS0KaUcI0V2=AF3gMd0&JS2(Xe,W7HMTA=@+e
/G7)JCE&.NTUbSbP92R_JZ[LEb78-(,GF(gYG7<6G<R9N<U[gf>,a(e3<O[IBIH<
+bMBDe/>^-<b48Q+Y084T]-G955;;3]K@Q(0A51+AG@.>>0PTfMVgZ7J7HG[23<b
#AH9?We,E-4-(1g&Z8-#(KPg=caBBc/6LG7I>A9_-?)\f//;J<0b+#?]O=:fe.M_
#AQ=Vc1.H=E0dJAgFKM_E,AURA0>C[BEM#6Ie][1UIDE1a-:(E>J[eWgV8EI5NM:
K]Z.JDfcF.5bABV171U_X36Bf[DV>KD[L9d/,>aSXEb9FY(\3e_:HP#bT6fA,A?9
IZOa=OYFV:I/W2Z6E/KQC4,6\4B(WT6-CP41+[aYNOKCIc_+U4A-HU>1Nd(5ZPW3
eU\36@4M-:-Tb2<1KUF\+-D3NZYX^B?)c=#5,S;eSHC<]R(V).g,D9HM/K>SBE59
29R(K[Ta&VD3ZbZJa3)59<PX95>Qf+(Ga.CA1@TR+H<aefdY4W90I@C.S(D<D&5#
P4R5H+V@a0f<2^WO?ON[dP,)DUX#;H@J<Wd4Z@U.Be)g3C3J+S((UN2Q0^<BM6GN
E+<VVI^\AW_Tg>N^S#W[?\4:82WHI)CU);B77J,E:9PVX\8LA9.180OBK81&B\OU
)S2W/@7E49K<GZFda)OW>,e1]YgHBcXCMI#5W<BVYPX8]3Md76.E/QK;=8L\4J+@
WT62QI>;=bRY0Ba?/DKK,)>)2]M8JX\NJ@P83=OL:c6U/_SRg#R0Q8eYT(34#C@X
>BQ>S:L5a/G=5e>dC@]N(VDNAaGXb+EZ;TCXDB\W/e=ad3^R<.BUOfWM?P:>.XSU
e3]_EGd]gA)M.=+)_.A^Kc7_NMd+-:>DcHP[(X4I7eGMJJ()&04.V(EcZV8,P_f<
Z)Y:S]1=L_CUQZWV<WQa@=>1Y(S8:e5Qa-1+^?]K7e8O)^S5Ga1;@,V5bS;E1@DV
CDbZ,/LF0<bI;9-3#:EAVWP:T45H.,#TXZ2^ZK:QU6ZPS&][e:3VXb@=ZC/LV;,3
#_5dQJf\8@B0[N_CC[I>5V3WgF[1a<4Kc)aILbV?,TS)HU]@)Te-O3EBT)=U<U-]
Pf0GA>6^g_17WVD<?9=3.E]YU43Y3/#J.EeQdbS\9-/K/=)QP9+ZC3@]><\)@U(2
?4YeVN1-TVc:D7:FKc8X.>6(0VfSMINfgbG(+P6\8SQ6ZgN+?)/9Y2dGC[#I<C[9
UCd^BSQ-.gC9:+RP(B2;KBSd^H0Ka,Q</>JMGa0X=5]10MM7KM\cQ/^]F6Q4#3,;
VbM6<Y)eRO)0Aba0+O5+4\:43:0g\:COIE5BR)T2Cf\9P9SAQX1459+PZTV288)E
,1&0?_<0;0Nd0(TLTMa6)7V./M#d=9[OB34TaK31+X7M]g_..aRP_a=0X>05M/?H
&OgUL?cOPAYf[S[LMfDPCYZ78C\_2@,D5#a2T2Qf]A9g+c#WC&PO7W.7R.1G_aUX
f4TT<2N172M,c4I=NOQH[(bRLN?W<d\3[[Q\Q6X?)UKX&,g74<ZBOYKf4X2YJ@J^
2E+HHOeT1T2V8&P(+Jb<E-CK\Qe+U&7O<Fd;g8Vd2L7TDNW#+;0<<Fa3Eg>H3T[S
Zb)IbZ)K@[@V7^;QQYfQB<A#2DM0)f]&5?(VC-dT=BN_F6-ZF.7gF<ccGJ=g?V.-
aB>ba[CA+,Z_K>=BCbV[AFN@4\Q0=5@&OKL4,bfT+0\(CPC,ZV=g,H@NLD@7?/VC
RR0KZ,0;EMc0697\@WH1\G6BVQd#=VPeQ^:^I_(IQeL/,d9J,_BZ425+C[6_[XWT
&PUc@&?U3C_;_g<ANd2DO3HU(ZN52eW(6E/PUBAcb;T\#(Z_<],DQIN_1X:c#V@Q
@V>.^1a8R1,AdBA87>X\eU)?]C:,YEYPC>R#f-3/KLTYTSfZYA:8)ggZ<1]<=:(=
MEa_G&:_-+J9&,d&(Je^7R-I]1>>6>+5N42\SO@#UN#+[R5UO]>F\A^:99QDfKUC
7Od-]E<#/)9cCX^:E:GXZ:Q.SbR_<eQ/NQ?BO6?.)aMF6e(N&H5ZfNE90cZWdBa<
.)2Y<8GRe?HWcJ5f]Oe33J>>8#SCXG-\QaU?Q+(];O><<4)?:S8ZOR#+eTC>bQ)0
HU4Y7<YTU@4aZSdE@J^6LSUZ(U<[SOM8#a_Ca0]V@C=(A+61gQOdQ(H3-F;XFBWg
[SJ/IOcaZ,L>]XbNBCPLW5cNe-A61bI.CL:ZT1RXHH-Sb#IKAUT/@=.?Rf@9W=3R
[f@W7LBZbOL1<F/9YNN<6S@EX^N-eSB</OCA?\@]J1OSBZNLDWJ+O5dIC(I2@WZ8
b^>6MHdV2T(-IN-@C5-]cB^(7^]EI1Mb;&SAB6./-L\#AaeUa6OK(@<gPFCFG6d3
P>E0O&\77J)PcSaQ)DSa89&Z)>0eReDYBE-RYEe:d9[<#UBd#\FWY?CLGGU9T#R-
:dAP0(C&=S5LeCLgZg:?XUg8.KCQ(RT.,S_c+_Id#-PNfO0+b=+?J.H)J85<)(0)
+_0ec^88,281RdWDc-A3;D.8),6D@b+ZI.471P39)0,&9d:NMZMd?Q3Pg7Q1:MLS
)L;/QE\0KK_7JY;[G=[]<cK#0g;4RXf-I1bS8GKP;P5be41^YEcb=.;6PUGX0&5#
)&Z:G+^QSc)<V.)FZK(-c@/Q+Y4]&+Y.gE9Wff>#>^NbfP0/NW,\>H(,C_/H]<^Q
/1=0]T^6/25b)aTWOUOKP2a@2Hf2IF/e+RH>]=,e)BDcT<d12(e)=\:@eDCPPCIN
d963GJ<)Z&?ZXYR>5a[5EM1=f)7Z70V1QWcOQI:TE\\Q+[;G6VZ\W4SW@3NIKIAJ
R^@WC,[B+/;\WQf=,[b=^_>M,3<bM(0>48>FBD]]03fbKG_W2DX8.Ae/8&_=74Sd
@SaKHVIXKMNcb/.XcbJgNfOYdROb[g7\;:LES>#+<?:E3(;U4b+V[KILT>TH\\;)
@T?9Y4:9#_&f/D>(R@ZIcU?K1]9KIJI?U#IS];b[V=,-2XG.c_P53OFDa[ca;SX;
YE,EW8\]];c[J-:F;^?d9G0J;V<F.G:A7A5bcU;G6K3Q=@a\MBI&1KdD0(GB8<0c
a[Jb]3ZOTaKb/@9_=UdPcQ]RG1<Sf4a_VT.)@NXb74Z2?TQ4,>:+5(J\K=+JGZII
S[85E8X^[K>:C&OO3L:L+X:)>;D-C+=;6=.ZTeM35#E/^.1/fTWZ)(<V=LI@b.52
g^J^b]@:^0OCf#WF8:R,.2(H/.;(Z.W_]d1I/IX\6T]<L,0>cW]Q=(CP0@E#?e^G
_)J0K[.FA#\A[EW0TA2IWJg^4\XO(V9VLQb8XC9]85]KCP]B?(NOEf;\O?AT&HZT
)ZT4=KLK:(XHb7KMF=_Ja;D(X,4&#MX]NJA_,:>E_d=5+e\7Ic(BLA+7d@FS:9-6
LeT-X7^,Ua\?Rg-P,CCTTC87L\4O);>,ZX\7/U-Q)JF2=@7GX8)9CcF>&G+W(g2f
\&,g2H[PZ7Hb9&(Y,W<AFFWc5YT8V89X0RY(-d.e^6SX)(WVU;@]3TGSc5H](GUK
3@0)d-_#V\(g>IO5>I.Na]MHGg:YM:2XU<02@6&QJG[<11,TgOEDWCbKd<5]F9-+
ecaMQRJX7U=3#Q<G8TZH)+dA/,_6T?(A/N\TS+g-[L(XWgKc,b8X(fF[eCHD.;=\
H1.e98&-<&.(968O,E\FENTWZC/#CZ&V+7:S-YHcc,L>4YLcJMR(6DTVOI0>M]:H
W&Q+=5:\YCU7YQ#=gcKPHc[++3YBJaX.B=9GX&4934f2@,O^4LgN,cFBJGL8<<Zd
8(G.<D-a42YSUO9++9f-HX=3=_<(VGO)\63:;55^9#TLU7>Zc,KaJ\#Y)CWM-4:^
E6P)UHb]IdJ2g)eY]W>)8PP@.IBN&J4\R9#?\_]]K;2P:THOTKF_D1_1a?I@CCb2
6;_4e\6ISD+M-[XO&KCMI<8+baX:QVJFd.V(6fB@?K[0[2>E[dKBK[:BW=+0-<J-
R;gA(8R29T+NJ)Ge(@IPRGPB#ETeZ)-[)f=,)E@752/Y8fcI1bJ[(@U\d-D9OdBE
JN^]LbHB?4H9_WE0GX<9><WaA>66SUX5.W96?106=7B&e^;587.UPM3YP]-#?Xbc
_AROW=Vd&^.a?.E]F3F\G@PPM0Qa=0K15JJIG@(e.M=S/EKNeYSR&P1:8c(.H91_
&5VIZR7f;IM=Nb<@^Jd;W-Y+EW\:9Se?[0XcPGfF)4b/d<(/#4f]##)Pf<c-g_K,
HA]d.S7@/;6S5.Wca,2.7S0dd[Q?<Ac7D8QBTVc(5[U6D>DWC_/10/(8ZJ3,J-T&
<E@/8YE]8d>);,=#+S2[FS#Y@U8,F5@_:+HAQG?@+;N0P.#H7Oa.cVCD?@RZUZ;>
YCQ1G6=Pbf?SE6?ISBK:B-JI\+C@].76g6FMHK<]>)GH@7NWC;(\L#9I)J>\/_G>
DN)<fPWXNHFE8JRW+8c9.WJ1[5:>D5Z3EV,1]F7d;4]5gTNJ)&QF/CQF6eb)4B.Y
LZ,Hc^K=((1_?g7_RJ.R^\Jc91RH+3O03EG?c.d8:(eJFeE_Z9cEG_&0aYTYXc+T
WY/Q4.,IPQeXN&&=HVN2[@K>e_PB@[-8?\TIM;J??>eMHW#9Y7CMDK#WYMADJG5&
B2FC5^@,TT[4/BO9Z,Jc&5(XTcH>S3aJ\IS;)^gKWS+2=C^XICLXO3OYGeaE&#@E
P>g,S8&>d3g,6:J7E:8a@^#=U1M1X;GG,7#G=0S4KA]J1PP_Dd+g7cS+VJ=g>\PD
ZNXAWO:/Wbc+,0OLQ&??J^YWYDZ+0WWNdMAQNd\-)NMUGHT>-0;:+]3;dVB+RU2f
?0M-S6O<F^.J+ZU&KD9QZEGgBV+I1-BBW(6KEVS(E,4@7R&S3D-9M(,V#M,Xd5V1
KJV4=0g@>e0Q\B[/VXKMgf[/:9fDLNA]#XD8PSOb607#+BO4>MaH=9#8+f[VK=<G
9c=8EUJBIZ_D643L[:S167]>X5d5U4d1LCJYNLbg@Qf5EMGe-R:7GV7YZS;#c70K
C9IJ(c2TPP4f^TU[R2dC\HEfSB8:OTD\KG5MgPb@9X0Z1GgB21RO@)D?)S4:MG0B
]KSeXcaM)VePQO_2S46;F+]F50\8R2e29XA<=c;DDIKeS1-U);S5c<_C<ENBI@C=
T8N,<\_BcQ5N2BVbS6QBZ45c=#P4V8b,7RH@?(B^.UTY\X2<Ma@I#BCK0;ZK/,Z#
M;<8BY/W=+^MMRJR:5>0Q?NVXSP=:e0O)HJZOc-VB(cQ=ZcSU9YeIRL;<2SQ)PAA
3(L)&?UD?8,PS4(9G]b)4<\1NbdHBc=aGDfY4?Y:=ZL2PJ/fbFCfe66Xccd7SH&3
3@Z=;Q(^CS\.BJ_fFWLF0Z6U0CHIL=d<MJ_?O(RD[HD.5PO]_Tg3PcI?X>3c5cP/
^&XA?=]T4+bGBMgb.07,2N^84e(\__C#76F4NGZ#2SNaCI&f/:@cA_PMW[b?3JF_
)R6)?)_c]fGWUDX0-0cg05^,L.,A17718<Q6f1[Z6<1]16TPJ?HDRP&UdJ-:.N8-
_7g29_\)G5fb+X:5X)0#S_a=97;,TbA-&AP7[D/d^@cJZR-7_;/73FX0Jg+_J<R^
CI\fT8&-FG.ZE(;dY&a;EIZ:6/TEZEX57b.O]SUO3@GF7a?\HYV32;5J,I9ZCL20
TVV5@<2fVUeFN./A<P\A57FM.VQVJT30H+KM6_cUC-8(?5?O;:CTN2VJI.d>VC8/
8>EK\ag(V#;QXNYGa?@A8]AVUU)&_?4Wg34X6+^@E>7U-[:^1P7.>J0Rd=0ECMP_
RLYaSdWgS8N6ED<5V[-[LBE5,@.ZOM5.<X77^e6)4=BL5X9\PbMHQGb+<9D7#:J9
6-\>BT>IB2<d=@3X_UP:c^JHg8GW=EU-H>87+HY(7HgaT6Z=)2Cee<RVW/+])4b(
N9<OKL9Q[3XPV;UYAeZ^?FXcPX_J7;0.c\-Y)bLZWBJ6eN.C]S3T^.Te1>4P[_L3
GCVV4FcYBKPd,BR9-,6b_/)4C<WRV-0I56N9Ze9F<#fC,+8\OC&[7V=)A<J5A&Q[
7:MT>DM\f#IdNI1Rg6=^.PPETFQ27DE49_f);d9XZDSDSY\[8F;d^)eH@IH:-9]9
c-]X7SOZ.?Lb:>K^A19&-LSTGS7Bd\f-I=f)M9gIARJ=^&#Z0@99X1[9TLb7S=V#
Xgd_@DKPJT[dWF-OGA>?)eIDNd^KJ0DSI&5Bg\g43\BE;6N-:6KZ=a#df/G_1C]:
861W)8?]YWE;d-7cN[,+<9J5GU52:gH?7ZR&I^UWZ(K/(aICI4YV468PD=O\2(gd
;J,)3eS[9f3[BbG5UbV,Q\X-W.^B-\O7E_+8bYf7X2&aadXPd-1#T)3ZaZb7O+(b
f];+Z0V5YBQSc^@We]@/^dEMgB4A,2,O^d?57QPA3a#S9c3VVg;FE#Y9)>;ZR6XG
PaFc_Yg^]XS:DF7gR2&.I49>#=VM@0IcH^fRDf/)GYM6=T,[.SgY8QS?QM=JTfL@
gD^0FSRdVeg8Lg78Ye3((dDZgU/H9>9JYaa)@KTZH\.M#JQF&DI(<edC<c2AD.#5
D8MTEZA&XT#GRSS@PZadg=;C<A[\@c+;)<OFc7OGS;/E?O)5_W04ZP1B+/?K)TXD
]=C2>(<9&N3,FEU:dZBL?[aAJ-B6#A0Le:WE/06IZ2UTZ<N/^P+P60T;4</b-C:9
?UUJTOJ<1/B&#78LF3X(g/Q[V(I+De>+ZS=dK2OcQ?OSBE]Q\6Y3=<#3eT/7\GWZ
Uc27BB5f2[T_,U;:AeG6].2T/0;g>?CB5VPc1R,@3SYA+AK/Uc<]>6=G)Z?-&gbQ
5M0=dZJM:bVVO.Gg+eO=2?D15+96?a0PETP-0\UK7NF#c91G#F8K?gLf\_]eQ-fA
OSLc]DJ:4A@8GB+N?)e,#.fP=QRCF#=>BH+P>K+FaY./A]SfFQ77aRNAE=^N;PP6
7T,HN_9#+T]A+^aO4M5(+.bAOG7JTA31=IF_@dc6[IKd85IE#^g57g;\UVHGd4C)
f&dNdR(\NZV71-I_SKf4#7(V8]@cb7;@Ed)0UP6PK1gWC4R5C>J/-gKG3e#N0+D>
FU63Rfc^8-(./]:L^FaEVX7ad13=#Y/^KV4fb^RICSIE:ZBMXA:UW1/2HSCB&Le2
[a9T0/V>=,J@XR_gE2Bbb-N&-,X:B/c:+BF>>SH:.44,GKDDda:1-/^V-9F.d=?K
#VbB(=a>(-Y.JU6J:.M\LC>4Y_MTZP?g=>L+3ABSLW9fLPfc:IcG;e)HP#7FC#R5
1&&QUYL2\M->_8Rg&;3G5]TYJcbS2/(6)L&f_7&WI@YKS@V#KDX@_#I#RM\gSUG3
4Cf)5K0:XgYBO_dWU>#SPQ8H?R^2P/B=>AI)GY3#TgR1BB9>]Vf.O/#-HFT6]7SA
IK78))/)^I(RD6:g.c4F\X&d,dP^S+SLU-G_R5C?E8b&^-;8B,RD4U5>M5W.e\ab
cV8&]NeG-_57Hb_T6(9<4Pg/f(b]32ZES,A:1::^<a8L-4Bg48\SGPOgU1^Y]e=P
IS/+S1B26R)APB1F(D7?D#;<050b4?fa@aJO2]KU.dM8?ZAHdggMHKdT62dc7-91
<>[L(OXa85:2dcP3F613@6c3KJ1XXGHDg\MG1=XYK@Pc2,Q]RKS[;d#HcM2O;cGV
Qf3_IT.@BD@O.fX-MP/b]8bYVXQMVVc/-[]CVDDSHLVa3[RV3N?S^C+)]Y7f^)d4
\_d(c=S2O9DJ-AaMV\AM-;J-B=7cEg1Jf:7b?J2EPe#[JcOWP>1[R+@c)=b1+T+&
43Y-7I@V.D(V/bU^3?>adWaAee(26[:5Id]03.AC.24JB2&V77(VYQbX#K4K]&Ca
(Ka2G@;;A<SXgPHB85&SX?2&LJIc(C=H37R<H:E#aCE55B:DbVDH1&S?X<eLVN/X
AKb/([)_[&E_XDf,B:g.^:>/4PS3V2:3IU4K]SB.XMgfL+:O:9[^X?950g,7R#[E
GS[b:#_>:F(S.0Y3[&R_P5(7#_\<\TAF(bcb@SJe^1_F?eXW+1JI(Q?2F;-eLYVF
4SK;Y_R4e:RD^d)5ZSCJ1C3J//9[Qd98Q\QA,S3#5C1H03TCV(?HFXgXVaWS<Z[-
?^dDI\AROLXf#b?WK#>DEBDVW0B9^0?I0Z8OSWGS;@1FC4XGN?X.PQM&1QLO-CG.
/8@Q6K#O:6.((#(N8bTWP=;_W5X7S<JJY-GWd27R&V02<&(.YT<_W:=YU)+Ng95g
7_bW),(MA;MFEB_DGRX8d[#WY^ASW.M?e=ZJS;R8/A8EAN-(1g)8=g\E#GTHNCUB
J)aW:Lb)dW3AI1IR-5-Decb\/RUETC4Cd^LP0:g>Hf2ZCZCb./)a]A0e>TM6Ze]0
N]V\YBWO2>7JC]M):a,?ZBg539#EBCSeYPYRg5&:O2eG^aeAU:?W?Y>-]HOV,4g.
_Nb?/TM4G]9Pg-7405R/83O+gKW36bQ)=7deK(=P&G0<Y?FBZU;-e4+PUM7)Uf>^
WgEB_<>5[X;],>3.fa2c;YKHB2Rb84V,W&O(:eG6QaQRT.B?H&VF0>]9D8F=IFZS
]b3;YK0CU4MKT)4@e8FUPI^Y8+cVRI+B-XGJ4-9YX3f0K=DCYT3#CcI9:..Sb&bU
eT0UGSB&fFfc/OP\JG2P::TcQ6,CMc^-JRZ.;=f?\?VX5J(8Z>,;]0:T]PM.DUg5
0c^4@E4.NdB73MdV-U]1&7D5+=f(&E13&4H@[QC)0Oc2A^#LYC+6YcTJG?LeIM0C
<DO=0@<)/X:Z&5]HR4HbJg^F2N-5AaJ9&,G&BaHE>QFg?YJTCPbaYG,f<SGNedTa
gY,&A7^I:\/Bb+#;A)gg(1IOZSdC)4CCW^<Tb_P7RDPFYP[cM]?BL/D2W3>T,S4&
=FILfI4)]D[a.>@&E4S+DE(eR(T.+9JQIe.fSJGO8+:WSI;cD(dO6.:-A)@Q/;b6
,?-R/-NU?A,7UB_KD<C5A?@L](dcb_P6E?YW)-0_MN#gCLG]^UcWdJB>_:1gcX=P
[.F1Y)cD08\+M_)AbAe>1Y96D>cRgHR).9DEg6:N;;UWKV=DOYRNL)a.,T+#W_2C
;4^2ZCRS#?,UEOW\c&c-bL9V<TY;@P84RK\;8REIWUY:LeM)Z@Ve#:HR3BZ4QJ_&
:QKR\5+K3V06/Y[SAJTJYW^IXSJJ[0J9F#EDAYO0O1cT\;&M&-W^9CK5O3EA>CR)
-2a.6G@\:_BdWVP/=U0WGW)c;Z79EE@CMV5D,1J8&bU?+fH7A=+D2//<Db0;OgfX
JcJCQQH&UIa]f2[RPZK?<JS&XSPUDCJS61I)<\+)+d^@Ib&]-.WM\c?Q&^8Xgaf8
[8I>@M&#bQ)&c6U==.JQ1GP>_2g>O(;H_#9?e(I&=8c8aU#JW5fELCSKY7#KZ^D9
Z,XP:d#LU.eAI-NMW8;,bNV&5g-:&)Rb1N:Zg_]AUGM8dI?A?GBY&IQ0B[KWLZb.
8eCMCQ/DWNdC<=)#_Z7YEF,KAbQ-#V.5e5?2RA+7V>)(b0I)/??d&7VE:DaQ+0-U
[a0HEF([\+(>L;(fVUgf_eeMVUK\A>LfUR_+22Q72NRJ033D_:a)J,6>)Q3&Z+9c
)QLXgd.;^-aDS5N4\-U8\)aVeI.U_90U\Y7=5T4NBO#VHX?;UdKbfXf^5FXL_S-,
d^GWUKL;?^eTP7KFcWZd_85FESB#SGO45\c68AS&Lc/WD4Cc#e43]f=J[?]EfEH^
bXfP/U>?)FC_eGM>f.Bb<I0+?;.TcV&(E/61dDaYRK032JTMT^,1_gMT<VgbMgKX
6OKVPTKN[\7fF4#TNfUX))[LJb8F+JU&5GCCeF0:8Kff0>fSEGTRSgMb:@f6N7W_
,0MY=4N#Z>>JRHOb1c,e36@-6T@4#Cee+ZLW:\[6X8VI7Q@c<FXA;;:@DaD:OKYM
,^#Bg,cWW7&)N-7<+OZG(>X:2<I;X6D-g37Mg23\8]V#?;OFW?1>XXM6[U7N=<MQ
9FOR^&Kd-eFHL>QH3AT0BEG6dK,C12e@TDc,K5>Da,F+@XS[&M-Ig;[9eD[J&L@U
)BVQ6Z(U6BIH7A@BN+0ERHH)M>1DSKBOc8MSNMROJ[^f#1V]RA29[J64,W9_XJR)
-dgL_=&B44\[gF[?.B7\E(ENT]J^GCYB(>YA=6]<3<W3:/Zc-:1TVW?+=6A&:D@F
gD02<&_DIR-P=WYd4(F>gNaT^L37\&bQcMNMEK:#e7OS<UZ1W:/G&4X=cb7^YAO0
6>I=:@XF5Xc=dKCVf/B7P?b42PK@FdXWR6.;,B5fXU,5D#GIJM&8a:FaI)N6:F;+
.C=ZO8>H1+ZMaJXX=I4b,.c73;:.e2c.Ca#.#V,M?)#D3fYZ/e()]WQCHMCF?FK(
0eSGBF.b5FKGB1._C[[OKa+Le11>1O6@5P4N0<I92,5QY#=TN_cT1I_;4bV:g0O+
@/V4S@GgHPOR0dEKN>>\E(,=Ve6#bB[7OZEC3NA-7^HNYH>aZ6g+<(>3TT6@:GQ[
:0;D_1^T@@#Pc6-Pf4MTTc+DJF?c/?;-S2R-W(3LQ68;#,)=75fI.0&[0bgQ2S,6
3C2:DHd7>cNc.F/P38e\)6+.<;XE[MFG?=LdbI86CRcSS^<EY7F<GS33=(9HfSEb
C-?I-RWgJgcd,Ag8W8/8^O)YFJ\?#,A)cQ:-:d,9b]4<Oa@ccEA>HWaA+6PYW)4J
+S@4aJ9;QB,#&D.c2#.DF/G4:^[K)N45L),LFdM.>#DaZ331&B.8_ZdN0d(a,Z@@
25JV4/_08,dK:Y0IGVCE^R.M;>)54)A_GD87+F9TWc_ONEbU#&0K^I+Nc@KIgL6:
,bfXOC_9N(a<[.YKS2b4?@0RK/B=NIU3PDWJS.2e=:N2TB<acN<;R_REK3MB1&Zf
EdS4ZZI4;F2)QT[f[197=?,c#SEF,b@ZL&]Kg2C3H)E:0OXT0]GSV#W:/@aAbf^?
3cRf1@@Z1(8#BPNQXS&cHAa3K5+=Y8QaYW]DNS\RfIg]U9?35MGGO,NG[W;B4-Q3
bNLG+#H6V5geT]3Va/0e@?5C?cH)[#ZQCJ.^&X1O+^c^G=_Af?WCCfE0M<Lc;ST[
1WIgJSBVAG1T)S/VMbc;>^D01[a+F#4A>?/R[88=6,ccT)g,L_f);U:5>3/0#Fa&
f>a::f-49-[()D7&?Fb:^KJ8&-;Z&\[FD62XR(??S6560N6e>c5F.&&NW<-1[V/b
O29^1=e@fL>3LZEf]Ve@E\IQ1Q;dGc54T#3KPEc(+_,ONbL.L?;d.UK+b](H^O)L
aKLW>UEPgQG06G34PgGPOW2#TQP&&bTB7P\?K67TN/3#)M7d6.2YHUASM1\;VD]G
Y[2M^][Xb<++HMH2=-fC5UB/QYQT75PH9<,-7f^BFaUF((<b(A2.9UOX^e6cQbFS
PVd1&/J=>.?XTag\VZdO+HX,Qg_NB873WcIQFP00]W-.BQ([&6a?<(KA9\N>;3<f
Z+:M\V#gNEO1>Ob?#&baC0[@_K=])EXK.b?5UN+3J9K7(;,R/^\QLe?]CA,=&ZIN
e8Le@MN_>@=f4LN;eg@A4+0W#11851Y_PDKM4NXHAa\-4&VcAXgc<\N>NHg><FIN
^-&>,bE=;40LCK(&<YX+#75?,3Y_Y((>6ZMF:\F_=IK;<?]?.3H?\fN(6Q2KcI?4
981Q1R>5cF<\D3ID/W@DEL1&<KM3?[fNI)C+I?>7TIBP:(NC,<eLK24:4fY8,eFE
]Y:=--e+;&XV7XPTB9Cc@+eW\WOfU-<Ye#U3EFY_NV6[#0//A?ZR>+Q[X9P.KSAQ
X.IaB#8e8HaHQM]X:\d?K1JHC/#((.1b0?LLT;ES9<E?K_@+c[KY6@/\^OW7BcPD
IeW3fAXFc]#]@dFL4R,SR.Oa0Eg^\_>M066GJX\_0+EGYBZ)f;d9?K\]-I=YGL0]
-.&AIP^GTKTUbBU0bE\c6]e8Lc=3G(.NEeR)#P=OD4H-)fKEPeY7>4]E(WGGM&3S
HgJJ0W:@a:b,GAHT2La8^dK+a#eER@FdLK#HC:,FcN#C0L5FdK-(/BN[\22#4EO_
<<(L/>1KDFF(M/=<Fg)?4_ZIWa3^L]baFN,_9V@1ZOP6\=d@\(9]MLaVRV)^CY20
<5a[?&F/?9<NNUJD>IWGZ9CT\I=R3<3Tbd(a^f;BNLMT.6W6RB.PHCP?&Hc\b5OZ
TF6G&FA7_4IN];>(9^&_V7QQ;RO_[98@H<6]5XNS=.E#1-K:W/cD#YJ8#/:3SIeL
&f1&ge8_BRQ&X?2-\7.56VNGaIL[>gZC>0#Y:d5OZ&MVZN3(M8_-Dd6RCRLfGU5d
7d.O)8RT,bQ,9<[A+BI_)HB6\PgOFD2<=DNJ9A_dSM0Z@,:#=cLS#EK=FZ;EV9HP
663:8[?cQB_1]HPLL6[:IRUfZN^,:T#&:CCP=aH?G+LG#DW7P.87Hc_UCR\cS.@<
)CB:NPF=QT,U<U..aJ\OK-#bQ&KI.ZA&85^<,K,D6[,I6VF4?f_U#]8EY3#^;+J7
HWI@I9EG:KBAHSNa_+g^a_]/O(M9L3#N&Vb+dKEA>AC_SZ(RJBKPVT58;7DHONW/
7MeMGbO]@FPYEN2Udf:6LHIf9])/cH9F27:OG)1/0#6AbW?J_#UV=1ODTC#.<@4A
&A)K/B.(]G:5Df:)@,>cO2+;7/OZC,c>a4BA\b&gGaOaUN[-44&;b/)VK1<DM7.#
VbcT/b^D)AWYR/V(a[683_P69U2M_&7TeWZ>g->E5S,X^6.#7KU3+CIHO3Pg\N.J
#_9Y(;.04g1ME,&BJg]R63@6H=VUS0T)-&;H@:c3Xec#34,F1;aG;F7g?S7^b2+T
\afC1U4.4;KGR?UYXHV0<&K.-RW;7X8&H4aW0>Yd#aTg&WI3aT15.a(D#ZNdP7Y4
5#B,4Gg:U.[+][aER\NPFf&MIbFN>/PO9OXSQ9GV?cPYR&1[58S5ZdWK/6O)LHK.
,K,_]?S8)W>OKC-D\7QH_6;FG]X+5O/XR@J1.#5b4bJ<&fHX_6G]SHRF&8ca=T_4
K&(((GeH@XT+eX4\_O>#,HC7S&b9_P?g;R87bcFH<WV_OH_F.TO@;@AD]1>L(eMa
4d?X_3]f8b/4>FUE,(YBFNRD@,e\7(_ag4[-Z=cA]?005X7U=)N9JX1W>fS;7LF8
K01.?:3RbR12J[MX&@ZPIW5KS\b_NC4:S#27&0@T6f-\]8@X@K1Z+Kdc2JS=:gWW
GT3/YW(dQ(ZT+K/^&Q=],65T]6]9GVXE?[V#dd#6NFX^P,((=JF6V1-Z@WP&8a)2
]HV=^RR7X[R/-LU+3R3-FHL&4@7c[ED_@956:&NK/Y?1]_#C^YL(-RGN=;Vf?&PJ
#Q&OF88Y2S#C/I<7ZdeR5S#VQ]G/PFQ@_88,22\0MF7J4Od?R=E54efM6YYNQZ04
6H#T#(F:,E6&)O_M7fD>LO#QDZab0>K^X<:,FA6YJgPd1.(GEb#;AX,;\(N1.\[3
(Y]_+VNb1=@,JQ2=[)2C?+YO5QY^X1&R]K_3/(9B8T>MCIUME+HVeX&3OXUM?4+Q
;=3J@TPR:cKHEb(c;.7804YPHXU)/#DN/J24/[Dfe?G3.,:@6UBD](<g5VMe?;9L
1?6(+d[QEJX:/UaGX4HO8f]?S(.T+T93J\-b:UO#,>D]+.@aO=U5U:X6IXH@]:G]
T/aF-gUN=TV0?-@:Fa@da,B1#TG&HTe9N?#BK1]&AXT]&@8WUZ97\:,BP^CYE&OM
L,&gS-fe6#EPAcf@G:IdEP?3241</7K77ON4B,Q4V(>,5A^V_O&-J9Na97BFJ9E>
]5CW_^c=56\H=FAQE,fT6<N=1f;EV^H)cc4HM3FSfAW(<1MVZOJa48>S?8=EIc(O
4+G3<AVQL=P6a.F^e,7RP51W#:7TM=UL:AACQ2#a]C+fV,b@1GI,fB4LYW>C6Y/P
]7H<[=)<:<[&(KCSSNKR7>GN2>?I5CYS9g3FYcJ2JN&V\4D4c/TY^_D:0-EJZL3a
\dMEU>KS.4-)5>@\N4daQYgb,X6Cb<;[PH:@)dg.,W(G70?PO8IBb)>@];;II-,R
T2DOTaU3K_VCW<]IT,2U+.5X)\MCQYdM)1E8D=8=8UW(<eMf85W7NQ)>@.5O/^04
BIYQC0^/VBW\9A@R0/?A)Re0e]8-KE891QS?e1RM+NRd7038=]A7-OgRbEV^fb2=
^[MbeccQ\X6II6]8:+#R_?<01Bgd3@8AZ,F9SE54G7)FYIU0COb+8&2ab#7X7TbK
RXLb;@VZA.P8)ALY78WWZ#W/AY6AIaLQVe,8,>RcER=&(CUMAOHcTH2RC@;FJTeN
&ALG?>I1X=KP\E;4]LQ4MZ:5P;4G7BTAS#23E<..NeEIW@1+DPQ8c)c60:[TA5XV
]R=&RITY(LCK]^)9PD=1S[JKMCN3-bZJH(4HMca]U9e\0LWF<2ET[=#0U13?Q_3A
eL1/XB)C5fA2^>gEIC)a2U)&1EPZG#JDCK#[c:AUK,TWYD/TK@^FH590:?@-.]BK
G(IS.T,.E3c4&GbNgE9fUSB.6+>4AH6U<_R:AH[\fWD\0De28FafXeF/A;(&FQA2
(dXR38/DUB_XQa.:G;[J-KJY8_-X-;P6LF</_OgDfASMU#f+f5N;&C.8D#&GUW3Y
fUJY<IOf-G_M3VE?@Y2LB(4[HXG3X4W2+&B)U@BXBU]<M=1_NZ.,S?a:VGK7;g6/
?2OS5W<GP6=0W\+KBSAA:E(bJRZ4WR,R>#/dKW/M,D-cL2.2Q(U52@HdQ54##GaX
PN8WUT<?Ncc[Y;\P:,<=R8BbFBVB+=DR^<+21c6U2K/a2,.a(2NK]a9-SVaPV[U9
XU<A\R^BS(CN(30CSA(U]-0;Y\HV9#efV#D6G>)?<(<Vg:eCdUGPfN2T]dOWScR4
ag]Z^-BA\^).FORbG3))5cSN-1g4DcB66AC,MXTcI;^61S:7F6JFMWZPc2b#W?[]
5YVD?16fYXE8Z?M&6=W\#T,4ZZGK.W&#MgCL\B)>G--.]M6Q@M;_3N3--K?HN\?b
I:G:20PTf=S6:(CO.9(&NcO&eQ-HL7M+J\(-BHc?;Wg7U.P_3V_^b.U_c[W6V1>A
AMMUaL<f)-D)gaE.+]_,b<A1BQQJ8eV\_OBf)2d=O8fUO7E@e>SJKPF4=6I0XN\<
4b>G,fF=ec>TYH(A0=e7985e11_6\T79+4,G9T_6a7@G=c&LBZ#N/<;9^V)=DHg8
bO^3?b=S#:9g#;WG:^Y8ZT2:)X[7E6UM\aBZ;&]#><ca0OLdI1:ZG2E/GdU-V<gg
E@8d\VDbYNZR+3CIc#EKBUeI&8((Z328]^<8,=F7RKX;aLRZ4e1fZB:BVY;3G0&Y
JRT>I=0N-R&-VA4\NSVV^?BZ=MXTH=LFIP,c[O>^\.CB>\L4TAB?cSPZJ,9/A(6d
D-N.&gPWPD)^(KBG5fYbfTX(X/2;Na_HR.JF.U=5I),^c(^D@R)9<>6OVc6+&4EY
_d_4.X#RYQ&O7AVdU=)@<cO4JYaDIV?M([ORNbC0R?8M#VV-CV]6>\-^?fD9-#76
-Z4K_3#X4:f:N\<:fH=b6R)T_LQ?1a\N/QBBLe[#TB<3>4,1B2.6+f_9I/aTF&E9
aK>R[b,d)L(CI@WbeMg3Tf:?[J-gL9,-A&JYI>^/TVC)RJS:W:L?CQ,5CKVB_D;9
::1gCYSM&5b\-=-H07IgN:=[;WJRN,=U(<#X_?/\8gFa(89Ge4^,gFd9TDQ^YdK,
2IA]2WCSDR@..KDa@=GUW;W\&C+f/5I:G:#IJ0G9[3NeP4.]1B<L#OF;9L3RT0>U
PU9KZ+HAM5g-E-,9#=:2&?0-cJ^[[NIJ6(2BW6R-UG7-Y\<?P1>#ScAeLNM&<E@S
WTAdc0Z4F(3>5Aa:=GJ=.BfP6MV(+-=9U_QLRG#1U,Fe]@.B]?9aRY0/5FQBS<a-
\Z1QB&Y[-]Eg:KaCFAaN-:/KJ2e#]:??5P<PDD<K?6L)@F]eHL.2[O3(E&+N_/8(
g&P=4M6-_/^TBg39OBD7/R,:>PU4Xf04(VX65Fbbf72W3/YDP.<:NKeV#5K1\eXB
VGEM/TaK+cR>.d?NX@8MEX(/DRCF=#PO68VEaR;V?a=NP<[H&LTI)X7g(;c;e04e
12aARa+VgV&KEC1R<](<+MaT.K-Ia8g2IL4YWT7D&YW=/KS>8BKKIc_7&,-HI#d&
CWAY?aTBA.D2DC0R.P]PS_,@gbO3O.c;;P#LeY@1aGH7+XaE.JfQ_Ab2ZSf]5g30
86F^OR---Tg]24<>ES0LU<:)N8N.RA[9=[;KBf)ZU0U)C:^MCdXBKCVBfTU(PUJ#
\ea=^#V#a5c0I?-IWS16X]0b/+\728,2F_<4Y./-=XY\E-Zg2DFH&MS+-N=9_Z]D
F8W^(XK&P7g]\;Rce81E4dH9Dd=0&39@16?^]3P0e=;6Q[eC\A5NHR][g0Z0eE61
E;g(GCE&OUG.b1S+5(:b7+Ya/5?bg7bA1KD\dY/_3d\Fe@?1.APZ@YSc8NJ.B-^K
a&?RQ75-<69gcaJZ@cR>1Og9d+?If596Q:._@>>6?.V1UNgeYgEC^;_+4cX]e>];
;JJ;#HUAL+GNSN(c7?E<&?a0f^P_3>)0#D=AR:_]=0UYKcLSZeT/G&4)Ue]UFCH5
DD)JDBN,<HCY(1#L8N0^9ULA]./JdWFXT1dOS9]4EbYDYMB\aZGb2LYC3HYaX;+R
?_6+]CT<Fg.7ab_#(+]R9[VWH#7WDM:GQAf08^3R3f@Pd)R3BW@:RJ,225\[T:#a
HbT,1KB6O.__FE?.W8D(+;_e;:dN+eaI2K#WGMCKF]LM;,,<;ca^55KHD04dZ;Y[
f(ge-.Y+P&T<L@D(6KgQ/ORM+M8b8aQ5)@/6I5N7#^2]e4e[4MI7aS.)Y1E&HQU_
PYeSMHPAX.fN<9f4.2Y5?.?^1_+;8?d^[#=CG889GObH_E97RM#dP](+WRF]^a,b
H0QQQb4\?gScVYA+9^eQN4BWce:VFI4@Gg5.</BE2DQ:HcR5F7X?/(;+Y(HWdAI/
0>Cd/>Z/Y[/W?7TIcI?\Nb^bQ3bBIJb=aP;c,)Lb9,/F^RIUPN99P;58I+>.@O8]
W1db-b:7(Ca4KfNHWQbbWC2=I;T-5;5E.G]?N)NSZ\e0^3B(KV6HCbcR]VN6BY2E
WgTgB4UfFC<Lg<eeC/^<&=3D[X1/=T48d?W(J8J_fPgb_6eLRa?c,NVL0K>G=8?1
;e8TJ)P-17LIW7KG5DYY/IB.<SO@Md1K=aH1:cXGcK0VI-cVH^R1ACY:8c?I]4YT
fg]I+6^ZP/UXa9]OOCEU#>9U;ge@[:egaG-K7.,784,S6(;M>V6/([]=,)aT2,1/
J?2JD5)R7R>Vf2GDC\_58,4W_YMd_)fE7;=.\/1E3X2TH]9aSc.2?b>R.N6UBN1.
/L@U.ROVMDBU78d_e+T<:R&KY:c]Q+5NEMF<)dL<M3QNcKQ>4W\WEC6b0Jc_,65?
._Gc2D1dX2@AAU@cLdC_Ec7eGg^,^3T_F94?1S-[DZ.4FRJPIDWg+/eaUB:)SZBW
TGaKUZ_D@a.Jg6?H(5<c.W/e#^,:aRFcMBYT>,)&I@TTKFFb]97:HM@1Ad5,:[7H
)W#bfG@J1@OM+5T7/=b&#E-UN90(9WP9\U+(<JI1@SQfg&G8GfSNDH<c](-O,Y7L
AeUNf,,>U1XI>7\[HWc0&Y98f]49A_ADQ@\Kf+d8).,a@D:R@c\.a76(8/+M\]2=
E2^^7-IaA4X5JS#3ORYD]Y:3BM/[VePSS66ZTf\&\NM\&CMA#I9?D-c9=TW.5_J^
.94;KdN<>6P7=M\+^QV]deVTMNRYVSAA3=/>JX^+;#;_d=J_O1(.97\NB7/W))UJ
CJ#K<=A08=A?L27X#;b1Aa_M:PdYGEMP+7?1VK;7,1Q]^]7OP6Q4A<04<DBM<-,R
)V&#K-14VVQf_AHVdL2I+3bV;eE.U@fHJNbU_C/d/WR3M.RER9Y#b[,Ge,/FDe=S
7)aYN@a0[Xf8g0.)UMfg[c9P@:;3UL-MNUUL3F:b24N3X\+0c=5;a+&)cQ/e9,C7
bCG^.#dgXS=?5YR^-C@90B:W0MdF+c7.K8;^<IRG[aCL#1.OW4&:D]]_7>9V&J12
?(AgaE+G-I#=>C0?WA:O(&+>g.<[=<,H(R;]G9O@5e^RVV<BC?ZFZKK]1a[/IdQC
HPKU2_GRC7#KB)S83NDSg#McPAX2(Yd:X06g,7fBU7=)5YY)d+c2QJJW)9L^;S?;
g16(W2UCH/1V/T<_15R_(>99C&Kc>3ca5+.EO-FIQ>cM2T6R7MOb(&W=Ra#-\Z=G
#GDND]\[Xeg@K[,[>,dd1K/:FQ?V-)8P98Z:+(D[_.NIaB).\HX-JOF..Ag9>D=Y
FORZJ_^f>&;M1MKFP(YXL&Q6RO9]ETB_5==WMK[3GB43a9YV=>)[a#BC)X_G)/<f
T]A_4e7AQ.R&,5:-2_0M@2JeI1KaE621IZ]C76bBcJ<K7W:/4dW?8H)dDa#c/Z\9
9:b<LCO)V:V(Ud#a#OUQZ+;Qf[@9-R&:BOEJ]V:_\3FL^@-R+F\WY_+1ZV:45PR6
Y^S6[;K9Se_?d)5693aTAcaHa=1)I^GGR\85,0LCKLb3H\O-#UePR2=H1g,6ZO34
K=4.,7fYV?57\L3CYRM<[Ge33dXN:P(T8^5=eRaQQC./XU;GL40+FbZ;#\-(cQAO
(KM&Q=EO)ZA<4Na,I:cL(KY[#4I<K<Z,dX/^QPFW@RA3HY8g[G5C/aeUFb3#WGa2
CR/dMCAZT/L45KeE]eWWbf(?G^M]WDD23,[W\^L^E@7+;dLKTRG,2]>5HR(-G\MV
8IWf56#JYNd[Na)-#BS-2LgDPgdb_fDR46/+&Jc\Q9??3#:-8M+?@d6C26_7I#O8
VNU6e&,OBLW\]gCd19bLQ2760#]3BXM5W.aMJ(0TYa[.T?DZ61a.N&PQ<PPUBS^]
QH0CBZcNNP?\&/RNA:fJ3C/UZT0A4g9V40A?fAYS-LATT\27>\I5f8:D1;[2Vb<Z
^&Z)_RC4g].gNZLXYL0QF+?7RXfBXL_(JKdQ/1b409Zd_K)@:W7Q>\#9L@#XUJL-
&Ba(X<7EO=ONCS)AN]SZK/g=_E2S5VP3O4HdfAA]SWF[8OIb59XY9NWC5gXO.E?d
P:SE2YQ6Y,:XaLSN291;\.>56YP+,Y30G;Y&bT&fcB4V&,XO1)->b87?L[:V6GGQ
_Fg@26;_g/BBZ<GQDP]->HM-).]B^cM@@PS6X_M:d?ABg\@UN>eOH+JJZeRY6SS[
2J>,H7E7M\&[3]U84TFBV8LB>L2Ha4(ZfgWHIcLca_PIAEYcf[&=Gf37VC-ATE9P
T4WJ)-,<AC1bF9S.O\Kf=Ca>@bG>WD++OA3bUOFP@+8eHE95KA6P#-&CKfGX6Q2&
0#LY8#R/:)YP346>&YL7c4D(VOKdL@Q5CYJc#P\_W65SQ(Z/6,-PXGT@aLMb9R_]
2V42dF7NBQdV#e-/HR+(g^e&PP;6c<Lb+&>?D_FTYbI@5J>S:1HGO9Gg1M6C6/4>
D^+Kc,DXX;T?eDYRK,3\/aI2:0^TPCV5OWWKD)RcfHc7^ZBgJe<GCMYeED:DSB-1
^#M&WEUQ+<=L8FLJCcQ-<Kf^3dZJ._U1;Cd=5HEe4,6#-CXCP>7O_3[C76HHS(@4
.9Z,6WGfJL^A=\+#3?E,e4Y?K,I-V6fc0DW/be-^UO-10f(L\c;I34EK1^75X_S,
,789@1&.0WD>@5]PTM#+P/J]A<D;P9.B?@K#]K4;>H_/SIS^6\>M-+3P3\T7RfOA
\aV3;W,DJ+g<]8fbSMcC8C]^:]Lc8TS<g]:OOI(Wb>+aHYAWbgGbBN1UG\8PCY,0
(O/E\D9/c(3RI1MIJE5D)X[U-Wa@cN+#97VXd\eX1J_be]Gg9)59<AX(B+OW2W1)
a3bE&O:-(]-e27V)1QCT7K+\F(4)H+FZ87KM&C,b8.gG^A8ZdOT5Lf?4>@94FZdb
:83FP:[2-HD#)/\A-L;T]@EaZ>XGR(VOZg-+c;16R^,Y+W.2-de_L1L&[<e5[U@]
^AbK+e)1SeacfF).[3>2/A6fGA]V,b7:a?)9fb)EZ?^O36:0?&5ZIM;09e5SEZ&K
>][-+0gM<X8.0JDKS2S>>.\_3YIg#1&b-_DPB>A^?a6>\-#cL&NXOGH6I>JJN(KX
0,e9dPffa8?fEZY##5B..P<^0FTW[9<QM]6Fb\Y1J88(.<\//,IZ:0)I^D,#[fL.
;_dN8FLfJY8-)76VGQ;[#[7_K.D[G?1^3/X&,#IbReObZ@X(M2AJG+C0e8B\IYV>
D)OT,Ae<Xe);/Le.#=BIAT6S^B:VR(A5[GWCJPCU5C?)U\=#=458>55NQN5BF<+)
.HXE5b;bUQ3bM>A-7](BA5N^e(1gaD;>U[0UP[QWUfU/N>_U7&>&SI2EeDFI7MDB
5A)<5A3N9+/UHBbPXW/.U#K2PDVS@&(OO83GgOZU\X&;;SPANT__JBIJd4AX#8JA
F:K59=Y;Hc<#(d5(2TMUBH8PU1fagO[W-e.WZ^E4S[#;APAZ@&Y+,6\+O(6L)d4(
^[]e)F.TSHOQOH&;G7:^=KDO1/?548G;D[6QX/A07U^gXXP4d3bW3C<)(3f8,=G9
O#M^-8[^^TIWY:H)FUXE@?dfP(Y]>B.XY(aE_93_,Q>9^((QAL4UNLWJX\fd=.g#
?&810UP(^bLCGVCOEAM7eL+L_-YPaU=ZP)IX=H8@BbE4Ug&:(8=HJUQ7(K2BMLd^
T3;#J]>KG8<G]5?+B7Hf-&G[Nb;C+\L;-J6<+]:^PBdg4Q,>]bUX\:<?M@@U=(^U
AfIR/9IL&\0Q@)+3D>T7F+55JF>5-AeJ3aPTUd.NE#bXOJI)GOT.#J6)Je?&+\:=
3CR)/aQ/+[B&Ua]>\bGe):7PTDa-&]b5d@=--M&eJ-047Y(Y:gQ,3d8+&cCYTUB\
^/8LS8VBXK+.Q=@??9D?_MDK1P++\Jd2)S@.Z&fZ^T<L,F^MKE()0?HXN.Qc0PC?
fRbfM\Oa5MM\>X:PLf)3c8)M>;&BM<K[76C(7+[3&;HfO7R#[(<=[<DL9D\4NgVJ
\I(T[_/B5_,3D5gPK93WVHNdMA^]^a04/A?U-W8Y(dHFB[5X]4;9_OMFFIQb?)8R
?)[3G\MTc;NYMJZU0FIc85>DaC&S]),e,Ud<O03H1Q--EVO2bb>6;:^10M,G59SA
8dJBM\DZN;8Nd>,c[<(IbPBa\=N3(.URY^]e+b-6P2]bJ^=M3Y5aEH(Ye&4EaUd]
dR164M/CP8b73PJH?;O.PbL[EK#)+[157aH+2@H49EM^K#fWAGUPI#JRf0UW]G:Q
ad[e__4d0K9b=;Z7.9W>2-OfgP^+WaSH[BK(6N#C2^F?[4Dg0]7a:H30a0G,.P<U
],?GT>J.([.]YIN1MNBMR/CD9[4^D3X/E,@(C_]HI>.bSc[+c4a3A;F5<Kb>Z)IG
_^)F<3gI0)+SI7DC9-S))V)D=KcaULYE9==L4HWZXG,W&H))LYCGNN?.66:AZf-.
:Nf]I:b4M9)/YW+TMWfH^-dR(9PL2/Y?ZG^3d0R;0(S=W?Z/83\]RLgGKN_WgG[)
/(WV>,2:VNO)[D-4R80>dADC^RJBL/O:A1M4XEK^CHWeGf4@-dc3gaN1-.DJd;?;
U\RFPSfEb@+RF3^KT&0.^\VF/4LGT,d?;3\CSZ38,UF3VYd)-WZLSTOR7<@+3>N;
MM?XO]V.C33/P4G7(AP4O_3^aeI=)CL:63]CUg(ZI<gUJgIb&-I/4W-3+E0d40-J
Z]G]c;eQR>WFEH@7)OVBS1PRG7@HTIA1;a=cT.gcKZc(bSf6V_I=8\?WSJT3F[1f
;^)KJ&B9#SO/F]<>_XYcg&-b1,5@62dg=M>/6N&IKJdDacBWCZB\-a4CV?1>E9V&
>XTcR2VUc;/XbPD10\d;+2XBf(K>,;TT+KGgSf0<E<_7>J0)N,1]]C2_U.OUUCg+
d^,)YN&GTaM5(3]6+OG/7^7f3c+J.d79^S3gLK#JFY3eH](XTG6L\<JNc9E3]ZM[
^,14:56P5B4dL;ZgXW;V,]_Z4IA1OEXa/4:I@H/,9F4C2C]1,eNB#5F8O_S>gXM<
YZU6bgM;=WSD\;O.XQXW0f>Qf\?HO?gWeFdPXD[.X0K.b@G4gKbZCF;fFGSU1>3A
dOQI1&WT70/^STXXX^,b^bFAKE9c82#69(e@C//gAQaC\f6eIDR960Z7\_=:A?3+
V?e)XDX>-d>6cP;89>b4^U+1W&YaaBMAH8X_eSBYA_[-+a9OeK=Mf,RcgA_(5G(^
2649Y]F,SNND>ZW)00^BPfJ&RLA]]+?8@RC9EWQXZ[cLBa@_X1-/MfOJg5>Y)g&B
8RV_WCdA3)YQ0XQ<8:B/7Ff,88T]]/;_eENU=I]V-ZFE(U#YL;@3MK<SDS[(G8#B
99O[/G\#Vg<XFWS2eKJ,M.<(25MU&9?@B@67&UY@93HQW#+LeCZbZN\E)27DKR<X
?0#U\L_A#>P,^IZa0W:^<N-82Saa>,2.(0CB]0gUL6RH(Y23,JN@/X&+@I=[@9UU
&C?^[<=A/M/G4OVMVa6Uc/-#CVP,N\F5@W4Je;??X(@Cd,R,f]M(9;5IQ]:5L-OX
U,b^IDfZR\,)]Ng21KKa<8a:K.3=KQ3Z3a__faD<8&A<<U[HacQK=D(A8HU4D^I9
beTQgDZ3+@1,98OPa;OR+fR-6Gb6KVO)GL^U3,,H@+DT?1=b>4C7/g1O(C=^(-4[
2.G5:4H0AcGVXMU_RGL/AZ+gU?U;,V;O1W7N(ODNa^<;=OJd+L;SKR\fcT#2S59Q
CDM<GP]=[,]57c3)46-CQ;[(8>CDVTM_D[\6=Q@R1)f<74[R@SeE67Bd,+[V5ZI+
/(X9R)&Hef@W_\fU>AZ-C5])SXH8^b-6:NEL)1D_.3gT&)B_(gf&W>)&)R^J/gUd
K(Mg67QXP+==44;.U3;]C31Y@.:E[BHD6HLAdPbbP8=Tf0712D_0&g8fFP@F2[QM
X>a[aUa8;+7[Va?;H^YR>Uf^/&\WDGSda8I5>H->D\_5DZC\/&KY&;+VQXR0YYM9
]4=e2L3VbNOQNf#&ZH9JMcWKD@d=M\@@5eLOYP:3XXfK#IIZ]b8acTP5FIM_MV3c
e<d(X\GAaeM,X\-]:,CYRT]e-1G9L+X?SVCBT/DWQ9+@D^^=>#Y]Z>C+7^/(a4A#
d51#cGX-#R6=?\0J4>bVJ:[<NRTPNZDKF@^f[\b<SM;VW#gP&dR#)fE.3,/\D70?
6FHHTKWA^Z\P9AAN9bW-__A&T_,=>Lc,M[US^g75]/3?0;./CWb-SY,1WOS(<;d?
M<ZLB^Hb(YWIbd^3]3V.HK.E/K.MEH+7V?<28=5#./HaGIfJ+>=gG7fCJc5YBTbG
7Mf#d7b)\_^]#g0#Xc0E7XKfJ:dW#52:DC7D??+.RgH]g3D#(R3IXG:Q)[KD;/;4
TDG,YA]+Xe0)RDT?cWF6/.gXeA[,T(]_:RO0KECDaB^:L0Q;W/.)9X+FSJ<//)bS
<NV:T\F?]LRab3,5-12Kd4L]#&X@1P<[ZCD_O;:,:OCX1_&V89Q]^QZCbU;.2EVB
Z[-=f@B[330_&\I^^+,7\<)Z)JL5=KGA#DGAg1;T;U\VA2ZTB9bA9?#DE+M_3eM0
-G:XM-J6AEFZZ6QFI55Ab2eTa:DA[OSG=Y\M^0]7X;=_&57U2KPMJ@O??O8@8+&V
.8PH2B_@I[,+K&/OA0_-[2/baY\AFcNZDVO>>WXM</eR,/c7\CN_RK9-J7-VUYTH
E.Y9@E(Q;57=Z;55(4]gMH/D+>-9;bVeQ(T@:)>C;0N?Cgf.NQC@J(6>6+=X+LeQ
-QVa1H9.>I6\9V>^CO\C\QCBe4=^MfJ(eX6[IDTeA/>bI/994eN>0P]aI,]D^G:=
/1M>bX,4=F>GBa#_cA(<A(3O8Rd&6L[:J@5_Z=g:_eW;J_JV8d+]C5dBDc:AWF+/
EQ-=7+;c6L9c9)2GWZBM)++4//W9LA6/V180(17]8B;e^&bX>ePU1DN[0>9H7ZaK
c7(IbQVIIDN&E0;89WTgQ+W:8;c,669UV/?,2fXA]_V:VDQ/?.NP>bgS1bE)8^D7
3K7>1[:6QN,4OD:+U(:WS#ef&eSW<P;B6EddB12aE,R)Rc>25#?N83ED,:,OZGD)
PCAbHaD65YZg\A(&f:\Tf)AO/f4#_Q#;P=G:KLE+dD4UU_[(CU2^L8eDKRC6P9]-
.>7ZRA?>1KO1e+BB9ZJ8(D-Zb&f:2[@^H2EI5]+YI=&5c^26bb>S:#aILPYFPVWX
#,,Z+HU]7H5cK_97/a@M]EE3VP4g4Zd_5(ZR8/L3G8T[R+)]YZU@/)FU^2+(DBdW
FJO)2T((c6_BKJWW,e<>X.gR?gQ@WF1D5I86+J0Xe67,BV?2CZYY#NadB2&?ET)3
07]80Mg3Uf1Y-NU@0=5(&-/U9TXfX(:[c8g->Ce(><=M[aZ#eQX#=^];#0./2fB+
28\Tg;2@R))@fHa@0f5&E)Bb4cUQbXC6P;MfM>3V;0K\_Y6K,A@@(#A^:QX@.33@
<F+8ZYKJWbeaV=UVYQOGJHETIG[PdE7/B=R&-C8,ZGN.)@7\#1ZR6H47)J.=RW]J
:LACQ0B+8BRRS?F[5\KSGW3#OI>&+e&/2[B7(+J1^[Y12S=&JY;C+CG.1fH4_)5=
FT9X/.;ZdR,N[+aO_ZZ;,KCKN(;1;F3JMRdVM3:M/H.K=B@HLc][MX3g#aEUWMfO
F&Y0fa/D-]O/N^?Qd+N/^97HcIT>WJ@c&+,CcF-49GSTG<.>bd2+XK+:V\D5+>^a
P>#e\FBHVH2#f;,1gPU-a,ZFDcQBWf+&>1TFJD^O4-2],^2MX@45O@:/@01\8_BB
HTI3>S5dZ@08KG/3L,_=GBaSLR0>RdV42fRY>Q;A=L;_RI-^W@ZR^9I6FG?]4C5d
OM?K:NJ4=ER6-eI)>V3OB.#(gEa1C0=gN-fL\76V]Aeb[SMN1cE<S&P4gA-)J6H[
[bRHU@@dLU<XSdY^T0#fYA8]gA.3#Q2QBd^Z(B7;)5Y)P:b^=B;+N7AD/E)1Z[K]
7I/KLD1A#HN^?A_(:DdP4;2ORE.0]CUSLO/S,VG;R7cTf&R@KbB^<C;]H4U1-RN_
#?a>?_eF_9d^]<9GE6:&.Cg58P/a&W=2TZfLL)(7FLScI5YH?.ZbaL::::;_G5Y#
MU\NKOf5T]g;:PZEP8P3(@)[DR=\N-S\d8E],CL3FE.F(9JR,OF@0WcT@aT^OF37
HVedV/SW29?@2.JWK]C_B#RQ]X]g5Ncab?/eIICCA#T0<.L]1A^bW),)HgD@:H;K
g5AXVSKBR;=;[PMBMN^Y&f/TJ+(M<ggK2d@@eYU\E]7Y1f<OXSJ=bfJEE0PC&0P4
30@(0#)NbX]//9?[)IC]XeXP_cg;-E[XMF#EZ_0KF7)S,P-6-;.8/(5F9I_KV]D6
PgBe+@fZGEO#)3YS:/Q]TB:U47XeJ:(ZCH?8N&6Fa/88T<#cNU1>A+<N,1Ka,_:C
V,Q/TJc[>\-C0cJSM-[72CFJJ&1(<W3#-aPgSB41MG?71#?ZWTDS^T(P\6BHgPb=
1#;<#,39X4[=T1452-6Y2aGG1(dG_Vd2/O\(:-?:?XF2-B,3,\6,IdG_58V^#R,L
#D&>ff,SY06Q>IC0cII>W01W,C7:ZL<6&5+V.FNWG]\YJW:AVGLI5Nc_&/SQJ+eY
#^U8ANg</Ib5^e;E\]9&0I.VXZg3bH/:97\<f0^K4ZGMYI10F=,.EV_gd=AQN0(/
NKQ.]^YKWEa:gLG8:Mf1Hg#-(67+de8CF[2d8d(:UY[.F:JU2,L,IV_VO-6JZc,W
<GdNF/9](P#750RfKXd@&R,5cJSV]Q@dU&=W0>=5bI,_ZS#]@.WfbB1M#C\RY=;V
FdcL4Cd=S;aV2:OO&>IB6(02AO]De;_]YQLX4Ne)&;g53#F=VQ2>HN[>6FTRN;DY
972_;ZU__dG1.eNX&&YdM.4deU@?LC-5[]4&?eZARTeMd(J>:07B:5+NK2HRCBK(
\,D1:V14XNH0Ig6W09L[H-3YHBFRPCWO)=\+W+?UBV31#K9?BBN;#Ag1;<<0Y+N/
W<#TO;)Q1H1<<<f;aeGf#A]JF;\(&+//SV_DDIT7JYd&L@97DOe-T].:^4CTQM^V
8S./:cC-5X]&@R@K_+SR9\DL^P(-:01Y2&L]>1SL\?6C^#5_c7c6bgUM1dGFS0IQ
QgaG5GgL1e/652cRSJTP[XPe>4E^XQ0JKPE:W,/OG+,94XZ:^KFA:.NJMQIcW^S;
Y2;RUCR.=&)<92G7T_]8Q/FV5ODO+FO4D.<-@B>ZZ82RK7C.XceCYW>M82e?AQJT
:S@#6[N5#KaF)b>NKV<=(5-[\-KA?56_K([fUQf1,4\:NFD=D\9QKS)1^E5D??Bb
A=7Y1bTX?&=#UFCLGe-+W]6AK@M90C^a>E/AP(8#-^7(cg2+P6Z8d;M;.TUJAT3N
CeYEDc9OG#@QUQFE4D@G^6eeO.f7BPEfKYZDd\[0L^/WB(N25R0>D)=3a&1EL]fb
<eJ#>;X2gf@TSN54S0EBg.@T]H8?A6ZA0FfX_F4a&ZLfc2TbVNOC/W1[2W6bZZ^/
<)D4N5G)dJ>e\MDI+,?@UOS?9P3#HW7FTe[#[B\b>/WNE1=;g:U&>QWgf@6P;&24
R,L;bVeKD;d2@(ZGO:Y8e2MRUJE63f5OSaI_[SE2RV=MG3+<<Lg@J/_VH+b]#:0S
OO.Ia;/=c&JAL\>cgI&R2HYY(][I-=+bPJ@3Y&J;E)g@ICG#35.,(3C6>18(#O:d
EXM=WQ>-H&2ae_AFO7@J#V>1DJ.-DSc(=[fZFa3D@-#4-8LA]>:28\/^(6Ig[S9U
3]@DVL=cQP.8OaPRFR39[47f)LJ6[+Kfe9KPg5E\)Q8]SH&@&;T>V;T@O)U#HPd0
00,>:?E<<M4E,bf,TI&JMf88M)2:VC&L=:W9@AWM6d741I;[12Y4gF3(0A]YO93a
abGQ2T]:WCdB(ASQ@^,^3b&S,3@<YO(1IfJa3Y#9-/7QTC?_#?gYE[9.bBV.:NP?
SAI^eHF/#_M-UQZEUEf7ES<c)@215&/@+.1<YE-^/>V6C;F+?U1e@fXT7F2DP>#K
3_.S<dY3N0>V&F;K04I.KMIW))Y^V.<_(HQP<R.\[G0_?61:#(BV>P/9-^Z\Jc4Q
FII9PH]/XV^#MHIWIB@afBU^1)Q);CMNIS5LXU</H0.ME)g1#=--<5f5GL?PDDT7
C3T:8Q2Pa2]Q[:7IdI16E//503OIYM58>#F2N2NZ/0V5Z:W8_<?a3FW++1f0+8/^
cKWT#H/?<>Y?\<0.K)GOc),73+RH<H,.Y#M1SIbe=M)ML80HXggHJ]627TJSSZHe
=O/#eJN=&eSHLJD0L33<-W2)\3aM3cd:egU-R)JHQAP?4K:7G]?FbWK1C<?]A7fE
\>bN?<0J\UO<9IJ]1eW83bd?5A8VaQ5fSLg9#3)?ZZPae6MdPC0CU7P=cTO(\EDT
=9fb^eCg/A93egY?UKQ27K\+4^V6c86WVI_)QeZ7_bSePQV0AI<a/b&VKFO:XaJX
MY0WM(GbY^5TFdPN8SRX>g\76Mc8^aY(#(a];b05XO4YH#3:N+9Y)FC?Vf3YEB<R
8SgM=:OLQPdH,\1F.6I>L-Za3.P]-_R6f&+H:2:Oa>=\LU,LR#\4C:3GWY195e\7
:J;>Nc<?TA)#,MJ+R+EHIDI,)[5NPc=8I>IR:-+VDA[.M0_@CY0[5D#ZJYN.\E9<
)E5\a9d</1g]2X\e7[g3CYAKNPNUCDS39\X@;<d(J4UEcO8LS4GDXaKX4a=)3bD&
D4B_U^OA0V(Y@FF,SU-)OM^JDUMeIMN-5DJNTI#\X66Jce0+bI]9;V4T^Sc_,\f2
@SYd_XdN<T>(g3;Df/WeS\V>@,L2?3\)((bJc;H9BBWQ5(M2A=NPX43N@_S2,5bB
4_WI@&eYX\WGQaXf7#>;O#8Z5B\b3<A6a.Z4JO^)gN8,:Q<FDE6#HY)e:7-\MZ9?
-O3]@T]BgDINT1:Md;RbB9.gHGTB&()Bd1M=?/XUQ-_ZZTJ/gFQ&6@&A;eH<1>-3
B)?\b[^fM<bDT/7^-TdUbDLMZO>;&]CTDO6W.=Q^6TU2TWD.E&ZFPZUa6.JG>UbR
V]]FAc3UC>[&Q+BLgJ/2NB8XV2.]FXWad)8A:CIY3ZFHfIX@Tfb7d:>3D,>Ma&.K
\5OLaKQ)a/\3d@LEA-XZMN>NMOV2F5gL8H.G]8@WGZO5MALaC_<g\,fe;.Z[P2AO
OJL:<Ba\2T#S<0],C0]>8g#=8CRUe7G9U&X#ZD(=5+gcg/KBWeJ2@b]GO72I&FF-
<;<fd7S#]F,D>M1Z+-d-7KbPWdI?5KO^DUEHQ;]ebJ/#GQ/J_:73:J+DdbP)(K&D
V9:gJ>]^[SXS./\b<V7282/_CWJ7F[(g/&/Y:C:3:34AH4g4a?d=72-D^A.T&MeK
)>EAS\I4+3(//&R[L)49>C.Ae,03\-,VN8/,T5N0&PEP^8aG92L70g#g>#J<_8+2
Ba0_[4W(RFJSe;^X(-_=M>I/E\Eb\(1HWf.:9474KZ>,[UQAV.AXFCYEU=?F?)D9
K#TgTGJ=CCL)6(][@/:a9PbNAf=H=[DV64B#,e7^Cf::E2O>D6fW<&f:=8T,dTUG
9g5&-Y]X:G43[)g@\F?2K2SMNM+gUc+U5_.eB)V&FbQcQ(+8L[>U].=A1Ad.\eP/
T(7C7+Sf7?-W2&<5:<2O0eW:(VFLQZCB@5,F?IIO#[E/E:IE(XWFYaX</68e0+7U
E2Qg+KWZM416Q^4D1.SV3&(a=5/1fg-b+d.a-]JX(J9EZ(0Q8[Y/YP-]F,J>T&-Q
X+6Jf#:#:eQ-F3SZ,IMXPH3_(BXM<c0T[K=GgD0-cM#EJ7I8U4.@;6b3\)F([dB^
RRMKT>5<]R<>[eY3(>UN,,W1g)fcP1IQ;/..BC-G/M4R)?>JL3\@U/b^0?T&BJ9\
-d//HU@&>-L?WJ>5f6G1Qa+d=H&++UEV\I=1RN&:B0H^@aL[7H&1@Qb-B)PE2gHG
-186&S9DDXAXQFA9gI^X,3BRdXG:O7B#W<S+;/4W^X)&-f+a7@dN,YYZJY27#Ud/
5#dJ>J56^464[BcXY2&KI&P5]f/_1ZVMB41SL3cK\^&YPff?.fVEJ]DW0bRS3U9(
GQ1b;cA_B9\\FU4&;.A1G14YK0[HN]&LR)^bVA9:&.g7TSJZaJ=^XZ_@9d^TQ(U]
a(bZO\\Y;<SB#>)@&B4CP&H[B]?>C6bS\Y\5:&f@;).ZO)B80/V[U_WE0aC\XM#G
-g)6.R/ed:1TM;K?[VT^5dW]T,Od]&S/JI=dSePK^F/DaFYccDL#.VNV0EIb5NJW
6=@G[a]f.J>#;1Y6Pg^>I->N.9_SRV+Oe;;RCfcY<G+?IK#2=Y)YgeYYHe/67]Dd
Mg.b3e>0PTL.CE)5WALJTb/aQBeH+QJOUc-=WBIdZ/)OTKHY#B0\87+\0c_B<;@<
UU7T?MG]6OG],H/<fa?Ec_?Q69See&E,L,9#0T#2P_I93Yc-&g.g;R2;U:e8D8bd
ZA@7N9#K&Ac)/Gb2=^S0?gfA\&a(O.\>aK6#R3[Ue65aF8.;,7W&6E-N72-Va.Vg
QUIUWS/\</BTIQ95bV8e:N#Y7.G9>HCF6F^0G#XF<R.Wd-V9N(X?7PO.L(J=-^\@
,JPMEB3838)LJ:3_U#,?K7CPca1YRQ&SEY<X\QUQ/TC(UDQ&B67^MBF#P(&O^V.6
6FDVKT1b][A=bF2<.0(2P3g/^P=Md)W_N[.>5b@T71X4\WS_T2?7Z5D1RW,TG&--
#OQaIO19ReKE11;:U<(/B/96#e:(,9?MfVV@P>B#JZBZ-IOYO507F7A\P8MB6#&T
g5)(4a#8a58[+\\ITMZXDP5?V4:Pa6P#H]Ydb9P.C=/A+40[Z@46-73/]Y]_:K8;
^B1W<TU<Y7^SVT=&FFK4WIGK9SM:PVCNW2>&WR?,8e^W]G\6#?\1LUTRXS4@XD\B
>fD\deC<L1-[RC.c)&<=PTDK96XeP<^W#>:Abec=agcMW-A:Agfb,D9D0C(.<[[@
^_)C/7,8d4[[G=TZ(#7d\Mc<S==EaNKK)A87gQTI(0JP(7>\>;c=;)c:>:4;cYgM
D-a]R/cZF?DL+W?#9e249PT#2:d,H]9+GH&Zg_=E),0@R=a?UeZcYESLeeK0O<Ve
+?3^>=gV9C&XVaPd).]>8DH#RQ#abJW&+FD?_@aXN3AfL7e^-O.UgWZ4ITQ:bFKU
5FL=6RR;9\<gXJ?dbGYTZZ-O/Pa-=cc_1C28B)Ec+JY?[W?,V;IaD;V?8_?N3AFQ
[AH84:--XTELJ2):Y,H][bW4]QJ&[QZbN-YQ=;a]GE8XH>ACS5YGX:[HL7/<HMQI
)8:XNB5854_NHNd/BK?aG#BI>-Z:0L>3C\-/KD+N>T(0eUO/gEK<+-OOYd#=<g96
Ze-R,).ZOT@5Rd^.#N4F3G>#eY@/E;W-L=:[<Be2<+K0(eDPA^]0P4&K?:Y>Z;W2
XX146&7A\d[Q/EUBLHFMI[F,?K682GP9I@A4/)9aGY6LN(Z-INS5J(;g&7Ua[-(2
\7&(c?ZFddaP/J@/9.JGMQ^.#0NBC;VB2#M(3->3K8FLM\@4[W,JG[MAM)-QQXQ@
D\_dXW56aKI4)E(A(Kg]IBYXL;3B^fT(/U^9G@G.;__)8Q#;QD38#4E4N2X\4O[K
W?F[N88IWI;T=L4]#XfBaC9fI4f-&:B;VNg2eA3;XH=,3g_dE1TD]Gcd+aQ7#W5M
,?#Gdb3^eQN()XW;>(JL^&1\@R1U4+?.\&(.Y[]:b-QUJb7]egK..Q5H6&<6:M@\
[59VMcA^Md\Q11\9(E+GU9YOV<6N_;f/4[\U=FW6<&L_Q7;:c?Z84)C88?&I=O]B
DJZ=Hd,f?Y)T+DR616P&a6?-RU/G:<VDb6>@G7ZLZ,e+YNI7I<^L->bd4f-1aQYa
^1C&7,^V=5A(OaQH&#-OOWO9LYW_AdTVXf:&O/B6Z3+52X53CRWbT.8/B>=,H7TI
Za]GKC0/c(6P-+M<TB121&<b/O^,)/PZWB[6HT\SCEVFO)TE171Sg[OJAM[F:Q_2
LHfZ>6:RIFCXf<H>TPTAagJR>N?b,CL-L5dCcNK.fPVYL5_9]<\fQ/DG,OT>F&YY
,P]1cK\2eRUd9-3Ab/W>D6aOSCb-S0?J[e]Bb5(^UC:WQ.a_C^.gK]&4#O.R?593
R#-Nbc6c#D(^FdP^6HNB(Dd:&-f&L>N<Q?)M&Rc\#NL^6U+R>9S>@4:I;2V^CH@0
[AafK1D)4RD+O873Q.7a#=LM?ea[EKA3O+BQ36I35)N3]04WYMA1_/E/]HVeg7e;
-_S)4e51@Q4MH278g3\.c:M+/+RM6NMH-E?^Gd>:SRPHJ5X\B^^26SQ3XZ&XGAI]
HYe@H,_0ag8]Y=NU#HCdMM^+WX?/W5R=[H#-R5bLAQAf&e19;P2ARYLQT#E((U3#
B6CT.dA5@G[OA);cU:/(5YR9(MSbT7XXN,#DWf^D3>W+>E_62F.OEa;;;9B_c\KL
J_@60=HEb21LN;?KgWXPF&4EX5<SX/K4D4D-.f1^;5L>Dfb47;D#X4bUMDKD];9I
R:MRK-_J\.7Y+LCb+OP9JL\SK;83,:/5H-(8)7),IB/7X@/+A2;7NNYg/4XeDC22
]d7YQ?5K(&^+L.P\XU-+Qb@F+R04O,cC@\Wa]2^G-;.WRP=>R]K:[+04/QR8,85U
)cSW<-7O)<f[7\E&,aYGf@4UP3a\>>,cYa:ZN:-&^=X=Tc>M>J6PREUW81K2-K[Q
682e<TWWSC6L][7^<Q7g6-bR>N2f\]4aI.V-cAIRZ,UKS_]K2U:IU\e^7:c#c^J=
;_:-B\=gKJHA_Y;b:35DL-.Y]=4Y/&gE0[VX=(E&P^8Wa4dB/0^T+JOcWG4<R3+a
2@#Q\XYP?]H,M.+5->E=8)4cVP];<XU;?1+B8;P=DBYUcE[UP/TA?-8e:R11B_BD
6KRE&1#9+CR>7?[]CdC6:a:N5)O,A@8ZQ_=-(f.BI76Y]RX/Z8]Df0^@;W\RI:6X
](,XFJAaCWK;KPKc(-&2^81?]6L88a+9a83-_4;ZZX/:P7E,C\E1cC4&UFLb;8<b
>5Z@^2L6DX;5DJ]E-3UeKVDg;,G?:><]GI/FLG3dJ>9XeRG:2cB\V:P>U)9+:[Gc
9N&5?cLdfb3R)O?SVDHUDXNR&ZeZC5AROE\0^B#,RX1OBGSS\c3--9WXTJ6D]>Ab
FJ84#420-EL.O.7PG@HcLf;7T;-P9#\=3G)I([H(+@fXP/0Q7#Z=>K=HD45;EFaZ
S;dJO]:30cSa+gB\)3-:.@3?)Z(NB+-PAVDYAX<F5eYf;N?):Mc,(UBO+e5K8U7J
/HDeIQL99dH^>)Fe?>B_B.&NZOBCE^B^PRB9HcC]VQ>Q)+CL_J\\C[3O]Q9U7IFW
3&[/T[&[3UNNF)QD?]#N^-?;XH=OS+DR=Z4g_0V1HVAWJJA]T[(U(-S+QNZ^LFZX
:Ve&V/:)K?f[LUd4]bT2IeI?3K@0ZHQH+3#.)U.=VFAUD/(>?SBT]4_c?<U][-^O
X<@>>1HHd@6aRHa_:Q=QV,Y+;Df5<D7<+g&e\+K]:WISS6#_]g5DI=7IT&0D5AaL
UUR_L?BBMKQ_g)9YIQR8XcBA\aO,V^IA?gZ=g65E74]dS<V9GbB)=dC0)2\NAP\4
A6HU<f.[)9JaS<,cX255>N;#K.6e3Gf5DPXC/6N,4)U/,_CF-4YZ=ZB90(G4>PR?
+/3K=5deT-A#I<ZS\R_KbS?80=8dY>0N]5]fCLbRLK[NeOBCHJ5f,)R7)dPOF<^T
BKX^@K/Q-6ee7I;<,a0N?/<G7H_T_RH6gGQ@VDVW/&dF^(fPMd?),2gVIZ.Z+f2b
6,F6&a<-AN)Rb/&G@5?]D=bRNb0?P2.3KDOIfCDO-:G3-X85B^YO]4I,d)3Gc9K4
6Ic)7KC=ZN.0+2N-:[B^G,I^VZF-&f6.K-=.>Qe2eBY265K^V[,8CZVd5O-=Rc&:
2U2#dZ:)R^WfVJ:]f<&>;Q]CV\e^+OY23QSc]1@=]Gc=4/YQ.UQ2?aeX3\@U&R80
,0;C:_,(]P(WaNBb=cMS9LW_a9X(d:T7\Q5@@OgUH#+C#d7]J]KY?84A+U(+PNfK
e6MQ_?C=Q,f7[#D]Fc-MbX)KRQ1X/>Q&D:]8UHd(NS9[aFX=BB#4XQDLG=YA?b5M
3aX(-2.LJ#dR27V9fcOJFKSFQ)DJH[M7g=S>8<];bNMdF7I-[a6F2Ka7T-FIe3I/
^&I7:P)gL,)>37aKDJ<W&9(I:/@RdfBO^\W95RKcaVV8(]>(dKAED?b,=PYB9E3a
F\R4EG)<e/ecJYbK]S?T7_6P-H#ACSAKZ6)2eb]H=J^NeC5U#0E[S2Kb#W/e0c6M
\)Y_V&?=/12)X8d=cCY8LS&<2V9DLYd/aG?\V(A>F3T0.4F?3?TMGBcNg&;UB(W_
\/W1N?>OTQ@/=0WN<,+[.01M>=B.IF(SU-gU:#:b(6RbL,]-AMRDHZWE[<P4UMP,
fdNOA[)[)3920/aGC5V;>-S7bfG(ML9M@]PEaI#]c?BNZOX08--2EYS?fC&?-:e(
ZaZU^&6f&K[_ddQfQAII\[X./aH>/XOf=4QJ@#OK1XD0d21(.M_X-g8H^SQ12@S.
6A/+:;9KRZga[BdZfR;)VN7bN37L(D[IBK_G2[^IEfKSUNW#-M:;dMRAbA26Y0Z+
AK_SV=2A,_>,QG5HH.GbBMB-Q12N83;GO)4+=F_/&E+=EIX?T95?W\8gPH\dK+/d
:/<EbM&KKeM2,5USeb.045=[)II</NgbE=D&_QgSO_Z\N:WC0If^L5S;^_N?FY/(
O0R(+c]+(-QagBX.31[^I(B1@99[QRfF10]e5M\2S.G6C4_UVX35b5XQe/cdL>aH
S:R#-((/N1247T&FJ(c<V4O&ZAM?Z0c_Nf0C_LeIf(JO2H@LQW12(EVU0:JT8P\2
QS[[,fccfbYV>VBgQUVE--I;ADXV5@2QSfWW70V)]_\U\Ke+4R.X0AQc&978DKA]
dH6JEKgG1\F_GbKIGIG:3]f+eEH338UFaGScSHG4E=KLS#c6Z+>aI84F+3@;B2bI
@]T9:4(,TAJA;];#Y2YNT0(;V]96^<O9V#b&GG@E\LQbHR;R65D-KKU_^c]<BTPe
Sd75VLWK6&(dEVV_84:EgJZ+44X5cU\5Y=EK.YZBDF\14Y1DU+1(U>LTTF=MaZ]f
9U6X8K3M;/MbCO;T/2\UBR\Kd2=+?O.\[TdO=81\a.aF?V[BV=cZ;]B\]C\TG@LP
/OIY5#@B@[B:\J0f:g2KUEKKD><OMR2PgK3DW)UAQaUAPE3V7F:0Yc\8I:FX8A5B
E+19O<1-/=BR9eaLgWO&+E]f<?[/5b:]W?0(ZSU@^R9b&^Sd7b@\@O9MeWH>@<?R
A,2(dN3&=0I4>N=_(L+E^CJf-@EI25R(,A?e1a;?#6CWG04D>S:d).8W:+@ZQJ7?
@AFULR9[E-/X^MH((2JUOb-@/?DU<S2/2Mf?1)C^>MP>1B,fTUL#<f8,DF0E^,JX
BNd>+LUS+-Ne?Ag=4Kf]LMa]a1R>2.\fR4)c-W\M/MF/F[OJe=WVJ7C_6M>VXT[=
<1(6aH1F>6/g#g,KA5]JG]d3072FLHEGGDR?;GMLWK?E_3V1LW?[:V4[d:-6e=6F
Zc[YZc[bgAfV;>RDY-+9(5QA4b.,>>WC@<:]KI6<DL;;Y);U#I@R51;gEHN:OJ/R
7-8Jd],8_Hf@/FeUS_U51V2#;9/]X2WBT7d4bVL0bg&Dfgd=Q6e8?c\7<DFJe(V1
/\=)UaS.g,NbI6K]]1BZ@/-L&CJ019(8f]EW;4_UQ&OLeJTE;C3)GI/.R\=0O5D\
>?>-\K597>70&/.XTAQ(H3-b,+_T;64+f#UI@>CPCdL(@aU[F^^R6IW<g^g8YZOB
^:).<AX+=Z/3):NBT7[1I5LN_MSJ1]FNgPI@9XQf?f9#=^TT-0c;:7TYX+-(fIcG
Z8OES^P^L2CHFcQ#&We_a,(7^DY0eS19[.aBMF3c8,Y_;=80:NJ4:<8E]86\-1A5
,dCKDV9A-@L_g<3/ZB+?aa_]Uf7>.#5[&O<?d3-F-EdUaH<ZY7F3DN#GaZg@AHDW
XI)&K?g7Je5YD\3RG13YJD3PcJgPS)+LCbQ:[5:dWSe@g&2ZMaAWA@J]MB#7eE+Y
^Q,=1^2M<1VgZ15eT#b?(aV,(SXg?O+AJ@X<;U/dM?T4-C31U5(ANJ&0H@?>4_1R
Lb9Ld3JM<4a/+^&3M1E#YB?1CORHZ7-G2VXY]1\HX?-9\044AK#K&[#E,[V<fcdQ
)+P]eW/bcD;+@/GCP5]2W\9=ZX[P]M.ZN&>[\9dT+E<e)OP4EC]?^^M2^;SRNX16
MZg1(G\L5HAZAJfHSC[:T-6YH>:eZ1\.97F\cR6K=aGN>-GCLHQ9C2RSK;2=5(O-
E)Ma=JMO&4UW4a@&KfG:Se9].;P6aXI+O@PU]A06M.bL]@._&>+/^>/dQS6e=?TM
>X[;])&g6][/Y.GN>7E?9<ROXf+^b9)E(9EPe@TE;+(DA^E=8MZH?HD(QF/^2(d(
<-J\gN^RAMRW[ca2#e_V0ce8A9>@&N0D<T>KD#d)g0;f65W7fO<]_BS^>gQBHe9+
f0K/0c=E.\/DYU7RJcX1D]fDO;+\1B37aV^C?b[:)98,K7<Zc\]fHI6;:XWKgKY@
&E89V9>d@8ffTGR(c7ggZC^Mg1Ybb3bgE[6.dTg,-E+=UEg4@P.ESM70HQe,Db#>
5GJHP\UEU<HQC/PVf2(ZB5:]4LF)7H0.QJZOfK#\Q=SE#gT/&9dD]e2GSQ<]+WS/
\UJ6(U<?N#RQOGM;Jc:b0J7<#9NW=;7eOJ=Y7fV37KZYc:NYUUM4SV;RJ02Z5T9_
R(1&a5I9;9U/S+Z=aF0>L5a8Z#R>K/M96e7RWOe9.5<7d)?ba([^\c2Y6H+d1X?3
K+(>UNXU0UKe14@;4G6?d:BaBVC/HEP0&XI&75]5DGBFe-+IE>Ad3V/bfE[M4-A[
?;[<W\K7EQ,ZL\Ea;B8J^:;a:BPEJN)(U,DZ1??Z6e/;e2Y=B2eOcR0R#aDIMg1F
F5P_V^&Y+8@Z8M._^<fGH>=@6]Z>P1PBfE)X-eQ_^Vb,69d84/;[-;7PKFJT6V+F
9EQ2(a,45J>R9fLE/8Sf,a).J7Q]7NfOF@f#_U.=UI/2-.b?YaR011TY\fJ0b\A>
\a(9.FfJ2RL^;I10SX7WC]ea?U69T0GL3e[7P;YRL1c+-VWWMWEH-8-D^c\S]7-(
XIaMdH^9+#//2JK</3B[I24O/2b?(R)+,#Q]1S3\KT4KEgaX>[[a4]:KUHbU/g4:
U7CQ(+-Y4;^CL0]W>UX-A]0GQ/7CD,7b0[8,-)3&0g<GI6(+2abAM<YBC_Z0&^d,
eM],4a,1FLRN_[<_BEW)1./X2(])O,E[).[6VY[IBTe2<I.APG(P83#H?gV0,RIR
H,W6EUHG_6g6/^.bc]6G&eBW_J\@>/[G<E/KD?,3DB;).[.1Z1OG-4:2ILO&87dd
CIV^_g5&a-8.B2OV\^8Vb/\(NOAV=3g@J())G>;PbL6geafMH>J3VX/]W_S#P-0-
aGZc)e]3/YeaML&/T\<&[]SV-1QQH^](f1SH1ZIGD]:g2e/fY5]eg4?a>a4__G>A
KU8>[5]dM^MM->gQc:PNWK;Q))GJYQ-a.U>eKCX)W<O-V1J^agK<_TXM<4QUR1(a
Q&6Ug<OM/DNP?)@AG0>NA-Xc6AEaDg^>(@U]/>3#7.P3>@P6,,I8@KE1MNc9RMdE
#EZG,7FSaX3U@PeWFPLXe-a:6a]=D),,Oa+\b^MCV0+40@/Ne+RW=OP6b+H+Z,9b
ZV-IQ_X(5&)L)X.@He#A=UV0ZF#.&<JA@;K2^#_6K._^3FEP<2)JGE=0#UU/:RZg
DV0A\Wg-8WHSGDTT?H_,1#YLRDO\I0[d.0Ie4SV3D0W9GTW,^fMN(36eOE,K+]&U
&&;@1B;<a8EKZa/60>7)ZL)0PP>X[()Q0aPd(FAe7@7,@\IK;Z1T30LCad\?J9C@
b#8BGE[L)P]VL@BG2Zc@.A>=FW40=Q14JO4RT3&JeLG6A,7[\.56B(L]=Ld&eBV\
/^:NaTF&S;6Y9(/d\NWId63J5>YMHbPK+3I4VZ<T18IL-[+1VS=.G6gEaLXJBMCB
YB&gWc3DTgG#GBd601gC#6Ag][gca]@\04R(3dQ+)Og,.#4/Ka,VL:M8a-E\CEQM
@;TR#>#LV_2;]&dF<6X?D6QEJW_?G/.3eWKT3aVW;ceL7MaO2gb>1]AK+HICZ6KE
6H2VR3:2RX[>F84:@;@HUN)2FSBORe+48G1UE3&=eYdO&_W>e<@,;5T158WMYRf7
Gf=YQL?@AI&BgFf>+RReB?\af@@OMLC5BSRYe>QGX>Te<??6<>2U#XP;Ggf=/UFA
_);2d;)^Y;@KJ.DTBgY3O<=b\>X9HB<cAG@-K>[O9Ya>8)0Gc)aN:c8RQIZA=Q84
G.dccB)d?&G>Y97bV_U]\dV^Fg&\^QVB_V#_B2b95_W^LQ#VRITK6YTPa6F@Y^IY
4cQC/5RJKH39Q\7/#C>4?PSK^?YB@7e.gO&H=>UVJQW(U+26N^8g19H+Y,Pg+N76
;SB_]fgG/=Z1OXR0F,9Y]BOKIc>80P>ffZ/D:ZHB,^a5ULAXF3E4a>WTX&DXGQ^2
d<.P(cD:P[YZUMUQEP>E^g;5KC[@,DH2:1OO@<@8(918(e.XY_3,c:2>E+/ZFW;3
#^G+^fU3-g)IUQH,AZ7e7Xf/MP_TM4/fE2H=SR:7bTfGCI7Q<0U0SN9^:4VC&dDP
D2X^.N,?eW4IcdB2-_b,8X+R3L97AZ2.d-)d2:#+-KFfU]&N^Af.4AKc#R]55O]c
[+N^BZ59/5ACYSA;LG3b0bY?9BbYP,G12]QD#VU?[M^T\Z8RE(W3MI.8XA.R;;EI
A5D/J3#3W81G,#PFCVMJ8E;d:S&6\_YU:/H^^VDEbE/#E\fNCCSV@&e:F4GeJGUC
[T-;5@+HLM(<ff/\.LdY?9B:D=,DcAYDSb=<fE2?g1_3\D[dB.5a?1JCV/Xa#)1T
?JPFD,KH(^WB@5<CNUPe;.#4>>HDB#61Tg52DcU]Wd-CYR]T1O>KHeb=#V].V<Lf
f@QJ9;)3TgT&V;9)QdTG5EAM_X@/9E(YXd)\,e6]/+BdIS[F@+Ca(dWX:14N4W?:
MHJ-RERFdabT4:HWMeE0df(WFfeGHCdHIDRBL-76358&+)6H][IO93ZDPB]L^a9+
Mb&4_\J\Qf\=L=S809)[c7]dLfRH?\c,#P,CE<,)aT(I-bUX]1-:EV>XXET-aeeF
J37&COEYJIG2J9c<[6D/a+LY2;UCV/47RGQJ>A2NSP/A3RGaYVbeZ^(c@FPOWFgP
WDN^]1NT?48-WgDabK4QN[]TG\<C]B]-CK/F2c+5L7.-Qa?7#VR\)&;Nag;+X#L=
gN+]R>/GH#+>BJ9/.f?UT/Q>1D\T/Y](N+?I-Af7\FXF+:Je#?HGFMF+Fc&)gJR:
(,(?;KRE+C<=I3V?8K-H#EYY,A437(//\CgPLR>9Eb5U+a1>0O96aS^X/UB(?&#7
GX(_HEDb)P^=+(>M38(.JO8aQ:ZMMNeRaG5GC</)O]S(g.^OdU-[Oc.&<V^HQ[07
STe)04.2^S/_,PCf0#Q#A086-7gWYIV-/NH\YSc;#LLXc:H0LTa,Gcb[gD+WA:+K
?b2,U(cKZS64&@.(g6f1[/:,P\[a[3,>G@52XR?,</DdQ/G9_8d<6O5(Ee3XDJT4
EG^W=?2cO_X5FHIJ(HgG#g^Gg9WH5YPR_Uc9XHJ+X5V>/5Ra,HTL_2Hf<^-)5A:R
5I1SUL&d5S&b_?=5M]?HIX@S=.6;\NY:B0QJPL:72NU+/BO5U1I@bN[-&AW3M63?
UN^AH-I]<DZJaDJ??220U?BG7;)>Q8-\]GB_I4ZEJ9XW/<.6EYK>;,.\#XV8VEG9
]=ePg54_[S1>T/JL(;KZ(aP1-BS96\N9=KVaDM#:?8]bU&,9KAC<7LS7IV:-K\[G
TBD4FTMKH#L<]JY4L,W]@71+/d6IM\E.Ta4eCA<:ORZbbB1ZHPf.7f[9G0OPHCH/
T7Jb/HVB0,PV+OPL,B\SMa&P;;W@7dP>U@fd51-@Zg#Z?22ADba/8?bD:[TUOfe0
V#-4LL6ZQ7U6[=(EP22BXULMJMf7?\TX_K?1B4b9\AICa5E2[Rb3;1C.&a]&eVXU
fTGS)aT6RFPSH@I360g6HF5dO2gD5b5]]IC1V,1&SJ(P)0U1g4458_]).^E:C21<
3WD>X4+Y6I^XE\8YJESR0_H7.dG_d<ZfR-5gDJFJQWBZ)5[=:KQ\IE>0f[Mdd/5-
C8c-M3R;V,=J=FJ^]22DLYB^Y\W;P2\17>>A1(=/.].)/\C?FGVRE2La\b-d:Va9
H]OA5N/U/J4g;21T)=dQ&\&R]&3C37@be4-gd+?HffH[4<W-5>Q+>EW?/.AZORCP
@/e4G->DS>Dba_<\\^Ie>3-SXA)&aaU@-Wa[CLIMeX#\(^#_YNKY-KM2=eV=/ILT
XAOG<:_P?.DT9bO#\N0Wgf&&=WHJ^b\^\R=&]cNMM0L=^G];<UacQ-:W1aODDMEg
-1Wg50^\FF;YP^.NG7[N(@EeA&P4c22,VM-A.E<KcTE]0d7@2I?VP+2Y)E]HA4PP
Z<]AYbdM4@2L>QD\Z<>eW]HO>&.fggE:K.CP@S0bVZ_G1R-BW::66-V[LF(#(fY#
F??##33CR3,aP/03X?Sc,?S\adCQd9UB3fCDH[B<SQF191F6@/6bYPELDDYWLfa-
]?-bZ\-V16#Y2;Y?G202g/B)deOHQ(gK9PVT=2e_Oa9K+Rf5#P.4L#2GTE:LC4&,
-,22]&_TeB=\TFF#&6L.F?0QS,=U_AL=6WGOaFPX(6J+=&Z>f^EJ666^E<AgI<Md
XQB]gWUcNT.+T7+BH(Lc#5BT=HW7YCW13Pa++#6:GSH..+e,CS,M>4:&A,0+=cOb
D<C0>fWF^D)2Yf2#X/(S9MB+\G#=U#cIDY&-gU?,L<(7<LGf@-CY#@[P-JX]G>ST
POZ\D-6<^[P=^;aa]LdD7FQ2IB8T/5A#?WQ_g16+38EZLET[PG##RHYC7OCQ;g14
U_NQJM9dZ2a#]Pc=NK5:aZ.efecFE0FGL(0GfFAMD?Ead,VXKD:W8BS1.Hd-VZ6@
&6_aAbI6b\T/3#;@3;cg=B]4&c#DMbK_<Gagea9R4JM=-c.2(65E8>6<I^EF]Z4b
J&RX2N;;4LRf=46Q6AaN@8HPK;7VHa<[CPQ;Qc,N(W&G#GY9@HQdFC_fQ3(HVOG/
V-dC1dSf3O[=><K]VO2Q3X3KG#9,/?)A1Y,@4E[DK-Y.F?C)MP@bAfd,-cgDAI2)
[V^:]1OE<&G[J]b]KD0=S9UM14<)Na@;Qd6Z],=N<<JGA/E?aIeFJNOGK-a:G]MD
Z-N;8TQDbLVY9(D31C\J=8DGN.XHCL@cTSZYDUD[DA-F+UK7BMZaO0<^VQPI@J6\
-,==20&V&#JS/)MDQ?K>6+H\;K2(LcU9Hb-[@-0L,9S]UN#\bLS:F^T<3J(YAD3\
.LAGP@QTTe(aEYZ@//HE^CIU=;:Rc((V:[(472S(BK@e8KAPS0OJfTAF3<8GU)\\
>g6@XAT.2;(+/1H>-9WK-W0(GL=,U<R2,Sb,FRbf;(YEN[0O&4dHH,7E#&1:0X;_
?L_PJ1H^KE=ea6PF[3aH=YaV@R@Yd,5)YbJ[fR.,LE;:/0(L__7&GVb5g<edF#Wf
QbVG1adY@/DIB^AZ\gTYR7?S0:^Zc3e8da=,eb]_AI:I.bcY.Ug>ULZ^,-YHL&D,
<&1WF24;VA>T(RMKegAM&g\MSgF/0NP6_285W/TBSHQMVW&@N)EbBP1X/-HLE)BA
>PeJAYT(VRVd^6;D@2ZL:M]bQ_LDFcZe;3[bN:UC,d=?AW>)dCD<+Mf9\M9bNP58
?(DYJ)Y6]V.HeGGUBSDI)5d:LGXdPR\O:I;PfAG8\+QA^#+X3X>).,\S81QM;X_]
9TI6>Xc]C5P8R=@JdG0#O4QfYV1QM=RVg75,gf\5C=U7-,DO_fIeaWG_[+^-aReV
]D\<KN.VX@ME_@/(A;5K2=g;aKV-+,85^O[9/GbB/YScZ:T96]C=Ce[CGVXZY-/S
_]J1L17Ia9?,ZJI5#:A63=f.Hf:c8L.Wg^DeXc90DO\JB0[\_-K]GG;SIbW2^[W)
#C;faCc04DS;&87TZ/,@7>8#(T11I6a]FFAG2XGI:[[>]J+AdWT^&#TTFKFSPUgH
?W[+;N1O,F]cPBFNQfYH&YT^8,ANc(_=f#8WQ^c/?E?7,6e9NY3_W>M7XK_+_91K
[VW?H5D/06<[XU3+0B&C5gcU3[Z(+#a5.c?@VW@A(@@Ic>?3fK=P;P;D.c^-0QN9
Ub+YUfcQ=JR=;<ffRaVS&A)9SE#P-?g8]OJ(6PA=6:T]5Y?X(7WQc)FCBUPa3b^V
3,^42+6e)H)2JG-b:@N@FQ^)[^HG/LVA&HgIK3X4/MMBcJc+Q?Q_8]<8]g.Kef,^
SgWHILKDGFMS:dN7CJH>K1^TF\+T1G2#1]Ta)4;\98EEa0&aAHQIY-T__[FF9G>A
.PG+DLS>[GB2^;WLYR[9>WeJJ+/KA<^CGQ]N0.(-#2gc0IF\^V+_&CRg(/@Y(3bO
cLK^,0N]1fXCP9T?\X>-6:QLLN9_If,:G0aUPcUN;,/-;QPaYZF+A[5KR8HgB:S7
IOeQH.cL4b,R:Z9:7C7@BN]:6I)257WYT+B/4-OdKY1O7DIAX@8.PNMD;)ZO3dO)
&VO5V];30Zd9XRP:N_ZeM5=&bVJA7GU@BdNfJ]d0.:8ad/:]N[d.N,<3g7QZO\9N
3U?P&&MT_P??abRN?S[X8g]./Ac1WJ7HE-/?,&ge>=5W8f&-OSU2?T?M7Q0QV>I0
>KZJ3\/(U0HCDecH&WfL<F6.2E;>_K#bd1@@e49UgUOH(0\=aYSR.)[VMTbMID2<
,J@JRUbP1P:e@)695K4)6CK#BMTK9dd5eUF=aP-gP<_Z6:+RbT<V>Qc:/ccYfBGd
3RE_RD90+7ZH_0cb-J#NE4^]a_9OV]c[EZL<[_cY\Q4MbDQBgfODQ&Y/0]ECaBXa
#[E^ME(D+,bQHg(/71>e1-LR([D<J@XMFL9NaO:Wa18Q6_33[RZ;I+d3EUW7+Y<]
\--HM2Q#=FQAECD3_M;4SZ_=?,0^,PQ+,U9]TP\R]6?))(@YT6-7+:61)0M^9c3U
A#X=g/AN?b\(0KCAX4H^HCfU1H4>a=DJc3JMWJDQP59PDRO]JC>V56Yd[/=GK#0F
#1)#a:5cT^35540SPd+WSbW\Q(2;);<_>O52<QXFN?+_ae]&O\D89IG9#66=P,J[
c25U_^3#A>#&CJ?g[?P>+^RV1NWf=6MeH&E.)dc&+H\^SB<ACAYg>T)8LXJFOGg[
^;47/M3#N3NGQJ^,46cG6@FN-(XG@<Y6PJ_)73AXRMfRaVKDaZ(.eG#?]L.L^^MD
17Rd];(>+44eV]FNg^Af(A81b7#<a-IgKe(;;>S8-W?]N,L0TgC]A(@(AY4=S-L2
>#H5gL&/Q69VfJ@\QD(>3([ad(PX^5_65YUSd9T/Fd0//#:EJ:I//69OdS9:Y<VP
f5R12Oc&/:IBDQQ9;Zd1:bLG/LC-_cbD[8O=UP,:A6?OB1(OL2M2^8E51JD5g2.U
SCb.]=^O^>UTd;.US)2U]O/1_]:RX<g47-KDK_faDg1+0VdaM;8\[^EYUW1BfZL@
HaVV\X]A&Gd-(T+\a-1@QF#WIU8WIWE.f)DR6_)f^[c^7?R[_.[:0B<9?NPGAB3Q
gU?\D/3EFE<XNB9OD].:MS[g&UDeG20cHXLS;;-0W.MZ]-7GT=[;OO/?O?(#H3TN
f7e@e<Rd_@9ZOLLN2&a_VEQ1d:QDY>.#IdX@5<M,)4K>gWXW-E8#7RK07L\cIEKY
=R88TFP_3[]?QG5X<:?CRcD=M(INTYA<2MK.+/U7.2;[6JOQ]a,2gYOS;&b#C++<
DcT)0RCR9(CgH9A8+ND#EOQ9a#F^TU=06]]48MS>,&=2..T?-IKaE;f2V;Y^[+gU
JA7Z[W:X/]R(5^3T.9P7&E2/606XG:Ia-J)L)/7UF3aGM.SGYZ]a7>C\-,QY]_OU
&eOXVdM.;<0P_+BL8/KB3/-5>V<_XP4[#ZLG[WJ=f6\<>(+3H6eN^<>T38PTI?Z7
.0X,Y;R[7451A8N_XB_(;/B7&@X\7&>F,]RVQK#VE/7K3?R;b:..7B-PDBZFJV57
.KSW39NUcTU=.PV<OD7IQ0#RH;^Y;_J9H-S&MMC4SU+)QSc;0?gdLY08,^RgK]2(
E?3aa4WF+0BZQRB<H_G0+YK6?>c,_+3+R_cb;]a7JH+e=.U(;N,.W7>],SZcQS,6
Kg@;(CQ7P+ed,.Ma(F1aONR\GA:H(#Q#GSd0NJ;:ZV8#4Q9IFWf>gcUgZ54/ac6Q
[__O++Df:O;e43:=&<S,_<,-37&OGG])VV.a9&](+D[G4eVf4WcU7(0V<PS6gg7P
FWDX0&ZG#=]AC/_M@C>]@+DSP;(.850YBg#IT8QH-=M5?+fG1aZFb<F)?<\T)E\C
C)-7gLH25)H/\XfC8aOFUP+f)fT3I6<BAOR<]6;C3X[Y<4[VE\P39/S50,Ad(,&E
aLP2I3,O^0,2]00V&b_MeaHeG5d@Z:^@B@F.)B<7LY3-fa)db0+=J6bM-O/B(\DQ
XNJF>&;/E6\He>L01BTd)DI&J+97FB60#)KZX3V.-NTdZG:5)<T+\P5g&PZO#67Z
:#8A3>BLP4U)b:(J=B/bC4ab>T9YR2Dc<ANc8IW</@2XQ]O<G8B>V2d.R8@31_HG
6)(NZ:Uc3A,D@YcFccP\>[0-WfUg,[PI<FO4PDA+.P=\::7?6SY+caa=JB5+RRLC
&PdBS.7,\MX_LLQfU_9<LMIH4::1KB-+[.[7;-:4UG@@F+\9L##-<MNa)&e_a;)R
H[QVeWKNDEXX;:K?@WI66@[XY71SX,HZG-W,0gXFRDg(=[J<0<f;e;[dbP&H4?;:
-507MgDZB#fe_>:4B1GW4V7dA9/K[gd>X4H(^9:Q;TI1GgYdJ1](/(a,&YZ[J@35
8;=A.+3T-541P\3A7O-OVR815E@Z@TI[V6O>-U6cLP1F0GDZLW1WAW4R-eS8e72N
L@&MI1?9XXdd##\@-g.:HaU-5AdGN6OD/f9HdU[5Ha70.=@0-/Tg#D)PS?B16@+g
a:XAXY5[b028Ob]<aQY_#BH]c7R^LcH42Z6/<>W](ee,5E&_2TQHB-;CWJcJS,PO
Y2CadEdM9#eC5.K.#eGQc)9J/c(f_dWXeNX2J4AFLOH980b@gg/]AE774b)dK2e?
]/R5VaFf^YDBCDd2+J/b3=37U8aU;d;cUD@50gdNK8-;J_XN8>e[\^_38XKTA9W6
LU55G5G33a7ea9Ica^<Z7E(4D(a;Kd-e-5\f?TN&g:IIdXSK/J]KR>9BQ)QH3[(R
5MH8-_+JQ859+HQ2:N^@_W<\LSOb;J,.FD.3-=8Bd(_\WVTST/O@<9@b/@7QBDQf
6X\)8KU9,2O>E+M]e(A<XdPHE3=.4a(R)9g8.[_LMa[P]LOf/JS19XXNKA1R8IE]
NM;@1&2,Wc^4NNK.):Y?aWI3_OKA-XGc>YBHT[cgBXV)BEDHQL6QDcbKU4?)GO(R
D)CX#_c./D#AfgT/(+.PDZgaG/368>B^dI(ggMID\6&R&YLCZbbF2f,6+W.JF0b:
:],&T732>YVF)QC+]X)\B2;H/^@0Q]/]R^7fKJ>UK4eB7[)Z#9,X?@B_L+4:DPD4
.])<JXS@([@Q;bcU9>W4<9E1TKA=.+@>Ge[gG2296HNJ.QPKe[)30_J+#DO@c_\I
M?4V@3S^YY:e4c#DV[]B:0T[[,RHV/ZHDPR-]+Ob,0CD+b8cd(aS+1D?0[ERS1B4
XO-\:03G2XKZ)d6OO_cAIHN(]OS5>HBAY1e)6&.97@abX;=G;6>^a11LK7f+)\O0
9M_-0HAF7NC=8NA72B=-c?[a0dg52:a^(EfN@883?HIG8<fXg<:J^UA:[6.@72eF
)e@>>\^-:VZ0M)3_J>>\SI>V60+/Y?U#HSWEd2RNWP1--+66gg\95gYUAR<T]:B&
T36gQ3d+(2de901F[/..M>-Z)aPdH3ML5FVVK+EfA8g5C+gA1IgK10.E1GHBK0<]
4EfIAUe@XVSE9\N8ZWXCG]UO0Ab-VI9dV^ULXe06]_V#^JKZ=Nf5:d85=9MKFAQQ
_.?MM+=CZG;CBeC+)#2VU4-GBA-<4,+EfRRU]@^@d-13R1I9e2gY@DCb71>TS#^]
a#C_VFA4La@H-\3A;g>69<L,#-MAE.a<MS(#S#78Z-Y.>NN7=D&JZB.&]S(H:]MV
2JgGeFI6^IRPdT^4FPe)RU2.K:@-1Xd:fJA16=PU24,BY]bU6&:(OVa(+)()^K(:
&\Q0ZJ9T<aU7X>I>W#>:>W0?5&O6\fbN39M=L&39dOabJWMgU4Ge7bWdB\N9ES;)
:X=\6,KJQ3AEePG^O.K/DGQCL>-fa=];ggLZ<>#E#3>ET9K]<HW[E^XE_eEOFBa;
<@F<O25e3PV+ECV_S^\?]ESFKT@=O0ZA\-0?P9LK9<([@CU@C1(-cPH?b?3Q>))&
6c[/g.CJM_f1WgTTLZ2[Wg-B9Y-(SXQH.f]g#-9FfI\a]PdO802#g/9R_gM+\\EP
V<O]&+EC?Jc#e99(D_K24\Q@S^(c=,bWda(bX[5-,L/a1B6/TS[PTF(K\?Q:V);I
g]Z^2[IB0eBISZ]6.\H8,68\29MU\5610^WIEOWfV2\5]#P8IN[<_D[=JfUAE=-e
HC^+CbPVUX8J@(H,cK[44,]+?2_Y9@=e=^d1_Z24Od4bCQcP8:D_<70R^_<<Teb0
71Q3^TGK/-P^aJ.9g\)JG@RZKAUH]=:fN1FbL&^:69;DMZ7<D[8#L2HI7/_T?\d2
b.--d>HE5-Rae8+@cH^)Y9D#=cJ75FKO/^;gD1]=/ULDE(eGR7ddREN4GQ^3,^;#
@>MPN]R5GN5a#ND/MY3b12TM>].K91e8\YHM\(#U_STN4#;@\/Y7&)HBFA-16XSS
BUaBeDRH+\XO)T;f3WgS_:.f1(I;Y)4SbT^DV<1^7R8#7QS8@\KQa^5LQV_RWdV\
9R<8ggIeb?F7/9fQL<<C-65LSM@^Q+Y^<X(:5\[_.N&Y5S_P:RC#;-GO2JP?KQLG
/&Q,+(Y\OYX+ZC5gW[/--ZI\E,.E:LWD?d.(U&fLe0KQ8dSMJO0+J]Y4-ZaY0N]f
&\SMV+=YH@.Ag^/Z,X7JVb^f2.53Qd<H90A7@B=8HW_AKD./L]X1.T+L_a9-J0]6
@O5eeBX,LZ=aKHIRKJ_aGP5]a^KGHW_4@]9g^V(ASdWO:Z\N-A0c((S>=.L3f]S[
DHFNd]Z@EJPUBUOT>X<^B?P<K2SF\]=NDN&<#X=_dc3G\>WO_/ZY\;14MTN:(?VV
G+(ANU0_P8G5@c#,Y8FAT^MNY9+^6ZeZeg4a3WdJY51M-6c2fERK62E6bT7KN,P.
HBPMa(,a0EF6e]/B=_b-.1.^[6QHN5(IL<W]4KVPYX)V+E.CFZa4fEQX=a(C]3f9
X=HMO18:65C@=O7P0gC?3d35(ZJ:^,E4]1QSE[(WaVe##(6?6,C\+2J(,L#@^LH+
,2ND;FbS,PB+QbJRE:XJBDT2+F9VS+V8Q2\b6YWOJP?@RKE8e#4F.df7&aZ0WDBg
7=:EXUZ:5+,5-I:0W/I?6OC@M(5?PNEG8NN>ZL(O@N?L763P<++BJT]&7eg#[J1(
\agXbR1O.=EKA#PDbSF+S9e182L6XLZ,a??D@[d@158R<#aI5L+L/f@]a+PD5B_)
^9EV.TU<O6L+P.D8S=XSbGSa]fO>1B3UPOcN2/^M?N/4;FH?)2FK?TcNaSW:;AHX
ag-ed:IY:.b+(72gW/<>CSOVBD^QS\1<J1QILd&6U=JgBYK5=bc89bJZX]B=(7(@
T.^<?(XN5g6U[_>]M83,N5c5PX2V8W2V^=0-c1-4+=N;7DY4M4LBX<Q5Td7TU2K_
Z<@>\=20?F^56Z>U(9[U[K;-ZUOYI8))V>,.FfX&MP/3G-GXSW>ZZDY32_dI(Y7A
>B;AUL&cKD=fHHYgESMVY:^GKN^=;U)2;\SPW80BZ46BJ)^#L@cD279FF=c/QE@E
;&Qa86@R&BZMVYR>]L,g4W2D3c#^L6^cd)AO6b0e2K\fHB#+732N^NY7C4Y/_KP4
9^.JaZgP>&M[2&Nd45T&gZ,TL74S.PL>9TGNH@aWVQNA9eAA=)2OY3\eZM4@FC^W
f#\aZGc>LI_V1[TSBR]#b(CAU;fE#/MOZ1dAEAOBT5Af@E1N^K:93&0U#1c/f1^b
geGVMCXMVH^MPC#]dMA3HF]1NIbKbUM/&RHX1S9g,WRCX3^0.S9A7(4/Q51.CRXI
@E[J33e(Ra=7>FTPeCV2g[KXRdK<-4>eP-.NGUA_ESWO6#,4_M^RfTDYJaE+LJV<
^ZGc=5E0de]OPURA91]M0bT1T(gBg8+I8cHN0;]XLT#A#20Td#6M>dP]2[T\OM-5
17c^d^Ha?,]adNP:(F]L/ab.4.H=Q,3If>;-2f?e=e+WbSbM<LR8]bPBMB2<9<A2
@@L]b^Faf?Z)0B[g6>,2S,bOQIBXN8H5g.R3)X4OZ;M^U2+F/J9\]^O+8ZG+SGUD
669XZbg>=2/NT[_E-g?_TGKL6>adK0A(b;LZ3A6KLWb\fg:#1D4F_;1&3EZ28.XU
6Og,QB\/4I_6GQD6G,JHM3DNC/M6=Vf<(H=/C+JT83]77X4b2DVYJWJ+@N@4PN+(
,C2,X,3Ee8#6?2D(TfIA&(/E>89cQJbRB0>VSAf;UcD6eO.X/.&8Z(JY5XO5U7EU
UL2U(fD;-J95B(96YI&)(>INS;gFZF;D.,??BF\-/^8YX:R?.7O<R1a&N@gbb=f-
42c=J19D:@&\V^/8J;X>L<PY5FbaJNAf[d>TQR3AdT+M)Bd<,Tg>XfJ:0?J_5V@W
HO-a(OP]DASAIJD1Q@AYJ1_b9>:NcROHOIS.C5=\]KQ\?/FJH0T@\AW\QVe?_G-6
2,HDBXJ#R<:9_+<f,/?;(S.OHAa+cS2\c2WW-27[EBK8Bg].AH,M2dX>(+H8)O6_
TFL#E;\M?c)LA5YZgf1@D_NOPLI0Ef\#eHXY[P]W;O2M[,N6G86Gb/dP\/+LfNCL
P6#8/75<VIG,4LeKW8c+T-Y\>_+P\_^e4gP4YWRd?;?+#Pgg:X1&O1F4->?(H>>g
a2a(R]E,]:;C8G8+(D/:_/4=-BI;;,XXca+P0_Uff=6NX_Z#\LGHJaRHSYGT=7gH
CK<e&E^TQ2-X<?;_5@Y[K&?Ha(LDgSU]#;:=)3eT.7,@]A:#:7]6ML+OBVS9fdX:
FCg;=dF;a7FPH8?:<N>MSIN[0-a89/PT?BEB1&OBK>I;;<.d#4FPD<>(4dSQR#4,
<WX+AfY-9d(\OaT[KWH)aN(KQc8Ud?ZgUE,2LbR;AeMg&Web&G@M@Ia1g9(T&eOZ
@,.eP-PP?9+]=\Y:K53M&W&dET;<OaCVT+X7#XW<\U/64\Bce/dPfGbQZ],1acRT
KZP>R--)gCJV)+]#8D[c\eU(>[H.7B;M:]_3;0;b?a)[DZPg&gE](&)8[HYgKJ#)
LfNH)g-@]9R9DH/6IZ?DPPc85;44a\X-JFXXI9K4PDf8?EKI9HT2e0\aOQLN^W1@
^c1VMG&V[W\)VOd:MYN<BR8H270A4[P2S/P:/QDYa&__)JUX^9E(&b7adLV-gWT=
g3G9IDVGZKWcJe_W&9;CJHE&bP+S5AcV:QG9P-ge/-X_@bRUHW5G:8S4^f/1-[9)
-e9eE+;>^P8E[Bf9<;AGX/bGKL+[B@<7,TY](cG7)HcD8V;OVCN;<\AB_^,L-/HJ
G/S=TG?74ML_@KfER4CM@;Hb3^GU/=?R1T(IQ6(]Db+.7CfMLd-V=RG8=U(>@+86
-94cf;6HH6_L9T0>Y6BF4,FAaR\3_3NYPX,&XV4#/TSd^]H9.89a;9Q2/UL&2[1[
I0JF:LPF1(2:J^GaB<VDBI.1&^&.\)4=-[D8OW,c^1K4I_^06V).=F5CBRQ;0__5
PN/ZDS8ZK+8b&O9g>Q8+@HLZY]6=DEYd6DNOWA5K8bD#O+&,b_e4_G(@_;e:3[cT
a(8<I@:VOe&PdQe9<IRR8Q9+f-PIeb9A.Q&VG^G?aLgH#K-CL/WY7<#CUQIG/JM[
DQ+Ud/B_7Q[Y0S9_6S:1XY.&KS;0\WXL)I[FC3@.bEF@K-_VX0-+K&H\Y(-Q_U]\
.<@Dg0b&;9V-_I,G]@e@Hf0WV.#[bUW[N1Gd\DD:S-:)>JXAbO;GL3b)ML]:#0cY
T6(S3/IG9IZc=/XL73c5fQZGJIC7^9#.?BadcN/]d3CBN&5,.F>98Z7f&@H?Y<&C
DGHS+@2Bf;B>4@[M3&?XNREaXgXEHeIT.YHa,MHUOgG,IV6Ve0DO9O>[Y#;KR@>H
eO8)IJB-5F^bQF;dIU#Z3;LI9SV]?RTPZ)).\6:<HSW<.\gHb9LJdcG65gY=^#,^
S0IPJa=XI023@X3G0STGDYZGD:I-1(cN_/4Q:)_S,-R4ZE4F5I[:1VF8P]4A.OE_
:]YFY(Cg-=8dC6]NcT(1BWIFEAPL0\\2Jc]Cc;Dg/?7/V,IW-4L0JP+&Cd;A<[0X
P^7_H=#=L5+f#e9g[.)\EOKNCBd]WND=C>O6RVbIf-^KV7RODJ@R4>fb+EG6JO#5
00)g_F_M2ec,Q.6D<HSUc1<#UEQC@YMGUYc6I\:d\Y,?fP0@K0O3+R3QB&e;\?D<
9Nd=-2,&9Xb=d?J6Q-JVb,FA.1)0\JVK.T#fG)-8G0<,JQ6:TcOR&Q8+_U6/IL4I
@6O83Q(b-(XLLKV-6cg-Rg-]S5>([C2WbT^K45c7dcO[a+O.U<PD94XD54CO>?#O
H#dET5fcaFXg9W>N9]&^1]S_EQCUL.&>E12VB\IEO.KP,TAGN60;Y:8[?BUWaZb-
IZ<+dTK>)2d<W#?[Xa17cK-8<1K^U?.LOK9OO2UXDRX&6(VEN9UAUSb:<_]Z^)Ve
TY[c1[Og42(4U/E\K(YgR3cF#d:RX)GSRBC7X^b0eANH0XRB,DY6&+fc7RUPg:[\
R?:DS4/1Qa)?L:@4XR&.6^[4715ZA)V1JDAgY@&#;bFII<VZH<(13)6KGc=LQQ5?
b6JK3.>6e_]^.WU3U.8RV]/.#0E+gVdf&<(IAaV6HD5aa5Z-J(X]SffeA&EO?A4?
e(#&RLL;=?F7HO+VWf8g(&UK<M=,-P[<^>E8;E,B7TA#.=fWU5T9-G:gDCJ8M3e7
I_B95IDS<>,P=Y]=1UUOI]GU+84B]DPWFg+(U4K[aD4>2aFINS2YT4IW=#+JP#[L
<S(&M7cD(18eFFQHLAC7E<AcPOF,ERCNHfRQ^3#8Y:\_7=_&/-30C>1<W5(LC^&O
(:Ae,7f;&/;g=\\5=A[^;Q-2-/APOTd261Qg#CD^T#LFEG=(O-FW^9<aGeQD8:e4
Wa9G@#]PHUN<ZE-VG-bS)0XV/;]OJFX[WV]ZMDU&88.62,9a.&U/B8cT+&KW\^KO
[#>HIe1&b\45IdTP<>G/<^aTF?B9.ZX(E+:T/9^2eeCJe,8B>\MUKUQ>Z349-KB>
&VY>Zb9F/&aQ9BA::N\gIUd86Hc]WAYI3/Veg:=Y7_Kd^RN3=\>c]G(f(bg5cE<2
S(<_d(f.&_?@dKeH4NSVUA3f38cQMO9>_A#EAaa6>3<,GK-?R9CB(A8/)3e1\,V5
248?D8C-?\=HUMK\WBGLY?3@3DgeBa]f&dK_5<2LB&0fMNSN#I4/cgTI[F8JJUMV
X:-:ef>gQK04R<bHEb2=;2P@+ec^29)_?(c0EP6A?Z_7.-@?SbZNLXM6L:_+DN)H
TV1=32ce7H:1e^BLfW7IE0BJKQ=cAPaMFF\];A@4P:CUVT>F>/HUN)>Q+g35MZa_
T,g^4?Y]W<<F<3d4M])1C5d]2]_A>BeaQ97=7g/XG?9Q-1bEd9K7=,K(g^Ae_X_\
C&UMf.8P8,._<S#:UX#ScT(?=KTe-K([GA[X)<?YB-QbJ[1E_4K@V9..8<P?F?W]
Y8GSK<U.333]G+1LQFN?D4UbNS5;1b.^5C13-7G2Wg(.0LBO>4?VT#=]D(If.T@5
J9M?3XGJ,T&>+E9L9O#M3/-K5:&1^;7g4J=U;0,3?ZLZfX2SHJCcTU9]ZX<9BNI?
+0I06/0A=9+U,baA9C1(<W]YWW4[X\)-D&I#84KZ:-@5Rb8^aXaYVE_-bgbfUWH>
NO>7/X;1I9PTVgHFJ_b;3&\\D\R?[XJTN0?dHV4Oc/9UC#\K2TK?0#@]DcTDF31O
A-cWf^@E)JdQ/P02>WBOB;TIPaaa^V[N?/M&Z-aP.;+a4#_A;fI]G=UJH#BfCg4\
_W>5\-VH:fNH7N^6_(ecFA^&bVA1&Y8(WHQ18Q,A<IPPX[]c+_>d8))IY6VJ5;I]
;RP=7(PRfH@E&:?&[0KP35J9fG,3P.APc(:GQF7U:Sg5/1.CCOGYcR-7[L&,+<6G
?U8CE92<@-NaUd-EHdJV\.YUH:G9^Y._DKI_^KKQ;,9U<ESadVNQOD9S1RTdc@eY
N(&[J6MJ4/LgS&/@M3dJ\K&?D7N/:Ib)BgO^K/:((]D;A(CIXZY.,ELB7O:)GaR:
b@@3aN)P0Q.@NEU:5&-^BPM+8A7Gg1L+.IG[CBMO)+Z[f:J?O1],d.J26@EFYW&V
OT7&fd2cDF\1G3gFPZCMD#,38:GYfK\DAIL.SIA<b3-c2.H(;+9S+8-KE1D5</24
.+3N]9>.afgP+..BHAW7/+XAFK[O+a+J>\K0[:P\VBY,Bc0W2=\\(BM9?@<aBGJ4
G]@6MPKe3DM5R]QJeAFESTUAV/([,B2,N_^0/B3)]V6=:87IS./)JfT8RJM.(E:1
KK&<(CNE/]2F5JI\-VcULTA#PKC);AXMV\d9HO_-LZd8E7=Y0>9E^;F;N):&7RE?
6ETPd#4dZRa-8H=?TA=ASH_2NIP+3-(NPD_TUJO2W<E(-X/eb/-g]U@)3(8[L-Yg
=80SCBYaT3.,L8dM..&SQ2WAF[]TMQU=VXX@Y.#0;bJ2ECB0N=(&X-1S;=b<XB61
a#GaH?YgT?WM6]MYA[HGFLGEM_^?@8Le>NP<[3\[PY+CNH]gU-G5(4Rf7=SKW95R
RaD1b5A>J3:b&;E1M/918eH[#BOIOgfb&V.]#ZG?6C8<g?[[;;Z4Z38T;:,].[L>
[=(<c@\IJMFO@U3@^@K=Ta3ebK@FBP)c(U>4]d/96JPKXH(f](cEFJ)e3HF4;f>G
UT-C>.:C>E?./1[D?Ye8]#S05N=N1K_::Mg8IR6_,<:>R)J=^90=80WP(c)4#OQM
+R69XC2+gJKX@Vg:I[P4CI1,eO65>62+dbVg&ZJ&VaN+/da9?3T7@TT(Z_4e:>:Z
R[.Y]7(C6U[+T]HOaFL8@YHO>Q<K5/C+_5JJ__P6PW>&528gW/^4:/?fB=-9F.Sa
-_T2=01Cb<8(1gVSJQ8OI?bcX<R)dMYBF3O=JLN9\4Fbg@g<L;^<^KKW4Ac=RRXR
X64bRJJ;4QcFUPDbJ7(?ccCG2TV1gKU<:368?DE[EL&IUcHg11/V,O.TCdf651fF
0a(3]K>g[;E&:0HX59/7FZ#W7,dGO_\<P\c9A\6J:DSfM.YQD++:WW;T8f_a[M[V
UC>,U)=60Q&gMI02\bO-I)5]Q7RA3c-[CC;6PXK7AbB]-+&4NXc@MQZP<a:7>1;U
B@P=@c<LYWVACQJQ#3\TIW/:9;&Jf3>P<V9?+HF@^6@cM1Q4[5PDbgW(;EbQ@M+U
MSH/b96WFc^.cc:7a)dU6GL4Y]JU7<Ic1:E#8^9GIfS-Y=Rg_1)a#X#YK0f.P(RR
aFLd,2,dLUg<g@@^ER<F15V7>3_-T6a+ZdH5XcR4La?AW#-fD2FbWOda/2LMVQ?-
c^-3_]+95eYYZ54X8^Y_.C@Y/a>210>E7IF&R[ABaX](R;H\fLB(SHAI__dLe@.\
>#)?[D3P68JWWME2DBQaYFME)G5:OHg(JSU\/FK,\4aB@71O(LT(V5CV=]FTX<S.
K,Sd<-9L(+dZHbEH2d.:.0K)G:8?P[U0-81C;&eD1583c[#O0OZ?TTRU?RdKCR9G
W9HU__DBg7\LbS4e8M\2aP<RT[Fd7Z@PHA=SOKZYF7\S)KJ:IXX1P)/X344@_@Ma
RDF?dC,a<d5G-/9c?Ob=J,Q2RObe//N9-N1Og19^0302/_M6;<II\?bG/]C^eY;e
N#7&Gb5)U09&b_O;/@VTeVN08\f\JR(O@eQ^R_c.D>]U&EKL@ZZWX.],UMK7a2##
U)\+2^[,TM>bA_5T=::^BP_U368f6BbMN2D/A0a&[geJRI]aA7ddRgX_EFHgEPa8
>be&(@>+QWI0/I;5):6PX@IHf1D6/WH#=LS9TH-4=#_]b[-cAT9R446B?<Tc2S97
Q.P5<Qg/-JP-K;L?EN7;DY,/cX#e<Q0R-YE+<OHHPaEX&MPFbM+6bQ_.=5R9_69&
eR_LPE7_4LKED-aXN^T<1?JP<8->KAZ0\;],J/:?+J_@K&FE\BO@<&E]RU6XN:H;
gfBdP^#VeUBIgJ0Y>bP^c18?)X13O8VSQ9HL\G=:fP;3+;A.e\[c?34D\<\NJYHY
?d]FQ^/@GL:b@@aGc#V=;bfTY^7[C-EFQZdcMfd):&7R4B0^R0/=AaaXb82<OAU3
:-7:,1XYa)_\11OAH9/VUMdb,?9O_6TB?Z9bB)-;ML6[8):TA-g;JA3MFKaT^Q]D
9cP+W80EgVW]P]12acLAXeGe.U^NR[cO)Y,7^5#_IW.UVQZ].NaZ4XX[J3?UNcL)
[)5?@_bP-Wd)0T7ULEM^COaCWW24.c-f;-7(<T)+f[],e:\KXFTBb57W-Y(^VW&T
,-EX2L#K,XI&fb(-.5PgI9\0)5.5^D=FXL_4)c0^)ZOV4V/#]:>/6YLF@bbC&5JB
W/34([=d4AWLf<Y2ZHLbS#Wb4=1+W?1Z.^LX3,P:/3H0Z.;.KCQW,+S&IKg-)]Zb
EBNK>faA)X&5dRX4IWHFX&S(808=G@1QH@5#B)_/?Y#b,6TT2#:4&bXKfV\+8#_^
Y)L=:T<C7NNA]Bd\?UJ1\_f0,e6<7VLB2M)=degNPDOSLH9Y&97NW[M]T.)&,L:<
88JHBgAC=3T-gRXX^H-.3-XLB&fI^\=_bDTTfAgIHYE)#(40JE8T6Eca(R8Rf:@\
]JSTdG(1>?\Ff>&S3-3Y@f(c\.(B,@-_^HB/[()X#^b0cIGAW&Fde59\9\6+8U/>
LKfX-g#MH8):f4CZXFfg[Va9c3V)2a#7fGc+/Z+Z\P;3;^M079)N6_AcbF6)R=a3
);?,F\YFgDL@b4fZQ@I>P.(-^2(-CSY5J0NKdM\=Q;;&(<WKa)C=>2aBH>WIS4/E
^_?Kg&[OOC<XT->?GDARM(&D(I,O4GHcX4>(4:N?ZBCZ:KfBa:XJPb;.]Ie-Y)]I
c;RXYe+^NC001)RcBZMR==WCD/N2QWIBRZC0?KS,GE>=aF_1R+Y3Va<V?FYV-R5.
WC/#b?MK&3Be2R9KQ#Y?)^C-5cQ@\XE&-+J/aKR+URK/\N+#B(&c8AYX,f<KQ-UM
O<P^16DS0Va8)S]Je+1P4T6E#<HNXV3#X^1g+1T)V)0C5Y?:/>>f#Lb2;A9>,:>(
P9X.N,#gZ5V>YBg0V;8<VO?Sa7XO[-I7JDHG1:;g]Y;HWcP)a]<2PWQ-.O,bbSd1
[:4?A6)a/2FP_gC8663E5_H/3,eX9/)c-ZcX+49Ic0_WNgS<U:9XL6UR^MH[RZI7
Q3a85-@)LCVT[<X1U]0a^^UX5OLJT(4D[U6;fN>+a4f_KB?LgWB:1<5Z?BT+)>3\
KdYO(V&#^cC@FROX+[L/:2d5M1>T2T@-EG>L[<SFM1Ce3eQHHL502+]B3Re)YI_Y
9_e^S&[RX/5O&0L,bYWTN\aH=#U#2:bP]WA4A8ZD/ONDEGA>Q42XFORd)_934WFN
AU.^7dgb/TXOdQc;,[Ye9M>.B,-32)&&YN?[a9TPH;]eOeEBT.EH\;WG_200^;&a
YOX5I/7>R157@@deY:6O8b723V,K#@,dC/,D=VV_fCAFH-3J44KL_,\BLbUE_RgX
3-eVIf(+)e?@dX0c?:]e7OE8\O=R-eZ8d?5(f><>OL2GU11+C,T5>e4P+U4LV-+Y
)aZRSO\.850VPJ>]X4&ZC<,K6SBTF24f,Oa2/:_eJ^QA_[;Vd/TXOT.<K,C<D<;B
A,+BNgSG)bO#Z)H?C;;0eX[QP/4.)-;NPVB<SA-6gJ[Y(@ZeK;6e+G=+FOY31?8=
GPKKN@FUJ[1R0<LB86_8FI7Ze[P<0(8fJ7SZ#L]^S,4S=gM7.V^b=6Z:TN[X>D#5
b]JM5@@1G/[[GQ[FHcGbP21&^LL8McLH@H=G&CRF+.Q;V8M(Y(Z/7b]>CZJd.-H@
B2JeQ;5U4E2+:)Tb:<:725_c?W/&bPY+X#SM)#R,\?aJU0EX;PLY.,DfPH2(]7,,
#cW)LL19R;T#WG+f-DVSL@@O3XX6C<)5Q8)GSVJWYfQX.GO@J/I6@N_G;JV>>20a
NJ4]&8.9;f-BZ5bge<S/+aA-ZY8e-\-?[,PDA-9S=0TBQDK,RU(^,#N63R>e+:WC
:]HAR],HXT&PGH-BE:<f9WN@gPf+,d)N-+/(UFJ++2;Rd^PEVZHN,AbT&WMU3C]>
dcd>d,QBb^^\M0^GY)JRCYb?S1Y;JccDJF&c&b?+#I:cdML,#C-gb\H<?/;F\D[a
1C.O>9=ZTUdIQ6SK.[(-@9>CI=GVIe9#O0TW5.SbFc#SOa4[L,RD52F=65d\Y.b<
fLfT)L2.&_DC\@NI3&WKND(P(D0<\BK\fY).JYY-YO@GeB.;gYYQSK\aVTcLc)@.
@I_MB7HcW4^/I-+ZKJH<a6.PQRX<)N[)[Ba+R6S/LXE7I:cW#NB5De>73L0?];=3
)YN2LbSJ.X5Z]1cWHR6&ZW993/:JN2TM]WBHR5W=XZ8LF1gDY2U^B]>KZ?7&I6>6
&P6E8LA^2+OgBbBZ@OFHLJB@J)df2g.B>-\+#8,DV)bc8;0d#GF&/=c-Gf2)T?]^
\acfa7V/Kb;g+Z&PBZ)e/dF#R0A(>M[SCUd^P8<7(]/.]&+H88\9]U&5c)@[-]_7
5QFGg^0JbN^aU]X3KZ-6V6CNHVRVWb]#E<@;?Y-bH#5IeA^HWd_N_NaA9&K^1[e0
QYe(DGgZ3eX-&7-3K<,D9#DKf)=6D&N>BdObGDV.XaN?+[=)7;_e14>Z6SfKV+9Z
C&:1XU6Z+@YF3f6M,/&R))8g@_@35A5#He4MCE0B/Y-Fc>2E-e8gYGNSODALR/4d
K62\cd+SD.&5CE]>T12\VcL&;ZNDWbU-ZGOYSU_2(@eQ2X1:.U<DW;/C6?KfKZg6
Ud0OZ576:B.HDDZF@f.CI56Wd@;C.,D49.[@)]B7LGcCF^f1UNI@N6LKXM,M<F6W
4a;JU&4N7Y5);7,__S,DJ^J[Vc_TSA(g0?R\8bVVAbE(\B#[/]839T[b99ZEZJH#
KTI8&_+)=U\BDL0=gF&Q#@X[J)9G,SSgd(>V,(KER;CF-=B4D.5._W6K&(T9465,
aJ>b-7?4\B7JZZcSQ9Ab.ZWRP1?3Xb@D8WOQC;d=3G,F.NgZ/Z;0]-@.6[dC?fU:
<@dY?Vc/PI]4ET][f-+G8g7)IA/8dcWc-72,=)A]eE,dD>6JcC4>D<VCc?XMHB90
(b;N.)/&QXd84[I:_+YIbdREc5Y(/.P8C42HW9V9+4ZdS?@?JD-a_XFR/X\dbGc7
accV0<GRZI)(Yf34FSP#<?KP(g++GCBD02QLC9Y((UP1DZC>DCMWd3g?,L[SW?9X
0a/54f<Hd@ebVfDRH[_DP3R>ge#@W>]VJ_,N@8IFE\2Id/_C/b-S&G=+?df4]AA2
P#E750=^&YY#d0F2\=Q0EfL8U48D7PFVN@VZ],YL>SO/N0)E0AdX)F5)+S3W7(/V
HW+1b_D6aCSb+a)#,/V\f[1C]D5QL8])P0-,Bc,aDd<Ycc16aTF.JS:Q]YF&TDZg
_b1A3c(S_(#<_-gKKWcD3S:TZKABMGC](,W6TB3V>bKPG0b_E7G/UK67Kf0c30R3
=(B.B\bD23K=+U&PQA17\7^(MFINe8SN]/604-;b1(8Had]8653+PY-OR2A13D0-
]:TE/\/D15@H0ITW0BM?@)<CGU<WTe2K:6RT<c?5O&0-OM^29(50_N\V-ZcZ)_EJ
[&[H3Vd]Pd:ZeT,[4)dP1M+e40SLY&B^OaASAfD6=bKG.1710HRXWL,<M<cc3-V)
NNdX;RXUTBc2PMOGe(&L5IGUJ24E\6>4E?_Ffcf=]E_775A<T5L26H)?/Hbae91U
KdY6<Bf-:AKX5cD/#6J]Y9DgE#0K+8EA]H.JNDbEeIIUDfHJ#&gcGP[dBg5&K3b?
.C5FPM;P6NXMDF<ZU<LRb\I/^Q]X,8GQd7\R;0-9+B/_D,][Gc-dcLDN:C6(Z6\5
Z?:NK9(/gV.0T+50aAWRA8_5DN4[?+:P)0e8D/0/Z/WCOBJ9E7I\H@<8/:gT?D4Z
d]W4eZa/R0PGQ9=UM7^#;TfI+bRL0;:3ZBMK^GD]-agg\(NTf<5>CQ=T3^7#2I=4
g1)#FUDYT@Be\eOgeO-=(^I[YBaY5,04+HAE\OYPCAISR=Ye]P7QBR6_J)8B84>E
Z;>_MgK+e12T,WFU6MN4(V870H8&E2_63+&ULIU.T6?HWgC+2&[e.C4V(LeNXSTM
3SK\VaH;YXfLIfB=5GT5_NY/2:#7?\:M3FGW.X7_S,214X=9IV<2?e>]M62:01NK
UNf@9(b?cg(c#g85RD\5bK2VTQbM3#YNOc[NVSIH_BL@a;1_K39S,4ZA5IHYV0)I
JMG[XDSD^dg)>+T^,T9E4FE:a7aF0R#L(_G0RO-;4P)+<-.Y5g;@Wd\36]E>=#)M
f/KN8;3>:-N(^a3#d(WGIUa?c9g_b3<Y92C822WaUB_>?RWdFR=V_8TDC;LG5-6a
+2NM7-L8ZOMd8NZP>MI^1cD&M<2\V7PU80B1ES;e;&2-3ea(S5&[EB>6;Sg;154Z
RM:][_4BVG</NR6S+K3?T;<WfcA@BL^)aN@Q#+I7IPPF+PL+\gbRZ11B?N@@=-IP
9#-\YB@0(P;\^9DT2Feb&:2X/4Q5X:dMUb7D9Y1cB=V#:/7NLeNNO-@E#]ZF(AG_
REf:B8<(F?:e4:>b1Q/]40O6=GJJU+[QT4?VEg]HWB(e2TONS94bSF4]PZ7;\,FB
?.961(Zc#->##(JYfWUcWX@cc39cMSNaQGK5V\:ZLfR#<9c+HM=>Q&Rg@5^.eE7&
P9RLLGI]ZR:4T^=VR[]8);:?NQ2LLPIgfSSGWTL#69e)I46QH9g>+UX4:<P2,-Q4
N;+_VO4_Lba3^?\TggQOFS^KMCRU_E3D^=KC9eC<ACUH_fHDgf@+Sf3J9]DObT(1
,Jd,BV)XFGORL11Ae847/)]41?@@N.1e#8Nb5Q/37OHJ.M<cVPT&(+T;.,I(f:+C
^PME(.490^O5eLHfS0;6_S^;(];gBE81#1OB][Y:BHD3F@,dfDHPKY;E[c^3B.WU
K5&,c>_+4g2:L#)GJPR8C_._UBIC+>DR3Sg-:20c_#W]=Zf\^cY8.fS&B@7T+A.R
;+0AgKfZJ&KT]M+5JG-+)F:0&#PLG=@-5J?2,T^J:_#EaWJW_.&M>@U@N(<D8K2_
We^3e;ZUAVP>3I_WW,EYfG<;<QMI-?7_3;);Pc\<7=.?Lfd?FFHQ\#gY6H;]9A8)
b@[YQE7.-OX4LDJNFMX4,GK4<9OH7M4P+IgXTHC8\JEGX0:FOCK7I=P8SFPEc&g+
a_f8D#9X9LP)Z;X5-<deJMDSV803K9RBc,QAD708dRD4V-+WI[=@g^.85?X)FfYB
S>cVP_9)G:4;2d@R6P95FEMg(S_)EVKRH3VYGRb80[94K;b6S):fW\8&B_L;0/#,
R(@LP>GdI1_N7L1=Rf=47]CSD;Y?CcRQbA6/;8^H,c35fgO>ZYFC,(BS]STDX1H^
/@\.^e5]4>6AS84RSKPeHM=.ME#SQXSfOZ;#ZR;5<4ZUMdX<<TV<++fc2\CB:H3,
,P=-&/_LZ75WLeGNA>8J?G0.KOP)5CYg/=8\&[HcH>:20+Y8DFF]A&0Ne7#3H?F6
R@&MZ]A]_3(6RG>)\J8Q+Fb@_GM.ZW^IV,9XWP3?J0E245YaHQ[?@0QI<-]d<77V
gBV^gZUbP]Q#PPMDcg@EO;+;AXY=cY\P2f#d[\&Y+56U(9f3(MSMd.O/KSf;(6H]
]^FRd1/.cL7BTLK3MN]>,F_\L))1.^OVSES,]2K/LGFDLGYg0R,[=f]-U=/1Ja]M
LffVTcaK[4FP/g<>H]#-c=_23GS&S-P7c>[C6UBQ<K:4@^I@E62Z?L&e=ZTJ]\@=
g&@([4BQdHCSR=4[_B(Kd[GbPBQMG(9&bcCT4[2bdA<B?fBB3D5[VNa.WQTT.G>A
QcM4Z/L:^?SE;:/TYV[9&)gF-OS3GbO98fFNN:L=MH4,N3>SJ1A5MCREF94_,/c7
=,05f(/gdNe=M,]41F.7E-&d]fFD6E=e2_;NLa[6]?0N,.(TQY5P(MPH1NDL0CU7
W-[+Q?c/#R#ZHVAJ&@Fc/QbNUU@O.;ROd615CDeeE<RAFB-4S8@daU_A(]gg,0WO
FC]&4a#@ZV^FdDP.DV40g@,,J6D0:JS2EBORUDT&Y9.P\aO/V>8aNUVf[a2Y:]#V
^-@d@A#Z;@S=PbAOC(cZNG0_R?LL.HQ5gVEF9>G7OSgH71)D=1+ZU<>Od:a=012S
fWcR^#QfPbU2T41@]JRAQfOV(?@#7VT^MG8I_Q>Q/He_GJ1KW_eXabJ)V_1NA4Gc
;?3eUE\28VDGNR7ea12C1L)FXd-ae)&[6e-C>IRRLY(1/3ITgbZZ4Yf2USH>[b.4
5@#=ZgaY.N<DI=G7T>6V(A8050>2UU&(;3=\M,DR89f\4AL:/CeT_I7@[&]1.;A1
H3b;b\eN@@]PY>G)X6cCd(5-J-T;)?<PVW?W)bd0+W>HbI@B&b87<SA(G,BQOQ91
_1FGE+2L;g<eEGL]Wf1c0EbVSKf@;+2L3I&<MO.STRQN=&?gf/OLf.J9^=_^Z6AQ
:MfJRYI+V,DS>0eK[V/>\^GM#&,;)G6;^<O),^QcS_69LbX.^3..;cY24<1EJN,O
4X\R>Va&^ecBd^<E[@GZV=Bd.TW_NH;X=,Fe_VE/8:dd#F:CPIRL<77VVX57(18^
00g<gJ2P]VAGL=g-?B,<7_QJQ3/&=Ug=Q[6[-FPDAF7QK+Z59@5CHC_I&:fT35?J
PLC<aGPT.SbJ:;(/cP8/SCS>L=X>B,10H6G5WO/XH0(]+PN==O#>IBdK?B?g>QR;
77QU6,?OBY@P+K^J_[bVZJEc@g@(=+f\8[()-\d<aDM_MS=;).?\dbMFDB(XCe#8
N,&W)g[8AdPF7S7<T.E6F2.@:db0.>A&@7OJDW5@719W3g=)XC][2\#a/5Y(4Eb\
-8bM^]U7<QQY#GY.@]Fc2,U75U&EfBfa;OdB>J#;4=F08I@JVbT<(WKL6OSGdU_A
Fg1RK1[JR2+9((H:UG/#2]b5f)\DOXb>YFR5dYPTUN>2_FAG0#I-^SR7P]eP-DD>
XZIT?U.S;@e_9O5_6#dKe/8E^Faa&5S_D>HBd<I)KK]9bcB^I6R/YDN[-J-UaR)_
US_gR)VX2WBHOa/H)(_K_(gF^R;1(4;bL)Z2>7^^cVN&gY+<>7Q@fIF/&#cJS2\]
<=V()S8=aYB&f]M[V7_HD&FROH)R:/V79F=DZ[\/dREAC53/f.aP:bW+B3):\XJF
-@:X/YGA^?O&)1Pfca^JIcF2C^#_0\\A?@:T[V;^;<XX39:811+#=Mc@3cGQ3Lb5
bLE+RB,=0M:DC15G/ae5SPE9QKX,S[g?FW6U5c-:NDMV2U]6@&,P/5^IAd&AfaNf
ZH26NQ+K(;B,EaHV3Q,8&;DC8]3566BOY@IDI;17HV?^dZX(5_A9<0;<#YAK8^-8
KRRUaFYT&g/6I9])[(\Ref#Qf.4P?8CRZdRSb@9&0;1gV?KWNGBDDKRU+B,[9:?.
VHT&&,aMPa,-W+VZIe&HJ>IcEU\2L>P)P.3W8#V5^B:K8a66.gY/dJbgMF=0M+dG
7CNcJ-(B9VB?1Y@H03,&Y,@;aWC+EVQK#Ze1XfB@WKNCJS8J2C)Z</EU?Af^K8R4
QbPSX9Z/e]4AdM87F/&&=PUS<,&f].8IN,K5OOP@CdP3F+G]#@(5(^#3#0,Q13>5
XU5Z&fQ3M,FHIKW+E1EX,6\7.d37@5\>UV9c-[<MOXQ)VTXR/C\-e4.&P,7>:VcD
?(>H/a>GNQ1M6[#:g8Q?,6ae<48)f<Y1:02Y>OcG_dM(U_SLUX^78Ub<_)JZ+Tg@
>f:R=W(70g.bdSG/4[+]3E+>M@^GAJ#9VEb,#]:1Mff+(I5@>(g-<_Q)BT6,d8dE
@-bd^T\DQ]\ABI#?^TITHR\fR#6[FIQC@4\R-TbXP#8D<37IeI2EZ_\WOb,#W:1&
e+]08>OJ_bV^ec^VN&8D^KK/0;EWLc\1FRSAW.gFE;7#<+5HcJ0J7B&]FI##LI?O
@?V9C+RP])SM\/VLP>QPgaTFVTY2dMRB>d78Y(1(QeK-TP9:>0CH^3JT@-RK;ZP_
-R<=F8)8KMcS;^@(fY2@;(IL5TFOcgX:TRd-+3E41JPG,=(OSXY?I2Xe07MN7g/Q
6@1NR7[I&U1>S8YPLdc26]Y[4b0\)YHJ#>XUS6G@&,0RE8PVUD=A7+51+2\-X^33
@=)>LAA=P<QOfHAM,LG3d+BM]WBZ##Ta\\e)=[d8I>fUNEWF-O+Ud&2W^5Jf:7Dd
e</5YO0@,[XBCY>WfC7VL\NBQ]dJK93?56.Y-E3fW4:PU?JYP7M8FB8S^YH;O:ES
V.-[Jb6JfQ3)0Z)1P#;:e8<=0Sf(:e\Yb[04R(@)9XDQ6dN@4FU5cU?G/)[/EcHQ
C0.bf\^^35KYDW#OP[c=E,41#F,(&[&b2+9_2PZPWI#M(2ge31,OT8IS4SRT:_>A
(3d7Q)?XUNNFUY,d4@;/b_FXB>g?&Jg-fA-O<LR3)3f;FV]bC>7@ZE6K(#]5)OVP
>#6&S[49KXc#Q=8GS:#7YZA9>2Y2Z3CQ]95L#_IA??=JIg?DcK.C_6/PL/RN__Lg
VL^,F5a6dYB7?#K3_J<+([T8>H&F()&NSaMB?5aQ>YR.@FbD4&302:T:[W,_VI/M
D7bd7BU_>781099\8e4-V\e5UNeE_J&?b3TOBg45g)g_^[5/8:4@RZVZe0PCfP:U
NX-R=aQ[_CRH8B:<IfB]_eQ8b6MKPde(3\-3/]CSJHb.V--<(D(=/#VPOcQMXA5L
SG>RH34<?O#@HT=7TUHGR>dUfX^M3+eL^H5[SN<ef<EKYKC0)KSW60Z?>;<Y@6=/
FE6>NHb[<3bIg?_>PM;,?CP4K-@WJ,5XSa-49f&R[X@HT>-+EZ_\D+ePCDH]_cIE
NXU?OOR4R9X?@J19OF]Ga\Yb@4S-=REcO1^/L9H=dT7fdR7a32cM5fee?RYQM+Z;
_cNH_:H=e8d&0QBQ0\LH/@6AF#@Q++=.E]gcO[YR.6+eWT68CK:Ua8/XEB70QC7g
P=D_bY/1S_\FdfQ\OGeQf0)9?6a:4AQc3D_X/6b>]/,PeW0^QB<.>LaJN?9Bg#L>
dCE\)7Nd?GKNKO1=#\3V0X0M0B0LD+bF1Z1Tc6aaU-9.;DL/E^Z3(^I,^:dN<2MJ
Q0Ib\f(<O_gVGD3LSG2PI7:aKGf7Y&/\aTBH(OQOcMQLZ?>S<[L0OeZf];K)AU/M
GB.LU80W1;.=)2UNe=,W6>1/]0#H.RFUT40=+/A?gOB&MCXQG#/&5BKDXKD(^FOV
>0JPP(<<3cT2:5e/LCX_^I0IUL_ESD.=L4;--RPfgdP<R^(;=5+/-=K65..+EV8;
]+68ddW6b;@&S-g4IfOBGDdTY..G^aGR2f9,_+c6Y-7W>@(:M_e1Q9BW\.&(??dP
2D]2@/5/SUcHf3,e?S^Z,/=TXRDO\e6Z-a[TE1Je4_+ZTRE3;J0f^QI@C<>@aJ0Y
dI)H-HF=+=5e;?Pag\()8-I-_9U2PU((GI\,8XV6;944K(-?O\8XJ[)9>f\E>IKX
++&7.g4Q(N:U+8Q&A0f59UQ42OEP?d(]CI.&Jf+0^\e971IW=ZH2QA1:YO;:.MS;
c_b5\;F#&:)aB-0/IR;d7\^C=^Kdf+-[[[QgU\.ON);ZgWeFT&\5C0<I<,9PMS^2
,O8#_QF,3R8K/TBU]BAWAcP6a)(=;YFbe26F.<S&1U_a[cPAE(D?&,NIXIT]Z;E5
H-d+M]Ye95O18(U^;N+ca^6<B-<NdFbIE<REY)UaAC(XRG]a\1UZP\4&K;5<:^LN
9R@YeHU7EeIZMDG3(>)B;)B7[dU[TMWFe,DaF0N.O^+B5/(DX?XP@.dM4-\ffZ@0
;/_cZ5CQYN2^6JDf^(BBLT7fE_M?@C9>(T1JZ0FX<E#?3&N?W-JYYZTb;2/CGMb]
1JNTbgb8U?Z?<#)<OHCCYA,SN(L0[8N=DCcS0dT^S=CD9Q-46Z:(>KYB,2\G>M/]
<LFB9H25)@TT[b#bG[HRA)71MH2=e-XAHQcYKcB(K)?FLU0?B=^67UCb]9c.A./?
af\U/#L2022[&1[JZ&e(L_YDb/ZH((2<A@W+8==VJ,\G-0=VZV:\+;V&/DXRPL6K
5=NQNg9RR;;g,E.b0YNW68>#90-YaaL_27OS+I#3I@-GQKR=8eBTT3N:YNFCCFPI
06WYMgW2?^/^,-YB\];8@)L;GcMf#)/0<#O90>La0HS5aS\8_9QF?O<13_ZVc5&F
E^Z7+-R8L:IX?FF(1YMc]AE/<<-3<H.DPBP\Z;ZeSM[=F\.2[Q;PUWHVPB@2O51-
8>-b5@<FcZYQ6_d91,9Jc_P#U[ZYT+Q+MIN=0dI9)6)fUReO5RUH2a_9]929].V+
N;&>g=(Nf;gD=@)FCa^2KZTSbG]d@7[KM8I@eZ[[a1:.1#QR^5bYeS^-CL3U8>c?
J3^HB=1]e>+NH\be/X8GZf+,_DF0[[41+D]JN2AbCZ9fLA24IdgOEa=7AdPHR.BF
C_/gXXCL::9aKPB[]>bd=OS];@/f4B)d2a)TNJZZ4)3Hf1Z-gJZFV@b6^bcddG2/
Ge#5EdEf=eKPdSCTGc8FG\/H=9UZJ]35AOgTgB<<fO^IIP;9#EX&d-1SV+b:gW05
([c9=?25fb)7Q-.39]G2\H0_+f]S]7Aa28:7:_#a0QQL?DI]SP>M2;[P4QGJ1e0:
/](P^#C46W;D&I4c36_N27Be4QT#V\5<9Z9S6H?GD@VNA/dPdO9c2bDJ]N]_Z]Q&
[#/E?)g4N5FYdM)Y+U/P:PI:#J)E7F;a>5#GIA[<aFZQ/R,DQ-f[\c+\#Z)aX](5
E;DQH1AWR<\,V9Eg_Y((4(T^JVf><6A?+A&P2+)2KD?]=GE8FEB_\3QT:&bX:V@E
R29f\HDa#NLKJQE:P16E55B:_\.H_O;A=afVda:0G&^de2RK,W)fe(dZCBZ-TL,K
N(@OcYNbE,;40JDaA^I>;W=K(>7FbBP:.XHWI5B,W@<M;WdQ\&)0bZfCPJ^8I@Vd
._/@V/29-__L4PJN<dUIFEQ]aG?Z:KB[H[ZOGFdF1ZGZTc2_:;HV&gYFS>?MVB@D
K?a.Q_M3.88FTY(c3A8[R9eCW:(VKaCa^e.e802SM-4LP^@AEebE;1Ve5F3G7GeW
;7RU2X7LNXUaT.bQa?1YSR&[HAR#YPLN./Z^LQff@+ZCI+PETQN2K#\Y,=XL4ZH_
JD=M;-II@O)HWKO)KSf;8YJOH1:Dc6?BEN3OIbgAg4(Z62KG/EYX.LOUJJU?bE+G
)G1eI(?Y,I/c[R:<R3V^:aY.gE>7Ud?2C/D:.(2<Qe35,eN6(2<f=:V\W&=S-RW[
]UPO\cPG?W[/>T=&-]L&1]d.\F2L7G[?F.[]NQ@65NI:fY:X?MF>0O3P<SP1H?_2
>GF=RR/0&[f:0S+Q>QbCB=Zc.^F.,M7A]#d/SS1^/aA4Y@D_Ra9&)8M;#7&<X6cK
R4-P1TId;-P(U1KG[5P2Rc2-UY=IC2D5A>W0(gLTV[0M+a&,@?3RY=_<c54(\fDD
-O9MO04[T9CXTE7dgbf^HTD/Bd;8@#R:FfM>JaASXD@OAI=b.MQUT>ga&-(H73L5
DWWeY<@^RU\OWMaSf;@#E+FJ(Rd2(]2Wc0\(?;f^bP&K2_;V>3e:<X?HQ.J1FG>:
[fU:S_A;RRFN=D+3>2d2;d6+AA@QX-0NK\>G],UZ>7=N>&ACPU5b<?_V;5Id8@Xg
5,e<6W_?CDB^;8QG3SXcbNFECa:M,H-N&)\TM0>GgU;=IEA2KPPINL3&/1aO^N6,
C/[DA;(a4A:B;eK_R-X=ce(:))VXeGLXY\;_S#dd9:HAME8D.&5&X#0d;XL_F+G[
a);X.0f7;_).)&-3P:WfZ@/ZR2GBHf9aE#AK6=dD3XaC/WR=ARM(cRRJTeSCU)4X
,Q\QH(^;N#N1aQ#D-N?\V+3KWgdVeW:]/2(EadYgTFRXJJ:PY\bf;IfLSCbC].A+
[/VSg&cES-LRVB(;fb]aT?XN-Qd5AP)e,6@)ggC<\dg1I3JcTcZ5OY-2<6#C;X;C
:RcBaQ1B-GU;aecY4B?_K=4#P/TgcC7+A\-ST+>F?I^GJ<=]^PB@ec470B/P#1^=
6Tc)O8^^2+1-5J9N379,(DA^6.:8N]b+DMP:5\Q6\6B?e>8L67fLdE4<^ST:LMN1
83eVO1L)^HJ,[+(GM,-ULYbe4E@12/c+(A3f]3cFX0ML6MZI7=c_+/8Cf2FED]D5
f7G,CS:GR(290[/.<eC:\7=]WX7V38_eW,@YY+gDSV7]HSE]aWYOb#9]0O4Z&N_T
=+6WeagZ&QfH,U3#16T>5gPJ:CFe(#EJ(E&6UMI>4V&b9:a+OcZ1eBG4ZJ<gPBHY
YXQQW6^_g43Mg,dFWU74<^<(L<(BcEMB65,<;MPIY&-Y<2<SXKG_G=#@1DBYIP,[
5]#acg&T?(J]8(aLfCdbI<>HE3RYfJ_\f\QDPOfaQ=WYRG_.UGXYGWUD.8;2.75I
EOY_3Vc2TPBQ]AJTd-1^]>82BdJO]X;+/23&&b^BU2E<L.CF=X5BfgUK>\C?+S2V
[)TD)7+dC4XcDQC^02\-Y+-db;.#O100:R/5DbRE2<0Z1JR],>BVc#GT/N79+4BR
JRD_UPEE((UVdT<>L\W_80]?gRUL7E-@S#J/#XI[+NF#>P.ES@4J1&SGLRJ,/e]P
8c?YE6&Vb>FP77agB-?c[bC0dL,&+Gd@GD]M24_QLWE+g3=5^B+b_2=V&/)c2VQV
Q-GA.#DMNF-.c7<]T[F;1O6^IMI;;@=X=,/_J4:/3Pa1D-I(;<dDIUIR(>)4X=_-
fA([XC9-/\UaS=a\Sd#[YafK.:f+);7a/Q.cBYIQed-/R&SL8T#fT_>+UPLTC)X;
N8fQ@?S_Sa:RWSQBVI?R_fJH@W4[K@=BAK,G9g\5)F])LYF@HM2Ga(@>#gV#P,a9
HS5[B?ReWVKK+^=Bd9M[)_X+^70c0W-bb.BdAc&<c#\B(S3f5:]-N>V77_:c4=L/
L(C=+9VBKe9g)A#cN;f#V=P#IQf]Q0;IFU<EJaT-;B<[KH9eO(A4AV^dF)]YGIe3
6.S5IN-N(P#X=\0f@+J1,4\?ZD1Fd/UNH4R90:U-ETgdGe@7g#W:?X,YI+dJ@.A&
WMN5Kf,6/G.1CA9U0F>2+BWDBQ;3OU_(9MHUT;4=MP]WL6eOe;2]Z.BDX,GHJgR5
S\(;68d]90V5WS3H(EJ\P&:O:\A#PH]I.QTUc-J?QS?L7Y&K#HA:3#-5d&?dG9GH
#T3MIYXVdd5fF&[7WU,LUe<OMc^5?V[=g6,Ea[P@<bXN-,M#e<T_3&(Yf\>)7+G;
/@0]+&NFDea)>,-/Z:W7JRUU<6.fM6Jg@</.83UMEMT1DLR973W62DfUe8b3T3WA
:DfX1F9#HK?@F0.aDL(bF0EK;L)(&YCgL?/b_Q;W5&Ma7e+1[@gGgL7YZW6(e1eI
;TADV6X_+XZMDf<Af9@g5[;A^@Q273\TdYeEV=<N?6K+CA4:Z8U2OZCf?9]XPL59
D>7+\(@&Sb-B>M0DAWdBIO>CD.1(HT\3-7^K:W,[fZONc:L.^OJDcEA)HJX:.E?9
fCP5]ZeD4L+Q2/bP;.dCOdJDQ6/d]g=3F52]W([103JBSHLb=P&fb]L>a#2KN/BA
cb0+)VaKaN],fe59>8]=L6T3E8WNYC@(Z1&]3FKbgb.R:LR9c2D+c7\;W/XL5VVJ
b?<RI-+TMIEN,6+8IO]fB+9WB[I1\SS)Y2P4efE47Z;L9f0E/=gfP2aAe)N#.,P^
HCaC.[6&>:B.gQ(1_<@:0@7GB=20e0IFWJ<3=<fPCHTD3bL#-FcAL?/Q1Q\]659+
3TUX^JVae@/ZfN-6L3C().RSDdBVbU^0M2N??Ff^,K5?>G-@SSS;I39+A2Ae4+&_
.eZW,L0f^/I(BXN(\^c5[deTZ#4)NIE^fH(S_ZT7+UAb#_Y)Sc:GQ0EeF.X;-,@5
62H=FFL?47dWJ.RA8QY\;cSK<7#<].73_E0UJ[Qg_GNC+.L0fF-_>DO_K/4;Q7I:
9;X[R8Yb13Z.\?Y@P-ERE?b)YMKg(TSHT\+U=:Jc-_3T@RSa#EX4=8P,QT4e[P6f
W0c.1Q)9Ha@@>BK79ML49Y]#+W)S65&dZD;I#?^d3B4d;8YMK2?##:M]X<0#[FLL
X3EfU;<P50FV+5Ra+YOC\AYd/MN[QI)^R29-]QgNB6^2:^P.fG-Qc:XIS(aUIU]G
/+V9f6dBFGG_JcMY[\3^,).fN07II3<dD-<c&W4O/[.L)Z>eOA,DWR1Hd\7.P<QZ
_(C^DZPL@CH:]XGV),M9FS/TX#F4#S;_g9@gd\a?6DFd<d,LMH(C,X-VC^VT/4=I
B?5LNcCD9MSNGG<U88]f3PDXVC\F<=?]aS_Nd]O-(g+fWFX#HaY[d,1/2_Q6K=Vc
/Sd_fa8EcTHI36E:2fN1RV)LR9AUY2KWJ[64a^>>/KP/2MR#KBQPE2\31=/eT)aR
BUTYRA8K8d+Q>#[0Y]MSaNY1U6>::[ADIEL<.Q=DAJdTU&4ZeWK^8<?H+7LaZMIJ
/N2F9S5)1?^8P.,c0U(H:T(^>\KEE0Y2A9;.cC,)U1(2<YAQ@D:HM?B(ILCdM;WK
U?2)NG?U&-Mf:>7EWeHO_KPEP:H?BC5EX.c)d[L@+-H6SZ<PU=UCV)de.1:@<1SI
cJ\_Q:-]1S_.1&Ve^J_=XLHb)d<6D:)EGfEF_T8+.(ALNN:^DP:#,K)Z#T;7F;Je
;PfcVfLA3\V0JS,b.+(W,83&W2g:[_OTa1H;EV3b5M0#6YPIF/eB?/Q<8e3J27&0
;@8]C=^.\2_[W?7bZFL&WM>7f3/S:71WFb),44,)><H(Db;S=;2M9Z&a7X(,OVFJ
#cQ>Y:_DD+f[f-6VZ:+H@L1ZG1dR4=C&Y[8+(gRM3IE^be>F]4YMASDf/BIC7aFU
-IK-FPUA70&ZYN>T]dgY7>@X79fXd<Ig]B8IgN>Yg8W)LPR\T_8AdaCUBI&gIH+3
3Z\3\;XO1-]U)O,+U_d[LXfJ5+0eg#?e<EB<@cZ[\Ocb?fXdS:+aX-RDTg([c\38
e13#NEM)-/&aGS>#fVDPXRP/b^[WTYOUbW7d7_R0V)UfBSQD\N.I3Q;7O[D0/?AD
7cA)0&_WdW/<4Iee9f.&REE/&2(UJ8gLLY#K+#FL=U=J=[bM6e.b?#6LB[^48-@V
bYY7<(e+1:R+P2#?2AX^RZ=PX_O(bE-E@DWHB?c2Ad^VVJ^P33CNe&4=6\<_EIb#
N.?4Ha]IG]9;LK\2_<&g\>M[V0<3\6)^WD0>[P8Y]0]?2gA3R&A3^5W(BM>1I4[)
?N\XcIG91M-RCM?>5PXNTP1T/J7RfgI7ffMH#3dB]W1WN_8VR+OfVbT,dO2?;ISH
;&SVY+5NJF=EeSHbS#JU?YbHG-M]KR;PJYW(A=9@(_7+D85PUFMKK_g:]+T<D0Ic
BC[cC(&31AN@YBI4TCEfETRg5CW;KLOd.Vg7WM@T1SB5:-;^U];OI#C/J-JS=d\4
d(@0RJJe&C@G6>XBBLXOF@,45_FXB;2E1g]R;E5dQ].R29#^&CW:bbB,[4Fd&^fG
>O0a)R2PH72MO_(W#Z8@90_a0(<N)XWeO>].dFWg-;DdLg-Y-N,]IEG>Qge;N?&:
J_fBE.XYF9;#,8N)5[-5RG\LR_d[\VMI&.?=LL5#:QfK_MZ<5Wb:HQ7O\QGMGPM#
_c(KZ/XA(6Y@e4XT1.<?4^FG@aeQ7F[1<]:a]WIgK)T1].GP&4FH\5KP5D+\6:CB
g:T#SVM&^>bBeY9ZL71]_V8?Y5)QcVQCGM2V)fS#W)4N#IYEF(;KDcH-],@2@+M\
Q5U<72-J@K[Zb?aQFO7H(6A;.VN++,Meab?#/#XaS:0X,3?LW&9VU?ITabZ-eDZ\
g?dbJ]c#Jg<<HH?RU#\3b)\/TTdGH@8H9/Yb#;YcVKQ]BL2[18FL0E\4gO8&@10f
3M0//bSP4Q:b>3SG@G>Q;K6W:g=,+d4WB)dT8^RLWXHaQ8W;E0TKX&Ad#UeUK#RG
cE6]&VAL;G0e1LH;6RJEZF3bM?9bP_[S?;2:AV/?A&+C?3=C0)73E#f.Z&Y@Dg,J
6-;a<WcP)1(03_-1,OBa;S@8\L;[TEIM-N+9AD5dafKb:L@YCa+ABS^+K+c4C^86
,=fK5L2U<G02C_LPJH_XI/X35d29SOgDYC<T<,D9H(?OA5_^dafR<N]Y.9f__4/U
E\_:BbJ/g8C3YgO-(SPC,fEBg7I09M/8Kbde]FIcH]^AfH#^NQ.fUQ>1;.b7[.5J
Da>#.0g,@5+C3?6^PLJ[gb7Y273Z)Q34g_N?@)EN8D0M?E_b3R:55PKc\3\KT_HK
#C<,QYLJTNXZgWa1U?FFWM0HeG@Y,S/8V]=U84JWO+P]0I78ZRR/_B@DQ3JK5,?1
TL<<1a2>[P(4+&V>P=L2ga7^L;#e)[gIMB&VY1EgJW2&g9/YCZ[NCAJKJ#M):(d6
L2ZF66@/&V;UNT]S&M+46?e>^B24SF)R8dF,V5/,]eRLQ_V1:_+,&]YL,M5I9?R^
NI711N=gVJ-XA(=VDWgC0VE<\fXGDcYEc()23=X+OaG9GQ)7A.1>K=,<D\C+5#(H
DSAPXa6T[f&.B>LJ:EHY;.C@VTXCaUG8GXbYLU+Z[W2#578,>bOLaTV=D<#B8-DD
4JRAXa7fB+J?03JYa_9)Ya+=41_FG?UNVSC=;B[-_RL&G4A[S.;.a88NVZPG7_@:
?BK(GLc,)YSa5#ef;B0S8f<Wc#Dff/MY=R6f6F+MG0JAfd#=L+Q8[N]e+0ODW:gc
c7O6bDA[P_gWId&W/26PbQE.?.4^=\#a0fDJ95-(.D6@^Rb21^1.XE3#U.<AVcYe
OXIB&6N37.V;N)\[6^JN3X8<H#MHb/,+5b&1_bSK<+LB\J;8>#.LK\PEU.[fF_I9
,+/Z?.+.S3](CDZ\/?+R/Dfe2XM20SbGH\Z6W;26F^52g+V@LG4J2ZYW,LTU:feK
ND>0M1H(18,a/M#6,E(X>?V_8C-&@B-9K#?\)_P=<:<;\dd6LL2M,=T25MJ1:,-Q
=NaT0<XA3K9E]05[=0e5]9[7OD:^A/^_6f[f<VC/>.dVd@b#;BDHJ5W^LQZASVMO
RQB)<0H9O3Cg=B:A?Rf:(YC9[VOeER+PYF]5,(R&/^;3J]6g@U?A@d:H1U/DCce)
QOIR+a@6IHHCZWYb,PKI?8XD@>,/^f;57#L>[FR[(aYecK,\+44F==#H:b[@f,R4
K.\aG1^BZ5H_VcPabNLOS+Ne6K0BV211^3@BD#S3JWX/\g8fI;>\>A\,/_0=F6WJ
-JCQHJX798W0GCV_+)1>L;cKa#(DV?(U7gU8=6FFSR[1:C]d7K#fcEDa>bRPC0L?
#9\^E+2P>NK6N4M55>_.+:]#A^Y)f;O_PUVX_-6B^d45c04:H).SDGI[YIJJ4a).
\D^SV.-L10gSG5GH,5B2.04Y5G1XE,9OfGEX^##_7/O6S^REMc^dGP3Na6IE./#L
^9K(fKHf1\H^^SWHY,H.=.XfX(0bIfHS[8RV;99@JgJVK9@1.K0RFYd9Z3I:.g?I
=0AWQMaXT_@EAJMN?\J.dOQ;?aZDNC#Ng^6_8DNB3^L73g.KE[O@5W&A8P+E_P5:
8&bGF/_RGGT-F-,dUSE]7N9?2&+0,9PeDKQID/7?M6X[89&=ERNUS<WZD-\\,.#;
^OVVN[MZD./e<?,LdB;[_G+(YaEX:(QU3K-MF77AV_A#,:W?E256(UPV_9f[^0/@
,OX<eQ\--/@.0P;Cg2J_cR5+gOR;[&_9LS&K@Y@.J[1J7C+^]@_H?HVVNW/;:fC2
&EK<QF,@,fD206SM__3)dR^GRLMA4=&O)CP+XI(:+DMdN20190ePE)S:[50;3f.G
00,#O_MF(E]@GBM^d/8CE/P[fOCc\K3(>U^a@1WVcDFU3MQ&UK<g._@a7:[(Q5<:
B-YV+)>IYSI#1PS>CPX1U[B&fP+(LXP_5?Hcg=<[/MgBX44LJ<;]WZ+e3a=fTEI&
Z9PT3Q,=A=9_)><ZW:?5_eHC#M-F_0>VX18_?<^D;<R^:@b73KF+9BbOT7E4([M(
eS[V+c7-fVI/HdX5_4[^[PaBa+aS)aSH-LE002MXAW&,_e:00\K@bZ?@8Kb?A^Z.
;QVB<ZFZAS[]5?5(<_=.+R95c?=4.O1\V:(.XI3/L8>-G4,++J-<==#I^5\(Z;@B
:SOP>BcO@<D&^\2<QG+/Jb?PJ&#=2V9<I:W_2X]XUA>XF7#5aW^(&FGK6+c6(0Z+
gW-#P.#O+bHA1\V#bZVEb_7=X9g7AHTXQ6gIFU+?WY&(I)[M.TY;[V(c]+&7fWA)
bIcI8,#5>24+)^e/O,aF^71<@<57\5Q,0ba&3;,3X3@c86ER@(BX9#cS^:@a)V?P
<[Aec35^(2cKIH]7aeQYFV561UD2)40DXc/#?,e,V?T<(:W+QF^+0W2,]>>^V4NR
QdXa6:;<A8^,@2_,UQ\#6M.c=JO#G++N.]V^L_c56L.:AYR&G5\?GRA7MQISa9IG
UQXD1b4A=SOZC>;<8bXSXZ3-CZ\gM\gASPf0L.1b1SI8IYd)87c?I4=T+\.CGP</
7SM0(FEJXRZ_09VR-[JU9@?Y,Y^MFRX?KSgM<+H,KSRCAD9-I-.CQeEEX]PU2OBE
KV2-(JaR7.A<2M,OU4aIH;N(=W;5U+Z\A[C[&,bE..218YNT&;=_9)_[MHe)>Z]2
LSWB]eBg0MDfR+?)<?DgedaXR.M--gd1PgONL10YRD.=_Ag)6-fL_3;=:Za#KD(H
(DPL239#>4^)2?F#GMDI2RA(I(WPLR\X:+)cAJG^XX0Zf(<eZHCb;=:,/7\ccA5L
,=KJVKc:<P#,8M/^H:4UU]NU0g__QH>N_9>2Ed)f]C&e+=b1]a5-MAFK<XK(D?0M
TME;DdN^>0=C;([DPN&R)H:.S-MV<cMALGUg6>cOF3ZDHW?_:T0DFJLSfgLgb)c&
39de\2VN,C,2Y15TN/HBe(WFc3OPff,25M_])1;aZW#b-(=L2RG+I.Xb+bRK\+6)
;R/@U9CAX6@.,f^6cRfaUKHCM81-O4POI&-QM@H6SXPKHM9Dg5?c1(d0:g8ZeFJA
9K4b-.]ZW0dgJ0Ff#Kb(:f;J+K1<P.K?YN^VUKWfQ(<@_a(Q7:<KJ#b)a3#2?IB1
dSIc(3+QXRe@2WS;D\6&eTEF#JN@7,B8Zb@2&9OKG\6#4[4-WM0dM(_^4-X0:8&c
SY99-;eeV)L&Oa1UH]=^,egES_G8ZY<<Z0@B<C-]^GTX.c.&+/G<;&:7F(A1@OP;
P3@-1W_CXQ1^>[ZEPg1<@]11fZ7.G1-D^/O67P+:+=UN>FB^#:MCf(Q7;_^PI#_f
aO)QbB#\0g1TM_S4]8?W.G-JcW_eW/C]=Q-LQc]3)=0a6(7I04CgNBQ_UFX5,/O.
d3=4+0L=ADd:]OZCb89FXNTd(&KK1NP;L,b:;TS+->R.=AEHBP-1;c@6M>dQ0Q=/
MM>1^-g9A=4;<]+^Ff_(=TRcd@g7gZCOPI;2YWVd4)dYd^,fAK4+0(Z.TDb0UVG.
B?QZ7LCV1a/YBfX6gSF9O[E9YPNddZMPRV3[AbC4E:bI3#VOCL@F0(?-5A,V+5R/
PEYb#(;_GN26L7+(OXb1AaWXV&<A\=0HDV\\.+-BOZR/U2J=-.cAD.<c.\_173=6
IbC)7aIaaB5Q[H(NcaaPfF8RfX:#3?A6<G<H_-XS<8OL4YK0=6KaI)QXGb97=8Ne
^J0Z:4^E/T@VNBQN1ML52U#NYQ=NXK.0&6CaI1(QCVLZED\g3&8SX,6cWJ1&KW=;
#1Te/9:VORQ>4Y.14.6a,=]0F2KGAOECM5FDGgSa=/^,1(C:Ce+7()Babf]5eacf
8NfZH]@PHIY67L(Sdd/]Q-KIgb6R)Z3dT#ODXVIZe2EaT,-Ge#@V=bR8V]dU5IU7
c>,:2]8L24.<JV/a[JMJ_7JE9#3&[SeeZc?&[SPZAD>,\]SEaf,aA?\7MdaT9>ac
69J>b<G=CcDW.GM#QEZ5YZ+aN:(/UHND;[Rf1@6KcB(@559>PJ;TUKg+(Yb]?V;=
(@(KL8]FVRP,4-?Va;/D0VN1_QgF>W8WXg5M=Z\&Pf.1JJ+,JZ<W,,?KfH[-O5/#
bCR,-AGeE-Z\aGZTC4F4af@-T.7c#4C@]bS86/O)SLHQb6V)VEN^]ee[)M&3Q7CY
]Z(.GKNBUd>_S[VIgSK,XY?=89Q(d_>C]\X[?,E_G)<#d4X,IZHBOd6[#QEQ_KLS
1:=\dR)1]#5+:4]ICJOH@_^GRFADeHe7^:A9WX?P:IMJ57NI912+7A2bSNT#PVJZ
JX.8LNCa-eG3,[T&gFEUbU7\gT<F+,D<;a5>O2bI0-b9<F2GI^fO\KG=IdE:5W+X
J5O2RdT.g/eJ4@E864:Fc&BTH[<=f2^D,70HbBdd1WJP1_Y&:LW=LF\DM_2L/d7f
fIId3&GM0e6/5OC^G@Vb.-NF(<cPe3W+N.ZOf]_QF?4ME?6?OL2KFCc:>671QM_N
-6VX70]1(\K.V6_b2Xg,[@QL>D@>P5:TDK+[>TG,9WaWX@f,?fF,/S,>f:DRJ^[F
QdZDB<+SRP\MRTY3L[RDPYb@b@J#AG9KV&LU?KC23+E^7,7)KN:D#2:SdXJMR[-U
^6=+U.>FF^c>:VZ7b)J2HN86f<0aJfdfd5GVKeZf5CNJ#KUS(>WKF7B>JET:0A=(
Pc06bA^/SSXd:()@gVL<+0P_A9T4VfdI89X8R.1Uf(#VZ)CgS=?EDEU/Z5B&K2d6
1IV<GS]RN^A:;Dg/AgV;0-LQZagKbO(UABI3W:E3RX+<gVEfY^8=Na]HBe9@RBG^
:?/,],NNF&HDIZgLD8fbILP+Gc-Ee<SBbGa5>d\]L^B@.-;5UHbEB8CYDHFUNg9_
:C,&GTJAc^MaQ<=eD9_2C7Dae4F6R;4>@-33R-ZaG4P](egP=6;Se4QLNI.9AT+<
5>a9O[W6=_UXGDICg)7OIM)9>V#A^]84F\dVQ\7M68Ab@UF59gL]<]5O9?C>MT8N
\@296)HRB6?eEK\+1eQ&E2[\Rc;a+^\4d.ESHB;YW\[1);[6JICPG6[)W^L/e\^E
S,O83.6\6\1a0&Ob@_^WHe6@CX&P29,9KSLbGH&NggP2R>ES^27>N]J#c/(E-fB.
YZ+Y4)5XfY_M]Ja&]@cP[]EcBeRa+U>&XO2#a;W@3f,&8bK_O[UX?:6ZWQVOcAcH
VJ5)bEY)SPO@#EQC8<.a_.S#;=DWKKBJ&P(9[?BG-(e9_ed2S5aM9=Ta,FEbR(-4
S)ZQB+\8R7GN2YK-#63U+UT)Id;.UW72:6b7;A1-3X=gG+.;\F+\gP-SVD>Eg-X0
V:^cGIPUUPTDK4FgGYVa7dV#;OcQX)c+,[0Z&R9HQ:0,__L.,^b7H-gcKLDgM?4P
@J9HG:f8C?BD>b01ZG.,Z^Yg+?X(D+Kb3=>aaJeD.GKX=.UbU<TAY(X[3(9TXEJM
H_)YIa9ecE[^Tc3b9]P^V,H:15A)>[aK)8:V;RJ6D6>0^[_eX03[<Ye@X]6d..S_
Oe2YWEF2<@R1V9(5H3#gP].K2bT9J&[@RWd7\Z2VZ>XJ)#5WH<,,/#ZN2X@++2/O
c^BfB5]2fN\S/<<K7c;E=+gS?.7MGVX95?]W>;M.Z/#30/7?D(\eBU45I[7d5^Y#
=-3W.]1<AJ==cF_<C\d#795^W<Q:O?],5E40N@E&9K:eCS:W4d-2(KX2FNQc20g0
W\;2.L9C\,B-/eL7H&-Q>[]W;cU;f3?a)=3BV0Z?AD+.<6NJEI_[O;R-RLKOTfd+
6Z3a._F2KFW7P:YDX&BG?SE@&GALB7fBFa6ONageH.W[1ZHLD[-bIB2^>F#cLPL_
,2^T5X9BM,BW9?eMR@GO[9<AcQ3_(gU2BT4Lf-EJ5I1YCAU^Ie?OGgB?YWa8:b+E
J\.a:[2cH&^,<CG<T[J0>YSZ^S(=/N(O2EH/gIKLS:Tf\a/YFQ+2@d9_fNPd><YA
A7@F4RIS-RK1@b./DJ6:LRQA5(E\;352T0<U[4b02@ZFB52a69G?BZYH+]T:J09@
MW\8R2UbI#YPf\a5.@B,-ZS).[7>]3>Of[FUcKc]f9Q>bD<RL+7VH/PF.(W2)^,)
9d6VP@F.B_aIW+@\/-S5Z&YW1QQGI;QF-[S?Z.;gC)c\47Ff)@d;:KO#-MZ7_5]U
>UAB:OH3S=>>3@JLGWN4Y[FH2aPAL9.5W-L[_,YV,Z39f1LN))34gIT0V_c6J-K:
6/&?d0e?<@&\PE0a;4/_39M=^?;XG0:X:A&I\3dbY8)6]<)bcMKbC-X[41)1<Y;H
0dIMT&1-S@\)M-4_LO0RDU&F2K0/I27NF8&23UBU9<).)6e=WLSD?.LLA?&O-]R>
8RSI&#?c5J^8,Uf_3N^NVYT.CPDC8dX/7XF?LOa#=RCU9g(R3Ag<BPg+FXZ7W_^U
<268AAc)BQCP\J#7Q5#GC0:O^_T#@0OZM?@OS8PADMHY>=;OBac-GVEObcd;ARLC
+)b6HM64;BN,NVO^NTQNHS@gKPKP-5-V;eC2)a9+/f@]1&@<C3a9Eb2O^ASdg8L^
^<:V^T5)KD4\CR@4G)cbG6NCU]JbTBa^[T]#EX]d@SF8U<5&Q/ZF-NI.#9)b\60a
Y.1^V/WW3A]Ng#-SPc-,D7^V2YFYbQ<OBcWM-M)4R1gWS67ONbCVNBMDR?4Ld6\/
4cH-FS?LT9>Tb^:S-WFI)^>QXU=XKE3+;A8f/TP59f,)TPY[D]Xf@G8[B[F]\+8(
g.\c19f&)c_1AC7@UXe<fN-9RfCcWDaM(IEa09eIdY8X=&Nf)HZ/0=Zg@HJW?eEG
b>E=CR#Z[.f/Ga,FTa91K>;JMVI,b9K8a.9:X@D4]B7O1BcC95abMJTVc+MSa-f<
KLI>-8.K7b=<3?BBfYA_C-X7Lc.99()?7A;?SDVB/dUR\L<U)4@BH=@He1F]3_C\
IH#:./&>@K:[aAY(cW7=Te@+E_]VW8Y-8aY3MEaN=a)WY+@MIYF&3aH3X;EL5PC8
Q-PAgPYA?e#+IU#/YM/GV_S,P)5]:R@AeR@<K.L&O\<Bd;P2D3^OK.c3[:HEA<g/
:7bTSFZaXLGf1]>SbU:>WNY_0V6?XgWF\d[KdY+I:OIY-\F/1ES:HaMY5JP7R7^^
Y7b/T6;[-A?E]FLbg/Z1d;2cb61)V55]&VFI=&@b\V#K:V.QXY[K&E_caPCHb#f2
JR71KP2EOX:DGK?PN#VD\ROVf7+LC&-gT3EPfY+@KB&ECgbXS;4J9P:0f]=OY)f0
4d\49L\>:_B]GdB756]B50E<)d&BM?=fQIKQ?>:Aeb/.-RdNZF;JA_C+5d[TfWPF
+X.2OA&d73MGQH7>eGH&B.34YbF?aLUQ<H_e?M1A@_cMP-,IPOA.JK\WK9d,>I&0
;Y4U2HNCD[:fA_,]0+6XS,7)\GNTT/ESMIZU.3^6LWa@,)ePY-_I]NLF/]fPP;Zb
._@>C5@?GR29@]6V:=Y@2c?4\AeD.cgRNd<dRT;BV\Yg840<5d87M6aZ5?JEA&[J
aOKXL<7JgXKQ=gE.__5C;3DeS-^:<cg[4HP\XLYBM19^6[J3dCKS?7-=U>CQ7K1+
MT(?Q9;U#f),ZJ^SQ_I,Oa/c40S,:/0=^.+<-<5TA\G\b=aWSEER7Ge)g+IF>dF?
Be8ED#/U7Y0IE/RC3\dV\Y\5Q&dG5BE&N<S<+1/D@]0bGG?RZW6,)X^FYGSJNY?(
3/\:@8da@B@W(9>YG=IXTMAbZQ;6E@QI:I+M^-)[6K@9=bOXa/;9a&K[eI9[H^77
HWLK>Z>OBKF:I?.O@HN<?>(]dOAaf[[-+@2)e-?:DPWIA),=fC015K]JP:JdCeJ>
WE;Ye#)Z8D9838N3d97C-dQe02G>fFP8R6Z]6T,S1cIPAE7[Fd,5NEK>_(2<\T@c
#AP-&F#79,WW-0<MDB_83V_+2^1--D>(gF;J.c1[M9O,3COB#-,La&?_GBUJDg/R
R6B:57TNI?a,Y6L0_-76#_=9E_UV/_;;2bE4]:Q0PFDHLdgd7]N;gXH00?_U+2b1
A(dK^@XceXfe8eUKBG]Yg^cB#[g[H>[[:-ZE(BC::.ga+#.;/PAH=/I3UVZF/+[/
1&A@JA/:6@9d^-f+7]MRdgIVRESf&^TX@fFeFH:1O^G#--#++=(>f+7R?/LF[#)T
X3N3\H[7?TA0dA94d.b\S1U9UQ)-AcWa0TR8\FX/+:LE#QS-O7[V))CJ5>PEXD5d
D\fM)^&0NH(e:)Z?G\e5)S.,d=2f]W:/@G^-Z)A3UF+4SJ,1dge?8[5>d(&A=>;S
HXM[5]:0Z(c:J#eZ<_IgW[EaFEV)#gC:Lea05B5:8gE5c4+08YKT]G9e,Y^Hd/OS
R.,f^(S9V)b4C9-Mg?YKQ:V+VKeKed[CK(7Q]4H5-F[V-4Q&ZTcXBAMRV,)W;ga?
-Cf:fg(6,<7]bdTY6WfC0@)-_&\3Icd.Q4N<^Uc8-&MQCH--Ce7\8Nc-[\NEHT,(
QPfAaTcTMZ[@4VB5^F6,e4TAeH&.VEC\g?)b)\96MMRd&9O\1LRKgXI;FR:@CLD.
C(LKXV5+>?_N,^;<N_8c>3=_:/G6?c,[SO,7J=/BR1OO;H0.=BX(DF[DS^QO+Hb5
]30O==c_B2;+3L6BCd>+gb1K6GPQ&@^aJ83]1H8.61=df88+Ha0+)#CC#0S411Q(
3\:GE,K0&1ONUJE]R9+bF-g?FaGd[487+>?&#df19C(P.5ZdbV7ccPfVF[#3)e5g
YMCYYPSSW3-aJ]GXK0P>E.=JFG1::OC0:8Q01#bV0#9Yd_df--N\<>XNWD_Z4gSO
?3_124RN:Td#8Dc]@30SAT]?/f1/FaTXM4S@95:(3[Kd.-\&>X,F^8GLgCcR\7#_
)\I]@(>]@Y_^,dgR6,_A;-C#0RQKAb-5=a4)+8><ReE6bBB1,a3WLd46@._O5(,(
-@2<bNZL9?4],J.\UEJ42eYC2E_YU-g9#g<#fG79:N2D1c^H:2B<VMB6fZLd.HcM
bN4<][3;c[CT6U(VOHg5aA:SO(-M#geU<9V<]6a2189J]F?]=YMB;];)X@)NNBCB
A;4NA(aV?(1@YP4?QV#CZ/?5]#^IOO.a>.bDO6M69a4DMcb]@L0AF2.Hf&555(&9
+2)IZN:MOAG5WV:&VYP#KJ+M62WBIBaC?D[K_bP^5RbYRe>:?@E(QR7&-,YZ_KF+
#KU5\8-G.W&,2P:a@^M2(5\PfdRHRY[(\&B4<0XVaXCEaOEEI,+5b5dc;4TTJSIH
^FQ8N6Y#;HHEZ6BaD6OR^H;\;[g16^0Y=1Yb>SAM_]c=;U;.,IP]3OZ=Dd+7GH7:
.cQJKF;6/4XJd2g]]:)3C_D11_OO)R8O5Ab<;8ZO[0ZBO&J?NQ@C-(@1&XT4KBW,
S-I>Mf[XZS?5)UR\SN;1/-I+Ec5&<RUUR--2@AG/Vb)c2V:7BAJ=ISHe0LMRGdMG
.RFS[gd64J_ZaJf-:8\T[L8\Z4RD+8(d<5+fM9G\6=Q8FLPaO7NW.29eVLIb)BNS
BLbZ1-M37O<aTGK))ZO(.fg6;Q#;FGJA16=/g6B3(3.3M8=CTR;gV1^:g_381+TP
/0#WEV1FQHCV^]<XWb99C\W>A6#.X>T,+>5E88;GTaKJa.U(CC9.FDOfYOBQf#68
+?&(/),5&QIZ[Y^??R.B1LV[-;eUXa_g=.RDbgM1]IJQEP7bd=AU_?5VaLD+J=E<
)F,AD-KdKADRAI[.ac516E?+IIXg:OM:gGM(QPU.J_>I=E8^J.I1.)YOE@-Z&H2F
^4E-IROB8dE&^RYaD:@V_@63-;H#+&M.;UBZXU(c929CXF),MgWAUC(\dg-5]G2.
VP]E7JUaJRc5]8#2@-YMKR2_>9:KX6>7(H1SOL-eA#_U^+YV6,O9<^/O>;WG5L+]
HQ+\L14SbMF=:<3L)^91N(VbA(,L?5gP)^Y_#[[)6#K_@A^cA_Mg[G15V1OL-;RT
#EbIN#AD5#/.A8<W1S4@HY>-6^,N@#=(ZQQ[I^,/\D>g<=@\93;JFW_&OT4.6V,D
eZ>S<c60;_K:;<L&CONc2[>Q4eZ6f3&OMM1E486KA83.ca=8f6A+5931[[W[f3>B
aO&.UA013ZL@06<Y&3-P<G55]A#\0@f&6/XUHbCgf)]QJ<8AEcS;8g:_dZERAMbB
2?&GBQ.U8)O3]DH,D]=MM3E7;G83B7XYX+ILH)W]7R1NKU68H:ESP>b\L<e<-e<.
O&0B49Qf^&)FUC)?7L6D;(OSd&:M_bAS^8D<Aff7H2]eP6;DP9Mfd7bbI&CL)7B[
\11?,[5)b4J><KdOHE.NbH.^(H3-5R(:cH?EF[A@-A^CWf4B71_GM?YN1@6OT.Wa
/MN0>D-C4SO;JH0>_P-+aSCE;9YAOVb]?KH=V6L(_8;BPV0[_.WI\Z-3(AQ,<6W3
^fVL3GZgUfJaZD#\#)NQ0dY[E@UO./9@QPU.(5S=UH90?OFPMB^<c+Q>d#gJ-HE0
b/D^FZP5Q;B]=@]fDY4J?F@WFBZ;2TF>TDZE=_GQd<<,P@/6S>J6=GSSF7_f_M\9
#WV=;J[ZI#(BME0Y=_);R=LRS4a(2Q)8>P/3Q6RXS@M</:G,dV&1b?8FU_D6R<)O
WfbTWIBN_b]MPMU-+E)Y/I8GL^dEfa&[(bX]S_>E\/FX[dadVMYR258FL$
`endprotected

`protected
=J2#ae^5S]VU<c-^ae37d(G]@J9VSe_NA869)XI>Z_eGW:X.S<1Y7)U)UDR4BRSS
[ge)QW-C>D#Q0-&B4Zc+Pa\MJ&]F.?e2?YO:]/dJ&__GD$
`endprotected

//vcs_lic_vip_protect
  `protected
Pg<e)T#U6,U)L,2I\A&5W]/Z-7(MQ3N;>5&e)ATPF+9PTTRE.LC&,(6LS:OLTFDT
=;7ETNW7UWFE#-cPSeUUN-+\FM/Y?#+WT@H:]Y^&XKD-VT0XMJ9U&;+>5g5<2319
7ZaCDN6MTc^TDY;>JFS_W\;PdP3cAe18R9(?11\YA:^YCC&,71P:_GdF^g[G,eWJ
M9fQ^dG:THA&JP6:g-dg##?IXee]<3FXe+(02FPfSQQ48IQ,Z/L.aYI7[BE;ZBc.
.T#QT5bI796WB?a3C-RYa6B=H9Y)g9H9,eJcaTP7W#3./QfKAN8Jb6(3c?;1=#&:
>gYfU;>a_Sb@+?SN4F?d6d_Z(e(F(Ha,X,[f6_VK#3fcN28])C1THH7],_YA[WQ&
98I9E3)WBc25&EaP02?_3a[UDOf0a#F<=YT^,JHF_P\69C(N]L];SL[=AH@PYZ&;
g7LBS(EJ(/VMS06C[USM7Z,_W>[T1B6_.2]@S2fN>M@,2XF@>cc0R6\3\+dJH7H2
.=N1K]T9ecJd-3AZ1gTYBBFITH)W6>6)SJ=_AT]_,9.D-;WaL+EDX0/d]fZ-O+TA
f[-;J+YU3U]G/=N(b2>LBbYeC+-H1CF7IN]B.>_W0;W#CDE<^;?2Gf9E9[D<E>>+
[=KR&ebH,#LW]aN)0#_2>c^E?NK0;V;gMU_+F07^DE?aKT_:B4O:P;?/HAGef+81
I>>RcL[Jbaa5G6NbYTC4B^_NegT&a(@UgTV?QJ0Q20WR=/_<&Sg9f@U_7L:GC<c7
QQ9AW2TE<L/g+^S.F_4g7^AUVW>gQ.9T@J6SZc7f/RX4DI[_[+C,2cLaaBWXZYJc
6BMG<WXGeZfP31UId^0-M_7@=J=5OI9Nf1XDGe,IFYJ1[>a\F&/ZGDgZg;DM)]>K
eREF_4TWA(DG>0:E]Z^3U[9T#F6,;WWID.#QMc#TEHe#e]4\>13<]GK5N;\7A;;H
_fSQAdXF_886c=CF&622++10L63d\W;J;B/<b^=O1DK4XB07OI]gZ@12^DLe;RTf
XRW/9_MGR4.Z?CKZ#Y_/&b^/K9,g0V:,70GK&^_X#>g[?.18](8c^C=T5V@>I=>:
bb25H<C1J#37<RJ)#(>1\Q__MSfKGA+fATQQ2F0:0@4^e6edE09@0)9&>P7Lc[F,
7BB@-1-&)2C>:0>/VGbZ?>N<A.-T<Kea-#-;)>b5MISO<WW;P[FO@b0YFUQL&S(T
K?FgOfCZ.^/R<,XU5ET\@8ZY:A8/[b:EA>]/2J95.A=8GGZ7ADCc>a,GN>Pe<<?g
90V;G_,G(X4(I>2TLH+@/61)Y?D&=[)bcLTPgaH+VZZGbP98eBa)J(5RD=gN\/:e
+>;9d,d^E<ESJ_EaaNABW+MO1NL@<GRH@-O@Q^5\GB?=/O?:UaL=&GE[H>B7UL3F
V/\<g:_0dMfeT\SbfS)DQ#P4Pf>O3IK(()S2g?eQB7fVJc<6[&CTGEV69J?K;/TB
+2Q:_[21TOM4=8d-EBZ?HF([49G(8ERV+7+U\J-CY5:TA[S:8@(<XIXZ4E=(G</f
-W(8/VMac59Kb=TMX<d8La^).b?9L\@KID/P&Q/@8b&#8Y2/T-HM)S-gAA\S^..9
B^Y225@PS5MX-E^DMYC=B<aL2(OT(9f.CVg:H)L;e?ROT\Z-);][MXQTT_#9KOH#
F;Geb@OW>N<,aFUQ<aKMYZ]f9?8UKR8&O0/^P3Y[c\)G)?XaFU6+[a3[Xg?N#BGE
/W4C7a6).d=E7@^DFW<6/\@-K^5F0^BF,FNKDW^OQ/)Ug3UI=I4NG^PHeX9W06HG
Y>ZMgCdD?/gNVQJ7)KJOQ=>I><<][bQ4@K&fd?]253Z^>W2(O@_gWB=/9gY<\;5[
g?&HSgL96UY7bf?EX+[Fe.,,L?8gLX&TeIFT;:TXc_SOAXX9Lc0L9a>CdQG1PP^&
D#fE?XWT3)G-R_G/aI+-4[G@fbe+f:Q6_7PNW@;98EE)#N-d9FON@#9e7YE,W,:T
_B5<XA>f?3I7A-@O7cEDffXgfJRO&e9]V@]1?_ZOSG+U=9f#&TS_?VSF4.YMOdST
AZNI&(:,04APGS-P?#7_3D]<K7M54?KM@f4I;06JgDO\_I,eW6f6b&(UgLe4WA+T
(SNW0<I7(3Z?C]<SV-+Q@fC.f;0I?[VVd\#QT[QSO6d#F\f,0SDL6g-LW#RDC(S2
\a;Yf]TCB:CfU_N?^ZTVIK&NSLW:.-eAS;gJ:F0TBGH=7a4_AQ>7AW>NEC2.?G12
NY5gP]2bad407=[/:F[8:4U.Q-]DM#748E_PCg8#0M@D&a&>E?[4?e>&5aV6@242
6&F9UM6+3806;I.a9=6A-7U<,EY12?OUAa4;U1g+=H=97cYZfg<G_?@^>#R60(7N
ON:[e1g091LBYRgN26?;LgO9cD@W</57X9WW,IYWA^gABIH)ABd7ENKY>GJCKIOC
/+6#QT]C#2S_f#AXeER;X6Y3LU5NEcH/I4UT<DTMMQ?#BZV,Re>KF:#09.\(V_?&
dfL,LZ0e\Uc);[0WGE^Q+e[NeMNB_<6V1AS;.[\\Gc^5]<81@&O1,+WF<@=;K>]^
D)McUIKD\8TTU?THUfXLfa(01Lc>)9]]6IS(COGH)=6ZBWfgcV^U39LX>M)6eT-J
,#_\a>+:+]cW]\[YK.dad.:\B:.3,\S[eB&DSUSH\G)YbFWH;7V.#5b2^,?-:gE/
U^KeB#V9YW9VUbd&1N>DYca(.;S<Bg[\=12-L),43IR0>RgCLc>.;QEI5^K>A=IW
4/W#]X=+>([a0C22#aJ=d+X/TP#@e35SaL(N][M/8O39B9HFI1)YG)DeB_CT_/YA
JeXL]8I,H,DX7F2agR&,c#6J7A1<_Z]PURga[<@?0/f/IfJDN_D/_XI&c]/R^/@L
dY<B;d++#87]_RELg,ND,_J7-@O<b:6HPd(Ld_KLX\17]&+G9Ed;>1/Q6L]5?8Rc
J8KaIES(-\U,E@cf:dN94P4;RK,>9<2-\fc-:]/3\MF.+DU,8ea;Jg(#16<+cJ@;
a^SL@0Nb@;0K[XV<=dK<^WC?)FLVJ3OP,8#aU]Dg1b8Vcc0c06<d6_BU&Wa_fSP3
dWEW=DAB>[4<Y2W\&4H>2Y0G]PYdQNHA&V:FQ00^SdFf:(IKC3Da8.;D;H<[\bb+
cG-H^Hg)SJ,K:\3L478,>TF#3TEeg7:+>>JH.30_@9+M@<5N(Z8/OZOdRTG_,#X=
Q\&M7NV-W)]][NYX^@_.Ub>6@X+5Mb)Rb>V-^2YAZ>1E;:5Ca1V1S,5fLf1[TB:O
,I_)6<B#F\6g(;?G:=JMFLU<-Wf1=HH,T8B=?V0RVX(,77?#EA2Z3QKBJL9OY(9N
ebR)L@>&<(J+?I@:ONF/e)7_0--Y=b->=F3>IB>AEaVDAEe,+M&g)0XRD2W?6a:S
C=-H4;=QOdT_I0K4[DfU#__[X]MY#bI6Q]4BgXA165&(a>F>6HY<Pa?^c7M.GReT
K)[g8CP[P:e\e4MTOVSUQd-1=^f8Z:_AHSTC(W18(@@d_,1PO0a0L^[K6XU^\+&Q
Ce>QZ,Na0\G[-:c7QM(SBc0UJIE]=4JdW2KIVU:@eZ6,a18@aBC2GHIZ:STLG^_T
M=W6RBDEV)+;_>PTJ_0>S;3S@TbLGd5g.1==VDW@B;2MQD:.3TYVdEOg]S7F5eP+
J3(M1MA4\Ce-cDEdd[E?g>Z2=+8#.?/^[K?H>YD;S07BGd(K7K)_I(QZBUT.J?H;
K64XAW;DFOBZP17&;UV^+3?OI-IBFE?#7b5YCSB^&.VCOOY1c_Bc@SJ/L95Td-S,
4:<+]RgX\e,49EcB7b<V7ZM5f/XRPI-bPOMI)9?LU9U7(1d,39gDX35?=+V7K)A+
,;L9#]TJ4B\f>CTNTS3OH4+=DL]bU6T6U=[.+074&>DYXI-D^KV[PA5OA_47,S6V
@L2O3&V[SFVX^[>]?35M15]#9]6]a=g8U-H-5K,S@QY7@FQf]<A:(1=EAFYd[=L,
g6H4\eHF:1/@?FRUB^9+eH\WCb)8.@IfBHFBS^N.V-2QNA@)9)N_9>\@.?\S9Z\O
SXNa:QQC^><J)eM>>c4+/,Z:^Ug9OUHeQd9;,F3)61W0bBQ,2G@e(N1HVI/@AaIW
0:Z;(Q[QP6aE1BcGA7_CX]W6A,<7Q3N)fCdQ1P1FZ>bC&5dC&A+5bNQKQL9PEGOC
EE/?A>6G+fM/NVYIcQPU@?LNRQ=cf@P&KH6ec\Y21(I5/V8H]ReHSf,YgWH#)7BJ
OT>QgVL+^B.g5?9O:XRYKg9X;dK:@?a#R?[_[&H-LUZ6d?ab1X9NEXYCY^3e0EH+
)5CL[<Z9Mb2]f@0OI[]bF_62LCX;14/[&DJII6M-_f.&]>LA=N,GK3K1=9L#G4NH
XNT6ffIVR=7#[&Q5;FgF&-A[(_WF?)<8=)e[AbXEfU7^#S^N8]L,?<R0I3dFHC:<
Ka)K<<:8Ad;fU,NG2C<1;<-XC.ILUJ?8_)E;;8&?,#BDO7W8/BQU),_ISPbbQ-Kg
G.0VMdL6=,;9b]a&]Q-T:Z(?c13_)I\be:6/f,^2>8_NGQ-9YB-D@_EC)8c7ae?=
G1P.TIc4S]a7?I4LcAJgYO)]5.H[P(Q\C2MCZS:@_UPdI3a+Pa&\d7\dM?JD@d[>
O\D,-PG]X8Q,;(1^ZN.:c7&+Q1.)JJTEG:A7#Z7PX3?.@9@];#[O=Wbd@fPge[(B
3#+e>Ze/fE)4-YH[A2)g/[V^C,UB+]XeS[9MAUWCXdX>c9_&6eBT\A1B,5QFWN47
9>3C#EdgF_7C3@4QO>G;WOX<-WfLJD>FXd6FZTHLbCN#.ZGN-\<_7-Ff:.^-:^;1
,15E&EB;?G3>AJ+bRfb;C?R?M?T5\H6JQ,?-]OcSfK/(NbG)XUK3:(+?Mc9N?_77
;dZ?VV)9GD1<E[U&_ND.?&/B&4(&+J\:f_P8bT>8VBW>/+c(;FV9:cO<<04b+FN9
N_=RI:eD?G@fL6:V+eH+@UJX1RU2K[C(<N:5==B,a)&ZV=Uc[^>Q0GBMa[_@UL@U
CUG0fG;eL<a:5ZXM2Q21Q\aeP_9U,ENUe[W:(]/\K?Ya<AV>YCD1S[>fWdJ9aA_M
6YcgD,_7QBF[KF(TfT>\cN>WBd=/F+_fD++T[X9..X>J_A-,[g,G9,3c+-^7A=a(
dNI9D0+&?M9M;U3WSP(,34Rd=IWP.e0TCcUROF9C?UG6_U2WGVS-#+YDd0T=&/3/
CYX2db/_8ERJ[XWbd/^OZIYIQSbN2=,FO_9BDT.2cM_Q=>^e#F?7)J\EYI3QRA:d
K2(SOfK57V,2,cW3Z[6W^J9..5a0&FZ@/3,I4+D#0P?;Q?OXHYaRReXZ/g_EJ#PK
;T<fT)=DUfAGH&0\[HKX1AbBR3LZ;QY:g#727<._b0&N[RMBW[(US+cYRHcJ+e6;
4QL[[71UM9?TLGEQ;b7>W.,+-3C0If;2:<UU,dT[Q#WN\]cF1dNP?)dc).C28FJ.
QHHJbePF6A:V&=-#ADUbcNOC[TKX2HPBNEF9D98^g,^85R(571(//MW,B-VcX^,F
PTgS(&gQ.TP&@,[<\Q55(.I=McdOA)-=&2Ge&R>_62DSN:c&We)O.7,RE1K/gB7H
B=F1\8D>-&ZI(/9?+YbADI#Ne&6cZE4-VI>&=D@dgM5B;B,g8P2N//DdZ][+=^HQ
[@6,Ha)8a0A#Wc9Z[bVJ@8Q=&0.XN6bC=cK8C=2=eLVDCa8_LL_Q&)WY-1bESGfN
&=M5D-Fbg)G)fBfUI5F1F[./P^LT&N^;#.[H7&8D?T27\P00Y4E[,e?Pg.D\0UD7
X+=RBB6&1E_\A^?3:3AX1EGO@)aJJ:GQLcCLKH3aBX<R21L>IZJ7_A_3a:.>7X;T
2<C?B<[#aI3ZdHBG8PZCcR^YZ.F2M(YC]ZS^I7&-BQAG.]4?55<)/4J=eYDaJ)dU
C;eV)0H.((DYKP=_CY#=GI<6=;2\^TKEU7@OMb<H@TCVMEL>cXD_WS)F4dg\A/R(
\-5Fe2?B#R)?J7#eE@\BRD1[cZd@_K#M#g.D;521<D?3P+e6_D/<;0J9E:9G<T4b
652K,=PR<0R^03dQVND108[:R\7#<2-NaD4OK^7b>TOR/)Sd-CO2)7RMULVfX.>6
.TMDd7QfV6R==d59(]fNAE8eRM/gL38:E/088O5;g4U7TaB&N8fQf<Fe8^2LKNcX
UcE6[B[O0&9-[W-LW02fTdg7J@B9@1OB<O0L?V_R,<GIef4/DQB/0c11HZ)SBE^B
S>O^UM8eE3,,]&O8-OQO-7)I[VQ_0^6e#[7^UQ/Y:=d1:T2>1_:]0KHJ\gM;J(UC
#>@,=\M-<6@294&PESG3<KR9CKSSD30>&W+Ue#_ZeM3YHI-gTeHXMLYOD/JTaL\;
+G?aW>9=8;5[S]8R8N:5S@QFPVEK7??R;5XdH/([J42WBTPJfR^0C?C;4aSeQR7N
2b[NL/@]4JR;G@gI<@EU_1fdXd98Fa#_-@I6>V+Y(?5VGK6\d-A-0Y@=R;,+[@WW
->;ON]G#MD7a@Tc)^,N_eJ?B0?SSE9c..JR2>;WVO>c<SJPR.<BCSD:3=\7X7=Ba
5,EU-3G,K-L5e>b0ZLB0bVBR-]E6_<I+WNES;[G==(<V?@[Lb@:QAV#aOe4WMfe(
>-ad7LCNQ--D?Sb\CI+?6U)L+Z/a\NUW:?RWX0)&WQgCbNWO=,0f081_H(Gf,T0-
-bW[MB5SY_P-SHH2ZM((c<+25OPCS-KER>JJ\<IJfF1=bMT=+Xcg,;]T-:BP_8-W
DW.41^PRUTO[7JWLKQHDdg6:.<0IDQ-RS?H_1W7d;H?>RU/J,TDM),3HM/+EcbeV
^3.@)SAJ_FQ:7WTPFN6][IW5I4PJU(TDaU7LU,R6]IR.\gH4f2Q\1J4/KTeD.OBa
c>:I-8NI[(V+7_\NE,S#(OcG]2N_,[1+;##9g8Jg#/3Lfa(/#\(5-<V@-3QH6b3g
agL/K@5&=06cIPJL820(N?bY6MXd)7;WX9^.#>5\VS;8::8X]2.JH+(QPBf(9XX)
ZL?USTE:b##bg\1JE,2DW&:F5OZJR490G@6&@-=A^M/G>CEOf7=-AaJ<IA#K1A0O
4SV#;2:,LbF5KJO),[_O=f[))I3F0>gaabVU.P84\W9792LZNBWWXKCKU,aF)\&(
&J+0+&KENH[\.D_7G[Re0]Ab\R/20FX,OQO9Y\\W:QFDM/GA[e<0ME.-efC.I@[e
[CDY;&&ca^W,D3H9[B>&V<c#D/LTNCN_<@B)aR(/U?:L)A<6D8;JA8Z:[aHJSU8e
N-VGE]ZCV)B@[.CAQXVR:g<V<Y4O\(,RQ80GF374FfaAJbZ7CD(7W&J9F_=W^3+9
YBD;2RL=NPH3aSB_=.9a)1c1aa)MO?-<88J)0BYA9G#Cg:BD-MM+F)B&WUBJ_CPY
B4WJe/\#aVM\OO#7MAWKXJUgYJ]D9[;OBPE.UfUeV@f<eEP@WS^e:9<LEQM(</+<
[cTKBWWFUZO3_,HUBI&CbL_2Kc3)EG_0=E2YPHbE1ZW=6@>+9\2a-M.LJT>8MC^H
YT?@IPMQKc1)eVRbHCP,f;.HMH5d_1WL?^@cRA-3B;.D#1D6.C,[\a&J^[B)59A)
dd0ebGPeYE#LZed;?\CF-2GcWH(a?Ob/@PIAP<IMW9YW4DZJ2TGWW9ZAId(FENRX
6SBPSaTY\\]7M-Z7.>LNfFW#<M-(Oc=bQ2IdU/BB..0A>d8TOaB6egJ_Pg>\ZHde
88g)J;a0c+?_VaX[:>8JW14d0T)SVI(2/B,@HUa:\:LHEZbTTP&#WcG4,S<B6PI:
@@1_C23H<JA70;&<6CMY?d\Y^)HLHL2f+</L.(^>4:^T7(I>F5\cQ0ETV)De5]f_
He9B1IgSMIT7]dGbBFW3Q_CTE\.]VEgS;5T-DGC(((dQL^@5:#<XY(GWc(f=d2U1
c-1:GYaX8UW6]-g_C(>5782G]>U2GPE7,5ce26dSJH@G8B29@BG-J[Ydd_0+>-e9
?IO#M/RD0C):./-a;ZgU;J4G/M7<[2[+WP4)9[6gZ8DCDOd.;RW^+eO>GGE92HOT
>Vd5>S28=GW2gd2AH#5FS#c&cTW#LJ=V0L/EI.Ic[Kf]N60))dE>O9SReVIE:\f-
+7H-5O=S)@I#U]1N=06F/CbOUTef&b(EB;UK@TQZ1/D8D:W9<-Zg&:UR@YKG;Y:f
0VX\/^:LY&=L\9[^=e3QHZbTP4-IBZSU(@R6_aWC@Id_#7.dK(VI.a0N>M-,JQ&<
4KQNRF83X9XKED.MR[@7f[.8AcaOE)\H9SG98R8@N0S3SY[0D7<aJV<9e3#Hf3P.
R:L;/=XZY[YAZS35674LI5,7CKIMfR[>8cDZeMM_QLKCW+WCKULM6KUc;8,f#+)2
PKP\dM>=XQd\RD;<;>c&QF)N=b[X7cTV/[^RP/#F<Z9U&b\W1.PBXcTf./>@R]=+
#?#5.T2cd+<b@>bD92R&>DKM0VcgYdeTAP]3,I>E&ZaS@d)G+LOf[I>U0f.3f2Pc
B0&6[^0gW6@WI8GbS]LEbX[MYGNT/_M5dTQg1<eU[b3=Q0.<fa#.TR^J)^J[I+.X
gD1+7(EG9>HDc)AX00_M4e:X?K5I\]^SEZAJ-ccGB_-7M^M^MHTLc6dJLCEE&+?A
>)P-2]VM+B+LLZN#MV>(dcJ^#dNO:#3BGT##0+FMEb=29@2#dXZ9>Ka)[UR&e1/I
&Y2K(0\d2VS5Dg0MA9R3,F=3IaQB->2Cg_F]&RLIaJ6CW=\,c?AaMLccLCCDJSY7
/Y##[/Q:RSD_cUHA<(L.X:IIC6X][[eQIeIYb2QI]\4HJSWN67).9d;L)[B6(NLM
=3?aN3#c@<0+eNS+Qc5<>@Z<X9]6@#SO\QH+]I6P2^U@9gWNPe6XW;bWKdMNQ)5_
:@)TR>dGeX27#N&M_4e\773FX+=+]eE-HU[(L0.UeE,Z:]]J@55bV<\C.f0bO=UE
>g&W497[f@EE#\IS@/9/(_JO[GOUY;-5F5P8RVZLCf7cddRaR+.XUb:d<:SP2_LH
&6fF4<,T)<RSRACN\8LK+8-[EG>HRagf<U?2,\RT\4]RESX5V=X:)GP27(?;GI@L
PEc^1I1MH+XEO6RKH0A7@Q)+JWXJ\NQ^S81&b5>]d+(KO0LE5LZ6GR3NIVVbVT?F
)6Gc)0abd\F[S7;>_#7)A@:GW:2W21;IU?W[H:K)bO]95/_C[1_HQZ-[06M6\U=L
7[<4cZ72C#KVZ82/#A>cI>RcOV/W:Y14+gQcZ11D&BNM6L>G)_P2GUE0A7:?U[eI
1F)LSdUHVDO;LOe6YWG2.?4K&Z>5^Q6&#L81B[E+K0T?@f>]RYL&8J&CQG8^bQOA
)#R?@KO\Y4?+=@ULOa]/I/R5?XIcG[RLC=ffAH@,(I.b<L#Ba0R)_ceP^=)d7>GF
(]?D+TT1L=^M)FH@L&+PQcB&fRFQ4VRV7WC:2]R>4SPP3THMddQdMO2P52W>V]M&
/]G1T2;e&D62LE4W+40f1GF4A<e]6Kb,=N@a7>=Eg41M^f;4J(e_GV8;;Ea0/F-0
/EB4L\SY5WWe5@aT/E-.>5#<b,JPLbQ5\(XG\=RQ7/;P,?]9f5KR0((3a/BYg,dK
7=WP@Df+>1=RW.E8+^Q77:IURHZ[a<+5=,L8@b4UfP6LNfWQ4U2dd:Z#2]Lg(;;W
4]3JS\KB<8=W=g?0Q[QD0?M7>L;?_e/A/;>JgGM#3FQ#a2Z[1<WJE3aA3;.:[OBZ
bg;3-[BP,>KJ\V3dNM2O.B=GQW6PP\&IU);J8d:2\d@3QgV0X506H=#U.)CQ--4a
N?eB_8dVSM(9_82@E@^,9+9Ab+U#,4K5fH7U_TS=g7Ie9.(Z1MVSF/c[AI[:TFI[
_)#4[8#0-A@Z[M((ATe38>cY\TQ3?QL?Vc(Y-LL3X,FG)(WaO6=OC(8I73>]L70^
eA96WXG,,W>M_KI,)&Uc[W5N;Jfb@TJ^+H.[B33+\FE[0H^?E#g)M6]gcNL6Q#,F
)K8>EfVNDA-\M>d;[d3M7Y>M@WVN-\\CSS2Y0Z>0S/fH(KH(80,R?QaY_/2R[e31
LV=6C[M.5KF@&E6aB<5fR>W3XS(7S9HZK:bBNdbHg0(>&#(Q6g9KTb+>?S,:#XG;
.dNHV.^?_a2<K6/EYK_Wa0,IMZ.BI;[C0OHB#_aFH1Xg-22=IDJDYELS7IM,bg3^
Q0(5DG+?Y=>^&]G(OCPQN,T.MG<GR<C>SN0MOQ8b#EK6TO/aG8#Y6]3&BVS?QBVe
?8K4bCD?K8<95=C6F_cM4#FQaR6#Pbf_+&TcD8NB<;dV\YF14_f+Y\gTWcW_+b>2
(WZ5/U7SNUZ_Nd[8A7^-,P5#b.F(T?>IU(?H6GI7aJXW:)c[J.Gb+?((FF9Yg(M>
-UM3_C4Rb?:g.Q>RQC;6:d/5CNEAA&cA6Og4:K,_cCX)(DX_L<?VY8J[\SELag9c
e83S26XY0],dDB.XFQ7<bF@abUG/4H26.:58]O,.#<]5LXT]<DY#@^a;6(D>Yg/3
R,=VJFKfS6<ZdYVB<b(EH@D1>_.R9+-:OLFafc5EV=Sa-9&8T4]6=E,Ta4g-+(93
@QCaS4F476.aGdEWUU<N(Fg)A=SO_/EUA^MHKK>\MEO[8<=d;&#<C3(8Sb;gT0Vd
S5+336,HU#_F8Ce&8eFJIXK_b(gIKG.L#c8A^2ab0NPX[aa8N?NE52Md^HFRV;8E
=/--MFf&5E6b0^ga>+T^O-#.dM641;=^G6?OQMYL95e&RR&2W]f+8]]4L2+9(3REV$
`endprotected

`protected
>eI7S2>c/(O:O,BeaTD0YHCF(H3Q]#d_RC6EQ(TbITfL[b,YUb[I/)d]d_O:Tf/U
WPWGbG^-G2/:.$
`endprotected

//vcs_lic_vip_protect
  `protected
b@N7]<I-;cW)]@bUB:MQ+^dA59K9-TE4LI<[I[:bFGc&283]EgUW2(-Ze_??0H5;
K,F^[R4Td+MO:d(D@=1E92Y+f=]^J\@5XIMT<;ZKZU7c4^4\0LI-P)3:<ZJ/1?_2
2M=84J^7bQ,DdQP]G2PWeSQ7-Ca0eTOMgb&[Z;6LWCL@UMEb9\?Qd(FL.\I&X<;M
aP6b).LSd#S0V?1EPUWSI/KE^O?)]4eYY-:@(/[e,cT,R+fDObF[0&C(9O,__#7E
MI7&#TZC[[2P_])\E_G0G<8=3V2UDVYdIUgc=EBa]9Z9PdfS4]RA1e/]RgKK-7d<
cAUQ(K=:RDG;Of>(g(MaJ0dS(^gU2KL/,.?04LH63bIK9/I5(O?1_@VBc(0YA]2W
L)G.:<[YCY8FKSF[)c>^87Na8Y\,?UAN]S\]]HHbV]YNe3<->>U)&.HF27Z=VS0e
AGIg1Y=eNIdb\)/6#dCMc8P00OFEGR&K_4Y@]@+[O\g6VDV#(D&E7>NQ5W;#?QW6
0GDWgRT3G@J+.5YaAI&X[a/.^5<,2]\)#-UW9_L/fdbg&INE3a=8Hg+4<J-_.dYV
)N9O2dS_fg>-4-_1RHDS1,YPA-39U<V7U)AQKe@JR+93LTfAUDF;W]<)3[QMgADN
fdMNZbgI8c=0C#DM04(&@]9-,4WYZT=G-<W(/?C))]EBO.-+@J65;bT_:EW_a7UM
)cc&^NPG_>K[g\5Ab[HTAS8g;Q9S41LUR2D=&:LJ+g#AHJ;/BF-\66\XAAMbd;:3
B5@K<gCg\@5V):<.XWQJffY1?\F]CX&I\WX.?/MCM7@]Z,?D6\6B^@L0<]/d7TC&
<T?5?Y]QT/7/\8.327FW5XH(A^CK^4QB08APD:>>8=[??B<gYA)6U354S(Z&,J3V
_(V11/NU/GCFZ-AOY0&.5LQf:V(D?.#+1d/3EUCK7>ef#7E7_:P&-D?Qc_d4#]A&
,YOLH?;G16CC;X<TbFOf+VA\9#aT>45)gNKR-#Q>:.<]4J>3W1Qe+aJTI4+d_K;L
_@-dL-+&gVggZBL[35L=@&Ig[U#[\^KXIX&PL>3P2NHaAP,;7[g9W@O1<7bO6VG_
0\SHWM3ZD;\<691?V#e3)RB>_fP@bE(3G8aE>9P#IE-X\50VE<9;6d2d[TMX@V25
A\gSL/&XF;bZc.YMG.<J,VL)\@e9?HeH_dJ^-;F#X]0NJec<&::+B/^L8EGF?^E]
KPKcPG_,CJHIB4W/X0793H001SfB>f)#A1L6(+:6(ZQPd;A4/#;@]VC]8NP5WFb_
)&SL0]5@@NRKWL?IJ./A_bM?SDaPIT+T(Q\/]HAU())K8H0:?eIF0>43&8OFV)&W
]T+UdJ5V7^6X\#eB8<<DF@[W5DJOdKV/0Y83W8WQ@@R5;CdV_YI^VG.#B.;+d[F=
U=S2f.NAD(GX.HSZ8C\]L74EK+4NUFdcKLRY5#?I[FIJJ4TWNILUgYX;X[1LaA8M
;@3:BQL+@R^(D4_<VcT.?f]XG\)VIeOQJf?dV^RVCG&@3^Vd+NBdL&[,CZd7g#EG
?]<40PG6c,fUNDgBZT4LaK8PRIZTSDXR2O(GOGe8#=PKdFL.;OO<?LW/U]2(c<)P
HM3IACCTM1#38[YDI<1.7>HefL@1+bTMf9\ME9W/R)?&,:E[[/b][O]Qe@bY^8..
J0ZOK>1#ZLO)AaV]\ONcQ6b^NW0-8V2]TU7ZN>Y3>g\@8Of_a>:-\O&Pd=YY0IH&
gX?)L?,;\9PK;0#8,ZP)>f_XdWJF7_T)@V+JE:6Y;@J;AJa<e4JYI,AIB:9DDYe1
)M9=;c7[;\0O+4-I[ccD:<#B>Y8>&CG6DF&8CeFI&0X(V)K:c(B2IJ0Yd->2JP&<
[bHX.Kf53\,N+])a<FP#bC+\65L\0;^0JP9TKABYXG]GEOG?&D,gVd[e0L4@(/gF
/g<V-W+f:5H2QX(A<37WSgUS/,Vf+g2#;G)789;).b#Rd?ReL7?,8ZYg@18aN9?,
_b^[c2U>,ZX&]&MNVG4dcKd?LIc,(MSZ]&OS1K6KQ89Y+[\K+1U>180IF+bA,Vdg
QY;7eH>=a80\.?4>OSJ<H;.Q1,P0e:NNWA3f<N,W@CCPO]&UKI=@fG[KSc)f:(0L
UF/^::?77QBR#+0UZBeIRcU]Q&NVA;^ZbdD=+F\>Zd8XB1\8JV_ec+,?KIdK2O.0
^dG?_U._>c8+PZf7LV6:H3_B2<c]:X)4([N=/4ANP9NU+_dVLKY^g8eV/[];RRZg
E@f_&\Q.>G90QASL<G\(K)Ad:+dAgH+Z+N5Z[Q1JJbSLREKeHd=YHNT-(Va0:HH9
-17GefUPSM#SOe3Q9Oa))AUc/bUFD2c6?[Q+:H?O.@aG1DJ0]>bFLI9[U88gfT+I
,MCc;ASe#QIN4O3/?MM?dQ\f0207G?GcB+gfe1K#9a,aIV<-R9.DTH-CZ(U\34,F
1,?4,aXHSI+JA;#L6MD208/QOLg87fA_R/M6(=[?;86I#g:4PZe(1.d=-<RLM./1
4R9;_)X\H0(E2I9P,>.>R;>-e9L+@&BV1fJ,IR-[=K3S4KC+Ue+dQ^0;4K:W8SBC
\GWFMXJaC3bW>eTTZ+_<<8M;c&ZYKR82<Hf=WX,3_M8XfRB^N.=&1(.b8R/]0EC#
HZabCG/8g2NQ=;>cN0Dc7cG;W[f;W)&H\^-MBFTfY&/cGZe?+4.YLcF;aI^.C1TX
0fbD4K,5eP>6F&fP5HSK82-&<Q(NGURK4;+b4LZOK)H&c^&I\A.D+K(a<Z>A1W@L
M5YZ.b>_fa.\5A=;35^a>0F^BOA0#;+57_]ZB]=3F>:[d79c_;a12;Yf2eHId+T_
CIeU>7Z@[NEH2MPM>1O+a]NVH)g=V-.9)dPaOK1)<<Z5XCU19\<C8GY0;Y^ec<E\
e/N&G)9-MQZ?\O3M;]GNg/7XE)VUY:YN+c,XG@NbB:UP)]<)@67:a,#JGSVPFDMP
\<E68X(#>b[^E,Y/Jf1gM==+[F2,LX@3]JZ15N6B:H;DO[[DafFbf12]Z\=L.60Z
8/#]JRJbV2QcYa=YSEE(g3CNOUSde=]L=bS2ZE4T_2/RZSBU@KMKVP2]K$
`endprotected


`protected
LTLSfA>d@>LMb.D^e(bMQH8?fGB,4@K2=2BIOIaU,[aBAD?@I6Mg+);=G<:8WaZH
cZAOCO@FHHMM.$
`endprotected

//vcs_lic_vip_protect
  `protected
NfSKcLGZ]bZ_ee:X9R.IX[UBC-NN?f,#A;@3TJ8fN&L:8=[A3&)61(6d,g#).HSU
@47.05I)<S)EA[)]#0O>;^F@c57#=]d2^)8AK#EfI^&\/:8V@1N9=-f>C2/A\K:I
UdTY+B>8DZM.]\6]N[ZSE/H,TL@/O.O+1\FeT_=V_\6?8C?cL64].E<UZ86T>Kf@
KA_b&(V<QE0[S>:,/)#HBL8[GZT^FbPD-2e\LD_d+1FFK+<KE3/2N7C&7PT^C@)f
E9A^d\:/.U_H\II/Z]Yg263KW2UO=]Uf^B((>a1W]/#a>Wf4(PNW>#W7MOC_WD.3
1eB3/OI^?P;Z:T\4f,:TM@:PXW5#JP+,]ZPge0D/1O9O=\XMKPMN:b.Xg3BCD5Z7
cEB_444DEObCX)9c#]A+d]VUYG5EffbWW1eSQ[0UDL_M505O/&L,Tc/1L]7@Bf>f
<SBQ&3\=-?^[1=d6@=LG5)A^W8:ZAdaLM8@FGe@6A)JJWX,2>40d73H)6@:4g49f
Kd_^3G_CPM7?b<[D^2)@,IK+W;TG\62>R&1[YVD70.;c1GIU5KN2QR#BE\CR)\[E
aJYP.;fB8)EUAY():IPRZ]Q-GG)ACH;R2+-fD2PC-9Kg.]@UceP5NXH#0XB:Z<5B
]:aM56d4,[?-B<Xf.NcZ/8O5YJS:f)M)Q68c#DNGI<C_dG)(18W3DT2NA6OKLcXC
A7Oad-,Y\dfD/NJ1FYM_Q_2RAegZ#<BAa9A@D>4\9[_L0BP.?c+<PXC)e:RYH4g,
-O8cgg2O&;cN5@US^NU^eeU9+;NR(8V.U(f4SK6>VKOE5E@f>e-+2JG);HCe]Q>Y
GYI6_CG7<V+_fI)T&KaD7#L>:2#V?&@[BC6;ZZO9^O2gPX-b&DWC=)I(@CMSdgg9
VNY6G&>E20;^_1@RH3e<]3+e3X:F>g0?[/g)IENXCJ\UVA2G0]TYIXC54H-U@(64
Ze<R<e\(>KE8K/CS)E5b0^&<=:.VHLV,L6?7U;:E3f+S/B>^E-30&@C^2OL8J_c=
K4:/86?0RZ7:QOUXe([2DG(d0XI4g=OccUd6?JT9aK(:&d;ZbT9OOZ^MT]://4>K
WRV.8[KN))8Ecdb_d[R.36)\?CHgce9fb#&?.R<)]g-;Z4B.3XcZDYb6&KJRD&[4
E8Ke(T\OR-b^IC&=1ePEQJAE3OG>8\]>//RSIO-13.DE[)b36A3_+=f^?I[O@MR2
T4TG+g8>f4[J1-[1;VMO#bW-LGHTH<)cBd](M\Z+71e@(7ME:_>DI;[cTKY35M_f
?ZC4Ke87&EgB<8JAE8;TQ#Z^XC+;U41#80A=K2/W^IA(#\-dag[;+6JT4S(RGQc3
YPW+:OJ+<&L(#,Og&^g7=GCP;8Oe+eF^W(.Fd]FX/bd5=?^e-N0F@KgFPCK.8(9d
=94FV/>MNe1#0SCMfL^YWW8P=0E7;5EYE.98WSg\PfMLHY<\_ZVW6e1.UX:M4V_T
=(H<NSWQ=3G;^I=gggR97>>/bRAAWMAD;;3;_&??9[&+=<ZQ3A^\1<-ND9ee,<[S
2,(JM7\K=[HWAbDMD/OD&bXb=KP24#H-SJYG/_;CS3J;b\LV#gZRLA5D1VdgbZ]f
E[<<7ON7P18YI)6A.daL/O_2BS#;0egW7IR2/[,UbJCMf#TB77)4W6XSb8H?>eBe
XCWVYG?6&9A(M?Jb0(K9eZ-LO.HP)ME6K]=a;E\.&EU/JNNeS6N(38GPH4Z8e42f
<NQ0DU46;;K+K^CG4.]H=MdO3Sa;eYS?R3:Y1Dc&4-0aSEG>90?Z?FJa7J^F,5TY
3<6.]C8G64HC4e->13g:1DF<D+GZZW8QS8UY;E54V+Ma-1ZW>]D_GdaU;;LOX\<5
3dN=5ND]-8bVbdcET4OA#e)E,:+([=HM]AMM-2B6aNUW;dBMJ[6./-fU._BX]8VU
WEM^MY&,K_U3OO-0ERC2gWO@9[&QL<6_,#1\7?e(\:O5V7G?W65(3&-2<b:JX1<R
(+K9f/3fbOQd3EL),G/+CF/25,X^]7gAcGN,F(,d5+A+:2=T54-B9L=VFCcH-C;g
B<_6N]AJP<MAX--]f>[>TB4a[(\O+Rf\JHf>;5VT#AAJ(Uf,F1+5]>eTAG<5A#O4
[ga1M.KbI,L.G/4)@>=1>)T,g:7#Y2JZV4FPUC&Z,:)I30dPXd,A<T+]]WK0=Z^;
(FNHgE()5eM&2YA3RfgF5)Y0T)9^D_=1W/c7>I,gK&AH-#IG6<F_X;#[;]R9-QWP
(/,<&Z[;4W>I:cO]bWAK\e@5J:-R3g\16LD/JTMBD)eY>SSLBP+T)N8N8(0bM&,H
>aTSU8(7:cE#81H>MG]0SB3NW6[Ue401P+9]6A98]YUR4AB6U.>GM2XXG8^UNKaX
4Z([/A]DA0.RRcTbCc7dCa/GW0BT4:EdV_?#]V46d-3TS+VUae@OT,YEEB=f@SLK
&DF8C8<DC6,]8H[7.6>3,GLOB,Z/>_P(Q:A@I>2d(&,>JIaJNCcX,N0^T0SfDHF;
1&6bb^2]@]YX,=O8HE,K<^[CD>WR3f)V09eWX-\#WSOeR^fT5_^X836/GEVLD[7<
-DWe20ITIFF-[9C8:R154M4Wc0_93O&#G]c3RTY=F_@(4J1-\>A/LM(/(WA(8KM4
5<8A-TQ\/gFL49f&VA5<T07)C0\<44YI/XG;18V\:J/Mc,EeTLXZLHa:dbbN(6WH
L/><((1aC@:MR>Qfb<3QC^8A/?0>:W^E#L9gbI/N>d8>#C\:-<7WK&_^G/(RD04>
Gc0QVXB/7MN46gX[g:Kg&cK0P?Fe^HO:Q/<R25NBQBAM/DXGX,1G8WBg=L.#d<Yc
88/W=-Z18M/.#J1I<KD=^daZ-LEC43ba5[J:M_6I229c^@>eNJ&2;PA(NP;?56&f
C@b#O<[Q[aPKCN;CD;&P@CHFITYd-c#=G6^DNZAFdC@CY8Qd<+040c?&.()7?[4>
/^g[EKEb_Y/_D#P&/U3>))bWL^TNDB:?NCg@PBGG)A;3AQ)Q,7C0NY<f_FHf&L3.
I\f#4;X;V,5K):N5F\CJK\L6@e,/.,MYP1+^0ZcSC);325aJ_>MQB)J?EEHd@K\(
Q=C,)Pa[1PTLU3EN;Q7_.OIK@egbS()S2T16N9(M(+2VCD,FTMKJc#0.)5JC#AC4
?.Z[cc(56XdS[+6;K-P0H0FOf;W9D;CY6J.T39&HSJK?Z7Z\3ZMY8/IH5>/;(3aM
ScH8L8T?eU\aQXP28421a@2B0SI2:@\4#g/,)LFDS,#OCRI6JMAF:cQ32eIdVG;:
S?0(<BZ93PZJ4=f:S>f//cW<6P;]YH&?U<^0/F2)b0@^#>a7@ab-66B-9W)B/=45
#50+(J,Q7AR[.VLV/#[e#JK//K=eMCR3J:b2>OMBR;]4^V.>c7?[IIG2A83K:f2/
8#F)))aGS.dY@g7I+Wf>D-?VVR>+c&A==$
`endprotected

`protected
M:E84D-K0)LUCJIeIHLE/WG7)N#IY7/Vg2-Ng3L9g_7,MNY8@(5\+)^4M1=WcM+5
[[^5;bLVR>[1R\FD,P,Y_)G78$
`endprotected

//vcs_lic_vip_protect
  `protected
I^g/)-KcIJb9@R3^Sb+:,a56CMTI28a>_C+S;3QV1AB,e)g>]b#X7(G@)VAC\g:P
RH?ga.XB#-?7D&+/>JJbEE1CUe/>)3-ADO:B>V##B7-S\PR]?_[Ue&).)<039gHa
&52e8f,_g.W@fFLMLc5S9HZ-dI:9#Y]O&dH:5QKcc)2\If_3Q;6H;DS9W?5G8S9?
=G\1a?\fFR0K.SE;_)]Aa3/ac+bE2A3.(0D>4,?[1Bg7Z_NU9\5/GCb:aAELXBA\
J(8WL[cRJAY/#2E23X2;B=I_;0W^J;]YI?@7IW,)4c,]^#9##@\&40gZBQ?;V7X#
)bH&X.IDJ7]<#N/D[e?L)UN3D>e[^ff=#_](6:M;YSS\MVC]O@MJ9RVV#O9\_[A=
-XV:PP>a0/D+)fD.H0O8K5#Y^aT6Y_-N4A6Y:K:\BD400A]Z(1MHO&/>e9YM@_K<
X0?)e8\(D1)V@GXY:045367f6KRU6AZUF1.\-R.>F.ZND-&_e^_=L;VZSLN)(^Td
3VJK>GLSV&M9VJ/;LT.XGY8[W+FeDagG0ga]T/Y:=;7Fb,8,I-=J.d_L;UAPQ2AD
ggT12EA]g)5P=]b0L@e/-2<IeA\-]W-#\_@c^1^4(3WfFIIa&[AC^Wc41Ra>?W)P
g1QGH-RALf8@W8;,:e4IR+5VT?P9GJO8#>[&IB1XJZK7@&&(MM-_/dfMda^B[,&F
ME+X/]2Yg(+?H6EgIDY2-KQJ5,aKY(E4aPK2I1@f:dHeWR?<_AZf9S1=edRAd^aD
eAD=6;c55?f5H4E62-fV\gENDQ?0eAW5\gfV83&U\eYJ2M+RNS^K&D2d?:/,PLCf
>J#/U.7&]b44-\?H:/cKI[.Z8L)5Yb/E_gULAgTBHIfU76\K1_T/YX,7W=H(3^_1
cb,XX^dEH?Nb9aHc<D,H6S7I7[WD3W<KD1OH^bHHA[KNI6W]7JPG.&&DJ-ML_Id)
SRG#A=KE2[0391O#def4b8CEd?>,0W\[O@<E8QF@Yb,aI/5/Z]_S(I]IdO,M,G8X
C]KXLd,RN@aLcB^ONQO\P6=UR7.YY)I>OR9aKV_R)6BLge2_]f+db:(eF)P2>ULS
B\Z9D>THYE->6eEVN\D0/?OEbN)X6gb;:3;^17-Q]K(FXV\JOLVTc^>9TK1T+b35
^&8bS(;?3Cb;/8KHHUNb0a</L=V^P-R)F/a>>?L0cCfOP7+9a-B,7E1V@922ED)C
2@8=Y7f8#U;0TbCW4;aKg9:+CR?=d\;MWK&M#f(6NBQ3G<H5GKFBXC.+Od&;@?\7
RecF9=M8>Z/H\_)EbV[dD\&dZQW+K1]Qf(>,?cQfH[G+4)#3P7M^eV(d5<^A4,]f
=P;([D4)Z5AITSA1S[:I/C>P1\K8bT5^TQ08(12F_c&,E6_^Ea\H4DV#<BRJ\L@e
8;=.44CI.__/89&]ZR]&T)\K&F(]DgdM;YXFP;KW]XM3GJC/:4#7?\ZX\=8=+7<O
a[1N,QL6BMBKBe_IfL/BAf#@CY]U>:J943=geeNYR9FNXfSR)_R.bd<(2B/LN9,Y
7\FdVZK9B\NDOA7(-L;5Wa0XAM/N5@9H-YZ[CEYP4]O.7:3;^A,.@W?^K&d_.?UJ
gF(8=,9C^K/Z33LZF?.5I^LO25FfR66H5VDAS?DY0g_)1d=X?(<M=A)+)KXL\OHR
ZM3VA>,F/QSZ-)b>H,,/bM>:cgJ97Z6a+>&Ebe8fKB=86ZI\GH];c77?GL\8>g-?
382PQ?\c+QA9O>4,]LeZU\)C3A4Kb1^edNC^MeH_7>T36CZ_C9Rf\+.V@?J7Dc])
QN[20KHB:4(DMg2BI-.Ie7,RdZ<cB;c-X2>RK,8OWA5?_@8HJMV(&BS_6/LM7C7L
_gYAB.ETS^\84TJ8,>?;#RX5C:^H9ICD4H^&YOAQ.-9-aQ[D:=3RHZ:C&;;eZ(Z;
<A^8f9g8+;C0G/Eb[gKS2WMJ^0?4M[I6.U>SOfG^+5G1)J2RV)R33B\2WZ:W)X/b
_3<A7\]#<0>C[Z;6N[:KSYEEZfB+0L+8O[H.IE]JdWO0RT/=9TOPORb4]^I<b.\<
<P#..3QdB-\R]-X.d1RU(0[0^R9K\0ZGW_-U5KTIeU<W&Ma#XA2GRfQ>RTN16#KN
J&aA4KeLR&BGCa4G\gO\9&+#^_^[3/KO\)4Sa]1?=JRL:0Z\/XI.T=MUKeYdc5df
_62V#U&IT2>AE5UZ2DK-X&3TbH2X_56MFdF7-5@#5g537eB7^/5_=d5-Og,XU_V#
+@IS]5WBFI3:fA5fd(E5(&5(A#261XaPR;S3M3bYHE<ZQA3R.-]deO9ff?/g2T.P
\&YeK)IECb..,6VB9_[5CCJBJ6=/Cg&OZ#_]3YdDU1GE+;+SQ+2?J7_]-[;8C?,5
:fQI</#(6TPGYS,U;LVD0\T07K-Nc<THTD;U](-J6@E[c<17ZFeGK<Ff)JI[6OA,
fAg,c4[DLKb6):9cC0POCCGQ<&^?727ZbXEW#c.#8>AM\93QW.>T9:EQe)])f.<I
/F^WG4&)Ma[=73A[;5.d>]9>.U@c5RHKOC\^RW2M;K&JEFUOH,0<\G5._26Y4N_)
S_(TFN\ANGVVOYT4MU\K;5^)Dg/f8/-;]J)V]Z4F-])+c[:=ZT6E;dd<]FZ\Yaab
:OAb1APO8,N/;(MC[LN=.CQd6=CI_)S(a@dK050W;fXfdN.=Y]MLc.0U2^_IeB8]
&W_YY[Zc+S7@S]d\Xe5^5e&7PP.^(bP&RW<&_KOb+QfUHET+Bc3YL@HE-2FWX^JI
)c94XeP/TVVM,^&;b-d8M7C3g=f9::2TI>&(T-RBS<(NE[2VC?6NYFI6L7)a&IA0
#O8257OQ&H/3N&@Wg=[Hb:=f]O:[F,H@A^MQYgea&VH63#:X^/9UCD7AJ+Y>,N2X
FLY#B,S]U&cHH]<?)#6N<Kd84.S-Mab[0Tg&gUW-;9]CBR/P/?9#1WO?]f>P=K5M
a4WHKQQ.K;.Q+1\8d=_5<d.O\[VN0,7/8WWM&BU[THS>\[\4f^^SdLd>]TK<g&8Z
\/:)B?,fVa#NIKN,bJMDE,]Q6(bVQYOeJ3N1^@T/L#Nf1G+a\9EAC041^^YR)ZQW
=REV5fZ,&7EE(b^Qg].7J^Qd02]=&L@ggf3__H_d-X.#a^5P43GN1#daI@A=GHaS
Pe008_)HD9W@,I]7Q2aFF[AW^V[;QdEDL+7K>O3UbCUAHR=0;H\5d]U=?SM9d1Wc
H+6<?9B7HO_?A]98LT5;f9(K.&^6[98#[4LUY:4?60@a2389@<Q:0LN#?R27H+QT
75fG]d56e/GFO30[Z9ea+A9ccUF9LP+L.>[\M9[G>N&IP57,+0_28Y9G.[CMUW7+
ObFCOH#J/IEBZWcN>E?L1D5gL=O,P@b1(N-QG7E):X;C:D=b)+<SOOJ7CM+N[Z<0
P:7?I3PGY(<0NTSO=2aI1A[Yg>DDZEHg#\^gHfBKN]Y^VSUHG8(OMd9fD3@:aU^R
M>MU\5J&AO;NC<4_NE9+bOHO^cCP5?2V/B0)87eY-4G0KM@>RP.6?]?Q[G5J;_-=
_]aKME^W+T7UAO+-FPXf2KO,U&3AI>+3D)aWE&(fHaSP]SeI6F<KB9M_>G.QJGJ3
&#8IVX)FGZ=Sc)Vb3IO@e_<_Oc6=C&BDSUa2K1R/M@HXUK]M5;Vb?e&PN5DO+8dN
0PM92SfA)+R/_#X2Qg.68X1T1;Ef,D69(,P_4fYA-:MOE9Y_A\LY0GJX\Z<O+_3e
#Zgd/C;YfVMZD_64e](GQ33^Rf<f/.C.W^(Q9CYB;;K]W]Eb?;JD+\/7G5,,QVgT
Jgd4M&&JG9QMLJX&cDKO?MO6^Ib\G3R-a1R2Y3.e@3(@27^;2gHb<N4-TR)1LXaF
(Z=W7]IX=7.#35<D.N=gRHTNG#^V).d+UFM]RX,XcS7a7C3=:#C/[]D)F)H7gSA1
ACFg7d6S/@EXW7(;;[F=@T>B:2deP=;8=)eT?_#L_b-]10H83S^NaI0G)FPBY+Ie
(KcIO68VIb<M-eI5M.cC@g&(.Q983P-)I0T=MJ540XI_fNaQUB;3W2LgQJ5]Gb#@
gF@aT7O5<YMaL<M([N3YPY,cPPZ-2#PY^(51B+^2+,N8&SV-TTC?adbcgE)A8\2<
@,JK,>H@(eJ??-#NeV\>WG&FIS[fXYfN=>-R+d9<5PI9&EDSR^Q6eKSeZQ..9<VK
AYN]\(D<Z<DULg)&S?J@dMDCENg5OLI2aPT?g&_[0V@->47V5K/C(XZQc1XY7_c=
<1dHRfLL@HI:L3]g?JeWVR20(>_44QD046514LH-.LbJ>7Y#OS<>Yc2H3E:GLZI3
&\Q4B2P9H[\@3f3PXf]D-L+9;-e-+b77>a/TICCXa.H5V6#^X[FMW?,&8X8&#?OW
:+CV+TDQL?aU;_dODdIK?7,(49J.fPH_R79e9X/VX8V.Ra.PDLI-H4U=+-RM.@5H
05\;K(T[?[cI?O55eARgK3@.[5G/W@@HH0CPQ,MGGQ=UUCFUBW5QE&/aAfK1#(RB
C:/W,GV/cf;E;D,33S7N6a4WFN(N.\.8./O=<=DN0K#AaJ9.5.)Q.X[K^48C_A+;
JTfV.=;/=,C)YK)1VN;2fJE]U02YQ_\YRR7^??F&3@UR/63QK#[PZ5,8J-B0QG[e
NbK0)+H+-\0C[CN0YH8VAZPR>/G26412MA>;[P):4KIR)J@4K(C.e)W6^8f=e:BI
).BT5e38]A>4^_N\:><IUfXcTDEb@R-FL94U&.:=7G.#.:/9H+0\V#XS@X;DU5[&
A/<P^V&?+a+_/(6?g3+RLA/#a?7Zabb-5]R\CW]+3=<Q(d3VI@[/c11&>DK<6L\<
:[c&1++/1I,-T4M=OIG_X=R_Y]A7Xe^X\JeQ^<]9Z[g-+]\;-X)K6f2S&?4Q5&9H
:49QcPX];=G:)9</7^)MdRd#/XY9SMMfJ<64b66D,]1)HSNcT7SB[AbQLCDWMK&U
GQY]8b]323(J<RME#UbY^5_W[?NALJ]S.2_>b/4G(T^fdg(JaY:3:41X+L0.XO3M
T.\=ORNUW44-KW)eG\KCf6F6G[_),X=?2RUb&4O5?S\TG=AcMV8O<12)9>]Qd@59
eMCQ.(VK;MfXU&R@Ne=gfPTAN[ADO4bX7I<1YII2HYM#b&HX2b0N5HB1Y?;2-]E)
.HWR\3YK=@9dMW#(7WBOA1gRNS8>:+CL;#aYQ[5fWYP:&9N^O8@dJaJ5J.CVF]_6
1]11RN(5D/?AQ6TZg;,bgQ(RU06P+W[\b03<1Y;&[f?Y6],D.88Y=F_2((IPTV[?
H&\>[382#\RS)2C.U>?K=_<C6N-(]6H5a;g5^@OBV@=GbQ-I;_gL_8[L\K@+V(5b
2?4Sa96I+R#/U/AgK-=D4\Eg4g+Ff3</FG0@HTb7C5__]@XPW,4P&+<GVJ@a/)9K
__(#)ScBW#<e3]P56@beYAT3MCXUU#\15M?M=g+M0^O<K_2a;RW)[?4V(f0bQ8,_
CbCCdW3&a5<W0b0.RPQCd;;S5bc>GcOaH?_f@B\bgR5S3/19@<JC[>=PH9M.OA\T
]gARc,@U4M-McS[CTCO2/\WadN&9>95eCOAA,BG.PBd,K=[[aJ[Pc?3W>3P6QQL3
B1YS:b<O2^;.;\\#R&]VKbbQJ?EWEEJX&8BC>A2b5>1LYXL8Ha_EC>NBW2Pa<UF?
a0R6SQF[F[?OBN-:\&&T+V@4^bH;d[/K818d_@T(VB=Z^8<#QC=_&.gLagaQfW/X
g]O<E4;,1d[PEddKY9K9/UT8d)88EZ;c+KJ6E2ee2eX.GD,eQ#3KC]0)+bCV.&KR
9b>I1PI>:9C&L+3@15EeHS.S]-@P1CTTD4@PSUZ.H_M:7GSFF6B1f.-[A7@?+F?P
,#Kf+-1X45K;AFPU+51VZ](YI^#BV.,:662@IdT?)\:2\N;)N[8c)P)8#H+^?:C1
V)IUKHLD^D77>dK9H>PeU^U2J&):g>IfafJH]/V475=I#2\M64#P](/GE]_AR3Xf
#Z5gg,c]E4e&S-(L]([6OYdFV8,@WNf2AD1RIBg&E/:87Kc\U6S(ZCS=##3c,b\H
./d#Y#P>^14IaDP7.(Y.e47VQ.Z#<KRB^Y-&@d/5&bHa#(_.V9I?EKC7ZC-aX<Y8
bDfe)d<Eb8[NFE:aK)MX&?5:^#QA@;AUcV.#5,d\<efCM1)OgaGY_JeS0gWKL)b6
_7;^\V/+&WEUUYWIP[QB5Q@)K\5YZ:TQ48A-UCY5K<NXO?#9PR]Kd#bFV_Z8H?U&
_Y1/_,3C(?>S>;RM9VV6[M;-a7BOZXM6BbJdD>7^#+=J\H8DgO4B3@_a/52FV_4X
VcYE[IDB7YXT<Ng4>#K-H7B0HLa=Z>P/>Y;Q,7^Y.K.Cgc+g?g3fWeXEOdF8L0#>
MTU?CbN]Jf[FCd<PX95ID6cNP<b])/8;Ld]^-7cT^\IN7fB90JO=>PNJRLU8E&Wf
S?;<-=Mc/B0GBDgLYY^@^GA1(@]@R)Z\/]B2X9FJ]BA<SB^>H1g4,4]2d;(IG-HG
;RC4Z^W?dF[?48e.LO:HBcX[TfY7UKDM,S59;AY03fa7Og/5,G;IWOYTRF+U@bAG
^.f:K&J+:E>JA&c-#Y\(a)IMY4W25]<(T_La:f=,8]2]d3WN9b+30NaYX:C9I\,6
S\YDF]E1D-O,46Hbe@WfEK#Z<DZ@bNPX7OJK_Lc;]G2ZbP58LM0:JV@NG?EC/4<+
D[84&]0?ET:S1f2<cE7:LTFV8TSS2b.>/g#/OMVb=<CMLf7U7ZKecE)INEf.:#W0
&)d(K64fP:(4bbRZJ,IE5_&F,LQE_2;(-=,1ONB^Id3)4@[[>7>1ZWfaYP9LHZ(U
1T(aK040T2[[f@6/g6baf=HgQ;I3A_[VDWPcM#?@Hb\>K0\&e5_20_C+7R?,07<P
HLdX)?UT)<AVT#[X5Qd.O4N6[B@1]R2T9N,/HL6EMVMSI5gIQgE+M<(/->TZfYIe
(A/c8Q<N:;gHfZ.E7C6QRGW^B:->NERRL>;V./VW-?61/FVgOBa#NQ\AK2=7@3Y5
6a6)/f(dECg_b4HVDZMFAWND4M^aaND78&bENI=@Y45&2_-7;G9Q^Zd^6_JB[^c/
+&d]^bce>7NfK[fZ)V4()12[Bb1)RbA?4S-/:O;;JeIQQR\8Y;(PQgY2QWI7dcV+
LM?^KH0b[](C:c5IYST?6@@@B8ZV:>G>7=dHb#9U[\STZH_@IY4=&-ON?W5G;Sf,
9A\#]GEeK9_fMR-7]RbN#+N,WV0YC/ZN\cD5B1c2,S;5\?JH87d8B(4@HBD+&\;R
P]-V5c^;6cJ=<N=:Ib:#:MVY.>2g7YIe1=XFC;R5^\2/?P31RR@aK;L,f59>cL-M
UB=0_Z.5<H6SaFfCUdC5gS/L82WC>AU+1I\W=^7^<Yd<+[,MT.#YKEFADESa7GP8
,;8+O9&1OKI&J3JNIS:cBVX+#\JC)a]ZFH;+dX0&V\H,DM&5LX=P=HFgFFB0,W[)
M3EY?,[7gT8CKMP14&>]3N92O],D2gMF_[C2@^fLB^T]X[++U:>COTF@g)CF&QU:
4YU:O<E#:&VYE]]T.(ULNLI]d_>E7]_^/_+8Ta+a_KX-(KWP9d5WP)00Og]E@CC&
LCGb(gT7R(M]<?(@7A.O^GRSZ\8W,e5E7YZ5Q<7=D-03:0aS_g,\MFda,3J;gQFQ
Pg&\M?[cB1;A3FeI.<AYc36PACFPKXeUaBYG_(.YI]NIR1d#Q]&VL89\/:QW?LA/
I>:#@;3bE?.#F7ED.J:a=[TK/S;,E(XA_c9b89<M-F&Rc[eI^N(1c)4L/WaQA]&X
)M=8H=]V\XNS?Y26&K/PTO_/=cOU7ad<WY7;1XW+M-+RB$
`endprotected

`protected
]_)XT-PVANI7gWT^cE,:;[J-\f1d>4&C.LW[deV.7Nc4,ZC7D.2L4)E9X0c=RBU]
f21ZYJJK1DMP#/B/(UHD[]J-4$
`endprotected

//vcs_lic_vip_protect
  `protected
3@TR7DR:@:[W8Q@EBVeA(R]++UaYA:36^I;1^^U]LSSNF#cCe6A\&(/15[[.A4Ec
.cVQ^_)/G>)<e-B+:EBAO1:_^BDG82E_\HC[>:bcZ/I8e&[2H\0/FabSAUUZbT>>
CS6TBV^PWFM)O4AIPAC#8Jb:<X]:e?@GOb#UEF_)\@YJX-F:NGW2b)+dS_>YeMHX
N(E-,27fK6^VGc2gW^G+]&_NTJC;21N[J4+O7a4>/:2-E)H(-0+gNK.dNa036:ZN
@b^KCGC7QXXTaX?WVZbP@VS?12HVa1E00\d\76L.A\,3PQKXE^7--37].[PVI_0b
Lc7IeLg9E9eU6W29M-ee?#H=f>)A7YRRC7g27R]5b<^^+G=V;RRLS08XVMedJ8L&
&SOgg_SV6#)J9I.^a#U2N>WQ8&\<O6Y37Y(_-7.SeXd/,dDfFg8O?O@XHa]C-NII
WO3;.d7g>T<=,K6<X<\+4?1^)182Oa=CG7c3F=aIZ7b@N.?,8I4;4^)#P=1dA;9H
.]KN@_K[DR)/)J2I&RP8Y\0JWTSY]ZJ?f5N8:faS7/6)[J2YN9R[S^=F@+J-&/MJ
E^@L4CN9c[3\>,a+Z4,O-;3GV-U1bMU5:W.K;BQ^\=U6S<N8\77Y;A(dUC7W6A0\
1+S<XX^V;+@af/6ADN9FCCaKEMSXgRKQTXT(6>?]X]ZAV2\^PQ3Q^K&I6R][84D/
Z+S;EH9e3GJ3-_VdP?9.(dN^C??-G?:\3e>]C0fge;6(\<O>,8?Ub75AW&8:TaVO
Z>NH5TIa-E)Ke25)BHDU3A\Y;d/+PB;4#CcE747E7]E8E8?Z.a1+D0#c;AY^Cfe4
P)UZ-?e_==cG0VYB&Ef<^90Pf@RG<3FbFM^.;)NRASEF3+>aH_@T+N<I^B7[T.bb
:LUB(3Tg^#:aFXKHM/3A3fF?U=\65&GBPGZ3/5@39+=U#)fXCbOTUFNgFa>R_gJS
gMCNZMPZO/X,Ie00-=Nde@L3GSEI1PYRZCTL,9g@&N6Y984JbY+IeZ(E=D@#0SJO
cQ#(9.CV_-dN>ZOEM?WCg?77Yb^_.HO&^^3-/D=4S8KJ,>KRZ)BL-1.14+B@@+Nd
3E.\GFFC_-11;Y+>B(MO3>@KO2LI.B7d<N-gJGgXP<<800aaU2H:4edYI&#_<C02
OUF,,7#/6/a+^cH\1N[Z+GII^AC0a5-@G9E?Q#>666a]16FANA>M80#>HDMH^0/D
D0KYJQ\DV]XBeVBE@WJd?<Y@&#]0?-Ec:H(Sa5].fXX\f26V-S]&_:7W0fZTF7/M
6D;H7C^JA],[<)A/gHb.3.Ag>S5YBIcL1MNL;GH[SJKD&YI?FT.gAOQBAH(/7O#K
cT7&4,3\#(YeZD^B]U<H+5#Z_d8XV=5]G7[#:,TS//Uc6Y<;0T;_;47PZ0#L];:L
WD/0>U.GCB>54G,R3TO6?O?:gUU/ZUCP&[)3Tc0)[#JUF[Z+]\#ESS3S;X=X@.KG
96/<-F+CJ[2(TNRT,65/GT7b:U&QDD)/W0LF[K_aD2aaMD>/GgcU31N#(G#7aH-&
P>cBR8V7X:+4,T=Tf\-O)7Q<61.<3F+2AVT/MA:40-;,TIa@\B_YT[W+2@<8c?I0
AAf)B;SXB_;;&]eHWd\&YSFB/K+.ONN^SWIb+JBUX/bNEI\?Q21G<P:>-^Tg\-Gb
#.b34e[\0\_K)R8aBR9Qf,Gg,?5Tag[];@e9eTHY,&O#UP54>[f+:H?B#LLbO95e
;NDT)]e[ULJCHa]&F=^YHAD/C42@3_TW?WS7T?EQA5#PffZLBICPU3^3Nc^VAY9G
5EKHO:VJB3ZS9V-&CV8O.J\R#OcLE,1NV[N/HBMIbVZ(dHdZP-3#JE=(b)>+eFQH
Y/T6]D/)UO.V#G6]ESS,JH[\RfW]-3&JYFF[E+fPGY,/b0KCb\3&RRMe9^<,A<5^
cX0BN3_>NefV_.H?A(O5\U;IM_;K^&E)H2_8def+5V^d#B_=4-[L4YG^c=U@5fC5
6K.UIM(HR4\)&N:&6^eaZ>&6#XFERWK#\,RcG,WaFH<4c@Ve1FR7O&3:G>AKJbPf
)6Z^4V987=V?@.([YU=eDgGfL(gcZHGPETe@Je/aeDU=AV5+G2Y&MQ/66G.SRY@f
g@2^G#NM8eH9Ug,6^eE<ZK[fRP[;RXO0&/U8]Q^c6LVO,IIMQeD2#H)4ZJ[+-.&0
:XQP33=#>P8WZ\J27Z(Ja,)fLW8>AU+/g?=&X.^]_9OP.7Xg[e0YU[_OJ#L^_)-Z
S3-Y;Zc.>K99D1F6[+D,]9U4CC0N4Z?V\2CM=G\L@X)LOSCd[[^dF+5GC)EP8PF)
_[[E15B_MZ_,5_Z>(Weg;M0O@QB8<JXPB+\&WZKKZTe2#L0#fC.83bLXXe=5cb8<
-U9^\6LPH,M<BDBK,V+[<1b#b_=a-F;=&a?<H1+>V+R_SZP+aB88d357[2JW6M[_
ANR?e^2SXK@YA>0GR&_bHT.+EZW]e)>6/UCeD4-OUMYb.CC2&0T_3cXG5/S?cM0e
XSNP,H]U<J3].C-B31.geGcC(,3Bf06R&d0ebLG;\;.ag)5=[KbDU,DO=+#E-K;A
JWcM(2ET;&2E[E2_>A.g^Vd@UXf]59-2=3,7dW/WXTQIdd)(>]N(AQ7DgaIBY,/+
+F26?S\KD&8N]&ad8b3L3SI],5DHQV:7[eZ@NO<9M+&ZI+S_U-QIcODR@Nc0A[+,
\bE/WBJZ)Tb:\8BN\/L4BFJ]-\#LX5WN62>eUQTF^@^Rbd:ZeZ)NKX,B>JZEMY0K
CWLa3CT&=8A,N@K\L>7e6Y>8=I8;f>LH-5-8:eN-A@S5\W4+dbRW[>Jd(&RK9QJ5
9=6EU0F_2<5SbFKA2V1#-dcM:]F/-J^[7-1V5-^-S.cgELgdZBX-eT2gO_K.T-YZ
X=cG&4MN-LN+W59@AcB/HJXSAKP?Dd7:cHM>0R[<Y9Q9[_W^a9^#a@@c^L/QO(,g
=/M[aX]DZKRXS>7H^T@>gRbQ-B^=@9M\)HURLga0NB\3<TbGD76.(W4;A@UB-RLU
#7fM41DGX=D5Bf6N2Y>PZP39I^Q-7ca4E4c\;+SJ)/G+)+QTK5KY99fa5YBLD_E<
eQ6?[XRZ>c(46#;?C_Y?U3G?2Z=9\7U/g(_8GEY\+PGE#80fVM2_2Y3WXVO@^FE6
@XLbO\[K\Gf9CWR],L)WZLQOS2c&aVE^&Y36>&0#\f_BL?/4WCIQffIbY__B:CE3
2=gZ9WE#/O@@/#&#P@f_5@:05Q6/7e2/YJX[?AGG&#3(S9UQ[82)O+eR=+JY<)4(
dWZ#AZ+OR,6Be&:_N.QJO)\(H3&;Z5a<QQAF)<63Z5?1b4A265M8FKE4H<P&DP.8
(N9Yg1-Y;2[48&P]C;FEJ+34eX3S)N),c&N_#a/IQa\3bg[C+<;F5[\3bC0NT8&T
\fKeVa6+,S@Z_1M..g.N>;LbR5>A.e^CaO+X,WR?X_25PQO5F<R)=WJHOGFIMOd^
f=,V&G<P&GDUb+/L?X]BTDGJ,4/,>T:W3f2:PXQ0LQ4+27[RKNc]^I_URQ2fc^=2
NeWAc>@1D5UJ5[C9)IGCNN0/E);WR^+^M[<J@&<+Id#.0NW(^1GDD8b-0,:9Zb4H
AS027d5UbENHW9.K<fgX_EJ.W^@W6U/^K:5<=C42YO@E5VD<\]2d-S08fa).Zb32
U)4b>+BIZACgS1C\\E..8J-\.UFQW5Yf-0=0I6gDF_]>Q8IKM]UaZ<,[<NBM3da1
=XGJWE=:([@IGC+#NcXf0QAGJ@FffF;D?QK=;Y>Q?=16Bg36S+&.XXYg^CfJ=g:a
M)X3f6UTMU:QU@-7ab=)]1cT-DIf+\WDB(_#>A4#C)NPDWD\@\3DH]2::bO.B[9?
_5/JPSGX7;GK722EME/U]-X?:[6FS-XY[6Ug[2FJbF5Fg.CK.&[KZ&efC8f&SU(d
?;YM\\4\aaXQZ6NIMY5e&C>a(LVVMU;[-b0B8<JfNC3eOff(_VDaJ-TSLB&RW<[Y
<?JL3+a>&VN8?HKOVA>aWHD3:6GARPZa?Y&]X>@0:ba//KT57@a3-O9Eg/CAK_96
=-BHA.SQQ+GJ\.@\^6@9L-DZMB_gb01BKR3a;fG;^=42>3YSRO:F>-A)4<U-/TOZ
1SUJRAd_BEH]aaRL<P6J[F;4P@6+:YAXAH[S+]R7R2R^#I=GRUX@Tg93YZDD<JCT
)adbcQI)2]+M4,&BY2@=^QVRa1e\4fE)_YcT@fKX=+793UYeYWO2=&_K98FZV9<8
::.Y,X7&R3;d@=NZ&+0Y.a4,.0XEF[7PY3B.B(9UYebHXTd6CEe71?g5IccBC\-;
f[5\_JH/Z.)C&H:1?RV.P3TAbX][?9A=5cDg:MCL/0JC]b^B<U&Eb;&9C_bfOI@;
G_ML@6[_f^8:7d#2<g<Q@Z-\V/FCIId?D9F:_3H?><W#,5gDcBW2+T&IAbL,VS,)
U;7[aFD#VDS;g,K=?:MYe#RF46:-Ib&R7,b/_7A]bK7M5JbL[C\PRBX7P,Z(_&47
T@edP_-06)c@/(&+NXKf,6a_9#W^?Y<XR,WU\OVV[XUDU1BIWJgaRO02;\PPP^H=
,(CaDgJDC2(+19a,1F/b:0Y6eFHPaF9HH5RW59?ReZ_C#W[N\77&fM&O,EY527;A
S)1:eM6#X;M)>&Y@MeHL_>1P3f#V\WeA&9L0]?8-[2:/A_QN&9CK14feaM5@g8T+
2X<Be(MDP0U@4f.O2Ofd(H120M57R?1T,C.>2WI2L8H;NO[S;)^gPK1BXOQ^[(3)
1^;8GA]PIXGa^[;:gK:62ML,gE;b-U[YW:U5g+[V4.(91S3[02X=_T0:,8AQ#SV?
CP8eR5D.bU6+,1:W)&DE1>dK6L@=Ag1HS;]^=f>2Q=c?R86Y#:9[(FdNF.LN3^bf
],F#OU(?&\.POAJ2L5f^9V@XH-TUU(^WJ5=CA]-1CNRAN@23dW^E\;2\K3D#d85N
4abcFC\GEL-6IW5,f[VOL):\fL?:4Z]JS:4f=]g>+JOQ]M<<L=<-N3>9J-PDZLOK
+VPeNZPRJ2IA>=A^-+3QbLR7562b@C<:25:N3+:7P<TPURM+0.S?&WTTc;7(]#ZV
LfYEd^><:>OK1c@Q2)bOQ2(:3DTH5bQ?J6N/g>fWCW4JK&^G/eBCQ&N_&.[f=4B]
eOYgXFNKHcU76OQ^TDPUF5aZ<1NIcGU<b2@^I8NE9OCU@D9GI(,:NgJ+AGcGY@dC
LJ__5C:50dFNbc,QLf7]::A7?_EZS85c#bN46[FD+1Af8Y.4FD):<@3::#TA:,[OT$
`endprotected

`protected
TB4U,Q>+fM8:W=Zg92E5.S-\K&U:=[+@gd]3=+&P0e>G(Ff<[Od9.)Wc;&a?N6KD
]L^;:;2P^H9:.$
`endprotected

//vcs_lic_vip_protect
  `protected
.=G[KT/SVPX)1^=&-E:9<7+FUCZ#9L]OVF]G#]++H9<A?QE@2REd4(_N)O<#d_Jc
gM:gGL@H#FU3(]]UVQX=>P)_W]&]>V9I+KA&@S0gC/8[CTXB4[1f>QG384V8g[^8
YFaV<-XfS,(_Y<g:4U<dD8/2fgY=W).EJ(&AJIAYG>/G-7NA8]EdJ6;Q9--6PQ^g
,MG=&3d:IHZc\(X:@\.+65S-(SYd@Yc@4(e4fWBa;F\P];cb(GAV<YOV3QC3S#28
CM<>4NeWZOFAZTE6)^\\1\aOU28<RQ95UNS:?Hfe-@a\A=[bY\_LTcAN;bLMGNZe
^SJfH#H,];K&/GGgY.ZTE\TRV33_EZ;_cScgI(>Ha(S-8EG];A;;SD#]J7;>DRM9
=Y5(--R;[EKOFeL,3B&O8dM3WJFc9f1QNUX,\XE.UfMde@P-RPI.:YXDN]QOF#g_
5+W_W[ea]?(ERWXg[1JU2U)(_N=_]XUE3#XLc_P(5.>[()BR>3\=KLFNK4LF#>?3
dRUfM9)LE?A--_Zb9ZA3?faI+;1,HB:/.Gg>?6g@MUZH:H+_N,5?^_6:&ECacIOK
N:(1aR)^^#,1UZ)b3##QV44A2;cAf,:.]R-a_9@1QJ)cC>;?(RW5\TA72SJ.O>Y:
\?AWG2SaaG4FDZ(T,F@LFG\e^I]cHW1#cWaL:3F5#5D0HNAZLgA.P_EM[QBH>_OW
@7JT+YVW;Q_cC_a;_^Nd9=6[,KMKV>:YI34C,3=O=RDB82=acV?U7b_MIV_ILd6B
U]6.90FLRZZ5+I,f0:eg](UOOf@e/T#-XdLF.HZ,Zf0X?1HX:KOA7QY=bg=SG8\e
13H:d#8:cF&OC?&bO_:FSbg3;83S[_4cXcS)/J4gZ+&gU\A]GI4[2eQVcU;FV>EG
aaEY_ROFY7.:KA++.:.EBb7:EE;AY8/HSC3=0\@cHS.UT8Y\4VEKX5P./78ZT?MJ
Rg+c-X7A6LgL)K#LQd\]PgGU&YHN)S;Jf<7c8TPC/a\Ha+C>8]?&SFZXKW3N^#6]
\R/:EBL:;:2eOJMQc]&[>dg0fDQSJ6Rc2a5&3OBWbeM59gK9-)f[-CK7CP#Sd3:f
A(>.^-3e<a2X]RCaEAbX_KgSKc&XTCC:K#P98MNKf[E;(@P)R0/=_cZ/H8I1FTOW
XS>H=@7^C;(a.+[ZSY2.8@:BDS+<<fIM8C9EXIeB?6EY8)]DHFFK\\9Q19TS49b5
:UH0(LX(HGT.9E>N^<UZ6MWbEUY?dS7c5A.@PLPI^K3afX=U3gQQQ<S[&S5fN&5(
VP>=&:Gd>@:]aT+AcAQa4,<.LZ4IB>VWS;=5X\I+8&Z)36_B3bdB;S<ME(FeJQ,A
R]#((7Z2<B/Kb77FS@Mc0,Y(-_)(G;H-SX@K6#,=D\1^I)VV[YLGYa<Q)=@DL^#6
)<9YGUR,C9+@4UG7]).P.g1a_LH=CN<^gbDNa>R6fI/:O+<I8H^^f@dD4>2WYQ,g
BABaQ(B]8Eg[F-]DWSM)C_d)Q<(+QW&Mf69[1/PgZV<e>,8;[f.#:b[#9JM1]#;]
T-\JNKb,NSD1D/f2<HGV@_4I<+OAHR[G4WH4-FID6>)G&;&PG>1Q]EcA-O/25:0b
=X1UZ\eZEMD&>H>5JJf]8\<:&WgefF4NFaM7gLdL^UYGE8e1#P]JOF0SC^&0R9\;
<1I]E9NE2[de\?B<8E:8KeF3OM<]9J6_]&CEHg(:T\G\F>;NZe^AKc.F2G+6DX:J
VM7bUO.P_YMULZ>PcK>/U+N^e,d.H&;V@1QcUT2Y.]&R9c86+G9H1O]Z2VD&3-Ng
Gb>(RUSH1\-deDE8M:8:VVM]P,P2V/V6Z&T\#2af)P9Ha:U7N-M2UF&dd\A3:VMf
4Nf7Q4L#(?@dV47BBJ3VO1/EPP732C>C+DAK[XFH?WP-JW>.=UM]L)A>e8^&E9+Q
dLXRJ4J#CbB]EI_-[?\W_=]M)KeL>K\T2<Q@LG_\>4=Jc#\-8HL+9CaRB4G[+?N7
VE=+FdG3dYJO4SZC\&gZ7J>59LQB8N]S<MVd3O[VbLd]LG^S?;Cc&#BQKM4@:LLa
3U:-X:+EbE59GMgPD8@0VIOgTL5e2F8SR@<D)RV=SI0;cVF:c(aMHVF[O?bK#V>?
:PA6/AE7TN=dLN(T(Cg^3PT/_a6HL0gg:7Y1^PI#XS><;g:5H4g>JQ=GOf[=)EMJ
/]#YfB7,^cA/M@+1Q4)&;354c9M=Cd/Y^H<g(CdQW2FS/1V?H<Z9I:(#(:C=J3\e
B5#XD#;32X([4GecW4>1UA@LL<#cWQG&/CQR/P(:WLC+AOG8TL.7O)Y7&+Z/@KC=
I66g>X+gTP8-43ff-FIL_WQ(UWcbLK@4[=aPJN+A7:&Y4dOeT]1[6ZCI7#=:)I,J
8d\9VF]:d6W.(:[W=7&P>9[4FRN,<+2b#A>gA0Ug?36FB0P]<a9.7P;D\0RG:<B1
WPK[H]G6M<bc<4N6>Z]>EF@@gV6[IUCSgcUBDJdQ@e8XbC2+FYd,C[\8=.EC7dPA
@TONG\K7Y8_,RU^G3^ED#\JNK7C(W?L\d4.>C4&DJc?,Z#FB6\4?_C1b9:XWDT1N
e(;eFTP6/OLP6)]YfU4JXc>B,7):D1X0aL[g]]Nb+KCf\3HdfMJRG:#Q@(O(-U5D
OPLL?LR\K[TD<GY](F39Fe.7]SO6)#=60E.e:T+=2?=/<HK:L>4>NET.1D,1Ab]K
RdB_13&DWWVFKY)6NFYV67R3CNe/4Y4\^LAS,_]HBA)R9==?aYKG>8OU;4-9=g:]
-;74(e=?dF[/(eRMId(.<H+QE]I@G^cD\V]9395gV#\;FAKR#:C/YDH8d>:PbS6g
OPK,&9G7<]/.B82ec.TG\KV2PLP_d;4NLE^<=HYa[31=WXMg&)Q_;5K-^T.gHG;-
F1cM^-^QH(;]:?e)F(-]=DS+c7\EA]<G@#8B1Ggd.\1cJ>agIEHaR?(UdIT70[(G
8,2(WZ3TV.7\U+,)W:-:0Y/(A@>Y(8.-]]b?RF=ceK;;PF.RS2IeePPP#\#.4PY\
U5Kc;E==USc)K1B2\._e,A@M+^^gHWT5AGcf5RW;YV]F<F,)D#(+KLRTd28,+=D-
A<?>71c6++ML2QGg2b:PC8N/_6F?CHXIL@SS7V>7Sa<cXOVH@WSOcDdAVG+=4BIa
.>3(DX)e=CQMNH#[b+0e(IMTcdfWeYLd-3_N-a^3[]C;.E2Ja@+KA9EU^-B4G\>R
+M,I=\OXaT)5g0RaJ?,&eb_LWJ95c(&U,===6D3Xa^794/GD5,&d/1]NcLE^S&\J
NY57@3X4EfSO2_+[4bK7[K32T;D)WR#RNF#(_ec.3?E]g(KU?2:TK7SNHd[b#c2J
H)d(SIADcM90c>^WJ^@2)aX3=<JW3ED3^6^+GL[U\/9R-M_;1Hdg^GEMZI+PFS7N
0;R9egVX.HZ4IS/d7_c\7cg&T-XeI/S6ea0b#dYZN@dLR.G_9g&))6^<NaF13MPe
>9YY&=dH>63Q2.:54;N@1B>A4B+,6,YU]1f:F,QOB?g3d/WJR=<f@/:B&0[?9c\B
IZge.U6R&ZdJ7(H?O6<?7.<Ig(\M4]LWJ3/E34E@b-,\3Ug<fA)e9+-&=^F+38A)
6MR9bFda135Z;7(AbcMM^<TOYDb(K;1BIeed5F2]H4O=ME?XgH0e6Cd.E[VIYT9Y
BTTC^&\N_f#YI_^&E7A&J[^3#NW4W;X1]X]I,8K->N3=HMg@>II]&-)2QU=X0AX7
8=W4N:gK(U0?=FZ5^V&D=PUIaKZ(3Z4;VVX&7c6IM_&P/PI6\._@[P9[g?#2,Db-
@@gR>05fP#E5R_8GSGJ(=Rgbe/_/RO&G^AS&#TG?RLM6Y0S:\.7[M.+gV-C-J3]F
E_H+HE#J[9L\C/;6:9DbC<.;AHY>F&gUKSaBGa)Z>]_<(PgbPJ&ID)D<@47?\dOH
A[Y)TF>E_UWF7[04MfSf^\6/>/+X:Ya#)([)0QPHCYaXTM&cH/cJ__)]ca7[08T9
??)D&_+/VBba9(^B0.g+D1a0J>8X7N:3>.XL#TcT:73X)<4+3+_&OWW&a>SV:g]c
TOA.BPbE:QBODgc3333@2]aY1W5RPYQLF1H]Z<@O_LF>Q=aB7<EZ[D;SI>XI4:.M
M^9RVf2fO-WH1,PRD]DA8+G/M9A)0)X>/#ZHVE2+#/)N>C^eU?]W&YJ]g.c4QNMA
f98H.NL40[7/Z(;8Ag06[OPXBCbBXASZ/f2dPe(&0-4DdgOM1ZY/:cJ]K$
`endprotected

`protected
N7OM;JXBa+5>M:\AH<.EgbF\T#&_X1OVGW5)dO,K2Jb\_DR:9)T:-)R]?Fea?c_?
GagZ>A\ZUV.XfM6IQQP/.F=VdPg-880^9HaT9O-I.#VLG95@Q91?MZR]K$
`endprotected

//vcs_lic_vip_protect
  `protected
@5_dQPD]D\G4M;58T^UPX>d5_@SL]@X6G563G/1&IEIS]@>7X@)Q6(&B\8a0E_7,
\GdIeU.cUO[-ZDac.(1)UCW35bV6].[aISY;-&\NJg8+XY)2N2=QYGZG024J0891
EIUdc3&TL:WdeO#PR2+J:M/ADO=8/<,b0f\+_[ELId\7.4UJaO[[^bG]):9<I=;M
df2@XO<4L@\.&eVY8O-),BDV#A\3MDeWX-?M:dY2)3,,T^NBEV0HH76J9.7+J3K^
UV9234MO)8PQF,fIMTA\[GNa2BARL,4FKgZQ1Yaf0=X)916OH)/DaV9NI]3]QY5e
)Vac>=C+UbQP3DBSe_/#[-AH[aN=#&[Qa#D+;F1=3;\Dg+dB8F/[6,J&48(S];#4
N6A2(Z_Q8=3=SU5K7+D&N).?32TV6b4P\^LK2LO+RMOgC.SDfYXYG4&?O+#[:^HK
;[7NLa8-:89Z\.2&Gd<O=IDN&T^=5,/f/I:IAF\^@WKH8=.0>3^6S>+R[WMJZe56
O<0g5ND/E4Nb]#US5)Lf9f^)ed087>XYbM5.1L[ZQL<\D\R>7,61FYD#UI/NFF/#
?NGVRe\Y7JNPPeW28ENb\#)cT+N9/HOW??HV0J7]&4CD9SORdgXUOe>+VB,QOb?;
)Zg(]N^Y5Y,ddaFaZEEH[S:(MR;)3[g9[+S+f<dN-=\[)a7We#VX<^JXMG&+&:&Q
IW:M+11Cf9+1X]5_D1^RPY^>S:)-P^e-J@AGK.K[\+bb7I>2JbK4>96#)JQO_3DM
L8@@/&ZNIWVaacU=bPEW<W,S[>/>I+b/f#WE#ccB5CA\JTbSM>;C8S]49?CC\FCD
XPTHDg-\Sf]7f1[>Y#CQJB/<L,a;XZTTOJ6Qb335[#A4#CGa#4[PY[5:;fA;GV?)
C/RE]>0fS<H2;3U.:+G)aUc)?<^#J3(]<S+-@<1+T/24B#>aI=6^X#P?.Q/]0cbX
I#VM+.?H3_9FI?@9GQ7VO_b>\/FDN)Zg:D?QA[]KHW=)AgPS,F/7(<_XX<HKKYfN
0WA2f7Z3b>b6=^>]TE0C98@L_J&Y>dP9H6]5QTgg]>P7V)I2d^MRScFU+3H?Z-<M
_W;XG\BeUAD&26gUK+7RV_Ae@UaAMN;XedP4f5.XF;Z<E1U5@cD9)/QF=dE33L)@
c7HfUBVbWd3V7&Ug&g#HG]fL^bJcR#?K:g(J@S7gT@Y^JK<A^^F-BMGeM@2R5ccO
;d\[]<?b.41/B7_N6P?b\<TF^E+_6\A7RQ\([\b;.3GE5/0dQCf]KS7H,^F4((]K
);R8.&,aSZ.EF]KWU(HHJ:IX<:VOHMgeIS\D#(f;f]ZfA&J\SD&/#\TYZECH6c.;
-A?[[8-g9#PRgRCI6X=?e81_6,9<9>S&8gf-)M-#/OE1Bd;:)DOCF^CA2)fY=<dX
[AAGOMXMc-7+&D-NEcY?Z1AF)A83:XN1K;^QDg^4?=#)9,O9\X0_.7d^R:Y1[JfR
gf\eJ9S7H;KZ59:<?Y0WJ2Z]F&JE:V,f#V10(3OCg0OYeN./JGBR#7+0T+Z0;41-
F3Z98@c8SJE.Z>;V#2XZNX;CW7fH02e3TSUP5;d/L^J_-(=MSQcWD:Nb=U.ES3Jg
I..Q5N-Y?7;e4VCUWV-O.K?Sg<g9;NNR5(OHdRC3g5S&^0&1\VWc.>6SEK6G\S.0
?4ab/7ee7]aV3d?YH+7+M(aCc8;M,<0Nf,IaW4.I1[#^@J/2)&/W392S@??W9=B-
SNXF)&_XF-(FX7:Z?_CA)-S,_RKIXX.(Y[[JKJ>.U[E+WGY>CNM4:#;L[eePEXHW
A1b9f)R)-2+AaI)Ne[V+)A,+#QLW+ffVdSbE>9##PN<G/V&<+&e9TcIE___MIa\V
.@JV-\e)d5A7?Cf6JEO+TLLF,CDL=UU)P1?94<eXD4fAeI4Q1W/fC,4JT0BVIL7I
[<;^\_3:LRM33JWOB+0BHU5URGNJRe>L17eY(F;_<RNN<+)1.GcF3K1ZM#K?TIR+
741aEDI>/f<AM\gTf6T7a6EC.T;CJ-OA&b5T7;3cH(.WZfY;>4?78_U_C=)ZDgO7
aP[Sf6?(,8D:77I_Q:g.QYEC5$
`endprotected

`protected
))JZFAR65NCT0):][&WT/[M2UBAbdOAe(&Q]21H+Y3D@e5R7EJG-6)).P#+]0L]A
PXB(dPT8JZ^.GD1<NWZ;H]aULbD:TUECCKc04&K?))6@C$
`endprotected

//vcs_lic_vip_protect
  `protected
NB?]QWRDAMe[^@(:ZB4^+-.&2UD+IHH,OM?/gBac<[DD_e3#a8O&/(3_&[N&BQQ0
<#38\fO7GQ[9HA/1C5V_A-A:.N;V^JQGHKaZ][:J#Z,[<<aKa<,:f63.D5.T]LIP
V,R2@IMQRa;[^G\AJP[T@#D[DSUGLbG.--7G\M1XQXY3;Z5b>-.-1&#=L)b=B:0I
45##c&70Zf_c3H1JIgd4a(;4M3/1,cGA^f5/e\E34#BT,1/7Na(&F2W(O6G7)7<F
cKIfW#^DG+R@2[CK]&=4c/(J6,eF<OMb+CU\MVA##H4-U]95TC^CXae)?\+cOG6R
O6;V?@1+F=_b+ZDC/Ia[>#14c22CP;4R,98XbXH4d1cd2H3:a5f?<KK4CBbPg]MH
9+9W<WAgeM,;<?A;=5WF]6;WU]ZdH+0(3[1K>GZN,Ee6gED[]=_PL>d>d^/YT.QX
+bNAR8BHD>N/_U;aIa\AZ;+216<.;OVgH@E??+4:<Q[7)ReMCAag:;=d0Y/W/(->
RY#9)3,.Y9Ib7S#d(V6H8<5aITEgRa7/U2-<GSGcD0S1,P,H\ZM>0\UFKbCJeNPd
S[[D<N)bSSf+Z]e-S[P1Tc@;(S??]FK8OJ[4?)cBB)=7>\5e\#ad.\MPG5]d&.=C
(G=Y;Ec3Og>+A_)XGCS8E,_RZ9f.#C/a9(+#C3]BT.0MW0LMX8K\@1=O]I=f\IDF
&NGa<E2EDDXQO7LI2SCOE9_R2$
`endprotected

`protected
.1C8,H5WZ,?@N#\:/\Oagf20Df_d0^@.NU2R1W[<2_V:>7AH0A6f0)\SF-P9/fNB
N/QZ=J0P9>^P1#^:9e\DG6206$
`endprotected

//vcs_lic_vip_protect
  `protected
,YP39cg+d3[[eY\NY,S+aS,5K0G1Og:e;Q>M_a<2Y<D&M<Rg?9A46(:)PP>TZR&W
QPLQ,0<WSDW8^&=4?AXZY[_3>F=C_g\GJ+,44(@Y)0]e6.B]-6G&81_DN2Db\cP<
F-&S\U8?CB1+DIgQ>W)-YTKAJ=7fN4df>-4:3D16FWS)ePLWDT^[MO\#(UUB]1@H
c:@=CWGEMJA-Z?\52&4\0;PLNFEEZ&MD3EDaDN^ec>XY_[YH>,/MO.YMd/+^1=.1
c>c7-+FZO:CFO,TU]_cT/GReKcSgW.b48d?><bbYeEX^S=eT[>\aN2aBYf@TaD6\
JW,(F)?#OPDfY:&/PS)L<WTFbM[Cdg12ccPZD_G?:I?g,3/a3Ga=D=J4DBX6D((K
IQ@89QBBX9eaV\_;:7>MdV#NaT+NYBJZ9FG<).2>@22@ObQd)8[Q^A4KYZ,f,b;9
FU;gaG/eRR#d8:_T>OI+0g>[I\\Ge3]4]T^)P+;>/&?MM1)+3961We5())4V?SRP
HM5X7NCZ0\_c8CJQ6@IRT3[]Aeb8H[=NT4BNGI)>d6EM#A6)[^Af?8-WeT:MFMINS$
`endprotected

`protected
K>6Q5F2OJ]f]bJR0OTgIcBMcQI[E6V]VSWE,[C0-53ZJ3V3>#FH3))F[5]1YH>L?
,MGA)0UJ-1>5&-4=<f8NSEMc8$
`endprotected

//vcs_lic_vip_protect
  `protected
7^S]689S//0C_HeJJN/I?]GG.4>DB<&a#._+6#4Md5B>S0S0,G7L5(2aU:Wg/\MF
b3Q#06.]MfN_D6Y?147YCL8(AAYP@,fcWK2009DLI(Q((/aaAbF:[?(e)O(bXc,g
BLC7DHX-g-U(S8TJ9<EeN(6c40V]g(]/,e1EN;S]#e6\I477D2#>7Pg8X.?AAM5&
fMBfXe+]K+Y,PK,D,BKNE#^I0O+#eG2(JIX#0#E.N_[LY_?A>:W@G<7#M+54b\[4
+2B-@47Ie+S8?Mf):fXZ_4676S^:=.W22=8gT154Q[gb]a+8(6ZA,(\?TO__RCQQ
E,A^<5_gO,&X5HE;IRa7N28)-5[NfWb54A/B+K0&K4()KAW5+UW+g(4M)95O<ZB/
:bD2&DXK5=EI2PWG;H8BM</;(+V&VG5WI^HTaD;]6O_@H41BRA8/6_F8aX&;)Lbg
Xc,Uc(\EU)DZb4M3#7,c#BDS<,@G4&[)58CbCJ;(H-5E<TADd[b68S5Me^.aICO]
Cd)?B.W^1]U[5;e6LYeU\54+_1+W;]Le:d/\SOf^C@MW8f3N8GE(Q8.-Y=b_CMc\
)T?e>/FRUW4GY(.#.YQ?aV;]BAB&(EQ0,#B)[#B4V[&;EHQVLgfZQJ/.R]ZOdG,6
#IB.-faZ7BXHY-/<E66CSLJ<CdH7bdTWQSaHHE2#HX:3UX]#BXQ=7=6;5DEJ>VAQ
]?a@dOTZZN-L]V,I4^_f<dM0K7(3QR8X(AZR^RP?+K=V#f-Q\FbJWG+RNcKL#CD]
M:J37/7HY],]_RP=[Q2\A?9)I_eQXR2&#M=L5Ja))YR1g]GGRKGSD)=]+LeT,X;;
<H(VUY9d#_4Mcg2/a[E^^F?/V=ZLH,XK0+W0<.GLDYW_eW@+fT?:_X#gV/e,M;Bc
M0a_d-HPS^R#K7Ue5\g;0=USE=143IZ9e(3/[-W4D2>2;>EXOA=3;K<MJ3^(;3P+
:AYag2D0S#DCBQQSPCbN7E[:YUP5^ULCLd<ScQ;+@A3Lc&H(59EXg5<?9\E/>C63
FND<K)@d#&=\M,2dQURHHBebc0;=V+I(JW/0[;BT5>Q@O^[?:@-.@OV,M<P&,/0H
V^Pa&f(KXK.#59EUA69V.#.<ag.-Z^1,G>aeQ2:&S\R/CJ;^H/>&K;Z1g^@\_L8+
;,F-9DV&+.g86O5Z(>J^X:2CVPUARg9XF;N6/5.ISN^,2;+A&_??>8#9-X=^;)W4
)FgIC1VHC9>34+F-JA>;PM/B&f[I/CBRRgJ,4g4#9U^d;&U4YGI?2[83d5dc3>Kg
SY8A9U&SCI<AEA/5Uf;D3Va];A=Z7b\E-_GD1LUcJIK:MEFDJ8N[[gN-,DP829;]
g/RV-8#+)<[B7N8:M+J_]fD[E^GV@CVW#[2GRb&U3DH^e4JI.@7e1MK1#L0)6:d=
(:47I/@e:ON_1b&J&NFXcQ1;2(M\BYc(=dAN);@SHXe/,.&83HJa>J96+ZG8O+S3
]0:NX+8[-\Ge#C_XEPW?&Y_0NFCH85_<TZbaUE[S@?17D85V,,^BK\=L6N+;JUM)
GNLB\G#?QD+9;-2aBWRf)_a2UeRCB=<93^@Y40Sb;NX7@/[L7G<,)c_?GTCbBXQ\
cS^WXIUNW:-[Z)XUcM=MNU=b57Ccd(OB>T^HK>(bVC5HRGa(NTVEELB2cQ(J:<NP
a]@^EH]0TI02GN8DQC#eMf)UGHD1PGdA]0SBSE1\T@e);8(MN94Vf\T9[If0e(:@V$
`endprotected

`protected
+<I3&3YB;AaSfP(#H66@Y^KL]:#687P@#/a0_.US1L_f^G0Q#H,]-)eN3Z2[#0)>
C,A[eVHe6dP69G/P\,@9IRKL6$
`endprotected

//vcs_lic_vip_protect
  `protected
[Cg^MOZ89>YVK@WB/,;A#FQ/Xc_B&JW>V0GHXbPI+9;1SKQW=L024(^Q-AacDY?M
g[Z8LQ6aK(/b-V<#L1C#c]Z5,HCBAL9PA.9OC_+-_7cMQX60IL<T&)Pb1eUG.d]I
f<Lf;AS2N-[:Pb1@,;8aFSCHHOG:O)Q/FVU]Pc;^1=(<\#:7<^LQVMZPQ,HGf/-1
5Z)V-LY+dB?:)E>QXB4SIYLYV.2/1K\A?EbPWdHe>NF.=I>NUbBeON@07.VN,NAL
?dH8^MH-Y+Z7,\@.+Cf8C?2,+K;(+2_)T=L\@6fTX_^c]TSALRgE+<O9RNDc:LD[
#FLNO8E9OW2QH?9N&@=f3@Y&__]_fFc<c:45;d8ZM@(8#1K<KMa.C\cGAb:.]T\#
;O]<)\3UgYCYE1@K6BH<<;]C>SYf]+CcBg]M2F?:F1L/6+^#>.U)9ZU+_U;\FB6\
bEg=ZA=KSA&+1Q]A#?]QU=6JM-4Z@>T8TNa/b=6Lgc>3IT+;Q-_)T2@TgG>I58L;
:#U_K-BcJ?5+5a:>)\X&_0IB3g3#eX&NT>+AF#=7g<O_(FdXI>eP@8KNL\ef87))
dKYANN+=9L:fa=)=TD)E;@ZCP]B(?V5DR0W;GUNFZ]?AHD[.N(WM>C#FJW@&EWIB
eY^3ZDe1,UMaV]4\QgeNIET)aM-<._0+;YX;FT3C]2PT33]7MP.VAf#T,;BMc,d:
NDUI9)2#bWa<9c?_1-2G3-[DcBT)e>8+ZJ#1CO=[A0H3=>A?aTF<c]Z=&8(DE4FP
K0QaJ(8>6W9<N@]3g&QU4TAR4F>P_.R)deP6RQdA8?+c3?D.;CNOfZ(OGeY0Je^_
0=^^gG@XV5>4?T2(F^Nb><cOJ7[.1O#3JH#_,DGUGF2S,T)-<H-.4Y/H4(bM3Y\X
+.b]d-a2dO:4EGH\2Y+?ZDTFG.9XS#>MC(\d52.0H&M2L;BUMAFE>V<VLA4U687[
c93CEN#<0A.#4EG2g<7K:#P_[9XX9_H?-RD4(;RH/8.2M1DZU#K-W6Z?I<+/?;5Y
(N.=87IO<IS]MA43]99<HaO?c\M_Q>;VZ0.2ZH&b78LR_D7(dg&T(bZ4WUJ,/MGV
f/,2M5N#T-9JV\9P(&H@gFBOI6W(3^98&U[c(],66f_Fba_)Vga5>-gKS]]KX:dG
aSWaB4FO^\KTPR8>#F5E;Pe5[:B#Xc&G0K&0]c[D6_84-OCP-&:#ZWE<F(0O7NYf
7a1DR8f5V;#1W\f2_)9GB]NOZ;+9=^;<XLJ_g]32VD0F]27#2NC/&#O9Vg^0<cNU
O6P5A=K7HW5CYFV;:.Z)7VaX-NJ\=_\,FSPD76/;J:^-5NX4<b)1Z#5]#86aeZ^e
Aca6?]KU3>AF:<JdU.I^LOV4D95gNZU\WJ:KM0Ye8DIKAW).0OHM<1eCc2(RG0#T
HR_g(7B6(I_R;G+bC1^d=1A@Y#UMSfW1BM]Ld_Gg?1N[3Pd;7IZ@[gO)&W<F9fE2
B1#Va.FJ3.K#OEcCCQ-1:Rb,-4?A.E4);A[_9b3Mb;4[4]7ZSEK-B?VWBL4gW#0]
->Y4E//]B@Z3(CJ,JV6I/DaB=\3-;CK]MDg<?^:Q<>aW7MAg+7KbX_f+W0I,2DJ\
b8gM[@UW9[5g+OOP)dZ+)49\f5fHD\&3_.8]&IU.e(9+(BD0g1&8\\6;H=.34[OG
C(Qa&A?(UW.QU0#,/IQBOL)RTLV<I;]?OL@WN7-ZL3I]78VTEb3XYRIIEe;]_W#N
CF7fe3>5R^<d;@G;=()N&>,a(bNcc1gP&9DLU^A1Y2JgWSgIcEIH/1Nc+JJK&/GP
ABgVdIe;JHZKf(^VgE)).?ODLU\36V@=)8=L0IecTaSGfU()2U+dZ,+75+@&:&<B
_N8=50KR;9LXC[0]g-LOHC?<RWU(+bSROX&]EKVAV=6+W;4XV:HA<N7b+8])D00&
A4Y<d[NTX3,PYW]H3+e#CgG;FVB8NYN,AVM90@f(,,_aDPSQ2895U;C.WMX+U7=E
QOPW-W5I1&TA75Ga_3OgFMBI2MLD<#]DYJbC<dc7K7+:a/1(.XWcMJW@eG8=^d#g
J1c20WPG+[(@[C2\a5G-Cc(L>6JZ1a7b9(QQ1(\>4=X7//_)g72N8ag]@[?AY8AR
.?OYEWBgDU^;YYLUAC;NQXc4INH7LC0.T)a])64\RCCI0&=c6M7B6ef+,DV9E/YB
(-c[#<V6@?SMRN8\(TYPVC6^#.MEJ9,2&WW39[++BU6R&28EOKY1RZ&Y[E&F[g30
?6E/g;6_^;0Sc@&7^.#=FCH0\a?8MST#cPXHbS99YK1Pe^-CZa@NGc0M;C,?5;dC
W@SB3V;+NfIVK@Fa9SecR<e<P[,/91^XfVLM4Nb:612)SRA+0GEfeC+\QKGCW8Lc
OZFHLUZYeHX:BV^W<G+7&A_dCNA_a?ZKZ4HE:/,5UNYXd13]2<GL(6>M,Lge.4[,
G&?4Ge0/LJ6F2H8(d>DBS<.;WK0eB(&J=afNR4<(862#T6F9?X[C0RVILVQ?[.Tb
;J9R5:I-/&J?B&Y0,,9=[d@WB#ZHAVRgGP84YM73^Y+?C/.;=N=0<R3)f\Y]ZE;b
=8-5BAO.FG]/c/E5OPb=@Jf_Md<B.S2W_I:3\V2T@)BX1RCc/NF[I()<\]4IAH5[
D?b-=HTA846a9.GV+\C7YCE1:>()V[U.Jg@O@COD6.I\@PR-[5b81T\KJ#JBgTCT
SV86N,4DK5H+1:#2[QFK0&PLXgE]dQOLP^+)5ddJ/:c0f8=M)P)e2f]:.K3b8_0M
/X:g)1>Ve(<2N)E-S1VaEcd=-<--SQ<a4f\K4,?7]VI(>M9gYK>&O1[.VB2>_Ug=
-JC;.#,++[AH#&8;3e2aX2OA]-c#\/RTD=X->:CD5Gf1.<P?I@K2,b1VKEIS/\^7
:NNe&7OQ_dE156/U-?BOA)C?gUN?RZTdgVb]PLe?3C@1f[C))Y.6(T>faZ[cS1#\
X4eb3RN_M^NO23PXGBgT1V-R?UT3@B8W:eIC_VH@21Z(NN>Q7N8OM_2bEJ=4Mb=S
f+K2#/[5D><O=&,G4F5Q_]2T0\\K(4C(YG.D=-5Bd-ZN_16T7:3U\:+/fKFOD@e\
#1dUdP[HA<^CIddaD0;X7cdZ;Ud6H&;5S/5AQBe>RE7SDafYET^Z_#@BeZWeOG_R
>;^E(?<U2(X.SDR@Z6SL^=b-RE@WQQ,Re5\4f.][C:cBO.c?.,J][C0OCK,#&Dc1
.^K0]TadSH-7AFP2L9.,[,S8V5D=&J1_&#=]BI]X@Z\#I+=?edSM>;1P:NNE6L(0
M3gE-aX6[A]_H[=H.PWB[>?g9Q<Q[?>C#6=f],JJA)\_;;OD>dJ3:e]:T5Ne7B.C
ad.4<WcGf(L0JRE/X[LOSAB58YaR#P?STR>53JP\bG.DNH+;#dXJ,L[]<0S<_M13
-+;@EPOW_GCG_R<6Q\)gc8Dd/39<:&(KQMW-gacCZ;LW:a,YO[E=N3AK_74f7(S4
TK-6?L)^_2Q]W\9WSE:g6cD=D5ga(-+5&.<H(aCfb&9>O@DDaJe=/c;#9O\gUURL
.#6/II:3Y_V)KZQ1>(#@FHMXb/AcP=<\>IM>&EeLBAS_L87[.5Qg(::J)b]CX3@#
_a5MK[@a8DOcF^.bUCa5:E;e?]<^XNGTe2g.Mf7AO>-4MTVD(3(2(/0^]YEVOO=H
3HGSEO4T=H:C:HX+^Z+?#e?eJ8D[BgaIIXAAIC6)VRLO]ETB_U5#5<;L-Ba[7bA8
E)M]UXCF93^X_T>;GG3L#,DWc#,)\8FMNTSeD/fBec.F5ee8;LS<H5#^2_H18HfI
#FTPD:=_I?7-L5RPf[(4:QXT[6eC^OX;5@L&K9@MX>O-X/EJ=WK/NX#M\HGQ<&PH
_&HCJ]G-4GYQ3:gWNY)_G>F6Y<I?4\F\IFWg8-93G3;/G18)J13Z>=+<\&5+0SCZ
,D2D:[:?Kd>GTK).RSQb+I@.]>&U.).=-f3&Ud,V>E^_Q=af#Q\T,=f=_6E+gJM8
=.)[+UW1bG\1(XGGKX\JNL.^>W:F4VKTbH.BHJ)d,WG8H:XFUGZ\7WV\6QD8MKQK
<Og;#6P5]c,BDW;&aQI@9?697;e_(PK:O40/f69#IGDO;gWg8[]#VDe/<MR3\b^@
;/aS,aM:(\)3afK9URO6N<>#V)S((Z^^T3U>BS3;N?-N?,9Q8;7<X9@9]c1,X\PR
_dAP7>QU@5(?#T?Q[OUdY5,D)gN)UUZ+ML^B^W99)C^U+=(UGNa7+7bC:_Z=b]44
(CO&:[Qe?WZGZ9D^GFKON?60=Q.=S2>HcfDI,Q11O\c7P]3,CKF9Nd0O_Nf<77H=
ZK3WHD;J&74TRJb=cPB675Ta\c+[\YfM.FPAU@AO1A\I&+K8@NW.#@YJWQ:NTde8
K2>>@F:BQKBQ8T=7CK39f\O5[@BTXCd,ML4,TFV_==Z]=fLBY.;O306=WVY&;0@^
PHZ6^FbO3[WefWA&Z,5YcMUN<KU0XBMYfX#2IMEfe(P@H:^JYDK63#)OLeAKe&/^
fZ955K?VV2dZAgWDMR2-b1;Qd]SG=)M+VD;T858/SR5;#P0@?9+Xg.(J)IT,/,gV
=LPC><ZbGfC-]EUP\6RUU;#GRDKD\WDQb#U/O_5EGLTdc=V@8+F9-AXDKB_2@YQc
=_&CO(>6+&g00G[\R7Q3JNFJHBddED723Zd-,>&#M=OP<2\&^(B6RB/31KaM4M1&
)I@L+9[5)&/^)^UB,@_2G@(:a.UYgAa]UZ2QbF7F1XE)(FHDTg5P7BA[C,[Z#=:(
Z7HSN&SQX^?(10N4?50bUSF157CLTdQaY]X(S<7C@)CJ8&P;GPTDL9TZfO6P^,4D
,))P6_>@cAV@T9f9Y)d-CMQX7SNf_?M81.2ZM3]98M-8C-1,aV#VcTZTGOX?#ge\
RLH#Y[<=@L6eL[.LN5>8CE8YY@K\JcCXgXCNcYWGD975E6.cc;CQcAP\=ER^[JLg
[:?L;^9OO]V?L1+FF/dMN-0aZB+Z_E:1MS3G7V2C?7,g09FEF>;fb_R8]IG?.2+(
L326_CQ(=LD]:e7[MO23DZ/S=?7/BHV?XAdNgX+49M#XTBK4dAW\L8DK=1a:[R)<
]YS;4J-1;g:WRHKeQ:,JSOSZ?REcTPZ#IF+?&OL]<6>1+ZVa5D7B5@gF,G8MKD[J
H@@.8\,5C7^I?^@1F5.URJ+17M>19#6f<d&7HP9)b4;R7YAP?XNB7>6Cd8=BJ(=#
<<INAfA3S(Va)]_\<Q_@eULG1dR/QGJVcM=RYc0+^/<LYOCRYUea2-MO#8K:9O=O
BS_=HTf7]AWdcE-.7?<_/1R8&gOM]P:E7bSf;O.-0CZY6g[@U?gM&HKGBD;,;9ZW
SHL)7R&P33DPB[)49,V66/R;#3OCWCF);Y5#5H8\Bg^4V<-USO5_:Q+/4YA8c.^f
GP-XbH+YQU/>9Y1+7FWS6@MKP9==4=+3Sb#IAca,CQ]@V)LZd,,:Y2bN>O[1,J]:
CQdXYQU(cVRQ+fJG45BS2@]BdFa^e)3Na2]Pabe&G^ZdWOGDO#4gVZ(7g^eHE62(
I1DU1&=e.Q);7T4DP1A+^T/1WIBLA4]L<@9V\0JED-L1L:Q:L,3d;W^Hd=b;,d4Z
&Ue??S3>B9<5G>8(\RGP<:U[<b5F5:aA.)KL&M[d>=N9R95=bC3#FX1Y1?_,I)1V
6#/W=-=30X(3CCfbG(](XH:9=.TFQb-/A+<-DP-2NV&7gSI,+7+L)\=c(4S_JI2[
d-,THebgK@EeM-F:WFC3-7M\K[HRcUB)85@2^F@A[#ML=cbT3E3S)UegYNAC@;_8
P^(CSfJVf;U5+S;G-DV<,WE?J5J3UC\4ZD8d>(cXS7(6<)<F>PMQd9QPQ,];@_B^
;<J)aR;L]F><X(FA2OG<=4FG;c/QRY:B+BT_X.UL=+;BbCQNK+-V/6RZSN/&G_=>
Z<GO2JW(]_]d1A)SbYf+))7YYPH-#7bbZ[/N+a6[PeTc&<DPc(J<69(aF].(cP:F
X&&QEcF[?[@\HD]/>RL7YcUS;Y@NS6UT8W1.BCdKgL?MW-X8L)UL8,91:-LP5;c]
.#_f]^S7=MHQMd\^aL4=9?5M41S3Z;2JT0T2)_.+Ce7.5:Y;M682U<I@HCI(Y\@B
<2Y>SP?E3B1A]EOF11b_:+.c\[?2[eJc/fBNJM)AIWY;K[J,9^].P#,VX.0@fA6;
KbWc4J<[YG2@VT_=eYb>Z3[ag3(-BPZIR-J7LPS:HF_c8C#0[3+/@c&bRKCIGJWc
76-L.]6]4f_)9\Y1S(VEG0aX7_&O=d7[fFLKL^DKF4bSK>K6)BXKW_U#V+g.G9&1
7.C>+4)X_KF;&agdg>?S[4Zf5^,BQc@P6.6\V97fIc.HR;C0@0Ma/IG?T.^LAXX^
:NR=0=>#++MUR&YK//Q3CK<X)OP>3YM?YW<UQO>\X3Z.MbK7TOFP,LRRBUf6:fGZ
4cWRI9;._0[8=1.ZGe+8=NJS^BDcd07&FZ53GQ5a>9b^A/13JWUSC?Ug([T<>N:+
,BX0BLDVEDQ&RN&W7D:]\Y,Q(=7R>^Y<;I+e8]6F47e+Kf^d),T=CNHGIA[c:5B<
)^>+:_EeZ:b,@O[>gCUF(DEMX&<O&OYJLZ4(ab(NXcd4XKU,K@eR/ReT\dM\UNIe
B+fggFM@R0F\FaMd+KA8+?X)X5@4S&)@G.EGG#<5\D(1UfM8e>c9\B]5Q=(-D?0U
=+#MBYQZ).M:WbYdIYMa6gA3O@/I<XE:H0)1#C.6:+gTbXB?;3b\83OJ-B2J,@)O
&38IXZ+X;)XZ2dPbO2C#N]N4gHNLfJc0QSOU6^c5.\C2_UZ[=F.AZZS32YL#Zc)c
8QBD[,2bY\\.7S>Q7_NbBW1(^S,EOUMZ?PNRXEPL#DX/AbgPD(C=9)@1b-#bH)R+
,&L,LO#N(Wc1OfZ(LOH:\5KWcC=__RIMYJM5E3dP0N6Na?fFJ<R(b<JIUAN^2a3&
\C?LN&R^NGII^+1E+b1QfJgIX^HQ1S;:&H)V1:M/_=ON]?L=6cA?[Q-/DWWIG._L
=8<<cN#&Na7SFPD<PM;)[V.UUNZ5(+SQ-UHBQBF_0O2<K<dT2aKZ92>CL47#ANJJ
f8GZ^9<7V)A.:QL]O+37;ESKX?eJ<3#BHc=Y84S7\eAFa>\a;JL]1)[B>,=-e+8D
ca=P9@(X#014>c)L5F;?faf_/Wg=b-NbN\A2LJ\8fV6TB;C;NIYP59]V<MW@fQ4-
MdE7b;6V:BTKEOFG0JCS63aOXAC+A&^77B3=NcfTC63\a[;.:47ALM(d6@#6+VdT
LTMbL#Hb59X-Z1K)^/MfW_6.W>.#fOLa1J^YY:DHTM@=4W(g#7D147a59dT#De&B
,>,S;(b4]/QQ>14L19KJTd;K_caK4VWN/UP(MNe.2P>X)^2,X9;3\YZ;&,gOOXa,
9L&[>>^ZQKZY>ZRV6XF4=gUFT+)ecAeRZ2NFJ7//,2L,U5+[V\ZeY[L1:B&=<KUd
SbV3A#FS<O#Y0FCG9?RGAXF+1a\06=<GJZUQ4DTN9_;d^>Z&6TN:BN<cebd#6cLP
g?\<@.,]d7:a08XV@8@X[#Y<eTH(Z7M](TJb^0?cE]TU6KE98=4)DbUY;(bUA6K,
Gg\E29=A\UX=(4bWDPO+fBWNC:Y4]O>gB8BG-f3UV9K+DFe_DSEC)BVMcKBQT1cg
(.#TW6FPW7KRPF&RQKJFYNONAQ@8N8dKaB,[gd/UFfWbM/4Da\;#fVV1bIV=OU]E
6HV1[S[\O>X;,YXV<T<@YAG7c)6e5.<Y.DL@KPSPS<+1[:Kg(E8[6P+/Q4:WKT(/
BT/@+873E0O<7\d[5MJQC7<(M&a&=<95_Q[QD^5\&eQ4aJ9]HXc@e1=BXefG._?Q
GJ1_Y<EOJ_Od12,7JGfR+/A7J-&J>J0#Q))#,(NY_Xa0a?>,WSa3=J?UVVA&J3/:
3.G<,:_PbeBYU_b,3OH8.;Fb1gX4=H/CY7Zc6aOCF=NHN;F(c4<=W8)T-4^0g^;E
[>DA-V]Tg:M>ZM^b3.C-ACZ8)Bg8?UIKCMUP#IG<K)OE3Qd:GHECV-(6C5)6c<GJ
,ZXLMMSVPg+.L#.#GX-N&::a)]6XcRP_^8CDILZUIAE)?V0Af;cbAR;@KTXPK.@_
bBD>FA@EL5=@(LB<Pc<ZWQ,XNMJ&&KYg&28LCUC[?FC<dK2XHcL.PPFNO\F30eb[
,eGNCQfcQ3X<(a,[WA+[N)NH\S+Z;BT,K.d]33=81_/N3&ZcJ]6X6CV[A1f:#J@R
MAR#+\]BY.fDA[VgB9=8#A/1d[]^Vf;:EQDQB6@)W8ID1^C:(Ef_G#C6L9G\dAO+
XB.(f3W,Z;T;9)ICI5A=T@baQXBaC?,7,C0_-[FR79Le7,:Z-0P)0Z;)BIDKNb:)
O8=:SK#A31Q>WS@2E2bD8d3I7MbDcIIETN2]RWSLRD?Z_6F?W#UPP6JVCUS[:8#6
2H=.d/\Y8M_G;d8-?g^3]E/6Z_4/FgJeJQHRL-J:<gJ;@X3)E5CbL5NQ0KISI;=;
43_f.;&TXCS-/2/#Q]SVPIb6ZD/FY6HNQND.Q/UL#=HTA,g+&53fDZ7.8/Q.]eZ<
WZ;107\DN[0/1@-C?H=M)JH>G+fH?G,=@44[-FEKX8L)[e&eX7J<LQ\=;X+f31=&
gU&P0;\K:cSS(Ba]H#MA;dgT-cN[)5_c-PV.2O<eG^-c4WbSI\a8E#@RBf]<I#;G
P&S3^H>f>4f\N^5?,Q^PTbg,&5b9VGK@2f5db&5XP@b.AV.-/E:T;^FSZAIEe(Sc
;UW8JF/]O.^,]7=;97VHM?7WA?Kd1V7+1_S[B>B5(O,b:6GP-TLP6d8+>@@gE<a^
[E&Ne.R:<)a_#^5LA?A9g0WLH,cbH#T,DPD#M0-]H?[S07M4+fd0?=BUg,,>^Jf4
@DHUK;XUNFK#aB:_6Sb#FMDdC)XbBJgTDe>V^O-I5G1gE(M8LaO_<WH?J:AC_cbS
8:b)7X4QP]534R7]<,,1.OD=/T,1_U_:_e[O4B59J(3M=Y?--BQB.]@-9>@Y<UY/
4b^VK9S+DWP2HF2J(]ONAS[YTeCf6-D(5(PD/_d,O_4PBRWKJ^X&OZB0O.52:@E+
(1&6L4X^^UONN1CL<Wd2OE4(F#?<G8bJ3HO,T:P:OF)ZLI(]<0Y]A#;O;.RA.gdY
,fU8HCK)C3T/1JbT2\)LGbT10.&EBL=Va5T#Bd81^\QbY+CAc@YR7WYMYJHT_eg#
3)?43#A/ec6C7&;>8LK)g>ML?R&BWB>9IC9SbFg7&>5+^P^?(Yd@3E<\?:+F06&@
6N^SDL+?F?@]:_,GM(#Z5D86GZ3UIQ?Z\ENO\e:X)(9_Fc1dC_\b71dW(\U/&9Ab
O-f37.dAaa_3Y]_XTd1CMca)55_^[;V[0L=I=QcD9?GPZ5+HWa@H#SEB&KAZN8+U
ZQV4f:7F:4@EA,\M7VTN#]O5\.RUA(\[/Z#^VfBQW-Q,@8/XY(T;.BZ3)aE>5]-(
<.T[bZa\d)7^deJR-<7fW0;=cBB<U&4WH7B#:;_S9^ZUOf2d^0WL[Wg>#A+e?\Nf
;O_LZIaBU7^C_M;0=8R2[]>S926ZU;,^+OU:^b@]eV/MDDZe3:509=eGDH=Q<CLT
/V\aYQKT)^)2?#,+MJ&X,NAA,/_1QfX)S9eSb>\=6_X[OZ)9a0H0#C5PJZ=-1V84
T>S36H@Wg;6F&-YA^D,VeRZ/:,HfF.P)?+aOMS]D:DJU3E?):MBCV_4HWQFTN&XS
N_#AdeCa]+d&/\&Y7.O7],gRM_7+T=7\]X+)@WfJYe5EPVQ5I)8RBeaEcM2Jg.#G
E[KU15cf/a17?#+YYR0@cI5FPQV=8EZW(>>S[U#P;ONST2]#&[G0>8_E8LgVJ)?\
CN80L50-Uc#d]c4N]X+5ee_C]R12,8K;]G71&TV1:,9S?XHM::W[?HaQ7bQCM,5O
P+WCRQPL.-_XE=dMCR/M6SQT41]S4\fLS1JY3NSW@L:XfH#I7;Aa>I\9>+M2=SW0
KBXf6SRF01LRP?]O&aV=/6OZ3:UWR_2NN9K^a@[[HFWRK045ZLDGGL=_HD=_HNNP
:\,@10Cg+3;)X0E99/TP;D<0I\3UMPQGK[7@6O[7I&X5CV[KU9IWQ4B>N:Z,G)S\
W17cKL;S17e\QL4\bB.UcT(&<3QW80+>@^L=LE?Q#?>Jd?5Tc&PJC[VRHJ1BFE)e
fGHbP>D)b]K^R4E2NS56)COBVXQ0Vc^V/b:U6-VH75+A&29ACFYG/3RHAML=.YC<
;S&6#X=LY&Ne7GeFR-Lg^R2:,7eedJUJ-.T5&cA)]@JK]IfX8Dc0K\?64Z)E&FW5
J@+P&f1d_;IeQ_(d9?PdKG-UH>HA#d09S((R7&#JCVN_Cf.@RHaO[MA;Kb1I7)Xf
@6N0\QJ2J0V;U70DERK\Q1.ZI:UF1>X5R+E]LJ7F0.UD3Bg8_d_@D0:/8MJ52]&B
2WS\UM<,Q0XP=S<97gd<WE4,IM54,(L6+AGgZSM@D-JM6P@.IOVGdPV2^2M?9?2C
a[GTPFYF:OLgWV,X1QHSCYW4gWe,)d>2^MSb6J=bI>HXTf=L];67f9?2H,WE(JJL
\YaN=9dG^Ec#\cd.-J:F351E7<c34^1IE/95V.4KBceN@V@1DA-VM=\R[;BJ:VTC
6,XC[cYbgH?DH4NR_WS:BJ89,P-XcEU[Z##05N\G=Ob@c\c4/b#K<N:W9d2LXK3]
^K(0YT=NQW]Db0MB&SXLaRLd>[aB2Rb037IY#bZQe\=_I<;Sbe4PDS[73bS=&K:6
+HX4E);P<6Ae_@1&4=[=)1;3Z)a:V<1P:0?L>KC-@&NSa:fV81LRAD[_8-c/@@5&
d4WO8\]5TCfN?^4Q,]9b]?IVfYBd-6JZ:.7)>)3W2#6;6RYdL0L-07E2](;5,Bg,
5,Rf2Dg7.&7FUX>P<\d4Ta)RW_XG+c]Zd4LcAC)>HZLOd.^LD>.G]-T6Rcg]66a^
XMH^NC5+-0]@a.N?Q.D?)-Rg.8LYDA?7B9,cUZ=[DJRF.LMF[+-SW+0JfgP/C)[.
dAMP(OU7L42=LE]K02]F>_1.:S#12R>@K3??0.F,[)6V=^8>cRb=I03P<577T8Yf
Q2RD_M?#TQ/f@e2f8LG=<7E[]B&Z4f@Z>F:V](J>TAQ-<eA/QO1?6Z3WHJDAEJ#B
f0L))Qb+KFbPAUEC:I)R<E)A^Y2@E=1?S5MN98_TCMQD>UTP\SZMVEMaV(fP:1R^
<C27b;R^^Q;C@]BFFNaNKMCADANZ9UZ?AgT,_;F5DO_4[L-#MXXDBP_VRJF&J6\B
aT-0T-G[dBNB?1\^QQdaNB:,O9LZOMIgOO0Z?IPeL84?d(N1<JBK)UKS(&+O;DcP
#C+MWWCZZba)d1e7(636Eb^QZ=)4^;(8]S?/M1.13)3R[<M/?aP(:1eJO@I+<P.4
#R&dC9D0IdUHV6^XTABKV4Z5)6]cAf<>#@Z<ID3g\#?3J31f8Ffa-]W7b[MQZ30]
)ATYDPa:aWYHQS[6Q:ZC&2PMUG:^KA56QI/Q33F@(fJC08daL8T9;gB67[(2N(;O
&OT_EAF#YLe)cIGGR=8GT?IB5MbT8RP:AHd&dcV5VB99R2WT:c4dPDI1PCV?/_OZ
;GVVfcL-Q<I>D;BFfKL@2&&\AOSGc69EVUW_8=IGf18PG+RV3SdJQ;KDbXUB,\Q+
59F:=(/O[;81;=2_I&6F](4cMZ<QW&DbH7TC?Xd[5ZG>4b,RD+PZWF)TNP+0FcB0
Kf944cF@A27,VU+0OKgcQ=@Recc<\@D]5>:U@CJ_,^]g,-P:&1;D>N\a(N\Sf_NR
]FPFZOLTR>1e0&#1O(99AFQH&2R,_#FEDDGSLWc8R7I.JN=;MK@^+><6g(/<7XD8
USZWEKa4QL>:C4a.E:=^>_>GO2eX;(I@SdXeYfQ&JBD9XTKfM><3A1P[K-KWAf#e
2V9^gIGNAgDU:,e?X&A1YNBI0TPP7V_5L[&2>Z@<XBGL>>XBFN&,.:AO_[fDTbW2
0g\LWNZGDc4PMFg>7DM:8:^ZEX-L6A&;L6)QQ\XEaBBa+JKPA1?T;;KSLd[;)MSe
5C?bRbB1CV&0UbSeVc_P[HQF6\.E+b-JUX@EC&X,3b0<dMgWSA(20K.KdU&MP<cb
cI=Qc/5^.JQ]fL<-?;gQ(aa8]U<M@TVf6_=JRE]3Wea>DFWD:OI/04SR]>5G3YY?
4IVTBdEYMHAbK?QC7H5(VfS^.#/FB1I^J,P1D-CW5._W88,IO_H>H8bZ[#eUfACW
g1(^5^cA_P]K4V,=,e04[SX94/B2L[aMU&3SKd7^ROb/^MgAe2XZ/e3,LSIYHN8Z
Te+7Xc91,G\g8Ag@EQLO9MFQeT=+.STZP\eQJ.8Y4^Af+^08^^IUS=ZX>U_bHC8^
,e8.IQIZP&[3;SK;Hg0=HO_UP/^NZECX):E.ddV@6?TMJ<=P&.X8,=E:-\P,ZO)7
&K79O>1J;HA5aG;RKBJ6H)_:HcXZ)>_cH4=3eY)gF)9ZGR#G>=--,Q2\(&&60X/W
>K]N9KVI^&45\3b[C(V2T<3g0LMHU26\)R?(E+,(2664Uf@cZ^E3U&675(6GH=dM
,(9H#_)S7J#f>\\RWa2;00b_VMe5^-=9;YQa&=07bT5>I;IW9&TW#fF=JaI8W7@+
WFaQ[Db82feA_(O&Uc,Z>d7M</c?V)e>5L]H<ZL4@A(J0W\\.N?++d[dC-7:J1[(
^+fUc_)/dLL0^Y#2-E\O_505bZ4\<0Q[b^CRN)^I)3.3&d;JKNUOf,aT4gGaJURL
c^IFOYE7U+HAa]:H,&TT=GSe=N,RT7OM>fRQ4>MG466aL[D\2\F-;D=DZU?(G-MM
ce4&]Z-6NBD6:KVcD/K\O+d#5Z4?)PbLaU@9Ua#I)D)=R#0K+F3Reb244H#[R?fE
>a2T2C-V0OVcV)XNGI;Fc\\H4bPYK:@DNX=L/#HW3M#U6D4//R>8/3O/1He<2L:1
-OfUE(4Q)/beVb@B)ZY\B4</K5TQb[cd=GdFfZ-FU2R_AdP9TL=)?4W,bGE7+c4I
X(3b1b8f0KD-UOU]0#?a:gA:_9I.MA_Ve+HR\5]O]@;9QF\fQN1UKT;7B(QagZf:
BBBG<fFCSL9AIbW7\V_O8bLO=c>S-Y1gV5Me4G00/<Q>CUP#Icc#,=4XCRP4-/&H
W=Y.X//9?8/bXe=81SU:D:f6gVV\d\/C=NH>]CSdP?c@D8U,AcF;I^.NFI-S6UH;
)/Q(E.DTcSW.;^BCQ?=e0]7VD=d&5[PC(./RHeZ^JE<FRS&:<0._^eV5g4.8;Xf7
MSF.,/YMZ<9RWI\OAAS5?+A^f5SQ?3Lg]aP-a^\@;YOc3IML&&0?fWV)Z&\bC98e
4SB7I[MdS8H7aFEO^Be?)HS+WK]?.\,MVeaU(3:T=V__B7\=gZ^O4;dC^4_GU:fR
-gRZW)f_]g+TZH?YC9N:9=^6,8;\O<7+((3TDPY3-/=4bZM84OET9FNgFI09M66;
8Z\8)LgDdLEZ#b-cR@KF4.3eN3MdA:cJEgGE]W\V2RI1Ld[QH2K.IA.UO_<TLD5-
[B48_1gF_WWY7XW#>Wa/UXbYVd-22=YHS.O[#KX8B;caOQ;-0>5=,=DU/;G0B#:b
GBBXHPd:KIM;>\)7]X?;B.S<+/E9@B1Ac0U@0W5_T(?\d#LXaL&X:8Q@V>bTPFRX
;_;1>9[40Hc15OENG?cRQOEIEa8?7(S]?^ALR3J(5[1dV&H+)P>W6KBP/P-+[:87
C:Rac#<9RYTb#>^A&gOfTHMF:VcfcI?4:EL=_QO+VS6/&;R\cSRKN5&8QP^3Bb2R
7#=K9ZJfH_XT]Y6c,J0+8V9?]04#3aM?N^(a\dRT;DBb1LJ0^U)@geHZ];[=OC>F
07>@6gWeWGMF@^[YLcP7Y-cg;F723,1B82O?PWT[A&d[J/M)<M.+.MP-0=BPa-,.
<d\@SQ;RUN45aFLcX.U/_X4@3?G79[6]J@LJW/=geAYENW2XM/F-?6C+N(D/.g=W
KdX.c82U0PcLgDPW1I::cV&UBU[d[[UHNQD0R8_W&6VLB>FVB<LNL9P?]#6NcQ(9
]K:.]JRY&BGA-V;V+EIOHHTZU5LaX+^fPUMI]GC[LW#e;bCJ]I,-A2dESB)S\(;>
B64dC0+RXE^:V>F=D=^_Z7=-:2<0E3/_CAR=N=)Paca&=EMP]b6OB(]DPVf)4bLG
bMNe&6+eX3RO@JY)D1,TS6Z1dJ0[f7\\?R7Hadd9_YLaWA3e)FU0)5e\YTPF22dE
3T2U_:U:&cF6@0J-914&WMJPg1WTc)LZ)]eJ]cA2N7Z.c:^QO)2:DVc+FL<C5QSV
5(F=L&Y.If0(TP]@GM4YFIS#/P@R/ZNKA7XHTb(8ObS>KL,aV_),#0.Ddb;<-48S
D1?9E<W&S]<[Y:K#c:.-_IYgM18gff_U56M=03A/7RF1U8Z@W<XA3QA8bR?:PJfN
eFK5eeOgaR.])CDEZT<9]I3.O1)]^PVM/6?Y;H[2F(cJ@NWd6>1b>&0,X(F15\23
WVJ0WYcQ8f7G_MN5>,YFM>a[^WVcBf4#OQF()-4Y<EcJbce6(SFNCD>XdP(T:CE#
2<8ZGAXbA6+DQ9QFMdbgN)6:C\HSaAB+))VXX@1_EK330GN\Yac+6&94I8B7a?]5
H2P5H.&P5ac5>U@P)X=a:-MU-O<E3IP&9e.dK;#5Pg#L-1L;E6HZ+:LL2aOY.UXG
JLEB\/5DI><]C5&/SAUgA(,cH6LT;Y5S:G-U5T>B-EB[^#YC+R,:U(GNf+O;fM8V
<SCcg?GEXPDN:&B(K6FaH)Eg1,:(;THbG.Ya/3Ge9:T\U4M.AMGO18K6HCQ(DG1_
3G.7&d7gAX#cTbO1I4N720XeO:82W=1B,1V67\N?]/1O=17aL=H&@X.cJeOFP6-Z
PMB+=&cP)ZA4T(K\N^LE,94d+CH9^..)=:E)GZ8^BT#ZNK\c\4NJ6R?.5HZ]TC)Q
\SRV<6cMMKUV61&@C&EW7a@aN(QEN(K_40P)C#+)U<1AAD-T]O,WYZCf=CFL;Q[B
,YCP(d;T^\F<cG0QGJ3:@Q>^>X4<1UHF7,E-P8\V;)e#<g_B.gFE#(c)U-b5TY=N
U7-W-67>_^?\R9DF#44a4,Me31(/-GIY[bbO?T,5L\]#LV]QSbLWNNX9[G<)=X,<
I[KU?VP4FX\_C@@[;/XcT/7gg.Y\#/Z=KV&(6\4\CVdIQR=d(CB0eU<R0=ObU77Q
BU.F7E_>@J:L(^H/3FS292G_fdd44fYWY:0DBCGJXO:AP&eT3_4ZGf8EGWC.FWT0
a9eW^Y&UNQ5_J\/dQ.\2TgC_:C7e)EC(UA,#\.UGgcaEVUDZWgM8>7]V_Pf/YfU,
9SH_b7<528#K?)f=54cUaSO[L_[F1RA2:&\:H:=8@<SC(NEYC9X)FS;)I#:gK46e
\:L&-08LS64Y.TYRD2O4<@0.C?C;a#eSfL7\P-9:Z.=H;Y6O0MT69e)1CO?H_DG^
4P;.0?,#ZaKgK<)\;Z1EX]33DeO\_^FZ+U2QTLBKMdUZB:S+R?.R#9]GD-b0UIaQ
JbgD>;UTR/IcDW.3NRUC]4Of&-[(J2-SC:EW4GQF+?(@7:68D=V#JLP5AD1b_7NH
[+UG+C(7Y=_U6L@Q;TN+BD35W.K^IB;;YCQ_[<&cHVI>6R&:[G^b8<]#cC(;,D&X
F;eYQA^D=8M8C0YGF0eRG]O+Ed77/_FV[8QK?S(FgLQKKLVK8aa0Lf>aF4;cP9<;
=(aPW;S1Y:)bR]\.GW;Na4@RX@N(-T:3_&E=<FLEQD8KJ6J4YNWRNfQ(6XD57A+e
>19QJ;PV@OA8,MX\)bc]_:.J8g7cW)R9VH?ZTefP/HgYMN=UP/&Td=C:b+b(THAX
F):#dU(,1FDDPJ+/I;J)aP.T]J.Z2:Z6->-&9=Q,RP0)3BMIQ9798I/=<&DeYbSQ
1FAI6;]5cadYOWMaT;Rd[_N,,T45X^LSRX-HC[O0.e;1g9?CO.R6TfcC^60FeTU.
D-+,8cN)cb,F1CfYN8(]G2W;RT@Y/@M]4L19@;OKT._\<V0<ESOQX_^Hc5Y[/4H9
]XOEFD<19Y26-f28JQO?I)<95?J4C<7W=):#+0V<cdZ5Z?CNN<QR(^R,LV6b?B..
(Pc:bdb=^bQ?@@gB_L;_.MR=P^e._X;O5X/g3.NVIH7,>4<P#eWTXP_N?P<R_&c-
8RO;6c&)g+X0=G<7;g_7PTMXCJb[aK@SaX<O&?8D4K<(C(F9MJ;UGKT(cMBGJC^Z
?E3F/V>0g)&,?>XE>J<f@(BA8L=^2QE+-bd,7TQe.f\F.DT#/?LQAO[-?UX@QR5c
F\\b<&Q@I#0\fT&dRYb-+C\L^[265.?_+7\IGEMG,@a;dCN(4PY,bJMcA@:8IDNC
&[TI5/F1,gX7[QWFS468]3HF:c]Ub41;U_321B\OOb]Jb5ZEdU[OfVWc.N1KQ/5>
+NNZg9dc,4<1)/..@/:.;G2=QUU,CS:D5bDA?R=,;Q)#H)2a8=_K-+g\]NUDP]-Z
-UXD1]+J>f&XP20O=JD#NR\/&EU1/QIL)[P,MKJ&a7c,G<@gHQ/H]2N#4-\6]0f4
(@e,RMa3^DQ:DTM(43&aFfIET\Q\K.L==L-JL675(IKd(c;(-f,=[^Q:D4Y1MdI8
\[4@_H\f6SR@4JV/QA-[CHVJ6.g^B,-<A-e>94P2?#.ZBU_-+E66<PR0V=;67;M)
RZWMFf:?W,10g&E3d[NL)VF59=<;T8(#SS=21fVeC,EbOM[CF^=gK8PULM0KYSNM
4[TfKU7^bYQJG=g0YXIZO@_R>(bJ3c>Gg,>4RcY>02#@<I+Xf<G2U&<,N+[FA^Z3
;Eb;C_a,KOG,]>U67[ZC=.&@O>CCAXOg>FNE?5.C)LZSI<#W@HD+S8[+f)FK9PYN
:O2ZVS9A/RWR#508_SYA55R/CX:+KX/[=\Gaa/I6b7;XB1@GLYSa5@=SQDI2B9_[
b?=Kcg=d^(XJWHg5:+d3?Z.KA+7->RB7;C3;I._OYI1fE;R8>?Z;WWQJSWgDY0D=
(eeKS0>_L#eUV>SR<\,1=22QC252:-X\E#22JE()=2-W)B\-3,&.@@Z(XXb8g0>;
@(XGE><;+gd(,Z<_N[..08]f#R#@:bNaY5Ed+8e)?&gYDIK(YH&e<_S5?(R-OJ^9
-[9U5(^3M8HQU#)bO=W1>;cZgVM)YJ-][c<3b8K;)&cG\X4,X.:G>2e.LXA]?)PU
0f@cL[IS.H_N5+96bQ2VDWJeV<-dYI?U^f&VNb:SAe@AS&:Rb2-CWY]71#LL,_HN
QABT1f9^HOK=O@205ZSB?VJP)f-0\;ZPJ/0P@c90M7M)8CD[K-Z?D4ZbNPCbg296
A7](8#D,M2S]8QHMYCf?YEJUJa52CcCJ9\4-E&6]3dY@#>M8=T__fP2^_bfHV+-e
gK7,OHXIBK#&gYSSN@_aYBFbURQD@_:;<RW_AQ7]G#6dZG;>PTU8EZa6NUQRNF.V
T[S3NO_WZ>:PWWUU;[9K[+EV1Oebd.9+_a/T5^g2YLCg]<,TBJYD@5gNbA1g)cBC
;Vd8G3_fdQgO/G@X7cf_CCJ[FeP7Vg8&</UK=O_<-@>3OcPM:D@@+A3:aBV>4YAM
54<A^XS2a43G[.;Ig&F:fD5Qc9Z&_\bT[9bV<dLHN853CX4-EQ)Q3YIRD1_XU^M<
B)7^&XH;\N#6<@Y=SA1HP,4?C<9<27RMC#]SIE9JB_@_KL0TJYETJ[Y]:H?eEgII
=YV#@JeAM3+R+Y?8^)>bW5[O[F((aL&(3D.9L?YXUPF.dK3W,-1T&e5I.>12)8N@
^9b#aC:6\eU5#7:070+eL?2W/QO&O,3[H?.5N;J7M.B@&H_&C&4E<[?4Q4Z,EA5B
TV\K\^d3&)Ba..[[[F-^=#[(-V?2WU[Y6[8V^V&HB.:OG_O>04.;T&I&1@T4=8:#
/fU<,)Q29;(N3[70Lg^U8B65>gM_3gMB8EA^bD7gYF6?(RLQ+<@.FN]b?:UNfP_g
e.F3Fa+.YZ9Y>6Y0CU6BC5U=[TE&M)L<Be170,YSR+S^6PJ@,Ia,>GS>=[7gD_@(
\=YN+T8R7=+FRb4:QJRJ1/?bc6SDVYeWNJcW5_4_(1V.@7TLD\:[;118OccM=RNK
EgFN(21)..<5-+\2gKPQ@=L_;L@;V6D<aMS0U]>0=;=D1FQ0UQfSe?&g-05FYI2Y
6GRdbSU27c]b=NTDWL8G,>_POc=cSN)>N<c@&#@B^ZG9XXF[5)2HN7?e>VCgQT[-
75XgE]BdKM,NfM.3N63e,Z<#a,1BQ4;>]cH2[+K(a^H7\4S<dUS3=^<aU.a2,Jf]
;S_B5&@<aF?^8GgPM?8F]_bL@MUBY(UNd3g[IEG8\5<3]EZa:._@X#+OO&VYgSRg
;gM>^_]^L8[<BA([0>Ya^:fE+KYeU?GdQ4KST<>:,]4JCC1?:&QJR93GTL>#.@@4
-I>Ra]&WMRcIYeQY_abO_WI=/dLP/+ZLT7eCg[eb,9gJ[Y11L\[6a147^\cKgLbQ
YC7BH:G:QbW2bJZ2.f\]CW_.e2+SB1E=?G6/Gb9(3K_MJC^]/Ueab>-X01#]NcJH
5QUN=e@O0DH;Q7J=/3RL3Q=P/e5]JBd,+=-abc.<NI4EbQH4XO2YcY5JU/K(.>Z+
IDE:A>_@<9=DB(RX?bfgd@g.>GM>HA-0CY?/\Od=C@b9-EAb_9^0KU_0:9/@,])]
S<T@NJWFSY&:EM/UOX4dL2]3V=]SOeV]NL;N,CLXSH(9+B<H8[Oe/18UMEaE+Ub3
6Lg?7>^>J::2L5PKW8dQ65bT[BMAgGDH_)/56C=3,-J85>>f])@&=KW?5Yc.#8@3
>8HgPKXTTO7d6PMQLQa5&;G>;:EC_4ZO4_[8a&<Q0:F6UFBF.(TM@H&^aX@GFIQJ
-GaFb,Q8:8RBH?F5^=KOK/OE(XXRA^[fQH3EAB/(C7Y(98g?FL2UE73XVAJ<P)a#
YU6Z;>g/)_2[X\4ZF)+:X<4-+,G:(T5\=4?VF7=cD]^+>1dUd05JZKgT,Z)R\_b(
>M^e+(6FC654S\3;=J<W<8=&<f.KX]5.d&?B9[?4JE_RePJgNEPL7[WQKIRdXDdQ
RC79>1UH(8._bZ,=D93H5)V5SY6JfI+ZUAF4=#a]T1@bAGAg3ZXW?S9(CUBWMD>G
M?OLVcFDW:B7fL(>bNg2PXcOCX<F4@\)f/]91J[-#C3[HODBeg^WgfM(6L:-YS6U
UX\?H(#]OfcCBc+/<[NYa:P@3:\bN,QOb6[#CTQ;7^9T?JB^F;Te_:_4;T2cV6E4
/#/8;E&3JKTF_O7Wc:6e^fU9,e6g1K3=60+FO.Q5<gbA6/<@JXFA;19gbW?GJ)@1
a_M^1_CMWQ2Q?F3(M,PC+K;KaZ_YT/@Ug]L-2Q(TNC:WTCc9I@1E=Z=agK52V-.G
)f11>_Ed_e36&#6-)gA>-2(YN&BZ:9Jg)R-QdI\9P_47=6ZNC-)c4ELf?KSW>?R8
JI;cb/8I7ccHB1UM>.V]S&I/0D6g0:TV<=C(WV>@ACXOJ,<VUeW/^Z1];YWf6SEU
HPN:cB+1:D]79SLC/MD=aV]KB(Z:\3JC-0S/-BTQ^J#M3.\&&a2ULX@#-?8Hf8U.
PcZ_KJZA=&.^fd90ADO&UMZHIV]ce0QMY5R?S@(A=Z:g<XcE>#c;+E56R@(]Yg6C
+X+DG#OYf<D)GDUBUegT,+BM\_DBF-#@N[E-);P_2A;:417Z<+,\AP5/5F/Mf:Vb
@4Q1/H]6OZ7@T&M_VFH4HMMIO)G>#L+K/VFfEJ0fT)Ob5\@03X.A\3CPbU\>VSf^
9B44\K.YU2E70HE4GCd4V0f#2L9=:AKfMKH)g)\#FI0F6&7b._/YZZP<bU+YM^UE
AFLg5[8?ZWF9Vf6TB\Ka3G<&.a2Y2T>;YZ>#NM8OVaHI0GNMRU;eJ_&##GW@59#6
:OXSE4c+]JDD/&FAB4=7]\g)L>>OXV(dd6fZ]MQGe4Ld\)4.X0,E>QF-WDXEcNM-
b[G&@EEF]#DK4@3-FP\7X>]O.F2LD^BA8G>GHG2:eJS<S4:=-\QScD_OLT#0M5[_
2+7UN3YdD/)L_8M<VRVX)]c;b)=(M?d]0;O(e)Q/V/?,TVS9S)XCMO?.&-FR](/d
^CYfbD@QDB4d5@0+/,6^ObJD?2O6Z^;ULg4H;EA/<4a)b?cN+a;RL_-TfZ/KE]-e
\(<.eb6+P7baY5^AYXa0R@8:ObgE#13K-,;UZWPLfK&gA-0NN18+)BDBE&,.eMM7
+LgO[^RL)Vb_E&VH?[1S[?Fg&XDg,229[FG0Tb>H@)Q(-2]?cC?b]\F]]_@&\2VO
;YQ#(Yga+3+2;W9La(b+=VCG=V)Q)e./&[#NS;]_PJ?T+LO#_^C[8+HW-ZI9(Y1I
f1W2Q^(H2]X2R+<^A/7,N/KV<<b#=JKaJ],-c1,ZWB[733+N&>5C@4[b/D+3O.Ve
AM&UG.A-9H<M[.(HB>L\+aZ3\7FQ13/VOLH@8-VLf8T5e^,_c,FbH6fWKA.#9BH#
<0GNF9Lc,CHVD+bS>&JZZ9C?E><<-C>=e&\1HS&/I8V1(X8ZOXOP7A1M79c>?&#^
Wg.GD[[ZK,c&WJ(.a9;a9X?LB9(LAE^<Y?LP:+[2@I12M#1B1>3YFI<ZFQM<704Y
c&.&5\:eeVTW[Q4D,I?cT+F8dTaVf(cFUXLT6gAI/XVW3+/MJ@V]J2Y0N;g3TON-
7b0_,Uf,3e,L@0E&;[4+67K&+BXTOP54BD;3>P4B4L=FM<7f+:ad[eYD>7X+Y&<+
7<BQZI(9N<><JOG-Rc5_XSMX06Q\T0._\?g^R]5ML5?<WD,&DB(\,7TM2PS-7.?I
cW8b10XbJ:fbI<<?.?BKZ+#a_=T.0/#aVH/0M+_9X9g@-GXg5-S\-H<,H32_bNA+
<9Q-)E&-ScNSdR>YbR:],T7-N99P#TQd-I[[R0SDBGZQ9FB<.^)1=DS-.L\fCCdL
cf\EX^G(]C@(>8UDKY#=KG:XK/0K<W_.1Ode<,4#4\^ES5=]H-QAH29b?#5df:Gd
?BABF[NT,&-^FFcW@(9O;6AI&Rg?^^,7S4c(gNU_U)=a@4O+VTZeUY[2Q4Tc&XT:
Rgg1&.\@4Y9J7H=LRZc:-/HFWe00?H-V0,\_[658.>6PT,U(Y4^2Q4O5RR(IC\M4
OA6De=VSIgI]@:,?FfJH_U-EYdDZH78)-Q,_e84NR5D2+.D5O]fe2-JNdMR#.[8f
G\]M>#:7YaEUW;]gTE;K(U+)Y_Nb>G:<,g[RNb,/3B#^#WF1UcX0X]2/I8B97F#U
0_JACeBJVLRRCVK]8YWRbP#WSJ>3ed37V)GAMMLZeBI-cBEFA^^>W&O9>e[1b;R[
KDW[7c=168NUFd-E(X+Lb+;G0R9.&(9,0=BEF9HR4^_@/0Z4&bg,a(Db:14a>G>2
Pcc8GSTS-6)E6\+B/)-+PF;L;@A]YQe5,OUY8WG35P\adH&>@N^<]2N#17eS6:1G
;F/@999)XT@<Q+4EL;3XVKN4D9\1RI\XE4W\b5Y/O_cN-D(81N]E=[R+W/X+.4?8
dSDT,:AbOd?-Y.\-<4/#8PALGNJ?ZV#>)2]P=Kc3/^.SgHR65fJ&_:7\-9B2WPVC
L/eKP-\=,1bb?SP8.Y?QE:6;PG)8YN+<J;PWVQO8bbN<24Tg5(VcKRbW?XP].d/Q
M-4e0ADJBH_4\NJ1bLbf(:b/@>^EQD^WF]OPS>Y&1SP(^Q\)&f9RR#e7KQ;ER\[1
[=W.XW9R3fM?;-O-C+NOO1@874a?P8^^DSO7EI&0H&dTGPM>Jc^RaO80@)1,O>JF
7L/^Gd-.P^=aPCU<.]^0cLd\E&6Ad;8QHdefB)>Lf^L[BgX\K>,FX9](39]^c9UY
d^JWeMAMX8F?3UW<EF0-C_8b&V,TAfKaG&5&I^MBQ;8F;2YN3_E>:;=d[G5^O-fI
OGXg><bgH98,N^g,RbA@YSP\:OO=7R4eMCIKMg).ZOY6[RXc;L-Q0MPZ+RC;e^V2
7LJ?G7=gHL^_V69FfF2cR87O=90LAB^H&?[YGBL_GVBX.&FA?_?FT[\(0U65)M<c
dT>BPd55-I\CbFT16.]US7;MR;E:C9eQ4W:])^UQ3XQK&WPD4L69+WXIV.0IP5/b
>;;W)Ge(RKRO]M?N0OE]]a[B7DS7c@5.)NG:_Jc81Q2EagR]0^?YVNJ\NI+NJbED
B:U<4_=;R7/-/[8393E?96;(=,02FcGd][PN6)XfE:\@&(d;IM=,f\Q@BD/;\J#?
7(7PWgJg7A<N9@;0FVePAPS0fJ,6M[0S;3[bBFJ,7[X467<.AV;C^G=b7TEK_(,g
Q:<3O2\Z38ZgVDUR/?COH(30@).99gCW5V],C0=<=ZL0R6+@dHB:RAMKe[M>Ufc:
29+;A7O[>Sb/-QM/YBQ>+#+4>>_;S6e9\Z+E^6L?C,;:UC&^/4)H5a>F4IRT,eOF
)LN8UF4)b;B=VN>2SLFf0M04\DXaZf64YSVAVQeF9;^T38)Gg7J_UM(Yg+aJaZI_
(e+.M0^[\:E]V+eL02eT5ZA-[Kc&_g5#;MF.&8>[fc?\KQTeEB6(fA(G+6@4)8)c
[7,<QK7BSeXTNSCO,?d-4>&&6+;ZC2cU@,,,XOAMJ-5/f^/&[;A_:FBIF@(-8ACS
=O1gGM4[W3LBFf]Z;Jeef44+ZIM5Y7,#b5L6./X/RUGI[;(8H3,1+@\#>N(3TOR;
B[Vfd0-KKfZ25Y?A72=,FN=_;5eMGA?5PN#D2[M>4)C4SO(#;PaO3M9?=;d_1:e/
c?C2@U_/f2N5F]@:@WJN&d7#TW.T3?_S9LaA_>80]RII[b0D)TDRSIX.:Y\0Y:\W
CFV)DZ@;fGbYER43>I=[A[ATG)(_H=UBZ8R3YG8W.8KcRg,+9a0O]e1M^b-KOZF&
fe#VR_Zdg>&Y226/a^X4<XM.AU;eB2:b\GZ72QFMRR(2/\,eY:2CX.;a4[ZL1(?&
D?Q_??Zg/2g=a-ACUb;7&^-f7+1fX0gSg@eF,LU5)7D5?]UWI-8FU_Xe2\d5(]J2
-U@TPT?LdSMVU-U5UBEO1CK,a.Z;f=C4)/0P;]c,7^(HDg#@:7YU72;N;>P\ADDT
QA/WC;efHF-E68^C,OJ--]N88bY3;8GeX/K(bfY,;[d9=#Fg5([Wb6>@fLSRDWZ_
\DMNV-3GM#Y+#HV/TQJ]@GT:I&Ue<-bA4>T)ePRC0U9MI6X+(]K^R]#L9Pf+B<^J
>g3WO7.&NNbHUbaEJfGJB0XR:IARX,#0S\XP;F9_^)2SAg#1aK7[T=LKN_5STe0V
>.:IZ,Mb+GZGbO]0UMMZV<.+SFFL6_HaZ>1PXKVX+]FTb^cTH,3DN2G)6/Dd.#KS
:</6/RdB9.7#V<7LJE2?6(XED)YQ=.SN[XRQ>LPbC:O8/[0]N1#W@26QdPSGaMEd
N5dNb,K;2P+aH^H5XdbfccCdQ)=(MB<1QDY9#T&&EUW_ENLCaKT?\U=#INc0Y[a[
9)AFF2+OP\BXHXTQU,aQ\:><[=YTSZ];_Q(BeK]<)_f8Q=,E)bSSaL2>)]G;_>#>
>@(&):FUEd9Ba:F-g)7GYcW0FJ&]O_]Q+#S/#Ub3@I]Kaf>.+,IF_H)TKeeQO_M5
\\.B3_;K1A?d/0+S]\7We(dRFC<V(C[TS^/>D?4KKY6ASQC8GXTP2P7ZWKXJ;7_Y
N8A0Z,8A&D,0K8=_MW(6)3/=;PG)1VD#L7@^SM15[=]&31O-&ZgYF0=;,D&_@37]
HMXS)4B>Y8fLeZC0H3G7&AAULOe<6.];TF@X.C[(_T0W11aB90]b@@(&>?[G>+Q\
Qg&:^N^B>Y1837&W=5(#2+[8L#.?#6@e)N@f[J(2S6D]ZL5A?<P?9c#(,aPV?)P^
)GD?=&X&8,d(RMLCbY]=]B)-&a?(daU009K/bcLE8gf/O2d,NBN)99H4)53QSK?R
Pf,NFGDKW#(5;MI&1GJ:e?1092G46e+QOSO3>V8H3fJe9IYIF6??#&TLCWG<e-dQ
TIe_&;3Q&b7PDCe+QF_KEEPf)8.3]]c10OE,HHV(bf<V1]L+MbZb#=WL@_cQ83]B
D?a]D94K=eI],,NE6@</SKI__EcQ;MRFAg.P^=6<-.:bI#0gP<2XTJCCTGESf\WR
J[:eOR8])[BGJ[6RSgJYKH,FLeDDZBV1P&W-3g79?d,PBV7D=?#SL)],X46+K+2H
D(P#@cTY(VCC<[fG9=Wa5Z14)J(VG^DM\f38UUa0:YK:Tde8=]<5Q#I&Q:G(eDX^
PX<AH]K+:fRG0baI4.-#M9gfN0RbAQK4V.#a/W3Zf4Y:AfM)6FO=W.K8He9@4.7H
FXU#H>CF&^D#c1:4-(-I9E3Q[F[LT\>X]BOHFT1YZ@/A9f(OSL:\)2/,4HP(AN]B
@-fbV9ZF\X.H&I/ea-HWK[IFREQFbL6N4H6):b9HUg<Z[T<AHW^@Z68]<27<\T]Y
9QK_Reb\QKaZS)f5A0RTF=a)KXVEdaZ3S2@QfVJ=RaIAcc@\a]d.:ADM4+I_\)bB
eI:KNGIf@_2L;ZNgc?MOYg_6<S3gE/-XbM3_0GGYV,7;HE7KPZDSEM+XFZf0R:<c
U0A,S?5)d4\86J/eQd3;S=:<(/5:BL=<&DOH7@8gVVO;G$
`endprotected

`protected
/U1U&b3ggAUP\.]8AN-L#@JYFS[6@NZ--62f11c=RUH:PG;6#XdR2)U3J0<7DSSZ
L#bPAOPVW;7P/$
`endprotected

//vcs_lic_vip_protect
  `protected
1//<\0QE2C;I7S9C\gf5QO-6Z)=]C?5ICJ=\eYgH/K:F8P,P5(4U&(E0&BD-,N+2
@9Q\bVY-GUcJU-g,TAH01P?,ALJ1A3Ie;f3dYVaEI8.&#6GBPT3Q#77\LV@PMeN;
\S#Y,)9D;:=^1b\d_R:3\:V&V,Z[-U#ea;KE:]ZEHT5Z?6=1]e92bA<H21aD8<)1
=XF__gU=;6@F6.W+2Z5=TPB24R54W.-:8L,0+@IB5d6A:3;O<;@.L;;Oa(WF7FaX
RKV&BWC15ACS:.>0L?2OXWJQ019^PfbTgb)=Y#f[&MX82ZBM>79BBMR.c-YgMPX^
U9\PVY4+Y(A6]4F72,/XUJ2<1J#Ne@61(eBe00Tc/b:HbNDdKcOgFMS<B4Ze1[;6
]=J+E;.=HQ?>Q7T/3GTA22Mb^]5B(0.MCH[\4e-O>H>Z:(^S/6S6?<TA^@\JPcB@
80:Re6,(JFb=EKZ<9824N]XV[H)TU393:IdJ/ABU\FSE?J-B/]B08eB.KdMDA\66
:0a15.PB;1IbRD,;VMJd+M,e^>\,C\LFKEJ8F,SPIFOFA?fKS+8e7#K5LKD.J,78
C:)GeZ5V#YaRUTQGG/B>ECF_^BZ)eD>T21Z2R[G<AHJ[4+R)0(\<PF09,5E5Z?T_
4G1)P(L>Zc1c2\]:2eP#ERPc<d,(S,&,fUfOC=KYCP3F^;H+]3H#DY^Nb)/?:XH;
CK>fBC;./#^Cbdd4SSMRc-Y)aQUJ^&CNV;[E0SS#G4DC<eY\dLH^&DBA^4/@bdZ<
Q?=gZ9V8D7TIM3fYBBCECTMN)0JPK2RI08RM>\>8QRGN12f-+Tgg8bB-1Y)GM/XB
M1]AR-+WOd-EH/2;0&TY;g/.PUW>dcFWfJ]&H7c3L>O0b>8LJf+D@S]0CFLQ5E7&
dJaC)8b2T/PH_4.GH+L:HHV(>&f2J#Td>SOgZ?BB:1^(6-O,7N+7HT.C_WB@[MJ2
512YH(g(\H,EK#[_U6Ke\d?:)>ZF4>DAI(Q:>[fd?gL+8/6RHPb)CY77@KK5.A;D
WAQ>+F6e<@YbX+H[-J665^cA+E:GR]SZ_;D4Je?g/VQO]EIf;6;@DZcTB3WAO/.L
2fFL]7gODK6ed,<4#]F.<\.YS2cPQY8f)-MBSg.cZe7[80G-IKa&^D9]\VY)17^M
XN/;FC6_OS7>WG#K9MDH3<#WGaNgQ/^b+WaKG.U7<>gZX^[HSJ6R;KF=-e9W+];U
=WC0\6+J7Eea-bN^+46>#H<]^ULeF^5V.^LV1_0?]:fQK-]\TLRYbN#g4J_c^>c/
XG(&&+4?HcX<RCHPgQ[>_#V-,)O[7NbHJY]dP(S\G_R@,-V87.SG7YKW[XW(TA9X
^:YR8@R&8OH=7DaX8Pa/>D:O#fe^SWV91Qf^=J]IX9B(YCNSPG;EKY95UA5_@WM[
K-IJ+#f<#X2feFNN04Sg0Ed/_GIN5d<V]4J:F)<Ga6@=JU/C5;+20BA@4T,/+Z(f
L_QE9KEdK.H)PdNe-+dHBRF8:@\L;TEI):_C.6Rf.[eUfJ03FdN@S-Vb/OT&&MU7
/>[@O);V6+ULQVGOMVKKc0aJ9?aJS>UQ8_8@NQF2O,LLM>MZ+a_BUK=/]5N7NFgE
W1;NgVc9YW([6U&/>\c4[6-_H-2XF5_(fR&CYXC?,FLA(12e8,0ZXW\MdX+RW_N^
SA2.RWH>((J]>)D@:RV>?0e_NYX-\Nc(e64O5d37=O-1aZb=BR^JcYH.I(<O?10^
f.OFJ1_;E46-NN?]-)KI)\VCCb&976UWf_&[b[:B^-6WSeXe?;Ue-8W>g@7@Z7D?
eE0#?S\_C7,536[[VN=B<)gcF@,CHcK-Q5]IAAMQ^<JS.27V,2)HOB4_FO#S]PDc
CS@L?/_aPc]6V5FIEXRV[2b7X&4GW9V#=V)JSUK\,-+1gP=0&B=KGKeB>0SE:MaA
+O\GMN&J6;YOcG/(Z[N_GB5PBV>47e#I\+\a.6=,;[]I94JNRAU5C]<U>-4ANHMg
,+@68Z-7_IJT=ReCE1g\.?5[c-JaC;27,7,O&e[DeV[-<9-M)2=G.6:.DH__I)6A
XMPYe@:E.WKNM,Xd8X)deD&HMb1<SGLZAQNX[4Db9[a,M5[D/c)9/3BS486-607<
)fZ]e;K3LLQ.+4J.B_6P[S[]C[TW^d;_]3C05R\C^CS3515-08IDRa&>XMH<AZd=
OaAJ&\0J3+[Z8dB652QZ]J5U8>_</G?I(3GMM)&&A:-P7,OYCBU-<Q5VgFK(/H1/
@5RbP-#Z]S2Hd5:eH=KeQcQ</?7Z?ZC7&6ND+XS)7\YKLQK_&N.>XcR;IcW5b/J0
f:?g5?_#6-eAV-;ZG-48]07ff^_QTWABQJUG2(>aUcPB\^7U#Z,ga7E0I.g3@;()
bb[MM:#d8I;eYT7cSW=07\7fMX+93FdEJc]gg2H;QSX;Z)F1@/5D.[HS6(#]b[?<
0G;@-U@AJY)@4SU7WCLFA6c:Z-4,beDGB.HVCH\[V7[L8RXVLMN&egP5>).aN25Y
6:8W]W.EXfD_<(\ELLJ0F=>YHFOU]3-@&2S:O+\-@5QDG<4R+cefIY-Ba/bL,IO:
KA8TT1+J5HULG2)0WGTgWCM)1Q97SE/e;C/JPP7P;EL<6:&<e:ZXSU3f9KSG58HX
#@L?\SC)UV\E,Zf8TU7b:BR1&+&1[BPVUJE.SXFYS:G:3[I,3,VG(B9IQ>Pg)-GX
6)NNeOb?6)(LK&c1g,=gEVdU:UK_N27W/QL@F@&J0,XKP#cH:N2;RC_5^7(KH&LY
#AaF9J8FT6EgC(GDV2;&8<83CQ.HaR+ZYKWTf^HNF][,(gW4THW,4JWB:8WA1f]_
e?Ka[QLD.,N]=);-=VXMZ5N_gD)IK/D4/ge?E9MERgOP\DYATPbJ;,Y-9K+2,=-K
H+M<2dTS)=9=Q4JBWR<:BH]A9K&,:+_=YC7_#Aa_N6g8GUMBJ>7W03R)ZW#JE5SD
/SWY6+_8UJ8fdcF815D\5FH)T\LI;#W.S@X-2Hg?N?:NNeZ-DVIYL1<I7<JdgW_(
dAZ@;87\>.)-+05NOb36W&1?Gc4W55gSGR,OgcNL8ZOO\0^4OV+fRW\f);?4[M&c
/QW(53Y:,-A<Pf>HCA<-T9U+>#9dGf76D(EWT=(#LG\/<dK+]eVQYX8/W?bDB,.@
_Ja,)LT+=SFE[@P4J[?YgHc6N)bd>V5cU6K=-G?GD84\,,MLd\Q+fM.KX:PKOAG+
c^TR2c^>C[f5US7+6M,EALL\ZeJYRZ?^Og_\06N8AA1A;f-8[6XJPZEO//Ne:^SG
<S(^(IV]eNG5Y=OgY1T5Jb@C,\fM[IR+\LfRVf+D74;&0E=J(DUQ4Q+S8a)c@OW_
X&IBB;B4:J1_CdD35V&cTGL)/AN1aGK1V.MZ>Y&U[a@bQbI_gY58YUPbWNPf<+g1
6V7-[)M0KgY60_F)[6A3[e7Y8P1W)P]T1(#cF0=WT)=D(+Q:OKMa45Ue4<7,A80H
JBKID1>+6F@[+2A+BV&.]SS)811>&bSP##/.H.b_?7^R@P(D71T15CJTYM;>97/H
aAANd/;D1VB=XWMc)JGb1F^?a36)eD>AFVd-LJ6QR+/bEM5=I.3\3?X/M636HP)O
DT;6LNR>L+AL(=be(\.6I,CbXSOP3:@1F6LG#DR[O&FQCVFP:Y](?.VJT=B:(HP?
8f+aB6cL^9OB.W80E/C^DXNF@7(-I>YQE7A6T@UR.T6RNDdOM6YQ(1dZN[W=gYDO
,?C@:g&WX9:Z\V=eYQSU3-(g_>gR[_\0=bA0aNP,+&4@,90V>e6aO5D->?]@F5JR
B?ZQ_UJXC0QdF?Tb]8.SM]LW5SOE6M)8MQLR]8:@#D,8ZSY-2e+_9:U06@UcMB4f
TN&2\+bd_a1]A.efJ7BYS+PM3Q#g.TA3\T&VeR&-I2#Z9c>M#UDC.TVSGEGc,=Jb
#.8T_04\8C&^L.L[JIQN:ET@c\G#]cLb/.gE(bRGLB?bbd3K)A2O]FQ;YV_6].Vb
MCD^UZb9S/#?_(449.=+?M2V7Z6P=e^^:[N:Wf8Y.X@^5\SAe+(;SL.c3^7ef9\W
LOK4+#/a<OO)9&<&.;D54\e]TODYW8DSKHPL/-U#OC1X0E7UL6U<U>+N=0L5^AW=
45-dRaZT8_ZXO0[>I\8R5@;8+D)X^a>^fUb]W7]XPT9SV7;3d#Z1EZ)O@e[J)_(T
eE.a1CXf,Vd\&Z2+)cDT=a;;D&B+XN8Ff2JXY85?dQEHe9bDNfb\Q@JBg63AN.P;
c59NVDJF29Y<2FTQbadH:WN/b(0,<]C]=7T3d\N>/g^RbRO2CQ/LXULIP/#ZPf-(
;HJF,NV\H4=2UFX>f/BR[B0VW[Z,K:dD(M:>&NgO>J^;,,..HfC[aeeO:DB4c)G5
&0Dc&cZ:]?-\MbSXKfgdL2#K?.OJ+=JARWVP0f36_:C)#b4?&6Ic^fIcJ+<GZ+)V
^@IMe0NJeeC[N3:Ra?(W:]+b14D^&XU\O9SDa/4a2C3?/Z-N_Mf&ALJIAU>G]6?X
KQ.E##?X.FE4.SM1HI8/-UR]GN<>;d1/0YcS9S220+[0\?PE/N4QdNE9R3g2T#\/
5.VFAB7QOQgQJ-eQL^2YUN[O]00#;._]2O=Y3_f-CF3a.aMQ9-g9_DNC=FM1SF\/
<FeG0(D6Q._4#7;;I)7VPR:ZOXG1.I<NW[+-BVE4J4ROO1HL.daCYPMM:=YYTUdA
JW]6930g?4H3QaAgV&VXD[-b3R=II6RM\)g2-P1M9,NJ<FOa_>@GC_LaX]1D0-f-
5>WKV6R@BVgQXcgSA0FJSY5,4X],T_A4bgNIK?1,[TH]49-,=[&\(_&SYM8F:#?J
_S1X=^QcAZ]<_V,TS]4P)8#U?..<bM=MB1)HeZP/\ADX\2O)^>:,dY&N.-876&ZK
90#CbH/\:8\Q;G\QY#//=RCc:bc9b]d#0)7EA7:OKLQeC)1.\8OWbWCb07:bN/bD
DFB3R(AA\bC1\@e(O?N,KG2#&Y-((0ESTECFND+^WL0:H<;8UO9\#EKAMZ#>#B)F
7##3#VAde2&P4)FS;ZBAEG8=N.S8AfZVBF]fQ0(:/^PJVX8:GK#UE0aMFfEFV/CD
[_B>#O/.S027CP.CX+8fG,d4W#4&,4UO69eLT8Q]OMUF[I08AN?&O,6OL9Ce#P80
9]EWR&\S\_])8F,LE=)-ZeD68?_,]B)K2==D64CWc]W9[YJUc7[]^d3]2/fITKa/
M=@Z(#Pf0PNN^S^PB8\<?d16C8)bJg+:?K;NV4,d1^+<gc\@Ae1O=Y>LR)+VH<N(
fc^cTY@)\T=><cQ^>?D,-BPBU:#4@F)D/&@4Ie^>)B9afE/L()BA^QF]MW:@0Y2S
\QA;a&RFW;2=5gdBd/SQ,f6-++<,SHMg1OBP8(D1ZM1TUD2+Z;YBOZ19;#/9b<HV
NaUH?bCPW@5=^f5KP#T0ab.(+6W,(/J\bJB,]<53^A;7-Fe/.&,O8AFCWf2]97SC
</e(PK(fN3dS^IRLG4</MI,V:+]9)D_/J#eZ.O]Q[AEC^2TI,G-g;AR;0[SQTFCG
W2cO/F_Pf?,2QAT@G=(g57G7TWCR8R+(V=W(>4Q,cTTX<SPJDLPB,aICK?3Z0K[9
f+4MT_MGSB8:.b)cH3aC>.9H5.T?.d_+5);c+9/Pc/H:Q,#Og;>(II[]eZ,E/Q/&
9-7b^14,7Z?FYQ21+&D?E,LK=PKUMNY)83^Ig,?VDVD4=E3d9[=Y@@RNR]\b(\=S
U>,>MLdgJ+30:G)RFF;^d).Ie>=@Va3f+6fA#E,]A<e\GeXcO,IRU@OGU,PR68TY
LF&Q>46fH-DD/f>Wf@JGS]_IA[(;58?L>$
`endprotected

`protected
YfD>(7396:/gbeVgeE8BP:?FP)]74#ZS[(5.X,[1f6P[U\2<-OaK7)<90<YIFU&_
6/B;cNR@B2;g/$
`endprotected

//vcs_lic_vip_protect
  `protected
8]>.,Z,0I4OS,2gEU:5&RFa65.8MJQN#YaaR2BNSA91B)GJfN6[+&(?JIJPW>K.P
F#R&Yc1ef)I;:(E@I1aOE#O4[C4<#BJTQU8=HA3GF#FTT0GO?SCUK;?aIBECF<@Q
IOK:-];.=f9:S.Q[V4(E;@VM;156P-YEO_0F6g^2>aZf;.0&>-IHPZ=S+F)=#7C<
O@E,d+dP9,7UaTaZ1YQH+9^\:R51UOV?UD_<#3X]g.BJZ,KFH)<1Rg[M_),e7Q_=
Qc9<@=7L[E?cMNT,)e+ba,Z31A_7)fHQ-68(M-R^e@3=X?+af(?:ELD1ag)_eBI7
K4g9D;96a>->Q9\d<YJQX6YNc#PX8PQ68P).Y?RYG-MJ5B:.\^>DH<FeMI,[c647
@<g^SB,^-B#+6eaP[7<e#O9#EP38fINJ8@GHP1=8#GKb808B9Qb.e0H.A;]R0JP?
)c/?WV+<WE/fA0+FJ[Y=HgV+##S[4O,b;JH2WLQHAdS_,)>[98VJ(J=a4cD_G>/B
I507BX:<9;?Udc\0<aa_0_:+T\W?6OgAba#45U[<::68NbGC^#Pd__M7TVgbJd7T
3K[Fg(/__;(d#,gb6.e3.EY0?a]247>Q9D2KZ]>Ca/_#:J=/L1V+Y7)8VT\f;H)8
L+dWP:UM^++:P1fG,e^3U2H6aKU;X;+,PSXB,36XI&gRFY,eVCQ\5FCVY)]XcHHa
?-T(PPDRK<MKIKH]\L)dPT-MePS6g=T[OKT:)/?)Q<733.#5^SN_\^[K.faMK;D.
SB7V^H-W(Hc?_629M@CV)<4UaNbe\ASYDRV^-Q0/7.K.J2W=HYN#>G2QVJQ=e[^-
.>]CT;Q5C>(gb1J5bYJ<48PO^5UgY@RDK4(R&\+>ZLJK:(e>=KF0U8Lfd<DS8+c?
M,UWC<6Qf96aEQ4L-0M&9,cV.GQQ=@4,#&21]E[/J,TJ(b_PEUNb9BBQ2e;)E(_\
7S)_OEDOO.K)N5;(\?N#A9M<Qb\/^^IFF-U)+OVFXf<>,V5De_U26R2>IP+0=:RQ
I)82:P46UIX9.INNEO2J5HfOLT&MTf#H,><+NTO5H],1R,.+Y)JbJe7,+V;&AQQb
bABFPc7K>>\\IX>/BZ3[N2RNZ5.WO2,N&ZbO2@2PUW^PRP(gd6?d_KN/K3cgXdAB
3O1?U+VG3fX23S@aOORR)KQ7S9>&6G0g5LLA2A:.MHf19DUQ=B7GF>6]b4R#&ZgV
fP)6a>?X;9bW6SHQ.)X7]V>Ua(F)fA?:gANM(&bTVFMEdb]CdOH0@#f7L&B3/aUg
N9K4I.3:L[IfR.6)b8Dc7gc7N:Wd1ZHc-(#a\S4R9[95-U/XXX:32,?ed6\N@#c8
4;-RA,48BH/@>PYI.:78KNZL\=SX<S\TRLUU.0fU)3cF:^O;?Xd_fgOQgP]Y:EAS
<KCP:/W0gX01B^@YA5@&2,DJA+:7e_abf#=V0,1Z3g=U]L^K3CZ,A3A^[S84&\Mb
:;05>H#5[,aS=8U\RXW;-W(dSHF<f)&Q3;:&<797RGHVb)3.>3P=2)RSJ(ZAOA(<
:O7g&H;\OU<6D/@&gcCQZF26R7_aP6Q=\.5<5aBJ8Y6\7U]7DOZ/?M+3?D?H(:#@
CbRf2][1[U:353--)C.PZF7=<2cd>GX/=CV3YX>3&/b-VHY7-5:UE_RI>4cSgMUY
73Y@BGL[B@^:LY/VQ5O9-5?/)_HSf&cMI,-=]L3J8D8#Y,gb<43,?A;J2_+1C16b
B?d+OY;A5;[AG[V#g,)a0-b7BILK8J9:+Y61QH8X<dZUY[[J9Ef\.#+L>6DbU2&6
V+3aL5UW_EX099I95\M@fF.6=KYEgJP)D.)\@^A[3PCaA3<e.LLafR41XY=,3X4#
=&V6-F\1dE\Q>.^ce[G1R4ee8eJUG3VfL\)CGJUJ5XfI01Y2>9.CO67#9Lgf[Q8T
DX:c&E=<S,-[F860Cf2Gd(-DeX?FQK0cZ+BVAP9;+W#b:Y=2K-C3S(WSZ@/+DU&Q
d&VF/A4@;62f6>&8ZW:Nd7FZVA.PP?ZSU8EMGa4(>;)-/X<KfID:M8B:Y.#5PN/Y
J3;@#Pb[C95,LALGU?#@1:9XM:_D/=fQCb<+K+#+4bJgMNKB)M-BcWUVV/-Y+SBN
UT(RKY73K>\MVa2=a3W[CKSc350@AJ3AH?5.I\QZ0R0af1e,WPO@eXf4N_(601eI
Z_dN39B/I9b4g\F0=c>60gDFLH_FRSW\H;?Oc4>;aG)\eT4c4c85f#7#B3gCQ[ZI
PL)E&\+XX+LUL=^g)3N1=g1PdfZc@Af)FH+_R^JM4F]dX;<-dUS_]:CLJHfNT?C2
P^Y99R<9ecO22W6Q_-g7MdXQY[;?#PJAE2B-B\RH-KX8>SQWR479:GV^UXG.<PgL
@#7A?3gWd435(Kf0TEBfI[fP1VOR)5XKY7I=:7XT22fEB:RE7bE4#_d\L21@:KC[
AJA>M76fEX=UP&2PY5)CJ=fUT)QGNI8O)@/4BDN3JL#?H7/>8e:4d.fL#.AdEOB6
dT<67N=U/8ZbW&-2W<eQbDVQK..I(0)@[E92Y38[eYTd(KMAN6=;<W-]SE.M#9gU
SN8Y;EdUCdg-aMH<EJZ1<CRML1/G66gBg.bT=]Z<XQ<SC:<L)_,UO[KfM7B>1UI)
WMcbM-D[QbIG3J4/fBWYCYXSN:G6RG][0P6?U\A:(Q=4;cC9fH-Y\W(U?1(9^Z@(
Q1NZ^Y28WFG\I+VUKg+:??fcCNBUYb@+OaSC.O.:ITZ,6CeD4D>MB5Q:aGO)_g8U
#F\<9].M\d94P9XU\AK?HAaU:H)S@L;AJe_HL>IRYN094&1J2T8&BE#eba?#YKSI
+H+?W]DA96\;6Bg3gbNBc:@EKT9S:S_;0VQT?I0Q[35H]Ea3(UB[VLS5e<1dP&OG
58cC3N;[G&)BYRf+_HE)0Ha+g6g[I(9-51<1=Ug@BX\fO^380gL<A+?QXUJ;.HIf
RD-(dg88=CL]:C>5+AR,-K55Qb+W:3X6#\(dCZgT02d8eR>5/[VO)^_\0bfZdJIP
1D(S,GZf>M4K#Z&U0GLF\Jc]VE,R^7S/H[AP(S89/NfFA,g=O,d=1H]WaL1g4M>e
Q,[]WFd3<C0&:,M+Pc15H^8_)Z_@]2S3]0:0bEgAe85Ue88:QE?[43/eRc,V2J6U
I<LVF]4LaUMVY-GbN1gRdZ)_/R.c,[XH]#FGMUP2;=@1F7YQC].C;9@^J=P]1S\]
+>bDb,_9178Df4U_.\4:cC]f#gY3W\>A6dV-VZFO-D9R[d<AAV82M3J1AX7E_-48
bSc&^(,4L?=^R40U5PFK:#.M29U#[@YJ[:4E-B(50-QD1=<S-FGD<@W[/;L[PZZb
AB9S1,f:1bE0[L3RcMV=Y)ZI>4&41N+XM&V12ZC<\\YSKK<dDJ\WS5TSbMU15a10
Z#6CEH(Q^AS?OHGN.3DC+F;X<]VB4]5Z.^bFK^bOPd\c\QR&<K((X#bC-__T7PNU
_X?_b8_T7gO@5gfG5=_1CHCd:,-V<L/+FQZG0Hd[1_IQ)gA.a<FJ;-6/eY^\-e_e
((T@T\F3baPW>RcIQ7<]c7IdTa=#eVPSQZ9&:VGJ57Y^^NP[IE(T;#,?TN)B8@g=
Y1<T6C[VLEK,.[L-@/KX+E9<&Y4L>1;892:#_2JZU&KO]A]O=\cCW&P,#BXUMGBV
#^YCP)EMV8AJU/H#]CbOUBM+9@AEMfG7:&L<3>c;Jc<aS9EYe=?49ON,AG[;_\E<
d2()&fcP@9ELR=;U&]Kg),KdN(V5gZ1E4FVTEZeA8U>126.M6FZ//gBU^)+TKCGZ
\X-5;J_JaF#>3SH]g+3F/WO<e/6AZ/K(X+.LDeUf^d4>R,Zf;Sf.(9\8.Z:4YX(F
)@P:9g6C,\7Rg.DQI5,M\LJ+T5RJ=.WV,S?Z/K:B:D\>:NF1c]^3:?MRf<@/2&))
f)&:LGX+Q5Y4.E1)NgQQ#/dC,IQLgM[D1X#H+OM6aeCKCY)Y2F?/,BHT/3YaZ^d;
L.cEQ(L+9E1I_GE]3F:7T[JM.bC^?gOcR3;AF@1,X&=fNHfFE7a,D>?7G6KWUb)7
Bf>_@d:T9PN^8P5W;a\OYBY-e1(+gV34N/0N@-6)-S7S.>fT+/CV..^+8bSR=,D?
L&?:FGT=dHRVC>.VBaFcHCD9Ta]K6,YG_BbOBX]00B?6da&I5+,W[g_NOMd,A&.#
)8E#:0d/VYCOY#]Y/GS[1KK)fJYJE/F4S-DU_K,94YPaceM,_@7K7S8I+GV\3c(b
I:cZB/SF]0H1>X&;MZCODIeW8QgOV.a;H;[e\]a+3>Q5[+HDJ4:Z#5M#84:8>-bR
4_QIBT(-#0d[B9aRA:E8E(W8NDHO#bf>)1e[:1g)7P(6VF,QJ[2_FgTPA38HV01A
@70?gF?^dJ7TgG+I+EY+[0K5P4[P6bR>S6?+<?c4ffS0<=Z&X5#dW<aQ=8\MUQ,M
4\7c/S=Hb]gf)W]6FZT30;GL;EMaHB3g.56_e_=6S:dD?_7Z[MO#La_\3+I?O[Dc
CUG1SS9L._[<??Z#<N,KY4bCI]I.<(CSdG[db3,_YaTdPceDDE<J5fG?-Na_LQ(T
R?IH7Vc]#d=M.b1.ebOZG<[F?0==f,SfLXf5dca7Wa2?:[/fZ@ae]KRMQ9?HP9GZ
SQcO:,>Z.<2GID&Lga;0C\Z;X4b>)9adE]F>^T@U9]=[TeTO2Q/F2#X_5>PEXB:a
1)/+][=XV31dGZ\^29.;7?9_J@B&FQU3,.H5.\8+E&SOT=d_C+/4.E417.d;8I_3
;;0cB.JR+.^eRGB7M1:PfcF_OEX2[OEYE]+H#J50.:Q3<WI?QPZN6()MWde-K4[1
d<SBJB4&<Q#6@38S.c-^RX)(FZWW91Mb0;c3FTU@55S1a@LDL,gU2-g=M-A[B7ZR
BGCL(<b;\^#RY-1WUPN#NLLV(DB^>bbI^9f?/Z&6FgMg\.MaWQHe[:RNVL3W-g>L
=2>>J4_3-#L+3fT^<L6@eM9W)YA4M.eLg_g)36Y.&cf\EeTV3/FRIJA^G[8[=e1[
RBe2?3\;EK4#VXOTb,Y/\](;09UNR#DJ]g<fg.Ve7CB\,BXV1BTQN].>BC[7]P:O
\[99QV2SF;/f?X;+TE0A6@R1B[51P?\([6&9(_F@U4B1SWg3(@(ffG],@_Jf@PJ?
9=b0LS7DW]&6A_YZ1Qc8[.JeFBd-RU[W_fZ/](8JX73&8^5CK#.U72E>0@TMWTXf
gW[SH(>(aD0OV]d1Pgb&3e]6:g,Jb3A&(>BF/&\7VM?\)S^X_DIgB4I??8?O0B67
Vd<-4.^S5Of#f1;P/V08Mgb#@Vfg>d5))-=WY^;<_cC=P.5M9073P5:UV_XQS+4G
eAeD,O/((-;LR+L(?3RBV7B6=]A,</Y(P&B=#_,#&WJFA4_e+-C#@<;^641WKA;0
23+P)OF7)6(X\IRGHSN=c/?PQ)=DRS-FVaWL<?606@&RV;4UQ/I-6EJf@Xb?QE9N
e,L3;b)QX<ILYEPI0dH1S:87<UPM?(.e\F(AdeAb0=J6N0ZKE#3(:1/ZeR&L?(d5
^-3M/gPFNI(DE=NHd78YNX[KO1\Q]4[RU&^V89XS7HfE:ZRdM+H9V2_8S\JB^W/e
E-AJ<O]+&;b\[WW1^eR<a(84L_\U@6eI^Aa4<YY,T4\F?9c143/N^\8aVGT/ZFJY
A&@\W6IA[)F,A;JB&L2a>;.H9>HT\?GKAS4,b0,Cd09DL#_F4E:Wa,>7>C(]JXSf
D;[/]</Mf0C>KY02Qd=:5Q[f^TQLT:[Q(dN,gaY]G[/]C01RR#9Z1B2J/M<&#>W:
P)NCB/FaB]g5);HJ:CCSDP.RK3:QfDKGYB6AC7]I=,HYV_/dg1YDb5CWXKT:aP09
fH=2(d[VDLI3/]DT7?f=X30gGd+(-CC]C[d&:4;V6/&-[+3,N&7_R++R^]2+aDA>
R]O]0#9U2M^/8;?NB_S/6R;?#DCdA9S2<(@FTXB7T)9#;58Y81BJ:-ScYT3eOd^#
[]@gW42,_R&]JL2&)@5W>6N^KWZR(<^VP_<LY5c[M8df#_@cRW5#\]H]VZEE0FC2
(,Z7^E,OgFKMMgJ27JH#CbUR)T@9@HK.d3+B)W#)VbX2JMEIeFM]+/c21?EeJCE0
?@F^S@N\M,@L)c<;?J>(58#@2/Ga>a^W7P\0#;QCYbNYHfb>?X<Zb#\/\9#8\K-b
H9(eW5B#IUaIF)[gXO/H^TQ:)RF5J/dZ4+=X^S^[FQZ6L<M61E7&YJfa[K)F;>^=
^IA#5IR<W5-JMHGTGW4QZT\J4P:bZ)KaSe/8]HY\ZBE=4H7Y]SLNe@fH;V[1f3P3
G6a^5ZUO<=<8e5I2dXg.\_W@1U4(2CV?8I#J@</#=(KKJ24[K5SBE=gCNaWMc:ga
UB&fUW5>b\9IO^fg+Z0g;J&2JK<V<:e+d]BB-DOP;2W;^(MK\LT2F8?F6d-.LgDA
+H1/gHN0;<GW+0,aQ(NIV(I_Yb=NAbYN-@K_&47=GK+#a9>/9.LJO6^STB:/F_TH
@Y)F/V1I::c1aOK<]ARc?ER7F0YU>8GO2OEH33ISK?BMA^._7Y=)<PPccHB4L5Zf
SK7[UO\F0EDLVe>CDKQ6gc#7?\8<^&;-EQ(V^&]gT7H3MJ[D]aL8;)ggZe)/8G,D
45K[JY9fT2GEU;E;Ceba-Ag&0F3TN>8\5O/<=<AZB-7-WN[]c=MC5_V#FNV9R&5,
2:e8<[K3=R1-Q6c&-ZXe1._\8gP+PKX\fB[^/[JMAP4Y4d<IO,I;.8gL@\Yf-((R
g(9I73BdHEMJF3L.[23^(?Y=&c;ZdXbB]K[C97I8dSeSLBX.f4]M2D4F8Xg:e[F0
(Sa^Q#_aS+/];.DK.a<E.-S.7,1UHING,[YFA_@IPJeM<VL&/T:#YR4M>\+A829)
77;WI+WZXTW,?bKN/[S_B(\J2X8ONeMe:[<URYg?V1#2c/5L874T;>b/VN].S_cI
>PSeBIc.]F60eIX,^0S#T?0-7<a=[+]]DKa->?CF()SD[2]9NEM8<BZ@H+(B<WN3
ZbJ5c<UFWcLQWHN,Se33)AM)3:Pf;?X&(9V]&<65K,4[\-TcDd#?PCd\-D-F-<.4
APX,<SbN)Z]^?;V(O=eXOVBXJR&QN@<[=^E6f^]JM++>SVGCcXW)1.;>Y)I1+6Vb
NKR=KU>WHb>G1RQ]O)e:.4a-@&KLdIa#C]63B_?,A=F;(TJ7AYI_GRY+_4g?CJNR
;,f7d/fe2_H0#]MJWAcKKTZ>J:CDcaNF&3IZCP7+O7U3C)BWS#/6I:C,KXe:S0<e
[,\/[+=/69fDIA1:[O9S:=(MG85.:<CA_(^;\d3Y0L\7a>H:g-c&GU_4D-#:_7Q>
5G518;U7PSJ>W:4UG#J,8e_U:b:RSL7=3&(TDe;ETI(7:N1/K256^1@3M@BW[+Y>
5H2Z@Neb,+8YVaSK.?01eE\f_Z2?C,G6-D_c,IfaYCJ@KeBDE=O39#K303?RA?U5
N71gQ1K@@Gc@\B)I5\]g==W6Fe0C3bMT2YeUQG.,&[<g;_)AFLPd.4EeO>ZTER5E
aO7a-1D-2^F5Qf[OUa2N1b1/9Ld<))JAEdOUO+#^8&#]5._[I^4J\#dAI]@_3?_N
f-]>NG0J[VE/+P?8D?0VKE?\TFNd+@cP2WJ<?N2KO>\TQ>G[)?I31C/b\0703=0+
9E9[0^cS:6UQ/5,A=Ea.;U+2+J@TB<QTQF5SYS#7Y<.<XLY.J.AEc..])2fQ5Kc9
.CeT77-2J>_Hf#+Ac[L4]FCI7NDL1B=92d,JX+<K)O^YUae_F3?<?O(V5XZ^^EQK
fCV?)05=ac1FC<WTI\)5cJA.X@Z79C,c7&5WC/TYCc[VHYYW)AF-[4),BPMIK4\L
2?[DC9N5(;aL1NH\WKR4(c@1^W?M[YGWFA4#M<&I5OZ5Z#aAg^[^:S[9ae1-f;LG
9@U(S8-/?f^d^[]=gS=EcO2G>CR@.CNCFZ#NeLJ-),BeHFRAS?Z&ecSBd;Vb:S>O
=AA>9c3R^#W<DOT9(_:\^+J/51VD6]AdII4D:]f[8K4L59b>FF59?>Ra#2Za4X)F
7E1W2a0K@,F)T#^[#?]\0V_(?dQ0/]Y@)6<A:@IdN9J8#>0EP<gCDf,SBQZ2<SO]
>Uf297<e&#d10L4gF@ATeW7WM8?V1bPaK5XRCER6BTX2U?..a1PeY@>9afd?J4]6
]SC.GA1;VJ2G_Y<L#K61>V>2KaOFKYc[94X[44KR88-bAJ:,JH;;)BAA#/g66WB=
c8Z2\-7+,.TQZ=&PPK3]X,N-g_YDO727Yg1fC6>b=0EA-WD_>CGEaRL?NJR9@fZg
XM89_#VF)</KZd6@[PH+OST-ZM(P.adX_\VHOAG25#W&J:/1L7bQgBf9Y+B_7T#)
da1H[[#_H<Rb7#5J4K#6HBR<c2#A/?,<Zd)]aO#B>RI@4,P8NE?;0QH90HgP9>Zb
B9\;cId;:6HcM>G]Fe/CWG[G]<.LJ7,:2?HCJ_RP@U2J_WV].###IB?fI?f2[^+Q
8S,#eZM_QKHAUI8PF+.YXZ0:JKL(F3OVEE2Cg_CI@8O.24;]0ECW#(1@>IeUT[>G
0L_Y,)aP3e(Yg4P)g:T8c-?7_DFXZL^7F:H6>5MRGWCOSYeTgR9?7S^MEX&&LV^[
-6+V5\J9?I\aYDdeEd+VHJT2</Z)X9S8^c>d_U8W_+<&)?Ug)8^E>=B8+Y^Pe=T2
(8D@Z../[Y(=D4ML=\Ua2:CL\VIO-O3L+Y=@8-1fcd<)A_P9A;gfVePHfU+^NG2-
Z>Uf)3.?2<L5N52H]]gJI/Z_;7DF]P.#Heg.8+ZC9JDIE6D8cJUgTf?/(CJOT3Bb
;G[.RO)T3ZfgCKYdbFGVgbXZJ10216B/;<76;WEJUf0<+eD4:2P#ZU6F4fbR#I\,
Ee<c?AKOMAcW4<Za-#BgA&[+;V=[OXSP<+CLD[6FSZ-PI>,OPEKJfD>)?ebb1O<.
ccPZ^IfDZ&YP;G31J(>1fAI,H03AC6cWJI-YJB+2G]/CdNg.(KGY;aJ3=R0cf=NZ
SEZQSbD:5E1:AU3UEdD)33d^.Z:\;@=HVJ@8a-Fg@V5@?Ea.8&9).KSZ/1#]6,8/
:7PZ_>e#SVDK4IJ4]AKEaX@La?+\39^^YXC)gZP;H1]ffR=>gQdX?0]M:=#E-9DS
/[,3O16G-?\[Hg/_?K+b]Z;9BS329)e&M3UEK^@S_2PTO#VR\J_J&WJ_BYJMHPe;
XP.K90V>^5]DVW^NLAYA+f\J&I4bWM61OUfg^aSSE:(X?(D&DLBbB1a?=O-:UgIZ
1=g;LOK,GbWB1B244,<;7:W=3C6?FX=-?R77/b]B,^D6O5=#S37eZ3V9PJNVYO:A
=LOD/R@G#3S#Y7bWU5MNU.a)LT&,B<SNM^<A+C+OY9=0I#:+ag)A-a&[:PCE(H9(
S5aL/TR?.^B:V(59ZSST/548>M6UM/a9(<-D@=,ZeS0(,U9AbMgLH2Ua0SO8E@;\
PJ)e00ffA<ddd5b3fJO.^BFBe\_b&)-65e@O,f;]3R4_7F;\+CD37>A)^XB[DA6.
1(L#.)CE3)XQ&]#OXT:<A3d6M10K;VA\Ybd<(fA>N3Ob;Xe[0>:COCP3d6@#WBCN
6(ZP;W5?B2,Q^GM?1#fe;;2?b4N1:=Hg[2IBZI@<Xe?D?6N9.^PFR4E928D6GWgY
J(e5=;>\a7cL)[XVc,A<L9gD4+I>P82);2dBa>dG1CP4dGW&0LXL?O4b6T7_U=NB
H.K2BU,F90\36Ub3R>F49?aN/JZU6T0;08cJOS,f#J:8T1\?3W8(U0=+([=LR=(Q
JK)(BX)[_D.edAa+(QSW36NAb08b8d0faO)PO[RDgTdS;&@I8a]T6c941Zg2ZG,J
O3fM?EA;+Pf3,cT0K7<(=T93fRRa3?3BOKBKFT6ORcS-10&7Y#2XK_e;3FafDT+_
&CAWJW0NL&3JVE53:T@T<+E)7Df-Z_O[+dQ@3DU@(NK?=2R/SS\Of+-Y&8O]QHNO
8AK<d1D3WXA(TN\;5DgOS0GHa/_(#^SW/B)d.TK9-D@&fPc0++eUK&4(L-X>Nf=4
CL5OF>)bcSa)LBJ;[gJaFOBaPC\dPa0;YXf25E>SZQ&J2Z^T\P>5Ug#:PO4VXR\Y
a-G()QHN(\.8WLP]Z;^F17Y^X:7L2<Q<TH\M3C,EI#c6=RDOQUQ><2U2#E(6)]SN
S2FCbW.C5?BSB3XA97>:7[THFSP)<SJ_6^L.J\]c>V,SB)W70A4RJ^/MW^-NGM+3
f_:79AM]7eT6714SQHZ2F1N:=eb+bOf97VQN0b^P@?7]=\:95RB(d/HM5Q+PK-C:
.ENBD.aHfVYaA<V-0X6b7T:.4MF.K2XI@cV.WS=10<L9^Q9US2EPe_#EUUQ-4WW&
7]#B&f)64EE8;Fd;d982=B@MI>GEa\J5F:a9\9eX6&Q+HYC@dD<:TSU.g8JCI#@d
G9T2QWIcAGWV-7-ONFYZgWT\f5Fc+@D:aS.?I3&Jd(HFD(3&d3_?g#K3N(6UG>M2
SQc,]26QI[XVXg68BJ(f);fA/KH/b&aTXVG&_QYcFKOFc&Y)bQ/7[b-?9gfN_HUT
b2fM]YGD+]?&6c=#fa.W/KOgaW/#T=c><<\VFf,=RXO/H</,R;IL9TRQHE/R;YET
6.0?N4;6F0SCPK2K>##]N0O6KeXdL4Q\FL9([A<8b:+)ZHc?8=Ac2CYfNE\b9ZVL
8.AC.F01<+_RcD=N(5d1X]QH+[^(:-Q^/b9MJY_&7_LAQZ\83@,X1^e8+NY<0EC[
5^]S\Cd,FHPVUE[Ke[65Y(CfaDD1&QWQ9TM:Hg\N);;I.eIQ5\@B:3MbWO^X:T/4
;0+<],6C_-GI=R]?+#\-&[<G&dFB4_E5PIfWTW@NUJ4[H3D4XO+3>65L^MME):gT
1&S97W(P[,4J/C9(I5()eMH62GIU#7PC(;6;=FS/0\U9J.#XVNSN-I6R7-M;I/<4
5]>-Ba1T8U;E6VP-bg-RNR<7LZUKfK3(;gJ#^b,Z4S(<LC/bP09L/5\)e5Ge]X3K
/]:F/\TF9f)IYdX:BITM-fD&Gf_K:DDg?Q^cOC7..V_74)[;X4^+G\=Mede]D)\7
=OP7C=d2S,a.I)2.S4&C2=f&OK2X<VPQUG#487YBYRHSf>OJWEB/#RN:/W@<>6?I
[O]WBT0DBH(gRb0,VRZ7KTKgI;:^-)(J93[X79WEX:BNZGW:W0..eU-0<\_&f13(
3-VZ4H0c#5+NQ^4,-SV=R0KbI=ZE^GQQcOb?dCbHWf#)+S744U:GZe1;Z50:<<XN
bTKA]^/d>GeP5?Od<FJ8.AF(@fFYMU,(H7UAFZ0g=[&==V_#D+<7c[0&.^IQ]?X3
3&4+bAKJ.>3ES>gd^Ue.bWa2S;IN6<Pf1LaYM)W.<bQeVC.e6_gP=FF(9DI,fcH/
LaX0#1KL=^HA0d>e;Q9?>?.^];1N;#D5fU(__dg;U5CKNZENgEd)#B:\(aAdCKSB
=PYAQ=@R=(Jgfe.(6gU#^[1YaQYZUIJ<^&GK_SZTLKK.X5K5?>CD4-(I&CTe:F==
+-F-]/ZZU515b]7Z9P3/T=G\Df?RQ5_1Bg6](ZG3P^:#=:WeYRF&,M_:TN8Y_0cS
^E/D9f@g@^X03,P0TZP(g/6=KE#GfM2RZJeRHO>HZ-+NF:X1_(2;f(#(2-UZL)<P
N8T)d;&]a2UWbg;1-K7Ea-CW^S6=(FD]F2-P21g-ZC2<E\B8W@U[-R1U=-L:UJBD
7VQO6UfEG#ZRbTL=SSC-VLY8V5-eN0VMCQI>Y2_Ca8#W,[^YBA>=DJ=_NEZ:HVEN
+aG7H_AR\X5>M.-C,&_0V.L1d5+YC:LPb3WQNW32&R;,S7(H_7^cdRC<6]0:Va+Q
Z?&F1J:dI88)F7.cN&1)8Id9TO-c[GTGM?Ba9?+>032MQaJU+:/&Q)J\=9VR<=]E
bH1GD-R,88=2):3c1]/59DU8-+fAg@J[S<:/HXc#5\X4c5XEQbFCP1B9_ALIH^BI
>gIe11-2W[+QQZ<Xc06T2gW<LfQWZP,)@NRD;Z@>8#Q.?XD_0RHU5dg\=aMZ)U_b
eFSQXQ+[R\)g&N#[,O4>:)TaEYU01A7<820_E<CIbEQQe:MGXEf46\1Vb4(-)8:K
B&ec8JDaf2bR05P//c0V+=E=XIb&VXW[fBU1=Ndf]IJ8H5V:#;K-]cANA^I/T/X?
g7OEe;Z?/?+-5>GUSa>:b+X@H_e](,<ASOZ_U@YZ>WPM/@-35(d\ON&Y[4VaKAZ<
>\#OK3SUV)e3U;)K(gfN44=JKIb(-REbBEf@(.8Wg;&F+-/eMM]eV]?@C\3H)3N/
DXJYXVQMLAAEAQVfT73@e,B5=WA24NR]fX4-:1>fJ7>0?c&cU,7GH@-LD1-?><&+
I)g-P[W@<c6F\0T\AJQE0[)0B>36X0g)[&U(#Hb9>F:QW]5PI+N.gJBAa29OHNC[
\a+J5>VM1=-U][?>)ZRg6eb93,JJ7+,#e;R@_JO92aO;RA_c6QUIC;2W2)ELTQ?@
GU;7#ZOZ7M;07T)HOA?N3T(_P7LZB#1V]KG>Q0d6@Y5QC)ZO-4V0WTC-[:XXI1Y<
[RY7;&eR]]e(T+82W(@S7I9E,:\f^^60.8<Ga.SLY,QFMNEA6N0=:gg]4W;C?D50
4DK54e.\/TR4QUAAN,>DfHW/X(Q<\L8c67)&2L[GKY923eb:6&[OcKE_@3ON]?aP
+XT6.G_C(WN@W@WU^<C_QQ,NICM-Da42?5bI+RV,M;M>&faH2_CNaOF2.\G9OD1e
-F#-+:U^?2A]:5/2+1CcOf9S_0WDOFI,R<<&6C4E:fM#1U2742HD</1>>3S:8UNg
]dMLS\(U5Q-EF<H,0=E0/WVX9:8&,05X56W4&Q782,AB59dVNJDN#>:]^PbBJ1I;
=BIOM3F,12D?,bO,PF/FW1g7SQc(SO518G4NHR\=#(VT<\>YV>fV\PG)Ea\;<[BN
QACY&cABWK==bT(B-YXaNT;,b6@gTZMS,FdXA-aNG3IO)gX@#efN]d?\^(+50C=M
859M1Q&MZ(bU[T-(<EXYN>-HBd:].O&UVI4&4^N4Q(52M#&,MV[I))5A>9F,=_&8
_8ZFP67BRfWWUTSCfD=;K96DY;;[gK,P-EaYRDQSc<Z_VP,Sa<?2_@:+8]aHdF?8
fPET@]cZ5EA4&BFH1H(7NPVEC&L/X#9e:),/543ZPd,dCU&O28P]MMVSaB(4W6JU
WLFGPNe]DUIB/eR&?P/C6W]?0WY7614-5YAObEd34>C<TaFQbK3T(C=7YBXf[KW@
8>Ib7aA.Z(NDCI-6GL0,ZDHGB?G5^7+U9W&d7Y[d..2.#.2N/B3TT.YW#d(QR1PV
>d9S2<P,(3Y@N4Gf#>&B@>cJ4<RP&&AY#95&]YG=eS6L-fb?JQX-:M1#J<X_BQSY
d]5NVEeR^8[cOOe/5MW=)(F8gPJKRR>LSO:+]M&?YA,),U^=1-g?S;R;@#,79=AX
DXf=>A00L?OJICM5I]4#BcA00K[MGT?cUTI&@XS?aL4ND>UY8J9.A/fCV,D6)]Wc
>M(2fgMUf5d61-UDUU4Cb^S3B/J=;0,W:\[)I816=HF]U]2@1Gf49;HZQ\[4:SQ(
Oc/#]?U9WM79>#GGE?9/S8<TO35Kc@_WR)J6X3a82LL4Y#NFgK,^E:4DI5F=]MEE
#G_.#b#Ped;<,/7ZF3N?>0@EX/U;4d.<)=BK_VD6=e6.P82,#0&LJ-8IIE1?_1VE
Acc^\/c\3[b#]5Wc&-_2cQ<g=F1C87d(2TDRLR.=719fIPHXC]/86eCV)<B^W0W?
YEL02fN5=:AI_EBCTFBO.;KPCFT7PCV2J.KKfTTFg:<X-?B/(+[S:1.702S:@[1>
dK]RKZ:_9YgcME,J2HV6)gU,#WBK^,d5H#0CF36-R5_d^Wa&R=7[Y05::Mg0e5<#
[;S^,SA-^(#]Id+SGOJQ=c]T9[PK_WBB=,T-U7.S5bFNdHPU3[A0a\75)6_X4bW8
X9#U:WE;/2b@,C_<<MXV:,I_WSRL,JV(baBOVE7I9T_;W@?d)@b@FWNR6NV@YX#b
V1TJg/7I_C=+L_[2EP?@G@f1S^J86Haa,@[G?T1a[HVOSYYO67,R/[ZJbT:UM?B/
O9;+F&^\YB:.>0:KF<LFUGN]@[90#H8[92-@=I9NB@RUTTLT<R]@F[_1cOHQ_(O1
Y)#>Q-5VK5]A?#HG-Z^-Y]]YZ^X54YO>H:d6bCP>ZfbS>R26.??EB9U?^HID9bf2
,WE(8;?[DE55P70YH^BT1VBQ6>3Hf7K\\e^[/d<T1NF2.MAZ57CLP@7GDR3I/7Jb
+-90/>4d_MW_;Bc[[2:#_U<g.O=EcL)aITH1]4d;fQ=7TD3\0TZ7c3/CWQ5S/;2.
M[E,>aRO/ccF&#bdg7QW,UQ?/F:3?\]N/_JEcL[0d2Me:AL-Yb)QW4RR&(C8.;-A
^c/:E@(I2AbcB59WTaXS5NPI(Ye\:0?VH^K6KSRIVeO^#,B@W;>0>FEKKS;6P?d,
]MK=\XI9\bG4(R.>SEg<.2+@T(#?deGd>^e-2]GW8e7YU>+73N4KQB[VJWQT3R\d
IRgQaW?gA_D;V/\g##WY#2cJ+\3?U>DN?Wf16)BT)Ye_YK6.@0S102Ta9Q>V,<:_
1.aHMA8c]>0#@&<5&RV>C-)V9K;bB>MG]UCVOYgM@_=UFI]GDAW-g&^=fO#//ae;
^6V@6RGb-B6KMM-1COPERDOWL0SF)&e9J[9Z&[1O;-Y=Nb6Yd9/&b#)APB&0W?_7
EL5(WeL8KR=Q5X,?J7V+OG&E/e,<JO2^HJ/gF?M&Ag;VeL0Pd2GWT]-\LC4dC(^D
2S>,0XdW/J&b=:X0K?gbJ9JH3K3=5UJ9f>.<>BBPF5/cAf]Y6F;D2D#>g[JAY:)f
[XI7eT>08+S>-=g6Gd?3c;3XTXf[K,dHeH]V]bHcN407P\)ESWe+bfJ=N<ID)]\\
<+@d\Z@.?T\<=UH2d/IfM?^:2ZI09I>aU]:)TY\UCMS7#WFND=d[E=>S1g=+gA60
BDIS/:#:fWQ_17g?O[OFf7_Sg4:>8b\CX@<QX-JWa)X@[=d_g1D[5^D#c2f,0J0[
1dU1XFBX]fc/YDJ[d3f3K@bHX-@7=)P)JB(Zc>Re(>L:BUd983=b\K[gJ87N9CVV
B=-b@=,;1OV-5A@_/[52TWQI.4J=2#ABd6dB5bga=:?,a(:1P>3=/9XgD\W)8O.d
71ab(1SC3gZIWLd+;5)Q;Wc7VXQK0G=B9@6T78=,f^eW,[+c/1L?YB,+>60CbYc,
fETHW,e8Q]7,N?[E1d^:^.@K.f-e(R(gJ7#@@BJ_>\f2c3U>\:__^c21P4K9aYMJ
&RN3UA?TbJI)2-(@FeFfCH.4=[I+Z#)JC>@cC)U#;VfF1.eO<,IFbOcMf)J62Ie,
f#c-BS)B]D1^(@:TO2@]QQT.V&8#X&LFLb,V33,eJVQ[He9[fL<B992c58H-&EC7
KK_[EQMU?O4PeVG\DN[dOA1Z/=;-^TL&MC8[+e#@-SKI87&+)OAcIY@OU=&7=>@@
/I-bR+WOG>_+CKX&AdE38XYG-+&\<KMaY:<->.2Z@I#YX@Tg.FV>S((W_POWCZPb
JNA?-HC(M&L\7)45/8/V@^e905dJa@T,_O&21[^8(DPcUREg[8g_B,dZX;.Q/f8E
065]81Ga+DK79,Bg?Sf.]=cFITX_F+()J6SQF+(=[NfI;<7N&TJa/\S&gf.74_BU
B6FN&:89NB@<=d3(-cQ)@@<NMCY>3.A&0.Z6;J]:bC(aCZF[7YH<O&@7MC[=G?0U
](UL]=S)+U_?YP4#^J;^OI.#^:4YPYVY1e5TO9-ZIL##A,Y.72T3]>WTN_KG-PB+
Egg#X#fG9CY^[,6X/URf9?]@UHc?UX]D4aO^9X[b7-6Ic#V;50JfXZ3H/,d8>L]Y
R2XT0Z_>)3)+(WSBg^V.d3=APaC9gU2@\#J/SIM[D,[T1caT&cNCMN32KB79<\D7
BMRG;ZMd;f8+25-Z\FRbFW9;f/-P7<_[WJ8bY(4:HI<SQ&^+T(W5c(KZ/UeZBJcV
Aee9ceKZQHML4aPRT:IOV2.0c8_X?CgW2X[KWf((D.a1,V&M;.b?#aU_?g03TS>8
8#32C-:/dSW5U;JR,V(DZWG_/D(N)M[VEX_;U3V,.H2\;43@:UY5Fb^c/N70SSJc
XSL,M+9&>5d.a]-^0,UHH^LC99/<)Q;#./DFReeHe__;b&Kg>b(/OIR?:O[C;=&^
DB2C;&SV?H(8/@G+T5Ga7&H)RaZS/DD-SGL9>H&\dBcYda7UEC7ZcfS3fa(37KR)
9Y^dJ^R4^GPM>daBC2^e#Z#;g,K.>0Qd?570>M@OVc-.;2HQDfGH>&HTP=@BG=@Q
QEMW-V;G:a8dOYWKYBT#[dJQZRaNB,aU&U1&8]6O9(71&dTXTMSNT,P6]@LbJ:B>
/Rd+Q]<cZ9].])]/R=L<-Z)M)SXb_#33?9Y@7bRe3&1/+6\[R^I9A5Wg2cYcLG=e
EXJe<eVD-6^W@S7=aQTB>cO/I6R;9g^O8VQ1A701\H]ES6gI8V(0aK5<IJ^2bU5#
ZdF_TX2&1)Ff,(SET6[1RA&]234Tc(XIO043b5CaNR^W+?cT;&2;^;HNW^3@CAQ<
/8Yf<b-_MY18^->+DGC]N)gE-g-8Y&6SI.KQ&7N2Lf^BDS.NXa)Db1ZO;OJN1J9?
:21SUbHFL<AF:deND.FO;7ITg)./D1]S,bga@-0]:91/>=a,&1L\V.6cafA80?PR
NRWKc1D\dG<17G0b5XUd5W=.0ILWW>L5B7V2?^2_9J3]?TO70f0M7O=<7,K;]Z-R
(P7f9^1c,D0N.A5IJ5CGag)dO[I8JWX;+<TM:@\7g#U1[a&O+[Z62&+O3)EEbWQ@
?5g9]:EJY6,M=<-J^AP2Q=/H<^:fY/bcGU4H/IeDUGZ?\-X,=3dRQH+c5L\(B&V3
_b(WP7^ZPEYgL8HXG;AOLI[2BP-0N+F+Xcf[B6LdgX?ROJJC#:Y.AM/7\#COb,E=
+dLD(ZII[6\EVA)&R(I@3aJZ[Gc?3^Qf7UGX5PPg#6P85O[,IQS-7A>+BVO8TY&4
Vc#S:-,2aUKCF?eV)Lf8/\E:7TK<[17YT&VGGb4fbaX<D:4eEBO,I]KQN[ZLe#=R
[30YV[TaC@<g;:KP8YXC#fMQ4=,Db-#aNaN=+@]fI6-5268/\J\Z,OB(WV89ULf\
HJA3NJRV8,E^LLgbD\CXCH12\H-8Q<=^?,^KA4[fT=O?Q][e@<_6c]4@M]C3VdI.
FPFgd\3cCQ#e3Ug-8[CTO:P4/a]B\?&:6XT]a+LTL6QP;VA2c>8=S=8g#3aLO7C,
52(G=E6@?>,fR>/?2+7cHG7fTEO?)>Fc/Kb_:S@HK)^R^T>OHSE9&>;Z;2KCA))_
KLFaL@\?,L@41@U<PRNZ63U2@ND3gARWFP6+OAW^6=V2-#D8((Q[K1H&=8bPQ)FY
A?KW6@^@=BV\W46X</,NY)&YV9X)Q#](^1XR>0>YV_IYV24AM?^+.:P+8G<:+2F-
(VQD7g0b8QD-7^29LXc6^E4[#e-CBT4XMELc-FNbdG92<,d?W?W47/CEH_UDV^5R
d+-_f][#\A7KB3_(3]&G&9X7cO9N8B\/8AWNC:b=cb[>dH28B1,ZXMa=fG&?2;P\
XTaBIW1D4ZQ7H:;X<J-T\=(Z+MY2V:=XME^0.dIOF]Q^+1dZ#J+ALHUd8ODJcO5:
JWP4-aI8b9S4+(PW])5b3e=V69ZWEdL,2/Z]R?\(ICJZg)Sb)K9-:U6gH>be/b<.
#B@b0(R&]WR_^a1+VC4\<XcAV,MPfR<Ne.D/FA^YGbYfZg/IZ]C?S:@YaD<U<3&O
YXa&5KEc@a\R5)/JM.YVY.=A;;^2SADXe;:?)<PRd;\V8bQ1b;R@4&(U-e,,Ofd#
0f=#-W3W7)4,3#dV6A)ecD.999BQ6-OcX)aL-TCTQ,RAT_UYa\Z4=gb/J[b8e,.7
b4#/d\YR(\DHE]G_W5OD6I]QeB6C:H^4](eI<R;L?V9O/E_BMXM2U/-HEYM>B2#f
M)fT((KY_70Hg1;3dSXG+e+Z>_.TV(8NU]SA\-MN&N1<G12.OJVWLD(E>]:/9&HV
_IG)FC?e^EQ7?-D)ZgNJ[?W,I@AaWeMCeQ_\N1U/=YB9SB[R)C(9#R[MF^Xg6MG1
?CYQFC(JAW+]CW-U)CEMX3b9YD?_EGCN-IVK6F,28L2c:V=9K:9?];cG+E:S,44J
Maa>E(PA_#&XM_[Sc-c(3dB=IDHW9E#B#&FQ@PDb#G9ZN]I1fCL@>V@BKb\Ef>+3
QYR]gYObEB7WL5dULY>&5>C-98\<JF6O?YL5T?KD04JZBOG(6XfF.e/U^K-AQfY:
#7D]4C=K#.Q9aP:_f67-^[T;O0GTN6CCH]g0C1YT/BMbYacEA[gS7+7a(HeG5J<<
AQXcVW3>XQ,HeI&BJcPfSV34V.X]HA/cHO,f8J0K\d7A\33b2RMUBO7-;223&N6e
]dSY4dSd@U@gIQ(G=gJ+.:6bdU-5MD\^TZ:DQ29G>_X]>)Y-+@Y--.M5S71d4U-1
^U@:9BS1][3KdB+I..P7,Cb6;>&Id2_DUN@XB]=BZQ4fSdGPfY#QP8PcWRH.)B,J
,/C(\U4&C?ON?X5KSP+eKXU,7de(MI\9?2,c;<QQS09]#0aIG/@M-0;6Q4]9=?RC
TR\FI,F:ND84&.M3RY),8g:UXE63O8H<81#fTME[04ZQPQB;WYgd[F),_Y0XV^OE
PM2S9:0ND>eWGG15aP_gMZ<;:ca<ZW7Wa>9gF/R;dAXL^HA=0NY,Z5&K4:HKNfLW
aUT_9AcCPg#K>7\@:7_-+49(ZEKQSGeQ(OW^HG;<AQZ(L?+@V-B_6+99g9OH2><4
9=bfHFL\-?IGL(./#11:e>(./R__HPGLWeGfP<,_NG^K<\SZ?5]T-8F7\><J=gYY
aIa>0FVF6HOC)GOX\fQO<R8g]T-;d=[6N/:,IFN5\7L_>IJI2?_&f((dI24]95J?
HPIU\O-OA-]NQ4dcUF@@U7c>X\AXW0bXC(;FO3W.aJQ#]8fVY2C/a@EPZN#^=.FU
GM0/O;;=c.:35Of<L9=1bbN@[SK7F6&g:H].,__c#KQf]C9cgUdXSRM6(NQG&T4Q
fGB-K-Y>454GEaFgJ1HdTB(&YG>VLN@;BZR)I:Y@Fad&9SZ;OZ/BRQ@dgFaO=^GH
+A>0LVAd_?A/YN4(d_b_3@.g.@^8EQ1cRUJS+XVZ>I(@2E<c5[891\V[>TO?Nb-L
0,7AR^24fMM[09F>PDFA\6#S]>4:;\+agHJ4g6Eg2d1VS+F0^-985I8\5#<X+>,F
\LXFcL.?M&US>PILN<YT<c#ILf01D#,7HX5V66KZ0L)]@Hde,3U=cZdU[V7A>Ef(
7\Zc>8F;FNRO;C)G>BPZMP;3T-a_A/[0VRTIJ\-:;FfA3E1I[7[&[#<Z?)<DK(-H
4;GB5b2bCKb^OC].[VOS#_1;gU#9a6O_)[,dP9GIOPI4MH>R8PIE,8ab[\Ke)+37
C_(I:[bDP5B1ZW]PAJDL0RFd.Q4PgFg+9DffVY>GV@>K]BK7CWENfW)<ZfQ.^-YY
(-1b^-#WSBA/]96;V>^J[&ESe/b2#6J)+@KV&H2OA?1W=OdD/6RF3DP[1>3;]AI:
>Zd67H0a9GO9-LUbMd[YZ/FV^(\RPa3)1fB[LZ-+2e<7aZVRTK^I-J7R?6-ad_cE
CH6H?/I)fXK@A0a2]6?)RDA,IE/C7.fA96G<g==W=>T/2dL+B5c]+#72WZLVUf.>
42+S28X[.GGB1Q^\:E:.3C9\34^eGE5V99U#:=aV[aa:1/7AL&Y1Q+GgG7febC_9
B@U+<-V?9S1S^\^>REfeWXH#]G?\#?=8dT;80<J.:MD0@_E5_EOPR5@EN+KVAE:g
3eFO@7-HOe\^_1Lc18R=/.+JU<XF-T,N([)^R6-3LLRJ,2gc[466Z.SJ1?.<=?f/
IgAJ8T8=?_5Pa0Bf)?-L(X=7,ARWT&^\a/?eTQYNSFTY+IfbM<G)Xd7N&Jb72K@Y
-T6L-Ic<1+BMX9LO66\N:+O2gbf@SS,BZL?<Nd0f/;>g#GbA6,M?D&.E?cSYDdN3
<+eQG5Ub<d&XE,e4FW)OdT<7A7^7E:CR3Kb847R+B-0;]#+,BETF30I#_QG^4?F]
_&XVLGA+,ICV5;@NP-(KL^5cV>W9CN9d4Ad+0>H\YbC=?[#H;M4PWS0bAS]6Eb64
?cgUY@JeHS2YNCJbV:Z.c=?IK)HNOH0=Ag\&^g^NCHPX6(^Ua0F[QM+9fgg2dQe=
QYdHPf:8\1ABg.QfYD_-4YH(UH[=9)CEF0,CXJ9X\WZ2=Uc;AVHg.LbBeeGCfXPA
KGXHHTW;;N1<>d)?=fI(=-VN3CUbBM6=(W,?:)RM/HD.Q3?_bHW)]d]=.5JK41:6
NRE8Wb&JI+OBa-3VQ99V084)1I9G?S_;[BRcJ3B&8\^0NB3b6fAUEc)3\4O&;?FJ
F;C]YKC+0Q?RE5\V0?Q+T<2fIU65X5UO4VG=a_A&S(;7,)dT)S9[SP7aaNWHTJ6e
Y#@YN1T\7bcH[U.0bV]HXJ(BT5_1&gAER=R#FUV_bI-C_CHUEP[c]V@=9L:7:VT\
f?=?(d:.2>e_C?B=[f@V5M++=;1X80O;^AFNK+(2S(Ng[c5H;R?8>>I;>5SLOd>:
^3WP^IV(IK4G4Q1<eEUc9>(&&I?I-Q)Y^c]0gXJ>O&G06.L>ZIK0(]]Da0@[d=MZ
X,0-;C0JfJIN@A6gHH(c/1eIXb.5dTNe,=dZ)&V8&0e1M+PbTG9F/g23a\N_:2Lg
8,P\R(e=M=CJcC\(@UIa_T8Rg8cFC(K>3dd(?dLPBJHQ2)]5KCBH-TYKTZ&([D;B
fQ#D.&gI_L<2Z&V(N#K(=f7GBd3b.[d5,Q@BG3QYba79TV1fF1UYaW?J>02&8O[,
=8;[fdV_--,_F>d365>1(KTXZHO-JeecdAG&EIdQ,VL6GeZ]@07=P>^Z(K#KXA-X
)9b=BXOdM^R;2^+]XU8V&84cfK8)29:17H0NG0A&1)V<MNK+AN1[@I,/F=]\:0KF
=1T4gNC]2CD]8QRZR#;O\c\dH4TL#3^8e>SWgce?I4C\U;5\SI,a17>?KW]+DbVZ
=3&BaG4AW1_/(KB_I&+S;^8:=F+9NZBM,e7>X<&OW=&96S#)f#[TRU;f&TQP25=\
#bDK&&&bP6/E(?U[Kg)E,g=-)._#)0==LIXV6H05PD87]+)F#-+cI05R&3bZ,=U7
YF;K1RM3aZU\>^JeO>A>\:EN.&KX)G&--_ce+@C.&\[5L^1S+(>JS:RTURKH=X+B
8aLM@#HdY_)Y>gR3LHa13?f7O\O&gJgU0?I535Q2V@a,A6g\]^>g<f:F9K_c^W9.
.a:XD4_4acB-R3/4KAD7A(3@aO:D1/WA_dc4?(</d.T4_-&E^\3-4W>VBB0K@9;N
I-@5E5R<_DQT(?Ke9/=;/[d&?BgDgGG_\EfbV9WZ/NDY>GdDZbMT8QYabY&8.fd>
-=FR&Y9[IS9<94EQ@6XB.J]I;FeA1RR@K3FAY#ba2LPWOK7DWOS1K_]6E85Y<D_P
BFCQb@32BGBZ:ZIHBe1OPA-T=U\K4)Y<Ag+/8LbQ.UL?^O)@=3VQV);YIKW>SSM3
#3+4\bWUN\Z3?OFa:&MF,Z(HG5a[P.1Q\K.CSQQ.cd?eeLUYLaFa2K?/[5YCA3PY
1OSPeK1+M+ad;+\P)BgJZaIVH_567?ZB8e,_##;-DTORI(ZC>_8/L4Ra.B:NP7fP
b5)[DHXE5c(9GC3/U_^Y+:-NdcdD.LD;/PbL[W1^K/(e3/XIb_52aNS9P#K6A,W9
+)R@CZec\#ZYBVC9dB#UA(TLM@1C\H4D4H1a@3MR#V\[UUHR5VP;e+Hf,dGWE,FO
BfB1GWV(bL4>,bK+,W&Rg<,5Xa>V,E(bM?gQ(XB+/2V+MA(QXF0E@AU3(?=+aO5d
RK7[+]T9-36@-:5#4f2^gE7[E8JagB6dJAD(FMF9\S5N56JV=(9Y81REe[N>SaL.
]4-cR.(;B;g<Y2XDRQ/dFe>+d<X1\C/g^@:WeTSD[^X;TPSHbV#GSHTX+D(be5V3
OD(B=EZ8+3C4M+a3RI^T:N55Z(\:(89DGYS-[ZZ508UNSH<<M(2]Z[RMU(J8MEA.
Rf/+#6XeF@_,LY.eaN=?H[9B9[N#-GdG;S8c;0I>D[1a4+I;A,4bNeUXXQ#US<d<
QA,;_bcUB+KbGB4)T=\]45>[CgJ(0-HNEL3H7@^V4&<_VZ&>+;67eeB0_PYc@BcP
S(N+6a6L>>@H^<?VD+EVdbJPg7-B8#Q#OGZ-)b<AAfG4NDJ68-M]]CE].,K6Q)_S
[=\&+NLVMF4ZTP#4HU;CZ1<AV(>[?b5?cX.,8_<g+^Ca8CU_+/9EXZ-+b#5F)5f]
(DBK+L[\6-5+E&L>gc&8=67e_B?Re[Q?U2.-GLEP#SOH&2LWBa>Z41,/XNC^#6>I
NA#^Cb4_Q0UVX;-ZK[ATFI+YLe&DW/C0-[VMZDdbdP4;RJ?REaATc#^3T2A/R7>K
8M38GD[O9]7dgP0A8BR=\2]YgDO/;N-UHd/.a\&c&=&c[<9VE?VG7X+4N6>S1/,\
43PFcf>aGRC_?c1W5fVW&RZ;W];+<(4/;AY\PV/<XC7<RTF#T-_0]H^D<,NRD(9]
#Mbd\YgYRQgReGLf5R89ADF&gdITN>IgQG^+:CL/AgZG:CGR3.d1/b8[]?4d]T3O
)0]>O628T\HaHda8F<c0c^T0_I]),O_fN_W<^1Nae3J=X1a15M85S1edD2T6]#Sd
5C<#W4=ga/>.H(V0#F<gRI\:U-[PI7@I-WW42>HH\7b3=QP\S/Y\@Ac4:L70ZQQO
ZO7e&ARKG9U^:ff2J8+_B?)4WZ1Oa9HN)Hge36WUOg-,[XU):S3&eSNK=>#;LcYB
34:;fL;:US9,K/DV;9:2FJO69(8CeggTS-DS7N_C[LQ90V)S:BR3aP^UU#JYOF\I
M8P9bP)MBdF1:3>.XQ;],85MGL7IA#g7K^Ca>E(dEabGX3^Ff#J71XOTMY<ffK#\
JbZJRL9,#g7[ZA1?eZNbU)#F20464K&&eZNTPGI3=YO]NfTA99G?\V#]SHZfZ-@5
0g@aM1[MJ#B;Y5/OT:-aTXD9[IW9OTa6@O34__Bc=4/PfNKfIF3E5E.b^2Fe&R->
YPg[8FV>/#Z8d7IY:)QVJ=?NIMW.eI<[>L55:0;TcST/0G4(5))DL>?B+eOgaYHA
N8)9L(=a;X/G[M(;aTZ[H](IA8OM;&E_CE4aZ]-FGJ1>H:O1&b/<7c5]SEXTg3?G
K_3,[J@;e^UeB-Sf<3#g[fbCSfTS58=<E=5^.@B3aQTB1L5Qd^7B1_43d7A3L)D8
X:KP7X3QVBMDQfZ)QF=UMT;7X;[C>9H#YTU2ZR6R9>&]=3a^6gfED#?W8^bQ6(;H
ccZYZHOJ0>QVDNQLN7I]IDEP?-H=PU-=6N=PA2A4[<,,6@S>cRG6,C^#\,E.[3T>
?B3J5A0eU5cTcgRc(MB/Q/UWDHQAOE3?(P.R3c(Z01a?b>ZXH=SWQ],(&?IX#PK&
c\,?7/+bT9_IJ)SGY28=WJ]c-88O:TZ:B\#AO\(XL2>Fg81.8-,+,#8O(\:2EJGO
@F2M#eA@B(:]I6LSTPFQ.;Y#,KU63Z=][gcE1#I>?J/45Sg04<FOJRRf\M__gI;g
=U=GDM@4WfC:#d&2Q#Ld(CYaa,Y\35[[<\DB@;/A\[Y@VCMF4;T[AU1=:><Q/S:e
0P79)8>-LWcYGKMD]SgB\2C0e^@bT1N;5EQV<Xc49^P6aA,BQbMW\LT@7T=9Mf8@
<.[RdFEdB/R73O:1X)<6::5a2HK6d,D4_#:N@0=,KN2JLQU_Ug<G+fRX>>2I4=G+
VJV+=ggL=0:6Td\#XBb[AFD?-_Hb:HENLK=AUB(N2bO03dS3eLK/YZHU:39CU\]J
JQ8dQ\Yd9MV<ZDC1>1b:/8<36[EB\GHM#ARQHT01&DeMfOGeN:M\0T8HY;eO3,-A
6acJS80IFN7b])0L?2+?PQ^2[5U@W?HF#Q7efU0e-6C,d)c<)gg=@T[5bZOSM[8(
A)G4NdNSa_.)LKga^-Se..,Xb\_(^4f<]V8T^D+NJ=1[]cJf2SKQ@<VbZL0DeGcJ
&PZSMXg)4:&?REd37agf6QB56-8B_Ib>L-(-XO;087.P:,gAN3B,@6)0gPMGD\CP
gf[JO3e3)L7\FRdZ1C#00DB2^&IEd?[,;.WFYOTRZ/A]Ga,1,FR.G#IK7M-g0T&Z
bWM38K)+\9>^?3F>;4E&U>E)AJP1WF3aL20Y8e6N>Kc?:=?[8(GPB@/(_&[eH-K3
G-0\Q.f;_P^9#X0?N3EOOCJS_2Y=D&PX^HC&W@U01#1g1XQ?e@=J+1MZJJ.LK?HQ
eefc6#Gc1,\6YF]3VJaBMFZ4^H3A4b)=;VUE+OR.VEJXJ&2JeeX4\YJB5847Pa0M
K?Rcfa-5CeI4da=_T]JJ52PgXG?Q-+dCU#aL#/b=,EMXY)&_&Wa(:LWLAW>d-])S
?Z)SAGD1VK8]05G<aeQJV&Z/ZDZ&XQ@#H]fY0D0:^<_49@51[Z[MVU^EeDd:b-)G
J6_MXOaAZ?[?RGeZ<F=9ZO6PR?bdBLU/DTETfP^W4B@\:Q3P/6f_-BdHN._C-KJ\
0f2g[BWHaZbECPXMc:7(dcLFBLXd?E.MO-NT)beT=B4T&/fa1XP3XJN+H^1bNCD-
0:[\C6;f_S^Ga+19@7@];Eg<G3JCB[(ORUW_bY1>309BNN:\((ND69H[@:aQ_R1<
>8^<1F8=_W?gc-=Y9N)>=Q<O)C15Ad(T0L_JNFP[E@bYBX?N0g_I[BZcQ;eU4dK?
IcPOJ):a0@Lb&&[Y>P/^KI[dYdP-0:e9LY<A=.SGAa[g?[33b[8_;R0/#]YP+XI<
ZfW^T4O?OPUE#2g[D8/TfU>I#^(/MM8_+?d:7F\W-VS2a6#ff=@/2H\5Le(?PM_P
ZD?A@(Wa=C58/-)==EH&8V?]]\#=&5]9M4,)G4DA@.)3Z>;@ZP&)>G+dIQ^5Nc/f
fX&^.I[P&=4B(I9KM71+J4DHHEc+afe0G1C/5=(+4A-V>F,KXI^)?E+ZIXWdPDgB
5[^g4=_7YZSR2EKIF(L2gc/;J/:b4bW,?\GKKI0;62/;R31:@\R?.>cN6-O)/Y-G
V^&eOff_^-.b9;J(@,6c^IV&e(ge0)HfgU06>IU,K7.+dM[X(@CZG7cA-7==OMUC
?.d,:SU71bg-aTa\(d4b:R+9QMS48,]IHEB+CcK9c_-D\ga_GeVYd<WCG_9f=fS+
g;)KPB(HbZ#-2&1;N,;YfRBZV7]WZfV=edY;A<+HQ1NfR\bN?=#:Cc:>eWQd<;7g
28cGVO>]ge+E&?DBZ>:G@@L<A#fX\>fI,2B-f<5HEVG1PJ&Z0U16/S@9JZO2/1^<
G/;>7g9cg,^FM(F[(J][1M/LU3#04]\bd]#E7L9DNG3>W=dc&Ed+c_;&g,\IGJRO
L4;aJR]]3^B[XJUbK4gDQT#M^V#gbUa7_7H)9BXDgecZIG8g::^E<-2cQ/g6XT5_
:L9C+W8P_(9B1ISZEXIPTb>FM;bD<K2(CWY.c<bP-@e2f;F>=:&)BT0>EB_3CIDT
@TMHg<YCIJ^PgJBB45/YCb/MB&.aC@.cdgH6)0:P.DdH[b=b>0cfO^ZGVB+<Q1>2
_QUUL(-We76A?<&\ddG]d_XXd7C=SQd_G@TR&/T<3P6#?BMM)gPG+5f+K5_Ze80P
N(J2,QaR>I7-E[IG]f<#C7H6KT3Tf1(.Y@VTKR/caBX;EZCG5?TC769A;T?eQ1Kc
P=e2+F5>[PS3HPY);1WN32b1+X/8f,8SU3Z?g+:g4^(O):S>689+W99[;8]+T?Y:
-ac^LF=&)K3=UE;&(^Uc/fGL/8??Nbd8:)OOHgcedaVQ45\#Y#SQSZPeW-[O7MZ^
UU8JA?/2c9(YcJGQ;LFST.CW<e)ZcH>)XeVY3I+]2R3R;^>MXZ9:dN=:RT((<</A
dM95DFe3L?7Se3[/+<da04_UZ-S)FG8d<TTF3AX[PXQ5E_Kd17:^Gae+,HKT;(g7
O#\Y8?QfTL(93(AMF_OLNa,O-0[DX_6c9QPJ3<bQ3dS<TIBM5;f1@[Se/#I-)I\c
OJ1Hg5-G..WG4LG-M^=PT/UG\K:L(U,_Pf_C[92M4+;5T>()NJfY=706(I>V?1)N
FID#eYfF=f7@H:;CQNedTf^6Haf@ZD60GK=U/@:2\>RI9CJYfIB@O;82PFSgHT6O
<Ya>U9[>&Y8O3V&JF7C?/M\L(Sf]]0<+LO.07/g?X)&,PA5>]b^W7(SX=\Kb7=bR
0[E(/c2/6H6VGG?XYSP<9CG7B#B^RF;(Z@P9)G[R#]KLJ#8<J\RPb5Oe<:gR8L+O
]-MBcPg[6_,DN182L]fTA>EGC&J>3c,OX>>,YTWBKTU8[3A.,99F8FXWRA3V1]P5
=M>20aFF7GgZfP-UCKTfJd@J&&d8W3ZPJ4e)V#]G_>//>1>/QX>6J9);10Qc_5.J
N7Z((^IH^DbaY?8CagRfg>Ceb)Bc&]_>(WF7,.bC+E@Wb9(G/2B>#J,=KCR:UFU,
.#/TdPYY)Q2T3CK9,fIcZ6H&84(@N>>3WB?/RQ)&ccEH\P,+7:^7+G5,Da(2/b34
A6O@6LKTFS+=F?]F&30PKdR+5L)Q7AK;123./;,<F,C>-\LN7EAMRRBH.Ra5;;5I
(=]:C[c64.e(BYf0SUAS2K^D\=L7?:ZbQ6gRO#9Q1/D4^BcMQF;b]FQf:f>=ZQ@<
-6.1C0L^BK^4X]^DeeB#G6c<23PQ]>)]SU7JO.)I7;2_RI5ADJ[03WF7W(MgLNH_
dH2Q,cdF7e@IP.0P.,/F-AS+3FRFafA-d_V:BWdC(C/.94_1UWX]g5I1[P529Jb8
8Q@<5+FQ0PG=Ugc9g;>ZR)Y2(;gY=[=aG+O1-MD1_5NV164[G^_aE_?&KcL)0/;V
D.WMLG)eD.1>Q.C^)S9>WOWM/I^gV?B:A3@NDW1O]D-caU&>TKJ+fZ7f+-_@X^cR
XQJ8WDS^V\;C:H/B\/;,fFaf-ZbIQ=BMPG-V_^R9;I@VLJS6dAY=W4NR6HJ;9/OU
)6C/c9DN:T&T_&<5XC(R=@A>JL4>O4^E1;>@<Xg+-V8cb@OKT0<B,40B9^MKZIV6
Vd9S3WgCNMf+K3LUBKQ-=7+TVTI\EG;\&#-cEFJ(P38e7]#e5BRXTK)QdCO-2H/Y
RI^L^:8&Q;1[a:CW1-A?,Y+KS-(A9-STfB+&J&TeT>CM/Q:\6)3W#S:GJeU:(2BQ
A&BfNHEW^@?BI)&\VfHbWD#EJ@MJ:>GVB\6a0ga.=DL+GCG-)LOCYA<LMa3JL+Z\
RD.b/+CP_^@7>g&Z0&C#9d_;cW?^Uf;:XS1e.(M)]1.g)<X4(^J)]a8=)89K5)&,
>,E6;1U>A].:YAR0UU;#MG-+/K)G/fT128&C:OaKgHDQ>6bd:D?8N,aXa3NMC)2J
<M@-3(5X,R@LR\3GA:aYAf;,Na-FNKGGdCDQcH+QX-YU,;SI=>>Nc6@1S[6L^ER<
;f,-TG3^E^RW=NW\)7B;BI>=]97O9(&(N>2B:57TagE@E-FC&(^0IdWDKfKUX-fV
SO1[OT&F4\=1/[aCG:L\[H=E32ZY^8\f-5S5>bRY+OVDB]aAH;PIXQbRNW.@H:JA
,12KNIS1J&@bd,[>UO#R7P7U9]PS5?JV;09_(NKg(B9IZAN/Ha^WU7U@4Z<=[SH)
JCAgg6V=Jb90==.76e4=PRcO_VeF<&bPK1_C)N>U>=:PTe858CX/EALR5WF,c>-A
)TCAX8RL/#21:Peb>.SI(.JK5@1/GP.g[@\#MBDSY>__>U9KA1D,X&F@SKO+MN;:
9<-C#^g:PU3BGbFD,;;I9N2Q<b,J[5V&ef8e8b\fd<5O2)KD+cKCV=8MF/F9F_^U
E<F8DLFd>Dc7[WS9X6,HZ<LIB<4^)MBZ)3/C7CZK,^V2.WPAB36@)Z32MR]Z4#.6
PAMKVXQaLE\VMHJLM3TeSB@V;a-EV]((1_O7S+BPSeCJ0>;=B32S60?W;Z]Ld3@\
Y-IP8&AR&KZBc@g,W,V9S,M.BNJ/4??L;MbZ&M+XM9dcFF(-TVIScT?d,@:WXeWG
Y?OV7?-=BcGC7+S;_;79UUE5c0b=W90#N/1FNYE#W^c/_PbKfRd7.7O_J\:^TP2C
;@aX3>3GNgYNAYLF=PKQN8JORBZ[X\PB6-#/V.G>d[JFVVS81ZLBJARZ@;6[RAG-
5,:]5361Z\TX;^6?OSBI/f9\&VH+6Td(()[^[]]31<AeFV^DPJ>K^0C)TH,F5^GJ
_a4a@-/2OV1GH^&;K\Cd[R/3+/1b@,dBAC(b,J_6/3Kb^K_d0fVNB+(4V@..45?V
TR/21UbbYC4PTT[1cV(</-E:bHa_I8?f48T4(]6?JBBQ5ACY]bOYSOD3B#)94F#I
>\4MaKc4D8A2GZM40X=&e/)2.J5<cQK=83<Z-)<KR)0_J7-W2NGPf4T:4Iee(^+d
afeHf&:>Mdd//\L00/]9M]-IFION8Z(N7aQI92GAJ-1^<9@<Mf[f4G[I1H&-:H5X
TQMY#V,I\Lb3@b8dY\&?PX(O&WSO7#AS),JO65@;a^ABO8Z64c:WIN52HV,Q+CaB
JJEMfP&NP_?d.@3egN)SP@dF:@RJQ^H:?2ec>@Z=SDX=?6g(#_F<RHXN9?=Kd^d3
=Z_CM_.:]d99V8PDaA.KL(F)HcfG#)+W3\V+bN.4g/Q:C].ddb=a:XV@Iac+SMKA
^Sb8&a.ObX6H6]2ZMICK.JL[WLO-M7Nc;@N2OA1aMd:?<F^NCGCW5KJfIeM==-&7
9S;W6P-RGVF<>HI7IWPG-,BO/gM#FZ0ceaA#J41]9:X6N)a^KU&09T,]M#Sd/[&O
?;;3-OAJE#.P[(c_9&Q:7\T@caV37,BQ[2\Y&QRD/ZW<^F1F;HbQ9@Q^PN>[AXZc
ZW;>J0CZ];H=DYAL_T(9>@+R6JV.==>Ze-=I^U<HC5\0=]XbGK:#R1893eNO1KCR
ATFY#W5K+4Id]KLb3U#Q;&CZM+^C.gU9@LV9\VW?.J71G+O2A5Z[D5R:[@]TPc#X
QA-/O)eBQ/7W;ZaD9P2>GeC.M6V\=)?S>TX/&7RKE<FbZ[BE:(N56L8_YEK^V#GY
f9A/F6:^3-]-R;/0/<Q\0c\@?A<5J:aF(K;<O]f37gg?I-:=L-<:G\:/&?2.]GEH
N:A_<TM]GQAc2d<8A)f<S]K16.IZ(c=:;_aeER@5aLP);4ZM53b(&Xbb0029)DL8
afJ:4(A\a\.[5APJ3N7:5[O=-b/K&8K7VB903UC,F3D><],K0c6;T\)R.2,PE[?L
<HX0]K/Tf82.c.+6W/^BPF)IKZ]_g[XJX0d0GYM?;<,;g0XaEe1:[+W\XP8\/+UZ
QN)AIFS.?dg02K7Cc;AQb\,dB:4MM\G@Z-b<ZWL\SgGdCHf8@<#ER#Q8O7b.ZZXA
QeNVf4>GA^3FFLN=>(aZdCZPI;<Q?2.CH-cR:&O\PUEQdT/Lb@P8gO[)Z_a@SD40
a4bB+adb-Bf]@e;Y9CY(eQT]@I[@cK#(PH0]LE6:)C_M3.KFFG-,O<SB9T/8OHG^
.WQ0AR)PID5ZC5OYLUf-4&8\JW+/aZ(GH]K-UQ8=bH&K.PaY:K4f\0AS7\(SA\b/
_D;(G^7FNf8_1S5=Q?MC(=QJ^4OKRD<E@W5FLJf[=][<L3;51^MWc@WWf=]AXC2\
?1DT@M<D0/gDQV33.=K=F:C\21V9@7(5-.a<;\cRL\?2_>2=:UM7[5?]d7/Ze:QD
.LcZFf?VJXbEDdGZ-dS6;9.AaH9&/7f9I4\J9>QA5;B.,_aa-92/VO,RY9RI.+>I
ER#b,N@Q,TY8)eIX8VgMWD)3Q#6gLZ=]bd2ED]:YA_eQ+egBQ:+^=Z6,.7MTWS^+
fR@426<;_]=5^dY^)#P3Sd>[A?bVL3[DB790A-e6A0EE&0)9@;5?)P4W].]E+<Xd
9;<#,c8X\0Q=]LZ,H:D./:,C#0<^.@_NX7SRB>ODD4NaS2-2DU#c<RM=M>V8>;YC
(_3A2BE_LRcG+TD3^S@W1ZU+2=DfAZEeLd,M1W4Q9DG0>.S?MP_-WUAW+M[<McSI
RF_KO)F3,51);NbH1?W),G]XW2,UeTPPKHQTgbR&1PZN>B908d2&c_F=FR)]+L-=
7A#^/SdX3F\@>>(O0ARMg>6G]aR]M64L>X4RIA1#Ae]6<De6+I#;FFdgS@UW?4X2
?1FB.V47EE:FOA9V9@7JV7?6N:_0:=>/1f07D)3@eS[_ea-E6edVL+ES;183\DZR
&H.1Z6B5ODRLNE(+IQ9@_ZQ:^60b5^7B[^aLR7;,8PbG.]Z6NG6F\C#]GHP<9?7K
5bARPG<0G3VV1HA9&V73J=QaF51J10J1W<A-fWA,N,L-E[P@YX,J2S[@EZ_3[Y7/
I[I\J:Z6?c4SbC8PP:;/HITW.G)I1b3+>.TDPc8U+b9K9eT;Xe-7ccW4eM:^=,[\
2U:ba+B^ZEST-&M7^V3)cKSD,YgDf29HK&:XS^9#aG9QE7:=@1NG97K\I=Y.f&:B
f-5_J#C#6cC@Mc&O-]e_-[,1J9W3.N]I+22&(N(Y@OD)f@^.U_cV@?U^+,/2.Hd&
c]=@-AGD)2?7NT@?.C^>O9g\/#A3?TZ8QSK]POe2J+ZI&=Yg92d@<_7=@ZPI[@2U
53cXY)6@4e@Oe<<>#P_TYX0e2<gG&^EH.N5c2\L[\O04.Od.S(1T67R@Z75C21^V
S.gP&;?A=:M#Q8S=9cKb_C4Qe2VeX?a>USeb)I6^)e,cN<8cP=^S2:99b\3C>NJ]
Y?-0M41+<&)fCXH?+bLUDH/]><bHF]VE74&fZbe1)+,96KPBSF,[]4M>)->+B6Q?
]=f8=C7;cLIB(/=Fa\LSDBVdI_XHd2O,IeDOMO7f<U;d6)RO<>6/,QP_/K\/f>T#
d8^48\W\@>P6W;?IA.0C87b>SKdIKVT4FPDQQHRGXSZ6+dH@2BI5Y]WVTb]V\Q.F
;=g?=Q6_&(P@&U5,gd&9S_HbN)7LWZE^e]e>:.1WV/Q#cD,Xb[.@SVE0Q@ELg9?-
d1J0dC;1c])d_K:SD:3Z<@Q0bb^VG;-fJ(41^?,,W1=2g6:9XR(2164GH_D(BOER
_[+P^FA+Pb23X?>C>MHcF9gd;D5HPf)R_P5[H?<5K29LX@&SLJH@H=@e]80Y.)&L
WI=8BL2]P&TA=4Me[/[IM(7R0E?N4\QLU=5Q_;/^E@;.I&SZ+AAR;<=OB@EQQ]Uc
dK78PQL_fb._LX07P/dX[<dX+3\\L+9W@<e5;J7e^]g/7+6b583,+RQT-4YJ8]4C
\P&8W-1VX,;a7WS[^C.];CR><0WX-L_CFFQ_=YB.E4CPNX9b?cPG&:[dcKZ)F6JJ
]TDL]<;V^b4N/#)4gZ8EDL6QH@\:0&R9I+[_0-<-L28W&8Q]H?bf27X7O28fHA^T
P\-+KM4+[HZ,TK7Q]=Nda24UGWC=b)<LJ5>P00RgI;&6fBJcA8?LCgYITReIJ7;Z
-S.EV+11&_K_]<NII.ZR2dM>EJg5bVF7Bf1]D5CN7K-.T(:<bT58eG1f?B3J\FGJ
+@;>311BAP5O8AX4M&^-#8B:a3&&\IZ.^gF0CKaaPF5<8fSO8P#0RQT,fD(5&NFB
EWAP?54@,4_WfS;:R[U2,=_SW]BTJPM2D,<3:J&QM=U[Z&eECRB:1]-?P+Xf@Z>b
DBG,5W>0<fGbP[g_KF3)?M>RC+CDZ>M&L]P4Y74g9dEc^a#EWB-\KX;Q5W5FP8;A
Q0]TPfJGAad9;/Z4EIf+?(=8ER5#<Y-N4e]ZGXE@=D0E[9]AC95VU@5S<;RZ8c8Y
gK2II412YLLM2/ILR@NBB-]5J^Q&g.6B402KX-Zb+YE>ZD0C3.\Naf\ebEF(7?LV
Zd@fY(T.SC6#Y.;OZ3\aUZU+PS6U#2_<Vd^WB)D;PJeO+?M]^.DOgKY3G5bBJ>2G
LX9,aDa[5GZ3SKB7AW8].Y(VN_fN)cf@cRG(A,;X@9e3gK3FFH=_M6W9LEZ=MR9_
_M3Ne_M_==1X/.5Lc5c<-6TIVd/_1)GMSHH?L[c?,TN<+Bg3^KIWYefOQ0f9_=c<
_bL:]^VS,.S<W?WagI]]W4O786G=Z9BP0-;<P,(Z89LDYW>e?I99ROHVIV[6C=g)
B)=.=)EFTaA&HIR@DdXaRYZ6Zg@@,V]K@/;(+YQJ16=JRa))Z/e\NH3K)K0WQIdQ
YV8:9;/H3FT#24B.GM7>(;8/Jf04#N(O1,G,C2g7W^FfaAJAg9PcQ,OC3cI(Z&Fb
IILILP\]HPLRH\?0EIDK\cfT6.g)-f[;fX;-aF6N:<253G>R0SCT+T)-0NACI9=e
G9c/>[.E7I/5MNfeEYg<;dU.7>APbFM>0MGgI:Ba)2Z2c@2e8@_-9]EMAML[UZ0Z
A(^2+P=>+69A0dJe2>T)IWMVg^]/LWG#b1bb&]Cb&f/OY.aH_4FWd8Rc8.HF,+5f
ZKaENUB@A(K[?,;L<cK#6<5<(dHQ:;)Q#[<c[?KP6U]bdTeOHWRKVU8@:4KJV\B-
7SZ(>+D?0a\b@K]9BgH94)VCV^.ZIK\7F[](\PaJ3V[59,81L)^<\EU_/4I59Mf/
\7YDW#+P>ADEB/?).M]I\[O=YZ9#Eb&_?S,D8f&GT4XdX1QTF>/>3Y:>^Z,O^JL\
LD+fX;<;TAY3/?7/D6W9)FMTWBFC#\?#=U<FW&6:a]0SVC(BUVGN9>O.eMC\b_cP
S+\[7NA?QA)J8<&A&I4D.LL+K4LN9H+@0@9OBgW(>FIXVJdeeQa8\;c9-A+_c8X1
>-0GR0;YL8])4<f[^TMETcFV3>-,DVGR;VM\b@8MO,4N@5D_:+M\:-JcfU)TNP&-
a]5aM_5T0fg<bE4Z\9ET2K[D#<3O4,7CbESS.&T--8OI?C,gVHD(+]E^SJ&]_U1U
RW?N:06G-;7_3dLCA9a1G1-1AH/INM2WJcW][#b#B[e.I/7B5[_TT2OAIB/c(I;c
2R6a,U_7,c\a=XEVMVcL43N#NJT9]/-QX#)L;_UaK&[IWYV@faR:)YQJgF]5e])O
RI_ZH9b?WAc#@Ha5fOT_:\2I<EF5@^Y:@@MOR0ZPR[3???SEO2)&883QP72EM#]R
NQ&?f#10=,G@a^7T]e0946XN\];JQB@DKAM(@UaA\))@/3Ha.bBV?:X591JC^=V<
P[gOYaC^[ZCG86R>@gIc\K^H3#=(UP.3e+=00X#b1]0<3M.Ya4I-VQ2G>BG[RZ&B
Q[Y8\S)CQT42=E8Gg@@7,<KV4D>.JTH-DSV>LV/5]4I2H+8OT3:1HJUAAc-GM-#=
[JYbEEG_HD]#BAg^H4-&8H2-1JRE=OGRSLL8cV/@\>?+TLHQ-0=dfS5.J29=GGdN
U5<,1Z?c+Yf5B(6WJE.\3?NaaXAg:ZcfESHJ,-AGHYS<=Qf:&8<gQK-LI.TDIFc6
-;#\1d55>gED4VD-^TU:(fFD/OWa?3?H[Kdf9+\E3SU0S-?b,</;8(OaPb2HBCLN
_1M/S#41)7b,TE7+c0Z:9L@WUNCYBcW;gE+,>]DJA7@6A2KUAW[UgVAW86dNLP).
;KO5UHOTQ9H0?d6Fb/J=4a/,P/O\RI3e]O#]6@(@@K(8aF#ef:D38bHISZJM1)dA
>Af[5eeH,/1B,B^9XR]c-V7[43a^BGOIB;_L_<NF:;E2H^f>A_L(U]RX3SK_HPS#
)Y<4d#W<^F2SEP=?9/<=Pe?db-L+KZW15dad^Hd<1JeT9WZB.C#61+(I)9:,c;=7
b4:?FCHcd733XX(KBS:<e5N2H0\BNfBP<S5VUQ/3b2<6H]C4:_(>J,XTY9-gfE2Z
LF]Z2XRfU#ZX@c6Q1#3R>NI-PLeLXD.Y+dZ],:@V68K)>MWU#_L^-D[&0)H<Z3NX
[b^7]&I^HVA]U5<][,#/>CSJBU+=0GJ+1LV4WV,XfOJaA[@UKPWY6Q>:^7E04?RK
7I2?STXEPZDZWTNZ\4<F)G+^>3?eW#gWY4>@]FRY)YH>A(:(QUVXPO(c+HUOdYUD
7T=W=26EPcNcf<f3^/f3CfRd9ZN&V(\OA/46SH9E^^IV_BYD4W1(@HfBR9;_U-[E
:KKR(V;2..CHeYR:1100KRXH&,1X9[\FZ@4PV)R6+IIg<@C//]aZ;Ve1Ed5G(H,U
>B7M2cdegC,55ZY)TVF>8+E,=]\/L=RdJKAW;LE=f_5N4UcG,^b?J@(P;PfZ8AMC
g&(FH+.ZW/:c:&40D[X:AbW8=UM@>O>fES.9\^J@1T_4>;<DS;b:(Bc]e(IQ1K8:
K/>--#OH)-JWIKPNJXaQ>LMdANH5F3+A<]JIc=>78#I5\IA(,&X#QB18S+@&a:Y9
^:>ALST50/@_>5Qb.3RNfMZ#)Q20(b,/d?,G#3T#[g7-[BF8^BcW,Y8^46a4SfB<
E9JOHdUD(HGd,DX</+0.3E[a9,K)E/87dZYJ[-FU8-U:Q,0,(6=P2^YZ4\eK^Pd6
Cg.>,aN#A0f4]Xb)8#\\e=6G-#<GK#S8g-[.FaW2/ATTe\/I,Z?gB^XQf[8\Y7=K
(CK@6WRaH-C<MPC)(;Z2JNJ99g<^S#dd8,VZ:PMM:G77-)BHAREQ&[FDUA>3+-GL
W#H7,^&MATDd4#\3EZNKEM?>fUT=Q^ed&F0C\B]-UHbWB3:?=b(ScPML2\Z<6+cS
H.3TcJ-)?((3K#LbUW;4N.Aa8b&&^:^4_WcS3OU6&#QTU@aRNWV,YC4ReUN7N_EZ
8&X4AX>5D-.5e,L-P#@G^/Ae<J9>>7T>WS+=PK[U).Lg5F[>O:a[RPJ8LFWGR-[7
20Y]^FGJGO@EUFUM)I<MRTY=6QFBHOVO/g-V5cJeLC#(JJC6?^K_,#WKZ7G4O&/P
.,2VUUJFNCLca3.XDT).DHSYQNOBdT_,70Z)+AG,RY6)H5cZ\[bL,ZTX&&aVJ8KD
RXWI:S#Z,S_[fKQeIc+IORL5QGbM1\_g@M5YF_-?)+4)EBFXZK(KN<?J&H^\P2><
QA;14Z1;2_F2EH,+F:Yaa8Y#2L<bdEIN[OZ3d^VeYU4K]X1UOHCE@I7I],GWLWO(
0g1W>fbJ.&2IBH6):D6.:9FZ6Z(GFVS._;?9[bXBQ_DOa4:-bf8eY1V&_gB)K\<M
;eLY:=^BL.(f=JAZb^?LfPMP:#H])C6F3FJ<EA4e^0]DQ^GS6EN4=@f.ag(<g)Z>
4AcLK1SPc596Ud(<I14IF150eS;bUS>0ET]419U:&Hd?D14CfSM+A>XN82/6CRTd
SfDPZb-R(703I7.[IF&)T^P+d+.(1]Hf@91>BT,(Se<YZ<gcNACSL-F2&D2^?28F
W\Y>+S<a,VZ^?Z+O2&+f+4Q+QHT(-b;>W_F@fKSDf^b]Lg>b=XN;^J4H>?+MY#SH
RYHVG8FX@@H45G3.5(C&<f^_=>P&1HRC_-9eGN;bM(.9_VfC,Y6C;Sf.Y9@]8F\H
4V1ZF[:D>E=#CIc(S<XLI7c;TB-?=:QUO\4N\Dd?LRTGEJ29:01<JO--J]Y?GFU/
]B=FU/CVKV;T]F9SHRAX=.MVB&XFe;&SFYBWXXQZ(HAKLHJ#d]);K#S9>+BC1:&<
&Z.U[A:Q=A.dQ^4\2<_)@/2gN+X5NC[_<P]QR31aNV4d0cdOf7?JLIG#cVI75:?X
SgEb4MP>a.4)@BGRO6^.K_A(OeP1YJC?/0XfF9VW_LXcfe&<OC48CIUMaVZAP(0]
)V4TaDPV<#M)/]ZG#O&NB7c.7Z,];>gI2S^]2OANS;79?<,4MDg#^:-fMLA2KNSI
fg]+\6ZANGH=E<7M3QGL7:G-,W#W\V^SFCf)?d5--/fX>U&<[^;]C#g7(,=B@&1a
[J.bQPe0FFIeVaV+:-@cX025bgcLVWg>JG+P/b[Q2K.[V46Ua7VPbGV9D&HU=FJ6
JR)1e@[g7G_bUed>e\HZfU-G8\CED#;a75L\L@K&N8a4A).d@QP:;O@4DJ2+2)84
8)U+>IA=Y7_X8bY9UR>MS2CK:77;FH]Nc,UCJ>CHcI/.Xd8,@f0W-QYdI,VE-RL8
@Q2JD02Rb7WAN=>+U\U1MX(F);/)Q#9=V(LBYJ27PF+(G(,g:[8fcAFcMIJc3e]>
TY)ZP.3+IK,Qg8UZbR+PfIQ9E^e,<82b,1W/cAf=)9dJ7+>GF<F86<CIWE6>\<1Z
&P1eNTW,0;N0O_#ST@CY:g6]?8N]MHe&12)D^S\)gZAN^P5E>e,915ZO8+M[0UXR
;IA/fUX<V;\TAE64f\c:&;g,#e-U&6C]AYV.L)H^2V4c.6L65#+A+.G07TZNagX/
>TA+ME31&e,2e0eIc(UW6I@@WQCQ:@T?&(EE^LJ[6V.aKb/U0/,DD@:GA<+a6K[b
He&GMPY1HP9?ZeN1f.4\IW0_).P76W[;cQ5JT>8WS62Y>N1DJ-U^,4;&,-eA6Q5_
I#KF&b(d<C]e:-IdR=O/?HbX.]+Y<QI3IbZgR-a7K0K3QaW6LTN4+CA+7bUR[\Sg
Z[7=1H?=7VLSRV(2\5F:]4E:KLQSa\8HBc\g07))EX-FOBFWXT-H)YOIIC\6aH/7
cB.bME>e9ZT1]F;b4QAA?fU4DU(8MB8W7e.8eRc#9^7WNBNZaEG9<1gUR#[JN_eX
c9E#T;=D/R2&_)>H=Mg;)?aR&]TR=082^26f(/b;-HZO@M#.;7+]>aLd.ULKP>=V
H9gV+NGaObCD3M[Mf3[PG>_16X-Pa9-[HO7\]C-R^ZBNQW+&dWZX;JS]6GB-@Xdb
)@G#&>5Y^EJ0HVG]:^T4M1=NCQ?I8-P^31@eOb#FJA<828D=TFWDREd#5K45ZEKA
#e_<2UPJP97HS7cXZ#X;K=0gXL;7I2(\573fTY+2)F_S[IZD0C?#0Y6RA#;.)eMd
12&E)#R2Z3XeA]4+=W+ZU1gW>7U6941b6R];.Q@\M:cc&?:7Pa1[:?M0ZCH_^87?
dC;\HN/fH(/-e[HL=1Q#RgQ9HgDIf#+7?)HeEUbg\B3<IW.87@(#KEGUV7;G/+_g
\V\Z_#\V<QD70;(LCN9Y-6Nd#VK;+Re]\R(IEfD#\G/8DRQ<]<dKV^LQ#C\@KB#3
_1BFQd-.4JM2,4#;)AZLSSYR4C49[<Q&6@FE@VeDeRfS3#Z7(bb[c1Pfa+CaH[M;
44+5fG,(Z4Q)KI2B7.)?]NU[QWWeTL2gZHUX:/,KA+61ZKPaSTQWZ2/33]C-E<(g
.=g([S6R^1I&G<=X1?>f(MAU,MK[1F[_4B15=W\Z+7d=HPJXg,2S,.PWf[e(;V&)
@\D^DTV-faa4W?-\RQG#Z]L=8G/YBHE;C,gX(cOaG4CNa7ZIK/ZF(4b.;:J[@3D9
4,T1?4XfcA0@QbTa821:&.G->NTV/cCC5)G.gR^Jg>2KAJRWA7gLCZKQH[Sac,a\
1FQIH3/XIaGLE9?6H--\c]UO>gDDM.g0;^KC82P^)S956WFA\)<c5LFK8I1J_AW:
HLcA?Q@gZ&?QRK<+6_;66<1e2=LE0A0bcQ:7L;I?8,^)^BHMLT_&:6e?+;bf6Q/C
gQTaCW9Q-^9>ff0LP[PM[fXcS8EI=cG.PKPZUJA/(&2&=L0FJR)HH^@f<AWfe9U^
&C0c163+ZF3N)ZQPd(>)g37_bd7SW6;XdL0@6A/W./9KB.L8<0ScWVJE1Lg@5c>1
475YN:,SH[H&d^4Va:e+?V.1c,SB8EBc8&3G6GCV9g#:B#_^gI)1_@MHBL?5R0_&
S:d(F\f?)A1[2QPf#TFeC?9W50O[^Z-.][@5Oa6P21F3QWa>#Vf7:G(B3C5e7c3M
>/C#O0)R4B7[EX-C-f_UPDZ<eYA):AW=\EDW[19Z+NPD<;C=QJ54,H7<D7KX]@29
>JgE9K\E?Ed\X,5bcf40H@3ZR1;PKMLO=@]/K\5X.ZQ7(^dP)^[S>e/e7[64#TJK
P=V6;YXO-eKLa5Y>)bYgK3&/Q&Ie[D1>R[3(?#dS@T[NJb.=&@f8/5/I,6ec&=aO
P_F=/&e#ZM=MQL<B_+5-1bQT0L5Q:&fJ_Dd<UU<Kg:V2a(JQM?^R0Y>DX54HTb]Z
Wc)O;/]L(A5geF@1cKCT#[J(>ECTW-ONgVX,+,.VMXRJ@S4S@^XIWcc[P/Y0;,+[
MBP?0:#[+c0\Y_=N(NIY&DF#JBK__ZG;+_W.XH+9C7XB_4G]U[gbcS&HY-?W9&FJ
AR6dfNfNb/X<4M+;bMYI>?DB>[DfW,JKc6SC=;X5d0(;_eU#6=NQ7>Q962f.UaU6
[87(J0cdaK-aC4W>W9IP.0^[d?Q;@C_.eb<1DS=L\Y62;f11LMJ(NZF=Sb<&_@,G
fS7++KOJP0>N]JQI3NFW,L(5gZ+>]FELQXH[A<VgXO09O[9IB.J2X&b,gdA\;7/X
JRM+Na[Q_U+#1[gOG-+N.aI.,D6#TfJ&^ab87fUWf^GSL6Y[Z4bHMS(O<7P>KgNe
ET.gL>3V/FUX@S)N22.(M)PMG[,gI#4C_Ua)@9:UeI[D;2,S6D99&T<(B0?:,4Yb
-e^A63=SR+X(+/DIG_\aLT=;=/D<1Q,c8bK4IFN<_54282]Ug@8:7HW>g+e,EWY+
\NLcHK(c@>O^0J-?Q_UH,3-^D#+4c8G.cK4)\H]g,F#/:M\DIB_#LS2=563=PF7a
\J8R3Q/A2d8WID\eMKK0@830WMZ]/g2DQg80:gMX>4#P(\P-ecA\/64DG38(b8K-
WNTUPQd:^D.:5TJ.SdgdQbD)Z3R\?KWcDXdRO:Hdf<D7=a/H@QQT.B96W3TWdN;^
&>B)5R</eKRdJJM.d[?47#P^T/PQZK3U-K]Q,XDUXM+8Vc__Ce_(&bE1Q&/HP4.:
=)AD/437L24J3A(IU95(:(Z[5RT^43Rb7G[83@egRgS6(AbQa8Dc+^UPZ;I48L04
OSWTX[@2N3HcPL&SQ4Gg@1SGdH^L:92QB#8YG/b(+D(_9KISWLT?Y_X@#_c+:a-+
0.[a7Wdg??H<@I0^6,]QFTOM39]O#]_;V3V9e#.E:NPDE?b]0d4+8:RZ=1cO;[+V
E-C]OUB[/?:DMBLFbI5d0R__Z6)G96FVg0_DJ/52+@W6JN4aLg4C_W/68FJ&JEV4
B<NCWF]?G_0f1/<P_[18]:>2<@fOIL]I[5H(=V,I[[887d5+^#9+[_@&e0efURfd
BL6R1?38(WBgH8D3\ZU4_.L_G]WK./-Z16NW@F(J&>\2C:&X#=cW#TMH\=56TU_P
(M16BKI:V/N^Z75]X\_9I9]GU9GGMfKE7GT:K1-&7@?b@e^7V^HE_NV;=VS-]CD#
MfIGR#Jdg7.g)><XBS8dc0E9eDUO,VZ>,^FBHO.bMaWZ)Ue]b:QV?T?QVKP8^@EY
SB,eU&59M3P-E55?].D.,8?.#gR26eG1DO?aB,5.[@a;-QB/9;N2c975]\;PH6WZ
A0D#52EX>H(_f--^Q,K8)8^@<HA-5E0b0#T,0V1EBLadXD^4##[ZBc\0(Y&<X/76
fU_e<POI-_[5#eY+TS:(T[W,LS]/K+VS_F6K\=8]Y,+4_3gH]:g>&&V:.FbQQ[Y1
V(.;bH^HH(?)L;2bLe2E4-5HcaYL494<f2>3Y1_2-O)F3+d6?B.bV9EC4D3><O:/
>I]AR8b1\I=:?YT#Bb4D.>4GH1Ued4A/gE31ZCH@A2ANSQ8-+KIV>(/KI]DCDBHB
;f?G.cXDVKF-:XP^@UP[<g9N4=SD0E=YaH>ITVY?H@4Ge(]RO;C;E;Z=R7_<c^Q;
[A4D3;c[1,@&,_Jb<#c98f3Y?UC3U/UJGH)gJ.g?.<\=Z7YC/79B:=eB]4KP/W[_
@g=:=8S&@ZXe^c29/ACa;aZ>UBV;Cg/^EQ&_.\TT7KX+^dOGUK-=a2(Y\_0.C5_a
-3LNZFIHScXOO[=IV+Z&a+>(9[18[.J\S#KKL2ME)]I>EI/),>BXBE>S0C/8PJdU
OH])?\e+WE;Df)0#^7,F-3_S)P45B>+-5S2Sf#QJ7Y#8IU_B7Lg-f5REIbfd-F1c
C,Y;TIde,=QUd07<9.\?O5KM],L;N>S6LeP?Lf+@76D185Cb>TDc4R?>9^0LJK/,
@g,1P\dLIWV,^g+SQZ8C.<N;#4:ffVA6S6&?ILNVWF;EO(+:7-Y]JUN[KK_P.S9Q
/1fd-8=60M@/,0Q=R[,c;[TfY\@;aH7-,_.Xd]X1Z#BCG.;0MP8XUOWG?TR--G=-
+MZ&fe+#^Ia0(DWDE[GSP(]:FOR;1?NK@0,M.JV)D7Mc_8.K=JCRQ6R4METI<U?9
gcF=Pg<35fIPS8BJ-F7[?A3=d\Q<TFB^]R.-F9)g\WL?&[)VXXb_FQ-3<aZ3L>7L
Y6\c+C<K)O:BFN[USDG738(>)>I<cD>Q&@4Se8CB(49X?Qg//@71DLX=U;]&MBZ#
(-<P\^H,d_(4R^21Z]Z>Q;.[<)3]#D/c42J.PSA7QB_WN,cQ+a.)M8Q,\).A>M#G
^A#CT[SU_H-U_:Z5A)NNd?M>\\BWDL,4R?I]?B?[+WHBeSZ(R(6S+_]/H:4V6\CZ
JKbPBa0_e#28;ZFJgZ:/,9WGE1Y3[<6@f]3:B8bY/QgP(^)VHeK_P#S4E79TWKKX
\Bf2g<(A>7@2M;1cT4BH:4^8T9(FBX=@b(/&d(Bd=7>+f<^2OF(K=2\6W;e4;@+7
35FS[,OQaA[N_f+#+g^gS]\&);KT,Yc2Vg4Uf?4f7eS(NDPP#=^=C?D,A:U9W7bS
V<BFCe6eD:X&KacI7H41)-?TAf=3#N?QF54M+47O94E0IR?Y/abX8GH>N#XEb./3
\dE[C61BdXbCT6RB[d#TaP7bCegFUb1HY/)WJR428-]Pc<+(-S?,@5\US5Y8Gg4Z
<1;eYTWE6(e^dN;<;SYUgT8<8-Z?;LfbS_P,U2]94W<MJTdAMdbBe1#T#d&)R.\F
S^3>EE,\&W<L(BBH;HMY3II6W1EK\a.)691GFPcMdbB[g&#\)@12<LWcZQ_;BE0\
[e_91A5ZHHD\V3E(6DU7FZ)G^Z9[L<;AJe<:(B?b/QXSM@1N+Q;05F^/d6B#EH0H
/5H@U[0NF._EO+:f(<CHP:(IQCb06_,UWR<#4f15:<<EE\ecO_e.-C?ATU7&,>N]
6f]XLZX==+B&T&b=DHdFRCZg)IbR1W+<G3AL)WAG[6^2>&4504H@)]G7[SaO))]V
:(W4QJO9]7<HX0.gMb?K[___4eS:c4bTZQ&C(G?-.\8eA0>#[ONK^)7B,^N1L8d3
T]L9?OL&Nc29ae-9USMH)d&VU<a2]Wf^T+J&W6N<gFQY>g/Ya[WPKb\IEY/d#J9R
V;0VXC8DGX8PY3M):?2L?+L/_U_[Z2(QK#_F5.BcB]UcQ+Pa:Ob40&O9V/d:#,DP
-^;UHI35TQXfe8LXIF[U@e01)?B9KHHP4GL&O4--E<SWB\fKE@S(G23D-V@,?SDe
3IJESbH1f1R6;S&]gN.TJ#SK+dE;#8_RTT\8>E-T:=(O<6a\U0:@)?_DW[;Ub3ba
fNKN48B&HO#I<S3^.D3e1CW22b+W&SL?9AV)bUeC[LKCD/b)\MATNZ=ggbU.XVE.
C/=2WRHD+YZ[RNY.]=;&T0/,>\_Qc>SJY2RMRXC0Y1<8#e+]VLc-\[]M[LIa&6X_
g^MRXMK\^Yf0?5[/Y0M+T@36)26c663Ff/fOCYX<[+cXZ,(?RMF5d#L;4\f0R:Zg
-4OUXA(HcM27AQf2-YLR]b@3C-TJGXA^.MdeO=eAW1FIXggW7<<RH?/PcHd:b?_?
eSLMQ,MPS8]UTEA<7212^_I/9(aF<U=W6OOQ+HcO2^8bA@H9UC0[\XN1&=@HF[8[
9=E=Pa-+cI3P7_=(b(G>3.CfU72T<)QN4E\8W@2P]S#UO84)ORC8Y-:VA?(0ICT;
PeAdXA.A,C=EAQ(J#gL3\D1b)0EGYAQR4-FCZVXe:g0XW]6G@RASGW+2^9aT6R\9
_]R#/cgg-XE6Z:D;0Kf@,=4RQ#229aXgHK5V<Ca;KJ.DAS=F(.L2c6D:MT_VcTRQ
T]_,e#X,1fA)7][UJ&VVD,UEe.>CXQO??-6W2:=V_f:BW_5ZD,T?C8Z[T[J6:S\(
Vg=DG]#e@)FG.M<K(J?9-?:6I?E&@(=.ZIa-&S&@8\d0&LMB=.Z+H6gG+W1AC7D2
_=A->bGb?_Ma;).dZHOR5<>;)DEa_c1I9[HLe-CaU8gSU(RHG<W<YX6A^?&+,WSY
?P9MCLGb6UNFI_2Y?g(E//7UZNR\\.WGK1&&[\O-W>F)CC?KeY,-+,a=_Y9(>=/c
YEJ6Rf&=.X1^d@a;85]MVD3<YXSc@#+?NY]X^C;>_K0U4#/].3H0E2b9O:>4?cT[
Y0af\HPdU0=<cZBR<AAeWQdQ</ZgO@3E4(BfaB6&\;RD6C]:M>Bgc,d&?1c#?AY2
]XN+g[DdZUb;M-VO1SMR)UM.@d&[AdIf)(KAC:(&KZ^SBMfDd]]S/(&Mg2-2FS;K
KV;<aL).S0:7U/5/)EW#\#7@D6^JM.L-A\fMF&QWX4U.F554<]?SCO+/PAVb.TbJ
JcN_,.Tc.P[<C1Xe[OcWN@D?X^_^fQ-Ef),W]bL5Z)-ME90aP^NT6QHWf1a9>@8)
bA0TcR.fRT#AZ0V7=;;<ZS-DM>#LIOd-B,+c25JOY_U1@I^OU)G8HCc=9ZY#QVK<
d89&?K+)ZeOeeJD11V;3/>c7.V3UN]d/\B=gNac=CBDXFJbU+-2.Sa>^WDI#547.
,ZG0SX4W^ZXM[#Dbbg?[PO^O3()-J4MUG[BGUZe46KL^[ZeE<I14E@17LG#\F8&I
3d3LK7df]N9+3/(Hg6<J.-R&f_+I@,);SH@O29?PLaT7NWGP?VV<Z00[3UYS=9T\
4DK;NK<SEgYR3WOFd?=LX(CS@YJ;NF15B6-fa[UIBI]5\60/RKNP1CLfS#\g;)V5
S]BAEY.4@VK5W#H(Z(ZUATSKTg@U-Y7O;VQ6fXO)T:0]6_4(8UP.+7P_Z]6GBS(?
7;NF2Z:UN5TPg>6_@1\\A2@SLUg9,HA7W\cGN4KSH,^]_XM_g9/0D8E:dGW7+DN#
@.1fDYeR,SXGScXNFU7U=D\GbWLK>Z<+GGNJ8<:?48RO;8DCdY1A60B#SNQP23JI
()7Yf\c(VVb,4Z2+LH5/b((?9#G=ZeHQ2#]_]c^9W4UG#&8=8(PNd>a4S^W;R+QA
A2U@Tf0-Y/LeAbc@VRKG9Qe.,HgZ_+.3M,H_S--]QQe;=0D@#-dQgba;O<\_)7N:
H\QJE[Y,SXR>7K2OOVKg)+5._+EWD10b_UGH4Z5WEabITP&L>?Y-Rg?K-R]WWFJ6
/8BGd^4<dO0E[-a5g73g3efH.YCKQ9,dC:NHM]MT)V_EWRC,^Fd3SF3c@[A60;<O
KQ5JQ_dD/&>V+_\VDG7^0ASV8HCG3>UZ5TbOcBe0MMFZQ6_b3fbZM?:F^S7YXI/e
-?U^Ue-<NC=H,I71US&aDOgMZG+UGE4E\AX;IBX(BM8^OM@VPX=@Hc^D>3<f3CGb
+[RaBV9B@/.b>e=9I^._;?]T(R@,:_<b+PRO&#O28CZ;Ob]C7<:-(R0C7?7[+YY3
-c/KA-a8gdG6#.eAcW#f#d1IY</PUa^3NL:-=M[0:XQ,+H(a-^L[P63Ff;M-\^[4
\4LR>7TC;3)BH)J7\<NOgM,&9J+6S8EWM;T/cC#V-CUG<.8/EIBf:+,JM[RN-O]@
eU(P>V/9Cc;P5^:Z<[XN0V#2DgW_0,#OVCXYY++-#RS-RI;TA:d)QWKWF>,J^gSE
fXg)<V3T:N;KKbTQN:/)[39C6Gg&I[+R&3BE@\(3L,R4EGU@5b&LXGCc>#,W\&+E
\3d/#_)f0S&A=dRV,;\d:T2U?40D0eMTA=UQQbK94F^;?,L<D5.4<eO8LO6R1g7(
U]^-^eJdJH,<b;?Y^.TQX?+]bFX84\aQG/BK)U:I@;5b7U]V9WHI>f4)5eD(U?>^
F1,NAUK<U=B@5&?FSfL:OPHcAVe5B)gOL_\?CR[_R0T0<AI97]74Gf(D66FA9HPK
I/a>R.)#8?eCNFL0>=U)C=WJF@D8=^d8D:=RXOd67(U/E?Gd5FdD<YVD\F2/3^@.
;4VVXN\[H+ICK:c9-0A--WL>G6UC?8gF^R1#dR1)W\#:See/A;M@5?f?^gK6I<BV
(?GRCfXcT\X@Y^C-SV##CM<AR:4S3,D:SNL57IK([2,.OXa9KOEf?\T;/03UBOB-
AdKe=-/Z4UJKIfe\K4BMURg]FL3I=S&MPO7d&W6-N3Q?&eB0/IL[1C60aagKX)bD
K+PR3b[:eH-(;UgU-Ob6\PDR=(0&YagT1UTT2QR(EHE+)]Y/5P#(N2M-7b6).\T)
YN\AdPVDM4SF\3@<4I4f^Q^<[=:-b/;LUPZY^4IeLR-)IPb8d:5)5&K=>c&>590S
0gEDXY.fg=D0bd(?1S;L6c0DecEb96XfLFe:9HJb=Z-EM(OK+H#ac&\S_H^.VOc9
/LW95MM)E,I.9YC\<PWY@OMCX&Z5?6b//geC3BKcO5[84PE@>+81D/-P#LSP>U(#
T6[<FJ@d@9)cVgX]+]F]bfeR,.+PJ\:7-?c2-@;=c=60MF=>TMQI_5QB_Q9#0TbS
+XECBL]QYgQaS7-4(3+I2bEEV1VC_G;G^\bcB[N:8>7KgK8T2>bVXVYQA.Qe^)-L
eCI8J#5e525LZNKR8]4U^@N5+4cGDWVd?9AN4#AdIgXTE5P-+E&0X&,D\\XY..5,
C^_ZG0<4S5Y]MD_b4:9A4HDHec=FaDN8DgdKcN&9XDV@8),8?PJ[+.U[^afIFV&>
2C,JJOZC@-RN:-65@fM[ZYE@2(7M.&[<5AGAUB]E2>f-.-HVBJ0[_UUVd=95X6.,
aTM&PFP1GSQ8H+2Q7=;;X5EX,Ba^]<Q5bMJM18.>40R]DEF.egaH.0fZIdH\X1I_
0dX(L/LF^R8@IfLLB7?&BP\;Y7f:#FX3/=H(WSSfbS;KA?CA_[-U]YDA@P#WP2-X
3>\P(Ec]1#TP:L++.ZX&3AGf32KI+<KA08X_I2-;,Rdff9dZ&R64Y]7JIc40ZDA)
Lbe2H7eg^4CCMB2]).;GP(b=)769M)U_X\,1(=fWA@^RBN].#Tf,6LH][CAT\&b<
&+?9KQ=-JYI+PRLIVW2RLXGI=Fc6gcLcQ^MO:TG.M&a(F7VO:]PB])Sa26bGE22J
c]baIB>?@62\/:a:VJLMDV]QfR-Q(J4H#24bgZ#(#L@/,JKGYUKe@@Y)f]P(:N<D
(Ac(39HV3.YbO8PA1)Y2,:2:\--Ed1,QCZ/QQ[/ZSK5WWMXFFLBf6bNL8E,&6AU<
90ZO@.QD2H/UYFe/QEgYbVH.L32:WGF?N3?QA>DcBVLe3P3+:1d@[9?UVXQTdG],
]#CGNZP7ge/OfeH<)0ECJB7=V+2M3d.T<]bc=?W(&bR8^d+=RI++1;:2&(2M8]&/
S7Y?WX_VMN95/)48;U@+.D82NF[1NYR2fSEI@P.2M64YV?0c5a4cVKXMRgfFMf[A
>HE.cE_UP(5bHMI65<IZ>,_Td<4^@fMPI-A2b1/_E^>9cK4C4.aOUODOX<;=K03e
L)RN,/gW+5+[GUIT7OagH;D2K7]GcU+=fc#<IOa.5X\6+H&ZS^9;Zc>VP>e]ga,R
EFZJfQ-^6QW:3P,BB;@LO#-\;4XBH^9AC^KB.A1I<(MU9M&Z4Be@6G16C8G\-bUC
5N51gNMEJ0@5M->(S#_eNK>G/:YI<WPf.E)G=8HT^-=1I/5);7DbOcIGH3E92K+\
DY+^6<0cH93D[Cd\f4-(6))?Z<g+T_Ua\3e,SW[3+5JJ[cLGecETY)8NJ-2VfCd6
@L[R0A/^CN@aTcLfKBTe\W-\fEW+<8L-b?fQZM+QV0dVc+S@9SC@ED?AL;9RO)e\
G]8GJEC3V5aQ?dE,ZEeaUV^c^1H3)/1a3I_.EG)/+aYCN7Zg[b4YU)Ga.OKaC6c#
?RNZ-5-P<eZ1>I&RV/,g,(-YO:&2GA^:D>DB8R?R3QaY&;.CAZF18R8:g-<da83[
AgL[^LZDCLdeIeDg0/QG4d2Z(Ng\bMb2[7N[DG,^<<W-ETR<\KZJU0?_@5aY#?Od
X.6YZ]XS\g?(@VXdNYLV[YYUG)dge(EWO_TAL0(8Oc-U<bIFVD.I3U-\D(5g3?d;
bfUOE(0BZ,I1AZRa6O@/KPO_e>/,,LPPIB=6fJGdBRQ+QJd5Jf8@Y2R3^(7<^@;#
(HAe=.?9Y)OK.c.@?B5OM5AH8_W.U?SZQ=C2O0TCb6/55(=Q_/WBP1(H82<AS6B>
ZFC_[eZL[77=cD&=gPHP\/4,H_T?FK0L<eGEd>-E>YJJ>g.O3T?-cd=,P;bYZP-6
NKfHM,gca8SO]2=+X@XgEbQdJPbRg:a+^MNVWbWM&\UX-0X=7RKXV1Q5R:>9d.JW
:/JQ5,YHV)[>5b87EeWa[=a&[=[AIZ7/2=Ja(,=(d6OQRTN4RA/W#JTCW8>e0Z:d
^caOH9&f?2XJdEaW#6N_FB]8=.>O+f8]\(1Fb7LbGCS_@7;QdIJg_L292.CZ3EUG
/9e/.##aP]/Q^Id;aTP\Zb.;4F@Y10<453]B3ZNWAQFFPP4e2?DL@PEX2P:UZ;/a
K.6dO6:DD+LfOXVGH,2AePDdX]Ycca>SF2H<D_5FJQM=+JXbHKJ,TZ:Y]?d?=fEV
@7LF8\gfa-A8=[d[J_;b4d61K/Ad+^3GZTP3BAgcH6=16)-dN@I78Ka&0M#Zf?87
dOG),<d@3TLW/O[<R>5=W.G-cf7F-7Da@D0_S=&-#^.683=MXLS_]=.Z&DL?d68G
<:#PM;\V7>LW>TW_Lg/]]@1(,YRgU_9=#AddR;=\)I(5?][O?P3)V:M7@8@[DROF
Udb+QG^0cZE]R&,H+C@Y9B7=LSWWYW+OHfC\E8-AZ48e9)K&-J3GZH4BE8-Me#GT
Sb71:SNK#;\4@Zcd_=A4JEOL01ZB:R-QACc(ae=0bY4A8b4=JYaFX&44+aWF\aeA
bP&)62-H9.=&Y=d0f-@1JLPFB7e7&ZFS[eT0NSEE#ND[GAQM>DV39E?bYGUPAH#>
\RR;.g(3;f]L_)<bAF9JH?@WDL;g]RO@\cf<(^46^CM\:U2U\gLM2c;T8OIFC??e
&JJ8=cGb]H1LB-;99bRIX(<2#Te4^b06_\I:]FW6/\A>[aF8]HAD<I0B9N<ef03M
<f\E2C9+#)24eD=;aA;5@4Q>2\-P0YCCgM:LKM)MWKIA#9]Q-<-RZ<3N2MB2d4+R
W;cf;[WCQ5KJF29P+NMLI_S;?<Y)--L2UC@)_AU-2g:\OddFM_OfC)IF)d=V(JXC
K.;9=@&1#)13AVf,\eZFPN#0I3]gH@6A9_<@WM^GTX-IQ^.0_RXET<VAN7#;MR+F
H<FOV@OE&O^22<b(7\/-_3.g#ON\O)\0[K0W:P0ZOVGY+BZ5T-[_:D6XPEWP>^N]
SJaDM#?-_9d\Be,a8_aM>ScA52<cfXMI?I=J/]IT\d&WOYTOeGeI+Ee6aK)SD([S
#,-dUc&,f&caXCIcEHP9(U0^\2+<<=ODG4Sd[9+d:C[WeCaB0/9[OJf>B/eC4OAe
c;A7=4(E\_4M/;@DVb@9_?>Q]g8&(Gg\.EHSa^KV/QMF:Q?_>1K,<b;?7KR,HPXL
(IN[AV5B?9AK>X7<fM^E-Y=LGe@>bD70J0,RVZ[#9_I[?>eME?.8BL3SN=M7CaeF
&G3@0]5cG\QS4A]5;-A;IU_,7A(1->.7#Q@HE:V]Fe?71Y-db;G6fcL^,@([2#(2
H+[=Q8#dP=@KBA-a0CSHCQb#4\]cCA+^7dT:F&,cV=BGL<D(gNM5W&3fHRGUEMBO
CMS0NTde=A.R\UdM<180#,@Ga8,[>C<&aAGbOOCJ-S?O]P6HLZYa]1;eF7#;g8L:
C5ePPA^@5N:;UVV_F\4:^NS_T(;g[D+\VTAH+K=P6+<U\g0\g@gbA5_PZGUDc7]_
F.XTK=WF3@-E-bK+ZP54XJS#SY<gJ02;eGfG/&_B8e_JBXR0Q:9O8EUc-X+G6E6N
(S9d?/)Eb&&N)3gQbDdCR^KZ>XdQWM]54XUUKP7QB7S?0@2Y(cc=,XYIJD/?cb5#
_:Q/<R5NfXRC,Ff49?e[:R(#YNg-B\Z(&E0SF:Ag.dEC.Zae>D&<CL960X8B-/_&
))dG35;YR7YbECF9\A&IU\?BUUM#<M\P5V)@FfXa^XXA(1J,,7UfADadL1ZcKER[
fG.G)+77IM(d0.AgVO,1V#Z.FE#.Tbab8K.56<K5;f0\J&<Q+gU4P,g[_T,\++\e
g=3PS0=Z.=[F]HaKMIL;ML59O?U1=dBAaZ31OGQ)ODZ9HWJS>GLCFR6AVH=PE&O1
<X8,#&4722g@PZ2FZZdEcVCA?M^2WW7>IB]B&b<8-1e:EZ;[=D9^Id/]5R/aD+-.
^.6dD-0BSA:DG[,\M7]C.2EW14d,_[_[7QKV;@0a5OTOeP>[81FbOEZNT4_V\ZQL
BgTR)[gU#]/UPFNJNE]HT((<7;SfUYC,5#BSGSOS]XJSFH-Q\(4CO8,d+.JKM7-^
#6J.^9PMBO(UP]/?P8U9c\5T7?XSR]0W]HZPBF@V=2KZ#>:<#P7272eIg550DK6;
ge,N6PaYM8_F=&_Y.-18DTO20]7(4BR\,,c7&WRaP]6U#\Z/6/Y=bD]OJd\&/S1@
^16,GA52SKYC+_g/#\a^=.,TN:7QZ-T?=gZE/(H#561G.LQR07=T#?HJ6?]@f[Be
>A9NS>cAPP3Da4M<7PVeXOD<7:\IV@D+&/1J\851F><IRM_aKKC)50a2QR_QQCD-
&\(=7b^IZQ-K(\:8-Z#E3PdONE;UXEQ_[A\1ce[-DID,P+1IBd5:dB@:6O;WQP8B
8R/;EELB(@,C)]#U,+E<c@&S)a_;f,1N+(O<<^S(#fU&^d6,=P(@ZcNG3Rb:\+a-
D.e]LLB1BB(/:5-</a:-FZBCZOI@D)b(Fd1DHG[2A#[M+8-039II]+MW<M^S7LAZ
9/+Xf63UAHCGd(,N8RTL>fA-I7Ka0AR3-W[P-++>ZVbI[UBFN;Q\2.;@8>0fT2IP
6R4b=&9fb>\9^/8HK;dV@2A78A-,=Y++N^^RE,eK0<09UGJ4,]E<[cUN@dCFN3.c
6PFJ]@+H.)#Gb+1+P\YbJZc2.;^J8=Pd)TU-#O)gP7LGLM1D=[g(+8DDE&c)aX:f
52\a4S&4b4VfGP;@CNL[#U-\W?K<d-1?1H+XE\WL1LRbLbZQ?/3D;MY]^ALG\/SO
]S[daX-@VO;1O;f6A?c22/c,.gQZcfUSVJ/USGIb)K33g@)gcMF6^E=ae32GgN#-
Pd_f/T.9d5>-_VSI9\CWZ@Z)Bb?O9R#KL=<M7Kc.-F60\/7E]9YVSTM[#&DO[4\@
^(T^<>O0GdD-d^P&W(e;:N\7PA.LNY=L]QU7.B:4F2QQ@R]D#X0d:ZK<>Seb.S_G
VH,C8YK><RQH^A=,fb,gH_T3KA^Ld__XYQ)HGB<+)^+#8dgZP8H5MFOG>8cH/JU8
bb,g31BdL^2[fTf:>656#[02]O0)\RKVE=aBT1&7faPMBB6D:U.VI=?,FH1KCTCD
FLUBH(U5=ZUT_,YM?,AQTNY-6c1d=WWAJNBb>X.X[A-(B[H9FL)7C]9CC)=G7]]b
SJ.C)H[Jc>DL>8Z_Q;OXJIVI.IU4?ZTCD+V1>BINB33.-N#Cd?IP5J&^\Q8#Q[bW
c\]0c;K.^,fd]1W0,;QU?9\HA^T16c^V98QO4fOX[:KP90.W@#PRFbLB60_Pdf9^
]CRWCFT1SVL+3OIP.XDd<A_P7ZTJ:g0P>BEKHAE^X:&P6+MW3K?#?6^g@O-VN)eG
b@SZ,NSCfPG56OYDD>gYHc=LJ?0_S3M-?EdL2S<P(-_d4CK8Pe1^C[>S-W8]FVST
F@g[4-Z8\YQI122]QVGI@,3gPe,TFL2;50@8]WdAFOIgCNRcde@7K(F+\\GDC0eD
g/cb7g(5S^I9d1#@53fN4#^=fEC_P181^R2bC&.KXHNX9UeJ1HYO?.,QLeGATI_(
_F#P<\K-<A]2K5TU@V)J>(W9,]=)Fgdf+=6R#@J7J6-eEG][Y0N;CY<O#1a2_7d\
^++dZ/Cfe9,<K#NZ-RWDFXXGOTCR\LC&;S2[^[=:\M&T]-)(]1D>7.2.<7AQ)Q).
7J2+O4S;65>;@UFF_M6M@Mg3eC]E35L(ORcJJK56)eTe=;/V?e]1@X]FN[M(<DD:
24H[VZ3YX29#L&Fc76\6E;<-a9&(cL.Z@)(WfbJLL1YEXXQ0FBTDR+NO3(E2FJ@5
#WeQ.,7<P\gALV0M,<g[A11c)O>Rd?GQQ1cGf6a6P3IfSQf+Q:-\(DEQ<EKU/Of3
=[@1eQ,<>ILO?49La(JI2ZEX5_,:IZVbcC;LEIcTZQb[FKJX<9PI6AFK8eG:cf^H
)\KA4EX3OfQ:J/_;>[Mb^a:A_bU\(-(^1H@X3][c<D=3?&BTC>,MB1WW+?eD-4OL
2U9)YFU]3\K.b&WX&4b\\I9dECXTdcUN+=<NP7WbW<X\7e>a.3[Ia-58[dS2O6SO
^O9\K@R)N(T]:X7IQEB-&cZ:<9GQ535U+:\QB.:TSQPVJ#e4(F]P^MSJ62fI2<aE
[4HFVg.@e+eM7fR(3CSR)_FV+Z&JNO)?>&Z6_6SJdQGP4J&D9_eA?ZQ_.5-U5:0G
?E,O[RSG:=_]d_XKB]+WeFN882E-X3ERKggMDgc[/V&E<QH:D4[HZgSa5c@.UK;-
g)d\Gaa-HaIEbFc@.E73H0]U07PgCG3W;TO@Md0G[DP5b5:1H]XC]dWTC:XG+_@5
D3_e-?R8KVM&\3c3T=&UBQ0NH+B:)>PH:F/UP3f\@M8AV.c0<RE;JAG#\E=a0<]c
Q(8EJS:WTW5L1LdF:A_J]OJ5S?-Q#>-NDYM8\2KDM2_;Y-4JeUfJc\X+S;d7L8@2
S7<bL^E14U(T4NNaL0JfAg/=+\IGAT,8d?KT_aO,YH\<E9ON\TM)_e9YC8_9;<4:
0CbN-GI55CT&.bN_eEbfBGdCV6XaIc&g<?a88D?Ad]0NR@<SCW\G5IO)-MP.;.80
AdJg+/:CD<Y(_0<LC#d&#;ecNE]dM/WSfHgcZcDSJSSW[-.2SH6/R)&CJ&e?KV=H
g^;[?UQR3eD](75f;KI-@CPT)X6GU1@&a;_/N\VCMYFR2Q_eX+6>GU,bM7&6Y;Y=
Z]XUP:D[eFD0_OPWb=#AU,Z6YZSG_RFH)N@PQ)BZH[eIRB(2A)#DCFYW9#M:7YD^
dUfQJ1&X0]bKce/<:d&Oa_ZfX9V6.TbU[@cfD-23I&BC37:D/0Ba@V-_B&E[?]dD
(#+I4^:db;Lb?1^-BBO+YScTQWEebVG.5[a4F34TI-C[9UdS=D@;PUT4&?5UC6D+
DIAbAa6BXE5&.K=JD9#0FU6FM@.Sa#]8N&Kf9:UEL^@-Aa+a8eN<Nb.-Q#7^,_ON
NCCQd<T6OVVRK/;<,2</RV1//f6N:cL\dP_L_L#6V:ZDA/CHPLH5.^g&=YC6]BJ]
LHH\1I)O\WMGcd<:ISJ]\M:M9W;R9?eMH[<3FR&[FLZ^8bN7KEd&aXgWTV<]fE13
Lg7@,]RS@SIX7A&=BR6?>J:LBfEc499;,#@H..5H>WbS7Za90eS[0P#>NY8O9V4A
PNVAN)]+Q^Za8A:>@aQTdCK5P^HPO6LC6P5>+_.CgG/=9KE6)]9g)dE;+0H1FDYg
gJ.f))BZP?ZGOX>,LZR/IBY&NTA]T]QU(40&>XA\11DP,EaF9\Q6B#?e^YDVQ2#5
eU7W8F)c9[:S6d6)e7c)54d8d<L&5Y9A]>LC[K5/g7W_aTMWfM09QBIaBQWPKZ#U
19=5\0\c<Zeg-W+.;PK(ETEdC;3GYR_\:fE]9aDB.CTfT[L.2+?e&<@JaBa=4Z7+
T@/7-5.K0-O2O1O#YU^K]5D-(5d_V?g_IM_cQZ8W@JXg0\5^VbF0I;#_/[3,LGa\
0T9Y2;<ObL@Mg-?.GbeQUQR1&W[ML)7WeV]BWeU24_c-3FHb?=eSQC+9A[gXJ+e9
TeaLRgb04.D+&=A?07Y[>ZB&.(.R?/\4U-)>aTJ_+e6[,3<)b2<W5,(N+RU]bDY7
9;TAff>UCA#A7DaHL3JY3J7J4CM0POUY0D_6c>Rf#V&ZF9Q(R@)MYcW8N_,QU&c:
/S+SH1<M2G@@>ZCaS^RY>VT/eGdU>/QF4eY3.?UWac<T.NZ&;Ye28ScecS+e(@OB
2D./H)-[-KN.LCW2VZI]^LZ(88_g1:RQCdUIC.Ba,ce5#[^F<Ea3X3JNS4dV.8-b
_4CJN=:CdF&6_)XO3ZaY\/S6?<SSg</Cd&8C,H7RZUMOfH[KdfHNHcJNI$
`endprotected

`protected
XMF0@Z@g-O.>Y_/d6J?TS8;]@aV&JD\?.g>g2Ua,_=?=.,c7=CY.()-\JdO2@Q_F
LC5.&,OCb<gXb_OU+2Idc_;]3$
`endprotected

//vcs_lic_vip_protect
  `protected
QV>]WD2E)95>0]^7Pa3aV0@#?2&-9#+23TfWP^NNA<)HW6GAJ)6T1(6H/,0S-d7+
fKLVT+;KX;+b-CU#c2e2=UDWAD+_&c:X(T&0M):JAfb.--#fLI)V4f0=)PK.[@bG
?dL@SQ4:JU-85&f-5\d->Q_TD9D/]d=5+LfK>\J8ZL;gRHG6e[f^-)d6JNV)5D^I
-_I+Ed44,X;CO-=/MJ9]R(5O_F>BLN:Cf;D0M2_H.N,X)4V?Q):N(3J7P2;A+8>c
PI.563-MAN?GNTD8&Oc99X?/E@6GB\9BLE3FK0D(G24g@F:VFU]-KbWR.9S2IGIL
=+]MG3R\2bM/Q+0b1g;H4U^5G+1ZW(0CTJUZ<XgV8/@[=[e+=_Nea&aPLcA0S9X@
a/(??3?fIZJH.+^bIY]YZ61[S6cMV[eI4IW,2W7CPE6:LSS\4KQQ8O1eYP:ZH>>e
&8H5e18Oc=Y/JTO<B.JY:U^2#dg>Y3>YEf<]f6AJHg+FB=Ud[>IA:#EJb7L+/f&T
;BX:T6Y9]PR<c>-M_4II]8(OV;eDV3YV67e0cLP97:4?7]K3\e<KF7a.fAJ+1-9A
&;KAH2[2RQXeMFbRQIHL>cOf]Z60D0.7S-Xg0167J=?>S/H:cbD,;e4NE>L9MLN_
#K&8.[E1#LL=(,f[dVXRF9KT/1J=0ILNSJV48.\c]EN(=dR/YBd^e)\W93](-+7,
9d5+Y-e>a0Kb^Z;1^R+6+F&gUW@]E-I9G^5B_-??M&Y38Gg]6WGb-IbUN\fA/99c
Z#<LFKUGgFB]<\4Aa-W,R=AaT[aO2[3&7URA7D=JJ5LPbZ+9K,e)IWdV5DO]P+)4
VW0<:C3_/II6_U2?da;f)8K7CJ.#3,==),YM=S5SeG_+X3[3PS-2F8<7A(D2IbAW
cCfbI\O7GaN\00G5+L=FK3Sd52Of@f4O+>1,D023[^;Q=+ZfQ3LYBbS=T:J0Bd9A
37DE5Eg9][3B1eb]AWZKRUc/7AKd+C>N52GbId@(^Z<b8_H33^&^GH8Ef+ZV_gX=
8EfH6gTg[Da[SYXa[<NX/_CLXS)c@_5X-2>6@F5R8]8X+Bb33F\cNI#TB+NCM?f\
;UFaJdXM+6HSQ+5B&O-;)cT-2M)g]KM]C:1T>e#+.IZYbaDGb7L,L8G8I6=/>aM#
]-V5JM0.;Y.#6>/4^R<;4(2>,C?Ra.a^e?>XG3B9RL;dHd18(SXHbWE56PKYPA&-
d(>Z]fSI#(g3@8g4#-[_4O/V_P5\bOR4f,?O+IN6\6A5ac8\^OMf2-[&1#4/0[Q5
;dL_VdCK)&#82U;_ICMg>PI,SLa9;9<c9,@IC<QN7e]8&ZWLgRa]TQ_SA\P#TH=#
XU9E75\W@)4;--0<RM]-N6T^2;Ne_bG,IYX^e_7YXTK;M127D^fR)feA<B570OL]
(W,DA8&4OEHNATUfeLO+1AT3fIebW]BC_Y.DY-XDaJ[8?cA3#73YMD&fZ9#[J59,
bG.;ea@#R-=0YEBK3E/Q.D/7Pc8<L(BQQb^&FF4:BL:TIG8EPZ#IF<]AC]FS_N8[
_A/e,MX#FK-VX:[];>2LOK)?04NA.0Wb-]<A,JI(Vf[EKgBcZWb4Y2DB=NdDcNV&
9d0#&DT7)OY=-TXE2XT@_KcS<MYV5=P-@=2EG[C>@d7RAVKW,bI9eYA9Q.RT3L8^
PZ,:HR6GP/A//5f/WTLF(8V1^G&Oc<geJ@_:ZZGggebSg=DRBIQ-PU:dWKABdM?;
fe<eA_@a:JEB>T.6eV[gBS^>QZ;bdI)X2EL?#&ERV7,WcMb=Z/.YfE+gWF<PQ6Q)
FRE3HH\MW\_N<O113b>5_N]4OP?3;B;XQY4_BcRUE@2)D^/T,[#8JPC7S+;F5(ZE
)Z]Og0bI>-[HXEMI[GRE-K,g1+?TC6g8,?gKX==6;-<[-Jbdb]\4-=Ug[>4@)8W-
+43_+8;#]GQR_=5U[I^MdE(K@b]D5<M:@9B>U]<E@eT8Mg0cEQ06(e^<_TOg>K<[
J=ePNa;Z\/\,.Y/F]&IU4WMeKJ-J8>ME/DBdU82@,=Zbf7FBD82US[=,(d^]dg.e
OJa2?f5-GFf[.06Rdc4QLLV^W/=)AJH:=85EDTW+NQ554VE3UN([+[g7e30W0?Xd
B6>,WCUOVJ,B2U3g]X-MX2=B24Y@QAL7H3dYa]0bFKMc(#PD2SN#ceA6,5dVRFU+
92(PQ5Y]S:SNbNFMAE=.WEN4OJ#_gYe]U<,#.MF-^1c05I[X<Q]fMLAS]3Y5d#Sc
^C7gL;@3JD2P#[)dY=AU)W.5HgSO79?[V.3=LEP[KIHO3R7ECfO7&F)?)TLC,,\S
I4&5<SI73bY]WY&&2aTCU;@^81X_E6?1W>ZM51+TQ-2P?&86A]+2<[U1_U^L:5A]
A6fB(7aB#4PV&-0OHI-JQ2Ac/X//9.@I2?aDSSMX6PHEIB-\b/CZKDJN^6C<A1Y#
NFgE,T>;YETVR>I>9]]Jd;J-eBTX>D&P0WZQS-<<6X^_a\5M[SM).Ma<b#=.cVKH
b037HaTdIdaW,SK0]=W+A1aX1IC1egGYc5<Kc1J0-)WG\PZ\EgL3?P_3Y2d>.3]S
)_fgV[:GXX]bNH__Y^eaQ^a?5gL&C^GRC5QE8_B/K9^gKEKf3C>6Z&@_b^H?\ScJ
W60gSUcJ4XVS-J6LH>BB<GaTb8/WZYM]=[&@=DeV-[]<MUZBG.ZW#Q9ZdGOLcH,1
@@;_[3P\L@,^cTRFE3#4;3E_W3&ZL3cE9(/I(e<&CAR6/N_TG=Qg+dV(3MZMd?@5
&dA4_dUTE\4:N@<-B&O#Q2SgZN287K5)7a3gWA[)O\W64d\DM/;34_142Q.T.J>_
dZ(JPD\,\c,&^U\,e9G3_f0S\C]<5)EU>N#c6XB)#[CP)@SK9DW2+_WG()BUf2Q^
^gMHHfeXX_#36])KCJ#=>0L&GDALC+7073K^SD35<3O4P#C#(A=a85J3)U)N2G0a
93fJV>07]g6;09)?-cU9X]9>O=6(ADdDcXL65HTc,L>0bBVHg\.:Ab=,ec4<JAL^
5?db&@;f>Z&]UE;?9TaMPeN1/X\7;(O]-7D]4E90S4R+GL3bc(5G1G3GLR76-=D@
X6JJJVC5?)Re=2F?K3SQ;e,OZ7&a/[/N?)9E+\TPMUQ,][8@G7MN.8LD9L/aMD[+
QF.[4,050,dA6@dI0R,@#W]>@f:SS&1J4>Hc:J0[2SZQ;@4.IW@^g^dg?D;4^0+A
-(X2O.]M:6MK5f63cLIE^)?eXU9VN;H&@I>P87H?(&1PJ.[R,RU\D+E2VfC1<<A2
<(bO-<AV>,c1:RC/?;&JXKD(0Z11Y?Vf.L.dS:EVRb]X5@M,>@RR4CI&HLgT]?IM
_61;#:d[#(eW(JAY]>TM\TDCI3g^+2g4_B^5DFCJ\5MR^M@#\:W[[/3T5R4O3eK-
Vf?OfR.d)N1VVGM5R3FYMHG_AZV55dEcY&G6(:A2IgTb0&IS6C0OI;;R[VZ+\30B
&<cB.9/(P]/NGE4Zg1?EW;,Y;NeDe.;+M0W(a969UP[-JSM(e=>6=BY(UM9ZaCTY
]>KC8;-bTY5&>M;cI2AM-)AWIdE(6PK]b<Y,]5-1+BWRa?1MA.UQP^&Bf(EVC(M:
@cWNab:JOF>;@(NYO+eX7:;ELH_bFI#0dF.S7)WDM_/O#OP8gP=;O6E)<BC/<,b6
X;.IWAT]ZYe(9e6BBQFW=6][I2fB79C(GaX5D_O8&DF#<,-H,:UK4[SeV&#2L_2N
6_aR#VU)+dUV-,58PE,7D)WBbM6K+9_N8Z@JAJ#XgO0Bc-d27JMaH6I__?aO/11U
W-59@DZ9Z&/37(Q<)A1S1XP)BGLRX]1b(7Y4Q&^Vf]<gb>Q]D^C&2E:+HK^UbMYA
8)fU>DS.5GFFg,.5\3Va#VC06.A[1?V(d(f(23@g8=g1)@V<EN,<D>VYG@)dH=OR
XaK@O#ZfCBIY1)[Cf#?69(R].^Ccd[@I2aWF9&c0IV5-7QNdWH0f+H_KZSU6QK&+
4]H/#D#+WgI^IHc[YP6AD_/2Z>V32/56,RANWH:<5;(K:A46DM);N#\fQWGT\OF(
YL4I@V3V;@?DTYFA.V>)Be.NNaM>ZK;f:2OCFWa:G/a7f?>O<?76_E^YaH(3e>+S
b9KZaXK8,O3[AY&L7E:JdS0TN9Xb[=GH.B&6<:@L2/CgCA,]TS9,-M&QZP=N<J]Z
F;-G1QOU=6(1AR@9^Aff/?91Vb+)0VV0>a0K]c+6X,MX;+P:2CZH^P&L&==+G<A+
UTG785_7bP;T8_7B/B&3LEYgY?>-#f>]BYJ^6RA]d54AW:MVaGg4SNaeT,#[N-81
@L+^#?6E6;2=FF4XS+QCf^N)RPO5][5bDXWKRbQA,GS+-)Ic)6U6?#0J7Oe8^4V<
:6Y&E-f,D_O\?Fg>GRWc+F@46].&0^?Teb=#2DaR=b4TS&H40OU3>PJEUG?8=ING
P?>+1\ZS.(1@DbBV_8,D4C^82NfEZDW&-1)G[NB(_7A3^>J&C:O<g67c3+2@_0MP
#LbbgGA=9gB2IfFTcGET0UeOE(F:4BHYd5.a1]I^P)R^U>^HT>Z+O=+bQ@f0IdD-
d)e]^,.c.Y-,JK9?M_eEHB0-^X0-TdTVQL.e(DJ@0+T+,-,&@R/d(AI0AGX[1^;J
Nf?CWFb9^D]QS=.^5@ggDKB+VZ#ZeK/5;V>3g7#7Mb,76IK]-]985I)egWS^/-;9
@/(SAD>e=54RM-)LMCc+\Ob&SNR/5?DNV7O)@_QcZBgI,dB.&>A;;7=Q(GdMG:NV
KTW0cGDd.dQUOCU6e>;CS^KI[=CSS2E]:J,U?^0YX#cNWW#;\bNSO:@Tf]]BD7=c
86Y@f\a;JU?P4Uf6D[NdYVDS)9.94L25)\b&;/?bRA]dJD3^gCA1==DJFHB-X<=>
H?A44d2H4b6X5LZ]YTC<K?Y\96NZIZa17#=OFO#VWCX;8&-4aSD3@g5I,C0WQ/9:
fUANW/^D?-.[Bg=,ZDVdK8:SK;OB&9?_OK5<4Xea7M[TfUaHF)1eI=JYR1+5VM57
B@YG:d\K8b;G=3:Y)-6RdY.e[6#IUfS-IX??\8B#+^E->^]WMBdVfc+@1]QG-APB
c0?/d;N(E6b3f@SJM1HbK>c@fEP7&:U)],2<-QU8X=0SFXW;S<W^4Xg&W6d)aNG4
99_F)<#=.bX@KYR]^=@L[9VII;HSS>Va@A3GJ30_-IgIB-@TBWT],_b8JA,[YPD9
?#BNK6B9):6Q0GSecN7LLPGF)CCL9JdH3T=U9IeU(,X.^+<\7:OY3^(S7[-4//Je
U#._L:DMc7J&_ISU^F><PI)a@AbDV>cW^6R[.+U:cQ>ee?X2aG/A-(48_\(A7AJE
_>(Q+F/[#BeBI72,[Y^/X54M@6&OWO^FaW+20-H[A.N)X^W?gFO6g^0EJ+4:?AbL
UOQ.aVVM1X;cX,4.<<;>5V[,.JAJ>WN\.H^gg6A2?dK=;5XACLX3X:5]+Uf+7ILH
E>DcC4;V-=ORFR_JOL=PbO7&aTR2LYWZFe8-B7XRWZMRSEE_Ug,6+c#ffI15Ig;P
,6,W;Z.;=]Q6B+^RCDW[>(.S>UNET@_eVIU_ODNaVC--)e11ZJc2[J9W[5BF2=UR
RTJ=.8N,.,(La?a@@XOB@8MYMAFDFfc+AggJD6(dE>^3HbA@UE:J[V@e:fLM:?fT
<9Xd@],Y6^4]TB[?L+?eFfD.>WbX_HPg]L.Q[TBPIg.9R1^gf>L8EFI;Td?T?cO)
^H)9NA])g)a9VADZ#b>117^4;Dd.6]9N9,/-L/7f(;1-gMG3WO9V63KOSNVcc,,:
/&^PfKBYWQ[LaS]S#Hb?3dc]GR27a823KL/VgJF[CY96fR5RH#6:8g^V+P;cg]2c
FF3[B_/JHL,69M6L4/JY;IRJ5I\)]5NN9#ea=aZ@JY[1I4B7g<Dg\d3/X_.,0H4M
I\F&bBgRY6?Y_?III[gOaDa1^?>A-;GY#0L=N9PRUF8L(.[CeeP1[8S197We?\4U
T<]RV1S>>KC&<137;QJ[EFUN6JROUQebX[SLRH^3g<#.G4P32M;&cfG?[;b-SR-H
J7.;2&c@.acR(=:2B0&GV&AW#P#O5H4K)9G.=J^e49&8Sb.D6C;b0-1@Z_PaX93c
&X:L&>OYM^:RIM;8)JM2fQY]DKY6OH#7-.QAR_)O\@aEDC/d5SQ5fQ3]MTO.=J><
IO4>?aF?])c0X1_[GQ..@c4=D35T/&JC6P3S=VcN1_THLB\9<#,=5)aB@AScCd[;
0_?a8c.E@[XC(6_0TN7a)cOAT(,bRNJE&c7AcO).Y]g2dY[VK_1cQ[<-caWNG=a<
38Id1@=^Z++C=D@d_W1c>?T6+WS:]T8RMKDONWII1Dec=LaJ^SZ7cK-75@9&#1L?
@&#L(G373eNfPGLN+&KR)ZATBE@QFGbXb49b:;\L]1(JNb_O1bV&ZILaYMaE,IW[
;[1QR&-/,ZZ9d1<c&XgNG5Y[+Bddaf#3TLYa/FS:6;U:KcNbY[3G1&g^3=0,0;=#
D_P<VH2KY.MDd,_f6OFV,dY7NAa[^S2;_G+FgWRS9FRgWUO,fY1Z.&-AM]FVD(L(
?fC]<Q^1@--U1E:gB:7g&H<:c45^dee2XEJ89]F0+U^NdeF3@9Y-ZQFb&X_V6;\N
;f5NJI>,3Z#MbZ>a9\7L.>;S4=2CUc7DP6>1)MXcHVW(O2L)ZcP8M.N^Q72.&,>&
;A/&>X0M/f:/dL1,L7dZJeO^:Y8caS5@dfA6CV:^/_/9GHIZ>3gcV9,)22)d:E<R
WBK8NG@>7=d(+S#7J0#E(0L3e13PM7bA_K&;LW-C;aZ+;JGfWXO6CP0,BZ:^KW,T
^ZT8+0^ceO2N.>EPcLG-6P:5_Vc1J7+A7K,D]<HYC9CWZQD@Q]Z0SF5W+.eG_16X
?RE12&g3I^HdHK^0.bROXQ?8?<fXbZ[.T9gEL^/(?+#e@ZF,1F2:)f1M+\J5IQ)D
Y+R<;a1I_E:._KO\7O/X78&CEAAN\V@BMbOZCJEBHYU<LWA,1#A8Za@R7?&4RL61
U=(P1#V#gBc?BL3/Vf2B9Z(G/#RC]QN9HG.Da#5XRU,R7Z^Ma;89g(:WXg/YKS-@
-YCLgA/=:^7(U+I=3]]d;c?]G3=4d[EH0K3T1Ke?ZK.d;_V(Z9>RE.@e<:=Q2aI(
R#0N5PGeNUO_-#O/,4gJ:^(9O_f3J4NA-g03@>/XFI_BfAI1Raa^[;W5\S<=T_=-
L-W;.A=\EC9,d(+OY.:f;.IX@\Y@eNR_NM<N/WL1dJa60aH;2J^]JAQUff.4D?:&
=K4:eBOLC[SfZ/4R8LIAUZNVHOHcc6DaM^?>&U^]b4^\I:ZQ+;9f3MI9^J;(K/Ya
#ad).(&g0+>6&.G,#KPf?CF3;N)_fN8]6LN\T/)90&2Q]bg_L5TD1T893MP7U?MI
6M4U.][QS.ZL2PDE;c<3a6J#=]8T_Z=?S6JS(1UC6aCYSSb8_@D@=T.Ja,PY)5C)
R&4COF)1TW&Z]L4\8ZcCSH9:1HU<0([7,P?c9WcbIb4M.3R>-35L>K]HO)cc/d&f
I\<#4NZ.bZ+9EaA,R+]I;1#I5KULFGc8K5JcLd0E7P(a&8W7)L\a#-d&/@,+?FV5
-;N6-I<<P4Qg=fP2W(J^U\g8<7AJbE_KGJ_\U./d@[>+Pf+fHPfN&D7C)FY@^3Dg
c,<<VE[I7,IHYb^@(gbG<]O7a1,GR3-O\d.2OG19HONDWC_@@7RTb=2F7C?Sd#O&
:ELFDFBM?):==9.0]P-V_1a4NT9:[MZ+-:X^TDaX)MY+/QR\+dYDa/b9[LV@7\[U
X-]\\15:E)4,0eQW2ZN_KZ&,W<Df;<5E[=6^5Dc5N8UOc=/M[QSf:G?IY)5)Y0#B
CNW18gF9d6OG_R7WLHR<QWGUH&H#(VK05>?S.\@]aZDaYH(W8,UWDAW?^cD1<3Z1
<KFAE-4I4T-J:V2g9S(5043R(YgM:&28CI9RQAQ]W]MUIPT^fEYD1FX#>-G8J<YV
YR70[TTaH&N=U]5:bVUO5O6UFDM1&;AP?&_TU(\F;,.>&7]_PSO,U:7P)V?/2Nd]
dbAHTI2O\]:)2<H+dEH&3FVfO32C8Z>2bY._>(X^RLb7^<O(S&,Z4B^M,b+R>C@L
(U#7G1]8]J]a7Z(EV-/CNgP@e\+=D@g/DMHI>#SgD?1JF[&&/PTc)SLRILP776^)
QgVM.4fV,cL+S[GH9Z^YJ9Va1NXP:5RU&.11aVeY1TXdV[ZbK0EcLDE9\gDXY#:6
Y][b=CSEO1V>4\WeDW#3>XQc^#F<#T8Q2G:?d,_7QNEgD5Pg.+-D:&N#87O<PW]6
.@H5OGdTXZ&ZM>>R4,F)QD8QGJB_7=_E+LC-D0O\QAY[G/OgKB#Y<=)2^^H[a:[H
KD^0WI>V_Q^a370UeEFS5f9TFYCa,a(<E6d>(D=.-=e17^C5TAW;FRd[<?c&(+@C
A1S6>8O72E>+[F.H,O5bAWA(.M6L,&]Af0\-a[-96#dP>G=IIAXb2U0ZS70bMf.Q
+XA)SQWX8?QH=2)08WZ#HB.5)d&8\Kb&4a=>,>;7EV+,e[JT.aQ8.bTY2Y,#5-G1
MbV7aFa]U2H7f;IJ:AIfX2eQ?Y[e=\eg_ZO>HY\GTLXI:ESW,32<;DV#+c]DFbS)
:W6B&9542-WNY]\fM2a9++I(1G36;2LY(0U?--J6\YY:_RWIXW?B);Q;]YSFfY+J
cJA8GVAW\0N=/>7&@4Zc@[FP9BSQ?ET?PRdOJ^;C1MLF&,_+-6Ng[H0M_@#?.#MH
R:g8Nf,89TcVM<T4/WJV\-LT[V_G6f+9gQAe6G+51fB]D);G+I7=?L=++Q^We&EG
ONVF8)f3d=^dT#[C,BXeH+N1]aWY9fR5gRC.a#f>(Y4Vg[a=KJ23PU@^,bbFB7Cb
Ja)FC\#PeDcD>Q);3]?&ZL9+7gYNZ9X@PaZ.+7U<8?bFFVT&ORWY]SP#[0X1Y5>-
_ETO(aU?7/0YH(1RSf19cMEW509@9D\M>+]>@41g]UN(f#b7Y:N;ME(^Ha/X,I(.
1UI1MXH<X]MZ0>[0)366dYX_78@a(R9T)CUD/:&Q:?cB29=GbQL+QF&9\G)B.C<<
1;7c>_-OC?5R54#=O1HNfR7^MW\2gbb-//F2?BRY5&g]cRAbAV3KHWNAHE/OeGH[
&(9E0]#HL]=fWd+4;:<Z75(7e=2J#)(E@YL/_31X\2a>KX>H[+g<FMM9GAQ>Z1bf
?]d@M@5(W(C@/Q.S66K)-4=_Q[P?CJ\#B7Ibg9d(O](/&71\FU,#S1OJ>DF&7=f^
L--^U>:[9cTJJ_CL>;B<LH<WAB:^8?5Na&0^fQ8V#.)0<QUKHY6M]Te,0L?^\RW2
X41eP0T,/Ye_048KN>U9TBV#Rf38A>P2PL[I_T9EJ^<RM7V9.4?PE&\c(cZIN5@g
:JdU6;96SC9bB.FWQ/TVJCBX=90[HE#)AC;MI12D3&3<8e>L?O1+XTMeRZ:&9I;4
NJ50VQJT</C,HR1DNIcE.>J1+F=771C+/-.:]4DfEJQ2Yc&]0CZb^<9?6VEF[g)Z
O@_C;+P(DCQEWE9C\DZ&B-H98B<gKc[1H)N<V([BK1\)M&_PbF1]E\HEM_C4V;=V
CW,E.7#c\<S/LBY<1S[f2]251[e:#E>[,CPIV7fH1\Y,E4ZKCf4ESH1aRMI3d2FO
I-3DadQNa@Y#TbdK0?3e5H=IG^#f:FBX&,CV-fA>4LL,SYg44^-&[bSVJfQ&fXa)
b+2L<<WYeXS9U[UP4RW;:OG@HcH73@X8,LW/fZ)H/0&^]D.B(&\?gKe2H)<NTZK@
@dJKGYIb&?eeV3_L4&OOY]Rg0B9R0Mb6JSOYC[X35#)f=4BXFDGA(W?0E5.(Qe2f
Z54O\VC&Ne+1dGLWDJFXSC84ZAONIP=8[6&[>97#M((#5:Wg]:0ZE_-X:BQ#e5VH
UWb]aYBY2219H];T_8J?WT2@-bKMc/A[,?cDC5A2BdW)Kc&.9#FO8JALF;e3He9(
=@&S&,G94M8]9Z+?K_<UeI6g;3^^ZB@)3cI?J)]I^g];S>fEV,I4:dB<d)7-ZBV=
;;K3d^6O>&>E>,](@(I+=gE558C5,9Z4KFGAE,^-M/CD8<JPXgI0<W>b.A1(a(G/
4C22KI.#.[6?\3bL0IFab-JQB]K(T_-F30?E_JQ,6[G-Kb47-g]D<O#2/[cQYP1G
921ONE(VRFQ1F+09_&@?Y+68W@=:HN]G&_A@eT[9E;\O__W/32SSd6-Q@a-S#c,;
X;ES^L(]S+1X2)fME21H;]W1G:R8<1e(]=-f-Dd@PPd#=@f;P(<A9/e_P-9N2L#W
DJATIB@<J?6,Q>c7[:ROT.bADgdJ]CY(]K5I9Q\L9&8[0YJ96UKU]S??CZ6gL^RI
E\RH-=.8]MR0eKVLAZ7+bAREI@4_.[DI<PPPf^@d;G>IcQD<9G^4NT#[ZDY:I:,8
MO_GK\[YO5<9=S^\cH_]64R:S&+G>&d8[f1C_&(MG[Lg>GSB28,\LRFWg5J4@0;D
IF<cOIE?LZcURKUI&bXCU(8AbE-@f(cRKA?-+CPgWZ=7EDge(:EVYD1_^3[4(G\H
g-H:=0fL@9\VYd18M736G&]e@_&I#)c96UIgP)7X)6L54B5I\&f[^5g0>;SeC[Y3
NN?Hg6a=0T]<;;GYZAc8\e/46ZgL85<ITE9;3F3ME)-\OZ\@X&?+ECN(AIE/J9Ba
E;bJAX-gXba77eA#I+8N.UH0_\UFE60+K(WIGV[8-:=3LJcfZ.3Kg_/,,W].P)0X
gT?g\]FCKHdGH7>Q>0b8H97(Z;W3W-(4;V[Z@9f7]BPMDRHZ81_DL2.E<e#+=\X2
-ZC>;TO,TQ0<E(:4QW(,gP6I-\#6f<,]03TNT0-V2ULWMGdf37M(b80667?GU94e
AMd^YEHKUPYKSRVCaMK>F=0_WJ7I&&d<HUKP/])3RgZBOg3bN;)\:A<J;e,;E18V
I,-e9eeX_O0Oa1fg2c9f(JS561Hb<H\L/JZXFJLWR4)^BeLIQf\A>Y+DY1M>c=Rd
aJ>Kd=7)\ZMI\FXO\d3Y>6_=)CW+7f2^YM-::BR6^Rc>T7Q,a&<c\CL_M;&g6-]a
e7+0H28G?O8;0^CBb)U5<W_I(P2#bY/6AZg1LI9D>;9Ne1aHQb<W0gYN^>3H6K5:
\Hd[RA]=eZCM^K#0dfSW5RaB46>Wf(.WUVPc&B+#/U;Y>6cW(3D;U?V3Yd0WNM^2
1>e0gCgP0BVBJK-a;f.WAOC2]#fVPRd<2..2R]K8ID]DJM/@:2<-135:^FU[SFc7
<C:IbWPN)=Z5X5IRCab>C8UK4gPCV4a7@S^cfR^b<>AMd4NABI=)bcIQ?>DQ\0W;
c-LE\(T2[_1-:Q^H,AFN],(c:=9MH@5#0P3>N\5.BNO1XNUC)ZD\W=G&NF0Gf<=X
-IAg;)TV/EMQ\Q>1M@=V_PTeQ>=?,BKM3X\^E21LJI6:_)@WOTZ-D[Fa77XQ#dO-
[CJ\6>AC]113T_-2_Y<UMCeU:0=-<BW8#M((Y7XO2V:XN-QdTa^]D.e,,K0[EXb3
)1,Y4b3cIHIEC6Pg5\A(;V8QcL?_?JBPOH\^<5d@MY:WF6@QC6;KPQ^(4KODFM7f
ANbS4W[>C9a&^]_VgLNUQc=IN<3fMM]ZMAJ^LLKCWN_)BA^MIK4I^J?A9/9H\FbA
RON+TW3K5@V92V]C\0W>=125V3U09Y=/GAPY^5I8H)\DE3O(JfZbf28L,6V6UHV7
ASbK?645+)4baEMZfL4,HMPC<J@\fMa4Q-(1301X(/Y4-Rb9TD(;d^N63dUGCB/?
#IU:LB+KbX)8)5?ZU&)cg_K<#XXY#_SL3,W>e?D6ULL<Id6R+RQ_CO@DgFPU&-X:
3EO@E-=NC(KF=\<^XU/#Fe,80U@AFgXE[;N<#Z8^g5eg7,A]I28H5)0TJMFZ0M9R
FQ;D6+3]]_=5cdA=K-bLcBRW&GMb(@FH(:\_TM<7bCK@M@?5^]1@.U)L>]^69U-=
),(K1b&3@22)>c2<@f;MJ]T?_9ZT27DP2;,\3;4]I)HLEUL1cOO-fZ<eG2QR8])S
E>=B3EKRb_P_,VRW3,>K&RZ\6g-//XBY0\;46;dP&FXA6W8[Yf@GQ@S4KQ;YVW+?
,3]DLKQFKELEGPSC5/XTTN^JQ-cDX_3QAI7Y:^6A&]D_,X;KBR_SVHK+R>c_,V9L
9OG>cUcYfBZXJ?c0cY2CZ:8\C..1/KC(9U/O=M+T3AT8XMJgc-@Gd^C7d0[WSZ1<
F7dKKA,Pf4@LF]7_O4\I7e,Ga[</.X?CR:ZY#dPFP/VVU6278OUb/+UR=?K;-(;D
,SQ9SXd4OZcT;AA1MF+&;N)#OH@9_DWd#D@#RU.IefC:EaRYFQJXY+877f>X-4RN
E=C,E#N-J.OUMY>_K5F)FO,7&2bP1#c/0-)cN6/&A;O)>/3@U/++\+L+^98_cNYa
:^d@+.CD<JLMB:CJ,<bP:#YbO;L6/LZ8WZB?Da9DCO]gBD[S.ZS(Q\See<Q#Y)EF
Q<e@/GcE-;AKfZB]PAO03]Q^_L_;&fEU_^;W>,eKCKJ&PaBL@AK(EL8=MB1CELe;
:)<ZRJCBEf+^LQFBdXG-9@4_0Ag?3)JJEL=WIUF]bBUa/LGT40U:Pa@K737DMfC,
Gf54DIQa>\8[LL?A1(WOC7^G[FO#?NKS[@F&1bCTIe3bP(;B4UDIbcV=XA8+MCDb
<KgPAeIU+XO)Q2O]6@6YVgbVC(a\^:b&C[:7XUac^DE+<-#B04I0dN=(\[Gb9?)4
5).SELM==I0@ES]SHZ<)0\RL,MKNHPJ4]L:\_U/PD5HXX9g\]FRRW@U)Re+[0QAf
P]0197G7HG:dSW2S[0AM\Aa^\4X7T6SZaU(eNVN8JLbcg7\2J5KK(5/YD6M-@Jc(
G1@K0I(,Q(Q;S_))2gYU@?Z0H^-2U[&[<g6I0K<1LID&G=7fC^NC9=BSIR,PUI9G
F^GC(\97?/MFbN&ZT@#f/],^CMRBFE@S>UGVNfBIRf&BB[SDS&FH]D;^HeS]L[QH
3J67<@FQGTY-FB(X2W7MEI47=2;^&&6gY##@5_Ra9)NKR[MdLC^UeeeL,KRR(95V
B^6OT8RG6[#d/[:4_?UAZSa+>LZ_7B)S\7QKQ@aQb;#96K8+IOe@dRBd7&?#G#EY
[^:3+CK0Kf\Q4+CZVPRWP&TaSX.6aEDfPL\Q#V6&75.5Y@_=;07A4D9a8T(WZFXG
B(C1)96EH)/;1?W+5(7X<N5../eP<ZM+eBB<8DCX,0K65^NXHN;B]W9#^GWUINgN
<\@-XC.:0f9V2=e36I&9S#1]##MQHEbCSOK[JWAMQG_JdEf1Qg9-34K:;M=PXQXR
IJQ_KZ1Q-3H9>QT1c7)=+-;N^#6P2/VMAg<Jd\gV5YgQXL@^PYB.VaC/<PR9X/E:
WQ>1Pd6IM?bY4cB1(JD<T.-97SYfEd9QY-+YT<e3D),=]K;11_?,KI=SZE0IJ#c_
[?RA;Q>52D7e@N7/\ACgG]SDB^=,6<]ZWD=:4#=B>Se\/\BFW2-DD&K>G+7#F2(e
EGacI3.(YF^Ed5E:QN@9_,b-)MG1f=8W>K8a=ag^9]9>fGTP.:8QP&OVfe<PCL7Y
8/9^TWY5J/cZ1NFP:RDTVFDT.ZVWLG8a4+^=f0^0?4HR(Z/VAPY=@TCB5\>W(0[H
V7?YJ(fd/?L6,>@=(E#JHQ\e_a:T0<;dZc7X(YZ0>&JHS_:cNN7>(3_Ha@6@T^+6
)LDNXJY+JH,HbXKR^M1K2RgM-9])H7.59dW+BFBRBO2ZW]G7S-L+f-K-#6A9UJE0
a?[=XQN^YG;=SZOH.4dg^J&e8CJ2;_O52#b4?REMXLB]=\>PGM)&MgVQ^BVX=QK[
5JPHJ>6:H&0&(=T[@Ldf=?>AN04&2A9#29[R>2&cGV4.?9e?.ag+-YL_M?M(J,#?
RGHH[:IO?<X>^@2X):Q>VJa8#?0-;fB:.UG^Z;=;ReKN.T4E6G//5NIU5f7)>Z&a
eOXEdgMO&PXZAW8#dT1FF>.LT94JJ+K-7aTEBTMDQORWK-66[W\:BF_0(AW-;8CP
W5;>QKPGZYY4_YC?;bfC\IeD-FRXb,g+#XJ/9WcIFg6C(D;(UAZ^g8FHSEJ.S]7G
_5:3N7=V>MaD&A-5Q/E/a@)ICb<H2\K8=X9(=b?PH:;6\bE7DCX(OXV]JD+:7HO_
eC7L76eeSeJW47WV(3Md8dY4U[((/=SSNd0++\YdaD]XQ0cC)P2BK,Y@F1UKES6+
N]N2SJ7OO9[FKC8^P0cfW]K)Uf](T09-5E],?R2<<Z\I=JaM-_@V4d4bCGQPWD/H
?7#=_T>5@J1,A(LP&2>@.ZZR_0IA>4O:DG++?)-(ELWSEdS>=;KC3<Lba3T<a&1)
[EOSR+;C=T7>-L>F=T..)3VPAH]GFd1+C4;0Ab&])N\0[))9\8dVT;]FIXYc,V0S
?/bS@_[A:&/.,3M_-J\9(G33NMM;RGA?bVAZGWUOH8:3)g_,F31/(@R<2+7@#K/b
[U\6)@H84e<MP,AIb]fe,^\b;[+\C+W[SEdF]EXQIg78WP&5,PXTH:b\)?K:<\AG
0M_1a=VT0\79?<NSP>C,8gCFBO)-QUG#O_BA;+=F3\TfV\Q=EMEc&J\gRB5S0?O^
WMH7CK_D6YF]9MD;^FOM6Y@N]R7A&[J0X(Gf_BG3(TbM7Q&,(g^2.c7C)>.J>GE&
1)CO3DaK8d1/-7@F]agDU]<:e1_E4K/A+\ZU9Hf^_2,5\=]D[G&UPTZ>cg9=(0VB
@gUQg3M.3I,f:G#a2P]DFIT5C.JD8]cD^0Jd+d9eP5Aa+3gC?A_[dQKMCO2gAVK1
bM064-^Q/G\<T&cX0[>9ef(>@gASA1>.e7(8D&+5&-?KX_/4d>c[[fQQUAN0.CT8
fAU,g[>S>0bfJ-;B6;>3U(8D.H/\cbT#.EN;8>LK7@GDPEbD_JJH6b-<]V4)XBfg
^KJH/Xa=0W_EB9dW-_Ya<d=1/fXg5)LU-d-VO.?=3MZP&]),-][UAa,,cGC>;3^3
(.]_??P\3XO)GA0ce+YMb9.7IaH)FCBF&A4?6T+G7,QOXZX6->eK7<)L1V#c9M4/
PI&T:AS,Y?CFb@:Xf^cC^[N/3Jg18/./#.),e.&9B+gR1H4M0ZCFH._\,LM8/P[/
6=^OB-gWKAPf-1,Me\NT)7c3:JWFgEcKN^I?&JPMgc/^9.X@f[H12^FYb.8JM/2N
A1F-YDFT,9gZ,KTRD>TM]9ZL1:[F:VRG&&84PZ-cb7=<GXfT@/&aNO3PbO;PWG:3
?_N#_+(#HB<Sc=4GG_;/Ic0&9Md9=>2.eD?K/]b06SeV7;8X6B>3<-8R5aE[O-ME
(AM5C@7]JH00(_<-K/+X3JCGZSOF0W8Y.Q1[^QP5]#HZ6>SD#0ZM;JfC4<YFS3E.
e:f&U/#YJE;]DgWX<;CD:?9W9SE,JU/c)6Ta=<f5ET1I?781eB?U_6+>=+Q[)2U-
-(c\e<f6Y:?,HRBIHF-_YS-AWd-3HZ;[1;G\,X8ec[4cDFJWZ:S#QU4R9&7NagL]
0E-YHf49/e[D=-Ua54B0(=^[#1O8.S9I]=08MQV&OYOT5UZ_WT-Bbe/&;V,U80f(
\U(bd,#7XD>&DSY(_QWGK1_:2>F\B?GXE,F08\E?+>;?8766]d[#2;F05Nf4Wd+8
KZ^H@CJK_XH:4aW8Wc3L7:KV/_5=A-5;;d;YX)1(58Hc\:223DVF)><JSO:5I#([
>U\)VMGdA><(#K6TX/(eRR6^>?[gVBHZ4.5\3HOT-L1V0^N?3Y3g<LeHb7KQ&Rgg
<<+7QAM.&Q5cb]4&_]WSDE\K)]d:3=cK1L@+Q4M@@^?0V5C1&,26L-<4dWFX:\AA
1GgU_Y<gL.C^BG/K4(0a,AM2X1>U)C?PN8<M5H^&HGLA;.A;9_NEI8@WcH^3>VNS
]K<EDgg5>f(&1&T)fa,4>H\+462f_Q@XM9#K<^eRg8?R_Lb9<OTMR;f4bZYT5@.N
c>L3a=.1?_0^DFP+[eY.\)81^G0eCJUB/^e55JOHRCV-2].E1+-DA^)c6O67?3,3
H&QJ7B>?4\a#^IU@SYGX0;_RWT6Q8WS,?(\WIW;ae2JHP.b5c4(P<6E=DK=33AD.
?:>0TdV)RRU<PdD.a_cJD0\aV[R_]N]\6D/@:YJY2=;-+[TRZBL8MF4\I)<IVSC6
X\A.,;bG#RT5;//38VLE)^YFc^@Pa;#F.W#B5WCe5A8<H1AHCg,8c[Y9,Dca8>5@
Pb10])f4@&abDML-3/AfH[S<g6gfS.IY,;93[W-K1CRM9-B7>IB&U.1L(N,,9LWR
FOKKUK&[PI,^E(XOQ]=YMU.I.W-JZ]eE;Q,>J)Pe?+G@1]EGOJ0PU25gR\O+]7I<
[=?\52V?]cB:,aAY-0RG9]GAHWPV#Z?UJYWD&HJ?OB&#;8;4B7)_+AXW02eTXbL[
1]Ja-2^aP[[O=59-bFUf^_KJ@G[RA?;cd4E)HaE#M25E.>+NP?PB4cReVe4d[cg1
3=Mde>A/6;G22RR1):NA\UUZg?5:?bIZO)fTLR&KTQ7:/]beK&:V7&-<2?MeN1&V
DMdG[b.I8_8a\+eGZVP+J=bTc,_,fP9+.FL;Z\^YKSCZUL#Y.aJCC.CEfb3<=)/Z
b(4W;0>7T&&3,32QG_Pb7_(gPT<(_?W06MW7M+aBH-SJ;Xe0UP^D_9VCg]?()c8Q
#7g/ON3:AL-#/JOB0WB2@=aXS<f/@LSMA>A\V=E3;-[XeZ?;97Q0=@=4GaOG#V>Y
@U]3.@9JVd.ce)T:UEI<#;?^(,,G(A2&b;c8eF<V.eAJd.NO]+LRg+L)TV2&b@[<
0.X,[]e#8@G-OX@R3Z8)E735M<DH_5:ASP?.D48C9ER@4_+0R>[+I\VFLe9bX.aY
:3._9Vf>/+EP^\<L3R62]&UV-]56bR=Pd#Y93JIe)Y+.PG</:+aB4#X@62(Z(f</
@Jfd]/PNaT3OLDL&FF/^-fR0cgg:>L1)WM5\f4DcDH\+:PaeDWNOM8S[SdA/XLd6
fEZ?OELBc@GH1.Z)MTQ)P0;D/JNEIV4FN;+TKX9:-=KNeOH?TFQ9EH_])0_L+/)]
)&9=;97T(G2e8?4Ne/V#N4G(Ue3c8A]035#[/=<=/Y&gMPMYb#,BJ7PCTTOMB\1=
V4.&d-=H;^<&c/9WHY_\FD7&ae>f=I-b8T;H,;2#M6&YV[5^\Ra5_Q_;ZWSgf:J@
&)K9=\dJ-KH529:\I>f1_KeIUA9-04#3/ZIGHU0\=-9Ve&\?e[+f-S,:fL\eKN-0
0c75(::Hg=a-4F:J6Ifd]A:#gRAZVB<-Te>a5gDSOT])]g?f7?E;8YBZ@DOYTEZg
Ac@X<[SVfe,Y?HR&Y+7VY=G59CCT94e>A:#Ped=@4I7<H\LgUO+8T@Ue<(9<XTf@
WH/U4+7>g/HN88N5#C>E,Q/\T>J#V6WZ<F)e4JD#7=+ZE&I1BTDbNUQJIYP:STcM
].#?[#cC3\37Rf7e5Y=4QTJGQ#1EQ:UMZdIdH/Z5SF(73d[OLdT]1^;T^4#C)FE@
gA8UG@4-4@2c?A5EN4-BXC]A-X+:K\IVI<QGDZFYPE2,=?W@#3AG7+8T[Y.G[5K.
\_X>/]E4()TdKd^&LI#J@3I@YXHV\55W=]b_Zc.&a:C<V+GT[F=ATg08gf9&b+e2
KB3ZL^BcZ)S2H?48L7<F^/4S>CBBg2I<25/J0)Pd;Y+b7ND))4HK9[PPGF^J9ZMf
_]R3=+9GaON,a+K1#^N1eY;/+;1.)25;=bg?QF05RB643#fe>gNB.&0dRd6QBIab
DKB3E;CH5:-AFe9=A(N0e-4J?\LK@36S1(^bF7Lbg+X.I8O]NZ77://&9XCGf16A
LBd/-Z4?2_Q3>V#AE)W4>N:gKOJ@4S<9X/7NX^CNSQ;<__(<&)A1X#<-][3bAF(<
NXI;fc>8@,Y1&L+Z<3I(K;LTTe8f0B5][R4B_?JVBOP.Jc;-0B3WbK^G+1+Y])cS
O_6?W#5JJVW&Kf_0_5C=#2bE6&[6HZ;SBeSBSVb&U;7OZ=\Y95/W4c^4,9g+/AQD
]K[CO[BK012S80c5\<(g&7b,>I(HaXP8V364]5=)/U4UAX8#7\1D\9AG#AKbbc[9
[,[g=1YW.Q5X#L->K_IQ?UDXL[(aX)bO7B(K)@/,A(BGEIU+)\G5A>cJ,Xb[014b
.8JJ<.d[Q_ba7IN,<gR^?M_9gN(F,0GUW9bC52WeW8KF5Nc=?L7_.FAL)1UJ(=2V
BEE1L:(U=aW-,?cPc+D+:)PA<bIK&&]??[cB8=5)4+.TY>:V9?&J]S3>f#1N&+XW
>WM:(QJGI:W4XL,1U2UKbXKE#@MGQE2FD;-c(->L8X[cT02F:f19)U^f\b@NA+^S
_XcT)](@B<+4NRJa.G54)+4L(558_R#Y_V14cf0ZcaXZ3d_a7E#S1&_5:gQ>\TI8
/RRAPe<__CL5NOaWe,3+ZCbH0@NQF=IZNQG2S4FTG[=BLT5I;T<1C6HL9)T)3WT]
7SG-9;+TN?>K-=EY+M)(UDN,=7b-g.EJRKdMIUDa??E=.SKV.ca-Z-[_C:9LB7I5
&H[PJCD#C5E3VJ5RN.()PWNAb5g7a_EN1\=70>f3-2I.:WecB(L@QF0M#J)3]N#U
F8cE=fOX.S5(J4AND=)cgFCI_UBe6XB-]8UEg7fLJU-F<T^>LB3ReH@5D3VAF91J
K[eM6Z>:g7PO1OT)3WOccL1OVTbAbS[Kf(e<^^[7]ZeR.^SGLCf4;EBb?]Y)KLOI
gE/\VMP45KON0YZ)>1V;g=^1bb:0L=0(\9QMIJ#G2JaKPd<]f#ZB5+DOa>==#G>?
4O-[W#;_LKLc7JUI>#1[;)Ab,VcZ7ZQg)4P6_FUEMDUSTAF;?&(IS>Y[4KTd)g/5
&<D&]I\Pd\=0\G-Q,,F7;R9U0^E4U?MeaNNQN3BJ&MB?.THL8Mf\@_Q\O=Z9\KH]
,d.W6(Y)H<HLd[(@65(]&JR]3CWK:^2<>KB7d=<>JWfgA=CDW4D\NLc^g[8HMNd,
N7WPRfLRHOW?:_B-Q+Z8ebfAY]SHJ>b<,T0;dYdXZ-3eM]NdJgJ2@^4@I8=#ASIC
g,_Y#bXXZJCU^#UAG8-@RK^c=FgA:]FB_9+W67\-TQ_#W1aWScNb3S7NX=X\52-]
4N,V.R0(S<bB;G,:-aYWP\gc,_,S?BKZ^-&1d4+T>JQbf^dJZ@U<711(>^8I#_dU
.HDO@.X860S-&F0L6GI^G;GAe#aTHUCK43=./:YSeGM4BANLWH#T<Xc2FR&EV?Oc
cA0E>=fA&#B26VN;BcNQI__#EeXQ:-+YT/F2H+_)3.GeIKSP3_W?Z8/EFHNGT5AL
Q5;,SAR):4_3#^PXPfX<7PQe,VX)2-(M2F)b9TPCAH[A(MF0ZJUEQ/&_XPGQG_S:
=A1J&VDbdJ>-^VHXT>YSc,;G929OC0YQX@_HT4HP&A>E[8SE)ULe\O7_SP>#BGRY
OCSa/4CgPX8(I<d+dIJfVP8#^8\?EfUB^.A>Y6Y?GS,/GJE79d&,,NF)g@(HC?9[
NaZPD\IDAIO.bF,c3]OFYPU.<b^)@5J3SU.)C@-ODTeXE/XIEQU#]1&fAD+^bg0?
3fF+c=G:WC:S-fIN/_]aMd=Q7;__)(2((NZEe0N8GTG/G1\40YT[8TDeCARBY_R&
XDZ^SLc0]6;(F)F<AN(#(A)G)L?8XC\GU<XF[RBV]^N[+RI/A<FCRZ))IBa-DZgX
X[IZ(.37/bLa+)7EQ=)<^QA(eT]UaR46_=T4KGceS_514UA,F1OYa6A]f]1J[2+V
8/<X:NCU#TR^@0C=OC[CILFTMBdE-a]_RY?UUZD7GY8OZPV7Z<)WA#9DGCD&\XLC
\f:I11G#[LNS4ZO2Q_M8ERD=@+<<NebBUO&G3Y:_1W2PT^-6,@VaFFA;:dCXJ[Eb
BIN#67b#2N^=_DL\/Sf92\F<F7dCd?TcT)2[WDDb9#JY[Q\(NIga.K5SVc]F=eb@
bD(QS_g]G-6G,QdF0EB#Zd>E<<AP[@GAZ&7eD/XTKLdV556IK.RF.DH&9Y;e[b8b
(XDDNW\.5QX1B,,e2-Ca]+JO>G+BSf>[A2Y1HD7]-&dA1IMHCRM?ZU=TA282JF&8
c+CDR#Jd\f1&;X77dA4fCG;\9@(7/e>Eb(a9)KLCE^/L(J4&d:8=C)K.3K=HF^ZP
c46E3[Gd>S6/Y^^OBZ[_?ZEWFg<LLc7ZM>YL,44N\g7TUVV,2b.X75#3C-c#M.d#
,Jf_0aE&aNBg<UJBaeEIWIL>L;S(1[:7:X_WXRQ)3HJW?a^?aX+]+SOG2@5>4E&J
a5>MW7X<;Y(NC?e3TVOAKXg[(5=Z@RN;Z,3Sb,CScSb[.(>DJ7UQ]/TOWU?[<b++
[ZHWb+ZP;:RGZPBeOaML3>UHL4?+318f4DFgJ7,EGVPZaG]<;Le/^HP:a^M^6R>2
cC.a-<Q,K</b,a49C5G^9YScV5KE;/[aO_C?58PVD0JdXSe7caIYS2Fc_H,,S&6d
dAI<3?LGbHK4gB1Uf3B.&(TSNe_b^.fKRG-:COM2?I4?(SWf>:A;69VPF.\>c]9V
6e)b)=JM3GHag00+LH^I#O1U@g^ZLFG0+0M>6O9D2/MEf+-#4&\V=aN0)_YM2)J;
#YK:@;-I.OWN(\dEFE7aV9g/0dgQ5D#Z]GTcFA6=32SD>Oa@]7Pe0=X7.g&RbW>?
<@I:8aSQZW@7_&\#g;<D&-CC#OC00RD<f]a5NV?@J0OZ?:TK:X[HW5SNU@W3_=U(
YO=<6/BgL6L7ZE3RG[^d5W4>\Q-&#+#&c,<Z_E>(,/Y9fA]+OTg+@Q)T@^QbGPTQ
e6MENJ^Ka>-=6&bVY<XV5G,XBO/8d@WQD)5/);=DbIPT1LDSb<IGD2^VB^9.fO8[
gN=bW&6/C4F#C\DB]6U).?-<36P\6f<fYU<ZBMB>HZ.QT63U>Z^4ZC5Q7f^Y7</7
[CeQTKC=LB[WF1LB;-,IgQ:;eAU/=WbYA_^V,#L@ba;3NH+UX1eZa;b_a9;_a)><
\^\)-^Q_B7,T[H:R(bTC)bB<@?1EbX)T0_Vee+f]NQ1L8K+gP-^J//b@SVU3R0-T
.]dA1CP=U@KA/XeY(:[c@/@H0>,&)SXWdgXCfTc3FHF)@WO2(b&L-/dKf.?;.?#]
YX.?PUF#)>V3JIbQV__-W+aLLO9.-4-<?\.IbLCMe9B>KbKYSA0<PX8e\L+GJ9C\
.-O\KOT2<^fK7AI)Y4ASS=ZX=RBP;_D_H@-]29:<_TS@Xg88#QR,&]W[Y7J(aQB8
5g>AP0\edg0P&8Jf,&2N=\.=#6IVg62]8[)OFL:6&d5D6\+E+:?RUb77gO\[a_FY
YSU8Z5-#]0QZOHV\8CR004beUNd[:OU(M\A6Gg)?_=7T?0L&)()L_NdJ]W2a=d@W
+aY[Y&3OI.\:SFC_(ZR:LUXI.X_/_>&b;K[NHAUV\]Hc=0g)4><HgO;K/gg=M_N7
6.+@VHJ6,5DCHdTO.])e:-BXQ,,_,]J#1ZdP>L6BTN-O=0PTBNdZ[bEW@HFJd7SR
(Z><109a@3aL@PGJZ9_d5=a>QOdC(U:RO(CfQR;H#,0&GT@YAb03\W8>E(cVRP\c
5Ff4L@<.,EL69]@6.aS6N7&6eOX)V.YK=3&BI.5BHgR6S@9^,54MBd9F#TP?28Sb
;H#\SZF<<M]3,F17OQ)RHZYK,3\\((H.bS=3S6PQ#26VabOFfJ5LC-P//22[4Y]X
0d9G@I=)A3+RN/]4O#Q+W-(_;UC_79,I-[Za_ESb\;SWE:OK:V_SR#J4O0)-WN+#
_^G=V@g06?U66SIC(M(0d-d,0CLO,e+@,B^BTdBc5>gd2:=:T\^<aL&Dd2\97&7@
<1]3Md??aUK:O@MF:IB=6W1Wg8G0V;Rd9-<9>G\3bbTQ-Cb>ccH;dJ9O56G[#O44
-14[R)K4^gILHQe2[+AN)X;Rb>#bg:#VQ3Ua7Z/1;PX&8D.@&Y8;;3OTQL#5@DL\
K/YH)N-M/R4PgcTZe?GHNe=S3HHTAZe;AE_(/gV^,UD@HbAY4=9a+R9fKO.:>KZ-
:BS21XUD-9CcgU?B101G45K]NCTR2C3gT^U\OR86]X6b=b:c8eWfT<KW<+//b>3]
UCWT&(GT3DG;Y-?M_7a;=4+OLBD3L.ZPZFV]N9gHcD@9_A04BC[E.>;_g9a)UXX+
KH.1-_\/&aV9HA2BN9/KN&GR5SL&,:()gI2J4?5),ER9UP3dUL^b>=.g:aKRZ]@-
AB>D26+G8HEY_;X.OFS4Q&E@_:;T,+<^dNf@#?UfU?PIF#W-&0cRA&U5NH3Y/#_6
P)EYISK1]c-4e@=e0\;,4]_@T,YJ)H4UI#SN[fGb?)g(g1@+,G]81aT^-6K8EC9a
67I+L4\dF)W].W(:CeR;--]gZ6S,PU#Me)1J2c<+be:P2RY2[aVG\PR@I,XCeIX@
0HDNa/(LAT0TA<CK1T^)T\@(D6:ZGR^bFeLH>[TaK3OUIgD:.GURNA8W<O4I_QO3
D8V+NJ-BXd(795@PHJA.A>H&a1@6=)<\#6/)E7GUKb-dLKdKKe,UYM^,J_aOQ+4N
5LgR=6A)QSd1FC[9FP4OX;@X1?f7M:FB3=dOJQ=dVREdQf<1@<EOIUXVUEY8.DUU
.]VMF.c?;CKTKZ80<+)>AW(/(_,gg-F\)-#GOCTI?:6_0_KVQf3\NB2C+10,UITL
Hcf9^[[#,;Q@]UXH2AIeALG-f@UG-.3[_gO8?d/FE.ZWe8V^+YC91V9)/W\eEXMV
V2P.Ace#R7P@R1UbM]-JK^P54c)af(M5+EZ+.]-/<52//-(Y/BL[CUN=M=aJe/SH
e3I_L:dT>IKcfOUeBI^c)R2@H1f3C<BW]17-/36L/CFV1GV#T_](Hd^;b#BDfT^_
6APC0MPA?Yf,C1:<L7GKfMS<\J_TABfZ:A7G332+IOgRbBZR.-Zd62,U?)><BRWG
TJ@W-O6/eY-0U.c@1e#PcKYZ2BUCI#4SE<&@MVUCO##NJ+<^T_NP:J(S/3JU0DPC
e29IEf?-g=\Y^+:Mgd6@2UY?0RVR#CM]7&[#3b0^_B4@6VKU)T@Y6ECA8D>JZMDe
Zd(S60)R-K_g-\eZdTA5T=:/B/AaEV;^5fBTSfX>7N[-XVf3._Z&KYHcAW)dB19\
R[N[#_bAR-edQ0)WBgg-CZLX9N6cT5&-e.8X3@>Eg)\_I;,0.@HPT&HH><T0Vb3S
K+S>34a(FQb1)-daT>-<^(]FY>4YNJ#E,CW&<A9CBWbT\K6;6:dGDJU0:/K9(^LF
JM_378J12-b1+A#_<dEaIYC1Q8NAJ05\;f0L&Rb?[S/B]H\-5.8;66V:)cg2SKRN
bPd)O\C[BJ4SYIU)NZcc#I\6\3a^=OgB6[bbf\7HB)ZM\<a_#=6MI[L@VAN4A52\
M^W/531VLDHV6N<]@8MU\aZB4.UK&[/]eY1]ULZZU<P5GT3Y0,I+>MIb[GOPV:4F
NT?W\_W5gCG0>P0]5XE]C=\_2?e8J&:UH+ALD0FaKGTaY:&OS<Q9@;+W?,0d.J>1
11f)(<A#a[H(QdSZbW6AES3VQHC3cFR[]QX]D\RaaC;PJK>QgS&YA3\D^XZ\a,A7
6gP#&];CSJ51g)_eaFf+S4))&e1N+J__UAW69N&IGe88bJ;=6>B(cAUd<J#Y9<CQ
:J8S5_[IMMGbBREUSJI]HHF?=9+bP?VN]AUM:gB)1)BQE>&ZA7]V_83.3[ZD,8Z5
MR@bf(G^[NMTIR9+#_@+<@Ae)IZJA05[aJKQ[\UNTaLC60D1[[GS[?Q&bdga9?Lc
EY;F/O1K4)-@U?4B:V)D6C/YccRe8O]8OMFLZOEXH&U_JMQT]/_[0LCa[b&,>6D3
f:BDI4Y4&,2;G.[3Z&(UZ1E758;>+PL4^G<8:IEgBT;VZ5ALG/_#Y40b(,A(=[^,
1I6QG+c^ZKF:XPRZf_NbN:E4P@1KEE1d#DM[X^(g7:V1YR[1;gO/P,Eb.)]Yd__Z
)[d0Z79<U8MEgfg;J7G=Z8U_9#GRKU1D34(@O9&TA/#>YT_N4I5\Vec@8ID;SX\3
:X]B^=62FFXECFE=5c:54VRc>&VHZEI.X.Ve)fd#QVfJ++cDIa[)FdKNR<0>9);4
IP4Y@VK;O,fEDKbY9B@0gMB4P1cTFUc^YYaRP(f2g>0]+fZJJI\TJEc&9_-9TL)>
Hd3C9@QY9ZA6b.B/LLNQ(U.CdI2:XNE:b2.QSOJ3)S=;DBDe6W;-79A)J&.4>We3
Zb_ecC9KKe<GYLC:gXF9YZ<c-7T]^Hb/f_E7)73HUBag,<f0EUU\@&V0NbGO#<U[
R#U;>/+_IUV>FEAO.[e8^g/+6eQ2fSf/F676?8607174U,XS4Q:)A]dN8:&I\H<?
-<6,fSe876]7A1^e]>[Dd>.@+^5cD>:PHAJLA-;f<?59U<1[J@.IcO<NFfH+d\Q6
/^I#d4B7A24NJO?0L==@N;d)3/_C4eSG13@2#@bHY7N^JBV6CVf2M2A4I\EQ5]fX
3IaX0.CWA39U0ZWO]?DL)f@:O>#C/+fV(Bc/T)02DJg)(,#]4AaUN@1R0+bbB-)K
88eVD@3FNV_AW/=&BBP_<UI64=5<)B+/48VK33ABHVT#KY]4=N<]gL6103D#98LB
A#C)L@6X_.Cd=SH89,;]:W.]I3T[Yc]9:0M)B03>B_CCH?N&+5]/a@Ic1Z?#7^Vf
NM<6)[deeIK[MA8:)O,<Ta9/aB&F[#]5CAeGH9X9fF#A0[JIa50SPC<ed#;2c5\-
;[\<<D]JR-VRZPZS[CPALRAF3fP08ege[4-OX0K#0<2ZWb.#2_Qf]&#Hb9ID>OL[
)NER<-7HcbYS:f3-+d51G[V/SE4Ge^5L+)TU#S4JW7Z4VP#@)G/?2E,EJ97G:bE1
S_SCZI>^7BR,>E-8cKDHU;KaC=PDN<_\2)(L.bI37H([ZK7JPVd7?fYC&geC5U@U
H^=7IMT]V^OM/CUM+eH9>&]f(3R0\c0:KaJGdG_?cB#DS.0Z3,a9?EES?7GG:/@T
g#V-P^)=YN;W#[Z#PW8:=@W@BV#V:Qc:]Pg?[>0?gI8Q+g3-B21Xc=;UT#4SZ0X.
B16NBA03eH6N.;,ZU;4RRYe5,+IW.<?KI<fY6Ta/WE5A[4Bd#MNDXRaCbU]cW@ZW
aQQg]#Qa;.H(/.;F3S=]d#bV43^4GWJUL^(#=XRM#@\JOV/J)>ZBCBd_#cN2OK>^
C:J>Z=GSb552L;W]c:IUSU@IY;e<9b(?WAP:ASP/ATDH^f=D:D1W<6[5&P3gIIbA
4+;IN,M)@[FY6QDGFQbA@@YCDF#B7)Z\\)Faa#K9S@dCTIE;FXfJZYfK&7WA;?L\
TH]d5)b@[:X;e3;[)0704+/(<[0eSI3(7f20I-Q5d.KQ(:O)8YIC?M?<0eYY(5-G
7?//O,QJTeH8fbH9MLOK<)FQ6&NMDCHSVJBBJgAU?MEP&#-fA+.bS?,+3LGB&<X(
fZBD:[JGLOA)^C>DO;/<+4Y@-LQWX1^1S8HL4bOS-P>7:_@Z]VR48f9dd+5gbSHP
B(MDD.c1-BOfLKF,7>_Bf6,1@#0@9KJ)H+CbLJV-fNM_;V\M+;b_KSfaG&TKLOW^
64<=aO2?[K+O+<G:_G.;?dFF_7gQ?W5gU@SU(CCgMB@;XH+O\X.XBDcKTdKMPeZ4
3^<6Jda.\gYIbReOHRH&Z8<)J6J3&SAJ@dTISEF8=M^IU0FW5FPNG8Wc=C/g6@Ne
=g4/ZU&/C_7,(.1cfK-6F_,VS([1:cKE53E7W\W_?+a@BI[aF-\26P&KL<=^G:Te
6&&:144,<5U,b(dG^+4a)?3b\89RW9O&aLRHd(,CJV1D>5:<a+/ggR.LaY/.+LVK
:FW/>ZbX1RfX5@E-.=OF=5/D=T=\C+79]6W@]WG10LEg2=e=3L\UKF6=fH9?,N@Z
9&Dg?<^UK<6G51<+::V1NC&HQ_4L;7C4O6a#LXY:52b/eB)5?b<Fc6<#bZ8O?1?V
\;J1GH5TcaA;7cZLA+e]ad.RB())_W;]=Y&dT-gId-7c:c;-E;9EDK\H#OZ@WE#&
W(fU^B-D2GTL:0SH,@9eY>T1MH<#SQgQ[b:YOcT)aHaC3^ceReOP<.\VK<c?W9:8
cQ3&264:QV(A.F@.NUN966X@)Z<SFMTd+2?bZ@PM)-[c]99CO4E-+Za_a:Je(_gY
=WBMNPK<_9a)S2&JF\[MKg<cDM<.dI&gA[\?g3G21XP11\a)LcIaUc)X[:<G/Cc[
GUA_R]H&Y6TK.>-^d;2YGgFZ+QU-CbZ9\7?MEVSGI9#9MUNK^>?3\KNRO>J/geY2
3fRNHY_Z_H,OGQ<HDgN(4^aSN;JMTKIe);,;=\@:>782g4#d.(9F>1_;H(gIEV:_
XAB_02Z4L#gT)U)XdR\_P0d,CO:JO;EEe]=dA41ATa2A7-L0A[8eT/=1C)aEB1a.
</^KD@_>0VJFS,df7?+UUH70ZHV0V9?#,9(388VJ3KIa)^A]b+G/)[[C,bTY7?GA
[;7+<X8VTcNN&C:X_6X@:Pg&9S^GTUSePGP?B7I]7-dN+C24(C/=[Z<6_Q,Tf<b&
JEHcRRDFA5cTAT_Lga;\K1IWBH4(K2;7WVYaRNNF5R)?N^H]GW+Q8??.?.7TS>R]
U/g>fc4adD[SLbGG7+/_KH0H../AS+D;Xag)d6AM)<QB^.R&8.GGA>&,[WL1?Xa.
]AAfUb=d_:Q)C\U2D:d;C]@2@RVeU1fB=<=1b7Db0K&3+bFc#-8&T(Nc@(S-55+M
5d7F\B#-+G1da<0.Sg_)T5Ca+C=T,g4P08^VD-W3>8W3#<E+6-[A2IbG1/L?S)((
&:B)R:PXXFJ:bG92aK4:)+=[\JXCY)TM36,&geX]bA?BWI7BeCBX[Fd,g=D?,=\D
CAW8YQT0BU4/)F,c5S3&?B[;<L/H\V9]2XIf--C.<<(dBX7)P_P/4)XBL\M?\>V9
a>[)XX)/Ye6bHOTdTD/UT,[bAa5,0?e@Rc+_b7GL\=.bMAWGaCHQLNHV).M0bM]1
.,W]^:B(.[8NIJV#\(4]LC:;8#;J:].).GPP=)4HJ4aKG4NH?6A#I14M1_I<>9/(
^/4120K]R>ReL1XKZJgI9[.03A>f4NX8_6AF)(1[A?<03T1f@CZ?JT.-<e=&=?DB
fOcROTTQ_FU:MF_T32f@K1^Y\QW.P7U4>LVT+7Jc-(cg(TSf-DIU\AM(WKL1^Ee<
_9=QHeW9PAOY58eRR8Lf9VSR]e?Yc>P;Jg.&/=W.,WA8MMH8[^=QPA>6e.\.;<O(
=_@;C^c;M+Ce[^>&Je#-MH/Q5,Y])W#DLXcVE4U-2(,>aL1b5E\(bH&H/(.]01-c
#WC+AW.00Kfbe(ZSe.:C39GJ^(_3WWF#>;MB10Vb[7L@.;cV4a](TL^5efQ\\4[S
-/B^K?TVK;;(91NI^W)Q0DRJV(:X=?<T<?feT):DcYGDU&/dIMf/ELR20<HCERaF
F+Vg^7Bd\/65D;W\S[<=dVOOG-Z8&U@ae6a4+>e]2f5DT\D8V>IM\9#]9(cA,@M4
ZR[/UI=.KaFb1]N5YbJV=7G(GL^JLBa./67ZO+RM4+@BT6aCFJT@f+TEF>NC\R_Z
IRXA\P9ST=^_Sa^9b4:c#VFAeWVDQf]2CcN=FQT6e3ZG,=B>b5,QbV74;9a.bXQR
>86DV;SZ?dN56GCQe\PS:@]7>#dPX4^\g-E17gDCID/CZ;7=LW)5JOHX0aWO=EBe
3=ZG)JYdE7e1Jf3QbI(<<3Q>#,>G6G3T<9LN<:6A<Ae&5@(bHO^P@O3H#4P3_,Jc
^B>06:#VgdRB)4MAP]4Za[>^fD<[SBaAb.=gd&REbX6b=^e=&3WYM^Jg?Q2)QJ.3
0DUBLSI9C9(LJb_P5VON)][JK\)gGa_IG[QNYFIbAEL^,\.gS^[R#BGC4c\#dJL^
fPF04]]a[5,E=5:STH@50[AN0>FBL_)7,geGPGA5UWUID4)<.+;UGVd(OVVXA=^6
D#G?W?B57-0eGR&Y?K9&b,U@f<DeR\VM+bCZg#89.V)N1+7N1B5222>OD-(WI_dK
EfYaEFfRfeE<YL7KCQ+E(?#:8PdH@4NA^T+U:@I61W3f@F#B#DceTKCb\<Ob#V8L
@RZQR3(<T1,YF)Z?\JG5CJ]3FVGL=MZ\O^H7[0:[)SDYfI>3Yg8.bO[JCd3W+Z9T
Vg+KJ8@J0Ka3P/WNF\IA5d->,>/L]DP_]TWJ?5625Z)\96+I7?baNa,-e.b=00B;
_5QJ&4:0MP;-6F8J&b<8dfBV9?X7HIH#g+6^8e^),<\^\UTb]IBB<N.Q7<72M:.B
0Yd/5L>8L4e1&eDFVK5H8aPWTV5Sf+_9VY?+P5CafQCAH,MF]Y--eAcI8\J[:2eM
]&g.X^GEMbI=FbNXIWF1(&JZ>N,<]PcT>DR:_6TS^/:[]8-Rc_LEEVW@/8fZ4@Nc
CGYI;FcQF66cN>75a/ALTE1=b&PeA3Y/AU)+-KXFGH17+WI70fWe0Ge>6@3VO#fe
e;W[RB?#,?JDN2Hg<R(f-\Z3Cc_7N&b2DS3eK2KcQ>1d+L\D2BagD<1(8E/1\:+.
\E^YL9A=YU+;G6E=0If<N5C&e)3e]aW9V@98I:0:eb].#<;FeSB>2a6[UgOU1W=U
Z&D9U&H7_(WT3GY494Pa?cWI1f;fS\dV)_<I,27ad3#-cTH,CTW=S/W(F8D?5-NZ
Y+[+]Y0Jfe,<AAaG^,K;@^^ea+WB>/e#W4IcO6ACJAMAa7]AP(ID+R&>Y]N(<#R[
.02NY96V<RQ;JYD2,D8ZP85B3VAHM\+;6GI>K=)8IK\24(Y#=a1f7V[U2^AAXEF6
1KE(Z#2V,-/4P+5ecU4eATU/a[Y@8GV^R+1;(#Z<0Y8D_B_6XfKf9H7(#U/R^LaH
2[F>B.&YUYJKI-=Af&g;QPJ5JDUBPH1Ra^MY803)Hb1dX9Z6<20-EIJ5QeE.#BH6
?B,1NN3]8&S1)IKHfXQ4D]Mg:)>UQ^NM??3_QLeD[3cOO5,Z)\CRd8A@(2FAA5bM
N9RYdg@3(CX#dZZ3N&=A@._W-;46+M#A0ELT?:]&E:C<&Q>+gHgbW+#[M(@#c6UT
Uf7DdW?2efR2(^U(=5W3TPA_S+N&QXW?^[[.F:FdfS\/ZgY8W>XS1cC<Ae;eNRa[
\&F?</fW6dIfSD?Y@_I1HJFU>D]5NJY3(4/5<#(JLaWQ1-KLH-SQ>[#M?MLA\b.#
CDL=Td]5:>WTI+Z/R(;g><LZIF067:d(W9eCI.K,-8ZS^cY4(VEECDBAFW,RKgLO
HDVg(QS.0eeFSY19W/I<Z)]ZSZ\CKS\GHLe>:PTFF)+gU)^[_f2e;6QT+Z7=G>U0
/01P(BaXK39L0SFgV^a;)C[?,.IGA#e+>]S=]])W<PMNU;NVGG^-f.R\@NK/.TSS
=0FB.76acJU3LT(1L(R&1/B&&+2#.H1NG@aVe.\^5HJ=^e<U\MIfY#@M?,9Z.bV?
Ic=M.1K_RJY,a<]AN#<<8SX\R(gcC?R2314D4LOCC3McB?W9NF[U+?_?HcL2[0?P
HT36]I^6K#bcfJI,]RI_S3BV8/.\+:(MX]C?W5=2G6[FN#B[.T^-bbd6dX0[[c:/
E<90V,W-9ZE4Kf],2,8?GPHS-1Sd4\f5;:M05_+C3ce_KQ1.C]Ee+Z/g0DNaPT[b
[[P&50.W.H3cfJFFRK5WWVW56dP2PL?[^d.E7==&N=7=ZS87XEYS_Ra6P(cS:KXa
(GcBV-UN)SDMdHJ1VP=P=;eX(<2@>:fHXf>61=GS96/OEZ@1^E3RE9.#N,eWL=Ye
2;AR[Ud.,@Y;aMA?Eb<2?\2<@?\3IPgYe)J+6DB1_2R6\NLU>HWT7J\ffKM^4b,1
0M2+4a,B-.8RMMVM;dX1U6BU(CL\NDCZ<-S64P>UbJ\0=I>dSE>Q9969C3H#\aT?
NARR](/[\d<,_Lb:E>3Hf4+0(gVTBM8;SIf>b4ZOe<O30X]+eAA4XWd&/dQ;),^,
4OJQ59c9/XZWeT]R-74\8&g?BR,Xa0A[(I02>WHHM+d#JeX\:ZgdR.KGL-2:f0[G
;@GZ;QKaEP^JFISF#,-ODF4M\4&R3WF?[7].U];@S;W^/@+0B8\3Oaf3;Z^P;?d:
DJZWfOE,Jc)2ZR,Bd1/g=2I4H,1ICIFZZeNVV?TeP=3?e&-E;-VE1.I0Q_fQID_f
,PFWZ566eK(<c]GXL]E0H]H+@,Xg<fHT4)3_4fN[,(^PGe&Gg\E\gJN&7KL<+7d=
A1aEe157SLG?,/g(;/a=XgW<2X&LQ/XFc^0DDc?@b@ZK,V#CH_6A3:WL-.#Ta&e)
=WeOJ1X+6f@d=fR9&VZRGaAR^[ULH-9E^>>f#==(IS5B0JV:c,dFC_]YN^>JCZ[.
;)B5bQ?b(Y?LZE5NAE-SD6=YF8?+5fA0aVO+eg(>O]BIHfY]Je@QE-KH)HJ179[U
;K7MC,?>^d[_ag]R<4V,^H_S<<]PSa-)fe/<HDc(>[(I?Z?FKD3_28fQ?+,3,5GM
CCYQ\>MEOeCXb,24.fEL._W+C)@13ZW0:/ZHGR>R:G4W(E1VRRF3?X<4V,R]gaC4
X)Q)DbX/AT+^-7Z4==QB2-#[-)4QY+[A<3N>1GPE;8@;A]EEdH@)dI&DGJ1ZK0H5
A7UdOU=,EJHfTL4+AY)(-@?SfBU&EU+E8U9/+B+U@>;\YY9M<ZdKcVP]45RCYSO4
@aLS9R+eZJG8c0>M)SJE)ZP](Ea[FE89FVe[#U)D34gAE@daH^:6^ZW\TAL6\5?T
X2VPHXc))S(N+d0eJZ?GX0YHEMDNf;a3I=MJ:YM17MJFMGgKMQ3(0dB7XN0[gcUB
/+AOSVIVF9G3>(+RONZF0T[>#dL?FV]66MB:&=A<2cXK5Y&PbEC5RO-.V5:&Q2R7
A4?NJ?HI@FGcR/C:f8@^OV@DR(P_R_OG\1OE:&eebHI]F>T94584,aDO4E/I2.TI
O70N:+@I,N^AK3BBH1P/4U?H/gL,@V9;8=R1K+9S8QaM&_Q_Xec;.\_H+>A1W?-4
>?e.#+dLJ#1^HOa5BL(e7eW#fg(@-^ZH4],E:XW9?)>_dJ8IG(<YSAU[[S+N;J9;
?S#fF@4-7(;9+5D,T+(2f7U8]0H/0(C\4:W3V]:_9[/Zg?XZ1Y9II>cLKKZX@=1M
I0DAY6PGZ03,2TIR#UG-5XU;VXe2SgP)N.0,2b>Y66)JN7/+>4MN&dZQC^e41d^W
,aeOM=]Kf65S#GWW.)L8XTJ@7a3+dYV=TdZAeW5Z6FD:5MV#@6K00N\;]=Q?gNUe
C55@M^V--#T]/D8^YT_:&O_Q1UR<B^(HHK_Zfb<^)39@cg_D7dHY4:V+M_+QK^L,
>_4#bbTFHSJOeMNTR^M^P=Z[)BXJ#5/Qc&76^,(TXfPd<J81Vb,].;(E-6-fQ=13
8FF\Af+<-_(cWPc#O^@H_BJG9+_<OT=f^O(4F6K6dPO;AK(P<TFNBAd+?BD&7-#Y
]#.YE@IPM]6XcFXOP]4//bX?Z(;<UQAb0BH16@0)],?IH8;bUYQPP-dYF@VY,\6=
aZ+)3DJB9^UT^XDE882.=U8:_G]KHeRO9R/UHNWQSPg\e^XYc;4dR0MPeQ,9.2+V
(ZA/[TZ>+&2ZMcg#ad<&R]+dUJV9IL3SOA73^7/(2D>4;SR=JD5&K\b];Y4[+Pa>
/04V&=3gAY60CS.#J.7Hg==>?@(6\;Sd=V[]M.XKN-@+3W_RH8b)+Q>&[0,HZPC4
N:)&,>G]Q#J&>25>.O]U&5#U=_MFQ\FcaN>2XLU.Y15;DG9_F+51FW<BG+>dGB]b
IE1)S2HVZ_(GLXNQ@2=EL7dMC33&XH-aU-2>]Y))KZ#]bW[YJUUH1105/;_^,TX#
ZT/K;<P-;0<1O8<dKK/.CA[)DSL6d6dWA#gPX00G25Z\B?J<K4?d-70;T3NC;YU-
&F<DGHDL]N3C@<O8:AW[eR3R[&>.7c+Nb_1aUBE0>580JU^UTD-??(8JR_<e(WHF
ZWFYM#N66K?Q1\<F[VA#GJWQZS(Z&4BLb6A@Ca0@:]=_WQbG0P8Vc7)V_f,8NMK#
C&Bb#ATKAO^TZM;DLY0Q(gSZF@FeYYQ]b?DJX?H8_HW7>_ATFc^dPM98UE1A,=-7
6S3C(JN;[JbOYa+6)<(65^^O]_;Q,000@#a7>UgQdDCZ43+\^,=]61RcgD9?)[QJ
?]31=\BSNBP]\?5?acD7+g.)(8?Y5,8BOQbGHW7_BP]+RC.<:B4g<WSY5F;@ca=[
2E[?C4N[Z7Y&OPT)51/:G0PNMF&1CWN^Q:f2HWaHPS=2:I3Zc\=6#UUZg-][4Og(
H2L^.,+NRKaPIYUB6.f,5-1N2bfPLPL9Yfg,QKQXXeTT/c6=+4)TZ;+a9SB[Cf-W
GHZ-2-gW?d4YD\=6ge,Q9^.64.bJ:2Y4@VeF_0<S-]289Nd;H(@A_&0.16K(9Y0T
=W40B5\.fATQD?KB<g8c11K_[&;POD@5f.8;QAWMZYXgL2:Q;a71?YPC1-CfD2[6
dA(fEK\Fc<3DBF@@U&E9&N,#(=#?\B]fRFaQO/MM_^dD]D3:d&3cYeA0f-JF+c2\
STT[Q+AD1G4R-Q\PH.TA(Q8TM7b=K12&8BUC?YTM(845VP:.4TUb-gYAF@M\GYE_
/3aZY:]b?EbUb#X<8bed/(NAQfAK\FJXLN,5fU^=E5LIYJK++3OMHa[^5=ZdEWcL
.a>KVd-L3>DW&2[CQ3\)F>#4(7d\e(VYdcI)(@8aT,(IMHOb&ULN4&cOb>GM30e=
8^.(7<NdA-Ce]64@J;,VC<7RW=34=59,XIb,Z>NZ+=(,/BdYg3\@4DX0@L]FT;.2
;58P0(0[.EL7Af[BU@LNCTN-25]NP4-@F)b[1&+4B8JK2=&c0)\1JNQ0^Y<EaI4Y
3Q#:6@Y9ZffO2GeG>eH@BAACKbC#P&G7=:QDV.2?HQ-/,^?><3L&V,)^Yc(3.T4d
@c0QFM_^.7P5Cg,aV]Zc1f07W+\De^51;.N5gXR=d_;0RQJ9?&,<7d>AC1.U+2?<
(\-/e1LF.WL<P-9;OM.a<=OdEJXY2BD_,_fcT4=PYH&_f961(H90g?STEO4ZP]CC
c.X]63CQGGR#L4W:><K4+E8ZU1b_/5]_dCZJ[5[f48.BW;Ub?fcD;a<\MOIZH:2\
]=1ee[U6(E,(<dI(Sb(S-e(SS/.(/&5MGT)+=gSN,a&VWMCbcH@Y8(V_[5M99+LK
7,JbY59;)TF#ge.bSFH[ZJ)S)SM>KXK04g6-L#1QFS\UV/EL#RUB99QA:235,1Z0
LWG^&#XIWc9X1>P<)g\NUe[CL\G<a<,W-,OfXPG]>=IJ5bF>ENL?\O0@,,6XCN#_
6GG=&RQDZ\Y:9C;Gf<eTSeC#eP?Sa>@6KNFMd1UbJ9HVdAD91VBF8gg:=CD+<D^D
=YOb^N4YP_^HRMPbM^dJ^/X..&7@&aJDf<<0Ta:VG=+5]<=/Xf5,^&&WNK,?c0LL
;]8]XcWN#BX489KI?RB1KFLDSSRdLDDd+Q[b-JBPgGERg>F<fg(-QGJ6(=\L@1(T
77[UbMTZ@I3Ua5V;T_TAD-W><6B4Z6A[dSC]VJH1f70a@Q[-NEg.N<dZAF2:&&K+
YN1,cTQ&cRV>=)S.4)0/P@LL_72LDWLXWM=I3X.O)>#bO@-[B/6b-82?1KP&]8Q8
2W]QY),V=ge,[5[.]TF6B3e#4\[R>#,a^&^BSQCPM\dRP6.Hd(X#^K=d.g\S/-J>
[Z;G64X]6V[TQA:=NBAGJ0I0eTG>#[U6I_=Z+>&cI:b,H#T.aF0]3SU-1AM\Y(LE
LCO6N+1eb:?5[2XO^@:;cON\M^#W&3D>C6&K[G27EPRCF1HdOcU)_^K(N.;D&1W-
;.g<d3HSJ^00G5<4WPR4(_:,]&]A/X5@@Q.M>IMfVM9cHf@@:GEPT(9Y>aReF0J7
dZ;a@F,I\K9DWCK:#+2G-YG3:1-a/[]&YX-D9f,EX\-/aSZGR\EM@R8/LDO^b@,N
f3IfPFFK&_9_W5.3]1KPRQFIHK@J6OPUcB:OM9((65fE753?/P^e3V+YK<d--8I)
gYHF<MDaGPab8..?Z]07-@A>Fd.D#gLa0J@]O];)QV8<\(WaA]X\KH5Nf4^d^4LJ
#8ON]GRW56./#+Ob/94-2ZUP2U6I9faU<7)1-27fZF0B&3[aO87\5_8&6U:AY0@d
5V=J;TJ0A.a6c<7?,bKMHD5D50<#T;Sb[=OD5<H,J@(=]MZDVcQ6C4b]4LZA7X^G
eP4EHYO>AUE-YTUZ,aLSKN6;]3?E>UMI#cIbb-S]85\gU5g;)O+d?_\Q):QNNDD\
ABf7_QCbSd8B=?(4e64/5bgGM(M2ZW0Lg-.@NK;F.Ab=Y0V>)#&E;ff,fICPE\VK
82;g13P5^K(S[?f9g<:g>#J)DfEYe_YVe5?/g@6QfY.K[4J&1HLUB(R=N]MT?D/F
N<^/>Zgf=?TDN,B=9=fZFKFR/]?/N80OSY5\_1SfOR#JZ,0W>7NCT6:\V9K)2IdS
]+CCK/OU>&2&I]?d4eM@?.19UaU;K1a?Z1IG5S))f>;/T^84?6:F+\g]:_EA/)@>
U6NWS/:]R7fe;5J@g3?H&0EZMddK<87ZVL5/.1.5J2=HLFFSMP4AIB,#;DG4::&-
DEeQU/LZ)d>a?-[H#4MSAXTC78H3>5d_(11-5AcNQ37aAOMEUg.HP&eRELU4SR\I
+Y\G^2U8WGD_Bc@\F=,G\f\-e1DcC=WEY]3;\FX.<>@M;1T[=RS(\D;9.0>(gdXG
G,J.I@B1fR?gWSc5,-)/48W-UENa.-a.+#;UY.bKMYdUeC2c]3+/X#:0(aFOYKCI
FA=[21@1K/^1#gaSdGZRQP#QC(,g_>@5J6^(IbdTMH\&:V>L<BJ@#5YcUeR&HI+N
V=^HSP\4J)e4F?]cJNcOQ#X;VJaP#P/MSfGQ;GKcB6)LBfAX[3UE2?6P2K4=.=[5
HJ3c[>bA]#,LKOAE2aSIQ8=(0)P8.IcMK35N(]M#EOH_79^ZVfBW.Ba_UAX\K>)a
A@B58dBa]>.5ELc(_?IT26.NB8>-eV(P=:T)=QK^_.UMS+@R9[-&g09L+-YV6A2V
&)/>O4ZG(ee4>J^=2VA=^<[H/<Caac/@2D5MH;^+ZAFFP<JfW,9MW:YSACX@c@61
]A=,KdIc<Y,))H--FA@HYf2W]#Y??[>?DN]0DBb734JIB9LfNM.M[2+cH+>[;0:=
e=&2#J8@#QFJKD:=5=4CBB-c;8e:M5#?_)#WZ]\K3E]QSSXe+0OO<cMZFR5Gfd5b
f27+:5L:HC^B964FLLE77Dd&cRCQFS^+3JAE4(Y9AJHg@+L7V1E9:WTRTN-])I4U
==A/J+)X_04P495VRE;b7Tg>RXaLAV_W3Gd3^)a7bXGS(Le0QZ/X59bW&:M7G2d5
_53e<;6#S;EB&3>]J6ag=6@a^XeSFN7GgN(8IeI]O4,f4^4@d[+5X6aA<gb]b@V:
##4=1<R4U7J>8,P]ETKA.[G^e1[86dUScK8I#2RUbGBT8OO/<R_QaDU]FX.^.EVC
MHCZL):7OT5I([Q+V#3G,3>9HE?X<YZcT4<bOO,([Z(B1G>51&V_-^7LY_QdcB7T
_<?@Y:c;eR^RdO7;EEe-[XdXVET?/.Ug)e2b515Se,W74K;U?RVW</c]C]/N@9C>
7K\6[R@FQ?47.5XSEfN2;F6^34I]T+eZK5&O>U5NJA@,QRf(,&2>^HeM+MfZ>W#O
P23CJN?&89_9\^D&GWHI6/CD#]Jff1?P\3Te;a[BA5@0N+I;)#F60Q,_Hd9.WM-.
GaNd60((,_+@7f>G&a-H=<Ia[@SgXAZN.dYNX-42JfUKY@GJD:MW_I393HLXQO;Z
,+XM=eVX?Yf>W4\7L^;K)]f<L4d91+T,&E9W]d+5Wb[8PZ[K>MIg>5P]VNR?>#L(
cBBYL,;Q3\MIPBWJ\X@.V,YG5P>[:HT-,)G:8Z8I:UYbcKgSg8Y;SIH+d,1N8(dR
-R4?X1WJf+cVC_6-K,>PKLRH@M(2+.e&0,UHf2L697Y([@RI(PONHE_4W3c]A9@N
;?2aNCSc78YWXb3c\P#&T]=CM^AGA&0fbgWdRdWCf5+[A0a.BV+f<XaB@YCQE_H8
H5?L7=g1AP3-F:T:E/ZB/8(QQNGQaI6\-)6d<G?LFK1a=?L;)<C/f>eUD8^M((9;
BGf0c202:U61^;[-(NMYF]1gdcNF7F5M4Qe\:B;A<D5fY_82cHLb3+)J.,1AO@S<
<8H#XbE9c)672a<_9a3:gQ[:^DbJXREC;4?EF^G\H4Q=F7&4986H7@=9EW.3M]4(
2O3T4IW606S4:DH+0WfbO#a8Z83:+L5BE4.#(JQG/&(aM(PWbN^^fB_BHg2Wd=.>
Z^;?A]bd5bTSWMN7Y9],:(1MZZV<PL<RU7F4N=-3A\bYIG=RCMCOVgP=eZY^>XZ5
7]W]5]S>S#5/MTMaJ?6Wb<_FcMM&T<DW8OYM-:C8E8T+\/SO^Cc/J>FdBXL4?WYf
A<B\L8J#9/EgeQ3G+_-)fbD--Ve6-(X-KQ]1APC\UV+IN]KffMeM-XT0L:ga;/eI
\IA/733J(YCef--AH/-/J3?7S13N_3d/./Y5g^-__@@O\A_cSd406&e0/f@@+6<(
=\gbC+0=>fVRaD6.PRVXH=OBHc-?c3F5W0FeJ<_.H6(K0\<fU0SAJB;Y.P,J)3,[
B9)5IKM&\@]3]YRV#1].ZAUAC+aa9J44K+71b_Z/[ZI.]>Q3.JeWeSCAL57A0]8a
[b\<HMA#GTK2T7,e37&\6=UZV)&8-PPZ<:LR6B(>F^]EK2+V]PY5P#VV7Me_XKPX
:@d38UF:G+;+QW[:])M+<0^2IGLKBM_5HM^\/+,SC^=-H?8;W^Z#Y9171J2C-WC7
5[MQS^)=#Xc2G&.17W5PFKWESTD/Z5V<P+E7JPdPS::72A)N[X@eN(bI1IWL7bMQ
\@RW>K7Y,<2>(?EG)]_ES\STBa#UFIg_,,S5(\EM:bId[:_=86E:U@&4&DDIDXS(
KDCR_[U3K-IeU(++b(A_5\<ab:;8.-O,4E(cCLgCB@Gb2Qg5cZ?]O3UP]W6)SQS>
V6L7^]N8VB&&<\-JOgJV0:,NQ+Z)NCU12O#@:.TTM.LSWX/g([L.E9K.MY:>#9eG
35@^f]9;<SOR0-#cHHCQ/IEM\E=EUI0>L.HeWb:]&4E#-^e+9JA@9--MKGYcZ/[I
>Q8?UNI))-U#^W)/_/0RV(g)/(S-=C9E?-&5Y=84_#2KR0Xc6U#>)b)L4_./I6)P
)GW6Y&S3):?+,;9SBE22/(g&<&QL=+aL_][V,gS.#X6>J36M\e1ZRJgPgS7OZgY.
WGbHOE6?6GWL5dW_6HDEcI]G0&We#F(EIWRE2JJQSXIL=U;FgK&EL]]7d)7IAb6[
A0GO4\3QeS>TKc95/I5^^B#\J7+@-)cXOM=J^P1a9?DJPXDSK5\DXa]UYQ.DL901
6YQ=1J9>\]Y/(S_=>^1I/X7_B-dUd6/2.H@RGa.a#@<M1Wca2T_^^\&O:Ge?&957
Mc\;?OH&D]]a8+WO^]]IMJFcGV#LN_Z:\V1<CR^KZQ6F8VP=F[)b@YT=,J)](fVH
a>]<MHe45&7:17W7)CK@@B[FN9+_(Y&:[77L,S5E3Je[#9C2/1OC,<619ecC_60Z
GS[E=:^;E/I9]<#-D2M2PD4G0R-Q)[AD:A15YWJUHTW&cDW4F\.NZdW]5W(>)&AL
5XMR;2a569C^;O3Z3aTWD^6CXZ<AQV[B/X4cPSNBWPLL<=;P=B^I1LKOCF4)Mf+X
JXMHPe(<=O^F?),09#[WbLCJgFa7aLY-C>ZB/2P9c@/<O.AW<EOP0,,JV^I=V4@1
](Y&7;=[MHL;B8#MaW#M&-?PJ\-4>?5YV:NZPg:fg6D\RSdbgH):K+>Gc7H^3_Gf
/?21EGN0[>JY]cCYH^(OMYQO;<EDFfA8[(/T6a-]a:8TXcf_e:NH(PT;eU3F.DB5
T4N]\6?c_H0R>.E3]8VFfFCA6HM;DR9ZQWJ_#KS^L:HV]IP#(WMcEN2]Q8O-,?3K
@=0ECb@B73065NR5#H-)GG02<caG\^@f>gg?A\QBHT^dQA9E\@YN)TRgd7G[JM/e
AE18+PS\,a&T,@6L/L_HP#WK);-=E>,XXOFgBM#\_>2<YZe&b<>gZ:(g#^NM^&Y_
2_YM?WBb^@W0aK+(#^W:IG34#Ec\ZTd(07UfC5JPHIFXG4R)EM.g)eE0Y1VAGA;G
&J5KN_)D2E1Cc7QH/FK::Be:W8.Q<:HV4.1U-_\Ne\]@V_DY,EV=1Q29M#3[^;dN
GXW_eSHLPQT7b4069N9UTXE#DOV\6:8_;ZTPPeI8^beF/(EIQ_f-eZN/J;[<?@=E
fFS&V@PaPF=?Lb?B+F=c:OS[BWHZXPK]&?gM[c[MU^L@=/)EAMZ1XN;,D6[TgQ3<
DOH=9FV?^75eYd=)aB-e)IfOdR,B)>a4G&O_],RP#TAS5cHUEV9@G58809/374&\
dEHOL:<MZaWQ?DC4-X6a8YOZ1@AD>K8[<b=0N@OM&IDf,Gf6;H;1d,SbD?F4-29Z
CK07d^>_0JG;:VYG&#N\OZ4J3M[<WBe?e>TW(02=2:b>f\,#((,;/Z4,<]cM//:A
W=BFgQ0=0I,DZ+08^[AcK=29C?((_?IL^H?\^M.&:gYdTB&)FCgK-N:A(<7NT,dW
XN4gX+^O@GYLJ^.V#GZEH7QJeJbgEQ5KE0)<cY3Yd>0_=]CFa^,FDcebVV0@2N9c
.TJ^#?E+,\S?&][)>OT,g[dW00f1MHVM^6G6>Va:[FAD,eV\Lc_(\gITG>?(8_K,
Z1[J_M\a^&6/FJaK]+P+02E/^/E)9HF9&fgKLHC4/J9ILd^c;<U9Ae>A;M@A#7>,
F[3\\77<>IV5f,UQ,^Ha?e7OFPB.@b2X[1c16[V36CAdb:Pd]\R3Tc)1.9OC_AFF
A)?bD]&0YYZ\P+QG96V#FZ=UKL,WS<3>:IbU#2,VPaQ_IAXNEQf[]CQ.[MV57Sa3
85ZVOC:OXW\gZ,J>df3EcP#+1@3#f<?:FSYC?E()?HXCI+\)I</ZeTH+=>@HC0U7
K7@0UgW)H^1YSMHGG(_JK?]f+LD0[e_3VgJ9QLN72@4MZgJPd+0(K\VQ98d>B1@R
^F1<9+7VTP(CPP>AH3H_IMU\ge3D-V.@/1F:bJE;:-Q79cW^G/,eJUZRL<F+K<Hg
VMWXCcZAD(M_.TX7=3Ib)T1_6b&+2W=IC^K9c:;Le&Y)/?4,cII3#(::CR+aJXKZ
9Z6P.DYRN,TKe\^U-#KK17,S?BR_JFTNQ5fR(b^4J=b:P,(H+0>@K-D<<E(5]#[T
b0@GB(X]a3bM3<3Rb2\B8\a?[\>eE<:3(acGQdg[(\^Z^SMc@+^2eW7=25c-(?@_
AJ.\7;L&5[:fE?Y+P:78a.G8X<UEA0Hd<216geD4bFX^Vc1Q\YZ\[2bBfGf,G94L
J<6^;+f+I,ROHW,gdS8GZ,AOL7Rc?e+ST38M)[cALb_L4XDFIY4\M8IL)MC,b;NN
<3Y^d@&B(QS9(X(-,:;0/Z2OOS9=\g22_9X[_(e>@/Q6GJ^D>3aL4P>U<&C\C-ZM
G=PHg/)4LS]O.TU_]VES(QcTC8.>,-;UFTH9];cb@(<@R0V0]g#S:U#Pa7])03@A
b>1NY@?/G3\5^J:6G>[M;TX;ZQ[g1UL464AC[EEI1;X&.D</4G_Ie.e;5=fL3K=J
\RR,c6cb;Z[g1NYc0&5MWI89BQE5T[AHI.X54[ZS0H^7+:1Zf(&W&C4]MG/+HA6=
a]d[S2B>P_-g^JC1[WN@fF7]\7N=AZNPd@H^UXOebC2<AIeTg+H<11fCO>N0XcGQ
5M^;IQ.BZJXTY^6>+e2J;328?PEN#O[&K3)<6.7T-_Ca01bJdGaM)+aW8a)IFc:?
b]:+7OB3Ff;5#b>YdXafF-.T@b,_N)9eb:_E[A9-S-\/M>H4WU]?aWa+H8P<4B(8
AfcL:N/X31&RUXV.5OSgFLdL,bL.HTJD(1c6YccQ]<HNa9<@2=,BUDQ>-Ug5?Lb.
\@XXSQO>C\:=PSgVJPB?YYDR2\E#0.4f:M1L=V9?X.ed2L1Y-7R9T;SKSTNY7_;R
@9^aU^)Ab(W1g.;F[g),#)5SH=Db3Q,M,ZE[NYOb<T[T3.VFcc/?S2SNDUYSK&Kb
W5WW&D9@Zf,G,eVb_8.>KA[23LV>d?-gFfRCNe;bZWIDd&ReX:aDKL2)Qa]Uc@-N
C,((YTJ@VMN@C0_BCQ:7U@Gg[Gc?[68,J?;9=U;JdWA(VX^98&Hc=8DW[W2,(bdY
5b&3@FW7ff:d3+BSbBVG&WBeAZR<b0X91_bJ0I5U?cLgH#OL<[+=Y4bIF&)QPCG]
;]g30Lacd45\(G1KQ1]aG^MA@&L+MB7.YPR9cWQP@deEQ2KFaQ(R/4<^V^E,A6OB
YL4RNV//:SbdC&L3@QdD^(MBDS[MfN<O&<F6:gTU_,g@H,UQ+?:eUg004[-SUNG/
1EcI7MX??N5Z0UJJ4H3X867;L64#Nb=LU1_;8:-50ZX.)Bag,VZ]:I+_XcWY<Z,U
fb[),2PLS+/S<SEQ0V2&)SM1?:BMK(+FBGAdd;)LQY2_WR92<#dI8ZMDRgg&>LS7
e33U.84da\-)FDBA7:Z+JP2-DFMUAG\dR@b;DW@MA-O<)1&Q0QO.2[,(/Vcd=ZM1
VfY.[M2U2Yb;ff^T2@4));,]:d[FHK@bW^@YPV#QRG4B)#/8W)V#KLHb+RYa6:SM
5VK3G80^[<f]W11:<+R->]-Y:JTf+aBT,VLe^OS.c.#4dTZ_^C)\IQGT,STb?_\I
&@7P&Gb>25[U>BD?WUDY_bAOB[gZBG1Ye2:#H6@N#9EI8I.XWY4D<K3ETK=I^2G2
Z>NK(6YQ\YKLB?IGSM21fX.RY2M;bP\5L+DQFKHf+H4UA+E4e]<aICO-(gM4+F,V
0XGRI90SZI[g3Q+XR<T8ZR(.YgcE3/5[=)[G2A;#O8##QM1&EP7HB;Z+E46NG8_M
[54I,D+;4D0/I;?2:a5cLCO#9:=6<,]4fbbCa+B#JD;N.\a-f),V3L^ZUdg1F1Z3
ZcI4E3:/[S&@\YbC:TV+4HZDYCCVe]PF4&=.O7^KORQEU-N==HYaJXZad3c0aRKC
872U?F>-=-8AW6@Z#VH?_E[U+WdRf]/X\aJ;\f?#b6?Z;QOJ<dEUAT#N=a.823&V
g0J->M7RI)_TLcg0.1dM?b](Z><3GUHA7fJ[R,5cQ^OId_N:bLU=Cg.^@WYL2F=5
a\J:O4S4a4)3\+(\2DOac;88QLDL+gG72cB0IN:de:OQV)f8\6)M2?\VL^(TZN@[
cQc9^M]bB__FPFOR)gYU&dd-0+DW6;V>(>\SXWVN<2ITNXc7N3ZVbH7O?,?@&\J2
d[,FU:CS)P6-R@4]=:ND\)\N&[LD=XHWNAIKJaD/d31((\cbNaI=29?@IEMQTUG[
[4RBZQR9Q\<-_9K6V<>)1]eAe47?<;dU-gT;;V0&5a2eWVg);>NP-2HOeBf_Z8QC
\\SaH;7-/3JQ9(cT40<g44<0V2[NP>#&U6b\&;;2?>Me0M.A_XeBXGP<MLdIJ8?B
\H9dWG-d1ZTD^-1P0:gNQNaE8(46b4S;M/e(Pf5WYdL[JO]YNJ;b85)MBg9d&DT6
D_5+ME.UbK9bKBPY>AZ?:.HaO/.03K=\B+(6WBC]088I\?WCb1#BOKU\OX?eSZJ5
C=MMQ;_#?gAacH>K9;Rg<3<\PFc.\]FH\=1bH0cBDU;c8N00;a+<SZ34OPSLE,B#
J=]=XC\g>2=Hc\<N9<@>[VM()_<4QaU]CKZ2/RPUXa22Xdf9-(Q/=,e->dN+#2ZZ
_\V,,I(N[FTM[)-0KUge_,[gF^cAZO5;@64Y<a:.V?=#VT2S>0^fE##FOU/K#6G,
:&O;-.99^b;J,-;&2P=egf]Z/\(Jd[M-[7G)W7B=0&K-\6\;G6UV@[).IRJe#94W
67>AVb-/0gV\MaV)M6[,=f^U,+E^)QRF=]@JH@^&0T\..H1+&XS)38deG50AA?>b
/(;N9L@Z;K/Qf@5fM6L^f#Je(cg8-W]:<UU]@:>^(G^2gDDfD.CKZa/+O=13Mf58
H)=2gN@GSHb5(V/9bUB4O9U,F>[;=ZP9VB]DZT3aM\Dc(BIP+24310B0fVRXV20/
U[-ST197d_N]55F[N;5]33[f_.:0T(L>Mf(7^.dUb00.LTD]BeSg=MLH+E[ZK:T<
0#)<&GM0,F9.=C#a5Z8PL@WH@b9f>S(dJTDB>W11S=d7EW(HL4DZQ-=_1JLf#)@-
&(PGg.bQ+g7cMbKf\S:9.?V15DVVb4;71UT63&0Q>^[+XDVcb.+;KeC](,f&G<FK
_JN&T73B<(e@D.SE[@AP[RdI)_\6Of=70A^b5#2H10a[;N;VHPVH[QSNGJW-J[;@
,)ONJ4)XHIgY9,O3#G93_FE2M>Fd[2>5B_f3_dW<?A9.3&^^EV&6\E-#MM7ZBb3O
X/[0dZR1VHI6<;a>_+]0b9,_XMGXR.+F7f#e-3;?_;.E9(bBQ#3b7542O8f[)77#
8B/26_e>R,@E(KD#f3L9AM\7eTe_OVLgV#L]7GMS?2(_>X=TH&8\N&=YIf8-^8E)
MUQZ]X)GT@3b:5TQ=E[^665.JJOQT4+=R^;KT;TW>ELUGg43?ScO&>#,7c_SHb9;
WZG).+.16&^MKa.\#Ya)N+,D02d(;8LQFcONdX2<P/f69Ha8.AWUgD)PDTLA8EQG
fY4g;E_+KE1K+LT,U>P.T6WaRGV#&GR^59Rd;<824>(GW\Vdf4.AB44^5,+4JES;
&c.fZ31X5C>H&B[GIbP5_S74/9)Z_D#1M9U5.=N,HW01Y)-4WWd7Y=Z<3SM<^SCX
;+dGWc_SQA2[Y\W];ATg[.,43(M#g;12K:P9[(>MMZMU<.A5EXY=,M6C+WC#(aG7
6>F\@)WJ1_:,S)\1F.D6@F_^e-JgAdFWNKedX+M-WPLb)-/S+Mg;F2cKUf37XB:+
0fB&OEe.SAAHgJ/X:5UYOA&g)LFC<Q,aE(3WQ7c\\D.?7b]NBXK_W]^-GIVI2dN&
8PCU7L;>^&UZc:TaZP6ggC+_7@@CUcM&4]P=\N8+RQR5eROg53;>^4K^6F)[864g
[D8-KR^_@X<Ug2O8^[&.b\R>^HCG@P[]@.d[<e8ID,,2O#\YDP6W57X6NQ9BBD)#
G0fSHI/D&F0&0c<O1_&L]JX[]-E7>c19_e2gIV+J;<LTc&N_Z2X_Q<TYOLUA?.)M
3QLED,U&(CP;B\>KUd[Ee62fO3@?&J.2LAC[Ob>/#W61&)ES^UOC2cI,@))63AMc
R]@S/&cVR>9RCf]Zag9:UU<\2MdMR]e:DJ6&=e?L?#^;>8;TU;d=PY@g1bH,S/PW
e^><=<3]+cagcbbe0;JCI6=N4AISJ&,QQ+K68Ee_:RAR:EA7N:ZNDO#0c.RVR6?,
+]VWW#6F]]=_T@Q#7YU3^I&1_(-I3?2DT\?JR6>&HY1Q2O6&.7Zg:AH<481/.92b
HYNM6JZea+\b0eUV)YW4f_\\b,ZdDV-H13A>R65XI:.ZA4f+L96e&4C&G#D&TT^>
&4f1=]3]^5-G/WZJg?[&GcHI\<c<.BSN+1R:2f<fW=R^Q5A0HG0S;UD)=Ab&)VMS
R:<9B(W]007@@^/4Qgd=cDIWT3W\D1M&65L:,^eH.KN>ZT+<+d[Qa)1<<Nd?>S6f
66@@LU;-_-HW1Ha\M-I)GF]QH]LDNM6FK.K=AbTKQY2CVD_1,7NMLdCK6dWR>0Ga
]?V/R\LLK.RCHGJ>1HWd_MM-56N_Y^B-8#ffYc?6/:Zg6g>S)b[@RO;f;5CL&Y6c
24)T(XG4=C;H26gdKe@:_,Q@G;X\?CXK]5e(4WE>&5bg=22HdCccQX9]0RT#fNG2
I)AO8?EQA1#D5QCZbUH:Z3UgANT;+aSK[:1G-_1Q,g5.4V+DDYG4[(0CUg?dC244
1\B8HKO8VbOM77TTCd(]Z]d;6RW=)9VX:24O\(M>[VF;HWFTPX0,&18;9T/D-B+c
27,]R<b7Ide;I^N\0GED;R-S-XX=;DJN6#\@DUOJ:,1(^(J&ZTA_a-^/FYgP5(0.
6>;&^8cO:KNSVFWXC([-G/&MbRc=B/5COOHaV7I9KS(23](6DOV&IR]ZBI#A5Pb:
Ue^YMB(_.?&H4_SY)_VgTQ=<L/3:#=2]((5VH.R(LCc:_REF99Z51Gb:-BKFQ=;8
E^BYBYU07c(&5b,fgG,ICW<&4JfPaT;0_XW+=0+M0CL>A>):/.O@IU6GQ\:9JQ[.
daH#_AXKe=BV&89\-1;BMd\ad[\53]VHL\ZZXXbC.MI3bWgK@FT\T5]P&2._46L?
:]QD?g?/=6;5cF[0-a6[;\ab.,C#GG+OaZV6ED+C0P^<UZ)3e&L9J>;M]NM9MK=4
32HG[O#QQb7]SG7H<Od<;,02KL(-.+.NQH_0B]HC5@L\Jd35a3-2V?JH<<,2,>PM
2]-WfaWK+J39LID4)aafUXDKWB:SXR=?aT?gP?]aP8a)C;NagM.TeGIWg@J9CSSU
=ZIUYHI]Jc2VH[dca25WVa[5U67&M/gR59B(.#<3K]PHV_)6.ZQTD3(,:ZcT+_1]
)9G-/9c+=ZOV_W7.a^#V,Y6?,QS<^b?IYN)?UQ[265&b?]^C.Db0P7NT^X_GDd)]
5;Y.&eUbM.c]X9b?98Y>G]-<JfXZW6F-?F]F)g5OI:HU.DY<Y_@08OO\3aSD#4?D
8_c@5+Iag>7R\]?O([VALBF0],PgNfJI4^5eRX>[M_U#ICY_V]g1&W1RHVJ71]U&
.F6eC\@GN=^6Z3Y3V[L[:+5?e?V8fB8KY>96IBaa0A@:fP.9ZB_I5NX:EM,&Q3D@
Yc.E-R)0_C>I2XA@GL,gd_=C@_@(I1;6RX8?N/::;PUDB23MGWNJAA][A.a]V]:-
g=K0/CPV<UeE?HZ6EHK7eLII<K4&:-&MLB+21#LRY^?I;S)R?GL,D\@eTM^4FO;H
YR#+CR:G7:+9e=N5gC+:Yg?ZSN&dc/LW0b0,-fFKU5<.WKM,/c7=)+#.0U2F0^b,
J(2.E2W)NZF;]&1<bXM@-A485@CJJI-](&II14R&cAV^^?&^2N<DSW9+e>;>2J,H
dGILU@;/^PQ#\Dc52I3KIU\]YbH1:_O1bN4Je7@JVP:-M01KS\I@0b(IGAeQ8J0b
D]\[9DH54]FXZ4[WWOA<-7[K:>WSNDg5@VN^:Ic^@W1-+c##=W)O72Hg>REBY)NA
M_Cc7##&OUE\8Y6\eO=3TNUb9E:BFPMV24/-Y<[:M3[&6VCH2;7A_SR[df.,(SJE
Jg]#926fJJ1X0HMV88?d+ZB@XeA[)B8_Ve47#UJY[[\JY5W^QfFMb(M).-JYV7.E
g.7[P2-#4E/UHSZgRMHM8f1K<1-a:-dY3dF2L>CI&A--1AE[#U6KL&P1)=fEL<:D
C?LbVL;.:)ZT^[c1PO@JHA(FZ^0=G8/))BB?<,W0YN,5)#3&A8_6M]dHQSdB=H0>
E5MDF[g@O??IPWP=CX<f#V>U1H/H@BE:Xdb[,[(YGdN4+#.bY;WE>6a.3.R0UJMK
e=>3FQ)RK(G4DFTZU25=;LN-,QGHU3OUb6TVH.G:\W0a70N#+\/GLJfdfa084(85
CTTBf-95aOM=D7=0:Kc1Z[K7T55VU7TNF0C[#_++B4J#eec.7?#+HUO+d_fNRc.C
DJF&)g1d\Ib:==(7(V\FNg)1S&fX@8S5/7U]0>707f2+>EUSIR1>?8b6YBb7I(I(
Dge:X[QA5/05SJSXOO[\.]Y4];Z8.APa6+2#cQG&>1ICT>:^.>MGGR1TfCI?#V:.
=bB19ce3.Ie\/IIdD.6@]&P.NY0H3\JSWE..BE+IMY:Q0]W2?8I?&+X>R9E3dS+F
W(fSKJUa+.NJ0d+:T<gSL-)VA5g-+4F.JPKX.RD\<<0BS)\]JZGT[@2f[PZdA2?V
[ZJD&+>N+U8ZY7@VC8?\NFP0:.G+-0^RDQXcOHG#.c<R3Cf<:/AFH:<T,(]gTScN
eO[-ZdIIaE-1U]A#JX.0:W]0;(I-D@f8E8>Q>Q2I6[T(^L&(B^1Wd6MG]6TZJO>B
_ARM[3TVg/d4[T3<F>B;-^@CRcXY.K9@4OF>Z(RTdQD.<,XOWGB1Q^O)MC<Bff9?
,61,5d.8L[AEfEEQcf[SADJf1eU1H+U66IJ5VAKBTZI4U,b:bLH_f.ZZ3-EOT+4b
-QO&WJ9]2dfgOK)PRM^[aP19<0+?&<5G_/V)A6fg#J(&@/7bYMd)P09F^#^fZP-0
/e7g5LFbOOV^d1,F5(&FdQ(/e3^7H_\DQ?LK)EESgINSf2(@KD=<C<>@WE.THHMg
D1VXQ#e.eQ>4IWeWDOHYY&3/W_NU(5X<PYA#YCacAYKMXV,<g8BNe]eK(f+IB\b;
T?L#N83:VK_9ce==P(NYPA@1^aL;HU-JV^bR#9===d0[2A7J\+Za/acWIaKHT+A]
g)FA)N078U/I<\YFZUL+>f\gBX1&4P]3.2,0Cg=6)9a)YO1253=:E.6_45K2d@\\
?=H,#Lf1g7:ZQ]()GLeP_#U3<]75K0f+C659,I>--PaMU&=g--W705BCD04G57^R
ZMdJ9f?Dd0-&GSb2L2^.WOH#_RC85dL\PSI\_]R=PBdBTBVFO\1?(^\1YGOIPE<G
Z]F.Ab]P<OcIUUN:YY7RW;9X<-;OS=.T.L-C88##IK69&,:/gWCfeAbHA50,Fe?R
.7,IF[8KGbL7>LI?U>^#)M;K]#E><U&1L/3<>AfgV5Q,@NEP5;L/N0^1_4.V12W0
J^/N:Cc@.T]#ZDG&5/O;FG34#M6:#&Yc7Z-2:S2AI_>;JRY47^>(UfcK1ZLZ+.e-
4C493c8;@F9g<4\<ON1T+4V1GV9\0\=?[#fWS.8&eU8[)+f[cI5d6_P47S.HA7fG
KKIYWD+bL7??Kb.>]P92?LJ+g5e2GNH?Q3?bbQXY.YF-fWP?73>-AeQ/?TVZ-C^D
CU^)^<@Qc3VdIC&c\7@Xd3+<QbTCY3;<f;8>cS.O=ZVYT\8&8@WdCQA=Z3PJ_SP8
873^)1>#@:D4::?YG-AAHWVfc2_)L1e+6f4>A\gBeUSH?&-C73fA00;B])fAF,FW
7Ig&_)+:#T]S#Cd39BL[3OP((6048==M84aF5,LCgR9BXc@dbU)5)3]5U3EV?g(8
a-1d:-)bPf^N.GGcS@a&cfS,[H#@UcUG1eFaW_OL9MIH@NB]ZC;HY-SCHa^D84+;
?2R#]Z#6b#?VOfH?d<eSNB4)WTWQR1_7+E?@]/46:X+_/+[R2f@^4/,(\&HLB=DR
c_#B(V9KR?=bGWD4eZG#,(LB/+,JI7=,Z3,SN(XEg^<)g>Fe^,=N4BDC;Z1MQ>-8
/b3IJPJA.VOE<<9RS#8>f)Ec/W]&=ae13\TY(:8HY84U;aN<?d(#E+T3:V&R_VgH
W08F6g<=^XdU52_<_\ZAZUPW=2Y;UbM<FXLL=GB7A[(1g@<,^PPV+Q?.9eV-0MQC
2L]O#7E=1RH22URN3LNLR(NQ<dMBGTCY2U4#^?GTLFaB\Le?7F^,>?93NdH+&f23
&<E?[a]D4a\:ON/&bJ&(D7D>-I,9#dbOS)?Dc8LU1:[.]H7cLRR4;,BPLBC;89KL
OP>PMH&\f;-[g:N;Sd[L:R,#B50>DI5&IcOXNH(9;;30T?Y9?A,;^aQ_PR=#X1Of
9<@EEdO6GE1^77.Z<XI5:Wf;K?W[1LXQ+bI&6C)VQ[<5R5b<[L1OaRO^9G;5=W:C
T)VQUgcIX;S>V(@b>UA<J_9W#KF<<aK3Ha;?C.E&]/QD/T.9#S?6U:J7G,4J_KZ^
NSG+;OX][f_-eN5g1&7N.G&M92M3<QV=T,B]G^-AGQg<&-af-FR5^?VA]@F=Ma\8
<)&Pcg3.a#(@+g\@SFULaJcd02^gaX^G&HXPPd^87VWaFb/]d]&#K@<4@R>N8fI#
Z34eT8-+S&FYQ>#,8f]RaT][)Wg(6L#^>KO)0]\0BVI(>UKPUJ/D]KM1gALZ-f0^
MUZRQ3:3:>JF<_dCRZW--E(_LfU2]VTQ?5:=)\<DLS)_,_21URA=MU]&XV0eU1L9
@<a#BIOf8KJK?M+_QNa>0-TN#g&\Ge-?^X@OYd]3.D.Z;J+4R)Hc:f[^Y:LQ((5S
A4B+3a>4A-R>77]/N=K(KX(b&^M=QWG&D]U<J5I?#O(4#39\@.:B2U;P-3>NXINF
73GWQ]J6[.JO^c2:fBKNMFQ9[FdU-OXL4VGaV&H&WF):6J<=(gYAIZ0KOI=NFH&\
OQK[]DC)N+Wf#EJMDKP(I6fO>3T,CL9TaW#.^-f-._?)W3DJ@S\6J/I0GM=bOV9c
E_]4I<B8A1^gRZN4eQ9+S[9G4BBSggMYP-=.FM4E^Y=USf?TLH=^P<7X\5Q9Y=:e
@)f\K0Z1[C8(HT>_(CP7)JdLN0e([A&MgNF,b;FZaKdVI6IGK(b\UfF?CM[O&E#6
Gg9gZYeBR,#^[)YB^H9BN9I6U(-&b/2I@-:G9KFJ7:_5CF^dAK;A2&_3FEPMP5P7
bPQ?CF9/@eeTOPJd>c;OU]+8<1.b(5./^ZZ]SX0fV:Gce-8g2>4)9S6E-B[0@L.4
>@),_3+G]@I&M+=;d8>,6GQd/>aFCOEGX^,5[Q\F4IQ/d7[J.]J#3^+TZeg<_05?
#L>7MS6?8Zf-Z6BYa43;..4=;?e-(\)BaP[3Q&+O4B+bES\SK^OAZ(DSWYPd<WWN
K4?2dSR0f>(@P)C+FRMCg-XCN?_J>3(RE0QD#2L/;X,323WDeNSI9+6B/,Z9A138
C&2^bDSQZ)1PNR;B.6Wb.3M6D0^66\(Lg/:<HCaSCXVgDCfN9b78/AO[Y\7O<^/U
XI+@^FCD7@8G+/-a]T@b/a-SK\LGQ&e2Q2WS1+5A&eJ0Tc]gX44CR>]OIC?W#AF]
f=(ZdZB+@07X6DY#WGN.MT]1CT_S(/;D/YaUHOg<EY?Mbf<K:aD>:(W^@A89]6&8
Ma#I@@8R4YPS4>AD[bVaUMM&Ob27-[ZYD,McJIZ&_M9>gV#;9W>JCecE1Z3DZKfJ
OF9M<5L0MN,fb[3f+P5CF4BZBEP:)8PWZf(Wd+&-)M0^)&X(;T4;Pgbb;bc\^OIH
X2EJg@dBLMbT.]c+ge^<=\7KU+\(:-6&Q44=VE<.A92,WF2BS0HXS;CTdH0?g5^Z
d/We4T8_+#SQXc:6;2WbU#J:<NgUFDNUXK.+dFZP;/OPa+BFASH+QYfH]8(UV4K,
8N4-/0_30?1))?3dIb63M?P#5ZfAgQWN[0\\=J;-867]d.BbVYOU26:SM\?BKJ=d
gRZCJM?:,:VISBXKbf17[,f4Id->L\gA>3P^ef<MDaS@Z+F14cLg\aL5-7X1-JM#
<3/(8>)?34fa/gaL@KOf@,WW.=,PU-#4=<]HEN]fQ5+ce^7MeZ(MVIf47D>]K7EF
V:bNe>M0,Z=gZ@TYDgP9^,5CQA]C9CfM.)P5EAG,KN/(91Bb,):Ge__?HVc40dd2
-a;;#>L>=6MS5ASYc<DRM),dGb<:CYfQ8A]d[cD;_BH/^\7bD0R7X0@^=6JdZWEU
R-gQ6RO=6MF)+Z07YRX,1\e)1Hf9cZ3&AM-a&cOM<+1J)]-,9W]dA3,.Kgf9O^B)
6?H<4BI)-C/[3NEM23&.8a(,-^:g.,R5VM>>F+?4J\.@)YGJ5_K-<Q(2eTLaa<0?
ZBc6@eW&R=1C3D1[>NYU4\>5J<HedKBNIK@b8Y?]9e9]D;DJ-,C;=C@4+?T5;T_6
.[ZJU[Dg4J+^33WNaCAeg=,D,76g1(R/G#STX,fFX+.W\Q>9A+7^R[4,.4L^;8)Z
OO1(25(SH9TF&TBgU/Ca0^:1:47XPM#IUd>Sc?(\d6?Of=K.JJ7W39gf=O>aB#R8
EPaZC[YL8Xd;K4<1GUUHWbafa@&PGddP#LcdK8U2M;&/Hc:2\<NBLK,=Q-^+0&aU
4D<5#?[<H2-A_fcS)c>MZ^/J5Q:27/)V1\LLE9aOfQ8>_N#>,G1Od=+fR\G;Z4/9
=<5]N^S^;ZZMI4P,DPB6U6J@IBMC/VNbE=+@4CAEb7W<(\T[DU/+ESXTMR\<GXOG
6ESRAK1]@]+4)f,PR9:Ub1O;Qg/T4>[CEQN:E2DDScg=SXS>PWTRB=RJ?dVf,_M3
F8e[HUOP-bdc4d.TF6ODB1Q11VOf5ZF8/>GB/,U@ZQA:S&d7OKZ<,U^3>V@;#U:0
8,EGAPDfOKQRDYe_EQeMVDG#GYcZ,B;<aLB=.KVFN_6eS&8Sa]fL5++<XZ?HWf9b
Ac3\F29@SSce8W:V1\YcPGe\4\-=-GI56AP5aS=<.[QG=B]5?@_Kg0F,0S9@e>U3
E1^FLSIC65YJ,\5]MYdGRI[X2TaPV2[,&(N]O<ZEUUJE9F;&39U2UD.>08MO^KRZ
\2V]_\F2;8_e<[_[0LSPbNPfAU;0dXc#HBGJW(@?CJ-3<7/E3YGY0L_4JL:bQS.M
K@Va^SL863a?60eFD/Y#,-O]Y,Ad&X.Y+\@b7UO5Qg=FH=e)5W7ACN9b](4N<RIe
L4;W3E\>CISIDBGIT-C&eG:0@]1_QB</@K[WZB4fJ+E?@.GC8+f7>1X]AXOg.^+@
J>ac]Jb2/DO33-7?PG6P[Ff8c#&1;+;J8&+#0UHR\0K)X]gQXe8,X]9K^W]OQEIg
;0K\P[:QNT/_WaN(^>U9,4]REXT.L.PO[#=^/(b.KOKW4LE0LOaK;Va?_X85H&;?
R1FcABV80FY>(Wa89C@A9X])0Y^=2,-dP(&\7RY&Z0&Wa]^A42d9W^Z&DY-8f,7c
gS<933-g>f&<eBWNONd=fI,Jcc\AV1?<,H-\ST&;T2F._>^b3^d^>,_IJ\75L1S<
A?^=@4gY@P9Y(B(^N3-7&[BcGI7Za<3@-.PJg412&XDZf-KR1?Gf\eOf\eDWSWK0
C[42MONM&T>aOeB,_K>_E,,@:;XE,OQA@ad9;);#9AdS66&Kg_<)#[VK9SDD3LP8
AZ0#>g&?U[L3EH]A#O@(@Jf\2aZ#/6G&e88gRb0]=,JO131cX\?O<]=Q1HfPOLTX
?^57+W&]WK?<J3B\QEPODR5S,+-,#ffa28=V?M+:+@dY?=gQS-N>/+)6]:B_I\&c
KPCZW3>>DPB7?C,JA-MS90FU<>QCVRbOZWaT4)]D_K\8G@b[5366AJ(+;7@aVH4G
g5.L/Q8\(aXV:6cTD0bQ/3J^fC3H_<HI1P-2@<H:[,RC&.MIMH]T=[-_2;9E74OF
#QONCgAUPFI<VN[XOAP7=)edDW?70+Q=[;WYg5:_@Y&O^@R49ABREIf7V8K-+9WI
UZQ/LZU;e.a<62P]N5(Ke,b8,IBT6--FP7J-WIPHJ^)&T>[V-Z05P^6bAIT#([6N
ZESTf2((IR(V+O_3LDVK[8@HQGf=4=4PG.1;^g@bIge>cJ9#FX;XX:TSKKP#^VU\
@DT7P?)AFUZg\[(<YeQ]OFE\F;ZM(3&L(eKMM9Z\.[HBVW\=H?<a(WU#A^.HC4RI
;dDaS->EWM//NY_P)HFS>K6VHb0c\>N8WZ==G?>8)BBcfC5H/X0/Y=T=+6)c3-4;
Ec.a\T_\<RF/?QRgU/d-@f1,12;N1XJQ_32]@+.f?.0-I5O2L+@.WgM/5M#^g/)>
J5J[-A+[.3#NFP5:<AQ[Mc+.R7,?#W[Q.7dTV7AJ,cZgE-Rc7SJPRW:X\1QgK\DH
#\db22)e@[EJ.S0]WVT/7e9R@@4-VeY;ON99a?TX),RZ43d,LF4JGg)A6c1VMgP3
9,XZLFT.H4c;FY(3J_I?b_5Y.;MLMI.N4;L6VcZKE<^ZO\QNde)Z90^Q&FI,FQP#
V/0AH+W4SFK^?E?,<60eZ]]79aN:@GFX>c^RH)1RHgBQ_^-C_=fSZA:VDJ/MPG8O
?Kf.3:7gMQ.@6\JJJYKR[(_WPRGH5J\P[BZG<A=N6c)\DZ0:e,)\QEa;FeIOI(M<
U\GZgP_(L&f/9MO,0<&A=6TW8:65A46[&(_T<f>a4dDK-@B8,N&-O1G5L\K2X0>S
0AG+?J9f?dJ)bA70G4-dZHSNM4Y5:W7Yf#bX+1?A2a+05EO4LVU4[G:cHgIN)<E[
B;#D-F@:3AT_=/;^DOP26bb#A2Y63YWT4g8AfPXZ-BC#F]Y7A>XJN(#6Zb[74B/(
Jf_L_]>^eSaM.RKIXOSf6T]cd)ObL#@OZ3G]Oc=Ke@Z_+&,)U;GH/f@#-[@[aKE>
J7AR2.R3KG7g,+55#Z\MW_/GUaI<E.XC,3=9<,0E>_41:&UZ)28ZcFCH&g2RI:]:
<+d28^4\;/=/@^L2^4]\c+fFc1Ma>[RaMWWCd3Z_d4?S=<BS#:&T;<2g-1@/5_LX
EUcUS@XQEZJ>,VHcD-V7B.:\B?JQ1\@/8QBY<>]:_]cc\?Wb]@cd[B\CNU#YfAW)
1G(+829CHB_Ag#+ESPNCQB+@7P/>&cG:U0J>JYDGfZ348_W#S5cb>\L)c99B^.;0
[0;:\HT(:>gXf7VF;HS@\#ZJGY<2=gDd4-a(+<=P+@S&F(/O,<56;)cbMbI=EgKP
VD=V2UO=FY;&K;^7D/9R5C^IYK)OfYONc#&^H]0/gCcH:LP]\+34_?G&2CF(C(Q3
MFOIG.G]#1f<+Gcc)&@^J(Pa^M.[N7@G0F+F467I1M97:SL#OYJU0_-aC7&aG1=.
)E(/?X1SCQ0>;/TD/UX?0#Z(+8P0[@9XK+5O[H3Mae_+gdFc[DD:_Q2:8FLB]FM7
S>#+#GGba1VHAO]Wg7;Xd7)2cH17&/4L5<7UKT,c4d@VV](^EVD,^)]0/2?4D&/Q
[.53,)>/T5AEXT\K7,L)>[YEG-+gN9:KWGQXLY7#BNAOXc12-&Nc)/V/5OTQAEA+
?Sa5:^N4DE#F8I@_YL?gSf4GK@01O#XVg])E@_OK&fE^M)_fgS??@F9<EN2edX)a
<fO;9^)dIdFMbGPgfX/<Q#7,]=[\^CO?8\=11M+96M11;6^</=(]--e?^N\J-;H_
7c:SE0^450GRVZ9>+/#@S)NEbTGQ_\c\FERTH^3(;0-O7W2Q:9]=,JGa;7)5d<^H
-IN6fN\HI2MLb)g&C4bB;Q&\eHXR+f+&9TAV5bTQ:1aX8S.:AJ:;:Mg4Ge2UH@\#
.(L#1c\?Fg46G>YOf5,GO&=T+I_1-5#;M.988IP<54U?=W(.a/f]eNeM+6F;H>A5
dUG^cP7gP?2&G#>5Y5Q2OF#,e.3b]S(KHR29:Q,(d+Y5/cAaD(8UF?POXaM/fZSO
YO)UW+:E&#V::YFIJ<IaKD3+gT2D?aG/L-cH0ZBQ2?S\X2]AN5HR_^6g,UHWIVdE
C4KLge\/g/4LL<VSb38T89[0D)SP78H@_fX4dS8_XFW)N[+#VTe4=WYcI_9c_N-=
/&]E+cB(YKCWQLLU&.Y&e/R1+A+J2gB1X:Le9VB@E]04J];gQNSU.I9:-CAM]EYB
,@=-/c3cHF\I/C^K0Me-P>LC.T(5VXV?(>2W\KcE_/EAVPD1WO?,GYa_>,bV8b@M
\;<.]OL7d1LeS\1DF/);1TXc.)V]SQ/91g&<2XQ\E:LG6/[<]#g_U7aO4b35^O=0
dLe=4[N&[3AKTA:AeFA)V#EZE>JKVfCPS.8MD6\BU+S4;I6KI:^Q#=P5ZaR[BVg]
RJKJWWDP^_:V4W(8\Sf)>[3e^N-HUH9,V\UA[;TF-PBO1aX-HXge&[]MJ[_5,gJT
8=>Z<a9.Q)IQY@B:BN<a]E>D&Ec2=8)FF&NFB5_9]=/^>9UITEe]XHR3K#cHOGO=
-&ce;2fX2cSO-XW_L5,&;D2^-.T_D3+;e=gY?(_8@8O>\B;NgZUIBFcLbO;W.1PU
aX]A^@O7.GEAGQ3eT?,\7?AcO<6[./+U6HHcWEVDIDWD[(QNMFVX4X,K]E^M-bM2
OMG.;Fb+U#]?-6TAa]M_B_(0VUZ\X[07>;<:_>F/1F=/-7f8/U(,3gF4U/:]27/c
>f8N6;>&C:A[:bK)Yb?D>W/Z3aWe),@U.>I8<aU\cR8_-DNBHFX\->RS@:+VB.KG
H=1\MEMSgG(E:f18V#d6,@JS]^YV+Y?/U:W.K./LG(/1@RT=:5K3]X+L21W.6#42
N@#6K6ga6e&OC.J<R=ZCO&cb:RC4/fON,_R>_@.11Kf55\KdKIEBV0f;Ub;e[^#0
<f<]2K#GZEc?P7DG-D1ISFY]60#.)H5PRS53,O/N_/A3M\>E#4.@BQc4BW;??:Lb
C4MK98Y<b=,-4^4/UOaC/&X=,_ZfdgGf9CECe;H&L[7<[T^Y;8A52D_5M_FQ\B4:
5TR(B=M5(G>JV[JW-HY/IDYG.-(FL(F0BX\@WeMUY&]X(87_7==G.;LKb:V:.bPF
aa3O.EMTOMcB\JM228eJIga+Z7T@AM5^ZY>6V_f;G#HYUTKc^F(=UIX.N[Q[698U
_OC5bB5^D8-1_5J,<6Jb&\f;Q5Ab5J[9-M#cJ3d(7B)OPZbb=EG4K8;@8OD;0,F9
6\9E#)3P8SX@:9I9b[&A8(N.=F5D8VA2\1XVf5>UH:S&/4Q7OA)O+R,95-EDSgP^
@]M1S:?\6,GESKHcQZf89B?3K62@?:(V/ZfBQ9S,ND,F73=#/F2LfP7_94O-:E;d
-5H/gQXO1_,_:c=+,Y.#R[Z]1LO+^?M;2#AG;UfF?+P@D1ZaJVGYAM1]S+E77a+>
(.I=;gXNc4BJgE;F/SMG[1S>AdRQ4Cd^[W^B6UO04KICXKI&-\A,.0DWcS.?21eD
).g),?-.F:31Z+&YJ<Qe9TIbL7?GM-87,(;7/eL1B,J>NAcY75#=gUTZ7A-FW2Ab
[IEJa6@N35b.CHA8E^W\KPJ7W#7ZYF&7B.UOd?b6?[NUCKS@-2):3a.+LXE[THVa
;afWC#>\US)94F-<V/C5>&G9d708WaQ-(V;4M=@CaeSWW1AV.L[Zf-e^bO.9.DUP
7-<ga)?E\caHIUN2.R]cTM=]=,T_<_Jg4+NX8GA:e_L@1,bO\9#&-W?Z>>/FaNH>
5TI?U_LN0AC.26?^@[Zc]3#_Y(6Y)OYS;3&M:5?_V#5CbTO,7R+IHfe&gBP1=#Ne
B]a,#I&V[U91Z):1?eeZ)K-XI#.Y6TC&N]8GL(UQdHAM7.-<I;V\J8D5CK#FL8>N
YRH=2L4OM4:g?:TBFJG)@+1P>P;>gTFHJ/G>b5#)?#]3;PSQ/a+2AA?(Q5\.O/=[
Z31S(0U,f@22&-TAW46f#FR;51Y&5a\N8cPYL\\e]M];dJX6Y7&Hag8&@,O=OF0A
f,-Re(ONE0=Db[R:)93UTDOYFEYUG:1W(1@@Da5f86KDeW[M=K#7F;Y<aALBN1:/
Y#fM76DQ5b;A=G5Lg,9;B?@\/@18GB8eW1)2R/e0[VK<e(8E-:.HNcMA=YOT4fH9
0+gJ[1UG<04\3ZPZ-?X^0_?2NaA1_YA(-N13&LX,2(C7B#W4Y0(D6;)55R>.EN3B
HA.6KAWbOdf?KK<4dFSX4e:8M.I#PICW3VaVPAI&E0+98.O<C]3VSf;[&BdgIR2?
2bI]UbYQ63UG=;,^#^AJY>PIC5XSKZg4Z)?6KFE_@\H6/B)6S-L]U#6T=7Y_bcIP
&_N>Z)^?)/SYNAD(e+AI]L,QLO5;#CU0&:d?&L3&S--0McQC>WfSDC#WW_6T;0;:
;>6VN&)OJ<8&/1[JED8cH>66A^U&W6LO(4^C.+-N;;^^d42K^3)G)E;3fD:d16N&
H,S8\JRObPaD0cX-FF94KfA?5+]\18I?IaHHggPKF9/R]V_J=#3c8VN+JbM?:?<M
BNA/eW=cg,CggE<b6eDF:=Sb#]H45IO:>J13D&J1QeeaB+?eDBB1WHZBQZ4KA@]B
V,TX-#FSTC&NB>.<4;C+RS@B&XPNO[@QQU+(ZL\[G6+7HIK69]b=?Pc>3R7A<b<S
,gJg&gT,KU+PD&B5&b&:#B=9)U/Y>9]N+e?EYWX769e9#FPF)S]fZZ7,1W2g?F4[
d^:N8&H33K.[KJ#d>1N(gdb]3Z[6a#@SW^-JT6EB)8H04ZSRbXe]deReV6YJ0T#H
AS->#(G/b5d=:e9#E1XW]1#(]b,\HVGc]gM80>X.>M4-1^dT1->:(R8Y]N1(;>@g
^f0&4Z,0O-KJ8XF:&(R,5e1I^fT+:S=T]5AB.CHI[R+a&3?#M?Vge91(0:0V@MaZ
CaJB-;/_6,;,D:.<eX-YU9JF20&W,(3IF/PB&SaT-5<WC91GfaWQQ3e#=:=TPdUK
PQYB5&(bRNX+#V_N_^_KUR^6A1^fMO26C@,Z_FUW6\(]Wa^S1)f02-N9)NA+3<_>
=2eM&C_OXEWHK48OT/XXg&bXY,RBc-4LT)L;A\P/6_AV[9W-J@YBEL.g^B/#WEWJ
I(CSQS-;_)&LYNVALM=Y3(f)E&O_3KYV:bLUV_:C(:+MWH3cSWX9bJCfII#0,/VM
CXg6M=Q^H4\764W997gSWSH(U;.[UQ3>\R6[D?L8XB/7]590V-^ea8N7RCUW#U?g
Q82g^C6+W1f5d;+;FZeY8g^VV##FLfQUQVS(7>aOD7S2PJ5:_O=.]?#&FZfdL@E1
(=T]cVIH:J344GB#>MO&.>6.L^6W^1S5bSA5)P>E&_HSS7)RE1((8K61.TB&+-c;
WG5@H9Q.FF]Y,>B(L?9?^FVg&c+GAgg=RZe;<5+U.Ig\,2V(9(&TSINT(YaeJd:=
&F_V9#C(VW9EVP774LE^MQ#SB-+FS]V_f[^C<>3JIO;(8=CQR&7?=?+_7<Ce18Qg
H9bG(D<UaU>-YdIQ>aJRdXN6+PN01AT7Nd4?c3ZYO:/KYFSAPa)@)Ecg/B\CP:@Z
L5DCJZc7SZVW.M[YLa?D7)6DHJ5.>7-=)S.6c/;U[Cf:F+?:8FMKEb6_eQX1@6)Y
?,BJ7&(9FS[>6C6ZA?-F6F6@&:]4-2?OJ+69^g5AI_?TF@,a^<T+;cRO4.dO5;A9
Id+J.50XNPD1:N_.a=)RV_\GQUbA>];&@.IIBHK]08@VcDTY#/B)a8[0K:9YC-7Z
RdG6E#:@EVPZaPc9T]TCJe/JX0@C/DC_(K=8eAZZBe>3>#,F1EMYA//>2ZS,XD#7
1+9c;^ZKY.RE2-UC?F_NI?Zg.;]J_8\^B_##(/?F]O7N2_IHO9U,O+PG&_4T::fH
&PPX02T1b+^=,bA,cMde)9cD[]RT)V);PV1IL06Zd:N3:29#79.e52PSgJ;40a&<
M[YYL9H7[;)EH9BB<fC;>ITUTP:gV?(,7gO86VM0,Cee#NgOP\gW7ENC]SbN2HNQ
;3aK<2;2#^U?@Fa,f&.7JUZ@:IS71fUQ_QN>QX):PVO,BBX^FRgg3,D[.NX-\2U9
W2@+VfT\06b(J\&#/D\OI]:S\6V0N=?(I-UFff=?]N91Q278Td4+;.XO]H,2aC]A
7+;?2NPBO)2]1@cBT;+9gT_P@5)H7Y0)0AJcc_eJU>&?KJJ[9F].GBW@+/PBT:T_
IGb#4X:dHUIcaUf?D3eL2<80g+f];Z9,^ZF#WZNDMa+;1N8A59W07VF:AC2Y@,L,
P^?aL;4MBA4eB_&V?+4A\I81E#&91UX\,IUCY^C>=a[1D8-Y)+b-:NPeGWQ4]#4I
g2;A?BZb@EE5N]DF?N6@_1+4X3FgY;-_:74J6;0#/\bTc[>YARX.5>,3b#KR]gQI
6g:Z3;[Ae8I7:bS]7.E,[@Hc-bCgaQSfMcP3FH9&OEI&TNOP.QJTf-;>UL0I3DQ3
:OQAG_(@+bI2IFJ>dTO-bG:6a^AS;+ZK9S@N@=#ZYWHS[_&>\^\>P&P^?fcYbgYR
PH>VMb+1WBK7AeK_6F9/2#LIT-DL]NfX)-7SPF2.>IVLP\K,;-30>3]>L;g:39_a
@G@&^8V20Ha-gVGNKdWf9LOD.?)-4@GC4QQ@L_3a(PCTa_,60Va&:=Q2(Q2K.5gZ
ZB[gU2HKQS?#_20M[S5MFTKdJaSE.ec\X<a+bZQ=UQ@A=@/?.=4-Y^:&f,ZCg2L;
b24V4(>f7#I[3(T=\bE10O?E9ABQcNZ]7L.aRTFa^_20,,:FKEegD4O=cFCXa1S.
)U]:AIG^JN,#0/0HUG<QTV#69<:2;G/&Z@Lf5T^;J105E<XO.6HFd0&V-b0?&Rg=
>1F#79I9H8(\edN.V^@A65&6fRHAXN2AM>dH]7^C)0)WW4(F\_KP6U:PK_(IDIM^
Eb;8S0=2RAG6Bgc0^TBR:&b[D]MTe;c)^>3VP8WVI@=g.OZ>/1,M&\&Y>Eb74HK?
&NAS&#eJ=b_Q9_cF1Q\?96B8L,,J9:QYBc?+1Ua#TVCH6U)GAW.V(^A8P2<8bf1_
>=@eV8K0N(O1A>&C/3XNDAAJ?[b8:(AT;I9D3MFBf-6Tg+aU\JV&6/e?\+R2VEeH
#F@NAEI5P\N1+5>H,ZJ\Q868I7M1\.S1+O<_:=f\>]M(L<>^\GEXA#@2C+2b1\1V
c;P2=6(J;5]MG+WKDFNM;7WW=.b3NGAf^_F-cSDHFTVb9<+=&9-^CM2_[cGQCe&7
OE5\)cGKd(g:I.<eR(5-_X]d)eYL1\-dOSI-gfJ=8UFO7gaL[R^P3:2Y?G)\Af6g
e+OI7_d-;f>)e1f^dXGT7+ABcH7)eS<g.<4G+f48?KASd??Zd6Va1F-.bBd\(8IZ
LB2,G^6[SgQBK8V[B1FDE7NR,>O#0);3=(KfD.E8R@_K3^@[1O2G^A3QFR7G+.\2
&c]-a/c9bcD6G4<05XG@?A(C<G-GeQH[]4//E).<E,]@IILg49gAed<cB)6#fGg4
TIF@M9<IYKTb9)2ZgE,]D;14eZ;@\,]&U84>36H]T;#KR,I01OK]-0U^)R=/R<^R
\@K3-/4I;LG45QdSUFZO)?49<(XN=c/a-F6LO&RW4g63<@d4HEK.&LB-Ud8[ZDeI
NWc^Me\J@9M641@Nd^Wf-7#8JT6VM,Tc7VQ]XV9T-#B69d:J_QAS,Jcc&KX;2M4e
DZ.c:3#RJY<<R19YSBZ+:Ga9:e4N.+aS)4RcLW8Wd5g3]V/F@=]?O6CKPBB/#fY1
B1dON^2_:K/-]HM,fN+PE)F=Z,\WJZ?L//R6V27(bOZ\T_(CM>c9=Y+Ga?MAP&:E
eTP>Xe8<cgJ]RD]Ac1P6;K9J9aUaR?7OPO;a5acI:b0PXgJCHR(>Ic24CCd2#4/&
JNc(6FBL(d+/(3R93J;+)ER]U]\=Be8<QFUOfC.F=,I6)O(8@9#EI-U/I,aeDNH6
S&@3MTHe_Y1_AcASUfLL^D0;8@)MB9d8dXU?1K38=9Y)6XHab>=W\&e\8<Pfd,@9
^@a,Pf\N&67?;Ba@d7Z?Q.?#IH2DL/?5Qf#&Y^.IM_.#/_4F7O&O<Q,:AO;)@C2U
.bQSX\U?5E5f#)IDN/)WaG#F@/]L^CT(N6+Y#?9<8Z?:)a4BF<0,6X#W1Ld=H,@C
Z/DLP;XUV&LRX5W.ZgT0^F^&,M)4<^8#>ScE:YX,eJb@Z](1\91af-&?3?+A7,=g
4F0^9L,]8b<[YZJe8HZFV@PWT@aYL^P?aIPaCD\6b=DcLFVWVE^=&#&8(aR0Y-AG
(#c0IO=V4E#R?W7:QG1I]E_JPc(gVIfHJeJ:af6Jd+4,)19S3GG7:[U9A_3B;gX;
(B&V_N_Xb[X)c69EX_S&BV6E#M_?D5PXW8F</AcH:=6Db1D-W8cZ:C)WUK6.TdVP
V<)F8J3(BYF&^#=B,+^:\/@;#aG>H+F)WT3a]3F&=MbD_=?VZ0cC+D^1DQTb&;I9
9a<.<FYIV+O@5f0B5LS11A=Aab=-6fRSEd]8WLNe.O1S>]IOC19BfS+ZN8=dW;:+
OY?(3ZL.QB,2\I&:^+^KC5\<RJg8_N]gO)QKJVLTUfR0W>31QH[0-<(/M[B)4g#H
ZFGgDg5O7-TFTd5;H2Fg;I(Z?<#f&&NISc).6/R\[<PAY#^U;d(CK8Y8?\.VA@LQ
[K[b6d>K.6KCFO[N0TGW+ad4cbP[Kc[L2U4b/A3X),>I4,.Aa:X^59J5WBM5cJQd
?4GZ&CLMN]P]6G<6OM(]FYFF\4-1&.>EK7]07]Y@N]dTfK5.ZL+J,V(9edR=W1a3
(FCUKH;4W6LPHL?_1ZW^^Fd4^a.=[D;1?O:CTd<+R7X80,;AZ)=UJDe&dL96P3f2
++\#S,fb+/F0D(+QF:=<IMV(>-G.d<[.Yg\K@>F/TA](Q;0Bf<Z#T/4R[bQW1A59
CIUC1PZd77FQ+EVW8d6P[SJaaDH(O]<DJHV(<gTMBBSMbX<d1/:4/:OJ#82.BR6A
R2JGJKc0RE?)8>#ERNFKFEV&>ODTa(/;PadV:AdX@eV[e3K8][E.WARZDP@R4Fb8
JM;U)SY89.]1&VDDO1,a>;Z0QXJ#Z4MZGP&J\R^#d,c_OI8^HK^V+[Rc0XCcE?,X
EF9JP;Z84;aRV18^J)A]KOYVaP[MB?KVS0Q]fA^c6)=&W+(86d@c2V8/geGg5.I0
6)1(+ENTFY1TB[SLL?ELJOa_<Bfb6U_3IgIR]eHX&4TQD\8&,WFKANSLOaO/b\W:
7@3?JGXa;TX<R9RIM8c?3_f+2<6&[[bMVaU<#_3+>/+BS=^eZe,@g6J6#MP<)JRT
LS8cf6Y>E4(@K<,G#7/XC&S/0Sb=L1Sa+TPA>]VI<fC>]<N2K\gEbD-_(NZFg,^B
HBUe+XIZW^23CSZ4N4=M27=fcB6)2a#bV/gg(/T,g&LA>ea[A=KJ=/,+bOTe0cX\
FVe:MP:D&S/e-.IG9IT4YL=>@MIbZcF4K(DJHfbeVf5IWKeVIQ7a3g;H^T31J\,g
,a:LS,37BP[a.EXK#2;K7D)\?26FQA_a&D+cSQI:8=6W,S\XZN+CB/e&JJH,N?IN
,(S>1eFVO^6T&A_2NDYc4]/:EdR\.;P0;6B)gDcd4XF=9V:dU5@7d^ZQdAU.,(AD
\-?Y<.N&QIF^S2F:ed,#TVY-5=?KK#ILD#,TRaa0<&T<;WUNAVHY??&6FeQ1H(7Q
<8ZB/.72f1(F_Ld4PG-0<Q:fb)fedV9]>[8S5;e^(9(d78TA3&0D]f6/,Y81W3]e
GX1VNYB(0d>:Ud?YT.AF=T^,f4#>P5cR[VO1fUPJff30A>=f3<Q+JZb9N@O^<^g[
(1ffU^Q3T6#7HS<?&9I@BC:W:Z-,7V/=PBa=[?O]BRXaL4GR)UM=bP;bVOeDFO9^
CZ5J>_aV_\7D/:O2V&MAWA=<<J<6I&#VE06>We>A&E\ILe)0V_Sf62Xg.+-]/WAB
:LWAU:CZJT0B(&cd8Z_b-RZ8Hc_0Nb#UgGX_bQ@FDaY,bS897R;[E:G]A[:I2#[H
S;SDe(-Ec9I,.:[1-DJ9_+I[Rg;FNMF1P5&F]IX]/F4[O<0_[7bP;eJGC^9Wc552
1P,I3.EI5WI.RaH[0P4O)6.BgYda:f_F&E.+U;/ecbeAV6SCS/4L1RFb;J(Z1NYE
\_)HgLK+f-_]Y0D/d&Yg2(RLWB>.S:8OT=b./JfA,L>J12&<>,P2:gZCcUfN=WbS
d6YLd+_^f1IHX64#B#dJEY_9S<SB?[#Ga@LIF7QH.K;V&<Gb&GJMe?ZXYMFXacPD
Hd[YGcdAW@+><+NBT(gM3@d@K,F0]=b=Leg+U>95FEg5_>X4f85c09^MB3[<b^O1
(T0IP66cF@O^-RfZZNTX1KaU>/fCcf0/R6D9(NJbcH10bF>dLQH@Z6>F=5L.Y5JO
4@AB,^MBOfHX4;\f;N0D8)\+66V9_Z7]I43(2/>F].=bJDg^A_>]X3XJ?>R>-23C
E2]CXR>/R<OGQY4MB6eI8GFc8@BZKSY7Z@<.,V<.f(&SW34H2ESe#[Q][L#6LJAA
FVN3]33W:,(Q:6KG^&g<P3LDc_ECg;WLW+3LWY+:841\+,;\)]K:TVN-X#;QC>fV
-&;?/_H38-Ge\dc3@/dNc4=@)PKBLFHW)dg1;S:bMOR>P3?Ze(>If>]GP5+[VSVf
I8af#+N@)\a&)(V7e38(]GbdUR59@?cJ0MGYX2I]+Q#.6;ANV;eG[PSJBa_S207D
6-9(Y,<1g(,c^Ycb<Q(H?]GeaR<3=>B?QU6NUa96VFX\dMeMa^6J<J.E.T(C3\S/
_R-S[Ba]CgU;VM4XU)A#2Q_A2N@3+8Se+LA)R&)<^&0-R_CeS-[TRS1PR:Pb=P?J
AgHR-<S2^3.L[VRNTI^\&]aOTNZ;0f7:43I543e>W\;-VWea3(S=\G3:HNGcW:]K
5:?2e:@K)RL]H:_&EQM(<4edXNUa>C6DgJVXIC0^MSK]e=Hf0B[&)\7=(>cg)4@/
eNcXR:V.#PWNSaHP+L1M;6&46Y^.9XOF<75aD4B8-9<P680>PI(H:4=PMg@Rg5T=
4([bOgHc_[2TBMe2UHTeL?3V:I1#7TVOU1-_=0<N\e;FEKfI62E.>fK(T>7RW-A5
O/-L]=DI8[CbC.A&SegAR0R>a#?[HOP)]R8<&=;TS1L?.C2\(0M2_IZ)/V9>CX<E
8bA[SdZd9C3LWOCG8]f961f]IC,K&0aeQbbL6W+;dFBAF_QOF2\S?&R9:Ea/U./f
0>@fWBO8/?YQC2OSPc;@=]<8MPJ(>4L,WYK&C<>P:0-eNMA5VB1T06.0C9?C=Df7
GYV?^2A);S;31PI25]K+CU:D\?@b?,YGV2;W+8VXc88afB4)/RD>Od<c)&R8/914
aA9=\KDLRR9PC4TRVZ#4G\:d[F^?MQJJD>cN>9;3/2NW9Td9Y(R9\5MRAFb(1U+/
4TL3CT\cb&=7KT+QD]TJGcT20.D?>=C16I?)G5_)QBI=U^M9eIKJ[@^@YE?6^KZK
C;@D^/X9F1NH,6947P#2LP=G,=<&G2I(EB+Yf:#:LP_8EKMG)RNIf&;VWNf;[8_N
ZMfUeAfF\ZH+AWR=1#8eQ)H5F#3A,QR&a_/PC>ZN=4XU)=6G22N;2K6BHGJ0b9./
&G4@51PdG-H5Ga]a0_(f+VA>dBN@f3T(\^_<,EB-D3_D_E[0(9]K3\73DC&TY7UX
[2deAIf/P@1#L8S@H8Ag[L:U;FMLAdT&UE(]b46Be.3,LccN)12eVU\/<XB:P-+7
HdU24?-a90B-W.;2FC>gWW]Da@TG->e4YeX\=U\VY58?6@<N0;9X;f.R]LI0?H._
41#W=MTC_N-H0]F=_DG4_Q>5C<LQ4JLL9@:g^OJ\eFUL5P+;+=.CT0eT;&8&6J)U
+g8PB8.@]]g>\aZ?7[07KGB+,E)JM;#a\aN++[U5^-E,]dS-H,Mg(Hc\7I#A,>6/
70H00&6cXC#.LdH/J5,C=/54g:.KXK]57S46.+XBbK,=V+M1;.#]9<c271A(61Jf
P?J944,JN=//=b;>5GfObHd0<-TPDc?7M;6&ALdIL@d0[a=.P\>6B_BV5X-&CNaL
_&F/gX1N>/T=QEL\aM/XdG[K=(?-4P(=LSXfKgJZPB1fQ>5E&(6JT20MeY#L[-]3
S5c3-:.N3A4(/^<2fB-@A8O=D308U68UD3ZSGFR),_LKYJZ9d/GPa@Db]S,_(3Qe
PTFX6C[)F2#,)D,3WfZO+?=.(<//2_U(:,G15(\PP\;dKESYT6-Y;+CQ3&A/GeI[
FB4]?JC>:^SX6I(X<,^)H<.W&7R<YHPgaade_+EP/^TE/J=Q):OTWJ8E4SF)L[Z0
>Q#/U2^:RJ4X3Rd/2JR5a4JcJ1MQ_Q]DXLML<F/d>\Jg.A)6LPa&bJSeO6fUK2O]
.KR]-,PMX3@;4+PX8Y/4fI?Oe:fM868b1,9&82NbR&9B5KI<cZJN[-M4Tbe&XaQf
W#YQPX=@>[RB3XWN8ZTIL5A<]J1.+f7bEI)P-/YDJ4T9Y.YW>gC-aNLKVOaCg-:6
A+3AZ((^d7.53[Y_^I2U^2Qf<G?a8=<(g/@R#dU8.R0+I8Yg;WUZU-75&8Ie=1c.
DO)95Mc=cF>FcFNZ(AGNbK2<NT7D?M40;0GJN5/^8c6CgFEcY<6G(VX&)KFT\OG>
?>g#1g(1OTN5F6T=,Q#/Dd/@H3EQbJR#KZ]K/Kc0Y[)UA15]+?Ac-&/2;0@3MC/5
^cbPWdOQ;LOYXeb-0_?,C1U&Z-+9Rd^1-Q(OA(GFYeYU])Bc]8c7PA18YbR@X3[)
2H=ObSIAdf=O3EX5&g_Z,/dLT<0_:8\[ICR3(+[Q7C<([[2+^YRDXgV#2\BOJ;38
((=S89R.[bN(+=b&_=F-AJA1][1#-,7XM0)43_YUcQLZd1a/ZgPe:I/2]-(<-NKb
aP#:8SLCU.gB9SD^7?9a\3WaD2Z5)bNf3b4GgMG#X<B#9L0?&=Wb;PSc_9B40T[-
[7M-G)[<[M(M5?TXS[(cR<BL<aY5-c9&G7RRZI(:Lee)((?O#E2fF,)Z;eRB2;+)
HMV5]26P)P+Y?_c1d-[bPP_ff+R;,S3R8FC?WFO:KZBE[\da]&[QX.gc>(@ZW>dM
A84KGW00.A/N=87IM\5/If505INL#g>DcAWQ^faQ_4=c9O,WA/M@.gD2aS02QE3N
a1PP1R55\I_X^6QMG7H90,?U6+F4N7b)fL)/aPZ1DANUFbQbM=^M\4]_\[#C1fF?
L&\JB0bA1A+,<0+Q6/AOadY#<0X:_G\Qd?0a1S_5F-g7)2;O_PK(1QdIKCB+gFHA
5c;6T1U^Vd6E=Q?9]OU(_+cOe8Cc8C7-HMFaU06^SS;NY&bIa6>CW5Ud1(<b/_-.
>Q3]4,J#ZK,Y8SWMb2FaU9;@287R1=CLP67NV+TbR:7X]4G.67/]OKUb>\)NEBA_
bcK;UH3@N6>bQ\6aaX[X0VaZ_JC@?<,&<O9=T55HL/^W9KOCbX7H>4CU;2a:Z.E\
dZHa,#;f/C0dNSQ;75<>K7OUV+4G:KP06bde),\==^?NG4a2UdW7LK)PR^5.KH=S
TaY/8HJ7^?J]BHCCa6,:RHRRV8LV1(BC)[UH>:4=:LUJ(AbG-IQ9<EHT;3739=,1
g,H/#4g7HS5bRQ88gIRG,[Z+>-N>JJX.IILXW>bee7]4=<JHc+LI:ESDJOeXbF<G
>V84PX^IZd&[/B/M6KE71IefL]cR/[:RGQIH)]/39=RZ-0SG371a)=9JG,DeY&-F
_+(f;A.UV^T__Q#<GbW&]:\V;Y/N9J3CG[CG?4SYLIaD-<(8V(bT?7:5&/^Z9bXR
<FN/6ED0P2;J8Z2,WaBU&ARCPCOcN)2=UA2QH3]#dPJN9];>dES;?,)ea\Q,;O[L
/bS2Yd(Kc?ITJ2\G6VK+EKP#Ra<C^PVJeJN-,IIAL;JHb^0&V>-0d&WRTOUW__Ra
VH)&,S0GP><J#aSE5G?3&+cPMg:L.(NDf;R=7)dSM863WV<@D\VEYN)Y=O)LPJ4^
9f>//)AP#IT3&HN9=+.Y?=aAIH>(-a423dY5Zd:Jg3S5Y/gTdH&=9BKbZ[.3P,UW
^Eg:G2G#4IK?MMP#@S;fUR,:9T)S>fXG&QTTU7/3X>/I@FB,<4P@eZH5c_e>E_T7
[Zg7?NZ^.V-<OSb<cP7;1Ga#KbRZcY#:2F-<f#f)5GR7+TfcJ?/]T8H13E>]7]N4
-QFX=d_6&A3QP;E(aBH>V<N8;QC^D48/DDCBP1FLEJ6,:E]HLd7OKbKeNXRF^0HW
B3AFT9PVLgbN7D+6)aNSJ_L/C\TTJC<]b0/M?:O5,9]f=E^3DAWe=B^+E;bIcZA=
2RH,1QcG/I9T>\&E^a/-3X-28R7V@8bB5gX\^MO<DZ^(\J59?GOOS@=P]CM2N5>#
>-HA6?1IAD08F\3+R3R]N.YbU/NILY=?8e;;J^&0fJ]9BU&UD_<\Y^-RLg<17:aY
>251,<SLI.<)W#9Zf:e;:?0YO[#f>>K?ScFT/;3#3+d1]FXbE4YCSfF6a4@aKC<L
MZPF818(Ce/<A9PU_g@@T,6F&ffG;5VY5d\8[<X\\+Ga]1=_\^KJA[]>g.\<,fMN
MA\RaNC#d=Tg\CE)]E4+P?^AXW277gbRORH4??&^E^d_:7(Y3IEB#BETK\>FF]?g
-I8ETBV80VNBK.7GHOCfZ0EYcEFNa,@Jd4^CYA52_-e#;Y#[6)^H64.=E=CQ#)K:
&Y37g4SDMX5&]\d>VVLQ2]SO9:bD.;^D1C\#>I^<X\gX-@AEV2e6_HYK>T=?Z1C3
29(L<Hf,U(D-ZgAJJH(Q)aR=&)3RSO4FR\4MSXRGDZ.8^K--\<J&B#0Mf>R.@Ha,
SR+TLEa;cQ7ZL?(.P80c6P9TW^LO]Q1X:ffb>7NKPW&Y<,C>/U@D);)dU32bCPGe
3_G7Y=CL86E&\D[7[]d<@Q(+Da\F,ObaMJ[.O,T3\LWON/K:fKA^eL_K4F&La7Yf
V<H6dG7e<bHV0OW-:ID,IeA3RVdKXN#L]f4R)Le;.TC81>ANb,J?aG_HbacK,2GM
>A?;&/TK5@NP;WK&<4I)LMT,KW8:T/AaO[4)R<)J5^DMfED.\Z7MWOV&fTV:0DZ#
(?eG_N?(JS7?GOKG.V<2EKH^ge1)[&3g[ATfU^a2_d2X476RZG;</7HT.)<,YK;2
-)>6R?KcAE\T#?6(PHaNIK;39CbV&,&J^>X0T?.f<b(U]T:VM4(X6b=91W^CL^DB
?_0:>5FW#+_T:U>?gTL+42GB;.Q_/>VNU;AX(@<F>-bc9cQ))VX#;:[O)-8_egAC
B\,SX;,5TI:ESb]3_;Cc_;)[?[\L>DXU_-=RbXR&,ZZ?dYO:XCD[/OE(-bVaMFUL
S\S]ABG<2+75?Q3-d2F<b4b^TE<#DHaGd#+:5FgO4C2ZZ6H0bSQQfH9OcM].2&b,
QGD=E@RNSZ5Zf7;+)<=b5+?9=<N+e88EMPJfH(dccd1;:gH2eH[K5E9>_a-BSZ+S
L:0>E\\7b=a2?b&O#AZ/F7@5cH;S&b0[P<5)ZP0##WWK3DS0FALSY<C/D;7L8,B/
+6H\eLWGRDc:XB:VTD&+W35bUfAaCI?17K-_(^4b?b:<EEb:7YG&3fXfed=3dVGZ
\PUa+FKI=W;,[AbKB@=GB5+-0L1X2S?//geeSaC^;(/G,JQI4-=].4B6RI8AR57^
,gFgU\W9G#N^=KTBC.07a_aDB7(K)N3[bR-L?X78\CMLSe:;g8MBS(R6ZS6O4YMU
E6bMCQ=:eT?PB_3_A=HgO7MMg#U1O;T(d=I&7daT8f9-T3L6D5ZJbR2/4KW[P956
@(#?[L63[^1Ye>7CE@))&>^RZO:-+#GB[HcZ8OS<9HUCH]g7_#D8R17PEd^HZ2;2
DM?E19Xcd82T#D=69a,g;Z&KEdMWQALMJ)?-N90>7C[#_c^]7,X_#WF4N_Ba@b0K
&GTGL7O#TL)\S++dF=A+<>KJF7]/EUa1,Y]Cg=.+[Y?TJ,V_9_VR<X/(S,40BHF9
d&W/?3MU=@@.8_P#QL;JQ8_861@fJS6HDAZ#dDB?E?K1YS1X=A=SDI@gA]F(Xf^a
B;BgO97e&KLQ\O679KTa@[T3J.Q,cR1\^g);\7=&e]H[LLcN\UGZ[WP>GS]^#,PC
[4cVa^a]6&a_8,&(6PK=2EE9;N_M?][K^MM<IgGIW5&I:G1=?bO[Ja#;18U1.XQK
J@ED[X#FQ(SEaY.cD+Ig,[Fd\<cEK3+=f#=^D\9TP.Z\]-\075P7gK<BG62fTeeD
\@3<C+fI/P=MT-EI#(,O_bgGYUdA<N;:JRaJZN5<B0T[UDdZ32>dOJ#3JTQb+E\L
QgH3WLX^^-@gd#T^fRI@W+-URfED&37@KO.2S,]VE##[fX24Tg7\>G1N/K3UaX>=
DD](72T.)[_ED823QL^D]HgcBF</d0.B_P2+#[fM:)?)JFeSg,G33X=6c)U,HBEA
ONT:Ue7YZ=(3&&)3_9gWP0WC#_BdOFXc(Tbc8.H8MBc^=ff&_H#e3:-6VP.5P>d:
V@28g-T011#X9+ZV(#aHZV\)<D]FRggCN/6.g2]SIF<aM#f]e&S:CSR+b==Q-;OJ
(TU-@@a@DEI,5MTg1Q2NL3Zb3?gG[/_(Y7gTdBZSeWc8e<A]3@fP[C[9]a)S;<-2
>00JN,(KHD[;_@(SSF-1Q-M\@R&7DN;[EU;;3KE)7aBD_2U^I(ga;QB+fJDac0#8
TcAAPHK]eD,TI,)Z--C/F-@3#GfY(f<3d_.AFQ2OMO<cN#gLa0S?FdC\WO6Q?=-<
<=.+QT<XE,X6#SM)&>aK)C6-P^NL+&.L5IXY[N22F^CSIUfZ2]4;\XX[c_f_9a2_
7;1<N-cGc)5;(/H1-3EO^/F+D^><F2_,\^LKY#+@=N1MW<B,@5.:EK#K2P,1(Qaf
dI<B1FB.XD^-f3JJ6&L82.94;0M?ME(UF)ZZN>==g4JSRKf-[KKUR6C:B-S0Od\<
8f2eWOR<cPY+b]SRe916Oab>8.8>]>:.>\gJU-ME3CU3L=XEF2_/(F6P2O9JPAV&
R?+AFK#A5.f#c4<0X6L#O5UdB3R<(3-0ZC_L+a<e1Fe>NZ@2=L\D0#OfE5(LS__N
<Y_1ICG_^SYfOWF;E=J=9TG[_U+WYW,?^H[(e;3RL@<=Y+S#U14-,G3ZAC=^bb14
_,@3U0-VVf\5411dNGKGJ8(:V?LV_4LLTL072_@acC9Wff#BS6dd2?ZQ+4&)X:C>
J+@SRJREJdU(>IWN<6M0HK\YQ)A[);4XTefIH2]e[NCe<&(8/)2LABVRbPLeG]_Z
#=ZPUO5;51:E9?N)+:\+e:@aK/_B++0:K?B8Y12B+NP-1W+T_f-7USNS2PSL&_6&
fGM\Tfd\+#\5/:/BJ@Bc6[[T(7GdW^LZ=X_C]4g5\^c&Ee1+/UG.fG4R([H6H#\X
B2c-WdSa@UR=2Y</A,<B9=d0XCYaO=],TEB,IF^LHKYX@(<d:Le5TQ]=Qg8/<.OV
JD\.PES[ga.4SY6<YYQ&]&JI1V[R8]<O-.gg<DNe>gAV=B(WR:J/(U(9]\Y&..2U
=>2f>]\66eUZUK_=K#b@J[XVc)</FG]9R5RNX/_0-22Z+;Tf\]5?G9J0g^<V/[X\
WbC\6(6LSYGd.95K8;W+aH4cC3W)@S@LO)E0BfU<eEQ,S+K5@_OOYAMW?>FT\]g(
C)Q5Yc^<DgU1eS,a;1g5#bTfE-#3B4Fg4VXFVY?+fIOQKXX7:CNJ;NOa)[OIaJ#R
NS=(TWM6D&J[UI+QAd[Y_?<OK5J8H__+Y2<9RdPT6g.KMfJO4\A+0:S^D<M/G(.E
X?@Q(V7L_VUWTV@+f+OV@)ZV7KP,+8XKNb8g_:>:<8IWR^gWL;O&GdC.O.]IU7b^
C&-LdDbQ&VcgL1J1=[);4+,]8(G#D]O72B+Mg@7f89V?@.VX/_T:&;Fg=);4]UBM
7NO>d:X[b?Oe8M\_0=87:1L:7AO\VWCYgD&K1(SC<Y3562O2NX+/^VN7JP4VJ&a8
FbM_UEV(N\302eD9@?TW+R+<5Tg&#FEaUKePBa:RY-Gd<DG7T-5ZF[)N9/DZ4U]c
?Pg<Y#=R@aGI_Y<@;4H_O>4.TW#RVQR.V=6I]UR[UfGEbd=bH57F(H?;UNYTbA0V
Z>f318->ITJ686K#)QOZ?#M\&&.R:G,,#R=1,H#P1I5=dTcK;cY)SFVb3>Da_I,^
_1I74X?a9+GG7BZLGH?_a+H1J.@aa;P\9R]eE_&<eD^A>23WW=bSS<^WQZLH@GYR
Z^eZ^d?UT@HJ)@R]^.N-I(gV#8@PWVOf-X,6F5.&3d\55&2f(C>cB>X#.4VOO=33
bea_XFg:Db?Ea(8D@9\;dY.cL5\G<AKT9CCU>EcbH403T#eIFP&(]MGd/RK@2YRG
UIQTXDeFE]+2^J:4BG/6_D\_;f>GeW;bd/QcQ(K09L&&+9I(7)?Ef&(@X[^PUAJH
bZ<#=d1O]?b#4+33],.++.8]#:=;bXQI)S5\;,c+;)SF>5B+I2KOa#G:2J@K(4ZR
gfSZD#R&CX9EPK@=aG]9A;Y.X/@)KAVTg.53=WJGdg&gC#(GX>5]_G[5_5fgf(=H
Og6=/Z2KTR\DF&2&9:[7g80C6IY\Kd_\0g+]+0dF9[A+6ROA_<AX^_17=gD<e;X3
55I8@CAJc0RKZg+J-a3O.(Oa-d9>cGEQV==(A<\:(La\WJI/ae](-AV[,-Y;A:b0
..:[<MH]9Ka)E2(WBBE\\(6V<a=0fV.IEO:bL]FcASJ?X?I&]&&eYYNG<03,T>+>
T>Pe\/[5cXO#+=d.N<##.2[IGAC6T9d6-^4Ed7B3Q64BU]L[_<@a50Ma:Xa7((N_
^[&f^>(O4D]P72,dOJ(Ng-FcNGE.OUD3>VgN-H]bfgTDE4F[K]b#3+\E43f1\&cN
9^_T<V_eA/8GBXK5#,XT5I]H1>gE48eG)=,9IW9f,.7Z+dB<B+X6:>16-Q+V^7,Y
.Z/>CYZ.CV>OB7BH=.:5EEZ4DQGD2X7E:47L0Td5P+I2CX/&:V)X18\a16TX.WK5
F-R<DcVCAcd=d&,M=STa>,_,)fD7Y&=[?KJT,VPZBO@ZOLD0N75:TH]6=X=N5(TO
@cgC50:WV[^5&TdcLT5IBgR)1,gS0XTCWZ&7eS3#_GH1X9=1d,cgO#Sg9dW#VJR7
R[C3bW_eZU<940A]4SYC(T47IHSQ,YIcLfg9Rd^2a77\(Mg/RgJW)9I1@:e:dZf.
E3JAaW\cI8gPIS>IgcFY;4-PPX0^6CZEQf^8BW?/#J6HTg)@3-^aGWFDTaQ5S<+.
eE.WOeP\=#9R#46Wa&APO\^6M25.LQ<I2/=;FETD5-TRU5J-OR:Y]Ba]L]NTU-d6
dV.W/gagb5E&2K:.]A^3&J]3gaCU4@C&6E?K.F\P1\NGc^(c@ZB[=+J3\RT.E_>@
>=c3&OQD?Mg1&JMHQO&IA+>0_6([)gdWaQ??37eIe?#081C;fdWOPWZ8aLSgU?&E
B(Yg+ERgR+Qf;R:d;B0UTX3EP94aZTP]a^+,/[4Ke^fe3?5>@Y@>/H2S3a1-&:fV
CLY(UIEdA@a>XXFAXNQRM4]g:666\Z)0AYDY;ca^L,P&V4K<BYV@_#>5QXf8a,.N
1AbVT>G@R>Xc0WbR=3TH,9DRYD\J,.GM_:-7U6>0a8H)GR(OKPdIXB98bcJUO1Ua
E0G,FE_WYZaO?TI,PU?d\dX0VV1L1L>=S39</?fZ2+\\=-M^([b71\B9f?3B;49_
\S:gUN5@VNYJ40,_e1@LCX)Ea.,>Wb)J,HX7[=/HU&YeRZAIDKBd+802LFN1P]YQ
O]]&)G;316PQA/FLgODaS;^OJB6U_M\P2;/G1>[afWY5UWA>8aM]d8MSgH,U)Ee9
P+#FT^3:Kc@\a)?/_-f]]d[FYfB[fXVg^&7IBWZWNDR7XN_Bc@GI<b&c4.[Q@?8U
]HJ0=VPD:FU\3;4^81+@6BeIAe.)&^YMF;5,A+,L3[(DD^(>HD:[(Tf6,8cA#V]Q
J)XaZ7f.2E\SJ2JSWe_KW-5Y@Y&8JLWU?Gb/bKR9VSO=PR770Q\McA+A8GC3g&@:
_<&Z)KH[+.INReadF.O1b.;UB_LDIGe_+G#W.eE7@L9T-G5-cK_0]STf]HE^fO&4
08V_<[SRL1/T^G1Re95]->g=W\<XGE/G,H,2AJg\K/GO\eIA[X;3-_^VF8A#+X=3
<N/8:<1I7/G6WRN[4fWK9a.?&UdI67E0B5<6U-fc5cC5E16a]>X=+,2c4-?H<8)M
:J_L<\T(7TXa0d^Y1DNa+;PQ2M.ZCJUW-L_b06E<A0UF<<<Lcc,FE02CR1AD,;ML
C8a_^Y-TSLa]/R?<N>+TQS)?B-94<89.cO(/V^)A^I>2Ma.fg4U-K:E0>4T+baQG
eM;;aQK08)Vd_g>2Ia&L+g_c-b(9S))4C(OU/5bc+RbL4.f9Jb:1c;M&]CYZUS&@
>+fN>K(>a#-VbJ>@?SS?0XeAP2EgEeZY;Lf87aa1O+<40/.UBFB:[R[URM)6=?Yg
P3b@CXdO9B@?O9U^8/HVB[D#QNTMb96297_De36]\07E+RZSR@5BKI?aI(d\#e5S
T^3297,OY^DNQ-MV9cIR<=XM#Y&LM^-QJP[CN/L79aV3G2Q?5FCe7IQ>YWU-;IR6
.A>B[83=,?X]YPb-B,;,01W)#Te<RNSTOBCB.RT2YBaAPGCU18@EDSGBKZ8E;[>?
68/OR84L44Pa&?PI7BB9<9_NgJ)HO>R(:R+07K1G7RT6,W?bFde-DL)Y(GCGYB>D
aII/e-S]aEI?SU/8Z>G_XY/d7@@g49GR0dfG5UUg<(BS??JWDV_KDV#c(gH&CIdc
0fK]Q.(.?[e339971GS?@O#_?&<X#ND8D?5^@7;-8L9YRXI-<,C/8+S\Vc&]XQP]
b]A5T(G8WEZ&5+V<A&8EZUS=41:)ENcaXX8NQRYHXWa(f=U?Qade>Mc7XDDfCaKJ
(JG1TE\P:1A8#,;4L/]D<8eS,aGG^=UO&UFN?M5U5&Ff)KS\J6.QWVc-&DTPcb[+
,M&DX+g^Y-8^J==1FJ5\aOgQAI6(;-D9U&7.?9-b:\ME^AUAW>4Z_40=Q?Kf?SSU
:YHEQ),>.8fCHQ9OMF@Ob2bX1.?TW+N,ZZ_6bKQQcS7+_dd=T+?b=7G:GK3ROW:T
5/0P&Z6e(CI9feY6a\a55f#CQ]7A987,:c4YB6/#GYcK9BCGKZ.&1Rf\2X&A]Q4,
DW&)1E;_=5aA#aU]2U&B2G7==V23MFW?=b4-9\042.QTb\Ng6Deb&;HJF.9()=:H
6:0NP\+DR9Y?a&6f&EAQUW&bVbd(=-Kc4]C=D@_OLWU_IROJccN?4>VaEbW/C+@Y
fOA]=9>G&9>W8[-D;B-FL=b[7OJ#2LGg:Z.WM;-OW\L6a=F?d+,(N+CQ6XTD29&U
TJIE)U=aO,[WHa=gM21(c]&S[J71?B-]?SW>a]#?B;V?&f/[\/,H6(5e<2L,YH\U
>B=@bF,Y]1&:AL^RL8L+1+\bD:gFKUL.::T0_b/d2aO2SGf3/L;>M6>6Xg-+Y[G\
I;:cCAJ^A11?fBP7\9,,26JW3)4C]SM1e@L1GXZD:6H:LVIXeeASg_&f88KP[+1&
W0d=&LMHM3Ma-^RL,#ENG@(-YKf0^f(Od9:@gM2D4>4ZQ_7MU3IB-))LM/aAbOb3
6(#^dOeA+S-4c::TR]U)g?K8#;/8(Q9?X)Q,USENV[=B]Bc+K3d)DTD8Nf?NT:)@
c_bLf8;Qf^\0#/HDW=cTQQ3[Uad.0E>J=/M^1+T2<2cb4CA8VWcED^V2TRC]V:SY
U?JIgHIO+GRC3ZH5VdM<#Yg^>0Z<ZT0IF6d?<J)+K3]_F.L?MC5LHGFK@_S8AaG4
cNS1d2V2Q)f+.,=JX^KO2[T_6&B#/_(7:^;CQ6^#VfWI:\5Y_0S1:P58dVI@.2O8
d7HQ=W=\)+7GaSfEJT?Q]HS#_f-.JL[R-,[:YgM9f4O,EC3M&<U7YQX2Rd9I)eE6
3R)SB[f2LS3NS;[g9/]X6J(\A)X,UeA<42&(Q/R-fOfeaG6=YBR11M6dFV8(f2;9
Q/25PDT1d7@Y8@;O.JIXSc?+-LX69,P#J0#=;TaY2HZKdYJW?ZI@Y]c]e/d_XOS3
TAc&eFOf7[<L<Q:P<@J#T.SY5;3HIKUOS\9?Z/,MAVCaa:_cW4A7)4AJ1K7>TX,\
a_4WDQRW&>d<aW>?@Fdc7[(12CG?bY9aVT60H48a&]FSZ5c-4G5O79F8KOWdO&,P
PHgG8O]QG]UKX>&5d_7J,=@;fL9UE\2]OH@P0=f==,5eeOG@KNHJ)b:Rg,<Y[AM#
SVBB4I&18M8:=6cON3\(+=19B^Q6(cEMRY2Cfc5I)L#E8I/.&OVN(\cI/3_>F+c_
3MM6C@HG&))ZTe#O1W=K.Ga1aNe,BWDd@Q?e=K0ePd7;:eZZ(67C(Q2DT#=1&1US
.VaHEMd_d[3bQH.:\\5H-<?Kc=W21;\HJF?-X(+P)>S2=;R91ZZM>Y(O^J_?MD(9
8RDX0cOY_L/N[GG.SL>^UU5F5?SgG?&-B>F\4K7g?4g2,Q07CGBU#L70K7^I[T(O
R[Y)I)Zc(A)G>ZR=0G,BB#@:V[eV.:(ZRB<V4K81fgQ<HLbIga?]1dSIg)]PQ=_K
M5KB)b/N<,^X,^V:N+H@\.T1?=>+bSI+=V)VTLD51gUEZ0G\^>-_Fe3@+>DFJL,G
IR]4\_]M^+O9;F+,\-A:T4cRf1NN+F_.7eUPW2e64KE?KcgE.N;Y7M05H=[X[=UO
(9L.VFR)QZYFTX7#Q0Uc+SPN1@985gPSM=&J:X\g)Y<K?f31fYC+G7@[95_QSX@V
9WNVfL^0c>Mb4N5MW-&22U.U8E+AO4eFSE?+:P72\_T<JM\C207WH9g:;@TT;B_4
a+5g+>X(90gdQY(9<#DbC?BH)\AbTN,;-.eLS-]bg:bK@dcd-7OYK,Y:QY7,<PD0
8?CJAO+5#]/XKOH<K7B7L[]LGcGWF?2CAI;P)JKU>38.)6NVUQ<=YC4ADHVHFRSg
0&;.]X#_-FA^(eE(b:W+G+Q5^Tddd7;1X8]@-g#ZbE)ZL7dSYGHcWTNCPB4-A3_+
]Z^R_6=YgbFI,bSL2(YB4#D72,4Z=\19&6S2C[0&71&36QE=MKg&L=HNVT;I?&CK
OKQ,,TGW;d[^]agKMQ?W;e,eSfD63@Yd2D>Y7G@:MV?COPLA.?0TbHFT+Ne+I3+K
@=(6C\[1]W:;.H-c-GKH/XT-1BQ^9OW&2YVQ;g=5#ZN:[R#IBBN+WSGO+fUKCI9/
77VeC+OBe\1<C\4fb#f0^g9[4,>/=X_3_^/<c(?F<THT8,9_.OWTW5<6fg[,PO>M
8fWJK_53&c12>_T?[Ab\@HI-[]F_\J>N)P]V>[)T-=g/L[=b-(^(P2U_).;MAXg-
&2D9S/UK\:4YNJgaW7>?Q_b1[DedYUL>?JJfJafJBUVMMC/J1X>-+]QLRId#;;/,
5X/.<HH-TSELBC6SeJU@Z@#[DHU\_80:Y8@;4WS7;8@[QMQHI^RDc9E?SKD(c1(+
b+f84Oa^LfPZ0f1?<O,YWL4E?2YG4HE.Wa]LH7#OEb?9ALH5>ADP-OF>)aNf+#>Z
JK4)G-C2?2;G/\2\#Y&_;S357/.H]@.?Sd0OAG,[d;_U=45P\0=#Of0T6TIMQNC0
J\<GD6CMCbEHDa#\Pb@3#NT^B9+4<54=,DW_:T[N(CX,dCKAM&SX+RXZ)<<Af>E5
FT3-8]+^b.8XJ\2,>a(RPX4,/4ZOUg>^@#&50-C9SWc_?.UfSR)KdTV#1[C.PMGI
6G\U\@2FQb1Q2L-R9LTQBQZCH>CbAE,d6eHXb\D/:5-6LR=XZIK..7FY@WLM^))T
CO@8bF7OE@ZS=@=_O)#2fT\F+Wa1S8XME[NG-CM#;FBA4X+KAE+@IcR_Og?a.4F1
Dd]VFa5=\BB09G>W(R;/@?HJY_)XWd99IW6^;+7J_9C6O^^J6Yg:.EbAU0J>1(UC
[\UJ)4V+Q3(17_GWJXOHB./#4<^JXL3?#(G6Q6;OR13c;cLR)70_e\O.(N>bJ9_U
?^Z,/Pf=E.5^6#>2)K\UbOUZ@1MEW9PD1T2W<,LN6GA:\fMbg.@:/89.&Z[0=TJ5
_,M8YZ7J>P+,+NFadXb(S-&EYU=8V:797L9YZ#Q,Aa._La1+0F.,Q5A+-[_@Z#dE
/(ZS8R##A,W?gdRI6DU/XS?S\0SV1(DS/Gf8gdTQCeUY4UNPD5Z0J(17@UY/V/\Q
MWOK0\/8g=LL7N[/<XBBfX,D/@]a\V097?:OFGRN0b_b;0+,E5SK<I4?9CR1g^=R
:Y257)^(7dI:(^b]gd3<XA#8PAIAU)7K)5?8]0,c/XT24)4E]K?A@WUF9<g9e6&0
Q-#NbZIWM.TX2/4EcB;77aRg/-N&0cTf-T+J:2^-2_LQ;,B\#X1,0#0#SC15:SZ)
ZO;TAW4N-94ga1RQa&,[0TLS8_WAZ&MB8&1.V]YT)\;dEBgc?NDKFE7&=G@Q2OPQ
Le04&b[Q;YQ?:,[Ma7.V5g,6Y0;<+99T<eEAPO^L>-\,c4E,YQ.Q9TEg3:6\c.36
B\+<Z/&6:,<T>G?J11PG:QWAVAC3X9_R(&#L<(Z(g0V_eE/82fEK;O7<Y\P/7G7f
_HEH8?V^f(A2MRV6bFdB1Ab@VSg95E>T0MM0,R/JTG^ca/YT4ATLS^30QMa;@5;K
&W14T<+.CdgU;.)<:#6-Q/_08-H1+<bSaR</>,KM:-fLNSE\(M2g)(3WR)0]9fX-
]8_Ga5T.FZ?34:U=[=4-cYG1)N<YL=XD8I:23&72O>U</K@-?_5Neg.<J^2e=\.V
03-3>-UXA#[3M+[)b-^&(H:Q7=b&(?U@Mc#Me^BUXF_?/,J.RQ(-)b(^N0@?OWS_
2FBX?;D5]J@8#P2O?AY+HIePN:JLV]35(_2?IX0.AT4YS43U1A:^0@8C\H<TL-&8
W)-1&^(<2cS4^fW8]BH;QX]RS<.,4<B&92W8-B5\TBMA>9?XB]998P2,TK;UGJYC
N4EXRBd2Y9)RXM9#5F<S=/W+7WZb=J>@#R0Pe;#E[#@e,PaPBJdI@c+(3QIIcR_g
Vec:J>;]/5e^Z#.g=-\R8]FJ/J1,<eNWe5R@@A;HV7MN=>E3)IUD.QDP#9-:_5)f
\YeP1.@ZG_/BUWgZMdR(E#)F7DfL5I4fg]09&MbDA,R)K5ZT/UEK&XFESgC)##E-
9.6=JYgg?_BRYM59DT7Q4[:<\bB/M7Y7ZU.<8:a4G_g89H3ZZ,X5CS9+R6Q)[gTJ
Y3PE+6.U8W)\4@(>3QBL@A<68Z[>5Da7T:SMH>\BIF>O0b8W+K#9FHaMVg/)P3U_
b3Z#Y69@[NDc/0\O)>aA0=RBJLIG.WB5B:1WIVRZVQSc\+g6AHgc75/66(:;R9I&
N_-492f=<RRRfRUB2YZJ\#cg(fW2@M^(<](EeD5ScIO0)P\T\HBMfT56?@:O-aBV
IH(8A7F&Ted@9TX83LABFX&6.,DZ1RUB@K#eWV5+0cNO.8192^&V5EYd^JQ7AK(d
ZG_)+-_BWEOFU;JKLTZ^ge>2JS[e85N;.\cJXCX=L2f,JL[/Ve+75+c:;;T\O/U/
^DY93)=O26D4d#P(>HSPa9C(Xa=gW[6+^BdZ(XP3fE^LY=8/S19<XZE@cIP9Z796
:^-+3<5\a0&#]3.\cb-P>?KXMeBC)4?PN#;DWM(XPSPJ7fX,8LVVd+XKRM_a+:WF
J2eX07CV[+XX5OMOU)ASHC2-O,5UaHZXaJ>4B47WES:PO[#b^_g]g?3-K=0d,:/S
@?&UEEEPKKO@#,5LGbTH#?L++6,\aSRMMMUQTe@+P.=/B<d2PZ1gI;J8?B)aeITV
,^/LI.K73Q^KK[](X#ZVIWI+2<0DRLG2U.-+_G:<9faG540+G?P_\dg[f5-1Zc=7
+-S42/OIZCF]YK.g+L)=0,DPH)^1ONWZ=N6;IbQRF=\BOU1(?2OL+g,1^P3]BS+6
=Z?G\R,8gVXYKaTA;P\,c8a7WQS@Y(+89=TIH,5K^fHD35;4b,+YS]QC.f0,B71@
W4Rc^FP=N:AdWe?D=3fGb:GCC.YORNE2B3+/Y3Db=5cd#HJ7ZD)\4JACN2R)5#fC
2F3NT->8)\M#JeP2YM,H-@eF#K;SPc_OJLL^PE#gg4;&,<b^H-VBGLCN12=d.CK,
HR]#1,)gd^LOLd,b6f5L6SeJeM5=XZN>S[8.7fa\P;_Ed:(KETMHY_K\BU;UCJY:
(aF_^1W)3U#;\E;b1#5TDHRMfN?><V)<gM4VU9M;.C_=9\H4J5P\KIf4+H6CHW-Q
>U1<FaG.c<F[SKIc+YL0,FLRCY7DF:1W&3=eCHP9Ge=+R9\Q^E7.?7D50B5#FU&Z
()<.]F-.=Pf[e;B@DX[],;cc<U4N\U)aE4feD=^V(C;XG3E.\^\12SRZPadM(T[>
(-XA)g8OCMXO^>a;Q+_ff5E3V\)===3O1YgE#[?AW=3>:)1U-b?0R,aL?02M&4IN
QLVST&_H-1QIcd_a&44GD9Nb@g@ZYI-.6begBT7\ZD,B\-V2<E[DA0.BBJV,?=Y8
RF]Y0M=_T2<ad:IgLSTS\;WC+)\BI;=B(@RT5^Q59<BNFKIGWQ-#HZ=H;F4OCM27
>JALT6<agF8R)[acU[5/9KZ6)75-HV2e=35>->9f]RACeL1Hb+d-g-e&2BIbE.bf
<F;7H5^C3g.[YWZG.T\b0L?=;:@Y04HL+e4+X-7/<X1T)QQ=BJe;KROe[H7&:MZ=
b0&df#Y?eJ4(3)YK7:BPdPO6D6R2?-2?D2I^XX>QS(=&NTBI_H(;L+PGe32;.,_1
IWZOZZBQ=[D@V@KY^eaB@BDW15R03H2?6cg5)Kf:5\H[IbN\25Y58&<4aSBH\37L
@H8IbH1GYNB2-DO6FIL-[<^ZJ.NdTW+(fb8Oa0&005Mf_e0ZJS:\QbF2[T;N+);?
M[bD@JON=;43d46M86;<SbbC@^6PT\?;GHP-3]VffcQ1ZPU>WbKdXJ\=3CCYHLMO
6_.V/)4B0^4;H\J4RQ6G7-dEA&M\FUE:_J/<MN)L3X#DHf+BYa#&2-];0(]^EZf_
[187W0<3,R4FMB00]FSb#a9H]IH&9adV&#M\0.#c+Y[3=Rd,&<8a=ZXKNK24g:NS
KTQQLb:8^[F#]XV32^,OG@]#MBWRbE09(EPc)dM>SI9(I.W:]8UR90PR:IEK@XT,
>(7G0Jc[gUSdD1WX.11UFbC5,H)UBcUdL<7X19=9O[5+#H[cW1:2).gN0\(.)N@H
Ge=[9=f-GB@5J@Bg#<?gE_PS[]L,NY.Gd)9N59-O6\BfE\\R#I^03D9ZAOFDXHe@
#79IYXX7QdHBLMV]PG+0\;U;^BA&5JAcF?^<Q.MZQIG?SECI#aV/M/-KC@4e<;:T
1C3aC0Q>3V2dPP&.)CNU=4GPbc@=R)F&X2;(([:X\Ndd&Hb2-WVW/c?TI4Z)LY<b
))?[&(f7/F_HNHQCfC+?HdF8Yb:,D&K)PIRF@b7BEB<.VT?5J/Lfgef^W#U[#&XI
APF<(AJP^V><A76[&+4W0Z(06dc3J+^/LCB+e0g6__#g;&Abc5W>)=]3ES?gTO)M
JQXE=a^cB+-PA/dd=Y3X&K7[1cf3YcLS\TJ+b_dAU-gVfZ?B)QgO0S;Z?B7,=#W)
YB^+)eJ2K69::c7&+UN9^\764_/ZD\Z4S)G@e\RJ57J.TC_;LZR24A\@AM0A1)W_
bV0O:[N\EWJXLg1.RbO7H\L;W]V&<?(cg^E^ec30OXFe8+DJ1;9dKJ.(2K]/P#2g
J;B@WB7SFJB@PXW[A4B_J-DQF-(FVNB:8+JOQ:YQ9W8D#LHeSRGVeIN9/DfD[XaX
,A_/NL](6<g5#cI:VL9BNFga?^L/^#<5EF<WaHK=:))AT]PD:=a@2RZ1(;9VaVF[
_]\GU>9S5NdTba)[L2N_K0Od]W1EX0JY1=9X&Nf9N;JJ1d;2U.WOR+Kf:,]050R<
=AQ0Ag2ESIATWAd?F9.^Z2YL7:^N86KX0aaGV5EY]C+[EOc>S+#8>H,UZ;^#+e[8
1a/6Z<?#gIfS)53gV6BDH+g0ILLWUb6P5W0G)53+^>;-FFC_AO#I8BZ4JO<EOXgc
Z(AOX+#U[@LKZW_V<YKcg@ZZ6OGW3H8:8[<4dK.-QQSJ)FIH1,7,,<#)H55a;>B^
IYNaA5]NZ-7CJX&7,c=b][[6Ge:1JU3])46+3^ZG;CW<_9;+BGS]LO=]RBX?HH^O
QgJU/I\IP\@OTR,e+\-K2^1ZcWV[S-6Ee@T\WKKYacY,<0K^N.[QP;g<]A]0I2cV
M1G;\[3bgYAU5SPKQ[:=-aPb(ScaEaA0VKAIYU:Q>J]6CbJ99<)95QCFbT97^@U,
b23Kd.a#/\C?2+d4B?JG]M&aNM]P4FKU057P87FE5H=\J1b?_[&DcYXB@<^ID-Yg
CP00R]\VA@+3E95H\63D8/L-&DcA6\TQXgaHFHg^gR4]9RbYSdG3_6<@XEE/aA:J
8G#O>.C4I#4PL,LPa)KL564b>O:F1,JL?/IO8)U.P]+KR<W+]/6Ea;FAV.2eNGR2
I;[c9A0@#HSWX3fD:Q:Z+I^C+/4-@C\JW1KK(=1G0S\L(_+031]f1QW7Cbb@_XO:
+:5)#D),#&>DFN3WXdC4W^ZM+A&UC44B],YGU-,=d-AKXZ\:5ARY]HLI)&X=]/[A
G^K7fGg<3HX?)U?28@F]LL1b\f,<FU=DK[;:>/&)^_-Ib,HQ/)gU82fg=MZ?]_+6
<.eB?-KJC9#Za#P7-dS]-GV(ZXbceg/f)GgU8-XRBH2)O[BITB)[\.VG#M&8+(d\
1TBO_BZb@G81HQB[N/K#1[dXJd_[/a^Q?HXg2E8f5?<b]8bXdEgHbfddSNKGC<4(
S)F(\JbX8L:9-(,1Vf6Z5AH_<+DC:H0NIDDR.<Gd_Qc6c/R/0&5HIbL?=)AJeF\G
FV@5=1JGVB-JL_,_fWbBK2+CGA@NNeV(QV@;/FbIL?b@&SaU2B>^_9BPRe#T_TBS
((_CB4;GfbV\)(,L^6;a,U#A58MGV<EIN;98R4PDGAf0+(D]8b18BY[0<NH^X=(a
N@d&7b;-^6;YV&?\C?51ZT/3;R/EPPNY.KCg@aA2MgRF;QD:E\:bI6Te_&72)fVc
Ca&/&)XbN7L)_HRF6F+:VP:?55=Z=@=O(RH0KMDCIGgK<3>KfYRU1,=XMD-c&[,P
.c>#,5KZF.-)WYM649EPD\ZEA)c3)2gbVd/Z;\O]b\7,1@RP4)g,3-g:9#P0-8WG
0H9Id>QaMZ;3?:TPZ:XDQ\@/WT@7?d>9B,@H2I,>,RT0>NA5f0F##(TVS7+V6Jb7
G&:f2(R&FdG#9#KR&4P=;Gb:1Z?_&DUVA.bSK<;LC:5_FZ8.LZTQ7:#]]@HBGF<e
T1(e&^5/UI=&aTC?X[6(OYIGEX\DT1<dB;8DO]D+A;a640YOC[^I>b6L^+OL=AfJ
TP4U,QAJ?V;MOc_6.70LaUSI#^fW;2BDHF^H_a7?D]_WR([7[)GN.O<<R?/<7D.\
</,.0NPf3FJ\U_e88:gEP7(f=3a3IMM6gMQR8#M7;DI472A)ITJR465\&BXTd3S,
>V^;T,e5#?>RH):20#?\Ycd[,FL6J6O1NLI4Oa\AD\_7?eHcME36GL.NA/@Z9JGO
(E&9=Fff@]-]bS-6[EJDD@Ob6g;.#]HMPS)1fWbXdeVg<I)E0LT5\&9I:g/RW&T5
-A14X\N7DKPU+;2Q5&0b-O(@>&dS,A;2>]cMYK,@T=1(^?K9YEEfGPI/Hc3@Y12J
A1e8S]gMPb>W<PO.7#CEbK3f;PSa1JIRY8Ca@2^VO?f]bH>R[H#b]2K+<S]dcbIK
,);^16;C8,R?^R+OEHe7;_?52LLaU(I&E1HHV7HQ;F;UfD0#,cTUgcS\IQ^f^J5A
c.MC^9[EeZ;;dRWN[D2Zc+gYbL=1:c2X6EN@FP/QEYVK-SG^=g5e:L(8?QeIJb_2
S]II&FeN-NK\gT<O@+(Z;MSH.B#GX+?NYTZN=;fbId96JLUc9F:FK:8Z^G3Ag:_9
2b>2RH_0eBU<2?e/-0,Y^(R5?_/D97a(gRYZ3WJFXD.5)[5X==FE#\_5AO=@[SZ1
F9cX:B-K)QZMN=fK6O2G8CMD_)Lf_<f1A0[O46P2Q;&TQ>0]ZMB5+QBf=^Qg+gDT
:C=<8(OcKNBIJbM/FX8,#)C(+IY.7Q;Q;N&OcLV2KW3KTX4T:&&geTQ8^:LdGIO5
-dN,?99C3=FY/7#1.R?83^-fL?LZBR+.71cL.D[]eIN[U=Y/Z6A\V6Y[]@ZdDDY3
9K8P0bc_IV[OTeRW)RdbcWJ77&L5+9\Qc=W?:FcS<Md@b\ee^K3<V7O,fagZP=@Z
QQ]9afc1+2WL,^B-Bc(:#Kc1KC]>:/NM;.3Cg:79?M;aXDX:1.HfAVHfGY26;N5D
-ZNR(:0<Pg6)6M-VY=^-VXd?F@9W:Jf6LBQY5.@@VV\IS+8D]+(ef7@[7ZG0YQG_
QOg\AegI8?]X<#dYbS=aO7(-VJJ=K+2L;#S/FOdNV]GB02RZ3[,E>HA+VUWIgUPT
T7V47&C9:b#AMb.MZQ#,TD/O_R1cEWa^WB??8Oe:VFcZYVYe?dPY+:K)E>&@V4d:
^.JL6ac,XH.Q?7NG\@B#WKd9P7d;RQQ[=3NOK>1&C]2)TZ1IT/af<O03,:f\8;;I
5BRC-AWb7-Y,b7H-O&feW3a<EC]+\/1IO()F5&0SXMU9>=_<7e=EaK;;S&;dH_A(
#+b)&3WWWCSHbH-SFfTGa3)NW,LN\R@?-[<A4dVH7@EDSY[4XIB,Z85cO-c8DBUN
.(H)b(I>R?QE&+.(Y)(MB4#1E)YC?#]ME4>P:#?f@BY5f9JHFC/J&?]7CYRTc.Wb
H<Z(J([fPb,63OU)1C)30A&T<TF\Lg4@4O7:&.HRH[Y@IH_B1Eg.B/WR]K9a/W[7
<aVD=8/;dMK^Sf=(-+^Z@e<R,4dD_gUNPHe0d.4CJW1,]QX8Ofe=84+e<aXK<BCa
1Zc4PLFedNN_&NWTZ[@bN5-GN[-F)WfY?,HGJDVfa(4H_DO[>L_<J..W@C/NXA^=
?G1WJC8JW?5e1-WQFKK+@.S7bF)Za]:[Bf(XLQO65@S?-#CfQQUTA.Pc4#3#)\5V
\U_2@CNP^QYF?=#IY=UKLVdFM33R+I&bc5(VaJ#&1DS;>)7VQ;O#bSJV_V)eH.UB
=U@^7H+,S=,@N>>MYM3-(0#bg2,3K/#RXRHU8S_TSY>@(g3e28Q2X,5T4?P3<SPO
FQ+G+9R3X.:PGT0\bYfQ)@2WEEBgI<^)78@Y8ZBL7b>E1VHF1>2KS6VH+F]Q+\Oa
cMNV)^G^b@)L?g(]1G2RG5,3A=4Z_0S,0g)Z(LdU[Tb_K9?.d,]18a[N2D(Q:eAg
+Y]^Rc+&[>8d(V-P@-O1TXBDP-Rf:d^/O24Wda-V3DUYZQ>\ZW<gH^VC)9<8;8?f
W5\7._H-&F]e(@W4)4X_1L)[,IB3W#8-?X3(OVabQEgTFgU]CDc3\?-9KGdBX.66
7JLGLc^Ie\:HDcZ7O@&,\ZBcE]b-M=e)bLeQf[H1:CeJ@VK5a,Xb?8T.4_H,U_O4
,E70-YCPY>8]-8_E.)P.aBE>5WXW3>2Z0ZYF/RXL&<DJ[a.(dI6EKI,aY7GNN8(&
,D]Z(@RDJ12c(Gd;c&)QJVO^D55M+g=_\QN93T<_G-5PXI<\_]Ia5ZdJ]BVf?Z\=
[2>8OBL+\a,/\W)ZMG_SLaARSB^B88gNH?;+LE^eH3^[P_826<Z?1?Q0;Pa(/9.E
-GH8>H0(NNY#=/D9_BEW04_LXbC/Cb:)=APM/G-8/7a9MF;_/8N4YPdN12gJa:<=
>>[CKMR,.W;D[[dHAJG/23f869FJZE7;BW/_G6eM[GGDN_P8;@U9]cQK?D1H0[BT
;O(aT)>JZ=XP/BO13S1UR:)QQ^,F#,GTZWE]bag.Vd02T[a5D=40[fM8gK4R)eYY
/JS?<_GZC<JUeDQf)&ff=3UQP75ACX9F4/KII5eNT6MacC1BVeF2<T>LF@5L.</B
3JGS]VM:VBP?=VQ-C<&Z/UbWF/#cHX;I.+=c//DM?TE[#e<8,M<AX9c=YMI&eHWA
<bAOgIP<>gDHa<_?,1>g&BRR\EX(d3g(6MT?a=B+CP\W:>#d(eDaf;=JVW3E>Y#/
FOb^eOTa5;/F,f90H=.b.-?d-AK7IXCP1,T_Y6)eS<BW6=R6=99S7?G+T=JD+Id]
WQAGfBLD64^C15WgJXM[#eQ75f\(]]C@)5+@E[[FEe^fXSG\Ggb19aSQGK5a7?B1
6D:gW[_;D@e-eS^=;\29J#@YN::eND?f.PA7.7(7/\H+W/9;Y^C5Q=@TO&EgB_0R
)N4NQ^>bWNAg.Y.Ua<g[Nf\<GV>X)gBJ41I#_&=Bb9M_>-QE61cZFM+d95G8]HLW
bH::6,f4da8FKY12@(\39-:P6M;DNFB\)Y=MY=<.&cFZb3F95N,T9\;C=5fgZ+I1
PCMR;Vg@;K@[T:A\)b,:#MQJSTP=<JbUddH/W#cdY;a)Xf[+@VbR;=OaFcfG&2,9
0(=1DB@4fAXG@_6ML4O1b\NeedR3R-@4R(SQT,JN1^[UX;;#9N+2ZH;=8#fabIPM
<8CJD3\eHfZGE_/YL@c-NH@1&4@1dI#f\;@/c51M58b_Q&#DTW8DXb:Ag9/H0+QK
d&:U_aUEU[+2C4#5_]_][fVN1Q2=+2G0E&1bRDQAQQO)3C7=cXZBg)P3#U/RJ,:M
\V.>)=C+B0<f-aEg5MTE86J)(?TUGGgEH0KY5L-MUQ;XSS62PeT2bPOLR6X\3dAH
47cY4]O#,.<dB\DRO3Kd2e2S]M#ZJ]X/B-#IAX:C/C,f)@4_Jb:K^SB4SeJP7+8O
<(e;UbW[R\2L+&Y>=87:cFc=VIb&:06Q.KICO2H7QLTHN^)+U@eU;,Y?;eUa[C1I
2W)6dCVJFX<>9+09[F(JZ5aI+J9>[ER4;[=fQf7<2W[V+Sd3PeGB>AfBH^=-VYZ8
AP)-]M,ZdXY:TcA;H1N1(WHPJST&bD:=\ZY-4=XTZA]648dW-#T&g7N36U3K,U4]
[Mda\LAUT^_OZ&?a3b7\;^57ZKCe_?Z-fP\PY0/I89SDaN9WC6IB7LW78)g86EF]
f)-Y,D..Q>\BfGY+9Y&6_OFOE,=-_K\;F@OW>W:GQfZY)_PfP6)BT,=H(M^deH(L
2[/]fD//QA[AKN)7Ra(P@?3bIM=OC&N[-)QHZ]N@Z5,@UC3PU76a>TQ^+IO2OQ],
Ba_WR<0gZd_5PC_Wf^0ZTCe>]><?S:QVQY)?ZMW+L8]R)P4LJ9]@)g3#^.d0#GIP
UA[23Dg^M,GJ7FZ+SC2[LQ(QET/C++d=Vgga>_VP,PL4/Ma)7G\C/YH2@^Pc1S)]
(2LC(-S&./G1^MAJHdM,1Fe:2+,=Q;CB#gZ2T#:@WM)B9;L[IJMG\,Nf>fZ=aE\=
/&LSdb/8F74;64&HG+Kd8)5C^LIUCS1a?9]K\Q,1eWB#._4gCc.d7;A+d:(7C0\W
8(AV=(5.1eFg24R#B(NYgQ#G-WW>[N,eW50-ge5Y;fGUF,bK,B?Kd@aU\UcBAaT\
^fQ/JR/Q1?<@[L+C;9K3A8dB41+IDRLV,NCTC]B/=e:<\RNfM?5g>8WcKX)7G;b[
1IAc&)JJU3M,@<,OVaA48BM-D_ALLc@A]M80Q\?_Z]#:De\-/-RN@BIXWG.8e-M]
LWD6E0+]CJLO1PRUc)bAAd@HU\#4W_.S\X,]Q[/Jg@)><@W?:\Z0OC0HQF#R/N7M
fDNa#BUO_9BHUQW+f(FWFH34WI9NK?O4X2@d6?R\_@?XB&.:P2M;(K8agVE3>PLJ
64DJ]eV/WfI4dMgFaJ+5eO0Tg4RQKX+c&(9PKQQ;PN7PYAJdCRY5VCbLV9-F_.OZ
/IV)8815E3TdB=+J/@3+V)P4JbDdc=:^/HQJAGB@V1F&c0Y1,9BQ)?M3.I[<J9g)
1UIJ<JXeK[H-XGDaGTM8]?;_OH>W-AgN[5>RTI[0]YcOME^M@\^Xb\4P=22a_9JV
e\]OI>ALNf,BX^\LdNQ\[#-M1&Z#P?KVWaASH?GF+ZCg/^OWJ0&8eW-:8Ob)P#MX
3I+X1Xe82.39P<HcU&\;02RQdgT.<:5VLH;<Y)Xa;S:P+6F_ZI<B7_?K<<8S^c-[
9J@9Y#Z&g][6A^B_]DD:f78:43KF@NQ]48=agK+J5?OLEW<,cC_UUC(BWMK>6@g&
bZf9(a&=EG?[ZaM0XRV.]_&48J53^a(]H6e/4,HTAYD>3T&#/-M58MJeEVVHEbc0
W1>,]1b,C+D&2?NS:54?_QIR_[ZFY.5M9NZ&P9JO8G-Y)+5P01UJ/T\X]XPaPg@^
e\6aQ37M^Q2DSN0aNQC-O+FHZ4_@?KWf>gc)2.\b?2-Cg=J)]01b9Z>Ta)gUX_J\
aK2<:W4T_M;B0AO]f)CFYEK6C4_7b8@X/:8V&092aT).U+MdKeZ2T<Ea[-@?ZWe5
5EF?=5F&/.=O5\TUFfKM3GE@&X?:#bb+79d(.5,9?:S+9XK=>/f^T_4T+I#>a_YS
+G/2/Q(>4U6fd/],,3],6AL.1BY>G^6/&HV9)X:KA?-F(]8_Y7(a9S2C;I\cAKaF
4-62Df=Tb4D9O/#+BLF:O[@^TQ0c2&gG.<9c6aLV.#RN]1)Vf,YW7A16bQO.Q\P0
.)+.dFX89<R/Eca1g?BFWF.HH5T:CYUZe9A7VLH_AX6-ODH=7L(AF@\8K1_7^XWP
CLUD.<TG6H3ZeS.:f:Kg11GQ4#JS8?)DE&BIc.d&6P@PO4L0)L80-63[7/W3AVV;
A3&2:7P]WfZ;KK]-5P\K?80V;B:Cdd(9/1?D]aDSKD4DKfO;E2b[,6)@^@KeL28\
G>2LSJ9I68>^PU-J_7@PKXf9gMT6;EM@/-MRH0a3U^UP1W0M,PKWRAbP)9[DN&P#
3IeR[3dL>UQV]VL@GF<IbOaJeOTDEO#\\b;)#V_](eEc9_c4/?XU_g_?;J0XDcF@
ML5@AeHZaQ7b2GG\4(YM^bW:T<HANKQ3D_X=R6SfE]S7g1.VeW;HB>J&;[4HY.LE
EZYR0_TLWJGR:G1YWK\52Z-,.MC/<f(SJ9@.@E(8FXPT_7>?1=_>:5)a@PgT=9=L
>D0Z&1@JUeC3]F(c(Se?HTf-UbG9#U9fg-_DbI[D5DE7X3.I&6@^Q<5SN#M;DM5.
9E7IV6eI8eZ<Pf<Y,8+?b>M/DB,;7CgdO?BA65QHeS,WLZ;,^.\MNgJb+)JAc4L9
OB2U/.I2Y=X_8[^M^MH7;]gE))M;@E?F3Q#e&_)^?NXeRB@_(XHT7#UJ94N\(^>O
5UPLMdCd.T+G3;0b0#MI+R=05;^3V4Td(;-&^FS.=F1@V@E(72+6R/YWXaI]1.-d
TNOCY1E-=-K/.:RW)c63M,fS[I_+5C=91_C#)d7egT4bBJY/5,#P-g]@g]HgdUaZ
HS.5OYI>D]5DM0dZ6bg8\:GdQeCDCS?G(EK?K<bR8?)K.[?FP\/;cgee=.ZAEB2]
K5A:</g43:5)G#g)^Gb]1#L3Nb/U9d]46QR+a9c\Y1Befc[Xc@P=#)_0eS/R19:_
PO+3W(I>0^G0QS&#-0/IP(_b-&>?VOIc#B5[=U<U)VQc0:F]H5UGVaMe,3F;_Z3g
eY<6V<2,8>AGJK64<OE2IUX]U7P<\d(VQDPHEHFY_OY4VAXKaIU2X&AI;R:b3CSF
[41e;#U<b[R=90.F?R&:M@5?N6^UP2N-26_?AbEbM.D>Kbc0JD\cD\:6(fHUeQ&f
B0W_c<9&611+IWC60<U._K]bC4BAZ<46dK5SESc(\F+=JZaBf7FSKI[/UW.26\)9
O^7&c#MVLK:N<=RQJA-3SJ8@G54K07@QH/8/DJSEDD>7?PA&E(DT>C[H4]76>M).
B?4&a8(6,7L&Y1^NE]=NJY8:=SN8AH])J5:@=7I(AJ<6,/YX@<e[2B[6\2I37aTA
2/0K5B5.0-[c#16S2&O&RcT8>^eKWIDUJ)G4)Y+24;Z/LD:G?W[<<Tf<IeEBCaA1
(G^_-1aULaUC(4dK[J0L@DbH;<Z(?@ZS3Wb#c0FObgXX-]JJ1-b.61_S<0X\7+@N
M+XDedVXeNf]4#^,]gRTG_Z>O(@5Fa5/W#DVTO2fdMA?)V[[H)1VC,Jf<<JEWd[E
HW3993R<a5UIFCB]/S]OA2dc)2HWN4^98e9dDU9AB\DR][ZCdaMBE5<8)>ME9fIX
N]+\[-(4E=CO5f-)d:=\)EJ+=BVdZ08+TO):66a(/;EU=Y#,,b/VVJ<1A,\T_6L9
4[9.S+3;O;Q@H&Y[(\IH1><:0V;-\<&D?14LN81M5fQKFW9ReQT37XK8C]L?Bf=9
CSab:P/-cS@DV/QKea=#0L:ZCL4/L6FdUC6eXJ(W,47NXFbc#[>)_d.O]AHH^TET
5^I^:8QE9@/dETIQ/W.I#0E#JeXagW(Q^CP&03_/F&NRK+5EOPQeCGZPY:U#S16:
#]d\#WM_NB5P2((MO6J6@-3b[H<7T2_;d&6AM;_ZT7T)(ZM@cE7-K7SCPH7>;0WC
Jb?cSRbCZcP0?AJ)OLX#6VaS.GE816CEZ<CfS/NeG/HZ=D7_,GU5T((63dB@ZMW:
d6DZ>&_6(O9bQO+-?KC\0L[&??[]YB#3+1D<0b:ARBf)YFdbcb,Z0e;Z+CH19>)-
)O4GM+4^4H+<45[X+0H&d5aZHZ/EgWGJ[7eE1W&[;-B&I^\4>g@&:,I6E(SB:H9N
d]e08B[_IA6b3UdSAZc6-#AP(84_KZB/7)eIe7@U9?;&DO@KN]EfV&\dWQdXCd54
6_237aXP<F.BXa/M9E-6T8b+BO=eNdU=GCHPP]<U?<OQ^4P4J/-E^F;e<9U\BHI[
?cg7^G-Y)Z38ATPe?;HDfN]VdY7+YC<IYI]P:?P+XACD,bDKN3RbCRUOH&U?4N=Q
AYJ#.VHA(M25G.W9V;GV#Y5a:P4@E4,PLdLT,TA84gc-Lg,YcB-cLZP2C9-&AgH8
7=<VHF34=JfC<.bIUFcQcXD3EP[G]I-[PdV7\#NBG.^f(GG=g((@]e])SV;3ce^F
J.+RC.=d(\O3(J_@(:F(RKEE.)U>gV&NRU4SIBJN\-]4U0U5P1MTN^SZ<J2:>e>^
8cfYK5T)K4V0bEMLL+2#CR6g6HJ&TIYUT\A)O82EYBVf1LAHN4K/Dg(cZQ54?C^>
6T_:QM5VC;T+f^g<BM4KMeGSCVCf\4aOCK8N#MIP1bA08#GG341bY[2L)O-ZB;#?
?[(Tb?MDeb:>?Z-86EI)6aI./XBMFLFAR-J8eS-0Sg^e@CQC(PBS-DHQ&&X3VSJ&
PU\YQ7UJ58WKbb0MMNf\Zd,4HG97bf&=bY4gdXVa=fDQRaM3BW(dU-EeR2ZXd=K/
V:C?VL;,V6^YEf/e:OSY2H,&]NHd=1#PWG\LP&-BccE-3N1IGM,Y/5&86gf1e(L4
6[OCABQ251HB:M6fO2L)^B.[A+QEZc^6&=VKe09L@9;02BEVY_HO;f(Ha<TJ401X
L<fa]dIYF@7N-;-+-+b0#,[YC:2DOQR=UPB^^\SDVD(aGDf7L&G(LI)^<GEKX.8)
K(EMX]fX5\QV&L^M3>-XQW<-Q3C?U=\J9M\+HM-/^F4TT0X>L:?bbHHYJ8<0QH8W
FP;M:0aegK_\[:?UUQ\RQF@@(&)^1]+d->KJ72^)YN+BgY)M98BQC,FPJRK]1>gT
KV\;JB]MRSaZgHC(dL=fB77LZ4[=60.7@2D9+(0.@(bYR8VMggb@4Y;KOb:,TH9U
8H5>)g4H0290a-[.8(V(&<JeZ:_IWbcHeT-L47)>1PG0FOP3=YX6R<<@FRR-M2dQ
<@AYCMV/,?g_+B,XPE[-;H)774GL\9M#TPfTZ#T+V+,0&gPT9/B)/YPX[PTKU\A>
?DJX?CZ//8WAE)V1XEEb,[#,W.__MWPFJWH.gE&bH)L/@gQdf,Kffa?-J3KK^11,
@RQKYRKf0+cdK\/(BLJU>eSY[TYKUQC\.:QEgRK4I-(X_+cDYKR3Iga[A\ON<3IL
22K9=cAD&geeR.)SM1W5V1I#:cZ\>C0Y62WTKO</_XVH3;^31AV[f4MKVCK.)K?I
YX-:<]CIY,<f&W@X0084Y-/XTC:LOOcRXVDgO_D3^+b.&RE2CGT__8g2D5X21N&G
_F<ROZE^]d/N10MZR3Z#^E(_>SP4c3V<3;ZG0:]&=>C<B/RF;bHFW2_O8XF9D3]H
<:UR(@DRM1Md#=BeEEM\@[4+\,d#\1f47;JgGV,8,>HT5I.g1PG<7Mg/dX/gDZN[
LL3EV8F0B)C5ORaQb-LA)J:7c@^1IDA[@bZ1@7RHA/FC+13E\ReW9G&GD5SXb[[g
&8_/.F69MU1((H&>AD4Uc-)6=J#f6Gd@TWA[[d7@W]=PXX-^M-3V;M1KZV,&[g5J
P7b-DZ)4Z\,LdI9ZZI7IM4gJ<G2)eJAI]5]._ED7M#QW6.=>@f>e6^C=(:@M4@28
41W_H;Sf8c,)#@L/?,^7e1^4Y28@I<=OYJ_;94-9I@FMMD.HBG4K2(X<YG[#d\AC
[a)]DK<9KS5gR\O3a6ZQ6<C]3KJ]/&4AI,GESB)+LaDQ5@+?.>bN4QCQ/US_g[fN
_N^.S)L5;]_Fc-^U++a,P?_I)5bLNd7Yf4VDEC>Y@G/57NH769_g@EPZ5^)=ICU=
,SfEWCHe&A#.dOY9>\/0&F6BSUJ1?Y#)=fJT+)P0C1VS?Hca[C@\G<)_=-)]YJYD
HIe406#=G&HOH5-7gVeFM.2@Q.]JgBZOE:2(YD/Z^JI^LQ5&W[dHbR?U2O#KZVTJ
</EdHd+//=GSA=9M#\CI^]aK(;N[d,K2O^OJU?1c1HeVaC(QO7CU]9C:7RK48.T4
4_d8C\>@YDU0<ab^.;[bZC^;]E=fOZ-<W-5WF+\a=8)-Ke=C;XJR.T)VYbFWFFJf
a3&:KUSLDg^4fY:S_d=7cLJLgP7#FdfW^Zd=e^^G\2&TPgP.CH<E_9.WV2[WM(\N
>P1;d>Kg<R#MHPBDXfdC/#74>)fD-OP8\S=W1/BSS93(CXAT8G5A?^8F&1gT@AL?
LF<^^5D=\d&L/_d_5=&P^U4b3Q7Re+Vc_eY37=QMY#Z[A(]+#=H\f^QRaI)7],-P
VWYK+.Vb27&gE1Z8#eXW/X/_^6e2A9?_e\J(AbU8GaOEH^C77IJO,#+I&>-S.2NM
aU4V36X.9SK3+T3.UdL,Ec9^(_RfY#[I)<(L;UFRE6eC;PN@I#CI9f,QP[21bUVR
NFAV8H&XGXU/>ICT.F;dC0T7TP:Q1,-_ZB:L,I)SAZ\?GGN,cPSef2<-NM\=N&OR
^VTe-1@X4LbbG\>cJ0;:D8\PJSB/L(KON5dIHHg0MH<TebA2_Se5,P@f15b_>Q=g
TY[^_c03-RUEM9,a?\d>OLPLC=:1,bQdK+cG?4WgS5gV?HTV&;ZfP^2L/H>HKaU-
Af;LP36fT@DC9S4_E(e32<)P]e-bS<c<[:.cF5W<gc<HQ\2QREMOFIJPL()+O;>C
<>:,WeHV[0C[OGg)X@U7Rf/A[>JYX(JH+[(,_9O\01HJ4Sc1Z7_P>7Q>2SL=YC6\
Ie.9\HAX)UWXPYE9=M=2M_NfCeP+V8?fPCX7S14U)#3fA_YcQe3=dOa_+.Z&.\:V
[2a(#@JN_?\bE<KJ/=5V5=5e:AQ-J;[dafT8255FFG25&BD^63TO[eO&CJTIa@E2
HFI;86[NVH^1PeJg^.Y&2FUb]L-I.SRDJ-0.?O1L0#)d.OI?UMGC+\?^O4eR()Yf
\^,?eM?&CbSA,/<@M#Y@CT<(_gFO]A^1aOTQVK7G-2/798(?UNUgN?H/-(==@E]X
>FN.NMR:#<>;,_\(0XL@ELO&c7_[5GN9WV=2^9]5BWC=4@eDb;_c8:#f[TH3WgP2
VY0X/(/#^XO<.JMB/?83Eb8->VVPa>8HT:_CP52dI38F(C.HXH6FNgB<U9\JI]L(
KgO.5MZG,,NPASAR_X?H[b[H&VgBA(.?4O7&S7J8&9K1a<IF_,X26eT^-T&<CO8G
P96MHQ8R+?&G_I&EVO2YG_VVQcUS#B/#eD[cDc=BW3\1<I3N.^=C9(&I.P<YDaeF
8YG.9A0bO:@#a[D6X@V@YOY2c^-PE+gM8B)RgH6S^/JN-E^H?>.<&S=N(,fDJK-^
R-O<c\SE=@0#7]G@YQVa?](6bX0UMgfB1cHZN=-aGRW+Y3b>_GS,&O>WYQ/bS>>,
eC8V29bfDe#G[)&BcVf^_:8Q2T7MV)/RZBP:-K.a.ZVUX7\V@TTbF.a@04;=(eW@
-,0-[0?(H_eH=aROKK:?)G-7gR-SaHdXDgLT>2M)5+4OWAC>J0GM^X6JL0NZ]EE+
9)3??3=G^a-SNVH/W5(UI&Yg0J>6^PSg-gM>[3[;=LEKM;]c;_/aJGWMW\gOC5M5
Te<=9D<Q/9+.c]&S^/eM:GE=cK4XVe]:WPN??@U;cB+,]3M_Z@a4GFbe^\a:<[?-
JVN>,+SN(Ra>T2F&:?YE&3/3VMLIWbgF0@&0N@&9E>UACPTCVMI-R-)M>S0R=Sb^
5<T3?cNEDVT?2X<6=A6[XeQa.CS>591LCV8UZ42##.W^M(PE/CS,W^((.@--_GR=
Q<TRe>3+RWV[=>PNE1E,eUfN#IG?30,\UMJWP^9&(.#>C&P3;6T@IQX1KD],+(]H
\=:BSJZ/cH:\DB@E42S6D(6315/\/I0b3Za><<QS-@U4V7g95c]M6+DT\aD-@>VS
f[FL#=)^cYM+L?T2RM_EOFEcXb/\QXX2C4?IR#5M;Y5c\=:/_=?:<>S,Q;-3+:\2
+:Z=7XFOIXN7WPHJZ40?EOaLfOD02eP+K)VO,AXW-V-?_dNFa#AV85L;B<A^<@17
]KTd48HXP\N.AZ4&;3.7YM210KKa3P-#5]GL=Y#._9(&41<J>.B]baA0a4,C6V+3
W@V_LZNM8ES#/FIN)b9@EZ]#eA;--2A^6[W+<+EF8R<cC#SgJU-[;N&FP#&.&\;+
WG46#A2[@^J[>EbbaE4Gg685B\:[b&4F/NMJVQbK+C@]MTD?M&=@YX\Af]GgI1eS
O7R<;U5I]IAB[]@A2A>-gbK960/KX1GY#^FU.F5_/SC8NfeLQ#1;[D?F(PXGERHP
M#/8cGe2MG2YEcZ;^#F-ZZ?\M+@)8H&)307#9bLe6IN(38Ada3Q#8]g8GW7+:=0_
IV>(bM<9-/T4Q[4M8eVU3V9QC\#E_E&SE@M,3#gAM(LC)JES?WJ+EH4.]7eaQ--U
+ZR(-6e(eTGc^L<8bK_>WffZOc03I\@V/HXB/X(7SBY(+-&YTQ8.47S>\0<dO,)Z
(KJMQKBd0,fX6#&]#;Kbe7:Ke:d_c2+M=65<A,R-<_72Y,2b)f/=.8U.8+#:7YL&
4U=(8[J]Y+^ZaX_[QBX@Y21g:g&/#IX:5YAHc<Tfa[:2-a@FHfF8L54>d<Wd))TC
VHRXc1P@2XX/P2<6(Z]RX6Kd9WX9)\4YJ=(TGCaZVMU_8H_K[K>1+FW9&XMA>=L-
a4N,K]167)QO?gd:T-3PWP)R-B)P6;7_O1AVY&c^<Lb:C,S;@;K</a&<dY,4\WUF
,:ZAO^Y[&^??OQ;d#V49gVY/POTJO,R50BA;\g__3V<-bODS,MN,/D(K+0YgQ62H
-b-=4,.]DY&PYJ<Gb.89B)Je2f7RYBQKN3g?J5][g00+XQ0eS\-Z_03.O3[)(V<O
NXO#;2P(1ZLQKFB,^?gM8P)8<;4?I:ZbM1>XG9?.5<BJB)M&MSK_5a+2F7CS[_<;
Ig\-8L_D;(T7Re,61:82_[8<G7+K#gD,\8c]BX]Y-0+=&RQ&G3ga)e^LdgLIaHKb
f.?0:K7LbT[9cD?>^=D>RFd8[.15QLbOO+:?7dZ5&92W9ISNKTDHBI]Y<\,G,Q;G
B804LfJY6^;W#YNFX28[;<KePH+dPf.@_ba/P^&570:C^<]N-RR^a4[DQ2:a^W,E
^+g]O+AY[-:bgfO.B-(F^RN>JZ3NL59/M2^.^W^96bQ9PHSL2TT.TW_[+bIQ6V=L
\SB=6W3O6^=3,L+68)JCWb1KELIAN3VS:F_GUgO_0ZR>VXK:,a-J[&,AA3<+T#MW
dRAKJDE,AOA/Q@+PFe_,+N@<OUIbC0,5@6Ig166JSB01;A2,[E&#,U/MFGf5?RJe
M3(FVQ=eaR1=^ZQX3D2_EZ^<J;C+UZLF7#GUAFP),==IXBXJ>F_C8G5;&^R=8\T&
c\BK]gD]Y=_[5Pb62NUQcUa>3=D#[RcQcH^7)I[DZD0CUWZ6#bJ105<8Ke[\RJB]
^9YG<[W=K/=8T_Z-T_:E8R?HGNX<VBb8fP\:4+,7+JMaN7F/KZSA4JBAKIGSd#Y3
4Z[/bU#V,?[ET?MDK6QQ[HFg2ad8ZWH277gbH+=Y^I]AWH6>GaO2#]X@cbe<@\aB
,_9<BN<]E,Eb5:ae>U+84:Z_G=7e,L>K_\^=]Qb?;egD4eca+ZA;f?dWFAZOLAP,
0^I;5YLO8(<L-UZN&bJ]eW^3Od^L3CRW0Ff1T[CKcOUa]Hd8\H3f[_DW>7+gOKdM
9O=@a&NB9^-33X6GD6./b<_4S@-JT1.;If]&LGRJ(Eb?DS/=7NO\\#Q;NN@b<;2_
M-TQSL1fQPOU[4d,]G>Y9F?LU&.U4BY,T3G4;1JM8S=a.>>gVVYBC60198VdI++G
WO)4d=f_\+SY377:\A0<#4.IZ]@^>\)/U/YU<9gg0E(I,MGS2@0V9/MXZIE83(F3
UO+3IOAW@<MY2KOV[QKS>WS\KVSP&-VMS@e-aRO7^CME2TOJ6D0e7A1#>)WE(,-Y
<?VF0@c_+P/?(_WDO4KY5OO+K9?Y,6J;/ONY.=P;<LX@G^7YSf15/=IV]1[b_1;f
EJ^:U>BK\?g;CH-;NZW87f,(&4WT?+N836Af<eB?GD734\^ECP(N/aCQ5\VKO91e
TC^TON,<4HLbJ^[U&[V_aXI,(7;TDHAI3+^_M@YZIAH6<75;=7B1G_-NO-aFe<?5
ab87FV&d.TD^?D=T#H03E0Qf6Z]6ZJ9Z4[Y)a6O(eF5;=6]-@87S@Y=,O4&;NbgW
G+;YgG6QZ>YL-.HMBZX3SJ^BQ>,RUD+a8NNQ)e)@C:.T4HVU#R>b@2Q=HBQ5bKd)
A>VYCTW0#V^RO1#;I7g-dA+^?.;?dI==1B,a=?G2CR)IXRNAKW+<4aS<I#dWXI6E
N[XX>2TJa-4KKKIUU;A5S;^#6TSUNVPB=bZXXZgYCY4X1MA-<10--3QOAT(1G+(6
+5F^HN^66fV^T39TVRe2E/>d@\Z@EPE<aHSeYf4gJEXF&E14VL@@/\1L4@5>EgX+
U^1GTAE5OL+Q,KMDKD[P)8>448/CWEH;AOHP#FD]H/IT2,6bF)149:[ADg4H4<Z+
/DgJfC_LLFP#:;Y?,?.)2:+6QgcWWcAg=Ja7cERT\+/UM83M/3g7:W/A+=,(OJO>
LJa_1d#9J+@1\Va>,4I;dBaK\Ca;W.2a&_14\c^2?UbaE&]UHWeZgM?J]FQ9eSKU
VIF#,OgScGK&R00a.Sc28F>.V:DN&PAcZOS0UcF&dBTJ/BA,(;T;6?@/5gFgFO;C
?F1-V=PfV@EXgD6KQ]bCK]FSKBK9:;@[SI?c#OeeU,ZN36IDY&84[eI8g:@f.EL[
GKKaQW)=85EEBYP]a#WCHeUZS3]S1cXU86U?#K>fJ.RK9TH41PBDWHU]+\ff2?W(
ZeZ&><gO:c>T79I1[,G+;7dF;=R[\-Da[-N[+\]_X]:U)Z;PKN3J+>=9Fg=;?fYF
3GB?_X).M<GFdYMfJZD;>Z5d,OR._AF^N(GCg<2Wg3OY8LO#I&=9.;V;-1O5__fB
6+8<<aOH#S-9fRAX#bOP<_(9VA2^:M8CO3X\HPQ8:.TJc-a9ZOC1eWQY0/TD+.KZ
-0ga8.5YNR^ZfaZ=bV5&c?EX5>DAYVPL)6Md5X=@X9g[GDb/?B.MNAM#NU\;MK7K
2H+\_aC8,_e586W^a^Zgd3#<BHSMaF]?\M)0;N2Y@B)P5REQd^?=NO=YRN+.e-cS
EBb55\]Q..1\[B#U64316S1e.T6f:KT11EFIEdFJ(0eSd]e7HBQRJ+1@TY&NA4e&
B(Q;)ad)0GP0/=?;U/()8A#2B&T&4:QJ8)8=QOOcQ[>4IN4VLgARa1KZYV=XKbU]
Yc#^SW:>>K92Y+gBd1gO8D:M&a>df5((Y@84OW:H@bNTfWb_Pd(.Qf_&MI0I[7\,
b(1V&9(f1YY=8QC.(NXO8<e0Ke0RP>7CT8CfG@:6Z3T8+NHfH:,Tg2GcJM4)/2cX
5dOJS)#D\c+>50:a2<.M17BW^N+=?+O.E1N99:geX,;d&c66@Y<;/5,A=YF,&DT.
g_B31fT#OF0ZW0S5D@2?R5_J]QL\?J,0DO82UFYT]MGa=\EF5bbc3gL;-7f0Q(V2
:VcXIU@\3D.f/=B7_]V2<Z)6cTg7=TR1)gf);4ffT#G0S1\9b;2\C&Z+f,RHAHS#
?U(E4G_./6ba\WYQ8X(1)O;+6=?C_[7?&T#_[?.S]agQMZ9,T<UT&PCAG#_ed1,,
2XIRDFS4>6d>KfWL;^NL0U#U7I:D7>ZZc\:15/S0)G=aCR^d6P:OPC?),V@A#LH-
3RSLUMV4(/Vb99\U7H(&\&G2K\#=P&O\SLUd4+AdAfI-^#8\OYe0-5E,3O;Y,?V5
[Y;>7?7L&#e0>a]^I<UB:K\K,F5RBL2NUR3CW;+CS3#S\:6A7-T7A;f__ARQ7<Nb
O(.3N=T1ZPd2?3829R>R_gYRMSV#F,-(Hg]JK5-_]gS4?3QV9QY_2T^V<4:-f8fO
C)Z63B0F?MgBM31X6&LU4EK\R>G.d/K^K/AO2;[[Bf11NKR+49a9R34e3Z/=C<6K
d;M=a<fQZ:JLHZ]ZY3?@N+[42196S,g&Hf/dB4fGeTd,;3PB-)+:d4&T872JB;J;
:T8(>SNE[/+,YI2D0F2U2Q;QfM_3MYCAJ6[:@;M.f/0f-LEMcb4+\6/.=E+=QL^=
56XV9(E[V.S;IV6]]6:0W_eF^FT_bXg\#&ZB^)VS:8J=S.N^NM&[FV?5G[^E+8BK
N[>#_ULe)0-A,ZJ0_aQ^<,Z_eLF_KB?b@&HK-?P5+?&:K-7BE8K[OV2KXC2YKGEM
Be21=3X89/CQB/CG#BR18E<VD\K/^#\UD./<IB+FeJN8XI;&>V>/U.eNH7C&H5_K
9B\3[,fB9T/UP6Q.KW?QK3F7KR@0ccWHA29KN+Cbd?-a8@]]J5M&<CYNdL7NgO47
?M6XUUO_,-d^Y.g@I/.2Vg5g28/R/6U73c2^+/4Q4+&[6_>X?I@#;ceLB7,#S<V6
BL3V+=UQ\^Z)/31#J_eebeW?(JMLVd_0bF9;?4L#18E@>XIC5J9)EDaJ&Wf9R^YW
?f^-C2HOaT1UB_2X9-2JUaWd/@^TeMSS_T&A5D1^BPC?@[7#8dR+YEQQ.bc4[&Q>
Q#^.,[40)PKXO1_]SI0&<2[U4b<<F6dB>0E8@REGNfTgQT6M&;[E,a_<B=<=;VP4
]TGQ1A47TT8R.D23Y/Uc<#Z-Vc^\O4+ZJ1>#DU0UI__2/5N=NM-C2:)7W:,RdgR:
cY\b/b;R&C:^5.Kd2=64>#M&)GFf#>EZ&H\HAX6.-9JV/F(,S579>)]6D8K[VV/S
b(6GKJ7U5YY5I1f?L2#QBbQUTR\E-f>D]DMNKHf31,NN:e-gT&4UD\4QNF1YZ@(e
;PD^1Z=Y:?&Y-3;7[I-?,)CSHBfd^A21bML]E6JDU(T\5ScgVA?TX.O9L&7DJ(M_
&X)66QJF]4C(<,CU.aI;0MY+E<gLXEQ[eQ<L4_;O\-/8(.e@\LfKbL)]5GK#YNBH
J_=\NWQY/4Y69XSGIW/[#OZ-RKO:F.UIAW<P0V,T?R-CYA#,.ge;AP((7NK\Ig#]
-Xe#3ddQ#[0#)T>)<MHff+,M/(Y)G5eQIAEL@ZH?NBYY;)V2SFaWL5WS^T+YI3[7
DD<<AW-G&EgN=8R;XgV,#(e2J-A2E>R9QJ>Na]Z)6.g(FYfa)32gOY6BEWaI6#5F
_d_OCMZ,fSNKbB6aR?Ba,F[GNfA.;5)1Y0\?L9F4U\X^GNSa2OG^7Kc&@e9^,eYX
L;/_FKV+7a;75I1=7;^8LO-]8P>W43P07e?^EX<)E[&0E7GINb4d0305KM8D^4(;
S2\[7#<<c6RK7150QKTR:,ZE3PbOQ5DU&Lg]7&RVK;QBW44M>N#-A\X),+:NcGA.
R,J6NM6N9?O171b>PcMDK]dF)CdS;UA)NC5e^_K3&L-UKQ\_0&52=C&g.CNIY5d4
a;_=Y@+^M+g//;F^Y_IS.FU#:R6T]b7++6-abX+/04[\6\B10+;L=RH,1eBWJ\PD
+_aB=-=#T(^UZVEgL4b;[a8J7QK(.78cB9FEO<,;e@dN@B>(;W5?7fJf-WbQ[f6#
VD.<;YVEFdOWJ2#c)L>BDG1WB;U:>X\6P94R6&9-W0I9J\3SB]@?\R[GTA-Ng(/S
b\ZbW0XRN7L:JY064P9a[YV3Z96JaSUD:-O^@bVIgaN1=M)J?#G/(GIE\7<^?RCI
)HDYQ_1eGZ3RH]>DOa=&[D#BZ/(Q;Q.L+^;0YEX_>b^fQ[aBf3I]ZZeGY/VVKX/Z
:;KB2^DLJL9?;A0IaLC(a\9(;Na46:.O25=YC70FS.<c#8X@4cK3+8_OTZ]0S]B?
1:FVLW(YBa\6\5?3BGN#^-JH6?[MWb,CQ.#TCR#BXM,4872?,F;W2;DDe,84::]<
O-&GOLSXT(<9XeHP<^+?IC?5CFd^IAB1c[K9Q;HVOJPI,#QG56LV;^S>Y(Y067dN
A:85)4U5PeAH]Z4O5acY;19VK<0>KYLf-.#:.RNK]52LS@I:+/OD=b;]M\=#W:U.
2/:70GAX7]&W-DD1Y?VKeV:VPYKW:FP==E;D>[5GQb3fTJ=MS@fZ8DcUdJ1N.3&F
aC:PYWWBTKdP:b9,PbBF(7./:S<cCV,N6(32b=&-LTPMNBM3F14=VVcV6_8JMI<Q
,[IE:\\AZ&&;965g3UZXJ)bZ;<JS<M_c(DE0OYQ-.X05Z5Z5A.?a738c)\Efb5F:
K?=EE(14WRQ(Y4XUY@Vd;f2<CdOQe/]S^1Z<NO<bYUU82+L\AZ34MaPDM+3fE(3>
:4LDF)G;ZD.[()Ed5WP[=_NfI(P_T/g=<KI/Y<N4(6AFV5QN?_B9@\XR8D?Rc]]N
A-IE/D4?X38aAQ7UO9[HGJGe1\3?S.@7c?2;0S5TPFgZ4K=+63SLgMNA=-dZL]@0
#[bTL=[8]#-A9:d_^gVW,ec,\0E6+U#RY&+[)E[SK=IJ+:?gPMAbX6H4&J+>V/(3
0@>K4G7D/e(L#HNY2VX(-7I9O_e8LJZWN(S4Tf6K>T:RaS4OGWd&CCC3(E=9KV6>
Q.ZSW-c25Y#H5Q-A(=egWEeDB6f._7K/=f4W/8S=W3]@(_C^PKH_:(5P2>d26YZS
,O/E9WSOQ9X1U,?W7=0X7N9EA1/;F#f1C3DXZO8:KeI;;MXP,X;V#Pd.fa9Q.ZNX
H7[TZIFfI].g8&W:APDJY.cS0TK2P3KNU0]^Lb/(>cD-&>UO(TLIPDZ9gT]aH\fd
UN_\Fd(ZdaNT/Y;^_XgB#YbJ3bg.WTUI22YF&-=DL(:?0C;]Y]\K+[e=KUO2L&[X
/&5DC@1,PAN(<3;49.,XOef#73SRV8g<Dg;f<XD.(;b8dP#HY0TUM9P(>)7?20@<
=MDXIV0Jd:T_<-_GcCIX6^2bJC@9^N]bA<\AG8T^6VMR_Ec(:Z=J97?Q18#ZHN1A
)TL^1:6K(K2-==^L[H-1IY+)-/MOOE#GZV(4Gbc\A83@EK:7CBUSBXI<:8gUJG17
W;e9IfL;CaHF0)2cNDUI[gbTOfOTdQCe;8\5b=6,D(PXM=KA)eMM=fU#>^W]Q7g>
RI71X&\BDg_5B8X\OLQ5]&6S^J;,6ENRQ<)(fZd9HLe,X@X[+;9[.-M.C443EeBW
//H6KB2fDEAX3Y(OP+cI<a??9-RHIcG4N/RE93MP&-/+I^IF[)?T6d0d;VE8BF-5
MBFePOVH_4)@S9N2CNRFF[CJ26ER&#GZBH[8e+V#Q/F9>bU2B_97?d02Z;U67)N>
IY(<4VEV9Y^cg>BQRB5K5TV4g3N\Ug<aB6a&AaQ[KA4Q)+cLX;c,e#F1>>G#MY?^
cAB_?fSZd6TEUY>^/L0CXEf+[K;@:aDZea#8TC<T>2=&+Pb)EUNO,Z#:dLV7]PA]
QF9\66<J+CS&:ZVOY.;aBZ-K[1;IKR2dcEbe(^>]dNQ.aEGDFH.SEcb]:X\.#RC5
ASIJ24.fVH_O.C:CcLA6Ca[HaMLQ9QT<(J&@KPC&W(fcASECY+\9=Rb85I@KUN@:
#6(YWMA1I_&?;8;0J]@:(&?=\72?^[2aJ@KA=bEb&;KA&#XLTP+=;8UE_+6IZYL/
3&3a55bWd:Rbg9^9MV[U3,]+I],9CFPW,g1UD/Z++bEg=O@3RD?2RQOS#\/]^0#R
<.P=af+^[KYVJdFO7X,1C6Je-L=OG<]T,U<^A:G?Y@U7T:36,#[+4)Qg?XSW?c=Q
UWM\FEMVHH<V2A-59?d,<^X##V:W[EgAa>790R5).ZI:\M(NMVU=HN@T==MdXJ9O
B:Q^a:3=;W+X;(a9CW\.M=c41\D3\(97Y4GKY\XGA48f5dM79A@ce<-74D#PY=GI
5eRC;I-/(+O@+O#A@,(E><c0PdR_YC57E7(fE=+\8JFA=@,\d);GG_7G3JC.1LXB
(&5/(0KE&V&C?+d5Q]D\4W(S(?P/:e?KZDZ]T\>d/NC2,;T<7_S?WIA7+b&,^>0I
\#IN4fZL<C=DH:fb4L>WF55ESd<_d^ZRUZPAe]L.]d(U)\dGW3:f4^\T)&UK&;22
]W;7W7QaPfO<>O(RO+7eWQBA^NWU-g4M>aR4fSFYKBg^/4?2<0FWTLKX.ZU^)CaA
IW(.gN]6E1JNQcER^9LBG>>CVOM2R]9N=:M]a+cWV-PVJ?0TTbHf-d=PC.P/@@RC
4BVVa:,:Z0B^;@Hf+7,-G8a4ONW/NF9K7Me2,W>-.9U8b-H,2UW1;>=N>aK2eJW<
gg^^d0,G]50f+<ba4P29B\G0U)IJOf?2cASYJ,4&.A<U/ETK6\Ad/L-ZO-g)>)7a
AM,Tc8W]QB)5&139].aAZNe(FX.I0D8edCP:3_?3)_;M6(?,^4#T_&[Q?.8:\F@/
F>5KX?\8,@\B3CEGS5UHNJHcg(9B@P,B<5^H?F9\aF#IY;g-8\L\Z-CE7F)^K=IC
]E^0)7T]M&OMR#ZJ]F9O\H1/PaWFL][/58.]:ZU+[//R@9JUW5#QZc51D(QM_V5C
g87JI7a3^\04e+FO\_CY2AD2JA?UYNLJO3IK9_X6^\]K7+=#@dWYBH1<2(^PW_IE
F0E<LdcgR&OGXIeD(bH.)<,PXG2XAG5UMO^afBG@Y#S1K&,>YIP<ZGT=cYB:\TbU
CK4&OCC0?g^SNg+ScVR(g-^-)2N:+1,8dK53ZG(T,c^GBa3.HVGQf[W1\/VH9LWX
,0,e_#3@]d];a(@_[>U^7?6ERYD29QAg(,.d@QMGQ)-@V&1a9,KXJaG5#A>@b4FT
MaU/C2LBf/^&)^)#(E-bb+YIeAbS7B4bSOT;2eP)#TV+g)Y_,PgU8fb>3(#G.00>
S=RVRC]E&X#@=d^8cc8?5<OLO:S/fXS/<+RVE,Ab.M)M41e22(4HG:J2&]4AIO21
QP7IFb_9+gGF<SW]C:-<Z4Y;XV=LVMC,7]&&TCdVI)Qb@Pd8]VT)1,GbO>:3-M[f
8=I>Ec_A2KVT\7,Kc:V(+CWYO&LVQ[DRI<Ad>@I(40,HY2Mf(RGGKRKfa5Zf4N/D
PZJ68@5^[JV/MZ_0,=#EWJ2KcN)b;10DeUgc31]eE<3@EB_^(DA9O&JPdZYF^9)D
\J-ASLDFC(M][Na[#97eV/YHU8Z>@/U6>R7)O_UUcf5d>/<0A.22D?P?[g_5E+HU
d]#G9cOH@@78e_3C=1-I-HM+)G#BcP-DTK0E\/g6gS;EEeS4d[_aS\_O(ZBdMX_E
&M,e?KJVQ#gcGM_Ic^;HPZ-aKCIfH&F=4D:K\d?Xd\c#9e;6EE85TW<6(D#6IJA_
B0PUT>[K]O5>Q<>K&XE;2=5b8\=)&\e?Q-G0(T;OMZU0><+Q&QXGT_-8=B12<CJH
]F;dGeC[Cb^]Ke@GYMGE;U]4,F\bgWfQLbY.+A7(fSf#52b6U5P(HZ;e:AFfGe?<
TScG??5B)1b4:=YBG,&fBZGTcd-<c8cX+_@Ag>S,EK0O9#[[\(45^GXSRe0TP5QE
;P-OWN_3=TgIRP#8aBE^+DY=AF_FV,@W#Ng9K>\2I_C5,c,9I9:V=MK?C:.YJaF@
C0]5ed?e4S(GPQ7[Xa&eBZEe[T0,OB0SaU3:_NK)RH]5QdPe@\,5==8.LaS/FXM-
aSANM#BICVQ#g,bKM?NUAdE;77>]->82[3(SH@J?PKC#\KTEf9(HB<E;O&[A/S\a
5?2\EGYNG4Q&K/QA/YVO_&[e3R[CdTU:;_SJXge2BB&Jc1S)Tg5eD>PX-XH7O5)L
U[JU861Zf<=-KCb9Y,B#-CUBQVAO[V[=04Q.9>9?7U;-M#J9V<+d9__CO4c:[,^#
dZTWbe@JRe>&\Z69]6>3@CH0G/e-g_c#4:a&3G=E1_W8S,c33OEa0_W+UfG+<W,7
#O,V:KC-^B.O7JYeI>]e8&SV::\,PHPaYB1QXPI7fQ)^.U#&,82_HT5H#/ea4Y>I
gVK]:1bFY_V0>Zd1+;B+)+9<TDZ<Y\=IM0O&WGd6BRQ_d:WA(A47FN@=VUc0@:JU
=[(=c2R^Dc:@&,X:0g7fSL[&O(d@Z7MMgB;[g@ITcgYbCJB&W9?UC3DfK^BfA@HU
^]7d/W<F<9RAG/]#6CT8=<Me?X=D#+=gPeKRF9N)M5O2bFTABEO.eG08:F)IeNI#
#9c89NDZT/:Jg@2T3HSUWQ/LbXa?82?YT:\e3:.a7YAWf]TNbPf?1ZKILVf54],S
1O7fP?,-_F#,N8]>:L9_#3ENaDfEd-JacgX\\5FLF.Z^T>)VLCHVMe2\b_bC,SQ[
\g)YI6/[5/fYVfa=,b#6X>[D#dQ1@[P&VcX,5fB1N[7^G1=0Uf1MHUXgA-]Q:?<M
^0P@=If,[Bg_ZB7#^2B1a)8[MFT+<XGaDK1;6F3C0CEQZ:Zf/eVDcM)S8I\A49-c
0^TXH#]I#RI4H6\U[=.R)d5X]cNHRKV-XUV&197,><MJJDCS-XDT+JT=X]GE7Z-Q
U)A0@L_]H.2OM28UW?/HF\C/Y^a4#Fb@FRfe3JZ?c^E+3](5=3YMCd+\Y2bL[+[V
><5#QeN#5;F1Ha?21/B9HCWaab/0W8?]S4QRDQcP,[;SeAbPHbRbD)2gNe#PbG/5
7S=#Z2AE;7E^D^?.@(9XKO]Ce.[[Z2/PK8944A;_7]c3RJg@Yc(M^N+/&]2NXAFe
aPgSS?E?g1)N-1<=U;+1EA)V]cNcFJELQ98Q^)+22/2GKU5TUc9HEXL-XTO?EZZ2
a=VRCWg+3A^#60PgONT2J?g(@9,[,ggY+:1S87C_H0T(eN+a<TZ_LR^@,=G;LHdJ
#If_d_Ba9>L8eUUG0G4=647eVK>8I=^Qe.&38S4dNN4@dXJZC;@A9]\W:(BA>=#b
COSJQ7:\3ML^VWLUMbaD)/NGJU20b2^\L0HX\D^JGaN04db7()dQbQA5?g4SS[4#
R)\VVaS([^(HX8]Tg#YC23<-:FC=ZXYG):=F^DE=3L[.=-:79SZ77?UX+8>7,0K.
P>>7Rd<XR/-KR,XMO@a18FXYG>Fd-C#2;MP0OW3Qc2b9@-aF:>JYTP_^?0C(X53a
#2&]^P8.@;:;G1X?cGcJBUFZ8EYMf;W9]Qc9g[\PKf1TcE0FH3S.;CL14E)C8f>\
)3E@,M@>//HN\<>73C(0:dM2B&DVNJ;BZ.H=ZZ4LH(K^A6N;,^X\VLRfOCJ8G1:5
FU@WJ1J+HWBa-24<3?)Z9.UMBNgNg(M\ffeUKYU,H9,EB+/f+0=9L6<=NZ/(GS9e
2C<5^O[bRM5V6cM3];I(\D@O4#<.APd6TC[H_N-cT6>ZRIMC(8a?E=QX)0DY@fWC
BYYg-D-E+58RT_QX,^#?gH6@YN:+):]+fV3C_><<,=+,MKS((C+&:D9[=X2<1O55
N[6UWGe+]>R-,12][KY.I]d\]NReTNfSL,>D-9Y67bVMVc++1UF6P1A:;^]:@dg_
\65@X2Q5=Z61Y8#V:?0^(cgK)a2>VaG;K-Tb+F>JB/,#,8?=H\3f^8J-/c0GA?QG
2aU<O1eZY<QIeLAgA:c9\OeaTf425KdD=F+OLD)K[cJHaW^J+G<0_#4>4WFbG2c&
),=<cH,bc,]9gEK;4Y?V()cB2E.a<->UF/8;f>@^W4QL5P8,:[9[>\,N]).?HaH]
2<DTUV?BL0ZR8)Y]AU7B8HdTVV;K2TEL@^C1IdCO3Gc2EYDb:#;^>N37Z?EHDE_I
VQD?/@35JC3N_HRe@X/H8K6CG>gX0NPIAU^&][:/cZBRHWON+BJ0\.9_JB-LSDS)
TYP1HV[VXQ-;TG.6MV9(d>N;fQG]P8-YH&)2-M==V<;I:,14YI]Jd7C,N\[\Q&LF
,(5QA49DPeUc&,NN7g(MeFILZ[70<4P.\=NWbLbF;:HAHPHP4(JK[9SI5AI;D+Ue
E&<F\Yg&N+;D\^O/V7=ZS?^WDLITB5-g[GZ1d4X<5DV,a3+.1:acY:T272geA2?T
<YC#@\YW#01:<7/X\1eFeFDOI&,]4eDEHXe@2^d:N#)G-08L6]A,S:f^CVHJ:DQ_
bQ1da,_^AfH/M9#cBc_(NUXUTaNIJX6\)X4@E#._6#,YUQUOIE<9&3[<0(>1AJBV
<\(7.U#3-BXT.OcX[?-2,,,MYHgB+8cM=-I-TN4YT03SW9LJ1+8/g.V&THK/(X@=
Ef(^I1)BQV:=2=-:7_L;ZY3Mc6d(CXSJTA/O,XgJRLY?XG^[E^OZ]S?Q7f?SU]+Z
#bY&ggS-X27SH36H:#9/F]9J+P73JJO^G]_PNZ=aUg<b^9YGGI[8R?IWg#4c/[aR
+:d=TbKCegOVVMJ#+,GP<:9cfgbTc/:\6;Y&7dO>+?)-eIU)H/Gd7dTVRQGE\>A3
0>Z8HII4b?X(e2GL?7b/C1[:\-c-L@UI<g1MBf,2Fb>PSF0/)@ZZ\S\@6>bJSI+0
IND1TA&?)5SU0MHS.P:52a(/7:O).?4AZba+UI)O^PFB^C0(6cS,MI812EM@NWU]
P+^K/(MCVFBdL,5J_B3=0]?O?GZV:GeSWTS(JEH8A.>?cE.fJ[G,OGPNQ_DCL@G9
J/ULJc9PcIOcgBbe#+-DC9=C0WU3W+SM4GQcQZ/6Fc3Z5,,@([2X>SBM7L;GKaX&
ZY)Ce4S6>O0>/E&.;eVNedQ<[g6_@dDHRg.H(c-f<6GW;C=OE,[5G[18:b3CIM#E
?8Ug<2>KQ[QQHdW>5[3HLeM]He4Sc^>dU:0/3Yc?e5XX?g[YK2V\<fX;Lfe52668
I,2]3G9C.-<)(@O>ZS8dXg)g^XQ43WU:JY1FCQ&&;4X3FAf6aLKP#_YG(HN9Z5R&
6AT+#1P#\Z>9c^;#d(AZO0e:Bg2\]bOUT4#U\L<U;9\d#H8=WL#aM:>LAN,?4]/\
H(,LZQg=)<K#):HT8I4?ZVD-ZSN)MEXMa4ELXG3Y9(f/2ea.R26VC2G=4e&Vf8f5
@cJcAYIg3S=f#.#_YHQK/\&5@gMBQP<@[,]eI4;D(bWZ=/LLM[+23P,>OWF(7UMW
WD.Z-^S8(-a_DO1G\^>g<g@31_AXK<55BOBFGG1ZbV210F9M1QM00d?6INX7eBM7
Ed8BPb=IU.)>cbT,5O[W2MPf.GC[90/#R3bWN=G]\NAc91VAfSQR[=f37OD2;UOE
)?Xe\#DG04-,8BfL:Y,L\fY/537-,_O#R^?#2=G>=Y;89I3=?&#DdGK^T9]P_CaF
L_59MdI:LLFCSW@g1P1OC5\9]PbE5=R1K8\;ACT;2^YAS3^e?dG+.e2JK:G,+7cP
[M5XI8MgfX59TZ.068ZH42FU#AYaX_Y6,UB;L404L\OW.4G-]0;ce\U5K-(XJ#a>
K2[;O]_67U;0E+2LEFEU3RH0Z:>;CKUC76UR@1e,<LgFFDYJa\E#IfXT.U(PQeA&
N7HHGPE&4CH9E0dRV#-:aLH50LeCP?a8caN.;,TY)<>#UR-ADL506F-I2(.LJ;D,
66::LZ\IAT-(K0F]8LM#eP)MaaCLfd9VD&M>T9bDH0f\UfE,c0W)>IUcI,L+<6e+
fGV<G/<9];7P81L8YX[.N@dHK/JT;_.TYcIJ(AJB[M(DTa=PU8#0ZNC+@OC4EM\F
^H&CE@gbG:0-)(=Y1-.Q@^Wg?6HS4]G590+:f:=dE7:K+KZ[K6F.f^=49M:;&JNY
5eKd?/cP5Z#C36C7ggP&AOO>P>INV?<2?#XdOD9EDK9dM1gWd>H-<#gEf8^[?R8<
5\IGU]aX=TYJ_/#L3G=B\;4ZP-X51G22]=Q;B]3,-&1SGc.=ZHZI,.W.TT-_-XXJ
?0X=FfM&25NG]#>Z<CP]f9&Q.&R3J^cF=##I:=BP+bdY^0]FM+QIab/XgS31<_Y0
X(G<TbcUa;(C@(W1J-8FD--W).<J1]Y44[VNV2DUK<)AWBQ6&U9.fJ==K<_5IRE7
7Tc1.\bV6e+3ZKKc7cFD70BPda,JQB_.#??ZA.2TZ9eIM:WIgKC=<4.12-^K\^Aa
4IQ56PY<23e+dWIS?9OfG-VgFIad+YS<N5T8cG/Z-Y-G>MMTD3ebMJRK-J?SY:QK
FGd+#D.T:a\Z0f4S[;#D8De3Db^WV?=^C#BF[4KUG[Q)S7YL4BRSH<NOMQYF/UHH
W+^7O&JN<RG(UIN<[YE=?@C5\KCDD@8&Hb>(d),Z8+:IV>X]?];OY[BF+A8\Z</[
R:e&_G(2EIEAKX2bS\5VA,R609HWT6C_P7d8Wd&<;U)M[V)Q=#O=-UQTI](DR1L^
<f\,,6,Cb(/TMUM;QZ:eDg8&?QLLJC^/GIaUQ1H0?SZ<&+Z7[@EK.=?XUNT0e5(d
K;dH79B79d/bTG?VUB?),.0,0[0?@0fRK^6=JT:3;8<61bX\dF37>0Hc^K;D]86G
LIP.GDA]EfQ?,ID+P[5S&)E@KDJR.ARK7)=dW#<>8YZP=?50)R7_=&eL.OS_Z2bC
eY947(C0A:KH\#7SdGMV8e?C1&Lg48Y8bT,9W2Qe2K+Z&E36D60GEKcc.MV-2]7c
QTL5PXK@YcWa9T<Mdeb\Xa8LI:;[6ENYWd&8Dfc<JN3<4UJS,PU<8+PV\_FDO2SU
Q+N=ed1SILQ//cG1<U9Q11S;L<(c,8L6d2^]Y;D+?LC)f[2<)C-?K\4a526_40d<
>[\<CN[6)YHHO0[W6(RL35a[b\-cYX-M7@F+_S)RGN._Za(b/8-6:[b5T5#a_1F)
DfX.TU:R>:#FN[F>Y\H_a4^+Q@E1-3S?PD?XJUK5+gX;DX3UbW^_MXTIEEI00cgK
2/)8;_P>:7+&g?QT=<XaI#=]Tb-<[?f;E7a0DR2-)&SKgT2D:.>GW,^G^?_aCK(S
-/<M<<eBT,Og(=ad>7:.I&&MbLc<T6-gQV/:Ae2\QNeDgf?53H]A@)WRF,GQ&L9=
14^e_2#a0\Z#\@_H/->H;X6^eMO]K-g[O(TgJ]A)DOUd)PK\S#,?KHE#AQ;&fSB_
>KLPf=a?c&\?56H_-=<-1>,e7NH]BT6O&-,GNPJ<@0K<PF>9UMa<86&S;gM1GW<?
Z<,\V./W8KEUW]/RW3>:b:U)K)]>bW->UBO:6K-6FW?G8LDWG/=4(e,,Z\(S/47.
c@7Q,\00SH8N_?2g^-MRP()EK:[-/3;&e?^-+f<CV2R#g;_c.e0:UQW=BbO>ZX7]
[c.+bXRA)[=fJ1a1.ZH&TLM(M+6A645JBaXX-QQGED_4RH)G99\KLR;SQZ53YL3\
?IcbLTg7KgYNU9SY;>(5AH[PS2Y+D2A[DHXe>d>#&N>LJXB4QgfPQCK#<04R4+_a
@O,MA?HM(gVNQJbXY>9Bea1FA=bgF7+f0:[5296MYET.DZ:]GRV[12KD_P]c[PE.
MFbG/&\dJc=\J;8GK\@S[\TaUM-M76LFZTF?eFcI7,-FdDMM0.g]_\;]3c]AOA\:
_^;M77I#ageNDIAe2O6Of#F9W@e.;EAI:P:D(:e(;3^DSO[bB1@#UVKZ46YI7HS:
SML?3)GITJ@HPJ[Cd>aQSRVF^+aJ@BFJCDcX(]^J,UI5/db4eO)JH[O_\?9407-b
WT[P;YXAOZ,)g\F&?KX):5>,bBTU;R-K42+4@=NfN(-\[14ObgN:EYN8Rg8^]4Z3
47fQ:eEf3[DR9D&J8RD\6J[..6Db^G2-8HDLB9;7>3/_5U[f,eO+.R0.HG#VLb((
4X<T_D(4RH&LeJg7^e]HD6/+S3CZ3g.+-fe]#)a=M:HKc)fFGEXC8I.AVbD6GEW,
T#3=eb#O8JNE85Q&#1UPL#PAO<UaGf..a)(#=U@(c[KRRS>F;c:=.^g;),#bR)7/
()#IDg?KJ7BKW<9,L9ZZ7.&RPXEDUg\.0^5KR\.\5+#c(4cV[5)1UJ[8.;R_QTA-
-YZ0M2PG#)#-\d9(0T5-bXS-8P:#b\QXFVKRZ;1ZI6A1TBXW6,,8VL[T/[@2JePJ
?a<2:Yb.MOEH]Nc]P6Fb-TAG@=2=(:ESbGEDc&UI]6YJaNP,9VRd;<a_3+:^Y/6\
=c>\A=M(#E90.ca-T(a&f/.T\J@[IU2SZ,g5eg59@+bA<#E9MWXWITLX>A:<IdK4
dRJD^f72C?/PWW@>ML(@0Q]:#(#9CaDF>C7J1_ObB4Y/#^^#-[G)<a&1_P2I/V95
ea6dZ>24#3//&4S+/&/>,e[c&>.=CQ=2_(6KMe?^G)_X5W+HB?PaB6@IJTca8+JR
aF-JCV5R;>W8SICJ@M\NCcD0bQaH39PX.A(Qe^12+c9>aI&(\caJ/PWU>\),H-4_
#>5S7Ya37T4c0SWF9+]ga@fXXL)NL1;(Be5M;-W=YSPdGSB-W:EcPS,cGBY/WM&]
/]<<Pg=Z+YfFb43BVXA0N]b.D#6JXB\Vg\MZZTAYI^D7US&B7c-VJ65#E2LJ/RMC
@cYLg4f/U\.+YgWVLC45(Z^<XN.:K1S6TbNY1_J4];Ec<8C8TQdQX\.aV&XQJS57
MZE^-HP/g4g_GS-=/\FHT^+F.R/MAJ@fXT9FU]W#MIee@3cR_FNf6U/+,V8B++,:
KYNJ+3UZRWX11.Q[ac]QA\9<OYF](;W7_08,e3f=,MJfR<+a(WH^U,gKUS@:/>PW
DQG((beMF?[MYF-E881aU9HRGY),/0.TA1P9ADf;2F:cD?c@-SRIXT:@5)dT7b]D
+\55+V]dMcQ?QCdV5#DS_FR-R8,S3QS(9SJ8]_eDYCL@,]Y[1Lf9bOOdI32O6\0P
6_+TWPef(NGDf\.=:/E5S2L)1WW&+8S\DG(KJ/fd2W8NRYf]a@T3Td)[C[7M46X_
dL-&;[3R(bOCKE(Q]XWcXATR.W2N?Ib(Y.,CIM61SIaC(/_<\Q368FT1F8b8[>\b
4^JKdX6(f[JGdXAXR]V)XTQ3Q]J]X[G9O^=aP2-V4fSR(^10c.Z]W(?DET2LdS8#
6,#fP.2b8d^HOb^@[,CBQ/1Q-];=O=^9<C:PLYWb4IabK[I-bG6^L06[B7g)0:&H
9&,V.cOUE.<V\BJ1c:1,W-SWYG9@>[)GZN+GR-73WYeZB1bGM57b/c14SCX:Y9QA
Z<E@?4Rd[8_d]-]#eU<MOa=\+J.J2]I+T,,aGQJ;^2/VT&25fE57R;#\^4W-31Q1
W2ZXS[#,e6D6B.YZEaTMNSD^S\[].U6G3)6dR5Y0U(6H2f[B.IRZJ2=d4TI^U;EM
@\\VINPIaSQSNP2g=[P\L(6XPCF@9#<1F,b9]c5&JI[,MM:7BML-1-@dKH8\^2J>
Kb^A/BgcE,>FZ;SA^2/&9>MP/6<M0<;ed2FA)6E(#[aDJ,[MfC62R?<KZ3PMD,Ha
C@[SSBf+Q@abTB/.<E_UYfH885B<>13:,N1J2Q.e@X@bXg[(M?GA3@-G_H7K8KZ-
>gLGY20?VGT]5cE-GGX1BHf=.K@[YYX8?=F;LKT+K1GMF5I@ID3&Fe]9:;6Yba42
;-R(X\4C&#]XYNIV)V4(fC([Ae#dU(,S0&>@W,dd3&T7cDNX@;5KLCE]e9(CA2#@
Lc;23Jb9>1AR6YOOA)Qd&K^<cEODE/?X&Z#>ePN,5+&2B2&1\;M+G(5(]B,^7]fH
[+V:dD[42#T;d]HR]678W?cHb:&G=L8OF,ea]Sg?[HSG]TAY4c6JfI^.RZ-80Za.
GUY]NcNS4SNW;>#2L/SUIXRD3=N)A&>Y<2a-2\7JKSX-U1/=FBcG=HM/<HN<Z=2H
4SUKO<ML[;b&.)#OI>83O:3V02IV_6S67L#V?B?2L/^AJCe0?/8eIFJ1LeFc0@23
G+1I9](#Mb(LAC/L,&D]P^\ZW50VNQE9:<Ac#J@\GDGc9Zd2/4f8T9)(EcPCB_79
aNb];9:K@0+8L4ZXJ4Y5Y]ZII0U_aabU),8J@=4WSeGQe1:=]@T?EU+ZZ1bG[TG[
EC33RSEF4W:Kc&6=V28\ER-b#=7@a0]_?1-JTS..PX+^]ZX-?Q6+g/3AXA&Y3BG]
JU[g\gDeHF?_1LfV+P/^QQ(.=N8N;5gP3/VP8>?#,ea8-7@G43KD4Gg0)^AdJUP?
-7DQI#<M(I+Ya5eYYNIdIVM]<77O<G7O:36PYb7(O)=O(6J4X_(GNcU0d?A/:b4,
7<3-EX:6>G4[RHOIfEfR4S9.5g7c\HMB=]]aQA>d]8@;Mb#9HdQLP@Hbf@LZ,?e?
SG:OEQN6(GfcL[09-+EA9eE,W5GgN>EF(;;ZH^:e&S[T3LG+LgLU,YZcaIRcZa:A
XP(Z8)f:^D72bMcY0]@DUOf.INa/&,eZ/_F]g^f=W5e6,bC)dT&?8A4PKSQ1UKGZ
H7?<WSP\-]O0b+Q4cKTIfDM#9T1e8IT>V]5F/@MKV2\R69UJ&AVX4,6==/V9E=[7
Y^29TV1SCB@<@ULK)BNO8LO;.:=&7_1(=X?b_e-d;NYeCT41Y\(.)b_Ga,(JG7K2
>4.>a:Ed0K7&Md&;SWL,.=Q(+a-GK#][,6ScJ<G^dc:#W5<1)(7e5^&30R8L-GeY
;afD-Z5ECId]?:0SQfTOXSUI94/)eK8=<B4EQ^)L8f;Y#DZ/D=]6K#XT1Z9:_#D6
Z4#eaFLNgQ<V7/GQPIP=Lc;Ta4H6F+R>3GM+.=RI&.?W+KMZe6]Y]#C[L8HLX1A>
PE:DD63-e8b\>X&-Q>))d75<)2\(/9([^-7_7b[5D3]E;0aH7J1?\/:7E6=2_528
e,:C7^f-^4\<1;I=,Beb0UUK4=:,EaJNK_X>6/)T,G)gN2S<(?@DaUJ=GO_BFBNW
22I[>E?9/_<NH=O\1d6T:/57]L.gAT8&gbMS_2\[2W4UQ8/bLIN+##Aaf^<F<dJU
\XEU^6<A<DL<KfQ,XYXXQ^_^Y>+aJ[SgH):]=+>#T3.MEKN&AJ;P\3-Ca^(G33@&
b);M)&C3?S+SIY;?cRXgK@A<F?&XcUW25IaGWKK1a:/D#__AL&4#W5;/(@/YB10+
^,RYc4:aQ(HccTb<O+4]<4E+LHeW0J1/2#A@9Ra3#IdABZ&Z(]bE2ZB(B92BJJJI
+eAW)f]X=0d]9-5a\3FLM7#3TbI>:8XIOGdQI57HM@#ERTC:W1+a>[VMQ^>FG3Q?
6I>HO@?1cYb>?4^.FA+O3ZVP62EfG+c.4,6NI\&]=BT_:b=FI3&W-5VV[-g6XaA0
F_H4>/P9E,TB73T3fCP:OBc+:L-[Q[&c]/BS-]DA9Y142F;XcV#d@HHe>=E\E2:+
fD-D-LD^e4N8/=,/Ce/PI,A8X#SV5IVTZN@_4-0##3@LF/[HXC#7S/8,2SB#fJ2,
VcdI,4YCG^8DV4984H2V)TQM.O5)R&[FY5PfFE+,]M#9BL4YQBO_SB6\+CRW6QIC
C1]]a)KXc3=YR4B,@BA-5fM[^/3#1SV:7eFb@><fNV(b.6J]>:0^JRXVV.OWVVCM
W?OHBT88[?DT:.&d0L.PYPd_6=g@7P)LIbNWA_[W[3PXM)3VX)_G&)gY<==C]CRE
,WcYE/-6H:1A\IfdSU6RQ_7d2]>&WTgQ4;IYR+;]2[HJ26R48WT_A@>@;_<Xa0Nc
(6YZ@b8fOD,R?PX1ZBG0C[R+BI<a\AQ.T[9DLKfGY6I;R8NC1U#>\bH<Y2e1,+T,
0a]_YJST[CU]34@[bdCeU,P0[_(,&)S>ND.I=(;3947Cb)?d;7]c(Y,R?2OdAAA1
KM\(gOc02<AL@J[/GCCY@T+MKYG#?5?+XKT))?G01A0GV(@I5-K:U,;XYg5:W5+(
SdND)EN.Q[(?L=7d_?N\E7:MAS>AUNIOfBE(T#M<;3J25Pe37TTLYMBC?)g\g>GB
<W?,G&bK5.N;]^gb.(HE2;VHJ;F[N?ZJ7I+\^2>W1)RMJ=9ODXL0EVA6#-Yf[X[B
_9^3U=&NYc0cDG-P<cJ._b+WbV_TIY3T?e#(;Sa0HZC=_4Fd1HT(=\XR=V37RXcO
4H9L98+ZPR<.eMDO+894Y&Tbc:b^0,+;H?-gfAFC@0EO5O>][gE_)[\-b2X7MgNB
eMc-&@&(<6#cP5S=>24W:&IQ@6];H,/cg[:PKN9Q.[O)77Sa?C@Wf.,A18D#2O<g
812=+c7\PALY8):T&8:H@O__];Y(Se[D:+8F#f+)d&.,X1Q^#1YH++H:]e?R[b3]
AC]81>EY1O#Zda751GFL?^YZJ=UL(.De>aaC1G\-JC<>5U/Z8:U==1WI4\>G1MQ5
SeS05cdMJUQf2Ig2AQW5RGf\+4,U8N]U7PUdR>G7]c,F?1@fb4Q:KeFZDYN-:E:\
.8[+9;FN@2HbN/2\?=\ZQgEE:LVf0W5:6SA[T];(g]5G73AF)P_DDfUbY\,2/d2Q
/U6;TK&8OI<Q:OMC&LB\,H)UZY=EZ<&1UP?8dM&Fc;Y8@,W;C.GCTUVS+1U#GZd3
+f1<PU\H2ZH9-H&0K+NbE1Q,NNIZC][,G]])@)\:,A03[KL;e3A.7\4Q6Q[<cZ2K
\D\cMSOPE0I1W^f(TTD@&0LYg:1:1TJJAd?Hf=S>>2B&(AVaF)U[GeRY=JgGKT:I
K>=Dec.BE]6AH<D1,fDE/1[<6MPN1=BZX8.+BQV+>;)Be4L8-(:Rg^?YP]@7/Zee
:5\IQKZdD>24J:/TUJ>.R>;/6XHY@AbLM=6NE#PCSSaX@B@&C=WO<L?CGZcD+S,^
/51ES;^1O[<0-].-g37Z\OS)#-a[?&3[<_IBGTc\ERG=Y-#<R+9=S8,c,=d4gR@4
U&Q;(PK^^QE(+0@--81-GA9ET4c^R3?HJd[8a#M),dMRN]K&b5>d&.cT[>V9bW<6
1.fK&/?Hd:1,#T<CSJUPZ<5DF81(&D:fM7-(UgP4EOg4N&XVUDKE?.8JX/ZeO9>G
_FLgYK3cgET9QE4(97_)6SO/a(@c\F#OZQA>+[7-E)W62A)OfRETd<]0T2\]3a/]
3#Q:6Q&[N.A:<X5Kc6aB:Q/28;2)BL[^L?]+XTJH,7UW>R6\ea,<OMDWa#^6?[D)
QHQBE3?H&_P68_;)HfK8f7b<R2;2HLP8Hf5.gMMPFbF/^]?7K7@HdY4A\\FX>KFc
+AR/CK9<,cRM,D73U2a+V4gK0Oa-Xf/9^K7dZS;TfMM?P3+NMJ.GBI.ZeK9ZaWg5
F^>@62RQNI._0\(GNG4(b6ADZQa\TYDP[.2,PB@T9ECZ0]>CSdPA<,9P<VR>eDEB
:9JU2><Z2c0bOTXa,BP3;+:_TB\:X748PSREK4O\BMP6_UGJ8RS[1VBJ.,Q/gR3(
c+gS/N?BL-eL@cASF#YZVF+__VSC.&M-#dWKb,\HIfH>e:^FbL)=-6A<-OX^2+9J
/)20A+=dJE.7T/)9-3).aCRBV+W9+^9Y4])9bB/1TL4GUZVKH=Q>b\DUg_PWOY8Q
T1)[?<Q\N][]X#:;D)Z58R+HE>[K(M-2e<3(d]R-YMST>#6=V,<FSGZ0XIY>9.K_
SBV=XTYTS;YISa0f>#R/D7?AaN2V@@7I-g[fH#V5XS.>L,Xa/-P::X;cI;DYd82I
R,#@8D/B8]0A0?^C.HMB,EN/3\V<F(^Wf?3OY_E_P@.g3[M>YXLZfW;FF9aTE)b>
NBeB)]H)G;#58+-RLR;6XC8[7aURCCJ0CG(0I=RV-MS=.OH3J]?@>A&\>T29Tg;f
9E?#LC\8K][&;=4.-7)-TSHE;=ACF088fW7XIRCb3C#[ccd6_](-NTb9?1IV.CL6
[A\L<eZUWOa/U4FN.:R7aFCNG^DT7872AD.9SB<e0eZM1VIB(EC+-E].#B\UF]=U
=#;aLb)Q?XYe04/#DZ9Y^/U&JC.&3RI&]7_XJTMJ+>&]<[S;0F)/egM3T(999,Oe
+Kf-HZE)d4VbD4BDZA<)O4De/U/Y#-AcC]DI52;&R/:<./TERU#2#T+,AI^]8(gW
,54#:aS3JKE4CPB1eWAdf<HR;G<ZH+dH75//Y7[<_TQUS01M,M[=Ga4Ag[UHdB5f
Y\47<SUf@^fL1+[c21C/aD[CK>DTS9H^5A@a99]KR^W472R.<<(?FY1JLJSPG^Y-
KaLb-WXX^VNIXb=.DG=aVaR0T8?H/?+\?:R2?O3Q&^<:NAAW8A&1](RQ@7#_LX8T
&VX5FggSX<\D+c92X05G3.)C_?DZd6-QPNW&g+;K6U8Kf<LKAD6;a(1JXG2bJE^+
>TAN;]1+MMW\TH1_U+\Ne\ZU((0O@>/OI<:#TFd?KG2A2\DH_:VT-)+H@K&3LYeZ
(XPM=HC;_^4.,OTR]206_62.RE#],+D)X68dDg7H:.7[b[THdHe;5>9EROO:8D&N
WJTTHW78#JJc;PB>>YfJ=3Df+<&fbfdILeIS0NIg(D]\@>AL\IEFQ2MM]TQ=,1e4
-\)L7HO>M;7BH^WFE)VUM_EfBOE1KP1^>YY#,539CIE1[^Z[8^1,g;fI9XNM+6MQ
],?&?\8)=Lg[9bERRE3>G/S461g(;CIL9Z/X)(gADE0DHWg\Ef.]X;UHK#GdfE:P
P:-;^-63&IVO:8+.S)Ue?R+KQBa\RK_c-:]G<WgUc?5?^Tf\4-APEDGdU9M?5T5M
I)H9NYQ^V[,)GfTO_AdU^O1K[;JcGHA5^]=g9<2DRWZ/DWg0JR_S^/<cYHGe3&Q#
A/WR=18E3<NI#Q[19Z]3bSW>/7[S<845bNR\V6g1<T.;^D-OcdeHWJdE+=^Qc+1M
F=O[ZHOXW<XE-IS<K.fOF=0=AKJT\a+S>;,/AWLIA8De?U\5.;-1Ob(&PH&6BLOI
e;:VT@ST(Q6J#L^UBIE&3Ed-HKBf6;GW8H1(R4U=5a)WI9:QO0/1L^]F6(.)0eX5
U<30\fP0_-:/Z3D=^[2+LaPO8AMU6F7W0JTK3#M]8S3FaJ41IbGd3SR5[93dJ-AK
L\g>RIcM]Y)C+ID)PC?FC&:fK3NDF3AXBdVS,>/.+^-Y/?P6EaC,-9D28A&\6Q4C
CJAAf4[CQ@^;G6#5(4]\bEBR97D3.;=6RH46+8[](:S3<M>;KT0I_V\BYN2c/_V)
O:?[e]IZK5V3<BA6_FXO2I<Z\g1CCf2W\&O=+UbKSgKDUB8:;KH<5MFX.e<&bI78
f+C4^a5()a1SBH4Jg2[F=_CKbf9LcA@+79+2b?K.c5A2@<@c2>R8c.4C?,Y]J[6U
3LAEI>?CQ#:N37C9G1a@WGEfR=18,Be./^Y,C0eEJ\fE.@eXf;8:FI0FCC;Ae&EI
S6#H<dP6#a28?D0\IT^TTZY;F)aCXgOKFOMd^1g_<1X-e0U+NYH.C6..37eW74f;
E610fIX7_30f\MK>Ja+DHdBJfY&<K.4Cf@NW]P/LD]6^LT0eX:JdB3LULT?]_A#Q
CT]dA;B.D:5b/#W34X/7B)N0\@F(U/Jcf:&67F_g@0Q^0H\bg8IRX;?&=8Hf#TES
fKJ._bCED2A_:5^NBX/e;4dC5PbEOB4#59)YC>b;JGIT+IM9dg0VK#U)VQ<)be3?
.Ng451cCUY=:)+>2-\W3I^K5_>W#6g8^1C9D/aFML[W:DR>Q5:#E+=]d<=]:YSW3
BF?43X?cG(#&5@25:#&,Oe=BKBNXP1<@OWPeeN#2FSbeVgYA)?ISNbg\687H/8Z>
cLO=?D2,W[<a0>C:=\<PX4M[=7b\AcROI83\(J]O0^F,]5]UV[F_<@\M&QQ]XZP9
&HSSFS#K24Z7d7B2dT43DLI&?(O^7+\fH<62]K\\V&9-@B4.gRI?)OYaVX-c3RJD
88;Z&4Cb/+2T#G\Z5&1&>cKg68SJOZB:S^bPb<>d_[K96f;A/fdD[gC8>4WCG(V?
?b3;c?](.c1];K3@O_.-=88>>C1D\B@QebH0,9]O#WQ/:.H6-RUdDE,IKL4@Z;\8
8>ES>UK@_,K#=@KGU/SDL+70e(.)=(0f\/e@1@2J\_ROG]EdNX(-Mcf6=X:P:.VG
P2Cc[ACCE)_Q=(KE0X^[G(EbOfE@5H];I#H<WSBbLcDI;5#YX;SfUWFTY\-CS(#-
bH<VdPS72d:NZKE2JBTaU((O(\;>cBc8H@e7YfNc0;dZ]dN?[C0\WLaH7>R&DOC4
[SX&A\9JgG6C#gH-3:+)PK/DTX3LZ,I,8D;E\eNIg13\J6>E,61Ne_(WRG;VMC[R
>da_BRB/\cUXTFfANDfT07NQFd91ZRHBe=#92MFGcVZ(.94+aX[NfU=b#=.8REJH
0G#]0>^E7Z\.23Z83G>8-Z7ER0@G#KQB4:FeIbg5=[Ega#-]UU55\>TG[:H>Qd,5
dXa?>TA;JX2?@O#:g=G5dc6M7bS0g,O:(6I\.UO-I&d;5-GScO@XKSBDCOb;0J4.
4KQ2CJ^1,D(5IHaF3\#>cbTB:?:JT0:F]MJQT\>9()OfL;0M\-ZCY@ABN.CG59d>
U_S3-[_SfFMgc,g6,&+M3@XA/fIOSg:-&N92AVX1,7D&N]/>D@/Z>X^X&[>eS6]]
PIZd+^_)3.a.KV[gCRM]U:9<-@,;3AcC=Z?:eZP=J#&\_4MBcE9Ng.2eF#cZc.\8
b45g_:G=bI[TL-Ug=65+6\ON2LN07&9HTSa]DNBVa0^W[#KH\10BWV5ZXO6^eg..
K6W=2<__29C.dGRNF1A<6G<##OG6D67;&g<I?4_-U4+20QTF<&fV#JK5ecN06ZZ&
[b1KE4>:YN#DR;-d?b&[USCUb0_b,L.)XE#R5S)&:+K-]TMG;SdA1R)+]A2900=Z
8S-.N2XM-CM3Q]0FeORY6<&g+-FgY:0a.+feA9UB++Vb:Og\HI(S7#b+IP[=CZ)d
/8QUSG/(QC<LV-[a,b+R\U\I0K_=6\LYdaERVN4G#DdI=CUY)cO<cY-\9^@/Bd/U
#^(?N=1P\2M;TUa1E?DTL>^KEX#1)]cPEc#^@eS4]>VV6GS-K=^[-U2^]a_2K:OI
C#bcMB7Kfg^C8<KWN8;>cR#f]S@E@7H,:A/-&#DcXc/SBH8&(B8:=F0VU[VU6[G@
]dD8K:[18VdXWcPV9c1(8[C42?F0PN@VRd/XGa^a>ABI;IPO5&H>A,4<T8GVWXC7
K&f.SSB:?;@D9\5<K/b/f:=MH_NS&Q/@PW7N+D9;ZHS1)c16D@AE=X[49FU?]BF.
AWF\#8NL)V668H?=-fG]]a@cU#D776Kf?<3VS0-;PY]4L9e61cMeH2CE:5QQ+;Z;
=]/RZS;M080MB;3]3EXGc]>.CD5YN=1cAC2]K\[6^X=;[#H5bSR:>GUR3;M(+I,H
IF4@bK?=G=eX87fQH:aP6<g)73]^4<(0#65ZR1;:5P9\7^Cc92ScQ=,1NLT7>f1e
M4_F)@&>7U5PQ>_0eC3cD)#^7;V2>dM+aLSF&^WS7\TS@\88L[A;;QO,cQ4YRYcX
&-R4)5MdI<TT]K.@6P0H5f.MB2;ME:T:NMU+fH.61J&I_]^Xg00Y.77M:S/+^a2S
VB,gO3X]U8f-eNcD+[JK916,@<+OBU1UZ(=.D5Vg3_,@@KA4Q?>UR<@f@2A8_LK#
RLSTD;/RN9[V+g##EM/Rd_N^K/>Y:Q393=KT1XK&T3c##K\TXT(+eW=K4E\9Z&#\
1LK/Z/4&S)a=].W&g]N:<Me.CJ>2]c]MH/bJ6B#C).WV11?1AD)g-fM@8P18Q,4<
EX4Z@ZWV]_5SLXD<B?_2GQ@TSK@E5eSFBd>RG<-P^J;U57]0S8E5QLH1JCR:7Jb.
7+/\@0ZOFAE+0Y^f_b2.7\811)D33<YS5(\RX2B&AYGEI@3f;DXO#]8KF+J;#b)[
fA#]5A=X#/]#<X_dN(ZcJFYVO4e,Z>^8+J=A1MW&Ua:C@fbgYKe,(\P3>AK+NK[S
?(0dGV6R=._DFe;C&RLbV&f\g@d#ZT;D>;:Mg<7]LR?>F^8,feUC7cgV><(>2RFe
(S3IKa#)+4>5-WCG9^fN]SIIf3.[@H\O>U./,7D)[HY9@eK,[JK^1@c?XH]7GfAN
ed_OWgY&<-LB+g7,cLKL]RMa=:<<gX6AQ2@LFJ16,0@;F^ZRIF]N_)F;\dE_0T7d
2];9>_V.:\+Tc\N3c>GUcP)D5[/cd(WTUNX1U50Lg,FI\P.-T=UCBab^c[FW-E3+
YD]^MZIL6bL[H]AJgMIP0,PaaUYFF7-GV#OEMa:>XTfL[@_KLJ+Q2UbcURH5bQJ0
AX[^DJ3@AcL,0GR57J0W:?CB=b\>eR[G#\4fO<65P&eNP+_7&)P/L#H=]?B##IX\
)=QH[Xg#IQIY8?b^fB6A@@<\de7=0.Z,MPHd;[_B&4=E^c5=KOTGN=cLCf[f7(3;
0W@6;G]XC;=?>(1#aYbON[HQbZ#070cG[F3PPS(@Og80=N?X3UB>eWERQNcPfZ?K
d[gVP^OJ[Zc;GDO04BdD6W<+0?NdUPWgV0S1]CH_8ZgWN&@fOg#0V/X3ObJ1e[Q:
YZ5_ag:<Z\ea4(]Oe_(&_4LPZ@\A2\C9+[b:Fe&L/,\EVRbOb.Z:2OEOaZ4Mg^BB
5b&6=ZS659>Y^;LV)<bM@KIJ&8GI@JKNegB20O8P)?d#)8EO,95QA=_<+QSBVG@<
K@@#AZV[RJ(=<;cO::JSV-aO@c\LWR@]T#b3aG0RP8W8^><)&Mg0<(,#QQ\.S?8T
d(#BPUBZ?,GBC)72e)9]Y]<-;MDcWES=?FSV#@6]&HdXF+7^?YXDS_&\H#aW1[b/
//MB@LdJQPKAM,101+V;f?V5Qd8dQ<.)^9ZebfP^3,g/76RLL@bKeI+eY.14YBcE
6H?;R]Wd88OG7T-A/bL#6#:Ua:@[O64W0]LABa>/6#a:efQg4K>_^beUe]Ff/2d[
;,e@5eZYGWd>c3=7UL5DHMJUeg\\@._.^Tg_a?DQcUHN8dTgX-##[fKRP0?LLW8Q
?Z\X<P(1Ke6VG=^1#VT\7(FbXAX3AGQdK,RZOfZN<U?W8-e]Y07:3...JeE/_f<X
XF.N,5eb[#,130&&/70DEC88\9/e;9dPdPZ(5NPeT#:,=3J[(OBf2X+TK(:/T=dK
^@8/K0)[XDbJKe08eMY9?<-^X<eI#TQFKF.+?T(Q42:gd2-5b(W]H==J,=c\If(4
?&RN)FX#69K2Zde]e-Hg<IZQ,51/-VW&bH(NI0\2YSeFF.;:B)cOO)af@aPFDa^U
8]X?Z^_Y3KLPbG/=b@)2TK_3O&Z6dJb2P(_7\LYL7_Q4A3[W5]R&C43C1<dL)@ZF
==d1XW[P;a.WFd>.Bde2B\WA+A&&PS>79e3D7.:EP#;CL2/2B#:D-@bYSYW7FME[
61-D1aAY28c=J)NU4ID#9S0LYQIAa6^_WFbg-CT)U2#P-7?g6eKZ:<0AGN>REEBN
DB2J:8.JEDG1SeG@;cX<VSW5NXOIIT\0F50NWUge,V0e;gI\3UDQEKdHE:F^,3?/
M)\.60@V)&W=\&09>H;5:@Ib6X?0;\(@5efGF(0YF+UH&(EaMM>MSB_:FV:KEQ^8
O]Re<N>gOH;dF1GW05Nf@#gE,8eUA=dH)2I<4Ad<+[X.3N^UW.2dgVMFSQHW?0NY
O]H<D]M0+.TeWR[>N?0B)2F,a4YN66IY+Z0<JAMZ\:bWH+d&;f,<B#DGJb#KE3;a
],<>D8K6]U+-/D,\E?[4K:2g2Bb/<;FNT<aC@Gg04RN9VQ+1NAE3PIX+#V@SHJ^F
YKaN:BT8=:&GMA,4<YLbH@WX+Q+;4N#,bG#-EJE5=:^7b8S<J2.(?Y=?c@T]AfEF
^BX2RD]91FI,;Bd9Y),_>30PDH1J_^1eEC<ZT:GUR8+KE<,2Q4TadUV6eT[^VW#J
BF1#V?_-;D[(J#<J-KOJXgNC_.&?a7RBX7=e:Wg#Y5?GARNA92::J>P[7XQB@.a+
/[ZGQR&^F5)e\R_8VX^_4O]AR;0#U&J,KSD2<1]g^b,Y_F\HL7K3UBX#G(KNXDJR
AH@[_(R&&KadHY8ad61?d2L9B?=8J8gMZ4b#)AB,I99JQ,]B3#B0?V2E+fA6XJ[8
9]N+Z4@TB-52H39PJ@A.[ZB)TW[;aY?f34V(e1S4fF/(fC^VL?A(08PM;Mb]N,LE
bd]TA.#?D3CPO9ab@+\Z-3FacR=R\O1YFJ,6Pd/>cAX#^gJ5&4(<\:cJPC;/V]#,
A6]Vg9CJE4Vb?5R;0BZFdQ/PU58,R=WEI#eY]DN]?9TT].R/&9J/?;@?5_L4EHBZ
V)WM7?1K@:3(>BfW<@\>Jf26;b8D=N_<+65#H>\/#.YXP)\+UX5+E?3+WdR-Y,>Z
^XUQ-GX]R>29f2TdJSc(F.WWBLFb9g8?NgH4-_EHDTXID7(F5URSB)V>;\^?855]
63MXOQ3dDS&@=8PO(UXX&=#VP=#=^F2VNFGP&S]K0df8<<Y.@O)afTBdIW=JJ\K[
U/11\RUEX;>U5R1JF\Z/]bAf\(=-\f(_<]1BC#C2R8<S\QW^+D6Z,L_T6;W?ZJa+
F8:\TAVP-MG&;>efT]5AB(5[^,U=P=P-@::JWC_b?0)8fMaG<GF_M+U8X#+-)E0>
^O&7BKW5PC]:=.1/JZeM0CUKSADEWG8O0ZKcGX+OZ620-O50?@T^D199(06A[@<e
5KbL9J^CEAdLVM59MQ:20,Zbc2@9<eAOXIH\&_4^OgaUf24ce\ON;RGe3<@P&d+,
08?Cc6b+JH^>dT_#?ZAXf&?&#Q1R7MRafbV</5D+,^J9=/QUAZRE34,L=0L/#+0e
Pg+-N.W6Jf;NBY\]-^,d;E]/<=748YFB.\G@M@L,_R4^Bf,VO]OZ.cGbJ;&G+;@>
N]1Mb2a\(XKZW-PMd2HQE.SPM\KK)LHSKd9H=2I5DP0GBeNK59R(14.F&3F=IHgH
=(Q/g4c5@7^FRSNI2#ZQZF#4dR3bObFgeGND]>cAB&J6?AJ@,:A=3;aTFCJ#SJGf
@W)L.N#2Q?0X6<6/#I=cO=:f9eGQW;2]R/cbJO;dW]>bH=QCL@?#H0d\?N(L+g0N
H](M.@;cPb>DeBg7@88ET<G#GYJBgaRC)8<V/8S3G2G5L)A)1)O[N5b8CRL,.CP>
)D3JX2A=CEIZ5KPBaMH[,bAF=)E\]SK782SX93A2aB_]\AETF,gA19BO[c)A^XHF
(Wd)WXX/4\SdZ3IQ5Z0e-O.f(SQA1>I5-ASc)5QeGF^27W1,GE4R\#fV?c>_IB\I
Y:e04^dX5+CJ[CZ@6cLC..4O)d0P.5JBe[eg7,3L6Q8R8Z(/\6(;UD4@=EW<,R/E
LP78\#g)]GPL;EMN_JA&CR4,)M<9]>CW<1X0VDeHN_,P<C<P5.&H4V8NQ)0FJ^^6
8NW/\0H#Ra1Z70/>QM]IfR/1V;ITUJaD?YA4a#bRX:4J.4=52@5Q>c?IU-e1>?UX
C:c8RQL>+J^-V+-+Jf<KRZ.?@A5?Q1J/O0Sccee\RU64Z0b>M+^X(NXILX[&=7dE
BTbL<0?MJ8)FbK2YNY34>T,0&S6/Xg33LT_\;34e_.G0=(g9(aO,P&4=AIZfT[KB
3Hb&.OK?.(A^fADbbB4-BO#48.V+U+\\^g7(PI]9@<>/@TdM)083;S59f_M=gX_I
.GWgTUQZI6_UP.\gEdP;(YHE#7dI58bH@\7)e5B@BHR&EW+U8V2b#c/A=E>3d^:?
Pe[MdI,Y,a/4B\4KNbQA+N>64TZdCf<#[b\/>g8b=f-QLV)JA0;I3Y9/DI.e2O([
,AdVMA_d(X[5>_2DY6?d-UO=bSK8SY6?^R45BFB7]0D)fc+<J@a2CILLC)e?CJ<<
JS(JDQ7LWfg1(Q8@,JI=\NdHe04-(D(>bEg(-8X5aIeY2HWI:[\,,HI/FE>>_Z7+
?B7HODa3W^]6[P]W-X/S^_MKM#>Z(RK[8,IJ6]J:IO0=?]GI.?Q2T/f[T2M>c0JC
X;+NUR/G0VDK11W#T)+_D#:QeH]:#Zd_\Rc5G^X1RGPc4Y0c]>#c1]cP:f3eF[0-
Kc/S.E,GC&1L9X[^7S&,)(WeH#_<OL34ED;LVAS?L0/2aZfU4O7DB+,]M\;,+=@/
bHZ)G&-:L5E.K;6?M=^e>aG-dC??^b0T@4.LO<fYLA@_9UHO857)CQ\bXdR6Mf0#
e.O]Zdg1@YBTd8#0U/,UQd_WJ<L#:Y]QLe?E_eF2/(1#V2&@A3caegJ,+Qf&1?7P
-SF,B2dB)A6_3,dg_Z2WY/G]L5[[C.JcN<5C.G#J0_)X_A\H9SPd9M6ARD,W._D_
ae5X56MW/#@\:FWc5(:]#<YSd05Y@d4I=2g.XBHUIMLLC@#2)0(@R8?\FS;53SX)
V5@V88D(@U70?eRFNBEV\>L8M4ab;]+Q/KeaG:De:I1>H?K>S@&0XI3>8/dG9K71
BV^W_<RY&O>RH0e5JgTF8ZD24H0D^G4g:]HRH/);8.Z;Q^7MH3-BMTB:1C<bFA(U
D,eM#P_1YRgc70NgJWfIgdKH(YP9WT6?SSAG>f;>3]1>]N1MHN#b828[g5W^H</9
.W;@GXQ4b_[23;,K[[).BD(-GRI#+QL>T5ADH_;(Jb#E8)(eRQgfX=/c/K0RdNDM
gBO&f+:fgScdPR_=R]GM2\&,ZN9?N\O?bbaOKOV]H=JI),c_@WS4P7OX8(QB,&R9
))@:0RK7?-O&V_,XN>JOR/dPF,UD\<c=ZC:,;V/-N=adcf1U.OBDTK+BI>NAeUOO
aN\G+\\OX8Tc--5f8fbGX(<&VW4(U[Y3JeB;_,V.9P@a93WEF,S?d@+a]Y9)Y_#?
>RAH=9_.F51VECKT6ff1fZEa17;.41R+c9,:De\[##?)\cQT.f?Pd^SZa5dEMRc/
PHc-P/dR=MRf.eCc/63UKASL6#.K?==>Tgdb02S=604cHRS-&7I^;)M9DU/[\-,W
):]0_H&c90PUaO:f,##4bP:b_M##5EIW9.VP\NYC\a>RFO=K@1M-^NVAL^ALB.VB
13]IDTBaZ58[5EX+Y1;HF8F2-)U2>N<f-_/UcNG3?1(0WV8>NI-\9ZK05#6Kb5MA
QG2<2FTGD5IY=VN_@/&HdY5/9eY_b]\<a8Q221d6DO,UC<^RJ<\SHB\GF85Pb^JP
F.gJfCUe5?D&C0a_YF-68U@_V]S3FCJB42JE82eRHf6,FKXJ1-WNA85+/29ZN?2M
4KF89g_SI>\6J]H3MLC@E,#[O>&\=\VGK?FLWY.CVLPP\cXa4Y?\6&Yg8N@a0E59
RLe][T,\UeZ1\D\(@R-_AK)+MF66(7//OL4,-M=U_UH2OFK2-7fB3PS/XY^,YPKM
JegJA[+c\Z:9;2:[XK[Z@8^1Y#U&-Y4I#R#/Q#b#B5]S-gM\4TTCAS959B0/8La_
/UDfU^.Z^CO?BR9eggEJeA.8B6YW2L>EM0aeHa[+U4]M2=.\GMa#8COXCP:2A&,J
9]3NOfC8b(7Qf@@6I1>e71#I^8[e5U>b89g9<-4UTG4,:HF2@EO3>19bW#W.c&/G
fA/UZf-]Nd\3Se<<ZOF?AO;A>1K\=Id<K_[KI-VQAD44OLF]8;W9-HG(2]=5#C_M
CA-6VfH]CU#P(E(HMIVZ>U3@R-62G[80.D95,LE45RgaYZR=_a]\FQXGNd+7XbYK
9WI8MEM[CDc6?;c?:[IdBTAR5B00Xf-;YR>0CEaFMMLF:#Sf>JQ<=E-@1>0.S2(@
[a[]D:BWO)]<K8SGBQ>?PXHR<gQeT=_2aG=B4]K(_7>,B>H^GN/X.8F/D_b+\2M)
UbUXMZ7_TQF@7g3(f#_-EH)7R#2HV3ffgY.KA[/>c.SF1^Z+VKTEAcD8c@8(Y5Jf
.==.,+9<XAWPL<Ca1T>Ce>QYLXER\gR3A&a&4F?HDU-1+[PbYfL=c2VL5.c;JP?(
ed]KKg\[U+,+KD,D=?LE56Q0RU;SW:1&dW-RdbWcO)RdT+(1g;KJ@4a3J>e+N37\
TYGD&[_GOAEZ(<g-4O8R2MK>IN_>Va8C:>TEW3[T[f&+6QWCY#BB,NH3:7[.b^@?
WS_e=eZIHJa?<BX6F]b[.TMNHQ,g5IN?527UWK]I.R\8dgCMH99Fg,U?d&HR>7+g
f^<?=\BO1bT4G>7KKA+gC]2G@X6Sfe9PF5d8WJBDV.V1G/NYN+)KH(DY:a;5MRWK
^?O8KULTKL3KDf\&Ye@.TX1TQY@?fT6B,g8<[+]=2+X4\RUN19<3bOC>6=2J6dG.
?Cd34GU5gY1V?6J68g?R_YbJE@W^HCN<8/LgL7&3;Q6Mf3.)=bdN7:#?Q>=F+a?:
0EU)UD1?Y6(F=R6].HY7JI];+\^:I8.X.Y&?((3H\UAU>3D5;:F/D[=@L2Ja]N>V
L^_eA(@MK&[U[=?0@->U.N&;>-HM/5:.GL;DGKP#6b,7LZJgcO&V>#5?&@DMN9?:
9fP3))L1796.4)86L8@bARA0[VUVN7,DX-5;;:&70T18A:dYK>L7#Cf.<NX+B2fC
_g5^3;3LT(+3[+]6Vd+IHS(-d(G>IQ-\-A]@eD#MQ3OYF_]OM?+EgC[DYI7&-=W2
;)W1:1/8Z:,?3c&PS]HE0bgA[#]\Y@GKK)5PXRR@]IZVUf+#S0#V4a:SS_S;YE\&
MR.8P0SUSY:EL\c#gIbMV?<Oa</_-;/?=XDD;[T8(S7<DN_dYaU?_UGC1gPJ-<9-
6=2J(&)Z94a#d##+>6<FffX@;J1-g0&H50g6:K\=_C]#dKga<4G>?5=4EI2Wg#9&
DT0WV1Oc]#ce0OI>SZ6,_@-f.ffQcTDDa/512N4?0b,EbA_B<[.\X)\(0#MO7_#E
.64XDdNSgIWd22RR-bL=.5I2<^VB#JX<>+>H=D.X>-C[&M6?[]DRg3UW7fU_7^D_
9@L]1;(Ye3EF+I7,(_]27G3YR?R9V5,aSObA\^X_J/>H6NWJ-I5];9d:GgR]:2,;
fTa8U-?60Q53Q4,^]9<bD(EOfAd[5-[6:N4E933>>&ULg<UY7O-/&HJA8@a:]-Z(
2A;HRV1EG\6-0I)Z<__FId@?3YFP>8bXXgBf\]MZfeNR.d@_NE]D4\1OgIS#eQec
)S0)5O.&?C[^-DaJ7GQ4?6NI;X>.&L46RDc8bD&BHJQeNB^,6S&BH-fCcOVA=7>6
EbE-c1)(S1&9HHN_f?W&+JcJ8=4f21Q)aPRL=@PX@abD#-QcfHgZ4)1+Vf6.aV<#
Zf1(Q[\[B@Z\9<FELR6LA1?YYV#PVXYFYR(N_gNc5ZGBN#2_fC>9,+/I^E</OD6a
B8d=\[ZRdKZ?d?Zc0Z(bF>[KaUQ&.XLXLaA;&N[-Z5=[&1AJYH</7)8GC_2<J\B1
<#AaZVRc(4:Y3/]T=6)(LYAXcd\>.QIbT#)P>PG7G.c=#74dNKS>(aS/AR)ggH8;
#2O[S38S9>H4NP9,RRGY9YP=TCL?\b;B2)1MM=I#1Qd]H&Q^a?6S8e/ZdYQS/H0g
JN7g@6I/:^9&1Y(SJ2@)--VW[QMNb17F?e;3gb:/JcbffaBTVBO[L95#(67<A+U/
?.&V<@cC[cJ@V/.0&_<ddG7^=+I=OYRRWA/QNC1Z]da&A9;FC.N+[^1>()e8_^a=
#M(IA;e0KcZ,:91Da@N/ZXC3TEZGEBV/T;S/G<)ZD<]I5I6ZAR2DRTW>.W82H,28
H@a12K)<2;UcA9\0b81:Y),B5]\bNfS)e4).QaD_[][0)X/c)0g+S,U[(FC<./?@
N(&2E5^K+MW:Te_UKg5);<RR?,<?LZS@#?YLLcC(BcB-@IT,77<UJ^8M,H5:0S/4
A2BK:Y0Y>X1I\P,cOM^Y6TTcM&.6V(<?GO[3\;W/-C?N0aG=fgM45VJ33g3Edd-W
Me2A0(NUg#F(M6+:Y(+_cNK-)6EW=H]A:VBX:;Y0,RfPMG4EOPO:D?X<8-b>ePdM
S+_bXa3U)5dEP^?LY^fMY0SIP<,IJ)gS#IJ#6e>ce>f3?bKc>6+]XPJIJ80>@D_F
P.d]2W,a.L2C#?_/G>R#CZ;[VDL(5/0OC]3G\R^]5U>[X@HIV5?+I=HK=,b2?g1Q
dU9^1f+>S0d;G@.AM8f)EA]T>J1PP5OZ(>1,)cg:<VgB_[-557(\TL6b#Q/LHNd_
2HJ9Z<74FO=OWUJ#RZb]-#>W5_&)dU2XLga;3P3X?WL2;LA-V98GG#b,fSTK;cCY
_-61cBTcV\Z_aV.N=3^9[(9CHDTE+Z,0;YT60b=Zg8K3FNZ3R]58-58g1[N9cP)]
/AJVFX8XAZ8HL+E[+dRMMXBVgb-IB>M^5-CMPb\aM]=W.AZ=22gR<TB3Xg:W6)MJ
ZC&0a&&GU(B(]\a^2D,>?-1M+1g^3LX968Q-E62CM3L)IR(O:IJ>eVHGD;A?fJ-W
2G&Y6=?@0PHFJ<IM.f0,cC(JTM?K81+V(^&>S@U>e]J>BW0T:eGI+U63E9cXWgaF
3:Oc@UUfV(M=-OdDL,.@@dX.7OOC,N/DYYS,8HU_#BIfJg8Oc90^_)?X0GG&K,O,
&9X+YP/b@>W);9J^JX3\#I1ZgXTZ5W5Vb3UMGP>-b9=[:?.>/(2\1R[(39]M^7;=
F[O9D-dCB),SaAY(7Bfc\Y2OH+;GK+.BQ3a?O1KB5]B=>)gW;/]GM_Q[8[S<2)EO
L0X??^,\ZX47289=HLPL3V2c/GE,^7TA?9b:X,_A/NI9JV:Cd/938F;PI;F0b.dC
R_D8.FAAQe1FL6.YU;Z+@5a>(b8NdYb>d=+c,E)M(SOK@HSSH0O.U#=3OYb(]XfA
GFfg3P6g<14V(QS_b\CQ-[PHX;/a\\McUI:JUOA1V\7e+9&0U)I22&6TX<X2V:SA
WX^,P>.S_3>45RC+7DBeC1ULTaFf</#CJ,EK/=SKR>>ZCK,gIaA<ZR5.;S,>L?R4
CQ#-A@fA2Mf-FLb-O\XRCNSRG)I,fN-\1T(>+(L[=8XE5a?RfJB&..,bUB8Cf]8H
/G?XA8:_N9>[L^YV:4dYG_N[<7b:<<gc:M0L((VL\:J2D)N?;<R:I,CLgN^EA2S=
R</+[@HYG:K1Bd;S6R@&>LB&:Q@Wg(@0cGB[A_Ya:a[f+/PT8AA&QN<^0_42g0:f
]929&ac2^-(;_.d0Ie\EP-F\8JQR[/b)Jc-IYEL@I,8/1e>^\0=Z3b25;52e4/UT
T=QcAK[cN=6SM\UO>VeB\8DEJB#)U2?BIVd9U<)I^W>JZ[+=eeAS]>>4R@VP)ZU>
N==-JHBbHK-?RD7DAYP0:W]caKU)=M?fN[IB,:@90LW?5a<XQ6@+[MA47<,]14O;
\&(<T<MQ3H9D[gH=P[R1NC3I;Z_5Bd4/Q<YOeVC+@HSaZV4Z8@X3IC2@SV-);VU?
\I0Q0O[CD86O15J\\,>^Dc^YN<0>_G/HDJIJ5DT#;W[H,V7a.=QWZ.Z<=/O(GSVV
K->YTFgb:HWTPLa4-,LH=.?;Lf77UI:Qa&27H08U.I.R.5^\f3W7a_SBD&.<./R4
F=fO\gOXK;8-dJ4cN^99AK2:EFaJ@1L.RD2D3X8dbW,Ra?>@T7OCe<SY6V-\GcYN
^1Y1ccf+aN@H,GQO1C[TdZHELA2@W:J;,N1K#2#Z-4?A@OVKAVYgNbg)L=^,JX.1
VT<<Q>66F7AdXQ5GJU3^ZFL)1[6?U.^&_QJD,>Ug?=HAK1XIeb#QbCD^)UF?-)^a
6d@E^V_=f\MP.cU@7-#B-/#HDSb;e4Kbe^(]QV;_N3L>8X/B&9aUf8#.E1MRfUGZ
Sb8S-5]LV>KOI31>D?O&f8&V-#3_AJE+ZE+I:eCD@GCaeS4YP][;<XN?eKXXQ;7?
&;([9FDTR-XSQ[5AJ\=I^O^8>IFcA8-e)Ua\^g2#.7<I0A>IRcD&GXbPXCNT,/+Z
B8:&8_eXGFF^&0N;RH+D-KD@Veb/VL+,3F_M6\X:V<W2\U^:b4.K)fL9GdD&,YN9
U0O8cS4#E1W<,?Na&K./_F3U17We5N4TB3fH>1,Q+SeFIBEaKbD,0,gIAP5fVa?e
G8gCOPYEOBN:]IPW\HD(KW[8)?_9G-@+;_1g]^]c0YC?_9V[VTTR3C..27JZ(LOA
@SZJ^:=IOSECQ]aNdPLN1#12+Hf1QRgWP-@S^LBIFCMCcP09gU5J[M/M+8+2;7TK
a[DZacV_e_aaU]9E#N#D05I(,-Qg8VGc9/cSa]N[_;]+b6f#COKT3F]_6?9/d:(0
TI:?0OAH^=97]WD29ZKc?cT&Z.2[F8)>1+A1XJT8fe]L>N+@1Q-?[]=G(DcZ]_L6
>DJ8YJN_WP\EL(d8Y8STe,.@,f8[g^0(PBTGJL#J+R]N+H1=G3P+_\A.1YcH,gPC
1;RHH#X/\BKKK#C68M)9(>1\]N30ff,^DVSM<;T8,G0;gLM8W\3XgG>[U@4XXSF=
BF252M82IPQW@MYL>K7^3#D?@C>,7LCP>C2^N.MNZBZRg^QbGZ\^g+97VEHU^70f
/^FT.#U+6)f6>;W<BNK_I3.-9-_2@]b@DI:]7YEg[/70Q6Y2I+)5cfBFe,^1=?+S
e^KX46C[@f5d0<DHP<::]W]0##LZZ]a5_Me7O96N)T^]T#Je.6SAQH8e2;HQO>+W
0=YB11RCAC2,2M=Aa+^3VD7DQA.SBfLYM.L:V^:U=Z[P=Q2OdE.9fUELf9Ff3g6P
#X\Ce8)SEF-WdQ5OR@)@-?0V2MVR3e4E7O([9U(/7OU<AKE521Tc+5U8cb]]:bG5
f_W_-IJg?6-)U&XC;J8bGZQd@88YIg_D##GBc)S:WDEPNKXc#H<)7?7dH)=(R&GN
K\AX\F?aOC-:UDT)27YM2_.d<[SV2Vf..7+)e91bL.ZT8&HO[PZJTD<+:fB].=-E
0O\d_?3J:;,FZ,\18MfQ3ZgaTN>,QZL2&5.Qb^8BJUHOgF/8G4SF&N[_4[P8SIJ.
)5L9JfX]+K<59=7&:L3\?8ZC)VeR&XYP.6)WfdT9f8/gJ#@4/;U[[ZZO.9;^bH9b
_d0E#P#[]L93\344aK+5T>&5,[XZ[)#BO9QXF(>cQbd/ZNKX>@N?,_7OLFEAWf7<
_9:?5;??:YCgPNY45SRE^W/O2RADFce@bG_2>9SBe/8c?Jf=GJ[eA)N8JV8,,];-
.^L;R(K9JJ[V0dfG/M.DDC7^1GDb>Bb#+0;eXLPKEF@YZD76W&/4.#(@>OV@Z84_
8HX<@E0dAG.6a6b]HQ?5:QVW;>3JOUMK821[2U,:<X7]BVcRb9\/0d_11)S8FfZ5
R&TC2HP7?=0e#)R;RWV&@<)?58P,aPGS]8G>V2@XF=Z=CP>RZNgfY>)Le^3[aDcN
(1/,#SYgb9I4&a=<ec6PE.=?4S#U\HK&G=a./_B+B#_G-1KT\PA(S/H>a2[P?F.I
?,V@;J3FCKG;_[7g[8QKBgR?T<YO(:dPafO,[G&/@VPN#:C&dWX:8RH)UC<)+,8K
]NMWc=V8-=G@(H;SVZT(>AYH;1N>LV1A.PAg\4ZUHO8<A)bbd#g:\gY/:HF6RZa4
aCITEMZ-KW05OQaPM,+8/e2Q,46d;g(2>63gI\HKe8SIe8;gf93HXU]0R^V(U\,(
0NV_:fD=/JV][_>bH<J;KJ.[F1[99CeeT478_Y)(RJcFQIJC2&W/W?Ac6Z:LGZ]C
X8Y&:W/=@gf;,-]=S]PZ-B)NgOZ>JR)X^W9,W-K0@O7_d^Ma9JI,(_O):dU136:7
@C,W#9-d?O[BBA;0:XWE9B=BCEB6SYCMT#C=J97bc@gfCW?O88^8UWFf0H60Se=I
9eCF)3gPcL&=6X)S]X;Oa<P3Y9M7Tc0[H?#Z>Z1e+[E+&c)NV]Fb([e#,-1514AU
RP4L<OV\@_-E6B3\[^JRV703V#+(KL6Q,11#V3;K=EeJ.b:(1HJ\P);^[VeW]:7F
aUIbT\/-N(?bK#aaMK?FeD2b^SFH^e)>e&3IGFQO66(B,B=R>E;UT@OT=OK5OP?/
XW)DDe3T16KD-J^c[KL5C(:4<eY7BR#\H9AC/;?ZR9QIU6#4C1+cd)N_WaE]1.Z8
N/5)^P\/)?RKIc<P5,KP7a7/P;d+A(a;2T\S;95LW(42\H>[Lg,50516RQgWVXH=
OH(/I4H]<XK)11?_H6M;V#-9]gFa\S9g[G?>IC)5L,A5K(f((72C5Y#d\EHOCW)V
>cWG4^c-NUYQOdN-PZ-&J.0J+1TQQd4Rf&[<LbU=)DM04F8R?f<.<JF+XBV>A5MU
eA@eF&O@]D<g,7_MPL_EQ]LD]W0X]3CKeb+,12f])^\9aZTVG;aA,][M&29?;0)g
f:^Nd76H5)+/f##;&^>;1^#J^(OJY73d3R/.XMSO9/>6Ag,A<Y_PEOR2FE-;=6/E
[#;dZ4X(Kee8Aa;>D;;:[+4-EeG?-BA?61gV@[/.0V)aaDXZeDM7CU(P03JNU[&@
Z=0F4#\LXL<^R@B/4ZX:1MMGEc:B[/PTRP3E;-QT<8F8_CURRI]c38DN2FY77PM0
O3()TQ@55\-D]c&BbWId9gZCJL_c?X:B/9<];b,aR=@YB-3d^C=I\@FYVbN.2_WL
VU>0<Z5U8G75fSA:8AcA728P\L4Z_b@_9,:UY\AGC/\=Q\4=74IYL8O<=9>2VCba
31KP>HZ9HAM\7FV@d+e>R9D617TX.OC4a:dA?b0H.^L<CZdSJ5KIH#4_>(]NSZIB
;=\0FX_+1NMS8<0C\;L+<6aY0]H3cOSH<H3K5J/.8O3F),B7WRfCeNWN])[/Z0&(
<E#Ob1BEC0?\d;M5O_<5:OWN.[VZdQMbF(I&M]4X+.27SF/OZ[Z4f70;H@N.SFT,
QJWdNFJW3IAMK(d#.E[NUYX81PT[La6<1Y8>W2UEJ^?@:DZaCC)1O7+MS-;__<#^
2?,M7]cbCc@ND6Q+AU49:&A&O?=1bgV&M>;7.,OG^3CN^AQCGY\Z5E8bZ<DHa[5N
YEYGd19>d0?>N[K4PU[MWg[:E_9JX<TDc)Vb6M<:La7EaG=WbJ<BG3K:6IIC.>@8
dGCC<R6f@/<5A\0XHQD\X(a_Af6aB@7-8DDV_:fX<3Q;6HRX8;C8BHXI(_X^Ga1]
^Z.?g?.RK4&97MB&PL,6KDW^G]H&S8=E?&MTXI#b?7ZH=1Fegd16gK7_\gCP9N50
^CLHDOM\,aNT^9^GWP.a:eIA4-cBT\Be(&.V\X1fS7g6W_H0EK.5[f^;QHM2X(L&
F]2<H>UefF/C,,F)b+>/I>0\-6Ic.4Y7B2ZYcG9F9;9Rgf#[EZOF;(/aDI]Id;DC
-Wb>/(JD8-@BH-Nd=LZJYeV+:V91BP]DIO#/ME7LXP-3BG176O#@+#\WC4V-<\^7
)8XH..VZfeFBKYLD5WI8;_X7MAZc5@HQ.H&-\Z996H]Le&&R[>DbPG/6VZF2(GN?
M.(SAB4D^4PPVV#<\f^04T3=+J.ZYg^E@Pa9I7RFE(_]&gIT2Y]4(N,_IW9b]0VA
OFGNZ>PSaSP&(_47gWgL[G46/-_.Ec>YDLb/1N^[#DK01=8V7,]IQ\EcaCR0NQ^6
C-5=?d(?@5>A&[KE8TD##+a(=F])fISd#23UK4(.YIWO@@)<gO\O<=6g:[BN[Z8#
N0f8.I;JbQ9]G/6G8??F>2X\_CSYe(>:GG=.__C?R2NA8<<X5=_R0Zb.(aVZ;JeG
eZ@5WgDYNBHI8WKeY\fKI5_[RO]YcVe3/.;#L:O1Se1+UV/Z.OQHZc/1R6dA]bf]
;g:>QbR=f^e5P=DU;eII1HCC2N6&0GOf6W0aVaJ4/)D7aUa5<O.X2K+5/eDT>39C
LcKaW(,bV1\&d=3U\FeP/RX7C[@#<TFH[6-7PV<0<>NV#WPeYD<+ccYQ4WHN@,_J
[^#W[EFC_?_>1?Pe#N:bV[1P0.HQ0V=C4;V][9/G2UQKJX0#>-IX=I)W+P2&U?S/
SQQVH_6^D0fX\AB>Xc.WUWb4]-_AHHUBff_P.HJDfOcP^X31(fCZU3>Z@\6\Ud@/
L0K=9e^V+\>3L?NR>:1QRObNF.)3E[/VZIC)Sd7AK65SPY,+)BD4MVf/OIZ#M)&P
)GTI7.[UYef],)JIZQD6PD_L_JdY:K5>CFJ[e^eHe=H?f[XQL[B@8c+33g^P\[DX
b44?LNCT7,C]=[1,D(G7eZfT7[OddaS,M-8JIX@Z:@B9fAd/9S7CXab8>:2[O]0Q
e2DI\O:NU(8W&HRHag>DJ^e_d+V<:9\MO..0QH]Y5ARL5K\BFgV9aMYD:?LgaSLg
>NO?MbaK?T&CVa_R7\Ra>Z;U&Lgb@NJdUZG[1P6)KFB#09?T\Gd5^bS,5KS,.WWB
V/ZLQ)B0J8==4VNY3DA\7FC=15Vd6XVL]^d-KNa81bUggf@^bVL_8US@Z=//,:SE
T&fS>O\1K<33RA<Hf,=TfFSe4;-AN8J:0H4c8N]Y)X<_bb<6>;gWg]_NA)@:W@WL
#V).F\?:WF8faa:X;O)(_[,B,PCec?CGT>EZ(T\K-Kd(UVRX/22R9cD)VGN0Ue36
[H9g50Ze8S?g3Cb^3:.8/R,2@>;V5A8Q4H2P=ZL:aQ>#NT0;BZ_QHJF,0[IBdb]f
^5>NZ1,NbX_G?;_+,P3&E=3d>8f[R^LYM+.c)+-7@C@DG<ab^J8b6[UL-d3>)CM9
S>3U?:5=+QbgfJB;,UaEU4fa31bZY,;K=7W_Mf2_gJ:cCg2+&ER\]Y(<K<O?eg<6
\].MI]g>^=BcXM.IU5K_P^SR59=7O9Y0[eS9O,P/cYC^a?]J=SCBC1:[JLCg4#7O
)S:K_5fOD4>;aaKNF;86@g.a;6/BHPGI(V)a7d7?R2(C:>V8g^],WD1<.WbB6?C3
_;8agXF<^dALLD.IQQ2B=LNg=-\c3C?6SKZc9=4\XY-V12IUQ3JS>=:-Z/S?&4Jc
ec\KPO78?b@MQ_-[HBf/S[1#YG/C(U;f7E]7L=7^5F+-T3b\/]4:dFPO(&99JWf[
A?PIUA316K4=0-H>46D>T:.(?JOVEI-#<0agA2M<)A;U^C7J=[fKU08<-M2TV2Q;
4gbP#=-f5CG#T-W5Yb02I5d/4&A&7\KKcJCg=.W>;1Y6B[Z7QaU7f7c[]DMV>H6+
5c1F6g36UC5DJS:/M<MJ6bB6N[VCRJ,X,[JNY]<c1d/:-_IUTcaHOWZX]YX\.BD,
YVWLDdW[/4\5;\N@3(8@/aY6Qc&>efOGY]O)?U+/]A=XS?&]e;<IK&RFZ@?3&RY-
BQEY#18RfZJE5WLF_DP@SMY[/Q:V.g6.-+K,<;UgT.X&]H#;0--CN=94O7BR;4Dg
1=6-4NGIgE(53\bc31=B5F2eg)OMMD=6H@?;,gHe+9UV)GNKdWgZEVS<B<4D?(_M
]OU.I6>M0ZA]N@fV,8+9WU><.(&VL>U]U(a];?Z.AG<3c2.?HM]2bP:G3)\c8bdV
]#D;DYM5dL/0_YL=?8D02DdRg^=QFD6TM0F[bX[)J_QeVb7:-):=OD/19EbO\(5d
KN@?Z2^UNXG&a<]YYBe,[?-W9cPY0(8ce+2R)E20>V(SM-,Q[59baRR?[T0Z4_bd
UL^0g5I7gT<;Y2Y.DP-AHOgFS+4#b]1\@C75-_DN7[M&c3F\0<29+cgc54Ib-a1G
g:RZM/MN+.Eg-H^=K\W[K.H,RMENIaH7P\;5<#/N7BB_;:/=6PUAPM/7V9TDSUF1
ReD0<K.-<XD2H;/#6.?7FMCg\>T/dYG9ZU9^4-P4eaQagQa8N:KK<:MIb5eK5.2M
4U<E<#/E<5a:C,E(bS7g[?9:@NBFD72S]a/;//?QYK/9b5K(c#6AEOcV.-ZgF_eM
gFN]WO-FbHPU<g6I+Tdc0;V/P9YJBXb<;[adZ.VbW+0H=J(]RAdIbV[0II;(\+0N
;agAPI.@c1d4Ke2]C-_=:H2Y,VFVC3)197(P&TW4>XJXIS@cIg7#-c-7[Cb-^fFg
N/AI>&\E>.7C<A0>S8e(CSYPAS2UU+#e9D#NCc?[+2KbF8ga[,dGF-/aLB=1-;[L
:TM7)EXUO\gS@80fITD,:&+#\eJG#,ff;b].49OA+0U/J-R0(F,)>@X:+;QNf/DD
5#e1KM)K=4FGLK4Gb@aK5L76.G2-?RBVbN;U1NHM]F3=J]dXO+FWQaCNGb[6Z)IK
Xg<PKS8^VP9.g#UG&03#O<V=EEM51dZ_Sg\&+GeWP<@Z\><2_0baC<R7SO:c]@O#
QR68GaJ(LKGW0V5f/3aHE<>)S.[H)8KNO\(7[d@1/dSB[^g,M2Y?gJ\Pdg0Z:DOL
HH-9FQHJJ3W1ZMag=_V@I:^fU9/AX8+VebAL[=>HZM(6>O+?g<R-P,H?]1E(CM0_
-\QQNLKc^2M7@/M?T3G9J[QLD:@dXT6-B+-7U1A5b3_M5<H//WLK6BI_\,60C:?C
H,C:N9,D,CC3^0d?Kd\#cKK7fcMKF>M@+(H8gTABd&MC:5;]:J)aE,>3.Nc&ZFC&
=f0YV;c.XDQ.^KZ?B12A3=O,[]8/G)WA_ETMb5IF19+&&U@SD()02:29;fM#eW)X
>>]a<[S[]@FVEMX=TSb3V@:[>JOeFQ:Yb[MU)#2?U=C@8Q&;,JR[N3@R^+[(.S=A
61g2L,<3/3K=8365?MJEC\ET<,2]/K84_3KU<CJ+9[+:]DNX>^C,f+0VVQb20^Za
RdcDWPI^,Q#B3KQZYfR7LL:+gP<AC.4X/ZR\>9^ga[dE_gAQ;DK0+U4d&_LJbO?\
=(Vd8HHF1U;DPN.a[Hcb3GU>:^[DR2,MZJ#c>.8THXKC3ETb=6HMF;3_M2E^4Z/e
5=UN&f@X96UcO53VH5dB,[^XO(JFUPJe2OY,[B6@]?,Ib_JGUNGV(LXDgaKGDQ,?
NJNL-T#6(#cB<1I7fXDAGYY261,Kcea;aE65>W3fXTC6Z>P/1LZ-e6V]+G+XOd<>
.=0bSFd0,BSC/8_RdA(8T3U#)H(YY8.L;dN&Sg_@gWV-?cA_/SR4c\4;73e,W45)
9]AaF?+5Xb:_]0]dE>>LSY7g=TDZ0(QV=&#MgSDP7^@1M.;S(JCWUX=^HN-Qe\9#
0.6-::0R^U23V)+C=R1NQTIVKKE5<c2738\a[?@^\^4+/3aJH.cHHa/S+OKGIKcK
);c<X8?>7^\1b2O7.LgO0FXN7(QC;?B2g4#5+ITI\d@_<g9\bDc5(IMbWV@NS0YP
))#4cf,eNL5aRBD.8P32S5/>c^=5OA37T-beg_\:/LXIJ(:;dS2XWEP(Z=>?P,<=
gg#B1Gb6&4IZ(^YVN8dI21FT;[S>9e^KG.W+EZNE@(d^6:gfTe+(KZ?8^:dgfH+B
M3e@S,B8:<:P#O+&R]4cZQeN5WYB^UGPJACQ0;2&d<Q^D?8:aS>9>a<0g_]5KOR.
X18XBMCFN\,DDa_GO5e&S[S52b@GXS.7:84)[9MRa:7;GdJS&]GVcK1W&A>0(a8?
)Hc1.f_e,G&^3&#QIAM4NCG)Q,Ybe):WT];7C@1DH67FZ+PM[bY9LY\dEZg5VcPc
Y:2#^A&U4d5Q;<6^bfZ.X-^5A_E@SVgFPc;]WA^BL:).?M5^OZ<-R@FYLe4Ea4Uc
4)KWINV8P;67>G9C0TI4([47;^Zc))E(6):FTM:\(Zd7aUULN<Kd(:]ZC.)G+A3S
=QA6IX.@(J+ba\<f)?^4Q&ME?G88791F9BT5fI(EbQ1?b>W-WNB-IY9C]CcNY-8^
,-4,BATI+\f_8XPKUV3Ca25N4R=/FQ5F:+5<A3f6OCN3&7#g>FcKZLYBP=E?DS6G
S3KK9<5,)1@g]AE2CJ@.g]S=)Idb\,.JJ()9M4&EAdRXF-MT8+4I+,=da?TE:6Hc
H?XU>A#dPNXDA_.>dE0L2=SRIUgHcc>OgN?DWDLEH1GY&FQW[^R)f+&8LZS((S/Q
VPEReYGd34.J=9F3_VFR4JQf]PbaQ8\HSe+B/7e-GIM)3aG-++=6./KM^eU9C8YG
I&K-LcKTHQ4PeBdaP);=_O^6NVJX+-<E;1fHea?-K@G41Bbb7Z7#a9AZf4#?6gc(
cSgW_R@7Le8LXg\:ceE>Rae7E13F]9O-/T]gXA[IWFFILZ:?W08>#?&e5(TR0YOW
WJP\X@-Jf1LI(4?(DZ9#Cg>DOS3KWP72Z?ZU&)=IOPE33HZWFgc-.F-_5F<Lg,-N
OQ^X)5+FEHE0(GKcS>+O0-PJC(<+faGM.7Fa_.C-D]-M1c@+1#>CH(Xa4C8cLc7/
YLO@d)CPQ8,H37F=B15D0U^Sd-O)9A@):e\)ECDXUc5e7MATFYR8S&IXY#E.-R)B
\TL_IOF#^YB/,c98FYI::<+80gPFD2U:IMK#/,P7Q<6A+S;US2)4=e\4)YF2Z_VP
dXQ&JfX0P;g#T,TP;=XE:S5S=g31MOfd1:b7:g#OE.M=^-K+ef2QGE@\DcIe\f&Y
I^1I_\c8Y,f>(PV)P9;a7g\1]4?7?OdK24ZAg<;3J&MU[>I5g-3U/H3H,T+>^e^#
W72+1>W7:_6gaYZGZZE2:(ZC<[\fc-GF5;EE.YSbR50C,Jc-DKLY.E&AR\(g>;_G
U@g^SJ&XDBJL3MR>0R_Mfe[TO1Z:+G@5\6?EP70[37Ta2:QFLdVI5@-Ca)-cBGR:
R4;V&H?Ra#+W<bZdW2?(\#,3PcZ<+:?1=^?-K:WOV?(Z_,62b#):dLgW@GbJYZKJ
1dU:a_a^=NT.XH=<C.:ABb8?&S;c79E#a)>JO]2NQ#N_Y5e^#V&4U99c.6C_MU4V
UH902O9Q.4B>;BX>^?5LEQ4@7D=,>5fPL#G]aW8D.=V-E]VL[LPJSN-KZd-RL,>9
WB0WXgH8\6G8^(C\#LABc#9-FZ_g[KN;53?Z<aNC#BEIK&[2D^/g0<J>PD4<YV_7
6&W^D&HJ8@gMVPYV\5]C.&cB&,SOQ?>36VdB^TIY\]V?;G#(O^5Q(K5/ff?0MK#[
JD:YB:f:1;Wf&0EU.G(]g0Ma?AJ?S-(G36(.I#)NgQU@S.TY^dQ26E)^<1(;#R5M
aT93&5+\VNTbA7PV+F1C@H5<OBQ5W18/XFH;8U734d,R;8X#gg2eHIOU]SII\C+?
Y.-GS^L?Te7,34;YAX:(2@fP9ZN<P+J+\5:aB\EaUKU1Mf(]YNN3f;4<?+74Mb+N
acEOa1?&1F[-Zf4KMe?,OgU?/HEZ<7@E+@XNW-a<(#Fg&66#E.]OUbf,UdXXA?GN
&BD\BAWAPGc;Z2XJ>_S_9;#]Rg9@aG;_.0cCU-Hf-]d;OG1@IC:)>(7:bdG03:BG
D9ZU6FO4EQ_+<aT8J7VVZDOF</404Z=C#XJf5Pb>eXA&>;Y6)Y+4c-QEP8U3TZ>K
VU#R?1T>P7)S[W8B:SfPDP[6A<aSE1b1[I#G0#Uc5b#.d7E;C1ZJ678N[E@BM>Y+
9>:a62T-EGQ;VGW4)RRT&_0<2+TDECc8Bf6e-FNdbX,7JKfbL2/eTJNY\XaKWZf:
3cX]QY7[gC?XHAfO03:B]de5C0[XR]RP>2P_D>UALUPZfYU4bEdL\0,HX[6D),Ac
MPM[1Hb8QbJgIBQ</XS\U6S:\&Uc90MC@=R[Ug.:b=cG#XOcE:0H5Ggd=&+^8Y+4
bIL/bE9E4ZaJf1OaIR-(@Tc_1J@Cf^^#QIPIH(C-&Y[CE/>MO.+<^gQ5<S)8P@X;
b_^@=6+&0[Za/f(F8.M8BL-g,-B8aV.[P63H57adg(7I2fMP=U<9aXTUCFP\[#b9
.8(G+e)JX7e-YTfLLO@.NLYP=[L>-(INg9Dbe@A3N]]]EJa##ca;SBL\K[46[-:<
7AZb78.Mf(F=LD;C6EF1T[YE23WV?7,Q)X+g@+MJ\?#=(10:<@CF55cK&.Pb6_Wf
ABcOOgZ44J(0U3W_D)N_+\=6F__#f\?FgUWO-5Q6^<\46/<WML[Ca>8C@)ZC2W\3
C5N0(ZFbcPA^#B4gFc#]T,[ORK=M)SH=4e-@X2GZP(G_>fXSO=W&e?TB/)JCM^DI
JbBb@R+eeDgca#aLLcR+bWaWWG@a,JAd]HTF5(P_:YYRE]=cLYPUE1bfUEH5_);d
<^f;a04=ZY=a@<)\#dKM;D.4>_S8JUO/CSE+2[_0[Vd=U3,2,>DJG=RFME+f?WKS
95[-Z(]ed?ZB>G^2gV[KGX^.D3aH8MJB)8D_/BHOe9.C(#<BYQ8R1,Og>N6SJ0AF
V>I7,M+G?RABQR)&()X/OaE#>__JYA)4Rf_cB>Q329Af<09#UX\Pa38;1UK@7fZQ
?P[M0FbY,WXSd&eX\ga9,.Ec9f0^B<@Z#3gWD)I)g\\ET6b<U3,b5Y>XNMLG4?)C
<Sg3CbFPWJ;UQ:.-cCCEGP(YaUWU@AXK7J+gDFGI#bCf3,7UR4ccaae<_M7>>_0&
#5NcgYYIWg?K/ZCZ<a1g0/DId6ZcW#g,;DHHQ,9-=H>g9T-2<Z[X=4P]CbGL_?GJ
AM\82+UVWL#Y/c1O)7IR^XdJ1#aY1+gM@OCa@G5G_bZ<L76c=@SI:8Xb2Y:A7T?W
g[M0FR()WfN\.b\RcP:G,LSF71X]^L5Wb:cG2ICC>^&_Ned]XPOc?UcL;VO9]&AW
12TSZ>6(&I7Lc.eNITg#dgdD91PFbV_=cW2DFZ\Mb[=LFQI\[CAM#Z;CGcXPWeL9
0BFeBERLb^CfN[;3(bLC(,@WJaJg>A5JQGG_(=U.;gE@+6bNbgW1W@4.T-QP)S5^
F]TCX7AS8(+]T,FbKLY^J/a80[P6?[4L7EWW[eFeMcT&bGPZAf[CX]cFdA@Nb#@H
f1^4]XF\UC-58UW-Q(:#f=d+I[KVdB02-S[]QA\\85L_Y#;ETb;/RK\C6a9K[#G_
bMBb@5&H]XK[-U@VR5G\BYg/]N(8eb+H]]UaQD+F[]8X:@P_+KAH0F7/e12LE^B1
->Q3G(H+Z7UE]GH.d)=R(2beZ/?]6-O(VTF:T#&dOCf@Qg)b9>5J1?MU)6QWKXVR
7RUY.<4+OSA&TGS=M]B(2RK?-MH=MQf.//D91M1B6g<g6QXQ2Q\T+0G7CM.6HJVE
\B\>>DZEc3&1N6S?F7QZX#M2]:59);#</V_(X)M.F&C_SE+3B2[=VB?;E;b#b/>9
/F9H?RGY8UC]UAQb0;bN<aF.5W5D2-_5#Jg=H&/32dV),OJ<HBP.L8Ka]EGE0Xe]
JCSNGJWeT+5,+9N<&dcK(JJ@1G0Q]25[dEYRDPN:MX00G(Y9-UWJcWH\VcT:@[IP
;MM03NaQFKBPX.?<NcHMMDd#CEA8H;;H((T@ef/>]8?K6_-2KTBN;P<5FT,-L.ce
^cDB2,3GLO;57cPS<fZ:;J/-G<D:,Y[0.[/(3W=X>0M]3.cI:/0#<(1=-C@J-)UW
]/?BO:?_12X-JVZgH,b)?-B7JN0VBf/2NB1](KOX>KDa&=@gRUKe2d,2/BfKY1D/
E(]&+07(42.0e@4M5LTCRENa:M[N-VTFeGJ?:^@(3Z6A<VBbYKdJ(,=VZ8Lgd)fJ
8_1&<FNTZM1cF7FTg-Y_5N@E6TeP^8>L_CF_[>[Jd9gDN\/_H(ZVD;f5_Q.).X^M
R0A^@Ta+RC^Z,V#b>HJX</RdFI6/6TL0HA++1f;ZP3JFF:X\[/;7FE>KV21G?:M=
#P(1Sg;G1S>0W)D#N1G./A34O]T;K#=W77;;@BH3@B85MdW8MGeJeOc:(VG-eI(]
R2@E/gI),9SG0I#23K=gRd#I5]CMa36B63/PI2BI^2N-bKG1D7,a:J1]J=_g38I6
ZQ)\(UBTG\DG@T3g2C&R<bE#U&?YHBM@N@I(A_8-C,R(9VN(D-][GJBdL#;0M8@/
=^5A/G1aK84QgS@2NCPL3LX=I/W#O_@O<93(CJ@L.ZGTO@.N,M:Rg)8MA_D\FDC;
L)PZ]7XJZaHHW#LSCQ0@X/Q@d,GYF..+H^OWc<B,GV4;D/YaaGHWN#SD=ITVG?5L
L.&Rf13C8E1>PZ=614U>7>.ZP#)G;8/=LN4e4^(NA89A^X>]9;dJE^>^J:D=R7\3
VRXK5EAf(A9,:dQ.]d2UF>H1:e]DH=:O_bV[gE\T#>GO+W_]_aIDWfSBHQ5/?YLY
e@>MQ/&6I@#7[R)T@1]Yb[:/AQdKJ#0G-.P8.U1CB2F,^KDWY+[>SO&1YaOUa/NT
19^>+g/+AW;ZDM2E(P<JQ,]U=5HV/0eaVAQ\8=WdSg&\C3U>P/c7\.1QKHf5W;F,
g,^L&e5bY6P]\aUXTbD<[-,^gG_72X,4,3/882[C\8KgOLOd8ANTNd[CUMBRbWM?
Y2O3E2WdAL/&5/=IO:NdHfK5^fX-&&WO=&DbU1S;&0Q56>c=EHU]7Tc(P\DRB[;_
9E&(.+L#LO3<CJC1K8&6-NHf@QEc\].(I(;Y@R,7>+Y.7Ra6^3fL8d^76^Ma(+b8
SEWU+?W,Bg(I?BD1:>W)b3@]W8P4]cV81X#C36JG^fL)Zb9>Bd]:M-AfX?,Z0fMJ
C2&8<W=K])K^YE>SDeDMcSA-Y-6&R?:OC2OP?MU@18J]0DO^63,<?BNL[>65KJVC
0WeG2b:a;bfb7UafI^.F4HD,8gfU[T(EE5UT7=_97e#cDC^5;,8S\a[-;20N(FNR
E6/8Z7#W:JYEfJ-A5CB=<b2S/TA^^NDCX^e?gN)(bNZ4dC):E),HUWI?.>5;cGCN
Z^Qgd(ZbGKbO#BWaXA4^MF(<CO+)f3d;EU&42::X50#6&X4:/L,S0MX7=:53YDd-
f9Eac<41ER5MN>IIA]_+XDJT&<H((3;8NacRe_:_RP57SBMR#6+b&eL4L\Z?KUW<
4F9&AZ,I?WXA>@Ga3/.L-KA\?K,2?784)E==NE/]I66^(^IIZ#f-d78a:EdSe:D/
6VVXK92=.MOIJG:b2UQd7<cc&BT^Ic^A)Cc1-K7>eG6C;IG-34GUXFe.V=(9K9@F
+UU<#-H\VfGQQ#7(5C^Pg9DU8^5JZfS_d?f99Z4N1\&)dLb.AHXd^aVZR1GQJ_Pg
KA28ES(679LX?@#cbDfeP?&X\A]eaUO0?RZ-RX.KLMJ>/GUc0\=gHI\c.Y,dgU,>
U8\bJW/SAcAV9S]97&3#:HM2CGZM1B6R>e81^R=Ib69,S].NDEX7D7=JK^D/f/TR
P1A@bL@1RK1=W0=?/cZf?#-R(DMbR^]&/KIWg<Je:d12PF5WD[]?I>\U:]&eA/(/
KAZe=HO0QcK5A;AD>0+eWg2f<:_cD\Y##F(FQ--_9K^CC0P3@IUE38W6WSM?&L6D
fRU9F-bD^TO6L:b9[2?1SD0\R6M6I(3Q2(/I]#]eP@)^A/aI]5KVYI]C;Zb_=[D&
3)8F)C,c4F,NVG=_07?aU-b4/L=OB3+5Ag-g2VR@@8)Cc250IJ98]O+DW:RMGLg;
PB5eLc-_<aH10.H:_Q2W8211OJ<AZcVg#+K&QW_+MFB&?59+JI#>82+6CYgDa(KL
4_Z^.6?M/5:NfeMZU)-U7Ne4<fD5L-b6IG.6dQ9]9NFg>@Ab06/,=A[,5;W(I#A[
M..^ffSO5:B@W;eSO6;H90=HOE3@9KX0MYN6/C+7bcL=d@E<]UgfE.[V/&>)L8A=
LTQ_aDf3-G]aZN,,.NXA@V]V55=0TaeF3-LT,KDBfJ;gR^Ud30M>8SRAV;:81RgP
Y9)<6P#S9)&=L==8;LT#A;c)?U#J(ZdT)?Gg^4ND/cHVK#IQ<+2eBJ9_M;eeR3KQ
TQR6D@\81IINQMFQd-)2SAO5_.ATK&6f#gb=P5N]@e+F>IA6CM85K#QU<6DD=;<X
gVHW1gLSE;]Lc]H[#33P<^e[TV:Fdb9Ae@=FJR^]7R?EE3.L7W[:XdV+;FG@+DO^
+XL=N-Xe7Q<..]<(?HQK#bX@P++-HVgB.61[E/82&6-_U3K/JH/Y\C0@R.H5O-(M
)R4_XeEU7[2AEBbT]F&2HDd04^-)CDH745X:bDM;>e,eRL(S,Y#1@3QSTGF,V.dg
,H]7&1:f&J3BccOJ<FMG-YUg8ZI3Q&:3#YQB^;NX4+?6H:IW8gKJ&G?6WSW;I,;-
>f-6X9GKN\;7X+HB0O#GHa<W0LG0JK&L3[ZAR_e9+WPES_M#6/fO.0^T=1,2:PW:
c0(9aW/1C(AYa0Sg=@V>@<eFcA91^9#1M>OFYfQ)&H:E3-@,S9;b><A15KZ.;;VA
MdU)SSJ.AC&._K<&C99a[;9#\BPS\9H_6>BA:MQ67WK\V:1&43B\&V>5eP:ZU==I
dFJ)=166(_IOc5X<-_V]gVF:V[=(7NWMe8G:E>U@QDSZ.9b[)\\c.OYEdce/c#<\
T3\+22/X_4IZ#aKS7Pcg>8U[.Q=bC125FKcRMOH@TUT#SI9c9WG6EAF:4T1U][EP
)Af.=W8[:43Q0A4TY?_JJgW]Z07a1)J0IA]F7]?;=_b#+4?T@3VcEI@e^#4V9]S\
GFUN2cbKCbG,K4BGMNaU?1:9PKbN,03F69:2]2E8bVg(3/?N/;/.eZ\Q11EXT6Z/
JW,\@;>91DaaT2&d2A<\Tb^A]bTEc[CE;I.U]1+^S]37R#79Ja<1ZcB_;3+<LgGd
GKS(<CID#LeX6]]Z;A?B[d2K?(B_CdcN>BA&HKeY:C+#[SY.9H8EfS:OeW)L/NTO
]3R_8/K2cU;d<\LF\]\eAgR(a6cCS?c<dNR.>7HV[XHG1JabSf7(&DXf@fG\0V>S
eZ^S=]TOT4fT2]M_@SW)O\d&JJ@>\c&C?72^=BKMcfT(P=-]8C(@d/PE3LZ].EBR
UDCJ)NB6)0:0Z]<[TO418V>S_6Qf-7]_G#2@-&O64bBNee=DV.6UU#\)?YggU2\+
b+c^<D3Z+D^HTBA3BI3CMRFE=EIB,?g)ALH4V)7(K-&H;X^4(P;?55UTb@\I\f],
.2Wb7P:aFY6AEU(b&BRW\0a\e.O:f@a4&=N^9,&&J2.6GgdXR]\#[DSc>gc#[6YY
1E,L7>T#\;IJa428R#&cER?):b]S&B#R3EZ;L6C>Y+03WccK_T=F^D[JB@JVdLPA
V6/,[HKC])@BV/X]>9;c,g##2A.3]_>1R_aUL2+BJ0YdM\^_[;[=]5WM<gQO_+YW
-f^IDRY)1R8cIZA__J@8XLBPKX#_M/3=ZTWP,:KMUH;e9\-7DI+3OX+8T::QV:69
[KD#OeDF(g17P^Y4_X?)LDIY87MR=9T,:\I1Jd<7EP<S(OXBEa8>+7VPXS?.;6:c
L3,MNaPO[3\=HN&P5GF<G9^Z8ZcZb4>/@W4=7(&KWY-,b\[Y00:1F\.PcF=3-W8T
(H.PJ0d,>30PO4e#B;),4+);KC_AMf[E1aY.9[U4^#7IDf12E3TUSZD0Y]3+?TNR
.3@P>UM;NVS>]+8/e-JJ/]H=VaKR#.CaM#Fe[bY(8>=>TWG@&fRF&J8Y[E\/TX&e
82R)aAf=I/()\(JfDYJcN:S#fTT-&FSOTS&a4[2gdJaaCMJ(P2H#?I:PWKGL=gLU
-Q8>0/Nf:7b[U?.WCM=AUI@2V,^#OG;K[[B<>@1B6:gKI8g.aA7Y\47:)I0>KOBJ
E]0)Q#XT<7SHFg?S2A;M3))^+JOdaG2ME#PM[4(6?b+Ka,28b\AeNcDIBF_4U<@S
ED?6@)Z5CfW:QA_^a;5S5&RHFa_Cb@[dCM0#&[=Ef@2_TX^VbI<Q0[NC_Y@9e]F-
U1WIG9;(VA-YM9U<AVN&WHDM41HL]9Z\V\:ZQ864KWb)fM]Ue-WILN<Xa<.OQQ)B
_XaXa9a#(B9IdS[b<IE_B.^7KVbV&c(Z<XQcC,g09gR?J27Nb8c[+ceC,Vge88eM
MD).:@]=W>Q-g(ed\DB4E_LSDY>)>NJQIVOT:YV;-3Ac_;/VVeBYW2E8:[Kb8Q9U
faOE@L5^G80V#\MEgAZ@KH)d+cU8=^UAERV3Y5@RN+]HAc)Z35@P;dV@V\Ua#Hdc
G4fKW6J:&^)e]D8:=,#T&OQ@?5C>Z<.>_Q13Dc,+.]\=[3R)(bK=F&#S<B=U@9[g
SES^EFN[/CD:V>RX5L^?NZVT/2]:0RJ^0=2;1CT;cO[>VU#aWFSZHMWcSRE9D[4C
fKRbY3N=)@05B34Q32f8+b&K>DSYBcM4TV:A\XQX.N2Y+F7g\gc9)\L^JYVHZDY[
aA.E3@Xc^@VKY\CeO.9fC(aSC16D&7C>/,Y2,E_ZQMKW9B_fCM+Y9/AbNEOc)5cM
PO>9FYS35a?:F7AC-1DW[c@/5P-)&;&#Oe#RC>\LXQ@?23QD=+)R<Vf\0B1B@YM5
IMFb,=SNC?5>]O5^d/-,2VO>aZ9e3(Z)TD&fGYTCAOd#3<?Ja3:+^\3[T+>RUcZb
I@cY5^Zb9;V):98_,Z6U&eRBM/N.1/.[G.LGF)@?4NVLe;;gg4Dg<WGF<C]^Ue@f
+ZZ<V]7e3J7=0CbaBgN.2AI-_OC6^8Q\(NeAH@]0WdO0c@a]85E4HIPc_]3Rd(_H
G@dBC7e6[R[RPM<+Yg2MZCJG3]5FYaLE.ANCecgBICeWNAJAZOA7[aF19fLd8^#1
NbST0L=XKQ>8=W_>HWVFZBD&d7Z;P;DH02YFF<P7O\LF#A[1da@.8S<d0?f3P8ZL
cN3R#J&]R-^+c,EYA-V[&>cM+IcDACOf:XE)]EcS@K/L,X[bdZB=_JK@Gb9E\1db
_I#-:LD]V7f,?JEHJYdR;P9Y^_DJQR&C.TcLDc)&Z5XS0;M[-HIQ5C03F3eS18(C
d,RP,C9R_?WTN=8eU9Y;,TfTF?dZ3T5b/UP<3XFG;CNT7RRI2[Q]BKWDX2S93g-g
7U704LXN16.1(]NbHKG,+eO7?[T=<H1^C95OCEM,3J,HD8,TO+-^a7FBSV>4-=-\
4P+0>>YQa#a]V(@S6-+O2)BQe\5(Ne:_N,U,C1cA>Iag-03.H@Yg?.4XGQ:eR)5D
O1?S(OI^S:TVVBAa)DFW@2]>&IgWQ>AA&D=+)K1Ub-HRRX,HOD7DE?[S@H/b+41,
fZ7^(@bKE[YVPgg+275>T,O3O-cC]@RBf;JXPUFVRN.<]4?U[EG4gX)bJ\@cB+</
\QFYg>e0^NP4?M.b7Bbf;3VHF086S@V_^V>RID4(AOd/Ag,[D2:;5F;gg\<\QWLd
/-\-7TMHaeZYdVZ7TNM1bQ+G7;E+cIT^QX+A>V?Z0B3GWcD]R/fSEB\587TOg8[J
RVN,APgCT=Kb^Y,9RO&1UaC\E&T4_W\N9@?Z3Ld(@G#[4AW&WfIBc&Na?MY@M7MC
3de#5R)RX]HEO1,V2EaKD(HEc,\,3YbY(Mb+5Eb=EPR#N3_HI]#UU9N[ZK2C[IL+
cO1(b2AKKeKA?3?:X9P=[\1A&]aO+b<QeRJ>db1K/50Z-aB,Tf4P;)1NXUFDdHYS
@S9d/MUR+2@0BGTI^f>6@/,4FJ[+fH(IY/75V[NO8aZE0SH&?E4R3@6aPPQ9TIA[
ZFe/#dG@7&gL)@fga>R2OK,)(Y^Y:R<\#aJdO\J)\W6CU_732d#LJF2439URe;gH
_XSOY)R+9]a@:&?bX#e(GGP1=161;?958NPK_X+9;M@b^6Y^VT3HbXOa0]-)V1-O
3V;[@&1,?LC[3eUUGS:MMZN3]eNP&7a_]G6:cZdL3dN3@(DFG>05VBfQ92dCGH.L
>c]SWH@UU>+>,=9DIc(LI??A.,FV<&5N3eV26f,We=_W4H:=++29GII+Y7,.,XJJ
@Q7+J2D(\6=Zd^[EO5:>-L1-A1KJ.,&=&?]:)A\)-Z]<N/^)]ZCPWDf&-#g2N/(S
d6HeAg;_YA\c<ES2&ITYUb<5OYTZT=&Ag1,6X9WF,@aXYbg^<JNU@QFPMa&1(I#/
A].9K]^]Y650X^]&][-O@a8,^M_]R;(78X34MV11K&@a0Wa>?QaFEdDd367/A-\H
4.M3][;>Q:8MB[XIgCASc62d^N5N?J110S@>W6/YYTMOLTI#N.fMH2=3>5Ue@M[8
Wd-GIA):#FY1Y=ZRC9CHY/;QKTOWQPKf_GU.Q^2#2M4FP769[E^g2[;_)aRYR=&5
55]ASaYe>4JEQgA]8EZ8C]CU6fP6g007E5TL3#==Q_H(P=]e]bWf3G?2Lf4821+)
]=+G^\PTT2]I@I3&71AP\73Kb0MGX^2E9FG?BTGeGgSVS:I.L[:cU3BTVf5+N,MD
?XS)R4Q#WYfD[/K7;B/VRfNBRB^M)KG-ANB][CbWMf0a[A3:dceFP>M,M/QBPTXB
\\CB3M^X9C;18PK3?^,(cU(DX6^\f3C)3:b7YbZNeM[APd+/7P,)3DXUNWeQ9FIF
QM/;[U431?T].e^H2I88/c\O>=#W?Fe3g2D9<O5@2e>I?(+TBBN\f]9XYWfYNfg9
?D8a^5[:93GYf1>L&Z-&J69?abbDfG7<?-<dM[6O?YO5=H0O=b4(/+V^UCP1UMJ<
9<MR(C9P[Q]899c:NV5\<>5@d34^IQ@.J8^c62bWAY4bdLA0/62[5PW#F.g@&)O.
LS?BGg.2\(0=K-Y+QN:ZL.UUaLBG]\#WbgW:;H.Y8UNDJ:09&Pb12?+RB(_:7@]A
aN]RcK^^UcBZbT?A&0e=;@80BD:+L/:WO;S,6Bg#a^8)cIXN;D3SZ81JO-ILG].(
9+;;1bEeCE?=.^cU#91e5:(a2[YD;Ta.Qf,^Z:04:/=DJVPE;I7LRd+D5B4IBNa<
K0+d.S.M[3(UHZ7]I2+3Re(NR440OA6-=B6JbaWAX86S+13+7dSdL,GXQf4D^K10
\9JbP6K&--cCA<\BQ)e9bMg.g+&cbFd?/EQ:8].):f_[bJ)P901eP-BgEICOg2:\
Qe11\>HS[G)RHV6\CZH3_X9,IC2JCN;&^;f=2YF9Q9/;c#D+#VH664M#[G<D/ffX
ROG,0JY6e[&)SK&(O@XJa&9C_^]fXG,dc\8^:dB,CW@fbeK9Y:4Jf07H/2NP-3fB
CQ(_(<@^3?_-+eWGW,0Y#Z(37g-<=BfEHRd#aV\\Qa:XZQ#6aC^BU,cR77Z3TMP=
M29MOP/gUT54ZK)g+3@0VBc<6aPZ/WH2]RC\F],MZa@D7)S)>#(Z/4V/(5+IRQ+8
01E-XU0;I=b]SFS.#&Lc^[E[D8&AFf1bX^Z^,-KV\Cd@2OJK_?&UZZ6C9bWN:gE2
_J?EB;5-5W>4,2K@1+-[K@D>9d74V+BA7A.Q6gL^RX;R9OKa<+N0g/.41LR-?L+C
0Hd.D(0N]BcfU=3)0/R==a/NZ^Cb72FSJH[U)ABG-FKR)fILb=XS;3/1\B3Q[;Q,
@2[7?H)A=AK5.1FN;[B+](KN(,XD:(@V@]L1HO,705;)@7=I,b-V4293X<Z5?Ea\
dUE+0TPH#7MQd^CEYRf@]-7e#&::O\WR:UY7ECID>T,7,@(:@NQDW4>H]O,?6PLF
]d2G,L/C07ZX=2M\#(Y7P6M9c;8PQ3@[&NKSOSc4EXgZMgN/O\94K:.Wd\YXf7@S
W?U<D@dRPTH?L47f?F.)Q&/dFa8g=(g&EY^#6EVdK,S08=^;X3F&B#)=7M)<\-+&
]:TPKZW4:K)7Y8bI>ZQDO_9P:Ma78+_W(9.L:0)0_;6:L/Q+;FNYA60:24F;f@>?
e4QW9++U40BR(KWT:HZM[gT()IJG9RZ6UXU&1fI^]G/5X=?TTe1fd:4QPR743B_I
R:(aWIHfZ6SJgS<+&4aP9SCWd+Vcd4f\\D;R8[O:ZE^Y5+:L/U3ZE[GH>:+FZbH4
K,9P\G@99CBWeZ[J6(]-d+ZZ\E9:R-0TfYR8d3N3N7B(QWeF0@[T3PU6.F0:_VO+
SDTe<NWT/b@)4SR(4HNKL_a\:5+5,dWI]S\GN:-PF0bT6__UHH1BQ=Da<9?P<K;f
J#0&],6W#Sa9=.O[;O9OL#>E3K23B3S##],Gb>I\aG-IV-2\XV79adX/5@:+U^Le
WUd@ZB4-aB&K?<ed5G(OTM7#?O.OSg&7082WYY0&2d;Ud,+TJNOP.0Kaa0D7UM+G
fBDY#?6>@=-3CWT/dO\V?>,2VNK8FB)Le4;aefQKVE2_4.SAW8DSJ;.D8F)OeR4L
=I0Y&T<eJ-@4Y&_8eV]dW)(-gG=^c16<>BB\dIP,0R=VU0,\4C0M2/Z&-Cb6]WS5
:g(aF(]&Ke+2&^[<BG09+U]]Z0JNbFKSMBc=Xc[/P9E?g9=4gB:=.PJ/V4=A\6YJ
.2:G&cT@O?d+A;TI4+:&0dRO\L=f1]@_#S/=fdIR5^XcYNIVM7&g.SOVf00eP.Ee
HAg]EYL=5O33.(LL^VfC8H-00F+DagB1b3ZX:<c#;#=?&WUZf\f26PP;M:?e^]M3
_619IT]8MM=[K<?HFH[PTgI2)&]D)Z5fQM&99]=FMB.1YGgERST@AFZRKEK^.H:@
Y>(J1A]7I)7@<gH40_C@<A7H6#g7dSf.AfaTJ&3D4@+NH,[LedA1XJ5\4R,R.F7U
Q/)(+OIA]g)39bOD(f&ff>Hc87Q-\4/CW_>QK1aYV7[T#cdZ@\<NUG=;(8/S2C?8
/4cSbK4;[6fW0d[0<LG]ZRVXKJBSRZ9f5;<8A[ZXQF@aB&<;Z;>0P61:\BdI##2+
TcBB5CMd?:ZCUdBE_;b\@3W4:4C&F(gBP\=3?bF<[S6.dT](,JU6:fP9NH?d9/?;
/2@1<TbbKeIQ51::;X/fIH\Z0eGNP[6bb\)06J@(4B[S(a+@81/(@66e@A/beG-W
)T>+M7V0,2CN&PQO7WG)Z>eN8+H)UJ4BeC09D8ObB)5P64EWBNbdF=4^FC1=;=E(
]d3;C_.Zd\H?=J/T&7Q06a+fVE>_=>-F>P<EW,]^QX^I-GWbR_Da7(3[?QG40g)^
;U;^^b)^?:V9g8X^G&d4PdVb>S/P6XdUAQS=Y45]<5Ge<+C([P@\aM05O;_b<O4R
EQ_PIH,I?@<OMM\a4EC1ag70JU-<GY,cDT8D)<4@UMO6bE\gcTdQ)B-S@XAB7],I
V#Qb?@Kg;GMC06.EGC9L#2HW/9I)N+P_8=HQ-WCgP)B)DZW0QcQ&dT>c^X09:BPB
A>0@SFNWW\>Zd.X4LB7]YOZG+H5#P^4<-_:HH+#ZFCK#>V6]7K3]:F3F7R4X)6N3
g6&/g8VCLWG,>Y+ML/8;.]#ARc?Z+>&a6NdD#P;dJ7=Q(TPaU>7/d8]>B;&^FT/g
\2MC9P:I95#O>(eO<Nacgb7[b)>YcA?I0QNOZY1dD6AB:F6]=IcQVA(gSf\/cW,A
cGYMLJOTa(:@UfZ6G34W1/A<d\6VD2,a22P;f]1F#)1bW[+C0a<.a.OEf[c+WDIW
Y&1Z;O]T?,./4SQ/^Q(1CAf.G-EDCV/B:AV-L597=#Q80)>,=[eP8I2,U_+?G3&0
^O(VJDB1L;UccAaTO#9TeB/M=2/gQZP-=8I=<Y=?TUQCFYb>B,J(.)33TaDJ0B9)
(.V>dSHO\V9]IdIV9=VN@3X2a>fZf,@Y2J9c>RJ_)GKRKLSNee[L=Y@GT4R1>#0S
9NP;[5_3M0BO+b\/Q755?L+GL8cea^GSE;0g8#ESP/2Cfd@Y,QO8b+^Y#,_;^P0b
<aEUde3I;gVLVK_NfO&fCN36\U1ZPR/@A=ReFgg0fSa2OD]FG[@,=a+?AB?AWNbI
X3EX+4X)C=E=d<B_<AZOGa3.^T,2O+Q<0##LE5TQ1&Ag_:6BDSX96-MBU;,]??a_
]R5e/Y;cM)2FE<F>Af6O4a0Gg(;28D&=]3=6UA3U5RdSg\>^-a_)4W_T<T493&8-
fcA6^d^^;a0Y]eIK_;HU=DUa^(74bSgR;V+JB]Fd4d=CebgLP?(BR@8][)]S6O</
Leb<gAMZCP3>?>L(Fb[E;>+Y+NXbDaGQRAW=FdR[BE2DXJ?8#L)Q.RQH_EN0c&@M
4;6.g_P?J4GB5HU-?@Cc<Q8,E)-_cM#GWg.[6F+HPC-I7eAUQ\XYDbX@<S1,?K0D
ET@-,V>9IMM57\#W=8]d><^_7_0-]^.^W-3IHE5#JGa8;QfI4LB5^4cF[EGUXZN]
VaRF-L>V.B-Y(X<d:IbJ;]ZMY4FN[dW-BW6R1)P(LO5DU]BMY)7=1[]3U.[KREe_
aCb&TdX8b08d=?Q\1L>P:BL79JJW0/SGXWQEE_c-^\#8(/Z(V8I(XSbQNI-T0SO,
_&/>4dAC.:MZ^+EL)9Y\-Y(b#&X+b7<WQ.9I.0/][+B@F<>57)aCAD^QCLB0+Ua9
H(G4c1Z0OKHT-_9dJU4AfU,FeRH13Q[@IKC#\\89\XTNJ(J>W@D^R/E^ge^X-=&G
]<YIYTa1.Q5;2EW#F25DICRV2J.D/8RB&J7Y^Rcf8S(3;J?f=1)\4==:e@HBYK,:
1TZ0F:].U#:1@2g5LR7:FY6Z022HaM.bZdWBCSR_VEMKN1_3F9OYLI]GP@6ABJ3D
>I))[LKfLWa8B90C8]RZCLWVVU0^S1CU4)M@?4#CWA/?M5Y8&):3.1I[dD^A:&U8
ZPg;<F8V9a&OY1PR8A]393KA#BB:gVU\MK<+&&bF^-SG-53gGf<ID+[PT>L\B;GN
SX;U>L&#6/^5Q_+bdM3O]#X0PSV15g0UMgYdH=W=a^3]E=GW5FdU4N)K6GE?VU3,
e^4RfCV2BN^/;&=BfWFJT9Q>b3RDg57^@,7eEI\AEP.FFU6b5+@[Y0d5Q;f8H,W<
Veg<YeJ.QOC)[BOMK2FYbH+,-VWcKP#]9_<3fXDK32@_6T[@&B;dadOYTAg,D>4V
@1D;9b&cg?@<>U(O1\7GN5]bX@7_Q94(9TIGc>YL]Be.O-Y9<4R0:1GSX3QG^(_A
:+<PKWZgcHHM3AF#f/^S2YG)F;VJ<SO0c88W+J\Pc#JX@]D#,D6BT1C6U(+aFHGU
-BdZ\I;He)(FHHYQE#[[JZ=8e-&Z1?J^ZZ1MI^e;,-XbJ0895);TJW4aEQ@Y4M,L
7KUa1,8MH,87]cO=1@PFd#O_2F0^K9Ya6]g>H)&e>R16:ZA_.GX;_)/\5E9IfeP0
ML+)1P(4NM2DHY1+eaN6T>fQMZX5LRNf9Y6V[A?db]2HeH[(]EAfSV[cHL@]da<<
I3YMaI3-?/Na4TD\A(;Q\^ecUV^GU5YeD=1CQ&5V:b-dD:T3OAJ8:e>RE)aADH_^
O\Je(;S(9Q7I(OeU+T^3LX=.33.aX059V:0T#T3?De.-=0g&JBUWSLc=Nd6dY#28
<GM)bZA2)<Y2:7.=.W03-gAYK->87GM4C,O<P9DV/66Be;_(SM/KRL>SU@,61EFV
6Tb]EA;L<O-6=G:FNSPaF,:cfW;Nf4H2U-<3ER+K2<XQR0+S?Faf(N+V8ga1ff#U
bA0H:96F:]NIVG#_ecV>W74XIU9A2P^d:b<Ue>\e?9DA90]9XV&faN52cf&CQ@4b
J\c_Z.E#2;g_b?R_8V2/W1.=96WdZg]]M&VHNW9S7YTI8[YY[@(UDRR7De,b1Z_Y
T0^W7E7/YGBbA^D#=B[6f57/8J//CM&(0HaYO:-[Z8^MF[Vg(0QQ<:M(F;Q/EVd-
(;2Y?:7f3W@gV9;a1(QS5f]5IPU,VK?8\7+N-ePM)T84OWQ/F=Lg45#fEVfM.95A
]VCR+g[cJ^^[g:^-27PSH3;L-MVGWBWCIG9d@DVdYH_9)MgOKIWKG9J]T^1b@4f+
Rg/f^\6e?.3\DVS@YSAL4Q]H&6eS-=>@4;JP99+DAb<W94EXHXRa/9G_RA9-Qb2[
;bNfW.HZK8c=X.]?Z7L;_1VD,/86P2dfZ7Z=A5Z)Z:b3Ue]:H#g=F32XW:RPb:\.
\Re0-,BHE;5e8EddR4,Q1]]^><U.?a/?VKdHPOLTQ1KRA:KZ#[-948XJ:JBBP)>S
#FKSZZ@WI2G1C-NfgV^OUT2UBeMC86d.CdD):=20d3.5VKD^a7W5Z6TWVTNWM.&\
8-&I@Ya1:;7g2)3)>)[T3D-8QE4c002/@)&B8>R?1[+WZ=NU-=,bAC5TWIVRKa,F
ELE-3^+,..Z8TBHD;U0IS0TZ;e8F_BW7N.f4[QCFKX\;F+N1(aCQL+=B.#Qe[fc@
_X_f3bC1KRE-5B2+QD@S^Q)-U[,?C.9#LO[EXgO]8.HC1CdF=CE08Y4>Sgd,+=GH
F<_U#G^ec1ZTBf6NHQdXI#Y_Y^1IEG1B5VEX@<+>AQa<^H6_BYI;/^<5F4WLKeH]
>BNL18(N#5#O3Gc4?#06?X0[R@aZ6VKI1BGK-EcAHNX^/>WAK[61RZ#UN=ICY72Y
d#E-03+dUdaJKV(8#>Da.]feU(Z@IDL5YRRX[gE\^RZ51//UQR)C[b)8gKR][1//
^C7>JNBE&GgE>X5:B657IX0ATJD8T>\5OT13d/.0Y,V/cf=XYbCR;[WUVNYI09L.
#49TELg,gR7FQ7WC.ZG819+ZDU8Z>:T7Dd.DIBa1Yb;@c@LgW#d>RX0a5,XKAXUa
1][?4DaLHI9W;D?QIWTNfeUgKPTG?cAK(R&2B:1847Ma7N=Q#fbb)-,[X\6LK1Yg
()_W,]<6\88>bBE_C<7bVN_T:[>CVe]+G4892Ab?X7b5LJMdN800[bTaTKI1F&US
??,56\-QFYfVH4TFA.4+PN^H^dS=U?/O&WRI7;7.O,C+(9:[2_XS3IK6TM\QN@HN
\?G]=4N4&]d1C_\^-Bef,--HK3agXVLfV_NV0]2-e\_W.fbAV[6&DI.^X2<LMgbe
H-H;Rg&YY1eA4^agg?HO=/=/Bf5+AV\[P@UR[T:4]EV?>+9PO7YL+G-_7G>?)S)E
TEZU3cd>N7<X:VZ>=VH<a+aA@W&2BS,JH5[Ca1#+-G=Y3L&IB_-<2WLV05e(;B;[
D5)#Lg]9aN0HEGYb6EKC1_c4^ILIdN8b[G>6JNPP<HOI7J91N,EJ5+:F1^5J?M+.
OFPa.N/cZ/MN]dX@(QZ-BRY/,S4?fRd]+Ua=Z\5D&P/Xf6-f7WOWB^gUH1+(UWV1
[?D//Y[A4Yf4HI]a49\Q/dc^QK6PG?>SG+_S:_+R\B]#UQ1(RM>]\M(75Cf=>/P@
Z6/[RF/JGSc11\/4f:c?cd)6DVOOZZ/VZd?c,6@KEX>XdNG2,UG2#=:3Tc]:5URT
E();S\3JB?/LIf[G=A3CR=>?,eZ5AbT=D]LKB4>?Ef.1>9(Qf]L#(QA\]5c^9QNS
@V48-21_3O[NS0+14__&(CM#K;2,J<d>O:HJ>C0FGg3?IF^E^\:&353-Q2)(8d8@
b3/c6XH-MGDCG]TJ1GI:^.M725UNG=H#(Uc)L]&EQUGE3Y4\GTS;d7-ITQ#>dK[X
N.,8T.Ga@I5GfR1^MW&<4BZN1aO7.,ZS];1UGU=M76#CVea@XgTcAAN5)IdU+N[K
OJ0P+N1?f8URXCEP,1/<.B0F@M+PP_Lb:aDCJ7V3N7dCE9CNbEVB-UR-:;^?g<1/
X^ZfBE?\<KWZ2+^#4\(?+8WPg;2^.Kd5S=;MPY12f;\+/N==C=:a]7#8[/I?/Wf5
QK\64Pf&8J2fI<g/&U(?M]aSBgL/>UQc1[dR3#P1Y[>O8f0S)7][Lg2II.4d#4+_
<O5J;X=>GXZQ(1d(CF;W\17Q=gM7N,:-a+\&NG09a;8a14<C].de>_O,3X7?4E=:
UJ1RbeBXSg(cd_/I8TKWS-&<CPN_6<]&gYE[X1KBNT_Dc>C[;c+S7AM\;>LII0X_
Q;M([&dSBf-;NX/CN_P<\=P]g2Af70H@M2#L0Z&3d:QK]:D4\S@,g15)3KSUHadP
:,BfUEBK(f2W)27ANX:9\Y/N(2P5T_c9e9UGC2]8D8^?OGeZeOe:Yg.#:2?gQ>_\
<KbZ@4:RYb?9&1&D_]MS]P,1QS7/b&N6&:383B:\PgAd[(MbO#K[b=Y_UYK_gM(;
aUCH<RE>R9[;8>)KC/XOQ_73]Y+52;+54:<Q-WTW@Abg.,I@RAUWH&U/3;KI][ZU
a[&@+cMQ+5@dS]#GUF:fE6(G#FBZ#JMNeI8a<97Wfb(O6:YRWC2Wad.@;Xg6-5@/
4/0?F_@:NEP9,1K9((KA>7C0,NA9RWVdcBTJ609\gLfQ[(eT^[G#CNX8G9Of9T^c
/U-c)U8bgNP46P[-FLE\06;Pg_3\AT=M,P^:2Z/=gc0H0(a:MMSdO)^ZfQYXOOJH
P,fe#5gSWBe#6ACVg#8TEEa859HPcO)4:OL\&+AOfZ&1a^P\TR?2ED@K;cO+SHSD
M[BLLXFS+fTg\d<=RdKLWM4f/BN/<+_dBYZ&AMOD0?^V-F@/.UZC672)[_PW0DM5
2fbe-X79Ua:bGSbJZ.&O<G;4-0[S@CD^6/;)6D7\1eW-F+]S@>)L#W.Q8bIE\3\;
<9cR#c^TZSHJK7fU7)[BS.-QD?#R-;gJBC0N-V2,]3M,A1JOLVV&Pb\Jd;C1gIBU
7RaKg8a\Ve^549W0]1?UIg)J.J4d2=EVU(+E4JDb_Og381^,K94T+K?Sf[DcDef.
EC6A:UW;KIMRJMS>d?EV+7I<_K=((]cGMZ8J0Z.(b.cQ;B?J_W83<B+V)FA^_/LC
8V=c>[FJZP[19GJQY^VOWBH5U\VV@D;;GV[A_dbKa>EHe8^X8DRB.<WL\QRT:-R&
dfB.X#C]PRX>[1;:>QVK]43K[[ABIAfI;^7:OZ^-1?DRAECN?ROEOSA,EN>Z,O.c
74I^&a?I&dOfW\eH/OW<;^5[:<A[WXO(gL,X\gbY]I<]3<^8,V5&_UVHTPHbf>eC
7/5fTKZ)FHB6\1E@UK(T6J;a)DGg=]Cb_ZY@49L@X/XOO,D1RH:\X=RNBOfN#5-T
J+bTLJ(Q.5\5_N8E:FAG6W,+g&3\04E#.K_HB+G,RA.?(KD=f<9)B:-AT?6CRffJ
LGSRYgAO.ZNOWU=:_LgBJ+<N#;CaaS]52L;b]]]<Ve;O@2V;:H+]F8Ig7bEKTL#[
dN8#ZHA9A:AWSFc8P);B2>9P6\GUMa:E7U@QI4E7:E-EEC5V\;B[We+069E\VY>,
C;LT?W:R=<[70cC4HfI91D_MF&=4;3>&^3<+(C-cU,H6X:(&].?>M=gW3cHA[]E@
G99/WF-:>e2@HRL:+.L-W:]B6)TPDT:/O:\@:=OD7\1N3^(_]R/@[(OE:V6.0W0=
Sg7YA0_#f(8&S@+.4C/SAb)47>^7:f3?&JO8f#NBP)+aMSXM\&^\g,gI2P@NZ[^Y
DJe\6WBc-67afM>A==,1\JQ3b=]d]dMX7Bc#M+=HU?4/PY;6F_J6R-G9P+eg>^<S
Y9[fCH,A9MSUMWa7K?/JP_6F(<7SRYL+C858<#)@^QDI3\1db(TE:/OA&B._6>8Y
O.OAaEGf1Y<\&A)Y8)^)#O8gB&?\:=3.A1(NJaAR[0.=C99SF+H7E7+FEQ7T=<CP
-AN-^8?LC^L<HHH=EI^ILY5:A2AXVc9=I.EW>_ID,^e>]L&GD_^(;b@:TFI]Q/:7
O>5RLa][G_^:Vff.=#W#K<f_+7;8AQd.K(MF_:R.QD#4ZK&>_A25gI@PBR/OeFW?
Z@WWB8U6(E[a._V-bB[O8E8V(c@\O\&GR[356C&O2K3ZV&Z_?+O=7#3)Q-&1&c=7
0Fg0M:#Z^4CJ.:N66S,)#6[M[NbBA>Z37gc3aNH2T;U+?\2>P>PRgOQHgZ0f/P^5
:bCcBKVd>CN(>X#-RHJ+THF7Hf--AAO#MbL2+)45cI5JJ#g/afd63?WQD=.VEOC<
>[I9R4NJ<-LXO4JAME6(G&<f5NVU6\2\85^[KH<VT)[X0ZeRd5=@VMAI3S\WOUeS
?807_MG+f9=I<cVB(6;bL-QP@9[Y=?E_YOGaf\)TH[ZK8@QgX8L:9FZ<E\K=E?VK
R^O7AOb)MFaNH8QW#UL1TDF70J6W1](U]_;);^S2SV_dIY8,F?b(DTG:J@@EN(T0
],X3dg^E/@^7:]^&;)IPaGTM/NES4aQL5[^TaO(4Y3.6ag8EcQ@6_XP92)d8d@Wd
UJ[E>fX>0;e\<R01.<GL:]L_d8@_VVYBMHPKH#+^>MYU,7__fcTXc@Z>U8H.J9DB
F<@56/G9ZRc]H0;GWD_AC+PH-JQ186(X,HG[>--1LUIN@;gI@;S[;BM?.BV6USb=
eL1<UVCPHV_C7_4NONXFEFXU6T@/-967<FS]cSc)D5e7BJg[(bNfg7FUe/LC(b3?
A7;<U&MdT-T[OgTQ@;Nf/874UHY:06-_:aY5V0)+,@HP2/LIPLVEFGM3,K^:B=?<
+XGDXVAJc?,WCYITfVacaBI9<CA70&TGCZ_bI4@+,12VWWH0X6B0Nc(:YT4.UBAf
Z5P6YYNU+-[+E-5>J[e35T],L_dKZ,H#R9=9M10@9QY.KZ\CeTL@LI,Tbb&YBNKX
1Y):(J9a_S-U+-T5cc]^1>IgD79[T2_VRI3W0MJ#Sg6[FgAR#:E)URM?=5MBHg],
7ULg8>1>.DZ3f>-48c0;PUWROVZAN-14;AIX5YCG1]>#(7@5&6/;=V7<_BR\g<Q0
NR0^?aXcU1dJMS?DSe17APVA\T]Xb5G9[W/?H1e._3G4M,F20N.LGfT@Q@H1c\_:
1D[@;S0Z<PY>YQUXT)Y7?OD3Tg(09J4W:;X[:G[aV?S56/;:A+)CUaI4DGKPD(D^
eG;I9>aY&RN,M6FFMKLNZPU5)1Jf8#P&Z>[+O/([.0OV^5F-cCGZ2Z[G&C+_-fJF
T7=;8^(2#&N.)DG_NL8PMb2Z1C-c&U-RV7[3-EFPI@+HR:\_[,]8ETcZ:+]N)cRL
N</.OLW8<L@WO)ZFU/DfK^-\7+fG)GE^E9HR3-GFUPQANCICH;K<E)J[4(e.^P6\
N[fU];R\c?\fc#4#WFRdKHN,MT1SDg\2T9U_G?6SZ9^]:(-DWe1?_V\\NN]7>+IE
ESL]I4IV?-M2]L7eH5SaGTUQQS(J_^7FJaG7=e<@#d[&#dY]HL5GC\R9Z+&6<JS3
<3d.7?C,#WR^OO+TdSB#/@&=K.66LV\G>Y:QL[XK7;59<ZJL?-(OHLP-+N,,\FB3
/MVCaYX4K-?bZ#UeBYLF._XG)+EQ._UL_#\WTM+993PX^4-Cf))-_2AA\8\O,IQA
XdGc2<58B0K^c^K.UdI3N7gNYeU,4b=:2/RacBM.Hg]_C]];QX33V/2f4O=6#V)Y
QX6_XeJ1:V(,065#LEFCJASa^eL?34^P6cM70F6A=(b2a6S.0e[aKV.V(>2e79@P
>=:TS>@5d8c963N^&.c?d<fc=I]O&>aO,3Oca_gC??e<(+QK\_5E5aO)VS<J_8J&
-TI&/]I)T2]<X./#<HOQ&1CS04eMHT7\eg.)KLS.#6U4/0G021:0aA#XPb=S=D0,
gKP54&#Y/R+00ZR+YAL4YV4=]6<?HZ561>+DJDN8Z3-SX1^@\2W86Lb5#b;HP8^)
?(Mb.KT.>P([KY+ZYHY.71M>D]<>CK@;9NI_3.f)P0XU>PM&/=TV72#CJ[3?gJg,
I+G0@U.C?E<&f4ADX(NTP0EFIc)]g[BWCWgCJAKEBU&GFTNcU]]bV^=#^<<:39bJ
eT)ZO6<eJ^U_=Yc>?+=Q[IA7@O5-0ccV3DGKgI)Y22[RP,1PIT\VI[MSO1A^Pa]]
ad-NDgNddbWN30H_NM2FaaCf:_J;A?>)]X/57NX,@TbdK.X3WN[X0&K/OGS9+X0G
ffV7BL&c3=V(N_,X^B\VA0NJCSXf2\TNbc4ECK>E&[8XP)(>3V;71>M39U</TB_7
eVd2cJ2<Tc?I</cBd#0YM0K5aE;EZ3)^e)VC[Z&#Wg5=N.X?(cUWgcbH(L^.(O+A
B(b(+OVWUUf1:K>NU^4)M2BUbTST9HE:7ZD[RF_bA?T5E>W_S^U<46Ub[eF(OIZ5
gKSESb?R;bHLK#\91cUC0.6I-XQ6d3];+R8eZTAQ,YVR^LL4gc[\7>>4QP)3U2YL
4(8f,d/KE]4_I2(8X\ddK95fY(XU;+Z7L4>bMPe8L>T,g/_4&Le5FJ[@/Y_WM46F
+B1ed:1eT(.9,gcC1Y<D=>F3M069R,De)(fdGRE6(#Z0#@==S4=d3.gNNbZH4@U:
66_b\R[P64S?B6]A7QVUN4\R]KN5O1gZKP[H.HV&g=X@3Z5N,OZGWAgaafI[EY?=
9H&T#[>0BB=X6e#4:bN;LI5IS]>?]66^TZZHWUG/9G3;IL8gVdMdG8BE[ab[M30?
WTaF=YW,=Y6>@gVBc:ED^04ZafdVR-S#Gfb9N,L,GROG<ZJ(ERW80=F9YC<c-.J4
KQ=0KbU)\&&)bMa5-?=3OKEMHc\e_#\Ec&bf(?A0]F33TY4)XD?LAd_RZ\K53bAf
[0O]]g<R.:8G8A><GS5&T_1:YW&6C_#6OedCa]-QUcY4&:-^FA=Q:G>(CFNRFN\C
Q>>?6(1/fSWIcYfKdCIQFb+4B,-eM=OXU=6+?=\R3K=;b)_I1Vd@,2[dIC/:ICN>
>LS\d;+[+Q4)Y_IGLAJKV[ZLWT3aa&/Tc(e]G]b5\]3TQTWSA;WUE@5[D/(c&7XQ
O2CK9N,MaQ?cF9cT:>-A0GGfM/&C(A?#45_HVJSCPZ3PL<7\<@H__/?FI31e]9S(
VCc0+S2_M,#>0N?Gb>\=WI,][_T)2[:QW&(,?LOa@Y>]0D0dSY=40UTeZB&g?8YY
a[Y?L-V,USKG&8b98bZ9H>.[+g9?.dE_5\[bA;b4[e4/MW:&>J^04+:OE6G/Z^UQ
DBWS8#:;)553EGSX64+]<XgJd&)Mcf^9PI&e&HVBM-[_5cMTF=J&R[,2X[bcL<-1
,+@[1=Gf9DDcd^VA^D^Y[,CO;Ua#Q-/UcS,R&.LKc91.cA+@e23d:A1B3g1[F)+)
<B2A<Of3<B=KAEV,_d[aQ(/eP61A90U07gT7Z7\3/&L7@XPI4F;EQC;b7:4c).+-
/.N/.6WK&K7930=H7>)O2ce-G/07O<<5(K3S\Yc@TWV_:F]C/6,A_T3D0bdQMa?Q
A1\YVW:1gC,NIL4e<R.^a+Z@L;a0ADb-6e:M4P,.WYB,J;f[&=VS@a2fJe,_QVH=
P+=cKJLM4R)M/f2gOJ?DMO+cFbX)GUH?#Tb8Y\4-dK8eUd\4DCZDY]S6aK1IDeJP
L\L.<3;^1g_YH:JS1cDYRTaBV-f<GUM&<08-&B+T^48)(VGGGV18OHc8UQeF_F.J
_\R,5FDFJ.a=EBT^O?5=+LTK5?L1V6I#.6UMM9I50)S^&g3fIL2gEC(fa-.J1KYH
fQ:F6<>LLMHFCAU7[R=-LgF#Kd?TR+.Q=I1gL(<.-CEH4A3:&WOCf[8JCJ(ZOf3=
2_+JN0_U()0ZNT;(e5cJBG\SHE\6DD6-a8gQ\\>U.E&+7_Le5-;[I@(<N\Y9c[OE
WP?BA^1V(>A:bL,/+?HdGO>\fd0bO]=;PFWG2a^LXHNTEV-?d?Yg<O94e?U<44)b
&6_3]:[JaARM^LSb>?9<g/#(=<2XJ9]7<DXgS^S_<BQUSf-IdC)JTeRTS43f,J]Q
GfNZ884(6:5:GS38XEN+>-LAU#Q,Z&0?[Mc08[7;LN]e:_G8/U(&7d]b7_89.J&L
/N+e7OMT5,-/K#P];Z@EW-\Db@(J.-9?0]b41WJHgW.Gge8;(IIL^_3\cQ?cKcSM
FGRM]LV6ADCBc0bJ-6HKf^F4TZ+0@[6F_3JDBAW[2HZRMgF8R8/cP88H:7=7]^HR
AS5cO7)3@];B@\=d&GN:BF0FMTA>W,&Ibb;+O98&@eUSK[\O.^PV\+.WL=7g[^1&
7TL6IfK-P.FK0HLB6&RZEWL_aWC0LXK9.,g6S/;<?ag+(3;Z]OB:-IR9J4bE+5PZ
IHR_D#-B-8./WW=2,1MYW^J(25;W#6cF4GKK[_3\<(edXK)V6g\I])c3c&#OIY@c
PdGdX^8E@RN0_-F)1V@GbO0B\I_G8,IB/bY\:23=PQA0\.X0L.+Y6bNE=I^:+&I.
4B6ZgZc&.JcJFVG;e9CXJX<0>_,@#X1M#8/HK;)^G53RDd=0819:26QdOTR)-Q4S
?#]H9&c1]N[&Pc+(37\CaX95(Xc,KNEcE/U\\M81;EPYNN[Y^KY8O3).0X>8XVKV
I0M-bac\2Q@[2)C?+0f)1V?,H];9J6Z\Y4BV[(4Y.(O+[;>cXT-7)9PL0R__;+XW
;I&]1.PfXb[6&0GDgD]Z8>Le@=,cC-RONW/cD[6V7eK:[-d/Lb=-Y(N<H_V[KaFC
DgTKCf\.POD<3+<)GC]QL>/Z&J^_DgF9M:GXf?9?LZa(D8UR1D:cCBG87FL3P7?8
I2g@:S8aagI2fAKYUX3(a+d7L-2:D.^JI-]_MDAR9\Y@3_L7;P;;D9KS=,-;8RJU
?_\5eHWaLc.eM/XA4E5GIHV]=C6QS_Ye^I&E.YOOLG[>E87P6Uf.E?N5D\K5,=Ie
;^JcSB+BD2:YF^@A,&&X:fAQ)E>N?)E8&ZAE,.+/=H;<9dI^9dE\0T^bL6_QW3d;
6cS@6Pd9>FWZ/SUTQPW??>YBW=FE3<g(FP8O<8)&d?852@[VN?ADAZA@R8ebUa.<
1H?DYdFd3Ka>\?T]bG+73IS^W^PF6,.f2Fc_)gMQ[-6e9GQ.\XaRF/F,KbRH8.E\
[NKPGc<RZLA+J5d\XFJEM)\6e)WDe^MMPFAFbK(>aPX<WKO41FWB#\/:7VWU#5+?
@1QSE.M+UC0F1Q8F2WPMfbRJSA-VN4]+6/41E3.^?5.\-&S6FHI([W2F0.D31g/K
^1L2PQ\cX>^4VB/b_^62>;TQ>M)B(S&RMI(QQ(717A-7W>-OA.?7-J>):;\&=bMR
OP7gL/a#_V+C8IIeFAXTUOI/&Q-M1O##7K?(J\>E6IH23(G7?2I9J>P4V26F_Q4W
C0_>d2^18g;B\HX]A8O(<bbHPc5bU<C^DA\X43-#R;;bN;/_S.UAIMQJE9T2WZNL
<;@K--A&f43(+7:b&52L;3U(P<<,ZNDAARFdHJ[?G4-0I/K]0Pd<1@&X]e7Tf&&<
KfP@gdE:^]?U=[4;9_&G2WMc:+.,9N]ZNd,0.aTFL2/,5g):=97JJ@#1g22dde/_
<LfQRGc1UcU;dE=ASK\;=Re9b2@aW\4;K)<F+CJH<.?^0+[HG)56#5]Xad>..0,>
Pd-a.;6DN<O([#RT]7P,-:CJJ.J>IXOgKg31CC>.<2[4=+<b[f_Y/W_/QZ>C\aE:
=Q.>>,]:KS&6K/I;1d<GM75dgTLgB]XFK131S6PI(fSgIg_^[0Va.BVbH<3#_#HQ
cLWFVeHK+-VZLg6eU^IE7BK)2.aE<0GcAV[(#=?e&-g4;Q<SV@R(2;^C6EGa/509
\_4d__]cS4FV2+8M8G@IWINQ9?/+QG=TIS3YRH\VMb3bZXLYV/cgdVQ2feFQ/0b5
X.WP<NBMJ7A.S9RVG&,.AWQ#W)C-XS8#PZ\SFe@(<84XbYQd(4e_EYCXf=L#YgA,
3FZ]-RJ8Zff.Z1\Z1><FZA=]dM[gH>0&0X43SO-0c9R6JRYF/B)PgE<ARUES8SA@
F@E]\ce;@F_9DAA1[=X-<KYX#HWJM]1U<G]eI^M=<O>@F]>#HHfO]Ac\ED>P5+JC
IJc6LR78(J<VO&)Y8I::O2/C]cXAeLU?P1O\T44;7,D+A#Z5)4PFB5YcEVgRC3\3
6:4&g071NZ9UFaJSZ0A,;UOgOVT9[bWbN^[BPN=3;\4Y#&K##HP-X-TE.gT:SdfM
AVWeGE7#=]]e[?+R.@R+2N1[]=;7DHgHO7W?aVDQF)]3B[a(ge6(eZaTeO71e)C4
;1;S]c^4X6SdT&[:8&Wf81cMYIRUU[R7d]0L4+J\6@5e9\+N52PPEB&aPN_Ac6V(
SY?^Ee/>b]R)dC,NDXAM\:CcEg:]5;F&0RQ/bZ(BEJ9G5.OFI0UNDeD]V5BNR[]a
7(-#^JfOca[(/&#Wb[=>[Va_JA?<9#1VADIg@)7G.22XHI,a&<c<V@&3PEU3\@[.
C#<-1Z511?V_+@O=VTBaI.=gZ#O)Q5+I3T/\cQWQC:)He2U,<@Xe>[WffJ(U7>D(
1>JL.)(OG^fLI@_B98QE,:3QWKaVLNS,A<Q289Q;8(MT0C^Ife/#cCFeL5J9G7/e
\FI0/V16.B1ODd^UW77eL=SLIdSYNIXCB_++BfcJZ4([A#(bgE=V];g74NA?ePVD
/gA1Lb))2S:V@c#O=f@M1e-b<#e=KbJI4A<BW?=(S4\Qa4M>K=#]7b<Cf\;E-VJR
RKIT4MFYKOOJMY_UQHb_MN#Q8U8N:T29\I#d#;Cc^N^cY7R#9WBaK@dbH@:>AIcb
3+V5>:,QASK0#/ARW5e0IU9C-436FS;2=f])cHJRa6#=@b/2_)&7R=9Bd)V3E6:<
3O54,X4L[_S-Nc#ECQQEfP(:TT,X>_PK\FT.7^MADKP&(5NL:e3>C.Id-A;1c5]F
(UH.?X^.D-KA=-b?;cUb+HdGMcSN?0eYUbV3:?Qb#.gZ9^:4KC2&CB>F@=3R04c-
cPdRIL<1E3&f.M(PZKXN5FY?@#L_5g]5QOf#2E)X>7.G\a[K>]MSPJe4[T5RG_A1
GFFXAZbHUO_])a/G]2QeX6,7-bGa:.S^MeJc,agY>^Ig(H[ZaWH#9CKE\@H:<2A3
J,f(PY0/^@SD60@[f7Z[d>Q<;+TD1bTf4Q<T5]RH+=^A=_H7U-EQ9:[\a2>CTSY?
A3Y7OO?Y,UZgdHTXCX5,ZMTIR;<Z#G\[Abb))bM@g[M_AP9FgB<RJMa^@K97SW3K
E-\ZE8\[eYJXB/XLedLKQ3;^T@L&17)eN?X.aHE1P4b?Ab_AQdQfTfTWB\25:?Ta
JWB(>SD1d:M\D<U[9]HE]9X;@IJdDU&Y4F\?M-Jc<-)O5O,U>+fB/Z,f(2Rff)QP
.:ZVN5FH)62+M2F]eJd>53M2HE@9C_cQC[:IB@):V0.G-46VB&VZ+RfAKHQ<d>4<
ZY3>A=>X9<PB13]FGG73-f<Ec#5W6Y[c@=g@\\ac59fC(9&X;0[B=<fOVSPWG^08
WW_L0C>VgD59VXD.EJPV3,=_H^W:YKbLW2>35ZIU&_DE0E,R(P)6FO?N+PK.=Ba,
S4_J-G:EacEN9:1aT0Z^7A=;VJ\dbOJ=dYEe:)[SDJT)HWAZ==WSSB9USf3W,9A>
ZA2M+<N[_^\R9M->J6(-Pa9.<D#(/+KQBb_T[]I?0QJ=E17ZU[W.C[5bKAc-c0LW
W07/gg^;VX9gTU[4WM<Q.[V\S)X?MS<_(N,G#XA0_M4bL^]CHK?62d4<a_K&LeN6
]NGI^=BWL8HM47gISL>AecO7-IF)Z:eO.g,W]6O<2Z7J;;3&b)XgEeI2;Q:COVY@
fZLKNPHIf.[NH1LKE31\d=P:/g\bL6?e<C\WU,P\OP:N];8@^7Be30S=/CE&UP>4
a-F/Z-3c\^D9Q3R3)0+F8e/K+b#fcBe##4gbPeG1^.96P]a)Gd]_,cd^HT9aYB+Y
^86^[2\Ab07a-BGWJC<;HBZJ4W+[N0;8=T2Og@AP53W[;EPS^0^D?SQBMW/HaZRC
@ZB_QF>RK,L).6S14Ng\&C0E.U@>cR5A97MbV)-,V/eG<4Ja7_03[G#eIQ2b<?QJ
=YD;G/?K7[]G]cA04Xg&R?U/8[e53EYOTg<Z9M\+V-@:B4Tg9(QR,(RfM1B1bV7.
(?>M-W4Z7\Ff+cG_&d0@B_G[Z:FXI]9cdYOQ]^\676IXgSfYGIbYNgfKEb.S_UEQ
&JKI9S<?_6F;?VS3TZJWX4453=+M?]=3-Z,PYX=Q,=]aSALf&C;AO8IDO#:FL?NJ
Df,D&-S,KZ0&>@0<1fS/:H#/^(Xe>^9W#f8)J&,S;S3.X:&^W2@Z8VYb5:@2MBSd
BMQ1Td>1S:bG6#_A2WXc>\N5RFTe.<KB2eR7)FgFCg8IcY535T[&S0Z5XTA-I_M]
G_5P2J3WcOSX;/=\\d5)O.?R;3O8PNF-&^OXb0&G/_1DC):dO?K_FQTWITW:#[-a
AT(<?c843NB8.M64R3^9#6P3?PSN+1-[FBYBI01;(DKY&I,VdLLU7T>b,FG-,d0/
fG0NY?-=\BWJRJ&B7J>7TgO?<W:fG0E=Q];_U\)HWfXQ3@-B2PL=,>\UX0G0L>J5
QB6I^8MU^K:XZ[2g2IIcfJ6H+MKUB,:5#^/O77g4ECX:c;K#^,&abI-X+d23NQfP
a;\JO#Z&AML0@SL#(Sg2_eFcX(c&N,(M9_fIe1b?eXD241@ScTVQeg.=IB/T7:&W
+E8d<-FgBN>PV+c3&;._c],L9Uf\>3b9NJZE_6=UCE7UA)(aI>FOdS9\^//\1(cQ
&H<.,BN8TS9gS3@^H],/[/4<OZ<P&e^fP5dNCNAD8LO=G:CMH4Q:_TN,[8E@G4(3
e\Ea<_b>SX1>b;dd>(W]ag2bKD0G=^TM>/d@3-IaSe(AV)0:3-,^Z>Ug9<2WX1c#
4_T#I8[Qd]K#OF@H/&4R;/WT]<SO[_WX#f>Y4Y;^#eBbQ7G9PS=_>=JGR;X2ML4F
Y5d;A?0-Z3QC_MGV)2_XH89)dE6efZR)A.CBK&]&A1B],-B=[=aO^#[HEXeJXLaU
eQF.YZT-J]).4AKB93WT#g=9/LTa>K-)-7-<\]Pd3&g3?QANT0K-5)eFW7Rc(dT_
<8VRG<f8D#[H=C8Z.9d9IU_YeA:/5YKS3.>#DeT@Q0QS,@P-LY]g-)8/]L;>OPc5
04#_2X(bO+Zg=V4V.<;.S/?9RN8+XgZ3b[Lg[^&,=aBJD08-CT+S5b^=\#^:_<GV
O3[ab2G(LL_4K78?YVN1_c79@JJ2DcL#[CV2)3XI4cc6OSMdQ/HZ#8H38aeDfS)-
R>.PK3=YJK174W1dQ/V=[U+/>KSI8L-P=Nd]<7a4(O#9aUYMNdCEd^1E<V_=W(O8
M1]f8UU8=g65<Oa/X5GMf.F66R]9H:)ZX@JAcZIY4WGR1E_c,,G3V]/fd46d9;Z/
7QWB@[Y84L=[,E4fAdD7O,DB(>Y__N@PN)L60#ZD-d?UJ:ff[gO5BAE4:=?<)NNP
:JESe(7X(\SG)E2T+L6D&OU7;7dW[Iaa:02^d-WeYcU?<bYXLTC0F_L2LdL]C?PG
\ULOQ2=HOSX#U5CKQ,f]aY1Y+Y,1aJ/&/a8^U<AFUSgBX.I&3bJ54Y/)IQ_0\B&(
VF7[^YgV#T,>^+#aVN/);^UYV#Wg60G)e](aO64(_>CXUNVY81NII)=O^NU6)2T=
J67WG)>)4X15,UE/CD]G4]3]/f#?:c+(8UA2D7QB\f(&1?7MS<_YPU.gX,V].=B:
UaFb^0:-ZINH+C8)UBDSNU2>3d^Kc4AVd.H)VbGH)N(C3H(/@0Uc0Edbd2U\D9ZL
QAR]U7[&0)R;/)7cE-bY-^>SDWQ-=(2N?:62=dZeZf:e=O=@E):UCL>P@E]H&(I9
W(Y3D/8_2g3@=G,dQ85+MK@R<PKSDE@/#R-+FX4F&be,5bMX5P\DgV>-L6cXX8bM
Z>BN3H&c)f-35AAf6K3Q/IR1(Q=X@80+P?N[GbRLR][>=aT[.D.dcQ:,c(TT732H
9d-7B54I,UH=Z&)?&9=d\O?SW8B99_]:LI,c5b/?/NH\S,QQW9S:2e80F^c)527I
KI^\8M9?4U\XI2IGD4<J3N0[E69[R/]#a1S#W;WP#+b(XeM:a0LR.0_6Q:9TUL>5
SWL#c&H,F)g:^&E7P.cPIdc;.^aS7YZW/7_#EVZZ6-@\07C6ENO\,g2S1<DW.T4V
N(5\OT)8I3bTPaGR7V\OYP5SdTGNSO3MN]MWM<@@@]?+&N^JQ<9&2gY\(Q9[3=C]
Nc?FEId0JTME3g>],9FDc(&GfS\e.V?]>#(Q_N=IIPCJ8Q#7W)f4(B/T>1JeHg(]
-4M9062J29;Xg2FZ-W[)FPDLW3;[=efbXK,+/EIEbPb=:QEHC+(1K#:C.^IEc<2]
J5V]>FWV]O,LNA]R--AZR[_S/cI&/>GYEPB6<Ib=BSeO_B]F=fF-b++&L@PP5QIT
W8-^M8CB\FCP7YWTb(PU\/8\4YTK1OC:a=]W,5f0ZU,g)GSa.E?F\Z#P&\NNf)EZ
8#NPKR2W8Ug\K[71V-e>:XRK?>XZfAa)/RN.?/#>\?48.G,1T-b-.V-):D:2QC8-
b&f5g,_-dbM8ETCQD3(B[V&b2feTFc+(?H<f)#8,cXaPO^A9,5c:NE3-X)XS+;O,
HPeMZQ@J8U-gY1OMCS1J#17\<Hedc[ag&:aN](1a(FP6;F@,&\D<\eQg[1<9+?b&
6E1.X&,/C_JNa>EZeD1J)\JC/EFIaYKg54g1Ie7Z.;AL.c0\LaIMWW;EXGZ@9WYV
H=[[7HgDS8_=)VWbJVD&dH:0?76)^#6PU0^#bKgIFfaY,SIQM6/1C<W08AeU&100
3&VJWKbDg;GBUHPb#YI5^V_Y=5RY4?Rb:J-Hg+07gf@&Wd,&_dW9R>b?4a@)0]=7
E+ZRDX>/5^C#_ffAY.@W<&C?L^Z.MKY3E#<N(FZg#]M12>eOR?f-7=:Y/24QE[ZI
S#N#cbb#EaTL.H/@0L?>WX9ZLG[EX4&R(QT\R@O_O1T6XHO\:OT[<\:^FaM^PPfg
+D\OaN>,IAaaf@0=97G)1TV9LU6TUFSeUZcV_TaW(?]NOdL8338[VXXV4SQ<.=7E
eM&-#VV7(JHH4P\([L1)13V^7++D87RQf?UdFAe0UZ)(DG0QWU00d-^XTaON-?^<
=8]3BPH-C.2RII+e\dEAV29[-+OKC+Ad]cIA5I+XC.,>D.YP@ML0U8d;H?]23P4G
OK3)O3He]Y_0K1,#KK):fM94JIZ)KH;(@G)Z2-BbC^A/O@)[:b1f>IV&cZH+S>WJ
?f<De)2O^<aeO2d=5;?U9=:8c4N)NE(f8),#Z-R@9T^87_RcEOO1g:fY]VZX#SNQ
.?CDeTeYG-dQLAdggIFWcBM<[?2R79AZ[9@8NYC#WWXPR6EBXO,ZfPIf3JU6aVB5
YP0G.IZDF7N@UE.?K@4WK&66&a:Y@:?=_/&RLWF<U]:UT<QV(0[(90H9=W=C6Z.M
,+O2Z\P/1GPRX<,eS6Y-@BA>^e,QNS\-.(2Z:+=B_X^SA+.7gZ[W(Ge;<>GPYEMC
cW0XB2U]JAM)1XQI).)aLA0G&HZ<S_P6,OJ3K(S;#J#=+39UHaO)?A[FZ[.PUbRZ
-?F5D[I\Gf0^VT[2Dd(O2b-QJ5E0bCTLO,^/G=B\XfEQ]90L^RGT&Y_GUTGgF-)I
Sc]/ER-#.gB;\JO,TDO\gA#->DJBPgVAc-=b-<N49_7,bWV_2)U=9W-DGCX.-LPH
:AFE25P0@Q2DGNaVHI1+^FcfF46Z#T4GVQXGRJ^,WL?\bSD[&B+e>\XAV>d-;93e
gH7S#gX)HcY2_90W;7cLU0\HMFMH+Yf81J-8<ISa5M?d1J,7;Wb<W@f37HTB\_?R
bS./U\AG/F2)_@aW8TWYLN-TF0>CMe3?Sa6B;[c7fO-F1e1:,>@TFe/,_J0E@JM\
=aB/(GbHSO&cY3V49S&HIb&b+Vgg/6>/T_V2F/g(]D<>:P;3=K-^b@5]d:Ef_BB#
3\S530B]3)9agV/AVB[+_SFXcg#_75B/^[D8MV_<?#I93=<X&ZPAd:aG:JM@\/)W
]61VTX,9N&EA]U(adAW1?9-0\FY83BL1F_A\E;6-(G=3X.(S(dLX7,?#L9#6/K,-
d/6E=#)Wa&.7C<VcJdMR<dWMfRR[=@?;I8]T8#,>8M8,S\b)C)P+BWOLW6HJgdG]
3Pf6e<:^[T_=#cOd=P6V)NfH^;&X+E,@548/TB;9;6aK5Y#N25K5bURe,[[(IK]C
R@A_;7(TL@a71,bd00e[cBgBO)JLP5+3dc&.#9>a=(<&PR7@^#_?b>@B7<>2)?M8
;+U^\^C:+I=-@gb\IS+0IK#.b5GGV&(7.],)TADC])ZSEW)\7eF@&&bOCO(JR?.d
>3d;K>_B8D?KQ0Zg:aEX@RLK8aI<bU6#]T/bV_f&<)K6:cTKVKUXb()gT9S#ZM8T
P\(Scb;:+8Y7O_LdUG0/FU:W=;H^90;M(T;OE\gcVKff?I715@R(=Zd.AH3G5]VM
OQ/I[,X+AdF5adX&f\8]3UIWJe1H7K3W>2(K/e=[aMCE1L#Ng(#WHA4=4\X)H=8B
[MKfG/+,2\8MdA^DI0#5^Gb35)9ef-V98]WcPB[EW&^=fI)P7]>OV+8]:B-3)>Q\
ZXNQbPfMI(H-4\TWe/^c=T(Z&DD&M-4g.5@USLZOd(DWZ_ML899;/f\14eSZ2-19
=3?@e1MW@&Gbb?VMKRPV_?##cc?g.+J&=+HDZ<.eZa55/<8E<C@30AI2.IH9Y[.a
=8<@6IDI]([5N2/_MULfgN&4aA/<;8:d#7UEV)ZFZ)S_4Vb7ZV6C/60-WQ[F:<e0
Xa6U?dI74gXb<#=R<=;JgC40g;K/BYZM>f&ZY-:e-68)2fc8aTE>.XV),@FU4EN[
a3eSMgSBNNgfc0c1VWL+9MJ,CLTXHB7JWA27EQJBg74Y>WQAa+L1f^NgGG=4;aTD
R4TY.EJa_\Vf-eD#6P,YQ/T9_RfZGB1S1fG^N(,\B^-QbE#ZP(ARg?bU<4Q1S4YJ
7/_>Z]/.L]^FH27PF=_?#.c<P_K^T)9L;cb06/],P<GU8Ee.@9HXC@P?5_c#62=:
J<FJIZOQS@5Y6W63fHZ]d;QDH(::/Q_>T]&Z,V#cd:BG>,1LbRX6d<+fKa>Y2VB,
F\d(6)a-.GF+W>.NEa6=g#b>,J=D_^PC6;Pb/J947+:ZZ(?(@V=3GE(0C2D8#:S^
JIZ/J(].J1d;eDOL&1N^1&g^U#de.cgEfX+0#Q5aX_YLc;T5eL#7BB^G#3e&,^V6
_GN\=_0Yd:FPA,A,7P0)11<\9d^?G.^YKPL5ac5?/d0R=6\#d_X,1]DN;2=R=IME
#5N,\I&R7P>CK4&(gQCH6N2/SKJ-F\6I2AfTdBOMTF)3T4GJNaL?PNCgMP=;b(+c
CSB:@5K&0&9cJK025B<?DU-0<b&^XOV9^d(2C2g#EZ?4+4C-Q9;MPO3^;0_F5M(M
_^SH@372d^1Z(=ZW,Qa/0<\PgR5JZ,P+X)Tg=T0^c^EOFgZ32a(13f3[P)7.BV3N
;1N7^31173H>[ZAVI0FYK,Q&PKK:e,?Y<ZEC2N2.FZDBgdZ/GCa^4#0BB,Age#XK
V^ZK[I[D08ERGJ(/N2Z[D2I,&)O7A=@Ag0<2=EFT9Y=@E&I4@;P3/d7</[8P1OJ2
UWaf@8&E?APNb;X.P;1CEa</?.J_eNC/&&]573=(<HQJ6RGP3C18dP&bVB<:?fH>
eL>NKG_f#E8a5PN/A-(LVAJaB&3H[&^SJ>@0G7EL&\DH?b@24U[4D9K+^J&7<1AR
E#?<)1F01WY]=eN;SW6@0UK@I:U3W4DEfUCg4?J[K0.a2dQG3A.R/Lfe?(:K3P04
Y<NEXUMK8NcVZ)N3O>-dHM^-#[.^+9S9S(,>FZgCE/CP+U]@9f>\Fd69b_IGSKA\
:A(Lc,YX6NeGe),,E(CMW83;FEBb7CcK>>T@bV>WYBOa\YAf+=X^H.2YcOJ[4?F?
7[]gCf+?9P+#/ZfDcO)6<J0g@J<[+@G0SYJ;\3:(Z]]N\@:)M_bYB70VC<(MS4PW
Z#\=O.1YLNBP4D,K7CM;A1eT80L@>,[E6&(5XPB/6ISE4+1SX5+MI3:TR<Dd>I>(
?0d95K#6K2#TNM]AO9[0.)6UbEDXbCZW+;P+,5\-<fK(DAE_78B6[70&@F0HSe\7
/Qb;?-,KK0D_=#[FeDe#IFX3I-DKWSgTA5UfXCPcCgWM522@#IZ;IL7U9eMB2<B3
.2K+-NSFb3(O&H]C?(_=dOfc<U>U,>XG#N,5Zg2VPTI7IW)C>D:NCEN#ZO0R_4/J
H1eMH-[M6b[CD>aN(4DSPMONUNQa+Y0VPP\c_KUC,C)-O]H6g#&c.L?c9Nc1.E(2
9(7+Q6F)^VS(Q&g;f1Zg6XCMHYeK2,.&[?;UF:MDK7&0D-2fEF^@7(fX^(.gR81_
c?cY9/d53KUHIRLOfHJE\:=-07]DJR7fJ?,\F0^b5_THM0GXZUXI][OLF43Ka.0M
0^M(O_QEPU&H:;Ma)E/QM?[GA7PbB5gLOAEV,LJEY,J8ZPHT;f2/Q;gf9g<0g5)2
fC+<+DPT\M_fT<1&;>@E:?0W)-GOS6eBST(8I8:#;U:e=R?AAC+)TH2a@Q.RJ0#E
c)eU;LFU>EXYQRTAO+X,<IPC-(;7U=1QQGO6C0Kd[S,+3,1CQ&)>eHS.Y^,&\Z_P
B&cdBaG(DJ,[BD?M9?8EA3EDJ3g;VXO1:ZJM:7Y:_DE9+8R4eZNYE#TTN;H&8B5b
@KB1<1N7&F-;]:0&^Nf(=I8fdfH0M^-<-+P:FSbD8gfWSOLB[<T:64(>W;+LW<R+
WLe0>^0=:g7K=NKc/D[LLgOZa@a-e.b607(gP2ZV3NF6fbE65VK^g+1P?M>(5cN2
O.I-TaH3>08GfdIYK,Y2;J3?<_L&UaI4W3)MG&ZRT@@f?JL?QU5(WJ#UR/YS<^1U
?)(/g>UIJ8[RgQ=NKBZA.COEAQ.^)@_DQYbKb1FWW@-HSf+QQ@NaVe[>.LO^P#7W
_.QWS7L@2H\>VD90?ccPEE7:/D7:GM_AJaa\<-WLYD(&2(-N4Pb)82RTbRIJP9bH
WODfN\S4Sd1M-<5_0b:+IJ0ITV65[a;,Y7gIRBE<b&OL+g1O7G]_B5cPPJG&S4U8
=LaK&\^ST6M[5Z8;.7IDHg-JG[U4?:4R)//?TcfObX/[]G,D)8#=F/dHFCU9STHS
(B0OK]a<GT7g&(T3#.>c[+>b,gIR8a@6aW^UXGP-=VPgWZ]fRQaSL],I-V>VHQM&
TQ/Bf)DK)bZd+VM+g:]#OX1[/)8N0gC4>fULNZ&0W(bJg8Ng)-,3c+P8+9J+W-]^
Y&E8<6fIVE5&/KHFaE#TY,(AKV1>c5SJ;f\J?NX2Q;:I]W_]CTc#,P695>2#.Dc:
Q/QOMa0J.(3W#<cZ.7M,Pc6a>#)JSfQ<;<LE^1E3QF?d<X]T3U(K53Gf>DdDJNZY
WH<)X-a79LR4PWJ402OV&PX6DC2.@HE=DR3dD@aZY-PL;d8b,RZ+C=7DF.5-:Q\4
_U-C10UQ7BF,[dbC([[([#QH.X&O-\5YH5[C+cLaJaKPNT3&3?MfR<JK)8DLMSZf
NS6&0c<TA(9X7KZW8(,SUKgV,JA4?A^#B(J6C,Z3FEJ;]UR\ILcSf8(8L9VR,AK1
e_Y[72TLW4IQ)f?D:\S\5gc;NY,G\HS#UC59KVd3,:>4M/geUN77XEVeb=-_W,,X
/<6#eV@9f>^1B;.R-Ga;Oeg]6>J&(HaHb/Na]W-Z0K4]UWB=O[:</W=TH:Q5c0=8
@YF&S(b9=D2O1<2UY:Cc<-aZ(dU16N<42B-.g;?aD)Jg;IA7;&&B/,MQ_[Y^eV@+
U39T2XSU[>0b0+_d9YT314)CR31VBd<PP\X0;D[XGZ+C,#b5+@74BF895E)2/g-X
XTTeIM7/TgB4=cYf>OLU3=2@]C-C;V-5X>+e_CZ0OM^AJ-;YPUO7_O71PEQe:=<e
]Lg6A=6B36)-a:@NcZM>0@/T+R#(?IQI9@be:E,\d;<,PFIGJKcaA]+68R#G5D/N
>T&;2/I((_YT\dPf+CKB)1-U#b]eH^O?K<[6YK0fE3WJF+@T2M_5ZLe1J<HDe-J;
b6d74-#\2],Y,ZT\CSHJ#K4D1K+)(&gQMIDfR8M846EGMHdGWfYP0BREX(2FB:K(
dW[/YQ3^fC3#B@7:M/A2<-SW9aUe;J2EJVLDDS:;PP]#Sd=fM+15&8&V)FcT7:YC
T5CKOM:O&@DcG#d49GJ#WD>dU&0?\;FX?&,7c]?[F<TG5LG^OA/OB8SdbU-Ub3Y6
.QJX_,;1?[He0E4GgfEY-)>,,5d9Cab1?LGX^E,X<CVUFMHY)cW/E]QUOLI<O+\;
>TG.HZPUA8Ka]]XW461<U5,9?-9K?bF^QWM?.LD?-VC_W=fRX:W/TfXY(dg2d,Te
=WP1Cd=WDCH,@62H[V?RZGYU/TbRLf+6HOBGIDKb]\WW(M)[XeX1@2.A)]BbgX3c
HX?+g/#a>5VKW\1f@I4#[/503CLR\H6;TR:RT6H[LY2STO@c&:+LB8AD7+6R=DfA
J.).eO2DB7,2D72<\5ZQKM_K[E5.WD.5a[_3W59L5BKXJ2aaLJY>PO5dZ#d8D>If
)UUTNBA>F17N@PgZ.<V?DGI&:U@<ZXUW=LeT/.We<PHH3:7V+ZdKe=#0>=)WBdg3
2I9S,T?YP62=3<]SY^O>)2EcJB\5IVfB0WQ275L]>)>3UQGL9+ANI+=0[2dB_4_1
7C]fE>B&CU/&66.d#7\f__;D<Vc;QS)@<S@<6=WcBJaLeXSL:g@F&QWO89;Z;Q6S
^Y0)BDJD.N),>>V]P\4,(YP,/AdSX+O2PY3fe_=5YRCG>L?[25:;#/G6G^UgX#/L
:=2XbLC:@H^gJ^3b5#B&[Ve;dYTW;Vb5>aJF45AW^g<#FHNCc-:]&MT@FDf@JN?O
TXS\UeE.HN+3BdYeNI1;H,8d#f_C[#?NM#5_FS26R,J:0TBE:DfaJKd1FI>/N4>E
H3NK0V(/T-CEZ,5OSN==Xa/6;-A(P+O+:>XZb0]_S8fVMdXE&A,RRB3L7ZF983IA
Me2P4aW<Q5-WBS,D85S;&?=+HJJeT+d2O;TYg<Og-;U&-M/\UL.cJCCPH,\L6FMF
/0(P8f;G)dcA+L<R+M(4-;F:OfYPaN5XU^PJ9_N+CVJ;.#[2E<1V27RZOH#8T<(<
-#;A<AVNPIE&TZG8Z].66J@5H(cWK];0Xa:_EaYbJcg9FLBN+Y&=f[bgS&0&W4RJ
#cS,a_EWeV]?HYKJEVB&LPZI6/UU^=OE>HY2L7^(P3\aAI+ZAFdf]eJ)cY<F,O3^
=2:CPM\U[?(;LK,ML]-8J+=OBWSY:7,?T#eX;A(3f2L,NGX0_C<eX5)/O&g7#21X
Z&\(2O#JB<9-f0@3O<#.UcRM-JB[63Y30G+b-:DaXVa@CU=.L@f8QL.W]EUR?OP[
B^DAdPK-#4\^F&4A84^W\LGXe_J2<.EdHB^O=Z=07LbIZ+YL_X<_f.;K8X)A;O#3
YR952_A;B?=XWFWJ>/DF<RNd;d)+&fff^^BIfeKAVXF;XgKb6M35E9g=\DJ?+L<A
U0572_YUa_\?,Udg,@6VL\[L;^^/d^2NTcV>2RHCI_9#3Z3P._:CZ,gHg:._TfcH
>F+0H\Z;<f2R3:De0-eM/;<;F24XaJ2-(D37XdfFKaL)/M>f]\(e1>V@g8LHV+RD
SSHQ(-U8>QIF0V@gg)be,LR&F?]\&36.8f]8.4f:XVW()X\X>f?e<\Z?c1(B5.(I
aJ2YWE4J98Wc9_]H8VN;.-PG2OH^39]LgP=dA8B(Qa&,X@VM;S<F&Y>_D;C@/)N)
ZHQ,,a5B)J^@@B,AfWBA2#NT+GR_A:XfU-WYI,J[F2WAC@RR^bc80)Ufe6B9T&9P
U^6-e5)_6S:LN,c;eZ-8JAQ^b>QP0W-O@&e[\Fce4ObSg;NZQ6a)bFU72^OEc&d@
HRDK))WQZb4<J5X5K:/)AI.3S;7>-=e+:74b8e3TXS:,TLSA=b0?DY0M)ffUa#Y/
4:+)BG3=X&6cA_#W5K#\-a5cQ@Q>JMM+6(VJaVRZd7&JPS,_P5X5X\]g9RB0T6]K
fV8VQ936/3=E4W<=/9PR:G=e<FD9RSg5LU5OU:IS92?Eab([A#0+5LG.L+X8]b&(
]W+ZBga(E2CBQ8f+VFPB\<&5:Jg6X@/aA;G_\-Z<+\Ke>BbC7\f)/KNL9U),F&];
EXQRJ&:UP.YgBdW6-eCc9WOKT&V=Zdb\8UC4YM>L)DFRC_L3\=bMMN5?#[.0Hd8(
YJ\0>^77+M)L:HINFeMa0XY5/6H3cUU(8cJJVc3QA7SR0G2eO:SIAQVdZFOeQ:#)
P__@>=]ba9LZGdMAXQ/W9)ABH^C\MFT/[K_^M#J0SRG_^,;U+8BA:L&[8?R)R<#c
NZd)^6aM(XA^OaKO=AOf0H17TH,_^.PFR7FZYPW]_+[T?EE/Wc4&8NK5;_C4)]^U
F?;:R+8T-N.OBa#)Z;R__HDCUWT(L=&0Me64NTJ?:9N6K4#DfQ&OZ<9<;@Hc1>aV
GPb80_0QAa>3-8?2YE&?W&BHe5(9/BBDC9PA;71<N:DU/R1XaZ\TPAc^/^aC:?5B
,./</)_HSYV/][]fA&I8Wg56&_D-W#gJ.:.&XG2NQ1AgXd4/DDA8C\<.BXPf[10/
<(?ZKZ-bUIW>/O(;d_e8(],f\O^Z-37,<&S#:\9^I>:a_>YJ_1fM=2cfSGM71M8e
Z]BaHOTW@H1V@B\A4;P?T4FQ483Q@TZ6LbI6P2L<9?0:5bCXX4WR,/<,.-W[K\#R
)5-cRUQXb^\U)KXRUX8IP9Aa,)ZTR(^<S>Rc@NG[S<&8G6c=1Z5?.6:>MFD:0H19
<e3S=L.P@3+Z(^Ia5]BC)D,I/Ia@Y<1.ZJ@MT6[#fAOedIV)aS(82#B&@9M9aI:]
e[I-2[aUY(Sa;F.K^:eG^LTNB.H\d?d[W8fKTOT=FSca70H6A3_SL>58-;bDCF@H
6.5WN=f_#RE1N7e92?::a6GXW;5_VCXC/A6)M;D74:)#48;XVgKefA3[YJeEV(_^
]=)YM7&4^;3gEH]Pd@O;-4B16GLWb,G(Y]P7;-15CaOCIP_TCTF2aLe.A891>],P
DbU1_GI<@W:(gW@F@&3]B_K&aH+JB5OI1aP=U)0/&gVHBWYg<fOHKI771KT(.O&@
L5HZ[TgWZ/],9_:_P&5bG_YN_RE:\9&_B.K?@H7FY^e\02X6/QFOWZ@IY5TL.01]
<1-LO<(Uf_(Ua8?0e#,MJ>ZI(^IHL83aMX[XWRQFL=@J)@Xc0Sd1Af-&NaPCA-B3
K:#D9NRSD,Sb)=,7]\]N^N+GJ=R>_B8L08C=)F&JO9O7COfEZedUb\L44PMP6T+N
@dRdC9#E/1XDT69EK+TAK+O3=8,8,T?A33G0b_S,62DTXX705(]OGB[).MYG5.b)
S-]Y#gV-WWUd9U4-3&O?O(be<]7:@cg947dMEWQc>G@7G4E0@ROffJAV+V7@a=,^
6HY=c5JVU0QGKFB^C:VVJ8V#/5X:MYY4F,=cY>:\#)b7B>_-\_IV.C7BK&Z0bc7A
9.835IcCKcYe<)Fe06dD27=I^K?f2YF-./PK+@O^8;gN0I^&4H80WGc;gQe+aIa>
M?MM0[G@U?UKD.YdN.8WdX),IO?>e.9Ha7QBGWOO&7EFU_0G+8_dD\,C4?5eZcQQ
/,dFJ-=/H0:1\M@V8-/AZQbb[-SY8@3)XS>H[DE0?8^\)0b]N)2fAO3fE1,>GUKQ
;#\gN:P5g?)8b^>Y?2:==6K+g=f5YHgT/9AP>Y7MM\+(@8K(#63,9PQG<>RfYSdS
^=-D=ceb_a36-?2\H[ZL/SA;.:GW5SVQ];A9cZ[>3)^/6,^<BQL.6f4]@Z5d+JIM
AId]\]3g528BOO(4C^JaB70LA=b<g[J3;^>P+5.K6UQ0>RdR93C?R)IOgO+Dd+(E
50#Hd4gXPH8#8R>93/@aQ[]]PFVC^75=Xa36eV#d.D>DN2_L@=<+KG/Q)X\-d?0W
\b1(S(O[a&eU:,4XW-:5=b_b>9@/+\_]_Yf-E+.(+[6;@1Wc(YE_#39SBE/FZC?:
7_H_1cYMH=<+_P.OQI(7_:](^2DeY\9W#DbVfRaMM7>.FD\dd^REe?f35?9X71U)
c)@-[I7V6K_:G[((SbH+LJFcTKUaP?^gD_.LE<X5NV<Ff@ZO\I=V0@W5-O0cK:d.
R9_ARIH2ZAE3650&A>GUWARQYd\Ng#aabeVU#c7C2NDYfP.+::T5+TZURI2B=-cV
8b@RgEI)3L6_N-_H89^SMJ5T(>fCD9^4=<_#K1SQ;XgVV7c2R</:D^RU[8NURLY@
?8RX,P^=M8T7aUPf#))4^G1KeYGJ<]D\KL[<<:OR.FY@A>5eGM:K2Sa62)NG9.K/
bTBf835-Q3PVFeC-7)>d^SMCUfO):/>A5NXZ2#bO)FRS1a[L+R#MNb4)^+2WaP(-
:aOT4^5LW\+C)(/WYV\<&N@F+XL\LaI@eULcf[UX/<K,XIHd@dL_8@PHTZ[DQT(S
=NfeWO>[/9C42^FIO>PM5TX(.D_LR,HQU,@P/TPe;60+dUF8(/1f+C=J09M0>UQ.
Rf,:K\,M\CdC:RR>P<7QXRWS/Cc4\_]LQf#ABTF+HB5]Z#M@eCH0[NPX:cDO#]9N
V4^;U.V\:T>-1V2.)SbR.0C1e(.FU-;G>Y@Na=/E<_UcSVYKfgKb<>^Vb0]bC\9\
X+.N^E#DA^X(<^8I(IQ]FI_BQ&@TJ.+b00(W1XCPB,+F@EP_?P+MCSIH;NF6-,B9
/b+MD^W]eKOBaAV@dFQ&.C,;V&0U+9/Y<YJ7/44NWCPR6&cVd(3QPgTGOG#5)If,
XF4^>IL)UM0^b:>_VWQ=Z7=THKObaGcIBJ5RA&(c+XBPg(M)X[2-[6/b-N(KOIbW
=,<5WDOB;@3DX13P7E162A454LJIcM44\+Jb+\J_ag&.76T3[P)?1RDHeA<;F_[B
[64]:JbH8#OC&=H+[JeSRE)^W(Y0^=b-J1.60cWW/ON]d(S4C)?#Yc2:V\XP2d]A
VV1;V2=aA];G(N>(;@0(1SZ+;Y?cC?W.Q>K\Z)3U)H+2758IG^^dJQ^a:.1=f?4c
RUC-Rd)N-7bG2]Q<bV6^-A\ea(7\P<1bZHc_SBYD7O7:G::5.<)/;5dJ8BJNcB>e
^a;<<-EPIIFVXS3N)W\Zd,;@MZA^20M,JZ0e.>06JWJ(c[^Qe:EGX=L<W>SJK\@R
DU,/1XR1\dFL-D=g\f#6C9FfU2ZYE28O6^.PU.DYCC:USSd32P,&(2E+QX]DH?\S
1.3\f,(bJD]?cM>>5P<M/96b8+M#>4g&O@699ZMd_9:_MgV1>FTPAP.7,Y7NB:#4
S,\APaWLBYAgGN.I-VcF-S&RT3XWM(C\#A?HCDS@P/B]:JFMBGa_8U6ZZVUDK63W
=g[DMfV003&UF-++X8RXg>8_=^2TB8?&9FT=[+H&=H1QK3@4ORJPWbM,F)C?#,Lf
?0Z]f_NUd9?bdL#;Gad+ZKISH)=+:5OU)<)D3HP<-\d199Ee.;gN0:_9[/dRG/b)
6H<R0e1B0_a\;:-P<ZQE[A2IWE]-M1?N<;<#:2Y_=ecDDBT4=Jbd\]Y_Q<JQWgKF
^9TE)RBeUHK@]PK[LFI?V;.<FG/L;2UE5E&JRe&6#&?LU=ERH>18^IE#1a6?Ec.8
eR-adNP=-U63]N:(TKGQ&=Pa517-S4d\&UHE,Y+9F#0MSFJTWF5a@+1K69/^1T_/
M^&@fP.J((\I#f_bb]Z4YB)e?b1+Q/)5dZaG=?2dTD?dg[;e#3f,5.L6ITe?6XM@
<9317R#Ea@.U+^I_&966A8bGC^S(BUP,f0C3T<a#N@@UL3e5-QXB-_3=+D#G5UgM
b&#Y&cRM&UTO1]DDb&H?P+,C20FDI?3g&CV:&[@ZAObVJS[6e0MHe+)T/XC,GV@M
VKS^LFKJB/TY&BE,N2gF8e[9W(c,OgO\LdM/dN3^K/QSdXe1[?gg@8bDIY1FeE]T
N6@)+?3gdFHcFdA(9FEf;R1cTFCQLG/S:OE6N25=EBGGQ.2=[UCYN]W?/<,dU,+[
:,^e-6Q+2fO/c=dK.H?<Z+2T4)UB9dOe4IY4QG1X3cQ1<+@HXM\ScBXc8#0/-?S.
NLY9<-4-VBSXWI4@MD12)f9\\Cc,5/[E(^,]3ZAI6VK0Q2\Lf;?:LEbMcT)8Z,UY
:>MH\,bKN.;-@7\g3J:U-GF1f^GePc_:,1]O=1O,PWZ93O,X9d(8IT<PZNS/20,\
;JXaC^>/?O<;^\97efI3Mb,e@RHBRfA<EfPN\f69\Acdd:T#YHX#4LZ,Z&[Ra#,;
/@B(LP\^\D]DYI0BR?X1[N]EH\&;7?=OV1]5)3EPb,D.Y6/Z2VPO[KF>SO>AYe+-
@;\I5;87D&&V.9b6JQQ[4PB\4e1c0+>JZ&YS6T6dRI/;VKY9@+[YPL/>CbIN<;M8
#S:R@-G9WGF><a#CHW[-6)6^3^@/a#02Me95<J#90+REU&J7fF&QYT6L3Y^V]W-(
T58:<4d;F],,2>.F+58KE87.[F+DLXZM3-0C9LFW]3J]<#d#Y)@8ADV>FB0&SY&N
V0^1NZDTD7U0ZF3bB]Z2?0FYd6>2H-GZGS,f4aHZ?&2(7GKe[02:\b:S7S59(=_Z
7EU51NH,)+A65#L92W7223MFSA@4+R/MMRXcW9>A7\>2aHH^QS\4aTNc;]WHA=B=
9c<8U[__TaO9AXeID]9&\eG&HIbVRT:GZ^C>C)A29)#1@I^23M&=A8+1MA2&,Ze:
B?UaZIL3HKM52SS8SEg+J52K-_^6Y)CNU[:5MQE<dH8IP=(T>D[<6I+1LDa.ZBSJ
_HR-e:EO>)Y&I=;A2O^Y]RX/:CeT8Z2a-^;\NJX8M_;7@;_](UG(8McAS/ZYYYe3
_/P=.KIT^VO&.a,&2D9PVK\d4U(P_VMRe]G-S.Z#&9>5L)\R]YB1]C4<;0Y?/UBY
d2DBGV<cA\cCH(NI^g3Sbg#01ZPc^dPYF<QNZ5PT2T/,4X?gHgQd_SBQCWdIT89I
KS@V,BR;]9G.\G8FbKK05J?5]?;OU@UMM^DV+/>eXc^@-L#3O(1G,3b^Z+Q;S8U/
BHTW5\=-](d&g,3_)I])HN#3(aBNf]9L&_K4TRcZD^0)<3Q\.CTbT:)LK-AIV5?#
>C/fB&-d_7<7\3:5V)^RQ3\74D;R9)C+TfTBR3-P;&.ceVKd5WZ/V@>J5b\7ML+:
TaB+B#S.JVG,3JQGZ[cNVYN+TSILD[E^X12&D[>@^g;d],W^1:=7H<CeTOTZ@2<d
,Z(=d/@@aaBgXE43=)gOK/(AWIW\5G1-J&3<4775U6^(SM._V>e2(9YYP2#(>c3(
JUHM19,@;9;g,&XF2\?ga6>R>]8>+Y[F-ZT,c.&GdK,0DIUU]T_I42\MSAc\?G83
)8.CMGR0BV\c4Y^@TGTX]7BXQS_F(;C#-e1bC(ZI^8TX7IH1(1WT&I;G0(PTF(9D
6MQYQ7^+Wc2gd,#+AKC&S>g9d5BDSTM4cZF\)SN4-]S77@PNRLA7Wb417^,5.)a=
QY+?OML;LH;G7[NW-MNQU^4GSVd38;R/Y+^Z;FKYLM@HcYf8fIZB:D#_(a>@UV>F
:cfNf23\?VeN8:Y.b;T9/@;E-/:ICG^H20Fb4X,9:)6F1J[CP_XS/-M>:GNY-A,M
E4Ge2g7)22<g>3L4EaR)>UIgRP+D0fS^ZEEdJ(Y7OS1Q3,gE1;N[B5F<WG&,AZc#
D-2TWeCc1-[UY=Zb^)L+W\I;(6FbF6)gJ:<<.(cP,POY\cU92NSRM/?^3@@9VgG-
d\;c3)X+?.;>\G;3;KH6+/Y0GL0ee<./CX-95#U&(D4cFJC1,7G]-.#DgI2Q9(F9
YCD5-)[UHVa2VD#fcV+-Rb_2,V&fF3&gMD[3JQR6-DE0DJK^>^E,TH9(M2PQ6F(<
LR2WUBJ8C5/ZW\QYK1EO-XM7HMB3)3RLVeJ6H7;1dPJJc2S>KG0>Kgd+dcV#0CaS
VAfF9?Y&C]8G0Gf,B\38Z?@2,MVYg\&Jb\0TLM]:CZ@APfSAa6bD<2-0MA[A9T?f
&?AIV6<VE]e#2D\MW1[HUKRZ76]4-GE1,43f)Z,Y+CL38W@H7GaKG==6\?2=E=8R
b-O&].?71<A<6\e+6-<A&Z\C#IZ5+P-54(@e.+1+Je&J0+7K145<EST(8:0c;4XY
B]Mg:1Y3N7cgKW]C0dQ^XW8P\\]3YXXKTWaLWFATX;\5Gf;SXNQ0ZMJS_()CcW0\
aL<Q9_1g>g097FJcPTgE\&+W5OeSDMERX4e7@]V)+E-W>^=<1#V?#WY]TN.d:FBM
G^dd]D-Gg_R^NR5Z)7E:L#bXMJ(_])A&RBY:,cabPOXeXU-:Z,YRFK2WUG;.GM[c
@#<;GJXFDe=7B+U&3?3@D6J.[X:.@J,@8WecJ,RM]?1)DDP)AF3V@0((8W-,O;Y.
?(?)]Hc3b0334GDXL(;[]SB&UQ24J^eR6#MbDKMNOP4W,3\@ae7fN7fb^?-LK+L0
W:Y2>R3aYIc\WBRe6E3H9(35QLTZHO>gfM/ZDBIfI16GIc/F-;A97?I-K-&>LJc>
Y[8MGNegV0VCQ0?CZ;>.KRP-T97#VQXIe.MJ6>?;,eO)LL^D+#JJ6SS7:^TM.Z4e
P7d?F9e)6P77EAJTJdH5A;.e2.Ya(T;.>GY:8\d84_f^E<d\ZK&,0:IFPc-TKB<&
-PK-W;BN\1Y0gb:Z>.QY(@WL(,JMZO+PJT<50?[bR:K#cH]_O[P210(MJg/UXF5;
b0:<4HR.FF:b^fa]M)3YOG</HLSJG:F>-19;C_#3Q+EG;Z1GV4U/R6_>/\FWXAGS
O\&1<d)W;4WDZ7N:.Y7O_8]3#5WS#d-=<VfW,5_e+O(fG-0<CWMVZ+#P;X=.U6ES
0,-LMT6^G-O_#_LF.A_]GK&)GcDZ.CL&Fc3OZ@gA0Ec20,/>AE]e09]RC?6THLX5
7EM7NIU<f&0-cM5Fg4HZ7Q->TJTDW5-8D=HJd3B0:LcP8BQOYAKS-e\A=YN2)O57
=^3GSQS02.JNc4V4N\-Q+FRRD#2BX)J6.;.OP/SN62F_)83&JU\eZMM4N?GT=6c#
g_U55TWSa.8Y]Z\B0<bG\g\H24-Zf,A?21_e8V&>QcJJ1TZ2BWNH61XDdKd6CQ&]
F9<CK>SE]7UYOD],I8388V:P()XZ7PA8KF,M.AG(5Wb[F;=7WcZUO]d7#NY.0Z:M
f(Cb:IV3)K^,)7HH9:N.,YLM,B/]aZ<@GY7#/LZ<fKB6>6?ICY4ZA8Rb>G+Vg;^U
PP3:];R6(-DHP\..V,PCS?a\-T6<d6#D\e8:/>E.08S]>dNNFgZV6O#a8Aa<I:U9
;)F>[>\HH2aPE^2:)YQ,DPQEF8IE=]@#LPNR;S-568[_YWNAGPg3)db:PH#Jd(Qg
H6EfJ=EK>VF0CFa[93^/a-0<2P<;_5EEb@WbZ(7aTW5^;T-8L/]H#TZIdU.L90N/
OMR9g<0?BVM4dA.[IaGKG4(UM\YG.dbB7b?B8^YCY_2J8f_91AQLQ<3Y&>];6aVA
H@3#-aMR1=4+1M,)^5(=:S8?QF2(J1))G[^K,]eXRUMK=S2c<?BU#4_&>3^GYgYD
dR/RgAc)<a>2gg-fC/If5N6=NEY);;W\9HVE<?8=XgR#IL1a9_H;D?6SQ3F@(1)S
VPc[<P8L-??NE(HL59,(X&-2M@/Y@BRD,]@)Z^ZOV]D2NQ[/JQ@&X+cTF_B7)49^
ZBUfPSI+&-.?\QCEEa^(4RGeDW3@OdU5=7N\?\^BGd(#=HfNW@G7VSYO+8TWG;32
]MC]c2UGDXQS-;6[K-4.3)A-1(TA-d?#GO0MF(NHH^d/SGT^<_R)5]cZ;fQg[?bd
SWBf3ffIM9;ISZN27cFQ>1]H#L.+:-;PU0d)fc+>#1M-=K4MITX70/3RG-AdWTg(
Q\HDS4F<GNXUEMPEe93JXg\&T^6ICd71Y^7_a6OT5cQ9d[P+#?,5QaD<MUadJc-)
D-7YfQGI\0CcO<>E/5]9UP?GG7BI=O]HWOW]2;R?:;)d&?C\GO(TP8:ZOC]dQCC(
VPa.5_&\4,CH+eXNaf2Z=3-?N#OfSJH/eLU0eW]]af\UX<f4A7e@<JZ4=T97Ye?\
ee(08KD8/@Bf<^/-6DC#7SRE95PW17KD-fJ[MXAZ9+4R_]HUAf<,/2]INED\6VN6
(ZF-6+caKLeNFY0B6JHA2V_c6=BPTI@^>X>d[THBLOLRI98PPb\SCcH]5FGNF[+<
U,JSYF+Y^>3HMPVIgZ-#.<5-,fTQTVMGFTPVC\S=]J:L,_X^I1C)5TMaRa]:.V]0
KD7MH,+H=53F[<0X:]BBT+>#;:D@e^W>XN&d(UZ>:ZJ[c;S:?UD6-d,V^[()f&C8
:KXO@\^SW)5>fUH0_P#>6MK..H:BXMF.g7I=:GW4XO<KX_<X?_;Q[f#I<BFf8UGa
#/+;DTd3@WY,4YTQ=f9TP,f,5c2?c=DY.+9CacRK3C2M4&82)^GJMST#S,/TU6KJ
#J/#L1+21.#c#F\^R.-^RV:IKDWN<e\XP,MCa7IR9=Q[M?8F57e#a_0IE_4UEN-a
C@UOc)>f;CU+O4<SO-2^=:fAYQ,8K_WF\/Jg=Y0aTe8K>AH15RJXBQ9XQ<U9-9LD
JB@WXV=&4bcaA_L3?L.F)52LU)1GL@;NI0DaO/FUg(B;NIP@4<f1(5e4BYKDW9+W
IGY.R4F/0/=IVVL@RN;B0-Y]\cD(#1@U<X=LfQ)J<gX?B2PCaXfW,Sb#;:(FP#OT
E)J_;/J73I79#HH?<\;P3_&&@3CfDT.;(8@,La0E6B<eS3/]6)ddeP6-0T5MM__(
FA]Q\WA\Tca>)A0TOdIde(/H7X_gI#/KIc?9?HfL?OXB,9PIWa>CZDg>LGI9>2a)
U[IWF<>8M;=+W@ZESMg(LN/UB.?WNX/9T_L>dQRG^YM&4VG#DFR+\,:V@UCVTNc=
SbIDd0Bc&DYL9-Hg=(cLE=23FGIb#UDJ1GCBHYKY5begFKCA8KG.8#KbI4MSV_KA
@ADeF3[[F7M2.=055^3Q5BOG-^QFVF;U@eGSYQCH\X8-ZU\W)RfI#HN]2O0da-MF
,:=J-&Q6cS.RSI,c4ceJ)C)fGa\>2YB(eE5Q)\e<HMR3)UHN:S2>1K-,2a+3868Z
9L31>>@+R:>YGV)Lb9H>1ce(J[UP@aXBaDMJSO61CEgaAd>4I;=U10BN#C?TR^E=
ObKL?H/;Y_)2F=b.TC8];a+e;9.6+F3\#(/@]X<GEK3L<eS(5V,R6.[SHH(N3b\G
E(0?->SUBVUCdaaIPdH;#-U-_0c@1SMMV53:.0V_A#=@V)Y]TOUdZ=A^?UW=]YeG
[U:913T\3a.RM^DcY[4Z0N3fdR37&TR+M1T0Mc<)Pc:OGZ<bKJ5FAcANGZd(I>,.
V6HPMGga]R;W_NEeEYXL[Q<YQ[&Rb=A\[9OO88^CF01CWD->G;QM2B;>F01VWRV9
CUe#X=W1A70P@=e/-Lda#SMgG#2Q3QM3.cGIK[dMZ8#bD<14L+]?;3.6FJT>QA@/
fY<3Q&3fJ_PX=(5N?6MHAF?E#DS?A5;RTe.H5P:\,fd-0##\6^PRXIO/c933.#[f
8gSS><d1TK5eOAgYd/HdQ=L(EV&M1KYMP]871ZbN=3>MO=P?ZSJ)\J_P@Kf)+1X1
^TR#K(X])92887F0RY43Q[7EC^2T515f,.RHTg^/LLP>?M<,4NR1T).)4Q^JP2J>
=-I_@KY:&eefM=VSdFF>H+[gWf&=6MACE;f>T5TNID:;4D;9Ab,fc#^)IR#<Kde0
b7^Ed[&\+S,E:X9#JVH8NS,5^>TX-3:KG\&Q/FHUG^3&_QMaN[/b(\IK67R,bP7;
b30gN9E)GK;d2UMN;V6-^4>HE[L.FE,]AI<BdCML9:IEbK9=IX(/UHX@0H-cYHQa
e-IXGQHNFE0L_)Ue,H?PL4OHM;(U/?4IX/b169JbV?9#SbD@Y)Z[2>=^@a]aROA)
dD_BCGF5>AAW)YP#Z3.fOK,TKXCB@O[A-J&_cF&dS53gMTNKFLK>XCF,#eHD>1g:
L9ZI0M,-3\JS0W>8)L[/>>@bG@K]+E2<#gc2<HCbc>?815H:KQdU\]Jd-:LULEN7
U0Z;V^\R;g=H#9,<aBe65Q6bWRWY@c:>VL/+A=^__UXaP\d+7c=_7UH(e,(3B/[W
2NLBC;#SX[S-&-<I\U5#_[)\RW#;>?=Z6BH8eN-O,;Q)5=PLf\BeCO]5eCT43H#-
BZ;[9KWI0K3OBcW#d&6aT@#BYN:YM_TQ,<?EaC_2LDQFYOfb8eHRAca8+()]FAMI
2XJ31GI&5./NM2B-+[NEGVKd9,5[L(@\SaZE-XTSSR23+WFa7,K>JWbe7T9W:ITA
+cLZZU<GBc\R\;#8@+-S#@CeUTA0OB)-Zc7g0YHdX/4^1</Og,(BV+d]++7(,UM1
C@C+QWOcK35UW)V);UIC5?E8>VRY1OP=ff0(#OMDH;3I@IN0;?2Y7MY5Ed^U(ROJ
6]ABd3#<93.dPLa@M,IU/2=C.]1SALTW):;N3P:8LU+E_a/:;eYeTPfbU;W?S9>V
gaA[Y/6XRPPb(Xd6[CHTJVbVWWHLf>[A>9\.UXR@\ba1IL(8dIdKM9Y_2NYSH^A5
;:0_3L,6d,1[-V>#ac_YWa-+-OEPF<L8M4V#>d9_7VVg5LD,&G^FAQX^]>P8eV3g
;;<11TK/GL;a/CE(&#K;3K;be5T+ZAPAaM0c[5>Y[H_gZ1]VX6B))X0Mf0VS.^6=
^K?B-=eXBRD?ICCPa(T11EFTMdD?GOR<0gKH#UfNGL#.BbWbc\ef707L?UZXbfA.
7NO(G[X#9cP^Q@[44.WJ4fdBNL@\WgaEAUKT\JS6)3GL)5XY.F>65&(+]B][LX?M
+(^P^(PgR^?\WNBX_1ZW0J&#fA-ZbGcVK>Y867DH>&fG-GG9PR/=F;/&DV=DQM_X
@@?3MK&V\NXZ\,>11ACJ1BNH;=:FTY-c;6J3TGdaAQ.U(0.+U3Z_b<V-[A>\c-fK
)1=G4MD>MSYOOLbGVgUH0,NPTC.=aTFJbXBP1aB>J,1N1=cR6-f>Ud34D6L7Z++G
Y>BDZG^]/)fJC#;AX)\-9:,1_<)G4+1)?GC_^UADaGKC;\/V^NaE83KO_cS,>^RK
C+443W@L2T8[_QL6A/WXQ?X&BHZ6)dI,3?1;(A]7KF9\>KK4dR;\1AOdV0TC51)g
>Y0gaQ24_QQa\/a.U4MAX:2F8GH;EI9,CT0-U>CCE(_R;C5XLg[2IL&0Z;(0350L
?4035/2ZZ]RaL(#a):4V3HHU1HfM-HUTfD,=6NfW?Q;6V8?F=cI&6f^<KfNYH][H
=^6[TXUKY^e;;+UaA,-\A./K,97@8,<4#B\V^cgJR(>#dD&1=JK9NE._A&+2NdDE
H2;:bgH=Z[4:2\b55a#DD)eGQ&QIKX)OT<JYFRFFaW?>gNYd2eaVfOP_;^Y8JZ8[
3RJ7/HWGb(K\68/1A\1a:WW-fPJQ10F+JGc_+8=[[(\,8.ZGNP(/@8\M,FQBH;P/
=\#(F,03J=._[@QSGLa[KR;_6_cW8JTN(<4/&V,E3R>S]D[&e1OM/HO=Kf6ZG.LO
Za8@)G_Qc9QCXK288P6Xe=d2gUMeW#b)1DT^Y:UR&6@eC.N\O\bDd6-MV1U9f;fa
L^TA-=U,/+:_&gCf3YA,FR_eMAaTbg@G01M_<c#,--Z\J?dK>:AQ9@BZ\?eXV[DM
CaaLPE97gX\L]DL,I.YC?@8(2e[6g-O-ASAVQT-X#WMI@5#08bQ<WZLcE;Q_7g?_
RS&<RG\F<H)_H?.>V@5FB<b7F0ROIH90-AH-..+8K:SC@1=NAO<M7gSae#7THI2N
fc?W8FZ?&Q&UEVdPIZON[BW5^&@7PE7a.K&Qf\TSAgM\2-U:fW.<SbKe.4\d2)CE
N9)cMLA37e]bG,_gG[gf2PA5>D[K&E><f4Pe+<;eQR,G>C.JbOF1,N-(?S-6ND?Q
@)>D(aN^FK]VF<DM#2^A:aaf<c9S?AB_Mg_cAaU#c-/NOYK^(+R,@W1U<XgG^DYX
__N((2M.eW.8(O9Y6T<,]1N-b0&/SG6.dZ.cSgXJF9TBKb[<XCgD@_KN12KB?b>c
T7,fOQ(VSB,]6VD+#^TJ6M84<_&aC?b-UTfU5U.]GE2LI>?G4=P=F1Ug:Q;4cb<e
0?;0\_&[?\W[>)F8J<0_F/9?]2I-a]G8LdR>G_LWe3WgQ:78,I)d7S-UFTOKAJOB
Z/YR52H:;=(MS.,XZPWgF^Z?-8=4fb&BD_#EH239d)ZXBV)VSNC>61V8O;QPCFB>
VB/SX@RDLYOPITQ+R+D)BE5b&I+7.dD=@SE_b.KJD7&XC6\9\()^?VIOC4+U^JQ2
1(X>H?@H,gP&17d6g2A49&Y3>_+Y>g)H)2:^7Z;-aA.U]EL\P5CDYEI\#C2,fYW_
&:P0<)9DY23ZgPW<c\&F]MOLVUAXX\8TTJ6QYDE:W2+bg=U=+MY1(b4C.B5?NKfY
Z8d6RZT8[ZQ&e,[5;R@_W@f)U^N@P,&MNO7aH#K#C>8=US.R??>cX>)\Z[S..+:O
g<@BS0ab;T-eW6BC;#XGCCEU]V1B&RHIQL=^UF>X=[YZ8d^9GeF?0PHU/CNf7#4+
@]ZMK#7]U/dGd6aP4U+7#WHWLR=:g#]bd^fAM/gKW9OCG+?d8HbaEJN1eDK0?\+Q
S+JG18@LYdE9]6HALY:2YL.P0UK6J/[O/G(B4CFe6,LR#)f/=c0A(>_fgG=0Q&\#
a+IO6_BfL&cKT77KOJ5R:c@-Sc<>c.SgfaI6L3E6OgF(7-c.76?P[+5]UeNZ6MDZ
-_3IY#&O@8?RZ8LA,Pcf>^PF8Y3D+dMH>1GG8B&N#+bg\Qd->^9(K+])LHS]0.B4
aW+8@eEaI\FC6[XHU\(/945AUZ[bW+PE-a97G-27M/L9eQZ?KP]R@_6W2g)HTBNU
UGONFaG,VDLXDd@NeE#^bDc@DBP^[(#X/d-&ZP_#->eC;?1<KB38(FQ;WT67XgD\
W74E<I-<8)aN9:,0?6DO6H18;[4RH@5^5R-+e@E5)+H?6/a[DfAgYfSU-P5B&1F+
U^X>VB5RGa+B.LN=OO;>9#7Y=V<Q/L0](a0Z6I\,LSdYR]S1L^^PbO0WM\dTV-/R
U44PC4/:Fd/OZf6MTAJ[(R,QVcWTP5:H1/<=+af3aO+A<QJdebC/>H0WG5OY0GOS
+@;HA7#Tfc8SEW08J\+.RXVA&HgU16JcbUN81LT>K)Oc,c#)AL,f_]4S8;<6e/eQ
H5_74+b58\&>FZc+MI]/(Z05QZQ2-&^][cY&WQb#.?RT-\U^>3a1+?OS:1/T_=J4
IETJ6(+327U>SC?HcG&2;SHf/FR:URA#)G^YCaE;@(5,IQ9X]+_@06.)X^&N6/YK
1d[(EI+0b?+ee[d[g1S.f;+eLPL(_7K:XeIHQ<S^P<c+BQBdP6LeGQd>MSg0c&H/
7&0bWdF4F=[<3BT7d+[:Yd(DI+-#R(:YgT@)]FXL4@@aY_PO9R6.fY7:W]9-G1(]
K0Xd6^]=)(N7/MC8=,-H#TMH&V/W@US+GHVb68@CcH(WJ,SSV+E(5;S1&Y,HgW83
GQ.C^:Vd(1ge[+MbRS6=Lf(_X][P1=<9WUc+B]9g]7;RC6+U,B.2#c[YY?Wa0-HV
aLaOL;?Y_DSH(e@;X<a(7fDc=ZIAbeLf2?EN_9=CT:Y.dU1TLQ_&;-[Q\J&QFJ/7
R@QH4Xa^f)-KFIR-L8?6(Oeda(WMW:D=QJBc+X]]@/E/5.HVMZ/L-;U+CU3:VXKb
/]0>51(.NCaR&U)&49gCWILg10JK>=BTa/9gXS#HfOU8DN=df,1N7=)-+aAEMfUC
?K#1_aV8L<N9J#5ZdI;\bL76LGX&N=X3YC#S]=G7U9?0XH]Fa0WS@A(eL?>ZECU:
14U#0BO3]F^(dD.Z0-=)BP8XYD6]R39URMQ0b#4DI>B._WXQCgMBC;eX<D>-VL#W
E;/UBLEEK#H\\O0<B&2O5VQF4#H@17+dPRW7QbJeEQdHJHRg:EW#73RP5EE&]?W6
XV37XfYFV]4e908K]GW-^)-T4Z=/X=LIaE6g#.cXFGJH(EMI8Q?0AK<I3c]/PP(D
S0^_+#_=<-,PRS_E2Tb9NPK.JR/BES:=.fJVJbaZRKOKF+^C0@c>WOBMGZ1Hf;/Q
AOFbX8?E=NKB+SLO3)9__C;KRQ\?4Z@].9:FRNW2F9I@0:<SRfRggK:IGS1WV@9D
=UL(3TbU#G/J4],gKfedH5G_FU9Oc_1&L12GcRRfMJM-+T8U9&YFd4UQ,HJ^PA_0
E>)#a3fD&0R,G>.9MbfCL6YE)94J<fVRZHI.PbKIg6J(^(@]-;2=\G5V[=bIJZGM
FOcI^MLN:P+DYE2dLIHBaRN#>EWL;##@d-dC;IcHU.D.&<KZ1<RK-&61D/[74:1c
22PEETBeOETBNPW-[-O7[5c.OgaE9VS<XL9Q:4;PDPI&+2Jg]->Db/b-(^>a=(gH
L#g9D)W@)KI4KZ+B>YST-gHG@eeNf?<[V3W>R1]e8V8\GK_F8=;W??>UJ:U>+T5#
+WA/ND,<[8@V^B@Nb+X?E&CL^9]dUVFIH]710QU:]fC5ZBeJSRg593.K9;AV>7;c
._^/]e#KIP3HfAMZNI?#adO+A2Vbg=Id_-7<^>J]NffPQ5QUAJY;c.ag66WT=UDG
W4P;F<gabV<&;PTVX=<^7+]STJ0;E3Q1_VS&6/-Q\K3->>/IUT#1QVD5.d04<.BI
U6,UP(_,DN[/+)Aa0S@LS2Zf\N>QBU>X34L&df<-2dYN:27cI.3<5caA.,d/T#X?
6M\b?KgIQV(P(cDYM)=cR#2^BLT]NU=?4#bc;=>-#ZR,C7FCd7<,gZ6#L0g,>U42
RE4JHJ9RN[0VBec>OSc#AdXH[(MQ9Ie(dBF3)#5/9.D\72NHQOVBUE)1A)Hc-92a
:AX#@G9BBbRU/OAEH]H/TSZUGJFecL+e0EW721(;O4()1K(K>DW.g_HN3I^H;S]W
bZYM,V<gA@JI>RFL]QHODd5O\]YSJW?ddXF[f+)MfUfE?cCL+XIF9YV1#@UX-faQ
9-]\PI0]=G:#6P>Hda3M\0(Vb&R[Xe8<ODTgVTAVQ[7B.&c^D,P,Y[UgBa&IXT.-
[FPb0#TY6-NcHAVWPdRXJL93T^QSDc\[48P@D^_PSLL(QaOH,3RK=(HY.]RYO&Q>
YGec(\NS:b[B<R1bDK\U/MDKBQ_43,[[/N#CQ@MX]S0I=a413_A\VJO_J=&ZKQ,K
JC>0B4.(8NJ_JGeXg&L1#).AAP,:]@YS3PN;8(GK1cY([,f?bWK.R\6BBF#M8DFP
](TNGf/#\3B)UQXN@P25@26X-bE33W]7..<+A1fGLF]6)bF/XJ7MT[JWX&>^O-fG
(b\7+#^LgQ;G>0,,&.(RD)L);;SDP,f\=QN__]C#;=>4J(P#UF<3e@+,#I7=e6(?
^)gdWGN/C68MLB&_-;_[K+3_,.OcOVd</DR1Ua8/4MAeCN?Z@JEIY,?5gD.FH=/.
MaC@2PTW(g&/MVT_a-;;ddD1La1eK@R)aO,&e,e1X:eT)ZPR]Ha]\^bJDcB-GN_]
R[6]<T5K#FC&T5,.P<EEd1T:9.0#^F:fdg5(_58gaWZ.)1;,,)2SNBAO:RMSD2K>
I5#_Zb25/?44e;ZfA5KHVK0[)CX>,_cX.5IQYg(#3dQA16:LRdA0.@Kd>ATZbeIR
4EeV2C8PMa++_F;aX?V<K09LF78,9a:Q[XXO->4gO/>F3aR6>VD1?04>C:7;554\
T/-,U/cP+0UgTBbP900/a.4/V8ZH2f\R[f?_H3AO&,7:.TIVK(DC@#8UgV?dFcU.
SIPMN/?S]JL4:LH.KIf?OgI\cPJ:+#GEbeR+Yd6_4+&0-ce4N(TKf>PN#cXROUNg
QET30D7[RCe-XDa(Xf,PXT.fAKN;CLM)Y&C:BI>E-#N.+cd]F_GYG88;23(cgS>T
Y6MGF\D92AUW?VL(I(AB?G66O4<:+<4I)B3B+ZD<XZFLEBW;UgY6\[-_bg0\J?S#
Q8_FKY2DYU@.e8Sd57MX^YLb@JPG;He6G;Qb8J(gAI-TG3eGCYO9YKFAE)=HcJTS
>O=_+.##JG#aUX57N\[_?K&TI:ID)6gL[B_P+9T4><2B?0Q<Ke\6gHLHU=eL#bdG
>a_VVD.IfVAXd3=cLbdA]<6\;(L3a@BD/.KF8Rc-K(W[4Z;)1+JBfBG^8X]V_9Af
J1LVOZVSXNSV)<b)/PZY,\KN,#6a;_58R2DNJ_+KAA0Jg1@D.1cce;S#T2cX/0Y<
A,e7=A<03OU_[(IB#d>QG17bWLdGKYT;:aF51P2Kf[C[EY&9G.IbW9afRaKY/#)D
QOGZ;R7KLb[7]N\DLL<>Hg+U]2,f/75@8[FV@9EK&-IIHE>dNP?S]A@dGO]7YA@]
JJe#N_)eJ+I7Y+3,Z?#HW^[9[UPCO+L]dT5=<cW/I4&32&L;_)LbXBBF6X,]=O\9
X^9T>QY5+;PY[Z(963V3c>^5>CC/I\U,P,7Y@@Jc/[<dgB.aL?1,66^9V1GaEQeX
>0Mda=HXGf<0Z<AI(8D>,^<6Q<;MdZ8B0X5MK\R,;Yc#4?9W,b6g9d#N+BM@AD;(
a[V/Tc34BR>>YFI0J:)1N/93;5^+Lc26E(?FR^AK359:5KPWXUAA/NS7VX?fH9b6
BXZ<I/<d:73f1CT>?QWbVBTO^0g2\(T^;\=UP[R=ee5LX0@3bb_BK<N3d.eN?EQ?
WffbBc.^)13].87&9SW),R<YFTT6MJe[_P=<0McHG0gWWWBA5.XC:D,gb)34.dT^
B_X@W52eCYOfA&<97R1C9YD]CfQDXIKcMZDCc+;_7JWcX0)aLQc4L?aKO?PKKEBQ
NA<XS<>#O@T.T3-4D0:@Y+-4=dD.2+Ye?Z4-.AfUI8-)VV;Y(CHI3(>f)TLHGYDL
B_5H:S@3BRD:(7@f7=G/6;H-CW^1M?8,)C&Df1616#8a^9U9785f^\LgFL)3+b0.
<<Q7Z^0K[/);ZWMPI09[EJ(PceI3R+51=/;V6?agB<[eFTJ2+HOFE2-WeEdVZC7H
4c2[6+N5QCGDO@4(b^bQJ?\52cXS2cR7X)aL:[Z>).fef8T3BC_<ZA,g4-ACI7:<
484U,]>HE9>6IB2+:TPD@WZR--[A4@(3b^N>AaN?S5:69^(8,)VX]BN\NEWCIe0<
&],Jd;+8;7R#?dN#W,L_M>X9.UA70b&0aZf#64),BSaQ-f;<65?S?W8<HKZ.9<KJ
df+gSV7^N>@fLV5AWHLaG2dYK.KEN1_e7]TX#:;D0eD^FR#;2OO8-9(.)0HD+47)
NM:9H:.d-KSU_>/U<<@/9:<8X7.2+,,DJ63WfRZDW\-#(K.G?]HePY\:H=]aV:Y>
#QC3C.8>\?P8<L+;S&cM@F\)XV3Y9da>TDT]K:,Jc);X@OJC?RME:Xb>L6gN\GeO
397OT7W7H:[aF=UQTT/=)_P.g=DX+/?14X?+4)74WESF^CEUX0HHD\<Ca3bK-@[9
3D5/,;a15N7&P]2)ZX?+4&LF:;2XYQP=QQd=Ma(XUDN;E&@,UM:(RKa[G33M30[(
G:0EBd4YX^<AFeccHc(L<PCXYDNYH-=N_a1PX)cZ(RUMdDI;1[1DMeRZNA=:B,G<
C>/<_G;E+:CJM,2d,8K3))1A1fF&I;:2=S>:YdFV26C\d/a8GZ4ID/Yd22JLXOS9
&d&@2+TA:?M^/PWM=\(=+cf&=EFCZ(:eSOYPbDWOACT04_]&c3-242fSfb>SI;HZ
Q_f_9#45]&=2VD],+FE?PX@K[.?9-b3/D>:]3=6)G.]W;)CAI:KG9K8^5CF5.Q\I
LI(&\)Y3VT/0A4;WQ@)Ee[4&E:J=IL7IJ+2b@<J9[C=dCNUKe65,]VA3Ic58)59d
H^XR18KH()24FGQ3/V>bK+2J7,XD,RE=BaJGV,5Q4NEda9[9GSVMLFY0_S;Va03L
)_R@FaK]\c7NU8#@6d6CSWe:4#5GPg2Y=JZ-.b0UVd-DL(7cR-P[:AC.7VJ6ZeA[
1_3J8M_M:BFce2]+Af;fTb.#W+R49E,KFM3@bVcMSIK-Q=AIY<=J9?WXObASK[6A
ZfF9b+TJ&P#K(HG4./+9UZ:YQb+3-DJ<+@?g:a82XJ16^VW&LaFfG.HfDX?b?=TO
<a;B\T_-&=b]_9A+cBf8TVPXbIK#-bbJ6YS&bTb,BLVDLNQ[Y^2D73SOT&ZF;efU
6.OT0QbDN<C]R:1O#:EcJ@V;I29E@YKM-6=B)N3##7eJ=_D8c?P]&8(:4[LL,8UT
P_-6P:E&XSGI-?C6N]<<;53)JVE(21X)QD[W4:ecV]P,+ZAe2F9db@FKLF>B(2)>
Q2W33Ba246B[3aI_+-=0Y6\3d8bT3V]?X+25^b?]:R8,#79@=/bV7A0Mf],EQ>MC
0EIf_6\L@BA2Rg0aeG>=ePIQT:TLDf<]E]K7JC,,)8V.QR_LDe^e7/1\G1LX@<;/
^53=YbV1dQ<MJZ1Nc/,(.f<.N2,)9WIL5d0<?M6>528ACF3VbGg?Ue4JB7[S,=?8
DX.2YF&2P9-?e(X=81S7OQ&1.3PGW[@fY#UQIIWP]#B8),)O:Ra.?OJ4.a<[GMcS
TeA=H@EeAKWg^Z4@B:=,(gYKdef^.C+SIdZ6Q5C6[HUUe\>9?J,dPM]MUAFT6O,c
#K1M:[&T>NL5PT]Y.R8QD.^^TQV#.FKNYW,_c?-GIHN&YQgRdC&)YeB\eL?>)=Z)
F#HM>_31&N\Ve^J>\WB^O2b[/EJ\L#Za6ZAJY#IHIHJ7;b2/KG/&@^0UKa@,,d)3
:D<YOa]PU#HA=:aA[;9Bbf)g.JGP_>8_H0UQ^GGP_[I]8EG?<7dgR[QDY.)W>5b8
Y<@4K/WYDU7S)U&6?RHIH<8X4IFA#.QEY?.ffX)J;<Ff93H#G>RKOJHeD6\E-30F
PXaERN2HbWA\E)Pe?91C4&;JR20d5-[L@X#d[S^#H)CPCN?a4Sg8g1MHRBNUQP,V
g(G:?9@ScZ&)J^(G.9G&_^PX5>CWZbfHb[2^TDWT-P(WgQL&JL.B))TO(TC.@Og9
/MYZ\WX8=dHGPbXYG?3,+bC@?6eM:b>AO-9FME:]\C-Nc--:8U+UZ82dL,?7M\c,
?OE5;)ULM<bIW41;0?R])PUXC.9P]RFC6)S\b?GO+g#+M4[B0A0NY8MeSedL_cLK
D4/MU9:4SXQS@3#S+N@ZQ^Q&+W(F^e-Cf58#aaWB>EDNA)TDTE#L?9f][fR3M4I,
-D(O+/T7A#0W_d5LJ?MZKG^f4\[WP2T6>JYG0.f(6H.D>VYDf:f+?L;6^^fK@PP;
#RHF\F]E@]7#T9_.28<@^GLH(/L-O=Y:b<:I;PCH;#U3Z5b\I)VB_c@&>E,7U6SU
Y[IF:7[VZKb4+6Kd&4fII)E>38G5e@0OMFW_ZN)>\C8/;aV#O0HYeBdBH?#>Z3aG
B-T3FPGI96HZG_aEHF>4JF.g7#@OD/-UV2U[FCF/3N?D6V>4K81?+c[U\W\+5d3&
>.=4VWd2XJTeFL=58[cLOZQ#Z@]a)V#bE_SI5&8N1#0OZ<V2BJ&:-,NB[&FD(J_I
&9\AZaK2R^R9]^G,]BS:@YYA:M4MRGQU^@KGe#[CF)d#(GNH)FKLaWdMePacd0WM
D3<cT[0^HAFWa:[0=;TbA<4X:83\#^B5X]<?5:)g[+R(F]_gHMO]VB<C=UdR9:XQ
NCC[7>.CT#4eDFYM6AD.^IV/HEgLO#BOHIKJ[[a.,HPH\\OW30BbeMC-:)PD2(JD
6\B-a#ed52?9<&7]4/ZLCC97MF(Z()Y9B8,+O95LPTG,6&ESU^Wa6S0X\.NEDV9J
[/=#Oe91_&FTAIE1>.)Pg<=QaAO\f)JU^+,NJ^MF;_CC\>;)3=HCc.P)JZB=#1LC
Q)4U0A/VKb>OK)+T2#EU4:P7aafW9e/;TQDPSL)TcAHE/O<3.P-ea]&K?;?c5J&5
NZZN3E#]+65//Ma@4SK>OLV&fggd0SA#;1:Vb#P#P-XW0@cUXPaePIUIAI-S:4:S
:G1GDJW8dAK/Ma)cKGF1LM7=9MX1.eU:_5/R2<dS94=TGHC+Z1]1I\f\AOSgb:A[
Ce@T/ZE@LTdR4XZ9)3_FFZ#9<bXgI;#5eaH3O?\,gD:8<#M=:ZJ=+@51(K&6a2RM
)N3C>5gE#]>Ie;KSQ?&XLQ36).VZ?]_R,@Q@-OCB5^#SaS&&1Q2]5@C,8O1FEK(&
34QR_QbBUWL3UMX4/=7)GF&:F7=gD5+L-0dB/Y3[UI#B]I0PW=//.BbH,0=-Ma&S
LGNVG&HZ26,F_)Ac<MKP<K_M#3&T+GO=MZe@ZX8ba\fab>gD1>EI+]Z&VPef0-;f
g)M>d]41R[g/7V@-@-f4I=9.Qd+]I0?Ae9AIQIL.D]5,HZ#OX_.I==--O48UD\^:
06?8NVAY\]^Y>@5],<TT=SR_:7]NSbQ@-&dO0^LgaE0QTB9U11A@JZ?Z_6+ZWX/S
d_&&\1(8Y7c@GS-774-YeM2[HSJE4K+XW^12(8HWb(<2181c7^&)]6:Y)(2ICV:+
O7VfT/DV_;gJgM3PMUR?+,\++_#D8d[(#Jb?9E#-.2HZda)&T?=_eTJ=[L4LD[Bc
]#d_:_^:DK?a<K#+_G[C&#D[2K(/JM@c2&]3(aT-SM(4C100XY#a-c.)fEZ_P,3@
GG0;;a.P^<8Rb:UU]#22SJSbUD9D;Q2.-P=UV7b(3Be+4Q<ZVO6LR#=@Z8CgLAOZ
#SZ-H6>AI82C3JA;=<aBZc0ec@L6;:8H5B_.ZG(_=bOR-.&/^U=Z^KXU0La7aJ#0
52a-.7[C:,aT0?5>;Y-K&5G9g^:664[<PF3dNV+#.+7+YZ[_X/UQC\^fO@9[dAM>
):APf[S-?U1&WK>)438BE(+gFC&7Ff:NA-:Da6bScO,fCDB[b+D+)F@@I[D=&JG2
L.R\.#-Q8TV=aMfTR\Q2JG&2:?)P^F<?.FS32QW;-ZD3B.CD[FcS\K03<PI29=RW
3N?9M]ecRb#]a,L>(e76;F#aCa@JMSCGP@4fM.W(U>>cG7:?))JSCFL(bLFD2Vaf
f4X4IBV9BeW3#eZ8-)@g[;PMJGKb7NJ+?:S#bPBQ[_Y29?c0P,\>8)KA6)5Od&/[
a7\>GE9/-3-;C8g8T1J2;\Z2f8;T6<g#c5MS=A1+BUFF>T9;:/8KOR=Fc7:<UU)\
QLY6G5(2;DJ<PaWX#29aF;L=)WW@gRb2;\6<_.NUIEdb]C6^CZM=@@SP;<C-N?bb
&,50L-^I5XO3&eIb?##GF)E+R9e?:b2(f,3G59:O#()KVUY6P45NXZ6LH:L7?:c+
JfR@^J(&46P&80faf:-\TQaa_1HSIS:\YAECJDCVefdU[d?-a9KZ+gb64A1CDLHI
)/(NLS<XG]=eG0.gO@d0)G.[:7:M3D<3N^0[)JE(e?81d#D[R674dFdZZG>EBFK5
W1D(<g0Lg3[B8O2B1;24L5=7\acHWS>5cU2@6YZ+[XL/(B6K80).(QD+Ne<U[Hc9
4IBI3b&_2J1BZ^U>Dc5cOR(_3QY7J8_N.5S,GPZE1[dHI(.W]X#XK)&.)4+(]>d7
HT^=aNgV9OXMCH?1[KGIH]J+THWaQDJ@eeGdAa)-@GA>WfM&c1W+_=[O4+/8.c\c
NLMa22(7:Dg#</SdHGVOe1EXTE79FKMZ_TJgK;K74Y^#8<J?Q?CA79T)+Tb2-5c]
UMCO>R^G;:QRdM9E=<RSN6[VJ<OMBZX1a(R2M=aU\(?RZ=+fC1AGePSf2W(](0-6
T;HKN:bL;=X0M.TdQ,.DL/3f_3]N;))V(&J.&d@GV3^5L;POEJ7.3>#J;e/2LSVP
g(P9>^II9I<DNX9AC[7JCgNPO?RN6<(<dBa@f,AbK7+\R1#g\,S__fYPP(X.U#DX
J3TU[JOTRfX[X,SPTB0DN9E)?G?5EO>=6eE:XfW:U[<0ceWFbJ)P;_2B9>?W\2)=
<72e[:;]?dCg6B?3cEL(-Bc\,d4&4_]=ccNG#AC^L_bSK@5U71B5NUgK\ZLOFf&-
g>a11LL-_LfN:g_0c&JO(UO/g+J)d33ZW#0A\OZ<L7;P@EK2,P?@)LFS]7M_f/OQ
N&IUOXCWG3[C;\>LV4f57]5eP90;\Q?c?02/a?G:GSWRDM;Pc,f-4C,CN10XYaTS
]df[/>W\dTgg3Gc<(SNcY#-fFW)Y<O(#\29NEf@9EO9F>bK>?YDU4:4+@+Q6QJ+I
WfO>22KJ0[>^(285ZPL?/EOS)^L18,ec&(a^9(?>eeYC,8;ad>Tg>5M5&f=QF9Ce
+=CA9#C?9(#(KGU->=XT(X9/_XBH/+MfLB##>GHXa[<GY-:77Y0(1OZZ4;F(HU9I
.6ZUCE70.3@E/gHQaXF3_\GAZ\=GH,7.P.fHdD3QYeO.0/JL0g]DEWR(9-f0(]3)
gG1^]\T^RdS)ISg,<3Q@LHR6+(E,RVe6SODCZFF2T7eEKTbJ()]96,4SbUO]6<1V
2L_SW4SG\M1JAKVYV5]@(01ZY,<2d[664UI2],1\2[32U8R+.R6BMfKTIN0Ic.O\
dMB#OCZLXN3TeKS/GGSNOKY_/?[\E0@H(c3HRdHM3N=c[,IJcA[M^M)U[/^A&\XF
&2(([-Z;CP4_K\QW1QgJS35,]<fg=-GGcc;R.E,eG-ReADOV-&/fF.G#Z=4OcTA)
=ff#>G5Tg8,8MWe0(^e5D<EWc]RBVOL(JQC2;A)C6[99YHFc)D/b#F-+dLQ)-8YI
)1\N+WH4HF^0aa\5?0&\ZVCY[H1IQEY1+1(8(NE3WC&3-^W?R0.Wc=&L(1P;MYDV
9QT9bF8W(U4NVD)/&<F2\d8WGK_-:<SY7T6IT<72ZM,Ta9EJdMM&>@CLOHX.XRKG
cY@D8B5293feYZ_0U+=Fg34d;DEPf7K=)]URS=48475gNgWUEH3^YA>bW<^fg=#H
@G&T.I+6.9P38&gNd4Z13d\#/,4^.f&]Ydb6<6/dU#T24aL5IZ)LUD/OZA60/VgH
H&^FSNKC8.:WYM=d@d241@4;R^W4?=+Df_);eW+.ZBBC:,+.EESPIFGbK:]B.?9-
KSaf1Yc^If8V=AN)WH^.;eXCdc<3GJ+<Y/O-4A=VP3:_V=CY>7N+Cee7=?TD+O>C
Gf.#OC0UDH0UeW+bd1O1fX&6(eWeB4>F.F+<fV+FYd=fO1ZgWDN+S<eZ)5ffd3\A
WU-HP,[R58XW3IK0a(P&F6@13?OB=AEBXUECOCa_WTG()aKdQ#CQU5FJXCT9,H[,
./[1,gbC?H#cEd5aI]Q/HX_O)R/;Hc:;EdZA@+QMM;1d.T6bLYY.^UY>bNDQJfQU
?;)E:UVPgH+RW2UAdO0?VBaf9EQ6,Q8Fd&^E+@<I.DfUN<G0UcL[\C>X=.SY7^&5
(S&VGLR;3eI98CP^/N8VQN+B+S+b8T(cV9VbIMOB-b=YQI4E=@\=c9FUD:X>OWEC
GXRMK.X;150[W7828[G3M8W^--G<T3<:RA?RN6DFaG&G,E1IF8EdE/QQW-;94/C)
)<E3_7W))/.W9U<FAJd5JL^Ub3S6C?(NQO27(Y4e]^255T(Z;?<ALJR7E(V:Z)c(
aHe3L(:AU.N=)@;)9Q-YP3J?KJc(C9WbHS]e,W(&SRLCgYTJgdaQ]6>V0K/OeTPa
MPR\COBT?+a0/I>X#)T@)Ib?UR=QMa.cU?7YTHJT^8TK9#;Z-,,J[LOVC^FGDe:B
C<ZQWC.F&O\SQO=\7f16S5&2FUSP_9NED2,2LZLS]af]-I4Wce78=J]P,fXA])=(
0UHXP\P&NU>I.07.@Og)&QY=PN:Ha8-V+<ZFLF3B;=5)=K2K/F02:Xgg>;F5f=R4
YXY0X/-2^/MF<9RgQC[=g4f&IEYP0<L0A;2-\G:C,)N4WANAG/ca/UN>C11L7)9?
)&/cXEYe?<<9-O-KR4<YUL(C2MQ1M_K=?gO06=ZVR:LBMK>dG9H/(W<ESZV2_5e?
faVX-GV1Xb?Q[6KBe]>efAOEF=#Pb(#^B2^W2]F\JF4;4GJG(&19VL&VP3VeE89S
7.F76dGdBQ=UgJ.@73I7N8Kad][834^D^a@>PO(/dKT[Wf/9VUKYN4&f3;[@\F5-
:K:_&5Ea_(gJ>1WM:gf2b(&E\V=P/,\Uf\PgPP5MPX90C[Y]S7GaPP)657SZ0NHO
6=,-K,<>Y<ZP1YD9/0)+VUXe?E70IZ8#MaaFA+;Zb-:(_GcT0Pb/GGe?H(-DZF#H
SL9E@a54KF=Xg--a;(+DH6XY+/,[67d16&=(e#F[W20G<W-HOG\b=59W]IN)T<&)
S&HH6.IJgWIG5)&a#VP6?L=Y\8F6H7H7#AIP+JJA=e8&)fVVLa13?V-AE+:GSN-8
UAD6D;2,:AZ.B3W:ScC2<?>CB@F^248=.;7H0Yc[^.RRgEH_WHM;I.gZ7//D2D)0
+@AU69E_/EABNWC7Q:BZ.Ye3.8W<;EX-,UFUBQAZ+@LZQ\MY=7g8QQP+?VN5ZBXO
+-21:WD=[YZ5BWc+Xf)#?f@fQfV<)b/7\JbF&Tb_a:=]MEDROZDA1+0J;VI5GHA=
V/.8a<8TX/E]2:H,fPge5T7N6KY4/^<d9Z&e,O]&C=]RM3W#YaK;?>=KL<RK@dM?
#JP(4\0-(g+QAeQU/QP=N)bC1^W;^OfZ,L:@P+ZPZW]Ka)S):<CEUKdOLL=?>A-G
85f-#Z_+>9@+(LHM<60L+Z0NfCYe_?Ba_dY7dL+ND63_Mb1<W549B#\/>MMO5FJ0
g=STRA[DaUG\]_egD.E<+KdQH54FT:NSbYV5..&?KeFc3+dFP+XZeP_BQW6CW-P@
ID2FWeU@b>;TT.CSTUFR?X&(5:g&9;E8cL_W]@MDe5F1=,4RSD6GeaH5M[<JT01[
SUE<W81J)Y48D0N52O6G,A[D=RNBP<I</EL-e&\OE.ACDVR_RKAVX\+U;_[E6+8-
Ff)RYfTQgO(+(Xd=1)A_6:BHaA(QFOND_cS-\@Ze144>aPaUf^bRA7;SX2Q7.KS,
QSNO/U\E+K[_T9C-?)g>\GNOWC-.gO/Tb\H9LL>>deea8<X2DXa51Vb@LBSe9b3@
\]1960cAb:Z8f&?E.Nc.b&fBRd9X2@(^f7F=YcAWL(CK\1&?UHAQYQHMG)<H[c#8
B[gbZZ.Q&b\AQ0Sdfe<A]FS-Y)/M<>TQ9/Wf+#&J<=IC@?&A(W&aP]^a0:.>0a<P
,XaddT4=2U2a(V_KV/.V6Z?JF=?#?GM7Jb57B.)F62G0J[I3W(da><1&A1,8DA01
Z9(#^4Rc.R.e<DJPBR#-34g1W?XaG;1Y,Z2@6dDeKCME=J_>,gK&,.P<R&)5=cCN
(XW)/DJ1=4T@#ga+]XETYPdPF0E1Cgf<a^UBMZV[44BO;.]>C4,AaQH[8G#3T5I-
1S1E^TA;HYOD@b#M.?6GLfA:@Wa7M)T,eA1@;3]))>4Be#;MbQ(?W0)eSeM]6/QP
V/+YNI4O,4X_aE_Y/VHNATBNG\Q&2Uf6#S_9T3P.dDbTa.-EG,ZJgWBg4;^6#dW^
-LQ7/J5JaU.d>0G7#[cg+@P&e:X2aVV(+WSI4SS0b<:7<;LXL_[LXQY_gZO<F.XV
049;#D-I3P4.@P-&@OXHX[eL?FHNW9G6@>P#.C5+>;c:&a7BA3F/J?NP+/WO(:d_
+)aRaIJ35.]9P1ZX/A:0d3QSK#>HJ7aP#b;Q<L;5Z#>@NRG/0VXbbg@-b72.:@M5
[IJd_8;<?f<Qba+gSDD^5I9I#fO+(6Q;#SeYMKM8H[J7U0(HUA+cY1eL?_b5A72Y
(CCA)@#GZFP;#JJHD6C7PM4U5f:c;-J(GN;G#3U?;[9J\VFeTbH<Ja85\3BU[8X7
R(ON<e^;DXTCB/+V4A?4<I@^[F]0DfCD+?LI[bgK(?(:]ff9bVcR)_W&CI[F>.6:
V,LOA28+B[>1VU\WQN?[LP2ZaXYJ=dO7^&79NO];Q[eH6_a1=L9_<@TPJI),Ad/b
1V&KOAS#5L:b:UcS[N(\?5295\_-cB:Jb<.52b]5:U:-3E?XI]#7<EC<E5NK_UOb
cG/>H#;cDB\R0#4BC]G&NF@ee\N+MfP?1DdFF@_>383/O)KJc1Y.HPSLUB7.gAN,
/Ic+K8CSGH&WcVbIY_BYZJO_@1<aSKNO;G(;J#aLR6AP<742BZ8][TQ;;28[@>.^
^_T#0+491K9#2D&f0FDQF6F]e>IefCC84Ga/TTMR-;F>GAYPVCC=CYefI=[K)QZf
becb#M1Z+K4:,@=e=#4d;74T1725K;P9C3AVX^[A)Dd7E2EDe>/4-E/[F,gA6XU0
W85Pb;A<2)Hc-3bD:.=K9Z>>6[BA+CO^,d=e3g_<Fg3R1D02:d6OF=/AFaFe6OEX
=-\V2WER?Gc8L\#B?GK\0RO/GKDYNeWIa_N@@[FB5=/49N:3((5Y.9HX[(&8U>b@
<E:^NaL3:^(W^dN<AWc,-:A6:]Se8+\YCC3?7GC\W;G.BbTQ/M5J].=e2\5?<O7)
\R7aON#7]LDXc7I)d#BGZ(==0eT_+VY[\/g_DFLJdBf19ZdZ&cQV=U@.KNX@]C,P
e7K\8&gbEDLb&7,DA,WIDfA>Z6/d5B_J-A.<Y_=2WKFA]3WO-&]0D&JQULdgZ>(R
_NN7M<E_:OgIB?LJcTTB[57g&;WV5B]PWS3_cG&A69d>3LE0F-PMK=R=?.9HbY>I
_#cXMW^RAREbGW)=.I<(-&FQ;>;OYD?://gQE7@K:^>\+0WJbOX#S>.LG\1<?AgE
93?;D23.@0AGK.X@UdH&CUB9]:Rd&1+Q\ULe\J3bOL?))+DFF:#O,g30a:+ACS]5
>H@OUbFb=&a_BT:[4;&ddWP1N0c?1X(Q_YMWROf:O,QZaG#_cG#Ra:f[>]c#b@AO
@Jb90>baH+2_YF]+M_AM7V?C=b0_)B/gHL=C>?YcP4a[,,Y&_G5NF.,,@X=g(PG/
8#UWNgg?SS5H43c.+a(D@YF3C.3OJ4WO6bS78+9AGbGPY\72:B.7>82GIcNaBVU3
NTEEb+UT&bLGeY]EG-H0,MgQd[\?c,6&eE8(Z6U7(450d<VMJX_(-YLMU0#6K-9A
&)OEPe&aW25B8NTNNg6(LQa:M9CV7YU2U-H\Eg#=3)OgH.3ZNDYD5L<KaOVZ?QTT
ICU,2D-Vc/IG;VWdTIAUe5[AE5N3b^-&e[OYAe2MYK?3V0^07OB.<?cUT55X/5=B
3L/G:Q.GVFacQ&7<,_FR-^X\bW74CW9B4G78+N^6_2LaKJC4B7DYKV_Tf))@^d3P
Z[KA6/Gd;;DLc@GPM-9-SE-6):T7XBU7J2.76C9dC4V(ea49C/6Z;#W[.97RPg]0
=\Xc-O3P@@^XIOWF3VY9b8d&b=C94BT@SX+A8L8aa>GeWQ>(P+gIV_ANQ];(I@2V
XN5]LMgSF@;<+8655:XZPH;<637YV8a@/8I5ROT;&9S3#<<R4=cfc3\LP_RbIgNW
2>T4?#9GE#[_Ia\5d9_a.a#7>Q9e\JaPdE<8TY=eX^I4MH1g7FWMRHg+1)I4IMg,
7MLS_fGI.1[7-Sf,5=JFG7P:Q5b[GLI)0P5BWAE<]EMdSUM6?QW3(7/HPL,FJcFQ
]55c5M7&cg)d?37I&ZJW,Q#d0Ze1f;Ug38DX/9P5:;^TLU9Y:<;1&CL&</c2ZLU9
YQ_)+BgE6)9Wb:0Cg]DCIBHT@OdZ.9L5W\f6d.T8O9GQe]B.K9EdT7PgFJGP+#.2
1NA(;];5d\\Y_<;)2._;P,X)0G>R[F/J97B3g13XD-S[PcJGUE&TC@JXWF&ZeHc<
[8+Y4HQ-2>CZMWNgQYf]DBT3_&TPF#1]d++8/KafWa?6ecLYLE4#BSJVGe5G4G;O
N<-DJ6a+#T[O+1Y:2IU6W)-.Y.N?V(J:ARS=JgL/71^ZT\f[N5V2=7(W;4@+B;5(
7:M-6X69.XP5RD^G==7KO]>gC_-gR?\[0F0(LB7WHQ3NRbT&2]#_B=V/+=A^g+/9
A<4#(3/1DZLBJd=<,K8[G#(@[Z(-&_CDKC9(H.J0Q2GUT&F7QFe2A,SRK0C\#HD@
2+@C@V;?7e:Z,=FN7a/T_U1WJ<f]_AN,c\2WQ&^EYHdM/f,<116BU>MQ[O9YF5P+
6F(9e2?YZQdF)Yg<F;.^&CAa<?22=9E3RILd[OVb]cRI/9ZO4SBFed+](4A=H0#Q
]#MAFNJ_8L=TU/6FKY@F^LEW)CF1>W)W9@ORb45VW2/gK2Qa/1+&fH](S@<Lge.H
4](T(V^IVJ:cM+<,Q&d]M197XP,EBUad<38U[LHRSQ4PK[MG=;128R8L64c<&.R(
EO]b<8Q.<TO<&<BDDc]3Y3;X_Y?4PWW7KOXW1K\0-Y2RQ[BdZEe:J]SW?bV-T-J8
)FJbKYR3HgJ]e&8I-(eEE.A)_.T:3b4,]-++W((38I3X;5TD//&5(L6QWJH9_8NP
OR9]&83T\CUfZ;OY6e[L^a&Ce+EacS3ATYXWce[O8Q,Vg5(J16BgbMUN&:OK\NSd
([?@Z>_46=3M:[Z&(g266Ecc_^/c0CfLD5&O>:EBRZJg94W5K?070W4/H,X9-?:@
8aD3_bEB5HIc5=44?ff;C;JB(ZNOGL8I^71=&1H5^8Qc__:X@&W-P6OXD<:<2E=P
3U]8geFPP1-W8?ZcS)R/McQ8XY06DbReI_APfZCRE3ZOd[87K5<Z6:>NP<aaIEZ=
]b,)-<d#^dc8>?K;2U6g-EN1,d;bMV9g1RU6)CCe7MD1Xf0QG0=Nc_BFJ]&W2/6_
&TOgbV-fL+eII)a]))-^;XaO+a?cU43QY-UdB9H7&QY8Z@F\>KV[MW(CaJ(0=Cca
3eCK:KJ]0N0ZC&5^&SC=&P4b)<IMEa,W),/R4+Fe]NV7>@dIEVc-XSU>.54+?BYM
ZbGX2LA<1GJ;f>MNO16DbgSGUD<Q4O+W1gCA2@G15+5CG<Sa3;Lg\ZL@&2.:^&&a
F;N(X[HD<EgY2/=6>63P9IO@;VgV^M<4MGNW=?E<ZHCIJK+_)?&98/R/X._59V2S
1-+RfGBO0,^XaHO7AG0M5POPE2V:YW0.H-^a=_W6([S(f?QQ<0Le^ZWOPC]c[VfB
=GFW);/[WD7G0e=Ec-KdP^ddPNaJLKKI9RD2I:\84Q/R#BJ+:a#_W6C^K#RXEZcG
RWdYMdA,3)M?)_/[EQgIcMf2<?LfT=_6<M1/;,F/:-N<Nb0e?R/3g)Vaf,:&HR.>
<2DbG_3TJ-;eeWCR77U&a8QC3Ud=@WVA?Q2(TVVD;@5P3_eBe&X61f0I<);___Za
/@&MGI@6M:X#JKWUDR?7+O4<cfYc3TZ2&WPCTKaDc1e8MTZ3UI+)[(J:+,FK#\F(
.LAJDL(dFPS=)g_DEOL.B(eL4[AB&NNf4ZZ-0,5(0ZNc^eR.K,3<M?gHJd<S\,-]
/<5M]NKcW7/[+Z71>KJN_(Ad/UO7H3Y>4N8=&B]-a4eZ1T1Va)e0GCg#,I8<dc\I
e-:e<>M0cbUVAQ&/DdEPD&/5=[G(UPT1#[[QO?)b58OV4?_>D.E9fFG(23)Wg^>W
:cGb@NIYJ3D#@^)N)E)O<5F6ebK-/?)X>TbdQQ2GC]gW8PDH:HI/0B5N2P/K])DK
I8FFW#Cd;Be3+BSdW375CF1IfX_QDVWa[NfYc(RZE.3dQ83VQZ8,ZIT,;20Ag=-Q
P?<4a&X5[AC7F#,,C5&L:FbB8Q(F;VO]#E)E?Qa#MAD14:84b&DD<e;M^dF6,U]C
4dOAO[6A5eVP6P5HU@Vb6ETI(TEe:ND3G]+:gM@N=EM:ZDB4M#8XQV=0Y#[Lg?d.
K&O&c5=AP/[DC85^B6\VF]9UgQ+V]D[MB;QWORPH=)M(T4,&P;[6/_I-ZSa=->FX
03gdNH<fUP.9#4-0D3,R_a0\b=2?UGGS<TP5[5d,FMA5d=Aa2ULP?-+=&5Z6OP25
T0b0;I_?\H9ObX_147cC)J1[g+^FZ4fZ6Wc.]D+CGU@fd0.6HSe^6QL)2R\@M6WM
U.5eG>^JcC4bN=;O?QRga.RI)V9[D4:efKVSB:A(gP=O5?(@@7RHb5,9gg1TDXBd
G+7&BDDBe.:5\+[;URCO3H.Daf8FM\aH@b>8:?MJFI^N#3R,2<1]URUTb8V2FO)Q
4U-Pf(Q8M/>Z.D;MQ&J^KD]T5[4g?C&NX.=SWVI)WCG:>/?E_(JZF.71SDP)J]T(
cMO?>AO,d#;.0BJS>W_R]B93#&,Q(PHc.>fIcb[E&D(Le\]eg(Nd=b=UUF:ENaN2
-)fZ3dc]()&16N_Q=daCXXcEJK;][bO7@bX5#^J(N/ePSJ7C9,LKN2Tc?=c]_cYC
=IVe[M+fe)DBGAWD4gC#3_>A5+D20fd+J/7L5)<H-JOW=Z]QS):eN^9]P.1+ZT,d
O8-98-2K.dXPb#H@;b;eERK#NW3MULZ7Q_,PELJ=2e#+\Vf3RTRW@U5\#?9EDY;a
1d3fOb(Rg7INZ6[&aCD>121TR<75YU3f2V/V(]OeZAPBX?+B=V(ee>6GH&0N<gWD
Q,+J3#0cgg4a[TXUF9.G-:GJ.HIAC,CT(NR97_c/KQ[&:MI56dLeECa@?.>\BK,J
M>JY]FX(QO^e[>Wf(E\;YN/QVf;)P7P-3P+:D0(&0\R&<de2-)Od[NCcQJA.0>?Q
KT;e:?4\U-\H-S#Fc_agPS?<4O0e22,::TFG20?)6.VcCX12Z^0X3S[@JJ0bR=J,
==WDL<:E^5GII6:Y<cPUa<3c:<NObV8;#LBQYUc;X.//YKZ];J]^A\NgR_4)EaXK
cV:B;b<;<DTAKJe;[DYgJE5ET+Ea?E].&dB]V;JXAGbCO)85C3;L:KN43>V\VD<\
B0ReKa[6#F=XdNaSH:REZUI&g7beN>THHJUW]c]^NGb]Na.>_FUD,bG8O8TgE9f5
@&P,^7_6deA4.6H8Ec[&bb2&,&)#CCEQCCgC<?84)df+TF)6.fNU+S?G)Y9ed-4;
a(Y6P:eK+QRI8e-SSL27D#5A1ZB)/eWQ.Y,T#AX);_435KMC#H+B-R+LT7Y8d7RM
-M=PKbJ?db6b;0gZKc)gI]:)Q))-A:0RE#G_38AT7JQN9.0HU=J5K(c[;@FO\gHN
VM_URR:TdOX(B=&,YKWY=d4#0Wc^KVcH^1L(WG+^;-KSI_,MS^,cLVN2:Ga4:CSZ
^,\XPAB<(IU3JdITY,(W3daDD9I/?Y.Q>^0/RF(OT-O<+?FXES\5CXE.J4#HZ_.8
_V4A56TVWO.V5\K+D-@8VH)=^Ce\-Xa)#<)0aBea=,-W#;X6+YZ^f9D?77H<25EM
<GFQSI:0&].?YU^<,dF0agK8d,[E.E=^8/@Z:+\P75T>1]AK<=C[I6cZZd]446?.
U1TbO2=40S@-af@gcF)[Z&7@I4+-I::cH\UMM5.FR:?geFd[@.HC_?LXUO#(&#6=
QZ,3EWNPd1W93JdCW4FX?YKb9SB=+Wd,Nb+HVQT8<R/ZI?F(B0&R@G/)/MLS1HLV
0b@.(Y<PC3O,I\4=D,&K)O+2WdD[dd@bHDf[a\^#V2W4bI/4G20WdJR+[FR4V?L.
0D^W#+2H<;Hf6<^;6T\B8FZR4e1.cGS0S&5F6<;Q9<C]/G+G4cS5(4fFQeb1L2c_
QX)eOU^g3=W2:0c?5BN6JcO\\6#LF780R];#HS2IMZI\2>MaW^)KP(\Z7#E]^ZCZ
=8,;.aYYE(/CTaTB5+;R0b\d?ef<MGD:VTV&a.7eaO<UIM1?&AN#1gfT-\]_3=Pe
LGfUgJeES-4L)F<;VcXS#;B>]\DV=W@#P8[BC9OX2c)@TCK9F&#8E84YPWGC18FC
IWTE.9IHLUH@@WDW+6>0a=(AV)Ad\0L#^4]0K,.V1b(NU,c8@#,.13?<7-+EY&A[
M(XP-&OF?KWUfUN?,LS=0,RO(Cdd&G835g49DR57#U(7-J])Xgeg_Y4=)HBW(T9Z
JVQS.FFCP^M.EWb?8SOL:-70557)]@XgDO7gB,;6++&:.ca98F:(V=(8E9S\)Y3g
H].^,V1J;,KLA@F#U4\&-(/R@V5[CT7&f^H)IZ9D:Z\Ia44OL<:X@=JL\QNDLaN6
G-EOV24gOE05VY:@D>R:@&>RA<#gd=L4TW_Z>.d<T=Q:gFD/JP.0;7DS3)9+6Z;7
]?M>TGK2]FCO5J6G]b5]Z7EQ:>TV6SgPQcZ,I=AcXA[G,L0SeB>ZW/,1VUS/S_6B
<PC[VAG>N/^e282UD>>Rd@bAZY:g@^4@N==GC3Ta08@/9P6fQ<58689AYYJSg9Df
4CD2dQAXQ3c\ZT@U;49&[F-B/7O2M&1[)U\4^68-DbgUMHDAg_>Z#P&-4FU/,[\T
H>O,4EU+7)bA:O<ETD97_7QHYR6@C>VUKBc3a4U2X,_7EB#YU8WB:71R^(E5BX)C
OTQ(e&QcMD[OQY->W6G&aDfA1R8f5_)Wg>,BJ;a&VWdE5eW9URG=+LP)c&6[L^D?
#B))8A#8DLR#TDfY\Z#QZB.=30KR@@cL.a6\6YP^M=85G;VP/&CJ#S:/GW?U\^-W
GGVL@8CH(-L3e[aKdF]]2_(&K#eG<.+:-)_J??4fW1E#L5f?97U\>U?WJPbE1R2P
>]OIF40QUA)V@EfP8BCMQO7e\_G6@8?F;fd=F2\I2.V2Ke7TOWfXX)IHMQ<6.X7R
IZ()Y4LPIHD_I8[,O5J_d3)OPb_9:^4P[c&Y+TbV8(e?&G[NL2a.21A<O68).TL+
5fI3\RYY)cbE::\<??dI6-H@[&4=<cfR(AOA&8XQP4;C2W[#@)d=F]8=a/3)W3#I
L/gZJ#;U:1K8PG&@f&#76fOMc\C\#,\X7f)Ra-[PU&C0D(^K250&.:^-0EfV8;D>
;6\F13fR_dGFPd;:.I;4\M27e0fG>1:9c2N5Ic_9/(VWgG;J^<)QaA+5f^27fAN_
PJc&,H)f<,U86JC69B2-_VZ]a,#69KVSO+O>dW#=[F;a>67MKOED:ZVP<b4VO6[N
dEb2Hed[f:a)-.M56<aRKR:\PfLa_[7MN)?gY;[-L\ZA<LQc?MNS(YBR&U],J_I2
a@P\Lg=9f37CN4+DSE,5=&_OSZ>g>0D_(MCUI2A@OT2#[<OBN@C5M3-[>PC3,HAe
Le8c7ZAf2P)/OK)OQ^gd]GaS?VW_4DJ[/EMa8);G>2D1TEbK4N0OT&2C5Z7O[89S
TRg^)Y=&UTCO[\^<E;KL[=B?Yf4/f]CH/BdSc](8[-U9+4D/^WS3Q1c.2^9\5_;P
T3.ac5]bF,-d(UAM#3]3[:Hf)GKGUPPEJ9B>N:+IgYb_DV.f/72:?]>X5_V<Ke./
BS6.OD5@6<_d73=I#_@YYbGRSC9C]YD,,_F?MRV.L>B2-/51ReT3Z1G]]X#M.0bD
SE2.<\cBO[4E<IMPZ5@Q,7(]S,9Y?4/H=I-=bgSH<LFc[+Y[5)c,[KUg7K8Y5GcI
#>bA/_IB+[IJeBaf:3BY]P:4HSb:8W^G\/87GM]A:+f/9QRU(cR0dV10b-Y>.Q#-
PC4D7eEQ\Cd+O;VOB[8Y@0T;)g,\ZB#-eB6.Se-5_XY-G^NU57g@;/S-HdS#b,H#
=D/E(f^V6@9Y]E@EPHG?>ZR0&e,STHc.XE6TfKb88e?5=GO0a>^U1N>G,KX7LIQK
=VXG\TXJ[5c:>2IADfB6ZI9?]NXU&H=d;B9aJ_,1-9[EQ[S8)HGJ4cVa4cO)fBf7
\&&C[C[ONcLPZ5ScMWJCQ;D^YPIB)P&ZeS69e\e6_cS47TRFN-&D&]4:\CC:AOXf
eC@^/bZO5>aO74-YeA#f1K/3eT7Y[_<H#:QWC#_<]GEQQ\2]V@:+b7N6=[fe-:Se
TP)>VGW,V,2G4d?XWJcgaMNOUI[OV).5f&&@2ZgI&.Rbb[V5.Q/dDM5]-/>>&e5.
)/@a[B=2RR>f&KU9M(Qa,f]Odb[e79.^,GB=43Y4_f])@,1COeG,N-Ib[G>Cf&G9
<1<Zf&K&EKc1b=I,@R0V/4gFY(a9Ab^f?,Z+&c[IfZHSC9G\?ADS4(PK?&\]\4[#
#b1/P3FX(C(5dKbPg(IN9@#4VHNLKM5[N8854=USIW3WQ1IN\]c+S@Y]OI(=FLB\
Z\<c7I^8L5&cE\^WKfC]<ZE(A9GQ)Q)K2?R<7TKT6#H5BA<1HW#)9[6+Jf-FYN13
U2T_&G@\.]PITKF5M[aAZSg:=SaA4;;T-:<LS@f/+\4LL=8(Z:QNd=8S]Y3>7-0B
0/FgO:H8JKf6S,2U<<;1ab1Yg_Xb.AOJH:1B57S9/+b=5D\#.\4bCdNPPD,1OJ68
5I6>?KM58b8,ae-c#OS#RSfIDB]XCIKLCEV@JaEP4ZZFZ/DC>Yd^X>QYR1f?[EAU
3[3PNAO[\LV\5D5Sd);b-F;)<)9e,:[a?N@T,-ZfWGb/JIbRT/EV_,)24]]R@a?M
3)TC@D+61AW]+Cb1TZ03PH^)N8&)ON[<#V3=?9bGOL.-?V]NA[cSATE:aKH/9R9K
)]Z#?Z2[_TH;>U7ZI>EU#C./#M9QGI>3VFA+TAZN8@+&<R^1e#eEG/8?P786?]NJ
MA2\ST&FY2;@5=7;H#4H)@^?CB-f:f9b8VFS(=g8SJ4IFCd0L#f56R3UGS&3V7Ja
D;B#KPD#@3IL)gP.DO^1MPEA)G97e3[XOeTb4dT87Q3LP]#QS#/8U-4Q/=4CcXaN
,PJ=+G5ANBb^G2O;;6UL8FVCMV1(Q8]QN;:Z.(&#<D3aRU;3#^DM?+0WI]gM)dLf
4c:LIC3\AC3a4^N#YfCBaW+<9g6QP&Z4T?<]8Y;P,cd_ZXeC6=2]T:6PcA=b80XG
B-CA6X76UdY,AL)&]BK[W#U9L[95B5DP0TDK-Ia8,^>dT8]QO5Z/7T8H3QfgNM6G
ENZ3A6Ee<KT9IKBeK>fUV.H(C831a6#]0\B(d]\3,67:V?TH)6G(b_#+,KL;)d@B
RPF_=Z2[0A>.OC=1VDM1+)c[B+EUe^2[ICa<TSYBCME>eK&7U7V0>QNdf0S317IN
2>-F:fBf=c]gQHT\<,I:?V+0:b+e1JJNVVFc8&C3F&22;I57g7<QV+:a]914QMQL
YHJZObHZW2I.A4e;cgNQX?Y]#ZT\#ULII<gC/NVLff^RZ3M9<)M8b4ADDVZOP0?W
/0ANMCL0RAR<3\_gBN5JDG.=2a[ad+7M_S?_U-a(6@IYd64P&HN[K)ARE8+(&;<T
F@dKJBSC+KBIK6OLKCXg?PB1Y1B^4HSDH;d#5#2Yc>(:N=A?P[,P<cO7<e?._=K(
9YE6d\&-aSHV#@[<cIEN&V+GbUUCgLHE2=XX0FXeRULd[K/GR;e=+EFeBJc8=KX3
d8^<6#VR^@#Ig8-\,1I;CVJ<,PA/(UdJ^/UT+1>,SSXH8G^>8A/Od8fI]RZ+K+?J
/V5SbE7ESAFcWRNV^g+3??H;B,,<>V7>2WJ7J#b7+,c[=baKT/_K]73K1^S#<E)@
<9_PJ#9S5E:LA5GWI9Ce+0;F+4WR)3H+A>[AeC1A12Hg_@NNV#@0R7^5b:BaTOI6
;8gNQd9A,-=[ZcB:)H9E/>^C+\:bRB(cT-)8D7KPQ2I8.VL4M_bcJQd<3_\8IN>G
b.IET]+4(B#/4bG6/12d775V41F<dH-.X.+;eXAf,WAbaB\]1+F5)T0gXO):>VV5
Y1E?5PYTYP&<3@HQ3=#\PZ/gA<M6[P\Z3)+dWIK+2OA9gbA6;2=^?/V2]T1^d)&.
6-+g.(QR1,VDF5.dM<82Q+B=f85UX9BTUM(CV.8^d8H3]fI?1L^7NV/FK[,Z0VcL
f]4PaGQ#5G,V1<NQ-7Q7CSN/If2(Q/#L[cFZMB>@0UB5+Z8JCMOb4K,(FGF0^Ke&
>=2I.ZEIL/]VY6(c6GU>fQ/TL8(XO?X_g(IWd:IRM-43TO.<e3:5C:LP#KdK0:6L
W67(D.XASN523ARAZ(>W7-a_G>1D]6;F,eP0C+&>F<Y&(5MT162Le]OTB28AV(ZD
,0(NJ4KB;V5K<CA&>0b.[9^1^,=.G?=^<9CRK1g;BbS.A<C_1.<Sa=L6?HKdMMa=
&0X&(G.F0L&Ib@eeg,1PNd3b<6Z]5.)=AQXS\[7X:P?UXZ/aFf_MGDUSL-+;3#T)
?PYYOAH_G06-aV5A>Z[>c?0X-D@^,Q<Z572Y>FE6@F[^ZZGD]YZG;-FEd.6:LS@^
:9>&4=RN5aW[XW.Y/9#(8ZeD0;(\]2YS,DNdQM9#:GVPNa9_N)]5JgNdP,^BO&_Z
e6Ec\.QWVS.8S0219.\DG;BPX0gb4g0bb6f=K@@#<=.=<a:a2YgJ4]4B@RUcbe^K
I#OK0Q>TP(NZOTB(UJ=CJ?OO>KJXMbJ+V2_8&\e@^V85:^5-2)@;FbN.S:0]H=28
/7K8&8fgM\Wdd<,=&+ZF8Og0L;\Oc[2gNHe\C?R90=3_D(9I/H0\fI4dXQ[//20P
+MT3_e^;7425GIIW>PVR@/ZgR=.Pb:M<a6WbTIDE#Naf=XP+TcKT<KN-[WY&U?T]
aAJC^68\/cGDYeX;+();1FcMbgYT#V894,RUG,N(CP31AgT6^aB<9.#eJD08(B9J
-Q]:K]=9Q<Rda,.eM7/HMH&>KN1@#5V1D_HPCOM;^WcG5TQ6a^7M1:^H&[_W[[28
dFZB\S+c[@D=&^9=AS<7W5Z]/<W=P3&<[AYcL[a49f08@KAQT=JC0+EO/N86=].V
_VKA#62V,eSY\)gEH1^D][>P&-SY87+>.V==78QP45CO1OKV?0X9#H.+R5^2Nc0G
JXJ4A.J12b?7OKFCN7[[c9GM<cDg6D2(YaM:JW]#EV-1g^ae)(0()EEEUU,a^C#\
P34G0=N:5(UEB:8S+4@TAgF,)DPJ)U1L9#>7L1@QJeWU@.^K;dN#>58ANa]a^,ec
fB#95c3fJC#+f7MGcdJSX/05/)[@?S0TT_I(&XO=?Y5+CE/g>M3efK&GATAQIdT5
d)GAe:1Af6Jc.d=2WBWSC:e(:EfLC\Hg;1U&TJK@VWR+-->5G\B)c[5E0SA?g)0R
?aLe.2=g45=_0YJ@>KS4G84]9_F&C60?WdV@PC&\0D5<<1V>9LGQ5UX\8<c7-:1)
C]NgDRb]1O\dAB?;VJ_H.K<bZb.O/GV4A3]1NA=ecQ?]<Yf+P^NZVYJ6&>-/g2H&
;;DeO>C;b+YC7>M?S/b)I?:NbYJ7Q[O8HY;V_]@K]>4[YSV3D,QD_?4?V--b_?a:
<P^:\M6RZKBF0.gPd180PY#N5UI@d)8U3+<aAX1>M=:0aIT:I#I1H,E7?W37ACP1
H8@e>-JaRV/.8.V5/9&M2eW83,7K]G//=]EHe&XA&SJ9<&I),R[[W.De5MNf;<5S
BF-AcS^ZcG8CQ[&22_B2]Ie7,FHR#J]7K#&@g3g-Fg120D<[O,0cR18>1Qaa&=Q/
,MbB@&C1Ne5<<QYCA:bGZE&1PfY>/;E@XVcPN/W690A45H<F^:I74,\[fH+0GJ0d
]Q\OY51L=19@G][F7_IVP^b/Y3bcaQAF2V]e?GNWI[--:#6FLE+XR.X6:>B]H>O-
c[&J&gVeaXB]&NC26PRc9P6_L8Na_dODW8_RMXP6a7AU,.[9T1P2]\AGZE<=B<;@
_)&6M)5=&B=,)\.(,TX[#Y5R6bJL>+2[+LA3Adg-F&5-M,/X)8c\A(RO47:Qe>#H
_dA]?._DU&(;ab_VQ<H6LU12BQDGWI[1\^X)[D_X42-_?>H?-Ig2[bUR8J&<H<<.
+T&]VDYJ?AY816<@H,HbB:3.(5S@Md(#;(&:JY_A]GOU>8Vb67(T[=Ra)+eB:D8>
G7(&0B#1)0bW^4Ig\@AR8C,A^>=:0\UIB8Kd03b<C3L+2/O>dB69(+FCN4///[/S
1D+K#E<^BF=L1(Z,M3?dd81[dbE9A+5<\T?Hb0]6?e.-2G&X9]G[D^=7;25^f6a9
gY6(1,:?,QgNb<bGW30<I:D#Oc,=8PI&SWYDBd5(c)>[DCRVGCPB<P,aXT,HQ.@e
:Bf-Kb6;T+&-(Ta>IHe/A(BR?e]D1O0;+2,,PLE]&X4.1bPDcIfB#-6a?69&H8aC
?eX3-7T6N,VEd-O()SC#ed;@<KUb#L)c0.N54-RZC,??/5<JSE:\U^Q;44QAQ#+G
>T)CJ:OI9Q7XDCZ^/KK:dgXS15-05(8+)6\&>L=<A_@VeVd0LS9V1D_Q&@>Y0JBT
0AJ=.:31:],2WF^@DWW&@^-3g8/D8PCcG[EVI_C3>E;9aV0N]Kf&M)fY]PFWR>SL
g61Q6_GbTCF\Hb(WIM<eI7+2Z?EPWL6B]XP+&UO7F22X?=fB.KDWWK-Q+LO/M/GJ
Ue,U.bG.WMaD8?O3T?XOHD(D.6U<3KQ,U(#>Z:A=HW=:[-f\MM?_9A9UL-Ef/A&b
f6DA:&N0P>RR:C]BW21M>[^3Ufa-gRDQGQB#=^@#<T#2O,MZ/7Z2Y58M&1).F1TX
WIRMYg)4Ug@0(\1RTS;-_ceH)E/a&L9gUJ2(/LE=OR_9eX,EYS9e-S[G;187ff<:
#4eXO?+Ca8R@DP1D(.]IM/_9d4f0@>@>)UYXaP\?2(_X+fLa^0M;W_7C)W7VgSH9
BR)W;B(bXP=XJYOWT6&_N@d\)aJKLL25_(KLfC/QV?&>_]IS)bVb-dR4/ED>Ja:/
91a(7)X5Ye6,f:B+cHCdQB,W-Oe.82]3GbA&^?8RRdF7GA;8(GNcR,W(KZQ>#D?F
d+c\fG0P98FIZF3K3>,HQC,W2eZ-K^>6Kfd&]B\=b10L_eZ.-W[fO/+gF9GMPRD0
>gS@[#ER_U5#>R>?R(Q#]5EBK#Z?,W:@d;9A6EX.ET\)=5W(^eN+@EBZK&f.BM&/
?Q.WQRc<W&U.3>CY(((Ke6\8;LLIb?H7(g5&^JJ@I)afJ.,AGfC,-+DN/+T?ab<a
a[ZA9X9<bR&HGIKVI1&@RgP[fWNHL&_1/<\g(NC+K?YII\EKeR:Bf-BQIMZ^I0:6
JQ<A2U3-:1cJRT>-\2_Q;S\Q+)W;P/YY^KOc-DQ#[D[ec+7>_cYCN/SO+K3K=UQ:
O9.CgQa(B@X@ZM^gN_D/OW0b(YaYX\BT@c-B6?W[TDd9c-9?XJ-K^0<MgK?gFfc)
#d0fIBVgST;PJK]?9&2-\E<D+5Y?5b1@CAUc5#19a-/(#=<XRf^XR/V228AIVZGJ
&C0R]VTD#XGDTE9Y;KLO^bMWL8HKYcU+\eVKP/7-LQNKV91b3+:GK)#[7/]?9QO\
^F..S@gB=C?Vb6Y?d(L7W>gca,5b_Q@]EW,.JE4+=WPBY/C3=\[<[HdOEgf0N\[L
>M0Ub[>4L]^X>L[07&a4EH#Q;S1]EIeZ8F9X2?2[R<#S)<DX0cVg/eC1?0/SaRR]
48HS]ZB8>]Z@F;1NATZL<N)61e@1)WW1E#B-f&4Q#+N#AQf<Z/(JHWNcRR<ObgCK
+6//Y,I4U6SW9/B83\,cCKHBf_[8UZYVW+&:,7C:FfO03K8?V]X&)_aXf\6c2f0L
29YRZ8<JTJCN1G2IB]\:ZI&REXg4c4GNYBNMg<S2a8g^Ab1L0079g00Z&UD)0Q6>
E6>AJ0R4Ub4@Q::DSJC1J,_(adH_fD8+XWIR@NL<8Ef):\0HJfEL&\WAB7YI1Lg)
Cg+?[/gAR^F(0-F1RgA]bGL#,+4^+ZLf+O3>\FT8\2cI2JB-eV.GFXJf/B@UMMTJ
>XS[fe;\g\d?0\QXC1IT5bF_=fKVZI,H3c]<eOTURM-45QQ&_8-DEH+6\:&#baL)
KPDS2TR6c^6D]8/Z-MPdfE(1ZXK?ZC1UFWP3I(N^0:?>FA,H\:DN5O?O<O7KJI3@
SCR91RI].7eN>,;?f&QAU>;E-4\ZRBKE^[:8B5TJaQO9./)aZ>TFY:HI8#D-]YFa
O42[6Q+5TAeU,/:;?=/.O<A]&)Mf8>S9P&PUYWL,Q+Q8EeW3d\MULZ\<\2C6=a7N
VF;W##KO1)5YeJ2a[YU<Q0Ee0M0(3Z/]@0(G65D<._Z\@HR>/@Y]bD-B[Q(V^LfH
&YHg<4Z+[J@/(Q_Q9K3C7AR,58W,;;J=,=V:Z@=(&Q&PREfEXCRPT_EUC#KBcN6U
?Qe6^VIPMN\0JHa,Ag2XANfNBA4feE-Wf_F5_dNPHZH5cW>O6C[Rc090KK;8<Qc/
IM@eC]_/R:46V]T_-Tb-FOWFPIW^<HJH>;JCHA//cQ)L-A_#=Ad&>a+-2GE8a;.O
c&18V\2?f-eY0N,FEDZ7GU1.:1Ka6K(G:aD6.=CObY7Z?+Y06?e@C+dGONQWA,@P
@;JfF&;Gg#CH);B^g<CZ;U^(SAR0?ZFVd:-,3AOE1NeGT\H6=:6CBg=4@QQ_4:P@
;7N3c)_FgP8)URWfY<#R9Y7;B,526c]FBWW01\e2fQE+A8=TP7AH#P1Z&b;?F?@M
#XBgO67LP)+Ec7fQOe1(Pc9[)4YVc6)[QE+_HV)PWa^6(CgZJ;2+W\)ZKZ0]3_V4
MCR@N_^13.2+247_[8BXR]NI0cBS;3XCQF_EHC,?cUe^I8L8W#:9N<(#/WZD>A()
L[<Q5B(]2<[J6[W>E#(AA[^:;,;,#TA^AH[G]0^aG63g;ef0^IFCKAU4@.F/ICNe
Rfa_OG_A8If^#ASCPfR]12PS,>1[6Z>aMbPJY0)Ef&ND???:^.]/U1MT4M#D^:5D
.SIf4]M7...UO3dZKfOW62bgW+T1)I2._\8g:-ZON?Uf[>9dRd9BG[JMCJ9+Z8gS
5MR(LH7,X1:WcH.45F585?abA&YZ=@J<WWfPaKYJ_?FI64OK>>c<BRg-@c[W-_,e
]059(^AGR-YKCe4=bUY\._YP&>)=SRI_IABEQ_0__2#g(C:4I@^gPF?GV=;1<63a
]RLQf?I(O2?8\@[B[]>eUR#Sa?(BIbV<#)5D.=+/QD5HG,)EHZK)IJ?K&5MYU=Q5
UD1J]TJ68bX5D;b>8H7QV7+ea#/SD;V=JD-5S6BR&V)DO&CVGT>RB@P=BQ].0WHI
MK6Y?NU^FIJeUR&5P++/BQKKFY[ZUQ13UP^[M91P@P)-FfZ^\ZHV(^V/EN8W6:@:
>M3\^;.O3T7<O#bRK3L)\XO>7SCJ>:cJUVc3F-RK(ec7@&#G&b:gba##XE@@(^9I
5/e.LTQHF_NESV:FNX57]S1DDVQAdf[ZFH1G&)bdTQS(\Z7<7(TFaJdd43e4P,^U
Y^/I(/WUY\8U>.<RA<V#]VQHe-f.O8O>DF;8YeI@PBg#N@MC\FEdNY\YDL@1#-bP
>:cE9Y]eCMD.>V^#a5aQRR_<&96B/\ZMb3Xe0#_YRN0<1dQgZS[V,KO[=K+Y)C^R
XQG(JYXb.N\H:\G@N.F:2.YC=Y?YEX+[K9]Y.W),f=B<DR<4>NMH:\L;+4-1bWS7
bbQ@e714I1AV^;/g3@4ZA;b)UZ-E\7a^I0Y^@,R>R.>QQ5)cZ3L:(+&][0SX/fg-
2C@ECE#C1L<d(b6NWffWEE)U-RJf4<c1GE9RCCBT:KDT88-BQJ/a\W4DUQ_GLW=O
2W[N7+&IO95QZVVFc[4Z/NOU?:H20g=-Tb_+HB31Xf2I9a/-D<f.K-YF5B-.b?)1
T:N_T)FT.EQ+I[P>#:2(S/WfDEVHM=XfdDBD=L-F9X^ILPY@BJfO1gA82c9gOZ50
?C5X903cM@d8R\.M??&-B+6,9g1L27,FQS_[<fbYee_0f/&,M(Fc-2\,1EW<]/_G
E>0TCKK9b]#N+@:MWcLO.&Q(TT#D,9&_OR53)NOf]+E5=\f(,PA.BU?@U^7<@;8K
P/2E<-:AA<b>BWg/#O#8MZ<^,/WGFUHC.0<)ZER^J2>7ES<EEcUe42gN;:>O4#DI
>PFceS=(LD:?F\VTHR-NJ2SaO6<KDI(Ya?.PaeE4WM38US&fL7()L^gJMBb(d@Z/
>)JEY>@,[J@6PTPVcX?ZTTgX17,4[=_I&g_HN4e@N73:=gHDBC?fPZBYN[V3C;F#
_e;.AVN=,_VS<NL6d=HYA<^^]PHX-&W:aESD(K)5W,I@A5H97\Ybg4]^.9[O\e\B
OT8WK\S<]NJPgK7eAVb8C3a\>/]Kb^;V+2F1IQGHOWe3O_,X9,=5\@T_L.7@&KST
5I#ZKSQY0\?PQeVO]8X/e+L3J-&1]Y+G9dLZFaR\;4]+?01Zg[3U0PZS8[.fBC(;
8a-6OYSPX=.5LA+1FB9\Q?g)2T//1^gd71KR[Sb8#+U]S/KOL3^A=C8C^A4J)NL4
VfTeYKAO9@c9K<Y>7?AcP^/2I@b3_J>CH&f>^>MWQ2WV14.8gH,_><483)3GPXUW
GM?0.H](>7#/HG<TBf(89N4Z)]&;g_<VX<]BJ-/Cd=FX#XCSYHJQ,>,-CH6W[aXc
EWD&_>Z^bVd/GZFP:/D5128L?F^e;I4>>SALB0&3]QgDH..ML&ZM1DIOP[[g/L26
SVNBX3^FHgE-ccLGZO-;UK30NMWV^>,&L)>f)390(RKJ.?L_D802VF3V;G1^?ccC
UZ(YFO:(FeEO:M_fXFC8(D7.CI6ed9/ebVI_FC@OcFEDFOYOb_0-bTdX\ac:;5^-
-2Oc[I:_aITVWS0W4(<B9..[?1N,d\=dRQU^#Z/,X-JfCTQ+AP#ZFTPg(6-ScPQV
<cAFV>V&ZCb@FE5V:Yd6:>GbC#^VP)2:MU23TTE_+K-RWGBaf?R24^5L;<_###<a
A:A(GM7XEQ+c02,X&.<R<_aLP++P(]H&1f2Y;N]-KV]F/#O;M:dX??2-0-/_cH0Q
P#^cf7,WE?e,XP,T>f65J-]QAE6gPg/2C&K>JB5[3UbB,WK7A^=9;-^U&CJ?H.;,
\Rg/E#/CV0PXJfVI+(5?ILKV-<6/MQ?BfcIC/?3;.-53-#BAIMG_gYB18:ETa6/d
R51aDW[[S@>B<>3>F1[Z;QG(HRHZ4@7QD#Z:KT4@LKfYLD:7769dA<Y/IO<Y?J]9
O;SMIaX-74fBW/Ed;..>A/baO(gfL,45Xd-VX>V1\[U,+1L88,#[AG+U^G@4H-VK
;=_=OB9#RX0/\,QLC;)W4+PX2g\DQ^-2+IO8C<8JfF>CE@SQKX82QEDYN#AY#F?<
CC)1^8_=Rg/NBAJ(+#UYR:a&G/gc[aCATMNM-(:K]R5IAf;SYM>=PE-<@^c@^HK^
^=QWRRB^44.]e-eFg.K5;AVW?7Q=X\RcDae#\+2d,K_R+\RGIb]#J/U3,VRK[P3[
9;]K\8/=Y61+UFe;^?L?/^?W-O)<HD,^&D6HCKAMa,)5)KK-J)TU]R?ecZ=c\?e\
)e,<BYRBJZ3E#bJE.2:-,8G[S/#41cO8E5XK^R<^1.2@S_025G/G,&=>^H(ZUFgU
+<#-0\@.3A=3+ML@.a=WH+PNNbQCMP,_@8PWB-_a75#:E43E4.Y^>6QC=c,UXR?6
BH.2L969<71N/H0+K&4_B/]S1O#dc5J)YGH^N,<=GXV9Ca=>SUUdY0DL3=WLFY_\
=0=WFADR(g/4\83A=NZ7N:PZR5NS]A0SC<4gb+?g5YV5/gbBWe)Q9^K/J?gUF63a
>Wb^-=.ca<F,5/]GfJD2+I&MG2IH.#>fP@e0ab&9g_+KY#@MMJL?cQ0V=@F#V[Ab
DXgJa/GCg_S.W7>X=?F>eNNI@e3ZC(fYBDA4c3,;/@U;5ZP[U9-I5-YP5SD--6I>
C^45cWJW^7ES/AE?VW2+YU=(4,HKF8.A&FBF2KdB&3^,78b@#6cJLRQNSP9,YfP4
gbR@5/(2LU\;>^8eRHKN_573H=ecBXbIe29A]KV:LEL6SZg?T2<QYK&^SY[c4WV:
23He2-L>C1a,LA(:5TNYNcaKVY98)8ZeS-fB[?<La?O2JSYX4,R90Ue2&M&VfcSJ
5/4a1AaYJN,??+f2e1&RZcL]<IP:HJZU\O[Q>Y)]5FObc&_G[C(+XPC?36@NJ-<Z
N?+531>ZQAKYA,BK^F4[5)T88@ONId[0L)0@SGVS>^XWQ2:V9[f5T7=DE_S6XJN#
);-?9,bSgAV:-2X8Na5KV@3256M)@[DP5]KI@&/He:2?[)]Kg/P,(1TaT6R?HK0O
3cLNQ=3D9F)U7KNN68_eXP[&O)e7UIH/gIA/.a_S,4]UCFI^VYAa:1\9^Q>\);40
B)[GX[/[ee&>Vda??#2P#T-TJNMQ^FCYAH&(bBH;cOQBG=[BeK?_\<JYf]UCEX?Y
YS,_d5Zg1N)ADHA9_Ig.\2:4/?]T1VY-4)4+:^4CZG?#D<1VS_LX@1Y-d,eD@B@.
Y3=L6T825,GagUQ,Q7d40bNd#;^fL(,WI_O;fPUJZM\:=8DR>#Xc9Q8(L7DG[<DL
@Wf>U5>+Y=McJKD7eZY)/e-\Uf^9P,E]:R,SPIS0VM^NbIgX8@?(K,=<G2WQGSM:
bJL-U;K8WJE529)5F9[?=^eg#K.Q?8T=,9<YB^UZK<N97=dJF62-Lf./KQM+KW;S
\;.TeEb5^>:_D=4180U5OE\YO#\F)W[^,_e_.99cX4B#_0F8.VVG#CW&^0/UYD8@
9YPE\&]_8\)ZUU/96:g1961abSOfU22Z)_P@NT7ccEHA0QCbY3]F,dBP[=7X4<1Y
C)#eUga)5Ge&9H8>BBL.b\9D<PMKSY.<5]:?M(L4J6c,26^_WC5W=L,d+R&CaJEA
MNL6B\_8;K>(&SF40OfF[FNb_dN:PaW5badP4\I[EZ3TUBNKc5ZTVbA2\K\4/?/E
PK7KJN8cO6B4&O07=2YbN4-?]/(&ee_.X-e@M+:CQ]gbPR7Cb8I3BWZ=RB:5Hc<Z
;P=/aHI,LP3LV+G;eGLWO.^(IL7.V8;RD=]?8P8[4([;1.OF>]6.7N)#Rd@OJ<@I
[g@2_+/A<KB+\7PHK:R>Y6g+IVDI:PT@:A8_.^^-cZ[=WFRE]@(\\Y7IcQ438L9^
2ZJ^[>ZR_6?NNFK6?4E<d70/L7GSN-]4P0@J4d>)&?I3<TT7O<)g>,CW,c@:#XEC
5(L-_P^[NNJ.-b9^(#)ZP.eN[SIYX;O99THNXc9[SgN#,.06-(5U>6:?.R#cJfd8
LI_#KFYd##/&Sa]KM-/MV&N8RBgFT/>,K>:WAULQ(L_aCP)[3:\8\b^N/0->#]TH
\[b6RDN(R6eg52N\AOXHGXM6&4NRa^f-I6DFRCG:gX9)b]M12<<c(9QO80fcJ8W=
3]I3^5FH[LV(1Q1@D3@BcNO:a^JE3;#N]=#2;cg8T#La,T?[8J0<].#?00ZLS&0:
^X?Q5O_[O(1b7aaJW-Ae/I,[\@O4):].>.2ZO@KFU0<W3V?;KX#8B+=T?@LCd]X_
e90:71>\XPe#??>Id05RR_<QEGG_H..WE3TUfGJR?-ebIR#/)GANVSV[GAF#Y1;e
J6@@g&<>>)N8VgO]1=Jg#;GU<//+ZVX,^#CM]J6W9S4.^8A,S@gePL9.U2cQCB/7
SeMc+;dT9=fR(K)cZaK2,a\MJ:LQ[>62OWE?,#U0)O;XSTI]Z,GP;e0]a&U49&\9
Dc@eEN+8<UJF6gfI280Q;&[_Y#SfJ61&,V#J-EB0M/+JF/MZ;bQF3/?[Xc5=L+\P
RL:eTGRe?LB=?]HS>/@[W+NQX^7PTAN):4ZAH,@;_gR^R=/6S<]c8_B\4UE00]YR
X;>a;7,SVO^/d\EWOOCeNE3QU^cW>=P3]Tg.[NaO#.8):^+7aZ2AA,9Hg.,EB4cb
UO)Tab^U=?3fBJ32^G4?PV<0c:;6&>)/b7PVKbIWH25N]g,0.BSW(T)cOU8C:QM^
7P6-5/\=_(S02-=OPWdY&Ff8>GF-@Z.dH+H_<^9eU_>2?XU&RcA#LV/3/_^<IKE/
@ePVPQ2_L_/>cfIbKWXZZ]9S/26c02\D(/J0gX]L6VLdC+:McAbM5a_\:#Je>YYa
+Z>D.61.QO7P]1eGBgGL=6KC9P+6Z]+e?BQ-K4YQ;0e7;DNKF&/2NQ<WBF/Udc4U
B;WJbgd@c_8GX?fSUWQVg0HYN52D>NX^6E\Gega&BT#R:CQ[Z_aGY?EYfQ_PP-0Y
02NV1.]a0U8eGE&4[8UD1TG,&O9(-Z65D-7&R[c-TM1gAS]RCC>I]FLRDHL^WHO\
L=P\9dYO#7#DOF,4&]_-AG,MFL<HC,eSf;Og=DPTT?7XSZLC?K5c>fca]7,2Z0,/
?cf@AB#NX8Gg)GZcE<M5K1;/V>J4PZ6FD9PD#20AUE[^A<#,V]Fe<LC-(,.g[V,4
#/A/88KG5\G((e(&-LV3[VR>A+>SER,TT[.WAPeZ8^_NG433_9,S/R&S6KQNg1=^
Vd__S13/<;159Q\DL#+7:)<[L,@8::H4KB]&U,bNHP+L7Z,[>JRd4RZTUE5LMLH3
/d#gFZL3g&Z[./?4;YaXaU\@4#e?_TRZ.d?GI]1HJ<UccO@__@B06OGfKQ4&Qgc,
W5EX5<,b=+\O-O+#MT1a.:PLZE6FT,VR0g8II^5O_E\_3DH5EIW(CaL;aX1?LM1a
R-Dg^LF\H:^,-CS1+/LM6@M)5[cRe#OO=7V)^5edEU1#7Y]PIa6N/R>7A<2Q:6V4
C\KP@SZURe,3fg0a5[FZ3LUeQd2)ZR1DA1[,5RSUW/<:\Vgg(HQ:1+7;,VO0D\3A
E]8>+/8\KDP+,&bJK(cY@F(LPD4ZaU&PaX9OO&;f71]^Z<If^_cK.G;Z-0@fN_K@
1K5Rb-M[<B5,9gcK8EbR)]EHCLBSc.e7\6fYf0fS=(TbGa^LQFHXH0S6MfR)Z-f@
eZ>HT8Qe5GAM)M+P1aS7CTD1LA_312)4=;9:f9NS[Q80X)BeLQC^GJYa]A\X=G]D
[MAdD_1TMf7TU>0FNc;6)aCHME21(#)#8>EC=3<P^N)S+fII\6>9e;(c_K=\/;LA
F:b/\X]4Yg+.N[-\9W(fZf[Y<Q<HR+8>WW8ICEE0M:3ZFAA1U1WWQ6aRX7(SUa]d
W9W09;4J.G>aNKHDMc>cdXLfc8=5W4+VVXf.c<_FQ3=2JWE4de(7HUK>8KHLK4>-
:IJ1#UA(-d]IE+KcT:A?70KZ&5XK.eBO;A)9=N)6>)3bSd(M.5Hd,J]?Ib0eM777
;Dbf<DQ5,W>/H+YFCdGPCcfR8bDC>WNYJ&(3gHdO@]T1\+;(6&CX4UgS[.O:(3aQ
4BC)YB:]8)780.P8@JSY,@bF&<BU#9\^2^P#7WaPX[\VRVTFKE:WG6f8<:7dI:fa
S^G#J<T-[\H>Zf@^+e7><N/<W6[16,&EYe?LC]>-G6\ddG=4V>17F1F4=5BEA=Wg
d3b;/][F\A2&AM/1B2C=O>A:1N87X<DcN2A060#.CK.A=fB>LMW_4:XHdJd7V-#/
Tfed^/)Nca]U5a(5WMZ2ISZH&3R65a?DX(3XFQ:K\(WdE4b]aY_cXGg54e(V&=e[
J>=2LI.FPa+@(g6-N-I(/e.]:<=@fM@RL)NYEC11S#DJ+W7<)?&O23@-Q-.[/E[L
@9L]UK\bGVR,1I;I7cNEU7fA\SGC(bJNNcda20(Q4KIR@@,cWQ@LW2I2/K9b^(LP
a<Y)e?S.#:&d]Z?QT>2>U4]+UbK8^W+UecCg^]T[M<T&Z1-RMM>J@>8e57g[5[=I
d6F=YDdZRT&cF(T(E2:WFB-GN&PSZYP/V=+>)\X-AEV/cafGaP5HP=H[L[FD+9U+
/a\()WRZK:>^#A]\V_)T/VfO0B)42X351;V?8H^2;V<2-_^&7_WY0N4E^g0Oga78
F]DD58>FHK(1KJ:1-7;GL><(6J]]<X,b^BVd>?[+TDFXBLaA[/L7E,TZSWCG>edB
@7^JRZGL0+](#\b]C>DGO=+#<9(d?/@Rc-8U-)Yc?&#6?0>KR5TK&^LCA.I:e.4A
HWL:d7&N7R42Z[;F6S88:G^AC1(RKQN>8CI7T/(^=#g@A.,+1Yb1/VPP9g17e=AA
X/=?#cI/1SWN,S4c<WK(-4f1DEVRX(NJe/W[J\IK#@0#Of2f,JK2>e@.FWB]8\>X
D6[;C/CQP52-UN40JeUNO45b_B=JT<(-A3dW-D8;:WQ@HX3M7/WUEOD^.f&G_:;R
?_F4Kg_MT[a,3A=b@DLNb,d=RM-SPS?fU0N8Y7_7:Xf>:XbFD[1NT7/4E5c+:IG#
F6F[CDOCC1IB1E<Gc<>ZR:.I?\bX1B^4>QL04RI/#MT&]<[QCV_17N-<NWQLd.TU
Q66[(..<#N_3.3^.)2)++QJ/8aUC.CMN-/E_d8[8Y21]:Z9&XI^I@7K9X64VEW<Q
O[<&[IVR2+>KT18EWH4492S</)^SR5E6IVMS_8BT05eT&Y(5ZM)AS36MM:MGO3@/
--Ie@B&2J7P:f>/:Z-4XA>[9,2g8I?bU6DQ4VZ&#89g-A9cFH-\T6)KCeZHM8?&G
-gGKMJO@;/bRB1JH-NI./]1>ge:#UVY^,U-A#d0e=W=b]@HeDd&\QSY;L2]<K:3+
^>[-aGFFZA0U4e6PTYbdPF-+Z0IFbc+9T>UY)8XC2/0V1]4=ZNG5I\5R6.CI73a7
(D:PDe]/T#.0N<EJ4=]1)Qc3TgO?6G1YQbWAB\X&P[(c-^7/JNEeS[>&3[UMMDc\
G6]<A@-K[d8ZB_/N/+^,#3,_NU4TDB,B=A4fK#Y,Z4WT#cVH#DJQ(+c?7SF()G\;
bFU#6T9X,@HZ7gYW)=>b/.^T3+;4f.dF\HENRcbFI/eE8K)-/N5(=NJ=9N^S:<?T
Wa1Vg]NB_bCWU8,F#BF\bP4N3,^d+CP@cIK?F&<8QQ9>X/V@6(#@L&#SG+aVQ<f2
4+&XDQ[@ADg+(I#aH2YB7JQHb;PWV)154L(B)FH&&UKcI<AR+X2,U;?>S;?5M,.[
F8MV9;]I3;O=&5/._aTW/g4A:F#,bQY5JF]LVZc#R[X](+TURYc1aa^DgL92ATS?
+C^8cBRCMYa)^X?8+JAIZdVI,ALWGRWAT0=EKWg1U-^T0[J8)6g:^IH/ZB7KV;7K
^=/,WPFALN3?@P?O#YAL[NS==d+KW,C@]BC>C.->72W90=<N)/=-+:EG@P5LXX-/
cQG7TbH0(Q-X/#B#)Ufe6#BWVcF&#(V8E=S)]W13If9TN9M-R4C39/1:AJP=:g#]
ZS6bM4F0Kfa71=K:SBP.)I=XG<?fI@[:Tb5NV7TcGBC@2,b[LWR0C-8XE9#2(T+E
6bSe2I:74I[?EBNM]1cSQMD[Zg1BgZ.DU_V,^6MEQ4J5NVE+.Dg5>O#=0<1TI7c&
W-4X+BE54@CcLT,\6Y.=#H6P2Xg\Z;M)8>M)YCd^HCN+Db\-faMX,,E:e)UOJ8@X
FOX:P)2X:Q[\c\J?ag0JKgBL9=8YQNXYRV^c>Va4&0TPfSA(+L6;aYKH=7I1[#Fe
WE0>.[I20KRCEW<,aU3[=E&Xa+BD@;=E6W4BP+N_LD?8#0@6?Zad/],BW5Y[]HNE
(aB1S?S[>;@DVC>=T<2N\A[VXV2d9fTY(1DS3R3W-?:<2D>06_>bI3B(b4ZTTES4
QDR[cB1#A/OGY;?\g&^P_PY=/8Z6U5\#(<2GZHYY07?;T3:L6W+5W0:N[0f3T<SE
Ua6f3&5baN(MHCTR0>gaG[C[#U>PUTZ?VB8><PW(If[66(P/6C;:H<NB36AgBITV
>PJ(0+?LLT<O=SIf902#.6G[RbQJ))M+\QZ4H(_&ORF-HM\5bHWM:0OT8=KA+&MD
I+EPI&O^[/^-EaNS8>.6>A?Y_6[S?^7Q2D->@JE#I6>/H3+,5-B\P;gO@T6J+8Z)
/4HW#O)/=fU/9T:ZJ5.#RW6_d-+ZS8TBWIe=&_ZU,B(#SII+cG+C(LD2T_6807bZ
C;.)g[7Q-VXY4D8J)M=BXF2I-WCZ><Yc:B88K0FFF?-/SM1d3]5U5b)T<[aF^4fQ
=gMLN7I^T7.-feK430a)H&Q_HU4UCUC5?FJR8IF0(C.O2O7(TE,.=3feCNHV4QZS
/.(.O:+_@VKa.IT?E/eBMRZB8(\SD#KF7cK(c82HVMCWD+bD,<g:-]D:L3;48U3<
41BQ6.AA+/R])_-_74/UI#3d/T3XUW.;@HOb+<68Y#1;eW.?S3.B-dWf_]QEQ_\4
--BB>Z-cH=T:/Sgb.g_,FEME_N(D0]Kc0L6d7?bPC(f&\-HAKWQe19c+P.CN689a
Ga,9,M1QK@P+IE\X5=P&Rg)/eB(L,YP#(JCE9M(G1a8G9f9AK?7aJL\:@+gcCFd]
\ORHF/_I?3\a@>E@[)[@)Z.@95Ed^L60U.@#B_(E#a[VSgg_&c\8.+(94dW20:6U
cFY;OLEcaR3FO\@[U:3,]4OZQbS48gT:?MY@RE5F9HC=81JXacFYFf.GTK&RZPV9
&[<:XE](g-g&5,5Y+11,W89D?UI+>BVfVIG?CH_G.e?Q<=PceEGTeK0d_RY2f7A<
JVK@c#RKS>PW95GSb5+6@NUC2\MXRX>+EO_Q,F,b64TObL<YTY5TJK/HN_Oa[>=Q
8BA51H8WV7b=R+c:./7U:.N8>RVQc\H3\0.)&C_NREF059[L9d4I)XfQ;:<:&bJb
dMT;f]#^1K<.?9<MT)N400bNEPT-=F4:-7_/NE<XO:(9YaR39#VCDC1I#L#&J5,Y
KV_^.7YeV.:JdTATP^RQ_1I.3[PNG.Z[X+-MeYJB:N?bZ6F+D#T&RSWKD_eWB4\^
LP:.;e>]&0O@F.ZOX8B#KQfK/F]MN0GIFfFV&<MVcEYgAB[0eZ.fDN9>9-68B-7_
ZXX1[-cW0NPCP&2QZML45c)F-^\Zb:_dH<P4I;00/cDZ3C4B:TNR9LEVFHSgA+?d
(FWF_I?W&M1FR<TbKQdI];\PG)dKZA:RX0R:_AA:FEQL01:18-=M#@E#aAI<\&Ug
>J25S8T6X1E8R=@B4JSdfC9GfQcK.@RZcUP1JVYUC>7L^[6VFO?db(;J0/1:.@4g
C@E=,<NZ=gKHcA)CK-V;+e,X[ZUK\X_4Td6>\L2PU^8C@6Dc\I3cY>(c03Le]YL2
_c^;?0@S\\HQ8gHMV&[L@9DW/b7@A7FIX?OS<M(N,/_LR206R41P\QQKA<.TN@M0
UM4FGVS2=@b\9FMfTW\O^2UdWbL?+gggU&98]aD=6AAg@3G(X<B)_M=9=>+[GZVH
GHW4#\/7?A(V#4E,QY0fNc(ELFNc2,?^aeg)]Dg+6;@J29]e7a@#)[BE^Qb^V_B@
OJg/I[>S(57N]Sa//.[&1Y0W>G3AVRaRS2^aaL.]O?M-4Ga4=DU/U;Ug)HFF0MF+
.Kc=@b]=d><(,=&O>7da\X4-X-(1RAP1;CA##=@:S/#0=,Z8g.>VgN;,].\S#Ga;
QT@^TKO9:I8V1TN,L\PX7#g8@MG8WJ9&&DN[g>+4&8Q>.fcd?&f>.\H,.+8^IcT3
5.+F^W@.,BW5Q@>HO;^2(U>4c-\SA:#Z.F\/OIf@MB]5<\KF;dST^?9.)=YMe;/3
(M_&0ddAN(#4C@JK\@WG85[&#Z_E#1Nffb-SX<gR+VLAR0E5[0:cV:,N9L^fN63C
))/>6UIgP2>Bc6aDMd5>7NAE0=/6LaYQNH1B,ZT0U4N^)PNR_JL<.EE+0_cVD[,(
CGY^18+dT8K>2;Ye[>GC/.<H[X+3Kg,A)Q^3,(KT1971[@BJ\fXE?];Y@4V6.#9g
Q#b>BZO(MeI:I<XGTXD9V;:X<TKOF(&HU@99:@dG14SYaFF??ZOD@VaEYU4T1OX9
b9Aa#&eQDLP?<5=,;&eS3^XB^I7-YD+>c9+HXN_[I3V:1,M\N>fJM?G,VfX\aHPE
]\B(&Q6_?_WVFBRAO0aIE)e1<e[GP+/(gK(\H(A_348<IT)89g:b82.+SR_Ze2P\
9+3Fe9WO@CHa#U_La_JERUX>5>0J>\8ODeD^A\=8LU[Y3([_0W?(U9c\^(U_S4R+
^ZbX;gD)33AHJa>^_>I<4H+@.^.V,R0Z[Dcf_=>CDO_6AH=QbgO0edaVdKPRO0d;
-;2ce>I.??B\9ggSVgfe7-))EN[/(L1?NKA85&[eIFT855I^^L]JZ+Tb_@:M;1XO
[3<=b3c5O6\4M]EMO^aJURLY=?9\PLQ]1CgdIO#ETI(HJc(Led0fKPVBg_V,6[GV
3)1-1)c,I[M/RB#b_FCOX8C\#U]#N&gOJV]]PeSNJH1Va?<9cZG+S;1@?8)&F/.[
b-(f]8U\HUTX,C)VRV&S)EZNfXJ@X:GAMfa25FPO/JY>SYB-M=ZM0:CRH?VFI]P\
XYa/4X7FMRb?)(R[eNe7caAaXc:,J@^JYI=+20BK]F5e].93d\0,IB2ZD#\c>,d@
,LR-8AI1E1c>LV&_HL1E.4N0A5F--Z?eN:0=b>#8YRa-a0GM5-eEE\&VDINQ&7(>
5&2_Fb.Z&bHM69Xb6B7gF>:>P?VX)5#/Tb:.dLF4Q24LE[b4#)V\1<b5</S=@]Za
c7LJ=G/U(X07H;>/>6BcF(.NaF<0L?0?T(OH4&]++fg(--?HLGI2.8&R^<_Z,.#L
-HF+d[Md2Q+:>K(-KF4&@DP5+E,JSO^0FY5b,Ibf@GcHM<e>JF2\cK=ag8?N9fdT
SfSGC:g1XD.09IPXf4O:4HRR(P@4RLIU\;+]O@H9QS9b^5;M?;(,[(:)3b<X\<86
4.3?/1MPOI^5)]0.4C_BL>Y+Q60OH<#6cFG^7#EU01_+X?^K<PWfVbbE=d[5F8^X
(=Ad=6L^2MPIY=:N20:\7/CF[ZLM:ZM(?O.O]H?1A9^cQV\XAMJ/(&;ED4OcB]Og
\>>5<DT:@aT)3#UELJU54S57U8eEXJ6d/V.^;6(&+T12.f.bF>^.3\B448F+W]g^
8P+PDKDX4EM69ALVT(M0PgBK_(0RFSK:YYGg-)T<aRe_/VI=TW63TDD>Z#)0bUZ:
W-K6JCYXK5SAQcOJ3bE@98cIQ),0X-W)J0NNY5;AcQ9F45;Ja-TQV5S=aME/>9=W
O=eW-PSSdE#OW^98Q-f?[_=B1f>4-MK;L/bXW1D\J)c6&[E]4/@JOI1Q6d?C-,Kd
TP58ZH;e)4?eLP[d=eC^QKC0]T8cA0\0897=@#CU;S/8Y#bVA_FWd^T/LNdA(Yb[
2;c<)Z>SY<)Z.cc376aVGYF7bbbAOBH(S551a?IM@gNFH_910g:(1;7&TbK5F^Yf
IOeOQ)CY>K((+XcA_E#6Pa1T9If,&e9I@c8_bUb3;_N8F.N97QST-^J?ZHHKL[^,
F4:0aX0@2&f.7?HW8He<43AaaI)dg-Z];VL6^SR7>G.0\RbJTQS-QDX;V-IeI36f
0HOY\K=Y3FGf<.@TBT-\SGFb2GS;A3PX1@2_Y#\Gad]Z@GEPPC2CT>d>D=I@6X,4
^bIMC_<:d++F;25e^?6J56QA&D#K5efD>Y(>(^g-=;W=SdWF]4FCACZ8^+/QKe9f
+^:3,Y<8M\LBEW[_2QG2<<IE2M18CJ.BILVC<I+Qc&(/8\0Oe)><VEAg&#<gE4VZ
RJ?;G/=BV36(#[&P#8-^70_&bJ+[F6--W-5>(ZV)HbCfD\]3/S3MWOUS6=PfdR38
2^-HTZI^5JC[bRAfU.e_cI.]7LL=H04CQH<U[^A+Y^J/O;WfBWY)2C[1#1[NObdf
cLdT(QeJ:(+_Y<\e\Kf,H+[c&XH/(>?J@?N=X_WLNeT#PI23c&B+=9R)P>V<?;(=
dX=fW^b_,Y)?\HQAf/:I=ZKOAG.>\I^F4&Qb-Ca&&YFYT1HSWNMSe,PQXEBF+9CN
J]0;CLI(6Ua7Z>N9af_=@(].G2dFb@g3PX:YF>EF11F,O#Y0FbZfgb61/A@fM>&=
SM:C>BA#7IY-JW?D8SMXg8O859PP6.&8;CP@=+U\0JCKW-b33\3f^SP?S8A4ac1I
W02)E@H_V)F9@e7)9[3>T74<YN<8BID=Ne0(U>#KRBJD-<+X&+W;T#1H8_cZTd2G
Cg-?4d0TM]P3(:Cd9T<.A(\?(S,:Z.Z[g8-e9[cYB@e=;=^Ga1(@G1/?3-_PL0(F
_c6ff)e5>K5#5d_>b,XJ<TDC1f(2YX6@IX<>eBOR]d_5[W-<ggZI9XeQ#F=fI)9.
E4Q?&:IdF:+a;:P#+:GPaY?A]+N(d6QD^YQ0TS+Y>F6+][>dZbCFHLO\^]W)C/Z,
.,Kb7Z.J:IR0#Uc?NQ]Ya]70DVeLQ49-XL]E0^6RV9#F0/c0K]LM+W^KcV316)SD
?f\J1_O<T/g3^QKRK+;P6LX=3R,H;T>NN1W7:86DfedW1Gd&-0+<S\Y,TGgZL+T/
K@H2_+R(=7KFgT=A+a7c#^-,bOI78;NeR9V;W44173B?PP9O1^e]GZ_.c7a,g6Sa
<3EXM0Deg+,f3&O.a)=3c1W>9/GKJF-aOT[YA:,QTUBYJcd3CB\QHb+&:Ta8LPOZ
1Q(@M_LPeY[_<_IN+0GK[86X4=QU@QgP#HgI;):8F^bOTWUU;EHQ1<M2ZUeU[3PV
cKE0Y3<L<X?f0H/D]6KR2c1fV89EF(TU#MZdf:IFZDf^SXI9.WZS\:=Hb\EDEE^B
U#H5d+MHWObdV_e7YBQ1MS&YQQWd(L<NK5;@S#AeF-FKH[MB\8<4eDB=J\d/GQcW
4&:SE7>+8Lf#4aYU\750)L=Q;8X^FC7f+)gW8c,7:EO>(+-9Pae+O,7.Z),N(99H
V=DAKG2T:E,Z.B/Ob_V92f6U_F^82FBYIEb-BfFSS]OMGKZ1=<d)f#H1PXDQT,ec
PZKCVR)<dW\;W9T)B6SfE_e[0,TO8]@(PMe&W;DL#UO[J1MeT<:E6YT\L[+6JG&@
:Q:[=dI0\G<c6\6<+F0JAYR4eH9&P2bc5X>.f/I=6XNM[1+>++GQ(,.X4RN]/TBR
5>(;@X00_6QOJ@c[C,/OR8@Q+_LdF+.ADF7F]6#YJF1:f90H1\4R-JZ,VF(>OCR:
;4bVLL92Vc#IRZ#TGZ13[DQ(f=94B>Vg58Q.V4QGb-3(2UR0W7,MF>-K>-\[Df5,
5L1>>0V:S0f;I_V1.\QOHWa&@JA9dS-AL,KTL5B,=(663bWI/6#cOSW#:f)QN?3[
,Xd4\,(PQVYHVFg[38VSZRJVdOJNZ]SJ5W+W,LM-3a45g_2cR1VHKN4O[RgKU,1U
>1fG9@LNH[(FXP0(<G[gd\.;I^^B(JB:F-F2/1CNZ38ID>,HR<;<CP:2d#I;GAT5
Ia:e555dXMCe?#=bBRM-C<aKR#cSI4CWC?R508@#?6:9>[_\NC,I,D15<JM_\<2b
N09;2CdI28D4\Z(S8H#^_[.WX)dW-7ec(g]&&/-Sc6RU<1]_V2.7[ZTY6Q2@RQVG
[V5aH7YKL0)K1_K>L6&@,<O9[_&QBIQ>MVWYX(NLKG=>^R;aUa:U05PUR^35)TW[
^RJ#f@F;1W[P(6Y_81:.PPC/MP7-O.e-e2TXU1(@5Ee8]_FL+7(KYGNXW+EB#G;6
7AW0)GM.OdX.I5:?2>D(2DSQ57[<D[S427TE+EUCKg:DG9SUB0B-YfIdVb,3L5bQ
RJMe1F#S6>ba-bL+Q.<8b7J_V:ATbYOJ2ZdDAK4-F,3;NS;HH^Z;EEGH(7^M@2BP
6Q.dA.#JB0R#;\=)\,6MW8g5^_.DGNX653:?g4+4D-fbA]]H9[TX;23L9Q?8eGIR
F>WP#M?>L\2SYc.0T?bI#g7P@<4L38&AUEB?gF:VE&F0cU-]#/8\Ne=.QCKeWN-@
T[:JR?LC4G_[1&UCP?MKUbJ^5)ZT52WZA[Ad79?)0#LU2>YC0QZ-QR59J7KD6S@/
C&N3(L<-,>3.4D:dQ^6ETecZFAKQI&0-2^g&=WdOC8cP2KS2\6aD3ddKS(.8KW[Z
E^ePZ70PX.4W35b1#]KR?2?>ac)J^-JREJ2G>\<e_S\VPDM1V\g@L@)HOXBPf(c5
#EMaVI-OgcPGHTI#QWdWAEZZ5..)I?<P_0L=;(UR#WReeeK3#0?W(Y?;ADS&8/Ne
?5a;;J_GP8QC<RebdDbQa#Q[O+X3DGQV5fD^M9T&ON-2bEaSJ7^4O>[0]42UV,V4
)O&-3E_GFG[Z\5A8CR\2d\[CX0\.H5NU=2b988TO@[9&5>bc&W=]e(H:LTG8BF0R
55aR<.XE06,Z\?MGNcXHAPQIb/[JU+2NDGF_?74E44)<NSWQ=8\d0_aA^^V>DM1M
=RZ7N.K3N;BU=-9\cSe39/W8&>eS/B,O4@Df#AT)CV5,^@0Z2BC@_Zf.JFAfVUH4
8^DKc.D(eY.4W4Q2aX=C:9Z/T-5D<RC4<5Y0c+8GSd[<RA_eEPe+QYc85^QGb2[@
4#U5,I/>b(NcfEK]A(#ZU/bTO^+-+Z]LS./Ca__L;-QXe(HUGQB4WK,5>+T&VP?_
g#Y=YOEW)[Wa@(TQ-W7=NU&W8.-PAa0^^4,L.Z@RTRA-a5Q@LZd/f?E.:5=3=e5-
=Q^13A;e7<.^UQ1bVU(d(d/G-?9]9K=T8fV)KXgA6,IYAe6::@P4U.SS8R.UB9C@
3#3.Q+A^91@R]df:37eb7@L_XD(DN@V4V5B;3f:\=S^VO-4;[JE-f<,2PZg&HCE9
gO#]^_RDI@1]@fDVeC\/VVcPRJQFLgS/^MZ6F#Gg92f:5H6/M<3YGc,<8JKZf](D
VP@J\G\F@>d.LEHFDUc2E:0B.8GME]EBT(S1A<]67K?):XBWQ/9.#,3BRR,H=<>:
5daHKTfL4,\/dM\fIE-S8S92I=UD4Y/7KP?[d;#BQQ8;?J:T1R<Z.AL@[_\-;P<.
?&G0[G,Y3@@&+QNIPecXQ(WEG>G#4UQV^B[Z#,RXPHU=)_NVL5IcB]5R4[SMS+G?
U)@cbAQ(#IUT]/Y7cMdbfcWYY.12ZR,1]ZE:/>/6bc5UI6b9?=+H56=L,(VS8c([
<C_YZNGR=[^>2[Yf51@Z?(X/>._NCc[^J]SCW9S_b:Ic=B5ZM[^TRH-UJHX._>RQ
e92D?=VTR+6BJJ?[78A/Q0fNaJ8C/B7-(DFMSIFK[M-Y#95_D5]CI;OHWe[e&d;.
R]Ia9=,E@c?Q^8EcTVFce=Fd>&S]QZE]Qg=3d:0Ae+B4<(+;SPX^J-/:26c=6C5)
S29d4Q9Gd<K]3Zc@VF/]&fe6K\G??b0dP707a/9b+\?gL5\,:K0?d2GZHE.ABdR2
=@SAV-?V]=2LS-S=/3SX[#,f7Ka.2\YFB7fa/fG+_CM94=WSIUS-g3?(EM\S^U08
/RU&8DRMABD3EKYb4EQ_)F7_X.UKO<\<8&E?STe0D.X/=<;:(N8d)\WCIBZ,Yg/@
SPZa]LP>aO2J2;&_f]I((0&SI&fN9C5fORLa6_U]@,WSacV6E.=M@+HV=QJ7>Wd?
c7?OL)9PUA.G8&d]I41VJH.6=UNW\(0D[WPQELJ+dcg+f?SbXOW6URea(BKRYR7c
Pa&LHFa+U3EQ3aFHB<XdU,3Y_NDRBd?OC1GWVHgT/E<<FGKd49g?2(.NRTOa66^J
RHd;)4>H^EL]>_OL)b/76OZ43=&:CG]>5VXg+8dLI=7RYMK^>^Wf4R(>4:6=:S+.
-Y([8W>TIE><A9.EY1Jff,[VC5N3+W]M<Yaac((_e+1H;NI2^DHeX=@CE)G/7QME
FGDU4TJAcY/9HK)&GV.d4?&]e-HOVO@AIDRG7Pb1.>43HZ_A8&VNG+^Zb-]83fHG
ePKIM]Xc\D[F5If2080B0C&57F0_5=WZ,>GSX17Z@@@(^-H6;[PcC78bRe:YYgTN
@B30&Hg,Kc0J/MYC[e,L44X-;VbVa)>1SRCe94+\HI1F9e]c,ZaJefDfcU]/)K>c
H@[&:ZOfGg?#3FG8I<7+4HQR8_]G9M;/CQ6fb(EGII?LH7\E(Q]+EedF:YJ<#;aZ
>VJ\_PC;P17Y.;X0)5BJ-&95O;e7We)PDJg;XQf[P:6Q5.3;9&3#Q3]1cL]QYFF(
(0Q0H0&/^3SfL9<-fVTY<D/>NC6HO,]2UECMTL62,#(I<Y3c>,2519I8>aAAF7/7
>G60<GJc\,b7QUJecDHFL<fU<+_,fe=ML^)ASGBcTBJLHW9ScGBGcOa^K,H9WL3O
TeEX.?E3JfHg,6(RTd7G.JYUe)CGN)1ZZFJQ1(f7IfCGg5E+.((-eU<-DTZL<Z3L
LOOEIM\dUc6&()0P.3GYNT,fU,3&5fX-DT0<P3Y&a@\JRSAfe6Q?1?:]16W@D+-_
<@7^BV=-JgPYYVQ[P+?DCKB@7@5e_X+Za\D,82gWc-];VggA2&V(Ee7E;(5]0dY.
](:WIVM:<TCVfN<=G.^;Bc^E];IEW)7/>:S]f;6Df@6RZf2+>KXWf8)XDab+HD)H
T[aRRf6LXVR,,PgG,.0,]=3X[S0G@W@Y\6O(2Z;0D^.[D9DR>CB0-E]C<.RM9+Md
+KCZDV)3+N^@,@P3-9?5@fTe1RG/_ScRK[?Sf>aP7=_(L]RPGXQbS/f)A&C1JNG[
5=1WI--Y)KFSc;WROd1^b9H^gH4T^9<78:9O<PF@G\O2L<1S@P&2CHOB9]D7-8<:
LO[Y3_dW<O@=]gEHJ-dKCb6LG\)cAZcM^TE;OTcSH(KE>\I]T7#&Ud,3<G5a+?Cg
HSZ/-0=JE1/<3V>552afUM7X+^2&#)):W+5+Y&,aUX(Ud>G>7<D54>WS4IT@C-#[
;S4NN<.N,-/V^LWL(6][1KVI4[X4D#>Nefbc\K3THMDIO(F&XU+U(OcZ+:BFc2+S
.-&[)4SJ:-aP:7B)O[]-G07,2VSU=cQX^S7YLEMNACZB]BK)E8C#R+[_.W2=ZfIZ
NO?GdE2HDEEGU=QUb07XXWQ[TQb69M[46?]S&T@YLB<2I#^Kc7@aaEKc:+)ONQ,.
#OKP10#EdWSIdJ0J8Z/?X9X2Sg05:<2L76O1.&XAH.YYP_0+cE8531#aYIPc.)P4
#SJZI1XOL<G:+_GF)32NCZ(ddg.NbVQg/2HJ>5@:IMBe3(-V:3)XP_8fU.):R^_O
=<-Y-#;Ud\EMO\e67RdD:(=D9@@;)/cX-N14Y7L4VU=,3d->3H0?EDEFLK#Tb^Nf
4/[(LJV3P,@a..(S+ZX._J^;BD]b<e\2FL+J]S?G#^36B:+c;C/N^.#g:0S(dZ:;
OU^,ANV73P6J1BR0DC=Dg\T[MU@</1ZRW>^_ES7,F@018N3JecE@:CU))AGHZbPK
5EZ/]PF(@c)-Ve_R-EQ2W>UMV/Uf9.-UHH4]JL2,M<7;H4X,EX(c_IX),S9=-K36
T[7,0^\J-S>LXCU8=(/I/RZ=WMY^5ZI4d>,\8.FAL#(0]3:30?>)PgbTH(cS1TZS
^7[-#=.^.(<?J<(VM_X#g4BY/bO5,Z8Dg.V3+a=efO.\PS9<Z(>Zc8]e)M+ML\f_
H/WA(F),C-ZAP>02aMbHKUWSOD=#WOU@)7,=FaN<95KUBU<]7b6)eQ?=CXP:FMc(
X?MN&WEN7?U(#<.W0=SP#JM:aML4PE>G2P2[gBIZXC>g68,@?+Me_/_bS::M+-0]
U:>-Y:2.cOVXC8JRc5+Z0-2TL;3c74.(aZc7@WDI[N8ZgQO.>8&2)FOF;ZW^.NS@
X2UAfZaS<..084K4)(IWb^D#:=B8+ZLbe=c;NEXRGJBB6Jbg404[][@NX;Dg]BJ6
.W>46ROJ\SAP_/ZF&^&_+,4AEVO+YX[3Sg8e_BL_)\WeR0&XTd51YMg&\7341F-^
EBVZ3^9W.XK7TO3K4=g3QCYN^]OQ@?Y3JNF?VS9=O^OMZ.XN7^NBAJ\4Z81Hg_PI
:XUM7eMO^:58YP#.\_-+5M11VW,,5Lc=RKcaHSAYZBC/#7BBPE[VJ(^.:4]Z>XY.
2^Z?(/SGKKbK-RPB<C&G]<#_09@P7UXg#0RP9,^#/AF>8V;Y,Ra5YH/&881KfcO&
ZGK=8a950./_I;=G>a[.2)1Y9bP5M+L7eFTG_]@#R=(AJMKIOY_^,3/R]F,Wb:/G
F-;bAR;OWM:P;=If5TaF51&5Yfg&5H]^>a:/TY6C1dCaTUOQ6V2IIUY=?0WdUDgA
9#AGUEFC4Y+F&C,G?U1^K-b?+#U<EN4\a#VfKD4ac)c\/NT=SBE>X/-#H-]6L7\=
UAA<H@WW8NeEc>;X7SQ&K:JRMJ[,NNLE,P24@cOSc:)5ABJMPF)cH.6FT(EA@Ld6
E]f^b0Dd5.@/?Y6QQTfcAa&20)66P=]L)X._/Qe_[D7Xb/=[E/\SSL:\bO;O8FVG
-Y\:9\@ObAeE/W),#?dU,M6e(Ie5F]4EOOD7\MF/R;Fd5BF(4GJ&?7_0U_eg(S-A
77dCPR-R(9,JJ#M#AaS;aU^]=G6T[(_+1NJB]GUMe[H[R7=B=A:F_)]#FK<5YfbE
OaUdcN]S^fR?Dc,)XDYF&_O>5VCH:YF-Y69I^WUbc5]GGUFG#R+Z6(@>#A@N][8M
>8/J:WZ;5@1\_X]MP;#GYR[Jc(E-Fd99?.5#>;+^V70D;Z=OeJ#^403=19<S:Pgd
eWZ>U7L2TdJB8Ld/H@4H(A..9_UPPYcc=ED65eb(7X6QV6(89,]Rf;PD8:g=UD/9
-T6,g82b[D)X@5V,d9U<QMWSFGe<?Jb)accRY1O)2?AJ>C2[+C9Pe#<_Ta>AF=[c
6Nf-_.-())KF)C7B^1^E[-1D^C(KSL4DD.dc7CgA05K_bY--22f56NWRg9,N6[+K
S^?;aEP)W)A[(Kd-#8b^.W)3HV:6RAT/\OQ?7W768#_Zg4a@YHE+,..8W(C1MfF5
XTY0\4cHJ2JIV,8bAZIR[OXZ.^UbQV6W+UN#b2IDF,caXaUT=aPR<AKQSH3P+JE+
+...?:Ge_81b_,8dQ#/[M]4)(NV6?9#?#.N/^f.-ZQ39eJ)?0F[-)a)DAGKb3DNa
Z11ZXG/gfe19gZG@1Q1LO<_D))=eC:AgV:[cH5&O<B/cN:RY2K.78RL(@BOHD0T(
0VJK,.?,^G?>gT40d#NJe;aV02e#KCX0gR>NMPLAC&^cZ.MMH?cJSP76<GY4=_<G
>OD^@)<>K46S29GWbUEeI[(F=0]UId6NXdK7ME,(+fb#^ab,d&^MVU^GOJ/I#Nd1
FP^E&bV]\NBZ]00^I//IBPNNcJ41/K@eM8^f3+GU=OESSb;NHFISg?W^GZ5Q6\:P
GgT7TOaFG)VUN@,GaME7RN7Vf72<-)+Ac<Q&Z2/C[QK+]N;(AYLEUdSB#P]E=aC^
\OG_\RfO2.-6IV1C88A<7BYUBg-W+4?U0g#AM>Z9^UPLcK#\]UCe(8<P(T6D>+..
.,]Q)2QY0<;ZL:SM<)R?B?;_2US/B12\6WL1&JTa+O)?-L,[H;YY1H<MF0CKS3=5
P:::fEW\MY-))LgEGD)<D-G=R<[>XSXODcQ-4f?,S990JQH.#H3M<P7Dg/c;f^21
S428,Eeg:.(-6_VU8#F21Y=#)>OacUCAD-7eU:Bf_?4Y.QYB)3_<&>2[aSRS>AY+
H_;8dJ0KXR3?]=7E0LT@+Ca_:4(2[+_IY^bfZN7UZ->R(-Sa,645P+Sgb008MS=N
c>-W=D\;_46#J/\b-H_+/P2cJ<3ZG.S1dY<0588.b0F7Q.b9CXNK82N8]V(f56)S
_;aRXNJ&Y6c7Wf]3[EXS9UD5B&:(;]I3W?@T=SB\MFc2P8<FU;RJIBYP5U)=0EOZ
UgDAb)T@K6=QM;:6\fY)<\NZ)G]\bXPV@-4#T<3ed]=6B5)A/96^L6--g@3RH?VC
<dgLdgeP<2FT&L[XA91IcdQ/EEfZ=F9O<@ad\=<<2FHMd6eXeF[I_E24PK[C(A2+
AbKBRQ,,M06e&#27/8c?#<cEPWU+EMO0K3;f.BC=@6_aUCHXMSZe5ZA8TeG3:Qf[
9ES\Zb3R=X=aOO\KI.bS1^.KeP3#_G)A_#Jf=.]:>FHJgE>0g0.-[SKR[Z;K.AT=
_>FEGedW,:=J;5Ua43fMa3>4N4E;EeME)[cIM;acMHO)Nd)I2W[-WU+EI=;c05Ye
0d>90]-cDJ>H[YUOEKN[;VG?>QJe<)@;LZZQR[W\(17:)PB>/8BN\B2<2C1DNfEJ
JaKW=NdCST=)R7#GWC6\/IcZ)(LZZ-W2I[T@[Oa+ZWbG6\0?(9(Z:F)?0EX?/ZQC
NO;,./8A,6-?6e/3^bdP69Z<6^>f\d0+SOZ>b>)(-L6^]6#<;@LVA#7:7e3IAG8>
NMSSHVFC_63[fK;HgG:K32e:#(<9FV<YBWR&CW8IMWDA>:M]g@F00X0]+Wb#F\cF
/D8c(g4AVg(KO6_J/:>X95#@JT/E<_XXULV+3D2Z&Q]L2O7^#VG73V]#FF1V@23_
0J3gQ@c23O=aAdK#5O\H)R7)9Tbe4c4DA@E7SG9LUKO0)R]4dF8a9K^4@eK50JMg
f:fTE^6Ag>++C[@K\G&740RUeEMST:a_6+Ld4G3YOMd)Hb2/+?DU82AQ+Z[@VM]=
\;W4I+aXSM6Q&Vb@N>UG<&HUbU4?Ra4QFb#\@-b=RaB@_a]?#J(-RU0GQ28[\7N8
L7GISX\RRZ9_d<&HG+\O6TK,],]c4FRa>M(fQ_.1Y2,END</Tge.gGLQ8TSK5O/d
V&>6_8b?d-eS_&9;>ZKd]5^W,EWQ-fVe9]eS^K=dYF_8<D4)+])#AOfOMbE,De6G
V,Z+D:PY@d&_;?\+g)=X/KX0#&__+YK>Z^@);S9KRDX[&P(L)3GT&CMbX?2</U4F
#V^3<Dg@WYc3D^\]U^^H1D,_R8YdPc_S=XT4AX^,a)A:\T?6SHITM9fLgf7LKHW)
YFATPg(@D?U#[DZ/R^6aZeH62;/PJOZS2ffY:&HW0TgO3SIAAa],>/>?\N:DMH;=
@bJMePV[L[DPFPKeY6UXQegTbb?(VMWXNI=:^Y2E+(G0]&Vf6TZ-_gCcf.]-1^P[
2cB>0FKTJ74IT8@0=0A.?=&U&#M<9fUYK>YRa(+&;Z/<L]?L-0GdPY5D^3S<#[.Z
WAPWORS)7I837CDJ]-)CNdBAN\_-K1CC?4FgSBRWO>SPPK-&-ALOY,,&[a&S3_[O
/EN?A=,D1NQNXOWG65]ZggTYfVF&Dcba=#=HXd<OF^J?[A]VBDL,]46=6&_a2c7A
DP[<GU]:4dB75S/LOc/M.dZe2NFWY5).O8)dMb-&7CBZR&cSQ^1WA?3MYNfa&;55
K&C&@XLHKO:3M#[F4&D4?#.A-?5B^.G]J2Fb^-SFd.7J:\f6#HV:]K\_@Q6PPVG;
?Y=4a^XVHG:gc,W+.5,[0[E:C+[4)??g2W?.X307#Y-c(&gQHdPYd^3HC80IECWD
<:VWM=P-&@7M&aN<IPN0AgeYEg]RYCTQaDXE]/]S\Q^T1f[)dCLAA27)[@A(#\7H
-/XR?dSI/TZS(:DTdP&f^8C9e1D,N?A?PP2b;#=ZN)S_T\Qd(c7]<2P,<]d20N>9
GF.H5-gMI,<JdSW3:W=I;;<X45Q-fC0Z@SEU#K_524GG@3I(L+Z@J4eLNGAU)I2:
RKSbW.YdCe1ZHXTF6XAH(CCW0;)3)Ac2#;#30A?2VBgdGff@8BV=UXe+:9:HN>Ta
#@B6=d)CB_&>g9LXJ&E@AU@L_EdIE8&Z+B,9LdARg9.@US]9g=7c[g;@9>a?V>a4
aA3MDgCJ.3A=P.?MLH&L]ER0fPT:4EI_@BVQ=DEbD#1AAA5DP.0a^8>2H_70[I(D
N[V5N/1)d3Y(D^#c6KG/R&PIBKe0(,)c#a2W<Q_OP39>4+-6g/(/-eD+AQ5]53N/
I>+ID]G7T7>Ic(5J<&C>7@/f<S4aOJZ7X?_@aX^N3MQJ6/=\D\;&D=K^14U5dQ[/
N#+-O^M8e3dc(5\HTSA[_66ge<E_APZK=aU5Ceb(9d@Te=C1\dJ>L1.ZgaB;\aTQ
JX2H_T,<AOW/bFO73AVRaNLI8^:aPaVSR5S]BBS@F\KAJfC?PPU.A]?<0.\T=.3F
aZ2AVU;;d.;W\YFF(,_8W@-SH+WM=XRA&db(a.dR1g=ECK?51K4]1@Ha@=C>08D2
NP+.&/5&Qc91bf1;KE2[c/[KdLG]5c19U/VN/5=d.dXgT<,?,/U;\g;#G+2-7IHN
2\Rf617S;1HN+]fLB-3(V:5ZHC0BK#,d28WAQ/b^-7T]Q.LgAaH]D/86,Q>[e9fA
36PCfWNU0KTBI,OX1GR?MbN?<G4d5U7XKC2GfBdB/2Ad\#bLX5@#<D-e>LF63N)L
@O#f+Cc>2[BdgG^CL8U8E6Y>2STF>E@B@6PN.KRcO@W>B(5>_<EUgY7IZ?bJ;I&2
-d8@+PAXE^EW:_DNO6=@b(db[HO;+>La.\Q?>Q&3UXFXNVeNe+G#0Xc\EZWW_P4&
H9Z9T5V802CeD3RS44;3Q^QC3&(g,K4ON[gRE9<6@LEa3Na2Wa8Qe7g..L0_AC64
=eF>6IGd;AG(KQE>/UY5\BK+8Pg#SgL5bU+W;HML>7WL+)^P8/gZRE#Qb;DbHJWP
=]63P<3NbaP,\@MaBDM7-Hc3c(:ORGDc//TTe9,MND@^11f/e)XL]cIg\1gZRMSB
G=+)fGHa^0K@49U\L_ZbEM;B0)^EENTgHdbM[TVV>I.]6U=P33)U&FE_8EN(&,6H
Y9(A:S(6U1BB@2+7ZCIUI\&e?[(Z+0J2(fEe6a.CbVG36-?ID_4XPH:N@[034Egc
WHL+\.>-f3gO)I48><HQ84H?I?K86&[7F(T7FIT57Hg:_GgWJGSZe7X5dOEOJ7HM
>I5dB^V\&JQ.65[9L[NbV=47)-X0.OSWO.PNcR[ET57V=@]3_>GOJ+c8E@eJ@:[U
:E&aa?:NB>e],aC(S_@YD[_dL<__WO-T0/gbEO06eZ?2FU^+H=5&W>SA:(AgPSc,
4>#R482S8bTXFV_7QAFKM54Y(YH:W3ZK0I??+=4P/98DX3?](&-LY[;P_bH,UTa8
V[E\.;)D>8WY4NUe>@.N/2]WS+L?VSK:+GB__9.;7HaBb0LS5TDLMRO#G8T+,#<G
LZN)BSME=.9)KK5=.)AKBP3^-;(OJ(,KO8)JFe_U.WRa+HE.Cf0=^DGUNHY3)V6+
+XMb4gZ^;2d@M-FaB=EAaAdMB?S7-2CfOPc7(,PB9X8C.4Ubdg+#>7-JNK^e\8M/
O):e9IY-d;3Y-Tg<10C]AYF/O0f5FE>#.M76e5F6/^>Zd=.3F,NX+)ee.[^I8.>^
.@,FF;E^.I4(Fd\WDP6FF4JQLVXS9bX/gT+fbLV#MAY7cf:>b,08>R##>C.&fVJ+
eR3REE34P6XUQ1<<,ZGV/f_+^^R6bNb0@74I-[3[G_<@F75[2>@)7F&JcO9X&BC[
HeGYZ2@C,)O[<+R(f^07I.CIQ7)IT-9WgV[E-_)1P13SJ@,4L&OW35RW<\T:fd):
1)KJb>#J=OU6e_Gf[.40-(+Ue<@TfgN[3SNXC2fFAKbd6NR<4.+4],Zed##=/b&A
BDQ,#P0RS>LXf84_@QP>._)P(aVbR(IV(&g2C,\;\]4C(;S&Q5BONL+GVffW5Te/
;XX.cF.0M2)3_,&6Vg5+GG[ZK/I/^UeAa3JXa[5dJO@(Vb,ZWETZ2W\CDK6J?7-F
@TT>WO#NPODA&P_V0#W+DJg^&K#XAG,U1VWfbgDCSDK2Ad))I,>T#?^NgMSG(DVB
.S7>QC]b)N-4CQe2HTW>3R7-_#.0IZOePG.a+f,,C(+U#bGKR2#81TCbVZ>JA^8.
E#NfAG[8UUHY7(4D:-0Y13;c<Da\HGdFEc@\HS0b[Z4MC2L;@I^OT5cd9;1?U^@c
Ub)d@&SAGH4>D-\HK,+AHK&UOegSXfgg,;IXZOE=9,&@K;fN:-+5L>^,b;gdQ=+U
?7R2@S&.c_HH8V)U/cG3#\:#)a)WSfcbc/H4d[,N1F=92Q=F^>fbJJ\Q.00X7KC4
<cag@Y,]9cDdTALDUXDM6G/?L\1[J#65Fc#O=SWV[[74a4N>QfAXYI2XG?[a?1A9
[DR>GMC]P2V4EL6:QB/^M1L4^+9HLe0L3[/01U?IU?(5.S9;C@/1c(Wc(fNCTEdB
I(PGL:8E?<eB]RDS<bQ4BN<\VA]T73a0eJ=VOEaAXHCe0fAW]F[44WfZ2GB8g-/N
.-XA7MZ#.dH,fJ1&fFX.81CON(:[Pe-EHU==M?N5-@eE)0=0/aS_ee5c?O7_]96#
LWGG+-@EaF<=B53YZH,3WbPA2DcAV;]-Ig-?d<[:+-,K@6_.2\B4>6TKYfc0U_N0
5NbZ@=DIAN+U]P0-Kcd=YZ@BWSCJEbd3V:5^[>S+@.MUCO2eF4eH3SY7;^dH\gL/
;74H<WC/N6VVUJ+:Gg#a:05eLED@86KYPGM2f&bN@T4#0P<@bE<[]UQT4Ja)ba=Y
XDPH#;4\:bP&C8L5ZI]<FVf9_XKJ1cO]7(YOC/Y&Acb0SED;A6)Cbc;N_W?dc,7N
I7(\b&;S#?YX=T;J&L_a?9@b34EUB2IBB=;SFH&gMK[#@?KCEO)-,cXWD9YNc688
;T8S,J5/GA7KGe-#SdeV=:#L_:-L>H/)B8;?62X;1W_d97>)?MQ_UL5Wf#NEV,LJ
4eWZ0/R/6E3F\[&L=gaR(D/N4G)J3JN-U8M0J?]T_4R??CTa\(XB6@#PRf/HV_P;
ZN1/>@U1Zg>0<=K29G,GF\]D5U2@T#1_#KPa3ZEc0(eX]:X@+HQ1X.I/#33X?)fQ
8dKbC+X&N;=_bc[\(a?.S)ZV?OE=JTO-c[dDaIb[O=H0<T:?+eL)[)Wb@1LTC:X?
I,&DCQNC]+K>^^XF4Y;EbA^b9DWF)OF&e9NHZb8/R.28KI_@+B>768EH4-L]+^T(
I0^T/OIgIQZDAIW::(LSXCdWI\;60SCQVL-V_WOaBLDA4=HZ:7-R#CfAAL=(ad-S
_..A.X,[2_YV?[gEVBP]8VM54[R<6&E48T>DF1I0H[>?5B_B\\)6Xg=e_9T5]561
@(_[^F3G>WDQBFB4[?2-#d\[\NNc/)Se93NX>^[,Ye.36F;6W7Og&CSR3,EbRYMV
I8>A3?8^MA]4eVK8D:4HI\;f^f.ReQ_fDg/N.1WANJg(,8SO)7C^F@XC@WJdO<I(
aE,\^cd<6L[C>&Z/4D0=2CI/fZ78T4=6SdMR\f0EQH0OKC0_(F6N3^(C8=-A?f>\
f+4=CK(KD)6a5PX.3([JP><F8&)];2V#C(V>Va7R]6NU;1)5T.HP30W.Q3BI(LK7
C>(QcCLRT,SFR.5WW1F]>S^9/;>)UMVbJ.K7Ia/7E1)EY\#>?Da:2](J]13aT=cH
J,J+c^BB<aR#[_<G.7FX>Y,_dS@_fB;+T7;NLXK1HKW/T76X/J2&.K&dRS82W\X[
J4UWf.=Ke6U1Va],N6/6H:-VC[O;67>V[Q8RAd:e>LU@1fO><(FR^JBR^9>DBf/#
9G6-IJZNPN_3IgL#H8\K8EPYN)g5+CaP>?1Mc;=IU)-M1MNZ[<S\1c#g/LJ9>QB[
>Y)(Q;TPe>F\>DC3aY@GaB[\#5L.P5D6)0TOa?f,DH)gUb[S9[NM(\H70#PC96-D
A[B4TS4HGEQYB@UL/-SG8#ETDZ.,6FDEY@+FRFbKYgD_HDKcbZC?^+BYdb9A/;2.
3^1TKS7^c?Q_2@J&KSQ:[-@I-93P7(,ETL#4T;#&N)Q_+C=E=>YaZ:c&2BX6C-7]
GG9M[a747g03#BKJ@;LOPQfCPW>>ecR(fbXI??Jg^5bN>W]N#2:\,OK,#RHJ@H(g
d4NIdYaaIE(<V6a8]UMZH>Hd,^V8a[\^PGF?gaA2[)ddO844)_3QJMPY@f8PDO2a
[P&Z1;[RSGGTX^DI-@TJ8#UYE>[#]gDce8+eW10;YRa)E82Q/O([Jde&Y@]bP&/_
^S=ReU,E62#[RB\9:>XB-Z(1FM/N&L&J<1[Da(1V:ZWN=L7L[TAc\<A59F;2e9Y7
b_bRE0H]3SN:Q95OV(6WHNfW\MF01;_X?8fIGT.AB5J>4+dFX\.60SXTX@Md(XWc
S-SPY]SN</ZO-X&?IB#L&J(Nf>4+-E5<#X?-WXJ=fK@5;U5gMB>gVU46O-3&\2B2
AP;U6U7(O?5W<203RMB7HH.ASMK^UXXdc7W=JU^65+0@AA4/0Ff]bLGXeO?I?a^Q
BcGCD>\[>dF&+IO([N<Nc]4f;@645^U2bGBfH4O4DfBF-)T8:+g;E./#>HI&Wd:N
@^-XW/[THF),NAO&1AMNF?X9M;8aO-/c6fe.UcQ=V\F;I)C88F?,;gaL+@9S>-C.
Y:;D(FU/+Y&fY.[6=214?GJY)=,IYP:(76N.MH2Q8HC/MI540VS[(U8d@;;GPUS6
BgDdHINd?bV_X/FH&H5L\DH]9TJA@>+@M.O?(Z1N@PE8H^_4Y8]L+R1[SU#CabeU
DQI1?,(8I_PT>Xd^J6BA??1]WGUdBT:P:D6dfd)K4/W<YbL]fQZ,<JJcXJ;A+TI@
gWU67f66B?Xc=I;I<1P;F:2PE/d&>:\5QXf6ECD>#&M86F8E/[Y[.W<(9YZWAZF9
\ZC/:e/IYXI]+f:?]5d+3e:<5RRZ/H<M&3MUL:40^GaC.dEVLc=Q/a1,T&Wgc+HT
<V\;1RLJRVGUc8_PZ&FQ[7A[.ZIN1::+7=)H5S1LRH6P>4<:1C7QCgD<\S@(7ecA
R3GW^V7:RF<FG+VD\O.93^+4+-/^Qa8dG;XW:XW4=ZgJ[S(:]2@WN;3&>[RRA5U0
.P7>A-bf#69M++E_QP1c-O:d[@R17D#8T3XYIL<6c090=R/N_HMa1AISI:d<PS1F
HKJ?)c0TfEI-AOH>,-4d8EQ3>^Q?Cbd7:NSJHV@8D[?6G&;)(7X(Hc7gPX@D3(:2
cT,H8<:XNUbADPNJcU:ZZ,Xf5#+5IaV,D]7I]=]P6]Dgb_3Yc5:=dCRIb<)\MN]b
K-^N2DN]efd]4^>8^TNUfW;Z&HZeR^=FK_1]YC-C+[g./<.gLa;Z5R&HLcQ3CdVM
.8#1(>:V.cF)1CE[f&<C.LWR&_:b^)GEGU3e\U+#QS3UJDf41#->\V#.EaGS_7aD
Qd<(0L971e2eJ]/#aCYY/TQab[8A+0Zb?5R(L:BYPB^JX&E6F@#+g;fI::FJH#f#
[E:PaIC^145<X5d0EWSWV[OFGPIc.YQ3d[Y^<.<6TG_S<fUYRZ,I5d(UC#+DPIc#
A-[[-P74b]NH&Q/2BANY/MDTZ2aDa9/C-&22Q0&f?JG<[_9(7O]=>PcRY0_(+(f7
)]d<GW?a9O1QL41>D(;;@_a@_37HEN@HJa7VO34)@2[=K425:?5Z>/OPC)XNFTQ(
/J9,OPHAZ-VeC2WaYNgQJ3c(,,.HY,NPP451]NHW8+K1;Y^-16U@E&#(OfSD(N\)
@+,-fM.d:8@2XP;&b;:VA:e&&OWNeZJGSNd9TIURHLH_N>U,PY-K7K(A6>^/_G?7
FE<c-9-@6^gaR)5)=/3dJZ21a^9Z3U/d9E?T2EeIZK9J\SOWN2SXARI(;#8fV6D;
P@\/8A\)WVFEQ)9/F-[gMT:+,#-FX#?9a\XXb&_8aDP0cB>Tb,\>ceg+=)dF:BF:
)JEeP3d4/8XeWCfC+3IQ_?\#=ge:5FF,=3#@Q,?aO1K?4_Sb3JCX;5>RRUFJDM,F
TK1\2;#[_bC?0ZF2_BH_STAZZb^8Q6Ba-bXM^DW?Od+N;b9--ZeJQ([#,9f,V>G]
bea+=OXb5(;75b+4QE92Q/IcQ]7^+[d/STSAZM<Lc4<MYGN@\6]X;Y(Tb&975SUY
BM02P+0X][0:fEY6]<3\+79a<6\X1[F>#SSXT4A:3=.?5Dd8e:8)g7N@\E+C=9)a
Ge);[_aTJEWL.ZM2\9]a+.(L;^;H]5I_IN2K8+0+QD1C?A[SZJ.<]6_Fc2P-+#A/
feF)ca6II_1?7#I)XRdQX;/dH2V@ZJVZ00^21;J+E(;WKRe6U\V09CV5\>].W4^M
UABC36OaJ&ZeFB-HD/=]TRJJaC60Vb([fbM1-eQ;g^PWIXQ797(?#<@-D(\CH=+1
UeH:\CBG?E@5V=TIOHPUVY-Y9JU7/WU<2A/@S3L;dXH1.6cTQ\?1@aY\3Id>GBA7
GBSF6cQ//Rf05K7[e[F17MT8,;A]1I)4fSYY-7#4#3#,Nc9/<#Bc[RRa>ERZWL>^
&@V[Y1D<KfG;cFUe^;W-YLH3:4bFU8^+AMP\fbA?.W,77gZ>&>XF,4KEMN7?K;P[
R[F7Y&>Ca__0^.Y4\7G[YOd.+U#gIcJH>#@^c_P<KF,cYWEa?R=92faM7)C<4CMW
]\;U[Z.4e^[Edb^D55C?-R+Fb@Gd4>aWCAYb<56>CNBY6@@Z6LI#1aU-L-F&^/DK
b()Q:7a2D,6I(CB&:?V.U>,XVSO9Aa<08e1B2NN@PDNYdUb.LOa:TP^RNL17gA(@
,D#0MWYE&]UG7XS8>Zg/W\H&D+ZFMQ-KDV?d\NR.XW;G5[2e8R0T^)?XTf.T[e?+
-EBE8NBfO)-QJ-VI#.J:50KfC]ROcCEb1U)AK+WT/dASc(>F6=0UK;0UaXQI9:+>
eY=_ZTE3S7U6ULY2-E3^MRQbLD@(O9HN2OO>aWaL2TeKX;R&8gI>eEQBZW101&<E
M?<gf_?=QRcS^D&]?87=&0OFd,+L9Z4FQ?9LEO>AS8H05SW(7f0&3\NBV[5OT[4D
eY/V=H;4X>J+Y5[Hc-FY_6f=[C2gFNHAc,f2?c;_57EG/L_,&13ag7c1K/0<>\^F
7)BIg64.&2WJ>_.OT;Bca1L1?N/fB8SH>f)>8-X=T\0J=LA8</eAc5cbTC#II)QQ
PKOcMFf)MRaPe_K]dJ8@F#.e\R[D18fUIP;F#E4#)J0fJHZCI2OX#Q#O)&5-^N?<
V?\N39SCALH=4O8D]1Q](\]RR9c7+<16I=Z,C0)+O28f[@d.O6fV2;DYIWADbW?d
R=,P3cY2#N1UM\Z521TegOR>M9Z)L,B9530cU0?3LBV_O,DM;3.?98FG<-dW;deS
;31.5(99ZDT=UE:^;TG4#R,.Z>@gB/)Y6TW)gZXe<PcMVg-=GO4A\@3Db?:GYJ@c
5QGYg^SJU4@aYPGQZ@D2O(@JV5>cSU)&6]5,/ZS?IU17a39eQ;..G^X/;J\cF\Dd
H^bZ#<eO4&92G&&<Q?NgF1S85I@3H]A9VcDJ[XV\X12cF4OQH/+5b4fF<:7:.>7S
G9H25FDG9=@Z9A+2>[C_C;I0>^@D&,K):_JRBCfgQgQ]6)9+G;3^4/EJ.^9V-]_;
]fVD-W/-AS@(I1C&TeU11&Xegb,,VE<Y@#e5V^F-WT.P]?C;32A&VQWV.;_D3TY-
\R6/;bOaIfGU/H8Rb,b9+FEZV>)&GNYFBTg/bfb0Ia8QNQYd@=)=1?Ie/fa_JMWJ
QOO?0FA?N^/5+=7N,N?R;aRg?Z-1(V:2FBB5Md0[U:Y>;/99#D2dA[R/ce;5e2\&
VX3dH0Wd8^G[VCa\B;C,@XX84)<TeZSDg\S9bS+b#/J)FaK<4SM[EP8.#;0RSA-\
Af/(>)0UZbMOWb6;/)NMCCR;\BYSb9_@1<a>I5g_QJEHQJ(#O4T=SbGE9?1QO0eP
T>NaaS>b0Z3dc)?PYI2cX[3PM;F/FK>VL@dI5>VegP8-TFW.0_d[XL-c+aCb&QK[
?EMJ4a>GWI&)Y3[HdQ=W(L<,bd.=(&Gc9Yc/&A./a(LHa)J\E9B[f.[DG8_20>Q_
<=\4e(5,/cZPd-,<2A>Z0)YKBTf52(#]<?/^[?29G4RXFYT;:C,2&@F>I2H<+&eL
eT]/)-\c[#5C^=04eXHQ7?E,3Da:1I0f/^e_Ca><&3((\Nd#M\)KMa<eKe=eM#3N
c:Q)]QGPU^JB:fQ)32M-?;@PL0BfD6Ma)gQ/GHT4<7KCYC5YK,0VI&e)Q0,A4Ha@
<-Qd0+873<.R:\HDb.8G?KVUfJBZF?J(ZKFUFU&Eg(-cA#?^CR69OF>?A2b/V[ga
:O?JGHDCEE@eg<a\VU(^WKQ#\N@?D8T>-^aTJa19Y]3<PA#_-;O[7g-8VEKScYQ4
6X?F)(N@Y49K\L;=Qb]23/T[Z4g106f6#13&#0AVT\2DD&4712018DY)KO^T/@R3
@AF[b0]@3YW3#Y1;R+1aH&.1C;Te7@GdZ?,>>]WL<Q9ENCc=MgcE#8gRL#H-\a^R
U_:I9TKS+/JOKTTUJ)<R_QQ;CC5gL:gU0N1\O:>WN\e(7_<S-a4Wa_cb1)]M40.B
(3E_7RJX[dNJ(<4,7Z?B/Tbd8;I=:7T4f-;)&4S2H;G@Z\G)&9PYW6ZALP0G.^71
QGb[0MbgBT#3LJZ3ZS-b7UFeL<bOL+JI=,C.a3Qccc]CP_-#XL&=f-EU_D4dD^PJ
,7:>Rf>A0[80?(@0_Ve-[XAAOYB?D@LEU0?HMHAAS4g<1:B2EWX/#>2[YdN#WTM0
[LR<KB9-21^8ESH[DZ\a[?R8_RD5WKQAAS(B+/aO51K#4:4G^9PDND1Y<3CbT3T.
b7?Mc)((@UN:E]JB^3b=B&L&W](HK6@g#T<_@aJ8:S^D&FD+5TR3+R-_@;AHH(,V
P\aD7<EW,[N5g6MV6<E\\=eJ4VB/)&<G,G(XNg\&Lf<GQBKOKEA,OR?W_=JP:(PP
](KEdHHBLZP<.-HSLcG=\ZSgedX#@H,BgS]/2a31O^([Ta2\(C##&]S[a50XC,eE
FcCGL5B>\FD:aUSaB;M++0X<:?e:N__F->OZ7?>(>[B#=ed-M3,XQ0F,DB12dT(^
dA_d333B_PFFK,M;dB.G(]?J&^-Z.FW,C+c<;S:UBJW3@aYB+.WB4CCLER3f7-AB
g(bPKW.9ad;RY=[Nc)^aFfI(CTSAEXGMVF&-(:5P:R+S/Ga5Keg-F82cL3@&7#46
QeEC=MZ1/EJY5^X7.3.2(9/4QH\3T@@g+_c_@\91g3VBHfd@5N1@/X7W5:^NC62<
PIfU).c;aU(?aH5WI.+XVH9G(X3-5I3g2Yg-6bI,3=gcIUU4U)\W9JI8:bcF=2A4
<d0>@FE6^f&\;b28DW>L>e57Q3V-Y]c6DgV^_D\+^57-PO\>##WGE.QQ?BXFDGbF
4I-YIHT)H:79>XMSF@gQ,U>1f=-\dQ?)Sf,+768(T_S\K)NfV#Zc-,\92?5)XZ#:
;(^Z:\XH[#YOf22URMO)VB[Z9[:3)TN67HM4dXVIg6(d0IZCW-_/LRQ>cgP&/K^g
,5<O#CR,.5::082NHb/N?O)^8^]PJBJ]3<?C?]#JP5KX<+AB?B5>-VXBeD7HB2(&
0:S;AO4B#60RUV.5IW:=.C<[eY7:/d6X@+#0NIN<HX3AcV\?J[Z.Q)4]M-PbNM/T
<77.;f9Te4_P[#&6M^WABO81PJU-+HH:DBbGa/&fHSY0YHLC\@;5C,Paa\dONdd_
&Y9J>4cbYGK.^I2PO6aCWCg,S/+H_XDFQR2Z^]@&G/56->:f>WbS/)P.H4K21[U9
=V@6H:XBc8-<Q,9)+_UC_S-]MB+_;O/cVZ^NJE8T6\PWY\29TXM\PbAM#(a,_2SQ
,P3@g8-AD?)++ET>G,N+2>2&7D((c)>4TGX:7f#L#4V4:XQLfC(Y]48YVN/\,Y4,
9BU@J9F.;=CJN1FGQRc)JbDA&&_0XCg:8,KbQ#VA16dBI)M/B@19<7FK=G^.6:Pc
@MU?<&B<?b6/+&VZKeMU/#;L/-d^1?f^[9\OgT-cbGMQ;aRUJQ>:VE3.4]KfJ<cE
gLf9O>1KA/.b-[]1&:bS:fNF6TB5+:[_B>7[RR.([\@WbIgc4BV#(gI,B)4<fNaS
25V&_+EZCM;0dK19=5CY@94)\08BBdZ0eMcg^ESd=)CbD_4_>W]4@KT=A7(-K,Oe
E=)+0W3DF/.WBPZ8L(4_7Z9R(]g.OIf<Z&Q\+Ac<OD[72->X]\+a?J0]<:VCA?1K
dUO?[_8Gb2OcIT[&a5IC;1U+4Uf:M7EL^+#@S)[X[4_K)7,GJ)31M(8(S.JfJTF[
]4X6K79RP70/a]QBS3a^W&b+8P&4),[&@,H<L0:M2VVOaSE1(QG:G;Z0a3JJ[XBI
<B6[&Ca4e_4Ob[:ZC/aaH(;JJebO7VSA[_CHLJJU[FdgcXE7F02b7OBd[g#Wf.d4
d_EJ4O@d:cMJd;P3XRI#=X@c7:?>R.0Z-;-bgB59A,49S@Z;dA/>a4AI;bb#I.P@
E?B6&+CL>FebL<aV^EG>NRH,5aX6dT1IJ5-SM<gU/BK2TDA#CXb-J+D:-KJS[3V+
X4aCU5cg6CE;G&^E/DC^O)a9OS.L_g?S]7#TRaEdJ0/BE5bT)N0LJP;/[:07,@8[
3D>:5K8Ta50ag._eBQO0#gaPW<:(fREL_<1P,N88UaG<BfNb61Me(=e+IS.b0=Ca
B2bd\V]/\/M:QbW5gUB?3]B@c70;Q,dMRaPJ+R_9V=407B^.d\H^6AaQ>7F]TYd-
,TTNG5:MA2e0DD=f41@LL-Nc1Z4U;e?I_QaZ)-KO<F(-Uc2C^HP#M];(gM[OX,P-
V:Cf?&g/YNVg3,)3;fZc.e;E;L;)ZJTWM=MUg2P:[688^WAS0NI9J[YYL(H4Z2?9
IXgGD.gF>,e4+C^QAUFY84>YWL=4eN0.7EJ[#F3[\;:)JXOH,^/YCL6#[dI[a:(<
GR6DM5J[aK-,TB3;[M/SHAH.=R?6bKX0&_+Z7;R/9NM=K3]AB4<\A>T4c[VZ^ZPM
#-89>A:C=_[9@eQT(I9D@-83aRAP4ZI@b\4\PdJ7K)M4J-G[b+1]]1FBEXD]fc#0
KCEPGJ?KEG::T9]OKc=.,?4WWD5EY[I;2,#\B&G/?9]U5E-92,B)fd+N&4a4(V;Z
^9eB\aGKLB;=+T;-+aZ77M<IHXC\1BHZ;WS./;RVYS+ZW-[;3aa&V;g:7_D2KgK>
9Y.>\O5?HUX>.U-)B[Sc<9EJ_DBU,116IX[.K^>?N@7;XZd&N(#baMTM=O>Ae_c[
fa9>HLI&<8;8P(3>SW00b=@JJ7\N)PVT,ReV[(?3V;;>=>Y0ARZ3ZH#fMa/V18[K
)[,<.-B[SKbZ0C.ZU5f/T4U9TV&cPPcL3^B#5?.\M+X>.GQ]bEZ.gT<.O\E_79\]
cA2(Q7]A\PQ^CYZNLc0^=.3]d4QfSe]16FV;DGH1(_>=#1g-C?;g8M&b\<V6=<dQ
=CV#PTZ1MgBa:+V5UJB[BWH,CYXcOR)\WL/T/RCCC;H7IeSaW02gg>Z.E]PHZNd_
5S.\5YI-:8I,OA8P.4+5DH-LHLdKX0gg=YQU=NNS,H_b:IN1HaO(-@,f@\D2Z7J=
4aNPQ)PE>aNJ>8Ha<cfB5AW..#ZK;M,K_&D8YBUZ_M#GQTT2&eEMB0TZ]Yf[XEIO
&ZE6b&1,<[+N\:<=:2FC]H(ZgCOR+Fd+4eW3?)1,U.JH3^f1E?]U6+b^FTJ&0AC_
+3\Z&Z#(?9HS^4(_Q0XM/X2dd3dEKG,E+UW5LZcZCLI#cZeL&.fI)Yg7NNW92Igc
N,WBXUZXBeJ6F&gFW6ER=&g0&L/4U0HLGQG/CA_cS6R.>79J=):,-S[f1_8f2D;I
dM_.)N[UD7T>115WE72:c1Z=N[);d\A6).A9>&;YMb2UGHVD?YIHRSde&X)ZKO3^
CNU(E@+<V6V-=P50KO;Z#&BUO:;Ve:Z+7Q+cZ#G\684g7-_0Va(Tcd;M^6[A0+LC
EIE_b?J848OU<RZG+:.d19XM3#PdB?;;Q6N^RUbQ>&D8-5+6^C/F]Y][K+07B+TE
5DJ#_<>Z^;+O]7IO<Q^fVSdI>N8\9-LSR+JUR&J\6KZW2>8B0GfLPKWe>JZ+PO(E
Z#S0cB:(=R7-2UP+UA:PeQT<-I3cH;U_<IM;ABc&5[+]\Waa5.G.TL.,fE<a7_-H
d4>U95?e@#9J2GAf?f(M?W+ZGLc3K[?Z7IILd1L(AcR5<:)fgUI,^XDH(>LW5a@F
[PI\ZX2:^W,J2@>6Y:ZXG^77.;(E>c?:5Z5@[73NO^<dJL1E^AZ(#O/ARV)Q,45d
e7ZGN;>8,DXCLK534A>KE+5&LYL-R)X4RZ,OD?fcO)<gge1HRdY0H(32e@</1LY[
OYF1IcdW(DX@c6AK;I7+V;38fOaF:GYZ<XIdDP1B?O&DQQF9BF>+@1d00SYZL50H
c_E339I>K,T_[cF<0J.864:>>:4M3Q^;?7-5;#RPI8Oa2+BGLSYE447UY:beO(1+
=<+/T)LaIW.IJYZL7508)BNOQ:>>,aE8\0Q_,f@N1\Z<\:)Z/8/6;CB+&]KKZ)\O
b2c-KCb38S4QR(b2,<K_/9?AHeI4>T>E[=Gc)431P3N#FFD0KO=>O^&T&J)HHg4@
;d^L_^+dV7cU-R2>a5MYBJ<==D>c1f.A)+F1#UPaLcZ/4)IC-7&2ULN/bGA3RQ]O
M8J/X/CN58C:F6&6,b[?G>-6W.57RRR_=4-KbM<M#1bD)G1_&W]g[U[-9./YU^9g
)ZKd+?[_\,aOC]K^b.K,CC2C.1dD8WfLX\D49O;A0X]g\a@.6>^3\KH8&X0D\Edc
+(XB1VLA_@+fbb(7D3YZbD;>YTA11UP?\;+7M[X1B#6Of=P63eKaZ5(-5He4=.#6
)/6Yb,?M^)U;R:c&Q;N=MJZOEI\]ffD8f^D3gA?C,_346g,1Z8-AeFIMPC86Q]g\
ADA:Lg<U;S&C@_<c=B2W-Q\>+-@4),TK^4JWWa0-H^>+^ddSKG.HS_[XVIW[;E#G
#(IN;-XOHZVN\N@QPDD[cb@7LgLQZb<;OOcSYBBJ8Wd)E8,YKPYcTO2+Q72fVS75
_SBEN,\9YWP+^fM^U)1]=PaPCaEMa(::WC4<+B4A_#;CfX&NKW-K?aAf181QKXG,
_aH[]X3@?c(<U^NV1G[Y@\Da.58T=32e>#,N,J0X&C)3IGRY5H:#d&S8-8bAR.Y+
\K\G\>611.&/JRU+V3@X22(Z)WX-XB<4QbY3b.c8eL(9>WQ=FdR\PcbD<XB@-URA
cHPK)KAX/)ff70eEIFC;GP.V-?,6cPaS^;c.3aR4@WQ/4f3+A<@+IebZO:P)\;G(
+-Pg7U<P)7P1<ACfI+QR7YGg/NXIdbYQS#7-BK,G1H[1YdW)g:[R,B@\E=C#7<5]
,_;HD8aU7Q08-NLQ:[MSD@Id4e7.aEJ7\I\-@H4BAL.^GUd.H[-c]_NFa7M#aF=S
6)C9g9+aXJ43Z,EQcfG\];\\L<+&8f/TJI<a3<7RZ7R,gY);VD4R^MfQWF]7LM=A
]=;=?#03;Y:Q9MDQ>af2Q?E9BPS[TUIgfUb(GYH=-EFLI_;=\8^OD(ZEWbG=BgY@
,=BO:8#V>GF6fb8K9NdEb40Qe?Z#UZcH3(G]-_)^.KFQ#3CH;=d0c+P=7C=)00GU
g0;N<4gX<?X^NU2bG:9e5ANd(PfP_\C,R?HVffb\Bf_e/)E>7_0QI^L?HXA&D5b-
C@AbSFMcL1JBJK4<4:F/7/8G<3W,Qba1F,A<J&Rf0/cGBT5ZF637Tf54/&LRZfgc
[P:Fa@A<^KY+K.HWH1/N=(/Q,^Q7[_H[-\:E^_#8:A#e9Ne?/@5Z.6^cZaMc.YH9
,&FA]L#M(^VV#7aa3Na8dd#G6Z0+a8DI6A((8B#\7)Y@DC&aA_(,K)]A=@IC>#,J
bc@B=:Se0F]0,##./2]:_YUgE5_I[TZO>2TB,-0X2ED\D5GQe.?aCIg[bSEgQD-f
0Ge8V[9]Wc==K^CBA(_GT,ceW8P=Cb-aPT5LGP\IIZ1<L7eTZ/?K(d:+OW>3R+&\
Od=)(^C0#5eJM=D.QE#J7Z/7X;ZT51ASCd_dKRS=WXMJ-+^,.#O-)-9:45S=(-C1
3XF6W8Q\+=]WDXK7;c28KEL3Z1agW:;MH+b1TH\<RgTS>>(+WPFVLB-AfUO==^;1
4-6;]Se#_5W^bY26fWJU_7+=R[Z#aYIM6Q):Q<gH&0/aL(.+FG<If:QD1=D2Z)7\
4+()@a_S:6B@O@[CB?THI>IE\>BKRQZd+[URPSC0,GfWdD[=A+N=a<(J[H-C/)XG
=_H#J0GFG,]6:DW@TaX\&Y7Ce=#Jc8@bL@>).=[^-EWJCQQ9EAO,]MZ.:J+0IH;e
-gMFI[SY07+Q38LIB]NDYd>4YP0@)A0F,S7^&5PVM;1SDP0.6TM;^5SP#O#)?29L
U:ILAZED[gKaUc-=Q=]UcA5K>?YR<dA?[7T.P-BMBPaP?KT79U(-:F4MY+Z,M-BX
eFHEef^&=VIY^P[GgR+fc+Ie0_X\7>[N;QFaNQd^\C>@.#cV>,Qa@ETfLGK);Z,[
5Wd(T:803OBV2f?e)JM59adR5]<_BcTV8,:DC,^M=IU6PG6EQW&DcT-3>Q#VbCZJ
Tf#PX\R9>UBT2K_<(G1UV1DP>6c[Ia-GEA]VAF0&--g[ME+E-cL<&bV)8DS0;YTf
(><]_XO;cgc===<(6VF6\)CG]1YK\WDIdf5:4K=aV;KEDEgeED1Mf#g3[(>FOY_T
EY6.&0MPfC(OdU#:]W:YKV@2^0HR.E@0b<85<4SJ^C8[V+U4EOE=L0RJV(Q7cB-G
1^6^LTWEb-_2N=@:BcT)A#Y52EU4aD+,g64Y-#L)CJCT6d<,FY/,dVZ:0/;]O]6C
V?d]HaH2f)C7_F+>3+IY#<\g(JK)2/E&F0?Z.AF2]H=]_Y85OTaVL55Q()fORQg+
-AKG&>9MPR&,)BaL>S<CUS(ASW4c;CKV3Gd2BA>@<ED+<)2a_9LSQ.^@N,SAfe:8
.^XFXU2P#RWOCE3V@51QMEBCXA;VXVSY-Z14.<gUNKR8N9;bVR6KX2DX/c6MQ/S#
V5\T^,ffO++c0M&&QJT1KM+\(KL5/@L+P3:Y:g1Lb&>9R^Q:T)ag?b?ONRNR\BPK
7^\J_1C<DIBF]bMZ3&V-38NKa,2?[V,KC&#1IOe\NP\X9GU2gc2G(?.-58.7JWUb
F-O[5ZbD?X,0)=SOMX=KZ1XN93c>>]BW:gf&/Ge1F4C\/+J(T@4_84NPBUAL+F54
@T+RXY,1@,9]&@>AZCJ<9@DRG[[_9@KL?9e;6)EbX,U8S_]))365Q+OYI7V;P6G@
-]P?Af.@\\Q7-EX[E1JI2MebX+O+7/W\RXZR^DbOZ?WFDL<Z?0Vc=3)A2P>&WF5H
YF/K>R/O\&1c51+/RcGVb.+C0XR+.JfOOY-#SE]abdeIFO;S&6dL]0gbBT.5(1_B
SZdDEb3CQ&KN?/R(^YbC+aeH;>F/SKL1/)PB?Y)B+c31bO#BQTC=I2/EY7a47:L/
OO^Ab)E^HVD5&9D_WQ:2c#NQdZNX,B9>X+]8P85>b^Z&:2O)MXSSBU&_S7;W7C3^
>Zf-2^Ve&<.ILL6ZN]&:XWY6<J>T9,H]#fabY]K[J:#?JUYMCY9>XH6ENF7Cdb0^
0d>[B(/IT7\_eA@E_18DDKB4WG=5EFE))S=R+Ccf&2f0=X:fG7dD68aRB_VP?Q;(
HO?^EY>TO&-?D=IbfN:]K/Ye@W?>2]&BUEZ&I3+RQM64P,UXCZ,8JNIHCB4]3bCB
G[[7a>71FaeTB?O6BYYBeQ4M[[?.831)N,)S=(aIEEPMGb<P9VbO5]MOc68=E96R
9.HWUYg1_ad]Zg9Kb4@EKM1):eQ^(+S30dG2?dFY?OK9,f,2>_UXAKF;fTD@aR.b
^gUGXW47aId0b:TbQdDH_1/T#)R)L)Ye)R:NdGY1(#,GETe\Y7;dXEa3Sbf\]BD0
&R?G]B@_3bH&CQ+MVMUT4NFeZ_0?Q5@=I=C-Z8(_d6M;&I/:\6JeG)=F?8KQa8P6
SO4cfOf#FE#D3bY[D\FY)FP[0#<YDU0U]O)b3e]?dW7af9<Ya,_0+&aW4E\8F^EJ
9UcIHKKGg2ZQ#Y@,-_MS^G^DP]Dd2JRA3FE:bCDdK)QNA&c+C_bPXWVBVJEbMUXW
gXdGU#aJKfaBZSMS4c0A>C@KX;e.RLI>OU3cMIHG<RU\POPY5LOfKT^\If4RG,Za
S6e1]WKd0)&C9\SR5aaM,33JLZ(#4=T0e1T(fTF3#Q#JNR7FECSCAcQ-_ANJNM4R
/YX-H?_O;]f1/\Qb6AE3QML;&R=I/KZHeY9B#QC.S3?HW+]G:ITG?J:Z<IDZLU,>
X<:Y\gYL#=a[7df1U<_2Adb/.CNNg?(bAIVg6TcH[^D\>,).dU,:URP>\B6\T8OB
CQCPf[FP^0OSI^bF6L\1=/:,^1dXC.<U,,B_9TE?316;e+a9b(N-cY9V14GL7,9f
d<)SdN9T0\-bBIG6IBGeENXD<)aW8=P:WVO0AI^V/e1(UMKX/8eK@R\[S>C=gDJe
P2&))Ab7(P?0G1(E_9(?Ad/<cYK)A?cY+Wg-c>Z?&c_]a&0,FZ>>eYKEZ.5Ncc5g
4;@K+CcV9]&S.>HAU_a]5,N?8:AO7D1MDF(&M/>=+OWW(daX<BJS>b<g^-8A5-9(
Y&a1ZUI^#eYN<F7UJ?7BOG;/3Ba00YN=K8f5,>@DF^IO1A-_.](9/J.M38Ue_aW9
5c+W6a.LfHS,V./17,1U^+\HEg:(\9_L.KJH:L0FCM3QH>X;E0QJI/Y3QGb7aEL7
;1\==E;ITFQG5gAaW?c[01U^9@ZR;FX^>VCSDG]gR5[K<GV#,[bA]M/H<X1#_</0
)R8B7(]]#Be=,UZKa.2Id[c]JW8;03g0OfZU#.De5]Af+[B-J15C4SBd[EIS\W2g
C:IeaWe#-aGEg_]XR6+40<,bQ4c_O.:&g)1X2_LV5_TR3.QKNTJ2?IZ;HY#R6Y>c
J>.[?G4EZJ-/Q?24c9L1M)1P&3G^-a4\3B>=P.cI[:Z0,[7G&-798Od;^8:Q:@6?
HE=JUeY=Kf2=cBH#_6)_0Y9=8E1G?X?5]_^RZ:<.dTHdB+I+cOOVDX6>9Df:R(1e
K;F.X<46Pe0-#1a4]JHH0a(-BJ14R5SH>:4JdXUbJYN;2[/UOD_8<EZ\-J^G[+2?
c&K0IP)\O5:Xe>6OY)/N6feZ.E+@KX>ae1\C=RMDXZ+D<V@[2Z5b/e\<)5b-3ZV@
;Ha17UM4_APIK]]O&A]IN:Ab1JSA^E]U=R?1B+FJJf4:?P^(C_7?d7RHKD^gHDeA
QXCF7RVHaF7/(OC+?-3GK?O]A8H1GT-M]56YCTW-9S=],,0J@/V:(GEB>K2-X=^7
cM&Zcg0(HE[Ad8?8,:POH#/Q1J.1VW1^[T@9A:gJPLD)>Q)OdJVY:?d\(L#dNP:S
H#g/L=\TEL&(/].GD]Q)ZA]8[Z0KRKYF\@)59F=W9;-[0Q?5T2R(?1:=_/S3-7O]
&FI-Z]=E6G1A<.1Ca;[D)2BF&d+F&R[-<1PH5SAG13,PN7ZO[_S.\50)gM)g_8XH
EWA3(7gT?S,_B52SeC=SI,<#KH=^PM:@R:(3\NDAOBKF-./TADcPNe,QaaX1=D&H
3YaKFEdP<d?1Md[D@XUH8;FDAXA[>_fR=IdDcdI0?_)X_4VfO-)A?H^,^(]2W1_H
V6H7+1>a_[O(4/:;<?8[-&/E,UGU-180NBGHY4_S1dK2.+GEG#CSK9:SKU-LDGRQ
40c_a-/;WX9LO#:bWf5SZ3_)e8Z]O&>[#JT1ZU-UZGgaV,@:;JRP#S<+BD#21[dX
#Q[/6Ob?AQHSJG:A4CeE/g>3B>#,PKcQ&K,:L,@XR9H?O?<L_a2O7f.+FW7\;(@)
^.a>&PgVgO52MDZf\.D^;@0a[O2e1WGH4Y5YO>QO>6@C6d0UQ<,cFD)d-F2,9;QP
YWJWb)EgcFN?YLQHF9J/V\YK:,-I=LHXd?[7/44;dW.6R:G7@T6+ATCB[AY7G9:e
4[-25Z7[386?1A6N)KHO/Y(:PE+9>]8WE=/g+FT[D+d?7,F9N;7-5A/I5cJ<SM_]
ZBEQfCPLJ>VQ.TB^^OIHY<b@OM2_CZc2caK8\Wd_ZQSAD#V:5UE>SdM[/0KRb98L
E6Pb2QK5,/:+X))8>GS[#,)8Mad5;N,T98?IQ+]G=+6\JG5__dFa9?>.a/6MNWNP
fZEf]R/1;[;T>_OF?,ILEOYPcTK:>d,KWM:A.;W<fe=J6HZ9(,Fb(9)OdX3WTK6(
SD77K\A:5E?MDI?F425S;PC8N[K5)6QU8(BKcP6<&E/Z;],0[;TIJ.HW_G-<3VE#
V=W_3a0H<P/EdITd5dVVGWfAQ/PcdQ5;A\M^#F3G^YGZB<CW^6[;QZ3,PC+8,Z8_
<Fe/XR\?5TWCUU8_N_OLHfD+b/9O+E^=e[FNI@U?/]AU991N82AUS+:<#\-94?U;
fc9a(7Aa2Y@KaR3M)c4DgR<&Lbc-c#Qfge.aEa?S,LcU(eMc;a]_00X;@#F5.#6E
:Z\+e2IaMJ7)2?(1-NSSJ/7\@AaZP_1#=_=fZ#L04NPM)53.S+M(HZ:-(7Je#bCA
5LZ<U<C#Z4c#T/)33LM_]ZPDFFX]A3K4YHfOO3gU,_E3\QD8EJM(c(BM_+fLf>U7
/Z]9a->BT6W^Y<A6(9QV5FA5(g#I3&P6F<[&+fSO>>^.O+]KRN,#GgN:4HdT39Dc
VZ5JKRF:/dd/483E.H21SCPR_1ARdO9b.]E=0P60+<^K8WANEEGfPJ)##K;&:KM6
6,9Y:SD0aVSK>BFH\Te+T>\@/>c+PN@Y03@Y7]XfTJg0&c+dM_b?#?QX&75>72IY
D51Y]ZdWN3?[L.ZQ(3-,[Pb)EC;/5B0]g2dDSZ=]YPI44;+R]NcH90VVe?<-THe;
6-N\E#36/2CB#BLP6X/DUL,T5]?a\ON8R_WY.eNIAWMbAW&-8.?7E6::CcMLE+7Y
@PV-EEM>\780dd(c/\SF@BUA10Q5QAZ>A4:O&X1@-;CR\IV,R&NW=[B&))[3e]fd
URI:0\c]CP2DW<C^=IeQVfT742Yc--W[VgVCSHfMZ-FdLMC]2aA]\&#Hc8M-GEeE
9f)2_J[79;0[:a[R@38X(bfRc,(=7g68P1N2bO:44I>,JXGDR1.HeV1gD^@6&[EQ
ZJAMeU6-\UJT_f^XWCTM&0V1QV3Q.(Dc24fQ/;:V:LA\]?7_:)Q63f:I,7;+EGJg
22#H3?0&F+[<Bb.UHM<\CDbL(>EK3:-1fW+,WIG&A_9MHFNKQ5ed8L>a)X]e#D4F
OddB=HcbK-.^J/P=.<&P23Y/38<G,eW).90_C_+cc>:gKdc]G)2J>M])UNY<c7IC
[RD<g&2[4BCFe/H#W1eA]1;5+)Kg.[ID9SV8XSWCRJe?S@A&#,aXQXG-eKb#)W6)
1-^X)WRXK[TDV95KZ:JP42O=7C@(BW+MVL@<14,21c.3=WI/9X)cUH34C)c80ZcN
HJR7X8X\8d_8)NXBVT_BS5^I_RbVE0TH1D=?e.4ZgG<3X3+O1MX8M04T.GV-0XQ:
B]W/98E^;8EE(EUU8IBJT<.M1Eg5SaH[..bBHQZcfA[MNW\)GBF5\;WFW8?\MG@:
GYI?->@9M&c9QN=/\&ACYcZ<Ebc(XDPD73JD/daYV>(8TC)-<I15bJXeg381a_?g
B2^?R4NIN3@M.I<6X0M)SbId1FgW4H/T,dAE4P2g:0].)dM([#2STVTN=P883?[8
1d>Xa-=PTTR?J8<a#78;_52U17gQ+F6aJRR-B1C)T12M\.M4JffT6fB7Z,a\SIbd
\F3#U^bUb>R-\#c29P&8Lg<QaXec><D0/G78A46;Qa?e.bQXIWT=34;R4.W/NL=G
bgC7#P:]_Ed@&.d(bYK9ZMaaN0#DI=22,.8@g/BI=eUFFOb_&gcAMT<WU/LWgLT5
+B7M0PESd4==G8KP3MBEPM]GZO2YQaUe>P-gQE&WV\ID_8X#fOP1[QcFA]DKI1^^
.R,.EJ[#@GID,d^N[6A+VRd53#A#2bcA7-M;LBcG^U/1&P?:8e8g.?4H9XdSSGHc
RQ7G=5;)[)_gfRf3.cLE.AQV/:VZg@(;-KY=J;,d?PC<bA60Gfd>TPATd4:[9-#@
M)gdf[H?:M@OT5:=M>Q(QU,4>^CG)7Y<5aEgF:W?(>HD#6&S[EJdWgC)@<&UE(23
[:FYPV#b<?35YKN9^[3=VV0K\]]Q\E8],[(]./>U+ge/W;>6]OZHJ>@\T6(66?cb
2[X;TV4cX<M?aPLZH,YP9A:->)7W=X-(RSd.d[N5KdJU0>b_.M@&A]3[P:M]f<MM
6e7AT>ILO?2S,Q]:^1D#HUeNMFg)=\;/Yd92RU>@ePECeE3GVYeYJ-<UcEM52EB/
LFW7VDT?S9d\;A?]7KSbQ?OI.M;VUN&@WJIT4R=a_MXJ.4\.E&B[\5#^>Lc]#<4M
F&J(1b+YX-McE[,dR=LbA)P0,NXSAC7W[O6:bK.2/]gRVTPY4E4#I1A\<V)c7#V,
cE:4\JA8#c:8_f:09g<29MNfC;R9AKPg+A+;JU.?5W+Mg8a.91TII531@=DFFUdf
.eWbS2/RcBU-0OO3E1K:,gZD84QC_,<\70&WXS=E:G&HC4F2FUQ&,85?BX9Y)aYI
Y<.WKA;PILDS+H;V>,2>4a+_Ma/BE9@BKg/)K1D1.R@6NI7[_>1a_MSa;J6^,A_f
JED_P+RUGE-LHXd,[ZAQ+TMEGZ.Ha2>>E[cST4IWS=PF:/R^V_HE/DFfM&Z-DaR6
V@bJSWg,V#YUKPE=GEKT/gQE3G#-/bJ_@]#V-R_[?@G8T-5,]FVOeBd1b.DYOe=K
MT/<K]D:NfTJS862=Y2H-OQD(F^PZ_.KG)UJ<KRE/6_62-8=FeA4,DK>SAF0UZ&I
PK2gc,Dc-O,aa8YWfUP=IY]:M6;HLG_HN7bbD)(b.B^E[LB>??MIIgBEg)[1c:Z7
a[gK4Me?FR_26,1J))YI5bc]))H020391X\U+UYZ19#W:=K7PHP.@>6@Y4Eg^^DA
caV(f1<K_5Q-T5;SSS)gffRI197AK/=OR9?X@N[7LK/CR,W\cN\&L1Rc6MGK2J0W
TCFUM1E#DUd7PD)=S5(P^5.Ma5/,W#d\g#&B\,gT\DE\Q<(>g>QH\+L^\;R/d/-F
>KHT&fe91-QF);7U739fNDHL?2]>^=:YIY0]AS0Ea^P;TP1Q@/D18U29]]?R6X]X
acc\X5.#[Je#8,(K2LNG?AIDHYc@M+f7GeA5ZDbbVTE.eNTMde_7gAO6);^(:II>
(=?WL[DG5LI3F-MCTQZ3LK4\K7=I8NV\eK6#GS,4.-A&9+2MP=0/5.AO?+@e_JUY
PS]R.4c3ab,[SH2/64=G.OL.c;\S.1gg#>HZ@?LL,a?JQV.P\=L<>8MegR76RG\Y
;Z8C<(5LN#7D[?7YYS=)fd?J)8[KPWA;]CF#CQT7__b]BUR<)TG1T.L_M2X0NL<Q
d,8<fMBfc8D#398U3+M-MQ4[I4fKZ,\.4b26@N<1?W-?.C\^+TG&=U8F?I=,-T_b
/>ee,>/I2X1_6^1J&D58dW8-1f;fD8E#gYb(#)3&(=)5IZ3ZI2R\ggO2OF54N4Af
A>bB-Z@)<S/+3N5B+BF&VH,TgRYZL?<.>@OF38YPMGM<fG^X/TOI):HY)?RcD&O/
K&ZR=b,BVb4,0V2YfZ]_&^CCbL,S.XJ[@NC4;d#a41Z2K/XA9S^8e#15d>M5Q3ge
G61E[T7<)c@(BOU1b&2a<&&4eZCZL>O6bA&VL8[O&(9W7gN?#?_/&[GVB=/50MBU
,gNZ7Sf#,XYR6&Pc0c8<_^fSWd9P#a=/J4#S66:JH?9,S+<@2AKC6CLSG2KM+1&1
[PTUO@d4PBY-D7=2d]R8eH01c6fK\1<JFTcA?;G)a2+d+-@LGINAA>PIK-UJ2dDB
U;H7#G.dI?J?YRFGY)Y,ZK4dd(V.DMe4X4T;;2^W-W3fS>1<6O,_ae]RGW8\(E3_
?KeV3>^_68eUJ2KS,Z-e[.P?F00fL]JKJf38.Ff;_be9FOc2?.fY4;O.J@NM[XXH
CE8V[9S4U],;S=X2::IC=DV+@^U,/e(T.5MQDHC5eef^8ccMM8]g.MBB1Qe.+Wb4
.>#&Q,H69_XVC92UU;I)X+JO>cU^^ZJJB2#Z55HPa]b-.6:_9/>D8:25>HVH&Y6-
dg:bYNM_?.H^Eg-ea-)P&U;NeVOB-:F5gH4UWb/:MH[1MAU97_\I83J1ULMcc_WL
)e/BI8WdDgZW35#]=IUZ2RO<_T_f<Q?TN);.>gS7dMI,S=V[X/.UF&FKX94F.Sf6
QX[&I5VT?98HQ(g._b[3Bc2gME,Y63#Ra2d7YR>NT:/2LYX3H@:;EffOdGHX[[R,
SMIgD4,/-N;BL(-HNND(Qb(JGeAWS+N>K7W^OUIN1/+X[D5bS<UARH^OKJH[>&8;
(^1,WWX?Vc[.bW32\)AX:CYfV?[e@bdMKA4??>KM]CRL=V+7SeMFfZY;GY?BS-EC
=(M@/DXfNIBW+-TM/GHRR<]-#^JDf/=+:2V5\6X;(67]f(APJTDXe+T1<SeYCVWB
?KF;IFEbEH#O:OMNGfB_FY?dO@H.R)K8Z1P(.F4C<JB0L=AV,D(RU1@4D@.XdWHP
URJI/Q#\R0X]&L;a[=b,Y68GA3edJ03:B_QBJ&?0ZMHa[a=ZEICeE]9\0O^b[3,0
X5LY#9;OZ:<-TUcPH.bLI0B)041NTYWNIO-g>b5I2XIF?JJ?<AQ8D^SMA+&0(fK=
TLD+?H]1-D#5G9\6>(.g@+A^CYg^+6H_+[7+:S15W+L82D/NRM77JNR[&9JCRF,P
^Udd3gXAPYZ,=L6S4.H5]^)D4L^B@F]ERF[R:SR3<[->&@_/+NZb)7<6aZE4OFLC
3DgA_7I\HfG4cRM9]2e?1J@4=KId4N9NFP6<aV8Z:YR:QMKA=.[dG&WM.OdN=V>K
U5\Y2eJ[I;+6d>GFH<)dT\5L=SbU+_P6>(/=g6+a44IS7_@1:1PT[7DVa8Vb,a,0
Ba(B;8_4/KC4.W4JNVDb/7EC-e8BAB/KRH&>6@N2EFCfY?a0c+I5UB@DVU()?\/A
bNB+OA=6QIdF9OgNT2:P#TJX[H+H<EJ6eYcW<@:9+,>S2QOaA5\4(-#RAE/ZT2EP
Qc9W_89_TCP]c#CKFAY1Z#\S?/gW:1@eL:.&711@9\e1-MUDLN7:eA;:_UP&acV>
HWPf^Y^@(,BcfPK)a@#PKPW0fM4LK9M>^UTPbW>YC=5=T](5a6HDW@aA>XdQ#cE-
DKgV6B25ZVRQUT,6/?GbbaONDV]dFU+,U<;BaIO2L<43[50;ceK.TF&GUf:BJZZH
YS>f67(<bg8<@/^G0_QbgKc/3ORdR+7P8>HU?ge-4V;c:P+Y,UcOUSb<1O,=2f,5
.ag>V8JQaG>O;)LI&#:OX(.Cb9DC=)c[<?5VaCO\Hbb+=@ae.456c<]9X:=]8-D?
<#Sd=]#P0GTSN]5,\:3ObZ5_O2Id8VAY0a0?P90M?4KJPf.TZMbOYI@(7I\W,UZA
GM54AEDVKG\aC)WJ71;e.gIRAaeYH8]86>ceDKGaK=0CV#WcN&P71d0<-6eEJM91
+UfR&R1WKSQ.?Kf>3Qc@HQTUS=cb?\?HY:g@8.d]d]CZH/WX&&e(e[I1/dLTSFXJ
4bH&fS)>4>SRFH>J,bT5D42c8DK&XZ,?[X#3;966B(=(CZ@@EC7VUbB3M\bBSf@E
V0XT/,0>:[F3f9g3AO:_EG:/+4-AVIP):)2c1]a<@Gea;2<?+g,B<GRML[>eYAAR
fbGA<OVEO8,BV,X<4P&#EG85>IOSJ/OJ<;XP1Na).dd46eCK[FH)e8P\2,^^@.Ff
CT\FBTU-&Ug]07a)&/\F=A,7#Y>e.>?A4OB)Nec@Z92[+)B[B@)c4W^C?ZcRgFQ5
M4L<]6O<;7?8XA.F80-9\)fSV;/]5F1<645IY1J(+K[Q3UP_RIJ-;@&/2?-Me#Tc
4-0WJ)&8K95&[I+[N/:a87_P?6U;Ad\9CNd<ESFXM,f[6^Wgf@Mc,&@fWT^M9BPK
IdV;4?)O-/@4>,G)/d+/@<]Tc=<<7gB^-B9?JE#9XeQ)2;U1O=QX@Qg:J=,ScPAb
&/=7U\e.9MF]TN>2<H#4E[]S_B30AZ^E<-Db>a:1>aT:2NcW=6SXL/,PS,GWP)KT
=HZJbJM3Qf]NMbV67EeF><2B[C3Y[B/IY5b2-N);Cb//QP&D?BIe5K>RVAff.e@3
dR.<?dG;NJWgHDA:,BG5A>GI.8bXW<6S[+d5d?37eK+Z+.),c?G,7>R8C_4Q3a2N
,;C?eAGc&J;9KLSDG[EDZ[A,8=&DICbLBJU6Vg(R9Y=\4eD)Zd8LP:<S8\?Qf3;R
)cAK^MJg1C<D\2^=/IXU0)9L/(1S[gHfZDCeSLR#Ia_Jda^@d>0-])PU(2g5+-08
:J+bSQHO@XFV,BN.OX#]B^2QA8[XT#/e5.0SW.5>ScIKZ8&a3WJ:dbQ/;MdJX/0,
KXOAT7.g27+PKIQcc#8g\N=12)8QU;+KW<T4.2fUd3M.UO?0KM2a_V;4aBZP;05U
eQ]<XP6NL#)]:_RW>,BUMfDX5=RF/S6b3K.fJDML24QUG50LfID&:X(>g+#;<ODc
\?4#dV6G-7[0WD):IQ<,.3U>Ygf+aM[>3GDY76B-1E0IfVI;/1)48XaZB:aTPeZX
)0-:IbAH#)FUg2Sa1\;]=a,7_A),:39VBB55,()5.K-)JG?P5=&ENBfXD7\A1?/8
@S2[+U5H&AZgIdf-_\PO;/KggDX5aJ5K&,\<4_Y=Md2OR,47E5U+ZU,J-J?e0QCZ
VVZ>fU+-/K:,CW>#<T5Y\XEFC9=LY:ZJE(9)2_/Y^;;db7)6bfXLRA[ARDCK_4]A
<5d(.M67^Z@65+U.B5,WW/e?=U,1QUW[c+?F7XEO>ZS2c2b:cTB[JO)#g9:SWdY\
303L4F^1#C(.;/[]YJ8(G=Y)GL[Y_:Ob//3_MFQPb>W/EG4<5<?+,-]/0&/@ES:V
b@G#F5_FS(fZ+2,+(K7CADYKfTWA4dWD:30a5+8+>SD9fbDEJH)[O.c;#:bcD,\<
=?UQY1T0D7_cGDbO]b:TN4PBb(?b8)I5GJ.eWXHVeGT6Y;M,]:=N_5ba@+P5b-=9
UPJ2dBO0PU,Tc&afRZ^,7DS2EL54S_3[B6#NW_7H^KOAL?JX.7#>M^JbOdYTRRc9
<M3NgR35B/[B<]?.bN;Nf4+9J[PW4^2\J0.2LS<,Z]8O#cS7,3Q+(2ZSR_Z_)dO/
CTgf/L<M.K9\R]4gZ(KXB3C^fEEgA_,0N\125(:6K<dG2&>fG#[0QR\))^=FPN_^
030MS^^(@HL;?YbNLO[)Y7dY^D]E#A/f?_J6TZVKR\LN?0A:T(?.340(T1A>)7bV
CXTXXe3M#G]f@Q5>9,5g,YAY33RP+G?ddb,@Z9R_SX-RJYcVZ(5_08CDSL7?:Y=)
#VIW2?D<GWKAgN\K:ZR0e&IM;F+3\9ZQ[7YSBZQ5K]E:26DN3bS#GTRAV/]Z+GS-
;YJVBX[bUVED?CN.Rc]&^LNC[0gI@>eRY)N=N?SgBZNCJ1-RJ[?FJ18Q<F_<[3GQ
Q9+=ReP:ga;<b<gSb),A+F27H-W-&:^4V&?<B>U6SC0]\W3HU7EL?+[TJ:(;Ya0G
=.;eN::B_@^8^T/8f-^D&A^@gP1O,T(@A5VDHe;b:QgAegg6g?A-5<LT5QGA=V4Y
DUWI46F?,KZ8V47=4PE9N\0dbgZWO.67:@BIJ>agW=ZX9-d7V]+3;6+dJ[_EQ[Ue
0,TQ4ga.@7AKB/_1dWG1Xe\/H=VfSWd#.&C+AQ9&CJ9F:@^(IUR=gP?Z&;A\79JV
QG20H#JaCNf4dTfaS54,<@e.V/C5C6?,Y[Z<)XUIF0,1:LK[ONA;VdaX?U79^cYW
H1Y#@\JeX&Ece#RIc?A.SB:[X?WGE[[0Yag)^gO)O-&285^UX=D6K7bgQ:8Q=.V>
2_24[AA?70;VW-)&3;XO^+V\b^eC14U=/^[Kf#g-[5DP\8F7;@C[T3/1X\3>\LcA
P;T7a35\a.[C+/3]X\Lg9([[4JGF9df_cAf=0?WE6F0T1KB;9LDS8db\?W-K&4T3
b,F-V,(16gfAZXUN(R6(WIBV=<VG3fRW_\:I(<VCEXN5g3LQ<M?ZV[=0D.VHJXU)
])MDW3SR,bbBA_Ee^@E_MS?FK7W:&+77;CYX<Ie5P-RA4RMCA;6cI8/=U;M-FT>/
IZg2SR_7c.Va>PFWg:71R,JMU3;0X9_G:J-Y46+9BXNE(f;+d0D.@W>2R?O?8B4f
S,gNHN,UAZRB/&]V:JS(@M38)QA<90&,,ZAQ/NQ[-UJ]DN@-/M:>(B0L?,<,N+eG
8S<ILIF?IV@0FHO40W_O:=&67-0M>e4af#?cZ=S@(<A&6KC@c@C&##4d=;9B<S(X
a&Bf&\PPQf:\a+B-1?eL59];RGQ?0<7(2VN<AVKT+3#FcWZ@f[3SN<C?_OJAN[N2
@X]\gFEN\caM]M<L539K9BEAG1f8>MO4@NHKFXN/e#_V>D/3?]RJ-@:#FRfQNF[Z
@BFf<N7HP^.H8LST@?9U\5VMT@+DfUU[;CJ)faK,bHZZ=#S,-_JLR?==)K2f6Fc&
J=BD#aR9:2@4&LI2ACg[/D,Z?8D1E<e<H8R#TU[[C@bJTAEO(NGK<;F=:Oge^FI&
_eFS9KK3_\>]Y+.&.Z2;KS^EN^SfSb34fD4NMc\YKb-H2WQYLFPWH+U_D-CWJ//E
PA55-@&C4/#SPPfBcLXXKEYJ=]#C(#/KV8,gfcBAPg;UTcD0>@A;Bg\A33&4.EV;
a4gWVK9)/Q[PaFbL;)\_]6OHM;b=VWK2[XUbX;X_[7e?V1UC(9@OICXWNdfgU2aU
BVc+O_+=e+QY@)>QaV)EaZb_+d@B,^^Nb46?FZ^X,(A#Nf,[2Tea=NJ:=2-HHe\e
/]]E--=(V=]<-D4MdL5b;JL_U1RVHIUS@YJ45_F8(TL724Z.e(H>2.2bab=S5aOK
Q.=aA)8fCN=Gg,UCG3H&:/KM+#;ce_HJK&7GF8JLgO4OVM]EECMfZWcY?46F?fC-
RZ<@(8a<2aRG_<FZ/=]YUR(Y>I40H3KFM4I:\,f1_;#/DCILZ6^eM[.X^/],J@R&
08Pd,)Hfa^)EO^>g8e]Y9_<[&5KIC3[^_>J8M3)cTReegFA])>8e;JENH)g=LS,V
_3APC:D7&:<@<P&2QIK3KX@?GVAO6,E8G)&7U;1)BUYMbMEGJfHJ/CaPeUQ18;N[
beEd_T+7;d)E2G:.DJ2>(g8-)I&9JCeFD95)J6T+7^W,A>I&adN;P7?7XL2#gP(W
\+5[Z-Q4L/e1XM?g6J>-E,fdJ)0O&PW\^b69,?G?<U\UHBOJD&-VHK5JK6TdW/D1
^3TOJIMMN=V,H:3\TPZ17+RQ7;>BS+N_f5d.9gB65&=D/;8XF[Kb1G3,URL2R_e;
e<TC@Tf1Ad8;)&1,LMDT7[Fa=6L#86F_X\-A_K7L)V=feBV^b?9LE,.gVXR]09HE
S26XCI_0Mb^7##/XWP5;5M9:aY_HO.E/aS=(3T82aOb0X/LVLRB>G^WJdgCc0?UJ
SdHJA^P>3P_I.HYO=5/2>DX+(M4UX#S,0gE&/Gc27][^@,V4(Tf<g+KNcXL4UID3
YbC&D]1VHT61>/G[H3:e7LWIc,cO;(QVd7=2-.JLf#YcJWKF>g0>8ULM2UaQE#(f
9L-e0^@OJTZ[Q;\.AS4&gW-<Ea->KU[c?<2U@[S59L,Q(RN_YLTN2:OY55^Ga75\
^T+V7efcEcaF?9d3)E()\beS3[,(+^a521/ZeS(@,MMc/Y?e\7ANeVcFe7?XH/.g
OD9(,#_:)E4H0N3&F7RQfY+I(0\Y=SZ^@NMQ^_XXA>g2<gYKF=--E=g0Wf]B:7ZZ
W,a0a3gddfBe_TZg&^#XeCfHbZX7ZX#Z4Lb:Q_#;WUeW=.I=T7gBZ/KWH9cHQ(+D
[Gg8J^2BR2@))X2&XC8@+S8>eWZL(4&E4X&Lgf@\C=8P_<<]YD22I=ZFIOVBHD/K
4(OIZD_eEaG0.._70),Y36#E):a8A/&ITG>#WJ5J7T)Kb/+eYB7.bC,B^>g:e_&\
<#[-[YQ;d2@0XB^dUY]IJ[/@15J)1\Ed@7&FZ)Qf[(>0\YGG)9d/JT6+3L&3+=R8
9O>B?D6AaBf5Y#?+M51NJD(Pb^a3@>]?(E;d?992;1_E;DQ^=8R:@E.cV-6:bBD.
IL.&@RA+;ESg+3-Z:d7H?^7(d-eNU=NYUXY1KLF8A8)SX>#0g6LK^\=\Xf05H\Z3
BEfZ\bLg-^6T;=P@./52167BO^JLMbfNN&Kc0RTc+4GGKCZAA>,)V(8CYg&f7\Vf
^[P[H@:5@3(#g59U9321gL;MX=N7F(#Y\>+T-,f)HM0@e6T9QIe#CC=T(&25U2-W
CG:@7AcO<K>O&58L7LE[F-4#)cSP[g5+QCRB?L/5SPQZO@4F_T929=C+F7-09cM&
?LS\FG&IM];R-M+-^22.E2U?_:#ZfL:Q2G.5C<ReVECX+IUEYU)-SOY]6VfWebUL
a1[7c)9DbMc82SQe24V+HYWAJWB[?=1[JdKGY7^4S],(0ZN[Pc&,UJfBH7E+;^3M
_)X[_NBM0ae>?W&gVa:DQ<AO#6U<a-#3\^MO^b<)ff1#56c6>6(e5A3@^BDZ;1:D
6B4,FK=[6<cM/aMg>B2F(X@Pba6\-(P7fHRAU](X,J1&D3,LMf;#65-9f8N(QBEd
E7T0@15AO6Z)]Z=GIdKGUH/4+Xb976YG56O3)gH88=HULD>GZA^Z^]KI6D;]QS9=
>;e5M1#X7;1YL(8M+K7[AOMZ=)MJSB0F_cYV01C_SJ8A7dL>^I7\B(L5LQ]TTg?H
8.dEH3&#PdL3^9SCMM-WHY6?F918517XG@0DS(87WPg((JS87g:O&[Gd]Ef5):LF
&>-3O3?6&VB\B,<QVDX/EJgR=>09M_FYX:b13F/Ra?(V76]5bWP_O8QXe+bIKT[=
ZAHgO:;^Z?8aZ>BQ.L:b/gc-ac-+6a.76[6DJ5,U9^PL9QB82VOS8b>,5QI3XOW\
VSg2J_X3,E>Y2_@EI_YT4I4[f&gTB/_P;b+JO,41aIcaJF@9e?];V/0C^;SDQRCY
6<A9_8A^c-5.N2E=>(-E:0&[0PR17^[,(B9WC87OCUVLa0PB,U=.=KaY?Lg[@)+J
54W>>Y[9If66NFgF[9UIbBIXB.JM.JXIdfI\@8cS7KJ?1W-RH?9YA4K66,R46>bD
aV0DS_7?FVK(Cb7C/476+V2Ie=c5ELIKNFCQSF:+>HX-P&HTLP=N)IWc6M6VFGJd
]BF#CQSA@DAFV13,1A3a\D2bNIY?EeB@]].eE#c8TL9(_Q9cQG8(/A^?Qb,9QSS;
O6dC3P#c(E-]8FG[<?<O_/..Sf-\7\.T[J\Q(@5Z8(X#W)28X9_&:7^FHWAI?M1c
/Q,Ye,P9c(c@-N8@^A44b4CfNe.;dBJF3+N2dOUcSW.K5GURg9MZIaV-17N^_Ta(
;64<e<WD/[Y5E?D(NH)E\68MA_UD/d1BBNY5>/D@<F5@0+:FI#Q:OWJA-aFS^NXI
SXRf&V9X:_L;65]))ERVeMcH5+7d,1Bc66e-.W@630#>>[G[WZGa^RL8BQMB_f:8
H+BfW?.F)Q]KEeN-CPgcObV=6&(8PUBPK[cJa)HVCaWMda8a/O;YReHO01,JQ_R&
6gYS2eWbc>LZ1eQ/>2agDFP_,6>ZA6SD\?4V0/CP0VBM;252VPT0<PBd0P:N#KL,
2BQI6Z?#fBZNUY:3JTFNFQG=XL:+(U@>CE6T&==Pg37+c;2A^gF(^QUF0\OKHD6=
e9fa)bMNHdZ/DGg_Rb3<//NPccK.[[6FX1T@;&7HJI-]C-b4QH3g78T@\,X>D2/D
&C5dF;eN:=Jf(GX])4ZW].TD5K8,H77J@SO=D:89#_6VaEM6GDK+0OcTcX8dO8BZ
U71DD6)bK;9cgSOF@6=MSPOLBR#9BMfD-eT1-IC#Y04a0,UeGD6239PPF2&UN^)C
35)X>&_UW_S]S(Zg^Vf6^f7Xdd,@(.fS^2GT(]&:<FU]-Q?G-3M]RIZW?::P=f@X
&bH@R]JdMCOP#><@)8C3,MH4S:d,-2BTX&#aZD1I^AP_]Yd+Ag+@D>eU4^I]=&_B
.GHA-T=Pcd7;dQ^M9EM7#b#RK?>a8X>Jb.,GN2VY1+d61f[X(RY6HIfQ6?##3^:c
SJgC)Z2U\I9S3cFUPJB4gJ)C>W.g39([d9[B=0L,-S_0J[EA+e[+]-MW4?D8-=HX
I3a7f(D?0Q3)=G?5gTC9.6eD;:>8eC+b3E=J_G2Y[(FN2=^f4]BY0.2F,U_CHfXA
M-;2NMQS4798O\G@PPM45bJ3,GdFIdOd9UD6[#B#[HD+)_28D(?+ZK53/X6K6/cL
(f&c5DTHbL&BWLOA4E1=K[HL><ZgS)>59K.,]6PNXT31JW:.3VI1SR;_YV=J<\6b
g,/;_Gd57&V+_8H;)E(1GY?L3+8=SbD6f),MN7gEgY8eXW,+[\.QUKO#:b[GA03]
GQEeaA4&_J18fVVC\)H=DAWeS+B#eJ#2XD4(RT]:;cWF4.12LTF4(HH]5e/;^U0;
D4)V+I6]05_7AJf_)/3K27_F;g[f#d_FbFYLL1\;IQ)_;G<MC)/1L26UUTWJ/\QP
aJJbX+b4IWWR=A<d[DKaLCSW5X53D1),ZS@N5\L:KefNO-H23>],9TB^\aL,&E7g
I:BC5/gD&(CB2I)33+)61F<9;E^A?EeR_CARW,Maf9<?5;V^RSJ(M<.5e3.E0(F+
^cgZH-c._bL62J+5G8]0\YBMV[GQ)O&DB/A/YG(FVLOB^&.&UF>\ASe^@dMJa#(=
6^)+cSA\9@_UMG/Q9dW2XDI5+OS[VRVdW7M\.G[Df994B&B@2@9@\T@FQ(.24-C^
46cc#2B4)@^bDQc]H<0AN#L0([aWBUC]B=@+ZM.&SZ4Zc6[,bFY)1cRXLLGUQ+<L
bM1Z&JRC[GPNORV+[3/e).O?E[LS5EOS>JT#SIQ[+eA_8;]P3#OG#G/cb#d^bU(I
Q55(QK0=Ca.4;KgEP.&^71K#9F>BP[eV:fa=,e8C#R/CQCcCeE:\#.MYZT5Z(#.g
#]@?<OH_7H/A9a[V3gCaBPT5C+DX.X@9],,ce/^UcO3Cc.PVP?c_BSeW(ce@Q(4Y
:\KTB4/TR]0:?/gJJU\B/bTH&GS@DX>A?AAU+\d09VI\L4;UIFA.Jb?SX8;;,NXS
W2Vc;A4956B(.4PLKD,YQ(FDUBgG2M32K8(gM<UPH@#A+U/A3,V0.][>;3QIb6Id
II15Q==^Q3X.\/:AS<g@ce).H:;1,WL)a>Ve3H,Q]P1OC4IRg+I8-5a,Yc7@=>AD
9XW1<8;MH]UF6LAYUT6?c6PM\7]dTe+e&JQK57)/2>U,_C;HP-2<\BUFb-4<_M8V
aA3U@8;HF9Q@Z&^-dHR?eG&H3SNVf^X_LfC-eM1R2Q]0-eA&UC[-M/\NTa6+]D@W
C:SC;YC;71M<K^B#faZR?#[VRE\N]G-Y9ZN@2OV-U@SKBg>=HEN#?.^(P^F?/P,c
GTY?/8_cU=.Q[8;gGP.RLdQHfU6&GZ&4+KC[:P&U^K>:eOVRbHN6L[,T7KRZ)#4P
[)+WC57>/J]_J7?#J_W?_Y0+e&Vc&D,OW(_V=M81@99G0NgGL#Pb\LXV:UN06B/.
@K?HIRaUNTER_g/3b7gW9d;H.7C(E/PUZ28/OgP-DSQ93D&D7VL4W(A1B:c>R7Qe
7]S1U_@Gb/F#_/(>eJUU+DREF?O&\T@fVF6GZ90(cF,<cC8EN^\R4SXU:#YgU.MJ
+(c7KM=AJD<g?XQWQd^&ZaQN/eac1_@ISW.O[\H[]faYO_SN>L5)#Y>SVL@>,H_0
;,VUaK>F1SeFXfN,,84[IE?=ZA2,6K47@.K[XL)U^cR2KM\E;.LXPX\&9?b46J5/
I.I^_[OZB\R2WH7@7^9OGE^X+3@?L:/?(e7:U]@[G#cY)fF+0:09b.WYFO8CP.81
?7,<8IIP4S]TA)L5#b1@W@0JXXAZTAKSNU)+Q2W5N#d@NL9]N??@A^&_);O3fXdS
Ua@XYI>=/CZgd.7U=+WbPd4V+7+g<?KGC^(c-VbJbc+HY^N.RX.O;\@R6M-f<-aW
@D@3g^T>P5\<.-PTHdbf0DT6_]C4R\?CYAaW,BZCe,cSL5b&MDaRc;DHD_9V@2\M
LRWSL5/5+9S0\RTIGRP+:4]HEB<Qe&>8X=dMZ,3?Bc_6>4+f?U+\G5a3&B>8+Z=K
JA3a#F9A(7NgLTXB+Aa(XD>#:Z4.-+4\eXM1BOc03,S9Q.R;@c;E-0J[IMRKZ;gQ
YS#g6&+-><A/-HS(-V1PH,Ic2\26H4/H5W3b,RM+V\d3BS#D=K[]dEB#BTQ^549>
d_05ga:gFA;aVG_b\J&e5BF^2O^8CJfLCVH^dD<@56]WFVW\(5bTP6Dc+&\V7Db\
bN?W.JS@NZAR:198Zb.<^]P:0,b-H<552Yb2MCa@IUeSSET,1cEGcU>@??I)6ef:
Z8LA\(U&)90<.S&fW9^\35>Q8Y9?]ALeC>Q4\TO?f,Y@:<U-dJ_6H_J@<ADR#bUg
@(S(@36R]6^L6:^8(US/BHAXOY\#,)1-;O0dDE?49<4&cS/,RLOWXKZH>>;?YeUO
7,YB2<f2(CP:P9JPQDEJX2>UP<^FeQ3^V=[F[D/-D(\);1ANALENbg^-3OacFV:B
a<3[aR^\:EFGF[b@c#=?\G\DFU:LD:(ULM>S>Rc?23a#M)AF<;D+5N>cUH&ODSPb
89F&K=^;?0fVe_A#XMP\>1F95Z[,4B6AXD-T;7>,G>1[QUd93LB2J\faM20(QcMD
ENB(?fK(fD<AY52U31d[B6KNU]NTF[/FEM+I7VF4K/5J)d?dLC)C_JB;ZNcEWLK9
g\=UNGNU91#GEY;C>d1@1Ja+bIMPL3W.1:1)#7H)QG[N0N/HP?CcC.PQZHQU><Y:
GQ5BOR@B3Y8\-54[V5]3:RGWW^-2b^Bg<C?V=].3f5;QI]CI_=;02D=gOJC\/T,L
SS7)KAC[;>>5YJ6-Q/0N<,Ddc#-&4?>>D(/+;JUF^;(HVZ-]&bcE,+MM[+PFd&^1
ffL6]dWH[<;:UEVN(b8(_VWXe)OD/?NC32deB@77c57C6]<0ab>7a#_#HR40X=#<
4=C3>]?06g>f-7640PH]I+6_1ID4V/HD4fEKLWTZe]SL7c0R.K[-UCT\):L3T8W&
01A3^_)a9G1c=53,41H=c_9IS3^&(7\QUV_a(-XQV=1YC=Z.\.W>3Z>QT=QA_S\<
eU8W<:(;]bg^F<6Rg;MBZ8eYdTYT1.UcbV(XQ04R_gK4B5JV9^JfI&\&&.FVI-\_
/FS;HJ=]]0WY<HCTYFGLMbT824+=P09JM=M0V[>,&I?Y/W4DXK/]\g2Q?@A4:&K+
7B6,Oe,0[Z]<;/LD:.]HSW_5Rc1VU[N>UV>:34Ad_S:;b].ebaL#;caPa]OSa:O\
WL-)K#^U#<gUd@)_CW)@A4[T./d\KJJaL9<V6_Kd1E=76CO()LD]RXJSDgT/Dc0+
bF;f6>2_1:V#,OI^UHHdP=gM7BSZ=\&_MWYIQK=HH2=:C7;\d[;H/RU\_6Y.BUcT
.fNMb?E+bffN&UOCPMPFRg1(d<SW43e5W4dP)]KK.12KM7gFE1bfXT9>;[2Z>^KZ
KC3FF/G6>OSG-F@,5_SJaH[II>C+Q9eW^7&<6<T,_^+4VKB_PeLePI0G8d)5&UP0
\6W2_Bf_M&OC.b_8g+dfZ9:EDZb,C651801?O9XVeOgS6J.0E:@WD6^S\B233.\P
/#:I-2P\3[]YLg+EdWHTH=_9I<EcG2Y7=FD(O;<<6T0^WG2SF71F==:.FD)97L18
dbdM:,cg_Z+,X^UXW]HbFX3#H6@+CbIW#_T4HJ+Q[.?-_Pg_JV[\=3KXc6,[R9K)
F.\TT6[^(YL=MI.SMeP<UBaYNHb1S8X_-W3<RKQW)9#&CdF/]HCNc7EFTC@>T]N6
]F9.V6]OaQEN<\5A-D.O44Vb7Rf8_U2XceKAP]K?bJ01Jg30VYH6Wg0L;B[]^ODD
Q,/H(;?dBb_ad)JT4A:d\a-\dXW>:cMa,><[N#dOgJ.XO#9:U<(^_.]QBA7-aY1/
_MO(+DNB9&)K(R1V-^X[DGFc:0).6H@c?Z@Q)>+LUVb=;Sd>_;Lg(>H_S_5#RB^R
)WVUd3YU<<F]F_=2B<,E]0\)V?W394J0+fPY5252X=@-X9F_6<T_M)UY7622#b82
CIMLBCC-)#\[:-5?cFW>RA]FXPg;NcYZ8G_2G&:OGJ#]bd@6<WgBcYJRR0;NXd(D
Z<DIL&:c7c=A[?CTI3d/2]D9Q0+fLOP_Q@^+]H+&;Q>+?[;7FK:-cg0)7=V80#2A
\dPO:;WXPA)48CQbPZP4<DeFU+dC_fLJ-AG+<OF>(:U1b,H3):SQK6(YCG;:I^Ce
2=+D8>Jb0V8faM<G&AB43^3JV<11R^g:3_cg+cE<_H(>)2XA:\FA]H.2cJ_R-48@
Mebf3JRO5T7F3Q094.W?_g8XM.3b00?NbO>T9&F_0K1&Y)8H5Q:C:Q[AQ;&,cO(f
4F=fHMW]V(?O@:[7N99ZJf<U[Oa5KJ]DB1/e).S\8gdg&6>Gd;+cK#W#X)SCA0eT
WQ/][D.X#3600WQ@\L#T-Z&UdC&gV/FMaBGa>@1fHUICBHEZCR\9]ga]8_&VT3-J
/#ER6DFNK#2MFPURBWXO?#LNY9=aeU<JNMX\c2gGRZ(O7Ka<ZfC[>XY1(,B/:IMJ
\)9Jd3/U=MS]RITG3S?L;7873NLJ+V)a]f_f[XVeFO7(g3BAbM1WJR)GUUeBS<Z?
M=O8[UOX.]_VGb,fY&JWdMQY\)(=->UVA();1\\R=@K+e3+Bb\cZW0G(_&8a0U)&
./a216:B;cBMG7/0MZTV(W6G;2NdJ(^f4TWF-RK:4:S9WF+YLA&A0SVK,YLg;74]
WAY/HWJL?GV,80WNV0JLJ3PFAP@X<3MUM^O6@-P:D\X0Zabc(H4RXbJ69e1U<68?
NG[+6JV]8YJ9G[M?>U\Nd\F]a/\16+WED?&>VNBO=G.5>9XZb0OOR/8?c@G[]f,e
O-]c/>/-PC9^9Lg_@<\GX-Y_cT3OXM\C9?_0bcD[eI?YHbC6(]U1C5ENJ;\RgYO=
M>,9)Z:\ae@_86E(8OWf#0Te>cKg&B+..^Y-H7HT)5Y/1X_F:;Ae5&NHOHd5egL&
S+O37aK.Y)0ILLY\c/=54K^Pc8fP.3d1BTVQL,K4X^[#RWOTHV3fbZ;(GNBCYB^8
3PT3R?>B4JNdX^f-AT1[ac#CMCNC#(VQ+cI@c]YV-7RKOY^K5fYQ>0EC=#caB<Kd
&ME(?,b1d:?HTdB]0EZF/dKOKfXBW,B0=B0\_4@(+eREaT[P.g)QNAQ)ae_e)]MM
V5K[<MeT;\5)-ag()MS8B#U/ON@^5A>d9)g&B[N0d]U9a>AMg+1O3DZ0#6f;5Ae3
(S&C)CYaD^abIEQF59A^.@cZ0=CP4#_?=Q83(^_2V<L@V48E5VFJ9B&)FK0>eR.Y
MCR[4?V=4<K[QafAHacdUB/U^Vf1g[5eZ.c-1dQ\KH#E>.g)10OM5K.31+(R/F&=
/0L(<J^_&T>)FRDU/M)d@f/(g]<F_;AEV@QSc?gRJG;LfI<H>YQQ4IB7<)=:16_G
L#IXa&HY4D7ZfA)FX[+]9[YD/JLJX:YMTH+Xg8Gf]Yfg0+gJfcFW/5\C4PZ3</VB
;U;1Z?d[dA/]1KNH>CQ]PHY,6X+gS)):,,DRSE(YD=<AOBc?b&[CP8NS.FVab,F5
TT,MVM\3>GVeY9EF9&/?[ZZ]Rc>[RgMB13R(I>5;@C2A&VI7Rc2cF#ZaeN_\YA3(
LH@CY6Nb[PA,A2a51GCNP?]]WcR@S)g()PV@JA24^egM7-1_YWNWfd&G-g@N@I2@
@-:&W06II6;7N/],,CR(7dI?\Y-4dG=[4]0[1.@gVR7_f5f86;;/c<+/TR3d73CD
2;.ZR8ZB60EY00<0@F0)BN_HR)ODKRf3OY01a.SC/T8U^^dVW2DCKUW-+V&\QMAO
A<P2;?JGUbF7<AaBa:g@\#8U38L#>]^\(]R7KY+5L776E7:We(QNdG=fVbbdO4?\
J=#3b(6>Z^@YIZ,R4FUW7fS2?8XD^26[A^@d5O58A[cNHXGN>8[FP<c^4@>>bG&2
d4;RS0W7FV2@c,/bMP\?N+W6M[M2EU8[K.>?HBPDc,dR_LY#46L70AHYf^f8c+b8
McG[08OUgW6#MRL.;XM(X+[YV.D]\4-VB&J/12?EFdDVW3\1U0CXf9=DBN\[HA,1
\TdbB6C]&<_#?\YB_fUJ/Y:T,O4A:CRP21Z]4V9VcLWdReS7/7-8b]MCbP87:aO3
9[[7IL;;5)LT@K.H+LK7CSTJD^5-6U5fJEg0]5QM35=S(^MCgC9Eb;98.OW]3Z<P
[XH#gIU&)=#GLO<HcEEO:fb72VBHK?Y+4N2=TdKIR^cV\ODd6ZL5_f01ac8Xg+_]
,OeQ=9K,[FC7/>K3GDW\LHJBYGREWgOee9J&@:M?K:a_U_Y+QT2S;HCd?>V^TK)-
WK;Wb:;R?Q;4eGJ7a(8IN8P2-@A.^PK=D,TPeC,E+@G[_@0QbfG1:?P=g@3;H6))
^BOf88,-N40CC#AEP:a?CETDM(5C.F4S75Vc81IN0<dK]0U(c3SUP<FbJ#eTP:-4
^4>Z.T4I4J=+Ab[6fcW\PU[d6A=f4gA]NT7dPSfZ4(0b&J7GM\<KBJ?a57V]gU@Q
5LQ/B,79ISd.Q>V](=+;DQ)C,Ig<b0eaNKa,\3>gXb6V63R+C4N]2Q]acH]7<)W/
?Ug7+F-2H^TKG/K20T^59NL9a>M09Y^fYN&7D?P)X;^QEUOfHfV<5W[+YQAT=a8Y
,Z6Lb_39DTG(fGS6dDfLgHS\8LYJWg^DgY3YX0eSe?((L,RJE^DNb/Od_\Rd5WO7
&WN:HAd0TaI5f5C^I(5Jf5O1XdU=,<CLE[007Y43+_5Nb:VgY:9\IH(cD?Fbf3-B
G<BW<U<Y3\MaD;#b3f^77C8OL[HQ>>aG(LF]LAAL9_:GZJEP7Y^Y3NQS_3GS\0A+
6D7Va@H88PEQFbUa8&E[>:NNZ:;\X60>X=RM3Ve:E)dXf.GgJ#bH9-GLVF[G]e]Q
<I8MS#IbWLLPQDLY,TCQ^EM[OOWCS\4HN/E4(URG4MEZ:8\0)#&:<7V#]0S/99:U
5JeY[-Y1cDXKZdN4(Z6aP:3Mb\FF-ESTe8MWY[e8.N3b\]]V&_5VJH,&FgEF=[F4
F0c2+(Q<D?G?@#H#LZNL)U[Sg53]:<553TTb4;gg3:G,GJdGQS9SbW)E4Nf+V0_7
@C:E_K[d8:X?I^0NOI,N541/g^8aQP+FBK\T[LH8g0[6/>916R&aBD4cOTUA4>a@
+^4W]dV\Z<_?NSG,T]DdcPOdT(dKXb2Y#4O&#58K1\+Vg9cK<N=.<QL1geQde0-?
e&f-&JA>_<I:&#f#KNN^VR4TD:Z9)BRQFF@L>DaO8B67+1+)IWV,N#C-W=-e;K)(
aK>g:FR;KAF-_d6g];U8>16eHbFA?JEU>&G-YVg6HCD]>?AC0/0J5]AU4MLGB-F8
[d58/OG_6I:;O_<_-+#Y@\;A:G+<;,Oc7U-#&3V/0R>L;Y^ae:+>3PC:M&4]GV6)
>B&QBKK>PN?3HYPV<O7=DO+^8EP;E5E+:gg+dbOVA<<XKFB\.84W1gb=5E1_ZFNX
(fAUDHQWVGJ;KCQISMe==:0.OeLcXU+Od+)0/+1;?-..G_>&()SfDQF@R0BB\/Ve
]cKd)4NLC7]F>WZ+gHS)f#&.J5/@\H0T2ZdHQ.P@4SV<S\^TTWJ.3<a07SY5F,e=
,W@S[HeJ54TL\\aGK5GC>Xf:WFQOI5DC)eUK3)32@a\(bY>R24LcQBEPH^aCDL6>
CEPK3TSG1A]Y;TUG54d-bM:@>.XF?&;d,?6P2I3T>dPC,O]31UT4?S@AN__)2>Q.
\LU>,,b[<#.FdX^=<IF76J?gWKMX\:-TJMaS(QgTLP;HR5=_ffW/=@@)eC1+OB-G
?TQ0XX@_8<6I^HZ@D^_Q]/9HJ)L_=bKT4G:<ETK[Fd+6UB9?<]RVSXR0;F@[#;8/
Jg(fe)=8O^bJ/K6#9-T,KQJLT+9)LF]N:KXS6cNNMP@CG\:ARI0@_2L4<@OLSW-;
>M29E<P@,OcB;ae3^gI2RbS-WF&caPQb6Q0e--RAEN4KfN[S.S<URRO..L-UKWe.
S9GM1#ID-\9GcKf@He(:ZQUZ-fOEFMG=)fDA(J^I(:=&49L2X;FS69(QY]OKAZOD
gXNKaGW4?+Sf7DA\3S>4[XW@D)FZWI?-2D\I>6/K7eUV-8<BHULC)BNC6HOYN8XZ
/89742M671)K7NQK760B.P62DX7bLWZO7FN5S&.DYL4(0BTPVe)BIFdfAeNg>A)A
Age4WP_K7ICLaVQV-^fW1d3:FB+&aQc1E_:f<);#eaWRY]0DZ#4]0L_B4\fcN).,
2VXe50CS6Ze<]9VB,PF#0BV-Ud2;01@OO2A-A7^5O0Sa.R7\WgX7f055T.#93JOV
ILaZIT<]JA\V>dF@cO)?f@WS4[J7=Z4@X.AHfecU8E;K@]O<LSXL=A1Tf);4_4BI
^=]BX#.FK1Z:MIAAb0<UTWQf()@Y,ASg;HEA98_1T4EB,Q@VEIACd:bBCHd&J?)+
Y&OSSB.QCBM5Ka,C1g,<eTcRB0J4G=eOKUF9VegJ_0Ffd>=ZU<?@4;c:#1+c=82N
Y@.4OacbFIT)9dd[8RSF]U^#a,cO7H<Z;8()(>.Cbd8aHc^bF<&?U]:4I=9:MM:(
DEHX79KQ--BP194F-XJbBFG]@5MTDJSD=^MIV^=C?TeF[WF+^T;9HK[IU+8cPRB[
93QSX6_O1ZKT?HcUO[]BG4_5&>;85H90@5]B,>U-J&W=.;?WTU571_ZZ6Y:a)2V+
U7YJ2+#f^;[eE-/V8S<61;a,XR=>fVA3I6<V(20eFE&#\T:EB&W.:2GB=N9.>;T1
OEeU&Vd_SMdNg4SO-dCT>))S[Z0DW74RU8&_/)GUEFTT-#P=XT6F1Z]@gCY8;6HP
(Y1X_VW_6<KZ^D0^P\_M7OIaDQQ.1eDcHWP18d+10NIS)V/e?Hd8CBU-CV6\8dDI
-U)^G=WYF:2)E/PgTT<GM6HE7UEE)KMc@23M#A#=1/HL)1C5ZWd-\-C=<Wg;#LP^
8cD)\?X:1?DUPWC6Qd0eRT3J>7IB:A;W]-@+eZK.8JaY+2@)7dV^J?Y.>,,7ELd>
\:)CFML=OSbQ;)LJ]CbBAPSP5E6@#df@@6[_@8P[JFWA&A8R@ZD1XR9dJNLKRJHJ
G6R/&.[EA;@\e<Se_a40N<c3=ZT\1fg:R6dD3-P^Qf&3IOKP\)AXQR(XZJaOFG4(
<@M.aU-9Sg83]6aCE,FLMddLc@A&8^2aAT#VBYeU&7)b.A7bHH_MAIV42TQ3.(b@
RCU^9-RPa=E/Y>Te&X,bd372JW\G+?)Z+-?VKJ.#UM>JK/bGK_SW@b-0\7gQ<\GN
7;VU95_D<AP]]g,f[3/aY)aeSSe+G6V/10&(RDEW[=2Z,/SA/59RI),,4OVU,XZ=
F?=;KVESe>\?FEbR/K=eggN:_#gY-@Ke2F6aO64@(fE:25+/N+LTA1T1J:E<KZL0
T1#4S3We7dI;AKF@)FgTS\91L[UI<=55d<SVVegE5gbM945.[;[C5(D8H5-01,b[
?,;G6A<AAZF;0)@dg_MU6IHJLUE?Q9^VVYJ+\.V\7KgMV-\>,Y>VZ.75#]GX#]C(
D(1&KB,e&c2KC+Sg\a^X#()U.3F2#FZQBEBB172SAIWJ@CZOXc#]B>C^)[T>=Q4(
>[DWIgE8(R>EO5<Ye6UO&^/Vc_82O;Af=YZ2cX@,T7O>K^b-UcIZW-?9ZE7#B1?&
:TRQfXeFEQLF:#IcYK@1MF@/R]gbOOfU5.9OU,28e1@<-T<-VP0KEV5895WE=e^3
TK2:b)-]<N3fKD+S>J@]_/_ef03?Bf/DLBa[d\B\6.edSUD=W@1F;DUZF0=K+B.I
Z9)gG1TJK#WV0D1_9?g7A,S;8@SH:2bPS/M.gc#eg(626KD&C/QNe(_PNOVcB6/(
]A+eHZD=Ce22]gPBOK(-TNP.#^2;_b11FN[5&98XQ@?:QK3c^SHIYUgE_YQ0&WU=
V>W&XeBSTPM4d-W.3@bH?Gg.+)RUUYBI9,Y([DO^SgDDfFg8S(MRZ=&IIGCVcQP>
^G\UTIX)H-gSgOF-P),H<W8D,PKC<^NZ96;VA3=g<^A,Z(OQUNgLf?;N^;bY3P+d
H53&]_KGU;\(9Z[+a:CN]Y_e@6[@0W,NZ.J6,O;L;BJ4U^JQLeBAX+O\9P,O_5&O
&].,&92YB?W_?C6\1DW7RZA8?-R+]J@&_KGWF@_0[TSHN[<1f..KG6CNf12dUIIf
R?2\58HIV\ODRc#eT/__S\E(bAcR>.aE-Ia/TIOPSe<]1O_F7AB4R7F[0,3]e3gJ
\)W?8gT)-1X7ddG)7TKWMHS[=T6<L&HK0NbPaF5RNHfDZQ\I#5D>D-\DH+5AF7(f
bRJ>B/IHe_S@Da69,4(c0V^P]GN(G(&Z;E.ZV4DE8UgR<8_Q&)gHAa4O6(Fdc7^Z
0,/V4X\J<#IgT1\0Bb9?2#T;Z_R/0;L]:L<Bc:MfIZ^J]?4&/((T2KI47WTed[VU
LN2BP70_J:RHO^S_9YUH)KVeF?b7(Y#Wf&[=04AK\NE:4DTJ?Ne;U##7BU-W63]d
_dUCD]2AFT_cR:bD0gaVFaf(X_I]F.VND/44[?/:/#@<d\-,F1QWddCFY;:YRW^W
]JeX9Sc1IBQPg8bP_Y9Rc7Y813_I>V1FVF52EBS[:UX9R.ZLd0N[a&3__K4V>L)7
1/<][/c.GHVD?DdXU-f\)aH4>79Q)P6NM)6AgTDE480(5S(7CQ^b\Ude@)=#^5T<
-BCBPcG81gD(AKDZf,X-db,Hebg.7>NfVJLQN1/+UC2>M4#BO8,H:=&19(4NB9d^
N^GT7TQbV\=M\_F1[#a/VJ1<]e5/RBR[F/0b0OD-KaFKfdf2>e:\=3\+_=Y]FNR/
add(6bc4ASRSHQ5Q2PG8N8Rb;T\_<.=]2H6.#M\9FEB19N=E6@XIe?dY1&6G@E+S
B4@J+O7HJF674\&c:ZP(UYONgfSc\fL<.@00</g-](N]U?S-]&(bD)eWK]NNZ8-8
EGR2Z#.>d_UU,_VM]:&ENYOf.D.V[\#Jd&8RLK[\VfX;0<:aTLT]XYZZWA^d1HA\
=>&/P4;PU:NJ1)]7g\)\;WeZ=G@64^_]U,T#@16F;gIW^PX1A.@8,f&MFYXc9=7I
e7a9ec(KU^9:OK+K/B#0GSD8c(BY<GC.33);U[AX@1(H#@;aE:\3:;_f4C46>^KS
E))2L&cF.UM1G4,O2e9+.1T@GAY<N1)NN2J?MH@Pa36>c8;N4O3](>;<IG9ILHD0
=11_ZKAYa(<R81SZI\._5BY[<f<cU0d5bI-^V&R6U@45L?19.4^g^GcOg6^ED2Y.
(#@ML3#H@PWdNe7eN=7b]@Z99W9OPW(a2(-;Q)2X9[8FI4eRG6b@4c\;b=_^c+71
;gVTOHIY[ZdCH-1a3TY+;_5=&Ef:Z/1780H75X-cX(_e\1>CF0cG.O:dH]M)U9;0
?/a3Q)PBIbN7,U_Q7@C+3JWd+_IRDSaf-R#F=VK#3.;2L[J=b2K:A/]9)(533dZM
[JdFRU6cY9C&S^M\GT9M9<?L5Hb,&UVX__V-)fHLb>\,:4;S/^e5=6G0O&M=KDbV
YRK,CK)IWU-X>R1KeM6^5/MFf(L&4_D\L<Odg?2?0MY/TO>F]_J6H@g)8#2K8aJ<
f/UE(=36VM9^TNU.TD)e?[,<8A576aR>6]8W:;>:#.FRLWXcW(J(S(\L_9ZIc]6(
F09,V5Vd<gW8H9T_[A3]e#SP7b<R0X;T9_=e-,G(E3UKY#M].af3W9J/b>&#:#28
_V=V02c8R8/9fcg58A^cDG?b&-EX?&I1ffJ3#D-H=/Y3,ARgE_25Q,>\.#EAgQZ6
[Eg\C04T&U6<^Y^[d.8&=bM;3>:4E(N>)b3:>/Y(7XF;GcHM\?2_]SR06a;0?(=0
,]eOa9]O+Dc[N2@^Y]A1a)Qg^^1<3UATGa_g(gdO&e+5UDG9e[VgAVeM&/a1U-e(
P#gZ)MGVWa-B.:L4(WI-eH;9C\3#fFQdKFf)c0=B]+f-1-dETE5QUJBMM6U(6a@-
f)M5fcF?Q8)PQN+2[eF;CDf>\/<BNcMJK7Q3KJ&c7c_T^84Z)_Z+fU4AfQdCgK6e
Xf-Z5@2/HEHW;;=)HS4fG&[0_Q4g4<IE_Y0X.[AMP87@FZAQ,I,Ig1RGD8eOGeGd
KQ>Z;4,FRg:E:?B[WMCX\^0Ld=NSXZ=3TCg5V(d?@AK0)GDbKI]JF_(S3NW_g(>e
Ld,7W_(W9>d0L^SS1BX@PFK0>@4/]YDI;a902U^^@+/D#d;eWd\M8MZPP6-Lg_bb
Da??RQgS;990fND0AUPF6BWNWbI-8,)cbFf?500Z0c7NRE_a^ddcD+=_^;G2A.UU
>SV&AEOERJ\V\S\5=;=[8@<0E(Hc+e=8\Ze:D^)[K)KWUCMSBVPf(JH:I[5U67<E
b?#bI[1K5?eaKf?1O-/OWe1;g7F4RXeE5CV9MdcaPHbUI&LI[]SF6[aN6N(1(8GW
f&(/HDKQ)6X;/BeA1E#UX1FJ@OL\6]QP8U634X.9cFI>fU)PVVgLU2,GV<d33O5)
UU881/GX36HF_,6c(>J2]+[(T\,bf3U+(Lf\d5F57R[?ffXN>6cfR2K]V6Za\K4U
-V.E0HNbT@IcIM(Ed&<V-.\ALPD,J.YU,X.DJESAOdfX\_a#bcFA9eDa.W?G/DS4
g,X(5\AS8FIg1aOWJ?<]X54d/dD9?BQ,@W9_g1=45W@\?E9;>&_Z2RgW><c:7W8>
P+:b2R8c+1FL-<QJ5#(ZT7?MWSQ/I#V0W2/SXHA&QC6R:H[(RTOYXXM)#\7V8[N=
;F7+)NWCKgMC7@Dfe+E.6=8,]_-&CWT9YB]WS)Y\9[U@c./8@G#D9:6Y+B))\d13
8>JIR40VL]@?BJ#/cTQ5X9d^4dbbg:G^N/JCJIM;.f3>HfMZ;K4fSC_YMK-Y>c?[
Ab(O9-9DWE@eA7_/H4.f^U4M(6<#7CEb>Z??/^:XgC>34\&dM+U\VV;3ET7QL<=b
d(c4-[9U]S]SM&5)+#97ZEN)O&9=EK:0CE<BP./_^PQ=3V5WXeCY.a?GYP6bJc8:
[OC6/-9DM0L4&5)S8@A\eC[HB,gS)_>1c.Bb3D\YLf8=NL?0=AB+d+V,a3OM<7XX
WFX15,7&NG2Z6SL^2(+0R,X:_4DF/+)SY/N-\W:d(1L.AU;NDdNS._gd)<BDA0U-
=9e5g2XV>7UP.^(\(M-Rg7V;8F]_FK9CCU]MJ\S@7Q@GW-3AQ=?XE-GFLVG/>F<1
LC3-ReHL=2QT[V8;M.Q_b>GI1geOb5G^Qa=+8WeL<74M]76LB9cMCd5<-\Y-;(^C
8_9gXL:&Dg@_#XGRU_I4CZDbg/E^^@7?EAE)0/dd](2\TcR>+#MXJe#F(28+7D@d
Eg<gCZ[g2I6X)U/V);=gZ6?J81I8_Vg5S<J<MfFcZ\VD(IDBF-3XA7WMORQZ6-(G
g)L>Sc7CAPd15dA&F6RF4OL/d/MK;F\6FB>V)3U#3]3Ad38CbKNBO2C-46I,OJ?f
1da@bcPZ]#eMKSM=OMJa[]6aW\-M1+N:B>4#&23ZV,FY#]J2\,MCXMZ4&gd.46V)
c;[TKZJ@P6WQK2gX7?-@X0,B>;6SS)(JdL/5>.IFC26.JLGN6^d;)0Db4_d,=b53
>ECD_<H#4B:+V?1c?H[U-U>^f@G0O;8_Xe?\1V#X1P<?[>E(J_[=[CN5:3>[2gJ2
YN^.5+U9H?76FWW[4M#_Y0(I(WJ-]QJe#7#8d?OZ.#E4)S]-8d3OV&-S&e>2NJV(
d12&dIfRU\MA2E3@/Cc9FHcZID\PC1TL.V=>W/Lg>=2a4f8[;>,//U3_Rg.A:QXJ
#6J_0>53E)\HOLB;V\,T0HLMXXTW]@#a/1M]:E-H9Nc,a?SA_W]4]T4&R,YKW[+C
[=G?D.[IHfC=S+CdULcM#O?Z]#H72[fCY^;1&1g#;gMJZ_>_9bC(LcQ-D?3+e^)E
J1K_.EQ-X0@/c<RJ>]66>F,O0d&1T]W5^+62;WeTVM>eU(UX=,Q?],?#QV2=df0g
;LF2VeL1=,L<S/7^[/I+99V6H4#_:V-_b0Zb5]GXEeSAJZ_RSO>VA[0^.//5c\?:
\M[Z2BQL>\(VNW?<8JVg]A+EKHRFbO_E#.<<2B:@gFEXWEK.+/.(#-F@:cGd68LH
>/=H=-3/BA0MT18Wf<dKCK@/(G2QJ_WN58,Fd,-1.(\K\5I][12P[?T_+_.\X&S>
GB)Gfe+3Yfb37f59XHW)[d-INd5Q(?Cec:1R.M/KG;9f#Q5bgG.W-fdTLU3]@B7S
V2O<BS>J[a&GW7UXaSJ3N^OSX.):b>E4L)++=_;LY_eZWFU4SQ1Ef4?g.BRQ-_W5
#;DZf=g>aM]/H;T+)\>HDQ;NdLI\/3Ee5aOI69Z.S_)SF1M>IL5Xd#7HT09/W,;.
H&c>4>#aDeC5H0:a6--B\ZN&X.=[CB23GVO,J)WC<ALLc8W)4\de:JPg9/0.7]G,
P#+W&GV6VDTdU8^[<ADAAOaO??=dL<<Y>]+2cZ@CSX&gUCZ:^PTSJggMB&b)/SRg
aWaS8LeMa>8b]:@a?667C2A/X8;80eI.&@V:NI9GI+#.5IJ-;&0ZS[U(^IMDS\U=
1>e2I=:\LO.U:QbD#WG?7?;.M/;#_B&a(LUOGF=DY9,1N]G^JJBKBbbgI&UP[@)a
daB:=A/bQ-60\ODMfY]A+f/1S#,&\_8ZL0c8f<Y(+P:I2_VGbF<)[L1.O&ZK@#PD
@&P:a]JB_-L0[;SV])_=0M-.>IMJc(IdMQK>H5C(?XK)-##,JC79]NJ2Be/A8>\c
;@Z0/^@3ONTX)dJLIC_B1=]8=6V+?Ef#<YOG<>bH)3>W8Z;LL5V&eI34>.V(K<[>
E_TD8]X:&QW[IC9/,a>dg3MY>X6cc/?ELA53;BJVQOW^GUJQ;6]^N=D/EH(0a20b
_\?3_<-Z@ee..).K/[G6QHG]b(3.?KHM81OgLTAFGHW+A4>[]^0_CB/=,TROIL0U
1-UKaZ=C0P,].e\(R>?C-YQ24f<;b=BN9((gd?_3cI#>T-+=1,#W@g0#R.UB8Y&:
eU5&]&<B#HNHANM8]K0)Q)adJC>R;=a?D;eA-bSLb=N0ab]IDP5UK&.S-NCYT)WE
CdWe46Y>P^\M8G\(K[,V30L^MbQbU<aGVa?d&?V-F:&NE\egTICPeZ&6BbX8[G?;
Z7@VJW>eMY]J\Z97dAF>I57HE>_P&9JdU@LMe<S5@.eEFT0@SS=#_:W,JU?WFcX+
],G8@.eRJVO+aXa5#&H)5ScD.\TU6N-Oge;XVY4+=3_P19=8d/EZ1JQM+)df8.^]
1M-Tf.8L]4E<4CIM]E)GABMHF6^b3U)\.<+Y[9Lg#eVVX2?H:YSO1ag5cIeGX)W4
G8L;8:NI_0GU+:=-O3R1DXdBbbAM@)(UfVa:::UeA<g=5g==AG&de0GT>?@IfJCR
NMGX,0aLNc-D@7(X[gDT;HZ(RVd)@MCYg@K0Da-JCRN</MBQF)I:Pd+2.@/#Xa/<
B8bORCJEL82EJEZ+<MJTG^=0+b;\g^=GJ4I;5<HGMJZ;G1YeGW^1W5K2E=NKgAFA
f71+;f.869(MbC<]].(R3W(&N/&O/UM4]d(K,4gZAVU/JOc2\\d9<?NM,CH7\TbV
P9d0@8N/7)68(.V?.@K@(H+1,</50C@c2(GN7>0FYaN@HGUE)>eG44aM//:]@@6^
NIcL87X;4U7Q4SXe^B(F0>WZ(N1)UGJZb5@M\GAY:8-Ia[H<R[&:Q^=1>-W6gRUG
DF>QV]TO1OWcK@A7T^#e9JdIF]P1@\I4_4?GdQP0g<?g^B;Q31J8N+I@(<XJc+WP
W]RKW6&T-,?b0Vf(O7#7.d9<05FAAFKX_T_V>fDF:_:]^f^F8HJb06^5AG;(d7O>
fS\3KAQWS5<#TePXOXDRG+gRWPaSKZ.AM7_]OJ26.AXe-/T.gLH7VK(BAJ.A4&9>
fJZ;Ya^g2P+6(5Z67;9?HUc0@:4>JTV4<G\(86Q@198L/(e-TFDLcM/ZR,/e#Rd1
SVH44g)A+6#TS=T[N&4J9TSCCJ#Of7^c_]dYM#^g=7?M9-d\U5[>I>?5E9V+1NGF
c0&g(_KYd[762KTdLdBEH\gYGRd4,;=2DF>]D;<52<L7)W)4T)e/9PZ@QT>#aFa\
2+C16@b^\_S#;Y(7FXUI0-__E)UDdNbf9JWB&MeRLM@N[EJH5S[Q^\?8851\NC.?
dKLCZMLZTGFN1cE99SZ?Veg##2P_L,+A,g>Nf[FZL[)?2YaT3_fXW3LHeaF,5J3+
[,7]KM?-Z-QfQE4W_>=/HHSCKZf19=He?68\L]0O]IK-Reb)/[d&VH&,Fc;DM2FX
f+8H((V#d+8[\+S=SXaR6ac8;9[3YF3<&deU4DKTbf9N7V&(b4[820C6KPP[Ef1M
A^9=G=0I9d9]^.0M@>.;_)SIGc2C+Xf)?L=c0TF,B/UG8K]3M_?Q?O1]bI.2FHD7
.J85V<^?/Tb>>\&+E@=3LW;Z1e]bGL[<H,d.AURJ@+V#dP[_K#8?5B>R,_K)-WCC
08;]D[NNC-;T:QI@UJKeEX1f^21?Y\c(6;Z>12C?P)e&+R<M;#aE++0E^gSfE8_Z
1fP]/^L^M.,JUQP7cH\,#885_T1H)NVOGd^05Z=Y4RcB<d2TAZe,#)R\5#&3La6F
fQZH>/:0c,OB^V.8HEf]A2cW<fHGA+DcdA<FfMae>G/1FEQg#Q;IdY9aPT\_eg6T
G&7Q9fU@.U240;[=P=54Z/#?LC[c1N<M_fJc.[eX6.]c+dXg3Ze10,2((f=/N:RH
7]#JLB::KQ9LU>VV,JMf8-Ja,HQC<TVCAS,^Se0-D2eV=D\9+4FGQ0f#HV-:CO.5
W=7Xe6?.<5dSK[6bS<KV._JO0T\d<VEJ,L-K(#LR&RSN_,S37@Da<Vff06D^&88c
Z)NS[I9HNP1[I2XJ?NU8fI6-A).B=K\,#9NZR.>),PG&[0F.&EP+J1?N[8a.,Z^;
3Y0)68]3W)f-gYIa5ADE+b=69)^U41F+GG<f\??UCJe\./7?AIHJCT<^KS0/a1/J
O9N/:0)3RIaeSg2H:Uab9WQZd,URb=R;XIcQ@DHIc6VE?BUfIA:J.cI:c-3/?GF]
FPB;R]62:)(1A_5UD-:[b@W^GW7W3&^(/@2S#@[J&>U[8@@XXD<L]-Aa\C8A1705
6TLf&=)bR1<9O1;KSM.4D6,;L1E<U>06JDG,YPd9-g&@29A]XG8&2Z]5eF3\f#K.
8d:GR3_#]NDcGSG&>BDQ91MH9W,ZEG8UIc-@MK;.g^;9?=P2O/XC>\HSH_ZA8#T1
)bS997g(DHX9Y60&-e[(-OLX/]NHBW(Z>B1YMY0)TeMXA2ULK=.&RHA&(<B(0f-3
BOF,0](GO&<74aO++5MB^Idd1;W55EcU@0e39HJ0g+We+X3b72XfG0F.7DQ-cSH5
4D^7IFC\L<@5,0d7__PEE6>/g_@OF928g;S[7SX-H,9aTD;KV+422X?;.2:0D/X6
8GIaKZ/cZA\fSSS.fZX\O]>^/N\O6Z\ECe3S3[X>HP81/Z^EHf7=WF\V7GL,=NGL
W#A7fX=,)+7S]XN00FRUJU0\..0V]ObGaAeB>\:-7-QYI&Z-L^HKMBQgV.EPF=GS
e>0=4+_?/&O#UD;0C6CF^KQ(,K&_=WII^:J>b/GBFeaH:N^ZUVV_RD^5BG<6-5T\
5-g.E]ER+U23L@bA[O^ZJ52N?XC&OJa7BWF&I^XfC>IN:3RaSfEJ](C^O,V/c9IK
<@=:IcA+[DbW<)TaIE>Z+R_PE_@<D2.?[]PL[GTB,1dWA9&FV4,3(\AQVW\=/GKQ
(,<0JDF./H?J=@IPbES5-L1M+YdE(0;?]0OdW8c73\F]1dg^_/T0c1WD4/__S>D6
VUX#1d^[MM<O?M:(->A^QQO75-2,JXa=H9RITGaI=TDFBF3;137eP^8\.B?e9RS9
X/\fLOYKO,O9A;K0>Q:<G_GP9aH8>]D^g)Ue7Vfe;eF9DKG[D[+U\0V.]96K4<.D
@C?.[30[[431S(;##LQGLN19NUC5DD881J,GJZ1S#<3Ta[OZRW[]EU#-(RH,gYeU
KP#/eS.]e&HFF2;S=@8f3G)SC/JF7Y6.48Jd,[P8.c>1ACMDN2O42Ygd.WSBG6MJ
4bJ+&6VJ-;#f4CJ3a)&b&U>M;0M:1N]CAXZ;e38>FPRZFYA(>0XSEYP2E9>WUb3)
67:9P/>\4C,[P)f4.fP,1?bWSI^O3](R),6Qe(5_4Z.3/d&aE#OP88(T9<S[>LS-
X>c_D,?dfDQDAEUNO/Og]Z92@^[WRe:+X>S>+1G:.+8M]M0eC,GeJB@,O=RB-L=<
I=+CB>^=)\X[,L+FEO=b5=^T2a^a/)RgD[DGV0:/XNE;Y.fJ1EP^#S4B^UHc\_#Z
)d(_N+9c]e92U>QQfT:Z#g^YR1a;RBaf&WG3E1)#FIPOUfWKFAFKKFN=c;+=7)gc
5CEa^<+M_G/JDTKYdaUVeJM4(@]Y6=ACaM9_;3\L=]5GaVIHG#S1=X,-_/#<-X&?
#:2/LUZ4Kf]d->_\]#g8<)ABP90A9)7fE9@(C<A_+A#C?QN=N5K=LPHfWN.<=@IG
0S_BgJJR=DE:+#G),#N?(GC7gMEI8LC(D#SY<V#2FMUIL]FFB3LfF#/:QO6[C5U;
&;&(A-+]RdOWX\e.=UbJT.=8=M\64;P>3()V&A1RZCc6(?Z<((QS+G_,a8KAG#9/
Bg1/M.MB\4dM&B,^V]JQdP0Y(;PVd#9^<P-/54#c#==7ZQf;=:V;2?_SYc&P]CgU
_<U#XM)\]FAP#d^]GOO,9>;6;--APeN4(X1IggSCU<T?A,PNUEc5>(Y(>EV#c&XJ
^3/Z9c=e@.(2E0Z9I7I.Y5IHUeX+7&G0<KK;_,R4_7T[:-]/,AV3D6VBCT_1K&FC
aWTF62#6V>OZ_Ub:/VbOeSA===,Q[6[Nc)Z^Z-Sc=@=RIBN,@51#_(gZ&4R5<9NY
6;6#OGU8d?g(5[^YPY=L/[3PK7P#Z=Xf4/S)CU(CHe__#:MAU[fI>c:f]64;^BT_
0OXD/(_WM0W,DU4KFM25,A_P9L,G;\H<T7A&5b]Z^)MCM+VD0;)S/@6_7Y6#TQYE
Y#1D?V]AI1d1@>^Q0=OM^#+L>BGW8)>P?3TU5aJN:8Fa>BOB<2gJQSZg9f.==J#]
KQ^?I)2gC^:E/D6@8GD3H?_+(.,CA/YW[K2\D[bWGSIIfDJ=YHT/45MP,@\KF^Z[
BK72IbC9B<&3.&.@a,><:;)&\d.bGee#3+DDN2]/]1&&M(#K#DBTc8]7Z?SR_+IO
NDK70f3X&./<?GM.d7Q\YaA22/G\ad(0&0XV;/OWD92^EC9>:5;-A4VcB\D]BY92
JOeQO(2OR-5,Q>Y<L5LZe^V->dVUXW4W:Q+OPce:A&CE1C0@NMMgSQ#,7A<XdEdA
F?3C->KN=7E#^&4d.dT&S3:9W3WMQ?[;<WU0FaL4]aJf4@bH_;KEL5Ja;]4gb.U7
3[cI(f(.V<gK\QPK)Y\BJ+.09\Mf70]DI[]/.8bFZYFJ@>WVR_:dKUbE._&-T1a1
NO]^9PC9,:-be;,+03TGaEPeF\#8Z0KK#?gG+2-4g,U8dMNCN:8(\XNMIdPTO0JJ
_8>#I-V[?F<gO(cC#1b)HNX2IR.f[H;NC4A3_BZ8TY9fZMeQ-=K.=^KW:3\YHP+&
S?\L1[1LW:(D-OPS\DE<>Xb(133-^CYFf>.6XGAPI+:I1<dX);1=#e&@T>H#I/@Z
^_L)2KKc9.^R&1WH3PbR+1C:6[KL258T,\H&+1P68[;6]RC&\e;?5-P^e.H3;2_;
QJd@Q4eK<>0BT>=W1ML/[F5HN^>S>0[P>IF?5O77&VT4?e,6<a\M6O2OP_O2O<21
gV[DbTN//^gG14&Jg-9Z_NdC5_>f/8bQ\,gPf5T2H8@\Y;EU2FPN_AVeYZI[B8=7
+P,UM\@_d;SQ#3c.II5\Z9KU(?/gc7(D<ggE@a\N&>aa\O-<R@\+@LWQKGYC#-gD
CTGbBba)GMHQ@+4]7-JbP^,>a?60F9G=GQ_RXEgK+]K/PW&.-REae#[C#+9)#9T/
B:Q_BT=<4N:cHE;\Ta8,=5ZBH7;JT[1G[&]B9C]W?VBD@N.c(JNK-;b.WN)-Q9;X
D9WX(YRLdRf0dU_Ef.J6?ZWV:W..Ba7:G/Q0[+3,5N+.G>AG^4Z9#&C#DQJE?MfF
IX01O8K.+HQe\bJ=f5bAI)9,@LeeUCR@MU+YdQR+eEHTB1;a;VFWe/UAB+aU8c0]
Xg^Ca:Hg-e>P<8;D@14AaT#D)&eKWd68T,<2GJ;SCMH.-JA+W?AC-d2g#dJR>&CA
2O2XdDIH#.=S6dW0T<//bALX,]Wc)\)U/_dJ[L.#;X/Z((d=<4eC=@MOK]T?><Xd
Q>,KA7c[SDSc(9c(2/e-X5^A##470eGaf:@@;Z2e0NX-b.e3GbU]a8AR;c^HG;]2
U:9:S]8X,EdL2\J;L_4Y3fI)Q4Wdd2UFH7\Q4@+3=6II\OGR29g[X=<F#]Q@QfS(
<60L.DcO@L2f<P/^\bNYD&\IYKKF[S@1UEP\Pg-)8FTD6/BKdPI2YeFO>BUW.bXV
ZBB_W0/]>gW,E7011SO4-)J[/K5W2Ad\5@[b:aC-f/>::_+#7<\D[)[+\76NO5OW
JLE7((222F:J0[C4PW6/M#QbN#-A;3Z+3-(YGC]WK1K@J)LeE=FH<]6+5PefH73C
IcG;(\IB3K@I6fY8B98bc?RQ=GC:a^8-<4U126M5T5e&W,cPG3eRb2GX6M5VTDAg
NT&LR=g05IK@9\B7fY[U\#7WW34.__3BJe@<1,<+[9Pe/;:27dKeYDU?@5)#G(;W
4TUW5VbP<<C=@KW^f[UA<46>0a)AABIPA)=@(b7ZfHPT:a=f0a,+W<NUUG\F)E(W
A^?@#c4OM_T\/dO.]85#I\C]DgS^:UXVW[3=3ASM8#WRUMf]8>WfS0c;f.Da&T1S
PD^a/#g.?I:OO,WgFX4IWV]->\FFD03F_U1cXF(LBY(_3ZKVBV71OQPecZT>[gcK
f4VSWNJT5:&4T2a\8;Q;g^dOf7b2LP]5+RPT)M1bVX+1NaY4I))&.;Wb/50+KT8a
7Pbc4Q?\Z;.\2ACX0=UULXfbHQ\.[3LL6#(TJT,C.=A^+PZ2@8M97d[5,?R:ebJS
4FZ7-X1.SU/4[#12f(6H[=/^)RS^.4T#3<3(]G0?+U#0B4T,RX?#J^6I6bRSS/79
9,TfCMb@eFIa<,L?]_J5d/Hf5E\:_[YV3H<JK4WT(R[8DYUPSY7G1_JBTG#<&-fM
IR@<V-3W/YegW#fSb(WZ\9JE>F<[X5#L84G<C#<g8;aB<3<UR]3RQ>S.II7UaG>4
+c<XK-NC2_=bG4cf55^&:FNN#8ED_;5<L9d-YCU>JOaNPGZFZ2WSa^+.XY<&Q1_a
;FNWe0GQaDYXG<HOcR2J>+,eQW;P.aRAcdQGaLS_LQ4J?O\IO[F#gbLU@]0/?=MV
0ENOOAL5IX9]<eb84#]9^5-WG#L;(=ZQ(eBeUd(SKCO&\<JbT1(bDY3];M8c/e\Y
<e\>5R4((<)?M>WcA>MJ/:]IN0>5WSg5:C8Ta(U></ZY[N6EMA3gE+a;9[OY3U8G
NX/NI:NL.>7L)8fG3J=&D2>TP+VF1IW)G(:6)^3Fg@4TFf_H7@gUa>RVR)VG3a9I
68M@#3GX/=)Z@39(EN>LA;AQMY?]4bbZ^-Q0>;^cbM7]T(9=61STCY?QVE6?OZD+
dRG()S9;O,)C#Q_)dZ_d[R+FUN)F<TWV^cDNJ7(^0:XNA^.g9[IM4ZIYCdKM_W.)
.gS/Y=Ka:LGH8>3H2YD]P#;LGdT+3O5HT)&eL,P<D^;BQ:Q-;J?NC?+8Rd#R?2dX
C8CB^[R#fMNHFVYgUBN>O#3=EG>f49Z(eK]d_74^Y=PXF.OB+;UTb^))H,\DO7?I
2J6XPDM.KCGb\dX&c+C]?O0+0A<Eb::aEE]Z5N7,4,-+_d4.>LZ1gb6H_?V9Q/1e
X/FBf5UEL9_>OZ&)eDZK+P4<^K.DW#VP552FcbbCYFKPa&ZQAW=gP04]OdbaJL6J
91>F(X:3.N5ReLaV<:&BeKcJ@Z=FCYA&=C,b498d]<P[I#8JJGW-F^(=8(2bQ)H,
.=LJ#dN]>K>MLXe>GNbJGSg=c4W6acK=;+UO7[)^[@.\+/C(d:NB3SgFWY@EN.S.
]@.#V+,U+f(GHC/_a4[4+A)P<aIA[-H\cWMM^_7C<2S47HOeW>;M;G#S_1)X,Z0R
e/M_9AL&QDGf5@5ZI(XF948QY(-UAOKLA0Q_HgbRK@2,H>_M7d9T\(YP[bIIE50I
,Q,Qe02[O#L-5EKQ.Be,cAI188fF\G0Q#I5e(Gb]2KG+dEU]1d.YT[#C>CGQ8[D/
M=;VZEXC(+RE@@J9A/afLf5LBG@CIDN_g/S_JNSA[/92#52[d])_UXEF\XM1R,6P
;WQVd92K<UV<Q_1(,Sc.TV?CZ^_W8VNMV56HFCI),ZY9;C^^,TJGbK^CW50F?dU+
-6A89g431HR^Z(/Y5],.2Zfb?XPBLWQ1U=8,1a#.;.:;+QPSg+/3Oc)YYgX=37CY
-FMVNM8V;b)A3bZ1fWG^f08(Rc^-J]SVX)=)5[&E9gc:EGS_]QMeDGH-/.KU(e+T
:Kc<&UIB[TA9;LEER/>^E7IGPW<2+aX;+E7ZFW;N3I/BI)/FXPW\]bR-/_Q[e9/J
Q[,P?@>BJWA;gJY^2S.AOJJ6C<VHMeVDQOP+\-3-HSTb1b/PaAAN16:WZY(D3I,E
@+2CY.KR&EL/d:(3K&[5;>Lb#,@W_TY<=)83N_P=08S_],TR_+PTB@]5>.4+8#a?
eO+8B)8>DKW0;S@N)QIBECP7\.GIF^P-DUX.S?ZG;[7>bH:H/>Mfc_.(X>>3X+RT
.FNc.>GOa]ae;,Xf8ZH9P?#e;TZE#;DDDI4DM/6YVcJVW7+.XD\R#N32EIdO1?W@
XDYMW;TBTQIb[TZCD+;<a,(7\#??F2W+ZBfO=G0[8_1,CTT^(DX,E@fC#bbPfNG1
)/dT0e#([XVe3Z^H]a#&d1]KMe1d3._GJ-gZAcE-=PT9Y2Vb+ASA906B6dH[a4#S
f3CJ_/VE5I(KRYULa[BaMB9A@]\d?Wg?^1-TdI>J0NH[S)I?T;9IB4Z?TMBaLC\R
BFg<8IJfCEg+c5;L;ZQ?&25.JJQ/EJJ4cXAcOGA9H,L(aDa.W3(.PSQRc;WcUOb/
PS&X#O0UW>3:PI8(.?c(_L>Z&f(7<1&(0DQHOX2^JN7)?dD4HL/.S15W-]&+F=08
4#e[_Q>(a,Sb5V#Y6K3971#eG2N/F(-X^(^D[,6^#1d#g@)c^9a6cb_.FOeU[?&I
?dEL_fg8LN[WJ^bH;Cf^]#E/DNdQ]Hd@5VLb07a&>6?Ed&c2^=30REISc3]d/8(C
2WB/BESVL=WU,6C-5&#bY=_JVU;;_I4g89gBX)0g[c_)Y4MSNBD.G(8K1(G2.QR?
/a>G8)N,OZgIL)A=>T[NgaCO^eD6F<[=6,7DDU-Y[1\J)N4DBTdLV0ZQfET72RJ@
ZH[R.^eI7Y-N3Ka0CeGV][J>UHP]>3_T9[bcF<HNdX=a(K9&8U<MA_>Z-<,,M>GF
Z-FgQ(/3Ac24:7gREgE5.WPS0&>DOUd8OV9#CVJg=<Y;\X^dW3MH-e;6N@ZM]0[O
B@@WT==_5I^cP)L(Y/SfO+FS?)6E]IRNQd)2QLDNZAEN:]LXPW@bagC)9(/YEDJa
]aFcDV2RTYdY+bW1d.Y+;);:d7.#=5gU&(#?63/S^VAO@<;_0O\F12eK@0-J<I=,
>?3XXeC1\3YaH>g#<&U6]P8QC(\678Z0Q+4g9(a5,BcI;03-9H_N>S:A^=a9W7d5
LeH(6(B3?\3B=++=(Db\YHW_21K10Z,7XdD:X#DcKVf<J^78gfBH@-DP&KP3&^_)
1e)V_JH-O81MKP=9F#2f)+)WG<@Q-KPO@d5=NCEbEUVKXUI?DMH/bX07\ZGY\)(U
L,/<:#24Tad2(GEG4\EQ(UGZ)Z]UEab535;)X\Y6YDa:SO2-/4G@HZ.2OT(0HZCF
-P@,e7@#+N^XRJBEbE:6^6XD6:bPZ;CYF,T,Z6f3f_9E5NIO/aP3=<cR-&DH1^9_
6KGSK(2X2&OGf1T0FcQM@??7_;V?>KQd>.@48E98>f+HVcRBQc&E/S0SF7,L84=a
?R8Ga5?,-QeH&F6FP+e^^WLFL,T>@Z-<)(?E,:ca?T_6b4MRL61aG?YHR6dMb[)X
=LS)LK)IA/:VL_U#;bGVJUEWXd6Z2OOQ+T:H^M^W::(Le>DJ_J2=6fB<B<-0YN[8
>8(?<I4P<4;CD__B./9YR(/?2-R@MdVb8WYZfVN3P[UV1[@RK#5b\XQ5eWY7b<1Z
DD&;IbTcc&[:TFXaeE2+GJA1;T^H-A9S3IW58(+.d0JU(<cTOV(A&&(X(QY9=7)a
+O45b-C(/>c3/)#39#KDX^L)UIMO)@/7?L5g9F.Z06#HTCdC2(.SPcQE1+..5-0[
J]1bEV60OJF/^-QVB5@IWX54G)\;>FRHT.1/[LIJ<>?gFA6?gU<0W:0,:;L@,Oa1
Z58^I[FeG(e1)MJ/ZI6=.;O)_S_-\YQ7V6PGKCW<)]5=;VVWAWe(:WgY4X/+_K7M
]3c4_FD;ga>7e@D>eO5F:NZ2^e]29#E-GPb=HVcW]..=&fbOEU-ScI[SU.2XIX8[
J7FY#,;6]1^47<\+)U2JR7J<KJ:E5JTg/A3CORK@P;(N@f^0:Q=(B1SQ7?>+W1GN
[V7O+V)f-RSJ=M_S=V[35JcO8f/[,._fLV-TP+Uf;<4=7?7ZaG6b3S5_KOEVMb8N
&/\CbC@J#8-Sa<\\SM5P(/HbfYCf>@_6@BWHZ97TGRNLb#7N#7O@HI)HXWCVD1++
3B-F5c2#?T/G(be+4^V0FT;N\Q)8(L&L3eU<QBPLI6(IBL?3G,E8HO97g;-KdFW8
XU.7>K.X4IS3d.#]8+;W66#F?^Udb+ND9M/XU.CN/T(7^]BK_&c.cY2J/ROW504U
(OGX^I9LH>1V]L-<][c;0+0e5Z6>FMV>(1\D)RJB,E7>IS;_7/\P:[#4980=cNTW
E4WdCC]-RaRS0C40bE;FMM_(H^IK,_2ZQU8]@50Jc:fA]_S]S.W_.HR:99I#&,;,
6Ga+C>5ReX,aE]<dO8SUbe6/Q1^Qf?f][?OI^8fN^g06OOK9SI@I@ADBEb+TI?HI
a>d-H70&4DO?I#9V)<UKb<YZ+Gg1-;=bW\RE_^T,+2bVdKEb4L=gV5C@E6/eKWDS
;5^PLWNNeB[@=9CXE[/D>+M3[3_+=L(#W2M:25WAV\([_)d6C>#Xc;QWB9)KeN0G
ST]D,?P;I#T(G1@(+c[ZXQbA>/R=\U<8QfO2P7aUB6VbgO3/c[.CFaI^gTeL_dB[
TdE0:?]0N-EgAXL;g5?a?L>XSH]ed>;Bc#K+f^YF4R<LMEACT^Z,?<JdZNK<4@g&
#->fD_EN6Y2<d@&Y=HMULM:CO16PM0IH,CCH,GRe&VKMN0)-1H.(5(NJSMf_H]Ca
XUTN+VN\SO^;3e.),b7+Mc]gJ1Xe?b@I\2SUfffE>-3?;[#W@8:NZ>=,WMfG<7f5
)Z4BdC6c79gaCW--A<O?L:O:[RcASCLVd_-KfO2YW&HL.QB.K6-59Pd;@:3&J/7d
eDI<&a<?..Ke<b#(:^ZEY5@/TSg?T1PJe;-#SS.V\/.2S==U#U66\;_&f#W8;M4>
UAI3P6?#1;#9Z@P/f;&D83=@9+<SK&UKE8F])>[2G(N9C2,UF8LAAd#07g22;NT\
Q=6:</E@T-,6.gD]90=.EBB9AEL;W;cZPPYX3dH0[.]NEEV,bSgNEc/+a2WbP=[G
RHHQ6ZL?BHc]YWGQ),@QH_X.G,gQbD^91=_B_T8\@LO,T=QaPYY5-EUQZ2dgBMfN
ENMJN8[0PT853E-K,&=USd,31XJY6RPZ;3)J#1fL@VU=fD=aOS(FfY1YWOR[\<0>
Y+Q+Ze7AfM^C+5)]Y+a[(ec84D5?\U>5YO@HDc40\A9N;_LY<)MX&)TCZE(HOQNI
-/8TP^TbVDF:AI)D-WZd\FTbFJb/1Q@O7U=.\[_?QE;=(B<4bHA)f,8Kg?39MgLR
B(cFV1JCK.+L5N0REYU+a&=b^dQV(<.M-Ag5&UCPg=gBeH<-,g3L-HTRN.3K=4DZ
P;H&OZWG8(a1,IH5If>7;)@;2[#C)Z_:b&NNXeW3cUH>NQS6RPX&<<6[]:3;4A/4
@#L#g5gb53?g@6#0\&DE6@]JcA&4gYXIaTVUeT)ZCQ2E[E:UEJdgW7bIE3EONWW-
b^R@4/-dSJ&:_aaJ,><DcUVXD=MGNE@2?Q]bO8:W.6A,WEG2R<E1]7?9fb&8dRKV
Z&f<@W,)2J,ED,UM[/9_I.Q;GK(G6C(b(d9e[ND9WA\N\E@@@^EEF^6Ta.J5EJOe
]NKEE5DF\)+5):OdaF=Ob>;[fFaP]7)CQ@+UZ)VaRFGN:H2)aG.gG<L4JTB&(AK2
gUEb(-Taa&X0U1&W):-I[9[-_M^0@2I@ZOSA&).Ic:WX,a,L,.J4E6a\b9H5WL?A
RCOd7T/T3(Q]7V^OFUa+7]L4DZ/BTPZ=1-T9[HWQ:#a\/;?@Dd4<fDHQU;H8f05.
>#5QY,B8Scb4GP@Ub961#G(YVFIJ-5NU3gd;;BSR-S]+bgeE/]1#XON0V:ZZ\XSa
B]7CT&^+)UHGaD=X6]H<dX89U@7N;SF36R\LKLUU2]&.&-.&>6V+5f^(c<0/B;d/
eB9TI)OH5c\><>F,S:XD>P-O13Y7W2,0@,2b[H:K@>-O;JdL6.YE>2&d>J2W+EV&
-;]R&_Ra,9\B;2][)DDRRCENRO.E4AfQ2P7)R3)G=Y^KU92ccVK<f@V[@c.&?A#f
N(3Y82EROfA6)JaEHXHNE74Y.R=41^:XKPM^@?PK^CTcCM8)#=(XMNBXc@F-?CdU
?I.4X<G#<Jcc\?CTH&EI2#@EJ#HV7f4)EX8EHN9[VXg+8]Ga6dc/-NV+^fKN?HaI
O.=QC8]5(Dd#HZG_2Af[I33PBQB&BMc?3-F_Z+cReRGFD]7<BO6#+[.>Ya2WH8BA
3+^38G><fCJE_,(g5=G#;dI4=<I=eF6.<=,:<+AB;[6MXVF1R=B^0Jd8/bC=BgZN
Gc9(0=RV9+D^-Pb9_N(ICCCOf^S8;JdV._g,]JeP7J3PN005[<(67^S?1MWF2D2+
7.:#_cOW)-YY[WIYKF@))ANT]b[W;69)H-SFfWQRCgM]T\Z.O\J](Q-+bN4H1[)&
P.403dPYA-[ZQY;(9WLII#R^SB#;Z:4KULURD:NX83,BB5ZabHFb=W_GA+H/XXT7
I0>H9bIABG,cc74@3@X2c)d-3d8CQ&&>(&A:\eCG3^-&[XDP+\OB.(C9[;8d?]V_
L4BC/JKC&JX.KD\>Z@2?AcS?3bG]MEeK0(Y-g?D3/OP_=,d;<(>:0[S3KQ[><[F4
a^#]9LRaO(O_@Dg,CMP:9ME\dB/?#1,YY,DLSPc4=.<_?)XXM3Rff@V@-.d&[>DZ
RdPc9@_8U83(E@DJW#(?dGK^/HL,6/4ZN/]:\K@ZO?8<[IOXB@af)gaK9?0=OFY=
<_9f&[LV0/8VUb8bSR4&C3Q\aIN^Q7f;RJH:CfRG,W=71Oc.N.XP-9.PU_,JJU[.
T>FZ3J,C>MBc\,@cgC_PQU#EGQV+60d3(a@,9bQ/VEX9AVNa(-H-=)=.Ib)d)N\0
DU/SW5Y;/BF]:<X^A#^8K&+@+Q+DK/6f+2-PZ_=3=d_<QD,=V_S:H)OI<535#^@c
:d_bVK[RG<XKH);HOV21[UJV,H6Nb<J/+>WZ:5dg.(DW-,YFaL5[A]X5Hf)_,2g#
\L@<VU+TSO0dEf5_cVMENYCfN;VFdW+QP:V>c@<^ZZ3YTKM]2K[&TC<KfA63J?Y:
V41I7[<Cbe40A@_IJWbG>ZS&90V/[W,>=03e_[G5D.Z#ZC8BZg6]G@7E9Q):LT>G
T+XO8GI/a.K>cTSQY9/b&CEId+,7;DE4C<d&WGCNTLP);?(-;BL:^#[<(60XOR<Q
QG.[[\=g9(ZDNCM8]?@@-4WD;G/0BfK,]9&bBPcM(MLKUNT+.8b+Ag2@^<:^UO[H
X:(_:/4Z3RJE1a#HCCVQE69BfOcPG(..gLT>J98T^^SLI0IT(6<CJ78=_#Y+/AJG
-[?KI:2];\RF(3Ie8bcd#E:b(b3L<+JbK21AW27VVM]>J9Z)3KDa<RAHRHHX6_W/
WNKR0(fM9,^S5G56YcQ89REW).SK7b\b8?G_(/RE4_)&F:QHSS?HG6?BaLd;WOJ@
WfBO^SR1IZd3#gXecS<_OHF[0ZEe:Y(dJ;SLc^Z>-6AS:24OI;Y2[bNOC1aCGaSe
BCf76/>]4f:F.0,c.0d2J)>1>-Y\OA-bec-T8T,57HPML<eG(\[@FaaR2-O>;QMC
>WV<1;3FND@&AQIb5]g94X#[CJ4A:MZ=.OE3LOYX#^F7Y3?:RP<=_\Y=>#8fdLV=
1Xd;dgMaN;=B3X@fK[ODR5PfO4]Wb;gJFLgCbR=59Y6C(3a;[6(6_KbaST7\(3_7
Z3K\YeG+#N1K)C7ZSLHg.1+\16CT#K]636Jb[:?L)9<470_X<Q,f&/Z+ce\=0;_;
,DU5c<]2=DLZ]?f#7:<-XHN0E.DAeF0He<#I1M8+FBMfKb3F;X9,8IW7b;SdE@(M
^EVaC^#Fb^S;6\40T=fMQMCP=Mf.Fec90@g1a5B;:X2cC(?E_,aVd?cX+L;8Z<a&
fN<EK2F0&OO:3a)KBV+b?=LMV=)W__E0N1Q-/[OXUD>c4-_O@5M^-TY.S[\>5,.+
(27PPC56O.HJ5f11V=+2Q3LB3[3e7_&LOSfLPA8.I^DLdUM]&T9)\HOT,8=;Kg21
X4HIRYQHZd^EN4@5+2\=/B775gJgKXAG-T._<4@aS1T9e&XQO,QJ0ZbMf/NYVZH[
ebXTbR<>g\&A722NPEZ/DgKS^0+a14PNV-+b)TKT^+<K\.PfI>L#A3:B#Q2?,5[<
GT[CX>4Q:[DZ9E=SFYd]gd=8H\EZ8R_c+MJWG5FdPKOLQ/DX&PeATTM&fbE4>S+_
G2<2F>BeCQW>Y\C]Z[F(&b&4cgeYJTK9HE=11=-Y6Y++@W6AODc>.?T:,:Kb2YcZ
WBRdHP0cg/;6^(^>9]Y)>aMd3fAOO@XA0_=9].29-=)R9.RXW3aKD;-I75WcA80+
gOD]D.KRd)]\RN,NC/a^KH=C1:F-PLPJDd3759@X,TZ8]=OBbQ7WOD?7M.eAO9g&
NH8M_FMObT56ZDdJ>@WS@96[+.>U1]I9)NOHA=TU]R)(BOSe)TJQ8YYGJY/cQ2dA
RbY=;B3QSdfZ4CLg4-CX)7XKe0?.&/SSOGeXA7Kb7GXC8+5\=7SBacR7^X#dPGNC
d:#KEVc_>_ND99)]c+e9B_FQG>)SeUAM6W7,EO?bJ)C0RY5<T)cHU:V+;c;[EaW/
MN/bY1N2dW+ZDYT-:#WFLD-9CGL81/DKMC:(7V3(g?K,Q^ce332)WE&T]8Z=Y=91
bNaJ7KC@>T)3D^AKHTZZ\X:UZG8\EUe2Y=XJB\WeVX=(+<?0F=ZP2a9RQZd]O]K+
ASa76cg7IaBARWT[Lc)61AJ)-g7Z8ZT0M\S\L<MKb]4OC.P=V]:>57T[F8C;8YEH
LJ83CQ0gZ,8c8A->F&Y>1#G-87]5147C.P2YS<bf7ZQ2J6&O-\_OIK7D;()>&32<
-N+Z_37(37ES)T]LZJ1cD>U&4aH+BHMY>G.YMRd;.:&^T\]7#1GCgR@H:+:3K_D^
g.I=8&-6\U_,C(c8Q1Cd3-747g^+T59J)^gL+S?R2\NdPYAGeJO-=;@<eDadFRF@
\?V5@0E?eW\>Q#6C+R8ZAJeP7];Ca,cJJa2U4?&_#[LDf?D;\PDFdEX/DJ]FO(Rb
X6d3DT0cBFJa;AN:6Q0BR>T3QLL<I6UbfLYY(9(D_]P4&W#4H^_4a@^\e-Uf;-(L
fMRY?W4A]XGXd6(-B6)b&MF?50FX/H@4-_[)ME[-fK_NE+6F;[BYM1XT1C-a6D>T
AEEd_K]_TPaFP0B80\g<VJCfMfYg1ZQPF8=D_V7Lgg4-)77F;C1\Y,+SB\JcD,M+
&?3^?W#06fMUY/5UXOI=UVK1/G[;+ceR9ZUQTV\0d\.b,(L6C)a&#/U?3F7CO++U
c+1FD@(XcMQ\CgSbdJfCJeCT<6ca:f9J4TYHbJNf&XW=])>Q+P?JR-EgJ7U^6d?U
W\Bdd9I0\G#ZJ6D2=3^f^2(_ANCZ6):BFG5(0^YI_df[:#XRA=UD^NeaO8BcH5M-
:.O3.7ASF2Sg+YJZ(H1T7MLJ,=8I#aTae[J=Rdc2[KRZ8,Rg)5OfO?[8:CW>:f,.
gSZQJTbbQKgX,BKFY5e>bE;5.]?+WZ+fV&R)+<Y0Cg>2RJ2HT5BONZ29B:EM<gDS
M6BK=Y/.ZU-C6(CQ?7W>1HZV^#1KAd?W&GI(EI/;COdQG;[8QZ(I]C,XZL(VBKdF
f_<SMDE1[Y8eHC#1:_HXFGMRHRG.YC(f#LGK?2V0GMDMaF#]f8XEF+52cU5[EU:L
Z;g??;\1<ZeP3>>b56eL[f6&5D4=6PJ@)@+7d_dC7=,DS,BU..K^[[WN[W5GdM>E
X1KBbX@#gF/QgHGf>P>cU1#[^acEYX9e<J0ENIc\RM51gY:Q93M>(Gd]\[-7]5OA
XJP[5SWVUOHf0[5-&]F(:78?)TKH[PEL<5@1ERVRa])@+&5+7eAKe5KGFY83(;:5
Aa#_K3_U^cHL32R3G6&7\<D?]Mg49)8)>DBb4c)5040cDe3,RYZ.E5IN+>QC\^T2
e8.H2Sc_c#E9(A<S)HbT,a15R]+=9L(2XNa=75FPMb.<W[EH<S_68__Ff=<B+4<6
5e>FKRcO&4AW^YD:8W.fV8[b[<1W(ZFJ;.Z8H/d8<26C5Y\9426e^Z^&4)?WBaA\
I?/\7G.e67,8^\/)cAK^aEDDY2Y(U-T1#4]b/>]AE8PYB_G_15SHZD19+?<RP;6:
(3T[d?1\fUZKO#7V80\)DUKf3S3Caf2J(3&HL]=9RLb?VW/)dY:ZJ<Q7NR>.[JT_
eC(1=3+:F(XIfe.1=5[O<a263^TX;1)Id+(;T93dcYfQgYI9@0H2CD>H;F3ae:\P
[MfN<cX7W&,FIR2[7NW1/@D57?DG>V^-fRNW[e@/+gSTegAIZ9=E4eE@(-JM#1ST
RX_U1f2KPgFJfFCKF#E4R.]=\TWM+,aD[DN)JeRWA5[SUYG9U>\=80[GON^1aa3N
C=P;Te[cceSbQe:Hc_@V;Id<=2BP/]-B,VY#EO#<YZP9K9T38/59R;SL_:/8G-Ke
_7QI[-(?(F_[(B7C@3MV\LJ;ML0&(fF[K.WTe9>0WT7TH871VQZEZ?F/;a2;>]<S
#8(>Y<<?@0[+We[GSF<R8>22)XL-e+_cN3f_G\S9>,HAL)2A)MV)B:X6bZ:O].P,
FU+4K-c9Y2QGG-<IX6]1dR[dOdaPc?XT.9\9MSFLE4RR#D;Scg4D2aO-C;FR]14(
bMN[a6^IKO(<-QBc3@gUSEg#NY?&D[8^DH?&EKI^0EHeT(QLB<]Y>]RLZ@C1)-29
e@NS(-=EZf4-.4O22S9I>RMV[eC@PA#T2&/15\#Jd#(+KDMC(B&4]MIe8g@FJ<E/
:bO[<?B5]I-G_UdXa=D2GWaPeb);fB2\f8-K_B[gO?+>+23gY,Na^.QgW]6Kd:6f
L]aA?U05L/A/FQ\M#LL/<88.FPTI.gA6Y;R09[I,^/0dTY<gD;NI8.U]>=Xd:1G3
f<c?ZNYdWO,[-BM_;+DfU9e_<J<^8&B/KV7Xe09JQ)>Xb9bT.>^MgJb6dHX3>J;6
LaGCbPI61<RXM\L7CC:g2dJ@HQM3J:;Q&UYO&Nc8W#7XJI;e7UYYZ;.b36bY--F[
,[KcH:X4C#f45:EgCBE^;8G0@):,@R\1>d[^AH3=@?UKF0CgTF-@Y;&(MAGe^?/W
_d@](G+J?O?3CZG?Xb#aMI1=2?XB_e[^]fZ>J\6XZ-?S5PAVI/R:080.YK:&B-c.
G^XeI)Z.Y=3OK;S=YcdAA@K_R)cS/ad52Og3:>)/>;6+SMFO]]@TQNHbFZ3_CeM.
ag_Y<A9feN>c5a;5@FAcBT=:(?SbV=fW^1NPMFM/bAfX)U>>/AUb]7_V)2Sb\35W
_.KeYL?PK)>LE5I(<bE?OJ#TGf/F4XeFUb#[@Y/A41NG.\Eg+O?)d,,3-<;J&E@F
11VI2/TO5g\@5XR+DP/SM6X@eLVb;;IS;XSZ@0Ma0NfS1>IKNJHVRfS[G;VR-].[
f5Jf0bB6U7<JGB)7,A;VJGMHA0LKA9)2gP9ZDE_gQ;\d_T)549_JE?D8XWd?(A[I
VL.?(3LJ\<J;Z3BAIE1W]aZ4_X-20NJ,XSgDRUN\BdA]CIS?_bG3TP;VQ&4KJ6\D
N,,CTBQ@g65_<BD7_S9@7WDT\3],fHLg(LYdRHEAKZ8<DR2a?b0a>-0M]QI^CeLH
FRGOXUf4d<)V8aGY2Q7N?_cY?A>>BCX(ZJ;N0,VcNQ[VSO4-[8Ib:@0TO:ZPOS/]
&=;MD446e>C2BK=I4U??2UD.&2_&fH/).c5DW_LDb,.EI?I7@(Y8W0XDZ478QYdY
\)g>f;XdW[ODWIN+HM#GL:O)#Gf-cP4E-KI,CWPX7GA[[a;&AaRGe;YA^V-N5T.4
d9IO\/-^O>Q6e6H-,W]Zc(.EKD2PJf,<JePc1Q>\,&3^G;G^X-;;b@#b3FSa;ZG;
CVQBUOU(c14)fP>&GHaJZb6f[=]AP4<GB2fU.4]>91&;:Y39aF6Q]d=_N-</JPNI
6f=D+GN4fN8BCS/9\BS\Pe0;I,Q\8<Y3,X@OSe5,?L2]31U14>#]LDgdM<<a38Y^
THR6[YD>R^._?&cM4/,SHL[BTY_19&RJ.FN:559LWVdS:cG.b3OJ.E56DaS1RS33
UV0BGFR?8^@ZccfW38AbgCKabYVXRV,97]F&H/R96;2g<I[3#UYU7bDdAZB[g<Te
;,E4NHX8)<RQPI]=gZYCU)/;a3-ad?dPRP^Ag1[bRNT2X.VMB[VT>1KYL\ac4&=c
YSFF+F6eHDDT0C(e;4L2gAV(<UB0RTPY8UT<)f287:S]?a(WIf2^Y605e67PLKBA
#-BWUKOJ&O2^c26SNRE)Fg?O6#Dg^BGP]_ZWT+,E?,]&=_JNN04J[;6^EDH9f(Md
9We<b.?D\XR58EWM?G]F#.,3[fYT?4RbKZ9FT@&f^#=c-8ZKVGSd(<g+)4LdIDJH
&Q.b&O\XNMcG/SH38I#FVD&XMJ-7WWW<T1#]P_]NRc-JNdL(+QR.f^dH;0B\-e]B
>6_&d9H_)<)](7d\9I)&E?RG+;f#X[]+^Z3/9d+F/a=.AQ4DYN2GZe^-J@:TH>(a
PJ2?ZZT[3ZeIC9G1>GV@bcVAg98J1U394BUd>QFMSf)5]a@62B>dY):=YZTBcSBO
3bT?JC[>RU6\/BCSC6NKI<8)7NJ@?P\,4]dU^U8FAa/b2Xc5[g=e<4]RHe3OV,d^
5:aO-S:U=?FS,)[RH3FEf;Hd#NWZVN]fAPBVf?B./H&GZ4\N)22Da>69+eU9]_3g
7=bbI5XPKD4Z3+(^&@3,&Q+/068b-/bNOW^6LII3.UPgV+SY=F;D:G/+P]<cUDVW
BKEPa&@gF[::.#KS=AS[S^=EL;;GS=MCX+&XVcZ\dR;fVH<HZV3</;JK^\5GK/SO
cU0SHZWG:2Q5D1=b#T\AH?0HCM-)835cI@HI+(XBTFE;U(<8+^Q;HU/KL;;,.Ie(
)+CJ]<:aLg1EZ+A>8TfM3B4E4G0]47V/F1.bDA-Zd)Q9WQTdG6+:^Ug):D:^7/C#
O@bC(LGR4]FM09QMM,F]IG^3gX4BB#+A^TO\,T=>@X;=3HXULI<SS-K.5I3[EZI:
844R^b43?>P;c4bf0.)C[G&EC_c,9GVA#2>8G;,N3[/,e;UWC7K78+=a[a(=F9I?
C1Y+-K5:?aVgG_P&96VD/MO-7d)9C;EYQF&PQV[.cVE7M<7-AQANO][K>bA-3\_L
TI5:1&eG;c9ce0bC^@c:U#E-VGJRA]9Ia(E@D[@X(^L26<2\6OO_11fgV7@:&UKC
D=UV1bc5JeZ63NAOU_L-4\MFe;4Y4L/FeMdHE?WLR/:efSe5aQ<6MRK^:IEOIM,g
0,POC-/5[S-A]IRaHb@f93ag>/e>)a7?[e@6\<CX0QPGJBS[[gZ<D/QV(Q?:2N>+
UZ381UHL@P8HYeO;[0W_BW:HI:W:DXI4?1QP-4HQPF(&N,cV00=67]],GGDKB@Ac
1KX\.S?BNY:@F/b99CH;4D<V/J#9-PZ.-Ua[7IS?BU?Xe3WDIF24^>;.QJQR&agB
B[Gg-4ZD)C+XI28IBSDI8K1_NP6bDeAD0:6:>:S7#.G:.bXT3-QUgWK\\K\\PMQD
?H.U:,3Y@5-RSP3X#ZRIgF7_c()2D2F2W/Z/I]:^@cRA_1YcQHG1c_0-Q6H.#Kb=
>-VXZI/NGM4TIgVC-WJJ&\N(Q<8/EN_NMNMcV?VT#XA?aITM+I>)H2\DDS8E_X<7
dbOX,.1F=OVLQ=7=COd[fW9F_b4JDHO--<Y^g4?M4DEc;F;&0[BY8UN9.d?>BQM#
?d(IGJX.g7a[gUCA<dO7223M,&6\dfFB:5VRf]DZ2>d<=EW,YM#&:,Mf3Qaf(<EO
E-S?T7.8Sd]1PD?.>&KSe<,5a2-0S5A;BWZ@QN8&g8e1Rb+&.99^fH_,3Q2L]NYG
?U;]?;cSYX?Q>4DfeOC1=-TeJX7XeEW,LbSg2O3:9#R+b_M,ZP<Ycea&4,NHdRd5
=&KYC/PK4R/9:e@QA9H@\d.RO[BJ\\BQY;GOA7_NDdN1?>1J#T0cA0WbeWK5))f[
[TV/,7[6(da^[fK#:@e>XVWfG5c(GI;V>AD=/>[P7PX)+1U6WdG3^V2GQQbW;G[Y
I#F?_?A.0)Mb#Vbbc6Mda9U&;O]CH5&)gfWd-A2#:d10T^8HZ6)_CO+ASKVWA7\]
(DZLB:5b+F<43D1\L1U(8>#E.\(2D:DEW]ZLEZe^cCPGRd/&0CM5>C(-O7?e&d:Z
eeRC]9]WO3^<Kb]CRKP1/V-52VG@1?bMG0)AZ1[2gF.C=FQ:OLL#Wa1-XRUFd5Zb
-GQDS#WDW&AgX0\-S?Cf\R(=8V+V?T0MgTE2URcC</e=E@XI#B/E(W3L-+CQ8M7.
^-;U#PL[Mc]DBW6^S8gJ8[R2O)SV\a\dWC8-cD_C93GX</^@F<W/_8G>Pd&QVH>Q
32aH9=[SOMGHbc.,_W9UZTRR1gPY9[X4R^6;;NER^f:d7^CWfa>I/FB?74]T-9cg
G=2++[cYRc./96eCM8gcM-MYAWHUU9PP.2/HE4@\08gK-:/d6Sba6-ZF<&8+Q:CT
d>R/[4ZbgeZdO2X=<-T^7K<4<SLOR3V0:F/>4bX_CTd[gV[(b?=)6^VZV(&-a[^_
=PV&8(S<[39KcZB0Ta.?,5BJ0_Z)\/SL>H[C5YfH^3Y<Q+D,33.8G0@NaOR)S;CA
g#AAKEM-A)58c#J>fN>aRG30H#SL,Z2\S3XcBOeO&ZS_U=aW#.URA<H5JfYeB)3C
4gd&2KL@XK#JR8:ED[S/?MQW>M_=/Z2SR9H\F\>R@M.d<8c[d-8f>I\__MgdaWK2
@@;?;MKdf)/.B/+A&c&KCB4b>\#7=01&/_0-,4BN>+SdQB3Z#]=KGN6E-.EYA,d&
cT;2ID4[06;Ubf#YW<(Pa?8[(;O_a0(_-UM7bag)&9Y:^4C5/L-)U/;-3Oa,JA)d
2Zb.DD2X9daFHW&7M)Yd-.LFP]FfILd?1WGT&LDJPN33?g@N:KXX:<XdUDTeP63b
BC4PQM&ZT[;6K^2Nd^Y:ISe+bCf[:W].>+F2PTL[4f=&#2E\52(6K_D2<?BS>PBJ
aB950O+bXOOd77/BK/V_L5A2FXT?8IX5DJeJ9@c[M1D6K9<^H9H:bNLaVb=+S\./
>1/^a6]>@[D8fLW4HD054&ELdGMILb-JE6[I25_P#V6&&H@D1+E\EDG>A720#gTb
,c/^Y4=,3NfT6d@FK@ZY+0b(B\TT.PNB?.=M^:bGIPWP8F5TJC#UG]9eN0WUYP@<
[N:@1O^>/QGCS[.\0Z+EOSU;\W2CFYT:0JH8:VH2QJC=)GXETBAV^f63F(^6(N^\
0U4/@:YQ\=37@NYaF6bXCgE75Q2e;Ae2#WR\FT@SG1bN-O-:[X744WL)4_NJ9R2=
)+WSU[JBQ#WC,(bf^5CJ4Y(&:FSaX)D.V,UMIX^H53O](c?;R<ZH5_GU6d3MB==E
dg<gZ\)P2R1[bP\)@-a_Q1d.B\Q#=Daa5W_bQ5.0O^@Q8(K3#2VZ]<bQ)ZK<1H._
7cJHHSVJgL?5=>@ZO86N;(^2eC+@PE07TfV.9f##g7OGH,e93U)WWc4\?FdYJ0?X
C1P.H86X,W-X35I,<YC@D_S3R<?bde0T)^,L9?a8E(4QT>8SK__-0=1b(g@-DTDY
7c3/V0P(E#]C(\/,VbBH6QS&&D4;)^YC==<W;?BF?\:>#2N_N<GgQF8O2[P14@3L
fMDS93ET.P3,]?9):fWB+KP=OKHV]:=[,M9LUB#8UOS7J.RDYVHOCQ75]dS.PE8U
L1:c_bbMR.a6Pe_;&Yg@T30C9I5^U^=>012.R6=Bff_NW/+#\F6,QT][=9KW^L<K
(-7)M31-NGC=fS^2fgJQM)#f7c^N4MJY#0Z=6IU-Z@cGKZD:GVU<\EP(\ZK[.L;H
WPaJ[5GI9>g1T1cSXT(cbCCDZG:22_g^3QWGN.F,7U.d^3-V;&-=BL5,\Yd[4F+I
LZRfQY#>@gXP87:VE&\)PD;6<=1OL1)<C]H?^W6X5>-L(B@LDYgN<SM9L]&75VSK
#FM3e);LZ8:;3<CP?7^7Kc7cQ;ZKK4@,eHbA;4]KI?V3Y_+0Cd(ScRIaRa(-,)U-
(CfF<W.)R9&N<f@O<8_5X>JX?25AI2OAMDF-=7R_=TSKZgOUTZf:-44=-+<c@FKg
#L])a0<:R:QE_A=^L]\+#cX];1]&@;JdJB41+Sg8f;G1WR=b>QLJ9V90aF,6CW8a
XG]A1NO(?XZ,RK[Y&H>+=AG.:_EP-DF>XJ:WHT<ReYC<[.Fe?cKL.K]@b#/:R9C1
CbH)U:ZV.43)\;;2I<cJH#5cYa9E-P&cMdT_QNd79P:g-Y(P<;(A9.Rg5B2SCGYS
GPgIKTG9.(N9W_K[QEF>>]_SF^d+R;)F(]2S3Z.Hg2U4\L>YT7Dg?ITb:B8<#gF7
.LVM)e?^4D7BTY?bGYH^I3BGf7-,Dd^T4Be[;;#GH4+.f?VRV-M^T[1dFIN_B>WO
WC8Z:cXX-aFY+5d(_f65O?b1S)a78g\21WY1A,H.c^CJbAg[^0X)2#U:]I0-cUaa
EKHA4I+<72AR+OHQCYGY+:T<bc?MY77B^25fK(@Q@S1c(9T,Y^FD8?IHO6/M//P:
3d6[ZAPK&1,;^C2E:P1gDZ;?2L.X(<AdI\JJ^GV#69gX9HU1^ZX:K7eM35^CNP8X
;=b5f:,)XF0+PHS62cV?eNCcUV23KY7#^#TMTYC>DRM1V-L;N5ePWZ3@M3RS(2--
ZYb-/cABUGYKdb]@\]:#P4M-LVe_JLU=)J,\f;4,JU<)\dcNYI,1RX4LGN/eOAM.
Dg[SJP/GL-Q0OX58G@4BC63ND>2.8S2bANB++E&3A:D5I?T,YC@ZWDEZ,(Od4LJ:
D0F\e0A/JR;H-EP2a4.KKbXCZ;1MgIO8S9dLFZ<U&A1a]JU<_0D1fP-FLXOML,Q7
/__&A>J3&+<V5M6L[T3JOZcGL9).R7Lc=KVD5_2L_d8OY,18d4&AB[3eRAd7Z/X@
[948Q@YN>Yd<VYQD,P<BVHAM^(,&GMJORP/^AgKaN<4>b:TJ<f9QcE_I()ZWZAJH
)fUH5@H+<+dQ-^B<SRWW1a/eV#f1(N&9E]H)Aa84g:JBZ6>XQ<>C4O@(&f19(YV1
XYY<?_5)?QeY1Od0cV9XbLcFG_>>(bD>_D?f:?D9MWHDF+^04P1DB5=a3g+fP7)S
_g-KF=c8S@[\f&3^M?VY\VM95NWPea-A)0/3&9GV2aDAR.7]/\R#CKb-EF]7[L\g
)K6BX.Kf[(=<cQFBBSecbg=E2R#agSPE\N2_AKUZSEge2/Ff_L+e4<&/_JJ(>1Ef
;fT0@\4ZYRJ(cMVGV0QSZ]7QMbGV===bDL5HdRIA1,0U_F)_BF@;P_90JaCT&?S9
PYO#K16SCe+BBAF;D?&@>;1S<&K?Ba<:VcV;Y^E3f3@YJ@^(^9-WXf7\d2D3S^7S
-D\67A0-bF7RKZW_Q0XZ;N]:DW.^NJa26S9DD),VE,@#^CA.IK.E-?g@gX,K39VN
U58)&e+70<KMgL(P>LeE[(\g0M7=KX<(V=R\?DO(HO#M-JN20W@#A+dgOLS(2K<\
Y<&932aB^LG-O<aI0G\VJ8T2bg-TC()27c,bbD:Hd2^T\_0G:9CSZAeBEP7O9_DD
]]b<=DOJRPJB9]CfJL97M9E1dS@&eN_9-B--7),-<M:@W-N1-6>ZGeFW]@TBQ,13
d(R^8E<.IC7.12gI\;ZF7D2D_I=;YM&3HM]4VJ@YJD?@8agGXZbR.9a<-H,SX;BU
VO7^7X3]&Oc(dR1Ab)5&BKP0NFN;Q^TE-7(>D;S;[c47[@L?FbB3aHY<GD^5J7#S
(V&6g@#<bg(A@/RN;DIe\K=2-#]C#7XT[Y,eb>ZWIaU=^KK:e74O&VAgVPcC]UUf
Y]5Q;+VU8#Pd,1B1XI-Td\OgZR09@T)3,YN<U-RJX/YE7L0K2-JZ#a9<EC=e(<2:
)[?EQN#KL1Q9<A+W6TCVe3cFFac3<aK=B7.g+<B7b=U#_/?1-VT\0@(L&IOTS0F9
ZBSd?P9e9,L;H1.@fX?=e02:]?6Ha6U^.M+)HIE&#C,baVGFHaUNPI[OeDa;cceQ
ZDfQ)fG]4HT)-DT\VZg)XSX\CT3C8(]=)Y+TM(SPJa_6JD9;JVBFgX_=8/(1YU9D
25ABNY7CNP\c@TW_K=4cO9J<S_Y2?;0DcW?8QP=\A)_X0AO5)C6QPOgE0(LH<X/)
/d-XEe4F:Q-3I&/3-8Ig;R[JGPGa;A)R/,7aB@MUG0>/;M9TOEFb13J]YI>0II;?
ZK:GG3NMSD/,GO>R+P#E=de\PN3-W_O9A7gUMWe?>+EQ6NP4,9fJ<^1>&BG,]6]O
U,62eYH?=WE,ZVC09U^<U_SN>YD12DDg.f9ZGN8JPX7dGcI-Z?#@T<KI2+&fQ>&=
,B/;Xg9gP&Fd57f5[T@6GOHD9&YYaU_7B>c=N</_^;;,7Q<gD6bARdXGf?BKBYJN
/0#-d5=8\V]#:,&X=+^<3R7/MEe?BSY=[,#AZZd4M8E.0Ed:N&FHY3OT&6gLTSRU
D6,S.QC_c:Q-VXYU4@JIGKMRQ&C/@8WK1F(NJNbYaT/NJC?U(QUCOTd5GVTRAKK0
H(W)4cLE=BXg87R1c?fOP<>c9c9I<^2R\OWTe/@bI[G,D]W](LF<Z;?99JGgFS-=
WS&@C?CUOFOJPVXYW^5#W3@:c#,Y0H9TH]U3eM:86a1[L>I9Pe\\DG9>6[S)?V^F
2Pg^RcW67ABQSZW[c:THd7cA&[Z_D5:\Y#,-F&O9:;0_Y_6W&:VO6/_bQIOX&MI1
-1eQ^1B_QI:dC>\:,QKK\:3TSZgI^c52M7b[b\UfOIc[)JF)aZ]/2XGe88CC42Me
32LLQ6YEXfO<3F)LbB91+/[^B<)K--QZH7<NACa]_Y[.YT3gg,DGJK5#:UV5D1F^
D]N/JA1FH43Oe.TR<D>M3)2<7fX6R/[(2bE;9(,17OH(gW.:>cJ>Tb+5?[5egeSa
-^_>MH_I])66@(]#IYad&&\.^6UG4ITCDU1fN&RFL@ab4GT._5^]N]+=^R+BGde9
EAFW=5@:QJ2_^,/4IT4CMF3F)>SH&SI1)KNf6\M[^g4S[gRX<)d+D3a)N\<9O4BA
aJa8K5N1XK?E[>ZP.O=&=;J@A@LAOEGIYO&]#^5J:)>H7cPU@L@H@g3^=5dVRO)_
1)E[3)^24N#OTcT]X,BH-25/URCe>1IGT=K9LEU>).;1;7@D._OIK#ZYS:\Nf@[\
]b.S:(eGa+Q_U;LY8YR:McD2[0/I]+ZP0,U_O+F1N:-<IJff93OXFf[S2,UZR;_^
G?aXTXY]@=.THJ=AH3Q#EW@(]F9:g>XT.DN.A&0HUcZ^fC;Sc=-FG1SDVZ7Ic5GV
NeEa(<+)3Sc4GM3^WJ<bVgJVWFQ@]C<>0f/FVDXD+0TNEWKI4c_Gb&/gAbAPR(FC
YBaVde#[VPH(;TACb[:>D5dT2P,YV>Nb]+P@^QFTZT:-;=US7)g#-&U1QbYRWE4/
U6U3f+5X,[4TN\-^f9&I9:V9?&O(3bQe]Ged]@79T?GSBL.<?4;N\HHTHb7L[HZN
3efO^:F]/1P9G1[H-#KTE.5Y)C5]>,15BAR@8GI1MO?;AaH5[AMUF4<K/,KD8KF.
&e.CS;J5:ZG)<SC)6M^JO1cV?-C@D)ZME<3&X:f2-IS8R\XF8G6-;TC0,9Z,D\Q]
&-GdQV_gFY,>aR^0]&8.Bc5I582N3EEb)2.f7-SA-.:?U_F1DRT?=LZU?b&;S:\L
VBPPW]TdD#V9(@)FEII8?KG3F/LN2Z=LAHa?-L(<88d<7G+RVAfB_P/[B&7T1D]#
U;YAd.Ja0@4@Ca(YQ[Y5^3EG]Z,[,U>H(TQ2a/I-SX\0DeJ)ZPJCC5#P;CBDE4X<
N]?,_f(5JA)6I3CF#\VM3/.OJ,91=CQEN)a8/==N\(2a\N:7gWeJ-OI9c1Fg9JT)
>&b:,^&CBP#2SZ6J89MDe5gGBf)KM8?P;-aK.+_&L>D6Q<HLe6S06e1W>@IDN8\]
U8DU=6-<A\?AeO7<e;;80QEgNNRX7U8;g#T<(24c]HJ;FO,:8bS&-T&1:a.&,]Q_
cE623fQebK()>:K6af/fR678GZfa76Pe_e0EFA@>I0+ff+GCFEeZb.(gF,\QXQLJ
/W.;3CA@)?6B.43[^4Vc4=M[fHLd<APP8UK+_&16FTTQ&J6[(SdSW7.S9GA41b1g
N[c7:^[c#;FaEFI9KA]bV-A_RHU;O:]5E^B7.<dQ6cYD<])c:#.@/S#Y_I?cKe;5
D/GX/E=M:371Q\Q;RX14B:KAD?IFJW2,^J=#M_DD5HK0b8WR4LOR#A-W?eOZRXf8
NYP>JR,G)2_HAIA^77>Y=<aI^HMB9+7;N)I-gVE.LJT5:L@,W3eANEbcYZ@+?:_g
a&X=X7/>?54,AQMYW\0Gc5-S,[-T50MS(Rc076>,I7EB8,DBU9T/1WbfNg8fR)-Y
_VeBEIB.GNI=2@g:@d.SG)d_ES71G6SW/7:=Y@TBQ_\-S.=f4N.@R+..Ze7N3L)b
e52Q(5^^D<J(d8c9EE/W;U.];.4TdTK8[;S,AcTI(R+P;>Eg+7e]&T;fD<.,a^Ff
D9fT>:38AaM#LO[-0bNM2_]M>5GZ4Z30cZ#>6=&W#)?a&ceGK2>^SL)]2He0=Ld4
QTK01RHH=(G,73Rc,J+1:-_>&X)#@W@2Dd;P/;=CScEANf4Zf(I(A#5OFMTG<-Aa
\GRF(.6O0<2,[+FO?4\B3#_BO-F)eaHBaaIXSY?Z#[2W;:)YVM_JD+>9&8LP-R=(
\B[,IR+]1-=^]M6D(>Y9?+QNPIRd^fFVg+N.+(@]E=8A2Jb?)7b#-?3D8QR>GXJ1
_HL>D/e0CG]I@gZ#>;WGdW9BZaZHDYcSQ?/1W3M];CSZM(5\MV.0cO+6^III4]94
5e]K5VE#4H_9-2@fKgC&-Yd^D#5__a#8;KSEX+NF#K2gG0(9[Id)^\:+I4K?@\\g
5P]-HZS<&L6A2)P6@0U_OIGB\Mc:(gK:G9N/R@=9[F9&Q6Q>(:/&>g8POIJNT[QB
JY.^/b?M+;Ee8D;#0IX&O?b:S-8a3&A=>NO61FU7ZKB_6\)g;5b<8F&aW#N+:2BF
D&6@P.YR,8@:]N+:YcCV^fNLRRZ5=;BSC@9W^K68=SGN^@\Q>EY]V^^1\P;X3A#7
a\bTIEUZ+dK[DN9&=W824fZRI5(gfPOGf+HAbW\OTL#;CG,OPR1RYZeG;X]5N.ST
E:cYIH9]>S6D@EA]V.L[;T@#H#J[c8aY-DE:AgGZf]HFR2W?;+HUTe2+[KCdZ5W=
8I4N=3^03df<O=4UFQ=:K&H;TYG4^Q-\<J[=TM(d[YD]0RABB?M9K1d]7QULUVSF
#04QAU>:(91A)AR(Xgd.2F[;a##5^9-Y52+IC:g-(K22UdO;M?NdD3M&:08Z)BS8
@YZ2BC[EH2OU+,]=:(,>fd\Yd(G,-\JWY1a8TCWU&OF.7NTU\VP1>E34R(MN&_a;
CYC(;a\([-XLTa\#e[;\OV8.=/>I1+S10Y]Q,NLK)-_7^.93PGOK.+AP/f/M:d1@
;1[9dK0QV.?>,_S\/05Wd3X==[fI]fH#LV4:cb]\UW#JS>F9>ULg8I2#W:>3D2WQ
_X[-KR>9-Y?5_0BD.&EV-Wa2?4,)6UU2AOUfcY4S)\3OBf;6D\c#RP4T[EDD>9fU
FQ9WED.f?:QSedHQ\#Z[eHK)dT>YO)a2dV+0-/aM:,;0#KKI4.T=L3.g_S-3]1P:
HNS,60FP@(Wb:T#I64N4g79?Bb))/1:<dMQ(a-ERcYTA]a)<YXd612&@@^O,,DJc
-F(,0.gZ3I9NXZZa[WO]3^8)W-0[L3f7LF.H]dQDF];J(<#I#N+)\>?&5<^Df,7G
&>G<FN<G::4eVU<J5QPfa,/[^-^c?<83TL94HX8(<R?g;N;ZHMXZG:V4G2;(4dC)
)a6@TaNdMJ\Ze/WV,)2VL_RVOC5ceN/&S(SP@D#1_(T^K>g>6;aS21OQYaQA7HNb
-7U,f@9/V/0,V9IBGC<VWUECCcGB-AH=5K/,K6WV>fCWW1(Yga/84;FOW@d_FO.=
dIUOUCUQa@G<X\AbKdAL(\Ob=,0Z0.1V8@fSK>H9Ye80F<TZ/F.;=KQQ:N7\BC>a
\D6OcQ24X=K#d8@&SPFG\36Q.M2+L+N4)>I(eg4NCWf)7NA3LCLML^#+2)?B8eSQ
;+K+6.8UJ[0#3bGCCc@>2eXBN;?]N;8RF:E5Fa&Z_K2<W&>6SJ8,cfg?Z<\&I66>
74T5<g(<+(67W?B0dW=8Ee+->6Ae=M(N@7(D/8We,A7^G&cMT4ZWFG??O#:).]3]
Sb>54g+4&:ZY&B0+,GI3@:SDF<(+>KVDM6:IQ?eaGY=gA=;<S:>+eD=T&,Qa5/--
cIBE8WZ@TFE+E3Y)HMZS1M]W=XDR]-(P:X1d7RYL_C8]?G4fDga>K\#\T=#WI7dH
1f9c()POXb_&0]._c.?2Ha>J.(_?/-E4H:;HB#1[b;?d/Y-?Z\[a<=]bO3d2Afd<
=X1)cAP)=\\[f7NfA0b.]::A>4@,G8/4K6fKHb<K@@a9#Lcd+V=J7WDBD/UJ(_9J
>Z@D4=\2,(aP<AS>9,N^#^?7&];0_VR+<&6JHI@Cc@[g,YdV<3V2)SZVF>C,cfI-
?O8HSJ<CfTC6#_36E3DL5#YbTJ@F_9^BA-Z6c@>WgM73Fba8Ca]^&^K0^Ug?[R?=
-2L_Y#@4BKA#cNZ#4YACA)9J88E0@@2+9(1QL>/8XCIGV?4H/Re>BRe:eQX3KL:L
9P,^<b-VTK=L>0a3:_eRSB^_d[&;fE:\6H,U[/0Y)QPO5HZVbcZE2NPfA-d,NcJZ
GL5.@RN]gC9dT_6>:U(6fbZQ1DPd#fJ<5N?1730R]L:27V>BQ[4]^_NZE#B&fF7.
))EQ]9RKFEc+(OFc;8_T2ZHC3G_Lb/(@6@8R1Dd?8OLXeC0C3ME\L)Y=e]#]b1NN
4+28H=Q&QL0]b20WF,^WBJ9L:75<C,3Nce@YO]0U0_++MO.:[Q);Z\U>X]K^<PIT
+9H8OX2;6MF1/#eC.MP&RaJQ0LQH@YGGF_.&W4B?L1FP#Y;Z^4=N<9cdVZ?5C25O
W8e]LDTT2#I3:=XM4fOI(<+4EI4GA(:=MQ4(HX,A\,2TZX-1IPa5-OKUHa>5UOP_
cAWW[@a17D1VJ/U>cUdHf0.d&/=QXGN5I[_eP]W&=+._58/=,F;H/4RQG84=-bgZ
@5I5RRg)<USL,bS2ZXGagV_4\RWTW=V#MHIW@I]g/a:YDQg()7.f3MVg&-II6X^=
9-DF,^V&g+cAV@T_c_,+B[JY(#OFTYWLRZeE<9P@K@[3/3a.HK52>0Vc/81.Fd1.
H_=4?QBJTU-cF6H0LHH\PA0(0fMR,_T@Z([1)WS<P/Yg3\B51\#e,3f7fMCc_Z0g
K@KBc9bD8&Q@-A\P<fIK)(7@X(>CMROT^L-E(5WH?])<4YNJQ@@+77E77]/1T9;(
[d/eaGT6ZNX^M/-Xff\5&?/KBAReV9W]7J#M5Df/F(::F;W8;7ZOQ>ZXSPBFcF=K
3_YNENQbW8<1->N,SX^R=cJ_-](.L?-WR]B;DYgCgWA4&MdG28=27D]5QHY--CBS
W.\42OHV=W&BMG>;97e=830#X;=6B-O@bIA6aXLgSMfPTb&f5.Dg-:G9[,PAZ;;B
eOY?a(J9+J:\I:Z2cM18\M32:CKbE,=HI0M9<PAAb2BF(_\]a1-QK&S>UXO[_a-P
_g8^Jdcef(M+NV9CU[[fc)Re^b>:e1FaJ5Va6MdP^L>P-^#I;b(4bN<^VVG.GBSQ
G3,UBN:NJ\7X,THe7EPL>;HU1S)?8Y@P99PV9]4)G&;@/3;GFEILJ1F1c3@24I7J
]I7U0TO=O1a(=e]]f)C+ZL#22966JSE/WOW<\&ZJ7G8I?3H138/2g5QEMK@NF^G^
b(V[S#2F;P=7BNIY_f\IgZTY81c?-NO^#4gBJHRGJbb].bJR]HDc=&\5^6RVN70A
,WF0&0a^#S4F<MG2ZIH=:4^eaQTfUW7X?98(/U83H;;8]>H;M?OKB?UY3ef0;YME
8OQR@)AB5K7OVJ6CM_EgD7C(=7F#>g87_#KYK;IZ?6/BAMXV<O?SFNb;BMC88=b>
8b,,fW@L=\&B,bB-Cf0500?f>T,RCe)<2(C33Y[)5^L;8RD)-V5RI]?:R;BY;Y7-
0M/\Z7;AV+Y26?,K;2.O0/c+S<)^SYV<T(HUW3XZ1=_JW688/7=III]#bcgAPM9,
L8eXEP[Zc4YC<3;7EggL.&+b3dHgdL,&6O1[P>=-=,);4YOGXNa(5(>W#Z>ET(H6
DMMB[Y)3RJIPB8F<YYadf2/I;FC]3W8ACXD2XbG3]g\:_G6Be+E./:DJ:S[8?f1C
MeRH=U&JY7Y16A/\7@1/RM?a(II2I.8G+eR\-.6#H5\64I8P^9+<)CUXN(SZ,10E
U5E6LJ3;/J:5Z9QPOS)_.#^S33Eef^_E9XN7/<S7)72&QgO0?,3A\dKR#6^[@QIW
K\W5^0AUA]b=[W4?Q4bBU;FgZXf))YcLNH_aVIXN\6YEde^DaK;2eX#Jg0c[.?4_
QE?Sb80B18^TEC+L_FE+ZH<.b/AJFN=U\Td9(1fZYFgI@>9(\^d^;Na?_^LAL#[5
=MI,BVMb\a.RfV0C3Oa<#fXeDc^[.JR-3>3+N15T@\/U&(QQ,Y^FU_&e=7;BS<_<
=GCZ<]3(UA+1/-V95:(XQMC[PURGdS626]9HVe<:?(Cb6bJ2D^,ZDc]?_/+PD^^(
U2a(QMg56T)c&A2:7HL8eM1#e6KM;e2^#UC:(;f/)]dZM]I2O+P&^g6ITAb;Q(2N
;-F7&.15R,YD-,35[D.ZbJBf#8P:@VDS84YH7a+^,W=bL6@^BIT1&PG0Y>eFN(IH
eQY]?CMOfGS=</d1F4JI7+fM;&SU=YAJ^9b0(6793)>HQO.=5]1N6LGE?R]1cLFA
D@ODHV3=?5?7MbaJ\2P#T&\0Q:O=ZBIbERJ+ga4^1U=&,PdBg-]K&4,2?U,HK;gZ
f/1&dGS)A28eQ#7Vg>/XKM2UX2W;AN4X:5c(0NSVBL9(cH9XK]bVT\#N-gb8O08(
Pa?:>HNH[WK[Ae2)/ZUK)SC25Z_.0HJ-5(>/1T,XO[2LC,[P&e2D(PKEJEN[#IJR
)4g-VJL5:QBR7,(+;/8.U4@8XI7Sg)NK^PY5)[Y&g;R_\Z,]CbZ)[C5W\/5SS,AO
?4S].S>X]RSF0?+WEZW7L;ea+_=]8)8BdNdQ4N4-BT@@2KTb[T?Z?7Mb.[LN&J;R
C<c/CgPJaTaW878#MIb8[[Qf(9O4KV+R1)R6dP^\>La=@5Yf&AgA@9a]e;G+D;;0
Qe?.&9eZHZM>98T3^0H:KAFQ+G\0@(_&(dC]?B&]K1FeWAF;+6:UMPXBPS?c?#D@
.#TR1HX_XM/F^80UUcF&C/4+AN1^SRRGXNdSG#\g@WD#&9e1#]TfMEFbO4;7FQe>
1,5=cK3,NU,Fc^;QYU;9K=:F2./G>H>c4O1Ag\-Y19U9HD18O02KIWJQ2gfQ7>Sc
EZVPPETFJB1CM52,JDbd<<I;f:-G(FD]FI@AK^_b3B-5.9=EJ,:)YZ_EJO;CW#JU
>BR<?Wa8D:K^B;TUW+#J6?cZ35G(6S2#dR9?MIR3c07Y/S;QOW&_+J<eCD-G/1N2
4:(-0eNNAAX23,HZJI&=]<+#R5;E;AS(FX+\1>;ZFZ^VT=g6B4a8g@;F&;(@W0T1
eR8eZgKZX,I9XA,O,1P<?aKMVad.AFSRCAR#SF<Hfc3WORIDRbPAeJ-a]Jda@(56
F4CY3cCMcB17Q7^)A\5,+]:S9gU57B(Tdf^I(B0b8/=?)KOUAQBUf3Z&F@]5@81/
Ya7&=D65eJF3X9VPc[;;]4]+2^W.2X>D_9EB=ONB0^9CKTb.,)#cKL:SdOR14+05
]X0gMMdB@2J3#O<V1M58B:&aJ(b,1;TN,2-V,AD>eTD<gHg-^WOXY-[ee26#.4(X
Dc;6C5ET/HcRQ4C5dScJ?G[;bHMO]=DgMN:GL05_O<dB;L6W04/T3SAF<]]A\D7_
f4cJ1Y7/5LSF=ONT]Kd]BFZ107/e_#O8#SEIYg=>#9ba=+8.20N.79\[VVZ)G)#L
B&>8.Ac4+6TL5/;;ZOZ\=<Q8I]5Q+7.OG]S6OU&>L:C]TBLXDDdGfeNb1T.B\a89
1&L6X8A5O73H/?I..+c.1af@H73YA#7G&;+CZ58]BD8VD.Ob<4[;.8A^0eHQ4DSW
E:BN_c+^52&Eb#T=,>+?0]J<CRK(B7J,7F&-;3@D(6PI>-0]>T5J&c[QbGU)e@J0
d;=_O(S9L\d_^c=dT07c^8HS\\Z.2M;_;6_Hg5).De+b@4)35cP]O&<[G6I41S-Y
/+O3:DE&,2-\CCL2<<7=J#.:f?cN<QLAbgCf[a/NT6O<#+XF5e_8f3dN^+N1;Y0M
GQ59=5C8>PVS;KT:(JcC>O?:NGG7R9TPR4&L5bT^a>e_6#ZV/^.;25PM&M\]d-<\
1KD)bg[PS?Xdd[0?&Fe9.0B=\fM-b\^26,:9A&63EZ\FKMKR_?H3H0YQI]<cQNVX
[Q[VWe34]22>#34^P+JM(_B(+d)2R@.H#PT_QEW&#f\QaAFO402W#>\=O.5C(EBR
PC2&agYc4]<99\dVPLV4[0JO66aJ[ZD4U^2FFbgF<^):N7NGZ3G4)<\^LP0X]e^3
6VQ,aSI3c,:JGDGI^V6L62#=&\R.\1MfMAHPBM3@c8b.EESV?aM\.=b##TQG1baF
I@W>E9gc3b>WUV88)ec^^bb,<fd2.]_6>7gU9f@/a0b#eJVVe[LZ[YE,3)CZK;K1
8>Y7SKO)M)<IFT,;:X<dgE2-XQT<T3,3#RHd7FL.8BX0@KcDa@:;]:9P)FYB:?Ig
?U:;a(QB(<FGGCC89,dN@W/9PTA(?U0[YbeC4&-F_=_KCe?I?1/c\#WeE3NE.M]g
a=D1b9Cde/EA6A:DCQ89C.0T]LTAB2WE&_G[(J^@I1:8CbB&)H/-D-O>Q:DR&_5]
&A[[T:U.\U3&2cI-3g>#9.Q6>PN0]>QI+cCd:6BVH^JbJ2&L]6ZfCb;f@PWG]KKO
gQUL\7:ZU/-&@3.MG&5&(9B2.+F_e5,V6U6fQBRf3#6d4Ba].6(@&;(HFM@P_?4b
+2<F7KC&GL\eH>]4Dg/=Af24(Y9EVSSU19e.IY/dMbBaETD1e+_J0FC\^Bc,-O:+
VVbN3)I8Z1DT@8B@D9V:ODK4X99D6RaY]^HSUB+?_b)FdD_KK^7R1QXadLUHbRR-
^C62]DMc8DDBW76a#?@76WPKD#-&-WKN5.9=cTAW(33IdMG9AFLHfN]<1KBS=W.+
fB9a6II.GEU)+Ue&+ZHe&R)]-&=DUAJg--W_7baP4B>]V6/0WS=DM[P6^9[#<,R^
9WV/c?VTC+\RKBVSX?ZU_[13Re)6Q<0XTK3OF0;d^S-_>[XD_Lg0938)]-Pc96Q5
++-BV[9QN^B,=V^S;.W?=OXK0TQ=@L8g<d?a/d?^I^cD_D(7Z03Zb(ISJGX/114>
:64.@0c(Y(D7f-(S-M7>P#5X2[4dJ@[F&O2CA#UXaX?cf65c7R:7IJ6cVR^ND02E
)=bYO3ES;cX3b&4Bc+BMILT5/.4W\Tg?+YO?KA0(TDHLeJ:;0XTD23[)+WEEBCH[
Z-#-G3<3./M)^g<:f,YLP4,8BY1=8;O_\D8[2FPVRWA-?3dDgc@MSeUP-We=YNE.
@_#E[;XB8\7-4#4G25)1SN(R#fa\Q?JL;9Ag6(?[FcO+J.-E<,aH^AfC+F8MPTL6
/>f;81K<FG6QV\X^24D9>.Q[&aaU,]0TgPLO:L@P.U;g]H,#cZK^-^DX9#16fc>@
7H^.Fc@=3/.3BN3]ZeP,?U6&CLXOg^>>V7/8SY<3fZaf4PJ6B[XOYbc@](?b2]>U
T#CR9HTTc7<C)6dIX_gCE@3TO@F8G3G,X7:IfAgDRO-e^Z.2DDCHQJg,68((3<OV
6@3BeJb+Kf&\X7&G-K53)5^\YL>LX8:C9dg@b+bIBE3VAOEY<J3cNCc9OGFaE6_=
8;SPUTWN1@\[/&R>V]7V@-KO],FG9+MP3J#^&3L8LC#Z.NDac(_Q;0e0CR6Y&[G]
&(4V_6/6b(bPcU&1=3[@70(E,,E.9<.U)4c8<;.[?bHJ=OWI&T:Ie.<dd_.:fI:<
+>RMgDGV\f1ZcQ6EUD+R^=&3X+_:^7ZD.[[Ze?5)?aU)E&>4#(=//;\.T^?FR)KI
@876N-K5ZI@]fO(>c8NDJRY2#E2^g.5K&>-V.\VdICD4&)3H03Q0ZS-g#GPA)dSY
2.b:TPdX.[;E;K\Eg<=H<I)SYN&:KaT,ZC,WCc1c45.\:N<TX@Vf,IGc?eSDc#+_
5M>PP+f3JR6W_W=#3H>f^XL#@V2MVM5fQa\R<+_e/^,<d-53O352e\V69><>bJR6
(V7&P0Vdb6ZDN?NfMZ8=P/LUZ_PND>W(1GWO[<7SF?Cc0-0&A]F\(2Q<T2_+fN79
/2>C4fNH<^LE<6H#6aG;M=W:QP.9#Vf;:KWO,5Fd\?#K1-;RTDRB7IC#c902.fEW
+?5bC]QBM6UM8GAeYc=CR;;WFBg81a_a-12baH[64gVM7eG69^/a-]1V7/-[;6^T
4(Y#C_c4-d+U_GPJQE4KC=UF\Bg(O7H]fSaF)0)_XV3]Z&+<c9>AW324^+&4GgNW
,c#0C^L1JV_NXM4Q3N1QAB?MY\K)7P+UCK@7&a:K<H5)>.cHD0T-U8VILa6ID2IX
W(8&cC_-PVC:WG<-T<68g;(Q<_>d3(<I;FR+DA#)-78?=C0-RaUgR>I@&=#QRb3P
9:85^F;1Zg)N,F(QUKMVB1++6@\R:J/1bKa9VF#ZI.Q2M_Q(J<b60CK1Y_;c)60W
aUf]2BRWfFP,ceJ(1b:3a-53f3PWQ[U87\J4EKK]T+7GT6gR?dHOF1FA]75,FZ?^
NgO-->-9[;^_G=SNS==#&9/9a0--RW76c=;bNVeRR/0)9?RgB2B3/Lg[S[-MgY-L
TGVJ6\#)R#.MGSW6f:c@U:SKDI.Ag-_LL>G\]ODD66#gT\[a6O:PN2^a.:.BK-e7
(+\7>9:>PPY\P:=>^ZK@2ZV=8ZDO2.8Q+:U(,#RK[#3X::f2TK5aBT=+T^?3VD?E
O.TF7-LdeI@C)De.g3GLAR2c<QG?#_X[[CGULOa?M>:?..:MJ1e-Y26c2M<&G/9\
,Gd.0M6?GB&Qd8A>8c0EHgd3UERR6<79.5(QIA]56HU\a:7e,V343(/Zba)AA9D2
38[8V[TU_L1>T?;U_WP##2:^M@;eUVJ?(F[,#ggJS5+AA#:\MR;L3c<Z=g3f]E1L
R)DW>T]SPL>WfM.T-a(P?J@?/NWKS45Y8cS1b^B[[N#X,=N9#ePD<:d6:U:@;PT@
#QfZN_;AbBP2=CaJPOT:6DB2F6/D_G50=>TfM7CLCQ,<<R1#BMf_(YTGMGM/?\c]
4@SN#?F=L2./d)E=Y;fAd0=]6LQF/X_@:4&[Q^WPJ;\7X;;7,47W\++/?5cR_Q&Z
7<MUX&.MgUQgQQ>_GQ)7(IHQS;T5b37/^3bTd+6a9aR[A^fcOdD8(.Z0KF?XA1N8
@E8E5&8BEJV4ZgV>d]Z1BgU@+D&Z\\a25Z(6,H-b)<<SVEXP;=Q;V41D4K21I4]C
2Sc<N\4&GDZTR0#FJV2ga93<M)60GgN/W2eg2N(KYbJ.##GBaCBYUN=5@<SHbJ]D
EL9&a<7\IZL\Wd+B[LEL,2H^7dU8O/-[+E4dTe_B__(3LPaLfH^BNERO.2YD>,G<
f(bgTDO94W.&f5Z@,4<PXO(5GPLZe@YB.3X>LA^E2B)4<F@6U3[G3eD+))9]dZC?
4RY\=CF-JHF:ec8)<d6980\S<f-QRD>QJ)ONHQ@GHX8^2WGeVPP^8SLALGH@b?b\
/6\aF;VE/.Q6@23T3HTRQZRLUKg,Wa4/FP-V@#B=BLa+KZbJJbJ@\bdH7/>.30g)
HF_4\1dCbLZ5J^fAY6[V/W/ZNRF&_2_TMQU#.cKb).7:.B)aK,+a4@WY67W@/V^?
4WMFDdQM0N9>5gV&:\2G)>_?Sb94]C(])/=^Q;7>caHB?YY#)V-3:KbM^?6<#c/S
6Sa3AER,ETP>4a?\-0eLE<NT4WD,=;J,4J\CU-&RNUD.W/De8=QCD;[F<-N/:6>A
L;ZHV-)^XBV-U9@R?09LPC6]\=8_52Q404S,DbQ,_L&B_,&Ia3dOD^^\#DFFJ?7F
;4)dA7O+E+4W51f\O5(S[FE?fVEOWG+a33@O0#=dSY2-#.ZFS<O=G2;<H7;N(S\=
R184Wd9,AC4Ufa##g;NI>9=G#Z4W8L^+@S@3P8J@V;?LD(<bY:1;X^7//V/P)HN3
CAf[;<RR9]OG/T+GL-G^SN#W>8+fNQET,9XQ.ZWYT_PYL(XEDN7WDQZTIe,/.KFd
?6C0A-bcS?0L0d@HaTH:-=ZYB1-1U/+Qg,:G(//C0VUSgc<KPHT5370&Z7;.+4?]
C18BB9V2HYTXU\[GAXIAJeC;_c8U&fCb@:_BP[@f/@Mf5X\&b/_57/:PYF.gLd8^
OX5RAA:W]J6H[\./\0:E<C]:f(P_PX,-(CUA3B.<#O<Q-AAXRddR)[c5D\PIM&J8
AMR6b;]+U/8DOGY?@_V?]R<-E?;4[N+S&,4>&fS);8#4@V9>AH=^12M=&?>3d/82
H_>3MXMdTeZ:>W#V>8Wg,gT5e2bC);WK/TT<Ae8G;><^VJgDOH]02\CeU1dU1R:>
TMLEb;e6GaeKZV1[;9cU0][f>]Q,G,B>74cNe@dgN29:(ZKaeBTV@VA?a-:+XcaK
H]SS^45Z[-EPdQ++#HdH[cXUbMM4,VY]ZQ/WEOTbK,BDg][(M(<\4\dSL>\ZWY#F
4DgF)fD(3EXa8gd.9Y(P#,b:M<MJbd\bCK]@c95a+F4BQ<;&#E;9gI[cgIA#)-<(
HgO)GU6Lc(K,KOeJ&QAWHacV:_TLC;9L0^5:<-R6FYCW)NXJ#\df-<>A6:^_Hg&L
Ve;\7,&9I7+NEO,6>1H+X?D:\:J(PEMJBFNZK8.YM#K;7(;gFW/fK862=G[Y16\8
2G9Wc[^22;L_B;X@O_&T(20^^;#Y)=2R=UW:<>KO<R69_M<_^g@YD03GIA0)gcDF
S&5)S4g89_0+V9IfW/NAF]&(FJSDM#TcT<8.:[.C:Z,TRZ7cX9TKaB.T;[_fbUG,
8gXL;V=NS#Td+.4?-WI24+#M<O;VfSR0CYS?)M/QF?FOB8QTbg+eB^eGEII_1JX,
O53;[VdbB\WFcKT<;HXCR4,AbWDBSEc#K=9,&f3MTc2)K_)O^4S9P5IMEdQ;GP)d
;OC+FP,g2SFR0:8^AAZMb3M\5@Z:fa#L#N2N5&T:B.5/\@H^Z2QJf)CY,Y-fPN>A
aeN9a)LEE];1Z/Zg;&D:1OBWFEbGcHAd8XU&#2?S)f?V:We#E:b22.>9Q.>X:K#0
.=>MHJ939?70aA5BcZT7LMX]T]e&E:9\/1bgP<C4e@,C7&B5[5:PW>T9A(<C_e3M
2-</TcH]U+@S]=\X_E7]PRA<#eFG43:7.9-bI:-3APa30&dA<OD<R]I&_6UPTK:;
&1eG#3,W>K&.MOXA29ZMYg/U;#)CgKY:d]ab@bN1Xb2FC<=69Mg;W#4B0\\ab?/X
3f+JgO/_NXQRU&KSV4_U/9]KMP\-b9XXVb<)&7PdcD3NL2>]b=PK9Q-K=-GL4+-+
)_UI8JXPZ+P?EXH7<?faJ^,7+5LN;a[E)f=1,Wa2=KfC6)^+@++;QB.=dON)?SQ5
<VN3@?#M@\ga&[.>2>&[6517Oe+7J(/QbS_V=-#18Y_<2(DPQU3S?>80(d6DbO\@
?HTE2ED^J3TPM#&,R?J4A5:HXK5e28,bE:/)1_aD8(d3ZDdHUc&DE4@357/X;d1(
,H)Qc426XZKe4FPE.0L<c/9A8eagV.)<9aHU-a;eR6(e>]6A;J#29RQZ=@/KQ-92
B_[(.]M?=ZA,d#2KeZ<eV9d,.AcGXQ@:F)e7[YSM\M#Q#.#A[]5NT6T4O+ZPB))V
61=?^)AT[M:_0U#gQdZefEX)UO1HQVb9c)/VgbT]&aX\e9]W<75BcGXfD33:^H_E
dIeMS^gd-7_EARf@V6[b\16DMOGS-gUZM8bW(HK&+I6ERI58g>GQ3S)(:9>&/6c:
8?WdE@b,9cH=)Oe1^aZTAKV8;LW#V08_UEHQa#WIZ@Z/_[GCL?^SB?d.+.H0Ib2V
FR\:)5e/FR3S],[\;)[YH+4?R[)dK8DEU1N[dbT/46KX840:KgS)WW?H6UOUE0bI
MI8A.Z)(@#=1\H>IIY=#@-6da()P1.,3K1MK(edM6Te^XF?fVML6ZP7T85P72&MY
5VN5XNM[:0c=RA?B5T]AR0^MKXI#(LR+;D?A7a9DSXfQDf2[_4?X,2(4PLV)5[Yf
#[5?Z@2N/(EL80BX1J\#NX#A_U,2A?7&X]cWUS=<97Q#8-BXXdcPY[=UB2\a;+Vf
B8PGV#ZD[&)JeX@O(3SVEH5_^]ZW\7U#eNBV5@2NW19J5U^g=<(fQ&-C-X\d.@?E
-7A1Q)O>OH7)EO]?-F]\\O#AU_OSZ0X>^]6H094M,gXP@Q&[:e&E1]9^SDC#K25=
RN9P=OJ6]@\BPB=/Bd^#(RfcdH(T5Ud]LY-\OfYJ<D1LBNE814W.f4<VccdW@2T\
?RGYfSHEe==_T5bDb<Y(=a3O]Z:;9MJ(=QQ&)=6/<dU.5e7CC\Z>,R@9OZ))H;-+
MINMCMf]VB=.\0D,SJD9JA;(^7fCJ@f0A,cgY+[6AN&Y_,T#KO=@H20JPc<VWU<#
2C[C7)ec^0_eb=94F=(K,^SAAf^XCFd<SCaEYb/J.L)4)3)DO^QBW:c>,/JNKW@e
20@2bHZ)NI>RgBX-#:YR_?QN)>/M^?@TWUU22(<6=G/1,ddRdQW(R?;^aZ&;4eGf
71_WANga#>P\HW,ag@]c0bP1D(d4BG^UgD/b7MO&]ZIS+ddBd/XU-7,1_I[aHR=H
X7)^42dQKZ>GZ#K-8RfT+_:?9PP_:;7KSJC(gBQd&T&C4D2RH5:/=e+<C6FG&e^S
DCeS;9(#&)FLJBad=5NFCE-5>TH/RSJRGBCDbANKTfaXZO/GO(1P]=5bKQM_<WX,
9=g;Z;)WUcT4K6^\;_D/[KK]aAcae=G4Q227GQ@A6DbO\/Uf:aKUODIWXERd?TB4
QH3/78B9>1@)#P-Y-DHW0.,9=PQ?#cAZ-d6\V[(@TEFI_8d#;ZL?[c0^QL4e?WD@
_VY&=45GM(b+Uf1ZeO04eVCH5^bb/2d##[_HND1Ed@g=LI2SDBGDD=KLcX4#O?H0
YOCLH\Xa,Qd(08)CHGF-[cRR(HF&:O,1/43_SAYabW]1OgBAfdDO@VR,;a.aRQd)
bFXNT.N1/0GJZ7a[)LPc(MZ_TQHX-6a;6:349#8,GTTB/E/^Wd,&1C\-WR)_G+.U
M(AS1Y9#_PPT3S]]e-3+YW7La16B1^B44Pb9SE&U0IaN#CgO()8=>2aZ,Q8NbQN-
bV\5929.XMFV+gbg[;baOW2R^OI.aA0XM;I2Rg2MKGEP.CDC.f+B+&B9aK:&g,@9
Z:C0-EB_\?K2/(T:9(\1GVdc[Te@_eNF_DgbBfdABX<F8cUCTX2JB\TH:c+H?2c/
4P_RZ>8W^C:V1FQ/&#(a8a/OSA6a;a,eKaEQ&G+AeA,K@F.>eVYDf:QP\2_XIYK+
@&(6IT<J\[#K,g/[QFZ:RFL#SePW\(J,4,#;[DPV)-C,&,]GQ;0@D=(e8<>e]JY1
F8M<aAbAU7O0J><MXI\+9fF];R1N95/-0O[gOQ.64d3Lc)<0RBCYf:5HQ-9&D:4R
0/(M>(=F>795APXS<-@LKYRL^@&5QW&6,WWY2<<ICMB2.NC\gO],N<4G_EbC14K(
6T@K#&<Y^NW-4&U]L959&:-dZM^5X.FATAD[4[Ff#-d-)Ec.]247-0:cJB)cX8V\
URb[ULcDaE_6;(;JF0_;9]VV5AXG:,64XCf.ULNWSTX-^BdYL9@S,(W?0c=#4<e4
4RDf\CDH[J)gf5LL:T\G14[5=EH)7)gEH2PORY8Ve_A6aAOT1NRgDd7N4M),S-9(
7.-OWXcC^XTEXO(-TX^c>23N&GQ<)7OX\#1E]^PNB0bTgP<V1U5XHQ^?cMJBI<6V
Nea7CJPVfGIMV40Y+2UdAb:;)RUd;]@ae7bBI+1QG))B7d6]@a3>\[GR02C4<&.a
#KB-Ff)H/:0RJ;\eA.U?/DB^O3V3T>.Lg8^7&._J7>cR67,G#(b?L^fgYRCSKQCg
<-J2AX.:I0XX5Y1d(,TC-<f3-,C:E-OC&?;23aIQf>DE2cZaI[1XGCG#a<[D#/)N
U2L:)4(H3I3S2@+)KQHC)SU=,HLTXb,cTD8)-JfaK\8ND-+\c--f@7=X_X^BVf1\
FRJ(4[7:N2?fAGO(+^TBdGc_1[@0X5E?4L;5fM4d+<370JQaB.SLG8C^;dLG@+^B
1=<[9WW_U1P,->FE/eBRU-Y=L?FV).E4Ie=3KDRF;TA/^&C_)\&Z0X-)daDVcb0F
\LI:8QLLI4gIH_a=?D[.Dea4966H(AIGgEZ4Tc/5[>f>&.@/&3fJ&P0GRc-D>?1f
WRKO(@V6\bf==G\5V23F4R-AR)198/dde12b<(bT/B,)VObCX1&GGQD@[N^(9<M\
\49\gK^[^:B&^[)E?G6C/?/gJfM^6Y(]_1E:@SU#SWAS@_@L;JF?>.6]R?O/=@,;
[He6b=01B5XD&Z=++a/.)E=&-51?=c;WK@a7W4Ta=@V.9???QF&^@3>fO\E86dM5
G1.X..XMeO=><Q/9^=^>&98FfR9WFBY]:VffZE/,MA-QgLHDCN_TI-d\_Ad>WS-O
UCUYW,K53]DTfFfV;#7>S]KbQ=LBgB-[].JL?:\@d:eCB7/@)2-V2>QC1MN=1fIZ
48dIVXRMY)2Q2\,Fd>SBZG[\T^)C29--:AMW1bea6.OgI7A0R6E?4P],W=V\A/g@
A^P69L>]MT&G0Mf.\9F6V_/I:g27Mg\dI0X+YRbFWUCE9>IEOPB9:9;P9-#5#Aa:
2W4SJe6MS@,,-gQXd6]0Qb1[Z-Y+=#g02/BFMfGVPGYf_=.abX[]a/S.Y+D(Pb]\
EH;TT1C?(N.DHEe3#\DJNUgX^5Q.FYa,.8Oe7b9AAXYEO;2:eR<]RA_@YOXW?6eB
66,3JS)&.FS(O2)76(]S;7V>9DB)_Xe7+Q+c)=e^2G)eZYRDM,eXJ\^6;(.CG5[G
BfP,E/\:/aSbFJcT1^&#+C=(/]Vg)50Nf0YC@))V_@N82X4gB^VIXW6IZ&QI#)QV
+Cb@@&?CE(\H;0>O4NgE?Vf)ZE3Ja&)U5_L8Sg.#[[F5\O#HF1CcU@0Eg[Y[f]aK
XdEfM=WBEI3,R-KPE9(UDXVb9BQP^JFC#V9#]?e8244;>+Wa3f[CZ_BCg99?W+DP
]@>F=_G,^GIdDYc@3,XWO\1.&G87Q(H&IL9\bgSOd#TWSRJ_([?R1287>g<-PV@H
b9&Mc@0A2BEf)16-<2H+;[,Y+E6_H:-e5MZ^RT/2THB(+71))]@a.<@_O3O,a#cV
ZIA/W;LJR:,Q9I=)bd>g00K9C#b4+g=P<[PTG\/b@D>>=9RTPgWBAccMPD.V9X&_
_<CW+\PE54CdSQA#CMN[^D5Z6G^<6;Ee/#;#>#?CAK,^/.3?^aI1bHK=63(6ERMd
MFLVJFf;_2D@1^a]DN5&V,)QLIa3c1J&-A#ZdAD;JM\7c?O0CR>^2^b)I&S57;RN
7NS822KR9/:WOVgS4M2R/:M+LCE#EH?=Pf@=IYA)FX=CM4S@>3:NDa;K/=;\ST<P
&9IbQ/=8G6&RFQ@(WCg+ECgZ<fEJOPJfD1\F8)]9gB7NI.&\R1A/Xb(.Nb?W>^/=
1VR^:?/NAFY/3IDAU&F/W:>g]a:2cF\?/2T9#V;X=f?MA0/eJA88VP@?3\,Hg5[2
9ALAg>fRA+0Uc<64]D&=X(EQRMX^52,gB#K,UJGU,e3bgV&R8VO,_31H>Rf-M++N
OX=.,/-C+N>ObO?H0B-@BE^\OSBI/)(O1^YB&.X@XV/A]8^^PCU<XUJO6,)O9IU(
)+5([;;2:D07+RC0GGgSM6#Vc^/.@0E.3QATc@g+V6P3.\K/(>a&2H#EH@HW8UQa
Jd-RPJP\Md7PbD+>R-JRB0=g>#[UVfV8]N8d9X_G.]TM?9-<<J2g7,PM/RDUA7TY
&Ke=U[B0b:fQ?R.dVf=beA;K<TY33:W13#1ZCZ,cFEdDH7N7U.3)A1:Y8aeDW^(7
<GMA-Igd?PX]EC8.A;5#(.AA1;4BDIO^DAJ27U<c:gK:A.3UVVF;UH45>5Yd9-BH
GT/A\a9N;5c(??2<?^e7CJC01P1E[-^P0M1XG9.=GT2(6^7)]_eYL0e?5FVZ.#H2
:Z=IEV^I3g<b>Y+dOUdSe\[L>T+W8c0,RPYU/-K:=[R\,ZZe<8e7&,#8#\PEQB68
B;LKX;=/dF^GHd&eR6L\UXA);BB#IM08gFa9JeC7+S->c(XT>N#@L(S<X?B)EL2b
T5(C)S<54DEf@V/4HfRJf8X3E>VEaK,X0^Z:NFOdUXJ-KFV5&/\g^+S,S_X0d4fQ
ed/MG^7.,UML@IaCQXT<>UXcL3HB)4B57-H=#3C>E\[<-5UZ\?>#c[GS-UeN9AS&
;X=A&S)MPV+65Iaa-\NS<f<H_X==_ae^23#d#g:XS65=+7XV4TGAc^7E25<PMf(E
cV?.ZCf)XQf?f\YQK1J#,X.+Ic55^YJ[RVd,d6a]4c1+c[YAb,7?4IUVXZT)9C]J
RO<_S=_RW-#GH#C0_5>NOP.M9a[UgA,60<O@<0f&4.63O9N0>2>,+Lc0E[,H4OA@
_-1\^(_BaGB=-[?):>W[b4Sd@6O2bC4OWH[T[6O7KU?3UD5M&PP=B8UNT/8.[WMf
&ZK38U2HC)H9PU9^(Ha_C5H/@X5eICR8NN#IFIG6#ENI9P5;FVCc&eBO9M9T/2,Y
>S<c8I78OI:JdXK\05G6,7Me\HaOU&@OXIa>6L^UOScLg-;.g\YS@Y:.bFM_gVdM
OOKca=Gdd^aTOgECLe;&e(cBa?38e7bfCRdDWT9=aR7L+.+_Z6gBUE-8#<,OKLbc
bAc,TH&_]Y,F&[cI:Xa@T\cWA+@/GbZZO2I2K6::O@;ebNHf\XgE9:@Q:=Y;^;^V
47063P^RE<OS4bH6YJW],A+QAT>__./@9SEU8e?:+CbL\+=@6g55#]G[.6=<.;b5
O/-M_geNNM7QK@]0APH-X7Y7&8SQR>fGg[,Yd9g>#+4[]S9AG)S?d?FgJ?.5[eL>
7Id,;IS+BGc3Z_LXYYY27SP]/&f0&Nc@@YZ7TZZa)_R8d6N\D1T[)19WH^TSUVda
ILgI#g:eWR)^POb;PB=:UW/S_0dMCb+Vg-9<CLPa[PaZJ.)[>=EF1>[aVQ?:8U0O
-#,-98cSB4/PR(V]6:95GfGJb^cP&#]2V73=Y;K/d4PIN?:O1[6Q(<[JR6H,dHO^
GV)Z13I:N+&4PeIa;T^\?LROKaeKMeg3.OTA\EY/LQ1&-CCWM1O(K>-=#)8W_DDY
F):Sc:3O6Q;58IB#G(U]&L+MPR_2DL[MQ^(_,@H5:.8SgER9FC1@1&U:)gbQJ>d]
N]9<#[?)&cNR00-:d)R7b1EF+f?Zc8H@9^NK&)V:]8Gb@7=(Z9PGL>Q:1F^8BP>S
bG9-=>N)^MXSacg&E&>5FV,I;/a^X>dJ#8,^,Qc&>8+APHN(65=P()=,].:E/X8^
bY<9H7+Q3H^<dUDPCF_Bd9/>28bL.&6H9<=W]e=,O9Ld1]/E&2WXH>ag).@_<a3B
AQZDDW[B,V_(Ig]_-NdG2bMad(O)&]VNCYe62^P3[T:[2/EK=gV6QETOM85G]AFK
96EdX#I#U<#GX)Mf3g259Y8HP:PD0Og/JJM7/SFO+f3OPM<#\U+SZ,AB2K.W(PH6
:9;C@9P1c28YU8M[5#BU1OF.M]3<XS7EF@U[W1Y\O\g\(&Xa4UBJ7@:0DW?PXLSJ
G1ZHJ//2FT/Lbfd([VTSJ;IYXI\UbI&g>+b9MK;G]7V4D8GU1:OGWRgT+KJ\+MDb
K71IQL>O:&:&PV(0JbQRKO,D@IJ^S1VKF=6e#0?CaV^b&W6G=/H5J;9YD&I,a>7Z
TXX6J.>&6<@+WOINB.S^]=e8O?/X@2?0=0XKABf,HaZEL2U]8LCG?71W)3;I:Q+X
SZ=?S]aDTZcD]@^AV8GZ(SM9ag[L1Aa;MaGV9WKNfBCB^L(0BAG2]6F?W-2RZ:\2
T7FX^EZ(//HgIQ97gSQ8B8#d;41BC2[>I.3]d][89&D.ARgZQL&,d#P=(Ue?UX]a
.+Je_,)6KPEM+b/:f/__b(23ZJGZbIC]d2_dJ6gJF1.]&]CERf:=G\GQ4]P2J(@[
CYYPV#:?#-PF(O>/BF-fgNdg?eEF.AH[N7<)[Nd,\43E];2-CY/97OO>SH<<PHPI
OVJTQGT90b((<ZFZLXU]#?(/[30a#b91W<89cXaXVO?[B6<J[LQG#IJ77KNH5X)?
EBH^Q503(&JDGX)#OLg=T1T8)NQE+,;:e_#B^3&(DLA^CBBH/eMVT??-d:(76VN1
HUB9&--&</0BR@R\F)d#M)cS[e7;Y<Lag5CC33M)b52JUE).<AGOAA/[K,FR,)a5
6Q==PH@7XOL2ZFfOd/dQ-E7b@]S)+@=WI1<@9Zg>67U-GTQJ@-f,U&Q;gI4>d7/P
a]GL6=TEW<A5OU)H6BYRbNC<M1(43QV9;>J6d+C2E#M@P0Z(2X\=SeQQeAN-FR04
49:4_F6IPC55B._C>V2TTe#2Z)bBAdDOCL3E[.8\K#F=<C;EJN;@4J-V_-)([)OY
<V,G7V[b,VHg5Cd0U/L#^##C4fGDSV#^1fU7[D(,W^+8H-OX(:^8&\YZBNX<>6_?
fMO<VcW-3;<J]V4N,;Ve;D3Ec]4(-eWcM]O053@R/+6\8eK=DYFX2/AC@8L22#TQ
DEKH;#H3gEZDf;5^d1#b1T#^)4E=gJ>cY(S2&S&]FHf.cGRLNW.)?Z-Y]N.eI/bf
KRIL8G9c+I9&LB?-a4XATJP_AT2[:2]bHgUM=,ZPPVI;fP8J:Jg@2]=O1^Bb#S2>
I6GHR0>EJK0Wf.[+Yb^MTFB4KaFL5e-0;O.I3JFA/,)@HWT.:T>6-BUX;b2d5LG\
^F.OH<^T@+679C5?JV9.We]?Ye=,?#N1KdUH8N<Kcg1ec:&dJWR8#\OB2N^5A?-G
fS(#GJ(-f+fC^@TP\76bLb+b\S+97&Q3F@3>f]>fVb]&+?&D^O13<?R,.g4;#;R7
MaW=CgK<//].QK];G:P)#(HS1.],<MMa.X.f.KJcT&/g-K8^8ELd3T#PGabATcaF
E5IBAMP+_I1eY0U?4[Y+RP4>966IE\]CL=W_JceCYOTc)XL&8<([&CKCJ;\fa4&f
ePF&8++&>B@23.FFDDK1dXAX^WC]5e:4[OCSK.WR;@[N+fC)C^^=@e/>K\/B=9\X
MY]D6e0Y8[O7>TZ,7Y,7=_[eK+7]HF=0KdBOf>3U0&U8M,HRVF8EPQFN22)ZA1D#
3:\1.MU9AEO>3LBL7FWQS/#WKCV)/\)J>>NS;F6\TeGKebF_5X:JLX&GE);4>aXO
>>[S3(QSM1fO7M35/GdA&#0D.1g;T@e,L\=J7[;aP/b@B>EU+3@S6g)(_R.M1HT#
gf8U1[VV/g4CA)?3+)T8_@4C4;3FfN1LFJ4bbMUK7B.5??f+T4LW#Bb1RU#\d>FE
)ba#N2B/AJLf;YD5[PT2C=]D/63G,\HPOY7bVXb&Q4CTY.5YLQ<E7FIUKeR29#MQ
VSaPN^^(F#A=?\GS\,:A#dI;#JB34eD2)6(Y3E<PL(Xf3efH+HDOVL4<e0&N.8_a
L9,J)\7_F)TWNc.NPGP40V2_#475#XbZ[G@Q98N@a=,.;9P0Z3TUK[:=aQ?L)/E6
f_fUe\(#K).8/A6<GY9481G@gC^6^&N;Z]VKeOKF90^[U5EX@IG\SPCgM1Z?b0/1
IR<BH0#MP4T1Z]751;)HVA.c+\=W>25]OD84aGKfQ1JR8/Ebc/=CUN9<IdT)Xd1H
XY9;a2]f3ZBg.aANV7a2Ya&?\)\MGaF\.I=6#g^:dK&KaU^.)7]<KJC?Q1K9WcQ5
Cg]\P259(EZ+N35:U(@NDO^=XS,7acS[?N[&>^GfIN36Z(2G/Ae(G484a3.CgL/b
IR<R8WLfe_=V;c/X?NWZR?Gg#,29bG?PKg>?S>(3N[MC88,L\7M.8Q>N2&;((H+g
0a3LDE=-aAE1-#,5)dS1W2b>M6VR./I;D&,]TWefN]0#DBNY/=1-K\/X&QJ4b95X
-13:<AQ\IR/MbB-.bCUN0Ye_NHQX<+##1HO._Bd?HRbB/]E]CTeDa]BL-R1)P?;9
OHRVPfVR86-;Yc>X@)X\(@P(Nc\NC^<E>WKT3Aa?&41-7cH>N;\_DWIS_b?5F5Q4
5Y23P#1\dNc5C(Q]>f:KG)\/b/J<3^+=JH^-+?C^MF.A#ZH9V_;L2_GDfF_d1CBN
G3(1#UHbG64<#YA8J>&eMR7UfU2V+Y69US=QcCTGI=EU00^:-9TY>be3GJ/\DTdY
RQBVYcR:=+NY\-&7GB7Y>F=#WbSe1^(([F\GDeA:C#/I)(XXF5YgH4GMU52CNf^Y
IMKQ<>d3F<(a1Bg#VF]\CZe1[_02O4VbR8G.?G\-72/cV2ddgT@Ub(<PbN]:6LE@
.bU^RDY#Ja(=d+JfX0KHbE_0ZbgZ0\TUW/T3FW8)^E<6V0C[I1eJa:X](LY]U;b5
Ua<e/?8<1f.Z4/Y8UV#D8@6Q\U;^:S00BO#00)<W84bZU.(+-Oa:\4@:X_CK2UP4
O1;P\E2\)G5^:,/C4C78;WfcDK/5Y^ZJ+6G<+D3_bHWL)5OFRMHU20I:275(Re@Y
3,.DWQdY-)]=AS[H++?;#6GE3]A?C?TbbBBB\&K3=]X,0,]V\6K+T?=6JZOV[XP3
-J3)^^VB.ZYJ-aRO-\U\.>W)>+T:/=HZ3(TS7>?aR3A&d8^dbd@1OLTQH1FQU:QC
+.O/0CMg^)fJ()FTTcDZGL]2//)?3S4WbKFfH>]N-KJJ,US&##S5ONHRd-7\G2AH
[UcFS=,8JAG2>CK:CRAg1=&WN:<CV-4]5J<9Q+:/+:d\fQ\M^@f4MCb@IWAeKUFE
7-b_N:&@f#N,L0\L^>FWM0]03CECK1SY(,_9e6,>[ZW+K7W\I@RgX&X@1W_^OX7P
O#XWV??R,?8GUU[](W4g-+YUObE1G9H[R3G;+5:N-,UI&P.Z4/:GF<TM,>#Q9J@4
FKQ@G(Y.ed5@Bb-<I;XaL#)/.V6KR2G?@@OZQO7_U>]_W3gR#6,KfGOC7O(d(D[2
:,)?IA45^UT+334a<e@C7J\)A6^::CM3O4VQSH+B&^0O(MFF8^b11<6UY8RR?3D:
ZGH/E(Zd4eZ.5N]d;_9[^VTM35)\ga+)BeQT2VX.dcD--^\UZ7F,\_O,;NU]=b(T
?B^/:6XHZ\.VB>USQMCFbGNV>5f(X&?5&YIL(Z1=V:\E>&]B?2.d1WUHGIF[[E&(
R+OXZ4g)9f;Mg9^Z3/DKM]#FbC#:#EF_.bV&5-(OELZ.0^J/+@GY^QWZM0@QOW4[
W4@7^;]ZFUCcL;VFE3b_#\315XVB)Y5C+dHbPf.L[MXTV_7M4bHOC:LgODIf@@1;
/51GI8P#:>FPVS1JY(-(QFYQ#\AbPT/3ATbH0K.L2D_]fTU53G/[c-2,E;,))0VR
#P_0b:+7?g\Ha4X_>AYRC5_K(L\9@@NUJ8,B=:970bB)85VCa6K,C0.-@AAPe)(V
2eJgV4P5SZ=O24QGODYQEA/5,GXF<YSfF7SVb]U^7BHaZ\]c@;@J,EJ2VJMAa2ZI
9UHXH(6f/EZM9-SO6)T=OR@6^cP.GM&P8I-/(6SUF=&<3XbHTRJSJ^B)48LUf&Df
^Y?AU@Za\PBEZZW2KODNHNLgUY._.I)fZ?YSM2U@N5??>)V52-?WfB/-Ad.&GUK#
CQ#KND0N?0\S=7^DFV(;I;22H:2?V<L.WdE\A)E3=g&DY>?AZ2;GURF)e7K1a7gJ
PD#2211-LaFSI8BUY30#RP=HTT46^fB##g@=2&gN5\J9V7fMUO;M5a7^CC@Q-MVJ
#-bKB(>TKg1bfVa?KVdUQ19deMf?YO-]794:\.;Zbc-.Y37UZ72P)9-NMY3HC^\+
V,@IJD_GXIZ.RBgd_/]\I/XQNN(8U.W.IdCf9Qb5YQJ[UNg]\5S0D<2,P;I>]+XL
YeBQNQCf?42XTM/MT?a8ET:1g:Eb923=#,J>7O/OX5U_f?R1E,LaZ4[RKC7WVW-g
Y>5F2]Re(6eJ-]C_XO.FT/L52g_)IYc?)P_Bg_X+K>7OA2B<0GJK]9L0b^_a4J;.
3LK(9D>D#ROD)>fDCPT<EcZL,CFH]+;5SIM#/.CYK+GeZ4B8/\12,KC(_P#a1]9P
MV=9d[:g]QZEF/Q1gGJ=K(,__DTGSKNB1)^QXUE5D[g>5=Bf0.Ee(SFS]9aXbe\G
fL<d:M(O,E_1(Me37NWT0^0FQ[2OH8X(8OR&g8g:EE\WA8>,.e=M.1O_N+c.eaVK
5M)ZK:3aCb@++3T86MQCaG;(aE>0XLMg@Z94S:^O&a?Z&.G/5XR]/C/5VdGN2(aK
>8dM98_Xf\XVO<)RGLg2EI^&LdO\7-6METagH^1Og=)3[-U2b:C0(AC9PcHBQ)GR
P.egT(D(fd<LA/ZS@AY7/W#b-@ZLN(01#J>UQ3;8PC<0#:O:>[AaN:IcOEDR23DK
QA==G)2]6D45[HObg02]fE5eS7[f9P(PY13[6ESZU3&:J8;7&bNT0@-K0CSSR6bH
+#ReKEOaaR@UaDL(Qa@ObM3ec&HEVYUa&dH.aK6TC<LPMAO2&3B],+aX/_P?VC=+
2QV=b4f:c=>cR9+.\dDc6P#SbO8OJ4[JegEHY68e63=)3J2BIXPZ=5KdF[Z0EU33
O[.E6]fSNP@fB\&>5MfD-UWEJ;ZIEJ/A\+20c]GPWY8D\W79+bQM4LHDdWMO?=W>
SVac4UD>fAU9fN7g0>&.A0bHDR:=a\AHYD++:OU]KL780IEg+/\RE)fJ_]U/;[fa
/Z.&VE[X-b:cRU<8:ZF[RF0##FG&7YbY_N);Y&T8PZ7f[LXb+1eE@1@)1Vd<SMHH
U.@E1AYe9@-K.A4@S-9(IODW(JMOZDK;^<GLdMe3CePDJ;RGM+8e.#B(Y+fWFc1)
d+<AR14cZEE<B-6Q9&NA+abJ+Qc?aGX-T961WDf7>5?-;0-&6=DSVWL=L:EFCZ8?
[>d+]JbP(S-Z2g(U[[fZ9):?b,(.#/S?..f,YHW:JX9V+a0II3eX;QV5R6=@I3Zg
<6T);1/V/,Q]1,8Z-W72bSI._4[EN]FP+c\>gC=XaPX^R5-^\NY9/6(Y=\/dIK\P
KA8cU04>Q4)WQE67eK,g2]G8Dc&-8fg0JH?EAJIEcWRS2a<AVH:+ALKIe3LaWD#Y
N<_,N&P#IMLDcQH0FU8)7-MWI-L/M,11E(ATa.c6Q/[YV2+]NJG-UZEdX1BXfE6M
gUb[WK94(VVMFZ4H2AWJT@;80fTXY17K?PSd[[GJeFI4f^(<FIF;O#4]R]EVMFYe
1:cG[cO,GM:=-[gPS:ZP7gVYY3U/,+-^Y=4LNe73.1L4YVd>MP3B@\HfY52EG9TQ
A1A9Fc:N#-6YTU/WR,9D(5JMe/CB:9C39.,W/ZLceL0IcP,Kc@g]?MUOA=+W45LE
7=^>?DZ_=A4\T:ZK0T4TO]>ZbOMEf>BEWE]^#1+()[7DQ7-+6cfE/@--VBP\>4(<
->IeV&EA=^RPbZRbV:cfTIW\)26^3B--;ZX]I7CMJ7^(IQV[F<2>.RWE/c.-4a]K
aa\W2<bW@3P\eA+/;=?Fe;90KF=[<bT:Q_>P39<L7BRG)S/G5:U=Q2DK]15bM]>c
[N)EQI4@AEUOUA3ReP#:Zg3PD&HMD,7WMKK+&S[A;LY:Wf2K9#DV=[566B&G]UDA
EBK;\A?e1+f)]/4LNW,):)#TPKDMDe<SZS(HK9E2?\a<2dNKX6X_DXFUT_K#BR^T
#W5T.aJ5N9d1>L=MAJE.]HQ9?VIQU<SC>U0:;8]78.Z)d4Z,G?gXZYGQ0)C]^<2G
?c&CV:,9(^7,1QYa3SF+,9RF3S,\.>[,J)23A(aDdK#@R),2>2f1D6<LT=H-fM@]
10//E0YN)W[e;5@,=C/(C9+eQYKG/Q,KF&a)JZF+V66@3DW5MC;Zfc=IQUNXB#(M
[W=#@W[@_S:2D;1&.Z=.<;fU:-LAT\Fc[g@.6>U-KE:UF\cWEU:S0H^M@X4K[21D
CQQ^\]4)a]g2:gd5&CMZWJ7A9E>&Ke#d4b8.J3>bc5bcS=NKMIg7#@JG,JEP3R9)
B@-W1^<aI)K,V50@@ZV(=EU\aF#D_=EACD#[I8;(ga:)/LSHNTM8/3f=P34Tfg[S
#B97Tc<7@Z<E6BZAYV>e>df,@b_e3RQRX]P;=8b1:B>7<66e;PM,QSGa+[^/c(7.
gYS6f@9Y>eNFEeQEC_UMDB[I>GX7@)M1bfG1M6#,=RJXDO0]Y.7]33A)gC(g0K+W
2<([Xe\<4G;0AYT[I43^J;&eTBFQEc/KEe4#>62;a&[CL6eM+,NY10M6bNCBf/AZ
^SN/EeOU+V0S<Y2TL_V=W3X:g0C5:/VWd<)2[G>(/FQa[4_H6I1ag:GKG[\[2@AQ
aK;&:V_^I.dE<Q5T1D,1e_@bNU/^A/d>K8GW:,)5c)RdS-dH\L._W5KbK;HbC]38
5@)Y5ZSB69,?=d(<3=V4d7U5-f-gK,-D[4/;SV;JX>.?H+ZP,U?6VSUM1\KU:UB#
&YCc@+:@NaFJ\2VWR2A7He;8MIVHJ)5T=e,Sf:Y9(4I,KH/E\1KeTN4,X[9:Y78B
LIS)Q90+6-8&4>(IWPUE3<2WUH\()Na\0aEI+K?(TN(\^E_2abP(PB=;^_Ob:\MR
\<\0#6,_ZRe<LVZaa@Pc9(2R8=_SJ3=\EcS<IO>EC=9c_+IJ2\B<g,683YZ&OAI/
DY)JQRI7&@SPBbTQO/^9(:9TIGYUgNgPTT9=&)U0L^?UKAXb^]0VH(6G\#YH9[Cd
gg=P=&P-AG[]?Y;B0M46C.Y;XQ((b5UB#cRNQ&Z:SP>?bT[@-S7=)PNPf;)KFUKC
-)\2fSDf4TX[3K8Qc+V[JaN2bF\2M-26:c]ANb9>->WP7>0>^JPMPae[QN9JDJE5
>TGIH=BKL\F.]Z@P-VA(]=gU^Y^0,d^GH(LS;\+<Z@-aF(L6;1RdL@UIGA5.I7M]
f0(?F(a(F]@PZMD8(R[a.U<5&\><80aRH.VGAaeVPRf\,V(6<;04^aGcfC66(N.a
KU5A,#)7WJg.]JP_X8W+6g[BMV&HA^f6e)S9@:-1^a+bJLL39)G/e^BR)Q#A3V,\
X>O_03)3\HeD\-;RNDAaX[6Z[V6f6+f>]=@Y9JTCeEaV05.b/JH..:eO3#/8f[N?
YHUV)XN[I39c^(-SF=7IL)F@&LL,c925T)D8HSg-L.aS=JT\K69cb>1)2\R?:E,e
.c,/,;._XVQB/LO=;KG9LY^Z?00QddM2>BW)KA.fdT7NE&QEbJH\JT/gWV(S3ecJ
;GXR+W^SMQX<KOX0>PW>^cFeVX==Bf?GJJA-^6#O1_PM^=[XN7NOXB/=>&0W^5S+
N/3-V=dW4AGe2:/b(QL0K@Ie<U1F,>#aBf<P,&)GfJd@=3(48eEg-)Vc7W:#2C9,
@/XCZ;e7\7bSE.-U#fF41Q1H)7-55&4g@E:Q/&H9Pa27RBK@1K3:H.\NN1d-<0NR
==A)[=+EM,&-96YGE3fV,RW>RB<KK&A4/_B^eL>ffeF<.F)PXP>]f_Y(<(P;6#fW
7SLX2N1)YS+[cE-_dJZ6=+9GgOVYE2^2INXHfK3<)ZKRN.E4O5G;(;DAWYO#,?(V
0)&;S5a82A_NF5?IO&D6cB.WB^H=1-WERJACM&\50/AT\Ka^=O,_(EgK-.[WSd2:
eGJb(P#^D3UC9PGV?ePR]X0H1B?;OCHN12F^A0Db5_Xd7FI:,R.>KHe4[eD6,+IF
b?E;CCafBa]/OIb#E^:G^dPXHN<4H6X\e8-g7Qd&NI4GNR&PL9Re3cd4&+Ec\gF@
BVU5a^/A(U;3+X:c>J.N/4WfAV1Oa;G/@=1)Z(8AEWNS1CFg7>&IAIS3cC6/I60O
CE&4\DVC:^8.(Sa_2eDGb-:fPNP>6C6fM@g<VKaOAaL;GUR7VQST1V-NNe4Gd_R^
4eZ5cdKcgK&HB-AS1_@(HP76SR2N@EWf>agPCCJM[,X;(9A6NNY00_YVJF8)ZfP0
L[G,G\2<b/2#1OLaA,#494XaO66N5W3]b),7dJGFQ2O<+SC&I1YCdY].QR484A)/
R_cC;#dI1g#(#aFIA+X25A#SUBc2cK<c_K)L4A&)e6O4EK=7a()Ef-,2^F\ffA3H
fa3[bMBSUS#MX<6B>CX?a)]TTb[PB,=\ZHW[VL+2\@4]Aagd.8#U<I7J\>;83S.P
:DNH99UMJcf1gMa0WWP>6b9BgS2HB58=(RMJ.6#bR4+;ZEJ1N([>1U\9U0gE88+0
#&<T\BYHPFbLLf:c&LXQRD:CA>]eJ=UNXY,1RU1/\d0GOCG1UC/?L[6HK@d,CL#3
B66\>:;Ld<[7#+UMP3>BM9&/2N>9ILKeCX_a_3dP(TLCMJa/Q2cDW@X=(>GF>cdF
g,7=gXF.HYL9J(DGFB73@d;a5[<(:/[C8+Gd]&H;?LKI2];OUPM)2PI)0F2UOBa/
-4NV0XT:@b7[PQ]WJd-:]YDYP-L=4U&7J+)I15<MI1&#29<16MGOU1X9g)3_QcXP
Pb(L2;C554WTA,-F><HT^9g-XNDAQaVgdP2X:M^:W?M&NGgZ-/(5:(7:_WYc0WWL
2R@.U7OeRB\a/b@ZZc\WcCU6FZ68FeR3M&>/L&J_gcC^dM4<P7T)75VZ]c->+/4-
Rb_aJ?;\KW1CB7Pg)d^QL-0N7,B)U<\THbPM5K9I-+37A61[GWQ;6]5CVg:DE#a[
dD;+cPY(-H#.-8-8,Q4M_6c:a^P;+4GNC7CACYLMdBfGXR9KS6:T]6E&OI<dJ?L/
6[[J)a5PJIP@bS>#><JW];[fF_^c1eTLY[\W\54^>dC0O3?aAB&X]BWRJ1DQ)B63
?(c1?VLac]L[>0;YC-2\L8\g&,Z20]0[5MC>Sb.&?;\015eS<)0Gg=A4-WEDSKWf
O@gDVa[<.SDOR@Ff9Ra>S(.;c,N,Wc&1#:\1BRCA]?eQ8F.1_>6066/.:2(d<#2I
:P>5N<UKM27fE&FWM@^&U)a;EX(&7WGA_KS_6=NHOZ9/083>bY>F,J?(Z4+9B^4O
cY-@/ac4-e^V\R:B2SAM-VEMN^g4UYAQ[Rd[;R;bK[YLRX76=e7cVSD2G4Ga+7fI
K<7Y>QH3Q:CGe;<;B.?APTa:-U5=d#08<;b4#<BXda<e;,)f6DHggZ)?VTGfeIP1
.-gc@MUTCU4)bSa9Ga5RU;]8OI1:\Hfb^a:fS+KJ^FDE-?,@]ffGJ-dF>BG8b+8(
+c<<C9N=SdK[36GO/&g_R)_X312SEPX@P(UE63A&2PU6SN12JdHLJ@ZL@d?3(L,Q
86.LU2#a?Z.Qe8H/R<(c=^Hc2^E1f#<R51,QC)<4Z#SWLOZX99_0Iaa6=/RdL2fL
E#_^BWF;-cCaMUR/72;W/E?ND_X221Je3<<-<4:,[IQSYJOO]1167_31]IE\]046
K:HG3,YM</O&7)F&?B2(+&CZX0./_,&U\)^c#DPUV]&.IWN(;<2Mg7aeVcRV.8dI
Z(&>(ED7I9^FA-Z(Qa2QS#B1<,c62>FK2Xg^.1cS&>V<^Wg:/F/bP(SS[-5T51N-
9[4=F0:FL#X]cT\SI=/GWN5A]dPMd7B_7dd&#dcBcef?R6YCP98N;+I-5AX<T.aD
DWSJS[-,Y5+#6S^4C8XGcI]ZY/<FDa(6N,5aS-fC(Hf9gG@?>CF25&4\AeHf@A@W
F&2+K5[^YS>dF3_/-6(?<<&@;I_BKg#-aGAR3Z61P\#12<S2d0NHARAZQRD_\#Mb
&b7H&OA?75W1?a,-@PJ9D.LL3CQ@S8c#e7W+M5B1XW;LO99?:N>f6@9RZcQfQAC\
g>f#_LFJ_Fg4AX,Y,0/C1+Lc=EYRQ_eXDc:-M6+BA(e/]5d8gaOTX&=@.DXUXU9@
Le.>P8]J[-WT,P,.g^c[Z+#)gHRU,L,G:[UZ&aed:Qf++PN&:6E;Q8Z7#OK+D1N-
eVfYTQUDSdJTIJOc+5Ne(39+_TZ4RC<#I:J3NdNNZ_dE@GCVbOKSI<64&A;S[Rgf
;BMe?G6N\KN1_@g:2b;g@@^:Qe/bP:H1YJFS^]&@/L;9DE3K:>Y21c[F^SY;.^)I
VTZb+7f?<+B)9Q0]#PL<X(=&-,fQAC+X62Af\-_dOEg3WHTM54292XC):1_^b>WM
=Y+TOOdQ0C(cTT1^@@bf/b#[YEG<[g70#TL^WFIaf=a6B4cb?=JSRZU7HF0QJ2C[
7ZfT,3?9ME+]@eZ[)bU>;CY6?KA\FR\)&[[L1g_Pg61NMQJ0.52A96;1\>-5,WDE
eUQ=4\J=SKfWg7Q@:74US.5^(]9I07:C92>4HGI9IfDT1_I30c^@bMR2:N[RUQ/8
f-3YB.<Y:7b0BB<X@bF/9DD#0(P11X9Y05c#R.=E60.3D:Y^-3E]a6fJZ1/Ye/:d
.UHOUD8R3T7>,#,ATN&-9UaJ>_9/C5_Kb[:+&>3&XGZ@.2M4RM>?0[+CQ1AR/V6P
]<1\&e2@eU8W5EK:9=M_<&OXeHL5?:;/8EK.FUIEE^8]?QD&7=SFSC[CWaH1J=LE
4(KAPOO[cD/D=ML^O.XLJ6F+YXSLGRb92U_;R-RX=JPKF1-P_W<09Mg4#gT--)c-
1-B0FM;\L&[PO/+dH2W[)TI#TE/TM+VGAbRMF^I9IOXZ\F#Y]QBO)D?;2/)[VT9?
Q:H.bBK).^IQQM5SQd,XMC(e4#[]ZVO1gU@U3e_)aDeZ#D6]J1.XQ)Z2YaVEcHH\
,T-^=8(.?W2Qe:])fe<?LBc?9^BM1=RQ(RTR>OO.;/eJ(@_cV[O++d?IZ>H#]^Y_
I+_KF.F.D]FEGKG[Y1((Qe8>>.VKP47I.9__F;5g;H@1,&(?/GO;NP6IHX?XX?0Y
I?e8/9X8K.B,:-gQC_Ja)d7^+SS[85[[GE3C>EC@,D?.MGF+XIZ_3DM4=9^2:)L^
Ld72)#0H7V1?\+g=AVQ^a&JLAb=E,f8Q?L99:SURI.A(61dHND.\f<K<=Xfg,>;:
2GXLNAPe,21QX.a8).+IT]efIb.)P6;Fc^c_Z5KDJW@HEK(9-C[_DGd(9dG/48B_
^SQDD60aO&WDEP8R..^,]X>1H^1,]:\DP1+W7cHMVEHE9G/9]7P=c&U8-C&KebXV
@e4bNV,4ES:7.agG2,^]NcI:34G_HHBMNU54,&]<Ee0X1,fJ[dY#6I+O@,0M-QZJ
RR03:/2gD()<-CUHcUJ[E)YdWcIQ4&X&,+#V+gFDRMZGYAVc4-SaEf#ME1g#([;?
Ue\Ie<RL\#+=F;fP-IdQKO@J_XHGH0WPYcY-I.D(8?Ed#]^)W[K#HV&QFQ[<WJJT
fA>?FNAFf4IHbA]fcB\351K7_aHcV^GdEG<^_R]W5X5M:&BN@a[,S;aRD&/LBN)@
b-OU?fER\95EEQLE85+]cVfd)Z;+4Q;WG:L\XT5.C<EN<G-f8HbAVKV&F0LW/K=B
C#5B3LF6Eb.V335QSTFC:Z&]H#eJ8KXbP.]QOJI9Ob;QB2YCUG/55Q[7=Q#geSE1
gU,\gAQ7EC_SNgROK0>=99:E3V\I>PZ@K\FIbPQJAJ?-36If7eLJ]_(MMBS;eKa;
g#TS9/\5LVGY9(@LQASY9,;)?J46Y^+?>f1R,7.Rf-gM^cf:I34g^28LdWH+d5+,
Z0Ke60,[29(L;KcL]4QB7?/3\IE=PG^]H.G69>,XbH]Z6L-4O4\?#Z+?R;@^47@&
#GYN+f\L&+gId,DdVRaW,VJ4QN:6AV<>Rb?PA[L[=T0_A.@DOH7[V6K/KL.E3+\]
1C;KIBG,7Sc[=&UL^^4TETO?SK:dFID)FbLIF05,@4O#V2CA8S4O:BPWWC^P@;&2
I-FL5>-U.<X2361W-XCN/.Jb^=(=e8PXb=:CM)+;b\Ub/[7AA^>WHT;5:bCVSM/3
H22CIUMD+_0]R+e3,WR><IYK]ZN4ZLNU06a1VQ1=L=5)F=4>&MN5A@<UQL4HEEQH
VM(V66NZ[P>0IQDefGFXO?KGLGeMG^LbF;0J-6FeGR+3.ZOHG8R4adg+1;DROD,?
:S(X[#dX)d[CC@MY<O6KI7)DO0>(Ba3;X[T,F(VWX=49^eY8ZUL74g3E]G]2FZ/E
EKHCR+L5^(5AX+FMZ/EgdXM,\NK1:4B\QO-4a^P.(10/)HN]0HU_KS5M=cHP:7eR
163HC5V:WEI,WXPPAOBJFK8EeT=Mg>I<D(O^dMJC0OZ28Z:LA\BTO:&B_bBYVBZ^
E5@c^O_?W09gN+@GSSaOgWb82N(a;\9(H9GS?)LgZ]>>Z24VI6N(6#F23J+C]H14
9&1#[(XJJM-X)[e0W4aeHY+edV)>353]=QOEE9UE@cC_K(6+YA,;=aDa8](@K8X8
-IEPAH/)<\>GA7Z8JB\)/[U;^?L[JC18>:a<Fa(X2ZA16eZ9L7D((M8-;ZOG<_H8
O,/--fM:Hd79\+RK+<D2X/Y)&)ZK4fH9;@c^C#CP7BAN6W43K/<[agD_Q)WeWN[[
>/<[GgAUeaTKPW#E&bVJR+A79c-@3]L,9AWH2ZARQVFH0MF:>D^_b95@85J;3C-^
8JTS]2VI@H17-Y\dd-dO:O9(]>E9g9K+/b8)Q+DIV2S+-]5UabOd])SRUfU,3K?I
-e3((J#6>QRgT_(4N[XHMTL2N46-DF[K5FKN;_9SH.9T^8&KW-:6)b;8ER4)B+91
6/U[W.:VYfJ7Gg5V8=<L_1T=c61&=g2#2VbQ4cA&O.].c9@C8>V@,@2?RdWXRJA)
(9T_TA^>KR\66(Zb7:&Eg_I\Ef0,HZE3OE9(/bX4]5>@OgKD^\eW3^0M.EF4?,D>
9RPWQ+WXC(Rf&ZR0<=IWegD<31=^e6E^1;0Q5<c74L)W5PC[g_F@O\T+HV1;bf.Q
RB9S.>5>SKFaT+cTF@Z=8S3bEe;gY9(M3PFfN=L]RB<E-VX-B;\[bN;S/(:Z\cJ,
P6-D:aM:?Vf_CLJ7VL4^XaTK?G73J8=]1@;@#<XC8)(B:K-7=+X4.&Gd>EHB684@
@EVZcb6#&V9ZMCGff;ZTZc,_EY@eC<#aFH;&^U8H-M.+FaT=>L1S_?8,3=S)<<87
XUHc?7dZG+5:T)73W7>:8F/F98-K)79^50;,N)c7S^C:cUEf/ZaC?0WQ6J.T[JYZ
,cURDN\8ca)KPH3RWK<D\.HY@eZFJ6.e[_97XU>J[TfJYNNF.D4E>IC.>V-)dKRW
.7Xe2=X3b\<SGIO@g^#9_NAA42;UDFD4TWM=;1c+T-3.(#?/0?E\QZB5FR(CSK=f
IH/DPZ^O4WW,WegIHGcWCC4;B)F722g0IFC;3cQBRIB&a>>2^0\)/@QOMSd5\+<5
QL7_1@(7b>KRQ)8>Ee<@XP3_X?CRAT3W9K0Ng-a?CdA7&c#@]E[c@\5VY(JV)>Ze
.XQ](WW>0L=YSfO&.3F_ODG?)&CLBbd.W/a5(2/8=aBX[\L6-?379FY=?K>f/_cU
,U(PCSAZ\AVW@?#J9FbTf+8TH[AP\>a]eR;;d)@f?.5d5eA>RJ[#f=33A.#X;6O0
/DL\TSK6;+X<Ydd+5ZUdQ6K2O9^<D??R3W64FgQ;\1<b&IgRE2A:NdBcIWI:CgOO
0E,&5</1K2(cRd4:XN[LM?O-[:bc8MQa6Ub=,[PX6)N/GMfcfaI55/Ka,WEN[<c@
G[[0@<4459,@PIdA3=9T(1BA95e^@H>,V@6?1YO2b5.I^-:@7UST@XFY@U)<5Ya1
;];\NJ9QRbO;[e4ARXMaO>ROP6ab\UR7WNOEZ2WX#C3B&8]O8OA?Y:)/./T\-<-H
>?d\SD3aU1/TSP\e7YMC:aJN&X.MX)>AUe@9(5ET9ME,E(I,.3CSFc/>6D_T1\&d
OE[>;\2O-PcATVHWaYK3[-:XB.C#Mbc:&AL^7\F0aO;UMIUPB#ILKOZD7<(SNW)-
cgI(f2(,Gg4I@/RcXb^5+KL1X<)8<WcZ^+91/RcWfH()0,8HKF(\6H=dB&a@aU98
e:KC&@.6>bI.1V4:W4d4KS1K[(=0-7]BB(CDN5EaDD\9Bg)Q=U<]R7V(?\[0g7MV
P9NESRY;O7BSQ-^J70Z3aUI3gDETIQ9^/b63A59N.;<=FW4=Z/dLfCR7IW4g<XL6
/0[Gc^Q2TJ#ZD?f@]+E_W;YUU-1/R1;Gbf_WK)aTb]J1HLO;Y:d]>DQ1bNZGYb/+
KS1.[\>XYVP=QA/C-BE9Z+6&?+g]X6YJI@E&?/OLc^IN[Zf9^+.>T:=+6&gJJV2:
>,DDZH:gf8AT3B;15Qb&a,3953SK#HC=<D5.a:2>B2O=?W[+H;^XIG15=B<-1G<G
/Z9ZI>1D16+DaBN;VSP7c^OL09TE4CEMaf3@9ff#.S9)@.3^+edB(:f:K2&N:EZR
8R?&/AL71Q=G[^CU,gPO_fMYHCGH4N4Q)>dF&]Z;-69S4T#1e7IGXdR133)>ZOgO
4V;S;R1\9+cW7N)<G4N?a,b&]O7B-_>QK7cV4&EB8XeNY\GA)HI)0cbQJbU_8Z4G
D01:\82I>c24c.Ce_U);KHE?#SO3F<WM-E3S;8SZd0[_8b#5Z9HL89IO#aC/YX[J
a\ED)eY&6UK@>b0:RZD#DR5<?2>AG49>-3aVVYAIAJIKVT\<PG0/B?1NT0eY[>+_
PTMWa\)WT<4>;?8cBCe#/V4)aR2E5@K/S+#6GCd7efAYQ:eCT[e;^ebA<[YbgdJH
f8UGH[O[,OM0:N?CLV4L\[GccA4M&b@D&S+;X@I+4f=-b8-IS\R1QV=J(_SRZfV^
7RBLUI_La_cADLAEF])H,4JH0Ng-\LcCcM^;+>SOVO55ITN26[^[4))Y@a\OG@c#
I&9R,(2G?-L;c69-#QC8.>7RD<WWM-3=)[eH@8@#9M;.(7\?ODdP=dEE:G)b87_f
3:a>(<_YO8eYf?FaFY2[<KU>[8-b(.c:D:LgQ2K^>5eS09E^OW;@,\.AYBMF;O=0
bT/KgUY6.SPf\,B[4:#e:7@MH:)g?:gN]H.3+=NFJa(6W[?VLBQaUG4YeV>G&7D6
79]8JScK[?,\Y>E).R<E:(<5V;3g+_aNHDD^YTPOGN>5#F+2e]gc4LA_C4I84<,>
_HEdIXARN,=3C@.]Y#Xg_RF9^4UN>L(abH[CAPD[F\A177dMZ<7ffYFJ?67YF83Z
NA.c6=YM20gQ^c>MbCA)b5GI?62G&HV)4+5&6gWbUOY=^&L&2,/^LE9E4,I\E@,.
RYMX?WWX&LXU<Yb^Zaf-Id,VbSe;Q]6bTT5?JO&P.CV23d4@-[P7b_&.T5I1?A)2
,V)O6>fcCWdY=ERc#T?4Q?6b]/KW25Cg-(CIQ]2.eMEWN)ML<JF4<D<.c3:CFZ@^
CM6[]L[9:4E<:2Q-@A3@^5fGgZbQI,P48QUR;YNbZPA.D#V<1QS34bXI#OE[D4U]
d6IJXNP_5,/@#D#fGC,I<d)GHc7-JL_dAeGE8#I[R.GQ2-?f/M)cXWVZfWY_fK1e
.)R9X1cg:SZ9.+-RMcaKMTHcUV.=d=EKH90QbY;4FSO;PTc-Hf(-,,WRO#3B8P.E
Fd17&8I>.^QPSBeE#=VN@/MGZJ&@DeS4<J^cC4+OJ-X+cW&^-+B01Z.(9=CHbZ1S
[<:gSDe<a(L_^7UG_Z>IZDAM\V]U/@.]@;]YdeLA_2?b.G/JGa@0N#N/?[T,N+JH
]C\gBX-XVCe?6>b;FK+/5;Z_1NF3+>-L9$
`endprotected


`endif
