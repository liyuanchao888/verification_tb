
`ifndef GUARD_SVT_AHB_CHECKER_SV
`define GUARD_SVT_AHB_CHECKER_SV

/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */
//vcs_lic_vip_protect
  `protected
I?MG)-\?:fHUCI]T@#DQfU<fW,9dF+V,f_E=HB#,ECc_4/D[=EDc+(1OHd)+_LU>
0)D8QCQG?-WT+Z2=XEH1_\<:.Z.C=?[&L&3H,,3P1Te(T2>4L2JY;[S6ee,eW].8
D=eQE^b?XW6U;J.5O&c]F&]e0d@R/fT>cM0<BdSe3X.U>TT.7M1(gaL;O\gC3R9]
:\FC>JGSN98]+-J22LbVUMVL(;W5,6Kg^285OfL7R\0H^(g/cN0]BIO+<4PQF5UQ
BX\\eB>XJJDP?+=Ac^H5)AWfOFP&2Vaf\\K52TE>S?C34XDE>1@>bGUC&+9BY<?X
FDU+<^1RR;:R>cRW17J=Za+]4KD?Y3.(IX,IO++]&-Oe\A(b4eE[0QT5)Va,F((:
VBNRO>\Hd)]D=:?JYXB6,P7;/WNNJ;f4/9G]CMA\RGP):D9bK@#D+PM41#?2,,.X
=GF\N,[:?]^O(GcWP(R)W)8[W@@BLS.^&;YC7EVK[&d=N>\->b:eMWMOP@<5eP6&
(93JB&O0BB-,0dA(H0Z,@d,dI9&+g\#-^Q9Q_EZ3Z:c=J7+O+0[#ZXO\_I+-<[cf
K<2U#H[4<(2NE>K<9_@):[gIfSJ+3Y[G<]ZXbU7,5NC;bG#Ue#L_D:#P7>1eBI3T
cZ5HG:/Y^F^1D75Q7VCG3I+B,N<I^YM0OHL.(D0A;4WJQL]),RW@Q^I6PPg2QU1.
HPJ]8Z,[Od&KLdG#:R(3LG->AFfBa1Fc7U@88ATVbXHQD:Y373<9A;XNJN+\gTOM
&-eR1,FIUKN&[FcQF@];3.]NEPcEa\N9AQ->fB/JSZGS)B1fFfO(aa<Bg9g>&cF#
G7cWQ6UBTbE.NIV-J^ZZ1W+VfT2Y>>eYJJS[Y@DOJg=7KK(=#=MN>6.Vf+WQNe;<
GA.I:T[W?b3A(VNH0\d9[V7>0;,A<@:H8:NVe_XC#cAe(8F>I5^a+(QO6If^WHV9
aGXJfNE_R+/=&aY7G>DT-(F;2>.c\NHg<8]4B?Cg+C9;Td#A\-]6B1^8^H3R1B97
R9?B#BYZ_aaA#X^#bOT=U@YcgQ.,E#/6,.BYCP(L#03)6\eD-:@)3]#J&Ze.T-Y\
,H9Q.aR@eO-cVCN-]A4B[O)S7N[-5f-H1CSB<?77f2?6Pf\7eXRWESgdH9P5B^>S
]?7+/96MJ+&==>FDGbQ4VZD?=2LdE\H+bTECa_=)0W6AM3ff^a2J47aOL;P4a4B3
5G<PfW+^(]Df\2MeS@D&>;3-9:Qf?Qef<7g5e>4WGUPYUC-]#d4^8.@XMa^,gYM?
#P>8c60G8C[-\8.M_V1T-I#FT[WMf3d23&M6V#a9g(/[/a;Q/1c31@VB8<XVI6,c
V4H;1#X..>I1fE+34/FB-98COA1.26PK>G,_fa5\1=2B<L30#:>X#Qf[EH]TLQ0K
Zc)^.@a>:(EXVf2;WK(:@_0.18P//.G0C2@aH.EW]/WRV34AJ_9^3PJ;#CT8A1O>
YaH)@>DHI(-ET,9M&B\8Q+.Wg=R(5]G.SD4N[cT=3Bg+N2[d5_CH\RRf#:^J=LC8
WR:=4,KA]8MJCD3VCAFBS#MaQSQ@cY?LI##-9-FTcY]LaNJR^=af?T78e0@FIEM@
X.VQFc=LRY92/M1TVe:(8E30Vg/X7fd<,_0X5cWEPGM-f-XFf&<cN&;H>\XHOV.b
UWg(e2YSe-b3c]ge?@4ZcbVI\4I^L[:UU++KI)MQ-^5Q;XC(S(D@_8/+>b,[2c4c
b/^=-_#,H8O/&PX,DB^C4N33F0:8fE<BZLX]S5-82);9:<_c6+U[BQ/>17G&OM;Q
W&Wd?IJHC\ISK<R7H;&Q;RO2[O_ef(G/PRI0IM^]X=ZK,77?e]aMRK@9dS?8^#EH
D[17@,.K5VO<]gGOef&_WWg-8M3E=.S/Z\?4AF.^I1BWbWE@Dc(@&Y1G].eBbN\g
U]R3K]7P9HQ_P-:/R94a0/?R]FZ+653(36U)C-=1c_b2+,PTNZ)fLKOT?4Vc\a/F
9^Y3e/LW+V)bOL>S]]+?GWVYEMQOIYF)[#<^^D6Zd/_\dOC#&ZXd6ZRaJ?.\KS[E
+5PBYfMV#c4#EcHg=X,3R_a3abVQeV>05-E5WBO3HD&Y+PdFV[U2CBIK#:YZH1HS
P[\NG1Q80TNXWNGOf(?0#Ya.AF^\8Kd5]\N-_#-ZP.BdOd5:b\/WA<b;>0@6bX9:
beLbNK(K^).]=,.((LA\P1R?PWcOHC7DW>Md9fI;)_#aFX<MOBF73=Gbg@dYf(XI
NISD9:=-Fbc0gO@c=&f.I_HXHEd(QaO9YUf4d4fD@[F.1LZ3]cRXTCK.5A3ET&?_
T,P0aI>9TBJ@+4;AbY17_aQ<-:TAS=dO_9ZZEB,G>@1QJ(R=JAc[Vc1K^\-3/f((
fBK)0ag1\N]^7N<;;\;c;G0LUI9dWJ-EN]CE==/6116T+.TCZQRA+<L0Qg.GcW(+
R.PG-eHEN\G?/8d]?f:&;.K<GLK#J8_4.L_<d<3(,=f4fQ1d20CbEO)N[1MUTc0B
(Bg9K\#,FK4\]TB6)_8S7_NWM;>Lc^T-DaPf(XU9<Ra#b(I^,#P<M@/X+36NW6/B
a7NG\#Bb\g=]/[V@SG3d9P->aG:#V8T0]VgAf4fZc-7OB93#ATOB@aE(Ug//WRVD
+?bGeAa)_RBC7K8/;IJMBUD8dNF[@DAU&#>96fgf@f+NRBQaC;#E@/GRZR6?@1bM
d#_<W>@&IO?GJP@02?MTBE8LD+C(GE9WbO/V4.BHZMdH6MP]A5fa4-^SMI,^?a5^
;HdZ0VN>IFEfHU>3CA<8WAFK[9#b5K88#VE]b8KMA3d&>N24UCFI3@3^a6C5L++9
1cI<VId:)8+<acW2-6G+/Sc5b;DP0e\fZTV5NgK^D<41>9&g@@)aT]S&6NbS80&3
51N)>_;8FbWQN4[Q4=T+^OZ[R],2S)V:=WA,b3ZCHbcYb@]NXb_G,A<ecB9]gR47
R((+-D3S>:.>A8d@^WP/O71J7]2bNOc>QFfScXcfOF/\EYR;YaC;]2&N45]TEL(+
<LMEC#[,CQ0<6A@S81V7.CC4H8gI,Y9N<@-Nefe5@1-_AY\41,aQ7=.YRa#@8K^(
J3bSHO7+&G62gBb<369U73MI=U+R9(P?L_P[:?3:KCFEXD93CBJ02.BEb5c=Pf(+
G1g,8E<YS>U=.OVE<fWdg>,f)YeC(_a[,Y2)FU<#IdC2;ESM/UH[e/FV0^L(Y_(B
e@^F=+#&5@S,b.77KN[WJ_.SY/<4&T\W(AXLf>YF,M?(WCAIG.X0RJU)g1P(beX:
H][bPOb25bd#5/(YfKCUWL_Ta_eZ)U5JKVRb1[ASgB#3W0]Z3Ng0NgHR?<J;)^U+
@A<C66B3XN)EL;BXO,2J[a?7G_O]^4/CGF11IV>DFU7?4BZ_.O@=S;(Ic,+^B](M
gMT6WeDQ\UZ[J4/>=.eCe3@E.Q_:SF86b-]O297+[>HKe-4d+#J7+8@O(332,fd;
e:50;U4[^\GG<d>g>aYMIU?,7#&XbGG^c-P;YI<dC4g5Zb0-G#.9=9gbb?T([;HA
aTeJ<IWfKZ&PL5-&RA<&N2AU@5BV5@CS]B\HU;7FD@@GK@&PNE2HOg5ITURT9W^\
N?6UCe-\;K.,]Ub-P1U3E.;P+#7IDI1,9D.Y(YFH+7@CK<SI7DOAB3G;SRSN6O@M
1d4:+M\7BC=0:#KS7Y4UYOf+(F0C<LDY4+YCfYM1[ac.]a/?[>]#]HPC]g0YA48Y
.8D:Q^K_ePfNNL&//b^^@&RJ/(HWQ(O[dQ[AGWPDCTU-(/JM_c1^1#C.YR[62I?D
10WZ8:U7=A<&FL,UfE_WLR[+c6FTF=PYf,Y=^ABKX3;9Z+:\/D(Kg6()^3@)C&Y/
OP.,dbR2\b?.R.0E?(.,fZ<acQPX?34YfPb/+ZTD1)6GdE]]H(gD,TA^L(?N;_<O
#4\UV9<^fOY+TOH[YM-Q+fcR>SAN1MT>[,I@g7ZY@SU]Lf]7R+PA^N+XLAXR)b)Y
WH6D=>NXA7-;KV<^3U2Y6HL0RJYA^,HcC=dc7F(::2SOdQMTP9A5EfCgWOU9MH.c
;aGBe8;?&+g1SQ<QO4L7).SJ&?)2e7X5?O1f:5eJF=Xabg2/dgKY<&20\8&6^=/P
c(TB9)VfO08_]aXVYN#E<.7.1T.1O@&GgVQ@DXRT>9[,(N4^=?[+dA[JU<TVa-J5
J56R4O2b(XSP-RSe?G,ABLIa/4U95XKOSDb^I#>9GNFSP68B,CX[F?ID5BXAMDRC
-g<T_^bVC63/L>V_&1(A=<[D[P0&K4)CWT(F#CA0JAU.(BE6@d:Z]]>WJCPagETA
,[(@B#I]NeGM5NcW2-HV5YB#NIebbec)RN3#eQ0EP-;6Rb>I<OS1<GaNIcW/,2^8
_4,O6Eg6Ag^LOf=)6K8Cfa\C\V44):aK4IO4fS#f<1C&C^7LG<)4]9RT;&(J.=V@
5D?TB]fX.(CM>?3.DHG0=BA=/#IeSJf2@;dZ77+JWOHJ[>eGQOb-J<&R\[BE\^.C
/D9=X46Pf-.-[.).C?@2ISa_4_J?B+1JX6OP<;#ZUTRSe[493K?eDRbRRU?/O]6D
e^URYB&f?R9UP;\ATO0D,Q4<]Q=<L:Q5VXXHcD+PMW9((P0N_8/FHMd3\\E<dG(\
:>\2>8804)HDf,c(7;G+J_8&:2OI6H\V8?KEB()]4Z3AHFUI9&X2&-g\&I<>&fID
=NR_>f^/GaA\#G3JETK1ac^<0TDW6c@07+ed>K<]54:D;<PL1^CLON/WTVb&+gb3
<E\;KbSgce>HBFX9NP@f2a8?<ZTedgWc[\AEf(Hde<X))ZG)LP7g-88VXLf,@&H_
&H.A]TH8T0>0.)?4K7.CX9Y2K:32W?35Vg+OWSa.H^YcAMMLaMS::DdCI]W3C9]7
G3[7_7&(YMEFDY-Pb9f64915Gg>B2++;(,fgKR_Bb(ES5]8VfL#>5G-/0ea]=,Ud
C>e.CX8X[<0d^b00aD+BSK[dULSVL)@5GC/:=P0(&@2DAU,SgXM5@_@=]C3:_M#F
agTJYO4W;BXY.2cg[,(0[:HQ?\e(aMafR1TN;&O_^;L](4ZC@0<O;Y/c6aZQ5P<K
3[d&,Q&DIM8FaJ6T8Z/dNP^&f>/Q]d2=17@7,_=P0?34\J-eSeH7KaKM9_HCAEBY
afgGL6MU6+4/QC9C[]d2_MH\.NbW.>S3^3/QC==Z,QC261AaQ_Z#a392c#?9&]Bg
Oc+SdMMR7#bHLY-DYQC9(QI?SH2+>E-O,,RO:#>\2>5aB4KccX6Z>A8.9KcX<e+]
_N@BOEIfTD)]>::UD27C_L[.AYE)R+e[>&-cMJa7;18VE\/FQ?_J4P=HMTd.eAe@
0FW]()J_dDcN/V6IWb6/@[\_bNW@W?5GeE.Q\a)FXC]@<eC8Q&[D4SI=VOc<aQS-
V.Sf5ZfORCcf&cN=&XMB.KQX/YE8((_M<_IO=+3:E2RU+XV_9BW,,]5J+Zg)#Vc8
g>+Q6MbK?//5MG2.Ud,NFNU(TSBe#S^<VbEX6M)4,@@4EL-3UaSTT63JBY2BD^J>
1Eb@4T5CfY?&:B;(aL+dZ;/e85eeeDbXNaKeg]9Y-?ED>&(1_:7f&HF4GP+>I+K.
\P@B.&TYSH(E_7+<3RE.JbZ8]\&-G;RSEXVIYGXO@+M?B\L=2X5PP2P@Ce;U7BFI
6(D/8_d#GEe?(UY+F#a:g6;)Vb/X\(\OR+^ZKDJ?V]Tcf;=T7>3CPI0+8\S3^3W>
HNL8_[J-GG=HU;B3HWWV2(6\_g3<=J0)WW/S5?3FB(6&S&;2GC7QFX(.GII&;eHW
OC6DMA<Oa(328NeGV\0G-@TK4#)\>(J.&5TZS1Y[F6F4-OdN:Sd^^LTA.J9f]O<:
9WA8CJeJ36_4H_2X).JC9\b8.U:#E=X2@]_WG]Z4F[Qbd87=NVI81d(a(b@HI4bK
WT-g6d()V23HI.J.[dC,_5K3Zf?bZV7OfG#Q/8-6UHg]AIVEF>=P\JW:#>C7Q_U/
[g.VRe,N(5Vd1AV?.7c^Q)_,^Q<]fHE5-([<;Ra(G\3a,c.CW-C]&G8#9L82.a.+
gE?#OcL?Jcc8:-.f2SeG4CTVf:CSe3^^<c5;;1_(8\KdZ5(_&JaL>&BgW_,33<S.
55\dS^_;0aK;:#RO7@,1>=3.L^:@@4=<W?L3#QVZC//1+4(R8HZRDce6:6VA=[3@
I:aZ=]_R-]_Y.cNA]b64NB+E;V7dZ7>4TW:--0V@6YOJNVV&K^Hc;e>GTJID0dG/
=MFJXB<aV_DF5IR^]X4@_1\Id7I=ZE5\VbB.,<);@g3&LPSF?[&aDc,ZW6bR:A#;
]<?#3^WV.bS5YU.BZccF5LEN1D/Z04U1K#fGQ?E@-fB&&M6L&S#,>#Wb^&EbP]UH
7RZN^M+W]+K-#e)/O[OREQ]N8RgcXZMB>N71@K64[;G.^XIc_RX]GL<UEfGO2WP-
ZVILc+5O(B):c-Ug.RfR2FH7P:H->PRICI,?b6aUK;DdL/KU=b7_X,95[K3P\BIb
)RF4?X8;1ac3NI=b4J^&EU9),eS1cSf7cB(]UA;\e^C):C9F709OFCe=75\WZB2.
4GS&PTXJ@+^4aI=/OCA-VD.P_O3##e,7.5LCeBf/cMcQ6/[9+P>a-]RF_b-]d:Fb
/WIH):M\5bd54F)E_WQDaF6;/Gg9Xd13JP-6bM<5B8,,[Nc/6R370GG1,QF?;PL^
Zg43L\0;B&)9E?_O^2Tb\-#,-KKZ09:+B43WEQ;FP,MPBQ(^-?W3&8fPRHc^\]Id
K?)VS;G6Cd+]7=[/I(GQJXU0DIM=@LF6>N[C::_EE/O)ZHRWFY&>U@O,7)5#]7)V
8[dD14CL8b-,=ED1;@</<T__eeEb9Pc1(6)^4S56RB4I9TKZGH&=);2AV7]U93WH
2ZNVg<ReLF6TWeNWRCE>Ef(\1@11N5@T]WcW&7S#bZQd;C,U6Wb#8PLd8J;?0e@-
:<_@?CJ&HPG9,)<6_O_UT)gKf;9+Z0#38((SXSLg/D^[MZ,X_<5;EG@V:?e>,1e9
Wf)D\EP.-KfP:I-R1S/c]T?08IE&54-PFRS50a[>,,b.Eg,@I#U42d:ZLg5)ZT)S
K+[W60VBHZ7cC,-Z7>2D@bLWI+d^>c23Y(#+PH+8+A7V6-I#/1FKTO+:&>?Yc2H8
DCZ15TKJK:H\K0dOZ9:>?QCW.K;5N/V(CL[38A?DLK)+JYI)O519<8Q+GM@N\>89
d^MR>\aZ;RPgSW[N33GMI3+6\T61Z]V[X;I<43DF@9^b@6L3d/,T.SHf6d#JP.e_
[5bPQ/&RS8Y5HCc\P>8NEIc/(4K\MdX6-a=CAUSWZ_,3/_ZcJS\PW2@R:H1a#/0f
XJBOMb@:b^(:e6V?G@FY8IVE02L=MdC)Me:GAF14eU7=.SS;JBa59@Q+GJ;@DK^&
,0)]C3&3CGgd=5WbPW,.[e5AU+>\8VOD+U6)1\\IM4cZ@V-/CX)fbEX)5O7dK85K
=?(Y;VOZ29D8e.ae=:(W1^,RKI[L-G7H=eH1D[D_V&5F0&AEZVMTK952/.P9+@W;
W@H1J:JA[>6QFe/G9[VcX==QL:8feMTcDJHLMKBg(?S#LR/+9M>_P@(ZePUEKCG,
@EdceVI1>,IU0D:E@],9SCCc?-g=EbfMR,B#(A;5RE;/)f>M+>Gg)E?QH;3g9VKP
P,##8--&(K2>(E,5QL-.AU?,[a](fDf3@2a56DaNU_R??b/>/9,-3[ceW6Fc2Y#O
?bD<3TEL+SgH<2caICM5?YC0/We[b.c@D)Mg/-9J<OL1cZedBFe-/WYC:&+-<>d=
TD:7D><d7P-H-$
`endprotected


  class svt_ahb_checker extends svt_err_check;

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

  // Signal level Checks
  //--------------------------------------------------------------
  /** 
   * Checks that HSEL is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hsel_check;

  /**  
   * Checks that HADDR is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_haddr_check;

  /**  
   * Checks that HWRITE is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hwrite_check;

  /**  
   * Checks that HBSTRB is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hbstrb_check;

  /**  
   * Checks that HUNALIGN is not X or Z <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   * Applicable for AHB_V6 extention AHB_LITE
   */
  svt_err_check_stats signal_valid_hunalign_check;
  /**  
   * Checks that HTRANS is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_htrans_check;
 
  /**  
   * Checks that HSIZE is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.  
   */
  svt_err_check_stats signal_valid_hsize_check;
 
  /**  
   * Checks that HBURST is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset. 
   */
  svt_err_check_stats signal_valid_hburst_check;
 
  /**  
   * Checks that HBUSREQ is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hbusreq_check;
 
 /** Checks that HWDATA is not X or Z   */
  svt_err_check_stats signal_valid_hwdata_check;

  /** Checks that HRDATA is not X or Z   */
  svt_err_check_stats signal_valid_hrdata_check;

  /**  
   * Checks that HREADY is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_check;
  
  /**  
   * Checks that HREADY_IN is not X or Z  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hready_in_check;
  
  /** Checks that HRESP is not X or Z   */
  svt_err_check_stats signal_valid_hresp_check;
 
  /**  
   * Checks that HMASTER is not X or Z. This is performed in full-AHB mode.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmaster_check;
 
  /**  
   * Checks that HMASTLOCK is not X or Z on slave interface. <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hmastlock_check;
 
  /**  
   * Checks that HPROT is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_check;

  /**  
   * Checks that Extended_Memory_Type supporting HPROT[6:2] is having valid
   * values   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hprot_ex_range_check;

  /**  
   * Checks that HNONSEC is not X or Z   <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hnonsec_check;

  /**  
   * Checks that HLOCK is not X or Z on master interface.  <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hlock_check;
  
  /**  
   * Checks that HGRANT is not X or Z    <br>
   *  When svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1, this check is performed during reset.
   */
  svt_err_check_stats signal_valid_hgrant_check;

  /**  
   * Checks that HREADY output signal from bus is HIGH when reset is active. <br>
   *  This is applicable for:
   *  - Master in Active and Passive modes
   *  - Slave in active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_bus_high_during_reset;
    
  /**  
   * Checks that HREADY output signal from slave is either HIGH or LOW when reset is active. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_during_reset;

  /**  
   * Checks that HTRANS output signal from master/bus is IDLE when reset is active. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   *  This check is performed when svt_ahb_configuration::signal_valid_during_reset_checks_enable 
   *  is set to 1.
   */
  svt_err_check_stats htrans_idle_during_reset;   

  /**  
   * Checks that HRDATA/HWDATA byte lanes are selected corresponding to
   * bits HBSTRB signal which have value 1 . <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats valid_byte_lane_for_hbstrb;

  /**  
   * Checks that HUNALIGN output signal from master dosenot changes its value
   * in middle of a transfer. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  .
   */
  svt_err_check_stats hunalign_changed_during_transfer; 

  // Slave Checks
  //--------------------------------------------------------------
  /** Checks that RETRY responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_retry_response;

  /** Checks that SPLIT responses are not received when configured for AHB Lite */
  svt_err_check_stats ahb_lite_split_response;

  /** Checks that only OKAY responses are received during wait state */
  svt_err_check_stats non_okay_response_in_wait_state;

  /** Checks that ERROR response completes in two cycles */
  svt_err_check_stats two_cycle_error_resp;

  /** Checks that XFAIL response completes in two cycles */
  svt_err_check_stats two_cycle_xfail_resp;
  
  /**  
   * Checks that HTRANS changes to IDLE during second cycle of ERROR response. <br>
   *  This is applicable for:
   *  - Master in Passive mode
   *  - Slave in Active and Passive modes
   *  . 
   */
  svt_err_check_stats htrans_not_changed_to_idle_during_error;
  
  /** Checks that SPLIT response completes in two cycles */
  svt_err_check_stats two_cycle_split_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of SPLIT 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_split;
  
  /** Checks that RETRY response completes in two cycles */
  svt_err_check_stats two_cycle_retry_resp;
  
  /** Checks that HTRANS changes to IDLE during second cycle of RETRY 
   * response */
  svt_err_check_stats htrans_not_changed_to_idle_during_retry;

  /** Checks that IDLE and BUSY transfers receive zero wait cycle OKAY response */
  svt_err_check_stats zero_wait_cycle_okay;
  
  /** Checks that if invalid HSEL is asserted for selected slave. This is applicable only in mutli_hsel_enable mode */
  svt_err_check_stats invalid_hsel_assert_check;

  /** 
   * Checks that HREADY output from slave must be either HIGH or LOW when there is no data phase
   * pending. That is, checks that the slave cannot request that the address phase
   * is extended.
   * This is applicable for:
   * - Slave in Passive mode
   * .
   * 
   */
  svt_err_check_stats hready_out_from_slave_not_X_or_Z_when_data_phase_not_pending;

  /**  
   * Checks that HSPLIT is asserted for only one clock cycle. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_one_cycle;

  /**  
   * Checks that HSPLIT is asserted for a master that has not SPLIT earlier. <br>
   *  This is applicable for:
   *  - Slave in Passive mode
   *  . 
   */
  svt_err_check_stats hsplit_asserted_for_non_split_master;

  // Master checks
  //--------------------------------------------------------------
  /** Checks that transfer type of a SINGLE burst is NSEQ */
  svt_err_check_stats trans_during_single_is_nseq;

  /** Checks that a SEQ or BUSY trans only occur during active transaction */
  svt_err_check_stats seq_or_busy_during_active_xact;

  /** Checks that htrans does not change during wait state except when
   * htrans changes from 
   * - IDLE to NSEQ during wait state for all burst types
   * - BUSY to SEQ during wait state for all burst types
   * - BUSY to NSEQ during wait state for unspecified length burst
   * - BUSY to IDLE during wait state for unspecified length burst 
   * .
   */
  svt_err_check_stats htrans_changed_during_wait_state;

  /** Checks that contol and address does not change during wait state
   * except when htrans changes from IDLE to NSEQ */
  svt_err_check_stats ctrl_or_addr_changed_during_wait_state;

  /** Checks that write data does not change during waited writes */
  svt_err_check_stats hwdata_changed_during_wait_state;

  /** Checks that burst transaction was not terminated early: 
   *  - AHB master should never terminate a burst transfer when OKAY
   *    response is received.
   *  - In case of Full-AHB mode, the master should rebuild the burst
   *    transfer in case of EBT/SPLIT/RETRY before initiating new burst.
   *  .
   */
  svt_err_check_stats burst_terminated_early_after_okay;

  /** Checks that master attempted transfer size greater than data bus width. */
  svt_err_check_stats hsize_too_big_for_data_width;

  /** Checks that burst transfer does not cross 1 KB boundary */
  svt_err_check_stats one_k_boundry_check;

  /** Checks that burst transfer does not cross configured boundary limit */
  svt_err_check_stats boundry_crossing_check;

  /** Checks for illegal address transition during burst */
  svt_err_check_stats illegal_address_transition;

  /** Checks whether control signals (other than HTRANS) changed during burst */
  svt_err_check_stats illegal_control_transition;
  
  /** Checks whether control signals(other than HTRANS) or address changed during BUSY */
  svt_err_check_stats ctrl_or_addr_changed_during_busy;

  /** Checks for IDLE changed to SEQ during wait state */
  svt_err_check_stats idle_changed_to_seq_during_wait_state;
  
  /** Checks for IDLE changed to BUSY during wait state */
  svt_err_check_stats idle_changed_to_busy_during_wait_state;
  
  /** Checks for IDLE changed to BUSY */
  svt_err_check_stats illegal_idle2busy;
  
  /** Checks for IDLE changed to SEQ */
  svt_err_check_stats illegal_idle2seq;
  
  /** Checks number of beats in a fixed length burst */
  svt_err_check_stats burst_length_exceeded;
  
  /** Checks that a master started burst with SEQ or BUSY instead of NSEQ. */
  svt_err_check_stats seq_or_busy_before_nseq_during_xfer;

  /** 
   * Checks that for non existent memory location default slave should provide
   * ERROR response for NSEQ/SEQ transfers. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */
  svt_err_check_stats illegal_default_slave_resp_to_nseq_seq;  

  /** 
   * Checks that master loses the bus once it gets the split response
   * from the slave. 
   * This is applicable for:
   * - Master in Active and Passive mode
   * .
   */  
  svt_err_check_stats illegal_hgrant_on_split_resp;  

  /** 
   * Checks that master asserted hlock in the middle of a
   * non-locked transaction. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats hlock_asserted_during_non_locked_xact;

  /** 
   * Checks that master drives HTRANS to IDLE or NSEQ when it
   * does not have access to the bus. 
   * This is applicable for:
   * - Master in Passive mode
   * .
   */  
  svt_err_check_stats htrans_not_idle_or_nseq_during_no_grant;

  //-------------------------------------------------------------
  // START OF PERFORMANCE CHECKS
  /**
    * Checks that the latency of a write transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_write_xact_latency;
  
  /**
    * Checks that the latency of a write transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_write_xact_latency;
  
  /**
    * Checks that the average latency of write transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_write_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not greater than the
    * configured max value
    */
  svt_err_check_stats perf_max_read_xact_latency;
  
  /**
    * Checks that the latency of a read transaction is not lesser than the
    * configured min value
    */
  svt_err_check_stats perf_min_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not more than the configured max value
    */
  svt_err_check_stats perf_avg_max_read_xact_latency;
  
  /**
    * Checks that the average latency of read transactions in a given interval
    * is not less than the configured min value
    */
  svt_err_check_stats perf_avg_min_read_xact_latency;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not more that the configured max value
    */
  svt_err_check_stats perf_max_read_throughput;
  
  /**
    * Checks that the throughput of read transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_read_throughput;

  /**
  * Checks that the throughput of write transactions in a given interval is
  * not more that the configured max value
  */
  svt_err_check_stats perf_max_write_throughput;


  
  /**
    * Checks that the throughput of write transactions in a given interval is
    * not less that the configured min value
    */
  svt_err_check_stats perf_min_write_throughput;
  
  // END OF PERFORMANCE CHECKS
  //-------------------------------------------------------------

  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

/** @cond PRIVATE */
  /** Reference to the system configuration */
  local svt_ahb_system_configuration sys_cfg;
  
  /** Reference to the master configuration */
  local svt_ahb_master_configuration master_cfg;
  
  /** Reference to the slave configuration */
  local svt_ahb_slave_configuration slave_cfg;

  /** Identifies from agent cfg whether a master agent */
  local bit is_master = 0;
  
  /** Identifies from agent cfg whether a slave agent */
  local bit is_slave = 0;
  
  /** Instance name */
  local string inst_name;

  /** String used in macros */
  local string macro_str = "";
/** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param log VMM log instance used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, vmm_log log = null);
`else
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param name Checker name
   * 
   * @param cfg Required argument used to set (copy data into) cfg
   * 
   * @param reporter Report object used for messaging
   */
  extern function new (string name, svt_ahb_configuration cfg, `SVT_XVM(report_object) reporter = null);
`endif

  /**
   * Execute signal level checks on the read path signals (driven by the slave)
   */
  extern function void perform_read_signal_level_checks(
    bit                                    checks_enabled,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0] observed_hrdata,
    ref logic                              observed_hready,
    ref logic[(`SVT_AHB_HRESP_PORT_WIDTH-1):0]                         observed_hresp, 
    output bit is_hrdata_valid,
    output bit is_hready_valid,
    output bit is_hresp_valid
  );
     
  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_write_signal_level_checks(
    bit                                      checks_enabled,
    ref logic[`SVT_AHB_MAX_ADDR_WIDTH-1:0]   observed_haddr,
    `ifdef SVT_AHB_V6_ENABLE
    ref logic[`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] observed_hbstrb,
    ref logic                                observed_hunalign,
    `endif
    ref logic                                observed_hwrite,
    ref logic[1:0]                           observed_htrans,
    ref logic[2:0]                           observed_hsize,
    ref logic[2:0]                           observed_hburst,
    ref logic[`SVT_AHB_MAX_DATA_WIDTH-1:0]   observed_hwdata,
    ref logic[`SVT_AHB_HPROT_PORT_WIDTH-1:0] observed_hprot,
    ref logic                                observed_hnonsec,
    output bit is_haddr_valid,
    `ifdef SVT_AHB_V6_ENABLE
    output bit is_hbstrb_valid,
    output bit is_hunalign_valid,
    `endif
    output bit is_hwrite_valid,
    output bit is_htrans_valid,
    output bit is_hsize_valid,
    output bit is_hburst_valid,
    output bit is_hwdata_valid,
    output bit is_hprot_valid,
    output bit is_hprot_ex_range_valid,
    output bit is_hnonsec_valid
  );

  /**
   * Execute signal level checks on the write path signals (driven by the arbiter)
   */
  extern function void perform_slave_write_signal_level_checks(
    bit            checks_enabled,
    ref logic[(`SVT_AHB_MAX_HSEL_WIDTH-1):0]     observed_hsel,
    ref logic[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] observed_hmaster,
    ref logic[1:0]                           observed_htrans,
    ref logic      observed_hmastlock,
    ref logic      observed_hready_in,
    output bit     is_hsel_valid,
    output bit     is_hmaster_valid,
    output bit     is_hmastlock_valid,
    output bit     is_hready_in_valid 
  );

  /**
   * Execute signal level checks on the write path signals (driven by the master)
   */
  extern function void perform_master_write_signal_level_checks(
    bit        checks_enabled,
    ref logic  observed_hlock,
    ref logic  observed_hbusreq,
    output bit is_hlock_valid,
    output bit is_hbusreq_valid
  );

endclass

//----------------------------------------------------------------

`protected
5:E>Z?aW-\L[V^-S&bHK#)Q6^E5](7Ef\]@fb#cSB7GN=A_-@g985)9(IP4GF440
TDgJJ^EP=LI\dId909]E<cTeVg4^C=f@LOFe;f3=>.&RO=9YVNXDD;L=1bY^@e#3
A1K(-]FS:-).DBb9A0f:;@_1KO4GYWBEfPH3[(SXGR1:dT:e<IJFG\PL#+\ObC^]
)>AG<@c1SKf1d89Y=[f)]T)RUg-;6I>4PfF0PQa\JaUP)AR6^cG((3P\aS,B5M:)
U>f_YSS4^>3g)<&+8DVV/X#FdER\-4GFTLQObdafCJ_)(+-bR4V.:_8,P<NKAEg3
-PfH([@_C4BW&BHSe1;JXdRcKLR3BBC&BHI=54FN:JC0.NI_P5f)5IV(NKIaJ:,;
DeeZDV_1>;=_7=^_UD330(9QcVF2@)\d#d_;AYA89;]RBH=bP5;>V+G7g]^S^<9P
dGAD#Je/[M3eP<_)Jbe)QD>]M</3PH#IHU7D4UeUGaT^+KK,@Q29YUDXNJZTd0^?
MWN:-5];8+_F<BZ/8S/30dWVdB^?Da?8E)=51a2)R:T)M)/G<U(:RNOG=cZTPTWP
SP51W@<aI[a&SNQV#\_aR>#dUK\^D11gVgN:W-K\^6L3F>:8V@1@<=@TCN#R@UDA
V?-A8S</6AY5RFHdPYd7K@D94#<KJ7VJ+OSEU_A[6OT./C(:J;J9B3&=a[&QBD0Y
aO>?]ZLB2UKcI<eF#:2<:&D\VFWF:(PaB9D@gEJHJRYK7IP0DcZAG?J.KeV[-=bM
/9V6HW_7d.H8;:7P+W\VT\X/gS)#N4/dGH20M[A0R^/[g6,E-,,N7?OJdKd5[e>8
e^D(I3U_J=@b10KKbC4=NGBC>a;E<-W?@/E_&-@fI)V+2KZ3PWMYeYf9e[F[K+1;
V[?DX4;VDJd[6WQd+^.PSLRCbIYVAO,La86<1K@/P@T)0\\0Q\EbU4#DF6<4O)O2
0c_=MTg=DG8?4@<YZCULK=/9]LO&0Z9[IT;H\_M6ZX?IO^<4KB(Q^d1#P#&O7##4
eF]SNT;1QT>_+\S&+5;G/aNKD8=eLL#6:G_]a,N8Z6NQ:,9<2,KCOd1aWLQ7B6XZ
._<d&IgfG?J;Fb,MOX\M7KfY@cT/>0EVK-V+36ADRK);0K=7gf3N7NY1<0@<DPKX
O8MI0W6JSYNX[\)936>2S;QKKN<eSSFa9[(=Ta)N>LK;QgLP1I409E:3+^566&V8
H&KgD.6DS+:[9=f?B7E[eYJR&:ELMTZ<PUUV)YP0)IK?]?HG[?8@DOX(4[U-NAc,
UaC=[:TR,/(Z>,;JL_Hf^]LTeV&fC9a3>7\JLC?G<P)+6JB@Ig5L0_NbQSAEJJa7
Q:P3>89R=4[1SAN><^3X&/c7PK0?9YcZ3BI,T,U8H/#>QECE2W.YKIN4e__a7)<1
F5@7^8S;<&^KYd,IW+:&Cc,4(]W6VJUG-#FQR\XBT^YWE;F&e+O0:,98=(^@F9We
W]a2Aed.aeAR49<DZHGC3]&YSb:]A88.>61\6<&)5>bH&G,_4;_R3NL+AZ@FVHaW
&CDZEaHB_Gg@/3H]_Y9VU)[6R0LbTUDCeSg,NPY-:5YCec\a.#272O)#.OKJGCD#
D>GbUYJ3g4?Vb3#]QU4_+SaIZU_4F7(RgCg:S65,..+fa:VGYf>e[P>0KYI<EDN[
g:M>1OJgU=Qb5?f@cY3(]SS.6P1;&dC6#c\,QHMIX0;_EgbIF2HM2PN@<.Y-#@34
OCC#5cTU)P5-GV^fPF?3cJaJ=?EWd+Z#R?XS05C<&(X66EJ+A(AQ)Q&O3N&@3<SW
=EA^E#4JHfJ1b;Q[HaON8O;_Y;H9?C/e6^/V>4@1cBI)6EEY2#H@DdB=,]@34[OT
b\O\8O[7Z6?-^J&T>^O2S_1U+D/6+@f<A,VFc=U)M#PY1DQ3>(gd1Jc3O])@B[ZF
1AVD0(S[GT\N+0@bZRB85IFa@:C0V\_-1cV>bEEP^H518[O>9:0>U/CPO\b-R/^S
L0M1cbfgg>(YDJ\<1C#;eb7DEa8Re67W,1^SD@G-.:]AHAgS>Y5T@NX-/W7)+/>9
Na.:9=>34]_00.DA.3Qa8eGQfST2,US<(BLB+B45A;4/28>I=O4bb[]PQgK2MK4a
a8X-X_f[[7=E6L<4g#@cL;SAGbb7RE(^R6QMJ+D9>[bJ7<IXRGGZQCI1IJ(#)O&-
L8ZW>NS0HgcP]fES]IXf38La#9Q1IaAf&(D?.19BLeK2>X-?GO.;WWY=e;F^PD/P
)?(M/Y+aS?&4JOe]^bVP(GN:LWZKIBeZ;XM.[,N7d3GE=U8(.Z,_JAaD63^RDN2B
AV0XBCK;4MQ3e=QFGLL6QKL7IS9<B_7KV@gY+,V6I;_0=Z4HP(&-D-E6L/U-cYQQ
/3:@_@JeI8WW<g6J,#gKX_O),=UaH?4]G&GTW@8W+]HOH?d[b2_4Z)6/KUG:UVTB
@#/1JV@Zb)LX;^N3-)2V47BJ,WQ+/<7M8L.N&X;U?<WV=Ic:,6BO5)/#A&CM3c3a
SI5.RO,R^VY;+:4@)SPQEH,fC]1b/H\&Vb_FD),()Y@Y]NUL9A4>#R<-/\Rff5>g
?K^@/J[&g2bEDaP(1-9;aI0VFO:A@I9EUgGc_R793Df>Y&17^\e2e.G(IO(3E?-#
<DD?9:&+-c3JDJJ0A5=)1EJ-14b^DKFTQO:a=/IN7>X\7L6KE]92(H?,NE@UM_;?
^a&fN_LZ0Q#7=:([Lagb8)E4A,ZR9FBVT=4V\N.(/J;2g-AC4W?&UY4&e[NLFS,V
G0a6-K&1dK.T[.L.cIP^JFQZXX7[PaB<P[T4:_^)f(^PX-SNSGBU\9ST+&N341;>
<^D+c92Q>&KB4_3ebS+6>KUK)E<c./;;VX/Q8=[PTY_B+AR:EFNW,3H-)eYW9-13
A5-W.G[5=3@/UEbN,82JZbY1c(OU4]J-&Mb\ZFTQ-ICPN[ce9SHCeAFTZ4f&LDD^
4NXLaJ:K8FHe;6ZOOV]2KUCKK<<P2f@(];^1ZC&A6D(-CI\4^<D4bcX#A?f#OO)9
N,<cg8[DN2C&.:VF8J-&,S[Q#;[Y.9Nc]K:E?K)1f:]Y<L(W>g5:c4g2TF>aC6#d
>YM5<V@SVc01J#E?R?FS+6T:KUSII_J-J4AfM<H2P>##5?d#f\4>W<465:(>B8K<
,Z)LI]H;NORa^IDc>?CBMDaE=OO8:)(L@Oe:Ud[:Jd+ea#(1_N=?]YUH93Z\)7d>
PeFCK2EW0#1e:A<BMOYHHT08F7cWMNKXeO&B&JT>5U[e4JNR>f@.V2)>GeW)Pf[B
dY[:CNQMF\:d^##5K8KaI/+.G3::]]+L&H,>(];a.V9fBB[SD1,.fIG=aL)J@B.5
XAf6B&D8\.Ub1Q571MQX/2_/CSRFBY+NV>b?IGE7S(=.);YVNUF@UM(U\:L#?HJW
C&<f4^:[_d3EKDDgM??X]gF@MZ@2@S>S7.KKD=e:TF-?1DM/c15Q]Z_WeEZZ6RgQ
)^d]@7GcO0eUMDUKD5<X/gc\^8TDgL_HgDVR-/^PZ&L1CBGGG#?79J4;bS0V87FK
_bT5FaZQ+>@L)W2V\IgZO?Q/0.I7:2f440H\MGIR9<&3CB:@g/C=)_-1gP4OCd)&
(bY_bLUO9H6H1\-B\=CK]-<ZDJ:/6-EJQB&-_SV#5)^QK\0\d-(6IX;E0f3X>9N,
-=cIa_N4RA5&GH&IMZ2Q7Y2Q(<S267G]5-81)d]K&BTIVQO,g6JQH6:<+e+<3B7Y
(YcS<GW8=G;9e:-JWQ?6Ze-RET(F?6;8ZC?61PdX+Qg6=R@_62VE\RLQ\?9]P3]W
)VME4?I940D7TZ\=)Da[PdN^O1?C6\8C102>.KUM#1VXLN;A)/cO?F&CD00LVA])
&;8Z4M77YB9Zc/bKa(e>cV#.[O,#SB,Q#V]]CcPF>HaV=_;[V<?-A8:ZeYU]V99g
9ZB9MGJe7\R?[5>#a&XdWefDPUe^</gb;T_47QB]B^,BK^7JT[MXLZBVb0<G]FCW
/+YW8Q:V.8Z&@>#96\<O#ZL:(ReJV5RGLCAY0_RP>3:EJgV=9RY,U2SF;[3X/]dM
&5>b&K6^0T(VQYf#-\N:GDb;C&8-YL\N2;I3L<2C.EK8R5R6M<.N7_6\WG>bZHL:
FL;[-bJ,FW8W>G>+Cg]+ccaW,=\aSB<?FMRP-5=UfadXB@NZD6+5T0]gX[#+[T<9
G=d;X+Q@bAY<a)3-aBd8X1F,55F8_9TEKNN:;:2LFY[fUgO<56&\DZI3W#/5Y+2T
Z,L0C>O6D&)V6Z2#GA,./[3,6>F-MRLFId1F/D?e>0\2D4+^;b(A#e4;S;U-?f)6
.I@:SHCGA+2HT]KgU5Z+B=F0@[P;MK-g;6UPgJQEIeNePR=Dd4?2,\YW[-?Uaec2
9(AA(;b,^R#V&R@HMDOJ3X=&<NX#;9(6@-OD,I-fDYe.1G=#V)C9G+Z??,&1-YfU
eWR&H;0)Fcc?&\@g]6+G#,L68M,WNNSD2FCA5=&L,X(e-2)4aO:-@7?GcKZY2c^c
C(>@S^OKI0(&52SL(a-_/[E:VUV6NJ_cVHEKaM:=RX_c_-SLdE>3=THG6HK&\f:1
L;\D:^4JSC,NfUYTK4^7.2W@84Zd69V[SK:L635=&UXIZc@S&]\Q(60g8C\ZWc6C
G:O-FGN8Ya\15QcNT55X^BR(-HPJ;7VGgLE?33J(RPaa5F.VLH[DRZSaZ5U57I5I
(QUE7H]QE,H_b:]<EggC)U0Mg\,;Ac3@X0Q[:g3(Z4FC>/IY5^]#4L(CZG,^QS,,
e\-O=Z)b,S=4Kg83+Z\gT.e>QU^-4=T4O-EKAf@6L?Ra?H2[YO4LTM251@ION^IL
[-/OC/H\+2H2&T9[=gOYD]e7>A(-U]D_((],a07[^QIX)1PPAgU]A^@07A.gc/+^
DKX+OJU7]+5BJGHJV>?b8;R_X;N5.g?<O-P3Y,,f#BTV+=J.@4^WFdO(39e;.1RI
^Lf44-.T6X]&Aab0A7H+AE(EGYb(/HWK9]V+&XDWDZ/V7+MeGKaMC/>Ed.bgfc@)
(:f7d2UU2LTS=PG(K[C[\A/a[+f^B[&1e/TMVe&OAWDYJ>L0LMJ_;+.U^\+X<V+G
M9W+3GIKgfDQaHD&a?0[D0T/ZQI&QcXG7^c&0/_44)09FWRQ=B-;R)7^+e=QG15a
ZaTU+J+K2#CeLE3SMCTNC:3[9Aa4Z8AP9M0H)2;,68E/[OVaf)IZc)6ff4b&7LSb
H7Q]M,C,ad:,JSEI,^PUK]S3&,,e)66HAfdTLZ;]&HMN#,>Y^48YAGN)YX&XZ+2U
0J9S8QbIL^A2])TDV[)8R1VQ-Z0Z<\8YC4]J_:_eUSL2,7#-bbc.1=7c<>W37P+#
^RM>)Md451VPY/G\bc)f9+HC4XdO)H.O/]eRe;/)&&JeDMJYbR/_P1<]AZ8#:@B,
?+R6L1/3]#KJ+)a2;.<0-dRA/Z.H?EH693=f2MO]d-S=(Y0-/XgD#L9a=CE7>9(6
PUR?SJ397_)MO5caPHSP^8N:/Ped\#]Xa^#4a[<76QKE/.@WKKb?68+[.T5GTSc@
X8ca@EBL1J1aEVLY1O@5;:2GSJPKQJYS][Tf9R4f0?<I^N7SL.ENa/9>OcVeR9LV
;d,#Q&G;Uf,)HgGM54<-](fL?4@U8=:e^+;P4PD,eMO@H9B?A(]>H4]_OC,d9c+U
?_ZfZEV5df08NXGXfJM1RDL,^@_PWYU/\PT5g8;2)1/R0Q\#/M/2P4)8c-Cb(FU7
:<V;3#;U1TfUG.]TEN\FG0/.N>98bI.@T+HJDWUFGMcVIe7IAA<)Z_A.[/Ue:d;&
c-AC,F:A>]RO.)F8GC#Sg,/G;F+?:ae?#WRH.A&3BdYZ<@_c74PXND;G\a9L2Z11
Z_KFd;gbeg#C4((C)aY@#?b/,04dgg^83fCZ57#>6RK+W?Mf,gFWL+E(@/,HULeP
6V(XV:UU@90HHHaV;O#aWQ^ALF5PY0N@BVJ[LU4F6WUQNA\EcTFKT[ETN52Z;Y65
LNfJW+VBPS>EMMX/DC9((CdU+MIY3b0eEgdKMDfZ0G310A/MJP,6JF,W<SRA,?cH
\gg6;<@TUW<EcC2bA^L)EM[+?<aI_OfFPX)7#3S1Ua@;Tg229K?R1E8d7FEE,NXU
V?cd[[+GIV+-Y#_b:3ZBFe3aX,TW5@0[-gOBM6_#CG5^T(=LgHO9gYV&d&bQR^^A
Y\9Jbda>;aK)FJ5-T2<d+ddKC]b:F&J[&.4BL,dXYBERNR)BdVD75gSRH[c7BHGO
_e>T#-J5\Y8G5S?D[I>8\?7Y+&ZRYL,?D(F-J.[(PN98F,/gKE>H\71)JBV1VaCg
6@c_B)(S:ZcYJTF#5YI/[;_Cd\_X@JOT]@A2&<:5;g+?eY@&5.IAe0HDWCJ2bVC3
:]26[O;KS<?-)VFPc/0W;6^Z9GG=Q-DM<3+D.08-;d@].;2^=GD2?5.McY3J3M^_
Kf,76GX(V/WJa=gWDb.^C<<)Z.@40dGMXDc4_S^J81OANFAJ;A@98J3QT^?\[-\#
P2P:KJ^HC.UFaDP5>@QQ-0QQN[YbT,g@&1efPA:3R=3Y4/R>3,(aCVAL5RT5<@g3
R1A8;2KAOeHBZ3aXP>MGNO2;@e0Q]\dSbD.0.MMLR8]_4=Z0Q??Z]@aZE]6egfcU
<&;L3&U&2IAS_R,M-5)PCDM6IP9?X:9agY]^20^1F9L05QTG7D;8EUR<8;G@17g,
R/&ERcA,DKME\I,4RC=5>OPHVH4?baSEKUT+7,AGXbcQ<DYAF[12TLB0:43_#aUZ
IF(TC#5-32<\:5@HZ#N@68M5/bG.7T5#:14A>c-F7\U^/?:I?RC9JI@;d\+<K3:[
2[fK0L-C,fe@31aTM<^&(#)]AfZ,/#Pf3VQ^G,WF:@H)/SL,,LU^-9eUb,W_ZM1?
)>SR;egJ,DdHIF/H=/b>0d<K@(ZO,.]Q(2fO(2\WLD@).)=[^2@g&\e1\/;5T42f
X?O;IAYQAd>M?O&Z8WHLTO(5:a@7/Z2I[??-aEWAME#::4aE^M&g:_R(f\IO&F)g
G.&Q/C?U@.03?\K>+BeT7R65NF8<E4]8G92BDLFb47f2ZTb/21QQT<(S7d-9=+3I
J;+0CV)]0@K7SI2TTGd[T&[3c?+4BW]V2+PCGdZ-&E_IZ)Q4<R3#aJaR6TRNMJ<)
0G;-SC]+#XWKQUQ6=5>99F44/7D/>_/bDOO\F6RE2YVC@>YCD0^:;3(?&7[N>_gP
2@:V40)I<2:J9WKDI;-b#,PTPOIdPfV(?>+3R/]F3gFaDT7,#f.>JW#QHC;JHeQa
\9d6>+HRDSKF4f/PTVd<UGV(PK]E#M<S=63<K0T?[&);DK>GNZCbZA>_Q0K?HaCY
H.-8PM_H(ABN_WQHW?PK/IM]V<2@1BJcM4[O2g[]HVT[RZ^#Q],,,/X\6ZXF#(;S
+S9e4UNeOCdX:QD@Ja@OdB<#)&0M1C)D.A,@>#2BC-1c-;L1de\;0KKK/VFJA5_B
;\V_@R<Y@A3R2bVb:fdAM-\O-g5g2V>d+QGG:XH[[g528g@Rbb0R+](QG_gI;BJ=
5=[N=72YUgd()EUMHX2T=X169^_8FVf<bgaBXQ1YQ0\f:b];V:Q,aQ;GB0K9(W8)
Y^(8)-bT4^UU/9GTEcR#Icef^((ZH1T=Y-]bET^Occ_Nd<aH(.DK25KUCG_T6Q:;
_]O2E>P^:R-&dCRGeYZ>Q01f2Da^]2_FQ_\9gBV3g(DbeO]<\\J3V&+_VECdY+f_
[G?893PZ2_7M:9:O4__65)LF.3JS>.^-J=^(:8-V[<E+8DZ-bCIdfV(W;F+b1.fI
SQ.A]eY,N3TN/K@1,dEDeXV0+:8Q(X9P-=N/63;TA@eU742.DYK4[Tc476PLFZ6^
PA-faMB5YP_@a_WdY+U?/S0K_&+f[Q[:(TUM@0/(3dN,e=2fVfJDYD?S?DUc-NM:
T5;Y)/0SY]WP>-]M4=VY&:FP.XU;(WcBI[K/Xb\UKQ@HHOfD(D2(c<aNIcX2]Nc0
MPCaR\P#_9S88R9Ac@=60?+,X4ZN#GQ8.G0VD:a5BdLOMPB8eO-6ZNSg]91OV+b3
1P-UEMdR?6N>\#N0#<Y7Y/;<a23R:&3IQZN5VI^2D1_5.-#ZB?&Y2J8=Md40bORP
OI-6[Ge+D@G(]8LRMHg,NN;7WN<IBTP9,Z]^#4+Ze\#f^#+WSb?USV+XCeQ-=QN?
D&W\M+PRaD9-RU]XP<[B9:+1<@?_R2K;J-TOEE9D0^H(C2X^VcV/BI+S>[bX@\-3
2BRKNU>NEB]ePE:BV9SP9OUKY\NPRe8#>.MEVN1@f>d&1S>9O8_+?+D>)LWe(Y,b
b79H?AV:,IfIROS\?YVFQaR6&eO<N.FXRQ)8XS]DC72D:,+@3=&4,<7[GX/-ce,I
P4bI<7WM,M.(^B,1]Ed.d,@=:#X07>&9BT:)6UZ&7Kb]Q,g/U<f,f<S#:1XU-QKC
bE6DBZ3^5L-FB]&2)JZ9J&:2>P=4UGY>RIfagOUGE;^Z/=9JJCYaFK^Va#a&FeLB
HcLX05acW7(5]fXWf4I3^a>)>3^C&-@/DMM_U5I09fMP-b8e,[OVJ._[\Q@DJ51)
5K\]E&KHTERXZ&)T1<K+J_g./&,-2X<agFcF[VT0H)_;91QbL/_&H5[0B8)B#EI?
9b+H4&HR_\14)\S]SYY:VAG)>TdDFK6>f@F0\E;XLZgL\4b>>C#c^=U<(XDcFced
ECae_=^RgORL+&Qgbd2E[FOId9GYOUW-5-.Wg0)d+\abF0XBFgU:<\\1@L/8I.?2
,Z(0?Yd\[2FTGNB=B=)GXd#?f@cb_YJZQNaGcd=]=L5:[LY8^S2&d5QFK/V(N8;6
B@&C0?PNJNaE/E.;:f2C_\ON(4[]1JHfL[6:MYN?,RfL(\/94#Z[cacR<#60_-,W
XFXG2[XE/4?9KT?+:aW-9BJ>B[K<a(X(.@d^5/g:N\++d\R<#[KU-ME7Ga+_:;,d
/:&5g=f>E9b2T3Tg8MBX/NH,5<&E03D+GTN9P..Ld#T#B8_XVgWeALe\V:fOdP)V
gF&?O+)>^74C+3UYO>AD&FQP/UT&]7G[d?0CVI48UgaSY=]9VW]-d<3S56MG.62>
#^6f4VH/&P[Y1AL+BR24@N<+FJ>ICJCW+M:b,-3P3/X5[YR8.K@JM^7b+@af8d]B
cP]+Q_6YWW+T\UUK0:NV8#(CgRP8)\+H@<:^fF,2aLJ&-+M1Y3[^SY<;&eHW=fd]
]U\5Fe[cC@OZf1)NKI,:E#(^)Eef.3P^d>HZ[gd0QW1e@d]R4:/1d#:<<S9>F1aS
[TKd3Y))Qg^BK=2Ib#;<K9HQ.c7>T6W)1SIc2IL\NDJYfH&?dUPDWW@5,b98d.[J
8<-2G>8GT8QJ0DDAI9G(UU)W=2-[Z9RWC7cC9<eEFZ<5e=LaD>>g^49-\5#F\KHb
<.;;(DZB9EdQH6W\##)fbI98dA[3Le]=U<AXL+<Td@Kb:(#EH5D&+-P@g&YF2RNU
EW]-P;XL;PB7ZN9_4A(/BV=<1>FWB[P_])XYZ]1E9>UUFc,GTc3#HGOg(,Q0JDMG
KM(Z3?ZU>L1.39>B3G=FG>]JJbLZaYc?5cE0GW=?<PSHR^>7[.Cc_G6YYf<@,GJ#
e7.;>aD<9<P]BBd.E95WSS#7fA3Y[IMYRBDBXEeaOdf4.f;=I]RBHCMgZP5.WI#K
,SW[U\NMA&]ODM)IN?DKYBCKcJ,&D.-T,?PW]8RA,9TYba==J,9+[eR+5^D2gA:U
KTF;(JPe-JgBA25Z:2^E/<cN=]5\6MLN.BCR:(?I[1&=GMKP5P,6DdYENG)/J9L<
L_:.<M57?:f\K3SF?78Ac06))6Q,;1Z9N\8KV,/Q/I]Rdf[g3Z6[3OUN56VAOV5Q
#GPSGe;>Z00ZNCD8d19,R#\^;+,g8<HL[Y\3VQ[(f)a?#-6Qb9GB=HB+Fcga>,A=
O#NKJ#8,K+/2UU#;5HE6d^S]6,3a&E8b/[BLFee5_F(12E7?2+3()OT#<2A^8QS@
]<8f38C)&(bA&;Cc0V1SAKS@-\&f]--5.CQg0Jc:cZ=1?YPg(<aM+f<.J9=dBc=;
D0N/.XN6);XEUN[0QB0-(73-:>N,P)PCI6?G_&=Y](-D9>3@->&b7B4V+e]^(0e(
,_1<<7[0U)@<PLDE8a6:M6IDee-MgC(Q4Me^M<eT@Ig,?c@(Q2O9SCRX(f_aXFbG
X,8SD\d;Bf\?e]-+#2AYWH1=482b4Re<,8daF>^0,1THg6(J5S^+9N5?9(;ebAdg
Z+LaOY-)-UX4d\2FS9C@X#CaGeP3^fER-(&63WCN3N#8YFa6(I]]AE_aQ36S^G<,
S4&:;X4WfBg9I<?-2S8HB>bWUX#2B[C[=.VG9.Rg[._S6D.R/OEDGF_)c6).IBTa
^R\NLF,SRa?CBY9KZ+#V6_()8M-DZCKf,c@fK1VW7#YGbZ^C[N2_@P]N?[>9\J3:
C(HT(<85WLHWNN.:I67g2LND:XDfb?0NI;[Wf((J,5Mc7<[]X,SI3]dP-;VUfFbD
NTN2)B8bOFMCO>PYLaa7T1]H@GeWWBJd?+22.C=S@8O>:1LVI]Ja==59R#NcF-<B
bcDL^D2)Lg+)7_=53SH(CD&VFRTG0))PM0d-BUdd]W2PI59W9ZR_]&@9?]a+S\JY
JN<S#_;>P2K,69FK+-&UaE7,JF-UW38S/F[++SZ6SHJ-Q9@U&D@KT/?4=Ob>FgJ&
YLW<F\C#R&BP_dge7-KE&\W2249TN+CHD1=S9Ggf##)RBQ+<ZR-+5IeaVS9QM)N-
UD<e-5&M+QS2ZZSa5+M:J[2B+=:2VV0F1E-:Cb5\<YgfAGVU8<-Y#f@PROK))S(G
BJK,Y+MBX]>YB)eQ@]A]_\,\P)ON=5>1\SeRGf2^6cID_R3MK@f</1FD>f+b;=.F
^H-OM&ZUWYC.Icb:GWX;[3P1SC<ARK7V4TS2[,a6bfe6BN5Z_X/M=[0]^^2=@,,-
6JOQM+GF;Z?X0I5:H\\Dc/,>_)a9Z5[6P/A/3SXB::4DLN0Q@T@.?8X9aAGH_[<U
0#<2RB6&T?VW:(QW73Y6:_;^=,9J;6WXbF7a;)_66KYH,U:>:/JMO</5W&1V?c/Z
Td6g-I5)0#M/g[CdeS;V=HWMXCNE2UDI,N13X<>.<,X_1UL^0;[_][c^,U9OOUS/
UV]_#JNTD\D746aO>E>,9GZEO^(,&KQ2PK&7fJ#5CBJCcX[Y1adXaYR5WYd8U,DC
QBc0&?-:PVdT&/87P8bd+OTE3;KRXQC&d/bNII5U2G?^+M5QVO-Y6c0MP,:(MbH8
1S[5D#]eMSge_5_B[4&KI6Z8McB?ZNG>V6Ug0ECQD<c[2;;=S@_VX:9VZTOgN+b4
g:gf^<aHc3[P]_:/Kc/]1\Y_H6?.d74-Q#58#O4F[cXXbN+1,V>=Z/D)8#:)d,B>
BP:Y)Z+#W0ML95QS#YR]L1LDBQV1C1b2.W\&\5XE5=LQ.>@P8dZ4:SEF]Qe1TcQ8
U4];?b-ZK/N46MKE7G?+6d/T./WC;BM31/VAL46/7TW12LRa87M;;A>6cZA-H&b1
K:Q[?/N><;O+LDXKYEXS2c>8M1@:+6O((-X_ZW-1N#T^e+&P;9\8LF=_2TYe?H(9
PKL2PfZ[?Y]e>:b:ZI<0EUC5)@.K.2XTHe68?Y0X8&OPG;e6-e+FDQf;cbJQ(O+-
Y2SOT8)0-9EOGg2Q^0LYWLGE43NXDO/?4c:?ScVF1f,#FPAC/d#138<^J7Ec#Na5
Pc=;\,?1A(d=C7C2Zf/F&&46+3@-[++G,1>[G)fbKgGCDeMAXKQ:g06^7XV.\+KB
)X+NaP?F1Mc9(B5P]EP8ST,:K65[J_NTQ4LD_06T8EfN_YYS]>VW>B:Tc^./V[XC
57c=g(C=+G5:U+V_#:W1_FKARAbB^^/\8AbaYLR4.<Wfc6]U1Q@+-095F:.,1^>e
&KD/P8C<?[U&H96)XPPL)BP]UFT::=(#)/C\O340,3&Y9(5S\YORFIR1D\^0C=_=
eR2P\3ZBKM#RTaEf#3KRBGL6.VUF@NGO<KQ4CWDYg+Y0R-=1(a<A_VfUIL<^^@Gg
;\L5;R&OZZ]FdJc;WBCV8690dV=[H=][BY:];R)+66LU/75cRdb4U>MB^:1bBG_.
=-RIO/-U>?7Uf7FM>^=_TF&^@J)Wg.Rc>+S;UON]ZRf+O/HW<+NODMb==GA#+c+1
CUYTbd7>;6DJK,a?_HJ-K=E@W@?RHQZN#X[-T#G<gCQ16MBe-4b39A#KdPgZ?RF2
@[SVCKE8V(?59.fDJR+XS/6\1,4,.L/[7#]4E#A&DT)XT+]Z81&8:Ab,R&J<G\U#
Y)[-&YQ3[;7-60BTZB09\B28J-BcTcbc#KT>T8,?FNNNeF/T=ZI?_9QXDa)@J(VH
+&bTAdgcFUXVZ1X>dTPcI##7L2XQYdc?FP5e/f=e=4@X@>a2/?];?D_Qd#KPLPE[
Qd_OOeA:A3ZK[;_bZIU<7<8^E]?_aCE6B;gV#KI3cCH6:LK,Dg(F[WZXK<1QYB-1
.e1&O94,91-?\A(Rd[,7445c2T@:#f03XAbC8RS2)ZU,A=.;>PH@9&Sc]B-6E608
GPR5MXN-/QdGCVVHGM>^F5YKPJSN+9YNQE:4;HGEXVH6GdfPYM:W&eaZ=3[A,^/J
TSbGB4^&8C<__?TPHU?]Y1P^+7Ga0T.eA+,40gef]1ecQV1L+Z<BRg.=C>7/88>C
e36\]/>S,bQ06Oc8c5^L/\AO78H4fDX-CO4\-J-/ZORFQPdG#Y&c(>B?.D[:gK1_
5F,cOc(#K9@1Q]EO^EG&dQ36)CbBSA#=N;>EN),)\29,c0R5S6&?NWI2TOI=6?]Z
T_/f:@1=O^_^X??;JJS,NOPfHBEQ)8?)91=QYAb#^Ae-X4WWeFba\+^ZKg=K;>eG
=J6<WA).VT:LNJ^F?:=UX6BI3fKXEGB&Q&>G7>BL^HL=Z&&G(#(G&\T/S>T_.e/N
:#+C4b+KX(CJL-0BTM,?gKJP\&+VP7LReJ6,MAB6],QVIPR,8C\.&GTe8T,<ICE?
X<-G-8>18;[a]DFgD<B4((/:L,)+M08,VFI=O>R<K75H3L2P336(M-227aOd.,-L
\S<GMEJ@TXe82de+&c.J1d6F^f69^VD<#L[+-9<<:CX[_&K-8K^gb[;U#?LWNXMZ
^gPdVc4T07;-V;Af2+eN[3]JHX9=0YF)JD2c_4]5MVd8QK:GXd&K&26F)b^W]XA6
D_HI4S3M=<:I^aAcC-dUIfRW=^^[+YT\]1T-[b1<[B5Vg@:,,fKVJMa=],/cZb(<
U,CMO-(;:?XG^e7(QK_=9&FO,f-J2-1VLA)T<>PZTLD0G4P^IE\MC5UBB<H3ILSQ
dS)VBI[@VH=bf&1U5S<e/62T2WP0L[R.(CBHI=:&G9eK=J^F>9SJ,CHCeK?67c##
U0^;^W#;gV(L/L:,W5=YO\T)g61F?33(?dB_S5S0d02M4NT0aCd]XV)M.g1D6S+T
9WN-Hd?b4UT5L7)F4aH(6(2>AQJ;_4O^DTK7)[\Ze5S>AYMP\@2M-6TH(Y_2]-d_
JIXBTaI#e-I&5,Q,:13/N1N0ceTfJAgf30QKXF\U7bB^XMe=c>=693UU:fF3<5M&
V[fERg=@YBF0GC1>=Y&S2([.;>eB9<DPA:+D5>TE62b(UIFO>fPQ<;KL<I.O/DfL
<R)>5A(^Z:<^@#_3^.+bEdFVE/L9cg)UEZd,\-?>bS<G.9g2YV9U9&V/)(D:0\[L
Y#4[S8(g/T=L7N\;D8U<eBL[f7Q#]QI<8gd;;^3M0d,F/H)?5cgdIM,3ecQMP1[;
VEdD]YLeH=4H7]f3L<7eJ-:Z01a8G>+G:\1@U47ZIYba&T/WVC.NNRV)(O5eQNLM
0GcLEbUI5BJLDY5IQd^@ZX_1MLW]Z?LTa>KbFQ3dQLA--9DS[TBTDH5,1gZ2;Q)I
C:bRf7FLXcf)-VCN>I,JJ?e6C_/UA2)b;Ld^/YPXR=18(<P5(7dJ1K[18HA,W-NL
gdCUX+[cF_=dabLAd2f>P7-c#EJ)<Q_H9V,..fd56c5,W\W?ETc,7EIK>:\<L,MS
JUfQK1PJ[=A8>+XSL[c:=+Me[MgF1GXPUQ@\+cFJQgT,A,UKQI(YML^,>]V9FZ2R
WEUL3N1X^N1b=&.PT+E_R0\PG+XG0B^F<S)J)g7CNg4Y&e7L-WaFFdH7U5\[0;Ug
Q\#M(+Z5QIbZPc-FMD59#D-_g)\M?[5KDVZ)=]1Y6^LO1YN:T-QfHd&VM48N-)-L
K]MMSf<Me@9W0eQFb<Y(D>)+A,Eaf:RX)1NX@7Be\KET]G),_/9a2CY59VD7E@-1
74=1-L2D^aW.M#<1FNCe,OYbY36-8L28K487Ta(0#Mg0FO0\A;#c-YI-G-ST>>Q/
FY1>gAB=TH@U725TNYag@Db_T:Q=^TAK+B/bY?-,Zd3#gCKdQ<P,K>?G-a<U+Q[>
.VA?]0H&58LX1D:SK/-706<]^F/:^.5/U\D@Q:dc#IA:ZHEGHL\N38_4IXA9?Pa0
>\gf[NO>^9HA_RO4?QE[18-#dffVg_Z.CK\#.J5B0Nb0:6>+.Tbf2TZ?,]\M@6:U
+FP+(.4gC]893eVE&1FGdY<XfaY.@[]S7E:Ef8H13e/UH8e7LJTEIWQ<S<e5aQ7X
EN@](&MSKeaVM?0_9]Q/b];aSOO+S_M/QdeGdDL&_<T<T>1UadGQbN7+K3=eF[HL
5P;\g_:aC=CS6QO8X8R1_LWKFL-]4;QHD-b@#NCdT#-G#ZNQ1YX-OG0MAfA9V&U[
(0a#2O:,(bJG/..F)EQJd)Ggb8EAf0_CMcUg==1cafcO_c_D;U[KJ^4W,/,bILRK
CZ_;<c,.@+3McB6^[)YIK8F2+RJ9J)@>8-;(HYLO.TZ,6/cITG7fQ0df-RQ;T/GQ
R1]/?-aWFBNBAL/H06f;Y[7UW(\e[8N=I;\3^6Ib<AUY:HAXU._5<5Q)GGe]L2#\
DAfG^,aT1(?,Od-@NSbS@\9-QTd/)Q#fR7J)719\P1a>([T@((dII>IQ_.C-XGb[
B:_4UP<^cHI<6X:KP/bDO1cR>ga]Y\OVL61d]>,E;P26V0)&RC(^_C6M41]fZCc3
VdJ&81=KS\,N=gRB#YJJXEWS0gLeZ]:^^D_I/7d)9O4T\36WbGPa\FcRZ#A05_&:
L8N]3[6cL^-gZ->)ZQKR:5K,agQHb635ZQeHO72R_C-6-W&#BV-K2.[GE,F>LM?(
\c:1[\(U@4-9[0SMa?^e&\f1PEP=]eQV:=YePa#7f+9J)&GDS?ad,)4fYFNfT;.8
.=C6:UNBJJbfU9PVN_dd_6.>,RGfEL_?NOPP[SNJVM6F^QK\U>HZMBRG<a.efKXT
Y^e_\8F:LM2JdZ@YT2,8:)gReY3,(dILd)g)2C57S+fF:I1A4RL0]H891Q5AO=Z6
B3/O?Jb0/;X\3QUU@Qc.>X8f:4C(?,.P[O8([9#<;PL7KU1bUb;=_C5eW/,?(>eM
gR^1088Oe,N[?Mf8GI-B4JBbCO7,aL1.&1FKcX)OA\b7,FE@J4DCX5Zc4+6_f;d(
-][9(Y4,5A#V.Y&TG>AZ05WKMI4B@V:8b+IT)_geY(I&V5#S/.F/0>af^GC-Q[)P
0)9<LY/Ra3I(]<.<D#c)XcFI204HA5-3E>HRB2O9)+8bC3J\SKeg/8[Qc6SC5?W.
XM>9RG]5K;?5ggO^\Fd>6?X4Wc@]9U-QU>TT95<]QcXI,VT1&][C2V\[])J6IJf7
+14[/16Xb2-@WZe<JLPNZOVc5^cB<XHJ.VT[R+:SH?J>J9d)78U5]R1;fcf#_2.7
^?5,5]gH+S/c4).J=1\N@RYQT4-RNQ7.d+C-V,9fTG805B8IHf&Q_[13L7db;4#P
8Q;1P3VTg\L5AH/NR6.b4-,HNE[C6-Q2#McE4>Zg(-AJ&AX,Q=?2H,Tf^GX8a=cN
BPG2L0,TE<dcEX>:)bT>C8TZL.:3(c;QNDC)[&L^FA)\I_\3>d+\+ZW.Ha7bI:ZP
8LX-1/Z@#;#1UQ74a<0\,fCX76A418EN-#;P&C/EW(bd#375=BCN-ZC^f,;YE0(H
CX7aAETd&NM-Gea<D#9d>,V,@<4E(&&GFbX50-+b:JfIH0BG8GT8I&=.d/I>9U1:
J8:^5U8H_6Dg2K&1-+-Y20[.B@Y)S-T1c86KZO>;3IKN^b8>IQIcf8?O=;&JZ^QB
](TZ70bGR+?]<C0TVHf7#_Y/\)R7:U>9+R=KJD\dPS.RZT9KO+gWVEQHCQ<ZWNPM
KVH=RD@-=8HHDX7(eFFDc?-\PfW4JI&BXCH[XDS)?/VZbf&]KN&ZEP^2gQ>9SKL-
&18aJF3If<U9,=QH7D.4.8;9<Nf6>FB.52N9PGTa-HFQYN-7.OV8(CV+Kc>U=c)M
,Qf#ROSKADbOLeW[99>]fJS(aO2Y&HM],F6\4F0:>4;9c+;#?J#+H^&.;R8W[fY[
.=.L-e_N-Z)dL^F4QbRL<-K\T(IL?.R.19G6?(VBE?=U/0J;<=^>W7:>#JYSSeeY
)IN/U,F?=]0]-e7S]8&#L(.F_MSDEEZT5bV>^VGE1A>#+:aK,L[X4HbWNacT_X>f
,TYbVAg5OR-IC3G=eZ??,,#5[2d47&+,U2M>+(FBge\f-\YGSgCOBQS)aD)1G(XE
+BDD6=?2DX\N2=FRO=3Re@+aFTeDJ=@:.6Cf^.]#)ESMGe4^?aDQ3N6gc^TQe@71
^ZH_QCSRa8UY8]).033TE>,)W<7N=<W/8,TFS<7LX-134-_19G&BQ8#d?7O@IUWR
K2e6X8>;K@BWHJ>042)<TEGU3<W=GLfUZ#3N/4+\4LaI#eYE^]?>1Rf0e=T^c-9Q
J)Te>4IfBW1+J>E&Adb^-59gW.R,+4H<A)2&@aF(BNWX5Cb@-8=1QWbL<ASB[Y7)
P@><3(D<,9E>Ld2?9,aDc9&7)T_C37Z#EB(e)bR,]5fO53OR@&+W[]9gZ0d,.+N-
=8],a5@LDgbfI+QVU.^S)eSN2TS\&@@]M?#;#DfGDF^\M(W1EL0LUe200CFRBUJQ
TK45P.II/<5-Aa2A3eMFLS2-T@#[,)?L#2-8EQ9KQPO,,EEA06,c=JKW?IX2WETK
W68\N.0_RGD6Z=6><]_BX,/E_49;V#G[0-WJUH@\MI#.7?FKb/I)J4?CO&08AS93
FDJ;B<?82)6IA.2Aa8[(H47:B3:LDE_gg<D:?3f@T12H3DL;K\5TFA-Uc]2?QR^a
dZ#)CIZ_OU,@P1ba,\7N>;JF;)NFTb^@,72cWeP,9]d<\LW5a11O3Y-P1HZDaR;X
UKO)&H_g1S.&M<?bS89TGCKOJG]Q4Of6POZ[K.V87S5MZFKVGVI;A9.gcW8f?8,Z
=](b-E>g?3[c9g\#1F]S3Ec08/G0[CXNCDBL,U88UNI[V(e.3,:gEA9PRdBQ:2LK
K3[XJ/,/WZ,6?A_[<#0OeP,7?D.a56fL.\12..0,T<>#?X4.E[(ZP4(>J>-CP4/L
;_UPC;/0Ya9]6HM/RM[22J0;&C]B>FQZA)9Fe_=a>?6)+f,^g7@_JY-bTPDb8D_d
L,_&@A:3;/&K12b]S<8M^\/G4@NO\gMFTII9g+?<(T?8N^\BcJ[c#S@=]?KeHgQ8
R\=M6]7dLcg1?5R(UD7.g+Ie451ND(QTZ]#^;(6<:bA-TNf<OD33H@?1M[aaF@UA
TOC<NbP?2D@HSMGXfg.E?(IONGcR_80&W]2R<De^P2<HE/KZfE&)dMad?ACAQJ<&
H6bFNd[?D=_GFOG;?dL_E6C23gS\#8bN]Y/(;.Lf-X<-gQbbZF;FT2CDa58-6[M]
4b/L8b^gZ]&aU-MH-_;IXL]#78@]#U3L,g31R1ZfLE@5dTB=e#IJHRWMf#/1a0JW
_DI2HNX17-F^):3J87R5C15gLB3Df-#/1<K^_)1FefC-GI4)N0XGVQAESgfg,OO_
UJL#,2:;FQ&F?]2ROLAg]?N)La)/cGefc.>aFP+.E0Me4Qe@^NFGTLE##HAE>2.T
X.^ZML2Q7--\f,DBR3D.(7@Be4\TGHPHff&7IRKZ?Y:Q+?ULC(YfHaPfaOAIW4KX
_==#@NdeE3M0,#?#060.;;@JBgUHcW.Q\(P&1V&ee49<@d-CW.Q/f5>E1IaR2;,9
[GeI(0;]:?3QCQ@E<C^)U804[ADUgOK;)S0Oe4;U.PgJBSd&OE9-RGc_AK<cMGb6
Gd2@?4Y9cVZ=W>GWRc>A#a__cGIH#MdA61U\VYL?6>(-.Wf59CJ-c4E0K.F:#RDg
2T8WX4M^aRBbccEBWb(H5@gKWA-_;\,&4[^McRfSL<L)-^3B]K.Z1HJJ+FG7TU4b
6[Zd3&#YfVAZ=A]A=LGM(,=Ad7<eW<JZaKEe=5-U8Z:/RWe-ZFC)gFDBI(V)/=>E
;BAYCYc__fBN.9\9J&a3QeZ^6@cK6_#^f]6H)3bNIO5]NKDR+518QbS&&88T4b-:
RU-XXOfW<I;B(1dX5BcG80;M;62R1ZVdW[V^K)-DS=Z;742,QJL][a8:MdeI<Q1=
1M0[Q2/DA.R1EB6;Z[Z9:&8:4\MQa:N^eO>(Be\e+:f.B_<]^.<WG?,49V7KR<]b
W_(6U/OXP2CP;]KO1^&?e&Eb:b_^4I1(^8]@\NTX-R^LX4CQ94SA2Q,8/:TMeTI5
1N?IGff331]ZG+(\;MM=Y,ZO;8<-US.=OSB^cT8\H2-8^C;\-(]DVS/8)LbQC#<3
Sc?7;STIAD30U2KdS9<.7+>I:FORX;:KeK;J1f4AKTUbF[>\Fe]Nf1c^>.JdIN4T
@SXbdZIWBMO/]13dZO9VM.SKELYb>K:+WFICd0&J6)NU09@J^M-WM6YCHB3/]PfW
GNM_RNCP0+F&e:\@bdc_>Z&/0C(>eV^.M91_274(G@)XSJ598.4UE_Z;7e3,B@:5
7X5>?RM>EF&<d&DfWdcYa<3T]2[XGUCD;A\-gb)@+<d5N:g_EKDHD8PQK(2e+&0e
aPfgUS.U#A^7^TU=_bZ4VZEFN;7/Ie8F5VeCLA1OG>&=0W\9OKf+O5U_Y0eSN@<9
#;(KG)4OL2Cb>HT/QL(>N;7a#U,GJbJS9a9>/E?]N];3bFUC;30BEaG8aP:_#E)/
Q,RNP]L(8#P.:BM4faLBC<#REEaPBaH.:DF9(G(W1(b+gVWE+(LXMS,D2[O/SZ]Q
@bB]R)Pg<e;#Ja<c60([>DB^>[H.gPKDXG8F821aV;8HTCDG\)L<AG[]9Dc6I>bI
HU5>:4+GF5PJBF\3,,OgE(EX:]+D#B@S4_V.Z)C/.1^]ca[Oe55#9Y&5-]N8Q.6F
eEXJMd:d:4G5UARNf9])J?2gBASgPP-#IE:A9T0>c2B2)Ab((cL6gRDa)3R.D+Pd
_47P[EU@JQ&E;_U&O2eVf?CbCH_Wb].d[]-?Qg4)5,F#IM(U4Wf\MJOc0Q@+/1;Q
&QJCOg@JIVf2VEU(TH)@J.27,2#>\N@STNR,AP1_2KA21,OcVF:H^J9B?\L>=&;G
.K(/T(V.,4/[,Ve1U9/@S;E4YdZSc3L.a4#3W0c(ga9R)YS?RT7869=H:S2->>1Y
W1YU14OUPXD\OAUH=JeRf3F+9Z2JD&XO_,e]G4EEJ]R9QV^U5Y<I\a?7QFRT.Y+D
>_aOY:eVTK9eb2RCKSH#T:gQ(2#=VeFKW&-LX\F6(bXf,&B4(T.PBK2VgA6EbgQ7
)A8#Sa,?BKI=JM8cKRgTe\J]<g@C4ZFe_M9G+fSKAA4+V,)D[]R@fbJSKJ#ER4_;
g1[EVe84fX:JWbXFGfbG&M>AGUEc(&A)gN\16_JLYWWC/8U3QQ4@WB2=U+AJ?b/+
/cZHad0e+QY4ND5[>bXM?D^7g,Q#UE4b(G@2MUZNdA9d^K_]c9(U&VWeDLMKTUAI
0&DH.U^6Z9P,\VH6:6Kca<<GU_UU#GE?2,4A5TZg:QQd<2ga@TA;-ADI.0UWAKLg
_2B2FF@LH)DU.QC^<+d6g>X>EEdJ26.X826@SNdB2cag<gg6+/N99O:Z^fVZ-9c0
WdZJ2C9Z@5;=@VD=B^3FLXYAggFG\O9.CZ(8.Ra4IbA=fWE8f?P=bgOLc-#K[PI7
&;@5R2P+cR5LgDYW^O^?G+eNHZ3X2)T>]EeFgE3Ug#U;CS4?LX<P8\:aD7W\B3&B
:8>:<-.-8DGRS6M;1RRU5)9Z2_eUG;0deDD_04d7dXc,=?95a--ESBd+]ZOa\c^M
?4U@NY?05_)82>Z_.gaY)8U(E\Q@b,NcA8e@#NE,>34/Ag#Lf6)&(G+9FCH=W5K,
7@WcSfJA>T:I>T8=@3g&Z#S>Q\Be>CN9/0>eD?0-F#[8EX7.M3](MCUPRVH<AIc^
UV9HL+Rc18e(6_-WAEKfc0#&FaK/=VZA3DcMXQ#UFeE3>FU@-5V,g5I+&S^bUTE^
UZD)-\0,+=;W]M>G.=DR+LQ8?:LMA[HN,^NfgZ/C7E7c(fb:+_4g?ATDAY[c]/1a
>DP61P7GK+;RVaO@feFU=G\STb^5C4)J]-QAL.NWeNeM<CT.C,_[2(HQ32gTeZO#
6BK#SL+,e[((QM9-F\\X+8>SNOK[GbdMUPKFQ?2a;C_XE&,-dBK#1T+XOZO\8U(.
=M+JN=T1c.V]&D:aT\PJaGLLa1M&;-,/I<TO26a=e7CA4DaG>I93[URUd+M36;5<
6I]]Qc8_4IF36D3A<DDc72T<[+^GJKX@U8:G]g&27]>-\Ce?++S+UdF38ZO5\U9b
T;><W9L2UD0O4J:Y.MLdHVMX6S:-AAb[G0.,f[-0GB7d(<:T7?QEaSZPW=D/G/OE
X@8-dg484N7(Y+Tb>81+-O.c_/ZT4bJ843HRM+-9K47?4dT[O+#[#E+LR(\B\gQ[
]a50^9R+VOP9eW,=FJA:YBL<[<&#NE)EV47ZC;_@gED;>>Z5W)g[U]LQbBa6C1U5
TGIJef?S2E=I6YgU;(#,(4JS/E>C-=3UIB&R_0HC0DfQ#>VN(\T1WTUCP4<W)9_2
XAAd&89=UAYQ]3)GJ[E>+Xa(CPI83H?@1IBEY@>-8PRb2cAIC33(.S3K2]6a_7:C
0cP2+@OKGKOcN^D??:?K^D<:4B:Z<>AY,0dP\T&)g1?MYG8.bCG4;GUPc+[JTS,d
6.efJ4A96J]#2/&O#cP^L3THO[KXI(X4a4@3WJ?Pa7cR#U.PX(2O)C3B.NT1b/UY
C>&>b<)e2g&]JC8@4S1WCa)7W,&7@&9We1b&>CST):<.BIK]f?]I0_Gc=aQ)ABR-
4^2;:<LD1P=OAX1=[#@BBRG\2R+4EOP\W37@^^4e;IH+O=3B&V,aD?8#;;&c2aWZ
9/)+@YAF]1#FDaOUB)#(Gb93GLB-K-7EQ7XJ+[_-W.OIS##J_+7^+G@6REfOERbM
K+7WCCL7[,@HJP?(H0BJ(G_FG.&;X)3G.f.,@4MP#GPCE^G=Q4bbRfI6]0a\WEf#
7#@JX3WV)&Td<E#7d?E5g^;8VdDT]CP8AB]NBZ1JBe-\9-f(E_+G3G]O./7W:W3A
KgU#1g/aRO1KVYX86eW(.\PY2b;M49-/-HM^42P>87c<BAfaa?Xfce]OP$
`endprotected


//vcs_lic_vip_protect
  `protected
,O79SJ2DUb80J0M+WZZGG6PAUD\]M?Z/a>B:V]NF6ea??DT#a4Lf+(G7?39&2SFR
B6XcZ_b^A]e9HDRC@G60(X;_4;D?F,e2cBbV(&/Fd5ZQ^-cE2KaZEbNfR7^W?LOE
#S/0BY_S0I3=4R#RI[ZO.W@>/,58.g(cOf9d<74Y3IKKI_U&QfC-XaWCcM:dcgQa
.)agC\6;aU&cI[S6&E9N>d\cfL\U@GMSG\f27Q=2(?]L:4BGTED/GF4O>FX-Y\1O
A/F4?&8^.33]=cNf6TE]Q9-S7RZI:0]C;.B+d,I.9,(ASRM+d_-C_5TJAMd(-DE/
>=S=fZ)KI5T>Y2A4SY0Y(HI#1TPOYO6K,OX.O#^4T^c;GeX=Ebd1I>I#1&QIT^3R
OIV&,d,PPUc5U1_PCW,H0;VC1>RfEWKOI9ID.T1b9XHG00-?EPL0g=egR#D+B&Ae
LES7=;]YHKa0[BS;#DW>2WV8L+DW1EaDF+<5\K@Ye+fRa0d^.5R.3=8#AN-(SCJa
:1aCc7EB1<R;FdT<[FCg8RW7JE/0G,W^34O]@56G^2f-,AIf&XWYC\>e4E7,_L(I
8TZ,(MU3a=ND<9U<F?ZKLSCbCM>9-<179B&<<cYa?QAXQ/(XQ[;YQ5GHYO.RSEK5
U;2/eZZE#_Q39CR;<J4L2JeLP6G3-JA,[d)-PNbZ0DW,d4)L+9X0,WFLNR?/H5W8
_Ef:23&G-;E=FZL,?U3g4=6V@/M/5V)3(I/K_22Q4[c/ME,fc?U<6ba:aA-A/ga/
:H6TVH\:)&#-[L>LC+c)?d#F9):a?ccUNMZb4V5EB9ac=Y-?]9&#gf[;G.+;U]M&
_9VOc>F^H^<gK\Mf8YGDg3\c8I:CIdJXa-&1P9S:O-:MM.G:_P@P-3)&J-5]]b_T
eR\YU&4O5a,ON+^1Z.27Lg=H2HSBR&_YO<=>WXT).4[d.-O(^>C\26W6gg5\/RDP
RD=c+[BVIfZ0e-__7=\^O\?_ANA;J)3=F1,I0GF;2((Yb?dBQHYZG9PCT790/F<9
TdDD@KBe@\-XKFNL:MZYU;gZd)cQ1_fLFRg#T4]H;OVVW2,dIU_;cEfMQ4g(bc[X
J8]9W9J;.aH7Y_<1F60P_f@4:LY.+:,La&[f@M1SE@P8/cA_TgGeRTSX3:K<T8f,
LR33OU-7R@N=@/ZX[N<9Ia=D?GFF0eV7SO1d=X.f>-fQB/XE>d@2>KT4Z82+a./3
fW&83-<X:GLZJ\g/BaUI#97-d,R0[\a_P/,V_SCB3-52:XMUNP^.,bQ=N>@c9AKg
F7:ST0OMa2W2,TF?F=ceQ1M;6+QO4:f3]f&>XBOJW<gMa&OacVQ.+I#&HJ<2R4X6
f/Z47<,:BZE>dP6O#8BG:Dd6LJG25<O[ROd\H4BWKVL\Z:1/=#BJGa6G(OT<PBUe
NL,dZNe@H]3M#6P(fDFa#:54M6]A=D/([/;+VaO6aG+?.>;R-AfB]G^DX64TP3:9
d2Z()bKQ^ZeDdGF-9DgNYT6OH-;ACe>QAFJg0SBG-Y0bBfC7&(fee5P+:ZbCMW:8
+3N(G@)\-MSE]S[?HBR/fgTa;_GIA>MIOXNJ539[:).#F]IB&B=Se_),?IO@FBKU
JeW^ZU2;Q&Z.A5Q<4@/dS)PZ0d=B))E4?40.[fCHST;dHU4/fWeAg7bHB51ATZb?
BUZBY<8^2QbL13Z(MG6M,M6:2EL0H[D#6JfR:O25c_3aH5HaHacVbHO1e^-PbCb/
9,g.?_gQ<e[Z4b]@5ENSgPWR.eLX&A]e7??_eI<9+/c]9B^Y_2bdGLc3[LL-OS^E
M8P#fKd>/ZFI\]GK1M/A@:V3C)JNd1b\HS>_]WTP.TV3H>O;BdPW4[Ke4(.X-MdR
K^ODQDPMN]HL?V25Df\PZBNYS>KJCSG?G9;OBVC1RVf9-g6c,+eJTa;G^Y8[N^]#
gBf_0;ec&W^3,WI9e@CM#PE6W)GS<B\D<VLPB>\b2_TM#K08f^W1];+eO79OTPA+
0RTO?MbUEDCR9:fK_N7#]H-Fea0OZ[+g+W[dRbScg8/10IQ8-Dd6D:<2KfG[Kf[1
S#0ZJ.?U:]VHZEPIKeP/EJJ&(,N+)BXR0(dJ]Ud,,GbbY],bUN(f;N6b_ADGD6/A
@?V8YAK3H#XI+aYTWKQ:J>6K45\NP_b^J\7+)ZXVB&0Q<g0b)?A<^c^gQ(fV/F-M
S[eH,(K<geUcfa[.RED6=_3=189BDRJ>/4:[>a>/VV>0KC9\I5Y7AO^H14/fU1,C
@SbZIY7O)Y\YK7<8fIZg-XG\OKGOU6I(Q8S,/W0SEK)]_[/_5e2G_f5/a2H(#R9#
FMd;aUF5c=+2U4,D:[LBU]5g--JD<Qgg?af,JLPFLI1,b.HT)0LX<S/SM;^<\DO;
P<@<I;2]6AP9fTc^?\>SSH92V3Za.VX(9Bbca:T92=b/QC.LQ5\K[O0-[9gN+a2f
F;Xb:=D-YLH4@daRCM]O._BUTA-,dgac=8>9@f0Z/3SHO(2X3C47\e[KMSE#,Q)4
Ab>FB0J1<FXAc;G=^(=WI0O9652;\\5X75-UdBKO>7(3&JaNK3)::N:7ReBbP1Y,
LQP,WT&675NX,>W]46_\RWV>:LP3^Ke7ZG3OIg5_T68;+_)0MP-6C[)+#H7e+ZfH
=9eS0LT#X;eHWa\Z5>b\<(\7G;7W6G)93]=Sffe&1aZAUJ7fdR,HFMT7A7/ON/A)
[(JH,&FCR6c8We-L;&I/VQG+7I3P\9FJ=^W:J32ZD@[f7H6JXUKP48ALb_Fb7UU1
B4LPCZ)QXW27CV_HEE]+7BX()^Ab[9bE.AKL1:[Ef)</ZV9(VaNIBGS,]?dKG]^S
OYLC.@ZY_U^;e;^AAP\2)3-L+=Gf:)BD4-0cN+]^3;#.;#[P<Igb[We3,MW@R?[?
7A]51U+;IZJZ]D?QY<6SY=^8PH_aS=Q9:@Q+X:J>dDV:+CG:ST:HF&IG;b?:@XYQ
MIF.cL19.#f63=UV?7JaT/IY@JX]7K+WPNPET.D<e9L:;9SRdcG;KCP>D>I7[Y.A
c1Y^X@[N9\3O5I+5\/)e?Xg=#DT;6:X-;T1ZZ_=&e_,+UG4IL4AaMge9LV-U2Tdd
6W<,W+FK7Oc3D>RIR]+#JOGU9B?-O.E1-1BbO@c5?&?L&1?@A7T>D6ZL)KVR/JTN
XFM,MCJW,C3>G#X=2^QR^&BPBH<;8X9;)>b_8d4fVZ;(;IPV-H5?<R_UDB11R4bX
ADYGLQ;FBQ=3GZ?KT-Dg+IOe4=c)9(70OgUQ+VQeMf\X=U:Z_OYY3g[Vf_RY2c4a
7QAS4A<I;_RX=[:F;0:Kc>Bb/7@WfTC^aJK^L+)#cd2WZ>MITD@b^2Fc(fX8-/+Q
JP(Ye^390,F7W\Z5:54B3TM^NQG(8M6TY5,HO+a628,+1S.HL+AJ3<Q=?&(dG@R9
P)f;DJ,MBWH>BJX==+#3YDVLNB(6S+.gK<4/2>O5Y9cDGL.BJbK=^W?cEM2JI5\?
IBDU<??F@N8TAF1E@c[<8\e@Hb<2-]Hg),fD^N^#Nc(];,P#Gd;HO5f:ZTO,BWNN
E)YX,).2V1e-e/.CQ.RD]E:RO:b^A(AK44QBA)c7a-f6:N\1^W6dC(:FOQM1dRaK
PSE>\AaJ^Y5O:D5I,\JEJ]7-LV82_3:<9@+R[5RQ_G\N^\aINWd2++(UBE1P2bPB
Z@[PRV@)S[L;#&H6^_)Z&(VL_fC;^3;FYKDgZ>/;R3[L;Y41K4ERR?SY0)N7,[=\
Aa++B1,(,>5Bg;T]6\#\6^f1(1J[Pg&d_9D5:eRL>?MIZ/5[WV^/A__E=-+_\&f?
BaQ:6gC5](+_&RGM5H0Y5?D.aA(da+:6<JP.G9Z\aC4U8gZJN01RPC<(H#.M<^:-
9TW=DCJGPQUeB1Z14C869b&<bFQL8JN0.JUJ&EaV_T<P=O6E1[HTXBO:-Tbf[8V+
AHV<H3SD@#OH@Q?WG>:ROCN+10Q8PGY/4+(b,,WP7f,DN-L::/Q<K&Q=J\KKW+T9
3b&0D/U1RLSE((S(GO5DO/48+OKeZ@=GIcQXFRAH+U6fPbZ&R6>[d]NVD?[11+GX
b[HP<b,f-QgaWE/F@2>+=C]Y+I=Z>1aB.A2b<<@FG<T,DdXLLFG>IKL59GD6+g1A
Wg1@V=N+@7.<d0e7YL(Ie1d9+ZTSV2-LG5(Td\FV7VfN)G&^I)V+]6&\&a(4:ZeA
#86bE]OXgX8?VE/53.Hf5e<1MN>2Y8gE5ae9M7PJU-U=fQZYaa)9VbF<Q_V[MeYB
0D2#Q]4bJYcYdAOQ@cP)[U9P]bWA\7L(f;S(UDJ<?/=XB0d(X(\.VZ]Z4EZdUH-d
M2VC>4AJ:D(JI.:VTYZN7YSEgE7VA7Ha1/M0BT[/L2-Dg>@b?aWdGA)N,#5[?C<)
7DR;Ud/A-.)_G6[AfI:GZ\HCf?@SfZT6[-;68#Qd2V8K51.@5WCH,[g?RJ=TAT0f
[^YHH@7)(;902)B8#VY>ULG=aCK5CKF05<eED(7PBK7BHV>E13+))YgD9@VZ@MT)
eYVRR5;3HNf4;M\-DX<B=-d91#XP0]JK-KD4P[M01&fgL,IM@6eEDE&6dPG[H0FO
4_f-_?7cDS1+__\UQceRRQ>YdZGLQ7@V0LG:Ofa42,V;Y(S>77McNd]1M-HZ2.c\
WcBEfG[ObC+I8\<\LNJT&4CN8I?<OQ=dbW&R3&7?9Y[J;X-G;+,G\,3N?#??Q_YH
.]KJ8)ZYYdbAQYXUO=:R]EW5:/\O27ef[>8N\Q:6JCL4JB\,P6aM9T:D]1NdDF-?
Q-;<c9+4ad7Ob>D2:NNLV8[Y(.Z;H7b+=8-]U@?Fc#<\58\FFU4aM>9^G?K4:A,H
]Bc@TOO,eb9dOH\B[A9OgPKTgX(,N9Rc_Q(X(fb_;Xd7:JHg>+T_,0FA4/cSIBHR
1J]OEfGOa<@YJ7f/\eN+GQ+a2F7Y9DP\_Q?H4\7NP2[1a^=f[-dN1O4-68aRVTXE
cSFH>P9?V;R3R_31M9FG((0D_ZQ_PF[RX4AH/?Eb9cg)2c2&f(.TPQMbbVC[&QL>
F:9LdK8?KV.;8DKgL+4/PV[L77N))PO_ZOdMbWJcK)Z#^>cJ94^/K=dPM<ZN8]aD
G<PC;7/G3LP&677Y+0#/.>NB/R7JQ]+>UQ_U_]B---B+E:ML.<@N/,0>GgcLG)U6
&O[RgX98V+^@fDK,BgJ<&0-J)39;_)#:SV92#IT_Vc]>KeS&Z?<f]5K[6@,_SBW6
TKN:P;c[<&cH689[N_4LdL5,.U;F#5>7IF?gc,+KEf\?6CQfScTGd<#MU;Z#Z1N8
0,E;^_ESFe?eC7]bNbHYB&P3ST_S0A3V0e:@<@/KDQI^[5LFL)#Oa>O^@Jd(B(I<
#7]\M.-QD88P8(XA1KcAX??:@-YWV6(4,;0QAgfRQeVJ0W28[7CRbWNa=41Q8+?a
9bDL+#)V@XaS&O-JcS>OFX#Xb205FLPM-QeM9fYg:6GTE1#JGf=(SQ7EdT\R;E[Y
)_D5:,QBSVGZ1baeF48E;I0Z:G^3UEb>E7MVL@VG:MQMZ=(<-T.Z?O>5-==d)T]_
.1_Qf[1dS=JX7S5#)g0:eTIEc?-9PSDS,(M01WRMG+7I_P+R6L7&S7,QR=OPA4RM
:)_.K+d1d(9/+1.RfS:.\XSR/1Pd_fVEaKZf>QO_(c8ULN)ge#f0+>:DbP0Fe8^I
VQ0a[X9F77LF_b^R(R)1RAdBCfBVB\.CG_OcK0<=F9+<3Z1Gf1YZ2OOAAFQb?e#?
X-_]^O9S2^J8dN\@a_c;\;_f7(IE=\V>#L+RGHH8]__3B:E:f=-U9GLb[W\H+gHb
G;N=W69@gNg,:;fI/\UfZRT-3(DdX/3.>#BdC-S]FI.I#28d4aQMEY#6PK,,I,J2
6QCTUdRa5JN^Tg94\@)b:Z2M&P/16QEEGaSL#FCf2BDA48FT27@J/1LJ&EK#4Z4@
Y>MMCJEN3;f0Rb(\K(TDWQ2^;<a3#N>-7&RA3Lg?E8,O6FIe[?E2SRWJPNcIG?77
PA1#FgZ?,f\S)WILJR<&>TNTO&dPTN4M&^UXL&#YbJNHYC6a-@bOa17(bM^X<fOC
K?e_06/VVOUF7],&,>0#W@Ke=SW4\+a^gD#f1;D8>\L?T<gUGcRLZgg8g@IWW<&-
GW_\C8NV3ZN^[5+]LJTKfcQ+]-,dL>[b1c8Z28B5SUeO-gf9e8-Ldg>?9Wec;R\;
Hd.Q+#;cBaW<3HBR<//T#SKIa)Nd=;SNJ_XU/JI9K7JH:V<>(aF.[dAd61ce9)fC
Z8OJ(F@YUB2KEDf;&,O/M0Y1PaKD9<HC#>c+[DO^7dN,G@KD_G-64H39=LUd=P@P
GGGTJ9X[7U[b7IFS#^S7W[c)-#TX)SFD#69=8B>gO&(Z;7#>>KQ]O7\[E1gB:/0)
NH[7DVRU7.754OY4FNTGC[KYAe+=B(MA#(YRRaAW:UM\e@.<OZNf.Ve#.,1F.9@E
=K94&aW+W,_[63WZM>8T;4^Q_+V8Ob3dXRU]=GY/fDPeCU&H6CMO2[e3OI?a(-<f
@XMFNUVX53#IYVL^W]K3d;]eC,@O<7DKHc1-VR8U,&)14f-3[=RgVE453:9(OMV^
/a:TL+MWbXFJ\ER/3BQY/^YbU)G:GZ>g-,OJA(8<5f-1WeA3/B&]65IcJAK-A=dg
Mad.?;bQ<M/H7EEAMd[#19</3d3BZMFf:L=L[YKe0e:2ZIIba\[//HS2@Lb63U3Z
?<SWc2PY^D57:@P+df>V5IW+2c/SZW34)G9HN/=[>V?.gJP2(1)=@_^BR1b\LT=0
McE<T6gG22#IFXL.F?=)#,&S.#0.A<ZQUJ_UWA;dPW+Q\0L[C+F_A.3>,?OOWc[C
/^ZAdM<\eIa^W3<5OB8OY;\@a-9#U<>NFQX3XJ?,\a9.01,Y,U5ROGcLa<-b(0bP
X)HP5)-IZYHRHCOG8,-JJ;7BHD.S2;BV6GLF>VSPB/FcF6U]d]9553Fd_aK4FRQG
#GY,GCT[bIKaQ6#\A--@5ZdSFGFa4g4?G@7\4TQ[9TZ+=d)ZO1dc8I>[ce/+>a4R
MJ=)3X\0g(@-3)+>9739Q84CbDWHee+O?SF]c.W9e^T7>c1IT7aW;HB6,^]S3ZM=
e4?:>I4a/&&^NLYICZUD)X46MRX9I29=FI;;+=ZJP_E?FZU5Ib7L:_NO93N6Qf0(
:@]e@_EI?<^6+;;<HM3W@CCWC-L;EFLYS>XH<@6>3HMX,_U6MC6[,8GPVQg.NdX1
O&:Ig\9_=Z0B]^MMZaREA+L2K=6_XLIX;,6G]S3;<-^KXeYgCC22C-00F-G-X;D)
#4g)#;3@K/Kd,f0+0R\6DC6bXB6/e:54NA]-f,MT,KFIXVe.Aa\\P.0eHg=,@75Q
:0>0</d6D:\U1:H#P0V>,3YTJT]::.3M-(Y(E3D+/QWf[?C0TX7CIG2<DaK-/O=O
()ML9C#[FT3ZN/GARDSC.K&]5dG7U&>7YPd)/bcUT0A#PZc;4<\:fTK+:f5LA0_(
WFAbN?e(3,^g-8Xf=CI>WMKe1bU5<<@&bODb+H#7E8+&,BQ<0;^&g^MM33,R&G0-
Fc\ON+PS(V#/g\>0dP-/2-VC5dIXL(3aG(,gZ7W0FD_[24dgHAI=SYA#YXUNe&Z:
2I@.<;]I(F[fa;<W:dMLAXU(=U)QZc@=NgTHf3G:UP.:75/2.a3_d(G7\5=K@[OR
82-.WL;eaLQD#5aB^fH9AR:].B=Cc>V.g(?1]KYcR-5S9)aXDA+9UPf6d\bT5DH^
[c;g-:8[B&:ZKaK[DE(Z>NIA=@LXGXPVb\e=PGG&5BfE;CG:=18gKK1HgBAC4ZD.
O>8I]7MQ41LK0H>X)\?;XDSB1aJ+XeF.]5XGXRa0?cJ)d,ffDe75]SaE4PG6QdVO
4dC&&+C1#e04&I=EO&:Bf;4>?-.cgG=(G<Db_]H48<UJ2g=9g:4NKa_),X4?5J=X
D>&F4XS_eHMQD5UDX+9.G9T\LZ0+cb(MYA5gTE.0Z(235^>/^(20Uf@K7_0Aa=5;
NXP)Bb_BBUA;;Y>PMD-#Y1;\M\X7.QWXPgVZK0/FK4]GaF7CA3[]DM?TC5>dSXUe
)g6W?b&KB,.FMFS&5.EF3c;^WZ5@f7>]CY>?g1\I2[DD&]@+B.c5<@[N8.7d]@#_
0af&U)7>,f(PefC:5-BB31J:]0@:f7&)#e35NK\3,]PC9)ZG-Z52<f<>E+P7B0KN
dSKZB<_TXZDG5@U]6NL#RLXe99.X3V+#Z[SPN?K-7.JH@1XO.,T6:VYeO?:J&EI?
3?,TXRe&KK;DE/#=9.O)?)&\0)Jg6R/FK6;DO@OLa>?MS,BOF&&L2LgdBI1^_?I?
RB7<F:0IC[Yc2<Y^&R+<KRd6MEA0bR?ELF=\XMI:CD3)(GPfEOBg5L5)FZ)L-&W<
GGI[1P2[H66e67&1]eR@a.?73E[87U6KEOA0<VP]Je,2L2VEJB/D;:[#S+U>)X8(
+S[7YBFTBH4Ya<-_13+-Z,^WG:C_/9Z03VM[d17Ea<.VC8#fOB0^K#;@QFf<-&[6
>;\Z7V?2g-).b<eG9+K572C3NKHLg>-)BQ.U0g5ed8V=VT;/?@dJ1D7YS9:fL=N<
\3F/cEcGR;NfF?WMb.]8+5T-M:TL=B:G4:.IHD+PK/M)BfY\R7aN??e^-VAI_aBa
\ZHQ5,NYAc8RGDd77;08Q+5R+HIZ8B>cRD3(T70>b-HR27>_PK,DIP0/F9(N9?66
d?\BU]=A@>/:6T7B301B/#-9&U0(4Y=#G.;Xb_(@X>fPNNe&#;#Bd1dT+I.98BSQ
YSd;;)XMC1gIEf>cf)aec]fcg1..g9Ag:FGdKZV2Yb5/L>bB&D9+)\KM(,)[c2Z-
Q8]DT]@H_WK;\^W[L:L].LcgO@JV<I(L;E(O3IO4DIV,8VVge8,^2+IKKBTF:GNU
T)W829B_2c/8<B.b,BQO-00C17J3YXO\XMB?0,A-81gXDH>NW[@0GV,>E9^K6C,V
-_/eAI-^T8&LECaQXNUR;K.;3<a-(X^McV#9KeQGNVF>GMMEJeA@gO1;_;:97U?\
0#GQ<1G?Tc-MOdaOBR5N&]-XJ6bY@A+?@TGNgA0)9Rc)R8;2Sf<7cB(-Y;.O+^=_
;a;;^4g89_0_^8<#850O<dUQbOg,ecB.3Rg/BgI3IgT6gEVCA[c1GU.:IAT5\(Ea
N[d\9/K@2;GV^G,LN-.7XN4B)Vc(WgX5;ZYUX;K39.g33H2V6LNIN-dII1cG5UP2
,[+8BZ[0NPK^:0dZBe\GB25SVHff<cO.d,dZZL:G\\gSf0?<cPNcJ?BL5dFB3=OF
2G(-<_>J1=2++=fL@1V493(5M;-QfMNd&f^5b@XfURJNWIZH,1(gOCEV&M5^X4D8
2T72UeO9+N:5/N(&<.0Dcg.?/4gI6fD=NfXHNWe@47(=c&G4MH-7Q2Ve4L.U6I5R
:+Wd9;)IN[a>KXTJNPb32CMZ42C_Vab.G)(--^E_)^d33LPZMdX#)d&ANbV<g>JV
9E?1_]MLJYOB/?C;QX9bR66^)[c6TM3O7>.NY1S7ZZ-eNF4XX_dXGda#cD8b_,@5
]eg:3G5/FIOC[0?VM/#=R>H9W[D]^a#LVfg#GFcC3@?@H41>cJHc&@0G@HVCf0D#
AfIT]2,>Y(N/(cMa[aNK>T9L]ZI2]Wf5I=2.Tf>@5\WCV]dS5D,eHMZ7)C/g]0>U
8UE-0YBZ4bD6FfWWGcX3e1XfDbWMEG7HW0FFO>&8IS)Q]<X-\?ABSf,E2a7=GBe2
A.)GLgVIXYD&<[GGDT0?+UMfgS-T)4aN[]d2P,1)GVZE96F4-U6B(f?0Q+Lg;1=#
N?R3/NFd19U1G^cHERH=9E5/T[Q,@XX8I@J-+aZKGWS;?<RI&f^c&b?KM:bWN-UJ
39=gU_QBgG_[_,(e2ONP>(O9a&.A9]+^L7(7@ER:B36\T036D(-AS:Q3fP4-&Q3M
C,XHXC]\5HR9&UZS1AO>WY=+eN4+[Y;+f+5[XGY2CWP:V/:LQZ,gVJ<73,H^1W,B
T?N13^-89&cJO,K6^_(\U6d9\CJSF01LQa9UQCQ&)IG:+0=@5ZY(fb1NA=d,6LN]
96SCVAA8/,4,Q<B8K&SCETA)?C>DGP36,d_SF0C?@f_#XX>bRgBg.8BNDQ[R?:aC
[#UOORIQ65d^<?UWB()\N>_P^6BOE_@#gB\==XHC=VF^(49bZ+IbTDFA6GFD=;EY
WBe&fc?TLARCXS?>BB6g9IB2c2S:YZ,FP-2Lc7/WH=T<c]Q?E^BNJJ?O/K5>0I,:
;_dJ2G6J-+dNZYaWMHJ,E4Z8OP2ZC(f,KA3XS@93J3b-Cf6&f?#)<;^:ZZd[KO(E
5WSU3?MFdLf(d1c^EJC)5H\dU.H-#60=DE#5GVd<+3c^GB7B,0_R?&A#B=+4Z18c
[UUFESIUb)66f(ZOB,X9NK,N46ggYG6]MMf[Bd79A<S/#[#a3R?/U-][V+L0<aMK
KbESB-IYgCg^8eV3J])5Z:Ae+#_@<>H+AS5&E;TM0W4^fP88I.72.QMBcL-QGGTP
3E1D@^.>[bF_;<.cVLcZH;7R7)b>P[=BXHS#JD^dORAEe:O[]I?;.2O+;N?.#;C6
V-8aTGLP@TOP#aTS4.TV@d4T)=cWHEA6>N,89Wf<_\JP<1;A@Z<H5P#[d\XdE0<6
Q,A3+O7bOY29#5^4eaGT.FdL^e(8J#3E[]g(bc.Zg4(]g/;_?JW#dHaBYG/?HYK:
X[48-4VJ\RKR@X,0C2]3<;A><bC@-JGH9INg56U0=Z[(TQONfCLOF=]bY\?(IbCf
KDJ(R3CPI(([;ON(;N<+]9X&/MY]c42fI.,?S1N:BPP)1#+MQ@CWS5.@80)];:)&
^N/FfRf0AKOI73/]We]X.&YUCB:.>eBaO8ZY:[7.J5HZ1G0-(>.Z8c_-T,De<eCK
gWTR>OTNJdC2\A1e6>8K:2;d<6aQ<;T)gA2A[(1@ZU8#b^2IYdY,:C)_/M_MMQ,^
S=)=&_)0c9^_-/CFKf,2OaPSSdU_Fc\dF;C^-\C0g#@Fa2Z#bVIFg^2L^]_D/DSH
^6^<P>MT3a1D)d12aB.+cH/:@[#7:]ECI#U[@Se[>75eb1H7eO8fSGVPO)@Yf0b(
c1gP:g/B\+T/_geCf1#_=.W:UYE9L@FHJGA[Y93fM-Ye5,,f10Rca[QUH/JG+;U[
J=egc>X\K6fJA,c::75RJ=0-a>/]/T&gVI;fCZ0;=fF+O3X9)8<eA[f?92R.c+7e
SJ_T[3A_b]YNB&>_@OOAE=Ga-B]b+HO?gg(e\RG,JNN@;YK\:-1Rc[&R(Z:S4PPN
FDbQ<-]dDUI7#(bB>?KL2=[91f)()e#[;HLUS27QIaHZg#\P5,88Y&Xb?Xe:_QSZ
H/+<-7;AVa<[[B\A:)aZ#Sb66S53XI4?VaVZ&db]S0K#b))0KW?gOGXdVc[.GKL#
FWPZFM=791DUAK+9VSI1J=USX\LVR37-L7gS61ACW9YdE+<?C@f_d2,NTOa=U;2L
X<PHeHd8<W;E3D7S.dH<&]eb7;.e<=?&[Me4QF1:ZBI([P.S,87=]14YL@V)Z7:4
:M65KH),F@.1;,#8;cNI\:Z9/-W)#><4AgV?f(.UVP(af=8X85dRbL11<F8Rb,ec
[F?BZTKB2b:,;J7Wad4d?4ZP6[:?.HT)>0g[3_^&\&RBd<FG@[U5,+1P)NKe6=8N
fYgcAFdJNLJ;/BCb7X<cE@a(]=9b72(W1<CF>@d2_c@NF/J?_R2>C_U#B-Te&A+F
OJc.U@3TgaS6Q1#,4fK25fD7f]<P<:2;F:/)a;PE+Q]5)WGE(XLIC0UB\]K;OO+7
[^>CL<T])14_c/>&_624:5cW[d3KO&Q91KCI_b>V&dLGX5,OZRg-c/39#;.]]M-K
QI##_S21J;E-E\#)#+7LRJ9I1CIL9U7ZVW2R-?J6^\3IAUV38VJ<C4_>34PH9KQW
UOI-FZ73)V6#5\:S0g7@BU>3FS;RB,>d(\TeF:MF,=SB@1\JGTSDD1?K?2<2fMV]
QLaV3)K0_VG.g.+T-gN8EQ@Q4)/U3bDW>,1LgA6,1b4]]HR+H<.eIR6?f:]f.c(c
MG067-C?\bBbFJEOSQ6aL_bGZZ14g#P+-=T27)-9,4M4&30R@IB\^J\;ZDM@L53L
7_-V>G3)>.(;aUL/KS#8UXf9+@#eJJ)P=VL?WBQ@f?Aa\Yc.GJcRA3>b3)ZOX9?e
R(+,UY5.7;gJb);[6D3@55ILHSSQX_\V:?]_J&2a#fP#X/OVF4UcWTOZ.KL<6+XM
>dNUNY-bN,Kf/<2#2HK^2J:ZCUCS]4#dYRA=6M8MY56-e+ZO;M<@2b3A5cRcD)4g
#/0:LN],2a;O69Z,ZD9-H=XI[=DNa:HIN@R0gHHgcV8:RZFZ&ALOAQ+]QAAE2dQ\
c;UM<=VEID/UF]c1P4N)EMQGAgF3FS<[?c6>Qd.e]GZLIAP@_3=&.FG<^2e;\#V.
;gFKB=HVIa=eS01D;..f5\JE.6/JAMHFd6ef-YP[U,bLH$
`endprotected


`endif // GUARD_SVT_AHB_CHECKER_SV
