
`ifndef GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
`define GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
pQlsCP9BSkh7OmNnHHa4hAnrs2IoVujBn+MQx5JFTe8opdix0+gAIPnX9NRmdWMS
GcbbrRbuOdc7driccENnWZN9B+BFusE8A9ZaYPcfhHkP5z1yx8yN3faSVm/agcgs
svkDWYq76C7G+EdHyMua+26xoMSeFxs4N7i0J0ecSvUPQVNw/5EP2g==
//pragma protect end_key_block
//pragma protect digest_block
lZpG13LUocqLCqMQNxVUwQWvpts=
//pragma protect end_digest_block
//pragma protect data_block
4z0PzsiRo19XSvudVJvsgfG8ZfXMdF0/tkALcIsHoLwLiMVMk1JHcnXS4RzkJoHo
kqDhte3/YLqWNjwktT7aCTm7VF2dCaMbigepvED1IvgiawdOwcUwrmyAEaGPk2MW
OcdEIGxuvoCN8pdL10db5CvpftvW9uC410lSX+1E3JVdz5I9VE3UrvMCB2moWOVQ
GtnpLLbkV1DFS23PTFmTHtWWzDXJOUDsZfebedl13d1vgOkomqLCxE00Ugd85skK
r13Z5ahdgTdbL4QwtGp9T07l3tf6v+VDawVlNbYGAjWrNRiV1Kkl3w/QmN9/dHiR
trt4hUzgxbb7sy3MMoU4qtNNTKH34HWIbtXKkac+y66FX4QUPalUI6E6FOGHiSum
P81r9jbaN0u3/78cRZiocF/IKom0rR+np595WO7lKd4TA8ZzHa5THsxnXB4/vuAN
2bqOXY85Idn1fxNv2Bry99SfNmHTkkQnZBX0te2u8IHIBZTp1/h/BUHkTbVmp84H
mjmMSMKpXv78zue4KWnPF9JIgoAcfmHxCEr8BuQUFPxL4z69JEaYMtNKybAyxo7p
O3IQu+qoJO5cpLVFh4EZXhb/rnU17ap2nCsKVSn6p+GhoSjgBIZvoD+qwOnTgrLY
ihTeM4Q8Qi3XmY75h5Goi6N+geGVCLE56mNpbZaoWxhJaoIroLsdGqkZxJKinSRr
jNX7ucdC0tzKU46GVJEDlpUWLE+Xp2IWYp2KW9zNMYUrOalQ0oU2ta4d3Asn7+V3
iXP01EwlP2BovFptxOnJFJt82IAjiYTtVMkFql0WszoNVrb7xKt6J8ZtE8J+qtJE
mUhQnNaOmJHa/fHXAKWHh0pCIMvLtRqK/Tg5d2WcapTpiGvUn+c3fXw/4Fr5wdne
Ls62qeIVjkpvmEE7nYOXdmhhGPh9dfJt07QO7afrfrh4G8tDNM+nXGM7vnskFLhg
KQkeuEMwTWlUzCVSL+4dghxVNppw2jDh1cbr/oDAohjDI6vLlDD6/QMDLFfcoq+B
cMpW3U6mzI72r8HH7cgM1CtZ6oSVzhbZT0ehoCjbIoE0NIo3QyhO3YTDUTUAlsZZ
knhkCxoLM2iuc9984QutDivVbygm6sLB6P9tcoo3h/X5CHt1gC6UQtfxV/R+R8ac
bq4JB4AwOaEozpLRVTjlN28QLtU6uPYh8Krbwe8kczmI1BaswybHBFqGwjvMfoUM
rvAotOK2p7ciiKVPCqYsZ/EO/YNBWCYGvZ6ECXIemHQZgpoIPbED1WBBHoTttPQC
6/L0wyB7L6jPPq9ON38Inal4gNMjhfrGzCZMsG/cCNbe7cD0blZTKewrseuffKQS
yoN9VND8ill67ufdXCLbW8+1tSpQ0LjvZ+NnE0kBT5CmH8MFMxXeWq5VA/xYYU9L
Ixl+WncKpaCWJLHadI+mYq+r2o5Ra58RBRCTm+eM/Qmq3jWMOp12hY/bP8MJD43p
uUwieIBBbPEcobubr5jf4m0Gjsm+muct870B/rvBGMQjlg2/v6JtCaFZSur6M7ew
y/zhgfxKiZtJ4vjyVwmWsreadpeaChgbhQzeoX/wFyMldivNIYqHnxl/TzOp7pC1
ZSiWRVIMrAlKFCCspOLgwtfmebLNbXTHSeUdPP2EbSUMNz672UE55EmqpO/hVfk0
JQIZB6rbUBkH1RuE6auLPaNXlLsLeXkw/FPsEvIxmFhtpQDhApesq/1wxVnGN8qO
rul050T1X0oljhgNy8XAxXZJEpAWXp65Ehs9peNTHMTkbzq5ntrTF4NtRqd8dQlZ
LUBEBPclBK/xZbpAzbx2IOdU/55xP6uBDlxVIH5Trda/MF+99sVl1mf2UWyev80r
4AM0TFbmQGpHPpCmnyWJZXwHFqK636caZtHQcA+ypSVdl1lmVn37HtJWdAeLFEP6
u+gAAR3ktqciR8PLAUT6j3vellZ58IgjYsNWYr2RXFUKC1h/FnGR/AAacgwdAqwB
bK2J8lvCgIn6HWe82tf+RK1zPp5EOaynhxS+8CZwytj63ifRlBR0GaqTIh3IbqMU
XqfOPj0wZdmEkULMKktfwZsUiqoBBiUfMbU8FQ69P/WxBZAKDEJvfGGuM8laXVN8
74cY/Z+kaiWBwK8YSbxyme06jpP922HeXjIS1Kd5oOXZ6Z7XluW/kXhNm5pz+9bi
9e6MgfK7dTTup7v3BCLZShWZ9AMmAriExg1elN0D6KamZuKW41OtWZqt3BGjIxPF
GkSi3d5qeYsZjzy80Z77W/eKErrWZ9c5ii2Yfj2I5DclF1wjaGBaGDWXmYM0zDYt
TQzolMPPfIv9k8XT3hwSuVOyAIS29wxJBX1GDCFKzPcfb+r83uQeW18kG1qIzEJY
M7lebGEwEJJ8Vb1Wnt99IaQd66Fye1hMpaD2KGSzIoSOMmRwSsnJVqShmGxYv6GJ
yzZqWcop+g0AyUJg8AsN1rSG/Sa6xP/l94rcSdzbWRHsyXRe2x9GK9oS/TcHbraL
tB06kd1ZgC+MtTX7gKoo8WpnjYKNpw0kArnpUwInf1a9/aswSb/NX2GKwTsq9FiT
ZlIfwvphy1lNutWchZrnORnYrxqz/hyVdv5iTZXxZz5XA7IIxb+XYkYfJhHrZybs
ZmFtqkY3H55VxHEg6TLl4xMpM1pxzGtf5DC2l/LUkyLZ0Ne5UlSbq/GK/1BA2Lfz
xSfOQRpraLRd6Ifjcxg0rJG7pHNfAOh65UHIve9AHf/evDnpYct8Gf9kFFHkiwlP
54ljR6E2SEE3oRcnKG8sUpKVaFmzIOzHnBol+moPLve8F8Zh+sVbmRQZbqfO83J6
nR2RxDjf00lIcFVDX2wyk+EZY9+dcFr7mZzig98vzk8Uvk8gzUu26cFAnoo1AiBM
dZplx5d14mF3I9/b4r3oVELzwrMTueJeCeOYsGTXWv94aC/eCfRRS30bjWYLwPE2
l+oEdkX5u+XNimxKh8JPWjFbUBCEjLLKKixpl/MKAk6+yZyT6JcCBS5vZaCCa3r1
3An7GWaJdIjNKvc/lBYv9nnBk81zIII266TwOv71HhtOioWzmmuHe0LX8Fy5ZXh5
3+U8omerss4R2qS4jaSbQGKLVh/vpgVcTkz/QYaJL/YxcXHvDH3aHhzYOw9GSzWB
gjJh80jmDo2L+eOFe0uRC/urztSkbzIZR/5x2DbMEnq8MtVdmcg+DgEL2uwvxu9u
49WX5S1vb5haYp9onlqoojEGWjj/mRsEM8UET/4Kte+nAD5sm1E8xLOdV1Dwmccx
KNhi9c2ezzP9Ta4edf+JUpMyOjxvtbfymUBszoA6/r7y0AG2dyBIodaeoz2ebVmW
nhAE9PnmkNkQAh4KtXEllSUIBzgO2seMT6K2niwIelq8jLy+/GjFGBkC7breqTc5
Q3cbkBgb7EKIeqBTMb90cP9H6mzHQSQtyWii4qPAiICd8wLX3+Qp7zI3X2Xx4gJk
JXcrKgggpSEfXKcRZmvK/1G276RBurURxHG8cp9cnwKofXzg6YMmP3hIK5DgqUE2
W0FIIIuQxdMmc0JRWdm5dzvV2YVqKhdiSimRlT/Zgb1cx9+n7lHvqzQOyX4ewH9s
6J1141Uzcy2+zHE2ViIAs9NPiTvTMAIwZEm62gtVsrLCzcarAscObxkYHDZDqSNy
2x2tcfs+lDXFm5iXQQfaygRa9xPS5yiF6MdDJ4t/q/g7SKtFUc2p26NDX9+F8fXB
RKF6yLKHUjjYb9MRj12zWKULdwYNnMMn+ZPTOMK1ddtbZyM/aNVE0XPxcTVddQSe
YbbKLexWw1G6hYVNuwpARVMSnUiESpPHlICdQSSePv0Roru27YAUSNsgAZ5+wnLR
yU95+bSLu/aNC5lHgRxD/YLRG+uf+nGSQ9eR0fFBnUcjlihkF8ccIflXlFPpKTVb
S+CmzZcMcE3PFN/xY9AxrUHRSTs/uXs/7cl85QN6PKkFufQ66Vl3pYL3ctKIATUJ
A2QQP8LymAmzNAGgf6wrOtDtULQX9VTCIxzRqDAxYba+GLoKF48eyWl/oMoyj7nl
SY5edDyyQdMsueGFPsoFePWy9Sukh7KfDPml09PhMGQtORFN1wTsdd47H050kWgj
9YHyj62WsIZgTle8x6+28Os4WyVzPIV6VtY6ffNHsSCSwSvvc/keeSitFJG/3GYz
4InZ0KQx21SPHWRLgAlAuVt9607QDX9u1aev+QqbAM/4Pa8JPgF7ECm7LlPitPQs
fJ7WDI8TqYD8ZKzmPJ2JttCPg8mZLGkf/Xgxw65BvLaaw86ClihdQauHD6a9kVKU
8MNFckN+DsW2NeMSLECvvm6PAiRFHAw7zDrYmEl9JRZ6RfzgEW+xSLaMjZ6Z/ZNE
KkLj3C//0t6KBWO49bf9yl3xfkiYiTm7zLKFJxft0kk4b2fpqQR0SjFpyeXdM9iy
mMUoHEzf2XqFULQ+zakmPOCJO/zcwSDQC2kiu4HLXT0r4kXzJUEdOfqtrMGZdNfL
AWSwAIhNdNAWfQ5YMft9iaXNqUC2JIBwH2mEeO/EDYByHiIOu/T3N0OokVx1EMBM
ryT+ikvO/yOlglk+Bs2+sIIAaXZH8THO/CTOuPZBmGcWPLaeSEOHEQwOLHpQUOHw
oN3Yth2A5X+hnMVnaUENlcDc/341NjmmHESn7eOaU2lNoZ5m5/wQ7XWpWMyOc5RL
4sHWIQGTIoj3nad/9XtRxVK7LUT7ga1NvBVU+Z0YsmNgcBmT1eZE6D0iMdiH9/ec
3AVxnuvmpI7dpUtO1CTn9k9+FZrF6kitrSO1XS/Iml8mdgt5/E3vCjKvG/aFxe3x
JLyKCRr/Tb1O+VPSCMLAW5SFKvJ7HII2tYIeC5k9HZ/z+de1A2R2IqqtW1/ex3Zg
fhK7S/pBAc1zG2GNTW9GglfYLZh3kd8PaSPST8JT0lPgDleN2XTO/BJEgAxI6zQb
JJXktj9RSz2i/rgZWJiEJA==
//pragma protect end_data_block
//pragma protect digest_block
eGcEmctXWyLFPbjVEBaceRb6wi8=
//pragma protect end_digest_block
//pragma protect end_protected
typedef class svt_ahb_system_checker;
typedef class svt_ahb_system_monitor;
`ifndef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_system_env;
`else
typedef class svt_ahb_system_group;
`endif

 
 /** @cond PRIVATE */
class svt_ahb_system_monitor_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_SYSTEM_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_monitor_modport AHB_MASTER_IF_MONITOR_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_master_async_modport AHB_MASTER_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_slave_async_modport AHB_SLAVE_IF_ASYNC_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_monitor_modport AHB_SLAVE_IF_MONITOR_MP;
  protected AHB_IF_SYSTEM_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_MONITOR_MP master_if_monitor_mp[*];
  protected AHB_MASTER_IF_ASYNC_MP master_if_async_mp[*];
  protected AHB_SLAVE_IF_MONITOR_MP slave_if_monitor_mp[*];
  protected AHB_SLAVE_IF_ASYNC_MP slave_if_async_mp[*];
`endif

 typedef bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] ahb_sys_addr_t;

  svt_ahb_system_checker system_checker;

  svt_ahb_system_monitor system_monitor;

`ifndef SVT_VMM_TECHNOLOGY
  svt_ahb_system_env   my_system;
`else
  svt_ahb_system_group my_system;
`endif

  /** String for storing information related to transactions to slaves */
  string master_xacts_str;
  string slave_xacts_str;

  /** System configuration */
  local svt_ahb_system_configuration sys_cfg;

  local int log_base_2_slave_data_widths[];

  /** Report/log object */
`ifndef SVT_VMM_TECHNOLOGY
  protected `SVT_XVM(report_object) reporter; 
`else
  protected vmm_log log;
`endif

  /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;

  /** Event that is triggered whenever the hsel is sampled for active transaction */
  protected event sampled_hsel;

  /** Variable that indicates the current active slave id, using which the 
   * sampling and checking of hsel asserted for valid address range is
   * done. Also used to bypass the data integrity check if no hsel is asserted */
  protected int current_slave_port_id = -1;

  /** Holds the sampled values of hsel from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[1];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[1];
`else  
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
  bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsel_sampled_value_copy[`SVT_AHB_MAX_NUM_SLAVES];
`endif
  
  /** Semaphore to control access to active_xact_queue */
  local semaphore active_xact_queue_sema;

  /** Internal queue where transactions from AHB master are stored */
  svt_ahb_master_transaction master_active_xact_queue[$];
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifndef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   *
   * @param reporter UVM report object used for messaging
   * 
   * 
   */
  extern function new (svt_ahb_system_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_system_monitor system_monitor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param system_monitor A handle to the monitor class of type svt_ahb_system_monitor 
   */
  extern function new (svt_ahb_system_configuration cfg,svt_ahb_system_monitor system_monitor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Sets the configuration */
  extern function void set_cfg(svt_ahb_system_configuration cfg);

  /** Sets internal variables */
  extern function void set_internal_variables();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the data phase signals */
  extern virtual task sample_common();

  /** Adds transaction 'from AHB master to IC' to internal queue */
  extern task add_to_master_xact_active(svt_ahb_master_transaction xact); 

  /** Adds transaction from 'IC to AHB slave' to internal queue */
  extern task add_to_slave_xact_active(svt_ahb_transaction xact); 

  /** Gets the system env/system group */
  extern function void get_system_env();

  /** Process this transaction and execute relevant checks */
  extern task process_master_xact(svt_ahb_master_transaction xact);
  
  /** Waits for transaction to be accepted */
  extern task wait_for_transaction_accept(svt_ahb_transaction xact);

  /** Removes transaction from the active queue */
  extern task remove_from_master_active(svt_ahb_transaction xact);

  /** Checks consistency of ahb transaction data with memory data */
  extern function void check_xact_data_consistency_with_mem_data(svt_ahb_master_transaction xact);  

  /** Gets the memory contents as a byte stream */
  extern function bit get_slave_mem_contents_as_byte_stream(svt_ahb_master_transaction xact, output bit[7:0] mem_data[], output string target_slave_info);

  /** Gets the address banner string */
  extern function string get_addr_banner_str();
  
endclass
/** @endcond */

// -----------------------------------------------------------------------------

// System monitor cannot be supported in the INTERNAL ACE TESTING at port level
// This is done in the tb_ace_vmm_implicit_1m_1s testbench directory and
// the tb_ace_lite_vmm_implicit_1m_1s testbench directory where we mimick the
// behaviour of an interconnect port. However, these task need to be defined
// so that things will compile.
// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
4S3kwxK/lHdIVOk2xnAYjw2lKUJLc2TnDRVVlaPPyCNdu39oyf+5zK0iOkma0grZ
U39h7pdzJOwjDrBR7HM+1bWm+Grub0YJPHE8WjI6Wy8o/T6J0G5xqC8ERyce/bTB
azYgWL7bHOQWm29bdwVRDXHYjdn/yn9vbXFakOCWFDWor5QJOcuacQ==
//pragma protect end_key_block
//pragma protect digest_block
CBMCz21kFeArdEMIRXzOmMozJVA=
//pragma protect end_digest_block
//pragma protect data_block
SMF1YVSdP1w8MkSsvDrsoTabu1CbP6ZyV1gWVFZEVokSdWO9vTjvcLOKtECH4O56
kCsdGWiXBEnFpo7zybh/ZjjynEH5FROf9CGTh6Fdg0YukRF9An0H//7hUbvHwvzx
b9SO4+a6+z0iHSUTw9IoYjMojIcTQSIgxMRa1aWWeqpEN0BJ3khbk6pOr+bIMSR/
0Q/dLZ/kRE2lDlXtQZi+xax8+87SicpdYHAFvLA7QKTxd9PPcUnh89k/J8tx3Ytu
imRGU6IPxtLCg1/GBTasb3DFPtBZU0ynAf6CoMMOC5o0ciMSXy3vnwCor0V7o1Jp
BNY2thOytiCLQYm+up8Xh05y9b9vLb/2CFVf36sTQEbKDl07662wtR09YEZQrSNM
90W5FWbOEXO4u7oJ5NpQPmnP0eNb86zE53vPral5h38eEuM7XaTHoISMhGsXS9JZ
M3MyS91dAnlKhM0PkEAWLazP0Z14R1+0XnkbvwFnbD3u5Dxwgr1/OaVuE6oJqZkL
HhHRi1meIAsoKaVMg8e1KQwoQnLTXCBCSDEr+7LPUCvsDD2zf2qakPZCVXit/wKY
Uh4qNfDFXpJjngfdSCxDMjvn7+YZQwZ99stq5h4XEcK5uNuv/Cmi10tmoIXqC5km
0GFbj3US3h4/KHFuFDPpU5UFIQQPUzcGO54ZXQPB1RIO8bmvMbPmUo2TB+9WSNlm
gUI+aqo4h/MiUV0mukk16IiYILFHti1J0jtBgyUGoZH0l80BMXlGQSnA37sfA1nN
wyrqBCNNSCDwYpw6wOAb7u8fhUyBLXFO8FChWcB+P+aPc8eEmEdwInkpT0KoMoiu
eR6VzjBM2uljrosAd47YgVOT1uDOEOxdxxn8BrecojRV5o3sRdZaYkCdXdLgv5GL
989ihEnOJ85iFVWzk130gn+BP2gZlVDc1qM6M1g9fSl1dsXpbeZHCr7QVr1NA0+u
glBkJgQK5jKJu7KHb07Oiyfk7kfiJsEEzvouAJOq7oMXK1qvSxfBbRQiDT4DTCkw

//pragma protect end_data_block
//pragma protect digest_block
RexNf21mjmwEBzpeg2dDfe8ZuYI=
//pragma protect end_digest_block
//pragma protect end_protected
// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0eD6cJ4RhJePbv7VVH4XBWVb2j1cHGwTirlgTPotzGV6Xg9G7FLRK82P1e0lLLjb
yWffn/SyNaopCxVwEz9lg4irWNqYVf1IftEGVBjbBv4PTuPPcu5PdOojK+qz5X6I
/vhnxWul2l3nvJdfFCX6FAYpaU2N68pOnshBKCruEiSDiFEirYV6vw==
//pragma protect end_key_block
//pragma protect digest_block
ssvvqaeQU4jJVpCXgJEwwFSwTnY=
//pragma protect end_digest_block
//pragma protect data_block
L8VKoWZ1Tcsa9VUsdiO/tLaZQcDZM7ebjFdh8hNF7VxBThczEjHIkvrB9fbBADTo
IBxFPy670o3zZjjkiwV+fEEopEwTUwsuLLJXEzOcO81DK9I6sqUstpK7Jz8YZGmq
KhvyfkHKq4YieKvviLD8XQwlztnJIqrDei1b8sCpBW9syFo8BuDe68fCUxD+xWhr
AZCm1/h1o79c2bfgmM29d3TQQ81zBVrwf4us0qcbfR/5QHC9iUCSHJse3030AIit
1RmW3hPiggW8x5FkYmXUz+KS4MLfmsg5ltO8rmnRQ/3lGEdt0n9wIBrTFNsphuFb
I0bBqKq9fapk2jO+MttF7ublI5TS6Nz8rriE3t2IxBwLsU3nnnZWQhTG5otBF1jY
L3U6bZsISBEdvxDFtM375cZY9xpwKKFqj1QDS7AbsnU7uMZFnBc7XV3jNUFW027e
i+yJEG/xpJmbkMt7qNGwAkVZMpbn3sl7dMZiq9dT/FN1qTs9U8WTR6cBg14jm2x3
ZeGz7K6IfYA3F1r3H82aFRLgDsFOBqRsJ37xDXXM2GLJHaDMDSsMEbII+4EH5AOW
AqoRlyGUO+CbwueWDtsG94RWfHe62FTz8V8m1WFeO31twSzFjETXBw9+QaNHfzkh
TLu3+DSH1p9V2XAe0doPCZur63Dh/QNNULp/T4jIFxceXMxwX2bNpwxvDjPWHwkX
uWIuMj9NxPTjC4AzmBd1XuLEVcV8tdUZw+l3jXaS/fDjjcOH0fAoTN04gLYIDqmR
V/eycWoOQkTC63TZQo1GqMltOuIEj8mcs9IjAs73NttZtsbSjKzLScgalKzcial8
DO2Ac4zPcgTb1TWXDvTDnQ0NHzut6r9MOXE93krvT3sY+VooQzvFCAESLL3vJcna
m4zasN5t5n3nF2L9etjvTlEaqu8QFX8mejQfvLLmroMwi/MABribzjRr4q4bYv/2
73DEZcdFrfRBUcORU4kPfilN+kVv8RpV6xK5lgLX+rvGjlH0JlkLZujPbSmP4bCx
wAYIVmPrT6YP7biS+PTqYAdIB/H8EREKioZavzpC7vVTUF0SMb89c9a6VvbU7mMC
D3+GZs0bTBURd3fFsTnqJTS6lJB2M97Cj6KdyfIWSYRyZegiHQPCRM+zDAZBB66u
1pptn+JVl8rM7oSURwRfd0+CQLJ9yEKeyow17DYPcaKrdJu7T/zulMpY1hkbtsvE
9Huep2RYwZ2iNObQmWPAFIZAMTzyP6T2KQJa0AGxgM8MiqTcqcN6vumT0WBBJP+9
QIe0bhYWYFtmvXvU4YgxfVyDrX97yeE4GpjjYGU88wojRSxHIxZZC1wm0NA+z8A5
p5COFCYEUNlqiWdB4L3yqEAOF+t1SLHTQVpbZ6/YIxopulBnyr8z1vldORskTqNC
WnneLcRrDpkfNcbveUGdLQ4ChWhPEaMtt5CozfiVuxoPmuVgmOhLlEDs8X5dQoSb
W2UC0VZDG9XwZBcRUU1uXgMapmKhr2XdsOYJ4ydH8cTBzbyoTol8gHtKGubgRUqp
0FLWdHakRs5YKyu2hcFB5hlfjxP/WCAY9+Zz1/tv6SWme9Vb0Kk/pXynv8zG2s5Q
x/3OpN8RIeMwX6xyn/yz8JPAL6wmjjcuAUwhKcbvGAF6e+UpzY1yIZ6/t+OtnTyX
Ldip4kNQ/+7EUt8Nk3N5rpGWHgGeB0N+Hp0JM2uFbZj5vgsGpBxprYiHGEjjBSdY
NhXTbGnOUtShb3RcjssFbBOYOFho+AXuFkTXDGkvCphsiJAiQKmHKe2Fe+gG4ci6
NOaakiCA233AtkmVIKo5KQjpPUpRZaHPdOtVp+wgvjZ35cW+KtYpE5ulFyt3bYy5
4kXp9Dbq4h4pU+/8UJL3LdIVws+K5v2QXJGusAMJClfgkalc7vl46J1wtgXomlnN
4SSvQBEL/HhizfvTtBeWRIvubHchCneEdhR10/zb4yNS8F3aTAobNEEjWVvzP96c
QkSUL1DRFBHXHmz5cb5M0CQw6rIui+Akqwx+uA2DSJr2xDMOAuZWWVrsPtqFgBeO
TrtQmZaVIT8hIN82Dfn69zSQVWQ1qaQkAX6xn6Dx1zlLzhT0HzVvru+MMEHztZBY
hEaLGh7fUbZYoXeWHhK50TRonVvcKUS+CfuK3XE/nXemrlhrVtD2LXcg8QZtOAix
iGevSR4Br6WtWBOP96hDIZkGo5mDpAyxGwbfzDrSd8M6bbLIxfLqfVhJsDEKNGt6
6jt6JWkaFKeZUxJj7iFSq+oHNq7BxYnbHI3a+HUBGsa5Qfd2LCh1rtXOSe0hG6dS
cYbalbc3mU6n5MiRAbL+YNPI/ITVpntVjH0bMW2KSA9jXECyZddIPkGhp83sHNut
x+2hC43GPVyouIRZYOyRN4LG8t7M2fYSxL7yDguar0MQlmzASuEsLgeaJcjqLw7I
7xQxWaRD0JaRTbufIHvUn7DtKxSMQqYw2TLRUoIcHf0pIdiHPlbRHD+MfMw0OlUA
NkHxZEitFxQhz9R2bVwB33eVROZs8M20ASoMkSa5mSrLKmRGKxIK3TC4PqC2S2Q2
g1EEthF+rbmANbdqEv43ePkbYjkx0eKxYqwyeOJ8e5LnUiR1CJomALqvBTfrTdAP
dgo/zdfzznqkOVe9S8kchmckgDcGeBzwRlRGoQhm/JfP40GZOjJ20pCNDfN5W5wp
wNOnw3pGvUQEm0pf8BPk1SRsjOIx8m8dHdn8k58A5hn+X/rYl/CtsXwp5G1uu3ns
cVsE/1G6doePv9wA/WGH1g74Z7saF6XtuVQ7aeSZfkVdLw9XBpX3RTBPybLl5+0i
6ZBdtNjd1jnokuxs5Z6+WA91QrtUNsx1sNu77xdv9YhnDek4+SQb7BI3IKYoBvA0
ouK9ect/X5JRLICeQqV0+voC9DNhuxyjFvz2Xg8d/23mOhxdXvHu3/TlTLI6yLAr
uRZvhrLx3Sh9lZSIdrLGFCfEd6OdxsUVzSHUBhPjgWArvrC50PeWAFpDJ0gmojY4
8d0ufWn+5ogV+V6pMLnSPIFowOVj4BOTY4n8R/b22RKG5BtyOTmezrDrxDEgMuku
p/jVqt9GM3ZWT5mWOpXOpV+yAOJ26ASvprYIb5+fdIg0fdFH1FNy5lPK40L0I1g2
5tW3pu5rqCHoKyI7HZeHotgfXTewJ6JfpltUUtmWY+QoyfTc/2O9fjRY/lbZ1VOX
8vNDO+Gi5MlF1bSSURt+wFzZFyi8rcE7nHjcG5PHeyK8rNpvSkYhVr+dbmDGgmo2
qeWww4yaBuMoPxsEvUzrUzfK/qFQzRVFk4B0yeD2V5LLz/qkxUPhCvFIkkZm3LqD
jhO3vbiRXQUXbhU18/Ciw4fyUTs/7Bg/tmWKAcd0DLgFmY0dBGO4NCGX0ySICFx3
/TsKQ8XhlFX23VspVtqzgcLJaZv/aT+NlViIYP0W7j/r8yt21yRDF3XAccxByVu/
feOnsfw5lGGqmCsWIIHFGdBIdMMSel29rYoVG/1UW7ytrLRTEEIM0asroahTosPe
Df8z4e1F5exM85fiQ+K9ed2mtSPeIdwgiJwKoTniRN9sfMspzpu5dPJmcn+PW2mD
4IcuOkYX1Mtx2RiPJ4/g3O4NoOT6Q0DucMxLbbdPy3KN2HdGwZ/sm5M1DZ2CmsA4
rq8cmTkOeWuQk+9r6ArsMBRONzDkrJrQ5FNZ2SAjQw6q65E7CMO8m9I7Y5jOxiu8
4c4UWG5z4L1pg94+z7fhvemdrv1VWj9MLfu4CilL90iEcM6xri0yLNF8FtQyL33o
4ElJnkKZcjzkQ7rZJbgSE3LQnguxgbi8fwe1F9TNFHeXuoTX1WlR7C2qtT8hpqrp
25xgFSL1TjLe9xUaXwQuCLm0ST6oDKo0P66tTiU0Xoyk2yLTjzb1a9i85j6T2l32
yDyxdZdh6SADX+tx0eH093MSgsxEUFyYLZ68TNqJLdRN+zTKyGU8iCiyC29GekrK
Uele4R4tyWqAmnDREYRifpdOw2LRLWjigfkkM48di25TzoeIGmEaH7yMBH3//nD8
wv+OLRsjqtu3dJ1q3rRW82R8AWbiQt6EmQBU/lM9VFg1nsQTbWPMBWKDraLl7e4O
mhalF0RG1DT19kwzTnUl2UQU9E4Bi3EdNvzeptVVhiMHLoks6Tx9dtaDFXOLaz0m
BN4s5Nq3G6hwHTSvbHzbchQRQAsQHfkXEHEiHb2vPlaL0WJEed3AcHnbbdaRjr+D
p+K2KpNbui8sOS6Fa8D0EYJET6a44ttvgb8SVKkHxagWwPrViYQyN/KCelLPEwvJ
L3W2p4iSeznilLWYojDnDq4xZxKxcKX/pQvSwxlk6Tskx4uTaggMcJrWsBrfo4kZ
endITAeCHEvuhbu2nQN6fu9ybjM6LjNyFsqZQW3MLixXr5r3zaYeWPiK2nl1EIeN
S+kB+ru+FbpoeVVCVJg/VibPfE0IgYaGSSQwFkrT45ftAVZkAy2Rt93Sb6QamzA1
4QYqZ9dm36Yr3uFWY32b3AIaxNksuAaUQAzSTyI6RNIp1a2WOAFtWJOzqio2qLcL
4Pftbr12Kjyxz4vQZuPc+eAAmS15CmUgBePoY3Jqi0v50AvvlS7qTeDIhk+xxRJc
Qc9UmjHvE0sGD1Wd1gOJYcLyU/hLkXPkq1gyzIAGfUXa9K60snCBmIjdk4WITPrF
SzIvX0YOO70mwsoQSIPRHyWrj6/nHie0JJ7aKeTmoHYxOrYXDAAwh6Ua99Dy79Fo
PI48UIVK3l8Raht064KzmezruEbThwvd/EtbCzDY14Ym6zIw8Q9BYMszpCE8G54E
p0z+jxof7G3OudcbDRuqsXIpV+worw/QfApEygL13OeIOEOSFNxXd0b4DRy1/bOK
b/Mg179TSFLjbwZ0VF4CeMmwJjAep2/71MFlg53Qn+GvovkWx66dg+7ka1Kuppk1
PvbjvuI6un5pWsgEMvZX/ks+DTbhVGcVrhVVhCeX0Ml6dz6ccxHlGnDrrYe3ADR8
wR8f42fM87+GAs0MbEV7EqqO7d4LKWQyuGdNEIhbBRjnrll4fKJZFy+t7RzIbvrs
NfvWWgO1XAu/wwqYarMrJ0w2JzMq9AG2GUu4Wm8lxeuGXdjq9XktzVeDmrnt2O3q
HUx+NCQdatWVvpdLrV9FTTC0zF/PShO2I2AHWLi3DbLF71JZK2w4rrbLExVVHtDX
NlCWlXRjOSPjC0hZQPoEYtcf/5qOZIGx2OzA8Mj6OSD/B9Ys5km3ECPSQ7qzNxh2
mbAAcD77GE83TgmolQa5FaFficmlCNs3YGfeWUf9LFz7jYvFMA8IZ/UOzOlE3URn
+NF5+cT/DhbUQuezT+AjxaQDWHJ5i8AN2FKbUp70COpjrGZBSj0TBvoYpaKWfTR4
9kVDlJjV1ynrqnYIHotWCLc9aJkxV9CpVSgJMVVDu2g8uGH9HWN/ipRZk9gcwQfL
XsB//QbsS0hRziEWYunnnIhqoKS7eqv7+p1+PYOWMbg1IWWApbnBglOt5TlIK5lu
uRW1pWDRJUSAqKyiJnc5h3rsRNT/EAoSTin4271Ma8n/RJ/6+9u5Km1SbXS1g7XM
NnEy7hWLU3SUoX36ljKn3eWYL8VdPtkv5X70IwICeIIhQUd+PfJk8Gt37OgJgjwg
wi7FTGIHohAHYMuh3oNolqAts90ixyNaM5zQcgRC8e7UIx5NrdnH6FkfUyen6XYH
hsuPJTBAvtFw/Oc2mtgDocMPGGdtvmHgvHIKOiCQJmkZpcG0C0zKgNuVKmx4j+an
L4NLitWGF7ZQmLUMhisR5Eg2ytpQrG5iOl41gJZrnHq5JWjPfJJ165eoQnpErg36
LqZOgH5MnT+JjJBzitl89fkpO2+DcGnRKVdoBUxh5F8bkOdFQ57NfHBfyS8KR4QQ
2h60dzNZoJ3r6Rv5ZrfxOUjE1fUW3F0RcbmiSri0YExtBDFNpDq6ng5LOmmZ2n16
ptb1HxL9vuLzRlblL7IgHbN1CHmqLYhvRfZ2K9qroDY/7iA/lK8yYc0OuP/OKYIh
xKIoJjlBP4b59Cs1NZwdjD82TU9QajhB2uDc8uGv54AAKIp3hoDIl6pFV7XJcBF4
5rX7uLgBSeVuiJ4vkNsvZ2EA67Pj51PFcZzko/oPXG09Zcj+bLTaViOtVR6nmNnx
tUUj/Qu4KI3qNIpieLRa7IOPK7+f7t6nj5CBySuxtwvJ8yL1iy2AR9Yh69UZ81ID
+UH9XIKPXdi3QUfHYdTxmaVuoYhOkWxp4NUFazlq3+Qp+nZL3BEBfm5l7CrwYROr
D0amTG+KGmfxvC91GRGfgMu6yPKb1pK7hKfxAsIw6skOBn8u0Cy1ktCdBP8ux751
Qng5DL8j2k0CNyPAwY5vxR1dMk7r2PjUBA9BoGnq6Lkew8JXVLC4ame6I6r1oLgE
lPPH+pXzhuHIPuwbCQPUbLLrXbUS1wiG2pFOccg2Tr7kxqUD61k+9IrgXFYZ53Ye
Dv2n4GagcKbuVKttuNwhurhRltV/y5CuBaCLhJvRZGwKJZrRjp3Fy0pUTTT/4mxs
3qmkspsAkV2koi/5RZMFQWZEppB8W296YmXDE22gh20yR2jcQrRH9GuKQUO+tPZk
R+b1LDUp2ffvqez9NyChQfUf6jITrZph4HxQTEHZHKQH3hM9hH8jTi576ouZEXC9
xIG8YUuG2mbd91IanFLkvB2VrPMln/A8pWL78s1qAU24JO3DRI5k1/FW8AuozVUc
ksp2w8NTQLCIHE7AGiaX6PaaIleg8FcS1vobhF7X8ncXOJQB2KvFmV3Jt3GuAl1h
5oo9tkk1udxyWa3Tj/yB/h4Me2HITPyqKl4zXtKwR99YkQUaJrdS+pvooqKoT84k
3uaY1KhTuE1o0E5iB1Ob1F+JhOeoGr/eV18pIZIwVQa8bPoVqcpo1qK8TE1tIYIp
SLkkGv6VAEK6Ml3uOrE4n6o06VMa1mJemQBpkG7oZqQw+gfC+ObKaLtPOZ45PlAb
DQJS4Pb2Wi9HQnwJ6Hnc6niJCZ8ll1aGNx790rotEoBJYqLsHkwxsy+BzoVfCslB
SdFFyk6dx08Bk810s2b8Zyzn8PHTQ3UqKQ9lO+zM9xFoTGMatsCnYWgBJjZ922MS
nujVfyCLw7nogtj9Yun8fIM59YClhHPpDP7GmLDcWh8pBLia0rLdyJRyF33myMHq
qU4yA8Vk0iciJrsmRoUuOgN2XJa/ONKD2UYI4Jnoe/eZ9x0ubYSulRKq7lIyAlco
Wj9L9MHqMB0jI8q7EIRSNhCiskqyVN0YktLtDeznasrWRd/3lXjUmLbAa4CYer+9
HcPOsTnQFvCf0n3t6Nkgfb6Ffs6m6lm9OLZmFt23gDtYuhEUFejPHQH6XtPL9NeK
tLTqcve4jz+p4xZcIzSW6xTOdfpji24igqWnVgV3ojN8iTEzEqIG3B+FGAIyuG5/
HLBsA6jC2GZUN88ZrpPnBEvh1rCHrxdfkhz19sQB9nylth+ZbGFmgTzsqOrw19Pn
8g0mVrW4Co6lB9qS5w3W/4ZZrwhuxunMBMi5wMhFW5Il3XNQ4GX4teI9oqxkS3gi
wT7jxw3wTPlYNfIKsL/XXXz+/arIEejBxMjPuadnkZFuYvz55jBbtt/3FwVYCbTs
MnNjyeXBnkcFssxZfIWyyQLORSIbnBM00G1q+zNcprGc6KLcP0YZoBQIozvZ2U+H
v+CDOkcmFvg7P5j41yCGFtW7eRXsTslmj+toMHaMwaCQn654sBSrhq15RvkifhJI
mvpw0mLTG7Tl6bShay7lTq1l/1clEG7OY/Vbki6T1UQt0gEgCuU5nEKjMIIAn4fA
e0MgXhvvPGQasGlsgSWRhoOk5+NLEzltxl8J20Ae9lLfv2FbNTypMVFyFwlynXiQ
gOZf1IECz8BcXDFmjpxlDNiXXYGhPLFldKLx1eJQb7bmopHabJLpCzssML3Fo6NB
yHAn7vQEqrlK/LJq8YiG3MJIweS5i0WUy5XTKYNFfmYTtrPlTHhlpLlYCR+/QR/X
4aUXC0DlVDVeq9AMOTCncxQXoPqJ5oF4xCG222aJ/BJ9OPbUJCzP1notsfya78Hl
dl4IMSo1CNa85ktcDEUbLqMXO8o1Sd8xMCSjSCLLWthrAfE5YgXv/3NcPl0lrywv
l3ix2SNaI2Q/sboNYFQg/T2WJ/ysrgazsjz+0B9YogJNI0kdo72oCHHh0lZ3Ke5z
jdI5Z15NUYTc+5SVtKIZR8GX6o2+zA7m/KERMzfyqTNjdKhq8185yZLQRGXB+9YU
H+e04daVDnC6mawUiD5JhWwbwCX6KwY/BBQgkoWKMo2L/s89p0loKIY7+Y/E4W9y
bJZKe4YzY0n5mxYkqSeuL4C1UoJKIDxQMMl9JpNCAT/x3jm9l/fzxY11K10nald3
6nDAmkU+ayEFC9FjpItTzR04JtB8p+MZ7iKHj3UpzSIaLvD1dBMNiWU+xatdVDsq
ATEu55slq9IyWIs5fvjhZeKGFDOsyb2FOmO+n2aX++WricfYDb52Fh8qFoPdfGxQ
/yxzLVp5/xL5m+wJ/jVMSaIWAObo8oQcj8EJc0SUjNqidMAFBxQVJo8eD6nrYa0X
TykusRYw2iVgZICuOM4EJY93fWwJ+8KZTtkxHc1DWomqqu8l4W3ArtC9jyxG6Z7r
Ae3uCGBQXbB3pB1kxHR5Z++aEsbeTadtKsvWYADVESlXmBzm6tST2ziCTkYQYVHI
IF8ARx67dPohaKmnO0vxJ7Q8QJF6HZejxczvvojRTxvzxZNlvunTCSZtLPyt2D1R
BXLHE2kc2HSr0SpsBu8L7nUOSkRRu7KOWO5hmngRukUdk0jgkhDWQnjFVBMrKM/x
CANdn68l+8W8orUJu+3Y+DXsc/bC4fs3S7n/WmkfuQtLyPsmfp8o+wCBoNOv1KK1
kE7j/htD7qGcf0gMWiifuoQvCR5K/Rzj8QjCyz9uhEFu1fsRNmqHDuP8EGM/ee6W
f3nF5DFJmMIpwVBO5lky077DZXzphIEjQOAolo45gr4gXmA1ojHVemQubo4TH9+Z
ucGgI4cTh0Dl9KwMwvZEyBwXwQTg8d2nD9CuOSpGBQyg3oJqfMHE9z4rRFZv5/QC
avg+eAM7zGOQleZmvRwsW1PDXUhrWplMkW649YLnWVliwqQjrvn9TzVEz0K1qXLT
ONQwE0dgDX0llwBGaoqVrcbnnG3GD6AoW1CkBfZQXLF/lAW9PKsouu1HFUfsbHUo
WwFh31pfJXORUSO/b5NmpAgVpoebwQBNFZ3hekdZmTa4SifXVvYPbpEEweHaSvXl
YjILy7H1KyQ+BJ9oupNfClQ7Q4BDa5QBn+Jn9IyfkQ6EawCkwKdnQkVdNjzePfFg
aXxiMNXnsQQ/3Z7PzbWXXTuSOuTycrCdIwJmmuM6u43fDhO/xR6QOKNa+RCQoXPr
QYQgpnltJmBBq0gUe+A8P0xN44ffCX/zQhV7775kkigJ7d5VnvHorvR/67AFP4HR
N8ZcZ/gzwRh75lLVKQryD539ycmYLKdTOF5JitYn7CeE7rMjX+KGJRFRk/cEQUkZ
9jV4NhTVe5n0p+BZvpSX4YGnYaJJnWYKobfL/FFN3IcMBsBsznZqpKPv8ED2Dy9I
OP6jGEPU2LJWqNJ4RgB6jv05JRR+7UlNW1U79mqkWEaKo2PH71MOuMDGSF4n5ui1
UDU+tDRgP/DwvyVY1jgcyoWuTcDII4ozdg/6dmo0ANs9Ay29CraV6FUtPsB7qRj7
sUb1ytOIoLzNAE0tqsJhKbAFxEIp8gM+o+SnEz/uC+kFSy/nMo82V975VvTzRkgV
8q89RqPnjz+TXGxa+2vJAbdWAaNkuOV/kNoM+qU0pXCabFamWhi3oNO96/LUg+L7
LEeEGLNnOfCu1tz+TpBS7ZCmm8P6qef9fm97XA8JVkHjTOl35Fk7g+8mOicV+zSW
oi//bcBxfr7o762nUuoXFZPeEVZEqrgIIVgl4Synsxmyk8V9g3d7w5Q/QoHtZoDy
Qof9FTS2YnsYyjB+G30iFMXdGgf/sc7QkNJogPy44+96RiDTaLIgq+K6JpXHF4fR
b0GYndPW9Fiu7SX6cHgxSaUdNaGDCFdsHPGT0SXlwO5+QC17LRdzWEEl2PHARVKw
wsHiiZzGOhdvDvGK8pyXWNdfNgtWe+RnZe3es5Cd340t/n9Wb0T0Jkx2kU+HHZMa
ZQvVJTSI8VldBGSVRY1j1nGSjFIv7k/l+Ac/49HVplOGQYRaz5EHJeiw8cmz2nyw
KuPLP/sP81dkQQkh/lgTKtJqz5aetWcTIBRdaSYpDI8KN72NeLflEhN7ibYEy2GI
bteal9sX3hPC8OuPaVxlWfbK0MX/CtVm+iQqVM+yIir8Zd8O+4ApsIoaCce5XgMM
ceQ2DEdOue4H30ddeiGiwHVrkIu6GjXz+UoW5rOqShLb0/x09Lr8PTi7hLAWh2bD
IoMgnO6HXcIWPhF8wX0jvlNh0EZAR6ad71Z/YuQHKtSxE70HqWIga1C3arxz96rT
MM303qugBqHu3XxD4NYs+k4JfnF8YsFg0dJpks3+HU85GsD4XQVChvUqm7OxzIeL
GoHlZkXcSzzRcnKMatfP2yw9qXYqFaBlqLrM0X5xPRNAxc5rkPNvhqPESmCsE32+
85TWlP79P7prXTf8RorryTEeNhdhj0amfiqQixOeTJkPHsOzVWw7JJI+wsu+p+vE
JS7oHDqaH7Xrf83eOPDOgVP+5iwl0VVOCJEOQvj32ys5F2/zP3CR8cVdN+CSWjmk
CRrFzZJY8GDyCAzMOvh+SXGATTo8oivTWgZZiQ+9fHnO0rw8P3DuEhwQsuyXEGx9
je8lj4G8mNb1Cy1tH0iK+uIC6d8F0ehJ6cEl4iksbn7x9dcL08pZUE5OfhDtE+0B
tNmsUaEv6D2hYbfwo5AVkPfN2934KT56RI6lqXfgJACj27h6wMSczfITh0kujYAX
cwNaIkVJbqbwaNm5RvSUOkQ8Fbt3i4GmNaksF5wQHwMvVUrw32MiB+YIoD0vNSs0
MubY8Ctcx+csFXzpZxIIr368mIwb73EyFxLf57/IEZn80JTixZ1Srl6jrprbpch7
6l64Ary9DXcg4klO97G1Rfae/txgfXlh7t9r+gZnJHYF/6xa5cXBETgxm4fuaMwn
pUTpLV8l4Miq5Ohr2wdDNlDV/SouWo/yyRh+lrieebqGyJNBJDWgfD5T+CYUUxBr
iSIiF900AxcDQ0pbrLGSg3Rcw4FStqpUdgZBz9ccOz5fMd8gEPWH7fvOCgjrVOkA
ba6wmouzN9AHh8MbXbgbzxGiwYECtgTp81Exr24uJ8mhHahEOe3mSo0SWh5GvPMP
qyDsOnZxUG+UM1DpFhXn3QEwpsj4ZL+bWUzd6my3veAhNu/alNL00A9qhFeVLQKL
f9nATWaY7GfDDYGbZU+WtGV8uGSY5yMSQ0kVPdvZwm714n0os8SUwepbQyJcJ7bb
noQmYP1YL0iTVkNhgXyV23U25h+NZyyLCx+iQth1Ug3ZpIIcgaT2phP1YWMTikBO
KxzJ/NoUTXvQo/nAtSq7LQvc3p53RimSr1iXqdoOcwRFel6XI6bouq5/+XypqaGA
kc2giLBhMyQmGcwYcXyH37uUvflF2GvbVCVz61iT7uVnc8HxnEOwzIl6kBtZM0rl
yD8In2XeTZBCRXbUiLEkUtiBjt2IbNSHZUbHFVIJs2g9Qgt+tcQFo8HP1ZaGgCZw
7i5wJx/IMXtO9EcQ7vXJPjY4SbsZSAghmCHgJZ+thU7fGgOiAH15xOTqutGTsTul
ZsA+qM3dXCfT+p0jaJXESxBoWwJVbuU0MCwZa/HU4XbmZT0CGG3MDXInBdnrN/kv
dbxFpf3SAHvuXCF4f4sIh79EBdOn2IeMo0aat+WTxaL4Mxp3HLuf5jL2Q700ARGC
Y1NEH97hUb3tZZ52QLm0VPgNAzuqn3cmlPrQ6OiGvJL4X0NYv332YY54qtO99A5w
6qmBJfE2L2mOEp131lW2vj9O5ecmCHD+EZ3bkIyRjKbEPMfQ6IP3YofoxT2tJHG3
BjBOwXSlOP4969o5t77vI9qYb8Ja5MzmBiGSlEjMyndzm0pR9VPyJ5cPAumOtMeg
5LXeWL+0UUMR217C7eCgiBw0/mF+1vZxTs/BvuQVAbi9U754hMNO+k8yMZrtaHfV
l5Y0V+l7ma3cz4d2WGwzbheORHHvixp7PTHmRYm8FMR2HX+laebLyd/pEhRdr/UV
PQQkS2pFTo+pAfhbqSm5hrvwSuZ6rD3Crv/aYiD+D9FcgbnVVmMfAms6NlChp2Af
wEi9YyEywW/7kjqfWByRm4fpNvdGrVNMcnyQYH7J9suNuRyydaQLLGCLoWKTkGBH
8yf9Z6djmtPdaQiFcB6BiybNlKG7LTNmRdeELL4q0UYceduAPwuJ7TKO6B7RGt1U
c2S0yj2IHY12g8I34RD8qFPmEYP7yGCmWFrB4r+i3ImLUx64LXBWyuvHSRE9PiGn
270F/zBM0oX2KJ+kSuNCXN46vTEE0KJx5bVPv5osKn5JaSpzi4eZC+gPb6xVm191
TmkuSXe+GN/hptPgn2ISmZaFWr1ZOxMSQ2d9mmAh/krmbFhP/Hs/fLQzsimQ4Iwz
ZHGLagE26Q8YehyIV4dOa82z8R0eXIwkUZrSwlyDSnRZmebHJeBlPTZ7lfoqD06h
/VZN2JKarnTq5tBhI30On8aMoRevaEz8c9p53JDRsuUL8/GL3tmbnMu7JiLivBmV
ddDmvVqK/MHrMdZs0KzGaq2U1PaqDhn0VZi/8V1fZwEmaFK2tA+wRLq4CwuUP75Q
QeiXYG8TOGg1fG8N5g7/8sbLjyFvgqRGNYU2+V6twWvIlEKDu4v8OLvWwUR0FDPs
+mdWfPX8HpdF0CXogS58HM1vqWRwWKY/TzmPILRPWY/8gYhHSOLl0rUfQce/b7WF
eQyA5eYRV9WY6Mr2hUaxt9qRJL160yQCkj+aJ5uyciN/cmDR2fZT6L5wzUq7W8u9
aojbyNR6u7bhri1AkUQs9azMNwaDrjEbxQ/OyWhKMdwdQ3GZFqzYU4TLxDNqFF1o
KCRLqpbIbxdj3LIEvBsHx3joJHBf59FNmgXCayrbXfnhRJKCkG9Z2Zde+3MSO3FW
FwVR1p3HhqpyDBnvbO64jD7ivYGZM9veXXIgKjEEIRhmibbeDQ5emDBwuyE4jaL3
88IK4xiKlyj59aTATdRx2ICO9WiqLE2GpoSx5a159g7n805q7AzOXl9sBOB6DWM3
D8a68g18kGLekKEWxfkXlBzwHxYrrFifkoXQCGU6bfqPFVRqMtVfVFljL6tCemVr
O67KmC9QOjA7PKbxy5+ybi9NdWc997y25T96glHc4U4mxhPn/7bTuksMVFAdamH8
G9mNhI/IOmI/FKuXmQirR28oDTvuMQpj/5R8ZmKxl7734B13crtTPYLj4iq1vkRn
ayiY07zPWXT+Ouu2Q4UlewOlXMYktoctb2H3EBUPC3LyjfiZzQIIq9Ufu9L1c+Bl
+9z1iznXgv1hF9AlvZphjJqHki8GZpkbszc1q7LGpVfwhgbkkEw2JPK/nsOvFfUI
lbspL1SxQ9aZYwttQXb7eHvycvxZj9XBYymlVd9SJ0na1S34qZOzOkdzjO0rxxcF
qhOJPlJZwUi8S5oXqbekSGTR3OEUo0gojJk8QSXVmunpgJoVnfAHYnI9zwkQwahL
3NjC9HeKgVoEZYGbqyki2v2d4eLIJkImic6AGSy2Rc6B+TeAoZXlBleX194EpyM8
6rMFCu2/T3W5hZ7YpUArxSEhPQwGUU5TGCFOGSyngxytWK9phXJlQ7PVmmjwZwqJ
1jr7X4rPC1DHRLNa2iyyhpzUlsFnwtN4pBe+jyFc0pXVnA1qb6v5imZ2ao2lZ/E9
qSpRSma2EzBJmoDrFXfqk7dLVVWGrsdLiwmXfii5OeWZxrPlWqGFkN3HZEM9EvFb
e6HSdWZDTho0fEY4GJZ/vVHVuFPzCtjl9HYbQ25ivvlif7bO+GGWjFX/LMkjaa1N
M8DG2645eP+mDNKZ2gHpIXlT6+V3bZ+Jc4A2l5YPdCpYcXRLMZ+3L8zpeqhtOPB/
tkP8EhCjdmC+nYikS3hCtpfHr10ys380QeZLm8SoHCfpt3QRiOykc6g3y7/3Nmdw
zxMcPhhf+hxRaoRstCnlDerm18lhlIRMTUK86bT+rdAXoJgAUxx9JXGva6WzA2FJ
HdQNnr+R7kil3Hant2Qd3xVaU0iKWl4+kj2YYFip46Sr412L1x+WHLg4zYvzQX7C
ZMSdk6dTmyzwlvPjBXGjTAByoeObQDxaHS3iZawTEOUKURzwppvQfom7hJDuDH1r
60CEi0DvWv2TrM/A4N1y8QxpOCGX+/8DWDK9p6/m63+5EJ27sv3HQTKBjyCx6pRw
/niynj4TVo/WD80eegThAlVP9dIJUHP1XuyvZx4oQbP0R8D6tj7WsC4oHjDE6C8e
tIfq4hpaMQ6WiGnwwryYIHeseCnU6DMnSYK/Gudhv0SDpxk+VetBQZMfUV5aF4zz
67spNOLSd9aKJxUfHd6yg+Kp+ZByQqXIDNz+qxiXeKTLmC7y6V+AKsD96vqg1X+7
h6eN9jb9v/wUNUEoM7gJ+qTescTvcLDT3G3e9BN4Cb7lXEF/OH2E2yXlX2FpDDkj
wfbSHaOwKqPqkXKTGSo/qc3MBIK0yPKEKxD+qdcc3Bwp+vx/4te+wNg/bNa1BHW1
PwUjNE5uMcA94p0woJbNV1YSmvVaGMSiIGLeY3UZmXXMtXFf07+Sjm176CpZY+OS
T1T3j4d8ZhpIXEOoLKtNsmNmOPfOOiiPLKfobymv51TPVU/fzfgaHt9pF12xjMDU
YFfiRCQ+xd73NVdVB4/GaM+i+V8gPYtMKdPt+vsz3yqYngPM3oCHucA8wUA8LCwS
Pe0Sot40oDNzEhuKODc7CUpXb/t8MFcjtIHP5frsMpI0uE5drsbJFpzxbJ0pGAXC
1riEAx6AgLkL95X0IiY9+NVHsdKL1GrheDNFNkrSilRdck5oIf04Cfv0HMlpwk8O
sGgCFRCx+lohGFaoaOemNEuK3+TTPGefFyo3GWP81jNIe7Luw/o/yyLdoE+O4WIA
z0espoAIT60u4OiisW4mUoBL8UZOdDWvO4o1PwUilMbBXe3n/cv/M+VBabIhoUT6
h/wypZ5qG3JjT4ZtZGIQVReiwu3AXzfFzJVR7DGwnvlNQpDNFz0vZMs6x08K9kLA
v1FezLDMgvzMyAikZz5tSXWK0kRRU/WqaO+DCacx6xzf8/nAtTF26wHBFzrinKtF
tlTm7xuNFBAGjf+nkCpZto8BjMyHur39ZnZjaxfUZjUbHfhLAiNlGWNS/0stm+2e
kkGRkTTd/KzWxxPqQ2a7G7p9TxasUkt73UdHDtVM1/DgD540+i0OLOJMA9OqhYkq
tUTWGvSCtL2sR1eHx7bmeIkjzevMwZLkgJQZL7TOix3MJy9P2T01rzroyoik7CmE
VR7XCsDtw2zQPHBOAN9jQgVF3MK6qUTWKllEd/mfzEObZ0VEHp5iEoc+tDCOZyfC
c99dQKEieZtn/fcL805H32rCVnqATzSDSNysJ0Fzr/HmWkt0aXJUnxojQDht4z0T
yfC2iBWiymFW0f6TAZeQjFKcv/BaGaNZ8cvjKHMpSIPD6gaKkpJym0EITLz8MXyR
cX/hwYDRT1y5jzxQY1C6PcBboTrga8qEkyidla/JRTRhOV9bgxWk6uhSVm6fwuke
ryfxXqQmpRnxC1+O8QCM2vmWyPjZYlNAuqvVcj8gxmtSlu0/87Xbk1hhLcBt8jCC
ZyXqmngDGq9nJCP/OZ79re1F/vcifOPvDrqFSdig4YM1KywNPcqwuB/fveqFtH1R
fegBA82xMF2WuUzZmEftfJ4Q/uXM0KR0b0sg9PrC8Yd33DsAzmDGMD6Ryc0Ftfcw
DTPuHBRB3bsUF3XLHXDaEs0IrzSZSFti9di6udukkRK5T3AhRFkw2xaRaxpBd76h
a3lmmHnKBX2OkY++eMeH76hTqkgG/HTNcYbJgbaFewH81RDnQYfAMu489M4tZpox
v3QT6PBatsZIJ4XK7uRl0ZkzoNR7gOPRupv5xlSyqWTnn7H4MBYFOexKs/JffAjp
0l4ujVMXuHSA1rs5KiHgs90LL7qKhIoIOO1RVS13WG84D0+UE68diYwDCF1Ks6Ol
DJDJdb0AtNAsZGfXQ6O36yElbeXRoeWUaNEvB/EUVcHpUGD5MybNtmkzGNO9jPEh
WGuWniocPYBdRSw9O04Wy8Jwi9mrvtmHngLGa3BHgPaMljDLb0DuRBahz1hrmhQv
AsqpbF0wbCFCn11HUZ+N6abwk4Acn+qYHoFHJJyeELQ6NeYofZZJPy2qruKisJh2
/vpirCNcwobJf/AbAhYEev0TLxsG/L57m4pw2rZaoA4XBMbCoIUc04dkV3x8yYix
GDzsAUmrue0hlmJcE4WBww8uFpsFzoM9LjHyAhB7tJdNrGhlWbEoszlaYv0IFEMR
wtbRp18y40lguXfTAQcv8a3SYGmYWOVQTZU7SQBodnBrR5uFenGT4WOCHnOD7qZO
0LqKfZKoazune2v199LI14nUsBi2590+isi67Tis+6tKbsfMIdVR7eqBSOke28o0
PTjlL6eEBdRrnCbdCsMTz9EoGJqwVbnGE2Uusoks75zDLeXIyNC/9NhMReGOwTlE
OXaaYlugnKVIoPmgOzBTxcwE89zk7ieVpD0+R75+9kbB/Gd5i7qGjYu1HwyETHVi
cq0JJmTY2nTHeiQuuB5hpA9pWByCCMtCR+jx/ixKPiGWIdHN3XHJevKJX0i9vL5p
aFQzFfRDSQ42Q3qeIVIwYWCCV51N7O9iwgpaZrrmKn58efROsaqbKA49aPaIN4G7
JFDNWDy8tx9d0xW0SWmmbCNXJkeERuaolSNjbwXpugnA8Kkj6ae12qHkpsj560T3
7IGblysaKgIwCqShaJZKQTkXdd20rz2WkYBQ4GnGNdubP8sohyAokrYXSn6Zh+K7
XGnbQ7mBFSzsqeILzRgt2sO0Hqr6Gz5LO5+SAFBA7wGMfuHLbsVCv6jlfpvRA42O
H2uqAkWiR2Jf9Kivb8V5WcoKMUF80eMBrk4Bp69O+pgLd/F6ROLVwU4i8XyFkH3x
pP7A6p3kP5AuNevQOD98jnyXrhtE3PMWhTS60ZHJPGaIOvSaNyr22HgfdunKSRlk
3hanB/GtPYLTsSms69hMEDGqbTQ+KjiPIDE2ygaYGo0N2kTmqcrNj1+sWiQYi3hp
QATrfUcEkbTHgRfVMOaxkcKTdEzVZAs6ZHdkF+AcLDzrZMta5h1SzhB+ptDCai68
UsgDsKF0f2vcvs2GJSbRhjy9JG4DcqlPLOh1yteYhck2oCsBbk53MciUke72bQkb
L8qhflaTu8xWbfDUZ3RNK0w1AHE5baR6370VQ2u+NaT+RPp3ZB5unYhIM+sw4jfU
X+dyY1anfEZC8PgipgTeaHFWtlNdcgoWRUPyqQPaiJfjktJg37D5EmGbMLEApeQJ
YrX+EuEI+ws5k3/XjUi4buJDGU5BTP82G3Pr86Av5d2NnpItQFZ/LefWqOhqBjNJ
ZtqQwCgTXvWDOoGtoCX6HRX1WAaZeTvL5h2UWQEgcSfCYbxIEQVyKEXeZ3PhpKRL
TCrOXBUCY743CVttPZ44DIJ5CN8w9Ih4Yfjy+PUN9VSDZKLHX1h8mR5ihguebSqx
ZzEcRPjdYu3mRud9U9rIQu/QI8JLTwexwEMT4X5ea5tjonwtkg1AwqcW9OUavWQg
nvhKzzeSXKwOweFlR8YTIVlXBEos4S2gMORxnS6FRlNrUavljM6kwPSLbQYYt7Yn
aMicBPaDmvCvANnEVwvrRdGJVaPWcUlWhIiJQ53r4/iCn89iBWsyao01PX/gzjpM
spxDpmHX9xH+ReVjj7HxNm5wVsKLyWtaErBv6af7WX7cgPbjHmuo3Zbj5IDgARvr
APpsCQgvK/uZsrrOH+ehZ4ZMDh6FiKLWJRCfIdz0gJWfLSBM/9bMVqbAhN/HChsE
EBBFIl72guEV5jh3YuOk/GLoNygBIgrXnlXLNtc9K9t7B502SJJ8knVSu6M7LP+1
K3kJRJG5fwQ1AwGkX6d3o6b/zDQyupngqy7wLbxl4g5KPIh7Q3PlOQAyTMpaaa/w
DwvS/zGdGuH+6oB8oVccuhp5wZWc2MGbIE+hdgozcDioOryoL80sjP1HGNR7e5fT
bknqvW6oWYdwfc2HAlzpG600/E7SxgamCIAlQ0TEIBVT12i5jlNBbfX4sHBw6bY4
Fd0eVxHE8EC+XheM/VwZqZM5IazOB9yYwwH+0FXRwum+SmZvnFV2ezDOZTz9TjIl
lPgyyP8nAaOC5B3pSaQDO/X6NKPcDxMS4CaeHofEg6q92qw6iUvJgegiaA7T+u8W
87KbXP31LEi0JyrXdHVsjhfG/JRj/QHir5EAheNAJxh6IohxEYr8cl7jmfT7dO/d
THGWAylIGrHfLnqj83z/+K0aQ+MzphUdb01x6a4X6va0ag0cOfNWVkAh39rl5flt
YSEUMYVg2ad0oJdPn+3XN9scd1Gx4Gx8tSDGzUigVMRHRAeR1B0PEG/SaLUrgZtD
NjLBvJWmUnnZUMTiTzy8PFiw/dehsNFDF8fcGS0sNjIcI8GZzpfwXglMQ53MNOb3
fn2zsMAPL+6xexPAg/e8WVorkM434TsbTGhNu748QuPKWLPFhEA91NQj1iWdfjxP
nK5czgFjk0V/TWEiFIQrnHHA4wxjkWp6AVKI4LH3sd6f7VFxQOsu9bJloz+G9iwf
Oo8GQoGdb9GREGL9Abj/6VRZ9IcMNFt7neMhI5l53ulSUh52pE6KGeuE04c78F0a
Y0ny2SMbOwNYgEXQGWbS8T0QjEkWCNrd6s5vQFK87HISTUV9elUS9KzfEVV8/nxZ
eUIi3Jw3iVV0TVhbGE88YrOs0MMU+X1cf3/LBQnHaJNmQbYeojOeWy3G8oqbgZ9b
IjoxRd6Ko93zLaYzVgUQNGGVYqZ8gdY+NUHU/V9o71abyPjps1PQ2jLGCsqRlRDt
K2VxOSN3hTydQA8ZjSjoLEPwE95i/MTe3/7WlkBPo2Yp+6O285N+Dsyoz9WX87Sr
4VjDtdOtARhNK47bevFAh0o9yAPPl77q9l3ZOUoU6VKXLLm5ys/dKUOYIXBJjeL5
Y8HlY7z6zqTCS7iVXLcJU+cVml5f7wMiNtU/vzoGTTgGYAmgDQhNs33/4PF+yVJ7
qHUWXpeQO+wqrrPrAoZKQDgiha801DJr4nCEHclxuQ4507Bp0vrb6dJ8OakIaPpD
A0ckFccusmCIDrUWWejq/5XdzD4wVoWWp3eieb3MDiS7n21m+euYyAWpIHXlgdbg
NmWDBXnUfA/mpCiyY/yxgSeH8GSWUvxBNxseBOEAo6nVp2WxpVJTpxB21w8Up92R
UsBxz4V65/Vbk580NqIgcdD7aSZ0MIboXLk28wHWNeCjfvIwol6fxwWbw1gKha48
YehKCSOrXCv52ohYdUvZlH7OVe4ZnlFkVXUR0XVN/Ncb5CvxGWypcEsB3UztBVgm
6euMSVtnO/kCqk98jtxhh75iUHEJ9IyuT1iDWT6KMt97tGo4dQSfGceY59qSc4el
akxCdpU9pkZXYPenZjS0jo8qc36h82XPKLxOXrdEK0Qg95z6MJnl4dzBArUnRrZh
wLfH/cPJNv+rs3RlB0/4XOWdEV8Hjk3NUl5ySgoOt3FaN306uuCe4tBjfDjPPZVc
VzjlMLBOIxEN5afRayZ5mHlnNWPLaQFyXwOZC4pviAQZZ/hNGLVs+f94Hm/2X6BH
hDYe48O1Sgzv7O79cHfUs0kkN+FU2THLbdHfCECfO1XOMr07Yu2C8ZRFsZ6XhRBW
DCH/Jn2nDfiyyC0Cv+MHMDyKtgyhVSoS4MkmFwxbXtl8+44x7J4YhDrHPB//zJV2
Rds0PT1jrkkPqjJXgmZTpADJm5iz8ohYfIzXALBoz373wVL2EXwvBlmrWg1k9yEt
abOt35iMyNIQYUuufN6fsFSt9aIW4qTUFfq2bBEJhkZ+Nr1EDX0TG5N1llbVZVao
ti+yum1oWnX35i8Q6VY1/Gz3qGhKCDAj7SjmlLtZJ/SvO4E5O4nJmEvZT2ne59Di
CHeMLxFvL9u/dl20vS8JrumbPLm72yUD61QbicIMK36I+6UR6D3AVBi3yKCHM45Y
V2941qYMFTTpGFfU6e4Yg3sOE/KShRDFecPciEep1QfcI2I+ilkitd3p4n5BLT1o
B14TOfVMltuCTYrdyEIzMB7mdo3LzAtPhBcF4kEVUampGlHz28psAJqdTDUo+J5z
2YYK9KKYw28YAaaq4/cviImCOAhNLGCsu3XvQJRjaxsROQScUBsthTw8D8hkCJ0A
YVhGZDttyH5bS8JTOf21W5CHOeJzzjFotwzL+4l6ggUW8L4bWk/qYBXnEuOFDWF1
i5FFjlJM131Gjm7YaLryCmqc9DExg2zAVYSzUVbS2bSLGMQ4Ct3GHVrMlkPBAJ5n
C/3lRieDcRTtmwBWyzijP3YtQ73vwMEZ02mFOk7YpHWdP4XnocFGqO0mi2C5seLO
MLbxPAa/XPsHAIHgHunNSOsEoqoPQy7i/k7GBUJY2b4Uk4y7DGklskiCy0KqufXz
5q3nFiyX49cqBzdmbrHM4OxKwTfIsTzzlYLLCFkDRpU2h7EJYByaYDw8kLexBMOv
ADfK2w421FLUcPPYeDb0M4/cM3nyfyynu+swFUacTRBiBLoCKD1IIAYIMLLm2QdR
o5lBAVFdFXQZ4vjxIiMX1Qj/FEFoF+IPW/Pq84eqo2uN33F6y+zOFYmdwJSn9luE
UWMej/Sw/ukU2Q/X3p4qnq0LsBMtUIOlysQf9gRatQyKXKSWJwJSLF8Av+K35fde
1gBVP1qUjDavxahZIZjKc6AMX2DxJDjyNNUz84Od0+eyqOTYBv/mpGzzgx8Eqx47
psLpM87dBbAvTlYr4CwtBQB3vty1K2cFhphORD837SiAV28A3128bT7zrFmv9yKx
wsa4Id/YRZulqKGEzYurCf1/UCsA1+bYGSVEdSH5+bfq83vR14lxTr5RJvIfNDoQ
kDozexT1aPTTByjQCyMUyArz4d0o4ooODlqr7n7VokwyRfA4Iea1XyVy8VFo9P1F
GsC8Yzp+2ce/07r2fiucQf1qguNs/cn0+zIecXCTru8xFi8kxu/VlfBGwwo+WbYI
4oHE1PROzalvZ/4fsp5O1UigR7UbmipPl25sJZa0r4G6Je6Ee1J9evvM59Xtxa3y
qCevldvaKF7UPpaKjpOBOOYJbSp7WufLr0SvzJtpJJOv8kohWTrZ/vVjcNcLp4Or
vthr9onAI69KRGSB2uDUSzMQ4V5bqrBoZUIgBqmtZhpr4/PPATt5u40F3vmrAz8p
riDWiQlfwp1m1mjxrJ4Y+LoSTHCgFK2SqlgnGu4NOblY2B/txtYiHVgHYPs2+l0H
ssweEEe0eLe40GovOZ/tVfbnuo9zEjgsZpJl/MD+z2eiqNn8PJHEU1aIce7Nb9zz
0aR7N40ujELg17ZDUqyablr8rwrm/6dXvBwzGDr3C+qNQ8jJxQaX/jFz/25+4cGF
l5G1PAU630n15c/W7QXNg8wTmeOAzWnNS4B8a4aVzI35TLtCudJVqsjKvcwKKbLO
vsJ4hMUYzwj0OxdFxZS04P6MtaZ5ycrz+9986axyrXcz+JayNAipwqzhaBGvL7Uw
uWnRM2SqjFaT2J6LRozdS+680m2GcAq/v2DCKvG/c1qF6jYKE1WB1HFdOgwplzWG
T6Ml4LEsT7egIfC8AfB2O0EWCfuQJKwDuNF7/YotvJKyk0krtOQl5gd6JRpqbYyD
gIc14ueOlalvvzBfupLKuCJI7NdlSv/EPKqEFx29JMNfslQAiZaV2AZLtvcbjEFr
Bmwho8v6ShCTfk2UuEY0zZcSeUhwCHJ/y2ocbul3p09m3/br3hNDF8FARrYaI0Pd
d4r/myVpgTNyu82Tu59CxOIQYRPgbsfyAzwVmJ4erLlTun0DsdroKjinzekWAznY
kG0oHKfdVLwbb8AFNxOn6eqjB5mhHs5ujeGA7rnXTTVQ9P0dixVQqwVlcy7CsQVE
h7vGTgf2gp1kz8hfLG1jLrk6A3dL0gFn/xbC9jYxuDB+vkFAwa3iw6I750RgBjU0
ndXZXroL0Mp+CwHDdjpFVLxlaqt8WyDEN8JRoqg+7bRtRsvePY2sHdC7Bscjs3QT
CaoDQVQBs/yCKKwB7mb/u+dW3hWvJxHNhA52xoA8srP0+eSxP/6uNlPlgG7eAuz/
SE7FRiws5zu2zjsWKgR/M+e9GsfP/F+zuNdX44eIWcU+gMExFZUhxu4UUZ3hRfpk
6ptzw0l4/iIDEbDN3/9PLQkyMhR2KQ9oGS9otzvUKdaLvPhoUscTPpLHiAenA7Yw
6Zb8I4RL63b0/cRk2o8W1szMfAqJ8Rlo/9mvkC1owPmCs29rD2dic4HhLRHq0BH5
nh1Ez+hPNTj0gnAoSjWZDZYaQowyxGJMWJ0ldZhoNHsSc39nIKXYiSjdYLxAyTGK
mXzUta9nsRS/Ra5HGN7SVG2ZnfHkTzTxNZuA24NMMuDG/hPt2q6ofh9HlaQtlG+N
S22Edk0jC4kFrnEqZj5Yh0U77VXD9yxt1DUv9eBSXePyiwqv/AskHPkLZaBPK8+1
ivdymMPE+NAndAvcEGPf5IrC+JRJ045oEpzq4vTPIqi7/3Px3uZDa63yUO6Rwttj
n1TB0m80Ar14WX8kq6Uw//9H3ov/HylV5QrtkAA17iUpiWxH6E8TVGqiqTxXz8Ek
+aasIMABmWMQRmxIKjsPfjCC8Gji6d6t9+sFMaYIuTex/43b+hTlntSJZvwihmJm
nK6KZEHdSwM6vcy0KKrfRSG3fVEGqJ4cliAPE5YNMKJyCyGsGNszsQdh8Sf+ny21
oJ4eGbkWdRnr8DhGXzJiAWxL7nx1Xsgh4EexSi7l1UCryJIelW0F/IkuHq0jDZtm
53KKDgYBUD2CXU5OypcbEcCUUKK2dIMbDU7O7t3QJwjuxiHOosncM1Ige0WJcD3e
6HM1cTYnLzbF6fhvFWv7mvKE3euRuxEmIviKTBS1nN8fV10U2YYty8ThdKstu5Ld
o56OTAnpw0IlJogVESL78wYOdxNeJzGacpGxN5xdc32uJSpo0hrmc1PVU3dPOeBe
kbVpSPF/kFv/ZTPlE69IdesJEdkd324+4MKnlO7LqoQ18PcOvvMIvDx9Ll6tsmYl
gHebHs9NFSPBPWVvcJJ4KVKhlj6EHNRAp7LzSbAQwff+7Xb17E8V7cHBGlINd4an
DrJuI+OOIt7KRO3IDZloYcAUSwhsHIiJ2/g2uDfWeZTXO5DJNFBIm7Syc+t41Xbw
0ArVdJtmU7pqkff+s438FTd0fvLgMpJjQgaVETwk56pgxCSzoW5ZOz1cVln/VifS
k7hySCEcxT5Kxr1hYgBZkASjtNa/fRVG7qrTLIkUk6pDGmF340HKUNaSyiVuvH+K
PgE3Pp0hIIHdo3sjRxh84NyXdINSvu1GbtXgTeGLtwe/CtRWZInZHOkI8S4eOVps
eIaed2PJnIC6spb975tm65g104HoUQT8i8yPAKf5fGTssEv/MnqffV98raMTdyk7
IwBU7NXC6PD0wuMKyWBAH8gWNqvGbzp620JTLO8gbm/E7serM2oTeNZBoevAEbS8
k1QuFnE2Qd4Ao5XgFrKfmm4JLa6HjIV21nt+8stcVC4U4LSxLWBVyYnvbA+K7sFq
BX/8stah1/KeKsYO7DpyxL0JxMXGgXySWCMNSLBG5iYB8T/bvYjDNWb7juPVcZu5
xYCLRZwm5Jb3wFI0fvZPLI8MGyiaDVjAsBdUPwzQPUfzjZAlNJubnK3NVmyTr98v
FwrsurcjXlmYQKcaWnJFk4m7Myq7ricrCGFlnOrApzn3z+O5fncrY9Iy2lHM2iWN
n4IgVXkSKNfW44sGfIzXaVpYptmuO7JnrC16REgOhVjm/0Z5dGhEcgOdSfb6foQj
FyCFiFAgWXB/Zwr5ZBqzPPJnrPNA1FcdaFI1/CThJhBFmbL8+VCZx+E4ogz7KIht
XGt32a8r3Ul/RylJPB5uA+w0wcQvVo4hbCccHN60lEwzju/0+4+q515GNcl29E7N
wROSIGfKJn2C9npVPrALicQe3BsVKjlkvxqR/s8s34nTIkN721SWg0WB5CvPqfrL
RZJV/FpgKb5CVe7AwtuRuqPcJn6PyOwt8LoDJ6ijli7MaFtIU6ojOEkeWdr/P0Nr
mTAdTwTz+glVSPyfKHmGq9ic31owZz+ePjItwpk6DvpPKyhWAZ7i73LTZWDnBgoV
pq1nCrb8nDDvonEkkTPDwHcOzmTau8GYb0Lh+4KvXdc8flgtKhZJP+ZOOfLlyGfk
C7mb99u+TST9Iovu8Y7lGEueAash60syBO5JiBIew5Bld5VGjrHGaoW5QaZ/zWsG
tf4ehiuJHUAR6HMBS92XHJhCBO5CDHSJPLVGMvqoEgWTqO3aqpolZJD75JajfPJU
ygDg64bEEojuDkeirSVZmOxVEFiO+SoXCK/JswUStkjpg/QtouaeKJTBZsdO9R1W
nCVsW+2mwXTJSIWYJbhr/GSKXMtktpyXuDAAL0smqkYc37ZhGL9s08eME+BT3QGF
mWf3+mNN404RTAeOc0YtJ8+/hyfHsZxlAg3Cjnd+Zv8F+0iqIHY4aWiCfSe4Pfe9
pL2bNsF4FQSDbY+spINqNMMkK5pNe0DR7F1nURpB7M/Yqf6t0eLtlLN+grzBKmRS
ZvPmdOCbHXJXpEVZnq1VTi2lm0UWbdeyyPKsSSDM5HIVUKgvUQluAi5cHxHzZIs+
6rwrJWxm1bjOMhkbxgq47247dTV2Gc5lCDnBMO3qn+sBrUJhCciWGgVT+d+9cusA
/1jo/Wd4ZR89HuRHKkB+/J7tj1FSKxKne9T+3fflJvQxkmaYwLj/KLndQwtWpIXI
nAyONQPo3mz6l1TywqKuT1LjLF/ZqVlXx/wwC/+defwOvHuDHxhDSpJfWljGchKd
prXR8fv1R15e5RCl9KP9TeRXk3Q46QNIZJVgtyTtdcoxcaWsDVw4eIvZMI8lNTDp
yOxj5jHN8HonJgog9m9oE0zOZV5b0aa2oegFa6ThK6aUfxhZrcemPJY0x504YP64
S4Ugt39zNjJ3TarxOq8gUiNoRrPsNHBGLTPaNdiyCLkpyuKeN5lzNAUr3flW5N5d
TwfuI11VwiiAx2wbNe74llKlgRGXbHHymp4UUl++m2Cdq8paL0ta+E1JxoulqLk2
XTXq4GKzHStcwZiN+OXnKExi9FjOIt1gRotH4KfP9LvUBTLpheiYUG6MvNVR0BJ1
w9GOz/xiM0FAUrxsg54tOkohbUiMGUY7pq4XIPQ9J7F4Y0qAli66yyd/oa/y55T0
rJsvOxg99KJFupqL42CZBzS1xNTK/O4mnoAfVDThSI2OZz143aCeoAtBK5V5sLna
A+o+dD12AWtkHoqEYRvYTfQUUT/MuORQpzjN6OUq+hObNnscWE7CNUB21BHlNWam
CwWTJPBU5UXZeB9TogskpAY9fVUOTeZFqLHsg4GvnavwUHuIPhZ7o6Q5gQT7gU5A
/KotR+pnS2l3H6t3dbe7R8JEHyZIrN4U3GFO+WXqb+8Ux6dhUp/dVjyxKjsYhWTU
cq4sgGh0ueqomqq+SGKvqlO5QsucNkkw80yHaNZQpmZZ6Db1l5fqPFxgd2CqUba1
wlA/TjoXkV4RZKTVieJ7zqBuIMW+MIHJHzb2bAoz1zKq1WJpMUFe9gm7k7zqq4Tm
mJHPnRlRk7EohDAHqmzMi63E1D6a05i+xfjqyhOLjp8uykgdznPk/pEwXjyQdMeU
P83mPYy6LLmCjLxJLu8etAObTxXLqUJubH3tG+2+Wv4kCEfTvKavxSY7dSJtU1aC
4UMy0j/1yFSd6wazul6jGkJLqfOU7ny8jJF3DvOCTESsX3LiRQ1ml6bN3s71NyuP
qlvnUVl+mqLz0Sjs3y+7sFZ7neabcgu6QtHCM1QRMmYVRD08qDDahP/7tUUT3+ON
r06E/phf4iWOCU8+4W/ogCzGBWqXlAb9stuEk0Okavw8DzV9JtV4Q04hLsgnYbBL
1InroWAwFgUmBXYBtDTUZAmyoVTZM16LFWQobWHGxMJTrIwn9BK9+yHHCHf72TWU
sEa96xOANrh4ejGDPrsoOyPu+4iksj8b7xBDemeKi3PqVbOFOO/WdrKGVuNwEyBG
b0uv6F34zoDwDfnD7tDMF3ZkfiFfeO7eH3L51gMbWqtt9HFd7GFNrMVBbaG59aPN
ELvPs04oKJu7yHKU2qqs3bWZWg03vIacdjjPqnLeaG7hItXO8JSkiznBydMU8Gl7
7bsBWo0eaRTzpA9MvePtUZfDOp/ZgvHCHC5KEQCt6dZ2oelqj6Z3LmMImtm1atc5
ZGZahwkQ7XaNGKx3VO4N/e1v1AknCO44LB3BnkCM+859ZkIbfRytttegoRGedTkg
F4qzl9buGuZVeV9xuZmlj8G1D43goOVWSM9F46lLq0v6b+fBl/t9vcUNrbdbDtMz
4woxkmy2KfFEfmV3JBlZeSyioFu6O/T7Wi949A7xRzYS+ocjKcSwUKL/n4s3IBsM
uFlQVFsL6iisAxOOTMK/63t0eO423p9d0JJn/VQ6PQfxzHlSjPIk7gp/X9CSBoth
0Hc5lr0Cm86uTrKCc7qNtvRzyB8fkSfRHTdU5s24H/RyiHL1XKobaDhM6v3CAF+q
7WtoVNh6kVZ84fdepOAzr1BZeL4Xv8EDv5ndsTYkAAcKb+j8dBIujC8YKhFiRZ8K
qVKmPX2a04rNuZzFGafucGw4FxJlZ+ta3+gJK1jTkssEZoqKPecgI+Wt7dbZuci0
Qqp6A8y2MeeroSrw1xlia2g87wm7bBZNyhU7XiRIDU6Duz0SU0I6stRaDl+8DBn9
tjfdaHz1Ux5oT725IAIrXHOztHjATD0qh4DhcGiaLCi8dzhOLYnuOx3IOXs12sj8
DLVr/QdRTyGFUOb1kkU6MI39E/jlFRwvcJhW4bvydd5dHeQWyzzqvk++i68Q+azh
s37ZNCFYl+FxhGgoYdm42GZUPJ6fBhM6CEOF2V5pGZewpG2WG0xsNAaxgWRYvP10
Ie7HbzjluygP7zwKraCP40KEDQoMWO6g2l7dgc8cIn5taUTeC2IAVnHA2f9k0ntZ
Dm+v0gzf/TLDOLqEcK+2SlWDCsJ3qNOdfY/8n2qlEx2LmYW8KpxoUaf6U87fHQsv
x4nak4r09YUIWSb8b6ro0syZFBWtM2qcrjYWsksOaqJYXB1lEZ821NqyGihYE7Lw
ZGb1cqTQFW6HDYFIGhBihlEQXfOgL5OUXnsUMacQtZDrSIsLePH56umf40urz26v
F67zUNiwUFqzsCmhKgbBO5BgZpxvFkgvX327huLChFyK59/aZuh2AJJqWrAbY3Wy
Y9ClfkWvxZ4WHcTuMT9RhIH9312zS9JQnz7DeGxfyDOF58GhQw4hfOSQxXPh6gTk
3wcjirX6M8OhpWEHiH/gmcR359mFNnW6z+396CZMKGz15xqqAO6YMdb7ax5Byn/X
QWvKkh6YszeJIHgWoEwfCNbcTGrSZ2YnNkZndJFsqqNPyaVeA8BIFL55zM9SIpGX
ADygLVaLBJGf+LNVyvWqUp2zw18RWqnvSC1wJnrAQ1J/bNdYzctsnfXEymOF2D4X
/3W22Dykv78exYXhmQwL/Z47oT1zp7rme0vvLS8Oe4DzLnsSh4A3KyhBFdoAuEAS
HGmXWib0fVOR9G1fugA7W8FUa2pg2XYnl+qrZqeOdJAI0MOVFBGGflURvEQQxjzi
WxyLb4OQi26iHvlwsy53wJFHYjEXlf1WFO84wvigXZ8jB2gotff0Mh6aQZgWHSgC
tkYwd7XfqE7rORKZyCaoEVMR6bwZt/8ZV4Q5LEOKuM4lijm8umu/fTavWWvjlXMv
Z8ytTR9umPWg5FBeTIap8vLAC5p+7zPWgvqVao/VMygTPgw4ApAIynRQFxa+o9W4
Ij2OSQRWz209tQv/8NN+XOD6KDzBWRAlqhQsZK5NtjvO7eOIl87kWokU6QXpG6Ol
C81192Dy9vMEL11bUIkk+iPkb4SaPmVYs6ZS4NaiVNZ0jOdZrba6I3y2lWCqsVzC
Ov/wBAprmvJW/rTldD19YX+aPzNy0Xkh5LuUWsNChwVDsWQYY1+Xg48b6xztvBlG
LGbckukz1HtOHNR2AmlegSGQgnOdV4Cd5efH/1NvuhMdb8Wzn/dV3fuW7mo4jGZG
PSSVy7TFUuRMgjXPYKMWZvDCgxt617D/U5/473dDAtMnXGb+zbmZFBCODT+CbiRi
cN4xdtT/zIzL76EKSwrmNL1wntP1waLASVeGyZQn/uADzBd85lnGGKX72nW0fG8K
WkqElaMVFlf1qVeOR/wtjraxNWfZJoU7LEUszF+tiNHkPR7WGwLHj8puiok0Tfhu
8RHM5qfBkPGWDFYkHIaPG3xmSlzxrCFPWXEu1g/LGgi5VtEaaPbfRRSIOoTvnKhH
0IWBTLtucl3rbUaUl7RXgcONdAdOvbhxHmwCLWKPQeGR5dEB0OhrYF9TFfecggMM
xGP0pzpcueuU9F92DFV4PsPlfFgTKsfmHCUuaLYB0VrbqrFm4hNPmwCBqyOQD+Kq
tFECWQjjI3kmgCeEt68UM1QnGhCQbfHnaJ1FVoWmtZjfKtqHMXqK38WAjYn4ezZc
o2k5pCiGq8UfbldCAXtnvjwduBL5q63jo8skKp08UG/S/WMZcFEa73qt0jEfTZ7p
XmaiS6B/dsrktRRTh+/tdFfebb2Ui+Nznp1zXq0C7bE4I4hxhrvUWXrPIUOJIuFT
/BFv25XFRFDY080h3BQ6MC/aH2hlpWWxcDd9syLDhUMtMcqUtLKhN+DAzFTOpxM4
AljV88gxwUOPvD1C3SwUpEluojdNyRHW35EYr8X3Lmec0gm1jfQmmcD3lr9WP5Us
9HCC6sUpj1fVuhiMDS4xxRWzxDUfFJF9NGOUaNZ3XcGPwljClPIi+D7brQeApChj
lf0uCi7R9qWR2vIPF2ogOYA4+C65cHP7fafgjZr/OcIYPVt0HOEMR0wfVO2O4zbz
hd1Jng/iAAcLJshvWkeqERd7BPED9wPHO72lt1zIVfAXuysS/CS94GWS4S9pheRd
ZIl7lnY/yOKke/SChMs7uqiEwmzkdMIiWmg9SD/KvshoIVqaZUVN6a6ox1eLosYI
mbhUbUi8IadyPuYzglbxIOFyGCxzwVNuOOLVJqlpOEtyzI8EnUL7MmdMupgufuJd
A8GCWnKie10d20ZiGc9pXyIkEhfxR5/KMpYgTLDDyI2drUbZm2GnuOLttO0sSX+D
n23Ke1CKxs42pvb8Xyif5yM2SMvhyNmSxmatqYZneJ5jlQaLCI/oyN/L3FKfsN8o
bDfrF8lmb4cjloZc6EFKazvzRHe5LxTD3B4tKGIiX/BsafS1REq1+jvE7g1yYpHh
hEOyriT+KertKDGN31CBeCmLSlR8c0//BQWYueABnWjm7pPXamVJCp0t0tPUW8rg
aL4WtA4Ll4X5GcIcr1yy/gSYONo2Yu1cqevSJQ239+BX66J71ukwRjh+7vAoLU1e
tj5tbCCXmmpe3OIEDYglJbsMBAI5Reuks7akQEpx2JVEbyD53YqkOoagLXocM67l
Kk64Gi8HUqozK8jCcqSXy571791Pz6DFVeD4252w8b2xXlChWSNpaS42aMg6iF39
0oky6ZgRU8mlux3ZWwRLitjuaAJP0alwolIxzcXm5C9HiTd5pk2ORsYIF1qMNGz6
csYSWBfs5lb+5cqFy01RYAO3HiS6wnj47YrNzWy/GHTOcpetHPhpl1C2aH24LPfV
yBTqTRBEV2wTE5gBzlxake6McgWnHZmHzsAW0rG2MH5qECEGHlLUAaTG3RrHwJCl
Kkn75VfM9kvQCdI9ImrEYr2LF2tFRPDMWwN2vhTJ7JAvE8crZdOLA1bPOEPfiYNy
n4/hz+7c7T2E7pEWDEcyPGj/B+Ywgh9y7q3InaRqQAkb3klQiUpcRHqktQotQdlh
zysVKki+RrbAildgv6mRIBqG2iJdp4clFlS35keBTbFoAA1HOEQlCgQG9qD4nBpM
40e8bIKOR8XB6R5WMSmoeO3v8BWsiMZciw7ZaBkbnMO7/aAEcRs32vNv4wJaQwaA
u9ve/RIYEETIrEagPx4Ji0sPB2dWDsfsCXJwVqcIQO1DjI+jbCf00/8JKeg32vOz
KWrPKJFeDoKuzPWUqP4Wn101h1CarbUWcuZ2AmgyULRx9xuXiDzSgfZCCxYc+4mW
SIA0OjlKX9Tqv/uRoW0XgpIN25canQuktfo92oV15no4k+c9fjL2oQYXnb7EFyzm
qe3oc+fQLCpZerRywi48WtcozP9LD7i1qUVWN6eZYFeDWwNyw2xAcqq0XoZ4BXEG
EimVHFsNZgyS3xusLywBtoIOIeaipYNRWasrJM9JdJP4F6pgTS6fCWwELzWpHzmm
Ce5DI8uMexpGfo1qXUsbmO1hYuTSjvTRB1o7WCX9HjiPYwcwjvP+CEQbvGiM3sqZ
74183I4ZX65A38n0CUXLOFzMswhVDx0DtCgbLFtW+gyLulpSBpIgoRTGT17KOUPP
z9n+8RcbwnsvdFmuNVz2IV7DdSEJNmAJpx04E5izM6F1c958ujaFA4YmWBKpvURB
ziw5ohXFjiuHAqPQ5zFSW9N0CrtpWYSG0zftuXmqWMypiILEf27gIWkgGui41pye
s303RY7zMYpHeDLaSM9IG4eo1vZptcxV/FydDNWISaABM6yEZWfBGDexhWsc2nqT
XAPoGgMAY7L7ODZTCLy7UBNyo8DUaaKz0b768zXwF+/phjELXgYvAa466mHE+94p
DS1TIDWXr9eHZJt5aHV3/HzlkePsG00L72CaorgCqPasxG4acMCLjeW01ew/kOWl
KGr7mO/lZrf2wJYTwMh2N3YVvntwsABgrYUd4c+2qH4eR9/t1zjZ0wFchr4/MLUy
unaOfKQB7ghiYTpwumvKNat5Kw2paNSFKTckCydoa4V8KSkGG45gjpvlWUlyuo0U
LZXBelU+qxF/gvmcwsYQaOhYMhQ2135bWhU0E2NKWuoYuZjh/Q2C3a66bFvYOA7U
Tc1Ee9JeQMU3J2W62CrwWA==
//pragma protect end_data_block
//pragma protect digest_block
wh1VvlpO0ZNZdIXHG15wfT4ir4E=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Jey0dsd6IiGI3v6bi5DqzVaehyt3iyre8XkG+fORxb3dmiOan6+xPffEaW2uufVy
elAoymyw+zmifc14dJhI8552GNojNrrUpEqdeDXHM4QbXrJaEd6b35Lvubvq1Ve5
nRKbZOyk5edloEzSfrVgIdAuQ4Rux2L3A+ub8hl5l/8myUhyfPq9NQ==
//pragma protect end_key_block
//pragma protect digest_block
fTzuY4xTuSRe2bWJKKb+XQhSPxg=
//pragma protect end_digest_block
//pragma protect data_block
be6ytsDF14OuB3SeEB65ImCAq0EBN4A9zuxbmVVM5TCIWnXRTmQOMGLKgkDjVoKG
4O/UBSNdMSGcc234MypY3ykJyvC549s60E0KGMPPcrXkAPy6OmN9VVXuDXHiOq6s
35TR4cjWkJZTSXG5oggXGg/VvAHjeHDx9HZ0Awb2Hsj9njPdUkRxnIOCPl/nxJMp
V46LnpBraPIu0TTr6oNFEusjMmLbdmx/L72Sn1rGTpBvGcQVtquRgkZmETkC8yI4
ziM5jIKYNR/v8+R10wE7odRrHbu7e3tS8uf6F9zn2EZVCt3dTIEPH+m7hQ1FaTMF
BVdnNWbCr+CkYBliUZtl0u05vxwGZqlmdNwSq+WX/XGnjDBWe6+0HH6ylWuUMEMB
SntFqTvxliyuS5dDkCrKj8KlFTFFN6baXtdsGVJ1g1bT5sEQNeMsSZCIJR3Wp0mg
Vkf1GJPnZ4w3ONcLHKx7pg==
//pragma protect end_data_block
//pragma protect digest_block
LRtDOJwYa/e0GdpRfw0EP6mgNi8=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
x0u/j8oxXzsGbnzEQxJIG8QUmDrmG0Y2hodRIMXH5NYg0hY5cGlHP4BS+ePruGSc
fxFPEMqNcJPRqMT1E6YCWRhiSevtyxvyP6JOvql1BpaMcKp2wRYZ0uhO7N4ARIOr
9md1IsV4IXAovk0fymkR+QIIcSlv6Y7i3ptdZLDl/hLrm7ZHz1FbWA==
//pragma protect end_key_block
//pragma protect digest_block
9/vHUUilYPlmavI51VVExOn5pkI=
//pragma protect end_digest_block
//pragma protect data_block
ZRPivKj2slJFh4KEVhM48aRcZhTxGItDk1Qc4F/iQW2aK25iTecl5Vv8+NIM4nFR
9XxhZJP/gZPCULNSoAewQtWxxL8o7u4RWVtYKtFR/JFtqoFCVNFSGSf7ZuodBEgI
Lc3esWI49IKMoNIw3+JBrd1e9EhMW56apduCmst2/xG7FjvTXX7mZWRRA6ann9z7
OpUlh4cjnJF01qadS/4/3kkXE8WoYURlmBa3ddBbfnwCONmdgcBgW1WDzDKMYuS3
vt70p53B+5SKMYIKHKQhr3AEO0/OFIvetWAMCT2AEWyuD1iW779oLQFVFr2ux1ZM
u07na/wJkpTRyV97UjDNDc0mYYXl3P5H6FZE3eB5C4EM1AGVQeyyYzyZPIvNVcZB
gxzrq2X5A7FVAnygLYuMNDDEkMancfJIq4OIb/w0dooZ7GNMP/pXgVR86Whu0K+b
LCGWJTpW6oox90V+B4U4FPQo7ClvLcf2Sfdhtio6bQ4wH5VplGPcdMZ/x/9fwqr+
cq6pcNci8OBgH1LV36Hds+RZ6VD5y0PKW3UrciJj5CWy3hFH65wFw+Wtj4YpWmZP
caTL9EiyPCG/LpoH9X5KSNSJho2lPBfEL0To8G7bZmfG12BHqxQg34uHw/AsWfYL
GWzK17YfTWdzOYAzZ8tW6+kGcToc1+4QuJ1UG8MzRY3ty95n6SbbXzhWMI5TCi2J
BZ+7gY5VlLkmkKfiy0b8PBqkptgs7ZFaC2zhm/Nb8hT+IesW0AMHWrpEQDtsGMnC
zRDfOb7yDPWQY16PX8+IcekyP+R+n4JD5exyYOwubY3oVbAopCLyy7bWArYx6BbT
mWSLERzmZ2LdbkK6OFmQHLw5jnpmQ9sFZCOvBYIrLFFRa7pzmcRux8en1JeddhIg
HbwWA2UYBpTDuiLu6MHJzWf44CYAiR3eB+6RZsaFAybRHfoHN76l9CHIr5VmuWQj
3aO36S4LtGYG+KZG4ThPd6ic9J7XRVMYjkgTXi6/0wqbCz1NYoVeIXkbIkF3Crpj
imSqB+IuV57DgC4XseDkYcRCHkyOhJ3AE90ottEu1XBrJJG0aD+sxnMP+7pMaaUk
jdairbybJwyRNj0ITX70vczt3/DJOeL8Nab7lcPrhph2zvMn+ZzDaQNnsgx3UH2q
Bdnt0t/XRDm837ntsEG0Vtfa0Q2UdMIelEo9jVFweZq5XC3MyOrXq3Rp+/VRZwRn
/wmYAu6cg2/DFnQ7G/IijrDaD0K/eBXsLNQegC1VsqeQ6HgNMVjFMEiYKOoSfiMt
HtW+EAH9ZCknuVjYDwExSsy/MAOsMu5lM+W/doIXu0FCoZUc1Hx/REYaU5v3brNQ
pIy0eB3zY2Z8mPWFkHdqYXmhfKcBTCa7tgOo+PVpqTAjBuA0Wx3vx0KR55jNLg13
gozGL7MQL5GdGfxoIfj18KcP58NpVi1mBnR0PwXOWJeq/zkH2rXTqXl+Z9Eyv9Fc
wPIGFdCWCkGlq3CTgQHNSoX5Act6k/ltSr8lzl/Lv/B9dVOnOmzMxyn0iv5gMGZ4
uatTZYygYE253RTKG5a/ofQ02C+oRIKWLp6fLYlLpz1IaNfADdjwI0rf8ljJ10y1
V32WnRpVDRNwMpMJ0PT6Lmak9NdXtkUGx+dg+zbWbenimhLI6f7LTAG8CZZqd/FQ
e4SZ6T07omQ42UUOBGRoEkw8OujHEUZuvoaVI8JOiBrz4sPN5zxHMtpTtWmkEeOF
dQJxSDI6VahCr96O28rnoh3Adci+UhVBegBSlB06UN9gJWfR0BxIKLFV4Qs3MNO3
yKx4j+dxyf0YDnO2toniK0JmtnBmMZBYO60+wHT+YYETEJd8SShzACYb4CQ+9m0b
OoG2GZjtpdOlaZfzeC4fPMjA3GnFum6GELbCCnlLw9QdOFi91ZdKtoIDyWPuXMsn
DMKrzpd2oRs54XxL0eIlPJAM1ddfSZsveXJxMnOcMbxlZfUzxtODtIhRF1ngjTTA
zvuVn/EnvmxiM9flBl0jRmJem0dLSprC97tp7MgNdc6p/Q03XsF5gr8GkIAMmFDc
xG/JbR3BpUZl5EYTYRWzhennLxFPFHKFoS+CfL2wbH90wczn15soTdgDZ2rvfdAe
4O0wQrKMHbUn6Ne85FxovVAxEOSlErs0JOZcdMdun6Afgs8kuqUA/qeAI4j8V37U
C3lTUUcX7d/pIQ3poF/eLq4bclkqgS97AGZNy1TAhCcjso2OcU8Bdijs+JKrRyt0
AL6GOHLrlmJp+4dyb9hfjOSn+cM/9pVOTiYrBHMoJnAg1MC4b5NOwRpNFMHwz+uA
EcgxsuZWNN+3PZQVkEZd8DdjLqt9+Wwiu6T8LwerY4DFf0kibEk1rykguY07B7Qj
bPDjNpfmAqJ06InlFWRiBJ5wuHEY2Lvc4gg2NZk3JPdE+dWqE2N6OmAgaIxPU4wU
TW23JCV6JSk7NHNt8db0IVPXMXPi6Y4qA/hvpTVaKoJug+Ucy3rLfd6tx+tZCnQy
xsTb1EgoD8yiz0nw/7hpqrqGsAwkItRMsyrRRfbRJvzyzlZm3quPotbAnnnE+vnv
WHe65JmY6jE4hx5TJTaddq9Nfjyufp0TLz2ZUQChO1wsP7iFu+AToi1VI/0M58VF
9gFmVKsUf+5hVMIKBUwBe3LQsMUSXCispICZfs+AEIuYouYfJUJtZtycnVnISpEC
hLs7wslOZNUCDBweM6NqeBYU1q0FYmoFs3R/XjJPcN/zLzXdSgfGJXdhLDUBxeuS
R9S4DcVYU0VX/SEFX3473o30rotAXZqlfOYyL4vW8dZ2MeQyjhJCaSkpjlMvgXt3
E8vecnEtqQdrraFlopcdYntqlR+YI2T+dOEKIy/AsRZf/rBfvDL0JxEZMK5z/7hk
kY8ceCyc4isqPzMGAvuCwjLptLOvXZiKP6mclXU/cz9xpja9JQM1iycH+yfh2ku3
8RCm6w6dq+X2FbgZ+ODk8Ig30PXGkU+7/C9tnb8cQTuvohUhIIPDWCwo/noYKVe7
DFpM7ObbuBK7YzsabHSbwLoi830atHXCQcg/sDGQOxd1sTJIRQXdXrpazIxrHaTx
CcEV9KRC0nkpszJpoP3S8Ma3MAVeyVNpm9UqUbt9cTb8Udjz1AHNSnbOHL2nIiW3
26YnysgM+2HaEb7xCCByXf1zYlVltAI2xXv1EgubLgq6fcVTX3NO/lAPtF+D1tYm
GE7Eg9HAXq3kj9C4uJJS1K22a843rX/xfJGi5WBaKcqe39LIsunvrzP+cCuGfyiv
IZnPmhgp5qdTH7HmusxRaSvI9SpgtjbU6G/GI378uxjwUFAeGWTtcdsrTSPz5TwW
aAFMpOGlAFiWybpFO33lOUPh5I+78ZMq/cjmno5GNfVZGj+kp8vCGeLnmrT/G/8v
g2EZSFiHGcjXdbBv6rU6V0Wl4ZD/ME74f4w8b3NqCMI4rCIvOaARfQYXopFlOOlD
4d3xd7kX0XeaEG0fMz91o6fssWL1uamoqf6t8DyOiiK3Fz0ry1raIOtNnzA5eVMI
6AGqkoNvsT5u4eW4H63UeayONSYzchQvIDQJm3pqX+NZqXQJ8+xInsx97mdqpPw4
0/+523lJhJ8vp9NHNA0j8OgweQpyo9fMas7lPUbto6fYeGfGqulnUSO7zOINVgI7
wOnJKnq/lV1Qk3XFxBHsBPSkkNMNdPu7iLne4ClZjrY98aTd0aI/oHTUVG+Az+vM
J2PDcym18rGwsIq7mlEcKx46k+g3v6zjZq5L1nVuPbJxOkHOqedFPJDyVQQci598
dbQqQx1xD6nfn2KT8PwGRtZJn8oykUGBBEXIeifhJYydtSEi4aymD8uCACb7UIut
ALcpLDUtY6gIbgood5bSmxTIpJmgMbQTzqv/DxmXz04M+xHOreCZFIG1z2FVf57H
hpflU1LEIjqfj9BnMvP4XSFEYLH0OlEn3NHcSG2oHNkqAIDiZjhMFIa0WF/PpoKf
mQ5Ec+gEY0nvUEWyjkp8G9aNtQOvzoZE8339BpXDnDzR55qI6j+NJh6VPF/QtI/L
wHHLYZsmogvg6t1+emSFVOS22fHtaGZt5Mbf69DHVP7FJOor1BPY+LOrBAtO5YQr
IocudwgiP0vivo3SE9TDfB2PC+7blUG2gYohPYUZtj0miRrpDGJYJudKNaBrEbpu
+HdJTIT5jDqj4SKV2rGyMRyYh89d6RCwc/gGMrCANTJwAYYnnaD+b6yyxNcWC31r
9z68xQL8rxaCsR7lTmaaCblr4x3kHBpZnT0zPVdI5acR6tA8/Wgy7wIvlm/demrT
kjt+zp8gSucgR6sx6h5kIuJpSOHs8sJm4/5NGnXnZJlWiIUfTC3YbnM1oaqJWjhB
9aBFXcgpLJA2bYUgYIySXiMDcns3TdaP607s/vMAxKvqkM1oiw+aPxuRP8vrNcsj
lDHv8RZBGE9Y197H9lwoz8P6MeEXGTFyMx4m/xNK4tYS/O030hALClT00EGGMbMy
1jcQOyLH866a5FQjxf+3JqtfhGNYo9ARQSbGWquXrk6TlVQoxQNaEJYVSrJAZrFu
2y2ZI6I7pOHaFHsPYgkOD2uA7cncCRGgIKLCq4M2ziUACtYyt0reRH+Ck0FkXxwS
btgCBXiYOt5QctLMIlev3QRfUrBfZFiE4DrrHF3fbsEwkmnezkbepPgeVWYiMKXT
0WoO2jIrppt2zugO7ejw8Rp8/GVlKNpnPFWPhZT1SnRlsOWJk4/fGz5ev1o8GTMo
8zyJ9CZn9jKDvjW7hKO26E3lOuP02tWnROyRoXY0LrmuBqdKl57wP9ZGsysP+Vol
HbxtMo6Pis2cJeG4R/S9jKPjP8s37OzqudNQoaHY8dgPXLxbfmg6ECH9q6UzPQX3
wVl20ieZZvXO/Xu8BboBK2lsuJXpczSFUhXujGRSnxiehPBlMEK9R0rz3gP1MZCh
YvywJioBUHXxsX58NkFahpifFjvUu9/JNOTaddqlrw5Tn8OwkHnmNR7iCtphIM+v
DORwicysIvzACml0Pc1fbB9we9q8AmzNv7DDwyH8c/DlK/PCFx9m1evxtNt8Rx3T
j70knIiF1hIUjWzEUmh58kB1drjkuLbrsBUqjoHiUplbSPr8vaGGVtI54fyKMgdu
Qm7fy4H8pFORCyG1k+c8MExttLvaBpNP0fEbktRd/q91LRJzjj+gl859PoNFI4kY
KG7t4CxFcxFgfshGZowPscus4p7KHtKUwb6h69nIAA/fFWOHQS8lqCyZXLOZCU8R
HE++CEzMk5dGY1htJx61bzbAVhhcCeDONOD1fuF5OIofh1OG9DoTOR/q9KvuS36j
xH4xt4yFb6kyk5382bqR3veGLGFOVKO2QKn6UhAXTd5WIKhKGbf7daxhTkCYAgC1
QhHb4+GSroUM9Ut0RDXBuBsaoBoPYAl6+T35NP1MKKcmB4iCmYPSPuHIUF7juQcE
s7/x2SguQub7Hd6cSnK6Z0BYI5v+luOYDPisRpxtoWRbEvdHzd64SyHwIF7iuDad
fuB+KMtG5d79Lr4viEzMcEHUzlsx+uO9s21Hxt66G5BXKui1H5Q5smuOZ+Z8UKZO
bXk44KKLSBbsmE0c3BZDiUcrqzIkilOmsU/GDdP1mKYbpI6C1acoCy5b59VErQYv
HXkUxY4t7ZDHbgMUF8NUGYF6mcM6DlcS3XH3T8dJVNv0zwr2acTjkCkVEHzN0JsA
RsED9jyqowQixocLO5NkB0WehAdiqGfh40F/7X9WfWdjWQQkPRL6uv7vS8ffvRT1
hmpW88DOgFaw2Wv8+fP0OcDBwKz09YFoPhmChWToZw3VJhyQObVQshFFq3HUotJO
9ouqyzXp5Gp1m0dBWDW/AyceasZLxlRQcy7DtWFFSqgO4K+N/YDwZPgTd3JcX6qX
WbfqU/yprG6W/MR8Gad8vMn32UTxsaRPB2bYEpa4votr1AkkiiiS/nXqXqkHIhHF
Xx4JrgNV6DntC/vQGrLxUMqVe5A+xJGGDoLmzIIXfXIJSyq4rQKzp90vNg6N+sGx
ZJTCHC3qTIGBqOaSNuM0h9W/v8FUXBYBoWzgOkEhOXzlQSuV91rj++uTqEayS6GP
Duc5SvEA0wcqr9m9iG8dEtcOieF58pY+fy7nzgqV2zJgtVJvXANATdebTzlmFFDT
iaeFn5omPPPEX6MCl8aDXrr8SFF2I4EFAAlGvsffGR4CAFGYEXtRSjoZejKHXL87
QVvM+ISG4rPGMrP4NrwGwl3ksJ+YeT5vXIWkwzqfTuirhe5y6RGl7INcii3fNSyZ
8LGraSt42byP75AgcWr6aasXhITOUB5D7BeL8cCp/mGleulG4e2M34QgkTRO2T9M
0gpxC0HfJKkG6SqJSzth5XW8Bk6MvkxUMvFmyPyrTklha5//EVJgWgzUu+17mx+H
UYIIEnaIm/yT2LvgMsLBlGdEF3GHjEINevnaDfT7LGfvoR1TmnjuS2kittgfCzJQ
n8yCNQ7LsJN4Tu7Uak0Bd7KR8wqNstiu8Q8ym6z3Ffa4mf/XCUecwYl0+5OtNvY7
2/kcyMVDNZvblwsDzngZ/XEj8CptmHUXsewh0XyY/0k=
//pragma protect end_data_block
//pragma protect digest_block
riSjIfzQSm0xiHBMtnCOwHmu40o=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NFCNlKPxZPp4dPUOafEYiyvSNfJfvgjyAxFoSTrnvYsDlW8RNtC5sVoUkM9uJQx3
uVC3p4aDCQNHXxJDBDElBC8ap74m4CS2659wVgqnNbPkkSKTc6OT/KDGNmf6HgbK
X9PVPUZkB45+iSyfo5iz7rc0hLuIyOquiRqGa6yIlF3q84yUx44CMw==
//pragma protect end_key_block
//pragma protect digest_block
2In0N2e2ydLPoznIfEvQMO+N9e4=
//pragma protect end_digest_block
//pragma protect data_block
/ekAhguQRxwHUEniGRXDTRsQ0AqnKEQAZYzl8h62RY+mtVUDLVCIQH+GPc3xmp7u
ir6y6ugxKXkXmCxOxCEoYU4T+fbv+jHQXBm5u/4DdFbLawvO+GbdNrUeozJwHYzk
20gRT3fmeDZ++ouOLLDh5Grq45H8qjWIGMbSeJaCH4Tzp7ODNZBamb+0I/weJ7mH
FduyZGVobNZ0O5iudeByylgvbHqG2eobAhXGjKo0XxCTS42eYL36JYz2eMTSWj8g
XNiCI+kho0xeAih5Fd+TQVds4kJCmGnHj5IF14Roorym1mE4cZWSpAxKZ1ao/C5a
Xb35Q5Sg9RWLCQan7ZxvMjg0eIVzQldW2MJyiraaehYggp8udlU7/gPj48vc/XvY
HTaxKoqls1cCAmWftUZVRZVKy5IZmTPSg1eEddLuv2VArBJT/ksg0AOticV0uUaE
Igw0oH5AQuYAhedG0aqR3g==
//pragma protect end_data_block
//pragma protect digest_block
eZnYubGy+U206d1kRRhUAmacbNg=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
zu1vhY4qtxbc/goPo3OLb+vUUjtPTUesp+3zVYav6n70k1Rvs5xK24Z8/nL4yioV
1gVVGWlTwJjVtj34uJ8BgyujnK1epLAVGhMhf/7lWgc9kf2vEGYLXuR5137FSJIx
Rz9IeYB7yPgwe+K3pTZ6UQ831bs0Tn8uOLya44bF2kBan+6rMO2oGw==
//pragma protect end_key_block
//pragma protect digest_block
Y6dLxu+x4Z2vzphDwznUQVEAFgA=
//pragma protect end_digest_block
//pragma protect data_block
K661kL9wh+p6pco11nk6ef/Hlq1wjbUCvhG9crRW6McZQHohRZggi/Nqc/c6eEMu
jI0bPfCar9a24flPIat7NZI4bCkrLb28TQG2sMvSsMRu2i7YcV1CI+G9yzlqGvQz
RodBrbltjMbWymFOLn2dxISxUBNpJGbDIYYJ7jCZIfByhg6rGerzPUwmujeduB50
MiCnEMEOPorGoI0PlhRrBP7g3f+3/uDqBkZJ/AKheZtwcqOq+6ZivtRNmNao4mlW
0B7ggeQpIl7EydobH8t8ecGe1HDLAc7lQhGp0PHs75YYfmaxN5VOkoHJRmjsg2sw
f+G0aadRXDIo0cdje3VW3XDUpaehpgKjR2ujA1nK8pVXLSR7D8Mi4HCmDFWqHIoc
jhqZe8UHAkjf3KCVGgvfD/Acwj97GUfM9YvOixlrrzzncj+qlIsblDierZsW6cPl
Z7PtYu+zC3k1xLDQXBLWUcCD+md2rRTbVVi9DuhgsOK/3PYvQaNf1arxQiTB7V98
3ZhwVgVWpA/GUgP++wyyUC/XbiTSbvOuADD8soyOlWKnWx3B8x6Km1n0YIc4nGly
RNUysXNxMt2raX9WZ5sucCQMv7O+i3LRCeddote0GJnJY5hAX9CgD/DGvTEEMStL
5FaMMC+eF47TXKkDfvAlPSYufHfeRedXE1x3s6gAx7H8W1TJxvIvjLc5VPDHm6fU
nNndKUzWolEvFqkxfd0AnGofUoSsGkxjP9cyRRkE43PjtaKhdCf3jHP+nnDXg5ZS
6nb5krDZQApv9KCZ1nxOY8NmabgnQ5iI4IxCgWzp08raC+5mDVTDPHIdgoemU+Qp
Io/84tuFVig+P9UKKJ4+TO6769tivEgpOB+EeZV49njjoU7sxD6TPnigGtgWSgaE
5+cN6o2F4GUqVaghyXWH4R4CrIrllTEm4MUQ5784/xyxwJZ9JZE2Ktuyw4a5iwLY
4pEegy1IqTBanYjSIGl835Fs59lL6QCywQEAMBOvlRL5W36eOcOKNf1yMFWeh/cm
7i0UkNmBoyxm114mcG/rVIYrpXJnGzQZyV7iW/E/0Ve7GilDqw58u2XiDi8QBvgm
C1klXKpUVAXs2B3OdMjCMgv3JHtq095nDiu6YsT6bnlmr/mNyb3wXayOxWxuybhx
URSBqGXVUoa+vhK3Etfa88/dILUROkoT0ziuECicY3j372GVb5kFMxjCg8DEoR9P
1Yb7D94RWXnUe89HfQ+QaDxYbPxfVTnnkkOEkkeuk2cOoxt6RPcymnCRYw2D5Igu
uKrAqITqzP9hA9K9anTX3pxTiyD4dWyLby9aSiGZX77UFF2fLcZhpPV9EiiI4Qz2
scvrhGzS3+HMvJLxoZqP+Js5yj5PJ15rY+Ntx1PF6AprjEYPw3/toNxXZoKijQOU
DN8RDFlWH/dLMU2f7XiURbPS6xkmoT4y4XrMxM4kBmuEk/sbrRuQSK7hmBOppzbD
xvDGxEnmIiyccFS7nRzfEzZJGRM4doZ1PMTmfZQgOh8627sYqgcM0OL2NKRhh/GY
ejw1rvIU2w+FNNQubu0pe53uwAGsULfLIbf5OFh7pTXLTH/qcLR0qDR8gA/11jue
iLdpHE8Wh7Z35BeuNKg6nHHrMzOqBDZMdfgUmfxGsbeh3gI/W11U71dfLsuEsJVi
BFwTpI48EtTHJ4vMHOy0t3Gzr47CNRUlTBAbvJv6gNjaN/oCVbh2D6DCOoC3/hiR
bMFDroiu67T1q4Q9oBwnolX+a9SxzKdRuK9EovsfXgKKIuCRVMV2Goo0Xo3EyoCB
A8/Ru/Le1JrZvd6uVJeUf3esaFedLa3D/0yP3TFQJKCikW0U7d1bkuEfrnmQuSHZ
ZWHCaV264Sr7rBx+7QIuC5/mfZEc1g340P9DLSVA7cpKZphiVmiHB62sY+epEYSc
YaYKaK0V4QNaSbc2U7n1GzzFCJveFmopM0KYETBr/NlJWlbyfGqlKfi8po9MKi+X
9RINzS1CK8wUNPhhjbV1tmr/y5cMlto1yOeHGRD+CsJZV6+mSlQphh2V7XU0O/WP
jnICb3EEcwlUczX//ZU8rl8yJSYlhiWU0uw0MVCkLjZlYv+36+oouIPJ8vPAXU8f
MWENTMNwhiVrbrnAkUCVn1/DyJwcB7d2n90DrezrYrR4VAP8O1tRn23pOvn2nLP3
4s13/mNS2JNjUqdWxE2fEFcM1LAwnn34MxUJ2mCBn2eL2YF3UBDgqW/KDOMCR/MB
uuBHig6aWn5XviQqr4IahwdExpFVKQrqJjRSDjqRjyCFXNlN75JWC3rJispG5eY0
Exnpq5Myk+M9yIv6+zkktcld+SD7ZW9vPQ0qlEo6BSz1XiRK2CsagSPxBl228WUs
irGAi+J/llQaUZUlFqqV+jeXF2w7A0jjKCWx4d/IPX2KjSKlR4jNJjRpI6beETtB
HF6W4tQ0nAwfi4XrPUVGH0l0P6Cb9e5ccYmET8FlAevEZuRhuo4RwdIXSYZCMBjY
5hodgxDRZIOTF1hzEjKO7Coe4r96qQew67O+8g31SiSnYULhJcr1UR4pro+kJOYe
9KWVMCzo5ALXltIscajCnGuxKA/B4R0Vi5mbIBdISiWoLZ5MJK1rjlBdFKIv/rjM
kAkdqV4NFUd1EZskJbu5bRctQqe16AZYyWtZAeftaPh5L2dbfBKWIPBtCF/zyEDw
rnUYAIELoFPsh3q+rkhzLeW0FTiMB1GX7Y0lGIO48SK4Xb5Yatewg2dFA+iQuW2r
m/luTADzuQCyj31tbTzRGZohmadmLYNg8mJrHjrdMXfAEf2eNEmBojfOTdUMSVdh
EreyVfcpoY603hfaLXA1W187JZtcqt6OVGAizw6dnEnjaagYHiEQZtmdbEpr2MkO
FieBLvvve0HEyttkBMtNRioFsHWfWWXkpYTqe1HEZ5716NfFxRrr2scNS0rMT6xe
HHd1Tkoo/7U8N6pPEBaxSkbav7pbJq8/QmIHnn6MgoR49DShInLUNKs7xHP97QQ1
881KoPs3U2/V8R/AfCohpdt5YhTr3wqDQcjNr26MCGK9MEPsKQgd3WHJugwSJmJn
ICsZNsw/50kgL4JMhgMsipPDuRSdnWS86SxQb4LAkvLHynhyK9izycve8xbHHXoO
GIdV5+oMvyyEhX7reSrJiTOLn97S5K6H47c6lWlJxYMHSgeO8suh6r3bgBD/B7Ca
OfAMPWj6Z3UCEqwAq5DcYhoe2FiKbJKOAAMoV5auHvfyJIMlqjaLACK4e1wxlZiA
pha4E+bU6d0iU9R04FlimDMiFL+ymc3PxkA7jAE0Q7t45uWNyzcolIypmnFMsQDs
1L+9u6l4cfIsHegDpPqGsPrw/xZ6c+wHZBpOFL7fs9hC22qNbBIzKMnM1LojiSJX
s1nEOqh3ECU2qDgUH/h4BElupTnajMkgKV5yi76XNV7twjf2uveJCIe8i6K/m+cx
vcaUXai0JqmRL+n2PW0SIC4QpX5IDd6H4INwA2wTSyP/j5Wizli+o75OqekSLZU+
8p6HlmcJknblQ6W4vP0MPx/Ha8RkExzKaJqMX9MpsTXES6wOPOn9+XKJFtMt2xCn
KcN6iVwXFyXl10wnM2Qjur3duYlpIqwI7MdJN4fcbhn/MyC7sj/HYMisnWojMLYl
DhoEh0gn7B18AXK4kZj2C7ouT1vyV+GWE8iMmErl/OmUkJHU+ET+TLsAt0lL5/D8
HKfUMA10EwtC566PCPDJfGzM+wRoupsSij+XinvDwNpNG6TDMqSbwpWNBvOjWCxc
ipkKKF16l6rggRUL7ps+/81HF6H4bn/tAF29edvLMJppeNOknXVLcUGKro6psSRC
B7tTyZKaNUdM+UqrnyVB9nhm7us1vJz7KXGFDYflIxTYRi3UfNEx+v4TgINuraxf
VVH41G5/IVEaoCKYlPawIl//Vz5/34dnYwGf4D60lVIZt6K7dI+CnhL4NWkyz4u5
7ltkNqZaS0VdhoS9VdSKWf6GUggtye+0BxhshhljZoNOjfmK23fCDsd0accAx7/k
jcaz+oVwAfQ9CsoxwmiglgM51HNQu7yjr/Yvah34MnXHZzGAtKJTLHr/xQk3ann1
6qNws7Y1r0zy/Fq6JPcCTOkTcH4eF7Xo6TfnoJIF02ZeBx6fWEafpZ+gRnLTEsRW
6iYkMf+vxAViwWd09zqMBv2kJ0D+xS20bBGWL7qKgV975azoSdI1WKdJUpLClENB
/psPFNsQhddRdNa0DXWlRPrmBTQX/X8fVQ4TG3d2hhiqJOws0Rk6PoENhUWV267a
f+jVFq85MROGKvxR15cXmqLyfUKfTYR9P8iRn9NPsV83PEsTAYf2/FW916VTFZwZ
EAoRtvGq6no3Z8Ajx5Q39bH/TwEES9UImZvfHpG4FKJP3irk4QLpLMYtltz6hTFL
8xmD587k0mw2BmdPIeQJbPRpmBKvFWO+gl65Vcv3PjRmL0FeLPdK0gw69KxT6bLA
jbOMFQAcsx4v8Lr9KB3SLmyyWmRx2RRIjZt+iBf0tKRH8+rY53d1Z7O3KDuOgTf7
MCLdMCU8WoiL0qyT2VuExWhouPn0t0YufN3yCVoTRVqYfe7r4y8px3gUqVYKteZP
zBDTr59dmi8Xg4yGJXE8MxIAEslb3a8JIgZc0lTbj6gKO4mjYi7ad+UKtY7M0XUi
UJBjgeMPvYo+GDdxSX1m5MhdqfEWiZLwUvVXuAozVg8b79MjcZls0uCAMhcAog2C
DqoOTClnQxik0cXsSWS5DmlMy5t6KvGLL3lswByFJ0fDansNnGoRyRl3VygKMwsx
J49rYmVkEFOwsTARmx1dF8ThFucm1nZyWOS26nJeM2sqeeiF9XQsPQyvx4AxQutJ
p4n/it/GLsh/tYKBmkZDXuIQOxiA/Ux2HLQZ6FRQOQmTh9R0ea2BMhtsSPHhlF86
IEijoi02BB/pJcaNkFWzy4VBEkgPp7/NoxgRd8NLGqMqPmgjmVYuA5ClxPk644c5
QGZyoeYlpliiYB4tPsyQGQM+cMlwHDT3ylops41wtQvF/W8WUOp1BxcSG/RkYqF4
1JrxVMxDJ1swE4ST0K/5hJAOBNml0loeIB7FFR+6SeXCtpHYKM3kYnI8Tv05aPWU
P06HGAQiUNPQ4v9sqpAzMT6eUEhii5r+Xdm89awMXPsL3MFD0BH9yKGnzrhbcH7u
wZ+FzVAafZk/NaPS3KCx6EPrxU1aoKGIJpczxiSHUIRb/K8HcQk5jEbikrDNpZqV
ED1srq/n5LmymPnvRZ60tdtnig4MzcTLhfJ7KsDz0sMM9WFt5/ek6gleNYOjzB4F
kxkgao2ca+2vLr6fP5GzB3x76SM9HjHziBVeaGZLjAqZUjJQHetVCJAQPSGOrkrs
mVoUHczI73+UtGFN7m/Q2UGoc+dAQRAG+QEarblK+du2lGVQTTU5WQDqDxxw+7KL
wD4X28v928OsBut0ch0TYUn5aRA++Z2uGHcLgRNB2lNKZKwGgpbsTHDprvv78D5B
MN+fMv84BVbxziZeRStzDtVNSizucR3sXSFBUm+yhkhaRcyT0adBvKLN7CqGMPHP
4NCOmPQXLHxi9HVVer4cuhNthTvmlhnNT7fklWqWP9nqBo8hTzmA2xDC4EC0o3By
5y5HaxoCAvyiplhqH7CuUjmpC4adNdgmfB2YaNDJLmi8eIaTPCxz0gaJ4Bc0JLpi
6ny5wYWRY/D8t9kV/+96brAZnQOP/iZ/5+FnEYv4AtzMG67CpZu6pmHX3puy5j9T
FUdAvFk3f+wgCTxAs6uJT4LmHtfJiwpU7zTii7RtoEAD2sFFQ0pu+tCYobdC1ugh
55vSENmd6i4cVaA5jpN4wC8mQgVi8V8QL5qlUojGrUDRJyaDXj3c5LK+s915DXgm
zTlCotdLGIoBDF8JHmZ4Lt8Oxe1RUrbkBmiI5oDfOcz/w5sQZra/TfyfhuD9S6fO
pqIdwLhC95YgXWP+vyw/EFgQ1C/lR/1BVnz0tLRV4rxuYefCRskAywqiEFp2lkTW
ZKjg71XnJfYTyw+6apPLwD+7a4H3fBr8aBU9tpF6vw9DhKn6hUlVXA1lbfBo0GQ9
3Oeu9Z99JqLobyoQ4frMjMaw+cw+nRvfMQNHku8AhiQ2IfYiBYddusuy9/buxeD1
gcFa3YYQC83k6e7GTGPyRHpff6eXLgOsZ/rxWg/vYbioTxLWGhVecwhvmsswI7E0
UW72C+C9NL2HY2wPhWAFBFkCoztINABOLj88Mqvv/0ykycsM/qJcx93bWNbJ/RcT
oz6kjvXMPsCSq9vWjbjrl/OUkG286NYx2ABFw4k6VARwSjLcKuFgQ8omHnC4P3NK
cylufvvV02yJT1v+/4CU+/zRl42DyXu6IkmdJ9Ef4TjhX2RLbviGzHFpI3l40hyr
VV2l3xcF/BBBt14UTxaHaMywmL1+NyZV4YQt2FjKOP2dujfLTiZw9ky7xWmKeDHf
2np5Xj02PV6/ZdshZtCbitqYnxdtqdaXIibRg27hB7ci4azHIHaU+VAmcDtjJXXa
L6EMkkgh8jX2JBgq0h10gdn95B15fZA8/YF8jOddEgiezKUZdeGS1ZZWZY3KQbYc
cAb8sRTPgLDdPUbHRouIda5ZpoQPZKWmdOKJOyyX059liRSW7ywAjM39PzYSeVJe
8Z4kUobSAY83GQvCYVL9efqnwNu4A6AjllFlKVMXloBsx7wxZvP+ZoDmNGTKnLca
+JUieLDv/loZyJFsN7+Zw79v/vZv9nJ8DPx3kxeybMH3gsP39l2QUAqLOiEpKx0W
qZ08zIvAvQnQU/9b62za2iXhBD9P9n1TSJSbvx8vszyJXiz/FvM1suEL4VrIzPKq
fE0G9nFofBXzs1BeBo3J3bu0Qt9HXss/0kti960YNzJeC4hDlgFfMn9kCb9CBrhB
rXwLx+F9sKbadfGCAM9kenJnPwfO8ozcGpA6oyXeMkZHeLY2vWTOgLsdaKL8dj7z
RMCVMLdw9i//f2VOMpUBHghHjtYwX++qxRAZet+mAk63zlBFTC4rTzbNNUQgztXe
k22GD/93Bh8nRdIu4oo3Bw6cH7NBgr49oWbWvtZBMTAFS0s96epslbrhwBKM30fo
n2zFBEciib3ldXCPU9/VgLCkrQ5QYQ273LX2gub6+1/35CCKGWhY1k7i0Ykop/Ak
Z37i0X1fYT0tFBiYN2QcZ+7rCQFAMXv88JshWJ4FGYuFDMfWx2Bt/sPuKUt6FG5C
LFqH8nMC4sHL8mCnB7EBeGItvvG5hk9xpnmClxpdusdxqSTE+4fQiaYGDZe5lNb4
4A3bjZiXIZGWg1TeBvVC3aXjXMkNnpVZINt2NOGmW6uH1r+KzC7PoTZfmuslPGjw
kaq6DhTRFqkJtJe9TJBRCGp/pktAH5pyvei7N1WlpCH0WqdGLr6zF7PFd2EOw+QR
bAJ1E/w3w9ras61/KW+ZcrtM1QsE28KSlj8ewSntzcSjwbm1DMCOUKsG6jd9/IYx
k8pozu8cfgYmObNbJvzrXv3MoHTqxklcCpYd0s/PFRaETDW1f/IgnZhBUBOX8T4M
aMxVp+ufIh5m/mrF9n2MAf+sPQ2llVQH1JlY8YVSfSmIPfGeGDfRa5tGqwFUM+94
jtkdtZl0oZLDqcU+UIC8qwZ9HllOq6xbKnJNaX2f6q1bCOEget0XGIc5f5puIS9l
3u5LujbnSaAgOY/IXg9qNL30zwSsxAqeDmSOhxXp4D2c1WcDaMKDwSwhyT/aUmXG
mXVHtf6vX02ruknef90uYJyCEW+AnGITUVoocdnAuQUQF1EvjSBVMhF/Zg7q/Blr
SlXZpQ6kVxCkVqJ5Vj4v6fatgCg6aQR/RuDy8839L5k5rDOxBPp/nIpRVLfYLZ6u
YzOD9VKlj2xTXOohPLVR0w8Mv5YtM7hu+Kch2Ei+G3y7ivPULUPwHKTsCBvIYGwz
yKiAshwA8NK9USjLHwCPfY/P7Ru8trQiTsxMENMb/dybmHUg1p2zfY/+cHL9oNoO
b8EzBSUnm/PKqGOmFxRfTvQWKS4hwmvMaKZHDGzyGbhhftGeSCfAX5F8bFF+w8SE
gn1+oCQ4mB3mxL2ZG/FcMW5A9lsl/3uIRCLbdXFuUjIruJkt/FI8fI5S1vLCRyPw
7T6JupxT4U5DEcF/ge9CvkiA+1vl1WxWymkly2czpMeqqciCBE2p13eQpsHsnR/Z
pVktFYWKStLmcflBLbKQRjtWXTsOs5P2OEXnjh6cHOmIvDBxfjI6AUOpE+aAH4NC
Gq/WlQ4JRJuuiANRpQfTAZm8XQ5UYVH7oritVn/Hi1jtMUAU++Dn6J3wsbR1biuV
VYEPu2OQcULe7U+MBv36tT2IBAfZEFWJvYoaMerylbD8x6s4u/eJmCRzV9Dngb4X
/i5eceZLLVKEbSegKVdCnhDWpUAuokD09XRZ7GSwCsKBQ1gDR6xvz+qcplGrko5C
XoYjbCj9re4MwAZPa2ZKwPNrZYr7EaOAuO8cVYi+Zy/ReUxMpaSpyZ3ErbtpLJOj
nEFu/ASzpVBmMiSkKRoDLHX6xBqka0lMffltr/vtYu7FsM7W1b2PfP9gGTK3iFc5
sSrFvW8nqOIcCSTbQVd3e2WDCg+WaXWqL94WRo4QSBizwpLaMx8UZ6x2r0HLkhCT
bad7tQFnN8D0GapNUGxZmp/GXtoYm9CtKtL92Bjy3Rl//EVAVMwZdA+QPevsvzxr
kR18RlXRiB/o06ilxcC810PqXX4zwrE4UwGwhQ+PqO2ftt2wB5NOrJ0OE6HNXGFk
o4mJ5qE2sJ7k/bZuuI3opPZ17WNsgxE/Hxv2mWN4A7SXNIwDfd4JdidUFczx0CHG
4sXVZCfp7Dh1IE6Wbk0610yGyUgUy+P/BO+q9fUKeeFCxoDWEZ9h4bOxBUWi70uz
vcdWbW1Xt17sN0jm9OvdLy4Mi9r1T2pEKtbOcXKFHfzdQ+s6o6mLvCh4ZqAeYxAU
4VvFOeYjvdWsjz0oT+R2eV+KHadihteuCUYJAb/Z9NEuKN/u+/3+arUW1g+qM237
nCrkVSSQiwi4/u/5T2zytX3ZvDeJ6mJNkWocc6zVADnTYdrKCs28Qqd6TMMLASX4
L25XzIynwOtTk5lhY/msYjigOvGydDmyE4wR/5AuQ6Wv6YGT4jOL//ohRTj0zIbf
iixchrAWzlEsQm6/e4mx2/Mz4DVL03fvgZiRgWUV06LDexFu/9jCeCPRYuO5SpkF
BTM4jC4o35riz1EogYDQ3a7R7YzHOpoh9EMRqqFEHrrcXS7G5Cf1ygzd4/ZROlfo
qbVB7YTpWSf/A8UhONmFkScv+svvbRSgVzCkrZL6aTuAzvsiOrjISoSrZ+KXQ/bH
9Axl6SfC522+1M9no/kMQ+JlZ2zfOu1Db7VqCb7kA4Jug6HCQXZdnopgXgPMlrQz
hZPPbVc+Nqz3PcLr4ItKNfYTnoxh3XLGmELr0/MuVy20eNADxC727Uw8v7vppe5G
5e+0K77tO90jqC+l224VPQopUCMtUC9ry3/bxDe2yCOlDGU6A5VV+3ZGyf3WnFXw
QG5MSbuvbNQr0h1xhRxwTNcHvbb3ciwfPTNj3H7QYg4I3ASLeB/H6sPwOnGAoqQw
xzMXqUlh64rEfudAaC970C2kuXN7z+s+3I3dAixOjWN6YshqyMxX/NI54QbxiQ2p
2q9tC1tvUFgejr2GJIWbrc5P9qG4aezN8xdFB5HGv0XYJd9c4+IsWSc7InjTmuqe
isEhS2UhFR8rFmE6lZfsYBMQ/DN6W+3Q5sDq3cmueb6s4KvygB+hFprdYH4sJ6Qm
+ye3qTSMBskS7sDdwMtHFHisGSBVc/oeer/iocjJrnXmi3pVI9hvcKIeKfvttcCt
42eeXVMqqow42t0JxybMseyBDv17OeCfynV5xsRZWhAVZRE1YgPAm7RfIFmZe+53
bQCJhCHeNZ778vRlUN7r7+HEfgL8ENTjQJ56Yqlc2G8iajTDVaUK9gl/WUjsOcw8
pA3wOkfErDPvNXKWQG3Xk1mfgSs7jTHr/N+D3Rvc2J3ybhMxso3F+40ICOeSsUfw
3lq27nrOFuQwgWTglFszuwtBQqx4uFsxTM7R4L7Wc6QMM13tEJI7KkY7phMTmDW2
BLCWXIK1xmwNopfhwk6Okz/J0vPkVDB3l4A2EZbpF7AAXXpWlvjxXKd8k3jYqixL
H39uEfMzbHHwTxi19uRRu09glcdUtwVKKhC1j6wUxQA2wijO8sbguW8n0iMdsMSs
pqQU+e7L0BUJ5gJ0zUjhm7BkCzJEXW6LNyg9F44lZyGATSiOddA3wHZGV1WCiZua
VDzGNe2hzPnbgHV4p5GKsSdIFEuWyevBFjGZSsGnwXOwqkQWBxr2BRNeEQ2YbApa
J9U7g+djXfFWePeCFPZax9niEtRrc2MAC3Vb5hUJgxPM1Y1vAkp25HeXqb7HDvvG
va1kseziLnDVQSfcVaeZSBDvoeWfBu8s1P7Q3zJzqV4f2cC/1hwQeP868ydYAuYM
cjimfp2g4EDLakel8ZMV9+Zp3oTBAfOeoWgj+/kV3EGiutGeIv+tRDDA5RbG1lkz
bpfVg7dWQ5FiuwOiZ+AB+j6NPxJ3TaMqPixIwUIFLYMS3WlloFEn7Tek4qFRr+rs
U2l+bNcydZ4OCp4fXVTSAviBBeR7PbVptdzfnJV9FOeUW5Tjd0hZYa4UQW3rV2No
kgNjlbchI9l/37l0zoCQ6w==
//pragma protect end_data_block
//pragma protect digest_block
C7SraC78RbJzFQ6+1Kg3QJh9kyE=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
4YiRk66wudfQjsFGohfjJjta1ocYKyJFrqU8lg34RZ1smeSJaAaVbLwAFkRmWbAu
SHt/yBTBiTkWWDh7Lup61uXrVp1q5jvr/1ZIjJ9oyKFrRd35h2YnXTEcHz6vK2E2
FG9cS+S6oHxWiZpZ9A852diGj+7yU8b+P8Y8nU3K8NmfuA2G6tBSkw==
//pragma protect end_key_block
//pragma protect digest_block
qn4Z1xQ36iUS8SEfA4m0CfuFxEI=
//pragma protect end_digest_block
//pragma protect data_block
G1F1+uIrl2u78Ta16LzBjYy/atO/TU+f5S6rT46dDL2g8jFejTJzXnyWTxZSqrpP
shIZYCbHz20vLAB2TJbOs8mgxbMYk9TKCUH3WIXlNIt8kZYmdP5gcLnz/Y8iW8D4
Ku+pTMJLbIFk7ibPrmcYr42oRsptgdpgCOpbBihahmPrTK9okrE9mNLrXi/2qk+5
tp6dN4XNqJ+wvLT7YNNOZuyWw1C0zWue3ZCAv+LVqX/EQk6Gi7lQ9mJY2cCmXU0s
vLOYnewp4v23JyeiGl0L5SdgJjatkPmeH8HJIa2zagDaVuMsjGXfttdjVFu/8eQ+
sGag0a3SyujGHqDI0460YCLHZBrrb9MqNLbMgnqu28TU57n/DHyGDk5FpbfkErEB
b2XkqdEE6M74+WU05bkpzSn1wBJvZV2MfFwvooV4cU2LZKKeIIA6CXc9D3fdlqDy
QlUWopCcdwgOwZa23lLRX/kXng3JxJsXkexoPsv3poj1On6ysR3pUoZs7LRkd+Eo
CoU8a06+BSEQG2vSk7vLelnLs9vdCfAXNM17om2UMDm8fhkcqCp06LOIuT+II24C
ndDcPa7bkDyG8SSISSj4a/s8a2zzV+zfa8qyQ9+grXELRPnOBjtSWkclDKsQFy4Q
OWI5zGD0Ra6ELduKERiEB1pqQh8k3KCkEG2d6yfkzAQ=
//pragma protect end_data_block
//pragma protect digest_block
9hrWRQCWSOxLC+D+jgPMBdviYv8=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FlmUsOltQNrwhPeUoF5MyXdKLcmJg/NGO+y8ms47PA56IWbYy3d86MCPiuVym13t
RY/0moCPelDWNqCXmSjcIWX4vDD7DTgp8VUeLjI9IEVMjUeMmQO9pTjGSF6xfvMK
aTbISJwkAdhBPCPS4Q6P/IAYwKUiW9RH3OcGZOpjioM9fbolQ6HEkQ==
//pragma protect end_key_block
//pragma protect digest_block
yNASHli88pHtW+YyT6qEoqG7U48=
//pragma protect end_digest_block
//pragma protect data_block
F+uqYcpfybMiQvgqGe8OpjszBk9EWuR/ULQFzh8ONVb95gdVbcrQQUH62rGa+X2a
+tDGU0GylkwiMNSIRLYd+lUhXKyf6sm9mE5yZMY8CtNfQhcpCGsuco6ODEAjU3vX
0q6G8Xs9SV6O339CrBlIYOyjpJ0PASABtc3Ei8aXXcxKXMNK3P4btjlenISX+VFF
wFwKEy6yqRqCi321peM75Bi6KLg3zEGxG28ACtl2iD5RcWGRYhynHg2oUKhqusPc
yZdwrrZjJBcf40chyfIuj/GxnKkAMotCgJIfHBaQHMTZM0FozDhnr5W613SvaOHi
rZwt22XHY+gDk6EDrXXVfZ1SVQ/S3/rHVztK550VCYHTHIdgm7WE2GFauK7CVZfz
Ukg3oOvdBt1OZdCC9UBSGeMHR2nlRjeB0i4seQOktMkOOaolxdkQ+fZmxZ5okhnG
1bDdmJKsg2vHy99/9mm1hXSLCP3DxzBZyLz+tMSbH4q07MW+gobKgOXol6vwbsBY
XFRhfkLo7ACgZaEE6Zff0zAPgMIWYQqybjoOpmVA+RF3SgnOd0AiXfvfLxzIhZLf
qhDeah1b9CYfG3VGj/n8XRUMvCYuK2qyoVAlBUs0dih/FEaQ1z8A6MijPkMi6G0R
Y2tADM/sOTalCZD+gXrT0IM6AuQquS4Sy5IhAevYG4XSSdIVg8SMR/89zagoDKMA
2iqTk4SVrybVaZT/uNXPPZVRXN1Yrsqc4wH8f0Xlaj2AiSqZ+6y8rqnOHTv16Wbj
RHZXPl4I3WJJ7NeWeNnK3SOs509qv+RcRS8mhMGYUvUhjMuIMpwusWl+vVjvvB7D
vAgBYb/p78AiOEDqz5uYgAaMDLbqMtpq1ZmEkFpfiCiXriqlDkW3INkqqQwDzryY
2KsAsA8u3eafET7dQkrNRGi5oUAgJmVdkoz5G4SSUgWE19BM8S2AUOF3RlTLHZw7
4UKPUFBHqnUjqcxYDV2pP7DbbFC1KUv3GFVeCWGorYr/7RfVtLNPZ3nUT0SU98h0
fc+iRHfq5x0BbaVz8uBfF95gCssplkfT3jKCbInVBLi08LjjnA+3fXF0YnBOJarH
qxXnniU0W8d3qIsI6XZZvxtptNPbQ81Y58f/+z50Hoa5fI/8Lf0bHCIBJcuTIjo+
BodTP2T456GH4DiAWZBpmiPWeUnSJ3y0hZ9vQESdAwIHXwvLqCBkFNZHE/MucI0N
cm7u0H03ly+1m8BDGT6gZyu2mJcQ3nJY4psDrQgfUCspPQMynKrUcd22jlxD9m3K
dNNdHbbz7HUbKgoSI8EjayUfkksmL8Dxlsizq5BProXQ71smWOfn8PGwOLumF7bE
YABXhUsUxBSRqIOOQukW6WWa+gVQaUCsG72SM/q5vQ80iqwWvh4qbKzCLf616vkG
ioENqpFYRKGfzRkd88dMGzj/oTioKdXy50umhEtgfWuqQ8cbInfBc8jpO/q2IRZI
gdSiHaR3d40vXP+9diDDKE1RX7HnicLQ+/3V2KIeEAWc92naExO5sLNJBp1rXue1
lJxHlABCJ3BE6WVgwTo6wKwGRW/NQPTY02bAi5rI3Y0JAyIHsXK8TYSMr7swgtwT
H0tfpxNuJ64SFqbw1NiIl67Ya2u3+iQbzXvn/VY1cmCi1WGtz64cZg9PKZ0dsM9i
QYpHyR7TyyarJBSjV04DrVsKNs+NOPIuveK87ZXjCMWjusuXCU0EPZxHlaHK0+Fn
IL0VosNSCm3RLENY3uk7KycSAgkbSNlEW7jqxHBz9rvtbrbqAtuYFrK26yBGThMQ
rH+Xu7Q0QGytT6zrTsDHHh3kNaX6xsFHoivdFFkd1ryVivsWUuYe8POITMsaJ88H
4RZR2D5BWe5O7EY0xM9IIa/NfU2XRiaUC1sWflxS2CR3FsCsfHdxolsczF8ezh4/
XjPrI3vPUl0PCtNO/hRVju6mv4oAkzo8ZfrWdTbzDnzrunAHwRJBNKsZPCL3XCVg
kXSED9u8anwkB+1OIWVt8wPiy5OLLeWJo/FFlu5fjKvzC8RDv0fyFBkBVGjuPfb1
YfZPTrHt4cu37m6LTrTTJh+ugYJLJ2bWBkIu1cYoPjQHjmVrWGINFD+hCgfgWS2y
/ysKRYTRQ0ntc/yYOum+NvBcOe1amq9n1Xz2a1VLkLmVX5vcAmDXRmXF/VvrlKhi
phD+H9O+IxU9qbciVR6qrQ/xH5/5JETJHagsAYq5wihKblNEqR9HFbiH1aQBpm0l
d+oovC5691KL3o14f68xrmX+2DebTZVi7/z+fd3e/+ZsgA+EWS+Jxl43X9RVI959
mXtylRSwCLR9qpQnKyMvlzBAzH9MD3tY6NsuiH2mY8DlbQveeL8MktHnA+RP6aiT
jbP1dFwEs3ROvl6OGeQH3eg9UkjGXmBTr9B+zhPYpGY8F7KemB91kb5ZiI7kxEnp
BWG6tjogEKlb1DIoVypKk9e+WyoSMicu6zQQ3SztO3NEzLBdAxiT0pm/7M2j8DUj
erH3myMn8q/WgrYc0uLzbwpiEG441oJC9t2UwYtPcfFqBDkXTroibVGkjZ2Sowq8
AIQVzr0sZImmsDee9TbgJnfP+3z2u4ZusMn2ChEgSZHbOOz+h+8lzrWDEfyeXbEh
RC0zRsjVbCjbyef0+7M5XdAe+G1gB8c21JyYoYav9UYk4pRqblfjyLHN2xj595gB
mhPrSsrYyN4oTwnLym4ZyFdWyo5YLoiPuMTaJ0WrMg2XRb6aeYYxCCogO1vysPzy
ezPswW2Esq+SvjsLfPBRWpATnr8wV7m/eU+pfzRmZFtcL2ToeJeN5eugeNYMBx/w
xUfu05QdXrhd9gzWcDTg17G/czX6Sqo7JaJvd4h9+qOjDsCZj+CkIgCARWcoagFn
KVY9ceYcwlSIbCEoLN055tofJ0ur80nu3TTZSPWcQqqzqygHFKDk45vxTjyVnc6A
1JkniXPo6vPmou3WeveT5cLxzvOkQ5uDTSkFOMB4ouOE63Hi4kcDSopQjQ7+iA0v
+0DpZrUQpeiUQiBGBj4DZZgny6rb1ftlFMISn5AukTg0Yoaohvp9MCB8sv4zxY/c
RaP5vfvHYbRVbn6E79gJC/5NijH5MzWJAk0UhsTWI0XonbQMoLPlFbjWpB4vbzIn
PZeUVxZkAvP8asuPEGhPJmB77jjKr+gotSdCBPQfsbMj0nLub8JPnJrCg4auybpi
VULNawcds7yrFACris1tdghbain06uOdhj+NMfZBeGx1D9zO+tt9nmxYlCAKnVrO
RRz3Cu0e+M6mllm9ni4tLt6w61gB77xySjR2OEZU8Yt6lCg1x5JdIzTKDWpVFcl0
N5Y9R6ataW9GnM8bfuWFrLDfQomRLd2tXx9jyNMeJZBY8VTeqCstGzXt/ByVsxaQ
f29H24NJdnU8SHvfAcQjpTZz6sUB0SPLhzn6hN3U6wixMjddayl4+M5r/BEoSAIG
TSrFEhhJPRvbLJKHO394obuVzlvYqy7C8VduKe5ZYVT3/J0O3OKUtbiFkpEUESI7
irZqqAkY8mjK+dN9uZ/VeBBOW57YZtiU1WkjUXJukZ6fjrTRHl2z0DKW4JsMOvfn
vAt57xb9Pf8WIF+XsW5SjoBTahaVUd6fX3vTuoOrZUkwd/kX8AuXpyY0RNPauFET
nO8XCciwIYAoQNl5cLtdtdJvjm2IyqkG2R11cCisNKcsi6pOte8bJiZF0Xux6rIi
jYsCznEA4OzVoABajd1szTrB04Qdq5LUUKgRkYkxhUb2q7SouP8/25umF5o7CX0z
GjLRklxnEWgdytnpV8ks+dKXhWk/vzBD6bUjitSr0Nw91vt77iHSeCp+6TxCJK6E
VT/jnGqU1GjCSST7e7Vnm0I1v/++9rgG8GWOqE85DTt9zoBNThMhtIaEXXnZfOS0
izk+tx2odxbsnr1h1Gmj8EspBeFRI9cRsrXGYCmHPaWIaEcr8zUKl1LNty59wRlK
E6Q3N31IgO7CStr5sXDilPo8dhmCZ2t+w4rw5Wv2x27/zGtVNaiIhsRoF/IQQvNP
oW8bblZbor36Tn3p+qznhqzNr0XWH8jddbehB6xs05rQMRWH+7MA2dTKiYSZPEey
WU/onkBvKHezHXdgWA8GrwSJ1XZrO/TQMcSTyax9AW1NgySX8lJEpYDxB2+VdcA/
kHroN6c2Uyi1xf4zLFOy4C8MFw2aGnuU3WYYlkfx8iqsSIpmyUYwGYa1hV27Rn63
P1UoB3rTp5O/RSma8elDeBpHHTjKPMStZlK1WUnVq4ilyqVtDp/Y5SZo9xshoVCR
6BPz2Zq+jrzXzGcwP7m6kxCFI3X3O11Pt+0TZmuTVe3buwmHakRDmw4kNuDuSj4y
hUQeRR54U6dNBP0gNNgWnRSkQfObVVtSSh1h3Lzta2/F3vWp2Pn6sF0WlwtjpnAT
QXm7K2oeWHsSNmbhYLdCicNU+3L1nYQ1pKPbIxQ3DOeiKge1Xz2wK+xLtwx7JLvw
y6rX3LQTJtOzTiHQWo6mRf0rI0yBZDl3EpO9YC9aweirgKUbBUoc2wwqgtjXmQlE
SHwPkDhHZJnoDthJ+DxW9KAVmaHSKIPf/d86nm0OXp48Ucyrydp+9vUUlqbqgK/z
TN2gOj1UmMy2mW6gC2MAbpxhQfvW+a6Q3v72Wd3SqgfhtkkQrCASSTX6E4CoNQNZ
1WASnwoHW4UXVfE1iCVcBKKIQ0QtWPUDBJVBFM9xUDEISKKiXoTzNqKEWvy8+BHf
kRJHSYjot3uWb9+YEGKSayQx2qdl3w8Apr+rl+xr4jibvpLHnkf4hLGjPQmuZWav
I5V1jwz8688gWtX3FmcHcsv51nr6+LR5VxNRcRdgx3v2tvF8UoTPyj++fnDnQ1Vx
9aCohiddN1s6nIvb/c2rYJTXYx3uyzpmvDRQzQssdKKf4TH6oju3lKh1wjsqLCcg
1Z7tsMIwzd9XyeAjmgrQ9bfwkWU4Q2TGuT9vUXU62TBRBck5cAcurTbBq7uhM9PJ
4Lfuu/1X5HguK/dUnAXlfoBJbueSeJ0ilZjxzgqA0Sh938+gMQhGycFGPNio9VAN
3akVwrFsdKtajivK6dGUbRPH31WGdUhfnp6NUV/uHiuySte8ghRtds/b6vzKc3ZV
icOqrr3g2H+5JeqSDVgYuYkszY9nJ8e3Q3J/VLSeaI0W3jMGNsiieupUJKhImpod
vfgXtWeNglemJZ/kVRzfDCfn1zvMiYYUgaoaepre8PDrm0MKERg5GY9bSfxGrJpw
HxFZYECCWPyEzmxvHhQkifxzlqBs2uOO0H8VWzNZpDpNwc4j5+jeVqBf7bHDLOwb
Y5mJ+BDlyhajWop38+NsSicWKwJdRP0zxSvZLG7t74ptJqWIhpGEgUrd1oWL5ylW
hkGGGV/8CZYCsPJp8/I0MlTY3nfz080ztVvF5JDJNvK4NKMETy1IW6q6v9r64tGC
M2+F8rSTZBHfvOIVLrsJqj0WOv/sTR/OEjpKcT+nX/QGn/1w9eDw2I004R+0KLgi
qhbFsqSRAP13W7rkxtfdmKuawX9+4Jo7gWDxIBfJ/hq23O0BydVELXqbOH8h/tpH
Q0WrZdwDOPwZbkLT8yDoGxGM765szNauTXOqbwsi5vqpLXSgKWs2PJ/gN6isFXml
x2ifQKYtniMcrZfhEUohpKx9X637rl3wvs9ZNM0ftglhuE28CBu646LL/ssJnTAp
HcmCAWsqwcr/vgLSWdpW8FA2Mr9JadBZPW4J9kaM0x0oDHi0gwt6j1/YI3hCX4Xg
HlDABNnPnp8XEdmhpFnMZAsoW7m3N5nmPy6GAB4t8De++V3Aua8wzvdvqX9BWaJX
V+fSk9TI7CYqt3JuFwcq9YVVnUA5BUR6jQt0qraE0TnGDqzzsBJ5XHJ1+y0Is6qK
f7iBk/Rd80eAQX6zHeizEJ7VGgpBkFtpzhJ8gP9mKAruVGqWvcYS8gmmZJi2PQnY
L4fiwoAaB9FzKZdZPC9hRxv5v55eU4KwucvoTdDYgedt+ksNsUdcgZiEMd5WzRpJ
K34jTbliGoysrPiOjf4lr5M9Kv9DqxfavNtVjc2ZM9W70P6iTm0+BcD4sDO7FG44
rkHaFMN3Awr5HJ8PRDv8Z2ej600at1dNFKMk6nT2lPV9+RilFZfhWPNNoZGJ3v4w
MoANRqYnppgCsJIFeP9STikJGNpqsI2NXSFYmviZrVca2iaQ/VogCCTcND/T17uC
Thqu8ggDh6iLIt6hxcUgUAvQB/jC1JpWN+hDVYbALCphtnGxJYAWtEPgDzKzbi8l
eGfld/3Sr7QIdeVvK0fXHx8j2/CLrnKQT/GUDyKmB4NZhZuXBj5xnFA+MyIU71Q6
5kADKZVmBrczdsk2wUzCG7UgV6hn+YY1EUJYxubsLphTXz7eChqSxAt2mE0uLe99
jctHTfwR4bLVbbOA3/hw/ykRJ/I7xjrKBMjAVlzWgFtWCojTp0Znii4rZur3jyk5
xh3thM1QaStbbIb4hOLf7pq7apBRfRHu7M+Upzd8MfZ7BIyD0HhoLAgqZcoqxZrj
oCsLnm1oapWlvCjQ4EJYML7T7UANv5I+TBLGc2XeoydKi4fi5zRE3Vc247a5brVv
BcamjSO0cAiuy/AozIP5FrisJg+TFAXHSYyJ8cc3KaefChRLTzB5fe5d2DLE0laP
a1wM7ZeLDXu23BzzHznjZ8nPRLpU47QIX3W7NmEfdpxj+hCbYOZS/P1W2rgtovvJ
+tdZcyJwnzi4NLo/3MyOd7ZoNC8HoA1L9xJQmVVSN9GAgRzMMofzE2yks3pC/+K2
S3icUexvMzfwYgwo359PRUbSBybQ3PQFNWfZ/7m1tb/8tOluzjC27N0Pv1YCDkEt
+lqFOj17lo2vWuqdnP7I3vYgfHe1N3Td3v9m2w6O6n/nPzYcjNCVV+/H/Z9QoX13
GCAtrIP+m3mXIyirypP/g65tCFNUkZzMNS2+LS4U9UwZWIJDhS+weOnvactIVNfk
rUNO7cOMd4x9lUliRxrBEdVkAmF6q4UA0p09CnKHCIwCmV3CDCPyD69MBjOzU/0x
ZpByj3+E7zVhILhiEegCiX/iF9r+iec85BTFWqIuwhh8KFeAdxPnrL3cZZA8xSeu
k1F6sR5T7cg1rhkwLYrT7a4ogOd8xHRcAdXaSsjp3i97DTMF8j+s4W3bznS1TSjG
pGtnulUeuVi+zx8LgQmiKDYjZbVOLRfeosG+9mR+LLF2qXYsNggsQQ15MRgFV5eb
ZT+5wxBQrNV01YtOJRWZqdZMmiG6iWagGswIWS6t8WtlA5n/d50hXoC/F4HpZSLx
Gp4bHjISKjV5hiMw25Joy253kLBFP46X6/kSKfED5HUifoLl+SM64BXRO9kGKKAe
/qnj8VFHnGVDjILBSUvJDS1xSTBm5qo8VagNIGQYL+ITmuMNNFM9AeRVKlbzp9tS
iAQrZ84cygMtOoiCV13oFapzSJ/IPD/zzJGAskQjqTRQdtSBQmuf+yh0x54sAJhO
ukl8wjJHNugwhAvtqtn98EoEnKfMb1kKablJprrSuJ71DM6fldWT9Ggw7f9tLlM0
x76y+rpM0fx7UMTvXtWIX1nlCrSm3bM1IE5HKp94LDmp71mimWZYnUPbF235tEOz
jTOPkWuSAk0vCL9h0eKig/SAYjHgAkv0BHs+8KKHf2Hd4ohZn6G/hwklYaDMbaGF
j/rcrYMU9xKnP78bJeBAhnWkBd64kcg3vbxjn3HjztwfuHoHXoYWPHMS04PLSRAH
0AeuY2LNupE71IpCFEXb1mIGY50LU+jMOjrX1L5rOqfPX67ftwep71k5BKzqAQop
eAkQ5FqPleUrQ05gxEIGleAi42wwJ0h8wTkodssJFdOtNkrB+fbCNrkRA+x/dpqo
DIiM2fp9dr7/PPIzF+/uBR8XFzfGKy6DMmdrzdG205k1Cuj47W3M7H3GEYuyi+fT
PR+w6gluZnSox/V7Sw6BBbD0ukyaxEb2Nrn/CgpLje2R8TGPCZrovDVtEVt6Bcka
HMgpYpPqsE9FBuvUdTk6CMBVfvb2pdhQIsZOFlwrs6Kgp1COTyQTMS5LfQbH+BqY
haRpaUn0jfHowFCTWaSW8rds7BiiVzl7SO3HTBDVRTsXWJ9qRAU8x1Q9gZ6RaMTN
D0Ui+UkcOR2xnKuOkv/StPprDakgPBOPB4ne4v5HsRQziYAyoyswQukZmMte95D0
GO34aoNQUZB1qKqEskeHcrR15ZDMJ1QAm5erWedPM5He9InxHCsl7l+gMAIFwTif
a+ZFiqDC2LuS0ETxzxzEDcoigur5ZK39mfqQYq878FGGgU7/hAnBvFtEspO2CLES
r5eYHRTIpiFZNtsMnXd2TNd+whd+edGB9H9w0gHp4oVSyv/Kh9cM1YzqxFRIKZkU
Dfih0q/bwzdAs0vFXOkYb+NdwUK9Pxk2M+DvOk0gbgqcY4QgZx/Rrf8fYIavwYKW
ZfNsXARVHqBlllsYXnMpjufntXkWAnsxj3zIRBq1/73bnj5yKWFIVu5Rr5hHCW53
dv+1IqI2+66IWR1vevSuKXJ/FTQ/3aDArY+bHKAmIyKCe/EFjlFCqaJuNYvIJtME
mTLAslOCjBuXfktck5eguedEie8ymO34edMicvl2+Ms9D15rFiZiUtPHzv7IHAUz
uRnoTa64u4c14NVj1jm8EUwykYd8e89LrYmf+Yr9q+OdRZcowQoPYALJH/XYW5bh
Hg+n0sF3llc0CaRTiv25b4k0G0/0Yj5ubdY+L2dlLvugo+TAUjyjWjqw0bho3fBF
79/oA5R4s4/eOFNbtJs1b+uFbmm/7kAl3fueULV+6+0FOVYSHhQUHELIq8dpJ4Ep
+GMkAzOEHPIb70oXT8qJnMf62ylXiAcRpGIvRd1sjG4I/qGMiLtuAAlUnaqZ3Hn/
7WgjOF98bs38io1yyBBYPw8u+sUORUaPu0CDbkP5bT48Zjk7J6P/bpeGvHUVhjeZ
jim5d9nA5G7R42Dfe7PmZ1X4Zg9EG0YDN9jYuah3yfc8R5Ju4EIGMSGrDOHA+NBq
F8YXgNijwmqYN6ldzBNOsFR2EakU9jVXD7r1JQcX51RKqhU8gz7hYwARhdtIpQ+j
tFArcfns3xmCHXO3GoDGEX5pdTY8crnYlWMbet53IxNdfCOI2Ia80yCotbzlpilN
mVj2vFt0CLfuH5kANDllbPK0uzrlA+chJ/8pvwO8UpOozdFxu0YPXakbHEo4hkET
ti0D6ouCikkCNctpkBYXVSW0syK7unmQWyahHYVPHb65zLGh1z+t04E1bXAXzLc3
vaJdiGJLfel7aPiGwpun9mFjlkPj+Tdcat2Gy7NzYWyPgnb2w0bY6qbUyjMtxfTl
7QBBg7mugngV0UT191mrsvi0mGjHQjztRuN1vz5M18b5FBRZxKJbGTRscuyUPCmn
/RxPpuqW/gU8zgjtokBDoJdn+aswE2pTTzU+r602CQC/XMdXaqWORXArcvaws8xQ
vKLBMTfvbAo8EmzPq45f9ooWCKjbPfKIK+AvBy+OZJSvS7C2JkY+M7RjHkw3yGs/
Onl71EukxYyIqvmk4cf+J+r7PuPTb79WEQy9LPOWSr5cms7ZEcEkvIn3tbQw7MsJ
KyzqpW79N0nIUlfL2qEioe92Cw7KJXgIRVlViE296tkOEsCxQ6gQ1Fw5q0FhZaxV
0ObOz65LfxCzkcfK2wPoe2HADlJfWyb4QtIzN96Mm0m7RVqYszfE+szGs6yAKfyA
T2RV3Qgy0sfIxxY4Nch7y8YGYGAcSH1VfRr+Gv/SGQ37OEVaM7eeN6xORMvSM18O
3YAWGPe+pRVQSr1yFFAcYhU+iS5bTB9HgXWihiz01HeOhg32tfr7zLBDjpEQiPXf
uQ9BUNk8h6G2tK6JWFoldGpeAYsbxrm35GsPk5zOUFzFspABtsGTTIg8w/wKiKT9
dfxKrkRwEKuUrIvDC3lBu8v+HJGscsXuPHjDntlf98WLGSWxHNV6+xh96cVOQ5Cw
CB21q5TwHlKx7ExR1T42WTTontPfv38Ymt3Rho/jQDbH84KJGkrCdyK+pWKkK44n
yFaJoeDIGyIIbQcBpPP6yAQBrT0GF9h/ybV/tCNhpqr3Ju2osQPQTnOYt7wrEiOz
REKA2r7Qg4LYeGrLr4a8JLiz+YLqYWTQWJ+tMCvgEX+vurcuAnGuW5sGYZKxmLxQ
SOKpWNSC82Y+DTlPe2BIxkCpievOvuttsxtUNRzs407eK0vsb3O3obx47dd4kQ4x
mfBHC30Zz+ECyFiMHGteiWp3/nn6TttXzQxrsuhbfco4DQr/1Owr7LN1PO5Vuvu+
iJsb4ukCjvBYsfr6Gyp/XZXIP+2DSa/OBs1Z0deu9QxjB1/dtiBr9yoNhpRTbGbU
Zz3AlApJD7zoB7vnKjZJ4a7fObUFdswsHdfXo9oix5Dbr7A9L6HXj5S69WT11Tb9
Tz3h+qF2CIXWO51hyoTZCfoOTXDPUUiIxH0jV3o1OFMRax8eT7+nd2O9+H7m3nva
ZDgCSfCPOVhA/L5BTMHWaXlhVYM4MZyd+02vPtOdjF5zCNbpV1rAvhzULJufPN1b
6QL58e+q1fc+ZdguCWXYuXbg3VMzpqAthODfeVWIKj+jh3x8NCXH8FGQyS7WyuEP
h33NhxN3/8joQd+x+oUvOFtlUg08BXXtzKwiSB26hxi3h/PXhV6iY7WC7yIWVcXI
BzY8d36wn8I1FlXa1n2F6EOIG8CgTxHjQsonBJLWh2Dor7mU34RXfIvM1ruLa1rc
0qLRd73fp/cS9ieJB7OdGB2u5Rkdeiumro0pbsUKiqC0/E+TT6Fj6tuqSDy2toxR
oQVQlZhstr99Qh3S3CQInwdyY06Z5YoW5GUNEWJuGtrxiNXY4GTwc26soioDHzCZ
Lw9VSq+fyVK7DwCDhwzuNXuHP3G8pyvV6r4+It7wRmBTwLhqWwwwbKtqso18G3Pa
clWxU2rCPseARgqUwv8v7g7Xumr7EFasSUTd5n71l331DZ/0HSWeX+XjTxsvDDzl
gmrOvCTptCr0YK/9/4iPP3qeUiBWCrDtGdXuIrd2HPpYUYWoPoJFuDUW6UBMYg7P
q6++ouV8GPUgrtKK1y4XRk9no9B4ZUsLDZq+tsEczZdvh2gLf4DxS7wTRBJ9N8OD
Ii8Mir2VBV61l0+xvq7Do7Tvxf6J4guXwRMyOU1ThkaJEQcaL7uHIRb7TOJTRsRp
93x+EVrS5e+eStwjGPoHv4yD9hRUo8I/zt32HHgfnBwZOImJSsNTdnuy+XaJXpxq
nVRywazYzFkj/cpHDtRAz139hauqR316m4t8+TE7+PG+9ARDAfS4dyY4ICdGLUxO
Yql85SHMIG6BvoRR6y795C3uE7g4TSxWiRcNv9w7UiRSuDMiTfpAaBIAa8I96dO+
vVN3yFZ6QE7wVzdMa2XB3MBX8I1WiehIHLfXePjYzU9g3nOIPHJTH9g2cTu/hAnD
tFwgkJgQNhhvpiROrqmpnzSO7+IlqgUHcyhMQC1ujhfIdqGxHbD0Es7WnnMI75MI
0QxUp7YOoujcHNAGMotqaRMu5tbFQ87U//9xwqfaAPrfEdeLRVH7xD7fADb6CCxp
Wpdo5N+7bveY26L8sLXxRvoCDS8Za312ca7iwXwpg/ip6V/ek0I59MrVc/QwJTed
RZkwh2B5UCtN4tBaLa4nMH+VMiE92pqIq2Gt4jv1Qq9hkvD4NXSuFyoxe7CZ9cEm
omyQ7A/r3Ec2zxT3Fy72v28jiycK1BblgK9XEmXqikjlVyR5QtScz+mSAsVPBXhA
hLEp2ln6k+FuyZZahSGAfN55HHljdAMrJRNFMwV1pYzg/jblB2JCeNiVUoRqMM/U
ZTITFFAM5tkNfjbdF7aQsdne2YXMhVdwk4g45ygQ1ypbRedA/5lKxZKiySwA+IYV
w2jW/p590mvCOQQ3XV4nFdk7ybyD+Ua4zK7YbwYl5oTERRp8KQOjzarIBZafPI1h
OC68KAX9rUZTIC915ESdHH+N1dLcrIOqF31Mthdh+hqqthnru0Crv3cVNgLKLIM+
riPwNNBvcO9YKitLCbHBBM2XTkgbmAx0PY3dxJz5y2YtMB1M06JpZ3nR46B6kyJU
bch+Gkz6W7+ko2MHgs4WMZBcDvQXyoolCkOGNJ0G6wabuarl/skP9PSL+N2+jAFM
aPLv0dquc3u+zvFi5lyUt4MnALHAOXZZPABUNGuZF/Fz3iaPxzDbHcAHZ/bN0FK5
SpY7NcMgoHkN9hWXfcsk++ePRcRXlUQK3UfAh9z2pFE5IER4cRh4PUX37NhSCC8B
b3W69h0PjrPUe/406Q47FSh1DX3fmb5aVpHlFlfWk6Mg4+Ig6vvL1JStYSULy3rE
WZeVf/a25y2AeCCUm1Bqgs9hW6r1gyNo5uKSUvCtC6KKs4Lkpap4vtCB8CBxqd9x
IiJ2nEOBO+061kgKg+gbNYml+Rm/bi6Lk+r12diHQronukLIsE8nSTGj3O71a4k3
33pa2NOCcEHauIZDLWdfSzK6n6NATEjTCmCfyiTysSdHrBilK5O6rSycsFRbQDKY
ERGK0UTV+t6lv2nYxGORMxGti6efNkwCaF/BZK8t7dnBcPZcLx9W4MrlwGSTZXpu
367GDxKCefcinBb2sKr/Fv9iouIDBqfKBoo+CvJhat+1nTm539SoLpxbbOHMc55x
EhjZF5oz1c5YLmLuK4SN2RgWDFyQifWIWdD06vCKowx/du4KV9/SVUL3SJT/dskA
AhnPs4cfgUDfWFCpzPwR6vbSulWRx2+GvjExJn5qpbKSUEzSzAVbXJoxeKOMPpT/
A7OnPnwMCvNGiVcZmuvDqrFbEdBFruXBr4vG/HXhVKWylP5W3crNqaYMFAY7PpXx
nhjvwH5kQ6A0zfIQ1cg7kPdJyNqFpdnHBTNeX6luUwlgkkYo1Zoz/5rCElmdLudn
WY/8aqJpGMvomHwf6Q+T1b2lzXJ1or1sDRKIu4ugNxPQXTW27WEBi8rZoPufVqhs
2g17fIgmFIHC2mbL9qROgJEdphI/W/alOnpXoNyxfMBnlNXQCpCznqWYPwkDf9GT
Gd/9M9aTZtFrF36MgoPJTJRjtpkBoX5C4RU2VnxigiB9W4prpmBXYZNfzu+oKTDH
VJQlr5D2cYjF1iY05lX4pje76Rwo2pwQuGEQ68sEXw9sVBHCwbdz+94M5RAeB12+
a99E+G33Dvnw0ieWYUixzaufdPF8+rin6+yEP/Bff0YLxzZ+WFocSCXNeZsqaXdy
xbkRDUlKm5UEdEU2qQwTyomxoV+f0OZQWsWxfbi2q+C4DKaHabsR26bOOOTzzL8j
vniPcllDjAuKJa0oS2sOaNT7kUiYqTRe/3bwKmpp4rI6plA+pSycrA8VNzxlWbA1
TmN7NFl2LkXIoQ6qBjyTHsjtV0v1934pGvmYDGuk22GDUKq3vLCSa+uv/br+uIU9
QotKLeWO2a1x1El621ysHKYhjyAFwaOVdaBRpxEemFv16nXTff5Aoalz0A8UFbtZ
fri4VhZXxaJaJyxENtV99gcIDTHVfAOGpxIpi0F0Pia2pDxEm4VrF1o5vad5rMYf
9G9haW/fvWj+iNuOrOtIo6iCM83KVNxPktgorRiOFiNAFk9d02Pti/OOuj2f8cx9
89Qh2AiypIUBUBgYGwhEWRB8jUMLh8W6bLtDwrpUZvMWDAmEk+E3BhUUSf2RMG11
NeH/EQ7hhmHwwHwTCGjrB4c7voWgA9d3iJSKY1SsTmHPsn48EwBDLw2cXMpbrwXg
PCm4ncHvgK0n1pxCkyrMDYbu8R49p7LZCZaLuBjrEZirHtXHyAnVVevzTK5Vh/7E
0ifm1aj5h2wz1n33z0kD3denYChctq+0iyfgHbZ1B3O9MlrwtBVd1muWI9S/xbxW
B2Yfz6OAdM4z0TU8wQoXVlPQo/fxHF+D0K3x/iL9eB+4a0H/L1GAvUTRklpztv5e
RaeYEejVPylIRS7A2ZiNL0/V4fihJXIqh2GWjeEqPXRwRhUwONGMo9o1gsZyeH2d
ZiUj+6g4kDxfc+1U9I0bKYIc2QoDBiPE1SNT1Dkpf6iOWLnvHLbl20k7y/0h5tj/
LUnC/z5WmxRNJHkdiIHTyJF/gNKxNGXkAjP80MOaaIp9gJ38SjXfA1h/D5+UC7J/
k7p4nQJS5YXn62iLwj4VdpHH08ub98G3NFWJEXbe6bLzCROpkjL3yTcrrx8gpdG2
Vcc7kYaHCFBvaTKpNNVbP6pfaqJL72l3a9012rFvlk9P2Dl0qEnscxNNlKAuLl/d
/pF6IZ4BssdqWBF+VFLAGlukvrMjyFKJGj3hCv1GCDdkJMJnKnyypTpwEPvNzBw2
TDVNn/SJ84ipb0eiIzoXipvrV1wPo0L2hs9Bd0vH54BjmoyKyQ8EX5cTHKdD3xB1
ojQ+6Umept3pjsaIJDUa5LXc51y3W6W7pSU60KR2x5gMhNIH8iaIT/pQhQl2HsPi
97c8GuRThqFuX0VTBne5OfqIHMxWfmtAeWNEclLn4IK9APOt0Gyee1fa92OXu2+/
Bsk4YJFMl63bzsh4n6xrkRtBZ3NAAwTmfODcdTagl06+iitaMgzlpeQ4zw6RgSkF
tugBaAs/1GdCt2roiJgWCFax+Ov6mzhyDNgj0/9SDiI6C07p8Khm6uhH/zdfp49N
clXJRznDnISWElmpCsR9YltqHdvHY1tHBFgk19HqrLOFP7H5f5lIFMdauWqY2qNJ
WA9OXyLQtEVPJXa1Ma1Td55nO/M2wMx5miVOSb2txFWcDBvsscK78ypZX0iikzuh
UHaDqaK/fKYuRIdZpVtVfWqdx8SoLbzHfHei83d6uBDKm4WEYprpMEZ0VPenZoWn
7uoStnTdb5J+j0H/A0fzfHSxHzkDT0v43ggbwvgW+c6zPs39OD6Xwxft0giWK/Jw
D5NKmTJxVZgRioOYP+DnSKGuMxeyJNQEeqpEUbNdPES+FNfGwKhV+6izyrgznZDc
K8Xe12vZJYumNwhl3ryCsQ5pXWdvg87raFgVda82T7Kw0XLMP4xS4kQhFYGrYd49
Q3uuvu2mfl0I1o/b+JlbUJZ+XaRhtxfvQjtUUWOEhD+5BDNxr8ZaNW4tL+v5uvyJ
qM9pdNRPNEtSAniPcQ6b6gvihqHfzoUeaGgsLShihWqjcZwPlRrRcCfhY7ReLxZ+
iRYN0YePfq3suyzNhaXuzPLXXPiKo1pQT3D8hRTxh6w5wb7/ly6PHS/Z6nH56RPZ
U+8MITzN8tLKQPC4uGoBlv5FAuF9a7DbS9h8BcVWwMyJ7XOF9dUqlXFHfXk0ivF4
c3KUX5HW1CGooScK66THLPppw5rmhvMCmC4S8yUulG3kDcTQkllcNq4wUx45vC2b
q8bvA2gzcDB/1s30hzDH72Y2sQtQZbmH24Ck/v2+HR9kLCahZylzWfyL0zk03mb2
aWKuX1obNgAU+9wKOb1qwGnSIKu1yBfJhHMJR0HcSq2lQI3fgUEb2t8RkoLf63nH
4s6Gxv34JtEA1bI+QjwFgqYDkJwsbNv6bYmzkrm0w1Ykyq9tLe+YQeHPPEhGssPo
GxlPIzoH+fWrDezDuyqFeDjFw1eZylLYNby7KxjaiPCeHZ4Z1+8aYbIcFk42vPPH
ONdfClxcdGDmrrA/itIATNmcuBi2HTNgS1/LhRKzkrg85NGJw40qSzjS1Gikg6qY
aq/Mfr5mWyioeZhdkE26KxDUo0dlyEWEYvof8WqIgADI331LjCK0yMcru3zG+nKI
E2oXIXPpsVoVamKifAUhf4mggSty/f43muUvWh97c4vC8sbqWk/c3KAowVOKiP3N
9fVmDE8fvjn32zbCSGXnMCKwkwkuKjCZS78+SganIc/a9O2AqFS8XnUeu3W+yjhG
jIAYyXEEZn/0tR5oaIIqRgKsVAMyiqbf/Sdcdzt96mt8m6MGJMvGu2Uh+8twLQ11
tvd74CHZfW2KvUEiIb3rdOtbf8Vg/hdR7ZehsBahd+aYCofFcVNOZ/EPzxWmpBKl
G/RCe2gVkKViqdOtb25ux/zwt/bPIquWB5D4UNOZFT5nEMAZO1SYUG2/yQ5gh7cW
xgomkHvJ+8u/tox+aVsRcFnoQjA19fgBd20XdsfVyYfxUkhMH2wQ6q2CdvMj/dLT
F3xxBCfJOwjFBeqY1b3zSAwbqnTGx6X6XzBg7WzI+vBSn9thR23J3OOyTlbmw0kq
NbM65lGSKjxjvM7iKzOKLfUua/O3/ZvVxOQ1AErT2PGSeyObvrZpMASdKSIR6cpZ
HyUl/roQq1kLPPlSshAIPoWgrvs/TtuSa/uRzaS+9sh6y36cp/CNFyI2FtjIoUHD
yhNKdCzoK8wiQsC6SG30FbZgnByCjxUhLWfA0FGenL8j8zDF3xv+lzX4TC5MtiN0
GHSDec1I13RZ7Ixlh3hA/gyg0uldt2I9rQuATUekPh0p6grrF8HX8SjrsHADIpHF
+5MgxcDLdKVzJJHCEsKlkjipHRipyVynUH7+j0o78gKvT/dvAu7BJVMDXI93NquJ
dMO3yFr/3EnIyeEMmqVWUz31Hu9EaHVafLENpxQfIU1nuT/qiPsnCIrEBu7oZ1vr
hUyAB/u2pb+im4/dN9m7djM9ykY1lgeO1oyviBoJ9aEOqc9y/D2/FTcxrXLnnyqq
0PX8pio2I5GnigsFiJBP9sbIhP28DzYZMQiDlXvmAhJMCBLloPixWW8MtWh9s3bB
Awcvhk1Sa0mhthQo31n/cV3zX9RLdejnr+Lvwyx/VMsyzEcAAck+5f0nntyCuRBS
FrS7fK4fCkeZR7PZOeEwhhScv7zocpH9CT3KFPG96i0XHTnLYmhNNFrY8SzrThnm
O4TkHhE8ILg/EnuAmzuqdw+3amWzNbxeIStAGEAicvD89cfiSS3TTKU3DKdXfSax
TrT1C2asChDNUdOHAChx/uYjZekZhn3qFmvodktkT2B+8O/PiOyhO8+jEBtyF4yx
eb0UJp46YQZkd+nVfLEJmDTMoE4q0pKMJKSi5sNXXOLnHbgG63iBuS8nB27n6x8m
WN9kOcW0YpSy5CO4kp04Az9A6Gw9MhtemA2b4RcypFqgWmwngJ3iNRUiNZVsBBKT
2mduiJrBf4T5l2aA+bA5vBvlK9dPoXakjBwyJIRYkHtLIOC39f7ZoAbIkItgzGcz
eie8/R8n5i/UuvD4SVx9PhnmQVYVpyLdJzaV8GwPsmUDiq+4Iumx/17fAS3Ka1W/
VUsekDIj2iJn2bsL/pv68NwN36NmMFQ0Ia3F8sGNlFq7mHUfJQai6ztxpe0vQ8Mk
L8C8HMZ0O87U1hkTUJyWWRrI9h++1nTRV+WkzqY37Bvq5gWHtsAjX+UqtKLph0aR
pN+VUe5qHxw1XsOq1imYc+Djwu495roFDeZycT828AtsH7Qj2Xc8s4i5eXt0YbQp
KcyNQxlx8guM9MKJdaLmNOcuhTLBGGIF1oqqlBC0CPNY4yuBB1er2n3l0OerQDeY
EZBHSj9n66OOeZVxESKtdgLEadMeL6R/rjuvc6opU3PI2AngWDcfmRX50Jq78iAR
LtNdg/5DmmdctM++r9aGMu91uIJW/Cx+6KnbMQWwxnxEb2TBwMKdC5JLa4Z/U7CY
OV1JZVt8pCCDKnMWl7pNFMWagr7ytZRytKspEWrtNLHPMiK+EMoPCbXHouwET6FM
XQUSJieH1Jwpjpty2c4Te6K8YMobDbZhkI4T7ZRKmuK2cRD0myHTp2Quw96Jia9L
DaR96Ceg+fZiUFwS/dTsdshqhwLBkFBDuYPkCQAoweumdTdCDh7npFSol2vRe4Ni
xT3+xWLPhDbDuOl+7TMKQtzpOwLmBEnOiBW6LNoiktXLoIny3XvW8VE0yC+Wr3iD
taHeIjLCPOFcVopeMnHWGpHDDfto+QExxg7GFxEkGt5wATYY2174EaOftdDXtLKV
YVOFHrTmm/EO5b2ztfwnWhF2nYgXzb1Wo5jfe9DBMpkZDnF7PZnI5FcjS4SRSA6R
eJ1D+ISRIerNkLHO09YJH/am3a9VCZuyKoNWeCGwWsWEluqz040iisAtgP5cB5Go
YARyDDqoK/g4lOPPpDcqzLeHfwrt8k+kh/oESYxSFs9h8nzZr8W8OaWRtuwhhLmA
sFZCfZyII64/cnj1qk2DuwDl9UFaOVXnHyOB/dw9OnzUsrpeSBkKpo1yXUjGChc3
hEPJzWrqdSpul7IbF7J4GOYVDwvGWhcV70pZAlAv6hIN8rf0gSdEeELnD5ror7DA
ykU7P8lMaBa4j2vJ3Ajac5CZvuAjdli47VUzEqCNvGQBasX+ZOpmM+jA1A9Hq6gc
e90Gat9y9yJYU6In4PZQeI8gcokHhSdxqfXFrEVBKVXXzcoMS6CLnHlexggufXFn
szYLrznwPmRDzBd7i2Y/eZcG4623iJNwB+L7+mfc8xV9D7g43VCnve3OMp6BKI72
UL3G3TvdrIgGVVmVzDnRc7rC+gUFheYZ2umfWOLynS9xAO33Hn0YtMZVTIthL7D0
NAI4bGS0ru1nFTSxtSg9cnf/xo4G0mxy5CLAVxQ3mgCj5f7b3JT4//Rq2yQNWDq4
3m+9+iC3HBvArShWudv5ovaGv5r1AURJ0ZBNfv9VZT4Fs4Tskc8cKwMMbZ8Q5oJP
ZZxqH3WHtbWx6QoGOwdjJITnjW+P1EcVwdjcwtgYEIA+VPI5DOVDd9H7uSw9ZO9L
jKYnoQilMfu5jJcR0rBWD4ivsySNiTckECDnUZUg+SU+WxZTq1AukZ5mPJlccWqs
sZUj1mCt0wua95RP1PnoR/8tG44Eox8sKxpGB+mwyejubUoF1ScZlR4LB1CSWhmn
3u6IpQAD9C9kLCpIBKvBGu8MqdKR5mhIUj0DBxZnXlwPTxbRnWCadkQH1z2F4iEG
y5zF4o4o3inu+pgZQNsk4HbK3sYc7V1v58C4tPSZmzJH/ggBSGK2TfthDT1v9Znv
eEQNzFeq38tTX+S9Uc240QuFhgyAK+NEmdlc08Ti9t0voHqPQTRBCQ+KYyyDuvCD
oMPEAA2RX2P8IrP7PuPV25KBeUFf8iHE2sDsMgUxou9tNPRU7LwukrfgeZwROQb/
AhcQRUBlfxby0dlQLMRA7F/oc/pgl8dhDVG/9B42YHUxCxXZaiIvG31OKaWak5a7
HCalqfF4ksmwUC0K/QyCG3VoMXGjExEOX81+7z4/MSnIVTQ49gO7DEKPrGsXxkXl
lHjbqbd+71+38yNCcI7M35Wl5dhxGQ6xTgJeV23/mEK3D62rzVnugf4yEof5t6iW
5WKFtaEjXP+cgR86vsqZVg4Vkxi6T0sIdGraOcFhjUT7qr1eDwe1kZFcU+S2T8eG
VDw+tp0aORsvQdi6ILVSASf02vbuFN9Z1ZcMl6BD91cdg2LKl109VA6zkscjipW0
2ACmD8ese8MEzAex89k8KrnPHkg7K5B6Nb7EGmMDRq9TkwikY8wI143RABbOp1LV
wfMVubICPcds+0kdAtJFxIxl0/DbrnuIEyvqeYvjbxoH+jWz64RYTH6fLo3bNqgs
C2DLcsSn86OhzQuAdwbNMP+TKT/W7fQeLmJ8FWamKo35m8BoZW3VJDPdqcqwUKR7
3hHvg8ZpNIXeUeYsXVY37hJwqexj4H6bA9VyR11K2Xb2/9MJBw+US+c18xnasBTb
gpRsxuv6k78WWWdxF25yaXEqTlxnKDEsLZqPLNOCNqDu5A4i8kNXWgpzmjMIQ58D
aF+GaBgnEWXEMO4U3V4TyFysSrUUtvDTyWzimTfd80N8/0+H8SomxL9niKUMqEMD
1KRT0XCOfs7DSwVquyBcsCKEMXYUf1pHWooG4NszjlnDnyCtJ1l9/Qnr+fNNvXGN
nXccfwzB5v6zReGCXriZ4EPlT/Y5gH3SxlEzNbm6jhUXNcmacJ1INqji+l6FtxHd
rYtj8/hPNz+yhx/e9ViBH6MIDYDJ4ODv55xL9Mw28japRw3B6ZgotPR1LhgIxVeB
Bt9yuH4naudigPYXYqQ4iw==
//pragma protect end_data_block
//pragma protect digest_block
gWTtKfWGxE+t0AtOShb1yEKwIFg=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NKGl7IkkyuHL9c1Bg39JU3IwPoeW0Nx5iELYyP5vNUgMv+M4otU9Hai9BimNtYvE
e2qpb04ScbiYq2nbZs8hKYaCxGn/fgDyy2Q5GqXKisRFfTsXJPp6mR6EmRnwEFyU
L4ddnxIk8JnRPgnV2cWqLBCQQzG4J/XxTxAOvTMehO7eUX/8NqN16w==
//pragma protect end_key_block
//pragma protect digest_block
JFB5KDYdVc/Mq2FSYuPp5jY0TpU=
//pragma protect end_digest_block
//pragma protect data_block
n8KUjnIMZ2efCU83GLE/NPBuZ3++q8AOWt8J2REUkyDXeuA5MXQuTA10UmBS/t0R
yYLaEtlvoOA63ZohWfmT0Bae3qckysO9h7mToVnP2qrJYmz0d/ScBwPrRqaCcZsN
72jmfZmro2F+s992TKebGIryXICWMB3Mg4sVoP+6B91VGpJ5u17glK3RLoAQldtk
WJGH0Qha9IxrnlFabKhX4WlI/BbSH5O44zsjK6VP3r7kPfB0KOkbrsgiBHlLg51+
U1C6cH7hhQYnoyIleKcO+lnWLVBHCDFUt4Tj//1/uzzYIqbEFzbLNEDfX2IP/8Vt
l5dnT5hsouvPvanwdHQ1FmS5CsaHBEwtMgig3JOnEd95ucxNkmm5PRwwine3KUHL
YcVT4DPoj9iA2uHgtj/0Qs8OhO+bx5AW1d7ZXflPaI97VOHxmgLEy/LE6IkJ+dYM
/Q6/cV1cv52neSvjCU+/i3yQQSgK8g4q+90cm1oi2hslKsP8h0lqVkBGlgH5igsF
ARrncDKr6gYGqgn9Bmg6SJvzyhaaptHZvcVnse1z9Ielbyziajz+OQtpCAYRVmSl
Snc32EaKJTAna22ldo3NoCFe812wDySmltOd374PzG0erp6S0vT9TqOUfQzo950X
Om5XhtAFONzq4b7ltidN45qjdRjmAYHaxEum2iWLWAEu+bpquN28NUJkScFyVpn6
l/FNRlAyHH9V+nXzbYLw17+rVqxBlS+6xXm3Pe3SkHY=
//pragma protect end_data_block
//pragma protect digest_block
nHCnSjV/b7mATKjU++5wIP7hlnc=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
IMbmDRSM1wu7fsodcaMBLrE89yjyetNdYv8zgkl8wmLA2lGMbm2W1Hp5DERHTCpN
Cw4ikrcpQCsy6pG/tHleivncIiKEsfuUcThBY629cw+m34IA6jLA13M0kae30x9q
oxYypg6grPA7wFayyGZ8Za8h9eevKdNudWuw4/WEHRRiE8WxSH6tQw==
//pragma protect end_key_block
//pragma protect digest_block
hrTBPHEfmWNdA6YkFr5HTNhtgig=
//pragma protect end_digest_block
//pragma protect data_block
bJAX0BS6EWVvF9inXI0cJCDJCP9qJNJ57AjUzLgCP/dO6FAKyy1pkvf+eUOzzF4Q
IdDkELP0irwdIByV/9zB69A5NkakE+ty/l1801O0XE83ptNw5RJwEUH7yFgYG5/b
gQSWgcuYXCsIKXdyzxFOCyNveVhZBZUcyZLBc1ak0EZ63QNSTtKN3o3zojId/0We
/v9ZhBf7bi8kWNVsxpCpr4UFOALvhA707i0D7lHust++J1Hs8tLxDfAcpZhtn0o5
/roqY2VURIkEASxM1PFgBprwFABCGSMKigo52TP80ew4jBab98JyxcI4jtAcSL3K
XtniVZqLRFZE6uwL30/dzrWWbOMe1G1I0Ye3hb01SOl4m6I75YGk2fte8TAwICT7
28/Or4PLwehM1YPStffE92NbOk7/8Q2Gh8D3e+yTKixzAr2I9byHCSyzzIvD9nff
J0+/QzmsgDgN01TRM87pQlFmMDWSDH9NEoVZlf+XPdjGX6mZjTZUkp/DUQhELrX1
0b8mR9CjVWhTnORiuU7k80DkVLOEg2yrlg2Dgl5oi4EiKXNr7dByihDuQwQYLF0W
G3I6C4pNcxGz6PG8QOZQdfYd0wI/bJjn12FG85fG3GM=
//pragma protect end_data_block
//pragma protect digest_block
6b8ztRltyypLLuZYFAFFaN5V2u4=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5AB0KUmh7VJwIzhm9ih8Bw5w8+jhDkL8q7dwJBtbB42swCespa7a7X3LPyaSkTBQ
gqwfPEjQXm52llq2x3KYKN4E8vt6YD4cD1K1agf8pxP0DLT8NXe/9PGKnThDCPgO
gfgAIf/u6zl/QObpSntSa2MrbaeUGITzrMalAG/ryx68eQG/nfXSxg==
//pragma protect end_key_block
//pragma protect digest_block
T/Q9b1T6js3GIgEvHMT5TjDy8/s=
//pragma protect end_digest_block
//pragma protect data_block
WL4WVStGT3RDUUUdWVAAWcSmuDSfGM1S2naykd9j6Ena6kUbutE2oghQwxTPmnSF
CUm85IBMerzKdJxuNMATKb+hPmJqxiwHl++XNQWs0hRUMniL9Pv3EmOqgSqKGQs+
Z5AMoSWPXLUXiP92ER+qphw1QBTydo+VaQmoBsG+Ju0ExEcMV4+KAvYYBXDd94ya
v3my4cSJQlSvo/Q9LYgp2Mr9oB9P8sCAP9Kd7Kzh9olM1j3pWCAaxvCHeWIjitDQ
rgDyPqkdVZmv1AwjmoA1dW/4y/c1yTAkqflAS3AueuaF8S5I0z1StRBvTeXHnO+t
81uWxbEE0dVFIU//aaLf+VGNHzJANNho1ix7CfcxdAyzbX2YFDH6fSWcJJGreLDc
yOqer+bMPZ/4JzW+IVEGMeuKmx6lMxx6moPCHE0dslIIYkeZgtPXtJZOnt7Fr2tS
G9L4CPSXuT4RHHS1GwBtfUMAIFrVcEgG19rxMdqz7ddyWl1GKYjBLcRnOo/fRJer
SohVW8hxk48l5HyU9mIx6rQA9H/2x+yyZE8UW/lkcp89aOxKgtc/dUzjHfIOuiUC
Ewe645rnHLQQoC5oJPF85wy6FZEjZVYPFvsHX3+Pdxg5kr0m7ZoMW6EZm/lhm/lB
bCSU2eqkDkCfFhPcRI5knmtu/artkcFOfdmDeKoz9dGiN9LXyk8KFPnhBCQg17j6

//pragma protect end_data_block
//pragma protect digest_block
PDqM2VKRfHPoCm1lOwF0mgmu3vQ=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
E79EW8jwazVFtd85wwVPfApaCL6GkgbefQHUtOokWU5RIuRY5sPhrg3sz7PunpyS
6Xp3HOzBnjPkKR5ApjXZxMBTfIgxXWbm8j50FUr9/sISKrsq55QEis6arTLimFYA
ohMWII5+PrF5uXTo/Yg6as9VtDJJY6xio6u0vm63bhFByg7tpQdr4w==
//pragma protect end_key_block
//pragma protect digest_block
Qisc4lgCYd1+RKb91H7eIh0hyYI=
//pragma protect end_digest_block
//pragma protect data_block
3ywJRfTfx4r52lNU6l2m2l7KHk1g3hgIE1TEoBSd21nZXKMCJMxqq7wsAzQiyuIa
lmkw/YjmeEiLDaFxyTvVCvm3TZOSLDl2/6pP211+84gUm4f5JhyFHfJol3i7FX2T
gA6db4NRcklg5gCv7gt7qxETGZMZxhcgYGFOjckw34Y10pNPWlh2+KQPErNcHf5g
IwS+cOsKau3hTyQb5JVcqiRc3zfBHpQVoqmX/sPpqY27iNmrQuDTIr3Vf8C/6k2s
tiYmMYJTHoE3AEfyrPv2+lQLXoaE2gDJE9j6KYsaTSO9OQiFLOGQraZ+ODUMOZ0M
/TyIrQiVpylk9FeuDzg72Nnh9j8x2G051MbLiv5iSZgCRVthju+a2Rh8EKGUiIsH
CzSPtAQ9kTKTXXYNpVydF3QRpPy6J8thfxKbLBvoWEL+hWsFq4Wxtg+aTpFXFPXg
MZH29VnUwqOEe7GgvDYGdwT+Sfc17Y+wFLXhVrfl4nNYu5aTKEI8tqewpyYtwf67
gEa1scHGvfaM/P46j4HAtpMb0flW4EQ8atZM7VasMKQyNKRlSVfsvSCoxciXzx9l
pa0fJP4ClHh519c+5IAO+ySUm6btXqC0U+1gFR7sgDitl5/TQ9JYHOFedjVCIXqb
9jSdodlOVgCeFVZ60IEMBv9s7rVwc/zAZnvHFhLfMdg4w5py0cYqRmpt02ub6aGN
dHTTmcEb0zLm/4IZ2q+VVcquhZOCU1Q+bF5xyb1Rrn86YOTGgFjDdhMVu8Ymu6si
yIb7PzdtHv4YfnBUEHNR4OYzL9x4qh9jNll0OaGVqC5Bfqi4aS9lmQZwEY7BGt3M
NAk0ysmD2k8aB3XtKO+ORQ1+ihu/5nTzwzIksZ9YpeZV3FA43pvTXfgzS2pHSRes
SonaNGomufMpIttYo8H+Ee4Be6nAeKf3wtYyVLqseArRjAg9D3pyFc6Eo0AW3T5u
f80eZ7eWqco06iPLs1O3txV/Veb4RI64R+Rj7n7PXNWr3+qKoL2iPZqCE9rfNek+
WZUR5DMpwkOlpfXmgydW5h1FhFAr0OWw5AWu6rG0QQbN2ia7Ge1yg8XjhPcr4RVv
8nkiIAs/qAj42WDADA+zARBqbusb2qdrnBDWsGNDr0dbCLEEa7vQNtUqCjRA6Dx3
FtbxZfuJzq09/u9wSS64zN0+QuDkEsWsMm/y4zT/A0is/iP8TFLxYOCFTIfOXKNL
A+kxZ/fbR38Uut8UZe5848J6jFIw6SeQuJSijEvKaxMlRB6xofzG+xiJ48yVGmSD
eGzBJM/sXzKi06Or0B4wMPfmrz+lE/Qq5T5mDXQDuPjhHr3o16iqj3Sni3lHjOz5
bQTRIYZeHo4WbGLJq00/xM8nfHXGJIa80t7/jxbwCbKumJChim3dbydscQDZh8jt
ka3r/Ecbmu/uJRdDKTxB+F1D1wVHpCOjbl1gI7l1SYMkzwEXfqro5YRb9OG+yZI/
OxqRQ7yAhKIiGFqffErusINTdZGCm2uxFKh3etCuAP4rwFDNHbP8r/FnHoZpUIfi
FVo7BnZXSHCmu2CPYF/LzNBHa4qMGJKWGSqFJfbyxCf87nTEZGTyIFKmTXqapvHC
t4D80HAXc2rcm2XxYYgIvzy6dlYA5X8dR0Mj7qqQ+xfBAkPMbbr4+Spbw2rOk3Zu
bqd1ZD3J+uhMFKeidq+XkQ==
//pragma protect end_data_block
//pragma protect digest_block
xvmqFP7sydJfXQJQD638zdNJuOk=
//pragma protect end_digest_block
//pragma protect end_protected
  

`endif // GUARD_SVT_AHB_SYSTEM_MONITOR_COMMON_SV
