
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
d5sH8sYk4XWXnOfr8pfzFwkmwjx6EZbMqQ6H5ITARg2SMJTo+Wgfxvn2bW2R6drG
dcSmWnY1iQ1ojXjf24Pm5oWdAbX7s8HFrPHufgITNcz74fR8eulAX4vfAGSxX637
MJvPy3KVud7dU02H5JiEU1hgXAKgrIo8tX4B43LZhPA=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 549       )
iT7OLxzt5iCCaKYJsw96fSeMV5l27EGpKfYpOmeAn+nvFOTGVaF9RKaCgCwzaluW
eGOG2J/QVn9EBbAUgEZjWM2WwFRnPRQpIMKQgObykS534nUA5iH70Uf4NYDkFfKb
n9nXRVjj0erKMBE7tRMVsW3av95MVoe9d/Xb4TMQiHX2LiZahPdAL9+hZzpyP1u3
m4TPGUb2M9d7Pw56bYRpA4rxgNQj+P99Dyuz9c3X6U3wGb5f/sxGLE9oVqfRnbm2
l+NjGwuFeuumWIH+LLE65A9ApNiquW5w9kvS28S+fuWK85VtPH5j4XNVF4hiUMBt
DcMyNamYhBBZv9fKwzA1V/LvR1ORcLBBbxwda5Cif6unRk51clhICKaUWAMDcXSz
05Vs+rx4ZkSZpTsnnaNp0byB6gJqFITJb+O0Mvo/UFU7uiCNM/7BALB3uoJ6532L
BrX9nxSZNPBYgd+eRNJ+mP4C7shzmNxpL6/vrCBFyvrDTyLkgHLadV/esvnY6sZ0
VsA/gUA1y0x8wlYhQ8vW2QnO0ZV3k9cFcIDIgreEd8097WShfqNe8Zmea85S5P9C
ZDls1wpZWe//u9F55xePeY9p//wvdxItQ1T8wr1fGYdMqs/58BKhUv5jIWE9Bw39
5gb5Q2MA5TXMxO1Jpg+SASd0r/EDTi/0vW33bILj2vK5Hy1009R1l9Rqr5CehVxC
0tFh+k1iU6FROVPGGWs0jI69JjZcGyM3w9Q4ttApQAg=
`pragma protect end_protected
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
C+1jme7yeIgqU8ABLET8R8BD/1sZdYznENE7myg3F8mg291Rv019JabRzNIl0/Pi
kJTh/eEr7euAujqVvLPM6qYDfotnBBdpGRhWawLbLAw4gF+nRn9cAYH8ABAxEJzX
a25Ced19X/Q3KPgWjvsN2Wnf+bZqrGlGfynhSHRtBX4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 789       )
TNqipC8RopnYstDc05cnWuGCcRkpeXmccpMzV47seednltQ3yWCbvrvGgadCyJff
zr3QMZXDaSwMC/3DAv7SFWIjOMrAoFg1xf25nDIxhM12l8sILeIPiir2ew//xS+B
srMmdfoM4b2KklUQk2XvQJlWkwYSfRJa60iKONFDOw5xAEjE8h9lKkS/7UjA4OnQ
yQaciC+K06vvvaqMpCOS+Y8MdS0LTBMQFN34y9AqxeneN2kX9EEqG8hxAJjNrzZi
L+HqKkObXIug9aHNRRSFOjNE6essyZcGwg2uTr8zxI7iJBBhl0p/BujPXFMLwd2M
e036rUHMdWFhMS82iUs0PA==
`pragma protect end_protected

endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KRBas3uB8rS3Sb2cWc4in47VD9Wq3TSZjCw4FfMopj8UIMzdJdiBkwFZ0A6tQRGz
zO5btCGiKnaDdL6zdtxojgsJ768Lrm4l5l785f5I9EV9kIDyCrxsqf0J2olcnrig
DkfwPfbfwieygomeH4tYhRBUSo/cEUacMp7C5jEIenk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1256      )
rj/9ba/FNnI6S7EV4Lsb0ct7MG3HTY7kbULTseLiVh234J6+qEj89jXBUn5CImBm
XIF25fdA4+AWscvmrGPFyXPD2zkK6EiBlrow3C/yeK5UXAE5SknPbLtLrKKf1dlp
kMw/3ElPI8lSI+RrMgArbnSGV4RHJwjpT3OrMTO/vAuzEL5uNicq7Oo1rwV4gNhq
MbzrdkGw7KG4RNe+WOylumfPQeFHlizBOAdP5jSxVt71y+CvWQfqoY4tS3MtwRxB
nle9osR3hWuuGwnUZUJVlcpbUTowNlYX365Z/eaAq12eivp7N30nCwFU7ne74p2S
ht0X6qFzsjK3DQ46TdSbl0v6J1Jjp5/4aGVrjkyih5oM9Poe4erF+nAb/2+wj/p+
FpgH0qOo7z6hq4CWM3UEuiEFs/LOdqdpsf2jz2MSJfh9HoubJ7EC8zsO31iyLJfI
zDQ8rh8yDVUUsxR3FQoHTPTkdVtlQsLhyAxeJldzZ9HYB/xzV2CJC56TKPJfbeME
+EWSbx28+GxIK4danRe+lyvXS9aVEOrL0oHBTvyZneu9KdWGj3YIYIvMhV/jgNI+
moHN4Ep/sfnLOohapl4rPVJCFmiAAOAhxdT+UFHSSwUi13rLY765t8icR0HsXvTM
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FqDsfK6r52mKcmqwUVY7u2Z8KVixSiseSkX8oiBI0H5H8bQ0Vgr1gQnraQeTT49k
uKUXDSqxDgqqhhsD2Vb4RIvkjy5M5cJrQN2knA4MDRn5LCurW8AQZFPbiyTb9OjF
2ONicYN+M6f9t06eN9weFwjL6971u4e9TD8kRGox9xw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 25280     )
zXdSfsxDEbvd/XDSPImWNeqGiEO80y6l5BJVj+5d+GRckrGRa03/gOzJd3Dgxtdc
1PC+kYLeIeOB3u/JmbKbpbjOp2MGtjM9EeSfszc1Xe+wGtCVJ4qjIXEzuedc7Ws8
2iNZkAoJy3mRTs7gjJ2y4QWTglOSoWTDvzlGPdXpdd9mUL4nC5k63BzqKyFDpcvZ
8K1MOD6MlHdj62a2n1ByPYpwIrceuKEOvTqkJIQJL+KbNIad6Cxnd2GTf+v3zL+c
NKknPkJZj2kykNo0bPbY4RIk7VGqi7r97p6p0+UJVJLo8qPrsWGbw9L7LWi+7XC7
bf2qk/KgvMeR6G+JfFEnZTDeyM1Kz1HyPdDdQq5WNJAWt46RUon3mfe86Qt1bVAl
KJmInkALXdoUgyfYEAcEd9vEsA3tb83lKhuGyQDtts3F5aQN+BrOzafxZhYkdTql
B5iaRP7IORBG04iXLvrRJ7LBFZeDi/uSi65mUNHQIYaGbrTMk3AsNAx/f+CIdtds
TLjsjFPDjYdbd2I67+TpxIU/L7K0SCcxV6+Wbf9AbEYWEHyeFwsyfbSn2gppt9ta
fSqhCusp9SxEhTedBLDNPFW45UM1ED/psxK9jjXCwPg/KfQA/WDIreG/RuWQ6bnP
g/Gd2hv78oX0cVCGlJBK3eHyKi4v5jKGtEObQgB6ihUHshAoXIsr4wtU3CItsgw0
te1GkxnRJ38hU6YFEj9yNKUBDDuHN4wbIMTfwMUEcImxsi2ghQ0gc/hpynw3srjV
COovZEgGFm5L4apX5oAEGx2hY/fbWuaS9ZqfYr0BjMlhNfADrfhfjGWgxJpfOUS0
HphJ3suGfpWRgjSnNag6iH0eKScXHhMLQYzvBrLGwoWQ996346H89wGSiqsjwrfy
fRENTt3hfAgeMjjVnpBKiiPrDFd8ptK3mYQlldSkso3XBy62WB1Kr5xkruLlMEWr
SBjnK+sTkUzt/pVxtJ4f6+knJAXd/WW6S3vbSyRysxd3MsZBPa9068DlsaBM2C5+
4gQB8WNKXgIUCpKXjTMg4wOP7utW/zFtsFJIOTTlktJcdGaB8d/Ia3NjOiOXgwO5
5rRxmWoRz15ecQbGgIps+hXXnYtRw05DlajGukcGt31TWdYzK/6GukJD5XRMl1ce
OI5tYkjh2usd69iFIWKUrkiTWlL6qqSdcRh9mYjdkPQIyH7K1UIHcHC6c9bl/Ceb
s7hNNcBXKv2U0CCTX6gOecILfi8DVhSUKpQItXsc4h3mu8lFwCDhKW1iIGBYW1uf
EanCMnzIs8nto8iL2KjqffRBugj0RJJQKDppanMrOg8U516gCs4kS668nrWKMTJQ
/0ouIdcRn1BdDKBxUksGb/rmJ3WVxQJrOG7raqC0ttM139ALJ1Jojx0CTZEyWVYg
KcTMTfIdXNAi/fD1wNyxFwlC96yuyW8dX7iWoyAFZOgOHRuQ3+AkGaSl/OI2niO4
hhApf74YrAIZfYhMypPQI+1EAf6tBq/Xlmav1oH5qriXh1M9BpfWKk2s6uaAI+DX
kSW6kfz0YNFCPIppeJADI9an2s3L0NX1RG8E1DzhTRX828h61QerFPZmvQytnK4D
1pnjhkVWTTUmwSVX19gnmrbI39WRg+9klM4mK+HbYTAWcukoIw2p3bTBDAUNSg4s
0YlNOs0nomaqQaecJBCYiVFCwh9IIvN8uVgqmtHJWUK4+Ds08bpDxcisTCHBNGEt
SQRcE2EeFxS13MLq3WSbvl+FNmg3Tpd3f528YUFKdO2y42XuiePXHrBr/v++lT4h
+57v9mrabLZ1SOgzyalbNRBXyJ+3p2Lx1g9gEAAaqw7ko6CZUz8AFR4LKbZcgPNC
iLB6fklA8g7rx+DIctTLlPMPUO8s0mpg0KWqDgkrQnLjCXAX9oND6QDdTIRk2Ni2
HNE0W4QL0AH+3R575byup8PRLuTBrbu+Ke5V2JFdr89Fz2gjxdCybjptvNIsi0Sw
vxHSFPZfsPR544S8ZuFptKPzWdmyD0jEPZ79HgfiAi5oGBbyNtJaZCfk/UTYmYS4
iCohw8xicTOr0v5XR5wjEqaqdKkU+niS2UioACfLUfNaYK+xCJuwR/Qy+mFSHFCO
LsYXXKMoWKvjuCenkOV3189Xgi8wAxhn0WNtDIR50FgVZKIcILJWvwIKz2A5x666
LQJdOILTKXtK4HnReJxQmM5lyQpWrczeWVo00GbJ9Vv9+6BE8ca7nDHRA2lKfY1w
88hl9XlEInPRjJ86OD74Oil95IFSXJwuwUA/XZvPAfgH0WAIVz7+NrDiLK/lg7Xn
7tLrY7EDkiaPu5QJLo94ZXZjG4HhGGHtwGZ9Du1P4DV87Vsa3SABZEf5KLBn87FB
LrfAOe9DET+kJO5/XOG/S5Lx9bTkqJf6/KfGQbqxhs0nns/atnGRBVqkbNMqTYhl
zAma1L5vEG+R34EMCDNJF3apRgQljLoJjfYI3rxlPuRFJZ10d/nU/0cOXmje2HEc
fSAAj7lneyd9XHabHu20Lqqjo+6hcm8FKsbBcvQ1iAFuqiWSRY6f82y/Cr2bKDrV
MNXJ1YyoTjHq19rFHmrwQdDnIyP80OtG3CuF9NL843rR8wS4hsGEhq5Vm+gK5uIe
o5Lb7STFhzmmD8iiT4CH37j1T5q+2HIew3jLC/cOPl1mnFphNMiUi5gyd31t/gfs
+jmXuy0buRXxlqobR/KVe2VBS47fEPCp2ATsbgii65lGvTNEqNw+5TOvuSkTYjyX
R3IwcPPCeX9Q99sVr/CVJaUpJAM1KqQ589P9YyQAFkpUBdABQqr0NcZy+PfiFap+
o5tuqCt45pKO2P4fzgOnmeY14CEplbJAhukMccoN2niWnllauH6qJo5iqtLKdE/H
4iGMlnrNI+iQfXrTSGfXASMEAhdX1l44nmCaS0FqbUtut5JyFTeWw2XQXi1wVaSQ
1/4NqX/S965YKBduzX0PrBs0bk1JwekZYTAcBv7BqA0h/XYNAM4j9Cyeb3Umyb0P
3+unHMeVlwdCASkt9DTSHL56sP43Z2FD8ftM44WbebCMJxwTaIRNPVUw+pokJ/bh
LFLQA7XCg1TEgnFmfoDcecMCKv5DvxaRpGW4tOEnWsLE5p8qy+S3DP2Srtd0QUS3
oHDzGvs1QTx3thVVIY1Oy9oUUi41Wv3gpNMOxVe8gbSVAUu1K3IMquKMVYWBxXde
yskcMAzveWZK/PtjjCp6XwiMGoXpmUh2kwsenBJFkmlb0UeUxuh7h8ydtc1Oq4py
k2zL3eCTc81lOxxsaTwCubGsc1VNi5Nprsb1ps8Aw8wtkohedPf2tKX9k37uvzcl
RFwqgHnY5M0X5vyNYigkBMFz9sbX6jjzhK+gcbLs0ZHfZ2Ksbxd13G7aRKrbaywn
E9hAO6S80rC9x0/YZkEUQfM87rs/IIZ6IbluzAacUOuA8RE8K2wpczYFjb4cXS+g
Om97SyGuDNRh3Nmkx3MVvO4+bULfO6041vkk4K93WHxhfT00XIac5f3BI0jfxa3L
Ca1QU52sTaRbxvtDu3MFeke5PlUluyf/T2DPGxQ5rc1VZYP4vZvHhEoel8foKMi2
+orBPk/NyWCwCardzry1KtvJp2TGhQCa1FSKDvj/xedUNAKOq55SGtI5JDiOEAPc
ygBUKCcxya4qy/YXqNJNG4VBGpIjlmg2mfTZOVRe+9J8lp11M4BnPI/+goH2U53A
UWu0vupnuoDAmLpkWba9QGS0MhOPTvJJeTYzCA9DfHQP0Dg/ERQrVX6l+X43jMZI
uUf5Fq6U+bzKmPmTKDRmfKUSEpDHk3RSvdZezkPQmVPnQcnOihqhuOrXdncl6m9q
TapqIgnWVqJfwzyuKPXdwu+TGe+BB+KiHK+52QXVduFHt6jaaYZyffgPBVy6vrY4
ABL7QZT/w1qEtIbODgoAivomMsiFF8gkND7NklYaCmKLSTPpBgCYSfbGnZWhd54B
ep2Nnbd7F62r0M8x3hfme75HAB5wsrvcIdh/ikE7e0B+syIn0w6MhqQKV+91UEtU
ff5OX0cBApkHb3Z3rFKY/HalXObj0dxD4QS8tP5zfV6Kql1MSzeNiQAMHtTWHisW
uiw0b/Nk/zPeoSRWmeznC8fFoKeJSkVlyZFQnAYkmULqqaYmOTgKRHYAk7tCYWzY
qLDoRqBoH1xn4kGmd90eivLNPYFHzWKPgGqh6H8kQmXuY2QVOsH/uCk4Rl8f0hXg
r9n9tIrtxFb3ge4UsQwnB0dH8aOOg+4A/p8gWfp++j0V94h4l2euRcjyijgKYqNA
GFZ3k2SSHJGMIgvV8Xy5xZhS9nJPte07rC/BRBN0v2KGdK/fumMNjOhYctaVNhEr
Lf63kxAcsCceKAfuLR6jKeCsQS2Zz2lVMSsDjR0qBQJIw99tmCXLN+TVvni08Soa
5BkqMjXS+oS84YfKK/CM4NZ7DQKphGRTl98i/zrNubc35OHSEQ8s8ZN/15ouHJUJ
kU/sGMd+lXubGIRSi5utrHhVkoFdK6vIxadGb7/gQ5+GYam1a/ay0rVf8mQ03E4b
Ku/pTYmxDN83O3CzmSZvjOvqUxquRQTq+NU3UX2YAOcAutI5iMwaHefrSTm/W0V7
TP2R/MGr8U3lzsq+NI4aGizkdlFRVdredlDKQRyHi4vm5Ee9AnIWNHxcqM48M6M3
xnObTA8YKtAbOIjZNTWUgunHsUVsU4c5hV7OUr4btc/m4FaHvHsgnV+q+doNHVs5
h4DdXvI27pA+eWBWUCij16zja86+HKVVF37VJq41UMa4fdXUtutb/H+7//1K7/Hs
xg/640JGRQa9RQFloJUJAFnDHcUKEWcAMLMKUmpt9CfunTieUFqVJAXHKpjsDnSL
VQsJPBAwzghQTOaVBxxTK0K/NQzoIxkMFnUlheVcXY0xehtkV/CZ9tWGxLWoabLR
1ZaUKhBcpIvIDU8uiFpY58L7Jmn4yigjcBdVr5t70yeosV1q2mYDmGWQkMF/txDF
t+GDNQAC9Q2pXltDgymFH9LIoQpDXBR5ExZROEYT93hLet2pgKFDEtrvQgy3Ev8K
REGEost1UhfvObcZ+oMU89ItrQ5n4D1v1YvKLh2msMwxF8B3KFHzQ5bSnU27QdLY
BQ+0gH/hscIHw6Z4P28b562LdgZo/ew8VrgvmQ8956H/yaj5PNrGUsr9mTbLcib3
YGd52Bpyw5Ey/+B9Rf4UzFfOerUVLViH3EcLDyl80dRddR2DV8fm0jTQWvDSTnB/
DY1+onqzbac6DeXpn47fJ9zVQJpuXi5nTMO4rBkdARSE9aW1Fj60PWNcFaOWTsno
uV+T1wCS4MU4yAbIg5zm59/55E0dm3QPV72e8p7wU8T6WQacsLNxunz7JMeLRELQ
M/QK3IXQgouOTT95Uv79P4o9BvpwQt3Gvsto4QjSren8sp3xqg9jQOnWNgZa/NXs
NUz4h0xlwhetsQWPzTRkxggrD3YAJnha2KnEkO8TfedGGsB2/FDjgNiDBWxPUHrs
QBa81bS0rrJvWACxsyUAyn/BtXGB+eVf3zm869JP+U3/CoQ6ZiBMUBmITRV2Yxj6
IDBpX4etdstoff9QkKNWr26jcGkYgWBPEjtqE06mw65KZRc9Dv3XpBh1sxRURK0L
v0XH0YILNhjvHDSKi81Mo3BnMnx37Y95XNlEbX27808ZtYrxgwEkP91P920VikfO
BbfDxBp1g7W4m9Hlw6s46G1z7clVkMWbFZPIIWKkhbeK1+gQdspvgCHZbN+9HIyr
iJpeK8X5E6JMwDmokrsdnnD3KIjo27XlAt03TwhFgeBEYbYVmWHccnjuNcrkMNA9
jMBIh4qSKFdAyVhxuk28PbdGD3dRer754kh8MNhijIG2TsfANrZMKitIebYH0sc5
W8nWJ0EXqvQeBDXOU/kQM/gYQNBrldkNIDeczLNi1oQ3G4CegjeyijQl7emjnVWy
ZubNNFkcO19xvY8qQjzuVl5egiSSZuGMG3fdm6rT5qj1MNWXsjZz7Ev+IvXbOyvw
moLHquMOiVjkUItf62HSkMe1oadxSoJpZEBXWPNsZ1E/qBzvaw8bmLWzwE/s/4Ip
kbPCxxQw5Mxng1SGO429E6MowKe5BpWGzEAbyU3kPiM7C+va20HBGJyWeKgLzcqv
uxdZR46UKl/zlNSkLUO3J5LSuql+67hD+PNGVBH53tPMiI/XvWrMDKP3l75Fois/
+o0iqW2mu/eP4HwA/oZQyOlh9OfC30OrTmVYWHZMKFpIEytWnyhsXyf0krxX3SdU
2zN1LlaOFEl2vE9h2+nGcN6JJAiGMRHH+jq7td2q8ajwcc3hdL0Lm6I8D3wcqJDK
Rotm7HNbZcBx4M1Oqs47ZlDb7kGC/Mr8zGshv0hVP7HUadvysi92HUqymljsmiG7
TJPefAzgFiSMHDkUNLpE6msi47MDMAiuJperOc6vx3aM3LU+ZQTeAMVGfPoFRVbU
SjD7xlXUOF6gWmXub4ACaEb2yuj2dg5oM6O9ot0esu+M3xW+m+doh16YOcUIBpJ0
sNwTaa0+QQB9oGmz66b8LO6Pmx5L96j2ZBFMuu7Vz1H7yyqF+pCkth0UB+RQ89Bq
zVViuKgwuW7BRe8s+I4y8sF6ZIUBUnrdnZgI7cKWudVOmk3yIHhxBdxplS0PkqsL
O49zh4htXwDm977bsFUkgYTJMxe98WodtErm3fwx12FH8YJ8cTlRQ+7rZe9ghpbd
AtJfdnvDPE/HX2lGfDg1qpl1T/nkYpby7aRF2WBO5jLDZ2uKBhGdaj25Y/rL4BaZ
xWNQ+e+LB0i2/Zpmfj+RhGexYS1z2gFti9Fa/fqAryNB0s8Ztez2nVNcjn8y1eNu
Rz7ubcFhqpuSPeKOLcsAiAEoWIosZuMN1fYRfbi7iWtt+B1UXbiPwUzHPESKnz0+
jUxn8/qmBpIAMSAhhYtN+LDugmdIT2MAPuRb8rn5DG9BGpqy5jQklYjmsWu4Euyr
ugfH/reAAGMP/GNlmmevfpG1r4AvVDWg8ZBG2qUecDVyWNxUzRZwde3OXUqhVLi/
hapBdDE5vYeB48tAnrcRq+DZrQp0W+bHn5mUp5DHMEJcmypWGDY2L+OtnziVE1l0
07qhFpo4+L69E86H5c20vybgeLUstBFyuNQLkHjOFTwLfVr1ouF8LHkD8IVZ6OWf
C3fZdzmuhBcaaKHkXtCOSnln0E/HuvKjQIqsg3CNDBY6a5tnt3gUKaFqi/A+i0z3
TQxPWL5AZRqZYL380TOxPlXbdW1YgaDpE1nIWjT8giMyN9iJGt7SDVL4VsA+LhXN
MMUzoOcu/MxQEL5hYesQYyZjQ5Fqz9D4KZa37q7hALZXj7yWpJeT4Ffddh5L67pa
SAYSGSOAOnwYVWyq49pHcna1TVzu7OQN0xkiCa9BY+zvCL0l8auebSgNLAPoU5cY
MlmCT/UH9ERyeiRDToohZFuwnmSv4azzDpaq5VTduXGEK60IEmVCE4qfruZh/Imy
wCOLdCnQI7ubcWocFXYBkXt9rnDCZrnr3MW5Ofpg8froH4cu6gU58W5/TvF8sW7D
L0V8MJS0TOWkFTKTPvdLjd98P3TVLBFkPQIuM7xzubvCk1rkFG5XbuW/t49Hk7fw
dbBcleeXchTmlrmmX0/PYES8s7eU68sELLrcIJ9tooKz/+MeRlGVxxPTIdxe4w5b
Ez1zq4hKyvIGxAMPAvspKVXvP6g2s7gRXvXj+ikj1wuMDiIUGt+iTpJWamWfROES
3kW2tNqE5QHSToCiSteAuwIs+0RwAa30CsfaSHwpD+M5WU0kE482ENLmaoiFc1Eg
otnaBgHcCV+qS5dDPh5SKf+K8rktApEF07JnNItBI7wrBdagJo22jZkVtVr3u2KI
vVp2aEGA8/mINdeXhwRaAmiUbusSWGmjb0W8X/C5aH0AiNzkICba4X3LN0p9K3h8
A1KqHTPsrRqzRa2XuWEe7++9cGIxdn3elM9rkwp4bVPUR8yPjof8sGiL7Y4iXXYd
wnPoBIcx0TFbbExcirwZdK2wGCkKHCwDBWgftGtM90mjRK3hF66uIEejM1Nrak0d
YHex7Jy/xuocow+mmPZr8jmCjnIZJbPmyXb6ldu8IYaBYwtIn23lp3WhSxI+NUxq
GI9l6egIREaA0iEXIYKKvj4hbGoEDFEDH2+GG9dzwBABrVXDGCdI+VXEBa71JceR
nCXr7WDK9zwqxURSpfg+f6jrehzzAaSQVnYmj6zBA3cLfvQhZshd8y1tTxAhxktM
N/47qpDzxlZ2P/CitfFG2F2s75XIqErD4z3/u6hzsxgk9/W8N9/uVqDxAGJtAGc7
l4JAtPwKxoF3tOFsMFYWDs6Gq0pvCfZbh2bamHPgOMx2mSMX26aUuzXmADdajF0I
QR9JEY/Wq4vv/dSz09Fw8lgvCNUl7KgmKr5g7pkAkC5CEJa0U1eaUMXIpywteUUv
LiopZOEcx8oAuCa7LdZvcmcwPBGH3lILeWc4AlMrBE5sqFufaoVXFVGOri0IcAKA
/F/ITVdYTVntxKWqRAdrhG9vGsBH4VRo888Q8Y+u6iIzwz8qPyK/yO/tIifHIKsZ
sAhqkvXRPdSWZIxaaPiI6Itzy3/sWD0n3/lv/ZqGL3+aTu4NaXelyghS5eJYxyQy
cM32d2yUcuA2qqmL3Q6hmvUSNsbzcUxfJ17MBVUCxczc1qNJM0BwJu2T09/QfbMy
4Js0CToQjVhOaN0O0J/tgdFoT/IRh1aQgTQsUeeiTT4y2HB8jgxX8q/Qhvh5Muty
PnboKVOb/ehmgzPGtHOwaN6lcjJ0pCvNsLzH7NJJZxgsPz/4HgkkofqHGC/t6Ej1
Zc+QGtcw0VDTFBgoipplZbEi64wWLwvRPcmaUWglcR4KUYAFxmkLgooMFyjb0tKx
wcbijg/CTRvzVwjAdqY4er0dL9CET0T1Fla3luTMoeXYgkxMhtKsJhnXR5j/fbZT
5J2wxqS8t4iNiqQT47144mBB7kOPfV6vbPMzY11oEg7E3m4o4pdpaqA3R8YHCxli
IjZhR3IHS9U35yWMiZx7azQR9jfmZhW0viMiaCtBPoaZqXoBvhxzpUw/PcerArQB
iIs6rqWqwY3BGoZ0dSoaV6N2WcUCgP08wFt9x4xL+CMdG1UwQ1C9qD3X4FMd19zY
c6RL7w4J3djIG+9vn51YxvyZyn7KJOPtH8P6q5tNzA0/eUp/0g9RVquTEGO6xW/y
cZpzGaW6pKqY8bk3SO7+LD7/lxeCGktlTcdddHUWMTxyihc1o6sk4PoHo7MeXpGO
xghE93fK+4j9swgPNiHE9X6vPeFBTRiDrJyp7Yw3gyRlDrpGFo/0M7Z6x6qUpNgy
I/DjipJmg5VEJJx4vuj0X0et/VuhQ5woThVbikKAo4XvSktgIOApnab8C2teDPN8
eTZOm5qObYtZfe7trbito953iYEUz1IMzcZhkX3qWVA5NfRM9IL7ITpJVxu0vxo3
hEvxnk1KcpGlQkCD6FOBdNfDCJONMwfLvbGIQ8JohhcWlBYVeE5UO01IW+yZZ7n0
3idGJewlbvshJRUen5BiT12sDvWu0rKT/2+Hy4D2X+cD4inc2qbK4G3Us4FElkLg
RToRtc/XxpMvltWF9OcvH3JPKQJCnd98A1IJ4vFZgrFT4K/upLAPZPAJlQnpe2jR
rB0vuaUEANME2SLy4GaEb5AAj7lyOuhpby8cWko4DyzfThKaq+HYcEoCZZ7fQc0y
Wc1KEe/mIfaZM5k+5Sj66Ss95W9/tgq813HmrajttbjmMKgQLRG2y9qAl+qZEaPF
BHf7xc0Udgzw/LUpJi4OxPnORAKAryC/U9JNic5+VAvGrbkijjLp9noC5NHEN9wE
FtybaDc/rTlmpOzgPCk3an9wZPdnJNSkUJMh9yEwvJGkkn6ftbRt7i/GiKn2Dzza
uApi64c5UTF8mW9PPxJYJHEJpXCm370o5x2PGb2yLkER1bZeJknSwCrRr9Fe9uOe
g7/b2WNZsnpl0GrjqWDNq25QJFlS4UaZM21um/757NAG85lnSEbh4bsbfZH6O5ru
Bsgxv25aAf8H/7uFSvl+Ex9VsSnbRzFVXessIl8X8UewpKheQMleiU2lo56u6ftk
TkVj2xW2oa2RFcgRm18xo6lx6FJhV45M6IjW1Y/Ytpz4H+trmZIbSGFNpa7NaVNz
wEmuLWYRqE2faYWw9O1Vjxfjkkx21JsLv2bspBFCZfNBed21ksC/sAwoeCCfJ4at
iuW8v1GRLC/Pjz4lfUr9obIdnhvAdp+A0oJUAMCjyuri4ha99lQO/T+wIDDR3l5I
W5AWIa6PXdXL3oWxLXxkztQ45A6Tsng9L4jnBg9KdvrZnywUPYQagmtU7rZejm9M
l8yfXFVIYAf6ZtsoSGGGGUE4hwaRBqBeNe7pHD+QNNf0OqDpV1Hp9Nlbu6Ve01ia
uOWTzzowAt+BduXta0mUSIYyKf23QapBkiOoLUIwvnudmKgsHXwdRebCf4nBLqAJ
9rtrinkTvbPb7wc3Mas1S5lqBypSUy4rQtev3EZD1e/J3p/cC8NgZOL5/XENDsDC
Osh1yLJ0Wf7lnEHY1IWufyA1nhoC+RqIyPnSerdmRtCBZ3KoQig0glExQfwFkblW
F0HpBfj/94WoPrjDdVWZS6TnSe0YRZWD3rzuw46rbBHds1zUQ70lbl8e4Jt1AY2b
e7s7C8ulPiBJkCEg3w6j08GjECKMQvdFNggaAw31VLtbKcjhDy8UnhZqXjWGMQl5
IgHO5b59dmkD5+zQyo/gJnOkhP50N5PGYkTDsvAXHl2Vj0eFuz8ezgb9tAGW6mCp
+YyzdOgxU64WJVLi0m6A41TyiWT/+OI15VUofmjyJ3f//B1JqTB6ccEDVVUA/iD3
i8pY1WqccLUxXZ9ACMbieLcWLbhLZ1MeEdDnR3b9oUubf4/QJuIz4/wOuIQwBfZf
GXbeLSdX+bsbuR1X+N4igpxvjceelXOJJim5TnkFOtXMT6/Zevy5sEnnUMrpfvR4
Wu7TcJ+vJJWp4knVT/qKxEDPW+HDqVj/4mHFjboi/Ghuvf+kfEf2AVlZJyF6i6b8
fkyP3FrvjmjlzhAfxwE6HDXcrVP+ERMRkTAke8h35g8sNfFQCUrFpb8LSHZeg/4s
xX9U6x4HYuJL69HdKxRZHdU7mdZM1PqZuN2Cu2zk3XTx2KZImbZGodMg7zFtXfDB
iNSbaUVZ5ZS0zJX7atsIpWCj+dvHFO+NqP+jbLbaAg6a2xL+qJzyK97N+pQGGlZy
T8+z0/YqJJ6z64aJ5WJozszmjs8nWqG3WoGnaingsW8cDJnW2P0cxrDnMrCVF1/n
cgd1/VwNwOdyzCjIKzt9DjO3TU4A/5GN50gm38ZRPi9a9Mn8py3kf6eqm9d2zOJp
FPRDnU3iaBJ8MPhGIQczZdjQOFK0kk7fhNoFYbWzUBRnPJem1nV3hDnkeNRv4hEx
OFZGdZMFBlrXSNaiD9CZ3HKY5TKbvjfs8OnKCH19yq+oIgpQpMNtysPj9JuBIGeJ
KivDRPH4fxPjhrw9aiWNzQbP2gAIrM5OCv9/eQDzF+5MW0IF+f6OaRXwwDfMHWYW
v8dzB2+XnbSw54iibEh9BtL5s11Xlz2Q1tBOKXulGpxEDBKwutFAJNKJt7hSZVC7
EhkXv5241dCVz1+B265z1M9s9cg9ceryTs0jYNfO/Z0p7gx9zcpWLERQprg+Knef
CpcJ6KmNKc46ZhbKjnkmR/128bF8dml0hDHUZHBdG9pl4ErQ7IGbc+vUWvuaC6P0
nATXos04J5RkC07nEN84Is2x9RwPfT8RRIgcvWCRlXUZVMZhMUY5CAy+RZYxtztr
6/CFCBF3bzuUjFnh2W0pLr66AInB/oabA1RFqMNn/vik1xJcEOKei2ggH7EoYnWg
QMv+q3J7Ge6MRmGYPBBXt2MryvulkHrGy3udPv/azclRFTaQ2xHPYjlPZSPr12Wi
Hgz3888h1gr4D8vRO3+wNeW2Qw4/DUWf7KIGiGtfEkimwkoOfzvNQxPVwTx+Va4+
C9cVfDK2Zy5YiqUsMEmBjH34wsesrokygmoLIhzP0QfRfzZ1e6oum2RYc3rmY6mp
ebpxDop7fwWFdci2uzaaNTO5XYmRfDwPAvUADd4E6DLyWMKCNqztvTrDqvmxqFzK
95cdDenrcwW46zO8xydyaBiuFsAEIW2jEVi8ZGfsbLC15fwZl2XpmkstT8lJz1S8
aiNF9dXMiZ2c3behYxeZ/ZMF/i+JCWMPbongxPobIxtGPuD7oeHyrhRNPT3MxIZv
WCHvCEv2FXZQbNfhLcu8ikFceeuvaXqwjAe+A0/EI9lopB53jcv57Gk6pbfeDh9u
GEf8bPABtOR0KsaBRH4z5FjSzbSEqdMA26q7nalFpGiVSEXa4K4DEYIT1C6qnYjW
1AxVh5RSmGvoSCNz0tccfGAI7IBFCN6LkD08/ucGBUuEIkilrlRVDblGKGbHlP0c
si8qZvHKfdQ3Q9rX8+c+ALigodKj8gdqLTIPyOJj3dnIYzvfCJqmkU/hR4Q4RZ11
mgg71jCzaN6qnForLRW1H9QeGQdU60FuUgyjXcSXcT40KWiYLU2OS4+54NAShf5L
Pk+u98lG2tOx6KSYcEXTt33+y5injKswbiq2VyVy8XRJ/Nx51pR617gr/lsvAmD0
Yz6yG+Vn1Aj576XRJBVVV/QW5/SiquSccxMB4bplPg4lM9WaDytPyTOyC779y9S0
tWKFZLjL/3IV/+kA1EuELDEjqr1PdXSNk01XBIH8Ihq6RDvT/dFLinp+cCTZiIkZ
u5JqtHPqlEaIf9teTRwEQKvKsENaMQ6P6uIKqoUCjEykvOGjWkSm5UZAm6MQrGIO
RCuqufTj40vdtfzQFBNTvHNUOL7LZgV2Ia0DDUtqCfrCMHvs53A60TZrIpguMTyq
J+2oWZpUdHV+C2u/me1GnRNUtVjZhBJSoNT2jrToMu2TfDVCjCr6XLbxJBUQQDZR
oShz5xAiG6j5NS1QtPShS5c86Q/fCeAMOjxuhp+roO+V+taam7XjTp0kzfWhFmq/
vVUq52o4ZUPjAwc+ChfKjrKgasDLaM0q+y9oB7Lm3mpB+XLiLhwutmK6hlpX+qWY
BDxtGKdfW+3m6eF/iAZuSHsERkIYc+nNKhMZZDXLOAlh4su8cvY7QC9PAQ0yggp4
ygiQVmlmFsmRCxYHaU9NPJ31ZU09zBLT52/qO5klxkr8BM8fYCucqTqFfMZ5fDCs
qdYtGySiyYCp83wCswG1xrTVf8m0Xp/ptcSwPArrpK9UrJsCMbT1HXmj0IAHypPR
VHTQj8IOjBQqLv/Iu5ySbfG7gX1hi6B173+g5FK7XlPpSJWZ5ZHBNv8I/1LAsdJ0
gyVOZnDsMtwitISbDi2CM62TvtIG+zKzSFDTs97LacwKuMU9AS1SYSAVYILRNcUR
+vIrpZAJOUxnWlVAdsuokvoY9xsoONCupxk0R8GfX9IzjAHkM3N7aarRuW95s6/x
tPpk9SEyw5TOQrP6E8/2/VmDB3XlPYl/CeBrdqbqxqIJHPPqimOBVk22ZrmNwe3u
5MN6VACCbu9Cn+l2PoW5S22wgJdAdL1n1VqIOpTSjYWTJHeo+SgP0vT1gCgQ0nks
kfMuyoXb0coqUOcSTb4Ijl/ULL8+o9JHA6A1O61GiOFpOMgoMbTuoDzuMmOU3GLS
+xwaRPE+br3slMk+pcUFiZ9rTQDhCx7E4oOOgAsZ5lNqmJ+zWKftW24oOWOBSVdh
uMXZolcyQQtcE/SPwwKtM7jTxs79MV2nI0FUAf+jUSyEdc1mwoRj+jfUFwyCiUZa
mHyIho8g3UfT+a4ZLHyc0IH9iUDo1HSR1/h/bFJfOMZarMnPOZ9OZ+ozI2AwLsb+
shTS+u/eyBImXB/TR87yg/V1ZEw0N9isUPVOYjblmVfUCRJ+k0RnRoJZjaQ1HbRu
AlfALz0EZPP1yAflHfqWghQVXJqtWXR2SrfQ8XhbW8x/ZTmExBZrO3iS6cxFBv4D
7X5ATyd36qLECFNwZPj7SFFKcySK2WrU2r04laihBQXZulFZlvlMdtFIlzDfDt3K
9Z6/94xLC9rlCS3F4rXNlPUO2sg8ZBP1U/+WVjD9y1QAbsGZdhFwJNyJ+bSobmFR
5UBXn9f4K/VZRCJNbTMATTtPWLkdAiU5C9XF3wJ2wdEdWohERwaRIwoGl+aF+HT0
Mmcd0i5J+tbpugbwBden9o8+qnWTrhB0Idioer9Xd/V9wXCDduHx1fzuvEK2EnOA
A33mLtRDXERM6JtNC/CVyQgiwll9oFq12AJ6g/M88ozo1q0aDw414jxJHy8NMTW4
+vrBpA0M4frtsI4VK0zltG6G8CHHeUcknmTnCE8yrTTmhsCy7k24EHxeDorGEJe9
UXa+8YHLgx/VpulCxGodC6bSkk1CvjSDyZhxfieA4vLpDqUUP5bQPQC7opktWPhe
6PoE5a+N6aaRlPgRpdAhgE+eIOn4gswXAcbUslWeCvCU2nUaJADDaaeEFqhQRH0C
KBnPJpPMyXsfXvjf3i4riiyHe0VuGb8InHACt2VbbQRpwEqtX9O951F2DFNvO6ht
wHs/aPO8C00mi1yMSCDkYujMgWD8cqEqc46v8iKouenFDMJxf4hbHTF403NWHizd
O4u7UaF8xpyXBEag4+H3gqa9rohioQjwgTuTkMVPMOqjTbqi2R4jB1EFXd+5C3qS
CCteE5DKczau903CF+eptWc6dnS8xVzFRi2Sb2l4uJWU3He0/+KHG66mUBuXoFo+
Nu/cPBDEzW0Gg5lKMl7wdl3GHh6UJrjA27pFEI37RuYFVRxJxejuRJ91cWfpvYDD
7z/5HeyQ5m4YkA1n89S2eXeKhSI2Xjd8AUlqi9T2KQ3hj9WzFcMhAitXCRFJElny
GaAXYz1ecfYLJYT6aKkFt+8O0wHKBvGpjy/kiTKfMIT6MbVN03FDwcgvzhF/jD9z
6zM81gaiXwSOr9EYZ6mDsalyum/EEOJbui9rCFUPpN0FLIyGCFds4FjZhTDJNIGR
IAbXWS0EOE+83nedZoiP6nUrwsm93yLD6ktk4UZC4Hu46Vdx09ERCC4vUIWplrDw
zIkbBZu+8J3lRfHQG0zxoQ1ObDJaP6HrBQkU/CDMF0zY5HD4t/fYaZ6y/i9P3n8l
ax5Gnox1k7ygmlVQP0uQWeuK5e3h9ht0OMorCEarN3LeKAERO5XGhFuEFJzztIkI
rC8XN49st35hDPYoF/WCh9AQtZdtw5xIu2KrsZKO98LmR50P9fYCGlzhAuDmnsVA
gbCShXgM60vpxuondJQgDJi7glRe2aArbyrGo6DeUQaIZ2wuv9h90a5LkIEuuvVl
kPmDQ+EhMN3+nvgYHPy2qEIB9OeKA+0sM4utZyDQaAexW849Jsf6Eqc9TMubkqiN
O7FRP2KC8I15a12qdGuejFfX5CCFXl0+zuaT3BR3rmkeHmzX4o6WdRgAOgIblzqz
weX/Azril+vcw0DjQAAXe5C3L1YMOCMzJ22iNv0YxThkH6+Tt98xrJHIjdTbM/pC
jRuuTYRufCnp8SMFQdkirsnkIH9qgPQpkLDVXXOe8jP7CjYPTwGdCAciqfYJ0rCk
eba+v/jHkalK4gMEDZNtYH7FFcLd8AGuQXrz2pMuQcPdA8sTnH4PNqU7zst3Vqzz
RzOFAvxYBBm4GCGP1CjAHVtdhMEELG3EDq9y0sWr35QHUT6AzpjVB7W293hspCgj
AtkFrZcuwp3Nf0DdgbSQUwUcKb051igp856rV1AxUMVUayKR8Kx4jXvgiHEY3dCE
b3+tRleY18H117ep5AezGIy2u6/37Pmno3Gg4fA72u7MwM9ODqDX2Ei0UWkuXbqm
ZSxwg/ZZkxp6dX2OdVgLarY64lslibAs6VnBDKkfxvbTSIXKsoFcSg14YVDkdFDy
GLRe1f1SVm8QH87atJfj9a0X63+PlwDvAdUhTuVJIE2zPBypU52VXESdU13T/thy
et9VB4RXyxD/aKNU87URwMZgeZM9r6iynEZX/HwrdhW+Yyohq0iD/vy6+J8jOOhV
gPEfwh1eFfa8+4aocIfCbYtonau4mGtO4BFO9l3P/tZN2xsm4X9IytucCs1s+KkF
A2gWC3mfLz6Uw2oP1QMd/d/hy9scq882ZooOLHXcpCvaOmKEdtEDV9FoGcnq30UQ
RXqoBr5SRIACXttD/Rf+ysjM8UJ/Tnt65fLpR2wU0pILtckKkyaWRi7Ou7ogUwNH
zKSswsyoeBgxKcegg2avaMI/DQyxiSrLB+PIqjLW+SgNMw1wKN7W2L3K5NF/C5If
ejyYW5AgWHcE61qN3tm9MSSdZ3+WFutm12WVSf9U+QbntJagmKvpF1+NS3k8yQS2
27W0Z/r1XPJZeT4ApKlcGot5tl/7pUPDgsNAcwvP3e2f1eOlNKxnMJqrnNwiCKjR
XPFfgIkAy6Jut5OiEJiuLOWW5q1RgVcaGujvxuHpDQh2ASu9Hskji7gH4cvGAAQs
BBsnb2vN1AWzp2zccLyz3TEtG4RQzxGVNo4MVsYeFlLSMlmtURa+noWdGedIbh2p
PRTQUv4OZg/Pj54gunBiSTkL3QIPqV15OQH3H91i3qPohuAe6bJBkE738ArfDZZ/
LkIIKYGpr/WYew/puLE2QlRY4idSJRasFmsNnFsNb1iTaAxE0NTmX8Ibre3W0ig6
y8IawPhwvG+SY1K4tSDTEtKJ+4GiBodd/g6HFlQbCuMyks+bp4en44OcWjNDVB0s
rbUnKCJYlVL9EyhYw9i37gxia+PbIWBQmy8bxWnz1F9+6im8Qw8SrfWiwTXnHtyp
0x6gtXG+KOYRKHs8I63NU+zz2kDEmC3BLiAPnRxg3Rg5QaULZmo84XYHq3Lf2CGQ
Tpg5sq3Q1QLA6z3Fmw6qtyUB4Ez89BX/DOnyEitqVeNwWUoWEkiAjjfKJQ+sVWF5
5auUJimUoLGVE1RQFO0GJGhRM9WJJ6xKy5qamSxryudOvfyb3JMpmfWWKttD4Gfi
CNcCX4LEclVg3N1NvDQx9r9oF8lVYsAbQD6ZNvjjvT3xC1nvomHJhjg/bU2MMNGZ
RfCuEz00WKp9zJ59qKmMdjJPgYOR6m+HbmoSzQwpw/iOv7Uh8UlDO3ecq2A1wEsM
bZc/ArDIs/ZcExQSuItqCo2EZYk+EVSMl8n9vHOw4TMUppYVDFm3uHJWsHzFyJq/
hdLdfVgsfY2iWOcUxMYPAFAVzlv4d8u5DvvrL8kixP3wov2mGY5L1Id+dD02RvvN
GDqsdFMFqO/LYKh+bf5yZafTIeq3PwJkJLy+4o41512UL3huJwWQ4ZsBubixNO9O
A8zjAgVLt4DnBWbhDlxnLQHGgBkMs4uNKCGgutU7G0pBYYtV0T10COdwpk+FrAW/
rzlUpd7A5Bt1vX9HRZaoceKOR/nkqitqdFav2Cmlhb8t96Dsl/CbgnMpAW90xer2
9Poc6jm77kQF+4tyIq9vKzaegpsJnHTDKaX84pLmBk969JoV5iBOdQXD+o7bw7lK
ajunQjo6zllSiHzcxCXUeBIi33BTHsB0nx1MOChgvmP936WTtf2mAvxPtI5RTBQG
x59ymdT1m37KLOk2JuyOKVKiN1p971WICQoQDNJLZYhqdgTqnkYwMEMAYfR5bqJ9
LSRechHUu6rjiKDC+DvyrdXCx0sFK80HzKmwEz4KdaXOxCb0nLfpHGJp9oa25tQq
+4OVP9vEyv/rWIRloXS/4advYaVB75xG4KU6iVPLw28jTLmaa5Oh06N6yXcR5O9S
p2h4pTDpmsyIcflbbXMreVm0JpQoczdayywg1oics4EF0p+5AIMN9rsIpIn+Rc1H
nIHNcvY/ZNk8RM6AQs8jPYE+D9BtpoW4hELFucpcGZfVYYV0Sr/vTtoIq0BuwLh3
2c7+Ac0aFajLcsFZ92RysUI3M7+rWczHxaCW4V1jYSbdln6N1KqxL1ySEjo1MG/Z
LgX8K43jCzYlORorE4QM2jnGj52+7ti42HkW5Dp/5XJYoVh/mf3aCzj0Y0OpTeqL
GJid74GAa9l5s3bncXRjO1aHZgi1MnbjbePfuEne+IqNH9QOJOICDRKXQ8TfcKqj
z6bHJldUXy+CfcI43ZidvVZMKoKMg0qx78GY5YPHw2l2LviKjXtXjY6X1aFZg3CG
ldQq6F5d6rv++A+rFvO+NZviHZLoMYS0Rcw1mQNXNmgnlgCNwo6ymGv5J1FXxsZQ
bh4dEN3+T6sFB1trouGuhmx5Ct/ua/o4tlbHn7uZTpboeV0zn4A/p5Bj7hlpaS8C
1W28QdBbgHg8jkExIAR1CCFHr2PgaeO/ZjTM321PEGYLqD39+2NseVOHCENxZxOl
cj10G0HAelXQ3mFsHz/XvyzAbJl1pEBkLBQU9EUMKVVi2i/goUGJ053vmoV3SI0X
WJ4uRVSWurRE91PFsoKolpIMcraEAnG5bfAXwhmeV7AXKec+RHTdSaumLlZ39bhF
sQecwXh0CZw2xQqhdFEB6knEQBECyKJp1UP9B5FixRc8R0+/dOOUNSWNEc+oSNFx
fBYBOkxJW0m6qk7j4tORrNyAGdVHgYY3W5CwnodyqDpMv9UWx/LzGnxXG/dAQjqv
l2nIvcqdz6WLphhEsv4k5m+/atxP9n+Giw4w5qo5JRH8FOLlIb11CVGkqix3S4Rm
vmJzvk3RvqCN+Z8O4j5zUOt3dWlFcvG83H0AdWTc4U/gl2Fke2/WySfzapZFK5Bh
Xgl5e75hPSBp2Z7sMyt/B7F+N1pxvO8UXNBw4rdp5rJUHrqn4EwLj8UvdEXmYtVV
sDUpDBsTwBkjN17Il3tep1gPtuTuF6QRXmQ8lBR9JGh9Ijllu/DNAWEThpXExvrj
3esGnmCqHKrUZRPzUqC7+ImpYAWAyHfjt7/IbUxWTTPP4SVyABppIK8fL9NGuZT2
asGK0c3RQ4EWqSc0p9BkFbdG6wKM3XeJrVFxHklQSCBIaVOglIlywHQcZYjFP896
RE6xY7bXWY4GDULYlwxYeWNXxGQSHlKfzp39V0ZNZr/+lHw5Xx7x9P8/Ue1drQsy
6OLPbgxedZ3FVjcq3Pmf+Ep8KPXZSCLcGNxP4nG7nm1wBnP5C+Z0MnBklE9NifUj
vyu+v+BJMIZEIlubpY3PHrVYvwEK4drCH3klmKS020J8xVwe9dj0dfrbptRrHGAp
fM/miRu748kvIwbLZpvlHrvbCwxtwRfliYruepLsykdTGWDkT8n3FwQ7PE9ZcLTE
t1CJ75bGJ+TkMrERasplZSK7WiaoKjz9tdG1/cKoqwGZ8rm+D0tRqMBQ8ryO9yal
vN0SkL18RnzjMyGOB4jnzAipGXcH7AvYIZzm/X0K52Nyg2WcqQWX44W40E16VB1T
/EhH1j9i9sF6DYU7LN0M2OpSs8U0llPZYeWpbgSSa/PnIcE+JDblmbz6GKDk/2A1
CQDXhaH8pUVZZtQPtW53PMKfZQwTR9uotNcRq1NwLNofUrk7KQJQncAGrCiZFZgn
dE68hvcoVsm//DzGvjKnhgKzIdmw7BT4Lz1lR2Wfk2BSs1J6nRvxNngLT2XYPgBh
pHVbxYEAXFaU7W9xvQXiEnAOWvzd2HfbjNGb6YRzQwKo4TJjefHUQeRijaUdfeYZ
oXMvo3R9dEOch7QXTs9uT9P5GQcq1oLgUBWLWenyy8RWbULTGMA9TniazJ0v3J7s
B+qlb6R7+Id//1JOKB8kme6u+LsJ1uIGD9oOWJKVilOigf+u1TpyP1bACtym50g+
yvvB3GV2dooBjdw4A+yyViKscy8Jksgo/pjaiZ6kLBuHY/GrlajcMiy53brDHjD0
IUww8w5xioCrEJ4X9+dyvvPJyZF1Ccu/hYblM+CD9Y+bdwHJ0ia+kzMLR+rxJoEe
sboD90KopwyjcxSxhJxXtCIXd6KiOHPJVGu+/LXsXSn/vIep3pWieM0Yeo1pmM+2
MQHBC8BMxIX5yWk4ZIAcpDwTDEasVqxtAekpYasJiwDDIGv1PHu5vU7+NTJAWMo4
ivwQAa0KGeFQ9qQ823flDRcKSvP3yDJ2NR9OUFm77kuAwFl64bpl9FQZoRZv2ssA
LjBvalxnMX9ZEzv0zw2xym2zpEsMfTDk3P3ZjI+8o2450WNyyc3R+T72CBnwUTXw
UUTyrj6H+eXmkEZTHanZj+eSF65Ktfp0RD10HPKDoDANlTrS44ktcafiEge34ozT
cg+qSfqnpxv6WOSpC+D45LXwLR81NumfU0J5GQY6ULWxaDHfD1I9iKSzK9BorCKw
pPtao9BnjlqvDygyFWAKg+Nt+WAo2y/B0aDekT/6Qogdi/8ToN2cBOswCbQdjSrS
+a5cDiMxZrk/eiNW3tdQg1ki+lBQOkGM7VegW/+tTLZn/Mtyrb62MYxNKj9Dfwgh
t+HFhyRG3ozSnMYgYZ/XoF+qXs1WkRcA80D1e7dBVWo9NezLi9dLT+lf8bRNK2pQ
vfyS/jQXxQbmjNSbj1R8Cq9XhPTtmYf4xHphFC6qzrxUARiK3i7uADeA3SoHbN0+
M28yZmrCYR5O7hRgaWuRJybMbpEg6WxHQFy5CoSHe72DVCzSDsLbEkK5gfzbuWNH
taBtL9SaaEMlBJF08RlGevmFS4dnOMWkEAqZVyDNwn/otU0lGR2zF9Nnb7WkaZB0
JzwRUqqU0KW+tls3lYQX9ixWa8NnwFZTpEPukYeGZUhTDiUy2auqhRi+hmLNh540
Z9KCsMx+CnfzLQveMknJbkt8Bp93UajMgcgJkZM9VAl1q2BRsfT7P8kXHDD9GfmO
rWxKCyvBNnafyuYVZhhQMirNmjbH1KG8LjvfVdCTCWHq6e5cIbZfWg7aZ/4S8K3m
0n46aS02SzeYQxMr+PqGwnblfouFgJSXMMIb8WUPKXvOIZJd4qG8I2UMH/3U0zvT
p+6dGqhEFZMGzFio8UPdRInTkFHttqDn/cB/kzD6DNAlP8ZUmkULaoCB3R9tivqD
W+gjOC09S+vfpn0Q69qMNW8DuriZMX4SneI8+CjVeLVbK8Hr0FAXaM91UCLJ5+u0
SYR0GbEP9vO/VxX6SbViMj4GVU18MNVR4drAr+LRmTzn8rW2WCz7DIXyl87Wd0/Q
HB5DXBjSsZ3vlj4eYv6KaWE+tzCl2kvq3/M9xX/DTfjHGoyzjWYVFlAE3+yY7vCo
1ye/VX8yQ03yDXBDM+PYgtl45FvG0+l8okG1ogdpUJMhH2M9ijScALIEMw0haZR9
JBCr5+dH9e0SY/9wGYdQ2LtkwmzeEihBidbzayB68Z/OKS1TvhQ6jy5CHb9dE7Ur
LPpoUoKleady+JIBL+Y0T4VHW11OwWPf+8XjfPDevBYqPz2u823eMpx71ZZ7cefp
55gqoyyHPfckqaPtQjrHG60K6eOGTifi/jUN5aYJi0zgSi3N/xOqCwXiQ1EfhhVy
0pOjbA/5G30lZDgsC4r2ejtMxFXbU33a6Q9DLm8ddmktcPipgzIb7I6nMxIXi3LV
5idOAjYC+FIwaVr/w+/paSAPqfkebEcBOoADg9xdyQsDfXeX25XkSmXJ6SNDK0p0
/8TurS5GmfJrCE36/N/mKqJRtq/YfCPmdFx8/hmEAEmo6/8KA8BJWkFSN5cIg7tJ
FRbLw4rIJaIRP+2ie3WvOSUp5TaukycbkIP39QKhD/5leSAGWu9h9gJhgfWRTQj7
rvkbuiSGJAdF4ZKbg+293vz5j55uaUppjIslNMt3N+VnuHjcEBCzVw7bOjC05S5l
NYSJydp76AXriXJ+RUyTLihb16nbVgwavA/Qzjm1U7BuOFSfAosG9+envApblg/V
RfE0ARb6hIU7C7o3VoLEpDQNFVokIwdTTyHvX44s6pIKC7zbDmEznqMoc2WXrFjf
QDUU/XR/laiuwdNGIAoKxef2ZeEpbXA5R791koC6YxiKgIsIzu0TiQ4PVaWOBSXM
yMyNwB8IdNKh+gOtzcOWVIYAohZxuoX+H4KL16BODvN52ZgYjkP32T4qYQTd0mJh
2Wio8LxXnxRhpCfjrheQcy5+MzO+CfAYeWeoPxkwLISUVojART32yllhxdvzI/CR
q98FxMXW/BAT1uLtOLCOKCFYrbwGqjJFcfqaO2N4WvuAqwCbN2jLIIQ8HllCFL/o
IMjIslMefTu2Bi/ooYydrMoRjmfr3VzfTwoYJbo8XIVmjL6lvtKVFzUeo+kwD75Z
aGCiq8sh9sD7NonsWhbgJjJ1wufdV10pyrfzWkwa9XrTomCbiqiPFM94fhuiDUk4
BRIb3lJO4OJbwUlB/k8MMk5yrMg91tjnu3ehNNiul418DRjKhwcHoNNyKQk1wcH7
2UBLPB5qz4y0DOhes9juEhUC6L6zx+Ndqd6u9sIXA+hlwEnVajbTqvm5l7zNTb/p
sHpSstN2PXjOjwJeSb1B5WzP8b9wU+G8DfxDpwrvpBqCOGKyKfmSB0ZAN1JlFAr9
/BGFNy+qVZAI74oLYLOtyTmwsM9vqHKLIXgygo4Ke+LHNq73rVMWlJJk3HKxtn+y
zBVGf1TsfCOAxM0G685oPEbztc8SugxW7YvFn1fonR/BzvjCDt8o7MzeP2Wp6L+F
6202OjFqFXA9dGr874Cf7SJKKCBKyWtQ0xpe/q1sACtRnSRzfhzJyeueuSSw+tzm
1EQEsgWjHHWb6TsrviGB37++NrgqfaNE+4Rqrvf+ahwJPS8C0r4XvbfD5jz1VS1y
LZ/zBYPWuylrm6s3A1YwqUa1sI/IN03BBywmn4BrtNaIuERxc9TSEyTPe6gnO1K5
LriKVnzgIGJs40Lxv157ooSIpUWozlKeTCBnU31V9NXYI/7bym7jLYJoDWfrwxOp
uC5P9dWWTb8lFL2AQpDTgRw1GaU8Li5WmDLkOD1B2vmZiPzWLu9/zridHpJiO56f
EuOAlCEy972M1G8Ql5NYHcyy9U1FOHSZLMOzobi3VF2Wd82kfrTUclt5T33SipX9
J2Uku3qYWw0MplM5ivzGBw0/Ls0689K6ug+VEue/NK9K6Iy57EEtGDERjBeUANgB
f7rFQWAh5XLYD66gGEdSXHfBJgG9xIkP5dvSb3g8g34CXefEpo9AWNnr/jLJmP3w
Oo+9NXPIXJI7jqMklU4z3dFkrAmXrPQZrIQex5gm9BNcSfQrrw5M+vv9o7yPeh82
pnZhbV/3c7qH7KHRqvpZ2dUNMe2TRa8W0P8s2OtDcgffvR8AHz7eLz96w8UY3VQu
WQBcI3TB9wTsa2cleCs6/6cAbmA1UnOpn424Z3GK+k78mv32d2+mS20U9u+9ePWU
swIfo8tKeepHhasjdQ8PU0MgEP+ehKRSMieFKD5WHmjqejc8seQje8YB4WVCv/Ew
2HFAaS7xhN1vgpSuyYuT3whDqA6GPn6Fpb6YcWoRj1qhQIFUhYx9hkqifEd+klHk
OFbLQH522Mts5Y0MomCPzseP7ZzMLSSs3wSu9TQzKwZT5L/Z88mcfP/W0Injdx1a
2an67+8SLvcsGrsENPPD1K6pIgJ5Z//pPx4FxmP3AsEoqLgUeJ+xaUV7o79W/CKo
48cfaJ+/7Eo9KMtqWRCFDpmok7FIvHme93Vtpb8nZITh/YABnWd74NFovbb/LNnH
DJQzDmMHW/m7jrnSAa2RL0B/e8CvPmUa4BoZETNdphNQZCcbsmWUdUDGzJdyL5wm
WNY9jw3oJ72XMoDCjVy5d3KY44qMsUveNGy+MkZ8odiOznTbhxocWBUR+jDPlJ/4
elkd8V4520NLeNH616dVO+/ZRwO/VG59BBgh03DX+OdTaLqkc0s3FxRc6aMuPPlv
Ldl8BX2EeGTrZAlCBUc4u1Y5NwU8+R6MULYvBgoOOA2SkZT2rOJm7WWxxihe12GK
v9c/2aPRURW/BG7BERFc1RD3bdzCCsddbjhhGfuWGrNOvAQ6xUIYCKN0aIMfuRdg
w7PbvNG3KjNf/ChJ5abbZ6bOzBTBBDI+MX4W4LOH6o101OllfmffzuAyoC77EmfP
uqJi8pLTcMikuJl4KXfEuWzwsJl7qpIJce3dGtxfkJxg8hZMdmJJ47eVWpq2atJ9
BtRmjvHjK10Zf5WnLsTFxKp0xd7gUtTss83CocvvHffpSafDTYlEKRfjg5xDEtHM
pkHmXiwsuPfEp6/2RcASSr+clZl1Hhfw3/uQ/3t8I3dvRJLgLsOzpaBcYuT6a0/h
aKyrC/RWOfiXG/ByQ2vY2/cPhbFwXoU170Nzd760eeYtED5hwuYX+Ip60lgpoov4
QGxYircvuFK8c/MbLCFCLO+6FkNYdpl1pThyEOZxJGAZ0hZtFyFkMQG9fKn+rKlr
sO8OmTi6P06sa+fMtlXK9VmLMsBZs0r9nU9KlUBqXWV9BsVltlcXddXEl5yKnyyu
0nIcfaiJ6Z9UZD0r9enRC7JB1+NvoajXUoYFAYu3U069G6E7YPqvzaGgYQa5EWry
KOFuyxxoRsmcQOKaXoZaZttD3rnrR52tlf0AfjqUGjnZ2DndISNdEKRqE/RJxa1x
JTmXp2jZMj4rnedrX/dDxy1pjZ2eq+9YG4vjQ59slTskLSj4oVBu0+2YvNTXJj8J
6cWjC09IVf4p5Tv0D38n7GFbqKDCpV6oBmuppAadnPJdTdRwvHml20h7SP7SNNOJ
ryqb42Qly6rsQGEk3jB2HSuK1zRenu8WPunV3hW1H071/2RfwOq9yh6/q7agCNL8
M7xj7lfQYpuDcn/gNWW1ylGC9k1dGWayegJtoSCo/dMeQlOmV4q9jTHXUYmpit6j
g0sOvpU3jj8BkZRrAEFSNHeOTkSUfkYD9U/QJSyBysiCSAv80mnABHwbCtKItKxH
TYS39A0j3nR9MlGRdvJJVsJtuQd9ypl0Q262GjvdP7TGBfvV6xOH1V9hi/4giaWx
YD4OMGRYlMlFsuab9lAseIn54YQylnWxJR6UP6fbFDHJpJxUxks8M0L+7snFsTh1
TqwZlhFEv7WaCZSRX3Mr/U3/YkrpoUSmglYoWNaQOQnaYvKnQo1MKOz0iox9Ojgg
cHmx8cASFdgzuv/CsRfeg3oXkiHp2ARgRy0JZ8qw2M3dzzckXl8wz06uxA27tlfA
1fi9wq7iMMQnbu3wwSGpUiqLUwyF0pM6/69pAzrAbxmqa3s8APBliYBbT5rKZiU0
IuCwoHxfDL8sgzuGqBvZdfpb51ClbZg2ci6gtZUsMbey/I7cLwvCGMgTW+quhU8M
Br5mX8qtzI0cVn5eSK6pA/QXaf2Q1poSBP8k5NTorWMvOu4C7hnzvbJU5b0gu/c/
orvuBiJMEivFO1cz87mSBQbDeekd0DQ4aE5wY9QSmHZ0HRUPxmtxF7qUVp9VJnJd
Ukk7o2ll6UdT8jvqDjwI/zkBl4v0aVwCWlMeQ9zsGZxeJ6R7iXH1RdZKnRM8uUKu
SG2WWEHVlPRqpD/WIfWT6RKDcl+egM7waayVlEk2KKfWEsu2mhO1QS/A2dtc/lhA
6NORDyA8Kzmrf2t8DuurEvduw5Dc6v76pQb4HJbhYpK5L9yupSm7w1UL/uEFuhcO
h+KA3C+JQOy5nnPSCTeXqWKYiJmaHihJJw/SrKvicvIkdPAAxjX01M8LPHErp6tl
/+qfhwuKvIFTwwBsUKVuG6Ua9bf0mZuqsV7Ob0UqDuScZ7RGK1ojOGIKwg7UDNQs
9OA3p7KK3O/5z2DzzpB1rQUzW8Lu9NjHPffAiyMyxknX9vnmloA2PnXhB3HqXUQI
pGOg2+JLDlhy0oErkUZ2ZrOCoJ8WOd7EC/zoSXWN0o8+cJE8VGmw49Ec3BnHuw34
Xvb6cWl3J0BTgzzoSIJt8a/80cr6DMjMqVN8l4irGyXnpQCN16k6XF3l7WkBb4h5
4DhVdnOKNcGTYcjvXRzpuvzb1VkbGsCmwuglZScFBgDenGS5pcEDSQH7gzhBaHTw
GJXqIT+aY/dElze5ZmTm5lifego0UKEZkmPMqnFR3eFmPK7Bh/Bksas1HT1ldoDQ
lfLO/cVUUq5gCGzaZJqXLQAwUiXXSGECABeJ4X6WgMFX0OkPQoKAAB8pT1P3fef3
UCTTrJ2PVz65C4Pw7Vykmfi4xkIhEryHg1Rt6RVHetIwndC3KaKECQxOTwwt3ood
Gcyw5lNGpMfeBgy5oOUHev2Lkzt2YVTf85OrAyrT2b2+S6hGOZMwqQes9bgw+uTV
OIYgYoxKSStxGSXYrmq5zbCFP5iNbecgzSvkJWty37lpeZo3HttBx65n0q7Umgle
rF7wTOzCspbxo9EnabJInaZ4N3s1bf/e0IpDXI/fxxu6irUo/kuZ8+55soO8ORoJ
5qN2Kp+jFSmneNoRRObEGgWyVM1XV6cPyhXrl1z0RppG+hPAc7vr/mJ089C3Hmnn
Bf+9MZIbtaNkj1OpR73+UCeALL4rk2Q+TGgjZ2JPZmxaYfiuArkIFko25yzLwMxl
SPWMXoZwqWWWAhEES7FyTGwgAUaUamelKdv8uavs7hFggyNHghBayyJ4kh7mq4Sr
zk8TUc6qtN3HUideDh7FQB+tfWswacnUrrdYMqYOEPDWPRVkQIvaBaj44g6qdKHM
aM1Rjk74psIVp5VFz/MDc6qkVSoy7abCs0JFwYR/uOWPB456F2U8za1FH4Q2aRVO
AekE5Ovk+7T36Jrc34PoBUSldxEx4aBmhPpW0N8qtI1gnZVA+Xqrbfcz/dkOQ08D
wO+kjIxIaYSLcZeXe243iWQvFvaHnPPdEqXj1lANs0GS6oLozX6g7LW9QqpUAvB1
ASmkSkNZ7lzQcKgfuS1K+0fLL3gFHI+06U1FNdB3aMaI9R8zBcnRXO/98Hp0gZIG
phpFYtZdt3Pn78nZtdgj/SF5K8eZsnZaISk905gnO5yqjz4D1hCBtFtcZiypSU/L
mN0m1P7sdh4+oo9CJVqc1Pk1mHuC1iXiXGqL2dCCUfR8CYAlC9s68u1WTX39FCO1
geSEekha1/6kG1HGvKBx6X1Zi8hg+K9apgxN+zD6ctp95R2esupCOV4C0lQzrGEk
Wc2nxwLawxDGkFzfLRhph7BBp58okcLnTGGQxu0xjne/wbaTWdSRS3hvRtMqm8ui
C2W+AQ6dk7iPktcEVuu+8t+3VFbif83dMvHLnE8eukQ7uzFGTx9NgXbU8D/8jIxY
2Z5OIv6O9y28ZC/85G09Vu108xFgEfqDWVn/JdMsLanx78CwX6WiBKGeuaJEfP78
tHqtYGgxW59Cni0O/Fz8TXka1CjAHPqvKhTfVFVegV1idXZF/muJgUpun2mUJG7G
DalSb4pnyxMT6yZPlUVh9Kg3VvGsLlVLbKhwWiL4Xrt3Lag3IROyNskhFQyxfrUt
NlICP9YRzv1VLvR8iJnGtS23oozvvWGp3EFMGCgaLUD/mfOeGcMPfO2rZrgZPl/r
aVCvzzZqxTVqa80jDscTq5lZbHFNO+JFlHwNXU4kBnMVW0sPJUbvB9ZyNnJX3rA8
SYnaFkIM63lpyJT1OElAU7voAbYg6G1/TbdKQUns6OXzzra0OLmWg7QsiLeqexdi
MGTadobKy9Rv1Krg64E9V421u9MqsFdpHtbkVTSppU4juIj7HlsG+1R/Yxx9Ir9i
msZSBjatrBIvQZrOV+e/U9AYvCgJArSf5pCuHkiBSuLVRzyRT0s1FUCppIEDB2w7
F2v+G4zu76M8q9w2CoHT3/2hPgBlIM/COT0X5jYBUKbGRtPFARerywaH80hOBm89
WuRULQaaxc8Q7V7uPkQKQwgVp7mZJb0rSQUAWAUD4wbgJrvzn3Htl+9CH81O+ZCp
05d6eYgrZc2FCOGJR4mC1xoAbNc2Op2vziST9w5tDYmpnoi8E3P81XHCFsk0q/Qe
ZXgtsf+ugMH6z4hkjVqRnLCX8AXuN5n/AJQeHRacVnPMnSfvbl2twGyZdUsQ0quq
jn7uSUar3nABeeLRLFPDQ8n9cxivJput9JaT2hrGxwnGvixBlModv8KqBEu+hHum
DKLc9d+VbALHoeb2ydbFxUT2lULjOoOlypVZHTIxc9YW/hfyiHk8+XuH86xKJecy
wHsURIqBxK2Yv5V5P7a3OvXY2aISUeaPlBLZiO1cPDYmpw7vly/a4LzlPAmS6cOZ
LkRzph2RhssNU6X4cv5RGh7RJYOUo5bLagSyJW4n1LupiIA7OjLjTgJjoy5w3r2W
2FX5zT3WxmUUeUwt4DLy2zdqWw4yUlIRLFm990ZR7c14Irn3a/gv7aqHyBtkJTBh
kzFYJ/H+r1y0fbprNdiywGWlSmkyY9Pzp02o0zuPwaLxrVvaP/dG1RpFBp8x/hFY
m6l2glYuexmmNzpC2vHsaMGUEDOBtrm9k9cfbi2bMR9ttqBk5z+CTr5mgLYXIotZ
vZf5DAZgX+iBODisiBDaPHpcBRxvPstj0cT+ryaio6pWHdPvvoxld0YraiWgSYYU
AgYwZSi5//WgpUCeQUwU/1eS8H2ORzpA7l8xYH9oNsAWUz/ZRAIO9c9uTG10tzLc
/xRt9jM7YKs3rizqyu7y4UK/CDPjxcUNLsnnSdbPEGg94/+H4+a0a3gItRPbSv+W
li4CYejKeUJBlWVuKSA3DwSYbWeXkv52NbEtr7AHLOqbxIe+CWyfqE+c+i+IZfcV
gfAF5aUkffG4PT/B095EEE/fPj3SV9jHc40kL45BvTtQe2YJAd2zEvTVRNRzIvDE
H1p33LvXVQ4/7O/s6A0cGaJK3kiEGAfvjF5MvaRsNi0yV0zW2d+jaehdXSdWnvr9
3eo8hYCKgLFhPWXkywpq0KkjqHa+Z18AGyICmFTOiMcKFs+NTNEPrjZ4zjdktMTw
itUN0PPz1VPi/iwNunI/ty4x6Ou+02Tmn5ogxkFIEw+g18FaYEIeC3rfHauxVzdS
RcDnheNCLiZDMYS5/EIAL9PBoIu6PXD4NU7gC9gpdbz+Oh9w57eEB0S8/t3jQCSu
pKVNO7ptpUfJTCr00TJxLFVEGDgta7HGzGC2odl03VLGdAKmVQTRbeUIE8von636
8geqghbfMiUapAPM8fjbFkQvUhFa8wi/FkYel3pbhb7Xs8IZ8yxRZ/h8iSRMVrpt
yvMT4MbFfKN+8LTxe0sZf3q/hti9yRPUw+9M60GXBLLTcqk6Ia/wG9L4JqXM8ZB8
0SIN6r8gPI2YTaFj+2Ibnq/8d2M7UmlVL7p10ij0U06ZMk4Ir5bu3n3y5EgQ3/m9
aXMK73MSnU/XoyCTnXDPWfejA2KQhqWADvSQE8tynefe+Beowt/9OBc4nNQayC9T
gRJGgraYlmQXPoQfxVes9mIBv4KthD3n51G2k7OKtJ5x9YdmQIq1eNdIjvYVFTP5
8fnccT7t+ehQb2vlJ6Wxsf96q/mF+4PAoVnNlBGKXz8m2AsRnysbTuqaidQ5kx34
rhatyd+AnWHuiRQoJ+ZM1rm8eoCmLEvuYGRGqoOxOwC3SQMm2L3VuskeKbAppR5F
NJr6/64VVZwgq3KdJKcSumE24VaP1T8NqrpDyYeVbSG0qm/g+k39293EO2mxsj1a
eR8GldV3vfpUiGL+1O9wpZ2+RaIFeTzSqixaz9M7XoXtXRG954FWtcsRHfutgzha
tvY6Z5zxdo6NGhXYULe6U/f3nEuLwpmlUiXUPP3o/LRjr/QUdK+spTQM+EQZN9J5
lv/ZbAlTevKNa3EFW5NKNUwNx0FfOM3nH7hhy5wUCKePJ+O0JQtYiAfACfQ4ptf2
hSOYsS2tLqDu4p+r7OPfraukYQR92U9LuE6s19+AYyVFmuS701yI43+BE8wQvCPL
W4JtsewUa51s3tpltCXP0QmO5/PX6PN6GYdQwjjB5L7fRAw0IQQTWLeoqeqMcEl+
GeeNJNj9QTB0ZnIn3wPcAY57BxqeD8WtW2X+hyWE1TSL7Ki7R4FNUFX0ntqfcu5y
FEN2K8ufHhemEgHvjGWD3AUHkTShvuomj0RvxrFUMByrbCqA+cCEHuPJSS8lxyTu
++dM//PruJe2zTjvF8GN+7sj5hUrvLEZHXUedLXgN1VpqhA6JjgbaMex34Twhyqk
9T/+7BKZKkKPheoNvJeNNdcdIdcmil7fF7/1qep0VTwJ01fM3OjJO69YIzRwXX/X
ur3bPV/m/fy36ub+bnMrvjGno94fJca06fY1BIZfNzrn1VmmIUfs5AtviQ8EE4mG
60TqIE+CapGRdAXTnF9qUlRnpKzJe3L7rDbAlpR4GajxYrVOjMvuEOHN4mWN2OED
ZM/T1Bj+zKLe0mHTD97Zrv+QnwLbAbVcpVa3CcrJ6ApG4EG3yYE6+khfgiq5T93A
LuQetkWqh4Nsgk7I0YyvFOE0S5TOEEvSYo1JFO05i80ByPNn74jQmMTBuVRL5qZx
2DewAolQHNCf3qtdIzOC8ZLDq/Gqn3Ko2IzqyGiCPMwNJr97PQucWwXuNBNJTfZj
CnfNMKBqHuoPRed1wPwzlpiDKz0FT3UDvI7Rkd6mjZM9gNrEM2rTxTEIavL/2uzH
eNUC2pJ1sncEwYRRf/iLGV9OPcfk0qL1r2yRZxhjjSqNegTtfYBxSg2tfWfEtaSx
tjc8SgZea2uMGti/3uqfwKUjLiTAW90arczVUWDm4wLEQz6Mg3w0Qbeo7FbwJy3j
sWtxDhZpXVDuaIlWw8EJwCAkdhtB8ZsZImb27P4qFIf1G1g0VlXPJuQWYDvTJrTq
lnnoMVrsQKcTIa+YdO3zbJ+5uVxWPxkkVuhRjN05IzsNj6IxH+gLHI0CDE8lF2g1
s+/eUXXFe8AGXSpv54DpwmWjuDLLPBf64bfkE+mm1mHgioUM0J30tn5k2VeOqEcw
Ja4bx7qpK11CFNnEGzyQD2djH47Z776WACLQNwgQTkUf3sjRePKhd43FZFTECB4j
+ojSTM0a0FGQMkPrCIQepYbhT89Bbk1TC+Ou9zwEV06HkNZJuEwfr2O+Z82qdhqz
mw+PHaBA+Js0uZxwkRN0yx22lhs7EWF8Gxadmf1uKxxlxOByxLQmy6U0YEEcl4Kp
3qezl2S8UEy5zMkBvBT6EtVW28ykvyFpsCEjpKOwscUpkV0irLnu23b4yvZL+Er2
3pV/xn+juUF6EV+XHx9hupacUt/rTrKDPIMuPDzFGmOFgnLF03E1nxRGBx640H7y
y31ssUeSlu+oC8F3cZDSjbemeRDjmcBNUu0s+DyHX+Mw8QSGUqslQCIogVSL7GIp
AttsKVEXNJPhkvMvpI2LUfJzw94m6T+uKSYRZ85/Eq4+FKlVuqodmIF+CRMlgtnw
H45eT2O8Muag5TjAKg34A2T02SaX0lJmJAVb4DSiZg5sHfU+F4HNxC5FGNHUsUmM
qZtkViMhzeu4eIm1B0i0jfRPSGA/0Xt3BHXo7P795h12/oIOvNcoVtYQy2TSJLYP
oAbcDfcC2J/is/ioeSI1v4sZXatu1YKNCiiS01WrqetB0FuqIMwpz5YR/8ygp9qL
puuylv2FxC7Ks+iNKOYBb2lERRM4UU82snbs5wo3MfWE61r6M9zqH4PhnTmkDaUx
M/h4+lWy7wU4N7txOpdZXmwuRRAaxUYOAALlES7s0b4eUoxXSDMjs4GfUBn2ooPm
4goO4Pr+sHRH+SQxScepynBCysMPG91CBF9PhAvt5JT0L5D4Rl/HqdT4gGKnSEB4
24qKCt2fuiJWoXkXZX567sccTLmhdqNaBAFP9/JHLW9ppTIF7JMhPSqOuRmgbxmI
tWRVdh60XZevVtRmKRE4/VvSD2gsDjBcR2L0KyWzShGiTyoVlqz7+4brXrAha5hm
huFOcUHMZjxr4Hs1dWsnnk0aiqbDEnkzE02tYWfRVUhATgTzjaiy1keJO3NDemFv
mPh+88FTxzyCR97Ii+EhqlZ8CmGCooPmzh1CVErZ8cV/qaw65x1opu5W/TgJtdu8
vPIULllsO3ovUMMWr0y9ghiSXS8bMuj9O789J53vYwRePAPlzEzLEGA2yb1oWAiM
XchygdTUnJuhjDw5EL4vNeKS4Mz5z8jRYFhtDgdpZ4JqJB5ajRi+KeExrBlMIdr5
FdRirLgOXTvFLS+IuYJDZdTDlFv+GjQAe1e3Qk2yTPk=
`pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_UVM_SV





`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
dFqTIh4iNlWUuDi07k8K3apXtvWR6/+vjy0eDm8diVgc+V1K4DFnISAHGYQ3zFOe
rgiO/AMM4yMzhH29n9sPEaoMQ/8UEeTmM3lQtLMcb+h43dOuZRfFDO7pZ2xNTF3t
inievCj/WXerHAJtEGAg8/Xp8Wulg2CX0STjs7Vr3kU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 25363     )
52ymvTPYXTmlI4UagXYYWQwU/DzMomjkeMN8pfDcpCpD9Ftpg+YK7ciP4adTHRsC
m457hNyH9/MT0F96jFwuEeR/Nx9lRH7wUaNEd633Taut5tj36/HoyQtNzJ1dDwEp
`pragma protect end_protected
