
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
W9scHVkUKs1w0KUit789aYqnCNzsAas3aUiknZnhC4iMydATrr1R33G0tWQmLbY8
tf9xdiWBTtAXSoJ4jE0g/lJJH7QdVvw9LH80qll3IrAacn64uRpPfsA5fI3bTbg6
Qs8lYUW/v5wRHnwbachFEOubHDwJyUiGIwRDqY3bca1xJdL/uXQ7QQ==
//pragma protect end_key_block
//pragma protect digest_block
P+4llOVywvdyoTqmQb3GWad72Ao=
//pragma protect end_digest_block
//pragma protect data_block
I0Ph99G++I43zn2fNXNXJX/HYOwAXxWHYsWLIijP1SnwQEoJ4QP3VZronAiW4wuQ
DqAlHqWxb2cB1UtucF6o/9cWSqLbO6IXbvNJDJ36/LhSXmliwFgzEsQrFQHNmX8I
Xf5fLC695sdAv0gqzXr3Lxl7/+AeBlZ72qdP49OAYBM3SZO7pwxA9swI0zOBnyBg
LjFTYuLxF4kgRtMGfPoOsnXRaXNyQvco6gF6vduxqpAx2aNzaGBRpjBQ2qC/kMjn
sngCLPO3XZccuHioOtOW6toawm3Njfom0IDPxXXIgHeKglBhjllXPmD3YfvMZjUy
b/EzhnoZeNduNG9UCR3InVryw+UkFTYJZeKznDjX0OcLtJSMmSyQuVZKdOmH1cxo
REK39qoow0RQ9iu2GP7gcQ9Vd1wVN7dZRmwKjSmqK9sOqlVV9mMG09U8XJ98x6w7
V75NYWiHiVTs1Gj9cYdxe7f/b8oWcSCBcMd/FmznO5+szUw9Ks/Ps22k6pJUKG0N
zGUHTgtZPVKeuHAXdvIcp2sD+9i2CGvMICsTeZT9Oj9w4j6HGc4BNiJpTqWp6A4w
SiVj5AGsjszop1mQRgeGzuuEQCY2H5OzJ1VxfrWDA8v0zSCYURmLdIf97lWtQd48
IUkrTZASb/KZKIKCXnspXcRKfp82B+GcNSGq2k/yIqF45A3SDWxMOcIwi7CTTdd+
bL3EYugsEDszxtzlyS6bVjMSOcgYnmA/7AxX3aLozAMBLxq0OrmvM6xwH2GuoT0P
8lBusbsHHXVCMV7L7YUPhn6AEDP9aGmnzUlPIbPdB94Sr1JoIfzSy+lO3r5HHzjd
GmZkXgmfKoFgxEpSom0vt6KsKfQGYCIAtUrVx3XpJXY7pUOwB5HcQo178lqdNH0g
blz2uTM4Q5dke9dHznjcbIYbL7yn4dIo73rLlOByLDe9ia5+aSZIQwCYDPTPM6dF

//pragma protect end_data_block
//pragma protect digest_block
W2pKL4o7Ubx05ZgzNT0hWwuC5uQ=
//pragma protect end_digest_block
//pragma protect end_protected
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
9VEhKrJFd23HK0KyZge498JdrANRzczZCxtP1qod+mbgkjlHR0RIc6+WakmweoQM
Gwac84hYyv38g0/U3otKYk85iKiInuW4y6VdDX3bx5N3WyRi8K6+z6LmphWlzHyV
coAQeZaARCMT0RgZ+9kwrkvhu4CIACo8ro7/FtSIIOUAq0sfqITcjw==
//pragma protect end_key_block
//pragma protect digest_block
YsrWUALpJxfp1RGornTbk9/RY+M=
//pragma protect end_digest_block
//pragma protect data_block
CsIrzPIrQh65FTOv5G/rVfO6jF4y2IhFqXaNjiPqYSPIomFnTGDVYOPS9nnPo81g
vXQMgJDLQyb8Rftk0yW9NDnToF9LeCl5S19N6QaE5Tmukg2nm4pU5jrreUzXT4Oq
Z6gQVhI2G997dCZVU/MTKq+HH0S5P6CFQanfvOokqIF4S4fSgwmsmnlAymVqeXhH
qJtQLvpfWwOFmCtzM+SR2BueFX+b211/YAbffaUjduxSnTFRCiLcKxCUOMvQJXTv
6KBaIetOIdkJQJAR4Sto8yi1YKYxIKcQLCaNKwUhcN9QeGvoayTYYdWenSKbuN49
qRU030UgulzbSMx7VAmFlDzA6HmnTTzx7XwBen+3qwNpP1FxlO4u5e4GU1qQ6IZq
Hd7LZ8GS1n+Bbkz/cubsz2Dm0422T4rc2kwZjcMJM3Q3yMvFFOd3yxKHDt8KZF6R
NMa/0lo1n7MxNpuVwMO5V5z1LB76V13JS0KsEv5qIvRgWhKiSwm+FIlof/q9p1Gf
/pAst63IzCFGC923OXiy0ZVr9SlRRBd0vZ3Fc9W36xE=
//pragma protect end_data_block
//pragma protect digest_block
fcpdVtCjBDuW7pyPv+qA0pBOjow=
//pragma protect end_digest_block
//pragma protect end_protected

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7o619i3FYZfV+wfWxbN3oExnPk3z7zLDh6oEaIhxBPEvMLgV3eo0sSnugWUWhJcw
72YYH2SvRVmJn2j6zla0Sgq1EL86y4CmydCTqRMdOAZBrJGlzBARRr7Bg46P1ViG
WsQvCSdTgrViSEV7XL6XHUXdVMnuSLejDTj+q7g35yRPkN9irqxnnw==
//pragma protect end_key_block
//pragma protect digest_block
jnuOkOALXUj/5o6pIL4vP6sTols=
//pragma protect end_digest_block
//pragma protect data_block
iLbzAaC4KKX1wmimf9aPhkmD3Lf8KhPkRyKnCiCpZLvtZg1WPKA8nlws5qEvB1Zy
hoGxZWh/ImaUJF0y3LquG75FuY0yL8tjnLCHh7AfmuPipgOtuHQ46L8uErVb4WBK
b9RRqQJxpSAni/ANt1AFyGllii99/ePQ4Fwn2bHe7PV1TfdGXV2P6ZBZDY3rVEk9
or5Wp7fW9PZ4OnKrD0jMQrtQmuy1gDwQZZYVx+sX4xa5C0uuRy0ZWPZ/moGvzyag
RQjmbqTDi+YSdyj/elemA/ixlUQgNE8WDsYztwPexF8Tdq3zQszHr8qKigW2bYU8
oPMfIyfMlgTuNw4Jtbt29sVY5IxSnKeMniX/QWK7CIbmWf/TzH2uQa3l307VPXjz
sEYzqy+ozGWZQVfVsXKiMZxE4hVJnk9mHar1nPZNV44qM2db4rxImFBL9RbiN2nt
R8vupHQGbs17CIMHTB1QD9x3h3aHfWpBqXzvM2gNuWfjncY54G3X+D5PfaagOkLb
sC+HD+tWYOVQh8Ojoj+4rw2IHxCosKCzzuR2BzncxTqCtX5/iY+Bw3ryFz23+fx7
+25Vqo1i13RaSMJfUkPO5chZmplpxFxEO8wF/TKtRhyD7uLJKPbHm46HPjx2Yht5
SAmGpvwi36WqGSeHgDd6b9w9tBbLnhJRw5zi72DaDNIHoxtUsvRZsk87zKACmxP1
Eb5LB89+vtnRHD1PGIB91jkoFow2fULsSo9DDgXbi6SiHHaSCqclnYmfD9QDKKlx
YhHUNvxCrqmwMW4QmjpRjhl80/gNScNB3dxztiTMgiQKG9GUSEteUqml8LAHzkEK
ws8p2+5lJRIyzKaHXm5UMQ==
//pragma protect end_data_block
//pragma protect digest_block
Tt1VsUAoT1c5hhIoeefXukvw9BE=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
jMhqNeuhvxcfXG7a8pAYPcFsjDbK1dMlzooSBBV9I2R943QcS2pSdSUCqg7OgqdH
snu7cdWrw58x9XHadD1ls7pFgyN1BvC6i9SC26HdiONvr+2utOBhbyHslwoU+agC
rMx3uugeuHVQBkd0jrbFY/3sg2OeiZMPJhoTwLAxBiMyZcjRCHZIkQ==
//pragma protect end_key_block
//pragma protect digest_block
LvJ07bxUYMf6pwMo5SRNLu3BE4g=
//pragma protect end_digest_block
//pragma protect data_block
XU2BzWL4Q11bRj9vrJA8KmE+7lpF4EpOvccqxaT9g7R78EUJ+mcmsGvjz1MO8Vov
IL2uV473ZwFrDL4PI1RwvYV2WOjWxWpFkg2Qu1KnwqmK0i1zLnHbtuvvVhrdDCwr
2Ja23PVpGI8P5sRdJsdoTxEgRxlYxogJXaa8t9+ihtLiY/jBKsU1PQawYSK8wtp1
tQeWAoSfTbFp226Mrp7bMwS4qgmiB46rC1lnCTYeAGHpPu6j1dkn6Jdv7ertRwCh
KNclyaDJ829alrX6oBv2rJM7fVUVADhkaVhTYM7lswtSd8DS6d9B0wPUdoGxKBpb
jpOycB8ifXBXonHto1g5Nd7/1dreRVi9i+w1nfHOYTN14CLOob6sOZU/HzEn9C9R
NUDsZoWmAoREZrPq8PQNa++PTWBEw/WHkvf4/W1yDSDcI5GCdqABNQexPA9jwoDY
sTPxfvgIcUZPy3+zjPE23yPTGztGBbyorCRYzyRgqq30p9i37n3RTPkI9jm84dS3
DyZyehyvAnVXXcyvxvHk7ADPw+N5eYi952AuyvNQCL9JaiXdxpwn6l/oDsDgJm7g
367Wt06GmjHG/n8KYZSrfKhkP5iRH1692M9x4rUxkxrjVSVvC8ynwjTl7hETff0p
XnhW/p1x6wSU0wi9L3fN9gqPkFB0QPanj0QsR675N11ydj4FRobYKcYK7tqArIYE
D2Clbh9PXFZlCHfraYMk/kyU0RZKlH8q3BIDr9QoQgOvICDoU7e9Z/Fm7lC3/EvM
thyfIVMq3AH0D8iMM4cI+WKhm2lQBbsvSEH/0jGpo7qHhA1g9ajCH5TMKI07sMcy
u+0D3DjraKppczgwNevUPx92FB0jTFHohiOOvxrDv9FkR0701HOqJqPtQaDkGBVI
aAtqa1kcPBOMu/arHYpaPZ+wB9mKo8pstautT9zgV3YCJZ0sIvQMSq826bLqQBBH
PYwgzkaToLo1UdoeNT9JFiy9iimlWpWF7ZoGQT7fc91nAIeDBMFpWIRUeq0tHGYO
D0BmPXJ2XfzYAhPzPp+bhqhobd+924Lv31+vqXLr2WEFdvyZ7fj5To5GpXzOHNzn
WjQMAkC+Krm8kK4tsdyyWYvuzxeMQXU1ujbRuzuLjfXXSbOIsrrYmBcccAK8n+ex
HYStaO8dNrsuJtBHmAyeZxiBs5HMZQgGi0gNFM7qI2Lsw2TJobQQXtv/qmoS2yOL
p9LOaL3c0QcCaO3/uuyL3N3icx6qL7SnSCuyTaW4PoqqXI1I4X9TeLJSHgRioiqa
lspkxL0rwNCi/i19NbWz/zeGvCKhMxyBU20eLT82xCEzubpbK9bqgugqQJq5sUxD
PS6mSPL1a79PAYTJXlJrO5b3JKJCe741TRL9DPrnU+zSQgGl+oq1KFEz/2DVD13h
RrzoCzEMYYj/xK/8FYG5IOfdDtuULVslrf2arDpPHo9wuaDrBs6JC9MyoxqkkFx3
XuQOkRVIYTswnXgbszuJ7zXicDVeGF2BosSWt4xc803y6JGvMigMK7gcb5yGKu5H
oKV439YmYuBJRD2M7BojYieZgJIqJfK/RIChwhnOpG2Jbh28TywBUGnjX709p48s
/Db0xW+kPMt1FIIMfKjbP3I5+7h1W2UsXANc0OyLsfCJW4PS8J+iR8eoe2PaN5H2
eO25G7LwgpPO3JGoHYyEvhDDwBEgq+zVkV/1UG1RtX1cISaRSDvQJYFfArePdDFO
RTSMdSw8YkRLxIkjUPyEekQVKucQnnYid+cOgtYuLYiqUroPqtSPhhbRXBeBt1bM
vjKPFrMqMig35p0LW/C1qglT93DoudMult25FrmCHD8CArGSoK+fhza0a/lzL322
BRg4wYG+nQuLqHE7/A1F6ZRyUPdMGd4Kw49Eig0gafXU2pnXVJ6Nm/IvBi400GYU
HlmjiJeZaQY0QBoVKfRkkjIvtj4bRhFH0sHPaVsQZJ23Po/0QrXF/uY42EbH4RxJ
cwpwuFR3gShsiCt0B54WPLxvrWtufaNwW9edgtnobnNa1fImxq7BYa6x9tvURsta
HR+nn+ng47dG7F58ANpFdGtlCp7pTRnYzlCrkQN/CPNQrKB5FCtjYRADDlIC+Mbe
bgEU8AG/zcXT242cyZ03rfVst+lVMW4D/VF9KEDbGgy1Wd+SrTJkdB3yY0Uh4RuM
bowDT+V8olo6Hle7cE6oek4nzZ3xsuv90ovW+MPEAvDe3yHwGkgE9W+gch5pa8R2
3/r7ucVMAtNjkG6eYi850zXQW1QztnkPy5w8HTxqMBlg31tKZEZQaulJ5aiiHDHw
RAgmss2cCsKFnzzMlYRF5GhsEhE0pdPY4z4MTfcKRDMBEYHpdeuXtr53jxyc/C9h
gjsW3NdXcFyxFpd3TzqErexEIKvg4JLgfTIU2C5Lh75VPR88gYMqzDBWx9+joZ1F
Jlh0odkxLyoBYVFC7/EQWIyptTvG75dY/t91uuAZRqdiI4xkCVQji0iOhX14dj/u
4BZlJdv8e+m9/tmlYnuPAvQBeStly6nmoSTe8qzI2Y+3CfXg/6FhhecyVuOY0izQ
xemTFZs1Lfzf0ccnXVDxusLAg7fVcNM3hMcskHr7fnrAWGcFfYoQkqOptGKuTnrK
eRElTi1hqhDgx+W8uTL+P41WW411v9+ZQWL6JxjqvZ+Sx3ZBsD/o3wPco41Rg9Ca
ZsNyikd2xpg9suMHKSbUazH/CyuCjiSc/48bQbNSv/jVuhciN43M1ihxQ/VmJrGN
fDRzcDf/BmBWzE188Na3eW5nQPvG/iBMS0zuJ/vUuSAS929BgryDnNej1+inuJFw
key7TmIPbwKBK/IlBAnyE1oCruVzSbgBfdYYeTjPC4xIrBL3fpk5c0y1Zv26yd0Y
TUVFg8BMxW1qrD79hzRENUF9yUdp0SntSjDIDqSHBwgFxeKtWZtQpyTvWSB3WxpK
IGUlRjeoRfguH064eiSZr2FhmvP52KJZ5wkxulUgp8CxPhu8C755vNJVNzZoZnwh
hmsXOIu9Pfboq3iOEp1TeL3ko1sIOMmhP6VlfWAT9dUPB25bb2lWwMRHp2rCV8Aw
AuEhUi3hZ8Xb0mLDI7zsp2g2qW8BtTzDlLHs01HyqxpPMv4W/kmBzY7AtUtw1x5N
4IiSb9baYLA/6qjF1n70BWgx7K9juqWeKTfLmetKIJ5CeENwQZWmMQsHV2x8szz7
2Rh2dpjGvP+8QrhjsiMjIHpuv8twD2fh/RKtHEumi/C9/wJfGswyZ40xkG1hAa0c
AvBJg9vLrJqmV0MfA/jk6veOs18q5q/DUjBd4pACnFbP+Y8VhKkXtUWI6hAczPx2
zpaZdURtz/h2LzY5yWX3DYUXUsartlIL49wrBjVsrAfl3qdDDu2m1HsH5XeAzK+C
9+YzhyjRo/KGLK6ati64wPQ/L6zDDRWdnsczAdZLuK858Zm+csdjdWNW4nvJJkrJ
PIBBYlav9TUa9KSFFHlAHqDaKpw1WmTPrwvESKdZmlofiIuwJsvXHUz/2F0M3mFa
JWO/T8xk9PQpleOilbPFcIG/bUWOt4xhfbzSm5eMBE/wHr1m146iVrNWHvOEyPdk
5Put9qIM7phUyWeK334ykn2u9QkKX+85cAyfpwPZZqBlgwSY3aHSb2C3Er79kM3S
kHtm3VEYkRz3w3ZXJoGRYjnOGnOd5lAsKjLHv2ZO43BONFX9HXW/mjc58V6m1T41
q+PnSVLRtBNJ0npI2OD0bjNx0THnPCCNZUwZ3m6L2PFgzTYNHKLYiKoNNXJlcQIA
CvVe6RzLVxQRy0TcR6vt87wvwqJCZrZbd6+3Cy3UV8TUmgg9JJFA/ey14gV1AC/Z
1L3Qh72JW5IZqOfRFiCdBOkZ5nW4ovkQiMxIob254TZ9Bgv5oiRHJgWPfH84p76O
BKKF2BxhFKMsmt7RLT6R+jEdl7JWWO50lMNBVivsVmvTFEf14OB7ezlycThfZZAd
sFfPxSfq+NyTSosy3grqEXHHkZtmwCVAd16wIwH+Qo9B9LuHUENyjaFivT+5Lugm
o8LLYJ05shmKoP+Yv6nbB7tyEJxVcUAHZq/uh1VdniV+ac/4V7I88ejkRvg/tjQC
BCjSyI46PN25VBgoy0mX60vT6NlWRt/MSyWoycmwHvVY2inVHRP4365VxoZriWX4
RB2dmJjcqjTgrEdz0VDSwQgc6BCJGarrXwQL6VcjBn2KwFAsMyDbX5cK/K6p5VPx
Wz7lcLn4LuETtNiZEPk0Z7md489yIKXRvhstUPgTgodzNh9rcc1z9wwnhmgfKUJ1
MvqAK+AHXcTglp8kdss4JneXlLR+mszLNDuBIOQ/c/qNKzUDjq6nzpTjO0Dyk2sD
QEv7MMiaArNoGL/HPaG1hyYUItfKADSYrK6G33DGVt+j5RSFQWmDof3POyVjCQjb
l+XBavKnt1iGepaGhW7YXyC52/1cZKoQ/ubeceDn9ll6a4USJreQkqIfv/8t7zVA
Swl5ko+1lR2mRR9Qztl3eWTJPBKapOTwETBTbdneKEZ5yZkVmYuRCO15mVUdXMB0
PvgdHx50t7nMH8IZ39HyE+++6fRzwJbI8wkU3pB4C1lmKt0zQJdls5JetZ5+R3p7
T6ke2vs/qTfW8WqZMZio/2m5roymr6+rwc08Hu8vyj3+v+K/5qcFHiv6NyUoDU8q
CA+FM+kb5X65V3ZydSZp/zdp95J318MEUFN1qjxvLOGjsRLzANAyVDzFrrix9nJw
aZft6oDztt8s54UmOh/QuEZXmSJR7JWVdqn/C7ayeuGZBxy1yCPZx80A38GJBiPk
o71SSeCHNCwrO02gF7e4h6tiAf8SxiX2kAT2wtFY7uCMIUtGmTItLHXslW/vbWyn
XNeRlzrLEG8K2epl33kleTdKKP8Xn09QvJZ958XUBVCd4mhTOEbqNzpqwUvJ2dxm
lc8p9ki5gFyAheNdOzVVuNSfz1Xiody26jrovPW1tOZuxl6DLiyu8BE80+JfyyJp
8thv6GTY33C7rnpEMxfATsR9+gXMq2cQn+l3LXXLgZ/q+sEnvmjjDjRqOWdws8XP
vC6A6D/gXyff4eVBmU4ewCXy2fRfzA8d96apeMuFvwceF+FmIoPGDBQx3soBw2Em
5jAUc7+BoB33zgwmHG+A+nx681xDb3J8IZQkmp7+CJ9F38VXzPz/XGeRw2ddLzO+
YeZQqlDUT4Yaz8haGLYzrK8g55kyh9de82fU5gGcsOtcMxh91ibm3tneeooOXV7B
3D0FQAom5i01P2XF5dSxeHNhTYv75cuKLnz2lirxEEGkPUvjj5sDPyyGDLP4RL8b
59D4qVLPFdkwd66SZhXiIjsilDm1416ar2/FXuGT9tcf2+FRoutgxZQdoSD0Fryn
3g242L2wQ7hqAeEGMkhhhbEPLs2kiQSNZnJkqfID28Sx3c/IH0aT9aynBp5a2mkn
J+M9HKE3Fbzh0+il7f7o1j33S+Qz9ZiCMwzxvWQONhm8wdhiAd9mUzoSbyQzaZ+4
D7QuVMwMOLzyTjYf0+J8cf+PpJOpJAfYxzbrycvNuQFOVETBsTH3zYKc9XK64Dz+
oByg9Yu6V1y/oCsnxyl0pGGamLjPn0cU9yJR2oB37BX4r9Wza3z3+YhQ5NECPQri
fNzsWHAwa8OZqlB/oqZKrpEdbqYjw02VpkH8x6846iPe6XChOIqWuK1x4ftLWjlT
3bqQzM/FBMXtHJQaHDSaTdFGvLcylyLc3IfAjsAB8mlgO97YtDFJfhC/KDlmSrXo
S+7vxla9IjbzOZa3kbJ1FVI8h4vIIYjY9ShLfI5e4h9RVbdIlYQ4HlwsjG+j793y
eJYxPY6kL5W9B32V4a1SC7rDl3A/C0VXuKrQhncUkAXO/QEfTW6TgHWwwj5NOpWR
TSiktbPzAK3X+CqR2OO6eSAMZrUJ8JfGHnsJIotl8eBlWLhdrRGcGN54AvWW0ju3
kLGUqWimlV8I7emGWt85otmTtalVoQibCnyR23UJbol0V96U1GmNpjMKeF46IZiB
Xzl0CK/SgRe5jAlWNFB52KKcpGAeJE0vhyzGhaPQliYYgx3koF2tAvV2JskkWCfH
lrrEKQlsMLkhrIi3Cs9kun9ZpPL/sF6MZ6/4Y8okrR/yI06ylzzu+vh0fFtA/+Pj
cCtRh5WvdJLssNs9XxcgLS8CBkc2ReRZeYQ3ojByEzlL7KTa2i6RoLJaixqH93QQ
G4ctY32y2Q46DAJOg4gb0IRNWmV07ZiZrfzPR7HzK2U9PfZdfeV4CtlpGFpjR34Z
+D0oyBy3KARsTO/QKYtMqIzVTUDRsRbK6HGTdm0NzUpcktWDxTh1T4llIcbp6KpE
/vxUX1PR7lPREJi6KebkfG/bopGoN5Dsq/97lMM0TeyV2F1hSro1yNnRwGaLG5Cm
XG3WzcbcFInEUxWvnWQetSX9NdZ8YwrGFiSlNPrJyDg2+QRXvQxA2BBqQxx9qTCw
Za4GZf2OXQs3uo+/JfpnfZbm4pTxYIbd5IsHNdYIdIn8t8xVAG8sB3k/R58RbYLp
GTDjOzCZ+7vlvnAFNRUxv2ThdZKMtsNRirHQILlB5UeC2mAXeFei1PtUdCK/FMot
V9ZbOQy2hwZGOwmSxRW+XuU9X9JvNtOX9IUGcKIHymFt/BGiKr3G7laF0pgGPHP6
O+tSmcy0IvHxiyW2w7+nmnkAHKyI6GUL5kI1YSYTc5pwIAcwKZYXlIpRBJqgLJSC
PkcRPC8CYWhqxKggEZL9M3haje8pg9irpQIlK6+LVPCYxDsggs2e3v2INzZ2XJGl
Wp2hS03qjAYU54sGdDjpEwc26lNYmzUofQMHdGIReeSAm5cH8ZRhazm8nx0Tw5rg
wsuFOkN/ln8EyK4i5dX0IJBZFCTVWbqlcDr1EFYdMykhDrGnN2NGyzZYmfefmCkO
QYfLBfOTQ8sZbfJBpCclFGB7qzeU7Le/vXLkmbw+tB6h5RwQx3/kxTlbaVkzsNr4
5hgKDBsGzI7yQCvIAvmwmE/DdcYCnPC2Q8xalMrZm0aGHAh8O672e06UFqMD9XJx
hvAdm6MEfptCpeCYFcGAMCfQHcgb5CUjtwVgSmdncdOorWwcMXZwUPWIekLh8y5d
O0FMFvXp5+NU2D2LMJ4bdLYwsXTBtEUUpDIyTYMUJ4TiMKYZCgRSI6sYMAas0/Su
tbVP8eScJpnhqj+EO9sivSrEyr62SsuHAZXqe1DcCYU4u0/Nr4lAF+m8j+yGwOPZ
HPSSGLPi8Xac6v6o6t3R4rWy25dfqzIFRwSDOy4ZBiGEhXJJAMjkNtkK23zQDJyQ
QDSCjndRgdBQ0or7EifJrm/82w6nZpGJLNzuuMlIJnEIJA/fU1Zj86KaVsa6Bl1h
4DyphFYMZO2bOMirZ3eQfDzUvpDPKQR6XWsugK873IFwax1q2aRq9+F7FlPMb0Sl
2WCH5lzsZlfmCUDSr8VG41QRPXL0JOuh6ZUg1WzWXyAp0ArFQRlntVD9CrfQLe5D
M12FH8vu1DYwq5OIA9njufNjDZNbkfzjUkV5RoNHFcrmUxCZktlr3fzZXOwqaAiA
v1WaU2lDOs0KeyVY0VTTNCpLxtuGsz1SUNcU6ACKUA8w4Gpc4yrj03bN1niox8TH
ln6heUeJhkd9lljswOS7Oz2HsPIA5g7KvXWvE9BMwTOCfmcXL6cUhRie6EEukkbV
gJcxhPIB1UcsKk7R94PGnXA2ct1bOgV1G4iddnGwCFbTBBu7xSqMDEVV912YzDwz
j7GY0Z39kwZvzW4CLsCGeDqWR08ENW83DOIgjDyO096lQrvofaxEbjO0UJq/TxpR
4khYxndTu3QlEoqcXH9CeuR1l+XzBACt80d5VFjSD4JFeAuDRnVs7mxZg9HrcEYN
VZv04WvB6xK/kEb2Dd3YApphjsWWcyR3+zv6hieuAfM8o2xPNTrN4pCdMAS2yzU7
fnJ7dVArFhT+3QHL6BvclVqCDrgVCvZ3CzbVb69hjTGR1YfOmChYji4mVx37YrbL
b/0lqZ+A8rDxChtp/WkIFAAKQRKXn1OaK0cUk2tq3oBApwUwUzTSQZyhbFNrR5hA
9tX8eHCnpCpYXZwgxQY5RvptzgDhovUGP3QZKvqg9lOor1FE87t4UMcaH+JYTL6l
Ohl512GCjxZtOgNX2DAMNWEU9EKQ/xQof0MiqkfaC+rnoRBLpJuXCKdLIDm/7mU+
L9GNFyUroJDU7vzmszqVhc/4DpI4Tcj2d+ZOYXTXeoss3Us+X0LnOvUq0c8jkZb+
WAo8R/D0Yiay0YHIauGZAP9X6slipx5vheMiH1c8f8IpQEoXO7B/I08r2Yk7D5yT
zJhiVZGZ8VdSxJNGFUvp0PZ/VwKaXdugldbomP4aHDPcsBmlJ4gtlFid3GJGNzA+
zJdtBIDm0LV4icnkKAAqr4D4gtZzMWPTEov1zCBf59ztICfK8kr+4V0PGBCEkzZ+
N2UFBcbz/kPBbXzyVS2hfJfvRZMgBIy/XONxzXA1fT0Vd95jMGv+r+vJUHK1Crdv
qiBw22pZSEC8jqbg5QOnALC57jg4EzqyMT79V4CLWvaEXPMnjDYYe2fj1XLKkL8T
ZxNrlWc1wiFFDiH2Qpc1NTzOmCzvvqfCX5tGD1J1tSQvzy2rS/xrE2mgSJpIEkKH
S9DNPkoYvUHu32Rm4jLCQ3NbXgO7hbFyjYY2YEOlwvWrr3j9U0FoR+RikM8fRX43
XDKj3sy/zf1CsLiPbBk/QQpGGQ6awEFoVX1UPqmu34R73cUvBqDUWLjgWjp9CdVY
92syDqtIGfE96Wf6u224XLW/MHv4kdg/ajs/7tOcqwTyxjTRTVD92TpXDbHFcgs3
ZhAUT81I75NxcEvQhuEH2fxL1fusjzSpN1K+TBY2Y+Fopb/dlMXFb0V2rU5izXCf
n1QXQXCZFVAZ0yj3Z1XxhszIxAGYgHVzTZP5tYI0HJmJcAapL5UGMWi4yuhW/liz
fFmrxhTRN0fVqhb8HcZ0y/on0eXN05ijXFdkx8WZVHgUvPrn4E27+18dVu02VWPO
YjZLRf5glyeuOD+r5Hnpf6SglpizNCPPDtjWVt6VNLAZXerxo7ZposPOwszdszvm
0oPbM3KqT/GNAfl4X6sh/QrqmWmJXH9beU5KOXiMSaJPqD7rK8qJxHhFnyzD5sSH
hPdGIpMd55s8pn9QlhJgR1vpI0F2dfAdzIs2W45kyoa9Opd3EqJAlqIVPC3T27Am
35Fla3E60q1W4SQrn3aTNzqEvD8JhvtPK/MkssX55DsoGy/zqNzMAQtoVAsfEesP
CJKEmqKJq+xKVLo4o4lgvGn6tJn/3sqvpNjVRqHi6oH+1PXAfa2YsbiUsNTHf7dq
SQRKVF8lonsX102htH2YnLRqW8LYb2yx4Rm1siZqs/ve5/tQXoohvk1xCqOHPxDI
Lcxorv563sw862FuwCb8hvdxS/oHuL8qnceOpwjFhdgW7z+wMVHLpYRutH71tPXx
7Deegk6cRKzIc/AG+wXGEqFz7YsRKDY7bZtzbevtuvscCFXBalazupA+H2TpbUOp
4r2+EiBgkJe8vnHEu9MQdN1YAtC9qEEtS8mjLijat0Y2qYZaFJnRHvXhvPx9BY1r
iY8pWIts0I/aHtfHo5QlRKEh3HOS2+kkng1nnx6C202o6IcRn0ciXI8tujHIpB1P
SSx2lHUwDlza9fUEWK4+xmaM3ocGqlbzbT6K6aaXZKw+DoRq/w1TW1IhPfq4rfkO
DErxpK+bW7c2qqi0RTPzeu8WSW3a/UmulnLA161UIQr5HspLwN8aFQPvmBPdypUu
/SeZId8hlTJ1KzaHLGbODLpX1MxyFGZX/FVANF/3g9LApKycbcu27Anag+nq1qJ6
pOxpdXH6LHsx5wTocyzDy3ri9yyzQk3SPbFQz+qCIjhEggwQ4rYUV4tRBSbddUMX
WD8D4Q6ppSZpZ1xGNJxSRCp/oQMA+ZhLLRGCaCIY72D1KFLljAc+Me4EwZB4E7Nt
a5kI9eFpl3cB10hQDz93idefo1WDRHCfLM/dc/7nAF+oKpO1qHdeFz7CF+7+Y+jj
vHm8Q3uj2JZA0vC6+Ga1e69pc1wONJYeNmBShBQklx1UGKa/Nq8cErX3EDSU9htb
hFuCxtMEaklq256fWo8ySuz1BdLvZQ+eWfa5wGtANz6mhnl1rImFKsvzOkvK3Zrc
e0pGZ0Tyd7VimE0LSZjhomKAgH9z1JpVetCfMB59X021A6hm4Updc8ZV440mdxAm
XXZJa0ZnZSwlfOf+gxJpNjAK15lLF2FS10QYtzKKcBkvHjTHBUBTHDCMIKSYsDKE
AJyy4vHd+6NrAMi8HnliF5L9zs1B+j1jOobYYvndCAtGYBO2oH53A/aHtOr9FCai
qbqyNyqvWqt9NzvKNkrGVv4avbVXh/kKX+NvS8mmu95u1nCLf2kwI3Fqfzt5ufq+
/DAwsUHb3gh6SZqnytLb41/eFAi2oylGQ/MdJyu2G/kLHxvyslfen70DX9enkTMn
VBMUmTnDAXS5XuYrFocbQ67oYoig91GuIQLhg7OsDPVFnpEmqTmQhiFc0YhMS0QI
bqx+Oug5Ejk7VQVEDyyoSSNjwNPNqeUzxDFWiNc8MINIfWWV4XJMp39A5/2fpkoj
vZ5i8bQVkhyqMnXkALsQ+m6V619BRsIulSjFD6rBj70Jh6ozAla1VH6rcEITwNsO
dqOfBYOjlZX/DhbT+LO1QqC6G6TMqVs41yQmKnmPgRZj7HG4f3HEXBNHkEjwC1NJ
lYeRpWURxxespRc7xkJwLLUU0Fv4LO+U7t4bGnKcBQjRxletIcWFvLawQOoDU1EB
D+XS7dPuX27Gpi2Sk/TYbcl9AE2d32OEX2imBqQAmlCqWp3HjlDWHUKRfhQO5+B/
VqyvoBlr49vRsNdhSI8F9cgnpl7JiUQnyXB6hyYg9N66UZxheXuoC3uHpNCtQFpS
ga6VtWR2EKe4OSNlkgh9u3LihwIH8JekvgaLtvi1thpKpLGtnOZ7rjxyJ0nVr1hx
5oinWbrANVM2fichNcmmdh9HDxY+q7n4P/w6hMgqINAO0wPzgdWkFLKa/v2daxcO
2h0mfohzHpR2RqsGbpXjSqbEozShWTUZ0r3YklMrHU4QxKe9G/kuQwPgIKnz0Jp1
STI2mwVNZtCoexTvk4/v2aZ8uiykcHG3+CHBl5yrKqYwehGIdF+plogYMzLF63Nq
kqcIa4xK8+55o1LawbJui6lNUrwZ4P9eIFZfQkRjZuSlQCfjMRWlpPL+FxOLqMjK
6w9RknMEKXHiNcZf0kC4ddgGbRNboj1+8CSNb2wFdxadM4flPVJNx9D0eWggBKQV
2ILRnkaanxUh3UaXGET9r9VryoJGrnmyIy2ToVIRsyixrgV9ewoJraawGHl2AVAb
Swyt3Sg2MqpiZFinuEz9R8vWETkOdracPXqEU3SVilH/1IgI1YhFozJ0jfwUwEHX
G0decwimJBxtgmZm/tO1xK8lm2JJFRNeAyd7/bSJ8R+f+3VKkxkp/nvOmGFWx591
m2OUoqNvx0/ziHh4AW0wSVTbjVEMIe23+T8cOg60tB3GMUuhRiK1T3zyQOEXAgFe
G6fBTUm7QY1Qk+N8fgCZeAS4jW90aG82wC9GcJicTuf8WCx5EwmfVpfO/Jfk1XzK
QvfG0aGDAkTZJijy3SNscXcqsgWetQuk8qZdeZI3hdGnby1VdyRGEDMGVBtVgKjd
8DqpvglW1hRqnG8wDUXfvGQI7zMimiW6rzSbtGtmT8/A8HqSiIil13/esR0DKPPE
jxA6u2XaLd/WCV84JFgtztVnSR8ATzzIBbkgJPBKUtZTBnY5znxsNsWcbAFMFf64
b/DQU7Ywfy0y/itLvezzqTjMSNz5ZFi6Osi1wwjFvLqXs9lAvfMLWepwgwPrEM0v
MkbiiTtR7U+3FbRygghOD+3h3ySbDVR8WEe4n/pwAjQYlrr3Rq0JoWb+d27Zwx7s
7zrIHmNg7B8s/7g3NevigbBR5qd+5sMKiP6jCLkIMoEVRF3vZMAiObYd+rL/yhAU
y6fuWXJZfsa5NSWJCPOEcRxcwZdtNTXaF+wmJONJnjezITnYvqbRyDCCJlWcetsX
Ki4v8FZ8hxwmU5T53QYNCGrX+ytieHEwLyEXO8RMNlwx6PA8ZEGA5YeHZjJE+78W
ERba1DO5BE9iilqvoUYzeSmvnDyuPNwhZkzt9fg1UUlE9yHvVlh63V9M8lpS+JJd
1jBjkMzHRrMSknkW3sCPL1XUWp+dLwC/GGocoU/Bcg1b8dirhiOInhtzqjDqkxGs
fynsernTXZg154bkAV5LI5gJytUDAGD43f5Ymna7tLSyBAuG5RVujjqr+fbFH1j2
pAh3QS44SjRQzhVH3EGnJXoWhXe+Q3XHZPY1frSAVE5liDxhtJtw/QrT8zkCUaCg
qKuUjhyDwuv7tayxlJpl7MMfVmwYhT2vH1wihyMXIEtikyP6+GfFBrjtC3/Plu/x
Fq9EHCD/rM4ccIx7annJh0O/RTJxvqFWvPj6aqz9kUT7CEH3JXWEsADQDOVO9O2o
yWyLEAibwR/XUn1r94LqlWkxBJeQ2dLOyLB38ogc7Uel9dKKR6PAYGdDNMW5q/lZ
m4+tSJjWQsVBuVOWDUkY7PPspfV94MGUn6CIgzG8zl1RFibLb1IUAbsIYHJ8Tw1/
clrXflir/ZT35PEBQLHBXnLpQ+fyhwv2f0RSgguKVrwpXNSklCx7AXEz32qH6zgu
Hd5ecMKDDyLoYQBXs1GFZKcQLWNtXPCTPmxGttZcQimgLooiu8FqGlNOyOP3SuMW
jX/TO+1bPDgNZ5IFPw5nzkUVrIG+PGRYVYHHbS5+3HKPmLyvuV0TeMjYfVTYaFL7
l6atCPCqjvxaoh1q6Nt+pfX4wIJ1MgjVJPzQH//5j+ZwKb8SR+W3eRerrgSyC1Lc
bmlJJb531TN4HlmAPOIzT4VDVQtgQxaE/LJiUfGMe+zvPGcOPxwJbp7laItT1yHW
ueSxb1RPx+vZlBjwmjv9FI4BoVpJtpRBVKL4JA67k2lDJrFkvSNPxfanBA32bRio
1q0a8VrslfZNdYZtsBtpHpnTPIFUSgZ9JkeaLdhVCNd/+59zNtru1IksC85d7YBf
zdA+XpBMRTqsEUc3EdNCvzv7W6MSAzACA2Z2S1MPnMQk2vTiT+y88A6oJk3NfFsw
bUV7xSQkqkqOsTt5QnBqqX860RRPLM4eoWjCLKnJblqa4KGSb3wHESN0MUQldwdt
R+zY/uUtlsUGNfS0x+zIUjdoV0HMjTBo+Zd/krmaGcnEX04jpcsAjQj+Pv8ex3ID
MhCsjZvjeFRLmdX9VgURaZZ2YAyHBi+8U3XXffPscAvb1CqADpmY5UM4pe13GeAi
U+ItqWSXAdO9Qxcupe0ZMK+ZaSmf3/H+pEu8aKvls5zG24sOCQpTAy+E72jE38Wo
GNkOk/rSC600gAu7pZCpHkDUtNsWl7H+T9PSOBTvATVEnvrJcpxRF1UmlRoUf76b
H61gCPYpBBkxuk/YyWDG/N3WphmlCDViJUPmXP4HhUH710n/+tKlw95tOFAc6slJ
cOOb8+AfvuMti0qYgK7efA5qr4X8adNqrTXUQ7vEuEetXHanVz61QMniTNcOSWUt
VbsiQaMOPWnGoKlwVN1A6iAdhr2SU4vXa63y7Kv5qFM7ZG/VXKe+98In4wIYBFbL
905F8qhEQ+6nAVIuN8joS1pPtD3EqI4G8IyAZ7qwMNIXqGIC7Tjk+66s8YGiimcT
BtLMJZoZPgjWFzACR5QISIGmawzdXfS99RMKi0H2lPmA7V+WleXvn2Cqfdmw88Ys
9dKz5rSida87sAPKeOG1IrUzldCZf4l/gJzYXrBH2X3Vd12U01MJfHog1TLXdI5B
V6AecLDZYJziI2tzJ3bxy9sVWvcragODmJB95noMbWvfO/pGxq/7XyIt0Xb+Qd9U
RAjqrsCZujFsL6fNRn0YVX+HFSOETiLScoc/jcqjR1b/hEwjc9c8Lkm1m7+j+fo2
9Yw8fU49QB5uJBG8UuYVePPFAzL8Lthy2LDGVg84QmzB2KLQdstIcG2V7ePqoAQo
dXIenpkvbXvYiyTwhGZCgSjrdXAkViTEq3MTK6VcDubmOJVjafn6CTJTEtram5AZ
sVy/ONR8v6ReyOlFy4ElsmwoVDYMDy2eKIQoaWC8IKkzMuxZZ8YVUtDogu/mDPJt
gbffELVISPxwuEcPYAEVi0rcPyD5Nn5gXs64T2qZOPQFxsRSnEsb4N69ulvquTGB
bYBUrFk1ldm0HFU/3M6Q/A0ikSNiOqNDoGg/e58YbJW9HD1L4Bg9Zp9GIQAt9qN6
r/GqVSYUkWuSP4Dxu/nW6JmAyYDz094CudGUU5DSmbvXVSUg40XvJhEtTD9oSFA6
d4gZAk25xd7wJZIrLmgocMGXYhAU48tbZsEWsh34A3cLhugal+Si64c+Rh5bAGgO
3QT5qD/H1gncXWU8pgBFD7gpWKNU8/LBTbPiy1KIFsDYj1p+eO4Gshq9macpK7mq
qGLE375s+S5LOGX2apJeiIZQ3gV86HOnwlto9DVHn0YnUWzXgTtANvGvOWhw0nkU
s40v2IiwICOc3EAVtwPCzKXtpGCSxeLEZrrjb3iLyaR3aqItyCzOJezsXmToVQGP
oaE1uMC76l96XW5eBKmy2HLZBxwfapnrB5uCG/rRt5CuHHk01bbXJIeIzNcJSUA5
dbRW46/41sBQs9/WrMwAAEWMEhn0BQ9p0k6kDT6/3+ndX6dSOtNlHj7tFxaT9X2Z
polWoi9/B148/tEptBFYNgJDkXnwa3NDxuoYcGQ846Aft++VD7gxciceAtF1O1L6
T8LKElLLAX04AD2oDTZAUXHJcnKLWUXVZj4CCbQHcLiQv2ZrbCpqnRsob+gxnKjb
UqKxaGBaLi67MRVRWjuZKiJXnrsp64TIaX5QxqMNSgT5ol+t6kvpuEL/d3yq78wv
wDoqDYysD5KCv64FaSv4Akdx2gMNLDJEnm0xNy2Cgu7rhUaokL/1tydBrZUFTYWy
TkTXvWmT5bcv1WPWKZcWGC5fGdMrlwrbcKc91L4Zx0kNuKVLR0CXdang3aL9TZKb
TzH7KRk4xanLVWd5CbtiJGSBVGjt5ewUBnLqxt5ONIy3HpNOt9jxcShAIVh8pKNB
nXkSI1qr6tT91IVhO1zRKBjU0OXs5kKnFeSQxQXtxEHCmnY5tXEnoVX/Nu49Gzyl
9XM40ytc7VvX+A3X+vmro0jIvfEA7kQZkNSx9Hs0vvCralbItNKph7o74CE3x07w
7PS9piVVQtMLd6i1uzDlYsIUzcqa5QEeZOY5P+bRDeL0iWZIX2f7w6yYaMkwGSyf
qQG8QSssOFD/OgTos1A38m/SNUBjJPKgBg5cyAcOcVaXpfG/9TaCzU+K+tPUfqSp
CqmdAM424Fdvr2pGZdDOZ0m/iHV/lEJvBe1sXk0/an/1Vsc4VTu7nHpfE1ChMx+y
jyXEM3hcRNmTDCz3cQEtD5XBRF3yjb+PC5UKWF+moPkVpaEMyL8qMgAxuIvq7XT6
9Kmva3katpcNa+W74GcbwzD4Hf2gGQDypUwWq+MT/y8AM0wnk0Obdv+sLeF6hLLn
rMX928hEvgrG5N4HWTKRxam3NUvY4mRdj4oDDn8aaU+hkV3andUzZXqFNWY83SOU
9oXYx4TnOHUOJXSOB4w65nB/GNXd0UPIVccfmKk8GXLa0vr+eI060vIkvknlP+Mc
OEWYieyMOKOSsbPdnR4pBjeaMKwGK0m55/kSGwuDJwpOVrzjiyv/TSFo6gR6YqlA
wDZADM8CQ2agDoCBT/7ezfr+7iY6Qxe3Qme8MVaJr82AqGlabiZm6YRusxKU60j0
Yo3lyWbS757bvPIIzljE9XpymzRHPYTZInCIbC1tPMh71VXWZlsEaaCyn1BHwSYA
JKYAP2eO9MY5Yx/ltW3a8C6i/UbmjH/GdEkqho1GAkTes3U6TkftAWwkayjNwShv
9yjVAK49RT/NMm5p/mrdd3I8ODch+kCQJiJwozgGWDDNawoFA2FATBIOrEmw9Ban
0plyzFAMCNg+fCV2WWif2DWmME+qrJebfR5xhqyHo2Ccn4nY1y8lUDzmLNONOxGA
v/hhEjjWa87z5b1VEg6pFFc1BKvhxpyDa/n/7H1ArZ0j3shf2Qspcjlt/QYYkyJc
aHhMxhAV34TWPB02QaaMbwzahoZf03+oeeTWVp8ePqPzoE2tWzuM0X6aE1ydbmaw
NLUngCQvjUVGUcWRMCCeQiBKtHOHbM0P+igwWX2kJSjO0FNYMCHRL3zNtRRGCsE8
6QgEfTxDPdhLk2MaNUohfYjg0wuCAJv6WIsPcizgu4P0gT3a9EEXytELkGVDHNPx
hGDgTmkWMQS96vcJ1CaT+8Sj/7ieLzfZcNdPQf80/3Ttegs1PB65BJnrYhqYU477
AVg/sctisPGe8OGW/bVolpCBJorpOq6gY4c4egpIeAFikTF0O514iWcioioHLP+U
HSP6gF55P64wItK1KWlKixj3/yQGwL3kE4RCXMVlHdvccncJk6r5BCItE40KJrRJ
CkLJokm++zKjywDybDskNC/qCTCnh1k3PBQJ0JkHb5ObWovju5DMfdOBArt9f1Hq
gYirEAI6WVaYgJwM+XgQdGvkpnCvCGnPC1IK5Mjsog+n23R452E+d0NfUu+fA0v6
xc+UQ6VDhID8uS9pQV3Xqdq05T3zqUtHAwk1wg+vNBhj5WE0Q/QF9YRLmtWCzz8K
h5Bijm32ISgQnHMxEeX2G3xZHK/40Ye+Y/4oTTyygVEqA1K0aKx+qYjC/OpCoily
/lELwa59d7EoK7qr3Vxf5MqLVMv4eBWOG+V2IjZ+IBzIJx5fhrm6lwYsZniPbgfS
HVfniwkkm7oqoBXATFyyJhi3hE3RTF77DL9eNlo6oCczrwuaZMzo1YShw7rlp5wZ
eMaz/wa1Fbm4iqN628OV0KpJp7OoUn5hm3V6ElyL3wy56odXAVP2ziAWytn0qUeC
bS/pg9YoWceApnXDo/Er3NyHpjKn9znJ9g5klvfeR/30PqR23x3K5dHXMklVB+1y
t0AG4zWSm9r6V/gAM/gYOQBM9hh5rK731aPVpUFrz7+VbLk1gfB7xBtg7Go/4IKF
HR/oCYyEGpg+b2aDTG+ZyJPSbitenCduA3emKlvztYhZBvyeKAcRJKwq90m3bSjR
rOqhcw1H9w7VYQnrg7reUZe0cax2UBqec5bm6sPKzjNgwa3LNJ5hn+gRotPdESoF
tc1bLvsT1D9Jl/WzBJ4yasi0aQjx+Y2i7bjw1snGNZtmkXHAOQF3GaF5oYN2HY2V
WoRm+Z+VSy16TJ4lZmt8PF/WHErF7mrPX1gfyeNEAYL5qyyso5k3HNaK/qKFDol3
YzOQ9nm7nMNingbRQtM2XUfNQvTLxgCFb1lpL3F00n4TuEGc8pAXyiSRqx1qtV7H
JOsz9Fm6BUkqVFCFxheXzIJulEOW6fT8H2xIc1Jfm27H2GOO3HgXwtJck52g9oBh
MyIa+7w7zU+hu7pOIxEaIkWqVI44Y6cOGud3Bgimm/MtRVJ0K/hywi68Dm8aoQwH
K2+TW6uF7ELCOtjldDxUy1wKeJuvs+v+/UU67QAzUdEXxx2Utt5WDQLVk1yI7Fj6
0yWX/taqz1aVNGFX32w+srpD9BLs/UNnvLGWcK/e80l2/5Tx2csEnBoIK7u2UD6y
AbMcngfilDx0xkjMma4eSCuosu8TxAJfQFCX4IkWCcEx76Z4eCB89uKtLEL+ne6J
QUlOi/Gscp5YfIuGkW7LoHGK9k4KE1um/PDXDgX7oU9tN9CQ7JIjex+A5XEhA6no
Z6vxEsMqRBxZ/MjyxUmMJi4aH70f69vuq7tr0DMC4THNZZum7w2FKn3jVz03Q4zJ
oxBBoVGGwMsIiy0oTgKpBs1MBj47x06KRaa4KteNktat3YsPfDElf3x2JF2V2Xnq
2uH9M68NaE4iaimlCJdewl5MPabfNh77DmJxRpxLbWfTNEUjEWkd52eqk0QQw2+0
QzpmZADg8lNqr3XBp2DdtRgrNTyoCuPsCQ+6EOtiMWsahKzluoM177rdJAbBjw36
vLz380QCNbMiDxEiQ0LWI/DT0B7+qsSEPo4XVlI30NUghEDVzGb7N/AxKmc6ZHFU
WfRu/mBp5f1IwlgTPoj95NulklWFrwruepmIdfqaNeFOcF2bF616ds9rof2bsLpi
MQtcnA7exlWtOho3ZxtnoXTU+MQgI8eX7WX0LYK2+GHFRHEOKy5C8j9ddrM34O2y
3x5G2dBtyDCbVLIz0MgJYgI/YxyOxLdlEB0/N27EU4dgBv4GM7BN+Ny4hL8NrOb/
SXu87o4LnRWtA6SGm6DGDCHya2cLMuYCPGsNgQnhizqg1VEDeD9cYo7YMex209yN
TJEyKwDEmyltKkSoYLKN9YE0/lFYuTUpytW6XGwYSsjyMa4KYDr/3n+Fq2EQOda0
bsaAkbB5cJr7GyTCcrTCcF+3FRLDuty6v2nkeozZPRjy1aLk8EE0uLLA39X5oFK9
0YTXozsOBsLfibek/FmGSjenYPo0x+OoGvP8dQwqNcn+ltIOTb69QhWIw0C6EuwZ
LMCxy4klDVnniOtqr79lx6r97zEjgPY91lolO+SRjFn7XC9Qx61CYSjzAbejZ0u0
y1JpZ6nXAnuMbltR7FncdE7+Jj44dZWy85rGDSi99aRUWsb+ZUIQDyx79wKJwlSH
Cb6xWrcUWzJ+DfnqIsW5cMVmMraqPPQGGk3xxY1Jff3OSvJfqrfBtWX7nWdzX5hn
kGheOpEqzXTOw43iRPRjilK58avrwBAMXPm/9e9KrjRc9Fd83fnNO9WTn6fUM+zQ
v5DqD+Mx0iQZmyWACnRCspc9pSkSU6/mk/E3sTqgAtVR4P6b2YmVpF5N2LASPK35
pJgCKdHkDqAMhviJyQN1am/hJ9sE+kZ1SOIrmV8wxTTu8w1IZIy3oEpphcuD3MyK
oB6HoXB4tDLe43bbqRT3CXhvTE+9vAp+wfBHEt4CrsEq1NN615DdFJPXsXwkHdTD
K1wkd6t5/g0pCu08tQFTyEfr47IwIJCRDoGGj7HDLPKxV3O90R+KbPBwMyUqTDHq
juR/0MI2emK1w6zAvJCFOJVH08//zegZ+4w6xMz7yyPOC3ugBqMkmQaQ/wnAc+K+
FxzTrjsmujoGWg8noqAHrCbKO3yBDrkht0YOeTIMxfyE/fMNpVGj2w5FGkTV3/YU
/b/bVOlF7j6f9+RjiWSu46tBRF48HDP2kqw8rai5TK48qQfmnjnSxyHnUp2jjXfv
IwcmxxjyEVwLoTLVdrt3cqj/6O2C8XIJ8x7yUnL0iomL8MSfqiaiI1JHdwV1dFVE
fpDexS+tndm8a79/Fz4UXuX7QcDZefSOGkoDcFpOH6ZPOwJVRI2lbELTvix5SMS7
VEqM+py1LJITXMxlTEbNfzoUCo7LsMseDtgLtMbnPzdO+OhrLBkf83hdnzri/HHp
Q0POw1e4bli6TgWBOhnF2gOoF2T0PiQVrI+OfEcqEydY5VUgX8bItgXOyZUS0U6P
DWq6M9TA9saPcUoTfyqxiJ1jlcYOVbKmc7Ki9fg4hNx5tmxUhge1EbMWyLMZDVDl
aZxMAIh4NI/n83vWmw3B7bNlaby/DK3zAYmvi8CQTZ4IfhB7hUdqJ8jm0HpW7bqm
l9ZLcgMIp/xJM2DYYcGJHiyE14f73jmCpB3vkSxIGdd5mJPN0ibRoIaYACN7EwC7
ZUpzh03J27E1ENduEak0iKzW+YB3SsyljMkZ49rUcA7MCWta4pazl2H/C2Lb5310
zOePuoM5Vm7KKB9g7VOooBoZPwyCdDFF1ELkOKO0h1H94s0iBOSXmH7UidGT9lxB
JooRs7DEUR+kRCCOGk05oVnVl9T0I8zrflMyJ3AI0wGlzk9347RRgrxEveVgo5aQ
nqNepxKOXdEhgTdwqPkbVPWtBuGvwhaBPj2/rDd00arjZJ2KGK7ILMAhcP+MrQPl
av9V7dFbRD9xNG8FAZvb2wHg5m082gx9I/nqhwkYLFdhHZdt0IrFYJX2JM614A3W
m5n3aCpPCHn7GFw41g81zuIxZq6JGPWA1WbRj+ZvxCk1dfw8R0ZaZyYiPS8J0GYT
jcORcSz6Sjx1b2WVUTyNhc6WOJen4PTb9s9CSVHpAcpAYgHCTaWGJPJKquOhqRAl
sz2j290zA7FKDowOxvS8YuslA+90lkArQj9EYapQXTIk0FwS4wpsodXadrV0rr0y
uuNZEPVTb33nWeU1hxcYMhY859Y/OGVOESSmczfZ7iXbahpWdrXuPhw61xf9cVkT
LsY555iLZAiUioASbxpcXFMzchzWsi3snhJ9+UO8po2qYtPY9poVUiY9BCjioeGx
d/KU4ifuXt4RBly3qMXPy7kOT5H+o9osImJOBSlhqGmnD6+Bm3sRvvN0bkTNBk9h
6BjvK8kdaYvqHk/o7G1lES45KDE2qdXyu2LXyZoJuoPFFwbfeZDm/CDKcl75VtzR
QTUvCR+rnLF+f3fKUyAuNdNUrE3VzfkvYV7zZsog4Tu8iSatBLTgvhJajCpTukR2
PZP6ztSRvbIGWPFEdNokZTtia7tcJq7bMJDglNJbzs7MOuZO1fe6QoaeyImv0NcG
Q1N9+UmTTSLxXufz1Bkcbv0She0mCs+F/DVdGvdxRZAD9rhbJC2s9ToG1xdKDdlF
Bqlj/PQ/uPFjqtp19P9Km1sdc9g452vA8SRfRo2syc0Z0hQJOyVJ7sN1a446HNyX
X1hQOOgFpN4XBAOk6XPJ9I4XYEElMhJMjbh6QNFVrk7R/HV0HMmiCZhdK8mUhrhI
REyuXBTQ7H6aMASBtpJMTi43qnTjkKAKAqGpeACTpGkYT5GHFiZ0WbcZyP7QpT4Z
5C24mOAo2l4VqZRLOkT3gXu5uzi7wVTNA8/AvosNwSsprqBVLPA18oKYRqKjxtFI
m2pddXEab/6suASK+5stxUiWXRWz9oC3t6XjXbvBZR4nTFtCPCdCp8pkO7+C2bve
dZuPCym+qFtxgALdAnFZ64xmzqOHJnu82QAZG6hG74DxMOdyrzkfHY6RxY7ru9N9
JkqxXaeUIwx6tJ/hKDx6M3pOfkd33uAX9ZzLNkKfC5MsF7DNzCAFjb7efj4CFsN2
7LJRiScurMQ4BDI/hB2rBrZ/R5mlAR/3wUsHnZmgycfiqBpm+arRHh8AeJUdSQCw
teZLu6gX+4tyCRcGaOAQdT/3JJ7NQTV+/CzgZrVVe25FIyR8N11vVLEd9EsM7Q8C
7rPrdiDqhXa36sGGhPATEqjtSbICl9rWvG0ZLF3wSiduEQHckdsIhUdGeaO1jm2d
O/+1fzKtu/oFPvCSgyrin2A1ptGIHze4832DDP79OtYsgq/ICK2S+HnQ9Nk1ciVZ
ALJgxXmKSW+ES8cY+JHuyy0Y40b7EO8loD0WMYSnT0F3lBRe5oe9Ap+JTd9cx1XI
imsRMV5wi8wCzUKGKlREPjeWCeobSInEuJ9xtpWaiTr/bIzS9+/q/wF7qJo9DAkz
z0JBBQTULEEZjzVNwQMWPyx+11uco2QX/rAfqbrOL/1Mm+Iu+1v78mKosJjy+9RL
muGzfXTpabPqOcF5jZ/W1tSAXADWTZZetSgb+d212wbXLOBfc434G9cbibAhPfUI
PFzlQx1gaWZyjg/YLD18kLmsR9tcMTymnfMa/y5tb9RQApg8lRgwLYyzYPWm1XYC
+rsPWNNryH+EbWqjzou9fhamIZtWi3UWzmX2Fs/i+YIO7BtRe09y5fO3s83wADF1
N0kreQmrmin0aOggzpFUo/W3NX7sTgCt6Qd9y9G9uA31uV4GzEABif7hRBH5f107
etNZYdCRQpU/48Ge9E4Rghy4lShY+ibyhld+fIIPFcsNEosNs0LaAQoOwmW8ZB0V
rzabJNZJV2Mletif1KkGRHbLFnh4fSIDCJGi2BjaqeQ21OiDcpAW5s5nrUNaSgdv
p7D5BfTc36tDC0Eae9pESmY4LqB3ppMl1F2/N3VQg9U9QaNzKdQWawlmQHPJEg0v
j5iSJO6U7m5t36R9Vr9pNfYvaEg6NPMpBC7HdCAh4lR4A3M9lemb8wZTe79SjupY
iIMNCyUu9hyOgUUysx9HalVgJAVbGu2+UnohAMjgk5dMWzTIiTCVDm0+8Kg4k/xn
mq7ydK+3TyKEhT5Yy8VpmjGKQLf2ZGZZKC5Fc2OTOJjPoZKxrWzybycMp11yPbBb
H6ZdR4lPn1nfdFdfrMYEX6rRWXQSDPlRP7htiFnCYJpyhuRwlPNxSUz0Nxnio/UL
IBlHUUqozGEjRpFL+B+XtMuF9YpHgOAUWQQ7qORrFmBnP6X3iYlLN1NZa1ohPZbA
TTuYKrmxCKOEfBEOlGenMsbUX8Qt+oxbd1AOmGs+1areMC0rPh5HlM3HKHKm4Tyh
EnWypbgg8tGB3Gou+wCQhUxvhSn/XWDNN5mqDtN4tpvouXZ0qGBt5V+4fWXS3AlQ
QuWWuedaGh/s3YT/Wvda4Zi49OX5/gELg+b3bVVIUQ5k7SNDv6dPP14N4Pkkvnii
F963X6hEN375otLgpZP7XQ64fp+mkPUfhPruCQr8J+mtdVUXS7NuCsAgKGT8eLY6
efqPw6x7jGmjfY92tBsQr1NxaUIAPSz1L07Kwp+5bhm9i3Z+Ue0hQZ3akJodxrX3
M6UanrOyqGVw8t41nhsc2r4O95rXZPb3Ih35qM/P/wtatsAGNCz94ryvjG4Z7K+F
0YY4BJHmyDQu3ihw2yLBIdpRcE5wYjVhrmEMhV1TSVmK862IqDOhpt7UZCoFVPKd
f/zM0luvLc4uxedzq72O1Hd5C3fk51L3ZPTzlOz7JHV/96V5ZtyJigOWX2PLKcQU
t/Ak35GOhwMrBgn2fOSH5HETe0m2XdoiWdVhiE/9R4PbN1LWIP4jcbcO6xvuU0T3
lWhp3aJoQXoqQSxjkCLMLqjcE/IXilgZzx1LZj4g9WbIM9i29Mbd26zdcDHkvopd
0psZydHl9r+UFAOrGPiAYVZIQuKuRXgBNaaYyu5OEYdT14BrWPNhpNf9qxsvRFF6
3+d1+wy6LD5Zw2G8InCp6wcQQWcQlH9rHEMhY9HZsYTDI0wmMgpXNpzgXrkDrtC8
I6oWn8BlyrQtGtpwde+cJZB2BhbLeQlMdlrO5huBGEWmctBFFgxcydHPNoFjgIz8
GwUQ4kG36G33/yVkL05jq/UWSDVYq/zJ/+yUpEEPP3105Mdn3ugJ1rlOeQt6Wz2V
uM95K7/SnM5Fonun2PbCQ5GyuJAP4eKyZ8Wn4Xx3OgZfga/fi2lwgAuxKnVX1uv4
L57EPtcpn6DiQ+/XeCfS3A9ylUpqVJZa+HOeHESovMrSRUTtVZv+V0u8z4/Yg6v9
Wik9KzCarrxWnQ54ZJejuz84mU7Da5bUdLl0bLsxjrWBxWjLBK1JOLe5p/AYuHVI
aiwZz7ymcoX6UM+c2AUXwNOJySrztGSP0mMWXpBOwmAEA/CLtmqCdsyE8QjfdDPC
y6MAinIEe+B2ZAlMax4eBDFqCUUfCs9wsrzIqso9az0VnegmxtlbIt++ms08+T7U
vNabtPhoOq87PcWUy1LY9b0UfIg+lWH5YF+dq9IqmR5JLdPpd1v6Jlq0SM6n8/wt
XK5nsZfz3JEqTdYPOEQdtH2epLaHWK3dFWQgaIUscTZ64eRKFM/dZ5X93Mye0QQJ
JoqhH9s5qADz5hiXm+WROhM+jYBLfi23V2eWxzfIG215r0AmV79BJtD9oq0GhqDJ
y7t3gmLymqKSfHjEgS8w/eFL5CuEoi3HVGgIjbX7Eq1b3IX/cqnKnCpS/zshhxya
NNuwMn0C3/gM81wzbxdsK1YJp8CzBBysOUjNPIWKpgLfaaPE0Y6rfprX3LlzpG2F
+vf10N5Ij7zqdt13ARpwfjRqycu/uxF/1q51yjOnDvRQlIAZYsc9rEoOBx5/AAO5
50YuUKyB4eVq6Bb5qxRWv+mhX0ZDWqyZGgLOM//zH6aWH5rPRqw9TwEPuXlEloeN
DR55NbaSAHXe8UrcIJaD2aLypwdpBJGd2Stq+mbt0et0Ff6ntMG0g7sIdG1EdBBj
pB9WCz77hdoegeN7WJHSor2Ovw3Ot1hHQoujhZBXHvjLcNXx0Nu7zQhajTo9HF3q
MJlbn4y94uvQ1TXg4C9RiWObbjEFHKIZqGTST/BJB0rNkWL7ZPqH0fuAFgAX8jfB
lJ+sPeWQoIY8ySOhFCskC6RFkWNwtA1oPiI6+oN4LWVJStsl1QsrovJUiodQ9lIj
nbg9zm3aKLbC+rpX+x3Ra3j0O35d+ZtgXFlb9NcQ+kWxFSqODeGhIxWIDDIJdAtE
/p6bvwCrFIfh/Hga6Vw77K8skddi5+WlxwGT8F/Vhjr1+o0bC4gA+RmRxAYyZb/Y
/OHIyhNbGtpmD4kUtVq2tJpZt9XVWmaPbU24XkENBUa7fG/cn4Rr5wVYIwxJ1VnQ
I9tL1mYiWljTz+/IclBVdPyPYBx0eApgy8UWxfUeCnnUt5kn2a5p0EPC1gXVs5if
puu7AUoujCXBq59IinIeXg8BbDe6U+yRu5wNoi0eZBd7QZ8UUyHAlt30pMWAy/Ox
eXLSaIQ0yoKgZ11wWPShuBnyFvZJEimp3l4DWI1TyloE7yeiOcQzAu/eRNayH+28
DVuXk362MMgFdH8rR25SfP4UXTfjOGOe2GmnpMJLD2Vf0Ie44aWOJXEw1IihRt2e
B0lCaahnRfZIBe0hUAT5wBOVGE4TFScOOHx5yOYINpYjYtScsoHY55OBh15/5YQH
yEVbADu6g809RnYUUH8dAaG/czFMKrSUa9R2K6R4y2tJmhKq5cIssZXiz1SrhnZx
9aZhfiPIhwoMwtY8tU2IeiuFyP1e3Wl0x5UkKTh2cHTQmEIoGEt2HsmFXouUgU6m
OPRrqXcaztiuG7XpZikovw904BLKpvf96MrIAJ2Rff+8WdeV/W1XjD66R3tuwIUA
5G7WRvXjqlR/OtaDWLuLHDOBDdDMo0mEEWw/hXZl94yjlCbY6x3+MV0TfcojsZ2D
/hjq5lasNleGX4rve0OlTbDvKEha/GBWG07SAtnS1HzlnMhvqb3KyEukcJXnA1rT
kpX5UbIC3rbyCnOzd44pYT9zjN6fU6GE1HdupZNRsCytfG3SlQR4Wh4ejD+xEcXr
MV/6ICXUNXur6GE3HjEhtLAklsj+/XxQLGLB5i0spavGw1MaHeu0mJraBJG2GV8C
5F0zDwKlGos0EDBU6hgDrDmqo49eXbhyFAwhYzBef6EjdaZhxRKbWgUI14juJB0c
l22X3KPL9L3Hm/7rn8F5MdJOQb3K0abRsAC29hfMs/nf++uWwaWOhMOAkKmyPxe2
T/zx33D7ZElrQ3/9ra7HkMMWb5NKdz0QfXysKRqd8dn24q5t5k2tTs7a4dyoRPsc
eRlxPiZXO5SIovCrxed2qNT4V0NSNJsYowCitmzYbqSIH0tVLX1hojrEanQ/CKKw
QweU7Ww0kZy1+KqHJK1caHeZUSwDmy9WfR5XOGto4I6rNjE6/K17XTuyxkwm6y1A
jWED8CQelY8ZCMRxC0kfBN27mSjyzNjm51kVAwKGE8MlfVRz3K09txtghDgXcNFC
vu9K/0UHqLYxmbCkmEe+71BlSNhSJ/IxviplSMtVk3UNXjEgpyKs1zjlk6SliZj1
eOGRHJtyRhKM+CQssdUrwT3HKRDUEnzwK3vDzCDuee1tQfr3A95cuuhJwfelTIu9
wFDayvdba/j17BRdKUePz3C0ueVObCsAIxwu4wWfmaVKYBVkIv7pfS+8HnwxfGRX
M3yiM56BF9cr09sAGgVMe1/30v1fDza2bg3YA2kn00I/X0FEVMKnpl1lJiXiNg/E
hwydYKsCfhJC7Zn9XfMO8Qf8/QU1V3/J1KdNqGziKSZYanqRg/cShBzVpJqTVGRd
0eatK1dYRHQ0QYVeKWIRvmLRCq79Du1V1a1EcaSXTCeqX/grQIwjLXGuadn7p77m
hig8YHc6tudReguMXVPMqOPsVJLYYmBzhxT3LVSYaPQWdw+DPj6IbZg+fp6ApgAd
dlGivIVbH2a4W5gwIZHMP20+YSd6P62ESSn/kpDno+HXsJazNPGf4a0n0WzRI9V9
oJwTjMZ6OE1hA/UUccJIE+2SwYMue13KbOiahusPQf7Eg6SpeYS1QYPGWdHlWcqv
Sxw2MI9tAM42T5JFEUPPjKA7KGX57Wr/8uqLnKKlUFZ/J7tdJGLlwmlnafIPmhei
CQf1PjHm7M+X4j1qWTxlRkdMc6qaziRQGjV++i+HRTwWZb9P1jIE1QL3/ozZYxHr
0PGbyF0bcWArpRS1qV2w6V5pXMg/HcIRGpW7vIqWObZrSEjkJ/Yybi/E++bMHo+n
Vr5j8Xe3cKt0EiYFOYVeJYx3Vth8WgXoPD5Eue3Y0B16Kuit0vSDb9ZxbZxMhGPV
41hC8RBQN6OUhdcISeH+Tl/xtXPBAm51cIcXnKhRlza9vpmFU7n5C2MX1XixzbQq
6L61S2XINSmI852lRlhnn9s57Gng9t7/CHVliD2QWVZbRT4xgPSxtc70XwS2uCc2
HidNeU3OQBoOscXmx7qGMRonJ9S5SeIb4ombMaX6s/9Vz5BuMlstN9n8PwbTu70N
/h2x8TWa3JCPNY3+x7Ak3pe+2zpVaeu/KD79SP3wEXrtWsB2ee94vMKj3Xe0yEeu
vRk367vsc94hYD8wTcjcSrz3B+pEVtcNLsDM3wxREk5DTbZWCiewZ8DqiL3EavxH
mFPgTVGu2Dn0+IofHDW8OMzUFDhacaNmsW6Z36+YFTLXx/GkTiCsU5/XsDXJhYOe
1i/6vVgppMROKL0H3+afUJvpIgQCrrbRjXBNCVN2ZcM/MaGIqEPEve1WcaOBlJA4
b7l8Jd2u0utiSQ4MeTxnVYxoujaMQAWPXenxk93f/OtrcmziiVHuNtFUaY0UnhK8
O9cZKkwvSNG/nmogcSA0CgCZerz2ml21NXPn9t7sy9ShU2F1pY+KJYkVRfgMNVMj
Q/CmTTYRzJ+w6xpS4/rd+blHOJhciGPJj4QFESqQL3nRz+A6xlSbGetns11ExjLm
RBm0wNBZ6P/KqinnYSHrFW3P9sKlj2+OE8chtH7pLgFfnjnIwp3UcRDFL0Q/wWrk
BbBNnwC4B32TbGc8oS6S0/OiiEeNs3gb1oCZLnWkHCTLVfWJ2121/EBoOOicu/9V
HmywdVbtUI2ApodD6Oj7fbtQnUpHVJITkSkYUQVz6QXeKl5o699nAIW3oXlR2tqt
RnjhEvXZh0HZ19FVRL9ZdhS9hy6PcsW+fPt+4Is54b9L+eoqCG9Pg9CEWGYQPC7X
4b3IJUKpWnmTSivFbE4nOnni7tb0Q0GlkBp7YU1FkGtev89hwkPopFyflxwmhc1j
q+ax+T7q1shOb8Yhsxz4OOspMBJa2PspeGCbMjx1Q7mTMLJ67iksEdWlGfx+Sffe
N1BLAjUp7Xb+I11VK3PGsFpAC/hlssMTYK84yoUQW/uAFv7SzqRj6+svwuSYJ/pP
Iu4ZfA3umbUFqzhayE2HxwbgTCDw1X1X2gVknf0QejohKelVmvuESOcjIIR35w7y
VVnkkDSbqCiBb34xGrnqghK2ubuhajqUAZ8czmrXWPTX1QBy9/CJEC23eVEBdf2Q
W8AOM1ySjWEnps959j4ecYfuKslP9Y6O9Shak20jmXei0wjBo8opNhr1Z/T/vUVT
v8s9jwaztzSUb4wMaIJq2kT0o4SbVudkeRESjAyT428KjdoKX6bNyEUfwntAbCdD
QGt0VTYZTg6ctG3IOL9+mjPHo0UN/fDQuiRA36k9mP0FQSJSU7t0GtrlQFxfVHQ7
E1rr10u8ZVee1tW1EMivWBvMLwmoYkRiKFR9hc62X/ZF9OPcxf78W6v7BTDBZVgP
q48NeltBmNwTsU2pus1Z9EmVSUPmiJFnp33mm1Tj2tiIonIbOOThm34sA6wLwuvO
NTPN1R9SbYar4V54mJKMrhsBLpGvd/mM6FuQ+L7Yh8+tSh6xcwlpuwkaBAapGtvs
2LaDGJcS0s0iyu7yUcv7g9CBL3jvPd0/6EggoEeP1OT2Fq2xI1pv5jI65dfVLE89
DI9biR8Yq+r1ZBVyyk7FfKgLAjZG8AP4zIf6I73kKTcGmIw517cspQwNhAjGyIuW
BFi72jmQGng368gyFBDQi0tTwZ7bJi1VN76tWlp1noVGZ2S9/uaNVm9CT+qvOuu3
P+Fp5D1PXnoA8Q8ok3GuolX8V2ZClo1iPq5s1o6uXZiNTwhoulGLcA+liCjZLnv+
UIvs3ZPfSrInK2N16KfrzxGNOefAI9u5jpvEb+T4aDdliocD+Mlb9NTUQg7BOa/m
4/+6QUcs9sZdAcynQ6+1QRWTbDj2uluOgYtvWKDIiVCwnRK7BBBhHQYedWwFXfoJ
bXBD02nx0kdKN4/J1OswOl8ao81fBTn4EYRAjX2YD3nFLHxBnPlg8iosPy2yy+4e
6dSHGVJzuaJ3OF/wnqV3HJ4zLqbfTLSmaHY8i+fQrWbzs1+zcWSCNrWEFhhBCoNf
f8W+UOIO/Jq8WEgy+gp9u0sVFY7ZIgHH5lrsJLvfRXfg6fILcp2G/w+3HKLpSSzb
dZrpfLki6QxMa3kf25KKipJQ1RefU9RzTDHCGVfmNuXce18U+MPfIwgWO1rKHUj/
PT9R+e+8PzeQgwjqlGgCtF5NmBuA0FXESDgToHbzgL0GC8mWKMQ9oRmh9WAposmA
p/tHeI4ENMTN8SDq2I/KF0ro6uCiJpAnq+zexNUk9pSS4vIh2Pln6eOb9Yjg56fL
SBSeprV/LltX5ScYnzThYAlDhgweoNAEhsWby4ZueMFckG/72+m+sUD71/z9QQPe
2pZ+JhHWNQ0x9f+TEh4DATDfUodfzUeDHI//m+pgxYuDa1LbWvqmPBthBOmm27jD
GZdaIH2oCJ23MPXGouoUtqwsFRjeF4tlT8rMnCyUIuQvJx5xxcG5FKEvaezfq9w7
GIdD7JZrrkFH2NuRjo/HjAGjjEvYz2rRekxunZCiYP+nTD08S9lrCvfA+Sysjbtb
EJyrkJgM3KcuTWKuTZq7sIXbEhH9xuNuPpmFwmPm87Ph/jW0oyDecJb+OTyUMWLj
+2mawtx2X/DyoumVM1vrSBKbtzNEr7IdzVgxu5fFsOGzYn/8uZRSWQz1QNcZc8X7
9S0CiytQnArszhXrTclp/DwhfNkPqWR1nWhH6kQN6/zicJuhoRe6cyuIX9q5a3Mz
VDOANbQLYvmPQiC/Qauf0pN66RZo6TlRcecVyJErv9vjiogR8Z8piXzXfY+93adt
hGO+wXnPHKtQdHq6XYrpB/IZy8lMXkI9nMj57XLZgGbivox2YKsS8DwD1hO31YVM
6CxJkk4DyoOA1RCcFjwY6356F3d0bgLqiWVvSx1sCI24S51nJ7boXu7B4CCe7qk1
hjlytSNyUNq1ocmfV6mcgGrqYSoLfgKZvvQrjKOPTZ8UCO6wAjIvizXUnwkeGTyM
IJFVvZObXM7wyZDI+/msNT0jU7wLtd9eMPDkX2UCWwjDyFD+TxgCXxKV8U7HKSl/
XkF0Fn8v3kjIElQqYhEhNpVNeGLJdnMdlpzZlqsDhrl4wKy2AhO09Xp0n3Fri6dC
8ZQ+oi1kb/oRoEBumh1By9YggmBRyvRcLLlvd/V60enI5cd65RK9VSlPu+7tgN1+
p94nGqnZPpatu/okElzo8xoZCE43Rg4rAvyfGH1BBfdnOFWE1VnkhNwg0jU39Oep
lq2KJd2KOc1XnqkB4MJ7ftUa1qUNoYmCtld0Ur1wmlYG+OmMAvaNRsqhndy1cN5v
xS0FW2QKEiBdF/YRsldcCo7zklw7jn6tzcZ20V17YWn6yBbaCQXJ3l+hAOLq0vKX
TVmnGkLNUUAzYZdeHIliK25FYyXTq7gUiVYQsYjzk01ZC7j3AGdzceFmtrhhXgwo
ZFnbu4FobJcrZcTBnuP1SDILR+ABeUoJiNOeYsTRqLdOor1v+TA0UN+MrfbKe78w
qaS3NcB3O+JVCsS5ArMHwCuZeelz67UT4f27hve30ueallHNxRNg8R190EAnnuNO
Wf/MsbzyQjsDhdwpnwo16jRVTIPg556WVp5iRdScEh24KpRm3M/ki94ll4wggU5d
jVDrJqkNmKPPlNVMXmxRsb1j5M9PlWqeO5QTJXfo6VqyfwxxuMPK3o8wYrvBo50y
8ZO/KA9KNy39j1Bpv5/JEuJoy3vIwUnXR5mTL7+NCMHRB9FLJouy8mOOCgPJCxz3
SW+1nhLEkE2lmIqv7V6Hnm0bctnJPpzwnyKuPg0ZN3qcj+5ZpXh/npr0E2/1iAap
c6nd7IyIg2HttPnbnSR7D6CCuFoUzpirvGzcDmc/6By1cjmFCdU0T77qZC6TEc/s
I84zbbXWyQtvOLpe9ERnyPdLBVHJx0/8FsrCT0tZfqHaFnIrr1aAOL+71aDj/V0H
rM1j02IXGJH3tRmeyvlwQ+TJBV5j1VYaLDekn2xd1ATzJffA/+ccRv3KzLvCpamq
0/1u/afPpfQlI+3CuZDSdk3w8sNx/0xr+r0OU8CFyeHfl5o99Yc1R4uU0Gy/srFX
rTyZ7w6AZeZ3FmBXOUpnF31gH/CAb5xceP27GIo8PaybDu8bf3x90ufWdfYOmfql
iTtGi+yEbTmcTns/m2ZrwQDU9HIGJepskTj5hAm/xKW2HU7LvNPzMiurXa1ycCsQ
BY0Ju9u7Ng5vZH6F7OtwKc77x+04AkF1U0+nCHB9Xpw/yJqy+MmUGyPJ3vqq0zFx
ajagXu6itJDdodfoTQgj316hklLJGlX8zh4wDahOe2C7DQVhIwjUjEeN88qh8v1/
aQY0lGsH+qLfOSG49rJHr7s0IT8qv8ebiUl/QWMZ2wp+4ofQ6en6koBgVmPyUr0i
C0lOYPeKyKj+deynUC27KGWf3N4AUvLze7wyPvHlzcx3KeMDr1ZOnbMddGNT7mV4
pz6NfS9QPY+wSNs7GCgBVq3gYVMpU2sVvJCEYalv1W0qYcznl3uo1PWpD4Hx8WDx
XX/6+AE4Ai9Jg9rsQjiWahzYviqQZmVqtyoNwuCErPoLBuzSHPwQdjIXY4a12WES
NuuxX2hzYWLq/tLp4tmDmQXGZVo6JlHd6Gwwq438vY/JSUJ3V+1QfSN6yxXYOZzg
eTwYbVuT0NgNpExJcEp9/L3Qb2C16psdMrxm4OG10shAcTp+YSOzWA5gEpnb+shV
UtXV9Hsfit5D4AwILs2/P6o13GLqNfIYjrifblHUofkGWFDOBhicLb6J96SfxbrJ
PAgcIyZwwftva3a5b5Hzm4Wl9iwBhXUj915l6OObEKjw2m6oE6bWKDBNsSyRviTx
v9tBmhJFpe+A6Qn0xeVWulZnKIu9WbNAEbXYjVoLI1VxGKx22Py11CxFrmd/vtTS
Y4g6s3wYP5s+Iq3F2nV0xYoVOe543hkdPKEc89ZxlbTHhjBLyVpGuutnAXncZe6q
W8jJ4H9I8b3BPeMpWmdfEfOCU1lNK22g6P+J7X9oHePoGkI/5r3A2b/GJY1Lvy3g
+vulOaOvcDJ0FuCAyBjnSgG4OBzbeXObkSqMlybWeePSGGxsM87FmVLsZHyPr+SR
vqgbblVSd1A6a4KUqoGO8LhUrGNCqC7VR8Q5XRBD4cbeu+x/Fm1v8PbY+kz8EPrv
qxPzusFtmjUBRRzsgI87+ywFXTcTSI0j3Yk82oQ8UaP5GfTK8vxg+IcpxSo+O4sr
nZycgZ86wu9PkNeGy4QkeHpZ5Nk0ByVLkXJQP3McQr/ubfoUoz9D9VEFifQKKGNc
HPEEhXO+1E4MV+3B4Rx46LThBK17/cG1NXKIJYixyXZrXJmCml/vXefHOLfVaecA
V/pwjBtqYbgW8KX1sXVeDmvoO+StJmn5qsmG2w5OWyleU4dGnSIgW4eHEeRjSFGa
r564eyPCafS8YmO2QylMFwMqNHBPSEQyeKQZoHO1yvJ876eARY9JypXxi6SyWxPQ
OXridRyqGnl5WBm1cs70NWRA3CQuYKd8Crm2XMJg8aZzu+7/zOLn+9RfssG1nD3m
rtNSiczZyMvlBQ+/SrQWcYGUjG/ZYXGDFaUgp9r8okLXEeCbezc9w8Gz9m5v7Tru
DFG5zr/tKuEWGsIWoklWyIc3wg0zQmDgiV+NwtSHdbILunUcIdY3SkIwP9D3pwjN

//pragma protect end_data_block
//pragma protect digest_block
/qS89Rd5J8C/GG9oSgNXE8vMz7k=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_UVM_SV





