
`ifndef GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
/** 
 * This sequence generates UVM TLM Generic Payload Transactions.
 * A WRITE transaction is followed by a READ transaction to the same address. 
 * At the end of the READ transaction we check that the contents of the READ
 * transaction are same as the WRITE transaction 
 */
class svt_ahb_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);
  /** Number of Transactions in a sequence. */
  rand int unsigned sequence_length = 10;

  /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length == 10;
  }

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_tlm_generic_payload_sequence)
    `uvm_field_int(sequence_length, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    bit status;
    uvm_tlm_generic_payload write_gp_item, read_gp_item;
    `svt_xvm_note("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    /** Gets the user provided sequence_length. */
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(m_sequencer, get_type_name(), "sequence_length", sequence_length);
`else
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("sequence_length is 'd%0d as a result of %0s.", sequence_length, status ? "the config DB" : "randomization"));

    for (int i=0; i < sequence_length; i++) begin
       
       `svt_xvm_debug("body", $sformatf("generating tlm generic sequence 'd%0d",i));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             > 0;
            req.m_length             <= 1024;
            req.m_data.size()        == req.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == req.m_length;
            req.m_command            == UVM_TLM_WRITE_COMMAND;
          })  
       `endif     
       write_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm write generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm write generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       `ifndef SVT_UVM_1800_2_2017_OR_HIGHER
         `uvm_do_with(req,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `else 
         `uvm_do(req,,,
          { 
            req.m_length             == write_gp_item.m_length;
            req.m_data.size()        == write_gp_item.m_length;
            req.m_byte_enable_length <= m_data.size();
            req.m_byte_enable.size() == m_byte_enable_length;
            foreach (m_byte_enable[i]) { m_byte_enable[i] == 8'hFF; }
            req.m_streaming_width    == 0;
            req.m_command            == UVM_TLM_READ_COMMAND;
            req.m_address            == write_gp_item.m_address;
          })
       `endif
       read_gp_item = req;
       `svt_xvm_debug("body", $sformatf("waiting for response of tlm read generic sequence 'd%0d",i));
       get_response(rsp);
       `svt_xvm_debug("body", $sformatf("Response of tlm read generic sequence 'd%0d received:\n%s",i,rsp.sprint()));
       if (
            (write_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (read_gp_item.m_response_status == UVM_TLM_OK_RESPONSE) &&
            (write_gp_item.m_streaming_width == 0)
          ) begin
         foreach (write_gp_item.m_data[j]) begin
           if (write_gp_item.m_data[j] != read_gp_item.m_data[j]) begin
             `svt_xvm_error("body", $sformatf("m_data['d%0d] does not match between WRITE and READ transactions for sequence 'd%0d with address 'h%0x. write_gp_item.m_data = 'h%0x. read_gp_item.m_data = 'h%0x\n",
                            j,i,write_gp_item.m_address,write_gp_item.m_data[j],read_gp_item.m_data[j])); 
           end 
         end
       end
    end

  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_tlm_generic_payload_sequence

/** @cond PRIVATE */
/** 
 * This sequence executes the UVM TLM Generic Payload Transaction in its ~m_gp~ property
 * and returns once the response has been received.
 * 
 * The GP instance is not randomized before being sent to the sequencer.
 */
class svt_ahb_directed_tlm_generic_payload_sequence extends svt_sequence#(uvm_tlm_generic_payload);

  /** The GP transaction (optionally annotated with a svt_amba_pv_extension) to execute */
  uvm_tlm_generic_payload m_gp;

  `uvm_declare_p_sequencer(svt_ahb_tlm_generic_payload_sequencer)

  `uvm_object_utils_begin(svt_ahb_directed_tlm_generic_payload_sequence)
    `uvm_field_object(m_gp, `SVT_XVM_ALL_ON)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_directed_tlm_generic_payload_sequence");

  virtual task pre_body();
    raise_phase_objection();
  endtask

  virtual task body();
    `uvm_send(m_gp);
    get_response(rsp);
  endtask: body

  virtual task post_body();
    drop_phase_objection();
  endtask

  virtual function bit is_applicable(svt_configuration cfg);
    return 0;
  endfunction : is_applicable
endclass: svt_ahb_directed_tlm_generic_payload_sequence

/** 
 * This layering sequence converts TLM GP transactions into AHB transaction(s) and sends
 * them out on the driver. The sequence gets TLM GP transactions from the
 * tlm_gp_seq_item_port on the parent sequencer.
 */
class svt_ahb_tlm_gp_to_ahb_sequence extends svt_ahb_master_transaction_base_sequence;

  local svt_ahb_master_configuration m_cfg;
  
  `uvm_object_utils_begin(svt_ahb_tlm_gp_to_ahb_sequence)
  `uvm_object_utils_end

  extern function new(string name="svt_ahb_tlm_gp_to_ahb_sequence");

  extern virtual task pre_body();
  extern virtual task body();
  extern virtual task post_body();

  extern virtual function bit is_applicable(svt_configuration cfg);

  /**
   * Translate a TLM GP into an equivalent set of AHBtransactions
   * Return FALSE if the GP cannot be mapped
   */
  extern function bit map_tlm_gp_to_ahb_transactions(uvm_tlm_generic_payload gp,
                                                     ref svt_ahb_master_transaction ahb_tr[$]);

  /**
   * Annotate the results of the AHB transactions back to the GP
   */
  extern function void annotate_ahb_transaction_responses_to_tlm_gp(ref svt_ahb_master_transaction ahb_tr[$],
                                                                    input uvm_tlm_generic_payload gp);

endclass: svt_ahb_tlm_gp_to_ahb_sequence
/** @endcond */

`protected
-e=KCHOG#9HU-[U+Q1[.?c@?>/B5e#afM8IKX4F]TVAegWSCe=6e0)#-6G)_bKd6
GF]C1QTK#3.S(FZ,G0VdEbfg@^bTZU\dIO?==-)9/>M_CW5G[.64I(J0\<X+L;BG
Y=TfH9>NS7KcIGQ;JCF@/ZXJGDeJYIJDUfK1[DLQYce03;FVa0.U+IAI62IGgXNP
7A<B&GaHU?0CX]cJ,dTeK;HA].FI2R>Vc1#=9K?c/-]U?L^],DNSK<LXb(c#^gQ\
L5:5KNVNPNQWdV-I18W;7)6eZf02d\^V>ACQ75>AFVYWa#GE#6I_632\D2]a_XGB
QTg3TdRN=DZa#f=,[-2]Kf\C&.+<aSV(1O@\YQ3.D7C911[<.dT</F.;K]Q>COG\
0?B@?_YJ6X):^e2gQ:RT&6JORT@_]4?YL46-KZ^]JI?HE=CVY?)JQb<IF(3R.1?2
S5Xc]IQ\Ae:g==KMcL^C);0@KFQ8#JJ^gM-=#@FMgVgTbb7+)\_=c.&B9[ST]ZLb
8M6(Q_d36e;]/CbQ7,-3^CHc3U8X/Q35Q=a)<G[7Kf&W0J[U]S;Se&UV^.=<F<AG
f)A;@Z_70QU,2_6WLG+3add9e)\\Q6MOK,Q>X;D(e^;?)RGgHa4dffU:ZZ(B.E=0
P4H:4AdH#HgfZ9BQH3\C)=D:&CJRAY7gT/UdLBJ3S6<92eaFgPF_@Q.YW]+>._M]
\:B^>b^7_BYd?O=J_RaHMc<IbR[1GTb/B@QVJ2CW?&BbY^NJd)^fA;;\7)G\IJI;
9XX8d:\(-PW?C^eDG1:FV/4M#U<e^&<0YJRL04bMa_eNK.S:BC6DG]:W9=/0,V#,
<SN(-0#6afNBa.+7I-V_2cNU8G+QXGcVBcFCJK@g^gb6CME5Z8bXP,1EJSgDM12+
X>&@Lc#QG,DA5<aR#fRAQN2Ve7#N9CCJ&-aKXg.eD>G[:ZH=6+K)2fZ&92F=SRAA
O/1M#?R&8gTV+\&T([5UQFf/?Ke.c2JN4R6:B&b6cVUHTf,C67^^4)fX<D87O<F2
[CW3JQQM;XP,EQX6G[WXKb.G#B.\fB5(Ub3Uf,^0J?MA#H>52fSGe(Q&4)e.Z/=6
9JXT=-4d#&8P,G_@a@HAFVc>#5g@Q-1-5+F5bP//HMLCUGXWYSJLX6<>N&B&)4D?
\N+F@EJRg.F.D((D^VcdWUB\3I+7?/43bBNW&-\QKI<4c4.YgSZ1g+.VUd7;7^]>
5MH4B#b631,&63K8>^fMY6f6a+]Jb_OQY1RVgHaA;.E5<<^_E[RMC)0\S[M4,B+,
7K=\NfV,A6Q/.X)E/JO^c3VP&cV[3E])UD#KZCO)2eA?SfP?RJcL]@?bH1:IL@63
cMOc3MUS.4-NBIU@+.EHD6=ZZBB\1TfX>(Sc[9APSYgK:CQ[cP1=18,MV8c\a=,6
6O\KK#UT;4VVVO8?VOY@MPDa_)L61@9b.8NcYB71#T37-._//IXDCAa:Z()^H@;B
_fdde^FMe5Q:b>_aY/FA+c]UINX69=g;6[)S808[+8;\OX-BUe7BX+f:QF[eRe6.
+A-:V2?E1I2&,[f>?b36,8-=cBMB=CW7bV7R.f\N_FM[O@9:T;T]Y7,?HG&ME(HP
ET++(g1fTJdaHTfcTONHeg1/GaF4cT&_9SgD\4Uc,#4[+JPOK&#:,R1UCUE+>9\V
>#THE9c32GMB[:,9N&;_<]\-Zg)=DCF#:\gVe3g2gca:=6)9O=+S5+EF^;H8EF;1
SXQZ4W9)I6V)RCM+&KZ#0RCI5(9b>VcTd#7(C2)NV6eOYFM9E0.F5Y\;&g-57KfJ
BP7&,bWMf0(\dKE/bRg,YTX9=/SAL1f\9#a97Oe)@H8a@[dL[?3H5ZGS7BcG8)]_
ATc[V(+Y3Uc]cVGIN3W7>7S^J0U[.G_;A\;0J(B2Z5ZU.MLW&BXbW_I5;@/G@2HU
=g(B^:(?_O]BZ_aAcOPbHYFSHN&b5PMTfegJ7ab<Y73D#f:f[^,#>;KBacV8E3D@
#&R,0G0^[]):L]FI4)\<+]CFNfbR^T#fUdDZ;=)X:C#J9_;/--KSC0dM^,M.JU7a
[9:L5[5+Ue>&GO1^(4Ka+.QfM\-<<V6#/PD>8)7#DfYBDf3;-Ed01NVZ?4L-S]OP
LSCXHJY9T\L4X7.+@0H:T?M_U/,GOR)@d-5L<BC8MMELD\>.FJSeJ.c1DX19\bJL
4[79K@WNMgc8].Y>2\b[.e[N=W=^&6a==Wag87;S+4DMIecJW^E;_1B4/1,;cQU^
IHU((D9XBQGD0)?:gT:bN_dA&>Y96K(6SC.(TY3.B5N#-#3dY;O9VMQ/0S_1R<9K
5e84S5D7PPOAR[ST[=S8);NT3I@_XI6)dK28F4G6V35NC?/;2P&TKZf\XW3ILBIE
6L3#G4]24<DNJL;CA>=DJK[:;O>gDI5P,GCbLgK5db:A(?Q+2#DJ-:B]7He2>c8A
&EdKdBY<[;WLF8\BS0=c2OKC^7ZE:a+=WQDBJPH1=+3ecPPA^R]NY@KN&EVfUe@^
4.PTd6@eGO<W.OT2IN>GEf@HJ#^4DL&JKA-G\YHHbf@f&6>4DX:YKcBc99SEXWg@
S+<>gYD5_]CQ?U#B-&c)9_1+/E_XPM._3OTa34P1IKY-+0YSSVTJI?8bNgdV0K/F
&_a.:/]6DP]0aLRC_<,W[LIL-CQS81I[OK/=QS)_>N1V1VAK?aeC:XB34b-1QXJV
YTG.WdO\A.V&TdgU6E\N3YENZEZ8,Z4<:_EdE2IK;OUOPSO0@MU1SCd@4g23V;@T
J>OTC3=g<&8-3Y^4RYM)]IE4a8#9)cTHF4Ic\L;/[eH65#L83@a7ULWYW(Kc:@V&
cba:N/eQEJdA:+2ZYQ.C^A)3^;.12c#[+2;2W?[B:b/^IQIfJFgZNQOW:,(\5M88
#\O_4PN]0,CdEHNZ4c?e?,)Z@CQ684EDZZbYc#F+F[@8V.X)#07dKX.6a(Ue\3](
/2IPeH<ODB2TX&LJ9-)O7]A[J<9M08J^g\<TF4SE\5A,Ye3&ZNMO^+36N(.U@N#W
[/D-APe5P8W-cE8)[D#(<[;MM>-V/H&fCR7)_UZ@W?B]4^0c]WFAYO1]5fKOB.,=
-,=F1Mc5(9FBeRS4+g:.PX&Z5c^WRVVA9L16>#/U&.XVa2cOR+&0(2aWBZETLLUB
#+fVE)+E@b1CPdKBcScg)7E3QR(\S245ecf^aUf)5\&3>GZZfaf?MT.7>1S,W<H[
C;U2_V]\:,cE6fF?2Z+_W4.9MD>>C4,PX4E^Pg0Pd&,;,fK3STOLcJ]a?SOCUJ8P
_<P?_\bJM9.]3J4+ZcBH1KP.GE\45F0e22;?cWa8AOB?#cO+U2BORg^;=4T;1><S
V==#>EY_MNH+I5P&R[d3M0G=QO?<@W>D79[JcRC0.E.UL3VM#;P0XG:8Y,0#5#3U
HYCP9NR8/Z/ag<EB:A/#):F:Y1IX4EOT5T47(HCTPBd5ff2Od5M[:CHYaDQ<cQO6
[EA&f(GD1ABYTY^0Z3c&:D-gB-LUJ;Oa_<S,L,T]QTcYB:\9)I4]MC[[^3aJ#YO#
_VMP9T^17J^fUJG^<FAR#CSIQ#G?0,N75+V(<W+Z3,Tg:.a,(.6MZY0@9d0-J7S:
N(VC^-5HDQ9]LW+2CZXI5g07V07?H2S)0)6acc[&Q@E)^&Eg01fb7/Z+SaO<e)4Y
M>6LXRH/YPFYLON8_L-cPfW\.2<@>ID6G&C)4IVJZ0W)2f^,FQ9PX-..GV;f=7fd
8bg^71?cIe&7aN+=+DS?EW9KI9d/-(Ba>M:I0;RCM6(E/S4R=R6\7Sbbb.X=KTgC
9/##L^^FD2H?S@;,#1V.Q]^8N3_SB<V^)GEN2fT@AObSEB8]=NLFHK66\O#XKOPU
Q-@(K=.HXaLO^EfB+fcF;@dQ(T4#1@-KVH7G(Z>5[d)dDTVUA\ceC[aJ#WN.H1dK
V,96efaR#36.DdQ9-I9606DAHV3,dO&BS?TN0]Fg0VN/7ES(53]T\d-;WY#OEL)/
Q=REa\PBO\c?J,V..KWg:-32M,(PFPFH4eVQe(PU\+YRB5]V;dRc3\5QdOa\fQL1
[>D9d&g,a]\810dJ[(XceJ=XEbNJf-S;Q\BO+>MN5BV3YD8cf=]Z>C+gBN4<)X6)
B]QN6f=bJZ:7<I,P@^[V.5P_#Vec@5>IBc<ZTSe/;X6?U8CE\D,KZO<K\dX5L+e;
].UL^6EY_/WKUY?DUUQYg\1U8O5d+PgdedB9MbC@6Xa<BQ?U;0IE)4])6_(PaS-1
5b/6cX@4GQ=30AeG(YY3+cI0g?,KHKL]VaQP7E>=-5:@)OGJ)4Sb-=Fb@L1fE8@9
C285BK)\aH;S<XM@5VIMG+8JD&V:4?@V)1(b?;8OCFHEKWHg@//J[VZdXS(&KCKM
RKI\Rc/HVAcMJUI^7[dPDKN_2[QG72P^XFD36f?eF.Q:I;/(gG^?=dMbPe06,(SB
2&/44d4J^4LfDRUHN@cLAP&fO(AVfZ[D]aJd>He\d0EY3dPKf.SECIC2gIK1AAEG
JPS94)6TPQ#cG(X(\:aZ:>bfcNJY7,U06/_S]U_\KCI6RcX7I4+8SYC:<g3D1LJQ
X9CZbK;NYK1;<-/U3c4;?M^_;XI\Q=;J3)K02JRJe18J2PRMC&a&WgK>4V_3>Z(]
@1,U7([7JON@DTH@FP(_U5RCWOE]?\D+[E??GbI,\X\6B;Y3gE313)IPd/?34#SC
^C5\_QU4>+4#da,UgYV6Ec:S;E6<+#fR?3F@3)^?MW811@=0U242KQ^<K0DQ/N>e
ZG1&7;GF_4c[@b/SF0f]WgEUKIED^AE/NB\1JfF3.<Ff\JP]2GW0?DOJ^\,M0+Ue
S=?)GARILa7HXC#(D7LBCeGOJ/Hg7P@X5f3\A.DL^6gTJ;)c81B-0RH6DbE^[/S<
6@JW^W^8_VE[E(cS^CJd#GDXRNea+]TZUAXDd7XX_V+BQ0\AB-=5Z)8JY@PZ8BfK
e8a>>K(Q(E#AA;==QM=JREQO1=aO^W.;TP(NLc,I0eHGK5QS.:L-;0c.DePf,II)
/ddEN#f_<YMY@dLLU@g:Pc:[I7I;f4Ib?DRGNFW:)FTfNNAVG(GH(_Y#.\3ERFeF
beQ((-D[c/P_G0cU0C(\Pf&Gc_dJMAe_N:XQ[f8HK[b7FBae<^4\b/<JbOJF&D.(
-fO#AZ^C^&:\VX)GYUU1NO9Wa#M0Te?^6TDCWRRT@;H(G>2/I(W>d]U8J9T)F?1I
AgaP-(>85YcI..eEaO:gI<XI;fIe^^O)F]S0))dU/7I79-bO-@6OPa2H_aT)40c4
Y92>\e>,+J;bTb&_D[EG<J[=W0JRJ]Z9&)R+;+KY8W7=S_;R]-58V5=\NXQ;>F\)
d>9C:M>KL1XeFg;0;DFbNYBJf,5HH(/e9Y_ab](W3d>LOY0]\3J]85\af5K#<U=\
=^[<3,-6W9gO7DH<YSdVI_Y(Vc&[L<>+BFT@SRIOVMF@IT3T+f:<J=c<b6?I/0R=
9S7=D7=3CI1.;V=,BcXKFOf7e8F<SMJ[5=ILX6=ZFI^OKQ<fG)Q<_IU\VA8fD8OD
_KdE3bdU74(/R^ZC&/[F#+D\XF@EJYAHP_f0P&PL&K+MWU?^7Xb5^HFcJ^=D8gb,
U>83?4FE+=Wef85bAZ;=c-[A\\M3]>N^5c82<?4A=ecTP32(F4M<C\.e.XL5QdHa
/#&)?I_aPeB_-S_@g[2gUg+HB:KABW.5-4>;eY6R7\P@#g.c(3PBG-8G^YF.#A<]
6_-PT?05ZDM]I[0MV6FaMb+5CD4T:WPcN1UJ.3e7UDN]=.H6^@]O>;;(^YE:XRc3
LCUOPO4,1&&ec\(;FM#I_LQ?;IR[TXa?>@>J:?X]H1?3EHNA]CJ;2XA2)F:6XXAJ
>ZK<2JE]<&38AE<:]>WTW7H4.=F9-^e,M(1gcP[@5(V^4FHg^S6OFILL1(T;@5,J
9+G,._-8e]81-O,J=BXFF_93Z;_MH?5ZAF&H([Ic;Z1^6Z?CA(#<6Tg6BISV6JcU
?fPX5L4PGSX-/1[4:,-]R#LdUA&BFXM0@0:#F=J?R9-:NYd/XGTF<(^g:5OZ9b&=
/OGRM^d<4@f7dL=>.))61B[=DD60R9)90bc-G>c6XU]J/Pe@5TbOCNQLVC?YC9aY
I;L)C]Y5KUH:(2K2(>FK,U9?T64G;_9SW^])\1,;>gEBM)I)6Q5QEL<0Z@H137YN
M)P0Ff<UF6a(OT2V#32T9K#QYaAY3XELE2=(L1C;;_;)_GaD[/_46;@C7R]d?S=)
Gb>M[G1BcXGV[1eg(TNS=fO:)V/[ZXKFKL<\,DLN/N:]bdL<L-e3(UQ9N_5A4(FD
GE>X^9#f2SS?Z928fS8IMR0.,g8gA[#OeJ?(TK?8f;=+3VM/d?Ifd_NfSIe6,/0-
01?S5&R[<IJ&D]\g&7CM+V1RNI&T\)b@bCI3)(:<F#@Ge5gT2?P@5K?&7f987[5=
I-<LP.UI8T2W-6M9c<gd;]7T3d#X/ab1H-0[/B679W/>>EMe1?S7,C<M=2@eCdS@
@IIaR1b@F.Z^[MRNb+T)EOMW[8\::+/B>DI&.-]I9L:>T]:Z#RNNdR:f#E?3-1P8
(_E1LRD,Z)@9ed;.TI=U@bGN/:.6W_1#(E)Vb,]Zg3:]d=FO@dP9PL)0cMQ\_aX8
eOOFd#CCOFNX>-8V&&,/(:I=4)SH4eVC,7abgfUY.95/^7G_41XEGEM;O47aWG?<
TYP)G#9Q=Qgg1g9D9>&ZSTTd^@MF0H>;JAGP0YZTLN)aD+&KH4ccf^@=Ma4@9:H#
3GP[2L^3baO#8VJ=7-&E)J/LIR.+BVC\Y^4^19aCf-AZZeW0.AIK#:T\3/T3;CE8
,9-^.-N_DGg^AB/HNNC4a,eJ>9]/]?M],I_3,N&EgV)N&<V:<0=DQ-:.\C;MP9X(
b#2e1HKA3I93:@C]],Y>8IJa1c?-=NH,E2/[F4I?X3(/g#U.+_X7\a#cR078,<a8
_W(\gH/T]Eg/2BMIRRLYMca=_Y4(,S9@EUL[-EXLNUg@<K7_41O7>4_d^2@N.,6N
JCY7BGE9N.5X<>QLQ9M8P-FYIQTJ?0.L_.U.@P2+F5-T@Qg/2;e(KD(CU3=IM(Kf
@GCR8:ddES-Ya_.W>Q9[\C\dO;;.GaXQ)_Z,>C/T0+BZ0ORc[Y?4RRDL8WFfKWYb
A2LS2=;)1+[R6L=JYT&TgX9WES=ef=@e+E0R=aZgD<+eDD\]#Cg:T:)Z?]>PfYR^
O3c@8c\2/)c.9,PY5>X6.<?L;#a?QW;#fQg6:>BEP]P(-RS3d3(]?)E/MH7A<Q]I
[UU6[b[-Xdd))[8eJ4E?P5/EMXcMaaaV^>:ZAe\ePD:QI42Z?@2T=-:4=:><?dCP
?-EFY^\._T-e/U6<4#&],Q;3&>:B:S4CQ^TY_>6#.GQG[Z]D(3&7C;FS(BDPOU?I
[NEb/fU0(K>L&b(MQ?L4U[b:4QZ_9cD/-@T]W>)U4b?BGA(3^6\[;Q/cG@KZPGG9
Za3D/Q_@RBBZ4#CF&=RQFRRdN#4#>9P.93:Y958N7VOD;4,]0582/6\)dY(((R,D
<<fBXC@,=XIUfc3J6[6MONKH7V9]7^4c]e?/AZ_19daC(^Z;P@c&N;HSbU?E923@
^12&[2@C;C@g3RSA(X1?EF2Z)Pa+X;KCVL0eSI:6]CB>YbT21c]0\d\OV6+\Y])V
.HDN\>R+@WYPYDd;U,/?2S:RX+LKP5B_QA_D06YUIMV?KJ<_b5>eE+J-d1a-/&<V
d1)1J34VLYgH:=SM>@g0-F46<T6J2?<98U#>M@G(<-/KRR+9Ld]=OILG-dN4..D+
JTgc0MJMI828B,[LW+GBM46>T;X7+@aKC/M-CN823<GI;U(>?,g[/;97GF5a45WE
OM4[GU9<[L5LU\(&g^BX(L_V_<8C)YB-)+SOYU#K:OA?G3,0H0Q90R9WO:.XLdSJ
2R]&Aag<<N7PAM/UWe,G>(CBS-1LbS40@Y?+N[Z.-)gY@Af-Q8>4.MEdHG>B6PXT
V#3ULHeNe=g@F][9SSFUXfO.F#1HT+?&D(5Id@].HM+7M+&+?Y@/0a66PMFY7g\<
L>U]/C5O2P]DU2K0Z>R&7G&:&Q56?H0L^D\c0,g&,g<cW5)P4X7IA63UKJW=C+5=
C#AZFW@=8QV>E,IP:JB(QDe-19Z=]1f06]d#IUU=B&g;9-.>9K_AFK=R5E\U]2)S
GbVR>e?6#<Ue8/?WHJ0#Ke;BS7XXC_LcOGdb?6fFDJ#5N]5>NO2\d_H;A<a]>a9[
C7Y5#([42aJEf+^X[#V[5Be(,UICNXb)UcVe1,a2URO.ZU_ZP677G[2P:fSS&EHY
KGC8AFf?ZZX+2L+:]TB,SR)KD,cPED2N4CT&Y3-0=/SN:F&^FAN,_VJKRbY?YS#O
@6c,YMPPL6+/KQNgQ=744UC[,W?1fU,;ONS9+F]9#cE&V)K><TPR:0U3LVVJS9Y(
<TV3Rf_&_&.#0M[5/SOcP]J^6D-?52EGOQ2P0L7b?Q#_WV<6<9+Q6<[(^>1D(CN@
T7O\-UE3XI^B]>2(3#DTD^:<SB77f\YEJX7HgAeecN^2-Gf>0PYOP,#fWNfDI5-K
_,V5P)+-[AIN^)5KFR5^7&Z@V-?YDgRM#G\X@HCLES+@B^,?V1X9TcY.C5:WI2B^
#)G+_\,F7[NS)9A_B#_:aQaZf6;b5?\;F70T-aKL2:J9\R:451^]B2AG1;[/36PQ
)-e+.b8LXN9#&D^@Y+^[Nc^K-4T)-d[CCXcgMS6^3@/++L=fc?#JDE:4@JZ3gS^4
4=dS2&YL2/)<dDWf)ATWZ_FV:G02E,CC_KLFcT>I).D<>O>TUS8]1JNYCTUOR4+\
1O]^4IH=N.W.Z6M(AR^A-2DAJ(@ALP;Uf3<F,>O]LO5=:TTWe.FWH)I@BCOaRP?c
)b#S.-Y#e?Z^M]&P54L.Ig=S1S;AE1F6++;BO?92]XNTP=V32#_\SB>44g3g--R=
,]Z.C>YH[5/2B,7B]caK&=@]4(dEPGF:UCU>6JBLLW#B)FR;K/]4G<e^<I=dKS\U
P8#^@6WP80e7VVD#O?T0K48N&)#^8a7fZ?B[8Z/\;GXeMHgTOG>eJ3>TCS>)2;#?
F:0:F2f/O9V[<bB@+A\Z+^(ZNa#Q>Z(F+N^[;74H8/,J9[>BbKZKc,<OeL8IM;Y#
@#4fK/X=E5Z]6>+HXIDNY3&S&@_R.1)REb(D2J[_W/9G#2^JT<FgDRU1?I0@<b:A
DV(D@e?S/F16Mg:HSFL[06c6)B3]&aUUPR?YJKLTQ9I>BNfMK^@U#f@fJ<VI0\]B
\Z;fRD#9=/@]Hg<-FYH:9]NN6]UWIYfF>6gO@:(g7>#XU+=<FY?G9+:CPBY,P8Z-
=ISLbG:E[#8@EB]MI@F9@d_<B=2QAe15b?5+d;e1ggCO:#V+XRb8/=?0G1NNJfMJ
9bYf]-Q=B24=KA973bc1#&@Y=84&J?QG;W;W5H:#B3]99UgYS-#:M\&6]^QNBZeR
\0=HHcf/XIQdGHgf(IZc;2K@g=P;;^9U99#6M._=ad4D:CF>I=#(IZ4ce)N?X71F
-L&&GFDW&DV^6RE1X[4:XGI[fD;/?C]SJQ>)78f,]S8^24D=J5J\0dWJDS86AT6Y
VLWMfg>J=WA.9>.C.W3G=RJ?]PH0QNY.bG<Ie23LADAAOWT21.?0dO.\fC7TBB&.
cHY]9:(Y12]GM42>QOaAL<MggYCRK^WG:,c2LPgTc^H=9T:2I44d^=7J1J-#,\J_
I;\&T@-_JTB<:0]?P)a@XNRNNU)L[13KFKM_^S_8.A)7[FO/.2W<0F/M(R[3N)-=
#8KeJ<UHXDgK2EA\b;;4.Wg]<<>dWFWYcb3OWJSX?]X3aI7X]+Q-dbO4_.GYPRSR
6F?1:eT>79fXdI<C]DZ?_5U?\__22A26_(;Y=?c,:[PLV:]Q8d7f:M5X.,TVI>-4
-HJ.5KUbRU&eF8HWLO9d:B[5TTb9J4ZcZX+8IBV)-Ia_V(]1YE34,9V,K<bK/BUZ
E@WgX(=:2/G<07A(ae4#5\8Y:WNZ6KW]VO62HU0-5LM8.>DYQ293_R^23J3)gWCM
N:]DY>gSffg:@&Y?eK]HBbTa2AP<V0dNZG<?NTbP&gbf.WGA)(f-)XC=N1T_Wc-,
B6Q>J)N0VVXV1Tg[Eb5&P&Y+.FI=UMU1+HZc8O]dcZDQ6O)[BWN@<^X5X_.A;(1M
F(^=aUS^29LXUb:PHTG#eKEM<S2E&:6;LNcXcDFcJ,.:SDfA;#N]U=)<S5G(PQ\2
GAR7\J9?g.c7Kc<UBJ=/-_Kd+/#g;^M?UTOD_S719\DLDUT.7c.f61,.dCO]IL4Z
I\TPMTX]a(4IgN6WAJbg^N4^N<c5KJW?+A?#X,1EN,X\]_+2d0TIVJ3W5\,BV,W:
@D>9^@P<CWVH.B32W>JQc_GD3_:N2bTV[9KKYc0SW]8P]c1X/ZeC5&^)U,]gCZPW
DL^YSFTD3KI)4X_Q]AWK&a_U)^f6:X\Y5(K[dV=.?6g3K:Z]?aQ?2LP,S+T,A2@@
5cI#X@:U-XXSEdL.AdeBL+ND/VKFc&/R\0E8;Gdeccc]=:QC:W^L>b1UERg=&T#(
8a>>;fM=?-3GYXM[C:M/BAgV/+<Z=U26c/bRY+T5&Cd9+c\A4)OR=FVJ>?C+ONeO
UJI)9^O/D^]c)9]e#KLc(eM+7//,BM12(/W;UKD^E5SE58&(\UA:S-@&Q29W/Z_H
+4N+[3a_2?bfG,(QA])L]=_K:b6B5AS7@824Q>)EIf::\OTfaRc3HV]/RW=W;U(K
b+LCAf>P^](9WBQ58<XWDH&KIZa>FV8EDHYI,>@>K:Ug]D#SJYc70V>5_K[]N6>Y
ECee?Ta?ZW()&YTZ=SSbBX@P(,<:D^8bOTQeV[^OHP22JS/CU6ZKT5=Me2DU.39^
Cf&LRdT;GSROAJ,XBR86<He^GH_JUc&1/A_JAR1-]PL:=GLRFaRBAP7[:+N8?K?U
H[[HR\S;Ad9<IaX07-:BZc=&7?EW=+)D,YSY4_P/9V8.E#Ng;d?VD3@Uf[>O7HgJ
JV5:deb4ST()U@8F5\<EN8F^D#8eP1ZNV3K>-3SO2=28a=O;R.8Va-6=8Z1^f]aP
BZe#;C:d\DIIdL#MN8OB[9C4)93PCGgbJ?aK\bA,5JaGUKdV80Z+<E.?0CY(;_@d
D@C1G.58RH)7C7@/L#3E5)WD4?URV(G0A74e(/^M:b6MdZBXDDQ2Y;Z1=Sg@6d@O
a<NG5\LBU:((/ePVRV?EWNEZ<S?@F.6&)=M:[Ea@b)#JP<W4E2-KL,8JG.\A0ZE,
UA_#[IJ>46QEcI?5[M0+?,IRG7KFS,>fS+UY0QcRTN7:eTRQSSb<_NSFV7C0d37O
E?]V#11J-48(aeL)E^/2&:<LN47IIT]K+)/PZ3a3E,F;#-8T8/FJ3B(:KA2V8[fT
c<;APUd10+V0dQK?+?#>/R?TGML+NO:U<DT3])cY_\DPW(^fUB[)DO7a82+^7gTH
/9&f1ZQ-B>D\08=caYNKWKC)Uf?/eZGBT2LgdS)3SE342K1MD,<AK]^JB57aaaRN
g8>,6D3S7]X1,L9U>25@O]0[D#HP0e)M[GFCMJ&5XZ3T?5MT0HI/X5;5Ka-U->a(
^eFUO,&#YZ6OK;.)RW\SJTL9O?cLb+-:[+;4Q7d0OTP3ITNQeNT[0I(.TE6WU;a&
gTH]Z2;QXNI8]QZ)XLadW2g\=:T#fc;FZ(e>URbaQL(d=gVNHWIZU77dA#a.BY(C
F;B,2A&7B&Z0O4bAV>_VY/#9fW/#0b0[P]3>OA4NQ[<IAC(3M=O9aBXD[+\[7&W#
J5;G=/50L]e@K=5V)R)1g:MMd3]H3XEA_Y)WC^>RK2bdPJbA^I\K&HD39U:cTO]<
6FgS6)];;5.W)KP3f81V09:XX)HT_8#0bNFE&O?QcfS..4ZVKGPR#5M[eRM<2OTY
T0;4YJH&:939Y[3\S-H:32E073@TPZK/L3eJJ\Y5JQV?H=D3AO&6cDG(>K4L)>MI
\]XX[&0)SIZ81J6CX4=GDb[.--_8JU=N2.RYDOWJf7BQfY&/0C?3C&_;?SPEDDK6
7Id1^1-d:0aLW9GAJ>V&e,)[?JRN[KC99a-&QD:e+K=-D/SCIU_@QX4<]515WgS>
P&FZ/#@I221<Z&@Z[J0Qc[.MTN;(G6D?,UKX[67WLTa)+1\F?\&C[;c+Ld;._KKP
\1/:<e[AUY?\;eB9/>;DI.T(6#e]a6#]I4+DJG=SHZ_EI4.?=bIO])f(X_7S<Y@G
9C^a+UE4?FH\KR5]#AZ&O#7\JN2<FACIgER&X:ZJNGWAF[M.3]K0eB67^<SPCB32
>T=1/_)EH(LTX_^HR)AW]PJE<=Q\b;XG.IWbLYK:2/,Be&cH(efe]/>acUeMR.O+
GP^PaEI0T&cIK.#DJL@5?F3O7GN):I=@V@9CO6E6(U[J\@EV],7V\-C>BHD<#V=)
KFZD/D,#Rc(19E^4GO+4]U0I9,3.+@:BN>D[Te:]?E>SKB&SQK6XPPQ4Z]dSO=d8
0>)@Y6..G#X0S\KI;gI39.9cJ,;Uc(ba^(0L,3aHR@65Cb+4RYG+Q8BZMg7<:?aZ
g]g.0I>=#g>0aRL6J<T=d>WUI++3M(IB/DM==(MPCI-f@a89\-G@b&Y1;4>Y0DO7
39Q5H?2B&E:M,Z6Ge).DVB9Z3&T3F,U[V9-gS-H)QfbO527H,=(Y(FXEBe2>Q3?.
3PS[=WS7>K@(V_cPaE@@8RN<?4Wf<9+JD@_WD;458K;c6eNSf)6MGK<D]7\-&BR1
D4DRR>C+O_>V]4LD0fCOO^VV]#HKE^Z;[[\(gL-VT8]e5UK)F?-VXEg#B9IEM@AK
K\CRJA5.XJ,[?e@XKd40JORLA[-B0-Z.D9<T<gYC+g#)+/GFJR]4Z^0-d3S1=/U^
\JXAHa>)]/H1AT:,M?1fEfd/>,4,0R0M(843.J>;Ae\<_6O9]?Q[Tg^9&LKcTGEU
1UZ^+GJN2<daO_YJ)cNFf?-79_XJgA=Lb@S\5>aec?@YbM:b.&cfK:aVL4A7M>DQ
eZLA/X4VBaL[-B)W\VfZ[fc#O)7JaJeUI77c8U#a2EIM/)(ELW?U3\P\.@,<J;]T
#VWUfQbH&&B2#541cV=LP<[Ud#IeL#S00<2R0HOJVeQZ;6#[F?DJPgZZQ,(>1II;
#F(LRWGF3T+3.H@1IZDCE743Oe<#SX-a+U+eH-.)dUf3PT?/bg@.[OMd+V5/U9MM
DUCg@UXRF2YcYgLe5McfbR);_P-L.6c&ID)P<Bf\[KKYa7;B3WK9U584\6.+XM_0
^UR_PEeMA^f,.5FKP:#6BDJ?#2g;9J4DPS/a\AG+@B@#;ETPIKf8I8):B;TB2[PF
E-.UMC6;WX1H^]@]+)Z4\YO(;G8&:b&;g^MKUbaNS>2[FRO7[MG6L[PAc3E6,B^H
Q]TdQ9Y^C3X?#_U=JTe3<,>a#f.][&IE/d8a@]SD,0<:-[UM[C[I@8E7VIN)+;01
:(Ve09WAAZMcP2GbQ3I3)\;e?b9OBX7=d\c3;33:HHK<7QA-S(,DgMX1:0WHCQ)9
T;K_\J@(L)\BMcMGcb5[@bcNKZcON3#bU]:LJX71K8_;dRPgJ9-JAB[O_T6P<\WX
2=>ABU(2_L;cN^S2FN;T7=<Q<<6NA;JMPGc@eQcR2fUVJ>MFZ@c=T?9X4a;#+5]L
+c)b^OF,]6.NT7FfM_9U2H=&9W5If74:&0f;X]8AaN(g&2W)Gc+W-W9[1)-TbU[4
;X:5a9e0a7A^J.]56SEZ@?)/;5Y#14fU[2RF+eb>ZZgUU/<Q4Q97\6MFD(KJ>H5d
_OH[<Ca(8)_Xb&/Y)Q?bL;cbEN[=;;EF.#2QMP]WG-&^N[/aeFCQ^[#<76LeF^Q-
D9F@T9QQP>]PeeUE3;)(3P:bJ^KWW=D^1I?I>[;H)b8ec1)]0dC,J&#DMH<OOY8<
O\Y\D-3Td+[PSJN=45]Q8;dXd2bC?CcH)I=]-#2Fde#-(<P?6=6GDaQ<8M#06G^1
BOGW(.Yc;Q-);-U4Vac?.)<V.3)=I?5QBXK;9c8OU+#Fg;2=g_F9db)19^&HfafE
,@42/N5gRYX@_+DV()d:-QMRQe(cE<bOOF_=,:AcP.93QefY<Rb8.>e<Yf))^O3@
>DV^Z641^:NWaJ/OBV;>GAHcRBA^8&S^G/4<OUbb;#U<GRRQTTCI/Af6beV&-GCf
BJY#WLJ)_;D=<a0->LS=BAg2-?Q8ec7XQOdBL:.-/L5)KbT&<HNS0Q4d)Z0L3EU+
f6>R;A6(N-IG+1gNS-aRPeFdF4<V[Eb5>1g--Pc.YH+-D@W;7;CQPg_-@-;D\;(d
a((^K(+d2I&1>/;PJK4\V+\<[gaWga0JH2#S+N5EX[:D[bO5LMOL0;#K2^;fG]-;
;B.[ScS1&[Z@7OFbgI;T^fZ9MM8UJ6L.V[][UUSBNUD[fMZZ@bNS8?cf;D;[W^?#
?a(@=QLO_-He-]eaINPINQ/O5[O&CLY=FGaE((M^]);+X6>9^^1C3eWG0\XBeV_M
Lg^EYE])b>BXaK;7HZS=U\Q6K@d5Pc@LFBR&NP^Z@4OE5H3MJ55/9-J/9A:E5a5V
Ece@;,egM4b=AeYPR-Vg\1RD,CJT5D]7ON\4/Da2d0<5:6_6bdTT9fV<L]cMd0K<
g6-N(P@[SR8/MFV[Q+Y^Q<_fAgQQ@R/-Mg6&F4E/O[Q+&FI^(f7X>)N;NNLfC)e_
RED+f:)^D;\bX/83b#V/_&I_A]+A,^[?[E:Ad^7E:,Ta9VYG4V=^Q1U4[3HQ.Z:_
N1BMK_1O^e;.^62b>DB+IUaHX:B3Hf++#_K65:g-O>\YYOdaTaZV1X6b,#70J/;g
&&7:C_@5Rc5_,C2P5T13c.6RDM=8H&;Y(&)C=/P1R_MXR(6)U]J8[Ke6^-2G3U4+
QH24)QQ@>Q^R#Te:dVZfbRMIPF4M56[E0UBJYYbK8^bTP:O#R8FQ_>D:BR@gcU@V
U7\H]62fK<2A=/PS>F4c2E]\&S;c<(YBa+?.;ZIT>=@e;5f.6=dA_0OGcV:7TG.+
?7b2F_S#_cKc5eb[fdY=d>C:G]c:3X?d;QW^CJRCLL6_Na4+V2V&d4+HC<P[OJ.S
N#6XfR[RPS@ZV)cKc.GVAa<#[L36fg[OD^16ER?]+G>KFDP6aM/KI#1AcA^^6-M>
F_+&8Mf[[N(WaEFX_(&H:#KO_R0:RR>dT71A.=?S<Z&?A4-7YRGQ\8]Hg^X:0I_K
1\fcISE_OfLaK,X9CSK;Jc36/I1557;>A@7:>^8O]>T#b)<D:7?YeA,1fNWS-3&7
A^#PQOO;,Z>K=8a0+37b]2=ZWKCXPe3(8PZHe(Q3G8.,gARSN3V\^\>_GVWE9d.&
X?McH]#NRbXc/>IRBVbPcXc]UYf[EZ,eC]9HLMFSFC&9>TC&82d&W?:E;]/b_PL6
2DRFML(HIC0YCJ48f9WfeFcC=X1.LZDEZ(e/)A-I/e]_eT/A,8Xc&?C0HNTUCM)J
QRJaTe08ZN2A>KF@eQ^ZgVO\P53_?J@c26_c#ZQBCW<b7@IQ2gTO-KB+>[-@NK7-
)VQAP@;#:Yf;cC:])/J1J5,D]9NG88YEG[>7[Y3#g0e>aDUf^.B[Y@c93G9]SR)O
e5fY\aA/(TL,5DZ(fgD2UTT8GSaC)KbO=EZ0,.e[d^QW;UDP^6bPU5_E7I=-<ONT
..95:6EW&H:gFZeD>YU;ENK@JU.aH/I3VA=BcLN:+_N,NN#<aN?)Z8L3PdZ0:a-)
efUK[-?N.61N6GeMP(//H8P(59Q8>WeY664)_]EY]6LP3G6^:X][@MUb8I1VbNY?
,]TT=&?2P2WTQ3FgB.f(UJWTZ_672c/e,E]Ma3abdR2_gB:PW^/2VHE&SED9AUC+
_Ua#I(L?e26+=6K:_eW><FY8b7HD:BOQ^\OOSSYJE)TU]V96T9-c^)^SVaQbOT/C
D+b<?cU45Q1;7;Q;8X5U[&gXR<<R;c3af@F&bTP6)+-4&.&e_+5V]/J1D7c7#L<9
2)0CaCSE9V3^]ea42\:QN^+cIIGZT-LDIe4@R8LcC<<)d^VSEF\ZI)gD6/N4EMbe
BBF^64->2V.:L>E:e.P+O9C2/b@2RUF-OF,0721dO=V+L8[C8F6\,XFc?FVB9TW9
-,e.[+aFN1+EP(.&BVKaR4>QeC)0a9BZZgCVcb+\6/M^c>40D-Ie<K+GG>1.537V
\VaYD_X:GDJW9F,;fQ3#-[YNTb3XWN.;:7XN91VN,[ZI+#1NUD.c.0Q?7fMN[He1
3PJf6aV@?I16(D?B9#\J1-,GOG40)&H#IaT\c)E;;:NHFbAY.f(fTg/(YS#_&W/d
JH-JW)F8F,SG5=OEgf_Y5F9.f(UD86BA1<-g<JCNZ(RY7Ob8W1R9TZ&4Sb\<)CDM
/5@Y@(B6T_)Hb:-cM\AbALDN4Xce;];Y>+9gYWW[4AY@BcS4=/[VV8P1&1eBO2+9
HG8V2T,CA3K:f\@,HbXHKcUX[P9>XBLC_gLQJ;OR5=[P/EZ3ca<85EbE@eScgJb?
WD]_a=O=.-S^6-(efOZ8;#:bIW&5gNGMed?[TP_cC+dC5(R>/,T9=ZW?]g):abe5
3P&:SM\,cZ#2J5JY]B-P>H5E)+e#[IS,<A&^Xa.Ie3b#G+;XC3))cE8fWOYV6I\-
MT+EN@A?M8:)U7Z6]D56>.)bKdd.5Hbf@&([,F[:IX>G5f6eP6-/AH?=g0L><R[S
<&aI5DaL>@\^d5CC\[OaR&#83\S,-1L7:(4KMY9b_@J_fU:MN:b^5&G?e<UdQWaW
G;<L\H.LeQGFf^N::QP)a#XLV52;D#)Q1>.\)Sf3P730R^0g3F7X2)8(?GSAf&XI
#3L&b\++eVFJ9-]G?&0/9GebI)0b:aSRI0K>Wb5T]J&X__B(bKC\ZAX:#>b9?8DC
6d@4OVe)(\&0ZV(JQJ/;\fE)6]c/b[8=AVI3I&>^=Q8]_7W2R?Dd2f))U&(K+FCY
K-YE[,eT@1L_6Yc9I+B:@3PXC1(PQIIU6d#7gL4(UC6INf_#KHO9@;g2W)(_&)HF
]U>c<WI:N3SZg]5O9LO2bEdUT;<2\^a9?;>:@WdYSBATL9=,f([L[\H(J&dR0E4g
[c+V,NR?082)_.L1R6\0(VKgaS0-T_VV1CXV5=1V&b^U<\d]G5UW/F8WEG(9+\2_
[;MFP5W[?,8N]cQ@e(^a>:>\Gg.Eac8_;FL#IY4Z2S:,ZFgG#<7=GP<:3^5ASM[;
-;4,bG)>J+A5.gBB[^c<3SPX\.M?)&>1V@4]T:,0H#5V+Ndcd2-&/@a^EXf7VB?G
.DLg_,N^+ZQcd??@XAD:^C@e-F<_\DKULBSU0W&5[P>EDDDT)Z\[2^U?S.0CRC&)
Y[c78964HP8L]D&&A,=GFMGI,fbX@:aZ>E.:aa]HWZ+;#[#DGG<Tg=@(EH]3cJ=1
Ma-[[[BHF?MaU)W:5?a.C18]+adcfa)IJ^,dTfSVJ.Y\OTXf@[JcGO5GP:\^YE.?
[dCZ)+)AVeZPD7KZ1@7dL#TMM6&Yd942Gd92dgUg7f<KN7WBL(YF,>8]/L@UL\Y:
Q0W+/]dfLg644H^]9D-?E(FXWP]Mg\[=Q(eV[KMK=>H\#Y@b&bJT@,(NH0GJ<GMU
[:AC1GV>Q>T;60PG-=,[LDJL/7GTCcLIDG0@KL4;)G),B_+##>0NRFW?+_<1Z3Q=
+7+XB:;)IM=4bOW4cC5;_b@eV)ODRYTF5K.R-@_6EV+cLOL.,#VN,1g(JR-(#O]_
G/Q7XgO=C2(F.cEF;<Wb1OOA\3<:IMEH?V;02U(Jc\0b^88>-f4.7R6JdHV@GP-d
^#_;5<O=Rb+17#Zf5^)_F9CGMNC:,TU7;#[WD7eKVQHWPfa@dPGL&V8aWCDKRcSH
-_T>:BX\dbS^Fe7D@2a49/Xc:6N?c1)bdC1O@&/4d0]60#a7)EEbbA[HCTERI<?M
JD?,0;MVS-@gfTJgBI<XQ(E]@8D#\(<:V=R&.2(cBa4B^T<>A\]RM\#(P,/fZSHM
ZfZLNNEJ0C&7#Z0B8d?]2ITOd.:+AHTTELdOQFLb)HU>9f;5=3[K4Bf35F-R]PD7
X63^FGYH0OG1Q1d\.ER<WL.SNTR/Neb05Q?g13Q,>;2H[LP2[1:8cPQHWH^V@^)2
D16fFW:b&P:9_)?MS(3Z__DR-I^QPD;YYN;(AI[D3D:/fZ7@81V2STCR>,;I(8]\
ZT)8VDg=dG;UTCM[;CB01g1^SBAIA(d.Vc4L1=9JG;S7D:2CKbAcF^G(-A=5fX\=
0,:[FM[D)\\5?:I036[B;;?8RR&H,XLC>W0bRDIb<3b_M,DeRX^.[2OS)]N(_LZF
XIM=EU#6M>XaR9.\0E6CPe,6R+)VgU:GHKB1@-E)KI-SQ/M<RQ\:=d]LP<aT5FKH
BQ([JN=1Gb7#-&8H8?2@38eV_b\g60[:SWWP3=X29:25[aYS(A]SBS0U#TJTO;B-
6+/MRA>a3fBX_0I/T,)?^@AV]d4;/T5H645dd><BN@5XUPfX.6<1@Z3IEP/a.(8H
@J&>#S/2?[0/MO+bZI&NCT<L_1P#,eSJJ=EM34_,(SC#\.e-3G.;b&Y\WR)J7N2:
XRRTHK&@S./aOV0?D@0I#dd97(X4#=8B5E:SVV1B1M<5J42XLJ7GH68f,@UAGgCc
=Q<.^]@LF96(C)d5=DDF>PLF1W3[IF4#5[\5MgPO,&0WE7f25(E60PQ<[9gc-0G=
1DV7#a=/Z-c94LN[.cP/X]0P=ZI#@[,<>&Y)JK=AP:8=-\Cb;5Zd,HEOHUf6ITZO
FU6gWPg4gb1O09_7EN_cbOQ/HHZ=gKNZ<3EQ>YLC\Y>?\&X?C6:.2[41E=d;3fQd
UC\JbR+I/M:<;J7@71QdCdG99_^=.);[WL.=[e3@?5B(0F+(?]2UQ8-SADe_)RdP
Fg59Z9aHgbK:R(BHbA[e6D#MAa>,5=fTg903X1-461^ZCNdJUG9-K<E(2-VLd(6V
H?AYVEd;A:UJ9aTWgANR]<G\<92B[E8GU=@OV^.<fDf0[I:T_6LT3aHae]J4:1[c
T0W3IJPcSJ?0J4GQ[U)RZ2^^BOU:]7]BZ&:F_Q:CMFUZ^[W-UC=OMJF)^HB5VSJ/
I;96J]HTG,;U&ZQ.C&LF8Zbc+Q>DKg;9;2Y=Z&C&QRc]AVF+OBS3=[-F:O-E:PX&
&D3Z0#\12;\(Z#\E:QZ5-306ggW?S:Ycde1&aN2:5])AY4+#YQ4L34TeGP6-/]-\
V#\ND63a_?^EC6VB\b_VONLOd@Z)[6JbAg&F(FCNK&O5^)Vb7_DC89ET?.SLOVVX
b82,d.TDgA+GOdNYG(MPWTBR=@4VH,:4NfYRATXCKPT9E3[@ZG8+HHWP<+LO>E[^
WYVQ4XdT/cf.d2YC]\V204:(\fD+\1>X\ENOID5B5aCb)0He2A0]Z3_9JPc;+XC)
DGXIb9^b(=YC3dN1NN2cD+^IZ/3bYYLecH<,>5KSS/#TSVELYUbd7N;+YWIL+YO,
>?AC1\T5Pf<8@S]7^I-NB>;(UZ-+X);JI;#BDJJ<@#?33WRO#a2(;]WN_Ff>H,RC
A.DNLS>F>SY(82f<LN1/Db(&_^:J63+6\2PI?S8+10DIb_S,)OC/T&R0^@8b_7Zd
gHTaaD8GD=OD)NLc]eLb=1[\2DRN68.;8+M@0J9gVd9aHd27C&P/<_aSCT3g1N@W
cIM/Wa?W^dNe3^.>6E.?62f>-@F(KQ-R,f8a^T[bCdN4)))6WVGY(.a\eVU)FXCY
)(eQg0,\RD<<R.D=@Xdf:+NQdPKG2_ca,7ag)EbS@97JCD0<=>\&?K>\G5HDR+&c
WfgNS&Ea/L:6N,#XJ]aM[UH)d(<bS]\@H-D;768V9?N=>AM^,#/f.65?bI-C,TXb
-Q5f.Vg<F-D#CCZd7FGfPbFQU,DKg4Q+1.HG],3_JT-R^7KdXQVM_FB0XENZ^83b
YK>:0Z__BK;C=b,:,_]f&d/f8RT=],:I^9AcG\MbB2S4&cVP6g#XZ98K^Kc+1=c&
A[HK&g=O_8J.]FIK.,[3X64@QXd,dNcPXCeDg:FEQPHQ@C#[5B+<32+:(-b4d>#?
G\Y>S]G1&.WU#/<1:g@9S#6IWYT7JbIVV8#7VdX#a(-()15La<8@07g&C^-BG[@M
\.7/C8L[O,bU-##cTDD;IK]+]7QS)\WM_:5Kb_951@EYXd@f7JIOQT)60DVX,.c3
F0H^A&bPL@_e2O2a062b52127]=5T4Pg?J/F\d7+Q;>8SQ9YE=YK0:P0IePd]3=C
XX^,<MGY27:EM2WDQFMC1Qdea:cFJ_]MUeX3.,?SU^T]EJb)P+V-4VEU@-fW.-.)
\]g^;=X=)E=8aE-gfL&\29;BYNeYg&79\Ye1SJ9I&S:D]45+-C1XR50C8G3Be:6e
0;abR:-UCa0:X82Y@1QY^.VLYQS]5WVLL(3a-80T:>Nb:9IQ-S2UEPYZI:UTB(R2
>(YJ0F9@-P[II1.7#:UF#I(RHf^9PA(KSW\_2Q68cHL-a\<U\N/dTLL&,@4_CC15
aDZMJ=P<4B_?c7aD2[.)((2:G\C-VQ19a5Y#]A<3IPO50]TF:P_=.CSb95ZBeXb6
OB5,[_Xd//V)/1@ef0O?6NSg9(1fc;cc-9WF4f\LJVP7GDc#6JQCcB>68#EW\.cF
OSP.KcT;#<YMC,WaWe.cIK\X:Y;H&c@H<JfCN?IYF_c8M\TH]S3K[7Y<@<FOX6g[
X+Z@+W8MK9DHe87c7EIEQ..Ma-,82&5?M(6A^cCb7@a-D,U1T@OG7eTgDWJFB/@D
@CcSMEEc6LB8+ID43^V21GK(c^TSM^T(WI)SVZc[7.:75)4H,@;aS50)T78+:OD3
M>+;eP7?b(9LMXAZ,)=fd54S_3&D.==1PB6>R.T<SYf:;#^+56a^O0S.GC;d,(BR
/WWYf[F1G]fMQ([VKW\@(?^LFJ:(2RP8-.HL),?>/dUV<OEA??,RC]FG0QLTNJ6)
_HLB.PAYb,150UGYEPBRf6JA1Tf:OJaQIFK&bc)<DLXa[^I^K0::I_SBC6?>@Q0,
GT>FP^K)2Z=7ZNO8&IAO3=a9?ELY4/_7[50[ENIW9XB;f;2PIL(WJC#LQ?.DVN>P
]TWJ4[>4@[RIFGB2C?Q^>V[X1aEW&Ja3;&3VDDH#/ENHO,a(NTD>f.#P<(g10.6c
8>,dL;&a[S?<K<<S4H[bPD;7@AD2Ga;[e#(RZWAg6X/4<Ba#G?],X;_NMWaNgeRQ
:#GB.P_E:6/b^4Jg3-6F3KT.27L(a+CfMT<e_AX#HOAgJNd.Z(Ke<F\aPbYF<\:3
Z+#F5bc64CGXV1@SYS@CZ1Q7?0/b48SDVP2UC34R3-6<fNc,2\O.6<LS.^+Q/N/&
<CQ,H]_YOLXSU25RC=e9B3b3O<6ZXWdQY1L)1FN[@BbbcAR>]L@Y)UU;BY1@54D(
^]gb8S7L(aK#P-,.)[,M7JQIJ#_I8d7D5/^[=<Z#fZ(_a89D-?Jed5K?g108V26[
1G.?g,MbY9KN1_?]DJXW_aWa6ITDD)QgTd#UFA_21ZD+.?85>DN61]VJR+0QacQe
RKO&7^DJ\f8K</IeLS@+HC]B)cZ:U5@^1W_@\:64OH1V/68dFb/b,D+4=)7b0[gG
]+J/Va71<]7<(7Pb7=QefC[2SQ&WX(6]?DCO>V&2\>^YP#>c9RM\R?90)8R[];8\
F-G9,G(fZ_69aVBL?^WHY69W\cRC\6D77cI>O]FDAE1bd?28eOQQ]>Xc512#c55#
SJKML6<dD&2N6,IUDR,]/.G6PJ(=D&6O-+__LZ<>Y9QCR<&HKQ63PcS#AL.CPT(T
1[0FWR&GJ]-IH3M\;KP@S=MI=M6a4Hf6<<bJAEWKM=+5WN6&?3U1^_TV[8A&PLAG
QMfERT3@cB@[;P9\+^:9J]NK?/\UdM=bH:IOI.]HG-RWHTM]9#S8-)J_YRYA2IU0
[9CAU)d#g4fGA4IR2f&9OP_#K,4-g(eTa3RCV.+&O<R7d]]<7L6@?[GfG(RcCU2b
55WMH?P.5Z?F<?<OE=]A^:e.014PS.:DbP(IRXAFA97cX<IXIe-4TdAFcMM>8dR=
.bb^<;CLCUed/ff(V5JLN_XORfdG7]OP5A-N3P/8=BBgc=Ee?BBEeAR@7>.Rg=b[
BF<1J@]WK#g1RY45<aX;PA)C>0Q,Oec0gOP(EdZ9cQ==O&Z/SCLH1/V-H@0ZUAXA
WC/10g?HHb5cd9;T(G/YW22(1\gEV<Q<3A&Lbg=.M2YW49E(F5X]\HK+<0B>.Y_/
H^EG6<8O>:R?/XE1&F^1@S#AQMC49_;\9#MbKIP(/J_]S,;=g;&#AP?LI8<2KJ<(
<^5<@?E(\1O&+:#>AG6EEN/]IDF3=&[U<7.3NZ/VB797@F4_NC12f-=+KFRZKcSM
H,?MM]Q1>[P&O#BFg?,Ic_#07d>gP5SDSMH-(@060)J.]W&CS7\:U6IRSe]cb=&K
d?H6c@F)BGY5JX+M4-SE2_EYHTK0_8>.HX3Wc@AF5A6;:aJV0?^HIG7/V\-.Pb\1
4,=CcJ:+)/\EV)3CcG?DEM+]Cg><LK)TJRN0:ANU&VV>;[#Va9P60LV]ZINV&KfF
db5c6?HCX[><T3NUf7ga+2+cFDecEP#+@b?491dO\2&,cN;P=0PWGBWRS2aE2;:a
=#.9_>@JJ4P=5)U74Q\T6G>d-,?]AKT\G1E6@PD3:?;WAbc5)I>S4Eb>^N<>ED\[
PLB\\5&HFf<-+I(RQ)f8]BR,b/0K\<LOM2K?bPfScO?G:T<@T46TdRe2(W13ONDL
Z&XU<0W=B;aN-eVISIKVLUK3g5IC\06=42Hf4BNFE8:ZRHCH3==(Y61OcM_XdSH8
4d)Z)O=Rf&4g0-cCL,TZ=P^a1O.,BPIF#0aS8SQ?M\.[60N[I]A99DQX,D1FB8I9
bN\_L_XZ8NKfTE[[HBFCL)Q+^BG&b9F^Y-VW,eE@I()dVFOafK:.cgATARc/9J4B
[AXSWb8#XQE(B#.\;Q2UNga4Oe#>UN2f&8\8>C^MP#9,A8bE?.c/Q3@CR8I.]GcP
4L:;U76&9.E4d2G.DF/,aVZA4MGGaJac8Y/YWNDa::9HCVbNM#;=X-QD<+[Z@D-)
?BK+]Sc9Q(Z;c1L5g_dBTM4,eR:>)FRQT\:/aTCLSV,N.3bQ^ZWH=?8Dd]-0RND=
_=;WU+\\P1;5:&55/K=)HVO01a/:KTX69>8SX+R]gM,MNXDO+QH2?Q]N(#e5EJE,
[9I?.V:;)\fgXed6ZU=g>BAaWNW_H\U3R(S_((ca7d:ZS3dW<TPB1EbDK(8R<IB9
S+I3H)XF8#X,Y#0V3B9.QbBg@aID@X00QBVZ0UJ[_-dQA6>,YC^FY_5Mg9<X7X@>
Y3)g(8USB&+V-Zg2..EcefG9)@U9e]a])0TbD[N9=D\eN2eOD)QAIQ6ZQV4_,d(c
?LC7G11KQ(2]>)d/f<)bO;BQGWU1WM>UDV]^?^Ed1#I0JP1C7b6\QOGYD+)EJR\#
b>S?29C??fcONd0ZV]Adb:Y-@#KR-9/CQNTa+)?NLQ:?NL(=^2fXK_8ccN;0-fF&
<gFI9/>CV<Ha7]54PU_,1SJJE/&dSY=H?+5TcAD@84Y990cBcd?Jcd1>K8YK=,Qf
A.bDNV#NV;)=-:-#ELabUFDX)10N;>KU-I#K;7,(OG=Lg5SJYB(S@T)#PbHg=:)8
]Cc-1O<VP(EaPJS8Kd:A(.3_N4dC-KHIQESd,2?C^2IL4C5C8)H<gc)fPK3:_7EH
?^>&VHQREZ;8-6KF/R5J_E2K3:KCPXRbg+7Dc.US]d4fD,d)9Ob6HW>6De)<f?Q?
4B.c_R?6+]e9=51W8C<M3L@LIB1S8?.FFd8YZ+Da#fIW4ad;3+#IGX:cBM/K+-5K
Xf>4.&]e/(7.OB6K9fH)a(/1_&,gJ;&f^0d=.H5\9HL-Q?;H\11f4&P/AV6HB;LS
QBN7R(N2BG3O4Q?35)N#^W5LTBL1WR4Z1^M4&-PP(R\?ZN=/6:aF5UXC6<#6<Y1W
JU_A:>]@V9_fBAe9O+bZI7KE_MSaeVA@T)1SNT\3?L9]Cce]G&KVBECF<]P2C60B
[J2#:OH]4b\:)QCCB2[Q\U^Ne;S/#LK-Y=]#U\T:I-=-BK+]PB8cGNDCPC6B1G0)
\S(J.J2aB#)HG)M.@feg;YEaM@[5beSZ)g5()Vf@X<:V/6/+37LQ=99404/f0<J6
4g_61WS^V/7M[426M@:)>.)S.]H0Y>cW<REF(+M>d0ZL5FVO71D3BeZBI92=B66X
0_8H:=\)fSbHTc][\AV<5]N[;G@aW1PF[OZ:a58ZM&V\6M@JV[29Q4)g0<PB<PGA
Nc-g.[Q&5Z_^eQHPP7U-AMg:G2ZW^2/KS/,^g+.MT#4)W>QHC::cND]9,>2;?C_A
]5>&+S#H,F4LOEU0fZ92e9f[A##9/#AgHUNPZUQ>9YL40[&LE&Ef;DEB]6&+S2Z4
,I.\.W0CGHW[gCg5R3gA2<IFcJPAPMgX6=Q+#1Z7?33]V\Ec)gM-X-UQKF6-4>0]U$
`endprotected


`endif //GUARD_SVT_AHB_TLM_GP_SEQUENCE_COLLECTION_SV
