
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
jluANltau1xFmF+t5SeRyUGK9tRVjigze5Y1qeK0eiKfn+ImqUzgvPjXeH5u6axK
6f7Ntkj7lwduETDdUjdHo4TsKtfN+UDT4fH3bNQeBwX5gwXyT8UbMrM5k1Dv2tde
C2Cfh4eQaLbeWoRK/KLj4ijzxLW5pN5pBKWk8+1Bx2U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 549       )
vQgwme3hrIRpgIMQH0+g0ZqwaKaP/jxmYNsPmKa308PwYbkDqhOIn09Ww8MGX35w
UddUxelg/8x/0arnD1Gxp72HEYbHMiSPy/o4gB7i7HEEx6LY2qCPT1K9ljrWIe7z
eIc2QKX/UHzqZieooVvavFYcRyFeJyaBKCuAWRAcogGZc3RjKHYbalpj4kkLsGBZ
+57tvxtfdEkAlgTUT9LZDFYGOFqGkdJQ4JtQp0aTTb+4Q3lfVoKsm9OobvNrsWW+
uBKHSv0AZIg6fk61kuWtrIMvU9dFAn4jWpPQvziiRVLzSsK4cBttRSOwZd8bu2uB
QnyNzhtDZ4xhRmPbRQMmS/SWuV/r6TJWmmc0veighPs7SF7O0WNuMb5HpjvaHX81
OoDzNwbtKHKRHK9bas2of/TMNaVK7Wm2tguvHpRHHQ0tMDNjdOcyHaq8WzxA3hZ/
kVybcPvxl68aCe5P4oEEknMu2/IcJL+cmEJRCYGXY0GmhLwReZe8j26Vozzg7YQr
8UR7iIsN9hDWrRObY3zcksU7+PMPW+l7uW40OE/InkK5p9IqXPFFNZcpG7X8UfTs
sacZKMZk69Iy6SVOmFDSc8H3A0aoBWK7XWOQCt2XDuPuTtQAynwKEjC5PO7gAuJt
hhgqhrJaG6V/TBruVPvxCwv23zWNvzAs60EGlrDkUSSs4GRAR+UO8YyT3FrFEYhz
1Sf7bAs6KrU1U4KkGvhewHFIbDcgBw0+UyGzBnLy82M=
`pragma protect end_protected
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
eR7I0z0rEST7wjyReSjdTnzTo689f16feUzcuhikF1Q6GiEbQnpHDQByCCYHZqGJ
yTihMc4//RnhMtxAQXbWm13DHrovCN3EXoyR2vQ45gptw0EqYn8E+Epa36aWpquT
1m8pdAwNNuqCe+STDHuCWLPL7DWTJWat7KbFVMtaNxE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 789       )
7y5TL5Jg+emiAxkisx+BLripIIwr/+h/kwq4XHALZqFzJqbeRdIz2JZ1bRKESq10
9+buHXKPrSuNoUUijc74kgpOUYxQEDpgkCdpQm/LdJb/0MaondQSRRWnoztd/sE9
eSNiKbeBPeMZGPK+D5cTjvBRQEwGmFoBrxpwQ7q56apTxYQ47uDmSbtS+43JvkSg
EmbjWNQW2FFCfFM63C6YPVS7v6s4ueeVEmlLhfxW8dqLToMkL79gnWWZKHKwS/qP
AIjUXe3QAqcusTSq0aP4fRrr/ys83QV6sm92vET2wEIr5N0JT2nVHQh4dnY5jdW3
kpqgvxvtHRcQx365/0Ubeg==
`pragma protect end_protected

endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
UT+b9o36UH5DbrxiSJT7aKf7o1lBhDXJ6FIdIlExDO8WLTiGpbVOfRDmUmHiJtYP
t6BIvmgaQt23UOl4RBcvQm1LP6kNcI97hIyvXnDCOodJMytszUp93Z/Ep03XxTgD
/uZp0eJ/kfVV2E/YGPXTupHTStDWvya4/7gzMH6LjW8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 1256      )
YTomvzuIqt6GNbUeF3Gj5sYet35h3K6OeerBmfOs2A3Y8mimtnKVN41a336+Lm5U
gCDMVtTtpk0sT0gGeWTBa5Xcx7f/mzfku+tqGLDSdMHR9CUHxf89AtsxygJYSVVz
QtrK+S4yT7H82xh+s9+JgcIx9AQyB+HJ2NMFDUTK1jCKB96fyH8+G0IhESzSNzJ0
TAd6TBD6yzrn/G7SB1m5TYP58rWUMJNpBkSB9J4ov1+1sqceQYDHG/2D3qfFl0hm
FFR03zBb1H530hm1YG080iifbVsWdrtuVBsEKBAGzZvSpvzTm9Z2KdhuN+hrtl0M
qwd3Vx39LdAl5dT4sKh/QDbHC11MjUJ6fAk3DGaBcsCgr5cF8ARmVszv0OVriHU2
59V1Ls7Eh9cs0uklRQnOGZY86/hDuNPib1cvyXqzwnNM9JXEg/7W2TcBaB4xiRER
RSC8bqaW1ry2Rc10K12bfU6ZH1t0kasTa1i/QDon373tmzYfCOM265wO9GJNv6LD
zk/oGsVXdZIbiG9MNXns4USfS3Dk5FQ6Zkz/pej7dz4AZNVVaAjydsOrVH1cDm28
Xu0fQX2dxjqYtoHS/jz1r0nLZgbnZw/p5T7xMqs9To3XXW0Hswpfdf3AzOnQ3Cif
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
gYxridb1GZfgN1cJ2mFhvo5sv9Toi3AW5tUE4dr8lSpPOi0SyH8xLFM+WiijUK/n
zl51aU+2TwBSDiaxIyuq8al3kj9vEca+hoYr7p2Tg75jl7emW70lter9BKv8BHmV
RD5JEv68RYhxaqyyKcjt0NYNded+3rYskU4qAHDX+aM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 25280     )
i2R4+jSos9virCUPjNN1E2gtdSbmotRE7LTMEr+1lRoQGNyrmiuYiuszBvRPqwAU
uvN6hv2oPPhZMWBtqBWSerhhQmFtFCmIY7Wy+jn1nwy1344iDdcqjGAqBS+tKEoo
GAd2Wkxs2h3VPmLxs5Q5KUZmnjWYKI8po1+ZX8Lg07lKVvjRTvqH8BaOApR2+4sg
TX8XNZHNKfRLX35/uIegToLnpmGZ3uRNL80rVy+ON0D/6QB06obaD3QkLdSzixmK
jqRrogb1IAhZBJ53ks23IwNv4UVJlyYd6DBztXSD6ZI3iyANuX8CSUSvNHgcZYvC
JYvIEDVIV5xLeKsT/uZc2vH6s3mwQZeNmCHWKdg1seq5ThzKJ6f6aKRwDu+e84ck
XGkIOEpNG3Tn0uedc38E8S130vhcpHcDR16AwFeK35W8k/hRsXtQxsNygjonurHV
6d1TN1DgjTk9XVp3F4Ku3dvafiV+o3MqEH2pfUUYniaM60OxmzbBCCs2xTwgKylq
G0mXVeoeoss1nOPmMz3/0b9NbHf969GMLlKMn2P1MFWnsUy1teN4QKTS9OI+x46T
yR+JIoGGaobzzQN/kryZj4jKpWWwL7phvCq0D+MGuJ0aWAc2YpmTdSUwj/NgR+Zm
kNVjiJlQoZwjZN+lJrrR9cmaUp3ctp0Msk8cnZXaMA2/DBlrjMruqR0BpKXEItXd
JqE9EqL/bVU1wd6Hd2SU8z7codpqFAU1wvI7fpSZforwJgOEAvVJGI+Vsc6kdUIk
5vzoeROc+OYhFQc91cjmY+pgSBKwHOX56octd2pwFD6Nd0L8KkHmSozmFePdx8En
yXMlYGUQycdVUIk/Qz7E2BRTeeJdzc+bnqYNt5dFpUZTAqNyAr3hTxTJEeznl30V
jnYpMWDkyRoSFta1FwVo3YxBbA1x390Szo56hWhazNewQjzKdeSQWs7XOBYCAaMI
014caZSDm7vxRyxnNYBgRn54CRCE9mzMNISUGqZcm0kUZqfzgR1YCHgFvu6L0D0n
XofY0tBIRa5FfaRZbGkH7cwkMxTanNhbrckM4l6yGdj4oTd75TCfk2+onae/mlRo
ITmJ2M9W+hTzgRqCd57p9IDJbunFYZpUDhg30DDZpMbiPuLwIX4abjremzuiwVVY
ZfYiqmh98USzFHfMEPuUHBYwJAWsH57PjIEK3N6QHc8JsmsVSJpF2EmuGd0TcAcG
mOM0kYF5u5+A9+aBzNbqJ2+a00CwcHIbYZyJNKXrGlT3AQcnaPPllLZ5CeuT3B/s
0Ig6cKNzruQoh/rfbvDH9hjvMspMO/icIw17s3Eq3WhD7U2dGEKTCTEzirrBdwv4
k3HZrVc+wm4RGl+Djq1Bjsn63QJour+5IbTe3cGYQ9ANcldUeLqK57gYw4vN3lyo
hYZYX28AzEAStMPGHbIskoto/J3M9x0hR5WANqoit1jXARg4mnaXfFYtJVMTiYDR
ftvhRmJIP7hIXzvb5ersvnooO3jbmI4K4s6di1D29MK4E36BGswSqeGeIQ0Xt1oi
MxoPj7xw0M0n+VCUBx2GYRUg+8q3CXJMR0DYXwFaCNju51HaY/ciHyC9i3UIoj3b
SH1ZSZ887d2iOgIdEzAkTD3vjYhyNddrvi2xvcpVEtbGX0Y890w9/anyYWbfRObv
ZT661Q6ixLaaHDUxKZmXzvd8Bznh5Pcf73UYEvGkcd9Fqd1jhWIaSBqzxE0kG+uC
x/2lx1uON0BEuXYqq6/YhitmAtsRHkctReB9/Y1GRgmEfakvbhQ78sq2VZWRYenN
Hw94GrztMCJomwlAGkqujR2E2Gcqhw5CkF2mxT1hPUoaUKC0iZrRbuAIUirhbov5
v8f86k93JLSTNHyHS7NHA3/in+TqJIDBO7KGhuqGnT5nA8TstZ8Cmw290BIqSvwt
Nbcwn2AWqJQM/d9guUhFin1EYtBW7wLTDUOSOWSP2pkpEWset7x7ADptpzDwsn82
9xAulTD9wV5U32+w9QyXFFlNTtDNKQIdjiP0JeCYBiBm8wIKbHzOew9DOM7y1SMm
gFfU1dYQ34PzC1yXQiUutev8lcpYSRqp4cNP1QEb2ClNPGpjxxxIOZa4d1wKvKSo
XLdeZiOWt2I+/zlfrVDdap7X+DHbTaUdrGHprgN6XAb0DiNcPJPPCZ0lYM1ihpmT
zzVZqN8I58A9LnkbK4I8gF7s6pESFBJjAty/G6BDkg3jgQrLkASDrqhGlwSkmA1f
+L0QbJLKTIUb3+zo+MtAE/kjLbstCBxE9Xe+xRptO+Usx5kVNzwhUixUXlBEUGgR
62YP34bXY5Cru/9EkRVPPMEI9DGOsAbWDvP2+9Ym7HT12gbFos3J+MVYc6MuIWTK
J6ZO45vHfuQTyEul4w7hw6z8gkmTVsgADnkr7eoSYCArZU4A5GCN7IpzsRMtk121
5NrDCtvUiIIbo63+x8ohSfC30usm3Gl34hTlq4Pdgvb1L3bfwnHvmbGufU2/SMw5
TZx88lV/TWznqLQhCeJ4y+txNFAAlc3XH6fdwolfHiRWV6Xjh2V5g0g8rDWwXU9t
a5sF55dD6wsWycgRRaXxms18CUSrkvwzA8B7ZvGqNIP/HqjaBLc0Wq4DDpjsWoDF
1KdoraO74GzP/10Twg2vvezryFDJ+kfl1DqKPU5/VD5yVcXmMA/fbPimuwZze+IF
IO+EJoBj5R4iwyt++lAP4NQ/ndoryVg4NrzJHPkplZ3JpmUpWhASUSpoi4zb8sKE
CtqEBqoQAAQpd+GB1WGXzUM6Ngl7bf6iXlk/qHOTkN9v+F+6mcsgRJfwD8fuUixV
wUuODc8dg7maxCYXv5TpJiPfQDLCiKvzyrbY3V6qq9T9W/ulzp7qsfJlMzVMXqsT
AcQ4afecKb6JmCVHBOxfgvTMNc5kdHiPnTXlYWfu3bpgiwF+L1U2WaxZMDBN5tHc
b6ur2O0NMFyCmpqBj1qviPf7gD4CKByzBk/K7h68CHwRxjknF/aqoyx5s653KBQD
adMZjBJ7o8oh1foLdO6LfDPcRviKwsA6N3+a/ab1D2sQwL39mwkE7hlTGghzf8xj
E0IC1vCMLRACG2naS7X7myMrjyQW98RpfMcT2sutn55sgGxjAdiJYaNx+iH/H95S
3CoSIS2fIAjeOMWyGGwJ7eC3x/esKwaCAtIe6o8UyLhVapm3BmGo10NYHtGmOX04
5a/WXtDmboAAit7YqjMiJyl6VOFqj3L8cDJewSg5VfF2L47/pg7KJ2LnzW2u08ga
4UfHvFWfZPPQGaJxMbzQnkheAK7Y2HIqusgmerssjV2MToBDfQfmYy1Y6cVv2gui
uICevvH5c0z3rofRnCUlTSBxNaBzciJT5p29NIi8EWuEYi7OibwsVbD+RbptrgA1
y9BVMgtEIyM7X+Ijx4QtMvNBE3M9YMUMw5hpXQkvIhKBYXyJR8IuseJowVndljqN
zt/U8T1hr7W4U0GLZZkLEUgF0brLh/RYignLEviFpKpUlloh6WGOa5NceiSKW8Dw
qNrN/8wKfEEZqrQYyH+0hGllUXn2OcMNtO73pvm2nEOEnX0rWcYgasvdNJkkWd/p
MKe8MNxHKjmeuFdZag+WsfGU1qAg7cWDkXCc2nOO3vHSSYdlD9d6ipnWjnFa88Y5
RxqqKFOqVR0c9H0wO134lW01/XHMpWbsKdltjzVUCrjTJiZ9sGPcRkXkoG1nK09w
BeaPcZTiiou3/DFBd5fOJNt8ltnODcxL//c0Va1FoZn29WRJUOe2UjvnYYZNyUac
bjbS4cybUsSrRAVJ3Wv8yY7O4i9K6Gs9rDpMmkh+1lyZbLItQL3q+cunEgnO3R4y
pczxcSM4L/4fnjZGMJPM54v4xT/swzz75v6BdPb2DYh2g10ywloOPROwthIGqDW9
o15qxdeS6X7rC1YiRS5fTqH4+UBUR/6rbsEuaOgyZ+3B0QBNvzYaGUSlegWk9QrE
MyORLzZiiizRzmj/9S+Uq/pLDrsqa1XBMmYTs23E1Tm2jbXZd4mCorh5Fi6Wt3Lb
R5Nd5P5h1DwfrEfBbITW+lAUfHbWUr+QAGURfwpOkzvOtfFlizO2SemZ1ygcfT9W
OJf/dc5nWLPQsdyuMz1gD4+QBYVCO8Waj/zcPee+N3ZVHD2iNWUSuLkGka97NTF3
G/oatd3X8y/jRVbev1M4ShbCgSOFb96FVHbuoF0X06pcteDlUKRiOMg5KJASbCxk
EEs9Oqm9tPKpe6lrsqnmW11l0r5CRhBnZdDvxYcTt4wtYPCPRmaPdyvEcs58SpFV
9JGfbGh/sYfTUUzM8m5EBi+/NTjwIvdrg0/iknU/1D80hRIV9DY5/bIVnFvzjvCk
S9wpKbjf845rmLFNbqLs++xiOg9g8o5YzlEBwfYMhWhhHCfUeuM+BzGHxJe55KjN
76ZdCTiAXORIuNUMr9vvIqTTcumeeFW/FwNhS7hefJ4wIYgXtxpKYnFTECR94PtD
pGRalgM87pkwdL+dooJNiFQs7tyDCqGXO/nppKzMRWWyvXCdbaghTUehSBVPQH+a
iWZ30s/MBicjVpuvtRKPAAffM9Sa7wAx+osLKcTQ1w67sZHOQjEZ5vyPyH47GjRX
psaUPIwFKiLPReNOJhKvW1wjgtrpazbybATkptzcZqtGmKuF90IqCeC6hhmbCxNB
KcBP76czJ4qnEDFwL6j9PUEt+eFAcUx3C1imRwU79Eqfov593n+OYwj3eakoc2LQ
ELULap2OyD0+323VjN9oznHTU/i1FbnfwiyKUtuARjsR1gLjPk/Q/qwB+5A383by
yTRDSwoG510oHi/C85Ujw1nmu1FJ1Vsy+nU96HVOlS14jaNCgqB437p0zLLerJu5
KSZm5fLjCyc+Wf/707S12ct8rB1UuTmyS69/RO7HE5QHP425u1LNjBv/tGfziyDj
TW7M5cyKmKiMZBpWwDfy2EZgFlwazhXJyWhcchYYOfWFAWhH4DqNqRsOMlJ2qMfp
Wp+gO/c1BbBXN92bt1G3JpV6L+OUAr36HjSSOCyElUn6eRsOOSntJsubpln7J61G
ZSh/xSrh2wX1vUoYEgyMo4rNkC8PPrZxcT7PlxjGQr/ctXYnnfWIblObKXVA9V/r
KryvaUmPCaTIbB7VBAusAz3SW/EJc12Je7Uhp6Uz1loMvLO3zhmzUFi+uHRZ4bWL
wdfEeTLo5t9Ud4UqYdjZ8NlFGUwqGALUPq8W2hb/0wbhC/KSCQQxuiMR0Z4+Im8M
GzQxDP+j1eAKTVwUa9dxFOjY2ZkGmxf6sr1kSPEHHqy1GWVPWftrd4Fg29UHMhXu
RtK6HyAx+CdPgJ3Un4aa7S6nNF6tycEZ4w8VW9fw57o/BLmCGKCZyl3rRARqFJgR
SZJiM/PPPsOOmWZGjznuDNDfARRM8rxtdoMiQae2/vcyp1LCDrBR7Q6ARNhPVKo+
KlekqW6u0A5I1tzpS6BtLGIREdfn70Hk5SW/MXtVzSpZQuQcV7Ln9QT+GXEanTLp
Hlog9fv+KmRVIDAXG8zfcPGyb7MZJrY2BTlOafR0h/eLRdPEMhbuB+/TF61Vl85N
f/OiyhvM7NbDA8sAGLda/ubb6VrmKlFb5w/rpti7xutbCocXrMiddIl34y5DwWQg
lRluuBhlWllKCW7jZtX7n2XICwo1Z215efgb8uBs9kywIe3LIHIFuYw+6IIMyL2O
8lCm5vErsIb2Q02fl88bxD85B7YKsWnWQC8ZQMhgX85Mtf0F9IwAlASwQrvb4v1r
iAlWLlXPb0VJNMfO0MV7nvpgK1qlQZzZZFPR7cAoP6EOQa+RQW8Hz/9Ljg06hGsY
56FuTIK8S+8M43IEvnWk7XKcPJ3D4iGYzidDGSI27eElaOzJupdKTfPyTXv5zXww
ppp8Xs4u+hl35Qov/Z7Bdp48jTDbTqzDsfGDSTVExaCPJVfxMiR1U2ul9fTFsEIw
Ukv/CLC4bA57yKpuK3uPA25iZX6dKVIf2UECUfGe1jbqIIBXewH/IrPS/HDpvzJ0
FEPjKiNAf6SgDuqQ+S/Zx32d6sSgX6LHTLzBGzBRxmFm0uGRZjT7wTGBPZc/pUvt
GJ20oVyDDqiJVhQDtmiL9e2yoIJLZjz4YlFcHxPv7CQheQC92i7QaMAuK0ENG0va
R0DrrHz+Xq0pCttY8P139YYxwa/Q7kmph312X1THOZaBA4f8266nor59C5MHcgrD
7Tk+5lu/LHlmT3lt8UIuboK8Dl8xAUHl+RWa+wPDfZrkuCinyGgGF21d2NaWMcti
cnvJXvFBPCTzTRiDwDRDTs/DLw/6mxejIac2bmmER2J+Cv9XIjHbCTjxEECsQGfA
neG3C5laryXEwrSLHGDeypf6j8+HQ4XLdLTWvF8iPZvuf/BbgNakAUGJRmKNcCVo
flZ2Qmi9OTKGg9xRqgSDrXUgYNb1n/vSC1lTSBxXIRImRfv+1a4XGt7TtbKpKXXf
5GDatnm8Ac6S1U/QDF25BQ4faXDYxmRKyU6b6ye0cB1qW7sc9thdy50iwouYcNT9
7GWxAyVtGpXpEusaREhHPwXPIQ70oY/EKbb4ksHhCleKp2MjxocN+fYhndYpNtsS
/xXYClnh4tYhOKdqvEVUbQhnNXoW72YncAKLZwn345IXxpADnCTihqEJa4WrmVPl
CCn1CkoZ42JP49cAYMWQAa0v4OpICDsW5Ta6Ok3RfHFTm99AaKvI06qQpyoaEEIl
gew06JNDn8iEOr5TTxx3V2+euc+iz7LQ5JqfZogyYgnRsb3lst0GUeS2xuyDJogJ
5BmV5xJOjS2qqVaUGoA46Xe19m87qSCSgsqVQCDVKKkFk61PWyU02xa/z/3352TN
j9iMsItn4rUMT9K1MMddcclNxW11flTcatUdDGn8A9I8r7c/1VJUdhbJKSZCY82q
ktjbq4EyJr+ETuLt1gSb+XeSeIFURtWO02d17oFW8ygz0YC/tDqkocRIDfcdAW/F
zzoZNz73FNKUMC1IoAh33v8I5M2kBZquO3QdYPesDdkedz/IohFaeWZ/qkBH3FLX
7jpy4plP7mEAi/4/2URSInSEcrqwR0TV7sZ1iCEjiNHyAKSVL/B63s29FUqWEhyV
Na8bxG+htZspkTVh+q0hc3pMaf45mUsd+YhI0NBGd0iESYjo9e1iWHgYY/kX8ll7
IKGpTYmH+xrY90hbVfMXdMzGE9JstFHRWRfTrsksTvtZnDDtmmgGZaX69xgeJ5rq
iLQbgWx19TPgbXYSuX4T4iWH2jYnTKKcrBHz/BqGWaHc9AunGF5u0drSgCo6ygdb
YFBEPnJmAdGEwVboRnxjFHJYiH2GuzEUjd7lqPwwjHdsprdbCxfnjZAfQOeXePz/
Y1vD/nfQNNX55HrnvHv4zEaLtgt7LQRuLTRSre4uwM81l6cGWcYp29DwBDZ3ppjL
FQdg7Kw5SQSLrLd10/S3L+aFRRmsbv/a7wVbT+Xnpi7fxr4J1QZoIZuok/J9puOq
ILU6udOzc80nJCYiFYjv2pW3AaGbtHG5ta/SdibnBQhnpwtYW6jEF8V+vfQpoZ1J
iY8paUolh5v+dtqQHMwyGbjd6SiNCfYKb5XUrBoy8bM/16EHMgHtLGuC/7qpFv48
lsPMSRcfixaWmNyYRSvXOTiSEVI+KG2zSfE35amWIvtPmZ7HlPkPVGpn79tvOjaa
krSiVhD3+53gr6R20y8rao0QGWsMmgAVpSTnMmLEsM8Tagx1OVPgnZyLxuJwRTLC
6PMgIchbhcR0gc4cDUa0JIsoiSakfDzWnMUqONnog/bbOOGFPMYVV9taJvjSb7Ma
f5mw19EnEf9cOrXA/kPGjxZB6Pj8aYxZYePBuizSEGFRG99V3bI4x8jmeseu4H4f
mSVMV5Ko4GvTi6VLFKyHGPEeZXOto23yuLmozoVH4LUTMlVhr3HXZKY+6AoyaZt5
5fbhzIEyzJ9mSOxZ469/RFlwlH9DHNkVHiESc4yPN7bob/N9hzkN4ogja8UM//06
HFz8D9H4wmaSQz3Ad4/RB/nxBCf7cUdi+WUyJHGw2GeyG0J3AcXhHNLZMVgi4SEn
ufZR2D1FlBP3WZ0vnc9mQWNvfRepQH4eK+Wj4YJdiNAPN/ywMX3msaabETdnALJn
t0ZGWB/prrFyLcmnl50N7VKzeLTgGQx9r69w6HFu/laOYHKGw29kIIyabryuDvCq
b0PXQdqYZoKd/qDlcE17h+kns9rNJL7MdBFtXy64z1o0zMFbMGrL2pnF6yHIPtfS
TdPiy9cwEpSMGiY1JL2y5CKBzGoxQDWE9yVWqtQCQW09ePMijNjZVCxBQt2Yr3Kt
9K/2Da90USBsUUFpz/oSR+n2/+mwbADSRS7xowvY/Df0zhuwHzuSMltD+HD9KaFW
LRJBVo73ESybUSFvN2K0KrRYFRgkzCsbNrUI/OljavjSCcBA9kebjC2G4seTifXJ
JAKhDxrUX5leve2eHBBOGeUy3/QmaaokFJsvbiDNnsO7Ci7wOKM41lSP+6Jmkvw2
IPCqoiOGJ6FfCQyzSrTbZtyzMEta4jLU60hBBRfOrBBzZrxCV+qCI/PQ4BseWcEh
dt7IiJhcD88nt6vXrdar6LULvMDIlBdrIojx/M7C0IilWgJt/HRMs1qUOm9eyMWp
6QqOI5gVWpM3O55KzmAW8K41+XpgMwiXhQg+8Dp5KpbnRCu0ZrUHuzl0F6zwijzT
fkkUOcvmcLlBjpKhxVsJfVEdurl3F9y2WQ34jcvn6dT24ZWZyqrmT5h/TOLv8ri3
fWLJ9CtXx9hSExK2U9Hoe5lkhpW/4dy2SQrf4sfO5ukwPs+KH6rcKn8P/TaegtS2
RwTp2ihkuT5uGIYy4BKMyc3nVena/+MYbsMs8gSQV2mpb6Lev+qAlfdq60YPwpTw
DonSW33vpXPYC4gzWbWzLhPWDHTnllj1kRrCnKIfg9yc9VeABL13pOf/11PPe4aU
XgtW3TrtcBZyDTb4lD0gKIM6as2fUZu64DmcG3O/M+0b97qazrtClm9gyi4WN12B
DFgmkSzL9V6TEVfPOLMVdEVQ5Pn1hV/o92SwaliRFvJmeqRcBG+84fxnJGwzrBbe
KOQBsdl6toyIFNUVj4+vpmP7XeVs7WWJRPoCgs+EjgnKZAP3NyUyzKDxJvsKn+J8
ejF1ALhRD3POHmB4SzfALDUhhVSa60fK9kWXMU5tYnQyU38U3lYxsh9B/2580+G0
JOQpCrnxAy2ZLCDdSk8F3+a+7whfIR7qIruor/mRqxGaNc7YltkXPXKS+IKsr/KT
+4fEcE+so9tSpzzE+UAJmPbEhAgGMkaVD2VnovNNfzP1sSBVo6kA6IVPfKQPoQv4
mQwogUOLE3BTbtfCtujHBC01JEm415GCOykzEU8YkNAvc7KTPe4RpcXxW0XYzPXz
+lRuQ7uOvTmkY+hmz0xGLVupn/99b/VpYB8YZxm475ht2rjqPm8d8K35LW7lqurT
NrDDbjLnB5wJutjWFBLAR8n52NA10L7HzjzPNEf/BWelpLaWzMmh7BzDxJVqBIhO
ZETv04mngfvqqSIOuPfilXHIxvw7yCTgve6hTN6ZIo6e/difQsa1kIMlRvk8GouK
FlLPjNLSknJLgf25bmHrx6hX50aju2fzbfZUoNIiPE6WUpQDCBRZQAMSDe3vlyq/
Xt/ltMTbMxb21JPJON5gCMI9fN4LoIVomjl/tduSyHTaqUoTxbHM0jho08hOAGfR
BGHXG1PqB07s3YviWly7NqaqWuiigw3h+FXZJ7fjWDJ3epVopvCf+VSBf6itkVH3
fyqz11H89D3NizRn8TLauLAfs85ImIM19nUGuFeKOn+zsOjCeG8cyofI14N0yyGb
KaS01UJhJB8cEha+jy4Ky3vz2EEIYSWrP2C8JTlLWiDiVDQn9Tc9mRoqaP4qZxeV
giw58yToIuErju/wetwD8F3LDf9pkh22vXYBgM+ltm9zxegmLO8JUqjbUhNwwKBD
fETnIyK7Eexo9YjBe8jL1lyJwZWhXdgFrDL6MFoxTPpC0UZo8Qd575kTbdp6NSBj
UtjIcG9d/75OlbREDclV61Asm4giZOSD5y5Gaztn+Pa4w2KZxa7RFiLUAdKSzHAI
zn2qMoS1AMne6jZj0ockRKDBbKDypZKUc2fkBw5zQV/lxOLb58aC1cuHSFaVrFQ3
bsoSDm5n9nJ8VXkI81Ht420S3Vy2fYVjyjqF9DawuwYHBnQ6L5IDc/bhkl2XODgS
+2qGXsiBzNUb9Iaj749czSknYUukFU1u4jhj+aeFyjW3vWYEi4pzlhThm14QBfxg
9r+K3qiaklYM2DdOB80WXCN2iC1TET5HbCs0sCO3x2Zrr8rYR6nG6t7lwDOOjFaz
orxb1HotqAtYqDiA8vE/QtCPPQSduloSUvVwAozhoT4fTaFjskzQHD6OtElCmlXs
EfYc+3xj5TKFw+Sed6ubbpJLelZNRdS5W0MFl6MMGodO+a3IXypr5TUmyMVgYFoV
oLvEzsJP4z8bSPeFmQcOej7SIT8NYkYtUZ23+MtyAa0oib43S/eFxXsefTh7Lieg
pIiVLJ3BiwuTInG/nOGi7HrKH0AXzxarug52eG4J40yiCbHnqn/nMp40UkEU9RqQ
Vw9QcngJX0zFp0156uPXmPo4mDDYrjZlW3R1BzsyyPqNcaz+0PmZdxWUqRs7dnoV
39HCIj4iBrmAhvf8XPDpN9L4jJ6SSWSQH43mGkO8wVkdG5qtotSz/j2w4+xWgcCz
xMApJUXn31ZJE6ctCoelH4MkkhwV2aaSpLHjDU6JhCdmAvtgBRDYXxPlcKdQGg0O
DAnss7Bp+zHH+Q7Q/i1mAAdvYKuXoL6+NU3F/E/jKw9/dIBFFuqec3zv4O5HMtaX
Wh3Z+yYP/VQSk3XgJiVGoyl8f2LDsd5nS8oek6VTjVnFSiVi3E7uhaJatbLLGc7R
iH/gI+RyXMYZG9GbXSz4jwGx6tFDrZ2dRem67NLfftH1ZwWUb8JSVjp9BDxUFAUe
33b5wVCM4zncizLsgZrstUyAv917j9TgFLWNO593ajTcTWM5Zji3hPakG8hCer32
rvL0SALqq21UO73GYR/Ioy9nd9rhisjNTVKR5Ia7coZdPnVmftNc7c6ymVsb7GS3
t9okidsWHHEzvJvKIwwP+YB0n9owBEMmS9kbvR2BcAUxRKiqGXHItdLxzOKmMdA0
Mrkc7E6NXCMsQguJXZUb2IMitAEOUATTywCaJ/L9sF79cA35lL0E644d3Ok8UD9x
yeZ6GwVfn5l/a1ok1hZLQ9J+CZRLmMcjC76eQ50dAoHYcnxIbUGtU1IJyjIoVP3S
/5+hpLQ0JUY06uzeIuxeYyC/kuc6VE9cakvbX4K6YvX6HzD+brEdU1TIQKYq9R9n
TDaW9ZXLc7Gj3NvQGH4d08AcrFh8W8cSjCK9RBHNa2X9IdkulAj0IRdJf6nXQlHb
2kibwPawUJMs+75iYN1w8e06rZJbagDkRk5se/7OovmZYMQahc1JyzntanGBdBOl
csPqxb3avJZxlH7/Ths5lBNUkh9cXqnlbUs9frObLK2m3XUNpq6gpxdMZiuFWNWO
VAPXyXkJMus/WHUcRs10EzJ5ciodKOiEIffJIfxSq6uza1+zcurjYcXatrfXuYtI
VDGvFy35N1ApN0e0Fkj+kxXZrcGxz8n1cWLjtxj00Zzb/KE63lwgHLeMzV92dYg/
cW0QPHn/SGlN192hGENsHE7qQIkTCVn1wzE1R3ru0okTWKADLmW5QVeo4ymR+kaR
F8SNWBKTjxc0P1eXW/5dyjSgbwd2VeMiAOV57MPvqZuhpcNoKRjQgyshizLBgboJ
FbM6qN+T0FnMD0tpd5Vvpk/5VNsGTysN63UTY1ViQL0eB1Y6/45n5gpooX2nFzCA
ISwURpRnCT/eNeLP6/JCNrUTno0Klye2+IV0p4b4WQQyvRMbSweBNjt3CJnCfgNo
05P1dvmVHeX0vnMXzu/15aJ+u+bNrpEtr7kQEXF0+0o8WPOauYeHFluQSL3JttMm
kOTFkFdFbYJxZqYTk9wSOchwCsPW2LTcIhoXnExZgXewXmd2YCh9BhY/trXCaxId
uNIBY/DKM34d/0PN/3uvRqvJY0sYJG3V4KuQBjRK7F+qS1ZIc8GdTp94EjH2OioN
ohMMYwjRXWUwY0e1zoEoWR3fxDUMW0WYlsViJCQBOaPKeKgh9F/jldaRQ9zIF1JA
IwgZ+CUnOok6iApLnbEwzs+LcuvUB0nZRnEC0dtFEf5v6a1IVUryybzWqhtnN7iF
TZdaxBhf7cAURYK7KzcH2a/UXg5DIXsYcamdtjgEqskuT2l8iYcDwSFiR9HCWX/C
pWTm50QY0NV0yD0uaSoOeSWqwJ9OxuU8KohNdnPJxUbmYMwhgYOxhzo/BaXibc9d
bag8a20l03EApIrbTSKV7SfujW6ycolzrncCWNBppa72AcCwnXTRs3JXBVzMKK2P
EKD4fpl5985KiNX3koChO9nt4ghPkfzsto29jsUOrK05lcEDikq3ecQ7EsVLUd0d
I2p1plETSIe9VvPdSPpVjdmNRV5W7Fnhf0V9ihwIkJ++yyjhWx2xAd9+J3BOT3Rq
8chpvadph++BV0hKQhwm49LfKo5uxMZJVDQz02vj1mEAXEzyjG1e4E0NW+GPjeZ1
RIpw63D0zcULDvWguOugrY7YyeCeynszm521w5EkUk7ayhtntFdhCPrB5zR7uIHb
iLH1FNL8PFEcJTI+p40vMqoUtcOP9/5ymtDAaYYfd6SbAtiyYCaT89K6opjklyxG
MXJzaXXi6JjZnzDPHAi9iHKjt+ZjniLY03KifXG96balGGRXbtQ2xeuk1AhdGLjS
wWAxwU9dwTBFvFc7g2q5ginkXJkeKKMPciajN763B6uylL68yaKo15ZudjYUEVjL
kauojQz9TKDHdSh6cadkcYMXBI5owd4ldZdjqyx6TjC5EWlYxbAnWiPy7RoCNvK9
joy370lr0hd1Yk7H4kiJBZIr5j+4si74fYARlU5k9fzz20X4Kw12bbsX6MnmyKx2
RoJYHjzZoMbSxKsr4OgPLqRhuwAU7vU/WDlC3HG9B25gwKs+XPSfR8LUczwfstxv
D1uEJom/YveU0NopwxNhhoB/HiZxSbogoVes8iYWwDK91BfYTGXpG65k8QEGt7ps
KkzX9bRt5aL6mpGpWgE9pVndKnSP/NsbsEem5V9R+DErP/R7tvufm8gOO9fYO3eU
osBYeul60m3l141DYx6Ixu5dkTcClQOHEpDrRMzUhRYjyDVQcfoaC2oEi+lfDOfj
x02jD1/AgV3TVcf9XQDVFmsVLqceMZm6JcyUkMmnWAFNvKuSzJmxg0U/wJ5FcAox
W5qP/bkH/fV81ZVzWTTiTd0EaNAmWDcbTw4Cma9SRAwsxlUzK/LEq1sfQdYvYfos
Ik0H1hbS3qxx95DeIJw1CQbG8Sus9GlQ/7AgFq2yf5UB85BHLYuWk6TUtrDAp9Gm
IWqj6jr2hommrLY8aOrHeBi7+L2plsv5LAyQYpr5mJhGOsPiplKiKmsMznh1A7vf
2ZOqeZcebu4Qa21MTGqtgH3HqtXJptKjgr6wFn1pn0TtHoZyTdPRW7LhhGUuzsa5
ck6CSdRVqhQRlsjSWvp7YFd+8g3KUVzdvoTSlTclwnaOUZRhBrhafhiVv5md4ZyG
d3jQurc6T904JygXfJERO/O2XWfQFC6JaZZMI6AY/M/zxJVe2TQHTdoCFvLnzec3
JvnwFRjYoY2BWfqn/E90Ma4LZdjK2rUgc1xUKhKPhsYsi4iJV/xJX0XmxY5MatzZ
h/dhVe9F3YeAMXhv8YcEDhI4rshDMHxQ4sPL2G0imbWElVgpvkhrBjurwVajlR4g
DQ0EFgADeMwxMpHmG3ZSVUei/Iy8guI0Zw/VMu4BF+a4Xd59s5uMgzOKuEgmv29t
znSJcWTjTL9h7t5o+Q1+53aBcX2ozyAalN2+Ham3LJRy096Q24SwlNcXpnPYA3nN
si6NihNi48/iGolPqY4KVrGDs/pENzq9nyKgAt4hLcPAjANIswyYaSha8jmLNsXX
9SoK7YIpwu6mGT9EeZH1j1serA8SI8Bj54yRkGwZmSPbkHf6QOnSFcBgObvqhWji
odYsvbZyxvHlZmq3s1c+iVI25+jYZqmWFqIEPi7E4TOuXfylGrYaNZSaCxLtFhEa
wNnzEkGeqjx7d1YxEpLM4DN68yIrGWYGKu5nDSMo4BsvpkWDQKWONkR/C62gwZGd
EEIGqLM9gdHmWtUIfinIDskdAZuwQ2zjiksfGs/6ImSvhD/3uoAZ38AEkPykJOCf
8vaXsDgu81iMhkNyTGKkvDZ3SNcyh6SLY7UQdKvC3kPAacg5RPtZGNjUfDVDNMdz
G1D4C7pDZtvX2frJmuibGTIlXqI9w247C9f5lZVHGDbHpujlkyLY7zHVfLuxBXzk
Bg4tQOAVJfFLMexTQpwd6O2/h+wGGvrx1woUNO5BYUptffBR694OI4RITfPYSy9M
4K9+YOgjJe0MMTQWbg7/zDqesIScMIY+CVsH5u7WrjnMMpyYqUd3uwK6dPcNs/zO
QoZyjbs+FKEIJHkXgGluqS+v+uLGFwO9/BrLxeRpFFyzoEoJTkQNhUaKb2ptCFY/
QWa18/pB05CkLpBmLJalH06ZtCjf9RIz1vRnxcHFnHp7HlJK1wm7b2aChqH0gS+p
mP+4Sxhta+Y0/o7gPxuSGAM3q3eR0A5NlZofu8/AwDxFDFAo+YiRpGbMTDY4OCHe
TZyHvhxq+yyLARQ6aao9sbg9nYKwBkcbUBXQ3OJNi0JmZCcQxC0uYXTiB1jXi1Ip
eKK73kpqqRp1hxGz0bqeHAaXwvJFoadeSUFoDFNzgh2qzl2nYiviGggrAnzExids
AxWRrwqT0qdLRWMXJZSeUbtRaeDw72iNoTbIjbnpngsIuq8JmpqecoH8vFWcy3j2
p/lTvkQ+psUl1vx+qLu/Rfbovnt1i/kiRyFj2CnlqJNFySwGnkf7iEJneM26t73I
G/mtOg5py5uKMIKGN3tiovJjJ8x4PqfAVIB7l7Cq6+FuE9eZiz4m9P1CPYsKicjb
q1mqkQ5OHxQDVrekPid3RnTMkbVlX2Vwfmd/zvwojbvdqo5IvOboM++9HbougNv6
4rwXPUe1bRs1BfkelT0WN8/1pStX8mcoQWipA281mqaIcUgODbGlx7NzPFNrKf7V
9leBzXAtd4zvdTpUTsKUQfThxM6RGtJkycQANazgVi/L0a6GEj38QIGiQJvg06fC
rFmneqxycn5YQaslUK8y69y7VOYaVnHyHUA6dsSlcWDTGvgsdPp1wUmja5D9LPt3
ThcchDeIGD59dmmWevrgX/L0s/vNI6sB2vOjr8xjl53DIWxcCO7FPaxGCXYr5608
Yt5oEpoKxmBdZJJIeltcdnYKqnBYEG0eSjCWTQzeCP3fqJTAf1ZEOjXTCqD2db0y
fSk0d8/IJT0lBls2GSd1J1MEcc894d5yp85gwUEHjmk+OMmI8TwvZRrbzeaImsc7
CzFyLdJGrYCse4nnhiuDJz0ruuC0e7Wl5HZ25Q30Pux38grg6LVwX8VwbVSgVn7i
B9GZ11Fjo1jqGFC6GBRBf/gNGg8UbU7eRIODrvjGq+oDN2zDO7tcno4f8jSz+gQC
vnmcANDsfmLFmzvkdy+IXgtBt88OObM6CMzeLY1OnR5d64o0WTsKocH18O3etKu2
zhs2d7KpZXl3ZRqf+WCya39eM5O4aaZPJ3Hpp54EYq7f1S/5DS7Gr3ITxL1FI7Ua
Gsg/JjmagSofiYzbAtMe7AXDdxW6inOW7Dn+hILA5nOtEVcBBIcA02FWHGjKGgG/
bA0EAEpi6A+5Tq4cLKaeQPm6u7VkYRWwacnMLQHV3s9osCByv8V5NaGxAb4lrU2P
pwcS5hFRIbj20DYfXyU4kgl5QclcOtt0D0Ziw73aUpWWLxAkzd4kYnwr/LDr8axa
9lsDdE+H22sI6oOaKI2XrTF9Qfqu5FvP9EDlliib4yxE5LAUbPRWmvTJWeBFEdf1
OTmF5QYjxkpMfIwKDl+s8o3Dy5VitXcyp5gkwWIdR5mfSbiisuGkHVrFCb51bkBs
DLq4uucE4MlhnUjYns96ejoeWndU823Eibs0kbKROUGWgez0iP9YcEncKdnpAnWj
zMi5uZ6lShvAzLFaS0Xwx+qNoYfN5bcsnyzuXcdndrmo48OJv1oRDPPxB/nVGEWo
cdx6l3tgQmEhERUkmMmcEF3ORdffh08W5JmuIrDwSSoJPCAtoPt79XERSTnoUKXj
7cauhYO+INtd/b8uoArYKMYQL6WUCFXEcIdTGD95nyzjxVRRygqOgcpS74bI1zQR
tT5rBic43yejHlMNsHTUU2xcrWt0tjpuTRAGuvPfCbTZhISePqJhXmMzkWrlIPQD
QUMJ0rOPl4WnXolq5xjgWuq/hY9FuGJspPCnCfz1k5Qm+8bIsW74TnGMM5Yx4BJE
b9M1ssBtcz0w8YJShjZ5FenV6YborCpOBLdiiiX3DU4WjXWF4BuUnHRaOkhpzpX/
t9nbdmOhbO2NTCt4nOGeVF4mqEBOFUxAD+982fPIEhT3haO2wK5KmSHEGcq1LenA
r15KHoUrgeI/dtUljjbXGdGxgXVtaxuQ/ApEF03L2+1fS3mp+1SNd+Syn8WwpNdg
OikjrltgCqRLs7Ryv3+Ig3QnlP6V81iDX+rNecsAX3Ap8ziJdfsi8BNEv+OMCIRP
xqlswKp+uNVOoByGHvhrFo2R4AHFE1rcuGJJwMLCD8C1bH6NNpgrLL4rmQ/UvlRb
lyk7q4nSDqu0A9rzK4KYNhMDh7sGMb+CQl8YlgYdnIQ8RGLMRIaDgRbzt3mNCNE4
5OXG7SZsai6Lt6OvP+SVXIrowaWHH9IAixgJUbuweBMju6Drs5tjhjMoJoc0/hpN
OttkS4uSpkU6Rcxu/J5ohpf8gVtdABw1X9DOD2dr/5rFEKrQcPuVu8vInM5czwLo
pIfMzcUUOO8VcmiVHspQBhgz+1VURrehijj6FhN2+FyxxAT0ULw6sXbIyg+rls/Y
BFgv8hIZay2TxrAFONU4jG7UPpG+Ozc6YsMY/9BDGLYXZnul76DasgiMb3C6j072
wPjto0ZJ4nIuWoqEwM3iRxSatcIlaS64LQgIeioZdbN7VUNUm77zKlq8GB7IRZDX
PrhpnzqTWf+P5paWhQaWVAhmZsII0A/1//JjUFpFZZy9yhm+dtKIDGkbL1C53eYK
kiIJ/aDoJF0c61OHsWz55YsjMwbcO1EVs8LTftbYtbbrT7q3A3XwOMb1V5YmpZcx
ThbxAdbMOjO4KR+YMWrOOsCkrAVq7ZTI7NgQJG2EACFolXytRFUNrdC07bPcOImc
G7VeGRrwT7pfcava8PhJQKDAtzMWzbbL4V0jF6mARB+Nt6WifQJX8g6FcLQJGzfp
TvbQVW+YNOm1i7BnsdwMCHJnrzQfM1Z5kLxb5wsMsCq5ESj5S2fJMMAXu0VzfMz1
1w0+3AL09b8dwGoB6tLmc7qFzlN2/Oxuv0wI8wB2rUVn8aOxuB/dWjMEOXK5LJm/
LpuSrCagyXij8QjkY3KUDDGB+k33P5BKLoXrn4r1q/YT0BEOtwpkVAFh3alR0dru
5AigOXVnYfnyrdG8FYlS/1cNjI5Flttay/bNf53OuJ5ClQE68zOc3geAfB2klb7b
YclnZYaw+xTsZeJagpNJwuXfxB9Q8VSNP8jTVLpNf70pBfaVcTiDWQ6JGUetyLTM
/m8HE1+XM1jwDzqSj+TSJsCzCMeC9U1lEQOLZa1iqeVBdfM/4j1VKzX4wZD3tMiQ
ty/yZIAu03yj/pMu6N0TOxblNGDWb0xU7OZuGLGZ0IVBYbr7Pr7OO2g3LjWpzGLw
+g348csukAKu/9Jh4YQoH+N1UtIQs4F1k+RvCb0dvVKfbtZ7k7oxoCfMqI7Q2nKr
ZGDIBgJJH/UI8XQJdA+1eVdiP9gCIUw6G2x54YzWxR4hH1XH0AqTSVZiNcV8E5Jy
6NRm9SDMkhkud+EuHdCDxE92Or/V6oc+IlPttv7THa78OVNJo4mK9+K6p8VCnTU2
Vd96CYSPioedV2eI4O4W43417MnQ+p2cc5HlgvQb2Ya43byJWne2l90XY+RwMBR0
lqyyMeL6xBl0AvcnSnE1WKW7Gx7iliUWpmJUkdtnYQDIBQtauubkiQHcIRb2vhoY
VuD4ZSRVuk089nATt/IoPRahiTNiy/1+HTpIYz8SONI9Rv5v7PUqStzT0o9V4jMm
7f2dEyHSU+D3WC/41ZR7ayxl8jgRUmwbjci5gGRbo2r1csnWDmp8JeoyCRQcQkm7
6OA8t5qsvfPgCdocHzPNjn6seUGBWr51wAo1X9n1synID6I2ZPEB33fsaOsDSOow
6d4sFfbYYmgVL8qSLHg/WyciljZIX+deX1T0pgK09u89JH8S6IPeSgSKmj9gAdYA
oxYcm8ZGycLPBaERovzijj9DIyl/GwJ9yMu75YUHt6o2ihkonTHy6lpjPrnk3ma6
51PBZxgKBHTlnPpS6zPkhhBGtVfuJrUR6BpoGaBR7YjJmbnmyBxJoLT4VNO7SkQH
izbE/QI9BDI4unb3/6dlNaCEESmOio7jylP9wyRDl6C8S/BEIAzAM4QaWzQPS3yG
bDVvWwOEC5t+3xmjP4D2jAIkHNMpFqRzEvJrQV0w507qklhX9rN1AwS4+wBHv+V8
u6ibcI9Oh9FSKR/7UB0PxNHhxtZbdxOxxA8z6ScNvz3ck5nhCEp2ARXJ1/FHv7YO
eO+IwZU5aWDbDvmSdOxaxCI4fNVgkO4LtYuq8N3V6mugCEQhDDtZzw0I0oEhJz5o
v490/n6UZKyleFwzNsrglLOZ4jp3qaOVLhA6tvaF/n3go2c6KvVEaCsn0gLexgcB
wrOFmNyRFpL7ohkaR8th1jDvmCepQrjeAzRnL3Lw/x/PQZNWv1CwGdAbsNPixiuE
RqldFA+tt3CusFjOIMCDROxYBjnV2tjx8sBDmdjBpstr3liDP1wYNGYy1JwnO3/g
6Rx6XexSzCnaPyo4ZHCD6GGaKO58ohGgdP/OHEfOIYxdhGNt1DfnJ8P9DMoM8NDI
9cfUS7G/pD96Cw/mIdv5iwLqCcf6+UVM/ABGfihyLTkClLyx2DrIe5Jfn0z2BfpD
gzlpOEGtoSEq4AhpuZ1p9NdkbtU+TQ780cJhvAp5s4zSwKlO9kMJJabAyiP+WPRa
rTo3e8v51KGOfF1DYmzl5Q1QvHz7XUOv9hR5NcV5KYF+9V0A8PngTPgSJrxq1fOc
gIhrS2b/mmvPvTqSbjJOMXyOAp7086WujiFyGjJWQH16eHLYmfSyU7Vq9nn+9z+B
qCrDjvbGZtvlfxZojIcCezfulX+ocwc6wooS/y/KmJkcpzbQa9T957t4oExdSu2w
BZ1rqYZ2I27uViH6grW/Q4YQOOFQo2LM38FNkUVswly9UBxnDc34CBZbzZ2sIO9D
AlIfxMx7BQ3x1RfhTnPh/mJTYeRIOpkK7U93xpGinL0ZrolrttjPEAKm9kPDPeTt
WxYMlKPMibap573bK5xYLFqOvnHXzYflphU6WOZMbK0WlDbF6w9cFL25prguH+Ul
kIItO9uJ0Ly1fyF64vLzyGz1K859dshskci3CogXipd/Yf+CRmeFF1hom3rKk3Pd
1LS0/zSwzfgej4QJ51DplwYnPDGI9Pf94GPUbJJ+b0lGid0gawF3i897IRE3L5IX
93L/xwcV3vI3pkDqMuxGV2y0d5NV6f4g4qktWDLPO/PDHJmTIgB533dHyme2/1jo
uQtF91hMKSuwq+ec/uJQaRHgN9bbRpZkXZARbhvDCulK2HUcAjrNUvCS8LVH9x0p
8xNt1lMAErwtdfgk1geSkKGr0scFbPRfOEJs2Fg2oAz3BO8KM+olycT1nDmMWHNE
14lZD9enP0nxIlX3BuL/xp4RzkYxhMhc1g10uMtk0CimUU1fkyTUJQQnQPZT1AII
iV3ebBwCbaEVFtZJSlph5kgzZOhcdrq/4S1KggTCuCC3REqlYYQag4FCd7GrlG00
l5PbRwKTCtmeLcMClHyHXUXamwKAan7UbZZKDU61YiKL0SPhRKjHGRcj7XQ0YYUx
sLp5HOmv6aVw900TQ/EewEy2K+YMARHgAx6iSkc1A3O+RNQ0g/A0nK9vanuu6Fjl
YiXn1mgfE49i3YlY4kSUu+WabeKC1E7nk5/Fh6lCvlzJHEBDyKFoF0gA3PHRN0qd
7amDjTn8CfJkwxFxNHNhRkKrG7ocMs/pfAwz8QytZdxZwAEbX/nI/Dv4T4moy1JP
gPYPsGiMGK+I9/kpaE33pQMRz0MDf4xOMHtd/u/e4tkeNn3rS0enJrUkyS7zz+YA
E1jlYWtC+8bW3D0ZBH+514mDEFjEAC9SHtVL1hrAEmkjzK5eTIoEqqpt87jA2Cl0
e8ttIM1pLn7457CfAxFOS0yYlajPdKeAeoXdmWa1DBqqkmkALHDJlQ6bAFNJ99rH
y7jr/MR5mEpfA7TO/7gfsEjluN8kJ/GbFVP3gtXKWf7c64XJz+3nalvb961PRu7x
xe/cEYuouL+Zl7WXZX4Pg3i1S0j7v8xzw2sAIetKgZFBy/iU2AlICHsxDQYJetZz
1yG+v48uIfYlWlxOvoJNIoG75Xpr8bz8G5eJb1gVLHeQcqrq8ke8EcZy1+y+l1Pc
6ZoANoJZqp5Vue2uyR1K5kw37ribJExM/A4A7zt3qVI+iKnWAYDgHCyV/RDDd9Rl
7ZqgnDBY5b8qfoVJA1fx6PGqnBpx1Vif4Q/wACfsxcm6ElMHS7W4+upwQlI9r+Ap
9sp52PQvi2+o/2y5jVUHfqkyptK7pxjqv8wbhLERJ9a7MsysNm2K3iiPla0wYFvF
PUroAVlUrkDyeLiuEZ1cEctWQIgApvurpT/6/cbsYGD6Cp7j6bX7kDMtC4y7UqpP
ooRzd9OjwsiRk//P1O47Ef8uZLapXebk2gRptAqxzBpyuPGYkanqIy9nGUCBqLZr
RCvzxjkEtGLpfiZcWaTE//Nvtdjlxdzl5C/kXNNRGAC4lXmL3PdEFTAgSHAdJY0c
kGVAAUzQQfdzYXzNSf53NZKHPcQ1QQBLgUVE7dsRohK3hqJEa3Wn5pkv8PYZPxXS
i+0VZ+orzwjKh0ZuoQaGtmxxzt858F+2KO802YJ/gs5PIW9BCZtkPV+i5tKGQDiM
17VTpj8llz6OAK65bnZ7hd6tsUl8Vfht06jW4j7Di/UzDgUaVI+fpc1SpqPzEcGS
t67XUqZn8uCY3gGcKVlVBMK5pxHSAj3p6ND99F/jHATzQ9Ez3ffG5s7aSneabOfx
weyZ0nncEJhLP01rpDXgB4wfS+yMu/vU1td+hmJC/SPuKIk8TnNiv/9lmrH6ewNw
dU5I8710YKU8SwCIq1MTVyulEKD4wO8wnm3hy3cWjnKzHlLUek0KzdY4WA/LvN2g
ESfjjystFW4aOxx1Bw9xvTK387f3JyVEU8r163knMOaCjXioHSW/if4VCwI8YNq1
CIH6A+O7twm2cfy2NTsnLfWdulGaboY5qZrbq1meHQFHiy0GCpLai0yJHBfhmLoA
62TqoivoFMEl7okF+0uCEHk08fpZKISrgdx/DPaPOZuHEQtAMcPWQM7F/jH6eLi8
SyL287Rmazyu/hKVN2UmbYnHOtOHM3ah4Oha0brRljeG1UV5VAt0XZja9N164lZx
p0aCswBz2O0JgOgZjBXVyk5i12a70kXBMSHnNMmrZ2pnftErEhhGV9hWTLI7U/wG
WQRek/KJmlJhBSQek6ZHm33EuyZN+2gua7DdYEvhzIH5BH/HGcXFJKowz4ahgXya
4S7sMAj+KVlCbxWJkMI3d7yEr5Q3Ao5C2g11CzjGV5wM/3amARqLRw5Pe5Utf95e
91FwW7xcKeG1ieybiIsqF3i/3YJjDsVyR/W6MgF/fz3KOnb2x+t29MVCeg9PdXxR
6BPjWTxN3zKh/K05Ey5ygTmvmW3djx2z7Jlw+713DmlwiSmtykZZQY+h8HVknDib
VOxy6xCmjCbaCEXuTjQPgGpCRmApBUpWdV85BBnqaJx7wzUjlYNdP0z9KmGZ6b4O
BfXo4A4xB6ydN/CKkV/wU/xcn8GPrJZ7jTvk7y9SqkWdgtEgqfj8VV8BsUoTNsLa
dPiYvP+jRmHYTauS+4DmWpGE0UimLTMFtOOkwpR93CadIGIV02bnYuMb5YKE5YmI
fIVpjUXg79MIpla4NgK1gU6UlIqEHCZCfn/P1HOXKjyFYuWuhKJJwAzIp0QJoDpF
gISw8iobwZd7tZ8mD5UAyxNrkK51m6AD7cftVKu/jcVxg6A0S8DvvXwRaVxAGlD0
clRCONpj2hHBRX4p7vhQsPLiV5kLI1+ej7TBRAPvzKS/fkUYMzo9+zLOcIHcxmBV
l14t4TI5JLieneKXuj6JYsJyICvDXPI/Xev9FO3cgUWKxH7ptuFel7TLjR3DDK3Y
dCOuhOJqzJN01cT19QkVvmiPAiZJEc/n79QV7KpJZVDAOm/EwsSpFlOCbJfpbGyB
Er0754eV1UTzy2SsGCPxyZz4TaxtHBul4SWZDksaAIu+y0ENVsKOKiyZjqVDNulU
Qn0JJV4FVo1PzFN/tF4BXtPvVgVfAlpySMIBqO0HiDOk+oiiXYqIrBem+BeQNMel
jKDptxhmBrWFERMjgKzZ0Z687C246PwXxRhqnh9t3yeaQ7BXu1ALGY/anBONatUc
MdWK06Ydjjvmqkdeb5UBFpHlScIoIzu4VlnhFhOY8Cy4VvBe6A4xmYQ1W9gIfEmJ
FysHWh34LIFHPvwrxVRZNsdPSjB97bzJYuzf8eU5uQuNDPAuKaOxbb9KEczEIPgf
F4U1KYHqnMLlYJqQ+uYm1tWg7oLmdZyPU+aK8bnhFLlM2+cKMz+ETENzO9R4WYpi
hIKQwkkWBwqn9LOw3kXx04I7YgaO8ZX6PmaX5FQWXGdFnXgJSFeWbdZbJrtSXhZH
Q2QMp1oc26+oHpMP/fPPgb9M0mOuhEGqhHj9axVhKYHOcsMogpVlKgiee+AIuUwk
hTBTzJRQYiEpe1oFazdmqA1zRvR1ocYQ+1gxcF6rm+JyRtJTMxcOObD7sMdka61y
oHgaufDaCifDLlVQPopn00Mmz3IplbbYLLsur+HA9JrEevOmpu/WfdHDFyKk7cSe
rUdke+936LaPy1MLBIQV5w4gHwWM9yRcpqQG1SyIb/G7jhVTQI4RvkmxnVDNIE1n
84Fk4Hv4dfCgtOyTfPSxFmZys+53HC/TZRGzAdZqzyT4zOlPuzyVAkn0qmByXKGg
78XzlHY1e7UmOgYnqmnDu1vBbKL9FpORDtjLoXC35CjsmvngkKNv5Kbrum64L/qR
NntCZPwUkpLTUB06sOhvKCI3Kg5naz+99KJMs2NrliHWl2kXBd5o1Vk++dffNYNR
DuvtzosR1uAH26WamNGVPlYbt71C9eSUJusmooTPvl83hB2EYbfUmPDq+yiKom/G
hsOVEq1mLS6hxEcn1jWRrnvrkRh2Nq9NERF0S2gFIrqXT4bFqwWdG5uPd3cnAGIZ
C6482Ic9rHiXzykQWt2rb3PpODpo+3g0zmuPHRVfqzZ2mdHaHZc/LfH6G5ksqZW7
1OGTtuRsxHGSl+e+1V4Yy8YVmqQhYOVMksGBoQrjSQEaBulcbKUNC7Mi0T+h1dyu
McgcZgRoBdvx5e4Kbd+qefGPLZBE5txvkAIhHnnsCpTUUZSIa1atPXhOllAdNyKS
PsNTT/bI5PKZkZd2Kehy4nDrBmMjLWTLLh4at/NBEnyQFnaUuLr5goqOU9ZiELdr
qSuBJwhSTeeUP0srFvDMZU9Jv8PzjolYR0DhsHPGsrrRqN+NTdBi0tZf9SzeUDyV
dwTQMPcdUK0OYdOcN/n02c0wS1i4i1mDVBcQCdf0mpNPBAgZBIgw8rFNXpgdFJ2j
B0BAg3p9O9nYozB8WSg7WfHLNw084zKOIV1z31O4uu/C438tmEgD7X6/EtPu4pKr
4/D76YLWcwnqQ9Jz/KAf5pJorB3z+WjKbZX048Lo873MUg6gUIFnwp9iwWETRFVr
m3IzEfhAgKJEfYpMKxoBnbLrmWGeehT45w2GFLeoWhmzuhYQ+G19UANQe9z/o6vN
PN8NU9LbdRbXmDd8R6txXcR8d9SaTIrraGUH2kNWEhPDQHQIvZj2PBWMQ25p5OYQ
Y2MUwdHJRCnkqtla/F1oUVel2Ok8GIu6BHtjqZz0upz+HWr7YdIelVuFJCXAjNkQ
9PC0Lf2L5QScMT5d8BiSnDWHqyNfIofOeisLIDBdD+a2T6Ho2S+NHCRRX4GTOr1k
aSYhUHzDvB+G1dHWht0qMyPnybog1ETg/N68b0+2QnMz16lUl1cJ68b5gqbf5KkP
O8FpGZTNO/a5p+McIlfpc96psOFuIiuhylPKTtxluxaFQ52VwZmV1a5cXU6gkXUM
2ygI8PwtxIW0bIDQo1hfcw0iBpqIwHBJXn2NuLOtVtbsSbka4CtvXIj8eQf5I3BL
SPNfcIQw6w5QOAUEghPLukRkWPoroMUSo1eFSAnX5W/drOezKQSRv87wLZGGasne
364ZUnL1OP3qnTV2OcxwM+p+iPMUKtLaz1HZmgBPZihtUcAh7Ohhe3Yku+5Dw7tA
tiKJbNHHwlYlgxdwdW7hR3sn/1Nki4p/4ppR6EL4gjYyB//JC8KOlfIVx/HrL2ee
kcaTZFc1GMtO/M63IcACG32FxoL6yGkyzRJR1+CjzKsDEYpTxm5serLIyfUnA4FV
eqcZ59zAmBgeW5nQRDCGRbHY30PidJN9uur6Gbrxc4z14rZVa3wr2H5Ploxxfrxu
gVEnPYiDLNn+FNjG69KW2dzWBrmIxI0uHI5M5PJX2puu5ye9WSMmv+LJTwo240cp
QX2pnTDzHOfw7+aMVEzAUe4v0wQzHB/3vPLFn24AarguIzmgaGTQUSm+SuFokQ1k
CRKwNlMzLpW/BFV1f3CXE0jjni1z6iLS605tCfNZg3d6uJVBrtb38C+HoZkYG+Zc
cxFQTYIJy2d3clQOtT3wvTXskkIg+iO9Keb8aDdCCH2gqfdCXNkye8oGBpIZqA7c
l6Bkcm6YB2pso2L0KwJyylmJ3XXrJNSNwwfBxDK3/oR0TzQyK+sjnlSxZCVK+2As
tNLUNB4HMZziVQ1BrSzXM5Rzq923M7jBYLNKSojLySObj0G9BuYYwsaLCYiT+Ug6
Pi9x0Kz/yNoMVPEcTiwx461NAWYMeXLdPz/gvOxf8xc6vSSLc7czyqO+Ee5CIgXu
oDWJl63SMPArFtompjSBk8rOe+L72l78xS1JjeoC7xwgxjPXpv18ss1PZwTANcO5
u6rlQMo+0w4F1+N6eWAV2EqoMDITdwib+9oimV3ztY6wBUgUNf9YnPqpUR5Ypf1T
avWrDQpVUdTIy84pmTHtxraWv4TtJEMxB1DBVGuqmYd8SukdsB64ftXSpp8oXuGU
a6mKrV9dmlZnB9THyXGSemv2/wJBM2adAWxOjCTWb+C5AQGOuF9Q2zunZS3kweqf
ueOSFVoX0MWnEy/5JVmLYkSOgc7Dxai41A0oFwmQxfTUa9u8Wtvr6dZ4q5qRnnK5
9zohAl8WHG3DxHn8Pkqy5iKb05KuHGgYIqhAtrq0uwGsyJ/ebxVpcSQ50RDeQ6yV
9B9hLH+oyKatq++H2SM9C+jSbJ6yB/k7G75f2EqhIMTI/Wip+o6dEON9IQnh+FMS
WQnlrEjASeo1qryL3xgk1zwQJn4+g5R/qzujuWeuFLpcNbSDiV6PRslQXgs9sgTf
J7jlRjXNVT73c/81mxIAQkrFdc2px0zIz7r50tplzXr4KKOGladZ93RjraktfNqK
+crn2Ot8rAbwTnCctsF3kmPy32Lu4viYtA3EqEzIkTxjz0QlYg4sXyXsoUEUBGPM
2kO6k4gR6my3CIN/oiKsORxrJePuNsNjqlIVp7AglcRSiaJhyhixwVgrALSypV2o
TS9A3b9sOP55G3+U9g3gpJUYAbFtpvvhX6eDmooqXlv8HZ2dPptu5jepfPl+y6Dm
JogYpaS8oFIY9gXUFjENHJG5IVBNqLYxVenvp5gQOCnFedEmYUeH0ICabPWmORF4
OtpQHqrqyTBsqjEE5qfCAdkngIbX9qkfcQwfl4QXRFhTa6jhFc9eqdOklAsJ7P4e
/Lnh7ulCyOJiui/x971w2pZn2Y9tKkquSLqS0NeZBxy+rPzYMiUDBveV5WiIqJy/
aMqK7Eos9JGIfVJ6sHh+c3qYWL8uHmPQbjWbI/jvNDs6eBZpo/ITsroS/m9y79J+
SQF9bU+iUxQualGlPVNwZx8eaBCkbpUq6Wch9FsmqF4d2fy4SwvLNtAZOLdb1LAh
ERYgk8x3hpZyrIZ879ZIxypOSye6q55O8osfiWA59pLN0PrVN6gXJ0yvk2iQTNTL
voC5UF3CYhU7K0EyBd3yUYDPC6BC60QQ5srlKuSGdTtyiPvBbt3ar1v4Tlo/qfZ7
MN0PIWggWvfuZvbRPSMR8GSqXxlk+2dx5v9Kif/Jl68ZefW7CCLE7+ol3ESbe06l
a9QyxNND7UQLTu9k7burBX7Wze5moqWle9oy48wC+eNj6jM9NLkNyDRbWR3UhyJI
xM6FkjEYbHceBr9Qs5zKOJO19vcAUH9cCi6V4H7AllITS5vqdSet0kvVPsMC1gEv
rrCGNnn4wP5dnioNtHQBveJdIEtYV7uYTxzFrlIMGqNJJOaFx4oyBKv3iS6yMhVf
ZxoNAiT2bs2joIDACLLcJOm+sIPqkUNgPxULsabXPP/g0r+1e3JMU35SiSsf0C5K
spQeBPWNDLoBV9atVC8nFuESZiod+Wym+WnpBGMBf/TfwUZQwPof7ZbQGKAji+5X
z/MwKeTycc9d7sf8+dJ9HV8G2ycqJQF0CQwFB/6rUz96rSCUmYIb58h75HIW8OfV
1eBYewB0NTj8yhg9e5k40WOZFhThziGV8jJz1nfFBjj0x9q7RenbWPHCK+8c6C6N
7n1ZNSIBFNULkRqXoW4xyjVlLNwOhD5EU9tx+eBnFdwjnYp5Uacf/FQlOSfdth2P
j8gSgbjnmaz2iTGHgvo/YBB0IpLF0Xhdg5skE4u3+Nz3TCpfLwUae7AytsSQ7V0t
szfTOuXMRQilVA62b2C1ad9AdWTC6uUD4KHoRl73oBgB1cC/6EvYEQWGW1HS8RRB
b1PjBHuv/oWrYm7JSOMKj2Y5RWovTVZ3+iPX9r/J+ovEfDyVXrmPFFi3/yzB3rkL
3WBbd+3qThPvCUGQHyV8Dy7LiweMQ9vJR1ArCu1L8KENspG3Epdos6LklIuxpnwE
mUTV0YMeNMcE4rL1mQociYvxhMBw3vI9BLcjpmUInhiyqJ+IHTIAehHzTjhLAMhp
Z1QUStxLl6lCdUcfJ5hUtQ0L2TpsvrgBwiC9ak2oOoYt9mzOkBVQOsBCqkGqFioJ
hkT/ZQPDnHl7OQaR5hFBo3WY3g4RyHHHuh69iRAJ20FHOtmBpHQByna/F+8XPYsr
wFWyjtodN/sC7gWqGRYB8i79SM/cdSEgvsrOKUTp9znU7qpetn5Fy8CkZkBRz6PS
03rzRcOXk4NrSwbctlR0u9MwVyGLEBrXXy2q/oLXqTj33V3tqQia5tuxCGTJyOX/
yoS2hFYb/+REf04/uwKAz95ifVlm2D9uUW3AyrFq6FqG/FdRPpk9MUQ/VwubBcMx
Epcsr4bp2ZGlxwWjBlHogOQJqEjEHgDeCXMUHcOKhaBYeMeGmKv6C2x7MWKEgv4O
JK72MNSJ5J6tiry5RrY6yPvNd0xdnSE0vcvQPQs9TOkviSmTY9+vGQ/u/jECAcUf
pR6H+5NegT2Aii6Z2SouFZFBSeA5HLxiA5EZBYNJYHU44PoEaeydv+mo0L/gTbuL
K3ezpNVglPENup0fO4zuUA1cOysEwW5DWuHQx3XUVTI/tP8n5WNxpJzt8xObSClP
hoeEcY17m71WTr5frXAgtM4Ex33MAIuRwFFtZxPnzV+ojD8ItfvQPXShy+iGYog0
OT+gBN5xP8hQF00z9rF2YhvzseMekxXpfxlGcy/czrJG7YcJfDAmPm0JPbCKtZ8M
XmtMgM5lHxxHY+O8dyQ+Ax29v7fpvLLI1YbNPf4F2ZVmVem5C7a6tx+RwAG3ysZ2
FJThRUFn+PykkhbOVL3+AtJRfwvtiYaYnNvHNfjNk6PNoZwkUOs/XsXicTMHCros
9pct+u3iYVhNbp2tg3vwfhf0qEx1FNMbFZOoilzwLh/oi3HKT5kY/OZ0oLvMNI9s
Rj603pLjQZ98evQS7Bo30ONiAQ3pJBt4XFm0YowI7t8vKdOOCG9uJAczigNzGDyw
sfLP/Hqaw43F7/MdvOFE2eXT9cX4fWzRkwJWAZdjIwGHmtKzYDflk10R3RYGhYoo
eQO6sn9UibrlFyZ8nMWEelUVeTRKvgrh9CJKoAaMVgoirO2nevL0Br+HasBUJeWp
6GkqO+CjPaF0jzFWey8ASetXgv+MvdaIkSRpIgCv5t4ojiHcYf9sdEaUDG+u7iQ1
0pxJzApLLfB7e8P/0p2Bl7dLJfIt5B6OdKGQa026UOyFMzBpuS8WQbyGdfSrDthq
LorFsGBKjOG4/m/B7mtq7G9C/uMptUpxtUG17vh8ajYoPTTLn92NlF7pSsUn+uz1
mfDFWgRYZTDKLr2oiQhdDvl24eTFzbta3ILo9sSuDeaW4OyMa3+CfLAq1visYk7f
e5Z2qoV/RXmn5Th404s9Cly4cm6zVXvc5Qwposil+WWED84qp0vFxCesgipOwk0c
VsNQePshmTkdKo/BowyNupaEL1EcnydSJtt0tb4dUhui2EGOKxLz9Zqb62pthXUs
2x8YEIQkf8InTGtkvKcZio9UfmbUfXlyZxMllRtJSYw32+0uYfeLdiVGvQgT2mkV
T3SDJWHqGBO/mA/X4QPY4Fs/6grP4MGOZfBTMnBhn4Q0UvHXWH2RyKXsTKPw4ej2
s4VJ8aMWtwIFji348jAgapewrVYMcrkOTlQ9XqQbLd2z8gABxFTP8j2ZH2xs70fy
lOBJeB1j8C5zvIKZ5oNPnGsQ6EOOSgqwwCNWDyN36pylxGY4yoYRhRi/eE4zWNE3
9ytlokYaMC2E4/i8b/HQ+CXyIdVKKau/AtJcAc5My/Ig6VEqMB/yH8pnSZIHwPhi
RSpxy+u8Kp9oIlZkFGdEI5X+3ZO7rJViHFdTK3ZDz57JLNJoA+ANU6HIyg2Smwcg
tpLedcbnHXFqh9+7iRMHn43q5xcEpHeXq5VK/CjOTCMh9O6sqdNejc9QSzITeRAO
EBORPgSWZ7GIFfJhExQ9L3mp0mkemGm05h/RCUknkA8pTIUee83OGx7tFKEoSgLF
bmWTqNS24I0UW7VAzJOigtTOLSAkewCpaKhfkb+ULSSruXxdAdle1n1U+Sz/0zNz
GdSbFwBFhqEOMfOw42qvTajditZ5tR+3e5oZVa0SImjQNH5pmkBOP44mdFpSnFjZ
ml1dsTtNdvcZ8FmlP8vfrL5VcNEIP+FjjXVJN7MZUQNOyE2CHvsaDj5zdn1lU9ZL
LKXWg389NekfqwAheOpXcX0Bdf5rgUR2JI16LvENrsiNSEAuKCU6BZLdKtDkOPMF
DDdmB2MdWHh952pX4BEfhaAk/jhrgJ13tx5HrKrIQnbpsJLjsAYbE21/k5NBUjYt
rwiJD7+J67KyECtLL3BvYhkfzf+gBklgbbKwqnjFH63t8pMQPlcsuBfdv4UO/NYX
f65P7yVuGKpufjHU1QXgiL3EIV2qClkCyjhXAu7/OSGW0nFANKFjS24NXzO7tsnK
ngLUflTN8UwtQJ3aLJKg3jGXAxFIMy5N126908nsgpulVGeF5l638aA5Ocv/le4T
T3Mix0u1rVhopRC5Xoo1g7qRCHA221mETatLs6oolpNPiEHR8mFVLF7GLARLJImX
Prsf7re9HXpyHF4l+0goiATLbE5R80dxq2ihZgyIxCDtipHNdl0PRwlEGcqf1cRY
6tf0gEoZQ0iQQF7bKKUuavwLOFYJcR+udnV/0g4p80R5WHjohFiG++DRoetvW/QC
16h0M9ucJlxSxIu3/6HwlvO3SZ6zpnvO4CD7w3wF4pekzv8+LdgM3/wlcta8uJB/
71hNKiQf8R9ozY+7EMuiQkLZXByTVr17oht/F9xTq7IzTLH03aoWTqp+KpRJd0j3
6d5kWSiSbG3Atc1IjJprEwZs8wjMaJlbJViM9j/2wq49Nl/Y/3zZFceQyYuEAB55
HBoHLOBwkhVZGwPYowqPUI3B4rRPv9XQLa12e0iLgDIPmiJ3e5NWO5Lc2+DsiEOr
74KgDF+yA5Rf15w2QXNgU+Ev78dZLyF9uH/dHjEqE7LvuNdoGeZozQiGnm/cptMi
AmbWN2j/gEvnfnY75yU2yPdh/ASdV8Ugt4fXJnOJXnvx8qXA2iX8GDjD598+6V72
laQWrAWHbsmfO8gmskxU4RY3qnxnCVFW3VL8qWMhjO/j74lGZLhQTQx6mEYtZf6o
kIYZ4LUQrMrqRU+YcdWUX30CfCsUBpKgeQH5lsodzROwWlKbcAn7DRQFP99NGh3v
8uNB4JbixAyg9f0obyystP/tEGoGRbKrfURVqW7ZGFeKgBpQtkgW6FWbyBASyMJ6
7yeNrlHv9iha+vMqIsJ8ymYSqnAJH4Kyev1KY3fG0WVBgLmNirhPtfBMexX0XULv
uwFlZTZYKjflqrgYoX3A+5biWgyc4XL5T1223lh0kzEEas6z0f7vPrqjz70afNak
lbenz5lMP6sgrEoAJe3RKwKW70R/ane2T4Z8jQCW6D53OidddS6rQ3AhC6aCwn1+
g5Pq1k2Jx7yqHB5A038RmvquQiYiQhty5sfYMFwlINj6nxU1DTvkm7GYdxO+v2FT
rxeD0boKNr5a5bcUPpUgyEJ3lgtb+OcZMkOKYUKKq55qQPho3N2rtihxdq+HzE4E
ukqTNudj0EQn6gSiRG2AH6lxKsl56ZLzQsObsjVLY2jOjKf69CV1rN244vC1Aeyz
1DRsZRCtcwe5RNP5NQnRBO3xryZOJ3fjGASkcWyTUJiUcve4LGVI5BF0qOTNqg8e
WQGadfIXJFbom28Fy4cxjr5AjHX4/qaSiNwn3JcY6bE/tH8x8fmlYd9rtRx47CQz
4mMbK3nhxGbhXlGdvxVdbGBYAAaTTC7qoMTMP5LGcIPjY7DFpENbhSdCnftuQStO
MEOAjqvvgs96aoR2YvqCfyYxEpbCEta3NyqijxR+z0UzIrnvNuXtsiAXYOp+mbnS
oDKSAEUCUcoNPSPPyywh4pEiH9yCq7kMDW8/THxEpOw6/SzMs7eEzLKnzTvSqcFQ
6YskAvJqiwsWghlJD7JSV3S6TKaXkDdTdrcOoR1hi5adrb6gmm3rr1svmvjjVdNz
xPad2uGl6HRKdKmkK/EJDOBDYnpqVkM92wA6LBRKALlq/Wo33sNhPfprhEy/ryra
MTLyMp/CTNfnQNd2owkkzEEZehi+6MsaeqN0l+xqM9kEWfuXXXfQohCGRgosrD90
SIi1XmugwYZ77uh2fXtLZHGgNBwKRaC2Y/ayB8TqPTAPIvC7mgnQjF0lkBmTQbcU
/ETV16EIkOx+5jSH8HsDKUVdUtMcPB0PJclqBhqdMIedTzxre7tRTbeSZPQ34BOR
SvYnzO08tc4lq9byEYP7LnUci14JflS49wEaq6xEB4Jexs/MK/nJ0z00zXRuxxNY
SildgIJDoOVrzKC9Yrlm1Mk1C8RZEoLzJBN+BYacxXEdR7se9X7OPF43oO6o1q20
8etbmMUr8af59vbXAt+s0mWYDMZUIw2B6OIQ042J4Pzu6fqPwbd+HA3tByzSLdJD
gj5rKCpHs2kOQQs2xwH/Dv7SJcYXWBtlx/nJOf5igb+ob9b5/q7t3zi/QfmlW3KL
5rxyIka8iLKJKJt1YPoZAmwmgkOoWmgy1yqTE7k2aNs=
`pragma protect end_protected

`endif // GUARD_SVT_AHB_MASTER_UVM_SV





`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
BFMtWVXeKmK7dmAQp3TIuFszLf29CZIEslaJRj7vky9WqrVindrVN5i9xr+mPMXc
GHr7FjDLD3zRzXQ4vMAbPYbU8qEUhKfPGZnDYHXWYITznlx+gyKZuyejYqI3BF63
PBYESKMhi6kZx3+EjykvJCeX3FwZPn8kne8Vfja0fJo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 25363     )
v54+TR8DDcuFBrJHy9499XFxIQKJCWEIa1KCU4T7qpZO8XNavD/WTXs0mDot9+x0
mMS6Vs6HQtFNTU9Sj2Le7KCmpV9AtmyZhy01AryTtOUV4H/VGaskXoYq5m40V2+I
`pragma protect end_protected
