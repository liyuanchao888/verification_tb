`ifndef GUARD_SVT_AXI_SLAVE_MONITOR_CMD_UVM_SV
`define GUARD_SVT_AXI_SLAVE_MONITOR_CMD_UVM_SV

/** @cond PRIVATE */
typedef class svt_axi_port_monitor_cmd_assistant;

`protected
GQ(R#4I,MV#@D^,RD^I4]f/4[UTD12V44TV<E8ZEf8B]2>De>L8B()ERb&;2a698
1T;d#5[])W>KaCU^:,V>MF#/[SPE#M@#ZG-Kg_Y.85Re+He;)S.Q)S#L5ePT1JE2
I0US++K8a^PS@cZKEa5M<.=(aZ\17^e(BGL)MUL0HaFa-J=[>4O2Yd0a.Mc;Q2EW
77>08#\T5K32.3B;FLLHW#,C39>faa1b?0MH[,5A.SGD18I;5PRL8+cSgH8:NeM;
1adW@L]<a3LNGO:e.8N>If6QX<0D\SMa/5W,WcBb\[bX0=@C?.]Fg;-[,dTMBOF0
2(F>>9G0BVTN_7?6N-J==>YJ@UdYB.MKGEc2@c46BOL[/#Na5@1@dc@2-,?#NG7^
8<E\1;SKA^<?RP)7[G7aN/AE7.7G.V/F]JOJ(WA#LEY#c4PdJ55dAU)PY6V2:-Qa
Z16_#]]EgCPe5f?8O_3Bc<Q?2Z:;8I-+V-SF7TZ?bP;DJ1WaI]CXH7VAEI?]:C:(
X/OPgg^)K>8&CIK1IW7J;S?@-2TO,&5#]7NbM@B2P?DJ2[S>)f?8N2+7(eRKa)b6
M-VeDI=Zc7@+KZ-gDe0_(HbOVDD1F3VR+@-L4_\\AgG#RL0:2(OQe4V3fTDfZB>-
]2?COJ5>M^6UTGBZETdaLEFXOd6(f3EdEe5[W091W[Z:&Ye:5>J=.Z6>\4\#>.g0
6[T#d#A;Jbe_fAU,1#V-)2IPgOF74:JV[JIQWOOK[NU#SLgW<X\#1+:D>P7CH01D
c-\BJZ/#0U4WH-A4\B+DN[><Y7_@S5^eMc?);\(,944^FN8&[\CfC-4,XKBX@Z^(
1Ee6ML[X_;9Y5.bf5)[S<ZPe-Z;Pe1YMO]?M15BU6_].N_PG&6+E09)>&D[WJHRT
2-]QEJYHV@&C_dd^aQ^LYY0IJ9W3YM_L#QISc6?2XY)e2#/R@XG>8Bag9>E,;U,N
=X0FT.@_L=0CK_6J>XcfRH+^<,bYC8M@ScB&)bNG=4)IPMWAFUadB#a+.f[^f[I2
?U-Me[.cIYI6dPa]+Td/QYf(;dUc=Ic8g[B[TB8GIRK;TL-K^.-N2>Qb?.OfDa25
FKd(VO3R)IfUTLb/_>Lb]2DFNX]LeeW9;JU+[c.c0L][PJ)3D:JT4=J/(@/QHYP-
>_+SX](8G\)G7/KCPb#G3[8,[M&Wg-N;_McB4F9+dg6TN5c6O5D<a#\a9_4LRMfF
=Z<50-P(IBG8M6TB@QC.P5/D@A_=WYBLf9bVDO>W5;L]-G/DR#_S]FFY&30?7[9c
=JM&MWDGV]46AE<F8@MEgafK-YQN,?4c?6K0SDZL#<0KM1LaYEU7_^O=,BQ>Z#[H
#THA3/\LP7\cCQB.H72S=\>G+,AJI2.T,#[EG,-9,=S9KU5V[&6W[_#<>6,:I<)Q
GNZ)RGd0.Z)f(/RLfMXa3B9<J4Zb._e8WPHDad5Q&Ga\:YB.eJGF+Ac0[7de0_<5
=#XBcT:;dfCY3-_F(3M7ee86F8e7a9dBS7..LPd:CMaR/NDG0O-J?.OD:/BTf\7^
/YMO/1O>O[Od?>IA4(L:\X@JI\O.d67BWgc&1Y.TgL)69PfMQgO&[-+AOGg+@&=J
TF.?Q_Cg.H&gM?d9d^76f0K9ER=8J5JP==8K21d8F1\5<-)d_>V5=75<,^dZ/?Q>
=?R9N51K&:[+AY1,XE+SKQ6<2\DaOUKeA(d^NL8=N#X@1\I3/X&aS6BW2_I89^:+
5XPX5ULbEM8JPCKW9L)==H/Q5=5C^WFLOA)Z42fC]M=BQ6G@Tbe:8?43gF((+b9J
(ZY]d-f)TbIE-5_#Q:L<5H(.;\CXAEZ)B0G]31bBG,MCd8bGM&dRD-F;<VFIE[R-
M:]AX?NaZ6M&RG>VRZH&Z3Hd9dV#,L[BZM_VOGN(>#Q429+W?SCdNc13>=McY&6[
0Bg;:(E>IKH.?L-ANE593H7E&\:)W7PPDdGOd@4BXaIBR]L849,2ff=[1Z4,GeLL
QH(cD_ScK3S_8??(g:5H,a2O-fa)/D5#8Va@W:F/Bg0>6L@Q-(Dd6-]+H/+&I3:J
W]VT2<e8a0-JXS1@(F(LES[\Q92U59IF4WXO7NfJYKF.0be2If&&;ZX=6<C\FQOW
L8RdTR8EeU<_3IP6<)5Q(cD7cGM=dSX0WLf&E;Q,YQZBcd&@_INe\H,#ZQ;d+GOa
-#;\QV?S4KT5>dP9-cL&C(T,0INLAH3Pge?++UG05&g7IY\TYV-1P8MWYRVcb1]Y
/Z^2X@CG(?)[E#Q0Edc\@^0>Y,-/^N0ZV=VedN-Td^5CeIH,33,J,H_E9Y5UOK08
O.fa9BFF=\4/+DfQ;&6LCaB@\5b?T;J947XM)7[CWBZ^N:bP?WK+6N4YROYEQ\fY
@>fR/STNZBM/6B]:P-QJa=@J(U:EL+9B3gY&&da;.U]1J</7AK321CNEO4Z)0Pg8
6G<Ng1-)9JQ?D[^>B,KFF#OfIK@JG>(Tb@ZZ<7Y;K_XXBcg-6)XKBFQSK^V&e_GP
C33#SOH\NT1M:AEG4(33G[eg([2Q=,MAb64f//9S#=U[<@>UR+BK[=5TSX6U:[V#
6UJJYYBEO>L7fED6O+J2g1EEKSFUEZ#3d5@M+NaHT1D@\L;?^OO<H=))eFJ&>78]
=P@7+\(UE/(X0AgQL&ZMOF,-a0HAOfAMOf1M)JZJ(@^O]<BB2+7AZ3a:Mf9L-O6;
0ELN7dT;Z)a2E>,OM57agP.AC=2FcXUDBAJ;GD5^X@]_ITPe.+Z;O(S&?E,fBM5L
-2@\geK<+=,CA&\KUXG#\AHVMVV1GQB/.Ze4=)CEdBZYBUa5G2IggXXa(:2VbaJ@
^LO\6[=\6VC=DY6.I4f)9^[O5)(USD?g3DXSSbaef;ZHaD@[[R_--DT^K?-Y:AL.
>P)3?Q)SU^1>\Xc7=1Z]AP^Y[bI[eESP@;Z_WQ^XM,N\UbSCaG@J34XUL13J+EAR
f,\PA#F;dQXQ.DfIEYITC\#;S\#YV&WX4\Y0JT:HZ@,#b8.UH34bMEY9])81QQgC
]O-/]T\-\GT:gBWe:XM^H95OOUd&GF?fO5U(=>@RR][YEAc;HJ,[M@8<MTaBX@UX
34DK4/IZ[eU2OPS_gVf7C)d+OM1^Y(ASLc2#Y.WP;8X#gY(ccNa3RXg.1M.XcHL[
Fe33MGQZb9E-)N--/2B<DR1e=CPT\=A+:cB&]_;485N1B4^_C;d[8^T6?:2T\(9F
]V]\@>KHW\a2Z_Q2K1]&aTeY/<@O(Y7ZD;CRd;WH<V<;W6Y+X<JC=3G351\54G9U
YIIPJO_)_.SfEJ#JK0+Ze.6,OF4_5I&c<P?3_@QaZMUTF?WVe?IM#--U?LA1MN#3
1&X_I.L\PEBIG8Y]Q35_6VK6/FIY3UKXAMMPeB.Ec6Z0NY?B4@=,MZLDUf\b?^=B
^-cV(2[gD;=P#?=&55;)@;-,\.K80f5+c(AZ=EF+-U-C^;KD<g+T2[O5WI]JKMH#
,E3[dOHX+BQaKfJbA3dWY,bHK\GK[_JcKE3OSYT:[<a;I2[L2;+,P:J7bDEDMaU,
L(>V<2Yc8Sd)9@,b#Jfd_WaAR2(77P?)A90P42-^<d;B=5&;@FDW/(G9g92>gfD3
]ZfOaIgOGM_^QZQ-&AcK3..@G1S&U.&&QL?9;74=+_QGSYZH^:9<d;2:&5[Q5RdB
LaE5(eFQ1IQ)E=Ofg@Wae=VCPU<P1a+T9\WdM+ESXP]A;N387H-QX4eTEOf/JHHN
4N07THW/4S@ZSKScCg620.H4dLHUH5J^1SP,ST(F.B#K#QPF?-442\a=SLI3&=TR
9GRE[/TSG9J1-VDU3E_N-OMeX;S>1UHSd8F#g/,@;WW^MaXV7dD?D7G4GY8\1fN(
:c]MFKHFXbcF293_MQGC#@&SD?4If9bc&g4PIT0MM@J\41@[UV1&ZA<JXBBZG3W=
7.T&_Xf-FBCXN2eZR#Bd-FRK&94[M8b]G5ZQ)Aa=e;^6Tg>S=cX&M-A@5e\Z,A/S
gfB8GDMG?F#I:61R3C,b0_;V40RN8aa#fLdC_/N^=[SPRTUHOB@5LM[C\=+0R-K+
3>c-A>VHeN8TO2D1\,]VN^g.O,_)\MEd\d1\Y=N.T;V)@Z9FNHR^3(><#GA+SHOe
E3T17d2;DUHNBXW<K[cXZGP1#F=LCQ.&@@dDW[.X0;-C+T<T:D@5W,XT>^\)^X5>
>c)DMH1Z>g9)K6^fZT,J.843?CWI1#A>D-e=Q.P=T0JcWCY\LZb^S?g;IN0Z@9Q[
7JCPZRVWV/M01S04F@E+cX=5-&aYGfMN-?JANDd5g-e7Oa,a6,70(a5)BAaF\Q[-
f@c=cWPSf(f^L,eGg6R04[I+\2V]IagKEGQH,Ac>XG=W,O)1#5G6?PIeYK6SF4T=
8JX^1BL4<9XB+dKc5-C0CX]J&;d&ZG<CU.+TDURKH5.KOHODF]TZH7M3YYb[R8;c
.,NBdSSN4]BNHFXH&E<^QBa0#N9Bb5B)(L<Z7OD@I.G/2YUM/F6VA)0_HFe?]0A=
\I7HH@/XcI6&&ZP@Y&NN3N63B;-,VAZVeW#f0][6>#,VY[Z;D163QEWP^1g54MbN
D+UccASSNV6@P?=[[(=De@30CHgX<\:d#2+eK&.(@Ug3a6a)ZGU:D)WVbcQO1TfV
JbZEZd#PA#7_N7/Y9.J041)fQ^TPcG0IF8+TXZSa]4#3ZSW+I-SbC2<9Rc]9ba^3
\/I@8a51ab6D9T191F4gFZYKF<Z1SL#g.:b(+C.GbZ4E>O)JY+,(L^/Z>H<FGb.R
L=)g>ff?&N[SS/3>5&4PGR>=-H9+g>\B]0IEFU--3W:H076JDb5/9X4ZZ[BWMAT?
D;#MXOPJ,?T9I3FN?T\6a3eENDT3^BgQOJV?2bM:TOU7TCBe/aHgJKIb+I->a6R]
F939R)#5]6TM&TW\V6X1Cb1UQ_.(1>[]ZV1ZY5(+L,7YD1:Q:;IW2,.2G:GdWdRF
MN51^MeGSW._E::IN)DdM];JSd5fHMFQ8VNA=1IdM)<S@5AHO0HCbYSE+X>UO/@e
5BePT3Z2CNAZJ_63:e&0JNa<(C=OFgbM,.QIT(cIKe;@G7=#77b02)65RGb(cU):
Q^@_aRDUg0<E(ZX1V9A12eB]EKL/03TB^9:1R/5,]9G0Saeb\(VXa7#P98V5=Q\,
&M1>=\;VJ:9>f5.cKE#U/cG#JAZZdBTb()^GSF;ELcZ9b0Pa8P,VfVOeR9R+L-ZX
[b\?63>#PcKB[^aREbGVf>a?X=\)/(5[c3e_]](V_?bIgFdWY))+LJDEb.-O>ZJR
d.\RU?aOM62;Wa#X2>SGcM22P)5R:cf6TEe?2(/beg+L/E7-4b@9&.1IDd<PX(A=
^7I9E&:J+,DeLJL#K?GRP6T;CMW5[A;gH@cBgCN9W.VZK>(1CWfB+0_?>VM5K.GR
(T(aC:_&2@#@d(_[P,SL?ecY6H.]_(f,P5TCW41KK-[Y2O9+g5WJ/I>=]06_DN)g
HVe-75(OZL@/RgLB?@\EL9daPK/&DbD>D?3E];AbN0VE)5-4ZY?W0W/e_)f]8gY\
#&U)1Kf&46a,ASL4Q\?<e4a\&F[9D2M6BQ1dYcT9-)(T26<0c;0g?82c4ed4/b>N
PZPD<RBDT(<-3Q@fM^LSR/6LI/KUdP:N51(5/cN8d[-Ab+&HGb8CO0dT3#33K0DE
.N01&6D[\F/A)\QbL3OJDR/&YDHREOBX@5eC6;a#2LA_,#@^6O2Z?ER^@RTfbUe-
\><C1fSVB,0/.;<g>9cU;JEFM9.64,NbB/Z&FUVV7b):.O34@;R=aDZ(2)#YVcM\
)>EQ7C]f_+2bYIa,Y1d7D+3#WRHY@6=Pfe#.?<=<,KEPdc^LU=V#0?=@<g]9>,;8
bG]@3YAU&NZBLM-89HD:NbFV#.B([DK5Q7OYD4A^_X]\KPWC@)/66;b/R<,N]:QX
fFSKK;NYLU_.#L=QX385dFKZHAZP)@OG>Ee?caM?D#b?8)9cfHH64VWQ?d+#O&,C
-1MR]Q,>HVU]Vd@TST>2aXI&Q6CC8+^Sf=BbX[@X>?DD7XF\F74E=^5>])Nd[,2e
8MZ=J7V,J2<f=K#[,9@=034C&LTVgN6TD,?\[g,0KIF[FDFDUK0:APZcDbJJdcGg
,_HCaVa1-6>UAF//;EUPIBNRgeWBD+,NeMB=0<_3;GX3bg8Ad6J]d/Y.7.?Je+O[
&Q,H.Nbc9]5Q>LC8S/AN5,NNC[d0-4#D-7]>T\XT2]MDKI,RgBQNgZ&,Z;/NETe[
e3@Q+BU4Ec,61RA^&;=K4cH320VQ=<TZ[Cf]FNAB\T(C=4;3@\VD8:e\9eGJO/C2
GCZF4QR?_0D[F9BbZBZaR\?2@J)EM90YB0LgN9FB7FFV2MC<FMN.?+UZ_MB7@e>@
1e8bT5a4XK_S<NJSedUC4ME2cUb(/E)<1aB9/4g5d/W,dP&,BZQ\F)E.FWEU=FW@
_G]>/Xe_+K(>6QD/2Ze1>J[@aE5c=R/FO/]bVSM[NS-7ZNC&[#S<-:8dD,>Le-g6
AKID+0]O?B><0P]YT++96-cOX+7_BX(7Cg4,KF]?K6JZ?I4)^:[6),d,M[4??b@]
4H#SHX_d-9S\7&3-)eOKCXTXF+9.Z]1ALSR&P<M2(#X@=8#c3^O^0b5\EMJG-E+d
\>V,A@XO-BBJ_e8J.B+RYR.-XK>.8,b@bZ-S)6_&CgHSL0^=];ccQ1HfV72A8X?Q
WFCH777EP/THIGU7_BBR?SM[(b^N9F>K_658;XG@@_eGIVXNRA-^:78YJIH(;-F&
?a23-eH1SbZZ=fa==8Y7gIG8(EX?;e1&[9\1E^D\@(11&8D^5G_)]e=+\OcV]].;
=P-HYTfBOgPA^2g#ZPCOK.45JW>+b4[H-HdY8e>T=fM_Vb.e]^UX=GQNT[:N[3Q;
.=WBR-Q^56>A/-adLMB9GQ8(d7>1E)_,C0_9O6+C^?,3S3ZOffBbU@fME1FHeHCV
^//D0Lg]FB;IPMLL+-5E@0-H[>SKN0CabOfK/G(:d9>TH9X&^SVT=J@QWA\c[\=c
2DQK4b5Mf.8T2)L<WM0Jf6=W&D,4]gCC)\V,POgGc2+[X48dSXZE8=9Je7GX4.<>
4JVPY/#,V(Y>Lbd6L#FIafDXYTd#9]XADOMG:Mg?/b9FN2.dL9)57)R>UeP?NV:I
BH-Bga5,dPaO48a7_@G+MN=Z4_A4X-(9R>QZ##,187N5#eI/G^::]]]gHR;Q0Ha7
>aP,EdFYOKPN95AJI\J/^@].[.7?+7A[K+MEFANRU-)8gZ4)H7cOYCW;)<d(6d><
NBMM02[O_YAGOG<RKd-0g.AY_/06;_.bUI^:c7>:N_0=?N+E&<fQ1@+<?g7OWaE&
74,1KEJcI8@V(6R5S#g.;EAPB-1.RRQU6FR5),7&5J[c4eHcL<4U_?&bJ6]526QM
+QD]I<#C5P568,V]XSa&f[(YeG(/E8#=;=.&D),6]80e(N[(:Y3U?QB>F\[6P@-\
_72(;6>)XUCc&J3geN0W\=)cW\Q@()dVA9JEBa=[I>\>&9c#K.+^#&cVAeJR19M0
&3XYW+CR4;6>gZ_e=Oa@S(BSHMRF?I<WW&<+ZBV&MccQd3J?1(CR9?7;U[5PeYGW
U&=gN2;C=PPVHDLI<CA/QGM-?^G1N^:G#fP;G9#KTM3-LZ,bZO(9[/1;[CKWBQZI
;N29IZK.;3T)&g1L/)LAIB#AJM/-07Z(GP4UW.b\U.XS?1IV;4DZbBM5NM^E5e?E
>H_L?6:8IWB+-NV3=JeNe^VQ0UW)T8cZMHE[<2^bCX,@NOWG:\S.Q,V@7V0&.BdN
cRR@?(SJ[PY[2F\b7MPF6fTf/Na_KF1JL7VR.aD7DCc&4G(:43J9V/4[UG>fKJII
I,dXUBXV[64.#]?4P,B,=^-BKUUTIfbOEP]VHdE=gQX947/JJ3&fXAX[@PR,PF7F
7THR+X?./+D+ZRH=&cCOEO>#XcMd>,@fXfc4I++U(ZO9_;M=H7YJWcGDLOaM&/W[
D8_Q\d.17\@6b5RdfY7^&;+X0YL[BC^+QNNFg:0dRVE?e@[Hf__DO-YUBYD]O@/@
MI26e>D;aO:;a=MCeS?Q:7DV-X:S:PDG6(<NH6SMG+=XX@8gIRHfSVWB>)CVc4)W
TLQ:f>CYf;[,84JI9EJPVc[5Nd>+JK[(afHZ)dYAIAI,e_#Y+]K-Q?7G4A]K>dQ.
VH]8>ReTY5XM)M35>g(F)&&PEKG(],PGXUEBWU,_3GKZ+A43cMaX6X:N12a-\N/+
G6-1_9LMLM/PSf[,#T\(b>3Q_.,-a&(0Q.P1\cK1[NA3RK;f:d_Y56bg.<f-&+C9
\(IG0;>14U]fIOa\_FbQ#NB[HQH<>,_JH&&\cPP<gJ5[8HeD+aD[Qc[PIM.b3\UM
[2ZAfFBW8>RN93^T663eKZ=\-@:\[]9^,J[Q?P?=>Ogg(&Q:7G<)3>V1>4+_aSP6
d@g\B<9?Db?&\H;EMc9QW#MQgC<?.R+[;3e=A]MfZ3V#N_:8d-C==&cBLD0Q21,&
+O=:5Z/C)_@TL0=YS+WJAR/S2GXWaLO6:=XRO?J.HFK;O3a]6X/7K.)#6WY=US<#
-Z5I#X:Ua8NfD<@dQ;Ub1.2Q&)V@M,+ZA@J@AO0IF77?)IRFX@5ST;^=#aH[<\g1
E8d6WA;=G#aJNWd_eMC;X?=IQZ/6MG?[/eSB7fcRVPBMCfX[KKWBE5TcK26<T,Q,
/:Z>8:=aA7ILI=3E,1I.^f2Rd#A:Ab3HMIdD_9dUM8#-:ECQG9/:g.cCRd3N90Ec
PH:c,P+G>&_TaK9#c+fMJQdKe7a45IR,;^-dX7OecOgD]5G.0dR(BOPg:]+,;IT]
(_BG8P]7,?-gO-LV8a)OKfbSN4A4,CgM)56EFdG&g=RgJ.a.,9g.DL?Y1/7Z+2)X
0:7J\Z#D0RaUT+>3cL#.QH0]C\Hc<.&-70P,KS-V-^(Ub>e490X/-,F2)N)&68YV
<aRGUDT<.L34+&ZS:UMdf#+f3d_Ra/]W-U#[,=R)Ycf\U9@YCOU#.,XC>NERLGg(
8:Tc;=a9feMTK23e;2F;(]:<X9XYZ1IE0Q/aRRQ1RVfLHG5H>gX1S&[e7?W3ZMdT
9GTf;,LXO\A>1f0:DbgeBNEBP?IRE07CP0BbDEH\4MZJ,#K(/M6T81JeS8J(V)@C
;0&:+@b.Cc4Y-4>NK(D/W;/KAL,TM2>4<P<DG_0g6E.?3SKG(D\2dV+D/d0CC8<<
a/U^@Qb9d)]RDT1D27MJ5IfYZ^21e7,T=[#=E.^YOJ=1;Y>cA/?AbT7OcL-@X](3
_+0b7[W:8GZL?-P?_N@WDc+]gYD0B3ODFDU3]UQ#(Q)@K^MXCZL?LM;623B_I(S4
FA[02U;V3208(c_=dJQSR(EP;V1.fR6BNZG<5+E&TeR_N^Me9V4eS)&V+DCX)=eI
(JV7?N])JX5,::bMF^->,c9=P/;<KLT2J:0FdLEC-4.JA4Y+ePa?A31SQLOW,J(c
<?e>Lb)G+ZgLMV^#=9BUgRe05C#\^9X&;;2g3ec-::EQ=#I<0/eZ&GT<TIbHF9=\
4/Z>3(V]@MZI>?FQ@&RU4U[_8@2aHfP&((a9G+8#UdCN][,Ja:E.eb<OV>S-O_d^
9e3^GI<D(NTfEUG@c(+#R?MR:8Og6)GcY+P(L8cNHBA/+:+K#Y=XK93?6QbBG2bA
V5,T<(\;e:=#92\H5,HVTf2b>7GgZA,cD2<<T55PWeXDCU1eE=XaGDAHW#)S/<QT
7.7##GA,B[.YAP0]7+F^7HBHgM3V78_6eaZCV1/063cP+3>I1UNDXf<+19Ga2M__
XAgR^LC^K]+K;;:,\(ga2&PN\?G[cdQ5<<dc9KV4b>[dQ48c^478B0WULJSB53H@
8I(V<JBbA28Q3EPOE_9]72VD50\#25GN39#T3X9cO1]?B(3;\OEOY5+VF-;9f:J^
6[F&>/-IT1ED,J^87W0&PE_PQ)7XgMg7TC(UDK(T0PR,67>S;c>+?L:)HUYHPUOB
gbPbK<;PJ>(:<82[f;Ja^ONJb-OfOT-?,FP:e,M]<3A?M1e?ZKFZ-3@^[4_3,XI2
SSQ\g.F<O[d0[O.JX;[0KJeWV89+@J/dGJTd=YHMM^U24G20]a#UCVK6bgM&\+>@
Jb7bIfJZX-2A-V6#)7S@eZJV=E1_BK_a/Q48;.Je;5fE)T?]=Y-dO)NP#22C=GS5
c1#X3a/;-0H9/+OS^\/4ZeCcbG1_cX21,M@;15A:]\PI90KOA:L/#5EdPQXN2a7:
\L@<Ie5[#CAOJ71N[EO>I)D=2QIX4L_?/L4I<L#5H--7:V/\LBT70Lf<&ZD(W)#1
6LAaf^]KG_M-]T:XPBC2E/3Y@O,8Ra&:FUE8XX[?#bO6edNN^JE507VM8DW-K&ba
R&K[eJVfAZ.-,T#f([7=81\HV779H-D]]134YTH#:-PW^g0G/K@:,XH.E<SG-3Td
0CMW9WW_X5(-ZPS_IYg0gSW[KCgS)Z(PZ?2dTOKcZ:>8Q\B(R-/18eQ-_B=5C+ET
\8a]A)Jgg9JBBPL[^OI#P/WD0W8LUg/bR9/:1?/(D+_WD7EHdUS[4_ZIB/T0L1\-
L88fFUY-Z\9DU+46VG65W>eSBXPJ;Y2=.K6REX[g)7c1/IJ[^1[,Q3L34/b6K.DW
DbIM#0a^]GX,9IH0W^)=1QCAeSBM(-@?)@C5<gK2\JFO?Q#.B48G=8ZZFX,2SI(#
9U5f2Q,MY0KG\K/Y4#^:ELJb5UD-;KHd0WS6#-+0]JS6Vd(]CQ71_b-0,QMaH6SB
J@cSOFY5OJ+O>9>0LP)[_1J,;QAG0M_[[X<^VNIf6_OYZd1WNA]LgMO(H>?+05T-
:=)KA9IGN#5K,6Kf\+a-C[C8]QO+TA02G63bcYW9XRd@_XM79PT4CcU-2LD7X?ea
N/Pb90@cd#E(T=fWYU8&V=@^J>P=fd8U]L:K4=V_O06+)MYc,VR52[BAG;O^^<\H
K88>J\@,-AaAL,N7,M=dYWDS0cA9@B=B9gOQOTK4T(LK.?eQaB/BaEZOF8F0Bg3N
b^geNeWaRIQ+;J,/[ED,UA;&C<^,\E4HV\?/Q4#1bO0(42X/:#2;5_gQ?-a/2YO/
KB,L)NG0P7^-d0@17UDc=-WabK\;0P0];;GHB#\fI+(<(9,7M[KR29O/3@\NGU:0
^R:3D1_&-@L&fbKS0=[[[be#/L]Gf76/V&]\SJTW2Y;?f^XcAV2F8P2&J#3eZP4d
7[)eeXDd9MK5LHf8VRA1D5+B-0d@OV(/^\>[_]5;6)e;-?d40N@.Y2KfH/VG4QQ1
B<3EW^H)5dO6C;X#KBAT)b7^4BYB@RJXY?ab:-^NR3&CY7J7H7IFcO;IOQT4\^YE
6#F?<XI^[G0^MK=(H.c;##.[\WGT+@R#GPeBEa^BOEdUY(,CI<@24E=O>Y.a>/T=
&>]4X])9M2D=&-[SF;B^Ea=#4?_JKNLF2E6LR+2T^QRJ(_?:2ND.Na@cC,/Vd6HT
^e^W0A5gPBZ>837VEf(?,cRP#4B-bS<Ha[^eE[4KLE(X4]aSXK15^#KU#P,Df9#2
H3>P0+KCWA[AZG4@]\15\TAGA->dF4<)GcY]LM[&9d@EVENDH>4,#R8B[M1_Jd;P
X+CgW-KA.FG5_I)ZSGMOV4H:GG@@I2IG:Q]]Z(;B8e:C3\0d&@af<U[^[=3SSBHP
PT.)G8YN50(dB[4SdXC4??7a4.?GTFM]R)LFIW+A)C;^1?[D=]YU]H&#-<Bd4cU[
Kc8ce:&M4&e^&W?+WF5R9@B\TZPOR3DE(C7<\A[:W+bKOS=A&M4H2?,->eKVB/KP
Acg+MI7TGPSD@7V7#]^IC[W/4H7DN-C[JDP]T0@g&f/L?\1E<(?ILOT,[:TESU(2
:Egb<O)4W5U-\ONE-b_.X5.:4(f;WN;8\Fd=N;],IL;B4bBb@T[XGVKbZ<[E57+8
e(DXG/(8BNK]Z(S&X842#;&0L1Pf<a<O=+d2]W7100E<>->db,[XIY<BJX5a>^@D
31S01I&DBg2>+],\9#2,=A8[ZB_\@(.\)?G7SPDBfY>\Y,d=2^Tc3cS_CJ)CgJG\
//_C9T<-dG9)Y(dQDRfSABHSAgIA[DB.-eP]b><f95/]O_gMU<PQX:SU./8b+\+(
bDI&-dX39f#aI7^#F)TdJ58I#AS<V1QTYU#W\#He]&<U3?W/1_Z<CRMH+eW)cHZO
DEPY6_7:86;Y[]@.GV.gMWY.W^aII)#4>E_7LGQ02PW(\TAbf<C_g6J(9QYQ(KKF
f;a.K,DRcY:14-8W<&-5IT1U58Rf@-f>9IA+636DEBLgUdUbH<1RW[-27f/BbU>@
4\4+=YQHGE931<W-2Q.)f06QT(]7Z;-BLA>N5YcBZYgMZNO@JBI;8L4If9#4FPWd
:]PDR]dObHEd<O;0gcd52&2W&Jg[2?F&+-_(>(TI(a1=HN3cHF89(&+2>NOI.[J;
LHSZ/C)B3MY8-0,L+c(OF-e;/e_]B:,VYB7E3EbK>P6EWK&4>#<e2CCJ23Ga.VBT
AaPV/2cd3KFb1N4+7OO2>]U,UQ]-:MI&&T(-UeXa=[#;6+[W^C<.B4T??A(76e&D
Fb=Z]A208+_5T#fMZ[07#EfacaTV;SQ#]9KL)5RCD(J9DJ/T+>CN+VY-]=)KB5L<
<T/?.69ABKaBSGV-D,TDbOGVI(OCOOc3)8Mb8RH<;fSJ.,X0Q=1\gYCPU[+),F^R
WE.f#A(1G,c^<^6Zf1&FGH>WB9(dXTfV&,SQ9+<8g.g<dWcb&,XB12/>B6Se7<cC
H_2NbC9]&+EMO@/C,@V]D#C<81e/Cf&<>L]RP8bM?CB[YN0_YUgK@D6K&MAWdZ7b
2dW?C)U[+4ccH-E@2I1J9SY0,.d+R;dSE]:(<cZT7bG;D7MB\_b-Xg&NW<X2+C51
eUU>_VZFaV)g2)?:=GZ5AQWYO06KNa>ScE]#W,_Ce_/R^-U.LJ\)T[Y@[M[2LX(@
/<OBfdD<)B@AJ,LE/B&>:KZ1.WGDMbH3Ud:+W=-/40>U;J=LESH[#0GeA5[XHR6O
?I3;f?EOD-.CL:YJOMZUBEWJN;2fbRL)eA)fO,(_:G.,<d/bL-;SVZKe_A/aH0<N
OWH73[Vc>.JTUJf6#7#JNQ\dO&#aaO)=8aKB.NT[@G^(+P4+cG2]8VZaWgFVe/aG
V0\A(=-9R//X8f,\Y10S#.ZWXJ9)2bI>)XD.VR<EEMF-#)3HY,#PVI/?A<&,DQ1C
)SSa\:0UfcC.+,IRZTAC<4&C:E3TB-1)V;H1P2GE@,1+G&QFJJ&&4f[_T9Z@GQMD
#@\@A^gY:@DDC6-A@(dPgcLIb4RHXI<5Z#RWc++;7S)(>:+,T1R\6KJ>-FV5Q/\7
K-b4\[O[D<I-D7I#^fA6VAO](5Cdf]HVbfF&]=>X_>2e.gG:f&C4IIA?cCPS+)NC
B@H\VB)YcA8_VdT3JH[MLQ,G@IEXA^6=&+eW2fTHZ7U\cHZKE1193:(/;bILa?#:
Q,C^?)dL?6T3)ed?[dSB)3d1#YJ)GHe910?RF?MbTO8K6;D&fbAX+H#TD=Tc/]dB
.179Y3@@X>Vf1^OD\7Wb\M,O<OXPgL)@?MNMP9-2.G+JGKU[1V=7W,_>C@=,HIEO
X3gBNGW<,(.,A0F#KL=1D?(8a\c@ed@[7.a])2B@.L/862-D-[:J@D(7dII9=U7d
+C_Ge].;ANO+g2-2R_(R-DK]6f&.X(58N\LTC[fE.QUGFPPbA,:H(>I82GG\\&S8
AQ\>KUW3<4\-FUK;fE\X7,_aIXI2205\.0\>#,699F&&VP)>FY);)C_>T)XQ--TD
IDg>6TE=2dC3486,R;FP.?:5:Ue6^Wd/O0X0QT496R;)#@9(I_,.?>CBGENJF0Y=
HSc]HDRUG4LW#F)ZBL,T?LEaeNM2Bf6/OH>.b7C81,eKWEfIJS9RVR3d]Z@G_K\Y
gP&JK=T_4S&^A_a_8JDU#Kb\2>T&eI4P^;ZZS6b@&N#.3c\;[H5.4^T,0beR\>D]
)3]X+,VXV7I)T;PL6/BTgMY8A(BNXSD4E[)5T.Y;Ne:3\aJSDB?7KQI&&G3dI;aB
0bDXTI\f/SP&IWIHQMY>(BgRJIMd)_/UN/M4A=g4;(::dC?8:#7).F1bP0[9]d;\
OFXZ<e#3?X]WYF\EIH^=(=M&1-@Z^UQ#0D&UCY9;fbD(LOAIfc2?8-Zf]4ZDP4.V
F#OfHQ,^I,NAb2)YB,dR5\\G2cbX,OXb+7T)#K,1PG?BT7VA=5:YP2NU:EK4&@L9
&-_=<X\&HcXgaPeW1WDIJG(1-51#>4&.50A-7TO&^RIT:[;O4:?S:WIa^#R>P(P#
_W0=I+[@g]+IS/=0K:(g^@I(KEQ?GO+&dJ>]+C(Ma;d5XcSZ>A&5Z;c;/Z?YPJ?X
OC=B5O=(OYTQHcM[SM8b8V@g/P:;;f9DfI4]9T@\#3;16K,1#LgQ&9c/.7FgDS84
C_]=)cfUV,V9I9W=B1S=OUDOHY=C[gUTS,3J+DY^]KL8&AXdLP@_RPIeLMZ_d;A[
X00:GS>FJ\d.\0Qb7f<Y=1(=4[:4MRWF9U/AB9[<TQ-Z4W0)Q2V<1M9b@HH/\O3Z
<SX91^-3^gX^2M[Q-\:-bg:<I>f/aQe,.@EDc@W;>APEf?DBXgVd47R;1_:^\AUJ
.;TO)UVdIAMeK^?/F-34ZWRN,JA9(.;V_8=):d>c/HSV]I<LVg#2/BL6^7e>6)4/
4:AEg@d)2YC7[15[ROZ+B<?df.cAG?(>LaT?1T9PS48=N5E+6g@<G:?N2-UB#,X_
@G8.&E6TB7.VHRD?&<OWHMHN_(F<34Me,HV^J<G&LNc6gd,2Yg.f-/YLR5GPgVFV
.^JWUW#D&N]I&cSTE+YR5;:Y]+,:OB[M@7E;0V,BL<b&M8]#-1&ESdd2H3DQZ[QC
aX<\/4F5\FaLC<PA@YDbK&MY6#ON&/C0IUXZ,gNEFbV;d41MRXg^F.11Q09dQU2S
/?5XB/X.dI=BO5V.]aZ3LfZ>E2H;@+KUcPD?B+H.Z-0g#fMEM#JP/5QJ[]F\;M9H
f]]b^2Z=fV_SI.8PObEXTR?5W>M7MKYO4_/HCU[B5GJ]JM2IVD(fVdZ<#L2J9-dY
a6LM?B6[f6J5g+0]cJ47.6>AQJEHfE1F/9Z74ec]13,c[/@WZc2bd0cXB5-1/1QR
g?MM9&YOMgb+^+5f7M<CS5A(\E6=Dg6fLcHU>MdWccDb(6&Z0dg+;;P9]RN(</-0
dZZO61(O)I?VIS7cgSJFNGEJJ2W@_SF?203f,-g?FM\/6LCVJO\BbZ8BbQUM:MI^
7\B_f57HKH)A7cN>-2Z<KSS3?d=35[R@1U[##3(6)-SNQXC)O8Z=3]RPZI97-0R9
L<GN9OOF94FBIbK<:4^JM8[X[,S<SE9>:6:U5e06)Q-&+W=7HJN8f.OI.@;X.?<>
,WUJLY1\6<F=Nc2,[b3dR-S0S,>&@UQ+0g(Aa4A@6<F[.XYT/S5DW_0McaS_&COS
Z9cK1C,^V@CX^YSN\CA03>#fZTR_Z^Fe>V7VH5<9;)]KfP:M>gJW1#/(bD;/a:_V
Veg9)BX?Z?_C:;[Q5Mc-58F</3ZSPPIN+AR.L;QLBe8G3K6(H2E[?9D?[dH8EIC7
D[MAPWT1<B_:3YC,8bO6d=0<6dGbBKP6G+eFX)&9,:2fe;#e>PCJDeSTgNNdYf#F
f_C_9OPYcTMe1HI7D>d3[PZ8:8a6H5DZe]NGU&U>]7I(b01\O(Y>CBA1^H^FZE/Q
KV)d:f4+,,0^5(_f#)If053NJ3#-M8b,<K:4FeF:&aI6A>XW2?A<dLdd+&=aG^;P
LBUIEe4P(@BGYfff3:>DL[;aGKWE17MGPa]e(0.CRNJ0bX/+/7Wd-NB0CHMOMeP6
;7N<OLZ4M-fHTMJ1U9&C?X0a7:#:VB0Ma;d(eT,X;JRSQ31O(KVdS;QdC7(_.2X7
Z+W4X:6;01J1O;1-<QFX^BSPe_\#U,O/;TA>g]?PZeg44AMeOdOC^>cC.#(4<cWJ
fI+<^G\ae#Y9]Da8-g=Y=GdKI:ZPdPb4UgW43b<Z+Y2[D-3?V3RG0fbAXQ_QgYcQ
gdQ?QX#A;gZ2G74-E+6VYTRPIW_?<YNX,:G[Q&5WGB&Z3;G;8IZ253R:Y0+MO#Z+
gC(;VH#MbP5<B/0d4?EHOR1bM#?PIdS:,T7F/#,ITPK4#])@gOc@/FHLK5[>G)2-
#<bIIVT3\1^.R:,8[2K=9<)B,XD?J6FZ+/7&(7S]XUc##(F4[E(NELYGYc:4B0aO
MF3W?>[1:9gL(5CVD1<=DVPO@&K(d68KVM646LdMH?fRGCd(GM31D,QEHI4BN_)@
3^XVgYdXI478=3.[-M/OHKfIc6YVDd.f?^b>OF-:]P98dX1=OV3A#^GaPMd[BabO
\YICM3KPJC:S<<QC\T4WZ2W@e;8fG>C=XVU>84H>][I<U]R71P4aa[U>1>G,R4?g
=OU:[8fQ?+@N2.#e^>a>C/-GSBHPEE3D>T.0G2-#eE8BJDBNaJa8OB[])Q)EHac5
XUL)K;_YL8^AbFOVAgR2CGT+DR5dN:=#81^f5JP^[fO\?<PLE?0>M&ANDJ=J<FWb
Yfg&5NGZ#PC.J1]Z)DW92RN^B:4^T6e3NAbM.#7e)R:KY,ZY+AO]CaAGD.BV&6)+
IC&F2BJZP?#:JZXH4?^S3c-UcG&O&fEMYf=WHKB4\)@#YP>K-aOc(\QHAZP#TS&P
(Ge(<4.Zf\GK#XW_WY(,EHKCJ;7G9,Zd=6:cP[-8O]bFVYXAD@SK^.;=bSGS7)OY
DA[AdI&TKbCgKa@7(YJ0d_++JNcK-/6&PF9R@.W9C^HFF$
`endprotected


`endif // GUARD_SVT_AXI_SLAVE_MONITOR_CMD_UVM_SV
