
`ifndef GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV

`protected
(?>9>PAHLDY?VRe#LY8:RLX606.f3aO)+K?R38-AT(8D6G/c8O?G,)Ka#^<0&1##
>=&<2\;ND?G]\;PG,SZ12GHaTQ->S0NLbH?_-/J.a_5A+_?DQ4]DOW+7&Odf,5.7
g[6DAQ=+KdJ(b73g[_2?X+O/-OXU@V:\]<DD&a,RO6E=RG06+H6B=U\+FF7SF@d]
(7R+G4>PP<Kc,VCUfd;cR(WP_.f)dZ?:SJPbXCG_[7Nf-^SN46.&\Fb8+0-6<VNB
<S^+1cB7J^##FegUUGTR=H3]GR0J(:b\W>>LAE8V=FJ)>?4YUbMed9W1]N;:Wg&D
3d#Z,4-SCSP2<FH#fcOI&cZ.^OGac(#]DbHGH6MQcH:]dNILTO])c&DZB^)NCYIg
]SO.b]W<-N3I\<&V.cS/^Ob._@NK&_2M8&R=b2N::)5;@SaEKZa9Y0T>&/LDU_+b
BE&FDXDP=c(/c#Z^+_;S69=XRT(ae3,,BD)WLPEKdFJ,K(gC0=LMW-U1d]2D7,d:
/G2XQ2g<fW4ES;UO7N+SDCb@_1ZA:\We=aJ4M1#dO;RXK5A(3O[O)\H1)<5?LXLE
1U8cAB7Q/c>.EdT_UC2f(93>;IY]R]J]H_BgH2&V34H_I58VSGEe[57_MF]&3bGe
0=2TPW3GZ#GE3T5D=:;4/):+A-DJ@8:[V8f0,_X2G)CaI8dBf<H:I<RHWYMaW;6B
0G3LK6Z^d5e2<:-cT5PIOb\TEU#(O)<U:VB476W:0QL>#\WCJMDe2-c5678D&T6O
e?bI#89><e=1B9a2+7Ra?C)f&ED44A[T;9VMU>?,,9RTKg/^3<0JJ(A/YFZ<K=\-
;1B<Z4c),f.ReH5@U><=Q=g-[1-]3N;]FF,^(#Oe(]I.JX;C@W-9]4:bc<RST3E,
=I&(DU70L[4R0$
`endprotected


/**
 * System configuration class contains configuration information about the entire AHB
 * system
*/
class svt_ahb_system_configuration extends svt_configuration;

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************

  /** Custom type definition for virtual AHB interface */
`ifndef __SVDOC__
  typedef virtual svt_ahb_if AHB_IF;
`endif // __SVDOC__

  // ****************************************************************************
`ifndef __SVDOC__
  typedef virtual svt_ahb_master_if AHB_MASTER_IF;
`endif // __SVDOC__

  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Port interface */
  AHB_MASTER_IF master_if;
`endif

  /**
    @grouphdr ahb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr ahb_master_slave_config Master and slave configuration
    This group contains attributes which are used to configure masters and slaves within the system
    */

  /**
    @grouphdr ahb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */
   
   /**
   * Enumerated types that tells ERROR response handling policy for AHB Master.
   */
  typedef enum {
     CONTINUE_ON_ERROR = `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will not insert an IDLE during the second cycle of an ERROR response */
     CONTINUE_ON_ERROR_WITH_IDLE= `SVT_AHB_CONFIGURATION_CONTINUE_ON_ERROR_WITH_IDLE, /**< Master continues with the remaining transfers in a burst after receiving an ERROR response. This mode will insert an IDLE during the second cycle of an ERROR response.This mode is not yet supported */
     ABORT_ON_ERROR = `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR, /**< Master will abort the burst after receiving an ERROR response. Master will not rebuild the transaction*/ 
     ABORT_ON_ERROR_WITH_REBUILD= `SVT_AHB_CONFIGURATION_ABORT_ON_ERROR_WITH_REBUILD /**< Master will abort the burst after receiving an ERROR response. Master will rebuild the transaction again from the beat which got an ERROR response.This mode is not yet supported*/
  } error_response_policy_enum;

  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /** 
  *  Enumerated types that defines maximum address boundary limit for a given burst transfer.
  */
  typedef enum {
    ONE_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1KB,
    TWO_KB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2KB,
    FOUR_KB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4KB,
    EIGHT_KB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8KB,
    SIXTEEN_KB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16KB,
    THIRTY_TWO_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32KB,
    SIXTY_FOUR_KB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64KB,
    ONE_TWENTY_EIGHT_KB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128KB,
    TWO_FIFTY_SIX_KB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256KB,
    FIVE_TWELVE_KB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512KB,
    
    ONE_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1MB,
    TWO_MB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2MB,
    FOUR_MB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4MB,
    EIGHT_MB =           `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_8MB,
    SIXTEEN_MB=          `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_16MB,
    THIRTY_TWO_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_32MB,
    SIXTY_FOUR_MB=       `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_64MB,
    ONE_TWENTY_EIGHT_MB= `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_128MB,
    TWO_FIFTY_SIX_MB =   `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_256MB,
    FIVE_TWELVE_MB =     `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_512MB, 

    ONE_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_1GB,
    TWO_GB =             `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_2GB,
    FOUR_GB =            `SVT_AHB_CONFIGURATION_BURST_BOUNDARY_LIMIT_4GB
  } max_addr_boundary_limit_enum;

  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This is not yet supported. <br>
    This group contains attributes which are used to configure bus within the system
    */
`else  
   /**
    @grouphdr ahb_bus_sys_config Bus configuration
    This group contains attributes which are used to configure bus within the system
    */
`endif  
  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  AHB_IF ahb_if;
`endif

  /**
    * @groupname ahb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_ahb_system_configuration array in
    * svt_amba_system_configuration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple ahb systems
    * This property is automaically set by VIP and must not be assigned by the
    * user.
    */ 
  int system_id = 0;

  /** 
    * @groupname ahb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

  /** 
    * @groupname reset
    * This parameter indicates whether a common reset should be used
    * for all the components in the system or not.
    * When set, a common reset supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to use the same reset signal.
    * When not set, the user needs to supply a reset for each of the
    * port level interfaces. This mode is useful when some components
    * need to be reset at a different time from other
    * components in the system.
    */
  bit common_reset_mode = 1;
  
`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;

  /** 
   * @groupname ahb_bus_sys_config
   * This is not yet supported. <br>
   * Determines if a VIP bus should be instantiated
   */
`else
  /** 
   * @groupname ahb_bus_sys_config
   * Determines if a VIP bus should be instantiated
   */
`endif
  bit use_bus = 0;


  /** @cond PRIVATE */ 
  // This is made private due to known limitations. It should be made public once the STAR 9000993130 is fixed
  /**
    * @groupname ahb_generic_sys_config 
    * Defines maximum address boundary limit for a given burst transfer in terms of 2's power.
    * Default value is ONE_KB=10 (here 10 indicates the 2's power ie 2^10=1024=1KB).User can define maximum value upto 4GB.
    * This feature is applicable to Active/Passive AHB Master and Slave Components 
    */
  max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB;
  /** @endcond */

  /**
   * @groupname ahb_generic_sys_config
   * Enables system monitor
   */
  bit system_monitor_enable = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * When set to '1', enables system level coverage.All covergroups enabled
    * by system_ahb_*_enable are created only if this bit is set.
    * Applicable if #system_monitor_enable=1
    * <b>type:</b> Static 
    */
  bit system_coverage_enable = 1;  

  /**
    * @groupname ahb_coverage_protocol_checks_system
    * Enables system level protocol checks coverage. 
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_coverage_enable= 0;

  /**
    * @groupname ahb_coverage_protocol_checks
    * When set to '1', enables coverage for system level positive protocol checks
    * When set to '1', enables positive protocol checks coverage.
    * When set to '0', enables negative protocol checks coverage.
    * <b>type:</b> Static 
    */
  bit pass_check_cov = 1;

  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to UVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env
    *
    * When set, performance summary report of transactions are printed by the system env
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to OVM_HIGH or above.
    */
  bit display_perf_summary_report= 0;
`else
  /**
    * @groupname ahb_generic_sys_config
    * Controls display of performance summary report of transactions by the system env 
    *
    * When set, performance summary report of transactions are printed by the system env 
    * when verbosity is set to NOTE or below.
    *
    * When unset, performance summary report of transactions are printed by the system
    * env when verbosity is set to DEBUG or above. 
    */
  bit display_perf_summary_report= 0;
`endif
    
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. When true, turns on the 
   * AHB Lite mode 
   * for AMBA AHB models. Lite mode has only one AHB Master and one or more AHB Slaves. 
   * It does not support SPLIT and RETRY.
  */
  bit ahb_lite = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * When set to 1, enables AHB-3.0 features as per ARM IHI 0033A.
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb3 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * AHB Lite MultiLayer Mode for AMBA AHB models. 
   * AHB Lite Multilayer mode has multiple AHB Lite Master and one or more AHB Slaves.
   * When set to '1', will enable connection of more than one AHB Lite Master in a Single System Env.
  */
  bit ahb_lite_multilayer = 0 ;
  
  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will enable AMBA 5 AHB protocol features as per ARM IHI ID102715
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit ahb5 = 0 ;

  /**
   * @groupname ahb_master_slave_config
   * Used by the AHB monitor, master, and slave interfaces. 
   * When set to '1', will consider / drive the BUSY cycle only with HREADY
   * being HIGH for AHB3 / AHB5 mode
   * Applicable to Active and Passive Master and Slave
   * Configuration type: Static
  */
  bit count_busy_only_during_hready_high = 0 ;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname ahb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname ahb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_masters.
   */
  rand svt_ahb_master_configuration master_cfg[];

  /** 
    * @groupname ahb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_ahb_system_configuration::num_slaves.
    */
  rand svt_ahb_slave_configuration slave_cfg[];

`ifdef SVT_VMM_TECHNOLOGY
   /** 
    * @groupname ahb_bus_sys_config
    * This is not yet supported. <br>
    * Holds configuration of the bus group in the system.
    */
`else
   /** 
    * @groupname ahb_bus_sys_config
    * Holds configuration of the bus ENV in the system.
    */
`endif  
  rand svt_ahb_bus_configuration bus_cfg;
 
  /**
    * @groupname ahb_addr_map
    * Address map for the slave components. This is used by system monitor for
    * performing system checks. This member is initialized through method
    * #set_addr_range.
    */
  svt_ahb_slave_addr_range slave_addr_ranges[];

   /**
    * @groupname ahb_addr_map
    * Enables mapping of two or more slaves to the same address range.  If two or more
    * slaves are mapped to the same address range through the set_addr_range
    * method and this bit is set, no warning is issued. Also, routing checks in
    * system monitor take into account the fact that a transaction initiated at
    * a master could be routed to any of these slaves.  A given address range
    * can be shared between multiple slaves, but the entire address range must
    * be shared. Note that this doesn't necessarily mean that the entire
    * address map of a slave needs to be shared with another slave. It only
    * means that an address range which lies within the address map of a slave
    * and which is shared with another slave, must be shared in its entirety
    * and not partially. This is possible because the set_addr_range method
    * allows the user to set multiple address ranges for the same slave. 
    * For example, consider two slaves S0 and S1, where S0's address map is
    * from 0-8K and S1's address map is from 4K-12K. The 4K-8K address range
    * overlaps between the two slaves.  The address map can be configured as
    * follows: <br>
    * set_addr_range(0,'h0,'h1000); //0-4K configured for slave 0 <br>
    * set_addr_range(0, 'h1001, 'h2000); //4K-8K configured for slave 0 <br>
    * set_addr_range(1, 'h1001, 'h2000); //4K-8K configured for slave 1 overlaps with slave 0 <br>
    * set_addr_range(1,'h20001, 'h3000); //8K-12K configured for slave 1. <br>
    *
    * Note that the VIP does not manage shared memory of slaves that have
    * overlapping addresses.  This needs to be managed by the testbench to
    * ensure that data integrity checks in the system monitor work correctly.
    * This can be done by passing the same instance of svt_mem from the
    * testbench to the slave agents that share memory. Refer to
    * tb_amba_svt_uvm_basic_sys example for usage. <br>
    *
    * If this bit is unset, a warning is issued when setting slaves with
    * overlapping addresses. In such a case, routing checks do not take into
    * account the fact that a transaction could be routed to any of these slaves
    * which may result in routing check failure. <br>
    *
    * Configuration type: Static 
    */
  rand bit allow_slaves_with_overlapping_addr = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 0.
   * Used by the AHB master, slave, and monitor interfaces. Used to disable HLOCK and HMASTLOCK
   * related checks when AHB locked transaction feature is not used in the design. When true,
   * HLOCK and HMASTLOCK related checks are disabled; when false, the checks are enabled.
   */
  bit disable_locked_transaction_support = 0;

  /**
   * @groupname ahb_master_slave_config
   * Default value is 1.
   * Used by the AHB master, slave, and monitor interfaces.  Sets bus endianness. When
   * false, the bus is treated as big endian; when true, the bus is treated as little
   * endian
   */
  rand bit little_endian = 1;

  /** 
    * @groupname ahb_generic_sys_config
    * Array of the masters that are participating in sequences to drive
    * transactions.   This property is used by virtual sequences to decide
    * which masters to drive traffic on.  An index in this array corresponds to
    * the index of the master in slave_cfg. A value of 1 indicates that the
    * master in that index is participating. A value of 0 indicates that the
    * master in that index is not participating. An empty array implies that
    * all masters are participating.
    */
   bit participating_masters[];

  /** 
   * @groupname ahb_generic_sys_config
   * Array of the slaves that are participating in sequences to drive
   * transactions.   This property is used by virtual sequences to decide
   * which slaves to drive traffic on.  An index in this array corresponds to
   * the index of the slave in slave_cfg. A value of 1 indicates that the
   * slave in that index is participating. A value of 0 indicates that the
   * slave in that index is not participating. An empty array implies that
   * all slaves are participating.
   */
   bit participating_slaves[];

  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Defines master number assigned as default master. <br>
   * The default master is granted the bus when none of the masters in the system
   * are requesting the access to the bus. Usually the bus master which is most 
   * likely to request the bus is made the default master.
   */
  rand int default_master = 0;

  
  /**
   * @groupname ahb_generic_sys_config
   * Default value is 0.
   * Used by the AHB bus. Master number assigned to be the dummy master. <br>
   * The Dummy Master is a built-in bus Master model that only performs IDLE
   * transfers. In the AHB Bus VIP, the Dummy Master is required. The Dummy 
   * Master is granted whenever there are no other Masters that can be granted 
   * to the System Bus. Following are the cases where the Arbiter must grant the 
   * System Bus to the Dummy Master: 
   * - When a Split response is given to a locked transfer 
   * - When a Split response is given and all other Masters have already been split
   * .
   * A Dummy master can also be the default master.
   */
  rand int dummy_master = 0;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for all the AHB Masters present
   * in the system, when svt_ahb_system_configuration::master_error_response_policy[]
   * is not programmed; that is when size of this array is zero. 
   * In such case, the setting of this attribute is applicable for all the masters. <br>
   * This configuration parameter supports the following values:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * This configuration parameter does not yet support the following values:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receiving an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static
   */
  rand error_response_policy_enum error_response_policy = ABORT_ON_ERROR;

  /**
   * @groupname ahb_generic_sys_config 
   * Defines the ERROR response handling policy for each of the AHB Masters present
   * in the system. <br>
   * Programming this array allows different masters in the system to have different
   * settings for error response policy. <br>
   * Note that when this array size is zero, the setting of
   * svt_ahb_system_configuration::error_response_policy will be used. <br>
   * Each element of this array supports the following settings:
   * - ABORT_ON_ERROR (default) Abort transaction on receiving ERROR response.
   *   Master will not rebuild the transaction.
   * - CONTINUE_ON_ERROR Continues with the remaining transfers in a burst after 
   *   receiving an ERROR response. This mode will not insert an IDLE during the
   *   second cycle of an ERROR response.
   * .
   * The following settings are not yet supported:
   * - CONTINUE_ON_ERROR_WITH_IDLE Continues with the remaining transfers in a 
   *   burst after receivin an ERROR response. This mode will insert an IDLE 
   *   during the second cycle of an ERROR response. 
   * - ABORT_ON_ERROR_WITH_REBUILD Abort the burst after receiving an ERROR 
   *   response. Master will rebuild the transaction again from the beat 
   *   which got an ERROR response.
   * .
   * Configuration Type: Static <br>
   * Usage: 
   * - Size the attribute to match to number of masters in the system:
   *   sys_cfg.master_error_response_policy = new[sys_cfg.num_masters];
   * - Program the error response policy settings for each of the masters:
   *   sys_cfg.master_error_response_policy[0] = svt_ahb_system_configuration::ABORT_ON_ERROR; <br>
   *   sys_cfg.master_error_response_policy[1] = svt_ahb_system_configuration::CONTINUE_ON_ERROR;
   * .
   * Note that this is used by master, slave and bus VIP components. So it is required
   * to program this attribute appropriately when different masters in the system needs
   * to have different error response policies. 
   * From slave VIP perspective, the indices of this array corresponds to hmaster signal 
   * value. For example, if the hmaster value is 8, slave VIP uses 
   * sys_cfg.master_error_response_policy[8] as the error response policy for transfers
   * with thi hmasner value. <br>
   * In cases where hmaster value does not correspond to  master index, this feature is 
   * not supported. In such case, user is expected to keep this array size as zero, and
   * program svt_ahb_system_configuration::error_response_policy.
   * 
   */
  error_response_policy_enum master_error_response_policy[];
   
  /**
   * @groupname ahb_generic_sys_config
   * Default value is -1.<br>
   * The Default Slave is selected when the address is not within any 
   * allocated region. For non-sequential and sequential transfers, 
   * the default slave provides a two-cycle ERROR response. For busy 
   * and idle transfers, the Default Slave provides a zero-wait state 
   * OKAY response.<br>
   * Used by the AHB System monitor:
   * - Set the default slave for the AHB system monitor (-1, 0 to 15). 
   * - The AHB system monitor will not perform the data integrity check
   *   for the transactions routed to default slave port.
   * - If set as -1:
   *   - The AHB System monitor assumes that the default slave 
   *     functionality is embedded within the bus DUT. 
   *   - The AHB system monitor will not perform slave address routing check
   *   on the default slave port.
   *   .
   * - If set to a value in the range 0 to 15:
   *   - The AHB system monitor will perform slave address routing check on
   *     the default slave port.
   *   .
   * .
   * Used by the AHB bus VIP:
   * - Sets the default Slave of the AHB system (0 to 15).
   * - Always the default slave functionality is embedded within the bus VIP.
   * - The AHB bus VIP does not sample any of the slave connected to the default
   *   slave port ID.
   * .
   */
  rand int default_slave = -1;
  
  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Default Slave in the AHB System
    * - When set 1: Default Slave checks are turned on for default Slave.
    *   The default Slave may only respond to NSEQ or SEQ with an ERROR response.
    * - When not set (0), Default Slave checks are turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit default_slave_resp_check = 0;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB System level check on Decoder in the AHB System
    * - When set 1: Decoder check for hsel to be asserted will be turned on.
    * - When not set (0), Decoder check for hsel to be asserted will be turned off.
    *   This is the default setting for this parameter.
    * .
    * <b>type:</b> Static
    */
  bit decoder_hsel_assert_check = 0;
  
  /**
   * Defines multiple slave select signal feature for each of AHB Slaves present in the system<b>
   * Programming this array for each of AHB Slaves present in the system to 1, will enable multiple HSEL signal<b>
   * By default, the multiple hsel signals are disabled for AHB BUS, Slave and Monitor Models.<b>
   * <b>type:</b> Static
   */
  bit multi_hsel_enable[];
  
  /**
   * Defines the width of AHB Slave Multiple HSEL signal for specific slave.
   * By default, HSEL signal width will be 1. User can control the width of HSEL signal for specific slave 
   * by setting this configuration parameter. 
   * This will enable the user to configure different widths for multiple HSEL signals of a particular Slave.
   * <b>type:</b> Static
   */
  int multi_hsel_width[];

   /** 
    * @groupname ahb_generic_sys_config
    * - When set to -1: There is no limit on the number of rebuild 
    *   attempts on RETRY response for a given transaction. 
    * - Default value: -1
    * - When set to a value greater than -1: Defines the maximum 
    *   number of rebuild attempts on RETRY response for a given 
    *   transaction. Once the number of RETRY responses on a given 
    *   transaction reaches this value, the transaction will be aborted.
    *   - svt_ahb_transaction::status is set to svt_ahb_transaction::ABORTED
    *   - svt_ahb_transaction::response_type is set to svt_ahb_transaction::RETRY
    *   - The info of RETRY responses received on the transaction can be 
    *     retrived by calling the method on the transaction object-- 
    *     svt_ahb_transaction::get_retry_response_info()
    *   .
    * - Max value: \`SVT_AHB_MAX_REBUILD_ATTEMPTS_ON_RETRY_RESP. This is user re-definable.
    * - Valid range: -1 to \`SVT_AHB_MAX_NUM_REBUILD_ATTEMPTS_ON_RETRY_RESP
    * - Configuration type: Static 
    * - Applicable to master and slave agents in both active & passive mode
    * .
    */
  rand int max_num_rebuild_attempts_on_retry_resp = -1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that the bus grant is 
    * given to all the master connected on the bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to check that all Masters have 
    * requested for the bus at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_masters_busreq_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify which master is requesting
    * the bus and which master is getting the access of bus.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_cross_all_masters_busreq_grant_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_all_slaves_selected_enable = 1;

  /**
    * @groupname ahb_generic_sys_config 
    * Enables AHB system level coverage group to verify all the slaves have been 
    * selected at least once.
    * Note that to generate AHB system level coverage, you also need to enable AHB
    * System Monitor using member #system_monitor_enable and enable AHB System
    * level coverage using member #system_coverage_enable.
    * <b>type:</b> Static
    */
  bit system_ahb_slaves_selection_sequence_enable = 1;  
 
  /**
   * @groupname ahb_addr_map
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_slave_addr_from_global_addr(),
   * get_dest_global_addr_from_master_addr(), and get_slave_addr_range() methods
   * must be used to define the memory map for this AHB system.
   * 
   * When this feature is disabled then the set_addr_range and translate_address()
   * methods must be used to define the memory map for this AHB system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  

`ifdef QUESTA
  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_data_width;

  /**
   * This workaround was put in place because Questa could not solve the nested
   * foreach loop constraint that is in reasonable_data_width (out of memory errors).
   */
  rand int questa_log_base_2_data_width;
`endif

  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_masters” through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_masters;
  /**
   * This workaround was put in place because INCISIV is unable to resolve the 
   * hierarchical access to field “num_bus_slaves" through bus_cfg in the right
   * side of constraint.
   */
  rand int num_bus_slaves;

    /**
    * @groupname ahb_generic_sys_config
    * This variable specifies maximum address boundary limit for a burst transfer
    */
  int burst_boundary_limit = 'b1 << ONE_KB;

  /**
    * @groupname ahb_generic_sys_config
    * This variable is used for checking address boundary based on configured max_addr_boundary_limit.
    * Default value is 'b0011_1111_1111, which selects LSB 10 bits of addr ie addr[9:0] when ANDED with addr
    */
  bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr_sel_bits = 'b0011_1111_1111;
  

  /** @endcond */

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

//vcs_vip_protect
`protected
+P1+f>FQS^.bCgXga?X]<TMeI96\e43>W,&QN42Hc+ME8(af/XIR,(/[9EGJ[:2/
SGGfe9a#]RQYUOceYH>&bW,^SJI>(&KfF;G4cX6=BJ?L2:ENf5((T320\,U_HA#@
NX,fY5_cME/^6C/QfBUF<:T0V@]QNFRCBGK&V]?#W7^IV=;#>2,<A2D6d:J^5D/]
[8XTCWW18_^HE?8DX2=Qa;Ba3&3[X]UU3;ZQB9B4C+IG0EfF=D,(M^eF[CEc<.Y<
?EgH(]+\8,U.[U=4/\cUSV[4be:7/#6aZWAR6If^g^&aD[c86[^Xga03M0/KAA]6
M_1YTc]<RBIAJ^]^D^1EcZ_4g=7eC[):KW=QD9R&65ZVeH>4I;D8FL0R:Y?:>F\Y
d#71TPWH,PRg(.gb\JKCe\UNW.7^Le=NMJc&3f,&bER5ZI@+@&])G423IcH[>AKZ
[eX17.\HJ0M^:U75P7B\;b[C/]-8^MMX-Z22IdHNd)Q8G\;7\2Ae:\.X08efYge>
E,d:Y>HAL]:LDD\Q7#b/d4<2?eRN9TgAF[4)@K(\S,65.PX[]EZEZ.H?QJ;,Ac@g
f_=)]bY/8e9_W3\/5R>T>Q[@M76f)N8IJfOTY@S.e^]6U77LKCDC=J-HL\.Tc8SV
3\ENAW[(@Y[:7fEQS_WY7O)9TfZeNA]/\?>]gH-WVEeA5)CKGHM76&,)[e#A5&W-
V7W0dWK.a4^Bb_@=574Xc50G>b:V:3g&<NBTcO.=S]5)+<1R.dd8]I0Qa.J>AET?
fEZS=Z:?S2K?99[=8TQ(=QG/(EZa3CV?gA=Ng[WKDQe-L#FaSTTV?O^HONA_79C:
KBgIcfNa]AMQ:>]<GS[e#0+MYf9UVe]Dc=KEAbCW7,2?_8ZgFPd6O]?PD7/b&B,f
NM_bSM/e@UcdV-A&F#8VBQTVge@+VQ1Zf1P>\RK11_[d_KUEX)-4=)O[A[41)>O[
M0W@dL=3aWB.SQLH&Bc^ZLV+@d(BT2#c/_]U5)44^G,PEgWfQDC#d6Q#,):;;^D^
\YS8.DNXefc+_&Q\a.\J8.8VePbWFE9]@-6I]^AN7feQNDBcb-S1B:ZNMD#Q(db@
GJ4gVfG)E<4[F0#<W2KR]/R;L:+DV+JH@9T^=#)S-1VZYQ,KA4-G9=(<gZB_ZT1/
=UU[B57)(+Q4C<D,JJ27\=9Y>[d#0SKN^I(ZV<H(e2g??&XaIPZ-]S?;]LSQ[:c<
9c@?CU)_BPBLP&E+FgQbH1N_+#?\PT8S#A^R=1475X1VN&+La=-0;6A;3fBgLFXD
IaFGgaI39A(Jb@PeWJU[=Y\@,gBNb<^R-QeKJ5L[Y:e6ff[(.WXH:gYP0HePC-c=
c:K>TFK62Zc76M\Qc0<4b)D+8<eQ7(V-ES9+:ZSM]Id-,LFASP+]P/a0VVBYab;T
7YL#-4,BgH,\5.)BK78Z;&NO&df?]A8P4O3Ig#Y:@?F2>dE6g([VG+&++f=3>K2(
\._;Cg0J6]6A]:9@U7X9&7[D=e#<N9KC5GL+@1;+[@9P+D(?&P<_P:+-+SeT-?11
_T5_+cBPV1@]YG:,QffQ/>Y?S6g2@1D/=Y16c+ZK/JI0,@2d[+d23^(U639;ScIT
cgDg<Y[?@(]58H8/D.OI_>)^?ba?L1LOe(-7NAM:LGSdUQf=G+T]A/]/JF/=:R0B
?KA<.X?,E6][?SFGf?&PMTPHWX-.O+Q^HP?;cM4U&SJSN=eZ)EAN4DZZ&Y7VYAMX
VK<ARU8&8,:(+)JTbg[MQH\O7[H8GH\?f>3XaG:9<FbJ,Q@g,gN/0T7f4\(8GGN(
-OPeT/SL80<^a,<e9?(cGN;_2=-,-c,+bG0B^gUE(&=,SQO;Z^U1>@Q<>UW49UI-
A85.a0U+dFTSS0(?)P?>NZ3-\H8)e=\3c@(MZ__GA055XH8R]<@0AedWLgQQQ+Z?
/YO>[:&eD0Pc.I?5c6BbK1X9101<_KR7bJ>();)fIQSE=I;;,W>2ZIFgK](?&efO
/XfWH721(f5JI<4=14cP^,8-^g[LY#gEY@b#Z06Lfe^^cTUb_(9c_F1,HYcB9Fb1
ba1(&@>+A-S0_5[M.^ZP?fV-87\1fUN>PFG4Q4ZSA:B\EULV.NRgO>GU5.=):;_Q
1<^M5F^CMRTdK&AeYU5M#gXT&O:^^UL:?[-c7M5\7PWZ=HEKb5#MHC<dNd,@+BJ(
]W[=>7<La=a[LU]P-Gg\LCP0IGBVW5PQ[_/.d&[)bf@W-,PZF3/efWU)<\Rb[.GW
Eg4DWJZbF-aeN\^@SBXTg7K^X(2:68M25g=-H?D&&JKe.QJ9=OR:B&+f3;-U(7O>
X\9++G]U)I+;FTef_G2<LM[9.DB0LG/6e[0gN[P:FDE&-d=UaS9H-Z=OCZ_A=AUO
@O>WDB:+\HTI2.A:&fg\gI/a=J[QKELWP-7C8U)^AU-\P:AJeB_+;G#<RPe/G,]9
/HTb9^XA6e3AV)5ObUATY_X<dZg>Z[@fIWO/I6M9SfNNBf1@[.VK6>ecTfNIY9#8
@O]SgbVc+-7UO(F3U6:0?0H/[+PE02;#V[bX5<b+B_[[NJK3ec:QWNLcS_Ze(e#2
WCbf?39#444XbB)#W<59;#94fL-JZfXg+4E0[=]#:K]-c[>U0V4KgT5gYeCR2FeR
5T7=?Y=&SLZ2>,E4D3eOTL[R7(@04YRZ6ORbZ8>gT5aLeMeL^gbZ_c(NT_AfA]^Z
7e^G)X37>(51ZcLA:HD\_,0G5D5a_Y)O:62[,f1<:YT<9JQeN]bBa,98B1SWF<I#
/D^Q^DZYYK4CP>aU6T-@6&e0,<&8CJ7&2/7+6E3E55RUc\2c]&>Mg[a?;D2[f,OR
[1Ng?b:X_;NB-)?a6Y@0&-7^Pf3XbNVT-aF@,ebGS3gdH)^AC@>I7.SN(/0:WVEB
4G<3P.5L86EeRUO1AQ#PAW9J>2@DM(_M4^2=:&=VQ\(>G<cLE=VZ.8_+U;M5O:@F
EI13dP\^8G-W]C;:7M#./,?#+HG77a:-MH,A(gXC(9c3#_IZ^LMKI+NX21;J-cc<
Kgc>CV>0Sea81Ke63?/U#_?cMG[G[-(^WPRTC7@QGbS/9_;3.NNYGAN0?@SX?8L^
X?bHgeNR[S;Ib=/c<3Q[<05L@OHNaYV2gUW+>B,N[>ZGTITc3W6XRf.D3=NQ,2cT
bf.E8=PH\_&:(5[IP#8T24[5B47^87TXYH?ReHKSBb:XC_e82>2O1JMVaRE^f;V0
1;^c9P&VfRG6-cZ(^\HfE-VS_64>@FNXLPb/d;S^H7.4I^1=Y1P\OO]P(#L;3E/<
^B;QX&cNEP74AXUY<YEU[GL#GK&?)O.Jb9KI5R1?fdN>E69#\@g<0dB#>OY29V/E
KG7E^.LHPAMb=MW\<^cgA503cVMN1QJ>bWe018PBHc_XBd8Q2#6[DW+Y8-8ND-R=
6E23a6X_Kf)b0)^78K_;P(=@.fEG.1]3gTQ=M](&=:?0_D0a<>-)JY(gAb4M_27\
GYWcUC)?#U/6Y:aNX2ZG<a&5@KegYOgHba)e9K1@a<(A:6-;/;.Y2,69_KDH<NWD
-B+1Ff(/KA[a-I=EbDHJ4W#5dHZMIdI<7S.Q9AV#KT&(@)BZdI+_Z.K:G:d7e@AH
W0U5Be]>;2.c1P-//fc[HN(#MLV214RJC[BK>RaaQ=E&WU)]#W]Xeea(8W,LQ2V0
X<eKJ3/]NV9(IGN)C10FTU^QPU#Vc5G2F<cB]<XW=5c7O_036H>b@#RCN\\aQZS@
TXK(7;;d271#MZ[[58Odc(;DgXIbA,87VL9.cI[L9c5E0RWag:OPYbf^TY[+?1O9
I]X81-H,ICTIJUJa3+2I9&/2a5K>4;J0H6^RY;Xd,>/V;3YFI60SQCd_ML_6^:21
RTJeKgfO43Pe0d3Y^S(Wc\(A^]5(K8=PO>7\/1K)D(#+cIBgTFHF]^>8@TE\/UZE
J/>&aC2WPgdS>H#VW&-Je1X4]1:-KacPU?1YbRKKDZ,g9WKG/Q\7;a>f3[VE>1OW
b-E/.f#PKCGd:5921;EFP_G\DSOD.7Eg)D1c<Ve]]H_VGI0fJ>\]5BPJNK)A&0Jg
]e5HP(,\;Q0;<M\4K;Y?GP18H?V\&\f><05bK3fKM[C\1,Zg)I,P^;#?0XBG4SV@
#(0gW3gF0#IE&KMCW>:RAc3HD^\J+<Wb@Re/53038B5e?L6G>1K]<9?TER]52+_Y
VPU2O#1\JM4.R4Q><ObB8PW;\.G\CE2;J04)?2>aSSJ+6,fK4bP(&e^N:0?F6(SC
/8N_+(K]Mg(R9INBX<c9(67<L;(?MgZF8f.WMdaQ.39:B:+M9[8^\FcfGORC>E+V
CXA90K;cWb(Q0U=-R1dL[^];V@E.1=)IY,b;gdBH:F_@gXI(/\,_-EL?C346dH+:
Cc=cLW685C,8753HAV@BPLL@&5.LFNZ^)4,;O1D+J1H/LG?P3gT]\+8M-bW5_e5_
2)JB##^EOO>UOXW/9bR6,?J[4\I)JVc724OaWK9^WN.K5GI90T+5/cHYXGQEHCT<
WD;ZZC?W6E;1Y=VeS8P.B4#F9M@Pb=]NRf:e](=dWT:^DZZCcgQZV3bC&M[6:7Y[
dBZ0ETWQDUOa3>#Y+EX9H38c5-,/=#/7]Y]U1MRe8R_Ic3DN9QI.QF7_2MHI=2K6
^FCaTEZMY=?<0(Jd34.+MO7RGXUWLBXDa9)0RUK>ACA846HQ-Q/QaI+,\J=9ZXd^
>8:,O#e.3I..[^5L//YC\3bQX6Q0?>]0R(6H;0f4RO<6J3R.cMGM.UTd@VN^YLVb
27]=B5;)ZPK_dg3JTQg55[?I=ST/X-Xc,ATK]@?2C[IM#IQ=&;2#>fZOf_>EJP#5
RZAC4;[#-P6A[S,4YFOCTa(f+,g4P<U3U3c(YZ90GPb]0LK3FG&<Fb+=3JZ^&,>_
4c])SKT>c_=\TZ9&.L42g;a-\[TY9+gd])O77?:@;J#<AU1RB8:#dDXeO@#fTYTK
1V/L63d&C/>YTa?N#W&TSO,VI7>c39>Le#9SU@27(=^,44LF7Y4\d&^;fFQ2TP:S
)b3@#f-[?XX;&-EUGKA\,9g?XO^OB^XB)RF)-XK_UL:,fOJK_@FF(VZ,>Rc=&&+b
1OY_3a9TMKQA[+YWN^<#FVD1#,&a(:=Sb_\QZO#>,dSYO_82]DIC75.f?^2:\,+A
RV9Re7(BKYA]Z=[N]-LR\/#[bK:+9&CRD#&bY)#NcIdSCQXP?W(g]6M[65G9DcK0
E?.d2g=^M[WJERP&+<63E+TbCMB0=:e<AK&@L7;5P-<P=^Y>-^4g[/f6S-;5;[DY
,Wc2Q4R)YVJH(###TG_2AP9<9Y<W=(J3Qd<1c]&LX^];.4eA^>3CHQ\dS.Lc&K23
d)CII&dIJ&D.8)D=(IJI;FU>=4V:F>GSW7V&8QAMGE1Z\K#3<AbT+J3DZ#7QbXG/
bY]H9cNP:M2Qb3Q/27@ZW:IKbWE(<5V6:g]/A..NGHVdQ\3&OKg=\b;Yg1^AJKQ_
LZHH)N<c]\O.K<J9_VZ6H,JARZZWCZJK,DBSF<(Y8Y->7#S\:V@5fQK.FP@c>#&C
03+IX+K=ae\0<4[=,<[5(g?1/F5N@STCV7>X6KJ=e=[@S]L#L9\1WW]VcE=fGE([
O_:XKfe9CV)/?>MH<f##Ac/-)(f.LXS6VPZZDXRb@73UGb-FX#MBG7/_OTJ074S@
S=C(QS(8CJF7#[7)[?R#0a?<3J.EeB6[K[U.:cb;,,:[Pg]a2]/B1(=C805Zfef=
RM2c+QS;gJ;fbQg[K7GTfd.?XeWY2\MW^FgNbTL7Q;IL_X2@2Xa5PAHWUN@2_2[M
Q]SMcI?DcVK@Gf&12E\^VTObUK7GB&R=aDOcbO+Z^QLT=P/PBRS&P3,+EEe:K9&/
V.-b;T(W,7\5cB?3]C3DP/X#bc6@3O;P?[XCQVG4f1eZ]01Vfe+QF/8_8;^BRM-:
GKLR3E-L(M-SIE#Fb[B3.=Z>dPI(:OF)f,[+8<FJ55(BEZ,ESD(1S=dI_U5Cf5&+
)IMg)V12Y@f-KJ-+105g_)<,(d08gHa^5>/_YfHN;eSf3Y9]2?/SEOX+K&?2A0+H
=>CdBZ5=5=]E4g.Bd+[J30F>1X[BQ3gbDKL9c,1H2f?MO&7TCT+a.(ae45(]XKAD
4cAJU>FHgc^ebcIV^J^Y:gSPZ2a]d5<SF\5]f81d:/1KWWR1#9aD>(Y83;be5dcQ
LXb3T1.4#B2TEfY,^V^1\0=e)dG[).MEE630F)^JPC8\=_JUML4;GeE>E:8Q2CO;
b8:OfQ?YdSKE#^<.BfAO:+\R6S],Q?8Qbe>O2JBf9+U<fBdP8G5C(,YH4Tf:FTSX
?4;?K(OU&CeMYffLJb,SFYLR/^27#:&#L]1e1Y#I&?9L:5ScA9,2_-+?_X(J<>5?
2XVF<eV)0ea[4>@Uc))8Q\PK<0;eJ>T>)fNe7;ZW#<<]aS@7d8@/;F9dQgR[Ed/b
_1;Q9ZX\N^UFT3(0X1?6Ua900JG/X.&@YTcYB^?#=O>T\aMKU476Bg>2:_I]F04E
D]5LH1^__SG(9O3RC1DZgC>XF\[aYA3^92E(<W3N0?bM-[7DENb@+@,3LUDCK,\:
K;53+&?bJX9034gH(Y(TPZ)[eb:?0,:e<BHR]((H:3?Da<\)AG78dV0G?Lae0?NT
HdFY05LYe&f5AJX?ND(CX0X<fMBgcC3R]7I(G.GR9WKBg30UN8DC]]Q6+2MS9cZM
TQ)9X0fRPF,BG<XV^1W-,[Y<)-b-KC[WHG_dM@^J.\_LGaD:-gP_Z<KA\]QPQS3A
_A_GF\J]E[aI0(I&)4&]P2>aTEgD@S98^R@=KdC_bLJ?\N#Q7,47AE:QS,aMTf#G
2L,JCe=^W.UPATB939@@HWa&;O<893W?6=DfPH8,3G,Gdf6aF.+45FLCdQCg68O:
\fKAOccFCE_2&W/W^6:BWa#L33T#UEUEJJZQ30NM9SO(#d1[.?^;f>=@HUG_e)G6
d.WXRU1gO0(DY\+6T8)O>.UW:a6/?dX3>_\;CH]4A>COcU//=5E.U]JP;7GH>@42
d><B:.3[#U:+\f)c,T6#I;=QKDF7J^O&\O5Z6[;TSJ\DLPL/,7f<]_&FHaXG[dJL
SK,=c0L]E8.1-+PER,3M]>:OgOQ)A5b\GaW=T2JZKB0TI>Fc0a).FT<?I;67gL8>
0U,L[>4&+5H7^?Tb)^d13EE(g;=@&PDL^A:?ZPP=B5RKZb3<WO.+(CeWG10cSEfE
4F?0Y]Z5Y7gMN3A@575=A;\->.S0<(Z;Ib2=Y4eb02KH9;YP/Y_W)L?IASgWLC;4
<R=gP>\RZNU4c?,Uf;a1c9N+.^(Z&LZ_53#&O9baN2)<@PZO>3THc+G/Md4^YV48
9W8?))e^3&8HHa^O7f;M&NK^KA:RaELCbNW+c,(^0&AI<I>6#^8BS&c0)CRCD:1S
eH237,]Z9T]OQ.c&^&1_?_<EL^=1VcZ.6;?Hf1.WC2U<2f(SE94RK0L>2CJ]LWbR
AY84@?5CaJ&ZJGfd@A1<]b=NefHSe(D_1MUfgLJ?&KK@EHdZ1g_-S[?fT?#=TX\c
?USgedSS1^IKG9bF?,7+:EB]8.5X>#(D[X-)&PTe?e,AWf:g_<ecYQ7LaYb7+5:D
;JR^QZYFH4R#HY.\US[5g/BR#5M>7Y_^0a6B2T8KS=aTD&.e#S8;2eABT77Zd5@&
Ld8.+</YE@67b81Z)gM:,)X5de,G2][gb#BFc@[^H(3e))00dRDIP8aNA+23@\?O
E#R8HGc;1+U?7JQZ\3^>I,O;S23:NJOKb#5B>_@DJ+()[+N#7V@.^@6M;=7RP+Rf
0Rb/>bE>9(MK,C)/W,K4CJX5UW3=WPQVTZ#^aC4<YOZ[<a)_-KCg-2-3S&6IJLWI
Le-DgUE[=^QA?U0:C2E^bZB1FWgPK<;d;D@PX1,FQG-(^a9bdY=gRc-ND+f7O[4C
YGPgYET@L6Ed&SgAE]1J9Q3>\:C19&86\gaB((;#?95L[K;V\7B<5@H/[QJ1G>T#
1K7.f0ZZI:cd.d/OXe74>0VO\4&LB0;Y5(4IR[/JF1R2)aR.:\G.]>363e?ZK<b+
Z#,#Z/+8E-Z,R@#1[:]0HGb@[6X9Q[Ag+](7H>A3YM-\?50a4,Y5116>^>g4LFV7
^J]7C5gd(4H(O&7YW#1,_,>S@R0?d,&\f4FZ[&BbOaaf9)ADYK&=;,5A]#FUQ\RS
2I[X.M_DaSgI&0)^f117B?ePN5#>c()4E9WLSDFJ]9_Hg&6K>Z_Fe0F]A\&6;KO-
7F&^gZEV07A;bX=;BVQ-+MZUDX9g)^H>-Z[=?J#H&3W<(],P:&FJd3NT4[0,e6eI
cLFR\U-eg.E?6:CSZ^[3\/0#)(F0??Ja<A=L(^3QG(.:IN5fS\8UX/LA</fE+(^/
PMg4)3C&8#=UEXSJEE_bTN0MG6W)0F8@g(Q2?4B?]cA0IUW<U5[5L4X>97<G2LeT
KN=@2/8#,RG)2#F[YT@;&^f(2#Z@DNMG_;V7\NZ:1L@0XX([N<Y<g>AfMLOT-bCL
BHbQ\X&\WfX]a0C0Z5YJM)TbXU/gG7ZD&_daEg3Mf8&B?J<@#EQ(Y?H&3IO#0?8@
I&MVa:^(L7<gL[;IKE+\GgM2AE71O3@9)T\\^7UY<[:J6QZ&Q6AMgNG1c[H&<)BS
#@VKYTQBMeDPC#ga8;b<g@3C.BOJ[,5:Y52ZT-5G]:_O/EgbP.(2:e9;QVa:]/6X
3a8JI.d09I]\VV0/Y_EL(M#f4eJV\;TgKHDL->PH[7L,\NE]DI35A5[4FW@HR312
ee/B6_A_(W)U1Kf?7(?+Oe3eQ;[?T]HLC628RH^].,XEe_#-cH5+ZB=Jb^APg9[,
\[G97POUEXA[Z9U1ZD<fObQ--Z&/X>8(LW3cK3N^&>JaOgK+J,eABX,6,LTS.:L.
E6fc,X;JJ^4F\FfG./-\Q5;>S\BJ)0>3d[H_)TK,>==;^U8?/(N7J9^4f@LF_TCb
P\6;W@M,g)\ZHX0VVWcO.7f8aC]W4IS\5SFcg+,\Tg)+L2V?f>9LA2[TW5;)e&N1
4H2N(Q.SgVQ4Jb0)_)(GK-XK,EMFC))H4dC(Z>TTW3235?F6H^^]=G9MZ+M1D)^/
;\/,>E/LT]69)e\.EV6=XM;(;W67KEBPLK4>W[.)O8[TMPGE1+JFa4U\/H4<cDV]
<<JN(VXU+.NI7HJc>W]U?RLfPa)LM-I/YX_BSTgH:-5M+8U<CUQ8U.3V3Ne;_VSX
P7F&W?&O0BT_]@O/R-EXF/(Vc6-@ZaGTF:)+LV]58AAcLV99L:+IZ^RM]8=(Q+4.
\_6DJ=Z<L7V:&^NYJ4U.?S;OCU57=.Dgdd1H;=+gGR^IAZ?b,PD5-)8@[?G&_AWR
,&JIPgK_NJ(\W[f5HI=??deJJCNOZ/HU7>D9M;NUS;a2_aS+H=>0CYa2IcKWAB=T
6AdgKd8Ug4,WU0fN];S;&dK=?=83f6cGX(_>dZ_48><_]?-C\LC58+4PK.G5HIKV
+9eL^@P4_+IUZgTE)d1e:9D@PWe2b+]+LBAWe<RY-:9@>SY_F/H=a()<0SUVR1X:
+#=HaNUXO2O(6+Y^POV/OT-8e<b)IZ5QV9M\Hb]0;13N+XT=\/<I:V./RfOQ/0Z^
-E\>?;^\O/UB;KfQ+S@J@9U=gEX/G(FLe[/:N.g99f/Z>RQ:06]T^C[KI-XE=gHS
1e#)_V1H[APbSS98AZ4<;8MePZ(:=69M\UTZ1f?[TMcDbdUZ8D5ZGGUb#UNdM00(
(?gW8CB?C]]U?3dYY75A+.OT>bBA794=F+LDS?^.P5ce72D>/9d]R]GcN)1(fY9P
G7;>84,/.2bF-H+b#AFSWA,DX_d(W@dR><Gf6@dS]eWce[c/FL+>9R2Q&G@>J+6F
<0d(Be(WO.A:I3a@]JZ[+31NM<0A)-+gF[@E0KdO&f;;MAQP8NbJ(/gE1]=WW21:
@#]gEKFUeUQ#4XPEg=V+4TR]8LJObQUUBR_ESgYAFYBY(^RCL40R:KBJaESN8e]<
0PZUe5^dN?ASI4=\3;<.N]#ecPc@D-2]CY@6P.KRKZg7a5\dRS>P3ZBc5?&P4dYM
\;P)YJTVY-P-0EBL]+dI2WeQ3.12/]4NW+ST:3[B0<VFQOR01FK7=8>8>01L.a\L
@TG2_3IGWK:OV\-&#8aH+.GW(C22?;TJR.f]#(WTeNIfTA,cKcfJQcP)^)A1GV<\
a59K-R,IP-LLMOEG.?/D>:;?4dU#GW<_^Y5VAR809J:,@^OP9c8WVT&HeHg_#23X
2R6V91Q946AV(HC6B_6Kc>2EJFe([A#TaSDU0TMVFJ;f5EC(R#>UB0DBT5e/JI_]
G@S#;N7F#WF:>LcOGd>;E&;:+]\L-K/<cR0I;4MDKEa<aGT/eU\;9)&.9;@fc[2/
(RGYHVVYIEA+9a?:#=W=HCdeD\f/5TO^S1.\&87;HU9e=aKbb>#Q^R,56,7HF8MN
faeW4,aR(FKM+^=N=CD?N<e5C]-,Qc[+2UG#4g3fSeLcYXf4?F=G97V2OaEG\+2a
QPK9aL;#0XHSR2/DS7E?TUeWD&4;(4W+H,P::8;d_OH@Hb;O<g]?92QP:LfXF:aC
Wd6L#7#NHU)(]9>_D.Z&,[5.]&Mg4X;?db9S0fP6LH@(:969/fOCZ5Z/[-81@^XC
O[U&53M?).NT_L4bDXe1>DTaaU6Q7WgW[?+-46,5Sf2C=_a91DPHKAe;\eLZA/ME
K4+:3](-?E7T+\RGgH&90PM;-,Pd6CZ=J]@J5,?XSW?bXC#N(B/3PWU)]DA\<4+.
]OHVY_.+RAfP4gGVYE7a.(F))[gT1gU6?^-6de]Qa>Oa0U7d5_)YHB7PA<8X:4W;
;GdMLcHbQ_-2JT###=)72<G)QFIPU+WIHBe]2e#1Dff2\b5SB2_J\89JL[6A=VaZ
EMQGc[#9bWe)a:J+S]2<PgHD9)9::NL[0_>IDNWE;3ZK>S(c?TMW9a[[1CRa.9UC
a9P;8c6c/AR3gX]=&)1\,&E]CSG2]Z6>F6.cgC(R-+:-W6C?dC:Q=Fc@)[UHHd?L
c+RIT?2HGUU<0N)9U<IA5(U5Y@-3V(#&LO2#b5b[2>7O+;NMA@T7NfCM@G[7?@)G
Z5LOA8,@\0PYB:Gb5A>7Z?L^cNX-<](=EGJBBd>\SA@G51;Cgf(#0_T7<G;6X1OX
LZ,Z<M+<O8PE_e+=/)WUY<Kg3_-HYR6caB\R9T_/51\KLCWOfW=K)g2\+4=Lg?;C
669V0I29(fX;).aF,2.XSTJg#&XF)(@,cf_YTEG4K#MIK5ZS[NaL5XH@_(F\5JYG
QPU;T;Oe]:0C(L]H0L<BNWaDL)9/@&#,:GgUcWd?]^5Z@<8(f/[<#YE0\+3(bR-8
_>YRfab-Y06806:Sa8.YS7R@DC;2g+R&LVLcDODGJ+eN7T5_)\:COS?Z,1@Z-N[Q
WC=W&B@ISF8@@W\L^aSQSG^:2e=96[eRf1,JF,DB5H\;0)I<#:D)aKOH:JPRS)_P
5G3V@K.Nb^/EBP=]:-._e\0VYRQ=3>[JgcG4b\)Y4_)\+^A</-Q[Z]Lg_MMUO0GU
?NX[FPC3Z7?+:fNC3S,#V&2_WC;4c1HIR7(0Q1(Hg[]OZScIJ=Vd8@Uab]EYfBb6
:X@K=+U#MaR]^[S]#OCeD&^CZYLBT-H<@NTCDQTE445=Kg7e)-a-KF9=?48:B76.
N:3^EaM/:2)585G_L>FA4U,1NJaL>WR^d@B3\bEHa@IgUJC>@]/M7[VDL+=GT)U6
:+@2UOBU442@B[\NM1E_JA^.CLA(&&J=Z5YA>]J#?ffLS9?b&K9W>2c>6e_MTHZ?
S(@:g.YES:QH(L]g4>VgY,a)>K>FHHAR@DJf)IF4He&-TWKd>XS1K6ZA=OH6BV+F
J>3ENYH[B+[+Ec+#C.\Z8/LLbIeb;OBcb3-YR+4PFS=,PZQcD:-SXS3^A.X893Pd
I-.,->K#M[A>Y,@E9RQ@>f\H,+AYINc\W9/:.eIP2-H<UF6;NOIYe]?UQ?LQO>R3
7EBdCT@PgfRXB+\]g@Re^K\H5$
`endprotected
  

  //----------------------------------------------------------------------------
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_ahb_system_configuration);
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   */
   extern function new (vmm_log log = null, AHB_IF ahb_if=null);
`else
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
   extern function new (string name = "svt_ahb_system_configuration",AHB_IF ahb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following:
   * 1) Allocate master and slave configuration object arrays
   */
  extern function void pre_randomize ();

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_ahb_system_configuration)
    `svt_field_object(bus_cfg,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(system_id, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(common_clock_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(common_reset_mode, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
  `ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int(ms_scenario_gen_enable, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int(stop_after_n_scenarios, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int(stop_after_n_insts, `SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
  `endif
    `svt_field_int(num_masters, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_slaves, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int (participating_masters, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)
    `svt_field_array_int (participating_slaves, `SVT_NOCOPY|`SVT_HEX|`SVT_ALL_ON)

    `svt_field_int(use_bus, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb3, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb5, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(count_busy_only_during_hready_high, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(ahb_lite_multilayer, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(allow_slaves_with_overlapping_addr, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(disable_locked_transaction_support, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(little_endian, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(default_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(dummy_master, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(default_slave, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_enum(error_response_policy_enum, error_response_policy, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_enum(error_response_policy_enum, master_error_response_policy, `SVT_ALL_ON|`SVT_NOCOPY)
    `svt_field_int(default_slave_resp_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(decoder_hsel_assert_check, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(max_num_rebuild_attempts_on_retry_resp, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_monitor_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_masters_busreq_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_cross_all_masters_busreq_grant_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_all_slaves_selected_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_ahb_slaves_selection_sequence_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(protocol_checks_coverage_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(pass_check_cov, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(display_perf_summary_report, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_addr_ranges, `SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_int(multi_hsel_enable, `SVT_ALL_ON| `SVT_BIN|`SVT_NOCOPY)
    `svt_field_array_int(multi_hsel_width, `SVT_ALL_ON| `SVT_DEC|`SVT_NOCOPY)
  `svt_data_member_end(svt_ahb_system_configuration)

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();
  /** @endcond */

  /**
   * Assigns a system interface to this configuration.
   *
   * @param ahb_if Interface for the AHB system
   */
  extern function void set_if(AHB_IF ahb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_bus_masters = 0, int num_bus_slaves = 0);
  //----------------------------------------------------------------------------
  extern function int get_num_masters();
  //----------------------------------------------------------------------------
  extern function int get_num_slaves();

 /**
   * The method indicates if a given master's index is participating
   * based on the contents of pariticipating_masters array. 
   * @param master_index Master index. Corresponds to the index in master_cfg[] array 
   * @return Indicates if given master index is participating
   */
 extern function bit is_participating(int master_index);

 /**
   * The method indicates if a given slave's index is participating
   * based on the contents of pariticipating_slaves array. 
   * @param slave_index Slave index. Corresponds to the index in slave_cfg[] array. 
   * @return Indicates if given slave index is participating
   */
 extern function bit is_participating_slave(int slave_index);
 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  /** @endcond */

  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 

  /** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** @cond PRIVATE */
  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  //----------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** Gets the slave port corresponding to the address provided */
  extern function void get_slave_route_port(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0]
          addr, output int slave_port_id, output int range_matched, output bit is_register_addr_space, output bit is_default_slave, input bit quiet_mode = 1);
  
  /** Gets the HSEL index of slave port corresponding to the address provided */
  extern function void get_slave_hsel_idx(bit[`SVT_AHB_MAX_ADDR_WIDTH -1:0] addr, output int hsel_id, input int slv_idx);

  /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * Interconnect VIP: If the interconnect VIP needs to map an address received
    * from a master to a different address to the slave, the address translation
    * function should be provided by the user in this function. By default, the
    * interconnect VIP does not perform address translation.  
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing system level checks to a given
    * address. 
    *
    * Note that the system address map as defined in the #slave_addr_ranges is
    * based on the actual physical address, that is, the address after
    * translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AHB_MAX_ADDR_WIDTH-1:0] addr);
  /** @endcond */

  /** 
    * @groupname ahb_addr_map
    * Set the address range for a specified slave.
    *
    * @param slv_idx Slave index for which address range is to be specified.
    * Index for Nth slave is specified by (N-1), starting at 0. If a value of -1
    * is passed, it indicates that the given address range refers to the address
    * space of the registers in the interconnect. The data integrity system
    * check does not perform checks on configuration transactions which are
    * targeted to registers within the interconnect, as these transactions are
    * not targeted to external memory.
    *
    * @param start_addr Start address of the address range<b>
    *
    * @param end_addr End address of the address range<b>
    * User can configure multiple address ranges for a single Slave as below <b>
    * Example: consider following address ranges defined for 2 slaves in a system<b>
    * set_addr_range(1,32'h0200_0000,32'h0200_FFFF) - Defines the Address range (200_000-200_FFFF) for Slave 1, defined as Range 0 aligning to Slave_addr_ranges[0] <b>
    * set_addr_range(1,32'h0300_0000,32'h0300_FFFF) - Defines the Address range (300_000-300_FFFF) for Slave 1, defined as Range 1 aligning to Slave_addr_ranges[1] <b>
    * set_addr_range(2,32'h0a00_0000,32'h0a00_FFFF) - Defines the Address range (a00_000-a00_FFFF) for Slave 2, defined as Range 2 aligning to Slave_addr_ranges[2] <b>
    * set_addr_range(2,32'h0b00_0000,32'h0b00_FFFF) - Defines the Address range (b00_000-b00_FFFF) for Slave 2, defined as Range 3 aligning to Slave_addr_ranges[3] <b>
    *
    */
  extern function void set_addr_range(int slv_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] start_addr, bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] end_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the local slave address from a provided global address
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a global address into a slave
   * address.
   * 
   * If complex memory maps are not enabled, then this method utlizes the
   * get_slave_route_port() method to obtain the slave port ids associated with
   * address the supplied global address, and the supplied global address is returned
   * as the slave address.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param slave_port_ids The slave port to which the given global address is destined
   *   to. In some cases, there can be multiple such slaves. If so, all such slaves must
   *   be present in the queue.
   * @param slave_addr Output address at the slave
   * @output Returns 1 if there is a slave to which the given global address could be
   *   mapped to, else returns 0.
   */
  extern virtual function bit get_dest_slave_addr_from_global_addr(
    input  svt_mem_addr_t global_addr, 
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output int slave_port_ids[$],
    output svt_mem_addr_t slave_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns whether the supplied slave address is legal for the slave component
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to indicate whether the address received by
   * the slave is legal.
   * 
   * The default behavior of this method is to return 1.
   * 
   * @param slave_idx The index of the slave that is requesting this function
   * @param slave_addr The value of the local address at the slave
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param target_name Name of the slave component that received this address
   * @output Returns 1 if the address is legal for the indicated slave, else returns 0
   */
  extern virtual function bit is_valid_addr_at_slave(
    input int slave_idx,
    input svt_mem_addr_t slave_addr,
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string target_name = "");

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Returns a valid address range for the given slave index.
   * 
   * If complex memory maps have been enabled through the use of the
   * #enable_complex_memory_map property, then this method must be overridden
   * by an extended class.
   * 
   * If complex memory maps have not been enabled, then this method randomly selects
   * an index from the #slave_addr_ranges array that is associated with the supplied
   * slave index and returns the address range associated with that element.
   * 
   * @param master_port_id The index of the master for which an address range is required
   * @param slave_port_id The index of the slave for which an address range is required
   * @param lo_addr The lower boundary of the returned address range
   * @param hi_addr The higher boundary of the returned address range
   * @output Returns 1, if a valid range could be found for the given slave index,
   *   else returns 0
   */
  extern virtual function bit get_slave_addr_range(
    input  int master_port_id,
    input  int slave_port_id,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] lo_addr,
    output bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] hi_addr);

  // ---------------------------------------------------------------------------
  /**
   * @groupname ahb_addr_map
   * Method to determine if a supplied address is served by the default slave, or
   * if a valid slave is mapped to the address.
   * 
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to return 1 if the global address supplied
   * is handled by the default slave.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   * 
   * @param global_addr The value of the global address
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave addres.
   *     mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *       indicates a non-secure access
   *     mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates
   *       a write access.
   * @param requester_name If called to determine the destination of a transaction from
   *   a master, this field indicates the name of the master component issuing the
   *   transaction. This can potentially be used if the routing has a dependency on the
   *   master that initiates a transaction.
   * @output Returns 1 if the address is served by the default slave, else returns 0
   */
  extern virtual function int is_default_slave(
    input svt_mem_addr_t global_addr, 
    input bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input string requester_name = "");

  /** 
    * @groupname ahb_addr_map
    * Set the region range for a specified slave within the specified address range. 
    * @param slv_idx             slave Index supporting multiple HSEL signal
    * @param hsel_idx            HSEL index for the specified address range.
    * @param start_addr_hsel     Start address for the specified HSEL index
    * @param end_addr_hsel       End address for the specified HSEL index
    */
  extern function void set_hsel_addr_range(int slv_idx, bit[`SVT_AHB_MAX_HSEL_WIDTH -1:0] hsel_idx, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] start_addr_hsel, bit [`SVT_AHB_MAX_ADDR_WIDTH -1:0] end_addr_hsel);
 
`ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
    * Function set_master_common_clock_mode allows user to specify whether a master port
    * interface should use a common clock, or a port specific clock.
    *
    * @param mode If set to 1, common clock mode is selected. In this case, the
    * common clock signal passed as argument to the interface, is used as clock.
    * This mode is useful when all AHB VIP components need to work on a single
    * clock. This is the default mode of operation. If set to 0, signal hclk is
    * used as clock. This mode is useful when individual AHB VIP components work
    * on a different clock.
    *
    * @param idx This argument specifies the master & slave port index to which
    * this mode needs to be applied. The master & slave port index starts from
    * 0.
    */
  extern function void set_master_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_master_common_reset_mode allows user to specify whether a master port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components need to use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_reset_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all AHB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal hclk is
   * used as clock. This mode is useful when individual AHB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode(bit mode,int idx);
  
  /**
   * Function set_slave_common_reset_mode allows user to specify whether a slave port
   * interface should use a common reset, or a port specific reset.
   *
   * @param mode If set to 1, common reset mode is selected. In this case, the
   * common reset signal passed as argument to the interface, is used as reset.
   * This mode is useful when all AHB VIP components use a single
   * reset. This is the default mode of operation. If set to 0, signal hresetn is
   * used as reset. This mode is useful when individual AHB VIP components use
   * a different reset.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_reset_mode(bit mode,int idx);
`endif

  // ========================================================================================
  // The following method must not be called by users even if they are public
  // ========================================================================================
  extern virtual function void set_num_masters (int num_masters, int kind = -1);

  extern virtual function void set_num_slaves (int nNumSlaves, int kind = -1);


  /** @cond PRIVATE */
  /**
   * Returns the configured error response policy type for the provided master index.
   * If the index is not programmed, svt_ahb_system_configuration::error_response_policy
   * will be returned.
   * 
   * @param master_idx Home Master index to be used in the lookup
   */
  extern function error_response_policy_enum get_master_error_response_policy(int master_idx);  

`ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  /**
   * This method is used to calculate addr_sel_bits and to convert max_addr_boundary_limit enum value 
   * to interger value which will be used to check whether transfer has crossed boundary limit or not.
   */
  extern function void is_addr_1k_boundary_cross (max_addr_boundary_limit_enum max_addr_boundary_limit = ONE_KB);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_ahb_system_configuration)
  `vmm_class_factory(svt_ahb_system_configuration)
`endif  

`protected
J]eFa6NW-FXHD(\RZH_1X-_dHPC,-Ta2eF=P;)PYU/EQaJ-cW^Kc/)680,U0.4[f
^eYcTE0a@J.H_Jg-)<MFC+\H^;8U[+gXO-\6N]F16QXLH5XAL>28IT,g24Adg)-c
O5FeD=e8PESX((daEV4gP;FV&V5Ebd#^:$
`endprotected


endclass

`protected
?E5VZb6eb8&O?dL6DUS,d#.b?S(/8/C=K?F&JFR\=E^9+ARRI]+E4)3G#b#2ceY8
4cV[H9G]#UJV>L0fVJg=XH4F+0SKKfOabI_#CgJRMRX9ZW9L0DJ93@A4M1_,0P_6
98DK15/K+QZP<&>,b>#(I1T\2-))QbJBR>C(a<HT_0W;8,1<=NPdC&^UV+3>\O?Z
Yf<#8aID:]DfcE^(+IG[a^a&Vb,A4HW7^QFZK7=K^M(G/M9O_Y8J/d4G^fO:FddJ
&e7T5cQaUf=2HDTAb7;(N9M)VXO[aSRPZUVU[/.^Q.)^>\eX^[O(ZcNQ/@)fJ18Y
?La2.TJeO.)f<@)YMLNRddSIaA=eB<ALS?-NEP4V[0\2ZCWNQ:f[\fJO=SJ=f\TU
=2Ng[bJ00EOJ#,.D6I7T&A>B9=[L6feS4V.S2HJLXb)J[,?0B>f\8P:)>/C_IWI/
@P3398dSJa3OFCgeVadND_?c#KCR0G^A;[8Df=@eW<\.FL#La)\aITeO01VYQa,(
91U2a??\e#FMLOf@?ON&8VP<OT6\7C#/YgW^T[[d2XT/[bUJ3K<)cS/8M9O/.1[K
cQG[EAE.17OU.#^V97)2G&,@]9F]<<ER8@NGgY-^IR1gaCT.XbDN;.W<O:J&g8K<
feL-ORIC(I86e8E3+SUHF]T>YKQ=H7f@\)gGL3DSa\X\U.Yg9VCQ\>Ug,Z\RHR5a
Q.aS_5Rd(3^gc#ZR=Rb(=3F>:L#&YP.+F_>PDT4/(Ha04bEK._0K8(ONgRJ36=Y3
E&Odg;)B113._d>1;-(MU7/Ub/4LbfHHHM+NJ64L<dVbeg9GSbAD1@ZZ;ge[.5EK
B.QaSP#Pd[K?LHa+6H7O^4AHT_^N41K&\.NJ)U](cV4^#gU3O2?38#@cGg9:_6SRR$
`endprotected


//------------------------------------------------------------------------------------------------
`protected
dWK:/K&V-1Y0;<?X71ZI@@OEaUTUTP@ae.:X>87H2HY)T>7#=^D5.)RT.:ZGG[1-
NAA[.EX&LY:<SZBR\(4^XYC=D_PNg\HF[G7WDU5WgR<?\UQgEH@<M[I3B5?:d>CN
Y_+44KY-WeL=12/3]c5<D&9;ZKMJ4caAf,AFA;BA>@U:;9C3PgG=]J6NY+>>4(?E
=S6I[4IQSW4BaC0;>&^:C+=5/&M_P2?LMcAWM0N=1+L&)3YMd6(E.0P>9df[5KE;
=+T0Q<ef[]2ENd]#6M,DE/NV(B.@,R8=6dM7Y@3+5;Xe_fZ]#3[S]LX0U#F#P@6T
CB.88A4EDQU^GER[N[PD7SA_EB<0gacdW./_Z>-&6R3(WZD;IY3R]Kg]D2GgY.T=
H.LJTaMWg-=dCQ>a4BIXD@?/^K=6N8QLN,]-6:F.ZId3?@EgaY3-,,e3ObM=4g:S
@V#<0<gX&1>NP<00^?GMQ2.b6B=fWD@GPC]=6HgVZ324b=W>FDZNDIVfKBRA-0V;
UcT6>3e(W=G+&ZRf5GYb2):Q2&#N-1?bYQ-CUCe\]4QVZ>43QB6f,Jc(S2H?9FV@
247HD2-S+G8+*$
`endprotected


// -----------------------------------------------------------------------------
//vcs_vip_protect
`protected
8#\0M?e\(VSDWK[RA,;X_g+[RED2+[e[gF5L\e)Vg+72X(+XNb7Y)(KB7.NTF^NW
cZC?=Sa[JMA?)71O_dWSgUeE9=Q=g8;U@T(1Ib)Q]b&@N@2;&\FMaC7O1+JcQVc1
6.JWQ#.O?7]&7T+DVKDbRN69;-aTWFb^F(8_HNW7AcgG0JL@_R+^R&D/>O4S::QU
X^0bc9()(GVVHGPZGX,7SVEL?;ONS:Xc2C]3Z@(XG=5[<X2ga05C;;c/GZKI:1K[
M^JVHg+OX=Z2Y:#/1Zf/IJ+P/f9M,)YGVaEMG/;7^;Q@]cDT?V]@g?Ig0U2#_]>^
0^&J(PLCJMG^W1HQU^gd+85.e-YGeZQa/d7_-Hg)2gWeLLQRH]0Y3T-BZM=_7XH&
,GA(.@HSBJRd_#Sc7L3ag\e6RZPG:@/G@.WAB]]#feSK_7)(R5gZ;R3659c0ZMbF
W/G;d\g]<5bJJN)M4FP0W@AWI#SMSMVb3bMfV::e^TH=gD#21G^-6GH^]XeN7<P?
08;\[e(70@9Rf@M;]<0K-Y.1\5+A43N^Qb/^+:KaM]):a\EEd#>9E.(-NRgXcKGd
,C36LDDQ##\\+]I5b[@B?&e&]R@;ZQ.3bUfBQ&BKX9^DGC8<#cI3QV8L77<Z)O\3
b7(eUONf&]KbUAc3M@8XIGc3XW066JC>D;9FJJ9IaMc,JT)CJK)YVYf2R\gIeJe[
G#])HL-(,(FQBJ025.=4TJ3Jf\WMUQX/X6_G\Bc\1/6NG.6^=R3Pb?+S&MIACXg>
@]OK\G/c#fdFSZ^09cc(D2aeJGe]WO6?IFDb3D0#f1?J[DV6X1aOQ5-Se7K1dY5K
S,GRT^6d6,)b3f)5<^?a1><?+H]39QKXS/:_@=CI[>(fVaG\4VbdNGIFEB<XR>Pe
g/?@48c[[&K@U@Sa[fg8/DMT/Be5V)_@P,I:-[&gTYGE<P:]9)#Q+<Q@OQMRF-Z-
BR29AZB<KC-EL_<aZEA=QCgIOJ2VRX+Ye/67U+)B30YNGBQ8MPCU>+.3;RV)<;WE
\(:gLcD#3FYNJ91JL)/@L\cf^=LPJ+XU^2I?DBaDSb</#>F+7FUb[d4g9N)4+7D6
=YC4eM^d)J]4E7-d/=2J#EGcg_+@1/0,)5c#+<4K;RcG:XCPfS5,&K5a4:fPIFg2
.?5)J0TUHE[))CCe:[+FMJbcWN>[/DVa.9fS5^C1FVQ9Y.c=;>2P=47/bB4;KY^a
,\g7;-F<E&ZJU7T+,1PF#]a,&7fd=._Q5()5_a=#874Z0+=.[.Z+QX+,A2TAT(ZE
\EUC\LDV:5P=(+<@F_8#_4\TbT6GV\0Ye8;7.M#J+e24A0NZA28US&-K=B,C2ff<
bcL<>bHWFGB4fCeO1<>=TJ?Z+Y9TO]09=)a;+Z]e6JS-:@NE&7K5J@d?BG&OANY4
eQ3Fc:H</L)36VT7>F?c4JfE;XIS,KeCQ:?[QRIZB8]a[79ZX>HA]<A&\eR5SDf)
ZN1/#44E(+_-f@;KS6O[Pc0Z]BHXW?S2DA-b2a3R<,,:F8aVF4ScZR(R8/AQ1)^=
[QfeNYc\0bZ-Gb^4V^?D/D__YJdfPLg8MA0O>G(#2UX(dWL9YAEP66EPPA>F3>Qe
TQ;OW(BaaT@c:ICagIT<^EIPJ/]PgK,I]c;c1YXbDDbF?E03I,<7)G+T7.8cN9Gb
YY:0W=W(a#0PMKO>268#Q]:#1;/<\N0(d^KO+@1.W7&6DKV-X054?ONQELVM.B]/
cK>)MON=@5Tg&,N+-^KQ\XN+T/#ZD)SbF,bN>0K.[W+U2=LfEEC90bPS,[0JDdP,
QU8;dc/YFKXSDZ=Y_4Y.]KYKKU/\FR34aLAL^C(FN[]-.OM1\L.AafeQROCB9:+E
68A047HC6(XQ7>5=I#7&NW)Q2@,f9F4]JAWe)V8892)>b\bU;)]SAS&BIE_KFRZ)
?e#b+fD6MG?EeYd[@MR2^;N?SV,PZ7TJ7ONcRFc=<_[GQ1.,_YH-W>.d0b-)9,N?
?Z<G^e[_WL[5LYf\9E:OS8<#S8L@GGaFRd6Y:53M.1=_H]2E7fEAbgfT\aTS8>[M
34dK07FdYFVTO[ELJ1]SKQ#\-0-E6WALHMf0CffX.?+CH@RgPgZ@IgUMG-cNfR8g
&<>CDK4_9B-gAYTg/0/KAYSRY4EgaUgIK\Be1a5B591+38SK/GEH6Q[DRb^JSX3;
2]F;d+9gK:-P3BGXKC_CK#A99KYE?HdFZ90Kc-S:]MSCVO@)BA<>)cZc5#-:(ZL,
=9A6eOE0Fd/1:SU0V4UTIHM9S4N?QG(0WJ:O>GYUAc(7[aTdW8:0_OM6YG)#J\NY
8M[UP(;PH&S6F6[AQbRKWRA_D5)YIA7)WWT3I>3TX]C,J>^WAO-gc@#:VN5&^H.#
&[@2C.R9C1K)PYC)Y4SE94WRRPAUF5ZbWDH5>O-FNW-7J_JDWa)SSCQ]?f#1,YLD
V@]AB?,4G_(XUB[,Z^;--/<+@5OcfJW>)A7)V39<O8+,B)L_;Z(R)5dAB7MKH7<G
E3PaYX2^?@0T>#)O\1f1W7,cZ;cOFQY^=::-C]9_D8\QS/&afRO==1=EBPG+,5dF
K[_K\C-Q/CbUKcB9:[XC4^5ZQX>41FJ@W9O?41HGcTf<&H3/M<Z9a\G8W)W_RY3=
X)._2R2JHb[+JfN)^0TF8J(TLQ3>@Dg>=-A9U(HU#3a]#-3FNf,<1eEO;8&INI2C
<CSH+S/WK[ZcJg6J5bKDHAPS19]O4#[8?.==UEU9?8;UEF&Q:VFfaJeS94RVD&ZI
5H=_]CK30XO=9=gLf\L629([@3A9Pb=T4c8b:&8T]TH7EQ<WET57;S3[Ne45);ES
M4f;JL>^&M/?fXf;7X_#TXYZ9+TM^4@Y7b:c-BMU?0,R7)H+g:LO/YbYUOLFYc,[
Q=I^L>V@TF_6P8@R.9/)A>#IgGNfQ14V2[FJKYV-;?^?g+O6#8<6P]R3Pf<HU_\6
B3Kc5Xe[DU6:HF6TIN2YCNb\TK\1O9V+:9@(M3OL\N])+]=AD];WE8G,BcCgc510
9^1-8a\AH6IX@V/:=_K\0Y;SJ>PE]8B4TRUI8g+P:LX]McS&[:;HJQfg/00f?0SM
5(R,]Q]N]/T[AN1^H]?6F^7VMGKffX2&Z+3QaAcg\LH;^a7-.Q33H0:>7:=f@@a&
9[WDJgGQWf0_S3^WDD+#[6:8X(M[9QH;UIW<1Q[&PR1K/OXRL3acZ];Y6>4Df^T0
HRT:X3RLfgJMOQR@9f3/9GIK1Md+=c(68aWUX1S,b(##.e_f6L1[^,>MV<O/=A>d
GV-=XQIYcBY=Z.=g[5S/:PP652gXVZ#N=++A9OM^Z]W;A.P@cc)Z8V@.Y\fU1g61
[ZI[aJa5F?f2LZD,^TLH?NN^;WX:cYO06J[T.6A)Qf/;R3K]^MQTUB86#?]/]MNb
BJE&E,0B9fPeJ+PMG:X:H@JU6/?)1(M[U3>5.RK:b^A0&../c=EZe0KagGNGc?::
F_KeRc8#&T->2T^P5N;60U1HR1@L-T#+CYN-E7<5,5K^>[]ebA;I6G>7?#B0NQ2Y
O+dV)+JdI4YH[W^1ZNW[?)&]@91(P/K-_BUgb.0VC\98SI)OZOCZ/4<C)A]b6S[&
]I2CFY8OgHNO21IR&c+g>)]4]-ZPQ7<6e2[]X:Ed?S+O]]e&J+DXRRR#^UL;_RUQ
<C9\#-0?+2^Sf12RPP;HV.7,+O7P-#32XgZGPO)ZcR0P[=VEK[/DL;0D,DL-eg12
1+8T)49NR-Q]e\b;g3?;QcKf5O9cB15SNW?Q08)SJND#SB^&BZZTNd.Hc/6[#g12
C-P^3UE&cbJ(<&HW23W?9LZAHBBbT0(B2:G&BDFOQZO,HI)eaIS_^[]GGD9<L[4g
=#eUXI.Y1<Ra[SRN6_[=Fg_O.7(OeDc_3MKU)Z><,(I@CKCY/_adePb9X#/^LIK(
-.)FQ35Q]KC@)Z9P[O69]_[8[)6b+#0LFA:9O^-T(RK^J[EUbO\O2]bb<+WR98Zg
>+9[)ZgZg75,-\E,N^9.MM@\WVe+Ug^K/1>/>U7K6D3H<I,T##1Q=[R,\XT=ANeJ
/7&8Ha;V<gE&4[DefB?)@I67F0c@-)aTAL#=2P6fE<+T^P;R[;@7Xe,8V;fJSP+@
N7^a/B#&\RDO#S:g[1SK-QT(_]X6E@)WOX+^[Z2DI-Ab-=Xc:?P#<gE[DJbH]dad
TbKcU?VGF7<TNILV5M2Dd-Y^e_@HKb,;B72Q5T4CZ2[f;V&Jg1DQgZa#[.CG/W^8
.8b)R,B4LPKNgQ2W2V:-ZQXLJZK4<ObS?e(Gc=1UD7d/O6\TPR&GI,g@HVAJPb/6
O<FH=Y/;4a/7F+79TU,E)8)[#9ESE7(],ZUJ.FXHO<663fNAF2H3>+W25XN,3:@L
(a/VBMa;^1^e:?V+OXEb4,aQ0+]AOYHf=+ZK84;Y@=&-e@J=(Xb?[XYS&^<H@aJ-
\eUVY;&Z;+ROA9V_/Z7EG+2G[/fG^d?gSG6A9NGB1RE6dJ8<I=M/e19A75UgUL5D
W;]+3@/S.3gO&7F:@LS.&=7U9R[P#W,3)b8#/6GGI7QAY)eg57V@T7=J9ZC[FGH?
bPHF=/I9MdXU8GVG?8H[4=]([<I-c+Z6F.Ye1R8@aRH(0Nb?/9L@/ZXE>dLY0_=@
@Z8^#;:BeXJYgLf/28;5VB;K9AJ=V4KM\OTAJOUTDPS,gUBX,0,=PAacT>+FHd_Y
K5HRER9AT4D?=A?,?@a:TNM?[;H-#:2\6aA=V)dUHe/4_3:V=95LC9@7)QOA&P8\
c5f&NHf5EM232(6<#6)<M&5OPC(LVfZ_6FLVf(V@YEN5[X^@F#KRO6I<)dS[YPQT
:[_/Z4T3aKTE5f?F\S1S5HJ3B\CSa[=4VVQ0Id>f[G-4PY.NPJ7+U7N^.&QCP\>U
R#28&:Y_PU(JZX]RNXNV4O.ND-@G,^E46ega2M?e<?c3T5Q7^\A4#?RNbT5<H7ec
3#ZH)c=bJR(J<]=C]=IX>0J9[@5.B<42VZ.Og9A_POeF=1>9UFKNVA6c?IISRG?B
1LfD5W[Z#Wf#G:ZKWaRP?S5QU[(V1.YZIQI>Q)SNCVLM,@X&NBL:E)13H;g+1F:L
=9f<c:]M__gfA8Z4OH^8c6)7BSCMA9g5eggLZ3:M^d)DD/)@5H0Q<cS4^_f(PMaM
-CLGaKAaa#?H\ecUIZL-g[XfeVDO:T=UBTfT&EF7-3KP;286_3H^,_@S2#I:4H#0
1/JM,EF&(AE6PcDNE,RgZQ?1AS.6IIc3N9Lb5ZRTA\)NQ./d3(RMCLe_Se^cLdVQ
\bBJF1_V_#3+=7&G4eZL/WJ,AdbAf34^=c[d\5@(aZ/MMMM@e[c)W22O4\0<WaCQ
Z/L<e#aOG3X42d^=ECSTb[D+c9H32Z[,?E<^2>g&=6CMb\6.7[CgR,OO/#NV37I_
W>dZR6?/#06Z2/U\5#)[)fD0eT;:8^WQ<8PJ1OUbJ,D1c.C<e+EERBNfAPUZ+=GV
-W_VITYHLfDKZ-#\99@97C]^6Z<Wa[Ia/1BH+\1X?e0MMb@,Ff?N&P8fAfgD7<Y^
a\PSB^02afAYb)B3=HFbIZ4&P?40V@.2a.9-TV_af:JML9L^Z#98^/]:F?CO))-F
V-T5_?;ZF7gg#P,KOBN6edgePEYc<9#+:LT0.0,\U(9=&\Of(fL;0T1bHB<]UW=^
cR4H<E.=)7:PXAe\T0T<T\PX^@VBR.dB:e9F[UR68-aIHKIXE[V;U/bAWV_F#.BI
?96A<29\7L\fNVc#@?Tg+6C[A3RI?->V,NHb7gKRT;-RCYDWRH^O?-Pc_1)+/L3c
DRe?:LNWQI_3KGFA68;LMH62;/dgE.b85fKg<PUG_X5D12d(JGP/PXI>Q&PKKXQ,
E7&#C&e\^<Rfe#ADO1bQ]&&+G<I0_I5U7@YP48;R==K4MXKaW<]7]L+]]A<[G#X^
ebGIfL(#c9JPXA<\+N2)]1Lc52[>].Y::R>9+Dc+(WLAY?;;_#P.OfUA^;B-c5Q6
M^->,V/W,T,O<T.&BfPW6ND>AZe.7H:X@=NW3S9+ga8QDH<Q(,_>(FC/C_U=^:ZH
1.:/_7(e.W;MH#-0^:/.(RO1W6NbA9<MKN^S+6B^,9X<.]@Bg4AKU=ISRYO-VE[_
?4[16eEe4#\LJDXO?f/DB<9YA2R(K9[LK@8O>?\^D78V#?KW\2+L,D-/9=NO95<?
C^PA@[U@L24]eFgZ;-Q2=<f5P>dH@]aKg^-S>HPL&T>NF6d03ML@Y@A4._FROf^]
\S6V+UBA,)Ub8+>@E+F_W,JdPCR[4D7^G2/TH92dMXf3YaFSK=Z7b0S@6X@EEa><
:G#.19^QF6Q>2&0BVU/JG&2gULRecH;^X7CfLcKebd_W]?d&P9O=D/I.88^BT091
<^N31\LO/URM6_H1d9AEM(F]Hg#09VS+8>0>0V4CL5c,/^R/S:W]0:2;W/8D4OJS
a2QKJ0W\_OcZ)EO=3[KcE:_)_CL0S.9ca,2J9+=1+<@TZ^C\4J_>D)D19K+]<f7Y
)N-G;-2]@IQAS+A10^+=?(#Wc_;/J#M13/PVG.M1T1M_gIS2LEPQe934\f.MHUN/
0/F]#1#F;@N)0[K:2B#D0-=I^66L=40Ye;+gTSB\SLW<O.&8YTK)/fK^&Q\Ufff?
K#X=;5=O[A0:[B:ZBPUe>B#+=a1F1.WF&+9KE=L@^bS\d9Ufa=M;UZ->.#<B9-[2
2_F67>IJ-P:E>X/I&cNefBH7T3gbd[7P;D]<f1HLd1T#d[YdCfP8XaUUTWU_gE.a
ZB/+5_e\_(E>+Z1MF@[TQ?KbQ6Q>S8@5([(Gf61Pb_LR@;MD^faae7S7Db8[]M>#
d8V]LHPMOb8d\<?^\Z;JIWJCHXBAEV/)5cQDcX.GU8TdNR1U&U.cQR@<BPNGK>Vd
#F,PLS98OOL2C/1CKKVc4AFL?EEcGHU&&V;N4?@OXTIOe/UF?\_C^\_-G-+JCM+-
7N8B-T4-Je>,(/(#0ILLXNUb75#E?/eR?7eNC8Oe69.QcOdR<GGV8NN7)0517#3A
[+?Q4fZgRHCV[4da6:SaCDLA-H+gaTD)_?+SE[GVTeb##65S&[D[-9+:ad4F&4W/
@D:+>WVT9+T)-F97B=CMR_;;(bGU5H\S_AeIK/_#-GZg32fVR\.#8P=4@>POe7SB
56&F@M/\f3.c\V;FN/JedEd1P41??,/BST(0UI3+(G)IU]Nc321c/L,Q-.QZS99^
HM+:<S9&MO&=^dLG[;D#IEU4d80FHWMNCNe(b):MP]7D^O?c[16<7+BDC]:1UD1#
K+LQbeZ_K[6_3A3Z;[b.#-A]K)CLb7G8H7:,ga0:>].dN;3W8=gf9NRXTO&90<RW
LP-J#LM3Ea\.3<G[eSD6?@RD\D-\NK@Id2Pf@5QMO]^18+KA?-7[eO9?>,HN1<KN
+58:U\@@GFbVTF1DZU^&G=1+9#bfR)-2DfEL7d6Q;RBV49UWFT2WY/(9C8fM.RLM
I_[4g(1F=/&RO@[5=7+S;<g?CcVYMf[4)+T/^K#S#_8E\>#NL7_EJT)3-Oc0W.G[
V)0cMQR4gX;26<9EUZE9826]c5VdfI19caR^<NaO+UKF>6W<;G_HBb-]-5/1EW9B
5<R6fHMBT;QU^?8KeAKGQ,_R^6fNT#\NE=O(WM097^J\E[4LQODROeE.0C@AGF^e
/\LO;TO,.C^R;NO+/A3>LfO.g&Cee-:;5=P(:f>G+404b=W<a8IF/fb).5(W]>a\
41-X:7-W#+W2WXfcZQ(^R>&5L(SU8gFDXYMd/+(6S++-NVE.9(D)>E[FS,[P6G7I
6:-=RJTE-&LP2DHIK>e^YYH.C)c&4eX?.^4=.V^X^P,O9OBC1X).(W][QQ+FA5d.
I0?Z(WV.FE@DMNg0^fPVFE5HeV;41>QH>3LKgT,X?<Re/.RXRW?afCcH_dH==_bg
fQ][[3W\S;>L[MU\,b=a^CNM@EZe#f7-06?H;P8fcC3Ue=&CWO;S/)]&E<8eD;cC
M?CQC(6OP,,07N?4Y10]GFaL@1eW8+YYbb#UO0)eBe]fg+5^F(a/,+B30K8a-<W=
;FWb-#+#M,da7/0^UNA=MeXNMI=g7>S[^X\U-G.fKB5VP\=6\F>1&YZ^4@?Y+-HL
CHX6EEH1SXL&LM\SaD#ABC<T06Kf;-QeQ5BD?d2J5QKE9DB);[&?VDg/@X9Z?0F+
L3>6FR\<ZF#MF)W2PBFDd//X[TXBYG[NRG1;/cXPeX,Vc]:;HI/@.LaC7,D9XWSb
X/IVV1bE<\,1,W,F0FDf2a-5Y^1A9WV.]Z7P3R?#]?TNHZNX_KeP,G&T7S/9WE)R
;<He;)-R].8&fd0aZ0L8D0X\eSGb()4XZ:>OV,>PM^1,]()G&W)=<f],N1K3U0H.
L7@fBa3==Y-[0U9R60d5/J+\66L.6M0FU/^,M[IOQ1ZdNQgAc8,7K798d5-Wg?6g
+6M347TH+H=aBQAP(K12g-Z([)OO;X6DV;5+3?/PS6/fQf@BQ@X6]W3VEQFeIXgU
Q8b@R7(&gd]6cO.5S)YBN+O2ISK^YW4HE4:Z)FgD;4I?2:O0b@+f1QE,0[/B8KN1
N:EO@,cQMW^gfLWEFR(?:1=9dV5O&^;UWPCQeU-[3N_2Q#@^ZE)13HCC2_MD4X6=
=TQ#F)W/c2V^e+;?g@UQ8Q_<;?&U<S2+8Y:VO]5L5G[]?ETQddW27OX]eBMR#<E8
9J:AUM?c#Mf>B<3]Aa#QW&3+\/5A^GX(P;(J_Y7FJW3C@<VDR8ISB<4:LHe>CZA<
QM>G+V&R[eG#.fI#AA2Y5NZ6L#1a9.IC)8a08IEH-f:1KC^E,-Ug846T4Rf]1<VT
?+0eEK_X3FbaRRV<R1JK>@Wb7D./)TDS7I7S;MK0U?5P.QeN,:BMB4R0]272WeC0
&JS<a+,KdF6Cd?)3#ZeW;(DFFf9R_)c^0]CK9XU2<,3NFcK)Lg&ECJ)[M(:WC_NB
RYL6>C<A:PA.3V49BIK>XTN8,ZY(RHI]UfL-^)TV+_7=N^cTJW716-;]J@+CHW4(
F=6@D&2Q^.Y2&Y[_O82FZT].>eW#83_J#(M6<U.N,3ULMVV<&2I==6Qf&CW))N,H
V<a24X4[:+Uc1bU5>RB-+ICG@:005fJHL<:1SM/_K=ZDdVa@W4Q+,b\[gLA:)C,=
,U[YHEJGT\#FYIUd9+]SXGK+PE&.;Y](b8OKFVQ4UFUc\c=-YV-4AI40[7c.DaYe
IJA)?/A>(6A:V^)XfEU.N(+6.-#_cNf7JB;3\TEVV3.d/T[M[Q#BG0L[@-bM>ZJY
R1WNL_>[;+Rb6Z41YB#[1P+-Jg5E&&dQLD6;3EgGW/LYNf^8bVdPSQBE^[GOD^0B
;Wb/EZG##7OYbN_YgPB<PXH5Z?.df3R&8;82=-@eY4]C<5Vc)FY-OP&F&NMM=\_+
;5dOX-=M9BZ^OFMRA<(D@GCLJF[_8XDQ[TE5HIMLEe9I\>b4A0TN,@IB)ZJ+HdFO
(7JfV[_6cONbMHeS:./9A(L#H>NdATE2a2)]Q=?B3CF4A/0dTM]+<Z^ME;D#[OIE
6EWWTHC6g#7<[5>c(AA.&Q?BMg.P/R@?a-Jf?N&?B.C.ec9[-)9eYN[TU[VA_Va)
<YM7egI5WcDe1@>.I>+gDLE9d\(HW@F#Qf_[O?RF,-fR2.O,0W0:.NcB9_AUS:)=
SOZgZRd;K:<6fNH7Y:MRYPTDKI2W0>,0P@#BN=XA^CD5e7K#eNLM_V3.)E\^NEW4
]:G+MYH3-W3e/=HeCZf/LC.?V>NQ4R7bIB4I_6T[Ld)^252_8cDJF>^PdC?LaA9W
99+_?H^-XV7]HD]AJ&(FLP<e;ETKLOJ/-f\;W:E>6gM;1b\P,3EB?(aVU8JJ^Y[<
=HfY[&fJQJ9f=@C+6KPER&S&,LR.#3e<2d\HVW;SVebG\FJV)TcbUT,fc_O<(L68
A@D@SRfD3-O:C[X_H.O5c8#VOG346<Ff/?e]AQK^#+9d#_<Q:C0KIM)(WH[6^7]C
&6:4NR:9_F5bIH3DN4/;^&6CB8YW\1\:LAUKX8J:_L#gcRIcIeFc#_3&3/aQ982C
3.a+4V8.O/#d_MMd8,bR8L\>^R&1XHDW^T>7T)8acQWQ<AbDV:.(,8)g#B[13Q=-
Q8LQ?gG5KI,;Y7dR2W22+_<1Na2G<P2.Q1II#&@-0R<M^Oa0)(gQ;_P=759D/@.d
2\MIF[83]]Y-eJ:RY9>FDWP[\T-U,5?#a]TKbUO+3H<5NbFV&XG;7b]E(BaIYNFc
F[KJS6:Kaaf0DVdfTQ]Z_5;3DBZ_6QJ(ZV.K9W&939XO@J,c8ec&2M[LHZeg_<-P
,;MU-UI\d6TK1#M.=4Ae:AV70123.4XLeFSX-V<JgH#/Xf1[VX,&[TVSdH[EgQE\
VCLc_VPG<.FR6BB93<.-#fT2Fc8Q@B#KQ?MF?)8?T9VHR4TcKL&\I-RR)Faac;Wf
60cADc;&/SI+83IdgDP>PVKUfH&dGBTYGB?CVB6AbfNc8<T)\7\Y^,-e9CeHGI.5
FLed)bQD<CNT93^XK86Z18RF+MO1I,^3a>8U17IXZQ#UA+:P[X_5G-<+JH0efHf1
KE23cJ.#605;40NHTgA^a:2)fC]8OC)K9E6=TGGI+1c[DDWJ0[156;\aB65@c.7&
(F?\RLCAD(TEFG[\CLHKZE:\Q^&[b+4)4VOT36.]49c:XbU];[&B#R@\^TZc@E)Q
Z-V<d?F/8UgUeU81S1OS8Y_0.c)8Q(62c+-ZW?:)Qc9HgG>+@a6[#/8XGQIQ^XNL
6;+7g98g@?=?TDfR=&]#&C/_D?GV9C0FLW4:[?3Tg?]N)a#ARQ6]S&V?=,e(90<9
I@BA?6Q6WRK7NBc,Fed>&73eF9_U@&Rd245#=+BW#\<b2P95JSHfSRT5_1T<7ILZ
:QW[1EUYK/<UL>&]9>Hf1H453;aJ,&_)PMS65(48/f2>)GH[a9ceCRNd&Td]@5^6
WKCH1<f29D@\]_W:_YP4CG<4=V8NeBVE#AQ@@9]<Yd=bAIQ1NV/KV0-#dfOB30HW
b#_bK[Hf>&)&[EVCX6KQ+d-,gEaI939HM];HeQN.-T)4@;NN46OKOQ8=;CAeR\^X
GQBJ.D;F?.R@;.G)Z7Q2C]<aBKfeSXe8@,a343SZ&-3,B?g7/QK=MT(E:<g)[>Lg
A?1SA/WI3Z>c^=(f0E#N10F,<Te0/HNS0SaQEdXN<LVScP#fS</K2@\MMTN(/.YI
B>#C1_\(.ZG9e9fb7:ZaR?L0<8L/TMJb901W_E#N\6fAZIZ7>W_6CeNU-&ADR@N\
.(3WIf1I7=E:-;WIcTEN3>:.3WU].E_88bVWSD958+Z9X=6P=:Xb@YQI.C5E)85T
X7dYFX,6,fDZUN_;_:1#VOCIQPY)U;L3BWMF8K8g29QSOcg[K<>F]R67NB)L?W=?
PC>?T[MQ1[)1,-aEb->X6,30b2bI1NFYEM0YUL63\M([F7e.\\D1>,=.YDD\X#W)
9c.YQQ,])@_TFD.W\b,(&J8Bb1f^b>./;;[IQfF4)U;TRH;C;@;fK5H<(E](W9/?
5c]f0>D/]UEdQ4F5aVVe7)RTe&2aSF=Y^[f_&d8)QT648EAUG.49L1Q;\=c8A)4\
CN[T;g+0#<.D3\&;6/P=&_8HC@)77Gg5]&\@M_(C;UVUBX2DdWdO<[eYT38@AHN<
Q-P^&cg):X?J@TK[0[LeS[(IEJ]f_,R&U+gT@.H&4d^fRFd+?ZTg6+Q((?@Z,^-b
c>XR3SH@[bC;f/R4Jcb:5MFXA40718KRIKD+#PZ9Z&b^GC8KJ?P=9\EXa,56)=.H
&Q/P6Q:3;D/N&D80JD3F?3\8M.dAZP[Sb37=90ZCdGObX=.]R&&,TBd:BD#P1Gd0
N?PV^;/Z9;-1[a<ACV]99V\_?cTHI9.1Hg>e-J5B]LCEMLQ/QAe?3#1Y2YL;@/+H
3S,X+Leb^]H6)M+Uc#FC_EFOL&Ka+=1L5C8ZCU-N754^:P\g(B_9_cHJDV^##8DC
M+\K?fRd@?(SdJW4ME.Y_1,/&]WE\4S)c0E11KNFd=XPZ#FS&EWUWeA]+2:AHWGF
BVL?#c1@65eW;fa7b(,Rb?@>NJ?5eI_ZTH1L&^OW)A5W]=.adVV;\1_>EKEDG;6J
e;c84&a1PfgT(_3FHL5;50BP(3T67H;aW>XCW9CR&KE<3\]H#W6\S-9cJ33\(4DL
/Z?5A^Va9@6a)TU;CD@-8Q[Wde>_0?K8:bW<c:H+ADM3aG45eGR>+#A^4+G][Q]5
,f-eaX_<)c=5WX]DU?F@L88d))PeOI(]TM5#@P8BV^]PLNU3.;._g)cS[UI5#R@g
a1T7GMTaX9@DQ3#edKT(c-g8L;O08NW,>JQP4S@EDDS;:4<7.4E]CMV4@O6d8Q;/
F^,MF+63=0/E#dVCN);Q+=<eT2DCPVT3BC:L-KHALg1EK=aR;gEa-8A04WB.TYd#
?NIYff5/Q8a3E?91?QM7^ELc^3U2HEIDFg5H5\(4C3E#U&&O6\AXLSLVD;3D04ML
d]00e0Y06CP//T:-I#.03AI9e.XPNd924Z_LH//Q8UX4=&#(8(.-S(?.ATd:1@N+
1A;a6(3XX9.3D1bR,;I?0cL1Q9N(HWf.eTZ[@U8Mga&dIEfc8+XAI@[-YD0^.J(/
\Y<A:X-INT\3g;QgcK,K/AZ@D.CV40^1>)Q;XbH9-eVc3D1TI@\gCMQUUT_OMT;C
HGe_RN.^QEQJ@2_?T30R0YF?S<[YO?HZ74bQ7O2IESJEVKV<U/,e-\W1@a@c54@e
4:OY=T_GMR<]KRMM9e)6a.Ee;XP+]gJ88HO;U/C1VTWTA1JELeK6Xc)[7T_DbVFD
N78,EI/Q#,L[]/)7(Y[B<CA:,cELS,S2+g]RaeUA+Y6Q)43)/ZJ]YD/[.cUI9D(0
Kd?FGCU21_4->VS](5d8&NV73+f,TY(7UV>bO@[_3,EN\Mb3C&dRCBe.]Y@([GV7
REN+T2&[=OKTK\f8\A(/DV6bfTTFE=OaddJ0^:bNbeP5]]Fa6]GG(7CX]1Y=Ba39
47O^N[9;I95FRCL@<<ea616A<,>HP3Q9?>Yg+1_cT-)<(OF^VY0Qg0Y1:KfCc)a_
K<Y,^-g))#VXeJ/eD7D<G3(2=>MC)?^c>T\ND=dTQQKL^S@N)#/LQ-UF1;Zc<;/d
V4fV6WRd6_J:,K1=b388[2FOZ/?:1EdAgY#b1\AX1\g/6AP+2R8VBJD>M,^LbP.b
2X3E0G[fL[)9?.B>N\K[X@a8\14-#EV<?LK10ZN+ND4T0dX/A)ab[Q0(Cf.+7V2(
NLQ)LJ5aN0]7,<V+9#VRa93NO&#AON1aET^<MbgB:C<(0S/c=&V@d4KVDIA@<HZB
-JV-5;MU0^=MWETd=9b6V.V.9U&Xb7W0\(=>:PA/X:VZZ;LG4H+=&2\?WbSCSZ@a
^bEaAdNRPBXR?X3)TOc<=)U+670C8VAGL?D&T<_<+D6NJ(N+cM5,-XJ6OE>D[(D5
JRgSJAa#@6bbcgQ5^Ld5d?BWD0?79))2U(fY.9.M6>68451U83V\NJ3d-9T>PP,@
e^RT@P0RFT8A^;8=FY@DI#KLLJ5[K1bP/Rf4Ve>WNE;&KQ,1=-P&\3,D.0FROB77
ALXdKa56Xf(91Zg>=B2EG7RX=3PIN4K^8LbL-@?3bTYG@6>/A^/O,W6=K93A1.NI
[9D,2:I\;d9EEC-@.bBQK\80YAJ0[0^.[NGPdA.V#D10a)bUF>\AW&30C1#7+VFI
&5)5<86/Z39VbQB=A5RR>W9XfI)=3SMTN_TU9#+3K.dBL^VeYM8UZ<@15)ZA:>E\
YD8FP-?QgQ15VXL58C14HI-9Q)1CI>2&VA;fR>?AHH4O2?L^;S@2/K[8,7<ScY/-
I/=D>G?#a?/OfJ,Xf7.ZdcC<R/S1][2DJY:T[6@]S(_VP]0&9E=4f0-;^RN=\U/D
8W,O,:[W.L=UF<A=XV5H:_GZ@ORLeQ_LZGXD1/+<d;a2Vab2?SKYJ,F^4]eeK4C\
J?&9\#A>\NXX;e-W1^&3<)e+4:_Xd)2OP]>)aWWL[E@:Z0]==YWX(/,1>AG;S0;I
D^3]Z/Z7S=K,@&f:R]7];&@OGO_e(HI@#D/U2dQ5-^-_/N4=7\0O9WZN=5c23H;]
#]:DUY3>U1@EBVZ+e1e<P2G(MUOS8UdUf^<9b]T/XZ6LRDNPX:c&gT)gO)3HJ2gC
RXF4NY/E0]TDTSAW/8#FIb_H9]O4,GUNMT=,7@T.]:93)1bS(e4G)3HE^VO?G8(@
[IH+R6C-D9HK1;BU#.f:OU6,.JO-e=a)5JgUR)f3f7[J1<(;.M@8Z]_fA9F0)g)I
YL5D8d;O&-DTU4dKcXWPdZW;N=^[5]06=Z0L94IY-PA[,TQ8eJC&3A[cf01^:#6S
DPJ++d(eW#20GPR4=Y0N?+A?]J8>cDcT53U(XS04.K[MUXbI3J<T/_gHf>K@4E7U
:UEHS6[G613Q363XM7G0fO89H,6[Q-JYA;gHL_@:>,\SdPLVJFV3I^[d0_0JCL#[
_HJ?<[bOC/#aRK(UQ+,D<J;&a+>MB@dD+a7G]eE#8EQ0DBgZ<JT[=4Xb\746V;<B
a9^UX6d&-XgH;SZbN2;846OPJAGY#KaWZ2&Z9e]0FI]XTAUPSKG=7UgM8GQGbL\W
]QGbgP:G2b_W8QF3#B)G/5C?4NfOE(?^:JK07WZNL4GS;35#I3.4cF,a3=,86gKG
b^74VM1O69A6AG3+93L.PIU&[:Td]MCDX3IRLAMI?+Q[&PB4.-OBE)>e#ZJ=g]@Y
GO=UWKae.d#-X95,Z]/T(.^RL#01K>VGM4EaFgE^6@6aB..:+,6eMXCU6?B4,[FP
)ZSE5E?PV03SMgb\M@W_d]M-P=H8M9IRSXTILZdN,WB1F)<1OBEfd+g+?2^3Jd9b
<N6=?)e9WG.K/NZ.:4.4fB;aF4BT74gbJU?>fE\=/+6A.=-.0^I80Z3P_=XO/,)1
4)LUKgDZV4=EdYI29(f..?\X\[/F)(C_0[([RDK#.KSBNe\>@b3HX@-Y1QT-R<MH
#1<gPC6gK;gW_>]GB^HVB<-PS>bdI)VZ=33fa]e7b@e(YCBH/Vb->c+J_.?HP4cP
4Z>#bTY6SNBB#PF5/_G??/aW;\<Jg\,[UJ7O-CUd\A&;]W#/W5faAL3a+a54Z@:_
-#Pe5BFf@,^GVV4F6E+d]@_AVdV&<HL9L3,H2KegOX@OOO:Z.^L.3ZNeT&Z[M_F/
N)JYB,b2d?=?AT6b0^SUPYL.Ue\aE6L4U+[?PgR^A(cgFc,U+cS.R5&D.f+8f_Je
5@0&99<Z)-b&KHVF=90_fJE2AV5_ICX;_Q;g\RgS.cBGJ8>28VL(^OWL4R2bf.Z5
fKI1F_U<gKR<K6eSMAb=H7KTI0_S44^]9U=M@:^@#JF6dPIH\]bc1..7aL6.,1eA
I:^;M]&DK8R2S+Y]bKF:a638KPH[A?TO;2,3:QTAE7fR.#YN1K10L#60O_.RW]G#
4:.e:YAL4a?]HG\B\DT9]<T7OA\[RM^5C&;#f;YTbRUE5R,44N;gJC,=XM<@bW[B
Q1-\&[BO2U>eCO+EQOOB/=Q/0NC)A<#RKMD61AfcX:</#6eLS,4]7XQ:W]Xcg+d3
)NVFJ=^;V:82<5PIMC[RgD;DBX4Id:^-?0YVfJH+.W#AS2G;/a?U&8(+gA[Pd[/V
3cI+Te^&g7Sg:>Rb0,Z[)[L5##-d_e=5WHK8aH9=&HH8CO(bM(d]bI:R)),;,c[A
:H(e-YeRD3:-K@_d/bWL6M_E@,W??_-Eb;Da;_Q)SYBg/#6a;?73@MXfSX_IX&7Y
NK?O#Xa^HXDZUG#S:I=WC3/Y=--/1R</@E>d8b_0V#)^O)Hb3M066d1^>6IJ)=d[
9<MME+7J75[Z\f^L&)UER/d,+2,?]@V)V5@20M@bY:?,M6:>c;9)BFgd^d\X_Fb2
9(d[H@3]YX4O)<&>a4K_,JS6EaOH^FeY1;a_AXA#O;<OV?+,7CYf0#S2&.E?Fa9^
H&\a_8)f=aY#F3X@,fQIA]\\7ZSGL8T^fdf4BOB=FT)(^@,-FF.d2>,>9;Zc;,c<
Ke3VPbF>>6e_MMNR:)L/0?F.1Q0&:+;a_e=KZDH2O&;f<dBA-YCaPgA8F&Y[10FC
2I6]ZbCLfNDMW]F_,GGMd84@W@L)XZN3-R9e.@XP7VN8E&);U5VHQ?AW4&4AZdW5
b&7QQX>0134c]baV>#:)1.TeCGOI)3K9]]TD1cTI6H8+_,)PP;^[4W^ITG^)fC>?
.5).+])Q)FG6P@cM[X^;d1;7DIU@\Y?c2\BfGZ&0eN3KYR4FN-Fb.>KVYc/2BH&X
V=0F.Ld?[d&AME/Q2V9DH/gfO:F4[GN53TRJN?_J8GT^]3BXBG-EOBb+S[12U8O7
-A2g;,CJa=Yg,CaF#W[5=>YR2ZI2Pg==XBXg>TD87T7J-1e^T.<,X7IQP,eWB.LN
;L6B4A8+,0_Ud99M-^3BH:d&1.1B<CFBWUC_TR[\26fL.W&O2JgU\O9C]09,DZ9F
gef:1NWdF?^:8N;43;&](+V]EZMQA,;?J.d;/>(f+A3+(HJ,#dYW)/^17ebJF<8V
>ZR7O]-JH7VH2Y&JCR47AG6<BA)VeR)^,5?Q5)<.6MLHW-7=+[/4TD>\BP2/TZ@J
PAX>.B>SLZ4QM6]V0U6/>X0M6EG@b8VY0dfR-+#(b9e_L//dc>B(Y^VLIc0((2VG
<JJOcdLC&APcH3.La9;a;,/0<fe0Jb+AE=2=Q>]_T^LYXT^/I,-S\9,594gGbXA:
NHCe,D@BX+ebN?#ETb,JeVN^&S:U=ZO8\fQO94D5D93QBDK1GSNH7@S)#&ec-F.N
LF#:<U\QXTOg?^e.Me96OV;5B/9&Tf4D\/^Z8NY966)g+9>J&cD5UJGZJd)6@O3F
71YKIDGX]262C8>Ie9=BO(7JN;:[XY?bFF#<VQSCEQ?5eZAZMWd6b,Y<E^&d60.F
b=f[LHM/@0=3d>KP4cDCIM163GJc&72\ce](EW];N:_=218gB^2&I.:f7I^Og#==
Q^HeCB<]DA(Af-8SQVOB-:.A+^+PZM@9UNA@7^;_3eQ_W]LM9&cK)<@M3b@fS.fQ
;<4@\Q>9KTfR=8.>aMfN0E_1PV1bVa7+OCQ..-4dJ7K?6)MN<0.7JOf;4d0-SQIV
8KYO#eY6]&R5/\2E21D+aJJLda.e\<ee+XAYdIN<V[\/P:@4#D/eL^9LaL7Z9RH\
fZ7=BU+&S:OOTAeDU28Id,5<WOW8Ma]3E9);BeZA7/0UeQUK7Dg&VAP3c@+0EU&&
\U#1>QaKHE[cMWbGIBGXTXEb_\SJ?BV,_QF>F1<Q@CIPgBC[Ud8gJUd4R\\J@NCV
AGAW^aLX3PPVO/.c,]BgS(PH:4UTU.[)TNU.EC=c_/1c1VFM4Rd6)>Q\<P=?4XN9
ggN_76EPJP)e9\<ABS@g)@HM8&VL;=4_fVPQK\NJLJP-+J#87<1cVDD_3TD:J\8]
Ba(CHcOB]]BfK9IcCW7W>4QZIV([.(3RF-DCA,^W#]RWCAS^=V5D+2&cMU0Lg5<X
?1<3=0N^,GMP.aYO+O5@gJ_Hg09JRd3K24]1d70g9Hg/3C2?JW:;[G)RBd<AA+==
F7V(+LN2cd2(Q/C5Tf7ORBae]a_YG6+S#_R7#F-BB(4AQf.-PU#2WC;g_1-F.HTU
Y[M+G=Ae[WWOU<Z?VIY=NYFVP-(QV)I?KRSB^=ZW6RE2J]@:X5LLdG@7NE9c:-AD
YD1TC&489b??EYYQBabEJQ=.?;I^@IFA?35F1YTa^#OI\<TKI(V#RQ][>:;I84[J
^O1CXM>9O_MJ<#[?HgL-;21A[WQ+:GO0QQ]V)]9NN?E&G]3&Mf0-A^@;K1c=cK]b
I8PI-<+f<TdCIWeU4-MRGU5U5LP.M_3R,;NFMWPCHg7]\UO4H9H&A<d<Yda>6N5a
;&bT0=(CNDP-8K#N2a.-\FRffG<28QRR0NJYT1.eNMG/+a-O3)PJ.B)>:&D+)N2@
Pf0f^/?&,T3c.#N)+<#Y:^Y8@@WU^&gF@3Y3PL7aP\W@)ZROW2S.Mc\?JS5Q?9;5
,\?d.;Bd=Tef8LE#AR1R3f9(U8e<?FVFf>PH<>\@afW#?b-g087Z]AT/<aC_cMCS
\JEF9#7QR).+O?+Y1bg#EP_.7>BT0F5dScFO?P(=S9X[aNYL,3@#Ng_JDU?L,#b1
,KP<cca5(bID_OH?g>DN7(ZEQVS@H);S.#<aAVbF.2K.U:RDQN?FU]f_e=JB[Q2?
QgB__gPT528<#;(?@,P9B0>WBd(WZCeP.L:;FeG08;2g?VG[3V@7W?4Ge(&EIBQ8
04,H8-E)8.LRa.0DIX><<E#T<&bZ)dL^HICUf#2(/EF^;B5VVV#b)4.A+VUXUGcd
GD(<:,R)2)QWKcZ)+;?#DaON8bT[e.?N5(TB@8I#^K[-:_d)/YaSMC-K(:Q.He3@
4X8A8DC@6.ggLB=bN#5[Q&W#30-F-WXUYWa/EQ;ec(3;M,2LRE>?<IafSFcXQL6B
eKe?Z=OQ=f\9>Hbc5^eg&W45(/K/<(b\>..a(&d=8>J(TD]F?=dYPE>bMM@:cM?G
M_d]@C6Q:JWYNaVWfg)04<9RW/a6;BU0Z.G8L8V#QTUW@aK6BQ;fK9\U./F/+1^]
_YPKgKA,X]QC\?XJb:\:(04D>PZZ_5)c-31,GI=8gMNCP2&D<2&)@]Z=DH#Q(#^N
4_dG6GR@GDd>UC:YTTAF=c:&+3:EYOPc(_-C[WVWE9Mf#2c[#XW1I;K]c&_3e]Zb
H3C^+\21(A+?EK=e9bJc@-S\G)2>HKea\E1Ab=PLP;)\#)1M\1BTNMMNKHJYLS9Q
e?_OP&^VHO^#VYOX(0K6dQGI([Re^;g.44E2FbD)DK]A0>DK@SIIGCe,?Y9FJ.:1
G,6V?^O83^I^/[J:<Yg^=@Jc<A17/4UcMN(K]0>1OLIL\;8U(bDJUYBR;+;OY]]H
fJIV)B)DFM-5F/,)b#g#QaYQ]:1^3C:YF?J;?Z;3JH811E#)&73QICCX/UH]+/M1
e-)68g1P-eDND12J<><WSGHa3=NOW+,H=#=+&9HbG7R1?OX3@Ma3d647dX(_baG.
ECOc=A-(H.)d6BI8FR#28M_+3B9VT)eGBDB]Ha(A]fRMV#)O6DYA\2^GS4]F<96f
[AN6=X7&)TH)>;47KD_^&(H=/HCFTDSS8c]KXEZ4CRPYX\:DePaa<T0&[04g=2a&
6^S4\F2f4-R<cH;EdfPaIdLaE+dAMA/X,:9QW-LNW3Q81ERebb)W=9CdV6FKXITb
2Ec>/[a-1&\e2:>;06fWCB#9P86,R]?N#J.:8\D(][ZaZ4KWdL.0V8[C?F/W4\XO
b-]R>2=[,.<QLAbS6(/O3BG1O:gIJJXDU+5V,@@4@a/@AN3(d/&9+fOU:6-;AKW.
R+TMS1_L5:Sa]&g5MAg0Sd&_X;;O:,IcKCdB56R<Ce[;5(I6e5Wda\NGf:ZJEP18
31WYG^@4L\0Zf=NX[Na9JT8dUY+H/[R)PZ&CB>RU9O=6[7=T14,Ig-H<UYTMbb&Y
e9/697+e0b/<a.V#+NO>H_Ue,_bOb;5=>a=HQ,?C&+HWB#<>CfD@.)K]E^RDA=)@
aW=CXGKCG4V,aW:D>-ee13<8<P<,YT30GANV5&Ag)29:@E()45e.H-AgN)_@XD>)
D3gcUG-AWWK)?U]MdeHH2K.5[7a:8;a>+,5.Q5Y_A1&RCRb;=4(K?_6+(<f?,TF,
UWTB6PRIS@B_]ZI^?gRf<;0SUI_8FE4eL05F=[LBL9\c7Q?f0=X^MA/bXI4M>&>)
A)8Dfg\:#7P;e?9@c>LDPA@[_UO/BUEZQ(-5PW9N,TV&5FG24]4e3EAH,E5V5E)+
Ya4B=I^R7&-EHKX_#RGcYadPScR6GQcCICC#Ue)S-<GGbV:O7L7_8KG<&0[B9CK+
.908:KO/3_/Hc[7ZcF=:3==4=,2S5NdS<40+6@^5W&YH+XBBFXH.f<:I3/AR2(-/
W?W0P_3WO0CH<W_K3(]-Df(6\P7f[J6;;e/^[]N0X-4,:?+R-Nc=1&]B583ZCLc3
BQ+9+C]-U==Q@VBD)]1K\6@<L.,FXRaZ^1#FfJJ2#Q[P>^AJ&TZI5[QI6+L.O&<#
c<d[-g-c+f_3:X\F:F?+/E\MS00U0H-@JSaN9W#0e78I-)SQ3#=MNPc@9?ELE_^H
-\4U=?g?FW(\1M+IZY3:..]3eQ@c=_?e0E1Y3B6efM.#JS>+F+2]=c#E8_C3598K
B#Y.4[9@_BfF804ZaV6G2AT_\0\@.]?>eRFIN1#HgHF6(b(E,O[E7#\NcW(D_G_U
:c^CeTP8QBd>UD2c<CV>(<QMf@)18Da=a/\AHU3HOg3b8?C15/f-5J7\(gOZC\F2
-5.HXT8_PC@,.2;c/6;2>=d?c8CNWV[=Aaf=/^IICMU.E)G1=[=/Y<&YL6AdOEgS
W:IdCJ8&6L0N73LZ=R.^1]@b+Q6Wc3>K;TRa[b@ga5+5_S_ScRZ-&A\7Q78;,e[(
8S=B1TcKA,&2BH(E5]f4&a+\#:6f/A.]HTc=@G_9@EaJY>,<5:5[dB_LDNQdbDBD
HgG\PX+69FNe?3-A5f0X&CR<01(6Q^C/d8>NLPY;2,5]@6U>dX2W>6&HNC##P.G]
b^<e29M8&0gSbY=U-9Q/>5RbQ<>O96_bZ#e(SQ:.C8_feT=8Y]=ae#<;GNdT/Y=?
OHX?ZNP4ES@Vb#g2\=DFN0]+ASG.c=NKT;?d:Z/9EU@:@3,R8ZOW)A8Q4,VC@NF&
+K)H2\8[aW,\/aH1H4<]N[)#GV&SH:?eZZDJD:b-N3S2PT52d&gd#ZN^T\ZQ+Q[f
/QV\YY:55@a3SD,5@].W8fKZ192SC[^-WZ^=(L<6U/>gDZNI,Y2WC)e4:S0:UbN5
,[5K7F#TH)Y]4K4Q=-&NA<5\4RJQDE[#X(Ld^/R/T^1:].4,KaU;H;aAe8bLa7X,
;/-#.dSFNfCN[9gg#0WS]B0=SAB\=X-YW&gT/3f(2b?0SKQaUb4+EdTU2T2=M(6)
GWR&E#SDfaEGXRT#[0V#B8<VfAU=dB]X/Xa3a<6#FIB0CFQR-1)Y6XXRDPcWFQWa
1CIFa.Ha]\aN>]CF+ON)SJ0TZ(^A&gP3]S+-<A)Sb;OBWU[cAM(^HD6T)D?>@\;.
J-S+4,aN@cVG>7b+Cg5U](dA]F5#7G_U\;]6UUQL@>@H,=;POF6?O/GBSHCX>1eD
UYC]+HWM-D1RP/7MZfXQ3(Af#.G<2KR]Z#5MAWY^6d@Lc80B#U;ER),=MKC[GX>d
\28fM>//7<=D=J:.DFQ/a37P+J3D6S<CT).-=,+TB3@(E60HXf@QA&CAFCD,T074
TITa^W>gD\53<28TB5-:_:@SW;_)KSL<5T&L\UM&U\U>>18W.gS;#]O5F]NIDMCB
Ne6GSeES(7JWWc/Ye0RA(WaCc=#JE&e6fE_\23Q9&,L,9LJF@XISR<2a^HE#YH@A
fRKD>N_E(3a.HBOGVXY7XR-.8XfRTM7g^HVAc#a]673;Jd)fe@]NIdPO((fX&;f<
W[HGZ5D9EO)AKa=CgVT/=<S8Qa8gYfFX\W)d,&;U0S_8cYAeA+A_(<91CU7Z/31[
LJXGcD5)-4/&O([B]BZ\4RNdE3d:Q<E35@DHHRbOE^JOW1.P<4\ADD@&6DI2c1^;
7d6B11IQc:BLO1FV<@?Jd;\\Na7NaV+Z8gGSc\AP=1LQWVLIQ_NZ#Y?1RAY/C+4X
fH,EdH?TR;<3U0?6RW60ZcB7(;g(OaX^DeI#GY0Q)T7>7I)QI#5S8:XD=@6I=aT\
@7/F<9KKc)7fYKZCP(Q>ZBC]YNcTV1_2@,QN4cYDE1<HNKGJ/H]G3]@IN6J)JM^\
]LXZ@#PX5K=S[e7A#)XS<1P/;NIWVPT?d5[NP&F(][0:+;OYRJ^dWET@2@\cN;Xd
[@T]E:O\gHXIML_U7RHX2XD]bE>;,IXb)OE2P\L4^g5He/0:?;6K59:<98@>2M8/
Rg13/7CJDSQ_2D1C^,N\PVCDL_@CX]CFCIg=?,:R?XRTS1S\05afKY1V.>c8N:KP
;AGLCbMf[BG?bOIg4)]_9IU?bN:8KGH?A;=<+8/DR=JTG1RK)<_9X6Qe?0G3>AgQ
;(TY;6M;.@848EA26XGB]>LZW\=Qd&&g_4O5f]69>68LC5D?W,[-,():0D1(E2cJ
TCY3d>Q#P0_+E90._59bd35:=Z?4T2f964AL7cD(^\;eTNW7<DaD3;HaSSZUTfN7
?H[9JF5Bg>:)M/4D(6C\Fc1SN<T?@_&gZ722PT6.[0.QOf(FH?BRJ#bDXW\79^++
QBdPR+LgZQMR@g>RbD)31&cUDRfXBN4RRL2W?)J>^4\ddPad2V<HS/b-O<#WPMZQ
&7?[WRL=aB^9@/>5HeS),Z^LBQ3/@KRe#6#:BD#ZgM7)P]I>@gNHL(]^<C5:1c&T
e4FId,+ZNgXY(ZNFPc3DR>-1M^ZI^XM00R#93\L<JC(E3#P9KMK#GY,)_^(H)R;@
\P_-]I8Ub26RDBGd0?;3^R2>Ug8=7=^6037+RPN/9,g^GBgNT6(SXJ.P/2NLd(;d
403N@M#+aCBVOgN/Y/14TMFGIH0A.7CM^BZG1M^O7:[3HLEVJRC8bagR?BOW\T@3
M&cT_P:bWO.bLgeIIVRHBK#2,.dC<eXY:,?4ZNbL>a@>[Y110KNAC4d^c#=8\0c>
&Q;0)ZMXR]>@8N]FH3YJ2?5Q(\M)&0aVQ<d;Mgf=[L3/GU+dD,aZgLeO60N=,Q+E
9)Z>8WPCYXB+bW_fNf7Y.Y@3T.A1U=)+O0=@NYVJ#?GQ9+,X)\K6LME/7?OZ.,&a
L8G@bOVbJY)(,5_?9BQBf0?Y578Q^#)E3,0RC#W/@<&2Ve,Y0<TG\;Sac?,f0K7Z
#INbR8<QXX>Z:5P18&<Z1;\ODdCaT1&N9KM+-K#@.@\5N&958^N./,&EF?e=V1RE
KDg_6@[TKcb)ASf8b(KJD52.GJ,T6SMHc;c>0<WQD2W]GA_b^^T1PC&[f;F6T_Gg
;<:08E@bIP,bEUbe1<bWFOK7NX/e_aN3KEH#5a?LMZ8PJW(^=.dQT@5F)ABgSK4J
QaJUI-0[Nd76F&]]SYdb^L=c/M4gH60VMDO3LQBLfa[/+QAAVUS8Q<6#d\Z/I.K5
(MU_5(NS.T<:e@#g@ef=U]W1PeO60?I/;gCA,-OI-O/e-/:?/NDIDXLR2)Y>0&.L
@8/V-WfOUXO:_5#aN6G/27.9-eJ2(KQBKf]QcHc3bH33(e()NOVH9[<WMPJ[]JJR
]Q[&HK,QXO6ZX3_1;_UV&F0dWTYJ13d]0@bC65(M]8e<^HW6&,08Se5<1,74LIPU
J;07MT,F0R@1LHVfb1>Q9DMWIC[Y\11FG4ege(aLWFD=T?(1=HbgEDNNU0:\,H&8
e63OD.>4:TN),=H-0B-C_C\8,I91^UWYXZ=:8\3W0Fc]T:#P=DT)?Y\G+J<?GBRS
b_Y<5LbS,=DKU21>C?/6dbVGS1N=b+^e#7?WR/T3TG4#5&P4G:)DYP4&+T-FIH@Y
3YM[BV>NMfI6QUDWeFa1_CMT]UO\b.PUO;ZOB2-@>KX=)7-DW6(=:9;1O:NM1_Af
,,T/0ZQHOcaHJ4G5B2#:5Ic6fTF>W#9:aaE<0ZO;g/<X9V_&=WbREDZ:YE4QQCZ6
bL9JB9Y#+^,FKJ_XJO\e,Tg(7,(-KcFHS^PT><+&OHRH<G34#+K>Z9ff7V8YaT3G
GdR&0BMPeN6:ICA^GIU^5R8LfbK(:\)C_]HDVH/S_QY?^LE+374G)Z5#WE.L)E,?
#6CHf4<#EH\TMMOQR:eC;+D#<\AeWC89b>5WR\>O9W8A=?U5LT-J7.^EYJfA/]9O
YZ]/J:U8/+^W07d0<F1K1>0Y<:U[?OQ+_9Q3-KX,DNfZXI#QRIg:BX.@TGCO#BeU
PMe0E>e.F?U,X99P#E&LF=cEW-=:#FQc5JB>#Of]#6K,O&56;aTe/+J05f6(+9]Y
XdY\[,IC6UBZYHd;G#<<M.IXVPCeE:0Ka7Ja@\WH(U7,g_LCe6EG[YU5T>IYG-A#
7[9#fd68=3BAE]9KB5g0T=#HO05Jb_,LWN+07507S_;g?F/eaOOQ<dDDV0]ES/Q(
A+3_TJ[>>?6[cDK+(QQW,b;+?Hb>S3Z9\NCdQ_QJ,K0U[Z>Ug0;Z]OZ1R_,fZEV=
UK/V<_Z@8UD2g(<])@1K[2<?+EUOV8G6&K12JA_c[e8;(]ddCNCTXC,(Se7e>,CH
2ffZgacR4_I7c?H0J]W&;@g7EDe]O>MCG_+U,2N\g9TM+a>&L)Y/D8A\5CG/ZT5G
\>/:A<YS9M4OX7Z-e(&g[)\PPg9US_9fJOb^;U\RG0#U-Ja#a;<((fEMJNVL4EK7
SY/X_L:a+E3#</D@0,<<S.gIM8.#[6LbL>e[279T=6,ZG-_9W2Ef&A-S@\>Q&S?(
.H3[A.NI2?)MbS>FeAbCQ]&M>,16-LbGDX+_D/2D89Cf-55T::F?(FBGdeWONb;M
>#>2Mc-M<2B=_d8M/RdB<ce20;TH2Ed^2&\((bT./9g:O6YT:.Gb[5d#-R-GND=9
A\@E1U>:,45,#8/&::\Qb#,-[de_J89_G-EM;:O85#@>&Bc.&FT=\MC5@F90.]TI
#0]7HS=;R3dR^8\?<)GSVYM_#/\XXR2)T5Gc2?EE\4;^AO8K\72RVEWUN0P;^Z^7
0L+XA:M7\NM:.I4R.Z-MZ_(Rf>_\]WcfB.]A[/I^6MYP-KGPPg71QWH)WcNE1F3U
c<QBI,E19Q]]dg1=A.DM3)G6RR1\/S07HU)J,Q\0(?\bgYKI\?EPIPc,>@\>G]JY
YT6^4L=(MET-)Dg@87G;W3dW;^]Kb2ZCZ=6J@e5[S\MKeOC&\g;Na,H6dGD6UFDO
L,[:&RX,DO42)CC.(E(]R_/&X?,(9<LBM:#TKeHO5CX50+8S@G\+N@UgI[N[H]#.
&9PGBN/Z(Kb9RAAV#Sc;AG]EaI=LBaG:Lc;1S=,.K0I\F)E>G>SdMZP=d8X>0H0d
QC4<_]>)GBQ[PbRdW?d6O3_&J^;3,IX4+@^YH8M:OA-WQ29b4c7^9.-)VL?g,7VN
9)A^Wb3K5NL38e<J2W791CY5+OIPL6D0TT)\MT?HB<41R.?))YZ]:3)f48d61HdJ
/XRCTa#^aF#L2&:M:+(N).OANLgf?T_YIV@.)XV#FM;37cD9=&\<]#=YUP(L)9cA
_g7+C@1(+UI;42=X,3Hbe^Q9=\7?XPEfbQeb1>F@+]3fM;[3H@,U5;JeI=9,7PI5
+O75V=cIKe1dRN4C/9=F;f];=M<&/#W#T4ZY&0T3CYcZ_39O&PZaF_MCD\RZ+W2[
6@?T8[Sd3cES:4.?I?JGa3VN++3-JQT(Z]aK,U].[I_b_/8#Je]#dN3@UcgQR2(\
b0JJR72f3R9f/1VKa_Hf5<,5W?8g7bE/#/A50<&Q_LJ@Y7J+=TJa5fK1aBcJ5D>,
G;d\M9-W=Z+E[:@1I=J,3+)]EdLX22?#54_MNcUZ=Q9);\BUN0eg(/[^U_O>@##N
V9H91)@UEX?27YfeZ&=_ZOET;Ta63+Q:KCeCa:aPA<QH.G:H>c\.<O(eF@JS7R#2
4[]TW.dHM1e,NOZbODCg]W,K<FJ13-@bR@O(aVAQ(1(\6[JZI=]N^PF>I1eQNX<)
ZXL;OA7V?0+@AO.2+A[aJ:<8e_MTJ<8]Ne]YgH#L\WcNM-1gYJPQR_^RN5(GbNE-
K10NfLJIT6_5UHMQU)P_-JK\b>R.@&K\DbJ6eW_FZ>GS:\WH-EU_I[0C[BAVOHM7
M9,,;K1&>CG_B43GAe6N>#ggIS>AWg/<;NFTXSF9:W=0VR.?M18.(H^ZU^N)d.Q@
b#+0U[4O_.OU9b6&;2;C=eBfH&=0RRBG2\cK9[C+RO]O?dK/:WUL+HQ\?agZ&U(V
NF4YF)^eWV&d=Q6&E8];]U.e(5+_6C6aS/X)>;BdAGZFeZC,(]TO\#RR3XQFe@[#
?INTe4g8f57eB1f_f]\:\M:]MN5EF4,S2aG^RIZPI#c>W2eZJb)TO51,dRP3=f(6
H\UeTETP7RLaU+@I5[D\,SA@P-MV5#cEaH^TVcYY+GbQP]1[0^:&[[?A2WLK-6bE
)#gA</)b7BC&#bW:;(D0cSfK2,D;ETQSM,(e(+Rc<V_U26gc\2=33)U4:\P(Z[7^
b_Z(<efXG/)eNQF^SVE8(SR#@b0WK(BZ5e\GP.E3&88?DWC3[A8W<RMRGWHOR;XG
((NOgM6dJG&--^@7QS;BJLU_+^RNFE^,9BUX\U0RDW?S=Of0JcYaUe_MF-fEQ9RB
GaaOX5E^84<NZJ8AINRM6:<]A54Pb_O57L->X^V-LLJ#Y>cI[(#0EEE(6_Y+;8(&
;6^\IMKbI&-]6E@<CdK5GG?BaQ3Sb,.1SZe,68JM3\IgQa5LW=UR#gB_6.HM;O[,
[c(75S-Ba@)JY6,J#],0L>C(YV(FUBT_&g.)KP::_UYOad)[FN4D;)G,,PE(LII)
#B^;?5aO8H?]57\bRTfAH9]]F^cb7-S/E@)Q8;C##+4[DAI4L\G+7dS.PN\N(XSO
8AW(,JAR9U\.MQKF^5ag(\If5,9Ec<a,29^(dXeNS_Og@8fKe@2]d/QXWSW/ABX,
UJ.34_I0<0e&f5@OTefE[)58e_eRe-?>T0CWNX&W6X5Zc.#OG=K7-VE),+[[[U=Q
a<0CN&T,F^9N^ZdWPJP:OH2??C\+=/BZ#)^(@KNH=LK&O3NT243F7AHNZC\0H.A4
8gZ.fAS5Q5-0b,;gO7YQP+((?29>)JT[a(68VDGN><BKTWDC1Xc+]&GWK_5BGTcT
;VVO+XY[4GA[G#X;Ie)QGRVH+:YL^A#BI(aWU3OKX-;OMY#^0bQ9;IULcX4WYe7K
S05/[<=ZcAa/O@Ha=<5+=E,N\#GgNOe<K8-#H@N@15NXKOVSg<9[R19^6(9UfWP(
6/?b_LK50NDN-O9Q;b=HBQ9&JA^bTOC/K>2:R^2C#4b]OfOa]BA;V9FF;-_L7.dZ
cSWX3+Y&d:(??^,]-?LGERa<VM?P@eT]#G@TGHU_V(MfGL._gc[:/\J]gK:ZH(-S
eKF>e+]7GM]X=E>GW.+4#2+fUJ[a62T,Z/7=&7.TN,8T-fW0-8N(:ETJ0O7[LQ&5
K2#86,?A7O@J<D#YSFR.HaZ_;7[e\A@H8YWKE2,C]QWc9N6?6M<-RTSC[S.I9^YG
:P8-)#MRX^f4/JdZS8D:Q[80X9C,48ba75\WJ8QQ#Z;8Da8K2MUEWeC2..GI0D@6
[1+Cgb_IT.@aWR_(O.gB7@:>[cZUdeGX1FSU6gT70Mbg0N\?bEFU?7?PQ0VE@cK-
8W8aHPD.c3]VO7L,dQ^CNXD.Iaa4ad99ZC#N#S/AXGJGN.WRabJ5RW56AUB\:>bN
T:19H5_O?L-b4(aOO2>5][/\6P_P337XQO(19=5SK2WN[6<@16=Q^<5.Q;@FI:dD
HTQC]GgLf==QKVRLN30dYL1IF66=<\^1<#;TfZ^KdL,Hdb=JIE[XGe6JISG1XN[S
\,6/+2Ga9NLJZ,3-TY/[/-#2.U.SLHYIcKTEB\O<PUcDWKYQI[;=(1Xag>#L#TF+
]WY:YCfKH74KJTaH^(f,Da\UV<>b(NXU=@-Ld#]dD_Ud)ZG4V\d.77JFH,7O/6B2
[J\/.FKMg32a\MZGWNb?/==_AG/DIA[8@3]C^U@[:b[GeVaL?Gc9=g)7FW0g+ea^
)g.([HS=a<?bb)TgQ/,^(b<f&A4#=38\&1g^&FB=3H(9:acKO-d4Z^Cf0LFP.bFW
GA?YOe13#[0823-g4KPF<_L0e=JLe#@F4M=E3I4Ob2-[fY)Z3(;cR4HUFW&aPLbE
eScO+&f7[[e3E)g:0Z8R_4YHL?N&RdIU3O(D5^#KDHaHVgF32?)gEAcg(F>G8>f2
VT7GT/[D7a63Y/5@2g8:Zg#g_O/afX:[&F+]PP.[b0<?28^2OC&2ed22#_H8P\]A
]ZZYJ-K5_?PgL?67b]Y?UF2Q/bf5W8HX.I@9&cL>2DJGK#O/GKUSeI(C3:fKd-)D
@Y1KEF\E-U&8N3^a)ID(5^W8HQVX^,\=M+5ESS846+:#0WTI?ZF4bLA>J?;QQYe6
^1.d?SeL_af?H=7gF\:N0B_9DQ4dIaY&]gEY&W=^aT6N3X1TX#59aGCO)_1,8_.O
Y+:_N0#D-c;4U=4OW1,P741L?,SYG)2T26WBd2-I5.^M69?42<c6TEEL/Z67+PC3
@XQIbKg:9?dVHE#>))+\=QR\:#8+&(X/D<>8T<d>;<CDbKW9OHQb)CXG^7U;OIHC
Y;;,Z_9I#V2UZC0YRJ;_H7#?PXedU8QRAUZ60JeX_C&CHGU,AL#EAeZ\VRV81ILN
EAI@DcA[,6\5??QI43[-7Hgf&a@QMAYP0>XfRLPV<^.:(fEC7\NbXU9DE2[:+XN(
1Q;2@C@(<7[4#JY=E^;KSd=LX1,/U5IYN(9KA_HS]d\,TP?R2AFO]9G3(XRCbUf2
g3T<g+8I)HM<84OF+R^cIZ)0=6ME_9K0:7@gY5BP7;ULN5>POQ,FL)Z>,Xg2=YXI
8=4KaLfLI@N>N+2.+94&57-M_c1eT/YSJg0:b.ZJ@E/CGC]XFgNZgHdE9aF946C2
)O.aFb(U)\K<BO>G)fA9g#EcF3<bEcFV#gWYOJJ\UD>.MSBMVHCXG&2#3g4E+/E)
14d(-J3K)gE;cF)0_LK>aM4YDa4]U7b<3+e_d=674M^=_0e,J^UO0IH<SCZYTfQZ
[&^Pcf4deb/\8;NF.T.fRf&8/YMg1ff;XVTDO-7c]gCT<(@^D.RROZK64(I+>@:W
NC>^N#JOL03U7faG65>cK85R7W^dT_KO_TRLQaa35Y)]dJ)U\Q]B45C0afcUDCP6
MaHa.7?UaMg:?H5^-K&5-@14QT)R@U)P<MK3(M,1Zd=+V-e5T,EDbV^:GTTbW4P<
5S,WE7>4(g(D09b_Ka;M63Zg#O:;_ZR:?Z@)d(DL)KO[.;1Za@J<b>g_Ub?FIWaU
W,OBRg(,_cI^(UY2Y\]O,f/d33/;48J>VE8C5cB19I>,BTdJRWLf#UD1^4S8Wb_9
0GVC5MQGgQBO7J.@6R7M?[II_:)1WDPA.0=O]/_Z38NEa++M\<_1deBT>Nf@LfE#
5K)/aT&ab]ggU_+<_M/_2.ca1J;UF?1-a6FYIXDSg=bG)[T7b^KP.F(DI4)22<</
cdU^.[QXAK1J^418YJ<?Ad6=-P[B8;@BI6<+3^fIL&)gdd^eLM4[SAFKdB(fS2cD
DTY:fLM,L@+E3^(e,=#DHH24M.5JO+DR6f@_fLE7H\P9J)I#cV8O.?,S>#\c;<6D
KDg#I+RINJCY5,_^e4:R>IgbQHdW:dH]CN>+&PZ[XgMf5SU3_3YL,?.2bOAc0AWT
^[?&94_Rf2b&Od:_+Bd<c[_3@U,??WaSP-8#E6C39B#W3A;R^?:I[#BXN&LD2_^H
9NF@+V=DR2TNGG0==abc)aV+3ceZgb\M^gW)bBFCF_8fU4=H3RE265KTU)(LNY?W
]W+E;U5#.SE=Z<)^,/O;O@B+QNP(W2<R(b5JgM4Ad=^D)D05W)EM\GILMN2&2I3I
(8M]-a3RRF+UHA:<KZT:2Ta747,RM)E,_Y02E>&E_/\^Y]R[,La=Cg]g8eLfb<O>
<=)L+<GVM+KAf(c-GG.Z:LXR?R.eg].H=c:FUD0Qe?D\dZ5[=M_3#ZBU84,69]1Z
8S+c+e)61:<S1^DHa4[CI/?.U,)Q-6L5[XGZG^#BAe@f9+,3F&R8RN=2ScB.HF\7
Te#LGGe+T1:?CbXb[B/58.OAA&6f87Z:;9XLeCA?IF9gb+B7EH48GY>9-S^THf3?
G).STB0cgRMD2cLEMdNbf#P_DDNR-J@UEVQbRU5=SV2=DVQ_UPgO=\fXePa<\XRL
2)7cHcJ4A0=M(FR7UBKgIA;&HH/,4S/EPD^;-<(2/:??d=bY^V02g.K#T]V7gC6,
6;<Ng2;5;MCABOBQJO&KN&JF1HS(9HYB^+c;D[3P3OS?A6+/6B42P)-KMJXR:?>3
ZV[:<YEV3R93g;)0A@MT_2&c^C@a]&-W#&:YdY/@=8<T3d6+P;T3dW.ZMf0fPf=C
)KQfTN-d3I0X<;7b;RO701#4A#,>PTg(4d8EaNC4f[I5c17M=S[>/.FU.@d\PVR+
LB?]<b0X27VaCAb]eA\0JFZ9:BSXQ[(eR3Q7^(Z0W,LA50Y[>Xdgfc<]@.\?)-1=
2JWg26C=,<f#bP5/ed@DcV^1IFO)(&DFV\2\+/d>M6]TAR_SRbYYXN46V1Q2cMbU
DM@4BAVVg0g<REc;6RQ06R1B>,WBEW@GV#H;3dN[^eJ;<^NX?BGI>J@WXP]@O@PH
3:1-7?-GKI9Ob4X#J,Y7R2M(]5:c/Nf/aeK=V)>G<dQdV:Y.V>6ILd7(A5;DMGSM
J:(8G)K5W\I=\6P:9H>a:aR/FARaL(PFXZg=KUc@3,U+NbSO377T3]IK#Q1:b7=G
[:_P9_Ya\-70NW\&@^>&UDIS#,TaB:;>FB#T;H3OT96(2]1N(GD[.cVgZKP):VVB
OLe2B]8M_aMP9f>\@^-]PYO;[]1P>TCZ/.3JO,#XYFY73#L\WKFD;__+8XUI4379
1;SfFDFHTT.B7ZQX()3U&@2a<=?/<D-P=&c/MfQ\=.c)I?Q,:g?D4b(dK<CRH/^S
L7476<YV/)](N#P6HQ3@N,5795D\LJf8)3V16PA7FHA8]N.^7IXfJ>.a1;?3f7D)
=CY(;?LH,N17\C\LUI]d=RSRM8@90ed[V3D_7W:Xb:cJ@2G=bNS=9XM2)PNb2g7X
?2_b;Sdd+AY0(:CTW;Y-#?9>:dGT?0=3W@bUEdTH3>3O_3R:F,0^S>LK4;de4^Q1
PSG9WO-EIZRN&\Cb;U)I/A.1KfU?_CUMXFK.[/FLT<FBgUbMH53-:D/R]BRDG.:]
F^#A/JG[:671)F>c2TSFDUbJ[N4;9cP4L0ORD])(@@fUa6>ER;fY+V<^9+;Ef]>=
bJPd\AFT.8dG/?1Q5P(&_CQdI-^\Y6XSc\)SVd#dUBSUQB/[EbZ&5Q++d7:KS]Z;
Fe#:B;S+[YT]0ZCXG:6.4]e;TAKaN=0b1eDS27HX^HSgNX^/FA)N(F8[_Zd^H/RZ
a__=D9I#,?0:cLMRP[c41[8&);<=5<>2dfTI+^TPD9=#@Q5P1[&@]XcYS\Bd>]HN
E]GU0+#1R];MAHG/;AH-.5&K2:SQ@>?6W3#BK2\>Dd70Hf/[D=TOe[Kd>dgCFVeS
8(0KRZ-B(g9-B?Bd:FS<P9.D2WQLVYTZ9#PI?9TfB65EAX1=fD(E06VS.aK6Z)O=
\YLWI?WXeQ/7^P;]/R9042@@P912?,2OHD\8/YL_;.fCN\6M,=U,OSXCPA_f>7&U
FQ(G+Ea].FKf8IHMTLP\df5f#R7(ScROT^S_/N_/QcC<[?RH.Z@->Xa>Sc5&(N?.
BNNL)Z87H0]RGYO6VZb=[CHdXf)GHQcJ\9MC@0TLI)&@OE7V=;d+f8Jd5,cH1+)E
AK^,\1\-9T/WRQ.6(O@DB]^fIU+8JbI2.YV7\.U\J^VZd1\eG6&HRR3U&OMddJOM
D9L<:a62=-R)T@[TZ24@84[^)5Z)L_?0M\,]fXP_89(If-X(Y8e9=YZ3:.&f,DC.
8S^ZdQD?-^J<1AZ6S]Wd4JGE1:e0KRRa6KK/,SEgFZ);DXfQJ#03#BcC@cOA5M]:
>77A]RfgDB+<;CW]RT=Y9b-J2WWc-KB2,[b)00<PIO>H82EXB1THfJ0WIVAGSA9Q
HPS=,XTecUHC&bd2ETJQ,=_(#?.5WEN(X-SYbT5U@YV<?gG2Q;\T7^V;KT\eg>UM
dG6,B;-GT?1&>Kf-^b,fc?=>/.)T9B(K>@E?[0Z.4@dYL,5,HZ.N16Lc1AJWDb>J
XTPUR>Y@fN]JI^ZD(&WbNP-B4<(g0c7^ADE0T(8YQg+g9A<>&I0-cB),#;O@gfX>
VA1;W@0MB_TQ5&BMJI<-\,U2-<U(UEV7_Dc4HD0DAgPO0e:eS..X7dg#BO_e9309
Q89IT10:=.<65_N7Z4\M]F&>PbLO2O5]Me^C\dT7\_+];@Od.>MGQaR?,BS9^PP_
(+GUWRVBOf3M&f@RcaeKVRbKZ[8X\BP9(Q=3.\_1:/9_Meb^H@.GYIO[?Q<+^\@^
aA.+X,MR)A([5:._&9MUGZY8/#c.AC.d+ab&bENa4N7G--7?64OY23+(KGT33D5B
+,CZ\G8gV9,#GOH4(1DXaG-ANC5J:Dg(:<0WX&8/K(b2.?gP]:9(+B]0:87A8aHS
P^c4@&ZQ5dFcBdfS,9fc,62Lf1g0[99D3?P:C;V5H0L#50aL=7d0\_aNQRa;EJUO
R4?IL&;KGCIdLO76aM/SY#M</9gI+@2O[N2;367gDVD(+;GIV6Xd71Be1\S&5fD+
QP^ASY9C_X3#[#3+:Z]3#3&/#ZKP&MHZCcR/dF]TWTXQbbO9\4L2HfVBC#SDPBg4
e>A+eI73.10B&FU(b/;+:X>&8cYVLb(f.@>FCgg4]0a99d.Z7;;A3Z,f1FGP0DDP
c=60U_I#:LcH+cAWLDc?^bFZfWUB>#\gWN_SNReL:_[SDYR,CY/HB=H/Te.B2U-W
?c<FT4gC?D;]fONXg<422BW2/^^KZNI9=+89/E7dG-DYDf]S(?YX;SN(R5]cME=E
5P\WA1JO9M5RY4(P/>c09:&L&,[bf-(,A6<,Ce]\Yf\FRf=1TJ+ZBL#(Kf4RYI>)
,O0+IB07@dD\-g(G._<_QK0#F/U00FXXFZ[<5;@O\H-+b@GT6Sf?//b\aT9M\XMQ
;Q:A:aB4V_Z9>RC?;:eQ+]GXH(.)&^[Bd:4Y9FR2XeD4acXcaFC4:9HL7c9,>bFc
D,6KLBadZcAK/FR3[,H>=f5#SPBQF161AKfca&Z(=[K4D]HX0;IcVQVH-71&#EId
0@5GSHT-e=I-)b,gEVe5:4Sc?9,<1H=^X/FT[Zf2b/HXK/e8NSRP14W:NMC]b1Gc
fUe#c&=?c[^1HbecYW?9V]CX^Z&^>:,_28/1#bGC]GCV>??;8(b5H@dMT(9-W#N1
X4+YV2[Z</]]>D;d?-(0N5fTBg3]F[_[O11((F<82QZ/fH^7O;##A0aLH(^,^Ze6
,O9+&SeAgIb5O.][S@M/a8G/JWg&82Q><1FV5Bc)E+HVg->U2H9K;\M7AL_O_V\e
ME?0fdUK2OER8+YICSHCOS&;-,.^EK=K_&B<T2?e_>#cf(>6D1aTd10;?+YM+^P)
0:P/G1F?Q(T_D7LU>g_Y):7--d/WF(W,8Y22.U@6_[@>eYW\AIN_>d3.2J.A1&&4
>T2XdXVP/?<0.6c2:[2cMb60#],CG2;AVcfN;+H041FICC9PJ8=_[_U/]cRLC9.E
+0K+.L?KUHR,?+&fD<L9H1)TV:[-U;9)\9a^_HFQ[C-E/;09\?KaD>Ef3<[PVZNH
:ZG9=.MT6=6cKa&,EF,QdVO?8K;EA:@V296:JCgNL8K0_M\Le4R-&F)Me=@)DNb:
E<Z-Y4bWRO(<O9bC4FeRKW<#HGf-:U52JIQYg[.&#CN^-^Z7Y?^/8IBQ?+gH6E46
UM\CVaZ9d&\([\EL\TdZ4TI#N.?KLT[S^_@HE&ICQ/XC5T9a,^TL_Y@Bg5:XRTFa
=aS<V@P/@K9E)K\4Z([98<R?GeZ.<&)c)LZY,@859-Nd_\NJ^]fA>0N83X;&,YB0
fH#X10S4U@,M/S_1=,D&O=fJDDRHIWM298=]bYXG??2>[PgE+cNG/JEY9E4PDM8Q
AY;_6ZMd:b>2U]S.1H\>S.X+^D+C:J(?9ODFP5a-+GOS\IIWWdcZ?>P>a66d18=a
+@5Ia?GK4F(EC9O&ZGNEGMU91)[B8BFHe@D5_?[^/BfB#4V=NG@.6^18aTe[cFVF
TD/GVTC=^9)P6S<<e+2-BdU6b5?a2?6I:U7_1SQN[2F.MF-#/^Q.<2Z/Sa-?Q2)b
-#2AW30H+ZQL;]60:/P:Zb)LbS,QD3^KEFRPX[5T5121^88Q?eFc_Y&B0)JIaPc<
_112QQKWe.LF_-:T1@=a62Y6B9WRKC-RJOg.GFJdBAY#.W=?1+@08FA#L<XC8J<.
KYGREBXNQ=XS..NE2L1Z-U0)MHdW@1aXW#+2F1\>b^YZ8Q^4GL--26O/C,@c#<=G
P;@JBS8R84=;6?(f8[WJ0-[&3R]4EWT:U/14/?dL0M.KQ?Ff0GT9,@(W+<BDS=4=
FD0MI0MAG(,T.EASPY95G5)gOJ(KFFI2NQ10H^H\774@RIMX7YUT,O_ZP>[bbKMQ
LG-9?D)JO25OD=2VI,GW+8Z6B/RWUWe34VCV=R-b;Ug<gN[E.;7=KY>P#H+@AF3]
>MGJ0Ue=b=&ZY5FG1\5_/OY5:Je@a0#\9@dF#Q@:Td7]^2=STF]X+e#=O_AG[K]E
aMH:^9c#(GHd>E/FK&^BN,cQP+)>)>:=SI,MDZWg+U.8:5NME\D=D#8RP3E3eJ97
ge>I-0>#cf.P@-&A^)GL0eAD&^Q#-^Kc?_1:YGZ]^g1a,>1T&@WJ.W3ZH0>+ebP<
Z:Z/&PP[Ya7cGPK)WFC#=VON<g48Z#:FeGVbdPF2N-<A_YZ+/B4D-S61/F38OeVd
e578T_dcJf+ObJ+>:6J^(g=95-3UKXIKXO/^Se8c@IH@B8Xf<\cFK)8^WK.84XbQ
CN1+@KWT=9XMI#6I/^(89B&b,F:8Tfc<Q@UU1@bfY_ZO5B=:[2O[?)^W.JHN;#37
/),JEPT[a_[e,#/+<O]DQ?OMF3YSPB2I25&=_/[T6:.fN)5dQ)DEZ;_;B.CI)[),
QAb)T#aS#>QRJV()=+OY,g?P3g:GZ#PY&c:L9YQF9([NI)I2#4fe.\AOAcB91V(&
\TLY^??Ac8=F4ZL0cJY@Pa.+C-0BPF2+29N,\e55.c.D1)_g-KaRHJ6\^dgdQ7SH
J6aH9,\BG.^G_./:98aLU.6TgAM:C3<OMU5:;+_&g<_fA#:[2T8Ra_<fRFB<=L:8
W1@:aV^M3f6e\Fg0WGaWHg7Jb?^U9\CE0dP:.?X30]#0VUaPAge)d#C5O<>Q+ReD
#L\/)U&#P,aQcN,W6EYE?1&B5?P]B-;^f1+O/LCON.gT;[Q[?H7@7QMU8fQN7Q->
-M;eA\P302Z[O?EA./1CU7VA4gUU3PFbYE7)PdMFCOW6#.I0OXYE@#XD_./@L/>g
:;(27eIU]WK=7TG5:3;M,-4SfEE3&KgP[gV,3FFA&<A1:67cTH#S=CMJNE&/SFP/
JPC3U-<VXL0e\&AQ&TQRZ__GL934H]<SPON5-[OK>)-&I&36=aO6?IHc-;:[VRVE
<L>+Y.5T.[]>D>#\((:X_1P-_K)g<U\];9P#ZJ.^Ob(N-M_aGB<T(OH_9CCF_CS-
BI6U6,]1?ceQ[;8,]a&F;@ccVbdHI+?O0&=N/I3N2D(H:IB&8(9e@TJA)Q[_AMBU
ZW#Y4?60PKR(C]P&Ea/6=,0Q=@HL>SNP8bEI54A?YdcE3/P<[V(BXNg[)A:/F9Pb
5[DXLW=^[ENB.ODNE.g7T5]Uc_F95B,(&CZ@5/MJ=V0:e0L_KTXSKbLP[9B_UM,#
2MZ<B00W,(F=WPRbV<77a.M)VU[<C]0.HfG73IX6FC^35?LDBZV6>Z&\eAQNF^:/
gJ>-8SSHC5O,>\g9;@^E,0NNTFRd99]@gf/A0\Y5+T^6V]CALU19f>[G&Df0&)3a
:7MH@BG:O6Ugb[IM-8J1_9CLe,\0FbO_W:)Sfac[_O3KIR,_?^5H2aI6,>\d7;B+
4cT(.MT3:SYL):M:1C6<1^IUKD?9FIE@V^:3KE29FFK-g-aZc:6L<cV>/?XM;../
:[gV\b>;MCB3Y=58X?aX_5QUGOJ]3/[9JQT=[-=cVC,?1(P?^bFPCVJP6U]L2WP)
C3+CLS9M9\/OC#gS4H,<2]bL>:C#K;^^<GI23b[B4OOZJ/;5:ULQ]cTB,fIO]XVA
TU\H44\^Ce:>gO26E^c-P6;3U7<1YY\=7:P4=VT&_6FE&3APab+,L6Z/^SSX6;(M
W>H3V3\,,4341Q]],+LV;V6TFdQGX=,3Z-<+3LW:)4QB@N#D(^Z9(7+SW5fWa7F1
[/R)E5)#.bS<g.6-7I33,6YC?]22PL(RA&EH>#O,b/G)#-1&gCeH1a(L#_Tf=R36
0L)AT[14A1/-/@Bb3d^WS;[>MO;TC.Z+Pc^W+#fd\8OQaD:4bGZY1;DH.gA19\0]
Jc97Y+d4@HDS\^gPA3eLV+E_VURKL]H58E8MRON16@_ff8Mb6X\4(GR2D;M+[M2]
FII8U=(0^UPP^4_&)8E[LCXe<T@0U2P(-87fQ2[\,-\d<#d^eJV@@IE\4&M:SPJZ
W<8@J_3@<(XGKM(.DS^L_YHIRN0gL-V,OO/Ag;\0e9.<YUV8.(?G(7W-a41Q1d28
#U4]OFe&&F6HW_H[3<-GHLJ]:_T5PK;W(^D).=#e.dN?FW[[^S+F;U[J\A;NZ9RO
?O9eZO:]<c>#]T4.J6FCa:Pb_#e8W\YJa^2\^:?0UQf-SMA.R1[,GEaaee:gVDI<
>/^d8L(_RD+?W2@_fe2/gV:D[TOE,UQ^Mg6,/?Ke9\TcLM>?RT,1^.EU\dFb;_]W
\VK;<#T:a,FRXYF@23e-V<H(91Y9(cQ<eac006M^O-4+]985B/E4b[I>X6RS)BS(
-?:H;)@N5?DZNfO36)N3B,eXPb2IW<ScRf&fe<.OO>b,,91#<=F8ML80=H(+]6)=
4K:B9^DLI<W-gQ^+(VbN^;2-6aKRG05b(E45[6gQ3+5[I,@WeO?KB6XV^S;:FZ8E
R>Q)8P1J<1J0@+,_ZXH&8S_34#L2SaN?9AS.&U88S>\_4ZB8BK)I^@cg\N9);WDK
/U(<\3>MK?75LH)<O@QI^dBe<a?YV&L)PKZZWE2G;G?PM][RHR^bU:6B8IXdLX;9
=2H2X(4]>@8[SX_XF#G4#^.3(J?+H=NQ+N8P_T0=H1;4-T7+T84<WS,J-fWRNE#&
6b-#8SAWZETPTR6,FR3?#2QM3+N?JVb9+3JH>+4741D@6BM_#5A2La1ORdC-47P=
b2eYe9>H6^eWM;IdbMP[_>(eebBJ_ccIFCW(GOJG3WFG4dJP^R#24Xb#a]gNWH;2
2,OJQ)F6ASSB2WDSQO\EPdd\\cQ7_G95Qe55J9;=?6?b):ZFEQKQSH9d(2YI5:J-
dcOTD7T_D@?aC>b19E-4P3dA1C[^WLJb8H)b?/N&@Le?O?.0AOLL>_HQcL:RII\>
<JJ^P:XEETGG-OOG<P5-3P<(?c&Z2-YFPg3F;/AV[88cL?>G>TcUG.S1aD;Ye\#X
PXMKRGJMNfS#U>cVB>R0ecO/C-4DE9]R]/8]>;,[H^cB(e(^87e@9YGVG,5]D(\M
G[]M__SJTAU=FZ&f,V3\.fB#W+6-Q((SA=P.JZ#RE7X2@gW^RA3YAdAXQ6)9?,.A
g1D1cY>V,8M2S)cH_.bC;9\(J<.HKNZB0F]WMB>c462;/7V;\gY<<K[0SYQ+#768
CJeNQIGC<U5(RVT7JB9[)D3/\;dWI:][6ENeESER]gXWbDD?G-V_;9bK<HHXN5d1
UDfWH.H?XR?5Mce7O>>b>;L(d@7dS7.UXTJ-22-OI^?Z:e80XDA4I&G1#We#\(+#
C0b4IAW-KA^JF;KYT3-2H5Q/TSTXFc+4Uf]=</e5?M6\>RbWaODJ4N5ZYbJ)3aDY
SA#R<PV)5J4U5eeOTC-.&R2I&F88Q_56=[Y@Y1YaN.7R#U#@W)M_e=@#J^^<D[R(
1WD]?^B9a8fS@;DE0E;[?VI?+G;HgO,,&KM=e30\\;(.\5+dTW12aTS)FaTH,ZeF
LGS)1;.R@O-.<8]4dP^ZV4IAaE)G?Q)M2.(#O:KgYW;2^96>3g:=3LRf9D4GgBUY
MJQ5MA--<BZ<N1^S<eN&XG=1U+0K#/QAe>cH2?_@C-JaOJ;O]F&T/MSFaEa7Mb@U
YYKMC+SFN&5&J=6WQ<DLgW<7SG]KY6e0>>A89+ZfU(g]CNH]0YTgWc.A_WRDU1g:
8XIcV>>:K?BXf&)(G\2COC5+A-SOI^.0,5Gg\,A[N-PZ9+]Q4KYaQ3LCMKfN_7A,
HK/ZSV=NJ5(IKD5ATI9L/RS8Xa6gM^+0If\1MX0D\X1K=2GLSTg<f]eNNMU:JO85
46;(LR6I.64GI4DG?VG=d6G9#OUfNCL-5@1_0\)cfDP>a)BeW-BRf&/S_GO/7\GD
g0fNb@I+NW<TgSe2N3S.A/N:?P.N\d(H_/F+V#BR2GY10TA8I1/?,NN@cT6TO8SR
g.U3VNY0;>\1Ldf=a>>0\eN.1H)+)FJE/>SUbNPY^RPNVYdeI3(<U/<g7H=.bO=/
S+P<cP[\V\._-PKX&#YDS<G6W\S_Z3edF\AUA^GdNGWCC>D)ZDIZ(/K;LXU9L1QK
(B^gV\Ud5YH(cbA23D:-C]N0[\)4#[N;9O]AUUdeJUR[T>N-UQ_O953eF,Ef)KKZ
(,-X8.[6;5>ae\1>EF<^AC?&P8bS>W]^.RHXLHT>f35)(c8FZ>H;VU?b/:L#7\g7
-#FW_g]DAD:C,\.,ADMJP?VV:,&YCQU</T/AeV>4:S5GM7dJ8@BW<EO6b4@46ZB7
QSgBCd&G7A_Ue;5SS_JQ18@SO;^A^5e\)+:#)I@#N?E2UOT1gACF3Jg8B]8aX2V/
X@YTbL6JNZ>&dJ6UM0^fMM01B/:D@N#5Ng[NaPUa\FD51<&GMS#Z<591),]^32NP
cRAL<1cAV:#&#[1-/P\@(-BQTc@=EHfSU+W?c<_CP#Q8dbcZ3fe)RU7ba8\gE.(L
I8[M[X<We/<0<N=V-DNd9N#S/fTTB?-^0dVfD^C3fbUXIW>4E-/G&IV902NW34+2
9728Ed6HK?R-9CO?a887\)g<UZ=3V/]B;cJ)O31&)T,AWGfac>6>[#U[T@ES,EVE
^W9&F^FQ_[Y260/8-P?9aUTf.,:_-K8LfY&.CSf+?6dS3@=.<^^4_/+-c_62^A1[
PN47Q63X_=/]&L.dR0O)HcWX,(-91W&??a5P<)?RLR7R<+HK^ZGGIaNfd,;DZ[+0
H>a+aO&HU@b[M;IcgLEA:.:gIgg;N\)[I2(+3+_5:BTIfbF_[8);_0KL?JO8/;b6
SdXKbX,ZZ2TE6BVeS?+@6EYa3<5STdPUd\EG3<TgU.ZJ=JS^Z766Z85K[]RRI,+X
(T+F8YO/GfAD;K8#2)dc4V_=A#^&XZN<;H(Pg&f^H?RcB]GV;;PX<+[2PO^RZ<27
41:0PPKUS#<.^\S+P^-U&;;]EIB,,.2G-?cg0YDQA_?4a.@243#1[]8.8(@LBPG#
b\OC0\)=BOVgXMJ4HQWe+1@82_3/IB0C3[55,.D#ZNWBQ#SQYg:SAB3H8ZSQ9aKC
6GM.)MNA&[F#CE=Q<B#XJ[F.))H;d#66I#98C]QN;=bQG7&84R@9=-NSg1[3#VBE
W,K:-_XS1e\E1P9SYVD-@2cP.\?ICYHECQL:8FQG#?A6aL+aJ(ePS>LXfAAQd8CP
1L)93Y9T=8.HMZWG#-G7gbc8P-82GPdVd.UQ,_W8e>AVdH^G,@?[a3=fB+Y<KE<b
[XPTaa_J>1&O\<LDB6E7a.&;U-CI]QPV^UbE73g0?2+^13EJQ;VRG_]b;c5a?H.W
-&S8eKFe77GQgQEP(b\FI\]<V=0,]FUL3ea7I4CJB/4W0]F#We0-4CQY?QLaGbQ2
:f>1g=&KAO&E<JW]1?1)=,/,L+,5E+++8\DXeAgVdPJDNc11VaDW1EDP;,K(]7+g
9+26(A4EfRCR_/X4+BC,WgI-eIFCHa;ZN:#K(]eXfSO<;#WHaY:..@QHZ,[7KU(A
:&dW+^.S9E9:B:HD<IBT1;PAW?G_<_^_0Y[;.gX^696X>P(O._ZF<SZCU)Ua3HOV
>A;9>9.YL0;H1<C[U3>>GggH:_J8E?LK@Dd+@HebVI3+U#J<Y[62EYD7UT[]M+CW
0gQWRJABY38:e@:DLLcbN0));<0,JM+];D+DcBNDNO4-&80RCK(6Le.\2VE=YXVI
-(dA@RXA;X@7D,RaRC5DP2EG84gBSB;_L-fFI83\45E8MLT@N>^IF6&GXdIJIYTS
OHTb1&5&6e60_X<M?YSG5&?KUSZcNWTd[I>ALW3(QF@1;dU&7@<J^(Z72H^;9.gY
E[<e(4[#VKIScK16@[H2+)?AR#c^HX33.1&-IH_P@XGQbCCaeIa\,B^=ZX03>;;e
A?03I<MWJ;c0gCa#X8E])F4c6G.#bAL:U=Q5,1Z7^-WD<)HER1bTBg[1>X1WH35I
X&\B6&V=/XIa;4O1QKbdX_;/8)=J#g)<O+@?T[S_#:_7JA[c)\U7<dU7c=IB)((a
@S3g^BSYH4OfdO6;8fD;:\T96Q+,A9LNH(+a>c1B4#Yce?[&DM3M\b09Ffg,#XWd
1:NRcRS0A<YAN&9>5d:9fG+CLSbCKWZc@;98[H#05T(,]d@caZZR3CBc,LXdU.>:
?5DUV@@&ZY51-_IJQ\3XK7>e&22UGRQXY9Aea27L2Dc22T^-EGDM8+6+aO1JJ)HM
([>fH<[Q#DNOLTeUH^IRH.1Q9<)X2Od+e.</.#M[Zeb)-VK8>M.A2JE8gJAGS,H6
K]bOUI-1W&5:/U2G^KUbf-E@4Q8TAK#JK:]Sa0>Cg-MK&f:?1J36L[SCO?AUX7XO
c@Y8aPfJ7.2N[P2@F(#_K#/<)T5PPX&?_02d?XDQV/Q(PXgC(M=VN.O/>fV^Y#43
:S-Cf((<HeNQMcdbT_Pf@aCg-N)[((-EIU?FU#acO+\5:.Gb:5/c549e@O(AcC,/
=2QVSOV^H0[@3?&)J6+Lc^e6I^_E_E9R-/APfX)QFBG]&/,HAK5PWZD:M&=TL)3]
e\X7_MGDNALJP85HFP2f:c-QbH0WPSDJ9b]IG^2O6,L#4/K3C(B?JGZ5>/T3KN+D
MDU^;>R>-H-;LE2.=XGT/STB+b;IgE<]]fgR16JK(6HUHV,_3]8/66M=9--Pf]:b
>?H1Hg+8A8#-,>1BWLUY.A/V1NLO/:\8,g7RX;@R;G;NQX6T9)]E,NI99;c@e:R8
SN1OPPb3c>Df]_94(,R+cg4\H@S\O_gZ3]QW-(IE#8D>>O\8cC5Q9CQPTEX@#,5]
,#7]5Ta\FD\@f:9WV0H[dO31HOQHLW[=1C4=_7<O.>:H8Xf2Y3JB>S9NH;ZcH>J\
G6]gIX>A18>.(F,8LSCHGR66E^#X7=6W<VZ[U(e-/Q0XWC#b6,7VMJ#)37TfXU2,
EKB&^a,@=F0J&3=JW4L9^P^fFT??^Z]H)MY6?5ZfU52GNA^6a:L2V:XN4)67HId&
6FCP9J#.cS5W&fNE92^ETdd=cKTGbZb22[Y;U5I)OR#BD7)3.aL624ZQ\(KbK89[
-F]^LOB(fJ.>)-)L3[6/VJ[eO/P\[5QKfGe0F#^SAAbY5eZJN+KFHY5X7JKW+GU6
WMeVLa?&T83566]H#Y?4ZVdHHP89TcI).QJf2)Vde/O,>9T#P<SRgHEEY;>Y>GfJ
&Y#Z[W\H@f7)Y&c^L_0)X,#GXWeZQ19<0.:4=Z6\A78.dG=PCPa,b^Q2df[Q+I<R
a(Z=XNZES\)LWG3=da@W([dNf0&B5N3:?#e))If.8>[9RgZVBZMNdMU2RXAG9fW=
g(1AQ6=>6M017[&J@Bd]X&;IfXF[E]&>=^9UN^AL?./bLN_VJ5<S^ZHCDS6.W-6^
>\Ac/Qa@=/G5Kb+1F/DS0#bS/7?d4NKHONQMCfJC[\/[^8-SgdMd&U155C/\JfdN
g<D<./TIb3aT<Zc@#3\,Wc>ce_.:6V:0F8Cd:M]>0P&^I+M-XJ.F=(D6&1BD3[EK
5F:ZR[eZQ@[C+eEcE+]<?HV&FfaIX+cX2+8BTJ7C_2JRI#0QaN6-=)37,,7:B.M9
QRBg8OQdeEMbY^+JPXE>/FTYA\HWBc,X__OK<M)V:IKG3T]4G5Q0eKO=[UaJ_>CT
LVJdX-,,M_M21eDTK2?4ZEZ=.>EJ]T=^,10]N)]]IK+95\(:2EA(/J7Ibe\E^34W
X?NDJNf:7<5U+3G1N]0CX4c0+RC/M_@T9#6+M(8Kca@B)&N4?6STJYP3=FPD?13P
<@TK,GeY+NF8g<bV=<I9+E@S<>a#fPZ5M8eL:g\6#KB9)EW.Z_DG(/e_AS4FNLI[
H5SHU:CGZ0[=;G562MaWeYRFfI9?VH\Q[Z2U(?\5@JMRd5Wb/KN43O,(.Mg#&=[O
bCI_;6?#[22<V1YJAf4dX52#SH[cX>?NU>HdI?93FK=.^GO/YT^fC;LQ0=_D^U--
,AO1agdXZ;_?/:F9I8=KUK64V51@\F</],Y\[Wc#c.K+;3ZSP3+J4Y8S;dQ0V_bf
f\M8M+0-[,\/d9B>FS9bEG)\ZAF-A>ZO,;SQ426>RfA^E7[?^T9U/d(H>UJ?Oa)L
);f[NCN2MPaBTeFX^;3AL;N]V)ef[fHZHAgVg,DXYLPO0)5Y5U@?H:N8A0-<g--f
G+@3@]M:K1W2K[9(4E\Rda0PDWF[LF99D#Y/3-K\M#Q;M8<Ye(#+,3ZHBO:5I22f
_LEd#bg1B=XYe:J.fb^SR4V>@@-g)XMIHZ/S2)\&O-D.@LZKAG3Y=>8X>XCUTX8:
0^6PcaZQ)=G_<NC&<&g:N@_(O<GO7NK+<XO)D[^2e+,I[fK(PP@F,AZ_,(YEQV,6
VWM^@)G2JDHMb@Hf-(AYfM4AfT1+D[2]^]C9bAWWZBGN_E:-30/Q:+Z^@PdA;7#Y
MeD,5)[>V,QEOF(#GL9W.[DHR>1>?LO2-e-Q2Q40b\4PP+/5MOG/ZaIA\R[WLHV6
3SDaRZ@.7b@O6>+VT6-P0JcE@ORH<0ZE+5SdZ[.)A-C#B0eJ-[d\PMN79G2XM_J[
^#J/W]TL:MO[^BPFMTF9S__PF3O/TXK:?H^94bc3B(-MNZC6:\.E1Mg4>]&2Ze=4
+f@(<c/Y.+RN9Q.W]Xf_N<?,c;D-(VT5Z9F(4-/f5a\7,\:89:4+SNQ,gN)W5L9J
b0EMPWG(-8:XBgW#XcW&XN.;2ge/0fA:]<P=33;_3_WfSg,K<7L.Z[L/SKc>B.Y7
c5X5Y+O@cJA;RcZUfVaN<AT?P(4OKe0ENF/FQfG-Rd_b1NI^S?d5IUI_>+:AFD8L
5Z546_;1.,Ya4>QA0?1(:fF?LReV.\b/N7AI#7W.:4+,<2H(Rc:gDR8T(:a<GG;G
_)<H1XN9YZ.U:R7090CH?A>cER&2@.C:F&J./^c211Zg:e0@V(>6CE-a7]\S7:_F
dC78#.C]#2bOd@<4421bQH6b1g5>,&8?^R@Ve.d-U;.Sg?@edU#SF7McP&5#B<70
L6+X-D1fPA#PCD\5JbHT#AC9@E#50)T84aPW,V\,#,;I=O@DH8<9fR9g?7BRJ,I9
#df6)S8HD.,[W:f6VfF,)P7(9d2O<WfNJRU136?cA,PeFdbHIV]F^f-Agg)2c5)c
S8(I9W4Sa?\SI-&HC9Q6=\#>M;:bd7)X(#S0C-UZ]_W1\0.,)-[AM:&7&eN+QU=M
DaNEgBMb/W_8)/I>=_X=QZ<8LHEeUQ:P4E/T[-]Y(bJDdHF39)7\3f8PK0I+]Ac1
/)^&F&PW2d&<7-c4,feD_CJVdV<=+IS=JPMCP_XCaRTK?P,9\GPFH9W/=UDB:6GN
+BbEgO;8.P=+_4&_YG2R5&&Id-N>=7Ge=8>Aa6#BQcP-U.0D=Q)Kg2RgEg;M8.f.
TZ=?5@I\P@.XF(ZfL6#:J1X.cM>.5\W-EG.;d4.UHe]fDQL_2e.,c>J)dS9K<;BN
^KfR0-2@)P7&Rg1b3X.Z1#K0IN/\2e;VOSYUKA9;&-CaQEO8c)K[c(@/>D-]D9:)
eJWTQ9RXU&,I3)/H);QRgV-6T-[3KOD]GU)-U6=6QcT:-Kb/)a11GFGfZI^V/QCe
,SLVUFY1GC\JC#+Xg,beNAa[,HS_@=5BSgNA?_-LWE909daAFNbKQXFcQUUR46+^
T\g4:E+MN@_g^8deA,O>^L[Af5D&1c^_7N9)H&/D->S_TE,NLV2gK9+<c8F_:c7Q
O@]5UUIXM<EL],Y^B0AF4#cOR(66SOLZRD0L<DA+,f0VI#A&HM>a_a^Ye+4,OE@X
:/c?P?+2E-YDGFDgOWD.L(=[XT\>Zg[1a5RPE3Jc@919\9OL^2557(;4I@C<+7NP
f(3+,&T2>B=a(N13ZPZ(B=C2.,&K2?5MV&Ra3eX^97E\Tg4&U1HVS@(][4Y>;8.b
H8>>L#Y&9O\Y@;F_Ae\?C8UcCI&EM4/aU@KK(bRVFTW4G\CL67;eLS]1I>A)WO,1
e8Nf1TW#fKXQ;g0GF:RC].E1Gc>JC>H6##71U5^4_#F;a0@2>G@B]T3S^2[e8#B_
UP6APZ6Z#[/FY-&e(/03Jc>bMKD),CTZ#:ZG1?cMR,aW31]@(^?[28C=LO^KD)f]
bb+__&c&gOV1b^#Y7;#cN\03H4K?MX&b2,DeC255^8+V-&Z5W;c+3=AKOKIfX)JL
V1K>06<<7PA;H@E/)QR4E>LMC_Y2.LT_fBe;4J?:c6H5Z#/S@7W[-V:R1e-BO/bH
gT6>@0#P;&/B:D=7E+=dA2=1XJW6)D1V@Z:#3XO2#e<>Hf6]XS@cc@U#g^+D]@@9
^D1QDdYQZ=[-MRFR:]f^&?+BX(=K?=SY0XXa:WW4^)\fg[/MfX6A?7#))/R3[QPA
_L1M7Y\&MQ.KYIH7^(EOGH=Ud/UWD=KM7KfE0[@LEYC8I]c8M^KA#DC=PJN.D)TW
B;:HI7[M<f3d?RI8PSU+Kb?PeFdWPXWR^G5]:9>97fS9EgF520<;<^;G1_3)BE;d
0YcVabC.fbJ;AAE;GM@g7+A>#-@8A\:6e2S@EYR[aTW2W+FACO?O#M7C0EDM?bQ]
ECB[UJ4IS]R\=96dA>aC]dP&F<]U@[NW-aC&Oe1=X+:aIbN.#Vgf[WfH@==CFVZ:
PY-NI06(FQ:J1=<<,N6&VC)80B7^UZMC3Z0#5,K[A+a<82LA3^,g./+3d:2^fgbg
4?a5EcSKAdHCU^19g9+V@4<5_Va?:1gG?V31bcY6H@/cQ.LTOd5>0A^Ua^5U@=b2
T<ZD.08]f4KRHI;4W>1/\&HLL1aKSF6GK4+7Y.9NYC<c21#:b1<#DM6f+0H6W.bI
V>Rgd?-TXR91@]1HL/fA97eLB+A4RC=;c&(aT7T.Td11EZZ)D4^6MeCY.W58ZN,>
?V=>U9Tg4&[06<NLcA6[MERKB0=4\MIb3Q9PaD(4#Y@eK>VPc#,fG1R9D.:N>QSe
6GAUFIA=Z7C=GDEcXP])g97,4a,)Q/0?PB2+e]Ng644@(A).&^-&d4:3Y[D5TOR_
6UO898?5V/NWId55Sc80I[aD)BfV30;V1@<6KdE2KN?6aKRI+P4G2g?_)D;?M_/b
Q8\6MXOJED?e&Rg3=O/9U8W<:JXTCdG8A)9N,1SM5&ENgd3.]4V58E.HYZ&>[2W)
b-@?+Z0]c@B.DY-OYLQ:>/@CWQSF+T;I5(/>#,HC)RU;eGLcKLSf/.^M/)V91@eZ
ebcaJ+GX\<8?I6JD=[6A+-?1b(NX8QV4TFZ0d1-:<0(K48TOJT^Q-_@+4Q3Kc;a/
8[R^:aSX]D6,1Ic>d/e#(dFeGP>93A,:G.gP?ZFH]fe+3J/K6?g)1U;?@)UfIYS-
I+_4^^\:6;EAMNHDIa=_X.dgK87fGg(.(S,>><8D24ZLGOIX@0;8U,0--MX&+:^;
3R[b]DX#B]#cF-^9,]7B0/@^=?d_XX][G]V[Qbd:C.:V0+(2TI6HTF\Yd]/Wa<aW
8+)O])5N31>S,W.L5.(4O.<If80bT,&IL[AeXB=?.BJU-74Oee,Af#.7YUK&5GGM
IW4?H.7@g&^(FX76X&>Mb8&2>Cd5.=UO.cdeaJfN@OM^56+1b)c^5,<2=DW.g=O3
5N\(0N)Q0?IfUfU4@NW?KZ8L\+^[O5Td.6U-U@1\]X(a\_a?/UMJ_#Y/4X(L_6<M
6a.QA5VHCZY&7ZBdJb9/V9[V=9EZ;ffZW@H>:&IbH.Z2&#ON5(E^&S1a\DD&IS^E
K)?dJcCR?.DOY:e;XT6;8#f8\:0A2@4+f0R=ab7,J/cb^F0^./<Z)Z>B&0E4?H=A
b\@>HPPVT?C2JH;aRU\;)Q6.UU-e3[Q3H>1+\C)=c<<1Z,Z<G7NJ3cN./d+,Q5M/
ZPb.RW>/0edMcA2->X(,<M8b&G^S3DbXWI9TX>G=KR#T=a5cB\b7O?N3=DWWc8aY
9NN7+AT)1f0_L<_.6Ac=P6_c;g_1Q@Qe+DWT7ZOfR]=cfW,@-.OBEOL^(_^_D&H\
KOTg(<E^Ic)/6G;@\<9L>9PK3\0)c/>?T8SOB.I<abZ,Z;=8(eO;@<b8^;LOf?XR
Z]dg]-SX5H6M;S=:L&Hd,(0>cT62;#27#0a0#EK=VH8M1LgPW2,:)N:+:3=9><LX
8]0[OEU]SH--Va/+&<QS&<+(]Sc79+.ZVJQ#BCg>Sgf^U,gf01[032S@)/-IXK8-
SU_2O_#.gP54_Y:BEQ1DT,_S=K&JEQT)PH;IL_L\Yf[,SL+A)gaJ,.O..1D-\]<6
^4YJ6CV__+O1J51ES:>MT@1,W-TgeW;:.0N0UM+G.P6DL_MYWAg4;Sb0L)W[TBBX
T)18U<E&4GPfK#4YCRHM)QZU1a++.CFDQ.TXPHFSQb,d164eA.(=TQ^dddf/QZMO
aB43?/:3\a9@YR<([:ea2.CPagU1c[4:)WNV8AY#(Q.+c4/;\9=68T=J._a.dcO0
L9ZRZ0dK,P&Q])8D.6BYBKeM<^eW,-8<YM-bWV>R6TJ-87<b?//FKd(a)5aGWWME
FacIB,b:#F@EV)__[_2SBL_U8-a\g+ORT.(_\FAKTAEIAJP+dbD#PD_AQVVGBXMH
@.DOS-0IZ)1]E.#&+&[bV55IM(,/4dF0)Nd@#:/[;IQ1CJ#?Z&DJLe+915JLbI2#
Bb84I=Bf.(E@gJ9AXc3,&H=.fQF6Q5-IcBNF[JLF<H-JK;]Y4ae@R/4S\B4^74G(
T_RS^)\?&[B.2V44,ME0Za+L&P9,Y0X4=YLGD&d.+,B@A(:&ebXbVLW58,6gK9eO
8TF?LHLU2d\_2CHge4F:[V9G0ZJG.9dV,R&_]9\87^8.L]BS>2;F/g@G>ETY9/:d
/=Q8a?^e7cAg^OFd?C4\HWc<FK-\F3OMU/V[&_>?aI,#JgD=2=1@LKcU\Id:3Z2P
JJUU0F)2\E+A+BAXG_bG3_BP[X(^OQF;42J@[>UV3^^]+6b6&,AP8SVW#)VX2BUg
MJCd-Q6HU.)A>);HD:Cf(L5MX/P8SCTfD#N9ae0#1/a/59.0BEXEZ08_:.,Mf?f<
Y[1S8V6T@WfD?4>6^bC.aK)_9K5Yf3RJW[:6TTb_FNF@,7g,/?\3T#<BZ1M[f,Z7
\]g>LP4NdT1#(VR[U#FAeIg0UY#2XaTf2E?/Z>@[JP2_f@9ZUMUBa<=aO<7KW6;]
,0Ye#aKI3(BgLc<41-\V7;VV<VA6<WTEFY\F-QZbIP\NTLO];gg][8g8YY>\^1D,
_KH_d@:_d?WKR7K&=5Q#1,XQeL77-QV?\&Z>)BC:?bOa+dE(X#BQ8ZV35(f_9d34
F]]c,e9c&Wb=/Q?QJf=+=?DN;T]NU9\?8fTGSQ5TfHN7C=X+9RM/)2+-PPPBe(Od
\fXR9@ZN:H_5[=-N[_@F2(\=bZdTPf)237/-44D83&[>/,UM>Y9I,T55X9@.^I-V
>Ie.Z7])Pg[[\0N^Ka096<<YW8[D[e5Ra#1_?YE42OZ[NgJ?BHY/SfE<M=B&,Qc+
RRF]&E6GE:gEdPB[S@.@JTg@#fe-f.:9:1CG6O?V<+0Z,DT-=<J/fW\\dOc7O-R<
UHW5\Sd1HQ1eE^2XJ>^f5W^(>O+H]?SRF:#&=b0X4PMB/4+Y34fJE-EK&A(AU+I/
7B)@IC/c@HP]/4\dgdX9#,M[J#.8:TcG^Y.D?eDbB<PB_N<@OZUK,a=^C<WSON.&
RE5607VMN8/E17@NF2;baV2d5;HAX]d,bE_>/+GMb\-#+@3S77?\aJQXX.-<b=^1
_eBfH8N.3KG<M6:ePbM;\5abG#LOLJ3@+YN@c/9OOK/ca>48GDRZ5Z_3dG/9=dRL
A=PCB=Eg4Y=C\LMebFB0BPW_9]B)@(dQH5@(?+Kb.#MOGSM]@&FOM/GVDM0&[4:Y
)M]R?e:d;d+KRGMLWGd>\NQA)^9b5/KPfTU_9bH.I<]&YY:dS6OJ>AgR4=U)-[QA
eI\>Q\d([aN=>a(_)G-L(_R[YP;L&6U3Kf:S6.JJ-OVe8I>();E64\S0cY/PdO43
YLTfU@<Sc=D4KLd0G<7I,OVYP+KL+B?-3HUFJGVPT[e2_A@G>S&NE]A[+Y8Ab9MM
&&dZTc+T=eGSKe\M[]f9b=]Q<>cGQ(^9ELSZfAFQF;NOD]c;7=I==W0@Re]A;W6>
bL<:GBIEBf=aT@)4.)TP,I[O)bIc;(DRD21K\)8IVedOa)ULW8IIfG8=Y,L@CXQd
S35&7.20fFZZ<H+-=:(/cSPUH)eW1_,3.9.EJES.bCdT4;a>6P2@[PAe>6_FFQ#d
I=N(]\MIJGR?QNJ2OcYH14@J_]O3IP\1B=S>E>TXdR:06SGf#Z\>NKeOK1IBcZ/3
66aEET(SK@=A[JgS8Q,@F#J1[M-G<UO.5I)UYeVTa)/QY-)6,_AEG_)(-7(2DC:H
X/-J#ebgQfEeS0,1.W+#?\gQ=\5//FgRa@3=QBS^S-93S\D@f6O#I.dUc@T?4)U#
KfCaFc)YTIE-^Q^CEg:&M83ID#^.LB62B._SN6+,UPZK@XN9KBD2b8XgVS#G4C8_
KY:3AScRMJ0G8]4De\_=5dK9gQ,[R7CEZ&3(^AYeW]^TQ^J6LK@IX(DV)+5;[)Pf
fXL>1HJQFe[(/<JJJ8(Bb;K77@3\b-)H5ZfP>M0,+=\a9+1S>NZ=R#BD81-MTLB7
ES[X_>W552YX[L_U:(-A1>b1S@6</Q\S9>.^^f&eN5=CXLLAf[VgZ7(E,9<-Q<XB
/K0G<K@KC+^54:<ZHN.Hb[P7G]-6Z;?0@.3GT4R6PC>ATI+O:-B:d86JKR0=S1&V
\[2YdNVg@f/#+C-UU8L)NQ4QSd),UZ0XN]f28K#A@>,Ucg1fO94C\Ve5,Md//]N#
/^?Xa949g+&:Jg-96MU\[G8EJE1P,EWFDGEMH4GGRDJ)9:W/gg#V;8S\>LG_F?D_
>/]YK_g]g9(]/&DOY1/(fGC<1A:)X;I>?W3Q/Id]C=>\CO_>Og5aD6C1fcb<2.0f
WWLU<f7(f?f&QfG74.4&g#,@DB=6<Ye09EG2aZ-6,bVF8OEHQOb^W;&aXQ;O_U8#
T7YbJGQ(IIF\2Q\A;LGd0?]58_UYAbAAAE,/GYAO,O_O<A4G#aFDH]_YY@52@<H4
>,CM.Q81XL[[,F+J.C_9/<3LW_#CgP/6<_7F\eP7.80TUC.&=2b132@Maa;^fUD\
O/>OB1E>;DUP]L4W==b^Z=&:>YIHE^H#2/EN4Q[)G-;cReF/)88N00YgAM-=>H-3
HZ[<\;[eaGYZG;N52-Q3,HBW\fJ@aKe46N]VQd)B\_GF-OGI\+[O9I9=YKVZH.E<
#/ZSGB<6@Yg;91HBXG=:_V^dH_5UEa/^N,U)>Ib^LeBVBg?X.Q3,4_)Uba]e>ZX0
gIdfH3<+-\JD0Y=Jd=aX@KMLFEJf^QO1H(]-N+gB5Hf<->_g](.g>FdSADYGB-I&
0#82?8>,(#Q..A=UM_JV#Kc16F@Z)^5Z]e6O=/NM;U+7SefIa&K80(N7[J/+2TU3
VE>-GO7J;3?,eAg]Tb<Y2H+@ZS<T8[A?fF<6R&e99F08gZJ>BK?cVN6.3PZLgAUa
f^6:fMgKC+N>LUW^_cGX8+_5)-T<+4.Y_CD<PTdBOF^LYH:JO/AOZ<BP)eg^CO^T
R,cf;gUCX67.VGPEQ?RY[5eCA9d1AO6/A1/J,,9:cF;82>cF95N,B1_5KZVZ3;1F
b#<(ZN:42HA_OXS:&0XCW9T6>;T_Wa6+Y1M6\=;\GQTbLAM7ICQ^4O/I.92^A3#@
EGb=\S=5/-UZa,GE^aLZCZRNNe;F+1P4-Kb+FQI./,TTI-1W[@03@bJ_2J6(;^-I
3U#)g?,:2;UNS1#C&1bb,C0>]\CVPfLI8a3^Y>MCNU;QLe-WA,[Lcf;H@@X\I[2J
?QNY;Z7#@acaH3_0CWLd4O1O<9.cU[:M]KGPe#X).X6\R:T&3(_/YAN)A8b,d&dT
(Ta2;A=UATU1+dTeI746H/6(ac.>#4f=SB4T4:UL/?KQDb(&F)JQS2E1fRZb:g[D
g,U=Y4[Z9-T.0d]Y&,7F4ZLE-U&bUN9eAX.U/d99aG=NN,27+18-0B+[TVdOPQFW
<#dGE.5JC65]&(NE/H#&9CbR,66-;4\+@cc\RK#96>:[eD(;ge;KV3Qg](@/;G)#
,dW;0gXKB/fg]@L[KPP,V+]gbP4HG/&c9g]F5IYJ6PIOEa=N(0;+f_(DAcWK//7U
-2ZI>WW-W;0fMP[:4A9B.[[H-S(N416&=L/BS.^U.MZgS=Q0S;V10XP?GgLgU-M8
\<TY65aQ>Z7Y58VN00=Ab8QY&&Hc2KAbC-1K)P#PAHY+e5O1ea=?U9]M9cI5KGH;
15_^YaB5=DU6JH,5>L).\6UVZP+.5[_MgK^,H4/A3X?8)T1PQ1N/A.@+ZX7:.(>_
Nf[WF+17Yf1(Fe(a7[ZFF6B7I93d;;f7#BW?:LcO6OJ7d&W8@[22^[ZgS><UJQVH
__3R7S]&K;DL:aD6ACaHIKaf68g>^G6JTQILH=e=,W66J,,I(Qf@Z^Hg,G>bRc<D
aJ9<_a8a5.57#fa<<]^VEg&Re>cIcF@N7#C#a6DJA;=cABN<Vg+I@/K]Y9<Ka^CA
0Z>9G(Y=VJ9VV6-U?>DJ.S0KJL^I7\1L10Yb\5d>1X,T9+6R;>53-]MUL)ET)ZA(
-:NZggae>Y1Z4/FAFegT#V]eKZ\c3ZOP4X/e@7C.-\2YP5Gc>?5gABUE@\J,F+G[
:[CAPc?;1Z<8LTMaA&W:+V6A1H?9YA/A(+?+T6,9gcKf8SXdJC?9B6Y^37)QRT\X
,[X/WM\LN]TI.M;_GH(S@2,+FH<JMO>55[&#F[4SNOZF/V_d&ZTgFScSRcCIZeDH
X?Zf=NPXDN(RDG-3R#J_3#5.).CV>dI9:fBU\)TS,GT2B>=\V?9)M.5(9@)\W6>G
96)4M5AF,,E-A7ag5;f/R#>\)E+9KFGMaD.QdV6NGFeS#eW?BKWWQf50IHaOVV-#
-DZ4dN^T72.DA81H5+Y,F9?;&a@&838E#1A#7D)//Q,KW,=J\IT@\Z+_=KWH]_>d
f+fOL/;N@DZ1L[>4Y0B,X+e=/2;H\AdT#+R(aWLE+e)B^2[V_9IJ<bGfWO<4M)(O
;&3+L^,OC4P+>g<UJ-<PRB>0/<L.ZC9@AF7Va[#aMC-g3/7LJ6E:EI.5d=(ZcVAU
DbQ/R]f-JX&(WZH?S9P3;c^,c7>22]+U09#VHU6UbO=D2g8TJc66LL(^LWES44<^
NI@I@Dd3VC>?4H=/?K<;+S9(4SS_c8#8Q=Y&e12J9Wf3@[27ZA/:Q\Eb@LB9Z<:[
I87=25/C;@b6SOJ39#3[FNMbJ2N[EQ6PbI,.A5-XZW.:_3HIRZ3eg:FG<deX^+,X
^OBaI+1@a.D_L9?6W3.gM)SF++0FBY8OEgCX-R/?>MQ1LHfJTf==S>47X/MVOBU6
LBQK>dc1/a2889MAY75V,AD[#7=5;.@[;#E7G1YBFdb^5F/CH\.X(@86Xc?A&0:0
=G]OP,?1K/&)L#+gW9PU:M7,:XZ(MCHKaG(,ZRZ:JKD1C_JV0LER9M5>C]YWO-E\
FCf_6Dd,+TOYTQD8=P+GL>EV>AR7&BbBP&@;Ud;BV0?<N#S^beDU,&DbSgNgUXb,
BWSXA,\YeU6=--^ZY((f@+6Oc7Yfb4S[eE=V4EfdC<G+U#a@EX.S>19]4eEZ1T3O
)WUKI]D;1#=^S(Td5UKGaO@-B8)W7X^>eaUR7&&3Y;44fZf.UdUaQJHG+6B?M2ON
.-[#C>B^C:(GK-]E+J<ga0a1[Qb6626CL3bW<>b8SJJR3B@9B,QF8c.6gB-<4C>+
9+?ZO@@P@IXJ#[)&C(dWE\-gA=Qf1IZ8]HZ:-YA?5BV?;9TLCD61K95Ye(8->Wa#
XL(_&6)J3(\MCUGLY]PYB3b,HL&O7CM#Y0/N2C=H4M@QZc\IT.1TQ8DAQJRV;Q\=
,Wb0IeeNF6^VO\?;WR4&&772T6b;f:7fU34V^:-TG^(BE=2/Y18&D)FR8T#\F5->
:.->H)-4M47C4KfD5/SY6;.;5Q/KV&-SPK8?4f7Y8-JZ\L5#ScNG^f_VD2LO?e(@
JM0V-\R4M7gd7a-L4a)5g6:^Y?)#d+_H1f0H[H0O3-<#9\0;cIY(aP1_Y]=OXYR\
3=H^A7N7)8BFHfB0J_L\T_ZK2EV0V^F@V-g><,+PT(J<bYSTQ6G?4I@/M]c)<>N/
VSI0Q[a<T/9[).]bFBQD;>>=3@I6?4RWfK2CM#?O1_VVVLf7a49F,[=TgU7ZBQ)\
a\NcW]R3(P+.9<,ef(U).;Gc^f\QR&C9DbCLRH\5(6I=6>e0Y]D:Ce8>QDJG\fO:
f/JVAP9+ff8f#ZNL[PVL.G3(eMA@E:6F8FXQAMb6#]7&?DPR1<W(&.g3C/CM(5IA
8XgX6[8E+27.E=#dbPY3CUF\4VSSb[+]HbWIEgN85.T(S175)A>W[A_8gcId@,..
UAAW-&>aP@R?-]H@[6JIDfEHSDQ[5USA<OY\>d(A1(5[\Q#Z.=62eg_D55IGX(g6
e9DBN6OE+3RUSa\UgM<L]-4Ce+^O[^,(?YVAQ])B_5,U_16>=VW^E<+VG_;X)Z:,
HP,LW#b@g(HY0/\V(PY&J1(Tc/BOP&aR?+d17IXL@0&FPQaAd]^:X8cI8QS0>6N(
Zf]Ue&0bI2e&=X2;J=&KNd8I..AF9OEX-\a#O4PYRH/=A)M[?H1ZD2WBIaIQ0[-0
ZYE+45HOKE9_9_COcO79)JGe^<RH/=9?Y@[E;b,OfBJK1c(^1Ab5)#Lf/J<V=&AK
(Q2fBAbeUePF.CLZ3-;/@?LS#)/@X[KJa7RS;??@(Re9F-@H^#:BF4V@N<JVAO6G
)5&>JK<13,&;FQM/I9VUfe.MZH0FD1U]ZeLQ3;G)^8+_);PbF5D@^\GJHG,YG76[
S#EONfQac/K:14d^7Z6=HaG#KDg.XY1EL5-UU7-)+UKa5DK./9N0\]MH3[=]05JA
eY#.^I,dB\O]M[d(0GUg]I8Cc)U.WZ^ca31CJ^K\ORaD@?2##cU/B9+fTIR4&G:U
CHUa+P[E#.]K72dPQKXgUYQFAc+(f4WO6)TS3E<Y9M;NSB#_I=F^[OdY;eQB56S=
^U0)[/6Hf(34A.?,0UFXM3e][6W942(J1;BaF0XW:#^d5HYe(UBDY?8VG]WALLBZ
MR&dU]>g2;gdSRWH7<HDK4gOBK^c1OVX1[)(D-_N?GW0406Rg;#/Nde@:_C1]LB,
,BSM?P/6,D^,6<-EXbU3TASO>SOYG@9[bK9JL)#3#)?2+5g]X8\f?R6):&O:?&?0
dHe;+IB4fKgQ]FgUXLM>N/&3^:d<:@aO<OdWG8G41b+7dB/V<O]@U@EJZKFa^YT]
SUf-IHO54^\H\+6Wa+:B<[0D(?aG;bF2KJH0]RfAdWM\[6Y+/(;]d<Na^U]BfN.8
;[F^P(P[G8bVUECC^:;N[#=):F9VPF5TCe+>4AA5T,WfU#S2Uc49bg/d1FGDdI]Y
;5HeG.QOf(3RD)?Q>\WP[#HN<1)[g\4(LC&fAP7;5CO)E\RHTQNdGYSIX/U,4_d/
UY,A62;E_YDH2(T789gO>?;2D,W#P/7^LF0TKM;K5]ZMPNXHZM<LEOXeU#fe2QQb
2+_g)+&#bE.4=&Qg]3CJ^ZL;]180[O\UZ8a#QD-g.>8Q-ELacO)b;Y#3>1;WN[cV
3Cd=e::-<UA(])0X-A2@>P=B;U_I;5;KKd>:FU\=AUYdB503^CNLR\8HE@,_G[^>
->C&<A3[U6_b8X#M#(DH39WZV5GQFG_5OI7Y.5<G2)a4CXCU08V<39+:IH]-A6c/
STA<H+/37-:Nb0LC^RL1(fLc.PbTb,Y=1J&db^)(0Lf3e6[)-6<<B;BB?./MNECb
b]N=Ke/GH2Ug2PI;#MEN4gI6#5&7_bVJ2,,.U/NP0H]dK[g\W5L:V?#F,ZX-07VC
]JUddcNe1OJRL-&gO8[[13gdY14O7-KRM^&(OaBCE1Gc5f^(P/-,b)6<W:L?:JOE
VRAC=[5OaQ6E<<N>#3X3Q@AS88C:@&=C>K.+H)QHJFSK<F4T9(,7M23VUSeD+&.<
6F,+_,=9T>E-3,X+\_9@VM?(WZQ(49?/T[(,:,cMT:DJ07Pf5a8aYR9H8(><W@;W
)6E-Wc<5N#g(>VQLb^>]N<>B/>+_9Hf:c#EN@1F5Uc\^gaE^4Wc5(7gOP;/I\#F:
##TdA],=]bfN+H-(/F<2M-KFKE8R<ca1BK9Z#3S(L93UXU^6dS3/_ZVE5e2gV1QU
EXX67_b9=UYPZFac5OL&>8@@.a490^)@U^M<A6)c:>&NHc;)#5SV_[J:#1Q;9a,7
.EQC5CW-^KU+a]^7JbX?&JD+Z:Y,;PH^]gQO&Ob85>ZV<?a&[RbFDTWB+5T47Y&=
G\0OWRZMeDL]bA:)D\>dM8FbRUZ<^/-dd)9[LH3eL=#D3HZ.8(;U>8BUC8K-PIf3
Z=_7YagO1J2_ZTC2^R3EM[)g(88_E[7@b,>C+a.Q.M01[I]Y:-O;g(a:.8.TVE6e
)]/T?PV;HMLfJ2^/NKP(M6MM72))U7UeONU4QV>DGf1a[WXJC6&6Xa]+Dbd?SBA,
fbcL.S]@:d:_?g98CB]W_,#_2K:5S/[Hae@OY]QG1KZ-7Ge+]5B?>]][WWP+YCN3
J&V1)F&<dUK(OU1Z\=[VA4,QcF9._C]ZYcY061f;ZE8P5FMB9HZ-0Q+MK5X?,:#+
;fQGc=f,RcI-J5eVCE9KOb-7JZ>8#ODQW.19g:HM(7:ZN9Z]QA(KCZP]WBOA[UD0
#PG+(4Z0RP5].=^SC_S986Ab;a7,RYAY80FP7b\H0P-H;OZ9H):@2BVE+dIG_5dL
G?NV0TTVW0Z]JYWg[B4BJD_DC>CeJJ@dSJ^5&8HVHR=@>1WNE5X#-&BH^WZ8GM&A
X&Z)_[C]KH0bdXLOYVPS)2RO,3QM^@4H>?9K;Ybd#D\F2L9YA?I9=gg=MR:Dee4_
],CIGb@=3S>f=IbebX9G?C1:Y4G4F;.7BKS+J[b?Lc#+JVcQ2]9XfY:,^@8ZH8UJ
R;3FeS@?X3E+25__b>cfP5?gEQWW=O6>CM;f?N:3\Jg_ANNO4?E\YP-:CZ<BRZBN
?\A0IV1IVHI@cS@[IY5#[JU?_T[B-QLK-Y-1C_(BLEK=dTI-\9R+EKBSJKY?AZ-R
(KPTP35M:HeV]/cdA8^_C,Tad(9DX1;0c-dDa39;#ZGeE=LbD\Z05^Jd,R4O\SN<
D&;)XaTNY0J_4D26>TMR:Y2(V#N4g-Ye4#f]VX6OLdUFVFISKB:OHUF8#F=VM_Ed
I:#_,SMYWS-a?CAD<4eP;;ZM1CW^ZSHa2RL;0=+dVK<?]FD#MJ_d#I5C,GN9U([g
>^C04)/YD]O=+\bd\_)4_+87X@8::=4]AGF>bI7>Q8QYRL]LH[?+C/T/Y>0Uc(A^
@H0@d6C873CJc&WMaR]&\J_2K.WDJ6<&7CL-dQU5DUI.XD:HcDAFS<7=V#Uc(A7=
//[8;9YX9[K[K]VC-9^)B]b[9\-c(B3G.O.\0;X_.F9gM_2V\R2:H3PXD5.fD&M<
A6f7M]bd,_/>^gd\O0dR<0@#V8O,^RQJ-HN:8><BK4dGW1a,JWe7AAG/L]]AC_Ta
UHLTODY\^C9#=V,1.DA-:3D:Z32BZC+S3faMeVEYHg\8K=G7O;U>KR1GQfHO4108
I?XZ2DO[Le)fLAXAK2Nf.fJ8(;ceKNK]F8^)P=If8JO=K:Ka5:^:gOI4G@Z+X>GG
-@KUPQd<YY=bfCYMIf1R6C#G_Qf>/DE]+Q#?VG=gKYA;:IT3^J4E<b9&ZFKFE>,L
d25Z+Ec1FLcBF6F/I78<(?LK8>(+(6:/fCM0&>A_H=:2J)dJ?:/7DbFEfSKgOY=P
UMa<-=/U-UY=W6Q2e9;;LIK>RO+JVOEZ6B/L)E<HH,B:A>>B#fI>B/1K?C3g5IUK
cB7#U1QYF_A@YSM12Xe.EX1B?-6@LCZ+_NJJ@QR]C.3Vf_TMJ-c<BOg=.Z0JC9g-
g1XGM;49[gUf;ODEGdI3R.XYA8X86<EJ@P.OI@J+PMW\6YM]ZeCTRRS[b45SA?(>
Qf:YH_M:RP(QFg+<g[?65?:]O=aHKOCJZ0^N6H4ZYP(6VL.1NYT6bdLKBN8=6Q:K
M56_?-<_+8f2<PRQG;J_\7UAN.M?OGNWDZ]DK2e#PPcUFR5G+a??8Qc#ALF]6@_Q
1[(:>UaIWP.ZJI.553>B9]&=WKU[A^Y4Q(C)2YW99NccgZI/=3K5GTQfO29:9BWB
\F_FcUf-IR_1W+FVIPI9=QfLXC,/e3S\2--c3>&d5W<J/TAW(@[CT:)K]=E;M[31
)G-H96;(^NS.WHBMS+JGR3/_04RDgCO#)(]P^^UG79NTA:>7C\9abDPJdUfE<+KX
M(RE\MB1XUGV)Ne&?bXYabH;F[QI\d/DaY.Q[]J)<))Mc_>G.F?K6QaT\WY9IG0)
28<gK(8g+\CFYL<RINa5]MD;&IL^JOfPSK)_>^XW\b)MF)@9-?H&H4e\B_Ge^.UI
.PWI\Y:=O/Gd-[)<?A0ZcHK[T9WCUHBTWH&++X;3e#d9FOKL7/IH)9dD7;/LX#DE
W9ZYWT#<S8VJCI:b_LH(8E04e[ANf?4M+,)4_OZ@(64Se\@66.A:+;B7U3,ePg4F
(/SaX-H+&N?-XHRbL#^P^UG?:R;X^U1AZIR9#0b3LAP^8(A;.b]RK>#)ec7=CKJ?
B&>bC#6bM@4g?@L.QdHQKK>f]g^KZEHOP;\7USYKBB><@\B-C[V,HGLYO2&.WC7?
Z[J]]a#L3-<F+?6@QF>7ESd2e#;);)bDTHBKbdC_,-daba/d<2XU+AP(HERA5:Q5
(5X/TKM>g@(Yd(c9=:0\Q<9Va\[6bagbG_F+A>deO5L]D6@,MX;_+GHB0Z5NQ,O]
[V:D/R(69+#E1fe&0:PWD0Lc5;]=:0KY)J]SM&C36-[4-_MXbH_1D(7=Q8=IT8db
NY>0RM7QMROUcDfJ+A4I&CC[eVLAI/RH],/F^I&3R0L/AV_/KB;f_5MfY>@#D3H9
/\a6,]97eLM/DdC)O6VM\G4gQ<8NBOFRR4\HH]088J/QPL@>dLUTG@1=ZQM\,ZbO
IOc7e@0/IXWPbM_g@V[\__]N#e>BN7S,W/D3?&<Pc_@\HS07-HR0eCWN>/-_J5OB
2b?=@XOK.b_/A^<6C[P)BA@E&(@LZ/\]cZ3QV=691fNKaQ\Of9,#O#[2M.aJJgG4
P9-aICZ0\<.5K>.GBcRIFXAY=H9F^/Kd>#N1+KADZ:;PGfRRHJf7Z4::fK=QK;fF
-L-2]]V?O(:T_7aKM>WOLGMH7.?=ZLKT(8O(A[,4+QP/N.DNRPQI1#K-MUUc7&)g
OF<W9T2MXP9e>^VRJULN;YZa7a)B6>;X8,X/V86>8Q1G0T4:=<5]EgX\HP)(T4RP
bJJ.,P(-#QQT6dATK-<6ZdP97N]LW=P&^<;56O;cCM:1=0E6[_:2Y43WTW^<a>8T
>e^ab;4]g-]CT1;Bd;d^dXW=IF?bc^\HAK7cMZ><,_4EY_(7#_</eTXEZ<HF7MW#
,K[aM7;9@JfaMcX;/LP\/(9\Rd(5NI2=_N\[2N=7G@Mc0aJEZ::ER[[_K:Xf1d);
56O,+P91+dC,V8_MJZ9NC70;O6J1?N<PFRJeOecS_R.3OT4&g/;LK1-T7MTdTEF3
g,TV\^e(W^OVK4T?V)2U<Q-)C(;0-20QR[8L7/OP1MDRW_P?3bBQF2;/g^6,F@Ag
?H;J2gI?G-9,W9[?D]C><AI>6bG1AJ1LIHV1UO+<Z2([5+H9K6RB@aVI\=7QXa\P
c(#KK>#.BfaUP&V+@J^/,OV<LBdg(&=Fc5GC)J7TO4D2Z21\#.1e\7=gH&Vc8];Y
^1ZEEAM&:07EOK-5c+&[)VcPXT1@LYEGdZ.Y<>W_)7A=/.O.Se..16Ef\SNAAGb]
(:c[<;e^Y:PB[9O>)#XAX@7SZ[JOY/P&A[KS29>R<0J^2dec9M36SQ7#aF]7\MIA
fSC/(#R9bWFD.-188)X/1QX.F.]NP]VK2:EU;6cKR7]^DZN+GTP(P+9L<B0><QOM
8Y6M8K[J?^YQ;;><KJ+H((\BgWNA+c+7\[Z-M<,QeKF0Vd??S,H^GR<2b2d7S.e-
E8X-43Y3fNXfOFOaB[UX+0C^d1;bA-&eS+-JPc@OJ[3Z.X^C(HXU=d.P5b@#A71V
OVVVSXD0(Q()R<L][X;bc0,KW;@6_#PO\[Ba]eQ].GTQ]f[2\3=WPXTP2.5T5)fF
^/+UKVW/:_4/34FJdGdd3fC&0KgQEf;OeLX\85+aGD\NGYFK8AKH&/3G23TE5>A]
78bRgK;>E5#.K&/#6,_#R2=W\I^#&7-A7d/f@Z]XT0g;@O+M]/ggM=#2(3A+Pd]&
5?2:b>Y#3;/FHSN5?NKKJTeY7A]^0>^VV-9Q_,UD)DS<Nc0M/&<#c5UNR8d;2G9/
XdYA0&eH&JPY5+FX<Jb:Y.]eMXOAKE@O[Ff+&SdB^<3NH4GW&M1G?C[ORM(<=)D@
[5VRL3WVeE.U1CZcH?C/b1DdR7G>=4O;-VW@R6=7@<=#DYHPKB:?/0M/IdQ<;;fB
L\)Tc+9dHT=d;7f3U=1D5/KT0\cc-<b;XM</W#5-P,0RH+S6G1QHT=f/H_6I2H2g
QC:H]JMMBZd1@4Q5R-L;ZVc5QHE5D;]U4)>ALRegGf+J_B@\\)b:E@9gGVB).8Z[
[Jg)[0OL@E_c-Y@H@C)-aQ_QH?R^0c&??UZ@V9eH9^.gE^gOL;YY@EMQIBE;F9V8
L[>X#BMQO@g6,3d399&THV7#?-<g;4;R]<MRgDY5T+2LMJ,/CH9.S@\.QM288Y);
WA^\8:d_/NGdT8:1=F6PS/,:G<dB\413,&>;86V[_Z-PG)Gb9W]T[TfPUNXRCe&4
gX5]/4QJJG4E]IaD/[eHWa0BZE,A&5M#d;?F?g^@-9E&.32@dP-/>K-^cTFW;TT&
,P5BaY..1C@WM1c6\I5M<>XARK<P:OB)EaE/;E7@_65#J1?AN7(5.[][=dJ0aBTa
W;1([gDDfNEeTL^g:-W9ZbbI02g8CBG=)eX]gd0Vf^/VgN/?WMM;R4RN#Q)72Hcf
>A2A7OJTA[>\.B89a]UFUfE^TV.M_+46gJ=2:M_U@0g<T56G0ZL\Gf5SLAM>L(8L
;Z\85f:Q)@fQP5\)g3fJ:^MOHS^(&:/aF(f5bY&I(gU7@0S>WQCF[&/cD+]M;N7U
PRBE4Tg9P>@KDYQ/Ae^[_\C]PGf)LH[e<bgI+5AM?B?X)W2C]QZH,2DgMLS+Qc9H
B//2Lb]48J6NK]H6&7S[18Q;@+;eK9QaWDZC.E),DeIV:B)SBc7^+VKJP_1R5XQ7
SB4&#CHG(c#WL]FU0>_TP4.9&X^O@LGK@g[-Md:V^/5aR&H=?)YU1-^X0AJc_Cc8
(T2)QPXN9YSWA?QK+IVP2KO>HA.5d>6ec5.:+C5)H+AN_8R#7/VRT5&SE]6;;d,3
SKQ?KDCd?NWX]gI@<ZJ-ZGC=_-4#>dOXTcN@]+/&M2f6f4)(\d7B4_8aEY4aBdgM
@aNa9&JDP<MeFHJ>#Ug)<I;8&3/.JW3R=BeH(C+O,W76_PFV2ZYD2<H6+/5U<(2E
?O3\R]I__E/b/DgHZ^_TJb:L[Hc<P-H7/-@1_?dOOfdB8B-e7BTS9ZD/-:-5Zf@M
F/]9K1D+_2E\-,dO3=ZLJ?OYAMO8B7^,e\QVFC-G:He00f[TQD&U\CPD@aQN<ZM5
D91;+?QX/9UKW]63#+QGU12f]5K=@_S)4W68TDPU2Y,@]NDM(<S2g?N\eS^-3G\-
PROD<.@0-:>gMT-B1G1;ST>XN7#I/TT-dFR?(b+]#WY-S/F76_F3Zc.X><SaT2K3
U8RVSI4<L6DW??d[75-N/F;BOcM07XH@]9II[[E6Df\KO@KeBOb@N;=4@0_MBQMP
&LbZYVXXU2LA_PQX?L,c;RWL1KFG[HcY3R;/4<TP4/WH<>.R]5a9WK]P?H.b&7,5
d7D778LZ(96_^;8#1);-ZcRQ^XFLY]BJAG(W(HD0R:<7Sc22U47cf\/9P5SO5IWX
/a8+K#&D;#1XKNTV7=>BbR5&QTE5>S-WeMHabB_W;W_2@&>7XI&<YQL?LU;CRG7/
TCHE+&W=3aa=7M?Lf/L0,_=g<B7M4.)M)>P2=/d4&RT\V3@Db:,4fa)Of2bL]/-(
4B4OF#6bHDXT+,b_^dUU2N2@A5cJ4I-TM\baYe6_f(b:YO3B==6gJZ:KZP[gH\Vd
?8_:J.@X4CC^CHMY:S_P#.9^5;T_-DJ+9C>^8(9cN&#44_f8a0WNWR\J,]Z_=5DG
+>X@9I&dAdY1@^(=5.cM?W2JR6cd<.>1f?A8aQSC7g?3(]ZbCQE?HCL#O18/]IC6
/4bb=IEDe4eG3bPM_RSGCQUWg^;&&9SKa&g60:2DQ]19MbLfCTE6AE=fU.TSE-g:
]CT2@9-ZgPIYIK\V+1I)9)Y/\1f93TdcW?V>U9CX<M<=UEJY608,OcQT\YFJTa[7
#5O?ROXc,0I@QYW@LT3++D?f51BKe_N@UZ]74f+[cGT-/F)DM3R<@#(=;[EeeQVF
U]_G+18S1cOQ[I]RLM0eF:S5L]P4B(b_<0&3T@A6UMgJ55#J<,:M1-?CAW#PUE;N
TL<O.d>Z]TCaN@HT\ZIU<J,5QE9BHGZf=ERSE@1::RP@6JR7@8)b#0(A]ac\D0M9
MWbS&\)cY/e82\YYF&.PM(4/4PDB[Nea&SQ76<C:H7eJde=e]6:Tg=dP9_?ZDPgg
dV#PTW47X(3)IUK9.(V&Uc+#\=;Aag(U^^_^GBI/3(7_S(,^F^Bba9JWOa1S]P4C
UCAU@gC(-H2APJWKJ,QIXW@L)B<K][:?gDHZ7O-J<g]_Y,6+;V.W2E1Y@GGZ_=4I
QAGJ:20(/K4b298(<e:XN.e>W6U9.YEUbLBH4INb#TIUX2NTGfb)/?,&=J3/U<^G
MfUaSOWKO&C&ALf_9/fRR5H8)#].gLeFIc+A;[</gFF\\Saf+RU+b,9>CL,N)6.A
&0?RAKc),:)HJf2]02Gb:I#c&WS1:<OREX:+Y5(I3^g6Tg&FRAZ;^SGP(9O0E+XK
E_/U,:fSR?6cBLZ)g^S11HPR]:>68U&@J0.[70FG0N]ML61_<_X_V7+5-LafTZN(
eFT;&.Y7MT[.YNa0?dM&RXT]4B+95KN,5M>+M?F8EORTZYAD52OG,\06f^1+O26T
_PD9LL/N22+M[0BF3bLI9J-g99>I9YT^]a)<P[\;IWQGa1MRLB.OC<0cR_NF@>P9
EGED#((YgO2a&Z,U3X=ZW(&V,BD0^KOg?M:E@.V9\)(]Ygd4LAD.MMZ_9d[Cf_NT
OFVOOSYF;GM#NQC52Cfa?TcVY#6[b)edbU?dGJ7&cHY^[L&Xb6J_OIF/SZY+A1Nd
5?c6F6e^#=5bUe.<U8bZ]O(^9c44F,J,Q>cf7LCBHa:TD(6L]DMga.KB>VV@9cQ4
X&6HPU_Yf?GC.gc_Yb1HG5(J&Gd#;^IQZCW&F(Y//+8V)gBe#UP@RW,WH]d4,BKF
L+-U:98-0;9EV-MdL:E]-JOPJ)WEebJ#Y4#Y1UN8a3eDIGO,6(YW8+50NbZC3RZQ
+PO7L?S_);a>L08WXNM;g6./:RTRJ^J(TD7a/.Z6<#<(<e>I1e2(+P>:f,a]_X<J
;B;M/4d<c>//OTT6;/DSL^(N@E_WWCW^b>.J,S_L,I+H\C@_=E<<,L]#VQa]-^/e
8&O1+?YaJT72KC&>aCb8K]EQJ&=]SL\SbU4A[-CVHTB-cd35WQ8OPQ-X5,C,PCT/
P@WWY#S:A=3K5&<IWcK\?.f.T3)R+??AEN\-7.QYLdEQeS5:=.U7S=g+\4;TS9+^
KD7,(5JY@dTYILYXK3B]S(HSR;GL@fTg>@=B4+:XKI8K-e\0e#6W_@1KQ5aNS;?1
1-WJa5PR:;9[I3^1Bf.4<aWXXNfC;Fb&b>[4.[/7RMMDWe7\Y]ZUdG(YVY=0GZQU
;WgNLBFU(G:RF\Y9S&ed=G,V8XY&:_-G]b3eS@8YCV.?@H-GJXCYHeb^75VIE\NN
)N-b_67<_MNIZQIULO+&e<M_F;@?8MW0W=UN[(7HE;fRXYca@Oc^X_7aJ&0Dd1.)
B,.?72LdV^UMTHIIS>S;2eFV;Y0\=ccPIICHW0KL\EZOI4bdbN:J4P240BS8;^:g
dgFUaZJ5^_IK62Z&+6;SFMU/?gG]Z;M7Gg3;1P.NU>.OPb;\]YYX;L_RC;O18#I8
^]:TF5aD.IaAL3[&5+81CZ3g^.K)OXJ?MM-R6XF7_EB\C>U@T)\E]98Z?UOO-)3G
UN.#P:Y]=f&F3Qb)T_LAT[DBa1f5cCS@T(+b6+D;5_&>1eAP]3TRYR=cHV^.Y?T\
5>\>HE^(;+YXFNCVf&b#B34;=<V[T&_7&aa,-7=J^DN=[I<-8<F5e:\,H?XC#fT5
6MKe]WBY##fBO+EBA&DL^-BNaT;+MYe]/E^>MFPeb]8D6(S,C&3)(8d<;)5eZFJ@
(RMFP_^M@AZENG8@,]74G7^D0dA=F=Md,]9Ua&L=[&I/P10RM32eg=F74]M:QH5D
U7H7Z/HRM\03,M=ZXLF(MP@5R7+>:\5X^f(S@^WT=E8J+@e=Xg?OYFFfe&Yb,+U0
+?R2Jg4Y[dKZ&10J:;C[B/\U-P#BPZ:[K4W@#a4P->N83TUY7>:-UZ^4U-A4SFSe
HZeDeJEM#bAO5gg8+b5;d&?>;E6?\]HJ]=)68I4fQ-ML\DYfT?eR0CaG[)9NbXFF
+94-9E:eaYT<?0>Y8?8Ie7d#6N8YWDQ<1P#K9O\D8>LGN-QMcBH?R/:<CS+)?c5b
YVe=:LgEfdOG/<LRGW76A\@Gg8@:>Eb]Zcf[(-/#UfZVf^>&NbNM1WI#H8.T\T4c
J5C.APVe7f2S,#e)?EEBD(\;Z949>/4UfJ1=ge?L\::03H<S-X)9ebR9d5R<b3_@
d]4A-A0X-eNgETZ?MT+,JVS2#;^]Qa1EKVc8PFHKaQNf)P0I0fJPYNIZ:]QO(:1E
e#:)X<D.cE@0^d^3bD<258((C8aLb9B,EZ^]OYC&S+3gd0f,SXF@SVXfMb,f0B>?
O4Y@eQZg8XeM__BHFf51S+4T.e;4(]Md@)cW\U0;(DONTAIP:V\FJ;cf#P_]1;6&
B35NT<d(U<342bDQ8gJ9M6RH-aCS<S.TfZL\1\<F/-L^cEH02>Q5U>X3ENgM^EF2
>2VC@;UO#]Mfca4,SC(/ZQ28?@We>_DgE5D;7.a88aaR+O:U]Tf&6B)8c\7/,2RQ
31AVM0>SF(34929OG.1TI/>9RYdHS9+;d(N3I]WLI7=J:1V>[E&\.6ZGL[J)W?gV
5J=g-3dc8YcP.dIa5BZ:.D6JW_PTS+H]C4D.<:S@gWK/@=#C3A.[\K8Sded[SE7L
&>E#];6&EgHF8bMXR5edJ&g<?D<;ONEdICg&;fc&F5X<;BAR/FV_X_@]AQT0NgV-
B5[GPa[Z&/2YKTTI3M=e0G1bbOB+8AGFaL1F[b/S_f&7O;Ld9D33Z&/QGdA3C+L6
Ca&L=JT9;.YfgMD+EUX]Q8f4aO;>L0U<N@]ET-8>cPgBNa9Y1#NCX?LU5JQ-#:T8
/_>-c8#CIEJ]0@PK,6(-K;U]1RM9]<\.W?(R#HBY-2SY/Z(KO[bf0MOM,N,KI>@)
)->&7;BSK]0_5W0[W5f:AR^IV,e>1e5K7/I5TDJgd3M4:Wfd63U\-:/,7;VO.JSE
PK-Ua]KaL:eF#TWX_]6.9C5X[B+)RQZ2EBE7d29\VX,b:(_aBQ.;cU#QZ9E:9a)d
?0Vd7B<SV_b6#V?:>2EeO?b\)DC^BRbJT[0:.BT:J<NZS#K5BNW^#AfQ-/(R(-@V
AK?2OP&bW)&Q0OO&(BEDa1GP6T-K9TYQJcc[Ca>I,O&K,:X_<VE&&>V(SOA&I6bS
)=)O,FeH]8>)e:5+S2X&G9A5aT:b]XfJYG[XIaGA73M1ZL2XXSd581)=gNC1Qdd4
AG3fceB9]N2_W(TO66@VTO]O6]/4BaV0@-(71\V_ERL[)#CPQCASbU;4SB=@g]NW
<E-WB^2c89Z1SGUN;K-a70L:gUcG+I[:fe_>gWXSd5&cSRR0c\/UZ[>1g.@>bL2:
Nc^9c]PPg21KT\=WDWP.F??(;#XI0)C\-[FT>R\M^dYGFCCKUg0L?PSXQ8UU#PA_
7b66dcFMa5g1>C+N&.H9-(9PHE)d>Pe_XPOE6G4FZH5\B0Nd#GT(GFXaE]/;]90P
47&JTLF[44.O.6f_NP\068AB7,C5^,<K61)bEV0A<93)A\Qd8cCA0<ISaL[W:2g/
<fCUObHEFE=(_BG9=2UDG+)^g6RR8V#TJ?@>M;BRFg4JF74),(A2aG\>A-GW8U:]
/6SB>O65>I<J?Z]9XV^EGO8AgE^^c8JDgg71(S/,>7YE9JI_ZPK#))]NcHS3-:KS
d__N:(8IPMfUc]QVdbMe3VQD=(JF7OBa^c+K?)^:8g5=[<fe4O8Wbe8HJ:IMO\4]
\N1(]+MQZ-,GU(_#4N.(^,2#.0[G;.6,B=I0]Z;VC\4X8]F9Z:2F5QRGReOHce7/
&CMcW\\)<J4#6AV))]XQ^(6=E6@D/K59WG=+gL7X,aO7]F#R.P23SCg4IGbUN/X2
24R0];<AM\KdA[&QN1F(LT9I-G(1\78L0[+R>_-=b.62KDILS>/^)+fe8SH\(O[G
K-IN@6XZ_@[f)cNY&[;V]?/PKWOJg7]fO4MW-3I=11?T\I-d7E2YN(,#T,L/cYYG
H@dg.d9Ab+<)XAFA9QXP94a2CA/e4fP>Z<TVB>HL&f:\N(6bDBICMZX:gA+PIQEN
UGKLP3W,Z5IE<J5-Hf#M6_1?T\X(d[.LbZP\4,cC>B>J&?8NWO6[0O3[9=TG0V\\
UYT@JPcbFQVb3GL7+Q)c5X_&&IR7<;K><NLY+e\>LKY.#^DR@7VaU&-e4R,8R0(a
]QTP-WW2&Aa^:T>&_6-M<>1C)gE]XQ,.0Tg^2&I#:;\]N7#Gc.Q9VCebdPYCD&V>
a)\&4-675;#A7Z&5/OWO=gg>O&:/OSgE=KA.a[Q=_P2HM,&EDUMMYHHB:I=^Z8I4
0HV&NB[F2a44dY8b0OdM,707A@D[#b#]=eJg_a.dL-AL60&#BeR&cZT]c1+bG<7D
#@4aJX(<gWAM/8>ZVSM#UQK\L@U8/OHQ=&Zf..GR69dg@&A903_?C3N_7_a0O;UR
HT>7F1J5V:)TZZ>cU9H39<O98LJaY78K_6NS0Z,L(f6,.MJH]GCC]L-]J0=bgb#X
=H^.-HD=)[#K#4bggDga,YLW)&gYedPF^TYcG+?B5B(8+b+T/?H4HFaXENCD(1@f
5M4,KSc;#9cZQASVI4?a<4+f697ETg&;5acX3I;bPcH=)XcI#R.&@HLV?J8_-eG.
=Z6Z0/f<b][>VVg:b)Q##Eb]A3/=4..;M@=)eR&Q8fPJ,FX?TZ=2CM8G4]#.TZQZ
geB:,FTOI8F9?3(0H5\5QRD.-g5L_+H;VBBC25b@BOXP;5V:E5D.^?56]Y0e#=U\
Q&6M>X0bXfXL10M.FTe\+D&+d85Ld&J)Y5a(H?#.OIWK>Y1HB95;5<QY/<W)c8VY
bL;IP3,bAA;_DJHDB@^Z4eB7>#dEg4Q05<H:b[>f\;b5\4?V;/U]J-e-5CAH[B<9
eRYBDd9NNUCOU@+E-XI^,^;&@.8;_YK\SAUM[GZ9a47\89g&=TS]AMLWSLYLfZ0T
3]@AC@MDGD[B3Tc_1Pc>64#1aJ33g1J]HZc65c;dQ2;f-a2-^X;EP,DO0PXQe8F.
:^Q]FAE^PN\gUe8D:O;\:4KKf/LB5VfI>1[3_Q92R(<([)A8=>OD6dA;>Mc1OAZT
T^(_MV)<g9Ob)6c)E_&U1CFVU_TP,NNH:5)5[e/4]PME^cMXR9[aO1ZAXNfX;^O<
e4a[GRKWT;PaP)KGX4(071c=[WTB\_>@5-MXM;Zc?[Z?TFE>SY_3<[dJ;1YB)(Og
VQUGN4Cd=PD4BD4Fg<GRU4YH,M2eb?K#1MbIB.7^V:K=U8/=G?3+cA?.7CEXD6;,
KNgf/,BBdedRIdM[RO:8665NOMOBEPL[LMUcFEfe6SB)IB1Y\U28)X\E7Xg8EeGO
X0?4aL,()F;JM3N\1WM#bgI;QOUH0>HW.(YA0gaeY=6^.4eN(dg(;cV<).SZIOAM
P#X)TaI_(2TIM^H7^aA@:W1>7b<VL1_Z1TRO6A(?FSV<D303,8c1?HXRdFD^,];(
FDN1@W;HD1=6Y-&MC7d/4.ZVBL76-28>Z_f2&e9TP+K26FTFU+-#+[Q;G#)^=\7A
+_G7(SgG+Ue-Rf@&)c<Z&2dHFXSS04UNR2R4/FZL)Mg.eZ;[V@M;f>cBPPgd25-+
-e+Y^>@61T0QW#U@F52XJ_?:]+6#/@HK?NDe?^GP_A>.E@EJ4gaFbLQ=@K4cS+96
6QHN/8E^/?F1-Z@8NOe3SK7R1B>JQadZ&X3Sf7RIA+YCF>GD)XQfc]b0PVG,^]+?
d&@g<]N1GIG@gS@6@0D>_6+/^,JGRGeT[EbYU;c0FXDd:6,[d+aDE^2VO>&YCYG,
eL&TP(\&6TJ>Q0JQ&/W9bA7:=V/dY;dEf\O[&DRCg9SFgM)<TWdG@ge3B\D51#CF
be(cF@V_+Ld)baUCXP;^<.=;DM<aK2PR?<]-F2M>08+e>+GKU:[8)FX^B-adH\EF
=@ZUFY&V.AMgfXX9-_&[#X.T7&gRPdcS&G+&08GH/?Og4D#BgTE:gZ7F1)XGS&5C
=_>O.WUW2_AWd\JKZa/?9e8beDZ=_A#YF.=O6(V3JT7#VeX5c#9O[+[?HQcATM=d
PJbg^aG^_(MR26I-BOO^e9Y@F)F1?^,>PTAe19fMg@1CAI(Wa>ff15E8a(PR_L1K
A8,4YKMWIgN3EbOFc&3JIKRC0+^ZG8EG>2Dd_71]XA/7a5MEA65a95Y0QK#=-#XK
ddSd3[OODGSEFK6fQeb1b4NBJ8-EHZ>e_E51-HZ0+FQ=HRTd@bMO_3]Ba\U/E-gc
L@[65b9A=MBMBBPTbIGEgbe_H23HQT-QC@B#W53^C,X_AINCPcc?YN2A5g7]?#(7
?V+/[bfOag^VK-^H<F<eS_3UT)BSP40[U@6_E0c7g&=YH[/Ia/a^&c5E\SXT(fM8
<,@9RPe7T+;fZdEUT9:ZDXP6,\ZT&[IY;:@2OFH/@PPB@97CLFLH()S)K^6BSdWA
V\@C/,eeLP1<M2FP>I@7(E[[I[+E,],;8\D1deY[XV.GZHg]dT==c00.?KfMOd<?
=[>4QB16]@R^=RL)/Y>,Z.<AN[.\5Z?/J@NR884/L\9(,SG5=aIU]74_Z_Ia0:)H
]PH+bL8S]_YY^8g\AWg;GY2Y<1+I.GUbC8]52J<\OTa<76SK7b;A/&3S8cPMdg@<
MA)(4Sa4JB#TgGg=&K]EIAE3-(d9gJ\OgF]<1X<^#.09E)Ge72+L3RcLeW6gAOR5
7)2WO((]U).9CP^.L=SOaXa=.^WG;a>aM3JA7NA/=/M@N=?Yc)GU];<,]]/UKQfC
H+J]ae1@P25K6G10N.c?KWW-3D6@>M6XON+Y68AHKB+P&U19\ICE/^09Hc&[;[.G
\E3DCbDea#HPXT4B?QMAY2:MQ,bQE=^92@BY6+2E6FODYDI[6HPH<IIN)R?4L/1\
g^Gba\]:<]]XZdUcLEQP/6BQN_f=AaY[U1QZGd+eQaJ11>_bNgBHZGC-6G3A7a3O
LT#5[=/86NLPI=\Pd;PXd9LHcPOb2ZC6J_<0R48N91;[THK\PdTEGVgCYY8WJK63
=/E?1e5-b-P9ZNX;5T]cZ(UTFVWPa[K_1\KdUOfdUbM:b]]T(#f0M_8186S\;B<[
-EK5_TaNO7@N7TB4eaNB;HFUg(LZ]6@IS+B9Tg@dV]fKD9Ng-?bUZ2ed><R7:#De
7L(/C/T,1+bJH&I&I1GRbQQA4(@S,dQe.>Q(8@J(GDHZ:]=/XK12dfdWMKfN2M8=
dOQCAY4Xb.D9V3IU__Cdf65)I;=f0G4Y8V#gUd^\gfH@P4LW>c7EA[0VA]OP[+WG
DDX>@ef,GF3gf>a@D;3N&]X+I4-<R=N0VUG&O;:7f/\)Pbf5JEaY^)D+JQ@6ZFH=
:PQYR@AGN_.NJ?1-S[)40/e5_\<E9,[;?FcV2.?@F9,YZQ4\#D@)4J^f#c+:NV32
cd^XYJEcYTO3APeW,?YJG80e]JKTaF8Y/+I=>-g8AO<]^EN8_dc(_YB.421F2ES]
ccC)?bZR.P(I]D<d7U(83UZ=#ME&@50Z=V;I:]A(3B2=^=C8]CHGa?)68F9DOX)9
bI-==0JbS\CRZI6LWTA0HYD4GCT8W<B,bf@M-1Y>4I.adg+H_#=^:SMRUC;086GO
.,<Q@_4;,<YW,,:VU5-ABPe^-(Ia[1I\27Yc]K/5F]a3bA(HSC;,^ZA7V5_LPKKQ
3GON,fOI#:bJL&=AWfWJ^9VIM]_3&^2=3X+g382GTfQ,.::9CSe.:RZZ]bYfNLYL
F2bba9/PMR)W3TbAS]S?Q:P3.^7[D]d,YGa(Z.DCPNLE)c+5gI:./U)cBNJFBc]0
f2/,aD8^P_@__()U,Y5-3F=-3:3^@ZDI5ePebG-#HcKK>UFDgTDRT7R1YNSg;df(
E7YegG=2^WG,8fa<^0f&-VDS@FH+(PZ80#Jea#([#5[^\ERVa0IV3;WYA\KSe7?T
1SOC?0?YU1._(JD\)2[;Fb+ab9_4KA((14S;,>]E?>\9D,VF(aB4917C4V<fS@.H
8<863[e_WZ:1IR)GL@X/OTF>NBdC_W=dg;BEW:U;TGd2^Q^1;+L(HP8L]X.dN=DG
+E_Wd2Y6C7H)R897,)(<f)&QTENd:f7-]^OfBP3U61MNgC_?E6BN[.]3YY],Z)HU
]5&__M20BG)B\8++cX@2X(-E9<L5-+CTEGL=Ha6@6DTSIS\L/\]WB#gG2eSR2BL#
6HOV@.-NKNY;&Y:RY2+I)2[04d&bZPE=?aI75.<-Z7=VBRJ[NB^NVQ.A0:N=K556
<J9DaVYLS[3:[,:<TPgMSOU=#>C\B(,R+6E+DB70:JAO_Q&#-IaX6?dXS.cOUSLK
QUNB+PA^PCI]X4EXLKc>FNT<4F-]^#IWWaV6U>,E999XgVUg@@f[Jee(QcI:1_QH
b=4)KR<J#);USB=agG&.ebTY@a.@VA=&09WCdcM/1?A^c#<Q;1VA^bA]<bG2Y=b:
W[;TFWbT,AD7f\8#/.@^N8]R+EEcUZ9^+U:/>e\?34X26Y]?/XV-:H\[K:]a7eXZ
W@E0BOZE@C49(;DV(eIG]]\gL/,BGNK,0L^c&1NXY_aN4[11b&Ke;#1aM71f^B<I
fTf@d;M=7]LGPYbG>c/ZG11X#^VT-,:eY[GNEY<gR1:-A(32_DbJ<deS/SPfcVN.
5>TU4DM8V8-V16TUb3@c?gTbd/MF)6K0//K+:C4F\G./[G@gTDNa?Q2<#K;:dS2f
Q9b3+bgfEe_T6RU+eL^Y,-TKLE,71LY:M+#7.2=&@SO>K^YS5:N8^WbKK1d[Fg+Z
)bGH_><58A3XM-eE.W2)[-I/U(;>\N@(Gb)ZY5@Ve)0d3/_)VH37OM7)X6?@K@=Q
Y0.?cOX/OPMTffO(U>ZDP_,H1Q@5fb6_b]/aK<bUeIG0PL3a1aY;F#Z=bT\J5--a
c^5Y;@BBXQEX/1#bRfC-5B;_7LCZ;C(fOJ;0_Pe&.4&Y#gK\-SMR_OTfX[^EPXHY
C-URc::[O936[dSSe_^1X))L+_Z+N]/>@^[B/E#L9342<-\(>XaW/KJ)][&9caAQ
gOdL[0M#\(:]_KG/#M>+0N_[d-]B7#gf1U2.9LdbH8.dC7:V\a9J+?]FX0Q,43.C
b;8d>ZO]1ETL=QPbZd(<I86OR#GeGF:GCKW.b4RI_DM4T>CCQ6K3SBQ\a@QbKI#_
N2dXH>V,PXeTI:L]BU4LSF3MV.Z<EMP)(?CPUfJN0KESd1B)8>X_NI.-Cg^?6)]D
(Wg5^ZgbC=3/B&B2<EZGYGUST\2C).DB;^gF26)dcTY#U[B9;?T#@VR8SP:<C1,K
VZ>OE#DPYZXDG-W,_\XfQ0Gd9-RIJ6d@JGfLD?VII.2:ES](T?0AV#M\+:A4TgbQ
,C<_H+0Zb^EXYE(&Y:;JV]CMEG8gXdEZIQ:Fa77@@I4SP0>N,a;#VUCZA^RUOWYB
\)ERRA1H5a]UKTO0,K=>:P@?H[YZDbgVAS7K81<O?[&Y\R^8I8QdR+67Va/L90))
d@9E,QfU?f14cRF3N2J6[DdG1XQRbQ.<1aE+#R6g^5&e6;c(CB(HT/JM+]7=6D^F
dHIRL&&RXAQLIcTO\/\@E]e8J-c1O73-8G+=f9XAfaVCU+H0&/Q+=J3+EU\H#RKf
,;d5W/0_Ne48IaK,[J2A.:0;BK8[:(_/KIReT_QF;FGMb+EAB0IT_/21e(0-I.UJ
CLCHWbXf:6?8U6_FC8HWFOEe)9N64f+W&a?Uf\?Ee4gFZD]Z-P4^8.KXBD-SWU/g
f2:K/MH+D+c)RfHNU:S2dV]AKN^22LK[&G93N(<=_)cN2S7&b7]]6T<6g[P22bP&
#XYaET+L?)eFeUcI0)FNc3A?,UDW7Y1A4cY\#eU5+#O76_HWQND9)aD71bPCHYCG
+4VRfO;UEPTgU,,b=Y8Q#(C,L4Xf>e-3AY;.C.4>9WH0@=P#A8[0M5H>#bRS2_L/
)Ma5B\<<(L(AfC^@DM9[f^@a2&U8K)gA366(c\fdUSd-N8;@^L(cHRGd>NNgB6J/
@ILa<):T>RXY-ULIdfFB??;[;N[O74d8KYC8T3PQ(dS&I=\QC0fT;;gQ+BH8(Z_N
VRJSK9YEg24&\Ob-R[H@T/O3+5YPB&Og?;6L]XBA6WB4B=@/;3C4)=;e9b26]+e2
PcPEJ@27Vc2,XU@8Cf+U=cJJBYff0gQQULeJY1gaSJ0+;Zc#fS#X0)[T2H[B\079
76?#+H=R4?78G\;)((D]/JHRfK[M)M7&g9AF(0\68X)a>4.-O([_BCDU^XbK.9R=
TZXAQ))O>d:c4891#N<YD<^=M&APL0;QCXE6a-GOT,HV1a_F<-R=&a4,gZX]bLKB
#Z#SKcVT>d<9VCeX>4./a_U8_30L:^RNKQ,-BCUg,_Z]4#X8eVW8E-2&_T\&O)2Y
>5)LEX,5B)BI028JVO(6+A7NU(baU>]6+IaEHB)C9Ia0WPf7.Z8)OQ5>WL8N[D\@
[J^+fU5KGFOCGeX>?U3a.7A=bUd^D(LDDD;,KBK8\f?[?8bP25.Gg2:L?8S>8=92
BcN\E..YTdS(a6J=e-C+.(JB<6M-e^\><E)TL3RAROSD<aE+M5eMbVMbg3))H&/U
SbgHU_?Nb)+TMMeY,4+U#:7V9K1T2@NW/G:6@c5e>P,cJf@8I\K9B03c2&SU_5ef
Y3#4dM8>+26XVXUg&@IL8:+R-6Q3]5EDB.IRTd21VOc;OCOd(/9abe_0VXd.5<CF
^7@(9Z.KONFL?OcR]CI4V4;F=>4@(A?X=9FfD86AF2XR6RZf1-WKSL//[VG()./-
M=Y/&[TT,E<O;HD]AQM[I1W@#SZK@G6)((RER/,U<Bg,+YW4<4Q@X\06Wf&XSBaC
&>bO#e_[U24U?5JFLH6_BQFWE\3aOZ94LI[<8XV2?)#E:UR^B]P#_7D[.ADL_0.R
AS9/TS19M-N^]@QG6A1fa.dbd3V&:e[-c8+:@J.]Y&>Bb>bf0YFP&WD,D2gTP0ML
61N0B&bJ;:;_F3FEbFV\-V/P@FSREf+>+g7K@#;CCL7:P_@fWdW#ZNW+0/9[1,R+
/Rf=/1c;c\[2>Y=464.?Y)@gAMK3A>,,4ABe5(GS[R2f>C.,<>GAWZ)eP6SZgb0b
C(QJ>9&?1_.MCY5)O__Y,+<dAJ3Jf5X/(UeWfU0R>]]g5^ILUNHDJVI2P3H&g0F8
/b[P-.L]a/a@5Z-3@I_A/(g/F.7[(6K](IaFY..DS6/>1&D+K&0QB9VAO_TX8=9#
FJ6@W6.8dKFXBST^];O-UX;T[(CX>FDD6&[/OHRc)/8]A=)G:0_WS<E6IG]?]f)Y
0;SX(>Q,K1Y/[JdBN3^]#L,+-PRQd0Q@Zc9+Xb#4S]E1[GAeFa5XOBeZgY0:Ha9S
MQ-:S?&&LK6e0Ie=G_)gO^g(74#10,bWZ)^,Y01#/VQ@E^)=:<Lb,;LBW>P:4:<R
N7Wa#INU^6OD<G)Z:=05,<CY>D_.-cfD;M[Y2>M6X?V3Z)RQ\8E1/,>GTINELaAD
.B\\[TfbK<\3&:fAQQ[-V9V3?IC[GN[^=T?_4@>0D,DJDMcKU(dFL3>eVcS]^;5>
LSUJWDGA=bY&<X<^H:@6E#Q@KUYOaQFDD_(5e\Z1BHW)JOFE-;RdF^9Kc_-9O#9J
>)XE=:=JSB#6;L+;1FDYS[<<XdTD]9c@aSW^[\PTXG5MMFRc5,QZS=F[g18/\+cO
;4=ES(MV:6M75SVfP98dSD[:,K7JN?IF(,&.H;.cO#f(ZKDZ^TV<N@#WV.G\YFP&
<RgT^(9gIdTaO=1AAgOG12EN5(H[b^RVWLDWe)KXLe,_ER1Ngb7DZZ0]=YT;V1(>
>&9E3>-E]?;d9NNM<Z:A8AU1X\,@Pd01CbIJ2LGNO3?L<,OK.:2R^)0A.1(];_#Y
)G=/fL7Nf#3#f]TAWJ0L_ECKG03:D.-eDVA5>75eUSG.g_\cRV+c>13072]54a5.
AaRBO,M&0@2=X_)QaPHM1Q-6;/UeO>SX1b[6eCU^NZU)=ML(0/D/]6?ZLdBSR0#5
Q>/MQ9^b#RIA8>;Q?b:?Q/&6TH4Q;CFc;-KcURM=B0B8D(ZS^79<d#a][Zc=b<]6
dW9&;I+2DL-[FBd5e0f&d?@2<PR<_<fS2JbE4O_@K]V(ZWK0VF.W?^^\_&2[,IKA
6Ec_^1SI],>HUZe1/QSYbC@WD0,gJVU_NT>/bLKALX7&/K?+X(\/I-:BL7d=9Dc?
<W<bE-BaW&b:(P7BH4D0O#>7TS^gZ.fb08c?ORF&4fC#JLE>4VQLd8S+&C]^:H/<
_3J]I7]0],X=d?DC\/BWSFAB^<eaP9eC;&>dVg0HKaa@O<IVYcCcT94;@W>2S<K=
<VeE<9ZJg;(A^84+:L6,LPd0^FIUPG<S&.;Z7?.W3?g28Q<O9AG7NDS5S54#IO3?
VNTMcPDTD?_3>[]XJSgS]+2d#?XdZWgdb33=<eD.Q3+\#E3:_^L[8e+^:dPOg+]a
_1@<,MOgDU0Z,/=Q.+G]fa&<]L_dcGAH?PLI_IO?S,6ED,cGa;dC)gcNe1D))AaP
Z[gG1?]=9RD^MgB#&;_<E=<&9\,O/C>T_#VTDYJNLYFB@Jd74#ST09H,9<J;GS.P
V#R6N2eRQCV,RAZ^7Y)/8\RfQJU#>E2(P]gU9VY]+-VT_=O=+#=5(IQIc2dAf&_X
+S7:NbF:bfA0DSg&daVR]L&LNF2),/0g(X>bV1_gaXZTVYO)MJ>fe>WbIYg+eXa0
9JVH,UOf\YR:E8^Za-de\1#&2g?dRNN#-<)A2@.ACcLHRX67[TKVf9>)^8)XWDUR
Y28-.&g+S.1V88+L(9U6U<.WW=Pb@g;PDZ^Rf7.XMONdMF=JXSLH_Q)7:U7\KG./
?Z2a)Q6JE,Uac.I^8Seg>=cY>BT9S?ZL1\bgaE_IEEL<;BW&H\18-_Ub@#(cZ;;b
F]ec7FWVa_7c.(#ULf3Xa-G.+F9_N_[OH&:C9Z[=#VT66:^U5+NME\K0\QSHecL#
MA9E3Rg5,;cM_81H/,;aSDJX4U.,IEdMT\CD258NbKdLZP+H3#UWa)=gF:J?UT&e
#JD)Be.\4H;VDd-bd6),)/V,0F<[7e/FQL-3T6NB5R2IVG&?2S0c2N476H#+(K6f
T#3,G(@Y2CALW(/aREF?FF8WOI>QMYaZH@+8=H4&K3/,TbLPSf]EJ:d3<_Og73BO
E8)[)5N:)EKCI?1),G?e0Q\#a^7V,/(^50W^a6TC1T1K9CB6^4B56AFA?Y;&Fgeg
HCaXK8O?\6bc-K^1XbUKJ(ZLB/7eVUJV@Q;Hb0<#>^GbaG@Z&HHH@GINTV[/b4BV
U9J(RR4;@Q3-ZC[U4a#9/0[G3AQ(JGbH9/C8S+YYO>TT;f6E;;Bg4@>LI->6I0RR
[H;Gd?F&H71d1?[BTDL@9UcYUY(/FSFdA5c@[H<C[6[-;SRH).1Y;6N-ZA)b+@a4
T5#B,@EJ4(?bc?,;9APC3GAJ6gU3.)f1R7]MOSHg9UYEE_.B?7g5?.,\ee4FY/N5
=b_8\F2,P9S<,[?(dGIX@KOLB&c0c(Qa2_F8DTGHLSE]^5<DKcXeK;WIMdJ\M;D1
b,?Bf=>,]IYZ8R,Fcf@/X4SX[O^:+3L#WR&_HL+W4g)_,?H#FZb4Fa#A<4TFGNB.
_fVVA0(W_GGd</4]W^Q5=[(eZ#K0DTFJgYaRNEA.&=2.6BGYSO2DS?f@D2/X#(?A
Yd/DZEBQB5J#EH]H=.JgZQcMd.cC-:8PIXZP\39PNTeA@,.7&<WdCCKXG6WZ9NMW
WB5AW\>daLU<0F9ab_J3UEC\-0:,L?,J#6\)d?9=g<XI/M_A(#/SA;#C);c<ZTgY
0=;S[)GY]D7SLa2BWfEXOU\;.M;.=-T5::f#[c;:3ZAHZT57be&@LWAKZe8gEbI+
#2^I1ST[/ZITJU)adc&Mf@X+^D=U=>f4EHRR<HacH+Y<R]R\MW@I7DZ26_)6A9,>
R^FYY(E/eaD3(9&=<>T\MH>d2c5\3HbE_=NX,9L4OWQ\W\J4Z-+T(F.PGe1SKd@B
cI9@?=A@<;X#\&c,T@X\[<R=@1S/Y.)]U3QGY>)8..A&)HU2R66I/D(8.RWHY8GY
@X-6CALg2&AgQ^RRH&M(bH.>a4<]2I[]Qa7LeU89.#;[K+]33VQ@3]/D)IJ[4KE@
040@0,Z:3FEIa#<=#5VI=9e,+XePJC-4WgGG8Sa(=<8]-20X].c\(XS1,C:B=YK]
N0B9):KdFc>7fcagZbX6)QVMeg8/=IS_9Z2,b]SLT\0]:+L6TLG98KYbM,I=Z/c_
a9:SC.5/2XGB)O=d,7B6BIX/g^.5)1M\5=ZPSM.5,&S46DH;8QcWM:E(^@F.#D/T
<)8:.[_gMSRD@Q0RDFdI6C(1+B.O3a4:OgY)A2ffJZRfTb@>3Z^G;2O<H&g:L,0[
E&S,[2#LYEP05GWbDeNgg,E,D?O;G6/K+SAg,eO<5AP:=a5(#@V[<)@+.2\MdL]R
.&G:UL_\SIJ4MNFZF8b_H<)(N?^a;>e]P/<Sb(S]4fRIbBH3EYb7GFeZE,b0cg/4
N<dI/>MW/b>QdP5b=,;dK2H72Z=ISeXP2S&RKDCe_81],3OE.@2;;JSO#EFe,##)
^\?]L[<)IbU.6H0KHTL>.M0=Of4?_c\6^J2)R/Z3;Ud0BAJ+57d3TL/_B)?2+6+I
D)50&G_Y.C?gWfN>^c9BS#H:FE+GUb9S:H:688\CeETdGZFYZU8&AM&+;0@&&37G
4WKLBWJC3ZI)4?OF4R6^P?3?RCPFEaV-&8fObIK8WO\&R7>#dd<Q(#+N;HfY,02I
E3I5;51JI1g^IdO6=>_K/I4Z<T).)CYaa+J0V8P6:>=LO:d)JO6Xa](+))290LY]
Q59J?cKJK@?H-^])(Ae(BVOZfO>&H):;4bQ.Y]8+6>c&8XCd4DQ1;34SeZL2.2G.
Ig&b]+;=>b?U3d2-J&+aZPeI\,6]GY^+)[(\/]4Z^H+)#5-;K=4?>OA3[-\\=+)g
\8F\=-S83gWZA8?1cWE/Y:TJ>M?PbB83WR^4a\HA0BVcK;=B^8(87DNO]]D1.bd4
G\,[3RUYK3L]dXP.4Ta&&86)&[G&7I)N5KQO0&fPDg0UCQ3dC?^X&f(3RHb68R#4
-?_B5FGgQ1FG.I.D#[=cN(R@ECPF/-e<EZe01;ZMDC8=RNI6?2-+)\VRN2]+EH3F
g4\F)<7QUNNe;3T-3d24SB@+..3II+K3652G]<.f>F>RV:B@QgGQ2c-TGHY9F&\d
JW]7OdR])Y5L3ST(I#LM>2/W-/&WLZJK[7.Td=@Y/?W&c)ZA<-_R4+3:LB=^A52f
B(]@5]#-5=^=G;dE^]B4#MLR&GBU_4N7Mb5-5&]@9DWOED/HAY7.Td:GC<.9e=D+
N1;c#;fbS>,W_ZZX=)K^[R/C4E+M\P<C\<e,dM31UBM@IJc.e(J((]1:_/QM02[\
2J7FVa]^1]_f\f]Z4Ga9U44RTANVeP-1F3;KRMBb6f<ES3]:G#]&P@K)G/@X[XR?
EN<bKJ=U=)L]4H>5YGMXY,P[,[DfBbB-F4KY&fM7O8&D&C4H_YQ6gc-J)8W]Y3DH
@0;<#)a+bFT\KE)a+=O&<]Z6eG?FgH:Z_;,WW:6#FR9\8E1X:C9;7D(P/E6/1:-7
+PZP:(W&G(X2-9g[EM05X[OXHJKW(R#?<K2J:JHOMa0+De0D9(#@2,5.C5W:_7S<
_3Yg^d:7?37Q;@S@\@a?9_dK7d=WKZ4X@6De^=+P+XZ]b@2-KQNV+YVBe?;4Q^ea
N6(-16NC[aIa_A:<abV7\7)3SUBU:32C1\cWdWbQWD2eB@<P2fW<;S@F[I&VDWfS
DcE<Rc#J/XPe;fe^B^V7LHD>5(5R-BODX;YN:LW]RY89e@X_+4?IEJ0Z:T[H4+B7
0bDTfKVU5RC(1\RWKRSMF2E]NUV\6b4WJB2/</XA6b7N4&Y4g6OcET?a;>cY1VYO
?f,J)CIa;JY?0B12f/D?^E.eA3472^Zdb>,ZO&,g(;:(EFZ:6RAc_)HCXT._B]2J
MD513CJ=M&=[aAbV#eU?<fR69N\BNQ0.b(G2>W,c[C01PXDCAfJHZM-f9,G2_.Yb
:32a]a)T;7EGI&SBF5EC0DD2W>)O.IJZY26DgFf-\6J,F:O<_gJS(\V94C=HPVCO
(PT]W>d+RCbX@9U7TUDU]AZR+8=]<G+TMD69DLY#BZ\HXS@[GV8GT<YEVacD:FM)
UZ[@GHf<\Y9T;7IQ@Z5VIP;7^N0#8d+\)Z6f@M0(<\ECL=6M=?H]0c0K]fO/9IP)
-[];gcL?b7e&<.1P,YGBOT,N7UUaH7eWRTf.:VNYY24Bc+<EWYMWGTGD<I+5g_(D
Af+7A;505]bL_+RZ([B@N0U^TT7P#2Y/NcU-D]84FaC&XI60<;C/4PSXOWQS#?C(
1E>>CTa\K55f+Ca+\811eWHX@G;F6-f@RI9fZ,BT<,W3g^MKg+#ca0@>4;>JL62R
Y7a4/1[#X1G)S6^;BV\WL-&H<G13&BIf:<?6NPfd^CWB^LZdVa0L>40e\Z9CH<3d
4SIgE[G42<>bH1H)\K?PY[@(H,TOK9A&A9GV5#S4MIc/-?E5WONa\49IT1RN_&U+
=UUAPbVLdP71c>\;U3_M+HP>MKL(69?A:@WK677MD.EBI;>A<G/7Q@.B,Yf>>HK^
WGZ7I;#^,D]b9aC;W2XfN-3>ceVcI5YZH<1\UgMK<EI?Jg\^^]HQ(_J((/7B&HLP
Y>J;I<^DH/&_gI#e]+Q^,&WZ-#cPC=-C4a.UI0a.DTdD1-b>d3\+6cO6)H5Q<@(B
41V2YY3aP:M@?d\d+MV[[?5S:LI7bVe<Fe^bW,/;)ffg>bN2TU4&a3>5#A12<Ac1
QX/g+@AHKPF7_IM06Td5D-AZ\/9&DD^JP\,,K0eVXGXL8HSQ+@IJ:?;5:Q@@D/3=
GQ:^OW(W6)ARJ)Vb6[[\8&M.9ST6&Pe7Fb:C^3QRSbC,Qc(@_PJaZgeF.UP,^XEd
5C2Y7d#6?FbfWa5&SfE]<2#NXReKf\12Tcf-]UK^.PZ<-:P^dUL_d+GMbTE5KMA2
&0H@1XQ25CdB;E(-Y]FUEJ0LQU<1H8-/.V&XEeRN9#Y1C(dGaQ:Q;@K5=c[V\I73
\X2<R<GV7cKI.4,Ig4S3bK9^@Z4NgDQD6FB8?;.6NfS?STIK3YTf\D]K8^e^?J/@
;\g-@/J93XdE;R/],aPeXbERL5DBJVVB<ZS97)_LAZ,I>_3YNa6(^AR4d=ZKLC=a
NZ&P]Pf^aU=0]N;(^41<W.HGF,OT4?]<QG8(Q9>]3VEX+3a(R5+^AfVeeLH/)AV2
_?e]ePVZ87.=e]=(?&AP01KMg]IN8\6bL#deJI>;cfXPKb3&^&X\7GZ4DPBgf05g
a7W8)+OE=Id1:E&SKH)]OG@+?^1:bUC;Q]S^Kaa=9Zc3A_CTDB6#[Q>;+DDP\b[^
=NP^4bP1aagdS/)Rcb-CPSD.cZY4;.^;KL5gfS3A?[a?P(__Q=TVTT/JZ<0\SCAU
Q;Qd]1A]3MF/O8D/U_/1RMP:VfHS+b&W:3a=15&/fRQ+eN:TNgSY82Ge7g>71YGW
5(6N?J@8GGcR]#AdB3_XUA\=_C#=b<8)<+V#5H(:bG54(INR0gd\<1BMU\G6&MJa
GA>]O\N:ZEC0K5)NV5@E>Q9268eH9H@6)>PCZ)>>]QQ,B-]KK:<(,Sbf&4S7N=;3
+53(/X&U(AY9&5\b7B;M7I4VFK[^g]a>JN9FYDdC2KEe-\6=/T.TWS_<af8Y)D.B
947I1R+,IYc#;ZLf[\(:,GD)+0HRV;1&R6855:SOZ4\&EG;-[E_J9^S,AJ;A/GT7
a)[5F-9\bB[2Z533e2V.+2WVX9&X4TUed^L1S-CXT8+eBQa>RdCT#KV#MK#dEAJD
+Z/QY^J\HK/#+O#c_6H,#7Ob3;RGLe/X\)-1SC57BPZQa/M?+:Eb:8]KB#+N;3,S
&(^:-))DNXO;U-d6H0+f,.2(23A9g55;U5Bf5Vc,-_BL-;H-KORKM)ALH+eb(55Z
cQd?/L5;?#(]L=9c?8V&)7g[g-?dZQQ<PD<BA@PS2O_SS\Z1.@g2>.#_BNbQVgFN
>)/K+FBd317KQBR_3=F8;dLaH]b>8cO1?TM25a-T3?4QLJ5I>R3g>>XHC;UH2T(/
DOfN/\4Tb8a_UD>X1)K,7C);Gg5#S9C^7_gPLH:,TbS-S>UV->NONN+9#J(LIB5d
df>-LT/Pf(QD0KF7XQ050Kc?WL_:3R\][e[fT.K2AbeL#SaV4QN<3,IdR:eY)PS5
KAKB_X9T[]RVKD<LRGN)P^cA1RZ=1B?5NZY0(>eaVT_XX>>cg(P5\N[+Z3.VcD03
7\NL[>=b>gC3;H[_Ma.P6E5QK?LFOPK,3R4^28:-VM-)N0ACR.F#d72a;AVdJb&4
]V&g4aY=4+,RY:+;9/g^6_&@d80Wd^:,8./;8R9/<6gG0fHU62#3(9I;]OHfPe4,
=C:/OFSNgX?2TeNXN?NYTP;_c68WYUM#V[Bd5;]]AFMI&&fG\3U@3DWCdY#DON75
e^O?00J5F_H5H5\_Q?P\0J[cZ@BbH=E,.)UF?NH3>RW.gfS^4.O4WN9QY2MeR70Q
F>c4BD<c[(FMS&0O@8Y[dV[3#ObIdGAA^ge]^Q]B=\ZPQ#:gVI-B]CR76=XU+U4R
QB);7<;\-g,+AGGD89d):aO0(DBCS[_S:Q<SK;Q9[84WJe0Qbb0[b<P-1DS2?K7\
:QLc4Tf6ebAL+Q/<5&W#^B,[((H]@#Z:OcUGBC?^-5R(cd,:<_=P8]4214UIYUC(
W2484+b_.&V,H7).@dIRTd(ca&L.OFa=Rf<bK?1(g0a?42_&_1F/31R(])gVQL6Y
>,Ma;?bP)dKMLgZI_ePYN;LSeE0K9OFKVB<]DAMH+W1:W+]1_bDF5/bRc=RZ5Ydf
;#VB&]IT\@?H[,d/23^-Md6TEQU)D^CTPKK1^,;.0HY+=fUA/c@[>@?,AaT:[[:1
N;]E\V\7(K;/7,/#^b.N/1V\.6KP,9<f6<+SbIH7gY^S>LOGR_I)Q#cPWRaJfXNZ
1M@d[DH[?M:JV=^]4K/a-#AMLEVcXO20+L#+>0;@+8Y[dN#Ie7]/9GPV:H^JBLC#
T<EG)TA-(TQYa]=&/Ee=T4OALa6:L#@.P.4T2d_7JWLA77+YO5]?aSg1@Y#E9SJ.
;;gH--:6/MCF1GVFA2KO-V#EO@C4WAfdEXK^)B4:DMc^UFa,;PI0<\eSJG2UBXJ+
>X=\7#__?^-:?;WFT22D]ZH#1R^6gc)L5,>WPK^#,Z+a@&^(3DXbP7C&>9S^L-LJ
L>^3<&<Q7.V:eOMIH69f)a-cC-ZL8(1>@+I]U4[@1YRcU:JID#J[N;ZgOL-+7g6K
]NZ8?BK_T6I:PW<-/)@#+ef<OWXT-G;)/_&XA;+BaCFMYW26((O@_^/Rb[?g&[XM
GPX41)=-g#;R^#B_dNKSdED_H.JfH:M@d@<UCgL@(,aCbF--A(SJ&B@ae[Se0BP9
5<;1V-;AA@[ZT-Cd5)/-1=NKZdfV[5Fc<?&\T]BQQA1a9QAbI=b:TFTTP>+V=>:Y
_BNbMg_9ME.[G//Ng?@09Ib:J7DQI][#LD_]/TF;0KR7_B39I2SNK]MOWd1Q^fW\
8@.B(\G82XAg(?30;g_/V2ZUP4,=K-WI1C<)K6OL@E2C=Q[.bZJ\;[0;U5X(f&/X
GS>ZT#&;Kg@S&&(<S@7C7\65d)+d6MKObF\WEU-?H8:M8CZ?O^GGRUa\<>;,,T/b
,-eUUU)SB>SW/F2JF?+U10Z);Zf;,Q7M8YAaT+5=2&U42:V;Tg^;0PFG-+5?c[80
#C.-F_I?,PVXcQ_.bW7K<2Y<+_4HaeSadaA#.UW@6P)^7Ncd_8\/b8,a;?YB5?,.
N+9E)9PY)X=;H2VV/A^&URK>US(d_)F28(G61@b[Ac>ZAa\dTO4,\_L?O?\C4.KG
2Z0&G6=W[+#cAJ1L8HeS;E&NHNWR;54#1;edPPe7>84@&bOV_#S]bQ(e<26g.D^-
SS?Of0cX:+&aKg_SE]A_fO6//gZe56597PI14W0dVD^-[J.EM5((F>N([#VHI+#U
CB+.1QI43gHcaC79D4\Z#NdMbRF]bXTR[0@-24_0<>:SR.,-_F]R)6,50>C_E[=G
?f53NOMEIbC+5cE]Uda<geW&O[ZNUE_Z2c,Ob&<.60Ff2=F[TM^+;78&QK40=?_T
JII2Og6^\\YZ:O&Wa22VG2YADPe+d(7KW9eULENO=8f.<FW\/0ed:4_E1U,AC]0+
.06BXf5V0N^QR5X?8Cd,bRbd&A+.H=H9VWf[0c/M#OWN5Te;Z/6#Z)f<CeB87+/:
5C@AbgC+cX(Y95;;)XOOO.>XNSQeeRVQ4Z78F@AT]3ceLH[0@g,#<VH^dUEdJ+Z>
KZ@>G316fOa3_QQ7BB=>J4<5]];-9e]W-fZJ8<:OY6L:?PINDBa<(NBY]d5UIEOB
d#KgO5TDaD@2]JSI9WXa?cdEV;N)9/ZYUa;<0b/g_P8Se\(X5I[5GJ?>9S^AU13K
Y@4VI6:Y8aB2.-WXRXRCRCN^.6=1M;6;[3P]9HWGR@:NVUEN(]5X>P]7e<beId5E
KNG<RX-@QIXdRX?R;XF_9],P>.,Q;ZVNJP3]J1TJ5F@3fIC-D]LV:8L;UD8-eZB3
@IUJFS&FBc1Wf/K&E2P?4HH4:]_>cC9GS<>#2gNM:#=UAN\#=]D1G]RJ[K&8S9K5
UH(Z10\^T@2+aM=+9ZY45L5g=S2[7LEY&^Ua(+_KIF<#Q^O/8/gE]gaPF(S:QW,F
#^bI+[)Lg(-_:1#+>>aI@UUX&O\DD)=3GR[?Y74()MW2V@gC_S^RQN7Dbf0RW0bL
dY<P+Y0^P;<?\(J,_8IW/PK_\9OX4@0?F7/Q=3g:6YMR@]AETY07Z1B^dU<WI1Jb
f@3aA-=)NE(O/4NP.[4JbLL:8<Z4OZOO@T=:OR@WR5?=d54DD9N_B-?f,3,?EL:&
\c4JG\T9Q&]];:TPY?EWCbN<B:>,N,\U&-fgOMacc-c\]<DFYWG(AeKK5c5VUZB/
8WHF7Rd\>1RX]Y[)f+W.A/N.Q>8WR0QKA=&d,.UU)R0@QQEbUe^+MaP].DGA<66b
,f[12WKJ]T(&KWd-J]4Y,HcR2<NHJP_,Z;R.-=g42)g_?U_999OMB3.?MQEPQCX0
]-LSQW\+UQ;61MX01],Q07:K?JLHJWO;c84/Zc2eAZ5ba2c;7T=fM+C+:Q[<f+,/
<6B@677G_C8cJ<1:7,g:4;AePJL]NCSCS-=TERQU<NO+1X&4@@0F^1+_OB]F?E\.
g(@#JA^EPRB^De_B-g(>6Y5,)6O8Q_DK2F>agbE9,g)48T/abd?OWA-,Q(=,bSGb
^@_Q2O2\@&dMXK>_EOUT7Ge&4M,E3_ETENBgg=8^b-2aE=X]F)S86MY>AU-;R8N;
J+AB(>\(KHBXbaEU=MXbP>>1]5+R(F/,LD(]eLOP:ZWBe]N9Xf=9c3STf5]I..]1
@?P/8DF1S1c<]P,AKR7^U22-UU32]?a1#2eHMNUW=IIXLQP8@99B+R>U[Y.PTN,\
X@6)N8b[X?N[I?[1\b;DBY,Yf?3/2=@JA.]OKXAD\a6O3&&8Vc[>(6E^d_\W/K#-
,Be1\E28]/^&TEaL\+[3\L6B_EST?;GYK5aC]HP7f2S5#S>:^AD&(/T>46]G[HIN
N,>Jeg-?W\-dY<PJHLK(:M4gf_]VBO8PDHReb2->?AdU=PWJ-\@:[61.59>+;aUS
e5D-f5O-:0=,gK@O3S)_K_&>4RABQ_A08N4Y)3J->F349U:[U6?+a-AZ&Q6Sc3W3
(V5R=F10/-[[\Y;+,CNQ&XDQ(_IH<J>;[W9J;+:f2).=.3#)CA+]OGW8=MF&Jc1@
1R/g;RVUc8fT@0?9cH=@70I7TY3:_bP+f^R\_@b=BQ/EGBU2.A/G##UY]ZE..Ve4
_XTJK&.TF:O)NeAf>Q[7TITL5c9(#ZT0Gg+,e<cMBLDXM;gb91Tb>4JD#cG6[R3<
<P>I4SNV##7-XMU3-G4D^gK-6+=2K:H.Td1d.[bDD2Ya&@]AZ6/Bd)L(UF>H;K/:
3XE-?8,<2?4EHd-PdbgL8M6P<gG.eSE2_09a-JB?/68GQ1(QUdV7[H(_2(La[;?;
MCD7#IZ+)_d7^^+#RS&3U]S9X@ZZB9C@K.\?@gF[P;DP2V+>.B2OTD-\(427cE75
f:XN8g:XS>1.]:-.Ea5^,aEK,Ja]NMQZ323T7LG[RHS0OU/4\cfPc+GK50TgKIR.
Zd1UI<cR?WE<25LR)W9ULeHVX=VHH_0\#YC2dA_<P),<\+9CQTUgDe#.ILZR:G/c
0HfIJ-1XgdR\71B4g:S9#SAKe7657ZZG\Mc(c]M+=B>T&LP<>b>>SJ-S47^W#6;Y
EO]0BVDKCFa61JLD7X.M@SMe7^CY^&4-YENgU0[Lc5Z8BgD<S?4SN0]T-E=3FF#/
#A+,\55_K#<OLWZQcU7T&-C[:3,1)67af/fV0+5U>_VF]HN1C(<S_cUCgW[W;AIe
4@2FY[M\@.II)/ABUR=PC/)dVT]aTSf<1V3\[G<1YK2^0D_Y>+28J85O_9#PX[C&
926X:O5+&eB6T=4..<Xd_XULF:F06XcP[#E)3Y0EIJCd0e5G00#BELW]=[(d2;cS
Ze08E/+@&cLM\T+TE/T_]RX?:G2gMI@BVLNR1]6e5H5Q2e[3&(KCY_6cD6g.YN#\
4@#b/><MJ88Vdc;SKB##ee;)E#^>eHS>f#Q_ZMP4(D@fOQb,Q@S/5H1[0(&MF^F9
Eea3@EW1I7<^.+.8DL#>E7,BD;Kg[T#?2R#-RFXe+^,2_eQdJO-AY4eAEZ6Q#?1f
][Wd4&O_#)I;4&O^:C?(T#KVZR+BHLF(;=4,UPO7+GD=;Q.JZTH25KXL6gZO0Y;]
SW-\HD_PLVgADd/\4fYNM-TP=O6/g>/FR(<D54R7BW1W/7YDfJ61fTZedUR?,]5b
22QR/GRV/ILHTg6&(EU^a#=?UAB+VLOcdWM4U;D/TF.Je>;_JLNY\68PZI2)QgMY
8M&1ZJ#0S6F5a]4SaJD0;_\e?f@7+NVFN27c,Qa#?75(LO/Ad(]DOZT0=P^:S3(:
/>3XR?@d)+EL@cJFf<<bIAe6f^;2LWFEbg?5:)@1,J<7b1YbYHM7<eALQb[Ic6X^
(\X_5@7^AG[Z?3(@::N),E7YNg#TYMXEHfK.9eUURUR]-VEdHfD33;cMB(0G5:D1
H[Yb?fR81Ge.PH]E=W0-eb//fEWSe8Ee:1JIKFDQ+e@>[gfFQdXFVc9R@OUJ>EI=
OOW5ecE=47DZP0_T=&b[9?^7<\ZR&PB.@(X,?9@:C^TKD48V#CT2VG0b:NOTaJ+,
]d2J@g9)XHdQGHMPV?O\]ePgX5&L2.YK-4ccG]S9EeJR_fGcGY,)?US./+FOS0HF
[-+OFdYPeP5E7G[-?17]Wd72FQ4OI9eWVV/cbG]d;(LW&=C8gFQb1#,Ug_M(2<#)
58ceMKFG9@@7CE#F2F:IO=NZSX?(G21,#Qa#^\6MM].0JD,JEHX1Kd->c&<_J5I<
Z)_d,C(ReL=b7\=G9]-F>YA+2Dd++9+EaI^TV<0RY\C5E9-FQ9^<d:eE_C6,BP@<
>Qbdcg&I.>MAJ+JERY/<5[D.a1(WW_:Ndb8D\?:dMGg2).@F2\4cOfEfA9XG8EN3
5RNKIX=a#\g7,TAaa1Q=]d7E9QfRHI8eES_I5#O;aUQUIb84/?(&Mb68R8DfH#J)
5NAV:ZVNW(&@^&GCS9ON>90.)c4\>GG<.EJV_D_@/.cY9AZ&FR3GM,HLD+Q2?ba]
#f:+PEVHJN1EJT0GOOO8bfSfD7fVDf>DII/.&g4<fOa?aM]6;A#:HOZPe=C5O3OM
(D>0-&F/@b96]-54XE\FBPM5a9)(0OEJ+4R3LIfSP:[B_@SWGa)Yeb,;)(F(1]f\
072d/<A-.D]UL^O-CVU=_87)0.M_[3+W_A?W,@.d+5L0E&M[T@UM(1S(d,J0ROSB
dEC^[G:VI-a\R0Q@fSM\0b>A48_XECCbT^_9Dd=5f?16Ig4:bb/]M3TT5&BQA)5#
,c6=:FD#2\fbg0)5[NI/6,/PY=;f:^U<NSBL.Z<c-g7d/>ebc.B3eGVXg+-,+<E&
YD9T^?V+cc>^QB[G_SNJLW@/:Y5=dBf>INMZP12IUZ3JP/?^NIKWYLc51M7G]S(E
FGS0M6YRUE&AeMG6X;I#7CJU?TYON>CJc:b5\fJVXN7A0YN&[Q@5Wd>EAg\B>=G=
(c2P#2M-L83g/XO=319&Y&?S8UWZ4AfHg.1B>@eARCaZegXP;INaM>0]0Je+bd:)
YFd1ZFU?.a=)@(\^[7B=H-4SfSC_#d#X)OV2#WNQcJdVJQ:9dD-#be?[T4bVN-Ge
[Y\+>B_-5J+XYK8:6ILfXN(bFgd1S0b61Uc)<DN]Ad[_.T-KUc4(B6=R:\eN)5&E
]b35OU5MPCJbKG:(X<+498_0:FDPEg/X(2S^6^c1NZ._gRf:ZG=^eL:3:EU0QM/=
4UVBK<aI3E=>L/Y+U1DQf>M3,AP2ST^-aZ:XJAA/]K42+3DIJa\ecWN<8&)IQJ_K
V&,:e,9\I6NU=DREd1I95M[cC.7_BZ+J<c;?f4,87/R#H1G?@KMeIO,a[_T[S<_R
cKg&-XJ.6=8K]aY6b^-2O6:6V5gd>/?^L&AcS3@>Oa\MQJ&EN0(1OW(c^?-GJYB5
Eg)5_B,]&RE^3?A6_d+\.F;U>C@>G72VVB--K&>+((+UIN<]]/\\C?MJF51bU=EP
a)/3]V1G;)eC.9O=BVJPTPF^J1RF9^O(/K8>.Ca4S:2QC=YIM265)/(A6RegRYgW
MdC7\IS^X;W#&+9N^JBFUSMI5)JA:::G/ZKMgNJ..S/b8T_8[</[CYe2-L;X,dQ?
CEa17]<Z+Ce?()RE:<fL<>)8AI/fE(;#;?([O5:B@,I[\f0_?V/,a9#IG3c:1V4F
E9g2SWc,A6_>_ZF2E6(\G>-6\dJM;IAdL-+f^AV&,?+O:1S.UC@>9P[?^.cU/TYg
7I^Q(PVadM01I&:-=A<fJ?e.>G8acT2P^5gD4@/-5K7;@7M^YJRUYQ#KN3T7A5bc
?^XF(M>UQ)H(=EGY\K/,:=9a7b38g;a1dS481-e74(.@WWB4XMfYS2L_(e171M9d
Ra;W@G6,#S?5RJc>I(c99_SS<KT+BX<2EfMPdH,gK9^4&QAXeL\YNX:/05VW/W+W
&M@K[&FTFN<7b]M]\7P3<Q#BN&TA+RVff]-)AJ-3C;B<I;c8P)>S7Y5IPX2O25gK
GOK@6e[9ZG,/P:0Y<(-D0]KN@>DXgWGF\_+X:]-M(^a\CR_([SI36X_]7g.KU?J:
74.<5R#6BU[K-+HT[L2^JU?SN]O#ef.D5-VCQ;ZZ4ZJ,;.)GY;O9RNVOOB]O?-+U
7fM3L^f74d9f]7O(&fG)a:=;HcA^M?9RR9cd9AC;,_,=56MTQaIM_;7/GN>_K??g
#,]&C7/QY1HU\E5BgK:3S^ZNYV,WS&:ZSM<7d9cHJGQ+3B[fQ]-NM/L0O=BJKBHE
&[9,1V0N;42G?c5HN3\8-+CVGB]/Q_]\+)Y.3]+Y7MG<H6&&+aAf484BZ:3O&4dV
_.8WJ<6d#N7?=Y=KLP/5\D968Y1BI<RJ=5\L<4I#ELO;>@HC)E2_ORYUGBTR@>Xb
R26)WcXGW.O<F-U@CLPe=dG20N/;;.+#b8@,b4P^/&8gV/&AZ[R+#)c1Ba(,ZJ,A
gcMUG-K&ef\9feG+<51GTS8QecVI<;5_6\bH1^g7d,D,K^bI:+>=K9H_aMZX+L-=
:CbKH74^OM#I?9/U?:4YJ(WH6/8;(,RG;9VbWQR^AQ=-c.EYL7Mc-,\O6NAF812:
KI+^Q&B&NMgeWbW:ZG63J)&7Y,4YJU2<Ycgf0Nb,8+W_BR]8=VHVKD^fV;IX(gB+
42M09f>D^.;J3a=#V5RMHfXE=aaWc>cZ-?,CQ^]/=ESG?M?XCWKPID2W+;YC2E&-
3fd@e,\8+?f;7g,2Lc/fBQ+I\<AQ.^G,[bPAL1@Z<P>(UTFAC-91AUWYMC?+=5?:
I\;?F^KUK>TW?N;gX:;5G7M70RNd-+PKe#L2b\I=76d#K+eI6TMWE(FT.NP_FF&>
&[:T-IC(TZ3W6[F5JT1bddN.;N@CSA9K&7X_DZFa/9<aFJ-?LeP@EJ-QVVd(V0d1
XUFI&fUZ_C@BZQN:ga@PS=g54d(PW9;D&55TMV4>QEUg1Eg#PAcb2DCX#?A[/=:A
2[=]FR+OS<X]dB-E@,#^T;4=JE>:&[fUASW4NBHa7PaYO6RFPJ(aK=;dcV5TAQ3=
P)ce<]?QJ_\X0W>4.Lf&DNA/gQP>I)a8DSLIcYE]U]f>;EZ[OTS,<:;OLG@c961f
DcZ09HAY34P>.M@29PC&O@AR/6?#3[aWc]6I7I0<L__(SVDW\D7B:Rg]YJ9LLGa7
5aK5_3>##6JA)Z4DCOaDR#(DV.?/QbOcU\5g>]CBJOS>EVIKUO3D;[]8X<4VLHF[
aG)fd8UBRYJ16798d3);)P]G05,X3U2[fC8<LPSA<)I#JW\@OO4aE_1a1L8W;TJ;
)CSBCD0N[PJD0HYVV?ZCQc0_a=XN<V,5Idc_766^N<6+O=55GeJ[_\Nd53FIGe^T
ZcbOJ]_aT(I#D<11D[+5)X(O(S::(E2R77W3D&C._ZK_-IUgXdZ=<N8A+,;V.XbW
\/cO8X@E(12D6g(dS;Q;-;AbNL:,P305FPd^b0=RD1L5C[EJUWEGF/R:ET@]PG0G
g[@_EF>Rc;89HT^MK3HJ8EVd;U(&)RI<8^gZVR49C-L-U7C9c&QeXZ-b7<WAJO[/
+P6YJVUUIN33fT1Z)c=91=A#=GBHS4UL^EP72);d)WH/]/6JXE+#N-QU[;/bKVYR
G?CcI<(>H4+eCUa<,E]K7IM0F&=\M>A-E[D^b>?KVL_#=?@PM?=GfgI51:,ZdX@-
Q+DT]7<2Q7.Y:gcPZ.56L)?6BWYU.//BOW8ET4FBJX/3-;^g@TG_2IG&T.GA^FH5
G,5&ZT,H.f_L?5IXBS/Te,_2,/;<FX=LT[fNY1RH5d#[[[Bc#\gSOXaFSNGWS:UY
J0Q@)E#NPA:WSg\Z7YT:ScbKRRIPKN[NaY&P_&1)K)IPVP_0SV8J4(PgGdL1TW;G
4<CG1Q?/Jc\FE4?[R5L&=&-cHc9aVY^F:C11^]JI4HUW_FW+O/UeN.cbgYQ##+gI
H<>)d7@\WA=4c2DJ<=+Q-/K-aFIS_dSLN@g>Se/c3PJ5E-LEWdbFJ^bETAGJSJ3D
,.PBWg:CTa^M&QQ,e-XX))O4FHF3)G6VGNB9gA.@8/6PA>)^-B,..=@&g1U[;RAI
_:PM#+a3c7Z=08]TE(gWF&&K1ON129d:3YPL:f4]gDR=_2[6KTUL)CdM[9^a1gCV
@SYfcO@4Rd9S4J^fQK8L7C7,==M-S5A7M:M3R@W>gE<?HZDZaRM904gX&TWOQ59Q
+g_?ZAc#e\Z:aFX2RY^PN/E>P-BXDHPY>V)e^^L]Ce&Z^V+\S,2SeQUaU^-O,bW,
&)G)dMd=UFXVfT:[2NUGQ@Va#LP@U]HZg.4D+=BV6<gA3.P_8#[4;B4OIdefIE<>
cGG6V15;UB:9.a?.-b=[@DY_[bg+6N\GQSJNA_VFW.HaXZKV;ODW/0D_@fG::LJ/
+PKTO7XK&853JO3CW;3[7485f]0N9^/W068QI2?0YI<f2V\&1_;[fgUBb=XQ_1N>
WTI6B:MfRgS)4eA.VV0e=C64H>VLJV#AR#?P6Wf#1VeZFag1T(N>[T_RHeGZ0O4C
TF[WC[1<dC78M/D=aAOdGGSf0N2\BQg<)W>abdf28J@=?VGHXIa[Db7>VIH/A&O9
=F@FK7f84A?Y+COXMcR9Hdg5]XQEg[Z()4SBGdP,,,UED)++<BM?^+NT[8^TVKH)
H,+U6b_2-5Cg-_D&MH&O#2_&=c5E:OB[T@D2J2#CQ][7,,<ZNWJQ(.1&]\V:/+F5
RL9LJ<+0J@C@;a5S4H,LLEGcg]G,_W#eaQ85C71RPBE3Q]S#W<5O;BR#[N0TD;-9
RR)HM;X,V(AL?]6]CP?=8Hb7VN0@>f6+2>7C1RM2[1<^##EWY6.+C(1:OTO:I49A
D6_]UW=^bJON\1M_aD0-D]IAeM-Jc\@/c0I4\:,+O&S1(^ZFOa^KF5E4[S9#B+=Y
9L7/TU0)dX(\T.-Q/MO[c]NO+)b@8WXU18=6EH]M/3D0MVbG>\Z4f[M_-7gQS<D;
Xf&R5W2/)\]66T#T?>>W.aL(Zf9,cGQ<U/@Y8.==?V^BS?>/&<BaBY^(/c2//a46
aV+)/c_V2f#-J(UdAd_T\+?HB60XcF(,8Yf6_gEg[W+TWS?O.JY]Gcd,T:]d:^]>
@)>5^(9EN^K-22F)P>ad0AcaZ[6)F[HSEcf[bU_Z21Z&JWMbTagINA;:X.85D):-
gFDM;E4/L7(3S_.+fJX9?19S2X]WSd5^UHCEY8PfFD^&0VGdKSB38[c2UY&U6FXG
8G5@(CQcQ@[IN63?EI8?4W?XON4IWEb^7AfIM7c;SN?)c)/AZVfPM@2<)1\HNFg:
M-F3)]>T3Ng7F_1K]A=QW<1X_Geg=adZ4J3QURS1B4]L4PV<Y5IZba#)Z#9W8+ae
9;Q<L5X,,7=9]ORe(,W\=_9W=M70+A@Ic[[;X1YbDX:)SR3gEE1X;SSF>BK9&[2Y
FCeZe8d[A3Z1;M(C#I,7++@a<DKHJ>d,5Ta4C-<>#0WL>.bg;Ebe++1Ie)0/_+:_
=<(NIR)]ZDCTZ)Q39GQCL_:AI[9XUOb20L4SG-HUP&:d-?_===PabC)W.O_@VSZ>
e3#KM;^29&^C@G5:?J_DSV+b).HSO0>aC3\?M]^a/1f6-Z8dKHGJd4LO^7bIXE(F
fM5TFgO?13cAE7/D2S?agMP5_.)^IK]HAD#2?Mg057\XEZBCS_?6PIec^XJg7=6J
8LUCM_+H?,O,&<W[78,LWYM_;K?;TV;OeN30:9A6^9:^Zc5[XW\=JZ(2-:)6cgb^
Qb_3R;1)81aEbdZa-ZQIGSG;RFFJb&MgX,BN,ZP(3g3a]D4C)85T?IX]LL9^eFWJ
=,]VUDV:<()Q=4[.b4O(&YR,<8bA6;)/M:#OE^^F:/8V]d#M[(?L>gA(#TV^XW6N
E^\GR3V,d>=0=VOH)M?NPLE8IdX[UX0fLg4S2Q8fe8:LE<NB(fW,M0;(J2B7bBcY
bNF(AA\0feAF\FIHdCG6Y4adTWUR,Sfd2;\<-K?>5]QQD3E<>Z:TA[Q5/[U6>1SP
Nf6P3G\(1:D@bS?aU?(a)VYOe)>L23RSbK4R_Z.;21)^[0XKLbKY#@M_OcG3TbQ;
SZ3T3B2://T[FKb0=[#?b5O4C-T,ef-,Jf7RRRdE,ed66BEGEe<JU5Ie.aU.ffZ?
RI^0gg#J.L&S2\?I^HdA[@&A&3U,E-1X;Gc,=7U9J&C.a=?<?<@:D=d;FV^R):#f
@&-aWI;_T[V/aXVW);/DIXW-_IO+C&6JX7Lc[NO0<:)@NZG8gRJaCba))#]2C=.(
C?:Tc03?PbBT1Da/.8JTfBYY]\T,Y\;Z2P(N-;FE6>_._J-J[4>8:.A9++:7F_?7
U(C<UdVQG4Qa2\Lc#29O\bOU[:\?KfPbLdEAOQ/&AW_b4a##RO4=1&(SP6:S/(O5
:FFWc=\IV^2QZ9N;TF3Ug46&Q_SI&B,Yeg6]MDH1I,RS9?LfdN4W\S1,X_:@3Ub8
5LF7OAdUYIENZDS[RKH65d<S089R&^N)6gV_WfZ@HL1.c-2Q20^M[4cM8I)R42IZ
5eDafJ4T\/c32)R)N7+..U7-WKAPEPG,Q\Y\Tfd/USR)G^FM\Z3?_67UI6_J:CO\
YIc?dHKb:;.=aT5?XWX.]7X1e):0YL:@9;Bd,c1ZfYO;2RO,UKab3L76,4^:gHN6
23SB5[)TQ0RV,;SDIe[N-dJ5JD4&Nad)(]^L^^ddWUI4?a@0,^/T4A/6fZQW&KT0
SF<7KgW8R2BJ@H0AV1?Q42OW#)4-KXKKT15eH]E0Z7+;KV[5CH@+e)VIX.cD8N1a
J-7af@[^\BL3G_f3#PUD^Cb.=>TDV7,=ONef58E&fCQWA+)G)aA0#IO+G>APV@&.
Q)VA<Y,8cgZ,91._>S-=W.G)V5T]94J\>P22>BA&K(Ye+H_.b5WSC8-@\DKIQ3@M
a->Ne)OKSe&+bB+P984@dF245,=M2bC;eY/?gL6D(P<\]dLCQH40C4aB(T@U>9L5
<g\_GXa:a\F19d+O,P]QTI^GMI=SEZ7#,4#dE_L1B.LR>=I&6cK@&,,(8.?1HbV0
P[BFJZR1Kb41ga_]4[f/_9]B/^aTcDNP-fC:EV6?<+ZNT7)GRLDd=F,Q:M+0NW;c
^=UaG]0+<Md[WEZG]9L](L86))-4.U_DFS60-4D.OKTJV987=]F4XNA;B9\gJ-OI
SYX75]&S^cEABR/cH],GMRG/O_(g,G[?C#G[38MWT<=K>eWA7N&O7JY2E<AGF1\:
PA9O4+7^G:S2E/42?4OBP\9&,FeDd(7):[9S^TZPEQA^\0B&FK3A/d:@/@aZg<SH
WW.RV#K<e\63G2DAb^M?IXNQ[SbWb<4:c^?bO9HD8Ge8gaGBf(8CWH<:O/<]UA)C
V5dbAS_^VZC&NO4N;gCgPR?0?QPO>I,V>T.5@-6gf>RG^T=g3G6b]YL>4?XIO=(+
UQL;0,9K]62#,.\AG^K//0)L((N+T=#,f;>Z<JG#Z_72M\()Rd+YBV_OCgP2/T53
8e>^]#5bf?O)7dL3f?aW;IXc(A7Q(0QCSbFEG=@F2_<LM/V28,P&NC@3V17HFWP?
OTcX\T]=_g#8;cVgG)G^1+?fJKP6eXg=IQeCKPY2C^8B=CED0)7/I\:N^]10E5g<
T^J<CN:2b+6S[R1ILg9X.(Pb4WHL:CMU7(?:A^aHE(8XQREf6+J5ddE4>14bf]NQ
><,YX(c#P6#^)6YO/(/?;IT-^VQMA<3VE6&&c0B78\+:(,;D;[M1A?;;E.?=Y+77
[\fYHX,N&U_DdX4F,.WSO;0[RKdQa[(/.K0#7<9[:WA#EX3OG97#\M=\NST(Y1PF
EA,G@Y,5HbS.UAP&,KVeO]9\(3eW6Z1dB/KJe#ad:(I^\>,))2PFXC2;e,:8-.E]
]S]_K18c0^Ta[M.I.Q--AcYdK=B/Aa<N\fI-6G(g69#L82#8K34O8F?c;3DBHN,#
K3?\TW)/gX@Gb?S-OVQR_NX-\ZdA=aMP65QP1#MQ0-cJL4/GW,SH-\Hd8IP9,P4[
&a>NNKDP/;/PGe1X@Y&5KSX.N\JM+F70<[;>a\aV:Xc8H_LQV^;15IMJ#84YJ2-G
7E@^;MO^A+M9H<7Ed>VH3293NLNFZ;8NQ=LGfAA^F,)NS53fa=T=>G87S18A8,6N
_7B0GT[82@0^eDJIPEf^bbf776_SdH3_5)T.Ud;1)A.86c+UZW)GcA7]&BYBPNTX
ENNaE4ZWK^OaU7,WOA09HY<VO&gV@JSY]\GcHTB4bB+5+;a_geTM=(Me5)_dR<FJ
.\4KST:/K28T0^_X7bI&<V[4M2#:GI2;fc[5158.O&9K3Rb2/,@\7GPPOQP);I;O
(P2;A;S#NI086.b+O6KL-_ATg?PD-WOKQ@6H=H__6S@9#<U^U#19\d^gWH]=FH^F
Sa3=/2()eJ+AUF\5/&6N==QM,[#6FZM\HKc+N7GFKBe^SD4b#dbW:5=+JB,R1J&&
S.@Z@4#ZU_X;VI=-4/,S@?9L;?1MQ<TL^?^A5JeO5N^a)IF=KRgOME7Y_V5)M3aP
WTV00S745LfLcg-@OMAI2:C<ZbBbI-@0bb_<a\G#,KA+E@-,KV2<D]2+UXa@BNg3
H<VZ/GMTf##^Q<.YKcJGd6W5#V31S9ePNd0(a3E6<)dJ>_@?B>bJ)Y-C&V,-.4e<
]DECc3@9R.:CLZ@2=G+L+JKXa_\0a2SUM;e0HO0O;5FI9;gY862(B@SYb?Sb7#>@
;MIdg8eN17@]g2K6Y\(1+WP2Y0=:E<[GCI.bA([Q#=F7dc-Id<3BB8/P2V4ED4+e
EY.,B@a?>K^ZA,P4LWS2_FS^A]c&AOG4P60g9dIcPC1eXVD>9.;Z.6GN9I?4fMfA
fB+:NO)B;EGF#0B#9:6b]P62bNJ@G<ab.;E7WLdd<5[K1,RI/->5YA7F8fM+ZOSL
=IWb2.Wf.=[&(A7O^1)#>(G9TZCC&+\V&].@VF.\cI=:.eb1Tb2=?;R+K=OKf?QG
Y_dYT7)ZQRfNg8+8aS;DM[XF#MK;S7T;I^dT4#0BJ_6IS;B37]g)AVg:ae,^&_IR
MV)WYJDf6SDReG>?R4S4C&#;A#VHa4@Nd7MG1e>eWJJX4^1)[:Vfa/C@\CH3#.c[
VS#_].J5-5P#/WO:H<T>O=PA\KLKL@O\OP2I-<dIb;aQJBaaW\,XQGU62.\259a:
>U_CQea=[=OC90LR-R\\b,>+0>Lb<:G[-WHQ6/JQ]1RF2L]620WeD5Z]fO3XeDLU
6?#bI8H#[_;]NJ1DXQTJ8H7IAf5>=(g5KKK?)E/\1)-E).KdVD)-P>;&;#A[d&Re
UBgb^B+BeBGRD8#=T.Ya?9LX[Q9-O>G[SUWS5N?4c;@b--V)(C_,a,G@)R@H#+;&
a_C,8+@TDI\EA:?^&;GMLBBBOL[;J-?Z-VTU;,+<W]bF2@:QHK37,E:e7N^.TNEH
>>TD^H4LMe@5)^[N484IP#E5-10O^Y2<Pc=W9]-,#cc=f#7+;-UP4?9^Q4-g_.cZ
BTLRU\-_+J)e,_ST[ZVSG+GJ7f<0<OgWFQ2D^C#,1DGGR>I0(&<[PHF;,3JNJ^1/
H0D;PP]R+&(<5TD>H:NLS0J>gYGVOM,]-?baEDcRPM]QA4(V.QQT=)>7Z8]E;5]R
OM;M4BAQ2:+b>E@3F72.L8bYLbFMQ&L@;a,.5C0A:Q@;G^]J^A_.RW_PBRFPUaD>
dde,B4JHQ>GJN&6/MOeN@aX1.5DTAQWR,ZTVNNQ@,gFa+f.P/\CPK1V/F#M<-]Y;
92#6a:IY2A,PR5;d/=:JKX+328d(9Ke,KG#1LK,96).IPF9G>]YAS4WMA#,YPY\V
Z\_GdY.Sb_Y1A^SO^^F1/T?(&T^W;H96d-HB6R0X<I4RA6:YQ4R<eCJY-gf<f&DS
5&49SDce_(7(G4:DA\8+&6@7H30E7JNP7NC[W@IW,H:FT_>8XP2TX10c9;.gc?<e
1]Z09,4P/Hd@,-77EL=f/a#eWLg#5A#DTEITSD[(DU(R&c7/3_.U9M2AR)N,L3#\
aPULBAaBVR+19OI1FUgMC8Q00X,X>-/^?K-GAU4_Rb8IDD+b_XCVdHN5=bN=X-e@
(2fYg[aPD345?QgFT=Af32N8=g3QW8JTF#--0B(=-[XKZU#7V:cY^=_GGUU=bZcE
=D2F<3;<>Od>Qf/(NFP<(#J<Q\cQ;TB.4?Acg)FC-9dZ[2?E9K0gWRU^RJ37Vf6W
7<bT,MI^)VV9KH4YO+@^N&X4+5D<?A^A\(X:,KI8b=PP1@:FR(WRMK?5FS,H&4a?
31^W12eGa:>d60;6c<56AZdGF>)).XIFVP/XGe_M@ZDM92EdR29FIJ@S)5eBLf4H
<dI427TD&O^31Pe0:8P\/Ee::7g6656Ee(_:P\@U0@F>=.-TU@.BA/??\FV2Wg,b
8F8[>(V-B/[<A^6].Z8<GU^4WW4&U]EA4(a8\d7N@eB@(PZJ=;G3E_3P4H_b;ELe
KEHG^L-;1(fOVRZC;]UC^86QU96fI45K+Da\CSZ.f:Y7F-^,d+BO_.XL1M\.:T+H
MF\8a+a:([;R<F^OMKPe,]&b4=4D1@9R^S#[]?L@/)4LIf1:>LVg36XA>4b7[c(g
_1Sa6H7a1f^=6I@]fd(O)TCa[V613fgbEfg\:N:/RD2+?WF28Dfe\Re93:bU]Rb9
fgBgY+>O5Z0WZ0#^=.c;K2e[&1T-HAI@M/\:^d>Ke8f0FQePLgfG+gg_&>NgZ1EE
5[dVD9KZa/SDNL_7)cbUb>3YIU/C7QFRYPaa7a],)S6_#WJ-=7#:fZ-J9@04WV_M
8Y9Ea7<d:S?7ECGB-?DG9Se3PU_:L+0a>^7I::FYbZG0^/SO&G#E5aO[,XD]&+Ea
ZE[YG6J_@,(7LHNb(e;N7Db,6cA[ELKMSRL1dgXXbBb@O>=0O?JQPb3SDG6H,VQ-
2<BE_XD=B1dK5aRQ5#AJdSVQA)FFX7K854H(;T2[C@b^&I^\;\#<H:^.H6:C7eP(
4TQ&3&?c[#JSXGg)PMdOfH)MeEJ@5&5DB.,HeEE4;d+AcIg_H03<MTA<d7N+?^:S
COE(L;Q=3V>9d8H7-=FEE0_3MEI9;dQ)D\ZRG2@97VObEZL\.)IHJDA@JY(_&&]U
>+QTX97dX6(&+CDg6SJ8Jc#<J<\]43A:D]#445b3[ebGI=[3aN:#]g?CC>b>1DN[
a80A]GL<H5EWS0(Y7R1U6WLPY-6\D=8\U^0a=/f(<>H]7)/FYgEbV:345SRRI,H<
d@16]W]TO^IUa@IG0QYO>C[<JeJ>(c#50\OKd0)]-CQ?(?D9[917,B)IF+J;]U@&
Hg7T=-3?+HEF-D//JECPKB,DIS,#gScE,c(5(S1<S/7^AOT:0af/f1@M;<O2J./I
[XUR9E#9CQ##<ecSWf2#?99O?b@@(380^19SQ&]c0)20>TX:0=_R8VD5V0H@C>+7
?OI.DOf^7QJ;fXTcUaC4FS[3A]<]9cBM;Df\WX62MX4aWRK77^;eWWS8/-.X3-8B
.MM[R>N?FJN9+e(]DH0Q&@,_9)6Ze^I#1()E3RN2[LE@g\afE1XG6#]SQMQ_6ccQ
UGS]f^AU1>QR&D5F_,D<S)\;^N7GdXHC8CMT\6-7\0W3#O+\]a<^UdeQJ,g6/[D(
IEID<9XS,/SJgML9J-3d]bDY:1:6Y(8?X=HKV.a_S&/I0GY3?3f8MTAf.Te,)YMR
GXR_Oc96Z5\T[]M_Q0E_.OUe],6-30QU1)c=V@#=I=N@/?3]\D]TXPc(<cHQK/A1
.2S)JVS]#@A.3I+WMCDH>7,_OG,\9\M;4a;L8TQRV?3>53#T:Q3Ic^WYe_bV@_RZ
&b.eHPPZE+>E/gE1Q.S,]XEP910Y:JW3b2WL6<\Q9b0HNb]A&4EA02Kf@)ef:JP(
D>:@VU;&M?(@g(5+eN=;=gNGCDM.Q[3/Y2J56K+QKF2O5]-<EF&.XY<+A;WGRE&C
RVQ<:ETH=/,_?3D)DRb,^IOQQ[[Z9gZId6-0H]e@O&>dHEg?=/NedM8109\HL^,<
W]U.Q#KW>W17=NY:]I@ZCT=c0UCAS;WX3ZN52@@M;C@QRZ,F(:G[[1(FX0;Q97;L
<=cKb2LYJ&&ZcNF_Z0[A=P]9=&0EH)ZT8[bc-DZPN&4YHN]e\&\2G-N1#fe;b2O^
LZG@gaR2^MDF7fNU:SLXH=G?3@P+Y9Z-F0eEYJ_9O5eT8\-b2]LSQF5/DNU/SB7)
BWL]b+G[?8fM:L+-F&dWNdYa9ZQ[O9/Q.\;^1XOWP.<TQP^)&CP6IH]V+?0G=>V^
7Ma?RBEAY+XZG347gA4fQGaR1YPfbK8LC@G6<2ZA.;c?0HP3,AZL_BDd8Y>;23LE
-/fTY0.aM91CI[U+XE&b.,^D(6L8T=5PV@@-bG[7_GLH9FUTSQHD?_]WKa^F&4:A
cRcDS7T6#_1[c2.FG9+L.Vf-H)K+HME?@SA:bKQ[.ScZH.;ERBA@+3Z9aER)CNOR
a(YEH:>84g(7B6b0[/.Q\E_57#D]40+[Y&_X-O9CA@4J9#Y9fb.1PZZ;R#BLMJL6
L-0EGC^^,H<J@=D90d5cRE_-I=LZ2:>K]/cBD9JaB72f9730G]K3;_eI8)7#&@bK
,?3D8P3+?]&_:VI.D(/3Y8]KEa4db?\[/[4>O2(aG@cT#W7Ic^c?aQeT#97^7J[]
/cO3I]ES[Da?TSXH933/@TY]1;;_4_6&<T53;94YDR:,gBBJQ_N<8@I+)Q_C<./-
Q36-PEg-E5,C5IHLH/[8+Y@Q-N0\R/8#@0^AB4[Rba=FE(Sb>ZMB^d].1:fFI]OO
5>Z>8g1W/AZfOT(>OY[1H?FLT0+IaRO>BC.AfOQX]9:TaLPNJY+QX<g_T_SDWe0M
g_7)@7F3Oa\)6Q)C-;U[]]Mb@e)[C[a9OQ\NDR(^>@e[K1>7=^&3X,Wb+4g1UaIR
22?D4.+S(+(fbR\+G-P:27N7:7^5:Z3#B8F^MJe#4&>^H^YJ@8)9,K_B_:#;\TT;
DgIJMFT,(dJ62\SHBdD3fKGb]S;9L_ebM_(U);)5J58K,\<+VNacZb(+?CZD&BOE
#2K+#fT\@W7?<L:+gc^ST\5^ER;I\1Bf2FR&^Zgf7ATT_KE5>:F-d@,HJcbID:08
@Z#(VZ^>P5Q_3FY=X+ff6eP5K/+Gg.5L=^_XG?E_eBXa=,)<QC?3DU;A9>1>>]+G
\g7b7(.SK.F5Y#FU[WGaXGH.O+(O-)Z+;AE(eQI;2a8(HQfW&],U09aN^@E[bd[U
DDfXM,HBGZ32=4:/J0LN&1-1a,5]EP_E<:\?NM/@4UT<\LJ6_EHT\9&VTF2O4gL[
aYccM6<d?;O#D?XV;B]1:ZJ5GgB1^C(G;)b?&D7WXPM+Z/T-\CGc4FDX,e,+a3aT
:g+N-.d85a75b-F2Q]9)bO5KPEC30#3>^.f@-<V:L=>K)M[c9__&XSPMLa_Vd464
PBP/&.D5AB.K@3LQT9IN<[9&@(.R3()2LMKJdCOB+d?M6=?21>N.Pe&2(WOeQ5NZ
e#b)=\2W59W15f)]BKUO6\N][,3g\PO&1]^2LT1+?g\=JYOaDATU;YCWd[bNN,]/
>Gd6(XQ1/&)@]_:AFI95-9QbMT8,P\3NSYPZS)g&VPL(MDbJE6c8,<;I;R=1B5B[
>,a16YafegC)E_Y31d\.R.Nf(e:cZLP/9V1cD@0Ab,c4SFe\9OJLObW2(=)_62=f
(cg=#;/F;e[UP02F]:?+]ZN=FJL@PO[#:PV^W))W[#Tb?+O?1L(W2[P98@:eJ/64
I2dID/=K#Q?JD4>=dFCB-g?E_RCKg3Wg;74+)ICMeC?MNW8QIH#SFP[@Ne2Pb<5?
_fAED]Y3?5@:[.5R,b_4N50);8R@V:D?S=;c5E)La8_:6Ng?P4X^?_eTB446Y;Pd
aa)cFDW+?(fA209Q)#OUY63V0CND\LHJS2c#:N,aDC.0+7UWE/WI7/LQAfVC48b,
V;b#C[(,-c@b0_[3:+bd[]7U?b2>Lc;<J2,6;?,[RDeD1,V9@GGVg31C=NHe<[<E
O0DR(,^>:5gGSbE?H3]NI<)7B)[I35BR2_>S=QX(M850ed0]=9+cBT5P8U+U@9F2
>[:]MI]K\aGLXQD==86;-@d7cINA=^c\[a.CN;KN?0X?>4C:J0[G/fL]W6<;X(K/
@R(=bSe:B:]24d<H[7.<ZN53<DgWEJVZ4BeD4P<e8@-/cfeaQUKEJ+.?BM/7&I-^
a3I.b:U;^_9-g/.-0<HcLMUKF[,]XE<:ZB>U&(V(OCPY>[FHNG./MC+L8f-P;K]b
89+,aDA9f7Gd,-Q;D\9Z^+ac.\XZ(EBf6=f-BCWOb>H(&:J3JYULID4)FY=:P@V=
GR41OG8LB]U2E@F4T8:(K6\e?Gf]GV9>T2Ya_^,R\W(g++M&DcJVNL?TA/B_D#ZU
&^_,.28UeTeb[@8<.&(90[ST>6CGN1KS.^G_[LFW_N48b//R+2OYK9P7e5O@4KS#
_1cU=^]9gS#Ae:Le#47@J8_VZRcNa^22,8W1,g<J]>V8IdMRdg)HX0LUIMHDc4P8
PXP/<=_BT@7&cYOU[5ZeXB(6/I])L0OHI7T>R#4@4+.R_ZCRc2TG_T@#<UG=Td08
IJI-UaSBRf.A..G>Nf5[4a_3IU55=6,<U1685,\LOB@/cR.<Nf(N1RdRTAeJW+.1
6RD]379IdB@4#5BXM30<R0&_egf[E)K(+2a-^5G3Ed\>gEc@G]g:].ZY\A0KQKNG
CUB<Y^:4acA7RHee4B5_RL#Y-E&A?-25<SP_L/4_54P;3YZT:a2UX<YNU#b=cAPc
HS8;A-;FCa>Hf<=86(.B@F><:E,I0AeC#:/\JYLE=?TbR2VVD19W@3(fIT./M=H,
S+>LR[<TB9SJTDb?4Dade6,TLL[G6CH6f,\OYE/Qf[cOg</gE.2(DP,R(=6E_W1Q
VZ>1W>gRL?+?c^c>Y_JUbGR4JU^N@PNaL,b&QDKV.TH2FYcT7MMFS=W7R#5:5QJ&
gMgB<Y[WBNAf=a?&aKbK&^@g,S9?N[O?WIV1\[CB/M_1=F+IH?cX)0\Cc]CQ7J&4
gg>U+3]V-CWL]719JVLf;-gL:DALGM5dN+?ZQ\RUB#]D;]18d0[2BMdJ-FdJ>Y)d
(F8b2YKTT9\2YMUbCC]FH(0\KL7B(L5[[3W\E4]g/ceWR/#EV4a\OC)f4IW8[P?]
R[CFK-)J6dOW-0LcL/Z9.MREYOSUd1(6ABL:W0\09=[T;WFS0_M.LP#Q^0ZE^#eY
L?b0[5T>E&Ga^]OH4(,Y:X4gEbD?#C32bd&]f<4Pa<I,Oe7G40RS?L_<=83?F&/c
F>S7?9^\BWb6.+<)IK-S2>UfC]I[&UZ^QK\Bf>8c46^-9]^5ZOGMA<bV\36-,RI;
0QXU+0H.=?.&TYZ04?6J2[3IPB&@7_<L=P7Y^)#G)[#H.bfeZ(;2:1X.850N#^>Z
d;_fWQ4HJ&ZcY&H0?YXL\4TfS/C?e.SEAHd<dE7Y/R3-3)4BFg]J?<.U55WK[J[L
M770FbKIKEY;JZ(TF@\OfG9Z#<Ie>D2ZJQ.:.c6R4-3[G3.VXE+dD.Z:W2J6WXdX
Db.;Oc+XJ^Eb?Q@[Ie.f\4KSA6#;S;Z[M:Of[[LWPGL/K6B\:Q89Q-.;LR=7gFH6
dHQA)eZB)1c7N#=Z.=&5^?>QeMb,3(3SYF>DYXE4CO@&@0^L;ge8Z.d6HE9H(XU7
RNBcH8C0XfGG<cR5P_P;fV11Q=D>9K2f]/[^CNgYN;WLYdRL)^EeW6c4A<ML^=XZ
TW[/TM1RZ(J-206-IWG\6^#C@3)L-P-?d[g&GHLHV60MHOA#gMSG\NT-WJCI-7aI
\DF-#AWRLZ_f>23?e.E1Q-dN73K<c2LXBK0:#cMK33SFUG&CKN/)HN4+de)R.b5a
N1ZKGJSUUW?_H.YP]:R)GcGC^B6=)NJE>01;BM7]a:=]YE)(KKOb/=c2@VRTQ/cJ
()9CfH7RR;QK7XH,aXP/Z4-4cNR(SKMT4@7b^>A@^OA]M42B<32=Q[cFe>eYNaa5
3OOdOQ?W(D=IB#&26J,_(_&[B9IJdCKf/46HeVD<F^1N\@FO?[MGO13W#b+;/3SJ
PU)CJ0P1G.F8f#OIZ/SO[>0E@S&1F#RBeVQ0U+0MG=X3?F151JaCA_TafVD^4P]3
TL-G6[\E[)NX_<@C<W;d05eT785=OH1I,Y<9V2)MUZ2&>W+VA[QF5U):LZAY,K3<
NQT)5R6JA+3U0/AW+-3YS>8FfaIaaY?U<F_GL?c,8<)[]DEY_<;aOE368MDcN4T(
[PRKS1(PKT^0O_=S-T1:\SLEE3B1]K19be3VYINaB1G/Ca?A])dCHALaXG_Q8BV3
^@VOc0[3YOA<-B@\>EDJ5ZDaI=0BKJ/6Kb62X-NV?L4L,<B/_X?_._=U&eG1F1a&
H1Y.c/7N&_.TIGb),IE-S#2IOg(;cW>@1+E/X3cG],?[b#D/,JZJV]:)K,9YYNM<
7eQ.?c]Y/4&A1)G..<;bN>F[-:5Kg=_D/Q&^F.QdFV\Be;1Q_1^f3;J9HLYc@LPK
R7PKJJcgD0?&6353VBe>G+_+,=&ED<ZE5Q0_]K8X<0,#E+&K>WWG5=?)&B/KL?:V
E?+77)29d^+[YK.e<a<S3cT.>NAB(VGc[HGbTHG,/Q5-S-3>W_78+g=/5f/^H:g;
ELEJY(OF/S=5X8+HEUed)U//0@8(6MEN<&^&9^+(:)DZ6+f\CHU:I3gAY6]\K:@\
3A^3J]+^J.LN-Vc)1023;6S+5::AaZ5LA(O]G38N\1LBE#5(O/V\PV\@aX9^I<+A
[<&69.ZdC8]27N?928(\.2=S@NWL#B[FaL234T#+O,Va(U3A62b2;c^7YQfcH]Kg
J5GL_:Ie_MA^I?Q1I7b28Yc6.N3&\cMY9:;]NaO;)c7Y30&(7I.[aV#IOQL8Z2G5
P/[e\c#OZ#D0B,=33?R5^1)#J?/K]BM/WBga/90Uf4W=F;T].,LUZZW;TX-Y9[+P
>+.8PI2fW+P4,(P7_F?V2<U^1@3IOg/</-;Z6>J+T[X,Y\KfE&9VCGKBJ_/M1MS_
S9L_PN-(:D)eI()N>U?+\MJ^NcRD43>eSG<#9f?]a8R16WJ89EWMRfJf.&0Z.Q&<
EJ1I\;TBS&M)WI@>)I,IB8>fS?P4T4bPY,S[;/IRJA:4I\/1NX-XZ>#M1NbUELK<
-4b+EJgOZ(=7.e#XUDPHTTGG#&93>.P36(JY1JX71)2TUT^ag/<4(f78fT+S?^(A
I4-ELKU3=fDUX+(30KBNN#F=a=3:^:_[eI4a;97B9.#G[1/eL:01/N<7,(b_Cc47
NCWV(KRER:Y^YO9-?SEY3\UL>edSW>/VfVUD[=&IgIY@^S?-a(LM7H_8H(HX4H1b
YZ=LdO-LDa)(^V-RK:NR[2+<XcH))]&Z5#C30ZbN-OFKc5:/L-RMQD/\]^eV9Y=a
+FK0;\DBeLJ0.6+(X0:]V\fA@(0/H]NWV&@],9(f?_RW=/ZUNNbHaT\Lbc:@/.\e
MDEN8?=?/+[<U@;<@b6<]2beM]2J][>Og..e_6X-G^KI7g^eELA<8#SDEQPPbL_>
5)PM\O74,DG&+UMB(E\5G_CU>_U+^a38SR9XZde#=f0gEAF[D+K[\3+C,#eU#YJV
]RA_:G2Oca2\Q(N#F426H&fdJ=5\T=\gc7<^NG<(cbZ;K]bTMdIQ>NIB5SL^ANaR
1J>T4R8fZM[HRc@U<eE\A+44ZWQH>H6)5NQY;[#ZPU^;TPVI=TLZ>g.g#KaC5-&K
;5R.T<J,I.fgLH/7P5a;4F+^7c/JJ57O+^6VOSWJO1?D5SC8SFH0_5H70\8)(,Hc
TB</^M&[F>Q2IGDU;-H&F[L(R)(,<[cdWc.R-V+#_B(@b#)I(QYC^RCbX&Ng+-2f
-gQ30G8N:#8L&_-MB-76Oa2>U5d:Q=bK(f<@B51f;>M6ZJbT4VS2?<GRaR^[cI-c
M1gR4R(8QNIc-fdCHC+ZIZU>b@=]S,.L:.RB<CO?H?dWI-?3FBR2G2g>-PGLaKEa
dQgKJTW7#</N)7fFd,6RMZFa7H91MC&eMELN=:PMS][1:7(S[:N6830f/FPBKbX+
,fPB,EUS)R&J]#2^aYHYg:a++O\8fN.Q:g/FK,F8WZ-a^YAT=4+)RC[:#GODO)b2
/P8d(W5bM)03fBUTJ:SU_/WG=8I^VQ_YX1[W_)6-B_XK@2BAa?WI&=J\H[/11>8&
J(]O+#9>V&TYgb5@-)5TP3d+Y=Z/P)Ne5KH(Y.XR,)X0#T^A:=/1b7&(V=QF-\9(
a--/[^3W7[#Z-42N<;AT)8XW4(@@);2E2J3?H@5ZbJK,\0,SJ]_G1K.N&WW5,d9<
>MYga6>Q[(;B]\@SVZ@.QB0_6ROGY78ZUJ^Eb08aAg?\9U=(GZIE>&dEHF8AE\-e
fg]0:D;8Q4/TZ(X)T?76fF87&4g7A=?D5[G>KJ.V/A.42W5>/7JYAMJd6,B^cZ0S
A#6)60#9<UB[cD8?HT2<>d0;IGCN^L)R9CE&F][UE2D2V5?f)A;W<gb):Ed);]0_
J0HEH90ZW0eE1)f>b/E:EW30HC<#W4W&I6Me/^8CM@QD.89@a-bReL26:I;7I7E3
5<-e)K=1,1CF-4+COcP8a^F/^;Za5:S_KJMdYNU(][afNODTXM\V:eW[K,10&WYA
D\E,HOCDI;fZ,J8@-GPJQXJ/MeE7IXM=B,H.MQ(gV6C+9B=T#1&O8_G#e99)a_#C
Ge&A@dHYbbE=YcNZ(L1-)>BHP.YGTdL4f36aP:;)6I[QYZ.@XRQX5-S(;UOP#;:c
YG\RJEd19I)KbaOS-H\9K-[aW4Eb[eT4#?)#K[,MS+TIFS?FACF](FFb:CZdN@GH
1I2g(O,7RJ<G],E^^8LTIOa^;(^F070>f/b_.>,GBVQ4G:d&8HbY3UHWaJ5&bF9(
XA;?+EU,.8#CIAUI55W,#Q+eL160F@2aXe?/2?(_8T<9H;Z;)M6]X50B_e(;:TE&
T[=e8FbdTECEO;]#N.I83=87Q:C\<Tg5CW4LUeK92C3:AIHfCXB@#?ZPg3F4Gda7
5Kf/a5W+TL2-4NLOb<=?]:J@=)]SF4,ZR<bK0Y&17+EMAGJG,6HA^6Q@/N[=NPJ-
:A)d=\3?DX847#MSN&:Q8X[bH#AG/871SGK;#6=dZ-=M?>O32D?VL(-VRLG1,Mf1
-)TA1X]<d@JFb#ULO\K)Ob?QIeUO_NdTJSB5&W-RHX18FWP297[+/?#1_\46P_0T
VU_T0.\f)0I:NBACgL)3\AP987:_WO@GVO?,>=PJ#Q-TOQ=eR,g7O<IY)G&?N@8W
B@7WFf+,W8HDc=KR?3-F?]OF(E,H,F4IF?IY4WX7-_M4b)#:)RH5N<d027:#[=aA
RNZ3#1^@P+c7U:KE--FKdB#Bg3f=<.]M#^P)d1H;c7Q8@#0=W/LYI-2?0eB3a2Sd
@]NGEQ5+ca2;:=V(WZWAg/=P#3NfSEB.<4b(6G\\E;W:,P1YbJSD)=eL8T90;Y49
+f;42b-?;^FV4F+MSCce(d4SI=U\e86B(Fdb3Z:E+VP+J/(_T[>B#U>2FZQ)+f7E
-.>;:2ISSN6FXF#4:>d_&UF.a2F2W.U1f^683Yg]Q<cdEI,>_>JMB)Ub.-63?JY[
<N?&1RG(AAFJUVf<]K=#[4O,8P.#f:^1NWXeF>>@g:8M)AA&GVgEO3+=O&@\;:GN
dH(PS/@GOQc-@,HI(Q4>D(@&Bg?PMBET3O+O7KJLJTU]?1=.V0-8_Pff,L&(M2J@
J.E7&ZC_b2bH4[BZ51A,X=QH/:5&f)5V^I7QN20B>HV2W;1B5EVN<PQ8L3e4O[S1
?^4XBCX-N1Se#]OaR@7dS#b0><VOJd>Q\]2STYMH6HU0PLV3J,gU3JW/XG(/WB@X
PO3Q+HY[QP=P6Z,3O-5b2Y7ZaLWbK>&EK9ScH+#SZgGf?cWD.1b.]=,6Y15:gX#W
K2FHXFW^PM1a]4?^:ZA//.\H@^6FLIPd;PZT=T6MHS(M[TYd>eCH<M3HVE](-b#g
>V7eG6]d7-a49dIZg#]N:4+8f577]2A]:NF)4/bDSDe)(TZR76M.Keda64[:+C@_
PR#d,W8N@6<,bZdc]VP/5RQ0be8@WV]])<g@-<V[L=?NY95a+.5cDa?NZdMV2SYK
RHEE(_K+R(](?&I1U>;Q,.FVR#[C/ECF_e=ML89-)g+@+6S\9MLJC]_XM3P-X//N
[5g@^[A@e==4U_.EgWb(Q(32^(71/UJ-&Qa5)4]BbfcU6MPS2Z0D&Y0eR65[5b_6
@PUZ;K:9Y_8TWVW(\;X^4S<DbUQAfb@E.OEX;/VK<dZ:Gf#RdV<R,:Ib9XP>LUCb
N(Z&PdGM;HJ,GNXJCG)3dZQ]fQ/MNac-G-:+YK)U<T6YcfR]BA/gVL^_SQ.LI_LI
2:LY9]Lf5b6ITR#?2BK_R:ZeK0I#^Jd8EBLKE38:IB_Z;_@H,-H9&A]Caa[3U,f>
/Edcd\b8.[Ie3MH?[+Q+)TO.;Oc/N/=Eb[F<9@BWZ21a1DB[K;?S#/30g+F[D5BQ
fcRL9]7>LR-;7#KA9.^e2PUJ:OV<f+gbUT=8BKTM=eM5>O\&@fUMLO&?Pe)JaO:>
C_CY/g4P:>4<P)6K0\E3KT4-4<gVFO==DW0/2OHO>A&Q>T?Nf?(IeeM8Z:T1\Nca
:7M.7Db<=W57)E-[71FA=],gK(I5O1)\+fV^\bI(4?-:4_gN=XJ/TL;_SC#d,@]N
MX+QPce02fBUO-@:94A@5E2.dA+=?fSLNd?77#3.>HNW?8#VSS-MK=&)XG-a+_LD
0f=SG&ST.K2HV,ef[?6U^+A_5-&U;^gWW]?T(/LdO_aLK=U#;=E<C(SQ#/ULE_Ec
W?R+.->JNSg?=CKIMb8>>F:M<dU]=Bc?aZ:I98[8ffUVY2e-/-YUdB9M:5/_-RNM
d7GRAKdAc]+D_\YUMa#1631)HKPLH@;EJ)<a<aX06KQH>c?DC9K7;OXL8.U@aHJC
H1AFNR?d8IH+HWQ?6AL(Y<5N2VS=/4MHE>/FAF4816N/H+0ebE8-.)?f_7TB4cJ(
65LZfW/L20+K^R9DQ+\gdM\d-A?2O.T6bB@(dAU([KSR2;I@97#+24D.S=D+R9&I
WP(d)MdW=<bFJ^<a)ee)3#OO:3C6Q]]Q9([BG\g5-VG]01d9e^ATI=a,J>BXJFgS
A]98Qb4#H3=_ag(+4D/7,UgVbER7V<2_5&>gfR37Ic@)VQNU6-BYe_7aL>43B\?.
[JG83430?+3ab)Z1PgEccTO<8.BfNeHID-/+d1)KBZEU.#M#cN9D7U>3:C\79I?\
B:WN3N[CQeLY62\JgH?a\Z9?(/e__,SGe2\c65/NLTB;:67-A9c@bUWY=TXbM?;J
.W\DI066[K[^L^dNSM]1Y35:e=&&JAB\Y:HP.U,M+6=_D/#[Q6@/>JLFM0Ag6V/Z
f3aY#Ee#8HW7W:@_UMA@:FcY_-0RUKI/L@(LQY&-1UcEQ:\0g05QXS>af]JZ#)NZ
;6[X]ILCcB>^YO0eO&T);b-H<[c,HRZA99OR/bDP@gVIOb5[2U(LXCC63IC/S@/^
b3&?Oe32OA^OO.TL9dJ^Z=>dPQf<aSM<(+R2[eGCP:7#@IJ^DPY=/LJ<^1;0[@8&
,BLdIKd>>C]I/;FDaBLM1@VTNDADVY,KQNd5<FMK?4<,g@JYF\gX,E)U_EeS=T#Z
HO&NTO5Xd>M#Gb1A?U-H>G0#-/T+fc3,7dO^QMXO)^cI5gC)##e1S@fX@2I1[9Z<
e\V(c_/PeHI=<NbcF(gMO5/=WB-XLL3@=3G<BfY13aa);V(gR;BL(a1;@MH7N<(=
c4YT/Q14ca)=0eA_(/D0DS)Ff5>OaEfd[EQ\\XG+/TLf3]W_TH_>RObHFI<9Tb:Q
55Z2Wg=#UD&C&#=a7MG1>)b<9_0aN<cOae9b_U/4<)@004H==R)+,P+9X-,g@BS_
\43L-_^1]-.Zb&G-,SRV2-Z7[GBdcU]UaF:e6WF3?Y&&.]U0Ncff^_0-R86M[7#O
?-GAc3X5R5^AJeQG:I<b+cG&>[WL;)HOEU+Hb1BEa^.M?;-SIg^bRW<bf0P>6Xe7
&B_-dUL4GPVG(Xa^FY1?^a?><XF6MJd/[9\1Va<V=a[IAf1\H-e\-:&ZN?;M91bN
^VM&O_8GW>5\,52B^<M3[CT<GZ3\Kf:P7R^,I.<=Ge\^?Of4CZV?AV9(1R:P0R2S
FDG[N7,AIVI5N&Sc+RQ0+Xc=RH\ee_V83H+:IEZ?4;WAU,)W>195(AY.dV5[BYMB
^G[]CSNP9K2GEd;MS0:+/aW0fE?\7ETC8_UHZ1a^[LDO.X7bU3Dc\HFQU#_[XC>[
)1VdQe(H?7EDI8_F][e7dc9&cg/?^Z]XNWC?32Yggd0FeZ1]LQ)P)G/S3PELGH;/
H<QB>gUY)\&VYM0Vd0O2d32.(7O]/KA3<(:e:TZ2OHgPW/.WH\5FK:bA\?450KFK
&^a+e](#:/-Bad11fQf^H8SOb@=:bc3/KY4.8P;Kb=f:A@INPfP+6_89e2]_1V#c
3ed(E1C34c3)Z]ZHY=(;GKK[][;?aVKU?E5MJ_;E,@E,FEVD\Ye>gf<2,[=D>^4K
\RgC\ZXX?#L+#<:FSfDYBY4:[g4Z(?@..G;Pe-T(78]8c=.7E..HC@cLHb_.0bD<
?)T88PEEA?M8<3_TfV\3W0Z1c//e&S,IE_W7]dRZ&+WY:Q(<;-KA^(PTM]NKY1XT
]/3=Q\FD1]23UWP]=Y0I2S-\\OZW4O6?+cU70Q0X+KH>f\(B_90E_2(@\U(c^dIM
PR3T@VZ6@VCg\&d/P0(EdX()M;SE3:d]>A7E;[-:H.E/8DGD8,&Y35]3XQKJeNV4
:73G=c7MA0g2=4:T51NB3B3dc6c]\b/SGFVJ&Q\GMK1E4)6D6Y>+Q9W-2(O&#7S7
&[GZ7A;7H_G#N^_I(7=F]L^]PQdFaZVgcZR@00[+.4Z>>/_g(YI7MNBL4754Ae(E
E5e&)0EG5Cb^g&>]ZaU7bgM#[gJ&,)0_8\Nd07bT)aJbR\fOMYdJeY+F/5YBCQVP
T7bH]\[Y-E21Z^G;+]OY2@MeY=]J=fMAT5^cY,+DM-<XK.\)8dOGLDLX_T4#^;L\
f/@:[a5A.8_e@<SX^0M3G97_Id_g(&dR>3Rg:OdLfbQ_A3L0-Y796RAW@)1[J01I
fF]Q\IVG\B#gNdc^=\4&=B_DR_,A6RDQTaI2Sd<d5gb+f@\-L11+T.WV-bgGOA3&
3W?LXX>bA6cVe.a4I3a+E5\<P@7#H4DI04U;9F\SbBZNWWH_F@=36Z8D(1V-J_SG
6cXR9g)N?^ME3(\0SG;R0X0-.USIa-(1Y@fBW#Y3\E@Sab3-S(^2:,@bD/6eCSLc
SUI]O9eKB.Vc7Tgf.[<E9E2f^/;Hg/;#(0]84cOZA_9I@P9V6:_F0e9Z\JK1BY5)
Xc=F@?d/]c5&Q.@BG;_>[XX8?Q9Je>@:=&8de3^.ga-D_Y3Vc\TW8#.&SV4B5D:S
_]e18Ff?#QY##,9T<d/6?L=121^d+1&f/@VKM77>O@EZRX?CYS5FJW-Q,?H(.ZCN
6N/c,a(2?JW[PfOS]GYY[1P#>We^,CSe&)?b3+>fQM^&.SP=G+BDJEAM_81MYU/:
WgFYR6XRgF]7#13SDfGeHa^42F:P1/E_I-f^(;?U@L9/KefBH;&<[Y=Rf4ASE&\&
/,Y7AH3\6fSKb_R#1NGc(5H6@Y<+]AFgR(RR+J2=f28cR&RLB7+91fH8@f:XaH\4
(O,Y7aEJa^SD#adXNUXL;ZHS50-Q?0H6P:@K;S4\?:2D]N&8&Q+aL5OTB8=;WEg7
Q_2A5JC)gR3d3??AQ:ac=4&HEGb7^@1EWEV36X\C<WBQ9Z7cbNWZ_aaTcOUXJYK(
fW1775XJ+4#_JCEDbV038c[65^#:LYC\D=9-7TO5P&P_6<X?\0JZE-[7R-50A2)d
f>+)\,>KcaE/R)cFN<.Ue_3;\#]W\>(3a_^P25)HIRK_<2LG.)gaQD@_(EF-GNH]
bF.?5L.&Ob89a@aXA8#+00]\c_+<M,_.WB45]KQ(LL2]]Zd63@>-&MNaU?<IcD=g
(g1O68dXLN@#ZP[O5;7:aQ=@Qg/2^D3C837N)IZOFSYNeHHDQSe-.0>A\c24,fH,
_43fW/)?9ScYEG3-5/RS3gaPGGP(C?JcI3<=IfdF=4>]?ZZ5H>Q&R\X+98?W&JX-
XUVXX<<7GgJ_#A6-VCbDBST-<G.eIG4g5bA&2WBaK/DP8)Wf]O1d/4VfJMY>T^F6
X9_@X7U[V-JG&G>+f\K-4I+,EV<5@Y?M.]_AbNE[_Bc#J_MU8^c&(@.2X:WB\,SG
a3Pf98:<c&(f8>+fG+WO&F+a;c3+_@#>^R[a):A6W\:)5cK<WSg,gZ\(H4Bc#NSU
,>Ve<5VZTaP,1A1I1LbZEIEc@DGaMPPMc.,-dQM)/MQ-eR(c3LPe/]e>>##FOLA&
:-L4Kb2W)0+),T7H8E\(?VHYVXWV9VNVEe[_EW<D@P0NVG@?\8Qd4>NOEK9cU]NU
.QJ.5?a1V+Wf>65OR3#DeFY2dA0&P)FY(a,I,G6RC@=.V0PZaCb&EU/eLY2c+W&E
WI7>&Qf50)3a/a,9E6N,#\dT(b:Hf&]R7P+:1WD+[L/040aLWS3W8SJI7X9EW7AP
:3ON4B/NO-^_7O9LGVSa\_dBEU573-_,7A1F6(RJ+9PW+RP2T:36@AMS9cGfCW@G
3e].DVK6&IYcBB(45RgUedgHU>QdL^WBU@cC1fB80MgGbP=U5e>DCU,S_=A[8T]&
S6>_B@0F5S;2[6\H>f#6Q\+)GYAWGIYX:ZG?e:A7S/5ad+Z]:]0\^2,?-]AG^Q8[
GXPaYee/0geSJ0;9<>Vc8F]H-+edE\&ZFUM.7/R#XeTG6L]\#[46S9_/P[Z8gW_2
?LS^JB_b^2,W#8GFWFfTA-4^9Z_7Ta,K>4UOI7G\;1WUN3TC+0eNIWaXH.Q05O5O
^CE?T&L_T?81#8@Ab6RBYT.6Mb882EWJQ>ff6P&5@TEKDWP--S,T)J(g;T+8a_.;
BWKN?3=QgY&O3\&8=;WB9Y+;cTD<,6,@<REe>W<=f6?MB>?[\#?aScg?UU^PU@.N
G+MC@@Y>Q>N0N71fcTN=/DRPTM/U1ZfNM&;Za)PMYD8HZF(W-J&3+gZc^PdOG/(4
<dgOQP.S:RMe.B8Sbb36QcT].^35V^/(M#-&cCJG_Q\_BO\<P>L&VK6UF7\d3QH0
B9NRcCBaSL5SM9dK?<2DP^g<dfE(OCVB7S=YC:UW0]&3=<X\E4(XRW?#0#0QV)2W
]=::c@39Ea9ZC:KW9Z6OH^>^dg^?O7FTQ7QG/#+M0VA\_#;=&aC_57\5CE42CJGC
B\.GE(0CNYZM,[c1=BQ2X:LT47<OV=#-6dO3JC31[F?S#;VJB2EQV0[JTFP+P@8(
T<Z5G3A>(_3\F2Sg<+0[/M?6]9/V[Kf.(DB;g\:ZXSWS8bR9=^d[Sd6>9fJ5J3>a
AAaaMC70>:aE@OCAKB=?^H<0,T4Pdd>_U3OU/U@1_[GfR4A0/Ed_\4U43D</#T2&
=P239Q>SX2O-=E+SQGa<c,FSJ@3J-:L\,D/=XU;O50f#<G:CR63e&be6g<>T(J)P
2FJDR8^N[WR]YO(ee_)bg)EO8b3V\##\;QebJeBDb7TY;/9?ZcSHa6@WHe+1S?4H
#V\LgAad40,D9I1[SgEWITE(N5,+g+PE7#9S8Eg)gVA9<1FFI>#]4S<60@=5]-JO
TN816TD&D5,G=B\L7\gNZQ7@fQ]BgBOK=1F4Qeb9gZ8>LY?#71=_[A<3\)C+A0f9
^(HUB8<=ZO7\c:f7_d<--;SN=W@O9LXH49aZFMXe-9BKSRaZ#+-RVR)T:ZHBS\/9
^W)9#WQX>>B4X&I[Ja8T<?<Y>f=eD+:bWR63XdX-a2]K+0I&fQdX?Egcb_#ZW(X/
d.8]K)ZdG)</X^GfK?e;XG&ONJa<CeD]c4L+9J@9?F8:/E;#E;RIL^[B^V]A,I<f
-fNF7cUbMBcPJVIdVXDB3A6^0W4KZ]EGJ51HA@Y]1+I9R,;O>>eZcec[B;_]#Ga3
>+fNBAM4)e?F72ZMGK>ZFTNXQPKXCA6Fe5bOfQKRPg_ecdREX5_^fZ7cdI3J;8Mf
9G)=RKS)3a_f(K+7gRL^D5]H?+TCP+3@Z^e5U__^OBg-Q1I\/D3/^B[b?BKAaf:^
Mb9/C-7C8/_c/fR/AFXbf=)3[98Q;T]L7g_eT9OD3.+>=)O,UE2];D0322&3V5X9
A]f&QY,[1&-A0&;:3AVUYHfP=JCZ-N,NdC)@HW6bTAb<:CBG.2KD)U?1bGWH^5-f
@g:P]/L3N[JHN321ICA?NI^3ACF>;f/e-HR#^<@V>4R<:FUYUKJcM6fY./KO8,P:
F/DSJIeU/PD0;TEYS@OI.FT+/_bA8QFJY84de,78J:+1KNaA)9RH:<T0]D1PYOO_
<g7=a7/8]-B,)OPZJ3M&/UC]181-L[<(]c-2OES[=4AG,THbG9U2&+41:fRTKPG#
GJ#[dJT2,3g6F\DNc=&G&B3@M.3P-#XWH&IPW)ZA0-<H[_GKJ88MGB(NSBF8B?)D
K#M<_R:,9cD3<B\LJB]?3f>,I?SO15-FBaBg0_(e/?O=9-\E1(<0<)HbJaR#P-UU
F=^X@2;]GM1>48)9Y2DA<\.OVN[=46R0@3AT6]bP)GNG/DBbX-@WXKBUVI\L=QCT
MNK:a=].N>H7ZcT5I93/KY[_\4gW8YgcB8c&eBb&=b71_]Ja3K?YE)[LeRZ>:.5R
S+9E9b7]4C0XC^<[b?,VJ(J]NCZ5LMPC:)P9aFCF[L=QCOG=J@FE7<,WM>dV]C8,
A>\abPPeT?0&]]ERPd>3fWRV5)gcY^+:d7L2?E+FeY1\5=IGB6.KR2MO3CRTb.#I
g<fdY2<]K91\WP2?PaWVBZf,:+N#],S9]A<LA9+EE4M^b2)[4[,JF(dQ>XDHFAR<
VfI9a9Z-.Q0]&_C^?I/GSX#Sab_f&+#]8-FLDXXTH_H@g)TG-1^#ffPJU,G8>J;)
eB^&FY8-(.;/VdV\c)R2<2.BgSF@<g@5R8fM+P0JH()PRdI=]<9U[KK)>;U>VfY8
D&X5eFg6WX:^75e[N8/?gW,<L#[8-=K6cG4I1f)1NBPObYb=,,O&KY8Z#\79[?\a
TLgP9?_Z+D,FC4.X(G+&1Y>>M+[NF7fLA5G8&??9^8_33DU>c:7FDPY94eS=LC4J
=@HO77K5-9Z@(JY3,MSe7ON318Mb21FIK#]GG-C>Q?F=T/]2XYPa?6/9=^Q\aOce
&5d5<,cU;FTVcCd60X#IB(XgJWT-g=JCEdM;M-N8SdFX\LJ,8c&[<J0T8aO/[a<2
>G2>f3HNVJ5LdK866;\X1IeSN254AgG(Z;1\G_YIfc14PcgdE<V1UO:Q[He.V.<a
8]_MWeYG7Q3P78c,^I2c._b4@3HIdTdB(Id_IAe]2Ze_dCIVc::+>]BFC&0aCR7L
OO,B#(H?L#fb7@NZIHCWE1DW4:=Ka;-R2.PY5>HFN2M8JGW+@dCX1=1aYf^BK497
?W/GedB+Vf[LAB+3E@<aE?D@^7I;44PPY)JY9L)2IAYfB.71\d1Mb=f^WfDXLEM>
eb.Ee&73cCeQ>eH(bf0-_SB7?^T>:;DNbMVY8Na6LX[VNMO->HWFSHQ8WaAEaPd:
8\:\T,RN+LW4V:37BOUcSdO^.XBY2YC2g<[4VZQ]FTC>#161),dM[:SWgH#>d_.[
FVMIVK]AD5X\HUFAV<O3AA:M?299HgeB,b8W/TbKM?=afa[:/IRd9QXL38>#12aB
74gQSKZFVLTRfXIB.T-(0\5P5Q:@EDXN<0]+0A+f[?c)M<aC6QBW3Y9&KNUJEOc[
(]TBf24(/CJN#Qf.4]8d+DJBB2Hf<g2UK[Y>A85NMc0CgK2^f).N,<7PVOP<^84;
01K8T0=>7fe7&TCdIf/-JQaIUDN3HbD+IRE0C]V+>X_&-0,WI9[J5M8/L=3U7#OP
0_O8cVJP29RENF49=<Yg^ED,<4P6#F\>X\&@>JfDB[J_WdG[:+8AX/:B7efXFBC\
.#4+\<BM1_d.-V/8H,998TMM1Y>,2<?Nf>;_>cKT76ScB__:Af<&RG8F.2/c;^=g
(=[94N06aRIZ;/L]T>FQe\(+^;AI>G=F://>V<\@&;/.=&>e61>?>YJ^b73IVRUK
]cL[XZ+X7(Ydd_GBX=-1YB(^FP+A;#5.4D5W?g=#G,0)AD?Ia,dY7b3Vg;@V<WI)
9.AIP([e.d<;eF1C/e:WDA,9O[W8ee+K0<G;2PAEZ5=eUXLP>8=aIW\-.(7>5@RB
@F39LfaE=.)J1Qg.fTD_L[S/a[ZfV3L:O?:X7>?b?1+K4d39V9c,;MagT&=ef&f+
QP)6:,+6@8SUd,8P&OL,UIKJb>8)+&@a?@6@eX)g:]79c.?[DV2P.dLO<JN23@6;
AeY08bd4MT(CT\40D3J,140/W)6>2/^Y\bF?QLe9a]YB+ZL#SK.Ze6GB@38^a6@E
&BS#C=>@RO/c:#&/NWV;=YF.1NYI1Tg1G7C(4>eE,e/6@J@8XgKSL@YY+_IDb\&+
148,/?1?[PD.LgO53847,-[-O]SU:9M.X[OcfG<8UOZAdTZB0c:ESg)5C5C30dUd
-f\?/;#-bFH27Kdag7P_<J81fO@eY2+UZZ7)<BZWK/7Ude13ZJ#[<WHagC-]:L_@
F</V[_HZbY?P)VX?^:5cI)[^FB<ZfN&<Y<<EPa9B4X&HV;K#LcW#)C8\E4L38##Q
c59?0OEd&K=(ASZ+&#C@J+bK(@=19GDI<+4K)H<+A9b\-a.G#(C7-R[R3CCMZLH6
FD/SC&YL,d[P7V,M0/DP5T2A6&14Q_CNXfA?V\0gdD[U2O\f&3MUMEE[LZa\1A(a
/ZX]a_5b5aP5AT4TMgfH0BXECcP[)/.PeG8;058^L.If^=f5WH:@e-f^1>ZYCKS+
aPF5>G<JfB]f.\O\\,_@>gODLU-d5D;45XXJYGFD?d;H@b,.EVaS:K,E#0Z?Z7Xc
-^;^]Q,]9d.)&<K@TPa_;F@O6E_]9Gc+V[e/CHJXM48\:AWILV>&CO>gU,B+.PSP
4BT:F:++_@1gSbb1_@PW1X)f29FeOULP6XWY6-efUD/0NB46a8GQD26)FND7@D19
26bX6#,,E8O/_9[@JS;Hf6\T]]7>^a^ca)45QaO5L1b,#_g<9Sc>Q(9LeR^gHC&-
\^Pb1H?(-7B<,[AcNN#4E#[E\M7#]:?TS#79:5QeWa4L6f8--(;9[LbU^_Q\NT\>
K_\A&-9fF?g_&90.fFNY<U.>#=(^^PJ&L<Y1J9JGZ(>Z507D>KZ\C[L^Le3dN./f
-D_)C;MCW),Q(5]ABg8)4A[RA:A&N(&GMOfFVZVU2fUPDP8FVQ?a#R7]=8^fLFVO
-bTdGMDSgX@d^NOJ8SW[,b7^KN:;X<F&V(-^G0AJ>NEY1HQUMI+A?5@^PK^B0Y#4
@Z39HgL-8L<)4?\>H.+?>:c1/(>H^7(V2,K,D+6D#R\(<L[_FQ8Ua0Z?]b9<.O+H
[J_M\6(ZY1^VKK/8:-.M]86<U4(@[8UQ(c?EW0\<NSCP0d/WP?:d7ANB;f,c.WC@
2IbPH8>b#NF.Q5U])9EQU+Jbc&K^fc=6U/&;/L.AWda3.9:aE0gC42+>,I/Jb_3Y
64?/^,22JLfNYGCS#LG>]H3WU(c+DAUM)LdEIL2GEDb?N.?a0gMOEEOJJP.#AMU/
RCBU0ceP5):N/KBLX_W:V=QDM3Z_U=0&^O1@&WP977>-HQD62gT>W&@C#,5+#aFH
/.=]<MZNNgLRK=IR:4:RN:FTg?e:I(JgGP2=EUT)FI)&\MLN]c1.?T,4;17.E.S-
1+KIe:#ZYE^=f[TL@e6aP/G//+WePK=VS=)f9_4TL^HaG9YCEf1AF/=G&J5+ZGSe
c4a0.1.b]&fIRUc<a[^4-N]ZfETP/[MJ:3ZHTaO-F^/A1C2]/EEM&DNeD?\b4?g(
4(a1H-/H[D/4XH8cL&)S0A@IdDN6V838;3</I,+;_M<d4<B+MMd8F8Z2(=;VTBbR
T(QZ6OWb^ZAAbJ2=_gQV=ZKMVSL+S1bL7;3LI@12:Ha9\?&J/NgK4#HNM=[1++cC
cM3VfXC#Vg2UA5T2C<7_#C5Ra30(=UY]VRO[KZBO4\O8<1.3)ER.L\H4dZQ4O#Z8
4MZ,;&c/fX#H=aHVAB@/=BD5BS7)7\d&W):1\+OGB)dIg1;bd@>&Y7gQ^>8M\W,3
+(4W36>Y(a_IN&^DF3B?_M<95dc]BX1ERE4<fZ1RJJ\B838Y627Y[:,\,.Z4dG,b
0@HSU-QGe4F+V=[HfP#FX-[84>cNY,-OXcJRZ0B=AJP03MTRX<#MJ=]\#KP___34
cK\#+7dJ4gC3?1N)Z2M:\[<78N1H)TgQcXU]+XDFe4##f^#^&B\<3gLJ6a:5=+Z_
5/[K:&-&/A<P#USB6)ZG(YA=3;FcIN)ZS/JJKU]b7#MJe2#]8</>&]GK/](65-=G
DQQ?#;_;>Md#/F6(QAaPQ1dFV9#[Z4.)_XeI3faD&?Re-BA(9-215RHgF,NEfQ/d
-TH6:5bBEd36274FZ_95MG#M0I7(T6fb:?U_.WBd45\URdK8IYHD8<O#7d-D#?&C
Nc7/dW1_LB&4&DSZG0C];13N+T]>fJ?T6290ORQ/a=[DQNZ&;#LbOWX.,6#_WSLQ
e_g<4Y4M(;20-XN9a^;@A,H_W=YAZO^S6J,((FCJeMU3XQM8P#MC_S5.KKb.fMJ8
MFRNUbTTE9YM0/>g1CgaNf=,>BQ#HSLPd_&OYNB#Yab#WbXT+#80K?)A0Ne95TVT
cY@I3DgRJ]...VMfEGE7-c,\3dPNA0KEQ<0;?/e5=WRKbGUBS<U\9_NR&[.8##J7
aGS5SJ]JC5:=aGYD),L/JE8F7e(]a],]@WV5NF3,N\3?N[c/O;L\6[)W4Z]#9AGN
5M:a1QMa.5//>dB7-OWFaeVSO5>3abA.PD8:P,-H0@DF-/BS<+X?@3#g&^b1D@A#
)P6.2#,eD8eP)KSDAdbSVWb-b81@aO7=XS6^RO3(E0Gg)Y<#<\BW#Ad,.E0MA5-Q
<J5-^X=7O_J&(aCD+gG:C4;3_Mf::0(T2ARBV;<A:LB8#]W8L9_8P0ZDN>E:.4PZ
E0bO?EO+R(b+>d/]5+g4AOIT5<9A>RW0F,R(2/AEcXM]KgCDgDNHd;BYNSSd.IZW
X@,EC+a4YVef;CA^Z#;RgD5-Q92B<&J^9_#Y&-JOQ]_=1a34DI89?:T^D1g[1dbb
@[+?2(]7FRV2NQS]1_)_Q,95K4JA?&-)PW/QJ?SZ[+RJdIeNg/KB<BOTd]FW7TA7
W.+JTD#JFLKcJS#_/V6;[[2V[)0caV4\aJ>V;B3--0gYZP><7T-Z>]6PB__RYI1a
bXdV7S&:.5_PWX@SYOC,XU(8;BE?Y377f\?18P)MFPSg8VBR:6^SEGK,MH2RM#E7
:EGc_Z)W+FY9APLcWL+5Te1Q4XWa=bCQ1GegZK:AWO1.fC<1?gE1]G)df/^82\4[
CXg=#?YO0F;0NVR:6))F/-=fa_:ZS](BZcVXN0YJO:UeYbR3=CLgN\ELf3^7Hg2_
>X39I+H==C07[MCXTVHgBCQ5eaGV5?YZ1DC_@7C.[dV@,5)4F:^8:5LPd@;[]^XH
CA<=GaSZSd>7@UX6babX9+JJOFI7[]TO17EX8=caV.[VI;L/Y;DVab>5X/H@aS?H
b3.G,JeKO0E3Gf\4/eLS-g\,5Af9W4?S:0W@EgOg(:>(5P/>DSDL1/;dEB-bY5d5
Zb@Id(e.+gDP>KD(2_d9c#0]S(OQ:P0&Q6K)5cG24AbEE5,@gB\^BN02M(>3bRV]
?5#N2N[Z6G#5gSB>I7.DA++39X<.G(fJb>G9[1fDcM<,76IM.-4V>[aB+)0Hbb[f
XfZ>8483Z8c;KWL6[Lgc@HA_=E+@Bd,aBBd5T)(_&PB>WAW\AP#Y0R,A\FA]F^/V
N(@<2QG_]5?5N/[\F^&E#b6c0(2J=[<L,)^M+?OB_Be@L8a>;Xgc>NTLC1)-afJ7
DMBKc1X400.Be=bP_NO4ZgJNE1-f^AFJ=764e+=<CU^=?90GD\=T>H81bROF0/-,
<U_09<.)aeKbOF4H8+.c=CQKU)31-9VJ&WIK839(4X&8fW0\]U?V6M3B@_CegJg9
RA.CI/1ZeOA)O,Ha6e8b>&BDeEaG8a1M4J).YEKT6#bD]e<9_>TI5B5E6]K;5_aO
cIPP<0)9PfgXUZ<KgW&Sa8E>WY30LX#FcRe-57gO:P:MDA53/3JVTcfe^3_bO4Q]
/6UE.9J7#]X6<J.U=4]GQ4D;<d78.RE=?3C<NG.IEO[7;-[Y9=,PR1+_YH1M@[:M
SS0<);Y3PUR](ONV70^/Daa_e5eN/PGN0&>[]?_1P6^>7:)0QH6](;OfGW#ZNO;8
SeBZ&)gZ6T2@O3Hab4Y2&Rd@dOKbfCOSUKA./F]ZH)T+eGabB,A.,II=(T;JI>&B
D<gI]E)88<Y6#H4&^Z#;T<C(IcVI.dFLPeRAeQfRBbT?f\P&GYJWFc-[E?]1B3I.
Y:d<KWb6K8&/_PGID_9N(Q@,b:a<[H<:=]T+K_[U-Ib(J2S+YfR6F=-EUeBD54Hf
SO^J5;-L5+^c;[6.NKS+BdN&\dS+ePR?<c14R=NcaeGQYFV]JV&XNg+;eSR-NGc_
4=XJdZ01]Bb>c4cYNbWa9=83Od<XVK_CM#VHT8T]_6BTVVVIXa7M,U74A1M^aD7D
:eK0FB])eZ_)cT4cAV&-?(:\DDZ#JG[U;gI4eFC:;_\O]WWcT]MAF_0NZFY^g[cP
S_G6e][A2G4b3;4gO+IVEN#^UGQ(e@<FEa2fR4_aWNeK&G?eEX@)7O+T7D/OCHCD
cYDF3#)RDF(#XbY#S>=(aG8)#.H)I#M1M2>1:^N1Y8JVFL^@T4FWSZb]a,Ed_L8D
9Q7Y04JN.&NRS[[CD#T5Y[F/5YC<7dH(>[F,I-Ka-2,05^<XYC@/UZ\F3BW9:D1H
>&c@=Z;5_F<J<@;Ld53IX6XY<OM^:L5592L2)HJ,F9,+KC0ZA4AG]D;&8TH72#<[
CGddI96&5OI>20TA,MN7WG.8WQV<8B2X[dKD1,4IE?1L:+/LeXHDAV;<J.?I-)Of
650@2M]6J+@Z^GS;LF+C?<B2g@bB9;IOJ:MNZP&RBTEd<F-<a1@ZD7(U57,&-?=:
+2OO)IH^_=3.69;0(&@]KFdW8XSOGS\+2VdY_:fCWcKWG/5WLMD.E9&Y)^aDRE)I
_f/BZ]98P_RWe@Y=eP^d(3DafH\DSJ_-I80,UCaIWA^PKEc4[^aF4.;=6^@FD/_(
c]9R89EJC=eDYFGM;QfL,d\X:#N9SP<bNVUIZ\E;<E#1FB;V7d)\c^&JM2N.:WYM
H+\<,bB_E=eLDF-d=F[+N&Fgg\O#BJ@Ed/SWdW1&RNL-1>7__,UeGWE8-PR@f)3?
..\[3fdF2g,<DJMH87(E;9GFDfR2YU380)]\VZ;/EBP4GX9facS2LHQ2<3=]U3>N
_S4A@D,/dARd(SA?,9P]9T[9/(g1eEKdM+D?KH<OOXZ1AY-Nbf\5J\bgQ]]c@P5R
F6b\[HED,Fd&4S4g[e5=LSbPa/MXA&0PO]a;/0OS8Za^S_UJ/C38418:LNF\86cP
6:VW9e<c)EYJFKT)/-f.d8>c1K[0CK^_NE-WLbD]?<0/EPLQ4HW1?S27Y9]VVI(V
F>:=BIV8gH<H\EReRF)2LK?N91H)&FFgHJ77aT?@2+P^-3+KJ,P/M@Y-FG(e#=,A
dAM(6_)Zd>P5_U,a6bN=0NXa>3,\YW>ZUS1S@HV^_/YG^^)YNa-S)g2WFIH[IIYS
NK)=aeHL^aP#?:aP=L;W&+P)VJ_,K>]<EH1(9=7H&M0Y0c[>JH1RS=8A.<C?;-/@
G6f#,a.CVO,3aeeJJcB3##PR+=;)NUeI0bL;+R16>2;4]6M]-FcUW,_?c@g+b@L:
O]MfRU&M#T9cNDTCMN/DZUB4Z1&#;3SNM&M\1&7)/g-S:U#R;?f4GdHO17)]]^5(
&.,GLXK,c1/gV6B.;\ZX?4<\F/Jg5LT:g]QO.3JAK,[7XAa,56F)DX?KdVETYV[/
Q9-/g.fI[(BGc29=OV6UcD9Bf@9(_#B[TOMGWd3EQO(5_A4E+?_>3A1C0cU7@8]f
;ZW(S1FW1[=9BCWBNS-0N[,WUPH@5Q]gZ5f]CXg5]W]37>2Zc@J,8_2NN)7SOWV1
.1?RQY3HcKIXOZdf_>PJG;KeOLfJD].>\7A2acbdHd8WSK,HJfE2\A.TKOK\U>0J
bQD?Z6.I(MQH&A:DYR@BA=5Q=d7TDKR44QGdBSX2=C/N?[L\<WVE/\[\fRLc=Kd:
)gAXA9FB;g?BJ.RYI?<B<V4Gg<FL(RTfXMfP4D->c)bDD]0D+NI3e)3UDOeADL3U
gV<Za1<XM9K0BA-7;:dH/[?S1E5K4O>=DcPVXL:QF@7\N:7=WY<)76(P)J:bAFOU
bc8OC5LH=OQ3g(B9D>@0S>/A_;,_FGJ6e[PSLDB<X=R-bC)be#RQZ;H(;6KU5fG4
:D9=S0(1K#TEe0:d:C)3ffL(T<R;>2YY&5He6#W_TX((P5^:=I)fK.4)RZWFB>\,
TR?XKE<5FF)F7O?5.E?36W@F0].Ta?^,g0/#GeYQUE8X7_3I\&=eR/6g>fH31,IZ
6ZggB<gC(.SCIE:,JY)<AcXF__K9;f^SNQ=3BA(4(7B\b]8(B@C\:)524OQ#cI#B
0N._FLV(\=/:S,^,N@4<UaPSFHA@>??;HT90Na0HUUB\Ee1=R9FFb#\F-b6CaC46
L039MC3NQE/G9:6MSe<<>3dU=.F0//39<JP5W]Tb^,#&B,DPMR[2\#VfW(I94TAM
b-T#;1U(7dKfEJc56aU?-A@Nb:bJQ&X4gbe5<@1=a&9HNX:JCQ7e4#g,JaEJ_3C\
[USeFbaaO3f]3_B];]0=3\I\HAZ5[2.RDWJWa:V7(7;25F_TE\W<>R2KBb#84:79
[H#,-7PU0[Ae;#<;3AY2,>+<1bG17RC+H-]O##R@O;O9-<J#Z@-UWUGKU_4c;=OI
-g3YX7[UN/RR,<T8QgJ1<+e_bVDY+2TePT]1RI3aYa5\+\)?6PA_>g7LVd^Sa=FH
9E5[U7c#bQ51T;df/&4N7fM))b=9aU5#+EaK@I@>P:[fU<da4D&VeV]S0?;Ve7g4
4TaK\>MNff/,IL[6JcTdY9Z1)NX9(/,ZZ-#7)U>I1/J,d_=KN-.HbR[[QdMMc^CG
?0JKHY:<N:S1H,[Eb+(>4-9/Q93fON@H1&8Dg?;XF7,AS;>43J^0dVD8/907fd=d
:dT.QAPDW6TT.:.=aMK^0@6(VB4)5^&dZ7>6RC^T6LQA38]_@J0/=C:K=@Zcb(5g
1Lf^fUD\K9dE8I5JJSe>04BSAW&@V:(]@@3:)B44JLA8SMYBBC&GI-gDAgHG4P((
+CI4\7;]6ZL)@[O._HV2HXM1]D?H^_;;>QE&,L8Z\fS,:KBO.UMXT)_c=Y9Ze@9F
IW=079M?G/B&HI<b+3Y\NU+_#55;:a^4#@D4Og-Y@40a;KH,?1-@HB_OF6US(.e4
GP:[B?V#77<ec\c4Y?SOEY_PO+]S36MRR<gbaPSR@-PJF7L^d+44eRd-_1),1HY:
\eMNEeWXUM<I?)2=AF-JWS:&DY9MFR0dNZ2M6ME(cO^.F=D(3Z7>N5^[=:ELZWJa
E+>D<M)7MU6BM>2Bd;F4a-FN#C)U,W<7>O51:I040DB4AE>G@2PW8HYF@4fH7J6I
#8d:(b1ODKA+2P#4-/ANZ-1aPKM\?Z?KJ3<g?V;?bDWZFTg;Q.U-L6Kf_#f-C,LW
8>);1CQaUB9J7a@Ccabba5LN=C<H=_;..g36&Q7V0&I<aW2SbCRX8&4?09K(7Q+Y
NZBCY[ag][@)LfDAYQX]4)U5.9bOW5:Q(I=BH7X.EW[44(H9.PAa2V3C3]V<GZ;I
ID/De<1[XN\:CXOOg9+J1CbZDA7E0)K-e+1gM&A[LafW9XG>K]LTQXLCP;9;4[O0
0;UQ^QT:8&+6]=+1/cZ?XF)4g8GIG#Mb/,C5I;]2f0C:KA34)^.4+U&GXBV8#\SR
?::AI4a-()<98/.)9ZO((43..)\&9Z0cLH8WAR(\Y_2(f7ZH]W1=@P8N.6#V)^3E
PLCTRWcG,aCNAaa>2d,MO&36eIfaIg-((K.K?KS-acWgd8>aR^/9>=21;/aK,C(g
W>f\H1LY99>eJd^#9O(312P\<RLHC-:3Id:FFR>S+.#0.W+abNXZ>CMUdK5?P[M<
S7f^3Sa&D+?\Y&[9<ATT[G_:<QgQ[HB@WdF2]Q)/#10cH(G&OF1KJXdYVR?F9><<
+GTNMLA(&^cf>8\XKL?_<(cCEB)6aS8e#X6:.4F,be^2e,g#_^]\5#4UZ0=H07<M
OOCV?[XUGU+519UeV9EbP._eIgX+A:DF3.a=(WD4E:e,)3Z/QI=U6&.1a+]&A=/K
(@QMEZY1dgK@A)QLLYb80L(A)f:RNB])61FU+];N5=<09fgC4&G7+fD5,H1E.e;X
Ed@4JC2]ce3>]d&d].),L_+Z_#Y<PL?KUA:B#LLO0J]Gd?8>/d?dJ)HT3bLG_,&2
6c+#(Q/EC@;fU.]<_C,7+b?g4(6?9L^dE(]\QD:9fc6dgZ,Pg.U\ReQdca=-FM#3
.Ue7,e=dX)1AMM,70aK#;+E,+\LAK<?VDO32AFL68PgW95)6?IE-9WAaAKeOQH6B
<(f<U/=9<1[2TM[&b(Of+)9/KWV49=L>9F1<9@V8K-c,]Gf\P8?:@b<X6)FX5gd3
.-JVVDc,R1:0>SLM8cI9\a6Y)[EPUfJEX3DN)<NV\&:S-X]M7WI^73=FF0D6@\:V
EVOMFZV/Z]cJRIXEYD:)gGYBVBOfQgd5P<:H<<RG>J,5<H&6AA;Oba&HVTYC,[OP
KVD3[QE:a<F/=#)YTBd<aV8RW/Ze:ZMS.:#@TV<I[fST)/G[<b2&3d/?L1Og_bR.
@Xe],H]D#@-XPL\aDa)J<RN3=62gDc[3K06WICFbd=F=@]0=,@<C)]fP+fDON<YB
+)8KDIW5\5[L&<Kd,]WEQPMIK]\8])FDE)]=5.(dePeMaMR;N)AO=g^EQ7#.5X/T
@H7WAU3N1U;[]\-]CXbZZ?<CS^7d8_T2F-^gU^9,+:HH.fU_,V&\;&6^&cNL.-fN
T_BR9DN6c(Y?]GbLW2fAD>C#79NP;:92e<R6PMFf#-VGA#3O&QUdgMa#4/WNf,EC
dB,1KB#9dK1.L;=V0@3f[SK4XH7P-F()c[=7:&A5(9D_:KF-GIDM?9A67g7S[8I[
JMUc=YFJZc)0VHN9a4_/X.Sa2_f>^3W;:^c]]+c<)4cg4>C+:2eZN/:#;WO?V3HB
.&0MVQ,-T11gH3EN9f7cf6/CeHUcIA34W@+#8TGNe822Lg&HA<S=f7HS3OF<)?@6
Se(R?)DI:O_@FL4.Qf;1Z9.9PN(MQ=9L,N4HE37:=DSR1#^[E\K;SCZQ72R?g\S9
8bg^GQVFcQcP,HZ1bZY^.YUgc8ZR[1cL.a&9S9^G#Q];D)@g_B2A+8,f,12d-HCH
<0MfARX.M?/=4\(H^?V42ecL#BK9?IGE6S4KIed_ET]?>f^3g5[@;_fcY[E;1V7?
BTMN<=aCf)M-aN:P[-WFG-<GBL&&#7N):6)B^HM&7E&EK:M;;:B4.)[PP:KOJF7Y
cZ#D0cNGHSSDAIS3bZ0:T3.M<UE.<HJHL^:)_?SfY_8f/C75B;=R7>:TP_]K&I,0
AeY\U2Oa7<UV5Z=3226<BeN3O&TN=9,CT8\\6#/1GEO9G[>e<H=&[Af=B&P9D9?[
^>\JfIVZ@)LaF?Fb,A:W)1N3>Xbb+F.6])@+XE<Y3RU^#X+cdHMQB>LUWMGTa44;
N-?IS<5#KODAU[&#QCJLPS2L?a1\86]bH:dH3OVGX&>?M6gbU3#\1X.5-3?0A]NQ
HDJH\L(N-2;YD[KQ6g(9_-F;A2O7SH[X<P(MFP:[B+(4E/\_J/H70DR#XMd@)F,9
>]/6H0)9PZ1#BN3_6^dF\JU>-LPc4(&?bSd3E<QM&aMS;-<Ub1Jf;@9.<ZXK8[<+
D@]/2=46/9O]N,T0ZgbaP0_5?\cVV507I4G32DI6)HJ[OaNcL.J+2]K1QEd3B-d[
@aT#OZ7OLH\43CU^J51CWX^N/>c^Sg2G;2W4&+6>@&GM)TTA-ed#EegL7K:4HP49
[;T]2@&O&#3)S4RaTc_CQ6fddB2g;GP>_T-;6/Vb\Lc+^UTL.:FKN?-IYaC.-T4]
J9R,PN\VE9(\+(1#@29&OXW)AF97W0c+]S2e=@,f5/5T>?fg+\>,1d:fP@eW?)J.
XA+Wd+(:g?E)\MQ:.Ga,LWgMB5SC34J&KCeE]7VRO][EReP>g4T0-RE.4O9@T?D+
7.2c):@T-^QUDXLJfA/A[?^(?LX\YLL#C)IE_BUZ;P23O^^_XfVP6ZZEX>,TNZ@P
>dPOb.R@82F02@/,\aEP/+c#fC7.-Rec:,?Wgg0,-2QDA46/BOf-O5E+G,TfD_VI
Te].I/M4=0;8V.>JQA2Z?:)d3:]Nge_46)gg6E=]3O)MY_S<K:.Oc/I1=8CR?TV.
;OOL;[[#?OV2b@V<X]fFG8Z.YB6V#_Hf>J.]d2d1L?b62]b_WDE^7O\03,;Y+9#3
Y)@6N<:<R+.Q::6(H=EJIF>;VLg6K0L?OYAf-B@:/=Z\W/97M/c\PY2R9+XBP+[;
SgeMH9\<0a.B/Wd8L,LW73AWQ@V7WI.US@fW[C/Y^IB9B+67</c:U,XQg7E8;K_T
TaDg,EQPKC<(OTU1[;&&-].#73.VLJ;.G0AX<B^c&M)3f/DA8^)4ED,0PNF+CPU:
E^80PXVAJ6GfNfA)1Pg[V^b2C)=8OZR?YaB:/418S=EN<68[9#8<LecY-.MVX_2G
J&ba29aL@e1Lb_SZ28B;eE=_,7)>dgcIY\9a^JGP0Q^OcgC3C7+.W>V#1FSI4IAc
+^@OTY#N==#XAMC>cd9c9UP2=_RNGUMF(_dTfD[g_)@5N4RfcQ[2#gZI=S<4)<8M
52S)\8Oc_GOA#Q=]<HV,&.d;)FS]G,9&\XK0SLLLfJ7RZe&Rc;^Y?UF@G/Y7M^cR
d2<A2/_gHZ3)2S8G_=f2BZV(a[?bM#bHA7cPI06,TVUgYQSGIZ(UJ?:T?JM4K(]7
AfI#M[A:.Lbga[HHQ:;_03S28J.>ABdR+c<dCB7CU(9JV79?dI?U)/;83_3:WN&X
0adeQ0OOU9/EfeT(8;FMgCJQb4V5[0U8b4RH>TdM:6L)19C.GbFKDc=6UA?VgQfT
+T\ZMg1P<N7T7eL\EffX44g&N2K0]7H(Off@+d(P\@d;^e<<Y@RVU1D[ec_^9#MI
FNJ@0\TG+5QIUc;3_FU-gDe@4OZa--EE(Z#=T:E2F9.)bIH&]L(T]?P8dR<JKf?b
#7/#QKV4&N:N@48G;8QO;WHUZA>Q6ec\;FJ9BVP83YUQ:PO@[O@,R6YX_OFI]>HS
3b=c&5HgHdIPL>dS33QOL0,.^#W^+QC@^S:G@@E]&:QPQK/PS,G?J0;0Tb2dVfB7
(KdY4/SP7I=NFS4_6:5=\#<#-3;f_fQ;#7\L8Y3;?&X,<)P]PO13OCV4=B:W<9&:
KcaR7L50IgA16SB<THA)aI.A1W.:S,bXD]^c@2U#TV_McK9Yea9VWJaACA?]/1aG
):=e-IH?;94\WgTfg3^W\3Q3M=VM80GCc4Q-fE7QO=\A;T9>K5gVIVAF)>)2ZPDF
X2f5K9@>NRLfR(K0Q&PbZ#EZLU^?7<6ad20MA2H=-0>P/S.0aJfgE\;:.BO<KY4b
ZK@.WVRfcU1O7HW5b+E8T6Q?,C<+Y+3E[db+OKWNbbc+8#/@H:,O0C=GF13YU#6.
K8d5:A1#@BJMa=9D[_AJN[>2].5c1WK>DX1=5ad-^3ESAIJ2K^?[-=OR(&5Hd4N4
_(UUgT1K>D\DE.Q<K,8MG0>BVS)_IgbcV^H>#Z9>6)^Y-A\L&T]E,\=@(Q4\&Q&6
IHHNRe(b08):P,<C0#-MC-NYa<f6DN71&?I:c0U.K[.9D]0_QG5-9fP)g?2OX16#
O0LA-caFV;KXJ_SOU@W^6=Q6d_H1E]bFTZ,E.>UKX3UTbKaFNZR5IR,]KAB3-S(Y
](LBFJFWFZXWgHSXMa>NCS>D98=,V<B@7)Dg<P,Td[/B0D[=gF^>H-A>&M_9.X=S
3TK3<(cBI(Q;O4,DI>I3L.#^AYX1-0^/:2;#[f@6WH\-63C&K,J96(bc3]L,GT2<
=K3S_g^Yd+@W0&Y]e&)2ONc)>JIE7CBL=Md(X3M8B7f<bD^8ULD:L.MS(5Q9AM-Z
Cb#IZ_VIUY41_-@OIgXD4)T[RJ^3Z>GR6P3e?ZY,D.adDWK_\MDRZO#]D5(c]BM_
0A22&;<FFB4.@6Tc52Z.7WgKYM_Zb+/[5O>B\17gA(8/W:5/P-U]7B9)&_,20#;F
3.YAJ3]LdC2>O9=@76IF[3Y_(#,4g/LM8G=:#d:I0(IeD^?2/?1\IZF55[b78@9T
c&NeJNI;N301;UdDOW:TOJDIMaVccb)4E#SC3NR>UTG_^5a__,79edb=]=E0]MRS
T1^2=/D=B/::V[BL]-=/+++.O0__>Ced.O@9daf<DYA&B<a2M2>D1?IAddcA2TTc
2.@TF5T)9HN92W77)MX([O^]QgfCP#XJ>X:ESEW]T3;M[JJcS4KEafO#7CO[2d9c
VaRKZE6H(0_3Q>NEZ]PAR_+<0TW&\Xc[Z=-Vbg0IP&@(N_X7f\EPKND@7;dST1Cg
5.Hc89F^g:PK9?.J#d3AK8.)]XE);-F5gcZ#eGO@B:OZQ_S\8?#AfUIV,>&=U5[P
DcNCcOH,KFBUQRRZE5Q+M6O1#0RQbD?951RQOcXSe.,@D5YFC5@NbAV&1>0fUI:(
Rd)Y[@<SO=c2?bQN4U0TYU=3[c9C62P=J>TRM,2/WE4F;W_4W\F0U28;3[4.b4aK
e;-b^<&HbW9LDTF^=9eNLE>>GT-@aUNO2a?7MU?,+6C1RM@/Rf;@1eG4F5R5LLaQ
\O^E,/7Q-Ig5&^RG52Je74Z<,(U0QFE,I3_)BJBUfIU+>[L2cUd^TFUPEN.<_7.[
D+PAGR-?I3NfG[NaYb2g<8dXPUVFF):O8.I(=d:_>bQY9W45Yd6)GG_UIKVfIYf3
cN#TKCQW_/\B-1_)[8W.cfRPaGLQR8[dePV:OOWXIa]/c6?d/J&JL@BZ)2RfP0fJ
I9e4,_Y3[\NWfO)8\RM9+dEJ_>W/6Z(e19DXc2F6-OH-]b(9O,da1D0)6W).(R&d
-N/2.7W&_MaEJ]OP6)&EY2d?c=XWb2V+,-#c4&8<IM:07Ad40U_7c6@M\+-G@I9,
g<3c]<ZWVQda1WHa(0a5fDT2b>4&8BX1\MUOf8IBa9CI3PPaZA)[N+3/L+=G_Z?@
g@<eVa(8F2)1:O81JJF#,)G71egX3_VMUI/#N81,C6Q\\L<FEZECCTRH]/8-XG2A
bBPVX;bD2-b\9IXGZVV/JD=XWHUUO]ed<6)W<990_]:Jb01c]QeHU)PBbACIT.29
/6QH:L)Vb40d-KW=HSVB-]F:E+ad#F27;WUD+71L^#XN:G\U&<?G[ORP15O.&<gD
ZC;):aRS##S[)fQ1;KI/Z8/WIM/U:35&]E]\Rf;5[UZe0Ua5.M-ANR^ecA_A.VKC
2/W2BdaZK[J0GI]MOUIV86f[RF]I#0&^SS_T&JU/C9F5H^,R1_ZVRJTS</:Q]Q#E
/T&8/#UR7E+\M6QgVEO9)0EPSCd61R;P/eP3WJD/FCgQVC:?FOeWJ_?ab[-eKc;)
dfI>eSQ(5EV.[O]Pb0AKGBM1_P1Xe?A7ORN96g@_]V+WUTU2XYIF:.BEG3K[D>3[
.P^^V54MP@a86DKP1E.#HW<]fW)FKceNWKc1]TJc0+-UB,#SA>e+efW4b(b>be,3
\&TTI^/B4Z\2ZObC,c#)CFad6LGYJKY_J&-c?\+G=QfcB.f\14OdY-fCK^gHPg=S
W<>(H\.1Z?]1Xa6R>3=f72-?:X4XO64b72bJ?SHDc/W)C#6Ud1DRe,1aMgbOZ#18
Qb,)FP7eFW.D:?7)a/8dA&BZFA8GY]?ZGLDSd^bD_#N^</L134]-35[aeEaYa+R2
M&HeR,INdJ_]4aHQ[=RL&P\Zg_?/WY2IfDPZ++42Xd9/\>;9A;\RIaCIWXQYZ.M&
>?XWY>U&VT^\&bV>@92A<WAP6@KK3f\(T?gG0f65@>c\KdB3),;9X[Zg@IfE.g(6
IFURU<=Q_2AJ\Y[1++gJHI_a:LG@#UP3-Q57NLX;S803K&],>76UPBA0)5:AAMa\
(R4XZ=FJ)+R(eQ,^A,442]L8VT.]P+^AB<=<5Nc^M5SUPBA2NVL[@?ZGA)=VcL50
=1/B&Q)0/1A&A8E._8SEO[1.B;X^YJ0>H>DHG,d4[8g1417970fXU?(aXBGCXaE4
4&@MC+U?SC3,MA@FXSDXbPK<d?b\?f15]_^1\;;1gL9-+?K0FQCYI?SF<]@TgK7-
,bY5JQ+:IROc3a:&DbgQYP/Ad.Y[c[C:PGZ])@c?)FOLa+EYOBK,Q?6T(E5.KUE]
^@&?L+>:>H(^@5-46P0fLa,H.47=,T@RPCD0^,N^UX0_]U5XKJ(>^f[=HYW/LS1)
2#LgV?.=-NT^;@HCYX]1[\aZVK+3PD_\QZ[d.LC>^V0FEE&S4YL01K=<EaIdI[M0
ZI[QN:1AX;@J_IT^Y^S9-Ka14UW5K^I>ZT>9^#FFJ0DC14=4FOLDe/;OK1538EPc
0)HF<6&&c,A+/G_8f763CfLdC&2JQWdCCTa>7g)?Y31CBNU#U,HGa5;Db8[)CIF&
,53e<9O\-KW)(4P().&(GW2#2:?IQ8VY0W)b60A<8ZX>?Z\Q0^@&@.EO<KW,e._a
g9JY3>WLYOCJ\8Q:79V1/,#TZf.]H./YJ:R2O;QPO,7@>-8f@I63FGS?F-e?<+?,
&_J6f1bH8@T[d=:IRZ<)0g;HPg]_IP7CH][:DV5K_HO<[H#B\;J\D1c-aW-(\_1R
EO8B5V>UC31<&0<Pe<AD-Zb/^[-NT[G=PM:NLM[5U)\YKI_.E?>\8-0QOM\6DF9D
VaM],UKR[]3YMZ&PG=O564/,BB.bFNc(2OPXL2-OK#\agV&A7\+QFW/N.;5X]WEQ
ZeG5W3?7.=Y=9/#,<gA[QX@,LJB#3[&FgP-?S<TL6+=/CO=\3:[6&-+#=DJ-N30.
C=\EN\YBKg5&,SBKg:1IM(9H9.\?a.DA+>\7c00Dd=>NA5=#YGLC^7]<e8I8C;4>
E0cWF^aBU??:]C9_R(ZDX+H@&3(dJKVE+:X^6/Z1N<G&3Z2<V=@#J2WQ]O6J-^X@
@MPW6#<Jc^dcJ#WO:2RIBdS#BX.dBXS0Ue8&T,_:__.:\cWB0JMXe[#2@8PQ\a?2
3PebDdF-aUB[e1bFP#KDa3G\&PPE]C190UQR,?WE(D(WQDR7#:e=HcW^MEAQK-S^
)F[Bd=;eXgSDWgP#;NAYU:5ENUc:fH7A;,f44A4I,HF&6:7K,#Ig?<c&3T<(/.>L
E2bJ=W?-KXGY)BdJ8E9WaWYOA[AgG)HZgP@WCe/2&bV:S-L,L:-V#=,d(\g)VT9#
cGP.-P_eTdb4gJ;Q95]8X7VHeF3(gA5V\N/8(e\Lfe6cSX7R&S@UN/T0b#c7FL)>
:@Z]\3.SZcgNF)_aA6@/eNE:^K./EKO4NcA>)4A)]:_2\KCX&4E3#RS^b>.Q8R1K
4[KbeaQ(c\GQ;<H2DEeD?G.4[a@a,LJZbWL:aAK)J7,9TM(4S_5RTB2E-(&73.\>
KZZ5Z;dKc&2F(QfNT#=PP1d-(/INTBfWO6;U\c?J<M1UX)Kc1FUMfPe;D48OCe(O
6(+J]U)VWT0X^?2_28U+V2X<2E4UQ^fb.O:KETbK,ZU\aOUYFVeHRXGLJ8S,9Ga7
P0HY3HDbcD0_FO-V;E>]I5B<=F1;cJ^[?(VDNP7YXS,E;5EQ^P^f331V+-=Y:B/B
V98V?3-5bE@&3>P[J7._a1J>737F8K+W+5Kd3[[Cf=DL:-WGNYVb?36JTX;IZ\HJ
,TgD)e_POY8WcDNZagYZYG?fV0Db[7,8\TV>0E,=AASU6LG4f-?[5D[2E\=6_B-e
]^[cU5X+IN#G5c0dD3PPJ@,WdcF&32R2?E#gA4SL&;^+.+fAP\4)6Qd.<NDTV<,@
AZYg]5VNCXGE4:dYcB:L7P)AWGBILa@.KP2((+J)H(3P32,_,&A87M@LF&a7fFSO
=2Z^YU6@J7X0E+(8@_J/U;5)7ITZ#VU])2FV/C;Sf;;F;dVfA(JeR14?=&OM-4Ib
]1O56;/Z81/KX-#3EM#If2OXF_2?_=7,L2GTc/9D3KL90<#SA;c@eP_.[7Y.:5(,
aWK4/(DI_F,\.QF_?>DI?WY@Lc?&-<T@f;#-U2VFKe=]K@Z3b8Z25Z.H@6M-+X#Q
A]NFb4N7bYYaWXXB6WPT5WCHHX&@;/FD@\f2cHSY-0g&MdcRHI1d321_b+,a9PIG
6Z4]7VU,8FG-77e[21).I2O\2WecJ.QX[I#5(G0B@10HL[:=NW;6+OUe28E56V?#
c_9Kg30f<A>e5Y2&-M+b_A>ISX-3WM)?&6/&C+e.?\J:+S?TKFU-H[E[UL+)YLE(
[?)GB;G:EDTOI475G4.fWX-]-=E0f\aQ/,LEbf?3N<@AE#0DXD[I3\:6Q>3V0LV[
bU^9:.HJMGN-><Oe/PS_)aN_UM]-SSF5,KFFUV=Z75cfI5G-/^0I4=T@#P=G6cgL
AK@C#2I6VS6eFe5UUTA^8P?AJKg^KT5f1e=7X\&&:YcV<Rc4G+P:EcRPYfd]_J,M
T_7e<TDeQ1>;JMK3.CS0-aFgSL^3<TJM1M[f9FS^G@?;,Y89<VI7\.[=0@__b#Mf
#X0a-25VT34MA,7L-eNa(2P@eNJK18JS:a:a;AQ#ACVE/^CEJg6VHF>\cT;K:P@J
AIT4:cA^&7Lf2-]O+I0BY2[FE44e@4QYF4>SCAQ1a//4(S3gc[XL.Q_YNXg9_C[=
1Yd86TAC[C&8^@E4A]5Fg:dVB;<b/9Y)D,N51R\3)RK>^#23a2QJKO0</>A3F?HO
ROY-B3,fa2e+(^_8X)V8]KIT)YPB@28cU&TE=^L(6[Fg9X,[e1LTX+,II/UXVaMU
C,;7-7_U,YR(G,&?NP+#VY23WALVa\,I,O2AN-43g&e>>1@bUH2,/=UB/JS4)6):
+CgdcPG[2;C>,OKG#M)<Ia-7Y>Y[2?c[)+/Y=OgUP.=.>+&#2^B>a]&SFZ7?@[;;
A9]O:b0@EcW1(M4dQGH;><LU3BPL#8IB?I.7&BR:^]#W]UgY#5RJ0<PHRRd=>/HJ
1Y5)I5\?Ha:c@=0[,D-Z#3CQ^SC&14EgBeC=3OY(\)/^@^FLW]E0;6/9/OX)P,IV
0b1M(VY7OF-AB4?A[29(cg-I^aC_B4)PV;MJ^f:WS^@@De.cE^.T@G818/=CWIUR
IYPAPJf1.GH1fO]Ig/>=2U)&>]J<_dK5JN/4LXFN>C:c:4/&AaR30@GK\O->+D\[
aJ[>^ZVLf#3&>L4Y;DK&L:Ba+O5#WX.91EV3DW??Ue2G#D2Z@QSHeOB&?_3c_gd#
)&1O9)<c/U>481S2O:<\VRZA\TJ@_H]HM:GDBD:OFagCQSE?BD;cebQ2>DE8)aLW
X1N:Q^UG_Dad/2/X:TK791eKb[_^J[3[(f:A?A>K4[J>WA;QOETR-9#-d]3g:7g\
c?GS0Wf9,3Q18ZH;dH4-RNKUbJ2<B:QJ&\-(F@KA##b)[5@Y,7J2BE11<M0=(@7O
>):(T63Q[^=@6DcVDX0,L?N18WQMR80IZ.FEM)4@d>7^48IK/6XSA4[G?0AY-/M@
ZMBdR^S+f@)&@3AX/CDT.-D58YKd>#;Cg3ZLJaWa=<K/DO-.]d1[M&<XL6^E-HXG
/?I4.YP4K;&#9@0,FV<eG>J5YCMC(M)=UD_2:\0_4SY^;[&(15:eCf#e\RW&A?T_
(9^RF);I#B[D:B<,I=L\@+T,W,WFP#cGMV<.</TCZ/fB:NNNNH3,PPMa+#C^&/ES
D-3(2[AaIHG.UY_I<+KaK+Wg8,&@BBKIgX\X]BVH\A?dV+)6ABZS:U)D1Rgb,YKQ
+^6IS=cTe>g.9(^bG>cQ1-+Wb,/:ZXHB9)M@-C]HUSM?H&aTL)9]@[;0<eY@08&0
F?44-G6(.D3N7.-[,cK,(Nf-8RdYf8QZ9MDAETMLdE/fM,\ca1NM+LDD(E&W7We;
\UMeY8dTTd?R7eTO^(Pbb=Q5Hd3_]76,AL-V0-&:,X#Ga.VOI\W<.)a/DYO1FS2,
S(bS9Sc-VJ[f:XX^0QK[.S6+Q?Ef,\KW=UXGT9)<3\097,eb8?4L<ef_aV=/E>;>
Y?#Y<^UWGP_FDFWUQLc9,IU;0>35<XW0<(HN5^MYJMVQV6?64T?X<Bb9926F?8<+
ZAa;X:b=>b6T(ID6&6f?[8BXcf/GdX/2B;Y4;dEf2Z+5Xc[@c@?FVHg7&BI/FYM5
#5(/L=b_Q.>C+U+EQ\L,43A-BK+=I+GSUc1(V8WPVR3L4L+ZDHGP?_;><]VF(eJX
S+A>:()FLNQL2B2(;eg]JaE-C&:#6:[IK\gdAU&=W0AC7dJ^R.Lde\_<>O?J#c_d
;+VQ?&FD3J3Eb^,Rc,X@=L.fA1/8O[2=BGA0gcE9H+D>.-X,1cPLc328SAL;UO/Z
-@>3b&K?QREA,Bb#S=O<XB8=YVUd3f&.8AGPG4IZ^afZOHe/7I&JFVfBLR83D^O6
JV32;JaaQJ0M<&TJH=)eE^4=)f.A:L:JRePDPH5-f.>_OT-X2_e.RT\HeWG?)&ER
9E&V))([/,9Y>GHV@(@#Y0OS>@c9c-:#8S3@6E1,;>P&>(]fPQRUdPM8]KS]4NQ]
R6eL<0-5_VX3<CW^V-ce(3MCIVEC)gZUUV2L,(L-_G5AGXb-(I+Y[Tc5Me]HIFR/
..2#4aP-/<51W^@eZ8>.ATSdPDUgH/Kg?e(M.bX/[AcPM9;#(\#^G2YQGc<GX(SD
CbGWWPX,B@]cY3Mg)ERN1G^e+^3@@;K3&D,]_CI0gJ,2ZS&T+)b]F=[J3_&YYf2\
\g1QA@BQ^Yff</:QfE0X#?9@>\LF,,HU1Y::ff(6&C#:;/f[A(=QQMIG#R(:]F.#
&-E+/5E6U@ga?4X#\O<@-M[S\:e0:dcDffFSXIJG_]P@R843Qd(Z0^QcCS_aF)(R
a?J,+./\AT)44bJ:B(O@6)29AZ@ISPI[X(5?FJ3/bS@..M?T0?[1@.UFGAP6NK>.
5P6T_^8B?6_6F6Z[I7?2)B1A&,0JNZ?K]1WcdBQf>GR;)F&8\J2f[Y^WeN74\U8e
UKf>N;@\;1L)G6[2J_cF@F[gDbc]((C=KeaZ,D\=BMLFII3-W/GM?TIgeDK.<H+R
APA,,1-d,g^VUG)RJF^X4KGKCIIRG@-<3DK7Gg.^>5_YF\fY-COYKS#_@UX.=ZZ4
A5B\5ZI3Q][40V=N8b9VBfEN^KMH2[a=.+^dJ5R\<N=K&0M#G=4<FR+1a,=+U7Q(
^5dZ:-4IV9DTa>F1GHRW<&P_bg[/SOFS]47.8d3EW:=@5#c:Wd77+a6XX9Z_Q\8A
4N;PK,V+@RCQ&<Q>DTW[b_g87.Z?ZHD.]-d15>C,&J^+NIAV&EbHM)J8D5382&>A
6IX02?&EAZ6;[&gcc1[ZT<TQWOB1cE-,:.Bc@(W;[Qc>S6J1=L1(^L0C)&@F\JL^
Gd79RL_^=6M<#[[RYe[7R-&I;UJ8cZPa22T<a59&c?FWTQ[c3QUK/32V;=8QY]fc
Z?N2J_H&,R-MQMf^KF@6ZA0IJ_OB0WI7gK=Q(GWITNJMdLX2+UON2B4+M4g,0L7T
&aGI_dcD;O\UNOVaOJDM[eJLT:MXEIJ.0FP>Z-.35SWI(^7FW&J/U:92VW^W#;/T
]8GBK?_O9-XMWdQLYS44U+A/&,d\.-9;e.H0TH8]7279Y)63#C6,T05bN9]&CWGF
UC4WBSY9^0S464Z:2RO)-9E#YE-b+W=;XK;44-DK#M&3BaA/NOL:D1YP@Z?=C\Y4
/OA1(5BZH3::,cW7IeI=:Df@gEbR-3SU)M<:AP;OTB(-A81(b0OL)DI9<<;eH(5a
/D)Vg^9M37FAUHaE()Y<N6gO<F]CRH75G@gV6<gGb2<\c3ZC9E/S01SCYG\3=IN1
?#2D[R(F@cGS8]gG9)f=#+P.IPe8:^.0M2YX2(OHcHd5]>)FF]-KCCQ6<:]U3B0;
+#Lc0eN6_4.Seg:7/6Oa_?=F^9O#W&9A67dOGO3-&Y6<G::<c6]71X74J+DU-1^N
>KD<UIDEO8PYMLB)/gA09L\_PA/]aL#aeQK-MR(EL.dFCb^I-4B>/B+=a@E<&85J
^J5DM6?BBU7Q/#>Z:g]BK^K&SAEQ(CJ.+-JENQ/Wd)EW&Ca0[cg0&JS#-XZGSbT1
],fJT\3O+&@T/f9Y5DX#<LW6Gg#/,8G(P8W@,VU@H]?OS_\Q7>Db<9V=B17JFb6C
WbF\.NbIN17Eb(2_Z4cbCQ9#dfXR_C\L<?eaBQODAJ_<)^O>T[WCQRd\BP[g[?<M
c^@H(Gb)9HO6T+6>b\.D8(XUC5>,)2a=?[b?=[K08YPeS?#?,E<N-)5S@5_[T,O_
N(@;@g8M9<F(\g-e13JZGaS:J^OVH6b=SGEaLA>5D]74>^9_2=J]LKI:Y+@[C5>L
8#6OIW_]O;[O^g@99dAI+O[?J_<UbCT2X.@ceY[S&JLW4Y^V[U7F\UW-R@b;Wb0(
7dE:(>5K#EEO2DZffV92LGNX@)SIHKIP7e_R)aV/1/cV7TT7GK:@F7T;LO.e7]=<
-Rc9FYX#g8EYUa?5V_9a@KYJBWVF9/QU]9[J_H.[SZ3Md@D=:Me+EaS(>S27aW9#
G0Y]6Z#VeN;0(bBPEb6></LM(d[<b1f/\f;6R?g<+1YIP2JOX7/>aQU)F>/a?TGI
7K2:C&68JfWcG#+.Y.3#[/NEA\EI&FL,8/IdHGa9NCceKQ2YP45>2?#(2=C,7F5C
/N?BTSG;S?T;Je)0L#]]#&2G&]G=G8cA8-gBK(QgIBF]+b23>a4(?C<1IOQUY8S(
D81\7U->CO9dW1+E><4UH9+#b\PP=,G;3)U5HYX3F)//##\(a,]2&;ZYBb/-(<Oa
Q\OMRQFfK546e&=4IVLTUcI03)SVcT)K6&3-7_GW9?bgFB8B&Oc.52,@359;=c0X
7A83-59?^PcPR6_ff]g1:;XV.@H>16[98#\1G_/\.=3PU#b0Y(\&A7#64S#AfdgJ
050YIYd<Cg;?^7C#ecgSIG)&RFQ?X47Y#;?0U)>;d+[1:DQRUUST&N/(6+EJS9CF
6)F^Pg]aPO,3g3/G#Bb&D7XZO[WeQL2ZDS[/0f?d15@CHJHXO&]&)11T(=(JK<f9
<7S+cW0b5R/-;77KbDg4G;bc(OV>8?/d-fNdV^7(BD,(DJN;^;HKQB,f;3Bd817I
92cWHdA7X>ES,5,T_X>5+38?^BGV8cJaDRHAbAL?DIAJ4U:_gcA?RRg3&+T0T&aW
EUU4MVHOI<I@dZR8CXeO2[2XO.F@1.)2:HW6g2#eH6.aC,6UIOOULJ.8<.@JN[H=
-Q@ACd26SF=ZK7(L?GRYH_G01D-FUGI+4=UMHQ0?Y/QR_)2<HQ88_-G8bDbAGNK/
12L3.IR8;.07AMGHGN+9:g\SY+<QC9E.aYEQc[Ig-P52/Ka>7/.,[(S78E7CfL]d
\18;<S>-]R8JN:HM=A#eZg.</6FF@>>;\XP<BbfeLG:IRP4P-)gb/2#_&P>8I0c8
E324.U4A?5.<db7BYJV[G0:-US]8I@B5(c,E^\,\YK,#;?YdZ<FUU2fg9>DVbEX>
XPe[(d0BM/]G\0)867T3LDV(K+/PVeY,a8W2[FWH-?[W)V59^Q6Eg&c25J;fA-B:
]UF((&Ugg@Ub[2.A9aGFg)VK9-@>bO9>NGWV:38)e,,4F+c1BSdP;c56QQC,J>H5
\:G.P8:M0?QCPffN9V+GTg8,3TN9^1=L7_==4LfgeA+FHA]d=EW@1W6V1T@-.c&X
YE,S)1^WU2(EA9Y]P&c10QEHF._NfGK29_6\D82cU&Ibf[QAKTHW.X&8BD8a&2V2
9KE^:H:J0ZC<VT:cd>b5YAQ=.G40OB,Cg5Ie_E.>J2FV22b#V[=8E=gS]=W-EB;Q
_ddGg^gZ&H\U27#eB@9^1QP&<G213LcA<-f(IYU9EI+2Q6Y8^IBG0529dGW@0PaP
D7-RAa^RI;X)==9S5P<.b:4dK9c\P&:=BMA\fc_XCC4Y51,7SWD=6T]D(@INLX,-
g-6^_aWU.gEU_?HQ@<dN0f=I+/3MT\Ief;KY[+ZBW<Q_GG[^/@MN;:2B191S6L[=
,8F/@#846Qa6J.Z2c7P;g?V/4XC&,.W+#8484==X2YdZ:X[TVS1&UHC?Y;?,eZ_I
c4.&[Be\BFL_SI1/),OEHW:gU@EO-N=>Z+7O#/61-aHP/TJH_3N1_^L?IKgAO#]d
7N)_Pa/I](O-(Q9PB\P]S]-cfO<99LZ5+GUURA[Lg2AB]]YO7F>gJ-BCFE(QM.T9
,MQTA_,&8ZTVBTVP:aDdZ^bBR.^1?CAJ.CZTVHAQbd_YgMKGf[V?JC7KY@COLX)4
^G[>0BX8)8[a;f\VWaNc=+ReWOaZ.R32MOVQ2M5c#G+-O09K#Cc#Z:09IUV+PcGA
-/A#SIaTDG:\07bAB8.:=/&e,J5dB(0;V&;^+^+]=GU/?O10X\gC[QHQQVKR]NQO
TU(96+G57f+@AgbOcI7C&7c_5KTC&3W?b=Wg(\7]fXRK#XT9B)(=]\6B__[G1?Ef
A#VXdZ_e08L=V9,=K&gGENbaHXXDY^T[M>Bg(N^QW<gdac17BQ4+cL(5E[F0-^0_
XJC+8H)c7CI0Y(bT)S]G#D\RVf][O+.=+.=SHD?<M.Vf6gdc)b/86R;=OBTMeb)T
ff2PRFK]I)YEIe/6<bcTKcK:<f0^eW5I?PN1;)&f6#QOHX9dOGROeZT\YXTNCJXS
O6WQ<PPeBW30U6LG(^Fd&c</8\@K6QC:7fIgNO+&@FIB;KK+^5\cD,GA;VG07Q\1
d<DZ(e8(SaBKgH(5[>^[D:MD;f1b)K/:S,B35[9CSY-FbdAc5BFEJLMKA-E1\S<^
#dQBCNV-E+bc2XcBWc)adQUPecY^a4>14Gb0]1CW6(9M.K-#6=@W^@g]HRCD?>76
7a=YDMBV[[O-9Fe&PYDW8/=YZ1S.d\#2&SOaP,AQ7TM@\e]4_f=MZ[ga^OE9B,>R
R;FFY8P:T8F99\L[23[6M:AJ&V98eO6M4^-JKUDTQ(\)D>LNH<bN>)D#Jb\_MZUW
Z2a>3U92Ug.^Y3FZJ#M[R+-T^PNZ^ccC)g\Sf@F5WM7Vb7e)L\#1B-#6.QTMP416
.S)T==L.5W3db]\VA6V.1<\/#fS08gMAY<1OM(B3df8SV@>=b/EYA]]eV;/W&3=-
B#APV/M2/B<\+3Q5.W9QH>=ZeFS^J>+ZJL?D.NXA:8+cQbY8Od3R(-H(F]9?6.?0
/d+dAeV+NWC]B2/b&4R=T,ZH(&=;FSI#(U51?HE>gDaDZCe2g/Ub\[W9ORE-7gJ/
BPTD0)#.::<cADdD2#BD;0B6N.M;VK>S)<G>T-U&<OA350bZO#MO(@0O9<7I7>+X
>Re=)]YUJW>LJ/8CK@b]W2AF.6QFH\d-gH283N:B]Q>cCL^D<M^?#4.(._CP:bf,
O55#??7.4NdP0aL75f4d_;2[W6H]gP6-25I+e&-UX@8-d].c.TJ<H.8]4?W@Af1;
C\FI>+LC1aF5.>7K;PMHOJ(#3[-YA9K:>+GUGc(,M5G:;TE<:;@Q&=)U/A7R,Z>e
(fVM+?\ba._8UR8HVC:Y&K,X^8VCH=0CL^BgDH2FP9)R1+R7:Q]&2:gg<DQafC,I
,#05MO<?KX@L_+6#8bfJW5\)0f0^EFbDGIAI/R#F9?^-)#([YE3>W>:cXH;KLCMK
AI=9C?.1MBJag41gFM8T03Nb1E-LC,Q>VWCdda9_N41<FMf^<Q(,bKfRK9J>];e@
\SDe6.+1gG,d[LKOI;Wd&?ZN)S)T2_W0^XYeQ57O\T]DO\-RQRC@cAGH->cM7Y8/
AOb>F[ID5#f::3FAI3+MG?B1dD?E5XQW]G]).5DX?:2U9^DWe1cd]G7HYAccR.af
/gUT&3VE809OK5POY[,=E+IC,U<566/eU5_:+?7DXO]?UaEFb;)Y7WX&,<&YB^e?
,\O9Q]GC8<G9O>^/ZR/^@=5AL(9FWKQdg]6[Xe/<#OTF[LN1<7;C=,4.0&JV@c1^
@86JPSGJ(\LJS_:3[P;gB9[=-B>F4U(7,^BeTT00Z>-28]I9_LPZ/BAQ9]M,e24C
--LF:3cYUG1d/W#GI?U4<J@&a5PGY]Tg_-ET3+_^\b:);\LCPcC]V@M.&8e749:-
&MX>&_]H;Oa:2?T@(/_OD[UBcY?I51UeYH9+)Y+Qab7,\Og58IOVEZfF&S?fHG3e
7;6F9G1g[--RXJV]Mf,_LY=[Od;O=YI#>HY,S[-?We??MB:M^XcKC?&E(&IfUI5D
@(:a5@X?bS]b1\C>OTcD&W42N>^P(&AG,@ZEF>E2@fF+gQL8\NfIPfI16g/6Ec9U
\Qc[XT5LXgJ&#fW5d?(dddW#\J.9@.SD?[_<V;<ALP8S<X2MSVc(Y3dZSM)?JO,(
bQ&YB-g;4/@):fc-#ODF>ILd.fdKK7g&++U?,g4S\(9-?R;M#0,9?QSD.WDWC,eH
c+E+G4CATdG&7-eUM-^V6+dSQW^LOWA/P,Q0Z&P]-3c2Sa7\E9g]cPDHQHL-]+Yc
c5RG_STAfT^VZIb)ZXNTH=EM,0GUaS^^CX\O=AMbeBe9R^LYN\3R\@<8]=+KH:U\
K&V??\QA1Oe4?;fDIa8./RWRA-1QaA(93f_0(/A\?R#:>CSC\(<f^WG./J\WPWDc
,JYV>DL1dD<VJT)VNW>AS35,_B-^N4?.,U]\g#RXaA@D\4,\(2H2/?<a02ObA5Y.
@(JD<FB;0GfB5GSQ3eHUK4Nf_+&:#(d0LA]8d3[\\=IS2EFYaRO\V\+^FX(G0N+6
S6_>8HJ7aRAKJ)W7DIaE4XYHNN[&=AN8_e=aL9]UgE:B#9+(,1Tc1/eN8_]TD,[W
21>=^g</Z)E]CdGbGNfQ6=PU=6C[CJ-DH+N-d[NZDI(79dWW_]JTU[//.C(Jd.-1
M>LW+e5>4GIJD[Y+Ff)ga)/1#MUddX?08KcUG2+Z+A?PZ.J)/ac4=48aWEX5aZQd
JaV]\?VT@0P.Y:V#P2eZV9BG0KEEg&8@EWST@cEa@ZYGNZS\B=XKB>@1M8e_ff>L
8CP?XSJfbe;,&Q))IO(JSNEMKfeAWNCcCbB;Y(BdD,[AN^I,cVR4B[aSVKdQ9>@f
.KI@A,a1JGKB3Sg)KZ,<Eg-E,JKG8TARQNNTHBf+5;J\SE.ZJ&>_Q:;Z<VO58)Ic
)GJGVe(B--?VLXD_<e3M@#QCFH99)-(eI&?S>AE)=1@W:[2^#R1@Y?aFSd<5)KaQ
8\(4;ZPB\_b20)>T?L)4(CDfKTS>XUC^aC:-STP69cc+FE:0C7Cc3<IK]LMJZg2<
U[IAGcYWJZ#2:QW<Ga+Y?B]-]F1(JV<&/)?L(<4,3#&W.M/@RIM<810XZCVPcD>/
0f@9..S9fSDI/<Ua3KA:fd4-_AG]e+,IK6[G>_3)c\J8V_,:GB#RfHVWeN<3,84+
^17VXI4KVG&:A+R8RY4Y=_(d8GHGI<CH&&E2Dc#]Z&16#@B^O(<T@fcQ2^@W8,]@
BRg<(e,,AQ38OIKH]]_/eKQC<_RPR[?RZYfP;Me\\18Xfg+f1^+]UYH50+10607g
=75WR#AH21(MNOcACagY,H(J#E4=RB#_XLXE]cCW\d5E4f8gT_:AAAc>LANE-BWC
SCCZY&.&g?BAcb@#\4OCdOGV+Be#F:L912,1g=87;5=@A6CF3],gA@X07UgZG/7#
7GS5d2ZN\(UgUgDCZQ=c3JS+_,15;V1NOU2]c4U&G^EY#Eb2K18Y[I?HQ#8&[:G6
TPHV[ZKA[Za2OEQ]KYAcf):3R@2[T.P[J2O^+BaQWg&+^M&U8cRGL1)[4E;0^;MP
UH=QXg=CY?O]-@9a#eNS+I94@?=I<0Dg,Ff8^E/V;ZcB;cR4P@NV(&4+9(a(H5<G
PQB3ZRYG=T&00/9G]IFIBARgP-E7g>&/[D?0@eXGOe1B-e=P2F8+BfT;1:EA=3U.
:d(SPV4#60+K1W1>?32;@4SgcO?O2#H/1cBe:U=^+<^C7LG6XQ:I]g,LY-D>O>9/
gA8MYH7F/:-:WO/@e,T1&:HI;3N=b)NU#&WF=AfVK(5-22)28Q>N2AaD(23g:C^K
<54658daABF-_JWWAM-=5^:A,[TS5<&b-A.^+Me(f[V226P7YLBL)>FPg@7E>cKd
](cNg3^F8Xg9Q6+8<?&2/>5S]-#U]\]3D.ATg4,aLXE1TJ<?;.EJ#.;;E0S1bSB5
#:/>@U:,]RFeQL/e/]Y<[5BD<FJ:TY[SJS2)K@&V-[d9UDPK^Vg+=[@CHL4UfI:d
cNGQMJB=R0<LI9A)9ZCHM#/GH6)=X39-)LX,aLgCT(eJLPDT17@f@U2aO;)d+8J-
#c,8fP8/4b,50\EW9=8&E5[09A1/J)-Dd&_367-#<ECR^)X/PY]aRM;RcG5(QW@P
F_;#I;\36<OfX9GSK-WF,(GJE\L_7XW@)FGU60c?24^G6KgV4g:N<HYROW,835+[
7)WQ5Vb[DA,3C:?PFdIS@Jb&8H9.:A):E7d@/5VVQF8&:aVD2+4BZ:2/D:9KO&_/
T.\e-e7/TN2FL&_ed\#bf[KbG7&7/Cgf49+NcZC5)/b]f4MfLBR<&F/DGC/D;gfJ
1QZ+7I[6MK9e=29c)6FDXT@;>e6,B-eb+Z>;05?d+I]d6,7,gXGe(e<)3=M4#\gS
W93>Y0EgGS]GT>Vg^J)X@QcO-aQ@ec7N<A>Y<)TA2-&Y/?#P_.YE?BQ>RU5H,6RX
_.]f&A/].P([YU((]Y.@ffSc)C,\T4-4f1Q:-d-1HNF9)VLS@_=YaZWX=YJ=DJM=
H1EK&U3=V]9\e4[TXE;E1,e5695H>dVHZUU0JAB\FcEJ#I9/9F+/2dV8X]D^f6^N
Y(3Gc+-F><-DA&Mc&Z#fY&+([P8298fVL-.He4M^JD-&49L)/_gJ8b>;MK3H;IIS
.F=<S/0#ZBJg)cXM[=R]ZYSP=HKTO575-O=aE47OcC#Z_K+A\gSPU1eE1cJVHF.X
KW0>e5M_3ca&F<3LR@;,@TYbKMaY;cTNM^bZ8H^9/65,BK#2?4^5MV\=\cSOe)>a
fW_,=:7ZfHT:&OK1.[V(9Y#,fWTc/M6(\9&.eF/IgCM4AY/A@FU_P@I+5F=dP2G\
N/_4E#5Xf3D;>;Z+:5O5?I7HS-;(-WW1E--HD0GWb79Y_BN:Q+&A5I0D2@gCG)gU
eYS(d&<62,CdDHK6[?T;C#.J.PJ,A9PHXRND)3D_&\U,SLVH6NY_R^DN1HPYe>DQ
,dPF+JK35Z022\32YM1HJM6a0F/@Pb-LQYQd9O38T#FZI<83MFQ^ed&-fD(C#B;P
-K4P8UR6QS@gIa]d\D:ASeT=7,8SLW4NACJ=@/&H,f1gV0/e\e>89e9c(4\<KN2#
&=P24H?[0=ALI=4_&MZQaWYGdF.P.cU8T\4T/>CL9@2,B3ST>06eV#<^aO=,BNf+
1f&TbYIGK01cG;R/b#g6A>0M95\Qb_RFITL\+6S<+^Z9T0PZLH0U0-RDUL=E#-^Q
7]#-0,a8<3=Se5TCC;HLg3.G7.g^P97[.7:S8F)W+Nb9^:XA]7[JKW50-<-YPS-:
2d#)^/()&K426Dg4F9K:YL6GTQVFNESVM)X2a^KI<#4]4cU:L\F@I&,3UWQ7/RM:
QWC#[^W:?I]./6-TI?X/3O>_e90CJZHQ2IJQFScbWTR/WCf-/.)4PZWPV0CQM^#]
;)Z?eOZRO9QQGU]^AS4.[[5;Ue-[+1fM\PP1,eJFA>2M[[P+K4+^]<f6g/F04Oe+
.L=P?E#]NCJY,V[3cP-)11WW5D)9a1L_OG;Z-:gd9>EKHcdHGPOZ(d-aA6TTgH/.
I;:[O3?&;[Y@.[UUQ#B=\<SP(Of+:T_<B76B[,OL>H-Je;0D3I@>,T7>QcP>&Re?
^bMeaH0R8Y84:Y;5HZ0^?DcJKTCR.MM#1\b.cdY77062UDF;1?gLSD,6.:>8NN89
U@BDVW53_Z:,MXFb-TeP\HWg<2.683FAD[T?Ea.;SfXRR_\KL(W)B?B+MJ\J^;#d
?8cE1QYC@CFBb.-eB.U1AW4&B&88\VI[g+28a00G7=F/e7X:3Bfaa0@accK(M6Bf
a0@Be8QeU4)PS\JX:Jf2VbV<B?.6].6,F3C4Be@D?E@->Yd.]=OR8,YEQT3:gD))
(.gINYX4BS4H9P;S+OU+>Z+F2FC60=f.]O0+_T/5;UZUL=A9^)DO,<S7cN5?fHVc
GK],M[<H]LbD8a;7?5?^FIMWA>BO5UX&OY)8T@B7#;;MaP0764D<K?3Q/F;L2@0e
-5+V@KOcJJJeO88cI\AGTd9\fg)?^)f2Y>^4,[:(B3=\L(cF>#W>cZ7IbFFKLM@N
Db?=O#(ZWb]&8K9aKF9OBF<8dg5-@56/g40Z_U3XM_18MQaL=+:\H&2X^PGbA<W]
5@E]U[&P_WH7^,WM/?_cQ(80J:O[SR;1(XOc;ba5QOa[)g^:<\K,2fHVV,V_gE;;
CNTW&^?<UX9QZNV]1W[dB3fZ^XfLfK0Z-9?]SOZH\T0CBW6F=.N,U28#IB0]19c=
GaK3ae[@_8-D,da@D__)?,];,1P@?-N;C?\FTLa04#:[K;F<IS30UG,XVYX.EYWf
S.N,Cgb0D;W,0B2VJS7(8L86,7L6+L5#)1e,P()fR^E1L=SU\SZDQ.?e@-;Rd(3N
Z7,?MaX5\0d=DR/4M^R&]]>+(946Y7aN2:3B9ML\ZF3f:_U=f-15.P0VK^IP).EG
62]AC9#K/^(/>8CFDAf_@B40MRS]E3G[_)_I\KW9bFWaGF==dHBU<(39dY,CG.@e
Q_VW5[_/L-5QEF\_MFK,E/8GLUgd&)BJJLO5DC#TZ@c^V[Ee<5,/W;gbN:cA\(W;
+9\Xgg9S?U](dXc<#Dd<24JTEZ>-Y@D8Fa:B+.fJ(+8#1O1U\[#HJ-;<WP+DH0#c
e^U_QcV=L\c2PB#8S)&F7G46;PR&:aEg-8LBBZ+)1>=]B2>gD;dc=@ZG19<f75FV
O(X(M+aA_?XY^);4^OZ<(f[BSUN6;]IZ;>@5/LL>^eCM?e&U6g0a-G=ESTA(K;fb
I(:L#-,MYKeDb]0fc[BO:>1J#.Z4cYD+f4U:J-+PSdU2\Z4C]UHA;+eBOKgN)aN\
dFXe4VV>ba#GRMXa@OfFG>bGa/(E<1DdY]L(gab=_.5Z:,J8S\d37g:a<(Q[0TIc
L8#>eQ=D]G>A]A&8KC\A^Z+OY,(<>aYF,ea)(d&(]O3=MAB:E[[LPgZb0]BVL.+B
\;faI;FNN7-FLB;\(R5G1(Ka>I/_CgM:b[W0(5b57(HNMaBI7OT.<\\\96+?0JM/
e;-D@9JJ/-gc,SSUFe=9Z7JBCCHW1e^&6SF\88a&c)8Re[HH3[-27_b.PZ)\^1J8
^]=_GF[3)A6AEPNe/)_H]gGTO-8]Aef?N4;7dYO@bTa#9D>?#E-3XU9_adNbF8^G
NF8D6-(7<Z@C>L;Cd@L&/GG3<dB21(1GLI?^fTON[^7U.f5AXMGY#?8acO]fJQ0B
aU7K&X)<CIO_dWL_Z,U6\0-&e.)E5TF7^ZDQQ:aZH(+BT,PWNMJ(I.V37]eV@G(8
/e.7TJd;;cMDUV@E&b@:V,?1Z]HLKf#?eT7TE?G(5^\@W?D+/6SO@^1ZbfVI^KPE
0dB1dG\PGf3Z5,UZX2_=eW]?S^bIEHF/O\QRFBMN-IBYXH8@NHBPVf;2/dc8,4(9
?GUbDAaf?3TWH,-CEWf0HY[ZBSIJ+G8#<5FS5])L.M^:9+WSf)X;Z7TK1Z^0L=@Q
W5[L3JROLcSAfGQYYWXA0b2f-941Ec,E[XE4/_+VgZ0/V32,2G00W,[M8c0DTe--
DYNgJ1H5;>S9&@)FZ?5LY;.?4Ec,TKYZeD917_FgXcS?AU4UAV6a@]Q3A[]_4dd&
MMIIb4V,gdJ=T258X_,R>02AJ.P,G5</<4(,-B/T+58YUXW^__O]L-^P-=D;/,(S
9I=gAB81?^dF/0;CKIT2582e]^3DN:ZWYQ0;2&]:@9@LK_BL4]8K:@#/45JFY_4K
H<\IgIWGR(+0M40ZDGDec])c=?151Z3R6PUc]0b0F/VZ=D+WEcJED+<#I8ZR^.5E
dObaeFU5:Q:C@AN#Yb:&f4f-VgCJ[.SNT;M;beZcd;3Z3@_AN;ed^9T_J0\E9YAN
>/67^TMG<6.)O@=Q8Sa[C=LL:V(1_F>W8>Z=;b>BE53NKgDJZg+;[5:B1<_6fVcf
EW&MNe0U^Ed)66I(?BWRb#Bc^E(&W)939eA;ae),GY[.<6YJ0)H^BQ2Dd34f,&KH
8gBJ6N<B_IT-c@A?HM13d_HML8M)aD#[ODMP&.X<#cG..;Z_Ab9AX)GFO^[@6[H]
.bS[9/c.LU+>.2b,4,=9Nf@P<5CbJ28c-=e?c4YCQIOX9Y[/<7<9=7f<beNBT3+F
6f6VJ<TSQU#bAKMMb2RZR4]O9@5TFI,fIL/BYS[LN@[c&afe/#\+QQBZ;OaV6KbE
8;5_7S=^7;OP;N]R5b5XC>3\T,N,2gW]XGO[D9HN_AL@N-7LYB/6,?V[[6/<X.;&
;#/I-/-c3c8RPIZES=\SOO5L5V)X;.:-VO6>F^bKTR,-4)AWQbb=B3X4G3A+&7G:
Yb7dV:8Fcb)Tg;e_?1#8,__?\GegY9D2MVL+/cG8L</,a_N(QXPd^P+>)JLP8)SC
OHJ-IbK.3KLa@SMYFMG&6321K^b:\gO=VQ&Td\\#S+WePDC:01T#^H0b+JN4QVVX
9#bW3.OBcM1+S=V?<,R6[+,eacg?ZC)\KS)9\:WY>3EfZRR3EL7@I=[_JE/Z-A&V
KCXHIb?SFO-I^RfgE?+N8a#]MW@R<1Mb]V12D3W]?G:&>5cRS=aA/,_?bbA(W/ef
:e:1fc4^D.G>bNV\2[cPDRF&TWW=,A,TB=B2;G:L^#K/\\abYHA637S04LYXP784
6NN03&3<ZGg>&V,,Na0X>[g81>b^f4:Lg\QM3[B<@=2)KDL>,]O)@UWQS3[Y4-V.
R&FUBD?<0893DG6^ZV?U.S(FcDTbJZ(72#ZNY5LKd&^-;?A-)0geEICJ=1:>T-Ug
bD+.;_d_^9IdZ.&Wc48^)PZd&BgW776Ia7a(91S/W\R(.QZQC^6Y2A)_-F@B,HYb
Uf.)@]UJaI_RZ6W5:6Ra?\1>AReK?[(T,c6=KGe&ETEK.,>1g(B&]>.Y=X(SAMN#
_.:+cOV6ZRGbP_Y@P<A+C28eW5J79;fWXM+U@K=dA:/@SN<50#b+K4@;/S:.VEFM
R9ZWRKcBQdO1;=O;B;Z:+Q#I7+N\40QaI8\bdNQO@cPGYLb3,d9T?f>[aP?2QGWR
3MIV/Ga96)@SC.N_W=BMNU4[,V8WHNAMcSOdG.N:,F-dfD,>e_gFOLXA=N[Lf@V&
(gO+/]g@:ET?5.3=Y17@@3GI3:UY.Wc<g:A&JF-]acDQV4TO^R.@_LBML+M;Yc=;
#dS6f^(;5b\Q0/d@g.]Q?.-9dGJP/R/Ege09\_RF1UFDWagC+2=P8<Ec416ec7fE
.b<B&WQ2#6LXD@egQfe3@HD60HQV<S?#RD<##c=&P/-gWTFK(@^95#\e:PA&8T?:
:0HT1/FPCIK1FLQ2_e@?_b[XH^#B@&5a-Fg_CGI9c/5N,W_c=35OJ_,/[R4.-24E
8-0C]PCM>+K/_:/BL=FB]:>O[Z?cSI5(W-C-CJ)IJC[IT-BcK2I#-.gb)e26ZD(3
\RFJ68Z-(D_dfF_+f#eV.L#-XfGH:gM.eRTVZdYZ7S<4//?,a0N0c_=5N,5HA_e1
3g<^^.bDe9KTLA9/DB,-GLdXUd4+82-8;I5Q&:AE)aGP:=;c1;2[JNgKQ:0+XIc8
.,-6#PX>/<:a^[M8Q/J@6<N,PCe<2N/Q>(YcD?7HddT;@d;7TQ4YHL2Je#dK#EFD
J,JUe>eHe\;&\df(d8@)-8/367T;4Q]X2HGfW_B\_;.#de8JZVPS_]>@dcDLRA)7
e:T;O\N(H^B6?a=_N,#:R-5b]MMaVK^9QNK=MSLTb(Q#/a1]<S.^gWb+)-T(ZNO@
>B7;&[D;K#4f?/\MHJ]Z?)B/+2b.O\J4fTSW)06F(2Ma-OFfAa<<4(CBA??HC>Q=
&[P9f?-4ZF3:Z0Lg[EHD0CC+&/@,PXH2JQAJ/22Zb/RZ,d17],,Y\A,aBIA^,4Q[
0>_R=0D2P@.2X4/.cO=W;^L.;ABWGY4#CbO/V/\c):ZU<,X)T#2c9)@cAP@D6T>&
XGF1[X5Z<[VYFC+TZ_SPJ_Y9O1B@V2[fDTfFH>e,N/LDZL)5_-a>g6a(1_S24[:9
J<FgI5dQPQg8S-0SW7Tg1#/M)CU.c.3Te[DcW__3<E5PeLZ]XffOGGX#QD2+?-SC
dfPR(,./W5HCR,E=6&ZK/X+]W2N@WIed?2)a;Rgbe#7YTLQ@1G43<)f<PN^4\,A]
))TUX9I@<a(R41\>,4fVd??CQd(SJ-0H_B/IeM,B065?MB^(H8c:WOd<(&[_&=S6
SHWc:XYPDP:;S&1.b8_[?7bJ\9P+@Od&#?3EP,e@&I7cC\Qf,D1fC_V)[Y9,7Q/[
3c/UB-)Tf(^,@<]cR\dX<YC#[]@)]:E/241O78eF0dV8SJH:fWPRO1gH?/HEAZ6Y
e6J6&eHc)OM)J?W>;=^.MEVbBZ&bPgO_D?TCB(TG+=B.1BEYL:9M?bAP_O?136TQ
S3WcPVW#T@DX5;+=BNY;59<VZ5PY]f3,72Sd,E#&,#DX3/JU/4<@Q2&0/1EQ^1fZ
@XVd?bGOKbE9+RbJ-;>Mf;TPc]F(EQfDKdeBVXTd8Fc/&TR6R9X\+d;dW4Oc)57A
8[b<2/d1NLF7&KeVYL.#HLXEUa>#MUUCcXIUS)M^VfEJc5>/B9;+TYF=N<H&.Y,^
6,ISCYY>P:ZCYa-R2HNY1>3H>A:aS\6Q97>U:KWC6CPg55V]]F.g^HVV3[a-3-MA
=_;.M8b=U;YCDc-^GVB#W>?M+OPcG@[FLG-#5:[gG9G#6d<9Q,JUUUaXAF;fB/Ef
\K&[b)H-U<:<9LN@If:\e/&B8)7#Y,8V+eTB/0>LX2fZ&U-)615M(Hg6R^1)5-g4
6<8#32HSXNBBROTXMb]_G]9YM]9.)T1WY4;8<PE749.M:dWNFdKT5[deN:3UA]:?
HDLIN7Z:(Zd_[f&&KC4:O68S0BDGeU^T>C5d_M]CTAJP4)DW8WS_5=E^]80P_D+e
:C8[,A_G?9gPB-C&R/;cc&SH6X>AKf7==0Vc=W)1(_S3ACR8gKNK[DHc^M];G#^5
3JUc9[GQWZDBH+gcGXgM7J41U]R)XffaX<;:UbVN]F=AU[\9aW2=.V6c-R,B5ZDK
FO4]]8>2(L;X\/YNMK)bd27^0HN)TPdZF&F5X6>-,;N:G#b&@<&AGK?OZT;?#FNQ
,)JS2D.<J8^.H/aQ>YD1[O^_1MeG8=cTYFK(C8..J@5f@2,)Y7)PR=J,^B_TX1d_
[(fP,U/W4K_VHZ[+(&aG49,)a.f-b=b9>YEb?GYH=OJ/R(G\:gSX9HL8@@c\+\;I
A#OZH\@C6MGBVg[0R8;6U#fF8V3FZ_XCG2=5HTe=LJ^IH5&I<\D<f9Q[AHS>gGd[
B\E;SDGMM#<HZ2M2O.YT2DGK3MS6FaKfO9E-S[8TLF<MdS6?G@-].MeAWSJNS\D.
^eENc@YT2V@[MU[75c95/STQ=\8F2PIRUPB]EQPZ8&3_]R=IF7_eATI4\)/g0C>E
S<D.3[L:K9Q2[CSDaX/8e1Y^089HX9ea/:6UeW?HI,WEZB<P?B_TXDA#;f6ba0AX
J;ag:QC/^DC8PW@7MV[+7H+#[+:.,_=-eaXMW.P9V7..@GGY/0g;2)f-,Z^PEc7D
[WA2a_AgJ3F7?O\IfL<a4UGHG4EfcUZ]2?eW[DKFb&/&,26-L+ad_V84&=4+/?;+
RcNKc@I1P7W_QGZM_\7L-Fa^93U__0e8?>@DDIId5OM:_H9703B;W2CP?_^IYDCc
8QLFEGPfD]31AG+1d84@c@5=5R7A70#@51FA312E<1Ae]GBO7@.-#ee\)Y.4Jg11
Oa3K@7dL;-6UGNa4UVTJ&FF@?\Ue5C[<D^WU4E-N-eBTR)]&>7ZcAYM+(O1RObe@
+gWfJUK26^.LYG(_]VL<B#P63Y;#S2-0b[IaAddfTX:@4FAde>ffI#5FC>/P-:5H
XPV=<LUf^K?AF[B@[T/ZLVbL;e-3H^FM-e<31SD6>>XNK+.cLQ>96&F,fFdE[80.
FI/&QIY@EdCP0Q,[N^[0HEcAR74;3&_YRUUJ(J6\-&eMK\bE<3fgaZXe2BSO6.W1
\S3VI)-J#H8:f,3Ede)(&8))262#CDN^COZ-3+IT-==IdI_&S-,_?27>MZIW_-P[
]@0WT-,E\S<2+CO5HE:RaJR+C4-P,.L3WOg8\V9G-+NT(&#5=e-]6gc@0aRL0/VR
]^gaT(be:2JgLO#T2?U^Q/deD^Z)]f?-TV05Jg0&LIN/O#)A8a?adb;\Y2H\A(ZY
&9L-V]N?G\e?1;MIbd;29>a+K:bHA52OPM_d5I_FE@/W7e+S9OD_/RM6>M[2[XC]
B84>?5\2YG90-]fV-N22TEK625R^,##_16F7^>W@)O1-=bK_2^,;;NIL_UT,OUeM
2CY<TA+G=YX98)<2f-STdBC+ZP463W\/(La;7EfQb3MOH.+eF\#A6.I&V,>Da_]g
LY5:&\>AJ1.D+]+U1@E;Bbb)?BVgSfB[;Z-JX[=2^abf^0a82+T;L7W7aPC7RB8Q
EG6TOed+eg7b^#gGHX[HLAP2M0:[_,Wg8D-BI:?_4W[8FK/4gM\>)XF962NBUA=&
KBfeS318-8;0LOZfdMbPXY(EGG=@c[GNZZ0P\9E_fH]5([T6JH]ADS=N^[Q)E^OD
0a9Ka)J3XD1B89Ef)5g?RE\Cb7WVC?VWNL=418&@=/.51H3\W(@(:5G1cM<=+32)
U>5Z/42IL)?)8gDQCbS97bWCU[0a+_-\\<Q&e_cETV28SIF[,]07?d0W^]=>&9N7
WWLc=0eGIXDcI;O?Ged>LJ^TDd>=\MZ59WHN4=0JA[M25[6&AO4X.3,73=0&/2X;
;D#&<_,=2=GG.4c3[ZAXD._]T&;MU;43=L)LV0ge=La^QOaTLM7/ZGFbc9EP\/[T
^dWPF9.GU)<T_@M_ZE#f90:VWUXZ0_VMIbT#\GX9]-;/Y?]VQG(9)-d/J..b+VCe
cH]9G]9=f&JV1IV]6QSKa<,D@\5&=\b0E)GD(/SN-P=c:3V3;<1;-[#=O.R-RFWI
O0VSJd5I^1F4YaKFTTa4QQG?S<[=Q()AX4L,/#&/??GR5G-]C<+^3+F6P/W[.ced
gEAD7E@_?fgEEM@8Y6UVHYL>QQY(M],KSSL&H\)85V]@>+W5fg5Z08,<d[3GY.a1
B:6=b@>E@F#\89dZA#.5e@1?^J0I6,1:+HQ^]fZgX?\,+G2?ag)00BP_8XZJc3GI
dZA.I\dXMG@,@3YLOQ?T&94I0Z?B-I<aG8Ha.H@g>SR4_34?P&/F@(,2P[a>9MN3
7DE8E1DNKN__Z?_Q28=C)-X.#\-4g2RR1(4DFK]Y1OdQGQC+)67LF=a/KU-OF&c?
>K-(Vga[?Z8(Q]+P7_BG&K^2cW/]EVS8TYG<?5I[AIee6Ne.RX:F0Kg+;YOB1@R]
R/3b.\ZD+G,&dPS+94U/;&=&2@5)(/E])J4>:O7:D5;5Y?^G49EGD\^Ef0=_ZcHF
aUH@Z9HR61-cFOXY1U)+Cg@NCU@E;)N,Z:(Y2e-+,;Q&<2?.bY,PKHO5c5TRSU3F
+a^G[-FeOT0D1aLQ,KC7B^4>JI;gS\9+N0a-DE.OIa(35fCO2[GD/eN,fEQ\/?4Z
/>eeL_@JZ6D^8?+a]@G=98D;,=T?G+7FfA/[JgA9:3R4&G+J28IG1@e76HU&__eS
>\X36;9egc?-/GFT@#:83g,VXAJ_)ZF[K,Qe=A1D)_[9fCQH\_CXP()J)07WY(=f
PBK<6X8fO0O/;I4dOaX-)GS=aETVL\OE6_:1_S<aC/+G1]6VIf2?EPEB]B2+bNaV
@/O=L3KE4O-dTU8;LDGa:X+2UEK1S<-CIU3]c4<W#A>53;>/\eBFe>dA<UIB\M]R
EOgRDJM2@XA7R-;@WBTMC8W[UUA9Ff,^2JddHbR1D462-VOa#4IE4T,CXEX-K<T:
(/0==E?2.#\CK3R\XA_&[MRPV)W^&FRDNT6OD=)T:,WDJ2@SWXYQ-ES5=)QCfN0/
9W=R9,(V-dAS9@DLL6M+UdX4YZ,b9gK#JCG^-7N2:W3+01\e.)18d\4\PUTf-MB(
3fW:(C_28\fV4<.R,YN<f\L_,>H6^]@.eVE:U876W0L<MSI7W:BCVB:G>e^g;];H
JLE/UG/@Q]@_IH<KE:>XS8>gAM@+BJ<W/,E4TM]N<5(/9[@f=SC5Fe;\b=G[?893
\J]9/9PQ[CCb<VQ4^A_)92V8AGA;3eb[N,39=^02/^V1M;Y)@gW[YX3FM>@#OS8Z
K\GFC3:4;c7HA::eW47Cf&4(<-.fJFG;[CNKINbV(\d10#b9U6Vg#<^dZ;e+)QMU
=7S^:L.=M[_cW<MAVa.8B-[fH?WIM[L)Q\P?XQ35F:ZgG:g),?U_Ua.dA:+&)E1J
KXKG0FFa8+?-D8a<+VU3.2M8=RdKd+4@.7)//7S5DRMN3[>B5bPC)(40]Oa[@TFa
@JBZGK&>)HU_C=J>+BT^7D6SYKOda3EP[U)L_Jd2ccPLYV[UH1:44)U>C3dVY&^J
d?XcB]C4C/-3g.ZfW-)[[DYSE53PB8I\\R0B-P&XQ0_H+/Ie:&?,VD,3IVA#970\
#C1F\NUFFPNJ=P.Ge9abE@K;JXTORAG.=U-b#FM)aSf[Sf7KSRVP=T=0BQ_@K8T_
O9eA,H)eQ0(#9TT_[),b:ce8eEFHfg+B3YP5EFI5C?FO3eYH,g6bJf;N?b-bM1OV
99XO)GMF8cZ,_(S@/G[LDS)##6eSJF#\9+2DGCILZcf67g.ACcL==G?O#O/&KJF-
.I9QO/HM\(^H<&R3]>\57P7V3NT5P]#ZUR5J6,f5@Ma6>#_[1.K,.XD6:-(<8#19
0VA4_>g9-=;2:V.,H&5B/Tc0K@)OPR]<0M)&c&^bQG(P2.DCPC50aMeaCfcML0N.
1[WFQ>[TLb]_]\G9-0A)EE]Tb&)49JR<FeEB]GH0FT^S1<#S,g-\Xf)JFURVfYc8
ZT3?YU<W5>=6?E,EcL8>AI.&/./B#<+MDA0bV^ILN6fTVZf^0_,X_8K\SS[Ue78c
Z[RfNT//T@<Sd@K+-1.3YO9R.T?C0T@e5Lf4eRL/Y-=ab^b#.9DaU(0O\XR)J5V@
)Uae/?1c[DBOB5:8f03=_VD>Z@AZ.MeQO<,1X=E=RU#R&Ag\TM]>C+3JP\R1J:P4
1V,V>1YQ2+R.6--+??]DY1:BKFY[\d+;b0c])EYe1UM<-K]WU3gEIFc&_gX>eTSL
YG5OeeLbZ(Y2\S[FSe+G6b1[Qb8BWa>K=bZK-dMHe1eWec_3.^)N)KZ9N(@0S68=
C:TX_a8bA=PY0&2OH]_E2Z<<16L[VW-a\37V)S8ILW740VSV52[D5X_g6fO)Ce9>
\U/4>?#Q(5(\>P3gNGT1KIM<:\fa,;H=+Nb4PNgc5PF(Db<@9b[##L(:U]S#METB
UHC7==[;6ZH@XZ<INCd3BZM\,?B&X;GOBOWLD],W_gg]?@<M?0YBC[5C:/^:[]aK
XU5QD;2dg>F[/#aRX7IXTc,:/&fW-5Q8@(9eJNdZ?L&?)1_U<0>.L]L,2RW?(2]?
7/LY+-1#e5E+9NaFQU0Teb5XOX@<,)/+DGfF^)U8S3Y-#4]cRAOA<<.;_2Hgb-KN
DUVf(?&#P<@1IP=57H4g8IW4R2eJH),@-#F2#8/E^PKDHOf)]^K^Q/EfY8W^QN4V
Q6:)Gb8O(2egdG0Q8S158.8J&F(TWB>&e89DLXV(8C=g#Y<NcB0R4A3N5g_Y0/U9
gTbLg2O;\D#6c3f(IR&C3C3E]Dd2S#?[g>L3)gA-f_R/6Q4]e+F]4&S?(Y&1D#?[
IfW4DRXSgbfE?ABJ9#/K:#TdM<]@VKfcFB)\TJ/0;@g0)V5B4#f(NGDfZOQ\HSOZ
8M3R;=I(02<<=YM[_,./@^)YF<[e[U)22bG]158-^?K0(]RdZ&AYV25H-K_R>b_G
RV+=[OI&]V<IQ3G,;JYE<P/AQZ6eSNO;QVLZ(A1&#8N>K>HK8A?>T]J2^g16V0A[
Ye(UA0/)Mb0J.D9:[9DBXTN0GRTfJfN.+W[B/KR:0.Z8YK.[DLG1//]GZ[#7?J#L
\<_</0H]_D.@e1TBbFP3K.5I6TO]:)DEg;La_-\Sb1/N.FJ75\c1<]]]CXb2_]95
>WB)W:^+=KL0A:ZFM6R;f6X77@DTTd2@T?QX;\2=6_)I/PN@gC]Ga4>06a4KR@dR
?N>+eTK9X,XPT(F<_M9?P;M81T7Xg(]CW?\6b8XPVR5f7.g;KP>?-\acX9VI2DF^
DS+\N.5J(\]7__Y;_6L?P\7&-FO1C<,-22_)S^RTSd<VRa.DBBRKSB0H=[T;:_6#
c,=MJ/,0U<c?7C1^a(^H/B^c#Y0-XPDfH,(d/FKMW34ZG:&gd>bRS_LQ5Ug6f6.&
(b<e__K3Y>_(<4^a1[NIQRG1/>/ZP;eTYeM873_fN^1IaY//bHF9bK6)=M:F^VHE
YKcG4\aHP&67U.13CT+d\\A4D].KC#M(b9@OI.PTY<S6Oa-^Q5H[f.aZ<&N_]?C[
6aHJPV4\<fc^+DJKH_8/S]GNS,BTQ:ZT]?].D]WNYD6g,\1@RMa:RGG973eW,+Of
EbE#63+Q58c-V_MG<d@B.e(BNc[7BQbF_?]B[e>29K>9cZNI3T.C[Mg<1..F1eQ7
^>^Z3CAbEZ/^ZNQ0Y^ZX@XXdDYN@U\SF,M\6-_)01e&Jff2=:J7M:@BMeRBb^I#L
<MAUfcEG-OO>4#8CU;+5OZ>(_OUMFN.-A(cg+?>#Y7^T(MZ(K\.<Q>PO+B;I<YUa
6WBLF@)_T\9BJ4Q/@ZI=RWcF@[;QXX2=(LRI;79[e3XB7Z2N2&Xf-b3fd/?(NE_U
aU&U[ZEe+;=WN=(e(aSKC7gPQ/4=7,GcIUZ,HOSd<A35]IMG;UE1=f&@U=20D0gB
:fG51f(1@Bf=AEUUgA,[0Uc9OD?VO+(@RDWGGX@c<SaIQ(f6/1W7HI+^E#;Ca.+3
0I[&KVSSM6)7UdFH(MU111CESOPRN#,467P\AB5@UPMeXfQD-cH+=E1<S0SE&[D^
HZ?#c61]ZDCS7EH^a)U4SDSRAQ+W/UBb;?+;CN1D1U+TYC-NfQePCG1XJbccZKbC
I+.&QgS86Q5L?R\fc6__IPH1I91fWITDe[(ea=@-IQ\\C)2:&?RIUK++&6<[1XH0
f-W>?L)A06e@Z:[0:Y:-T&4b_O41+ZS#.S0:H_?Q24a7FY.LK[56I^JWEbf?M&M#
(M1aBHG7X7/T.[2Q_]F=2aa:_#<ZA9N0Y.GN84#]R@5+CM93VG8RP+:X+MCeFH(#
-;X)fPZa@bSUY]7LNga_NN46.Og<6^6QWfFV;@9J#cQ&dfaP/[d+69HZ4?;K8@(?
S3aHKMBDDV8GBN8:BC_J_7?4?O(]/?8CPH#]+g@#0+NQ5I+=LCB?8IG?9XcLN#@Y
VfU/_XdOEAF3J)<9U7RIB7(V;6)(9(Y:-H@9PfOa:^f[IZK-/5?;BPfHM18(F^_?
P4O?]GBG-FY/=<<f/FG?-:bHfZ6Z1X^MP_ZP&aaUO:d\[BL[-#3XX05.[L:?]Z(4
\YW>>2NI.R:YVF>#+J(e9LEHQ#7<U>4Wb/bP5ADA_F]<)JQCaZ&Pd40@54>9A+aN
f399LGL+fYQ8R<6I^)-WdSHY\@TPN)]?A+eXbN96IcgGMCH.AGN3[B,4Y_>UMeAa
CLdgVMYQ1>X^MJAJ^A>cSX&;0WXAeHGUW./2U#0d)9XWbNUW\G)f;cKA<8VEJ9BJ
MbJY3.?,147][#^S,+.ZV2c]S3=-6Z@HbbT]E(+-COT2(da;-GI#S7-B.AI?ON_O
g#.Mb2]AF__<=LgI(-+9G\HP[1T9M7@PQPY.0G>DDVEVNG[-D&IXAbf]9gLM6NE]
T-M6AV#)cFE#J;ZUB>WJb+MRW.^>eFCHNY&-\6\R&,A+ZOJ\8cVE]=V2a8D#R+]+
&D(cOXHT6?ZfX);&H2[b:V_9O#d(eB,\<?N0(50/9W-IgD6FbB@a]SNV]I#659(3
T8(([JN+A#1/f9;T6_gP/.ZPH?L_)DQKX,H,2PeV6_b^8[aJF,]MBCH@J)P6S(P8
=-YKN,EFWaLGBSFYgeJ_fKB+G+?>SEP^W&,Jf;?DSc7f++ZB[5P:7Tf],2-)gg?,
@/NT7V&_EeI7P@6dXgd?UeY1U(XPHU:L]db5/<JI<RFZ,<YY52YMf_QS7A1H.N[K
Gg>]YVGW:ae?KD10=:/]d3,DQQfQ?f.KdSKY11eFTU9fd;IU#E)W>DYSS;/--G77
82^L?\[3AL<GA\Y[6O?XZ)dM&ZH;6HI9(@1PKfUM_PV.BQ-.)=XCN<BSb.#\eTX,
[DQD-3WKL4a,:1E1>6R/@5BF(DH>364VR4bE&NO\1+a=[ID@fS-Me_\<T+M_FgS,
1URQ8ZE(L90DM[=5(F\&F(GX-PfUAg?cZC3#LOEWN<S#=eJG^fU^fd>#PNUATX,K
c-W]E:2^0DT:)7R<WW(;_:+>J0?D=W?:/d-Hg.b/7\f+.&:[@,Xf;W@#^aL[/Oa2
=#J)I]DLAaJ_f.XT]O1Qe<X#?XP)a3;<C8LgB2/KW^><9K,X82LHK[6F?.^[=T9Z
GS_H+.6+D[cbU@.>RLXB77K>I?OK2\FQ,/6IFT476b-AAPb]<a:I?HPZa6DQBXCF
f3ZY[8L\^RGM(Qd_JO_J?56QGOYT1ZS1M]V9&TcT_,cf_1@]+A(+>IJPB56ab7\+
4P_=f4P7EbgYHFcH^9f0UWAOM;M:;WR&39^=V:1Q/VM7>COS6?bfXLRc@cabV<45
;gJIIH6+N@-FePE/Zd3IT#YI-1_S+EedY&5:d9]:@JM<&^DU>]M,1F,+Hb:RL?P?
--G68SA8#Y2C9HP8+C>TB@6@8\CJ0R#9f?LOM_RH\SX2+ZEDR&_X0/SP@7UScR6C
agg.G>4MFAU.C4JKKZ:HK).<@M-L63B3S[[,L;MP3\-5AP@.H31.])<[88RPAZ3M
<H1464/BDT>@J?0F2T,XG@?bgPb&.^UQ\[NQC:8LYgA_(PZg#5JfbH0gSR/YJ3;B
<7LNgCAAPJTZ64W++SN=<9N,MB5)f8CIV&6:G/^,MgKa,0QHL<PHM:[fW4T[#6aS
72a\>&EAPF#2.89eAN_8_?G((#TNFKcR7(YbCXM3XcN/bR#AbdAUbVTODD(=I;Z6
fDK)FTE1?SF+aD?@B190.5?K9Z-9ARX]/OTb+CR7K^F+.O;cSUe^T@S)S?8/A)N#
W?YC1X9K]K^+D]XJ?d0Fg=dDO8E60OKH=>O@&1\3<DeYRfU3UZDLQ,3:VDdFOg#C
^7d3XQ>6?6)4U:UZ/AO2:I1XM)WROEDB1UC&gBbV56JE)FN,X7CEB/8/eHM@&]O6
<HND4[.4Z9HPP(>NE#5Z[G9N^6WNcVZ3f4MPA_(d^K>SOB02YL:ba6=:5(9)YBD;
]&/??=N1VJQ/?#TM-#P\\I#a=?ReIeQ4>@e_;]2KC7^a;^OR82=B+36ZOXHAZ(6g
f@JCF]@Cg?a:JYY,:]Q>,:)ZM8VSB,S4^2=2+fAP;ZPQ<L14c6>L8YZ>NX-XUB,&
C</8H5cL;H&#b80WZEGNPGL(#(TT:fC+E8f3,-KAWgdKALT,a,7CW7F.9?LD507Y
SXPXa(a\8C7=VTgEON[:>E3[;e<6]d>>;[:Q+APLg7[69WBId?6+/774K20-C2&G
,[ZN<H1P16^853&-?=G>e6LG9K4]P;&gRL;^])-H]?LG2].9B^\\&1?M(D(@L8FI
XfY4/(WZaG&Y9^#F@aB)OB7<KF&;[Y&928>]-94QGcg-=Z[&I3\04VNa:fD^SUGV
Cc:9BDIXMW8),5UJ#;QR.7@\6.Z<G1,CBAVb+>R1eTH5>8SHaSg=,B<a[CDEUZ/U
7+BLHQR0Q;e-23AXH)D(K&(.[-HU?\/a6-6c/D<.0.Ff[SUF<7Ob))7HeI<3PDeQ
S+1U/9<338aP#BY.e>JM]FKHd[)-0g/<Q?a5N<AH:d4<b8NFW:?_0L-9aRC_a]Ub
bcQ,\EA5,.JRg3@Q\OWEQgFW/ZdeFd7(dI=E.+^02_FUN9CP<[eaZ<;>)[MK\-_3
DI.R:0>DfF&H#IEGK;4?P:Y4d:;^4WdC,I8HC.G3,Ce@Sg[IFZRWS8]5R:eT\0IR
:HHJW^(I74d34H@;(K1H74;(BNMTbU)_3Qb<5CV,9gR7Q5I4\b&cU0RU?P3DT179
Y@bC+M]UZbcUN(M&ULZO/3=]aGBS\5g=aO564c[GHRfaF0)CEK6VMC?MN3Z,??\D
SI\U_P+Q>)QID]G_fEDNI_4D,[7fO_^/J7#]VBag.]1:#]dBLXPMQ4+M)292,H_g
0Z#;e\P1=[+dg:@MJ7[APgTK5GP&N@e+_>aIYMKOBBO3gSHagTDG(YB:adX((IXL
[/J<2\/dLL_E_-JY9?g;R6CceS^gKP7EEA\0X0>1E>@J\S87([<4d2(P#S-Y[5A,
E/,-JdB2(g\1K&6cR-)Q5#c(&3]3:RA)TT6gK/RGZ[_RLY-/Y#@]9#IF:8_]/U./
gRDcDGS((_D[7<dQ[&R2P8SH][RNSPaUQ]-^0]OD8W0A[JEe+^N>]&:BJ80T(4OD
H#G[-];S_16K,?L.,GXb;WCSLO;SNIgQQSJ1U\Rg+BPQA;[7(3;V4&9P:bSMZZZB
IM9\3E50VB3(/PS(,,.#f3YSW9)8cFdT2K,;PIHb^>0[YdA1X0+./bg80UNJ<SW(
I\B,[OALCb>.)>A@WVG-YZA].RYA?,Q7S187GD#3-5A<F:,^N<8-:&B/=-[a2;.9
>\:U<?Ne_\F&W3PF^8DEbg4d^(51.CDBT;<d04cL8.><S#;H6dM,PafZF@),/4)Z
C/(@g#g,+\D.ON2aXbZg@\Je^:KMRU8d\A#.NRR1GJM,<\(RN50_^Ae5e?bV4NAW
#RQAA^GJFF.4_]U4_:3A6>_SF[]@W0\Qf?ac=JL+UJH41DZIPA]\\.N54WWTF6,(
S)1S#(\01C&31NC](0[>?P>cOXEXYIZd=\-#TIEY1UDD>UY]NgY]A_0^aa:&<+G\
_E4f3.00U=,_&Z^6@H,K+5>5ZPUJSFeN3Z4I,Oba0/OT^O8HA0)^6c^/(Q1\Yg#J
C&eWKJ-?@W;VL8/X>0SD/IaQeH2(1+:2RGC@^MI&U&a>LJAAc6E8EEX2Ua[7&<0L
T-g7E^D#WPa.g^W&@a<4^)B.TbgUEgBQ.^d=E5]&U)4B2&8(e1g7X,g:aVGV<O5^
,<?Q/T&R.1&B9SXM,\51-?-Rg^],+O@LAM+U4=YK_IZfT,,C\XgIC1:6L\@XN[:D
E&E<VgCb\P)7C1NbC&Q-(^QE_QWEHVCNRU]X7YXF@cL17SeU^:T#a+E+2S/N:7\9
SE@./+MKCN9RZe;8f=+dU<8>=K@GX[Z&e:VbUQ^8])[N<D+H9<.[Eg@ZCb?YI)7@
@D(X,.e_5RP/AA7:+Ce2RW0a(]+9[ZTaV6I?DBTJOZ-[IIF_D=bP=AMgU+g?;,J<
PRZFbD&ENW0(SHTN[,VS5VOWS@]>b:KB:7NLWH>_9eKR[J958KB>&9W=Gd(7YZgY
6I9BFTfdF;IXY/77/\]97V]CXe[(X1-EMAYT:GFW4?Y#IT:@XOKBMG[7?QYHM;XY
=&4K0Q(,Ta2<CDPTN&SJc6-&_IB@<fR@B]/[N;K_cWX>&J@6a\8^&EL3TAEU9?6L
<L+H5>M=+I;cF5B\#50f@fE(a8LJdAQFU>F:86Cg/.HG=f??]e>>?Z_#>:#Y9PWJ
&4VQXAZZF94_K1O[]NfWO++,5ZO:67g5IR.P3PCFH];3(:<&^>WZNOA?MZZZ(W:.
[TL,fVZH9b1)/<C9\de:O\#fa<355]BfVNEb?12L2J2<6;CQGR\H<]=767-M.&75
>]6+82I(@G\PBaB9>\B_O<b0N9TK-8B22,<\6TFc227JX#N:F8([_;==;E.DA.Ea
\V97D[A610E0[]f9AJ-Z=Z-F)bKe<+/(Qe3U4+X9G2Z)SKF@6^F<-A[KOFe5JY0;
61^.R9F0B4c6NTF0Ib\.YbPVI3O^<?#W+;X/fA=R)LH[SGZ&NgHWfaPR;0<@U.P@
Sb=86K<dN=&-L4.)?]3+(^J#NP.^JgSH7<]4530gPBCK_;5b/-^XHA>5X/ACDLPT
4U;&^QK(CP2Qa8J3][ZB1,e-#cYWBI4Sg9SC>[TU,8O@^,Z>GY4KW:OgM8VSg0;N
bDCN+I6AdB1(9Y0cc3/>O6f4adeNY+W2E\)4;52^R8#8&W9GS;BEUGf3&cObKFR>
RQ,P_<^?E]OZ5_R+EMP8&a4H:V13=&FQB9Y-,]fP-B(9:GH1,g(2ZS])-WY[2S)H
?+^eWLG;6@O:_2IUaK,N=/>>38I?5RWM->KVHO4:c;40;U-OH_,XB4H+d\+2QaT<
GcD5EC\G\UYTQd//QPY\eR_2[COB6OPQN\I;=E>9WKJKXFN;IH=1N9f#<(T4:),B
:F]G;:=@LUaUP7CdDX.ICCA=X)J[+OaZ-7(?=\[DO;7X/J8F2PNZI&c(BXd1Yd3C
DNZL[[V00^D8YO33].#LOMM?Y6Y@d_+bY4)CS]b#d@4O1:7Ag[Q4UHP4P^1KQB0J
+,f2gAL9(TL.TdB-L1bIX6R2g6</616A1RB):;>6OE[N;Ue4K_<E;J56O+XfEDV@
gSG;B-W^ZBC+F@H5AeBX9&26S3NK7O:YNdWN2L^&5TQ\L.M;NT)MSRfH@>\,_DB^
;#_>+1CMa1O70JY40+UffGJZRR3@(DX0S>L9=MRA.06@\<RX-HaZdCK=W3SG>eg0
c,JG;N\4@=65U2?+7ZI.BHVX4X(PF?WOa^+ULEfaVcK/X<g6UL=VW>Z]aN_FcI6b
F4K</MGST3U28CZafK#L[K6ML.S7F^3[\-V^G;?D@YB4f1#N]=C:1,ZdTF8<H1/<
2>B2-f7AX,LQ:+U^F2>OEA+\7?<3J_A9[AUQbJ-Y&bg_?]/H/>9d1^A)@7ENE4LG
QF5Oa:c#P8GX2V\B5,IIF[)@]5ec@.4cE<7Y(OKQ6VSdFYGEXMKbPDS5cS6_R2Ga
G86Q=2+[0;Ka0a-@aI>S_A4g&K\:I)e5#gI5&82>I6WR:<S2Vg84V#@1=H@1&Ng)
F^[O<0I(E6JC#E-&HA]JM,D@E_5)aBc138>+.:M]a)Y994?AZF<4>N7^RAN3C7?#
+O)J0=3[ADEcTORbWUbc)J4]6Gg/7G_,3-8>4&YM:QU7DHXJBE:Be4[=,aag\dgc
T3.[\W0GT2c\(Y]CWSSMPde^e:.]+:E2b/G3Iff0GY.T2GEQ-K.R[<BX&TgJL7,K
YJ7]5SW:/THAe0g^B7H^DG^FWS)OQ6\9JU4XHW.RYT/:SW(4f(<(KW,=O;QcZ:M6
a_>a/bW#CPPRS8>Z)0G:\@CV<0bVUH7UTGeO&5g[D;-Y8J#b3Xb)G0O2)3MaI6+8
@/-CdNE+_9@.Z@Eg\+>URE8T7>a/J&/Pe&;N+L//^L>g4JEWfc_)<a-,94dL)e1F
KZ<)&718dMY7fePWHXa6=ZT6O<<)>8-1XUR_T1#Z\f@LCL+)]=&2#5VHLdU@A=0#
.CdUFI3Q.XPOea96K=TGAQ[-WF@H]b&_IcF3(V?1b4]:ZJ6?:3KT&SZBILBgY@S0
?@ORRZ<G1).X5V4+c=UQ@\.6)\T?MZ+/XYK8b[OV19\c>::<6\<F510VI+=E9O)6
^>AE9++(XgcVC<&e@WW5(X0:Z?&&PJ_E>.F=96aR2E2TcaVA#DUBO2[&^QBC2Y/C
-[,=:b[ID+50NC5aE80Q4K7dV2>L#T2:OOg=8Q50c,+_06E^f]V)5VTX3+^ZZ>B/
.60-U\g3F7T?Bd.Ud#/QT),OgQf9#UR=b\7L_L&07@\EI9.8AH_Kg:WD2K(8N,Qa
812A&4a8I\a/-(P<S1W^41Ea<F=eF;0^Q9HPF:2LNfIB1,TWUfP\N(F5JR+D4ENU
ZA25DL_3;9ZR?<ca.+8Z8\28XF6AR_TGN3?-SID](P\30-Y/@X\6[D>#e1#GVF9W
1XGL:Z\@6)>bRUU(YR1JW82?)R86/Hac.>UCX+L6DNdP&H4RX2g=b&f[M@?+7egg
,H-S01P]eHgadF(>P)f#ATfX5PA-&V?D.E5aeHO.c=M1ge\2N/_(Pc;IR,[+#@(>
)X)K(.SY7EKF[09Y(W2)5T?Hb(ffK783WX+eLCY&.+XEF5dJ#@Z\+X+W.&g.G6LI
TJaQ#-?B.>S]=#Z]0N[=b:F,GD1_R.K6^4QbW&@fWY+>[&f=ECYKVJS6YLDQ]T=C
Td/^gG8I:Ue-T=]Ob(Ec?302g3eWH;TTX/dR#B1B6^;<X9#F?AG45b,Ba^Z94NeK
IB>fYP6dL):F1XUS?5FeX8I_5DcG<&CL;&R21C12L&P@RBP&GJIS(EWeKEY3fAeA
FP9KI:H;4P-Y.AZZaJN..IJYX6Z/@T@TdARb,]98].5,?F2TWVc=g-H2I=DMXd)9
X^f>PW[fMQWVD-Q8#3Z@H@b_?_I?#V&U7>:]-)BNXBc=-:]Vg=R_g;K,1]?.0_-9
L&d#dE[&^H^)-?<A/=#KY^O]>c9<]b@@F=V?GNF5BAG+70WI6>2=LMQ(b@,Rd#Y/
5g/)E?,K?W?ZS_[&93[2>+HLM#4+K8Cef8(M_HX12OM9N[EEKANA4KH:fHZ]Q767
7#,RL1<,g;,+S25.;7,@OH)O&(H0X,W?DH=-]\],^ZJ4B[5OT[FOc8?UT[&c;T>D
TD1QHDd<136]5cSa;0VeC5cGOa&<fZI3USXDSX@ZedR<=8_(C>A^O1;/AZ68JdUB
MGM1E5f&-F^O.T/^7X[RaBc4IAg^fLRU0O7AW3&P@30\cQ;#IR8H0FLSZQ#8bQ]5
8&GJ;+KY&PVKW\4A-@2F[G0)^I6#bfZbY^@@YB@_:,B\XIO9;D_8\DU6]e]d&f/_
]QXS5Qa),X/IYNRM>Q)8.^]<E3&^\T(Hg2H2^eW1HY8).b8R(g#e=T8=gUWHOT3&
^HM).80IMUd@J[&[@<QR6If4Z]VD&IF+^,=f[F_MV^/g_3#CT>8ZE19G0E;]PEIN
6>0PSL7BcG)F-=BPg[<2A=+@XSNFA6eSe\G4BBF.TLIWPKNQae>SB^EaS8YI1N\dU$
`endprotected
  
function void svt_ahb_system_configuration::pre_randomize ();
`protected
]B35657Oc0.=82:>E_<MZC1X(F0XK,J:bEOa82EGA#Rf43PD>E_g1)Nd3\E7MA#@
?DYRZB6SZ0MZ:29LR]HJ:(/]0(3GfL[56_1R=fe_8EBC?-[e?;;dFE3Y>4?2MZ&H
M:BYF91a\.\c#f5V_R[^TSAOJ)_6EG5/Z4UB/4#7XWE<=#I-<Y&R.e^04I/:\CVQ
SWRg#3\EDL5_1,\c]EX9K4[:>AK8[#UD4(#Fe+]Mc\fE\5A.Y:eVfVLPY[4:4[Lf
UHJ^J2T/:Q,dFFLD:K708>3#GLQ1I>01MBJad(E<aPa]eJ:XDT])+U#2##^3d[0L
&COW>@BB=4=.D2RGWZ&NZJDf^);?Uc^PZf^YL6]+OS/V)10_O;[:aR?XB+^1(#Mg
IV/[MT@b@a0\26[7H_WD6VJ.Tf-gSPeX:$
`endprotected

endfunction: pre_randomize
//vcs_vip_protect
`protected
E73=e=FL^;JO),g+3K_0E,b(NB,E7-J&Yg?GY7W?1O;I>HFJ\d:N((f_]VHUI_LO
,)V9PaZ;cK&@dA=7X2Y>_(fbPA\f9Y2@/&ONTH96AS_T=_2GR.MXTXbeYLP]Bg=-
:E:<+3&Y35Wb8\g@eI,>1?5K4@E6LbAO)P6XG1RG0@KMc+1Z8_e8YEXF(]_Z^3c#
SX<^)M_+4Q49V[)gM3BO^g]TEHVIJWR.MH\L[1g5]9[TdCI+:4AgQ__L2;)3F[FL
:<)=]__>X,[X:SV,&WI\=^c@;Ea^=a(gc+fAd^[+7_c\WLH3/[NaHQ?_S1Ebg27(
2L+0XJ4Z5:0^:W;(5?g.cIJO4FOCMb(W6KgfV1?/1fFA=<,>WYHD;]Q=(B:6PF^C
S1(e,:e)T1+XKD;WG6aKSL,][K8BdUBEN1[e(b4LK()f/==Le@_:OJLT6<:[c-6+
Q79:NP^Q>D)<<fg3d09(8./Z9#VB36BA00^#e,O.M#I#LO3B8>+]3;0F4A+_<HNX
[N4@@&]3&V_YEdfY4GR-P4VVQU434&.=RKJ_U<[877_Z7C.gRHXJ#9Gcd>G-_VI@
a9\/V/5(a,W1b2P21^OQ\;)/77X^=g:f5P@DI0A56.X1G-g[YP6F;YdEePfI34;7
-.HK,PPLbBWE471MMd>Rb:4:F\\RBRP0eCL;D@OdXZOOeB3fRH\#/1.63+S7CYT,
f[=2+CLD=ae/T+S?T8NXS>]6cB7=d6[(L6dd620]:YGX/[SAV)e1^]a;X=8.?e?I
[E^cX<ED@fU^TQ):[DO@ZQ]=3CR5IYZ^<Tb3_^9?UCSe(>4YJUC>/+0+@Bc^6<NH
X1W^(ON<g]W^B9QJ39?)/@bOZ4<+S)2<>WgZSS==N&5V&DD/G44a1^<TR[T_HFIB
9##bP17c7Y67\F)fSJX<)P0c.eNgB[Z#f=Gd4F2U+W2M)/d,T6C0Cbe_\@6#Q.(.
-B(XYdTY^VER>APaA<WP.Nef(F8D^X5)+&.VPX5aAVA5TIF((KSMU\F#X8:.BCg7
(RaD;MZaO+>JV,UFD9V3FI2E=3\^L#P)&.b;4^][fN/<&K9E#1N^H82aK(,6ZLV2
NGHTb^OBe#F2E,VR5Z2Z5^\>Pe5=H^^O>MGR+XE6ScH?C@:(dS?REUb)ZGg&<8IU
E>EWRL-H:?#3c=Qe0DD)bW0d-)Z5Vad7B+\4G2cV2TY\&CG>:(LQ[6(W<0ND#JM=
Q8FQ(+Kc,=aBWP9E;bBec7NOE.#P,@a[Z=SF9ObSDc)#@;=(I;C[HD&(8b<-J<,L
LTF3[C#C3c[K]F2NBT;ffM;8M.<Z2ga1P..S1/Kff&)7]g\/G;gQgZ?.:]ZXedU#
ITJD-a;3)2(d#&1C9-)H,@d@2:,DZSEI;bZOG,FW<^;NVZ?>Sg8De^,)BO:AX<eD
]1ePZg0F\c^^]P\I0SZDe1(C^T(7NNMR81g/M&BA;bbC&;a&/=(cBO,]2R.74M<M
67<9Zg7TLUEf+M[@JgeI9?IR7#/02M;)\Be\b5M1391))W1I=?<cICH\YGL91e^\
.K&F<^.:/=.B(X32-ML4&cN^T-O5\4X_1:+>&TU3T8b&XXCVRCJJEa#D0PbFe0>:
&GPW\P_M\+N)0g_EZ.0=2AN?&I1O4B6.fe],D6_e&@SUfRHYF]J)NSD=b;R#DN^;
V.7fI7P\H>/]b.LdOV4-DP:_)[Ba[E5TNd(fg[=/MR>&\73X144-c>&N?E0gR9K.
MRJWZY,:g0SK>RO>>HOAOQ\_-&\C:-XPNWRRO4^;X52eW\M@?U3Ae2]cg;Vb+g^7
_]R[eV7KRX>208,NA861XPd\PF,(A&X;;25_^1&EOdQ6&D?@6?aGaL)<)6dc7?Hb
;c?ZK3._7I-91CG1=0f4\6FL07B_a]dV=,,K<>C&07AA;D[2f]IA1g1J&5c8.XPC
LGIa>&RR5EMb1\,E[+ID(IDRYY4Gg?3d\51T[L.KO;,&b+3gW#[NVE^EMaVSH(CG
RD1HcZ/GZF[e;HT[c;6#</,dg>]A,cZ4(8f_/92A@CXg/Zf6;K<IO\J5/371;Z;T
3-Qg&G5b\B4,,K,,G[U=eK:SK&dPM6Y[L;ITe]W<[O-D,6;_/6MB349+7GAYH;9T
7V=M-<^N1+B8g2R.:(<EN5C?ZfRSc3b?QQaZ<#17G/4e-F:_>g^TQ?0FEScUeR9c
W4.eJ.YcR1#gTeb\Q=GJ6eL,DNP3)ZJ0EELV7I_Q_[/IHa(/#L,[Z4)-ATEUOT#L
-cD9([\H:R0J=1QBebYWaBX:a&R3+D6&.F)M[6#;(7VYKQG_,.bPE:(BR1e6.L2b
Wdg\Ce)8=;T/=68f8Ga;BJXWgDC_6A/(UfK,CEdE,871M#=J(OgAXbOb8.RY^D@)
g0f/7@[K\V4e)F<30/AIE\_V;,Y31MP5@.TK.+EUg0B6.+]gB-f\e[AW^QZ<Pe1?
ZJ)K^(DD;A]WZ6HI#a?R3)0N-6^c3GgL1R/3>,W=5d/IC5+Hc,IW//[Vc@>gT/<5
68JRaM@NMBF&\1@g]K1dIFUc5Q_&I>a(YfKM)UQA?aTEUXAB_9Y3a()VYRTId;YB
.2U3e9C0TFZ)84ge>,UdA[ZGRc?Rb.C.83^5cb34F&NTJ5,?9^;1\Q;a,6I#8>a^
;;7f&-2CM=:1]/?5B@=ZZG1K2d+]Ya0?;7S1(f;b\;]QQ),9B@e?e;3M][\N38JJ
>f#&0AE[4GMA]2CNTK7U?\-PTPICB.COEM,HJ>/^-7CJS[#TD5PM@(c2=-WRSba@
[]J0WR9B>9U[B#;.BW_7#6Q(HD.\SPS]BTBNbfe\7e+B#M1T/34>?^aT89]]ZYJO
e58AG-^Q;4@/FLP5@GHC[9d[_Va;E3&-78cS+7H:I+:9T8NVB_#bK)ZLC98Pg^B=
ZM]@^^4NRUAePRKVAW:]LX.QM#S/IPCSF_;#UX7RWOcPdZG@W_-Y;1_]FT^d;&]3
N=.7;=U,C+MX7A0Y&6DQ4Y#0c-cf\27^QQPN;eXY:d72K=2gO7c3)?V(gL:)UE:+
NDSA=5ER5g487J.b.&5NO9I7QFV00L)XK)H8?D\b>eN[L4>d#WG0G4>fK<g0@gX\
MS>Y]SXP]8TageD3]E8&0/WB<58VPV@SJea5KN?X3eQI94,?[Z9UPBC2_U@S),(@
,d+Gb.gc?YdEW]PHLDW2)cMd6UK3[TF2(P&X61]2ZJB#Hd&CPY(T5M>(<@B@]\+e
3Ue^-.)d6]6]cg).J+N<VC&P>JfOa?cSD-Q>]FBN8&]2?aReFdTRMKTTG,^.A<3-
&T(QZc0#5TFD:J/YX1=8E]Ib6cdFQ2^dZW19)Ic:M1W;dSed@(GAU6D3G-L)afG\
f-FgcS;;I3-dWg.DGF?M)>Y^c;g@a>HJ&;1M7IZBMAFQ):SIS6;c3cabC-(/NXWI
[0ZU6_:NH]</\WFHa>g,-+b2Cd(>D+;BgGe]eQ&HIXf0(NZ-2Y7de>C2IXGZ30f<
]R/E#Gc\RZ^Jg8_gNEBE4R(Y]I)dafSTgg9Ec<g)&E/PA,=.1W[-8_T6+aONFDZ6
2\ZO&0HTE5&J^I^(68G,=,&3CMaR[9dgP)JS@]_)&2JeHe##d6=1<1;POS,)#3>L
]&?6T\OT+fV-][7@SQ6,dE_3AQA#43;b.[4\.EK,d>Q78M>?U)VZ:(,M..\4+gFI
8T>b.)>=A^=]fBTT9eJbB>XIB;dRLcgF7G7#C@8VXH0HVF7;D.JFU-?Y0\-aDDTB
TDbf0BDeN>U:E@<d.VDC1Kc,0BOVG.5DH>I>/6F4XLZ-e(;18+F.W92#@2>;5M[@
L^D[K&g=I=)AeP;DS#(NR_00MQYJc,#\2ZO@A3UbLZ0R2=>RB6BWRE\E3#=EaVK=
DFK<,S_Ff5ad1KT>g[JMcQF1cF+7_I(6OT()2JgD7KYPb>Rga2;(E.<-0-4-)?-;
_XD#4Uf6/QKS&F4G-TSK?[b#63JBRH_b4^&C+14Pd#V.9bKb3264b-b+RZ3L7@gN
0;&+fR:N?RS\=OJMU8WAf@;4VQ1O()A=QUGD<aL_63f<S7[Tc5==@S+(&TVSKQS0
73B444K;_A&.;-\BTDI:17X;5^&(F[>-LO::RdIa@9,g:_Y-GBcf<F7da(YX.1d(
EEY@9Q9b\^+6-^g6H<F3C]&<JYg;N_1Y7Y436\)#d2/B-WBNdY]]S3G/)[3SHZB+
UKBPGXEFc2;VQF0_O(8DAf6S:+#IPDM&;b#CL#^##Sb9&>6R1PO]XEc=0N9AMSe&
XAgVBLMdXa@6g0Q=eURO46;?OY#f3+N2cdVfD/4-_;RCF4K,#S3Y<g[],1AbbPac
G(geTT\<SP[L_J>@b:&8A28@_1P13UGQTI8(N;PCVS9B(RT?#A,THBT#<\;c>+8X
ee3.POVBA^#f#]-7=-IL+LGeQ1c5f&7:fBBXP4_3#aG?S/a_b^^KY=Re[-K(34J(
12V[_:_]>W,:7K9NJ-HUAWBXe\W;gP[__5?W^EA(PS7T6VeJHg9=W8TOZ?EC.T>.
e58Y(+N+#4VRP[KC+XePeD>D.1(A@=ZB5BV/Ubb)IM<gcO])1LGFEOWJe+G=d;:_
MbX)>V];ZKC(cHTC.9P].::A2I_IS]AS/cKKaJa,L,EPc(Y>a][][bQAPAdCeN\<
\8_R@d)Z,BIe9F3X6#M9;Z@9Z+#863ANVX742J@5KOWP&+ZW_L#e-]A?_Z?SK)OQ
UQB^JU0/W,DRcHgKM4<TKXD@?fK>>)8:D#4[7,ec3g8:/J\P7G9-T3#T1FPAT/C@
:BZ4R>\3UY&/G-0:NSdK)KfKca)0[4[1<,cGf9OG\.,9.JVV+=1TJEf\C2O1SF9D
M#c=_?FI56dSH7/GbLN][14C.@RMd@5]WF+J4W7>Q#c3:<JA3+Ee)@Y6:BbPP6eS
HAUF]5cfe9IYc#I(C\c@@\Xe><cIH(^DI6\\cVJ:ZBF9eLgOBf7Y?VZ]XI4/a:b7
T&)0.>b9_EL4G&B,c+Ea.EbKX[2UCN1L/5U]b;Yb.VR=-,72<R<8\/.#eHI9)+7L
M#BFYVWJ\I(]7<MWL=J>MTcd2aZ6Q:Vb;HFC=\8TcL2W1,^A[9GUM280O=Zb^\6b
#0.3.C@=8=N1Se=d/>7-\ESdB&J+#gH=[J.W+^5^[Z&:9(]8W\E2CE-6.&#_9CaJ
7a<UL(\OXa4=L^X.XAM;[5#0^)MCg1Vge-CZgS&SB@GJ8HX;)V]=\X>X>FW9L4^U
bOJGFQ?\OMC>.[.;2\+JW@Z8CE,US83Rb6M\CB[.J+A\QBQ(OeQf\79&WM[Wd??L
I_2cB&6BTP,E9cL2N@GG)VC5@@e0:7IMXPCB;S9cB)TN#:5_8\1LL[]HRJ03OOdb
N1VBJf;-e@8M:_,M)EZ?W;U:^?>R<;NZ?>Fe5E&=YNR1S:&NE=V6WFbT#faN4ee+
(/1-HUC;X3<5SJ:bC-T6P@?3&(7EE-G8E<bPeG=B1YF)^G8-P86-L:N9//7dcBRJ
XH71;MMBA@_@E2^aR:]bK,PRd_F_[4AR,&OV1cD_.FP8_^ML4>(+CDTdfWdL]KEP
R7Y^NAcNC;M2=K^<9_+J;\=fCZ]2F_,?Y9+AAUVH3_f1N9aQO,H#++E[9T[&;+6/
;<?K15LF@AdDS40gG>09VLMMXTdM8Ae6JXSCWMAdU)CH_1VF-3A[[WMFOJ@d&2,Z
<c&-OK3(1ZVH<PTG=AB?gYg_0,bd=#XI:&.<1+[4f\5MV.c<WOZ0R^d0M3\d(HN:
d.gE:?T>EP-Y&,SH<GR_00Rc,I(4:R\_GL1Y?]^gB[=_(@TC_IVI,b8P;)><7HV,
&7DDb<;#OE=F(&[)KE6NXa-+?/NUKM2UWF-K>/76gc4,bV.OEd,WRXS1KUW>+TPG
31\AE0FJEAQLYG1c?Z(:c/=MGb\/(VZA/QVd@c7e2I1#,(USJ7>#].5W&/FN;9E0
@E:<Ke5D8E@X1O;e=&\O@L1N?21.5X4W=.VO.5aW@F0+K8\5ePR<Q_WP&0-:TTBJ
+XMP7DLO<AFd9]+5OR;@F-RYSFV<YV36>1-E0OSId+gfS(>@;c77.C3ONRZ>UQN-
SCEOC^cQIGFe#IFQ?,FSec.bM=/XD\K^_:[E@a5:_)+OS<(VN9[J7XY>_cSd^.P>
cEK+5)XV>@LZ[T/9L7)M^ECX]\d1@g-RG.?e+P,aMHF2MULOb4_#CS;\=^]ABbZ8
]@3SL[5U3=aYF;ZHB]Z1T1#LBJMAICZWXgLEOFB9)C3RG5J,]cV8[TTe(4N]WgGb
N<@9?CZQNSd&VG93ZG[Fg?>[-8[1fJ&9VR/2)3FO@HTQDU;g,d&J[fWF]I_:/B60
C]O1_9J5Q[^-dg+M?cL:@(X7/=5X?2]C?OL1H:H>6ZbMV:4A<Z]DN09HgH;d]B\)
NGCX#F<@3#MLN\\U7#3.KZURHGT1<L&<?/7LLLLRVX&JS3c[B7Y0JRHHVYgJHX8O
=C2?B&W/L+GUI4SG3dR3FZ=)Ma,<-d\BYV5]&WT=8)]21X>/_G]b]D.X.<SE>Te)
g>,=+/D4S]JT_fa)<LT)7]>;C1+Q-VIC+dTR&AE)<W?Ob)_S4IX;3=I8_M+&Q62&
-9bAGWd1P#]=E_TS6)b?&IQfVRaTJZP[064<YfBYfW(6U4KV-5ONgcKYDHB[3;@@
2G^:I[;98VN40._g[;-T/#A/Ub16)AWK&@14P[(bc9Hb9CUK?QgF4LPJX_&d2+PL
84ab962^[(bW(ORZ2)[fXBOe6GHXf70Mbe-Ee49fg/:I[8\FdJ2/-eEMIOe8CQTW
(8:6b>^fK(Cf#+#QdV#=G:a:V6d3Qe?_]cK3<55QW^C7.MIc2YJg7-SNSMDCR.UZ
QFb.A?.c@&1b7K+YB5OgO8E<4LLT4B9RHW;_/6BLP52YBb67#YZ+R#EeEA@+DcN[
Ve]c,N&Hf:OY>dDYBc^8NQW-V40;gIcAf7BZ2D)eO6SBP?=5;40_WBD66)IQELOJ
@11<:W]H8AQ,QUW?9CNb42+@B));D]UZ.81@XKB9#X(5Zd52@5?8Q\8<K#2\G8PT
-]SYd2?M_c6TZ9(;PK<J^\K3C5g^#X)P8/.SZ&L_V#EJBK-af8;2?J,T3J4+A+XG
+D71C<O@dEEc+_#GS3I:e?B>d.Vf43/T#C<\O8T(F>47b;6aF5.F:)]N>-Jbb1CW
L8#^c?]U].76]G&eH[7ZOM-RJP.D&@D(8/,BHLQIbZ7F[:LR+9UQEI7E)PTa^Zbf
dH>45[[+2c,b@g+&RJbeeYMb9=&4PY,UFTN\4>=Q96+^c)dG68#.5FN)J0_/W\GA
\Ib-5EZeOC<eJF5K&8ZP>IDP84S\L1U@.Fc.YdNO)D/VAgK;bV:7-OYQgEaA.PN1
&H=RSU)OT8R9?D,=dI9g?.HAg&?9eE/g,P^dMC#B9EL;=LJJ5NYb;(ZW-R0BU0U\
<CU_\aN]>C_/(CVD=\abA&=bR&W]=XA:BBfIacFC/V01fTZfQ4IA:g8T[K=+8OLd
75>X(^&[V2#)\W[>#:M..Ac/R<BM;JIg.<N2-B8F+_A^1,0-^2\Pbc&M9=g1>:2T
D=e(,Cb1eZ8127(/)@@Z[^8[A0dY3_fXHdMe0I&bD)XHCT,F:)J6E\FDFNaH8OBf
YVS)5EKN:W?.O6:XCab\/UE@5?dYS&LP3gYSX71a[ZYQ?V22]24]9K><5-2>HIbZ
O/N10#e>7\?69+^#>^LK8RR:MK9VB2#IDP2<1A:4f^JMVV_6G]P_U+Q_HPHJ^H&B
HOdE)/L(Qc+Y4D3:2CLT>f>>A(<?P#:1X_L6QTTBMc3Y>a1O;7ACE/.=N1RR[>-d
7FLN?a3e;c<0)f5cA@aK:+D0Y@VVUL#PYF,5&E[?ZK[=L,68?Z.>45JT.Z>IE->W
>a4J^a<FQCHU,fcCaM&4ZGMIfQTV9KWP8U)O)ADN,L)8JDUG]<:G1>.W<g=)+.,]
),Yde5;603<4WU,+8ONZTc)&KA\Sg&]=H;-/)VH9XZC)D5D/Mcd1?Fe<T<K)E+>A
]>?ZP8V8b?=&)_9eP18[[40bT)cATedJEHf6#=(O^=9ILeI6<1g)[@.4&Z9:C9[a
N[,E@Y^0.=N>g4]SLEbO9:?<KYQZ=2=^?QA84#A<[Db?\\@D/NRf5V.BG>^TXXE?
fRd4#GMY/EM2MLMfL?O-L2N^&DIM9.XcR1^gA=3EN1>K(f/5c66UY?]9fL9L8Z,,
C/:94Vb=I4,D9fgD]M-02FA=XW3+G,Pc#0AL)cNQDcf6<2WWGU6OMJF^5S6N]574
(HBBa?-J]^YfN,GW_PF^DA)&BXaU3E\V=AM>]^K+?C5AB)PVEV7a92[\<X+F=OU2
A94/A>YG@QJ7Xe&W5UNc_/Rd-4+U2A62\5B8\F/>M[&:0-5BfdWP;W.L:#fCP)XR
)F+3^]]8K_2=:?+HJbe2MF9\S>TY+V&c+5_[X-/&6X(9SIgRX91+b@P&PG6U/P]&
&^eB=SIM/9[MGV-S];;DeMYB26c[D7MTS0))B9F9LB3d:^C#,4aS=eL)6Dc8Q+.K
O_\.X?OdIK]H7&54=V;WVGD&SP33\YU_Ka<1\XGb^5BbDZ??WMS];W8#R<;,?Q@?
f)MQTI+OUGf7<[[R(gc+JA6UK9[@U0c8#0?da5N00g.T1aLEfPS\cT>eCUeeD013
Lf=H5/1SZJF<)=Y.10L,]ITeO91g62A8(F72=b]fb>+gAb+I&F/(4MJ;=0c7f)K)
e5#^GPc<R]VLfY/+\\<OP)I1KF:H;CDF)]<UU6P7JH>Z0M>A;]fg]K5\C^AKdagP
]PS(c;G6b3_ZKJL9DZf68Q;RE+H;Q^;F1a6U]06Zg]>.)61b+X+XKLBKS=a_1DI7
STS+b/aKTf&da&X4+[\H3V,BEc35IR_Da5NUGXC90P]:3BdA@@JWTDP.LH>-aSRe
[)C09Uca_8LQ(1)C&,&^4S:bFY-GCC^<AbT928de/+0UfaMCM?;)47;>QV7<.R[4
,MWS(XW0X04^55QFLDCVgP)dP@;fLd.b#TI^3OW_^=TgYQ6MR4=U6R66H604UG=F
=3M_9O,:)\VV7fX_243>a:S\,5fUW#\OAG+2Sa7NG2d99PW(fX\KP@+TUYa^<=H^
XP3ScH1BBF8f?<DBOH^-J(46^Z(GHK=W>e;O:<Ld]3?YD3cY.@3a-FL=4fT)S-:-
>ZKC_gd2ZM(RaJPeBbW8D.(-X6af?eX>.S85&=b0@7:#)6B<(#Z#9)WY2+gP5Z&E
AT72)P=L&K6g4S<5TSD#_1WPbeB/TG:+3K_2(DMGec,D;>GMFV]E+(DVPPg3=N-K
YO0Q&F+.Y)881(\93G]&3-QF)Wg.1:H:84D,K]L1?8F7e:G7RbX7gCFD?W36=\bL
1W4R&]B#4N/Z5a#PKDd-fT&KUF:#Z0f8#09+&:1CXCX<];;d.;bE76fZ)D.W_eU<
AZ3?21Y4N/_PZZXE+ALQTEHV+R=U?#\2RZ[Y8eD>@G2\[5K8^-1L2+U0OUCXd>)[
f(SH^\86RBA.1?FFFceZT,I3H[S@]3>bC^2]1eLKI>Y-C0N2VX?geGe=Y<Pd6(]e
YPgW4E>-UGc(YD[P,@0OBG[KHMdXZA1_227K+2=/cN;3G2<ZV1d;N+U)8>T+4(C?
dH8,&LO-II@6<#(A80OHGfE>b)IPFJdb(.c64Ic(L,?O-MA\_<L;f3[L6d_+\1fG
@aXU?8RRTK-L(MCT.72MdKOR-e?a?F+3@fKfcUI@AeT<D6D^8MNVS;UBD5Ib,YN6
2/W72&<FS&.[6H8d9Q(\T9MF869R.If]a=]4&Zb7]NZXH]gT?Qb+=MdHSBT;ES)7
eY6OgS2#OB;.8K<?8R.e[)</V6]dB)IW=HX889V?<Y>;);].:D+g.dT_>4SQYd?6
Fg(8/,3C2<d(Lgg=<FY2SWK^VVZT7b=R#L/Ve7XgfOVA#LMAN=FLIa(b<#Q[^PW[
,d)_cF6W88237&@eY-5BNG_[HG6A,6SJg.+8^dbPYcCA8-g5HPLFg=CVeR/-^g,V
X8Kf?4=Z+M#-F[5,]G94@g5)J6&aWD-.+P<\SW1H^9HeJ7U^B=V9KN48-a\Eeb@-
NGI(=X5=e^Bb.TS5B^8<Q#=N2=^8H97Tg.R]P:(_RA,d^<4VUf[caMUc_\R_)=@>
>c?@T<dG>@.+#+<-:70cC;Jd-A0NQa=3&IaWaR)3+3H<_Wf64FZ<b_U<]<,dE(/(
3f(<_D)?(fQ^BOG9eZ_ILKfA+HL+Qe1N,I.YL_UHVd?C24YAb@STW+&/LV^+-P@E
1(#T=(\@GVGS2W4C=#^,_T55OV3EgDTKCNZT\YJ+c_b.KYWHRSMT[/:_7#&E<,f/
O4F7\aA\aQTX(OFQHTeQF8)&#:)<BA?\^-gIJbaK1d=6-H\JO(P0aReK7aA(H5;>
NAO@W<+4#7+MNQ6SW(DUabg9953c<TbgQWA;<@Y7ZJK?[aH6_5=V#CQINN6bSFQ7
>W_H9Vd/R;JEIRJUBHM/T-Aeg7:aNVLA[RC.gZR==6G>\JM8S51EFW#.4RE/4gaO
<\#<RLEMJ)/1JY7Uc=TCMULLSdP[N;;_4Jd=<&K;^?HQ^[_(X=Yad;1QF5(=]JVO
-La2WM.F?N5L-d]IYdQK2T-A;DNGJ8Q#d#J99VAF&KgW4X&37fBd8,5bS^g?+eI5
),@fa?6P0b^=+40;:&U74g[+6eS::E72EGJ2L3[7EGOMR?LZD);B_5<J&:b-WB63
.(+WSKVWJKcT.HZA^3D#\T,6ED5916?g9>:9,aa6S)d,M>:DVfWA-#]><T<c=Zd;
f61U]:_]cJ=<YVP/M>3EOL:#JT)Vf\Xa6Ma;Gd_>8?,@,G4F>D:DU^:=eRHPb>I&
H^)D6g=<Y/72]W+UMY2FR)XdL,P^\_gLXFU7_Ha9M=K5bW(d2W7DBMAEZXc6]CP0
5=>X6P]@J#/4=LA-fNUQXSP6LB:?UWJ1gME(UP.&>CC<7;5@OS718ZfMBFf[D/52
_1S31-d@Rf)X[FWN>d[C8f+])BD[\\:@Sg(BZ2ZSR@g/BP#P<ba9aV5&-7LKM([E
NY4VD+VVBWdJ;J;IOg7YYLC.4CMafKT3566=X[TM)#5C=N0(cB44DAX<1H,/R9#7
H?@52A#/aT&bG3]6&TF;&b<.dSSc1XZ/BD?9;J+>(#K6b@-:V=&Jf26B1.#CeO5C
>UN:cS_\W@KI]efTA=/<;Q3;JNUe-0e?O6)2PKc-@=YB1cXd#DI.R794OE7Z3I12
G_LL9HQ.7VEFE-JVb&Ec.D>A8E=UHWJRL(K=f78(V8(K-K27B/6FUU2--F9KW(-6
McTLaM7>&eAYJ1^Z[:Y[>_WL/UJ()3P1[[d[N2<[Z-Z)Gf;L1<#CJNF=6E]3Hf<+
[L46U>OMJ4VTAHccDQT;KF\-<BET>UR]-L9/39^&(]ZDDN+=?4RSa?>904LNWWJc
<I=b>2OZ.NfZ=9,ZN.?SGN2gMgg0(g:3>&:P8[I?+3@G<=ZDg<N2<]:OCKQ<2C-?
<2Y=O2BK?6;V-(^_PN](1[?2d<EV88<[gT&ILZ\J8P09Q?MKA4QXfP7TL(0gD._;
;dYG2KSQe)SbA8IgYV3O4JAU(F86KW-7R9e\ZMY6]\AWR&(+e@PYf5,(T\a1M[.<
;4T2]A)eBQZJXf->(+(O,];6b7AbcQ57\cP.aaO;(:T_a\4FSMWF\0AKf7dEA6D^
\<AJf?c0LBU/)P&c2>A(ZN9:M.JX-7bABN+WQ.)S7/F>XWH=7#4g;HI3RaU6^#09
J;3IbEc=5RO_10AL-/&G\Y5E\ZT=JdJT\HR),48ge(YZH89/2,(ZO[Z:L,RVTC7?
MPVKG/M<E,VZ7F0C9^69)OX;O>W.]&8/TNND(0&IJ1?:>]X@)b[)C,.dHTKJH_4;
6H/W_,>;/5ENKB2_ED7<I^HZ/.E?Z5OG2?CX09.V<X45UE,:&YO3Se)V#.;?<b2c
LLe_BM?+_F;4??SDSPI\S\(:G345_0;[#C3O)gLf;K?BB\EHHU:E^0X6K)\bB<6_
=+17^fAf#:B]9KW?SB+3SbV@be?JdB&f7g?KM&cN/#1BS]Q[XJFS=RFV0B\afT16
4\UH^c(]1I/[;HTJN4fb-g)(K,c=IHDI84(-OJ5FgD)d<TNRW-LNWB[86+5B2VcR
,bb/26)b6IQ)RL>aP\:BK.)(>+f:?R3f.-aD;O[M)F@W^6/NES#aS7A]>[HG6,&3
[FS(]6A-aC?]+@FC,5e\)K/BEB>83(:4d]03?D4Z:X)^+90SG(Q,P(43/2Lg.>L8
OEb)LFJO5N#[bU^K15aPB7.0L5[]<K#)XV(FNb:O/R;S<a\:Y7(UFS8+f[FUSc8L
_5^O76OA)(OQX501Z6KEP@F[F/5Vd9R@>dFeCE<Dd1B;HR=88/R&NB6H<VU?e-X[
#bNdf:[E3:3,RSV+,#a;b,HRP3,T@K9;-ONU.(9:Ee5OG1Q1JIga\\MC:-<_JbRW
O1[VVT=-fD)6Gg#H21F=Hed@d3JRX^X@WRJ66W<d92;Q3d_B&SO]/&a166GBV&.G
BX[F^C)8Q@M_N>G1M-T]8e@2:B0H:P4+J^28LB2ND+-ZY;10V&-/dD0O#5W??cN[
L:#86+f3dH\F6_DP?4-eWB1;RXcZX.SFZ3U(2,7=.H[P,O.?EL3L,SS<HDQVaKN3
<7(GfL/;&D+P90IJ)?S]GRe8/.d2Nf;=:)W)9WO9XR)PCHbTAe3Ma\(-;f8g-eMa
5@=WKVBOGH38N0E\GOM=bM&Kf=Nf7?)Z80/eN4)C2XF^)B8dg]]a#4=\G#C\+ZP,
.NX>_G5BY-\>SeYPM6EF:)M+e1S-IPFL_,;3UFWe,.<I^6Pd/5[[NQ:/ffC,>_ca
g-6I;gU.g.XI9K)Y(b@[U&V9cG81H3?LE^Xb&/,O?C=X>VAReX0/^I3[X3[KJ9:f
dWf&598G#=9g^\b-7UVT2&)4[g,;D^V,(gY,)0<&<YEg?QaUg&1,;B=dE;LO&1[^
,0:DacE(:ZIRC:SE29RGYJQ_YBNXU5X>I&LCL83TKaYac-WSeed-7\]aLd@L(U9Z
^-WR5M?C&\A9<4K<)E,HJbAb?5+Zd:dFWH\2eYQ/;<^V8KL;UJY)@CS-3fPXf_;^
A-B0;O#U[VR4&>g)LD^e2JLY0&YC+IW[-]W:U\T@=#CK1L,,<:3=7#[aZ.4-)-OT
\@8-5NKV=[fM^,A>gfB^3Z8f&\A76E9KE^J6CWc\Dc#6(d,N9R#3d@D8#H1W\QQM
[X5N&<QSF<UOb+BW1TGSQQPF3AMW7CZUX5+[gQb_c\4K^(F^=7NY=WNf0Sc+FcH:
5b/eOIHBMYEdW0@L/ZZ]IH8KYgFY1L,^KH<&EY\[Y;&DaPTL8AMV^ETQ4f6ED;Gc
8P+:eAC?&R@BJab/P&FXc^SPaV&]MedKWe++ZY)e@>f&DD+XB(W&g<3=Nc=QGT>F
.,[#dUE]C55/D+[IFYS[bO>+-:SQ\NX@>]dEVb[3OT[IDdYAXN+PcFa#X>I)c\C@
9DV_^gHP9gT(@1ga#N&D.TK=W3.5E4&(?338Z\I?K]W9+3Q]LVN=U^.JYTQK]X(-
91?NC^B4aKEZ-R#0M\Q>&8)(=:@^E(-86&OgZ?,>5NAOPP#D:;:?KPVac,_1&E32
\Md+(g2Mfb6If@Wg<=e8V7&T_C7aaF9./^,Ld>3Q=8Bc0>5D):)9V,MY\83O^daA
)3:EC,@5@=Y9H3V0SW<D?@LJXbDg&C:\CIb2IPJ)4,JeG7)WIR\+5J8:@F#N9\,\
A2aZV:aH,G:STEGPg5UD9<=0B1^:[HLS4R)PdY=@g#Jc?I<(X^c.a.[6aDD(;KG^
deF/BLgX#2d&b@e,AZ0^72&?^<:RQ4)5L-AI\\M>.^9cJO8C=gS2.T_^;b;_M_Ze
8If8&)a^TIGIU(;=E[-W&]E,SAe.RD#b#O3:,M9Bf[>#Dc&J):8gUR:1Z@G>A9(#
/g1?B.BP0T]8DPI00+g>IfSSJKQ<QDEP-]MPA2LEW:dBR2JU,QJT]YDGZC\BKd#d
PW?D#e3;:9_Z12#UbH)];#JB6L::9(G)CcU95g5g4+:TIK[VW4E##B=[.>Q65-<P
1#?,Z2A^cgBb=X<F7:Y1Fc0\VWP(EH<N-6<B(,C8aQVN@S2e\C6&FG?&Y_8P-<-=
c?4?UYbW5e5_+E_\Db?bbA34)CLG7YW[H?-HY=QOX&gN70V-dH9PSP2WcO_VQ^fJ
bf:44:R?eOPeSBT4S,Vd-KM[+ZKg[F:<7;O,IP^Cf)#d[0Z]cPeeR(f/]Z5NB[a\
LE#MVEaWdTZP#.0OM#-I<SO,PK1d4;(^[4OW,c-F_)VaG83Xc[34(<QR_JK?eWB/
-_#1^b+5a).=D0Y@KMTA3/W.AQ7&>9]2;e#D2\KAKDa5gdH26IG:JIAP36dbfN2C
;+9Kd]4J?b/?;_Y8e^e3Rd&51EMZ6DgXK/Y>cfGYeNg)3ETN+Q+>H_4>?MH,\]FM
,cc^9XX(c3]OJ&].)+AV@8LB43dfM?J^eb@Tbd^]#]OPZJg3?K,/HTLD8>N9QB06
N^Bf#+=6R+S;CW-3&2Af:W[8O7RdX[#a<G#Cd<X,Z=.1=-[9RaBK0C_ADg+#b<+Q
6GHAa0.1d6K]Eg7aMVe2.6S^_4:JRO6\3ZGBZe2];7-^b=:DIE,URG#cFgM0Rg1U
L9HC4EFd,faT5^AUEObdS^#GZCf?UN;NR<.9=5L<-<S=,\5)SG<e6Y4_\U2H7HcT
Z<Q,G:a^BLPaENRHT9W>dN34d55O\:VNU9E54W8=<L(8W4SS^=<)EJYA[6.b#6W/
9<eURNJU:9WW;2H2YY]Z5HL:\SU5?eVVaAM<]8AMAY@_:+/fIT_U>gH7-4^::/E#
9Q_[b;4J2EHNG_,X4(_HK-.KIE@8NM7/HdPH2D,\<1Tb4ST#0fN3\]0[H6Q/>C>.
4O9:Pb1d]3S0GM@&#e@[V1IdeKb7F/\RCPgT>_NM-PJ1>L><5T.F4??^ZY;-)WUY
LR1KJ\8b..AfN6Y[.aN7Q([\SV#@YA[Y@3E[?LH102I]2TV^^MDG2L501[bcA_\1
U:1V(#/(7[^5S5K;E<].a,Jb#WPLQ.+6@119=g/YD/NMCUE5be@18Nf_&Xa/Y:1U
d6_]B&<FNW79)f^CeRN6?JGP7XVQRZHV3=^M&D[XB,T9a-9fD)/2M[&B/^JAXV>T
(_DAb<<?GV/Ye))Nd(I3a6C?_aG;&_:U?05;H3D+#RXW>]@aBUc@EW2EbcVN+6\]
W8<_Rd\)QU\.),4(A5<fO4e4J>98<XHJf9//VU+:2/XF0[/7FL[Gd?N4R7aYGW6[
2(E\WG>[_-ZXKH0Ta(SY17_+#W5c3bXOJa/-;+aE9ZE:2?faPHa775IK5TBXH@LG
<AWd7fXWF>&P5)/51g3^#X7955Id>gOf-6Be=J;\9]DWBeeX(/B83FS>AfW3QC7&
Ug,M&AK[cbe1ObE1N(fUSER#X2IAIE0RV859QY(@VAcT]E2A_#YcRF=J01FdbL^;
3@0Z;6d>O--T3FV4@?B_67A.(6(+3,R>NNdeg4BE(A3fc14R(b1KV4(222DW5@+]
MG;9ee@e1SF?,cC&6ZU+P[T]R(Q^47Ld-:E=adY9ZQ9SU?VA6Z#f7(\d=\&OF,FT
9?>[)<7g&=T1cPQN8V((@;c04UP_M.M;856bII480GV+M#<::^f+3Hea::E)21-N
2PR9a&DdM:Y7YG^.QbaYOEg?F)1eg9@LW2eQ0<XRf>2ZdJ<347&Da/dLcQ)Y_HM/
CFES9\F<a@?BcMF?@5E;95\>A_Qc&9)<3g:LUe6H#PN5FT^A3M4\DYT8KL4c3XWF
5)<eK=e28)H=FJV@]?URXWa19Z@dG&WY]?KOgegI/O96/)C.G_&RHQ;W#4gR(-Wf
.7Q6QMO\34?#?S>O3=FE>:L[M8[2_M0(14GfMG:Z<1<-JHS[W91,)Vc\;efgR;Gd
R<&T\_-5a3_UN,SP@1NH683/3aLc#J7c<@SfPHN0cQI2<IZ+J_(=.gH7FQ@S8I6F
Z_K&1^RKaNR-0#(]]SKV^?\0Z0Q#>.g6W4NJA92a,Kg^;XN/aB+#eUP<D:<YZ\.S
=5,O@\ZTX@JM;3T45=^]TKYBa)([EBPgI4W)K@f]e@2]HQ33</#NJc=-LZ,LFfJe
Od0TbAL0TCQ@7+]1Z02/JaKE2_S>&Q_IfYBf?-bG8CL??;:PYQQ0JJJPg0)ODU^P
CVd,[NW-M#3SG#[QPPc2/d<9Gge9RJaEH5&eW:.#]g?&03)6IfP1RK4gZ<Z;>->_
HLF@RQ@EDX_,9;>c4KKWZX19>(<7IXdae,dN(&,aTe#SVZ;a+VWffR1aKI4^H<dY
+5:e339<6I=cY[#/MG:#[6TH-H?#=356W,6GQU7/QeA<=fGIJ/(?O&/I3?0gW[Ke
696&_\UO=UILX=?0b^Y<4)aY:+\BdA1>);cg#Pf^e)0Rg@R(EP^2Z^g8+UDR2K;Q
N\\Y.YH?<gT^(YJTegS(5S/#UYL;b.];RLW))X=a]c+VQ</NL]_^R)S\B)HW.Q1?
/[&;-Ga0e^U[1/eC/9V_U7#ReH\)TcP/P?&1RJ+AK&C0A@T+P:>H2O0AB/fUMU]?
Hbe0_./geK/YUeR7EX_0b>O;=^43GMWIc5V;9;>5-a\7R[9IW+2KP=M-]/]?]1-0
N3-VY&_K=[/7&B3O]d17N)X,dMR&(A\]:,O)-9E5-cX_O^BDM#[/<4WY7X^:M6fe
-2aGQOUK+3fZ1YN:1=6adS)\I.,&74DONBUa)H#)._d@2IEU]RNg2PKD9T1CH.2L
cD\#^4A4Z9B0_ECP9Ha?XH4KG_SdVeg\7P1:b/0[\S[RW//YHN1,LU>M(ND6eKYR
).44Z89V\38J-&O1M45X^3<B4T)@Hf_9&ZB&>;d#RJfNF5/F:-G0>F:Q#BX?PV7P
,L;)YKT]bE[JPNF5G&\F)0XB&UeIJKS8?QF?SZ(C_T<AIB===\=f7YWF7@:GC0HI
M@ID0dY#OL9?5\_Ha^WQO8Z_7,^YG8_74]1:S@9&40[23D<0VbIDZSbBND;fSG[\
c-DK6>[BLY7R5IIaPQde#FJ#^>Q8If=?fDT?M17^QDC;Y)WTQ5[RSRPX3FLJ;8.O
SR1CU.5gcXcFg<M4^/_]cgaGX>.5W@D<8XEL+cLG1HD])^X@QDNbU5HbfaNA7T0\
ZbF0;32;.F#DIa3g8RD]@T9LW,#0KLcJYZNe9.4P>(a[LPAE.-83V]E3Q3bf?6+P
ZdWgUB>)2&1b]?WW]+F?G[D&e1Z\&RaE<.B2[P3&O=Z.X5S-O3Q?7[??1#-VM=([
LU=R0DaRRY,1g4<FHa,AFFR+YD7;GCU_YH<6I\@(N3[OO:a9bW\,g@TJJedD,QHP
,.LTfMAV;((P1dH6fbcSMXfT6^Q[2_/3_7fDc?5P=_C1GZ_>D1#HAOX:=KI_)E9^
Wc[N5U4efDT[d&^.Ff[X&XX5C_IGadIOQ/9P#X]#^->RN+=(:G]eKQAH24=;-\e2
VF8UMGI4,WHDJ+0.S5#9A0,ePcV9RcXN]08EFDO+6/:<a^FHJ+2;KN6.dYG)8AQf
Sc<<.4Fg-/&YL.I4^BMN_T&c>/5.FaZU_RA_dHNQ235.^b/9L5W7HY:6Yg^8IR>L
77E=6US7X^TEbcHT<19>c<5_O3,&=X_6]7gSb_g]9R1TSCgR]?:3^Y.ETLF)EC2a
3^e6&KULcbXUPEUg#,<7U7.IQI#I&Ze[U5feVCR1DUZ12/<COgC1HgI^OD7gZB6>
(ZASYHTI6M6A#>&F^6FM]0Dd?YVO+B_:E72.C^@E,/=gH[3Q>?-^_E2PO.A@R63M
2<Hf7A8GW=g;3N#ZC.UH9TcZ,1B6OUWSSI8?]Qe9/YdT8;N6/+6U<RJ(aA)]CZZ6
cY6(^<JTcV4N&8f-CU8(RCRV3<1B3JK>O6;?O#WI?V#J>I]HKYI=D]FKeXI)#9?N
6JOK6Y7Y)\8#8<F?VM9P1#N3(U+H?4>JJW<g=5Y(RD19<7eYb7>G]?b-dd^JSEQ^
#1.1(Q11D2Y2GIKP,VM:9TGdH3BXaO[]J2I^=F^+_:38>@E5^0473-ec^Y]=(RX>
@,cXe<Dg)R.KLT;e>9g-L124?,4aMBR-:G=KHBRgDfcL=B;B=R2D,<QSObUG_K9&
(\9RGUU5FdCa0[EOCNE(TCWOPV/=Z#L9HF<^(3f?7(PZ)GV-O;7KOH]8R)R&F6b)
[B_KZf)TH+J5?AB>bZ?C0/WV->I[V5CWH10PM[NeM+@):O?5(&a2&[XO?;R2@<,U
<1&E/J=?I#E-_GdAAR^V/@SRc6f5#7TeWB-^b&XWNc)a@@I>KB(XB+SMRU[0X[?8
UP#WaJTBZWOK)QcAV(La81Kg9WAcCU-Lc:K=0\1>:QIbf\RfVJVK<KJ:@_U98)+U
_BTTN,c(]MSD32VK/(D)&\;8XD<R?R:/NJBO4Og91I;ASM:-.a?NK(aDID;a7a\]
aJSbVM;RW6LKZ_2QcMDed64=Z;E)eUc#LNP<T--PdfX\\YCbcM78eQLUb]<JK8bE
19JZE1H93=.Z?0VgM\:7-W2MRbBd/IJOaM8N-^)df]&BZ1Eg@B]g?b>^T(4CX@fH
=1<SLd<<#48BdY>+2&QPaWK=A8@D.9I4e[BM<D229+eI++>HRAN:H,g\VF?Z#X@H
1-Q@2S7F;9M@-?b>@cK5(?05(57_W:EPAEgI>NE_2M\L^Ja7RY&,-/fR&)>492:3
J?-5W)Y?=g-VA_Q,5\<)_5+2Z74=-KdW&V2BEL#(f0?4b^b8Z60ZFfL]H@&eb,;d
a<4gS^cQ.O8,caU>9&PG,NZee<IVX?NP8&WFfFJNYH7/JRSVKc<W,BZDdT(<Z#YD
SH+6/>Z12STf7a^,1T\)LL)YAAX-GRZ=SY6)b2dJBHc:VUCR>/ZRFS1e9;?\(K+;
@Y8a5>7,.N\b2.MY#)7d+^1H1QZXQSRMYK<UQ64)1JbC2Ha3P3=99NU)dH]+]E]J
Mbc\45V2FP4Ab3/GA5K7LBYJQb&LA9WS-KLY(2:7](NPO;80fHOH/.#8L7E36S&b
HK-Pe2SSa_,))FX,R>bSQdFY3VLX_C#:=#f,[&J8@7QP=A7N?012TZ\Y&]:-AVEG
8R#FcM4FeaC2U1BR-S[@)3O,<[R/ReDE#f7JQ.>TXD;cZGNIB\(L?0>Y>P,6b)K7
cbaE/dW=&b78Q\ELab&(KCVA5W]\8gQ4X8UD-8:[KDBXZAAg@5,_OL&bSA1Z<+C&
N1TZ4)[bc8NBEg.UKY&5df2L05Yag\QPb3Kd\G(8=4)feSK7M[S?=#,dN2+3/YGL
ZC.H2N47(e5-^X]R@@16-:,Fdg4KQ>;/#@6X[/O(gZQ7]&d.AQbPN:OJKK4P+T)J
5Y3T+WMJ3;K;f?5S(IZ09[\1I).8.O^4GH33KDdE(eEg:=+PIU4T]D5V@GOB53T1
,;7N4[LOf[OG+,bQL^(dL=8>:GO,O>_>B(G1WX5aJ/@TbPT?#TL7=VV,@bbH=RaX
IWVKaEWWOKU^/B&@RK-F&LJ79ZTITCE(N>KD:BXJKC^V(TMR6P&P79&baafP4(ZP
TAY90I)54JbE(Nd6I6N#bA6W]4BSEP-[]RYNCBM#<,09<<gO<QX=M9<VbKcQ)56,
Q,M)I/WfCZTg75K.aLg@8SI^CdSTCB9\Z,9GfOF#2b?&?G_G?G4AWGT[6B?8YM0T
,2V[g(@IC?TaA;+_cER4L#)/OaW8Le7=5SO]JAHd/26PO_DP:A-@X_1+17MZ4FAO
[Ca-&M_QV6XJWe^E>X62T#^8b6bM(7GB2<c).M,ZP&]YC<bcbZTa\IX48&7JaQW^
aUeV[))YcN9^VD&,(d:348gA6-^d8\7E<[&NdG5d,f0>N@0b)6<9^^XI:;23-0.3
I.]ZS7GCS_8UaD1(CY@Z(B_&^SY01a\D1W5ag>f[_RL.cLWSPT6W&-LGOA<J/;@M
(U(=3,8BH-LA3UV\2A4J=4E=&11W)IT-NSAZ<&/=4c6-J9UYU(1-P=P>:74<M,2B
g,/f9<Rf2J+;LYbYdZ8H3Bf-L#1[SZ0LfC-_:/>AV-M,Z3M-SgL2]N(0&9Y_#H,8
d&J\X#DPWPPP;#;(LgO@-WT:=QW@8QAD>@7SFX#BR<RXS.ZU@T6XMBg:)Fc<_M4J
VIF>Yc0cc2QJS\2;&DePePHYLdUB1I/VA\V?>L:UbN2US7F8eb_;W?]2,CZXT/gD
;ET+edC?D8e=D.-VdKY06cbF^TUZB@42^]9VVJBEO:H>K5XK#gVbe=\TJd8CVOb.
N9&QAX-<Hf>?d4)?9&a/5(fP(U^+#8OI#A,\9KGP@8L0c,gJJ5G<eP6?IcKKGV:#
)S@FD[-HKULR[b?2SL>2<WZ\>V0cQ6e]HEI<gZ59XRPQ)NLfBG4Oc]ebZL9c[_#M
_S=+D2]16E#P^.Z>Kae1?A3+/TX\SG/APK]<[P9YV43E&(g;0XeMG71_Nc7S\gQJ
7KbeZXKAH[>cB.G?gVad@aY=T0Xb<_694d;K\1CU8[7;[9-PFG1+\aSU1J&S>)C9
Hg_U7S66)=&<H@+KPa]4I@@&_Yb<@fKYbR9WOD,WR8=P>:(c2d<HF+645-0,gf39
1S>KKd8MLHbL_@S.T>#d._7.7-@0#/2RE(&TUc/O>+J?F8,NPV/,H(_)Y)9E#^Ne
2SLGQ+Qc5;,W]I,0cbd2<_+5067=IO6LP&Z>b?6)I1)3I5TJ?W)Y?XB>ET64.)>Q
K3aHVSEN)#CY)N:JF0[Pd30V(@LA41dAY(OMZb2S&X0Z1NKZ,+A<^U(]e-0Yd>97
W+E77b&bdW\NP9)61bJ@N4IcdQNVPG]bXa><Ze[)WYU<-]SaEaC8Zc?g,EHP=F_S
HCg>I8LP5J9/2S&&^QY0<-C6BP\C0B5-Z]]9C02&XPEJOfL/9L<W4SOd#7#d:g\(
;S-KM-\)DSGe&TN<CSBB);#/>bNNDQ&Z4::V4gMdHA-8=3;b80Bd[.WFGAME&ZX\
[?3LO,Vd(f=O=CWU_4+YCKLPRT04=M\_(1_)M^,O5+U?4Z&?/JR:KBWRb2Q#<EK5
g>AYA20R?4gE;4#FIV&N3?^]#^Uc-5H((_b.]T)Nb+gVM<G_C?g=WW:ZVD2DAG3>
G.C[JW[7bYO(V4E<:gb&^XE/5V7_g>7#OQYNcf4WBU^HJ1(c9,IccGWV)XCZBW>e
1J4Q+0#T^O9f,@g6@,2b-]Te,JU_GIbV6LfY4#NF2PaL4@:;,9e0U(9K0@<6CP2[
#=_&S,NFK]9Oge:C[P3FG4:eaK#HAcCMg[PHg0XJTeZDCg:eP3V1&^3-MfSI\><f
7bY&ScH+(^JP=JUDTCPEIcT;Z4=La-Y+H,XGBKEYQ6G?>8d.AH9EVI2N732e/T5#
GTQ([E@PI.>F0EG6-G)08YXgYXRgSfY\g,Z;^O.d1)F.+Nb+D1ea#))W.,_8@?>a
_\NSIR>gZ?)TMH/d)TPMHOYYKH>CGJfaXS<]gC<#^QSPa\FU7aaV#.:,JCYLAN1@
R#V<.UGI3Ja,fNW&F,U8+\P#TYR_INRAPgUGJ5]H2QD-9RdH[X#;KK6:)0IOD@KI
7Xf1D&+?<1OR;^[1R^S,f>1-?9VJ+B47M.H6MXU\D\.J2gV&;6-F<_G45Ogc;H/M
N:B)S0^)NI+=c&6NFeHAg,1eJIY\ee\Dea6-/Q4LD)2S8B7KW77J:SJe>.Acg8H;
:VF_\bT5McTVQVI1NR2,YI.VF(<\8._1e[1&AaA[AHPD4)HOJFAL]-Zb4#U:;2c:
JMN5=C&:4]M:TSCT,TY+(R@TWZLBOOb]Eb<4,<P&/99B(L4@0a4=YU5e01AK+bf]
LR55/_fO75^)fA41ND4eB>Ob^3=\K=VJ[=Y=B.NKNRGJ.6_&^_TNaaI[QS@M5Xf8
E+76TGCTcK\CBH:D[FNMc<d6.bAQ.,@Cd05BN:F2,L5D.Ye2P2:Y+/:\gG1-Y6eQ
2Nc@WKLU>A&d>OMS#>=YX1g.,0XH,/E/e(X-^;WJF5G+-V]:M15@QcX\-e&&Q1ZE
AbHRQO;#^XU(IOAU>Df@1fgOEQ7_0X-?=dQN9UY/?@_/25f;VQ4]/A<RT3;1/:WO
MW5_?3C,@8_Bb#e2#7)fFEPL-eXcaMOFFGXZIe:.MBGJ3C>PN8&a4N02JLQD+U)[
93+BE(fCf<?\MECg,6<_M3I;W-c[9)(Vf362ZD+9/+W\)\6L0/MCJ(fX3AA>F^:5
feFPN&#[^JF^.[Y+7]d2K,8>@@^XJ&LFEd/F/3[fCA2(HDHUURP,^)dDK+.K1:4A
+Y\_?<G0dc\NYfJ,R2cP_<-bY^dRT5LCY9fP<NSM7;=&EUCCA_837Z,e;C//:J=L
A<3X(C]LOAJJ-bJ]UZJbf#45KX_+H)A1SK6W.\Z80RW-KVg#CfPL6TP?;.2\2\#:
U#^S0KfcYWU6<)W@N7.OA\78e:[48(3\9KX.H02=&H/24K]3>X2/]O9];AT)J&4=
/-c?T\2cZ0\eS/UUFP&2Pc[ES>bgFEGcV<54SX^e9QH:S,[B9)_8+VU_^V\ef,b:
[4Ze\IBWUQL0D+2E,JS&O?g]<O7S=B0E,JMd#UZXLeNAVPHHJL6=c+J@M<BYW>@Y
aM7bZ7QX1]7YD5?]><M.]PI72aKV6^0Z,(Ed[YY2:5M.62L_]0\+DG11XN[\UJB@
ROdKP56>0,<[4a\..Fe?TJ=POJ6HF9KIZ07P3GcOa/N:IWc;.ZWK?<K9KfPVTcWT
Xe6/X&8.5;)HV)c-NV2cURFEL=(O6XCN&;eg;HaM6\f5cbg3=QXeKIdeIA[+2^<N
F_(I\WY.cI3^[TCY-]0.1FR:#_]E(CP=4&5T<_9KE(KK\Ab#IEXM-^=;OC3@Af9G
UXEeM1/PCfb^W[QTJ6:2979YDHTS9Y_#X([/?=+Z,dPbEa=DbE2HbUW,WI?;Q@EE
&f#AS07IV@aHLTD>10.:WXDQ;,]E<8C/c=3cT</:9P49cA5VJ4b0\[T>C61I#N,c
QO-,0a.96I@IZ-(2<+BT)<&AR6a&#1@Q:R-fdJ_\UDDB;IcRUMdWW@3;@EPXRET0
YOU7>=#ZGO^2(+bFO\]dCE@)4gb8:/^VaVIWRJ<G;AW#)MZ(8RK-V,?@dc_Y:XgT
60[5;0B4[7&1UfR]I@bO[IT&=HG7K8O]OJ<c.]5gA,5Y)c=#F0K(_KI0,^Z>QbX(
W&]fR>CHZ^DG7_Xg&CG;2BdLfg==JO[c+DW9>&=WgX,I7O-21YZ:RV)=]2JBLd/)
^_MJ<NOfNX5W2>6U?1b&LTM:-STPF^(=cf?4GMS?]>:O@<-a>-X;[S:OXegWK\RV
&13GHUd;@BU#+fNQZOXSGHFIgfT2Q7(gGZEC\7T88+fX(JY)EZ(9^=QDPf[Z9K<=
8YN\/df_U:c]//LMK5&@=AbNL+M7T691LNC1OIg7PV&J-<0O&9d)c/_ZIe/CL577
>f11gM]g@<b40M^CV>ZU62HY=)YMG,NE-bbNH200C&C^A07\gDW[0eBZ6G7&6150
#+,G2.O4(b4GDd<;9IP<-^V60H+&]fa/3FL-\0)gc@SRO6_6:ES0<P,;=eE,;VTT
)BDC8YXb(QE>B^@\NVO:]Nc/E8,L+a88d_9c7\8?<N6D&b:a/M,Nf[L54c]>WC:\
;^a+6[B?fNdRV@#)Q)[V&Q3Y2K3Gg&KHN@ZTO9SOJY7M^^Q18)QCEZ/=>(<+YC[&
;BG^-<TIc[fL7d\#OJg/+YI[IIWXW.E,2L#A:3RGFDML<:9:#7_)cNOd8;&?FJPB
8eVC)7#T:g/1PWUDXZ[YX2L[V8</A>.P4]^e\8GWTPS&&YG4#>9ZKD&]_[P6OE/1
\/gFeS_V^.H9G4/^)FGO.K<H,g+-#cY.]a77#T21dUaMd[(dR(3<WK@UP4PEV[gf
SKY2_f5&dY8bV9:-@Q8@^SN7/-7(LSKP:]aGTaaB0?eT:[:UW./+FR#N0N+E_M15
S0@:c5^b#Jc/7A:[WVD\/FG-ZXbd4.CAEgeH#.N7=IUZ>_N);)<<;PgSF[_@#Z-B
f^7&U(^)/O7,G&8KB,8J[/B8(<GM1LX8]4+DBH2>De]CK@e\eW-UMS[d@L@Fb6Oa
>5B:;K#^IF[?E4-HSXKUZcZGS?4G^_(AgR5GP/,ZBRAEFVYT?a)U4YEQKg,d;FgA
KH#0E@Bdg<[HRJgZ;gH(><<V@I[)^#VEYU&ZM5K;8fb1c,g[JIEH@E1XF,W=I80=
]=B-R@1TIX.PRBFF?)#:3PDf.e=:DLf-HP(B)e1.GDL0d5P@+=<QBJFV=X@U#:=Q
:)b2C<S:L_A658aZUSeV?)c;+9(e:APPeZ6H/IaHV?@+3JFXEH<4e-<bRg7-\C65
H0^0F9,/LP\f[RM6d<aKfFQCKFfKR1]/X[8P3?c_?_-e@CSAI?a<GQe;bb)C6@Ye
,MgX;aC?g.bb-JK0I@4Wb4TIEOO)<GI>aH:7AO97;^RV+\GeN;M)5eIP@?4O6=NI
6?:L]N#c4Q;6^CLM)[d:^_>A4TX1((CRf;HdKQ+aAgSG;T2@f99H\63<I-,eYS[M
;3W5+K?#R?)KG=R9f_a)]_Ib<0bgFE,aKK2aLZ]K,+=7UT2ZQTf]@JdXJbO,,IW]
(S:C?&?Y.&O2Y5-?3F3,-dY?\-F]]g,<0X@QFY7FbYDdOS>PG,Tb68a>?YXL@:1#
P0^1@D=W5UB[@f+Z)&B5W&[e/]J4)&R2AJ&9IV8P;cFFUJT@JI[75[1aP2QdSU[F
#g58R?fU9H>V1T[SIRV-?@28KQWL:RbU;=V]5:QY;DGTNV9&2^I73b1A:QDV&R?1
[3)-(#QX7O4G@JI+?OOUb./]\BH+a<)]&-5^5\S0e6+5(06SY@2KG[(0&PB.HW\,
9N9KC,/1;&OHS8V^LJ?S6]cYHQ)/M.8YG>;YaXF8@MCf<L6a-NTNfW=D_1Q[S]O5
,?(E)GfSA0,d-B\P[b,G_fe[QSA1><52+CI04PL8N5W&BI7;Q2>#g8#Y<+I^+Dc7
J;.RPc42PWH<KP??2614CS=fG_WQLT(4=7)F44\G0&e=?+\e?(;L\(fAA0&]_^2G
T.W3MN^bIHVX4@6G?F3AKP=56N<IS&,V=TcePd@8;P=:KC.J/83<#?T0UACQ#=TY
V[;12C5=SA+IYOCEAV.()Yae;<C\(/&L<?J.>.?:J/>S&23,HQWWKL[POMEc8+(#
BRb5NW&B6PP,Wd0+5]#=IcH8f2cLeaWc-/Q]:ROGFdgF#\dM&8(9J[KC6771@#F,
,KW[G]3G\N4M,HV6Y/a-)-5YL9^V-L#OXaQb/FTf0/(U5GJa?I+7Tb-^GO8B#[fD
DP2,E/OO;MLW7#1C78MMX?f[ZX?^PceI3&^I4QN9GfaX2Y;_Of4@&A>P+2&9VRL^
Sa]B\_XD:d>g88Y#8XCANG_WR^)@@#f@E&2Fb4D7EF3N=L?^<aQa^DC(^ON[8.[)
GY?H).X<8.6E6Bf;X@JMGf<baAD/2XI>&5,65E^dc96M,EO;LBAG\SfA:T/AT&8\
GOO8D3DZ@_^_b((PQJ(3K(\[7<LQITQ_3BKS4+9=,4Q)Ib@,39:S\\8WJ5.W#b6c
dQC4>;,N8Ob-8W[>C3:XM#8]5Bb#=U_>O@PS\7+33CTM530MFedP5.JHAY]6A;ZK
C6NZ1c=8Q9O9HK#.+G]96bMc<1&G8GT]a>M#MH@(A1S:e0PHHRREZAL^M[V8S>55
e(C_fA,N,92B0A81a7P#]9[Q_HE>V@/)8(aLHW6C\^?f?cGc,gfRM?B0VN#1LgM>
KfX\T\KZ3D6T1T2_@OXd(/K(0?f@b3P1]XED0gM3E^7-SCK&4&c1^0<_R6:<_GbD
-#D/F-H@;+B>J.<#WC#3=AfJ)R__gCe:S(D/S,_^JWZVF6aE1gZZgE[;cfN4A&:e
I]/D&E,6JTI]X(J@>^f.Pd](-)LL5V,5[@>ER[=Zf_fRL-?1/Db0I5H1M#)WUaa/
Cd@UU\>Y_gG?gKY-E3E:RdV/=+9A=LdXf1,9F):-/f(RWg5RCXD:C/12Y0<8X+A6
0MeT14H_[U6IFfK+O4PfMC)WVW7BS;@dd#5eW7S<NA1QV[&+^A4Z4B0-\3Z,HO3)
d=bV]HE&b542VU2UeYCa9)&+EH8_ZM>TH-ZY&D4[W2>O2O>1JT/ELUED6f)W@W:]
\0Y3Q/11Z(\^\&7<4K?52OKfCI1)4c5G/8PVG@@/5/5HZ-W<UT9N?5PJWgE&O;V>
:H@&dfH#@NI@0?C@89)WX2_@Q/\):11aIbHTc6RS#bNcSL;6g(N=59<]D=JD^C+P
X@ZHfE&d?PSMIJJ&0JH8&;>1H&\9KT:<MBVNe3D&Cc4e7aN5,/&U;A)WV.#YPQ1>
g0gWTI:Ae@F/FU(FX.e7P>(C7AaK\G:PIJEd(A+\B<Yg--@Y^7GbZ]a/O3E\>7I)
/T,S,2JXKP33X6[b-EB)eTK#R&Q5\9R^[#-d]T#>a>B9;(2BG,:VF(LJIS94)5+?
W@_d?(5Y7.+YKQ8&9-(Q):->Y&^P^ZJ1F(A;V4K-1##H>CX<4Fd)OaD:<PgIJ(P_
?+],7Hc\A@+.Z/-UZ#)7GBLE1QZHbc/^O1CXPEOC)FA_F\a=FN&Eg^/^W6f(.)[G
1^&K.C8.0K5Uf21FW+HE[_b]WH&,#DFL<V[=WSgRV)(>W=/\J.++_3e^6QO-O\^2
36)-(M^aYf=d]X[2NcDEOO=L>5DX8+-;,1T1>Z+Z]LRVe>K_.DS_]Hg+MT>/gS/+
BS=#P3MaTB+9d33H2Z6JYY/^g.5K_AJOEC8P=E.dLef/M70:A4[b;N[^Fd-]U.#Y
=WY+9)Q5^ULT\LU5C@LcW\_9[X?\H\R[Q]9IJcRF?GW?aeBGGET]b=\McT#P]#b#
5X0^]R_AA.^=RJ#T947SKRQ5:8b[LU8+U]=WR_>Ma7SC2SVd<GD?TRYVA-Y_g:cW
VU.7NG9KPLb6Ye=7T;:\XKaZ;T@]G4496MGbdW?.>+.)0_UXO659.ZKbf>K5,UO2
QE9:9D;(\].C(FNJM+g^[gf^=#^JC?598SK[eDb(c8P)85\b(Z__^ZEe-;CX#b-0
H9ZeNcG7Q.G.:Rg.U#3UKW/.[Y.>0)#<bLZ4?2K(#,9@e/:>GH:\W.BEG^B:A.+B
:?P_d063Z[JY1Y[e,^W2@0PdR]5E=T,5W&B&\<]<I>fHJ&:>_+D5+5?N_AA#Rf&Z
FLbNTRdW2UYD(bT]5RGcK<AMbdM@>ISQAR?5A#=8&BV(-\6NO.DMN>XQL&A^<ZYA
0Q]U-X=B_6fg#.VF1T&.a(9<))Ea;@GNG?37_A]1#HH@]]0R:2H(a[Z,APE<@0L-
O1#A\bL0F,Pfc[<Z/KF[+#3P12(VHWd/cKS=/)K[672LBd@K9)+YW\=VE:)6+(Q^
FK6K<=\8aY70VE-J^Z3^8TfdK1HII:HE;\Za4A6<K(Jg^SG\FL^c(X5dD@N71<b3
J:3WSQM.GM]8/&.40K3ZT<ZDBLX5S2_eKYdY[&Kb94L>@5(+OF/5GYU:OP&ROH4C
Oe54X-F.YN[c71(<)b#]Z.+W4-089::G/4H/\1+4fC#.dfd6:S6:=DW:Ue\cI(fY
\<F-=X#)=DfA9gbGU4,YC=?PE:O+;YYeD)]_OL+MK9OE5TZ@e1S#2,Q1g6KTVHE:
+7+)]Ia&-FY:WNI,8O3H\d(Mc@H<ELEDJR0Nd;4IQPZ1?GE37eKH(42L>OgLF<OL
e[d0d@72:0#MS84+QN9IaV:FW-A+?VA,a<+>g0?#@a3NKe1B6>B^T)b5V-9?^->D
UObd>_=B5]a[0\5,K\[7TfVJ8Y:>T2KXR:gc:+X=eV&NL4^<[-9XRWTKAC+c+7Rb
c&W,HZ&4)bEgOEX(XLX>SV2-@PN4U[U]<Ie^Ad@@L\V@UZO^F^<dBD^?W-TcC]F?
4S4aB:GXSNV.[)R(?F]H.A.]UXEUaF;6QbOJJYN6CPA@ZcTQC,1F::ZQ]J>#+dJa
6fH\8ceDEIb^T549#E-g17KET3Fc(3gV4b#O^BUe/(BI0O;bDLX/CIEfY,cUfP04
)PM,^BX07R<.GN];OB)E_+8SC)e46B]XK=)dQ,VRfXU7DFNETV0-9^#a76P7&2\+
+?PG(Y3QfX,](Q5/]FUca-KE6>&0cb)VR64;H\H<d<B-DF18XcT][V?_NZ338MN2
&OX2ZSMDZ7+Rg\DQQ^b#^YXUBUXa]7W.0[S.c3fW\_SN<>SeBeO>PNYbB^5YVTdN
J(<EFT0F1[93ME0>TW#e1\97R[dM[.97H2V8&\F8DbG6\FW<_fFgYY475K4;8a;L
YH;[f;7W:6DVV94f.&6:2O\(?SO)/#XUS]25/Kf(Za>R7f0-5E4H5KY(YU/-aVPA
2+S2^Q6Ga?bG,#NW&<[;9Q<[W=ME;34_2[54d=[YIEP[b,3B^0>FG<8<bgS;;&=d
+8QO2c3R8RHc6Ub3-cNY=..Yf8XZ))M.?aY5X^J.NASB,9:/QO),,@3J/gI\JY(Q
6]EA,,#eK@?KZREccb@3@CR@(N[IE&]8NbNBgcNXW4a_&)\ea3Z:eW#-R\D=?ORY
Gg@36gLgES[^?d@Q/JJ7AOb0H:@7R0O^_Lb(9T[FP(EO53YCeAE_[UG@,TU?f]BX
(G&0+AJIL<4-_YSG\d5P,30a,Y=Y]1L7>C-NBfNXO(VS)^8W8HCG>e1&N[e9]A9D
5V(OA_#Q0=&DB#I08gDg(&W7P@Q+L8Fe3g:b@\aX33_T9[OVYA((+fO,=HXWb9/V
Jf4FO<AG_T6R..L[Ga/5O0+;?5cdG=@HL82Pd1#KPYH.9]P1WXW8X^Sa/./?WTgG
.c&;(#JH&Bg;b&5]KMeAS&J7CT-T&F8?);UE6CbSE&C8O?,a6ORO&V_TWX+Q@BaM
bN)+BY(?6ZC#LE;H5aEOH&c9SCT_;T9MX..92fX/&T21@@g;K_V_0Oge8;T18=[\
>_?FC.9KNX(.[^_A+&a^COJL63=c].L?/ca1EVJ<4D3>AC2a&6_6^LL4\.NIWMEX
NaSA5=C&]X9D+)>/aR@DSJ=&JKed7O3bb^eVOb8K4e];)O>R1fQJNP_Y&f8?eCZ1
?#/Oae9f9Y#MU/7/PM&:9-Q=9^gZNQHMN[#M-78(>95a>D?-2(cAM7G4e-g-CSNV
H79\SNcQM1HAWDQ8\B_e&XVaJ\1F71\1SQA=aQG@1:SOZ.NgTPJ+A&PQ_gG9H1WQ
8CH,bQNDa0GfS5(]8W=PP#]F@/RBPTeA\R&<]bX+4dKUP[O634Ae^.L#?LJ86;W<
8K/BOD[NaC^a&&/:b#\TW.BYRM.Ma2KM>1g.=/NPC=R>U,QGeeB#7W&6@Xd^]6YS
[I^#[Q/6aT5DM?OQOBCK?[CFEf+NK<X;T>AEK_1eb^e+7K8?[RZWZ=Y)/bX5Y22L
.S6W1TB67c3_2RM0LL&IUN31G.,(\M0F+fS]Q0C?1eaP\0\B556E;JG3MC&<&Y_<
XHfJd)M<Z7YI&B[aJ_XN]_<IS6B5c8L8C@QU4QR)K&>8GG?cS[,JA]a3\74dHJed
9YV<]5HGA);?IE+?FW.c\AMY?M7?Q.GE743@+W]A)?@#G]PH(O;PP#VO)8&:6LbI
7OMd^fM0M??YH3TCX_([YZ<7:E@@T[AG)OUK_(SZ9GG<8Z2g_8Sb_HL&:\@D_DO=
LZ2/T@6=FS\<cdM=23E<#7cWA#:+>cR>VN/T^9g.)Z#<0\&a:YV^KK:^#:Z/;KEV
71/IMae-M+V-\Jd1P/b^.FOZc1cc=-?Z=RH\R^IUDSRbfDH>7MR:.\+Kf_b<e4\\
;@K]0O=g;;)-FV_\4LA=T;ZPd-M^L@@8TbFOEd,SaC^U1<OQE>VKCBLa186M<#@Z
GY,>867J:3&+Je:AWGX]d^HX+1+gdLX.O12<.2c1E=]0)Za7^7/^-5KXYa:CdZ3\
4>_UPa0C/J/9cQEVCU5URE@];G>1bH3_UbA0UT\7I/[eK-G3eVJ06\>DKL/);C^_
#>>R&QX?7H-FcVfU:02WC<N3aHTPY>-2->M6^aNGJ8Z,a++VeT[-G54(7,Q2;#]5
N:=<CBG1G>>\O4]VMKbJ,>6@C;a(8]5E1eQETU6aaKT#N[:,KV0E-9<NdO:4Q--C
CHMcS?Y]e<F46A3/Y:;YXUFg(T5:cRAJTIY+c(.L0SWb=d76+FQ>1TKRNg28_,IN
QYB51c1R7SdU-XE3((8:?@1>GOOCG@A,YNF2UU5-D63>A6EI[_^Z#2=94V(MEd@F
F4S3_WPX_1<PH(VaEB(R(B;HO+U_U@IJ.aV;Q+<>=6gbO:B1CH-3/bW?dS(Z,]P8
UM8=_SeF).BXc:dO[f,JGNQXY0[7^=bTb9C:gc(JM]5g]3,f1f7U_>RR9T[EA_J-
fNF((B+KWKQeAaA:6,D1Jc-F7DET647J?:+2ZWOTO.c[7UOf80/P?KWG\e1GgL4M
ebFc\54V:+bT5I\TJ5Z_/gL)KfJQfg)RcZY1+e>I,K(6YQH3-K.LK[LP+F_>&A/>
F-F3[6aP&)EV5g:JU?0L3=/,62Eg2aB>e>^S&5_e<QPR@]e3?ZO0NKdC:9ZR#@NM
a.;66+U0/@XZUfBQ_>_0b>6+H>DN0++D7L94IbFLB&K>L,DB2)&YGL2E+FJNc(@3
8A2LQ^/.f@ZKCMd8TMg+IcA;^>7<W@CMNU;W_FCGD3ccA&FEZNUDHOfPI:0KHacF
]H@]43KCHA?FU01?0.P63;&<9bM#_9+_H69bfLg[g@BTb#e#36PV==A2E5eCT0;-
Y0FO;\<ZIN>Z)RV]FIC:U;P4a13aK9aIY0fJ(Qb8:HeFCH5W?.e\N0_WQKO@JcaA
I8DIVUEG.7BHEdeNDLBL[:H16<)FaL5d(M_76,[B^@]0#2F^ad;)RC>_S0&7U@5K
DXbIgd\0SD3.ZT/T/2c9X,fGYDZ;M(Q7?GB8Q1#E:Y?c>GdR8-I<TD6_5Nd1,<LC
NEQ(.;/NM53+#/QRG>)cLEQ=?(UW=U4=f]S+?W4AdE#cWREYR:FX<L7W_[:E::fV
TCBOTD69:_Lce-6/=;7IRN&ZB>I;0<1C?8=>97+g=I<3E4gH.G4+E]/@GH[,J6Y#
W6H.)>W:XY7@(@/YV^4#\;gAD(;<OY=>a_F/5[g7I1H2JZ^fLEZME-LD:1V2]0K2
KJ2:_);Yd)=.-STJV[P#4dS=9;F;?HVO:BW<MN?;bZ4?-YWTV11ZMGQ?R1V;IRT\
OHW=NYC31LO7^6cEFW^#\M:Od]Z67P-NVO/QF0EP<aY(5O(1XSX-.IKZ&Fg7J\aO
L_L;=KV1g<gB::JU?aWXV]A:,d/0d>Z>L>3bH_MaeA1=S9a4+&8QPC_CW:)#b#cf
KX3&CXWHL@O^RA^[ceB9X^F4/XY@\NTS3NQ:]3>A_0bJ:d2D0J<(<TdbOY=U\EO[
&T]O>+13b^NaIFb?#MD.gP+0L_a3]0TP1R[b(I=/g=:4g6WWN839Y/c:RNMMU5WT
<6<EB0Ag00=0NC@.E64#SX8KAV,a,OA@AX<M2)2bgQO4X7PL(SNK3D+<-Acb)fQ^
BDEEe\2A\34Q-QXS4AJ-Fg]:PK#]ZIbLc@\-1VZ=9,E]87EMHH:[Y5,(^C])9XaQ
Q=gFALH12c#FC]@b,G:;:[2SW#N??9,=R,V7/R6>T(P,SNgNg;P-Fe(1f_BM8gA:
N5GIO/BeM9I++b=8FD-;gB1C+5]IOFI=/Mf_-N_31IUPTJ2RK]U^\+eYH1\Q5aV&
De-R4-CT..E.H?JXR&\>Sf[P3=Af+\.J,?JQV?O-<9U=-cU-Q29R910F5<5^Yd)2
=ET\K0H\KYX6cR_S;eQ6V._;Jc;GYV11Q/29T9<+O]/^N0a2gg&\e,=/C[+R?/I>
]ge_:AP#=S_VNK,6=P6-\MBgaDMSQK2@(^<-S(H0]e_C87B>f]@KVYAZ4QE-FBWd
S7/3-=?NN)ERRTSe+]+RB9)6b;XLWH\UaH\\B5]S9Z3S^G?Q+B7E^D_&<2]PY.Eg
UC3J0(E@@8d3e69_0PT)-L8Z<SXE[aAeEMeQ3\,;H7POX6>;+C74>](.67/&5YF:
^a3B])\XL5?LC2Qc(#6-CD()&_QOa/.RJ[DO(EAfWJV+f>-F+-_KS7U6^L.<Nb_Q
S#2J5--dbX=,(>@[K-08>b8+]dJc6_CbXIKJ7FK;6Q,dR<SYIKcd2K7]CeS,Z<VM
N2F+5H=cG5.)e.5HDZ<3(IULL,E9)TB#L]H&0c#;Ig#171e/Za/^7^EQ<4@FT.3)
SJa)#D>-Pb+.HTF+SBG@DJe;7ccP/?VUHHd+3]TS<Sa<NE(6N)PEB:9TOO6/?Z=8
J<_U[WE>b+#+X3J-V/I@MKBKG=6A;P]<Y]fGX@aPZ1MZARHTS0P_bUHOB>:7.2_[
][#.2/7(g94=<N4,Kb./3D[fe83WWN<M=;B,;,dX:^PUb\^U3].\Ce=#HXTbSO^K
JY=\[0KEZNacO+SX7\)Zc(:5PBK4<JL:VS,W^2#3eQ0FDIE<Q9?Xg.#BUOdFcI[=
;,E^Gd[R(dHdWZNW;?2H_=(NTfWW&T>?Z7+(RTgN8F^bWA=50D@cSXS&UfU6@PK0
LQ;+Xe3=aEYZX2_=;PHM]7ZHZ,]]NJBdHL\[8KKbCa5MHc6E@_2/AD?be[,gfcUX
GRe@@QJYNU(P3d4V:KW+,aHDHX/S;843)/bL25VgDbB)1\gDC#+f634.U17a^9E)
HIQ1d7D@J)4EX4(AS:(6@WUEW,RP8HRdLL<cGSD\74cX)M.FN9]O9P)#<\LM5,6X
364UEW5&G5:RfM13aQQ,==O-V4#K0WAbOL62&\?4@d25Yca2aY/<Ucf&D@)YIL5C
[>Wd#Q<IC5QV/K44(Rf6]>^8M)<M3QO94_2-LI-D;I6;GR,J[a<064KP61HWZBP8
>M&S-)&--I5YCUT8,WE7JHKUEKKb]efI_=MS.]&9YE+2d2[/AVM&46@A,<.;S)?_
/7R/\19R8OBCcJ1:+b^2-QNA\Q.<3S>3B#,.I[&\CZIJT=3aSf(\1QI5OS<gd:>F
<CJ,WeGZe2AcTLAcK+PQ;(4]K_MQ]&-I^<X9d]6I_>&,J.K)#-\^V9AbLX[aD6EU
A7d=N>;YUP_^5Oa\7.PZ<6\FUKZN&5Wad/);INMJPd(YU63)UC(Q9fbT3WYL)3^6
:+^V,0:(HE.@QR_4)93babe4<?\(&X:+8bM]I#Ub5HH5eQ?Wd=2GdA3C;_-29-gV
-<9:>#TDJI+K8gJ.X;69.3C>LGI+BM.bG]DgcfB<;Fbe>LWBW9]TgYMeZTE0?3gT
&=Q+2JY_^9OE;e&1ObRf+XLJ-gFf9EZ4^dF5[(D^B;_X45J-07_AY,J?))c?BG:6
8,9MG@^Q;:&#9<PIT;KUD<<TTBM1<AI7gONfS[dKHVbX@0C@WPL9B5f2A9FZEg/C
WMLA-6Q;e>TN::4CI@We[1GA?MGaKZB#\5gD,97c#=]UC_E+_<:HOQ/@-Geg3+_g
SQ@;;3O3J:NS>5?XU2A4\[8X>I_57g2fF+Ac7@\^M?]Y0Xf05C#^.(.(WGL1HM0_
<a[X4S/>bX^VPZET<bYT4FE8VG?V^aQ2#Q7CAE6YS:F-NEM(CR-8PBJ#HQbU]=KY
-,<2Y=]e-&K2Q)bg_?-5ZdCY2+9[Z,?/Ia,QMRK([&LE6CP.MTK@3O]C132P:3NK
_DO:d-8K8GS<A]QUF1)<\0E\f1H\g@\cT\&VL9bBY@:Yg][=OdC&CfU(FKF8QQ)e
>ac8c73&LE&M3Wb.-219/]ObRd9-/K+L?^/6L1?[P\7/L_;UI7VD0I>G2^=ffSSM
5(ROW>^P:^K9H.58N3^W+WEcfTU&c5<8,53H)+OOP]a#IJdZ=CX(.<(a:H&T\&06
EL<#4NCXO/M:;?<^9a>UD\ge#3X9Xfb89O@K_+@_<(DCLL^JRVAf7Fe#0DU1O(C2
/2>O8:,0/e6Q261)KgMfOS>X/08?9SGU-fTa@4V3]S:JcUF3P7;e1I&([PI5(.8+
YG@2Zafa3f^)VI&^F[SR.A-)2WV\X_4T_6KY#P77A#R3C1>)@ZC82(?^N^P-YcKS
6d&VaS]gfNg_5#_;7ERXabU&[e(9?C),N#HI3(NUA,bLS4F&(/aY-MN/>PcT8O#3
.5)E]:<O(\3HH3(B8)3TFZd)6@@DS(cD=gSYJM3P[?a3.Vb^4>J,Y4V/_Vc\a=M<
d-\EO>8e9cbH:N6a6aC]W7IMOHbgG4@4\/5P/D<[<=.OF\b5DX6/=_c2:Y1:^9F:
W^B-[7LX)Y?)Y?K@NeAZfC?[,VY^#Z>.KUIT(^OGe(Je0^?SG@e.S7a2VR>)YS]>
XJ?BVL]P)@L25?X\1?34<Q?Eg90&_6^?aVT@TYJJLP\XER)LB82#+ZJEV.I]Z_MQ
2CLL\?03JbWR+I#F8E,7A8EEH,EaTXL;TFdVP:#c,C[?-KH7YGdM6B[:Z).49(EK
.D6MdW1^^H5R,$
`endprotected


`endif //GUARD_SVT_AHB_SYSTEM_CONFIGURATION_SV
