// =============================================================================
/**
 * Class containing the events for scenario observed in svt_chi_transactions.
 */
`ifndef GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
`define GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV

class svt_chi_scenario_coverage_database;

  /** CHI Node Configuration object */
  svt_chi_node_configuration  cfg;

  /** Array of pattern sequences that we wish to match against covered transactions*/
  svt_pattern_sequence  cov_scenario_seq[int];

  /** CHI transaction scenario coverage */
  svt_chi_transaction  xact = null;

  /**
   * When a cov_seq_match is triggered as part of a match, this variable contains
   * a list of the objects (i.e., strongly typed) matching the
   * pattern sequence.
   */
`ifdef SVT_VMM_TECHNOLOGY
  svt_data_queue_iter  cov_seq_iter[int];
`else
  svt_sequence_item_base_queue_iter  cov_seq_iter[int];
`endif

`protected
V#=@BfKWJcg+H&S35I1PVOK.J,4VIC?g1R3+D>RH67@d\Q/._]Qa6)]dJK>.K2eP
A<3C+<V7^O2,ZGIPgA2]V=K.2$
`endprotected
  

  /**
   * Table 2-9:: Order between Transactions
   * Applicable for only CHI Issue B Specificaiton
   */
  int  order_between_transaction_sequence = -1;

  /**
   * 4.2.3 Write transactions:: CopyBack Transactions
   */
  int  copyback_transaction_sequence = -1;

  /**
   * Retry/Cancel Transaction Sequence
   */
  int  retry_or_cancel_transaction_sequence = -1;

  /**
   * DVM Operation Transaction Sequence
   */
  int  dvm_operation_transaction_sequence = -1;

  /**
   * Exclusive Accesses Transaction Sequence
   */
  int  exclusive_accesses_pair_transaction_sequence = -1;


  // ****************************************************************************
  // Sampling Events
  // ****************************************************************************
  event  order_between_transaction_event;
  event  copyback_transaction_event;
  event  retry_or_cancel_transaction_event;
  event  dvm_operation_transaction_event;
  event  exclusive_accesses_transaction_event;

  `ifdef SVT_CHI_ISSUE_E_ENABLE
    event  memory_tagging_transaction_event;
  `endif


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new svt_chi_scenario_coverage_database instance.
   * @param cfg CHI Node Configuration handle.
  */
  extern function new(svt_chi_node_configuration cfg);

  //----------------------------------------------------------------------------
  /**
   * Method to kick off the dynamic pattern match processes. This forks off one
   * process for each pattern sequence in cov_scenario_seq. This function forks off processes
   * which will stay alive until halted by a the component which initiated the call to
   * this method.
   *
   */
  extern virtual function void activate_dynamic_pattern_match();

  extern virtual function void cover_xact(svt_chi_transaction xact);



endclass

// =============================================================================

`protected
XJ:IL82H047>efAg,FPdeM7WO4LJ7Gc?aCGUXIQQe1?&F^ZZWT]P&)ZH\C801@\>
1\(5J3M)P0F/R<@+Y9U.T3N&HF6H@XV3SM#42EG_>(G\-AO=]IU9U-D80&OZKIJ#
)=5-9e(Z7OB=OM;P&e:^3ZUD>LM^E0Z7I.4]<#]3^c[^gL_bNU?b_;IefaO,EY0;
J05=4<,=_Q#,0b3MZ/g(+W2#[>=:0aRS6/A]##B0MR[B<^UPZSc=>RdNLHaO?[BC
1+<65T>Z_&I][CMLVC1#JTD:1F7JWRPFKFFg>[(PcH.KYCeJ<e6J:aGO#T.W;BSX
Q7f;JMCg7YSW/\[GT53/A7/BEM2_N=b;;f#9IVDP8IFJ\24+?AbJX^SKcP-U\aF:
:NE;HXCOVU>GcGdXaC7C]9<N/V>.ME+4+a39J[]Ced;68^^B:4[bZ+KM<NU,MY\B
aaQ@X&IF=ccU4_#gUPfgLB^-EZ:)b]8+,IRB12FH@KR<ZQY@C+_85H_(Z/fWfFIL
A5U^<4IWJDWH0F7.R>f1-;+CVY>aSQ0DWUVW9L^BAg#QLJd4+P38GQ[/1\+CdK1.
cMEBCZ_]/DOSa]<]aPF##UDOa\6K],>(H.XKYV&B-8^^70F5T9LOW\ELBe(\C4_Y
[dC\_2dgf?R)E=:-?>d>b0D8gJ4?C)H,@K]WLQEJ+MMN@J<T5H.8CE[Z^+/?&7V7
2)&4_&=TL:T=Mb;D^_R/gC),c3-gI<C1&Y450-Hc5f]\c6]>H1<XQ2Da-+\O/4B(
g6CJW/-81EZL-=aFe=f4+30:?)b?Bg1S3&ZHd##Q94>/KQL+GSREacIf;1eIH+0G
CCF:,>5N3K/S^a^AXW8E4:3U;fA=,,</#fOZMVCAfQbS6NEG63AJ9.:D:aH_Lc5W
85RZQRFMTAJZ/;WMcOg0B4-I267/40+JFNX;(:eUYe>>J];C/8I6bdCgYW/2QdKg
KXYHP4f22:/HL(1L+c_TH,MD4=3N-_C+J[(IdfY9LeG]eZAYT=GSQe+bMX[aU1JR
D8<gFWQe?)+JFGbEb-6NB4(\LH:[X\gQZ2:\L3b@-J,M9a;-6c.4W#-DM[_Q?L7g
#fN#fX[VVJYfRMODfg(POZ\5(:++_7g](WD7gL)1Wf\DG(gK#<EZAG+TO[<[D(34
c=J#L@Y8G=]b4#[(O\8.Jd8UKM8fGV(bV^UP)Kf?e3UFJ-=JFZ?H:.JTCb^cB_e-
Xb?NH[JUNI>:<&A1RYYdTXXOPN1O#+O>2ff=8KH_:28bMA>?.U_@RUE(5,5(TH<0
gb?HWXW]64E</WcC,)3[d1cb\;^S#/,g]5fNT+N-^MDB\O,\J/;LeA/dG+.gY@(=
0[N0(V9C]&J/@79HOTVe:EKKFTQ@D\<15,)48RW84CBM5D50HI4DH5Y7A]D)HPL)
L6M58f=^^;>3^d\XLC&W(JPZ#7[+&R&#&)N(#[L/[H4VHKM(=F5E2eB8PESbEcMG
-4>F;KAc&+<./WL?(88.F8H(Z7GLC3IcE;=.VZI/aFb:70ARD;FD+=+B0Y,6J8Z4
J?6V>1KL1^>-3WRa&Z^P+@(B(_d#)SgDYGRY^,X./I)R<cO=-)a\ATSY]@XAEX7)
4@8&cUEE3&37RW5/N,7H5-<GNdK<\9gJa/S8<B@D^]CMX9VSUV9DP=?QM<@83-Kd
VfA+g99_QUdU,8OCM6L(UX4gZBPf&,I)@;ZI(-e#-,@gK6fPL2;=MX?<(.X57F@,
[NITbP;CX(#EYc&XN#e#5WP_DK?&5&\).I6dL;H93-V28-G;#?FU:7_J\Cg<dA&-
:[-O^^FR?T.1-9J2>gf^O#P@-=^=ZWQ:55:@U:3I>ZWQ<WgP2@;?,T>e5>]/H&DJ
D8A[.;aBCR)eCJ_E(0=R/gVYJE]J2RB2c]Sd+F,L.GLUc#0T^KCL9ZC,gKK5Q?8b
+5;^bM;[WcHGa9][GgC0<:2ZF0Pa8Q]#-]9a[=NR,>S)SX2BXee;C?0?X:-]Kaa.
U+dG/F-3.2]6bMA2W]8SfTGbcWgK<4bbVL#]@4XQIY^,F[a.A?b@Y)V2-7Q<d2dR
D#:B->N#-DMdJf1O51NJ<GgM03PZPA2\NZM=f&J:)Q10M5ECd>8[XeL()26.9R:5
Q&^//B\9UGX.KY&OFP22P[4/IDMTYe+V)dUT//C]NA:)=J&#PLWOXMcD=;XT2+Z@
&NEL3X)SFQ;^4C8R:F=5X,21G82(5K-[^7ILQX&QXF(<T#e;_GSce)\fAV<RM?_I
:0Y_+d^CI5,8MX)M@_&[\KIJ<gT=HOSfbQ&2>a8Q78BU<6D>7KRY3@K#.If2P=8e
M6?dG1-a[B5^KbDeQN]626_dM4O84T^LY_I3f1[[3T4FW&250][E,e#cc2AWfIOa
0&,[AN-EEC3/K+&ZTS:>J#?dc9H[&0Oa]D@=6bF#RKWG;=GdK,C@GA;W[S/YT3E=
U3/G:Nc65\L5YH,^(_\EEQ@4/fUS?1PG#d3GID2+0ef6g24K#c\f424bF8TUDUM_
9M]7F^DG\0QTDJL)=KE).N_XMa5==+[d(CHA(9;_RXaON?\+V>,+^V=@QS>6Z@:F
D4WU:1.aJ0G.MU6?+aPZb?I3GT.:Fde4W#Z0OFK:a6b5#^4#6#&V[-2D/3N5PW3S
).0cDOX:8VVI,C_/FQA6bcY17(ZILdcM?g+GEV-@+EVg4&/35WKI-1[_E^_bPfAG
XRdSAKg+(.P&T(1UUFaA1T+2]L;^g@.FLg416L5HIYd+B;L2NX_C^5A<e<4I>\PV
2_egCa<ebOH0O06&C^)8B/4+0W-:GC]G7SPaAH7CQAH5DI;S.@:e>7H[2I/?XQf#
d+fVG<(G4D75<NR?E;[VeKIdJ,5W0T-,#LG@0ZE<b+YdM@g(XFWYYdWHNg^@2\?a
=OH2ca]NWfK=^AUKJBZ]GTD=]\dV4H)eMLPbe742G8+JcUT:C6\#GIK89W7S)(EL
/B&K]3#GdC(J^2ac4Q6QE8XN5VBPKMMfDfOe3LN.4NQ5V[dCA>]I;PN];.#P.H/Q
ND&;ZO@9<1Q__[SDMP.X]58>ab5ZM1,V728bMfY=H[#[YHP_Ub87I4DI=6Z,;?A6
G7B;U,\8(e,4@L1eUO47Z-B71Z?MA,D02<2(LVU[0;KUEU_3I:6e4.^1:W2\<K/<
fR[2;3Z#@;/)K,f)@Jc3H490QNM#V,+R+DLLIK>LBSX&5#83F+\1OR7cOaL()0+B
.[(fRHb6<]>ge:Q3S<60O2cCg^Y=\cAN?A8Z65L]c.7=-4@SITZ<eII]dA9@LYLD
\>],\S77-;8K_^#;A[T87ZF+.:8<-e:ZbK9f3aS6FCZ[g)1(bI6J:3DcY0JJG(^-
1NWCa[(A&X\WKX<438)>_^?fQ^gEfc99^8O:W/M?L0HNRL]#:.+VH\7_c-D)0@^-
//RCK<.,=?1B4TVPI:]W)#^1JUa/Ld;S\>53-GX=>/1Y)T?.TVV[2bI\4K0fAV8H
\?6W>X4.EY9<0>KO0Z/JdBA3>\f2d.7DP3MUg-#GB#R@d(NW@d&Qb5.B>96d6_M(
\;9-4,X3ZBfNDeLY+fMAFUQ9DdT,CNR(Hc77<TJQ\7JaO9eRPfc)=(U6S8V54/0M
I8f;bHA_+d^TCd_,c(I;g(X7PM=Ac=\Db@4a?I0eWgZDR]ae06DHL816QG:EY(P5
#H</-:451;W7,N[-56_6^XX1T;O=QD0f[:M#>,/f&<5-Ld?)c74c&g@N]H3-1-_U
AY0)0@5H.Y5>(-(dHE4<]DD_K,e9g)a]I,?HSTaV/(6N8LC[c7B:_YA6@f7ePC;g
B4DJ0[(4E1.(^:JR7AD.Lbd^N.[ML9>\Rg1@0fPQ+S3>G#APBM_[(AD#c^@,VGQD
F&bJY;=T>8Lc;+D;f/?I71.71M#BSZ;5,1F5[G+De#>E5236eV0AD8Q)T\UDcD],
35U2/&]=OOG)caXb@?T++<_T^:&UPQ:T^,][cL/SLO/d30<3&\>WCTB#V#Lfe@Q\
):B;#E^.Ve:dE\KZ0NJ-Y:N6@ffS^Gb5X,78EDO5:feg7g:19NG?\9=Z]HRfUUTe
Qg5]c?EXD4ZPebc/-]66,)@)WTVC&5.&1H^EZH]LVY6dB7(=EFER:QS)-b)^RH(6
TW_TN)W-G\_O1b>_HPUMYO]POcY[0-GH)BAZY?BYJ)U:>=VF_D7QLR5]JL4-N668
37)EH+]Yf[((d9Q0H5QU<>FU-?ZMP;EYZ@fEH6\QLX][ZZ7Y99F,.7H)<V;+9H3a
,?:<5N6^25d7HG.\]P]9P48)Q_.DZJ56cdTE+.0UY6D]\a95JO?A=Q3.@dX0d\0@
\ff@g4.A6c?:?G6MMA@.]7eaRRc-\-B\NAR#WX^(-KVP@E:_:A\7@\c;+NeD@JYJ
3]QLFC(J-ZDA;(VEULIT-^U0#NX]+UMU4Rd2_GYfbTL.OW\C_(CBWa07.==HSc:e
_.Q5;VQ;I<,a?eT#[:)H,_g?VW)7WfWM>2IfgB>K)9f?1@g&AbUM>?Y]9FAEJg[^
HFIW(aLc(:3/E2^9>5&\M0YaIJSN#_@<3N;58;EeP&M&BJ-:c/P>KK);=d0;TX36
.L+-@cLD)Y>]_b8Y[cE;D052Ta(I6RT5\R-4AP\(Y)<P7LSH@(G018ZOQ3G\^Q)+
PJ+<J8aBZC1(#@6X:^3T[E2YH^(C.#Eb.L1O?2>5289R,94a5P3_?VD7;JX1[@VZ
d@aGd;SA1Z43P7bB;RE9OLT\N\6JMg;^+I7IeOB&IUZW#5<QdTT9_b=[ZbX+:,90
c[5&3WKNaP\0Z?QX]-(BWIS7(cQQL0O6V&G)O^VNYO#,05_3;RI76[TS1Af&DR:f
.DI]>1[\FBP15M6JMaJa1/)I&Z@_H^^X9QCO)/R5bW.:OKS?Z(+J]VV-X3VGc.b]
?ZS&:a4IXW>:(9-83Fc@W@5P&FD+a(9WcbUM2?&HJNN1P.H<bXU;=g/IG&HIC2U+
)bg=dA+2-.((8.RA04.#(W>G^aZTeZ)R+>FO[3\K;)Lg;^M031^U85)9NCJ+;YJQ
@O&;gA.53,.G208S-Cg_:E>18VT.XF7E=<^IAK:ST.^:Z@fU1]=YI,SH@W#WVP:K
EG-^Z?.O4e=APaGcUKU#B__F5e]H<@XU]M(OWO/d@L:,@1;J_,][ABQSD18CF5WO
N-/HU,4OOLF-X=-+]2P8K8[c5Q3]I?4c/^c]7^S8EP1?U885[IP>OBM5DYL+e;=<
Od6-5.V1]@dE?3V>@bPKRC2SX04]BdC#OMR1/&<Q(2?@N=]XY;Q,\gC_E4QU/NB.
?^3:P8H]D#eK;4.UaGNBXAN/>P92;7^9)UWOOM+MHb?YL#d,?]V;U,BJ3PISNf:L
^?C:4:5\<V/,Tc)=528(B<g<MY-<(ZISMV-M-SFDXA<:>eFAIML;a<KY)=4\T@+4
/=,#gZF4Cf^0f@J?48+K&[TO_3JbTM.,C.N=<\E(UcY3+e8\L<)M<(>WFMb+D)T1
PA;0HLGgXQ_=TfY7FgQE=GERG-fBgf#J6O?UITAd.,gU3g]MHI,0g+QB1E7#<dCH
.VS=BON1D4.TJ?Pc/8JJ=W(YgY_P-5SFbPD7TR/2[GR/0)Z#:9ScK3L07a#Ee9>T
[gAC?GLWf,FVfE#^9B;&+AE?_=-eSB<g+fg7BI9RGd3KY_dOSZ)gE_f9F&(G]+\W
3e0[[f9V[FJ:0IJ&eR<>9OHA[A/,M:fW#Q)f5)KDB6:B;HN0+64dY+DGNK\]:;Mc
CGfAOe/_W3RdK=)RJDdBSaK5Ng4?eP=HB&Za4bc?WV,?/THOYde2/dZ6g5dNTcG)
43CC^1,TQ?<PD:7OW8L92e_@WV:KJ\9-^@6K2aVX]2DU2=[8=TR^98Q-&PMU.bPe
;N:I9(Mg+37,>d[N&bcA6g@Bba8,7c>2<N>_+@WOQ68ed5A:N@[[cZ7>841E:=Q&
#U8^bKNJ<D<0?8PeagdgAEOJUFP\S>/Qd8JT6aS[4Rg,=D(9##_X<D2&561^FHgT
&NMD;41MQPI#8MWJES6BcTIYQO8@L:feMS^@)]>PE^60IUgb37VcKgZbLU^,\?)2
I7GP+L-;3SYDeJ6GA>aZC#FPOf?SY4#1\;/NOB6XaA]5QPb?3&B;FS3E[dL;YY(0
bfK-=-L=J62<\Z-aGXE3<CWO&Bg-fIVe;J#+ZGM6aV+f><^V>.a]dBU?WC0VZ/L>
>,33Pg<-6b7aSb3(5OQL&A/],+FY:NZEOI_Ogb?HLV(I@e:-C7.dJC8NMS<a?#f2
Z=8E,Y(3WVbTa?5TS9.K+45EcO.Wa,V.-+<@3c^0-L4QbDfeFZ1YLb_PICN1F_M)
,?ag?Y:)2S86<,c[\P>dR4.b4W5Td?+=05>A/Y[[6gURYfa9/#=M(:;&#2:E+(T/
Z>0@\/aNGA;O;RRU3R&9,92O^>=X&5C.MO5d_H<2R<K3>cLcD#Q4T?@N[=TDI2+S
/c\O?W@Q6ZABeL4DI\/W)^N3DI,VTVfDI004U6Z[/.TD;AN\-Z7\B0(T<Qafc:KT
7R,0=eB;=DNe@eO5OK+.f40I_)R#=Y&5eB?E5Xb1b;Ua_V7XX?U&IL?J71XV3VV+
)D]+DVN+3O753_a-.gR[]e<<=c2XNHX2_@<+]RK7Nb@-ZLR&<P,6:L8(;T#gV=M@
eTL--IXc;D9#JF2CRA[0#3>[IJKD-EM\Z3VW8[bX:7MSG5/>NJ18ePV5\M==:O)Q
A17KJSO48dB/UagYgU(5MQJ^26EV?H6P^MSO/_7B?:f?734(#0BJX/B7A:XQd@99
ZTQS&,;JI12UZRC41e@VD.\4^>,55<YHOCO5IERgXg(UaD;8X8YVC4ABW(1GJ5/\
#14bZS+E46<a>gPH[OVLIA1eX,6)Ea:4[.\f0^^3I3:c^<_<Q-e#1KD:6XG__V]J
#[>@>F/>)HY4)II1)RSPQWMDb,2@O\Jb/D4dL_.38K-Ad)=a\e=Y6/aTFfMg;1Bb
UG)R8O8^UW7<b3Q,OaYY)PdIG5.B&bF=#S8-MRG)bMJNMb&QMCcg4;OfAMCObZU=
Yd;4((.b;/6@P1eD[_AN=_@:Bge8b([=ZfX?H9:&F.1@5Jaf[BZ+FC5D:8@]QB3X
VZ//JD)=3Z?T-Z5M0fd)M;GeMHENA.B[Q_dCTOS6=d:))RAS(:=0&gFJ>R>&-,/0
)VaEaKba[IGc?OP;)&[VNK_,CO<J7DKfQf)OE<K>0EV16a>/H+fM:E?QR<FZ4(OO
V;Zgf^Sd?.>X<34J#^N6_aIY2>NdJ\>WXOfe,4g?7:K\6&HCZL8b9@E+a&]?QJ]K
/B1\B4=2M@)M)]5QUD,\E?@J.DCWC^[:#9FGA?@A.H1B&V4H^aM0YUa_30b66[&/
S9>E9AO,4;MKNM.1^0S[8J>(?CQ;aU-7afcGCJEDIEV&96E^2[\@aC1J8c[RgJ49
<a&]QFK_\[XTOaZE4J6AC7cM(2_8LG&DC3@E]/39<>);,g:4@LDHC_[>N:H\BN2B
_6BY_OPb>S[9M=B.6X.[4T1?.d42DGPbDMWNXBR\+8\X))a.8a<+3-1dUL9SHU^g
3/&M=g&>2Z3-SQb.?AEHNCGV+(>O0D<fL<?K8H=PWdE/DZgD9dJZ-H:J^M36RUVV
UNMg),d>4L9=H:2,<NW68L>YQ0fTK2.)EB+-[DB7YC>.SH0X8?PS4;=b]0-2UCY]
RSE--@>01SWYU6g:g)gV8R\=7/Cf)]I<V\QMU1b8\;U>JN^<bZX;45@.D3VG(IX?
:e?TT&X)8:@&f>I4ICET&169EWbB2-MbT;1CX1,3FJ?e?@?DC<\bF5QCJ8&+#CNP
,_cP]4cHgg(f]IZg+d8R0]gK>@\UG&f7\JO2N.g)^HUW3WBbI,^b48Q=/fO0SH0[
5MO],9T&Ya)@T#b0SOKWOMWgd:>VU3,=[J?&SH6Y8=-??HTe,-@Jd^e1>L^1fHUO
^=P7CNMD:JRH0M<E9><PJC+1^J\\^)fZ[<3VCaEO(0HI0ITG(F=O,5>CC)?a:/11
L?9TCe_)JI?M3BQe3A<UE@R>[KG.bU5^ZX^1&?Y=NNUE9dRBeXK.M^?d(DG<9c_&
e0/R8PN>4OM@24(?;NO2DB-HP_4+OZedc1[^9V9eULJgaHeA&8PYG:TbG?C94ENO
02dgZWU/3dc&_PG936VDbA9252DL3A=2CBb5e3IR\GU4cW:_G@A#(:]R/H_GDF1Q
c=/KWD]E:Za4\>[CJ=Q3/VQA/1R1.U(ae03CMWN&f#&Ma7L&7fQ=CgK&\3F(U&#2
g#OV9R0(IO-N8b0&>b6ZgL2HS]^XA#/2W,8)Q&9,XNBI826/DGB_cdd+380>1L,M
[W[1f0&&ORI;YFKHKEUc>A/#Ce[@&^@Dbg+[)F)C(S8TNIL8b,7bWRPf_UR3^EC8
BX6(8WS/U_a?@H.#(TZ8MB8b4;JUBcRJN<ABad@LRO\GBJ2L9K8L(CRcf_dL0?=3
[5[KKY(K<XE1CUN2-JQ..S4J]a\+RC;@>C6TDc,9\E^R0/8YRCHF9bGB?N&FT9?O
UbG9NHXaaD3.H1f4X+9)7VR.B?d,HS8L)D_8^;b4=?4PML+6:^]aAaF((Z/H]adc
d-V]fY2::Kg<)<=4Y?-?0B=;W:9Teb+V<Db-dV[,?;Z<MF=62=UBSc-3?FPf4E<(
))1_D\Q35V98V+=3fRZ>b:#=RfMXJOCSWTUR3R\QATdLC5.UL@]WEFBB.daCaa\D
LK_6JD?/^gSaL2NU2KGL)\@La#T.=IRN?[5,Q#5,D<67feFJ,VMOHWSCMOFG:,X1
J(TL#MA09UN39=_R-@9?[H0WgDd2a.#Eac=L-&/O5<;S9XB5RFUFf>S83D0PdIID
25RM@L6),45;W]I[[R7[>PWD]L02N0d76RE]:6V1K1DcLI#1C?OSQH5<P52&68,:
MaX;EJPI[U>+QJ1Z9I-)8QL-1(f44?7gVT9KSI9;_1N&MCO@a87_USAb5I<Dd;37
CG+PeS1E--.1)@Sb5_J(1+FD+&&bNWb<421,X(dY15?_P</-g@C:+edP7WD.MMC<
E^#S5,&6KcX1U/7_,8g_Mg5A^#REDIO#g.]E.6Zc>CR79gf1;3(LMC)Db,Se:?Y@
5W7_EE1FX==J&OL)ZFdXUK04Y:G>MBOL<AS;@=gf92BMX>1U1I_4P<@3[E_Ve5E3
<=]HA#RZ:7_RgR+XK)#)g1QdB8Z5EIA\+M@d(^@X6fAHF#;Z/afb)#_afaN;f=5X
cZH_OX5CfTM,cK9cJ9^]GCF[g?R63(<>S@a&2>;?d>eYG>QK&Q37Ob@f]g@8UZAY
RDf-R:?]^=65OQMD#^_]Z+[5:#A2)1DaLGED6)B<E4MCc;KB/KE484c4&c2MbdN]
FEUT5fGW1=IGKH(W?0K.7UAC&91-?>WQe1^[9GOQWA2P4(3TT)DOG4+Ngc234fTH
T3JQ+O#+NVC7fK,XG<CL1_WD2,<KLI#6Q4UR(7)ZP:B5GK>=9=V6S=.fDDb)=]UA
B(d4bJg^I&Y@d29BZ.MeHS]66Yc\4[&T8?EO>UI]:7SW+FJTM)@J:6WDMUfN:=6_
]J-W#faVQ-V.S3F+;fVZD\cFQS&L&^_#4^?8^c>V2I3Mb(\_GP9F]ZMaaQ]Kg[#/
@E:=)\GDX61>82GO]gOg8L83QcXdYFfMK=XfB#B6?5dXOTQ3,#SD8:Q2W8XDXeGQ
-9]+1WTN;Ea38a/,fGf0gF=P5#SVB)aNYB-;=CdPEA\FPdT(dQOYT[AFIOYB[]X^
MV-&6(#V/W@dg.Yd3>:5f>5X-][-:MMQES[G7U.dHdE@ZC_:+89^>]=G;)AZLTcI
f#PX6TKX\RG>X]-?aYKH>M/;V5E.I;L&3,7f^eTCO?O/#2R\ENZUB5:CTUc[f/<5
X3ZUgSOMQU#-YUJUALF0&>S6^M+d?cMP&15&V<+Jgg,<Q]\NJS8J@+VOA8Z-^f0Y
cOR^,H31IVPNEWWZR_UO/#^26LNTC)[&@4G-=;OP^Q_Bd06;.GJ+N=KT=c<80E[a
T4I8Yg5KK+UU18aaP<52dSE4UdD[,/]&D\=e15JK0BEKg]F/@dSYY>56?]M1b6VL
6(72^K&94PSW-bQMe()]Y:?W;00A&R8ME^bLUJLT?>YEHfY]cAZ;&dPc=4?A273b
CWNMg?+2?T+:_gG8:C5>_R#/NWVA1>Hb51/1QLWY(eG8XEB6R?RcVLcENgg]Db\W
S3Ie_VV2HU@9Q1K\WU]RH(U]-1GL:C,Rf)-^UYW#e-(,4=7LZ./,(NU0FH,S3E36
[C:\Kg91IP;[8[4N)bS24d=:059DLKS5+FaP_4\Qa:[d&BNTfNRMG@1OMfB+;7R&
:G<5[.Ib.HXR?P@F;F_c@0/f@:PLW?TY?:R>M#/T#1WCN-4C6SCP@;D^eP^,&B78
)GH+#XNS-b=_JHQ]M^TJI,MD@C\B0SYcB]W+;5A7R3?Md#gIIS/HTFY(<88g0^_Y
T7[J<g-5^YX+L6^:=?R=S\#U)OC2[;IR=1SZSKJNc<9(8AT39+3AU&KT<K)?DHWD
QB,^GC3\JA&UE0dQaOA4[:U4]IUe2B:g2>e/#4@&H\KB,IXEI.-,b#1@0P:0TARa
0FFST^bZQ-g6@S?#5CV\-G5UWU#feGB_]OPJQ6Lf7])=f2S6Y_HMN1HX?6PD.-c)
SI97</U[8BKX)eX5,8LCc9XeOb,QNHA_/7Ag&H]3a^N0N5]LB0W1>QfYM@-)26S6
13d4aN>gP2SJJ(FBgQ:&T&^a4DF3DG^d1ZUWHdNUWX>B9.f?O:/VYg]1:7?Wa:)P
@M23I1L?:FHV(?f^#7OG>IS^Z\daG;\]DBO+>Z-FIL_>8acF94UX#e-Z70V1Q8R2
\C>O5:e0-e(e-<:8Y>189&S5a6A3[EdLJ)>@8CAV/+-,UFbZ;a+JH.S>[73Y693J
Q_[6G/KAa30D14M>-1E:))VBFTJ?MA#:OEM)R\C&T]([R0?gePY\>d/FL_;M/43R
^^LFV26ELJaJY,[.C8[3ZF-A-VE/<&g+ED0VbJP@L3LPPCJ5g^BEbfaeMVfb;R9]
#Rg@gdaW0AB9)(+C.Y.BFYWg4E&D[J=R3JbSP@?,_L<LO,9@^RfH;O@bN#;-/5X(
+Y+W(S&ATEF,6S/S[[\Cf#6G=#MR054dA.DDc,cb#c)#caI/GL<FBBH,H]I;>D_]
TGVQAZ.S][e=)X@,fRb,V14U]4WLgfW#HKeWRC3bA2_&GDD)IJa>Y@:;LOG1c8Vf
:I5K:^2bGK8[?Pa3BJ71dA)4(2PLHYV[5J;QbZIId#ZZ&H6G=7ZLcSN/YL+)EUB\
_Oc&eJ\MKK]eFYD6KPHS.Y074&C?G0Eb(?_(+PbV4Z[<<bRT]g=WD32-?=W4aL;M
+UQbd#[O_/5MOT87E,,\T@9IC5Qf[^b8,ZJM[KF#TF8N7QJ86MNTPeZUZ>4Bb3SD
dKF_@7]_@3J_O39XR=[M/d/)F2[a^eTEC2U[IS)T2^->JI#[=)+Z-CW>IHMJ9ZO&
9DdV\HQ#W[G0Y-T3a+J1^MC5Cb=E+H]5?3O-H#.ag,X[EXOK0(&5\K]68WePIcb3
A=FHIO/]..RF@6648Z&3?;+/MWV5c=_e&G<16K^QCDd+]@8VceG1NTAb6=1T19):
.F8.dTV>,]P-f4WIXWAbYWX#\?WRS<C80KY+_f(TXZ2QQJPP=D&YU^<Q,5Ec5/HP
6N)c^J#b=1(<7JHbA]E/C.RC34H9;7dO8\+J-PG+L65[_^06-8O>>)@d>\OAab+#
K5d6]O6Gc=V^Z7.N(T90e/03EYT,P/+DB5fF>./]7ePV,N#QVP8=7A5c[]WL,;6Z
;=^;.T>7e#c54;?&8UD]7-TBfCRH2@c-YX=>5^3@S)TQ1D]d-L[A#AM?=1MM[eGZ
>-.B1H&/3Z,U[]c_WJLJ/I#WgYASN&/.:C=1MD1RKVBFXW3Ig9WU-MMAX)>I@TT(
5DV2]U4dL2W5a^A?>.]0e>A.C<9G.)S>P-gQ/e;RU=T[CEB#IN?b:&&4Y/>DbNb#
X432D<CeV@0I[2g(cFgg_HH2;]+#SU(eU#gLCRJ#5Q:(J2c9]Kd^Y>5KX,[TI>6D
1QRM+W.5&)BU/O8,K.JC4[eA4?E070+A^0O+=KW,=A_Fe480>^Z8@.ZbO)^Z;?=>
D:\&0MH_47Ra(Wb=F-62eRV#P#eZ\+HK=NYQ?@C;2V7LVQ7\VE=,D2c3/=4Z.(Y:
^1H/L#(<[D>#Jb\).JX(6)FA:Q3EPJ);\e\#F@1-bL;W;W4HVULNE<-ZF1E/)eZ7
?fXD&9J_#(2RG@1BEdS-+E5R=5\L9[CT)PW&P]Q&-GU,B>[A8e/4,If5b25g(8VP
@84(dLJC.eK/LE+/K/Lf9@>X,78=GQfZ6YQaR4-PLV.=NOJH@+GRXTE/EIGAT>.U
AOA3cScQ+X5Lb_;UD8P[1Z^JDMZ,24ZB29H-N)R:I2>?_W?GX9A/W>HPfQ=T&gI;
aAMG/T#07SE51GGcOc[L-:&,QfUGgIYR2JB2/HaF2M/QS;<c[W&a@)T,V=J3CBU,
@\4HYW]G_c4[,NPf+:TQJ(D;>dUTCdR61CJ[RZY&,.81\J&]DDM0LV[(ATG_/:2K
Dc1[^CF?DFPG.[(N)=42YW<S95@(9XWc0gMVbA=V1OIAA[(A4QDaW5O>A4GU)ON6
+AB;)1d3I0HSLR,5cf9+@=)SWg5UETZ9QTb6b&DA_Jf78EA2e_;5+IfH\XV>S30K
B@(H7J)>516G=?7f^d)D54R,>TXL^^ffT2\6Za-\8)P3NY2RFK/G[@\J66]DK-Ma
Y_E+bfY3AWP6eYN)LV.JS2#5Xf,c7If&b8>PA<?7_)V,NV;&\XW#ZZ&OE?5AWQ?:
)K#:eF8[;:>0+BCC4WM_T?BQ;3/@0?aPK_P,(d6/+/\Q5G)X@bRf?\00\+TDJAM5
N<J:[P=fN/9,8,DaU?T(^cJ4^NaU6.d,+c:@JCO8.TY?\>,BZfYB9]R&]#FJBC;2
R7@C5^1(eDZWRBH,_<.O<d4KB4I,1Y=<KTJa31T^:dU#IAAee/@@WRER\6^5c)3R
VPR[GBA-;O219YFf)_6VZ@,5>/VHKO^L5VC<;NXd00bUUg?]CS5(Jg=83>]W&]&:
;H[03+dPB-_EA=>/G^d,Mc\&5WXL58J<Sb6Y(0K#b=ZH^\2[Za.>UXbED\E?057F
RE,0]:b:QP2BSDe_)P:U#ATU3bJ<_[dU0)PJ[TD19,SDZ]C[DNe4@PMOP>PXXIZ-
@-?(_b]bNJ,c@7_#.?X:OHA.U/58?c54/+?69QPHL&M1MWC7+K?)d2I]R;=X_8@0
N:-<eAeT,MU/B?:(J5Ld;9&<Id#QY_(NIV#]bHeB,(:=1\&7Kb2YQY1AFU?@=ZB?
-#fIQJCT+KPT\bIV)AgaWZ?]J)aC+7T7>]S6Z^SaLPAJabSIUfZSOeKGV3BD<X6K
0FR95M+1-_5V-ERd#?7I(S=Z[XFYG1LB#7AL2HWB(+ETaY.2AFF?<4_a^f9e85a\
e@?09@/KIU8X>4;L;J?6X9-_T826QD6<fWG1XO^TSeWVX529<GG7;U/c-L+4Wg1A
1#\7T)]bR746R=33(QKT>F?7IWPbPOHF]C?[ER_4[?@2U&O-P(K;J#&3-YU^C;8N
0b@d?+P&I^M[,(N:#KLcb]4.cQ>b)F\YaZf+8a+?EU3<W(4ec<I\\,O&8TH8VYJf
C6cP\+?4P3^PgSYO8]K]@2WP;1?ZL)RJ+Y>T)c@<B4aBIBI>]7HO;A0EbFA(T42D
VR316030]+W]7e#?L;c40eUX_&_IROIA.LF>@DdWQ4,VLJ8P8.:gVN_<]M&3R-5\
b.E-C#SCSZ@EJbK&>(->@DeX5+\VKM;FZ95]GOd0+@JQgD6_V,c(a]9b&2E@BZD&
E39@E/K<@&A=+W:DB\81fcDGOIf=J4BBZ]VFA6+/^B6=c&:6Rg>?\Y9CV-&=3(UN
T^VPXR9,/UD(-ZG]JC?=/ZL+CJDe4#3IZ06eT@LeCDJ^1JJA5@:1/8]dZG_=XRKE
L7535@?S1_fJB^X-9_/\:FO[LHaK57#M=^)NdJD[Vb76OL_WMNcbbCRX<J(].4KW
Vfe@YVXM5R@4CGMRW4eU__O>,gM^Fg(81Ddec6e2bZ5>=P&/Wa[FaWPPZ,WO7[2P
NJOK3c.HF]&_<AfEQO\]]:.]\D67P]<:/XX(F9:V3M_S?JT-M@2,)93X2,-+Igd;
/S@&U3FGBKQ>V1&4Q2b_AG6-YLRe[)1:Z=8YW0Y08MVB<9F17GeG=+XX,9P>A<8,
6HTBedN5SDGac;958V:8[:Gc0.+]b(@M@0OE6S\=D=K](b6,bc7E+f2<,K\ATU)D
f-YP>^&S#OXY;ZHC6c5T^,\MO.c0=+/7G:SD7-PHK.AdDV\3\Z@P0\Y6_=DL^470
cec_:JMFXF-Q9Mb#2f2YF.13b>dQJF(]&/2:NL9UZ#(CfF_/D,CJ<YLL,@fUdIKc
Y>D9/[b29LLcc,K]B>J^\2>9LC^807>Q898d:P:7VUg-_^P&4aTM=7g[[<gIJ<)g
-e^Rd])0X:?4I892K+OS24e?f<KUeI?(S,f?\JZSgZ0VOWfDYd-W8?OCO6>?.\H6
\LE3UIA]Nd_V8/DFLU]-?@YD8M&?0J<_ZVH3W.6?B;YJBE9M1TJ5YLG#PI/cb_LY
T;T-g8T^+,IE[7O/>4.VPB&4XX;L0O36Dc#=9=)]E4]L,Q))@]480C.4I:V;:N[R
2PFa?X9CU^H.6Qa0,-(I<J:E9^P]?V4^YUQEC+9DgO(?^)KKID)6>YN,C)/Ed.KC
UQcYGPR-&G=2C-ZLA)1@ARd7edX+0[.WfgF[b_S.&8#-:)]]V4PU.I#[HC.JYg]+
:Hg#PII.9:RU)I8FHKRWbKU]&^dIC>>XbTQGg6Eg&YAS5[662C]#0W1/1BC>\SU-
GbSX3&L&Ic8,6AIPYYT,#8\ZVOE9&5@BLY\#CCMD]a2e6;0L?[+8<dd3KWgB]S83
(HU<caP0ZQ10a^&c/3NFY>@(2X<DH20bATE#NXGQ>dMZ2G[9Eg1N(3CF0Q,>.A\:
+)4^I8Vc/1#]&fXaeCP=A=H3-E3/c0\A9UgSbG(;Tg8RJDZ4?3_4&5BQfT:5J=IH
21RCZ)+[@_5cY?e./RENY)5XSX/Y(c7IJRE#OC8W4ePQ5E1E^H8g:,D);b3I&LZY
?QUL-JTJP=K59->1G<?N&P>b.Y;Q@IQ2d<@C,=>Y&](X^9(M<SV=cDB^_V^RW8MO
[IcKV7BUBd/2e?9_I1L;VG\C^ESfEK@XB5)8UX5A2RY5:18GF,X<00aa58aC=_Uc
]LUW@^C:C9/1V7);9KMMc;YTUBP9A_4X;bS&AS<JFFdQ;..5A>OJ@>.8A0R>=ZRf
;XL6LN=4VfQS;SIF_W.3g9MYH&@78^?#0>B;[d+eTQZ<?MAAU\/dg(+6:FO,39,>
fAJ8.MI;6F;FM+0fYX?R9Vf0Lc4CD@;+-bU8#>6+U+8g>I3S,DOT)-gSDB/^F<JY
#f+(K;+X7dO:D)R+W#e:)850ORQ(f9J>b447SggeI[SSLFI0d+_K<_YQ-C+KUQP^
6#a3Y-.T+^;(aVH\R+)SL>N^6G(AAOPQ@W]?[3&D_#>Sb0E2YI)&QN;AfMPLca@]
3a6LdZJc\ZJ#,ABdORZPD-GgA077c7g,-^;@#9KffI)<<3KG1+&QM=0OZ1TbKR47
f82F9Z3QGV6ZeN/9J<>:.[W:D)\Z[;aB+3@U9JGd:>BAd+,g<5H)UeJSKO8SJ>fW
fAXd,5D2^7HN/ECOR)](Z79?Oc7I-27HK^f29gFX#A;P=4Jfc))(bPX7B4,=G:\Q
@;+4.:9M??2L5e?#--/aWd[1@4E(,GA]MA-67aWPWRIb)-g.PB3CeGO97,+YXM08
RL:<06H9#=RXP/.1ReF[YVSLR9eLZ[\R@-NU9E#=S9UPAHXK-/<YQBZM>2Ie9N9P
c,;@-?TKU49^FF+I?JXV4:&K+^FF84aL6gWG6e_^VA)/XX8?b[,LH];C#/,XB,g]
^/BUCH9.-?W4GY<//66.0LA4b+E>UeNA<Y]9H,2FI?MRW;IK<4N<L/WM67]\2ZKM
NKd;1I[T9:)F(XT/?G-PN;Y]]J\YaFI&[a#V76G_@K,Y[>LgJ_R7&/):\A,<088D
e3+.,J#XdEdCUR32@(R4-D_P>((^V(DFUK/G9fP<a_2U\1#WeU>d)HC9Z4SO1A\1
ggEGMgKD6WPV(=aY()A.N7:bK5<O6UPFAgAU:+_384aH^UP0WOO7[S2e+</@JM6-
M:UdYY8FE(e_Vf<Ga<_aR,6.N83G7RAMH^APP1\CO@<XFDGVg)0,bgT_CU-R4\6Z
Gf/Gc;DK.?@JAY;TFfe,0[\?5OX6(/?[63WTVR]OIMdZ-_bG.^&:KL]0]=/-@>VI
QDgXU1PSb5>49#_d792a\NKd?/1@V3&#6V^WNd(MRS&W4UBZ6Z\KOY574+V1<7;R
K5dGXIWUQcaC(46+V[BT6b3D(Ng)Q2DXg3^;.)7[_#-JPAQgV>.T2dI1.#-@,1>C
Z[MI6^P:Z,.P+D@;G3D-SL_+a5#BbgU3>d,dCY?c^CBaIW&Lg:8f7TCIM[>.Q;[/
fHL,BfEg[/PEfDC[G.U/N^Nc4e3T=A;(_^/PaMe#6a)OL/6eW-N=YcEJ,B)C-SYG
[P;b#GDD&N41KBP2#4&c5B7#L@g.?>EBAgS0/#7P(&f2WR4L)C^UHZ9#;-A?S:QI
AAAN4(G@0UKZWBKR636C@S<eHg^[F4[L7:?;\S1CSOO:Q(_.F:\:Tg-<@R8-R95b
::O_,,Db_B1>;OWPPdKR/CFf)Cf6O^16bM2R.+8M_C6T;7@)MFdW4K3-Y2OB:UVJ
VD@IKU:@?&[E[JD_(Bf]&;Zb=8C(9^^EF[EI3I:b1C41WO(9[4)5/\M39^-:8f9H
0.^U1Wf/GW6LbdI-UeE^Yc^)(5@BYCNd8^[1.;1.W45a]I=BAZ1MEIE,>,FN=P:N
O+3S7ZJ@g<X0[/(=\^PL79.;=&dd#,Bf0FC-P][-KO2Hf1Y=^8-&TE7N3dgC)ORE
NU(g[dV(0gR32&P6C;<(K;eaMEUAC06-C-8/@-Ocfb#\DS7OPfQFaQ4JZ;5915AV
;Ya:/-TT2>1371)OOSUQP6/X@a(L0d2:W_CF&^_LQS6(SAd,?9aX:PF\bVVc4@3N
<gBUVCF),0K4d5YC&MGg/8,#\EDF0W]S<X?61g]O;QD:Q3\OLIC5-c8ZRf2)I#S]
0,C]Xe0b\<Ff#40HCG+AbMcWL96bg,D<=.E)]#VFC1FS\XEVH-X4aFD;]S@<KRDF
):]M#4gS,)GZ-@3Fe)=PWE^:3?gII;+PU.g^deZ<-5PfDAB)93M).SMaB@NG<_(+
=XbQ/aBW9N<+D)RHbH/DF>EU/[++#,.aY_c+=0P(eE0I)FF6;\HKGKGZd3-D4J)9
;a-PKMJf2;=TO<C9KEf_Ua0V)e_JCD\YI,)^1NH<Q.U&FC+U^K3<NHB5)38YbG72
@>#g^B-/gVg\c9BaVCG_&5]cb@>aP9H3YDM7_fDFbbD36LcW)<1B2A1QR>DHQ1FD
c3)&HXNUeVbdKA/R?7P;R7(U5T9a^63D0ZZOKSg5C.D=eKacS,0daeNQTcS]I.H,
b852O=Q8SaMKPfA7b5ZTI.WGI+[]2J/AfWbGPY]\[:W7LI#.(CQ/:bHA#JNESbY&
)cWX&)KU=P&VF+A&-DKLLf,U:XAJI:#;+<c4(UXZ/RHSaNdRE7C>cd)IE;)I1[&A
#f6@:3J/5O8cWRYXZb6Z<]A7A&EVQSUQ6&Nf7FXC3c_6QT</GCL:ADg]+PR,VOVV
e4e_BEV<6NN]LfYUHLLJ@fY)WAG8401:6X9=).#S)N0[MFCO_OH8BT+D_K[O:2XT
3,/+L=Re_AeXN5f\cfbJ5>>J#9>IZH\;dJUJ3;)8aFd3Fe8ZAKITQ6UQ]WZ4(&EB
VK?[Xb_U14HG@OA[bXdC2AHLX+;[MQC&:4S>MaTBG\5Mc7=NeWR5ISJdGK,R_4WF
ZbN0:?.OUC)Z\05TLMNXGR&.A5.X-C7dc(Z>WHRS]+?P^D325VD:QaQLJaXd;f@X
.YF>@E83O</Oa_,e.K?]bS<8]NV(-))WbPWHE8;5SGFB@f@_E_1/LW>F4MA9EZGI
LcgSG/2KIG7g[?D0)GJM&3fZ1:@[8aI^]5f>3VLD;R-HO&_P?K)#4QFO_S9I#[E_
006)_Uc/>(1/4b;2G4K.;GWJ7Z@L+DR+[I?4^cY4d:T6c.GO+<]XA/]@dJfW1H]]
4L@dS,Pb,@5DB_<Ta#+UY#CDebL:a89RKVP^IH0(NT\;>@6/N4)HeYG7V>=.N/NB
].<XND?9-BeNDZS2AU@fZMXHOP;c&.@D-G,d<U9:I6HIGL_]@<MLCO=#b2e&ZK=:
(36JV0Y)>AXS@BU/G^<UWG:.FZU@(/3+W\>a+Dee_^JLBM0@8COQPCW=ZfGA3]KY
2Y_B-E<LLX]V(]T-TZ<#G6gKDT&QO+3bEcc]\T+HMOW:9G]d;MXAR>Y?<#fK6R8I
H.-8]C#Y(9GO1S@>BTWRQ]G+b\/TbX[BI_M>^:,K8.-8cOC8TP6GY(C)OFE)F1_4
]g?+a?Qe3+JL8;O0@YV-#:DegEdHJcgRFE9J#3.fSO53+_?bR7IG=/#7^/X=:VNb
L6)bT>)_NCNL_PLf7+P3dXP3b:OOH161_g?;BWb]SPUSE\:UPF-\==ME?OFg8ZO=
T>;_GeRaH5a[dH)[PQ]0d5Mc^UI+\-2MHV.I4E@_e7B#NT,NB<+>FGKGcDISg]\)
BG8_\.7Q0G28S)c/c/_LN-H35T7\.cDWG0YVPO&1=6+]SS=c5[b2_\]<LY#=M:\0
fT>EW?<K:>1Z0c)Ze,d;+Z#LKL9b>JaXCP3A\Zf;D]f\P5<]7?3JG&\@#BR-4/Pf
fDC[;]9f=Z4-9@aa9ONYgORBL5QYMAPQQaMaDFZ1bVAEPS_)EUW6>O4NTXAH^(+S
Ldb8.O4#.S7,UFAfPgJ/SUbD6L&ZY&9;;QWEP0)?ePgaBGLe_?5&OHY<OB6=W3]7
d4Q<d(SB?@c&:eY.VZL(S7]Se;#K?-X@;;2=].4@O29H);]A0;)#9ARO^#SY@B_d
/gAEOdIaP22N=f6bY5[KLG_[gUM?Ya.DO41K\)3^6&K)[Ma.8RF=+NdX7)H=##]-
3BCS:JVOU>GQa8)C]KGJ(TZS6^RV/RHR2]N,D^=SeFW)4-GL\?^^WJ;K&2)e8Df(
N)RS=Y7:]@_0SD1Mb64a1E3DRX8[7b?@Q7VW)2?9g7QQ_OZ5.V2TM8)LUdSc4K::
:BbVRK<(WIE,)&;8B+DB[FK7;-JJb8a9O&]eP6C00CW;2I\0R[-15])AMeI]HJ/&
d<LQSC,(P(D@K7V7:W5YeYP3:Vc/HVS=\]9;KIN#GFg(8bAb/SUNY/FSW3?76McB
.BEC,EM2D)U-f_3f@>UNWZJAQ:06#X7&HM^A86N[^T[Ub)A0#-[53fJLGBa3?E=G
,GFSB9U7=M;9C7@E<Wb-4Cd_8[#+(VV^JHR&:((3FZ;DBPZP2,R-gBb?B_a_A6PX
a(F:Y(cVCQD\SNg^_M;A(48bac?3?S>(_&+UA44a_^XeR?5=T_6O_]g9K7SFTfGO
J&acCf4MB&>@cW]O:@H],G2L2P#IG85JBPD.EG[_95C<33be2V:,BF^7aU,dM1Cg
>1?OeUBB4aKNJ/F<bL_2(-WQ4MA5__JK)1,>S^18K?#8(bL#W.SV_(@3PC2eS4O)
Qa92P>.<HFI/eG1:W-K[fg>W\9([.<D-bH8QC)/MA=gd>.8F\\f3IVZ,?[c=PG>0
f3:g,-@C^#IF(QHc-YRD[DOI2&1^<>e(EJ)C2WQ2VO+T2Yb]-/;K3W;OT\==.]&/
XSW&X:Med\.:7&I.2)>.5A&RdL1,F?IO>MC?(.5dGD?S(4WB/W0&4I+b?F/T=S2E
47+^S-[NM+HC>U4[)JGTbfg;3=Q[DD]@83dQ1HL/#:#-XfdZ/X(a+?#I4+]FU5^0
T;_3C&/)[\Qf[J]e5,>DRVYWBJ8F4.IPcW,5S2(aG<Ce)^PK#]dOK,2TPE.]@gFJ
IB+a:ZHP:H_7Q=HI2U_^,)d5DcL2#KS-F@83=&4D-<660XPF,aaP[,7G](Rg0KbJ
+E7QZ1VG[_3D94UF1<N5[@8L/G5#]M&T9W^9gHE-1FcZ.QD6MU#3#/V#27I6(cfe
(VVJQ]NUN(a?\ZI,XFPdcMW^a1YdM8954Q3)ZgJ>b9@E@>-CSE(>\afGK)Sg+c?5
<?[#VR0#=Eb;c;.LQ;)&>_@=b/XccU]MR74MCOZD>X/a/WK:(RB3dHL^Ye\;fR9<
C)9RA;BX1[ddgg#?;+N=6EM?H+4EL=d98JK(<cQ.>42/>(E/:FTLVLC(Uf;R[eT-
YB]QKGP[/ZH99Z)CHN(b+6(EaW+WA<;2Q9M\S<3Y-dKdZ>1cEf)GEH12G)RdH5._
gG&1&&P6:^Y</A/21/d2VTWM1P2<U#PDOO;J(,3aJ&G&Z1;(WYL>bD7EQ,2=E7,4
8g2J]U3>C67QMCOL:aBXb9MQMZfDEVFBI>a?P4MYJV,(S7Y\+JdRMbV[&)4fYTTD
]dFE9Z6f3CWXO^M.R7NdeKAKZ_<X:<:3T/0PgI71dcbC+f]NS>C;?eeO/fHf<fEb
dTf;P=.<_#.fO.J\X+QQMN_>H\f8&dcX)CQS>)-)F<H<[=@Q#O)g+10+:6eP&GLP
9]Z+ZGUI3CL2LgA/-707S,8-VYMSUN9S7DZ,f#0_5P21K49;G(^O;:QbH&-U\6J,
LG=c+:g9C2JPRQ.E#YSP\_a[MI1]1,XA-b+&3e=4bC1Y[\/.83]KN)89JXE.a7OQ
Ld/aGB)USXdMKAgL_@^>8[4LcH?MU<-bU>Y3SU=@6]J^Q7GRO08S\_MgL.?dCCM#
/HR&2=8GHReZg;g_0eWAc5M?IU?X^[<W?<@YZS#H<^bQ;@FMDS[DN6[U.G&6Qc7b
g0X1@D]&87X)\Xa7&4/HV\g+(91a(MR0K#;J#U]4-Eg<7/_5JbccDI98dI23[:\-
YR_g&D&dN\JKQ=W1>,020-RL0MdB[P[AaI#:[B_5Y;MNGLbFJ_<ZH:)<D=8/I.=?
R_dM;-3SV\;f:L,.I+O<bZA/)FAIO=L0aL::6>B?V8>LG\Y(P>@/\U794P_cgYVS
>Y[OS)gfRe-B9NbOU.411,C6_]25a(b<>6\N]F0L,\Sg2K<6/1Z3&7ZU)BT69^HL
S03W<:c)YS^)RaEH+MaQ9A]V.8E7<_/a8FLPOPgBUe6?N7>U)Z+2\SA^BZK)g8&?
YTNbXRK87PA^D9A.YF(A4_c8V1Q27I9S)BAPa5)C=UP2SV?[]f=:/:\0a0,NO43C
10M(+B6#@>\T@)U\C9,9\UI7P?Q>0C9J(c>3=;b[F/MND\#>DO]4:J=Ya>I-QV.>
-DCL]aOVDMOBa]77d>G2A&4AH&U)]Qc,NE-/L[R:YP9AeAO)NTZd^\82,V]KS_?U
J_1VAFLF;8NBUbdf;3gFZ\29:e48c:9T=IbgA+=K&eX_e.TN&f6J1_,X(=NI(0NS
_:RHC)#T7<#8F?L512\:eVQ&42.d:J+2QU_S7UEN36Tb0<a7^RXe6O7+](RJ]:fI
J#A8O-P.(YbN#3R25F#2G[UZJWJ0]=NTXU;J78#dU[=?6WB&D\5;7CAgN_WfHd=H
>FI:3#c]_ZXHUU+GQVEe7@97O+/_0:E[(W;4b78Y-8;D:>VWO&3>VeIU5KWUC\#M
eWeH+UdQN36KJ.=IW^4B7c8;\[:eNBVV:C,DC6Vab6EBa4F<KRA4H]M<8B&MgbD&
9I3)E7J_49(1,W<>?[c8^@[R;QE>2\cXbG_B[EQQ>O;9/G=2J4+\4M^\ae6X8ZfH
)a)&=CLTIV#X(78Q:\53/K47\OZBcP#bDWL3@IUBGgTfZdD:M_HXgO;CTZV[>OaX
8@NIS7\a.(_FaJIAQ/>,SM@Tea3#@@^OB)U[gg(Z9V[@9;)5I+A]_[Q^T\Gb3HG_
SVMYPb;JcZf)-d(Hg]HgA5EKJeg1VX9V+=a[J4WaW0D-?V+f8.D^,TK9A;E\AWHU
2?+TWJ=_\[(IcO2R^5\6=>40,K-&VIYTKYV(GW_Y\5WdQ6DG1FD>^XW-65;1Vf;1
GU1/^/X.Q/eWGg[Q5=H5[WgW.F;VX^/9XXZ?/G\IVT)1aUB?YfL3)MA/P/>R>++-
,B:]XE0XWK.)dSNZO7_?/3cTdR=dKXD2gZ6C12I<HU^XdUeFDc>BRR<WYgB:=#O]
T:^dbK06XWH,gP#,[UHa]6Ub#78?BG?6S\1Q&HLU23(0Xcc03PY1OHG?X,3&AC/V
8<Ig@;+X8XcWU-0M);U?8J&e:+F@FbN,5dcffa/U^ZMI?2<bGf4+7:5C7=gXWENE
Y?0&7ID+WE>\fY^BG;#IRJFLd&E(9?4=CeB5BS5CU4#VO,I;.>P./dZ__,1D0;PU
R@;P\S4.@Z_.^IY+;dRO(gB.>Z)Z]HP?e&OI9fB45gWI2+E&D7P/4H1XKF5:_6:2
:3eER-6X:_?C-::CRa3AdJ[&>O6[08HHL[N(9P&cbD9LC=@YN>=2:)Q?/(<;8CY3
MP07\]Z0aER.VVTD@=_5;O.Db6F8R/YJ3O6NA#0#ZKIK+)g8LDa#]E&E-1^3FHbZ
f>^SDB0O\)X:)^@2IQCR3G8FA28+L[GS9dI_S[&8G52J7N8V>^66Dg6^KB41Te35
33e?aT#]=TO[RIDM72_OI;e,_XUDIIZ9-c,1OA,eJb:dX^Y5Tc3_2Oa^MEX@egM8
,Y6].XKDgOM^9)\Q7eg?==W.O)UF,g#,fY<PL+NV@EN4KM9FJXWK@J[SS]gIeP4-
ZHEW8=;e@f-U#O]7+@1K[b6c9GWT>^4K449dG>cU82K/Mf4NL>;a]2:]T)^IA/WX
/+@Z9K+X:;1aE9/L9+G(b-LYZ,KYHY8b7EEbF8b.H#THUT6a9R>Za(;3R.MM3,JC
fVR9SHCXVDdZ,)/NU6OeAB:I9K_S:#804P,KWRK7GaAGT>F@2QAa=H0UH9D44)JK
DLH]OU;_9=HO\7cO23)_28,JXc:9JDJZ(C6D8ZWZLE59QZ<?<2Ff(Ab6LY\e,A63
-#e;:>&E3F(NL<:&E-ESa\=&KW0XNW)(FCN]3M\KE>-_^O>:CTa^P8]ANgOE(8@3
D:e#O949bG6\/830^?\=I=C)(]Rb;8Z+>F?,7-+?g]d?-;S#>5gH7@X>0DFf>&6W
]0([^d#<[Bf[\cHeLA:JMc1(eEdYOf#:V;PCgT\YTHAXV=9S5cT/gD=5Y&-,-<UR
3D.4Xd\Z)M=AY_?+L.4@4<aU@#SWXQ2JK]JdgDSfJeD]&:VCQ-J<SX63D[3JXUN6
I?)^TBa81L#QbDO75<H,Af(W20Ra3Mb#Q5d._.g)DVQS=5DgKJJEN]UeCcC)19RY
bS;SH:Y26T^40S5/L^VK#-\H;U\5)\,^N#3_LK.0#^e;(9aW8:]gZ(BD#\6N=J=;
=cU^UPe1GMUWL43C2CO#DF_SMg3cX]U8>5:9?I4@?A=L&/(HOUJH.\gT.fF@fMAN
^ZBeI.#.<g]T@GW[Bbb/Q2IcX7fNHbc:OeWQ8a46G<BF@dT9,?;X=a&(1X/]RZ#S
<eHUbfXc3)X7:0OBM+>TK(K4-X:+D\YWUNOC>1[F[K#_(;;fZ_cB0B(WO5Af>K8[
.\?#UgBNP>8Y>,g-1@dF8I0S.,Uf_0^C)+3NX&LRc\UA_]A(KOC24O\&)N0;&#ID
P,Y)9D#-OU6KK=C\;:UafROC9IL>A>O4Qc?J]=BdF1EKdA@=36])adJa&A=>GNFB
XM/KC,YO:>[YDL4\WG8CQ?7Q^G=)b84K14DgNDQ087dYbJ4#<B]1Q7P]4X.c&JMb
GCNZV3QNec_C2,)8)X4]Vg#e]P>;>6_&K4(;;YSaJ<T9@01?^?KJM<]?P4]>7=EX
ETMeEH5&SN8[+<b@:5028P5[QAZC0b8#?XLXCXA;0:@63)-4(K+,d6XFJ8.Z+F@R
J&WE7TUGO\<AKSN0_05dNEV>MVegF9Q<,_WIQBVbC^SX&0b\D6WR7bJG7Q5Db6#P
QO??aUCgTQFS,#<QAFO_dAK]LWR@dA-P-,S@@V,5^0OXNe2XeXRUGZ=<gEYJ?bHK
a?A>gd_,\ZBJ?A>.6.]KNTd4Pg,TI;8b#2?LML8ER&SI>O+I-KX8RS,SVc=(e@_S
<gN?bX)8edYL2:,REU=;-\/EADVV38IC3R#OW+;I^HHa4HBgQcd(OgHOIQgU0WfH
/G.MZMggIU,-5gD#+Q@=>=S:VZAIAQ]2LG7EB6(e4)VK+HXB1OOA-PNe2XZ<MLe.
26CbY-AA(4a^BOfQ0+Lb86/BMg53bVH1GgJ([D^/0d/g^CO(=/R4gF2S@3JBb<][
@)JN1M_DUEKEI3_6\+IOB0gGG3_U^WK=^dD[;_VLg+Q65?/^MbYAeD)3ULdK(aVJ
gaf>N0Ya+##X?9V&I_]<(7a0X]?<7a(RQe12Y)>62;=B\_,:e_Xde)dGGb^d(UJ(
KXE-<YYB^AU:GT5=)(=gG/Od]7RXcgdP@OKL?7K4:3C=g&S_^PNAgf20>P/OZC0f
A6J8WZ_K-^>#_Q)@AfP9^-2Ic.K8Kg[b\MbG9GXQM\SR#9AJUc]/6+/GR^0a:8fZ
)2PXNC(/77.]X^1UE2M+&=LM@V87HPH&C#I^PHWPX=:Jf=N0KBE52X;+\8.]U/P_
-CP2gIIf4F8[:,QZ622,3(X>-W5<8_(T&a[>OB_P8eRb>BQD89gb6JELQ7)d=XRT
/G&c]_<B7U3gHJ8-70\LIT;O7MEdf(U_ZWe&PJ]VXI)XS_9eV22McUDA/R[:F?#^
,YZ1>3XK,?U;-G,4J(3@Y(K+_,H@.<_[M0+O29^.JPRV-9[c\NFTKRSQZ@#VLXe=
>,3,^WRU&L&E3BNF\MZ<3]e#M[RY&G^N@LEU@9MF1XEb8[fCU])Ad=C)ZgJPK1O8
FM2gQ[,c,gM/(183.[W)0#;aXPeR)9A)[+,WC\ENY1W]^e.=J:b-^=Rcb[8G0<cV
\]@5F<:M?@6E8>8Y:JHSV]1]676\]cL]O[H:EL,HNOdW0>fRaL@.BR\[(JH>:Z/E
--eIJA\D\8;3D1)CI=IJ+6#GG.=Q7<+>LR:9HbREN0VOH+AX@(CD_;O7-fEKHaRB
aZ/fQ_Wf0If>#f=P32=5bH0TbDO.c\HVf;(O#UbFASP:/.gX(G<:1_]];+3FE/cc
^4D/Lg&RHaGYeS7#2CUA.SI3;=SAc@C,9R0,.bU);:(#(X(^VXUJS&<E)3E86>dS
;=7Mc2H=7++ce/Z;]9Xg&QYUR51Q&.UA+=<LK[6gKHDfDYX=6A[aO(HZW@WWgCT1
)-K2-4G40T8#N;,TP(>M?6OQT0_-3&7_1AG?b9ODWMg15>W>ZBN^799KTSCS&c9-
;GL4+3N<[XB&DL88HZE@f@T:\ee[B_BZ&feL59>5B1(O+]7?LO-@Hd/O3].LKc#3
8QePd[B.AHbZ5P(M&UBL1B,Nb.#SE#O)O7(H]@b]/d@[W[_=PKAbd8@T]SJ(P(/R
g@FQdH36\6;f]>^9@)(L_,VIE?K\KBGQdKNFI0JZ&MTc5.X#KJG4R2<J3L4_\5KE
G4DMCJ]Q5a7SZ97;NTU7;V#4AEA?IW<+CIb6<Ub&+J)>;Fe:Z#PWNM_C^30fJ(Zc
a^QVcdb5:A^J1M>U\@)BZN]LE8Y]R8a#LP_5OT5BbMeG#8e907>@><9/PSA;K#_3
UDR5dP\)7</4D:PaAW#]S3)AB:WVGEXSZ6XS^e?B2XRP6HDgD[C.E-a1M095VS&<
dS?^-,d?XX^2MO;gaH[0TFHB;&@a.MC1,2K.b/0GF.MAD+5^bEBK[:ZAEe-SO?,O
=c;fb7F=<L8\-C(M>;[0?Q77WO0_+9.W.b2._[(V3dW(?\1eU.T-,X\G[B_LGU:)
6.b&6cbE>DXgZ\1WGD&)UW?NA=:Q;S/H2f7AH,S.)P@_N].WSYTPae.PD\/dOgFV
+<+FZ=:>5Nf6#X@0S\TBX?ObXa/8BG@8/&#PaML>-@BIa?a/;+#[TeZ73H:]d)[K
>M[.)C:;?B\>A0K3)^&:+c31@#fX6V#KV)e:Yf6&?X/:J9-C2(A2Vd9\X)K0;08D
8\BPG]FIXKL-:@_YE]622]E0X);G4QH>3O@C+#KFeg\52CDB@+Ad5eGQ3Ge.W6&]
NVe>I>.O@R7#[[4P3eTJ^Z1cbYZfA(Sc<)[6J(N?(Z;c(W^T\<N[43&@4Z7ZQ1KC
2/,TRVI>T<e@+R#7G0^,;SXf]Mf:\(RaX;9HI\&POdB7956=EA8[V5dEWQ5eTDBT
BPZ)d6^3U5eWQ7d6?.1T^AA&,X(F@FQYcKQRH4(Gd2YWc\?K/aFLM20A3]g8)D7L
&g3::]f/U.S)WY08<;fSR>60BaAgC/2B,?#_9b5SL:K:Y74WVg;<24,)@YBfIS7K
FPNb:d[MA#K6YaQ,I?<8<>C1=0-CgC<L\6c5&UMY&IP&>B]/FI]Y?eHdU-]g-aT(
g(gRFQATQQQB<J,g394MbX6H(DTa3DNY=)&Qb_6aLDI4L+F7GDT+GOaE1CAZ&R;.
0UbD8-<;AIHOM,MSW+_/W\_S#)-2[g=JfWW6O]F&4WMK92:_4-7;\)JbYPH\W0cO
(>)b?_N+E.:B670@XfFa[\(,Y^V4,BRC;(^?)0(>ILR3Qa;TUHD.XX2=UH>3[UQ)
bSP_IOU7Z-?Vd<9-.K[&2(F@Ee7@GY7S4UD8SU^E+&R#KX^VMJBP4H&fXZTae&Y9
P,95J\:,1eAFS9-\TT<+]I^Xc=8H-:YWVQRE]-MTAMDSJHJ+.]A8<XCc2J\.X2a3
R];433O<O<-ARN1SaC>3@/^5B83.1,GIX-UXKWQ;.gB@4fVC<\^KNbL0<aSePbID
H9[Ta+4_#[+^+#TR.fbN:^ZHa;PYEX=09(O89J)O<YT8E[PK[/-9=+<5bG/?(K6+
<c^U@(B-g&fIZ&DXaH+5/N>,dg->\CXMa@VV56fgF<3Z(7F3AE3C#GR#VRO6Lg+C
?1KS.+D/E;e^9ZC0dH327V37\.\8,G2eF.0LH\K9#P79=GS87.JQ12Z_T16:d80/
V\#P6]7LXQ/<4PPc-D)^J;?)P(H/MKLT6+e/Ba,,U,.;0X3U(<.C6F3F>4Q-Td+A
_Y6RaO-9Z0ZcBR+gfB9A=a9LQ:[Y9,5Ya#@UO7P;_13Hde&P5AL_U30E,TW5c8\Y
&@M?^La(B6A^</8++A/ZQ\W#Nf&?,(9=3<(I(R\9.>.+cB\g3bWJ&c6&+fZ/UT#Q
AZ3U=F&YOfd0,?:3XJ2_35)R_PC0O9=>c.:H\@^JOT@Yec#&1Lfc3T#>F.b61X4G
0^]ONP<D)gFPT);Y9UDVF<)dKM;QWGa#I5O_[3S^H)A/WL8B0A0c.<51,]2^3578
Pa&.DdCJc+ZSVgAZ^DD1R]DM+#M=I=JZ)[K>DZcK).0YX3<gM^PAdI9+BE^W3f.0
]#P40@1dSe7VM]8g)/JI4[F]]#N&9-F>P,c@)4#4EcKW?6]g.6-<8VQf150S]^gU
/&DT#S&&.LJ^&fFBMc7(_RK<+f)UdJA&D>e9c?feW4S2:BDLb?R^eNf=/4)TYRAf
D5_SIHcD@EDcc6<ELVcEF5e/SKBc4;[1#^<4(SdKRAe)3(E:-KUI,N@_&bfMY+Xc
<#B..\0ERBWdJ/V(FVV^(S=)L&[V,L7Bga0a/^97(3,F>1U)c^DS.geN:=c=fe2]
OeTL>?FG<g:=&)]IL2M/6+6()1W_Lf6CN8Y8TPVC+eaT[c.HRI<PM3b5UL?]X.+B
[ITe+H=ZgGS5R_fBUBY.YQUNF=8ca_:RAWU<QR0NRC[#^JCPb:.LILWYPCWT<=^7
E?d;MXfCFg6&IN(Q;AQN;IR0&c1@#GQN(_gE&baW7;(g2(EQPYN)X0fL_B++5)&g
#]SLfKgN-L(3WSZ#eI/#Fc(f\cZ))b_CEGJQR>^.C-T^WNP#-G3f3MP9dZF9.2O,
A(JbId;>?gDX;:B#@@(LXJ,Vf77=fJ1VWW>OC6BT&5dD<b7/B36f@#[7c<MB[6Z1
^@[=]NJZRJ=,;c?M2WJ&MD.;OXDJQM/Y7XI3,QO@;/0))FFZb+)L(0FDMI1-J0df
&)EXEW^4a1gC)#Q=@O9ML@D6UU[1T^E^D1E8V]D<^,06S<cO_RA)4ZSG?OL6edR@
(,RO4Ae^H3Pg@ed,8:6.YdLfb(cO.STFF>U^7R8ALNX>=INaU_AOYL.:NVAQaD?<
9E&4,ZIe()@R:a[[,_,Ee.(T>>GbCB_XQ[[\S[VVd;/\1];@a4=-7:GO2<d9Ob(9
Tfc_g?7<gIFb,B;X,2\LI6,+A+X3dWeQ2OKWZ[Sb:YUW4P<;3./d)I^>a22@\50)
)>I.Z<CV5,>#V]a1NPQ;ZfYg_^PS7W]cWFc4MZeQE>I(Vf3N4)V4]NH[&_<ZW3I/
&NAHTKIIe.I>CgRU_MI)@VO+-..A:b:BZK?6VU6J/A(WJ:5,D6LR/MEZTeK,JVeU
f(.?Q^PfI9G=AR/JRgd8MeR>:3+<+DL?#@a4U+C5IgJX)]=;e1)=+b?\CO5=_VH&
#OXE_G>G+?MWg6DU0[b,:^@P8W=++2)/Q[c0N.fQ&1Y-]4QQacf+XQe_[#:5AUC7
MA#,LEIf8#/>F><S&>T@,L^R7dS92.5V.Z=:K,#VEbWSZI75,+>A-^cSBKVV&Oa<
.f_FHNgWIKUfU?_P,GSc3_gX2V:JYSUZ^])\G/G\VV?N;c#f4TIR9IN0.ZMG6<d^
1O&+V+-4EVaaW^,eF<GAaD+K:e=7,g2DfHX:+FR]UTJdGINS,.]GX.QdbK@L4:7b
B9Y,[&HE-Q[/Y8=F7&fIaeAO3+Z,KY9K0)IT&K<2A>D:?3-cZQV^^8U\aD:,36NK
WYAUQSV(YHYJ66VbQEK(cW;6dYK<C1^C8K2)G>>8->_\V5V/bG,WCOGK8dG_U,&S
F/EbT)+PGa9eDE&]?J^2?_Z3_#f@GQ6@b\/#FbOK=GD-+OP)(.1:+W?=^U6LCabE
OH)AFOM4>D;ALFDbB?AZd:,24(0[Z]HNg+[LPR#?bg_ETD_e>#,RXP^@Zd#Z;g>a
f]<;MR5cKcKbA74EJK2egZJ^aG/LRPAg2>KL0[PIgcWYRdFaMO\38__PKZ:aa?D+
N(N@(=\ePWVRVM<35S6#bAK6AYHWD88eKRB5TD3PD<-7T<7=_)XWeBM+47S;\O:7
6H(eZ2Y=Z-#_aF,f58K^J2_GOTaZ5_e&?MBZBDF56,QH6AE;JgCbKKEFaU]/&N[Y
^=G63/3IM0A<M5#SNUP:S7_<LV&25K++]MS>L52;N&_cY.QTJA&;YcR_ICRaV2-:
^S+URIJ6A0U))EHIUH847<>D+8WWcRLJa_R0(D+US]64WBCaC^U_W_8)1,C=,.1>
fP]P\T7Ae]B;M.];f5dB5B-U=MQWPDBe/#+H3KZ(@Y#/.QS6R2CIJgNROX.@G4de
UCe9OE5#QXP+cQ+C>4=V)C_gSSM(7YMGZ5L?Eg4)7Y-;<1L47HCMVbZOPOa94N?#
\9b;>4+.6@WV;0\;A-T=:(eS>[3K1Y6aM^=-E.aIOO2@:S,?;V8O0ELNdFT:J-TN
(&<IVdPU.-3,d9V)VOGbN>YP/cH-;842Zf#<]0+2gg:>N^BJW&c@5X(FcK@J.6]+
:BA4ADa31OS?6eOR.V(52KMc=a@SCK[XD>I9[PKSYcC;_^WFc-,/>)[CT)I<5<8E
;dd6:<HgeaE9B:2]+K6J)UQAe9fPULUY0KKD0Y.&9_E+D<QC1[/>K9,Y2YK<M/];
9d;#e@CJ]-Xad/N_M,^>MZGCUH75-f?;D+[M]20Ie397<FB\:+:O1R415@_<80Oe
K?DQ)-DBc6aZ2#/;3?<L/7W8&7CWI@_?[OFb#9V/-5(c9P665?_2Y4CPWI36?BN5
A&Q&M#,Zb._Q[U/<->4EB7#PfP33:gZ^O@cV&QY(D:S_/13f2>A2+SOQS_8)##cD
N;Wd+D^[5>@CO)4F?HD^5W)f\SL?T<HVe\Vb7?IgM]60a]2ec\5=;.31R2./Z-A-
bP#Afcdd4bIX,Y<JBa&9@6?PM8C9.b0(N?C^Y,b8cW1)0FW7gU4G)#;13.EU;C@L
X^?N1F=fP,_f=<()<Q34X3DMF_3+8)BA2Ia>gJ<JA)]OdUXJ(PARDfO&B50M8]BZ
Nf=T.21Hc<QbX]CeGKd.Z7UY39N6R-C4]2X3R;U+8/+)5:=88KY>@eYL9;@:F_1U
Y#_1Z=d;5eWJe&gJF^3;5]0;:XFOP03gJ1gW3-a9)#SeTQb[@YPJ,f-9:YM#RX/a
g0\&gabHR\IO#Q#<d&R3(]c;7&6=>dTW&0eDG)dHgd^Af]//eS5gY.:FXJ6=()TP
Z\.^E+JAg+W1@:\#?L@EU#L^6CPfRY#QD5XY0K10e1E#X9_1EVM:X>/3D&/QN(S/
_.XVYPA9QSRc-Xd-J0(<-AOD7Y-cS-8cNaaa>7(gTeD5BVc.6QIVMUZ\/)6.cC+<
@(9b0T::)#20a\2Y60YX:XKQW4.\B[V&:CDQI9B+]KGJ7FdO>&X[?;E(2IcB5C3_
=8P&\,?>GWf9LV3SLeR30(32+PE_@^]SAdQYM@+e<>YD6;O8W6@_D)#&<T4Y+(X\
UO=Vg(E\9NLL@OX\;DZRaaPTLGAS]AMA;A5fGN/29FF+7\0V&]7Jf;cR-FUC#c8a
DT^_Y^e)fLf:@Y,BO1W9222dEIL?AXcWNc#[#]JNdgIC#X+VC(fMZb6GB6>2]_M\
R>T:8Nd>OXT)Kb-a/+/YTVOY,]:>H].&JNf4:(.3FR<--U=.9M@<6<cE,TW:;ME3
].<Tf=))W]1GcRPA25E)9]BVYG,NCa-XP5,=-_Qa>KB9<WA6B>/_K&_ZS;@Jd7,5
U]DT)bI^-MR1O0c8c<T>E/NbTbA]@e8\RI]00W<&-M)1#QB=31WGaALMM@5F&Pf3
\^KefRJYdg^5=C55_+/_/bF1b2Z2(/TE66S@+2)CLQ\-H7HYJN#9UZ9/Fe,A8]MB
^d;RLU(g?PZDMS.1\15fE71G]NRF1).A&Sd,:L@;2b.884I0B\<bUX;__CY,ed#/
b5F=)=/0>XJe0PK&FSQNL.O-S<?G]]+D>?-SF;@@A3@N_?LL@--_NXR35WQ/.VUX
M00#1LbN1BcNO3EaQ&IML@.D0dT:6WQ^fQ1g&Nb&Y)HWZPeBE^eUeTN_a+;9a3\1
;+(J)FMM3F.@7J6RQ]cZ8\SL6^24:O(,E:XfZE@E>\N,[N?Z:<NcS::#(N4Gcg<K
P)-??f;9ZNG)EK_Gd_3\D9NID(/WSPWQX,O85N_\7N1^QfOZ#gW79FWOUOP#1(Ie
4]c7?Jd=7g8E1;],eAN4^_R8#92Rg,BD^[7F(CW;gPPKC#&c&OU?A6\_HF,fcVbO
^CNLE7J5O9MQD(/NSYB6Udb;f-02F/MP(]_BH)RXQ?M5:]3E#76a#T[;RG2S]GHA
E=[,I@/bMK/3GC4J)8-T5)[[8(>:]/<A;9/LE2]-I>fLAb>#,YF0LMUSYH99:(V0
U0c,bXGHHQ-QFRF9-Y3#\I3VQM>3E/7UBg#:DRU<R-0HUJMeX26);Bed60YSDeKS
W#a1(,Q,M3BKcW1RVQ+\.@+U05JHR+6#^=6GU(/[LJ3S_J;>C/A1N1<C_6HH3gM)
/#f@^S7=W:8THRX:T8629Fc26B^?-gYRQU<NSA,&KS#)bf3gabHXATCL3/6D@3=G
g5bU4]4XVIHF^G_4RF9Y;0>fQ<NB^C36c9[]SA7I;S7,F5L3NY0;M(YB2I3=XJY[
#N1,ScJ_DW@W@07L.-D(H/+&ddC@N[Ue99J8bIZI.:d48aE#aA#G@+T8Ic>]b\W,
U/#:Te]O]9?Z<MU9G^I+c8\9/)5CMNJ^e^QQf80].ZeV^46T]XS26HfAT+8#T798
gD8,3_L,&W<>(#>A:;CYbbd_?X[6c:+>BN0Z>]#,;L?&14X;)#3-KK,IA+L>a,:@
Z2W(Y(;1bdK-gP:P?XcW0JR5_I,F6G?VAXUS)bgd?7A7Z[67Gc.@N<65;1^(dSRD
W;W5-&/Q8gFX3aXCSO6fL>:9])\R1NeY?U-2&,G4ede4JB0c,N8UW:#bNGOe[+5>
ITB,f4a46UVL<(07_Fd[fJTgU[I6&X/V0BV,2)Uc[+N]bIUDX#N9Y)#S1\)dKB@I
T-fEOV,fDBe76_TAD/1P+6--?=OH35FGC@P[Z&E)R50&cKM(dNM.RR1^E@Yb4>1A
+O;g-de4T]PYJG7)TZNfDad_ZS2gZ6O)7>+Kd:<Rg7F^V[+>/5XZQfSARgRF#A[/
O.OSdf.362fN:YG=_g(NS21U@W[R,eA8aZ7@3L,2I&@G#1JE7-7DA-]]@We7,(P0
#T<>RB\E8JNKaQ7_C,;:L@fcP(O:P__MHYe,T<gI\EZf6>.8/g9eMPPB3\YR]b&P
YV(Yf.ed8g3RNEfbBMGNd:aNOYQg)W33_ZQKeBFdeE6UKf6b,C5(]Z]:#EI>c_@M
dX&4M;_=SOBO2<R\EV3(I);/]Tc]KY_c/?7;N8\E1GJ@Jb3[#Dc<+L[40X,-b6M#
487H3cc?1P;&aNJe1e<UB8=BC1/@IcP2943>X;/:LDbg?O(DJD6?cS\E9@(ND8?T
a;_^K8ZQU8_cWc2dIF]^)(O_:KF(95EMFSJ2Y7G#=0Jb0?SEL?#,#:U.9[2<9_U/
@XS/;X6Yc0HAHN0YL2C(B55?)4Fc5XAY81=@A4=EFHB/]=E[Ff6b1)-gF#(0/.?9
Z#b\FK^<]beC/NOFH4LgbG]WO9K]F&K?+QeKI65W;&P2?[2^KJ\1\\K3HTRP-AdZ
B)C2Z-UJPD19,J_H0FBKDP_Za^fS+8(AGFY\Y8SWg6++7H5T2.Y_NX[;a=,NPg#9
HfeC.R@.4-;#(&SY30+/1C,J86.I3503E(#\2-P[\A)CP=ES+(gRJ324-fI).\Y/
SQdQU]VOHIJ=cC[dDHSQ,VX/Wb+<bI>c1(P&/A).H@T+bU+3CXZ@HIL2&BS1<)[d
-XHQe9=]>3I:ZDeTW2QSW4.?SXNGFRUNS4d76+RS[S/c/EV57BJ;MgM0/N^.WSec
+8W,:I>U3-,(B>R=2TET63UZU)KWfHN2XCSK+9HC?#5,:G)Yg6cJ?U?LY7-[eF]@
fW2I^#]E=34O.gSX+&I\R&3g?USVcF/6QKg;S0PHSa,01RKZD9?09=>F9>T3cUI[
g_BYJf2JaJT+dRLS3..([KI(6,g3W@V#]I=O?BaM_F/\HJSO7JYVOBL[.BST[af.
X8-KJc;([1+RW0ZI:#L-(;1@R4P81TL,<B=OK[E>:>E]f\\+<+_F9ON-ebbR4-=D
HANGe02ED3]Q(dJdZ#;14[_,>J,PQ3-Jb,W@H6gaY>G=GP.:/[?7-2eEf2Cb,cKP
E-G5XOb[d29(eW>D8:ZA0fV:fga6@O\T\5Sc@e3W3\]J\.)EDPJV1W&M[eYN4dM_
9b<IPERJS?UaX0Mcg;<?W8T:DcaJ(^^?E.3^-0VQB(];>b:ED8GDK+B>S3af\Kfc
#>@PSLWH9>00//33U&(I8@3cWA9;Gd.=A0YQ-].W@Zd9Z6][Q=>++a0^TSO-3@WU
^Xd:Kb]eF:I(Z=/6=>]&B[@0a5Y.T[H1.[6TQa3Y&\1S=SXb/g,&X:PQ,fXO4F+X
bEdDC+HKY@f3=H9eUbS^2J3L(+a3XRNMg&PcB)&b@Pe(5@@C]B496Z=(I6I5/gfP
AHB?AV@]GVQ):K9Cb/.5(T^+&b9LA#+ZIL:Q=@JZB_M?b2MK4@(\1U5VA?&>N-U2
eSI=SDa;3+:5.YD2TQMPAJ18W.<IK\GAAN>RPT8]#T_:JVK.YB)eOgWX6SL:QH_A
,:IP-J)LYZQNTWS3gWRdHVbJR0=UKG(U;\YO]5;M\7\\J//W=d[8&C0;0YD6;EO\
N.H=4:=4Ag\=NWI7\P7<??UT5-R8S?fRQ[cXLTE,^bd1L/]]JOgeJ=UD@8B9C3/H
VA<OTTa[.cM6@/8.,16eAVXH_H,UX+A4J&HH=BVBd5L6OdYf1^71Tg,KZT.,GS.C
?+,NJgbOG6e7T>c_CYOSUAWCIL<@9a>4FPgfe,;&.XKPB.H5USPb]U.<B1@S#eeQ
C9G-U_^/.@5A720b(,S>WJ3IK7>AYdcUG_2W.Q\=^N33#0)[6E\R=#1E6S>ZLdC3
Ve>F/P][+ZGG@;G&4L^R#9#&QZ\G<;-NF5UGEXG.=L]MfFKNbd,B[8b7Ka#XeQ5M
aJ8:fQR-;gF4-U3_:W.//,5df#E0GE=30?d[-.XXH+GMCUL8#<B@]^CbRF;.cZV1
Z2BJV[IfO\;&YEMgG=b_^,b^,3>056[EUH_=7]ffb^]&U4U@/gPT2Q_85H9Ug(UD
d?)aSVZS+95?6PVSP&]QEW,.Xb8Kc:gaHURPDYX2Z-[?dQ;(<fV.K+#N_#>d)3YZ
A):+3eF@[\fS[J1c]PSVUF44c-cYc,(6##YEE>DE)\?A9K^XJc?>/E]VF8[\NQ+D
&IA&/&fC-2:+31cU\PfaPM](S&OdGQCe-UR^.=F((EUeN31;U&Lf:[>5,^]0W-:e
^D;ZDYcM27d7.XZdX@I0/ML4aEINNGXLKF3J1)VFHLJ-PRR01PQV0<(eaY<?^IH5
W04g]QV?Wd\J5gA(5N1M2?-\C]bI<+D+A(NXQP:,6+(e#Y4ZDON>cPFD\K.a&H:C
UN7[HgNP7<VV<cC,XC?ON>EGaY22,dX;(@M=[]I]-SKDL[G?FLG32[Z=FHHWB#N&
MHccG^[b#K>_490;_bg+U9U+LD</Od\RJ]<Ge/:B>^.[_D::b3fZY9O1;@,LKF@-
F_aL.\=D,8XeTZ_ML<=]Z3V.d_H0:LT7BB:2&4(T>e#/N\)X4_Id6IB3e@L6bXTO
-fXLPF3f2cbT8DDL)Z7=/)Y@a.DE?FA.#&fR8BAcVO)4E\-/\#U?N-3HUgG](XU+
ZO09PSVC+ZffgMR[O#[Ce1I/:1ZM,&;[+b-HQTT9fCG7:,1-Zf(Q3^.148Re8Q#1
V#<:88<+A?I-5G7<VPE7+BRB/NZ&V,)G4F5B;8K4HCdNdMBG9U:1-,R7?0J#\Y6?
cEG#C)PK.-2]#)^g;)&HBcJ@TgC@BR@J???L4+=+^[8KVcfTc/d0K6/IQY;DB_D2
4DUAQ6B;KBXNF3,UNU?\#);+)NQCN0dV:\97R=^dXbc\.B4C9ZVd7AKNOe>F@/23
]7H4d:CP1,cg]ZU\fOc^B60]Vd5D9:LW@NMPaW=30=A5MIf[@_1^LU/,&GW,+,T\
F7Mf]IMF;MC@[JMFYB07&I12g4B^.1Q,[Mde\)Uc7ITVNO-K]&6UMR=[98CTLD<>
Y&EF#>C#4=MDNdI+U_We8@QaA&W?=.T2@&]+H-L1PZeda4TUUg[7,F?cN^;-E?Sb
,c>W+P,__fZ,gMB:&PG\[2d\3CW1f(;JC^S&?Wf)RcbFIU.<HQ8YfYHA5HGGQI/1
YDSND.I&<VJTRBOf5T3Ve.9Y#ED97(=eGFQ6.EcR>1NB><E/4DVIf-gC,UQ(6#]d
85cg?d[Y_bc8OI\Dd_[IM^B5/P\PYD5Ag9,;3>BEd&ERX1;_202e1H1fVRKI\W)R
1?\LUZH/DTM[[,+&&<;AV1HbF\3]]H_OL,V4Q&MbJ4dPF,G8a_6gDAfGYU-ZLg#D
8T>-G]VZO;8?ZF7XQW)7Y.L+aNRXP2BWWcdJ:1L[F?CI/K3FX6(W8H4M#G7T0LB^
0[+5:ceN>3UYY(Wf,-CYdEPE5>6,O:bgb3#D_.<f=S4K^X.EYEWJ7_X>EP,KPCdW
=9)K5ZAae>a;^fH(FBB0ZKP3VKX>D2eg[(^N2I10a_\:0QTAWb?G=.B9,Lc9Cd#.
9UDF]Va(4eRET;bQQ[G_XffR4+bJ8PW\5_W-=KICOd+4=BIVJa#1EA1#)H\SUA_?
fUU\JdZ<GJ/Wg8J(CK@IBVR314d2c#CBdPe[<RW\/0J@=#A8/b#AJU)LIT>S&_N:
CHJF3:ce-J)NW+80HbAVRd,LIg[3M_RQOSHJV+_d)&F32_T.B-OeW-9KeTT])HK+
=We:.9B-0Z+:AKV9(\RSC[f4>>277P\gOU@5)cZ-Z;QbV_2.Y:?aU\6S0]U(XY9N
F3I-V<21CUR39=9A+#JK#40a1+@dFRJD#8d?Z2:7a:TS\0D&6?7E[-D9FTD(-e]Y
GFLBTYWaO87[&CO62cRBYbGPS(3OSa4G:&.?eIV_8H7E#D_Z5aHFMF&:BcgM;0T=
+,?Y_V@=9MOSQQD+J=1D5##0M8RBK[EZ2++J14RLga),3)=XX<S+_XSDM0JS?+Gb
W_C:6:E\4>8d9)MUL)X7V-f3PL+S=OMgdV=BTHXH9#<V/L?//P<\#2K@#+C+MOUc
GW[)UXLb56H]Y:[7JS/XYOY4VfLeQT+I6+TWCUHH[\AaS4Se@>#Zf8aEf;C(\\1&
F@F,9O.)C8Z#EPEYF9HL^bHHbSMC/#BdN4APZT_=,:IPG\d+=FT6Q&@EL7[)&2bd
KC<VE:\3-L[A-FgHSN<@IS_<ILdPTO/@eJIG]AR2MH9]F?eJ=dDc;\4]OW3(#46B
,5FUTf/7[RQH[0NQ[abJ#;2JZe2Y7aV3)1S:MUg72=QNfBF[Sb6C?FVTJ.<<6,:0
E+-5D8Z2D_9\TgBe0H8(8a5/-dde4.-,/4S_7e;Q^1WOWK\;^5\0GO?^6P#X#=E8
4JNMge5\L1&VPTK^Gf+X,ea9T&fNZQ(bX/eLZ]EM;a;IQ8]S^U81d2H=/&d8SgI[
b8H@W\QXT&V9:()0?OF,1CDdOOJ(9WO51b_\&UHQP[I:,R=1BYX7;60O:g:8dZL#
]+Z>W.I55(15E^fCM6@.16Zf+W:A#J:WK,<&cC=[Yg=<ZC0LR;IMR3&V5cG2MG9G
8+b&4a(J,g,7=I]c;:L.QL)2,:]B-fG/L;Zd,Z@-VAI-\S@F]:7UDgf3AD7UcBXb
SV5M3;bL>]4f-fPa<X\^9W-UB?E/_99+2]3WEU/QU+H:Qb<JBZ&BG>@:VdaUK;f:
KW_4aQ.VKIE_A6.<:7JXKXfc>ETG<f68Zfc[4=H=LgD8L-dLNBd4.:JR[\Ge=UaF
7-^=F<OdG+JA>-E?O0XZ+UG57OE-G3)&-HNQa.<4?E8dZO=?WH4Q9;P0&KX>#Lef
G=21&XL/9d+@M;O[RB01fG-daGG>Z5<U8)CA-d<cZA(=H2#_6b@=<VR53K>:&D/M
OBV<U@&f;VR#bH(5EMgN6a>GeXebYfJ7H/?(5P/LL@:8<1GZR:]+b+JQ;M6/T40&
7PcL#LS@e<cE=fXbY@@eP@6BIfdC):AQ/aFg]6aI&.d0K45X,CYKe.A^FLMS436A
a(^#\M];V(VXa].MG,bVC80.cS=H0#BKB&>^J^Pfc4)@BYK;.D,NW^C0+75QV^ZR
2-_F/LOTPc>CYWK(O8XIN,Ve^HA;HcLR,g0<Y5U#G^b9B7ITQ7gdX.MT\<+<TM0Q
,(,/@S#?Q)K53@&e^111_155;SC??^4MRTc_(&Ud[6<RTY&CaK5(BWUfQ_8S#^F&
AgbTe^U2<2?GgX.7@YfEFV0V66cBVUX3ZO3B:AV<b&62EdT.5c(eV(eP?>W=N9EJ
VEVf=9+KLTV2U.HcB#egJ<M_4@D^1TfOD^MR2L^&8,L;>KBbGcD^f3U36gWV\YD=
84TaHGZ.R,.5?46I)SbN4a<]^6LL1_9DO_7D8/:X<g(?d_fMKKbX.><SB[V,>6HL
fgYVKY#>Y,FTWD9H<+1WJ<K+.&Z[BBF\53Ta5bS:E.c85[-81_L9<,Kf0N6e?^>L
a)RNZ\;)=T>D_VDCHC,HZ.f53BDWF9e#1V?;4&TU/_4X>c;G70K,3U<dYG-EB6F=
<PO+:g6ANCC2ZLY6/gG85]_Pg-Z^.4L.313Oe1V;O7=Xd9&-NWcO5V(eg0(\d]J#
c6[;.?@OIWRfJE1fP_WfDZd7W_GYK[-&V5fO+;XB6@E0\T4ZNZB-e0AD7T8)JQ.3
^Jb7,B[]RU\3;V.1PF3MVN\IB-)>;WII]U#PIFOa+dSYAcQF4Tc-H8DfcXbC[33f
I@,^N97^eCHH,;CB]PO07(cYM(&^c7Z5F9X<HaZ3IIS/B,U7XQAERd#aT+W;^,gU
QB_,QI0Ac7:13&dG36W/PcV)@SX&a=,9DgK.33[f^bM?W;[:f?Z/D@T_MFHbKMAK
^:N@ECRB=K-dEITGVS6EXgc-2Z4dW;Zc1JU3&[/(\SRSJ>9d&FW#@@)IMKF,/]+X
N@-LN^1PKH;[FBZ33U;(X&0>C#&VfO0RLJXgbPLXL57BW,]?e5_2VB^ZQ]K]C0SN
V(aGe^56LVfgP#4IeLK[fJHQOH]c2:NNbABXIAeQLg-6[J::+D_dRBNf9)e#>Q=d
&M)-T52^E9;FNAAbEYbB=?UDUL?>BX>JH9U]<<UXS_3,#KFVX^]V@ONd(=2,,&JX
S^8eK-5L[;ISNb\PA#\(MOeGJ<E\G<)F/P]8[T\(Ef0Q=20/1K]9+;-7TSO?5Od^
DSad=+_^0.<MfB&bPHBDOV-,,#)BQST&UPC]TFF49Q0VRe_>5cM9bb2Y6T/3)?M>
&e1NC@)JDW&EY.(>Z@BJ:+3:^8JXA1=\?Zd#?@^D=.aR(?X>:LQGP6T(]F23QggS
c^0/?()GgdEMe(2cR8[VgV^&-J\3)c>a_+&-JQ@L-59S1EO#g>:(<Rf]1S-H3M##
9fA/D768H;W16]>FHWJY5WIT^)TGIg1,&TbQ-&(a_&_^FW^\18VSAg5YI2aBA=8U
>KAOSK=[53K5^NXC#2:f;M1(:]RKFeNX.fe(E&)R[.8>(SQPEE&=:c3KA8Z/;1C0
9(#=feR4WP4,cGc-S4/TPDSXN<J8T++F?Q_O-TD?f(5CAL3M#Se#7aS\cX6/&1@e
LR?E-C1ISSKE#V\Q<K0ZQHfLa=2Ubfc##\O@8<+db3N0b5Wc>Q7=6<53S0]]/VaQ
GQ0TWdW-HN>WAC\B&,L\<I49CESXIR@S#0>W:CBI746C73=IeU2D<]V9//KB=B:1
/RV)/>SgeRbTD=<aIc)/IcDE1@>c5.&a:C6L)_d(ZG-L/X\^Z[P?W._YO3/@AbD>
QM-f4@OgeG/WSI^HH8W8YbBD4/<V@=c4R_Id\\MSdb(WJQ6BNfN545[/J]<]8?Ud
BZ=_QeN;0Xf1ZT[59;D-g:R4+=/7GSNM9(#W/O<0VaA0CIQV+4:..FP251V;J@Oa
/PY9#<C7,KHMVc3MdKJ(7K<[AQT\4?Fb+^?)N-1ZQZ(J1fYEH#BNQ14W1A<-^,12
2_a2Q.M1;Y5:E3_9>YAXD#PPSB[a?\E6WVb+<7g7M@9aGK5]0LEdQTB-@CaS/c&&
CBZcd@@ef<6#P6Q8,PfF4([SA[]VYBMSdeN=@,g612VUg?[U7C34VR)[936[ZfG[
fRROg]VR\WGg+fH#V;dV#^S1@2FV-PJX/5cBP-.fY.3KSBC0a-T1;d[,@dZc&3MR
<Y;?JMTU3KYdNC,b@FU(Ud:IVI]\4XVDEWR09e<O_0O],]MI/N4]+VAdQ/FRCdXM
f7dNO=.@K9DTEI:Xb:X]].4__-4@fY3e4<1CagO.8?]3c#GN,>MQ.d-TcY9Q9]N7
36TKO1MI5ZOc15I59F11EHIa3#728I4cGWBM9C94S4,dd[&JB)McM8/&9NeEP7ED
_YUeXI,gMgZ[?#DA?_+KCXY_.G-_cf-D&\eg#\=(=QA#(=>_d#Se(Z_HQ?50^VPW
55aKS.)a0Yc)3H>DB@_(@/+6&QgGE8ef@bA(K?PN_5(aX/dFSRTe]42_\UGH;JC5
ab8@W<G<U1e#_8.6B=P-8IC@?2J4TeS^I.6d/C6^&F,.B9e8g88@3V;N3OO_b/34
VH>#I,WE)[#J.8KNPIUD/daZNfCI1W1)FWSNN63b\U.,K70C-_f[F]14K#9XIRbf
eO6FWb5=@G&TV/U4X_0bHg13NHOGZW66^A]+LSBBMRV9)_O:GKbEU]B3eJJCV3H]
)KQ=>T-[IHK:T&8Qc@g&Dd^^#-/J56]@^-.=>LKg4G_K><]AJ^[<0@1N+g()&>d0
I_.+0@8<:[,U8_6ZE@aNdZa:>Q=aI(WUAJOTQg_.#.:;5_&<>R\2CcPTG0)f5J83
1b:#6,:L-91Y-1HfO+SMeD(-G[)LgPV&AbO_B</YD-/0B4T(c,c>C7_UPId8]D_X
8.O67ffgGM]O+M&=@-CA@Y]TY;?8ZP0Se+9V+70SI>-M[(cfMED.<1a])VA[e)@P
=dA^_(R7(aTLARW&a[E]+BRa;?[Wd(/.CKcWUYJJ8JQ4K57I0U?3<-,e=9HD@2@D
Z3G]3<6;PQ0La65S_@6O6Af[bS5@W&EVeROT_H&0S,?fF0.gd-WO=eG/576<1U:P
Qc0X@T:6:U>DN9W[_Y:>IUH+T+_SBU7&=;=A/&?>\7@4ba70FPXbaK]&6A]g58\_
_f#85,A?-ANY.X5.OU=8ROc,?Kc#0J<D:HK>(,7@c]<;aD>5dVW9,1/e]J;_#OU(
gc:.6:8(Rg2e8SfP3N-_fLRC4CW5DIW3g5U)EaK-_ONH9_<#<8Y>]=FQ^[3N<dbg
0Se6Z/-SH3DF.8feF?1UE47g&bDXGCaM#QNeK\T\WR<7-DEWaKR1(:?aA96A5X,U
+;D/O/>fEP67FNO&a?g594^_R2WI2YNE\X1Q(bW#WT,VQ>&XdNSF1f=VEeJ-GB8V
5/2][[C>8EI1^LXRB76ec)>4OUCP-;=9G].f;OTB7C,\(]OI_1<N[Z/#d62D7@_a
D8XKK(Z>Rc>N-+GGQ;IS,Rgd[8e+TWU<WD98JU9E.]98S88TMOfUOO;/88U:1bYC
#,R4&,-^+fXQ,OI&,GP.\J-B]H>.Zf7?YC+)Q/A?GCOYdaBf-EgT4MJ9,0IdWa_3
Ec<VX3OGXJcFP19KD3V&JZ>NgOU+1,RLc^GGS6[PcHP02(W)-a2(<eORA7@^f[K)
gL;8c-N78^26WBWR3O8TAQ7;2ANVCT_Q-^W=(JK;0K+OGe37FOg#e<S,a]7>D94X
/MQ:<eL)>KaO>ZDL(&Qfg;g]ZB=]BIJ#X4WS?GKE^B<gTQPA+Za5[GX#;GRU&JMM
bOBOYX967I@8]U3cLZO28#6:4X<^UeS:0H?cFIHA,0<BBe):CGYEK_^#&T?E?R:<
geC\K;f9L)Z^3K8OMVVSV=5N3V>]];E5^+<+C1:50N?UR]B1_HQ=d9[QW4T1(C,+
eOH2XXN&:XDP;61\e1IGCKT:[H:ZRA:+d.,?;fLRJ.:_0RN\:,GPA8Zf@12OSUKd
,UFb4g1^B+DN6^7NVf&2HI-+0UU_?<;aJT=.7=&^-M#[I[9g,A>@41QE=D:)GIE?
DK\GD>I>+;OZF?G(XJR#B:5IIQeCWe\S0d]?PD6LH\;8&@g[FbWdR#GT(RWV+=F@
FYg-BJMG;VFYXIe#I4eCKUa7G/E4\Ng#UYI/eON,<Mfe1(+0K<>gbA/[K(f=SX65
ERGKNQW\E45W.D)5<77f27MS\I20\\ecV@Oe2f>3&M3FY,?49P6^7M>c)]FM,AGN
JONI6fY0f&#SXJIQBCT]][RWg?bcR&f6,;>3K9.K.a30._[f\e;W&P>BVa,FPMMX
>,G,)0dN9^);AWLIdYX@)f-=P&Y6fZWWR.F2TJN[(aFN)V5aTF0<2(#VI]G59BFb
Z-EHCI(UPA9;6_H.03JI<f&0(EHJc@1E<1SUZ-YaFMFNB[8\FA6bTWLO:JN.Qf;b
)X9D?;4R0BW^Gd/#dMN+VLeH@cbHR/.X:;ecdb]dVB)3aG<4d^:YH2V2(/N4e21G
633f@5PDbceZR7R7P]8_BX]_M/C_+1)M_&YMQ6/Zb_69YDFH0IfNC2^6cg>UY[f=
7(M/CCF/FSd+Q:dUfKYM.P&/@UE51SdV&B>bdS]#]W2gRLI09@R1[>e200Q6DK_@
@W&ZG(9-d?F(d#Y=J8I:E]9#bfL(4AfZT]/<6K8XF?L_SQ.Y3]\KRXUL:@8,3(g(
(..04:J8DYJ-#^Q^Z@6Q8FJ/,4<B5O>LWGM8)S[7E/TW-D_fZ&M&(-:f<T8YA@Yg
NGb=HYV,=;H^ab7?7-D7#&YOUN)8M)a3I7YTCCGX69Zd+86&;0N\MZbW-7a?)67J
c<.(].LdJ0#&8_\OOE?a=E0LIf679U1T;@LIE^6=.^bab5G]T[f5,fBZ?3W1MG7G
eZW]Fe)#^#IHX>C.L@M]#HAc<\O[Ob>aO/F420XR7Z\6A>E69E[YI+QU]gCTc-RE
/])b&;7+GgB0_.OJ#Ca^SCAJ6>2MfL-.Y.,/5:=]BcXb;-DEZ6,.<16Ode&MRHd/
-DCQ..YFDQdRJG9DI26[CaD^ZN9;+BI6DAKaZgaU1;RMR^C0Q6G3;ZT.b20J:(_2
&GSPdG;UCQ1Ub)5CY[NP(.(Q.(Z,[[X6eS?,9c@_&fY)7SF^f2\d>f1,.901[3)#
NXH52=[MWd=c9/;T4/O<F.<Jc4,Y.CgbV#<Y?+Y1+W@AeWN]\L6<IDKRPc=)6<:Q
]K&H9X38XK=/76@D-N()UcGX&Za;3S_aWg:EM_3]H<cgAW_K]0XX6H6,Z:M8\Ja3
bU)^4V)Bg#2DNKa_.9O8K8fOH7:U<V_D\/OZg;afe3_J1.If>Qb/5XC[^RXU[D+G
]3ES?@[U.?6bL-4+aMb(\)8AU\7QDOg0O7(:-Y&J^IC&U#a1VS_:&e[+]+?gf/<@
A23aG&AegN6@FYHHJP(d:/-B-JS/._)]f034&B=&.6TZ796GAdHbTD&FN8AQV0.e
OfDF.F7A-YF8b.^SC(WfCC\2YRSJCJL)_CKZ->bS_ZZ?QYb-cD)&VDY<DE<cHg]>
BV\O5T0M-PMJ-_>AI)N,+4dc0G>JUIF0\;/SFYP&Z^db\#C:K/#G,QVJ4A[R2#7L
^K]\;?YUX-cf2&]/J\:M/9,GMKM<J[a[cQ#2QH(5c+]?&\0fe,3Y6T<L0;/06[@?
4CCJ5B5Yc\Y:I@U3]aUbI1aRVV4A+Z<75PXD#(^6ZR_O/2,-4AG9<Nd(1f(a]dKd
ATM3A#GX+dcbA#@^4,C50,YK/P9PFH-BO#+OXD;<C&:8M,Z3WZAYM:8@gXb&<ddT
PO5T=[6W\VegTI&0E@(GRGAf@@#a3&QCVcN^SbU<A0c\WY@)GXP(O;C=6[B-(:eA
&E3--7.=Z5CB5VfRc?[?I.,>Lb=&c-fBe\[IWaV:P@PPW_Sac=JYN?1MSA_]/-+S
GJ#3dgF@EbY:XUJ?Z]PdZ9GG^.1;[]02_6(4b=7aA66A=KUHCe]E8^Pg_8:M5V6<
9M=J.^eLaVN5Ng0LVL::9_5bd+>RR.1X(:U(AHY>&]XT.d^KI0fO)\Q=QKFL7DO;
.a2A,=9:YW6B@>9S]R)K(6LNVIFUXDG.@M0Zc-YWTNVC5EY.T:4:YeI]59Y(O2B2
[P=8:9e.>#H9<)]EIa?=]0<)a^U.UVV3XFf9+;D\QBfHXGY4S^7W4][?+K4PYC-B
65_IT^ROfTf0L<9PQ#V3:;/WN3K(.aES_>aSEA</B7PWf&WHff;7(]1Y3K@8GOe[
R&VHB=UR(#27\X3c8(AH@TW[Ob<3OM67WP9)XLD46e8=]HKgIeG13R>U,ZQKC,=0
WVDdH?/M(WA<0=]F:X)EFB/D\[Q-IW?GP:(A\)G9)HcfDP7K5<gD3.Yg4B3e1Odf
E9?H_,-A#I1CQb8DCW8IFM=Z_<Cf15:OV[\,VF=D&)3b#Ed(cbd5ISN_a+;XXR=0
e8[&SXBa5gZ]7YEQVCQe8)[C(fBd1+PDH-QQdO_A0K3MP8M;d,c52C2C^HMFEg;g
B&+\cS?_g5N;Kf]3U99#:HAcGL49CI[f,5;HR]ZIBMB6Q#[DB;HP]\WfFR4A1IAL
AN)U_7CU)PDeH=\<[g.]:1EEN3N5c@Tc92^7(H)E5QZeJ;893\1@a+?N:B>CR);7
KS^F2H\&?P++:=HJ>c)RCPJ&QbZEQae@)0]05^a)fWAVF#W/-,#/V^F53PCd/ZPU
_c/C]XTWFAB@N#&7Kb9FV(W2<Y/_dZEN,8?9M3C]f#+DV+,=/CHR-\E0@+8IC\A9
b[N&QNJM-DD<73La(YX?X@Me+0V7U965Z9FBG&,P+[Y6a#IQ64\d.-)2)/6Q8dIC
&R</VOZ65(_&Q[b18#UE<NYS28?;22DM<=\#Q)EZI=^_,##VAA=&P0>>KZc=V^9+
/Y0+e_#S>=EOM5gOa33M,WDgb/-,\^,+fHQ=e(&cDbU<:U.4QK[CY[.5:S6S_DGN
3HH9A=MgWF6=.8_I753Mf_DREUF:bg6g796aY.ZFd;JLTaf0/BRg6QUJE21_QZ</
>.>:[_aZCf>0cBcA8E(B&,T?cU&4H]eL5VX7(B#d.&UcJX+<<Z^K<CHFZ_e^U#/8
gCV=HG[2gU;-N;&=K)5ARKg>b86^X))F#4-:<<Y@X?_K8NfF166IG.ER.f5(8L@&
+[OcD?:OK&dWFeSP9,:\/CE0Y943]_Y3,]&g&+1b];_-U<7a<&G2&&@/F[=I@1_<
]7BP2&/B7fZ_F5?XP37_]](+G)DP5]6C@2PdV,,c)c8g6V>I3gT9++JJ/WKW>X>=
2g>2#KQc.,1fL<Q0G^BUfM.Q)-HYT:WN#a-EBGSQZ:>O6>5DMT,L2Y4NACab?20B
9:<T9f+RYZ#T_A/eE9f+ECW+4fbWQ5]V.D[+CF(EDB+MX8G/Z6@B?b+:25G\C(QV
N00(0Bad6a2V2/SJ_^0I+UP-C_9eMCgG]<:7)\N+[)(^UB[eN+P0W.WE/^R28FNa
64:3_.fZ0\XVe.8<9S2>5MU5KL_,W(6KPeDgAE(;M#=5<.J0G^O2EHMK1.V2Y8Dg
PF+D>e&,-=1F_eaZ-/ARYg)@<:O:9>SKVV-3<:-0P,2BcCeG:-.c)^7J#E6&GA,N
PFGSX;FS0c0P,K/?-V=2]#:C_a4\QWOJ+\+T>Nd9L0J5CTQWC3W=b;BNT/Wf@XfQ
#FN0DL6[1P@gXP[\=e<Dd;?Mc4G[N?\K1L@U)P/YdVI;U-ZJ)N7EA<QZ@M6bP)J]
<,4)IZL;_[ZB/[VdN&b1N\UKXMRAcZ=]0P+M=E9>Q?GTbQ,3G+82TebUH8YI;>Zd
[#KB<_QdfB3F6O+cBN65eb]T1B@TfHNN@AVFV/Qc-XNK^Y;e:O+:VI#[:K[V29^4
9T1O0\JRTf_CR)Z)eaZb1EIP#4&Y498KQc3b<Z=Eb9#MAHb/eQ3Eg=+KaRMX,I55
U@Y#KTJSVa[_V9DV(1TCBBL9\N(8(,_0DRT<0Od_,W/6SJ(+XGX#XK6/NMZ?DK54
Nbb:&;KQREgYLc(_=CH:(T4g_^0-7:8K(]45SKPN(&22fL[d3d?I?M(aB>Jg;=+J
<<.HT>0(9_YM_)(.EZ]#9_2\>^>dP/F,TdB,G7NMDQ5OXd/P[73G^KTAX62CY\3W
@D/T5H2USDCZC]Ea>+_[&HSNCMgO.5MJe;P#:bKDNPGcQ?A(f]9S^&33eTUR?ERV
d\0[][?Ye0VM)_@@5D2A@_5)Ne>2,^\E:N0WLUJaN.[B389WK0@13@\?Q.(UB.^A
d=403HdKO7MM&B2->9>2Ic0A3LK8>KHT;MVe,(V2)d[ZJ0Pc8IDY.:L1]QE9fUb>
f8D;)]Z]>Y-@[P/APa[+QE6R7GMVWgMQ52U[GQ[J>_SeWH3b2P91N#7O.Z\>4)TI
:8c)Y.F=OZSV@CMc/TKPZL3OcNf&V?a@ALWP&@]TV6UAH/&>LO:[dcW.@]XR7@8_
[<=LVc;cP8H?2#9@6NgGHf3K.(C)>?TQ/gJGcT[>&X?-]AM,#VP_2N<TMY@;;D+B
e)Qc10B\63Y]2#C+Z@SH]90&U9(N)af((O)2W.[IaMAHfQMCc&Q03^C+8b[a].Uc
@RJ6J).cGRaIcdI@/<WbG#;5_NWT+M</R[:(ZEUc5?Vbeg@.E7aYB-ZH_)HU-AYd
=d2XC/&adJ&8US=5J@,R&\Tg+P_GI;DJZHEXDKO0FO0#Q.HQdPa,4(W;Ic_XTST\
1E6ec]b]B\/GJIDLEC@0]LDd+A/bfZ5W,]S</?\3c_GB-ZM)-eX)J-_T_>_H?4N4
He0XcUC;H;\0c;cH9c/(baM]f.g[5I>V_D+6?;JX2YBee8]HUQf&F/?35e.7K>UX
28.3\Z9=+XACM4,]W3W:e)?WZWMgIL4)0V^(8e+K(J1=G#fE-_<2Y]U:cI&,,>-U
(E\,JVU4-\g4I?7SL]ZH3?T[I,Q4BZKP4#B.QN^&ZIUSLgbbI#>0bf7SFZ-BSNA,
WOHGCeNaBPV1;)\A8b3>06VK]I0R=VJEbGg.HH^?+>/P3Id9O5_dUNRT?/AgS#KV
IIK1<BaMN=N26J_L&;Xg/X/U50f3#<cd:6LE0-FQc^RSAFPOHB\(Z-],\48O=HR:
N:N#GPb:5]&?24P2B6?GW(4]]9VPQ8B_JfIa+_U+R:>>/#fR0M.&8cP43#>/2UJ+
^LEfQKM#E>2]U,]?.N0DePS1:LH]282#Yc96_B-P)?f1ZXV0>?I.<]R1<MXPLX)&
FgO3aSVa?:a[;_T=:\a@54(PYOaFV=.:M\CE&ac1-;/.dD+X+#Q-IE/e+PSM7eG\
LT;;:)=<Y42bGZc]gQNZPX9F4IE+((Xb3eM_gSCd5^-.5&>Z^I&fb1)ARGIR2Xd#
YcGAE#2)&C:0(VNT]L4QC4F44&f(7DM<KL/E6D71ELYfQ-8D/SO&07O2E\LLWK?[
/e:]J>dUAUK(?>LaFR<\HVH8Z+7,&14G#0^.J#QJN])_Z7#T7bNf^6[b-CfB=b9a
--2+34ZZ>D4X),D8&,JEOR1RC8TU._5__Y3/Pc4=6Fb8e)8VLJ0aDB8G0S-.fA5>
H#dbXGVNRY.-.;L;;[f0P1eaS]?72KDb;EZ,?>T16K\>?&f)_&cPP[-Tb47;S]aI
G>KOLNaJL@VKS=#AQb(+XEU=[_5L0^MCAQU9_3YeY^N8HH3e9>YDQb44Dc?HG/?<
[<F)fR/K6)BZJQ;SX_]OI^0>BJB\7ePUWI1ab6O4U3;O=RZ:\J6G-.-^Z-=(8-[6
[IM?7&KQ+752ME_QK/c)5A,1\:49=R9KR+GMd7^^ZJI1V,4B2>K@^RB:)6N?g3Y7
\Ma+Z[e=8,UXM5B?UXE<W56;UZg-3g@+DYSXeVXMW,UAL@)L7bM5QeWYd,MF@RX>
CaUd+D/[aG6?cHW>Q899+M88^<<TBMJ_(Y/A]MFJ8N=M78AHC^4f]9\5cAW>B2@C
Z_:L.(+6Of\<DEc(X0A&.f(>]dI5AR=0R]@4cK;HBLdgG.S^/_Wf+IP1TH:W[@24
;[:)&cIb,7RSW#1I_2&>QW8EBCJa@5fI&HDZ[U8IPU]<5K9I3a/TIZBWg)K?;:\;
_RFCdA@Xb75W@fGD7K?V2,3K,@0.M-d+&AHPGDb393Xd=)/f<+6+>gF/HD._#fS(
/)--dUUJIZ;77FOKf][(f\\/<AR/B0@IGW2g?NOOf_,U3WF/--gM6VCMVA.N4@3U
d#.>?SX7[_fQRDZ<;U^f@Z42=[]b5eMd=@>NeXZ)IYH2+,P#8#gU0,(RA-7__c/e
GJ&@F1g1U[(g#G608-]WI^B(&Wc-+8=:0bXXZ4+KOW@VX?>Ze77(2Z/a^)=GcA^1
@I8Z#NVF&#7bM&RTU^4ad9+6E6HfA0IN>DFH;,20D\L]&OeQ8>ZcNHgT9eg)G0>[
Mb+=X@XJ<d(aBYZ#,5)?59>;&,CYZ>3ffER.#GTD#K6Ne[Vf1OFbGL=]?ag_Kgcb
.cM3F^MP:ST&TSO>+[DUCJc?,CTe9-5aA_+LNSG,ID@1=6@[+.+:b)B,NA@Fc<QY
)^aG\E^=Y5T8=CA0I6Fc5DAZaH..\N-1YV?Xa21ZPc#:#49aEPQ]b(\))#JR&;.A
9#:#_]&,:@(E,\:\8e8e3GDY;2^Q9NR0H;31LQg=C?ReDaB@66/J:GX:FeRH6@YI
:c<W9AFM(SKeG4):J456V6cXb)UXN/@Xa\\J-,4[47.0X\Wb.B<cU>6V7^J_K4RB
]&GX)bI;gbE6S]^.;C<\7WFRK07D)7KNIDeEL]RE5O\^:]:MaQYLH9L_aBecY#F5
L)/#B&,S1F;[J/=@NHT&[3ON(R3d1]\@2[@JJ(G(G]:NXGC=3>)NEO:2,-VIW^[R
&8(?=^XH;;RG\PNd@dZ0:898+D:ZJ2PQ^SYYON2H=:2C>eWD[ZOWBaO_ZGe8-;]J
2W.KB3/OYSH#B\(HE99Cb4[:71cg3PH\OW#7S<>>QcecYRC5/(KeXUdZOBQGAK3_
F4Ac:AZF-fgUFc#E,[S[PO:S[_fd2X:.6N93b[3];Y9K:M/3K&(I(b]?ZZXA=.a4
33&0eO/DV&L^<WKL9J[TG#M^0#^=Y69R]&;=?:G/GcDc45e9WC]GQ2N\S\X&(]80
AcF@HefU;Zf;CFJ_WN5Z=,82Lc9Q_;6b5U[8a_7\V)f^7@@__+HAED/fLR2.U[JY
cE2<R7\Z._9,3J.WPS,K&-Q_V]eVN8(LP__3AYUQ+10H/Z7#Pb+WYM,=7ICH4WKF
Q4VOaLWUYFR^=O,68@PJUFGE9MEE2Z1#b]W]:;H)Z#/T\XID[I=.b,NUVa8&<LLc
AVL8I_+g^:&^P+3R,(Z80?IA)K26887aRA943<DENeEH^Zg]/_49La]M0-,>R4V3
C<]L/g?=GW2CCdMOa\.(BaN?<3.,fg[N_1-JB4##XTJV>?42WUSDgLUJ+<;Bc>NK
+HK_[.?B_5\6X_6R1)0IMAb,&WO.E?XGEdfN5G2J_cf/NSH#A7SRR.7XFN/Q8c-?
)W_F_].RcK;@a8JdB+J_VN/Q16.UAST#X=_)+^SI?I<_Z)T?MB#[3K7A[Q):Of<2
I]IX;fT6[,gaeOb;W,S(P4/JfHU.LM6V1GLa^Z8Y825GN^<R1dIWA_GVE#0@eAGM
f(3Ee\#O0P?A.\N3[dTD/J73_CBHZ^Jb8H>-93]Of6#4_e>I2E>8CZ3dMZR2VZ=I
_R>.f&0Wa)H-W41.3:c)(M<R5Z[JNB:DFK/3JUe6>^,BF(cS\>.AX,2a&/#YK:7R
=D7/0^dVGbCbVBV#^.&,g>OA+dZ@)ZGg^60,e&V&TV_UC]0X)P=ME;2df[KbD=ca
0&D1+(:TMKHHF9-XNE0S4>Bgf6?L:6M@5UX417D\F10Z<;5Z>:1Y0]>Pd=@?fcVC
ZHbMF#2gg7TU.R^W+D^P.OYcX4@,VGA961X5CX\L755]3;UYF;OFe]4SV.b)WAa,
g6SI6V<2T3#ddf[=U95G5+XbZ/;?R-FXML++/1JDLb+0K.LOC^b)E_aI6R-4aJ+Y
#+HfH+H4e\R^<5E=0Z3)(4(.e&@P>T9I-^f92.D>G,OO71<bAJLZ=+G>aUZCdGd8
GH.4TT?6Q,ad..PK0>9+V8;>HK0d0_RDBTP3dML/7V\,+OQ9N0.a:_.8>ZgPZ-XX
H5Z&8@ZCSg_3RgP\WC,;>92aR1c3S(VPDID96a(?IG0Fb7a0b\?;\Z>;cc8a=O2\
#DSUM1JT:JaFAEU/]T>YHBD0AF6I3.9fQ^QeUB-C)#D];a6WI)7Ld-J(Y^ZJJBc-
M)DYZG;J4/F=<RTH1XUBA(>-1MO^RHEY)<0g5^E:U66Yf1S^Kd:C(/ZJ37I;<3,0
XeP7#eR0/Hf\?6)<g&;Wd?>U^,DC\6F3&2U>GL2@K.2H+N,aCV8^5GJ4-IW3R[,2
P\MN_KKYF&f/8<J8aU>_H0E>8865T8d>5d.gee2Z\MF+\\10VK[0@\NI5\1?3YEB
cf:Z\H2/-B4NbUE]NaB<QG)HZ3.b2Fa)E)ALKB29>EW+^?Z0e+_=H)-A0;P\^C6O
Z35B=OU+g\CbUBPg?S.J^84AeR;]I:1L<0CJf<B3GL^Laf#7b[)[DBd>H:35Y?XL
D]C(Q(O72<X2<[LW.3R<gS#Q8@C2[X@NO[O+.K^LZg0ab)WeGd0OT[TTPY:\KB(e
:-+EUdF[O\OEYBVa&cT^YC4XMW&5cJ98TMQ-/2Vd:SSd8/Rc][S.-7OKf3d_II9]
T=N9cV-[?/8W=a[6L<,?W1]YY_.=Vd(a4>C5>g:9^-<FE<H;IMJM::_1>S)I)?U+
Z4_K5,bZ3O8WfMD(_b<X4,#3:=X^B1^5BM:T/;c-YX.1S27DRN(<S0XcP;A4P=eA
+2>9.<_VX^b\S2X?X8N(^GFDGIW&1dNO4MNO3^2BNP/<TQ2PM_CcL/bK/KF4578&
;Ng7EEOLFW[UXagW8+DZI/Qc?,=19g+26W[aR+QfVJe368S_cCgbR:d44U34WS?c
K:;,.dY@gIO>bKYW][-5E;f6@?eE]@D=B[K/(E>9fSH+Pc.JZ7M?E4K)3UR+]]+K
5a]f)B+K&:bFQ_I6([8O.:>c7MLBW3@T+LRb)D[c,S/D#P8(?^TSUE/a:S,AL]]N
a3Ff[(N]JRLM+6DTNg53=ICK(8X=-Qf^&7JO<N@H5Q.C_dCaU-d&,3Q^B<<EVP^=
7<+PH8M2.\aI[1M)A,,,Y<Y3-1[X#QS6=PDH[Q#(bb62MW21K)>ee<P=OKKaJeF>
eFLeGS(=4I^3;UfP-WHW6@UYM-7/;+Se5>:VDUWPJ<Q\<B90-PJRAJ3^10(cW30U
P4V?-Z?4?8\_f<[\CYGZG6CgP#I1&d.]5a([C8,>XYb95RWJ<gE1dZ9#&3HPQDR4
Ff1-?+:NK^)9bIe2/\>6=#f3F_#bCV-ETa[2g_@+H5=N0-MM9\XUDFg)2Z(BSO>:
aA+aPKB2?)T,0,?>S?@^J]?X+V.?>J4^7LTK31ZYR1@K>.;Jb:+#\R.5XEY1FMIE
KG(MGH1@^2;6\gXdOQdU_#8L&?)B>.)SNMN;=RHQM,DC^L?AHabDH;G(#F;)2#(;
54W@AOQC7,c7Fa9C#29D_#SWXAdPV/e81c5GL#b\?61WXa9-\E&SHDKG/PPI5.>d
C)D;/2#IB6?9UG0\PD&;MW=PV&TJ[(:.69TGfff>->Q/6)MG3Y>WTJ:8NTAFK+>E
@Z=2d&0F=BR6O;H]<Hg,3EcbeO:G,9b=[J4XCf2-Ve-6IbRGL/4@,-d=d2WCgV0Z
@OV/G9;T<;Adac[]G5I-3G.X&]BR2ce1CS,\^=JBNJGBVD2If=/VDL1g3N(9E9Kd
&C_1Z.<eL/T^V463,SC>Sb<g/)bUfD?LPfeD23-2JO>98_>TTeAa\9Ua<O>Xc@^2
^]6(#P7caO^e,I7C]]TIQB(+8PMaF0>ZM>Q=<37G&#M,caD;Vd+@:]aR.EgVcH,G
=9+MeX(GAb@?dX&);R=F0IG8(=dNA0/:YIEEPffJC?HX#EV1-Y,1&,OSIR6IQC-/
LP_.fVB<F@8R#RC#I1=1G4QWAN[?\;f43K0;5:WcS]_f.M09+c1+F3N[V0cdED15
-<,3Q6&H,-c0LM7N3>MT>5QUDV28Z-I^VGOK)#6[?/HJXZc;CQ_7fEe\93B76:ID
:R(;fW8Y4daTV1,?Z(GJaW<MZb4)cd_N\VG81]8d;?F(VfZZ5Y36_X,]@[LT2O10
=E?MP-6CYZ0)E.K]R(^c]/.MeFCQ@8X3<G;<55-::A8<MUd\V4OgY&\gg>KGU2&G
-()BgE;E=2?ee@<D]gEEM4IPJRG4@=;U+L0](dcg[GF0GA)#_0?5TbHU_1EK<9_E
Y9HM?W>eX07;=3GVA8J7S+9P91@+T^N+KAe=<2O@DU?9_1H/A7gWO.7bBRa0W>09
<[;(NF8I9K/7<2\/VW&^OB_NO5[,SF;#>1890@a_X.cQ@M/gSf=bKHA<TJ=5>f,?
&#50^g;N8+a<Ma]/U@59DWC-H-+K_]b/KRd?EMT[3LX)LIE/=(\.N()7:DSU3D<V
550^<I+BafR)e^fB[fJf>Ka+#U,4;>VHB/VP38KG^U93SVN-YDg2S6,d?:RNf#7/
G4DY##7_3>5+JKgOVPa#f-UgPV2]M_=CZBe1S3A+O#4DP29<;S9CbU=N[(C8)LbT
dJ4d6cV?UYQ+Sb<BcIMN0Zg?f/QMJ.8B8>@OD-F75-+ZE0a>PEdfH2c\:e/7e_fA
4+cI(&^,H7)[Hf<TMI]Z]DTNTRWRT9L4fYY-/C;UG.e\HdF#L\JV7eS:[Tc[?cH<
:/eB8AU>FgfOL(15?C/[L&J@+Od&3RZ/Eec?6A?Y,+4]6D(=NR0]E:87YFU9K@?/
TOU,^[1^4gE/0/&.f#C^I>c8V9UKX9aC]K/eYF_#YQCX1_S+H[#,?_]OS^a0.UA@
??\\EPBfCKcS+NBCE0TAQ6)Q2g_D^W;UGVQU[B0?[L,35K/O6&:APDI7N(>XGace
e(H9K7I[Zb5XZSQE=E[Pg8P4BOAH2@?)5:9=)GOcBX,VEcEFX10fDIQN-3^A;<K.
#&84A=?b.7O4?U@R[0e;M3(.eUNNZNH>4Xf^R=_XK?d@HX(9E7I7a<6.P.]ZEb[J
Z\.FD@KT[0DLG^SKZ7=@T0(\?@PH^X6SM_(aegfMDHV7;F-3ZM(;:?V;67PSb-Q8
6K,RS-FKS#EeB0(4FC(?\K?+@Dg+e+8UH#Y4Pe4g[A_@]X8).[:d>3e=fWV,c?aT
;5AUPCQVEE)PF1[4g)KH<87O3+70+LU&C4KRQQ[ZTP[C[8&M?63cS:[=cP9H0AF6
f<QV/2T.bcgGUec5E.AY&Pd8Z<+MaVDLH#&2&<X,/8QM+R5/7LRF.gL9(5aTS1N8
[,U11(Y8<@8M4e5436I;E0):2e7:G>0AMFEMM9I1<C2VE?F.F<V>0H3gYG.-0[Nc
cI;7GTD1,7-_f14RS=.G-gbG3JS4@c@\?UCQM?f]EK@:5bILEK;TFRSN[V+@F75F
fb>E_4^eJ^0&IJ[,VOVf0W9HAI_2V?^fWD<O8,\8EZgNIMB(b>?:L83G_SB_4#dS
.@>Q=G(9VR:KfU/Z]7#U&W=O<\0a^AO0;TR3<BJEQKS_8BG7Z<EW.g\/.ZEWaX>1
QMYP_+.)Q&>C-]<CP-eH1ECd1df])I]U4>DY758gH-J.1:6PUEJ]F9(O-LD\Z70\
Tc/\PUaR:g-gJW6J@6M7F:^J=1QCB2?A-4WMWWV.AH^aINJXZ5P.Ff=/3cO:R\dZ
[4SR.5__K6GS7-b]LUg+5N6e9E=?^XX#TS?Y+#K6)GH#7fP-.UJF30H>W&L3c]Te
(.7V\7XfPcXJZV:c8&AdYT:cMX9^9JV)&0EDZL>/S,LK[a>G&8B^3#EVDTMRcM7T
<)B?=J7K@@aJKBQNd3^DZAd>CX>@C+(.>].OAa8Qa[2HY@/8E0?[4A[-+H38[4dc
QY?afe:#1&4[F-6TACEeQa6dJJ2??f)NcgI_Y2TU+Y08G:EY441PL5f?R?8>I8)O
LO(?2T=:=?>M0-0VN;.DYX1@9a8_X1N/cVUK/PfP,V&=W+J<)CDf^_cQ<^8c^O>e
83ZS#+CRJ>>EX[LG+]F8>O[#09T4JES6P#SQE4;[]M@EVTMeXM0#91S^)\)S<9>U
4SW=\aHJ(<GZ^adBfE/B\cRDCANEJQ@QIb?2ab5FT>[0E8_>;Ogd32e,N54#F0^2
_XJ0ELS?#1.^CdBX6.^72gdUIB=T[0[<3_=<6bX8T_CF,>Yf&X^Eaf#9SP[J70f6
Y@Sd.K+c+MTK2GCd+0VB):Hg?Q0J#K34aY4BYGL(4dOMK2,[(WFS:P[892Y)S:=@
CX@K\H\?.U1NDf86(<,49@MAaN>=#&>>&U,0Ja:4a].#OSQ2b,/E;?<#A<>]?A/8
MYAHCM_&KOd]^1c<5BKVT[d-S-PEZ&;+^@FA7e,#JKCG]b3D8,3VBKU1b#NeYReU
Q[a]Zg-aKWHd:0;5K5;MNTJg/=?dZfJNC[#+a8.FW-:Z1<R2UM(XdXTbK=<293L&
U8LT>3-Q06aZ.7)8O)Ka/+L\UK<U)CfbQSGFM-W/[]CcG=.YJN.fV4geJE6#ZMVP
D59^gPB1&RYW#CF<1(3gV#6&-Re/M,:_J[3B[?,4Je@9CPTbW4&G#4HN]eYTA-OM
V7D->KCCeUN-M;gc9<]g2,b-3N]Q&P4A3&ZS-#?LH9E8NYeA=O7SDOX,2DI@M]\I
MLcRbW7d#;ReFJBY3/GJR4/>HbC3O1ZONd[[g)^F;EU>eM#C=H.ObKJ4f>cBSK;W
)TA5]N:^V2C6bEQ/b/D)\WOW#ZRK=9UEfEG-<;)Y&gR+C?BPG;Z1=ZP/6M_@5RL?
?^NQ\M9OI=O.4NSA^3U4A\P9T.D]L[-;c.0>4VE..AgB/],1C64CCaI3ZgHT^U;@
@###BaOeYL8Z^P_0L:^Y6#XQ>-UAgNJS[[([_G7L^NZ-H^gLOf8I<-.3dD/4D;ZR
dAEd3GPc#L8NX;TQ^L>V1M2;g+6#(3J7KVH^+FgJI\DJg(3WF8OXcZbZ9<VDbFA<
d#bZWP5-P-(0YNB,UODM4UTd2B9N0/.W^C-D?d-b-^:gC?cO>71#62-<3&LH4G6N
>.&#:.T.P8V9Qfe,B&,XJ0D88_\\:&gGKO+d8:Q32g^LD8FG5)X@G>[A0_R6IA=4
Z)fT0O7@3Tg(Y9QBaKJUG.6)/gB]U1F<T,GO&AK#XUXPS/]>_d6UFB)TZ9BTBTAg
&_9QD)WbJK;C<^H=/)?C?^&0HEY9]54H42<19,cOM=&EAeSJcda&(@UDF_efWc4\
>;JV9IUEgR#f;3MPc6.<93\Gb7Lg1B0XK[:/.BJb.P)BXAM8BIg4&;4Ub,3Rb\#P
S7b[.f1HCJ3]9D<FF,MDCE0I:BYRQEIQK<SUERIG?ISJP(.BIJ^e06\7:Z5?]_+9
CF##EC(CE19D[bVbN0?)\A@Y&BW27587JOARIWAgAR:f>(WWfC)c;V8@FabNGAJ@
@1)08EBEI9CB,U:3@-#e#)b]VRV_^U;&\a5[@6Z5AW7N,X[E;0E:(S#D2W9KeL2N
;(Bc6cIT@(ddPMYcBZ<QY7A65-X@[_./V:27JV/,L4g(b@W8K-,8TWLGZL>bI+#U
D6[>g(cP4MT(K80BF+)8PP\.MTC/UdQM&,8#G-N-IJCaV1aa;W2GV5;(Le30CC,E
)56QRD7NI)?>Cb\LD-UfO0a^7KUc\W:E1)^2.NgFaFRXdL=N=1D;,/&N#Zd-@5aB
L:3T8&M&_H)/d<QXbS]S4MFXKe:OcfF)K,08[ABJ5gGd=ALeGcg,JMLFg:#H2=Ie
Uf@0X<F.FN9NYdN8=IN]aA.R;aG>.Y8O)0=P6,U]Y1_?,PD/?0I>C2dXce<>#041
\L/[GP[\+\/.&(BNeL.8e^3<IU#bLE;C3Fd&OURD<)BZbV##UTR7)4Uc2A5GcK>U
adS)C?cQc2VKJ7P8_@dT:5))B.8T,0JE,.D(_3\RA(&IF1>#fLBL-eFA6]=PH9?G
5M^H[]9K8QH,O0WQU-Bf<NL+I1WZ_UNH_4F8Z2#H+(MBM1@IN^;&A5I^&X&Ubg4G
[>,W=SUK&#D>AeJO4b:HGO3SWOdW4W@J_aSBX2dEWYfJ&_T&[dLeYXFR8VX]34>0
O0<7WU&4,-UWbH\f6J&CX6O@B.8[5a:O.TTXF&WO8fD@93\Mg4LQVCTHZ]LF7JAP
+ga6P(.X;_\/14-Q2I1_ZgY<fWcD121&fL\PBQA?/+X/S;>\B)N>]N=Wa/NR-VS0
/e36@O?)X^TKeLV(K(04.Y,-X0A_a)(Z9_JQ8=b^=@ZC>#O7:M8D:#VCLdTWNc\7
_C0#B^#Uf:gP)I-U90UTDd2HS-]?XQH[==gSCTX<dA.S]4<ZDC#<AZ@5V/ac,e)G
#EcLdBaV?_=+=P:\^I&I:Y6_QSH-\<:R(^Q9)TZ+dgBC&BB=Cd_3Z4cOa1^O(b:/
J]5OJPYB4,?g44VOST1Oa<c>GN)]O0I@Y:>e@IIDR0-F43T>#Ba=)=>[f[N7FG=;
Uc4AO8GP;eFf^#\S<X^V(ECD;UcV912J-Z&A=-b?I]]:M^^JS_ZNTNB.>TcJ974f
gHT&9@RGE;JKg,\3CSH9_A<9fB=c=J/VN<CWbAS2/16XRF47OWa^RDIB2RAE(V#8
gF:#^4Od,]SSSNP+S[dPQ1LMI>QHL@<>F7KMA\.M2eBDd&U1PBHHI3\)J^JXKD&I
,#6SF[+1<\AH@Kee=E_NV@+A0HURe\J8ZG76E90Fac6U\GFO@W/&RJJXCI,fRZ7(
eF_d6WaZV@XOK/9VW)SWA[USOQ^?VVd82.LaY_Xa19_f97XM(J9Z>S@W-C4@-@IQ
9S<R&XH:UU6TfG5bdN^dg@\,?5T3^#HWSG8d=TC^A3aGeJ2E4bETfNeCL89Eb&Y/
Bfc9/W5BP.V@63#&CE(]^/\F2:C9[[F\7+35,G/8H?Q5S,>)O7/SE(Q<M7d68<Ve
8@BHUF(8?3T.#6^=LBTfbQ\SEYgA)0\[c(UPB&\#g4HJ;[#+&#E-1<ga2/6BQM@f
=;4HY[eaI^#QTTE[@T3ZcaPT5KNZA/=FdX)eeY]d9Z(Q31V\MX6a<A\Pe,<5KGWM
+AZe7O1P3cJ-YXC@51_NZ]bgH5VcTX_XB5Y:cV3U<>5,O-:7:-gR_L.WIUZe\4-&
O9e0KH3BS[[\aO5f?Y(\Z_)gOS6WJ/<2SOZ2E5->.XJ)#g6O?e:daN.@S]O>WOT7
[XTf\BgfXZ-K^OQS,RG=\YPL>(SMYL)MN;@;LU(/MVP>9H0HKQES]MRIP4TG4]OL
e.=OB((dY^3^BPKJCecA_OG>C096J?#a\[C9W:KD0#>2-JAG\PZ0b6Q_5A5F&D=S
PU#@C=(Wa0-\?O2V9\W0712T\[EaOZf]YZ/66]?6cHDR8g-O&._OC5D4Q9)N1N+T
(VbK3S2D[+8Y2(c6_14&EDTV9/[D0COQOF>XT)2?HRG59I^]4A]f.4MC2[R5MNT_
KR5e3g.:H6Tf_#@D1P9]b5b/-[M-ZU9,ZbZTK,d0+.LJKF:/cTY7HAOL--,^J7Me
/6^5:1X2bEE2)g#7BH.Kb@>NRCI65620\\UP+U]gF5@X/<9?)_cD1Q_+()g,dD\J
+>R>.Nd]Q.H,&DD3P\.T<J4&323_F:8OfSQNfX+]MP^\Ib+Cd#CKLE>Ng.22(:?B
E0<^^ce#9MRWKUTH]<R&^L3\VXgI/55/Ob=;90JC6deWQ+M@]?V+fHNZN/:L/,6[
aVX4.Wc\Dgd8\XeO]PdRYP<XTVf/B/_f@&ZPSf8#HC69gfcK79)S)6Z+CF(ZWOCD
@+IHfJYZLVNPHfG;N.[WT.V6<VM0RG[S]HeAWe3HF&N^HCf)KV6,(4OF<8[-cLG=
IT8TG;fd\aSS^Re1C&Pd)\cNE37]Dd40O9U[e0b>@CD(C>E,^V<+0d1HQ63FD2<A
N7B]eSOBA@:Pc9:0-RZEU/:RWUU=6?d+4XIJRc=3fT(Ge=+B)a#A.VJ/_>70[LF9
#KK4XFfL2bO6Vc=6Pa7[B(/FE7.2_AJeDf^Ye03\=J&FH_TUaFdbG(T5(Y/e<\W>
PINZ/4\/6e;],/4#\L0J[KI-^TGW_2(1@#(F/I?\LY8B;Q?A>=T^4R>1@bf+><[@
;:-8VI)Z@0[J4T<S?EEGLF#(QK0,<WA\C/d_O_335C+[?/3bXe.C7,4cdS2-]._b
[PcRO^Y:Q+fE3L):SV9A^<M&5P#SH:cg/#e5ESR]GQ;L8Z2C1:XE3XRXA/cMQbT;
P,5[7A-^7I6\b\2I78,&&#/@/d-G.D(VQN6XAE?VNP:HHSTdUW51FE,R38#L<PTG
^P7)dXWJE04AQ&22-Bf-cJ7YAI]_#65JIB^d_&:0>cI2Ab(7-7K[AI_>fE8We31O
E1#eZS::?PUZ]9Ma]c4<8Tbg<eP4RXGF=&QG-c.DI)fKO34F#/cOTP@AAadYFfZ9
O3X[@98B?D^Q@;[JXEMMSa?9O[WaU=(0P&^CJ<-g<4_-AU1F/<OOCfCX.@8=\3.<
a?;@]M1E-FG4-DRXe]Y0:TTKcffFF^<G_&N&PD=.8LD,^=)YgZ[U3?#36473^_:G
@()3e29JF:Xe?5,=,LO\7T#Zc?E&5P@V8M29AOA;.&?eZ#[0#&O;+H7bDUdJT9WM
X7LMgMY490FH.][:Y&NO.(YJW#)ca8bRN3AC90&YE@36.BDH[U;5>?b+[RaE8:M,
VG07aZ)A1D7599RFAG3bDO^G:EE;;Ye=FE2gM=[;P&ZR4+f\I5X)W9CYa+Y0UA5U
1=O,aO[&-S-77EWHaD<-)\D[T;<+YVf=X8?GSKccT:PIF+OX/,\7/5WJORgU/-;F
U\5U@E\M[H]@gGK=42b(5dB.-->LDBZNX_f@Ud+UfK(1:=^UTLK)G3>R3#P5_+V3
>T)e4b)ER@e<MU-@aL9?U0WZ?b@>&31AW7A5dG#=d:@+X<g/?+@?=U9-9^.CJ:2O
9TgE][5AF+V+eHGIR>?-Cd])6^Tc?6E0T[4TG\#>>,S_OgV/91:CL-S.[6A_8_:V
-c0<\O,ZDG);A#;4#^RD._We^FHW1ad6[8:8,^<0<e3O1aSGGZeRc_d;e-0L43d;
cN-]FQaa?.:FZa@=>de=9B,=._UJ0#\OK-_7O_f3<8eD9K1;dJQH@g/O.5ce4fP+
],09_2#OQI\YP^6;1J_3W2c4G+-@#,RKN//-fJ;IUO]>WZ&eF^WV4:DXMM[.ZWR?
UNbPc27Q8PDY[AY@QH]^LW\K1E?)D[27=;+UL+QdOUIgNAHB]cP-BMDUc<#W/Yc,
eCUE,)P[/X&3VVYPY;9?UdE5d^Q,00_?gJ^H#+2X.3@D#(3\8JZ6ITaM^TQe4KBL
bTVRH<^3eJ\a9+B0_J)\cEZ\8/(Laf7PTW_:7bXF01c0ZPT40UP=^+Z)Y4&6ZEg^
d3N-+?Va;eV+fZH2:38@Xc.OPg3Kg=3==6B-1(=ND[5ec_C^d\S6aT16S3dDZH0=
(SGMC#P9=Z)2J=4(A;2(dKe_Wf(:0-+D<_AM-GK+F\&LVA^b):.WM&=6#(DDCRL=
+7M(8;XI0\_gAXd@N+dJP3>V5&U)]HQd)Q35?8=)Z<(48d181A:X]e1gVBEd:30G
-JAc=GL3QE@ZT7;9V:^[W:UPT+[P,8(5dg,/T:-L^PHD\VP,8TKb9CB0?T(,75J6
/,g#_><=Cf=afE7Y6(PGK6>3Iee4MQ2OX--QK4771^MJ2[CMc&HA0KQ5a&CLI[Q1
<aHB4#H)<)V@DafU3=^5NY2d_4P;]eTCTO]:f5[59Y3]F9B1H+-1gTZTF=RL:MD5
<MEA>S4]XM3Z<CTL@6VHYMKb,V3_I_1P(f5]3++ZT@9N0f&DIg:^]C10]d42\86=
N\^+<^/_GQC5a&S[ET)_]#\XW57><@0EAX[P^0_5FQL),@;HF?HJ?1Q21.3=0&KX
.8>0QRG#LJ;P.UO<1e94U:/2V()^69QAE?5,SDS1\D3\>@+DXH_IbM8>MG8\AGaS
^YRfAdQ<4B;2V339(-[e@V=6F@2IgR0g&CfLLD_RUf&Uf8D+U-JG?;)&;-[++KSO
XYYP52YED2/<16>VaH[PF[(e8#>S.3g>X,d=E4f],1DP;P^=.RB2Z;@9WYC77gBb
ME>]I0b1VP]>4A5aXI>Yf)[M#K@8E<FS]S8N-(c5dMd5Y@Nd_HMUWI)P#M];&DD1
caF6D6b(QM;A8X9B\[ZMb[g]#>EJAH/QXJVK+eGATY,OAceQ69,H),#.e,2NHXM=
I926IHSMF82]-8]Qa79g1^\gJ?#.BW&Q#Z:/X\VKMX&PU5L@+VfE<U@4]1[M[&Je
8KM^5c+GE8V<\XN2=a#L]&#1(H;X,ID9XHJE+YPJ=B8V4\;NVeMY+OYg9U>+SCg5
39FS7&9LfRf]^5;/c__9;<KP8beSQ-e@[a5MKD+L,#3aP&;QS87H&f7IWQ5F_WF;
F2&^0)M^?9CMNN?V?.S[[8:?PY?<NMd1L;,F\05@5+_Y7^?5UXF\/PgZB:;<39\Z
U:Z2_P,bZ1aTMQ4+]B?=Z25B=Pe?RXP8(O+,\bOg5&3VEPV0P[5F6A[b(H)MOSYR
HX=I9ed.(O@\ebRMFUOW;>RLUD\(DW:),b([SR:R<-=@CdM\@+98bf7G5Y83#c?-
P8#T6>+>c+^F3C.-P-C\G&M5L>8<dS[a?c:cB8ae1W(.3+:H7BKH;+e;bf]0-Y+M
4+/Y014KNc&+MP/9L9]QM5;A\N]<N_c0(EGATRF55EHT[5=b,N^6PD7f.,L(CFF2
NIZbFS.,-6d@L,9Ca^+^aT,F+A+)@b73F)^MD,[2T(;:]@2V0TcS#>Ee]1<5#0Zg
&+KS0:I7TA3YIOCfT)Y+(7_@E.;]IPQcD40]FB7Oe/VW<Ub?6;ZT?9-H.Z[.5?+W
KX48_BS&HE>8YN2:FARA(D+g>8E_LK9DUZLR9QE5S:>?6&NY]5NSZODF<TX0[)f+
JWc1;<&e6)P8XROaCY>7d11X4<WJc:2[0Hdf[XJIY.c+FaN?94<&J48FRJ1OSRcU
.A&G?)4f?bQKQSHWg;R_0.SV]^cR@48UNN=ZA.KI<]UB&#9c7X2;M:V(8UQDXGgg
:D#3-W?7SOeSO(<@T+dS?0:-4+)=(b7G;>Ub&>Rcf.,6;W+e3&R8D2[+(8W<FgSW
LgB?f+NOcEL9IZ#&D3]S,S-5?ecJJ4fc/@EddHEc;>JIgG/0&^F#RcB@9E)N:U.Q
[]Dg[DYReT63baA6<<)8Y)NQ73APN3X/9B-DW[ReRMUIf8<KL]IdH>=_)37RYS<\
WAW8QBYDV\a-\cOUQU3V](d&@C+_EJ4^T_4)W_>.A>07\8?,aHLG(f:_B5U#6C0T
N?+Oa-eP+1S93GZC[?D6Gf>g50^3:,Z4@<0bPPLGKc]d[D/VJJRfW1f_AB3+&O:]
bH6SeaS>1Q-=<39ARO:1FRH=<c5I@#1XQ?X-V<5;5##B:^QHU&cMX\4=]M4c\Oe?
GM\CG+S]#dWcgJ&Y(<G+90UE6c55YNfD:+eTF0H7\W3&Ue=BeP+2gc+H6^M0)0E6
gfcb[Z.PMJ?XP.BK>.(Y>L/gWag;Q1D^\CXe9VN@f<MJT4BQ&ZgS3Y:#eSLUg[.0
CfV)(bQF@2_;^WC\U@\=YJ0U6O/)H@&4?]@_BXJ.Y3\g[DZ[U\3<RVe8^F@8Y9b5
JH0A@DC>Ad;Igg)\GFD)GO=@\13TWE\)<F&S7&&22YN#YSbG+ZQg0&X_f8eDbKF(
cI=aASbFe=&V,:2,<]YRV:Q>#25I7/b#Je<XE\/EDK;+/T/OMNQd5@MPI(0UO@b9
,;TM3N&;(U;?56/bLU8I/eH2F0+a8_f+\-#H9E=)O;&aRQ6YS.Q#R\I)g>c@GAD[
.5JfMAU=A#6/WYY_3+A<#a[<R8G\ZQKMHI(LTgZMH\58;(A8]^@:AHM\XJN,):Zb
BL^c1\=IXUAO9Y,M<51?-M<-PBOcKHVW?NW/4QG+_>#86=GK.5_VM79RfER?)b5-
3_>D-=)-&XO;Q3H+1\Te811+\MEaJS)H>98RPbgc-eN?(]J&/7D_6H_I7_@I0gM[
g^EZ+6S[CVC^3YbAH40^LD12S4>.dOUPH/cM:+[,NP,NcTX^NeCQT)U[7(82B6V^
;+?4fgcE^e:/2P1J3e0L#U4ZdGe+V@VX2::K+]?G9.5CSbDLUUdO0EGE]D.D0YAY
E/0H^^<3e9L4<f^IGQR58f/3N8[,@DcQBT3/[b&eD5N8;0-D1AdR/#L(G=5\-R.;
GCSNRJ;(>IRHN3:Q1PQX0g(Mg0W4SRGL60=QgecM&aDDV[c7TEd6.+(fH/015,C9
_TN47:ZW(#8D0)^efTCW)E6@cE]=R,]2MAB[2:(8)>=]/TS^3fBL3/b+IeNFb]J\
EXPKKa5N_/b4&:,DR/?BWOO.\2U>,G7+3Q#<d9@58H0(EQc1ff4F?\T\4:K56bEO
,;&-e0WXAfcIf7E@@>N]FBCBbE_@13TITYW<71R6W7DRDfPS[&D)E7Y32IYQd5N&
CB)g3S^AV(Rg&H_24)#[Fd=H(c=F,\)KFcT(de04gY-D2.g)XRb?+KL)59)dDWcV
JD@,NM._,.,(C;ScF[+JKI/RYFJOYDJbC;X.X@0H2U)7ME1U+WT:)A]?gSfe)=R=
6Z_R]5CJ31\D&-X0N)N6XU=cV[aA3US1/#-+Y5)@C8KE9VW]NZ#E[6?7NKAY2;bH
BdH\)J<.g6@MI)XX#>d/9V1X7&+]TM9\:5S0dGPOYJ.8BIQFFPX#-I/6P<5#4JH,
&DY25Jd@3_]&[1XYB>?.B5TZ[G?0Mc<3IMN9ZIW@D]U6#,I;[N3g)OK569b7b9?J
MG=VQS(S_7&D2A/bScBT=#8HeB[=D/(&6gR6Za^4EJRc#EP5Q9,1BQK=X<ddRFO,
Gadg6f3/3]OS2X9-E,(-(Pd[?\_/bR)\U:Ud:^9d_4\4&)eLH3A4NYET;ZYCOG,c
G=V0)T)9MIQKbL(=(>cJS>;13#+9D76K5Q>W(KZ35:_AaF(Gd<[6_04SHTLLYEF&
b0ALCE?acXfI<BWJD(HGCZ</UVJ(1MV0GQMPcZF8@F]1KSEQWb(OLQ1-](?/\2TD
7;1I>#2X)]1O0d4K.A+).-ZZEQU^[I.eaL+=5\)YEITW9(VSe+OGGF+(TAZ-0,9I
.dVONAV+MO6:cBFONS.U+7b#(T0g\JeFA:IS/(WZa^^3R:P(f@U8V>Yc<IgGS2YN
GECKNNd3&f2J;:[2#d\P8(6/.;[I&-cDE4;08c?>[6EJBQVIa6dARcd<_GNX-?QL
Y[Nd,<Cc\@c-6W2@F+1P-Y]^V64S?V>g/(NMBGf#NA9;LWC,OZ;]7d8YbK)T-4K6
YR?762GP,^NKNARR]8SQW_eG/c;Rff;&)VB0\Q6Q7QJW16e0_c2VZ3\2K.Z\4&6F
dF0)RUZ=dJeTd_+M.f@5N,O>d+)fb<S\d_:QVGE+#/GcV/,M110[d?Y67&&/PG54
_-I5E<]/7\.SI0+XI8>TWc@DDI-Sdc+3L[C<#>\23-_;O2cWK[>WbAO=U>)#KB7#
?b\NUVLG?E+B[;A<&O3>VVB\O,:5LICcaO#FO]XD/W6X0&R#J(8EHZ:\g]I30ZV&
0,:T+V-2&^;0>FSd1)<RF322^ecR=.8Gg(dIYN0dSYC&Q6GfPA^X,YX@_aWb&Md=
IF0eY0?+=1J+Q;c(2#3bL:HYTRI:F0KZWaF5-RgXPSZ9;f)S_ec:\b\M\ZOD@>)H
T;A\X?;2e=H6\gPAbHM@gHgZ-\.Q/AZM_OH4[\e&BE&Pa^?d;C)6V4@/:@>ZOa9W
.-ZWZ<0KaN)=UI[<Saf^+X5MX^c7H+b>N9A26:PCZVeK_3U?Q91WUX;-9O;E5b:@
6?aLT-F=&d&V]H^1]\2b7d)W0eZdZ#1TIJEY2@56NMDZe[VO5#/4^8d+>[)AG0GW
O;+f<>^9=AMH>#[(:B+[^8S7+#FE&M)caNUH(.BGW+28\H&aC,a]ZL-ac(ec#6<6
+K;)+?EeW=-:5g(BTQQDIH(4Sc@OSe?[.5+HR0aN2;M8?SEQT,+BM;[BP:?2)@g_
b9.[BPSC;6\GV=.^7.6#1M\0;4b;Df.G6TTLS8H5MPaJ/>4BD]NQ@O<(UQ>N+@96
C?g,#@VSFS^Ha5A)LEQ-HUU>1)OK?JB_I&/#WPC60J.O2RX[-J&G>SO4b2,b(IX\
Q22&5O7g<@\)[.B0eC/9#=.9Q0-J3,DLHdY_)6:Y/R^>.:<X>^T?UG.5-ggZ1V;(
HG:Y_H07NW^f]0gQD36,^TSbNC(+._^(dfC(YKZ#OEULM8I=2QP>Xe/.Y0RCJ@\_
FE]G[_&Odeg(TY9_)P(6Z.<(bg3bcHC;+BMfacS&ANPA9R_@G0]Q2C5IORXe=5+\
bd15;HP1YJ2?_2d@FMT-,;=3bNeEgCYHVS4(++SF?f8Y(cR=gZ8Z:OV^3DPK3,CZ
>f77Y=U:2,J1ZN4fLUdF2Wa@T/6;[?LE&a-6PMFY/7XD(&DS&R<R.]=.>&;^,^(K
O]Wd_K10?f<S_XH.#A]:ARTG))eb<U8G2>377\]3EHE\YAUYMB/UIcTZZ8@fFdKA
IA:3V1VAD[FB=_+[J2fZeE@TJD1DE&-^L4RHcbcJN@SIWW/a8I=-a;c40UeNb[/(
Ac2;]O,eIWYgQ&Q\6LK\aGdaI7VM1Sg:]+?Y0E>W@GUa-&D\0TfXEHeCF8ReN[I-
+]4#Ga.:C8)J)bd/<:B2/cY7X>:L0Y@RNGZS(-QbRPZ7,U5HGd6^2Y<:4TR+B/4>
/2U1W8DHG[V8]ZF7=.B2IfRRBVTY48D[G-)NZ\QN?(N(R-0DS>;IQUT[871/F-)=
UIFaS\&_JIGg3U[CD=Z1[RY7(572SD1g+U)?8/,T_#=E3Jg<(I8\:N?\Yb;I>_@3
c#f@W77G@[9Za8V6VKG^c^<>B?5<,Og,d0.TIONAIGJV;cIM3KgV/]^_._B_ZIUR
:&0RR3>BLSS-Q?HF/C(N00CL3R52Y]+/.DGPKLTJObMPc_+YY/08Q;JY(<>FU;Bf
;U9=@=Ag[Z5PaHNa727&ZM;PRTL^Eg2P1NJgMQ4Y)C_JcIgI/ZFZ/=<>9TGZ5]&F
@]9?MVeWe<O/B?#U()=C7D_DTN@Lf(X[[,T^eUIe2>E^?34Eb2OT,[31KP)[g:J]
5N.\CK#ZUTb&4:+K+1aX/^1)I?=(8.=T,P<NJgST3#aEO?(LPWC[eXM;_e&a@aY#
R@J[EH)I/J3RN)3-DDZ=.PRS[E0)PA8F/S0[?gG)]C:2,;BSOV#GJZ/,0<1K+&NU
)VH,,/=TD\d,JK39XgT>]SZ#,>>[G>F9F&@],GSLG<?^.A+HL3b0aVB.gMbE#M]W
[D=#S2PLDE4gX^cYfC_<9E#c34gD,^E&7VRT+XXAe/>DNE+X-K7OE@U.790<S&Z8
K;&8(L-YS?)3f^,4Zaa=1-W\[ddgB+2,#751_1.^^N-M85SeDSC_7IE9_W2@OdO0
O/GWZWGYNL&U[A3V4Hc5_B7Dg2=]cQ[UK0b90PPAba15=##HeRJ.f@@-dJ,L9&U:
Y5>I5].[-M<3dV#[;+KHY[H&G&BL5.5L:-,U.HI:][CPMWfD6[)&JSPX8X)S7I5R
R_(1>9H19&gQ=,_=DG?B/DB8ES(LAHCPMJ.bZ/;W)8I;RYIMM._?KV_(\7bH_JTc
:4KeDTTJS8N<8?TYQZB/]7N)3(I4C.UP@)a4\,M0O>YDJ2:\:PEK(6VA(=>?c;9E
CVA+LOG2=:?41<,.CaU_EKL5SbG:G,LHg,TUZ0199Z-[Vd[aa8g83c^eDZHLYf[^
0&1?AZTeM+68Z>4H&Sf6>/B3C/AOI_eCBK9M)L>NDTCX]Q#G@C)EZ::EXZdM)W:g
\K+dCHC23M9Q&=NSHf\V&DL;.Z3R_9#OH_A:AHK/?J.5Z1)N03BQPbJAOf;/9,Cg
)5VTIAaOM57Q6V5Xd1/\5&^3WK[FX>QIIc>(dC0P3J0-ES3&g[aCKMfK-K1AG(e3
S?K+fDYOMQcRa.ZYW,&EXVG]-L/JQ?;=4#=VHI<5/AgW6N<H\&5Q<.0V3HOAWABE
NYLHH0P3S9e1HZF+8ASaAfR]AKNfPW.@<caH>b^Q2SLf;4(5.KgN>gT/c)AD&<W,
2<#42O9_e<EDL?cEEd9@D?F2dP[f&U_G6-XVGYSYeffOaY.A/gC6XXK)QbS&/H(J
5B5,CfAMSdbT#a,)Sb_/)B<SG,<X8Q-@]S+IN+g1a)SQ/3,.&F_E]2X(=3IPRCB2
[S1<ZR.AEYX7gbd\8O0EgH)EYD642&;(P2.HA:\ab=;3&43;0WV>:V8EX43CEEb\
YbEI(.)gPFMO,EV4A73dP(NC8DZga/_bC<f5O(RU5_>A,F(1695P[G28+_?(8Y,&
<#;gSVJFW9_UPR7WQ3HDQK-dG[-[X(6/X@S:WbIC_>cX#IX2dFLKW-@(YPYJD#.e
2aM9F_)(^V\#TgZ;g^>:Md04&0]V6]M>W?Y\XJON;Te6)Y/?635X,[R#aXS?TWc0
CBDg9DOF17)7.JI_cH#6?a.QR?)=9NTgY?.;L8N\YWSY[S<2IU[0PP@8Te_cH-&c
a&#V1)SRf:L1#QT:KUOC;2,]YXEA7M/b7IA\RN/W>7@>TT;a#=V8PH<#+55NZ.<E
[PTK2gS<Y;J+bP5cIK6_cLc1_A,_&,_OUBLFMSRb7KYW/0O>9.8])K(b3,LPA+&]
=7605Cc7/J>9C\9cW//B<BD#GINcX+?V8gHSE[Fc:/6OMKMZO\AZAb?Af+Q^]4]7
9+&4@GXM?e-]Oa07dM<gFWBJX4WT.#@JR8PE,XWW1SgM[4:bd0gEM3)=4]fT15ba
793Rd^M6XKPe)(<+23I?:]#N(Q2O2\Q&#8-RQZW6QX098VM3)#59b>/T\[Q?0.T:
U^/^,=30.Ab]]4#f9/#>+5E)YZV#>_.c=-A/0cRD2J85A1O^ZA?eJWABH\4:9gb]
6(/H:4E:LGS06]O>ANM(FWL5S]YA9(WEff3P;IFV4;04e.3HX1D_:/OagCOIA)D0
>X<Y(0G;>MQ][RKd9W>gZ:S8IE>851Pc6FYaJ&=BfMMC+>aYWHCCSFA+>;UZ_-6+
E/f-XZ>La(;3/8PSQ.S=8H<gP(2bNY&2^MLe<07.Q+P,[:eC],@0O)<F0Lbg5fb\
_<dWf9?6^b<]-=[QK^N&(T>g]KaB?WM^\UUGE6I76]W)&^d\[CW\&8I>0&cZPF3H
\ICCT3Y\JVQ\1-^-(D;\6RD^Ld(H)Z:AW]#T4_P.8L#60ZT]ROOWde2HF&.+Ic8<
S?GNGZfEP]#=KY&5O@cT61d?fg^>bD.2C39W3Y,RX];c+a-(\:<PL/.53bL#0E^b
HJY7fNNb2FT#:SC13]W#UEbS4R<(4SB9bGG[,I]YDOE>TD^3GU=)M.&((]+/I:f\
XS_WJ(7dK^U\RZ@2fd0HWKQ^Lf07>0Qd&G,S8T5IIG#UVM7]6O)&=f.:S;4;N;AU
+V2O_0+@>^F4\;S334\7]=)#7#CBB-Kd=&1dcK,/>2e>G77JL]TL#\d8WP.M^)&F
]?5@;<.#Ac+EEG0^WPA#EH\_+.^)4C6ZI1U=)42KO\-VV]\][?(]?BT5;,EX#W)c
92[]#QR3^L[LK:9Vg4+I<c.\dQaae)5d(>R^P&QV151:),g,RI+9IKAA:dPDM+#P
=e93JMKP&KbI),AG5).0)&22IU_]F2SQ&V+^egSe&N,J^UT-:Z:M3I:WIFGg.P._
Xgg@/N.]NC2-PNX]4#-W5J9QI[<QGZ(0dc]@16?/D?DXIT?([@1B@103GUN@)<UG
Q2(AHMO,2?f)S71,2G_M-AI?\Z3/:MUT\c\,D4(Pg4&@f>)C-[CR;4HE[8,-8TQ-
S(;[O#bf_J-A@;XN0EF([DI586J[/dTLM@]T@SZc:f8(-;:ebYEQ/[M4M+>D:CH6
A3/b;XG0<_>4&ZU48dE-J1\f0a(OW7F:^)AbF-L3#IbYLL0UMX1UGBMXfGWe#&RH
<S3^JOW(OJWV3d2O#F?GKg5T^0M7:[UT[_::eE><Dabb+HWB@;@PUGPHb:WJDV&d
G0/0SGE,QD;W/\<IaS6F3G^M=V/A4(-K0D/,/Y8C8GF9_5H6GK_9U2&(^GO?a0LI
@KU2AP<He)aMX\C5WE@b_BAKg(0FIMWX]=.C@#6)XA3(KJ7cPYYW-.\8)bBJI@8D
D57+9JM=.MV2<;N6S=>GeQd<M++[GBOB,)2HcC>(>.ae9.b\P/V+8/Pd7g0/g?P4
KPT^Zf[7:9F_CQBGEE^Q?CJ&[F.>VOb<?3_F/T3M)d\ZAQ5e90g2<JeH1g\R_W;6
::VD6X>50FN_/5S<C@VUQGOX]H+49)B\BN6^Ic&GdBQb9.IOb?e>,N9.2\@B[C\\
;-)W&,#=MH2P;6)(&L@C:8K-eIX:>.#?Z&M^L@B.LI)MT1>T=7bMQ3_10J\SbS=a
Z]SGeYb71(7RG=H(/f:O@,XdH?U3<OI,S0,@FPSNAB^;#T]6BFD>-?7R77VV+cS_
94c\QeJP18I#gWB@L]R(DNbH0BZ5C1.OYV</K_Xd2/J3:JHS:5Z8-K=(-.a:58T3
aEZZX_V<;B)g;FQJ+-?V&?>\KW-0R@>S2)QXFR5.8JEa_@3Pgb=A98/XDU#aT</@
b/,Da&J-eXXE@VL&7L?)JV/3=[\8TV0+?E7B4ARdWA^Y]S)G1H;,gPG7ZSZ>fT+0
V+]:,F0E#X[,b&^/4ec]?URaY@KW^d6JK><Y5<UG=;(D<8X0KY8f6U+-+N75Q1H@
)E9APEHe0I#9?MY@#Z+/YQeBCS]/aD@E+P_d:X=92LBZg5?/<.>VFQRZ]4^X5Gd-
Pga[A5fU<2=YNXJIHQ.E40/P>>BWFJ.a+GYQ;46Bd65&ZJ,)W0V\E,Q(I.W4E;@J
Pc>>fV(R/cCAX^[Hc80X\8&]2S5:N[I/U/+X4E&RX[US9OC<Z1)Xa@6QB2[+AV)Z
?.Y[@.]UW5VNMMD^&+;OGOQ9a\5F]L;R8[TT)SRVD8=&7F6GCH-B?<0a>XJKF2d>
:_.Ya\SSFU-#da53DT=1T3Y&af)CMAICT+##aXZ)2J(^f/VaNKgE(#L>)c;b_6?,
YZf^N\,>A6ZHY?+GYG@+V16A&<KW<g9F6\M4IUJ#R&54C.]&J:D]62#O)<ED@=FI
NaKBO_EV_@AdCGVHg(gX-X316BD?9W[cOfH>g6:->@-SdE#bLCY>:aVYNEGM5dO(
5D68Ge:_K@EC_Va/\S]9?-X[HeKD_(TZFHSNC.[ggTf@Lcf>e_S6B1R+M&48K+6-
a5HMZQ??R8FKEYdUI#OaY7N^5NSa>LB>[)cUA9OMa-I_<d\318d:5cMSaNA2IQG;
ZM2_TU^c&_254_>&ga,NS\F[+G#S+1ILP(5dL@(&+bZ/1YO@[gI/TAGPC+dT-EGg
26,VZ>C#]LRM\L3S?a_J0IK@6@2?5L>R<d>LO)&f^_S9YHY(e:0PRZI_B;Q^ebZ(
81c[dg8)N]0DDG@f74HB73Y;K0<MLYN.0A/;T-1>51]VePJV&4D8/]\WKFOFF#TL
<@d\2:W,)gXge?O^A99236FGV,SD[>.e=dd5ZK>d>_[T,BfO:aFR_4[,6[F9LL\;
;,8TY:IX#Y>+J&4aM:=)6f;Y25bX1(PY6c,MgEfcaGM[Eg7IT.UUPSe:BA<Z1;O7
\@RK4X-:JVA]a4XK6EF(aCB+M?W[1?ZN&^XF?Y]_g.C5>aOa,-XFK;15=T?We=Lf
ITWR[ODQZeY\F5=--C>d7O<E7?0V?,bNd]g##G;b,MNX[K5;Je<BR,QeM>MJ[\#)
BZZ34[UDOE)DR-4bEaA[BYYQ-Eg(IgS-7fJ<[_[C=d&fB]4a5ccQ>Wf&=[.T:cL,
)H&5C@9HFe]AZ&fUX+ABL.\>ZdCSTFf@)&EG.fFZA/9/-X_;.](gH=K?=f2T0;YD
bV_2=V,+TI3ZfK):^I,V@O8HdK(G8S#EQ(cYE.]XZ6@0eJ#Q,BbBL&1e,Wb/S;_0
c-;V-P=D>)<GORLD.dB5/Y42RZT=)Vg5?P>T<a)80ILIbbMZM\#J<[5-CSR1DFP.
GT]+TXN[TAJ>_0I8S1KMC3E4)f8,b7LJHNQNZbG/3OFXHFY;2QWAV]6<PHgJefbK
\K>:>W3/HHIED<):fYcS\a7J+;AaM;07b1<<a&PQDH?CfUg;C>JPX.:/#T,98U3,
f\L6DX+Q2L\9;VB@M6AFT_>T^A2=V[a2/4E(A.dX2W^#.0?^&:OH]^P7F>OFV&L=
@/^>Y8AO=4J-1_OPW.gM1&Ma8B_ZeZI[g_G7CJ1P(<X9_-9F3AHC^Pb4cbE&gNeS
I)eY1=PLO#2=MX6gFf865f_[+8>6c>Sd?+@][TE\[V)YKGaVCPKE/&=I/dM_-HZ#
;UZ:e7NU(T65Z4V\61N##g\aADK>SF07_7::+B\-0][+7CEKH1?27bc\^?g,;=G#
(f>6c2:BZQRRe&_?PS4=Gdc/4:g/=0WJS2(S\_612d0=L\N:+^2:PKYJd;9Z]Y2@
VPEf)XI,9;9K<D0U@37_D[Zd1TfXP#[[6?Bf.A2(EZeRK?fBWK06GGC^8g1:,U6[
+#e^;-5GWX9.L2eREO4IB:dNY#IVK[S54b.Kac5M>0]_K6a?e_G-B8,CI(JW&&O#
X\AO/:-,0]d.#9@5T<1JVQ(^aPc#C#T/&G,Qc;L;II9-<:(,0R8WQc/g,=U/E^JR
/Kd:SM>178346YUfM:GaC:C-T?4M)fLM4,fYY7\-53>EFO;U3#G][,<\?A;U9#6+
_,GW&WF.=U#WEIga49&Bc_a\[D9&2IFbY6G2Of/3,]gR=]/>2:O7HdA0_FY4)g8a
+Y/Z>VI+X2/ESA)K#8aFOL]8(#F8R\[5DM0P+R.TRaRdV=1KV6eES:ZC:D-NM0=[
G\K+?9(TE.Q3f#241LR=GcA\G(#BIMQ[.R75:)H]e>P)f_P#0+,e/V085PG>-PDZ
?gcWXd4)>b_^d_1C/QT)R;[DTUC:QgI:LbLcR\,/V[ND#c5R[Z84@_(P1I-PRYSD
0](G^,DEM=<T[8[bb384IeQ]59+F;;8YOUO.@.WAU(Af>7Vg6a-CdSRD,HMgd&I]
\&#@T=L[Ac+3T&L9Jc2_.Sg)D4[8P)7.TFX(=P@JJ[a:a]&TE_OP]YH</1LA8P3=
IJ4MfcN3D[VQebTF=UN[2W(187OG5TJUdWSbZCFb\L0)d.TW@D,YY6H3d\?McIMg
CD/H[Qb3.TeR43H-1;/,1IE+QNB:^RL.@S6S]gZPF0<4e09^eP@1?DMWEL,>J?NA
M,12P4N7U?88C@W=P^<cLB1[?c;5HB^NIT&NKc?T[(V9g-;863@3W03c8/0=NDO4
c^3Fc753:91@AJ(aJE>7-D(#d&a@P+<,#E,H[0LGW[EG3<_f>#JEQ+U_[/AO9]KD
IIKXC3[32@XEMB>L13NRWCSU85^IAQUESQ78-GcagRE1I6^F7ZgU6\@S:N;.N0-U
MFZ4d=K(F.O.UaJO^aTP#D>3=GeHJ@#bN77^17U1eKg=5&dYQcBB5eAQVb,T&=CA
26]c=V@V=8[J0Y2Af]9T;J=OaR?A(VV+M?EIPD7(\SW.7SU[\46WY-,@@R^=f1/4
[K/@G()7?,e:X\]KDaY-DB/aN1:\cf-W+M^/M1#VE:J@M.d(<A)c>e-/XB+[DT1c
-g4CFZ(g+)bKE<afc@5T1TOX\L=;HJ>+=D)_IU9K&=HK@3<1f63:->[e32?\3D?N
<E(>^#(R0+5A5>BOZ8+-,7Q[6cg6QUKO&FW0KU.&JecB68>]7&Rf]@[S\?SAO;=>
MY/I)K4S7GZ6)MX-+_9OeS@XEU3b.f\V]U=0H;W8^7Q;6YZgIW\@@I]@Jb,#:5Z6
#.34bWK:0D-4IU[ND3=Z(J@-5B_):/JRfY(ZWb^#8_<7<Z()PaF8EV.7_8b[Tfe3
2OAAR7a<.7T/E;CY7BID@g;)3Y2Y:a22NNQc3D=5_-4Jd0:.:FYUJ(=54/T?.(Ae
X7O.+b9[faa_LWgI;B3RW6AAR/8@gUBHSZC[89+G]./RJaC-Oa7X#;JX+2;]Y2FW
7DIYdH\:_+4[[KOQ/\1#-JD5XF:WB.+W(:^<M56ZRf&5)NM69^0f#(XQdP+,.e/.
g23&O<cT5T>CF[b,:KEaD-HBRO2:R_K\XZQ&:YW>F2aMQ)][V]9g0/C=0&_]e1-(
O5Y]b9BLHEOaVf>@=3;9J/aSCE(87+b+aWY]Z&PAd9\GRB?OUCDW188U(I5C<8I8
BcPeDD]()02D0:OIgI?723CdOEc<AI#?787;AB-=FReGgRP+#RUCQf0+G>K6Yg8>
+V)GRB_OVAJ[a4_=?>,>INa(JE=7bX0LeXHe8f^@T^U+OU_#-G,@5RdTf/9bfH22
1)XZ=B/I.d[W#JQ3C28f\?G#WDD0Z-5Hb(3QNBMV@S@bX[SHY+[0J:VZM;]#_T4U
W<6aR@ZYL/SOf?;Q,#Uf5T^]F)<U/bKW=(:?.1YF:eRLa@5/dDZ^GV9cRQ]O_P_e
K,AD:17N:-d.R]@Wb(gOY>Qg]0#<fE)55f=G?K)0PAEOY-f[c?:BbM(e/NIa=@5@
1+G>[067=NG<]c,(,>f/#e)@G/g-E1</aG8LLE^:^:_(+4&>ba&a?,).LZAV(b0#
O;7D;RVcIKEP_9aU\5GQ2/VYa[[F0]b01BE+46[#Q:[eLHZE5_KP5:8fJ)CCUJ7a
PR8WPcVag+V^5CA#0,E@L?,fGE>>W)/0[e-VZ(CUa,XJ)-E>-^+V84/O+E9ML_I@
5+?eB)e=)\G.)WWZT,10KVGe&e1BK=2f&?U&1]+8NG-dTJ&dOK&X_(Y-;\976=>E
eQZ5>>Y,8BW@^@#3U^4,H8;)e^#H2NK<L]6&]=BZU)I]aTAQP9+H-P7gXg59S7+O
UQOG7(3EVE9(R008SS7[7UY.AbKIAD#SdZ5?Ag<\<[#X_UaNN]2406fHHZE_FK&c
K;^-))DX,IJR1g;(X#JZZ/VDC?\W7ZIS4^LCJKO_D@T>P9@HfUB^_b>,#@-e,fDV
]=,e<+=eTU,VEffV@HX@V1HHBC?@E/C=dSX-BVdZ<,<LFb@Z?-dF<F0&.L]g1=fZ
?0[;WUOJH,B1KbFbJZ/,WN5V#(FCQ=IcBDZTceCd?4(0DJ->cN-89,ZJbDT0^a/:
XN6FJb5/dHE^H3G:T#e#K-=WUBfBa5#E?&UC5>9\,<Cg.3E[U\D?6L&OTZZG?[\^
(Y+,BGK^9\33>3<)XSJ,AcQ)5BWed@D?1?:5??(K12+)\4,MDbe-J8;LUg;G[<].
NF>5L&RdQKI9H?NRd0EFd9>BeVVGMRc64Jf\QJ0TU4:c2;K:eRK4VNae7R/ZRa/X
K?#B?/T+@a-^)Q@Q]WRG)VC[bH,^:_e-]/d)?TZ](VYe]238FdGPe]2_C54I^5NL
N&PF]Q77<T]V\CXdDF(b=S5V3\@ece.-Z-HK2McUZIWYQ3dgQUSR4C+J])c=_AQA
>774eI8J/E<D<W92[DZX-RU;eWPU>_THTg>3>aIN).\DPF(YXK6dX7bJ@GRW&ED)
?,Z+]?SJYN]JJMT-8R/Vf>.#Cf5GQKZ-6,KXBe@Wa.EN#cY9UK+5,DMR+b9?LIV6
LLA8)=)/b)JY/dP_A]J#+B/PGT64SZeVb\S&:I>)(JB&a]b=SK/)3FN)VYSX/=Kf
\dN5D;/GI.>a;+J2XQ(FcQgH)ZL#HW:L\<=YT)0C.8g0_&.,8N(,Je:H,fA#(X9L
Bg&):KWLNO9=OP:Qa5\G_WUT7:Gdca+RY;;KC?5<LGP]B(c3+Beg>JHW_@&P0YC^
a<8OQ#DDH_3LA-5B?L3>S&#.g?6R@<eJ)RFOE5ZY;#?Qg]G<J5RTN+7C&@fOP&g)
V#FZR6)2c<GW^0e91a))61=10PIYN;ZFQ\W5QM[7+W]H-MA-W2Q/4]UOWD_;,JAA
4)8-F@YE066L,b,V@9[[ETZT1\Z&6Q1IJN^4@Y-_TJMbCaJTbUfbBJ0N6<6NA1C:
,aPb0=L>U8EbZ]]9OD]IS5ETA]>ISD?_,H9MHGXYcJ,YV@YJ?Hf-aH.?PK_VU[g#
I2V[S_I]O;V&21-Fd?Zeb-+NeP/IFUM_AVgA7Z.e<LP,3VFAKUPQF1F,:A//A#@U
QKPS&5:7RM4@,.3KW5eKK8W-2E2>e5RD5,I9AC-0KcH/,WKY_5,a-d8.O0gR85cE
Z/65MIgN6gF&]X?^[G.XgLVYYSBe9Y7A\Ud#dB/5O\ee[.ZV\/1B:a=b4XgLa&KI
1[[fRZb#c1?UUF2C2^UKV.>NU=^/Yee1U[>>B#\KL[f=;YOC-,R/M/_aAf7/W5CB
c]F-Ca/.89R2afMXF<Q0C#H6L<#Y)_X>Q,0a2Q#ENCA.+8gN6cg3=PV-(9fKXD0f
XH=),_\fL@P&9N(#;=R/A\0WVQ42;NQN9UZ,2[ZTW:5EIMJ?9V9+T7J0>EI^Lg8X
Ve:5](6HUe[(5a+O^P95CKCI_OU:J_EC4eY_RH(LR;XV^YabW0]4R)NY0AOVaC;+
A41YE-KMOgWb#L3H:f,&OC-4[YMe9;ZJW@G[edR<SIJ+ZAe@>+_=4AK].LI@)WHd
eFLa^(Y2W5^:=be2RA,ZT,VG0f)[OP</?;&+/Y1c<&JVb[/3bW(^0#)(+[].^8/(
9T@D=E61Z,I7O:&b^&10E@(,UUUY]=0<-C&+Z>0;f35fB->W4HA?X93/VUXQ2GR@
H<G_/Z]g6.[ZX/Da^U#5#?/8=S65A3V;207-BU2,83^9T/9(aU]]_4E(+P6OJ)=A
fZ\?cL3UGFUH57@2bN9gR??fWc9e;P#S1/JZF<.MT)5=^/&#LF;?SP?T8PA=+Kf:
c-dg]?5M:I>OW0O&2@RA-(C\EO&HG)3&]W/^e++0_RD:D,L6@PECY[??bP3KaTO:
5T\LVXWET8Q7Ic<9,ID95aaM4f.ZG-PTM##(ZY-Bd4]B&Tc\0&J4XeEM<c:BXBR>
37e570J<a.6J^J:TJB.7Q,EE(66?7V4E6KS9[X^UYL9+01D=3(35Cf/APVJA3+b;
HW81=^?]d76W>^385F?OZZcAd#])(]@<T7\Y#O\W)ZPI3;8R-c)VZ/R,@2G5XDaK
W.3NA/dWGB)#P?JD0U-VVW..CV90_5&eLT4d)\DQ4[V0e_-@&f6dOB..gYAXEZ3d
.#8:?/V\?-H/SQd8HbAZOPbNNXc2SPJ=EK0H@M=#QeK9P/?G.W.dK3WJ:(6bPaUb
Z_+_2.,;g(E/cFaRY;=4S^Vg<)Dc[H^C3fLN)@5ZHVPG3CcDDN4VHV2:CJS#faL=
X?+Q3CU\P:@e\T1NcXFUR8aFUI&0A,P-+.Y,g-1PJ::Hg=(3+3(eA/0Y.U7H6eHG
BAV]1#eGeX#<S;+]F]PPP)IN545XYBN#OT/I0gL[aVG432.b&:_ZX3KC4^8QO7+1
<9Na1W8bL]OXIS]A.N+2]<HP]Y)9WU/W5?^J<SLT]9_(RM0)5e6G-6#]BcOQ6S)K
5@.0X-f0;1#[L4.UY<0e^Y-ZILG@#9ZO:2K#aJ><NeV0.7E@11XgcH[^KXJ9C^@6
KfV?X>d,3>D1L]<a[87M5^M(NcBaBW_C8=X&1Bb_J_9bE_AbWM<O)YM)a[=J06MQ
9Yd3]Y,)c7-_SNA4W9_5V8@G/18&7?W5BYcf<^]K\DHg760e0TGP2VK#bbb.5A\a
3IObI-&dG[/(Q#4]e7-10;0Za\AUV(2/A(L:b9M[-7)2,=MA\B@bE7+(>0.6KG-?
)53fW#5][(RTf4(2H@0C]=F_2fW,f43a@\>0aF:Y+4UMDWfZYX@a(L,e71).Dd^D
bI=)P4bG,GKT^\dUE?3#[g/,TEI2^M/WNHYM.38^Q9Z&+HE#4G1?^9Z;J:EEAXMX
-HK5.e>RNfXT,1C<-<0DD@e=XAZ?\T;/=[?=,P/[Ne860T-[#7,EWERYRfOL[0K3
U_E899>#B/3:7ZSH27PLB;8CIYGUe29[b9H=2-U-DAc8Tg.)F=[D+Cd5^U<UK=Nc
,3\6JJN,Pd4W+KQ3Cb20e\T[0:K6;O/^U(Jb#b3PL1H_,Qec\aQ<U(a(9fd/fT2U
].KP)gMD2&0E2DfdP]<UgY=HQIY=-[<^BdEFH:3e:]+/->b##?+aXc]AE4Zc5#Ea
B/L-g:]1c<JQM)N]>]].b-NT7A>Of:E7J+XHE[59HX<a;8::WHb9SOVL1d1&J];b
_QI2<=CgZeI.?;U1(L-IgEEOfAV&-;/RJQJPab0Lb\g#WTgeR+LT9D#cVA]F+WE4
.Re?UQH7aOA+E^SE&5NGbDc?BKdcf2F167fM>]EMBG^dL2Yd,<fYWS-gF^fB&@5M
[1&SUMPMLe(4UL/(0-_NE5#NYc0E-Wc;?;N[U>Z+@XJZ(.M[==X4#]<#Z_8:PE=-
VS6CQ6?O4GD:Z;4A2/UX5N)0X>JHe]A02^J88-BFSKS1e8Q8ddGY<Qg>9BX9E)8X
#I^<-WcZ#T1&3T]740@-Q=gTJg_#-UA0B<UQILLP9;+&,=)?E)d95WL.a8E@C77&
52&Lc1HNM2V<56^NRfa=M>G&ceGdK(<JgYII4PK&S178NRA<954<2S#\?W?e)W3V
IBLgU_NCOQ8+V^#AN8CS@YRZXVUb2.+J6YKR(7V.SN6E],F_Z,/dNS0W02RUBPGH
beWP))7QHG6N5:9RP_aa_,P/U:M?HfYO-79?aB[9A#09&4K6Nf6#7UMH9bAW[WKR
NXY5P6/T8VS[:UXP=_C7/+.#^e?01+XQ0OR&2ObHX,1-#ZK,]Y<-?=/VJ3(31(U\
..FSA<9;I8:Pfa8\012(79VKfQe/d:OgT4&.(PNV>_A32(BFWde:5g3\5EOY2MP#
MB?MV28V_DNYL/=V^d#_K36G\?M\ZR0Iga;E4c<M^J;.]PUc;RMObJ-8EME6E4G1
ZFZKM=2>6Q==DgRbA3J]F33;]LYaH4KB].-4XA1DT>c31Wa<AX7TMUYT4I:\Ra/#
8=4\FK-JSO3>@O=_KG\ZICcS;gLLZE9b#29aP8#6J0,eP(C..^ZFLZ<Pb((\\>4_
\\+aaQ4,a579;a6650J2C5dg=E#&XW,\dR>L7HD>ca8Q1c[-B_7O^RLYA0B\#:I6
#,O4SJ)F:4\6NaWO>19S:gD&KS0+M_E;5SCT@cHHW=W/>=d5LV<ATc\5X#E/4]\B
Ua1P:c4ZP?9I-KK3YD3.6eg]QT,&(ScdB7A<e4=[4960R_W01I/b6Xf1HbF;?9@H
V)bT:)cCH?79XbC\=[Qf0)b<#<L/A96U6EW=_Qe.7-;_MScFC_P/GdWXLgBUTBFW
R&BAH8e=V?CV;29@-g2OBNbd+6Q8+LW311&TW7VEWO&@VC:BW^\YXBVB;VS[YZQD
WTfENBKD&4T5=c?&+:H;UPf?)8Z#ZFPcN2d0T;Z,^Z=/TS0WG9#8+XXPd;DE;;\V
YR-DG8D&b]05[Ad6[fNX[bV<:f//eKGIJA+R;M=EQD\[Z#\Q)G0df>b4gBgGY;?R
2UJ<]L_3cWT1ZPWI?/6a2aK8=Jb]9C.](YK?fNdPTQ,7@Af&+I\eO@K^Y-V=_.6W
E0UO8B^#WK_f0XLXWN4,2LW6[[=X[SM)+ITXK+#3bOg.BD5=7BC8aB?)Oe:\1f(6
1J]R/;c:Ve:RL]ReD_3EQf_La\R6&Z>.5g.;BIQ+#OP;EGU/WfV\T#VPK_dAf55D
gNc6PAQdX82K(7VFD(1.gcVIJ9CA/A=c#=6:4bX9II?B4HE<0.d@g,T7\6#67f^L
#06/H[CaB7H74B\[O(\GUID;]82(1269C<c<\Y.UO>@0Z_XJfQOeC[&0=Q]3?\?7
d1@Ib@:2X-T,>(e-;@6L]20e@0V?gTP+D;gWd<@R_+>IXg&?2/b&9)&f[1O>f(GF
]9O][[?+gc7T[eb?aQF6VON?(f-/Zc7=5?]]WYA/Y]EIS6A[-Tg@I4=4OCL&;66=
I1S=KBQeafG=]P)F5:N9\\38MD2BZO.CK,+8VW)5<Wf]R:fMS&T7RFaVE]aR(^B5
V0O\_=-[6NS=11SRR/WKDD5:O+>I&AMEZ].1NIM@5G(-CU\_d:S\(Pb[9gS7UPG@
T3@(g:(8<T,7<;+@Q0bSFTaR5FcSW,NeOK.G\5X2UWg2JJ/D@CPFX.8/JUbb9/f:
#+H59/Sb3Hd]I,^C>)\?^6AQZ/8D/D,0+^@Z7F(JAM=B)6+S1?6Z]bc?;3[TeeN9
e5QQK>0+2:K7]#8DDT//&.+Zc^=.#N_&AIPR[58]BCVfVGBHM82gc3F([EZeS1TX
\W9Z[6H6f#P]<N2BQVNfQ1+G;YdE-@82?)3Y&Q3NC4A2bRFD>8IQX_H+6/d5T?cg
-c;JBg^6cZ.dcdebC;X_&?d>c3908^US6Q<@3CM;PSHEM_E]fZ.cEFMg;d90X4\,
WL^@NHMc[E&KDU,2GL[HIKLBJY2L\G25ceHZa^9GeV_=f9C[ND@fa@0.MJ858PAT
ZE3\_5>4E#Y^S>LCW_E;82/E@DHDARNMBI9CU7UDYdLT[b]&VXS_;;2GI]LR:];Z
.I@:c9+D(H+:D;K^;ZBJMU]Y297U=<,?O08(D6F]ACB.W3N,Ka(?(SHg-=GB0?ac
^JLD2@0BKQG^U^+PU3f_+MI/,17.8&8-YKb5d.Y;P2:SP;WI6b3J+6>)W1c(IC1Q
1@T#F^WTBWc,=f+cVUdP4_>(=EJ?81Gg]3Z..UMH#3JVa14&1P2EZe):B=1JCY[:
XI9b2&20^Z0>SPPWJ(X,7CYDQQ#EWRX\f0Y=E/He3S\:][\=F+=DZKMRH.?]X0GC
,N>N<_0,KW#56CW?1J0eM4G93T2&1)cd.g/[f9N.D_M_NPbH8IYf_XTU,RC.5+Ca
JKGd7Tf.@Q&HPfP)POF&]7TGOE##KMcJSD>ZJ0NORJN2W3K?gb-7_DLCeVbfK=Cb
F;eL3F^GMeO)=)d0Ac=?^#f6UCIXeeIAN0#\]BIcG#4U?W\;OA&b.aG+dKJD08[9
2ELMga=cY/f0I[)JA._,gL]geUAHW_?(f<&[^>Y[H+_bH^HLM\#&[4=U.@VB>Q;F
N,^dB]5<Q=N-2_IRO8544&[8IV>)QQ9_[8GHV/@KR_W6.FWE#G^V@[Y_MJ#U>NN0
;]VD>D1>PG61DZK76?H1,\Y]E^EP.+8(-QRP=GEW4eV+EOE,K=Z#7J+B=E>T#aB<
ZX6?\a-/L+RSVV#Q68;(4_O@A27d6<AY7->(][(c;S8fFU>\S;THWDOT(Q21=6[W
:D,^WFK295[LM3\eZObGgL(NU;;88U4#c>E@NU/,eaJ3ebgf,P1WCC4RFOCJXKF/
U2,XV?IOE\<2YC?&H>7YLP6>GW08E-a2V=Vb4,GI8[bfF)PaX]>R(X;9DW:]>b]B
FQJC49]OH?[[B>:.Q:8C?=/a=^bFC0/8a3+8UZ#T_J3U9I3AVI\BEZQa:+8U35([
<ZgQD5NYJQDZVT)&LLg3&1Ta\2g;VQ2<WJ/_8P3+@)#/)5T[4(&/@d9CJB-R5@<1
a<\gKc@=<g).TDMC08UBCI6UD865?Z^fP[P[V/.&ME>Z+B8@ZGf?Y\;gf\V)_LAd
UdNU#9NJc7L,BJf3R&ENB3G6?Yd(N[3D8Z[fFQ2)I9.]ga+4]-Jf6:+_BdX]:\IC
XTJH(&96[#[LO@VFf=NY-W097D4LBQG#TXAEdK(S\LO^JJOIaQ?#,MEQ\,1HG;Ld
7BJ7>SK?Z09,IgG#]H9J?Q2d@WJ0BW:?7&/DUH&1;(E.Dg0O9<fDfA>M>8?-/#)6
4a\FXYJ?=)Ee1U>E+VS7F6N>1F(G>/3R+T&D&3@9._36f71JI/+L9EJ7(]/CPL0e
XbZCbN^+..3N&T2KQ<&dEg>IbL9/8\]</GO:;aaea>MdN/JFIX]:LOD06a\4c4F_
.UKGYdS;_]UD)7F6P(;7Z7MeaDH-:V2:JIRcL?\8PM;+J^914V&/579B>_1Z_S^@
,bg^bU[_G8[QS5+EZ-\>ENX(P]59L#71F8WPaM;,VS]>+W+4@/#\UJZE(VP](#Wc
eZIXLCbKL4YVF):Fa4]Bcc[18IAS:F[IMeBTcQ1OR+d7FWdJ_5b7+6I>,QJa<&f6
@?GY#-4&aU\:YCVTJ.?DA@Sb>YH?\58RQ/OE9EcV(V=Cg(8J.E:_A4QHdX?Ec]K)
KU=9MMQ0>,[RLHI_8YfD#UI:d8GObgSZDcN)]\)H,CHGZaa3JV^NA)e\S2];<W<[
ZBeT85X,4?=4ff,c<@,0T3A6.7Q6L-\(D9&d4_f[8;\5&PU3=:2((K]I^DB>]NTd
.AX[cP78I?K7>bFMR60^S[dH2FE>KA[#CBS9g</gJBMLL^?RG9BKY?Q;-g4\9(T.
K+ecCaTPUI[4(PX46](]W-?ggGK_^+G@EC[GQ[K[gO<_OT2>QM&eg@MW:(+D-EM4
S;6\a=A3f8JOE<#H>Ha:2aGR>3=GSM.PGRa<XF^g]]W:J-ZB@_,Z]J5NM9T7FSU?
N7T;DbWB;Y#MIZTP[HAg0(&D5YCLO9:4-]P0RK9X0JO&Ma8G&JARWb]?R&g^bN2P
MYJNcFLE]:PMc;UOH7cH(+6V/0=JX[Zc[JH#&b5fQd&UZ4AN48-]CEK)XXD[PLD4
a1G<.9VTd:KF=A3cbB)7XeAKMBLVc:(#;dSE,WXbEH1FOfA,?=-G_Dd:V;^=P<BJ
<Y92W?W_V5&IUQFHA<(.IW4Q^#F3RPL]41g_MXfA)IaJfV9@C:1)g5Q6BNc22aH9
b[^].[Uf-D;(P6[FB.18QBfM\+9EbM8G^T&0^XPIBZYBRNa0a:+Bcd+,d5Q_(P+D
.--.MYJc=AZ/La^^7MN13@.[YdV5LSY2H)Tg_BIRO<U)TMFf:\4<a_dF7a;I721<
aGEccMJcRI)5;J53e.,6)b2B)#HFDG:AcS2>;R6/_+?4I,C6aSaFN8L?>#-8Le=^
49L/I3MW_>G7RHW\4)g^FKgCI.4.V/NXY3FHIGWfe[[^#@WWeC_>PNQ9?QacdbQ(
VLJ<E<GDN)&d=)A53[CH),U-bX2PP<<;dWV0&GC2&4eWJPJ>IfFebY/@#S9E.MF=
)JO.5\.>B/4,80=9M)=gG+^X,G??_&0b)^X&_15H3+QTTZ?Z0+f6Uc;L+I/]LZ2a
O5)/d__U(@\db4:DbaNWI4&1Y3<PBgAbgHS@BL:PeS1a>MS6/-NLeV5-TIC^PWW6
A2X1c&eC-9YZHUM[GJ?c6C:9F1F8+9AO)-+C3);WD[+TG9)DFNAXN9:?8H+;FPAG
YZFI3V@R4_SMR(^MSaD^_:4\^FDQ]Sf5dJD,FT;G6aH5g];aZg:.96LMTRG<8-Y)
(XG+#aZNgDCYRagK>>/)R0[OUd)MO)]M@D,.,=7?1#Q^6Tcg_44T5)/2),2TG;QK
LM^UXee>[>f8KYGb-;,4BZ&^PYaLQUP[>ZV+CHZC4NCHgfLX4?S52@9CT:>,)94-
0Q2N#ZB<B8[A0Vc:fFG_CH+:Qa5M-fR^I(f84.FN)=5[^61PI@fRfVRU:HJ&OTBO
d9I-)J,8NT9C,:fY(]O+U24\G:3.N,(U^1C\DT7F]Z^YCDG_e+5Tb36XaX?UR5^(
V<,:Kc\>-807H(YIb&aA:7/2G;E)Eg8eECTZ6LX@1CWR_.O@USHgU#I<[Z)F4H?\
-=+SSRXbCV=44\@+>ZT>T]UNb.eIf56+dP4ZbM,VV&8@f@()&=:Z4aPCH;6QAI/O
\C2G1[aGfAQ7DK&b71J(G=:TCJH@_KV\;C>X/1AKT(:-INY6NZ.PLEV4B@4ZN_@.
2TMM\,\-H)--21-OE:+3@+ENY<J9.WD]c/IG&5,VV2<9K\;JHOY[JTUWd;#/@Z4^
U&RV,8PKdAfBZ[DPR^V3MITad/R)YbADVUFV56VLXa)MA_a>0E):;=TL->:c&/2.
MdXK&B;#Q/QH;-(KOU1?f2Q_?&7UOcaZg2b:.BE_K+I2@aO+VZ>Z?GS\7^W4PRS=
FYH>P\Zf):O(FVYT&Z6;2;&X6ECdAANL^7K&,<KK/SI.?:8VZC:QA/)@7bI0X01?
;Q_7JJ5,#dQ46?\V[TE=(OE</_OfZWXEeL7Nb1.XKgIga9Z-dYP@M;>>T.MX(&4^
I+K6S[D2T^_GUD1E2TK2bg(g<aB0I#.;/)>]c/0D3I\D9S+:R7HF:+2g\>,+.gFZ
H)SS?eJR>5I_fgQG>\N(ZT]BE&5/B85\,ca7O:40)[M#c=SK6b.DSgbKcOQ-L6a<
/B<7;b[3>Neg+I4>K-FU5/U.&eL9@P0>fd10,dT(S8W5RDE+Bb#5/Pe<C=EcXVB@
8+LD0LGSf/f6<M:?J^HN@PN/=#0aNYAM;(@31#g)D)]53>,)1NX+-3Jc/H&9,]MJ
)Hb0[d^G5>CI8I/9<7QQXUETN[_d=N5:H-[?]OaG7YT)2-Jb:&WLUbK.8B.+XDK(
TI?+2?@V3-eJ?efX,KW<5GYgNEAHb22Fa-L_@HV^<-3=K1W)TLe)fIX0Ga;V6gJ<
)N^#cV])7DG714Z/52c0EQ_KdJ>D.Uf#GfZ(LV\7DVPF#b7_B,5a\<O^0QI\.CHC
A>65J?DWC8ec8J]XGa5eZMV3U^7N#FR,bS5?R-GJb[9<\UNAFOf07c5MN+KNY/&3
Sfe)0T6O8W8-?e+a@_9cEff_CXEgJEH??_f3]J_9QaRScVYDd:,N@SJ7AU2_(T8V
[eOK;Kf_1f4(5]#:F^K\ga+;((>Gdg3?O[BXO(Y7He^;[^4fOI)[FFAF@JH5IL.+
K@-DTY#PVP87502/eC31^X[&c]21G+H[#O<TcbK63eZ&Df;cPNWJ_/K(H&cdA#H^
4gN5XeA?(Le(#dAcCB-E@Q)Z_>DXP7S97=U>91,g1Gc_?.G<KA4D1?#/Z8/HL\S)
e8^^:#]UQ4)ZZIW2+PML=J9TI?WZ2;ULOQ.dQJ#UNU4:,_1[bMYE#-3d6,eRN(;4
)\TS[cI(>9@c07M+TD<(_R8Z(9YaQaHA3F:6X88J,CYB2OFS<5N/]Q.:GIE(aULZ
5R^]<++SM@#c5c?G\c&V,?2.FA\)bUU?#,3FfI95<@)#SFP_^8NYUK7M9OE3;(?=
e8)c8L3W^dQ8.S2+8/V>f5f6/PXPSIdb)]AZ+gKd38E[=S8CPY2_+@X3#VIW)-_D
Jg_4N3S2&N8]SWEV:^>1WEY;#Zf?CDF5P:#@X.,d-\AXU<?fW_(L3P=2da\_e])=
9P1:b66cF5\A_(YeS(>?VF0F#b74\OP7C+V/?T\#=<257AD(-]JI^KV>2H-N(AX?
34)KD?<Da^CY0aAYK/1C^[@OBT7.7(1ZYRI(?T2GWWff8Z_-NS9<GK+WYE5I8+E.
7J2aG^+LB=QeR4<LAdK]+D//N]4ZENK0JDT4_GfKD:Q(JcC4D2;79VYX>5>4D<1,
NA7UD..[c>_3CA:?+7BWa10gKKQH/M&1cHM-g)C@3/QQ>f^7^A?fdT,K<>Sf4Lad
1c;Z<5<cELPWR(:d(^RdQMf8[]D6R:,\SVF[VM)<g0),:;D]-F\g1AAM\5caaU5#
LCUYEGPB7d-T+^]RM&L(7=MC;W89?c<bG_H_.,>eRPS2MCfcL=K^N44ZMOB8EQIX
V//8^//Z3-W;@CR\R]f;5ZX#B77]OQZ.&Be\7+_P,GNK.+[>/^e:&cGUL3/U&:KG
FZF)Z2[=1W(?49Z39@?T<eRY2=UW5IC7PfRHdcG;^V:-35:,31IGKDTQ5)GIBBV[
Y:dB,a>=IGU5NC<^Gf=FZEA@aaP1&Q\;-(OS@ATQ&R(+N_H;?&Lf33a\ETbO.S+a
3?5+V/5&R,92d(D9GK\U8?a)=V7PQ;1WbR[Pb]G(J;<BA>g2,;/2YX-P<P1TF2NG
a<B4V1]T?X_XKd3<[3.V_Q@;MB)>14(d6Z7==,;GVaBF_?&Tf61eP&DM9[=QNYSE
X9+=C+#:MS9OT2Z;P&P9=c-[9VL5QNF]/T=]+D3XLOBX990e0WbM-(E7X;[X_[7e
G0Z/aTKZ_^[9:P[N(7LKZ-J3A3]<be6<6&;]BbQ0RSCT/6-gbA?eEd3;W7@W]E&8
Q/F\[CQXQMBE4I&^Qe@U4)_fQ_(Mb8[FTR\EJNMO(fa(KPK@-W-5?1@8C[KfGf,&
KIB,@T)2#_LZED>,18G#fC&#<_0IaDP/XU_>3E.NKSd.FcX91NN=)>FD>&8<#ERY
&#CEM/f=RVU3:F]2,S><(c9,gW4T#)Y_MHN\V<2=]K9UZ.@I+N<f:O6a1:=F7^X^
WC5;97HgYVHPJB,90<<Rc^L,Y=4K.C6B0R8AA;RMXR2^),PM&AOYXXb9-REUH,3W
-=6NK@Q[+#7CTW]B9#+XS#E):JV5Q:&geOa6>^M,ARgaMc?Q:-5EUNAZ4?Q--/9W
99:IAagC3YRF7)/^&)EeOeK0__f;bGf[0VV63PWFX<YBaGa9^gJ60faf0FcQf7J8
baCQ^^7Odg@\b4Xb4-2J9fXK4W/0,:R?6\N:KBc@]->#4Z;[GZ>YT-3b0<5U@6N6
c?R2@5.;N8g/>/A4VV-4B+O>2-aL/NGKSNU(cV84ee>3]=7f]P108a8_]6R>8HUK
Cf^CcAENM3b#QV6AV4_f/bQ?aT2.eNVdUSEfTH\P,8M87,:XfLGNf+SLK7<605<a
(A;a-YOA6.7c;:1fB?_B=XS5)E,+<(S&M9>ZX(-aB-4Jf&:^4bM+YLET,03LA1AD
:L2E0PeJ-POA=&V-T2QeW/0b-.YU7:O.HBgG2-?P;XV6L:PSN-ZaUJ&2F^J^C7e(
2c(LaW=GWUNADd@U8ITILX^)FAO5<7?0,IT?\G:Z7b.UMgK1GWR0]..25D5^8U)X
]VCIB,V\U.&1KE/HSeVZ()6Q@3Z@=>8YANgFZW_UR0c8]DOe_a((:aY_^6C)-:+^
.PBS6+2034EAgR33[&1F5B&;D5WES;.6Ce5><(_^IMESad9,/d,D)];\AgY/Z&Q_
L=]M^[Ne95DV+-0P4H^^:SX(FFA2QfHK(NSa9@?Af(F0d>>AP/I<PS<;PZ6=5Sb0
f31fZ[FH=W@34@FT6DW<(G:3O-PD-55bQGKC<&76#g()2PZBD-]=D&<7GH,^RE4F
^\\>_B<\C6fR2/&MDLT?N?=9F<C.IZ;GK[F.)M_0d28aSJS_)RG+GA\G.^FaPW6M
R;E6L,\HIA\E3.,?JVfNOC?@JaC+83B:d,UQQ\7V[bB6bM.5&fW(AfcU15<R1NL3
(&)eTVSC>QMKIJV(U:?S>L>Dddg76]X,AZZ97F9+,G>3(TLe;Z[FKE#,N&^0gD.)
\4-U&@RM;8VRQE=f1U+._Z.eacN7?+[9[,a(4C]Z#@[(9:A/;eVY\>McdF?6-c#E
OJ2g>fKgbf[@UB]bR+AC_PO]2T)]\9QNV^TUBT/EL&X:5=>/2\]9AUX]De_47>]X
BEgcbg\<ZX2cRd_W\8>f^3V^KLDg4L<]9WDV0]XfKJ[N:HH@#>_GKDFJdFI[,5Da
LgP,TcPW83=_?gD6K,W&^.SJ8;SZ1<eHfcM-1(/f:Z&9L[QN5&b+[LR:Q\P)XfAd
P-:_/gE&\2(<K#;,CAf;XZbc105\VT06DQeE;d.18C[8ae(4?[cAKKf:=J,C>IKH
HIEQQF:7@V2T<_ESCCLRQE<Y/L-)3W]:,Q;I2.f/N9:c7bF,GKCUGO812O0YGf^#
3,P=4U].Mb=a;3P.>Y[-/U1S2@PUWL.JCVN9@4_F.dB#:b7-eeZHA<J5/AOff-EX
L/(I<)g=ZFW:/47K>^R^/f)A^;22Q<3-?EJ7S?6E:S^S9H^KP:VUEG:1;@W=cf4a
T<W/(Z3W^:<1@4Z/O(>X+NQT?1d&\7P3bBgN8]ga@&RB[:dZ4&4/(U9Gd7Qe^<Cf
2XV3U+]7LccBO>K^d4O@7@66Y71b>5=Y/_2]c8D3=5W_S:#5V^LRRGPBb.O7HST;
>^BfHf,014a-^2P<FRJSR[Ab(BJ_X=G)XYea:=/OG3Cb-He\\Jg881[a)E6GXQe>
3\JY=D4SDb.A,5Ze+]341Q^c&HE<ad-N5Xe@8&@)+8=:Jg&C0@]/^Z<XBg\0:2e_
1.+,EUU^;3&O8K2B)M@Y33>H8d7e:8R<dE_c-bEL=CI(@,g/fZL=/R0ZDOZ5^1LA
^2G_9_0?M(f4IcGUNPI9=J@ecSM=gN_M#Z[/,(RFO8,?AG@KdP1dd0]W?_VT/,&+
[VVL9(d)#@PT6CNNZ76O2Ba/_<.Q)XGUWDM]RTMSCX<GeET2:[.;?dC)a2]HJ#,L
e9(Va03#5#46U@>APJ:?_BNcIV4g(:8?)Rc3NM_^XI,C9d_.^=EbBPPRS2;JcMDB
bB_52d-J0EKQ_NX^LHf:>\;ZgFUNZ4:^T3e(&ebQg?9CE2^@V.]fF)3-APa?P4?)
N(SUFE;VdT.c<d/Lg+TW^@CZE7:7QG8FJ#6_E,J\_f#1E?(])X6[7?5f<H,9UOY:
_SP]P7bI0+DZ#QQL+bX]XN)B]Hgc^0^0Y=)#IV>J7bdGDa45(JP,d]<OFf0/b(^?
NI.7)894RE]&G3G]fLBHG0&6)J46(X.aO_-3+aVD8Y_+[c7bf)<IGb2@BGFMNDQ1
7N8dCXW:aB/^YeR,V&?U^9N;8-:gA3&<67:3::[fDgP,BfA+b;S/++c:DKR[S;TI
7H#fJd&-aRZF9Ue3(YUAYdP#2/?fU8AK9\2M-b\ced&&\-Y5\GVY@Z1L8](V-05^
a_[D0(Z1aIVHVCcaJTM\EFcR^]KP,=CS+cH@0L4AD)QM+f8/14((4:S<9Va1PJ1=
)<4eOb[1M1;S^8Of>H)+4D2BL47+E3X74_6]GBQMH;GPbMg.1-HXGG+J7CB?IIYM
Ld(3O,(bS/TYSJQKCQ;V]O[XOf:a))EZJb)W76[M#ZT/8\L?.XcJ&Ua^51DWF+@#
8Xgg_]GDMO<==d+^Q<@V9_(2?3_f6cXRPNICTY.#.[1N_NLR.NCEc1:c5.G[gBV/
V^TZ^2[EFPOgcbb6AZL>2#:.N01GR;8DQQPgU0QQ+6AN9SM0.>/aRB5KAg&R]Xb5
/Kbb<e@2)LWE3)LIL#=UI5b6JUL?W9QOJe/8ZBY]-IX:YMUID@\R1<ZaJIc@TK:<
W9+^T)&;/Fd((6QADP,3@1<ZW19,aFXQ0a)FU;XdL;^#HIJISccUPL<LFe:UOZ7F
_+@b@XN(G3A-6WgJaYV^PKQYWZ(Y\L;8EVI<L&[df3/+N?[NZL>8/)>B5GS0b[]S
JBH)?U1U]VZC7a.bcT2HA+Z>WNF)QV:R7+fV6]7]\X\]bfJS75+>+IV^.S7&C1=X
&E)b[9D&VIVZ=P?PR_^8gO&.-#16RAO8a[(/1F71\].IWMK2LP.TP=W_EPLMZaOg
T=/^[c2L[^8?E&_a+-(dZU64:V(N4+MI?OA-#C+::M98bg#8>DSUJVIF?7:I2e7Q
IRP[MZ1K/[fcLL,[J?I>&U8(,b+a;UAg70XCCT),X;8,9aH=D+T1,:dPAd,W>=^X
U8a<5=421]^a0M?1E3+X^=+)M;fY2@P+WNdbC+SRG.U^gE59;PHO=XEe&4d\[,e-
\?8Occ.<2)5PG[RW-4LcM_88G:<9U)YF5&R^#G\G\X7a:RP6f\g(V:;38J8S81X@
C+,]?C)UA=d/ALI>)JK6)bC1@C2c^Q2KefTSJPE9CHg=^G/b/=JC&,;H26V+Q4KU
>#86;^O@MJ:B73:.2;E9IaR[KJ(CJ7gW6Wb^L;;#80:RCJf1K>H+U[[cb=]3L+.S
)2L<c+>F2Oa;R5]O6+cJS9@OF.RXM?6DeG==:G-]B[?R?)9J[2OL1B]RF9]CB+<e
4A?)F5Te_\@/AGQWW^Z;6^c/SXbG21\.L92JISe&IcH\4cPOCgH7AT@&9GSWZ+4[
P)IU55,:H^KL^Q.J,F>,I[2,/:O_P<HYLfM_ILK(Y#66U5@S\.YUMTGe0Y)R>N8+
<2/P6Z<FU0SLR+Q&->gVZLO0(=H:3/0<Ba5047:\V/a]eC;]cFWJ4dK:2H2<;58;
>2_D3(Ua7Rgc)@8&=5?E\UYC3>,#e[TS<Ke3N]&@,X+D.#MPRVRFNbW^&@4J29D8
LE?3fIM>SW14eIXb0>JAf)2-PP2]@G9NM\/T<XX)T_0U[,SUd6R_D(E,J\O@8-(L
?2W);W,a1Z07.aFMd4I<N8J9A67[([:c^O69W+??<]QT]?Xb@33)O8JOT](7HG3Z
=?83<c)VVf#TfXPc;..L;E0+7,g8N/LKY#4D<gM<7ab74S9M)3,;)d_I)ZD)HQE5
?:L)4]gHZ.0J&01bfF_CF9Y<YDe?OL,@^_Y?a@;@gS+-SaG3XNX4^\0Pd)S>cC(d
N5OP#>[&;JK#IJ>XH\a5;.K(R6BY_Vg.OL1fMX3?7fcQ;>7ZTX.MM8,N1XeO+Q]A
WL7\4;Q:HI(8MVGJG&BNgH&@RN:7-e7\AXLY5>0A)[gM2538OT\BE2IE;3@;FE-Y
<LN@].-Y^-DTgfL8]7WWJXJ_SU<]QOERcTXBQba,K,V]fSQQ(]\9Q?1e)X>[5A)S
\8?aAcb3UD1[O#M(_[3\bAFA)WR-6EDVMBDGPdT^YM)8QZ8AcUcU.b]d@b/VULe;
KC5eVE;3/^TTe^dY>cf<8fFPdVF.@,];4GQ&,,8Z=S,]6:WgQSGVWSbU1+RAX1)Y
9&OJH:E@6O:V>Wc5TCX[Y0GaTDeO@VCN+Q4W94^C^)fLP<+=+-Se0fDR\H3PbVC-
(Fc7bY-fV_K<cA(c[3:fMRV8dV#aCgKA5bK,RJZ:RRY+gN2RV/>8a>_11O;X\0/R
B,?M7U,K(0:DW<9LCL@^MZ:cS1^\FT=4L##^5VI5?NYR-=SQK\H3U;(K)R:CbH7V
g]d\SPS<e\+I7XCR1-_D#&TcO0Jd\D_.c(A;e\7=(C[JeLW@+L;\IOOKA1SV5.^U
2?EOU.-BZR2#b/E\&Pce^8YZ_<Y9Qf25\ZEgcAK8;BKe9eD4=:@56=gFMeMe-1D1
K=aDXg)QYC@(H\c;#2;[b4ZWb0e>YXa)RK>C8e@OV#XAQ7(AT][Bda7108;C_[YG
c[K<6c13aP^9/45-YQ6H(V^<[,5)ZSO??JW)^+/QcUN,[VQcVUL,Q7(<Rd[&G,Q=
TGHEZG4]_G&\=YRFBSd(>S+IX[P40MfLK).YS]fQ-eV;W1UW25gC@@M(;29@?Fg<
YYDRLM71+?ULSAbOL5=#J:XU(=X^gb_85Oe>,1JQ5IG65LW.PP23FL_=RaOD4f14
Z_)64;1@>^T6E;[dOY3/W8QWZ)TPWN+49-8eBR2LJ#+6#If_:dE9M)0/I&06_G,>
@+AaWN71;N_?fOYTgZ@T/.N:;g09B>&ebQI[__5L.Y<JF2#\X7.=,VR>4\Qd8Kaf
V^J?4>NYfD</N2@D:]1P[:H>;@@Y(c55Caf.):?:2eG6QT5ZHKPT]3)E[-R]F7:&
fJE=.3_<LEfT;2:fK7JFdGY#[QSA3\]Ig]<J1ZEBa7T6_<JV5G3H:EXB;+g&ZG[Q
(0FgA13cOZ40gY&_WRd3U0aL=?=,GJdJ&EP]6IQ?3^F>Z_MV1Rd^UOT^;f8+;)D:
PcN1gH(5][?Z&-CB\#9Rc208L=dG#+OO^-KfM^IF+[E)65PcS5cI,+aaX+5PU6@X
YP0[9cH.TJ,^K>ZWY0V)):d&=/F&<f/eJ1&<,Cd^U^\JDZZ@ZB6]22WIQ;T/M=&,
3^^>D_^Db.QV\AH>7=0IY]_9b;ISDTX^DU@K\QFHE9R0K+TU]49\G>7SHga9PCQE
f5P;ISSA+,]=B8^MdGT@^O@M3315[1,/]9W1&L^HFX3<WUEU/_cS.(,E9H\PMNLe
#X_VCP5-b6]6_EUc)6QG+fYFfB^GPaQ9@XV]U<O79C6<X)Z>CLGA1RNg=;b0Z(ge
7SG4/;S,B^+[UD]J\UKQ[=3^dG)>N90&,eUgZ/.#(_^>fDYO,T])Aa3.ecbV:?#E
4#S#-V#1/6e4X\RU&&H4-dCM7WK[eNVV0Y9&cOT(/3OUaGSO+\9L0AOHL=G.7T9]
+,8aD^gaBbQO9b^I]dOTg=.2^]ISY<3QDDGU/6H9\eA10QRB[18LWX\6.?]3@4QR
G-gOI5_8TU(8<gVT:QC_3cVWU;4LR8Q(W[14CWT(=^5Hb-J-EUdR<T-OXYM<cVfE
R/@:HY.AZ6K)^L7>C;LaPOH/+=[IBQO=I(&7McTad+Z0.(eE&eG=NLfACg_f3acI
_YZfQ&0AVQ0JI6,AFTLWFaT7&>R7?6^GX:HX>;]2/]F.QV8);5YX]WH3GaMI2cUP
J,d12.AHLPY;fB3&Rc?=BFR1X8+b4X>FU9K#;F];ZY6G&.\-7:[;86ASWWP2K/;J
2T/Y,a7;VAB8U)ed@e\?VZAY2^.bH^H@D^4dd>YcZNC\NT6+=gR]V8D@N<X,QWG0
JCL4b=Xf6ZV8AN,DR85Sab&E+/5I,(#OK+E3L-N4Hg#WK::NS073=QK>NA?QSV@M
8YY:/.2@(3G=CUHQZg_bUaBH\H;N1>;La[0Qd9OXa9NdOW-FbQd;0]NM/_>]XG58
X:^P#,\,b;0VgRRJaTLLB[If3V86-:(QdY,53ST14)O29,UYdKY<6ZB9-6Fa\Z[Z
)2G:N#^H7e4J5=(8WSSVDJG#@>L4F=<.c@+UYUODa/A4MdJTEWfXQI6I14E/PJF0
dE\Eg#1GZ=8E6HK52-/8>F[B27Na0R3]g<fRHKe^G/]@=^??)/O<a.1(>7^FD>):
M&bH#2.X-W6=?>W5Z0]^?.U]<e7=+NaMa9A;<e<-RAQ>2g]OB98X[LgGQJQ;]V[S
5fI3U\W&JKL&2Oa)cTXbVdM8B,daEYd=UDCIcBW5gNQ9;X2[,4OQ1CAJ9Ke]TcKB
<BWEUSKJ)Ug4V4fUTd>bEN\S#T-<YPMPf8H+XRF/B>+KJ[6C;LR2^RF07=,AE-E4
SLNgEUZ9XeGf65G@Kc0&:&/Eb[?BX9#3-S?C-?&CQ,+@?JHeM@_7#-M=VaQDEBN,
^&5^&L2AG(b#,[:R/Y(FHe9/MVf#=C=L#0Bg59H<&_^>:[(.?@JZD_cZ,PDZ=VXI
#S<g9+_8e6d@Y75/IK1,G8WF.-D=g\MO?9L@14A[X@BZ<C;ef:LYb,]SJ-ODYPF?
\#YMZNKWXa?=0J40.a=&8TE&^2-N1F8K/N,3_-gM7:@LMb=/8567GN9AE2T_W,O.
8NfP)TdH(\\-:D((4JD,\,_1V&cHD/Pbb<<J,.-Za94FKYC=_89BCaBDd(KN.(P=
9]ZF<1@RH\>F)WPZbQR2TD]K>,+Vf->;P9eg_Y^&6D265N9\4[#_++Rag91c5/H0
a;@@,VLH\A^Y#UKAIAGM.B/:W[-_QI8^Reb/TI>-HW0?/W\KM:,5T(+:E1SUIC\6
K4;UM[UH8DUL5FXd<U[PC?3BFda9B[GOf&NL9ab<XH2bJ\=8R80D2(7>.\eGL@#d
@;@H<b#FA2<Laf)N0c:[H>1X9dQAHM)+OM;WW33C=#FC&eVH\7R5(@#^(g/VdX6f
CC>5Y,RFRUH0\-)043d;U>YVc3AePOcQWREL\[0CG8X\-B<KSe_4,8ZcEA?(OE&)
(,DD&#X7WN;g?gFY/0D(#EIB=&15(&Fc[-Cb=ZR87A#4Z]=aD;MK(>A5VD#XdO-7
ZWK\Se6^YOMYYI,CKMgDX)\DT;W4a93/971Z)MGHA&F@Y<&OH=ZN_f1I0D:7Kf]I
/g?;L?]+F]>5\XQQR[0V#d27H9/LH3(EO)7:baLA1=A70F/+B;@)Y0fd2eA,1Q7D
<VaRac.,A0=90(X&#eECDAX5acR[GR,c+0BLdN&)2#M4U.5,C]a#H^-<0]XLTB[B
7f6.M?++A+/LfW<XLOa2O/,31V+86Qbd,SDYWc/;(b?KB:fXNGAU=2;R@X41L,(P
?d0GZ5DY3NK)P<L<g.79TJE-YeD>U>=?+T<EAMKY]bFLNW3(6cT,@e]#3;>LS,d-
F[8BG.-H@X#RJ]0d>O<B4CgI1,18_<OM4FJO4O,UTM/,;#aW(/6K844:[Y)dc(b8
0Ec5LeQfR)5IH0E+1HEM8X,+QgB]Ma0CgS?HQW4gLI7C3,b:)7D>O@\3;G^W2<=Z
YL23#G0,YH?;O..Zc//L,A9K_U(c+(E-:FS2R4g?D2DC&Q(N-OZ9[J-C@7cV)_>I
8:I@ZE&499W2V^O\)WBGR6OV+N-GB4dS_g6CG)/@YXWNTO/@EBL7?6OH87#\Y+NY
a?Uc/U^0WDIF@(B1B09XA2g-9b)(^>fR-[&@]3a-fX;61<4E#21;Z:aD(]B5a)-Y
f;1-:JU]6DBOdB(BcOQ>]?1#]DCFZFL2QeE@+TZbP^RH5caV0gaS#HX>fE<#eZg6
\?U<DVb)bK\RL4>9GgQY9HJKfATZgR=e&4A1.>eS3c_f6PBc5_X=TS::cE-Hd\.Q
0?(^DRX=+KW>32ED0D?QALeV46LISO&UZ&9TGL/1>e5Y=L1)L(VJ+a_df6Bd-8UN
S05\BFcd;B#+6cU]<a_P[84g(VLaSXGYg[V-J8dH^C/b&Ce;-UI?FbW^gYCTA&<+
OQ2\a+RcS_S\bOa60ZH8IHU>YDYeSMe\N#?gHd;2LQ04#5DfN,)G;8(#;)N;F@PO
U63>eTAfUXGS=<:bO5?;[gD3fX9c)R+T@7Y3J;,5SGeY?a9VH?+C;.[MeG.e[(^H
7gKL5aPd&>dQ[[b2E4=HX7O?(Q/R1Z-Ycc8MCP<N@ac5JLWdO-?eAY)#GV:G38]K
:AW[0,@MT-,=[/1N\>U38>=ce)4fP+b.+>F<6Z/2H\c]F4G/5C-&ge0PeU0-Z=CE
Z=.U.WefXJ][G>FaCUV[(_]Z4:;]9d1QQ#&\A&<=#&CId>RTCTfT]aBNO15WKPD5
cG(R,6Z\-E=-ZTbP<0b5eA6N]fDb2?A8PF--)CeVJ#.LNDb=6T@dQ3S6[I#_A.I0
1T9V;?CcM7+[HCQe5NYfg&RQNT.B7NK[W#F96.cEafgN]?QP/5,5@BNP>\_:4)](
;BG+3Z]M;]+DZ@8VM_S7UeVZQJ<eL^GdVWRZEL+-eNN/IH7Yf&f#A@/9]S[&>N5F
^JJY/2P#^fb>XLW1gVL]:Q>YYX)bRd@cJ36V)-759Y(>PG>e2:?D\M.SB<LGO,N7
3-AA\C44C5&IU5^LK2/f@VQ[]b3Z-U-UXZ&FQUbK6V[\6KT5AE0Zd2S7-2=;Z40Z
B#1><[gXM)Id<ZLTc4UU=_1e^b.gKUd#eTDH@]d(g6dIAa(_:</_Z\A>(C:K5cE#
f0#H1L.W;8TDNQd#D2Y8,L)0H;D-\2&4DJ)NLW=ZTTB4c1ZT6PY)KL1)AI,4&EeH
_e?,.Ad1)SNMfM]3\>LB-(6W2_E#c?40PbF]=KRGOG@,-@1:=O,L<.56CNEMM<S_
KeEM]0;:b(c()LT^e7d0E>9CZ0C51&@6WeTXY1R@G>#6g?bb5T7DYY6S6CA5.TH^
&AcJ6#[@a1#fR6E+XD_-X/)-]&2(_+VZWTYK&GG6ObG6VV+XTR228N)&5UF]GO3X
2:P(SfJWb[(RQF^N@C.,T30OXGSDDdZA71#3F9T7GBC^gXD:RM;:)7NXTeS#1Q)R
:&]J2fe:(0c)N@1J]fZ+>:QVS&WQ;P6AS_(#<72CE/.DDAE#WQ]I-OMDJV2_f3#D
Z4X+EXc7[BR:&2+35:079W:LUdUA.UEO6Tg9;<GYW)X3RdVG;.\81T;ZGKaSE/E_
TE2DdDP&/67SZ[FILcXC<((\Wa(U0D?IHQeMUDL5;S3WVe0?@Lbe^.4f<=Cb(F?e
#7.L?0FBG6<J0\ae6-E-3[UbH@B.)eXIPNT(G:TLFKfG?TgNPKWc?[:fI1XC2cA^
Q64[BVbZ(c9/RQD)SC1.6Y]5-;LdH&Z^NZaE@PI]-:D4W]^/OLNRa#VBT_#T-&GY
cWW7T2;^9,-G>ZK+_PYEPM_b_D,aDS4DfG70Y^H<EA=.Hc(/.1AL#H2+41L@R0T4
L]EX24>ZG]0=M@I,-<b/OZFPOaG6,TT&B)LF^#0c?\5JQR^G1K3fCK0gGR6S\YeK
K9>JG@B?UcL9@9Udgba.bDU_QJ59dd>aN]ALf3TMO^0;GT\QK=O>G5G1;J;QJK8]
0GA_=c5;GV3RL9.J4JZY/58T4X>JL_0V7bEXTIgR[WaZQ:AD,CBBZ.a1IEP2@gV5
SNS/B66.d+0YT4E]I<7dG8)<0)CJ,27>T/b38LU+-0Q8V2=(d2c2fL7^DY#/@K;&
,M:UTG,@KN9gKdK/12BPOIdf3@;ASg&\ca:(]Ha3DCUUJ=UM/eH=>&SBW>Fb76f4
=S+K+FIb94=/15@E8FKGAgKd^9ZS>,JgLC0UDI7^#HPb>DGIJ>2(87:6H41.P(=9
I?-J>]BD1^DY7LM)<4\0_<S0+aRJA[;:g\]53EE9FA///]I6f2BL99+4d?&EU7J/
0:/P]c&\V;ARLCI</K,(T3@g:GOfOZGKO2AYDc&-eQ?1APV0UOP+DS5dJ^V?\,7V
Ig7:GC&bd^Ce]_&?Y&gH)4T=FFDZ=W[E9Je=S:2g]WZ>46K-[VGfdAEQJD<_.)>&
-FObKVdZf;964Ke0[bP(UCV0R,1;.7+>Zc+ZZ#:4>AK>8:eScHJeFZ279=_P>GRA
gaCgZbVdB2ed<II[UG1Re1-1]Yef+[#)(6DRaX-ABX&;aL]-S]gO_,AYS;Y>[b=M
<Z447O@V9F:[(a0W-&9ILP#K5#J5D/IJ:QWK6cN0ZC5g+^WXPW;FMA##^+DW95O=
N&fRdVYP)./gQO2N)&QeC(YBb)Z.MGWD+=M:CMPG^&O>KBX?YNW6F#a\E@TZE)14
gS/bc=TOTcY5(H;<eM;<V;RZU3Z,#]4B6LO>W4E-#V?ZI@d&f>NNC)F&_SIBC>^A
>3I-PW-ZB12[-/:Tb)CY]\_YZ/O,+>JHO;ZDF:L)7Q-(8X)>bP^6-?:&,_TAA[4V
9PaI>Mb/RU.gMXY](a3KY2@+.HAAa;3U::D.+SR\=P?2;SJT)+c7^5>=5J0\AcAO
SWF;3FA:H5B,f>O-&bU=@N.[_bOEJb&aJ84Q2V/KDbF#b[<XQ\2X3\VW?U@2GM;e
8Dd07_\fZQcN9GO,;Zd:6b:XKZ]1<ZB4TcFUVFf3>_@77Kb-T.d98KWSHNFQEKVW
\365c/S881>@PdLBYD[DW;A\[7VW0Z/-AO0.Me53Ma5L#F(aAT=_bLNH<A(.TW=7
;BTZK+BF>^5^S[Q1D>?g(AVI;<@[_;57[b<DfR5]d/.T=c./fI8-_:=g3b)^?1?1
8M]?0I\Qc(A?0=MX(#HYHR=DZ]I\MF+G+0e.[eZ1fgT(d(^GG7D#G5[Xa[UUXc4H
STH#H/:2A;-5Q;e^)\g?DcMQB>XcTaJJ_8EfUZ_BeOgEQ/baUZ3V&9bYeA/3e,<Y
?WFZ]7IW#V><.b+5(0[[/@g)^,dA+1:+Y+F-/d.N.6[CAgYP0XY.<,/C7bH=ATMD
3-3Q6OId1+e1>=+(E?K\3;e[SL.G]\6P]<Bb80eM47/@X,V+1,-E]?f3(Z:5QFG2
_=:PJ&WNEPP5BBZ82b=a@XV\329IRU3V&C3J/D>3E-2-Y)IKPA2&I(e1Ng;gG+R)
F;GDT^EV=XdJ^_cYI-fYM;O=e0<14\\/I#P3U(79RbfB+^L.Z5L\)F5Sf.=]_A1@
+(=XL)/9@;Hf&:aGZ(B.AgCFOOcC#)\Q<X^Q\f34_>dK+5:MLNP5geR7B(]?,PMR
;K(<C8Kd8[]&4O^XZg^[6:LaN2\b4/g)44V-5fJ[,R\[b1KRTE)B\YPf+4G=C]X6
0>d8Y#OD_X3b))0GG&XJJLWK\f]TEgL/7_VJWe[(gW8dC?f1d>5@F;ORB41ZH\IS
,5F[9;^HLD7eTMJ+6QJN-Mbe_<^,LO@G;KT_#BD3>KS5M#&C?S0ICWE<fB7@fP5F
7AKI\=&]7_C7Lf9>\TF0G#HL?T+JNN/>&FN7(R@\eB<3\De6<-PHXVHIf1;(W<B;
?AL]]91FXSUaOW61#fT)#R+ALZbbHRG/8XXcT6A0P9__TKCHE\UFB5T1cG+ab=?5
<B,[1H2=?_a2B^dMEH0b72S7LM[aX^/4Kg\>@>?ZB]QCX1CCT7;GYaV@.4_5TFT(
O.B=e;/32b6Wc:_47OUV83=>6f[G7;C_[N\D?I@+0\,[^=RW,]eYe-1H=cI(J]H<
.<(Q.)6)5e=?1^3V>BWg_[=/G3P&9AE>,.VVQ6[daO3.SM)F5fBZ=9FC+.W3;5d>
04WRGV>Y7XE(]aOCK,;-8@RX[27NeaN4bF-M@B<8_1A2/TGbNCOg)^+5aaKHL[9Y
ND5L/ZWFX?L.F_K#A::gb?]eIW16G4eD+W:O?3&SgOf&ZgS^<a[H4Q_ge>c@<&V3
N<_CTObfWCI-/YgH9]=;\eB22;FDG;3CJaE@RO_?33aHJ_4QZ^:d,AGC4O&e\@44
)M<EJO)A<<MIS\97&7YL12<Ga-A)UP?2Q16GWI_ONgD;3dPT;DPc0T+8])I[@.G]
;P:_g^-X5@VOJ^=_OG8X_Ic)gfD1dXN:_#Qa(DW4DJ,dH9U3a5.+WQ.@IA8>&GGP
U]_#MJ@>fea_]T3eYfR_2/fOF7+<9_4d#JI7/\P8;A6JB1V_GM?fQIa8,.LMd/H]
QUHXY_87E1H3:H\b_@^@&KWXB_IZ]eXBZIT#-?[A8SN4O?>.??8\b21DE<eZ@f41
,b)VG9K\7BV=JX/e9,bO[]DEWC(1MP\E7R-c=T1S1J7b(L5T[ab<#C8.cb&H(W1&
&<=K;X4^Hbg:DbBD@N0AB[g>#9<E2Ia6^-bdYOY6ZSHUNTL+Pe11G2)1AM23dS@N
F\0a:9AOSe2cHA@_cLYU7CYee?[-GIY9aBfN0&,+De64gBK82b(=21Mg@Ib+/g1<
T_,;(UF_<QMS#HU+T\^\4C@>RBb\?S1Zg./IgU]FMa(6N3cQ[Z]?-S/aD8F8Laa&
Y3EI&13aO-:b;DU\4VbePLBO;^E;caM^bTc,0PecES[F)<2bJ.3e?^<09P.2eW8?
U_ag0d]_d_YJ)14Q](A/J>.Y[)1SfFBOA4+fb5U&B7M82[KYVH5L]#&R>6gZ4ICf
bRe53.[P[G_eBUQggTM]gJY1)]]ZSK7L1BE<gG@Y.[VT]/gIT<=:/dBf.PY^8ZM:
9=[cg5>).<0,RBIV9KLGb2^+>Md5#SQfFESAXYJ7?+RH.R&4e.UBD^:MQID].]9]
UJ^KX\3>f^aJFa>]IK#[:N4BJcL]0N3GVQA<3NIgM#\[-U1P3&69gfNU).YT-dQS
VR;GSd=KeEC>g[JVOaGO=dK]/-,J/(=dE6Q_\@:NDY5<PNP-EDF0X]OA?E(gY20c
EE#gbQcQcJbIa@S)>c(cD(<L[PT,YcKD^+ZR]?aJT0/ABO5G-PG1Ie.,.J]-gK]Y
]JSMYKC[SXAR<66K]MDM^5=:-^)RGFcK9^NFA>HU.cYZN<+23K6#e\#K]_c=MOPA
4?+_U>:[9XPL<f>W+\H8]a,.QU@d]C(@C-76d>[g\[^:V37(0Q_T:^];K[g-EOg3
bD8^Za^b\]T<f9@(/KP3cS,W4?QEQW_ZMX-3(9<RfZI.F1_H,]U=a6N4G.AfP6I?
?I67EI6@-=+NN29A@DQA(CRF#]]7?67e#89I#>;P0.#dUWef_/IH.JM<8OKd+Y;H
O7/;^_EQK6T\:,T@-][[PcL6O:D]RNC\cB.AF@GbBKCI#ZU?\Ab7-_.44+-+a\XH
D#U0ZOAT-4E,)7#:5?N0JaS2(MaA7Y&&V(U>U(-;,eTHeNG2P2)B4(]/L75?7#8T
OB(eQLd(4,5LT[PT4:]I5?2HSHCXU@=cEY[)ab6BLX4G^?4]-b.d8+/WK9,(a7d7
\^=1;<FUKTM5T^1IcR6bLJ4&P\R/8-UGFP4Q7>?,LTJgRSIYaOg=We1AW=X365=B
Y\WIO2G]Z,J_Vf^9K,@fA89+CERCSMGV?X=fdD[.?Y>YOLJ2=K/5@G5\fNbL]HLe
\;G<060(V#X7:O,WQcK>:WX,HDWMg.a4dLaBS@)VecM9JNXN0N0Z&;((Z?fHZaU@
V)OKU&)XG1,)Afg_&6bG(dRFD=dV,OgVQ=8DG=NgSc3])A@2;b9V2-f:U910Lbba
Z#:ONN>PR1Va7J,Id6)9aA7MPWH(0:>MS]G)Pe_OY3RN#;0/,f;7Ga]?3WO:Y_-B
HbB3bGSDP2QQK0NO;LfAe&+TOED0g];@b&@)4G5dEDGPU4CaOQ(9.9],04T<B2-=
2]FR(_-BN^f;9baG?8.WFC:=9_X\^1OBA34e>0==&F[&0311O5FOP_)9d]E?;HM.
gTdJM0^G7JARFK=0^8V:?4fB[(+F<MH^_4IL=ME7A4Se&VXC;dUE#>aFBbKJ6#6_
KIMX723,JX?/9CDRE04dd]G50.RO\FIRDQ7?+_)3e07_Z4\5:01]DQT=c3><WLVg
Jcc&619:,7^.g-1,bP2W\9_Ib1>1BfE():2A4P@\VXCTJ+4+B^aA7GM_.VM27)4C
EY+63R50FLDAdO9JGGN@YdSUO^3>=efM0T<U?#P0B2g@=/G:^U;[H0#+0b5[C]=C
SXZW,_7QKW_\PIALgL,.JWeL4E_AZTF&JL_-e7UVR#>8?DUA=e7W<=)M=TR3LF+6
^00-@H0XP)ZHST#f<1SJgUgG=K9HAH8YD(3gT^0A;RMG>X3_A,c2#0a4J(FTNN?7
D=F;@/D\>)adOD_&D_#X4\fHf.NU6^GR7VZU.[XF(\)AY@G>#Y=;QQ:S6IB<dMJX
HN.15dP4R(DAY033HEVI1J>;HEK2fIQgXc8Kg.QLfA5QH&5.6QA-WR[2C8f56efJ
(KLE=]Z]UP,RN7)55456Z2).+.).ge8dff8DUL8+3KTFG-;\G3T@=I950LI\O;59
d[b1ba9[UI?NcEOQ)/bF2BJ/eK.?;4A)6b&MH+#_CIQHbHd-a]1]FV&gTg1(Y+83
-)9aO@Y3-XFe2e]:N,T@O0GPFGW,>HFWA=U65T=MfJS^JE;3AERR@3:WX>1+5^:2
@PIMJ7c4CC]M1?Pf;L_30LRgdG@XOMW5IX&4EJ\7?9N4_<=1XQX2eD^?#\-aI.6I
.e9Z/Ac9C@CODcG8HU]EM4YQQ#fOEd/[.1I[^e(Q?JG=MSDIC,b:L#@aGN>PcL14
/V[(?^BL]Y6FAEWXD5Ke5W5\6c\c@R]c5F03cQJUK+SZE?<BV.eAKZ8<IbLHV]/7
BWOP,7@WI9)g13I7I)ZK.fT3)M8YV.O(@cGLAeQMa9,MLZ1<bE7K4?V-a8L@^6@H
=@WM4.]H#>_bQNO+YI-J=)<?9CbP0@P2UYP9eL]_&BBN;M;RCXH<MdLGO5@IEfAY
L^:.^a-e7eMWPN5U_:EOa=ZgF[_Y-OG933],3G31<W?8AbIaFNEUO)f/ZC]H].G;
8DK3PDI\-BG^HLWfF9d5Mf@7Oc_N]&Q9Z:H)E(1+C&e_WC<@=G5P2WT/@;G@@f37
_P)NeMa=T<RSSQ@PM+OaH=L;=-)<,f=D88).T9CSO\:^#EORXJS4Sd(Q2YM]d759
L8D\I2.e0e<Lb6@I7;#NcGG1<EVO3U@Ve.T[FbbfGaRBNSTZ3SNQZBRIgT]Vf1ac
.+[P,1EL\HXEC]aeO49&(d@RH>B3BXPIJg[MZP@&3Tg4GT:Fcf[46R=cK>;#.><=
@WQ1-^[;Z91gHJQWXZP(_EGfgBe[-CSA(HE\<//=C+)KLA]F^eWdd01VS\;7/GBT
MRV\Ya.5@6b5E7).6CP>Oda;V>.d<7G_d.^>84O3O58^0YC;307DZYEAP.UG)N7E
&=7N=a_=b)LOQZG@-Ybc\V;\COTGK.CJGXO-C/<[@>EgDCO.5>a]eK8Q(P_O6C\&
V>F__+#+O>M[QgM3cAB(R20^ZP;GTC>#W.gJJ/7\O,L[c+B(4<#](B11dG#W@-M<
LAP]D1?C\#(POS7JXSYK6]d_@2OR2KKN\f7aY]Ebb4:Fc2?/2D+\dC/c(^:7a60R
[1-D2MA\UQ5^UU8d84M7e.bKE(cN4bM&EW.@FBCD0OM[)Y^0\N^c2891EXITVV(G
?KQB5EK==/+[&L(3.U=O3^QYL05ZB;g:&(\>#&d/.)[5gH\2##IeL4NPG@\^(g^\
d.=bWY_>LJ3(D93MTCNC/g7/7dL9WYLW7@ad@^BGb1_,1HK3KaR#@U,[V75AJZ;<
Q^8998QD3,]:>aSeXbTK1OT0bHJM9F.A1EIG0#WN<Rb]fdc(+?f1(-^6A>@+]9;4
=JPVLcNO:(O\JL6WXW.^b;^2HV9,4U(,_a0TY6cRFg^)R#MD;=/UH/J#,deK_>(A
SVO[g8&6P9bVKd:U[dB@N[C>HaE?c8A5HR\#K5&U/@9Q46V:1eK&J&7YSH,Y-Le&
N7\G<<WT1RA@WV.=dYg.3DH@bKGdE&C0b;[/5XgRGF5,&X6R@V,<KXc]8IG/?L3=
YUBDSeaT,W4FAfS-HGNc\.,/7@<b\\SY.1S0FBOA:F_Z:#Q)1?U6OaJ\9+7;R>Zg
A9E7B9X0;LT(>+ALQa=?-3VEcfG?Je;]#N5W8BfPaD,YM0TGX#/R?OJE/SW_(T.:
@c1?N3U6JST:YAaCbfaQ/==]_GMA,I_:T3\DCLE/d9d;([0..&/476)]:Z8<g+[I
DPP2f?9N.?&HM[1;L[CgROMCcLITb&6N8D+@<d^23[@@;ACI[]P#9UE932&>c,()
J7NGWU/3G-Sd5_OeOSBY/-cJ?T4)XN3>P8;PK.<TG+-b]36>e/B/667Y@-LVW>Kd
c_0gO^V=UK9RZ&VPFc_TcGC_],P@.70P^:(Cg.O#CSe)<,L=49>\=[83-;\K8I7;
RMV:4B-6YW,10Ub5P+9g5GYYA8(F9WXLPUK_#XA94bVR2E^^.3KRLMN=C46bgMXF
)LdH^cT4NHbg3_DKH\#e2G0.P^d5DX9bLG-EPgO>bb8.R^WZefdLJIPG#LIbBJQ(
RV#ff0=_aKD/ND4YINVT@L=YW@06V<_;feg0F@]JZ^5c^VT#HAXfZ+c:3WI:b/7\
Q<C)I7L()\G_IO=F,><-Z<,Q#(YD4>4d+)>:X?I[+SHP7bN[eDL:K2=H?/77f6Le
?QT613XH.@NZIX:LUSRY6ZcX5MePCLC5g;e^-4)29I32(cT[/5M16AcfK@fHIG+?
/W^O25()I7A^3X?e=<E:c4=EWHU=8V@b?VY8TabGP;,M8P.;XJH7-bO=0#c.(TA(
\^&?+RR3LPQb^0X.;X)G0KfJLYYa].TF0OJM-XMEe=L94#?9AK1_#Rg4RGN\@->=
)12H)#BEe&)85V<@][\BNCf@L\>b0L?S_\7c45JN)NG8.\<6PNf6e?;=^RZ569GR
;d8WNAY:8BbM7^FE>\O1YgSd,G>/>[J/aD(Y--^F[=Z>)dY4C3R[2@RWPL_+.PeI
/2MWTFTSMIYfEZ_,<Z))G6_bXOFg/L:9\gDB9-5011bB:<dUWM@L/G9/<>RdOM=\
A<N-d5cB]+\1?W\#5K36,^D\HIV=J-?Q2:b1.PC>TY^J)?PF^1:F4XZ?91c\a+52
)H[)H/fM-IS-B8EL=+04N.6P7]Z8/JZ8L0<3W;Y#IcHeTN1RcW)2fUW2C;T.07dO
^6,\/U@2-/J\aV1JBR^P0d8(:)XX?D(ScGB?()1\QF:9@+SZ[dWa#RSB[+[?6cg4
XO3aDN<=FM-40E4/;>S.bfNc6?6?7R;:,L=f4ER>OPbc1,A4WY?I\M&#MCAJ9@g)
KK0-gNO.,YJ86@:(/3<\O0X<4aK1P]Y?S5L;J[^aMGV:VSf].]YELI#e6&VVbb=;
JIg<_0>8QObH&TEISSD450T_>YELI)GLP?FI5&b>VB^XMD:cW/b87,H>W:6_,HD?
E@E<&J@eLdHS</950<IWE7;7[e90/05_25_<WW_LfBN<ENS(^>?3@?b<cN(4JV:F
SY<<WQQO=R@LF8F&QbIf,ER)F1LM\?O2O]1M2eK/P@8E\K-5.RWUfE+VG]LV>BeR
V,9[IB/Le+Lag]eA3,X@_/E@WXDMb_MI92XM;Uc)X_6e/E+?4R?2\BeYOeBL6&-8
D(3ggc(\,#eQFAP3=9#5CVW/bd8QM&MI@H/Y9]gD<bD+^>G^bdA2T4YHG5^NXBD#
U.G,=68B)836HJZ-QOD@RSXFGK:UVaOP&S(#Ub)EZX[Y^U8>M[^]BAB3?:9X;^56
gXZZGG_ZP&4R(_B^He2#A,dc[B,&HaMLcJ;E7[9aP03bP#O.VTW[PH9);E7<+Z5_
,<HI/A#=^aEE>FKEBJ4Pf=OgM9^WI&J)LWcGP03M#MQT&5Q8[PG8YC>#1HYd(=:H
fR?^X1FC\BDQ245NV.7cOQHG21.K0Jd:O4@4^I^#M#0#XZ@DZS_02B/+5#04WVge
9a]bNVT39Bg@OR+:+FI<R-G/Y[]g-F(23BZ0O.S3;.gQ@bIW@-;,4&).A;F[4O5O
639@^EF3&&U_/bPcf@)56?UJbSLFZ9^.c4-[OW+/<PZX,<C;>E):1cc]61a<MXB>
dT\fbD-bF/YLBQ;[ScffDBd78S&S3(53eEIF\U1eg]@dOQM3\?TQ).3W\6Rb5]\)
S#gCS?A@5W#3gKYS-8D1c>F=K:78JfG440<cCL+80A+V&d#-CCTa-F5Fec..2fbd
;3J_F&Nb2]4K)B:V9:2C(:@32LTOD,9>.C<(?acXHW<S:D38N3B3RbKe0d]U3Qdb
bRW[VJ@fL4Q>TMTT7N[J4A8WKc(1C0<EDW+7+44044#:SGLaF\\(c/52L\_,_X;g
=Y<(GO<JE360@=[b@,D7+SIZYc3A#OOM1\][:&O@W(5;#/2X^#VJ92.=5PP</N#6
3EEUdHUL:.5aCF\&<0GC6@(AMW9N=XHZ4_71?.[#L#1cH8>O5[]L\^;&YHcPQ:U5
ON]aEd\0#IM1;bT<P;YE=/,IE1JH=Fda)0(e(W>0@F+NeNG:]@:?9EB:1:9&dc93
3?Y@WZLDX->gWDLYN.93]UBT@.9WGY7OfL/)R/>;Eb;gPf<C#RFSV&f+XS#J#:e9
52RRJUD(15SSH=ZECba;1&A^,4bLTfGW_<-?bb_LYVJO;^cY]CF3Cd@0:GQJIPV(
bNaLVUce7.#09#:@e^EdT]T^SR02gTXDfNA=9#0N.PD-VZR+U#K.V3I1c(dAH/S#
dHJF<bS(g],V:8)3DbN(D_RE;VR?QKU6:EM=[NQ))?AF,=+Z[SA;=>SCX[/1G5+]
41IZYf]T#U=Y[D,^Ad(GY=HO0@7G)\1WKA3FUgS[1RL=Y+GQ@[ceO6VaZ3aA.g=E
A1=ADC49eY@,UBK<OQF=[?QVZ#&P@BacA;&a[FB_M#K./G69/gbK-0,./(AOd00B
OL[aDDHC[f:ZbUL4fFTHc<N9R9GPX@_BJO^c7f2^#G>g\@R[EG..]RMD\GWAbMQE
7d,8K)(FD4N<59I_>9[M1N2F]>QTWMS72AAD\NdM?I6TES<5[D^8GY-:_@RFaMLe
:fFXT_R:-U2a5P\]0X>C[a&:;.T?2H#DJGJ>9YH-\c[3KY;U/])3-N&B+)#)fDMC
G>RXeH78__V]FXW2F(:6He@gULa>)>0>]5#<F6EKWSOU[bC4J?DAS]ZJXV[REWAL
6<(WJ[/4cNQ4X\g+LF=Rb#9f?DU0C1b>7:&I2(_(Z&^aCG-AFS^^DO_SLODdL]3L
<IA^I(D(8^?6\=1)UQ[AGe5Ac]._.K(\4bH],7]VC&S&TGF=BOEeWF)1F5-2_S_H
)J23>[Xb\1#5A#[4O&:[Ffaa.Xa5_BfKJWTd&NAL^PZ-K6g6[<]a_f?<CG(fW=1e
2G7ZN9B8Q9N<^C1VK.3NG^\MLPLQ[X_SNPKQ;&[@E[(.bZQQMY=RH/bTaUa&0aYa
[J([W>ffL(3)F:@eU;4;Vd63B>2&MMSWYF4AU@[S&WeS:+E=V&0AKZR8)e<H=95;
@0gW-S.UEZ.@b<(bX.&6WSUY\#5__<+LGCY;_,7.c[)J7We)1Gb>R^/-EQ5f\CXU
5N)H4N,]cc1]H)C>4D,Sc=?TT1;ISM9?V.Wgd+OcRT1[^2OK#2Q:W2,e-N9[,GSS
(QHJ2,=Y2C6WBdBO/72B7)>YU8Pc(g;U@26CI-,50c)5@&UUbW\_4?XO,_3)aN4X
aJ@RLg+M12V0DKU6A4^ddY?_,\EM0)8@(<RCGB0@NQ):V=gg.g0)b/c=WPbFB&fI
@?[-^#VR@]M;\VLKJK))FT/[=NRLY9g[/.5]XGf)Q\AH\+bS.@&:gL_2X=F-@aFc
#F^a)LbBCQR4NPePO/,4TIELTY\^K)2d_PUf/IL-4KTBUMGdD-?-be=<fN^C>3I;
,U\,c2IMc@c+>>H2&;d]f^R/7\]X]<0W<EBR7O1#U]?37&:21b7]0)Ya/&36_[(/
YS>bW3CW1SP#H:HI>I:Q@+GWCTP@cUEYa#9X5SW\45?fP>6eB;2X,?a._/1)36GT
,dFTWcQdS(N=5]IP+b^?PG50W5^eKTS@0XKZ\c0YSR\[=Ue.TZH-M[7d@5d-J(+)
9R.#@+.-G_2NC(#(OLI>3XO#RUF-7W_aBe(>,096HFEQfO@)[-)W3b\D7ACWJGb-
>.+1TE7gCcbdcb80OCKOH,\R+K19M4Z/0:)GR+Y,W?AaOD-IS830KO5E.K4^YW/e
3S.PcC@PYgA/I8Cbb-.Cfab@520S[H\G(e8V8-,+HV]YfY>@:KRdR7S[84/_d/.A
aZ.K9\03>._R?&f\-d]WaA)O3F_b^5)0deV[.\8cV9Z8;D0K1-^b7F7\-4?7,::5
JNTXXZ,C?V>SM:6Wa7#V7)HF+/_aQUAJM32_56@Ob3fQW=U/)<+CNN8#H=gecb##
GQWf0IPGS3G1d[S?)H)feU72Yg?Og@HQT)WUBO;>.=:cf)MNW>B61@+\04FGHgU8
fT/(EDS.?=Qf&S[7LaZA[0SW6eCRP+.P.cTDGMA<SXK-SLa6YQVZE;eE,_G+7P1^
H#<N[=,:gVRIHd:^O5;P^.FT?U6Z:,I81O9]PG#W+,W\=O#K>6NL03WZWO36HePZ
+(HRBUD?g&PQd+X>5+,g72g-@#Ye):\T]?61A.L(Kfb_+aXXS/Y5OLNcFQ:5:W@S
S)?[O^O>CVCDc7cKg8NRIMBW]96(<:L&fd76@A:LK>=aUR6;5dAfTA>4d)e?=]P+
[?X<PN-S_JR]FU^OD_EWDXM=9=(<E/0-?dI+)#X(+dS<;SVTBQ3)XJ.@W@-f0@#A
@c(DbNQIH&.=RY[021>b:eY#Zf^8c+^[+V7O(Vf[0WAL2R79DJRO+G1(;eWSU45U
8/M>I6AJdB;=bLKO,I,#DC8GM6V2TG>gGADb-[c0SYdJ_P,eBcP9YFdgBPY1Pfdg
YYA+^9FWP\B>C8Bf\61BI[ccA+UPHaH&6.H41D]3+gBTZK?;Y1O#I4?)8@2+33-0
X)2^=/gf)cgT>b3f<U++E_^^\2X1g(aQ^Qc0PCa,C)bSK3VaV[E6>Q<P,DS33-?\
<O5XFf^&fb7X\2L-V,Ae3++6JV3UO8bL=TBG(K)1Y[U(cC&#LIL\RK.=T+^)BdES
VDTg2G+Y=_P:02\N;:=8^d[&-XYTc^_BWN88@#Abe9)@YAT\X8EbZ.5/<6+(<50X
MY6G]1P9Z#ce)LO,0BBNSW_NFUM5Ne<T>IV-5NbK&]3ET<NHf)Y0WW(T89)@U,7]
)]-J;GfN-Z&J5@X3<CU6<e09SD#+W\#NNRfAa-K2GV<)_@SE+P;H@HU(ZU1@Xb]G
E)&R0D+Z;XKcFWEF>@/E^bC2b5AU</6U[)MQU.cZ+gFCb<UPFCM7H7SQ;WSN;7bS
WBdd8S5Z]&YRL=S:Jd:bbHTIU@e&2g-6cI4098=.<A-(VX<9PVa#eBY=K;_\0O\)
feZDBe/68ZZ,Y#^d9^&E@Y/F<ET=KT=JQ-G87Bda+RO0NQ[/gbZg7);2P.N8@L?;
Ob(COHVH1SD6B6V8K@A5=Yg/gWLeKLeN/]AM.\c<HE<5L\U3_N<P=4/X5[cE+K+7
C=d?ER]NLbX+/-R)=e-Qc-F82Z:HZ^bSL[4B8IX.EF,&dCQe2)9KIeD)T^\@V,_/
U)7[WU>&f7#E;aD+<FZ5c@(GY^1HFEL)4-B-5XCRMe.dI.P>+a[V1:?b5I44Ec@K
1UP1^;-:8[EUd:\2]546ga-\FXJ\\4J4b+0>R&d>.BXGd<:M,IV1dQ2Q@^J]_O(<
.5Z=/^Xc?IF0W6<=QG.8^#,,9(^Q4\Y+710B)bX<^,[>/311d^<D=c>&J1VZ_gQY
cag^=e>]1DB<<SN1=0JGZ;4A@,:Wa&3R(&A=--V\PKaJddH;</I<e\\1+MT0aN@^
S4?Z;(MQJe]T@7g;QP3-SS/f+YMFN@:3:(]5g2Q:29R)&N(9I0JG\@Ef+D_S<e4(
UYKd(AK/Q2ZMA(:\Ld87FQ@_TRCd#)#6[#FH@F8#H]aMCV3FRI@gCRB_3gW49^XU
.,F=9eLQW>N/+\W/B,\+/3[>F^1_ARY8_D^MFY+fe@aUB)V_.NZPN_^VQ)6GX^.3
I-;0@V>]LCV-<H,\0_.24;87VGVD1XE@/7(/,-1M].]AE=+7-4?fa&dda+bF?7aE
3\\6>+/BZAQ^NFXf+8NegZH6^E:-,R_BE<(D(f;;Q2T01^V\AGd8P7[Z9SLNS?@_
QAL^62K=7H&@&70c@VB+0<HCAde.Q,?L@^[_#+(E4OfS4.WOBL5XM]_gC,((3?eZ
C=,5;Qa3W7N54,]/RO-WF>WIcEBA)cdY(/5ZI5/QQQN?WI2:Ga;=&&K_<#]cPYG\
0&<e\^NKYI50T\JKT8G@B?ab22#;KIQ-)3&>UJ>+:VUB/YZd3-LNT&#^[CObNdc3
M:@JC;D(:^H?@QJ5gE5T53E+#\1_0QVS7TPK\M6EUda(F(U&Q6;QK\#&K&QCLeHO
f=7A:cIG[/EB.-LK=J@;TJ).?HVW3N)_HN.VER,GW0.F>KN=R67d(7[_U-XG8_M&
-NG/,I=e]cOc[7_L>5B/^&J6CJV9N-P3B4:<EDJ,,=>S@bb.R_\AC&-f;;SJJ8R9
V7B?cO3HMR]?5^/VZS&5+,a0=]IYd.5b<-^[:1KI61cW8gPc+ZNNC0#>P)#O0Qe(
g8YKICa/[G82TX:VFL^@RD0a??UA)?B-g?0_@E73/(HU0J\^I,6BPNFCYUQJ2=])
K9eN;9PB[d^A.LW3FYU@8bZ;CD2&QRbBAEBQL8QHc>MLTY88BOgN9)61Ed,,+=PG
@.Z@^(bgG#]L(gM\3#MS)IN;-),d#T)<&+O3J4USc0UVd1MUA,Y)/,,.HVacOIO(
Wb#<adceM,:AaSd+K^Kce#S6@O[,3>&XfQ)<[fBeI=CCU7E.).RHF[Hf86LJ+<CG
Re+Be^:YcD(3+gE5#6G\L8OE5A&^9g^G1H&]-_DJ(KUUY/_cM5__PFCEK&C,RUVU
0@T?@_K6DLa])4VHQ>-G\.?I\7K))c;1=]#)(ELNRJ-<PGZ9BgR[0>DaYHg9dFV<
^-)d]P0Y76NZe,:[e:.VJT.OEaA@)C(#>&XPYd3DR,ZgTN4H;/<5?HMPA;G?VN1Y
#I>Rb9CANQbCWSJ_[f:KR-ZAX#N^ABQ#a16EMHFgG0ScJZV:L<^AGH=PYGU8cL&b
He-JTa;6/Y2Q0f09CU=N,PBa<XGCY+?;(&OFGCAQeJ5eH_E1gT2PUB?Sg)P#5@/>
),WK8A53L3N&PGa/6W2;1G((fd6>?dHX2S^XHcM.[U2_[:R:?.;58@]cg@86@:I?
0IU-cFT\B=J]94?.B:RfVR^G)QNf6QSAH>E.NP6@9BgHbFV#9=@1D#cD028J?7@&
0)7<[^@Q6C.\ZT\XKa4K=37V9V3S8M7CKQ)+3K2IY,L8A_&51aAR>B-Vf9JS@:8U
b=]XcHG5MTKX[CQIcHW^<EVeW<ZYLH^ED#VdL-/,&W,//GV<_[aPZ-Y?]9;8Y2;1
67V)RB7SCRMBCb-RU\F6T;OXS@1/Dc-\R>020)bKF0PdG8+01CG0c\gM0,\3HU]I
M3U\.e/;g:e1<BEG@RDCY7ISN>IQ^/,PZ+:&1MZGBZ+-3F9@^L@UGSB3+a^dIg26
VHI4X4Vc7Ca.XL2<89^+56N)F26&?T#=8DaM)7ZA?G=+NZ5DC\MYCVaS/8BD5aMa
OOROKHJgI&AU4X7PZ;cR-7:]#PT=;>.B,]IU)6C[[DSg_Be-FE:@0Q3DV#V.SCG/
BN+RDM](e.R=He+_5H8QBB>QE===GbV:Z(;&U>Sa1C0Xa1HJ67QbVY]YXTUB,QU(
<<D&KRJDTa;f_-J]C/A[e)d_K2?B?:8aGB.J5-HX_AKB/&;3=2[9DWL2]Hf-dGF1
MXcDb4OeVB:Q@@\\)3/_P-da<fNbG7:T.S8OLa/&+EV+9c3g72Sa/.1)X5eOfa]\
,18c7/)1:F<5-6f:c#J=#WP@@QLNX[RQa[bS-fR&?UI+,XAN>0]++(6C,8L65VV.
FDP&2\0(>8M8O(B^.#/UYX\:ge31,g8&JS6?R2Xd<T8_CI34798R-0D->>VE[aOO
O@eH]<I,bZ+GdS>[7T;4XP83SI/T0be\(b)<P.MJ[6FI=\O>K/-?IC8SN)J;JC69
=FX3_-7,?^HM>2bHPDcWDE?9&a8<[G6+;ZSJU@[G:D1WYEY-J]_&SFF5fFX?TJ8:
4GeS2/#W5UJA/Vc/A-Z3&g@B[BU(beP)TBM)QT+N\YU71?X^KR-L:gQ_]\-E]R:@
5I0T+^[,]8@JI;efO)aR^PA]>g<PN3L)f82Qb=\RHcdY_<e5aRg8T+cN@AQG\4KH
2\EM8Uc5C08J#/^_QZU7>2Ff4X[/#F6Q@DWEZ5VSCad(6DZfY81MP1R(e;/I#HGX
&3ea1G=]X@\3\^1KLVM)1_:>Ob<3VBLH]Z+I@ABccV;=STYTFH\c)?YPH.gP&F0#
T2]+Q2DDNBSQF#FFB[>&Md1##)&dW-_;bHOO1.Se]S7\_d;+U_N6JN8JD4H@K)3e
A]eI5J;6HHF?96HdbNIeHTX[9^Qa:\g,TKKA.C6^f#A[G4]I2&RH10/Zg=8Ue8X-
#2RH(/Ua(])3(G[<&SO8>A?OebZ0ZLL535LWZ/(+-8aOGQ)26==Meb9V<KSW<&4B
RgT=>SU<887R5Ee)F,F4]gEa\9JCA;Jgf[B007+P(+X0e;)^K=LX#9a+d5>H#,NG
4BdbL,JI,b=DVa0\FEXX+5[9D9YGb0<?MO#Z5::Y-FH]3g-I@^&EG_#NM-,U)aTA
TF6gDYd?:S_FT9.(I\I8Z^#f.]cKd>=0:ATXNP],@0#+:d0)CeYJ:8Q\@Y;d\97c
0Za>0_;^K+XdD^9C,cMe60&@;_#C.5SBOLDbZB:>XG,-<L=dU<X/&OGbE/),9.9;
#g+aU/,1H<1O#-4)=,_:<FMBg]SX=GEMPF1S=Z:3MJYCD6=YA2T\=9U\G]O<<MYR
-RfJQGN#GHCgXHH(>.cJ>e.\:3PY8;S0^380JF^IOe39,OagP=ZYO([N7R:W?WEI
8K(&1eAH.LI4WCG;>2R6X5D2B??aU^\+0?3=Z>1M][S:9AAQUJ#3WOaG434F?1O8
5;D6FJ7c^<IL]H4?I^:4R(10-dVaC=&4G+_S36101N>)Sc0d0]13F[@b_BD:0=)V
b2?)f?4ZG3UFe2R>EULOb<3SARTfGXZf;L@JXU>(VE5-d3cQ65[Z4#<3VFZR.,]c
C+4GQUgCQ,ZJKS^-F1aB(V><(dYEYaSIU#;(@F__5W^_8D/0G\6Tc,7+)61fea@;
0[6Z0Z<W]S)f79(J=Y2HWMcCUE#L^H9=-8EM4-FTIFS:YX?d+QL1Q..(GL5Fd4D,
YVRNbe,,WP<6Gg8_&:H6[6#H/T3Z5gWBb]O-1O+86&<Rg-XZ:R?AXS7;<K:dVBgV
B:J)fQL2]#8=/;/OYg6XKFb.>ePbF1,TbK7J<5#EP2\@GGebKV?,Y3QA80,/7SP)
e)9ZTP@TJ60,0Ic0Ff8]BcDE5D#](a]_B@B671)6H:1[[UG0;0+EG:,1P\SffC_M
daEF,8VJ+QV/>(,^a6NVb_-29@L]>:,[f[DNc:(_,HE=d2,RIad,ZVKHRTD@:FJ)
-O0QaFNLc3IPe;Xf4VDVL>?;1ae,T?#\@#NU/-<1JfZSd9C>&J9dC2X+aMHeEQ;W
/H).P,7:3WDO^\?K4A2=WdEgG8#:.7(#Zg0<.e(9W>?]XA\J/V3C5Uf_:7AHN3LO
B2:^08&bf=O_VMKMEWYAM+8(8+cfb2(g:9O<EX7P])KSK>KTI#)7BCL8N--\-dRS
82TLPRGWXJS=#A9YHbTUb,QU3&HZ(4MTb/XTH>]L=6Tg:;G[g[+f<HFTTA/eaKdg
Y6GCO&FSV_dBG\M/8_,L-5?g:#8TB<4IeO8d^8=J,24&ZeJCNa\Y?]?fcTX\SH1@
_+9&I7Ka.6N>2(@[SG9]CeZaVCK+[:V86Q+J4c0/0G&\Zb<#+5b1?.0]]/2-3:>1
G@EZ??eae&c(eCfDePX/.AD&F2761<QLa:\Rc;Tfc(8Q)8MdU?;Sd9S7XO=fRdZ#
LOH8Y\/UO@4B&9eeZ_bQ#<ER\4BA;<5F8\DQ97YT)Of<Dga0[b?RM[(5c6gYDNb6
A,d(SZYJ?:JX]@.N:SP^^78:&)JfKK7,+&E2MYWIdA#>/MM9db8g;^N1\D[YNRBG
A@K&J4#>,@9.4+X.D#9[:FLA2)?GG5.O=P<R;G>./61:B0.a6>]NCXSg<V6(I=QH
_:M]3;.&?>WQIH/50[CD5bf?+g5_?T=B2S).e>\K>Q\a]d39T\T@Gf?4VFPLPB&&
RJ>#JA2[^DP3f^2b(URE=PF#eI+4K]Q=DJQNa.U3IZV:3?3MRZARN/.JSH=d0cfX
2&B5\X@=&A&;;I_N)VSRI8(9@bFd/O1cgCUVZZY_=F[L)I.P&W3Q.Sg7D&>=;1W#
3E97Z_fEM/d[7(C692^)4[HL6BBLJB04P^Q3A(9daWZQ\R?)4VaMDF65(6MVJV6^
FQfBaELIJ(1RaR).,aa#-3fH7TaP9J\HB-G_VfTS9S,\#86631?]W:2A/48,E;da
B@dL\JD7>G+^D[^PZ6R1V=VZSKe3f#e65TGLFfMX\fL5^S29JB38]bS&-;a0U?>g
:,VTbM(,CZ1a&8faaQ=2a&D;;WE#-^+J7_1SUGCBX5PI+7#aFfF@+B7#W/28gT+,
SLb??RaSU[^#U36(BFB]^IWDP1ab632;E#M:/RaOdf&,@9TA6VgF+&3E/dSO=f_b
@(IOW&(6CebXW;Z0=?BTS^8?9Pf^ZGO,bSaEXbPd:.?S8FMFYd?R:9E4O6KDZ7[-
05A8]_Bb8-U_GM,gVIQ@<PA?XZ0W7Y:S59)/@f6KHKW5IGC^3]U^9:#AE,L&\>Hd
.<H13?8e3L\d8OR2,dg<3,^>4>YE)A,#a4<UW,8L2TXB5/<VfE&\XgC8\Jb04fa_
d.)RVbC4<^08()F?NU];&,/3YM-JF7U5B1SHWV(LHQCI3XAKUZD^^PJ;+KU)gJZg
1/a1[A7J-/=&&[f<ca0#..gUg)+<ZT+:JWd&aB?E5?^g=OG_e/0#aHC84#5IB9AL
BUDPUBM3(XG/d@cQF4[>(9#RZ=>1+@DQ1f2Y,,_.dUdU9/\<+,-Y4<8Yc8X?8-a;
S#DMbYe#VGW<&W\3C,762T./#=[;]ea=STScf@06H#&C;=YY;B:H-ge&3C])M>J@
+#,:/^O8;PUOFYe;Mb1#aM/;A&g&ZN8E?bALP&OLC&=BAJ?#0Q1ZEZ.1MUf-Ld2;
)A;(]d&:AUNI&>)RHa,U]+HP./6A+XUQC8Za.0T<dZP]GKaW4RLKDcc\Z8QX&XRJ
5-_?Q(T\9G>5]=7=4(Vf;G22>N1,+_Z/-[5Z6HAVQ.^6=9/GE75ddGB1-0?c//&:
MDU@aX>HVUSF,2;4^P.TS5WW@9WL[68VKKG?1@DgdZ;&@@fBK-V/SO@15:d8SS1:
M6MX(023P?WOe,>d=8a\FDL\NVY[NYf_M],-+@Y8>;]/>ZfODB#2C_XcfBW,)P0b
G#]X+@3./BRMbN/@cDgg+,XHD0?fg6R#&8NU#X]>BN4&-S)._c(=Z+/>W6ff&^J]
/^CXd?)^LKObgX1-@2dLaaMJJ:)GMNDgFAH?,IO9LO#f./E<ELWHO_4Z_fL3]cd@
PZY1@ZgE)4cBb9;6M1Lc&I_g9>WCe;C9\^D69fG+aD,@UH5\:<^&9AZS&2KEBRZU
#C;,S_E>]=]=X\KGDENWN,?BfaG7#PMVf?C=Ob@O7^AT-F&eGSWB=WY,PTEa]FZG
Q)U_45=>7_E>R,Hd/,6f]7-(JJZ^U08E>NYCA;+CQW&BgA0A7M0OQ(\HO^9dTZ?H
EH)BV@[DUMH6:Q-,WD4/^(Y8BZ?4(<H)f6.OS.WI;[+VR9>U#1AdS:f3^^3cbbV4
WW:8U9Y7E8I]2FZDdP<A0+d\F]Xe]@a;cUPe5Gd:G;K4.VHgWF,]NATZ8F9&aNY1
L)bcSQfV?PW+ABFL884a=)RdDFE;b6G>0bF)c#=KXdECNO1dMX:EV_UbQc;GM[KE
XR\7a_YV^Z5bQ73cRNRP]2VTC/YI9N[\fV.XgYTK]5BTC,8dMWK^HQY&H#20Vg5Z
E64&W3@RG@\#T;VP(UL[MLNP-aY0^NN;/4(;5;S@P[.HU_3V#L?776>\4FE6,@:7
Xg/g8(@DA+&ZJ=)HH[\&MKJ(CUQNXWXGX?WH[B)2;?;GAPF:5a[:PQ:Y>I7\eD-+
-fcRP/<fSA)F22<GeV-ga=4YZUF]g#=7U0&R,X/YU=6Y07G6#I/.B(:DA@V0;d3L
?-+U]F67\,_Y(cV?9dMD./AM+R=-/O6]P@Z&>Z6@10a#0=1#cOO_NYWFH]U=G:F<
-WE/?0.b5f0A@_dYbaOM<T@-S;+F=.IOV.6P#.F6LIbFUEPUB3JUPd\b.1]7AEET
25C[W[(NA89&6aUFR=Z-+XGEUZ_CN3,PUV^DJO45c,[,B#^FC=^DZH3]2O1&NJ-c
:&SFWVBT3>3CfC9ZTe:=>;LYRL\d4/(-W:R5>QOW[JAbQcFYf6/Ab4R;K9TN)/VZ
aT6g&VD(YE3SaL8T;fH,8T\9Yd#Ug1bLb-[SATb<\>AdF=ea#N)0MN);2Y[9O6d9
D^<W4FU=&1WQMSV3afXPWC6+0M9>/.#6D5?1WPDa0=)B??_\2FdP9Kd=V>);GH48
3--(P(dJXI^M0BCJKY52>@^]1O,/KA>IMX0bNCBf&\W3S3#7^_K&LEL494+_6V9U
YX^b]#X[LWB5U:BO/=8g&Fc+/]LV>d4P[LY@?aO;QZ17_/9H9Tc5;1dUI/KM]@(A
3>X>(\&2<MQHT[b)&-SV1S#T.?XE-B1G?<20e.#cZPT>32f5C)OY@aLZ\]C>LDWA
Ob0g\[1.I9bWNHY@ZD[3W<&fXa3<OBfNF#9X4)=CDT3g(731RYScE(@MX[_RPa2B
<+ad(P6]O62+L-?,D0C8V6f>FFTA@bR:1,6CL6IXX5O>\gYDAVWMc:80FE3,WCU5
808-Y67bLX^gWLL#1XJ8-cUHG2=AJ23DdKb(eH0c,bQYb8I;C4(;MJ^B+1dJG-cI
KA+MBQUeZ^R5dIabR(^<5I6<?+R7-)KXZ##4A_K3BUEAZBM5AQg523HS+^J9L?;I
QW#[9)5?N+;F<4;5D/cNb+16g+29WX^]H>FK[QN^;^W4CTJ2T:24OX,D6(<]7&/c
9dLFWQTAP<NTG8U?41A;HMIc&Z;I0)VC)E\f-_b4.eJ_E/>=]&)5<5>4F-F>&O.O
A3NNT\bfPbRa<K>8I,SbBCJ81E&7ZAO:J8d=R8<YYaU944.6GeS@1Fe0DSO08.7=
N^_f,.>;-^7BXf?g,IHO&Z>1U2XDGY^_P;cV-KfHW]G<a.[I2G=dfNO?QF=c7#C\
<6.-dZZDObM?0S<&a,BQ5K4bB5#6DZW1C]PY&,1VWL7-Fa\^_d_VN);#]MG3/A38
.7ZO.0^HC(^W:Qga8\M(\2Q6:BgI@<K2HXN<QM\V8#L3?89@_DNeQ)b=2P8?cXMN
g1[[8[W09MdY&./+c]+FIS;=^D.V&@.>-PHTTgd32WQ7bDR-bfX)I)J,T;=QW[_Z
#-;bB@-b;beUT5K<g)3>IPJX5=(+^/B=N4WXb&@bN15CD^=4H(Q3+,[Q:A_fFI3W
T2TN>_,/:TdbO)FE;,ZK@2#1F?=#;ZUHMbCIH@DHXL7,D^I:5-#MJ.G\A8d_A9/8
OdF5,MPEHQ=N1GNeK07N?M(OIRO&&JM]=Xc[F<+dCB1-g.VHV?CE0PZ1TB<Y=<A&
Q16\2:H]aV50@KVdJBF[XM8d:WSfMN=@I=-FFbg3]-](4I/LN\#2.VHY>OXcc<](
.D/c/9)fcc0G?U662_^#4J(:HSD<][<C)gMXZBf,#__RKWcBQ[PCP(&X3Ae=_U4c
LW#FOHIT+1Yag[;M[fO(Gf4V4=9K-5CURdURU^3g:a(GNEa5M.,8Z-X]\:D.CP67
[b^/UY/,=d+_H&]ZP>Q0&1<ff[4U;dBVY0T@3:EM7]FVMbW85Ca9J>c&V9.&JBU7
d=]c[.+9eF?LHQ@a\OMW2=,5&Z@]GPD4a?I[V[eHcR)F>_6\S6GTg\R^A-O_&5B,
S@8<6IO\JLeT/_N?UR;GMEY9X079L.ZM6]@?N:MLd,^4ZOT4;2a,XD?G-&A+SPe<
bM>&?DW#1]T<g=-acQRP,ba_3SZGY:W\M=Y7:Z/27<<e0e4Za36U]<(L,183SCeM
LW_c,.bG-#Xb_eK51O1QH1+AZ9#T/-6IWI8Pe<Y9?3C2<Td,4aL&FZI-]E@3gJ>)
^2\II0HGUQ6Z7&O\R7+O3HF^4<@K=]X9d5IK^A19d&ANN-3)JR:Y&QB1[UZW)TKJ
c):6,TT_NC6)_-GI9F9R9BdWSIS\/c-JFeJWbQ^IK^EHT<;H2:0-F[^-MT\DZX26
RegNBbYgQfPT?)\O=3?=K#Z0.D5V5F0Y5W&(V385]eTVLIC#HR)WH6XH9Q(MDA?a
BbP9FW,E?)D[KO=?@I/GZCLDc15EU=5O3YJYO5SXf>EV--gUVg+BMaJRc;c[BO0R
F/+ST[&-9Qb6^M:_U7=UZd.-0&(eb-_S._TU66bC?LUW-]-cN]_MWP_SHH^ZbRRa
Q+d8H?PDAVGab4X<Ac,E@M1:LU4WaPQ#_Qb>&dDR;<H8:B)[5C7[WDFF3cRU5#WY
)(]=E+@MQMHRJ-(Id,1+B_LRM30Cf7X,aO&Y<GK[JJ#[NW@JZ9E;dS9.9fETQ#FU
#^FK5Q:J<S04ce&F64NVf-KH.4I)EeaX363<KI-2B,gS2[M_0HP(4GdZZ,dQ^;,2
IR#F1YYLHNXX_f;<IR^F1=?EL)ST:O&c^::62e+)6dfVDMcU\Xc?;R_LVb6QOGgd
862Rf0TC^X5RKDM<Ed3c\QD>E]+4Mb//<^.2]#0D+Fa?RW&GW,J7X8)Y&UTB;>d<
_2LJ0/T,f2+H]7cQ;R&P(QT[OL.16&U[0Q>C2gO3/4Q5#@[#@DS+YIKRY\YfK6?_
UT^=/9R.4/QHAT.[7=-ge)BcbI@^#M3Y5KdCFF(1\CP]Qc:?(fFQH^=(I=W:Z0R9
Y[MCA)LAfP2K29,)9#d)5)EOOVWC7>:0=K[[S(6[?K=_JN,9^NbSa<(^f4]1AIC:
R>0:NR)(W)>N;g2,fZMF&[-4gFOTAYPA+@F[9IIYADJ?1YQB4\=#eCUTecYO-Xa1
U7S;^D-ded8T>,BM5W=7S7dQfA7;>G)dY5M&,/=9FEL+0e^:_H6-XSW4JCQ^aJPd
A[DY4#)<Y7]?Q&aKV^83I2e)(U9>R-(.(BO0,S(@REW=fU)Y>/>RGJFf[7O(;2g2
(ZVA6ZBU,bSfB++LL2\)TB;a;/:=C8P_@DTIXW>gdf/P+JG]C7@S3<.ZP8#e8(fE
K^U,>L7Hc11cT_-MR&C1TfDY9SE,+eO=bCg,,:+FI7_L@2ST9XZV9+8X9..79]bg
D7:/M0&A=Pe\R#SGD;c2N<Z4EK7[a8DW[4:Q9W[]#g<#EWf@-&#,-ce/]K6H&V3]
07\UGR.^FefSTNY#D@L]8CW=P[UI=-Aa1AG.^T1?3\8U5S<,D\6O(2A85Tb#[D&N
&GJ8&^AIBRe1+dRZT<<CL30f+JFYb)CceJDW=NNHREA6bg.K(gSV_C^Z&@/&X(<V
JA/WO(#cS[P-b(2:\OAEDBMe]B<7^4)Aa0b2eJf7K[7@5DPb+6Jg8&D;7d/18K7.
E[7;bfUdZ9Q4/^NGO0C==G1@95->?S<De;:LOCE,T(?NCY<c?:O(fD?V<7U<g73&
J5BZ-4ONdWGODZ2GOW9]S_77Fa/K-5ICP,Q\Q^DNRN[#5SBB8/NC,?c]?Rc)/G=L
@]EGT@>ggLI35Y>#Ud#;M=AeU.Z@SC)FN7@)3_G-MaLW0Z)=/a..P-R<VT3?[3]c
g0#-&,(G/-G,Ge>,c?CG_6K@c68;<H8eN;GM?aW;5^]FB18WbA(FL<V(eKa,b=8F
(<A^,_J&&^698?Mb4.Da2Q>3L#f@&5]BOFQ@0ZP3\/Q;g=CIeK@b:9EY7=Z;#S;;
3P#BS9-P2b=J(G9.\C@cMFX+R?HM/6,S_2\W^[Idd3:58G#3+F?O@)#83WF0L_WF
X=?_Qf9#^DYP+[4F#-<65fPHZ/>F(7Y]9dP7d<+NSIP#X5b&R)dFKR(9KRbf?IdI
;5V^MBL=d^7^/?^=YF::&G^d0;TPQKKbE&g<7U6[Md@c>YdQa.dCELH+K+^)L3G[
18A/.M]<==IZAO^M&B01?c8T^Ib@G<Zd5P4HZ9)?L_6Y=6c__#bV>@(]USS2aJ&4
M?0+?#ZMI8#(gb<::??faabLCWe2e6d=535IRY2/dH]C4A56;W5E<=YXbH6dH1,-
,@=.A6QV&[#>CNQDg[XHX:7-4B2O&0beeV[?f1)MIR7Dc:+J(SA]J,7a](ICF=dL
,2)YO^B9,A]FK[G,+2OJJ[TK@^aY=#4M65ReD89OFC__A:YQ-.T3gLV:0(4bE(Rf
YN>e\aWDQXZG2SJ4,Q_8cS@A#>(WGA>?>H#EgX,@cPJ<8WZ<[R\U0P@E&Td1-ecK
M?=3bGAEa<?@U6Af1K[YE3FC5A2Ff8[CTZ>]IMY7c;80=7cOWEW>.XGII(2\OI>\
bdgMZ/]@b0K#KWC(+)7IPA?(A9ac3d;eB-LS?)04cg@SKZCW-1ebU_c4FRANBa/_
7MJdYQ+GKg-#:E&cT(SAEVef.fGS2QQ]a>5ZZfC.;,b3[4GK/IP#^)-_XLVfF#U,
NN@4g&3DU/;cGJU.G\J>@=L)fHD#(KN.g_b)[&_JJfV5Q+(PfY[2YW<Ia[Ef2:T3
GeCEJIfLJQ)>HCHACRF_]EZO+b8f-ePWAS_U+]YKGU\,-NB9KAUM6#4RF;FF>#:-
EOR(DV>QWDd9@LXe<C6<<USCSY@5Q,WI?_A(0G#&2B23;;/ae^QT>6PZ14eBG[T[
:+WAY=.M#9H[IEH;J7IY:FUc]aPdJ5+79&88B\[b3MKSR^,#d+2fe^GObaZQR96+
=O&bY?eD:((Za6#T9YPB7P-1WK-=B8gU:e+TR[#M1;H\?N5gES.<d#F2L=f4e2b@
LDK&Za-#D1U0_b3&-8.@W_JI^Ae#H;OAH0X<g[PHc(H=P&,H3/cDdFDaZV5FDgH5
@#TS]R+d36X#Q;G1BRDL2KBC[GCT3N;R?DYQH<@+)Og-6J,OTbFD,d0=Q<5;=WTK
(D+L\fZ7-U0B]\9\X9E@^B(4BX+B2BX]F03+?]O4JSfcF),Xd_g?=6HLNEO09T_8
+7)W,)fb0YE_BMZWJU7Z>091SB56L@4FU]J-XU])P/[9S;EXSRfK(2H5XU7Rc4.1
NYg5-6N3NgC)<bZ#ALZa)^EbOHC)Y(L9dAO+)V,C_U</2:db41W^9R9-Y\R7+B<_
f>Z+0SabGNeIHa]TR5+4DJaJP0b+\8c_:?IOYGSe[<[4]78,KC#/f)];78_&YHVV
\0GDP]Z@Z5]0,gB:=1CVMQ,TH;]@]&.\>g[X+f;U,_?KaRQEe>MH0LS>5H)DU])5
+:,.YH(B[<B98^)HS\-=B8HU-A5(b^T]?PSYId&?@Q7-(eMG];Q]?WWV5R[FL0IT
A2#/cTTEBReR[>b?:\LI2G/(:?NA__BcT4GZS[#N<&Tde6faXNgdUK\GI63KCJCL
19\^U(YNGYg30cI:0Y&GO#ZbV([=CDRH)#)JcY,&-+:(P^Z/PaaafQd#0J@&1D>6
(BBR77.F(Uc1FHA4GJPcRPSQ;U>aEHRT+[b3EL,A-JA1E.-C&&W23GELE0X;\E4M
_IQ+A&bPX;\CC#R^(I1TRC,FJ02YKJD[NKA/A/M)da1FR2D0Gc@PFb,..bLCCORb
g_<U.<X(3,D3d_PZ3.C7OZILg:?34IeD+77g7G8c8#(K84<=PA1dcMa+]TU[_#:V
d5PeYR:W(g_L:5f)C5cCSF]H4OODJM84U.:7.8Y&O:DW[<)dYN<2)B3+_R9+Y>^F
c]bSHXJ:a:=JZ=2UD-&OH.c6J(KMS2cO3A&-Yd^Z,H/g1Z_LG[5/=[.EZaW7\))+
/6YLM?SV_DJT,THNHN,b]\RZ#;B(OO;Y4#I^JO,^d=8eXS@\cHL_:bH[]I.X3:\X
3@[LS8E8:<5+3J[W[6&]>1e^MgQ&&3I/UecH;;=Y.SR)OM1[;K;PQJPg\+9?A?BY
.APSgYSK<(D:WX6JG><7(4]51PU8P1dBB8fbd.:c<+;6@&#Sd))[JXegH=a=?A,7
9<Pb.3c>&;TQ(L5^EQP(RNPE3NN]dJJDa1&-X<\4f1(EI[_&#(a#(/_W1#75M)fQ
V)Q[NNc(_+5#:I&=ICD<,3aeY&<F+bRA>YR11072eWXZCSgX;VE&ZJPRXTTUbB6.
EF_)<=4C[6FN;+BC1VcI/c)4BKf/4^JB(eAVM87XU?Z<AXS<,J]5S^A\.?RTYd@0
GS\>V#Z;.46=S=K5VA@>=a8OJRU#T+ge9Xd(,dZ-7)VW)UB49FcY_PALcLaRe.-b
4H[H//J/bAdDLKNKdE2^(C6@E<X8cSO;,#,]Q\RdSDY#.L=9R8?aGT7F7^gOCI#E
D[_D?fE##cECGc<4BOL,gLMJ#KYYMbcK-;>8-b;53P/CCGF\(1;>A]<]S>;6+e[N
HKF7b7b/4>^JD)fSd/D:7:<3W\MHgAE8^CG57S5.[8MP9IPELB0TR1<f=MTE28:Q
M(Y0R0+)J5W#JQ<OM0M3d1/HB:.DUfe?-2d2&f)P_]bJ_dK08fNCFWMT&5bN.c1M
8^YA]@Q/YEUBH,WW+@O>^JQBSD=95)c>e<PG#7(:),TcE2E3I^bHf.(gfUb0.LBZ
b-TM.<(?I#:7gc.e5B#bP?0JG2>AK5UaLYF?UGLS8D]=g&O&5.ag]HPfbC:R<.20
/5:E7^XY0gH/;(#_O?<H38J.@_.IKW;;#?=/Oc-+\<4^W/D6J/a>;4&Ug#O^-a:[
RFL9?DWBC93L9eRH_U5d)F?)UNDMaR4^K+@9]1e^_JV=S4B=/_c0T+7g4[)#@85>
F29M^4[(g8(9H75F[8[<]bZ-:52BOC(c3DOZ>f(g8@AcZdNFUCg)Q_bg?HRHT9:c
K4A+N?L,T3FA.?54QW(Ma:D_X1K0FHT<E=4>5c8V,X[57)GF_0QWHZJfIPHTGc>[
fVLXeL0XM[A6eJN>g=P3@1a,,X/O9AXVd]@LU<dW4&gGdAZS:.UeIfE?Z8b4ePe=
dV&X@;a2Y8HUZ=&WKGQMdB,SQHIE2,5;FafMbAC537LY.fCe8aG&:IZDDA(QT,C<
?<2@&)BZMP7.XO>=bA[/eR;g6gL68\??d\U<(WW+?]^G[H;8f\_^H:KZ+6dKJOMg
\QD4&,:b:-^UGYA7I(c8A_7H5KUdV\.?^6[L0VOWMH?fXb+5.db^BXOd]VY7K_9c
7_N78GL.90RdX]/;POQVFS?DVKeK/+1<NW9\85KN>N5([eKLYJ[N+<QfAK6J&B69
:Q0X>U)gY-X/^0U^YL1^L&M+2,O;++4@CCJG4)\Q]M,PPBbN34b3^<4[.[/LJXWY
d904)0<9,:C[M//B?#d6S\3G1/4AeT#16KW@aG]b/J49(M0K<::7&KYMCQVF8HKD
AR<BGRG>+fL5.84HVe_0+E(:<B;K\_-(+EKS1I\JeBY686Y.VVTA8)VP:8Pd\6/F
6[c@=EMI@P_Uc^c8YZGB-b@=ILbSF,129ga(6JVYG_KLg4JWH2cEaNcWF+T3&TU<
bDKd63Z9@80&(O4O]1Q/b^[F5E/DUXK)-HV:+WR[dR5S.acb#O/_O(a#\&c5eRGg
a?G:(ZX@S42g+MaX30f9\Q-CgaKV8IL@f\F.(0&RTefCeB380,V8I54#2^b]PILL
Z40@g5FZd_7fDKOW7G<YSSd^8P:X97aF;36P7;NVNFNC(;=Z@0]][2?gfD+W1F,2
Z8QW^QE:]8Sg1V-3DLVQb8@)3@U3\-3PU(#(1\eW2#=JV=+I-d6MYX^8)WG68g,L
X?NK#[J.Gc&\f)XL,<9D7O\=dE5S<C<&CPHEc@CI>/60B[XZIeC?4-[-WNba-PM[
efC/D[aR?V?@?a;H\I-;]:1P[&A,477#9_Sb8+310WK_K?6EBTB3]IO[<K4@;BHR
()dK9Z?#6;P&(G55=dMPADK)#W)1MI4(6K=Rb?-a_QU5ILC=.[NQb4b//d>])^-@
\WW0;I(fU.I<-3:TA[>^ETPcF:I>,aKSHTF=.]X(4<V<CcN37DIE,-](2J+>132K
a9-C:E?I7&<5gIIgY922Y0PRfA2#_MN.KBW,SDgf5OD^^@2/W?E\_SPF=A0=#ER(
BTC@K>@P)=_&P>57(U=3KF^_I>(f#E+ZEF_Zg+S5VHI:@&g^0TC,/E=5LHSC(SZU
:5UA(b=Vd1?U7<3UMa+M>eDD5O(VY:HVgI<&#DPT.Y<e=<B#:<D:g._[1#EZKG.U
/BBY_79Bb6@T7>a=_8TF\O?PA<H38O+QRKE1bXX@W-)26QBR2Z#\4T+F^>SM]X@A
0(>[_J2638+6da<IJ1ZG:NZAX-QL/J<d1S^_S4+-gOO+9EI30HKa/WY);WL-(QK2
bBA\0IT<#aKSYO@:_a26\@S:^8+;&E;0TC_]aSc6/?M5g\3=F?2Ka@K(5Ac5/4D>
I)W:aA0N@S5YH_b-A46(_,G)S9Q5f+RRR:FRNFNY3I._NZ00Xg27U5H?>a>g/fVU
<C-Ra-dT;;E?E<P8gEO,(&\-]1#GMW?K4&OQX57Yg224.5H1c^gRD-9gMJ8dDS7E
;@TZD_-O.d/MU6KP_>IUdg6E)H8ON]cGL>\YG2S8_^98N[K?9bU>5eXIC@W3fG9;
GEedb]OCZ44T)TQFYcVHW-FALDG=,#e>DgA&S/3F#V7TFA2cTRONfGGVPaHH572=
UR?c^UK-ZB_,JNXMX:YBA#))UEBUa]LQ_0WWC/G#N#JXeO#^Xfd6_@G;&LZ>Ib0@
=/feDS/4bZYQ-78<&R8A(UYK=V?MQ=K+]?(MI][>K7_RP7#6I2@d^=Z/+aTCTV>\
d7JG:3d8TgUU-/IJ+;V36RHbfWWAbY8X-GP^#3f9LX6CR>Q.3\Zb56Z0GN(,#]BN
\\^Rb+ZZVXL3f_ULH,AcWLfS-ga<Hc)07_Sf1L^Jb)/\F^C]77),SC.CKR\MCUf)
DOYMB.C^JeT.\JMecb3DSVW2JP(4:GPBKP)4F9KAf-AB5VcJ5GJ4,M4-_=\1+65#
bfSF)N\FKTKLe;>W&(W)N9/V6Yf\I#T23O8S0A?MRc;L<R\HN-<=1Z?gC6\OGDNc
L,0>=?Y8SFD?I@4MUJI_DXZ-ER0V697I9L(5IA>a1Y+U)X?..(IcQ4,a,289_H05
,?:VDfASb_U<>&8==H,DD]<ca40C54_TSZ14f2ZV]7U^>R.S^AK)QP:dUDBW^78)
EgGIa-fe4H/5-Y7^aQ\?T:6(R:Z_cZ]1MQQG:]X:\gD\J=[1?c2g;:)Rc2Mfe9We
&F+NJ7KX:I-/c8]CG.UGIdMJ#]9e.)01X4<I^/?>,K3RB75K/>YY(O:R?P/75T6K
#X<1>PV;SM[_MSHQ6_Z([(_JYHPZ2Y.++(Kf;/IdQ.;SaKg<R9HTB_[#B+ggDUZ7
Z-6B+](9V_V(AbEYIgYN/=?@U-\=D=.Q,&E,=I4WT=T)EP5ZZ75#dgf#9ZB+9a.7
@TDVKRXFH>gF78RDZ0V\JR9ISV0B-aN/G2SgF=@NEWNC/K/#T7O+\Bc)[,g.Sg<U
_cI1X]7f(O3ACD-BIQ1]OD,/K,OMHYIeNd=/@a,f.ODN-,8BfI([_&?03)CJ0Qab
>UU8M7PD[?F@;Y<+FgRMLfB0+S:IO^ag>.>(@:6NBI,9_OK1cG14S5I.PMFKW(P(
8/)#1\\<DD)=cYa:,]DC99Eac<.cTL9-<+TLG?d=O=?9E2_aN],c_e&2CO<[WcO+
7beF#g,5=55P?aHK,RBG:)>f88//d+K0F3-X0&[N0e#//M<[+P;g..,HS\9GRR3d
^<J1bQ[LNTD+P1dP(A3XCI#.6YB89I2_;[,&4JdMcY(dZD/fSe(J(GUc:Y&Pe[#Z
QDY9T7eWe8c:F:/gRGV\HMK=+O(Y@+,&=GB9;14.7-IaZa;=1AePZW=)-V-cT53@
DbNZ-Ka#UKf<:@;8_C044:5ZRFH>=;.<TYY6U.a1]@FB1@MQeKJ/Jg[994B_\Y/A
4K1dUF:JeT#9gd)B3(J0+O2\LHL33#4&?&cf7#<9Y8Y.PT72WGVALMIfP5P[C]6e
F^YD?:8E5CNL(,?Xe=T+g2D7#+U_=J4g\g-d\<516-2V,6QL^,:/-/IKX(AA;f<3
ATeR0(:A1[):#,.R82]#/;d=c;Y:7RA;,(E?=LI5LU&Xg82(HLAZ+T8;gL6S=MXP
2ZeaY\0.M:6LBYYbMSN1SX(&G4=LR4VMCK9JF\Qg(RHLDNI(^@[;DJ^)]U+=2\;2
+MeT^#^C\/U/fY[bUHa(8c>]L7^W2ScAF/K^,X]G^51]a[Z<=PP&[:P?-8T<Y,)&
0806GdW/4^\Q-X>9^X+N]X6/<HA+R6M0P10KR&UO.;eU<L6H;1FL[d=_B:VSB;\d
1W93WTa;g4Z3Vb5&SL=[GB^GN<cJZ7>O/554aaXgfg>a^eG=#7R-)3RecF8.40J:
^Y+_ATT/J53MD+.f86P4)7BH_9AEYVP-eFN-MeD=+TSDM#)8UMEfUXZQ_Qb_7X;S
a^#g3b&Df>:N,6Q)\>@:OZ#0(JY5QG,/e_MOQ^P_?)L\Tb;Q)MH>M3MH8\44#Jc,
+&99I?e8WCRJe#KF<@Y:]>Uc]4?U/,?DIc0KG/cRdfUC-b,D.G.GNfMeDd<RN2d^
Ud+g/V:Pd6A[B9S=I++5=/Q<PW-)_ZL>b60,IQb\-[]M/SA3O=Qb)ebQ(@F#2g<A
V/I0WQGT1:H.>DWQJ/QaSJ1LPIF&6?KU&,eB)VY.?\1f8]+F<FQ(&9[^>KGA^ZZ2
>VNeRL5LABE@ScNHB?@dDPN@.>BCdEaHg.+E]&(2eDSZNW;/E]bMD=_W1._GY.I/
V<b&HS.Yd(N22gOPa:g1T&1,-:)bQR-6/cge1gFe>+.[Z.NOVdKOgM0F??]5a[;B
d_0=]SNH^\N)SU9Qc[,85_YI4@)PLH5SK5?G=XP?g8Sf7,Y<\gdg,H-L@e4>Y@<T
94OP-Q7,DC;BKP;LQ8ZA,Z@RA.)N>(#O3X]\+P[V][D<)&TN9L^LIcG3Q<\[\0a8
?L+.IefST(1Y2E[YCeU/9,7L8Q946J#[BLf-@Ua8VXNY^DEB^.:;))NC8R#4)17;
_Q6F]J@L;acF(YJM,/0Zb\W9YWHd<Z(WK=g[b\LaMZJ,[C&TKfTL\D?1OBYYD)3F
6Z0WgA^D[#9#/MVGc]>4.D5Y=/9&TF)bXBAXDHO8Bg2<K5e/]V6?=QA#OBTR8MGH
R:GUY<\68_M-+.G/8ORW<#6E>@;+]Y)g<XK4S/>W+TCHK:@MP:7_=XIDD+bT=C>&
HG>DF6392O3P?.Oe5,2?;cDVB-9FWU-/H_-2N&0N,WFK\b6c42N@_@ff:-d-;Y9T
bELCOURgI&UV=KC>E]\La@DUT1MWS3+52S[-QND__I)2fH^4UKd2G^S3aaK/M0&8
#a,+.;Z>Q;9^fMH_g]cWPaT-OdH\0L(R9Mg9eAJ>aVPfK+c6LM+25Kdf,^QE_d4_
aeca_A9a>>@YIO?1VYQ:6QRY^]b#,+CA2KM92>OQAe;EROd&c/V/[0^)0^#XUa=J
FeHYgR\U<T/QWB<,1+;E9-GT.#6J?AV[;A,&&1:/dZJ4L-FY&FU&1BK5>R89gA]U
LMgL\8?Q<X\+/UQLc/1b<AO]CcT4?\:E-O3fcKA0[8>:f<[EJ>EU?@XTe7L[+SXB
Z5BFGEBbB7Ocg>AFN0f42R92\5/_L]a>J?C(C&B[IEgfB+58df6Pd8.[NeF7>IH0
ZecB,U]4)&_J,Kc39fWL8;ASFP7WHd&3e@b2+S6G4[gWSbI4>fBcfb02R@];@Y\H
(=OFTS#</FCfX-RP#0KF5bG]#8UAV:LQUOE7gY:b\3fQ1SU0YEE8)DD(E#)RXA#^
GE<^Y21K7?#A+eW+[C6_/,cCKU3+BRPIP?;I<TW3-DB=)_>3,QA\)@0f#1b(.3]C
X9Y<-78>58@3VUN]PeKY-QSUcFZfB-I@14a2D)S<P>&;DZCK\S(05:J.5(/SZL<R
fXQF><+U8<^cc2YTGI\1,T[g/E6&8;6<9MAR8#/ba?9=_]Y:,d\N&fM.[T8&@?5Y
X:eDbGFK:2eY_NQ=8-V03&<N;#573Y[bWd@[N6VJ/AC/b,#4B2HE#S1=_OXRU\92
[?YeEWEa7_UJaH,L6]E)GYgd71b/#1-A^JZ(J-(\6&dNCGG&G(a/a&d_QFI&W(X)
AbS?K\]HV2/JK.:QOZQ46N_+V=MLE,8agb>eBf/HCG.93SHD1aHJ-^8QHc+#]bcg
T7CKJ1J\8aUG#e4DR60#@,0TXYAC)Ea+eT,D;8@BPe.9R1W4c-8A&f;2FLf]3FRc
H3@Ra5YCE&+8<@F@g:+._a&:P:19)-aM1fVR9A]D4;+[0&M,I:eTFT3YA&678)S_
<Q[XY:,<QV+-&)UK\OUSJ9b=L?TJS5JL2d)^,>Gd8W]_[4-4E:W[AR7cUOB2Z&XN
X\YQ:&3eM#(Cb27OcP_>#F/M&CR9D@6Z)9L8Fb2YT6<&d+,1_RJTV9Z=7WJ=.,,B
Q9e/@cE_40?ce:740^G5F6H,e@?RT4:+S]?Tc60>7QRb#;>71^Ef(2P,-FA6N5>@
0/0=[M[IH[IXaJ<\)ZVdS,@.>Z6Da_H=^fOXR[Rd_Pc0,?-KL-K(:558aa49_FRd
bONcbOGYXZBeUF][5d/?1WN7bU0cLgVU6<C49LgIRA7N[WH(CcR(BbGbY\U(THS9
_:dcOcIJ2(gKI1+<IKB:@))D5gB/(&DR,.193I5]QLCcR\4-dR60R,8[P]edC7^\
XDSe^)N8X1[U1b])]bJg3-)NEC[>-<PIe\9+06V@LQ3BLHcC=(F=IB1ARDB&>dR3
\3(LEfMSe@@ZSd)E>[&DY3IBcOe\cG,S?^QS&aO4J@KgQDL&a[E327^F7J_8abcH
O6<@1PY5SgXNM\1)WgK-AL:P:>;1X:\VdTJ@+Y:6QZ#UB@&N=[FH-7E]+-bI==(\
0<(LX6J-E,_S>SKCO4>b-0(2A86HE8N?N]bP,E^MM;;S(Z3_W)0?f;5<=@D<MgUZ
3e-@:YDI_92;3-g];9RdHU/>&&>M&MGWI&KWd1ZG<af97=R&8@?3>c?SK]Y?ULF<
cNX;JCDb5#>5,9<^6gaL\cd9eX\G2CY+C>3#=[[4g&Q;:B#5AH=QO,Z[_?gO([SW
8&D:K=Q7X_1^.:2VPUX6.??+H3M#>V5KX.@f:2FO,UA)BN;RW[ZZ/#[^H@OIB+c5
8ZO6.-V5JJ?@#bTe0A/cD-&8@96)Lc;KT6D73aXP>E=XMYCX0>4DB;B\(DAJ<<2K
\2gG7/g.4+KQ+E5&981c\7NW;P8]0f#VCK.f7A)RXA6-OQ3&B5KSM4=U)(?GGAS1
gWAUYE2RNM]./75C6W,\)>JJ^?D0H(ID936+V@G9Dg[YE8;SdD,_P>L#Ma)g]P,]
NCBI[R,COH<_3UGQ<T-+-3?2E8W4QPDCf8\EFAM;Rf1X@1b<K1K@a/+&C[+/NG@(
MX.+F^<gR;<F+b3e,.WU./@VG\g[)^gBDc+LEG,28M\5db;[e<,0@@\bJPL)EDS-
?7BXO?GY6AdPeTT3ed/[\U^8IB(@[8^#b66cT;#JLSXdD)_;CRG,&Fe2A.T0)TWe
BcZ/BQHK,>/[fDEZb<e4g[1<]gY2]3--b^_bUFJC5BN_gDY>HY@E283\GT:-c8A/
ST59^&.]Va([,BOMI^&70BPWGLEY-aRBI.D)HA)Q1L#NIefb,4GgfOC>)GbTOLEb
UH_gV3X6?J.:\V_a?()]YMMAD_6<3Dg[81d/M\91SFF^DQWe7A/X\BVGW)Hg;K5[
K?b<g<,\Y^PMcK]UG,g+]A&cQ6L-L;)MS9@bRYAP[?0)M(LfD<1fdT;5+2:(:11M
gHAM\g\9H3f5NND_3Qf\;cU&X@gL]^]E8CWK+^N5Y&18H@Tbf1<3X,He#g4fRXbF
SB9[CbUf1ZS&HKJ@=AGeD1JaWdJ/8S_YC@Y60+LS[#T4eAMD@(?UIBe^:SOCVAHF
XSXUBSG,ff=B)C2D2Q=B9JZZVHbXagU.edZN4#Z>=^R96:g:-E2g6T_7RHFf0W69
18J[BOc>93+I5/3#a2EP&_BS)?Feg4Z<4XI-:/F-PKSTDR.\^X?1/_Uf+C&S8W0_
3D>b=MXcPg+#\BX_-:VeT/H+aIKZN)c>30RG;83[Xa6WHC@ULa0OF[4VT1HdR9QL
HP3,_GTS-cgCafH),gf7MB3E#0(K-S8_T_?>8BNaZ/c/(b:9E&4/#H7VW+GGX^B+
8NECC)PPZI;<@]&cHA@-@_5c+A?AM.,R/42BeeJfE#[YT5eQPG3N5dAYE9H05L4)
PUDaSYK:#dMU,GLfb87\O2cQ)08)Gc5@gfce3T61B6Q.@2?9fI^8Wa@X#[_63]=,
61IfS?#UJ=L/,I0:.(.[ND\H6G\(68V_^G6VgCCOUSNTD8J88=IO8;(<(S0;-WeB
HM4gbIg&5+=VPZG.V,<FAbbM^5#?@<YL7D>a0PEZeU0YV0F9?P6XX),9Y[.R;MHL
XUN#7g@]5/?B6A,B?KfXDMQF8CBLD>P;;3OKG_dA(?@--Q+IQJJ_,K<@\f.B+g7-
eGea5B\5D:-R^.8,DPZ]GO9cfac^1_HE1QEC1W5W?&-JD6DAAVMg7L2HE2BLS.>\
PBXI;JZ4[TXE^JR?bf&<59<9]@-AE>-?D8c/691O.X,\VH91GR4HIJIHd8]NBT#[
XE\.OJb)J-gS(AU\(JeK>ef#X>T:K4P^<8b<VJ^](^J6)CL>J01,(Ve>;N;29b[Z
(4?50A6=Y&1:#]T.K4TJ+8#=MeRKKW_Q(0HE07V[>9/WGOcMGWZDf&^6Pa9GGcD8
U5UBB7H1^A+HMBU[N=.eS?JB]DS]@c/aSc2#6X4\M;;6+?)4HMTDQOD&_a)A9#fE
d_H-LMg=ZE),=SY&aa\7.GT2/eG/.H<13WQ(_CZKBfU<U[RJ=W+AT0dK.IaCQ1Df
/KD-O>:2R)a@a,<g2G0S-_B63/1S8[RdVQ+Y2<,]#c>U>:;#b5Z1XBZ<+<C\-9J(
bdJ2DGKg5P9Q>5G@0b?@7;T4+K6>+=W_gg63E<5NTI5]D#M9FN1fagGd^DIGfGLe
5KKPH&CTb6Y1#R3T?f@KYF(()c4?6[S]>A&0?@J]V\R3G&.1)f6MfK\QT#7M\C#T
U<Z]3D6[a&/014@S(aZb[.2c8+6G-3S/&_^Y07T>C5ZMC;81gA5^e(-0)-/W-YKg
f/bZLZB^UBK),025C5T]#Q+]W8-T[+b&+.CLN<FfBI=E^16(DBF42GABH#,3#bP-
^:_RV@D#5GMJY;>E_.9(B2L.ZW\UT=b97:LWS4B&OF;HZEf_:\+2_4H?H@aU9gOJ
3b3XXeZ4[U=,EPA03K_Q=a8I<E.P9c:Gd?4-SF@GXX:W1P;VZ&LM#SD][+R&c5.f
:O=8>RMFbWDg^:(:(H\U/YSc4#RI54^FO(FJ/(/3SL:d:g_&MY][R1YZ1.aQd@V0
U:YPTQU7&FV79GW)\3b+T3Fd;<AMM\&GEA,SO,+E1#9GNP?<_0GfU]c(B24E>(D2
2Ab[39=8-/aPS0/dC\+30bZ+cKBOEPf;+eH:8^J+VRIXd8I.5.S9EYc1\L><J)A#
)MD,EM9K_=^cW-3Wf+BW(7DR;.AR-PA0D##-0<dJCMf3UPYd5M?4eMG\DS@:[2K9
SeB#(fC2g]_4::Y?>fE)]\7L?)_Q4aB9N6=^,e@RfLA#Pcf1g?f3H98NMD0-bE]=
eg<B(N6)T;P^1-\;&MA(UQYcIR<3c67JUa4cRWKX]L))9WL5[^-;C=X3/>/=1>:)
O^g?_Ka,d-],1.JVU4QF(Rb5eRc#3EPA2YD>Of8JOW=[=W5W3]J=NZWDVe<UL]#@
&>dSRfdG5)EB)@J=#WgG=Fec,7R/+Vg3?g-[/<U._>=eaV58#9;\O,P)^)Y44CR4
1A99Y>R8&XQ&-;8=O7IH,CcQFAOH.3+\Y]LHAG1dYI]2>&+M2[gPHNg(M,WKYUIB
ZI7TLI<+B,(G_E@?GODaIFE[C2<5a#Hd3D,[7-eACdHG]BU@E7UIfeK?8Ta&gX8J
<T8LWUN#B,W#d>/TRVW4-c^U)/#&Q+cUCb)YBMPKAU<KZ[?DKKHU8G[bHNXK?A@^
[@)@&WfKcB,<=5AO,b5b<1?d;W;#V-K4[R4aG#(TOK6d]NPe2@>(>UIH-bP<Z(5&
7P:e88>#[P5G4ONXXWc2OWVOY;_]@cf(I611HEFA11a\T0@[b(XF)KN30Wc^PdZ1
JUO):T5W:<#]@?,eNO&LL04V]T.7Z/?Ig1QP<.]gN1)e3b]U1-7>9\;P3W,U)&(B
=G\a#U39;B8]2g=UZ2MN-\EWGDM_O=X@d7M)7@[.^?\8gfF(Y2.[B^TBaIW0.50M
?d];9H8ST)7)XHb;&N@ZU62TE^P@1YVfRX[<PA7219C^OE/DD&QHR52eW_^fdZU(
33ZP\g_-/037A,#KQc7?JZR4@=JPba5WNN^^;c?KLGg)E&TLWKN1#JJH=Ug0bCWF
f6SUG@09bJ<+61KFKa)bfc[eP1.@9+#F2BQZUfN[-)W#.=^/GYQKZ\=VG=_,?1TM
@9=@gfO/@XI@8RP7^GN@-4,AN]e-&Xg=-=W5<S+d:(T+WWM>\Z1d)Fd)8D],JECE
@WUCCe\;4J6#J9IeH29).bPR:J>8=+0YGXKN2G[a><LL3#?/09JQH.HD-?0:9JHB
))^:eMR>TD0fC=:D(/N(ZLVK&5aLOM&)CU[8cc8=34:-O\<AD)E>R?=:TeP,3gEf
XG)=OJLe:YZ_8+<3d3I>HD&C?:SHe79@c@VeF6CbWXWGP,Z4SBVMU/[8_gTfNGV8
a,^)eL3PO\\\)6W_WaA-([NX<cV@R)<F+<QaV;,D/>Ob2K/c5J_;^[Pb]#fc,9EK
MW.H^K?XX]5f:KWG,Z[ea5:9[&J_7YNKHIPTUH&.f,02[,WVY^:-0:[bXY4.d@9^
F60[[/]9;dG21^@2-XCKd?KZKQ6W,L6-.+g-?)1/F([@G[8.b?A(VMJYO[9@GbWe
Z+I2e2I?4A-V7c-M.WWe9c7L1;3=RfN0-_^dNE0)2)(ZWG56;c)RJGD+c;PF:(C+
T>9\/3>PRX,6K/Q?=^C8g)fWdZ7<]&=4gG7EGJ8<Q)4=@H+P9OW4<f>0gDa8H_.M
E1f[aCGRQS@RP/a\bEKHWC1[^[,YNcJH]65WZMgZDT8M61#CP.WRL_59./IR1)L-
0GX\&&W])P<EeB,AX(#,-^Rb[+//KTH;LCZ;9D8?NgCT^:Z>P2TMdDTc.1=^<9[Q
HP#3\RWX=FPU^NREdF(7=BId<JfD1H\3>e#b+61:)9#@S,ee30P^8db.7SfU_U:@
fXKgc,c5N,LbL+K9[KP,72QbAJ:C])E5E\@-_ED[.;+=C2C\J0-6)S&1)TSdS4KM
Q^dZXKHE5DNAdCaEO@;,JS_^e;^DTN3?]SO)H^HA5POW4LR@4NBYI//S\K2d-8+T
NU]f7ZW#C@V1/93SJgJ7VgB[0fN8W/94[_YGZASTT/gUY[eT;,gTP2eBNfHX?;5&
\\cIdVQ&P2<Z<)L--F6aSB((dc9[74>A?1eTOM;,0=T2_F@UO?A5TA_8_V/[ZJO0
>@aZ_S,;RcIa^(H]?c)[+1N>V_SE_^JDF9Y:DIfGYQag,V.ITS0;<>N,OT9LI=Nf
W._P-AbaMDTV+P@(gF0Y3c7GWM4WFd=0^aEAB:HT&1W3SRP[#/[>d2AK?e\)(+YZ
#-26Jde#XCH0g.5>5B4,2652,MT=Y=Q^ba(A(5F:f62dHS0I1SP#XeXQg8]9gKM<
MN0[DWH34H>#]Rd3TAB1RfE&8^HNc#=YN7BJ,(P.#:E+RY=.F<ge(Q83#W,BaEFB
L8aN^_((_[DTEdF;7>W1J>GT]4;6X.g1V:IMcHNbOIH)IcQ9(gU2MU<ddA6WT@AT
#c69U(9/5+(#O=K>gFQNd=FA)LE6Ia=c(,Q-YL:^0&>12L(c5He?dGTRO?fcc^6_
[BV/g7d8&Oc.T=YL?N:cTD0ca>=a=ceGYHbeO6PYPBWKP5+(5<#KE^<1L=:<Z>W,
(SS_QM<T;Sc<B_3/g599=FF\YHE/2=Md;g@F;EJD8^<OL8-G]_SP<Ud+\\E91U^0
KN.Q9d,R41b//,.;DTNHI<gK?Wc7SS_2>bUME6SI#@Q).8-0,B1I4Oe:#0?MfFHV
7K>4;0c#ac?7HL3U:(2&GW>CI7DCM[;Agf,8VGJ#g#8?f(:-<07JGfTWL84dRIJ9
WXZ@<)Zc73aZ=]O0.DF9eRJU[bC[6;91;HN+FESILOb#T^K-b0:2<JN[8,:LE@/7
IU8RUF_XYN/S]_14JQO5<,,UOgE9-@M-4V&4]e1fDE0_,==SfHV\C0f+._D_W)MC
FSg.9,1]_K@^W==^[5:g]U1-f2>/.>Mg(C?=CB5C3\6bAgKd75+4J84+[M>OBcaT
-NFB5,V0cQFb+9be]M50XL4(J:52T2M6_&VT=.BS;e:+;=U<U#P>+0Cd(5N;P\\=
0/b5,0C1.H8T1Z\?bH58H-9\d;NgZ.QU&#6(IJ1C>f\]691P;5QI5@>/I6.K&Hd-
8P47P.b&cR_e5T.ZTC]=9J6/4g80V12@77(=W\_D+TZPJ>3O&(Wd:XM_Z,N4(BQB
O(;#Z4A+6XRCSg&:?N=3@/SZJ)#g[><>[:f6MX\:ggCbDQ-/@4N4f5WTTM:Cgg3X
d=V3>@0IS<F,(f19W:_^Z.TG^JO=<FcM#Q+Maa5X?^Y0bc_3<O,>T:]3.+LY>:;(
F&5e/KMV(YK2FB?IOC]\X@e5WgH)NbE][GO-,8e:(IVSL^S:2PKU6/,W23Z#W00_
728;697B>Aa<_fHOIIFR98_I^Y3?G[7/([KJcA@>M]a5<[6PMf\T:7dO.S7&8Tce
f8S^#HD]F+LF//)W7SgbS1)AN-DLJ<1FQ)XI_eK#S.NZ1>0GV64FgXHHg&C8P^Cb
S:5GR,T@]gIG[R:HS7a:QXL2C^J/FLdX7E/fM,(N>HPQX]<LE8OOA[W6#+9(10Z#
(@@CCf&)?0L.YY2Tf7&>1WZeP<WWD]=XQ3SIFCc)V9FH9,)bW3>99d^S[A&70#_H
:RJCQP4J&J?<^#]0(gC8c71#aO;1LAMP5V0@VfO_HPK;N+U2[WF\[9;5RLf(?>(G
KK/JC;W0MWg8?GI/X#HCLQA66,52D<MET>4H+RX^3D?&DLbHce4>6.@a+M3H97E3
>L/XP52_:]beOM)_Q)fN8D^(<gVaI423geVIb.J(-G64JWB_X#ENaWV\S0;;RIO7
5\5&M8U[TOX>:GcA<B-P8GRJYL23>HGeGN^M@;R79<?/e.cFGHSN.:-YHM:\?IQE
^2=T)Ma^cB,3a6L9O#I-G19dT(:[6WWD^eD5Z\NSa+]]f2[#E6G5HC.Z>>Pa+/b0
LK_(,9G#TGHUK/MBP>3L?DfRHH-[@(I8f0C8WgLNYGTL6M@Cf.c-N=/b[\XJKK.4
b3D:@GBJ;Z]]3bH+R\8TPPD@G^7:@)ISN,&5=>214KX\DASM70U4W_^TP<E\&K8E
Q+0BWU.I5X4^^X2AV7/W&dR&EYYC(Y&b&]Q2Ha7=U-bbf32b/Y<)3)4_1?]F#?AP
@J\a)C/Q,#B9QO<L>>G#VGe6?\6a?DX1TMF,=+CT.A>[YEO9A4EG/8d\O8ZN1T<V
@LY]9EU2C&&MHCG#T/A^@gPd2/&5agNg?K1V)KIA;;WbSTD2I+.ccVC,SNa_G<cX
g^TR7B_H9,7<AK=@^<6KL?D0OL0\@<caFOgEM20Y3R<KOBc?WF^>Yb>X>P,NU(ZP
SXg5R?+@2ZT-BX)Z:c_6>9FWAAS[Z&1GBD?>?L+;R76@=[7?_?KPL]0G7,8/4&_J
.6Q-2AZ@eO2NN#5P;4SM?ATJ9I&/g;9I9;df)@DQ^O><c?5(.Z3ED#e\1K2;HRWS
);6J6=aJ#V60=4gW7bZAWaXgG<ZcaYf=f;O8dNP:)Y=G==,7R+75T&QK(-e6Ag1X
Ya:(5]N>HSYbNEU)IdNA=])CIaKZG-T/bG-+&L5Hf#CLTee\/@W;:^;B#F<N]NT]
.&KCSO=5A66)A+@;>0d5f[ON<6Z>V<0MU;BO/L,3_V,79.?f4/d8L?V,IX=^[&NT
QWUFB8bOM&I8DH7#C#,=\\?Pc=Q=F/<R.?TNd#0I,DAPD3d.3cb8L&Y.;0ET56bZ
_/g[:a.[d^^I:5B0P\(F^<<5_O7_5+g[OcL;PJ[44SB25gYa.;5(gG4c18-WWL^F
O&,R7[L@Q,882HY^aLLIc9SV;aHJ50:RDW4L/R&[J/#5c](XUQ&8>A=06U6S=MCC
f<,Ne),X_7CJZ2YFI42XB]I2YCYC[a8^[[-OO,a9(BAaP:N8G2\ZEO7E(UE,B^TP
d(7Lg.cWbM4#\&0PUA9ULPB)#>E4RaK[P(XM@WLTF7PY-NCY@A-:]X&U-^Qd_.?B
)RDK(Ng:Db.T<^Fg7(H1ITI(P\,GSaDJ:##?/E123g57GA#D?.f57acNH9=[7BL6
5#EZ\UQ^Y_YYI85E+F8:c=CR/+[gD@M\)a&S-S>a,26^LdQ-<FQA842C3D6X&V/,
gP)&\Y01^SM>eK2\5<<U1C(\)eCDTDD0+MWGI7Y/7\aY10KSUfe>04#2B5[/=&;:
@+^dI/_;A;JWfP>c0AM[+K&6DC89+K2G=W.g^8#d2OK:+?L]LFd>C+77Z=g\FGaF
7606;EI<DD[N?RF6RNECFD9X2bIS5/YHceKdVZ8>H+KcFHc5;</(TQ\1>^86YdZe
[B0WUMU[,6#3NMT3_VDV\/;CJ8,I=)0?4=5Qe,LbF)X][@X[T-<.;FL)&+JFReN,
#8A._F<V/L9UT#4<_4afVV]39XcEQ59@ZEL9=+I@JBI;(=fYW5XRC2M8N#<dFNBg
9<c.JG_T>O\0R^BL#69_FDG.XO1F,<N)PAd6SA;B?9a:C5?-O[_\<;TBK]X^[P9<
=f.T:(/(dgcC4^3^CQ#W76<cX2(MfKec_N^a[_@BLe@JQ40;Jg/JM3\N_,T;<ANW
+\7?U_[IU>6.4>YS.5)1DV;Q,#7.c>XRKYd3U2X1\-Rd+Q/:[Qg#c>.[4QT?eLKd
_<YS<NWE51JS3VP41LNRV/RO(5M&_T)8;f<J.;][>6Y7PfcJ,=7e:B1X86cG?(DN
/@.MZ/K_?M.9F69)RVc1B3:0IE9\gPV)JQAK>R[NfU4E@;A@8E^[6008?7AD7=G?
16;fH+SePK,,d,<T4_(ME[DTH:XcceSQK[<egT0Q75^TYNbNXc_g3:Jd^=504B&R
NSC.<c&4aF1@6NW>;5eSJE)@]4d[>gJPX^D];#^ePJ)e[1_4/#_\JQa0J;_;XM7]
Q7Y+AUf4+&JO<^DbA))^B.SObY,&DQ/=;LG(M4[g+Y_VZZTT:1:3g_cTB6U)IMM;
cK@0I[bP:DJfDb^Pg9Ie1H]5G?3AAL(PX8U1:>EfJZXY4)dd(GZYF#SCF=-_DP[7
gHC6K-2D2WOMdZB9MDSU]9KEC?G=dAR#OAScH,QbY^^PE[HYUOca_VJ.bELb#ON8
&gG=?HTRP&A](^N9;QN&=XSB=4c6DO;.CIJ1e4(D2O5?Oa@L[-?8H^a5=&87;>S2
PQ81c>C?63_X)__Cd#]2[;+1.0^HDV]0IAFB31HTFff:8G,2Uf6gPKTW@_QW?KE>
C64+KD\+fX1c4b9MM?Y>JbFA[828/=,GF#Dg>3cNNVJL2=.+0UFKY8=)N1)E.9Ob
e(.f;69.KWMK2Da8TVE/U3[^A@]72;f^b/;CC^X<^YND<Q<Cc6NVQ#>7_=?)-V\-
Q/(e8=IW4?(B4?]M^DPfV3WVH].=(/&__c[g_-MI>4b>8c8>YfO-+d?YD]_]\0,a
IE.F=6N^XP)_g;S1#+&2[3/(eP;a]-D_Y6c+Z_a_ZJ3\?D6d2F0&^(W1@/U1X\A.
3QVR7T)UG(JacIYU;Hg-?9=<4Y?QXF[8C?3^2\=<N;FHZD@834O#?0M]/[H1]:G5
6=b\K+eS,0@ZSeC(#HR&Z/MA_J^C:1HJA8eGJb[Y=3YL\TS5G1.a)@MD#_L(LfN]
;.(4?-0T7L5CLQ.SGOK=+#:J<4<U#WI()D<NE&?7a+9=Ya,/([R>dMZ05725=a,6
8LM0<+W3?[-[.1J:P<09:LOU_,I)<@L[>4DMA[JVC&RG68JM:@R-U@Hg?eUP=J+H
g3ZJL@OMePBV=:4719VYYaF6G<2c,YCMAdEP@b\OK-^2[GNN8US)^d9dDaHZLdJ3
cae(_)8?Bb1&/Od_GG?J@@W4)cBN@UW86KTARQ\99JM#;YDN,d?G#Ke^,D,fWJaT
]:EAeG[RB;Xf5,GJP<Z08EMEdeEY0H?;bcf@N10PGa(K_:Mg3-#6a&4\S37bL4e<
H?;]ZE/A0V5a8Gc[=N]2,^SeK_eVFR4O>gA&L)>M1b&RF_DgX(H)e/:ab2f9HV\5
=XN<=CWf[JTSYBaBeZ=BW,[Q85C_AZ+_E2c/Ac=9K71ZY-.D4?#9/P3Q;gIN.N09
XKUd:#1=RgZRd##g0(X.(cg3IN(H0Fc[XM0a;9?ZQD=B=3FH6CD=6V3O+C&R+/gG
gY+_cT5P>=X,6.K[b_#N50cXO^CZN4@f7a]@&F(E:D2XHeWX?<EeLXX0.@?D<A.L
ODgDU8PI&^,T#gM.CL@W<F#J6:41Z>1)7(5(PA_ZMf0gBKGUEVL1?A4Z[.]?B&Q1
eY-P)1A]TQ]X1QgRFL8EPB70cQOL8eI,efe-Q1X@>b&1=O8Rg=Ha]+YN>Z0MXVf)
C?eHIZSEbZO,Q6YG(QU0&_Wb-<QL1D:UP(;XUE4<P5b(8+?<3\\W:0RT)da/ZALC
.RN[V+SA?Q;1,c6R6D:TED(6L\X7TOP5V&)L7S(&aQ<C^1g3aIee^+f<6.W<K63J
Xea=0gZ\5Q4e-(HBA[,Z6O)8)Z=Ab2)#9Ha_77&1W#bG4.2Z#7(XN1#H4=FgJYHQ
LSHC-PTSfIMe>P\9VN@AZX:P3bBAUP#7FdWG91dIb<)R#PEQ,?S:;&GRYa7ANP<F
/&@@I>D5>(PQAAYebOE:=;5F=D99]:dg/>2fFKcWdNZ+7F+J[D3UC>F6TF-[2A5<
Qb7M@4JA:[V=<2R^.(T3NS.A8dKQF._RPB6313^8,dbaBH)5>BO2DdAcc3J[NeFA
95aDQ]?PJR)1G:43]dC&BN2S?GX(&&[_Q?[]Q.J:=_3\.)H)Z-g-Q\MZB^I+/YGX
_F/3fAf+93D]L,5O_ZVKYT07ae+F_c>gF]C)Vbd@J)Z+3RIC)X2&&FQ2:8>Z:D2g
MZdE2/:\:E85Nb9T]2DgJQ.5>)Ab;794;\0cXZCX2,,8A;I8AQ2->gXB\8dd9\S]
8H00^NdV-3c?WPA^AMd0gaZZY3QN#-&1:?GJb+e4d4[O6B.X>=X5/:WR.?24/F;W
YF+MQVII);WM1(>YNOJOFYM9OWcC@\;J>\<P7R^>PWdWc,1\+FQW-<>1Id]2HO[8
:PV&IL;0#0N8\[3TVW2-Z_NCV..Y-K]P@f0/BESW;#EFe\FF#NK=2FK\93]ed;GC
92?g)CA3>Ia&@CT7.b&0_??BA/JYdE<2\?Ud24=J5FQbH\G03f4Pce:B)WV#Q7I]
^SU+TV(18.)OOR9+4eZV6>0=);NB]TL7N-2J>3N/SZ)8UgU(P=3TN7a<?K;f\&.?
2]A\bKNZPRL.,A#ZZ&E#+4P7GWAXFKM)L&<]L)bF1PFCDY+#0&GJbe3eYX6;ZQ#+
f)B1(dBf@HcJKHVE7WaDITQO0(=5-#cD9gL[[80D/e&3H6:J;gfUd3ZV8BR_@Y:I
O&S^^U.-B/;1=YU-=5F0OeV263N?eT;OE90:8HaBJZ@B2_6W#UT8_@O7#?W@a:,b
R<PM3G923I259+YOf+2ca2O3Q8MY3F7[;5]+P5=e<1(D0._F[Ee&79MA&(&J>:/)
P)?3A\?-gV/+\3@L@80?<QX4D6/Y[0+UE7#W>U__VH1-JG=LF57UH)K6.,SG?8b2
..7F([>#E5/E4(g^V0A[^>3/H95/)e[CR-R(_Y,JV25)d_H98IZ];G:B<K2=G.<7
Kd]XT4EA&LO^;Y(\[RR8XMPARG.e&\;D2b?aO9/H^,E-#,30EV>S-],X>\--g;B^
N8;PWSJJ_A9bRBf/8>LW<Ud:=__X;M7bGH\_W>O9][,MS#20e<[BPFfae3?FYX--
94;2QV3,E^^_&;S/OG]?YR34\0>#N+M<24V9_W6[KVFVcKIU[]-BDH7P2cT0LYH7
fRRB.0Ce,a62ENBe7f_VA8X2_.2DBUgS)\\?.)1I@8=-9g8SJIECD)NMAMRA05;f
M:[2EC2dgbgCW=^aEK)]K@A6/aH6=EH,E0()&cGBHY[+@\F+J/5,e>^bR?XgH0RA
FNYNTU\F=ZE^fcVE+QVc1<=LPaXeaWgeFUDQ/]-;&JA?N22;(eEKFPa,X]IA)8YY
4:Q138O5P2_8[/ed3KBO8D2;TFbf6VI@=8MSXH7HEAWd;?9gQZAM3LKHE]@_/9:;
DYQP0[?F+(B<X#E,bV:9:[-]GPgJX_M9)]JLc>8IF,XG,,BfS<2D8X.AG\ZPEB8a
,@.I<7^+M5ZICY8<T59gJ8J7OJaEC0#>](N3HLb1\7<NZgQ5H4,c;V/+LGGQ@TUe
VNeL>f@?f3dAM5aH^>c:6#+_\SeG7C6E60Wae4@b;d&R;:fP46;R;\@4fWVHfgJ6
3KKTAEI22U:GAC+E>P]L0P\Md5\,1gQ(Ja]QVKD7X:/>^?AIcSVdKQbJ&dHGK8=a
2Q4(\cb/K)fOY:ZI>=AFRBW558K3a9<MH[Xc;Ec2dBc_<GZW=R2(..?+<PY0BOQZ
E_>f+e5[XdS6WXY:fNXV.TB,0Tc7297a;IEUg,7LA=WED6/S4=[OS+T8/<3[)c:;
G>ODNbWPM?&/.a]UQ4.7CDWE<3a-BV^-[LCP=bUSS/ef,F88d+U6&PU1,UG3@?c@
^A3INE#Ta@)&aRHGE6Z_>?fV?F_KYE9baS]EQ3V9LD.^1^AC+4T;.5D+XR&W?a0]
/0eAYZb^P#CD\+>VfP7BV)GLB+(:e;(N,GccfPZ^>=TLaJfI/8V(>,_-PbJd;+0>
P<O#e&^<X?]U&c\;O0[00<7=_6_fTZ.-Q461e0=IZD).Vg1SggdR4g_3FfF3^P9-
6=<dR(M=DRPTREMX&J?I1&&g>SR#d(#/B3fWJZ+e^>HaX:Reb@>V;aF.;UJ0H7^Z
9+R1_\COc]C4AI0R3U&_:0deCS?(+9@1<73Oc\BEg>Y):GSE3-HaD,1:SL.F@_dZ
3^d&+=:9bP&Q.E,.KR?ZIW3A-O3#76]7YFaJfa\]QbNIV?&\QJa<FAY:?D\POafe
ADFf3G.STaVTMMG])LHZ&d9HW#H>+]DUW@&gP\XNaGZDP=Mb46+UPfC1D/(MaAEf
[<,HD+Nfb;(8.S,ZGM4=[CI]HC&cLDA0Y7<217(;IOM5Q?ZX<^P./3XYI.Y_&H(O
ebDbY+dN8DRegJb7.\6KT0\9:DP/GRKZ20\dETC]\J;Hf(F?TaTCWL\HL1G=[_[Z
6:P(U<O5&68W#TgEV/E-6KaA22:RL(aC1XD]4S>G[c(,/+58f-bP=PNCBR\4a.HH
28/-7,,ePK(Q=ebS]>^T^V,Y56-J]<_#d?M3RaR28Ig8b#\YGUVeIKN=RA_.)7,?
+-,PPO[1?e[bD,#LL=F>5_>H7IUa>.9ER,V7K-XYDIG6/^ZGID(/)D#YAfS4P+Pd
2UV@Af5/)=ZdN^B72e0<f5dE,:-cT^[M#e7H1CU.IY9G))DWff3W1X-dSER6K1.[
Y=9C=<[Z;@5Dd7::<FQYFfQ)OUP3Y94^cP2EAHT+_BG,ASa6JY]A/M.e=deWQGL3
&-Ve5,4a2KDe?<b>Kc]f=@@Pd;CBfY7QWMD5cS,FKI8[4=1<?N]JG4Ue[(JG8RAQ
:51LW.3OO8P7^/]G#+50g/gKM44J;KT,U=(FF[;21_)fG_^SE[ZR_NS8O/79I]>.
D91?d,-EQcb;(.(SL]<(\65X6\UU(VQ>HYDH60MDC0VGgUJ8JFT-OF+T;6V(ZJbg
?&bJ43&GdgSOJd;C[7_><VXca?D#[9W^@[eLNYCLUSNdV<R&^S.5>cX.4B[e45aN
,I-FN\Z-_XXEbVFP>C(R)c8b==E#SH/N^d2JKEf]B;:#XZOBV666ZU\KYP__0Wa[
YEI<:G4[4X#;D4WC=&9OT@OQ=Z(+fIc6g&(INLSVb@K8MOgWd0gWSO?JZ[gRIJGC
;[ARgG[6V(VGOZ\MKc(X+F.eI?:S=FD:=IScBJB_d&C]CFN/A;P&1]YL]3Bg3;0)
-JJ[C::XPbPXS4XI24V^&&fD5M<M;VQb)]&)@(M+LO7&;-J5TBU)5[gQ.&PDPa;K
W?EB(-,A+:GH1a>gX^74>D/TAJ]7PV,\HdET7V?RW-Ng?KMAJ27/21J(UX^\F.IP
6f_PW8[V8,a@5a9:FSf+Z=Qe/I1bQV]cAfTBY=9,F><+6,TR(-5QV@^P[V8ab<@d
GZE..e+JB^+ZCJe(Q?-;.DG0K3/1Z6K&)-(IYEa&&EKRfW+Q?.\.,5ERbe])gF>H
P5La-CPU,U<N)[Bfa8)a4;1+JC)T4C5-bXR6cJUeZ4/dHR\(303TOCb:IE5)dB^7
Z0_6Ld:IVRFZI4+1YJcY[WPURdK(b2][D8Ncb:dDdWe82&U[GZUXQ?<S:bK?J]T\
,4HD^NeDP+F#-[cXP;29Vg01d?JB=HXC:.U<_M1U_Ha5WG/CYJ9cL1bG?:,B.f<P
DeWB436VJRL/^D_Cc4CGb#)Y>1^:T>2[aI?8&8VdO,&@a70aO\e2,a<GA4>AG@a2
I]PU&7\?efY#3K,W02-bI#^;88A:)a&-^f._b,)P,<WfO^,^aAB+.DA\B&TLM8Z=
)VJ.Z5;gKLK&b;^?DEU[POEF]NSOFY^P)@(;Qd[4#Z\Q<U,[NI&]-@ARf,gb[]AH
E9[QIR6_RHT\<HDeFC+3ZRfRe&)RXeEE)^Xb&F]-Pb]Z]^Rb);T4dJ40+NTGMA^3
_R65Q+=LI4N_T?bCJ6+,#JGZ).g[>6UD.22755EEH0(W8JS=CS20&#6DMIPgW#LN
,LA-^_6K#&G=S#E9GXFPWU2&W4;GM0J,R.B;N9FBW12[N7/Bf]#MWZ.C:=H<6.W>
WHOKdVSF-PAfdNEH^?,1[FfJ@E8([ARQbR865:30UdK\TFA(0JJ67ZHb@Z@[UU&3
4+Z0ac68M5E>-bX+W/f=2WB@JIYc]MPJTY=3DWM>Uf8e6?UPV#A6V]3Z8YBA52_A
W1;B;]Tc11P^5G,Rb.ffF059b^812e=:X1]-Y0^cLBa.RYHS9/#F-T.96=Td\T9O
EKNUCF,#gXe6#\0Kd<V/Td_9M9?X>)8.e5\REY1@([@=1V>1Q?49+H;/(?KLQPZF
YT)AZ1ga_4[HHH-CD<a<TG:eR^g,d9G_.I)YTS7B+e4.SQ=,Nd&E)HZ[5d8R>ZC+
P^4HL<DK6J6@U8VL;7:IDEO_7>]g^I8Xd3&JVaOA@6E?+;_O26\BM?]L;//)<G6H
eE,?Q[[b2Yd4:)QQ+/C1YHe-.(Z<R8]_[W&<eFg#XGOSb?@UZA<=HRb_FP2CTSD]
6.J(YH3]JXN,IO<X>O>-]OJCf3=(8DeB(<e.UVVEK7SE2g-6;Og-b3W^.0+V25d1
70e\5B/gJXNgXWMP51>?V06eIF/>bO]@:<ZX(Rab5LSE#MSU-&b.PL7>ZMD;Pc@5
SU4+X9Of[K?_L_e&3;U_/08I2UJ/<_\&BCUXK40+H9_W;UY<VXI8M<^O+f@(K3@H
+&/3ROR:YeO-2dOV-=.a49eZEKZD/Q]eRX-E:e_-H0,=IGdI\5.g>)I<R1CKN07/
[,6:cONaD_1aWB5Z57YQ@31@O(8OKX-;U>SYJY\Z6\31,[D+][]NRUe0DdO0VA^S
@FgC^-Y7@#0N#:<d_d:A&b>@Mg&:.KX-FENOZ3&GOLdKf[1[?Pe]KdY+.Q7e61+Z
I5[//X.EO7K^5<4,#BQAW7,HR[#A<F./bA?<(b33APF\QMT.MCG0@T2=gG8OOX?B
0X8YG<4I,O=ITT_?[Z2JdW-]C+WKdW>/b9Y?:UGTMRg=FT(R^NTS=VD<DK>?7Vg>
+P?>_aK,;aQ--3PJ4S1T4N1+49W8:YE(-K##La1(4]6>OA38FMFNVbNCL.<2@WS:
AN&6FWIU:0DP2QT\Zb81PF;2W(A14)KI4,g[(-ecc7aFOV_XG1W7<UG_.S=VJH9)
>4>)K6IbAYG_Af2;J<MC#Re,^#Q@A1eC(\ZB0@CL8T;DZJ@VZ&M)X@F=9bNAK=AO
Hc@KOgZUDg@AYX5+cGO_TM-.3:gBf_8Fe(FQJ?JEN4-Xd(HOAQc+fc+fZ:YK(LbB
IHcW7R-dAG_KB]d(P&9F(A9@MfDWf3A]#ZI:?fPbY@T?BH^9Hf5,4(+W_fSN;VCS
&_c>I9Z_CW;=,DLIDDI]M<GLL_TeQ;Z-=TBY])NZ6=HSRaP@F[BE9aNe2cNaU3,1
D+3]L236X]R7@WF3QK@Y87@M-;X9+NY&X+c4@bFb2/ef))CZCMR+:GS^.0OVVL.B
AMWMYQ07?WXC#(ReaR+4ccZg/HN3ZB@2/@530#c1^-@;?^eF:[Ja,Uf[C+T:BJ_+
C#;I@8[\,AE+A]I/DA&J=eIP-fO5I9#0;P=OJI1=+K4>cA;fG^CgD\dHfLgNBX/T
O?M.&7OLKdU8>NSZC<L>/5)VFLdI;VCg/]R\4[>HCESBJS[2_=\U\&4OWIAXF_(B
[Q/QXe<X//36eQ[TLZ<?:cQ0=-QB4-c^GEZZ>c2_e#9g)^1/(bU@2^Q_L8QG)dX8
##]UJ>)TTDF58--;BH&3@CdCZA(6G;dM.E7U.3RP,/d.:FRJE8+;.Na\5EU&3NY-
GBCH,LaC_551[BXV#H^:BE8J1C_XcDD[(UdWOQ0UO-2T<MXg9+Ub-@Ra80XJE3da
&XcYX7Z3ca1.7.&JgOS3Z+c?-Sg0#_d1L]V5WV?W?56436:HeP6EE6-LEV+ORFKQ
\R?7U,L&0OXSC#@W?,.R+,=3B2^Z(#0R)5Bf:0B0?I81@,N5S):_a8I,UBL?)LWE
HA&L.D:g8I&<^U44:B0_\@\dJZR8ZI3gGa0Cd7^]<VW5T>Ae\5K0(2B2KcLN2PND
XI(T>E7+<cdP<9K:,1/B8gY?a3L8/__\U/.D3/01RPN[1cZSN+G+M?DX_Jb-Q&5#
eaMa)8ZEe:1QQMRQ)E].WKBA<>3P3UF9=U\R;A]g]4#0)UDHZb@GaTf/3]6<RCfU
NJ,/6aS0F+6EWHV^UB;0\VEW9@E&D:HM-,3D=,YM:YI\9BM/&(X,@&3J?S6O\R&E
FYGHVU_DaGBAS,W<a).&fZJ/6<Wd,9IHfXINEFVf&C>,B-+W7<DT:GUFXHbAdLIg
A_LFVV,X\?L-H<dLeZa]Rd)ZZ2VHUCfX7f]#4VFe2gg0Zc?=&\_G8&KB;@O^9-9<
3C+;GeC))M/DB\c[,YPH8258@8LCc@d;LKA6Tb9:TJP&Z@#3-bS&:FZZ6Fc]c\F#
@.=fdIJCJP]U/804FDGaK\;PeH1Sf^Q;2aSDB;S[8cWME>dN-@+DB3/J<c8DeAHH
-C8>0aA256,Z\.Y^MAXD)L:fX-S45)0fMJ0?W]L-^1WF8D:,S-?I88O.?W^IQ(=S
Xe:3g/<JeB8d3?4@&gHa1BOfR@<bSVQ<0@RBW/N:<9SOQ12c4d2_e^J4Og^AH=50
JdMW-:1:Z@A(?Oe(A0KK0gb.2OI71-eXQ<XUeE2SE#IBWA[,9]Ef;+MG=90)JR?&
Md5@Of,V[,Cf@f8@dOI_-KKID(,KBRC48La,JD.U;\6WBJB.B<:d[=J>FPE6P[f7
1ZU?-/4923(\E440e6d\XWI,L_g-7NM(IYe)aS@O>b.FY/L=.1?UP^709GH_EDCa
IJ76<U]NLY/gMFXV(A10bUb:gc^dOAb9KKdU32UGX.AdQ^[OGE[+M<[E?g/@e]bT
()Y9&c9a\9aA7O3#NSIBeT_]D)+5](QfEFYEB-OY8;NGDW7aC5aL8/K_,DM,Q3O#
9[-AA.&b-\IQQWZ\]DRe,L\I(746I0[TI/11Y?6cO2cfWJHe6Y+3U5=JYB3;6W5<
/1[LQOO-7_]WG(.5eS3GG8;X=QPM)--QVfe19[HTb_Sb;Z8a[X_#>A8f3KQ0FKdd
[>;#7\P>5=KN:L63[\7QLLEaBIL#72.E_7-6+Z054]g&6K0C;DcL#EEQg2+<BW(>
eZ)S.MEQe>RYPHaG/@8J]#X[G2NfXA]B(-S6deN.TQ;L1K)#IL-V5=]8e_@[E62E
WTfFG<1_0W/#0II+13e+c\^7F7IR[K;WE\)ST;.;Zb)41F#65AU]7CdF\Z(7RQ\Q
AZXBGR(3JD#H_A?MV=<06CC2B(A-fBU.ZQ=9J\3Za<()4X?)g6@GI;.aS2)\<_,1
7A@\;MWK)UE(_3Vg]2#]?bLC_#Uc#?Y37/(_?NcH36-JB-gGC@K/>cOB;S7U#0>&
E0/BDNKX7ZYN29aB84I52+,CCF17LT0.4Y,=B&?WAUN#<2F0)XDX9B5A@Y>R4#a\
06I6:7JfH(cac?G5]WH&ZZcE,#=Eg:L.f[]:1]+/V(AIQ+01EJ7MdBVHHEg;@W-F
:B4EAXEN+,+K(WU9^\deJ+8,4YZ+DTY:ADa]C]1H2(0SR_-1P0.;GKZQY1cQ+6g:
-bMYT^F6>E,Ug9)cg.2ceQSJB):c6:,FBE(-=LQ-4<U9KU&K;_692N66E[<VX=WA
AB5E_gB50.\d-8141CQ(11Y\SD;A4DG2d0CG[N;FF)X\cP3,I8,&GI,g_9V3P[c3
P.GS\@FF-gIF3-5.Z\/6)ab+F[L2PIG(3I^[O@&7V?]..<>,5SJDY7ON;KY+XFeP
GDWYHIF#;I)>Td<\=fJfUa?KXRLMDe83V@B(Y1W&GVT>]OQ:H=&X#[N\>[I^U+Ya
,B&3SU9aUN1HM+Mb/3P9JCD4==C3])>,R&]F#;20(Z[CaZC=GJDFWP\fH]ABV^N9
8XLf0X4cOP4g:>3:WA1FZ=b6=TUd;R+N;C:eCa2@2V?aNBF5b-6[X_TB,P\gL2/I
MW/.KIUg(-;SafdGS,KdNNRK=\,HR](0YZ+[(U8V_])T7AV-:8Y\#Q_L51M95ENS
0+&eB\V9.NWA#SXK\_A3:NH+d]GTX6PBWI+#BEU77CD?V:#R^]\=AS&L6\^8S3@T
1_T;T3-d_@6=-Z=;(V.SfE67=,/?DT_OD8__,@O-,6Ue1I0@4&[9JSZNQIWN-B=+
]<Fd/#gZU@J(_Z^?Z#^g.DZA/,L?K0@dMc_9Mba[:9EJ,IQU6W)#/BZF>e>2JZeZ
#EaJ-V0JNK>#L+RUT?f5UdfX7N3DA@&H]M:EC1?BVg)U1B&8e,@KX1[2@S[FXJKW
)@1&&\a_HAcT^X1b.IBa3Qc5<=-2b.G[;C8W(2g[=T&^5K8OLfK&L3DV2Vd@GNc<
1;[-N+K?D\26&:DNR,fX)94Te&[4<3Q5TRK#/LM-;S62P6FOKZ/Teg<QK:[RB&9T
FXNT?&V1RY_SdEF:A[a7_T,c>NN5\+X(a<bQ3KX_McNP:5F0cbM18N#MZH5QFZR(
95IbAG_>ZRJ)MH>d9GLcf0V71]3P:46VEAa6O,+47V_>Kf=;cE1OKLf[Da4cU,P\
]04GW9+6:-ORT[(QN/9@B,5U4941E)_3TYSOE3d@^3B^Sca=^^7(PDS>GUf^ZIA?
-85_[)MZgP46ZQBCb[ZG0QQG8C<<?>V[(D4Z?c.HK,fEV/ACSgJXaUGKNIX1Zf8=
B_NYS>fDWF]B0;--LABP<E;26?E;5/.[b#>(8cV?[&-)W#D<.:P<RW>78087XNVa
]8-DS(24aJKR_#A9[eF[71_.SO?L3SeI,LX<,fbAH>0#CJd[J:8],?(BEG@C6F.:
994fd--A?L#FQ[T5Xb1GVLH4)7VeS#53_GfAJL1dE;;G5RU)J\&K,UP+c5WBc9WT
3UD?VcfH,Hd2f8N2a#OR.aT7-T^_JfJI4Z?a,)XPPW\>>64/:CMIFXM,65O@AFdg
;IHF^3GSUG9^(bTPYWe<<]E8+@/8^@);;C[4ALY3/:Ad6:S[<9=<9:PT<RO>c+XZ
W)KG7H=Q/VYU54GR1fFMBFX3J7HO_N+=>0AfH>Rb8N&QGERb@P7:PBBJ,g7YD(K[
HTX;==7>Df,(MWZ?,B1LfXZBS3ga@+XM[2L,g,b3(c-U,#Z94<@eS=A,-=,_9JGC
9#L<dA3)(V/(M)KJ)WQcC1U1b^SM^C#S)(G6E/^L6d<85Z7@XZ?J:X-Jd^e^UF)#
cA)eK5\\gH9SW\_5fH.PgUM^IeP2CZSDFN:2e\CHD]>V?eJ8fVDD)S\B;UV0[@8H
\PPFIJS?T<0?J#7V36QJIW@QW;2aY<,#9Z,+DATE,dbKBP?(8L=3YS5X:=&/^d_,
&7d+28<3f51BGdb[3WGGW6TW@c;SNS7J0&,W\QH\E&b_6e^E&T8B<=^P;KCC+WTM
.#&_=5@,?.SW06G<2.)LBd=,6O.2=55IXRJ-KN0AVE;P-]7G>[#=R504Z1&..&7I
R&gU,XdDQ]O>g7FHc9?Ya\LB3=9;#2=8bO?\OHSW_FJP)_6G#bJGZ),.>@)9e1FY
K+^d6/XRJ>FFLT1Z,9B\H0C-RR[UeO1G#d7>fH(\3]&O>e.7bB/TB_KIQ5A-4ISQ
2JY;_FK4-:4B=\=\_SP(CGP9F\N_;LTeP[PCNgY<I^PV=(^RZE01O0Z,?7FXe^GZ
@ED3L/U8;KWFET.F<KA39TGZ++Bf)WPM^2^Uf:2428-)1(G^H/AB&_gW12#@<R1e
cG\-e6(=B(VDd,@00XT_@\(.KV=>T/_<D:Y6ACIgQ@OJ&>9+?NEHTfD_c:01DcU9
LS7R)d3=25&7;SOYaZQ42[&@&T#1gTQK1(:;=U5\S[1-<+bNB6+T5STZO.Re:H<N
OL22A,ID0H.WPMP-9(e,[O_I+^1;d?/NZNC@P1OP;1C1?M?;DQKbYc36BZ85ZY&0
ZgVf1f?DJ=N5_?g>E[cJIcO:6E>,[WOI3f^8),aT;&\-C.INK2J/DS+gW>I5X]g5
e(I7ef>f60;LL4G[C\E=cJ,6DGRcI)4^EQT^T+/cG>#@+&/Y+2-R6E98>9SBYDQ4
=cea(#cdAYQ=K0<F[GH)bb_VZ<81TBFI6(4((WE+TcEM6?>.B[SA[>:@+QK^LWJI
Xb\QQ9a2HR/e9f@b.7P3YaA15YJJ(^VP-K7:M4C(11I=9R<Sdd[H.5Z7B=6_L[7=
D:b[5G2fZEfKd]V9aeS^RP6fQ-\B#,TD4V\b4]d.9F;7^09JA6.;2EAB+[4:DOXU
@bP8K]/7R5+;Q9(;@HQ-HHeDD5+]L4@c8,EXd@gJ^7UTScZE3[\G3N\\;4I7G;\e
>5gF@J1I(,\.HHDM_Pga8+eD3$
`endprotected


`endif //GUARD_SVT_CHI_SCENARIO_COVERAGE_DATABASE_SV
