
`ifndef GUARD_SVT_AHB_COMMON_SV
`define GUARD_SVT_AHB_COMMON_SV

`include "svt_ahb_defines.svi"
typedef class svt_ahb_checker;
  
/** @cond PRIVATE */
// Note:
// This macro returns the width of data bus that needs to be driven.
`define SVT_AHB_COMMON_SHRINK_WIDTH_FOR_MAX(width) \
  ((`SVT_AHB_MAX_DATA_WIDTH > width) ? width : `SVT_AHB_MAX_DATA_WIDTH)

class svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  // The Analysis port for VMM are declared in the ahb_master_common, ahb_slave_common
  // respectively, which needs to be parameterized to the Initiators ahb_master_monitor,
  // ahb_slave_monitor respectively.
`ifndef SVT_VMM_TECHNOLOGY
   /** Analysis port makes observed tranactions available to the user */
  `SVT_XVM(analysis_port)#(svt_ahb_transaction) item_observed_port;
  svt_event_pool event_pool;
`endif
  
  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
 svt_ahb_checker checks;

 /** Sticky flag that indicates whether the monitor has entered run phase */
 bit is_running = 0;


 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag updated by the active or passive common file which indicats that the
   * address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag updated by the active or passive common file which indicats that the
   * data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
   bit first_reset_observed = 0;

  /** Flags that is set when a 0->1 transition of reset is observed */
  bit reset_transition_observed = 0;

  /** Sampled value of reset */
  logic observed_reset = 0;
 
  /** Event that indicates that current_data_beat_num is updated. */
  protected event updated_current_data_beat_num;
  /**
    * The configuration that will be used for the current time interval
    */
  svt_ahb_configuration curr_perf_config;

  /*
   * These are objects of previous transactions for tracking the active time to calculate 
   * throughput when perf_exclude_inactive_periods_for_throughput is set, and perf_inactivity_algorithm_type=EXCLUDE_ALL
   */ 
  svt_ahb_transaction prev_write_max, prev_write_min, prev_read_max, prev_read_min; 

  /**
    * New configuration submitted by user which may have updated performance
    * constraints and which need to be used at the next time interval
    */
  svt_ahb_configuration new_perf_config;
  
  /** Timer used for performance intervals */
  svt_timer perf_interval_timer;


  svt_amba_perf_rec_base  perf_rec_queue[$];

  bit stop_perf_timers = 0;

  svt_amba_perf_calc_base perf_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_write_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_max_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_avg_min_read_xact_latency_calc;

  svt_amba_perf_calc_base perf_max_write_throughput_calc;

  svt_amba_perf_calc_base perf_min_write_throughput_calc;

  svt_amba_perf_calc_base perf_max_read_throughput_calc;

  svt_amba_perf_calc_base perf_min_read_throughput_calc;


 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (`SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Detects initial reset */
  extern virtual function void detect_initial_reset();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Initializes signals to default values*/
  extern virtual task initialize_signals();
  
  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Returns the expected data value for a particular beat based upon address, 
   *  datawidth and endianess.
   *  This is invoked for Write transaction by Master agent and for Read transaction by Slave agent
   */
`ifdef SVT_AHB_SLAVE_DRIVE_X_IF_MEMDATA_X  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`else  
  extern virtual function logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] generate_beat_data(int beat_num, bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] beat_data, svt_ahb_transaction xact);
`endif
 
  /** Method that is called to get information regarding the data/bytes for a transfer.
   * Currently tested and applicable for AHB_v6 incase of unaligned transfer.
   */
  extern virtual function void bytes_information_for_a_burst(int beat_num, logic [(`SVT_AHB_MAX_ADDR_WIDTH-1):0] beat_addr, svt_ahb_transaction xact, output int num_bytes_to_be_transferred,output int bytes_already_transferred,  output int num_bytes_remaining, output int num_bytes_for_curr_beat); 
  
  /** Returns the expected address value for a particular beat based upon address,
   *  datawidth and endianess */
  extern virtual function logic[(`SVT_AHB_MAX_ADDR_WIDTH - 1):0] generate_beat_address(int beat_num, svt_ahb_transaction xact);

  /** Returns the data value read from the port for a particular beat based upon address, 
   *  datawidth and endianess 
   *  This is invoked for Read transaction by Master agent and for Write transaction by Slave agent
   */
  extern virtual function bit[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] extract_beat_data(logic[(`SVT_AHB_MAX_DATA_WIDTH - 1):0] data, int beat_num,svt_ahb_transaction xact, logic [`SVT_AHB_HBSTRB_PORT_WIDTH-1 :0] beat_bstrb);

`ifndef SVT_VMM_TECHNOLOGY  
  /** Returns a handle to the local event pool */
  extern function svt_event_pool get_event_pool();
`endif

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();


    //-------------------------------------------------------------------
  //                       PERFORMANCE ANALYSIS
  //------------------------------------------------------------------
  /** Main task that tracks performance parameters */
  extern task track_performance_parameters();

  /** Updates performance parameters when a transaction ends */
  extern function void update_xact_performance_parameters(svt_ahb_transaction xact);

  /** Updates performance configuration parameters based on a new configuration*/
  extern function void update_performance_config_parameters();

  /** Collects performance statistics when an interval ends */
  extern function void collect_perf_stats();

  /** Creates all the performance classes used for calculation of each metric */
  extern function void create_perf_calc_base(svt_ahb_configuration cfg);

  /** Gets the performance report as a string */
  extern function string get_performance_report();

  /** Stops all performance monitoring and kills the thread that is tracking performance */
  extern function void stop_performance_monitoring();

  /** Enables/disables performance monitoring of each metric based on configuration*/
  extern function void check_performance_monitors(svt_ahb_configuration cfg);

  /** Enables/disables of all performance monitors based on the argument */
  extern function void set_performance_monitoring(bit enable_monitoring = 1);

  /** Prints performance analysis summary report. */
  extern function string get_summary_report(svt_amba_perf_rec_base perf_rec);

  /** Returns is_reset_active value. */
  extern function bit is_reset_active();

  /** Perform signal level checks during reste*/
  extern virtual function void perform_signal_level_checks_during_reset (
                                                                         bit                                         is_common_reset_mode,
                                                                         bit                                         is_ahb_lite,
                                                                         bit                                         is_master,
                                                                         bit                                         is_active,
                                                                         bit                                         checks_enable,
                                                                         logic [(`SVT_AHB_MAX_ADDR_WIDTH- 1):0]      observed_haddr,
                                                                         `ifdef SVT_AHB_V6_ENABLE
                                                                         logic[(`SVT_AHB_HBSTRB_PORT_WIDTH-1) :0]    observed_hbstrb,
                                                                         logic                                       observed_hunalign,
                                                                         `endif
                                                                         logic                                       observed_hwrite,
                                                                         logic [(`SVT_AHB_HTRANS_PORT_WIDTH- 1):0]   observed_htrans,
                                                                         logic [(`SVT_AHB_HSIZE_PORT_WIDTH- 1):0]    observed_hsize,
                                                                         logic [(`SVT_AHB_HBURST_PORT_WIDTH- 1):0]   observed_hburst,
                                                                         logic [(`SVT_AHB_HPROT_PORT_WIDTH- 1):0]    observed_hprot,
                                                                         logic                                       observed_hnonsec,
                                                                         logic                                       observed_hlock, //hmastlock for slave
                                                                         logic                                       observed_hbusreq,
                                                                         logic                                       observed_hgrant,
                                                                         logic [(`SVT_AHB_MAX_HSEL_WIDTH- 1):0]      observed_hsel,
                                                                         logic [(`SVT_AHB_HMASTER_PORT_WIDTH - 1):0] observed_hmaster,
                                                                         logic                                       observed_hready_in,
                                                                         logic                                       observed_hready
                                                                         );
  
endclass
/** @endcond */

//----------------------------------------------------------------------------

`protected
#4aIc+V<Cc[gB:_S@0Y,QF0+B=YH/DP;Z0<e=/\U&9b);-.(a2+>&)FNEXL?9[+G
NI&+&7-RNHO7X:4&XF\^\PKBY78Z87N[c01.a>ged4Q/ZEbb)H31K[XBJf0^J3[:
.--<LXO&2[159(49YI8LB)X,NWB3>G=dX@+KUT3HA>2H?TN\B08[9b-\^HD@^D[6
F[;Z,\ZPI)cMTXK=+2HJX2gR2@Xa]Hc=?Uc=E8=4)MaKE0f73RW0U8#OKOZ]W^Ob
&PAI08IYeJRCXMQCUKD<E,EWCL:1c@\J10??6K03_a/e405_O7NJQa&@QAWgF=DE
8?,DfYg0GWTTT@b#/Me]aTcFW5P/gB,D[9@M&@^eOUf9&&T:6BUZIW=1TPL,>Nb5
S;YGQ94QK\=g7G))f&79AecF6$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
U1T&e&cP(0?3CM)eY::<V&?V)fEb6UI?]:9dMQ+gN/2<-U>E2,cg4(A,J>S=aQUT
Y/6c.FgMJIV+-1L.=D<8fM]T9@=1fR#KcOXg,a]>=.Q;Q&7G(=b]GU[e[-[ZdPU(
E#SDdT#]2:AX_(AT@)R-Q3]gb4^=cYd]eL1IW@+?[\FQ8aUSJHBAI>KdcL@[.:La
+7fUBY((:6JB>:ZZ:_XWW-.K#C;-905<=Xf92_@gG;MQ=ZDRgZP67],7@3A^#:-(
&XMA\Cf5fA#1Yd6DE]HD\QPZUHDd3W?W=&fS#]S3F?<()0I#NV2QZ6])WV#+Y)TP
f>]+6-2R,A5^6,bX-E9MdV]g6\@SMS9A>#C2<,=&YQ\3PT[]T?2BSHbK(?8,b@]1
Wfg&IKDC09U5C8KW>P_2,C[0_Z9<b:<\\-1IVI&:&B.DOI4+L.S9ba&-cPO>-B4A
aV]VJO#EG@=TB4()NG#/(K>D\c^0HHH10-+UeDI9.(FG)dNIP2&L:]=M/^-Q@KS@
+KM:WV6G+OR_&D+9]#&R1T4(S\[.Fe(/dc=/NL\VK/Gg,F[IaU+W<e4MI3D21\@4
W^NJU\\EM?3DO3>T.-T;QPbMN6B6Tc2>T6+;P_+V]LS4U#VXLY-##\I#=RZP8P5f
O>3eaOWg.0R[JS_D.>:I_,@#TgdVRAI>)V,A4d<26LB/AceE-XGIZVM&KPbGI5GW
37:f#(O_GFFb.^73cHVa0?DSS1YfPg^5&DN6E6F[B88QWF9>Y>U+(R_e3/]@deXW
_K4ESUB-gI=;c=&[b\_)Z,c@Hc>Z;c#53L&@7A>NK;:X5RKR6^@^N?+?@YERG\LT
AQP;<X?4LW<,AWF#e>Y>177I9QF&9Zg;FS\fB/C438<LRQ,d6TE^f==SE5NQBD;D
XcXeAQ3WUJ6Q=<9:d:3UK88)4TANd#XR?]NG=YZOdaeI?a)Z<OKJ6F-.FYf2FLY)
B0MbC+/g0&bB8F(Wcf>9QTY?:\=&DUSbC1(cH.CbN343:V[J66JFR#@AZb:C+\.c
V1A)8/S7G5^P=#B,Xf0:0eDDU<EN[E[Y(P\)&PZ<_HI<ZRb)e1M??g_2HeFaRORA
[JMX]D_XU4KPb+#<19H;,;#3OQFWNVLJaI)@8?[@??N\A:4;1BaP]8.e@1T^@49=
@g)gcX3&>a<QNYaR(I&#L+K4NL=(/P]c>-^1M4E;b0NgNgb(YXC+Oc9M,G[)\>D0
=W7#7U]Q&DfCeOF4_Zf;ZXaMJ]E@]3W))R6QK:@XS2^Ba5<5N3FO+R?H6&\C3)@[
.(R.JgLGS2R-.+V120]2GDW[]_Ode>f&?:W&OM+S8=47+AQdb9T4&YF+VREg6W[1
=ec\PWY2BYGIC3TMBKC<2N7Z?)F?2+(4Hg_Ia&Za7aFYNROeT5\J>_CQW/)3XgW6
I_OOJ=Y7>-.ZP=J>96Z,@8\e=Ua07:\]99QXRC:=:Hg&a+Ja<-1@75,X.AH^\1I?
Qc)F^GUWMBVQ7M^aX0MM0d7e.@ZJ;-R];00>9Q#F6O+S3eOY(=Y&0Y0;afNTS9G-
):[2(gAaLL@;QD3/c;;D64=gA#R>KK]/R.-E7DKSWc(,d@(?;aV;.-(-&GI(]6;1
)Z0]F0cA/21\=fD(V0[,<X[])T[AFgfe_=b?5d=L_:V;&=KK462_4gWL0+):EQ,V
g#23(B_e5@a..@dXY;_O=SAI8HMW<T+M&8D5U-#5fc&V(WHefaKf2?X;d,B-FHQd
cP][4NU^.0;;-1R]YgN4SbM1F&1U.IJ?5T5UH61)e,b-g+^7)ML&YBT@a;?K@TG1
I+.N2LO&HQ?S\QT@9>#5Ve0)fA:O>+VZ(@>WKLH1QeOC8PUQWAc-+gFM@E86Y9/.
P/+HL-/764ZH;+:JXg3b0Q-e6:<cBD5;-(9OeX>D#;,X7?75bRI]RPN..G1f:S(L
T+:C3d.&5)\WP0C4FQLLK7<(JaHY&^GSHY-,W/KD\CMWVY&c2g4#9G3d0-(D,+>:
XK5<1MgBV)1OZ,>I@7\WTT-fJ=]L+]XeIK33S?1RVe^)UOUM+d:9YC3I-^f;8a/=
_9Z<_BfZIbfcdA4#ZLa\&/0KPZWLO\]-9:dSa:?/_Y,;(a(@?#AY,=]:-K5\SSE7
AW?];:=3R2(SY>:970Qe/0ESC)E&S/)/gdFR-JOA8GVdc6H]XS6&Z=d<CZI@B1Z7
;DYQEX/^,)BZf?Ha@8[&H\@)d5Ua79B#bPC<A=WcO-fD0ODTAbbOWWHgcH7RB&GS
AgbQ][+\a(5f[F[0]=8W1XQ.]8H;a@/O0MI>5=U)(ad+e/HZ.<#b6K0DR+#b8>WO
4M2YI0&d7J8F8E-@I#L3:<N.]WYM.BU=c^/5C&eQ,.L3;1;\T?9C)e^bZDPM@_3^
R0&E>L]F]#DM\#A8KgM6,TTS&VCfWX+^X@;L5[C.^Y3R;d4#&SN[3F3a2(_9/C+_
G<45WD-ODC=OLJ06?d1<dXf(AZ^BfN#agB^\S<U75:^ART:7;C/QVBI-/)XeUT6-
b,dS,@.G1NOML_E3\fEW[#Y6WLDO1E)&^P7^A]=4UCG<X,WN4S04+&&=]aBAd8eY
3,ZEB@[89O7_\A<1;0?4/.Q4[D+T[2IX92]--c9O8E3[0:,M?X,4cIZJ_.A5R\H6
,IT:Bc_Ed+V<>O]9L,2N]-KSD7:Je7SXP4gBYZP0K_[76(5FV7LTg?H)_g4?L4Ke
eUJV[f+bP9L\HD@aa5--?09C/M/5#fOH];1J-3,XfB9ZPT_?e9ZBSX<ZZ,7C54?X
2f&IDfaBZbS=<c^aXXJ)]VJQ]1?.(M3X^@+B7BN/I:d;A_=Y<M8HI=?<L-A1KH5F
bU=QYA/.OQY_ZYY7L^g^:=c]=,WeMeeePC[00)I3cSAY9YE@0P&80[JH8dM[BGGJ
Icc?Yc6:bUG[aGgf1D+aO0C8J0RBHI^;;^I\H/DfOE0>#/G&e;bc^A:C/LBQTcg9
>75YWCU7:LW\Ob0TQO&F+Z?7#F3gWU6\T3I_<;HZ?_SPN_,FX6-)HIb_>4>-bTbb
)I)V^e32A2FdeFeK-O=cM#F8MQYG_0G?EWgX;DeLG(169<K<<;F<9bU==QN_T=@g
JBFUZ:Wd#/SLa__C;,Z5HF>=N4A4]RQ;C#20/KA\W81;R)3F2^==^QBf9LXKb#@K
^8@D^>B84P/8>:138g(MFEV>04+B?1ZQ\Mf(?<^BMPT12?1P)_;N42K42?<89]43
Xd=b;T?A@CXYP@?<K1:<5Ee?4:L5OfW9RW:?#3([TK^^5E(Z5+4]?-79L>ISS7UN
PJUPZ29gb)(<P5_f>P&0MUN17gG&#K1V<S0N1;c\A0L?)Xa[E\N[(Ecc>(F&D+H-
LW8QeZV4Gf@)Nd^,>+]cC#[GAN5dQ0MHg/Y[;U_C<-(b?^_QVD8,?4SN)ACJd^Gg
\3QA6T5M]6\7)W4]:HVC<3.2HVC>\A=D4&g9]?@-/bfHMdH\90TaeG?,X7;WMLC@
e^^e4\O6AFK+1Y9g9JSZ);0\--RFM^R2#8NNbM:(/W\QPd(Q4OMBT\ab<ZB:ZcP@
=2[_B#MJ/RXd475O.(=F6,PdU.AF&R3B..+M;+>gEbKYa3cB/I)@W^)Xaa\_J?&b
Z=G),f.CgT_T?d\&C&]++0S(]A=c/O?J5Y6J189X_<H;Fg[<FBZ[TOE[9O3g;[[D
2(I?8F4@^P>Qgg,K-dGNKR>V#8;P^H:VK49X^7Ggd8Z.;RJ#]1][^cDe]FXcYd\W
B-AMbg_cHeP)KQZJ::A.7<&KFA,4;/#NMMJS0b45J7)eGA,PGLGJT.4a/Z:3S5(Y
gG,2TgV_GdC^EOCU2f0MJ4POI::NGRJV&)H>cdBT;Fa?]02I<UeLEQSb&/PN-+Ea
WBE83[d41EPSd;Q,^M.7/0B-TB?&E,VO\L,Y.LfP1,_.GT[K1QR>B(W8cNa:N4ED
d(AfBW6^[(,dKT@(V]egCJc-7.12BZYL/#ffPQ&eRbbJ3fd>[^4<STBDH,:)-V#g
E##+#<30;W?\ZAUcLL@:^<O0@E[U37W8e-OD?<8^e+6AcD,YbKEAK#:BR-KC:dR=
8HUb&+(8N&:W>](W>>@bQ+ZB@EQ7B\bJXRA,,<H;2PIW,_LaRJZSU_L(A2=#PdHF
1T0>F0H,?]]NYC+^OH4K/).>18Q#c:E=Ge@FMd83QgW8;.J2)-[<Q22[gIe5:=V.
C<U5N>^bB+-TJC32;49ZA>?9X7EaBCD^XCR&F67ABa/B^_-:AZF9J/MbfEb-?L\c
7X^JbbYDa3QM-DV@C:\RXd[.GE+V/9b^^+,_6CMU+eQY]0J5>MbW#WQ8NUDCOZ)[
F-R]3Ga#dKP0].R7BAMVD7VP,b4-,cR1Jc4\DI6-eDQ=HXY?fZ1.?V(aM)8QD3ZB
WD2G]E/^_]4FYP6a6G#C\f6CK\1US\ffMa:,;+g;4HOZcM1ZY)?1D+fZCe#b(7LX
V\P/TfU[MK)2X(^b7V/^C,Hg&:DTQf(eA4Y#L(64@/Y@P+/A>T=>0+#19=_a^?O=
N0M&Xa6,:,]gU8b.9?f-_2RPd5)<S:1]GRB>G-MSE6@DK,=60c3&T)\77&#V-db[
PMCg(R)P)YZ)N_Za(3Hfg4<(B&(A<RNba:1=>9U=&N5RJD47TN[d?S)+<Lf:#cRI
Qd7P1e-F=S1fR3@WXI_8N#Y81TQRdBA9]HBI&FUT5)&aVFV9UJ[:_^LEe)N<I^@?
2)2#d_,K]BT?bMP.>+G1W3eLTMH8FbFHW1V3T\W-..)L\Pc/UM>PV</?5^P3EV?Q
5,_693;G.MSXD#69<g=bZ;QQaD=d1=)Z@P36,.JC)&@Q[HObS>L:+>bO3+?5FT,K
Y#E+eIUf)+T<+.ZM(D1YO=;DC?-C_c&:\O:PcISOOI.W?a_[Q3T13D&9=TXUePKN
f@W4E;LC,S2cA)6X39-IZ9J:bIP(&ORaS#3d/2gHCAZ\HWEJB;EN06DXIV]DDfbS
U4GZ90ZI80(7Z^U/0/eW/bR4F0-MD42NNQ[PG<V1^8Y=f2eGd\I\+,]B(eKccU?5
C^P+[[bY##V@?^WK4)\#Df-C,/.b(@OgeC?,+V<94IdPF7Z<IUaB.4C1NG&GT(NU
R>H/WQg^PPSEHVNg;Ic/fcT5@,5W\GNWVfcc._3?^B2Rg.G3X@JdA#:gK9IXBZ^_
]X9_\<:DIEJ_Ree<7/02?,R?MDaU&c0A1PDaXLGG>:;7+B/6G-9>A#]2g29b;G4-
fZX8>1T-O0TKBS2&)C1[dBT-Yd-:<IQAT7+EKPCg#WMOb^/e1b(GMg)(F+LS;0:/
X12L,a+#a7dJ]P\XVMV>e1OE@05&MO4N#5@K;;#5J_?QB=dT-WI/C/.KW+>7Ig/N
H7f?R&9GC6U&38CG+;5YGY[@G01a&LFLOU+3-JU;f-+VfRb-VA-c.7S)OK>NZOLB
&TQ^BA+J[H[b/];Ec]6U51WV6]JgTY._4]SSM>V2-69,\GN1=9Z&a@R11IT8(bKL
UPEFa2Z(XeM>V/OTQ7#bO[9[W]]V4<VD7S>D&bA;ETBJ_f7OeF-)3[,eg[0T(,?G
UCc:c-ARB97EGH#)=Rf[.V:g4OTb9+b=Z[-M;Y4a.EV:Cb\)+#,5(caUe]feI;#?
fCZdX.\[fIaS,BXRM<MFK]Gb\a5QQK=[B[PSM7QK;U>?b2,2:_bIWc@<P6J0f(6]
>C_R&<WWW>(#I&G#70_J1>F9DY63ZA10C#gLDg4[b-8L21VDTK[=d#6bQ.;43]cd
H+7\H=?d+G?bDHBb::H&dA2e:/Q[ZY6V<JCN<5g4?-[\NR76)b8ce_d#[V(9_1JE
(D7=<H1.7/+?9_78TW?FXKK<<&Tf4)dcM18DEF_A7&U)?dXR3N:<;aP^_QWTB8fO
?c-Q-PB3d5T<204c4XX?S@K/\YN4b_5FeD[3f00We:@23.6#F7.+g^_YTP3E6IT2
TTF^9X1_-@?PU^9UTFDIV2BfG[F+]?LU7ZEf09aM1-XH)HZ?1;E&_8^XXG7S12C)
6_eO/O;P07EIOY6-cEdQB(c0cPd19&));TLf9>GI2VM:c+&19D39<a:.#GC=L/32
Yf7,@eX<]J]I9db__f6(>3bCM>1KDKSK>6O3Z2<Y3WPGR2@P]BIYPgdG1TT8bWZ,
L?(QT?LWFL2R5f/=<[[[VB6J?&fW2]GY_d42.\SVJNNA]:7;fCBYW+.0<[\=[3O^
H3TZ?J#LKS8SF9BQIg1R-YR_-K&A+[8D(@ZQTg5.D^K<fQ@V7A7P=a4V<gT+K3WX
J>=[_B7#/J9>H.AL-65GcAG=Dd_f3NbCS-51\^QFIYKb>NLeIB<(g.K\gU013Le<
B,5XG5/4O1BO8g^W>c64--=5dc@W[EAd_.[K@>X:F.PJ-[KAD>LfH_<]TO1ZOdd)
b<<f@@(I&Ma2BXDZ\FZ@(YWU)6Aa2@baa)&&WQbBdgT2)MW;gIcGSM9)a:=WN7(H
.bQBLg<eV1(;<c]b^VHd/=-EB;^UcHZH.4HF=ZR;=]d&_dV7PD0XcZ+#X#,9-XUK
#MP&=Rc4?eL9bJ?ZTX]MO0K2+L8QX]Qe2UO^/Td:\Y[PW9@6@06-AC-WfJAV^H=F
9>KIF=+-B&UIY2[F/4_AV:<4I_>EBN;:6-bB/+1fS]98V2;3^Q(Me](2_MDD,IK]
eVIKTD+@:2UQFfaH+C(aP.&#A##QV->FOP>7;A0(&YRX7<)S6/JU283.&@5_=-fU
_AKWb3HA&:e]Y\bC+EC.+B6V\1XG\eB#EK3=&Vb(@-YE+;f4C1]?=M@@(4ZXJ;PS
K7J])>3KMOS,^85:#9PZ4^X&C2d5:6)^+#DNIV&Yb4,DV&)V1Z1YVMHB0Z3#\^EZ
ZgW6ggA@?QXTA9aZ9T8\>VPH4B/5?+b]=#G&)1bL.e<<##07D\N;IEg/=[A/PfQA
,(-L0?AC,DEO,OaQbQJY>7)9f^,L15=[BRdHMFcAH9+-VMB;fXU74Wd2TBV0YDaD
OFD[6;@4a5_O?JJ<:LRN<a=/#.)=Za5Ta&=12M(/M^/e<Y0V9>&3Kd0A57&X:D3X
=[BB-Q=eJ\SgC==RSVMIe20>K77HBG:0eY:\Ia\D(6,._)MC(>UF22;R2RB7YR8>
\CR5GH=7:QQ^;<[MC)#]O>;^XK.;54d(;9L(J8.)4SOaQfgHSHEd/S9f]_AgPX\[
0Ib#H=<+A0=LREGaLO?.f6-(;B.,^=MLO_,9[Wg>EXYR#^1:A<Va>NB?>KA]f1#@
RJ?>LdDCg]-d>2Zbf&T5J27(KdQO\]FI?787S,[@ZD(CN&N-V3-TX\D63c=cW_CG
I(a,6CB9T^QJQSIAV./R#bM5Vb]96/-K),?V-bY:J-M1+5F6O[C?EJ;WU)@@-#DP
[0Q_L(a7YZ9(\>Y3>HW(_,V5XeORd],ZC7Y6FYZeT+/G+3Z@J0ZQ<Fcc[9OVg7Dg
X3XDGJ[FKB.:#0>>OL7TcDSfe-2@66WGReVS#M/<8b[C9#]OLIL(+?.IQ-[d)2c&
282<O@@??>KAGY9[;EI/[?@1WR3,OSeTg#gT>SIJ#<S.BZAE\VJeT0dSL;2GS;@5
d2J3JEB-VZI-88N3:)f2[/0/.b]Lf_:\Neg,M5^c1(cG62L\+N@eM<JG09MaTAI,
?4>.:XXI.J14JS_7WZ7bdTLW.DK1<WFAC0^.>fW.Aa[.WJW88S^eSKLA;NfI[V14
VA=CU^NUER^BEN1E_6\>JS3,WM(QU,H(136?L1#>HVf,eP#L5fA#?d/[799-RRb-
V]A(++J_UfH8WI6_JcQ\FaVV.(XfFf0eMZ5eS9;,c.??X0]CDeZ93H@XP6EN]<7J
R0@NDU#EYWKfY/QBc?9cQc1GFGO_bfdf2SVESQW&bWf/NSMc\H+IJ)S_Z-G_BY.,
c6bPa]WWXaH35?M3b&Q/B/6X&0]2a8<E2M6W#6;QXagAVJ>^+<dA]fA/d=b8;3Q4
Q15FZAYP&e6Tg(QO/G>DL+PP1?Y6\[f<3BW/8#+[?5)#P=XQT07B3\[H46D<:P_Y
2?d^,KAI(VKEH@&Pf[&eBeY>@3G[0.:1>Z...JQI[M)6CMX\P#ffPS^S4;LI4.-^
N9:;bUGDdXJRNeF:1?R=ce;4_=d7[C;C=fDTBfY@1A0,9,Ma57G9bR,XCJ9Cd\NN
V6G0fE^RFCVCW)NP]YRf]+I3<,;T.EG<NDfeQ<+]^X43UagFc]BN)/Z:Ka#0Sa7X
e]WHU5QD98).aHMZ2K<;P8(12Q#bS(V).1)KO^T_/+f\@Y&B4AcaAS(T(Ta2)4-5
F?WfGW3)RC8H+&\4Ogc[[OK\=D+.H^.b)/1G/<\H#gOaDQB#6ZI6U_\97N=(eAS-
;#b:OH55g.C]&gJ0W/(R-/POF=?()HGEYG[b9JBO5&;d8Z/&#SeeHcd/&F@O_#3V
b=aI49R6#HT]5-GIK?\UcQ/=&Ae2N@0MQ#g-&-?0^5d7]J34W-\cKZT\fG_4b7,M
9=)(H;EL]RMYdD4gXKVc].:=Lf62H=[C#,F2C;84f><Vge]2@Pf6<=\8GEC,+0^b
#MeJ2G:^CH[c2c]5C6\c86ESE,Sf^IWa[B(&^J9C4<YgYe,/7d=_/]ICD0V=Zd]]
,gZ+H<N4ff:D1ZLL#g5,T-KN>_-&]Y@^2DV<@1D[A5O5.;9b:&E1+7KC<-1BPNNB
@]BR=A@3AH_F)U5G1UV7:P#Y^-HE:KA@PeG9dSCBYLXY]KU9X@+3_4_IGR\+[9,e
J12,9HEU8B45FCA-?)5GM4dQ[>DO<E;;QDTV2#;E464;f;(])BVI.@e6;4>2H[B4
^e:R]J/5-AK]\-^;O9U#@;S^)=DAZaKIQ@)OX@ETNf/OQ3W[g8\85f])0DQU<SY6
V:I2L&c1SBN8=</eTe99F#)Nc]G8d@D)&X9]A^&dF58f_gcg&ONLMZe,b>IVT\[4
.a0c86-O70R6GO1TB-KP-TU:E1?S6PBO7D4fL>WB<8@7Id2A>Ycga,e?EC@QEZLE
,Q/RKU9.XeMJU(^8c]..THSg<EBG^GVOU(+<_(bH0[U3VXa<UH6S\5fG8,NX]>=L
DdW2:cPd-7^X@V6@,08L16f8_gfC_,d?LCeA6WJ8C1-O>4]P8^QK;-Gb3B-gddPB
<eO)2J8P5CYOT(CbL87RJ)@BQT82Rg:GN3fFY5bE-?Jc1ZO^]T8J)&K=2>)-+Oc#
;fKV#OGLO/39^=L1?g[L2c9_B9INgI,,I]R<Rd^:Y&W8OO+,30KC^4Hb-L(Y5QN&
YSY)\D?<O^Z47Abf2@Z:,NNd#W4bc4HC#6Bf@K;RF3b-\1623f]AOWLG#C_?SD^P
6ReWGZ;#FM0O</RPfQg5;D8Q;[YZ[@5)0C7F?#NIdW3BXY;2ML^d3Q0SG8LX\/0b
#U).K<UgQ1TVT8)+B^^(=#@B5G2^aLINZ49M/1PMI0</+09a+,UXf68YA0?4>g#L
:d._/M:4G?;:;b/9NZ;Wg:_2/S;;IcZYCd_=ZJB@^^)KOD0DD#TaYg;MHaUN]JgV
(V8=@.6^Y=aE4_3d31O)/57]ARFNe+d(;DBZ4WYe4@=PJR>6=H(LNO0,9J_M87LI
:]DKWX\]Re;<H<DBK5&R_F7WBR^:U@5eL945@=103]P>5M8a0+>fP2M?=Kc:gf:I
MIfJeZJVL-.-MQ,^I5,G;&D;NUVXgV9\,3P]BT.],/T=e]GYFN#:g8C.,8_Xf.eL
H]_QHAKYDLcMC7f^\&<[g7YH^?:CV;7D0)NGdP0GaJ,QB./3&1M5fI7?L&9MKN@L
0Bf.dVfT@.(c-/PAI^?,H)-H+8GP[1?/EU&;GC(P4eC2EFe_Xe7fKLST&0B0+&:,
?_(&;cD6>=:IZ&gcU50=RP)bO0bP#2R7X<aO/d,#S?5T)KAL,KLX4b(HH\<cZ(\2
;@#X@>GL]6fXKePcdUUPfPLS?H[E]4B?b8b4>7J@_0DCFfJ)7H1N9dGK_TA(a50^
?GF-AebYJFg\RPJCRN<gAa.@&5de2SU^,UVXY6d6gVGQdI1EJH6SJEI84@;\aCKJ
,OP4YC>KFE:]AFC3D\N2)Ma=_YU0O+S0Cg?Fg.aGFF+PKdO/MA)U8-W,BR@HXX_b
JOAJg@85#E\ZYGUd>W3cKC_W9f]>?K+1f61<#4M>e&FS-9TH]Z<&NXG#-c0&a(+<
4J8ND1I[&A&UPK19B39c#R;4VAXM:(2&&[/L..b.H&G4?PeR#H)X4d_.+Z#RWDO:
9Ff4;,a(=6g^F.M@PB@O&c8@c<&4c)9bD377:HEVR?YS8>fYX:ZH.?D=_#[0#MQJ
g4>O1CKC+F@-Ze/&R==FD7QR65#PP3-Ba\E6C[:2W2>fE.,ER(+MLE_]C+Vb,ZOC
7.D-1,Ud,&^.e3#8[fBYKb8c+Y.E;C5:8(?e#NX/:dH++\f4HI2EaO^aeEW)MdYG
44U4EU6CA-,/_R5+0e-X(@ef\UF&GG,59P]:I>W6ZNGRScfI(@d)IF7(gO6YSG\f
A,QV\=[7?Q+1H&NQbN.1]L8?dLPg6CL9,,>JL]R??+B(-(6dN^KL)5V1g-KYE<)=
6K0Md]KRH.F_8-,XW,@^DHSe#SET&Fd7-K<K<Wd.PH_@(T-<L6-YeXOS)B25^XXg
V@E)@dHgHg\H?_dD]P9gZPY.c]Z)[S&La7-<bfET[<?BS;gC^5C9A@=3aD/K4E5[
[FK,CRJMY.Qa\VAQD8]AgLJM?1c#D.W=gOP8W+C6#g>-7I?A<@8;QH3513.B1]9&
OF,BU;:.353<]5-I0XM&,;\DI_()]@>@_X:238[6\:.PL:fe1M&4BcOg4G+;bge4
+5Ke1PYCbOd_T#4?],:>\c)60I?Z#\1VH&)XDI(\ULB)460=.fH^B@9W-HI8=:Sf
K:g:W(&Ma_GfT=H9aSR3\?=gV&WUAaO/1KI(dXVg)RACcXg3X<(b<SMMN=DXcSTC
^1e?ObL47;W<M6N7Ka+1_3\bJJJC?52ag0)e^F-<Y5J;@gB]1@>gd4PgKUg?T_gW
74/<&f&FJMV@@>D5S;fT7,=>&AB<TSB#cN7C:d<5AcB-Ja3TR.#NIe(<e)P#3;6B
FXV,Z4]Z[/2:U-K@cOKZS[<>Oe?2@eD+e42;^2+<JcDNg)gO)D9d2WaXXC8/7F(O
:H+N14E7).E8dKOSPU]UDP2@JH[FM(@##1Q+9NINUS)e?g>2SbFPI]E4T0^LEMOP
ZBc->:)U?=6<&D([S3a5SG:>a9PbTK1QbP++#:L-C/Gb/>Ka+(PV^T,>>4gI7B<@
NbL:B5K@>?G/2HUbIEd0)UNI]d;>6Q#2Y=7[O,\<;M4;72J5,WOTgC0DgTVd^A#V
Ra&#S:3N@;=DBCDTa:<dV57>b.==D:8JD3F(.XG&.@YCO(cLE3#\XaM+aCVVe.Ie
e(QdM=PPFG[aU)BFZ:4e0493/G8COB5f@@WfPJ?cT0+&>b-C;TG/GOFe?3&7T6RJ
6g_Q;e6)gKP4E^0d4KV9]C=5,NX+2S)(S8+2FW9#[.<3@DbTJ2Ee+RAdK11Fd&6G
RD??5)a)]0B4X_/Q>+7-S.2JHJR8.1,H1Cd6O(aE&>D=\MO&9Q>T(J6]e15[??N^
YLIBIV.Y>Yf7E_gC-<T_9agb1J9\.RZ2edHXPTVUMG#0KHYHK@2&>7A;2IX.X@f4
2YRbD+(RXH\YB:G3TA^A1g=c[Q6+)VBQTd7Z^90SIV08;(W#UH47<[ee0C(.S0AD
(\\d_G,1WONC>MLUc^)CGOZ+]-g3B3FcZWGb/OSK:NLfZdQ?d^g/3&/GFW4MS:WH
3Kd1cOeO_7MIM:V\I\7ZTC^VcCA)E(-XCK\4;c&=O?IZO\E2,/=Y@6_WdZ#=fV9U
DOOd:\UI>7,1<E\WDdcdE86T[8@Q\F5I^N1G,^c<K<aW=HP(e\U:<0bYM,:=[C<N
W>HTfJF=c_#6cgE194ONR_#Ade=FZI./8V]L;=4Oc)&6S#29aL=-B0G?DbP_-TL-
3dBB@RHab(X?&3G(:N(SY;?d;0#&Oe-S)UI8H79HPYZeR?3_=\DXeb(<T1g09aV:
.1/NHJ7=E,LDON1<^0gC5+(8d7b<MFCUK-HCOG#4T-J9^[ETS-OgWTRQB6aLScb/
GQFF@=D.6fVYX=g/#0_K02=0U_<P2_.T0=deA<?YCC>/bd@E)BX6;>O#^BGCU5:]
.6HF^-FC@bS_O037J<[<Cg5?EDQc-ASC;6THYcHc.SO+D5CDfc@>Rf[_P8-1_DXf
N=fD56+]0ZGDVII6,27J3)O3Y,0L3;5<aJP3>[[g]g\AAS_F[=V4aU-JX3fJV.7c
J]QIBT1bT+eB^GC:4TNW?+_TeRM63HM>C0c&W^ZeNP]MJXH,K?R.R3K2U;fe?5IQ
4M4U-IHaOe8&O+;7>/6&JW(YSUe_45<f;L4\b+E4DEfYf;H#/TCU0&\5O/gSX?4W
gXDA\U?JYJX5_909<)<Y+d5WE/CO3M>>F05&&YCRSJ.7U8SOA)Eg=ReU-W=[WcdX
b=ML.&L(1V=JP[e>=/#DZd[aC-6_3:677)EGJJSe]-?SI55E,1HJQ[#(N5;d0<UZ
J1d6;fgSG+.?L&#3PMKHJcdB+N78Z4LK1ZHf_4c[,]2#<B3X.cKI;Y8IWOPISO[B
U^3b32T/3ZP;7_C0+[-GRce8Q??BD&(=<4N=7O(,Pc.E,CJ2d4T]Mf[@5ZR(4cc,
BP>A;ZJ]ZONa=ROT3B5#>#ed/IY7UZL:SfYO&=9f/:Y>#Wb,>)FKF#We2?F)+ZfJ
[BgF:9WUW^/0USW,:\^H_\L^;JOJ4E_TPJgU)KA(\Bc#=7^b>WSC3IEb.U-K=N,;
.Q<RHb(9XcdYKSKe3,P6JTdE+OCBAGKfJ4O.>f?Dc?4BgTcRbIcIE3@1-HKd0=PR
KD7#AU8CYP/V4R>M)0b5.W(ba@<]CK85Wc/cG9Z5Z<H&_]\4/J3bDGLSVI7I:I3;
701#>ODR8Zd-5Ag1.YC.(P+a^&N:O4^g#\8EOC-?d]_=65?Xa9^b#GLB.0FF/;#S
[d6OUO=e?4SETAQO=:[:I@G]\,4]<7UL)>P3E,<>Y4?W)52S7SUH^.B4<XIFNHFY
2(7IU?Q28.:P:-?J8\JW55e,IB<_.Z#SW.fWIEDCGI]W#/I52<R9W[,\59^\M-c(
Y<JfB@YFXYY&G@9W@B,ZIGf;)c&NE(P,[ZT8e/I;[TA63:/+#8A^/O.,\.JKRB@8
.#f07PQ5:Q_O_9TRURU[J03BacZdWEdIPRN@N4g]G(f.Q_VC#2d&Z9F=Y/6H-2c2
>N8eLOa6AKdU,?2SZ1KcAU1e@O=gXR)2F7_La)XJ6/VRFg(S<\GUZa<&1445Y7\@
SUW^9KRf?eUdF/L6e4<0a.>+U8#D4E&7UT+4\-,^^DB4[b2/]ELEN&Fc.H0TJCN+
_.TM;JDOb,@+Q0ga>PCa^Q#275XbP_T)KKRbXZBX1;fb@cXR:KEF3KB>0,35OS-]
O82IJBVR)d&63&Z3P)=_WceXg#Qa5NM9NX7>W)):8fBbWESg;[#E;IK?P_3TZG0a
2P&:-Q4S&#Og7e,cSXK.G?1@bH[0F(=0Yc?H^DF6AA>P.B.&YY&(O9,@=?0GEH?F
B0YgZA607U/],S3S/S1&T2QV^<fa9L<fPQ7S,gIccD_7K#9Ida36>Cc77cJLf)PL
KQ]&D]XdR.aPU7>-AAVIed?A7c/19Y1cUOJ5TQRa<>cJ1eFD=.QWJ<5CFQR48/f:
_#,#aUVD8B-dONS\=>/c^BZRHL;5XE9cU=B(IP^?RA&-&L9LYM8&+Z8(>@T:AG]X
XTWUE5^./L<S,e<2fe]-Nb;8#-5PK2(,N>N;:GW/KGR8?SUH/aE90U9R(.7&M6Ud
P2@EREYUV[6FV0QC]TSG(^4]_8/Va+FE8IPUa?<GgE4PKPR:f+S_?5V#S\fR90g[
FRL5DE06)>(;=g-7b;a\74ZHPHPWg3+66VR6KB1:a=2NESN7@0#GE3\_.VC=5[47
<S>4)7T/_5g+NQ/36Y.0bdS,+?C8T9:E=S^I=+6YHf>+S9;12PV#D]Y&Y/@#&VLT
THFNJCeR=+O-NffITN)F)0@I===NQ[JZF]N(V0eb\28^[=#)f(W&WG8FC+8EFLPa
CV3HWCIfAHV@J&]YLXNSUX\BK4gaL[2,/N:V9T9EH)@AKe=aa<KN)>5e2IYR^\eI
<g:I5CIGIQLagAUYRLT+F,f8L^3<]_E1eO#[_b_B8(Ve?\6E)5P5eMHXD6,N3DQ7
(?\OdDDJ(UdOeZJKA<(Mf-aIU1]@G8/+2B=>6/P-29U)I9Jae2F6==QVg/(89Vf5
fCM&B=bN70A#O<:(#\^(7)8e?0L#,)7fUeV#P&4DVZS5=(=52TR\HG7PMg8L&Q#-
V+NdR&NeDaGN04MRU^?e8b^QVDG[)Y2HE5<)71]GHH5\F4;S2KUO0P8]PN1?cFa@
F27GfP2F2YEZ&:Sb.C^X,):K;3e3Db;E7Y/R2(@UbbI/8:=b1_:)3CY)-VE;RH&Q
K,ZYK.McZ]0g[b@g-U..>fQb^)3(Pf2-KDDI0SOXdU]A[D&a[YXd<///]3g?0e9N
J3.c_8<WVZAb(LZO6Y68R+?42.,B(3F[@P\O8d<ZH.CfF)O[<8_Q81K?L:C(-A(X
\]3+2N4Q(C+CCAJ\cG]W;_=Re9MS+T-Od0f+-PRJ:AdbKeBG//;W._Q2F,-^b.M,
AHC,C.LCKKaffc(4XJ__99ES\KPL1O=Nd<#XN:;YZ^;VbfT:)g=6,Hf<>5^=2^Q5
8(C7C7K6B\](=WPc[eTG\1cAAA;ZD]UR6:7)^EL?Vg?=(G;X2/gV6e_?=WL/L&N:
HA41]HE?:>:PBSGMGg^cRZ7Y<?Y@G40e<aD[GO&H]URRGN/PdH9H)5YMHCC0,IZ)
;U?4;6(HSaKY)e4fP.V:P5=1MKZEN?D7/O7I1?AP2S[PBaUH4/A/;P^4]P(F=,#\
MIgB83J-Dfaad/4e\;V=:^3-25JAVOKcP(OTY;[VK>>^E^#>C27c1D&@#)HcECLf
W9aOaJN89T0@4[e1DAN@2&94:(JaOJDK6d/,<7CdgAEF-L/4fJV8KdbV&PA1+87g
-6283f<==c;JT96g+SXUD?IdH-I)E0OQN,Q4S2)A,?\;=Xb;e&KA5J#JcDa>89^.
4cQZefI,?J(6SQJ2N:3=AB5A[450ET=1T9T>5__]<Vg<L/:RZReZE1FS>M-//>aC
a:)&6VYL0U^P3a2_0TV>]O.fJWC;@+[dQY[7ATe2dLLeg4CBb=G?AG<aUOGBAU;/
@BaTVM^(,#Y1IGVVf,@VDQEB(NP0]fLIc7a,3Gg;OD:Ae\FCSJM?FSXY8)T(2fGD
8;3UP+dBc&2U4S?4g^R\WMU5EITa6VUV5@6/d?_]&I<>(6.HGb:IN1UCE/Y/+:VL
G3aG0LeJ3DW-df,8bgadNB:\>b#M4_:eV;NFfA_VFW738^QDc_:(-^cB,\/DZ^Bf
<_A447#PNe<CLYHW;RQ3^YM_S/bcWH5FVFRfIAJ2,=7O,<5W++-9XE>BEA9A;PC@
F4:=J@gBb=2Vfb:ZZCB-AHK,.U#9OYZK#O1+PHcd]Z]J1,URPO&1\cd_R>;19a6W
bJ48HeO=bJXU^>91>&MG1eBM8H57I+WEKT:H@8e6GB(;I-GMf2Q,RaffXS@01Y0V
CBS)>3X@J.T&g/bXGLE934&aX5W;#bW]B;#G3E\f/C9QX147@GS:9L9:HKf2C\TK
F[8e079XQE_SWL?XP2OW@Nag#\YD7;1CMZY@_0bPS-CeMO=(GTU9W)\T]D:XJ[6[
&K&8GKDfUa&H@3K5ffJg;D>QZ?)HgQN^G\=]f4;&4R;fMF&3_BQ]K]9YfIV^O\3e
.W4CQ4V@NL59PE9#91eb81P>&2>:9ecJXB1+4K=Z3L>JT)Y7(D71=OPL)N[8H,NP
Z\4ALS,AgI&BgZ18O#cL0<SddKgba)DH42b(PS<GA4[CWa-=W/-Z[QZCB@cQ#eFd
dOYT07I&e,)G-8CS#U.]1(Y<bfL&IGcZgZ;dg;2Qb9&5F#2Ee:.D9[7fQ2UQ.ag/
[<WL><?4EJJF<?W(F>d5G.:,^=9NT<4CI2B8HF^>M^5JH+b#VZAG0ZRTF0-4XK>E
-[G<OVFKUXR=ZaeFZM-X0LVZMK30AG<6;IU-,EZ^8(/J6<8XOgTLIDK7UB)bEcN2
,3TXM9P.U7aQZA,A6HGE\bJ3?N2:CGQAR)(>\f0CBPbDQ@/Y.Ec@c7,YKeHc.^dT
-J/419?aX_;1U<\;XBSOJ^J(P;VGJ^>O:ca9E&J-4aJC?,_PUA<Yb]<@;;CO?aF<
\]+[90#O_1Y&C_&6RHS0A\g;,DgEUVE3F0YR+PRKZb#L9R-Z60.YOW..d5??^1DK
6L-9cbS#UTCHEVBVQ_&9D@d<-Wa;I#&ZBZLHWYT4OAYIM42AAQ:NM+&RV&&P3ORf
EZ5+bf@Rg-G,?Y^c#eBM:@d&5d)Y[SWB)<][]b=^X+]B5&C1,f&_#eR_d,3AJ?P3
.84<B6gJf86<W.E+_\g;/QV)4]8bcUefD=0IYTM:HH\gV@UT-@_2<?ZSaSe1.(I1
JX:\+P^\NVg2NX6F(38,[fF,53^<85XMV8:NX0O2+:0LgZ6FS(_]9aF>B/C>fT#L
G??]WVL?4C&J(I4&K&2M3VQW>;A/QPL&2c:>,-&?@[\?>Y00[S)TJMcac^:C;Q+a
C;CX/-Ne+g#d-6WNdbJ>Z)IK?bb>g2ZR,XAb.J>@_<YVO.+253=F>MSe=(a1KX8M
S=6[B;V(M;TGY+NZ(SKda#U@5Hc1MUdOLV7@:gW.WW;.(KbLC9FP5<=8Ig=W6T+,
^5?160YZ-dDF1Y1e1T:D6?S<DBJ_-Y[J51\UZ,7PL0Q\4_J&EbR/Z8Y[CB4N-7IF
]P3Y@:?=H3EL.>Q21Pb5fXY&P#aBO5Z>08=SS<)&d[)+A8]4-&J[XG[bEBY5_,92
b?[-)C)+?g)Mc&3Z5?ODeY\-Z4_cdA\:Z+OTQ>+M&a6WIG#MSLZYbaTfY1HdK42C
9Z@S5A]-(OI:B>CdM1G\7\7B<fNb0S_<Y2fEf>UAPWLL3e5R?_gfW,@g@]EV/M&0
Y(.YZNIYN-Z;]ENaTdb9;gV1QbbEQ,1?b2LZF9@-=V_9M5.95Nb0KK\a&O[6aQ1,
#9e\?QSFY8Y:&PcLK]<X?g##dd-#a:9cK1;07EO1Og.e9.TaCBGM-&Da.6F-,F(E
/Ke:ZF-/T8D^F1Y0&T#BY)d70@KG@V@.E?3a@)F9-6.c[27LW,a;H26(\D]b=HHC
FB<EF^c,@JBfGNN1/GYRffafFG5+gW=FAb[Xa7PQfU]8ZA&bM0L3b,&fSe<ROF2:
0-3(L=JJ@6O=D2UUQ3^;+,6MV6^4YR&/AKe\^=PfO-ZLJUR)^<>e#e+,b,_<-AN_
5K][8X(>9=,-49G_W+;/WXI:A.WZ7A(_La]Te>_GP))dIE_X6(HfT4XIL,A[Ad(Y
.X^X>53I3+cN/_EF,S53:=G0_F1a;>_aQ=gKCBBUeZ/5RXg;-C_fWV=OK0dTg<gZ
Q@WcUP.d2]=E@0#48=(@<\>49QN&^HKgNF20)g0<IZSf)f>J[+QgDbeB6(]AE@JT
M@I1e[Q+U\__D=\CK#B>9V_FdT+LES\CM0=0ePK#/N3-E./)[9.L>9gP-fRQLa3+
C[1fH23YX]EB>^A/Qb#f.540^aZ@W]a1P9UUcPbC]DEeRK+=\Of]6f8cF>&KIL8[
Z_SS#41TA0&-ZMcGA9DJKO0I.W_(AVAZWC=cIL7g:Y^4g=^Q,e+:T)68;D58)IVW
;0(7g)_g?:Jd9<+JS(fHPRa-S+.[R@.VWOf3@E+BE</A)+@)5:?DH-MQB_0aJcV_
H:,9FQ8LQ1Ga/?L_94;4S;.._?]8CQ@;E2#9\bGL>?SMVH(,77HgO?8M7PS[1_;K
a9#a(#JMg>]8(#b5W9b2LZfZYC7,3+KWRHTS)7fY>2g_HHJ0c-C-Y-,88g<fY^&g
TO/2,NEKAJPPZR07d&L#aI5W1Y7QY=43<<:gKA0^.)]:>RAC>X=R6ab)L2+gPS[Y
[gL&A4Y\8WI(L2K_NO95aDLP5B\e46=]I4^)>1Z..F6RTJ2T:/2SQZ,Y#AIa1[_>
XdER/TUeOR)V9d:AL@6=.(?[+B+U5GHM1-Sf?F<ed=WWB0/SNf7PUWT/A?_1B#1=
e,DSFAbKLdGC#(F5SND-&2/B4Q)b8#\@@N9,_D<WB?Z50QO,C0&UX>^(f?a7QWg]
?OUbO2Qa++)=9Z.<PbH7d4NCNLFRgY)R@VV+S.F&cY&[Lb5.49Gg5Te/C/7gX9L)
ET:TB/-GgNK.FIJH9+XFfP6P?6=.K9,=:AP\]OEE[?2)S8KD,]4-PD&T[f);bJ).
a24@@/>P&dW#(=TO&c8<.U2d7D#?Bd2BC.X8[(U3e;dJ.(KO?(,eQ]6QG4a<3U_P
6ZUH;80M4g^C?=>58X2D\DND@=f@Z[H@FX(eR:&/=I3<SM)RYVO5HW&V/eBX?K.6
-XLH,E::fb:MD^g/g]_>eZfZYF-(]3C:N;NFK>[QUE31UJ0GRFS-ff2VWP7C-OZd
YNUBHF&A/d8-GMN,1C0MAU4+H@Y_8XBb:^P?H_PD,dV7aA(H2;QdD<ERAIdXQ[JO
HTOD1&=bg?[WPA?#c_\(XJ7HRSJ]Y@]?7^b-6CM\JZ@^1/Y9&_#:;H,&Q2],I6bT
TK2-IR-V136,M:13@eXU?9c&.SQYPH8&KR;KJbLD8TaTGd9U<KEE/I(<V#+JY7A5
A@b-H2=b;D.NCWcRGK0cO0MX3WK-9)Q0EbeUCRLNQb@UR,GK\bDd9BO_9Ng<c\]R
fGbF0?e\2\X^#G@g:6.&(f9Xc7OUbSJ];]#abgZ?Q67+TaZgH-N_Q4=fSZ=KD;ZX
HTb(]^Y\SE7)&\Y;96T8A9fM-R>H.E]87c#eF>(_?b/G5e6LL[ZE89V.MdW>1He0
?^6<KO)7^8F5dQ=+U#I=PB,VHb_4a3=K#26KAU,9#9IAF?LL7/Jf^VG99>>f?Z6/
QZYB&I[.YV8Yb3]^YYOTP#VJ^SD]8[58e?W)UT[7KJ3[=&W3a.=9(d=(3a+C9cCS
ge5Y[>U=N@;b4[Qf_(5UPC1<)MAUFCRf-NcQWPK&1=337->1f81/\2FMZ9=58#aD
E1X[f2KIfI^Sf_1.HQbO;bUcR0UYdTd)CF#+AJgJ=ETMNJ&@GIA)1gTc1+Da>6#>
,A+5-;SY#U5g31KUYQa5S\ZOA.D@b5-]EZV[YFINb5XC?U=6.EF7MZN0e4//[L;_
B+36-bN2GV0\W7C:\:W&IC2eP^)CWP]Wa<3gc_F^SeZa_SK.gCSP^+98e;=/EUH[
N&bg4+0<dGR^UcQ3O_5^>1ZD1M[g,@^bXX]WgZF#T=N_-VT-Ab2H+<f?AZ@f<SOL
@(\#MEQ>c#d0d7<.@L2)f@GXe,f]5Z?CWN78[gZ.82g@B5SZeC<RX.ZNC?U9Oa)(
).4MQ(MSXHS+_BdbU#4@>5QJg=W]/fW3TY)3QU?U6;U-8+H=f7Ib-AG0QcDRL,KX
Ec-gbd[:I)Zf<f?7QS01:Q>1IZ^\4,IWRd<>&57N.4[V7-K9>PcGJd>#OWH/aK0O
9d25Bc6-8,SN6.E1?YIP7IVVF\B^AG:D6_0G_=^PEdIM>#,TH#:dN2c<=:HQ#:T0
,0,R3M_MOF4=dQYB>1M1#1[+La1/QeB<4N0^J9Q+-E_A_X)7a5W@J.,-CFb?74KW
ga=VCTO]8]BEd,:@?=/-Y=3T7PQPZH+)1UWcK.)_U.fCI?\8_-6eET4@ONb9,<cd
5fW<F0e,,^_D?2#I?O\@K_W&VR_\;7b]UaL)Y;,Y\4AA==9JSbTY4<MJCPfcdKJG
bDIS4J+d_d=gP_:VcTAbceA+.G\gS.Zba)fO5N<(7+6=GeM3bY]CAZb?eH/R/^8X
+6[SZRN+g<&Lc7GN^fH<=2^3)(f]f=H<A2Q;3V9g#JW4c+HVI<R6#bc)BD-ITFRc
5@7/f]BB0AC7#3Q1BG<2X7>A2;W<SG1SDS]=[]U=V.&],a\PW-VD>+>Ga2OI(>e[
gWW#:NP;>40Of4-UH]S8:A[\WP<K[V90[dVAQNWY\</X^]?TYg5I5WcKK\&&IK8T
5LHKVaJE-R+<_XS)[3;b#9O2f,/@5]ZPGfD(_R<?BFE\3(FNH;CC2)(+&])_H9>S
I204eeHQOAGID8)Y[#OJ;.W,1^Kf^W>)RS(UJY-EP&#:6P?:E.SD(?aF,/WN8OD@
5U^=HbP+F0KMLI]+A>CLUHM<f+dQNbA,7H19Z@N=DH,#02C7RK^H#9_FW4M<@P]c
WaART&CCL</A5P0-:TQVJFC\K([;-g.H,829dTU9OEBVP<B<BD\A4\C@dK<C@PDW
eM49GCfO@O9:AS68Na1[B@,O\3;RF]RPSc3a>>\IE\L@DE(]&R5KTB>AeL;DJ]=e
X]g+SRfDbKAc5eL,b774E^/@P>PfN:G]a(WM6[?HO4(VFTE6W/@<#db>)7H;,7I#
f,,P@GJFTd^b\L:(;-U8)(PF;HCF#2&GEQ82:#5H\GXV<&FJ<B;V[df/RAb:5Y<_
?A@9_.5.:;(]O39+:c8YaPZ81(XNa:;d;@R,]WEY7>0g0-XL&\.5OBc]H;^O1+M(
eIQ>/[Ve,Ub(3?gSU(Wc[VDZZ8=+gB5fP;,A\A4:J[CeIc(d<6S^M,K[4A?X/:I_
RR)65V;0L;Dgb(I8M@WGI9@[D[_3D:c)V;&OZ=\E)(a0D26Z+-Wc2SC>40bAa#e>
)LILR<7GAV-38Be/Af@(6JUYPd8K<6ebdSb3YccV#V(RCV^dPZOgPC4X48?/5fNX
NHL3[6:0d^a[#e^F9P=93B(Hgg-.2g]AI0#=_db4/BKU3O&cX#gaXF_f9/=^JQQN
[QGEXKYD9c-85_([_[/NX?aKGX27^(<(E?,#A1W#YKSKIE01gPPL6I410W>ScJF,
A+\>44bR;F]e/]gI_VB?^^R/-b?&WS]P[J9A3]MXIT((cAWN&8bDE),(-,PfMTb;
69#^Z,aWe:8WV&[.8fV<J2/@ZCX)#U79\4@.QHd(ZgXd8^G;6+/.<Dd:-_L9c+Fe
X3XTGB=3Z&PW)4[#3QIRR_H2@RWI)N3Z>QFX+Zg>S(bQXE.9b<@A,#>R-FJ#U,Jf
5Xa\2U8@<NF?^+ZU]<Z)JabU6d^<7SY1_6V^Wf5c1&Lc3]DCOLZVJF[;/ES_^AXQ
(8IFT,+=G+?56HUB1VY/9[-e[5K_HXd3KO]aGUJ:d\R9:,JGA9FX2;M-dX^[EAJ.
ZR22b7LEIZRYJa+L>82A2OeC7IfEAaa\cA>g3fF0S[bKJ>D0B,=[^7e?./4JeU.[
P#6[L(26.ZXV\<g)^ZX.U7[^=D6I?1T7-:5P,feFg2ZDd4.S]-,2VXX:84TQJBb,
[gA89/ce_.#M/,SId65EJ=8gWB&-egL?E\RCZ6[]C&@Ib>8)+W.dYG(5481Q=KMf
b-SKIA@EFS?\C2EFeC?(H,F[;T/?GSGW]RPe\B3KfYc.2>DZ16](IEM8ETRa@8?,
eG:@.WI+H:F]VN&HXdJd_\QU1?]9B#<P7QMUGfXU(FZ?9c^7R5_HaOWN:UC,V<.+
DZ9IJ?B1ZcYWBD-)D>,]fKEBf)[7SRWVV=ZEdO1ON67O^cDDZd+\&J.08=F,aAUS
a2O4\\0BQIN1GY@,2]?58AD&1V:#Y8Ua4:I>0UTfO+M^]6a\gD+K\GVOZ<FH[_1L
PHb4M1IJRM#XI9X69SVR90BRA4;JeQ5JT0aS8bEGR/F2[T;1;5-9?C:,H4XS,)-\
YA_XD-T<4KWRB.9Z5+9a76_c0(LcB:P1Z&Wf0,&_)D2AM?N]68-9)a,LN+P?D,CR
^C7T&/-@\]=\c^HM>cSRA,-<HKgU;G.@&@c(.aBY^<>=T=(6G;ebfbL7_@.I<b\J
Qa12:1S:BW2C==G?@?@EYZLJYU]1>f?K0Y]g^Q47Q\4[<M\78eJU7+&P6==.a5)A
e80/>d26((5:AR;;PP8OLeISQPR,OTO<:2S,+.YdeSaR])2aNG<D(=9-CJP8N?D@
dK#Vb4Yd1RZMYCI=3[TJ48G<[.XKFMg^#??XBJ1aH7Z0RcO^LAcCTea4a@3>,dTc
B+bO]e3D+W#Gg^/7WC(d?S=gZ\5&03H739YS[K?(]VQ0^-7SWH)??MHY_ZgH,1.[
OgB-f#BK#B3R&^Q1T0;^=>NFO+;7b:])D1+5f0Z.ROT)c9Pf>9CRZ=fScZI.Q=:3
fC^>a.2_Qf3+[B3/9^;[49F]@6?1e[<,(P-J5P]59_L4V4-:&Ab[#R62VA-U[Xc>
0U=fbV6K+c=e9eMP)WE@25#cab1411G&BY\F;Pe2&S3#;])ID]gGc+0DM8GS9\SV
Ob/g+:I-f<a\@^9IUDO#:0S>-F;a3^BH6<J4)H.MMHCYTRd,E()aI]:K;.@&=bAG
W_Kd;E.2#,7<FeU/DQZL13Fb39]1.O5F5eHH0IT_SYTW<AS],)/^<8,,=g94WZG9
\SIMg9eS&O+gE4-QW>?=<f#?R7\Sc6:NXaJ)a@TE.N\GLK)<[&BX_4XIZYIPN+7e
7X,)BS3+56PD:2<QV>+W=(aUPCA^^gWN-BD:>>3_I;RESH9VYG\\:cCZ<R#e?SZ2
^<H2/N^)A4<dG&I9DK5JcKMeB/f\0c+Bb,L)K,UAKSe+=e^)\.6QQ[+=WD>V]3:f
L(c,d4QSXb+VFD?<LbIEUe)X5(C+_8a0e[+VK_#;Q<2M&fSb_>+bV6,JRZ@)RJ4H
^ICX)Y_d[_]P[8..^\VXLMb^Z<BfV<LNMWgPSH]R6#)Y>8f)g&dSXWG2DWd#SH#J
,J0VgXcQO0_CV1MB?RPB3]DD(Dd3]2;CFVHU[^1+XV4;AZ^dI6WYM8HJOZCOZE+H
<X_H\BH@]\fU0a2#dC6-U\T?KBTFXN4<5bX\Q/\)CR(0S9JJVd6UM=f7O8]K2BMQ
F/Z1=IXa?[(Z]b#Pg\GZdfKSK>?5LI#7T&]WW=M17Q-^4U.^T_V7OB[4\WW(V^@\
:dT.&_&_-P\9#R^&A5B2OY5XQdF]UE194T5.>I:Mc[^L]TfFM.aB7<(66#bZ7<TX
ffL8DIT#eFcIY_S?)&LHaMT8BcO0/c(K5D85KT(5JeSAM6HQKK/51=#DD>G;6MR&
BC\XgfBddKaRO_J.9V_a>ITa)6X-\VX\.a2I=#R0b:)1YPcC,_MQ_I4J89?GIRg2
#AQfdX+(1a_2ZG3/\]ENKTR+B3OLZ#Q9?5Z2d1#CNM/C;#X8\4HgdAe958922UW#
V&#FX.88\6Vc\a(.c6MH>6Gb6^ZT19CeW#Ud6P]A]fK#aY6@EEegQ.N,3HL=?fKV
f@cZ&B?97OU1g4=/2-g^/D_-4G?-CI])F33SLRd>dC/-5L\_U)FRLgKGUQC^P+G:
(bWS<&[NE)YPTZF(8_dNYN0FCD<c6]bI[/H9f.&^MACZ0b6c<-E2gWT;bT/PRRNA
48<JbQ2c8aW\HM/9(-51_0D;F9/0\(O?&K^_].FUd<T&0GEOMK:Y<+<?1HZ96##\
PgR1W<@AcEUg#NN8=U:DGKc1/?>(TLJ0L+N(NU>.#eEGL^M>e.Jf_34Z_-f><-3O
:);FgPSGRVD00WZI0aPAb#,(cC/Z:J2M<T2f#BdZ&(<)?7@>L;g)d..,(If/1S-J
S\KS102EM:adbc60XJ5>+/eT<=>RFJ-Y=,A?38eZ/deM<1XcdCV?29V@4-d#5S6T
)]8CaD[&U3c[+/fAJdUc7]\:KT+g8:GeMRg<&O2Q@ggf)8<ZdS(82@IHPI2PRc\E
6;=+Z7C_f40HLTa:G+Z;DAOg5M1ff^4?6DR#;8J]+JF(BGc;N]O[6d@R?LdQX<XX
dL_-A;/GbHK?dM7CLMK5f>8>9/LJ>XMKJ6&R/=2LJ?5\_C\&@R5:Z8Q)f&1HdPK=
?S&.,(#C4GQ.4J,TXW(4cc4KNH95BZ@8A1R_L>LV\86cc-</6C)UY=Lfd7ZQfFAf
0b4cQLB&I>>(NJO\-fBA\(ab^b/AO#HWOGM#0(@f5I/IZ-A]U3)?Y-H.Lf<OH3]:
X:8-b=<.JY;MbJ9a+8PPf>K(NTPWUR=S9\C])-^D@H+]ZWV]\U\P-O^E@(#91+Ud
R4V2AIa&S;AX.eBZAD;@BQBS752+<+U,8LaI=6(Lb#O_A//e22NY=WCdG=ae7[)0
PKfa.9.cbL&WOR^MH(1;?<E\.>c]5f=YD?[4ea0P,d8S2:@<?0+B3T?UNB<g(3BV
_9gfY[S>JX.7H7_Wg3N[>W=9^^QSV1cUG,G>9);HLW/+Qe>E+:[:8IX:cb^A0;Cc
0da+.PE_LNGVg]>U>?8^RM+3UA^,Q?O,I\dG#XW)J0KWa;0Mg;.\,VGR92HdJa8R
_BaR73#99:KOCZf2XE<8U,4a&^B.R;gd(YCXN[^\-5>FUH&P(dU;_9gO/cT-TBM?
]Y@R;^Q^G4IMaFc\CQA<d#0eF[[?X^<aI^b?B1#CY\@B:=K+aG5VQ:1[O@^UD:Z9
F7S;DF9=?g[O]+<IBJY+;&W<7b?6--2/((.1d,VTfWMN]1JL0U7405OQMKZS;0F4
/L?T-/7(CbaWTEI\=MZJJ5>J&)4O)=FFNc\J[3Z?4Ec[?.T/-XVN<B>(cMcUB.HK
+NETNB(BL0LHfS0U;UI5,aD5)8)1\LLaV3g^NZ&21BB6S:FYA_\>5/bXCTFQ&18I
V7)TQP;;3?=4(AD+=V[XZ<aFB\5#VF253#J@g;^f6DS+E@XL-\M6I.-U6F90,1IB
_5#P&Ye:3<7U>:H7IcACb;EPD+0SDF\R/++\)4GWT4J#K)HXb496UIba22KT=fLO
?4[B:G\e01ZDHd@X__.__(/MK<\g^>H7/FEI)f]LZcNI(1LGY/f.[LLa@d^QA2IO
OA5S7)+:VV&BX@:6SJb(+9:>JLI?8ac?06L59:C:BF>=FL9e<#X0OG;.F3g;&X(^
FQLUc7)6(WWY-XX-X6a75:e#ZXe7U+:V[@(=_>Q_2N,QZDGSc<^A^)PaH3HA/4A3
UP8#_CVC2K_JW&G9-bF.gZdU7c;VBZH(/OCg7I6bMW0D\eUg/@&SAGR74fI8K^#_
<@gV>cEMB-,\>/g/37&.QK?@_H0QNE6eXKbX&@+Q3NZ4Q/LETfLFI/c>g#6V2(TK
>BTBPW9Q?a:V<JY<;6[5<E?UC.1;CZMB+E@eJNOSM9TBY:H45,b9]DJV>(-B[7)3
?[S,#-2Oe-f>>)KM=QO_X5IIPUI+bBH;B-GM&ZaK:J^F4ZbF:(4>=NY8S/Y/^E\)
5&R<@3cK4e2.DKN,3Vg2PX0.Nc@5cSI^J5^ETX^L/E(U\S>?O?<CIe2VcHX8X-5M
9YK)X;&1Q2MJ9Ic62[TU75c_.\G<]:9VS9R97FI8[(OE9E#Rc5\3)LD2H/MWdF9,
.gX\&N?UU5c^eQ)5EG->:L<?&3XUNVbU7FLA+d5.LcHA5g0:23O3g,1)?Q:RK2AG
:N@L4Bb-8++I+KFIg4Z9>TVG,((DJ8K8]A4fZc633d@#Y9;Zg6<P_f0HdKOS/?&@
WX;2;5J0TW#IZA23S?7/BWP+7:G)f#e9BV<=2R:@7]WA[6,Kd)_#:-W;GCWKKBe9
17<e(W&GVP-XE+=PF\??N?K84O]Q7K13IO_8EHZ)SB(2g\0YNccN,SfG2\.<],K4
&29.?UdO:-&/:E.K7Z-6[=C0D(^07)Z0WJHC:;:B<KK7K#PZIRbXGY(P.4OZC/)B
fbER55VSg@=\F?+)cUbXF[&eb=PF\<SH[MdSSf\JB=W(cT1FP+XTDVD]4I<^35[+
2XG=N78-Y08e0Q-RObNJcdP[GY<(g#,O,?R50WB>#QW:@0O=(Yc3WP+<Cd^6@3->
Z.)[a4BNCeHf>)ND6>f0]/,UBdDGG27@[Z46)^S?8Efe^@<6<1e>GL,^K@9[eCMc
2T@.(dJ(YeQAcSZdK0Y&QZ@_@I^<;+@:-)JbGLT-V36K5a_Q\Ca/@c>Da?]5F1BG
;VS<(@E2^O@[d0L?/3#cc7N:&6DFBJLL4I2e.8@0<\AQ3;T)B[\;_36BU&KHb7E)
0T1f?4@fd6[>5[:>AFA7.YR(e;FOV=dgZbd@(fXW<)]U[;IDWL]NQ=,@Oe\BdF=b
2<)EMHKPQL)6@fNc=9(VeQd.=^2g)G/O=H^JW=a-U,S(662YN0,C\4-b:9?a)P,;
a6[=GVY/=RBB,a9Q1/=?,=aQbJb5]Ed:6[(g.K+X/cO6fO+);UTD,^g+R:O^M.R1
cEI8;-g&-bd<LPTWPN2Z6/_GC,FfI8#6G?1NUNO-Y@f_V6VSD3YUH/.HbIA0Rc+6
VI@)YXZ#Y(JeA2R44f7\&ITbBN[>B-NVa<3I5MH[-8=Z)_.C>@PQY@\@eTU[PL@a
OTbVR>6B4&>(fC?cDEO8b(VM4DSe-4X.c527D5eQO]^baCFW-#KG2_50Ab^RM];A
VOb_gUEQ.,B7V?:9T@3#<GTae]KaQQ<a;1c^FUVC6(<HU;W9O.dL&2X=\H+W?5^Z
fYde3Ng/[[HW=P<ER1E^2^;:a:8G,)AKT#9XE.bQ#.GNJ89dB:MUXAM>+)aH2cS1
4?CIEa:3XK.a=)Y;>_18QO;<U\PgDc1S_WRd5M]#4+#cd&UO-8LJTA\JY@.HSO&a
]4Z&bQL1K<:@Gd._3[U2/UPde+3)bYAY>Y/&K/4I6_V\aF#6b[9ZZg(0C#J4KaDO
OSSf+&Y\3\-=E]&OU>I&9\A[;,#0ZgBT1Tbc)I(5MJ<@IT7AW.e[7B^gW7Y\B-<5
/U@A[?=O+#efBfDA;e@D+:XWV_4CJLIQ^^cU?>C#G2#:4+/Q01P8#)e;>;T2b-gC
@aDc?W;,18#,?EN5fdG_+CW5b0T653LTSdWZ@Qdd_+?:G0\]IXc+N2YN+XVW>J)^
]PfAF1I@?Q?f#F#&:-SI;8HZO#bAU8NaLUC8=_9.;#.K2><;6CSQ6=+/8\0S+/bQ
&@d0ROX9\4bY=S>,ML><5IH].Nb#XB+,F(XWV20g]-dN8+SD]HE6>_>8>bZ9gXGG
51:4A/-,;P8.EBN95dC1MI^>FSY+1OY(RE^7M)?K8_#Mb<f:R-@LVY<[./@^R4Wd
QgU#,Q?f)]P<SW<^e3B\YM<SG@R.B;/=9(]E1XcVF]O;RMe7]&[6+E22BHP4:APX
ZD=:(M=)G4OO_](H_[^,V\K25GC,6EN7EER:e&dP/FQ,Zg>Kf)T4=6#Y9-<CFJ+5
A_/YbF7gT>4b&Q3&\.cDC+C/G;W>Vf9MdR+4c@=YWNG>?aD/ZK\RMT^UDI]dH93&
-G^3[Rc-/TY5PXLb3\c1gY5@AIIB&<=J&8=\G6BLT/Q..):@7>9c[,EfHW@d5@?:
VF+KaY0^GRH)I,N8DX4^S.TFe\0_HLHD4Ub5F@-.BI3^61Q>T@[RGFcG;V>TK:::
Q@VY/F/^bAUGaILfD=R69\aeJ7e/7;LS4?-#9]LC][B=I2-DIaFg^691bX.HGEV[
Q^3-=WZ]8Ga7eKY^e:I@b6fW366K&fNAO&F3(S;;?Pg-7-cW4;KbM=X\S[9,b98&
5cWS<bg9&M5;=^/3G#E;/BI<8a?DIQT)IAKgZDZ13c)BJOZ3e:,DFa(Cd:Ec+P(b
-B.WZ0B&+PD5_dVSELd6QT3U0J^)_2QP#5Q1999gME)9CZM8()-ePCIWYRR/6ba7
X,#-BV_OTb:.g^HHYbL7:OW(]1S,1OTgJ40d2/[;8Hec)dZUL^(;PQBIDDF_VL2;
^WJNA6Ig=Z#E?J0>FHeWa/SS+EUfR7ZbNeO>H>1I89e0CUKG)(#6AS8S-f>0cbPS
83CCbg2H=,@M355FCQBBK>D7W)bTVYC-Xc&JE]egTR@^Q<TJS7MELgR1WBIB;e#\
7F.]1@Y(Q)Xb^(:8CMHD#7N]:BRU+Qf,BE3OaH4HPD_ZeY]gDIPR4J;(/.-ACZ7P
/g&-CD7>a^V.YZ?&T@;00I^:\5:]dZf5,[VdY3X,.aSee<N-GaY0&&K2fYMAa67a
\3686.]B2CH0Y<IUK_U[OV)[F.=PLCV44/DZ&.C-,f:e+JAd<T8_D:V^Id_+>#_3
EdD05Ae\B4YaT.H)EJ&GdaBD\9geTP\fL7Z(FN=C<EMI_^Yc,W#XF<YXR>c(>f#?
0;ZB8<00I^,#O8N,R&C)4N(?:O&8:V)f4C<10S?CS?8/GY^7G.73311#]CRZ[d;_
8(ZW;WX^SZe3[5[KU(#F8X-+F2GYN)gYJ5/BX4H,^V<P/M/T+QI_:VY1EC]E8<cd
[U2QdA;8AGMF=#+0]^e10d/WDgbdCZ?4Y1<](&[0ROcf<C^MZ.^ba_?\CKUafcL8
M^M1NeZLJ#FL>(+b7(B^]8LI4aEWNG51Y)K&785-JfL)Fb(4(5^BL8RO2HT#6(Dc
ETWL:B_=FU\U\e,VEM?d9JPCG?L^,3J\L6REJR@FMMJH<ANb/gP_4&S5-g2+d7#[
O>]@)6P\dE@IM<QU,d2M6B;^_bK8,W7Lg\Ud,#/+b7S3,a[)c_KW1N?7()QgaU4\
K,C@B9CWB\GJ.^DZX73C.(/BJ+(&DF1V:^>)9<@Y.>+NgbQ,;3HT+>O].Naff]5R
4eD900]6Cb;1HWM>dYUJC#aT=9AJWa]-L8<=6A:Pff?O#WN09\1@6YagAb&gC)0b
WeV1P&g;780=[H?^=KdZe4VN,,,TL75?;#I@Ge?=NZP]-&=0DP-L+bV;R(9A)[f-
/3QN9T.]H@EeR09A\G@&XTR[_Y>eS?g.[1MF^W87;d\E;(U[:c1#U.ASW;_5G?04
V\4>d@2.N8);-?##[]J[0+0_fQF[bW@OS=K/WRbU=93fK9KQdRV=Y[DC@K)=6\]g
#390U,5T3G@0aEg6,RdH?VQB7-5g2f(9=.>ZXCBG.edMRWSZB\SZZ5ga/PW+,EG[
#@(c7dK+XD>UJI&QSO4KZ@[7aFC9c^\OHHS2_dTZK,,dO_de.BKM2ae0bO/F7C1d
I@29UMY[+eJHP28AC?M8#c0<BFCTOINB+G00&JI4M/]-N:Dd/=#5,(>e/g,2EAP?
-<CT17X0#b;+K0)=;)I?F]V?SF)MFKaG-c.OAP4LD>HQAa?&Sa@U>H;;^HWB;PB8
4S5/QP=05gW7?V;fQ:GWW:c=9A0@1_MZ5f>?BSZMd<N4NGS_4a:).cZfH+,]-(T4
fac.4C,gObY@PC+BeWJEXC@7=@37@ISH&_[f6//VBOT.ZQ5LA(3A2g9?JOf8:_NX
XXHO^]&8J]B?eR)@K\f;:cbIP/K@degCJ@dNW>Y806KM?_32;cff-6?)CXXCD0=C
FXL]A>.R(Z/&>M5(\>ZEbD<?<8:]YM58L9Ne@gD5:]L@VNf)/K_&3I:,If09209D
1N.^RZ4JN@<23;4,QNK>d23;d)8QX:=;7.c=:E>I_H4B.;\]06#@L>S,DGOBK#/-
L7RXd111AGN=Xe)YCO#=3B4fdegG0TV[eZM6=J9.B97B_=XC<+K-d.T=89,]AS<J
F.6_6U0S:&MJIEB)LP]L#1(-^ZG\gI2XDVF;?dC.IGU;^RWSN7U;NgEJZ2Z^FCJ+
ITI_VN(TUHHVbOecf<-@;FYWBVaO]g;YB+>A)7&;/UPg^1HVG6,G53<gR<OSLI(U
cLX1a<d@I?[)Z;Pf]F>&9A#0:8B/1UJK&Bf6_a5Z2:bR)#RWTTfQP>O^(VDRNO8d
PB=DD1OF4=7C2d.RD@5YYa5@4[(>7.KS0IQ\B^SM8YAXU^c,,Q:\cQ\S:4dQ_+X(
3T2/[04N,bSc9d)Q=<6<)Z[9D@=.Nd6>OEY@DURR,3g\(+;20],:-DL+[g/g^SVM
&2bL:f/FF9LbgEW-CS12;3I>DD4_BZ^XfUQZHaaO+1#c9^df03\.3)K1VRTJ^RFX
3I&O6_2>eCcH<c.K(8f?,SVR<f(+d?D^XZ05\DGOdW#)I&D5W.a.d-?/0LXgg<98
?/DgQgRa4,IJQ5V<<3;EB0,JdOQB,^dLI<R&TOW@#,Zd0-S+L8.4EOU\EA41Lc4E
afUP_^ba<2?GbOY(4\J=_:=.\&dZ;[^6O8:#5be_F5;C8-HKOS45]X7Bb;)/JDeG
42NO3MDUMXB;LK/FT]>:0_IGSM]_?=c_E>NP<SEa05_O\=HO^<G:\N&THCR9ZR&-
79IH(BO0+>cD0Re\5Z4=Y]UHcCdH?3&838E:aT4U^<W0N2Q9\OcQ[JJ^;#U_bMNN
6^65@@7N<QEH+WgYCF&8gH1DA6L@K^BF.<5D1=a;0\4D-PRbdT]8+3J4F^V9dZSH
A>\>[#f]A0=SM:9b3g+Y1+^5>W.C__g]SLT79ZQ>\Hc#H&;J\^eQINX(AH?Jecb-
S\NS;7?2KF^3g@/b5=e(I[.BbYfT+VA75W311AM[/.O=P^+\5&C/V9.c_M2\9+X/
)[@33?67e-WA;b1@2D:&0T9Y.Q-K(F7H_Qb,KQ-\V9GZ@IQcRaNE(c<eCJcHM[T;
^Y:gG,gB./#]]GIRb/SC&(Y6LI=-7_ZKcH+?[Ae16[M8_Q?B;3;]G80GI\9c[cLF
3-g?&A8R8;f_.7?]_dVEc=bQ<]C4<Y3BB0WH[VI,;N\;V-#E9N3F_GA[._UC[T^S
<7:?f_)D9?,:L.<;\A2N.OCHMWLMB^D+bAAC=WZI]@6GKLbP\\c_X225=F=I5?)@
[L23P=c/,KXF8D92e?E]AY[JYM[C:T\5RCJLe4Tf)]6&XIBB8?&a/c[De>\C44=(
>fe=ASJ./KV#[6)>)X\I;-6[023NR6_GDG.Q5/,+BP:3IQ#9^=LZ@I(+FbS>L\I+
A,NV\Y#DMcG2=--A-gPGR,Y(;YW0X(]\>ZP\QV+aQFW0U]@7EV.2AUa.<^.VNC(0
R1@aX>1L-[OIg-8C>AgQgJ#\+d0_bAY],+:GGeA<Y8:C^@dIT<6YZSOT9:N;aVL=
QI7F#D?(@CgVDUJ00PSJ\6)Ie]dd1dNY\=6dZL0/T62@LgdWK>UNJU;8Z^>dEZ:O
G;W&K,>_;fX6#Ff3W(E>d8F:I9.fDEA41X;Q90^8JR\,#+\MWe7-7_J/9IQ6KUO\
=;D<HKKWN3:+<F67FN,OO[8B+_8SFE]EB^9e@KNX.@;cD,G9dJbX6ca.Gf,GWUHH
Cdf5+-E1RQE:80UcGEJ-OA1JYVW0_5<W::V2P_GNc/2^HWZdZ#>F7XeBI8)2d,UA
PU@TXM(8O?,W&.fQ^1[HUZG>88;GC)(bBQgMC,UMeQX]].RJ8>@>_O271+SR^NE-
BS&g1edR/VaR#S^24NVee)P,<&HCcDDD347?\J1MDf5c@+QbP.4cBA;)=-^KG(+#
Q-L+?FVJ;3ZP=91<Pg@?/9>?aI,3C@>/dYgfR[IC1@=LFeKfH_B,9W7d=B+RXR7f
+^gOF5GZd\U(+>/[M1gN_dG^F/fVb@G5]a3U^=,3^gRCa[5,Z-FJ8EO7:&M-W(IL
F_?A/HTf.X3>#[P9,OV66,CCQXK;=URNK-O&X?EgP^P=S^4LG^X@DPM&,Md?&:;=
:TA:0[XYA[W;E907=7E_T/?4EOd5IgHZ50J?bB3=(8H]?5K4WeNIYY(X-:_aS/05
8UYS4f9-R]:XH)Sf)cEK;J,F5YGc[S.0(T[N7^Q^X5-6V+#;P:/Zg)d#,PNZDJa3
(0R[JWD.8I,PVd;A3U0a.@Y?<I9V/ad+b>,CB,)Pgb/GCD=K6\L<Z=Bg+EBb:K1@
YJe5OH2N[?IB8>Y(#+._0f=KaU40N@=87U.L)f5]f#Z,)4K+C]I[G@\>YaK)#0aE
e7A6<?KJ0=Sb85NX\G(E&83)T)L)VHIRXC5@SfM=_03A(cbJ@:U6RV<fZ0GA-^<^
L]G#A;#50AW-IAedQ_cBLL;gZYM1/P(0]PW=&L1A/,L532>DX3Y24La;_&Zf8Q/(
2^4(V9CgdDg&bU)GZ?YdPW4B8N&NY[/Se7:ALg]7U/7M/)<_F1Pf,e2O+H=S3]&1
LXUGV0=bbT>/1GQ9)31VJMJCR[Dca;M:UgMQ3Z(SdQXU[QD(1O#7aSWU2&Q.VE2<
d8=YXdWGWbTEdH]f3\G^3X:L<bGT>Q;0f]3#COLXe?#?9Y\]c0-0N4QY,.:2N<]I
\Se:;Nf9N:QG=P0-e66#]5P5K0@;Q&+SYNISW9aB=WNKfXP)?0+D;)e04?M&/])M
0fOA/#+.gE/CgZ#_XcMLH&TYIgbT,PDg=J[OSb;63T8N7J7HRX5KRR8^0(<+9,Jc
bT[9IDDXR2<c22R#Of#HDC+0DJ052POPJdKW#bORAD^;OF540Y&MJMKab\A6JN?S
5W_UG6JMdJVTY3_1E,WEL#[Z9f7VA-WP?/eRAGG;dB[8JGTW.)6)JZ>PH_UI:fdI
:M=?T][3:HXA:3U8X+gQ_FJ0:-cf]1C>^SODXV#Q]FgF54P>\MNCe)PF4<?6;=>f
4GKP?<c,aP/bbaE09,O5bD-B=:8+a1G?M5Ea,eBDb0K;L6WeYf#LAF:a2A.9a\@^
SRB7^>9;X5eZ[)F7&Ce>gJc#BY)@@_8,MgZ/[23YLVVYSg5Z</AMGDUD,GgSFA28
5dS2)-cd=43S[4)/2V2+>2ad\Z1S9]VT,\3/8[-2/\TfK0<UODTOFKdBXB\L+QYd
,3C/c^\XcLIN;b=M.(_]40[.:@aP_RC_C_.f7WXV0_5SEKBGC4)7ZH?a8e]3B2JK
O=PGGQQB8DZfX?3XNARV\JJMef0f6QHbIg(Y3?#)eQ(f+4B_YgbFWHd>K\@d/H1P
2/F@)<MUFN/]NGRRBT7:a^g+FVT]S?&b;/QOZHN5fc(;_LC-7eNc5=_-g@4HEM-#
0^J\dVNX^d.?-_6L&72;G^C09H6X[5O2?aOD]U/4=P3I.3J@B-WQH-IZ>JTb#+Ra
GXHPZ,JMFCEWaT3PG/JbPD/aJ93fFFFS9IFH-.(WaP(L-gT6J2gW7-:gKYV>MDUc
0,)2-OSb#e<^5&bbF&H_^eS5N4T\?W-JFOAUVWcGBf]Ad,fNgU(C>[bC+?aRQV]0
.1YU0U0,P;Y8<+bd.SV4X#Z/BBR7/9<\eU;AFd69_Q_b(/:2A^gSgB6^N6A3WO^P
eAZTKS;G7]4.E)>,=QPa#@=E=^-]Q_#?X@U_W@ZgJ:OYbf7gO&U&<.<Z+GgS2>-#
a[H6U&TI#VKHc_?KbLZce5/7(&AV>4=-Y0TXQG@aa&>#R&bKG(cB#(bAE]I<_:5S
>Z/E@WI[A&Y35GgUNe-QW=K(Ea71a^bXH1OI8ZY7+G#.(db]bCZJ1EeG/M_f+#MK
cJ[e^g;VaW>2Q[[P:\g2V4R6Q3@\1e->bfE<L<GC:a?+1X3\<FA@I3G^BB]W92]a
E+D:=6W^GY6)V)WFAGVM.2L+7^J>7UUVeXK)gg-P&/FS&aB(=0Xf/_:7LEJI[CC6
MP-Y]d51XU@HD][=6OB2;S:]#?9=F;RD3)P_I9L&3bB0R+fRT.J.GC:Dd]W(]+;V
1=gYVUL>c:O_(H:&?N\Q)_1[B:9M(D<[][/A>4-8N:+C^38^]^9</G)g1.A\G@RL
[:A#;12\.SJ@NIA3DTJ_.2\GN>#N,O#Z9G=02a+E[8P>KDD0:aRP==DVE_1UX,?=
12e08/A>N8URVF3.BTB.<V0MISFfEE1::KO/S(U,CbP?HMW2G5W-+5X4(K),,&AP
6RL12e(=P9Y3M&4f3NE^=Yd]I[4F.\=>3?-^CJc7>;E,ec#aF^5H49Sf/@>-GEE1
.#ef.gO5(XPE.CEKF67+;6N7]3Jd4B7Qe5a)N(J2<7_Gc(]f<DJYGY?<_\1Y/KE6
V+=e_YCV6QR(g0I3^4_>516XJ[geO20C;,.57]\)/HV(\MVD3_FOgfS/P]?T7V(3
STB(6@ZC_5+:6f:B-&C]RHW526@&B/9=8_.R3Z1cCM30G^fad>+a=dgQc8R\c_DP
+V?BQ\U6.Gb_4TKURRA=<6R?A2NN@bafTe4&dKOV+8WZMEV3,b]8gTGbfW2N)dHT
(&9Gg#ED-.F=/GVVOZQAW0>WY..SUaU(4^Q(f.\-b90>YI.;.@Z\7gdK;aAE+e<A
OR[Wd/J:YecBWTfA&F0&:^;(J^eJKRH_EPRS(C6XBTDb8ef:ADOW^BW4fPZ_@H5/
NK-+<O<J3FL\]0Y8Q5g\R1V/GDD^QAOV4c9I<4R@:JV&;R.-#;]()Zf8gF;bX?IV
gC#;6WcS<2\Mb5b_N>>=F4<+]::W:9Ve&fTJ<1?gUa^>]7X2&S.Z>>S2;RY46UY7
QD/7Wg45CPf4LbHG@A59YdQ1UGSY#&[,LN?@O&YB;H70eV@VE=-#KRQOgbEG0G]8
.U(QAU^;D.+^4f\aOZR31A2L+/K(Y(MUS>NX-=21-I2(a:W_^2N6J=EVBVP.QIfF
-4c/IHDfO0)5G[#01U\@^ELc.:OaI5,68VA+P&O/^-XCL2f?_XOcXV<+:@6OS8C;
[]eIMb7,YJ_G^DHa)N.1AG_X]ZXNU?BS@^J-IKfN0?_7+9EK^K=@SM(@SWdZN>9=
(:732Z1XVe[WGWb,AOPWQaf&c,2U[<\X,fFQa/=,E:XH6&4XZB(,WF;/Q5V+1=2e
bbXV)>O2>f6D]C><2KF&^ZRS3+,[EUPa7dXUMCH5_Z;gJH1[NY.K5J8;W>#(BcKA
+ADPfCGB#ZH,dYS#TZLP]NaG-4W1&:#bGG+@f?D>G2R-aVK>>44).d&\2^1fLBKV
g_U2:fM[TJYM:.L7&FU+0053A62.A1@J9Vg<Q=5\1-B#E<?VEYK\U&3:G,<E,V7E
YAZ-g<egF#9Z8;,O6g&)EM-YE6[N^=7aY:S/<._=^eR9-b40a5PH47@2cc&:Z];_
XW8-DDCS4J:7.8V3d@+&UA9dIH-(cFTV5^>VfA4\^UBB+(;LDR6-S:BBJ2CDLJH)
P]#2T=EagP9^X?3EF35/DdDaFaJEb^d,D4LD2WH=dZd.P9X_R/\IGFdAJZHeIdb(
HXVSO\-JV;e_aT-.9D.CXEPH8dD3LUCEF[VUZI/ID_6R9+?\e?QM46IO8Z<4b[1C
5&WMLL92cJ9dSSI_-U,7>1Nc<bSF-F&TL]0?ggW6DJB<eP-T^6/9Y)a:#e,Na2A<
T?]VPO[RJN1C7FK^fC9,,[e72BN2[f]<5;K=/?d?M;-d,OXT?I2BGE161X)C.]B9
VOBK#8Hg27EL_aS;MfO8>7DdW:5FKgVa/>-#:K;>a5)e@^2?,C@UX9?bb?&:@B@.
1T#6Be=+M2C;PQ6A,WT1bO(X+?ZJcOff:Id3Z^8Tg;G\V_2KKV0BM+13(,QX.a0&
>,6gA@G_N,L<M0Z\ANIO9AZN@Nf,DdC))LUJG5UeT(QA5#>DQ3b7^<UO[F(=:VM]
;aEUb[)B7gE7g]:F2_P8Lba_;3e6?)SULKe&R/]4C8M?1b<3U^?+3?>0>g42-=FQ
&<32A7ZWFbM3I,8YET0[#QObNM]([FQJ0\[5TYZ-,;H6cUM.dFF2PG.D/NV5),/#
eR<^E\USSZM+>a<>A8<JE)E?;Oc:1Y[@L&gDP&8Z?cR/2<VgSNB>VEB@>[6\^b>D
=0bX(b?P_V)2)?R]^W=EcYCB_f]NQ3Z[&AL8T^NS><]bS1_21\8@DZ>1[=DU[a+K
CA=DX8GZ]0/KgH^g)D&K671/cB/\2K<68I=?)G9gY(eRU>Q=:g#a72MR)4T)67?(
E&aC2)c+6[e+8U2:HOdVMRK:P[D,dAY(OF=^AbbdgVKdKJN><Z^#D1fgA6&E:Z=a
_Z:g)E9.af.6_+R3C&^4DJ60Ic06]4MKb(GX=XYg2Q4=G);PfbEZ[YBg3>\O0bda
gbed<9.TN5gb7I?Yd;O#9eJ5,,2cG#P4YBHfe<[aV;1ULZD_?F7DM,2RJN;6N@g4
3UQ>:e4O^027VTON/Ka7Uf>D7+T//XP[,U8UQ\6O-47CbEM_LMgfa;J:=3F?AQMV
AL@>C)X++J#fU\;f]&..TK&KG8^T88)F+fBY+C+Q/BT^dNV&XC>D0F9E?<Z5QANC
<@G0I3TMAcD3J/FEP?/T^9;[YT3?cg]dRd6eT\?9K4Mc1AQ29@HUQ#2<W<eD?K;N
O=)M<4>fd.FF(H6?,+M]aUD)AXT?ED2A^A30CNN_G+C6P;FA=^Ne6PL_<8Z+K&aE
V;\e)J&BBbcG,6E<7b+KT<^48f-\I8W)J2:e[1U2CC8A>XO_QHLdS&:ec\b\<KbE
1eWU^Cf<KE+-.c(^/Q+FP(]B>,?4255C)=DMJ6QHNc<@Z,#QH^1UK>#7<5VJ:cbL
\WA8Ne>.b^6.9?g5(1+Og[)61T?KKBPQRAG>M6^ff_<W3T;H<,773#aR@AK\>Y+d
2C^U.MdN#)/Pe1IJ(QZ:+R3QW7./f,4LF4JHcAH3\.;dK]dS(^^^+?-))gBfSJC]
&GHY.8G##?MH(P>;0#+?U5<MXN2#A]OIb7C.5MMAK<+b)f67;2V6@Y+gP<;@T(NC
<B,A(]?&F;g#.e5fGFK45K0^\aTdRcUUQf6Y8S<E.cX06,IWg40+-PgJPB@[0RT)
cbJTRYd)a#DNYS8G1/AJ+BZKU5PB.>R#Z6JT,00d?H@2F[Z?C9GL1G^E@gJE7dGQ
UR[<,9aM@_KBMec]IbSG/(LG,gJ1-@X<bMP8D(/57&eeFNW>M+#T[BccV3)^gMS(
Pa9W4H5O0LQc?R(<&J?I@3FN+7#_LC:L<TB&=eIT?L/+-=S)fGc5Y]ZfT<g217aY
@e/<<eIGL0.^eJ+&0=V<PfD+=a@NOPIM1ZQVF/T[/JY#dC+]_]L_^?Q_IJ5cSW.]
1__4Bf2eI3)N;.(=7-&=]1D0=KS0/^9cM>2+Z,5Se;5:N,OaNX_e;4YeZD@dbOM+
^#(@_]2KG4;e_9JXeVZSU-LbN)3[IEI_0)0H)a1=XcF)1fP+TCLeb)@63+;C=gC,
UN&g/@d^N^f7-fP9V9aOI0dSXE-?eQW_NcH_S?:dNR+KTS@8LK0(M1G;R\Ua.XHF
,CMVM2G6@I9&L3A_,77Y[K1.?+=\;GFSf/d+1(G9>24,FgD?3fOU+YdPXcIK))W\
3:a;)@6)0Qe>Q@_>M-QI1EN]\JE,,IXCWN(9Qd;^S#;8:<+/>3NcSB1#2)Q-IG?Z
5:#L,6b#C#WVPM[Lg^>O4/&:]5L[N3D:LdH9H;+>?M5KZHbOWa,Y5^8NT4bg;_9:
V1]YcL:W8eD#9O8,7-+Wb8a)eBa=7SeV>bKML+T4K>I<1.&VE7PE0c;c0AMT:Maa
+&M87Id:c&7#dgbY;&]O36KF6MET:36a?1A-=bWZ6G^P#_a)N:KJ/WCZ<bH/^=b5
b^40Bg^&>5XaSL\C9:eJ;@(AMG&KKHFIK1[b:<.P>:@/TL=g;8[J^-X#XPI_Z[FT
V,0XV3dM>2F9T:PGVR<;,.CHP(YIbN=IDa47M>0VHeG>6K=IUeeUNHgQ/MV01ZI;
10YDa&&KJQQX5,#X1F7He9]#g&bHcY7V0U@OL?a-(a,;265),/8f26P4@DS>=;,M
39)S]NJG)S^1KcE5<4f&\VVg<L+#3IN5B#:0?M6-U54U0:K29ACcb)eRS#MbT)FP
L4F7+,dL@cYcI6&_3A#PS[H^GG2>98EVdO7>VU5GR5AP)<MH1MZBK<PY&MY3//Qc
C=Fd^9RL7gG5C^.+MNO2@#(8999U&&83]+UMg?LSTAOY75:/EeWgL3FBY@H1MUR_
E3#BRTX)N6R)&XV>C^9)dW9F=NH_\,e-b<(11B(R@WV?7RdGa9W?GCK-=EUQ-cV;
[(:7)V4AJN8DQD6X8(3SLN_GDI91e(W+U\1K&BM36;eBZIB)U0&E/KS-fRUc3bXa
&\UT;C;;gKU;TV)X)PafEIB7DHS=TY:#:$
`endprotected
    
  
`protected
_HRME2UB493bQK:dSIA\c_W(2gd]\)<6<-QagA:M:-C^-_g#]:&c7),I=TMbfGDP
4a^OV-P#-4]:FX.g0We8<SKPV^G9:Y;g3?UaI&9H]BBfc^d(9EY=IW]]bHCZS4&=
4Y-dg7^FcXMf>c0\<[5843L79HYUQZMXT&ES>9T77RJR#RXKUV3H;c@MD>GP=\f1
](WeU#)0L?0EXW]fO[[eRF^&WO_OSWV0,OeD:g2?<.#3)\\eE\(3L8;K>fbA]5e&
6,=AO:MH-^FVJ&_<2@:=6(7\-=IP3S;ZI5WI7G[)>RJ^>/\1aE1]BAX?dS49#9Q:
eZ=1)Vb;(.Bf(@,#N>68G8(XV2<+fG7F03TdCa<6VS-]Y+.;NFVOY9dI?Yac#NH\
a->1:Z#93JJ=;>g^:O,Hd[g@--\E+#&URN2aHUV[RT-CQDYSV@N##UU2#ZZ-IH#M
g^SXU+fGN#TU0AY[V+<^XTMEUT)@@4S..K@^>N0_J>:]g_gE)SQ@dE&+JEWM&_aN
WYZWEHYI-f643b?:D8eH2dV#=M8>gCIWbM;E,),(ad&b5b&SZ0@6/3VOQ6-gV-UA
GS)/I;I/0,KHBLKDBV1HKKURgP9>PA<[CU59W]Rf]^BYc5?D</QXOX<&PEIB^]LO
22]4NW7YW7S)=,FG[7Y2_BTSBBDb;>.G+X141<1VNF@gN^=eFNVfZ1&^<E3:f@_L
)XeMc53=b,/G@1I7^ePJa[T0X8=U)@b[8C-JP>4CWWF&/9):Jb+4I63&B++&>N@J
]RW,K@D><QBX1C^b\GUCYV&+ED49;;4P-2dD()eTANf;:C:e4P\E(DYVe(TN;,2M
6EZDafHS(R9J1^ZZ/I1ZJIg7M7ME_9bTE9g^C:8>[Ebb+MTB\Y]:-KJeD)R1JC8K
g:O,D73MZ@U^/1_EU8OdA]2SbX_7J573J.>U]R\U-RNf,H\]JSX^(:O+],48O]#)
-S=NO^=JA=K&7I+/IPGK[YI>>fOBB4AD+P56<85WR6B0;=H=.+6B2b@4\_C0c0QV
[NYR\O0GNb_IB2X<_3)Rd),6&\3N4L=,WP=M/Ld(N^QJ^C28>5PgG(fZ7B-/G>S8
IPX3/N]H+9<9/4c(<<g&\B,RG5>gFC@0EF,.JT+,UN/AFQ?6^Z,@bRd>9YNMV9_-
V)PR6DVe/(?WV?Q@KT?8N&P=F\8;?#EOKI,f+aR>MGIEBBd8cJ-7e6FU2D4=]IbJ
cVW?)OZRRD.5V871gCf/cSc@Z@U:SUJ)X]cE-=Aa@^NETQBJHDMSdRg,fgGOO]AB
I^D4feX,I?fZK\Ee/LO<X=C.e3I1N0-N_c/+>ZMV[R7f?]2IfA,/A-]N?^_>(MMF
DX1]0JgPXMdWY#,Td1@(8.?4A9d]>>VQQPM]C9D9_4L.=NKJ3)7-,PbOga.Q+EO2
.H\\/NOE&a0O4We1d+GM^Ae\P8&6:e<Q=SdS/c<^UY621T7bX.f5bUEP[&e^_CNO
/ORU@A20^L>MJ:_8YR<M-a??JB)I)7=PE=?7H=[LK<RXFS8d2Of8>M8&LJ7F<aH;
L>;HQ6U+BdN9aY462HK&HNA#_W^a_C]RDB,FgMUVGPFJ?[5PMN1J5XFCN3]Y\Y_Q
?B26V,)4&BOdT<4@-FZaPD;R]6>9[(](D&O#JN85#O4bH&^<9RD=G@6,4&a>P7U@
Dd+8b62><@0gKYO@^bc??44dC_DV1.f<(Z9];IHZ,VIG&CS8JWT4RI.6RDLL#.PC
eST<M])D9+/8=2cf6;&OFgSa^/QcVP2);V^@FF_1fE6NUVJ-5X+^:d#b[E=KE06-
I5=0.:We/JJX2c^9]X)]APU5X&>?2G.8\cP4bAc+E4FF?#A4_KGWa1f@>&DaYD8Z
/?:7-:7KVV\8:+#_+O.=G?fHfE^bR><J@$
`endprotected

//vcs_lic_vip_protect
  `protected
VYU>Qag>2/MH5D#[+&fC9:3=M#&^J0ZbBQEG=JecU2b6L#]SPVYD,(X0-_Y.O:&8
GO3.AcSN:21<SWQ(WX0fX/JQG1ORVbGYSV1P(f2N]92E03N&CHWI.\U<IE\/2)O7
>0KTHL?4?S^,0bdHIa-COSH>>_HaHDP6I@CQR__.MIXK:L)0W?X_QI9K8+d&g\U9
#cFJQ/c4>JS/<JG),VHS_VMQUd7e<cJQG9AOaF]g_=K=:\&f<QN39EJd(X3gEW:#
\>DP))H48XN<D1@W/Z9Y#3(5M_C=(#>9OG9\Sf^UU9[_IS6UPQF^?+T@eeM[V=&P
4RMFL)d3TT]&c&D(g^g/f.T-/GBHKM)7d--@U2IU/#POf>E]9V[UX<1/#E0G?]c<
S5d4=O@:0AU-=EJUbAG=20Ub]&TG1>;Ff3XPK,(ZY]C4U0)P+d(-.S=6H35BV\<0
)/[RYccf-N[#Q-E1G@JfX\ea.@=9)g^F?;0@V)/HM.6@_A2B/CCB^.(X8[aH9GO?
-g3bEH(cG_L&C1Z9;ZP3LbUL->D7>;^KdYZ-=KN)(&9aRDAKO=A.GQ)c]H>g3I07
?S240\^.e24Lb(?12f/0(@Vb13eX^cSbNN_ODd]8BD^)V8_3M>gaYfUH<5UYJ3ER
?TE-eJQgBOD]#Bg[,B_??Y39^-a77(N75IHLVB^(2^+ce?bD9#:M-Z2Q[?K<6@^6
=.((P:#_/Q)[Be4#JgU=#V>KO](a^JN<H[Ma.YFRAEf80dKB<GbB;GI]Of=F1+Ue
_aXf:e,^:K^^33,GD<2=7_2dZM2fgW6==C8#1X<Ha]L@J/GAWJT:P0^If=aOD]XX
_OL(DGC=a#/BV:<165)cd#>;>XXC\M:2?dce1GG[]J2>M=Mb3&5Tc[\?Y-,<Q^>&
NNB\gbaAcG]CVFD6PdV,c6e?X/(+Zg6JGNOGWJ.\UX,F6H)FZ;VD(B>,/GdbK=&;
&&X/b;;/:Y-b\d.K75(C+AS+;VBJE8(KT(H4]FX.LJ;fAF8<PB0>7I6.KS]2>G;A
.C_OIQ#>B=W0&#,JG\gcTAO?/ORUc:,CZZD@KA=OZa<,YDDGFP]X=TF24#g4(?<Z
3<4W]LLQc>d&2U;1Dd03RB5RWB7b()R4:RVf?.0R^-&MO4QXg:.CF79fFKIf>,U3
0UWV;4)=ZNNV9\:#^6a9RW2^0AY2OU6B[d-L06ZVPD4_S2D9)=&XSY]879LfeZ-I
C&eSWBX=0X+]e?WVPaaHGIX&GcB&25VND]0:eF.gENQE-:\AcL1eG>bLJ9[6ZPDX
TZXa@-=J@_+X:-LJe&D6f7(U(MDU,WUG_3<K+1DU_(Qe9YK&)fY38M[7(Id[GW\I
.422HLM_4Ibg28e9;,UBQ&@?)J6WcB#N5;.6+?22<>1Z9)Qc@(1[E(gd#RY>0A8X
/fONOOI+K8EgWRMa[=MIOA)6<<83B>_]FIa2D=@Z>==&KO/EDP3G)XD#DQJUDC^+
e09910dRJFN=]+?6L&UBP=0Ie=gW/.,LNf_Tb?_A3Z238+)I]F7D)>7Z1<_>FdBM
I38)ZA1WFKLCbBDB_XbLCO^X+7@bPBceY=/4<9>C9O(LDS<agR<A[[H:J8LP.I8)
b;B).)P1e5;4RaIL)a\F>8R_C_5MX-CXH):B,^)^DFO,5EBF(dL[6(I^ec0G.CE1
?-6?:e-g<UHTJJdcD&d3=[8F4QXg9+Ea+<.f#CIC3,JcVK2+YaZfF^+,&UH1V>3+
=OOff=K)AaLE3854e379^JL<WOU6AH;d)NX^O[H+\&]L+)^4aGJ91_KCC)e6f=@>
#]:=XF(/+e&BT(Ve6\dc=dP4,^#-5@<)bbE&#;f,].00Ld>?@2XHeNQ72]&cY4-C
cV_a9KF\Ue)1?],dg3U-RCYX=JZC]7&9\O_2W9N7<:#T\4ZN#6-L1O7<JZ7f5Sa[
IJ@Z4Z-_,-#B7F?YE^4=-HWUMgV:_PJNFdXLfLWBQB+0;)Y_00@R7WgbUO7>d1eW
8R5XQc>SFAL2eTN4&4#]e#STT1^[6+E];#8-G1)-B(694Y=T?)WeR3REe&S-HcQP
>.1DFeOITKd<^Ed(Q/-0.BEQI)FdWCTF#[e#V,eG1GHT<gSFY+_XN8=)aN=QW)>a
0UV9#^S7<9Ha8CI7a[2C/0(g_</.4IQc,7X+&MQf#.Vd9P.H949:@&3?HLYIAA[f
5<f08>KW,FKLT]Z8LVf+=]>+4YfV.6+]1.eJD3GZ[Vf2MddG9@HJ5c;\)U_]O_5C
DS)FC/JaT6U-;DX@(d6Ve>A+A\)WXJZBRS[7J3ZBHSKFXa-33TdPa73U&N@GVZZC
<9=EMW4b^/32XcRa3N-e^8e1P=6NSS>Vb74Jg-[_^B((SbJP1N/cWc2F9<=NEJ(4
Q&=BaUd_QK/UL,M9;;dc<.\?[F=EFP>-__dC2DUf5<;D[//>FI(NNZ6@RSfVf@,7
Kde-9dSc&\L<(g(A2FSF+#\+g^<b_@_He^VQ;a,F_L]a095(GHd2?LPL5NKATG(6
Z6U8\Y(4N@7W5&FeI00+b>R9VB8:+e&FaU.3L@JdS.CPW-XC_+6(E^EU:ePb,]U^
UXOBDDG7KSN?X>3[;W#50eBBbIMQMHQ);Z]IK>2-D>a@\&5UQe[AONB2@+3I3/10
S:B7\V]A6@.1X8Tf3R2@R,>@A>5;V8(O4DCF-cWf+9[/;.<-I87f+X.N#9cfea6N
)\9P7G@7H;b2)0-QGc:[<>99DCNdbY8#_MPH)K#0F97gW6N&g=;U[ESU.9Je,S1\
3<BgWU?\HEbK/K/VKY_,b89FHZbVb1#Ag7c0EXf;FX&I=8/g-)gJ8#_M44KSYe[=
+,A+47+eM3g^g&Qd();a;eFDOaa?3/0a4V(_#>aTI=6LYJdA.8EF@fFWA,VcXL7R
M-].A@+NC/&#b>g-bL#P52d)LMNgP\Jg&YU#>/cD>\4:[d)^EZ0IQY0;/NacISC5
;Wa-G_PORcOQ70))4:.;_1\RYeEg6<-U,19SPPI50;6\(^c=J&W0d(?7Hg4D;8B&
Lb<IL/UU&7>_Y4&04[]b#O,-b;ZadBEX/0RZRJ)RV/&R6_48\Z9+EXNS7?gFa<3G
ZM/,4L=JK<]):e?PVIZH714)]M^1BSBY-7-b<65[XV=Q3593cc5=386)6U715XH(
C)&YUE0UW:\-DH:)Ab=0Z?W@CS0Q@?C^?:f_DO126GGHQ-Z1_QKb5c?&OM]S=P,0
&0FL<=.d<Y6^=?<T\^C_C^6.8g&W+-CFg62KU5DS#PW\Z;0Zc2Y]?@+DU/aJ.C2&
K3Z?2V)OPBd#6KT@W6;056?),W6,?D6EZ#H+PSSX6QBHa?]L<@,/+WG(NQaLX=Y5
YN)?WI0HO;,gcHa7g468,>+-A]_E,:MN8aN+W.HB00@]1)5]eKe8_;7SF^T@_C.b
I_93-I@S^\+aM,9g6G8G(N#]RJg#KKN(/Q1;f.a6K7HXegf^W=ScG;JOcMJOK+R6
1]Z?J?2-b28[>SKVdMU>94EN;AUg)#0_.>?K@J+eV@e&,^f73d;AJG8),e=W<,N)
K:MS8+3A5C>Le6eP=&P7?7Fg5XTORL=4WSBH;.O?EY8FTUPZFH&X_:IN9/Jf]BaM
/cV>QQ-6S0,FJRIVMC8d\<R8+-TH-X-/6B5Pgc/TP&?OePf9RCI;>OG-g,SPA,F7
Q2M9TC?;8fQ;HA<D=Z1F.Z6O1E(VDGI\MOH+?H.=3_>&67@6A@fB-eA8Zff7Da,=
1DAQH&BEOLcEU4WFO().L4@V=RT,3Td+L-M9Y=,:EW+63)Z+J:cRDC,dbXQ_R7RZ
&4)+1CXZLJ:&J7@1@_Dbf-XH9U(/?17M?dBH&MR.8#\+L]_U^fFJ66B,8)#cZC5K
eggDaJ?_6K;beg#DT,X\#,cZ3XSLYB@>#Be6KZ-8Q#4BEFE-)/.agN,_W3POD4bf
FdCJGGD/.;Y@+H8>IY&]UR<aDU__UGSY78KK(6F\0]-N:#U)4\DaD.gHf+._d8+3
>fS^YdN3bHGMEV_Y;d]/+W&-cM+:E<VG_.6dKX</72aGOXODRR,D&=<_1=0/@gT?
7MRB2KMN9#1c:(A=[D+1U69J>/C;1Z8S)g2CO#.5T7#=1gIWYMa,=;9[PCIC)02W
d;#+S(C)YHEXH,\Va(HM6)Sb.__U7A\M3LP))FNUG>SB:9(]&5KTOPT2(dI<JUZ,
,FW09MZ0X8PfXW_a=ZA1Y7a>HaO/MM(^9e2CdM/[f:1:KMBYCb8eE@YWE>8,E=53
]0ID^Z<FC<NS@^#C6IU;(d4-b:I8&AMJ_BWHPVRg42(BUF&<_Tc,,CFg@U=.;))=
bFI:_0O&N.&/<[3P4/G8H(4-4$
`endprotected

`protected
H#&P2C+K5NGHO]4EUW=b?,+R4\OgB,TWF4KH59\I\H5YBT0)Z/&K0)+9aYYMdR]O
Ja]BI\L_fF0IV:a3()?/T>;-NH<Kg=M<;$
`endprotected
        
//vcs_lic_vip_protect
  `protected
8:K1(]C#02:E^I09;+QSRECK]a8YMfL[f6=LRZgAfA[@FIQD5A]Y.(3VC55?1aRZ
(]^[Ng[O\0BOb0#0bT3-ZBN4(_7:-TT[&=Q_=D)?S8F472R<N_.aFVU6>V=^SBAa
4)f(0/S]97BF&bMMV8fZD0.LGQc3^R@3=+19_WK567DP_Ea_F9>E@\)VHY>GWCN?
WV)ITe]2DJ)Zb7(eR&0Ag&N5(E4Z=?c>XD0+f4XYCAYH?U:T^CgRK&Sga\HCW?.F
Pg+3-B)G++#25bJ0&8UfB+X]Z5[M\6GD406,)PK(@WM;YB0N)2)G;5H5IK6:<I>0
d5R]1)3e+4?>)<NG.FbDMIeH0/TgRP+HI#D2>.=SK=@04CeRX@Y-C?2QLf@4^VXB
<MHg<cQ:__&]Eg-bGIVQH9MA>6Z38JW1Z2Nd]8)>M?;JFPIH72:4IbT6C&I?MMH0
<1G+4Vc.51dE9g5J3@M4B-Hd=+&W=aFf;CS-M<P#X@2aD)T,)9R9R-F6Jf8AXHe.
5>-IgI#V+=TLd53,:L0&+WbVAbNCF+A7X]Y@IfbPa2R#Z>c38:O^/X]B-&eCDE:;
56I[J0E5#/Wb4YO3,@:dRYN5d[==6;<X68@#fdC<d6a4I2G>_V=FKdD65EY0BT>.
)X:7,,7]2[SdN,M>XefS;5Q##ZcKP8cWW5./XfOK;;bT[Z):X.b4ATY?5D/5\FYE
eMVf\B<G<^QD+>EM5,_>9RbM?^743)5bSH,48J0[@c/BMdTOELM9=JCA<cF&#(@0
6].275T<,,B6b)M-L>A?E3WHKZU3?K-C^[b3-R):2.4ESf:.;@MCW=C>B2)2N=5d
A<8.#HbFLd<=HKF2<:1R_fb,70L.WYIQG7^T=K\FcL@/9EeKJ7-.G8Wf1\Q5[Ldf
;KM@eI0_.6?[51&[IFffe/Z#\bZGF#I)>#A)XgePMU&eTQa2>3J;2gagWDJCYT5=
dYKB2:aJf/OE2-U2\6PV=BJ[]>).0PHN:A..3(g-.2TT6V3c5CLUXU3@>X^/?83>
OdU@+859/G?JgFR^6DIE5=J8,H#<;V#:U&ge+.@Ua+eKbE1:8MMfK+7@IJ[1Z3KD
>Jf^_,gP+VQ#U:,:UTI;JR_PN)DCW]XD90JP,^ad>/:8I?77PV?BBCRJK\;LeJXV
(>SW.;P3Y/e:9C^e+7M+aLf@OA^28.0#.\Rbe.)d3ZPFI4\bX.^SV<JHE?PGHDH7
X78e_]G#JHFB[O+f4(DBB7BJENOWI2SUNP1G>W-H[(e\ABeOU-b^],bDZ:TBS6B<
I#f/+^V1,c^X/R4T&-OU]47JP;U3\G.IFT6B]=Q2@M:Q3,]76QW>-UD\<ZECO6J0
PQSfY:NK-.?N(LT;N,B?Z>5b:EA:,25[@T^CJ>Q0S<,IPYO]FX1;>B+,7EgMY^0L
/_.e2c7=4Sf:Y;VGaCe)#^U?\DfJ(d=#G5[.VeLeK-K&2dPLSNdWCO7NY_gO6\W&
&f4(B_:4.920YVaIL?/XB+dV#UK?><4XK]T73,ILdAC-#X&7b2R2EYe^EQ[,@Q[[
C(d6M3\U5e>611P\KT?(UOX65b.6A75ZA^IN>R+d9E-=g_GGX)b09TWDF5eF&MZA
V@PIVU(/J#bTCId@#>dGORR+PMdHe]UNB)IVf0J_0Xe0,O-WI&/FFIH-;I?PZA,0
2^-WF8M>6@E?,gSD.@4VZ+gC28DJV#DJI)fDPT8GY6Ka5^5dY>?=WA)SSJ_aa,<D
BT4ZXC3WgD.cRTW,#OXWa\IH^K&]OZ,Ica_ISN#S,GS@=&S/NT9SA_+B/0Y&b_46
Lf\U3^2c#@SIJ501;Qca_YOJ])SbL-<eH3&,>gPP?375UaF.d@^-6VTg&_YL6VA=
SNB>&E#W469Le&2;?f#P=B5G?QfE1G.Q>5d8/?3T5+_L0SDM.5F06:??_1FPJ9<g
]/TPTWYSb))(;&d5DYaJY.ZF=7RO>NIR:XJ]>=UQTcDbOgHcT8:ZR1<P>4EQEb1E
BK;FZG@bGB)b[f_V38XAgPTXCP:\4N:(;T)f#GWOP@&Ja=Z6;3Vc(fN_)N-Q104V
7Y-b7;..74=fB:54&WTDB)OOKK.c7#Oe19&+[O=,(cS742+GUebcDb:(O7AVNQGE
7;#GTb\&dG@0[9AE&gP5.ETI(@QHH<I0(]04TfGDV[QXdUQ>).4,XGDbdFg#4F[Z
.#J;II+5DXM07Db0RS1@_-5F6,#XXE?[9.W@R_CU<ag)E@e]4D2LQ<cOES[I@@/4
+Y(HDX4#fWdIWS1VH10=e)PG(?:Z[XF7=\.0f7G;L3QQ]6]6^g>1fU;>^J-SPTa5
/9ZVS(df^c0#J&d\2K/_Ye)E)B#[([L<)>fBg6WdP@7HYL3B6FMQKZ&a:)2GE)&4
@gJLMce&NG)3A2DL&4S&B)H+N_GIY@L5a12_DAH2X-R.:^8:gDOYQIP4_&58R[9b
>_V_LEb0[f[Yca8:W^_VJ+KD?bI/1dHgQ#a#)/PISDHbgBW#0;X??5.0M2EE;,IM
1&2Z:,a/,XaZ9G<>SHCF/_JM[G)N862cF&a&GHBfU\C0;3YXN7f<CGTR0-)OUGBT
:1>69_Y?\H6Jd+cLd.+6HG\41M1O(,PQSNB;g7(&.747)gaPUJ6FYKW_9PU9Pe<W
E_ed:V&-V<b0)R,]\O]K,Q<T?6YQ_R8XcP4C/F/f+,Y7S.V#Z0Y17_PEcG7U(-YM
OPLB#I(F?cRKFN?&@Z10H(VCOB+N=f4PPJP.Q/OZO.>A=HPVOg2=\W_.[[\;@1=E
9CG42./:9X4XK@4<YeJ]JWDHG^Z,B:c16C(\DW[](/XL-d_STWN4G<VN.J_BY+:2
d3J45CbM4SNJ/<;ZbBE0DRQMQa?Y].HRW]dbgc8c)GGSG-^-@J4>@6S=G5W/YA-Y
+LER.1a1IDO);JE?X2NLQUBLW+>I&R2:AYFAd+P^TeY+,=D5N+_S07&(V3C2BL#&
[(98H8B@T2A+FD9BfeCVYT<;(79dJT5^4D<Q:E5?,Oe<\^GST5F;^Cc7I1g[;B&<
d9_g\:Z>;AT,^:b;C=#a:CHO];:#GD1E@8M5+9e@Nd(S>UW(gI<1TADRFWA._X,^
D1B62\3eVeD,KJ/<.D>:VQIHHX7320ge6:,6>,(gD3a,P<87\SOLCE7YZZ:D]W)a
BPEB1@PB9W<6_DdX(LTBBEegT9PUPCf_gM^b4_KB:L/#1X)e\YYQae5/_#KdNc6A
SLGT=<8/R?^AJ5,.3#H^IXA6]]IJ=Z\:2_]@AcZM/OX(Wc9R[P#f.;[Gg68KN=57
1;28?/I\R]<SA7R6=BM)I)+2TV01B/5PXDa@V)P^([)70d;2+E60)_6d&MG]XWX0
JGfYS3F6a1UZN,W0,[AHg=P1YH>EM7=f+-O7@cJ1K]W1(1\1&[C@:1B8N:Xa:_6P
]D/(>JRV&QQA3C3MS0[eW6\Y>#_,;LCa&G=O9)U=b0EZ\Ef&51PR9A/D69:8cX1O
05]fb^H,)5LIPQEF1UcP=-UP81NDc;^P>N;0Q>bXI=gcaNXBHM:e15F5NM^-L1X;
fGK(M4TS@W8GS&1PS9+Q^K2&2g>Z5T\+d+.>aQf/S79.AQb^GFE_OJI9\cL<=c+3
TAUHOTIP0L]d-T9AfAX(0QM/Q6A(L,\FaMU(J0)NW5Ld\d48G,a->e>T_:A7V=V3
4HIYd#RBcAfa5W&Z-0Y1AC_?LfBWA210@g7g@G_CSb&<;HI).93>F@27Mgd(I9CK
,RgcHY)DLVG2MP,TLR:>GIf4T1S/;^KZG)CPXC^b=)SHVePG_Rd)B6ONUAfd85(E
YD1[8EX1gR.X.8dfEG[S@QI-SRXDLaKNg]Z9e1<YX(96?I&&a@,YY</=1P&T8c<S
@AGG.EGPA&N>g5N3C5EYB5O5f?V^0LTBR#8S2_:\NBD>9C2E[L@&;U9fe]:V2ce^
18OUK/LZMIVC<45?bKa[\Y:/\=-L9J4eP3I@2f2_-EY08]_^-:Wa::VNb8)]a@;[
RJ5@AC&+JDBM8d<1],HeA?MM#E-2/8)F1Z0@#ZT[NW2/)e]#&/PNG[E^Z>F)g/S&
C@e2MBSQ)K/MK@0g82?+SU(c-U[8C=f8??0@?9=K\7<BH&U67VIN===.,#C09[1(
Xga;F^]V0/S\d#1#\cTW[47UM-NO@/LRXQUB[SK]NWW6CNQZ2I67cK+I>MSR##NY
RYa.Oa2CPYc&a,ZWP5Vc1a0dOTZ:[N#aKe5Kf8]a,FI.X/(F8#Of1N^B0[Sg4f/?
3)aGHSDGG3L?G@c9[;UAC\/M(7F+^(^D>4,)>].-BJZ@dGeO3P[f:6MZ5?]DF+a7
O&&S^Z^H8)WT8]OR8gDI4>Pc4<D[T-U0L4^d]>I9Ha&7f:,]IR:Z[.?HJ=N\<J0/
\CE=?BM<Z=AE&Md2E\RW<2GJcc/D.YLQ(NXL7;#4+#DN]N.C7\:-1>KDMZdD2]Ab
._D(gb;.?Q?_RE8]J8?96;4RMP<#ee:ZAfc3SLLTE]W>aOg.g,ZN)c6VP,2F4:35
R=.L,cM@BJ/.7C=[PafA>0#CBM0[[Xc3TgX6G9JQ&HBUV<N;9=:1(__S:bB(gS0+
[CB9@gA1/bDC_M,.Q]W3FRgG/_@R_f[P:.DSP83=O;aY4NHgfeXN/GUP[c2C(;5X
Z-@0F(E=b+)22S_C;1>-G0Be>9CN5R#H7[U0S2@B\=_DHP8=bQUV(VYA\H-#de-,
LJ7@TF&0?b)F[^d0A=3D,U1=1IPB232?DF_#W45XYc5N.gD=](__UZ<LdH0\J,[f
8O[).SZTf3O/K<F>)06M]QKH5WFgD938X;1YQ(Ja#g<,)@SgA+.#1e.XJ@,N4Y_:
P2Bb[,(PJJ?9EHYdFY2K2DHccPa.JB1Z_EIDD=Q5.I[,-gV7#/OY;eT&aEW6&b;J
(A>//53?PFQC+UIYO\;^E9S:C>;[[3RcfOI0D2cD=[(f=?;fWOS=9b.a\+,aDE9-
DX:7P;7NYSHLMD5I62,ca7<[:E#\RU6+FEQE8#YG2Q<H\8B_[[?[eB3^@J_B5V?1
0GNb_&5H@K0+^.X_42a6\?1CJ65OEYcYE^H-4(RDAgJR]F22>:b]fD4U42EdCFfX
GEF/W6d0J@>.62,&1Xc53)<c97M^0PZ)N;P56C^_f?UDc?A<FAa]P\ZD=Z@KYe&G
YYQGX,Y+.\4#IM=.cET)5W_)+_UR2)8e6YSOT;Z,e9eK:PS)E_[.VJ^)W]9-b0\E
0)e-^1f/VNO0.;C=[NPF-R+gC/g31;B?C3H1==6)4^K@MLZd-.6T2Fa01]2fPcLb
?2HOZF[,]9P^aPSO[4:RgYbTf(>4##5g)a<e&U:b@\=A#LJ_/b4JW;6c/K+8L)/J
;O@IE&LZG4EXG0UPdT,I8EPI6&WA5=F@C9_D5RE^G0.JL#bV5a5[;08,ZbSB,P^\
3N/3JLD0&A4TMZAV>?U];46(<_?6C]8(37,JG65^/M8<>0)II^bID#8W1f33/JJS
eNJQ]8/F+1&a?M9>Z3g=(>&;+PLV^a0\/G1^#0^+T&1gXF&Jc<.HAL/WR)23d<fI
TKY9C/><H=0D2\<@JHSWSDKW&S94FK5-I4JBY2>7_M;@:+7TE@?(>1:e>BQbd_3c
fF5P8SS;>@50b#[bGf>YJ/NaO5\b.Kd1\.7+B>3__)Q@/E@K[71RAY9>787@bZ6O
NdR_OfL6gGCMCa6ZSCMdP1(&d)(I+X#>KMb-1cV_Ue90LUZfdI@+3,LAH\dMUR#D
YM=9DbW-d#^,c+<0\[e42=26,TTL-4^[;JF8\?9Xaf?/PX377Y[HOTR\3W-bX2eS
[SBWC#G/V3]E4J(&?8VIC[^fFH#_(,YI1:5>RS5EC3Z:>,Y.7)I<Dc2-^^VI0,+9
5LD2<NT^M97[>MXH_cR\@&c(d>+bTeQ)/BbU.;Y@X9,2(D)@Pb5DC^VS<7Z.ZOd3
Z:=C+Ue?XU6>GXF;#,Ke8+]N)e7O32LcDRa#W/U@ADGFDY6X]94,&>W,E\]K1B1/
B6QNG;NM3Y2&4YHYUH#<N0/=#Hge[#X25SCS/T]6GPM?Y[[]b<4YBaFDJ[[X@DcL
:,(+(KXe>>d>1agLgHOTd..8I3+DCRY@[^dQ^/14TFH4K^)f2a];8a>Y_IG1_1@?
8VMf313cJ^-bMB/T[YGddU>/69N6G<X)F9-04]R=H:@bR18A(W]:;&Vb.E5PETAU
d4HO;#b-VX=_]VPBRJ+HaYQY#&1f5QAe&UUF&&]//RJ=\cd\Z_V]YRIM1QD[^F.G
;/\daDg?T]OZY9a_#1FLI(2?X/T+)IESF0dM7LW(aG02.Qc<^2YN:eGGGfZLcg\J
#58\RO]48>b_/[9+LNJV2O&(gNd(:PV)?9ICB<e.:35LR[=?SB=^>WG[@bg[N7a:
\;>A6\5.5gJ1YM3U0Mgf]6-33g45eO;E3CRN+_4KbZUSPBbfQ0H>B7gKI8DWM8)g
FFCJaVG:H9P5/0d8Ie/XH3e[c4@9SM&0<2_+-eQ.O&UC\X?+V>QT[)=5QFT]U)dS
H=/G>;VSL8JVSb91UY8.d[6LZ3b7AK9]2TW[eR183Q&01/;97P3R:N[VI[PN_=,Z
H]21:LARWYT)HeOI=UGP8P7([N4[R<W25IX7^EF_Df@bU\T1=fQa,>\MIZ-6_=BJ
B(ad8RE5IPVT^c&F6R?&+8:^.TEZ>)LIQ02:OVN=&FEfc;;@NI0(\P26ZbEbPJ;1
UVSB&48+UKZH.=3P)6gA@aGgN.VWNce=E]W?T[YGOWAG&8D/H/.g0J=K;/-(#(AS
:a9B_&/,eH2Z5P908d9ZRI2P6(A5#GJbM0@3>WTZLR-dZJ\WK/7#QL8F&d^,bg;S
@CL<EJ7H_e<e5W=XO#e0,(]46[V[F@>1@Ca6I#XL@[\-b7dR#e(27GA#T[K=-f=K
H@We=eU?OX[7#S>Q:--5:.Q[D@??\Tc&80@VAK#A32H8#EC^A]DC=53Z@f(=+G7<
(OD;3G;be1)Ra#NK6(DeYbf8@aX>\)2F8FL@,b\E>7KCQ#+:)+&]LgB=.PC?NABV
V#EX6,T7N<XY1)P[@S2P1Z?E1SM98K<W=#d&fK&f=(-SfNZ4W]NF/:VfH.X::L)8
0>V.0IIUTc4TM>:2f3GQ.+OZ-b,)1K:SX_3T/6Yg)9:g6V5FGC7/?LAV30>[fJ8#
[HPLf2,Y43A_U0PBL=55D)619:gMY[?g&H;F16<GcKb4F:]FU2O^]aR=bZYP,OQ<
E?V?_N2V8gG)P9W.YTWJNaI2.[S9>.]R7\=X=#;N9e=LELXJ9J),S#,^&0\?,8O6
=,Q&>2D2R)d#7Pa:e]D6V9,fC?eWUAEe#[XCF6&0@\WZa.JFA[G00CA?_+_++B#,
AP:GE1BL#O985Rg3bI)=2?fS2dT]aAVCc=0QI:WWV01CgQZ-5@T)#OIHfTR44a,_
8K#8=YQCFG/4f+>8&R,d,^U<3-=GfS<VOJFY/^&#d;C[Le&FE/aEP,B7DJfRE59U
&/<D7XD6=V.FEVN:Z@TA[)fcHC#V:2_?CLVNW>afDeQB2\L=f.G2gg\+gTJ6g[9]
36DS\UB#):,K@NQfVZMH_BHTb:d#DdSf\8WX]5)M/1:W3;;6T1&-[]?B5ATTI;L1
:/?Q3,=&E7]K6UP01F?1R/K;MTfX#ZLY7PZZI(F)5e^SJg66D&.+Ff?H#>;@-?Eg
WB>,U#0,#>G,f1B6f2CRJVVa[TGaAKEOPcW&1eB>YV0QA4bLE?gcUVB#LJF@X+@[
PcAd]2/[YC_B0#-4J:PdLN:X+MZOEUS[7IX_)3C0=D(/ecD6>6]He9ED=-YJS9KY
7B/L)NbJIRG[V3;[PbVQb97d-gB\b4AJFZAde6^&bYR\HG-<=DIfZ>M);cEEI5gB
bEC,f9:_UQL2K^]47(36A2O:He8^0F,7G:)SO/gfb\P7+_MX_=cK#//\K=VL0=U=
+06=g,5L8U:G(KZ:NV)CYKMTA]c&3Ne;R2)XXa8Kc2Ed]P[41;]<a8)W&7H^O257
T4G3=_MXSab:0OHG]<AOVP2AUc/,/NZLG3.g&(::NNTU0YFWBUAUMOO^X#edD\.f
MB+QRC+6MBM.CY0,a(414/_d,I1g9]&)cU\E?,,M>^0+dA7<a,]eHe9\1,3V?cJS
XA2/(B7)D(KSK#TV,Xdc\g4XR6VP(3#2)S:5LLNK5MU9/,Fg3[eReQ+dSOdG)>F)
/=,/RX7M.1Y&:YfK=D>d3cOOaLgPN6Z.J)LD^568ddZ\5[GaFF3?.I:NP,[3W8NQ
DdGO/H]U0[]IPH.=IA1^L)fWT&;e+###eJe@GH\J)A=aZ\<H)PY6^R&5]P/>g8M-
.S[UEGR8#)a-K099J=F4a,N[SDD/V0f1UCYT#J1P.5N0GM[BEQTWbU;ZHbGJ0(,U
]N6dJ>;H#;eJR1bHHSQ+/L<@5C:>+_EQJCCgEdF=<<.GQ2J1.e.XYI7=S+(bIM7,
V1_gc#g<J3><GQ+ZV&dNP_^^S5,JFBO)3^V2g@;)a,C-()KB4:24Q-;#X8e#\S>K
2fVF=@X+SdO(&MD=BaUU??MM/&c#JB2@XN=J_P?-9Mf2/_,TPg1J8FJgg;X;O61Y
R)PASS6)MQefP5N#f=#^BSGWI\Z)<50/<VFfQ9@#K:D6H_)I^SfTN]O\_S_e[U:3
:-4(,I?XaS;G(GUed9:AI805[&PVaK9b2=T<MY0J(HU3\>.-)]NN&&.1^TL(Q[dE
T;D:DRR=[(D?+bYC0PR4[&GfXYE2XS-@?D8[WcVKE)?]IP&;@]Z;M65X8TG&LFC1
=5:I/(0@HSN);XS?7G.fZ/Jg&2&6e977IZ.[2M<M_0d_XD3Z/@KFa5bF</2F^7^+
<IW\1?XAafSO^S,E7T?7?2BaVaa@=MHY,J(R^R->#&N:@M.C/+,^\RH=M<ITNgDP
2O:5I\B;7baCXOK8S/CKfN-@S3\@DP]Ogb7Uc;QWgR;8]1CL&B(g?I8d/fabX_;7
HP77:8R3H3.>Q^(c]]JOObdF2EUHOf)d_=G:aE;a/VNLgT/,SI<#=>Y,5+Z=DHIU
(TR/5+>EW,G5(E5RJ_W9[F,,13>:69;Q:H7TW]\_N@4/b1?,VYHEPX9^&I1[NY-d
aC.RG/gegVZH)A.ZG>^/a6;K(b.S,e(TRQHQeRf\&-AY/GU](R\&:T8W#=?ZPXT=
5&KKWdC44]6C]-N=G?+<=G2#64@-9-EO@cNL=)<RE3/Vf4SM;HXC&/fJ^gV;7]Q_
F;fRP=FC9GLLLO2>+)\K6Z;eQ&b0=)eT18DEgDI50)3P?O#gDc]@2c4)B18SK7-5
74Z<?C^4]E&G8DS6#AgbTC[\T1]3--0BO\K:\L)PeXS^@MVP/?RBPJgJ4V7-T^>/
^?+FHSee^>)6)DHWc4A-;_IGI^Z^.HG;4D.-cM(T-#6FBb4D^W16ZD:F+Vcd.bFC
R@6f.]W9CgW;e,Xd]698B^^H(^DPc.669C_5FW8_GIQe131Ye6SHG99E/7ZCA@Z+
+:1B>+#^XaMe(g]@JX-P;E#6a@0?3<W^;>N+f9Y=Y5=e+_2HGOP:6+dV3<7LWgJQ
OWaUF:AU>8I;W&.7N512>PddcWaDd)8LCN^cV@V,5dE0Q#^>W1?+T[W;DYO]6;C)
4N^.?<P-C<[Q_R:)Q)JG0WF4<H,HWCSWUBYS_\/:F&^R9.5S?3RGVc[e;>b_fY7g
9^\c]d19gGbF,Tf<=YE7[442d2J0IQS./)S5(GFVH,E[YFPbB-8aL&<C+b<#I_W,
W5NbZ^RVT_aNFFE?]]b7I)Z@.LL<gJE(-3=dN5BN8g&EbTMaF0,_C,N:/[QF\ZK/
CK]gb^VCO.K+g77Z0]D,5)bO82X\9a;)I-B6e+K=STP2.IUMWOPgY@bZ(Y<\P&?U
Z;GJ]NQ?fN?>AO/ZQNE6_)Bc;beS4AaU-#TV>-KJd>H)54FU5OJR+1\PQGP6MNe?
E-MFUb+1_5EMR:YQR\.9F<dUeaKR9IN]^L0XeL]&0ECHCM<gN9OL#S^I;>?GG/0-
7UN9@)-^dP+;3\2cL5Tf.@FXR4(/^\CMIAOS;1NRN]X8N3e_A[8&M/]3\?^^d&,g
5fNA]N?GVL3gC(Nb6U^7J\<\3b=\gR,aA(::^.7YZZCfC,R#aT.],#E,\1W:G3ZQ
NLU=KAXK/2eOT/.#M,+PR^A(fC:Y:VR9]0ZI[E7=CK3ALC_;f_AXP[=S@^A5eJ=D
TKV_cUTQ(SdVU5.db[baQO=D32330Wg1a;_:?OLYP@7TW]HC&Y5=J#([f#BZMV>1
YC0AV80P1e1a[34BU-Z=TgR-()<1ET?>#-cZO/-7U<1A^^Ta9OV)72TAT&7Nb93(
P9gJf#4V2P],8;_6W4.#O4Z9cL5#:TTHS_T:U(>\R#XWPc5UZ?0WWUAWD65=:94Z
D]e;1c?Y9.?H>-9#G+)^=PTSB0e]Z=2CYE:-BIdcB/f#3I=cMO^LZ2gO1fNFd3/G
)&]O/<A>@16/(3cI1?>KSa3^?1b46C0#P).-^#;b\?Z3HAE;PEYefS\#3+00Hf1e
-;;75V5V,0#MTJ<5<_9\:GBdFF[6f5;-a&S<S;Q]X^27_6f@MEH)CfS+#]?QZ;d1
#N_f;=_P1Cb.E)8NF<BVa&4R1)7f^20TYYG/=,5d+bP3J@C\/M^K=KbAAa)J@#\7
L0@fTaK7<@D5?<_E\K&GPP>=9;XAOW98CT^9Q:1/DK))X]e\fXY=+R<5TF\A@F7V
T9?D&YY<_dbH7])gGVBdGd<@WAY,?IFSeJEXH5-\=c.6[XdHf8W.3?T>,HSPCF:N
ZU6XR;201&A>6-JAF.HZ27_XEYYJN2&P[de,bMH4-09D[C5HTdIcZI+.A3SQO5R9
X_P&<9S87d?WL[/TF9#0Tda+a.O?B[YXXT0S4/06eZ+W-<U+_.d=(HVNR182GEZ@
;@S4aae95TJg_9aU+LAZ^L6gSd9LA1=-@..GV1-_1W:5_#b:g.fGDY@Z,,,90/)?
O8<2eX9@D&E>_Gf[<D=7.)&:VdA3I_O:g[7R]FTN&RR\V[(R:1KKC098[6)IU^c=
;G>5\O+B@M\K8Efc>+_>.R+gR3g&F=B-1Z8gdSgA[Q/=9Q=OG,0()9Sef3#+U:J&
>)K4_+d#_<XHU^Uc2V18e(.D(L@2;I@[BLCQB69db8BaH5_CJQUD-9e/,b#4N<LJ
IIPbQ6U^TJX;,+6JMf\J>05LG@V1YEL\8?^[:bHe:9(4FANcUfS6-<e0G=1=F=@/
GCC=P8LUbP2]E;DgOK+E7EXS/2OG_9V+8]7b[VVY&Mb>&7J,#+-62N(S9C67^S_,
:W5=SP13K)^TRADcO4A:#4&XQcF7Y^4>YP(Q35W9W</2C6#;:&+G9c8<#95S8URS
.#a-:U,6eUDbHFLUJXbEX2eYJPL4I7DA1GAQ:8_)/.3aJ+EDDDW+99GQ9?g4,E&O
YXI5T^@Q-CbD6e0P,WZLZE-ae@:]&/KgDc1GXEc@T.[_ZcTNP(Ddb5N(VWT5gT?f
:E2gVf)6Y5WdP^Q2E_;J-IBP,V/G[P]b9>(ZOYUCg_3fDZ=XES1eLYeS[E+C)XcN
?X,_QBe,9AW\A/>ee193\V-I(GL[R;3TBKG(:8G6M6g4c:I#,Y4MH8-gA_TOg<K8
&4D4N0VV<G@D0L0)g5KH6[(D@g[6LTd#cV68U<Y8ZZVA+P5NM5ec]TU^f)ab_7aZ
IfAZMUG\PN45-FHD@ZJPFZA]\DL7Oc:1VRR:gYB0]]EG5;fV4@CGH1d36;3FaY,K
\54gAP;,9GKf3)cD1TC]d-CG&)JH3bU_:cg.Y2[bK3OX9GdX^WW=98L#,4#M:[f5
Gc1GN5R\?6eF&BcU;GII#7#G/7Y&I3<BX3HMdGd-[_a>?NM\#S1fL_E,MV/_;]ef
K(g2Y4<3O.U#PJXJaZ\^X;;_M)MFQH@EE)N0c)=<BW7cCc4=##C@AC+FCD4W1<e,
K+^XIT>>.0[dfPS<GSc@VL)gaS:@dVEZREF\Q]CA.E0WI:8[-L:3D#H\D:5ZQe_f
/7d13#FM-U=Y?9]5HFLW+_JA5F;\@F0YVXN0KbOAa>>RT?8(&06E[[N.A>PS\^:K
3R90<O1R9+\CNAcb^fd4X+(OL\J8Y]g3-HX5=>fF\Ac;+:&a<-VeLC90W;D\^H_b
[_#;2AS8.SX<>HNSY<]18c5OH@ZdFgb[ceAO#=eg-N#[Oed>0&Hb\?L)QMV<LF9B
a4WJ7B-d#4..)^2GR?fTPCEKY0)TFRa+0__6TE8Z#D?,<;D/QR+WJ.8eK8XFX4]2
QNJ(][E_5B/c1U?BD#\X#.5#+Yc6+cM8+[,K-&cd-+,,?B@2T@AZU8YSOX=7A.+J
1]SAVS7b@UZ;B?Y1>E)Z#NG<;S#8@[W+YVAO[W<A@_e1Q;FB:[LdRCQ+_KEP4G05
.43B6=YWH=9Y\XAL++4dPS2AJQ6\\./_aM@[GIPe,7O/Ob@ZM9CQY/eR@++:=I;,
A3e#1&0TV?BVFZBeP@R5-dDWaLV.XJB)\@O,c-/=1F>FSKF\b3<JK;),G-2VZ:a:
V=EKCYbIK#(KPgW:)^_9cWM&?_GWWCf06Q2-cR5(W=(WQ02A@&6GZWBOT(A&618&
SR.8dZ?Q61_GLbN401cb2<TH7;)Of:FH#)?^-4+:ZI9:9_7)U^P&C^6]f?eYV+K2
2?DP10]B6a(7:3)9J)1MFP;VB,4ZSJM,ZB1:@CM:J3/58g0I#8T1.R;K4E\LK+59
]=g5MK#8LHF?5?b.AS.#_e[?KW3eKDQQIg;J.M3+Z-d(2)BL,9W,N0bO_[g]F]UD
O[G_/gKI,-H&W-XS^=3a#.(ZG_9<KK/4A&=da_Y7[8RP_VY#.NOd6(^0>2UV1)bG
&_)R_0Eab4L/I>aG?^X.2FaCK5KP6&PLBPJ+3.G<YA/4PPE0&U+LT6=+49Ca7gO@
HL>]RE6);;9V5P3:W-0-gG8-YNd\MVdPb31KGNUZC#)E@W-]IV.+Y&OHA6e7PTH_
E?2Kb+EK3ae^Zf=E5_G&NUE7<:[G+[PERe8S]M&^>@H<cYT+-d_9AD<dg[9LQ=2W
2IB;^7E[cE=<?c5O,HMN].6&<R(f+PXf;a7dIYf>#d)__1[IC#,1-/,XD]UHC-PH
B#7UWYQ)?Se;T<UT2Q<GDNfZCVB@gIKK=O75JE0#c751YE9;],cc2&)4MfJ0U__F
&O(D1\YCb?)YW?b\J#UFd[[Cg_Qa)FSHa]_S&]K,fgcX8LJ_SWR+2g=UDR]]Oa)E
e)FT0a78f:;Gd,RgR@3/IMYUW#78L)d_MC:WGU]I+a3P[:RYW2X;X]gQ8_=WH,FK
SP0DeZ?J=S^6=@Z=[5N,T0U3KG[8KbBb8&Q]^;Z]0_JVbCP54;,1NV:(<.]I(M:8
/0<1G+,]@S+/;JP.aV_gNF]5HB;,O(Q?(#N+:fTZaE@,V&(ZOUc,5f.9ZcN2<OPL
H.#N>AGC4Kb,_DJ.F+@M=-D(@8O;GW@FS:&E:5U,M5@43;9Q<gQ=2)7S/1B0)&57
QLd>FK4&TTI2N[MYX[a@T[3SG^9,#YD5QH<2QebJMF5-#S.&5-SP]Z,fJA3>H)B7
)/ZRf_:J)HV6S&/LVJHC=&62UJ9+1ZJL_gZReT-V0\;d53C4(?;Y4?SI;-V1?P6B
3ZcIbPCQg4FRN.^STKfL=J[V?W>62gD43[W<HdY@5-]SJ96O-]eI6C(YZPQNf^L)
<P5_3RO+g6d.M5Z_?;/989GB==KEFOCY6GM[ZfY>&@UPO@=H0<Y[<(fB1AZe_XXR
DVOf&6D3E-(,-bKdKEBW[F_SRI2]VNAEVb+UQXe[)]9E/-2:S5N#)(Q_N84#Ra^,
W</&UCgAYJ=_gA;[)gP_HWV085RTWQ2Lc@fI/d=ZBA:S>WT+VEECN97>/#J5&NgI
0f&B<5YY/cLH2#U;e:@eVAZGQP=I;QX/=?-2G[L?9VfHI7U>:DUT)K?L:NMKUKBQ
T/^X&+34>ePBSI?Zb,]0+HINJTGEDBD7)5VW((dU=YC-Q[V+JA7OdHY&?/RHCGR@
167T&)_L(507TO;>K_,ZNM5LA@C>U)Y5RW3RX_R5g]PD1#2]K@_#+eZT4JTF6)X:
RYdMKKR[H/Ka.?NAJGB<Z&0HJ@B)0DD]f>C0WdGLL3Y1,1ePX@U;JB/6[.Fe+)+K
U]9B2bE-G4X>J,L?PZ.fWD42)>U>2>;HQ96PFW/.Z.YOgeQG/@R8L#e)8\TVVSa7
P@cgaEN_L74R]>@JJY->d)L;)BXN=b8A/+F-ZYcf6=@>,-)X6D#]MS&f14,Vfc:,
PE,<Y1J\ZCM-3d6B<?MKa[BQUPY8:eW+\?72cNWU#R&E/]Hg:H^,(7..IM?)gdMb
COH]3P(IN;eKGOfZd1[G8J+9gUGSZ]JEf;_b3b(GW)_^^U9a;>+@d^L6<2Db=460
N+>)PCNPY(^U(:GNRN0>X:/_,&T_<E/[ZI9-EY17U4.V=P26Pa_1XP4V?B_IX<:9
&3<\2@;X^#ES_B;MEXU)B]ZD_-d)<Q2gbX+1#HSTR3U_U:]a9ZMC7JA/,\PZ<)NM
,CI#ME9NDNfKfdAa3Kc=K2GDH)56Ma6&dg=79VD#g=N^T:T@\_3E(b#f3#^6efc3
K#:96MIW9Ff:M&\e+fdbSB=a_MScW,,.S]UH[9:4-+)S1:7SVe.[b2BA,;>PS\_e
:J+T:X1g1]4@_6\2Ha<-ZHPXDAGLP^IL;<7-REI<9([>,AYfR=<^/U-KG=Q\2:TF
Q^aPC0=T\.327B#DHHaY0:gI7YXLdP,/<SWU)LC#f_/T]b6PA9L<V&<R@GRP^bFQ
dIcafHGaDe-=+&I[fTC\-BA]7E:)B])\+aX-,cW)6&9Y#?P7fdI9=MeRC<+-M2a5
X^K6YR]LC]PUT@=+.)f5(\8<=7_DGT;5a^JXL<60Ee>YLW6e>d-^TD):IY5YEGeD
+LM7A_Fe_gC70945X#<+,T?IUO#E/:;4dfH[J<<a=@I?^]27#]=IDFB7LcJb5+BM
dO=DA(-F<NdFX9U]?@6[7;)9gSXC1BTY-#]U0WZ4;9Y=<M7/0/,R&7;?g^gNT<GT
X,NB-bW>7?E)_eJ-UH5D4]-.g2YaMRTbT/Wg^:QE\;;5GB\SLS<HdAI^[QP;MNLN
9P<<Y;ZA-:E.>;K[d&UNWbOA+\]92X^V9&>+8:XRLOV/bE9ce?W?JJQL.T4-CKe>
<1\Ha2B7J1VW5/<OV5F:JJA_GU=SQSL+?79YZU)Q5gI1FC(KE(BKY.GfC98/._NL
HCHIAaLX-8b28ge:/D0[@dN4WPYZC#.Pc(DFd3.53g)76N\TF\4]C5D@8)SgQZG4
)3CL5<eO6X^dD79H;1.IKMC060b3/O5c4MO>Y5PAE_A=1FQL<2TbFA-_-F=3dZU<
+A_d:CQACSNLQ4G&P,aY2584UCWSA)SH.9QCFNg?RH?)=1Rd)>CV:_^#IBG@ccPg
W^Ub[1/>S4..dAdL@[9Y:_]PQ=F9M4?OE=K#G8Y/CR\@GAZ_+RV8C.O1Had#^A57
.U6<Q^bWZ7ITS8M@-BMO_cVAQ&\<A(<fHKBcB(9V;9S=AC@fJ.V0ZY\Q7B&7(O)4
\VC=O/a#?_P+.B62Gf9WWL]7F\,Y_O0A_GBW8Gg^GbD-[]=T=_[<ZT8\MAHeaDVR
dcF/\\\;V[0SP&R6c^H\X,?2b;WDHLc^N<^@N6S20&579C6<]C#aY&YNK9#NG85G
+6WH6ENT-=HEUWP-HWBe<GOFA2\J3Nf3H(e>OU#A=DLYH(T4#&K+K.OfS^>;R7-C
eK64>@K(Ua[WU^DbZ(X]7H<W[28[FY7/NE/BG2)RB\&bG4]Ne0__39TUEN;L>NJW
#cOE+K?.=HMB.IPKfU>)JJ-NL]gQ(Dg-N?_Oa[^LdeNSFB;=AFS>L0J@:58Rb(Ze
g))S@,RJfJ.(Z>B:A2Nc.C((@;f?Ha-a48#(+?.Y#;+PdFD-Jb/I7g83,W<F=JcA
/2fXF[gY;A--\L-Z.[fCe@MId,5ef0LcOCT_e;SP;QXddPY70T&M5>9(55/PDIaJ
ZZN52O:E;1(E9AJZH+VN+^Q4L?-WD1dG+9B#<UDD3HC#YSc9/BO)P^.CD,CVXPLb
D18A\2HUbN]3(DaUVC>OYP=\]T>3A7WL8QI,g)E;:6:fHMNa_O\AN.#_<MA<1W#:
.+4#VgaG#QHC6_<5e6A[X7cL&B2R\=\IKeF,#UeML=[(Y<eMZ][OEP2aTd/Ma#7B
IgHVJ8OX?[[ND47fUZ&?+(fAV1KSb3A(]QaN5<T(_^&J8V#52fK:,4TRd.L#fF?2
Yf/BK(]BME#9]I(Ca0>](K?7PNP@f)FXZF;-g_S<JV_OC[1N>bZg4M).YPd^bDII
SD/R#6P9C=,2TfKfV83f0V=U7>7&g;9S4B:gVL5DVPNdZ>Ye4=Q:e8R-Dc60f-=A
d>6?W9#3X:/DbA6gPTW^88U&_;-.NI<S)f[S/Z.;8_PT]E#@/@P-<eM?8CWf#/2(
L.E6Sd&S@\Z5^+dZKeF)3DJP/DNM4S7@+)X1b/ULDTaPcZDRf>e6@YI(/4)S;V(P
WR=5d;@dH@Ed:O&C^C0:(+8H>]BKN(X<dca)fT[G.Z,DPc;3SDc/OJLVSL[[_7+^
T3(WGA8J-]DW\b2Jg7@7<1<1;PL8?/;HTF=RHL=-YU)9_Ld6#RR-aEKSIc@\C:bS
@M?MZ);C2a9JeOdJ_P?_fB<]e]9FGa(@B)?N7V2;WdXAf0IKS6,OBTP_ee>_GKR6
\7<gQGe?fUJ#?R4U;ReE:_>-OeYUOg73C06P0Fc;591?O(-A](3E.fId9_G?&P.(
[?&Q6GB;T0WI)0IT(&GQ8;7,X@Y>.5b>76Z-+3>3JKd],cD^<L_XWSU4I-E>bQXN
NGH7H553P-6B.J)C>[)7GEHVQGX@g)RQgDP]ef]L:D<4ARJ#<:29M9^>;<Y;[4bS
G9FM/MNR91U8[(e1ABN4&g-\67JGQ;MURDRC]9;)DRa72AA]]KFdLPgP1)S?W:9?
/6J5]3[NfF?Tfb7L-I5dS@^AZ(M49-e31;XQ9]&B7YDZO&R8FV&Z0)@/:<UIIJV=
-c/f3AXPXJ^1YH=CD[MF\[8-V[TX>8+Q,;\Xa@UYX;RTCVI@)A&R/>)a3UX.S[R<
?9,\>g)1AfZU?6(]5Z_d-TK;U\X-a8IJ:2UL;fNCC70Y^>#.B[]VGaBdG4RD&/HH
GY]gb??g6E+#;LFQ7802YPd/9>Q&7W.1JZf70d>T>f#O3D>5d^[JA2fTdIg&#CEL
1@FXT(JLV^LCI&>cBY@IN61LE9N\QD2V@gFf1&5X?bV+\Z0GA^/C06Y=PZJ)ML-,
bH>8WR.?bD<&^J(^J(O<ZE-f4KFBY9#IKZVH+T_aIUJI_1ORR(-=R/>&35B,_EM1
L\9#(3;P8YZ?KBQ?]3_bd]^a+]M_]H(.2_6028K;(9KP.ePS3J6@32O0X;Zb?C=f
UG/^(+K@,aFZ@Z=11E6RGFCYNc^e7J1#]gPW8f?]XN/)EeE+7+:[GWQDAK/e165d
3,V4(f<@b=6#ZR)I_H=P[(Qd;JPXV::E(MJY+F4dafW)MRdJONGK1T]UD)(.COg@
[F]T:CCZX+Z/cKddKJWaK8a-Ae\BaH+Ye(W1P<F[WK4b2<14a;b#BK=V5(36]\BB
?K-)7f3Y:QeLX7NZ5XY>9VTfC0^/Q+[Ra@U=#BJ3N-aJ,1G3Y<QYL@C1@ZG#d21U
)\NUU3ZWH?b5Y4,8Q4W8A0BGK<g021H_[EK1&)aOQ\;.<X9[Ibg6Yb2Vb=C4\Vf=
EIAT/M^BKR,>Gb,2TK<X8.^?[g8Ga?:BIFHRZ(]0QG#Ga(@;GBFTUd,5@a@M:DEB
S]?L5Z^eLQSXPZR2E0c/ZD5Wd3@cP++@4S#W?Jb&Q;Oe<=(C55aSDB27/aBc==#6
T/Se\CW2VRZ9U(,2:#/L<fQgAdY\+C]cE@,Zca67DE4#=ZH1.Q)aW;d4Md\S1##O
ADcVR+A.V^P<W/b&f9b]FP.Z1Mc#_Z+32ba.f+.K#KYa8\e5U\FR+^]VITfVNQ7f
VHeGBfY^d#/TX<L3HT:D=[T)U#7]#g^(,g\ADI^3Ja-M0D?;VbKcQ=9U><&(0\K4
]Kb])+J.NRE>5]5#S[8f5@M3SV3EH#1ZS;YAAH+N@4f8<O:7IJRH&2Pa)HK[T#WR
>#1&)L>C4:g@YcNCP<Jb3)J@F&?4Zg_0.EEB/NIa]RG=<SR(,eEQ.bS/I,_XER\:
[)e9V2aDQ4b<IR1JX6R15<UQ^;+HUXIDS@2WVf\RR^)[S[5B4HSbO]R]MS,a8a7:
\5F[6_0,<4Jef(658UPDg9PYJY_3cT:72C3@9/_GZ2&3_N5Sc-KgWOF\)]&0OIJ;
(4\P&>F)K@^aCDSZdWbfBe+1NBg)Bcg0NFb8CQYfM6ad/gOgHXY-(_DGG=6Rf&DC
(JF>dd+gB0)EH5LME8AU[SBWad.L9+0URWV9H&.REL/Q@=CRD[+dT1)cFQ#T2N?F
)gDU4)+CbVbP\XOT=fKgN1C\D697H;J?5=NaUEXHY3OS#N4RaC5&VV]UbM&d]W=]
N5ITK5L1Gd.O:PUCECA[a)WbR[X\T(TMe9M/+(_SIN6S+M(PDMJ12FBD.4#<B)f=
\QI,9::GO.A_GQF(LaSdcO1H_E5D@WN1<=-D-Z>P.gZEa)N#77<WQ<EeTSX)]F@.
GJgN64c>JLU/>U,NC;eE[>XGZ+AU@T_O7+E(AQWb:\OO+@?6G7L0]K(I&FWO;6Lc
(QC7S[L@,^1#/3CBO(-Xb.4#-..Y^+[?#XPAG3FX=SX65M[g</dAW.]g7,#d6O0D
&0+Z([96PfU&-^_7&9.c7GD)8S[+XGCBC.aGR+d&4f3R6K@8aT).,=86413:La>P
fc,E+JKdQM^68IGJ@-T:F_3QaBPMYYJ)&SV5TIP06&+3\9>-?2QNbF#)8PeB#e57
^G^WZUSbAS9c0>_Bg5WN2Y,X1(9@7,>R9SDHX\/LA_34b9L/?d,7.IKZ+^OS4I>O
(^0Z8=c;X_@POOZVdQ?Fe[6IDE-bg]/]\++)]AEKB_6^^EU/O]A0-PA4N/=?#EdS
g6c:cRP\D7W1>\MW_9?<bVe3&(:aR(V09BS6G@R[EV@-PMH#(QYBCL@f6E,\<g#f
ZMa][1=gTfYO?^QSGMJ8e2d\Ie)Q.DfEKQ17G\MG<QDC[7>,?Y]46eK5g#G]9c+8
Y[.Ze&+S@(gDLEG:P^^XF[V6?d>?=dLVZ<2TH,T@Q[;^SL2RF5f>cLDBYJXXKH_a
TT)85IBN:J15186bNRe09@7T<b-=]e:d<3_/1)^0+g8NaIcTd>UDXHVGD.WFN;5M
B:6LgD\ZM),cUJCXE8c.+6U_5DK09eDHDI:MHFX]U.<6N#c^F6-YQ;3\?eG@]FEg
V-W(f)EXaLa9)d-Fg<48OM4bID=b8&<>35B:Xc;]]GY]YT(4MH5V1A3L_C\ef]@[
4a_<a3f=&gW<>D;W]NOL?(1Ag8<8?WMC2I9-IR-.4>W;bD7R,+)N(QX]C,,8^@Q&
BV<X8S@Mec?a/R@e,:Gf\ObA4LO(?KVJV<B_8_UR-_a.Vg0RT(.a;M^2K.T3\ZZ;
=F12OJZg7@8>]EBf&-bRQe^\Nf5c)V,2B8RbU6I#<IYbg\Le&5e6:VHDgEfO7AI_
]>0cL7+[<CJ@8<M8\D=HLOTOUUAZ(7]@]XNEF1IG8;>/\RH1;7Rg9I#4:0[9f6Z6
b,BM:-,bM/\3&G=#Z/<D<IS?<WCfN(,,MQW4]d>HNDML>BeBbTDH:FHgFVXKO4_=
\EV[,?/W0\AM921H\KX/#LeB9R0O]EDYc4g;O^5\]2eX7>(3g)@IY,_J8XV][^T)
QG0[L+TT+c:DJcX]:Z-/\NO+F87TJ;)^^0cX(WJLU8?8Rf2#OO,bg4:SMQI,S]58
FS?;eIf>2D(gF-)cOZDdIC6@2\cg?9U;DU4>4BD;K0\V\&N/DIUXOC0DB0bI<&bY
RdM3FO@<LZd-Y=T<;3>EM#(-_^:fEBX@SfJI?9]:3#MABDS^2.Ib+W)QBFR>H_^U
#WZ>50X(Od[5]1CCRD_+8GGAeOS==1.R7f5BII@#<O9F4V0:Hb1(;-89bV3>3<WW
=a5[V2.WabTe9.<;A.RR_+-5Ne[cD-bYELF>3fVb#eFKR=)4N-bJCT2a2f>+/:a2
[^DIE22AOQR3^4O3;2TU#cBcW_S_UKdT6>L<I1>HE/]52d5OK+f-?:Z/,DF/PEU,
EOEIG[^G3d=-;3)M@9P=QKA@7@fBYb(2G&<6#SL81<NZZ-2M[@1?dc[.<#AM:c+Y
>C+_0b2VN=(&@?&-RW_)GC5=^>;^:dWM,gPIf&IX/(DQL\7^#XbLO6F7;M)]_:7R
\LCbJQ1JfUI8Y;,P,;7fgR=dS.CT@&G^b4=<4Qd-UGeD25N-<;6W84JE.b;WS^1V
F?EWA>XWA=6#dXQ=#@\f;O,AS[.gOXLSd-M:N+acK#@\I)Z;>Z18YL8b4XHC3D#d
Od78FBeQD7P9RE/34fTGf].<&Y;d=Q^&a&FgKBB.bMKSQC<A?^72B]CS<#7HQd[;
QGU-9bTZ.)Y](;&G;CNVAL[,GIW4LH6X9?MCUGU#2+J+VDWLRIe&0dGI@G:[HHPW
J[I@?X?LVHdG/^OLS2YMJ_OS&b(_AK23TEQRKBC+aD,c:g7S=J[KX[FX(WN:C5HR
.W/&05-8QG+0QAA<#D]G-^)(bI:^=VVH23f\d[=ELY];eg4cK9S)H,=F(7/B&W=#
#&LIAg9]=(I+IK;RSM\<b\FPMIK5YIO,1&+Z^8gWIAO,A=+K@84?ZC=bA+SMI4gP
_0H9=,?f/\/?T.X6X&=#AG;Na)U4FZf._-],-TMN>77@N/-DPN+?\5[M/),]b,a(
b@[/V,MHgUX3g0NaAe3#AC[D7e=IVA[?9^813SOS22=(E-D1bECSDCK8QO^fRC&5
-T7[PV5[S=Tcd9/ESGSV+VgAKT,G)&TAXZR(0dSeHae)_(+I;L:J+JG.J1.Vcc\P
U77S]F-9,CJV6,HMf8SSXK=P6454\S+1+4IIeW@((D6II_6KDg7?2^bC&g7aD+2Z
@.dGZ3Yb832GU8,A8U+1:bbe7L^TCgeQ7^ZVSC_AKS=P?]5b)+<^W--aQA^BO:\&
F7LdOJ:?feXI&,SJVgIVTU7f/^X50S#,J2DF?Y/M088T;+DH]?KD+#ScVBXD&cX/
5(DD;N1\.1Reb(B&DT#?fgbU4<?YCY>N-GNIXE;M(ZG)<BN4&\efI0a2?K]1?70]
\Pf-N5U(=;T;)48S:[6^BXbZO&H5bE]Ig?.,cN;D-f)K3NS?(+d<>8??:Z64gV6O
afS/R.DbC1B<_Z=GQ/A9&056QYLO7Zd@N,^:C4/+=>?\.&=TBgad]YZ>1L.Q.<gC
S@dZ\(agO>GU-LL?dC/V.KLWA;=(f&XCHXJ0IUG#KKCLF&L>A?PcK4<W0dOd,_3F
UGKe9@>I:D^1P\5ANJFUHa1<C,O@E7>U[P;WG>WV:;/5>Y9D3S)6LNPZ^AO+Ac.X
K_fIMJP#NAU\,<\TF1(]EX)b9]STg1)[(gfLECHH\=d0F5de2:8DcJE3EbOX<#/.
bJ9>-9B(NT4N?Z2g];X>4b7DO,=>)9TJ:G9ZTK0WEYSMf@)&UHE1Y?BJ5Z-(-bWX
(ddF>EW&TCYe-6S#.V#LIHfaTD2+g@]+LON85P6SGge?&V?^6D6Zc<#HPFN1;.CK
cH]WU<\-0gA5LMg=b?]OAXMJc8^IX.Eg?0.Y_+F;/ATV(SVMV&ZNKaN&KE5^.XAf
0(<a(X-^ONO)EVVP@MF@<S#aOV-V1)++.]9-F\/LdMH1_<N>](MK#dKYbdVYCP#E
>e_8]Q=JMA:>e+Kc+8:AGOYW@f9RLW>7cM6,/9-eV>6_8GO-LO?<Te#;^GA-/A)0
6>A-9@DWYDKbWg1H<8Y<QI4cS3)=)DFEg4#C(T(X-f,7M]aB2Ve-OR&5[0O/R8^<
^P&0N=3g(Ja@_aEcG[[##DWFMQRQLYg:L0(Gb49B/8_@_QfDHEY56He8HJd)I+?Y
gQHAW/LEeQH11]I>&8YW@>VUed;2OKG&Q<I->S&]Y+H+(@.#b^/ZZ(0<YKMPY:W.
:?O(@1DV7/8SE<e]#@]O9(,L)JTC/HEIXfbFZ@FV.6a6-+99.;?C+Jf4;)WW^H[N
Q^gM(-<(MV]PRSJ/2NXfg54)YZ4_/LMJ>PAa6N]^,?fOfa<a_IO+;cFfCLFP]ObJ
(e2(b1@V.?-8+ZBDU[FMN::@<5]G4f.]cP/2_^?gK<124.&R1_1]UB=9_)Z4Z-/L
9gD-=,W:4\P[e:R-MU^_OGWcJ^C\O&[UKdLS&YK_M5#1ed#.P1P-G&E</g_+4-eX
P1^XFa&6f57[fFaW:08\+2Q=Xc..T]/X2J#VU7-SW1#UXa<J<L>HP<:<+b0&XWY1
1S.<)9W-W9FE,6>.bR@#8U)/Q5cK?\;@Z>;J/RPH42KQSX#R#2,JAN&a_O25+5CZ
A&fA_=N1)>J\5XQ9EB\b7>;RaD_HHc=F8#O8KTXNdAe7BOO;XYPA_W-^3T/d\2;Y
f0[EM2ALF8IDC/I-b/R4TP4WTRZVQ7QDQ?S->Z(7SG(BH\&?N:Y<1]849+3?2YF+
,9,4M+AWC3^M[4RA#U]5.Q^B44)>X-##[U@S?[5I)<954SCSMP_JD.E1<QQH7AbU
P:5[83,Yd(B4S6Dg(IF1)ZLDJ?N+Ba1bScB8eZJ-,0<1O-:R<,\Sa2YP=XJ39@<-
H:1ZB@gZ_#]2=@ZR>+IW:B,.6L(MMUdR@L9TKe/HaB6Tdg>=_V-9.RZf(<D[?Z6A
,[4Y?;D(QTY2gI7.(^H^bH/RW^&.D5D5P,XX(TAdBXOUO(=MHD&HR5/8XBc8X?@&
H0gAaLa07@e/&QH4b7d-XLI#(L;A(JGU>;aK5]NV)-(+_Z:-Z_=84L0<cE=?2dM2
CBCK=W2)Y];+XW5N,8VB8g;O_]#D;:a,M)NP-:]=9@609d4U&#fcH+:R8N=/A6-^
a^QU(cTdMg_FDK^,XZHXc\T&^RG?N>2H1\(aNcX5f+1G71;eH@57-M_IM#R#P=A.
:dS,e;2P2X[,,_B()^_I)RZJ=Q5X+0CTG7gL_0--]WI(FNWHUd.f>/9(;V&41aK<
.)SS&O:__G7H5EV^E7f[XD_a_fgY5TQ\g=g&MfU@@G_Q[:??1JM>KHPRM)&&Z)4;
><,O>R-CE=5aM+\NbX:8BX,BY)N()Ng&ZIB5?XY:^F\S?eb7g6?I2?<F-P(LLNIS
e:L6F.:\fU&G9=NJ=\&V5:)H3>[7UEFPIUgAI82V19G/>)JXFTaI.2D45Z_=bX\G
#YB@/,_,0TA3^eX73d_1P@611EdKe7O?4IA;abe)BZP)E>M[+#QQbDT.>]5^K81)
Jb<[;32+></;#.HZII;;+VM.-AJ&UEF..PH=##KN=VEZ[c\EPR.@UA2KHgT=Cg[E
.17PHcW3P/4-KWG#C5&b5g[f8IO]dBYI2E6aOa==Aa]@_X1&KEL3ZV-g(C(_O#8P
VG07JDP#\cVA&Qec+gIKe@>C;HBKO8[3OYO.IS2#\d8gL2ZCA[ZL/IFg(2&IGgN=
2?A39Y/N3-8<&\^Og),-&(?8)gGF6:53-]PD\BZOKR+RTT:)#750@gafJ42=WLgO
<HETf^QOdL=fSfGg@(6/:].A7,A()2H8,379fZ=[FHZSWY[>Q>K07(a\H/WU<^BD
fYWRDB)^,;)9fR>K0&XJ],c2Y:&6LPE=+/I)(KRBCaT@\-da-[bI7;QW5KB-.6e<
L;WMR=Y&O]#</c=Cf-GZgS35c:UT7b\I4,P/GLaI2I+&7A/7519^cEXJ&/,OTLC8
^NQ#L;4#F.[:cgd-+A.QWfZ:\^7_dP[O.2([cQ]ZCbI\12@=ZFT(S5gMH@+IJ?S/
6578:g91:]_2dNCYE9[?ZWa2f7V\]bE3<>0/UDE,A<I:NW5&Wf#6K4:BR[ZUA:LQ
.[PXBV>AU#5XQfTVJAPFP^WW3F[NfY[5eOT4D7(5&g<?dZ^46aQ9GOWMI.I2,0/H
CXN3fWTI\W,EIf2=1@G2^G7e4E9_&.?[gL/31ge2d9OL]^FU7b34JSKX.;Rc#O(L
F0MF7EW6CV1bD1OKG-D;@dd_OQ/L>/8AU#HNX0G=CRaa/B<6e(?ag8@GL8>2>dK_
X))DB;&QL7B/@@>3<NV]]5NHP8c1CZL=d:ENI_ZNYVfU)bW4.H);59daFaN#:BSZ
>]M<A0/AE9VMf<LMS)gJL99-9I4VB/58]ZDN>DU(MWTCQ4K;E3+BF11>1>@/T@+,
5K6\Xa5X9:=GbbcQ6:IeYO9/78:WI-MJK;8116egP9bfT8E>F<H6S7,5aHMZVaGU
-Odf[,B/Ub=)_e9cD+(8@8U@N4M+>PG;FQ+2ZH#3)fILg^a6Z6>WgKCd-I=FS3I?
7BV/-+L,I/aLB6J(2f/fD1KF8=RNGd^gV#A<VSQW2MS:@1e9e\@J:6gO9@7LDaBI
&^L5Pd@I1DM,M[95[J/PX@6JfS1@R6(e/eRZf:Bf?B.eT:&E7.ML[=01(fK2eVMN
?T]78J,=L8.1H()_Y;HO)f6,X[f2@5HIVfBG?X)cN.K0f,VI^14[-230L35SWdX\
;_:4fI267(F5Q6R?:75a=9f08H5E&D6YIP6b6G1A9ER[N9,&YaT2MQ9G.-Ac-MB_
@c<4<D<@2SM_J&_UDYENTN3d0gf(Be][WMR#=DS29YI#&afB>E26UYb=F1(#Y_Da
7CZGcd^0Qgf]WE7WEB1RI_5X&16,8gG?)9>^R\TS<J&L<d<20<^O^8[_P2:H/KHM
DdBadC@74[DYd_2OcbS/g?&BI:IcE;[E:JLN\#\cSO?g<W9gb.=4T@[.YS7^^<:,
gUPf8(H74ZX&1MIANI_UBf>:ccZPLG/_W^_^[1eL72,1:Qb;VW@UX6SZ[98W<4M,
-4Sd3VRe-:1bDBTF(d_S/WLZf)T;HZU:0KR47#d_L534,F,1RQ_OQ^LFO-aN;5dX
e#,(C[Q:6(2J^bRC8G-K>cX<,a^CD[^5TNbZ+;UCDb:MOfNPf(61S\Q([4)XCR5b
e.=Bf&ONE?]KWXK[D=410aE4=GZ_W=(#\VB3BdUd03C3[EcZg677GT=g)=Z9H[Rb
]I^e]_8RM:4+>14FHb>Ke6aX9dFUCfI/UTOJ,1K]PHIOZIc(A^)0AgWEc(A5S3ZQ
8VT5I:c7:FA<KNTZL_B2WQN>,NLgb^(MAQ,HLI_K=L5#e=FYDD+]M@IaNg\c?=^5
SNQD^F/OFAAeG?9OB?+2\e26S/WgXbYXC=AaaEC7:LP\IO-gcf9OEO@Z9.@gSa(E
::BA[0^3D6]1,b,]=V63.I[>Rd6V-1BYcXEB+CVNDO0_5dCJX(\6BZ>2?J@g2T6E
(JEfM+)Q#a1L5II:^gB-&UL\4](XQ6V7N0]_g2QXD<#;9UNF4.I-I,YC@ZG2W(3M
:SH[JT0WYDF)faRRQ0-@QF;gF?BHSZ8#HT-E,TRYESJ=f<WN5DXTFWE54G_;1=1d
>gbR)OCGWYeWU.DWY6<:E9D.HV[U@fQL3N_eBABadWRG[G:(YXDOb9=9_7A3.ZIY
XR,]]^/ccORJ8GU4D0#&7__?L@5<[ENL)KUPF;;.KcL58[#T9XA5[4@&LF+V2A-\
51BbP9MM=#53Y<ZFJ8g&/b?P8Ua](<U5RQANaOPVF+;d5agQ70@7PJ=3-+I:]DeH
#O^5;a:bf^MU(Ha&8GGG+\-7])W]W@C<3(O&^f;Ag8a6;OA_Y1)\NU3?#N:1FOa-
SPFg=.I\[,N8N1OSXF5TcC_0>#^a#JGRF6\-F5[GDT@QG4:;ZM(D\3S-7BG0<O&]
g&a0(2cE@V,\dC3\W9aPQ4Z#X@UL7e,&<1;==+N:T#;-RYQJ#+N?gC(2#9_UE51I
Rc?N&VB1OB[ON.\Z/4P]M4EZIMH.09ZVX_^UAOCF#_\]Z&0X5U;Oc)G+c2;5/E3K
aOK?P\X9L4@_Y#@54PA&9D=^]X9G8#CJB9fKJ4,[>X&@RE7LO[Q/YYY]8AcV.-^(
3KXAKK:dF+83.JY=&)W=fV.Pe4.E4RL.6bf>JfZYDBdKSAa<P2C0bLS4_9&IG^S9
QL)U\F=:gK4Vc_e7N.<OLN#;CU74QX1@Sd-&aYfQ3X1B9LB^(S<a#)NGAa,3SX96
]DdFA^dVBWd:He?>L&e1Z=VEe.TFDOUHQ+@0-QV4:+ZgOSJOZD&c^N)E(C;K3)[Q
]#TS0/HX+X\FY>N]Ob>.@Y.(WKUe>>QDP#]KT^/eMHN=&]GA=P5)?5\,T54;;KI(
?;69DgSL_U(\8A]P6EBBUZ(A0P.CfPVMXZXgSB;<:@cR)YSf1b_eWY^WIF^fY_N8
38Tb2D0JGE3.f)6CFMX4LC&7OD9Z[Sd_6;[D]\8GNgW_ga&O-<E;2+FYSdH3BWVG
_:65O=6B00?J<,HW4ggFPM\)cNTR&\XG=]DfgWQK@D=5E;NGN=;Q>5;Oa8Z,_]+T
g\gCYC^)?E>/+F[4W##E8AHDZTQ/721f[;Mc^g=YLQZJ#@D:^)g>c[@&4)5FR@^F
:,-0f,-.aR-Y9\^I@+^.L^O26,9LA^=D\K?1?IG07UH4QJ)]cA#-0VL:)5Qb6GGJ
[H@?)&&YZ4+)f:H4X7HTJ&L-J/74QX=FdG<2e.L-+bCNQYCcL+a.D2<#-NBLY5].
0-UG#>a3=[\B.Y(8C]GW;#O[KaUUKVc3?VB;8CP(ITW)cF6,EZgL#(L@8#M?)5[J
1)FEFgcC<\M?2YF49-CFC-<_)7dWM)O4T:2e+NF-(eCO_#HHT<X.O5DaPV_8fCT-
dK;?M1_&4dB[b)5_POCP#/VHH#MGSDg6.XSDAHgg0e6P1,cY^O^M0_#[E\cg[SWM
-M3L1RgWWaKg:SN1PPZ;_+d@2VM0J#cg^5H]0B5PCd/36:Y#/dK0RQE[N_UY)B_+
5T<3AfETA4]<)a-HUMD^-1/)KTKV=_7\^cgS2_[O982.[^\+KTWN=WQWO,HLgN&R
Q#JKGEQ98#U(M;PJX>B1K>ZX,=3+:Mb,9NfLcFd?M#U:542S4LV1/5A(=Wcc,?]@
NfYNN0&P.4,G?a2VG1J?G+eDa;[ab.7<.T?3A.eeJ((6)KFYS_+0+.fA98;-/L:d
]1Xe>_6B6B6;;:;#VK>87GIZQIg4]3[_&.LV=FCb(<gR)>aKZ_JRYCa<(0MKI(5+
KPXVeOU1gIe1,MSY_W=&<4-SVJ]gaD5@<e:);BPa^LJQU_D\0Oa(IfROZ-].^R17
RR832WF>Q3V.#<39A=1d&L6S<ZEL2CI,/f_))F6#9[a3LY@@J4+ReQU9M1AcMe85
JF-^<+eN5@b[BE&U0E<&-R17IFcB,g#[>D^>D^eLM./8Cd\YM5RDLeW4L4e;YG5a
:9^NVcBL=A:4a18QF>(Bb;-MR^[C0:+X)RUY=;#1EZLXb<HfF[XWBf(.GX515:-C
5[&:f8_GR84ERa,c9;cc+VLbO,&_X(Sg:1=[>bLfg2.X5.4DcQ@\:-R]#cTSY:];
X>4/SB^\500<MI8X3dS^XBNA/DDG[3dHV.OA.I9XB.,5Tc=\31K32)DdCJL1Ib@,
],3:YG\ECXgNa?fZ+4[^G;U:5L+JVLI09ce7E;d,,#K?D)#_;KSI(^>LQBf>>B.T
@D>GXW/5/,RT7b#cd&_5H_@NTNKS@K-CXICT)P\?<B/W:<\@<bg<DEA\,(O+<CFD
2A5G;<EC=HXL0[::De>V=\OUf2:M[0Qc50]PeU=aa)EDJ3g\Q.VXHD:5:V6_^X_<
fY8KgN;6HcFc#F?<]==0R7W<<(>Z8gf@?0J>f[[5^MR&5Z.VXf)L>O1a1V>,aH5Y
Y#[K9EfB)27M65]47QUfQ=7QNZUHF^19E9>M^bFRU40_:FfD0/8e#.aGSSSBM0WJ
](EY<BJ_-FY\Cc^NHQ>S,V0FI2\4WK+Y50A<N_6(F6EH<[8gT0TEA9\&5ST4g8^c
@eHLO4],9L)7cY(V9PDf5C#ae,3Y2,e;>_AG9D6IG37IT)c8E+EQK>Cg19L^LWXY
.@-6<(U8G,P7[B7/VGG3+IJM04>:QYH&<?^eOeZS:.aFSL,D04QI4Z8JV_D=#N92
@JR9/aO0]B\@)K43<4;JJc3;_Z)4T6TXR&NaB(]D\aAHe2>OOS8\F:;eDV3AT9:<
ENMD(CY#f[D30K[FgPV8G=eaV?JY]6I/^Z&=53XN..I2VK?WFFFB3bYA<ZVMID._
;,HZ,QZ?&FF4/edIVD2Sc+V/T5_C4-NEG#DEgGb@7\^#]GUD<3;eFZ^:Lb43c5=H
\L?]B/,YFbfF6WUIRP+21+^TTB1QGII>=&+KILIL4N9RaQ?eR[NVLW](WE2-XO82
W-8L&Y?e+7EQD:#&B\9,f5<U2^3Q&C#O(PK],-PWS(+A:.4G0#X78DH-bZ[6G@OY
7?Qd(?b.T.:C\fHZ=,6N;Dd/.aD<4Fg>\G1]:,^.G#,6Y0>M4B<D?Ja=)&UZ1[Id
8G>Sa77eCL+3-.fO)<Q.WdR8T\>(:.;K&C8XFR_K0a5>K&],LV3_(@bb#S)OT,U+
#[YbZ3HfGgSPE-&<5M\)S=G3:&2.,>@[Va4L@3.<+(2(,gE[8Ue2GPdT)gIc+UM?
>IHgF\SOFDY;b+\+.9CIFdYPFJO3GPYc49[4_GR&Z?J6FJGXW75U3?DBH>W85ZaZ
DXX(P?OdZaQQ5T&NK,G_CMYA2TS=\T-Bc(?aSUZ[FL+>R>977b-cd5()U4cA+S\4
28\LRX.=Rg=f<adW\2e:(0dJR^Q<C@GF9&D\SANC7TDZQ0YSQ3-:M_3EONT78LE,
((\Yg_==W>(XD^IZX9eAc&aN,52K2FQ]Y\8Ra>.?L5;KXVOa70HJ5E5=+g[+LA=d
]NI4K66J4&Q?(O+ON^VWG,8TN@:#gQfUDK_95cX]ae@@e<;1:.Z\4B-4/X4N1aOM
T693[R@g7\L.;E1V&eQ[T0IU^Ba.SG(+@,<#R+@4HZcUR=WMBJZe3cZ(?IL@4[&0
XN^#^I@+)(VW)d#;dO\J#\f7/YXT7S3GI9W/Q1.EU1<^dAL53(_A8U)SZ5adDZD2
->8GgY01ggLKHNI#<AKDEGR#?\b;DVZSad2+&S/^8<IO_YZKDdROaRA6[;(d;DK(
DCU[b)8QVbN:Z-W-322ASI&ecfQ)QVgU4TZQ[V64@6F7;X99)V#?cDA?=c,V^R36
R^ZT#/1AAeU<H&=7:/<dK[e6]B]ER0A)D;A3=8:5:)6a\8fXGdIGTPf1N2dT9(P_
aSF5CV4);gTa,b<0O=IL0=Xg>#&+/,_N@0[.8NH2gJ;/H:e]cf&.GK+dcaO)N2,#
a(5@S=bfgCfI@704CLcc[QeZJ3(RVJU(+7Je[1CJG95/6>JGY3C3d\^](dB^CQaB
D#PP9Ue(a65WCEIPW.20.M;;YFX]GM&^1?5-3gR#IYSCcQKHA4/dH)BRbM.]+;^(
Q/O&VcN)6G6M#C/201RIYQ12I^_T4I7ZQfT#IFD4+<?0;DcGM[5MSN@Sf^9/8gLC
QW5&HLE35HQ>faMSXdUM]T._[W?<)S^2M<^+LF_a;18D>gL5b,S@1GSNScae\Vg+
aF#26[&&,<MegJ04OV?a7e\CEB4=cI/B>USb@K046c]OV:#;#[?0R#Q@CZ40QSI,
7:95EMU:7YKL/U,M_+PML-?+RN1bg6EL3Fg:S@-\&TS(J?#g)Y=R+/@:#Nd1J=9F
E9/^S8)FTTT2_>DY#EFE3IQ9-P28,;AS0@+\Y>6NRGR-#IH.F7?F;RVIgD8I+,3)
J[5R19[&+Z=Wf_3@?b05\3:;:M@Fc-_1bL,c1RW:E;^:UgJef(8[[8Y-Fd_NA.T[
B?Y2)O@:(fB,BK(XM9ZGMGX=[ab@g-;dGH1CW2F^)PH<4+f0,#c-?078[EM1ELQe
)?I,EL#\LeF\3,aD(FS&gM71PQ^ZR>b+N8[b/EgeMfMb)#IRGZQ>T;2JDg/+e/:6
-95QYbZFW@PeRI0AZPA;RTAP?R,VQ.N&3&30:Z6@HHUM@8K;J,4ANRfOGL_5T9E3
^H-U9I/RQ&+ONLg<6XNT:Jg1L+I+P;_WSCSE64Fb:PJK^&d]D?]IZ1G]TVZ[M9[/
JH/2KMMF-47A]HdOFT?=F_/3#ZX7]MCT53I]<T6?;2)L44IfIbKeYce@;\ZGP#P=
RZ(J7AUM,F4NcR3&S35d]V_aDb&NdU:UR+#&dA1VM5Fe.MeCMdeaHP=:eP2#Z7JX
\@&1E96WWQ2R3U4#VLJ8H8V?=TM/MO42#eS-]VZ1EJ7FHVD,8@XL7..714GC=?U:
Z+?19bME:\_g:CHW1^J#^GP]^HUB-b:g&/>4C4HR6U/ZPF4Sg]/J^YTCb96VRH[C
aPLaIAI?=ZJIY6(da1B9D]@GfEM(6)(L/W),9\ZWYNDC,):8K?.bfQ4)4A144eBO
]O(M)<;^Z=A?1^CW)7d_@>@9I95ZOZ4Y&^0L:7CH)=ff=SVY=(/ReZ,gXZd<a42J
U[\1g#/;0LV:M4SE9ETNJPL/[65B(-0X2L]=95Q)VS-KPZbfDX]O/(-#V)42E>5X
gO,ZOd8<<L3V4a88<:6K@D9+FW./R-KFYedT]2:Qa0:XN8+?PLB=I?FMVE^Vg\_9
H=DFNdJ<>@(^<7a=1(4\9X8D8_RZ2,cGIA3][Me7HM8A34O@YZTZgVX[0FA#^-7@
)FN:E3ZNYP<QI=O7ZJ7SF@G>R8BS=-a?UGCcUY+Ud\7C04e,D.ZS=+Hc7R<=T^CE
bb2UEUeWB23<FD9=9(7E(R@OeZ;(E9fIKXaQ\=AK^YB?eX_X7(f>T7,:P1f?=N<J
NG>dZ/J:JGFUK__NT,@.&E358^IDeHW<PYUg0I=F>PKM8D7T@fRJ(Kc8#aEa^R]T
9Bg&?C4.f3[7=U5Pc\&6F#OEO+5FQOD?T=MQM-A3(\,C190W+DLB>#Z2X-UK13.G
bfgMYN?63^AgM_IdBe(+Y\#EK;DX_AQ7([LPEN_U;6\0^\B4,0F#X.#T;[T1Ig=[
QE847BT?70YT#91)KJdZ,3C/)cAVYe\3/2+VBNM?)NB<]U?B<bXK5,#B119/bN&(
U8Y6:36DBPA_H#;c90J=#fYEHRE@W;6f47:JUMN1@/)a5=8#D7/WR831fK]aVD-L
ccEY[;W&S49EHC=#_D0cPQ2GBd]a:8.7eK:4?[)#VO#@V94.C,3.7UZTTd7E/H7A
N[:QT=XZ:]VRRKDIT;UbC&XQ,X<:4Kb+Q8ZW</,Fb42B.cB>VZU7RJFCbNHI5XeP
2VRE[QEB]0#D0G@2NdQD0Sf/-DP+<)LUJPL9dP:#Yd\Y+?;(3bG8Kc&f.3&R2HU?
a96MSf>E#KNL:T[?F^P,d0_E9-_Ve&VY.)JHO@eLXZWL_#\cC@A]<KU0=Q;=/D)0
.)X9J.XBY^H;82]C:AN)fH4]e>b3HL4[8Udd(GF)P.5ZZA@NQ_6;-1ZcRJfg@)eF
e8agG5)/QWA;J?D)LA#+dUR(1aZ6TS<SZJfCYF;G>9WM6/=_dZ7Q[LM9282MOQO0
WK?:10EK&0e^YCS^/?T@GO9XT0g>=XRZL2<[OFTFUA1V/G6Ya,^d\MWG4S6P(ULV
.7H?&4S^_6cQLA#^0:RKDDT6>A,.VMQP)-D&CU=.W<AO+KPSOR5+2g#d^RgA=0@9
?C^/KD\7_4;Pg7AZ.AbF=C)ARYY:DP3&OV<0>_[2DS3&H70R[3f9J>_22@9P#C=(
3JY;bLSW0O.GHUb4SR)>E^Z#D(UdeM\T7Ub>STe4YF.B:_:1AC>PH7[a[(UH=ERU
V:UU8g:QCX8.>b./I6c?V1IZ<GD.H\?ZDRP,7bRIMNG:(?&fccF#O1fdc377[Jc>
e6YWfQA)@O=&N(+/:6YS5J?U5MUg]Z&DKdfT>MeG000FA4+KN(@dD?S5\<:0KLSg
^0&(3_3]=>MFV:AQU4J^XXW)UMQ\GR@bEePP72@(376Ne[3B@)H0c]_]]a.BNcZ6
ReH.W<+/KLE\OJF,#dg)?83LgaGR93U[XMTa&c;ZUBKW+YHQcQTaQA@ccb&[[LfW
e[@>.O\]C5SB\=FZg(Q\JY@P41-Na??YV;&E+LBCdH.^L225G/a13eL<B(MSH1YD
,e=Re.,5YK6B(#Z-_^>MCb:JUEVWBG_6e(#&-bKeK0-&JCWMI74b2N8ZY5LBOgLg
<(F->JNd6)af6-bOE)M#RSbM#Ec<gd8:GfTJNW9O_8+g-1([7(B<UC<5e,8H_f(,
&]]Mc52S(QBZ,4LGPNdY3/PN+:5#HTO2#/FOD)?<JHPP?#_\D53?aH&HIJ27V::X
M@>JbMO2><.8f/5+Y@bFP=cB&=3I11^=#caLK0PL\I@ZJ#5feW7W=IbNPaX7^#.=
_QB+I9?=>8R-&\C.Ga00UITTD]_Kg3/(?#&G^+9H(&:9C.6>T30K(>S86NA^<J=V
&I&#G77(_@;UKI2(Q_0;#X^,5Ca__>PNb1cV;D6O/0&L0TO9.e40)_K.a+MDKBEJ
OK)5a@VbS?1=1b/2G-[dH-;&:0B^T.^/F[>^>DZXCS4,4ggE,(1A8@83^Fa<AHF/
_GS&L#DCSXe9^)Ke@9UH3)EL)6Q0JYABQ&e4a[C<MYKX00W>4BbZ.Mg2LGKIc+0Y
I#\,AL(]a@Q[a>8c+g<1YFOV>;.89;a7XRVS.?S\<TR0?,->T#1EaHTC?;#PIB2,
.7V6(6[C7+?P&^SR2&B(JM]2W)-IXHUQY0?JgB=]c8#]+F?SXFNYL5?WDB7F<3OW
FXag2>HPg],Z;JJc;#DE90HH[-@V3=0Lg?CMa1OJ6@)T/>2b0A&B;_^c3V6=Pa[&
PHN[KT#VK5F-V=,[#,M#\2D.ZBe56.AX+gNG_dQ.7IDTfC]Vc(g^#-;aL/4bR8c\
g^[FG^>=R:Pe7K4R&Ag8BbbHW8b.X<LFO#[@9FL8>f47HIeNU:YeG40I&E;HJ:\3
20^IA=E]R22e2]<TWJ]Qf4.HT_eDUS,^f=dEO2P_;cVM@&DO/Yd]);3SWFIMK-&J
DDV]#8@)>b_CA_QAPLIN5gGC(b\.-,DaTX4=V-QF+D1?4NX]Y]8+WJJ,IZZ:D)Ya
NeLH?<c.dNB(>,9WS)=TdT3;RT4gaB0E,DM0eOA0^F9[5[V4EUf?S^;L&+f.R82>
f#(NL/bG#+(b2WJ:H-D)H<#9Z;5)U(dA.]bdaYVc)HGW3ORAK]1\QPX]2NK7=P4B
,-B?PBZDTE.^.?S_\1[f[N=]5V,g:=c:+U5UPH-Z2R5b[ZNg(5Vc4+\XSg()AL.5
\,.\g[JH210E_H]J?aT/UPWQJ)6Y8I1+:G,dLW#XA6CX_1cZNX8ZV)Y\F[)R/c[K
AYC4Ee];cG?L-7O0[A0#V/D=cC)Ug5.#,[)R@NcRT;NIaN[J@f.A>Q,9K+[74@WA
O?7BY^1fSZXW\9PZ]YV)SV18X5]=WB?1[?1U1>@O4B;P7?E@-CC?ZL3HCC/cTDb[
1EIcDe\,+.GC\9,-DJKEfg(1R:@O:RO90SO[8MLL3)eQ^[^1\=[PMX/M:W6>3L]:
/X/:JP<]QKZU,g72a7KZ<dR5^7cZg+NHRIU^^/VHE<cUZM_D;AIZ3;B+V9MLTAW_
)9ZWg&Y07fQ51UI7B8VP&?[V13e-6gJaKVc>)P@0RXH-Lbf9BK6GbF]HUU3P<Adc
X&86g2JEfHRZ->e)6\YBa,OCeV4_5TLP&[VBcI^GB5Z+.A:+8CXULR<<62FB.-c1
3TAO7)c.:1_MZ=<NN/]F3#E9HI-QRf=]=TSI#f-[?eR-cKb\,9F_>_Ad4V#8DbbS
JQR6C1ZfB#&cPb5-[\+I\P2X7Cc/fTK1IfS)[5<C]5e-(T3G1<aEJ;=Q:M2ccNC=
-FL\Mb?,@S6eCVMGNI<9d?E:e[WRU,-OgY-gMNg-Hf][T)aQQ&9O1#5d3]JTg>1\
3H7JKaMZc;TGF76802,]+F9C._GP&ea\5J+<C4QGKMZa;&;-#b=-2=:ML5GeP]&;
aW7&fVe32J)4DZ(bDfdNN;ID_Y2U7CfPZ<-:2A)4P8=1?OHSP?ZF?S8SD[YQWTa_
M>baR5^:-[O+DIMTTH9b\\3,7]CTPHIb::V1,YGfAFX-G^7,RE4B+c;aRSZVgB13
a,Z77a/P&],0::4YOL\;SR#.=A14BbRTcRLBI)(/#E54d4P.J7eQHSD0YG?3S?,/
,]JX2W72TQI-&9?M^KX.<@,G;61953,XG]d\A5+PNAQW2a=AQVBTZ92^^YE@e5=G
[UV^M:I6;N1ef^[?Ra1&-58[ST_2-00<g3bAe\QNUBfVf9(I3K@:U9fRa.6I;JaT
=_DN7b6D,QfZ)R5-4E>@4c?g)=@J.5dTX>/\OXG@(URBc].bRdc7PBG&V0gOS-Zg
D/YL3RQ#+cV_3;LQ5^O9ZYDRPdc\YJC7dIY&Y.aI#-[-3EJ<ZG5<TJ0+P=9#DEQG
:;>Y\/6[PIUM:\9(?C/>H9_KC.#FO)];;Z;C=5GQC)[bA-+N/Ve-2Oa<#9bGYS2<
YS)I&I/d)+=\BOa9SFbF];Q/_17TdP>d^bZJ73cB[EV;;>aOC8<=?\+(::HZB4(=
<[4B^U3#K>[UL?b-CQYRI<B4T8G=XKg)QaAS;2cS(d?bBa[9L;H[5L#\-+&J^/Dg
]C[XUcY[Ncde4aZE\LGE[/>9df7U.Bc[1eEJB4ABWE?(Y)19bX?dIE_ba=HOd+:>
e/REGP&DS509RKJ_Q+P0XBFC(WUE6?e,JD\1>^WR+,YaZ9&5=.;deD<M,6=.U90X
6->=Z4-.fXQY7Qa47A&H5T+K^F6VE^,FRRW-_,>b==7bgD:a24M@RMXS<RUR+?F]
f9SFAPg^.:b8J3b7;R]&53bYME5NV,Q0=0C:X8KH8^4:#CAGPG@\ZL4KVJ\P)L54
5Xc2S[]66H^4f:WCE<((NDMII=M>eT1QbW11.ba+&]b,Z/Z,=4?\Va#;PKgA8&S0
00Wc#&fZP3BFG6)O;9c/+[:N>@J[]Re4aGX8CCUdeT8[1/e\2X4(./=,]a\HE1#9
3X+Dd)e76K=++=V_9MZ;KSb<L]<EXC1W=a@B3W)@>N7d=I53:>-Ff[)IGB^=WA(R
(@HM,d9K,6JAabQOd&d-;)eL\gf)Y[eY]b><_82[M>X&eD4Y>>RNO0\&VU2C&7KX
B#(=AP0c-e^@@#6];VO@7K<P^)VAeVOG_#&1C.gE8JG4X&1Vaa&<E@&Q46I9\3]b
(FbCaS-eC/010Q_.ACON=QGd<P9NgHRS5V23H;K/2f@5B,YA(=0,&&aD;QD)F(eO
:YE[0P\Jf,ac>;\N@RB;K[bC+:IILT;)9WWKISF6c]/.H[>&J[UCdH&GTN,2(F,5
>>9UBb7UF:H<Y^)#UaC_VL3&83;-c19&f8857]+JI?FQ<V\3=8=Qb+[7LV=:+Q<A
)[[2B9TWA(6T<J8?b-]1GZ:HY32?J;F:86A\e(BI17A;KXVRVP\.0X1c_U:H)^4I
a?6<XI.@>HZ6VS:Q[W6Y6[@3K>IQ]=+5cRQQ(,Fd/SCFA@MeHc.-cWf9E)-9\UIG
;@=HG1XK^]P6fD:H,WA]/^_:6<d;c4NfNe_,f82f3BETID&?531+&gaT0/A,ab6/
ST<#/a(Z7e91?1W[BMYOeTSc6)K)(SK2=F)K&MQ&Y(^(RUGdA&YD&G)1D_X5A8NU
,&d5W[Q&65+5RP,ObB]Hf[LXBW?KODL(<Z#f4X-NPHOCgHB@.@a1]fTLG->J;Uc_
O2QeDV\AS[4=T)=bRMO@S:7&WAX-UIa.PPB[A/^@0J5)Wd@ZN_N8T:>DOZQT#CC8
gMO9/+>@8YWIF@+:EMK3^)Q#T>C99BN<OAHd]EYAR3@GR1SP0Ac\#955J)4W<1eD
/)V0e^3LJ,UF>A&#OI_Ob7UWTe+[-&e?feM90HQUG/e>6CY(;eF?Z.E<CC_gOBG#
+Ec718WdEIbTMJBg[U>7V_;CW.1fdZP.Y28-#RD]Y];\6>UC0NPK:LYI&^<0=T?g
dR(6/8-;5Gc)CT:_6H2_g)FD57..]4V&S8/Q[8QA=DY^D:LR/=9;HKEA.G9Eb:)T
,dgcI[&(@I1gRT?U(U1]=#8Ddf2#2LHVF56^<K+Lb?eKg8/1JDW<0P91d:E&W]ZX
PSJeW^1WcT_/1C)Ic>7Q?R/(RSH?KB#g6Y5K6]K>eA17V/:/CPCI9gPT;aTRUQM;
B3S[-X?2ZE=_-_1Ga^O:FJ+YgX\W.U,fb7^6^Q9g/UIW4(7Z\<D,LE@-A@d?e-df
ZI/QceKBRfSJCf5P8M7S+ca^R@DRC2-Z+6O?1;d-PHg)L:K0d9U#4Q;:7ea3KK>R
G+Z?EXB^4P(9>4Q4=(A;<F(>JdK4ag&.EAS;0T336474ecEEK(_O.?EIa2Q[MO)R
432UAJ1](5ZHN(dI5:.d#:P(P>/B.79bZEU&,DB4;/5=9C@:[(5UcK6c6_(f1aZe
\ON8UbXcR:TU,.-+U>J_HVA[A&/_ERXU@7/)==B9TCRYIYbVU@UT,_P>-.[:685R
F#)N^M.>EYSS@I9a[A:^&eE,0KN;a?>d[NbLgC>eVa.MVJ]\Mg)b23#B=#8GQVL4
UP;KQ?6@6f;SAC63+RJMA_9BPTW2NB[bULd+)V9;dc,<5C<;U]<J<UIWe<9ZdAVV
58@/UCT;0W9G:4/Z:.E]ZNeM=BCB<\CGXT)7@N=[^7Ef>^8#YT^SJ7aPW_FY/-NK
TW2TS0JE#40cG/^OHY]Hd?=<9(=AG<eQ/@LB>9R]V+S<O9Y2DF(<F4K@,#Y)SQZ2
VCP-UL4O4=eA?TSaNE8+OE;P7D5dY7-@5NCJC(P_2?7H<Qe^\2J-d+Z2RA)e]_S;
>c65M0DW>b,aAWMd@(Y)2<,<@,@(2e5>Od6dX)&TSe4IIS9-:EZ+=\SX^D@Z0[PW
[EYGfb0?[?\g_Q?#I,.4f_IU<KHIJIJYD>PY^XPTbS9.T#=:^Z=g7X;Z.8#[)_FR
bZf<=JEbVY55N/c(DNc@8IE4TTfXXMCbM)NX-L.1+HCQQ(-W(9O,OYQ6O7R(+@\F
Z^?->#E?BQMVBU1MF;.-(>^Jgg.BbU\OBKNIPQS(FEgTR^+KODSGMLBH=+G^L#I#
<FX/A4Ad4.Dc4SQ#R^2NJ1IcKdF9VQI;Kd;I#>&2P6/gdRbX,a6>W[A58g36D#?a
VW9(C_(;I)bI]GTWTRV.NY0L<?cK>TX=6-L)JRB?+^a5=^LUP?MdBUDcIP9#]=b9
@fH1c?3&bX^NGNC+(],1HLX:80NKSM1)D:1c16c1#D<Q[(E)QPTOa>WMV]9ZbLDP
@=],&ZacZ,E2XgXU#N;DVB.42EYHec3VEW,MD0&>7^-M?KX)TE5/;7,RR4=SI)A\
dG41aWMTN=5]AED()cM#NU>BP9R@OP1cMC?QV^XX-O0OE=77[10]O:6H69YP?8L(
He)9feCCK93:Df;ZEI/;VS&L/K_f&0R[11Pcdb3@e(>6OZ(L\]\S;1PVC/b=,3a5
_I=H-]HaND,cO^HF.QSWQM-Q8OF030\fI:?a1d14?GER8^/W#9TJ@VN=U:Da\ED=
:7JMT97CZ.O>Z,7_b[^^Qg?8ON4UZX[JbYdeO+g&L=BI&c)/N+-abgDIZ1Q.X7AQ
(Y^71[c^0_?5@OO>5eb2CUc\g.9R:)_L;N5FQQX>4#=f,BH(@e78NBgaL-U_HEND
F^T//1dIGg+g(f1:7>M2f@GEI[O8D&AQd[-_/Kd:YX/RI<KHZXXfJGUQ6D.Nf/^G
D3N_O0RW\>,9YDdR-K8X5UJS364^4+?bOWcD@WK_3B<K+54EX68,+?G-Te[+Na>E
I[98bTFK-+dfgbDBY@N^C.(T@OP)KfcK1(gGBWT,CR;PX0L<f.dNKDd,AeQ^S31C
AIC/)[69d^J>&,b2f_[Xdf9L2&JJR\&BL1JO]UdAX(_38Q6@86@A.X&1]?g&:Z;c
0D55e3/RFUa.0Ce[PIW&9Lf?gM-U_OU1KY31UcDg58=UTXZE0LETa[)>YeadaD(f
V@Ha:]&7bN=;HYP_NJC0.(TS?&RDUV\&<FUS#/JCbcaXgMYCQTAge3?f:7b5,4D3
V4(D>&4dD4g^JH?9+5d1#G3BNZ,b]NM+K>E)8#+J^K68?ceBH52[bc^\7=I,NK@&
32MaPJ(J[1I7ALI/g1)H3IbH1T>_g+3O6Q/705IS]gb:ecDYKE2Qc(HM8BC9(64e
aUC-\^Ga&005gW/]PF?9,,B47aCABI&(7/g0@^EVM)5ReBJ(,W:b(dd/RC/6F?-L
7cXI+D-F<)01e[g/&7,UgHI-AZAOUO6QS6(W1LOWcFU9\2<(7_?LN80[PH2WY)(T
f9]c??>gZT1/N;-^5P)7fY+6,P&W#=A=eT4Hge16LeO1^#M:?NG^:TT,)O(I=]eQ
2)@a=VT[-0fLQMAeZ]HS)Mgc5IccXOUb8(;ea5^145f/N&:?.TK6e3S+OLH>E@:7
g##f,]EMWL]JE@8GVU1;#<8UI[.DVS^I_KEEETGeX3EXd[e&b4WFaV.1:_]>>9R-
dYIa&.B;e>+RTZ,FDUNO0IZ,-2Fa.Efb\dN/:\g4@.\093WKSY275^LU_B]F>D8@
/acS5#WROR]e[4SgL\>V.61(&_C^a-Ag57SRA5+K=feKZ?@0NeQaC<9-^7c1?Q=G
AO^?DGbJ#&deGI^@=cA?HS.8g84/[aY/@O;Y>D_G#V/N90<X,e\-M(/).[LN&QIH
a5^>U)FC#@@8_OVcdGJ&1cFd73a=9\=PWf3,[M^2Y>4eR9?HPAN,0V#;H<,XHT2c
^\Q,H&^Ab=^K:bP+TAcT)B4(TVLEBg3D<-7(AG_IO&c<)BaB#F1U;0c-L_<=6:<&
14<,OT)cfeNXQ^.b-?UH[RHJ9V?VX-4-]DME=/VWaCIbH-KaERd2B@8e3d&G9cbU
Ng[6-NT.MJ5#-#bDVUB>/8O27gLQ_P0A45cOgNa.ZFK+H5W>/[2dd#+3HAE:X[=(
C)0W[PZ;57&T0TED91DK-VeLIZB-S)gVB#Hf.VNaY@WQfbLMFVEbFQGZ=_(+LJ1N
QMOUg_B(TfH<V7QZ]d@XJ)W>ZCE4g7HS,)4^6A@Ba0MXCcX]=C+6;4T1#PRZ74WO
5_-&Y@&Y7LKQ^CMc)&.gP4WEGLPV<;Y.C8+-CD82_+.R]HdV8eS^J.081fP//?KE
\>B&RRegG<GJ?eT>;#9b/&Jg+gNfHAb8+YgDL88K:NCMH>g^\_IScZC^g7KVD<C7
Jb\4,SIXWN,DC.L+-.H6IY_MYaC+WHI2f>C9=P2/DHOX=#gd^bB^0\cffY:>.K_8
e)SC;3F8MXIDQ#-?(Q8#X8-e:)V5T\@(&G2M^3Ug0KE<)X+aEVRVD\_)a4DA]]<Y
ZU?7G#K,25[JG<F#K:UgcQ8gb)N/1ME7W<ZP2cd4KY7;+@#_]3:bd(eb&<C.\f(F
H#8b211ZEMICDEP,^@18\E_QEgW[G>d\:S]E>d)gVKb#]aHO43aeD&\2+Y=-d@(_
1QR,+X6[Zf=MP\6f\+6&(/TOGcg[NX_d=(Va26,dE9QJ>LM=5M(\:L_WAU?2:]4J
_AAPB2NTe3>.RVYQ,1/7NHOcSa>cTXdgV=E+TK>X;S#E^&T>ba:fM[P==;21&WM.
3)1YP5g7@SFMTRPI83D=Od,+,5J0B@_L8CO:WOdRR-OQK)L<Z(S<=I1d?MEeUX-I
F&:AD26Yec7ZC^GD+DJY25#Z2Ag3I5>#?17LNA-?X)OQ4O]8[g=5V=EZ?_=dGD1+
@g&5#F?.>3SQSOJgIae@7OXQ2BdP@L+=-MJK4)P,b^/f_BU(R06eb;=@&OLA98,,
V_UMT+97[UZ0_8NZE0NQ:6.Y4PU?BY9#6XaYR2+0-D+Y]ff?/;1K^f0\O@O_@^P6
4LX1.0/&SHDRCHATA.+8#JbG/8XO78PWUdZ84Y1(O\)BLAI\:^1+dDPK6DOTXQWK
)1^-J,fP1KEdA^g47P3LfDO?0[HDQ;3gW^@?^LbbBN<8TT&@EZLMTD\^)3B&Q<8R
[K5EM_;B_Z2ag>0FU[X<KJFFVNQ.))C:DY^bdZM8A=?S/1]C5#>JMXKLWGd2;c1\
VQ/Yf2D4WEDFf,XBTe&#]O#?U7F(?9PPR5J8\Yd[;2+DSB;aA6=B4D08EP_>RE(>
6O-g\^,,L#cHC#P/N;f;DM@5MW^V0^4ACaT9Eb[RR>8/<1a5JBUHI6<+,)P+gQ7;
3f#AdCKfSd(B=&gC.BMb:^TceT-S;fdP-@D)VVO_=7\bfK7=G).W:.V;?6,;cC;<
e?,E\)e,NN\CP<AMVNeC:\9+&(c+8+MbVPH_P;AOGe5C\+M36XFH<1&RV0RU3c?B
A1bJ1(dFXZebe2\V/C:X5T@+OMF.EP2TTU5;A6\J_\dP))37IaQYFPF?Sf0G[#[e
2R4/:fQPbS3047fZd=-QgTA([5YVL<cA\MGIUO7#.#?,4b.8eR,&P0(94.U/T#>8
S;EgUW_/6d8+HZe-2K[1/QC6=gIMH1SDT</cVP+V-gHT>9O.DfE=JR5AQ5UdMf#B
F&L2.]G4N5.3e(6^7,MDS:JZHW[.2=+XOc.EVR80-&bGHTQN&L/@7[);;#C#dXb.
,5-T6FLWgIb,f&@62O1LCDYb]#M@U:J:NDE:;JX5CRV[/[e9g<c9RP/[T<IO3/Te
1NDZ;^9X2()82QXL\ca\#YXW8R,C1a&IbQX#,<+D+\O^]KS>P[3/N+c7VbXGO:^&
Rg0XT=)VFS3QcS_SG15HM_=UPRF2RaQZU6>35:eH,7Sa=Z[U#e?0VTM=4N7)X80<
a;,@LY);0Ea^F0:8+W>)R9+acYF392[3)5QA<K_e?/+;7S+5\->#e7UbfbP1QN9D
\e;G@&V?VL(G_@NODOR;B+BID/KR<KG1D/>W\B2P7?6d7>V4A;aFDfQQbB)1+J+4
U&WS[=\gLg544ZD+5^_;=M/&(FHZ,:TQ6T2MSa1)NSM2baP0I=-BJ@f]UZ2#M.=@
9(V6_N]W-=2,>)WO\82>+Vb):OV2XX(.Y5A]Pbg,8G<L\MH&JM9FSKf;cPege@D<
IO76dDS:=B=2(#JBUWS^dWS6V+WGcdVT3+d+(_24VYL+:5V:ZSL?f:05IeE>3DbM
53QNMK^\Q0gSUKIb1U9fJV2ZQgLTPSHaTC@UX.^&&SPb6ITM<J;@C1<.HGfRB]])
:]&^N_)ZNE7Sb;dOBZ<&@;\c#GffD[D0/W2e9ALS@&Jd8)Xb(;UEdcB])L-Z90Cf
L5QMg&gg;4b_;^-R=K24efGSS^Vd&_#<G+IYgM&X>.5]O3];KcP7BM1bWdH\cS;E
S[Q4R.4-#5Re?:,U60Z@TTX;U_PE]S>HINN1c\Rf;#N;EPG:UddRe40N^<D1;XZ+
GKIRV/:QX_#FW2@T91?2f/G-/.6b;c1/Z.F7PQ&f:3;2/T6MA/fUKD]IaJ]gge/O
J0.J-3GPA/BDK/4)7G:.>L;K8<IYXM,LY#8]@-\9F[Ka+/Z4c4KNJ.XE^@1@9+WF
#dZH.[E>5TD4L[f][MfHc.dR32K?.XE9\THL>3T?+LE#]5D8=McbZ&aR^;]Vb6CU
L]GF#N0MT74)4JV?=3,@(>Y1a^O+1(6Q9VZ-1Q-)#B^eLXA(XJ^>I7Cc/@D],dDW
_7\;9YJgf;GP7>S^EY/S9df:V:-JN/?OE((GKANd,+(FfU3W42cZ;TSU,K:V7E72
,.OS)=>VR5.(#K39QOE/X8X>7^;_DHPEJPN,0MZeRSOR.D^;)TdP2c@UDC-L@^d.
@N[cc:+bL4c8+Me95NA#MUY]8.cTI)OI>e+F\>Kf_e0b_^4CI9G5&K;,/GFe<J#(
WF=WDR>AdAR+,bZV6\WN=30._=cZ6,Fed8Z?6S?aBDD3KB:Be8ODBB?1C[SWVf(8
Y7V-dPQ4bV/.I##Rc,MPQ=Wb@4?G9)#g+82<02)]][[-UMS[>5f8WN,ZR_7DK&\D
<2\257ECgN?16WZ[Y[X;Z/G2ABFSR)eU)0V^]8,2VSGcC00S=GW:[]5Q(^12;NNP
@bGSe+1#6LYbGH]EgLFH@CdT.R?BRg(FCF?K^UK7ede7SN3,7=c^D2FP&6c-:a)J
#K4XJ=5N8KBEQF/XZ<>>HZ)IXIK/73;LUNG#=5CS/([YY>7&f8S<1Hb?L3UfbAL@
#JP@)&.[e-#L:T]TA7g\:a30Vg9SMT[BIaKWB\\Y280KSK>MVNX;N.8ebZ0A3?IA
..T+/LC.Bf1L=a>6DMgb4Yc5gRd_Z90MJ:)P[NeP^?Fb8A(C+MeGGSV@6:aXXf,6
YH+8)JefFI?,aA\ab,gXQ(:IX]K+,Rd]D;^P>P=NbW?SJJN70_F?Z,/Z4+B#E=Wa
R5VgQ[).,DeO;5.I0)[4KeaV.OB:P?0HITd2CdX,=]0_,4/VB,(^)I=L+P60,a@g
Z;,F=9BO0cAXV31KC>>KHRZS5[20e5#d?T(:.11RS\+OY=X?=2Lc9,]gKM=F@?A.
]&,HDe=-7d=C.M#G_\+OQ1[FE:&[;HQR+IA&1gG(H+XW(?]<g[-TW4AY[\O:>8KA
6.?a+PRRPb2a2=eO1HXg9&6a9(3ceNC:#UWDS0&L]XV\VF1S&G&Ed=>cBR-+W@.+
Z\b11]2PgB:^KgB\bPE,V@ZKJBSaI-.93=]HMHR_4J;,5W)5\TU-4@KLY-RU10F+
=/06H0D3K3R9M\#a><SRG^eD[d^9\JcVY7/8E)f4WUCG=Qc_6gDP9#Ca&\^2d+4U
W&5?0B3N)X5>)aV?ac?&61B8P)b?fWWd)19\1:KbJ1(6;^YaNbT.(c/<VX5c8TY-
XIHGVB/8@J[^A8]b0YVaJ8(g[KPD?\.>-I2;fb5S=1bGK8PK=UODJ63UMYAQ>a5J
O@-GNGZf1_GPege_Md2KK@ZBA<7I?0V\6#_6@QC=c\14/Z?(M0?[SCMIR?N5.<GZ
f(E#39ZHBG?8-_]S0BAREPE=FF6BWN?MB(#_N6C,KO_M)7.8&Gg1gE9/B?fa6d=)
0NHeC.:3QGeZa,a;MF9R]75?6=Oa#ZD+?0b,dT>c;R@?,a.KPCS(ZJ\e/2,Z)G5E
FVe8EO.;F/RDdVeZLG)bK</#>W^)3AS5)^eTF76S13_7DdV3b3fcC0CT>c/=X1)W
?Dg]53[3Ief#P]bD8[Q2GM2dL<^b4X-+R>QKN)52Be13@&MD_FQ24UfaQ=E7TKag
9V^b.VdK2:409^7I7#-JIOB2g.8MTD7#WX)DGVF\D?6(PLW>g7T]f=KG:SG4R837
Xf);9>bEGO\V9cZ1KJ^IUL)5=aP7J=WWAI33ZS\I\BX/dMGFc@9,#UIZgKCZP>(7
OH;T68Gd:(&GbXW(.T:bYbT_0(U:T]EH[@0+=>^aK&,M)@7-\R5GO>/9-?E8gOTO
KcC&aW)M)VH4cF.>XcU8gJ^b6<c/QL<b]:E9(aA9J80(YW=3[W:e+0/)J_;Y@1)R
6aCc7Zc]NRWQN48-GYB\.0LN/3>HG6_a(F9cII>eS,U5UJ1Vf6]/F(&WN8/6b0@?
<AC=S^^CDU.R0GPSCS.E8F\62f-NOS]aM2U/ZX<ce6S;-@8d@d?IGc?#8X\IYMF&
bQR.c+IT0[-X[L5I>OVK/<R)A6]]PB0(3)@?K+Fa34E_E:N08X72_5dENVX)Td7L
PZ1ZCCO1;D@,^33]843+W4YE=T>e/MI\.G=/-Q\@>R]KP53K4=?,.eD[Z/<&(XH6
GV?-.YKcR5Yb866c?:0OA8PZ5/a<c<D&J5)+X,)2S27W@0TZ,gKGa:<<_JKCC#)S
).cRX-993@gFEPA=CM[c;XTSN#Pb/4\(cV:3W4[=;MYXcaT@f)U0VR[:e3^BF_M3
5K,.3)S[ZeJ,W(Y\g[(HC#URH3Q:4/CAPEfM?1J06&BHEf6I(IT/5;Q#^6TS7Q_b
LA=ELK6^6[C]?6L@V?(-S1MZg5C2K,d>+UTMQ9;g.7?E2Ob>,^EE,TR=F11Ea6La
#W.I<;/e;/f3;@9gT[RUY9fe4UD2<N/a\_2\/.XOeY1K[^2SSVdD1aHW^-Z/C7G&
:O.71e-AQRPf@R3S(b465W#M6V]c=0XPX+/bQ+<FY44Nd/7WFEPS)(be40a_OR;d
FNJ0R(fCf:1S<X,J;VNEUIa(@-/LOOdaT]0DO.V_I<R8V_LYEOM<K\87YFVF0D.5
.S(KRUS);cU(\ZT1#O:BD&1=_SXb]^Y?3Gf7_[Vd2Y(@-Db=&ECR1gB_R0CONdYd
NI2GHNcW)P/>(]aD]7+L8-5-UJB;^\YKF8QKN+eBQcCB)?:KJKUg<.LQ98E.HQU?
&K8+D0@:C]QK\G&5Yc3N04W8aJH?T>6D2B]NYD2=/[RW27H6Uf==\6PCDTX7Pg>,
N]JZ8F]a(S4M(@C>^BY]A[[C(Ud8XP_[/UaPV#f&dGT5_2;3SGAS2)9VY#X#7)([
;d0084QAN]GF2;^X(CdVgZV8XfSI:5E?0d[+<bI9b=NKF)@DT\WgA-MQZN<0]HZD
<@EfEd-[=9;f.D<JbCW:^3:fEKg+.0=d6T1(Ccc82NFNYTcDb\(P0^N0H?(:8gdb
-LAS=J2c_]d0>V<+N##[J@;4cKZ9AE)dWbd#X3W7(@?UWYRCIUXH\^M=PL[Y+6]<
3&YOURT;8TO@dO;LLR.=NZe&d^f2R<M]2A<+<SUWZfd).E&LfgE&H(DHNL/9TLO<
)Ygc;edA^C;2aSCc71#)8K2LZWTbB200/Yd(8.WBN-gHCg@Z0>Z5U:_)IBH5ZSd-
/GSFP;U][+FS&0^<Ma;OE6DR#9(D+@@?U_Dg#_MOcJdKCN2f(AD)f:G;dFXaa/bL
P>Lf32CB=_QFOG<IXO5;b][J[M>]+IR94W&Vc+e?>NPd,>+SK;cHS^gG\:6KY4de
W78CWbQcWg_]ede-_RCOe/W6=UFSO&N#YH<B820SS+\<2D_5\)-C=S,9]J^OIGJM
0Hf&5L=>a3EZ2a>&QcKPLJE:Ff1P/R)<1b7=Z?ggY=bOeP?5eBSB#V<VeF(+?\54
gb,,+F_K#=Tf#;dNaU#)F1&e;W3=f6L1T>e<[705Qf/Y3?#K97]7b7\PgFB:JE58
A88fcT]49c<66I]?.6-_<#RQ:9;N5GS>;A1YLf?OP</3a>V6=aT5@0Z-D<)a,0fb
Ce2EVM]9^1N:8JfDLGF7_UNGJDbc(Nc.6JJV2K_SC^>:^5R(S)fU[+O/-G9EOINM
N@-dMg1MINR;b-OV;#L=,<I4KCg2V^_2b(<Hc>EVE44G>1QQO@1bWfFM(FS]3+Kf
GaUGPB..WQ^bH#^:[g86cdg[aaE23Q-;OGT:_Z,,IH&1N;P(B+c0]\Cg4DOf&>QK
Z\G2@LO&@2\cT@172Ob\_26GbZG?S1)(C+F]#@UF;+P_f&B8H.;C:T&bC\=SZ4\4
ZCY9:ATL==9IEAJ_NBT?dPUA2.F:5^@gN<-34C9X6^c=#@UA6N67.+^7O97RU;ce
OU04fEeK\8Y@CV0(_<]g<a^W[^CSTBOP.KY@4/VFFO#K:aBL\,7>>2L,,<]Z2P;.
.Hdb.gdL>VHb@Y5M93<YP?^FZfIXW[X3@LY?L\BE]-VfF82]:OWH::Tb-P]WQ0DK
1fP=)3S@eB_MD0d(P4[F8Q,WeL@WK>2f8g.-3/bV7c/P1Q2UcDX\C_J,&&5OO,UO
V=6dT##&OaLd.O,X5K71(SSF?_Q4EVf/SV1a&-LG]Ef-f:O+b6d6:cSgF-JI,>B/
[_5JV3V+g6:N0f_0fe):MP:_BR<?J0^LQCK&#3c4QF-)+(E>6.SOX&-QcAB=2A:(
;;KMXEDgN9/IN]2=OO]\^Wd@K>=,KU6?/N#)fIK1/#\[Z6\70KI5a8US3-[AC02]
5Q7^2?e22A;B(;A@aQGbS=7d&UH.R(TVY<=5L792>).-XdR;NF.J\K5f0]#N@#bW
g<:083fB=7^]SC07EY[d(b9d6KIN#H_S2TgDR,P^fP4^N;4aa:#5]:XHL7VN;M6V
Gc+B)fY+7S/)AE5?)DZK21(;ADQTY\\R;DMA=/XLgS\]UD<O2OFZ/36@M1LJ@>,Q
V_/OdZ&N7eaDQ-N\N9#)[LdJPdcWa(&V5]04URCJ#3N3_2]eMd:gFKbaGQ-eTL9E
CX112-67)AB\Pf/SZVU]^6QHdK40=5f?W4+/R&\gS34ed#?acH@e,),a[ZBT_RSU
,d4O/BfaR_R>XX,BI0XV<[9(;4+JK2@GHg\1AeD_,<KW)b.ZOT?bL^+AD\&U0S)[
7H7D4.0I&gHb4(K+ZC;E,@FL:&()Y=CUJ<W1/)C,)94&KS33M3HfV<D7W1A;22W1
TZJD2e?NWc_8/QP9g_&fIA3MXZVNUBAd[XT/<AY<Sb5=#FGABDgL3G1#[\J<9EJ.
RB5FUg@&McAGX^L=.R>GM>f&<RXX6BR>HD;>=La+^WO0.GP+c0eHMdQ+I.@R@(#2
JKY5d#GBTD)D=)7K#/[?,=>>De@GSEOO>1,UbUc\T1,>H[6I]ISa+8RM2X=_e\c9
MKY@:B^N+cAgFNCN@a\>2;S1B3UD+OH1V69L0AJJJT]&N4-bcDA<X^)>W^:b^dK8
=M#<VZY:;.6b_5O&@E/)XM3N_cRW0U?0&S)2,FWeX>6F;8;bBH\GWZHdV_6_P6,+
3BB)6G\KK?bQJ8dcae1+=PKN#Fe=P,LOG^L(1[L9HQbLDdCA28WfF6,VL7)Y3C\-
c7Oc\?OX^+02eAO_&OPbVN\CUa51R8[L7L@NTBA08E^^AZ2gKL)1)A]d^&VW8aa2
YQ5E/CX4D<_YPac:3@Oc<3;:2gB2_M^PIAW\SD4<X.[#dSJ0f5@^NdeeK7V#PBV:
3?LUH#<63M[2KLfH[[g?B]&IH]??VEWHRS2GJF;Xf##+2IY3eIAc+3>T(JZ(?1?[
:F-5<=TPgLP=MZTUe>-+1b5<:;;RL:TRaIQ>e(dL^S-PD;9:64LHWAUJ83CJHP+9
5A#=G2.g6A>F#[#a4P68M67eJ>0Pe#>,?0^0QW:1HXCa(1&7TN&T@ZO09@ADTbPY
V):L:bFb05=)T:=GeeAQNR?;I[\8=Q<?2G0\eUbgeQPBe4^5:ZT:ANTO/(ND-VNC
QV#1/HWWF(QA8LdKP=IXS6@ef<.HM.X6EQg:Z6LLY58(eK7.feJW.T[EYZQ\M\W\
CbYKWgRISB&M+Oaf(K?NH78:&+(IBUD[?25b,3N<SWC3M,T\YW8LR(_ab1D+ZKCK
H\[,F:-^(8bFF4PH[a5P0fQWN^:RHfD-ZFQddGP.T1Q0VJY#GLM;R:AR(O^)5L>8
aPI,0KaTcNN4Y_(PF?G,.M,[ba]J6f(d54,7GRffUD7e(EHe9^R>RXFD(=d-bPM2
XH3aFT(/DHfeKTQ?R3?7?,6^bOJUb:Xb6H1#2/=2.Q[(/_/\=XB#<<H\6b5UGgEF
VJM?Z?F:g>75]CQ8FF#IPLfQ(J1E13:F.?_Y2d#6]L[P:&F_0_4.QMe&M2H5Q<;g
BTWUG?U.)H2e.8#IbAe<DA<M?bfWG1OJ=DgABXGL(OJc>1<.:3XP][VYd;F&K]CC
>c@UP3405C\8#,JaEFa_[]+_0BfLA\_DO&S#_bHf?SVGg-G=,BeP5cD(:[#-;.8#
J88;&1;OQdJ,[(RMH@WW[WD09@c@/=<=ebE2HScV)Z(.EJUBS,@\&DN<SO(/GP)@
76YH.VX?2Ef6Fe/cOTDeH/ZQ=4<aJda-eUV7VJSP9Af-NeQQF,ZH]?FMN,^F6N@a
7K>^aZ&6JdGA@[dHQL\e>FC1L3E>SK@@KDU@PGVFMYB]&A2cFH[2\c8A8OMVaKN&
X(H=c1RY?RR-W/;)^:VE/bG[/_<)5<^MD99\_P2E;GPD#Q2B>AY9/UaPg;)7?I>g
1cYD;_]>NU:>3eI&R]3TP\^;F>83(#\DE:S@R/9fbU5C._LRLD.]E/d&]]RTYV#.
0XW9@a.3bcB;6LNaV)#_a=FU#(^?6((@5J\I(IPQLDS5XM9W#D9]I@97;5:&D5e\
F>-P_2M.R)A.G/d[X,DZP+(,?g:=(-+F#C^D[(^eD\a8Se<-H8[^JTWZIN@7:^+Y
#B/2_T^a_9_99?1aJ>ZV9dc7F[E1=AcRPU^O+Z0#HQ0S3,[:VIcWEBV>ObAGP\<7
RFC[^9fKSM8H/6JUN.148M0)+)/Hab>7^81?3;NBMR#FdNNbGbF8;\;Vf84f>c4H
Y,7E;J6eKHVSQK9W&<e>8UN#Ya=TN/^:f[,W\W)(?f5H#@I]K]P47#.g4:2@U(Vf
dd_\\KU>)2-^AT:4a5>?[I)19cLY5TH8LFK+Y[cK^7b3&B,0cfQ<,8=&RTFSfW4Z
feKEg9g^HKB,CY^;6.>E]8>ZaC#]adaG)3GY_S])9#F9Rc_C;+1c=&2V[^_UcQ=J
\Da3N,,#a2K>;@UbT.B3Y<cd038/?7\Z.7</AS&T.f1e>MNM;Z[:6+7dYffWb)1;
.a5=LPU8ed?g)ZGgM2#3&0/ZS(XU;QPX7KX(,dH;U].4Q;IFEOaB1>@^<0^#O/8=
LeMS?<B7Cc\T.TRU1KDeV-E7;XO^@WL1aH4^]]2c?=V7fbR;5Bb]]cZ/BLUK)bEg
^X1[??\;22<-]JAQ/#MOcZ7W4Ke4c>1M#U(GN=4>ZOZ?DOf#e/,]WT]Sd495fDB)
BH_\ceEg7cVU)MQFERQT/9^S3c^DYAfO\Y#07#aY(b1-g?;.RT9ZW>C_J@Y(G,,Y
\c2Nc6#:\\6X<VeUV#ec7#I&?N8C>g\?2b5FMT-UHWJ?)@LPNBC><:[+J\F:1[0<
B2N&,H^JcOA#\)UPKQWG47]E968R3g-8JE/RJEV(;T.,AX9[D>3PFVdf+d,O][9f
IF,TcDPB-FX[BW[bCcSW<S.L6M_=Tg1TOP@P4.dPf]+,7+b-MgMXc=6L&5FFg<5Z
5b(O^JPK[-BE/R4?]C3eg\2#J-C@/.aEF0R@LaR#MV=AWOTXQS2IP_>T?ILDO^&-
MA-]aCK_?LTBfb#:<(.QLXY.1CNH/\=L^_R6-\5dYZTPEW2^a+I>Sa7Y#dLXU&cX
7O;(eEQee&:WL1PY?:HBAV6O2Y2(KMaZ6)O]I,,XZA?.PX\(3@^IGWcGM0DQ,B?2
e0S#]c@fGS3fLK7=I,eZ8Kf/G7Gg1H\USPe.3E-5H#-7N>MdR\+3KU4(LAK2f;=@
\9M9QEVF_T[a.]??+UYB,+b=^\@EN+bfaQWN2H]A,e^a>N=VVL,aUf\97FDWQ:EC
LJ4S/_F-<Ccb4/UELJ?Ve@Jb,;4c9/+V_(3AQC:6HE>^#3RTJ^=Y2FZ[d_1>&TE+
NATQ:M0;^&ea.DI,8AZ:/79\_Y[,dVH\:ZO(F=:7e,G/B3@/[TFE9R[4NYF9>EUK
.Y52.7IPF<Rd#:9#SF:GHO>5R9:_N1\1@^RX>@E@PS?:HL/Y?D&;90NJ2g-DZK7U
ebg[:<F3Kg1<N@P1G-;9]2D5NNFKG#_40I/9>AVM(98+J:CbA/P@XQb3N,_(I4OM
9C=>;F4](D0+T?Me7R2G>bEJU#?W<P:,RXB<E7D>)3ZB==F4#94D15\O?,C5QMR8
]:=LUM&R_2VI^KLD9H;F[\-DgYc[e.;GJ/f8JD@Sd@eV8LV(<6@@JYfd2d0M<d#K
V0T7ZW+?O8LLYQVIW=<;P5(3UA?LV@GP;+_YbTHYO>K<.6U]P:TJN#&#G.&\B;UO
-SD@::8G^Q<g+2e#]<:6DT=?;(Wg04CfAC?LZERQN>V_6@.[=;R_?aEJH3./^T=&
8_C0J&c?J(V38cHNGE7[\1KPIEXc0aS3<4g,GL-QB=JR>B#J7QVT5V#([.[_1If0
C)D;/96W5Dd:FT92WW-gDO)A[DEf;0CYTLO.)?^7<4Q_02Y_IK(37&<</RF2TT1W
[>CVc>LHLY1\_#\(<5^f;B1GJKL4W<X.-+UEdH::<RAF.:A3(5ANP>LV@8&@dD^7
MHN9N#1UNE[^5N&#P7a2f@O>[+?BDT.7beACPB0.2V7^OE>QCQX.<(.?Q,K30#a:
V4J)B_Oc7907FFY@&WJV0.GM#/dR:d7A^;WB.2([a^AAbeJQFdDVY-eN7[-2OF3e
1GI:I/+=R9/D.FL[;9GI#_@eR>)>P^F)X9K.I<23]6ZRIMCLVS1YO,UcE(V6Qb+K
/X+.V:aILa85PV[67gPYUP&FgJ<A2EV1+K,D41O#@:]5VLSX@+D,&=CWW<c@a0B3
2e0fEGGf<,#1EA(2W,@QU2I7SCVA59(a,B@^HTZ&?dF+8]0N^1S=5GZFU9[GHYXH
2DLY,GMEITM][Z7#_,=M56)L(BOCSEW)RP0Y5Q?E(4dA)K]>OK&A\cX^Qef:_gI/
@VN[I0WG77SG&,11]d<1Fc>N^ZO.g@2E]YV(_ZG?1X_TF5dfaf+>Te-#@#):J.AL
,D0HH<?8+EYZ^8(fT3e:O9:P:<>O:I6WND9W<@.NMYCKQ,L\KDPd408Rb2B?NR\c
#/<;6bRV_/_I7V]_)#bS6f(a&RFA\TKOPL\E+]O6f-#:+PGQU;gWE,E)@a2I<,:H
_:;:GBGdS:YP6:U5HP,;+5C:YB/b8AYQ=_9YgWf/<-R4eg/(@/1[6FIYAUYLEP@4
\ODfd#0[/@g_S,XM#E&,[)SKW.SG&_5#V_T,[4Z[##B>9U-12G\P8.gOQHS//C6f
1>4H.1Re?OFBVL]9E1J@TI3T:UIHgZR+N-aIX&dA@b)aIfH>B(:&><,?R@HF,;V0
eJQZ<MUKc&?184C#SES#ed64-3PdPRUfG?B]&6KX#IOX4CQO=e-2<W5SAdde-J.:
R4(?(LbM<S9]FM7\A2Rf=+FZR:+G.AE(Q5GBB18]dBd[TXJe;0ZFL::Mf4S=644J
)]<<DNZc-9[^;6E;SE6eN#eCRCZV)fW-<Ha.PPI<;OP6HX>W6Z>-a_Ce;=1bS5^J
S0]ER>2.+_Pc:aF&@1a.=M>I-cYC0W,8=:W-ZY<CaV5:?XOI3[ETZZ=UbL<-773f
4)/DNPAR=)eK&D;A9.:93B2S_R^,cH>c:<M.a957I<g[\f/-aaFE4/-IMMRAKZ.8
/D.E>QQX>KV9R68T=cgV]C3eE/b(gfI;WC_36+41V?X\8A(Ve<#GQc9LC)fH(=6Z
0C1aPMLXNFS1M&GSA7WL.M6=UJPSV:79-.N7<#UeZ&Xeg1[_VUB<1#AR(19g?=10
9c/,F?#.@1_c=dQ_B)0V5?/Wf5VARS5XcbAB6&^\.ZPfPMd=7A3gE@WdM6gX_^JR
BaXa0XA-&^5_M8aLgZ1P,22<5Fc0fKU=OR;]VM_YEU-7e7/^]Hg6N>)9MN5-g_3)
Q@LeWRGRbUF[H6BM=f--8FN<K)FMde0QAY3gd+9Kg-cNZ-^G\SRf_BB:aGEF^H[#
6?0DNa1b9XSFg4)RXgU-7-.>174V>UN=ba18.)S-gDa6Nb?SIdH1789KOTV(P0EB
N=I;G>+CWd@_bERR1>\HNOENJMfEEA1.Q^F.aIgZ5_=f56dM/-F^8F6CEU-5IYeR
(N>9\4-BUZ3)0QK=.>FcgE)a[HU4IQ/<.&_F:7O&X4@,0bH\>?L]6G)0=B+@,K@J
CMa0S[ZK9D[PMKfF_&bTB1cQN9464RJgE&83S+&QTOOPH56QEPXaVIYIcS6^?)6+
]W_d#\OJD_0,U2?9M-AIBJ,#6YgGBZ4=T;<=UFI0NV3aGc-@Mg7W9Hb:18+J?b6I
N96>/:;W6a),N=Z&1.E]c[8O5/-g+ZBW&Q.Ef\\a2NFb#]9fHZ4[d,.&D2NFTO(7
_T27gbPa2g_7>QAN?H[J+eQ<DHELc+PE-\=R],KUf.5G:J<+2K?fR[Z>]2c3c=)7
2X))\Y6:C9I:RW#/@(:9:WEb@TF?\X9XV7Y0d:O)6D;[L+&A>f4@b:K#4N2^Q=cd
BHY]TLZbU+]g>R.,7cSKaC5d6T84fcA1H#^Y#G59NVLRC9^VA#/N2/7T=^Z,g;DE
aOg^fCKH.J3P<Bcf6XQ5e3(RgQ#@BK5/:;BYCBQAUY:bK8ed8/X:8\15ZAP[cKO[
BEU&3@d3a^^A+DI)@:@5TV7.-<&FK(V(:7S<LR2(Z5)?_VReD4)P=H[USQ&^]0d[
_@X)\S6#8<6dZ/Q^cX[OL:H\d5g\2:_G_cD9(0P]/6c\D&6U5RU0UEXcd3CTBL&/
G>9B0/Y+G=]>dE-CFRfF,7Xg/U7?5.,?L4^&dcVK>5_NEU=JO,#5A:>DA9@ZbYU,
7LTe5Pa.5,BIL3FB#@I:BU^ZTd7eKf,>1K7gXYPP_\F<.FE(<UKB3(,_D-8^951]
.g0RR&?c5.HB;fbNQ_;Cb__8C4TAUJ0Q])5FUg#I4Y42=:[aRVa\)?(DN+#gFE2e
4LP@+<.5(0&M68PEX1.XEBBPG+gW9dWcA4(].-S9GJ(H.OOF-5gXg_]XXLIMdW8\
bFI@SG1D5R96L?>XWCf<0^PO^925J-d5/TLN@K-F]0>/A7S_CVcQ)\^c3\O0=6M]
H+I1<GT(,c+a1TA2[Qba/^&NCI)B>Z?HC</7C?\4]2B_,A;3QPF3G.N,XPbXE\1Q
TDX_IKY1.E[/SCa,<Z7+TbWACHgEV07gd1YMVafe^+0d&G6d9QB46X2&AD#W1]TC
@.(N,I1DNX>g/KJ:eE0M9gRgLBRL;E7)3(XF/FbB-1,-7Q5E27&C>[c-0U;<,MVB
gBP_d3RaEVaf[+DaKK#+d5U8fGW<]dUP-G5:5>3#b9.<UCBTZW>@N5R_&7d?NEC;
<a1,7KeVgWX6b<@^gf=_Z20RI2\;+bAVSYJadBd?Ca>NSC_Ie+Ga<Y<&a4Q=3(;Y
;;Lg>VZ&>1]\K=Z_ZUZb0+EEf\^AV6DeW&AB\=8(39^-YRBBD9CWUd^._)3_0V<;
+@0O5#3?]0ae(8?P4b4RMgNcX19bcL-6RTf&&B&ALJ);Y8=V[f<IY;.?]Y7,e\<c
_:cV[;&9cM#/-MF_Ra?]]?IM5eILGI&0Sa\H2?W]>SG<NQJ@2L]A_M4LXVWCQ.?O
??@XZ90FM,G:Xc=+;)F8#@DE50VK^(\LU#8G+(c1VW#.PVE+Q^D/^>EYM&S::^1D
U6+-E:LZ<LJVa)R>@Y1D#,XQHcQG?LD_f0+CZ,QcJB0f3TI#g38H[-B8_2.ca/Ab
d.;@0A=Q&]/9RSJfJIVMH#E7Tb[;IUB-KAFD[H,AaCAaBK9cV00WRTeJM=f+LPgB
f(LMN#G3V=+EG?=1\N+G6(,Z([,IVP4^.46=#W2Z2^=-fD(#;VBVcW2Z:K#1_JFZ
=B>DRe6^7cNA)>]]-I&daSfD\\SOCSF1#.+@Rg8:U9>TYgg+_,V:^.0MO?(B8BCg
&,KTM,:Y/ee#8Jff\R=??V]8e\B7ER-^.gd)#6:g4eaSK^>I[1P9eMDV.24c.^-f
6,<\Tf_,eZ,fY_[UfZe<ZO80ZO4g0)gT&aX)<)/QI9/-.4cY+?JP3P./(K7NL;,T
Y:03DZFS1GCO2]E9(c7]]?e(d^aP(^g-IQW4G=@49OO-RZ-0:\R&:e0YP_NABM+\
WePcLLOdL7/J3NUV\B5+@J3M<[/a19L(UBFHYK?)FdFLW<Z3RARSV5Kg8EHcL[4O
F,DJc;08@SMZIDKLX[6.2Nf:ZaBRZSD-F\#E+3ddU.,/?;U[KW_0ZBU1EM2(EY,7
N?Oc_P9[M6C3YNa;a-G?@+L)RZE\]B(;GNed?VCO0OYcD?M>GBb?)/=R&A4YGXI:
M][^@3bYZJ_cg+VgeRYJDdF==Sg4_(DJX?JEP>ZMK&F\@2&=YXVe>G(_HLYa4Va9
S\A1.+B?A&ab#.Q3c<[W?O^07+X<X:L5)336E[N4Dg[1G>4T]e[-]69>4HP+/,Rg
T_L\[SNT7f&-HE5TNG:K98L)B?)W6E;WU9XUCbeD]]@^8DT.d<;A0e0T+^>4BLgF
;.?S?c#]R&PC@BI/HONX(?+d<(A4\C?\KN<GYM&\\K>&27-K39R(&IA#0>3-BXJ+
7Dd)5\@K+9DC##Q)/Fc8)U<F5I9]57dG=]@_<4)?ACW.)EBAa]JNYeM8aUcHP:)5
@Q=Lb+3Hd9bCbTX>RT9LfDcgE@](E;<N0RY@d([]dPGg5<D/g8(@O&OPVVL4AITM
1N0V+DaJ5bV2W.gV>12\@??N:cGafJ@/eHC?@5=Y@LI1ZL7^c9#NXGbcY/c5KM)P
>_&N2L^SREJDOFa:ASf=U/U\1H..F48GDPN=2M(9KL:QM?Ke503CZQ)MU&gb2_#>
(=E>CHPZW/0[&W)ZYe]F?Cb6B1RSI62W[^4U9Y&HCJA2Q1:Ib/N^PcfWJ_T2ON]>
A.<X78@QEd:.\]DV:(g@Aa@M22I?9QI+?9U3^R1>+2+:dOg?U=8GTLK>;R:+P.Z3
<?eW_(UadJE7gNb;4MRWQaC&JbLFKegR?(_KP(VV:eB/V;54O\(=M0+M6U8-05OU
5W0<LOg/0AL@8S856E0S(#Ib8Xg:eOK9Zc:Q06FA)S(Qdc+LDD0)?#?;_20GcT[F
Aa_1Zc&&b+=SG)DgO4:^f502@#=XgC<a#6>NL1QCNG2@dJ4_ML?P.NNM+b9=R27=
P1+LZY5[<(]C8ea-GfY8OZb>-6d@)<ZfGGWG5#B>XIDJ]Deg28O;>4ZId@A0IB34
:SOW7QG[d0Q?XPUD&>@/T,e+-aXgbJO=e_VA\11EUdJY<2+V8[;>Z6@<]Tg(:Z(;
;.FR_1KRgM)U4@O1Kb&ba#5-(L.4V54RL,O2>5Sf_dN?g001=9U4U3ZCZc.(@<H?
[;I:HK4+?47O/D/,:Z\U^&Xe8/FS58_ZAe[,Z2C4#\Sa#,^V-MA[(MSPO<AB;KI[
2-6<1?>F\85^(I.C>T6^_fZbZVFWSG))D>I0ZL=I4(:c2eaX&II#&PfbS1N=.P(]
/=>?=1Q1d#V.GJP=Z,DBFgEM++2]FITG8]AR<a\YQUIc=(;(;__eAJE]\@?K:^6K
X_H88QYdE.PEb4_N)G<\\ZgG86H]DCEe],724>G2dbK>Z31fA#V(2QNfKJ6SWLQg
aOO#)L]\^I6&b_D8gP/VZQb_(7<gY&=G\WMR5)0]D4]bWTX.-KZWU<1NT63d:0(0
QGCNa&<WL]d:ffe[:B@D;<4_2.TJ0.64;X]gNW4/PAPEg<88:d2468_d35@[cGDI
O;PC2E,dJ&C2GJ29S[Og,__#V]H9N_CCHV5\PKXVdV;]E15?4TCB8fR[.2[IbQZG
)HOKDS7)(V@3T4?9OYW./-,IQea^N#N(M_KC59T+:_)/LB.QCZ+9LM/)0Wef-bEG
Q.#]>P)18?G@PS26A^?]U>V&<Z7Y3M^M,a,GF5&XIcSE3\CJVHaFP[f=gD,54XeT
EQH#J3?dN-3R83Tb]5+Z<RVUF3WKB:cSVb-(d.ZG[TMQF;eCR((JKWE9>=_DZI.^
^Z_4A:QPQa._<&g5[?AFUW/8T7I</>XBLOd@&]L>\/6BY(ZG41b;XH^Bb@f(W4YN
CUc_7H(JG?NF(eD+.@)98AfVU-1a-VUIb1.aC7]>gSW1\be/>7bI3;Y>)R((.71J
+S622d)<-;1N7C+T,H)C5)[HL=KU5,N6AYg5,^5/Y;6]RF]W9PN&FL?X-#[]8Q9=
M;B:-]_3T(]/-LETGD^&-Z:U=0c27T6a9dHE-S1]]L-dg800S-d6)MJ,AXdb9AVE
MVP6ASe8@5b2Z9T?N\(V(X<6Q6DV2.(#?9O#>#M3NNL^3-Y<,6=eRL#TagYINB]A
NAc11bGTUd8QUYZN@68^0c(d&SPO)cILfX\X(R(+=A:4GU4W.2gZcF3I-H[69-7K
>eRd>OW9(RX5\cQJ]ZQe#9fa\>B)-Y&?Gb2E.X^DLY^:9;OXYSIY++8T<Q[;?b._
d.<1,bF<6PdMVZd:<;^bOT,_W@N_ead.Yc]b+1<+3=Eb?_ef+.)N/&.cS6DSdIQ+
J6-B_5\>>MP](b4LF3ID)/6@IXEZ^2(-?DSQFeOd.)gSW9:2-S,&QO+2Vb7S?K+7
66eX#9N=_[X8GHI4Sd8@OF@[N8H/UcF;S/1L-N(J.QZ(\@4>C=AbWGEFdb0P\[XQ
c;a4FdYW?OM/d.2[e\c<OF:>50GRL&2\OB^-/0CHL\:,HV#=>_=<X4B<gS41RBfT
,G:W9=g4VTec#2dW,gX46D0Z88JHVX>,(LV&]-UCNDTP)eM>6e^)TcVO7KE47\R1
HEO=Q?[;MPd1=4AQ:IAaaccD_=)/[La+H=WDQK9V:R3<O8W6_eL2KcI:R@LGN-R8
]L_BDO5Xf7-&b33dI7;2UGgX1M-IG,XbdS;:>T4F,#bVMX-M=I/ZRNgUCI8b+.Se
0N2WE1^\\7A&5XRV<95-CBeCN^973EA<><b>H+Pd.9ff;&0,/A983Xb<PW+bCE2V
9M3WMLDF?KAR]H?;?Cf6[QP(?I7T@FYbFJCe7T+4MB@OA3CWHKd/;N?S-FC42\cA
(.2V)6P],GUT^Ec8dBB(S?P0)I:b?c\;b.+M:>7b-.S/adQA[aLOH0UV?R[\8Zd3
CB.<5b],_(0gK[KAI>H:(4J[U(\^BVK/aQAG9VYV:9ZB4fF=#;)?(AYa?/[7LHOF
YeZDM.Wg1D<1V@8\KJ-gg\J1RDY(A8CW:V^[Hb,3&8c#;,Cg3XfIQLNPZXWA.=bG
@7GJ[684IO-V/XMK=YXW50+4?fWUTIUHN6YHXTW@57S=S;6^;<.Q>1SLC&a3]<]Q
b/15/LH?GUd/<H:(.SS.7M:XB<H1Q6EQf_,BK#B_f?-\K+_MP_=J94e0g=fSD+Se
a88+X9a)@J<0c3MI0M2AFRR#c,f]3FZc)cA#@2<g7dDV=&&NQ=P64Ne:fa92dXgD
4E-U3?PRL>H:,=8(EcGL&d(<.V^=[PVV=>#Za+O:IX.ff9Ib555cZG#FS\3\=T8G
J,#/T#Q=6XOI1]5@>>RYMD0f#\&X=5B?QN3NRCR],IHcX^MUMD6eK4>\A/<LH_-/
ZLFeM4MaN1)#U)c5=B1agb@I>6]f]Ze6OKdR)VNY.^+&]W+SNJE.QDT_H87U4f6C
be6T14EV7[^:#I5DT_^WM3\bEXad9d=&A#fNF<:SXVY^?;@,7CC#1AB^([@?#JH3
<[.eOW,aB)Z(;a)/OJM6X+-8S_7A&GJXMaCTRH#TA^QHYg6OXV?><EbZ3.FR7T4-
SVF.c&Q.ZU=T:V5;K>4J9DaAF<Q@WaUFdgJg1>8\\C?6<[:NCL//X1d=/_[##=F=
DcGacQH:L)OM,0cSSI<LUK_;eEB>O-IGR#XEF2]N=)]WPK;2D1^^O;b,#DJVGV>a
U-5O\YV99ECK6MTLH^29Yb@X/Ka5.Rb>(-[4@PgPFgNIMS0aa;?=Ca4/gI_g+IO6
7(ff2(ZWE-b0:PeL]QdS@]_Wa;S?F<MTT=/R(5)8=<LX/:VT0CTdQf;Y3ZM(-5PU
eC@gM2@_c^&>@_B00HXTLV/7^0Zbf260;VgSbJg2L?HIIV;-a30TE8RV8\<3Lg,Z
c\5D+[C9H(60eXF:5NRI0I?QbTSR-K@=gcO3&afe9<0:Y&GI^(RW+)Z?;JS6c/M]
YW8;@L5ZYHT0.WMV,5U?^VJ&BA]?7FM7R3-I.03X:Z\KKM]:)P3-E@I#R4_\Z@/_
V47U18319Q2^BI3eGPR5M&)84GT45Q7^d5;DObN&6^OfXH)IgA=<TUXK#T5_Af>]
NQ_K<<8&98Z]@\DI[c(O)b^Xd;_4)6_S]YXNR9IdY#Q6.)f>#DAe+B6XFBM]ZBb7
]=L1VbTN+G\],&c^cN2>66fe?b2QND7-3YOOeQBfBER^97&>9,?8WaAY=@LMK(dS
gD=X2]3ZEA7L<Qb\GP+9cRW]9MWH+RC?R7+H6;2.gW9eaCNJ7T(4GBcRMOCC48fA
8T=c&F7=O:=19/D.82cDF5=):Q&8_c75=2(?DfE8WYL7\.3bcEeO[@#RGb/FXc<V
:a4JD)F1db-S46E-Hb=-R_AQ)G](8;ZX[b;@^b>:.6&K^CHL&SOJ_gSeJ=(TZRJ^
DKf+):aaaPCV(ZRRT/4aWU^\R5PSPGB)YP<V]5U9ZC^#RR>aKB7P\E]Xb(HV3f=E
XM?C<12Z?1I\B_LJ(41L.K>HRX(:HecL/;E^6a9KHGg43T)aVaD1LfVJ_44-b+3Q
abYWX>D?):751D_?,FS=QcGc96W#O.PM2(<eK&YI859B8PY,._XEfKfWeS&DRQ_N
_W-7MCQYLPEKIS+2H3]CGT9bM/3/F9B?G,PH^TcK9LORfO7+5<WI,S3e3a=:C;OK
A]NE_Y;_G\=>3Y(DG+;KIJZ,Z/QC7P9+P89LKaEJ>(1C8e;N4ae&+QYC^C3&)O.N
+CW^3NF0\Bb@J>E[a+F2UM(MO8PT3J,2KZOfa#9N^CB/_&3]I?F/>^(a-[-M#F[5
^F;\e[#gcGM\XJV\\eG:KQL^XN2<)</5_G80:_UFN.WUI00XGCI\KXY+cfbRL),f
+2]\_R6?>.S+4RG?5R^_#Q(RR1R/?UIO4QZ.DQ95d400d>/+0?;:8X3OE_^05?fA
VX7J;#DgD;+8R:Mc#J4d0WB9;dI[M5A6XHZU&KS4H<c;R#S(T>^6HG,S-05UOFQA
b()H/4dXA4E92<<)2E@0>@75P;Z#MdXFO89fPNd=5bb&G56TAOaE<d-:Qe2K/5b>
\PeC/05JARRJd_cIJB_a\IdZF0W8^8L).7dS)<,/<CTA@<X]+C#/&+,SGacTG7MK
-<g3U5-^f/=0NB[X3)8CKG.6I-?122/+\,FRZR5Z;(&JOQY64]TWcb.6^]c6(1I\
[WEe^-P\7V4U=L#L,WYc=BP9N]/-dGEcd?3W0H3W_N8C\gO_da0d-4H__J-Q0?\H
1E1A=AP12D)B:NTUE@4\7->0(8c;;?V#11YB)Q5VR2f59C9BRZAB4fWbKW8KGcHW
)(#SUB82+8=HBCP[]?M0?aG5dVGT#,BC2HSSHITT(=EIgb&1G\<742O=^7Y#U+D\
IJXMEGF=<Bd8-:gA<R)a;_fa1SORLA3[1(7&?>eENYGWYL596.B/]2#HEbI7P?=?
;BGLIV90G]N[]C98FdfVe<20[)2BJ+K0)1-KV+,IKbR/=b#UDYDM3Z9J0Q))CMe]
14FWK\f>c7:S=22e[O:_ggF35]SZI>;;PJXg.2I7(3,^P@.<H=H[b2.F3(bOa?WW
XgZK^71R]JX.][MDZ1<Ve7R=UfdQK)HDZCA#_CF[ZI0^O()08:+;Q+ETdIaeDK4J
&/?+GWP37#Q.7BJMbE9VI[D(N-fW2:90eR#&7:FK,:8&MeS_DRdOR/7YJZA\e:e^
b5/MMYR79^WSE1)9Xg\8[AWNK,V;HI0NCc;#X9Xc=,Y#/>^cSOd34-&5fe\fBC&1
Q6V5+da[59b(Z?N1/^IOA?+LK4I9387cG:S[DWKfFNBU1PRINSDF1WJ1&E+IbOKR
)4b(AFMdTQTE1(2E6(8W;@H\2V_cCN=7S47)7O62CE43CRGNdA.U27aO&IK.[D@:
#STARV2A6)I27<66D1^a:C>\6>^\CK+O?40@F.BL;PHA9:XI?DbD#X]a;S3YEA_C
Wc?0I7eN3&SBELJFX)A)b\>_FNV\ITZN?H8MH^Hba#d:H?;7gO8e<V(/8Vf(CMOE
J?]^GUJ&/=)X@+GYT0[)8N(V;BU@BH^c+b)R>62dEfK.G[14JL\<59YM\77b(X+f
bR(PP-@8PZ#;R@e5+>NOPGR6^]>5Z>gdSIYZ&^d5&,\W\BQcA@\/bK0<9Y&bZ:8;
4<]>S+\J?;XJ@_S6Y)/[@HBKgLa38f?QO66Cc:?+dO^d/_2fGI[KRY7e;X2Q[Sb4
bg(b:+?]\9.a8YD3ZTP?c\#f2H+-6\e[7VdFfZ\F2G17D0J4bJ=&X,PF6(M5MZJI
E7#JKRYM5C&d?SZ)/;f_^c=b-GU:.\f^I\^HP/8P7X]^G,)^Aa81ZGVcZ7cV99:D
OAdT/X)P0_S6egeSC8L8KL4J=28TaV&_2Zb?J6+\[9.O,L-Ac7?c@0R+@),3_TUf
Y6T613._XQ&9gU4?=C]F\5&(67).LZdI02_T=8P5X@+.&BV0\a=(9X2F]T((-\Z-
-gFDfR5aZ#<KL(F2,X6&e6HPK;1B[Y52-2XMGU=#:Ia4?,0GY<A58R&5Y\JCOgW^
36AXN-6OP,Wa01:Uf_4BD/f@7d#4NZ]ZT)[OCO/XE694A=?1680NCZ;A.B<?F=CZ
=L3&V?bUe=F]4\&U>T@6G:>N^&O.XP2TF#Me#4-0=O&Y+X[K;\JITA1^^:RS>7-,
3d?;=a;VFd[<EMJ?f3>c<A87b4S#d#:R4-OH.]&-YGbKRC<QTA]^TM>4Z@_YeZLQ
G[Y7_AH./@25]UEBdD(0/?D3KTgA=BBE;/4VHfBB@UVf85A=<T\K@WRNU25/I=M@
X]cH@X;De/bOX3@7bdK/V0:BHZffNV@^bACLE(79B9G6K@GO^OLV0Ac1YN8C_O5&
(8LH+VK/\05FTD)X6&-##F=:#Q;a;ec2#bQV^b6bC2J/F[INd\eF0@.S>eG2:?8]
..T/5H;J6B9B5&#?MIJ7GBcU@K-[I(.^A4gVaA1JEBBL,D(A)g]JRKDe])MZeWgc
7236Y2[EJNI9CPMOV,G-.Nd8d;V[Mg#f(aG4+0gQ6\-;RE=IT#&DJXGP;c<4P@0D
CZ;7;LFU98KR?-e@JB[W>AI&1?B7:M8/NZcPIE75L+a)<(TSY8/N2<]LS9T3)A=U
O&Y\IE.T3H.Cg<>+JZ,06E2Sc^<H0,^\#4dP.fQ:\BOE?4\dA8bW0:c=8?d/6EXf
UWJ:QX,.8&[fggWKSbE(T3fE4@62LTOGC^Ig#IdG?]4+dZ_NZ6PBKbP>@):;DV1T
e=P?(W6bW\f-W<DU=4I.#+\.G0V=H@:M)NGJ-=bfJcfbcI.=PTY85gdGM:dZ;]X;
f<dQF<&0cAI5WfEP^D:#ENCNNX^M,=O/fFL;d-255A)_R92H4DY767AW>/2E-/9?
c,](6d[])F]<]&5cBY<:J6;L8U9<MR]KE^U_(O\NE&ZA[GPFZ=Sc2&39#RYaHTdZ
[dT:\EJ78dGJ0N;1.bE,Sf+J:2dQB/UL;1#c:&_C2JK90/X2g,I3Ka9HH[D&ATdL
Z&TR-(?6P3[YDX-;X49/LM(IdSgS+X:]X1QQL2;Rd]OO=#=\dM7YHXB&c#VAFUGX
SY]bG3YNFS=^(?WSA3=2+I19AeG\5)7GE&I7;P^45Q=c>BBJ7L.g6GD/JJ7XQWFa
Y:M/66O5U:9(#0B^A\KG?QdF:R\M_W12NPM_1SPEUcX#.4&,X;d/a7H#:e\6,(N1
A_@_EB:NHac)^FcA-Z-]5IE6Q)-g+]V<<;0/&ANU^,B/F75X[1e/0(\RUJGZ1J:e
-,8+6(f9;CK=@e5?+aW\Q5R\S[;>FJERc880+9SL@(:\4T4-PVb=B1EF^;:C1YY>
Xf@O[#MF7.S1Fc1RB6D1M0U7O@cUE6Y__NQN15K8#V]I7@LWBQ+<(JP=B8#8Y&ZI
c_#?0BdO^Uf.FK@_GIe+RK;eH/Kf_[:cPIN/f11(IFdVf\AW\[f[#<Vg0?S3aE#=
9g;e<4eT8PM.E+^/BX.GG^2MZ@fV;g>/1[;+5Z,V35AZNCP94TXURA+;U;GEN^-2
dcaO<d2,5RI&^M7R++c1KZ87ZZ]g>Y)2@9>^8(8=MX<X(7?d[O;SeTAg5_P7V^.1
M6eGL=Sb_2d&Q^4UVBAT.&O]DM9O&QeQ4I>Vc0_VT.:f(GXc,_N9aGT./@^RL^00
]=9UB<GY78cX8EbP^W[[<Y_,_^C?^;N6?QAK\_:+D,@F00dAB:OQ5CZEB231=G(e
G=+f#/:HNWG)UP(80+M8BFfVT90P-8@RQ-Yfb9=XIEU;MPNG=Ee?E)VId/fT-9B7
LK:8F,TX-.0IAMg\IK+0;1D0T\?UQG@:L&Me\c#8-dIfa[@;QIdXQ69Ad6O&aOKJ
O^?\?H[d0^HRK:_b+/gT]KJK\0/WRMK=&/0:9(&V-0^cS]Y:e/)7R[gY6XR:#X#)
S^cI85#c3<F(g<J[dF^<O[e:^^W[<.J4^:QO=9Y]S]?81b4cAba8_5,3R7+GQa=9
K4AZFRV?VQWDP@da\FY8&A@8fE=&45M-/.1&N5IA:8Ed:75?,+)MNf(ODc]\77U)
-8-L>C>.#.D+Vb]UV&)K8+EFC<O;P6NM,V\2R=XJ[HfKV>0cO&E63B85UH@ea(6>
L>g9UGU/@BX>>S=gB5+M2FBJ&>I/JO=b(AVRAgE>69Y>N5e4:0H94H=T7Y>U,.FB
TU/L;[-4cVZV1[I@ID:+bVgc5BeO_ULVL]70ZR8W(P&+BK9]B#g#VeHV&/>]#4-+
@g\\G4Q?,4F0BKMb:C^NaPYf9NAH7B4,7<8/bW/N,(HP/<?UEF4RH_dSaED<,)9f
5TA5.81#-<AW#1gDAB_O-\E.[2Pb+-]W9GO6^4UGEVXE#DW;faEQYYF0?.9F&?K.
^7.eG&QAC6Vg=?I:.3O+c:LMKYPOeCQ;&Z4T+&KMaf7eJ5VI?1C_I2Rea8f\MFMY
^KcA-4</E8E<E+dO5Y[2Yc?V&=d\^AQ<7;F2EN@KJQ.?Z+B@>e<O8&?9R,_V68Za
G-BfaHOO0I(@@e]LIID#C]0.2Sg82Z4LHP/fa6^_8OD_<C;(JK]ZPO)=C)2-7WT[
99N7b>#?>220&VI8=@.#B+eS0H+Q-6Za0IQ8C;4[b>+>W<#[D[VH8Ld_;2A0_PJ\
]<^.S@0G_T/Jb@00TAJbY2Y5^c#NfdO:Bf8FJMXG_ef-dF,?AZA.>EDP(edWWdI^
gQ9ZOT/LNW:1a:PcQ0XI-5<PQN,2ZWHaa9OB1<N-]J>8N)+^-@UW;#e5<2#AP>8=
TaWa:T/((X[<V5/7Ygb4E[BFB9aJ^&cU0V?(2W[Z]HP;5AUEYcD5aF3@CON/[3/D
]T@&6]-41RLV>35fLE\K2cT>K+J;N72M(TD6_;74Rb[6J:(S1^4)SP[B?FdUgT7G
FTbC79g>#WH_EQJdfbT>Lae6I/XebZ_eV=J)]9^=_7aX-F#-\FbedARDC&ecP8e_
,a/LR>Q9,L4[+D8(-5dTD:ZOZ+D][Q0eHT,)R&ZJOfg(6&R<KVRc35H]Bg,O2-WC
I;;U[b1H,?/FVL#Fa,aeCG_2+7^:H;6<FcZeY7UadMQec/+<2Ha+2QN[@ZJL-]@>
0b2f53WT51T\Yg4Sg6U+R>\e5H[JZI2EgEI5T:_;&9M^-LRf2N0D4N6JCdMT(V.4
@AZRI26GWVa5/MDKgI#9f1GMND/.CQ<a?EKX8^bW?cF0a5?0,6>[3ZCT>gG<KVQ(
R+1;gGK3CM#47O7:P?:-AO@;LVBK@3Q3A;2acBVHN\0L?M90dJ.7.T5Bd5Nc0H7<
L[CC[[SE#7/UJ(5Hc<9dGc9cF,VbQWN<G[.+X-1F=GB/@T,9U#3dINU^?\AQLY<V
BV[BG1LRS@0(1SX0[CU4VQ2^I),N7&AgIHag9]aC&E0PKE+NPPc[ORJG-G1PW^?f
L-OY;3MDZ#9#>?>dVW<]>C;R4b4(Q7X/<7J[IYMVH;SeCSR1cHUKDA];_g>@e8V:
UC04)F&DR1SH+Z-^^]U.M9U0&]O]L\Nc]L.<JH=[f/GON;a54;b\8>RQ)IKRV0T.
:C4Y(NN]8Sb6:9-<#gb;=,GZD&fRZ9<_#=HWHOBSbXce4&.DeW0TG>GR16[D8D4-
H]U8^[>06]WN&=@[[5^^E@NGGO;:[KLS9(F-3^3B]2aE3dRg,=\b0f/=PA:<:.#E
4CYD__F^W>JRP)c4^U^e59g4(C[.OK7@bA4[O(F](AV67\/>b[J-BBN1D+LDQYP_
2gD8,a:e3^/7ZV=E9d6b>X&.9>IgTL6@)7UEH1<</CD_5F^.b\Z9OQ>3Y83&=7<\
f_^VFT.?a0M4QXYJ6@Q-P-ML:F27-f\C\S74CQI-6)AR4fR==OX8P6g_8USXBBVg
XU#CA>a\f3IA3ZJKK]bEg,5C><UFY/5CN0[;>TAAKZWI&>PL93b4\.B[:ZIW,3RQ
&R1_<S^:a[d8VU9+1AKX)-#F)+?S5RLV]+P.:7Y\\R(Y#4/0HK6_fLaKAf^\^E)<
P9M>CJ31-57c2HN<b7b5c=Dg(KL[0SSOU]T5?5J/58MIeTS/fH_+T3Fg(LH<8[M8
O._VJV95P6J3^AJF#_7HV;Mag6USQ>cUDAIJcN7=L=ff3UHNHD>c&LfEQJ=:NP=K
f/JOPc/@2&/ZY28f)@[@NMNM6+F-4?#&G05dZSCZU.MMd0@K#[f?f[g#d9P[8+2Y
d/NX6=B(L5#b^f\<Z2f[43?SW8\IXCVHT>]KG&&4NT@EMBWU2=L0e&MeF>E\3FR=
?V419AQM#Pgf82\OQV]=QUPCY)]EK-6YK@MA2UC:61f1[2GJ/55NHcSe<6S/[LVb
_g94=H(\bg&7H^L4(S8+;<4^(01gDRY54@+<D]Od/QD?<bCH(PC-]M&)-^XZ<S7W
[E7J918@?WH@UCI:G327^5K-0;<)F8E5&+[150?QXbDcM0T89fJZ)(#LSLVNW,II
6QW=74,P7Oab29KNC0TH_Q<6HQM\IaPV0VI;1_9Lec-]fW=aTZ)>Ag3D=JKLc9HQ
-PQ)1KTNGCd->.+30V?U_71XC+SCEU#1E9LbL<bZVg)1^TS<e-A0^#fb(9#/I2D@
a^f0@D2MWc>>^7ccaaN)&^=IP64VXS4L(eEZGOfXY\<<BD.L@HcQPM.bV4MIM+@^
/8A/8c1ALLa,2E(O2)PPcF^=(/eBW-&-07G34+(#3Y>;>M>Gc.,6#C:>K[E@2_Be
O]WA;b_b>2U/:4dW?W00UBZ<8)ZdTF.BeS=B0,gN^DB<?B:]cVgY78TLU^P\+)SB
35IB/\@OXVWANIJ240f1:5eQBJ>]7I)bE]a@.,[D]B#::dS#XD;<_/^[L+,,[D<.
2IUT9Pa@Z.[cLPUWDY))NFTW-DQIA(;:c4_W@G\&VUE\K/502gB.YJA^8gDHQ_5O
:44e38c1UN(>&6>Z9>HAH]J>;P[[WXcYD#GQC>79cbZB+9N,eTG(Z?UQU-]\;9MA
;+BA>Ye#2YX,Y/\5;J([#Wdd:NEBX4H_L0_;9^2+L.0I\HEUOAPG@H;U_K-Vgc:;
Y&.9\a?4#\V_QeAOBJZd<:8D@O?Lg@BaGeT1IGf_K_eLPD9<&K/O,6c36K//MO:Q
bNM]F(f15ZH_D.D0A[S1E@WcOK1=X)4WD6#^SA(R.E:[&MKOY2TLG6eS5EY8NZ[<
^_>-6>Y+3g:HBEW9]bAe+X^ZE?6cMRdJaRP:_P9Gba+e3\TEA]dZG@1)LB[.SLD@
#F/X,LP?5#Lg-\M@J#)cgU)7()GQ:Z+2ce6c/)[g?IRIZdGHBNWC[->gS8R0?#2/
f<MbbKR2f,EM)UR)DB.bS])9A_?&3YB=-K&5O9>EZ^Dc>ICg]@0J-aCdVBBY(>O?
.^:16)E_:0\dIeI-a0ZGKVWf:(]LDFD4+OaC0)9;gH4[Y&<X(5AQc]YLZVDIP<1]
TY93(b:HNE718aG7?PS4EC_2GC5+LY6BP\Ae<=CN(,^2WB)aZM0ZA)+fG2II/W)6
_@Eg/BNJAXFWCQ^MSC8]&bea,HOXeNU#A2&GKP<b&4;MU6SF_JaKA]SUQH?/I_>-
E/b?+S/3MDd6V#1DH,N^TVVJc>)c;UFa+[DgHadK:)_0aDP#c]ca)\CL(9S,W.Ie
g^+X^8/Ea,Z?V+OKDgQe5OXaUM07M/-O+,PgFS+,(/08=45[AA;+:3>M(bU+^L5)
025T+Uc\0(IS.RAD\I2N91gFWa=2Kb?X@PLF+fP?7CbFF((UO5g;JJISC<-L7QSU
K902[TSe&PB@F[CEU_,7E<LZHHg:=\PVWc3;G3,]#B]//0(Y#-0a/+^)6+OU[a^L
&f<I-8HV7F#\2#5E^ae]0&_88MXYB)-/NMT6-Z&FO82K_5P()@MIH&RHAC^JVdbO
caf-JC\VQ(Nf.)P.TK0B:gYPT5\[;W66Be^UYf?M5d#JORGV[FAVD5JdSb-_e6E4
,+KNf4.ZZW_&^9-VUJ)6PXJAODY4I=e4S(J-QUg#:ZMLYd_A6aCP9&-<c6M0;AW[
RKV=XQd&ZcHI/EfC\12KUSA9)CPR,gX+0/A^\OCOFV74=I(LMV/_^IBZ(@E]IC,2
V<?;B==#U8,R+VT8/f+>@95[?.HX^Q4:ZaUfVYJ#S-gKFBB[c:_6O.LQ&A[2;-MF
II<(/^cH#]?5]\4WF@BN)YF2gOHI0#FRN)-P1,:\H6(?BH91@E-M09SQ\G:C_&ZV
C><89FB<_Cf\BP\?<;P5@A&;-U[MVf1[I?3R#Gg-e+XGgYE@)f8LQfVQ6V@SS6CZ
-[AT:FEW6R-WSS3bECY8DKE8eT)>7_U>(94[<#X6O;J]&+CY2f+H(D\27B^S>Y63
5JeG0/@QJ9<I#U/LSQb@[@c[.6&g8P[1.gH7O^I05+caLFF1?cf\58a)=MaU3<0M
RB5V89\1C@T)gT;[aX_-[&72F.LQWO159PQ[1>T(=H2).G;^8N:PNdAFJ:PCgNW:
09,fG?cWI]2,_80DR^_,9PfGWa#/Uc/VA>8f@N^<e.eObZ9C/5bCZ@664:[e7UJA
(<,-[SVJL9Rf=&9<EI/^#?&V4aU&2FWHB5M&E];&Pa:#M<><2L+/3K;1aZ7-:b=R
-S3-^Te3gLV:OUL3+MZ_\abGB9b1/P)L[OPVaAB(IA34DL[17W0H#f#4Ee6&DZ?7
:(PG[7gDGZ#&c-GBT/:.,AGEMR5W/a/=+9?3,7c#WQE##UK9IZ6=8dO^A,D9A7=,
]ZY6Wf7P=7)4^81P[e:+W4a0?ICC9FHQ)&2IIY+J>\-S9aN_E-<JMbHULDT,R&f,
[&2YO7DbV.&^.KD#<U.)O)>S6f?\2-J4K@+#gdEOd^>PNPXA,YNM3XLA:8)5&,T]
Ga0LDZV5HDU[@G:PJDH?U5)\U/&(=IB1>G=\+A9[TXP8/gE=QZ<e]0/#@[R89WRX
OfX@OR>b2]b-Z<8,^/AZG;cFH+.c6)WbNa6R(9ISZBI@+OE=#?J2]N3cK)D)bEXE
d-IJ1V)L=OEL_,UVE#4RUPD98FK,;Z6\F@D.+LgX(-J\J5NF8SeEbM6MMUJN+6R:
G\gZOc0cAaL\\XJK,9[1K[Nec4A:8)aC,E09L89:BOT/DH^g/gOg,F/KX0]D8P-A
6<cY<PdM_;00EHbB>MMc0)QD=0K4#QL42\.@U^fI:AP3OBKIe_8FN0=KU<=4:e2(
X7eg.N2Q;D5aICaYLKE(8(6]6LU#G&FLc,Qg_1cg_f#&W@M]Z&MX)dOb.HagD6GC
JBO<S_P>5Y?a#bIdMa@6<9Q<ZC(@SR35Md,[-89>I5/LfK(9(O?[N&ceO&\e=b?Z
Y=>DG0?4K&6Ggd5<_QRN7]8@8GF0?N2IWT0dd&d7U?dAPQ:7bd]4#;bUa4@25T<B
LPN4O=\K6K>eEU.NW,1eF/g6OVE>Y0bfBWZU=E34E0N=b^@I#V:S#<S8_,H8UND(
J=a^CD&cX/6H,d>R._f-S3+]^N5ebb@B.V#.B;^G49G-B\;63D)BH.WE;,.D-)67
T:2(ZT-[6:5V,G,JNZgcO[TLaKCA.bREU0gEc6M4b?A(8d?D_C>NZ(<g#S6OU_&^
P2Xb-2cfK6=)aL6P5^e82):PO>b+Uc--:HS[EeD?<).C;ZLc2\(A(B1WXR<.)Wg_
cB4b8aD3Zb#e;5WO^KeM4LV/,+AM)&1@+cWd4:O0HX.@I;)I8EI@.g;TS?6(Ea<R
IX1Jc^5Yb3-J&g,gJDW:bW3_7+45]c,Yb[,;^CdW_0TI^)U#H-1ZJG.5_CD/;XX8
W2HC45U;:W)U1Y<\eHHJ3^_WDZ.UD(6&[+?f>0=[<7T95c):@N]D+0Z3:\KOQFEG
)PQ9-&Y)9&Y4_[EJ0LB3JEK\6.Z9:<9/XDLccGV@aY>_,WZ)6#(a\\B=UC&IH29.
OU1_gfg2J.L08?BeFeKHb24;K8:::@LCU1<?TZ<Z8_P&(>1WFc:<,O#[0_9O]g33
EF97T?F<GX)OLT-ZF\9E?6ZNU+Hb):d)/R_7-)B@7+dVbJI\JEUP:0GS\:8dO@G7
_,)=SfgU?03efcdUL.]\:1E2:TUZe+,g.M+T@G=4<^S^U6-.:^<+/==21A<d2:[Y
F,E?K;>\IcE@[T_&B:M8-0MC2CJY>NG;]ab(A1Uc_F0X;6)0]R6Z8TQYP-@G&E#0
J/,HZNYdCI?N.W;f2])KR3KX\AL_8-MHY+HL,8DJ2?d@9]@Y4;^JQ\_7L,@7QXZf
1#3/-HY>L]Ag^2F4c(PX=VGGB370A-=VL=E34-T:#;<Xa:M4]:)8(<3gKFX=<3J0
7F.Kc#UOUX=9#333,f&@CaQ9Yb7M@/aE.Gd/_5=QP@OOa3^/([R;(8SF@]4[7+0:
DBTEN<<L;?K:;L[B)JY?]P/Nc1eE90:I7B;;=QBDRP7O24F4Y:-f3+5].3W:T?a]
W:a1VEWfGZ[gI3LV#+-W@(X?GB7IHAVf^0MJ,Af-NIc:-(W+&g@PPOQ/IVRI@E_=
VZ1QJLd-P;_e=\KB@)&d410dL/D<?-S2e)4H9F;d4;5f4,PFPN16R>P#NS@YScB_
>79@USZYV/S]^U[J+.ZY5+Z#T.X@V6J4_),X#]R1<89-U?^:J1cD=7UMASO=GM(1
VQ]ZUL8,FZcE9/A)I)ME#9JLD>4[9O#95g/\V=B;[43[;7F&ZH_8Qf#4<gBcYIW@
<WN2KIP8A1-)7E;QZ(Z=)@3^BWT[3d]FfXIX0DFVAI]Q]5XRgcUR=fHcQGPP\DfL
_2/Z/6C[C?TS+A/WFQAF7d4fK;=E^DMG/2a#.2(^R8=@<P3Ie<E_b]g_P,NJ0e#E
SdEO_S@WF,IP6\.RFV0R-Md^+Ac>dAS0\4E?J#B.<Q&8e_Qe[7#,?6J#@7<de(KO
&dA58JHXc8.&J27c<FD1JN-Q]A_bOcLV&9O6bgF\2@^5FA:D@FW]85YGC,_Id0&+
N3GM@C-Y6^aN7fcgH:VQ;JfLG1Ef5>L]GR-ga.TL7X.F-YK=9<>^Cd6ERgHJ&>OC
8H5M^P1,T8a:U,4YY)3?<:_<#SeA-R8P?.)+)JKAAFf=_;ETGR7O(e@>dc+eFZ.P
M_PO;.<Bf3+;VM/Q.;<)[K7c;\B(G48W3M(6IEf;/[6RPM@IQBfOaf,d3,=A6=CL
Yb#0)<CM80RKX92=4=QL#2EAC)d?;ZI81-#GS.6HW[_b<7aD,T;P03I6_cd5ZddZ
17&\(;_8PTS]JWUI5L&\1CFdSg3W+MMY#>7,7K\VgM^d&65f[&d]CYc]ab-TPG_B
.XD>e]^Ia;W_Y<:\bC<=C/X/5:@7_d[1@)0bG\FfJR4#RA\=IM=\MU>PUU5>7F[L
f\W,f7NgXggW2RT1a5(;_GZNG7IIb=4NXI<=J(6c/(]CWN>YZ.ZA,5OPN5(O8^:2
O^#0b=29._E2W<9Z,CWJI.CQV(PX,dBSD]IH7YGgJffRP\-)DeQ+-=b)U(ZY=;18
LHBVPN4DSU\<W3Lf9?e^;C&E?+cGN_=7QB9)4BXeZVfRIa>8f7#GC=(Wg@L\J[3O
+.Zb0dfN17Nb_LB#]dWIQQIe7H9eB+L_G2\_C#gN1SfQ,8JS,]=HLD:WCE)0MbU6
S&<41U7)5ITcgLMc<X/P0X9B_<AF/PXCJ/L,&6GH;\O\>)Ub.6,(7&4M^5g@X2MJ
f_>6IfR,;^LW(<FT:\F+]GH11gEZ:;UVH&^IRTC_CWDa9:[TLQZg\(FYWC-5R;4_
bf5DSLX9;f=G)_22?cEROL_J(I9DBJ4AH>4+H^7O[K7Q1H_NTc4a#D+NM>QV8;Z(
4IE;&8ce&6?)-LDUba/@0A:f6-H9@3cYFNdJ[Z=?00]U29D;P,IgU)YH4,5^@U]2
JMfd5fVgUA&KH@d8-OY/7(SBR&G^TQ\?,geY#&eO+(3c[T]YL?1:+V9e(S\(/_D3
1V\AG[a/2>J5+5NEP3UBPB&1BfX7.CgP.fcL^Ce]<Y+,I.ZM_0/gSUc8M4P?ZZ2b
@T-88VN):-KL5H#\MO:(MK#S(\JK#f>+b[d7IJT^[R<cA;e]._^UdJV.5EBQE=2B
Cg(O?W2PIRJT.(-]FG>F]&YJ6?AF86RY<&M,?N^G>BQ#[.R,AB&@d<\S)M\DO7\Q
9&\,6e1Q+Lf(CW-HQ(;B?<BbY&2UVY]/42AfdXF7PAHVbK1(5@@2E2)3Z<b?&LG.
16:BCdQ4_Q4#eDK<J4cZHe07G3Qg)TJWI(MbT:(XH4[g7E<]W15=<JRH3F:5OgX]
fJeOH,=c-L.4[U,.>UR0b;eJC^e-P3G^@K;4YNH4?/IF7G@da9PV7&LB,[2YEWXB
La(CFd1[NM-_WZ6G\):>NU4XY7/CgD]Qdf?+^9IeF<YSOE>:4=bG-g+g/\&HNB2?
(.<Kc2OQMMaW-WV&;(W)Pf,NYbZ?3gE,-Y\IE,BT#?Q?XFO)TAG1;-5egQG9?@4]
;9\HT:M5ERG40(f6M_R=9I>_#?e<\IcJWI^cJ&^N(4(WZ)&[,[\46.cIU:&J+(+\
,?HN2X?a@Hgc)X?>I4+=EY>H?SNR5AKOM.B[B@SNO5)M>(0STU]I+H@BU2aOTT:N
HA&:_6]=A9IBg>Q=\;]a]-#I))a5UFZbU]5@01X@MROdTGPd\F0Y8)#&GWLCV;\3
_MWD,aEc\BTR]_^dRcDYA1JJ0ga0BBZK1G<79WagR3SbXKa6)-d@7[VE2B]/;=HD
SeJTRc+SNe::NC;6HBU?_QP_M1gf5:H=E\IDRQ<0+K]9\9G5O#5K,6/Y>8I;=?C8
NFAY_7Q&8g^C#6P#I(S7/;Q\=a5LgG1Tc&G6E8_)3.R#5N4E/dK2<4X#6J(C?K0R
.5H;C258<PDSQ](e682<Z/1729e&ZYQ=DQ_>[@LTc[A.:&21<gQ)@fR6?fcdQ2@]
g7Y/d1]b<F\6e[-3QTOXORF#g>fg#2FIUbIBS21>CKdb#V,g2TR8=V_cQ85)N3fd
VcR=II?R2TR&ESObM=LTPDWYR7dWaAg+;5OEM?46_FVMO1-=:da42#K.UEBf::WM
NEGBc&A=fB2V6PWZW;/L[6A5#BPfX(a-EY5cg:H#:#_U219<?T)DBSPO3G8&.ZPd
eIQC9?O;YLfL8R4S3XOc:,+/>9_[db2X&S5PH7#<OD8H&NL5(\JeeBA3=Y7W,Zf)
DQb-QR6Ic0JRE;+AYeT4<&ObHJIQ+a3d&R(GF#14@Rc@0I\CJK>>@KX_AI\cV\1:
,&Pb_WBBA:(W)UF?BY>D/Z6G]#>ddFO/6EQ895#:a3</=e]N;A;/D;Re2&?/\0g,
+dV21E<7,2c(KK:2AIZ,68NA1IKIM9O:fS26@1\Tf-;-NLFD,cZO.=W2fMKQ2^89
_2#,eQc4]d=cPJMI?J5>c,,F)M-Q>LJ^[P]D-[G:^85J8#6O667Xd?bLQ3d2cB8C
d)CaIY&EJaL=,3VcGP[@832V,\Z<ZBe>VePJ^8733f4TOGf>>QIGW.e7+R3:.?1J
c9ACS:&/HB@DB/e4O\(W5Kf5CX0O&/JPg0c[D:2@CcEGZ5#;VD^R&fPI<VFANF.C
>C+1I5GY,4fV;dL39_I&Id+gRPaG1UO/,/[d;/+1Ud]8PD_FOdd</9&&(ad(+[+R
7HH<V(R6VggENY&V=P>f[,f7f-8Y&,\FZ[;R0b)a46;#L+HIEUeJ^+3A5cIQ-0O)
,875TJM+Q<7O^2K-Q2EdAZQAR1M_7JC6(BCWXc3B>JPA7/A5T)@A4ZNUTU)&Y/BY
5VDd2&Rb5f?1A,<6[U=K8-A(,,?Y.?^(74b15,2;;AY^5KC4B-XJdDAJI3HP-a2Y
E211>OH.(G6ZK+)4RRRNBPWa7d/##:O^_R@__T^ZgPe4IaF.YC4B2+7/=Wfg<_fI
fCV\e2+GOd/J,MeaYW#QE<D[=gP)bMg2C:NHE#/)F)&\Md&NKaVR#>6+;?2Z2XJ8
-V@K[522dBeE/X1JLEfScGB3,2RMCNb?fOc<2A+JGUWJ39<Z8+(:P2D0D_#(G@Vd
6VQ\<@)AWe.Y6B49\7-#?X8+[2FDTQZQK;/I=>aH+^5PMfKR-2?#IQ[aO<H5@@-+
>;LfXNCK./=D64>&R5IWR<X0LVNEH)22TS?7faB=N&;BN[Pe<&BVAH4D,M1(3WSe
TRP<YU2LW)\XR6CD[3=QF1BCF<3Gg/aT0fHf:_76gKL#I+C/FPAV1(QW5BQbZSaF
<f=^aMI9Fg_MUXIJLV2;X&bUY)M]a\[]NA=\ELU/G\QIE3E\?)5dg5f089[9D]a(
+I?O/Id[4&?c_V1V[b7bNPVEU<VMcT=TY]I7G,)+]?(U,5Q2d[-,eP/-0Z5G5OZF
,Bc0GfgU^65S-S]f[3UNN=4+;Y^N,AO5=f9,bFF1adEDOD,+P6L:1][(9e-(D#,#
Bb9bF7IX/E,I)VGN.)71bd0?&LEPMFBG[#WV<WC)JC>,:g[;_CUdMGcU];aa_^Pa
&B:H[f^C&bIP@3IV7A4dP4ML6Z9?VIb)\&(VH/+OCNK;g2@/Ce6L_^2>C+cD#TJL
UOdb@C;?FV(_?/MWX6;-6Ca/[U_8/VLS./A/L(U4>BNU>K&Q&NT/5WK\G2-B6ZC^
fK4(GNFMBWg\M-GeR]eO<S;8_G?\R024GDV@GP]cQMGd8D:W5#Gb]d2:I&V:^dgc
4(7&+H?cAM=VHfcX/(7WQ>eJ-<U/DNYg5W1HH/)VNNGUILM\3+=VJY3U>:Q]/Z@Z
3(dNIGI-KDUVbZgXB@V7/\C,4MW^KIdKWVe[C0NcB4KY;/deKW6Y34I&6FTY=D#G
f4<1UZe7NEJYY-DE^c(-8QWIe+LQ(+93++/+FPeS:SD6V>Uf\T\+TR;+4I3Xg-9K
47>=<\IVRM]_fbS+<\IZe:b4M/2:2<IRKeN?29(b1BGEdR1&5+OIV>[?cXS)eI-[
454A<9E<[>F_[VO6I^;6eUg?05F41=gX1c/<XWKN^7bX42>4Q@)g.>Q4[GC_E-aX
9V@WKSaaF?gg?=1bf]]#^:&;A<+T<4.CP^#Y7AZV[-M27:_fZ+5MB#X))/e3gRa5
RTb0NIBC>d[O1G>E;/^4Y.XSBQ?VMe&LVBXJR+I)>QK.]Q.2F4/L.Qg3T#\fa0CJ
DV?5b2gPBUULVM.ce-41Z1X9/BW:UAS.Eff94G]U8=:FUJD6)HfGaFM.<Q8&S;JF
<5N,3g45_IL@\MD>.(?6_b&?(MeW)5/&M.N^.CdF_f^J,;g38T6F_=EJ:ZA&3H&f
fC?9,,4C;EZZBMS-BB5XB911=3cAaT9+0TA^f=^,KK&Se^=Z6P:N?&OddD(D7P0R
6GECWI)M@#LT,]>X?1&J0f4<=Pd0Sf(G=AKYf=6aAbcSQ=YZdXM[^@<f-^1cB(3W
8@C+Q72Z\:)eQH3E6XJZ=He,VGZ\U,Y:ZEHDS)E0@@<@O57Q[geg+\cgG/1BV:/-
N\=J+,5PdW+&?9-].@JK:=?M@O?GQ>1fIFSEJBQUKgU7:8WbC3T1Q(:N9XO2f&ed
JP::?;0;;b?TJJbLbD9]S>\+B@M_7@GGG4X7b0:[##a]E7UMSM-]I)5_GA(9<e)H
P?>0RR1;YKZea:H?g+G5e71fNO:.QCd1?>c_agRgMgdXKJ;RRR>_96()3E9Ab,MH
AE<04f]T6WYDbCN65daDOVAOMIC0VO<->>^CE?7^/QPRO7/X.LbK<fd.+CQB^g:_
V_Ig8HH/?F;//BLQb-A2U,LQB,-#d5SXgWEb?R6G5\A^5>W23.8c^=BP>;QU;;9@
>PCJ[?[GRRH]EZ0C6gBFN;J-])4M-O/R4E&J]]:H&b&(c2:S<1GbH,1,,Y9;UIR1
84;RJV#0BI=T3+daU]HBL,68\-NELF3]?N6I<W[d7(MLTL(9ZD3ZNePSg9N93NXS
17X^SN;\]+eW?#bRF\9ED\(8@A&FOb/KGVD2R/6Rc2EB8:C6AdN5K:2GJ2(@<F4.
4NLCNT;6BNSe@761[HNe/cIa(?ZF:7&(/1GD[;0W5L_L;fbNREA0Q_YSCbQ1?K1[
f?W)2]WD(Yb9]<aCXNH4&:UQ[?FCaefdY\-+IMba@52#T7WB+5f\<&DPK)V;<_7b
)edFP7:1?(^O3H-:NG>1GNQK]JIMa-^5PWYf(6C5OR1/E(;M3QYe99)M2G6aGP\c
I3,,-YTL#a.ISMH5J5B2beJJ17<M^UH-A9d6UFaTQ(\B2gK2?@T?#5eJCP(:XN99
52f6AKaK3<dYMSeMH.cabESZNBL=SdT]COCXN8YT;^57W9EeOZLT_JTfb32SgKNX
@MJ[:_G=7f10KHCf/MK)b#IBaMg5@5<#6eXD@55X^(&F@5_N-U?d5/@:<O2E;g?B
(;?/XeZ>b6>F3&B+E2[U2eG=61eg7?eU+N390JTHEQ2PLb@fc#_SG#^1gH)3>::H
e.cW3FYV4ZL97+EHb>\d]-C?\]DXaE#H5W<D^4B7LVV=aE=VO)S>S&^.>FQ85>_7
T@<Qbg,J9BQ?L@)AUJ.FLB_;g8U?G?:5P>]3Wa,NDE4GFU&5#_e5H(e/)ALZ&fRB
Q.;DcM1MCZYH[A(O]W<@\3@TK+G,aVVGfL?LaNDX755M9.85@-J;U]bOMX#\TM\b
W?]J-TWMc2d>-1X-af-g?#,bM]7=+g<4<Z^d9>DTT]9CgFP/QGFCc0DK<<Z7X1B2
+11A-C(@6cJU0/9,#Hf1KZ7I,>O6I#O^FO=SFS,/c5MZf>8<8]R^EY<>:G[\J5:W
=Rc\D2Ig1+Xb3Jc;\)bN]<TTePBggX?Ha\8#RUM#fU9,#?-^DBYIGY2W]MLQ(RW/
Ye\&8=NQ1.fR^(50RD4[-a8\cFBN^5;H/3G&e8J;fHEA4NFc,_MX#eA;@=0\83E.
YW;CA2(7F<8N^.7I[5C#7T[E;&/OH;1U[adDQWRK(H)]U]6.T75MQM<EM]42,TK7
9[0I)0200S>?g/FCU#\BAAFE3JC@1RPKCVB>HSe_\cdg3SH^<<3e_NdFU-12b]1T
?>L3a3=(G:XT)Q85&AVAKfOGCVc9a)b[UXUddd)T4b)ZMEF>KL@QZeeFDGV\HV<1
e&H)U2;#;BNB?D&^PS/#4HbLZ^>(.a#aBfIIaADTWRZ/,Bfa\,@CKVXCJ@Qa/5,P
g>>)?D_XD;=F51#VZ0<BdT5G=D.CE(X^/Q+QF2)bC6#6V7#IT5+D]=)_<2X23ZZ3
VCVQ.5PTR,;R>g<2+D[66ZM_(KbPKQRdKFFUH1(ZB.a(OFRIII&R#D_Q_QJ=>1Q@
^MRPDH09gMef0]DH(,@f4LCW?eQ7\0b7EN&D-Q51BF\V(RWP\,W?^#,[S1cbG/K0
XL5@)CXK-)9I?^PGAN2<F\9FJ/,8I<RY<OH7eDZA+O3T8I=B<:&APc]Rb;-(869P
2>]G\0gW3I^G\TgFUJWYVf;4UM11D1X(V6(8,W_G6/D+D#33H;FS>1DWIXXWO0d7
@Q>[?C1dVHUcdS+O;-[5LVJFHV@D\I;X58(<J4RGeR1D<Bf=9Ig)O&_P+R^Mg+c0
=G&VDE>ZO4<>UQ<H08Y4b[NO]N.@>=U[B62?@Q3B]>3A9YM_4U/_J1/,?N4@e3cN
W(WKFL_Uag)ZS6#.=>Y&SXVH(bH^dK3LFO7UKfIP-JPK[98._)ge8TB>cY;dJX:D
/>96.4d#H&[&cXUIHL<;E/.BeQGWP651MdO2/LB=12dLC@6IZ<[C;;/2R[R=9fA,
V0JJ=C4ZP@>\eI]:)\8<N&7;IDZP)M8deX>86:b)P4M(@?0=@e4H>;GO7g^]=RS2
dC/,T,;+Ag(CE)@S,&UGD?dK-2T\CQ1+8Lf8A<:f=WT<)4LH<2cDNR-Vd6PNQ@>:
#^TM51e/KKRfO;Y\\1PJ\KK^6L+)Y4^bM]02(ba^-<,.]V&41_2PM,GKcBI.^IF1
,YFa?8(Z@8(LI1a,@gcc8GABR#RG>IY,;>?D4S71A/YX7;0/ZXD5.D,YUc2S(&NX
-+=QUK7I/Xf5,A3^_G7<57?\B.dL-B8UEBa^;(93]>YG\R])7KJ[PHBKN0WbMOFO
U^C\/:3d:ZagabdKY\++V>#_T;6g.Aa7BdM#H+KN0\_d8;DI9We/aRKe184U)44<
19bBAM51KDT-(g8Y#LbS[B;f9-/_6cY.ggd-0b=LgcR;cg:c2V:I&MA45/e5=XG]
JS<CEK6=+]a^Q,:U17H&(VBgY]WX\g9#9b8Q#A3bM.X&<6(8M9S&M5O9@VQ=3^+f
(6b:a?AY4dfW28T(?a_9MP&^cB=[7SR)TP.9O(7WHHKE66883CY]@O[IH^8ER\>H
>f^R=(d>AIR4&6H2=X8a6-X^,L8HH1Z.4C/DPQNWRYW0dS-4R#b_E>EFF(,J(9fD
fQX.X_g[8eOXU[JB#&B3TR&8@C,2FNCN49\SA.Q>].75XYXX_d5E,89=<Uc#EVG&
+Q&eI4e#?f9H?#e0BfD1#AER.ZDeA8e&^4AUSED_4RHVKgGXW=(5.U(CG<LC..:9
IR=K<b(3/_(/VD0H,b<7a^Z6=0/4_bg>WKe]4cT(:HAU60[55C.T^7Z<agVF4#Xa
<&BBU6eVQCO;-a>RNAf7QEJPg.D0e6dQ&_5=0CY.CFA)F@YbLZ:0[?;L(N2JG-EM
:OIA6I)&-[N:))dSbB1<QL^MD9.Fe(J#H9-;UMCBI0?;;I#2ITHef7U&/c)A_HGZ
EA\JU2&:P4TZ]P+PJ>]E5IHH5e,#M..KG@WE[WYUK@8E,+ZRJCFQBdfS.^4GHLIX
;=G.<F7_^0V6W&Z^J;DT-4OLIT@YMF^DM]Y^BYM+T7^IN?ecQTP>J_6MD=HLM9II
1U>HF6(E&??2?BETPD+RQ1>\bLRb,EES)0ZA=LG?MY1e4D01fW[:\)1@7a)ASUWY
7TKPPOG#66JH35C[KR)U^J55FRa.XQ8d-]6=^^9-GD_KM+I85^R9Qe.:U\,;37##
&]S,#LOT8.[II>d#V8a#<PT8OQS0K=X=(=]?_<20+\^_XHQ35KM]dSa/:b+AN:IA
@ARDcQ8SKc)#Q;F<S0OPScF1X]8G3C@80N_,5A4>O_XWE0+G9Te2P61_5]MM^6eJ
_HV-9Z4H,#\+=X,:[@.M7aO?9J(JR5R<4ATC<#QKVKNIJb-Vg=H^=cdFK^:;\--=
3[f@,ZNOHVgBc4d4SH71[?+T89)?6B2.^fSW2YddC3K?fV03-WOYB+PX@U1&VKd/
d7=bWN+e4C[YWPC>\K2-#=OBA7Ga6?1/99B\9JM8ST;\_I+;f=NU8#[:.<T>gMWJ
7aLEV/8U@PfdC4Z=e8&cP>6P41J4N/:bI03??RT9/RSDa16eC?M.164/3GWAH^&B
-QPcNGHD-4S+aC6aU,NB_L=CK[(7QXg:GUCfH/CP:1)F9R+)CLGA]Yf&S1OOe2F&
BX6PDaRM;]T4:ee/fV[UD_T,RRY9[T@faJI8G&14[U7#fa&;XC<NC4Q?Bd&8&VaN
I<4I_]38-4dFc[OP7bf4:4M0)WY:\A23F3.0cDdb=D+0aC;939bWcE##2==#LgL7
BY2ZHQ2YJRa?U4\:GE.8U\65L9]KX<TcX8<<P]Md-/deH:ZGNP>d))YK/4]G/f^0
+4N70@\+7V1SJZgRc44;0f?Yb5]3TG1<_,Ff>ZG<A;,WOOCM14eL+I<88CK^9dL]
<fa(CcbNLH:]a18TPDXHL6W]X[gOXM&gE-dLe\g_)#BcU\:^P(<1PeP\4F@X/P4c
)<]AP<Ka>C2_//a>X2W>E)U.<f[Q1JAa&M+.Af19BFTZN,f)02@[UW6:TMCTXVT5
d89L>8@2Zgc1B0H,=T7#.E@&f7<RXBV(9cDI[#)Hfa9FSRQaJ+&:[b_X4_a-bJ)@
DdH@Uc#cBRbUNI.NT&g<]KJ7Lba.5b2IaCS;S[Q]gL[HK3UEW6)B9M<,UccU=QP]
LNC^<3#AN7G#ag@V#^X-=^Rg<4Q+9=RO&OF<8geZ1NCUdSO\75_2^DS_:CW.TA9)
,J\ENb<g=9eJ;U\H6db52g,,YE,,^#Y,JA.=GEQ5]19R2_d]I(YR43)P:O_@;UW^
a)KZO^XH1#ce,2FP4AQSbS:?]Jb?QH9252(7X3VAfTUG8<9\8^0[<NU]MI\AB._A
R,E8JH)?F8/NM(P/g579P37L6\NeS)7YB0&C)2/R:^-^?/^daZB.N3b\W+L?\1RR
/>HFZQS\W3W41IY4E6g)[f4e\.[+fRSUTUK,EHed/H/N=EYB.__C_>ZZ2DfC9KKd
P5DGU[c2/H4^)TY(0)cLM61K9dB[,?CYMTQ@II9@E0;<34)g<B:[->^]5QKVAc1:
0b3B]>QE#BIfU9e(\,R2>[W#>gM(.>@5_#>X_O:OD3,3SQ_bWaU0;>#U2.I[H\39
;:U;4LGM>?g@<+_^gFBbVee&3O7ec-KT[E0/Ua+dF9.)]Jf]J/LI9IW0^?R+=#Pd
0Fg^#Gc#[\g:.T[YD8@=a#a,>R@DUQM@BF5WKY]@GG_gRVHgG4]eBL-c@ICXLZf8
5GK+#ZZ&>O;D0P=KJS@X,BIPEPL>dNFUU4=PN[9Y-e&[=]eT@eN@\LgcZ1)U</VV
9(^ZK?DbdIZO,HW.FbgB#)c;7.Pf@B)XENB/^+BPOaY)Z6^\WC#ODHU4/U;6McH7
I_/CP3b[EQT=?,URS/U+:Y8W_VIA?HU/GN67)J5)P:WR[Ndf92bBdFDPN_g/gb=O
]/_&Ta5cLXdF4-;6?Q.._-U4,?/63JHG/BU91DM>JX>5=FX,DRd=PP^V;&<)8bcL
:91;9T.&BWLUZf)b5:8N98[b=F)Va>9/]De#F#>QGYdaI_3LSI,8aK:#Z-\e]9:;
_DW>X[\d/81B-P&4DVP&NJO7(2_NX51g3\6CBS>R8ebE]8A3]\#WAN9(9U-Df8VL
@?>:^M=b.24P0YfQRcW2BL6bVAdW1031I<+_\S7IY5/>H,EE43)H[3KA<e\W<dE>
5G=+)5Zfg:53V\#gFddYB32CWAP/^[J<NGJL,eLYI@<SM.;9W\8/(&DA+YV]CARd
Od=e-XD#A4G/[gYaf&]36I;BOJT-Z^M=NHcfMI&cGV,@YHAQ;(d5_6)P&.RBM4_>
g25E/[,6MGJaQ(-65Y8c>dHfHR?;,YF19Y-\\YUe3,(3-A7^_\T3@D9P(egZ(P(:
0=TI05f#)#(RU1Bf1Q?+)_BMaQF&egPAS-4&Z;49Zfg>NYL#0Q<dH@bJ(];8RfR/
LQ/S0+ST=XD>M#ePKXPXMH1TZ]?bGYOR/f.QHL_UFFD,N;E;_VLJ441:>6ODdM]K
D&S?D8=LT(<)HIO7YK+X\1_RK]S>9LLL-B[G,-()L(\g,CI_ET<UEV#]>G>\4:M&
:THKfbE-1Pa84=1&=>.LfU.bBC_WQ;AL6-:X>Qd+e0bCG7B74E=A1+P_6+ZAD\R&
)-=Sg>,YIU6^DeOFF4/UKG,J0=P0Y8E-b9A6K.2Xd9&C@d-M^]gM[+8F#AE95b5d
,\=+\S<9WY=-C>2af1PR#fAL3=e-#_;7]_gG,C(C9Db4AE7;X.4K1^4A=BXF<6)4
UbaQ&;8YF4?L?4QOQ@J>PS1AU,+X=[_.F4=-E]4X.(WGN5aMQ(F_)L+\fJCS>#]=
P[;,7Y2LZ+6Q(^GRT7TT-HS]9:E_A<1:^dReGb\O[W/JCLO]+A6SG.SaEJ<P?W9Y
BJ3NJYbb#ML/X/YE=46)V&16MBUEe8G/NP-=BI+IEcO(59\Da[b1I()bHIG7RAdE
1bMQ/:c:LM-0[(-M:PYcb2EN:5(2[GK[-[UPZ0[IE/)cgGN<6?4O^Q>Fe6VU9(HE
<3(_IGL\7:+gX>#R0D^YdZ1LEG2CNA;Z;\>&OW?A?_=c]G0;C@ZW\7JU4YI5WO#X
/YgN:H8/bN>]HTA])E3b@CT8P[<78O(/FITP()a3C,HT=bGLNPN_&J8,H>>>e(<]
bDV(Z[^_O#BeXfGe,a1EBHP7M:E8F+#R=6/_T?DIZZd?\[;VE<3T98X^b2OI8E:S
LLa>;=RW9b/g?4+8<2@cP1I^/WS)J\]A66b]OJ7[N29YfLKI@Y#+=2&JI0R-&\YH
a<8PW74fIfZ.16B;VLY=W,Y9f@6@;BMR90;9\8]e3K@e&aPU?,bJD300>3IYJY]]
DO,GeS=Y;8@6AR?.b.Z3g^9?Q^EXW+>Y5>T<H7dNW-9@ffBgM,6YZ9^J@D,6,4PY
)B:.Pc5PV5M_A=TL]4OI9/Y:K9Y/03?&PRgY?HH(^H>gLd?cP2W-7PYZWFN^&4&f
X<9BB-d&GbOD0K#RVE7@9b2D,U29__fC1O+A3ZBFbB)U]F+b<^@ZU490A=0(,2g6
R59L>8L(@B&VRaW]Qc507>5G&YM47X5)#GS=HD04G7g9CXJ_8d>_P64Z\##BUDG<
3HT[c?a&W6:X>dWVcfg&[^I/PZWNaFSFY[W1ZX\R,=A\XZ7B>:?:VQTX?YU:c:dF
a<;A91#30)L#)b@URQ8HYb,b)IeI\b=bQG7[-C:1KTV@]gNVK,1X^#Yc>)WKHbUT
WCc2ZSJS\I;cCDgBJI9EcQc6]TKQ(3<Z6+a+I&8PC8T?(9JXXH9N#JF<2I9e]/.4
^K^@YFG]@W&O/,aGH7XMb.CJ-6-1U2/5VZNFQMLZ9HebX:?I\-2UHKQdB]K^/.Gd
c7QGD_.53D3He]\a#^_^\S=dgf6.YLH)_S+b@M(Ec__D)QX+O/>&\-EZV6.S?FUO
P)IKA33M<\IH-7Ife6#f>@M,<(&Ubgd(Y?3d^BX:<\2eN]D+F[:=RIG>GB_dV#F/
M[JH8RIA=^Y64JOO=:?3WUB3GYVOAFRG.Va01E\0Z@7;-=MH8^B&Y+_57f/DdC:L
[fW;OAYRV&-\#1OOUPP.WcBfO,2V1WL,C8fe^\RO51IY4=BZ.2<;@@N2A;5BPL>0
PTBBTa_4C_\&RPU_2;F\?AX8b4&UO^(a4#^>Q7dV82I/N(:(g]>HQ0;1&OJP+IcO
C/Pc_4,^]d<)PfT;Fc(C8Sa5bH(@:7+(?7)I?>8a2R/;VCYMW?@bL7LE/L]\^6ZD
)Bd<cU4aQLcLG):]?0fM;ZTBXSQ-deBg8UL(Y;W]?g6^TKD-,7\O^W#GEOdd,g=/
7?_+Y-8RGY[Gf#(5&I(caVK_#9D\ZY6.56LO:>1D_;Dd>4=H0gJC3e?TFVZMTMA^
-)5f?S^1T@;D6=38_](MbX2-BAM0T@@;]eRT?5#fGJQ]g1;+>_Z6T7f+T[L5Xc.?
:@f&=(#aURVEg7\_>&&A;F5,DcdE)Bgf=CS56\9IJ1dD;F.E/OUcDYg]A,YZ/K-R
4CIfA4J5#I;a)DK1&SND<K>DE;]0X:<G12b=^HC+43S<Xf<BZ5YH3>f\)M<Z@+26
T?R]7D:>->4S<-#_eJ-QJEX>E\#,FDgFI[PMFB]S5SXIY9LXaEc)&5G)VCC]^K>V
?2#/32WA\VGFQ)B3AcSUDI-5<K84Ieg?]#M5)\J3,AG1a:cJ4fA@d7V9=Le&OQHD
J5F_0C8+-fQ(OZ1K@4WG7bXLc2aP4]X,L;&WMP_0d>KQM1<\W4Hb_b?6JLO9N3O@
HP<<]S.S>G.4;0RbObN_Df[U5=L(:6D+F9V[G#VW6,>3BHQP:1CS[_P:LUC>gOF3
5gXAb;YR/<=)G&2[4&F[BNa4[1Yd<8@@eW0UL>FEf#(Ya6V_5368@I5.VMc_MY6N
6IIQAIED793bdaM2N3GLG&1;S<4)aaAZW6DRg^.&3(8RS3:596=eMf2X4[75Bcd&
,fR[L&2JF]UB--Z1/8IHIN;\EMG&/^AdK;g:FYe-S;1</PNFa)a#K>HgAIgf@be0
9ED#-;Me1VH=B#[)<DF[DRFBfV[U<,M)+WQFV[QgfLR\=XZ@Z361RO9F-D9S?:,<
.94a-8\VGe<LLA#J-UTU9@@,XL\UI?,7b</35[eN<a.-Q+:LM:\]C)D;<JaH)OCS
P(b?&a4-4@aN2GSACd1](,/?/VJgA;3V?3)IdNJa-))EgER+cPO3gfY>V]b?Y(=H
fg7@QdRC7.^1Cc>X7Od3(,f@XO_2=Z87)@CC\#(HR@bRc_V1U+:?)egZ\I0R.<\Y
(GCf>a7GXU6ae3=+#SY236-<4&OWFT)Wff-5165_NK#:MU@KW.M@G8QR^G6I9:47
]Jc4VV7XG;VX-#/Q8KCT<\BfXHZ=K?..GU43W]9A=HbR75ACE]&]_)/KPX/g;2GQ
:Y8TLgDR[a2D(.Y+d0(=,9&E,RKY14>f[:WN.O<6/#0\eW-ZM-29bN7T5?-KOX-3
8=:_G,H(URA/2(/A0I_BMWP6gVY@<AJ-5NL^+P3d?43ZEX(WR&UU-M))AX/ZX6-O
G3S#IVTgJBC<H8(I]0=K2d]EK\UG?F6A=U3eN/<J]AG1)GfK]KE,(UM4GdI9Ha2D
L.Y0Bd[U=9=M._QXF:g]6?HX=KGR@D30_\YO1#20][./-b59D>N&NeS[.?Tc1<X+
,DYdcCYD9/=50cD3Ng)N#?DQ?]3UH<SW97]KK@QK_,:9fI>C:e8S=S/8WB&OWJF?
.:fR[<2U,H)HNJb72NR,2bOBC^:eYF45,+8JJUQRW]/54Y.)^f>3:a3:JD(FT/64
XI8R)I)RR)8<Z5YBcEZgZ=3D&dJ(PL>+_C/aS\^e=9EA]cAd8U768<2T2Cb?W6,V
Y6@1/>0FUH;CeZ)NBY,PHJeJ#VC(Q\9@>/5BX3[f727BI5c8C749V(&@,H?aEX2c
@&,O/1f><2X,R<W5MI8^LYK=]g-I:IaXg7<F-:2+5]ZNNEb8I38BaQY-DVRK2eeA
OXF[NYGf9OD(Y7@cH9\aE[\L#WA:A_9(1>LII]#;YQD<S(H\U\CWPb=0Zd@IDC,d
HVQ2KX1X\075^]=M9,6QC#&)eI@#K+0>G^,-)\=\DQaD?(K-9\Bf\K)_):))De5[
50CH/27[K__D/WXC^SI1e06FbN[RO^a3NH&.I.=Y=[EYeM:VMNM@=XN)W<)JJ4OB
L&SHZ^2ILca:&H0:G)_ZUc6F3$
`endprotected


`endif
