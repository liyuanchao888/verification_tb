
`ifndef GUARD_SVT_AHB_SLAVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_slave_monitor;
typedef class svt_ahb_slave;
`ifdef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_slave_group;
`else
typedef class svt_ahb_slave_agent;
`endif

`define SVT_AHB_SLAVE_COMMON_SETUP_REBUILD_XACT(curr_xact,hmaster) \
  svt_ahb_slave_transaction new_xact = new(); \
  rebuild_tracking_xact[hmaster] = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact[hmaster].is_trace_enabled = 1; \
  rebuild_tracking_xact[hmaster].store_trace(curr_xact); \
  curr_xact = new_xact;

class svt_ahb_slave_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                            type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_slave_monitor slave_monitor;

  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to slave common parameterized with slave monitor, slave transaction.
  // For UVM, it is available in the base class ahb_common.  
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_slave_monitor, svt_ahb_slave_transaction) item_observed_port;
`endif


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Slave VIP modport */
  protected MONITOR_MP monitor_mp;
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_slave_configuration cfg;

  /** Reference to the active beat transaction */
  protected svt_ahb_slave_transaction active_xact;

  /** Reference to the current active transaction */
  protected svt_ahb_slave_transaction tracking_xact;

  /** Current beat number */
  protected int current_beat = 0;

  /** Array of current active split/retry/ebt transactions */
  protected svt_ahb_slave_transaction rebuild_tracking_xact[`SVT_AHB_MAX_NUM_MASTERS];

  /** Reference to the current master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] current_hmaster;

  /** Reference to the current retry master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] retry_hmaster;

  /**
   * Current and previus value of HREADY driven by the slave.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit current_hready;
  protected bit previous_hready;

  /**
   * Current hready_in signal value
   */
  protected bit current_hready_in;

  /**
   * Used to track previous burst_type for error detection.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected svt_ahb_transaction::burst_type_enum previous_burst_type;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit active_tracking_xact = 0;

  /**
   * Keep track of number of transactions since last reset.
   */
  protected int transaction_count = 0;
    
  /** To track if the hunalign value is changed in middle of a transfer */
  bit initial_hunalign_value;

  /**
   * Keep track of the addresses seen on the HADDR bus; Used for protocol checking.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] previous_addr;

  /**
   * Keep track of the HTRANS; Used for protocol checking.
   */
  protected svt_ahb_transaction::trans_type_enum previous_trans_type;

  /**
   * Flag indicating if we are just comming out of reset.
   */
  protected bit first_xact_after_reset = 1;

  /**
   * Event used to trigger passive monitor signaling that a new beat has
   * been detcted.
   */
  protected event new_active_xact;
  
  /**
   * Event used for handshaking between common and passive common to
   * inidicate common code that current_hready has been updated by the
   * passive common.
   */
  protected event sampled_current_hready;
  
  protected bit   wait_for_passive_common = 0;

  /**
   * Flag indicating if this is an active or passive component.
   */
  protected bit passive_mode = 0;

  /**
   * Indicate the last transaction start time.
   */
  protected time last_xact_start_time;

  /** 
   * Flag that indicates if hready is sampled for the first time.
   * This helps to figure out if sampled_current_hready is getting
   * unblocked multiple times in a given clock. <br>
   * Used in passive mode.
   */
  protected bit is_hready_first_sampling = 1;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked previously. <br>
   * Used in passive mode.
   */
  protected realtime prev_hready_sample_time = 0; 

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked currently. <br>
   * Used in passive mode.
   */
  protected realtime curr_hready_sample_time = 0;

  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;
  
`ifdef SVT_VMM_TECHNOLOGY  
  /** This is required for VMM where monitor needs to know when the driver is
   *  ready to drive next transaction.
   *  This comes into picture only in active mode, however, the slave monitor
   *  has a handle to slave_common. So this member is added here.
   */
  event          beat_level_transaction_done;
`endif
  
  //vcs_lic_vip_protect
    `protected
(6E57D[WJ_#M<C+Y/X\<2Q=O3bg3LDX7;BJgFR9/6+[Y^:G_c4Q>5(^OYLOB/a7W
L2+HE]PF>fTc>Sa[09&)5-5N\B#TPN)INHg,]T_;d+1L(O69)9DRQ7a14/fOI&.T
-PYYJ\0;-VDA1PACANYERG3e9+W-M^>/+8fe=a(K2/T#0/[acL[<R5W8:_JB(LGB
#3dD4N2^.W1RDCTSLMS56W_W-.3;6D(5D/>)=aM/.8g\fX/]AQI_A\31da0JO3S6
2:BO4D?EJC>QFcC)(8MAY&&=#N?#V3<60:+.()Jb8U=6.@.c96d/#YPM_GPV&8Z7
L#aDNb,--3/AN)S/27,KNJ.2DC\>GK7C5\W(&<cADH.HTN=bGE?I2c7;Af^Q4[Xg
_W9[[@N[94@H-5WFJg(RI?V4=AW:08]3)G]FD[eY&QPe-a[\:+DUd]YP-:BD2K3K
KO4Ge,X.#L4>3d)RRD:98)+e/R=3_(2C@=?Z5A)QPBG==-0_U^<d4[gN:XaYAdCU
I2bZOg001&)=ebQ2TTd(gGbee;@Z13^Bg,.?TeA3\(d\3@,/S;4)a[ZZX#A6GgJf
IbG]\YcS1\4bZJOI./YEV&.#CZWA^7L8bR;<,;WCIF++Y8BKH_SC\K]e)XZX>R7_
E].9=\R7CP&5XG<3D_b;f;+(;C8d2\cc]gHAa=\A;4NSaPQ;Lg[UJ&WO1,_5H341
RZZX5VZeO/V,O2NZUc_X&3MfHEBZ3>18\R[D9C^I0QGUc,E^M9N8&3HCDII]O@(&
g9?1&P7(3;J65CW\>-L][NZg9Y[f3g4b]8LDM2d=I_#=I:ZJ#-QDJ?HCL$
`endprotected

  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();
  
  /** Monitor the signals which signify a new request */
  extern virtual task sample_common_phase_signals();

  /** Returns a partially completed transaction with request information */
  extern virtual task wait_for_request(output svt_ahb_slave_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_slave_transaction xact);

  /** Monitor the end of transactions to drive the observed port */
  extern virtual task complete_transaction(bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] hmaster);

  /** Checks to see if a new address phase has been started. */
  extern task check_address_phase();

  /** Writes data into a slave memory */
  extern virtual task write_data_to_mem(svt_ahb_slave_transaction xact);

  /** Virtual task to drive hrdata when busy is seen */
  extern virtual task  drive_hrdata_during_busy();

  //***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
`protected
c)+MbCR3SJN(L_P9TfRK0d\Q7L),f0]cMVBI01:X9#^.N-cbFS6K))3),=0T1_+G
30^5-,UWF/=\c[[I(b+f[M^-A]SBPGKHf<)-SQG]BUTE-G:KHgSWE_dU/4OPBOe;
0-DGLJ;5KIBSO9AF6M_4/7[-/?2=.V4d^X?TeKR46<0TO2@;^_Lg<IN)7M=\MKd+
g@LbO5)MKQX018&Ea2E;944.GP(P;c95D-3bbF:S7/b(g(Z5a\T&U1/3N8UdA:aG
8Od]8g\dE;+G>/X2-G5@^aaJ<_F:4K+.QC^1V@d#@BSH.MNI\-/J?1SF;BcAadD4
dQ,>L4TLP/#5@[ERb=3D7S#=<0B--+c)eRFE0?KdKY2I(@GP82>Vb]RJ@EEa^,N+
d?RD\L-gO?a[aLXNUUB^9E25>^Q0G+13OWcY>Q2:B45[N).:=M]aEe)69H9gN:-g
-,V&1=WM7LMP9WafUbDUO.^R@EC.M2#K8<fKY[]0<J[g./1_MOG^G&Kf?[7?SV;P
+aVDB^[e7F:AOB.1OaC21-=;Ec/a)-.H=A]M.8@OdC8CAGc??46>dE@aPJ10A&?D
:[&L#DZILJ>9^Ia,=:+>3FYH:f#_Q&0>-QeOgS3c^0=Mc(&-)M01+M;+)(Z6,Q9Z
34^9F8V<,a7ENYbOF2-L^86C;eR<3A//c>_5N)9c[K1aaY/&C(IIN[DU3OLA5ec;
P#?WDFU_G[A(e(>B<-&5TM483IAacT@<bJ>(UQR6G[BBUc[&3+]f(6Ec=>JBWD4(
b3\OG)86^R5SgL;.]K,\8<IE5KY^]c3b;+W+V(G+F:XH3JbS+50D8U;KT[Pg/,4?
d=cA[5E+K=<VbTePMED3<ec@Z,gd/@C60[_)cW#Y@(Y9UC)KO>bG.D1bM5PD;G=/
^8Qb^0=?\XHUN/a<YR7)If):5Y+)b2-N^T)]bLR\TNb?(LJ:(^>3/5O,(d<5#W9#
_b&.KdAPIgW#RfZDb.>7e06[)_YV?]@I5CL@=e.3.[7F(/DXFHR4VbNCEJ^4Na3a
12d)[&UXfAd;(2gPKeF1E+(<^L?KMFITLOVD,M&WbX@ZHf.[/8CUOa3bN0G&#]B=
.OB]D]A4F5XH#5K_P<4PL6\E?80.T)c+M1&&PLMXE.)[bBaBRJ@d^,XEDVC>@6&8
K+G:BA_eXP9A9<YcU&B-W27OSA#3B\&<S-7[P.:I6#\ebRJ6bT<@UUI9^9NDKX4U
J_b8f8WY<H;):3cV@PZ4HVTWF1S+BH(I/^1@QNI?CFSC(0EOIL#S7.C@<W1?UD(Q
g9b/e>O@3ZJX+\aP:b,S7;1=.dY-@4dM;23QefcUU23CZ)25D.fGcKU5I&8W[E2K
T@)CaaKQP4#S8^LW94R;::9aDN=:>-V]4^c5CQ6?OcAY6>:cO2)B<LAG:M==O;3A
XD;JC=f(:e4LP0b3G##ZYZO4gcGLHWAON0.U-G;#LBKQB&8OTWG+0PJI[A1S&gBX
SL778KM=WX(:>bOLER.<G&f.4(Ud(&&+Ece<(Wg3NZ37=EVJ(>>0+FG#-XbIDA<B
(-6g=(BULFAIM\=//c//CC,78;V_>30=SF]#M9+]H1MATe9UM;3JCB;U.+2dY+WT
CY<J-8+MOWQRM1?=7H.L4?9WO;EId,O+BfS;_4I;L_]AD$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
<53&K>eOEJ?WJfM(cUDXVL&3cg.E9A3O2AFVf,<YQK#dTN]+//?>6(Y,F1GHIa,K
MV.9=.;L.^>6Dg79-e-_XfOJ/IP6LXfd_9Z-IS-8@L62c=67^RaJT^PCY>HJ_]eJ
-&LVb+G333>Q#I5)IUKA^.)cT)63_2K</Q,003)UYT]_K4HRBK^#@a.#c9C(H60d
5HXJU\^H_FME.^IJB<2ZU4-^?E/5(U/R<b>:W>B1cbSACbON5J_Ya2U;0\84\J]R
ZaM,>X[PV5eAaWZ.D^,2_^=f^D9;))WSW_4D:Xb4J<Q)JD5[=]3Y4D1<NK8+aK.4
Y=^0-@:)geC&9\,RXFN67_KSfK/+U5_]4T\]b8V0_Q:S_&Kc+ggFI;#7P&6.B9<g
TJHIO3DfP[V;/(@HVL+1C;e:6(09B_+]I\<FV9YLZJ.#4Y(0)=X>2Z_?1QIRW-S9
(0WG\1+<<6]bL2Y_^-gGN0S2T4S?B[BD)0Ta@Y.&d\e(;-;@P8#-J=eCUB8e^+a0
a:V9LQH]NO&1FQV)7@MLEc6X>)2&CIM9];.2:OPX-_PN8S\5Tg3:V9d>)_K3TZS4
b-6W&XV\#QT^LY6.f[W\-X#4G2YVd7ZP72-1V-Q.QOP<ZX<>)6gIBMSfT5ZUK/1A
3WA1V,+PZDDJ_([WHY,DBJRd.Z:>/0dOZ^9:D:Gf==1a;5_Z.cM#^8>HU.&Z_G=Y
\eUZdGOgTccIJgL&-f6SNUff@69N&A7)MD61Cd-A@E0Le=V&23Vd-aL,7A6J@5a,
NFST>S>C)^V4;?W3@P6=8QRE3#3.+>1.SMR\K5SDfUaJ\V5WJ.S^F?7U]FSYc[EF
a[MGFAVGXVbLde4PCX\1g:Tb8;_V?9WN>:F9J8:Oe8QIeR[>-_S/#1<VQbc:Ef5@
+_C&^d)d\@:V#L-I9-GKf=77J\8VT3IMUGQ+Y#O[af(d@2:KKPKQE]Q3C8S^cFWT
CWfL[#B\aGTb90,.VKIgf.2XUYLC5H(@LH3,,D;<YD^aV@a=^Y4dD&<8#K^X>QG1
a?]Sfe#_VF(2GMD;[?CBK#c)&1d[#Z)E>R7[A^U[]aM=MGJ]@d3_MN@>):c(8ffd
R=L1LZAT<KXdad/f=R1Q&F[8W>bC[TE5RV8/Oae_Xf0cE7<SHC@T6E\X0@2<,9E?
5\V[R]S+H3=GO,a8\O1?T_Ab=GRA^NcSWG9ZXcfOgaYIF=BZ7@@<M5B4=/#1/PI0
>?:b(;?J^BJ<R02413IM\+Z3PPcHPMaba^FMFK=QE&E<?(KRTD0f8LJT:J>aQ[SD
+1I?()<_88DV+BF^D=>I3I5KGO8aNKX(JZ95c_)C8GQP)4^5-EQgRc\)4DB=:H[&
C^f<g+&C4G,P2+cDNO<^RaZg#I(69/\<U[0&2)]R54KYMWMW_@)GS<@#QXY\f[V0
-36)HX19.PRWcCRB2EMWLQA[:cMdXMD7NC/YF_J:OadG>]bV(c17/6Z0:I)W<9L(
G&g+,^C>,W[W]JL1dRDeQ;bIA,Gb3,:JH#>IC9K-1:@G:,cY<gFa-PU,Rd\0<_A)
P)>23674,8/T93e,V)>G)f5\IQDYC+;&cDV\O8E<T4EDOB3N[/B^bdY@NdWVDfT.
H^caeZV@EF3B^HH15>_LKcbA#92>aeg-IHCSU<7\LV=V>dCV5&BFU#_BF0N9I<fd
D)IYV\6c_PeM7G.=[HF39Jg&33#\>=2&+LKc4H]^=@>:CGK_.[<44QGET[c#J\f9
>,-Ed\#A;RKgL919+B8<KGYY-c;K24RA6>S<81JA2^5OJV]:5G5Xf]3c0]R98<60
Y-MD5<c?,L5\+bY)aS14e>:M1PEEY#MO&##)+==,C=:L1TW4-TV=IT)#6/IX]D1C
XNP\L:G^d\f5B3aV3S#VHB?_#b,<BJMH=<?6#4#0=[;WN?G+d\d.d9AR)TF>S/?^
@R]7BV:;5c7:11P8P)3=7GLY:-AM5.7Z@PXI_cQ3DUUR9#B>bM[99YaS58-,+CE@
UFQ,#))N49@#)]BCSfJUc<M:@11&0IKXbMOAR-B-D\QU5fN^1[X-8,YSf/<I\[9U
F<7>1VfS5^H)(/._56]e5?HBd.G1_gcF(P2GJU-@AG2KT+D(a9Ya6eG=D>[PQX[b
:L;@DA8eZJ[GM3Zb:Qc0fJ5O8-U015P1.8TRAEG=].WgT3H?WT,Y;M_F70Y/;T(K
?ed@JRSIcQ(NWe2cKg[D5QZJf(-(XXHPg3/2X]+&VFgMO4Qdc67b(MN7EgQA1.MN
ZV>3<cKaC=8;,[I2L8.K[bZVTDO3IaHG\a?T,9W<LZd^J(PgadbMNI]eXa7KSWEf
IaJ-\T2MW&<R03(IM>+>,,f&8aN;;<W6V7SN^7[4^B>^+@9@>/]W]c.SF>>#-YTa
<T]TT3IHMb>;&4&RV&MKHbT\L>1#H105H5Xd-J/?UB_KCCQDG9B:^+2.g&PASI4S
G,5HeYT>SbcOd9B/]#N[-\L1VgMW_CbY>Q?)-.8W31:TdZE_f7?I6MKW<\Pb3#1Z
[1=U?R@G5TE,OdSQ)UVBUIB-4MWJ8PD<E2TTY<<NN;_V3WFb.,IXLA[<2E=:J[&b
3?FM2\#R>B\:egXb_R&Ea-&#L&WFJ4NK^cEB4N,7SF=NHcQH<Q?I3H-RTD_=AJbR
841]&UK#R6WSG_(FS4eH[=,bAUc<L3F[^A0gcfcDN,Fa^DQ:@-aL_+BZ9a0gHg\#
)AOL99e<MfgVI2^K;HCGEP?Xd(>d3QULUN,1HTD49B1abR[[@2E.8+2,c#ZR8DWf
b(=d,LaKYS>,P.(EURF47EUV_S9JdMf72L56&D;[ODG1aC3LY1)PP9&:#<&/0f0A
HJDPX_1,9^;TH^V5O+>_H0/R<#83/<@Ve_994_,)Z)T_dL6b;C-R/UYNJc<SQ-gV
RQ(^A<4WCJMN8c9[&L[/#4/f]P<Z]ITNE1\YFg.RZ5HPPeOg9#@EIZEKF1^:<#F7
Y;(g>APY:cY)&g@N@\Eb6]Z0^[IaJW2,#F<56)J.1+C#_3+EX6b@14[3fS>^WF9E
\R_>_[>\;b>69U[K;X7FRY&FX-09ZgW54+IID\fP9BNb\Xb0<9_UW@RbC(3G5+U;
CTd8W>\COXccX3=c[X=GKXKbAV1V:Fab1YUHR.F^N\:@O+TGd;:Fg?BEJcN5f/;[
H\#M(Mc)R9P^\]@519V0QB\VUAY>6DY0@>S:I^7FP0>?3,(&@=4R80R)9P_=C=eW
4?;/Rb&b#O[bS=[Z;d,C\]7P=2MDdc.^0LdO/R1c#Db_V/BRRK@--CL?<Q3a&0S+
-7]1Y>)/W22PS3<dDW[B-VRcL-G8N5-=,eG?V@)&H^EQa#^]^U;CJMOE.]I\[-G]
)V>MCSO6>6YLUE+&Q,M]EN#D(QUB=d?cX0#.PQ3[8<^OSM-KN:;]FSRY+>gd.D-:
1ZUN4eD_US,DVO9L<Q^g><d(?K>f?ZU8L8gZ9fMdE)cR.[f15@GB,dL_JeS8SJFU
MB4AMMM/Ceb[4Xa,BA6?fY=G8;EPF4VZC](c>:c9B,\aI2:IRQdGZGVNTX+cYXTH
3R^S9A?E(_)IMa2fb@]U;7O92NZEe#>7c)1_S^/[M,1E/UV,RP^K;7A)PU:HMET2
[=8JC8157Sca-.R69T,YU[#1>5bMfDL_/U(N/HKF,&[?BEQV2)U]Mc\LDPR_<)6)
[:^Xd?W,7PJZg3@0+5QPBa,^WWK.8Z-A]XY?K4Y3?T>Z4Y\R-BH]6^QZ3,7H;Be>
,1KMSWP+QY0TV;ed<aKMXWWIXKKRJO<6#^c=e0M90f[C:ed#0;1,Vb0H\6efS,R.
8\DX,7U/ASUVQT[Y@K1@f/f#SbU01HIWF<1fCe8Q6BF.=4aWM6DaQf82Xg#dbde)
K6]//P>L[8:+9QQW]7^.6dB5MGE@fN99HLZUcQ#X:1@23N[7GZ8B\_3P><VgFMg,
G/O,-#)(>,S_d27ANO<K)WD+HB^[eNe[/UKRTBXGV5NBId^=bC/fDbQZDBfAc\a,
4MfT73G(Jg:[Y+_.7X\@LVLfSdOBTER1;B4COIBe1.4.eYN9X99(MPKJA?115_^7
E]+f9]L5e?F)51e5)JT@VFR/G4\SG)4a@a^[b)0+OT2SZ0Z_ETXOMA0A?[Q6=gUZ
W6H4?=\f@CbfYRFHXQ[;;5Y63#9ERe29_8]TZcg8c:\LMLW3A;=f]5[MCJb:UN2<
M70f:M?Y=fOKQTH=&QWYJ]3QJQ#;IK^WY3-,PT/@BHGG(MCE\Y#14KeM6__/^L9P
D\/Q-2&P=+;0A[Z:/NJaee4:)2H33b=RHKK]VbKYQ#g4)0K;bDZbdC^GR6WX=/<K
1\D-f8e5LeN&INEADa4BaQaaa(L76I0VY&eSDSe^\gKg8R^>+C,_E]QVb;TY2,1/
OGFS@N^9F]3Kd;1\[4\9\T#DLeG-B2#d^T-<ODOfWa(4DA6AN)(d]6Ec?YFCLABg
F0-DN.MTROQV@fJZ7-g1EME/3RcN;MeS,)&dff48Z&cBb>D@:G.WHV<&[<D?2649
BK6D6W2X(?@.V+O:/=D7+UG)MUO0bAd.X^T/A6<GC@fa:F+5OT&ZVZ-V<9#M_QdZ
DfZTDDf_6BAO)c>1c@.A]aF/<fQS>4f-2gZe790cG0B+.e[+f==I\<-SK]a_7UUO
a5WFJO9^ZY(C=YaLSNReN4RO.\T8V@+L09Ng\:KT+eKe0W]N+@Z,UUP/g#Q\PV8/
eH^VUI8R1S_Q,2SPOa=ILM9HR&FMY9^b<:?7K7E]_HX?f1]U]@84ePE>8=V5EU/(
;WO-^@B<BJOM),:c^.W-_M&fF[5e;=@;0B-K]:#V_A4\ZH^]Y<+aK=J@W\SS1J3\
GW;[K+JR&d09C^[7C^=#5NOU&_&J=.8LKE[-74I=QSeLYVLCG<6T:;:LE8I-V=\/
)^@21<5N(ZTR[b8g5>RE)A<8N@O_4UO9D27-N/>-d=g9L?J(BNEFVQ@\&BYf.8>3
SUOCLdB;<PUD:=O]6fTO/,I-OdbFZ<a9e8L?I8@HbZO5a;XAgMOXGZCRPcU@4\gB
e,=EWf(5F5K[4O]17N8fC9G1U<ZIG)K&[b.1COc+L[T1b^ZD/4=W>28I.PK)f&/c
;_KU596UU3K1fccW(@-_O57=aZP=9L,8\ZI-T7+KK77NN<I>1Lb^UeY^;:d=^UNc
/UaRS8/aU6QTRYAB,3GC#aJfSURIb?O)-4D58U&4bGP,(K09@+8\gCX89J3MT1,U
g8III(+M,&-WE.Of@I2DeK9c&W#XE572R[(@;[9@\<IeAP?\Y<IeD(CX]_38[A^V
Jad;FGM@Z7.9YQ7WaZ-JU]#cHbPI]f80<<S01@HN[b_2bJd5HVJ/1HZ)&N=[801+
;C\N(8/GXEM4CKHHMRH)#LHQ2N[RXC96&?XLO:b/3NQ7H)O60<IXO>8[96?D:/L7
FFL1ZR=7JVaV,[2Z657ZKE@&DII2]OQ7[NgGP8OF=-9U)&=XNd4UD\-gfE@69GF=
MbV=R7(L):XILO(=QX?dSI?&fGCN92S381Ma^Z.0&.6K_KYX0SB8#NQ4d@#[3CM<
IL(W0b#?7YC-3G^f<=CQQd_QI3KD8E_P@XGbR.UACHGFcSZRQ-8666<b@7KCSb-E
1SfWOc541X7P5d\L9#]J_)U)51A/\U]TYFCaQFeG.&a+B/J7PP#dgQG(XM]<Z7\Y
)7T[ef.X\0[;T#;M+RYGX1Y15-_.8DO:,b-CU[JV=e)=1KX2:daJf81IE4(dV#RC
4@Fe5S8@:#6[E3C8LM=:F=+X5O(KU/WR/6K?AVYK&1b<)2MR=L+;IZML.NNe;^fb
,OMfYSMJN\H[PWIHSA.V:=d]NMUc]&I]E4PK1eIJ(YCCWIg3_?>VQT3gRcKgL6eH
?g\X+;d(TES\6)#@YBR:>FOP8()&MP6GY)=HZ>6NU3Z(@U.P=(&J]/Oe=UUcfae?
<W#Uc/=T\Ga/d.3aLZFPc3ZcKI&4@N.LVA=N-D49T[XCMY&<W21__5@V]-cL&@G=
Y:XKE;@5IJ51fPWEJ\;Q5fCEC^[Z,g6O,5Y168aQ3LCQ7N^YS:23W^LYJWT/06g(
PWXCL=8S&Z_.#H?I-W>T&)BIJCND(6@XW,DN&4C-)@4/O\\9fd=gd_;@FU<3;M/C
d\f;BOK-JURcG37Kb@B6I9)<YH5;\fQ-9A40SPX,&dFEQL5Cf,CD3H0.AgMPOS=W
2E]Z<f2_@-NK_O0994;C39@8(\&&(6\BV@-98>Z8#_T_IZeZ&@c7AY^-bEM]<Vg.
57K3d36Bg:[&Y.80D7QBV7Ka5Ae-T9cVTUA=>H=;Zbd;QI[RZfFec4+VVWD@fN1,
<H=#e8YX=/Q)=ge3GA.?Yd>Q-9BYKf&?85]H5:59F5ba^TZP]C]NQ/@AWAV.fG&&
4M6c;#+XV4V4VGaKBW[Ye997C<CSE:7eFG5L7LO\9V5Y>A;^SbPga&]GNbN\EeU7
(e(D>8,ZJa<)8g).M:#4aX;Jf.9gZ@#+b1BeV<3:>;NCJ-cBIG+N2eOa<f&fT27D
b0&^SI_cMVL3Q1d3HR]2-g49K,>bOg#FOdfJdIe6@_f&LXL(MLdXV,<1M2AEJ6;K
gfA7L8._@[:-<94D,a=KFT1cFRRB&UUNe0ffK\CQ1+),b@/JVP>:O<Ef5<S-,G./
^Z1bF)eGCRR)2L9&<3XV+XP/(;Y\\M0Kd.EaEg:YP@S=2_]KDQeAZ?B2#<?;SgI@
T5B#62#-\91A?^S8>9ZQ6J0D6eI;M2&8;A^SZSCAb8H[:c2,QB[:d\:Oa-O0,Id/
@gW=P<QEX^fFZbMg^1dFWg.C?IXN;dO1TA9/S7EJ81<A0F(>QT/a[ZEE7PgJE=\2
97S:eL6\BbT[&MK\I<?:U@(b)AME]JCBY\fRL\FK7_5]#:^K)^E^^KLZDe>D-Q6C
KR()<31L79&F/(KVbTS(3VQaDY#?K6X4SfcDHP)ZX/3(]E?3F@MMR-90=SX<:d:E
XNe[eF5;M[R\dJY4NVUcLQU.PY@6[UGF\DACFQ[19X7/XBI>&M,d?\QMU9ND(5S^
&PF4,MdT7:Q0H^EK)H]T8Y#Q<D,F\@LEK5Y#L_Y.;UX>+A/@C\D6T[S2O\]agLBH
T#OgDV)fQ(+dO>a-HZW1EL+=(?AD\DA1ZA6M:6J_SXP?fGfE=CTOS-<:ffW/HFH1
5L[^+5(UO3g7[-ba2POY&dVgY\bU5_PAI-^&&^#W>7eX^?WXEgI;ZVO[5WTL?5-R
H_-SeM0-Q5)-6-<^(C5KH2^_1O4H)M0g.#L-YfRM;GIHK,P_6T1JV[7E7>+Sfcb;
/\ML?bO8LU-15J5FV<G9:F_bKHea5<d-&g(-Ad:X9(>B:N^Xf-DXTE^ZaXS0AS@S
I.E=XOI##6ZI[O_^J)[M(S>eID2-(I:Z0aCR(LW:->6^?4M.CD?ZC6(H;A?8f6e-
d7fITO(1BDE=HIa7aUa]-RFCEOTC^D(??DGE0S.^7aYPa067\3cDNeOb7<0MHd+L
=&OCeH1,>:>2WQ8#TJ&4/_0RX8e@<?4AQ28/K_+QRg(<]:GAPZR\A21Ga7UL\aYZ
EFPW+NG8TeD91f^gDf?5<^:]Hf9\.eQO(DSPX;C+d_a]=[&CCJORAGQf]?VSV2Qa
GMa_aHfY1\=3/TVgP[G#R+?]\&FT5M,Uf3]A1#FOW,TN4?VU^DA(T+)YR=I4OfLV
2-Qb=#5P&URL+;@KOc:V?F4<\V8YTOSe.K-<1]DVZ71R2N3>7KYdJeV,8J^Ne)[5
gKaX(Db3F[VG)HCENeX^Sf&.ZX].,&#K+-@H;c@ASgX8^N\5:76Z@5-1T/&GDfK(
A.=Z6L\V;5B25VeWFEW4;(J?7]75+.9(12C@eJPZ6@0>G,AV/HJfYT->gK7B0&g/
#B#f:cQ@V5aA@9[S9a6F3MFB-])Z340f#GO3TK=B5\)_g3K\gcf/#KDF(RJgM);J
0F82_ML_fA-(A]/GS7CRENQ1O+(4><W>d->-Gg4gS(gM+I]85c&];L8/;[ZJb>65
CIW5JFfJA4(bg>UcZ42a5aU<^3SDGIaS6SJX^IeeLII=cfX3?U(d5g2a5?KKc]^:
65/I706a0R<(Q;gg;L:22;6TI+KdLSd1<7FA)JW]FWO0.T6LFLAEf0#fa6(1dLMN
5YVFd=YK3V:,1>L+?^HRcc34__M[6R0,;P^g2A0OCY5-0T-YQRA5#e?(>X_[8T?7
A<J824:gT+D=[@XcK]0:Z89+eKE=_7;[\K0,RVVdAJT?<GX)(8[?JFS]?N6Jfc.\
)-LAc)JZ5+CgK(,Xe;0)WE]TOPaJP=fa<(QI5]YgK(,:1f22bWJ4fME(f>ZKfM,C
b05)7N,?3Rf^DHc:d.1MRZT?T(cB^/>&MHMD&Af&-;@Z68;-ad#B\WA0-]X^c)3b
/#A4bC,0V[[+I](98@R^YEF2F:85+M+8S(O:.RN^X&1GCb5d;P[(AcH&XA7MIT8e
I->Q?67,82bM86\=a)4Jb-^a9./077X1>[AJ.#2Ea9<BK[7J_._=g,bXY0b/:PDS
\UDZRJf0U^b;aSO:D+6a2L.27eOKA(WDBP6C]8>VFS.\VD3V\B@GCeW+\f;DU>Q^
Jb\RA-S?0fc<7(2NE83-baggHQKOIVR\+73V<CC>)dORU@W&VK(31R?OI^Q^T+K;
<O5KP@Y0.N52&Dd8.WJMRe8TCfA_5e\V6]6[?DgPbFKN1A<E:@Z-#A8+H)B;-Y.X
,-Y\VNe,A.;187108LOQ0PcQ9/)Zc:;Pg(0H_f;aE>f?^]dH/20FV:U=@c-@MAL8
SCeBW7FS7)6)S4AE=YDX.c6-<UX8MMCFRT0g>c/f\O\bL,XGW,H:V-5FZP:KE\D+
T/ege#7X\Y34&?Z:\M95:QW6-O]ReLa)7WGTQZQU1H8E\2\>E\Y++)f^Fe6(8Ng5
KMC;X=OUcFg2f4<O?Hc(Q)TXCe34XXI0bU_32HKH3#N^WF85_()WK.RN.aRddF0K
G[b#SF+-4a5aAC_S]8?WVb+W-S)a0Ab-Xd+/&(_F:Y_a&.7KB::]F[1c7A-3JD)\
ZEFb9).29-TLWJ[6]MP2Gg8[#)G0AZD..aT9C:A(F8@9@3PW169RBBc7QP&JXF^Y
C\LY=VVMNNJRf4^3R74T\RNN,5]9IZcLV&ed=bC>.)Q[/JJ;Bg3-W4@(C00_GX?f
IgFaU6R?-D?1=1d><>^1/A(Lb1C;B2A_\Q7g\T,-<0:(3)Medd_4MgODbVRe]Ecd
C4S-2\)gLEd75NgP>LFU6a4R\]N8WH=Q5?XWgBTaTc]S;K^C;ZN+7]@#fcHIF32_
3-(JfJ];.ZC>M?AYAS?K,g(FB))/>SEA7g]+F:->QHHgVa9g;[2O_NF)01[V;W_,
1_(@,d(,I8]&URP7WVaO00:HE<XJ]EbXG12)Fd@,(aM0JPD3QeL[)AN9\dQ)#O1I
dC#gbW8,#;YU^@3ER=#&GZQB38e3TLX\MQa[;Pf5K^f;Q@#P<fA44DbYcS<=5-00
&W2b1F;P^@=eLeH;PgRG0-KS>X<_7KG,1c[?b>&&[B,,HOIX&RHAN2Z0HZ;BNLLg
F]g_3;CfDC>Q]CD=QQQ1U^P#K3OJ5SR^V^+28VT_>]bfE3#E3ANb3K,U_1CE.;PZ
J>5Ja],:-?IL4g?Q99U<eJP#2$
`endprotected

`protected
=4BYB2:+H+F91^_M>NC@1dFVT(_IZGg:YK/Y3,g[YM8N6FSMcGL35)Hb5^.<96+Y
)0^M#J#6;1>d?S1@Ag9]Q9FV7$
`endprotected

//vcs_lic_vip_protect
  `protected
?D3-EUR>T34U]E/TY8UX>.c;P=cf#?4Gg8&L)M8N+=CWCJU<(O#_7(V:IcfgQR+a
GUc02/bJa:CT7@OA8YAb2[&KOF>PAVIe;JA8:K/MAQUF0eX^5Z+--e[O7_a],PL.
O:0D3W80/#YPQLMYg@5Bc7db<)3F-PQWB>;W48C[-4:d#8U4_H1a<:S_8PK8#2K&
LQ>d#6,:L\5M=ZG+:39RfA3M?NJUZ=_B]GL8)MB<JeJE;:ISV2]3^Ff-g&WH)JC0
H,N#DF(D5@0CL:#R?T1d30TCQ/08e57(A=&KM<<FU)HFO;a&&ME<238&7ScUKd^:
EVMaccc)OPAWWXSc>G(9:^:8MgJc.f7ER7,;0^@E@f&4_^,284?bg;I1)LD@,2OL
]-6Ief43H_(J7_OHAQ&+cMRf]0)IA[gTb]S/AP>8LAK,WAZC^ReAS8dRA1P1(-9-
451@,\=?,K#\FfT.GF329.J#C.NZ:1WF[:JOUQ-^3^-0b>B?aNRA+T8W5E:;5BW?
5Q<6(9AE#]&#K\^&^F#8UHP:2Ve1D,1OUE#UVJD>G?RPL\<S2WPZR:74+6+=9DHL
34;NLbUUH+^8?LBNb[QA]F2V69/_E1;Vbf:[=JK@PV1U9A2V5#71eVd1NQ7(-UHU
Od+IEB=fGJ]2,/g/<2J5aE9QLLANI@:aBKM(4XP<5-:3(^>?.=2N+M5P[QId;61g
,3I6gU4CAZ\_9&@MFKYZFeF06_AC-#/_V_/6_LCb;7N_6@5CY67JM)^N9A&,d5+4
1YU+8g+73L4FCS<KTYA-,55#_d\cgfdX)4R/+1PYB_U.PNDZc1PdN0aWW[&P,Jad
26776+QY.S@H<72KZCZ5Xf25PS7e(QCZ(CZ:F.C7dfK(FH:QW0BJ.4\7@90>cV.L
F9?E@1Z8J.//_Wd@B0IM#+>VZ>:5P]aM2>XJWedL>=@[FJ3#69:WT6[RE2>]]f1D
/+#/;GT2;^TUO[Dc3G=/+Z[25TL#UTTPDQZ^IP7TNI4AGDDXaHU?NR<J1Q8?E,c>
SE0.)RVB^TU(QHdPW-B3;@]2<[=YLWUK=aTc,^(DD75;](U)XcL8Lg?bc5eKXQb?
OML+1:?b4CE;QRYX=b?,5O)Y)A?AW43X><cWRPF3F#I.H]6N[=WbUe&f&:W@@0M1
9f2L;4a8U=f5J[.OD[?1Fc];BFgOQZ/gL9ScfCJ\6d>V?HZ>RVG-dDccJI9SNDR?
FHBR3IC(e.7+CJc9ZeXg#[0[^\^[IJEK5RK0J;;(VD7DJ9LJcXE<3LB.2[gTEG9\
32L7P]-VgE\NPN&(U^XEe]FdFB(RcY<;,Q=H7cN[+=LgLXWZL9?5e+KXgG7@D)W4
a(d[GKg]&I<&[ED+c;S94<f+];=K^P/fQS,IW8TXV,H?N/_Fa/GBMU@:F>)gfQB4
VUX\4^e0;FZ<PTUQ7L56)=f&2:[e[d4EVW<9Z(WJBG?JKZfe_/BMW5IV;P&+W;G(
9C[)#O[/b<W@S3eIJ6C_=b=M>AR^D1:Y4D66[33<??AIW++G;JOg?c00-MZ>X@L.
ROF(B@gb\^GAA-dA>3\IXLBTdGZZD[f11MW-[[VD51G,))cd;+19[fPQOI>FLPJQ
O14Cc0ZBEQ]MEFW:^TIQ[_9Qa_ffF-84M.VaE,fN\2_6TN4)Z0DNabd8ELNXgTE>
_9RM.aEA9A/NMY5KC3(_9QKNXQa</>>XO&cLGNIg#M)-=_?#LY8G5OcO_<L.aAH3
/VB?eXGKS^aE68=1NDGJ:8Bdf.#-c##OD1aQbSI7^^^&H6;W.S?8:AQ8/Z_5D-+Y
@J;+5--9F1c788=.H.RBVBVJM0Z.WcRMX6)8a]C_G0MA4dK++dA/PL+<=).-XPO9
\0TDB2YO0=TPMD<P6?G?S^J13ZEKK=JT^c#cZ@?PO^B@Z:Z^B^+L)()=/MHc.5L^
(J5ST2P5],^W\YODOFD-Q7b)8+@gaX1e+P#Q/>]Eb2-27W&:f)1f?[9GaC-+<CU<
<[eaQJ:N.OU@]ZaQ<>WX>X?BeZR1FUKI->V12B\U3\V82b+G^_VREYWKJ7f0+V@F
[Y[4NX2,P..0Cb+PJS149Sg<:;&\b<>a?R]T1a,&Y/FH_^Y.R[Q2FOJ5\R/\_3]&
Xf#70&^(cP7TZVL#If<.[f45.]=184T-(=7dKKGXZRRL_D\AH-MI_gQSEJD_7KBH
&OYa&JNL0^=9?2<-N__ZQ+G+.Z,R]RN,LR45HR@G;+P.I6JK5,g)ZOe2(RUIICUV
<93SKD=)JKgN@bEF;BW>F;f\/UOR^bM/)7<[PW;PBL;M7]U^I;J_1ETEDW;dR040
/LU9L9^DcY=@XS;T8ZD@8J]aT5@,C6>;4IRAUPUE)b[TfQ2YST=P)eNM=3=,&U(I
]dN<TBA#7-&D@4<E&.WAbFK9N#ZXIe7[G1R]bE2d>d4#?^O24aWNSWRAKA):0UPH
:fVZeAJKEVH68H2H,>Ge<D\\L4RB(8KdF-EBIg8@)2?g;WDcfS&dK0T[])M/,XXX
#\.PNJVbfg\Ig3R>5L\?..N(Y(IJU=:GSG_Qe-4;.fg]TIc0V;L+H2]WMB@13^ID
cR&.578D?#gK7Qe2MUf<;@J8EOdQB-&GKWbG;_&OBA/&W6=eRF[D_\.FSTf&^R@?
Z8M9-I<_[W9EPKd4Mc6DIP=P@GP8=N6IPc-e(C20D4M?6[(T(12g4c4Q?e9@FZ7H
_9<,#0<7AM8c<b@Z-6,6ZQ)cIKgaV_b1a()P+1ZY_KS]GK:UJ8eaT=Sb&RN#_))/
1#I_E50^H_-f5+<<NeB@aYL5FKX6+fV6-cA)BR;3#N)?ES4:Od_DDJRJJ+(;WE9A
>BA)b[I@..C2G]7gGVaK=.KI24M-VVZ8,gEQZNg\G0JPNUGf\?dJ[>cCHg>1JFb2
2?5D8_-0L5N.ED[O<(U[@/4B-f5Y^eP00JeLNOOK+?,O_+R+T^8XOa=H;@^J,].L
M+cK_E1&?.?)I#d_e2A3a^PM)M,7EW<aV,cg+<_&9#V#T[e1O+8_V#S3MN1M0XKA
J<AX]?X45[7<O=970G>_<WgPEDc5\Jg;YG.DO^BC2F)<]f(7da?;dccZcJ_<UHLe
gOG1H&_/:7@;9QZI&LGdXKGKY.19_,_;c<3gMAg_Q[B82.caO?A(DFG071We1N>F
GOdXD_?^S[8aNA_b(bf.H#.LX+f7[4:DWE:><9^UYeW#1g-<&19C.-]Bb(@C;))>
7I6FDW>C9K2L(]3D.A7V=9JAQ/RZTKTQfL&)N<Z^P7S3C\<JMX5/3QQ=NedQQ_?M
[OEcD<8S9S8b8@EW70dbS==,g9>+#C^0OG9Oc#G??@fD9VAZ]S0&fg_:DJe-6NbM
8ZW4_9K22SFcS8MV\7f@0QI&1DY(ac?:((L,SMJdO[@Z3DaKXf-7:WOI[]^F3\YE
N>AZ0d5RJ+>Z&?V9BfY:D)e]54;;62D\Ib4IK>7>Q7:7RDb9XH:W4f@0#\HYI?/Y
\9MK;-)(XC+1aZ94O3QX7].4C<>6AXb9)+PgMebV/5M8??5HN1Pa5&B+/;,W_+WZ
[B_)ZV=Wg1;K&d?MC<<>d#Z#Q/_7PJH.\R7X@^I1WE1+PZ+@6<.LUE:K3WR,D1_;
[.C.)N?F=Jdff#]A-6=T-1DAINe5_:gW).IF011,=f@MX:W/VDH>^O[Y=2c^:YQc
[?D68<W:_aAf1/)#cUc]e5YgGe&<63Sg+8VdFIL&D6A&KcYc^>gDbeXc@6C_1@ET
=)(#[@<cA&aW21Oc=_#2g4MS1^#UBZg7^QO_KYMZf[GZ,#G1dQf757_.0a[>\Jg(
HgAF?##)/\c(_/+7+>6F/JUD=@5:7cSQS>KM[,W3>BG-61RR-gO(6LN4KX)L/QV&
GOG_^GST5A<5_3RedbOW?4b\10LbgF^_e;&)Y.B=5^C3TdeReTGUZ_C+3fX+W)[6
a#b-2X>ZCM\XEd,)>+HW4R3f]AA:=Y1dT2\f(c5UHGb,<M@QUNdI?(a.&a7PUZbC
E7eA,OSPadT2/-AJDM0JgB#C))dNgK.^^,[7MB;fMdY[QVFH=BNLBI6S2>SJd17:
L+>XCJQA0aBb@DV^UA^7@A9<=Ab9KE)6ceZI3]T-RK0_Qd;f&KeX49,PIGZH^054
DFR#3(EK7eE_M/a/P,O)=bY+V?1/CJZ?#JM1ZXL-7-#&c#P#?,U2O8863+Qb[0FY
33S36#-?N01^a6?7JOa[I6QI@DV0M_,#9N5Z8V]=X4d:O3MKI:F<7=gL-@dNVK4R
0SZ17gc:8NTUR9VXV-P:C^.K\MAb7Ee,a65GKPF?YX(d;FgRgcAJP0E<;f;3(5[Z
+5f8.][Y6^;JOe&PI38]N_]JGc-9L,1>PU_?QV#Zd9&P)C>2P;+6J^Qc4M)P@(WV
0M@ME.S]UV)3UX7>8_<?K<WWE,Z^5W3fbS9Vc-B&,,;3D(.4F6E_;Be3dPP>c1+B
>JYI?QIG-=#[5S21;B)IK,_RP)QM1Wf1NPJR@L.5<FJ?AbPR65fM_/HW5FCUSXIe
QB@V#XH<D5V/f?)9-;)]VRX9,EL&aJX?5HAF2)[7#JJVSOeZE^^[VBFK22)QALK[
gL65,2/E>f.2@<VU5c16+21]_fe4b[W?S2IB0Z&.14S.9R.U&]+0Z_+G(@@,^.R_
30GR09MYP>0V_Z&<XL\_NALY#SM#;6>S@\N)eM\89(eXUQ:3^cK-[e@IR?FILMe@
T/B]^#CU5@#=.K/Z3)^1WAb#8<Q]OA5c^]&Ed]24<LT@]cdA1UX.<EY+U.]N3c\T
bC\8HM-3&89)XI7c2MXJ..\W)HdQ:B#XF)K739YQCJO?4:ZI[U=cX@(]=GT?Va;a
DF]^-&@40FL(-F3UZMS>.e@C9,2<-;L#8?aMQ&+D\D1@94@Q\3/N;dX@JO6;[QDN
IPM-K7=:?Z\4<@^:@KN>_.+BP^55?[=:UN5^78SK524,?MJYL71bAC9NH=C6E/Ic
DcU:fRHZ9TO_C:[f/V5>>FSbV+SZgZ?</QWgN^U,^XRABe89^Ra1Kg>f>VHA]LH8
>2+2^O&59Cb=G^C8.;:XV^DgCaEE@,bKT]g](+BbecILFe]_gF\6b?+EG050&&-P
c-+ZdQ4))7NB7-DdPWS^>WZP\Bdb0dKX,d<X&BWKcdC7_;HFF<4KIK7EN:C(_7I]
UUH.@KI\(1=P0WL0]d+:Zc9LV2H^gf7]EEM>]QO:1fW0P,TK:#9PP.^fF5JY4,.#
S701-DY=Z#B\GHDY\Z-(fAB:C/:IfH#_G_X2PC]I.(YA4g/db=?W)C5B&L7@<T#6
:aJX1AP^68>8Z:BC6;1_-9075f1cBOX.adIN?2O45:,ZEFfb;86eY:A1IJK,bc?W
(V9c1Yb(0T4c/VRPLg3<?20)KT?W,,^VZ#8YgWQJeZXgdDG[1N6O9dE1EH3#XHA]
H:]U)L-Z>>,?V3fc3&_:XaE91NbJ-]1Z@&P6P3J)cT>JR=4:8WT[XGR(_cW][=W)
EL8U@SD2470,Oe;aJ#16Q)K@Me7\>L>VTK&KC3\D#5_&>QK]3bA?N0>BPC>4CR.Y
[M:YV=-OEcXN4bIT_6F8dA?Hb_]H8Z[3<eE^[:a3N3acZ[d)>3-,ED[Y1Q<dbJ6S
L<E]Bc_L>SDcG/SBSY)=(\dWG&)13.?bbCSB,BI]F]fK4&CXD@,[@,=F:>#L2KDf
WcN.O,#(f36@?3X.2dX@X<:EVO]6Xg02D<bPffIU\A>,:W[R^<5:f19\1W>3\)HS
c@654#(36+T8_;7[f=KTBc&PRR_#TE:0L?K[H>G4G_3@cU&8?:5Z5@#JP+IG&+@_
T@7Z8,HOB>&^SdIfgZ;#Y^-g.8>[>8:SC3#B9_QY#-5TIX]Q&FZ\Af[5DTO7B^N4
#3PHRI:I^R8/?GC2KQE4R[Sc>Z]04BAfd>^H&gW?MIg.4g#g:<?Q;+&]g@(CSGS(
6dbe@dU(;[#?&86PU5g9b^_g3V@4B>b(b6T#^Q8bg<<7&U?Y0daB5K=/6U#a4Qa<
TXHI^\a=@,[C=VIG8C6a=d@HPbB)M:-,YI\_f7Gb[YMKZ.F/SGS=(?d&b+UI#HN4
cWHY681K([9>7],X((41N>&Z=L2;2./8,IT\T.E1=WM#1cW-W[)dVIO<O/87HQa?
/:dJe;[/5eF7WS8Z4=&W-a[c1;8VI<]OG[1NO)=Y(0M:#XJ;F3C3dJCY-BZ<-]G(
7dEU7,O7&+dD4/Y0RTFH#JFfgNQg0f36VRg/O[6>>A(\M@6.^dVOHS^MFRT]Z#UI
C@e#:Q\+.c^(O+/;&#GZPCa07UY>U?=M[3(3=@8LZCQfaCa71&&e)<IJ8(L10O0M
dM9Gb=ZaF\PIIGEO];MZZK]Vc@ESd;9L>;&a:7K#QYcK[+PaK-Bea?ND]4+P(gQa
NT0.KQ2EVJXJfX5C.fc86BgDa)N<YJ7V2a+gSbJS0Y][@[BWMG<7&eF^X]94:L/S
<5<<HP_d#Ce(#;KK9IP0(_B6M9N2(BHFPdJN7<SU)9+G\X?BQ5bO]F4f+6ff&9G)
BUO05G3c6F@>Q)[R<B.Cg7]>[&GS0aVCHa-1P_,2#>4>J<C[NTE9?)=WfX&+(9-S
TEZ<YJC50QZ[9.UN9IadZa0(0P4[##Me^=eU@0X<1M>QI;KK+)PU=cUAB5J+-MWQ
3M<Gf3:R@1S7605R&T..X@SN+@I@G+__1&WE,b\&EBD\(+-.5@bJ&XP(?1\J@0TB
T9Sa<A8&<@bd.bU]K#X2YSX>V<OeJXOM::8J.^I4BBc>1@E-#9f,940=7_aT.ANE
6NSEKR5[+=U:<>cbFT)Yc[Pe&)#X2=#?36RT>7aKN59?D9V,39\?#WH3fEO4U2RZ
?[_ZC^_f7BQ+b.VSR(9ETWVFU-bc^Z3\#/FgEYQZR45Y+963ACfR_Z.K40RJ/N3U
+]:35:X<MBP7gDVC]YG8K5cT3MQ1CFQQ@D[_M0:(]+:KCF&0d?JFE#W>]ULYV/.1
e2Z/T#<AD\F(0:Eb?9.+/6UYQ>_M86d,IDY=gM)e9S/YE4/fe/1(cgA.[&7IBQ-9
LVD01CN;gG)G>L_M)0ARXO_;H)75X-D_.U(?PL+2[Cg8L:Eb\=?>b5=:06])b2EC
SEYS.CX2bNVSVc02KTT+5,XZ2NJ4d\S,=EXVE(9YF3AYcJJIZ#I:_g0DF.\:?[B,
N[@8XdO^;:Y,Q=K-DV1D8/eU6[e2:F3(]4c]L.LfW]LdD6[1?,-E&2QW2?OD#8HW
JgDJ9dYWWH5RX;L>MC=HU\/\GUH]fg3IUdZK.b-?/gY/FI(:e4Z.(LE4c)Id(BM.
VHO67XO^VDLD:IeA<>42WK_Vc(4&d<KL[;+4T?)_X:8R(4R&Md&F_.?VMD[R\BVf
>ME60&gKfU<fP4]f5398ECL>Kg1gNLZ>JFdN:Q?B5LZ.9FH<TNHSH^S9cY_T8Q_d
-],98KL;.ER;Bb__IEgfM?-/[)DEdV1Y)T/GGDG#(#]^+R=D?fDbJ6OSGGZ]=F0M
@>&)?b-.^](+>6V(,R6c-<gV4X0]@6d1dRfY,J#,@bBgeZ27:SGAT[X>DN;0LbJg
\@a_.GBC5L+95,OGd1caR0]PZNIEXFT7>0P;@+)b..[5Yb?B<IA1G&dG09;U:0-S
]-X(NH,[NON<E0MJ.R(VT-AD)^88FQCDf]MTCdG49BY6FPMfLH_YTeU=3/#?QADf
OM-.A=++dfN1+;]V;C?PTF.;00>J>NNY7eebJ>)bP_/UQb9KG81YXZDWH626OgXg
aDD#]\:1g.-D_6Q9JZN;?YHc2KKb5WI4ZIaSG.2ZG.+I1>):68@X76GSR0NS&K.#
FB<#0;C2CN4\RI=7.RbW:5)E_-^^SS8Z?c7<N8D1BYI:+ILSf+9\>J[2:__(+IMP
F]:cQ9;-XZSXdRHdb_V.D=@#2K)]dBa?dJWIS]7&eHdHYG)XUK.EB[4QdDBJ5>X9
W5F:2J:IOV<O1@:.0GP_:E^+g7-EeS?00N\)g,>G8M._9S=I]9,=3PA(EWb[TG[,
4S/f^9JYgEEF7.2?g:ba_=M:4b8N)1BW6UdW8#TW5AMH)YAISgM?EgQN5O1:&d#8
[:&5:5)BZV2XB6AL44<f\S,Q.PJNeE1SGAMW>#H^IV^Z6@]:DBE0WYL82_G_7(UK
1X9-3b^K[:SU=OIZ-M_:FCf&HY:S^@HQ;=HH[8](RS9N_bg=>\3M+U&=MGXePXP9
:WZAa3]A#[R.]&&C7f>0VA[M?;Ib9Z=:M2:CF&b=FM7E;.bER(a;]:)PBbB+1G;7
ae7WRP=)7_<JPUJW]GUgBUU0<bGe[bI>?c7-C(?;K3=25AU+aJ_#6Tb8N.M1/ZQe
5=Y8-.Ya,gB_LEC2V6f^F&H5gZ,ZM^Vg[J63UVV6--gf#F^5bQ7QMC-Q3A.Ya7Ig
[Y/I5](M]RM_)c+7=H/HXWQ02(dCC?M+PB72>b=^AUV^Y4W]UN+XfS]9KV[NXAJ3
+QJ#LQ30ZeW8M38fDF?7#B068N2D[a&T+GBH_7U&D,7RO.d8DGfbR5@BE4XR)c0L
J8XS;\=_cTA[Z0G<:b_HO652#\8Y[.OJ@b[1(d]A+@GJ@LEdB@TW6-F@ET?]d^E(
.Y.N^1]S:^f.4:+2LN)Y@dcdNT:Qg>>GA^/g>d(c9Rf5=3c5H+OD7&;QJ^QJ>;I_
g:[\K1J+V+TF\-_AMA;;F2#LXg]<?Y;Q5?=)3b409/E&CZ?J[6cB>;AYMN/[=C=O
QGST)\>^d+(1@aDZ<_P+=fHC8g8ZcE=5O2BUC0K\c^=-OC1<@VEU+dDCeH80I?73
1#:Neb/R<).9SD#MER54N0Jaa8L2V<)VUHW:gbE6>:7HXdLOZgdP0@V:/BKO_VO<
_?;OVdY:>QRMFMee4TOR5d=@I^S9(V2D7ab1cY__T1fGZ4T?)BI_fG0L,O\GfW94
4;4T:P1C)?C6S33[=;C?3-SS/,YC(JbKT[SA#LPfU.@4@(.H_H/V?=c7D_0=DdLF
RE(PMeOYeW>L:U,PaXPAKN@N>M9O&?(Q@FI3]F4UF4GK-G2A+LZFK,?)UH)GW^.&
TG]Rf^1T29APHF06=IV(g&O3eG79f_b&0YE=JVJ9+2>5:1c]>aS+6?C4b1SfY<bK
-/MXVQ0)NVC<T>Z;Ia(2XXG2_c?EB9B)/1(Q\IL9T,5;e9;]AC;bAa4Y6)[MaSPd
D6QR5^9Ye)FO>+#&HPDb4\G,-)+:Z:HLbfA.&?K=@Seg>Ug)[PGO)F2TP>+WOE_\
a#]?5ONM3MHJ?E\(XaHAeV/JL-Da&:SBM;c3U>3)e-Z-ggMg-N&M=;OcPRZT/d4E
G<Ua.E5-49M#S,S=X>TfBIAYE2\;\:0BB5+[,OL[72A-JbP?L87/;ZX:d+TKfeQL
VA3/C?&\CN@.HgF&F2P\NVP5VBT5VBQL;LHY-SL5e.P+2OHJJ-f?4G)XaaJ\1:W)
]9/HQ7W<4Gb#SC<GdaC2ZYTW;/<W^Y9F9A@MF#=A.X3GTY#-5ZD_(e6Z\QQTNZV2
IK,R&Sd?6]2Vg<T-Gcg_Vc7d_JXYO3RaH+fL5BaIMPHbaR\EVcb)Q:YKPZDFXK4\
/ZEfT=(^#6J^-D@+4]P9B==::/HfaE(JW#+ZG+0_<XT:DRAA-DM,ZHag6/&ZB28/
Ff0N0A=&49W:9BRBQ4<SL,T6bH2:^Eg:(Dg#FY;Q.LE[,f;4VYL?A[BKdAf)0V#H
[#C[c1I;@XCQS33N#RcdG:-.X;8d8SS3IX\Z4A@>P_;#&/13_4HV-R,BT=g?7_/0
b=[B4DV,e0.Q3<]??HQ@f+(2#ZC2Wd=W0E8Ud);5_92+Q#-YI/9:E]#RH)K=<:2_
#X-NaaJ2PgH#NA[N-0?)c3XMTO/J-]7\f9(WUYe==:#dQ_JeZ6EVX>A_fC;K5NOA
/__9ZY]MLJ_dBKc9&-FHAf@5;5101S)6MKFSeb^/He-SQ?g4:Z_KJcKYW#K=8-1^
Z3Z+CJ=P_A,[&IHcI?ggX8,UH#YV(/EadF;2-#,a,)&[F10?HI6:^,5Q5:&KGZ4b
.,705I;.1eMA5aZW<HA;6-R<E.>8YDE#M&b+[cBeSGD?VC4OQBFC.DP0g\W?+:Xg
&BgJ]4@6X):L>X&e;2LPQ2VaIS3-cNN>]bSW0)0EU-f/J(g\O:PW/5Ad\Og/9OTI
.JIN,UCb;)ENRK-S[>X_]JX[0gXcN=bMLZ8F3Ga<6=N:H+CJSM8YH08=[gE07AVd
]3/S8DS]=c+/L+/362X.g6fN_.W51#QfdE140L)e38&/.Z_&7?@6^QPA2I1,L=Ic
e;d:U]Y&#&8(Ib0gaX(@8:?:dG\bH;X?W=U1;[V5aH>Z@fc(0-eI2)cKOVVP58A]
=W:(OO>IaMN8O/WW4\5B6,KD8dYID7K7YI.M@f]&=3&6[4#a&2g@6W>IMCgCgeQU
#\IX8a5<DPZWagEA-PR#2;B@:ad.2VV[=7=;(I#HN<JBJR&AO]M.d.<7Z<RF:&bQ
X^bHH+/FD5OU?UPb=CUJQ26&_M#XMC[SS^MCRZO(;<be+LaZLA#-/;\89SMU3^5N
11Z3TW\3,>VR[a&[c4-]dZ4fBS60L;eC,16.]?)>Z[1+9P=VGBJS^fH&SU11;d_K
P_<[ZHeJ[#b.&g#W_:.0^M\H]60XS?X80C-)S<(-VXMba.7?PdO\PH^>_>CN<)LI
HgUbM8)V3VW@Jc7f/EGHI0Y&PgK+>0RAB)26d_IAXNcdY+GH^WLO/_c0L&Yd<a;B
MI+11WdXgeOd2N-]g:8OX9<&V==D8?9ZaY>1?5+FS^U6D8JMfWH\aOV6a@@Dd5c\
+KN9-,HVD()/G3<^XcIVZ9I;GS.BB(Me76]Cg8SC1JZ<-Xe:ag9Z[0\Z)g-GU?BC
:dM?cL\EWc?I,X)IZ:<Df-cLaSH2Y?c^WQT7LK[.JKT#>PG0I1Kf(JLQ47<3KL94
C/4?]W<<=HaX]Y2R#Ac;2QI_8&#9Uc_W+5fO3)MIOCR=1-(NG(^6&WW[0JT=d@K[
HK54.a/&8BaNT=)@0;;ES0E#B)bTe3DQA2:JZG2_LK,@O;Q,@>e:Pg5:\JW6F:=f
M:SQ^AS[[KLZ^4#><3+D.EZL&1L@C)cN7_63a>W]\B;+H]gGY7Q+.>Cb-f_FJe;?
F]Ne=J;5X0GZ9&9c4Y4],.9d]bbS68298g1&36_.C-,D3gSVW7L1JfbVRH&D/g/[
GO0PffMOdcB4C0&dZeJW4@@YU0[Q@IKUO.6,)fW]R<0+W[B/QLM@]D#A,9P1ZCPF
gQa:a5dP9bS>?Ta(gUN4aNe4e;PeX0Jf6fTX-2E>IB35?O@G)\U7@[UX4T27K)Q)
g04DCG<M7341geC@UOb-E5FTaCTWT2UL?U]ZH/7;1B4<a.B_gd^GObbOc4LZE./_
IDG,ABdg?TgR@];#SHI[Ked+D/4V&4.Hg4gOA\WN<8/b3<+BP]1P;AAN]SH61OJ5
2EQLOFgV^Gc;;RWSMHJG#UNGcHE0+dQ@WN&g?)KO@c@^;S_G&X35&S=QO/OOe.ZI
5FMM#_Mb7S?T1@7MEF#GIC_(K6P738N4/SB?_(Hc@Y^]]f?SCHN-1aERH^/1g,P6
#fb>DaWIGdQ4H_C,E+W]RH&.-9XATHJU?DET2\7ODN^\.400+8IE;gQ_74fF/W\a
,;&WMgVTR;@/7aXLFRU]Z):I.Q35-^?DbMOS)^0DMe[)(2EYWMb>QH5O10B#W?(E
(2Y^=1T>)(I_?EG=A=IAB?e[(f8Z#8GM(6?&S)647T/9e.Tc2-IT3gVT(f7P^R:Z
@:ZZ]N-g=eFWBgL9bUGD-W)^_Z;/DU?M<HRCP\<+daS_<Q[NP4J>RcY<WHR&)Na1
J8F_PS?Q&+^\4I^QH9G&8UC:\TV-QZ7)?9-QBPR1[-6H;59O)??de&P;[V,][.fb
I^I\^4(S]+a-KfX>/d:85P8>8<323\JCbOfDbFI)13beQ_H\A0cBb&A82dG]&_09
:B61g(4AR-=[&FUOgBNA/KX[F2Z233NV=af]2[2L+G3.ON+,LM2,g2=]+6?VZd>5
e5;9?/B_&4:\8D>Ee+I;@_3_+#C0f8@0H6_d,2e&fX;MU5CRIdML@E#=OVc9bUAP
C[86KED/&(b,92I^I4U3BaKUFI5_b?2J(7XN656X(gRW70H#=_:+2W9_\N#P6^IA
DeM4I:.54RHTSW1K=)f>7[5Jc0g.Z<.RB+N\^Fc-699GS/_cA[IXa.)/+PR[)Ug=
4Tc:WQEDHO?1bf3JUeIJG@RHC>CeVHQ39?YZSa(#QB:N,4g=L>R/HIYN(=:Z2NZ=
f_0D30b<]).^eF>Q4e/FNK@PSD<YN6Neae_E>/V1F>S\>EPH[UC]A/T]3e(KJ0N7
JaL=eZB.,a7e:TS&#ZAL3e@<,HEAc;TPZCd?CP6JEg+T^@/O8dcdcP@-]7B)F8:T
e],G7UVC@TOLG;:+9FNM<g<:7_7)-1gG33RZZJaI6^1P36NH>-a@C&#dSb53C88d
\R[TO&(\b&b@)3E_FXS5S+V,EA9?^dL2Y9G(I8fU3fdF[KYNP#V2@WY4aeHBRcWe
<Kb9<+UGcKeYBUV]4XgD+A=7Ff:M[O4/aTfZ#R5.-FHL)5f=XR=-9DK>NTOVD0[K
FT-.>Ab3=?c+:gg5=2(eKCAgB\E>@678&-#_6Q=^.I,]<&&U9Zf5C]\2,@X-K+f3
.Z;Z[e0IUc3P5a2J9RXS[:-4+&,<N@Ed982NYd:Z39b=O++S<\.LMKX;NM[I#HFG
C?NZ.E3<&(@1gQ_KW,356WKb37eWTK1K-N9YCZ5<NDdRI[F/Z?FA@W<]dZSLT4KB
-J,(D_4RLd5<?1cOR3S^IHV9TO0-R/RIFMSZ6-J56HJGU_CC\?[:0\EHGgUMV&e]
V>X+aEf46PT0707@L^3ee99K+GG3]VJ(GFP<Ag,T8?>QRCWLe#_G\fJ8/(7Pg<>>
8VaG6C<)_\7(4(5P2=[_QL;\T_=^S6I?:$
`endprotected

`protected
.g+F[K+ad]U+feL:GKaC?3]g(;@9-GOg:YJd]W4(GQbKU>45bA,&+)BSGYdM=4/B
K,IcB#U->1/Eb1/C_OH3?a]g4$
`endprotected

//vcs_lic_vip_protect
  `protected
:dS_-M=6S@Ja-@@.g?(6OWD:9^aV:e@0@Q0,g6<2LP@d6?H8If34/(VC4X,CEfZ_
53U@cJSeV?gY_&X_g_/AgNZ-,18U#7\//_9.HbLfXReV[b#3@BCEdX)\9#]@2@Sb
XKIQR_&HZ2<581P]c6GB8H(?[63T]Y&bBfJBSH@IW8U;?2W/^YI45P&(NO6,,)>E
6d#U8AgP@;L8[VPM=AD-ZP6<[?^6Y@^9UQ,H^F5??2UJGR3<O#2#ISJ_+fb1V:;M
f:b]+.O\]2W\=;Y]A\3/:4O9;)SV)<+L>R7&?@A.bS88.BV,@MQ]+EDTCJY66O<J
VFc-NaIV[&7IUW.JWcaCZ?_AR=0)IKQ]E=&Z__#BDK-+BNe.I1##XXQRaRT0\K]J
J31(H5PZ50UOfWC&_KTT4U[:]#RK6E5Cd?1=J_ED]:B77<8B=A<=M1O8#EY+YN<:
Hb6,Z><IX:SeX.^J56Y=Vb[c+WSI7^(55G\e7J?P0,X-7?+UJ.4LRe9[-:A?[Q8/
9aH]bf4VG1a-,d#=+TY:RH,8U_7B#,8G4Fc?Afg-SD@FGF6Pe>Ib5R94a.5[)RKG
]V@9R39UZ,^-U^=<B)0@@02#\H-G\PFF1Z&(458J)U?CV7<T2#e;4\X5Q0(+E#&Y
^Y/d0&NO4bEO#(a<Q+MC,9V=_@XaWAG-(;DL=EPDK5>]-cKW^7O-IgW19PYdg#.7
FeA,LV]5+RHK?1QE.fbDGPSI_/^?NP_P=.RE<21TO[L;TPJLL7?Ob_/R&W>8:(N2
LD16S@NUW+?VX16LXLSG=@:DT6UWZ;WTQP\GW^<K@8KSY1eQQ6]Q7N7.gMXS(.\L
Hb16^2gf9-?-(BDbSL/PCCA/JZT9T5QNd79E6f2gC4X9f.69+4WC:T#P=8fM4<NB
FE?G9MW\./=C\JRSTHM9T<GF0_:2J)7]I\8>?@<5++Ic=:]7\SDI3F2;cM8LUF]X
Z_1ALTbaSR-ab^94NE#OSQIZA8e3JM\\0e/<P\J.RgdY@18E@+I-1aW/Z&PH[;CZ
](R4OTaa8/:?F/\+_;#+>O7?.;Z8V\U(FIZ]W7U(<Uf54?),[/aYCN#L:=34d.5R
^fb<R(JY7Z#0-@DH_a4:FgJQ?Nb4Z(-;Ug3564TVgGJ#\^#MA/acFF=PASIIf\P[
?dA70W]MRS0S60^ab^V4a1_=e?LZVaZgCO,FW,AU?9,b-7Q48gaPL4dJ?F^+\4LR
GM7F@S&#>Rf:)H58TA&41/96>]IJK/PPg3RO5aM80SOB<[@VA[<\bF=S_YgI1Y>b
TX)e\?EEAHQU<a>+:Q=<B/;SaMad;2,_E^DbCA;P<c.VIVFf)Mg,#J#\BF^?LT<b
D\=NcHBG+RK8B<])a/#_9V0c?5Kg^7Sdbf^3,CMVM?(;3Dd?M#RQ4D;\E6aJf>a2
0/7715Q;c>:Fc-GR,d;@ZI8?;#^)3O].A[Z3#QUTK9F>A(2<S2F0G.cg(QaBP=<6
dYM>;c-#/;=R/2Y6M]R4^-57a>IX#.R:(+>SRWNF,\acS3NXNN,dcaPL;,]^_8\^
9__QBUdDQ:bW?H+XB[512K<U9AY7b[/CLd+0BZI4fb8K83=,H?X#R;9[ZVeGOe9>
-,\)_-(:CGS1?G++(-.K#DS&Z+dPOP,aaTJKMP0Z@OL_0-ed5Ic3W=)D94dK68Z4
D2P7Q.PD-?1[NcYY\&X:JZ6aFO\(eW2OA1=Jf(b3,VO>f+LL=eMa(0KZT-D7IK2N
3BJW;_MK?cZ?3-?03Qgb0]H]R=2H27a)0]4<R<1(3PP)?_.I;\aUa/9GG@,V(15U
WII/EMD#VASa<O/6W(C(41cU\HLI^SAWe^V<efGgb8EK>4]?9)=9N@/=5Rge<<.H
CF0X#V4D:\.O5N<9FeYUOC(L5-1Z1:IHZSW75H=W0QN-8?)fAWIegK;DWL7fV;O+
1dLK&/2<&Ic&KA\e?c[@L==CZ<F5<\&@c:aQ27+BRb=.A@[4-I80(A8,=e,/(+@3
MU5,6RbXcYTC6@T:.\TCN,Re3aS<9MT1>?7S?b4?JK+X\Y3:e_)B2:c4XUV0OC#=
^cYFSUN)D6[^)f_[@_+(7@2&c+&MKb23WD)5b)KQ=^#]g0f,@5EMNG7AU,Z(@bDE
S>:(Kc@3KCV,LPXK4->F7I?4g1Wb)cONXYe<ODNF4ZNIHU5ND@2&/:Y@e/(P,32K
RE+QRdP@+.\3c5A-,-eZ4T\__/\Ud,W)2FDA^]WO1c)cbCW+cZX;gKF.#B-a57Hb
QDA>We,@T^C@(TG=Xa&9e8HOaA5VV<8X6@,L+a^I,.V>1F.-7BVQ0NfQ;9^RcX/b
+d6dJB-aJA(K1###<>E0AFd+S65N56EN)N(Z4TZI6=fT08C.Ja[#Q85bNdVJKTV-
:d/=a6BUF?gF]SF_?W(G(Y@DA&?X,A&aF@)-M#2+94XYc1H0cREbY3,2ASGfKD7U
:5W<_.X8C6cTOa(&YN4D:SOeabc;d+,BC-9&bE5XRePUNFF5:T@d[Ge1E>1D7PfA
P73_(K8cKT#\[V:C\YCBR6+<PM@#Fa><L>-O1O#3NHSY1GEEMY]O(IW+1E@4D,?W
HbW&9_//PTQQ60<WR0,M,2-(;+Y-EJaXPCW#MVLP]&TFAa4=Y1WW4H?(VH.J1?<@
VLHaP<ZAX_MQ3#5E)7[INS^3Wg/F.XK>;U/3b]=0H<2V.OP9@R.eP/X:JK=]\LZ@
2H[BE]L0-NE/4#V3<78I=O8L0aN5eT)_KA=-50HRIgURH?:e>F\[MX&GA;SdgQ&1
A(c.SL9b;Fd\1],P=IGX@AQ<XW,--_YJKIW2N_85d7Yg>gL4]=QL,a=O>[Cd;ece
T\3FeT4ST/P-UT>4UJ60O(=+7N\d5WIP#SXT6;QRX4?OR6N[_YR=9>E&AM]_M#D,
BT;J>aG/bLXZ=6<8<;RZ@83@[[BaE57JEG(/-.U.X9O2a8T&NUBH3ME8U/1TY[^8
UP>Db/+RX8A:R9;D78N-FD_V:.gX#[+YbJ=T,8.9_Wa+d,KKJP0V-Va+5R=#5:,:
0cfT95e&cb&bBELX;Z3[L<^I@c?5;FO0Ua6#<^9A>WB^9#CeS99VQI<AN5T\#ZJE
Q5YPH\#>CU9_36]7c5IaP@YKJU8Y<#S01<:A^F&50T>(&OJD=9DH^#MRc=KYd=Ic
gPW8B<DE^UM58LHF4;88?6@AeBD^Z)EE>e:.6W/?9?H6RV)91f<];/--Oc6aI/@3
_fJHb4gKFc(5Me/(]If\Hba&e4P7_333736T<EHBa>K4&4[9;3^e<NaG85\Y&OCQ
53F]U<ZBOZ?P1Gd6&M,VWMVLX(<K72ZDc2;Ze=)W+1-^X.,Y5#Ie]B&c(b?^FKHB
,I/97OD\P?fe#HE_)d?825O\HUV>MP\LafcHKTHbb8D0CKb@)2.;E)LAe2,ZYa&/
0V(#XD6>^e<82LHN0_+fg=<,:Q2TF0gaE[WS#-,R6F@9,Gd[G92b\^2FgI#]?C]N
PcJ)Od16VQaKM9SI(=FD17&QW&,XW6?OV0GT:5_\SPQG]]Xe=eT<d[?1HS];Nc\P
ZXR774a@;9N9L=,0:bE0LdDGIX?:B][F7OPKUHTNL)J2.?f/[>)DJQ/0d#;-7E<U
b6_+1T11ST4EKC?CVf+a05^gX=LRH6&=41]CLKK-TI.U-M964=>GG;eJN<69K-:e
DWDA&eFX2WA,YNN-F-:bMK91&)g1>/ZLB&=9--Y&3Y<HB?R:,A8dF6(E#d)KK0Z#
?>7CME,@_EOd:_J5]+Q^FE7,;g5Q/-/gI-/V0Ib,8aMGLV0@)J3fe0CcW#Z-^1WY
#YC/\P<0.7cL5Q?BJQ3#DALg2\KcHddOR53V^]+U0<:D6CcUW5g2+e.CHY68<a(O
#D=B-[cgEEOS^:08X49YVJI;//<fA13A020?#/ZHAH(b_c\GPb5>IL.L.:FfdN39
&_G>526a4[&GJ:VPebc7P+@=00X<_-BK;cK]a@_0SHXN0DeHCCU:,+aHW,J11WLM
R0_Ka]<\Uf3RHQ3/\RC;_8,JRLBF/8XN<SYb.=Q5^C7Lg+;,;5Nd17Ae0OUbfdH^
ZA8fUgC[bWW.?70E+<2=Ve-UUMDY8^T[A9+WKcabDc_bg2C]\25<AbH2ae5C./M;
=F@S:<M535feZ6I_I61<HZ&@2(DVZPFa[[\Hg07-dZZA3N;97:D9G/207Sg9e)T(
UMfH_OLd)T,8AcE0ZW>>5RJ:4[+#[-@&E6&GMF1<@GR33J\]^;RGZT0>3X22;\+d
V+SOT9Jdd#X)MS+@(DF6V+X2G>WI2G72[c];:1@(_#RY@PNU@2E[VCPF?(O<c3K0
J[7>HBXF@LH?N)AQW4bQY]5a/eG+T4&dU,4FUGM+DPa7c]H/SP-V[N76W#-/3c[b
B955:,NI]650[Ogb&(277Z\N9A._a5Hg<TBT[6G;-7VRG0T1D.P+G(:=eHG:c^P=
[XC7#3Pc8DC>?8?\X,7/?M;_75IEXHfB<H^V)1c#F/,8>2<FX^?C0TH2[_CdB980
e(,T0C+MaA2-ET&#:H-_dQ.b5b<PUI_FWGd;>TW..H?3Z[D33FQ2^?(&<Y+YAYPd
?X&[>P0PAcg^M8[#4SdR&\Y^FbZ?7<M?Fc94?=.ObQCYCZWJSIScPLNOFFeOY?10
?JPM]/N/UL=W6^<.d#(O5>B4-^cPV-4<Jd6.9SULQ7cJDAVE8A\CV2-4TRXI>]G=
d&=<[(830\)Rc0Z.:>TZ\JL8Jf52:.HA0gRWaK\H+e_4-I8XISb9EKS,ZM&bSf<8
0/8#S3;F8e2Q3+RL+I+Z)#E/]e2d]83(d-^5RB[e&K9JNL=21TAbA=6G3<^1-0Df
L1H/cN;b&U@4WP+7NXJ76.KDC5Nc_=5RIJCM1ZcHSUGUJ/2/CT:_N1_EO37VV2M7
T2=-1aJaHMN#bLG.VV>A[IKIO\AAU<8eg3FTg04-?A7-XU]PYFca#M2P=P=_OW[6
^Y7X>ER84I>Q+,Y3-:aVG36M(-H8+1NN:ZG?fDZ86&0/)HeFY=B>&aN6]/74+O.]
<&/8cKbg1Q]YF2G6A>JF67</SEGL#3IKKcOSK&(+N6V</::_D,IX\J#VQ,bX&[C^
24>?Y2[>MU\Ee=0)UDCgQ=;&H3ZKQ7bQQ.Q@d3CB&[;Gd&N5[AFTg2ORV[PPD1/I
9BLeFJIe+)R@^YBc\UK1_W2JA26U\VQ+D^ILCSc5:RRZ^UTZ_@O:-_Wb]]PBf?:R
D(X7BN/.Q6H]bFI0gV&cGcW>&.T_G&R?_F:0&a1]5Gc=<a9689b(.NeF4DQCQ+b_
HRWHDEBD#IET#IGLV&088f3X/U/e4<a,47>(f87FL,UKXZ+J@FbOWH7KT/:]c+NY
OL;<]Rb86.Y&C)YdZC#Ac6fA3-N1+\_?QL?CM@_2V_SFE9:RZD+,^UWcJ]M.Y-@<
^+SB]:05-S&dE]9,8fJ=ccP0F)gA(cS,6B>ICN.O>4PgK:JbO?00:He_(]b3<A\-
gFYO.(K&4[V8U9CWeUDVe#IIIUIBD@\Z&2g8G\8@e8VRQ[3\SQdEH;QN9T[Ya;),
Z;(8P&b=21WPWE-#E.^5F#]OF#b7[/V9L05ZB4Jcb-,N_b8Fb376f6(2-1<7VDF>
C?QO<_032&U0LBN0:KWa.A@,C>RSYR\#bSI20BU36]cAJ,CJgK<9=aGP0J88^3=X
2g>=B@W6[;4-@Y8,(IJ5MIWJH)U>82&F^OXI,gLCL^87.Pa:9F/58UW6E_P1-e5]
@dX3/-W??/;9>\&K)\NX9T^?Q13(EZG2\?Y)>HKCTV-JdX:[2eSf#C,6/OF3XJ+T
?[OfUd<GIFB1UXf)eWadX5,<DbR;Sf0ZMPL(0-B8X)WP24egLH.O4-fY\;aI.Q,:
IaI9T^VNIMV-M.2OW\B\4QKOMD[dDK?f-9\ZT,K^:<NKd&6;)eGR7C8Af-SSB\a:
+6GYEgT/JML6DcV.Mc/bK5(OS@;RZ;H0YO/N8]Ede#)10XAEFbfO6I;gc]R#:WWU
&N2=/#\[WE5eV5e(K_N^Z2DF69L<(8F(\F20K=]:;.B1KMB\9?2BM>>GVKAe[ea<
7-a;<W7(@9?Y4X0R?^U\:Z#8&[Z#R8WJ,F5fKW,QaC?5W2.[H(/;@2<D1TFAOK@:
e+6I6aWd>[1-JT-/eQB<RGe<CTZ8H,)#WYJJ4&fSPFVf2bdLR+I:KD-K9NE=AaS?
H2[.2L22;C=<G2-&6D;M3f@#US\)K9>@f=IYTZUPMIe,9&Q[,ZVF3d]6:6e\-9:4
LTKCeY^-;ZN#;d^CcfgVE5KCOf^W?,,I1ba1W(PeI-S:efbGH7f/?3DQ#I7DX__F
M]9YZH:-^bE,/UVI;&PQMM@M1)XSX<WV?gg0E(TO);++4)G)E+=M7+bEg/&X.Q?D
).-PMG,[V]F]FgU[;>P]c38\YCY3]:R#YJ[N,<Q&2;/.J;[A-GTY\\b.^)NV/eIH
YY;=cNPY=aM:]\bP6HGc47^BYcL^H:NXI5XHB1_[dUES[BH^=97=1=\ND3B7,fIT
E^1e2B[Z?YG@[;4N2V?N@e]<CUY18-GfI&N&Acc8;8C2MEfK\aS,gM,g\+<ZR7>1
:\,[/),_1(bCQ1.9Pe0THZ&g?4)g1ba+GG<58S8J.Y#\I3+0@OG;9NE:9FU9T9Vd
1<DTfL(/Pc=d(N?]T>KBPdXM4]=\52X2Ra\e,X=>/O=@MdWC8E9)N:BT0JH,],@5
CDZP4CE\E##GFN0=aLI2X04RJS_e\#f7cRbeQY/f\b+Q>B6,B)R3F2A#H7cCb9&H
^/1EN)g5,0Ee/MXVG;\28Dg72OH4.W;T#OM2=T&<cU)ACJf>KK@O(7&_)d7:#I&E
C9P(BS)PQ6>8NTJ0b_\N[@>K7H=C:<R6#d9[41CdS^S+,bKYdWb=K+/_Z-PU,FZe
QaMPCKGW&5,:=&9W<[#5:CU=(8cNV)-1bbCPB>#361Uc2PK<+:;R4;7cbG##L&49
&Q<e^_fB8_MIb,8FIaM)1UC=WJTd/DOS&CGW.,:Q24WXTHXSAg;,9f5G0T_9)d[8
f=c<V6=/[W:])JM(8@<[Q(QG_8]dE\ZPTcHIK2OZWI+OZO,6Eb,5N+N;71(5SZI[
/Yd3I6.g<CIH0&aXb.@6fY3Y:-ZN1^YBSEda?D]N,/)DZ-edSQ3=1V#+\<:7W7aG
^K+Q2cSVMSM[]b9FNI]YGYGZYdADecEOC?\Vcg=bE)(Z><J.W_Jf7::/KDAN?&Z7
44G?^&9X-R+PO#g,c7+cBOM;A\9,=6D53)[,;F,4RR9N0;a>E@2](,OdQJ=e,6\/
+)M-SP7Z_\42Y6g]^6BD:6SF90g5/&CR5X8]-7#<KfA:R@A,+1M2I5BDZ-SHNQ^/
3DN+Ta+gGIZgR5#8#[JcIfD:JV5,gAG:UP5_ce(^b[PT#,XV)^Z?>ZBdfW.B782W
L36OFC.fKNGb70.<9SK(HNP<D1/F/77&@E#-<.KEMT<#+WL,<K4/W/KWEV-d#FQ9
S7L3f/JD,S#XJ#4c\OG?f=XF;J3AS/_Zd8Y:+2(MbRg:OA:KZ4#Vf2#6EM)#UXPE
9U2N2gKcUTNW2Td6C6TP.FJ#ZV@;_^0X/(OTNc-^M\#2YVV5IS1QDYESOHbdBUM9
<XT)KZ\RfI;a0<B+fdC[@>YbTJ]1D6:ETcaXN0P#D>.M8NFU2\G#9>9F0WH=[KFa
Za^/I7/@,E4/T<Dga;e9S-,8QQ,UeV:W_d.\8R<9N\1L96##TQRJO6@cPA-/O6gB
21/0F<4A)HHbgZG:@aSKK5-TYT7#B+a8#K]ZB&:D16D)VJFM[7;?6DAGVP625,&P
7U+e1DVf#c));KVWEgbA]8+RIZb(;Da>RBgI;5YUB.2\=H+<>fcL9NY7g-BS8bSM
CS5#_2KcgN<CQBab]0\)),Y]/e#=c:4#NE.2BJ>RfIL\P5PU:LY_Vc[Z1VXWSNg/
OW=24I1V?J)CFZefbC(9;0ePc+gI#_D=[K84VY0cK/IgKGeZ_9f0e:(5E=;5M<.Y
C<Lc5,9]YTD2BLYBdgWe(>aNc@.QA(,\MP2Q[A0?IV>Oc)Z2:4FC\a8+eQEQO1MG
//C(@Q1)(0Q=(>2LAKFBAV6+(MTLedJcMB+@G4.6UGG47eQFHRHU:,W.KfF@2MRF
]X#e]O?dgMC=bBG2Z[?,Aa7Vf,#dTf3K6/#U+U:2.Oc3]J;:JC:8:ZVd<d/0QLeU
ffdXfZ7\DJc2A2]bL(PV+EF>@B15/C_T?#LC&[dD.HCDD3a3NcE6Yf_f-g5FBd;J
-TOe<#Jc;A2IA6ccAIE53d@6V[TbH4CN:LIba3VH[9OSUM25.c<EC61;W53([3bW
-\5T,G\AK.)N#FX?EfWd28?DE13L&Y^K:9RN(6K\TO7F1c+@#[W]6(XL,YJ#WSZQ
AU<#;6bB>I=T-2PbN]<8GB0_QgD:E?BB2_YCg38^;FB.@af6X36a/YN:Wd_\8#eB
1T=a\b6#IE;bbQ=0.-F+[QKdT(aF)IXMFS23WgXV]BX5T=U4873M-_<-FC[c[GLM
ZE,7<XFU3)(1,4G_TIL:OO6GU)-(eJd,=dQS9O6;H08)e#c#:XLK.D25SA7D@W]<
5K&RS+ZZ95<Q;/MN5ENL:,NTEZ]>)FaLX1LC)4WJ)FZIF:QT?WFL]&V@g^?956NN
eHb1e#4gHB:C9?>1VBc=+4K>+Sc\+Z3=YBS2(5;QV<)5d&[4-15.a^9?PI3>,I.f
H,G.G9WbfFHN]Z)Q8:[V3(7:[#Y\#EDbBDET-3OJ+D7ORE2#fE>7:>9ETWfNEFM&
;XFSAfFYAJ-@1?^<P^K89#?E^N5@\;Y02b8KHG,D/H&c1PeXQBC(W43^WaD:2G:^
LGXMc-aA]K08SN?1@DS?CCZcGEQY:2G9Fc>gIc(/>A3+63;a4KZV2E,0/SgZ0QWF
6_(2O<+;WQ/BXRVU:E?C[^6(IY#NNKTY5<4YDVB3NTQ9HTTB?c--ADD2V?N-Ee_-
DLW13W/a>]]3#Xb?=]\=91J#UJD@P_dKN\]MZFQKfEGgB;aTe:&V\]82@L4>U.ZU
8?2[6MIEgS2^+a4B/F61IKNS;:,=0c7gU_HJ>a+1aHPV6O9ZM?GF65#0[;VE9/(K
DJ3\P2C[GeOF_.Q2V<3&5M,He/BY:.YGR=GbT]\gfP@:+9]/P,J1X,>?#1M;K66+
7aX8YM#g1;-69a56+H2eD[aBLRS3Zc_X_#=CKe<aOTb2UA.]\PeUU_>6Y?VK0E@/
:M@dH?;OG4IR@AFXIO7MD+C+P8d6aR9]TA(RFT@d45(/UNJOE#;5e#KJOO?IT)@d
-)]g^1c?6cV;bAKLK:1MfU#EW+?T#d@;gbZR@=;B;VY],SMOV4AXG9V;Uf15d)DB
=P8Q_1cQ5(563JMf)O=KZ/2AC[3/#7+V,+cM.QMcEA:2&\5,_a]A.d_P=AJ5>D85
W4P-4TI._QfZ4b>#d?^(=@)De7+:WSF]\Q]P\I=:aDAU].VZSPB;#e6<LPJHM<M2
97ZSgUF)0,]_b7UTA7W3O5]1;N[WI)LVg25UH7;9V>^/D+](^#5d.R+JXH)K[;)C
.\\9MSe4;Q>A:IZaF>LWQ>L?__?C@/7CX58<\B<P,GAR4-YPb-SI0<0_8ANBD0c<
4DQdJbY3U+Dc+<e(M,&F?_TX-a<M>fOP/aUGB4XH6;IM4]@g_Me0c=2WPB/5<bY_
5[F:PEAfKIc?,IV91,8IT6a5K#B<6)Kda&3e#TPA=A@XBQCWU>](?bUWcQ?4UY@<
2Ob\7ZZ9Y:?+g&T8I1D8_PJI):@P<:P8Y=GRRZV,f]4_L&5.VDQQ=+?0DX(_-\6;
,:-_J-ID&aR;_S;G/4:8WK)1b8IC=@DcO5?_J_0f)T>R\+ZURQ=d+Q<(F=?VcQ5R
EaMK4d/]MUM290A8]QI^M+38BD+61[bE3IcOQM9DF[XXD/]8QAN,9Pe>A[<.gYHc
eN[c.NJ&0=eLOGdR>S_;HbDJe;5f,#TD1C&;)cK./R=BM8NIFV-V:N(/^;RU.B33
S-[9/bfFMNF0+bGbL\ZC4QC=OfW6^[BYE704a6=f+GTM.V<Y5SRJ2;D9C2c5f0KC
D3;E0(.&Rf8+gbK7AIWVcKKMFUO(OHF,/5=/(DAKH/(C9E&A9I(M]>W6)<11H.aW
.=QUX=^TX(=E/HbZ2(.W3GOHSX_ee>-F5gKc?Vb>5/e?ELF=B0AOLg@GdFD,CI@4
L<bEDOMc/3/;01EOWK&a#I0>b7X.\)HOSVVORILWQ<_V-(&]8&D^<+<b<OdIA2O(
]1gEM4Sd95<Ja;?ZYgT^D8,C].5FEa/9bb+LHPace8E,XT7VI.D_KV;QA4L)8DU_
e)LM(FS^]YK)<-5)X/;EKOA0LL.RKY_OX8MV>9J9@.<PUV:UHKB^_;B:GH/KW1;U
Q]]_)T8T)<A?5(ee7QgGO&-[eIQ@>U6)O3#]?a=>bX0,94]8O,VgY];gT]b/#+bR
NPPEg&e,D::+5^[@G]F;5YSSIJ.PN8;EUOQFF3aL>V[A0)O/>#/>d0W3W:dHbaO@
[&GSC;LO(&ZSJF>0?E)LDB:TPNOAO&7eNL/@b()7C0#ee\Y.JM,?-07<X&[GF[gI
R=B=+=>Ra/2L+QM-S2CASAE]P@FMU<O2cN4[ZIg1DA#-E@9]M;5P_/Z3/@c.15De
+fN8TF^M],CdBN9I1_7LY<KAI_;F61P&;Z3GP#e<VPIG4+EZ=g3&dd^_\9/.A+Tf
ZUY&.2ZbDLRK2MCTQD4+^Q7f6-O91QRZ):+T<BZ[(XfRI(9MVI@V?6Y;31[:e[&=
SG-7HOUN0^SGRWfe9F9Yg9[J;aTW=T\96]LV<;MEdfH4AW1>WG)=W^L@C]\9=9Ob
].((1#BQ:c_a/G/?eQ:6,Ba1c0G0)L]:G7N^O;:_)LAT0,V<KME@E>G6]H[WN_LQ
7ZRBN,4+G,HYfLE+/f,:)gN-Z93T38[V>[Q-Y+3db:E00Q&4A-a)Z2c.Y?1?#Mb)
_PC9fLe+&SYEU7M2YXYR;^[,3E#M#4,QY([_NGCIO9DVQMWGJ_O22&5J6]Cg(C90
RL\(PN2;R>4QN9/5,c0,>^S)gXff&/J;=eMS80c?aLa5#geE>c/d4cbE.MZ=4g0A
()gR.N,(7=F7G.5RIYN/.K<V+;IPB]Z2bJa&DKWU;D@X]3;PFb^MU5^#HBL)20fP
_LJd^[Wdc7<&OP/Z;=NI_A1Uc4-(Y.M9bK\[E+I=JNT(0)a9cPH6XcA[DOXR\><R
3:3H/UEIQb3A[&DC=2Pf#2MgbN9T,eZA^J7a[KW,)dLHU6AS,RA=2;=\Z6J).HUP
N&>6eZL3c;SG&KA4I+eP?S?L-@Gd89YY=7I[_=^Mb>NcFcgU]QOD-;X+bYgaJ=T,
=F)IK/Y2O;TBaO3SM5Q/<C]<<d:Z+O3B4TdK)&4QR[(#^_aJ(@b?QJX:H]GLb+IP
P5#:IeZ@]LU;T]:TTQN?I#gU]2GGAZ+Z?D7PI+LL>Vd#4MX/g.]3/DVZ^>N#Bb4J
J/[d2ZJ732ET:cfOEY=U0.EKcWX,LR#LWIYY6Ge,c(EK/Z?ac0aeF(,Y:56X,_@(
MN=GJ;UO3gHdb.,(M2N0BMR:(X^-J^M8M+=UGJR3GR[g0)RCIeca],]^M,d?@]++
E821;OS(:-:gME=^RM9U?SW31b3XB7R0DN-#4OLFZTQ.Md@G/b<F#c3P<aYNcA^/
><6)<\<>(@.Qg3IcVc>gSW)[AA6N\1N[?XbY]=/ME7OgHRb<G2]^dc4>b?1T,AU4
d1RCa+GH\7.EX03Mg;XMTXZQ<P1@Y4Y>e4=1JZ.=b+JA9_I(TY,^C@]XV,&]P;0e
d&&//J9bICSPTUQN3>#?J1@Z8UF:[c7T\U+Z?.8<FYN#d0=Z;gcC1V()C/_9g8U+
.L+S0J/\C]3B,@?B==8=eW^0+4Q/a1ZNC0fg4#830])X?V<a@D4@Q.fKQ:<C^Ma6
V4(76WDEdZ&BTC#.XBX4;dW@b)f5L[Z6D1B=JF^X5N4]@E<8(X:Uf>(g,WOUSV1S
XQ.8UXT;d(c1McC.]],97)Re5[,89C+(JY.3U5T3F>=^LA(c;R>9F5SJ?ETgD502
0;WDF>-8_(,I;Z+d4#]?^c/Ra4P3aH7)>;G(UK=[L.(KI8eA0(:C&:IO70407WY3
\4205Y-/>Q^A1GE1_9]R,aA^R&5f.O?\Y@_=\aBH<1L#cG<)B2PD?>=_SVU4ID8Z
?.S^4:AS7^eE&Eb\:63DVe(1H++O[cR2Kf6aSVbWRM9#b;AIZ[2b_Ee?4@?#(7[9
KdAVa0MT6\c^APOM:ZPa_T>TP,fUBB7]2fdg^.\e5DL\?+eMKM:G-(LXRL.+W8KK
<XJJ(RReY)WN4:9ebW;f+4EKNDZBVB4CS+=6+[EWU>Z,A)e4:=bbDX.@OT#^HC[K
JaQScGKAa\UW=#Q5]&a66gMIMUdOBZQ0U(f^G[Jb.O_=ZZc^;G#ZT&0bPQERWU\^
@.W5c7Tb1_#;ZT^AS19.LNT_>J[aHJ^VU,15]9ce^G?I=E7H^eSNJ2[DaH;3B<:H
RQaL,23#KYL.6;MJOKOTK>ON6FHI;W]E?F1R\,5DL.];T2L3#e+>:</8b^HJPMgD
BGD1@,0OcQ3^cMgeGRaLD/.F)d]bI:_9C6;0=J&G2#&&@T#1b>e,B6[[T0;]6a04
[7\R_:S_.38Q>Z98Q(eMc3+#<.[f73<Z=0#2F_3dFe^dZ7,&]MSZ4>Z6f=BGCaVT
BCYQ?0/LNb02/10b;(SUSLK<[S@D2;GK4TF6Z>DELg04DPBN+,TT0U&a?f<-0;)E
]JSFPRF&4/,bA,M&RWcDQBYXCW772b3I5-,c[E\J_;=]eAK>W>H=b@U(2ID2Bg(]
?\UI2P8#[8[):C<\+SMOK+)N=&,82M6PORe/L=d_DB.&&](XU1J^HW6/[dAg@ADC
R0(WV^.\S]FXS>4#(_,M01Z.Rdc6b\+H5b9D2aV23bK@@-&\S(2L6^H35Q\8?]=\
/Q2,^2;QBSF8H)8g85)J[/aZ4=LW&6:D;\HYU]6(3FAY@J<74-O=[&JI88@.-9Fg
A-Nd:^PeOe#W848:HCU29>:(MHKf)aa\5_DbQ<&C;-]E1bPUMg_&a^NOV+M1+;I)
&_^[9b8X5S9R#d_3;S-7=\13@gH1HI;73;LgRIgM(+0(J7N6TA^VOO=c5TDBg#b1
G6BK2?=5+=+AdTAe-AQZ?1GRFe22-f?OBRY(7;0c\a6:3_ZM]/-7(X_0TMVdQO:4
Z+OD\^.dJMYbW/&)M6HP3N&P#8LF[4cE33@&cV7P.)3EJ#eUQ@2#[MWXTgU_/BMS
[@?e.8R;>D&e7\HZ\YVB>,0W.D1BQ1KF_fB(E>#U\)UBJ)NJ_0R97@3bMgBL#KA/
ZL:OJV./9S)HI1:2JV2f+V?Yeefcd;S)<X8HAT2_B4c7_UM@ZU9R/\@##QK2G3#Q
=@BV4d79R2&S@eBPG&e:Jb-c>])):Q;a??V=67RSg<+>:-2L/NeX-#[P<UP+CI/4
HT[#/HZ?2/C_cYQ?&G_YZgd,e2WHZ46Z.Gg36Af,[f^.EJDfbMTU#1(31QXZE=F/
,TfV\fLE9:g(@=/2\DK23__J\):c:3[YCRREMfM20@Ba=)@5+J\7A+eJYD_)D/<(
87W6#93@M\+P<XS:4Y=#NPd&G+g4GePWVc1/^\Q^:JJPc\2+EW@DK/C(S<4#Xb3f
2Y>PWT6WeK(8?22b5V=bQO4f4:+G_:5gM].ZDGM0b2bOJR9c#+Y\c^T]G0SLGK3V
^WTAXG\&RJDLI6Y&#Gb:^\MJWEBW0g@=4VT0TIUQPF,]OPN<Mab6N@C)_(2)>^NE
6F,dP_3f,7aZNFYV1d3beE2Z-N4I]YX#,[><C<1_@CMd]dTKN.O:8Od[1_T;3gLG
7b(6W<CZ)#-7N&M4gAIPK)V#((B;&R/:5?@cd(>H&:7)UYT(;bW@(HB@BScC&JFZ
e/]@Q@TDWSZTUQ,+3>7IM7P#.E.[CEKJZ-:]N5;ITZS/,DP;Y]g_Z(V&gLdN+P+.
8f8).bJ1SY?F0Q\SAQ\8=X(5/-KKQ;)DT(#1#P2Jc]_97S???b>#LMf7<D\E3R6W
dO+7S#I>bZaEND[59abAW;Vf?ga@f?,W#GG#OHOd]f9g(Vc?6b;\#eL&VHF,S.)/
<]d?TTD-(e)&AcTEM#cC@b@MgI.9LCdUa/>N-Gb&HX@eY3QV>CP.JKH]YNC5YA\D
4<17+<\:YR8TWaa-RF9Y(7bfE,#FM.XBCbI85Q;R#e&-.0^H3a.6IFE01]?OFEP)
.aHROC\T89=CJR\QK9+YAQ\7H\IDO200)=CJ=Ee>SZR?REKQfURL51SHB^/(8aHP
Z-B=F#GbKb)-DVHX<.),H=aTBTJ[2MK,7Ga5@29-PK+E<M.JWSK-6Z)R9S2YI>UV
?b&.>0a,GMFb=BA=J[S12KFO5ge?RER?N.FVeU?_\5R(g+T<O.>Oc81JGM#\XKR:
#L[7S)LE<^g5<H^\>:<T3Gdg2T]Ka(61Z=C\ESI^<:Q1O4@dV5#2T]--./6P61,8
6?_/S1\:--M9,D1aO,c;^O&=?N2R>3C45#R:W33-296P0<YF_Z4VN\?e9?C5)46^
0@HZ?34@K?cIQH5/U@CA.6/9LGY6LN&F)C:L<A5Y.J^D,J:3Pe/PMgG77^#NbKAH
YW1W?\Yg_gQMSGJKGSd9fU)UL;5B#gUHLMH3C_WC^Yb&R8JRc,&IK#VA778C>)5&
Y]dge8->MXaGf8CGJN,1#@.LCc:XRSFgX/II6FAF3]OE<caEe+ZcNM#d@:RR>,4W
eT;>N&YZT2)fQaeI/cATgR#Z,XO_UREg,1:Z5LFY(GF+X:]UY?GIF294>=S-=84O
H9HfWF5/Z:?UaV-FeeK:((/:PBc@+_OGP1K1;4(@/VG)=0:#@Kc4#[&HCdeMT>CI
]KRI73SH(^]T0.gSNQ\K5#d-AD4WJ(VLI,LgJ(B44B@NR=;4CHN7VA.9O4I87(:Z
DQM1]1]PYUTTIS8UaS.#+LE3cf4KBSV)3G5/eZF60bSQW73bUW.9-SQ<5Zf,E_9=
WJJPQ4R1UQZDN;F)_XI.E\PNE=57ZD2G3QB7]LS=DIJZX8Rf?a8M4)eW[Oa>74_6
Tb)<G3-&3Mc?MVVHQ0fabJ:Ee[W=Dg)(0G<YB9f<0aYP53E[C#O@^D_DU:0/W[G?
24D.e049RLX@USA=5fd.SeZ>S[79a?:BA\NG;fOO1GOWW1bD39-aV(;-/H1Q>/7+
>T4f/?O8;#OQO?[R.]g9BY?.e4_WE40)RLa)OD1KY>[+T3E?V/P>RG5;BeS@]S4)
F_;FTH2.(AJ>[;E-cL]CJTG&0UgaOe2SeA(.f=,Q,K>+5eW3&Re=>ZbT8(Bc[GK=
K),2Bd/[6;NRcCS^.SQ5gg^G<TC5SV0XW:TTETX&Rd/1B/b0d>0gO;W=J;EMg(>Q
ZSL@a&E^AZQMe>6]Sd?JP&b>HZG:e6X;,XS68:b:3E;b^LM6cRbgb3-D?^<adAS_
aHWca,T1]8QG8XURT<6aA])S-X/;O_2BOX-QVUdV7PbX=X5S(Bd<8Yg4AZ^Z+Cf.
(YM\Wd@&9gG-WW.]G.f>]Af\QR;9P_]41=7[[OEFLb;Yc0C[3Y?>9IeIW<EY+3O3
:;:[(X,UD.2Te1a\/7NB2Ja5GLW382eV5=M/#Y4/VWUB@L2W:^6^-7X#^b^R\0IZ
2>7K0UbgE()0#2beC[OL+_(;1QRMPJCd;fKM+Td4B67N-?FC:0-,PNULR#0N^7<J
2e;&JCbFOFZE)83e#eS+TV^MB#_1,^]1&+05C17?D^Ze/)VB?X>U_DPY2,cC1S(S
d?e.0&O,+F/dI6P/FaFBG]X57cEU(V&7Y]U?WW7Q54:1f::/U53@JU-;MURD&L+#
09B]aE8954VcDF?\@(+;_/F9@Ve4>2+CKT.B@W-D?UPW2fOT.3a:Bb582U)3#),e
&HTd=f8-3A;@GR.6,YJGF_07aC>U(ZLMG;YAXN_,(c54fA=([);N>a]^.VJK7),1
;M7YJL&[Sb3/#;DMDNS3[6)b(\G/B16ODC(bYcBI0d,_/36UH33OC,cC44D]OK.N
W:KMEd#MR4HaS21IR:]U7>L][^D,cbP9De9.:23>)DCb15ICO,8SK07CW#HJXZ>0
eS1+BW<+C&6U_d4:]_@4F>/EI52D,>S7fe_#(V4K?ET@c3.&EF;gZRH5>XeV:S8K
=AZ1Y@D#AQL\C:UB#G->)8#3&?HA5K>fCEdT>#>YS&/V9:Mf:A[0J:4&I-)BcPP0
cba=QSEe@W<4J(J5+CF](1<Y@55GKT,0,#W&)Gc5D33<]6@D):\A:eeT?#Sd:)dB
B25&eUU.B.Q2HIfX8f\.ZdbKN=cQf3X85@U+_5DbB_egX8>J9N<EDC&cK<()HMUU
W_+=UU<K>+<YS)0CTB3PG5T0c>QdeWV+L)fRS#cf^3N3K?36D@+JfX#ddHIJYMM]
bF?4C;\9)__:&OdNB:F#>I9#0Wf-)G8&96abPE)N@W8P;RR8SbbcV4PUI^Q8d@X3
\/[e.V?)dO6=LO(f]@&:MB5)ecZ_&[AF8OTa644R>6W-&B898[J)CO\:NE[De.=J
D95S>LF8.5RA59,c_..efdT-7XbX\b8P/[B?eY/YA-c/fV4ISU.KY@U0EL@OaddW
)SR>MV\81B877R/GNE:PCDR2I^KIIQ[+9ME4Kg8X;)X.fP=6<G#E+IS>D6_SQP_U
]W2&TN<-cKCXg[A^?7M?QK22[IF[Q@PTf4gKY2WV6Y0(fI9BG;-RD\@T=GVXN>fQ
d1HH?R[Bg5g&?II;F^-Re([<Z7d0,/Z6Q.e)[]F/(&BWRJ?5Z\)6P]>B]e+3V,Zd
=])7JAb)2N##4XXEPHaZ)d)dFRM?B5N4,d7NL]<bG3P42L2d[CJM[f6_)9T5eB/O
0#UKKd_=Z##-G(bQZ^PQRWPO&<A(>>d:62)NR1.A9OH_[g\WU5S\RO]]F:GL5a>S
8ARR8C&QS==Y3cZ=;K9C-f3EJP81V#7I_LZ0B&Q=.L&e^4@7&-RMM(5#<I\ER38f
FHOK4VFJR@E1QK58E=#K-RGU#N/]ReHJS\H_1UbeE(e1dAe4]MaNEE84I=P#VQcE
[cGXR0e5fLJbc8KPN7?FMa-JIKUgQ>0e>5-B+T-geEO:Y0#P.]FG0OR/TNRdaY\B
]cZC.[F?4V+DZ-\7GD,;HZ9YN)dLV^PVMR^<ba1[a),THZ;6GLA.IMM&4+JDb#M8
e0UBU-EWL864[]df>=[P[5ZE<H;ZP1([FW/ObQI(XLEBaREBKE8gN-OJP;B?-G3P
]MTUCM):2bB]Y<1c-DLB4)OJ3;?+FDIMY1Y,_K98QbO8;Z+99De^OLY7f=^eDJC:
OI=H>;QFe[\>bT2R)SYT9+S52L3UC4W7M7&P)>\]WQ#)<-:>R7B->7AUI_-QSPNU
8/EI@U4<,T:+ZJM[/+B&K)9#O;A=K;Q@Df9D,10C_BR;RB.7?O[RD<P+L3P5bW=M
#2)P/]/eNN7aLK&Yd9fTaY5/TT,KZ]QC2R?[f1db==VL#CH-@>=.Q<c05UagX?@Q
S0K^])&4gN5/VCBg+FNQ^@=CO-P>49-FC[(M^&_R>RUZ/G9a\Z_I#6\O;9X,g]8B
9@A160LdKC@FcNIG8Q.8G(2YE:b#9=QY;-/\Og@;P\#Q#;E1.R678DHJ6E>C_6c6
G;aO(G2H&LAO:K)2TYeFNOYbfL##PFQOIO&.W<I0(K_<A5&P@NFUOXI@MCPBc\X^
J(_<4->PB2<1KUWT_A,&b).gJ,YbN<\/-cWc8g,3.QHJDG].?EPKK:5\RQJ9;X#6
c#:M/Z^@Y7Y\KMg^Y;;O8bdT]^G\Ab(6Ga9-80eQ+(206\JX^gITAL]CE(^>\bQX
I(AM5G>LUOC[I2(?dGg/Bf]379(7RH;P>bd3LNCLb>HbD_J[HaGG5E2V>/8+9L8L
Z=CFJ#J&S#b=(aF<[cg^:HfTQYNcFE.[/b=Y.91+Pd^5N.5R5[BR4^>KO((XRe8?
GTEUUA;ZZK1#&QF-P-(2[_\b5)BM_2-_gM;2_?C(G8<TUY85N;-1O\CM(BdSQ3C1
5@_3geHJA4O?2BD3T]X[J7>(>?]#ZF3KH^J82[BPT9gZ/;K4J3.=L@Q@6]/4HPLb
GMeNd+:T2<3&HR1EL4SRBT.93(V/NKC:Q]cQCGNab3P^6?W0?T:E<Fb?87I+aIEZ
<MKAK?200FGS-IK0DUX1#G@8ZK77>\^7e]+BR.Q-0cc7b-f5I7e;+EE9SMc&\#:+
>^FAIT\cRQ_Nd0@EgQ@NGC8Z))(#NSS99#f>Ie,@SBfXZ.X@P](PYcK<Z-\:(=3S
aH#fbe?EO+b&a9:bM(CEaIA:.e(gIJGQVC>Z@gfK8)9W=/,Eb3,cCS\.#9].<3)2
35Y@VEE_05PdY4@J@&X:;eDUbN2GI/E04DSP/0DS-?O?D?]ZSCVcEKYdHV[@T1X:
5ePJ6<Hd2.J+IVH]-\KKg\4+90>B7/e([:^?AK@1.IIT3R(.eHIaS&37T_JUZ5/E
>^a^FU<1>/30((H\d0).Sg1OZ7]<_,&T\)M\fA.067ZJ^Qc-?R:-R1b)JYX\f0WL
&&OfF9S)bXX;a,>Q/[S5P(]B:<dAJcPb0@)3(I?C?EK3[Z?I2:6.[R40aVC-H^RX
12^[NHCHV@B;F8U[QG&P(]5D6+E_U&N=BU>FI6DR]D)L[[+[#b3AS1GT(c9HQJ,1
/34Y;GEcYLD8@@VDgRBW[3fgPU@ea1.50GW?3^&C3dJ1G<YA=#PUSeTI]]8<gHU>
a\7HGCdcTCfJ?B+&4YUM5a8ZVbY6J7CZ1,2N4K+(b1e<,D]b5KDO0Q=18EQY<:6]
2RXU6ee#+1KS_T>d1/\62AbgDG?+7WB7H>1N@LXU-I:Bcd&KXG9.8X&a;>A-(A?Y
XC5V4XfgX>IOb@CcN6Kad]#gPQV/aN-,PS2Q2af0SQ7cK+e7/0\SC#\-9,<NYL?H
/1ASNDW&@Tc\Q0(^)f^ba7?>E;XgCdT(>1/JIT?XU/\aaK>)^47\1[5<PLXJQXZ.
FM=9#ZB&^1HLWB@DYYVQc-0>Tc(=2SUdD8AK#/7D>e>.SH1OEU_Ufb43604fSW5-
#KM4gg5CD\L3If,g[(^@BfS)_Y.N]NPfT43cWHCT,XZb>N=.X6Hb+De7&);-\Ua2
M^PC<[\9UFB5KV<]R7d1:\a2a/aS#gJagW/9/Z.P<N7(XEWE=41FO5E0f?F_JQC>
[EfLXEb(/Z0W(-:Q1e)W+AUFWb]Y9G68Ub&^WO]<:EBOgYN>=K2Kf9TCgT<>U0(U
a2VF5NIe3^6.8@J<@dfQ80+5BNdN@JX@DfDa0&9b#F-?Y_//GNL?QN,@:8EgLI(_
:MGB+_[\3PSDO)7P9.#gHP\BXVCLFVI#/5NR=/9bJSCY/0[bI]D\A=KQK1_8T,^Y
CYQC>@W+3CL;G.D@-^R=&..a[5#@?FSYf592#&/1QB7U#Xd4b_(C:KQ&@,>7?fZN
S9Qg5dN3E:WC._b)UO0#;a&6I8.#-<Z(-DGaX()VYC6>9g3gaXa;a)eTPTG=_[U0
.cILZEIJ&H+GdLVRYG7C#C^FWb\CFDYBC[X>ND\>6#T]=^.K+a-fMcU):cH+(W8\
JTD@8-RM:;A1D6SPMadXeHK.VQS9K])CPD-I4W^KP,g6=<-#[Q.SHH^PUXF6c==.
JVZDKU+8fFWaRYH3MSJ-^,gZb(aP?;@(FEX2)g@f;R]g5J.d\PL4H\LABUH9]K_9
HPN#GUFAXC#RD^Rc:YEgI&9?E/5=:KM/0Q6HQa,8LUU2-JKd5E0eIg9c8C:[/E[@
&Vb,-AbH9IeJ0a:WfMK&PDPJAXR3[TY\B]KQ[Q40_&8dXQ?BSg\<9eO+]<#TK3EZ
H61(DO,\L?9A8F&-ZJ\0bAVOLfd](=g#]]ac@,R_G#48TP@2@C@0S^>WM.LZ;8.3
OJEQ+/a;U^Q)-.X[7;;P:Kc4EMW>O3/7P-a8B>,G^B:E]LXHA-F1RFP[15RbH]J@
b6\egXI\bD;Tc04D]0a.=F1GJ=ABcWGINTNQ:D-4I(XTUN)J_=+E32ee[/eaEME(
,/IRYad]<DNf/_fcG:.4\#LZ.g&^1+G+DA723-XEb8_5;cbb,:8O9<_UCV-=A\7<
B9[Sccd_Y.ZP9&C=Z[dZ2g07Hc7Z[.+:<-5<//d-f9//93bX(4J6K\eV4]AI3I<X
U,\_]3bL(2B3?J->_)++T<0SJbb)2<OQBg_[?I5EJGgAVDFO^S=5)VT(1(G&F7,#
#G\-S;OM:(gDZ]aVbF\K5[]&+.LY80K86@,OK5<fWE)[a5S&7>;AXM5Z?4_=WQMg
@7cGTJ3SIK&UF.S/Z>GJUHcA1QDZ>Q&#Ig#Pg2ZLZNE8cJ#Y^5gGL;=>eCB?]@K9
g<7Sg.2XC9&f6[d[,,<E(+37=c[-6ICYGc5bVYNa(eS66]QG<fC=gW3ZL@Wf_(;=
dK]]L7IQ#3-AMOQE\7Hd#06IQJ7[eUe/[W68g,O0):G(^7R^#F?5RXNLH#[<)e4,
O_K.bQaS=N#4cW.T7.QeG9,82]A1?eP]0C5QRQ)>(0GB5YMDLZ__BC]8<cAZNW+7
5^L(F5G752b)^4g_OcDb)EKKJV_?7X)62PO_Wa/289gF#.dOZMP7.+Q_+YG[F#DS
7#bYXV5R&YB=^:-(Kf\,aI,(-:B#^(0_fWR..ZLgX?/GEEE#A78bDf@ER3L>Kba5
b?4BVIL:#G./QBL;K]^C7^Bb#eP?@M,W<+/\SK?]09g7-:>L6>.AgUOC,)2/HOM+
7A46XI&N=[f^.;b,\)a#+DR\#/BU2CIC71FHN:_dbSJBK].41N?;TKd\0R7DS=2H
4K2gZ=A;f)\U^.;M.EO2e+Ia:FJ6T2Fd(1.<,/g+?)AbZ[W>N6G+\:D3A237b:HZ
d-9LM8K(L:8INU#Xe#,#c+G+0(R#ZG\?.(=(fA-:#7I4F<c_^_U)LAHV=9WP)ALP
=g@RVVCIdYW0C5=78VcUZU,.PLU:NePF6fT88L75GR(cOD<b^3c3La<>4^=;CM\^
KRQW^^I;U[#Qb74>g20UVgZUUTfg#0Y+F3(VQ(VZ=W\GAY1fL@e(7OS9F_A439E4
+-QFT&?-1e)F=/?MH(F(<eS3UIQAdJ)ZM+2^Ac:&8>^U56#JgYBVM?<DZf6c59LQ
dD5<aAE\H5M:-+37[TXVdU^f6\bJOL:#X_.>J-K^c\XH/8V5>3K[>)T,TZ;_)2EX
PKHJZW1aRgJf:O;P.<B^K^C//NW+CcGQ=-CQ7+8S[DJW@_+3=KR<:44IQBW](1A:
f.\T^_IcO>cJ.-86QdJg5^P+&-L[/SLHSY_dTSdJ-I&S<+VM?e1(L)JBgN[P-4:R
)@-5X7Z0V83Y0R+FR5YLa=R?9,T(2&EMcUO[GU39a,C;/,7gNHBBVKKOUGf[D.T8
9SZS?6+3=gM/F7[2QRM]^fOUBZc@e]<8LTb[WC#]N))X>R<8]e>JE2AG^._WG<LB
>4FRW/KcXCg<PK(Z\S]P_aNY8,>05eI5^2T[5g_W&a7=0NNL>+eA4+BOFZ.EHfD4
H[HY-5MaUX)<Y_;(Xf]#Y;7IN17&8:I8G_KN+1#-P[IEWJE21A;\J\<1&&HHe;Q&
:<JYc[5JSBZRQa2gc^#:I5,[>BTY(+52U7YD.eY;=KGAA;Uf3#G;SQ.TC&Z8T,9#
=b,]:V7:_f516:5d2f?g)1GP_:\FNTS^T-E82d@H0\H(FHV1gg?2_>Y+&XQ29ELI
Vd8,>3UK7c4\7N(8U1<N[E\]_N?0NV(5^bR2DdEHQ?Q+@Xa3/f7-@,X<-DSV&3a/
<Q>W/.eW^]BXJ37Y-JeWUeU1K]c=<HVB0B@\P9&6JK4#<CDeb4HA,ATf][eSfIYg
Mc8&#H1DU&YcNec@;#eaQ(Re@?P<^?6_R\T]a8O4KCKaZ)F,[-Fg,I:EHd_O.bf7
.?R_-CA]8<;BN=7f\@K/-\6I\XPKRFFLaF>L)2O_@eaQ=)Jb&5fYT0JO^F&.<?A-
E=KLgY;LIUMZ@fU1=aa5H@7P&NY^L7+E17Tc8+4R;WeY>1Td.^6(:\FVN5ZaKMNa
4.P/(LUY6@[+3@]gJ8<S.SG;LP=;+ZD?N,?(BJA7RYLZ:-2cR=J#618J8J&_B2Q<
NHb>;B63cNSHC#a#cgFY5FP6g38f6\G9:NG@Z>KLQ6+dHQ>0)b8=^>a&S#32aCL2
X?/WEQ(E\c<&,XQ/V4F8X3HN2e5B)AQXD(7[7aLNQ6B&+VP>#XEP2(;\cHfaV-TA
V=1<LD:G4_5Q06TOe.)S_aDN-1U_)P,^F^D1a0_dN,;V>=JF,TJ?]W1ccUGHVfdF
LPKP8V>T82,-IP-9YS=NcFQG2eC6eTb;/?2S1fE@WaVR@6P10ACVE5\RQ/?G65ZZ
DZfL?8YbE-6[gTRMF3TGX/QVA9cb>-?6)&;<YZIKREF4AUed>dd\LfLS>0;(M2(0
M.6++@MP,M=P:1-5R51c^T67.),F#FPQIH^C6-4;M1@B2^B8Tg\.S3#(FRSM?KP1
+Ie9M=bQBefUe8VcC/b2&6.YPCCZL9#69X_UM+AGL(4L)XaNd7AD:6g;eM:3[9Ub
#K:TZZ\&[2F231#,f_L0.P4#N4^72]6,eaXcIXdeG\>4,bKB<:b:S.#PRKDO^1Te
1WQ)M0eBIadBb+YEbfT.D>f/+NZBSM1f:X5)/+fCN>>fB16V>Se;>F@.#JOOERUG
bb8YbHI790QU]ZN0KQ;VX77/R(U43(8PR=65+9@+:YL(V1(O5W#/d7=V?\0g7W2]
(2W,5+&F2a-cZWUE:(21UNKPMd]:E3^:fJA:\,b0AO2e_+7^cWIKX.^<gCV8<JJO
Q]4DE?HY@-6SCNaKUML7E3FDS)X3G1Ff]>8)Z+0/Q:cDB/4_L\c>TNU1)W1BfgJc
3Q0<?#=4aN>N77(2H9WUXW^NGeTAJZ#8X1[K;Rf/0_&d>[Ge[5+&#5gGMR,]?HBP
&B:1GEG^FML<D4U&DdeDY3YF<a[0XIM@M;386YNa9].e5#0\DQQ<6.cEXCAG+eK7
<9_>P@:M,aS6Ba:G^ON=3fV\PB\dR;#,[9H[Fc4MBbbQBZK_f#37Vd90=J&K563_
>Z1O0Se,(LXc[8XOE+HFJTSaJ/,4X.[#@<GP^<3b-e\I6BW;&E?]VEdYRN_/&3X8
28=8H<.g5FKcYL(E]@83-(a8aaS-OKHX@S3F3D@<.bBZ\DWA=LJ)HfP52A44<:4U
0VdTZ/7:BLSeeMC<Z.0MPcXEgTc-N/-(7RWeM[H.c+b,Q3_DS120JPZb978+a&aV
J+P2ESO>?9WZL-B[XO,[gGHFC.]C>?d:K>gO40a?VdfYN<3MQJEgJ#VNa)WDSF.)
_MN;@4D:-7G0(JaBM,SM8C1)>8a?&3]S#8B:A[UNQMX?;\?IM,gcRWAYX#3W=H?]
Y=V0:;fVW\B-VbIF2:I&0cQgE(;[:#B?8\7ADU,^;.K&#.@bQHTL^Z)a?6\6PXc4
A#ee>7&g>\#;2+;C>-+&AcD4^^>R9;9Y\a3PHX1@S(c;-O)/7NTXPT>0g#HY6U:d
Ya25\d(7>14N@^^YgA>?1NUaI=OS^D/A-:GH0^_AFFY4>/f-Y5^VecSNZBeD=Wb[
G-NabfQFZTF13./(_+[28W/>Rb^#Sf2I,C(LM#ad.A>E:J>VVBFeJd4NXO:A1E()
//BR6+H+BZYbX[4;c429PSEU#=XJP\E[,JLKWSfJU^L]X1M+XR]aVAR.:A;@:QcL
V.RM?Q^P;;F)S;7_H1_+=gc;4.>58b[9AJ<\ZNC-aIZT2,Mg@GQbb_YJ>_^Je,OS
D/Ngd0d;Q:M@/ACcWKCCa:dM[;<E:-fddaG5E2O[5+6Nag3(]JZKX3G6TPF5]/S\
S3eD^RT1Y/LB9Of^.\b:S9KAT-)X4eT07:8OT1CUX4a&2/9P,#&cU:I:&.)QQE=M
>:RF3DCJaAf1DMYKDMdUJ1dWb87[OGI])S)^FIRE<Ec1aN=75DA56gD,R)@N[ZX=
5DaZ1>KY9Qe1L<))fOJS.7#9+^NfUV(c4G?JB462<12?W4/a.SM8QIS\YT6bNCb>
+:8SZF]M-ZQRNJDZCQW#2=e\YYWL/V?6PM+40dY@;<:@)B-Ba1KYRETY5.P&HfX:
MGI.2Y9QL#TR9>]Ia_9D#JOM7fEOb2f:Z4b>X96RRA6^6H(,C0Q+TZ=9a\6aXg-R
>22..-WP&=0K)F\_+N[_-L&,74;;/4bYRC9&F]UO^=^c:;13^RdA,Ga5?eS^5M5>
MaWe[EDSA\OV(MK1D0Q+L;9BZU\-.6aWM#;.\9dO7UNf<a-A=<gNR)GQbUUdQR@#
5XHA_b6^O7OPS,21@)Y;K:-Z=\;BDWdBLFU]0,)L9R(,05aJRME?78OG+gM65DYY
MQ2V]1FB1&4G[=#cGT2TKBZGO(^F_O)M4(c\U=55.R:&O4UDgCc4KFMX<-g9G(37
0^O5.<W-ZR##H\I4PcQ>KO4UfYISe#83d.E<6U&N4O;S@F6eZL1/[Wf&)M>,MOFT
#K[@.SA,(-6K:K7;ML?d/M.\Y=+7-]6X#(d8V8/D_D#T03.XUZZ8.SVHV:[@Z>Ke
Z&b&06D_>X+_J,+LU?&dT7SK)VFD-OVHWd/Of9\QN_VHH\WSd3>+)c037IQc8AbQ
UF88T1Of/3;PTQ:ZdL(MCY/-=4B0P6ZN;_ZT]d82),<RW[efY7Sf:-HQJQA^8gUI
=M_A<\]6]S2D1PMOHR_@^b]P<UD)3BZ53c;0Cd8#25+:GIMNT]\KZQE46d=.2A@O
RK-.338SF0[GV^YY]KKKJGYG7_8_[:KR0H4@#(S4@1V6=(V^a:MD;@,8/I\<Z8c,
.1U+8S:W)eJ1)@a4/d\bGUU&YQ:3UDJdAY+;2Q;XEPL[OOC\XK.L9U6M)X?=G-=K
2#&T8OBQd;_g=12+(TJSN7)9K7<N3\RCRfW<6\MG;J.<C-Fg][S8CN4D2e?AJZOQ
cc<+I+W421K)Ye/DeGc17E^X(C(?XdYO1VgKU4\6;[+CWg1TBXg&g2,;,^X0f\=c
#SKOUfO9c0L&X]<-JBB<=&Y[>-H:\0cL&@f4P;ca>\Vc-@XKMDW;gb6J3?=eEdF[
O&bH&GeP18K\::75<JE8a27@8P@X?UgXd_Fb#E8TW0cT\._dY[;?:46=SO8U8U>>
^8PD1Q8TbG/<;\OC)]IPUaKH\\Wf2;D#b2LaY/c<^,WSSP2+Bg-f5=P4)DC:,N9b
d:9M#;=YSHUfFU#J27B&A4eXIf@OAZNCW]LQ\CL\b\E_G6e&P9g&]S#JSLIMGY,P
ZB<FK\?]bHe1:B/RLSEg5dYa;3bX#9?RF^J&;V&E-UEb9>EDI9Sd3@\,.A7CW1#/
.R4Y_E\CECY3f]1b2;02HZEP>USG@N0)=P@dgDR=];\^Feg)3(+\#d#GQ5bRI/S=
19?<Q&<O0:B\.Df\7DQg2g-6S<[A9QY<fG\fLXVL]&4JMQ]CJcAFgX)3?=bHa\e?
3,fEB#L?][,E=:BWQ>Q12]FT0F@Tc6LFHC>]<Z\<\Fc5E8359[.\ZaATG_ASNLdW
W9+_M;A@UbHKLI0Y^7+O^=I+O;\,77B@0(L?RW1I@PPG_HYULdReJYIM<UR/)I.D
5?.JG(Y.LVQ&1C.J05U3dc]MPU\Z5/(0.WS8]bX[>6BAV/D&0<\5RE8OJH<EVTX>
)Kb6PeO7X+D(^G,=\&#8-2NJ^F/&/\@4:1RW/&H;A@:dV[WW.-(f2,E5C8G<.4;#
K]4\46AM&FabB\ZUW@KJ]WY)CFHU^0-V0?FY((@&c\Cc^de+2dMUd;SP&IR/-WD@
/ObDCHHY9d+QBeRSF4bgY[c7G&UO#T?):C\gXC,KBU#N3,P>7)?N4N+b:OL1B1.M
5fd,B<RPB.SZOCT8S0S;[dgGHb2/N,5=Z808:Z^dg,_K=H+;82(SB@b)8@WccFD>
VFMg0+HAR3@VP^A5?K.K0SB<#OZT_>R[CKe0.AXF1?=V9c:8:c7U&<0a=]R5GX:5
3A^T5>S?>^6SURZQ3\NP0\bDU:/dA]e8CB)bJfgb2&/M)K4WL.>#ZO]\]ZOE#]-X
OCB.&VT#4d;.:4DQM9W<a#X2@KL1FM=UGEDLP+A4,1?-2G.G_NdBFHGeCff5K[cP
=+\AV)3CVa,;NHRDgXS5VS.V.dHX<5fc;L2S)=_g<I3Pf=<cQ]C@aJXN>(?eCcfL
ERRg&XE4]3+e0B<f3TbE,7877#0^a.#H^Af>HH)cVLXcA[HSHL##9PG6A)6]@>70
\4]V3(M]MY:91Vd6b^8>VYCI^3IVTVBE1Ma,0(4LA6M3HO?eJ[e]0?=-NACc;VE^
.2.?M48L2#?J)=02Ga5)>8KOOg-OM/b0CbC+R+#Q\aZ5b4Lb3-Fag=NN=._1TGAO
PFE+a:K8?17@6Z9LSC=UKQP:bG,S[[U@O&9F>,P:&E,RP>TOFI+O2Q8&5O]F1)GS
bF=+)_cgf_b\Ia@A/:DD9:Z-/bM)AK>Qe^<a>=6&cEbV3?3(BZES7(N;;.LDVA81
9^^[0f@g(2E1N7.UHAd_R[R/#aQ]?cRaSRcR=KZ>H2JEX8I&VTLE(M-LbQa:#@/,
O7[@6Q+&O4//CA?MQUTgQ@JcC(PNbI-N:]d9e1Q]CVLWC<)KT.66FO.dA?WJ\EaZ
IRb#HHdd/-#R:;NaY.VUP(.W/<g9g8bODQM@&)6#:Z3X:M4S/EO.W/W\_W=OUXa+
B2GLL@Pg3Uc/1Z;Q:17Y(K#g)3gO,FHFH7J5RE<G<RMF[YWAZ\T+dHHZb>&=QIPM
3Q45JIVRfB_G5Jg#^[F1?dV]RNKc4bc?dgN\5>G0OAS^a2a,=\0G^<HM(gIa.G8T
,NfdQHO=UBa2FSH]KE59SFBX4Y)-OB2YfVOOV0c?2><IXC;Ef/2Z:C8DAJM=7PLb
M668/Q+K5F@I:99S<C>d.&+F2Sg<=^3/=[K(RcBQST3NXKg-)V?5.f>@d0A=^7bP
(&9AFIb?5;^K=f9T<bSbMbA.XBZ>[NdC;)1B=gPY0#RYL7,(-8@>Y#aQL^=KcG@1
SP,H/cL8+KH4/5[-f]8A[)2:Q+?@.&/?8Og0AK83MOBX\b-S&@#(VE?:2YWD1R]L
ZG1MKJI^E=_?@^3,_C0PWMFI69TLa<b?6&eY87G[IfSJ:;,MH4)K[;1]X:Y2W+U.
ZD.L;56_G@a[MC/B/GW=bM3@(H03APR?HbTd8[8>)004-aFIfbP;c5PAb\Y1H>/I
^7aR8.WS4I<D4(3&W^G.Z^Y>ab,#-V)-Hc7T</AK]BNL.3c\BJO7gK,4^f/2:@P)
R:b&d9DgI@3b><C4^5O[1J06I5#F^LU<I9\):RWRd9D/\f2@?J[faO#Z49\Fd?M_
_#9Aa,F=dE;Q2&R+Z8/SC1B2-CGdGTG>NeS_#3(KYI\5R4deUBWC]=3UR(S[FWDa
G5@FPLR6b[,OJ1C9E<b8a^7(fP5FRT?4.D-bE]/T(7)DGM[,ZI>A?g,)1U5D0E,\
M0cdg0)cS+BJPd\(S2[,Q/6:g-e#)E1Ig#>(ee>L@X5Rd]>=GNV9-aX\X;5/)86J
HVG/+JU#a4VMJ42_>7eVWaP1K/aRaLOS&1H=5DB<51Pfd,>3V9H+F:,)5J.12egV
7f0cX32GVNPa<Kf<#)HL\bOGab7:,Z/R[M6W^QdJ]HT,DJNa3Q2O]XLACXA><ef4
89RZPU;(WQfZb\V._Fe;/]8?[A\-BSf,HE^8BUX8ZJ[VJKD,J.()5B)b.\)b5L>W
L)>3RgGZ;c([Z:I3)1L;g&ACCSKUBC\8\fVY7<X+/[2S>I7&^?6]BJB--&;]eGBR
EQb(-O199Ka;EK6#fS6:>89T_DRW\7/WQ=N[a02(1ZW]?:J56E];.bS5fS]Z0<#(
R>\_HERb&TACb]C\a#Tg@SQVaIgO[I=4D?a+_g:D8KdO@JXa4adb+EYb-SE;=<RT
&&T;)eM#7)K5&\IO2Ma0V2EGgC--N4U=.,g/;5Lg+faZ>7/8YY>Lb9OK_>VQ7ZY7
2&]^E0,T4f0Bb97a4T_BM45Fd&A99)Y8IHR647W+B/8>J1e+M9-I#:.2P/H.ZPS,
_&2558dbE4VY9F)3K45YQI?3IDeC4#3R5-d-LWb.UEVHc4[]Db7b5;Gc/TaVLT8:
&;NgZPM4H0J5_RW#O&U.N8e2:P?5NY7MfUXSa?,30b.JB(c.eN;NgBYP+N7\8,-X
#UK,]C,O]E73)E<fM]KIbNF#):S0M1E=Ca@4^0D==[Wf7RJKfFGdVRI;5RDFB<:5
QXZANQ^Vb,>SGE&7>&2_^(E]:C>3G7@UI3)F99=0CM^N0X,g<;4HFaf=a.W5/+?,
5Q]=.?RdQ<g\=3/[30[_+T/?8>@IASY_1V&\S]ZM>[(M7V0+SKXc.@G/b^^-71A)
QceQ?aW)27=FRHXCB717EH,W:X9(a<2ePY<2<AFRQ[U7,(&@U,I/>5,-L+Qf0>[0
J5?E]1a<7LYX8704LgMb49c-5KJM;bXBefTPG\4VQ9R;2CYH8ZR_#FgE[JcD?H_&
4L[:E)g^_240N_L6=<8;FKU[E?b)6D0Z4J8f8/TF<N/09,_U?Va;N,_GYg3CI2\Z
#/P??+S^-[]2J?U4<BJ5@XOH53Vc;+LES#U6g7(@2_I5-6=2J,PR[_1,gc.eJ1U\
9L:1PX:_C\KQZ&#Of^&^f\DL+:OABd1WD.199,CA9A;[4[[RT2f^?+JRdKAFI,f8
<J^AR>V:+&)TQ?^6R+[([K;ZL./H>U7WBIXK[-C(Ye(850>H_gLc#J@<JfYHfS>@
B#3&C^5L<6#+:3XK[34(T+;_Y09.+?FL0(2NHX2Y3\(cWd[T,\&-^8J)IE/Z7@M]
Y3Z52FXV73/H0b+GVG>a9MWH35E1>A)27U.caI+10.N>XOTMC([b4S)24[D/8FDZ
F543L-=7PZL,Z>J.3>g671Q.?VV;5^U5BDMVCb]NKKA5RU/ZCZ.2JG3#LR>+QT05
O?:QU@U0Y0SQdO0]aF#dFJANIPYF7+GKK#K6Z@4=b1H3#DQ_35:O_@.8DQPSGF&(
A4,,R73\H3I>?5D@dH-7e:HY#B5_VeGSf<HGgY?eJ>#f^C,62DBLP^M6LKWIa6:P
LLF]XWB2#ZPeBcIJ]fb[UI9G7ac69KKEX55?U@^3]Lg>2+BQZNW@8c7XgV=),9.5
G=Icd;T6B\RK+g5cE[7=53@I.S&c_-QFVb_VL:5N3)5?WX1W5KTQB08Q)T<;H5[,
=bL=[CdL[WEdgbYB73AO4#8N_Z<SE/R#1bPGOeFH&TcKgORdRb:<f7RF643+)gHE
7Q=bG18KTQ6C?PBSfJJbdJY7(,#f=>.^_Y5[/40@?)EF8[7fB?HVNCETcV;&@<Af
[8,Ic\PVc;KHf+KgC;<9d/?#E7PZC;R?6CQ1W?;8#(\,fFc/:.LGBcG@-6]-G?+I
LA/)Y[fbQ^NN3YJ=+^-Y+Iaf;SP=@P7,G=2)Y4UCIODOUPZeW^:@T2<N1>cHRf<B
9Ka]=JO)4.afGPFC^<MR?WW?+8+gTUYcS,CG<Y6B,aJCC51A4TG]85fA+HdBcRK4
AQ&P7c5e0W2deK\6[9=QT@\:SVe@X#->@NKcdLKGW&ZDXeRO[EF^M\F_0X8_X:b@
P;0SKGC8d--b/TK(d(6L0dIBV,=.=Qe/F,Z?a&/dC-_bAA006^P[5c3D1ST9-#,0
WSM[I<2-MA(g?>CTC#XB[d/2K=HBVX0d954H(gR9><?4cKY8<E.HF.>?cEIW17Da
;?#?629::5D11,MYRFHN8ZaHNJ\c+<HfTg8Dc<D8,IIQ0OR>@<ARVPFS\Y+PIg>,
HWc>/46NVGSY_N]PCGXY[Y_:TLK2#A^/+&2,#04._+Q&Jc:\3BeNYIP+ceB3&/_=
JMO>a&S-7D1]EW[,5/IU=YV>b)R-FEFV+D@He>b&6[P[0a9c[C@d##VFVaU8O4X?
G)][Ke1JA(X#/E&<\1#P?>f;VWJ==3d(Q:dB5+B8D9/&?/=VUL<0.X]NM1U-@e)S
9HTL9[5_5ba44_J2W-OML?bD\:#(-8A]PT&[,S9F;W-+VZWU_MR(.I=3)VZNL;SW
U<G9BE[?=A8L>=HgUM_0<A.L<),/V]IR,.#(Y>#O,6>:-+@aKDZO\gWeddcfD2#Q
EdI7d,SOQC;eSNCLZXdFP.[#0c\7I<S[X;bLDS2C,R.dPg9>9LYTd1DQ4M9NC3Wa
Z.KL8e51TgQM))e>IC3:MY&:,dP#Lg(-Q4>(3U0aC+He=\Q/1;BRe2&H^@1-J8T1
=eK_S5W[/^3]:CCVaWcN[JdNCB?VaNEG^0)\XIO[60@#/IJ=d_fS24b2<MbOP[<-
-ZPG28gdG_+A(f#O?(Xg(fbZY,OPcW2(EJ:#9#C#X0>&Z@EF(g_\a?gb7?.,Z/bY
M[W_JR4YO#7RKXJ05;Da0c&e8[2<UIQH[#S)=#N5J2e4/9)G^^Z.B^8XD:>80aOd
CLLa:7:dc&OJDYR?Ga5[Z#?cYZKIQ>XR<(T9XI>HQB&bId2VPG70D2[V3Ig.YH6d
&)Ad.7M25U-LF[XN75L;RLW5\>6^1GF0&TZS8B]d5DI<)D>2@\[9_&=BG=S_)\[a
5JS\BH#5b+@HOF3?Y?W3O]4JKYd3bA849&e2eB&P1bAPQR4_0/CEFT9HM:D[[S)5
BFDU-04aC@YeM2bc^K^VT=6_)@5(e2C^XWUE=6]9/GR/7AAE6M#:_F<dU2Qae;[-
;3[1;GCF]#&JDWEKZ@CJb9d9eIa,6POTJM6..GG/bQV#c<3\a)BACF)YL=g8L^5>
e59R-?_QB7e)5I.fTOT+=&MIG^EK;O;Dc<4++&OBg+M4YQ:?.?a[J4Re#3JXO?U[
ES-S<:Lb>:DC+1DL&MF+GJW)<&K;]QN#UbK]Qg&=HSL,?aQX_;,.F_X^#(W1[CJ]
A=RcW[)E7DaD^0/Ra>-(0d&//gM^g_.P_O,PgFg[@3HfN:E^T?ZXdIGGS<b0bX#e
Q=>W5#JUX5g)?@WM>3CLT&(cH[g(\6IPa;TE--SaT#5SHPAeEOK-O;K,_4e)DDH/
A68K0I47HF,>_T4Q:F&)9(9;&f[1W--@D]C.QY9]E>9X3V9[4W:+<UdYAZ0WV/_4
#B0e7SK?bA>DMcH;X+Of&d5?,B8(5Jd1\TW&PF;cf++WV_GF+UT_0YM,T,_--Fa)
Z8WFKA55UP.P-VV/A=T6TK^fB:A4129\]HSc.Q@3^&Y3<TASYa8M^/b2>[B]V3W#
27&X\a8YQUYOEEZ[ORPLES;R:J?e\;48AId(>HT7PV507Se@?7>;R:P1SF;g--EW
/_g_5C/22A_Od8-HEWY&c8YR,(JE)&[AQB88<25T[T-N[/6F\33[4H0-&fEIB8>@
?e2,adIfSc+F,^G].-L=b(5Y8K8gW<^,YeB>M\A.I)fNd0C2/ARMFT=dE_F8WE+f
UE3W(@9.F+^FB=JRfe8Ha:SJYT?>=15F;g[MN2_YMP7)@D6+;_._8_58If\\B@b1
-DDT-Q5&BR6EFd01K60KVU=KbBE<<5-\=?D_QNCD@^.S8]BCaBQ4CJEX(JQ:6K4?
24P<\)=@B;AC3>--Y(PW\N5R(+G3M)P,_Y>+_C^X+dg<W(EA=.1MTHZE_I46W5XC
HaRB+H&IOTJ6SX7L:7VFd#J.7@A9(LJ1^NM4=B4=9+&gZP@4#K:7ZMK4ECIP+KS8
CWdZ:)gRI65;Rca)a3Z,c#KJHaTR[5-f1FcKbY3NJ^.UV3(9,3/#8PML02(CE2bQ
Wa=65,;=S(b)Ib56\9B?,3=.RYISYKQ>5YN_f^?e>/J7VGS:?cI?HCO>aP6OZU=_
<GMQMI?BEA5VC,>A9?D@DI3URV-(W+MbVQ,U5PA7@MP^F7\[DDGU2DH/U&[TV;SO
^I+/@egMKR<&.4_:/5M&7b?Q1,d#7Ja=6Me.A4/;&FIII;]99KK[JCKPYT+97\@.
NI+X@eL&&KM1KQL#L43N@g@=FB4WaX&=T6.F__C5(cKR=]SX03]c?V:NEP,9@VUR
<3f+.OKVV2\e+(cY(73W?@5E0SV#7Q-cOJ2-.KdKNa;^,W\Y,T?2.YJSA;d3E5QC
95cA+H_a<bCWfQ/Lda&5T8dg3M2GB4-]\9gV8@ZFcaNU.:[\P=F2WDf7V##..9:0
J6N7C\ZTPRc]?TAc)RBLR4A>3G[W;5N4?aJHTWJVVS#RCMe1>W#5VfYXPMf#LA9g
M2)KU(53@bQYT>b8LPL<EcL4PC:f:]UaI_#I,F#(@E0N#;eb>NY(SKERNY:VEg@]
)PV^O1=_gBC+Q\,EaN,]d3O]#C6-W-+8ZTF45e1G[J>Q/>J/>:f/f7YB=KK0/,TP
D(^PI+1b?XA4-cHaG2Z5;BD>e[2Og87O;eJ0Z<)5[0AL#VAUMWE8d^I(^KN_WLYU
H>a1QA-I+\HTZ+QYLY,Y3:TIZA/F?>LS2PfX^<TaRG>T:,:/XNRT.DC_^8^XN##:
61=OI<2dQPC=7S/>/>#3(Ua<c+CWJ14-;eg>E)8SfYgK/QB0c.7e3>XLb)fM?Xgf
D=V\;+69KcW7_)S+\<A.,T48dAP0;G\V.g=);&TH_?73]]U4<?HT/1?\6\g;WC2\
aB]\JWCeSTUS#[M>;:MRAL:W/Bd/C+#0;83d),.GM+5fKW6ZBR]?[9A47294Ea<;
F(;&UMZ/?6=PcgNY8d<d=BF00#63U,(&=D57OeSN]&DIN.N+93Dg>Z3PO?L5MSZg
?S6OYbO.agNd_X<.-dQ2e=[5&fU#FC.K&df88;fbCZ[_Fd87?e_W?#\eW6M1XHVJ
:I,I+?8,f2TP:9+JB2PHWNNa1()TM@LMZ/;]G>V-^RUS<bgcP@^HJg<+-WH?N_,=
+d\O[[>JZ]AC2L^g]R9X3C?());,[7GTK_BO,-.EQ#08/?e,03W#;^M9<FU9#&aJ
Q:TCEHIK7OH#8AQQR;f3:[ZObg^^5AbaOLW>(bC8Z-:JO3_d<65W_9THT79VND=L
IY^;2AJ_T\fdNT>N5fMA0]MYfZ-7V3aU/De37^Ug>FJ00aee5[M740.,H9eTK[7;
E5<QST3/fEW0+6b9d-1Z=QA[9]4=B5F^71f;Y?gW<V^VVY:aAG>&Le.(4E#<9W5R
aOZVC.=8Bf1?:4\S5&][fXS,N&c+?gQYF:I<5T3,JA:Z[aD2H)^FFGcFX=#.H5I/
5C3X>,+7-9;P\8K>(>9XHFe?RD]UWC&99RM(^_L#e,J<J]=gfZR1bG[S@S0F0P^H
Ig^1>0R<,bO[f?fC2QQSKIN.OQfc?V\+X^+bHdO\4/-Gef=^2(:ee?RE]E0PI77#
DYb^=8\.D]40BY<K:Bed]IJN/NRB+,S16\(cM167Vc\AO;d\A96?Vc:4(MH9.e.E
B(N_(:G-KfN9AMT@]VN=g.4#]^T,R.:cfL>2=_PTAd&/KCKNaf(8R#F=>M2aUPFN
=/gPPB\=b5c2Sg<K\OZBQ[T4#T_6<MT_;dH^HSWcb=<e[[[#4V)[U7R^/16F.X,/
CUI/KD9GdVD,CGUXFb0<0+H6d35X9d2CcbEEf-F0a6bVAb>I^]ET0(ab-I_3c5??
JfFIL]fRb29dU2FU&ORVCD/-=:S53g\@ZR=T@FU/06a=5I;^T:#AYfRTR:IS.)2C
6W.4XU#\F\M3X+AdAMNecL2FVD)9;#UA&Lc#eMg.CZ7V27EH=+#&b&Ed;:/:@?UX
2K2K83QT\W/c1e7ZE>#JGARgL.dZS7Jc^F1B&d(8f5&<U-[31be4UI2.eC8E-f&<
>2:8dXP5VC:\)#c:5AJ4&b?gbD=ef=4K;GU1cK6,(aV8S:afUUe@K(&d-CJ2CGR3
V<CX#&NFUKF6G_a/+5ZN\fGT.>F@e:<25d0_]KDe9e3-IH@&P^REU5dW()/fGY&V
83K<NLgZ6.&07C?BQ60KMXLF[NAPL+JI:D3@WS&LeRIfL^g?2[T&U?T76aTV]a_M
<+eSeb4&N=d&MLcB<0,KZcE(D/Pe\c)U@@Nb]dR+;SKfP&^+R@0:P8KTPNf7aNK-
EMCfb_26W;D5Q(-JKDM@LMTbN.COABJDD@6)_0O[0Y>?[d;O@.cdMX&:FccFHQHI
.U/1Q\MI]7PI08HE1BCV)9A;4/gBILS71++H^_^JdJBf9=3JDEI[9M:;49CX2OT/
@Gb<31LLM#Z5ZZYM,#1B/4EeHg&Y6K_P9b(VK=d37UfNS;F?S:SO9F,I_MA0F4DG
COd7O;G]12YN>V)bF@,(aQc_&a&-8RSdg+fA=#G[cPE10.PB4(T,]>].2f0_F&Ud
<HB;JNf[LYJ2BA6:+I]B1@4[?PJU0B8RCd)Y?G.G&3=F0=9F]647MUW-P=TBOY_f
a4L\/b\K8A5YYdD/E:D&;g-0HfY7&1Qf]1<5e@INe)/Y)^W._OOIZ=XL7^Aa&(]N
AF&Y/#3g^FEbX=2),0e9UFXOSZ;/-F14f]9a1(^eG<A7ZXSPC\F?]WET8BX-R3Q0
^&a(b>#aAAO\RY;D^BC)+cG^YEUEZK&4].(YT).RY?:gG4^^/(K?-5SBLGTVW8X:
&)Q^N8FKE=8eK\E0@^QI(JI8-I]Bc[)C^@bF1KD=(#9P5c_M;,ZM8[SeSK;ZZXPY
#01HR?4FLS,6_X3G&b0[D)+PP\8-I6>V-:+&4CUHT.TREKAVQ#,@YdSc;ZNg^ZA\
7f1QcDWS?S0f?L8ZbaKCB^NE[W4daF?/]XeCW@Q:RBgFTD+d>2>OZT4D?GK:L-9J
^)NI;=/eB[>9_9LcH))^PI30IY/2;LC^@38a?QB9.E3D7a=0067O(&@eY#G2,X[=
IP)FQSWJNYA@MBJ)IV.GN3.)@6G<?(A)C+WeCHC6)=MT0H1P@Y(.Nf51O(cQ8+Y,
33M4^<#W\eAJ[W=9B_VVKabg(-FSEGcbS&BTZ1J_&@N-0^@J9a5D+_/C:S;4)W/Q
U)[M?Z]35][Q=B3:4,02RIBgePeSK@b65FBWJ?IJMQgZ//^(@QP;.RWAc=GgbB8#
V,-9b642<Sa&;6(G[STQJQ\_Ub><UZH3;f=5P=KP2#UGRJ_Ye,\\FB/WQSE&S_==
,aV_6Oe<A]<.R2;U/2X0?#5TZZD&4Y:Z3=^T-G>MF1c[7c=JE#]):@)KB3.=GN0W
Lfb;,2/U:09TB9>LZV);]B1B3IUe@,<G-:&Z(:C7aEAD?<Fe&(6EL&ZeU@1eFIQ-
A(..?RQb5@,D^b@&5@3HI\3W#6FM<G?A4^VeXL/DQDgLf,A@&INZ@OWUE9;A31OH
4<IW6ZG@d[gO9gc2gEG_X?_3\4c4O08>-2]D[B/.7^+74+6;CVOLI+RFaO,Y>.-b
;1f+DUM>?ST5GCZEZfYEgb=;_E+5IEfZ_^DNED,ADW:Q1SOI,80e7e8RS0PdL[:C
f_NOVB8S/V:6H,RR?]9[,80YI3=GI+F^b8g<,#U\NH\AN.eQ]=d-2D6?gg^L>48\
.f1c&-:VVTN[e^RR_V_?=C9V>:(4/\JW:&SLJbHCZI1,I12C0TUQJM294P\;;MWb
AL>e0A4--P:CJd4^E:H6TfSE>1?E#fa/.Cc17OGWF&#,T/bX=)?MF,d;cM9F8CGg
BUC&_^6P42TgOCKS,I[PEdfMdUPJEA.E[#PF8<D2;8:aNT+T15]Q#Q&VF@FELbDG
:DN+U+eO8G_b;/B\MH\2FR_,X6c59e68:X(+:fdN>c/XaIR_#gc72N&_:ZK8aSML
)KLeTP2N+DY_MYTOdb:QJ3+VK1cD[@U/2Jfa<.<<Ae8\3gH3)&S4V62b1R6Y7MC<
OdIL+W_g)BPXSA7A[@ed(3YgVN]SI(W6=&WHJf#cX4J[FHR=\/F@TA.Ca=1O&44+
BQ0+W]GIBNVO5bC:c:(]4JL/L]C9[L1[:RF^Mf:;2,BX1fR>W+SA9,b;P0-P,0-+
D^(F^=GgU46(-3;c9BOc(2Bd;<^YNZZNZ8ZQF<=3](@DO?/9N#BUH+)NJ:H5R,;T
.]6(P+]]P[5XbMC5/83FM?BMI03f;F@GIM44?eB8NWZ--DWMNE7#&UVOIU@BgXd3
\G?-<BOPOP?.I=I\4XZ2=_/;NZBSaPdP)-SgU_RX#N@f<gDSVHe:[_[0=J2K^:IP
T@3aNaXB_;bV6_Z-88dBd,W.g7QQ.9f/fLCPM(J/X1^E0DILJCEU=CfB8Cb>J/eI
<?44=1X7JbDY32eK&6]G::+WPJfCV0-(WV@EP\be1J^CPZ_,D1#\fJZ+c<ecX&GS
X#&K-YYb<)d;99WX3M-ScI,a;CeTQPDZFOHG,]f:EfW=E&F#61]OfE-U5WJC2RW6
2/A,F,Z8b\:-bQ?e5.M\4E7C?:F8&-5VP](7a>eDB/(39R?C;Y^__LZZ?TMDO2VL
2S47:Z\[Q<C@-gS7UTTd#Nb&)8S9;W2OA\Yd_WUWFSde11^:J4766S:?58E@GK6S
GV1bE_e=K:UG7bXL,PF,DW9-W=K(K5LK9D\N]ZAB@3#;-de04)3;8+6)>UP5+,<U
9.(8]eN&_Z1eQJ=#JA5D4ObL+4f/fQea;gTC0F2W&effW0.5SVfeE=gdd:]&f9,U
]<faag@c;1gAFVfO/-b\<B]+Q43^Bb9V?GL.8MB9A_TMK,gW__#E8^-039L(KMdc
/Z+&\QZ05^f5X4@HP:=H.LAR]M4g&H)T):C@CQXW)eeTP[MLL31?^ge#&#aDMJ5]
XY04Y&;eFB=cTC.N-KSa(Y2f##@.d=@P;NaS0a?1NY[)9]6Je+WWGH[^]\JbERcZ
?cU<V#T/d93HUP#_,cP2?YBA2XbTVE6A&#S_N@<+_@HPH157P;Q6_S60g^egQgC:
;:aOJX-D9BYF1>:T=0N3ZU+dIc\1AX?d#c>/[Y,P,@HS5?V=&T2(.Y@>b8.K-]):
)]DdX>Y1(]8IHTGa@G13?R]=U[\FI-8\4ZG1=&_QMW+cAGPeGRVVAG(Oe3/;.F<]
9_+Y,@ZR^DSW4&[B>J]##??9#T^f&T^YbS7Y.6\#KBP;S>DV5e/,PVb.P[908(]G
0V.V:QgM0A1&aX/2AEQ>E.9M7P(1B/;Y+Fb@HE)B,0PMFZ/D8N<KEXW<2+2Y1>L9
?9H]FcgH2E6R+T=--G:TKSg71g4ZU?1=WN\Y-/&bC4A=^:QaEUdedBQGcB0I^<6[
[-?>c08/S5KaF7?/JRG22_)#d8B0E[1>Sb,,d5W-G/FEX2LFRKIZVD&.^O@=.:7#
)X:6L:N6WCQ,)VFg.8I69b9QJ^_e<)Q/f?U<WL-(A;J0TdfD5VP#Wf)S#b[::GM=
aB.ZL@M>cNg+-PgNg/SW)GKHUV-=J^,;&806\V3)+-eFH6,.dP\O+3?-F81]BRGR
b81af3ce;[Bea(.e6W(]<O]L]K5?UPLMGW]c8]5g@d/2@EESNH)YQF+^Ng30]:<,
)HNF3\bd#W+RX1/_S.?/D7A/IKN6IEOg5KO/H@,c381\N&8RTB<]L,W0YM,g6K5-
H2c@.RCL(.KHC,]WIee_;62?3@ATcJ3dZ=ACMKSUg?.Q3<84Q#,2\C>?4,WH>;]M
W7T]C/&P=E/@2]L=)V-M<.a.#6OAJa0+>K56I)1<X;5O5NYPI.MQ]RA>(D19^7X\
EBcZ?fGa@DU;W_HY=P>2^7B[#FNU:Zf2bIRT##:CZa(\P@_8_S=I4_Y17&HT80<4
RF2526BSYL99&Z7NC;cI/QW6Q2JO9SVe,1&\8W>TLLTXc6N@8LN=EX+L@6_Dd&((
:F^a\/EJ3H[^+/>XKA>7,&1Ge[PJDDX2V2QXa^;GHA6.(H?>998T<[\c6@;Ua_.W
?RQS[ff6&FL40#4K6]abC]:-)V/fK^ISe=H.M:(H[3>M0#\3@f/:QW>?>2Q[Wc7Q
A]2,?C@g0O=7XLRfM>_.Y5K&P;^8KE>LM5WE\)d:@?]F-Y/@#_c<IX=_P[OB027]
]gB>O-7_C9Q0T8Xda0S4_?e>b>Z:-aIaK=6?0[L8U5<M)C/Ig)R#:9UNY50B#4g2
U^f=T/0HR7B<.+.7e^,g>)B\bNf11OH]C,@[)Q([M-6D\CW7g[YYK7O>NQY:(MFS
/CH9T9TAR0;KgRO3<g+R+X]b2g7dE.,1E?TB,MTOJ@I+^eT264Q6:BUR)Z&CN7_W
#FCCQOEdC#FHH<9BU/WXCgY:-&_4&E461/9KVJF=9RaZ\XGH>:gK<DE/dU_JAZMZ
O/Tf@F]a3O0(dc@d1O-Z9IKDcLeW>Z(6-cN6T,-A?7366G8gU=05W_C-ISe3AFde
f-eI/;5A15fQ5:D@#EM[I92GUZZ?6?9AX2g-[aT3\bON375.d6N#_^C8JTVCY@;1
8?aQg@NC#cE@UfJ48,WF2S>JUV>#NSc&&c16)g;6QUK4@cRG-,90@5dPT+\(REOg
cf#GKX]H(Y+_(JaJTK[@A_BC,IS&6&4KPA5<;I12_A6,&\S:ReV5<B3RX(G[1.I_
+,C/e1?#.MQ+,4_5/e<VK=4<N\7;eMW#gRF]Z_L2;G^/1])&-R_A5VX)B[GcS)g:
.\DH<+[BP)O4(9]0@2WU1[fD):AP^d0^66,D]-,G82-e4@CC.@[Q8G]6@Q666gg=
Wdf]-EE>AIJ7)0XaY)1S#<g6HM/_/3g#Y.PE+]a@=f0RJKdfY(Yb.+369UNG2XO^
LIHKFEZc4QZ-[c0)]11\CA&17#ALcN,+.<dFa<0_acAX&_YS,/8M1dg/(&CX#Q93
.gPNg4(N7_8<JeC1A)VAA=[VD@9?H5NHVW[gQCG^G_4d<8NJL16/HH7]gA/eGb1(
0GR0B)I.P=L)#2bHCgC)8)gFBf787H8&RA5E.FKPQG&B\OHf78U[UN+.?E<cKM[e
7Q,_Qe<]fHIM:L4>SQ:[W[1_L5E[_Bc,3V/c0IfF82c1[Tad-I;.bTI.(eP,S&J:
a/1TfF_OHc4fLY3M_ZS=)7FO:7K\\&X(Q<K-5^RZ-fFCQ:eAV;R3KYJ]YX4N2.:L
=+Y\Z+aB>aR[VK+DIQfONGBPNULgV,E7,bZ\R&H0D1#H>0<X>C#VY:8&[BE9-:F4
e=1W7&2JgWHb4=;AJ27e[[/_YA,^;2_EJB)Aa(1@4OX]=NPeY:7HV:4I@?C1,X9I
1JfD6XF1BfJYKEWMXd7Ec>V&9FX1A\42M#7Q38&K#[TU+[R],-BU\=3RKBK/NK]\
@QRA->Z9O+DAKPeIAU6e_7X4M=N>LD?+Q5W];XU9A3:F50XVI?BC,(3&OOW;PY[e
^]-c-[[&3>1M2AMS_43I;eIU(N>gYKfaYNO#(I7L9eQ5-]/;cOD?XCEU?S3^YODT
gK^W1TG/8H@O5F(^bY.G6Mbe2=0a(T-J+0_0FJa9)W^:8F179JHUg/0Od&U(FIf-
g\5a9_ARbT6-G(#a(SF1fB.ZR/e>785-PYE9>U.JWT@&_96T;+.CDZD.[148,@6:
O4FZ@fRRSUVdg0bSgeYeeBQIa@7[HU,Y[XfgKba.:)f]+O-69D-]b1Qe+M3&ULHd
=F6IX2Y8D/H]+KaGf+gYA8c33COIHMA8H)-:.I[RYZ5bLO^L-L5ZFH;=e\,2AUJG
_ad[(cKgWTU8d>?@fHRC62,+\TPU=O=L@E6RA]>)8=;#22.S&EE8VWQdS<@#]f]2
eWTe^^_cO6dYd?1.>7+.30QYEF.IJAV1IeS_(<dR&KUN\R43+^2eTZ:82Z1fOUE/
#G7;@G6,WV/3#XWN(-2.W&dHZRWg;dF30Wf8<FZSOC,@?]3;VX9W+7P0G[.>UGPQ
C/=5cTVHeTN9N[K\#>/aG_.[>=43FN<F(d.SB+c2/AO^Y[O>6G4Fa]4LL2Y;DD:C
]af@&Fb4g0OH;IH[(8Ja^b-Y;&_Y^1)TQC;;Y/#F_1?a/[@_D[]baeG8KI;OSC#(
[D))M0PU?D;EI&RYLb4@AY#@.N&>C[QUGgKW9AL?GPQ3#DeDUHFO7Qd#UC^bT/4G
;#(&=F8)YUe@GeC,B1^&^2;KD\2L<&9Y&Y/YXJ_)@g4F&\E6ROXN9J7G8TEb]S&9
LdVf:,ePHD+_]3cL/695Ib>],<Xg_?G>/R8:Q[D4+H_Z&SUI<f<.-406a@X,A)f/
EZ/NP6.?KRS&^66?PES/.955MNa-dC?568e0Z>=;?MJXF+LI1&#TS,<:Wc:PSg5f
FRe8=GTN#4E=]f\=YE\1V1UHH3?S?a3Eg^@PNW/6b50ZEN]&b?8>SD1-TYGeeUQa
dV9WWAA-9fH_W]J)PcV\gJST?Q<Y-\MA2+L,>UfIfJQcOKQ3D#,@7/ecVGc1_(K#
g^FADY25bEC]E?.EB3d82#>@\6@(8cTQ9<#@9ea)OG4(ICKXb,_1:BCC#Tb7KHK7
TON(-^bO)+ceT3YH7\Lf//f3I=LXdHRKfRF_TQ&K=W[Ee?^=gf^#1OV]^?53IbI(
RRN6+;EN)Tf(5[Z:,XC]#&\cebF=XIX,<IcBY:PW&SSB=:YKGN9g6PWQTTI66_9J
\/80f[)EMb]^8/,3RbYc7T?=S^N?9e:1:?Ue]dWR^C,dE:Z<D/@UJPT/?PeEe=2&
)D0J?BL6ZQeIHBUfK_g-3;O2(#3]:fe\L+F=M]+4,U8AWFV\dG06P9cRGX,1Q>&1
[4<]0/J28VgKZI:.7;c7_IL@MYedHYY&(X=X,Y@@:I?ZbH&TH.2QdKB?ZM:6J=eX
WX]W-YGd2.UR+6,8YeDLD76NG:-D[7T5U@Y[;cP)AG41[cXc/AU4\PABLHA24=)S
[DFV#_6.2<<30dT_>dI1F@_V\C+3QMX:U[(YV;5-1:S&7>26Vb]&L.fJNLA3gNTd
?>eBQf5>c2O2G&e8EM.]J=]7L?>]O:#=acP/dM?+UT3e]@?;AA[9Q]YZ#G,]bJLe
\K81^0Ee9dSMFAR\BBLDcDPX3J#+??:bS@RBKTGHU5)213&8W]b1CN@TI>GR\RB,
51CXYUW<+;@^_6L@7&f1O#<2XTIF#FC->J,2AZ0S?./\;20>S+gf8G\SH.J2aQ4&
@A+/Q:?[2CJ<WTX<&H9e_abZ4^baB/Z3WefZ8f8^K@T;NULb/5,.G[KAM4&6/?KD
(W7N8SB&?(C)/WEIF<AS>G6K0O.X-G5Ld#+@g/#Yf\:e,EX>LeFPPD)MA]^)1F/B
P@].4FF05@Og_(G?P<]e5-#;(X>ZH_?5)(V,a+T@&2D:N(W^E<e+<[a@A?WGcD^2
Z+cI4[93:5b0cgHB3SIdDMK;N2=f>GUP8H9>B(e)JZ?#gN71-OVX6E>Mff=[NU2)
_dO_C0F&Q0MP0L?O5QH=TBEGPSD)2g:N.Q:@6@7P/_Q;9;70)B=T-,-[_[VXR1D5
BI>AOT0dBO15=9;&5OI(W7VF6@e/[Z&,eFO8/-CN>[#fI]a);H)OZd<>8W7U>;c2
0I/d^Q/A3eU:1+HR5V;7FSLV6]NZeODP0(WafQg&b#8N-b8Bf]+JUR5<&Z9,J4&A
96JH:f(Ng[,bS]4@&<Nc;T@K+Y4cS-YE0^_+Mf-T57QX&9>OF1WMQQ?fH=8P<9.;
XMMcLR[AP2^(QZGS[T4]L2^=X2b]R/5@UZ57T^CdZ42eTE;eU&]4S=^-YTGN)7g2
M>6J/F]3c3]O9..U(;L:-X);<,D,2[],#BB(;gVdbBdL.Cf7Y6gJR,P6?[;DIY<L
X-)QE3fN:8-H^9@@D&2f]Q7XEH6U1^R?VQAPQU3]H??L1bf=PY?PBV;MRC5WeFK:
>,11+B8.QZ69fVCd9Igd+S\PF:D1fV^.8+@9LW53+-N#J<[:4)7@7C[G\g83AON-
BPfS^7LS\c21FMTU-gJ8c@N.VBIY@KPOXP22^TE\+603;:OVA2FI^[aJeC)L23]7
d3@RB?Gd0-=,1/^M_.@Y3(1U-DU,I^fC?/87;(1AVM]?N+6EV\XN/;R,R]7==Y(#
(/MS_=RQH6If/B0^CeK^@S+LLVO9A5eKG?_I9e5d;-&PKcJP)#Yb=E(+_Y0G.3^N
AScc&>0HZ\L0>9JHJaT2,YfbX^^b7/a+HQ(<JH]<OVF[=B[]Y&Lg,902>/W/G>Sg
.0G<g@:LOQQV<#B^fG?7K/M)e1#TIC,LdPY6MCD:ME=a,470[^c6Y><U8fM6/AIR
PcL).[&Z5[1EAIGX89G;cWTW0N===1UJ,G@]B]TT&^DcbQEAH6dSIG]K6=LYQg2J
(bG;[>KE:X#3FH7+=3.<C<Ic&eE6Cb07I<a,8FXIT0]ZR3+DR[N)P>:^7d,PX#(b
e80K5]eHI0&W/78.:Jc63/#-ZOZ33>6@(NO?9/H-A6<2cgFBS:N)cA9ASgS)AG,P
N,DYHe,QX3.7V\dKFN?E/AD<5BHL<<)?XH16,]S75#(C5Zb,@2,-.bJ]eM_EY:70
?&L1L+YYT59Z9?X+\SR\2Y?f(1KcC7B;ZS#2\;ObI@[HI3E0#&,D(AV</EL99+#R
H?+4SVS?G9/:YV^<B72R<8HM<0;MFG;GQ/ST\UfY9aY>KBf@aMad@La05CDaZcW_
)I[>aP,^F_ZKG74YOE.H7JQ)fBSYAL)B7^>9]778AXT](+-IO+9f4-S<3VIg6Y/5
V@F4;cg4LWY.M7)dTcX]6ANDf?B^9b)b1WX.+c3dIB;T=>4DWM<3>700L_c/41C?
=JP7Afg:SW[)QC@0\?OOK0)\-WbY:G8FV881dKG05B7QV>?K]L8<28U4J((4a-_1
37^EDe\4G4?LBMQ\P6e-M>KG/[W@+TP[U(8aJggS9RfJ:#W[ZYSEc1.H^XW,#,fN
.cD>BIAE1.(^<W?=8W=.NY6_4deMdgSQ1C)Wd<T^K8^\^Jd\K)S:RTVG.0?Lc.4(
RCUg=@S)EdN]+,f>d^R)^TRPa6+[4YL#&6XA4+AQ.O@ST3eL637K9GNSLV\,R(\Y
=OP5c^_F7[BE6V,3A&AMSW#2JA96W3SLR.#,eeQS5)e<8Y(\I)9dc]b/LDRZ)^J9
e[[JACUB873UBU>H^cdLM7d&OM>be.<8Z7,gPB:#-cRGb9(Bf6DXC]AW+UL4MT;7
O-A-9;;ZIE)c-&bR#1b+OV>JJcYe],8N95WMVLTG9MfeQ(E/:(P(G/^04[-\=B=f
80U0RQa2K&2^6RXFT</_,.&7E3Y69eAa+AUMaRS@](-9REVJ\c?268_4J(_>8D#J
>XNPJXE6A^<I8/<Z6UD?-O</QR:P^46fN[L8KN@][XTceeT.(@C(Q)/_6(Y)+,MZ
eTe#)E;^BE3:W1QD<\E>+](W@?@3EI]SFU+_[_\^f+:]GgU<&cO2<0SPL8G:1:9;
8b\#\Nf>a?\3b-#[;GE[aMS+L8I)PPKDKUTOU]];T=I=E+5=@bZ6KGWJ7f4Dc4;^
LR9BM&([XM&4>+H#J+8AA;?Z=GUb2M[6N,L](C\=^ad)ROYI5b)Y6.XbF=V#2HYY
DG;9EVFRd-d(5QE+IcS]3(YQH;U)aM9AH=T=7\42(X0Z#:,9\[GO6-IS4A)B3E>#
,L]@MJ8IH4c@M)5)N7EUL42^594E,77X^NR542T;X(d(+CXfT/2+/8aX1H@ALBS#
M2C#fOZAJaS7[X<_gYQg&0W:-^H-02PQIO(N;P9RD7K;V.D7M0O]ObV#WJ/SB9MI
JScOD#PIBD44fbJb\8)AXaK&595EY9.G>f9_gS?<;VLBA1]RH+Ng3eV#:HTN4>X;
\G5SW2BEOF_4ND.3_:?HC&bbU&YMVMTJ7-bQE(8#Cb9N6c)EHRbGd,Q&Zb26E\2L
OL#=9=_]RaPI9LgKK+#Kc-XTaE-4:AM_&57>)VZ^=#_V4[L:IH>cI;IY;HQ;X?Cc
Y04H.Z,J<.^1ZMQP)3&WC)/];3YP-6RQ5=]e./BO&=:11I;EJRQ\U]86S3b+X6YK
aRO)e3PA4eSFc4,S0,^=O2]FM0P4:-PKN1Jd;+;8/O@ZgWS2S^\H<baA:50M:P<,
OAe.&&ZUA&PQ4,WL,?7FY>336X-5NK5e3&1,I6d8#V#VU3aM)R((7\6_@,_Te>Mc
Fe(5OV5Yd(4HZS>3S,ITZ]<)L&;bF>->[2cP79/;[4Xg(=><SX,YA@M,M<(fE[;W
/Y9AIEZY<W/NPNW2X9Z;MV=VTXfbTT+cc15Y8B1bAH[L1(BP^.Q\F:,&(c9(+H07
_ORQG+eBA8ZM82KY9cY1/7D[KJQ\cT@;<2\R[3_2V^.)Y<=QH4F]0[NUP,H7[a/e
[,^bL(Y^U(6b/e<ddGRE3^dd<b_4,OX4BAKSeHT<FDS5;UFbBN87Nf/=Q^M/:M;0
W\c-V+?@V@DTe<:@D-C26[]EV=OYCK3NWQY?TN\&:L.B&^4LIe11EAD8S;U2?5LG
08OZgT2#?a&O/EfTc9.K(.SPFHFOBB0/O0:7V6&C1-;AR[>J5@;9eZ]MSe3MD-_3
Sa@B<@Q/J40gW&-a:=dTf1>a>F+9ZPGaG(@C@g[:ZMD>EKdf,=Q:K<W1Q0VHbH.X
G+T\@Sa\+A>?RNHB:Y0<FdC[SSQI\aNXQeY[Ge<8X\<+GQ=6U,ASO)adMQWOHf,Q
XIdC7SIeDdX=9P;9eeHd3X?@0[RcP:cI+d&^4<3:RKD/:H4\202>I13Z:9WScggB
07<;<W;MDWEZ=K@R#f4FL.E85=+ZQ>7+6c6JAM7WFV9PCW^,+Y@d+,BA8^F3=B:J
0DMOG(T_\-+<3d]3O&5/)a]/a.BXZC<KFgS?g]5P>9(?gE\e6..D1(KXA6gV^?LT
.NB-S_dNR>SPS)([K7=/63g1OeUIBAPX+.[2:JZ/a\[XPFCBT^1P5Xc;Sda0ZNc\
9P=ZS6UL,0-#+(W(L:0Z-0X.,Ed4.]VKH57+J2_DFO;]N[4K)?C#fGB4cE92d]b/
4e<:ROC:4^KITH+f7MBaS(UC0dMa#I3J>P>=g]M7DP(?#;L(SfLMVcMe]89R9agB
DfH5dQS;2P:f=dH&>M5L,]Q&X#Ad-Re?PF47SP8^X>/L^f1PPEB@gNefR+?_b7be
E=6-X(&Ue287/:=6?Z-\-SbcC5\RJT]61L45MH-IR1JgX/<A6dda:P^ZT8/D81SA
H^M.d?,+K4@BHJB\2a\E(XdAL0<b2/?^aH5>87IVXaVTgY=b^5>g6QBO&G->;B8P
TI7O+IV(Fe>X/L?<2ZI3([[I(L\)aO4b@M3<9U7[R-V(YO^d\a\TZ@Ucd?3A:eg,
E06e2:95]>(9TR@aLE/<VZ#R?<QTfU8<Ged<5;>^UV#cg7<D5ZZEFTJX\=TG;?#G
Q8QC))AI.CbL1LL,d>M&FO>/TQV.[.4H]d4BQd)Y\AQ1FHg,V:8V#5TEP?L4FE<d
cA=L@]AU@)S9+N&#-H&OSX.HE,Q6CE2]&LL1T_YcHQ.M1f#NZeB[T6:gBZD9c<O.
JPFAQXVR0\S/Y.I\,LB//6.TU<5AGT,@eS:##QVZ#0PSE?3X7UOF]FD[6TXdD.CG
b?>ac02#.2V82>VTVb#E?FV/@2\BZ9=9PIZL8DfcZ^;/85B</M^)[LWJaDN4eZSX
ecIK[Q&MH/Z0Z3Kfc5M,Mfb\@LH>.+a<9CRRa3?[<<.B7K2)K@M_.,.&1E:T;gF\
4[\=P:,Ag9@65>L1f<b3;R9[MWVJO7]@GMggBV\P36PM:8NP95MU2^6gFbR.3d3d
NB\eS[84U\V)^FM(T@L[O8VgF(BBf(/3\/HYb3K6E&SgCGTCJ7aKY1(-/@JQX;EY
<V;@P07O0e[<W#\V>Xd)-?RT4Z2FU=cCb.9O6L;IX4dg6gMaJ<XeLA+K;CA.P.dW
,8eSfH2PLA&(M<2(]T\BeA4b,D+c+HXTFKdY_&fc.0V([D7DFLaR<&Z07Q+>@0AB
6J@_#I2#5;&Fe.1>.>_,XJ2If=64+cMAS2BB\A?T+cN?8EDF22^[MFG9&LMYXUa>
[?a5Q:&,-=dc^]3]/dA=C:dT+gLNS[T:+HKEZJ>)?FYB-L.b:PMJN3/>8-ETYTaE
9E_=5g)aKBP+)69^3Z,OCgR&\T:>:^KWD+7YcI6#+D8A7U^DD#YJSPQVYe^?XJFW
)B6-&LNX-W@UBcG+-R;3TL(SDNUK.UU@F]d=TTX:\]S+U(&-Q:]cYF/;Cg2,5GcE
.85Ta.c;6dUKPI[:,3_X^c9NJK5X8Yc+YKZ?d<X4)A2EM>H7a61-K&78Yfc3DK@+
W\S0HY@:3P\(UeJc\_+2-R_Y4==@NfJ6:+dQKQZ9)T_c<Z9+VJ8O_^8<fP)C;g(A
J[;R+F=Z#.,#>>0a=5DB9O=]CA[aL,H8UO^^B8PJ:\PAeg?FGIBF3FB3G:0T@4ME
8Nbf<:U_#B<R-9C^.:U.-+#&UQV=CY/30<g_W<KL9(@73?[GPM?Q<VGW(fa0&6De
3LJg26/<],T403EWV+F-cKOWDWEI.J[-W0V:[U.5@,[^<F(=H[KMK(PVObFg>;\[
/E?.98/?b\)a?/aaf(=),FR=gE@I\_\=-OLZ8_ZD4PV4fM2/CMP/#eM9;2_\+R_a
Ad\\,_MbXGUIGIU2MINSX_MEdBS/H:DA/5CfEW:Eg&aSJ?KdZf>.8ZQSdPcR0D+Z
OY]C<=XY04,.1++PZQ/eA8\29D]:_KM-5+UfRE-6A8]edK@)T6@?d7_KSHC6W?1D
XZgIeBKI@QX[D#+-=[X4[F,VEcb8Ea=?1YPUdA#N9aL;>Z9QX6//?<-1[CT1:.cb
]31\+9P\>FNF/U&gbH6eU_8.9)O>D.(3W@@V_0D#+GUZg/5;1>EEB9C4DI2VCK.(
(X&75XcS(M;^BBW;HWZAO6\4P[C#^E@BeGANK,dYZ[b=13S_:=)H04^TER1/4GX?
=;9NDZ#2M;&Yc]6KY:.,0YS8QCU&<#+;X?:8.RRMT;M>;eM&M/E4Q_&A9IfVV77(
8[W:SU4DT\O,VHC&dEHP/9>XL4:VW),^KG8QAd8.L&28N#?-;[2R7STB085CKF6J
]U&^4P0:&MWfed=P\DU+N\KAX5TgNb2cFB0g=>/5F-17RCLRX,8;5[T<?+8)JN;<
DQIT\O]DHOCAXMXP5d=^9MN\d(++P&3dLQT29>;cMHa@+S[4X^/#>aO+Y1QA=e_S
c<#1\.UFVN],45WGIAe=c2#6SQ@BSG\]BR5g]^Lg@-QaJd__[4#Y_A_L2WbR=C+g
f4DK[<2(&)[T44\4RQQ:3CcJ:6)1/Wd9F+E)f.7@Ueg8VX,DPZ[9;eS1acgbg(_J
TLCZ4)gENc57IJ</X<S\Ncd4_fPUC6:1P2c(HZS8(C)LgG5f5Z\OE?2R>Zd]Og\O
)7a_N=69=@#?3[f00Qc+@ECWN,N?KX)>D#Q&S7R3?X.?eFbf8E6KFA8)OWMMcF7#
bE6dFLNX1\:0e68L?Mb^fgI(GZZQK5ZYYHc0EfUD\U@MCGM@5&[&Z\\<ZK0&VB7G
J22Y=1?WZgd-dNT=/J_GI:f\4WX-2ca2@=>.dZ-4?R>,EEGHNP/9F)-);9EX->12
P=,7HJ).#b;F,S;\>Rb.1(RXRNU8-[FX^Gg8&CB/3]a+J3+P>K9\4@QT7+0Q0<J8
a/409G5GcKD6dK(BSM/Y\c^OV/E0=NME2J)G(7CdKK86MS\XbJNY(@?F;R7IKIdY
40=M]NL1a^4#g]WYgX/dWfM=F>0dH=b,_M#:N#)\E;-U#GV<8eM6YJgJN>IZ]83D
89/?dN_eD79MEP2B)5(MZ+9.1^;9,gUF?f.E6\A<I><LaUN8A3N\f7faeG-+X0J:
fbF2\ZD6WT_[4d>O^gQgI.d+>L,_]XX5V6Jee,)Rg57:ed-JZTN0:+MB)78S;e<N
]P?84XZ[bYB&&BPZCTQ(5C\8_[O1/0ZG]ZCUY:SA(ecER92fYV]\X3)W,FJ@K3aF
S-Y:51=Z?<SM:SHad564?XY4U<Pe.DLQA=X]HBBO5AO[HB:Xc;UX3RN@4FI(-H]g
()UcaG9:^1=6C;RN[?Va;CI52d[KK5d;U4YZEMK^>+dTPc)I;K_cV+(eTR^U:CPc
A1X?P61>0P_YS1^Q>B&a9b]FGO_cd[[>\HL?&/KZYTWZ[@-8AK[E>];e4#,QGN6+
Y]G)L:H-G7d/MZ@dL.566JT63H#aY)ZWP@/0J4WD1SCNKI:)XcZKHN\f7;cPHPCf
-BK<.UR:\&@4LbWN1;=XW(<((UX-f2D?3HFE[.<#C1Ed@02#RF72X_A;BB)2P/E4
e[GA<#<+CQ3#7^4_(]ZEg;<W-I@\8g7P7(J;-RWNC4-QKN;Wf1.G&OKFC&GUd=F#
-:5-9dRL/Z^>EKS0YcZ3;>9RSTgOE<ML^.QOY(;E7DGV#TBSPbL4IKPXOXDX0TC6
)+KUgFLb+]VA^g34=5\6_Q-4WT/QUX7acf4,8X=F9R=R\_.CSY5gI04?GI3(ECS.
(H#)1+e/Y3a)R/6TMHd(W[\(3]-P#K:YTLHQ#E6b#Rf<B8F7??\_6>LMP+=cS.ZP
VgaOH1UY4OFb@aW3#EEU8Z]/c/W/UT)/?&YR8>&1?T:PGA1MZ19&<IZO[D?GCXa<
BTYU#J+:d2(UR_3]@?S^J6&VQ9?.Z-AV2eTedc)LgMWa+<^BQ2.QaPZ^37T8<O@7
K:5-[X9;&D(QOCC=NebUT9RND.YVNDS=7f@IXDdCb5ZL20MQ_EMY>Fe#9Z+X?(/P
a1\ZIT-&@\G?AIPN3&1=8#3\DU9&?8OY6Ze2eHFI4EO9.)9eL?FaVb8(M_F+/+-0
Y2IK:ag@:R#Q?MAW]7MXJDR>E2:_>X#0/FNP+AD_S:]8_E8Z36IZ2D<7b/,^0?PH
8CH:QK),YT>?;<gM#dG(/fQKW&H0H;(S:8EP(aUP\1Y9g=GTdgS@#dRKb=[KUS74
#D?@TQ]C8/Xb<V8;QT<L^ICB5_12ebQ81dRa,UN9TaD7-K#EWG.e;-XEF>cSf/33
2e8[:.Va[4BY,+FT;S)>bPL2W]g#Fb=[QO,5_DJ0)A3K1G_51)G@[K:I.^+<)Jgc
EAN7PW7_ZEESF&IPXS?cdN=S5L]6O6eAeJW82CVGc.9V,>c5+?LO+,[0Z?[>22B^
\I[LO-H=QM3bY&P:P3CM@DFQICQ[aUFA=8@+4YdO:81ZV<L1]=WTDJ^Db2BO<LIV
7?g<\]KQa1MXVHY1Q:Aa=3C73YJ-9RX;4NT::LXXL1A13L+gfG[<HB1MCbXgeF@>
,H6P&Z^EddYW&FVOg3-fD8BcLH(N:XQJcI?U+-A0fPeO9\WE])5f9FEXL0IGI<f8
0Xa/eKRc9A,>8-1M_5X9DEgV(9D:3Z#2Id7=&A>P9\bP4OKS;8L^?G;8NHfB99J0
)aETb01W-=+L73(eQSEb)ACcX)9IRcUA,A#CJ<ad[C>&-S41@D+dC=>7_][_bLa,
9_fX@BT+TSeb#;[K&OfS(@;23C_C73eEQ_eK,+Rf:?F^3I+a11MW4OSPZeTB(W68
,>AW:4&:>bRX>^:gW=QH]04U?#K2e50GI^.&&^J,RJ5Jf]Va+):VH5cH:9;H_Xg0
U<Q5J&;^?=P>T@]YK9^)02R03JS=O&b[Q8Wd947FUZNR=:+>HBJR,JVGU-QXg384
]BcW9df+CXgLK@(B?3(a@_f1MD\3G7R5SBK\F&PX<fAe]W\_QIb#2@GcS-2^B/d.
6K>=cBB,2GWfY-SX]_O-(Z,S6;bE],&#gdb&.EATN4NfS[,;b:FP26:I&GV:]Xg-
0ZT&R?=2c)3IYEOIN&g3^BP]1AG=FZ^O\SMNg=(?Kg-S?<;TA@>>]OIL5/F=4e[(
eHOUK8+;5C+H0IN/<=T/ZA>Q/X]&3I+,G#V^I[_F<Z;HbAce_fZW&(6#LSU,<J.]
OEYLg7-C]83D,T^9MgZO(bPXIJa9JUc5):ZL6+TG[Y5PA&U-778-]8=---P-4I97
H_I>VGcVC\5f]8V#6f1H0Q3:EANG,\EK:ZE93#G;CG22^(<81@^O\DV=eDI=+dB5
DZ2(4LMXa?#cA^]c58MTH3)^J[/LGF)0-C-&Bc,[N;P+;[<<S-e#\fc5R]=BH_B@
XTA7-BRL]fOIg(N+E[[JDbb0DEV8.V>&Z@K49K[-^@@6,4.gL#WWd30D<=HPLY=S
9TbOdFXVGVb;E6bZL:_GbKfOVM^(cUbO))SY3DO#7UDG_D,a:#IYOITE>eE;V]7e
EYFSK_(\NCEI5ZeC7IXHf5OND+1_bHXHX#/dYge+Q+,T=\J>](9?VX)G0d)g1E(\
FeHRJ,,EXH_W510.aG+Y#YYS=Rb[02(KFJ683=7HY?@H(/-(L39QbT-AggCW;,AV
J&S5eb-H^3-T66&g9(7T#gIIQ>e)BT2A+\V;&D?R79;cRFPA;3#19?JR;eV.SSHC
P,6fJV]acEZ<W=+@3d.@912Q3JZEKaVJVJ5C7OBFU(+.Cc/3.<JY5K[<V0^X2g)g
aEXcA):1(M?1b5>c=>#=H>\45B2O\0;U^PBGWHJ.a@CL&UCI8KH^XecQ^9R?61J?
gV/dK=FV2-;B#ZCE7W..-4@([[=Lgf6/N#/66f9OQJd<<5VK;H\15bJM^:1bB&Q<
//XEb@P?WA)I8D\/K[)T:TWDf.4gV0M0IBZ22L=gW6cV\8OO_b;PO4)P<D6/4?R@
_CF75<GV.eP=4N3I#a@U?aID2<ADf4=[M=gS6Q,SR^O=T0H22;<9.]0BJVabXUX\
1L^=[I18?d(FWH6aPAJ.ZW(0IBAQOcZf_6JL+FQ)5@SA17ODM[\ANa(S[F.-Re.b
E64T^J(f;R(X_+g1(8.1WFHfYg<6>H\DUALdE_QIX84&WMV,.(.=]3#bS@0FM[-7
fB+TWfAQMeWK.Q2>_VeA-dK#CK3760B2I[b5\/(dFRIX;U]11_]ag9c@bIK)TSO:
Fd,D,?,b_HcV=ZEKg^<FP.(-d9[4AZY0&JQH7X\P\6a.H]-&URC<#e>,/K74U+VE
CJD8:3PX)>8Bf;O3gVg\5+-Z@U/77I4:DA36_Z+7RJL=1S7UbXY50b4e35WR\#.F
\>LJ<DV^YedEZQf+NH^AJ2cOLD03-1-<)/=<QRQAD&HT3QTJ)G?:agJCaeBaKLC=
5#cD5#9N_3OFYCNT54,#R>QD?VTM<4ZT\0];SW6?]J.?g>X)78@?4<\+>0&R1&MU
G#9&aU,+2A4L#Ed4F&<.d0WIfHMQ7@R_3:&NMcL)]fbS(1R@>c5S85+]\YTU.6PD
S:82XR<a^6;-?+N_NbL2]B[Q-C;aS&N9?X;a<M2Q0\^4B:dR[(33H-ESf8XLJN4+
7g6D/+:^Mc_Id&C22=PN-c-a3&a@#PC.8IQ@AaT48QP9?_JV-?:=-S@)AZ?eg:-4
Wf+MC(H@1(VPY&fB@\)J4Q>-[1^b9g\X2&cADO]gZZ^S+0fTdO/,()GYR_B466NS
6[)=0GKCKgf-(V>3S.]D=X3-d1.YQY+QKA[dG-A)e]0N4Q7XJ<H#Ag9b3?U8T4F0
Z#4_5UNI@E=2Pe&62d;D5A)>R)egHc=eZD+,b\f2<1JO=ge&_Z9:egC.e1UeT+Y2
T@YJGR<K:/[@46S2]7L5[T00,ZS><XU[Y/T5.W/P6+)SU)LXDXVa7H>N&;,@VYPZ
D0B,U8-&XS0bc0K=A:6[MKf_fGARa+:fc1Q2Q/@G0&L/H#5c(ANeG<UN4C><WP?A
+;E_VL-EJXE3ZF0:Q#>I0-e4ZMX_+,CUR15d^V<0BTOdHXY/eQHZ57XAB5NC:;FH
Rc9\^6&C=O=dHV.#:C]8XcA\Z<.CIR>9?:#LN6/(f+L)E+LY3/TV]^(Ec&OVJRE-
8QIH.@WOV>@[?4b?dVXQfMR,)Pc\IM-M0:\NZ1)<[0>^WG1Ac2B8>_,HJ)^c#1I)
#D@BX.NZJT0,ZE]c[3O44LeD]H2W,_>4X,.ZRD_OO5@UG/d9RL]7Z,4I.3gHCZS@
HB&N8RL076Gb=dgT[M/DTCVaK9WbaQY^FWg0&@0DMeJIJ@V;FJ#\\0K8:[B)X?#]
GM;X.B#ed5Uaa^437Q[ZO4O#O7:FJH4H=gb0#bD,@(=/C\>Bg(QA><Z8Z)aQ\9c<
ZeF;@1J]6b&9N>T1bEbG&)BC<E?(ISaO(VcgR4f732fG]Y>@_g.>^)QFA]ZQ^FX-
YU9P&LAM9ecF20L(#Q3Q16D6JKP=0[ZZ:YBfC0,(#Z8=8ULG;I8X&c2HDf:9,+XB
<V7#f)>),D,DF^Y]G#F&1F.)#F#@32^K:[YgX&-44SfGRBOA310[-T)bP#04Vfa-
a0d]9g>#42:,M+G&F.CdV[UJeR\/4&G;\>Z]5^GHP1e05&-V?PM-.-;?c6,)2&#>
X;H8MJX/^N>HZXY#S;W].NE@;[JDDY_&[L.FY?_]]80cA^P+6WFc6^d3:G2DQJAb
<P(c)1A.,J>\KH:d9QFS:L>\./8PVGX?HfagJHJ9gRg85:@IV),).#CbKa+9B<Og
0Za#<WFP/BTJ@VD\K7&_J-?Ub69?^>#>5:19HJ_N.<\?&R)):Z)S.QP#EZWFFK;5
#G7&]R/;AHY_#C#>.=5P0@<4>6X7ARbXee>NU7,#HZR)g8IN+e=B?f1aVW,c+MFH
Ta?)AL98Mf[5TWWHU]INNb;P7ZU_H5<R,OPRb+gMJ:cHKEX++cBA;YSUZTM;fK50
_J7CYZQ-I-^8.D;[D]>FA-7>046_\^B[([_KXW1PRUZc;C&IA48UG(8dXX?CJMY;
LV&)8b\HWU48c3MKUW.N=JX4eU7>]IFOVb<VE7KgBB:SU@c)7-D4Pc@GWXWR2=<Y
)8C0<EI(geT&GEV<=X30;Cd7]=3\[-T42\<X20b8A1:RZfJ/U?QWd._)(a/+=A0N
UPR8#YWF/>TfSGgB_XW):cP,gL4)c<4&SO;E-IRcG@1>a[g>@P/VE-=/Z-/B=7cM
1UCY.?Hg+20/UA^_2RW[=0@FI0N[E@/Y4WQJ2@aC1HW;bX[)QX2ae:5230M??5/W
O2&)OHGC_Se@#Q3.C=X/d;9AZ9X@@51F03+SJ/&;VA(;W(BH2-1M6a[GCfd#A:YK
cV1g+5ASUHG(JD/=67c3Fae\+,-40af;9=7QB;QFd-PLK>G4TSff4D<?cM>fd(c/
5+C/3)eK2d_>#JPKF-f-g0GFgRC<=O9O7=?2)K2QNEY&)aeL(G6bXCGbZg&SVfHR
c,.?X[ETMZ-7]L\I0>(;?U8#]f;6B.9B62W;aY\HGA&@J4+cVKF;;G,ID05OQRST
5O,<;\bgU&bHbG6=HW9H_NB)Z70XScL7I-6\ONdX-aNEM_D3R.J#)8-g;T/],CGc
-^eGQA-J-+:TFJHC/P4UTYX4dRWP.CM_7Fc2^>;FM>;d<[09Z:RNQdMeQ]OH,_62
4Kf@-3XU[P@,I2H&^&Pc:Z;F2NH+=7&_OWE#JeKdM-YK_=DdC3A,Y=KS\]0CbXX9
bc26g[a75F85Y283KYV]1cF8O>aJ[.@eH#/5/,T@_SLNS8<ECHbZLFLRK@#@GQ#G
a7U>NV9g\NdN:ab2e@&geZFWJ:VE_DK7N-)QJWPe(D6IZS1gd6S?T5Wa51+23U^7
;H-fP3+:&NY.;60aUW]a65YYQJ1JA:eLY8=J#MPT<dWQ2GK=N(]e-,+\]][,-;U_
b<@fI^5\.7gG>@,;gW=6AHP/PceW2M=9>-_TXL#UQX(GU00eL6=2#1S^)76=F65)
R(&e@UW76A[1Z=/YdZX,S,UOIH0dPE2_IC=H&Ed=bW#9_[F,c1-Rb428M5T+:2dH
4Z?M1AO9ND]@>(XF+e]0X.R=O?1QFT]:&Rf?KQ<b8]b/.E:W-YI3R6Dea_<N43+W
4]F/4g:Ic?)@O8@W6DE,_:37SA.NVMI-:3>+3Sb=X\K#(L<U.<.\854DY^&?7?_(
aA8Q]LX5:8+HSF4C0_ScOL2U7?DXUSCFa8T]_ARaZ+eJdUH@)7<8&T(P@[;92P#9
J.IDA-/W>b=e68KF;d0:g]:]2:d60>I.Y3_W7B_N+\=S]#;G-FeQ:TB;)e=R>d8-
YP>:04;Tb\5TC-]aX]J2g:9aa.KB9.+@+NQY;88bE0eM>_N/^80\SQ5S#f,?H>VG
27a0R=QFX_HdbB32NL)0,-Vc6UP?KKZD<eI82?P9(NfeLP:fNS[LMK^<<JVE(YG5
B:1U?P.V3bD)N+1f0]eEYP1ZBdWC+AGO/;T&?(ga;LbE;]0G4R1^&4/_]01M&R[3
.HP+X[P_Z_eN4@DOI](REM=/UTS[7U.[\Mc0\IE-^V/GHWbeUa7VJ@:U?&.M]bHQ
=I]^-^5->M,8)&DFfb5:Z+L6EKK/f&\afH][-Jg(Z.O:+SacE3BY4ff=7V6SG(Na
:/SJb0-=YW2:R2D+JEOO)MHU=efJC^85/]d^:>MCdE;#@58I>01YH?;,&-EF]CUc
R8NZDMD<,M5D=9H#OgLAMEU+JNZNTSRNUY#dCf+T#d:&ddP/[0CCY9IY7S79?c5^
=.IOP_Agc+M;UO81EFd&DeNe7;F0aRX)KTHbKZEaT42H:RTT-;TA]YDRb@RD81Y)
B1,/<NDO@?F;>0fN.FJAT1C5aBN[ZXA-4-8J.]d.:X0BGPY#,S7JDd:;-@P\CCUL
:M,-c\#]#:ECeH,f4?5N#<b2IU+f+V)M(7-5)7V1?&](H1G-De=eT:C3ObHGV;L7
D#B5TCU&,f5g\;RWVE9VOSc1\W[6XM[3eO>XJIY@)#U#Q<IC<WKAX#^1TBR3B+GF
24Nf1D18/eSSW+ON.)?-3;6)IDPWJ-1GSO>d#<AQ/5WOcDg80(2dPeP:FeTe-T^T
Ff.]K9L+<Dg=OMK]6g6eZQL1DZCK,UdPK0Ac\E2Cg;LU(>C7SBO_,=(E4],\1\@Q
/9DQb],G+W]XX6-CQ<2]^IEZIVUE14I]bE=H;.6.OCFRL;a,I)_E5YOQReb8J6]N
gTGc811VNX=e(B^R/,gKB+LBC2N12H_,CGAbO1=;VOO<c[BL>.07=1ZH(.#g#?N.
g/KO3+a5BJ-L2BF7?&OdGC@.Qf+PaSHDea5AWcN4-U9-3TC807:N^/W-+C0.KO(J
&5?_7bEJd[^AK?.J2<)SM=AWN.<Ua_\?P-CaM&UG?(#:15OY9PfZeEGBPA)5>X83
X)FWPMJ:25Z5<W#+LbY.0]2GW>F=VQN:gbARdDFFZQ#_LGE,d&)<L>>[^C[=L,,6
+6,/^>Ga)I5]M6T_\C#O7XYQPAfA71HfAd(5R=6T<U:Q-QRZ1[MVadD(2<E8YQ^U
2J[a6P87UM;:O2\TVD.?TQ+ZW,@KQ4A([-5:S>YCZ,/@ba6;M>WQG3L>4333SZ26
GH+7RECG5SI3FHQ:D^UE5a;&#MSH]4SV2MM1=f)O>1NggNAKTT@f4M<gE,g&FaL5
ZYGX-_98<SK,I\K6JcH?5?)_]bB)8G;&QQd?_U+;0@R&f&^NHMYM+V;=#C;ZJ?VB
#gacb\S=:6eIN/KgWHBg-<3[_>[4e.eX]9.b@4b&[F\aLTcKLb:FV[OV+XaaTB1=
6O0[b6Eb_LP#]&UGN(M2..QBS6PfO#UeZ&IH&Oa\)8ZIV<^2eLE)K-=MVM:S5?RT
ZVeCJgV_H(Qb8b^9J&KabC\71K0BA4A#gLFSEZP(GaOaXJF\[10ME^a@+,TV+,U@
PEFU/FR=7MI/0^4/g&dIcG@3W]PD^_RbT9=0M[,;;R[T7_4:]@#R)LYRHDY)9P(L
(b>7)Q>\9(2]OJSa^GNESc(N7?UX]F8?I/:+HW4T#XKK/Y^E3X[+HWJP6;USEc[g
VJYUQ-KQ@3;,OeY?E(dIaUR_QLZU-4eRLY5U6P1):)1-.TU[2^X9[8SWDZMe-1MI
7.P^d2:DAL1/+#1A\\5:.@OP^:FEZ^[(&NB;?J(bC,8a?:bWYc2KG#6:&K/37#_[
UW6W>@G+#fLG@\LJ&WVc<(9IF[eRaY;MO],=bS^CbcK-ERQcS5f+A5YVCH>1?P&6
?L\fBP+(C,[\0f83;)Af-1C2JN]ZE>CN6ZC/9=4W4YTS&I10&8_+9<;G&?c+&U2e
&+;Y+BDJ-/XdE+NL=QYRRF-a>@SeT?\O&WK.e4#a/47;N6+7OD/]5\Ma=XPE3[O\
-S.9NGeJfV-3..#B6EM-SbOFS\/Y/+bdd<:I.G4D3Ne09.4X)=/>3a&3O613XK[K
C@[a-7H7LXT<\65AGYX1]KIT=:.^P/;I+b&)N]TE9dfWQ?)Od]dX(F#;+)^A/GSa
fWYZ:d5\3B6?COA5Q\3Q&Y<&&+B#Y6P/cO>4);::L3?Y,Nc(H^P119D:<HIb2QSL
3<1S\^HB7LcX0[94XTX[IK3T-B;E]()XKHM4QHJF\XX-39;f)ZC?#UO>a)UcC1-R
DR;^#MQ/Z]@V)0Z&f\(>R6VA.GGVSGSd1RdAbf53-[4\6GU^;4&WBdD;:d7GBU1c
W/TMdH/#^_J./cg3eJc;gU?C(MaQ/R98LUX/6b_Y>YLR]IU&F@)C(+QGL+.=f@J#
9-B_c=-3LZ86D(#Og,@QfJ-O9ESa)8_0:)dcb&?UG3?,TMg>=G@JN,6d=J)b/MIc
6BP=\@2P/dFB>AcMbIb?LETKE+0[ML26ZFMT9D)D1a;ZJH12ZCfK[\DHaBUGQf,T
VTb_[VeT2GW8Y2;LeVG]fO#Pf(Y5E,0VVV4Ve/3;VODFL]Zf4\d/Ue7]<=;6ZR6\
1?8^492[AB./(-Z.,J4QH[P?B[RSI\Z[&<?2XK<=IUXX,c?1/K12^^5/+#?@M;dE
+3M)G?K5G45XSc[;QNf,cZD3gIEb#b.DV3c3T9[\/>4+_-L;F=67KB;^,P^O)OE3
C&T4GJR9FR(/=]DJPL&O^<Nc8VR>Q>RXUG4=]1[3a/O&/CVSTOBO)BE)=KNQ.d+E
W[.MJG1Q3W)e+YBWeT4AA9dfVT@V+0@<Td3?e,]/9D0?A<gOZF-@VKVJa/M6CGL]
,^?eJ50P-c8[\JXCFZcCA3W^J16M(Aa]bZS4N.(;TCC9R40;<N;AP)RaY?g<9;/W
0:gGT8=@[>TcY;g:Z]20?47?:A=#5fI]?>ZGF;J:/@&&eU[f683M\W5QDOL<T(#A
FGTQ;/Tf.N3FZ^:HCDPH.F:Mg^.2;)IT(LK_,<0I>8I\GX2@2bLEN4dg</VV>FF+
eaORRfR=XMEM;Yf2NYO9),bE):;.dA=Q8:BaFRE-CDGD7K#SgLTS6#@<g[d=.A?/
(]AIeB83;P#QSB6SIM/feI2HL8_RYNJOJ4F@UX&><BT<P5;^AA<12)6Z(;:?9D-g
QSWM[JSRD5b-MQ=3L)61UVWg6:V)eg^E#A[4&YD98&AL/@#HD+8S,#^.N1B/+Y))
V6D(]0:88M8B#R4EW?3]RG.2g8_B)STN<14,D.P.1BIb#ABCKb?KH&Qg);.L8/b/
N_[:W&06<:&(?Z)JAFK1L94NG[LbDO>@#P4a]_XLLZ_(SZ1M[KVGa=)<00T@cEER
NJ1&ILQ57Z\6P\_QTFD@YVbAUY.QH164M<P/Me[4-URf+d^,JL(GI#15(>dG>-O+
P[S^5(50U/MX6]^)H,TMX9(4:-[5fM4[K,^HeJ5N\1/O&aREQ_d+bU#cS?cA?<JA
0,N;XYI3T-/3H5SKAS=aIC20,GK)=LP_cZC&SNS9#[Q&87+bB1M&&]8,()e0E/5L
G0/_0-&Z]?+>^gKCA0&_,Y(OY_a#]9;cCeM4M_RY#f?E4O)>eE8eA3OE80>=</DG
IT[;6;d^]I[U\DFPf+KN#-S4:K@-51&.2.BW0a1cE3HZAJ1J]afU#g.5,U+b.7<D
acK1Q2(MI3#TaGCC3<E]>\\]&M+J66@;@?&BMa8f5H,X]:<?6M]O5QN>B\2Ud#UA
Z#]_@\e;UX:PFe=Cc:fZ7.K-#->e,e1)O\2QNQOXfG\&=FIIDWCW2UWO3g3fO&g&
7AQ1Hg\=U,6Y=7P#B#>UIg1U#DOINTH_WRc;92).L5M63cT>ICLQ1S@,DRZeKK=W
@Hg4=F#EaZe-4C+QTEN3gUVSA\<MM8Nb2L@6[84WAH[c7KZJb:e;E7-)Sf18J)XK
gYccFB79/;_K<Wb+a:SIMOTaVE;&PGReH.(\3C#3+]bRA^H]3LU0Cb?CcL\)ZCBK
J1cX_?0,f&3:<,F<S[_4^<T2Kbc[R/df1/?BGG[4TW5;RH?aS_N2C?b5W(>NRH-;
VM<5[1DY=-TU/g5-]?T1MPd4D/JB@_]3g)?5D?@_5_=Q=38L=?GY&H]9Y+^MX3@J
N[\99E&3JW7&dP_VI:)\c9EXL6=JAH5=I>;=T535e]8ZREMI09V(^72E3,ef&7;/
Kf8V_#MRI.9CV,UD=-JXTbf=TFY-;B50G#,0SEGbS54MX1V>+6-a]=6I.[B-EKTL
VF1P[M&2DC;/PYXCK(MFO4EY+82I(;P[:+F/)>@S]52BBE9<?[:)C<,)KSIc6386
IYG)7R^Ic[YXH_J(&>?]UD87J@XF>[#=8e;c:^WXK1+N_(f8-<G+RP\O+2d65S7G
9Ab\f1HcQQK1=Mf,W,U^QdI\GSf?<DZSc;TXQA[=cK^8dCU,SMSDg\0-O(,4I#J&
+NKg7SUT[>Nf?+BVc:7H@/N.\OBAZ?<AHGKf[W3c)@V36Y05C<C>\UA87?(bJ7H8
I<(\:P=a_2b+#LGX(@28B93d]aO0^KU0XZ>J/7RI.?PY44;STI/5cYg^/6#&VDW#
O>:RJBfKRdR<+2E38V1Ef9HJc+A>HcK?>#N@@\E#/QX8PdfTCeJ^)]8(fF7aOR1&
=e-2.M5GOJJ:&CBX>S^U+DG<^;/]SH)L@Me+[3[V&1P=0g9]_7.ZN48XQ_H_X2#g
&S(+RAbeV7WgT)bYYd@.\^Q3c,SP8B]ORDagQV56dJZO(5#Xe;5>_,<L?G>CID9F
?L]3-P0MHdPM]A@2TN(33>975#.6KH0&[#HZ7T_b4GR5RP@-XJ@JeUW@C&g6#5Md
Q0LFgT66KN\6;S;66G37#W,HXb>GB:G/\M8B217bB<5=>KL_0>K3(TV1S,ITV??M
UaP06A&-gD6M(\cCANe@a)IF;b[#35G6gXKK2N57E94+=KSI;>\?JQ6XFIgU0RM5
<c/SS^DeZKV;=&BbW?\4XNVDWMII^]RS/CUDCJ:6F#L#e]>U&=aAb9#_Z<HAD)2J
a(ORUNBF.I?<-&JI@;+b3EMIYe\a_]WQJ=7DcO/@^bAgLGXCORM(Gg:L9U&9Se(,
.4_5\6gE2Re4&4S(H+^EXCSWONUf;2R2D\Kg4#-7.BF(#&;a.-3+6ZCQe;c5>]9_
31WO13.E]W1[Q,S+HEV5(T9Q,X6N#2gQ037_]Zb8D;f\#4A0HVMO^]TSCUcReD2g
F3SIWIY9HA:WNEL:OZ]+DXfeJV.PXIdT/5:HEZ[62&SIbd^T9P@Z0H\>TD=KU.PR
[g(gVJ?R,g^_O4GMH@34_4[[U[P6#A[)?2-65U27X3YBI>60f4=gceX&6J)3Bg31
=I+\89/Xe8.CB,E.8GFGX+&S=R]P<[<c&MP^:,g9C9S[dC]gE&Z\^Ud@3F;;OUD:
b^54WN(Nd/KV55cADA1fN)@Xd]NH+\N(X>N/NS0d)&IF?#548eCV4MMJfB[&Y0&)
(>[Z#1D4^SfM-=WJJ3?bNe<N,UDJ=WdM@1e;&I0,4D[UJeDN[<Q=EfW-@QREN3F]
3,JJaY+CUI:4D@LE:Y9DeYQ6_.GI;XdYZ#eESQ<cN9XRB?7g?QJBCD\=B+Z(FXK+
L9bfDZ+VBX#FCOP0cI-+.ca&4]c3[6RZ,3]MT?>.ZfK5aM<M?P0)6A.cVb:+^,O>
Y&[9Xf9HKVDM[_BP-H-2D&39c4D7RMBML191HLF@V#JH7a,APO/3I[(NG;W7+(XS
e0./b^G?=+P-4M[60\AeKa&88e8HAIJ2B^W08)#PUR/G?[<MTY]=9e5XUc,(<cGb
_Y1_9E.KBXCBaaS>dNg?3CMY1D@bLT\&WOW_1^QF1a5R^8QT;PgDC4\D=;WM[QSQ
QIV</HJZ,])>g-;G1X>H;+g7MR>DH+e?W6E64TdESUCQWI.6e1+TX[7>,cbZYBP0
GRYB6LB;Oa&47E3/B?\V/W]FDEZ/;fG(5afD25.b\^F1028dT)/HSDQY6MeYE1Q,
PD/dE&7?gLCYJ6?g[b+;@^.-CU2E(?\:O.<V,aT6VReg<DLJ8aH25gAg7\4;J+ZE
F.<?^&3)Y8>564f?##OS/f-/HWI&BCYA#,,580Z>0X\[8XGCa:Pd2G@0OP#8J@FT
>+Y.dDK[?A1(d0];]MeaL#JI51<JNVY5gcGJ(7]F<R;R,cfD-1J)2PJ4BV4a;O7R
GeY;#1-R/],BU1U?S&<_8f29<Ed@=b1J(<dV?:)DKa@RYV#:?/G\L.206L;E=A^b
IDFNXZdQ\/QG+Kc:/<5AVJeJ[+@L7/Lb&-/W&B4RO4RU?1Z_bbb\.D#M1>8ed^^(
DM-AN>[SZQd?Ge&d=NN[e<-_5QKCITII8)07O1X+\]Jc-MR@(5F;M2[;__LPHEAB
4PPcMIW+1@Ab.0>B^0P\>A>:,P-<4SG^V=dedIgfT=F2+-eN-K>e1I#c-:-6gV:,
3#1_ES/Ic.]WW83]4/,UWbTGG6&VbQ6dFA#A^Z@TgGdN3)3T@<[5W=&E;QeY2@V-
acU6212cT31UeLg7U<?&JI-Z=0SJGcb&?7F[YFc&Z[ZOf-10^BI;X,J5P8@^0LV(
_(8XJU4Y.R+ZS]98&[+),U/EJAWP#a\[&OL#0\8U1Z]b-a4&RG<#Dd7d.&V<K-H3
&63#H\.MP>:FK,4Q?^bJ[0Z-OdaAY0eJ.//SU0a]@1QH.#fTNI?.UQ/J8(P_KMD@
-bBGZC>Rb.=0O1ZN4aNgPf8Ndd^MG]SX)g5^DdJUPg5V&&6L@U(\/[W7>#T:;9BE
@(2^-a_:I(6e3B=KDFTGL//ES.W@1.aSW8E;)V/9GGKHIfZYWM]R;dN6aY96GST0
L/(Y3a9a0dSEM^BFadYT>HEZYR@/LZg_ANaD:GCQ6J7.1(:.+UOcI:NV0f,LCB5W
TGUK1:92C2]?T^U\.A^d?cMA607[aM.Jga2E?JQC63AaXg:a;)NE8AQ/;9WfJ7E)
PeDH+-@=;T[a=M[0f]ZW=MWg[:Z]baZJUfM\=Y=4BOHC:C-Y0:4U[^O+g<G>]..D
>FSG>9[#Ddg3UUaXL[W7[-PTUM.3G-C(9aC9D1P_.4_??I5<:D8NZe<YJgFAb>Fd
Bb(TXVR]NUW@2G8[87Y1Y=4,bVE/MVd(C9R#gJ@2LGYVFG)2:.S;);cf6SLa6A<V
OSZB\A_]N2P3:R+WPKYd>92b798AI2N:eYSKK2C-D<d<.?Sd)D9ZB#-W>B+b^.^L
)Ja-HB(=GT03OBU0\eY.eR)6bX:B1O67E=?g_BP_FJ>HgVVACB>fUT.L76/>F])T
RR<2SB5^6bX#XC,H[6]\65ZDF<WWXU#0/[a@U/HL<0EAKBT3(?d0dgZQ<;f0ZQF0
>#=#RQ=5Rb17<-L6-d9#GR/HK>Y.DeI;^ZHI;X&Ff>AE]</<7e_K/64V]G+7Sd/A
c_8V&MYX?NZ[7VNZ)FEH=L##b3AW\;U,BO,/U0,M0@UWA,TC6Ab^(a@\febQKIg<
>=8KPL&VC<JG-:9g2&g=P-P)SW3.XI>4Y3cY?SL#@:.]ZY1JM0-7S5IJC2]3Z7Q\
<V/7]3aUf>VI=WZ;^HH&7EA\<)BadONERNT&06)>\IDJ4KgK/Jg(SRB&-L8cJMA;
Y\X5IB7L5B=.cLZJ5N_,:V#,C)>:dcdBPSRZXEPP3=gLD_P&Y0TbM)[VR6K?J6M&
DXFb)5_WY+GBc9.YBB1]-gW&>F5ZCG(^EJ,9?]2c?ge8ROG4g+^S6eR@FXS]O6#-
]/Q#4)[g>(?__/_g@P;&)@faYQSKEf)^3GF_eBb#R?L>CA4@+-L)F<L.IM7VC#[b
\a]9aC+NKYO,P04LL&+).IJ:eKK.=?+@]BKU7;/8[+HT&GGWA@e?I;cI;bJeV@9g
&JTcf@U7I6\(S-B]QC\.-ffYO#g?Y\gL-5HJ4AS;X=:g7CEG,TA)\)/WAHac1CYK
^J>9.).\),5RK;aC+-LG,g\G-K#&2X-63UHVeE+LN8e>Y:L5CcNNfYa5R#>6S[;?
Zd<4Vg?cU+9M>JHfV4<RQ[]1J0I>G\1;c>TU01&;=^G0/?.a&@2a(^?KZMKL/dI?
e#06K2_9=I1N2cU9ASU?cZCO/\?VQfXW^>e&d?=P)R1@OM\O0gC8YQU1ZEfc7.5X
Y+e>D+XN2MGcG&Y4^QPc-&)O)?YC<1S@0aU:HP@Q),LTTRJ8M=P7e2Q7:W;D1C>E
IA8a<?BbX9bECO;7?64FcWab@ZLbTbG7=1bYQ4VVaPNeRGeFY^R#BXCJ,aV.)L7c
<9/-2#7VScf^QV/1fXA4HX[)I.EMDac\G\bFF[>-YC[\N1-eb4..VQAZ<;OZ^,@Q
F2>ZE_C/K,KGO3=DV#-S2S(+A#LUagdF?UQ+Y^bT;V7(gVR#JKaIMF>E>>1F]BT)
5_+fQZ_(.A,Ec_W[NX-FW]c9CO8Q9@Ld?<&B]<eNbe/;E@c1W/V9,gJ-UCg-)\C^
L=g8G<WM6ATCeSKd#-G0M[DWC)J;P05(6@D4NI,0cePN<SB<V]&W])GTN#YIYf2e
&\CVS?8eRK0fHK,cAHDN^.E;:Y,7(=G#TC.)H#[O\JNNeA2aDL?J0_>7aaA:K[+K
VN@[HS+FgXRLMRJFYB89ESZXbJP_:9M-)6\<U@=,I((Q#O/R<=@O32II-Qb<^\2G
.]^C,J+^MU[-[gO_(=?;?PCaVU5ZILdOT(XIQZ_1C]XCR_>C:EB=)V(bF6-G#GdM
9b#X(Dd:OLKKB6LVE5(L_Q?e.7D^.6(>#U9[K6dSf=6<P;(C2T-O6_S^0QPQ0BQe
XgRR+/PP#;f\=UERCIfS4]\dc^3P2+YYZfTf]GVL8BDO6@]@W)0;]WP/gbT5KNX3
<2&e_G9LcDfC-,4:B:0g&=P=?D><CMEeV9O+W.I=b--GJLc]OLZE5I3LW:MMA/Z@
.NFGX9]/RaWE:@^JI?[KTKR+05>,:G+R5_=ce1R)BF::C)#VK-AeXKTW:A_]aWXZ
4_ZY.UYGgN&:N;SK_dB,&X-JRdR&f?)3H7O8_gP>)bPX+bB85+587Wf=Y7^Y6C+:
3.ZMBf[&SQN?^0S&)NYCT+Y9V^N;@^4&GH&OA&<)V\M]cce\2^9&Q,HV\PKS@>Ob
V#V(:FQP)LIVbH<;0\T;(VQ;fXd2:VJUP#4e^XF@a5PT6bgcYN6-<8(FP)dOXNg+
gN+XLMf9#JE)+SV::)]Y\7^5U&IAPVfa,;XTC,Z\4B(JM7^#5R).X@@8N7LWN0ag
3A/#N[7YceC<ce<JL^gLfN]S#O2SS0)d14:26JeKCEXdW75V2E[FbBbQbLA_U?]_
M/=F_50[92>A/:9B-X#M<-QR,Z5K.9E[+NgV5=#)&8_e3a&I4SW.7#2(0._-c@]R
a7ZGZB&\eJ6<X2&QTF)Pg:6F\aBJU=0(G8.KZD:&PZ4)c83Sc1T[RdU;)>?G][.W
.L>#f(b.2)PD^OOD_92.,2+17ZXSV&8g3+Y@52H,eLB,\3U6KRNIQHS3Q3<aaB1d
8b6e03CR6,@#;./GE6_L+?@cG@4.7+9_1/VGU\D+L#5d(Ma^85(0S62dR&g;F#/d
33X#R#(RCGH00JSZ(5Pa/BBU5SSUZDQJOQMOV3,.20fPSTZ6<b=U_>gP8R:7.1d)
5e,SA]@74:3+_WM>U+g:/Le;F8:&^X6-7:f1I86\agL_(HeZ_.)eAfTHbIX70LP-
?\22/a91(::E&1D3RGW&NGS]_&_JaTEN:CSMAPbV?W/QLK_D5eIW5a.CX95&#0PA
T6<LSTB^-,05XOZJS;ggD8ALA2bFERW4+FRb.40)NTK@8[V&e)#-LEL0]CFOOP/.
5d8M(M3+>S4#[(4PYAURg^P8LXM20[.BJ7UQPU,FB[K]/5fD#-3,^2?NOXIU:BJ:
X\:5B=RIWZVKI@HTfOJL<._NSg(TU4^CK>DfX?BV[G9K,b>WJ01D=>aE>6ZB<^eV
3d-e^^WM/=M?2-46QFMKR7?(G&P;3cMLGFA18A&#>YV0.U@b08T4c2RBa[M>g1<0
_/HXEH1JT#Y>I9_a6=MEV4M3d<V+9XZ:1IL\Wag;LR;847XM,]1eKaKaDd48f4+c
PI\g@f]FH[<]3W-PZ(X823&5;\_)Z67gdOK19_[;<J5C7O2C&F<H8623OHdc77fQ
fP8:Se<cd8d-DNS+NWELRgU]U_P[JBAT).VG7<)F4IDG6_^XW1c,,_R1M_PCI8Ve
U:I-UP3Wd]dKQJUB#Z#Jf[]U[V7,9QIda#.FQ/-\/^Z7g&->QA\::KAe1W[g0@5)
,VI2YB9=d7M=Rb2dfOT]cVe[J;2#(:[-N>-0BCG[)YQE4:?HG_&1Ogd0P7aSdgG&
]8Y#FFb1W9X5(3a1c\,/;WCFg_LECWb/B=+b+b@,N\FS+1CHMIS@;C#XC@HP6]ND
JWFF/+QU(6WBB10>cR?4YAYTEea:,812MNN#DNc/Ia=I6;0,#&.DC#(gMV2(6JQ?
>-EK4Mg:IY<_IdMNEaW)=]RJ#X)E:+S-7>[9V+7A=B]@1;@P<;B/_[0=bQ-1+67H
Y5^+1c<J1=YK^b-6WZeP-3982;B-@<+_JA+;-(<?9g?B?6M)N4L?38>IZKgQBN61
E:b.@^T/<7C<RY,=3eW50[6-?-,_,V]V+=;F41F6ZU?0(IEHc/eX8LDS0,3T]V0f
E.)3.fXTWAP+BX/\8B6RP=aTeAGg:@/?7fU,,0LQ;QMVe&6,_M5f3U_O+6EQ1#7[
3^0UP1[O97KNRa-YFZXd.<e6_VIW[SD?<GdL:0>F8T&\_ETJT181Q5e(.0E3Q_^5
5IdDCGS[<g(b#[Ob3CcNbbH&fb>Q+78O;20#@[5H8:&SILS5TIbLWH02fc@?D#/K
cHcd\W4B[GDOB.7\Y)3]LC)G8IaAX_BfPO)<dMG7Q5fDdaB;;0D4;+8O;f6./_-L
Vd^WaCLP?TQCTJ[ab/8bLTU=7Ja&1L=)S+cbWg;QH]F\CC9+gY)A]))#&5SKOF<#
.UfF&I9J[:c]GbM<X\MI??LRDR^-&=WJFY8LGc8#WEdgQD-JD,Hd[16C/>=eNda_
7+95K-d6=+gW](_E)Z^0V&(R0T:6L,=I1X_S@)@ST,F8+GQK:UTYS]7N#S1\15#M
(07eCX]QcLbB#VF:7&JZ[.Y8)JOSeRE9KZ^-d0H71/W&.MUeeHJ#/?I2V::D9)0N
OG[,;_Ndg0dD<BgQ(Z[H0HHaRCQ=JY\Ca1X[eKBLJ6>b(VJXX9F=6C&8/ZJGS>d_
LbS64:)[()HS@[(2)1)^(OT\[DR6dJ);PI66RYC>P65-gWT1KT(,P5])V:Ec#6)_
#)aQfR1c&_D4.F-I46QKG;N,?U,8bdKWY6B@c]ObfW/NJAPQa==SOU2FSX6U^Q0A
3#UT-Z^OI6-LS)^cd\3Aa,cI,d2W1dHDTYC@7M5TG9HD6J#L&RT+D-\B^OZ4X1KD
Ge-1\\(9]ZN+@9)bG.4Kf]L#[aI6DFbTE+4.VgYO]aEQSP_,cS=]XP]>DbZA-YPL
^[UP#;[OF>168.TYT/Cag(?&D:c-c+W>,6[A6PJ>Va,8V=,XfXQ:bEM)JSC.4,bU
XD__]ID3^O<FSZ=NaAXeRC<1=g:]GY#[+9g3J;3?:?a2O9IdVY\OO0/BU<J\4WM<
90f=X.^2cfY1,,B3?b(HE:A00+.5S>4O^NF2M]ECA[G-:;=Me3E\&2[3402&cNae
7D<XC-1NG5K2E<S#-d863P4fXDa[1/56(W<1T8TAdLc=C3#_/cKYd3-X3]18?HY?
4)CQNYB+F&I,_2IAOQ)FPLI[IU>IMe\17?bC-a5>)G7NO_.MH?K)YMT\Hf8ZE^#c
I=;VEd?UH0>&UC9VRX52B3MaPF1._;9LaI#T>92)6Lb7FW6;2e).>&b/dR<2BAB;
/b4c=87TW\KC:/cXEAKJY1XB6.&ND[KeA61JPQC^.eF=b8&L\03Z7DV:W]^0:A>Q
c>3Y4OI\[IG]W,KZAN9^)MC/?dTJXY#MMUPf2VWcF=0(]RE&:H4\?O<ZO<_;OC&f
cP-LM&Y>934e2d@&459?:@Re\@\0)[+e,3gAY.3+0Z&8?eF)77L2Z.Q-M;L2LD6H
70f.?:=9GSUOKKZ(DU.,3T/ZXYYfQMbC6:F+QSX;T#YdD>Ca<ANa\:CPa5VOd5<\
F^,8C6D^5IBfC4#)U>6c;/&)/)f]PC/fa=fbU1UARQ>HgDUO6-71eK7AdO]+EH-E
1/;<2bG&NNe^X@HV@V]GD3/#MHG/+a_7[Q-2#OcJeBL(67VJ5?;@FN^=GZJcM7WI
&O95VREO/D>Q@,8Yc&1N9W5gTdA7NBJgA;L5I_HML;QBYHF?Q32a@XcWG[T#UIFW
Id<BB/AggKQOW.HA;NA]gBF,QZZeb8.1A_dGJ,+\4[R=U+YaUJV,,Z-,8V1,G;;K
^cM=OE.S;_2XDWHLU28<9[-W(.VX-Y_,;J\LXPI2481W5=4a&MN]Z-SCZ>f<dGb/
Db</,]<;IES,-gI+\e.e5e#GU/-fVZPDBQY5<0eT?4EEVO-GC:].,2/f78T+^Xd4
1,,Yb\S)aSH(U1:cR^=.5<JW3dUZ>5MFO(_9;6&#AQRQGBQW.41&E32g92XI@UPB
UKZI>_[Y&XS5^](,NJ24]A)?Y.-eJCJMOE(]S)0J[YRB?,aP>VNT]#&Q>f+a#S^B
3GeOJRcZSBUT+NX6VV@RGb=fFCVd1U;TD6>@^KGDRCE6Zd7&\MEJH@dR>=.RF&^F
IMC0V^)\8:4Y+6CGZ;8ReQE^bB@)=;+7=3G:L54]+;>eFE:S?S#?24S.e7KRPRY(
PP^55A<<R5X+Y:]]9;&NVUB\TZHH<eJ;)\5V:T0+>.GBV)=a[V,[bUD>YW9JOg=H
4K<M2VVc46a9Y=1>9R/F2WLD/,F0+Y<aE5(:OL;YF6U)IXN/(Sa1BF(\#I40,XX\
9XGN5.VY0O-N,&O6g2]D[KD.\\(,WE5gg(I[\0bNc9>dW_P@3FOS-+/2Y-54:@VQ
<9IR2NOgB:6.bN(0V4>b44BY^fC3aB<^[;fF5#5JQT5a-;Q&F=XZO2P]6K8+b,g,
4@#;:R6[K5UFgE^TaHAMG24X:XH8]0XWD2,:3gJM7CbD,NDgO9ONZGe9dUX?AWC?
2=WIZ.<KJ5;M4DMF,U4<?XJ92?DD)\A-2^7S=AB2OA8?^H-PD7S9b^)3)#Ua5aP]
N-.Z@.01=^6dgeHO^[Pc&UD5^43=W2=[@,cdWCRa:Y>d3+)+_&(d6_1R3]<^CW5>
7ceU:PLU_2WCLe3+^]e/2_eK90_8V+3D:-d5LdWE1DLBD_&g]>/792CMR3>I,BY@
^6C;M?51R@7Md>NCW.FffacS-ZH/8T^DZ1L]_(fVX?E][WCY_c<c4IILdKUKS@H.
c_PQ-&=G><4HU/c;c-_=aD(0QBCLb#U2F\X_T/?5RAH>T:1EMa;b^_<;-<&/&SeD
0]I:Ze7ce-J;D>f\&7<^<<J:WV_4bB8OFD))>1AXdAa@)0\0SS4;,^/XgQ7BKIFF
;XISY2c7/GC]&;3g0@^@3J1.cMcNB7>42WT_E(4T#05U8?U\P^1aSPe^VQ)7g1F3
Xd92M?7\EZ7\R99O^V&1=&IS)J9L0Zg]77=68:c.R1GL@YUVUU3d\?Sf^IGFVe2K
O0H]^A9RZ16IL7GTDFbU.0\\#KfBJ6a)O@dS\D9Mc#7G31JJVOCgU-<?c,@);H?S
=UDX43QT3+QH&YdTQg57XF)eL?E6.]Y.2?@UP:F3N[cMbK1C3=61_.A-U]a>)=S6
[BN?C9HY1=#KS2_&d<AX8;A#TQJD](Pd9QC@[DJ@D?>C8KdH2K.(LH3H@;#4M40L
MTg<A]3bM1>=X3+GYe_:\KbGM)PE;MPQ/Qa2^HJ]U)PKC^E/K51cZ)f+B>81R,L0
S_AR4fS#aB5c6IB81I:5J7LB2aQdDN?Va(N,W0,-bW0Td77=cI9:6,IO6;)1O[c:
8V27cQ>RM^BJJ#4MAOTfN2MYcTQ_D(:Ue:7+26b&A.df31Ec@AN.2(M6)C<+eB_W
PW@5>MFKS2cM,&/DU3I:1V,:GP@Z2.OW>WE,+gOI<+8Q_C4O\AA@f_JJY.X@VFFX
WQ8ee[J030V2cRK-))#3/&)NA3#6B3M;PZK_.;HI6@@R2B\fUB@2ZOLYNJEMR6F+
28_26=295?\Lc96HY9Q+@SVNZ<<OD#X@G7KOgJ.4f;=V;>Y?Q9-DL?O+5+NM8U8W
PNL=F0B/X2b[eB(-AD?N,fK/CS;LfY:WAa<U[0Q@E4G@3,IN>:f:ITfD:1M\RLSb
<QU.PFd6=R.#bBW/I]UIX1;;<X9HbSb[SAQ3)4^_RC9H9]=(&6a.F2QN8\QB.0OZ
=L^;fKMJM52T-.g2>96Ug^Y9aK901NAKQ\=AVfaX#agebT]:Vd)S)NK1AFD,F25I
8FLbc_YfY<LC1f>L[7CMfL5g]-O-gV+,CCCKIWD62\[/c=D.U8e8H\6RZJ&KU,fU
9B.4TdO\WSV5G(,AXHL1_e]d]=b^:Xg:>:320/#^XHB5SQbOQDI[\BXO6ZDTW4J7
0@:G(D2JcW0>O:&(4e8L8;=D85:AIce=T5/VDN<56VCNOf,N_PLQ?E[Re]9b.f/O
GH/^YaZOdZ?[ZE8V17GX]@1fM1Q]&3=b0gYH3McDd#f??1-LePT(bB9bOHWIF\Fe
@^CN@&YFd?;]:LbU<_3JD)E6C-=Cc5K(a3\]20C-6NSf+S182BW4gK[.IdZO<W?[
\78^64d=D^EaCQ]b^11_@[:GE<Wcc[gg&PWD^8I+&=H0CJ<R#(bb&]A#K(QV?+18
dK&Q]?)NJ,O5fYL@]4;C479L?:NS4f^=e=FW&P+4T(W+)8D62QeG-^?D(1+)J)F7
1?-</)c/W9V(TF]9b:+bYc^U(132/Na>aHICXM\PKNc:;&a@GGeU8AV[^0c.aKN(
46TfEOf=[;BdK;_77ONV6)7155>.>UU554NQ-9QBA8,>06<?,--T>?YN)EW3#+P5
e8@EeS=_^d&0GJg,DF<.\(<&dBg.W4]1;C:7P=f1W9-7[\0<D@KA^V=Bb)REEbZR
a?YCa?ZLOC7N((bP5S<BCAY84aDV7D?c:?GU#)d@(/8a5<acUQKdRN7>>V7;]Ob0
3dc8D/0YPT01Zb>9#M:18>EZKUTH??S2:2cUM[R&EE&+;BJD1gK:8f1E#H([]C6b
:;8LD\?H<V.-\(75=N0-YF]AT:A+>dDa]gJUc-8dQYH-Md@c9+OR&4E[#;JPS/Y-
^=P]6ID(f@LW9_95-A8U]aWOEKAK3La#H7PbOD[V8F0#P4g\QcZ00OZK]B)R.U.M
)\O#O]1Zd(C2+8R4@BU)J3LSXYI?Z]5_]1C\K(XLI8KUYK3/]QLXE2?EBZ0HAKAH
-FGN.6]SIQ>faT@_6>.>>[;g+_R)cZcfY1[4NZ6C5AG77G8B\D>0Z(8#Gbf0JPcU
?OZWM,IA?d.HZ)8+Uc77T@7FH=GNg_,KYMLBX)8d[8V=98&;PN]-f#MTP=VSPGD]
03>^f3D,.QU(V5f_JaNZR8@.<JA@O1c\Va,D/SQ2QJ7JK,-A)fce58,7J&K7b:<]
3?^fab:ITQ&aKZ?K/>9C+NQKg4C<HM?]^9Re+-?)])D\4/XW,-H&Ida7&]ecPTUb
fSMNGQRFfR9\41;([4@/4UJG4K_.E3#a15V-XY\X#SH#<EE^)gEI<A3\2@Q-1H]-
6\>(48BA]QA1Bc9:J@IfNf2OF.Y3aS=I^1,#b_3dRC8)FJV=@@L)4EI?ERIg1L#d
N(YLJOBDZb7BZO[HA6N;X<Fg^G.J7^#RDC/&P\?7TOg7LOf#HMKgSV)bMfAdN:5)
bc,[P<RD.>.3QE>cC#L@NZR0\dg0W=K\7c=e=XK)E#W6YVH1+?E?#8SMId1Y?d1J
M]=QL1I?C=VXbGR)?[2+^eV^8K.dfDXXG#AK\@a95.BN/DFK^8(db:g?ab[fY2W)
[g<K]a_=Ybc)a9Z:/8:cMaWINIV_fV0O=Y2UX3XQ:O/+;;;251,[?#B=Y[&7M?Q-
VJ@1EEM75EP-MbAM.SLOcH:M2,3b,cI1(DMc\AP;Q<f1OSG.;;QQBAUeef&D>=R(
:/9CFS[V9V0Y)[&H1F+;C2Q@:L8e<(Nc@+R][.\8f).VKfe_+b:-4//^ZO5ME.I#
:N^N_#-U2-U>U:E#&(^[MY<7gUf^#>>>.Z_LYWN08XOX^0&8/F\X-UH8fJN)=,I=
DAL\f]e&\0-C^5;Q#VSF:1dgL_,>b9KUc:[>B[T(J8&\Kc7Ac+EaN8\@9TBW]dLQ
8:3I;cKZd&B),9B]df+LTX[S&Gb)=2X-XOLAIFBU[VZF4?=9XXf3Ga9[_DP2W8CA
P^/bDIXU<NHT\Y<GV;f]-?QH^GX#??I3U5HX5?^+CJO?-#&I)KGaX/Q4+QL:gJE=
(WaVGF;7GO&1^?GLCJ.1SW<8,0<IUG56CLg@O5#MEAfe36QRM:4.#/D/MN>A9YP9
YQ>eH9NW+5G345(<cD;RJ)4&5LG8Pd2dU5+M(KIc7G:<OM3(Q.eTA&IU/NK?QKI6
+/NEZ2U6&8d2\ID],/V;bCYg3agXgKeU<8@8-]W?dF>0/bY]E=eLO30FA&S3bT5c
A8WE6=OPNGa/a+B_\&=e-Z==-P@D_Y9VM=@)Bc4,3M5cGR7Ed&B#:09@:49J-?T0
5PX=cC-fBR4Ub6#;DgTQc;5:++KX;8D#O,eFL/-=N6d?^;K#17,MHC;AN2G31cC5
JVddYXDX,@?#+FfCK_@L2D_V0<6V.I^dR)#Ff8gX,f?\;XCa\d2@eZ8#RR\6eNee
,b&Qe&C_6#+M_.IYdD,eFd.6DS(d7(N:,RF<VMB/()?Y#AO8[cX+B(Y6g10ECdN_
Z./5D#0Q?KZ[3]TV[ZO8P(TK5_fE\K[H&0TL<HO\W5fGKLD>Wg]/ZBgQ+d?T5e^7
T9^.9dd1U^C&P9=HRI]I0(4&U(Og2,:AQNP#^ca&S-e,A/ZO68T4:e(J/c&^QEW3
RBE963K[g_^,_fY]Z>>MQA?[;aVF2ZKg1\-2f#0/@N<P@(1e@/NTV@9]3ZB<5T\e
T?CP]\I5>ZEQCe)F]IRbG0f>5.AMH=QWV8J1.;.?1.[+aX[D\4)PC[A#7&D2;c28
\0H4U\OFQ-e1bOAU2eeY\U6XZK=]M&bIeZd=4HYB<01X(3WRb[N.[a.W)UC866bH
/Vc\>bI\?>YfVQ<S2D203)#<;R=+594N=49)\2bRdfcC?#6K#_<M(ag]3D98Z?JH
B&:+gNc_5Ae]8HN<WX.E2Rdg+<DHaULE^TA^;If,g&21MYIH?@Z3^Z@R1>4We)DG
,&-W<-FDLN0X,Q>(--_3UH8D0,T.CT0Wg--9=#;53JZ@9B<DW0UPH.c1/eIf62LW
]a[<A#Z>PJ4gM8Pg=G_-\N<1J@>959X)Kaaa\^+N+Rb&BHWI)?4O9.Y9/gF;5A=\
<8UVM@BI;\@P(-F\V@4.>\O<f/\c7CW7K^bD,W3N\SMF2GZZQ+QG()d;0]=(5b,\
d=WK^C?\U6g-?IJ?&VN?VQ8TARDK7Y/0SE2YEL^]#4f0-L-P0DWZ1POX7,A@/QGL
+2V0Y),,#c/=?0^T524B-GUeWP3U5B\;CS@5PF^^KX<6+=^QD?Mc2FcM&?c5#,9E
J5F>9cDRa6fgTMJHEE-T3VCcQO\]S+:]\(F=-]e)+FE6RM?6_eYcJD[W#&WG04DY
XK:#f.(g+gK;F4A9,QI:+7(YR(Hc6W;/F?=Z<N#bW/fJSS)Dabb5;;66#-&a8I@P
ab^K]X\B^0VDY^DHGH;//NgZb^XV)c[R)(9_71c.EBA,;#>fTY1=<8MeT;P(CI+4
UO:EdB-6LLSS[=-UQ]R_d[A0Q2fH=T?EEADLb/:ITX6EX?K9Uc_b.Ea=bDH>L@SA
38VDeM]@HWXBKcQQYKIZa&;;IAW1C6@U(B.B1_;3]2)Jc0,3W0[Jd(N8cT2f]OD)
ga5_(:=;?L:9=A>5?1MJ^HQDZf#0H?9F^cA1X)#VXC41:3NRFf))[]B(fWeb(Z16
I6DE1EgGg18-]7f@YZT1@4A_OPg&RDGJ+>)40__@9?c67A&fD]0N\PZf-_-f4EE=
d[0>V<J9C?H(@f\e\NI?+.Z?7H_]H:_.TY&J#/+LF?9J=DVYXgOOZ2f7SE1-/?Jb
Q\cM5NJC@?LZ^L5\R<([>9c=c#_]GB?\3]T8+6f/;QC[)H[Yb:.[G<SB6>O)b:b+
BU,65K5;Dc<69a@O5Q.d18N[57WM70]-TB<(#\0W7;JR8de6)H6>/_IH?,MDWaIU
#5M&Y58]-EU;DFI-I2#TX(,4eKUZ8CM8,>X^O4+26C=1C-TDP_;Vda>WF;G>4F.=
AHH=8[)\:/V1WN4DN1-G@](b/XFdWGT&1.Q\/WB0^9JI;IWbRTTRW\]&9YaF(Vc&
6W=A0JAGKUH6N-ggUMC<g-7/[)GH3B.&3c78,8b;RU/ELT^[Qc-]DP_cII5GS:>/
A^@:]S5a1VPLK(ee(Z<T6N3W_YC>O95,BQ8]G2QD6##S/aMEE_b&SLA<&K]WEH7.
HC?cI>=)B9Xc4L]OIgM<WMP@S+ZROb)<7\3<)C27+(WUW,#R\#Q(PJ_JXYQ#8(7f
ZIFW3UGabdcT)5\DQA8Fc2O^:W##A\;Q[F.V=O<ST/5)WK)fZ6USgK.79Y5G\[d0
>[>f;;PfDB7U3&cfec&A8^TIP??6c/59U+42FR^G]N9M.b++REc[,/bW5(#9LZ?\
3QUCRG?7YUDg8]fYEHV(;cTOR_b1CFF:W^NMeMQAR.&dKTIZcE4:JV6N&BEa,PH-
C8X16OF]XLDBdfU4dbQPK1OR9HXMI[F=EC<:FX\S,YZ]/]UM1-51=\8-TI&+H&E>
E1@>HN5[U-771g,.9#P3W6T)A7PBgU]-6Vf]PL/EFRKX1^?AMg=8JIQ&:CI52\J,
YY_2<7fGbVd\Xe8?W.5b0@WcYb5Ke@68ESO)_Of)];#DR1cH8\5;G[W=:I?OY3N)
^Y5VI(7&(T@gN56YF^4&?ASae296^XJfOR-NC33eR=#8cYVg3e5JbEUZ0M/6bL\e
/AYE?P;W(,fU-+:=UDH1<\85AQP<W?Ge;3W<9#>6R],X;MaGNX3=5cR[QPa[&X5R
F9CL]1T&6AEK^;)U;TR-(7VFPXI->Z]XUf_T1f?>)SdSNR:d?B<K)c@Q7[IW.?M8
8=5\6G?W9W3O=V]g,7GF=)2TSGbc4T@I04BX+#38=IP>YEW+M+[PPF9-=S.,-_-d
cYZ33@VRM]7AELDNWBdOF-aW2PK,e,eL6=g8L+\A1)^dP-GVf,+Y3_f[5QFBPf?1
-e1X[?cKeI#O@.)XLB[ggQ.a4V70GIFRZd],BfZO;LK<NI-W0)UMXP_X\((]f]@=
gg0+WPS7XGFV\a.N_J),N@:ET43;9<0AGPX3?EMY37L8EIE[fUa#f<.Of[@L[\d4
EdTF+87]GHE_cKd;cc20Q(8M;AL^P)b/D7,X]-(WJZ8RMfIAO/69,(^V,c,8P#Zc
YJefYT^?EIPGUCFWY(/NPW-FEG=CCQZHRO5RUd9[L&]E>PDHY=[8=GD0gX,X89gg
M4-;9GWIff_4T(T/;RXZLSH5_Pc=K/4CY/<U<UR9UbAJ-V#Z+TS.K92EV<e+89KI
c((@eIfHBb-MYF#a-.E]BTVRWPA71HQ)RdO9gDQ;Z\Gf\I;e=CL^Ic\D2[]Q.<TJ
_T4HZ;P:SbA0Q6f56;+#KOT\SQH-E>8E]/8E?K<@LbR&46eADa=3)T&-Mc=>:95J
#J[H7fF^7CSG,e/&&L=bdCfCNH[UH.4)0_+Ja@F:_.&,IQZ:0UH&Fg28NCIf9>b.
aPUC>2Q5:f@XGJ9?dTEdN6NCTA\)KI67)Q-@2PW;TI>CV#F>I\V;Q1PGVP??9;d6
9&PQ_&.Xa6B@=4QZ3e[-WM@6T@;bGa;^3U2+SEgX/01XSAWXZQ=TSD>KeMH6c_R<
.Vd6T[DF_69RRT#WCDO5(,HfIUPYdDb@AEEGBKDW1OLF=)+REW7GLTgU+2TYH#32
Q?>_^L//37-]b=JP02b#S1;PY#]8&7dgeAaB\9c6Lb=E+7Q^7[,#EST89A=WB7]c
0>DcM:XbKMV/5_<#1(0;d119<OEc/04.7X/aOZP_.e6a8aPV\;7]<MH^?=[Lg1(4
\4c5+:G>(V?(5/A3;_]V6b/cf>R2;<2c<8X[:TLEL9)(fX[-(OZVB)J1V3^HXW3J
S^M?e+aMV_>T?-?]fEecd0&C0]P]9cc_.^e:WGM>-B</I@F-fM;X3-;,0E@SM<De
0ZANBb360_H=XWa.3A9Lag8WWL1R8[5EUNf83F(=gO/>E65JDFfLfQ)JEO/c2@?J
:dK?0(G#U<D_<#1#<:+#UL\0X3WG17>\,2_36]5-QJ_g)3(@:;XKEK[LfB2O_G4M
LR#T#61Q5O4VG]GI3_],QBA\U]8_[C@(b1?ASLDb;D1HRMda^6[eg<JM3MGTH<,8
NN7W(CU4-)YC#(fG@5(.:+?=R.@8<aGc>PbgaB+S0^8[>C;Q04=f)B/KgV[fIU3O
=1,dB;Mg0<?D7a5:S208;KK(1>ad7#d&)aI6GWJM4c.(&ZZd3L]51QGPC26S/SMH
b?7NE\UM>WUKT)4@[,3M8OaOJ;QO@6=DIC(LO#,C;LIX,f6;I;1QG58[UR3@IF-9
HbaP05f^[Jg66SKO_^H9E9#EK@bZ3DV6(&M4.Dg[+HFT&X-G&.f[=QVaS5SARTMD
[+M51X_=g\@YEXg]dM(gK^)Q)&Y2G;_S+aK1Q-EJ>(FX9&DI(Q=d9_fR/)0,Y5DG
/cSAADHT(Gd=9^(H&\KQ0W3@G3_eF2L9b9V1TQTRI[F]@YOKEV)aTYdTR:S;G\V.
1;-1Ac&LS?:O(La-&HE,5V]LIgTM\0CIb(ZJAET?;C1I=Md]6DY;;MUL?dSLPa8>
XDJDLff#3RIV4gY&P^<9P&A>P)7OHJS?.JO0?:L7Uf5A_5_P88?QL;W4JUa=J41V
L@=?TUNKX&C_MZgEM0WZfTS#?e,[6eZ>+^\CLJ]:G?fB#6,:;0S_:RL+EaA<62Z^
.^40/[AT]104\PSf\[),G,_X)NcEO9ZOVY?baBN1T#Y#bKL?W:@LU,,:SCf)+U@(
=(g5DeKeNf+#Xf+#g#8A8bO@S+]/7A;WbX9J=F&X]A52gKK+G4M:]/d3?N.7RbB9
/0)OH@P=9H)D=2a.0C8(TGKQ#XW-;NLT5ag>K7I9H^-7^0@ARE1]BfTF&TBVf\##
(W<IH9.>=C8QY>8YI&#^&JZYWT)I3[,5>HYZSNa]EOI]P^Q5B(gT)ZK>SXT4RgVS
aWMF&4+^b)\L,8=P?aUJ\TPQF3&M/Wd,>N&c;XT0-?d)aM(Tbb>a)VX/E@dOM-H;
KdT2OMGPTDL^]RX5Q[7LX=8Ag15^7O4[-HgJIQc\MFD]C>;Zbf-T1]B3&,gI,C4a
a?DJb_.X:+TAJXLL[QB5&ZVb[<JbWbf<R8EJ^\J^EcF.LgL+(,Sc<\=C(=7E>C]:
1_DYdN,eT>UHTS.A6CWW^.HH[1D=e?92TO\DB<J]D^J-Ue0IgKU])fDK^3dE+g?1
/X_YZQ>\<3#eD29[KJgP2L^/((@S\EHVA>-P5V9.MJ]FO49Y,e:MGU)]K8;E5?ER
DW^(Q510Na:[f]c3&7b0Jf#)[/28@CM@S8^bNH.LUCg3HNA:_gAE6X1KK&24S0Hc
P-&e2MWYAD8<b?MS0H1B3Z,Z.;T<^(BZf:N=V,NU\#R-C,a.J))UFLI9OVbI?_+g
HS;J=]d.-845g9BTaUO83XA700VbVF+2e,R70,A,<RMfZA_AU#[39a5RRM/>]>Te
;gX1R6+_6,L7R#2B]9.c,IVE\[^WO8+^T8/X8GD.:f3(+0>aPbPe4=ZJ?#G;15:f
#3b:E-(MGM\gWU]6H@&K4Na9[ODdNaT.O@0dFH][QFSW2MJ]@dNB6W)]^MGc:?=2
g1-S/_ZbTLH^._7gFJPc.V]Z&V;fOa)Z22fcP=1XV6SH9(:==0O.b?HB#47FP^IA
3RJd.bFV7H<4L:;.VDW&+#N:/=4JHEEFg+CAP=W1UN(=\ZW.Q79^990MUIF5^aI4
TM,BId5V4Y3,?/94S7ZF[QDRcSUU7M:18[1/OO,[G8U5Rg@[aEe^8LN3(PJGg_La
)=B7)2\Q.D4)HOKNc=A\&0Vb[2eER^^e)2F39#d&RNd\R#=IW5fF8)bI;2[6gXIY
;YBdg3A&>#ZWg?Z;B/@^\?4Cd_M4NL^;\0<]N\SEb/5bW4FVQAM(L=UZ2S1G:d1\
De+P>fHRPe1eVJgP#c(LH,bgUW>]I:^]b>[PaAX;HdfSY8T=:YX]6646Y&BA1e4O
02U3E?L&F4GG:RgCCL:O8NTJ.3B#Q]NC2MV>?G0Y;(YE0_2N[__U[ESV>9F9^@61
0.+Lc(DcP:BMPY,G46P&\AEc.IJY2aC(b8KTLL]VYbA<=fU]:5V@OC17H2D=Y-.b
],EJ8EBX]&SC2&P>Aa>0E7Xe#D;Pb3PYUR\6N?DYQ;HG66a>M\CbA.=-f_ZN1WW4
^Jg/Q0-_V9Q4P1d3R\_2#7@\_-E.-Pe77DTb..J1cG:<.g5T1B\;Z+[RFegHBS@1
a>H=eJWG2U=#BHcH>FM101V:T@UOLBNgLY(0>12/GEg5,A)[#.aH=R12N#-<5a1\
[9I2)H;0MbQPbML<++a4@[\FZBX?e^-\N\;U?fP9:8)eebT.b_L+f[f9B,F))Mc,
NV5KaQ;d09AeMB@fF_FdUGLM6_0-?32K9&g]]0TP5X6CaX&?GgJEY9I@(&U]4IfM
1/Rb+Z6)(Q>9)D2d24>FS_WW7&^K=9&Z40>QdA#g^2SSUX5/L6U7D;^_WJ#A^L;F
>0PEf8D(7^Y,FCE#@GX5_U=-2QeY:SYcW4^,O>[UA7FD#0a6=X[MX+Q-6#=+PQ4Y
XHN>=?<gGD+L@:ScP;1f<d(/#V8AZdJ<Q^[@8)fa8V,K+H#H,SIPc2#J<3eDIV[=
D07F4K4PGBNOdHL>V+F8.#c2^T;eJ6.b7B@UU0TAF8XgGe.b:BE-NR>=Q8_P>74G
+7;ZDL6eIW58I4A,,O/):=_+6<X6GKWcF]Q3^^YULK@4?5=I+BgbTCb0<PE);RNO
/DLc>ag5Pe0Eeg=-a4Wf>CJb<e0cd[FQTM=TP[MO7TT4:TCd,gf<3(aC9[7Y(;2V
.dHPJ4@4,NSFWAJbQa[<&7W\XP297I]4(;6BF^H.b<Nc21S51f#c^L_(VG<gRP@#
?]<NA65E1NL9Xde:SWG5B\?&@(\?YX;?P\-&fb550dcf:99?Z@<6+PbM/CIO0H,F
ICH2WMCUAHZHf1KGA/;.GIBdLJN;U,9GU]aQM7:Qf=S#c@0S9d&d@BQSABZ8T3B^
FPCM+IZNUEe0;80NB@QWaON;c)g_5EH)Q=&9&Z?g/&&[,?E)AQ/,1BF61BUAPBDY
]&/KDPVD>4<JSP#PaaL.XX.5OUZ)4:NeAA<B/[/D&[&L.PO]]3U6+7UaJJ:Bg9:b
MCZF/Y24](WWC(9.G;3T),B9IQ_a2,6&Q:>1O-aeC[+^T>P<-76FeJg&(c\2@76+
O1-G#gE;ZEK:>?;NeSYXLH;]Y]IB?[_Y:V2;]/?CI-UM6e^XcVg,,<,_)N/_;C/(
,4B:^&_3cJ-=NN>Y.1I)&H8S-cBND3M-SY2PBFIWggQP]1=<H=G0)f^7RD<:+WK(
d<@7_2=Eb=W.d1H#e2?2.e(NE-eDSRQ#6H4J]Q>3A?<:#@LI\5-CN_a#Yff(=I1E
3U+2Wb.6]8X1f7EE9][[LMTAC[a2aT9H6#H?ST>+#SFD/FE,P[=.:,Y1,=P,TBA7
=Vb_?GZbdXGR2ZCV;f43;c4BFEX@T,>+CSgPaJDgQB8_.U)S_U=9W[UFUUC69[[J
:g4:YIGP^]WW/[c07+?W;<a(dWE[BM2ZB0YKD=<I)@Bd&I+>DTDEJDEPZ.:Q/S7Z
PB^_G;deL3[2c-2BIN+N)F1,.@FaL7O_/Y9=5H:2=P1S:^C.#a]HDRBAW08>cG.<
K\E??S=#3ZAH>eF>]2TNN;e7<V]ZLF9K#>\/I5C&fN#DcG0550/[ZCD124-^e@S&
#)1Y^(UQQ^K)&_\H??F[MW)ZAf>LC])PC/I^2YW?S-3_&Pg?)3O?=S73.2<U#dV@
VA\Ue75Q-7;<X)-7Kg9;662H)E,\Ea>Se,1RG4VL9OZVdH^TJ6Cd8eSI+Fc8A_3P
+0427PUE<=(5b:NDE6S_dQS/7Ma.1]bZfI:UC<W.F<^KaXY2,]J+)82^95_+HW,H
J7Qd95NRAZ<VF7S+&JX]XXUT^\V.W=(Ea-CRea9S:I];#4;JM<b[;d5bZc6)3M6U
_g[&+0#8IL_e:eN=2^.=UIYFTU+(^Na,2[R]78eVABK+2N+J+<<K2Y-)JbJ]LTc8
23/A<S\@QV>Cb2;_T4Z^1Z:W:,JNZCgM7G>e#@?RP_NI5W:FP3WAN1cVHV?WV/g&
@5C)/EA<GX<IMXL8M])I8-DIGW=Vc[HRgRPd+CK88,gVCN_LH?T)dI^>4Y/f]-19
U&FE^X6Ic[IB;aDYQSPT[H/6N?401#[V69a[;WgZHQg:4V6].=<?/.+P@OIX,#\M
/4\Q/SHUTe.WR7H6W<c420XU6f];Q^+D==?,aLf[Xg]accJ3GOP_(&feXV)42W]4
?Y.e^c/O#[+1>V8Ga5QDg.7-H)+I<?RALS.&aLE#FRCC.@PF_deMe^]D(+:2<fH6
-+]U,YXJWB<19N,cDZ0=&JE/^2a:X./T0GWHHHEI53\W527E0[L#9L:.X(/OD97M
6IV5\;:;C,<7/[0&7F6.7:5B49W<H&3NDW^A7.OLU9B[DTJV<_O>fTTKd:5W#:<R
.F]+Y1V9X7#^IUPd<OG;02NH:C03AA64W0Wbc&<OD(RC^IW(GV8Ra4852g8?V;^?
K/ZLJ>V0\EBT.YI/-WNfGJ&RN^E1BU3@6H-.B<U;3Y=(S8WAVg)HJAdV1#7_\?N/
/aQJW2;EFP_)TPUMfP4<)QCEPV+.Q_@TOW7EUQT4#T1K?(Qa6<6_,JWHT-+f(R<=
,N6X/bb:+@Pd25P0E33]7.HW7DVLG;R80()g/EP249MB2>BB]W457M7(ZR]P4d=7
7,,)L5V((LM&f5b92cS>=eEaQ^49QR#a8d)AW_JL1ZJG[,O(E4>E5GHZNgERM@DN
[^/D8PgVUEe.gQD>\4UMB)<0IVC/+_2\(@a:J^Eag3G2CNAQAY8gg.Z7U&e@F4ST
eL2/SdX,\)RaME#P@.N24Y4+&eW>IY_C#_YEFEMP66KgSASa3W8OAWY]9_e\DF+<
0>/L.f^/(9I;&3J<[gacaQ+SPD]637?-##7QC;,AdF47Z-RK:bgg)O_f[6OET9,8
2R+W7>PNZ,O9aF<bFWJPX/E4/)Q&0][_8Y8T99V0WBE+?LM=[15?V/3.EHXKTM+A
)W73dg;B/>:E40Y^=+4S?LH#?8EI#-fM/+2G5SgT^IV;I]O_XTX#&IMY=:[CZE0&
3\,5-R.4^B)b;gFe?99:AX^.aI1NaZ9HX[&AI+KD\]g4_CA-@g([BIa2?IACU7RF
C0GF)8S>N(624V2ZWfe;e_D;Y7EDR8D)1T\b3IcYP#_Td9W@/H.5L9R_4PDS_4-(
[Xe>?L(\ZTRg&<2]Q,^4K#Sa6:YT)bVUI[JCYO19d4+_/MP>XC\?W?]@70T3ePTV
GLZ-0??\EM?7V?>L6RQPILfDZ8)BeZUO362Ned0g=2M?+^F1GcAcdR63aQ0MaJNJ
1bX#CGDJ_UT+?.^MJT2??FbLRO+5Q,bbdD=U)Rf0>4aZY7Pa:8K)-0C3gD,@RdNX
)5dEKUH\:(\&I:YY@fDV8NILE;I[T?1]/YCSJ;,FXUc66Q7+>5\;dJ9G97\VCX3B
4FA\T2:6/IbXa2;g/b9Y7;];O@&^6<467PP9+N;H..X1Z#a.,Ng)b;7-=BH28eGQ
@E((CFWc6cF3:W7(_W)8)cc-W_XUab1.gc6^cVH7E+G2a5;V+eDM.ZZR<T2-?/_3
?KL<0P8TL:C=(dC.RTe4_c2:<71D0J3)+?aLe__1:45,RW]c;SD=3C<--J/A-&6K
D8,_aN12,)4]JA>M&;F@:>-(8ED6GB1Q0egI@L@Bb3eOWc)NVM[S4E0H)I&e?8-a
ad5&C\T=T;3>+L;P>?[<(8LZ8E95g&a&\2P)NIMUfaU[9-(K26de8WbP]8d.8L>9
AY::_[R7&-BRab=cS36g]C6<S]4B#@KI;bZG&O0gfK04VSL;NYS=N5VWHD--U^?5
B#9-_[32E=;c+W:g6FBVPUN.<5c;AH>.?B5@Xe5.526UN/:ML/U_:O(g7>Y.ff=J
;dL4g5D4(DJZS0f/]G#.VKB4e>YO(5d/&GeS2g2Z\>VQW.4K?Sc?1[L(8JE)\g@V
FDNWeC4@\3MF:<W@C2g:<c<7OE1TE&_;L;NHe?4RCW^&<7EK5a5SR.TaMc4g_1,;
\e6EV.L7=6Z,5D,VdY_9_=A(U(#YSV&?e\P\eAY-N:_[cV\=KVA^2/P0NOgQ(K&?
X6/87TQ:7KOA?NDE<Z2H^0P8>Q,TG,d_V[_(=RePO#\8G3;cV2+bZLG7f0U7&@(:
f7=C1N,g8\G=._NgC=,XLW_/QT=N\D.5UR+-P,C)RbfAJ[Z4f,3Y1)@]JH[A@JZ>
(JSdW2eb18P>0_L5S&EYa]aT(@WA9AE4@C481.V52CdRQ90&C]bXFO:\1E[MEA8b
D_&(H.7^&7Ia/GH2VTN//6Y?<>45G_9A\YGW2P:&-^XUd+Odc3\c-CEeJgQMTMgU
Y&IK=,@BA<&gT9XM03DR\=C/<Q35]1ESC50?gZ);Vb]@#?^=cfGN7M#E/a/45be,
P6f)TLY:[LZO)0=2X@[(863VNa1WL2=WJ,NNN?>A7EZg-c:E/@I\W0>R.9DJHV#)
C4D6ER#Vc32_;R_3ZfI>Bd@-;IPZLX0DR>e0Fd^S#eJP?0E6/+9DU6X47-GQF)HA
UN[dGC>98g&ULF1@UN,;O,N.S7OT046NT7;-,G;<[HH.((YUfHV:HDP)WH#DK,QW
8YeB20e(TeU+-bP>0.dV\ScEc1N23Z4Z^DbK1B1BKF&_:;9[[(+]JZ91CbZW]bb2
TEHCND-GgJY#ST4<\0TI:@4--83H=?fDVAE63/@MS\PY@-<ageHGfROOV5=Q[5_G
2<9BPQf4C:Gb2@O<L\4:9JL=6B0>4WH7^N)b\,]#,7aF#+LV&ZG5(\DDND.I[Y?)
T.A6c&,QX^VVeMOT;=6XONbT3+P?O\Ng(QK)b.B\4AV9QF/&ePf8TUSM=27Q/1Z@
_cX:I&NW[>?=Aa.X:Bf.g4df\\SC.>[e3gg6P1)Y9U=eNG()F-C54Y?NbRZ(959P
cG6_TOTdV30dH>#K2@.0+9BCH6=65[A/1aI=/Y01YWZH@Ib]]-..BXO;1>SGTQ^b
M0^]V,fVL0U+?ZU=7UQ,9&be>1-1[F7B@46</&-_XUCDAaU_66(Ca1-)V:BQ)5eA
ITTIfa9-#C_P?d0(K)EVcN\C=4#N[#.e<@E-@.RN.-M3N/B,ARB3@JdI\,Q#N>d7
;S.X@2S;-IdZ-LF=eHX>F1dK^?\JO;/H@QP=A?;=I:S5?<<9_EP848H@PXP8C3:=
@g3B>:1=d4D_T986C41;;>XJ>7PZU5M]RH(]bgd/L-5FHU28Q>gA4VPJI9+IVeDf
54gU5)bC]c>#c/E2LLOObP78KUb+<Cf7:#V>/X&]?44[;f#dBU.6&3Z/(HdbK4I)
Y8L]]>^1CK=DO9fWd&D9YR?9UUZM#-(EF3+V5ge0eN(Z6[+O0_AX-W9,a9G#_N9(
A?@=YM;Ld80NE#(-P#I.GUSFSJ?5K+RK][HfWIg,;a1dF;GTE/679KN+2:)T]C2_
:7=I83LE;&@HN8@)J,,0#4HXVg(/TB.+>7D;,]XgIPeefUbTE<=AMP)D?-W<dE2]
XG_M+f_c7W?MKGL?,Z=5fD9ZR]231faVG3[69KBHbU2WESB27L,,bWMO#H3ggQPQ
<ONLR[^GCfC,BK77g(.XO9^0X(H<g</M2VUBCO#,?WTHabCb+OMK8;8\),Qd\TX7
_^.1RF;&JY]ST]Q0UJ>NW094O69(eJ)Qd0ZbQ9C@KB8ZPFYY)GF[,T+>&WK9H2>L
VM??3b&J/gXXG^1S,aZC_((ZEQ/RfB3_^a9,QUG\?QAL9g.&Ec2=0AN.-51EPg8>
Vf&)6Qbf\#Ga7#)/YH7Ea+2X0R&.2AMHYS#CK1g#D0I/H]1Q/gNC0ALCB];8OK/D
e@ZJ+\d@bAe3XFU/2H<4Y)cG,4R#D579aN9;=3U;bU2Hc:HRfb9H5)^gHS\G,.(:
f=TGT2@>5]e@DJ95-D+Z/Q(aR0NRTN]F3d)I+dM9]F1&:gMKG[RQ<A]?@-?2#+0H
4X;@:.e3.,5RaXEOdZJ]E#QSd?LFH]ARLW;CX3B-]VeXfF+dKH:ac0>a9].VcKD1
IU:IN2IO4RNM-:E4e&=PE[gB.P.W2;8=6\ACI1XSg#C7AE\-fDPFdLZcNDRO.&Q+
:=W+/6#7fQ;=d3Z@KR>R&_^2(g7]?DA\e,N^R@J:-J#dd>6?B46Y/-BWJ:/_K+Eg
PI^4>>>E]9bZSN&B;)YI>(&67.(1XS/ba[LBIAg9Y73NJWFVQ^70R^G?NTLbZL>+
HG[Gb+0Q0@/&:.6#0KE69e&f3[\^dSMZ+_[/1J/0Tf2Y/c6H7;@.Cb2N6]dX3cOT
05JH+HYb8Pa@L2/ZN#RQK=M)DG?\]5dPXcLa#[R.:0J(aJCT/SA)_7DN&/)NAXMe
]cBQLZ1.TQ,Y16X4b^eC6RNH]PH9P>=9).&2K9GOF@=KR;Eg0RIGeSIKb>#;&Q@?
I<]^KH)@^JKOd6F<fV=.5XdY<.5P-f^Y:1;^dDOe618P6B_OD#aB(N)cBJ8aYLIV
I>DV7Xc,W0:PEV\4KHZdB<c<1c<U4M+)XY/+Qc@;&,F[&@d<+=KBHeA/G=TS;)<I
ADLE&<A4/NCLM76)I0L_S-b]UCZPg3XO)R<2>T:8SA)A]U.JXY^_(e8<DM58+fa=
0cM)JT7JF\J>.^2QPdL>U+3TIGe13G8S^AWFJ9YYAbX:IJ?2^6ECO,N:b4BZ5eLU
DbA<D/C7V6NS0f4+8;>:;Sg\EfP0N@0[W8K>Ud[@@LW^BG.:P<)IKL18\eO+B:XH
5^PL.c<0JGQd3aL5+A-#6V_d@aG]Af6J[PbR3Yc.@/cH5L=]fR;;SJ3f@57Gfb<Z
K[1XC^F\7@1T]>:L5OLC?]fMB-ebQ.[a5\3P@[eWHe;)&d_&f#A0M<)Lc4gH:P+f
Ya>(g:(IC)\d1]\Ee4Sc\?gAf=D2a&P(OTMKQJe//b[<Qg@eeM5VUA>(ZZF3Nf_Q
(#=g309ZI)-DI3W)O[^P0-HAW=0IWS_,Y0;AYg-U^7Z,A;gZY[a]]cP#WJ:&LMd5
c#?VUWgXf):9DIgIU3?>&?ZB:=[,2Ma/L/[?BDVP6AX^4=^U9Iba;D>L6+\X>,UW
Ta5A1fD8cBJU2G2-[eR:M\J-N>Q9W.FHc_A_T+#8S3F0FI85g&>:VIRSCN+Z]U\6
0eR/HA8HE<:BT:fCL-=AF21,17I#,cRB1ef9-0DK?EW_<a8&^J(U5?]&G+#V6H?e
g,5\U/a5^//>b.USZ0T#]JR[3B]-a>2;24:7-4EDGH3cgEaaM]JR01EW+CYKW]ZJ
+<87CdF\ON(].R)=>A56_YI?U:VYK\=C1M#AcF,b=A[b.fA;3F.<D]7INe9Q\;P=
XIQ_O;?-WHWS0WWcYX&.MZW1G,c6_720:P#OJd2I^AZf6c)CJP4]CIMZ62X(?NVK
+RR[)ZaL8&eOaSA9P<:]OA:^_d4;e,HJ:]F9N+D=>Sb_DN10fd&-T@F36]XNC\CG
:Yg(Q]S[WA[5g4Q,7,)=BT-62@@(9SGIM>g)1-E2];:;e&]VF7W::?4Z;/:;5=#M
0SV12M?U/>JTQL2:/Re+E2G@XR)BV:U/I)X.R]32a5[KR+CE5K]]R3:FGFJgBYZ9
WCf#ATfb-=D25+4(W+<IC_9A,QTII-Qd1#Za[BEX94<Og^TJFK]A&;WF&BJ]IEBV
cO1LE8WH>4E?R60,f>1W7Y5A:cY.72OI@(U,KY?)g6CA]G]cDEBJ?[2@08JY06AL
Tb,gF/4/,WE)2YAg+B3e>/0^gQ<SdBMPC17:?<5a(7:1Rb-<e[=9L?5XUgfDPaG)
Zd^T\@a9WK\4=bYIcFQG=4aQD)QS@?,[]7OKK395C)[-I\71?SC8\gg?SbTA&O<E
X79_;IA4-+(YGL4\>e-4^[J\_7:g9)RL2[]/2,@<b/R)(\YR^WOd=)OgY\6.4V+?
],Z,#[R=O.0.VNc4L#?GJ3g&,(=Bfc1[=_;U5=gO/&&C3IZ_->AK78D>9<?]R+<X
8\^G4=Q:.V[U#M/2;&X9GHb8\3=Y03Y0OBB<PH=HEQ8dI9M(5]PK&UR_cCc=f0bO
FLfJ:>2E.g.d-fT=B37RdT^^Eg4NU3d7@A^[)<LH.ZY4:1R-g?-54\45L(^5QHAU
c#QbaZ6Eg.W+LPS8N#/WE9cYdENa]R)&K>OVMF[)TWZ)=cI\(3Vg[)DBEAfKH)IX
BOGR#IL)bR[7Xe:E,VCfAEbg7IC@8c>+Y>FXGa(?ScSUJ(=ZN/G1D)#)@6MOL)\b
),\RA(7-gbWcFWTH+\9?M:U/bUAP(1.Z4\I-1/WcN_A[I=ULSWK@+1>3?=[E?845
eMG]bHcRR/2:+YC46cKG90aN]:e,Pc]ORL_;f<U&R49<JEL&+Ge;0:JgF#WOZT/9
QM?TBaNM6bI.R]L<F?B)O,TOHPF,/0B]J>dJfeNF_c]Kb2N05;^fVa1[L[N->;Bb
3\AA>Fg-fG#87[+6GP?7@ZKVZL0X[=cNH6X5D&Wge@E5Kg7/0UQGOd_HYKe[IJLM
1P(+=BQa2N?>)8fPd6V_0X.JBEbTQPe2/Z]gg7:,b_]4[WK5AU.WHQ:7#RDQPT^<
aU7W5>aP>RJ=Y#VV&SaHcCB\)VBa@)5\ULSK=\<./UIZ;(F4LEc)[IeE>E^AX>=/
J26(-;I:^Y@1e76R2J?KC9O]GL/RMOKI7@CffIO,g#/D(C8]K;aV]IDe,1[X<\L0
W13@J]S\LO<Fg?I3e/\Z\W>5C>VC^baUIOSFOAKIS+8X5\JHa2NA[g[YS3.YFNKZ
^O1)GJ,+1AaDaX2Bd&Vg[OB_IO\WcFA\4R=Y:K&bW+A=O@^/OV^C?EYRDG-X&V24
;XfU[ND&c9+AbcbOEM/>?P07-DV[]I&eECFYR=TM[(IRB>5,\RC1MDBS^C9gFM/Z
A2H0DRD<&V^D;\fY)FAS#W\dFCg>/I6Q)aEf@K>=7P-ZAV09COEd>>2BZS#GAL<_
bd_IKaD7KDF3Tf<F/F&:QW>STf(dV_N[B^47,LYV9@fX6Cb(M>,3TdU;FWI:CM;E
?(KJPQ2<;:MeYI]I?af#NL,JLI]ZP3K,E./GD1Z_&SL(II7>eKQK:63&09X1]7VA
9ef,3)NYMH&>B)PM/16[5beNFCWX)W9(4]56#N?]Y+U<I8@UPMb_\>^C.:a/EUQI
OPbgM4V@0I4b<F([23\=N@f5.8[#a(T\(LHcF,VUb3P?T^UC]4>:<1>>81UQAM0I
8c<R37IJ(]b94SF_GNDGbP#P0cZ@&aK^T;>?5>dg.[)8+bL>DN5;_X:[cg3JS:8?
c,KZ^)9#)dPb[0?X@c:)[]g#B.YLA0=e8^X5cLA.86K_/_0)ePX>)>+a\6^I25WD
#,a7X&7G6eY+)O2NI5-0(+[Q7PULEFVH;2J^O\G\MLc@7)N=V#GY4E?g8O._4Z]b
8BF[T^HJ_GP9#/)6ZC_?SBW,KI:[GU+@9J@?f@+=b>c[PDfQ^)KGF85f:V:/G^42
f4Bf0D)]aWgXDS52\I8PE;]A[PDQP>.4bVX3a[)Z<\.C1?=TVfD.[0S7c6I[fY(Y
:f9#,G6W^,VJ;9-7E@e>UAb1P,,cDE1=cdL[1&<^X9gI]R;KJd6<_M_+2KZT]\d\
[=[LK)YX\,ZL:R4(FVRW/).778/SOgU^JV.MVT+@]\FaO.720])5A(SD_g#2-_+a
IKaBMYg?,E?bHH>VD)Ef<XE3T?J^EVEZJ(@3-cP<VCa7Q-=3)=YNM>(BKSO=#8HR
dcE\?MT]c5)#2IH;0WNL+=VM1A&a\04d+,PH;=cf>7I[?dJADPc]A2QKf166d@Uc
c>VggCR7,E,MHWTTE3IPc(@0\.g-T6V0:EZF1Ece&f[#W^<(CBM^^[>aC=6Z/E?-
a4?7RKRE;J]GS(b6aa0FaNUV?S)E>BY<g/C5GDT=,&)D>^&,e,=S2G0+QFL:U@DS
6c#:cN&26IWWBeAegNP29>.)^Xa+,^#(6EJXL2gd:Te2)AB<7cgAY6YXPCUO/J(Q
e5SIR0#3FbZYM763#=IYOJ4DfJ-Z@P]((d0)eKTH4&U0cO[@N.H-5^WC]7,<fF<-
#QY\.3.4W,?L(7UeU]0+,5DV7CL]8)<?2Zb5X,baG#^/&=^GJU98eOC4X.?ODTa_
W=TDLV+RG71e3+1\\G5.\CVbfK]7gD@-)@fBTcA[L33DX4Y.afWNYO=I3Y7^O>H@
KLdKa_H7L?X,D]4Z\f05ZX&dH8/Wc13gL0?+V0HJDXGD;3V4Q^d#YNW&MaAF.BTd
AO/R?5C=S<:(+#Q2)X<EON8=Z4(.^\8;FC(<>],?ACE=_+D9SB8Pc_ZVg>Ug/6N7
CHZDGegbB@[AaQ0&-93>[JeJO3T565HWbCCfDDI77DX@G3]6c:,d1b+G.;NC@49N
CNNI\a5#.F,^?N>f)bMLf4Gc&bPR=fG]Oa[5ceW#P.G[ON/WO_<eX/deEL_YTYC1
cA[T1_aQc83Q2MN[]^g]Fba9F)#U7FL/(4)_c;38OZY&>.E5,E(4a14E\XQM4-L?
KbVbMMMHNZG?5YM@#5@SCP\?-5L;e56W8?eSW8>GXgN\87#SJN>&_4X1WI;[W##?
f,=0]]00KTJb)EV:_W)@Vd0dN^3G8(^be[0_S4HH]VNgg,d\BAW8>c;YaOS4RW;A
&&dBb3D+adD3[0b/Q0g#8c5e61DJ</A<1&ZMBTT::RX.@=-2\5ZVJaJXZHFM])fJ
e_&<5(&JX23II2_M?:bMM4&G#R)9fJ4e8(<#:L#-8[]W?-\RF0S5^AMX\4;0.cFU
=R_f0]3E#+S&(SURVEb?02_,f-P,>+8><E,aIW]I8MT/MJA\[3(]Z,2?MD+A:F&/
8YIbAfL7_C&-B^,&6K7)=fP:a=-N#LBJH^9_RR4JI)IcD8M3#;0-@eFF&R:I)9a:
7)Z97&I6\4YG-8664^fQKe<b+1U5-\Lg:F=DJ+aPBUe08[b:01IDKgAXQb>Z&:9+
:V9+F>ELf=WJ02A^@A(4Y.:SF1,9PH;4;W&\0_QcC7H83/4.\>\=:K].IVc(NU7e
ec6-:M6BC=8#-U67MO^Y1.^-P]NeBBYR7+.:E1H15C6_K;<ENAJ6,]45>d(SYP0L
4P[4@G5J9J=9^]TL9_aT/]W]5e)9U5GE1LbC<[\N5(4-6#\0OJ&+A:)ALY7ed;;[
WMMVV:\9D=]S5HND:YC4V?ITE1@b2VS.PM>eeB-=TNeSH)O^Bc&@C)dLaOD3H7IK
L\T2A&T8(9]Ze:)M;^8^Z#V+eE2O1I)BAgG[U2&I5eE0&\#a?Q[gAJH6_(e;U71c
E726_-E&FB-NDRa_]3b^cZ>VMEQ;ZS0=R<V54<.c^NIHR.]\T/c3S4B((R(c]&/I
@Bb8SHgeaO5IfB3]MKSP-6\AX=85e3L.&C&7Y9_C)C@,R#Cfcf=Aa,Q\CeDVc^,a
a2TZ_KX,[XG)d]WPV+TK<gacUIF1OY.fXbXAV.EEF21_6#e3c(WFIP7KR3=V_WE(
FXU8bVS0/_d?JO3d<Y8EA<1\^G_ZZ.P11gN-,;4Hc@N&_cJI&BA6YbF7I#PO#CL>
AT.)@W>IbO6/U3>9>/2&:G1N=[=/J8]M,EC-MKH-.(?a0VNS]Z3L93;55NQYI>P0
/A=5^1N4];>50OKG5@GATDQAReQ:1-:NS?3MX8QGPV4IRDeOVIDW8T)IdD.9A3C+
L?0T@FSYY[Eb2F3O4CB+OMRL75HGZ)Gc-=X#?#UR@ML3,IWHQ^WB1;\^40-dZ=1D
)DNSNFEF::4-V.K&JZBV1X.?;P:(IQK#fPN[a4O&fC6,K\S;&D]&FY/SW8]LgR4a
#A:>Q+M(.FS&1U&:cO&XNb(R^Q7^SL[AW):8U#f0_c(N+d=;SdDIcXg(O=\/[dM&
R@8(78.fATOV5P)NQ.ZK?892E9TU8-S1a0:Gc>6P_?=gU-e7SaA6[RNI--D<1T@/
8/1aX34]TeHCSA@6f8RR@:?d4SJG3e-Bb]WJ2VHNH7?N4KOAT5@6FX77W.KHKTJ)
f\ce@EG=;M.5V<eWJLZ/-=A<+Y+fg3;]O]RM&6<YfJ>W<9I<?_Ig63JA;U\VK2/6
<G+3#,c]>&(fW5]1>#aWO@64?IW3DU8FaYU7Z^Dg94I./TCY9#W\9<GMFJ\>6IL;
)PN.=V7c]38<(<F4R]X)D:A&@M7D;@=AT&O-YZX>.>;Wb8IX2GL.(bI[XIBeOE:O
FX^(YTT7B#-KHR3<2e@FLJJN:K:UA_U)[E,7a.W\.Q_0PN0L?LV/geN7<OObU^5(
9&:4^GZ7Sf-;NJ^(_51_1Q=g[cSDc]W:V(f3SaTM:03ILT1>B\XFK)Ae-T7C0>N:
M[D#2GCA-AMQK7Vc6_=TROL6YL,B&R\fH.b5dSTf+><G.JOE+b5.D4-[:V2_77bX
K[&I^TVdS0D[f.Be9Vg)(8.NaS\.P42#MHU_1,.YD)c6[N1CQI\FbU:fTI=PKR&d
+8a.:16WF.FW-7?CI8.:A&UEVJ>_-Y&A&E8a(0g9fPQ]=Wb(D^4PPYA(-;@b1BLJ
8]H.(0SAU4XY=2Dg/AEe,@JGGNYc80]Y68-+<QHNYD&b]Na]2(F-gRK:H)]<VB#K
->Pa<2ZTY=@D+e6Pg<eC2NRG+P[OWUgSO?[&Q_fNZF=#O]NLXG,4AP]f9@;&58C8
-()cZTP3=.6b9^Z\[NMf-K:BC/5OX,&X0Pb6e^Ng?O>R5,cgQIZ1LE<d+Y9.TPcB
:cBU6=HF,\N2dC-,bc<V58[AS+&)DQLTOBZ=\Zd(=2Z2&R]]],C&=aD834c0UX1J
[@=NEc,QZ?1[-Se8A5REF522WZ5O6;<,5X]AeS19GE:g526K>_NLg\1e2#N?XO.V
XJEP:KM)10FaC,<#Na]GC5(7N3-J1>C<ZgbC-<aec=CDMBZR^gRGT4L=2;NF/?D2
.P&VPU)WFV^:8@U5)WQO+0=ZR8QU<[M#AWKUJ&FG)HXfaJSY0U=B\=Fb;f+CfQ58
0gfV0:>RAc/?aOa,5\_77_+eM(3F\)6:g\30]4?HM(>A+N4?Yf_/(DFCT^-8)[J;
().f/;9P0bYf8T/9(YG9DdC9P)6L15XLL(#J&/J:757b,DI]E]JXeT4;cIH-JC?F
C0\+#B>O1c2EW2DF1d9;ACDVg=ad]6b4)HUC/g&=W2gc>65R,.d+NEcM^KVeW_Nc
/0[JgF@>6O)/IB?1BV;R7=.0I/71@]Od&DedR7V+ZCcQ.b8I70)#Zd8Ec]RCfNOT
cPf6Yd@J/;)F#1S5eJ8OCL+X6ZZ?(2(g2JI^DD#\e.E>B(PY4[=b+(gf[=KE9])6
6#\@L;QDX_=F9I]OeCV:LBTEb2ECQ05]L?,E^B4B7QK0-/&MT<3;a_,D+SAeZEPC
KXdR\-O[Q2a>aSOO2J:C0:-_.MK4)BQ7XGPQ79gW\T4F0(C21Da6R,91?I]W\bSW
6)M&>5GcU(&VF.\A+R61BVM;/@+R44[T9GZ^FS57&FFNK1AKgAK_1B)QCO[PK:aE
fFA[,8P0+VDZ\73_Wc2;^IIEgD2G]aYKH)(^g6Z1=Kf_J?/)[.,OJ7PNAf0:/]>;
;2^7G].M6:&W;RS6Z-b8P<BT34#QCd_Sc?P5;QX<NQV#6\5d4,&RC4fQ6@SH-K-+
QP0^/aYY_1IfCVJRK&4Y,gXBC?@\7FO.4VUD6&HE?T2)GFZ^Q)1[GW]SgA(D-d[D
,&D36SGZZZcPV&)/>d?QH@1dKVO90-TNG<DHT6]:gQfN+9DK#d3A.-e#\^CLdP:#
2K>DJ\bbA,2CQ=87T</[Q3BPTNg/G>>d[P<cS63KSB@Pa(\;^1&E-<0d>=7WGB&#
2/)b.Ncaf^1#-JDC\gbI?H1]@C:HWOD)SQ/;6GR<XATNODQ2.6)SKGLJ_M2;5IRG
-0b-#;V,BgLFRDS5d84VEAP@Pb2Sf,)=f@,b6(I3<[@Ie:@JeA:TRUbU?dDOR9SO
LO##.#ORU+aUT8edURP1A>af1DPc1a7_g_,;SJ7H&b9a>X5DLId5J;,AT=N3gNb#
1PT:<f.Lb4IFG6V,3;WfE@.d\M<]L-6b:(5>\X-7;JFCKS-/W-M3M+fc9Z9He^0C
2V97,,F_+E@2+:Q8RCHOWB@YeH,]9BWB_RK_23&0f&a>BW15I[0adI;5V]fSgeFQ
UH6NQGPCL()WQ,.TTVBG/g^5]ae2Y321+_W@^;OT.L>dFOA@P2=]W-]Y+.#4IQM\
58YXdP#B;e@B.>+LT^YWVHU&O:B3=dPQ?2D;-bYXMDZ,(V?YN5<B:Q[Y=/DD+=@:
\7d+<IW@&-S5#KW-_DC7R]TSEOYHg&V,E2HG.W1Y;3H5^>M13B8H+f7IR>LSK^5[
MHJPbEX?CC-&<SZ43F_DR]LOa+L(977f@N=fJTV:CTBWE,g.:bT[DG[<,8Vg_)8f
2[TKJHPG<.,^/dHVa)DBaMdY8aJ8d[f<@[b6XT_K0_Ub^26E1].TeeO5ff0JFedF
5QOA-H/^GT6cg182=5IcB=cO#M4:7J<A,@c,eYXCQ\J7A)2fVdJ<.,W\0d53,//_
R=\\;2W?9^P&ET6>P+N0/0I^]6BQ4^=Z6Z^02@\UMI0Y/4@6900/:]JB5KXPC=UK
Y.Q5LQ1_50J\0JB,MR4b;<?,;E)9=2NQ9]/^?EeQD@Xg4MJG5#Ub(30:I#R=^9Z+
.@:fRae-<PZ#GM5?4WbTN/;f>)UQLD1/TV9+PHQ92K6:Zf4/U_T:g?AR>M17#M#A
U<AN1.STMK4fPKc7dfXff;7,9-<RfH)I.)POBSH8TI2f&A/3eZaBGOII[-bf+@fN
?6.dcBM_V@PUQH5O(48CRbL1X_g1O5,9^;I]bB,U(=M6OUcFT3eLWH<b4+G;[8f8
_4>/4.0+d+[+YM497R4/\P61UA:5)O\8I^LN^ZPI;fO2d1P3Z,8HMHT,&>d=IQ68
3>>UJL:T@4fO@:&_bW2/9MSM9A/N2Hb-F.+B)3X:N8[)NaY6X_K?)QPLH@8Q-HV\
+5f9MI?#5(d#EI>788N5MF[IL@&1I5EXF<5T36B5/Me/2NbL:Ed/7KA5aTbTGB[c
?8c+J86,AC].,PPfEBH/fXa0TKaHNMI2>PT9Y0=XUNcX@FNKHZC[N@[7MH[H&V<N
T)>0&RJ1ARVPYW_7BHQU&g#GOc=+(MTO+(Y.d6KfC\M4IVBDG1PK/L5AYg)=[VBM
#\]ZI.cILI5(3.6,BTSJ@J-B(2PF6NH@1Y8TYKF.[cVQa^ZMJAC7)RG&O0S@gd7b
O8,T?>A\H)a-UK/(f_KK6OBf7?;<E-J/;/1?S;.Q,b=V2c4=ZGU)UX6a^Z[KF(dE
/d+;VBe=KSZ6@1OHXIQ<;>GPB#P:&7Ea-4HPaKR0Q4)ZZ;Z[c#-XYP:4HIFb8>Lf
G<U16f7He4JR-I\Y)=f<X8.H;C3K/e&IPS].-K\=Q(G.fBf9[ESI,Kf<F_PPJAD0
>caGKfX.8PVfP)H79:1XA<(=Q;=RLJ+;Z&PIAV2A^X:=QfLR;VGKXOc8&8<X2INI
V>S4e&BS262W@QE8gPgJKOD?MaADIC;5RELC-L2FEF4>eU/O55-9WA.TL4->YW[&
7g98c@K&<B[Zd3IQa19V#BC\T^2YDKC\2-TGQ>cdg#IH,MJZ^dWVg(2MDG,7:9Z^
N[cbYGJ6HRR4g\b_e8SHV;OKVeRc:cdBH,=9LTL43-.B&/7^ARNf-]J]b5T\+X<-
6:>Q>I1@5_NP+2S&b1&><N[]6Wd/[/O6?JU@5I7YIaB>\KX>L3<WWY>f8;K0I91[
4K>gK>5)bMOH_)7TcN^^;@F;SeST,Aa.]Oad>CIG6Z@7()b_CVV1<gU/L0b09GDV
Q92B,fFXd7.5Y4E>+N]<8NOZ3=+O&T0+ZZ<.g(7@8Q[La1,G^e9Yb>_X@K_)W;?N
4]Od?SJZ-=/U_>;c-+JIPbY4c\ag/YXGBUg/b[3F-@7Xg]B0QY@UT.5A@=6(B6_V
7+(+P_,]^O]abL:>fZ?gOFHK]c0J0@3LA8;EFg]Q&DL^)Lb+]ae0P8J:?(#?Xb(B
U=dO:cF^Xd].Y4^8^WI<dCH-9:81,B+96[g)g[B.F=_=NT)5a&FJ6W:HN8:c)2AB
V([GH@O0K\3X-VTK_I3=W:_2P03&(17&^->3T4XR2<G[B]<SZ//))<a;:?2_eOAc
6?+G?,<fFAG/\O1K?38>eN8UYEU&EJdg9Y<=<4SM+B]NX>8eXFAfa.9@Q<=9.g?0
2?.L7,4P=CEbJ+3Q7CHL-S_4;ZI(Eg6+feCe=#S]7>[LI#7XQ?X(B^0;Of3beH+U
=(VK[K-I3@BOZf7?TE2.]Y&8aX[PZf41?gYXZ7SIYEQ->Z[K<@K0QI?L35Qdf.Rf
34I=,9T(N5#N_[]0GgbNSXWSe]6;LM7dJ^^+^0g?]<R4B,H^?;FWDQSF)bX_+?13
+];FF3>f?&Q-d4&A)XV(7@(O=R]\.@AH,0eL4;T2-2d_3C<1R?M6b<CFG6d,M)c:
_UHP#BP+<&3)eE3>S^_-4H9dG]J?TXY=\\XdgV8G6?E]8VB<YaC_KXB6YF\;,AUI
C>\1BJR;YR_I/V)aFgZc4=b/AU?A/&2bB-b-G^b.HXD,=RZTA4TJPANZ@R@:UQJN
a_@QS-^(W_>#[+0MF\H\:9:O[aD_MC0Y-ZIR4&5>&KQEPV9Ig)7U\PfTXCORY759
#]SCfaCUca;KGR^De,DH+WA/9OBBBJA2?M.QH0<g5J1N/.V[Wb-]W-XQ<3VbEg1g
AJ;a;V3XAG<A^cU=_aOWF#f\1WGPV0Y7^IRc>9Rg/?N6C31UHF#I6^cD:>@@LCW=
E4VOLQ(g2ML(8:Qf01Vb=L24T1g.A0</RNaDZLC=-b@J56+]\)5L2d8+FJedMY0\
@0EAS(/e+8a;&]5,FQVE[af8fWBdTI&&>Ia7:(&BdeA98^:N+-,4[Bg@X8Nd&L.g
Zg0P\)B>fcBMMZT)G9Z=G<(X<+KPYHT0EX[.\Na[]\CT9LI-F)J=(4-Q6S+-+2L(
247O1V/a@BY\CP&.I;30/1@g6TEP<N]&(7X9CQB^a64048d^T=:b>a8D]TGQa]PS
X4XO9V@>;1dPX.=5=6-<Y,c#46P2W])(.#__9,2YLK@gK5U:[gBU_I8)BRKG.H)-
[WEg\\Vf0M@Z=5O6_81:\XRQ4GgXFS04gc_NaZD&KOIc9bgVKd6^0PIg5/M/B&;S
fP^JA7R&.WVDbS,E4/]=+OR8;41TI,d&M@8Kdd-#_@af[WR_ZY;8c1C0E&?Gd\D]
53MaORYZO=bW&VL5BbBfa6]6C9U/<MG77TEE3DD@;PA?(f,F.0[^/<WILY,UbP^e
RINHY&;D@eB3HM[5F^8X]3178HB.0QYO8#0&3SB\dRB:7E8JJN/A#@&)B<a68;]7
8RZKKe?U^@UC^5[4WCQ&S;c:A/?LA,8&_ZH?KX\b(Y:1:_W>0HRc5G3#<4RI&+L0
Eb]UbWYb>C9Wb/>C/V3HBFC5N0Y8+I1fFU4@8)5G.)ATLYVVT69>S5O];9#C)E@B
JL6_c0dCSgV(4TF?I5eMRUA_K,53Z6cQJ<3:47X_<H<1gUCfYaD(E^795V2W#eY^
BO@NY\03/)Ta+B-()a3><b>9N(Y\dVN9HXK=FPB0H36164Z-YJ[H7VN&[_G.Y/+V
VMa>=EP=]:H9a/M@8[VKf3@AX?aWL:P3>JQGbF(Z:D:4U7>\AB7H/N@.H[&-]4-3
#^U)I6@9(/9EQ^0D92a<WdOV2;bO<bKG?/K&HK1GNR_d[(ED9+6PP,OcgM/<EZ-.
7T)0C_65,I]&ZSfDa=2<JMMae)<BK477H1CG&&<&PF9;GXdJ+FVdS7=QT/LaF9VP
KYJe5:X(Z.YcLJ@fO&O3<f&+RCS)S<3[,g\>/FgZYcYT75:).FVU+5(6MJBf4Y[&
\Q2327LX1A+->N78dcB0HCWBG[:45-];bfO\9>#Ab5HB()6#O<U@J-WJ&/?O>B:&
S86)^0Zc+dN&&#&:CbW+C(Q>>MVB2S#S5:1Zf]a]XOOHZ=E#:T.J_]?eM^N)X:K8
KHX;CL<L<W5RVZWLeH-:Q_\?;#Eb)f(;--1Z^ZQ=e\aM-c.UcVIL,cBH\SQ;C2Pe
L8S@58YbU(X@A>e/aTIE21.dIC[FS^^CbbNd[?MQP]H_QWfg+^9I>HY>?J0A2M0B
bJ5&]M>Cb7HaI.EKb:Y[77;:ZOV1dR-\dKY?)VRHDb9^L#9DbTgQO&bRcV?4\Cb#
4/O1/=HFR_H#c(RT>3V)60OC_5)NJd+T)e_50Z3P@G89AI2e@#EG_dH(M</T2g6c
6VC&F(LX14@IL4[I=ZO25.8cK@F_Q[2IRL>\.9N-O\:^+KO2^@&M?QD.;38I7U)G
5-OgeBc=2>[beTQE?G2A+,LX+VTXYP^g>QBRHGZ4,G5V+Eb)#6#ZY6)UL()VUEF-
ZU,/geXKdJ8/?.;9EAV95.)^-RT(EA_X4@=-daGZLCIA)3I37@4ffO7R#0FVDG(.
&?,2GHb_H^1M>](^TTFf@]KG7)8daUDC<g4Q;Y,eQb+N=EN>>CUa;C4EG:Y18=eF
,BeP8K_GedCCJ7aaPX>(@A)L]]MB7,XNA]7S#68a1HCDRZ++75,&7G3EJLHPGgL>
_R>,Z#fg,I.&L:P;29,6MAA<ED?S]aRdQPL#VHcT;#B_26GU8;?->S-JKaO/Ra02
a?GV?Ua61TaB88@Q-Q0&a<Kce&=^ffBC?U[C1A,R)V[9d==&1@7I_6Yd&^I;XHP\
Gb,(EBgT+7@O&<)?71dTIW^#<7JD7S=4A//0/UN<U_IMD92PL@RCJ\E27D.5V\e]
@]Wb+33O5#@GH6O2,+9<;Q/LO.:Ce23R?22&dd#4ZZE317WA6=3FM@Q<>:=?S&:P
):>4<H1C;6SO,e:TM&Fb_41IZSKQS):I3cOSD#KLVBFA)J<UWEO6LH&0JgE^HFa&
YCV:)AU,_K6@3-f-28ZSIZ?Y-Jg1K4E+fZKP3IL)<]^5+g^PE,WN]LXBD)\f/8NY
W;;GMb:3H_GVS9Mfg)FbI9Oa/@&T,/^8Y^VfXdgO0#C+]H>6\V+I>HNZGOS/QQY>
^:)T2VT+C2]JN=UQHFK.P)&_FF25F4[M7gQ[7I5/R&gK^\J/=9M8YTK@A6=&2@6L
O3G(Zd2HH;YfY6\),_6;Og1N0eI8TIYY-8#LcE3IEZ,dC1?@g&\;6=#IWW0:]/O+
S(RYe0_#eZ^Q932LS4@dDeQ-0+KOO>N;D,0Z1)Q3YQdM.3P#7Z;Q1RC<Z,(Jg6eY
bb++c.]W)>Oc>^622QL4AWI.c=;eJ&^/7PUBOCG+R)c19L[;R:K7.Q&a0XNB&CPA
_[bL@]B(5\.(-4EGdKB_bW<JN+RAAEI:fS+U4G9B<9Lf:QQT5#DB>b#[-#Z^=COF
X4HX85;JI_\Q74-b8YY@d=KG[3-JD;.O(B9f/a:<;XMW^-6C[V_\1]OIeD^K(e,J
L&0X<Ua6E/BEcfa08b/2WEF1XGQ)cK^NZ)2(>F\J9.RG8&;4V>A(>X>@c&ZXVN_X
V=HQ+29[(J,Qg5>.72U)KP0?RNVc;+..bBa-3R@f,AHL,[7RfF[AR(g8WTFg#dYL
<7S1Y?B;Jce[NY[=H,B_OaA3CKBPA>.-dZT-J5b9\ON;bNEB_0D_Z/;;L^(f16;a
Zb9GC>1CK.UdMMYMJ:57\3S>Zg,@[O&Y^Cg39Me?E_XW@:,5)U4?S]46L?Nf3P50
<7^5IS\-CeUC@LSZ3.OR2Wb3-HIM9LBHE7:5^_3HfVD>O+1J3;#>1dJY=X.=SE-9
baIE_E_c:0RV&A?bC=LT[F8;C^dG+GacD5cg4S\7A\;N&L-U(FNFBHT[>KLc3I_C
]IQ&bWH8+_C83_D=;IgLH==\V)7eZ?;-_ZEN6b0@4^;)XHNa8d2BF+.2-b8ZYF^K
E3#?#[L2?14KKD7QB^A<-<eX2P;3]/JTQOW&[@1VG,6Ed(U-B@I1T+@1_5J:CG.<
NJ-:Q8f5=_V5@_eIJPN_RR(g@<J@]L:Te7/F5NQL1LIS&fcT;5B1DCH/5fRG1++A
d?#B.3JD?)c=@b0AJ[L;267?#XRFD.D\:9=>BMTCNSV(1<B1g0&.Gb,==]006A>K
_L9Rc[aA>[<_dZd)1b[b:_FL-6Y]SCVF;@6]=d\.P]+I/9OW?@<)O0L;A;OBJWSP
G(PMJK:9IQRC;+MKXO96]W,;W/-\OdA,8:7E]G8_HF2EX4HR@E3<U;B?[YO0XWQ#
&:<aIBUg5R@\R/HRV4/a)f.(]PM3G)1-XH&LQR?Y]db,]fRPR;,C(DZA^@<\\Ve3
McD+]6-N&d]aSNO?1NM1U\W/AK&IdOE:)O+6U]<:DC&4MF[+EK(VAJS[?V2(:-7,
g6H^TF?LY40T)^XNE.15bK33:Y3W0[CFeJ&-7]<5adYfef1F361C_DJ11(FH2)DC
=GG-RFe-IJZa/W;H6+e1(0;K:#/(f],5NKgB#L/_:Gb?6WI#(O(I9YX:Z9\PCgY1
ag>K7B>2K=Pa8S:RUa/ee8NB(ZcNGEY&\^Z57OA+ZQYVVAU9.E8]Wf3\N0.[CQ/G
Q88aO.X4ZB>J^+7-H2Y-MS6>2ER,N9ZSAG#;GCJ-fWMb1g1;G=6O>T9cDfK1,SP]
0PY6R52C(9\:](#B8.@JIK,K\bPL#S8Y<3eJV6=G,+.DaE1-DU-8fcE3D>G3_R2R
Y.75(30cDN)BC1NMQZa/?J1_=FP?W/#MGK^&/b9.X6;(Ib><;\>?gG.U3F+IJL57
UQ^-VK,2JNCNQP)#?1N^QQc5cGS5T/@=->NLT@#dP]VMKZYfLHf)aX-\ef@aB^IK
5ZE\e]:JCY([-YYB[O.gfARY72YZ5>J\eFOJ5DIOfZ+.Da_V][@BU=M^ZE+[S4@M
JILg<@7X<S5,QG:CLZ2M^+.-^+cUaS9gM>:c]UHR#I0)V<<AC^4bCB:URHbV95@3
B3g1>@5KX?SAS@#86JH0WQb-EU96P@3X:V[C-9b:_A#>TGYU&5T++F+/2:IFH\71
1W6CKeP>BMY.FV:Z7[[)&PFO3MeI-eg1Se(>aMZ..C6\fUK6^^W68TJK;(:\9NN[
=+0bIW_;D??9XRF?B:)5LN^::FH_ce_dC?LI^EF@D6c#&M=W>>1Ja-(]DOd63e)-
EK&7gL93RN^DHEPM_;=P7,,D03b\,b,S(XIJ8/Y?0W5eg9d<^1cJGOAXG#eZ@\E^
JCaQ&J.Kd(T/1.RO2THR59PXEdf(QZZ;<22;AU/MU?/=:H^O.(Y6F=O1AfFW]SS7
>U_deg><S;db\\>ZD#Ia=C8Kf1C1=X#L)M4/eBFcD#Cb8&ec2B6FQ(_dHU>a<<OJ
:,U<Y7)SVJA.7YYIC+G:)?GNPG=/EVfF3a_5dcXQ&>(,&N;;g9-,VBg^D;Ke642>
R[#6BK<f#53SUdX=@+U5T+).I>4e<T[2ad[c[50#;)GJA(beK.2+#N_D]V:V[]2K
OC&YE@^<WIH:+:>:XJC;5KQ7^MBV8@bB0ZFD^&ZZV1R5.(R,5-X^6&b_0;N#IW&L
LO<EP)A:0-UY=deJa85O8P7f\F[0N5T?J5:L7RQST+S5109\L^80\E^HJ,eLGSOg
?Tf;HVcX9:PNYdf\2d9[dB&+N=^RO4YfVH-cb/afc=HdO_\]<^1g#<E]ONQ,#gc-
0,)MIUdKI\.AA=bC]S0F:PVg12]eEc>8.&NMAfY5W.5\SF_4b;/\?(5<8[QZ?J]+
@+@5gd29V0/8,;9Z;(UNQMK?7EJZ7#U\aK<g+1>Z>9eB&=BTKc1)Yg[Ve&Tb#R/(
EOD2\LDS3@REeI7TcHcNdYHb15S;<K#d0L8&7:f<gN:OMW15RgL:W_8W.M.:3KdB
:K+b3FeK\5<I6AQ]K&@)-CdPYfQ&g(06)ZOH<:PEaPI>ZbcfeWJ2B>+M@g-(.O(N
+8Y3#X-1db=aPK:EgAZBH/U.@RNe=,[+P8,Le6#JO/.C3[K_.36e=Cc@\deb&UcW
ae[O4PFR^dO1T&fEF@WX0]+dgN5UZe+@DTgAS_=E;:dN(c()425YQPVHDT]N^b]J
>#[dXA[f?&A_7;c,AB,g.U7JgJ4^fO,[_X6?)9ELMG\([@22DfDSDCV)Z_YPZ9UF
-\I>8G00NPDfa)Ee3a6M2K^0&=W(KKV9E14J2L:<)_^\db,8P/ACYWS[,a8T2Q<#
)#3\dQ=YV==B(1U@,S_bWZE)45AdL?8Y3[U1I(a&FHE74][/X3&.e0Ogb^.:+N7d
@O8A2[b<GNcfENd<a=><])Wb9?cV;2V+Y^[Wd:>-<Q1E@UR#L_3&ca9>S6T,,>=?
&W@V?ZM\0M?-QYD_NR)=E.N-5#D=&&._J]X2[C1:0]1bEJg0VOB1(VW\7;=\9Sa:
TH-2@/4-:)c3247KdaH<c@1BI/RMKL[#bA#O,@1Q<&E(&-ZgAHd9I\fV;d]BZY9X
D3aB;,W1TJ?R6O;NdCcg;.V?+KULWE&gJIa.F<?ZG=(0[RQ22,JQf32M#Q+]:Pa;
S]6e)Y;>H#]SXaeb;@[#G.\dAJ[dURL[-Y14X0D=U3J;F1T.]UE3@7G\&?.M@SXe
].<B;7MHd-P\O-^T8M))\2E?Cc+66D<RK.1-I4@S7C2TL@40]:.DSLNHLcW2/A<e
/_,#LD6:QU3+VESY6aa]=bB9MW/a3?,a)Q=;#81@_1^<9DU]Q^.=W)?IM#0f><WS
g(_>U7QT?eF>c0HWHd0Z3/_P^5MWZ39)fNe2^T==eJBZ7)FJ35Pb^#X:.&:/8[bc
-Nc0e4V^6MF3[Z[J.b7YS</K@]9DOD+-^RcBG>XMb6D4M\4S/BJbHRDVdI>R0F:d
\W7gKUY(95f:C<_^IGdd#@aISN_[.IQV^J-+:MNMF3+#gRI4^1OV\\#OY\X__be#
gb6=0V-)2=-Fd9c8I0\Bb]YYY,W/;=gNDLAP#(BQ8e>PbOO;:f4A[,4dD;WZ9C]Z
4[OHN)82.E1ER)NBB-P,Q:6Y4BTYBJ0bUH/9YfVN@#4fd0FZW06^a&dfN&A3?SQ4
@]:acDD5HP0S?[fE2DRFV/H6C2XOa:?8,CKd17QK4Dfg]<D0=(bFRe7RK@N[:43A
^fJ^cd8)XU]-<B?XXD(MAO(gR\+O60S7=ScS0REA>(;d9AJb4B2bcR,YfeJNE\:_
9GP,X<&/02BHAFMD9C;1LMWCdgdfaUNM4Q8QPMO#SIJFO=-G1(PEMLZA#6K9,Z^g
PZQgI;Z[S1=C/K(V2ZVd<JUW/IJfcf1c<<&F:.ZDACAGW911_Mca0F(&B\IPQ+CZ
7PgPB:cH?2[)CfGL<E_bS5(NV.<Y<XP(QYC;K_bVL1Z6(RdeF\b/cGAPXZ0.M,g7
Ta]@>N(]9KR]:,=9Ta#^#Ig]=Mbd.:eI&b>eIS8=?&PB(f-XM[CMF)2N0GaWgI2O
G5)S(,3]\#>_ef<-fC7GgJg-UJ/#XLffT?(O?>aI>I]#L(9_;4c5E4/G_N->GeOG
IH8U:\H87a=.C2^Y+)UXP=e49V)XO<X^?X2/@c?O[;H]Y4B9CFD#@dSgLA[FL(fT
6VM2^P,]9b=c4?]>PX?>O@?)6.R83DXD)XF-._8MFeXH_Df/QIX;>f^F_]).GDQ;
^XF?&<QS6M.CZ21_EDQEYc##?B:bVIf<2gWYeRUF@bT6g3KMXDKEN^>,_:?f3-a&
<MRNL:E,04=RMQg/+Z#[BCAH]@CBQ-aJ_;Z,\Hg:/XaX9GAV&Da0R5#>TO;<0eHT
c:)(_R+XQVd>)/81(aMSbT+2H_TIS@DM;R+)=bA5SR9B<FX1HQ\;-DgN#Q?(:DYC
RXIQ=M?#CTN9Z90(>D//Z^HH/8\^=&,\^25CB]D3gf^3DPTLdX/LC27?Zb@bK>3&
bW,ZF/)dbOPBLg2bF-TaTOC>L:Y&fe11&OQ@?Df>C\BHa+2)98K=?f0b-e@g2^6Q
HVA?H_7RPLbV)ZI[4aaN1KN0VYXf[C->?.V\05@3K76J6\SWPJ/Ce9BQX/L-,\/[
_OdGM_,/E,)7(XP/F&9]N@e3I^;H-&3^(1?bV4TgY-[Le@gG?fRf5,S[?Ud3BZVd
/c4?Z.Cg1?PL.AXH+U\,LQda]F(W_1_VfI0[\RSD&VCOb@TRNZ4GCG<#9g+I=PFE
SN5ccR^<.NXIBOd8Z@;+)K9.-g>^CdbT5FLU#A3K5@J&QAa92.@X55d,4Bf(G?EX
E/S-:7,WD,-/>J)]O)ZA#aCMA[AIWWfHb/O^\-@a?bb&J,DdA>E72W+E+J&g7MH0
e;K5Z>a;,:+MM1;_X0NJ8?H6c2\PD/0_.cQ7@?23+2f)3WZQ+Z:0>54SgbE3UPL?
Dc/:#3IDH\Gc+f]N/+MUQH5efg+\-WK#\2-K:Y-I?U7Oc#L(AJ(J1);a@Z1T&72N
^dR)F3M<<\97JeE;31=)77?Y^JWE@[S;c;3QHFMK4^/?_^#2@J1F6((N=7THQdeP
V+--AA?fLB#b68IVHT:dP?GZ<\R>FJGf&HULa0MB0WHXg<Jf;?Rb>;cJI;?#GR(<
ZfNZKJDI@K<RH8YP4g>>0RD^ESb)b-Tc\VLH#ZU;@#eUB:^4b):3P6USIFb=bfN4
DF(9F=+[CUU9/(2:@<2M?.RMX#7]UT62.WF)7d5ddeU+CK+@eFLYH@4)7DTLZd;;
KTU-JNP6_=f:.WJ(U<Jg;@5RKC]M9D&1H<3/_)^PK5B-^<=M\G;RQ_T]c7H4:R;N
0VcU0^#,)e>2f3]a:JWE^DE8G1;JWR7.N?]Ba46@L^1&,cT=^N])JWX5O&XPJgR7
e8=<bUI>bbXVD&Qb87F6G?@\D0UY.;#4e,4<.cTB[(TG#&LMUDHb:9#JYRPeQM<X
Q-+(<7B5d75W\A>gVE1B=65810VGR]=4G,]#;DW4)b9=:dN^:=XYT=VdSb5>KgUJ
3-NgIT@FOcGN@c;S7@f>ZG;>FQI1H.FA4D8/>/;TWVN&bLZJE2A[50?YP/1RLNJ8
FK#8H;O]JHU>;BNcQ6/3;dN++afJf583>97Qb8/BbIBHJ8(U<>=#;(J7R^R(7XJZ
4C_,=ST[5I4fC_[SeS1,H[AD/fI@W.L]^/[IG+\VV.QM\J=IRDJPMDg@HW[#,>[(
]5e6<+STF#-E#AJ=ADdfDR23R^+9=cT<C><]c,ECQ93VH+S[.;BU@E[^AK:E+W\W
QgX;@bM+TP?CH57Fa9@OO5<.^a0RX9)<:JY=UNE#?TX@E.>O=aY>cA=g:ZJX@MBX
I:QcUSUU\_3GC?=2(KRcW6c/B7XeT#R\G#8?<2=DbK84.#+N?bcLZaC<K6PS2QBR
agI(3D-P0=27TJaX37(cBP7JHGG&ML,:O+(ZPJ=Sg-OUK\=#)1MI:.G^CZ\T(T/L
H_\(E:3Y&4dB/^10J=.GU&_T3S^8NV[KMGN0VSTVTOggRA8P@R[L+Vd<\L(75H+F
a&-]4=G+,._)+>NP7cYU(8E1Vb9g1S8MV+06ZCM.,N/B-+W4^.GBSF<S5<ecRMY_
#[>(9,>]KgNXI&+0D_Q3@gC)4HaXH7N&TgBI;BQBa.1C]-JL2b^ORBYHB^(6]@H5
>e6OP]9)5YSL_?8TT(6I09N[(Y:.A4c\//?Se7T:Jb2[XUBW9&C([S1f@:\e_-Xf
UH,3eH\MbU1d<J/7#BHN(\Nc6H7AVC50L7^aN1U7F]a2SRJ?SgBJFXRAG_dK&7VQ
Ca7L)X0U1VLd-,9YEP<6g0Ze:E@,/e:cI5VW]<>?W>B_(XLF1AM=RZ^W,)32,V<a
9--)A]-bE)[\YXcUN4WQ>7LW<0a)OE86S<W#LGG^aOP?3VB;;]<#g[PD\]HCR,5X
e#3R]IDRHEc2b[]F\?G3FTLLIF4,:>DPYY+RP;)0&cLg(W&?X9G+SP5C5Z(C(;4C
H-6<=7(@2Q7/Zb[6SR[29Bb_GeC7#5=MHfV5D.&F,B:BYQ:/Oa;gJUfR:I4HE[O]
Z\5#WSE+9D[Z_BJ)T8IQ,aCH^C3G#AOfVI?.E/VW9HA2@?](M=:4F&FcCg2R&-^[
/ZN-+.&fIdKHL@f#a+3R+5bbGgM[RgK[H1,[gHECO5PP;VD@,J@G,/g-EH;R99:K
O&^M1c\P>ES<g(AgH.HZ^V1IMB7M;L=@gMRHH3IK=1VK)M(=Xfg=24.[I?9OR?_(
=CFOW<Y4_]7C+KabQ/4eGfd\c#)[+S/5I>cDM0FJS6EQgdHY@TeLbdYK=Of3J5>>
EKLVJe5Z(Z6=f_17.@YG5&MR/_:POG<aSS72NQ48/0UQQ]?)R@0Z@<=8/WX2Tafc
-db,_M?35QTAe4]g/_EXOF4CKe-5PdR&Sg,FdHV0>S2&5g\R3\-JJ;1GTX;_.^CI
gK:.5f5X3\b-NJ#H5ENI__Q+_d>@:VR\X@DU/MGLWM[gS.cOQ=J/\IG@R?OS/\(O
71gU&fb,DVJVO\@D7+HF?Fe_-UK._a#27JfSI.g7#a&1aGaaG0Y^X(4be@UI2SE7
1-e9eBT?FATV/[D(KY=U<[2)A<;dQYL_IT)eO+DGS:f#JfNH/#MVKb5V@C8SO[Y#
X;17(4M2)O+YO4(CJ(B5J3<-bS@D4c\ORDeJ0O=(]HTX2/CTH()65EgP#.9(DTaH
CgQ7aYPE[P9L6_/--B7@P\Egef8V6N\?NV6MKW;#>1,U9_E[Y1\g4KKSbZ8Q)9Q\
)I+M3bV\dRL>B>E;FY]6A1PNGW>[(5ZFHV3TXHaL[X.bQ:/NWWM@@&-9Y(+5&6J<
R2@Mg+Y\^V1aA^[@[.>06f)T&>#YVc2P)<gTTd1YQ6f6^9Q>^b<cX1beK^,b?fIG
V^.c3/<,W(OZIaP./>7WMC7/F6G>=RN.UaMc)P.PY\c:I=+/\KDGHb\FC3@9;S8:
Ec_D&5Y2NIM0dDJd[6e[]a13Zd)eZ1BX,Gb7Y:[_>fc5KU,K2EB1da6ZX3R?POM7
M@gZF(/3^)7U;5H;).>)AV)d3,<DDbKJc84K&:D+GB8:[&I_0_OP+T^WC2Tb(5SM
fJb2Y9<_E\eB#92#f8N.685VdPf+X1+,\>=GK:[WG)GJWL1UO39_g^g[;0eg9_-[
HC1fI9Z@bbN5TAS/f\=O7GT7\,[/3BWAPI=8Q[VOXZJ&4N)Q0/Y>8L_c2(<G0e.P
1=R@I<&7K9.NQ7?FTJY5=8Dd(A<F(@,ONK6I=Ng5=QY&0A8_2<-ZK_+g8OHcDFN\
)bR<3Q8T1NTC6#KR]EM8[\UJgUf4?FZBfK;PNVG7762B#<aQVe],DC);;a:2#H_M
(B18gf^RBaD0+Q\9PfB4Lg>0._M[4UHMAU#_&egf?Z?SL87/@SQ;\[2H7)CcTKQZ
4S)[N_MS69JUD4E40(46)gUY.]/aE,B<;47ID(e?c,&/.EF2)OAZ9WT9P#P\2gWQ
)dW7+1QBU#NDB4AC(-N;+B_S;8U0U^1_X4_8B3U_/AGc[g+6EXIR)[/FJ8J29_9b
V<<+;RaAfLUUeg;A#>S17V18_0@43T]<2L>/,R)<SgJ[D)2\AO-P78Hg-/PG5.5d
P]B6-5.=96.FG:a4Hge&-f.]8+LYI^9/S4V=g4,(CHGg?c_8T#(>QHRZ\QGGJWX]
bL^_O>E2.AWB>S^IHdYM^Z2fGMHZ+.,/8).9bI?K9P_Og80Y6AC=S/cP>Q08aG-a
gXZc(XCW>3eVT6bGTO_P<ZHe)3Pe(M=dL4U5B70I91G63a6]BHb-@5SV5PgK_L:J
aP[JZ1((O/MFH8MK4[?SD(?R+/V;=b;VPTDdCJHO8(>ZE8[PQ<_RQ<eDRXU9;^BK
#\]9\g@?\>4?-Tac.<Yb]12OW8.a^H:adfV/egG;d?KOJgOXFAT_cEORIS(\&GSU
W.\-@>)CO16G3K2bG487)(9D7?]Mef,-NFeL+;R]Q5XPS1=H4QD#<EfQI.a6FFBQ
L@<9GC^-G[<YN7&L=7eB2;=I6+H273/:A.1I>QJ+,Q?^5:JC@>]64581I>89O(PK
-0S7e]\X/N/cD?OQ,Cd.GG/..Y+Z<MHC@_:5dR#33&OHZ\D@O2aWR&QVMDGeQ16;
0_=XK&.G)Qg.c9H)10O#TH<Y+YP9;NK@TO/.TU9c]BU^eP8P5JDQOAfO]DP\Ve4^
A-(^875;+U4G2+48Z-?[c=,[;VRXgE/6;R)Pd1=_fV^7ZTM;[EF0]LX,OMeNI+27
Ma60cU#]=f29CdJI<>XH4X]TKQJ?8,aANZ&0?ePg@GXTM&^T\W190.Ad=PT9S(OP
LQN3N#a>af62/GU?G.H@VMGUb@I@WSD@\c<FUHH^&GXRId?e\P,,5F:_bTe)cJ-?
-<Ig,53.R1M0OAW#0/&ZW5GMY]J5KT1W<b<12LZ[7QP9<E5B>=7(V^7\F8PWK[fQ
YRG=L+CZ3(SSIVNN44S.=&g4IO9R1/(VY/PULU8TO?WcIM7Q&gWUH+MW?C,8\309
KSD@=V<X+BOQ[F]W^cVaL,(68M@Y>0a#a-f<@/MJ=X;O3&-1fgIg4eL_ND,ee4a=
8),_P@B6TVB[J7ARba5&CRA)d55FeT)1DG2G4cG]E5;/Md9(+>0SZOeOR5^VE>3:
ZE&-MJ3\_#M8>F#FZ3e0K2FScRBU5\8AH6,A8&f3GECgc1Z9?<d,\I]eR.SL@_.]
_^8JVS:3NbXY]X.@-2)Y8NDc8+&+KQI#A/P-VW7B8W==#-AfAIB2.>,Jc@8\;[gA
1DK;,@8cf0DZ.6R5eUPREO\GFTQS3:C<<6QFN<Rc:#/X.LH&_B\^b94FG?EH:K1,
4([B]XS\:BM9<ET2\gU<QeCLE7dKdQ\#SZcX:?I+0gRK<XUde@?eS5(,HAI76B>B
^fd\0=eCT?U>Bd0&N>_+<4RW_aYC/OXX?)f_:7ATSY/>L;>HO_N(E4,TU4=cD=\,
GZQ8M]Q+TeFYAD6AL3V1\LfAIVAf#a]=]^Na[E@B?-0YJSN&7JYg?FGNNMgO#J3P
W&TbT#&Z6PW2E1?W3=VUTBfY4ZMJJSg1UTa];56DeR0U[F>Q)C.J&>:XX4/;a497
]/YDPFY3IUQdG3a,7eOD[/(M0,C@S/Z&(LWY4MSg-aMBMM7<(W&D?c9T>_f.6&M4
N5XO-FE[I4=UP8=f6X;RcFg)&<1Rf(7=[5/4+&ePFJ9T[A(e5,=_R.4T8T;75EPQ
&[5^D063e@RHZ#Y548X)>6(0e(@/;dU3P4^R8<:H(g(b8HRfTLRI[SZ@3\J2f/R_
d<?[JI]>^bPUa\F.eO3?M[8:aRV9UH[OZU-<]U/=61UO=dL3[M16_UI_&.f]X=E?
0-/>RDe+gY;1N8\?,2GD#Uf.(Wb/V#I0]RHOf3_96GaQ/,DgHXKA;/V,VGeQV^Gc
A.<3HA[OcIHS2?UXU21_3BQ?3]T-]^a54Jd4bJN<QOUPXg0f0B@BOcPDLB:OWK.Q
/K12OGLR_E]N>VR0-E3]bB9>]W#7c<HFKXD@]]GO^R&J8\0cE>H;HEA&<357]g9I
^c)#YBbDLJ>?g&cA:(LO^QWKLR0bXIc2#5AWfAZKMQcTVKed^,<2aeM13=2?2(_e
Ogf,B&6]fS8;fX]M<,_3+f^9IIBT[SP2g1L@\(,1Ed4^;2M-/7]5HMc>3eOf#)0>
FgY9K[YJDcK)VI4)5/R0M)]0I1c&.2>3ZS2@I@1+/UCf;QWBSdDe8:E6^/gYe6GS
HB6aQZA?GPV2-&F5G1aB&5RHdX0RgGLaOD@a)Le?<32#DP6IWefQ:RN53>6gR+.>
33[/cO4bHS6S4[W+UR#Z1C+.I?AQ98/PWB4.XgDJA]gK=#b_LH7I<K3IF<7+.?2S
=BK8AZ4.<a#^e5T:cP]L,=N[NJ(U0U?c,eL\)I<@YLTJ,6@E.4,BYTcQcW^N@KY^
@[4ZU)JC,(/AJ<@9W\:YaQ0-e:UR/cM<Q-J6GQ(?eN_YRAX>L^2/YMH-DDZ;4YW7
Gb@[NW.Ff7OSOS(Sa[TC&?g(TGV)HTDNL7+F+A^@1fR6+-#\CS35\(SLFT_4P^Q1
Zd;Y0>M/38LQCTD[=10]U(Hg6K;c<^\VgH=>bZAG&A0M21aR#T\3X=NADWKH#19T
-ZP,NLTEI,2)UD(?Rf5de@6F>.XAG3eML:?#Z28I<:P?ELQRb\3bSEO@&O?BK,Y.
?;CW=PKX],M0M^7K/-P53F.PURHBK4C:3agZ8+]K3=#8<fSaFIEYQ3V6;.?PR[6F
258U29dM3ON<g<_0]@WOe2[G<J8H@\8aH=,V:)58GR_:#]]&JbZI2-QaUd=adGe-
fT4BZB1,(^F_>H7]Y[a=T54e<A+.)dHI1,bNBd5R<3Nb4=6M#NgFLfLCM4H/dX[3
EGKW_MHAGGe8[dQ_gP-P+#bLHG0C#12<]KACJEa^:=Jfea2gbUI6aRbN^,4Ba.Yd
\=baAdLOW@0C>ZX1bd^?>G#ECT9Rd&2U8UeV[S^5D4LR^7M:1<=2DC1VHO5Cb\DD
C8_;59Qe?;c[5a=3I95?\J19QD3PYB3EE0=5f48M/<4@Tf_C,W0b#SI23Y7XEJG5
2151YA2.#6J>48<&+7bbX)>(e\b_0Y\<cD[.I3P^b2/U@Q,gB7H-eENJOFBF)+,D
J8KBP9NeI0V6O0.&<Ud):.7eaf16MQ#a2HUG-]<R8VQaGC#K\d;T,#?PR;eJcaP>
>1@XR3_CF]3aT)X()N,0a.BIgT7H3a-3XK2&XBa&6NITZFHV,c3a@-aYI]CRF;Le
E0,Ld=F>N91]QM4<4XYF2eZAa33T.V[g6G),#<)G/+Mg_QXgCPOe/cDM5E>\PD#d
@E9^ggBIB(,N=>7+G7WPNZXP?LUEG)]K=NHc]31cWg>CbQQ9:[g53V]]WfTAgKRT
IVVI?4,JT9,TY=L4G/d[RAWEJ-)_KC0[d<4,K?R]UT5639\VeBS:/d&2OUEdWS&/
AMF.S(M&\_\eHf6e-8B-dG2.c9#_1VMAC)1+(HP28)]c:QN/FSVM5PW5+ab(I9dL
>J+<=]aA4&>N)2CMA9QJg6(WX#4.NJ.UFI+1:=1XM#aW=J=,?^5C)ZWc]6_O[.4;
T>T54&8[Zc?XT\KDZR1Ecgg#RKPCfB?>:(cfKC-),/)f8ecU66/UJ#5MG+4ZT/cO
FFY)A.1QWPK:T._TNIONGH7fNWg(Z,#:00DB2I5+H65-,69]B&L22(SFH^LbBL]V
-W8MP&DWDF#g?C;@9ZQ:,F,UcE,2Y71f_7.GG<eTR]bHKL8LW.dF)R)D5_,)N(7Y
GM];+FG<DC4XB/^\D5cHX4-68W:431?eJF-+aId:e1[_WOGMZfcO<Lc:\433WW?,
A[C[#1VgJE&01VQ&6c:1X3K8]R<U1##T0.E>XOT1-b&LLP(7?ZJFT=K0I3E9-,aD
+/H)=#ZOcLMG2c]6SC_+SMcSX6<2LGJ/b9)d-f61#(c,XG790;#UP/<=02NO2WS[
ReD#e#5;dcb5])1^_0^6-.eS0a<MGPSaGDA.:W\\CC#ZfFN2PeMffIQd4BbR^X6M
^#EB(<5dSL>Cg:gG7CXH7bc+SW#e[aRb#:3YC3Tc7/d#ca1NS_G.+K.KAO;-D9(T
89NABR7WUG;9M)\Gea:+<(E4;FE9KJa?0@9(0-gGOV@CPBGI#OO/FQH2+[^RQ=K\
VID/VR]1W8-G8;bLQc#+fPRN6CQ].S#&48892I]843Zfc.e[:0YSG2)V??+:EC[J
=;N=EX&^QS44(_A7QA+.T,/[SUT&\7:/,<C@J;0TD\d+;Z]MDYb\NBWEd(/_O,S=
=gUZZ&#Q4<B8<I;g.IV_/A>XS&H;)RH#g9;fX]26FR.U<=:5Y)RR;[a68DUee;7+
/CKKfecTGg[D=OK7b\CFT@HTC7N=M\<@9_)SV.@.1JN[Y[+(Mc?\]NLGed-JH80Z
^1M=HIQE[ff[E_W\IN((N87C@03Z>97A-]g)OES?A7ab&eBfbd2S0FCHa@g>PN0;
=g/[WC/a57&>6;g:.V_-1U_983/\F>gN4E9KY[2[73KP4/23A<Z8(d1ASH9<[?b/
<.Y2X71MKS_NE[//5L@PZY8ac]fAd>?-T&Rg/OQ&?Pc;e,eOML&9Z;f-ZEFF?:(N
+C?FBgg3A_>96b=g7Hb_Y#L&dfcNER2ZHd&AJ:UL-PaLKCH2K3@[.V6U68[_ZH5<
RQJc^2@DE?+9E0Q#K5fO8W&[,/KQHP&#/bYd,JZ)CNaX,LOXGR#GZX8F2-a-g+=<
OP>Z=KH84IO./8UN]@^,D]YET;I2LHdYMR9K\E6[@OA8:gE<@S,PH99<[Z4HN-&g
_(B&2EVdJ0dTWd<[LV)^G3WeAb/#@>CGLf;OM<6Ed3c/cD[WJI1P/ecYaM(U(+<Y
f2)>,P9^Q>4;]6?Tecf9COQa^Vf#C_44dcL@)[-]DaFVUf1?Z3EASJV7LA];-AeY
NC->^\X.cIGNQJ5&G8cFSB09DHU-SZW3]TXHL96,GFJSD_]GTP+\T;<T5RXO,IeY
^:fI)VYO35^1^-\6ZfT_1W3HXC_>REO\RfNc&=YgFe8E8DO)Z/Q;+8_ag.C[R05f
Y62CDedZ&]L;+bYN>W_@_P;2gK79PAA.()<;\dPLC^PH_Ba=>@Ra:J:KR-;P31AQ
UbVcT-gJ);eC_ZK)DJ<Q8O+B8#6?E4K+(,ZNWW-ZYY/Q,<<?&Qf-3)LS-BU[CO&f
X^0b\2F,:X^U,@@75O3PG@8\7,FdAWNN-X@,J)ddJZ+.\dIYUIM[(>3>(A#-T@91
4Fe,4Q7^1c[U3Q6D\0K@M=ICT_/+<&T?SE_#NRFBMg@4R;JS?@dLILK?R0)N>M3D
:#_CFXI9Hb._MPCSF4T1/-P?H.S[cNF5=@^[0:?T,754I_S==UNSTH>-)\f,[]04
(S1VP\.=:[IAOT>-I.7P(S-N=)DF;]#4>](;2AXQaaUc:OI:E4&\,A>f>]C]&+X9
8Ge9g2OIYS/f,8DdSOG?G^bWg193K2+FA(Y0&W6:C6MD^Gb#(QE,0@+AL59)+S^S
TW&X.L&]B7:+g=fS8Bg_6X+1.UJ^dS8>>=5&dDEC(W3FW@f)dg,=;1)&3V</VC9(
2Zc@fHH3^d-ReF]X/FN3:(8A9/+Kf4&EDQ<2L2MGBUAEc2B^MF^<TOH@>Aee8U5V
G)eZHI.;[I.F>/Z>;O5d_#](4>2+eg4aNg+gb?YB_c[SJ6^U.#BGL@QOYG7OAT0g
SDE(E:^/Vb-;fB[-R6.-5[[;4Gg@4KP<YZ@N05S[8UWb.&cG;3J&#:_E<E;N3I>9
TA9#g45UKNILcMH_]7B\HN/QS-Z_@[5b2Ucg=eZYW4TC:DMQ(aTDT2]D0:@U.J1I
Q3=.=_YPE/CT>YBY/+Y\GK(3]IA:Y#>7YMc^LPG\e&IS/W]fGdR&=_ZI>PYL2E,4
3<E(C,KBVL=Q)eEF@5Z.aZ.R4;]3H>&85LMN/:Kbf0^)#CR)^6./^;K#DC#QR&:4
.cf?f1)U/3F39:?T[#5bLYf6OCU<RM[K+[4U6B]6&DLTB\O#@/fEG\SND9ENI3(:
UeG8aM-1>]Y/YFgE:@U^dQMX,D7Cc)a[;^=<A)A.+e5We+]K)O.-C/^;6^VY1IS\
X2:;2-_1cF]PMf_J2,II9<E,,eTJVd:gbfGVAS+3LC=(H>^CC5TV9TNN&BT^&./F
gBE&^a3gd&3=)3>T<JV29ZC<dOVN&#-;AcRE[BRd&f;:OU2CGKU&\0WI8;X;8EGD
?HV6bO,,d/[RW6dO@IBHU_N<(Q;JC5PL_;H9)6D6dLC#O(&,(5]])EZ]R),g7?J-
CcG43^\BD5OW0O(1<IF#aNNJ@90gEK2CADW[S(YGSGE:E<2Y5d&/G?YYY^UYWGXL
_8C+Q5KIUgF\R>72U71UG\Q)D&?d4A(G7cHf1eeCME]BL[5ZRGIU=ZAY7)bR]5]C
(ZDZ,&N<&4+-egPBQA@WFd4-Z8@JFeKK#SR0)gEFFMgD-QT37bdX>W6AJbfG49gL
2<-S;D7/4G3/V?CC>SZAL8L+/KB)03P\,18c[G/Wc)L>>HG0>eeZ4N.O]Q8:[^,H
,-\#,@8IcF#VL:Jb&(N-Z3+,R,EC+JT+:27U+M>Lff_.6/Mb,/]d[TI<33,E0cBQ
>[M@KH:RBed\SbWc[fSK1/E.NOBJcL4FeVgA-8?Y,X&aUTKR;F59A@URAL,de\J5
gE21YW9_=FJQd?0\I/[LCbL7c4G9[4B(F#UDK3fb</CP?^=e[c1E)I;O08S:1-FX
5/SFU(L[&;)W?Ic9EMRXHKd,L<>#/:&f_\5YI&/aN\6UF?fAJ(<C4&D@W=\?)Q(N
KH]bDdd3c\b/,\f6Jdb1TPT&2LGHVLb_]\TF1d/X=c8GZJ>g3<e],DKQV<,6>0:O
fL+E[6F)CF9gMFOB+6MRP3Z+6-17GR0a(:WDN:b-6@TW]08(#a)>YPQ/E\F#X23f
A]?_e_>FCM</-W[,P#7a[Se5a4C4CVbV9///beZTY5c@Y^c?f9-(e+e59Tfb\.B[
5YX486@6\-3+[=@3HL)CBI3M7G0+W&>01IFLcP>S4\_VC3LY)O-Vb50Z0KBE9YRJ
>^a:BQWYB&[g:BE-FWc7b++F;&0(6E+c+:W0K<gW6Y4=<JB3&_FI8;U]2[7E^BW4
>7[RO9dUgacAS1HTKbZJg-ZCcHIaaQH2]B@BG]SQ?BEHL#9Z2=.(82KFB\GP?IfK
+a+2#UU&CgdLc;dJ8&aA(AY@STE&,ZQQ>_XVD,K^&Y,TUN()3aZ3(?/a[64PN/+b
=/1>Vdb1GH^W-H[TVRa@LddDceEXXfU@53fYC<QK-L#(U(&/0E\6DY?/6X-?TYWg
Y6@fV:dET[ZK?+P8;0fY;OA>@(B0&Va>0@4I4+VE9RW\7;AGE&)T+AWYf@53SE45
)SC@2IR:M9[3e@9PbA^JA)>aGY=&fa,XP#4HXOJUKD.GQKFR4XY<>C\2[K2T(;9;
+C1.BGZ_DZ,4K;LdUP4>C.,107V#U]>M^LLG/A^XK7^_eeeBYVZX/[GID.E9;(HT
\//FKHD1P1C3G::Q(GeI+3a1.b?[_:6fGPINfCEY(b7a(ECC^KHeW\P0[2)#eeP1
<=E&+W95YB&/ISJ:S;S@9cODDAQ@g_;deCIc.Of[7,4T4U9[9\\1Qc:L]-:[1<W^
@UU=:8d8CLE&5B<KF++RBe<cD#W_P_,EHfc#;#=TVTB?FbIGJXG=dZK]0@;A&6<J
aaAK:K0B3P\[RdM9c3G&R,9H&XDBca8cHRLBB/>7NMX>D2<3(-KVaQ(\;9B]ScB/
eVR?N+BGd21>e@K)@KNKX[K](1>H?ETFY#U5Db>8cOV4]06GD.T>(WSI[M<c/GT5
dJ?@76+ffM\0:#V@SeeRU5IgQdM3D:Bf6L7UN/SYH=f;._VTcCX1+bS\PcfBO.4=
d099G5IL12X>)d^1&.N96Mf[)bD&J0\EbD,=[J5/I;#;W@DC9IWF255&cA86\HC4
DCG;GSO[)#Y#-RLfPb:U78&5^:K7X1^:B\#aU7)E-EW^EfC_[^6(3PbR0?TARaAX
bAW59D>c1TK-&FY[/f=\S9_DIEQ@2G9LS,9;J:-DgfTMO#Y)e<Kg^7<3=.XO&\&6
T,bH8_V4;0-X.O<:L9BS9E;#C?ATS:C9Y?VcB8<2bIQM3X,=70(EDID1;\?bF[W0
FAUT^NQO+@LFP]4:S/>2-0:)7Oca1AX@102-DQgg+De/?FV^.,8A\<S8_X(JY]VP
JY=Wc?=RW:@J(fV-I\>5,:]#O61([dU@HT-R^G+DWdH4N]6T9NgYU(0.^bL7Z?&a
K9O5Ma=^-,P0M[?>6U.;+S)Q.;C\3L#)>>3;^ZJ-H[g3\d4fVU;MIa5a;5;U\KN0
DNZC>Ra;+[[MVf&TPW?B;]GcEK[@._,DO\&M,Ae_<CY3)L6e9.38SaM_eEQHD6UG
AdA-d;)URL8\eBOYb[Ua:E@N+FEeRQNL>AR9Z1VG^,RSRWMX3#DYX-I]+603>G)I
+#HA^\ZOR82gB#(AWOF[)>a2-0+.7L=1CWY@.VIPWJ-H#:BdCeQ&+=0L(@KOQZ:D
LKIM\DJ)PY#H]X>.d>FM#X93d=Gg73E&:V&9E/C>7=+OUeJe9M8R#1(CF_Z;#??=
DD<YUVgM/B)#[#I]8fa;=AbS:UGbOE0e)U\_0Q1KSK=?2Fa:])@6L4)L=R(EJd;.
PJB[e&31T,))5fAdXR0MU76&Vf^RAca^L2cAJ1_-0L5MCf77G8f:9V\2##?91#9I
9C:UBCfQf+(<_Y<31A&]DBOd_?-6,VAW&?\B-ED]\Wf<6,=?a-E,2R>3EVbd?\BA
@9X2cBC>+^G57U4AV_HEF6VcKa.@aWdC>baKNLDT1M78<)G(gR;Q,>ZT2N,,A+A3
D]:G&.@25f)F](D=4S]^:<\5)V([^6EBACZ0N95S@a9SJ=+_M[U)Y56>97^:D[A?
Rg#U=-SUGOU:f?)eG<XA_X[ACHJK&1X<IHCT5d4MZ:?OG)_2\CI^[]B0=WC.A0B:
EXMEX=e/IWZS>@BS#WC;+<BTWSQQR19FJI.Y-:(707_WQ6ZFbFT<^1XCfOJ7RC+0
KbfL4dT<WTd^];#FEeI8/:B7@3A@9U<R?dF0@?38?fCFH2@d:Y2/5EE:#9=GSQK/
3:gX\\7c1=g6?8UCA3R_;9GTc5>gZ@OA-cQ\:[FAZ_]7EbAE3=gVU6;VM<U6#/X7
7HBXIg:DCQB276/+H>0]1&ePZ2VDW7X-f89d3_SB@MaOG7.HN6^0<WME,(P]U-T)
:GNZ^F84P1G)-D19)e0^I==039[;.3cF#3TL+Oad-,C01.)U>.U?RDMT5GOX&W[I
aHKXEF/F;LQ\&_JDYF<:(dX.ET.W6Dbb27+<\BF5P=XOC+82[-Y(\=MPP-)C<.W2
PEAL/1DVRQ@K+MK2RT9B,B9;d6\[XMG[67RbS,S)<)0Q:3Z76-?cU&NW<J\Q7]=?
J8;6A8XZ;P/,IO3IJa+O<+\cBY;g;/C8A6ESX6W[AQ[.VJ]a;1g5V\EYU+(Q1P]+
-7W8d#T\_O]UPW,KdI3.MM1^5g1RTC2TeSL8V(RM8^QCD<FdK+Cag,2dD4?;_+0a
D580BKXW6P_@fJ,9U,QHM_BH:3/SOU.Z+#OTYG^E5Eb&4BA_FR)Fb+eg0VXME1UW
\(bQ0_[)HP>/?0b^cZ,KeQXFg4K#\L[eQ>7@KIc_b#5GT?/OePF+_f5L;5EL[K#V
N[ObO#=XG@G,_]M2\d1VLA,+@YU0@;\_ZZ19Ug[5d+[([dM-^WINRJPfIHAMQSI0
28[E:GI/e.<R.4)S^e^Mg#a<fT79M->&<:VeR7@:=;#bSG9:[3WfeGLCAB(GeCPQ
N8205Yb(bM\0IMT@gGP0I26MM>Z?PXG=B/#/UFgNPg;/?A3KcV2HVTEEVOLOO[A:
^7+KaVgbW_6P8SAaUGIE]f7eWR:)=a[M\&]?@7;KM96TWM9&c9:40<;bQ,)b8)G6
?+?LG8d,_b>>G<IDg102+]#4ZL/ff-CC.H<6S&KRJQFY6&YLDC_MgR&0J?I_Wea:
,d[]gCBdG2D?X9K-YK>EW7L&MDY?NM59aE=Ea@3<B#._6:FL#ZN))T[.TL^9aOMX
237>()W:b7ND,ed@JP2C2X&D4IG/9,CGGIggX]RSced[d=DeJK1E,G@X;;2BI^@L
S.0;dZ&1f.;NQLBGZXB/:SBDRd=MOXbZ+9))@S5)<PDDKSCcLWW>LUOTLA.R5+9T
KA-.S<;D_YO95+d/N/0T\d4U?4UQJ/-=]RA@1gK)4LJ,B)R:(Ya6@Ce<6Q</HYUC
OSA?H+.W_[SIN_f]1II;[=Vd-eE=-1.RY9704I-:5@-03Vb6R2DbV86R46VU5=P6
DfYYc59<WTaKNN[KOP[fG/Y\X^V0ER3?Pd,/=ZT_V:9]_ZS6fI<LAL<N#FYQLE/H
-Ceaa:=.:XXA-JW/NA,4([(+NZf9bNG.\\SWA(0,ZAH+KHdG_&4M-NA9]PHP\UB/
JU#DF=^ca8R<ZMV7UgYZ3+]eUN>dYbDED?VaZB\+?BI79#\f/4Y[+GQMR+J/BUH#
?CGN\MGE^1RA3ReRTPZG5ZDB-f3;d\6f1>5>N.=aBY6aBD7S/Y\_ffI?7;X6IFeZ
^QW:3EU@-9f1D)WJD5.C3dc7,VHd88dD]I\3C0GPA,d.-4AJHZDZF(+O=?AWB:0T
)/H(>VPG=DNfK2DUQ6C=ZJ\(:8TB@d[BP9Z3Ub&f;P7J-4=e+eVHXY0eJ_V25F)T
2:=@Z1BFY.6>FUbH/g41].0Tg^cI6Vf0KcW[.1#[aUI)8Me)c5<>NB<I5X\6>]L7
&/M;2O?UB)YC7>?;6b/.:9Pa&5[VfN]VA-+UN&7=;UEY>MdV\&_Bb-:NDQ3U>E<3
H3fTO193b:1D4POfd/H\[9YM0d\A/Z0]R<<749B7DLbN6Qf8C7NV-1fSPEN1-GTA
fGA,bPV]Bd[6:QZ\(7>O5]76Xb3AB(RO(XVKBA1?QCe/:X<HQI;>60LSSZ0#3O&B
)GaQF><S>1,N:cceYR_1C@_\G;8/f5(OZ7dS=@V@f-3c+AP_>3Y5&J\4QGSM<TU&
ASSV_c0d6_C)c3EI<G5bdZ=1[8-M&4eX<Xa7PCV[M+/.^CBP<[Hf5fYM0R:YJJ=:
0]7Nb=&YQ[C-RME(V+M0FM]>X<>_I]4N=VGKA5XB@7S)5gRFbW0+Y57WQT>cd.V(
##N&W6@8JCDdZ]9-^1;a]eQ7>-KC-Q5F_97:e&P?G#HARE>O9^;P)XgaHX@QKN_d
A#<7OJ@GJUO39c8ITaOF6OQR,fac/(O-.I0e3_)XZ9.=;8c.3Eg[/[6W]/[,T/NJ
,C_>_9Wg6-3MI&1@g_5F?C5G,3&P<MV22+0L3^&HZ>[f=6PZ6Nd_;WA/Hf(S8I-1
Zd(2<P)M_BTZg1:G8]IMcX\[cO2#3.41ZM,EQ5DY6/WBQ.Z1T5,M^^4SIaHMMb9C
c8@WU&G&2Fc/1cAHCOS81(>[MB^][Q==TXEWIM845ZM\M>3E]g9e+G6=H:S,L+(L
N6YZeS2/faM<^a=GOe(34g@HK_\FEPdDSHT0A5C#W#Y)>G_0L;.K)790f-)Qe[gH
be,6&YAaWSHM<;:=+VJ6>8a\c<&BX5ZLIKQ]1^66,T8SRYF97e)8WRT[#&.7]V7S
7PWH7)/0aeT>IV@V\1-TSD;7>Z_M]\)T[?2LDH0O9(#^Gd?Ncd=^S011=UQa^J0O
?4>[\VEM#aV9++>PLCZYW?+=?[AL.g^@ONeS[&GK&AXA>>;ZEb\Y;V4U6OG/Y/:>
-AbCa_D@8?+F)/R=O??N)KJNc01H.XJ_QFLLE,FMT7/\[=A6e-Gada4DABGC0,Q7
,NU#2-I6_>=T-@7-I6aO=&9VQ?5E,D5SeT=:THW=#.EJQ_4TBU+)>#ddS3852\Vc
_W3G4A,INA?8e9f]3[#B+GW<,HRUR75/\&\PR0f[5YdB&+@#?:D.?#.KNV<.F-^e
MYPXXWP<+gQ4.g6JS01I752LeDSVS^,X-@9[e)S2))M<2fX)8b-Z;-KCT0e5dZS&
R:)_7@C^/L-6S,Z;WW&O&ZGJ4T&W+(+ZLcA6M<SUe1QLN.I:WIfGY8aX#_KVS5SP
AdXV[X7>)/?:SM.aULReAcTBL8B8Z,_Hc][bT<8F1@:R.N@:eM;L4./Qe:@=61+L
TdQ:N;c3<WB3W7IM?R/2E=3P-I3?Q^8DdX1:d0Q@/CH]#M^_]RMV34XcW\IPMMbf
[(.1HAE/KaXJ]LMB)H&@b/gSFbYPI3I[_6-WUGDb1>AHBZ_&;C?O1YUf><&NgK(O
cJYZ0ea?P65[>Ee(.S[/@CDT>eA@;2Ig.QP^@NQFMa6\^I=^O2GAHd8-aeYC6&+#
e(=ZA3&/M4/.-5XWIC\NB4#J<TN)GK:3R?XDcd^aM(bAJFaL97-,SDCQC&9Q)Q_4
P(dQ/H,dP05C5UNVO+,GNB(1JVbD0=?V>8(+#4J+SCgE6M;6Q-DQJ,O]M#YU7.LC
ePLX_d^BZ0]4(27W5)Wc^V<@fYRJ5#R>g:Ic#DX)OKRZ8a/ggM;d>/)[&Wb>5E#7
e0;\O99b@IfL#(.&AeP:E)&_KCKEb&dJ.Q)HeQ@2=-^+=>R+DO#QW.:RYPMcU=3H
]IX4LZEd<LJN5B&<V5P;fgdVJQ;\V&)Pc(gVNM]H&A>Z)1;R](d@:9\P_eS@,&TC
a+OPKg6F6;<8P9&?2X.aP)XIga:a=:(A3+YJ4<e^@A+C_L/H4]T35FR4Q,/\g&Q(
SKc.,cXLP.(C>8O.DY]VGeLL;+d0XTGSU11<+cJ>c4<-X,JgKRU-&b_d83Aa3Zb6
]HfZ58.N[EZ(,\)F9J@M+<X:,XT2RGe604XL6I9+D:gYDF3QW-7LNZ&ES5A-8A&+
>_Me@+JVZdF@3H2B\.DFgc]J4(@ZE0#EKc?Y<4C[(]?NGI0L&&\:c/C9B/a9L/V?
1;K:Wd(;\Q+;2Z75_ZZCP5ZZ:ZXe.dOD)\<D+OZf4^aPUE<T)-5X#_W+b8R6GHDO
-6DgY),+X@\U=fOU,EH0MEcI2M8X5><[g,H[.a@\DMI]MPe/&/gZg.=cSW@S5=;U
#a)_eR]_#X6?K)WEZ?CV_HH7]/&80-/C-73@MKBE0B^PKW:M[2M^0T=5)e257O=>
A&7B[>]T3C[XfX5bL3_71;S^+D.E#MP4C+YE8OPf<YD,YXQ(L9J_d;1[OU]-4TV;
HF>aBPWTL<&+P]9>X3gU\&T2^&1CN:J=)g[,#FH5OQ+9M\#K9U^YHQ.\f_[\cF7J
X.d-HSIcZT-&#<FC8T;d>N).6I_aVIF,;J:9f=C\I/2Od2,ESJ[R>IHUH5]+XEPD
U:LDE;De(dCCRLD-TOIRY(5S2d&AfW07[VO=4C7H1@3E?,=(VbHea8e)fF[YW50=
eT78YaYQba11&GS,&@F8N&)<G=JRb2^[[R4f?(+NT<2LC(]L)8?L#).1<,;C2g,F
NL(@gTAf<GbM@TLNKJH]T>2O,_>aAa2AW]_/R\D,)Z)9;5=<T5W28/ZZ<9b,(B+^
A<VJUg4AEa]W1;(34-<-BNSL[I6a]#JC5=LFcM&(N9\9D3.D>bgC^SfdgNb?f?=-
d^LF].f-dPdX-CbOR72]51XIa6SJ^=4535T&L?8-N2.W-8bN1A62Y]Wf2<FV)S)3
07^?MQ)cX0gF><;.(a03#4Z37T86VNMOXfBR?4AP:N>KRAc#T-QQ2A&gW.f8Y[[)
ZI(1a;3R<SZ^>^9E.AfF<)ZK_V;>a1N[(+_-f)g\S9-9YL#EG6<@]6,;:b0(R4=R
W]MEdKLaG\9427Z>IeOC13:G3eO2L(ZYf/(#Pagg<9\GAM.:(-/U>O-1EVH4_C78
BL0[I)5:7&ZLML?f+c&.]#(@Q8P)G;bMRe1W7I=-,&0@5\/P^L,;gIPg>+XgWO\3
<[H_-2G:?VA.H]:&8>XDTTHCc+_H#T,)c&=/R##B4H3J?;2SgRUG1-^H4d#N/1:a
5M^;MNLH]<DePgK;??(J(Ye,Tbe5]2I,aBK.f,>D<2L4P315L5NH)Df-Ib3FMY28
g&5e=R6?(dRW)K/Kf[W&V6[O=[.@SML51<[cV\0PHI-d,W2F=M33b3E#=X(WaQ]=
RA+RL7<+_ZD[ZQ#P6ceJb,<XUJdSVJ^dW8.^UJUVU=N=Oed>e.N3,CTYO)9/gOG=
/J1e)?E@a3KQWMO7Ua_M37.VTN@;@6,YB<=,c+EYH1Q)d9(RH5+.C8cXM^,_dV,+
XXG_MFf<QaYHGL-HJ__deCEBF?+H8X9gI\AC;=<KC\9aZW.)7D4GRGb)3/_H:/Gb
A&+@5>V\_aQ?Q-#d</baec1>I8>];M:1/E83IA<TZ\[77KR+.4]X^UJ(bM^f&RYJ
-&3:Z-GVCDC@?9>08&(/KY_]UM2e@)2J],-?cR\E;+f@H6\fA\<2[Q:cVdE9O\1[
V9]+Z/XQ4,T^f^G6-_XP#Y6T;I=UPVDGES?U&4Wf&123CV;EVQG/&fVNJ3#:+:RZ
-SQC2fL)8Wa>dQRH/SA,3OVfcLS[7bRP:BLQ(EE7+/^OOcdd08]LM4)eRZBKF7>W
(c=L2IdM&T?YT_?M67d,cW[TT).f@N4cgbY6Dg(G@SC(@.aMLb[>L9Y#C2K041L#
O2d&J59S-KdXfJ_9]d[SE,9W9;UDBUFJaS1VR.-1#@Te[.aCPR4eU(S>_><M]2)<
2Y\8;D^g0/68BR1WeW>a.(WL,:APBQN45;-=X/WS#\W2(1);0RfUWY_MZHAZ>C#@
L6.e+-g[VG7#f^WN/107);V6@8UL1SO\Ca1KF(6B/L+#H;-+,_/JWP-VcE[2Uc4d
HJb0agdf.]0D<1(PbKe,(F2.E+GdP5),JEWL#259J;09>\U[1)Qd+XM&e/>##+Pe
LXN+d(_14P<9NaYT6D_LcEUC?c^LPbPR\>_)U.^,YR:NedAD9>DDZ#;A5H/c8++Z
NE44gAP+L2-BCJ(+3IR,U)cG4&g6\36AYJEQg,dSN,CFT;]Y8.3eHWH=1(S2@b6V
#Y-A>00RFH5W?fPT@5Z#-bNF.H+Y,[f[P><2-M_Z:P0=a35d)-HTB(E@YXWeBVZ\
gXH_S+RKP40C5^U37X<XV96(8QaKe@dgNY(aXCL7e^D:T3LbJ^_TXJ:V8L+(Pb.(
G5:#O-1-:4gKEU7.3=1,H&#_2;?TW&HL.XB4B=)Ee30+Vf8#BK[XG/O8>D)3,RR9
]Xc\g4E[]0ZGPaK?7L=94Pa.E:adK;^?U&g&[X@GG#=S9#1JJEI-XHJEGF7R.(WQ
FI4&2O278+P=:SRGTc9UA>O)V2)4N;2baaE7QMYB8&^B0U^VVG:1D_,,[RF<;EZ<
W.1fYVd]CG_X&FT[b>+)+BgIY>((/L&C#D6^<3825ZM/M#@^dU7WgW7,MW,I]O?f
@@,?RG1@3SFB,\c.5a/>D;>;60T.S:YEGW:&\@TB0V=SBXR6f1GSUF@1V&.Y@4)&
TT@8U#TA#8&9(O/.P2WA(@U/>C#[-7J#A/<+LTW;96BY,.Cg)W<//=Sb8C.?DJ\^
M>db:b#HWfX\A]OD8Hf)V)^)N8I:e5C+4#5>R-ebF9A?0RU)X4VV#<WS=D-?#gR@
U6U(XM;5VMLS:Vfda1PCRJ@;C4e,1#[)a5S#8fd58?Q2A=XD,+E59Tbc,P^>\f&f
4KF^5_1DRd1^+?BW#2Y:L0;YTYE/E<@c]X9b>+f&:IRW_2S9,&R#<a7dO8DgSCOZ
Z>YQ>HOI]J.;378^TfadOBP29:OffU)P_Z-P&&^ULPS[62^L/<<+<K@;WbU]6<cW
8+KV2dG,V@LT46^C\Q4@;ZdU.SO\7V<9W3W?3VJ^5f3>K(]EAd1UeZJN,gP-X\L=
=^14W/eSGbGT]NR^Zb-AP57HQ\&2^f,OR@C=d/JQ.UTG>YSAJGC>O.Y4?83]gSTE
-?.A..#\&S.fQL(YaP?ZbN<CDR=VfT7[_S_b3>N;?>V5@IZV5G976#=@3(2gcb2^
9L,P5N]2CU1b/bT.HCJRJ(-Ea=dQ0T\&84BQd1Ba1G9,gS)4Z?5]cNICd4[Z2Ybg
SGgfG\G.T.,-\<3_IRLYdZ/fXJ]UV?P??Q63&B3:,)L;]>4).KQ0bNJ\5#Z^AE5E
&WD/0:6>V,6_C/.8\\BW4b<6>G(cRbU>J(OJW4\XWCa#<S&B_ZTP3]#1D814GDM1
5]?HJ3RCUMG],I/11N](S8EX+=f2>FY84&cI1)POfd)b@-2(OTNQ9VO\@?,=&4#W
(LBe>I)R=TXgQ:N+35)V2Rb=L/<5#<Ue,Wd[XJNgO7(IB[<(?+-R5W2=8(G^<F_O
2/I5)(XJZA&,2gMZ.SZ7_2#W\Ke+fUD:b?.>-fF8=.;WF(XQQ<+g+0[_fVCB^Hf/
0@X6FGB.[KYGb@GNID5;9TKA^gO,5#9+;4#R3&6<NUP32L6JP[S43F^G\/_I9T4>
LF)HN1NHF?R=R-&F5/,+e9O7&VF(4>B:)2[;OHE=b)O>??U#QP3+g\[(.-:];\GS
Qc4NK:W^SX78LTUEQ-H+:U4(d\ZMMd8dM[+IXFUOfT[Ee[LY_@N<4Ug<YG8>6S[8
,^JE[NU)]EFadHTg^CJ(Q>3)5<NG#ATM#5D2C6T=.a.aPg2OVEfHb\SF>K&PU]2E
g9G(bEOA>(ITA=Wc;\H1gXf\RFPC98ab4]C1RaV=c5W^=RIOC4EOGTQ0Wc=)YGJP
d2+D/[3UR@PCZ-0Gf^U,gZ&/fNHC8bW2-Xd-f-8.K;Cbe6e#WB9/@dLN:Y]NgHOP
/dN<a4XK39gVc8-C:A).NZXe\S7:bL8<#\2&2:eERR/M-P\(:MN&Z8/YFIMM)1.B
:-AE.KK-0A=)7J:T.A;MJb7(Rd>(W\T+XQ._(Q^0Sc[0DeJeY=[7BAU[6YdM?[=(
04OQFbCce1X#DdNUQ,Ia/BN[7P3Q-gL[[-Y^Hg03:?VMP(HL=-9S.RFZ=e&,0e9P
N2RSU??(KELNgT09Z^8beLU)06KDIXJ&ag]Yd904^L8WCfGF?4OaG+&7X29#RVZR
D0EG:9bZEG&PF,Ff<[:[A^UfJM45Gda,;\U,8gE4J8eg3K#+U-2dDD0]a\?@Y:)J
&f#M)W9b:,U0S#7V@TSI8:<GC0d[VN71;[dC],/<e8fC3I(6TJ=-I.N\8_,KGQ][
WQ6Z@6_6RbW6d:dBU<Q:b91D:AbbG=CC>P..e)H(aIdU@.4HfV,C7)M,6TgNbe)^
c9RHOB[[[G-^8199[T7+c^SE1O.@E#;[QSg^a)?FIC;4aJLeO)Ib,+HJ:-5PTCY(
AMSE6>8FSf?aV6Dgb=aSaJU#9P4MUe>EW>6363f<f^/S(88AXNN-W0P.6N6BAcWK
4]CAX@[;a^2&Mf]1I/U+d0G\HPVGaZ<C^C#DQBdb=EQ<+#6Z9a?<aFfJ@/Y]/R(F
@QG(R)IfS_##<gUW.F_@C:)A_2(YS?<7QF0d+-c\=PU,RVTPU\/IAbW:fVcaIP8C
V^WPR^3.=bOSBY?AHBA(?N..:dMJPO,T;ZN\77NEa#/=ggGJP5d\W7@B);U)1XfM
D,44M_1.;V4&d=AQ:-,NQU>S@gB^W-Q:#-)c>5K@7K7ZG1#E<0E0#>NXR5IdAW11
U5T[P.GL5/]/+d;FYZAbK;U_M+S(P=GOT.3cI^F3UBPR2#Yde/58M_9EUePA<\U+
:MKD8dP#TPH\;.)[ZgPYa.E\E#?5bbQ<SP>d_R/+W-PPd2gWB.fIf[W;9)0A4Yd[
;X9QC+:V2V,a&,Cd1VdS+3^A(d<4+Q&/+F_JZ357fF]6]gC;XOAVNR+&Ybfe_B<Z
a)\be^(cMG-]>A)9QG/M59<YX/)+=#^7OC?+[=gYe@dS/.6<(5=J6PTdK(V;a+6]
85#a,e=&55]Z]FN^YJ[\eZIDI47]B1GAZRA&.bcFHCAPTbC9U2d9PLPU(->W-?,G
K@>c;T\:4fMK?d?GJJSVM3A;5=(?\Oc2:9N#=R6R2,<>V]GTSa=ca:0\F7g@+Pd9
g]fRYb?D](6\cH(@=4Kd.._N3eCNK8+X&K=K,9@d<Z>b>:79-U)&E9-]R6TO58Wd
Y)N\W^A8gLY5IMC8&G[a]9a_Ab_FE6CG&I?4^2.8(,Vc#Za[(dUQ#GG:a[\97&;M
=-WWYU7^AKK_CO.aRSP4K?YOQO,]QG2]MFWSBde:d/],<O#g#gVLKFUW>2G#9g^e
T=D)V2B03_#[/@2WJ0We3QI00Ue7?@#4@.A[X3?RE3;6b:IU-Jc#)Ad6SL>H3b7]
@Y=KB.1=3PJAIJGE_HE>M+PZad0J>a\NX\Jb:1E1[3+X4ITOJRbeeeXCM(gGKLS-
_03N)YeF^S@Le3\PWU+]GS9XFJ>)cTR^U<=8Vcd@UZ@fceOgN?-C&Rc]J:U09UbO
5eZR]cB<5^0b),>/<UQb5c+a90Yd<^ZJd)C@?K+TZ6ZM&P#b)5;eFJLQ?ZKK<8Cd
C[NT=:0[;4NG<fU<^.+C5gZ:=D\QW@M65NMELeI8=Yb+T6A];A]-.+:8W=d:0DYW
G11ULE^?U7O.>012]^>:[0Ree\UgD7cAHb/a)dQWCS&Z3T5SZdLgKKZ\1J&D,1G6
Sa@.5_>,RcKg:L#WO&/T^X3B49[=/V8XB6?CZ:>Pg]H[R8bD1@XP;RLQEM=JS(dA
0<1YSAacQ?2ZeEO<a>RHVF1P.bB;1^2;Mf.B;&62;RTgF0/YH[;4W_:CK->NScCN
84SZDAU//9SKT:FK;)3XAeYJED19P],f^&9G^aTbcBKe^Zb+Q6A>)WH6,:JAb4YP
I]AV4YG#&9gHgW/K\K)FR6W0X[:T=)KIYXCKRI/C0W6X7&K2HZDOZc(a6.c6]A((
cL-^45YgN_gNS(>]XKe5RKW>fC&P<P76T(G[4(dK;g;>:B^M1SA=dbHS.@a1bea,
MYGX_H42YgS[5>KHM0;J<^^1^[1]6Z66QH>(BgU(Z;a]0@+-[U]H9]GgO_?7MZ[S
]?49NI]4&+M=A:XJ3R7c4-e;UFT11BC31KCEUAV./B+\JS3P9D5W\N.J3,R-a<.T
#WP=D0f\T?UZb^)FGfP4&T5>c^<#@bg<:YA>N&^>_N:Z@N&FUVaB9X_)#_.MCPY4
e/1:MJ@4[DNUNGS.HX_[E1TPbZA=NO0UHM\4^\-MI90Y;@:1d=.b0DWC)DY09&/0
eDIeS,1+NM\bTcaAAg;G+-7bL(Q/S0B#]L?6XD?a;;RR#NQK+G0aWI1dc@@HOZP]
..8f.R<S>&I71b=<4eJD9\e3K221fVe>Zg(OU,eOPH7-A2A(OK?a9Je\61e.cAg]
4c/&>bEVBRUR3b)dQU+?ZTTb_^Q&HTL>FV-_P4WIX#DR@4)1I:PT?eSCe7IB.=9-
O+EFW;gDL1-T@-L:EHa>TZ/L[S5ebLDd;(\d+^,d<(4Ec-0#?HP7KTH?H#]AdfRf
DgQ5P&?FO[+MWCCA\@/@1eMK,/K<4[D89XVC&/.0>L[G?f-FP:O)M/eBC?BI@0,T
WY...#SO/Q1XSJ56DD_66#d,;@LR@Wa+@F[><GA]69\H<POH@#3KI(PW1GY(#SFe
EbLJdZ.V0#ZEHHTRMPA)KB?TB_G07W3;T@_R,??N(=_@1@D0IG>#g;QG:T63?LMe
],+Nb7#=J8J5HPY.aD7CK_DeOe3e9/YG\4/C;[d\G4cXgI2f(gZfWE^_3#Md]f0D
9caNWK@-FK(00c+55R[MaKVF>e=LC^1A,e:+QaX^^QG:BC2Y63,g8R,.)VT@/e;-
_=DPOJa0HX^b37,KD>+cY[9=^@R=SD?K-c#^A-WUg/,[475FUMFc5?#S2aVMF\(D
)^eVN.IA5R2//d[JM<QDEgXI2Ld;EP@-TUXHCCa/VG+ENUOYcf5B);,0K,9GOTcD
3775?K<>&,1=??_HNVZ3^@139cdKJ4_V?\7NCWd,?gC]eHK_IDH,JZC24ef6\)&>
A2IK-B3Q)N0SA<2>4YGGfU,<2(O]?]1\0_?b6RO2/JEadYTFJ+X#HXXZ9G[,L;PS
KPc?X&#F5W7-&U?Ud1(O7U2&.PAF6M<)5B:(#5ObMAJ&73^PNB,[Y/W;?e=I_91N
UIf(>D_08H??Ke#DLRNEM8=V92LgCX\3c4D6PdN^O_W3#NY0,+X<;676M1K9(VQ-
G^\DVLd>582OM5gQI;Y_:-Y_\SL&B[7+Z;M.,]628E,_f^T6^8P0<K];R,H(96T+
Y.VMgg@78aJAU#ZI8WE78RQI>5_SBW3BK(36YbNUI=A@<Q#^1>2(fGeb#Ug-;;Y5
9Y2HSV;O>W;DP:CZG0I?51:F@A^X#J;/XQbOJ<OgQ-SB6c1)LK:YI:OPI1@OAZF;
ETgH=+,c;OY8/gYS=>V+DS;4&=05=\Y=,.OQ:O\-De@RbB+FUOUM),89[AG,<UQ0
\@)K6QPOFdK7<XC-?:7-T_\P@37S)78I2]S&B5H6F,7@6^X?X=&Q-7.XQ<L0]OIJ
1NHH+.J.d=bcWXa.AUSO&?gUg<ZD7G+:XfCL&2C(C^M4UF]T3c1DENP5OCf>E79[
>)QYB@^IO2C)H(D6CG2;/D8E4,afR=D2T<Z47/NY7>R=A<QC62:,5;\93:.GI:N)
P,B7AHEH/6:0<I,)ST18>JNR4-69VCJ,=:0W?ZV0(^fLDdP39fWaG4ZCg37,@C)F
PcK&HE\f7:;CeSG6[2JHO&6)<UGG,(Cc]?UPCN+?-[G2+S0N&eB2R;.U6NBYA2&.
S,25I&Z1/a=F\,PEeaHF,EH7BP1[;=H9G?PFR8bZ<3.CWXP213^GIZ;WU8V;a9C0
.H=@KH6]L\94b&V:9fPdUC3V9DF@DZ\^#Dbd6a4\+5d?IF>:3@71eDF<)VP0.8c5
>:YC@()0]\J.>Bb<EZSO&,8)egbXZA0ET5\B(@#.Gd7J32)MT4YWVL4f,4==?Kgf
ZPFU1>;#TD_5U^<Ff7bIg;XD+6/&>?3JMD(QX9P44FPT\7)@/++,8c+e[e0TX15Q
d1Z2dDgXOFL+8M<4]TGN4#8G+K6H)GeFb4#T0HfE-)@F\gG/78[.2PJH+2(#JB5-
>)34._8C5HgGJUd1#8bG:Eb<J?KJ&[\+S14CWDK1\4485=G/3D9MfRc7ZgP>,O5>
\B@^3C^+HB)P2P_37I(1bC7MV5[M6W6A1SOPAUP^J@^aYHVL1JYLPaK:):>]26&1
U.V@f@AA2=IL,G9f&cJ^(=5PO]YT</&a<DZLD#M#^G-0H13Y(H]LAN[.SA\:+)73
ORET;\=@E>BZE#^+3HPdV/#fJZKe+]JC-0[F?L#G9GCLARTS3P3^MNA4N.;>@g+f
G\[?)MF@X#_>cY3-XA2NR=S2]<@0/,^^AV\eB;:X5C;P<B^+R?a?X7?83E&f@T=+
A8,fB>?I/D+,fbPZ@b#@(,JC,)JKbaQ3;4L6B#ZA,N1<GJ:?a)/CW:e[Na/LFA>S
eA=6?gPF^K@d,.Q3_HR8IN1N5+CI[IQNNR,#e+R9Lc,QYBFO;[,1Y1eWYS1Y-H[#
^R\T)eP&DUgI]M@__Y8.\#[?0NXAK(<FVV@9AH->cPaC5YgN6KMDEJ3M10b;WD_A
U7]=bAJ_c=+@RBUOQ[VDS77^+@+/&SVeVb?4=I(C,+1X1,R+f\5LN.LN[/LYecXL
HRPUU3WSI).TJ3a9BB1?G[G.;=e8S3(?d8g51.=GMg^[13P=U&@Q43Kdc&?.X9);
W^1KX1&9Nb+f=(6WaI?[J/J\G7bH:OGI<_1^.SYe7@f9N>V1(.3>NK&UL/VWOZe6
+b\Q/39SdAIbD_R_/[P[Bg:c6aS+)?c#LIc25VD<KKJQ84g8=e[e+IYae@]74HQ?
_TAg<FVIdV2;8NGC-Y3GP,@5L:dbQ9;Z7706eT_WSJ+cTM-:9H\<:Ng4[OfI/:]9
+E5AOf:e@ge_Ab=a_QJ[M752[3N++M@DFQCbQV3beD(#dZ(URYWG2d\34J:NYX#I
5S&A=PfTS.#60-@P6TWYG#Q@==2MAd;,[A</TPU=0=8J:L>(/(Q_aI3YN+SPB1YJ
&-PWHVG]_KZ5Z#16/MgJ/Ea](f4<F4>)53.]R,<G-4,O/4,7AaQ0N4^JMFCN_CHL
#QOa1HRM7)GCD<#W(4K3]BB88G#)>T3HQcMGITHZJGEQN1#0<ddaARH#)fcd\+aV
\T;N:AW6=&^Y]4-]=cBWR.2LTd(Zc_EC?_ePZOS>eAPZFKS^a^U6_-F@/FLEJAN<
8#cCJ@;:US.K]EKG[dI,,I._K;g_)L?)=>^7R)>90457\A.S2ZW\>_V^ELL<KV)\
.1L[LYAYW1R/(\dV#V5^X8B#:f<YY-3JKLfCd0VW__C)E,YER1/M4W)N;F1A36_6
]eS^0KBRW0G^?A.bY)[7FA2^HFG8_&@#3C1MV#S##7SfA0,SBK,c2HRE>L#QM80D
:C6+1=PVMP(eYZ24PHI&A,W;PEA[d;eBd^-9@\6EVT;_[f>JZE+=69(5AN;5X,WH
_K7@<Y6VVg9IZc?C;LV-f#8T=/aMH6d8>,WQ8(&]ADg:0(#J4(CG3-f)R/<O+:eY
I8RUJ[05LUg2-/]_f&^Vd4MfM-]GS>ILGH&_d4(DS<0?/=+EB&FdWg(&>D=+0T>7
(c(2TWP;Ge4B51BOE5_]]0E:;b(Yca^BQN>;R_dI.>YTQ(_]7cb.>XBa&DD,BGH;
;[XLPD><MTA;R(@.HIf_J>77fQ..;b^[3[L9N=MP?Y;,c>,Mg04.=g/WG/U2U,ae
<.N]2\1<He6;ZU\b2)2T2<L0fd_bSY[12;<.MB;1831QF:D=.I07YVB1S/C-QbFY
6+gK=^F=TY_YU&Of(]f#1fEM99bEOe38HC;I#25IK][;0V>&@ZM@@<Y7LX1.E^WR
L/:7S4<^dZPM8gCE\:8&7Z6_V7_;T>?&X0>;a=gc^BYHAQ.&(DFb)48gQB:.a.--
@X)G0+,UdcV4HD.JC[:5:N=7\BOIXPN6f)@ST^V68D9YWc6c.Z,(cQfIG@J7U-T;
/CJ+[Sf=]Ecg9J.:NE46:IRG6=-ZRO=T/(N&\>2O1<LSV-BZ,A8J>#R6RN3RKBNM
P,@8_IEPb]b6J)AY:VT,(8?T(Fg6/()3/8:#^:g[5ZK2TK2ACa>g_a^N2b]O_cR5
F-Tf?cL((^K\e^FKC+:#GNgLMMf[7GI/,3N-]_HL_370@aZV.O^U,3-/AN>f<M+#
\1UB.(SU<\GODWP)F&;6#fJM0S_&a_P[d.2J1@MYZ&X>_ZHPbQ_.+QC]BW,J.<Ec
6G)BF[A=+@\f:PM(RE(NGFV22BHV:O/;9c4PV:[c&R<C,:bbO1[Z2VWdVE5EFIbA
CD#6U<)a]\]?D5R>:LRF:HS#.>2Y;29KOV-Y=ZOX9Q^81_&Q.RR6P#HEdCdV4b(d
S;]WePIX\@A\@^e93cdB@[d]>We=:K2B=e_5K)G\;/<^fb9OV##K&Nb:V]/-E]3?
C/R3.W7S_RGeZB.(LN/c&,_edVSFW7M#MQfPO_GWV07KHKLW9aPY_g;d[[A56cNK
Z8aL5aK#dVEc5A7e6<^I8g@^2?gJeL:<-ERJ);F@KQB+>SR\@L_BQKIYa=@c@4F4
.;R/4V9.,0FJ]3N\X#S1P><d5ZU-C&S<f#9/&/#KV\b[>(#8\SI1<+0M;ECa)4<:
<I\6DAI\Y-_B9-Y[ZDcbc+9LfS7NOX]W[eD;SR:21<81HQ&dRb-S7E5P&91Q[+9Z
Ba,9&_LJ;,I1@YFV68QO(/<RQANN;LA9J?;eP9=3)2>?/g(7f(-c=fEI&;ZgKK9T
&>?Fbd(e#cMC)L1I4&VL>_fg9AGb0C6K=BXW:JUP.@/CUaTcB:#:XaG4cG#f(H,N
5@I?dXd:fM)d)NNTfY;cRC8_WfUNBZ+e3+N)0D5.8-61@Y[0RWg;(0_FW5#T>NOS
SRSF=J:D+PMg>&N\@SH+SFSb67C:=a]S,].&?&NN1+2+=+W.=^+);eFJS/2+=VR0
+<OJG[ECQOFR1I[XJET?Z)?Y:09H.]Zg;E&g/S()LR^NI#@VIa9&J9O=>3,2#TcR
[1@FG0YcHI^N_K-e(86N97H.5dB1L[N1CHb0Hb7#Q5Y6=J.J@V0@cX:))c8X\=dG
E_3C+Q)IdQ/@)QB=bB?Pe+7E,W&fI.N9/.KP>B\=LVR0_N>5I/-23S<O)ZGUN2:.
?L2+&5WW7,ge^I/A.&S+0]6)AZW/Y;3)NO]XK.K/D7B4/T8c=VgJSYfgW[Bc3B0Q
IU_77DYHBZ<WPLD3fM)8HH6@27X+TWD;3OZ7^/,8-9YBZ1103A(=^[K96)O:-,/(
9=3HSbQ/ECfFV(7SN5[LFe@,W=3T((+LQ\[IUC8cZ^HEbb7>]@K&R_\FGg#&8CQ4
;MB?VaNM<TNEfbZRS>Le\c<d(&IX5CCBMZQW1#E,-\g3D9.GUg):13QeF5ed5b6?
T2U4d:_QJBY&I#/^PbS>[6aPQEW:7,C[9[Jf5PG,/&8N.-QO]Zb;:O1KKd=fLYY-
KHIEEEa#Wa;XB5TY/Wf_L:4&W:fgE3eV@,IG&0bV-?)GUJH+B@MOA?R)4(O=]UL>
^Y8Q5=F6+A<@:/1@KH:2KV[R)41,8:F9&::[5&ILSJ:-^Ne;&(aFV)FGYFHaX]I+
DJ=5-9I<H8>JL+b:)8Z>aV+FaF)O/fbXQ45cUJA[\DA5M-)Yc7OIH=[]75]Ba1(.
gN4Q+JD,NZ=_BV0(_a[5H4KZC^7b&=++f]7,PETZ<^Y6,S27M-/f0/=^J^/cSOX=
#7&dD_\:U09dM?<8S[=@]eFIO=]4O,abDcY/];cf7K1W\#724>-I8e?VHBbg0/:0
U>7-(^.IU1N,dZWYZI5>9E&U4J:?.dTC=B.I9N:Wg8a=Oe9/?0NgYY_O;Ze9V:M#
FW99=&>2(6,V.\GSFa3[))KBEADaTbOO#M,3H?^E.(W_[EOC1&89]Z>5R600,F.Q
LKGS+La:bF^YP9GGd(3:Y5RP\<0;1TYP_VfK-F<6fbB0)JAX(76J=&2&#[[#44A<
d./.Z-RXH3J-&W8J+I,S=T1;0V>FN#+),07=8Z,RG#(DEddB797NIB5BP10;JbZO
abgUGe\6F.6SdZY45LPH.Zb@1OFAaF;94MaaaED)B,&.0-f\EW85ZgE/XJg4HT-\
NfaRJA4^U+&WLJJC#GS[G:OK])IBF(b\,\9cF=EbSbZVI:@#VX3MdSLa&/,I.c8M
XcQc]9SWC/<Sg+L^Z1[dU-::</+/MOS0@<NLSGF\A_3\1@#=AfPac-\A[?X+9V7P
?696GBX.Ggc(c&=-cDE(SMDK+>ZT7ZWB:L9;(E27CF?-6+[Gg)@Xe/?;_51D@N\(
d8M&JDGeB@GPPaQ_P?cagbCGW[=+Lg\>GGb0,9K1b_G^KbZ#LF2)gCBK&&MO8V++
5-T+G\cYd#-,1QPRD>]WQ7-OXGL4EN>RS_==F(I8O7Q3L#TU;3g0;Ed]4M5V5D,Q
,8G)G=R->E9Y]-^^(^0g[.2E<b3FS8CWHM+514?^3V^aB5)88FV_2&+\,8/L0/6A
c;6)X;^-6@6Gf<;[9Z^-BQF28:H?,gQ[-./-Z3VLY=,Ma:P\S)<?(^dC2g40<;7)
&-UJAO,LbERe<RH0<P\AEVGeA^7J2f6IYfHGgg]0R?@7H:I-TV><7d>#W?F&;aHK
:IT^1YPJNd5d+8T<Ue/gLJWZKY5Y8Zc^1ASZ?(JeZgS&?6S/bgec)Q>R^DGR#)bJ
O[AF#JCd(R#,[_\VX#Z1<M:5+_V56W1R7_#>/A_5bL))#\M&(R(077KcDegAFZ?d
>ff@aLbPM77P_FM54G<Ke\,H-V54Q;fRN/Z&NZ\[Ug41e]D.<+ff_d<LTZD2fbDV
;YQ:XV3Dc8:PZM=-AEP5L-ZPTHOBg.)PcB:YOM290?(KJI-9[ce@(-)3^T)=JI\b
F5;GQBb;0;UE6K]E;Q/>#W^JBVNQgF88(Tg<\fWV2X@@6V^^IK^We9F]JRFUDX>e
.:&Jcb-0#B)6BSYFNT5VBA56Q@D4AAESV.,<_fO&CBJVXb[cMQ^6P16IR:fI?6+e
FXVb=3H(@Bc;=_HY510Ug^NU-L:\]OKdEZ\CM>CL2XOU=+C<(66;H7.E9Ua^#_]E
^+#S[<O<AEef#\Wgf+[GVCaPOPZNfKK3\(?(O/XLfA5U4,A((/^@Q?XBN,SX2=I:
BJP4=YQ+8)V>aV05QHA?5UCc.DFC5EA];G.;3Rc8T,QaMcT.9NG_.YMN^8CdO\DC
2>-PN3bW?0c>a+B<7((331U_NcD1@^X;_L6W<J=G(;fD]VCgKg]C[8CFJc9Kd9OY
A4EI=3g/A\H8T@:/Ec>;Kg@30#La-Nff=G0(B94W;3-2ZgP&ZLg;R30/_Z<=BS0E
f0^1^D)X+.?N.D8e;^4dCE@Z:NP+6.:Kb8Z;++C3/Ec@fXK0^=KDRMGJX2YY0FY@
C?^F<g2@:b)OR66\D@45NcA\67DWc_@6T>+MQ@+UFeS2>eGTWL4.QX]77C<d(9T^
XZO#D9AKJ_Yd,?cg7=ea,af]78M+g)@XO1McX]D.\.,YLZP\0@eO<>DDSR>JIWS:
]TA=8/PfSTNWf85dGe+X;^?Y+^EGETb.8T2AXKJU^+-@&_#0;[+Saa/W.QP,EAb+
FAY?7Dde@0\]>:b^2-.K@RXE0U&270S3cR3a#X_CUPgI?GJM)3IA_,cCg1dDR_BK
.8\R7&a?,E(V7FXG[,5C\_^O./ZgE]\\U]<cW1?TDgY2=YR,adQ[R1/3J<PK_0R?
DL3F?M(<)3Ug>9d)JSKWR,)]TQ]5T.KWX/Q1CHM0=2;b[9RMVH_6a^#TbgJV-:K(
Xg>#I]d<A=SdEc\=/TL=<CK;MUHMM[.^[3+XV/),f.-8SFP6.PaNI[0(;70,]J)R
HQ-LLRbYMU3-eC.L-9ZJ.6521S-c=7Ue?]^1<C8(#Wf:3?1=M@2QNaCM^N6.&7c>
6I5\_eD,ef83]T,&C:13V8(&93G1gG313VCZ-+@dBI/7+:X(cfEI1a1,7W]M9_d?
Q2D/PVbJ2L36C#?IG3D8UK_H#(Y_08@LJ=d>LXBT]#_-\EYZ@9CY1G7/eGDSaWS\
Kb.)bNf^_Ob?2\UGP)TG60NU(HLLJ@&8:5J@0cJfVY>^W5)H_JBD&#OF6,L(fCcH
_g@C.2B)<cKZUGS;CJ]d#X8[]RZFXU@c>_WL/P,)\_<bFBAIb]E14bRN=(V,?[BW
Z>O1:dB\=C-PdSUBF,P@Z5A>3C--K\?SYM:.:RfYP]cO/WO?<#\dJGfZ5]@6>]2A
DCK\+AM490Ua=2J+:8F]RD5MS1@0M?QKeLY+OQ2Gd[]dXL6WWg9g<8AZ0C>=2:RP
5XZW#B<4EfJ:(_ZT:bE_]Hg;2PDDW?I^Hg\@RH8LQI4M:eZg/[3P7C8HbW&W>A<W
VU46=?[Baf\c\If]GPW0_4595I2Df)VP=d:+IY]\6-UZWa8>H7:+2;C&Tdd9MSNI
g<\6+SW9ME[@XB_\]RW,&8Y:5BZHMgSJ4eUQgXHWH0aMZBD5->^LO_f;(8=gAP59
a?N\gD0]MYADW]:;c7[N#EFC,C1\S2[GDOY\VGe8<;:0Y7#Lf7XJ=RTg;/MFZ4B6
deGTe0500FEZ\K@[GP_?PDS>,GA_R72JCPV;-\?URO^4Fb;K>Z(^6K\Zf2ZS/MAZ
-98d\]L?0gH.A,E3/K;>5Y7S_5,VK][SMW:P;P6YK9\0[DdJ).PGOO/U.ea<3Pb:
@Jgc<Y1.Y[6KQ+S2aAA(O25:^H&dOa2?#U?3V4=0/LGOIfP9DNE_?9c@6Eg,3NDG
:<8g@XPK\3@G:aY0&)=?[UHC(6f_cHR9a\@L81@DcQYf0]\g3?9JO.(#_4?AgR.d
#1AQROH8ZGOUfK2]#U2COg;O=\K-eIfe?]0,3]g[?OY&(bD[([01c8V>\&VggYfP
9RLbOaH2JLDWERf\P:=.+\Vd#)R^<G&PS7>)YA[_31b-c#9KX?D_c@3H#NH@fP=(
ZY1T.RgE<42cPYF;S669XeC)0g14bL<ILYU:SM;&-Gg2D,gIaC3P^eY:^<99I#DE
2Te-<UBN;f;9=&32]0+36:1OY6?Z6I>f=aZX-3PT/YQST_9665?-0Y@V:5(N?fG]
Qe)AK^3;N6]2WbE.:cUee:UWQ;8cS2&[cPP0K3bg2UOEe/Y>b1<Y+/b1CLg45bS[
;bFVC5YQK?8^9,CNB.fYOT4.Vf,:Tb\aUNF&9WM5,<K<4)8G_e0ZOG=<EGRMeGg>
Fgb7F:FWHS]UY^LVfcSYA-Y9Cb>a]KGWW&)Pg?YCcb3&<CgB?Ad<^19K?:d_[[=L
(/>JFA(DVe+#H5(B@4YZI<\S3V]:0[OC6?,^_RcaHON9#g^>)1>,e\LbX3b#NOM>
\gP.VDJAMCY96@=2M#(dK\@++QgDHMSDMBJ>,4_eCa[XWI4#?/Z=0[>[TL0=He7.
Q6UT3BCbT>O7G8geG5\B3^2W3GQGEUD,3;WKg)DZ&<cF7(+6L3AeC,dJ9TP]UG1f
>CQ#H9I8.>GG6D+I,?7SA.O:dSJ>2c#f:FV]4KC0YK.7[<X?5VN;<#13MHfb5g(d
]84ZX=BEG^V/B.6@[W8f<&&PFE\@?V<e6NA@g;O9OF)eCA;:8BRO&OA1/?:FWf>7
4N.bTgI)LaH_J,SBWR_,Nadb3\^P0-(5KC[(4(=g_>F?^#+W1:/9gL8+40(gS</B
)Q)=R#AOQK3K9\C#K_/(?1;b2T2fgH2g>^L#,;SS-d_&W0_U5>9DXI6P]K-],7bV
a3;,(X<AB+TJ_Z?7\ee3R5J[#.OF,A[@M\R5NCDEQN(/)3+fYJDcPBBYa>7cdR4J
XH,DC)C1/IYb6&?(4:L>@>8AMa&4#L/,G36B1]+-G0FTJU9Gb.+P9&FF)F^@B:&G
9<4(.AgUV;JJL:ITcK).E8C(.@_gZ;./\]GQ(6@CI=T0ed2W-80<5&QaRa]G8.]P
U)D\G=]cdY[8e0->UIN/aV:<W-Qf28/[_./+\WO[Q_VO2AW48Y,JXN&3,A=AZMP)
./@eEB;,(A4Hgb<]U:7gF_cJ(/)9=,]/e9f[\OT51H_a(KFDACMe53^TFL#gJPG<
L@AG,&R_B<6;Z2K,MDR+Sb0JNd3^84,9=687XHBWTS)<=81U<CH@I+U?GSH5LUU]
1]4dES0<gFSJ2W__CH5VR5]IfMc#/IfA=J>&DR/CW:>;2C+Z^/[O/.8eW-\UB5,0
#;:FAZ(/US;/LMD4F6;L?ZTG?-,N\WBI#4^FL7R@?-&M@LKS(T3[&W?\<@b\+f5b
a+CW;.D-PJ9K^?B@_8c)UHAdTOYAE3\Q+fOeb@,.2(dAJ7,e221T;g7WL+WW5aI2
>4e\ELF8N09?J9[G9T2cd^@G3Y>9YT(;N]1L/f7PU7:.f75.T,]WUA]?ROA:=<2&
R2JMB/GIbNAg[+.QIUWU--&F9F;N]#]0]CEWJd3J&XO-L/eY\#H(G1(_66e@F\50
Lc)XaT?MOD3.>R/O>@:\^JBABIWKLML@G5><)S^_N8;&M.>?O+1.D8M@=C5gQ)AF
FI0W#Og&]07>/VL<2PZU&0RHSH_.Zc.50,X\0G^NcN@K(c>@+1/>5VIPWY=_N.#Y
M1Y=g0@DBAHDX#_56]8KdUT:c=Y.M?0##)/IK=7U(Q9XQ>K(<BM_QNIGSA6\9WbY
gOJSd<HYNTBKCV-FdfD-aJ(?.D\^LCFTTSP6F;.#5DGB201-:&VX3Yb=fY#ADWDF
Q^)AWH)-WBee@\V:C+Kg37LMRZKR:(VFf0DH7^TdM8C,9\gN+,Wd71EQ_6S=EHI[
8@,Za/@\&fU7+==B6dNBZZJ\O;;FJe5V?I_[M5b/>-W3.^2QaJY];B1D^CZ?C<OP
@WDFc._^[JUaQBcbYe5LcI^XOG0_[,bVYVa;Y:AYG))R80VD&cA&(YN?<cQ3E-=S
@LKA^Y,)/8+O]>Z/O3L0&W2?<0FY,9aBYK.-d^Y)SA.gJ1Y(fHBA0PG)Q#9066#V
19N^D]?FRU^VK6[^50=RA/8KMV/<0X8@R<Pb@MX=FAR\>/P2+?S0;71\/T0H<DPV
,8?.aF;]]FI<+25VE57#+05V(#daOR5UG.(L2)Pbd[6>K[F,\\G\^V3_5<=ed28D
@_\Wc&Ud?aH?354)FVP&F?@A?47DP2E#-=60&f=1=g8^2/#JE&:F[67&]/,NJOJ0
7]JC)#[QYf_/:M6O_KQbWfBSc(\Yb(LR[;782J:@(:1DN==[W[e[?PZ(HLJSdFC@
DbdW5]eD,]?+:KOSVCbfZNK)[L5+/8Q)(+Q<U&J_-.P<S#A-ScJ2R/BT(:8<ZS2/
#.^R[NNZ)XZJ&IRe8aB/4NOV8/V5@5(-8gg8aJ#TB^S97,V<bZ+>c8,_18_GRXCD
>&Q0Lb#Z#,?B@=+A-_8;;e6,gY^.[C58W,#eEPf3a8dDJ>QV<&#E=dXbW;@bA2c0
<N:L&LEP;gA9[4+/=Y-_12?IC>KgO@EM5YbcG)<_=O@S^]21[VFLAP9I?W0K<+Mf
,?I?B81>9&0\C[HU.D^&dDF9_QB1>C4B,fQdL&PICU8aT#c>DSd1KC12)Q7N6AMX
^1[TS3JcTBV<<^JfOJEJ<#3=K0#+\4Z^gcN:R@<\c+dgbg8bL9a=N3R;2SE2EL-U
#f@8.1>eB\=:>..+E,7;72dS20,>e.+BYTA]1TH?(10MEE1=bAQ9O=C&f2LBR&P+
.GQGZ6Z\5IeP>Ae@Z(LZbM&Y>>YOG:a6f//_P.bS^@LFAW2NC=HfJP+H>.HND@R,
8&.?Me\@Z=ULUTe66AfE#5fB+LV^S30V6E.&O_6(R6<L2M<5L\1,45GDL>EWcaL\
HR4>[_7;=ZN3\@88E.J/OQ;=MfYR]2OG1@d\ZU6J<ZS/Bc8EUC+[/8ggY6R+_<+5
S/UZ9gWUA]W>Bd+ZHMF0F8A,HWf^JR@T)[:OY\VKd7T#Q3M>ZAXQ;g>-ddg]R-]1
/4dF<^4Ja2U4T8H]Zf_/?R_N4L7:2eZfS22>JA,E>H.cZE6gKM\CS:ZH._e/6BMT
3V2;Y]SCB6Ad>aGSKFLcKXN2/)e)48M\TZ7MY3HKdXbdU>;6]^\&V)fCO/OPH=cF
Y./DE5;6Q2@bfIFdRR_SX5M]QZe?_8LXQ9P^AVbM68VcHaX:;^6_0?_S^@RN;9([
0F:\eIa4:AL^9Sg]g?2>HB;F649IL131>R.\^1?0+BW)M<5)QI]Z+CZC[\.>T<5g
@.2WMaaPd#B9a(VWJbANC@:ZbQW,W,?-NRb)IHB9#<;(DFcR)=g^Wc3X=UFA\-QP
_T:;;(4NO]?#:4M;H1CZEg>CH,4I,-):]dM]3897?AUY[F5#1J]XQ_;62bZLGObX
4IaF2/JTHQTD]eM?S9/Y[<O0(DI9--[KCN4?:M0,b-T7CW<b0N2Z2CA9f<;C)&N]
;^2aD<f>K7SB)HAcUGJ.Z.Dd)_U/=AfLM\b&Nc-DHH&aL:QdT_,PZ,P>gD3bX@-I
MA31Kc_YLERH;;>L_M))_3C+,>6-@0B3WDC_7HFRN1]HF0N[/cXLRMS,>-WbgQC5
]2W.6>NZC-7LYST/4^>/IL.=4f<PfCQ4,T5NEC7^]C@Ef4B:O8^P3Y:2De+Pe)12
)7G^]R4T8AMd3M;C9@0AccJ2I;D(aP1,S9.2AeNKQ?S:U<EC7<#S,_[aOO^;AaHX
1A>O>&60Kae?<7R+?=?fdT46I[@+Z?F4YOF=:GR4(cF0g^;LC?G-F533:EL#]I2g
^YOB)^)bFND_N:8U37Z&\:0?_.5I_?_04#?F[LdAIXXc\OP+V>\W_[S^RDFGaAZS
_P6H\\NHB4H&,I#SV,:b_cPAM45#S>X;<BE?,6Qa/+c1;X)M][[2[WG,S@=<MM>)
b2C>cNLMA2^D9]LFP>Q2@0&KecW:)9RfNaF]+a<OQ01bMH(<5Icg^J3S2QBLJAE1
ZV4JM61#L.8CSY&=HGM8^UTAa_K)K>cXdPg0H9#/@G?7][DSC_7H_:YPPCV;BaLa
cB6VQMGd4[R9Ye2W1BXS7BG-HbIM+XQA>@N-(IGZ3gQa(W^+?1I3XR(?3PF9agB+
UMVHCI>IKQ(Z:H&@&.BAF0N,:@QV7>1S64Mca,IVP]O0C#D[IPT5]-WAT#f3Rb)d
U;D]2-J001PS)GWVGM.Z&3V(_7^_Z/.9NCO4ZAKB:FKHWOEY\F6?O\@:W-;1bWLW
HfWXV=3X<gIDO>CdF>6HNeL:8b9Jc?5a5Y\EAFgC9P0M<D3HG__fJ>?Rf59@1@T@
<Xc]:)Mc5g(R83JE@03&gZ>8+V>AEKFREId?0RE4\-3PQJYSOK,7eQ::Dd(5MV_5
SIYI1B3V2AB>L316Q<dPS)4KVWbga?b0[MAFKJ;:-./#,EHK+RH57cN,Ia>.NRYK
?J[B[4TB#\\]=+<ULH2GeW/@<)KJ69<^U\Y2g73R[Cg2G7f[F__SF)f8>YH)6JP?
702\#LC/G+[T#E#Nb&gZ<ZM(GYZ@DR3Qe6/ce2CFF;0RZ+&F:M/)QKKacYIY:WO]
OJ1=,e.XIdA#gAg)eZC&)J-.29D+A2NF>=]N15/?2eC8S<A,f6;V1)cT6CJB&JVS
,6<]DS#bCO&QbgDQ1U?N5A/V/;Y6CSGN&UTLa,H56_PH]db4YR>GKggQRT@66Y[F
AA#5NAAA9\QA/FND<ZFXbNVXf,,W/e+HQK]URYYY61^?5SZM;;9[56@4NFM7=GdK
Wf-3PQ_?#+b/WSDa0[)dI8G4162JLbDL-I?U-1QQ#]-,]4c<b8YGWO-RJg?0/^_G
TN9E<@3QA]A_8Z<>:2f)^,4dBOC+ZKg_HSR^\cD5PG2[JR<Z?4<@N0S(IU]0MeFK
^86c_/?DP<UJ)L9,[TGa9.=4<Nf]E1W2NMHLXXYde]A/d^..J32Y4ae9d0V)]YTI
EcPANSMZWV>V7cI[QN\UU;/@JC98RUc7L(HK,C[K:+ceJ2Uc7TccINY#e(7XZ;K#
/P\R[[cR@TFdQ>.c@[NCT26e2+1+ZT2dDYC(Q67bM/96(+c5@([Q3BA/H><Sa-dK
eEY[N\0c&_?(<V-f?cC&N>#f^3MBd:Y+I#1?+33(94I9f5];H,Z4/@dUST34[BII
7&4P(,.Yb5ZREO[fgE7U71\9@2NL_<0T1C)9F\[]FG#HZ;>HE2/UecH50H4gTY1E
;fN@PYHM)ZL2PNAO69gGO&G_W;59X\-RQJO360EcegF<</c\SO6AAK+6<8?\V(@:
\AC5\KH3R5-#_6DP)KbbV,Q9LHf3cGbfUfcHX26OL:gHJI=eI@OgdTEEeW&gKdCO
91<M[57gRD#SNJ]VFF3>,G#M9gH;Q5+5&C&ZP05=dIc,a+7:PB#Ia9@N_6_8(;&;
?.V1]AVEJRI>g8<GQCaZ>,]T;0Ze3/,HKJ1>NUab,YWJZ6)@?,4O:0@E:NJE@Q_:
-\2BC]4#@/,3D6:#2\P[FA)/#]7#2Rc;[HdLCIQV\1Rfa+JIfZ/R-0<5;JdNeYdC
?C]R<>F46=cJ/+BND<0?2JG&WfDgMJZOLNU6?(eWOaS9R+E;XWK-ZL/a0Q+?-ZQ>
ZbVXacGgfdHL<:cFW.6[@_Bc5LCOX&^@+,KP;-CGYA^QJ^BeZ2<-4FVEHbK=dBV/
PW>8WUWQ3H](92+K^eN(ZLdMFGdg2/0#gc37\?=UAZOM?VCES,TbM&M:)g/J1)AZ
[5:]S6dL?(^YX6L+J#WEU+16YAG3P8Q;QF(c9LTS3-_3NAOK+\:-1V<F.S=?WB>5
c&NMOY[b=g70e_gE?&(>8Td)E(,Zd/C>@?.4U-W>\\?C.)b,_:EN8<9aND#Ybg<#
<\V8T<N;P]/-J-gJ_?=CWVSOdEc]g@S[X]^Qe&WFg<RA0651LOG?L0:.SSU,g,:V
69Z/YY+O)[>3C;J7P5:B5/ZJ_gJ3TB&)L7;&+?Vc;+c&#)S46=P\g4J<BP8>0KfJ
.=Z0X#eM)e<@^8e([OFa(Z)]3&?4QDfJYD1Q\X&=e&(MdYZfCM6IK,DR>J#)RT)Z
DRL#M_PI3<_;^5:?08TQR59>6J(?J3<1VF8.g@=b80K^WD/6KfOJ[(TP8TLN=#QD
A77AV9YEb7&4B:E111PN.[WI;G/+/CH8Df(#Vfdd\.>0W;b9_^ORBMI1Sc\cC5<.
)\[(b[M5+,)/N)TT:<QdS5c#AXP=^_51T/5VWR+14FD57+9#c)-<Rg:#LB8-^[VQ
EKegaVT_-3/AX5f6g/M)MU)QF\Z=)KOU:(4R8C+++F;AHdQ/)@6@^,48aPSX_O6/
\HJ?-+H0T6Rb=QM(B2d(L\B+\JQdN0Lc_\:EO=3Y<#.A#0E=K+QK+Y8CPT:P1+08
ME21H(52A?6,)a;#/D55JbN?fH_N0QAP0cZLQ)DC=Bg-+T1298-MY[Se@HY@I\a+
Dd(AY(;g=d7LWa1H[@[5H)-6ePVb2VgOf^c2VB_)37dVIW[fNZ63a]+4Xc>9+Z)I
bY?A6=;cY9_GHW\[1>M/V.a4?;QAf.XJWV#9Yg>5VYWG@V:-Ge>Hg8WWA,[O]c3Y
2I/d1XD.b8]Z[#bTUIUW=UGaU0+_3&=))I/#Ldc64d70c3B/Z+bL]<b58JFI:g1E
DS>LP<RG9Wb&2)?I+E3/04<>A>7Uac1.ZbF3WP^W&JHSUW2g/-]@F@RXHYU(DU=C
0LMHCLWY9_A-N>L=I1/C+S2EN,(_1W+KSL8(>X=\_K[L+A-#)+G>[E.AFHAJ_b^C
f(b^NM8=<(\Ff9J&bZ7KR^L;cFG.TO>(80UEBB177V9dQaMb9L<:T3S^?[A8&5X6
2^-]9.5Y2O9I(5DAf<91?7=a0JY.Eg4?K.N294]+.LMXgPT313K4K^FMbEb^XX;g
LHZT81B#,4g@:ZJS\#L:N[4aM5_4-@B=</PUML8SE<#=g(KA83SU(P&9bMFO4f0#
+ANF8g5-Q<EVIV99FbJ:AIRT2HMH=?MWHLE5b3EOO#.2=X]8FYGCO&>))(H-P5.E
X<8&#Z<N[=]dUK.EPNUC[-82>&)Ye4(9&>8bbX?0]>VaU]19.I2VJM^27JK_>GD=
,2]]<J14N6FXVA),Ib,6R7_^WCE&ag^76=127Q&:JgS#LKI@J6@8[A()L.S>KU+;
Rab7SXXb1++(17[=8BfBI\A?[>O1<H]<K>##MTE3@U1:13C-=7Xg&/O2C0.P-E=G
S42Ze&SU1O.6XVS=@6M(^b]fRZ_P[.P6JHN@N_&-NY#A5S(-9:H(O]Lcf]:SJ4Le
\26GCDWK06EF6X;^&+fE_Z3NOL#H?gPKg&\L;2:;]2;)M6>93X&aCR>^S/BFS,CQ
1[cJg1?CB/3g+Wg0cZZ>49K;_,/+Y^5-NbfR8Q(=PQ1[9.QK3[SaDaR:BVBW1\FX
dc>fMW/:b)CdJ-7_<TMP^#dd<94;8HJO@_=&FMN0AO@&Pe:+6FV,_caX1A2/4MNM
I7^Y9,#)Y@dIBWXg0@c.MFNUVAGW?4V(D;Y-Kg9>]Mb\(f;#958EJOO5@.Q9RTYc
:6=ROT?^6fV/(LM,,V]B:a2f(Jf[;OSO4K9bKPaA8=b<T?IZ06/3EHDM,>FYd&PQ
1D95RTY[1?P^I\^B66##UUM^d@afdGX,gEN8T08\1Dg2P1RAgcN<dVd=CGPbL,G^
eG48[.G@ZH+[H7EGXeUZDVgC#1V3JZ+LEeGXfZQ9dMT>[]DLXG/XZO<UcO7FI<M?
gD-;^K<93>_12BfQTHGd=,WSbAA,\/d]Cc3(@<L=.#M,\RCO(Q@Y=-N6V:YF:I\e
3O;[K\D]RTcIc\dgcJD\>.b4_,8>[#a4.,B#fJdM?UMbJM-eE?N5[,fdF-E]K6X#
8.DgJ)9)7c3;=ZbJYcMJ0CfLed(Q)J#77JfNbIT5f,X+.2]BV_(EWcUc+G8eR+df
2Z\O-G,+FP9LFX/J9W6g7\Df+4005+#_6EA&Xeg/(<J?:#_4Pc-9b;\V\A>K.[aK
0a\b;IC[FJ-6>&gDc5QZ3TDDcN\K.c3@aX/WXI03]Kc-OT:S#c?5MS[84/><TCC6
C^6f/-^.?g79NVVTZGK_8Zf/KJ1VO(;F.JAbW8G.HEd7_VR8d<3IB_OL2?Bf8cMS
H3THUDX42N03YZH1LV<=&F\(@J>\RfG#YH5L^E\Rf2,&26-B>?IZ+N,D8P62=>M7
,@E#]]MfYOV2dQ9<=>27/:O9?H([:RZ0M?fI-L_U=70dU0N84PN(9N/aMVHNVZf,
[gFW[@Z\.a0/OL5.4[:\fRLb0.d7=-V;,]>[ASS?-NWBX^7LKB,Z);QNC[_gGIeO
JRPL@P,KR&5_&(7VUe+A9J.N:7g0,E7&O1[2Mf3S)WX,Zc4WTBIX?@N9NK,;cc(E
DQD:5fENeX(dXT&T>\3,TWae2G5/YV8,MR>CL?VOTT7&>Qb=[:@;:f,d7IQ.?NJe
:gfSO?<[B^GWag4M^05cJ^KSJDg17RW+=@Q&?e0^I(20B::D63fQ>^/EC(Z+IMD9
6HJ=4E]VBWA=/1A;T715A<#,cZ[B(7aICMWHDP6/N.<E/5:<RZ<NI,U4J^8=aEe;
?+\W@U]J97=^)e04N?&?<8VQF?S>G]98]IQd(MUTEcLLbOb_B0@,TbOPedO4gY;<
G#bJKQW?Idf2C-)A#a7MbAIQ-b5Q?T#bLV3#<=>b2X36))VJS-24G)bL.P83RU\E
cdg:IBPP[LF)=R+ILWO22:S+JX.VcMHEP2c;^?=W=ge<Nd3cVbV&&Sc3?c2-MS@9
/4b34e_.#a>)K#1JbNU0R=B2@=>#)HLW&ACF\]6A8J_&,X11?)-5,]aG58/\54gQ
_@=57A&WPdeW+TA\(f[3c4?.D?1:B&K[XI:.Y50#1,01+T5Mc7F#,YCgK,Fa#^gc
KT=C@1TYV:=?PYZP5VeKFFf8JL;LCbgZ1Y_OR_J0;>14Z2SCBKLZSGFYf:(Ng58a
B)3Q^6C3OI+dMB?a+Q8e5=Y.Y(FHg:LWS:Z+TAS&Yg0,YL/Tg/2^&(f3;64e@\(H
R.HMX4LC.Tb7T;TS.Y>]aYH-CLeM90UNS/c.@Za?cI5E?cFEA+NdIUI>3.W_EKSZ
bfDQ3=:?WT0<39KDVe4daE?#4Z.be<?G7-?>M54?:4BHgPIV?6-N]C;_>5YD(0eK
3Ye=H:+DK,2eCQReA_/>>@e\S_^5dAcCeE@(\131RTN0)\-b>Ea<A=CdObIU][_2
>/VI[H0f-+BN^JeD(Qb6C91ILV&3?P8D;b1_f_7fYSD#?387@bJ.d/Ve3\^)eR&5
AV1&-V:R;;++PI:#@2TTF6b5)P_6/@S4?&YM-+M)BI7M7EKf\A0_Z0<bOH(1Hb#W
T=AXdP39KN/NWc(12X]953:=^:R(@@./JABKfBCc4F&E;SKL=<LR-F+-^g)[(&F<
aBb#[UO1FLCObBO<)f)FJP?3A+9J<d[fd7)20JgK0/HP>4_Y=?87gaCI^2,G;G4Z
fW6[=9OJFC_WJZY#7/YcBEQ,E17-e,(9&L2YbZ[DUULJWIAJ+;G+J&A(6d:35c8+
@eA;Y910O[UHB_2Z>-TZV=(gd5f.NJ3R=FLD\^\8Gc^ZO02M)L6D?,:?UMP7\W.d
C\8-\ZD;4_;].,R,:M6/N)^TM&;^FgDaFS0+JRIQFb[bF-H&KdBAVeFb\^9U(5\c
5J+IQ_:A-8+bf(b>HKFEFS6@.&fcRBNJ=E[,e(Q)[:dJ?\UJ&M1:UM><W0T.HbO9
0(K,#P2?>\XP0F@)5H;ZSN(/;LZ#@g#@W>.2f<5?cM9DNd,@PD8G[9\.8a@a4)<R
VNQSFW_[(;Sg8SFRJ/8bZ9]9+>bF>J]eNY60aaN@XP_XYCQE06G3\5_bD1)MRAN]
79f&38QNAZ_03A,74;HA+Ve:L&7B#a/TR_:?e::?b[\IcO.;bD:YK&Q/+Kg(aJ,X
WP<:Y3<?YS:G-ea_Y4X_9QI?B_cH?ABH(3be<I<3B(VL]a<L\a?DbC:K&<fUXPQU
0B7eba6cP63_8<gAf]J#H5F3G;d(;@a;V_+-Pb#):9(@CZ&M48\_5JB<dP\4B;Y[
G0@31VZ(2^4^ROMQ.U#?B+V=.<S#U9<(1#&[e9V<ITH.Je63-9KHdK-U#[F_KS,K
,4_FQHEQ4LDR6JW^(,7,?cH@T+PeP,R_9@;c82E=-<O0N_]RETU\PUU9S4aaG1(0
R#a+1UK@U3^0LM(.gR]VSHSM+1,F?NcfXE<+d8#]6PB@;^aCXR.>K2C:,5[a(PO#
.<S::#G04K9DC#^SIVXF11VWf#B::?X,^./0<M],\G<P:T,LVDY]8.d#P[.?)0#+
X#=W2:L;.SOFA7_K5b^\U=+\f0B#X^PaRc^M5J\5?a9Z>c^=EQ[UR>&S7G1^9\c-
O4d2AK0TST(B&CfGOA+b(:-Zg>;\G2d8(@RQRg2X:5Q2V76/VU@8g@?7eF;K3e(;
aEac/MH=EaK7.Q0YN_^M<,IC=:X92FGXN.>G?<bV4WZ8>ZWA:W9FH[+DS_,AK.@;
ZQ9B0b;.//O;Q[@:^4K/,B)4229JNW;67@B_UXB2)e\52ac2,DGO#:6):Ab.7H]4
cT-37@.df+2707//afX,T<JF[WFSRD-#9B#P5b5,Z[cDQ&&ecHZ19:8g331.)3/W
T^TE:U>F0SA(=@WSNX53E07?+c;62cLWc1#WYLYW00^4d5Q&-FC1)=FVRPU3P;3I
0g:VU&^Tg;__;d7RIQ1@)bLL[NU_2dA96@AT7.K-50=+&<1&d>A);P\IH#<PXVD4
2V39RE0C^Q.NR]f58H&bN(B=A1]^LDA>LWZ>[R^]bA#,1UB;D_BaYOC[)?:/-NWM
M0B6^3)57U.#/N:e>JNOTQ6BRD(0Z_]5e\LPL+E#^U,K\>KIS&8.KUJVXCUXQ.Y-
V+>\]4LC=)&5Ug?NG1-eF<_5M@4:PA)6C6fHO#T)WY#<BS=+27)QfSRBV]OW,+K8
9=HX[S0D>^9ZeTgg]E@2V_E4R(6??V1F^:9:3TCQD)A;OTIGbMf2ZSLF5L:AHJ[.
<4F9N&4\9USX>(#@LI66TH&6^.P3IHeQLHXTLZ2DXbY1AV[P./C:(Ob?TNT+(c8J
;P0(dU4>8^&R3T3]?/TBU[ga_,N>Q(\.XN0^D5/D&LYT/dGecN=#=NeU<gg#]c<Z
0(BX^\M#/:@b?a5Z4Afec,Lb]#d4OZ:9_SY/<Z;F&MU9>KP6G]4OAQC?CI[fbbM=
6<(.ET@Z/96Z17ZCE+A67?H>O9Q&bV9U-EB2RJ:=-\+2D,=6f3;]EcE=5#^6N[E4
/6:&==B-ZM)[;IFKYZBeCVT\WJQfcY]a:EO128=d5(D+N;_5.IXK7COWeDZKb/KG
#OgVQD4XYf\69@,]6F)9L>N++@.g3)Q+7M)Q6QXT44gL4]5Y2-)2D:#5J_^V+,8I
1c0Y,N>#b;e@##RT0JJLCbD:,=ITV.O_QB8+A.1N:d.b]+6HM8P_@8J^:eQ>R]HQ
/;:15A;.^IXF:@^CIRV.@36Nf:,H=[Q/O/+RD71Ie#AAa^II6C;ZB>7[_.F/e9>d
KK2HC5G[/9Obe@F,]NVJ@9M^2ce5EYM8MeAMfJTHgfdYC5;e\U5gc6UZE-9Nd,UF
]W7>8dfCP:EP>SH#<-D.-0L[P1b8](OTVCUc(U:VFD[/L9OXCY6F_DA?\K8#XP8C
RH.?^^?SE#H:+BYA1c/=[#B[@4O-:?VLb4>aEKR9Z4e_eBH@CCgfY;#0T@@.<E;G
^#^fM6QZ&--RDd2.b=dc)/g(8f=OA^,@7MgM75N7,H]g;B5NA_Z,3O88=B8G6T-;
f&DFL[[K0bUf;c).3++GTB<7:Z1;9TYS((HFZC(=MES>^_GcXC9(W.0/.MP^JSb#
;],Yb=3WTF51GGTQ8^@0#(=-,.b?C3-F#2)b(=JEcKJ@D)#eR048a2fe,6(6#[bT
O/K(J15ND5H.;TeX2^)VR#X=2P,H]EPU:$
`endprotected


`endif

