
`ifndef GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_AMBA_SYSTEM_CONFIGURATION_SV

typedef class svt_amba_system_configuration;  

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PDoESi3CY3lbk2CAwwTIPqjv5iBzmnyi8dk6BUz4vIqVT4gsvAzpb0/7li6xj0Pg
hi0K0jZtsL+OErGBytT85cz+dofZWEUxXkmSikzx1ZO1Zw9cELzSIKxTTacMw0BX
c6wz2t1DClwsl5h6fwCUwHw4hVGxrLow1A1RY6BaPKc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 2132      )
g9wmuAbkXhhb7U5tH8nfrAgjheSzMNpJrbzuPvOVwg2uwV/d7o9LfO/7MXWvpJ0D
/+/P9uphFxr8ZSQWVpgWGvUmnN6jCxjjuejsMNodl5/37+SS3lzDlVLaI8oCslUf
GVPj3NRh78I/MB+1Z2hk/s3pCYItvt0ho/6LpRZ/950vpQCtEAwOaiWiYKE4ljlU
4H4Q8h3nMnWuwnOTJdN6GHsFaAHGxnrTDWild/yx8g8jcv5E8a04AqJS/BhODgzJ
KZR5lmlySMX0+nSRQJZ6vBLj9t9pt23ILsEg/ae6e2rxOI1y+XhNCg1J2T83jmxc
4+KOinRuBTmfQL/vifEdDU8IiM53BwuvzCDncI68C3nnpoE10QPTB2JWI6nokHMG
0g/cRVfIqxsy78qbY7wlSZK+UaLOd8vwgSD9/CxwnTEWjGvdTlhFTjhLS/kWSJMB
MDTs7nqeifUunApVC8bn1zJP4sLwfQ8dMWFcgU7DguuUl9X7nWdJreWJ7Mk3w+P3
xc325KTjujG1fvNfQqOfgXoCWzDsHXo9Q7RBdl9W/jT8O6GZvMk9SPDh7dV0UeCd
yLFT2uz+MKoWQvlc6baOIwKTqsLTGYO+CoLBuKRE97HJSO6RJ+fbbMFE94rbw3Yi
H87bfYliZmRqR0DEfSejvv2jffAXolnJ+OGi3min5dxi8BJ2k941BTVQYcQRsXsD
6gbbSuzqFUtuXGTIVoIc10VAqiH9fqnOr4Bl3y0tc8NJUGQRnFp959YgfZA5fdZo
w0LfZddlz2PcGEjcIzZoffMeEzRz3kxadFKOUU7g9rrvxgKQxQ+RANEpW+ACASU0
c6wDHV96Co0wDLdmQBjgD0i3Y1WlgS35G4j19Al4EzQL0294wIFQW+tn3X87gimB
/5+PckgwP7lkCRloLf+Tp2lHt0T/w/7f4KCN2YKlau1EzXaYlKAncuXHWQBYRHzg
m57+ntgefJHR9A6gxwhe6Mu6xPvCM2EhAJMbJt5FotH8m0jN4TvwafEp2OW37JmN
4hHU/UzlIuCXxyYDUCHgPD45G9BCVI5M6zABT/xgX22HnT7vs9NfrmQqVexIuAHw
xPaZGD7J5uml31prROocv+BoziOieqeYc34EG7SW5DgaoZfc1KrZt6gvASKPMEvM
OCHF7mwx4GaldmX/EY5T0nbqNTZFm7qMs4Vh1gQkEP9+ukeWGM22kla2Wt2qyHSF
9JRbRbEFkbRmYx5adXgA2ESpVNMQmWEl9O9LxjRiQ7oGhS5OGT3J86IVTfWHeVDR
SDjic99Wnegsnq3jDmXGZCHC8E93R3USy9nYoUlmphv4rHRNyAUreJXhRLRt3RJ5
mPEeECYVK2+/3hwSltfvRZZk42uX6wUxVjP1YecLn8Pqfe1wieAHTqEjNJkvdoum
KWdc1lVx2B/LgBua/wMwElWuvm1rEQDmHvFg7JWGfi5nPapU53ZF2rJ+fyqNYY1Y
8hfnTX6cpOipTSKndDqP/wM2Gt7r3lSm76WG7EZc6stXqtfgT4dHeQkqXIsTBIEZ
n95qkn06RV7pBKC3A/QYVOsPM8KQ/LLHfvUmaWYaRFnF6WXgHE8TIWDzzi/hhCJB
4vJHsbpsfMRWsGcnsU0iwhbIMYfaliL1lvh5GIalGrg16cuUC60SZyl8ivl5EMbD
h5pKmnFIZ4qOmGCzwKak2miU0HKOcZ6Fj78ONCPCq6+lmxtKApuHZMrOUZipzlij
153FRawRcf24kluMWWWnPjjxUC4b9Bd40BfMrvdaUzVySwEoXmtU5BIkpJkspEK9
muxOOywGS4Y7Hz57eFCAkbaJci4RYSx4BWRt9Ux9hsjW9DtBjDHp0nz7zrZ6ipPR
/OfSkNBDeiYglP80FIn0vu8ThR2dQl5wQZhCfdbi7PMPa21edZNrSLehQVAuYGth
GdV107fMkTE17Rl0S2iDRN0rJbW9WI56YuLxLF6Y8Ebq/OE+opdO+tuDuCiMqVqT
m4TZoWucdaNGSOqX11YdLV2m7WrFdN1XODGhEd+MTW0Wd4Wr8SEJoVUkNA1dnNlY
lWDSW2rWsoaAywNdFRN7ZB/SDYUd2WSLRvSiuS8jCtdfo+SFmXGdgWuS3k6s/8bL
fI4iDDTpB1jtfH9jWJTGzuuEB7sZu3I+15wxnRFbRcBfZsHMAWhtYlM5ytzkEDdn
erQYGdLHIXsfa7Cyvu/1FrMorXpIm/SaY4V3K1KQTbybTWkmbj+s5NNXT1kvJULh
Py+Qbcc0LppZJEVaXoqzanp3dhtia9rg2xQaqrHOQOuIerv1twF+5zZf9ZlaHLvp
L6tqrCBql8qZorNAMUc8lc4ndGZbmVI0jhih8FV3fANItMPvRqtMF0xfixz2DK2d
aniDr1ayNonBz/LQgGPW504NgDEbYgan3YVo0k0noTVR/OqWYvROBRNFIIzTmxXz
v/SfTHB9DxPZc8GVpu+MRhT4+XZTQKTHaK/FcIFEcGYNAkiiJtnkcRKwEwC5F+Uk
CNrzt0GvRLL6il6tjM2RiqubU7u/aCRPFMhDg9Spgp57j9Qocc+zNi6d4Zat5uUN
+5IXGdtsjUeCN4L1qwZ4TSK0zEgynpeY5EGnVkaRhJCRhGSMnO6y6hAka42oHjIf
6mNeZ2uc+Hj/zqeJ2+KI1oYYIbMt6kV2gy3hyURbS7LTQJwtAX1N51FFDP5OD10C
COX6q4HyNRGGjbo24b0XXgOfhhfet4MHRYpyR7QNLapI0JjGv3pF/YwSNE7BOdDh
YbGOdYVmu5D6NxPcbmesxgyMupWF3bd2oXCZMasae/1jPntg5OPI1VWJGhvWHWR4
TKhhHE8s0TIS3qJovgf3XbrQFEnfm5gz3SzpnNXA/RA=
`pragma protect end_protected

`include "svt_amba_defines.svi"

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
MIZaTPhOq8eq6SHlg8uD+Ld8ed5vFove2vvEgyQU0ueteylV0aEbe/NQKPRydT26
SsP6WZd5Kz6aNH+TlQwZo/JEFfw+1U2P1NkwStSH9Q5xiFURYgOVjbpm+JQ8kNpy
UaXewGUPVl1qJxuZhFNCsRTI4b1YLTmN3C9CZAXb5wQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3141      )
M5ZsKdnXmHdDQ6gTlUCzbCugUh4vXfIaGvM4VZ24Oqq+M+q13hpYpCpgQnhAa94e
9u+msywvdGvvH8GuwasYknV0pBGPGFmShnqg1XERFtWNgTT7HTcNFoaQ98xQ4sEV
6HGp9RWRmkTkkQpC/CSMl4fYe7IQkiFSuBBWltA1jKye0l6XEsw3Rn3PoPVEDlZd
kjnOveFT0D/893yTdTDyT+Gzkm6uizmf2FhzAgdMutvZLUu36C6xJmc3w4Z3VG5q
hVe9R97ZZk8JQVC9aS9Ee4DbfWuyqtPQB0Hy3R0KiINfWZhUzjPiR9Iu5yP6+/ct
f77IYrgBbAJAg1Q+wckV3tHgPQpJG3hzmtU+xh/GXYeTcSgHI96MxeE5uq3AN7AW
dZDk0SpESKGPWOWjeKfDzcIv9BvfTGhP3I8ka8ccmQY0WPAk63Th0st/wNXU5SuE
DPliDvdxo/B2oQks1x6s09naYZlaYUcVcYfXhSce//SH6JDZJCyQq5gFHMweDOfg
fM2UDS3imn/BxQjJIpIkU+lHPsrmmlVauNv74JsiYE93ov3arKqTgP0YwliCz5rC
Jfzy71we1fJu3NgrIPvWdBHs52c7QybukxoYDh7x5dPgYUIsTD2aLkGpRfj2v7qj
5N87i0k0nVaxcsWaU5e+VXqg96f5Q9scgW50amwxXPToHGm0HIDBhg/eWzL5G58y
HFAmuu6RfsNarMnfLZdpsZ0MnQFFVDzrzh+lYq72qnZiAYs0TL6+Pu41TkL/OEma
9UV5InFEp2FWz4Jof0/1DenbT7YxU5YG9/GOZizGnTIaF1QkwTtwyxydyO9c4O+A
UFaI9Ef6Xc6bgfr+ogYk9xjyOBAh1qZ6embwwyJc4mBCMRWHz7hFjH0A6YLE86o+
ForVq4kzoYizZN8toh2eRnRLjfW9rGEFYDgW1I/xt5ydEV4XGmh+k8c8XRXFSXQn
5+KrJ7nXp/W4+rVW5qX6Z06t+RX4W6qtYpqPn+oCcKxF8NYrpMkQMc1l8whUJgmY
9TStOvtWAFY4hhWrY9/EpBIagd7C6pKTjMFOePzqz+4rAUtifqS4hPqlkZNz6r4N
rFiW4rHUxXd13r+KrHxDpVhYBIZG3eSmEt+FjzP5KR+/7ZXYNdjKUdYmPCT5dWtZ
RqZROkoTKDaZ3b/ICBbnRKZvNA0RFSy2G5WSweiMaUKdlct/H9A60P7Wc14gxDoA
Sv3YyOMMMyNbqXEXqdg4CPQzxAZ8BZWUtrakQHNNxLm/3I9i5dHZtSHpf2/6PVSi
R+tr/0ORBwevy286IzkMIFJ6cw7CI54rlpLaXbeyAYcwtDTM0x5y5b28jf0y3ior
YN5Fb/5Cr4PuLgP+vWf70w==
`pragma protect end_protected

  
class svt_amba_system_monitor_configuration extends svt_configuration;

  /** 
    * If set to 1, the system monitor issues an error under the following 
    * conditions:
    * 
    * -# If the AXI/AHB/APB port to which the transaction is to be routed
    * to based on the address map is not specified in the downstream ports
    * connected to the system monitor.
    *
    * -# If for any transaction received on the upstream port the transaction
    *  address does not lie in the specified address range configured for the
    *  AXI/AHB/APB slaves which are configured as downstream ports connected
    *  to the system monitor.
    * . 
    * Default value is set to 0.
    */
  bit flag_err_if_addr_not_in_range_specified_for_downstream_ports = 1'b0;

/** @cond PRIVATE */
  /**
    * Applicable only if the system does not have any master where
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    * Enables the AMBA system monitor to handle posted write
    * transactions. A posted write transaction is one where the interconnect
    * responds to a write transaction without waiting for a response from the
    * slave to which the transaction is finally destined. When this parameter is enabled,
    * the system monitor disables data_integrity_check. This is required
    * because a transaction may not have reached its final destination (slave)
    * when it completes at the master that initiated it. To enable data
    * integrity checking for such transactions, the VIP correlates transactions
    * received at the slaves to transactions initiated by masters based on
    * address and data.  If the VIP is unable to correlate a received slave
    * transaction to a master transaction, VIP will fire
    * master_slave_xact_data_integrity_check. Note that it is legal (though not
    * mandatory) to enable this parameter even if a system does not support
    * posted writes because setting this simply enables the system monitor to
    * correlate downstream transactions to upstream transactions which may be a
    * requirement even in a system with no posted writes. If a system supports
    * posted writes, it is mandatory to set this parameter to 1. Reporting of
    * orphaned transactions is not currently supported. Orphaned transactions
    * are those at the end of the simulation which could not be correlated to
    * any slave transaction, which indicates that some transactions did not
    * make it to final slave destination. 
    */ 
  bit posted_write_xacts_enable = 0;

/** @endcond */

  /** 
    * A back reference to the svt_amba_system_configuration object in which
    * this class is instantiated.
    */
  svt_amba_system_configuration amba_sys_cfg;

  /** 
    * The upstream (source) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB master/slave configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int upstream_system_port_id[];

  /** 
    * The upstream (source) port configurations of the ports connnected to this
    * system monitor. These can be CHI/AXI/AHB RN/master/slave configurations
    */
  rand svt_configuration upstream_port_cfg[];

  /** 
    * The downstream(destination) system port ids of the ports connnected to this
    * system monitor. These can be AXI/AHB/APB port configurations
    * The system port id corresponds to the value of amba_system_port_id
    * configured in the respective port configurations. This is currently
    * used only when AMBA system monitor configuration is loaded through
    * a file 
    */
  int downstream_system_port_id[];

  /** 
    * The downstream (destination) port configurations of the ports connnected to this
    * system monitor. These are CHI/AXI/AHB SN/slave configurations
    */
  rand svt_configuration downstream_port_cfg[];

  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_monitor_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_monitor_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_monitor_configuration)
    `svt_field_object(                      amba_sys_cfg                             ,`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
    `svt_field_array_object(upstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(upstream_system_port_id, `SVT_NOCOPY)
    `svt_field_array_object(downstream_port_cfg, `SVT_NOCOPY|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_array_int(downstream_system_port_id, `SVT_NOCOPY)
    `svt_field_int(flag_err_if_addr_not_in_range_specified_for_downstream_ports ,   `SVT_DEC | `SVT_ALL_ON)
    `svt_field_int(posted_write_xacts_enable,   `SVT_DEC | `SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_monitor_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_monitor_configuration)
  `vmm_class_factory(svt_amba_system_monitor_configuration)
`endif   
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
XnuwrCZ5u25qZY4FK4CzXjGOuJoy6brQq1dFMdwt1dolMvFG06t8s5hNBaEqeC1R
9dFFyvj9S/D1QuHkNMRwxXi1BJMM/3G0IdaANkczw2X0fKl7GdPIQ4LMynd+MirI
H16ZGdzo077ff+hGsokkeEd2bPYbFKLtAkA60vUYxEU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3787      )
qxvXhQhhxVH7494pGb16zBzYCxsJdILECpJe2EPxexBggjKvrkOJbvuYhxwX1/PH
CnqCER3TJNcNgpnkIv3WAeAu6JZu4k6OCxOEjdf8Db5KoJiG6S30INRveCgfsgNo
/9iuA6gSNRK0h0AHN4KIc89HkgaiDLK1vaucugax2qYgnm2mOd8dkYRFD34TkomT
S0RlDWBm09XrsJEr4Ld/HITD8aTYcS7uPDjqdgNhiJrUUcwY5DFqut1cWmWMlDVZ
aHLH/RgrU1PahTDZULSNcoWZ4JWI08lboDhdEIIGJwIPapj21h5WgHsNLHgMkWaw
yzqN8cX3w1BEfiTTXD9YVNa+Kl6ablfPRxafZaW64AETu876BWGMfezKCIv/X04x
93x6X4bldt4jk20fdWoa6IJuxA061DzkevGZsoIzn4cxE9uIDSQlO/7jfqV5FGFu
vcdcIfDtvakssDqkYYjYZ/Sth0M2wPcra/faLrd5i76goqAMiwx/8UINiEGoQoLk
HUtusvlhzIVmBcZFPvV21qJTGyhmQyp41f4tMbq63k4OzxWhhoN5QIgIP+wtuP1y
+aO9yRtiYV+sMp8I12b46gr7ttGEzkks4beNQbzjPQieHZNjtwyjJG7C9tXwg/O3
krzXvvC3sde/LrHyRIeFNDt2OrT7yd0bfwZO9ncKWRkakaqVMitXZ+4qNYjccGF5
La0wiLS/8jy7HLChAfvAjs/lwYHXuGmQv4RZ50XCKlWqFSwceDCcRvKIqUNE6bKk
3gEk3w8X0+lbMsgAqCoB7YCUG1mA9NCvqQObZZz+++YCx3zr5pOSOEpJVsdrnMSf
qEmuM8R8IZNGRAmc4jIbd7P+PNgPzcglFCKgHn9b//g=
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
O+aGvt2+i3ys5V3+oGF9TVEMpBf4yG1D4K13Yp0mbhxoIXDyet0YJBcb7lSv3Tzo
JPhtk8xd/BWhlS/IlSSrPDOiLMa9QVNWMKBecYrHJRatIdzFtBzzeJNf3ZNa7Dgs
RbUEySGyV/0C2ERwCNl4boAR/FZOnzrpz1pb++ee0Hs=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 26340     )
0eeOAg2u55iz4jZZO9Reg3wT+kZw58x1Y4ywqPVxb/pjlfFEnEX8NQsnycEtnGgo
TJ3PlO9Pywj93NV35SEIzjJ3xIFH225ttxJYCh5b8RuS4Y4YN/o0J7w+k33nWvMC
ILRjUKyJ/fUmtGrjJHiH6r53uX/GTSdfS0l6H/30DFHs4FVzzf+K2+bnvbDXrWxY
9V8iO0Ap7ZldJScSzGQt/iFIFfszvBA12+AOYAdqSw5TPJy9/RWTSnmgrSAohHbJ
PZXRb40W7ksLCzJo/rrJKkdy3yL/wlJ2ejLDWxhYqCKH2EoOCgZyy4o4eJHrbGhW
020yxPEGYAmCyt7v9PRBaT11ywhL+QgwBdMbRDodOUl5vrMSYlyENDE+w0FzPejE
PTwiY6blor4sveshIbaFAi27BGaQkRCaOm9xKVscDZEscbDwLbkJRFmHuztJgWbJ
1iQIrxl+Zs6rOXJowz4bWDZgJ4XxHL5wgA69ewgm81XFvIQ/yd3jXG2RRawNhu3U
G1NRmhxW5MuCSIuoKD5orR0gUT961E7PpqrQNF51jAEEERhuoXdR4Aik7yLhcOwb
i3v9hAOpYzzAYk7j7y4n2oaXIzsHN1NJuQRsj3Q5/m+CjV/eWgd4X/YWThkCJ6RK
2fKfx34Ko6iSFoEeQWuq7gGlPQkwHR9lesPGYHjrnmKSGK2k334QClohRFm66FYM
ojtxz45VyNUnsjV3cNcNJhCThPW6lSw/RgOt2jpnrzzD6VPE4JCiv7aq1Bo4It1V
SLS8/jhee0gVwJHJBlYff/QntiszcLHnmH13qMJt4LyjMhb0rETKYtYYHr9w1KsA
qeix5so8Dyju/o72j1WLO+4GVjotBG6Uo5pFPOw0wCfZB03f1QuxSmRV5xILnLl6
t+Rv1IthkxRa7Yc9YXrOb2TBT7UBpdn9pA0NjuDcyTh63ofutL1aPNZpLowGeuC5
UJJsUwPLCvvTKeV78hoyJI9AwkViwypYb62qEtNyJ/Tugn1ekNLxuyZc9ZGAaDRp
upxho7VOItqNretMWoIvTcSULu5hVzs5pYgrR0NyWVMne1JOMLF+a2hD1JqtRCyt
n+qGxCeBGY1Jhjcl0fmVx3BU4vplcBm2xSTrkIOCvQ+5Qr8sjx2yT2SncAtZ0cqP
vltOKTJhOwCjmomB8R6wA054eLuyXtWxdz4NgoOU8IKT3RojE2/zI6DiHYpkgeKK
Tjn3vOIr6h/rRd0aO2h02M8PV1YVIi4UUVDY8vwK6gUKUIgCsaRVo7dMRmCW1yVi
L+PUcA4WLMxcfzcQHpEl7ZfDU9x4esGHK3eyCfxgcOH5CQMBGtteO+P5Lca1n2Dw
TaMN1DKp2s/yIKJB+fjhryVa0dMxI81C/c+1J51ZD9d5UnswbPzoZNR8ZVE273bi
pIa36YTKXUqZyZ7v1NlXlLRi1uo6Jz/+3eYjkvhbfFCuNbanETxEZy6bAowrmWNQ
PXlK8mYq6ll+uYHFlexOY6/irlEfnUUyabGsDBKsD6+w3d6Rgc9zi3ohp0U9GMbv
cKaUv9re4jr6Eqx2uC0KdfWqbGy4gJbbZzXuyjNOuuHiIrIqrkEUINbKta4fOR0q
aOGKCIPueyrAQbbnE9snGA8fhN5j5fyiVpKGUeK4Ch8jPodeIYrhJ8D4vcwbRTyV
iSYsZPNciHHYhIV27GKoB4ICr3zOelDT8qsH1/7/jDEU2Gh6XzjylJPoo/9Eq6eH
iVryGwviRkCIvvsHG3k7B6Zokv85Y2GWNmeEaaFWquUsI6FKvXcqGAu9VV7AXewL
H9yulEgkXLTdER0631frr0kJ1h8z75cI7YLr4blSTQtzFgriRJuXtGPZycaq91ga
0k/Z4Tr1vIMN/hqxeXfI3tRiN+M18QPdGhsAxY91/mkGAPZb68RLMFOuUU6KcKy/
+5s54TosqXb8SeMixqiNfFiq5NlrddczXEkzNsvYFNLezd9/NHPrf7j5p/oNYkV0
cYsilLVMTWVyS80U8hFzW2rUy10i5aM1eq5adelCd6+LtLUMe4FNG3zDPuM24Vvs
2B8S6RTeZUdCYfRSpGwFhBQCfWi4tndfCUTK8IxZykPqvy7eQ69g+R2ItzxwI24M
g80YBRQsSdH81v4uJ7wuq6nPm0A0LK3aWoqqxBDI+7ydjVyJV8J9LELvV7W/imqz
b+S/lW+y0WVg7Jh/7JnJptklryW9zhAhRSDI7zOjhJpsEl++3aGNux1dfrqnyTUY
GieHUhiXcssule/b9fiFm8HT684/Xo3cjJE9/cBYm2fcBGkl/qge7o1+ExWyt/Zq
6yO03H09NE75MJbXuYZJ9JZUAY499tHtipEfDMIkL/RLbmO9xyg4myPUe0QEnQZd
1wPHbWv9SpNo2nrQdMyqfZkMbYPewryIv99XVbx+FL5fMfe+4vuHHYrpJLdX3+OR
JMKyCa3suq1AIZkdcAxT2BZtbB2OVqw/tc+obWqaDJIKnnMkFhYuRjC7UTCjVowp
Femce8Yh4bf6nYVkwJGQHAdGOdc52hnxsvZnH2wded3M2PqUS1OUdoH5BBrEZ7qi
Ks4IkYOx00PrkrhpDy1JmQOpzdVwXkEMcGajiADUwf1l2YI9BBwdbX1N2D4EfdOP
ToI+r9+DWYJ+Ptq5PP2kqnYHnr+RVbsDqxBFbrBzbbdt1MlMA5K736gSM7uJfcqV
ZEJPZ5k+H83HgZDgimuXDk3cX+jRfFm20pW5IGT6vnKJd9llAJqD7FWGINbwTPVm
g6O7I64h76qMhOvSqBFdOn3GrSKzyi7F9clkCX7DYHvZIuJ2D5rv9yimx8ZmEdPo
e7RwjIaavD/tzBnmLimomr/sKRAaUBQbbJTwqOUmUnkg/dExl7xyyrRdLY3uh5ng
s02dYlMGmIOov7Xqm5SbLE5i9Lc1u5mPPyiqBMT+XD3FQsggWzqlNirt8A1XMODo
MUktaVxWCbxgjwORndjTnXgilfD5+uDRMu1vWpOSszc3j3JMcFsw9ucWZ8KQMpLC
lw5BjYWPNHZr93hVQAvxuoYR5uBMyHVTXBLH5XnE0uyzpzxq1atwVduLltWuzJ2L
CGQgSmfBRqE8zxQ/7+bV3dxhAsZjNALoeR+YYp0SYIJE2EgSWnpH1Q11DIr3KXmR
E8Qpp2bcYP2CM4k6UWlvauTbe8aZbunvKIyK++83Q6WWjvXLDSuUKEWzAqAvD6Py
lk/3mLIzenu0OgciKloQVm6uRD+tBwJd3zFfKVXcxAZ5+Gkd86uarj87IOSYT9rs
lNZR8D21JjR/tDO2eluKgblLEj+NU8nwV/15T0rmqRjErB8Mw2V89uX3AOlybIIu
sQfX+NAEHuarwc4Py/H0WJUclj9nizBuQa6itulNCU/tOd/RqcrjUHKjWCnJwuXc
NOX2H4fOYMF2hopxxAaAaWTtOpoM2aX7sIspq469SP99XVD16lBr0OoJL/SqtZaT
trmndBmhMJDTiMwsvt//6GslBXk0iiISJC1wL2uxe3OY/jxPl1us8NA25rWoE2dw
w0fgPcyyrmSEpxP4XYo0yEGrYy65TyPSdOt482J6PLucW2ZsvVto9RoLueJ8Vc7a
XylZ4Bu4pAsfUmOIXqH8K4Eueo3zaDsDM+WJ4r4Xqw7/SZvGm/tNTxECvpgwyQMJ
tMltLNdUtWzxzrWLZGGSPhe1boTQj7fDjev9T3Mz2uop0y84oBMalGDy+37biRRj
fVXrOm8JZiFxeIlH3P7kACz0CqJegEYmbZfVQtHZ/ZqmrY7wTHwhfuWjeyXLKBYo
atU8xPACV++L2T12bCVIbAtTCSbUxwBc4TJqrbP+rrlpw+NFudwAnlqtwir8yltu
cFH+9qAGYMvK+LzQu3Qpi8z4WH/bB/45Mc0noCstTKbfHmP4X83ZsvKmW7OC6M4f
+Tr13yBFypL7FjPQTF6uHrrwBrxzE/l5wNrnakyw+dUTOgE8cjD2tFO6flfY7jvP
zHEcYNCHjVDg5dmafcCgJuiDKBl0mNoMlZncXMtr51EjfLAsIwrMg591bDn8/f/S
NeS+dPr4f2xJKUUR5nVgrWniVkhXvC6owcggOKY8ydP1p+I7Qy0dzqBqnc7H+jap
4E1SUJndFf9xt6waXM/eKEwgAmRnZF8Zr1F1YmbO51538PCoxtB9kDB8r23mG+FC
/L6EEnkf+sIKG+SjiIEF4ff3ipOUJd8/qwaksxBUnEYyr9tSQXzo1BidWa/zDiei
wRj4U2JFc4FIGQlKYvf6a+JabdNdMvH7w0KaaP2tNEd46HVToxZMztYl0SJW9CtR
r0gDtzOWZ9VQbn7OOxEc7fnuXstwAqV/ecz76cI7D0CdGfYvb9/5VLx6LoL5rroa
5xRKmfcHYFvqOLTlmeSiC7KoMAe04TTkw661yo9+oa69B43F+87Va12NzTAQg3iE
TZIYotusHT2vRKvxeTut7TO7hSWuUgwl0eRECLwuC8s6cA9/xkD0qJ4xoLIKY5Y+
rAuYzQlp0QT7YVOHqOuG6XGEb6KM8XdyJy+3fY0/uNQTj5a55VUBkHzqKb9R2r+A
jezqzIRkKjtfjMgV91A6BS7TYfjX1M+Krs157uJGPrnKWD6bg/Dovboh+RvKClmk
PridFZG3oyST9/mGpUK3gyDOzWXI79kiUy2fOvDC0sTvs29hLfOO5y+I2SViFw1p
uBSxpJnK9n9Lfh1PzSCQVTo9FKb5P8djkk8O0e3RId+pmdU5m7YlJHjZLGd/Rpu1
6r7SpB2D408PeAL6Ac++h+WNega/AASd7Gf5/8JxjNwgLyXhIrJeYc8PAJ6WEKNI
fEMWWEYo2tsRDDD33UF7fPwWcP0LBoTM+Cc1GhFfWXDw65NK3UAOxRYI/TqYdA8j
tvEdoacWg+vyNEMkgk0wL95BCzaRM5BCAJ02IcVZ9bUdyh1SA+icil76RPW4nzP1
sqrhy1pO9K+pQhlSlDw+lB8+H8Xz9umoF6zono5JohFw+AUKz7AkzAegO7qFXIjA
Kdxbbq2hYPkBEn0WkQB9shUjZ+rSTLYqNpC035a23O62MabEA7uSBMa/Vxr5JL7x
XukJok5ZNKcd60Z5xWqEAlFVRQSbBWe4V9nujkYhjVcmUeFTNQPSQhSr9v3dLdMI
VIbfpDpYFiGHhVPs25LygoimhGxXrR928Ns0Cnox2Py7Pvs3B9OegnPOZQmEDWTI
t9f/qDigmnLNiptpiAKeLPXdqkfWgccmqK7vARG479cmInsWAH1DboCpJpkUSeaG
uiWsTsUo+uAHSFDGxgGgSM6vb4qP46f9uzmZbMA7yAfueEj+7MLGjfjF+x8JxKCx
NvJfWoURh77WMR+98LBocFgU0OcCW8CKoNiETU2MDZFBsu6RPyo8fpeSn1BAVtw0
EIaapMfnwubsFIXGY5qm2bJwZMmN3bdjZvjA/V6lSa4YhVdhY9Vc5mYvjeFg5K8y
dxzFFp0dIlMdDfrgkq0SMPlFbbbyeDYlwLa3yxL6JPEQcKUTlh4VkmMTTaYH15eN
mpCknDZ42tubviBdwpLzfimTFHMhRRrQBvdpgunmB5+sp3HvhcSx2TU4c4Zu87UO
R55pljGyjBT039KxABTpwMzXJgywmYjnn8HV6DesHLVT8yYEQYtmWjyjiIdRId41
vtSwSka/3v6Fgu++r8FYdECsm40L8qxGWMkUQADctwEQ+DGgrz6lmhkWbrUtXgZg
NZL2MXrWc2EGkkOEA1WodFsCQy6wy1sdsEaVXFZTC/HE1OEPA/TCGBGny9WsdlAd
7iQOO8VzyMALOBwOpT+KXuvEELFF8T1Ev9o0Tubu5by9BDPRluANk9Aqwr4XItsc
WDpIk3ZcVIh0rlALdrqzNGdhjM7T3oiyMjQOu6o0XRfeOzGcYeMfMsr91cDi6fQM
m9p1xxWm9SFZ1uyk2V2hG8XM1wRSQcM6+oKqFp9DbIxB04iJSwihsLlovGENsOET
jQqGQwHnT9rG+hg/FJTWwIBuFgPpZlUNrLGvihbae5BCmvMv2oLwKvz5GD3pR/cr
sGPYi5NyjTiE/PepENXqLEAELTo2nnatvI6N4TVG0to/4BfuKl0tZxKd3jEWHOcu
fN4cGQ9/QP3tn9YVVsAfCJzN800dTOh/kiP2DpYmfrSyBugUHoXCmf7dRJQ/CCGR
Obin7h/LRLaKMFPZe9YxZ8IXc8QrMjsvYCf2tIqcQcCbN5/hr7AsUlXtek3UxHG2
mqxZAmM5aRY5G79JlCeKXxcq/IoFadQqaTOiQtKtOPFr51ABgAczqTgRhEjPkOu5
fT1u4RahSEj+4XV5es274cmP8l/vSyB8rAuJexGnVvtIPMjsOvDnkFZ6wriwbc5Z
Qbaay605XPYZzVPcX4i3lzZDzYiOsAu8MnlsvRuc/zTzXO2My9EXU2D20yRSyyrO
oCAg4pCqwKK5+DGxVS9tNbi8JpDcj2evToN4t/QxwLRDmh1eoDpkuEh3kRhVfwT5
gd5Y5rpP607wxB+431bO+vyS7wqAdyg3NgrDK10auapJVfPobm66kKZMc8FSWeYg
4R/nSTIm9SstKVzFJB4ZkUu/Me4Ii3MC3LT1ptVznvBNhwAElmpy7RhkUlEknL//
JxdbWLmSJdXv5FS7I97wtGF4O7TSFzZjVsnzCmt7JsDK0aPyIil3Iz6fADT+Q7tg
Wz4lZ8oHGs7B3LM8ACj7fxlOPT0rZ5Mlb0YrEHdKgPSRdMjBy7dLy9BDlwfqUIi2
pKGCst43iiGrWMHMEfCyUhJHXpVjDi+9X3TIWFXWEH1WnarwcckfzIQmKnrZ2Rzs
sICb10UGp4i6I9+gN9XTdQjzyg0GiPtHen2oDNHxnjVrRmpXCuQ3N1zq9/g5aq+c
/XD0nUIYlIa/cSiwhMf0WXIMLLMaQawX0Zg+QUfco/YG6voCGgO2CIOYuYW2aXfW
YMlYd5+krcwqu0tt+6OBhhb6q6vERA3cDqiTyBgfEdvmvj7KFH7BALbdrwplrWGG
a52gB1Lz4ntmGqVPWMqfHJa2+EBb7yRkhZoHumNWhtw3qspJmXJ3Mc3xfVp4cZcL
pepGat3v42qOp0FZxesDye7K7in51CgqZPx7e4aHdHAQokvAoz2EjGc8QACKv2cw
3OTac38s1cZ5dsvgibR6Nd2BXP6T+rHAL3sPnsv1Viu2HBsruyukTIK39ohZeoRD
RSnhu8usHRNJzPqFPRWzTV55an9+qtM39iszvixqRsBVbszHNOew7eKrenUyG0KE
oP/21csPPS4+MAhhgYXHlSSBaWBQSmA+JQDUdYXrup5Xb4460jJoVTXwscTrHwyO
Jwjbx3+QJMcm/5i77UFVa32mnvbvlQS7/ChZljNScfiY4AfocdppFrEpas0VfHbl
jCc4ycbPLHnQvX/REQjc1CQb+AWMa+YtZ1RfLNobo3xpsdIfxH41qXG4TyayVQAA
VJTWqtQQiDuI66OrlOUNpoP+Gdsuorrlvv4RQdLIosjx9VGk8aNrTlyZIajgZLel
6vJdypudK8ZNlBmRyHK6SZ3Be9ENqbVMiLa17/jd/16RVxNcJjciLb0pybvyVV6r
DWr6uYdz5V93JQVggqVIOBtsCQvINULVZbUbWflB7lwj6moCup8zqsVxnNSBvtin
1yCE4rQIp1jni/vo3zb3NFIlVRn7zHQ6xKQ9TPXTmF6ypABXXfmVXK0TDCZwvtT+
YkRxZoNiuRi7KXZI0Vc+TJcODCl5ea20Ee04dV2Pj7ABF02eBuP5z1gqrhPGmaP6
poglXbkKdnF49yWU9unf8WIDBNEaqheJStHbsYN8hI3pjxF8kUEbUT9KAKDcKLjs
5YpwcR1XyxZhw6rUOzWmSJxqCt3AV6OpkQdjTqwZ5vzaqC0dG9GOvErTJ4aUA2nn
Okmh0MoS0vh67ottrLvC6np/7E67dgi1ryOjqHld132HFyFTM8c0Hrqv11FT118L
t8pcTap28FKW8mP4h5WuHKwPtDXqaPCx23Y+TV+oCQ86QB7Fad809fJUSSN1N2fk
wMKLjBTATTOxokSV7nCh9o0J5eu6/hJYA6A4Guj+7KHRL0ZymfhzkrYVeRw2Oi98
fWNbIiX0rT4ol2l4kCS0abYBP1fImrRCrlImJsRru2fZuOdBaOwkTfzEZ2s4sHVR
ZS5jXS1K3FQvIp8iujS1GEFLpw/YBAMbvMVlD395ZjTv7w1ssr8gMaCSk0oq3D1z
lIK9bIri1Tm70vz/BJqCTBy+wJrbr307sWwqsRySyYrRfegshq1ZtQM3xvFubfds
M6jvQJW0pVMjIuvrXf4revWlVN+bV/6UxfoNpy963JZ7rUnnCj2QSHaZURlYG60T
PIKcX7w5Ixf17KekAQEsAH9ouoSlwYP+s7uvy+DhbkM7TrxDKSCw1i92x1vDfbg5
pBGv9rmSXdYWpSbmYcmxv0GblEKOcx75QUYisolvOJb/TmEZSbkdFyuFslGqBJL3
2stEVBzLyqAANcQvcsV3mi1/38k/UaoXkDXmz8bIWSznXOh5QYIE63blDcByESKa
si6wCgGyO06OMDFsDvrakuRulxSVdEKqKGhUgjM3WBee7Zgh3LdwmsNIzHncW7a4
v3rQtKcoNld5HCNq+6zaUwl/bR92QOk5De00CTCmhxvmZbRpACgjcHFZil04/z1j
I8N9gOVEV9S5j2+HizsPVQ4maKbRWYFWtL4k5A3VDjd2YqpA6wzynDIcreK+Z2dO
am8zDogUliojZyY4JSDlf3cIKOpF6oSrUssTdUPPwQxhw2Im4OcDKlsOHN3hTMwQ
L6Kx5irvemP3aPaBs3poXmccY1ahN1hOjt30ValQZpr/lE2buUqQBE3Q5jb9wEy3
4v6NI5m6GVMQZ0oODllcrcU0qM9WBfn1nME5TbXutAMfhpdkH2Ei3nCeGC1OU/Xr
FmuwJn8RS4apR3H9Jt5bvETGLIbeXucGMlpZAXyyKMp1dd+UHGFXciEfVA9PyZ4N
/wYsyU3NbeSnYAL0d+lA0zKUmvdkewXbl4HvpTgGN9HMMcNDJr02AP7QKrXVOt3R
SZgJofjjGrW2txIJb4UUWMDZ27OOg16qLoy3X0j8U5Tb2V9Pjt5RGG/8mhy7QgOQ
fRklRnnFdgj8IcSrI5aG+cZNdnuW6qrNWx8n7OmUTMFmUnufIcW//ONGjzQnN6SA
rvMUXlzuBU4e6kQDUQ03F+ikCV/cVdGcXNKQCMc+coEKg0ehQmoA8u2asHbIVMY+
Qqq/H4MGVBrcdYiE6u7WdIdWJm1qQEQMFDF3lVkmeaxp7evYGPX32NsRh6/pXf8a
yP6BXf5w52gyomfH4zsrbN42cbUhof12VDWQ7oRUP2fszjOTE5SBZ2VUeb5+MBVD
CZEsLPxyx5YMxrcidjOa6gKBEzMylFMhUYnF5eNJBXTY0JdcXDu5YV0a+8wEcZmr
0zjKFGb92eTzrNblwrWSwyQjmWPWHFpAHfXuM9J6xzBcig53XPLdrhQ8Nf68F/2s
xXPGKYYz/7lQbTnbdIhN3F2Mv/T6fv7+A4lmOcyZ9MlRFE/Uuz6yylJK09Zfwzay
cMTSU+PMPqs41KSkLDmnVWGTU95fUelt5g2394wsBbYiyLP7WNPSifZzP5fko+Bm
4kvPjsRPyuQW68lAa+lVcM5/8RLaJp+KT3NBjmEph1fQAxK6iolJ1Y+CQW4EzAU9
llF5ubpwo5CaKysTabyhQivM0gXCRYxXz8xvZhbgi4LhJdXI2Pavq7GJxsEx27XP
NPEIdITnHGpVXdPeuU/gVqN5LcA3WCVqfFEyrJYVvY5TDHPrhuzJQFk824BGv6/c
HjejUPSNE6PqJXalx0ODqa/mlg5fRE+kNfkUjbHZw3w3FW15M5axM+sAu+vMm3JU
AxcnyiE3kPPZkE2TM4OnwwYrvQSQ1FKYlwdvpW+rIFT2/xkl+mo82XjJgnhazsbL
/EvLMp3k6LzY20EyeRkw5qP4WkJvqReIH0PWjt8IMxPt35M5V13Ff1TLlIrpHADa
ABe4Sh+ruiy76Tc+2ouPsrtGVmk3kw33JkK6YLLvPMdgDXISHRYa22bWUyMYGPmI
2UkGSYR/IatWGIk+Wi/0x54tcAMRWYSG8xYTR8Z3+tXaSh4ydsZBZ+Tdtc0wGTHp
qH0kd8oyPlYToV9mK6H39B1YLqZtgNBaWyVt58AzotCesGiuARFFtUrVxStGgMB+
oEC270cdRqP5b6NNSaN/KTvkV6uztxTb+WVDEcXLAHJ2Zs26sK5GiuMFW+XvRC8N
Bg4tRGhQvEZOz1PANHNAUkNpEy4oFJ0RuroJKtbFRHcAa+exjvs0vC10vulzYGWR
QuiIh9DkPKLYLBvypP9XINFNFzFD+lbBfV5Isye0wqd/Vwd7k5mvtE/17kDHlq/Z
BhtSXLzlsQ23MvLF8s9slfkx9p9kEkqD9UWkiVqnHL5X6reWweEZLYeg4LA172jn
vlExxTjiDZmUCtm5fPqcYdDtXlplEtS1jVtSVVyPBzI+33h0vgG2x4Eq9lj2ow5Z
pCiJx0MOx9u2ZNfQCe2uUcZR56yc1JByrbfZYgBdRTdOEAR8bV72+h5Kq5xvhGU/
slAaZYMeFSrQgB7D2iSw6Z7tEezEcVExNiXxS8pQsHoKOhcowfoyN4S4eLBY7WKn
zKeAx71oMtkwejwKqMXB62vCEh7aRDMuLOp7IsVwX/HClKWC3KkPjLV9G+tZLo49
ILUl0MgZtpIG+P8Rzeatx1EL+vcLynVei2fVl5+P8v3w4pCyW1lX3+4sKxSBVMKk
rLGwXdOtY0yIPsQfwI98frtVMLRvGAjnpejKjkW8rqywyR531vQMqxK7OWCGdxv6
XvsC3Es52eSrEITUf/PgSxHq3yJCPISfCvSr7aqvQeAxnEW+w3ve0b0Ni8w2oEUO
3oksTgPrRadmdENjE9SK62FK88n1Z82zl08cMnLyBeVwjJ8qdH/9Cba99cOi3Nf9
sp5wQE5tr9u3INDvvi4vuj1Wb/8nYU7q53G9oknOdx72xw5XkSLXC6m3P6mac+fx
jp0iPByBVQ65P4vbBv4Q1sGOI2Pu2vHQeUTdeZKWOSxd/yd5GCWxjkJ7W4CP/MNu
q9jJOCHKdWv5Fv+I3LHC21cjTaW268kSUJxTHIiiWNSYBfELAdythin7jkcq7Kxi
4Hi3TmXlGA+L46yviBIjwcpWeSpdtrWK0z1z30o/XVK9m03mP7AZ058nXfV944en
YIvY5/wckizcRbSOwRHoBE6vDNaemupquHxKiHy+w4jIOWGKfnQDSYzyvUxjAzSs
bYCEp9wMGnvQF3WyOoa5r58TkdHvnkk8hw5JEBgRAiHTaBidonTShHZ1Mh1dYM31
Jv8BHwqzy+MskYwTV/saX9QwShYebNx/eefkkdElGn6YZ5h/6dcta0G3i3jDlOwW
fIpo0JMmmzcCIH9A+WJiKzZz+SJkwXWgr73iCEWL/qyYK5uHZznjZTP57LtrfIAH
NFnw3EVlucGVhyfFJVsbzgYBcMJ1jqO+Yimw+H9CB01Id8EjKmpyF/uvNDKBXxue
6w7tRDSdUIMnL0uFjvNcT1BOKqVRtzM8NRrkW0AvJQjLy/xPgK8anYBjVDMC6txv
RN6Y5Skx3M4RwdnALm0wS/F+4kg71KGCsucNtwNUSHfpEQb/da6CRN9mYJqr+VGl
ok8rel3MHvMenYIX+Dbiy2dUNYXO/CnbOGgaPSGMT1W7pAkd/Sh7mRygKD+wGTq0
zyYqpjnUmZ5iPQYikjFiON6GtYNKr3/J8GAcLVQqZMYLeW76yMbKDm6Td9PhkfZj
iRqgul0BQg9iDauDYurkjKmBNc97hXGD2cJVCDVSYsM5Suj656uBQmw7omPRtCl7
9mJUBOUvxJ34nbLIH5+vMX8ankMK2YSHN4dalmTR19cij57NTOnERiUGTps8VGi4
NZbqazDmM4E4GN2aqRyi+kXmrwAikH62Gn2ftTDnFawzbYWesZAmexyfm8fP0IAo
8S0TJ/5Mv6uLrH2FtHAhuCzHlBWMM/iR24TqGAzYjGje+e/sjNpo3Xmp5+3BYSqN
njy07l4Ynr9q0FjlHRfd2Ve2wQ/OklmtbGoSMvA8Qxtuuu26+J6QuDTQWeQ0O1Df
OSi1T9tCuMykDT6n0IpcUP9PY3jOPMehWKUCD1YE/CHB9Kaf7ZK92u0YESJhmNIm
ix/e5rU6L7somJajrj8EbgyXDXBkf0zcRGpVBhEolBPMSMYYKfsCAvfONRET5aKW
2gZmdDOoPObGnJLwEwXPoU+ZXrhvUAPG3HpE9IPw/wRsYXPCeesQD9AEmGef+GB1
GAMC/C4sIyA949kaqkGEGHxgNubwesUPmr5gAGygSo0nBt5I9c/NMvT9Hz/izyGb
OxycheNT9oyf146+7SKL7I7Lk1S7ZzL5o9QWK00g561rOD+K/7wNacFtv+ycMEe9
1LCoeIBFgTvfijvPmulz6kn49El9nAK/RZeElAa6Ryq7BLYiAPzlkHr24qqPG6pR
RQaxe9KBHCeP1ngONaZu3wR/h9uPXk7jn+MzkA/ByGFjcVBLZyFzAXjSTQcHZwn2
C6PQWNYp+2iE0nAlOZU6mBWILxYFRbwSAdyxBDFB68MSaDgaWGTtq38JSzgObYYB
dZ6ZnzphZ0d3gi6mz6DCkPNNlJ44MI3hvxfVacd4FyXu+OOvE93Bsu+5R0v1GH0W
ts5jxVzy4dGjkGOVT5VXjHI52QjjELBgcPHpYSPBXlPSIgmJDuDqMAR3Va09MugO
/TODJB/vDOrL3ZSf5LwkHxFMP8n33tSV1dwecM9zq9ExW+Y+J5TlAxIJIvJs1vqy
NdJ0VlBhDSChw0CaSX3ddl7bSFcT9LXhctpoWDiS3fTU3WGUUGzaLC8TwbixiX/d
Ny/KHLxH3OrpKQkUCXnyjRYjENqBm7vW2MfeijlYXZQVWIW06L99FJHOMAQyBBVH
YzOtOsv+oL1Gq9I3OrnwOrloZoAX0ayepDhQkSUBT2dn+Z9J6S2AQMD4+jA13dSo
MT7ZnLtyakfip63/dwbKBGuw96JRJTYFjhRQV0WO5l2YFYw9q07Ec+EwHWgpNv8K
+iGoJll9s5TpBI2zStRpOsyxrv2BWMsTKzJXQbkdfdIjZ5xNGiFh8vt2cx1/FYVx
aPyLwhnIONnDiVmf9wipKFmS4yQ7gwxM6u09EWlcL7qO6JJhJJFUAwvn0FISvOLt
s9+ekw+bYfpF6oJp1/q0XsxL1tuZ+x6gK4boo3KRu6fpHIzqPblG2F7KXqvL/L1l
V6HPvrwDOPARLp4WowZYXMaTLyX9dp4HMAEcl5/watcHU3y/3Pi6FQi/8MMgrnsx
GHwqhwboP8scjm14jvdbGNU81t9lrx4ikZaS0VENZD2mBBwv5olnh7Ov6Me5IWCi
O9t/2Xriqqr4wPTs4NgmQ/UiUQGMS+KJlwK48/Ywc8jS1eui7BqRxCqqjyMFSDa1
89UbN6pH+t+Q6DJj1HkbKiR34HZzOoRWT36sO+yl3msk8pwU+YLrCEZge4zCQibK
zjtVvCTx1Jl/0DX4h7gVhnqVnm7mvc8kyVQ57uwF3qdJpAGKiFPqvVxbZzHau2kN
f/M9JplRsChYoMAxQAV9TFtJ+miJI4CmZIrmqEJMAogruxurolUbyR5QLkPexVg+
aAZB61nDd3kGCuNl7pCdaL9kdunzM4YfnlDpK0SBq8O9rjNzzo2jtZpBsuDryBht
y6SF7tclip7ZAM8wciB8R0oGtx89Edha/qx+vo4dI/KYNfva4J8XMwsNNGjCEMz7
8hENW4GB+7PHGaHBEA7FX6/NKBPwO034L7Crc3Ozm3m/OKKu5ZJAzBK5U32VvYyN
ENnbhRNU/HYvA5WiMg1FzGAyTmafXYOR4LOEW2k82ICrwoZHjQT8eKDoX9IOzAZu
VF1PcCmQFM1LcIEjQzcoCDerZ2eNGr4VM+xgBHMtoSWSN6TsoXdV74mrPQGbkqJS
ckweFmEeDUUwxNtoZcc8s1cUBw5vFEQhAqPuou3I218Mhigm3jityPxbiG66VlX6
fYzj30V98T8+luXXLpFShAfDqDWEFufeeVNvasJqLOpoPlKmtk0V5m4O3oX2Coo7
c3zDkslvo7S7NpWlCFhDOZAEnzrNZkJr+TV5eraI3+H6jVXqEpOvGrCPU8O1nQmU
JWt9AiUOqlU3Q2LQ9D7jln5jU5AADYOgN3b+0U47TLe/YCBXCWGPW/Fe89WDFNN/
13NQCtdrbLNFA74xxg5SI4DzlBmSmdQxzJ9YurDSuN6RZfbEDE9Cm1jwZFLCMGbu
5HOPY9QS0/+YbKEtGNumNS6o7Ihl7hU/KyEZD7jmRDB9jK03Ipcv6hbzDx9faet6
27g3LujiImALSOBTAF//+gz6i00YKwZVE+qX36clNncWQxrHYBK+NU+/rzBu2bC6
SXpmj0cS9yEHi+rb1Xz7L4GjpJlVfHbVM3VjGKhmAFFR6sExYY/KYD7hXORkvRDg
OO/awQ3eUQgxi+A+7NZ/PbSDWGqlbA9ACHVN7oVuk945NVNyXhsIggYp1ribyv5u
P7HAXnbqPgZmDYkbErFT4you0/scGDQS5al+slDpbrNKvyYuXG9aSoTfUJbY/TwG
w5nbju5G0HkGJHLsLnmEWUku5ChVCZwQ/5kp8aKlFYXuTp54s1Kyk0UScBuaCNbU
mDFDBZTZ7J1pJFYA95ZiCuqxwoUM1ZJo2Ed0PU8HCOwzrIBVjMOozKr2ROEtozu0
oR5iNdwF13FU+0oPZLkCJK1+7qBvB4PwOfzdfMq9eh8Kng7TOq8x7cnqRYIR8JgH
a+dU5Rv/J+VJz2kiNbjPhpVn7S4MU/UTs/PD3H/G9T7Q2Oo9XeYtONNkv+cGNTcD
Wgm/YKOfLkVmy4QtHBCRwd1VHFGzZdWNREtIoHFUElFntxSB0jQNe5QAxlGzWAQB
qeA5nAEhnqnpfAvm0M9AHUjNprfP+dBslQsIJXtImiyz+yjACha21LYLxOwsb4x8
eHKvK2k05dunh4XkDlCenHnGY+nP2F2gCknkgJU3g2Jn7Z2eL7aT0YznF1s8QhbB
hEjxUHzfTLa5+m/bBlDGJvpWKS8/OQDGRI1JCQ74cj6A2YIVrRx0SWEgQhJGt7tk
pgfYKUBq1N9BB55GLcYX/W4hRIgmU/ps/tYNROIaToZCr///Pyyjf16ZJ7d3UpnQ
SjztPCWQJCD8aQ8AffKr243ZHtoR9mWASJ+TvCbT/97V84Re+eNBuKf04eCDRAvt
PCg1Ty9bq3ZT9PiCZlsO1ba63QMy7Hd81KD91h8eYiSPSPVhiZJberNMAQvXoGQ5
ynOhrTkVp2jzGV5tJ4xNqROdfFfZ/2wqmQnsiQDTgMCJfX9HFUPPKMyt+2gMgjIv
/8jiRv2Ym9mwWePTGce8bJlKawML+7e02SHT77lyQyAPPXrvlWGi5JhiFIMt4miI
3vBoiXuNIwbXiC1KTXsyyUU5SneZ+aTCwzxMZT93AzXm7CpWLvusOYIBbA5d9AAH
hvjcmU52O6E77/r1+RRg43ejm/Flaui4U0Gdh/WAWSdxX46WrQ/x1zRVqvLEa2tI
xaef5KFSbWcsGgVolKezK4EkLmWOHyF61yM8Bul0wo4KBHeexsc/J2+5yA43uxlf
hWQmT2jo3fkBn1dIG8l0Pr+be1L9O07stAbyCrLcFptjoF+afpOPN31wbaMaOr0h
CHzd7H/dtXNJscd3yKSmbeBQStrVqfC2Xjp2u4qT1C8800ekBCUIcJY1aBIg1uh0
Cq75ODnLQKLlYf7tGd8DvjQ6YWmC+dkihghQwmwUaiAvzlPDqgcPpl6AWEs064Gj
etkwrWPfN0TfX/mbO0P8oovmvDLUsEqGcPpUDj+T6agyjlpJtqbmdwtzAFTlXLCU
UKENcBoZDN5e1chYxSWzX9O2pfGI0yr1wKMltMbOiIfg/jopm4IPREogQfXU9Y2H
FeFQgNiOU9vAVJGcTLjWQCyiLUIqmKTFElhCjGh3TW7KGwkHH1PnXSzIeZxapH5N
1DvGqCacbboPjaF2HpuqL40eBopEnJT2Ccv4Kxqh6Jz+vcsQdtwWN4vsKK+/kFaj
URke3SvvjBX6yiTrWMMaA6aNPD+wLGPTet9DGXWGwAMUCBtSpGyiYM5L/tS4DeTP
U3UhnNLEbma3c/4E51vKm1nOG4hh95wV269gMkEEJfYlodUNQbQSfxYqobVhMQts
VpPA8/KRhJBR/eTZ3OvuXZsbknQVZGYi6GJVlGB+jvJ/dHV+AaGVdtlpCXj+OlYG
GnHpLoyc1a8Ahg97XYKYDMeqg4pCdpK0pZ6xVfGA9Mj14BECB6COx5fLPAT3YfQ5
I+dgOT5eSylAW6VRcFls+4bUq31u0/Ekps7ZdlW41Gz6xgJs37c7iuSosqujj53z
1MKcN0kd7GjXSNtvNyKN3eKAJQURCp9v0stTxMMmXslJ4lqid8lN/hvAJ8f6cpPq
TJcnoJ9jaub1dDekuDPYu+hbcNZRwfdQ1XgD8bgpfLssUquTrWhA3crgE2SH7rHT
v0BZ+I5DN5NwYHxkNASRzvSpVHJB7rSiwcI/h8u41XGH/54qwHs7ACPfhOORw5oi
f5CN+6Ik1VtvE+CfC33DBjopfo2DC4Z+QDWIK1AROd2U+gBefoYQb7/LeUu9Fsuf
LU7CIvcMCVEkX8dyyFeAY60hpQ9WvW4AmEnsgYUOP5uODSRe/WILA0muQQYFR+1O
HMkN4zXQGFep0fHS2va1AOfgNoalRg2XDZz0Jch9435IhJkh375pNfKVg8E9OwX+
83YvpQWKbrQTVFMmVG8Y69bq5BMeiuOisz48ERWCilmqDm5Kwh0tl1pwkMLaSwec
AKTm/V6tRuHcYIahawHw3QCsHbPX8cbHoLBJwj2DpnXIEmlvJA74VYDOBJNzIHft
qHL6IILPxXq3NCO2h82jqke9zx/yVuHFTfhm2+gXap7W3MIPGV6zDB114bzy5FVH
eBGwxGmcbx9QHkywAch/EAKp12h9Uj+Ns1zPvb2RocjvwJezgso9leWhB8wJsI0x
JpWkkic5Xntp5IBpu8e13hTDnrLra/OfLmjvZmIUTQxosEv8pn0QtGlg19aFns2m
4b4UFy0YMXqMtjPE9A0PYqlIdFotpXlutlbDi0wAfJ1HvOOKVvtge9eaDQwnPGiu
XICNkgk6tPeWvHmY1nz0xASlRTJ2kuuDzLSrdAYplRFHaQsUWpzIBSLJhf1jkHj8
tl7D5MGyl1LdXd0XwdXVTyrZD6Z58YQdGNRMPiziLOfVVbzrou4f785GSSPwQ65J
o0nX36lndDVHbXutcCrhciyjvAwddu0D24K254nkFRn0RZqEIvh6bn6i1UOOVQd6
Zh/SbFEr12YyV3VekTC/4BlUNtMtKR+7Ly19U3ovUokgt8jOT+yCbhrXeG9/7tKS
AWDLOs0WX1iHwZKbKubRT7wiwqwOt1OYv0USDDWVYylbLNoN2Qa9/jZIqpx7B/zk
E5GBMQlb5KxxPh7s32L8sK1lGfd4R+Y9vz64Vr7xPgskSxyK5FnUuE89GzjobAXu
2Fx8d79OVT6Al/0gB2hR6K1DKT60x1zceQAvslyVjixj1VJuX9XbDI6Jn8OaH17p
6qcwdydHHcjzKiKohhIsc30pOgP1/iZNrDrMTDVL9AhMgLnVEj6Sw9VmUIMPtsYT
rGGgbRgJ9Fx9tWErmKG1a7CO85fPo0gypveYJKA3vAx5wa+URaUnBT94nI41R8BD
5knzwiXbJ5EcVlzDX8IXIrugVp2ZBLot0gB9KmXm9L6b3HMp8dUsEruopCyL0n1P
xZznpW1ZtQHhieCrvRygv7U33Zi1m35km87sd7coY0Fa8k9kK3VuzN/h/ASVSzaC
AQqrZ2/7S2qIh9sPDb+RwTPflSd8UfMTxMkHvZZJMyxGJUkwLThadCA6JHdq0oW0
Njz/dlwX7565RrUILvsoOmFSdxncFR0XU96XCrb4EJ8ovM2d2gLVsYJbExm0ZaKB
qEot+1ZUbu7hx+xVhomIRTzcE85HmjIpF0f4tG7Jof3huruWuZcYTfXcWDxmn8VS
58m8S1Rh537YKEn9AeaShonR+hSBMBapL/W3txnpj0HIFxq18jbBCK732RRixqy3
hysxVgH8GVJJlSukBGSbPbe8bqq6D4KcFexZ2nDifioNpRXKwsZ12ycmrdS4Y/wg
L/Px4mmkZ++2+Mtd5MZIGWITkcQZ9TTNl2Vm/Q0pU73dHdJCl97kHCWyTOQ2Z1OW
Mi5Xf28mdp9hCf2IatbSyMPpUmyejQhfKB0UAEOl2ejs4pjjZakopYvl1kHCIqnm
eTgL5Y3P4F8qDKSm9QpuFNJw1sEy1IQWbpCxmho0UorSyp3chYk9xtICP1/Fa2+i
wnXHF/h5TCnmU/W8hc6v9J0rsKba6289Xj8oFVR16BctsbQXompV/3PhxECnDuXZ
NCJAO281TPxcgMeQnp94NB1Eo3h7NkQ21S9LFbAaj4x5PWavVoD3MRtcs6bCCmML
TTCS+bS8zuSAxhumyOHNX5rEXa8fgJwmybaGHEWZcn8sKGj/xJ5Qh1pnU1VrMv0z
lFJiqPTRh85SGKbTKlasdTDeiB/NPOTXokWauZR9ANyHZu11WJR2QdfozpRByV06
O/rG0PU7r/ejJsTJBuR18WoCZnJ1mJQxW4fZ9F/yMJ6oNVX/X8NrfKRZ24OC/ReH
4ocG/lim9atc9QD3QsX2U7xDh/216KAUZeYBFb97fcmrDWsxgFuWFDTEv7ze44Oc
/7ihhS28n9XZANsYh2SMfb8HDlujJ/yVBr7oMusXAUwoIN+VPRtxX5kAQdex4Ri+
RSsRBkGFwuRdJgwbGGo+zGUpSP+pGIchfYoLnTvO5hsDqURWbxywTHXDU22S3ge7
n2rdv9FjlrEC+VpNTCqmOZlitaKj9D2SNlqmUw4X3vcgBTz1QYLqBbwdgTRyAdjj
IbLLpeZjXKcKyp6h8ypDlNwalMkO0CO2kJ6Y0yuYrNU1DJaMlHIe04WLErQAznxQ
+/eVVg/m6rxU9fq5ch+tdiUzl6JgjiWtsK9FW9X0xmP8ESoX8oSKVhyPrTP6cMHh
yY0Yt4S9XqrrllK44kigwABYbyQamNqGw3O+cEFz3qbhcpC6V1eU629JEaQF+EzG
KYh0PjKtdrtOiiYxXUhNU7cx1wTG48fNfPtvHSZK+z4h9U5otmjcstWs4tavgX+c
ByPHvQRtfG0UMUoVBQsvbCfARsXU1mqHVX+s0pxKPOVDJMaV4bN6PQPIE6IQrPYc
tIPBH6Cvk8Cy62/DLPU9jKQbeC1ZRoj9+odu0RXS79ukv3CHfZo/wrJ3pTa1JkdZ
VKmJnQyniw0Xe/hr5Cxwjr2qjGt6YkbOaWBKEW/i/Cx2gE9CiGSlLbVhntpGTBYh
1tv4TJl2mVsD1Itks1g36o1wgMWrnNs2jfA/hVrfJS4vUPyt4gah24vvHrsj7avp
qhUXJ0YbazH09MP3ZdUZWXsJn5r595l2HubgV2PopuVrb12sHcoZcHMlTmBwxWSX
QDAspAWrdrXgy32ufpp6iJ/BnAFMdK03KCH5gr/tCPYBI5e/xY9zgRHjtoPtxewQ
58BEaCOM9pc56huE2GVwWUnCxymi3EyRebrhYT6Gs46kx/aBYHk0aPh3G7u6dnoG
fIRnQD4xWEmoQZLjhWks/8DXxKLgwIyKu9lakDHQ9rvTDww1kH+S2PDEp2Ky9Jwf
eFETAS30ptayzKcWaLwz0Z+oJIXNvX1lcVG7avbkgeSoMLHYx3hLD2/3ZStVQD/g
wIzvPy6mjBt5/eip/DGU0PrFX54LzdcIjviDJLLSp7O4xHR2ld0QBD6K8GJkIp39
ktDUNvGWRzLN4wCHjAq/PHgij7nRwQdeTkOXGpqYtlwATwH+NTSI6ivWhGJa2J8r
vR5K5oj6/vw4qmlqCszYBaTMhpiUyuYxUl929bNPd8QRQkVNLH1IBQ7f2UbpDORM
/5rJjs3jMe+r4VzLmG5WOr8qi4BdkuSUtW2BtLiHLUMKfUyn1gD1tpB4NDjWVC6Q
1sqpQz1AGbZodX7opcoKFIz4q6nXQboHXC3N6aVhOMaNKGkUDE0ac5CYJC+GOemJ
dWxEGTPxMCe6CIi2XXB7eub3H9A8N1gMRnNWdLvaK2cIPJDsNTZ8zupNgmULDKK4
/jXVCgTZ/LxdiIeDnS9UByqQFrOX7jJkMDEKSkteb4M85hw5NfotWbECiglV+6jl
MmZlpKH7JoaA90jR1lGtif282LvGd4GDwbI7vgE6zDRezWnybAJyQipus62wRge+
q4hakX1gWvJxjoDZwDRlVuSVvjfSuZ8Z+pPATELrMWu3HnL0qyMNjWhYG2EW7JIB
Z3QAYUj63QPV6AHmS/wJHU3x5+zlCqQiv7QOR3X5kMgiIQdDVWGMcfwYrRSvgKJU
kbr2Vyh/1kqBYyBCKJrYXg1p8PJshTVpvbdoLcr+t3JGUN/DWi6I27yVzVtYXPam
AWhbfcSJv71xvb5DaeD6ehsFFtGOMD43JILPjfxF1Gtekhb2fNtd4HlOqEeEXGx3
zIFH1I257BTRDmLW00sHBYdrP7kuXxurLwgn94ZWtcuLza29jul/fx5crGUY5n4q
YLej0nUmdDkFAZ30YHNujdl7Nqds8T93bwVZuEI9ThhIB9YU2rh0xFuj4iMKk+/S
/aNzBZAG2ygr1qVD8ZLBSMLTPD4GdxiOL6Eh0E+3m3YGk6c6Fb8W1kIkdfJUtReo
jjY6YzsiVi9ahY6p2z9h3SLLpvSn9nvKqPHsEaN3lBfPdCpPrXT+xAshVj0mLUG3
sUM+7BA6fYNj6v519TvV5H+1YAywDObsDTDlillZua4uB2dGgQYm4+JpqSqUKi4/
kXrd1MrAozSjuIO0q+b8T45urvhmz54gX7HsBohAsHWNLRZ43jNJj+7ix9qmgy7b
Y4IkEykaNK3/A88B346y4Fy3+yZxxFfFsv+0elOtUlxxURT9pkdosePH+12+m/CE
1l5qeTd+DELqpsJzaV2/uxAmp8jFvn3Qw6062ZbCDpnEDPJaOSub2J6nERtTxs6q
2840uaSDp5vPYunqQ58CCIqJ5LisvbaElmvtdv1732QNKVc7jbIp+IWDgfcPsZPC
DEZ8WbfGgzNTVsw8qdueiMUl79NNNqMXCmkDrBTqe0eG0dZwVL0fGb4oTFHwR4lY
cTcshc6jYeBK4RCaOanhdN5UwwlvSQpV8kP6ZBHJ7rkaJ8yKsnYnApiExiiNxLWI
+YTxOUPv7NhRD4QSGL3xP0XFiAxF+qeiJuWDSjhmHFP2sBFeT77cYLAEKEQ6Obf4
86QQwGZtcwNypcS0sru3wEArwWvq659azbXKUB6UoYTny4BuVYlM6Zqjev/msZli
CfOTIQDNbhxhDCSPFKFiEGKSMeI3oG9rdS6jY49loJCjj2D21uI/P9LyMg/2bIud
I6Sv7rWsNfXFMBZD+kiD0QZMQCap1cy917ayy4aAbSIL33TCHdi8sP0be7B0uIH6
Dz8yAhMHX4Trp5LGG2G6oP6v1GuQEetfGIs2AwB6z5zyAlvo6bADSCoaE7zKjaVP
pGW5SYDalqM9Q7ZEvT25IWAQ/ByDKUyN7xOlcWdvFLCEcffydJvq/DoMdj6yLrN+
Qv6n3SeKv6r31UzzQahVDlYSce4MVivAvT+FdBX57uH+wW47I6tnRl46PkQMwP8T
XNQ5roA+RwFEEFaax90uHMwA6ym3dEqB4K2LXJT3fqcpgRomHO/4s7Ocy+oCYSAO
5KKN2yCW19WOacKajwr+YmOH73jAcYuIVC7n78N12OSFPUB+Ix0eCE8Oc2BpZg0r
9feHKcOEKYyvenlncs7DKut8iE7yFk4hLGKN7DfSs/1D4+BYODFzj260OBiQVbVq
mJGcSgCBpf8707XMId0o3G0cSN/5cPJXyOOUM4hD46fGd9Fky41DZ9930TWHkjB4
lIAGDKpIPaCAZ/2yOuQ5gce/ssxShpGkViWW2UkRnx75MX96HZbr0bSVkHmUperV
cQioUzPDqOb93fs513NwkldKJo83juhRV7qYMHfvZZYZFBroIbmLt4JOV5TgpL4/
JPlA9+6uWBCvehbIVB7ZdhKVGEEDSc+bm0jBBrCXPr9FH18djlkweLGnU2T2T+fa
SbZ9JsL6x2gh0A5Ibl9MCZsePGnF/e+JmaNpE8Lt2F/9+N0dckhvv1TkUD48Ndjs
qe1vXB51/mKO9BkvivsSmZUoersmhRVrWrF5+kawaEE4/mh8hDjci7fW54TFgCIK
84tAOwu5UahXRe8r08GGzAZH7vVnaiBW1knEfCeo98JQ1TRkVfq9ULjAqS4FCX2v
2DfUNpp+5jNE6SkBMQNgoPHvjgbUBJdFq/3fluil7yntqAbQF3qrb1hsr28EOYrk
20w+Dh7AWN9BV7zXwjkU2nWnsblSOEComfquYFhsfE8TKWIw/klWcfzaQxphhJS0
vvoPBsT7K7ZdE7FzFrL+ctQRYs6oJZ5pEgCbnYwkoqlqjHkfNslEUZNCcANB3wj8
nm34CtjY+iFUuq+cFINV9okIBzOBFT4A9iTTWWcBdP4xeNvbxeb8c5gHizjlXvTc
qghonxxosgBDktb9ShQbMjzibhGSPxQPT0ezCOrFO7kA9zTmSzkOkdFnAczrTm5b
NiOu70Y7+9bDK/ejc1WoU/XNFpuN066L3sm0QcAniQ5eZHAXsOK92ypUVB29Hv9X
qpkNoiEWlnbjA3gl4cXZkLYn2Z2YyO7ptX9KItB22LZT3uOlGc+U++1HjuV5CSyQ
QR8ex8gMNnSQjAOSlVVRXOp0wPKTxoOxcVF20L4YjldX4pfCAKirIXQ2+DZA8gpf
GDUKo8Dxz9YPTzcPizm02TXGh+slsVMPiy2V84hWK+TQWgX10jqRdNDieiUi9A5m
D4vVcmGfTVbHSttv4Y/Z6PCGBR4rYgwiezbZjygUOvIY+kl8b6w2yJE9a4oS1WKP
ts03MHpmDYX6bPuv7vVgDscZTqNf6qEjnWsaEkumNt44ZxLzUtqabZvdlnpVlYiE
Cvznp28SZg99q2PbomvZAnz4XukicCR5+AMAwBOAd2eT6o5mTm5sPOGU6Z++1gHj
NK74Sxo5LnercLd3BZ16NssoU+wnsh67b+AC+XVls/NEV/L9ORUmb3lhY9qRwlIP
k4FjTqbI5oCjSW6V1wySgOFPQ4jtSa7fg6CCzOPhcAaVb9vNiqy/OnUG0Ur9Bm4W
HD8KeeNUv/vjiFRkp/0p6mp6aOE8J4o4C0g1LnhgvVDHY99FvptkUpfKPYKABGTR
z6Eaok6yKU9LBUMJ3vZlBvnY5NesXqyqNv2yERLZWxAl64CGGZ1wLRfygHm/YPh2
VkXiQfKgMBkf0drNleZ3z8O2Kc0xeyrbIIdaVsoJ3RCzP/melHYtfV7zdDsOGzCZ
Q68HdyTj6SWJQQhjBYQIiVUuTxsfBxM6fdKkr1bxEfcw1KMml+qfHZIdqBtUEhHW
FgrJCfekLLMtTmPSMEWcI3q2pQJixa40HIbfixb5NK+P+vVGpWcW05wNu2smI2on
r7A0fGpWzjXwqjvB9QP4ykgZxZ83PryEpR1HhdLe7WQwRCxTzVugqqrubKdYdhF4
I06q8UzVMtyRfL4DQa1/cTNIhczuODzWPXdXoQ8ThKF6nrYjg8u311QTZC2YHUJc
DVV1Jk93bXzLTjUvXRzMMWhzz7KJzilwPV8xCQ+/es1VqyqcDeHLZozfY0H0IcXg
vDbc92BKAv2fehAsV2poT7G5mIBD9GKNpEY5JCZ/dSSEDaVaFNdQyRxIWrShaGql
f7QOXy0fAPbhiq8FuPD7MhN2yAveUkvZGD8l2c8gS7zR+2Vzu8hM7uU/4pFqLXa1
EjovS06t2x6dWHro9fsRY/fI4u8b02GpwM4v8UgWtgCM+JhXJ7Ylesd4p0/did4W
utwJaaJUj/KScBfelZp5OaG3D1Qwywi85lwIJfkrybJqzwaEv5i/UrkqboN1ZbVK
QXx6CMeoB0EB8MfgncyqFqBeVTqkj0TnBridmG+hxJzgmc6KW/s1sFljKLdpZ9CI
Oe8dgTaOq9rQ+hLGLWcQQcF5l2rorrgi4zj+k0+bU3T3rJ2tCmTLzem2UX1ajucB
tl8Nmv4IE1gzE0JwIqHToBPQEN6QeEpbs8hInWXlpzZdUOlCO0AwX7uwynOhp7Hg
lYapKHxiYjk/vSH7tPDdw+KVder0il5+bggbx/3Y4KamxJJWANxEK9611kQkPB0I
ku80X8jXh4SHB0Yovl8iQutITqA4HCGUglTYmpKs2fj4gX3sUPGZxow81dOhWr1o
nx41wD2j7OfDaCL9rJNol/4ilQKfmjtHmbsneYsTS/K0WpH7WUYvNlTxf/wmOGp4
hTI5OZvs4gPO8G4myE2J3zOkWoRTodh/YcyP++1WNqqL3K/0NjYSZWtD2ic14moW
zz1LkLGvFXXrP3F+YzLtDRAxUhPhGa3V+12ZTqbxkPhp1d3iHjV2AWRoI2VAY5wm
/yXFvGAmjplvh+3UCMTH+tyYsrx/va04vExYobUsY60DvARvqG8DifHBhJoofMAx
OGnTv/1Zn+8HBB0O0AthE46/1HkxZyLlsX36qQDkCU8ZxceM+gsYuyGxviBqrLgp
lGYjxYzwfcYCoBmtQrINB7bcHRe9lJJfKmmeIttnnbO9youA3uktznMlNdXe7346
Tn00PYH7dKQATacmr9zjuBN/acxrR61X7c6b0tIyrDG1427jx5Z+oUDtabHjnKbB
X5k30rUI7NxqIX/ECyNB7m9DgMgz7+m79NcAj/C2xkAc0KzrMHovTHcEkGWfsydy
V7J8/k2e8NqThn+UxPxlobv1XzHUeMdVea4QWEoXg2ye77Gjr3r48pB0Fo84Zub0
zKSKyR9ImCNo8TMeY1W/Kp0G05hZ+uoNynRxLfdCKiegzxBRbRigBaKQASU3RaDn
MYd06rP7WxT1BdY0hZzL29yHvEswNAmOS6BJw/G8VZLwnLBaqEQ7jFv98mZD5mzQ
qtxLzhOqz9nMxxk74yp/dv0N9q6aLIwBGJpT2jslKX+mk/gEokG76130pk9GNNsf
boSgY4rwP6o3TnMMmi4qQlE2g6jmXdKV4yOlD6wi+G2z4syDBk2KfIoxqR8XGAbq
JSTS9K8l9BuBmODZfBJBaPMSDdeqHZ80c/esphnIHIIqtJxeff/q8pKMj+Od4Bj0
7AioT6rSwEKwlaWWujzoykGWB1/qHKhOA5IG4Op29yKNECe20romFxZDqNmV6xd7
NEF4DUAQ65EQt2hNXV3zpPTYclSbNYxSjR6fcIs9OnhRQF44F0koxsyoc3ajqN69
eJs5aYnm+IM5Bzi7zICP681+48crnFsy7Kuh6qZ+BOpc5vNoN9t5FJhHOPr5Movf
7Aybg3GW3B+GcbOTpLd0x4CCpMCRRl96pGGP9ulN6IcopuyLqO7oRyAtebmhndHp
rbyVJKQRNGZ/51lpdia9jPLzvrQX4/YANBar38SWIa4oXxZN7mkRWgQ91kC055TH
ejrblFezmberPRJj3ibWU9K5W1KaUzVomx1HhtlScjkUXQQ5DUuxD9n7JSuuVUsq
Z7Cr6m0giUiTf7JIjUdzCH4Bn2mPpHvb2sBVki5QEIid0y0IWXg6NbD0j5bauwK3
ovk4W8oDn0nK/sdGBpgxgxlfQMk7rPFkIpiMj7mIYSKhzcsxQvlY8PAczIO0JlIo
Vlqtet6FC6CLJd093JeyiDFKE8rkl0Puoo56GZXw6oeAVZUisxtrmtzuowJdBVxm
ZNMfxSyMxwbmqkle6WUgk2RxRNKNtFLuwZmt65HFtb4LzY7c3Pvoqqq1oIgikIMr
fHT9ixyLrpuWHvE2yf/BkxDBbTQxWVM6TZJ/DbMQVU3MYnmPu2gBaLnhSdV7ninu
UiENudHakKOPvGfkFqhpFAFnWdhRX2K82e58oa4pd2Z33zsrFizPvauOvacH1DVZ
neddESeiLn7+zfRP2lw9WAIjjmYR3DSngQ4EO/F3KMNvG/9d7FgHC5S20ZJzxu/l
WDFqAZ9QYBE2Z/BoTcMeO8daxiN99HZTBA3/kv3QG7TI6FRMTg3qMnF/mN4XMBU+
8JUOyDAYuJWwHyigxA4QgUJ5a6zFt7JRu4CZ9qsUIyedn6DFErp0EbjNZoL9hG4G
D0E9aSHeTzbmXxGp3rAVssf9BFoh7kBEml9pROrxnYNY/xlc5cCN52DMWSfNBitN
bw00a0k7aMfSCsBFZKaiuTcUGNa3tFsgn+6zqG0fPkbw3bkWnWSHT2AJ+hfgX8kR
P+eSyU3hnbW3DPABmfesAgtgrsBCaf3cZUWbpbRmGbCs2LMMXhzyPDOhYYjnqRiT
Y3XU6/HfKGsUQJLmOSUSg1ckhw1r5YyUshW1Imjy67+4WWxY3D4RzUQEae8CjrUT
y/TsD47HpYDeYYLoP2nIWogOYQgFoLgawCGW3pJiTQIniHuPWmH7qMFCtFfJZY8m
qyfZkcnMqFaivdIRyA0cnbkl2pPfdZIT3CezrciqRmB08NUFBCv3JoAywnDL1J5K
p47JjC15x2o8NFgg6k1fPyGriExTf8aGJs73rRQr4sZ+oLxMASx8i4lfvwd1Vo1h
FFxJhTC7GNB1fXwgAuQoCogTFwN4XoetHkeHVcV6+r2PJmX4di+oayGVpidCBHH/
tZVec9N3tSmoR1RQr5DcbEyRf9B79PxJD7Gs66t15WHcYhe4scC/3gtVFclgczQr
NJaCfENJyH6Pu2mvCptKhaWpyOUEIN1oz5UURcV8MNeehkznLyR9Dj9xbo+mPPH/
AyKYiXrk07T5cdq/HnRsqmaErQJcIO/X0HFFK7cduXGdIFCg8BZ+nX7rSrdmbfGX
EoVlIYgrKTh6ts5sRujepfMNoN8MhxVce50oyNXrKut3lBaNy18LkhGyJnBYaOMU
NAAmm86aZlT+fdKfeF5evFHJKtno5PNv1GopDdoPVG3MOIV3xd9emhsjxl37Swhh
LoPvNkfWFWOjLzrgVj9DEsTiXFJe/eelNtIkBlGHqn1PRrxOKRFdtCaYcCnmuc6u
t+cOi8rex+Xt99CpzwvNazJNVf9B3uaRnQ5XGekvn5K5q4vi66G0cu7tfW1Y7fLW
18GePCwaNKnKRXyNN7IcijL2QxxznOgDnZlw7LlCuVFu2Kka3jdSDpF+wXChusy+
RYh8QIoHwpxjGaPk/KzinKoR98e40m5y6T5OemS2KhWnW3D4KcrTLcZiA+vJGp0N
RuOe9qiH1xVGcCzlcZtOkrttVSuyw4L3lcd1AbM6wEY1z6l1SNkMJT9HVTIst5Og
dRCRl5032WlKBWA7kzevikKVpwQ7Qs682t5WPIr1E6hs2IXvlhgflaPmdMydig5X
zQHu8zSSam9QGxC6r9eS0Kliu/XxUQ1BsQar5FxYUztCiLzBHyL2E1tQnM9Hy4+a
WRyXum8Xi/wzCVecBs0Eaxv4R+NIKLopyu8EfR//7X8aX7PRZJFtbb4G7+7JrRUC
REMOT8kI/XVKLUvXTczOLw/8lCsdpnKG7XAnHtGwxyc9eEXS2C3Xe/TkWK0XAC1E
/Ke9mvpx18g9sp4V+CP9fpcsmzOw+SRDg0fuKyBgry+MFfip3TS4cBF9IIoiV+JJ
ZkrifCsmSAfWzD6CJFc9Th/Ok6mzLZYs04sUqYz8MMlKIrxiLdWi+KmfEqUQlYVj
NBNfWjPUs3fWw37zuaFjA6j+ppD1cAVfvxjiON5xdEIzU8BTBi9hfIdPb6jbbWJr
R40qXoK75YYdwyk2gIZx5S5/laQxOasJ6KRrv0TtuiLMCnm/z7aTmAuypsdCCvGL
lwhuZB0XKtsu8P15KpiqRcKCm8AcKsEbrRI+intpMXtxtZDvSHw1wwhH6cvJMpP6
m/qPHmi/A9q4oCTzHxB9GBfoXHD7+5YJijgF+FFAST/SriHXbMBE9tc5GdjUmylF
U60Th3MHTgp3c5m53IXBV0CVTTe4wdqNtmLoJ2VD3tGpKq9ezh9TFtmhyDz9sXj8
UtyjslnOF2CIho2FZHaQQWkxijx8mzv6fFwBzDB/8nrB5qNnOJQmuCTPtUHtsjLB
GK/Kiu70k5rSlgyou2hdvJtTytRPmdzzQ9z8NU6jLunPC+Mn0xNPHiJBlYUb0i7A
Ix/CBRyrOAG0k/nozygl+0pvQz06bJIvlCW6xDMCg4ZvDkBdTVmwmSIW6ONf3CzQ
OBtqVpZ5a7RUmhgonoujWt0M8KY/3OFMQ1ktMgFz5GIFkiDvvq6WntUCIv8hWmnO
wpUbA9xWUTiHDa+vkhLCGUSoeP0VW9jnVERsiQohRAAbZp/cGiI7wWWfrKKcVyuc
vSwCl6oZklg65rV/tTITtFkSxmxdenMru1gAvad1pugLQNRY0zAlyomKTTEKU9W9
IYFDZdS7YoWWDN5Bxsajnef8C5UQTmGU9QOQckvToqRBnPwKc2e4A1BKQ0lHFgY+
AqwrQABEl1o+qayoB0KpT1qUsaUGcFQ6D4tJgIXbVUB3afUs/lFTjUCskDq/l5hG
uAEFOB7Vc+HP14eY+rAoU4G49PTz2/c1ZSHnLF1OcBASOqG23AexxfQIv/ZnUS5f
4zSfy9NJ+NncYcvTmHjm2PapXr3LhUOnOIQtQ5fjgpWTHIZG0Rh/O/3RsEw/VCim
oATLMK9X3Tv1DxgYUmYd69XpSo+KVgcyME6xWa7ZsOeXrbxxiGdjwZ6jtiXoH1Lm
RBNhaKA3Ty0jpKIbW+xlzkduI38IkK14qDDWp6U3xxVsrxxU4PQGHk+s2DnVJ+ZN
U5/1icEIEoEZaY992+sumCGzI963vAe1kfE6qGybnv8c9dfwK3vt0ZrIftTyZ+Rr
jo1hUAc7DQ8wmZ89vnf0GReAWzygJMc4RN6buk88wR5J5BCGcpyHpvXaQWdE/b3G
gLahXziM+nOGcuFy0F210HZqKTBV4YZcwKvCMITJ8peT8Kv06lyDOeDjn9/KnDbi
fcZ6U3DMStMIIqSku6jkhSIzh0SjtWQSRunHroUIg7OE1ptBYcIRKXEv57TXPRQi
iOj+YIakjs4Po3HEjURixpb7mt6ns89zLqHi0/kIg+wHvxgfJ6cz22/hKDr76Z4c
hPKm1tUSR7QMN5b9NXgFUYny60Zjh0Szqj/xX25Z4giKlEgu5wCbTokKAChLWoaG
sPfUv4kFYgj2SMWm8sTayx7fA91oCy+N369kHc8sk1cz7KK10OC8LfQQaBQbkHDT
619qdEOhKiojhYpD7oI6ED62x37M2jKMndBS4cdKSXoj1hD447gha+I4oNlxXRXn
IIwwhtjeC4PBNkSUhuoVb9hMhQ5NWN08pVKsebuzXs2uxKBjZ360pxowScBgZEF+
Z4bR4TeJoS/BPd0jjWLdM0jadjAZAOBieV5cJR4mgVcT9MqaMTmuOVG5EmoXDGOa
+cEJY9y5JtrD9knqZhkfg2ahKeGo0sYonXvI8kOsFsBJVvRFzr0wnU0fu3tHZ5qn
7qqzzuKMAPYeihaDDeva+ME3bhFbbN5C4VyRBE8wlIbpFbmbXhgYqet85yjOGL33
eLkPxLnUrNTWubcmxwsb809jA1N2/W9TtwF69JURQLNL4SP+5mz66luaBI8yCoqt
2sCx0yY7LH+FLrxFo0qdVnZtXDe7CAKHiuBo/yeViSLhNTLyv9GRaYQFqVgr8jX4
Nr1rJcMT6YpCsOP67zE8tJIZa3gZxhxN9M6ZgNsv3SoHz5Bux2Fg2r0qpilGc7H0
u+TJosZ4sGxq/lCzQ1WQwcAoqkII8rbVCsbVnCTwZKrzMt1lUs6VTVV4A3AM/6ZS
GUdjP4avx7FWiLYRygB0e+Aq19WQbvaFSoC+wg9SAq2PXoRJ92rUBCrcIffNLVZD
dZ3qVcjAYkUbRn9ai6JZhWKQhr+g5xR/PKXPlleLc2n2mrgHiXwXLgJuIkyQBh9G
ATCZ0BhHYuYBcF1MlUCSPo6IyibEReiz2X6o4uF8S7C/3PFSqB9xsHUiVs0FFLFU
LdvnlYyNPajlD2T6TLLC/318UslajwrZr/m/7hiTIkyuWp8JY1TOdS8GIG2kY9JP
`pragma protect end_protected
//------------------------------------------------------------------------------
//------------------------------------------------------------------------------
/**
 * AMBA System configuration class contains handles of AXI, AHB and APB system configuration 
 * handles.
*/
class svt_amba_system_configuration extends svt_configuration;

  typedef enum {
    CHI_INTERFACE = `SVT_AMBA_CHI_INTERFACE,
    AXI_INTERFACE = `SVT_AMBA_AXI_INTERFACE,
    AHB_INTERFACE = `SVT_AMBA_AHB_INTERFACE,
    APB_INTERFACE = `SVT_AMBA_APB_INTERFACE
  } amba_interface_type_enum; 

   /**
    @grouphdr amba_generic_sys_config Generic configuration parameters
    This group contains generic attributes which are used across all protocols
    */

  /**
    @grouphdr amba_axi_chi_sys_config Combined AXI + CHI system related configuration parameters and APIs
    This group contains attributes, APIs which are used together for AXI and CHI systems
    */

  /**
    @grouphdr amba_multi_chip_system_monitor_sys_config AMBA Multi-chip system monitor related configuration parameters and APIs
    This group contains attributes, APIs which are used to configure the AMBA Multi-chip system monitor.
    */
  
  /**
    @grouphdr amba_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  // ****************************************************************************
  // Type Definitions
  // ****************************************************************************
  `ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname amba_generic_sys_config
    * Controls display of summary report of transactions by the AMBA system monitors
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  /**
   * @groupname amba_coverage_protocol_checks
   * Specifies number of AMBA System Monitors in the system. Enabling AMBA
   * System Monitors in the system also means enabling AMBA System checks.
   */
  rand int num_amba_system_monitors = 0;
  
  
  /**
   * @groupname amba_generic_sys_config
   * Enables CHI system inside the AMBA env by  constructing the  CHI  system env
   * in the AMBA env.
   */
  rand int num_chi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AXI system inside the AMBA env by  constructing the  AXI  system env
   * in the AMBA env.
   */
  rand int num_axi_systems = 0;

  /**
   * @groupname amba_generic_sys_config
   * Enables AHB system inside the AMBA env by  constructing the  AHB system env
   * in the AMBA env.
   */
  rand int num_ahb_systems = 0; 

  /**
   * @groupname amba_generic_sys_config
   * Enables APB system inside the AMBA env by  constructing the  APB system env
   * in the AMBA env.
   */
  rand int num_apb_systems = 0;

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_generic_sys_config
   * Handle to the CHI system configuration object
   */
  rand svt_chi_system_configuration chi_sys_cfg[];
`endif // `ifdef SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * Handle to the AXI system configuration object
    */
  rand svt_axi_system_configuration axi_sys_cfg[];

`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the AHB system configuration object
    */
  rand svt_ahb_system_configuration ahb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV  

`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  
  /**
    * @groupname amba_generic_sys_config
    * Handle to the APB system configuration object
    */
  rand svt_apb_system_configuration apb_sys_cfg[];
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV  

  /**
    * @groupname amba_generic_sys_config
    * System Monitor Configuration
    */
  rand svt_amba_system_monitor_configuration amba_sys_mon_cfg[];

  /**
   * @groupname amba_multi_chip_system_monitor_sys_config
   * - Indicates if AMBA Multi-chip system monitor must be enabled in the AMBA system env when there
   *   are multiple CHI sub-systems that must be monitored.
   * - Can only be set to 1 when the compile time macros SVT_AMBA_MULTI_CHIP_SYSTEM_MONITOR_ENABLE and 
   *   SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV are defined, and there are more than 1 CHI sub-systems to be monitored.
   * - If set to 1:
   *   - system_monitor_enable in each of the connected CHI sub-system configurations must be set to 0.
   *   - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations must be set to 1.
   *     - multi_chip_system_monitor_enable in each of the connected CHI sub-system configurations will be set to the same value as
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable in the svt_amba_system_configuration::create_sub_cfgs method. 
   *     - In case svt_amba_system_configuration::create_sub_cfgs is not called for the AMBA system configuration or if 
   *       svt_amba_system_configuration::multi_chip_system_monitor_enable is
   *       programmed only after calling create_sub_cfgs, user must explicitly program multi_chip_system_monitor_enable in each 
   *       of the connected CHI sub-system configurations to 1.
   *     .
   *   .
   * - Default value: 0
   * - Configuration type: Static
   * .
   */
  bit multi_chip_system_monitor_enable = 0;

  /** @cond PRIVATE */
  /** Internal queue where unique master_id are stored */
  bit[15:0] unique_master_id_queue[$];

  /** Internal queue where unique slave_id are stored */
  bit[15:0] unique_slave_id_queue[$];
  
  /** Internal queue to store unique id for each valid accessible master slave pair in a specific amba system */
  bit[31:0] master_slave_pair_id_queue[$];
  /** @endcond */

  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level coverage 
    * <b>type:</b> Dynamic
    */
  bit amba_system_coverage_enable = 0;

  /** @cond PRIVATE */
  /**
    * @groupname amba_coverage_protocol_checks
    * Enables AMBA system level cover group for master to slave access. Note
    * that you also need to enable AMBA System level coverage using
    * configuration member #amba_system_coverage_enable.
    * <b>type:</b> Dynamic
    */
  bit system_amba_master_to_slave_access_enable = 1;
  /** @endcond */

  /**
   * Enables complex address mapping capabilities.
   * 
   * When this feature is enabled then the get_dest_global_addr_from_master_addr()
   * method must be used to define the memory map for this AMBA system.
   * 
   * When this feature is disabled then the legacy methods must be used to define the 
   * memory map for this AMBA system.
   */
  bit enable_complex_memory_map = 0;

  /** @cond PRIVATE */  
  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the AXI system of the AXI slave ports
    * specified in axi_slave_port_id queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_axi_slave_ports = -1;

  /**
    * @groupname amba_axi_chi_sys_config
    * System id corresponding to the CHI system of the SN nodes 
    * specified in chi_sn_node_idx queue. Should not be set
    * directly. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int system_id_chi_sn_nodes = -1;


  /**
    * @groupname amba_axi_chi_sys_config
    * port_ids corresponding to slave ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_sn_node_idx. This array should not be directly set. It
    * should be set using API set_axi_slave_to_chi_sn_map
    */
  int axi_slave_port_id[] ;

  /**
    * @groupname amba_axi_chi_sys_config
    * node indices corresponding to SN nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in axi_slave_port_id. This array should not be directly
    * set. It should be set using API set_axi_slave_to_chi_sn_map
    */
  int chi_sn_node_idx[];

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the AXI system of the ACE-LITE ports
    * specified in ace_lite_master_port_id queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_ace_lite_master_ports = -1;

  /**
    * @groupname amba_generic_sys_config
    * System id corresponding to the CHI system of the RN-I nodes 
    * specified in chi_rn_i_node_idx queue. Should not be set
    * directly. It should be set using API set_ace_lite_to_rn_i_map
    */
  int system_id_rn_i_nodes = -1;


  /**
    * @groupname amba_generic_sys_config
    * port_ids corresponding to ACE-LITE ports in AXI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in chi_rn_i_node_idx. This array should not be directly set. It
    * should be set using API set_ace_lite_to_rn_i_map
    */
  int ace_lite_master_port_id[] ;

  /**
    * @groupname amba_generic_sys_config
    * node indices corresponding to RN-I nodes in CHI system. There is a
    * one-to-one correspondence between the elements in this queue and the
    * elements in ace_lite_master_port_id. This array should not be directly
    * set. It should be set using API set_ace_lite_to_rn_i_map
    */
  int chi_rn_i_node_idx[];
  /** @endcond */
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_amba_system_configuration);
   extern function new (vmm_log log = null);
`else
   extern function new (string name = "svt_amba_system_configuration");
`endif

  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_amba_system_configuration)
    `svt_field_int(display_summary_report, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(amba_system_coverage_enable, `SVT_NOCOPY|`SVT_BIN |`SVT_ALL_ON)
    `svt_field_int(num_amba_system_monitors, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_chi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_axi_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(num_ahb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_array_object(ahb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_AHB_IN_AMBA_SYS_ENV
    `svt_field_int(num_apb_systems, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV
    `svt_field_array_object(apb_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifndef SVT_AMBA_EXCLUDE_APB_IN_AMBA_SYS_ENV

`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
    `svt_field_array_object(chi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
`endif // `ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV

    `svt_field_array_object(axi_sys_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(amba_sys_mon_cfg, `SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int(enable_complex_memory_map, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_int(system_id_axi_slave_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_chi_sn_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(axi_slave_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_sn_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_int(system_id_ace_lite_master_ports, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int(system_id_rn_i_nodes, `SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_int(ace_lite_master_port_id, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_array_int(chi_rn_i_node_idx, `SVT_NOCOPY|`SVT_ALL_ON)
  `svt_data_member_end(svt_amba_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
`endif

 `ifndef SVT_VMM_TECHNOLOGY
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   */
  extern virtual function bit do_compare(`SVT_XVM(object) rhs, `SVT_XVM(comparer) comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );

   
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();

  /** @endcond */

  // ---------------------------------------------------------------------------
  /**
   * @groupname addr_map
   * Gets the global address associated with the supplied master address
   *
   * If complex memory maps are enabled through the use of #enable_complex_memory_map,
   * then this method must be implemented to translate a master address into a global
   * address.
   * 
   * This method is not utilized if complex memory maps are not enabled.
   *
   * @param system_idx The index of the system that is requesting this function.
   * @param master_idx The index of the master that is requesting this function.
   * @param master_addr The value of the local address at a master whose global address
   *   needs to be retrieved.
   * @param mem_mode Variable indicating security (secure or non-secure) and access type
   *   (read or write) of a potential access to the destination slave address.
   *   mem_mode[0]: A value of 0 indicates this is a secure access and a value of 1
   *     indicates a non-secure access
   *   mem_mode[1]: A value of 0 indicates a read access, while a value of 1 indicates a
   *     write access.
   * @param requester_name If called to determine the destination of a transaction from a
   *   master, this field indicates the name of the master component issuing the
   *   transaction.
   * @param ignore_unmapped_addr An input indicating that unmapped addresses should not
   *   be flagged as an error
   * @param is_register_addr_space If this address targets the register address space of
   *   a component, this field must be set
   * @param global_addr The global address corresponding to the local address at the
   *   given master
   * @output Returns 1 if there is a global address mapping for the given master's local
   *   address, else returns 0
   */
  extern virtual function bit get_dest_global_addr_from_master_addr(
    input  int system_idx,
    input  int master_idx,
    input  svt_mem_addr_t master_addr,
    input  bit[`SVT_AMBA_MEM_MODE_WIDTH-1:0] mem_mode = 0,
    input  string requester_name = "", 
    input  bit ignore_unmapped_addr = 0,
    output bit is_register_addr_space,
    output svt_mem_addr_t global_addr);

    /** 
    * @groupname addr_map
    * Virtual function that is used by the interconnect VIP and system monitor
    * to get a translated address. The default implementation of this function
    * is empty; no translation is performed unless the user implements this
    * function in a derived class. 
    *
    * System Monitor: The system monitor uses this function to get the
    * translated address while performing AMBA level system checks to a given
    * address. 
    *
    * Note that the system address map as defined in the individual
    * slave_addr_ranges of the axi and ahb system configurations based on the
    * actual physical address, that is, the address after translation, if any.  
    * @param addr The address to be translated.  
    * @return The translated address.
    */
  extern virtual function bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] translate_address(bit[`SVT_AMBA_MAX_ADDR_WIDTH-1:0] addr);

  /**
    * This method creates the sub configurations for CHI, AXI, AHB and APB
    * APB Systems are currently not supported through svt_amba_system_configuration
    * @param num_axi_systems The number of AXI Systems
    * @param num_ahb_systems The number of AHB Systems
    * @param num_apb_systems The number of APB Systems
    * @param num_apb_systems The number of CHI Systems
    */
  extern function void create_sub_cfgs(int num_axi_systems = 0, int num_ahb_systems = 0, int num_apb_systems = 0, int num_chi_systems = 0);

  // --------------------------------------------------------------------------- 
`ifndef SVT_EXCLUDE_VCAP
  /** 
   * This method indicates if any of the sub configurations uses traffic 
   * profiles for generation of transactions 
   */ 
  extern function bit uses_traffic_profile(); 
`endif
  
 `ifndef SVT_VMM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the APB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the APB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif

  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_id. 
   */
  extern protected function void populate_unique_master_id_queue(ref string master_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique slave_id. 
   */
  extern protected function void populate_unique_slave_id_queue(ref string slave_str[int]); 
  
  // ---------------------------------------------------------------------------
  /**
   * This method will go through entire amba system hierarchy and create a unique master_slave_pair_id for 
   * each association of all legally possible master and slave pair. 
   */
  extern function void populate_valid_master_slave_association(); 

  // ---------------------------------------------------------------------------
  /**
    * Gets the handle of the SVT configuration corresponding to the 
    * amba_system_port_id given. The function matches the amba_system_port_id
    * value given in the arguement to the value of amba_system_port_id of 
    * AXI/AHB/APB configurations and returns the corresponding handle
    * @param amba_system_port_id The amba_system_port_id of the AXI, AHB or APB configuration
    */
  extern function svt_configuration get_port_cfg_of_amba_system_port_id(int amba_system_port_id);

  // ---------------------------------------------------------------------------
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the CHI SN configuration within the given CHI system, corresponding to the 
    * given AXI slave within the given AXI system. This
    * information is used by the CHI system monitor that receives transactions
    * from an AXI slave. When transactions from an AXI slave are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding SN node to facilitate
    * performing related checks by the CHI system monitor. <br>
    * Typically, CHI transactions are converted to AXI transactions using an internal bridge
    * in the interconnect DUT to which the AXI slave port connects. When
    * CHI transactions are sent out from a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. 
    * 1) Configure SN nodes in the CHI VIP's configuration in passive
    * mode and hook up the output SN signals of the bridge in the
    * interconnect to these nodes. 
    * 2) Configure SN nodes in theCHI  VIP's configuration in passive mode and use 
    * this function to map an AXI slave port to the CHI SN node. 
    * .
    * The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts CHI transactions to AXI 
    * transactions. In such situations, the VIP will use AXI
    * transactions and provide it to system monitor. It is
    * important that the SN node indices provided in array are not connected
    * physically to any SN port because this function will disable sampling
    * of any signals on the SN  node indices provided. The configuration
    * information is only to facilitate association of AXI transactions to
    * CHI transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the SN node.
    * @param axi_system_id The system id corresponding to the system in which
    * the AXI slave ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the SN nodes which are being mapped reside
    * @param axi_slave_port_id An array that consists of the port_ids of the AXI slave ports being mapped
    * @param chi_sn_node_idx An array that consists of the node indices of the
    * SN nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_slave_port_id and chi_sn_node_idx. For
    * example, element 0 of axi_slave_port_id maps to element 0 in
    * chi_sn_node_idx.
   */
 extern virtual function void set_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[]);

  /**
    * @groupname amba_axi_chi_sys_config
    * Sets the RN_I configuration corresponding to a given ACE-Lite master. This
    * information is used by the CHI system monitor that receives transactions
    * from an ACE-Lite master. When transactions from an ACE-LITE master are
    * received, the information provided through this function is used to look
    * up the configuration of the corresponding RN-I node to faciliate
    * conversion of the AXI transaction to CHI transaction. Typically, ACE-Lite
    * transactions are converted to RN-I transactions using an internal bridge
    * in the interconnect DUT to which the ACE-Lite port connects. When
    * ACE-Lite transactions are sent to a CHI based interconnect, there are two
    * options to connect the CHI system monitor to these transactions. The
    * first is to configure RN-I nodes in the VIP's configuration in passive
    * mode and hook up the output RN-I signals of the bridge in the
    * interconnect to these nodes. The second option is to configure RN-I nodes
    * in the VIP's configuration in passive mode and use this function to map
    * an ACE-Lite port to the RN-I node. The latter option is to be used when
    * it is not possible or is difficult to tap the internal signals of the
    * bridge within the interconnect DUT that converts ACE-Lite transactions to
    * RN-I transactions. In such situations, the VIP will convert AXI
    * transactions to RN-I transactions and provide it to system monitor. It is
    * important that the RN-I node indices provided in array are not connected
    * physically to any RN-I port because this function will disable sampling
    * of any signals on the RN-I node indices provided. The configuration
    * information is only to facilitate conversion of ACE-Lite transactions to
    * RN-I transactions in the system monitor. Please note that for CHI, the
    * information to be provided is node_idx and not node_id.
    * node_idx is the array index of rn_cfg, corresponding to the RN_I node.
    * @param axi_system_id The system id corresponding to the system in which
    * the ACE-LITE ports which are being mapped reside
    * @param chi_system_id The system id corresponding to the syhstem in which
    * the RN-I nodes which are being mapped reside
    * @param ace_lite_master_port_id An array that consists of the port_ids of the ACE-LITE ports being mapped
    * @param chi_rn_i_node_idx An array that consists of the node indices of the
    * RN-I nodes being mapped. Mapping is done based on a 1-to-1 relationship
    * between the elements of axi_master_port_id and chi_rn_i_node_idx. For
    * example, element 0 of axi_master_port_id maps to element 0 in
    * chi_rn_i_node_idx.
    */
 extern virtual function void set_ace_lite_to_rn_i_map(int axi_system_id, int chi_system_id, int ace_lite_master_port_id[], int chi_rn_i_node_idx[]);
`endif

  /** @cond PRIVATE */
`ifdef  SVT_AMBA_INCLUDE_CHI_IN_AMBA_SYS_ENV
  /** 
   * @groupname amba_axi_chi_sys_config
   * Returns if the mapping of AXI slave to CHI SN is valid
   * @param axi_system_id System ID of axi system mapped
   * @param chi_system_id System ID of chi system mapped
   * @param axi_slave_port_id Array of axi slave port IDs mapped
   * @param chi_sn_node_idx Array of chi sn node indices mapped
   * @param report_errors Issue errors incase of incompatible programming
   * @param perform_sn_cfg_checks Perform checks on sn node configuration
   * 
   * */
  extern function bit is_valid_axi_slave_to_chi_sn_map(int axi_system_id, int chi_system_id, int axi_slave_port_id[], int chi_sn_node_idx[], bit report_errors, bit perform_sn_cfg_checks);
`endif
  /** @endcond */

`ifdef SVT_AMBA_AXI_TO_CHI_MAP_ENABLE
  /**
   * - This method maps the AXI/Acelite transaction port_id and ID combination to CHI transaction LPID
   *   - LPID[2:1] indicates the ACE-Lite interface port ID mod 3.
   *   - LPID[0] is generated based on the OR of the AxID of the request AND'd with the programmable mask defined in por_rn[id]_s[012]_port_control register.
   *   - LPID mask in  por_rn[id]_s[012]_port_control is by default set to 11'b 0 and therefore LPID[0] will be 0 unless the registers are programmed to take value otherwise.
   *   .
   * - If the user wants to modify the mapping based on their requirement they can override the method defination. 
   * .
   * @param axi_xact AXI/Acelite transaction to be mapped to CHI transaction
   * @param chi_xact Mapped CHI transaction 
   */
  extern virtual function void map_axi_acelite_port_id_to_chi_lpid(svt_axi_transaction axi_xact, svt_chi_rn_transaction chi_xact);

`endif

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_amba_system_configuration)
  `vmm_class_factory(svt_amba_system_configuration)
`endif   
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nZA3bk2eNHt7sBVLhcRwAdspR3R/vUqn6CoYkbC1OmDJzMj58y80mkMgg7dQGlpp
tNjTGKdQkxaIiD0/JADgOm4JZrbUv7jrHjkZ/N2cnHoPC53nc10TdZzGa4C+rBfT
SNFFZwHFl4hwFQOkYrV/wd3Nq/84uBmA0YajBJQQpH4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 26954     )
zoHuFjo2x1Sx30ePk5v6zbc5AtfmddmEJx0yMGsS7NNeL0Feaf/c4CrsReAFso4n
VdnAc7N59HOSpAfEB8cXZgGHg/FLjcQx2JUwInUrGrstqbi15/fKgq2GaDgNl/vM
v9qgAhmE3WISSToOgBqcq8EZklqiFKweVB2mTonCZI3onEDp/cwTYlG+g2L3jL5r
8Q7/xlBPg8idQH5VbR9F2/bh96i83JSG2wNA4As8Ur+Ojx1ePdw+y/heGFbRzpXm
QzcDdlNk28sjRr0TOiQ83lEmVmRcZfXc0//t6EVN1j7FyFfMou/7X6zbdKDERZPY
4KfXvzB0lImL+lP7iGH6MS2/jfUxBMvrOfUfL6R5R0hEQsJdija1hXeXWhsZTC9M
Xyddp6FqxYI8XKj5R4nUNUBhyY13+1Xr91q2+PibYaLAb5VDQH2kXsgSRtvcnntA
ZICtp7Edq+CG6grWjoQUQZUy8w98wY8S8QejrEWWJvCb6X8qxSNqhyvW5SPJ2eXP
dwV7R/iIpN362ip6IwW50NKgfrTEj/Dux+yCfUwNx5xnzlapPq38yeMBaIr8jf4t
VVgLpF7HSgaMP+WC0meFAkD5YrQpaggQ+JrWAAjxFRGimBrx5zia87iWXi4VCmI7
QlBba1//0HO9csFZtJg6j5U7PN/jelmfGgJDr8euhN24XAvFvRk9aZVprV+v3NAa
SMDpTq405nCi5uyGnNFXFCkNPKWWS8rVxILSvLCEiPIo5bNXTzMo0Dkfl66e+SlX
8khJGHnhICMSQ6XF1tZuoW4tuneJFj4ie+GD2Or/5Rzm7kWs/ePOaNArZmmpP0q6
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
NE6V0JkJFoRwE2W7B15dz/jqqyWAvV5fqoUso4xWLk//LozN/idqZcDSQY8ZLcJ2
pW6XKfTtEsk/IYeosUE+LLWT8goLhVqQnk8DqJ41BhbpCwQbk6TKd+QEEPa2HjPs
b8P4PjGnPkg1T8zmEHGYqAhohxxytBQ+8qfQ5tiwsOM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67119     )
TyHPw27ll2/PZZpdERVQ1fPTl+9nLl4GPSVV2ZrJEcdNgeYmjNPSPeO3RD2LdN5G
yIWUPkYivm6acMEkRYS5wUze7ZkOz6eD3B9huMRZu5SJvXtOu5migBm38U5rvmPM
KpPJ9U5Yy8mDknW3LVwF5HBxBrnh/Mb/Tb26NgJWZxcvdfkYN2RIHNd3mwKZEAD0
tGiJBLJIe9EfcAwVpBVyUhhXopgckYSbMdukW2Y2JWHmCMQV407DRXw80+lr4KOH
xaR51U/cfXtyNT+XEk0j3pSvzD1hrHKtD1/dDHkVGSGM9UB97nBK5cVspII0EBF+
EaxmRRoRPVLaXzAHyL3s1uKEbMlEhAJpUApj7AF5YY7sAvgVuW2Z1zsyHjO1MyMQ
B2BiI8kP+s0tmOmRWLWDLQiSmPLDfX2rvNj6MBCWzv8Z9/rQsI76y1rAKFRILv2S
3bOIQL1+pstR+xWYUyouVzIcERxzE4aRK5iRCTK72qZhcUispLORAgPv+mlfoENl
D4F2S1z5WdW1SsvyWKeODAvqqjggGuqKAxgb9f7WYtho0D1tpe3f2LGPyf+UnewI
nQCiyFhQ9aNJL62kl/H+djSerNmtH/WGTclBXIXGy0bTje/8o5XfKgaeKEj/Do3T
x/YKa6/UU9THokaqaYiDAs9pmbDGflBTP8ZCX4ovuJxfMSkyRMblMd6l3EJJnakT
q+CRwrrOU8HpPOXQVwux+TxZVowWDAfmRozk9EEzKnmkqrLza4AfORXwiV/6Jwhk
HkxfyxJNA7odfdp+25Wga4r8wajCp6seIsm1j/bErzZY4+gPuAW9Li17EL7qIM0o
E9CbWiniF927ysq6IMYVcMI25acD2dX8icA6+7o+q86k8UisBQwRrPWOc1jdT22v
DrT7J5FdSRtGari3bhwmcOWK1nTMRgHEL+YhJb05qg1N8Psbfe26Hw0Ks/WtUSLP
tynz9UH7DnCYJyVGwKZATjBQ0nP1/nssQIJl+lGJlxtX2r0JV8ScE9UpUTeNze9Z
j6PHJceyFXIvWmUr0g2rGgORGHIgYfaoFkB5i8ezaxQvPimb7nsrVNZLznEGuItN
RUczxtZ15tXbMgqiBHhNOYXlOFPAvpMTL1KLyfBN6orfE1j91C+MF4TSoWnxLpf0
Kd0TGGRm8kqlNyHcaxwO+UqDgtoWU4OddTGLyume7KrQZU0JbH7ue0jl77yDme7Y
CbOlPQam3vBg2i0z3Kz2kNTWBVI0GsI32GR6KIiN24/gYvKjNGS6z00IwE6TA/1a
AYt/zzZQngxZoRYI4rvsz9phH8xc1HDsE/C7w+C97ocAPzP9h+/dhb0doIwRU25u
nm+EVCm54SYEtfDJi10qFUwO1sq1CoLzy6iwrkpiEBAHI3njD7h1hVmCahUgM2oI
pvVnjG/RajHtTwFj1Fal3OTAC7lefP+irSBsW+qraNIMCJo/jw/gr3A1cPD4jseq
Co3WB5PkVfNJ91t4VK/SuwiOmBmIvoT0MFvnGwfSPmAsSXdHJHZlk4s7TuHyIb4g
0E9BMfzEcfNlSBG5+UzO4jju79HBrCxEPZofNy3vhSL7pSv41EXnhVXOYJbzCUIE
cYkpiluKXI9ozbHy8CewxxLemzDiR8Kf1XjPvQ8SxiLHmNcg+XvIURblXXk/KoSK
9EBbkNohAcBasAFAQBnMlCFh/uQWC8y1u2ngM9s0/kwi6hlFwnZ9Pmi0i9iR/KSx
dMQQz6+SAl2NF6YHwukmStiNbnuk2xQoi0jQVa/Cp/u4gm4DHsj2wC8xb+5gTIWx
obBc9f4mByoVGOaUdRamooY/0aSgDtx3J1GRZYMat5x5XFp4sporJuVlblh4JzMi
ekZIMIuThk8Cbqy/T7xxRlYuLrXybIAIh8fQAFzpX9u4bPE/AaLNtUsALCIsCszt
7uixmhw9vTc5ptFB0Ds97hbxG9BcZH5YhPdq30d0+j/dKEu6NMo+Ingts/Oj6Ymo
9NlEkeeS9RHoJ9bXbnwb8J9pQN9fTIBub0TKFP7jnXXChdbpV0B9NGUo2QtMBV5g
36R+qc8sKB1+fjBheZM4iXLrPkfLRlLN5JPH34jWBMgADetVz7d6RWNSJfUvui42
mBcMEUErU+7ZcZnpreALWAWuyrszZoopBmlVDvKr9X0y5oZX6PMhTPog3WmwqBMd
XbaSKM4kBWVAr8w+9mGx+NhY6SbNR6eSArorrgAJkhx1G0nSAuMLAaLlqO6WIpZo
jZXx8/rS91onc9cudKGOSIYm7ts36hg+ziHK70GtswyaANJQNJoP9sopMAvhSjsP
3fC+WE/fjJFH8hbHm2Tb8elxxteDnJmZpV4yqtO9RK8NPk2nmS+9vHF8ZmCsRS+K
PbABWArSs0BJtlBEzMSDbc/tD8jqenZK9c2Cn2FWzsPAhHr9E/L+j4niLRy+5MRn
6KbZm0GCx4OgBYSnpENuRd7wMP3w6R8Sys/DpVc4Yh1+79OoQ8XuKLsAhgOiLbsy
RWQEBVNGEGzqCS+iQVWbSy/49ndLjYCVJ4u5Wu8WEifUeAOHsWubW+vVXF80wTcZ
lhA1GL4HfT2Ii75LpCy2zpaki3acYJhI3mVwsmdkP750G3Wy+7Q8vo3ombenJ8RA
m3t6rsC3nUfXt0fjAYAH8JewoZfBmOWmfnV/ojEaTuSmYiUhUFhTAzMgufDd0Dj0
v9tm1DoPhrfdAW8U074rzL3oDDUCy9eUgVd5Z42nFgdizNzLQZ8feRu76DCaMKiM
Ux4TAoujsfuHfR4uiFoiOgmyPsU6PYx2mRIJrQgXBD4xwQ2HvEe+JkigNmdkbZGq
QeUzlVAex4otnx2uq0XyC5vbrjl/4l54cKjzcmInPlpBC/ystxe+ZN3mdi7eNcvc
zDIHbVUSfCIyR97hro0fDV0McD07fTi/5VMkC2rys82YQq+cjeEOqadDro4Tfdo0
Y2o0Wgarv/oTJmmK7wjdEzInFKMumGczGIFAyljW9fQbjnOocmHjgQSsmnuESYCL
XEGE50F+2SNxg7PbgsaQ7UA+uWKZQTbSY1j5Tee4ho3bmSgkd3T4FPv4q69Vwllp
MtQvC25j3IjreW50VLY0r8EFJbUIGEvdJDNDDMUWndA5hmxRdrj8mq8MwiuhDp+Y
Vh5khi5l+mRTQwfaDRnx8MLhaTDgveCdDqPUQvrRMT+qKSFszBJXdlLrPoB5MYaS
5TVWwXZwfOZWEHxnlubCwRmjYgHtllbW1vKCAf8wXG73/WGYOu2jU8boHGnI5NmV
hjsynV4cRoNcAI5iYKik5QEPhYIO7zJbNupozlSSrsMgeFEEE9OrL54quFyy0/yF
A32LJUpcLImCUcHUiNYW/yZJlvRbhbhf1SriV+dL0c/VvisPR11D5ThO6QdCKxJq
ylQ+LEnbpkAGWH74CnhzPXbLgXWJP3bs4CJa4Fn0BfUfDzbiO1yfdeBmC+5OVyi9
yl7z8md6hgEtkvoC0Zyl9Palt2jR9w9bFqm2lQADGRInIr3oD+XkZekeP6r4yJYC
o4yn9cAB8r4Kr0Gx1Qsrs7W6Do0tiUsk+7nOqMF+/PSRHQBbmvV2+YtQ8sirPBEw
kD+63UDfQpE8JRuIH0gnyz5n7vsz8xKOqfpzVOL2120SfmLMVAzYykqvx7xyBV4q
JKh7sMH5/ZUnwUEZIrRRzfnbq2vlQy10jCT3y6y69G3uMP/ekQI3iOd/GY4Nvc5z
YZpPh8inP6xV5D/lp5ySqzA3FKKUnKtXoY9fut3BJZY3QCpt188ZQnAxNZkitQXF
mxAkf+GhGUwe5J6xOIkL89rP83lF0zDJpWnRIaQSv54zh04Xa0/x5LoK5Z71xtlz
RrT1No4xGX1lUaHXmujlR8QX5+cYToH6Z3pTxGxOgE0TGcBn+N2IkXeeS3Wbc/gr
l13lZSETWiplI7o1YsDKFHgwImC0U20HBkmEZpRWiidKagg6PBD1SJbblEgIO/Hd
j38KA2H+GvqT9LPcfOSwlITw1DU0KyVSWrJwVem827LeAqyXLRUz9h9AorR2iGD4
20+zZVNTeIS+l9mfnaOtb1fNN6vs1kasbOPsJyMlD6Hg7kBEbwZgPNT5Io2Zorrr
/lCxeP3GgFuivrX5QUpAdu5PkGTTCw23o3H5rqLt4wQ57EQ9MIR0cM5ESr1LKV03
MdL+dXCD9UQT25/Hk2TC6A/U5hcWxaSySYq6unYZKsx4IV6P8rO9U3UNfgXm+1XR
qb1PcYJQLm1DLcDnyVflAir3imjXhmlgJi2iSX3kFCnnxRGKoth98znAP7XbQCQb
4GOByq3+fwK0a/7Xn1eVKrSja6yFwqmKsgQYDMi95Sh8jN7GdXGKZQXapBVXhMNG
7Dwtn4S2BXg1x1b2gmKyruHUNeILkFfNihFaVJV65zUfsQJqs9jAsQP33I1kmNji
e4FaCp1KBT3o4zzL/JxnlY/yRZQrTDQ0tHiSqopkUca+Dqpk+9Kg109U2oir5AOT
xUdF4KWg7x3gRJ4p/MrNS/YIWEQ4hbQMMGLEVfdIZ5PJKA/z6udCTugKFu4CGekr
6PjxhQUXpTUw0D6blKTz54PK5X21JfE1hXfwfWXPzWLK53kj+P8dtH+lEZr+C+ap
hayrtxEZqVghbI4RCk+v9/dgqV5FUs6X1/xBSSM8UcZadpVgFkbrd3sC6TfhHIrx
Xzw7qt1kRs6tH8NC7zXwTcQKTftixYI5wfsbBXz3rHHIGkSPN9MUfmuu9ncXgjcU
Z+shvZ1f6a8ZjSVKk4r9qfOQ6aLY7jFNX0SldDY0kWpG2Krem6T+xiCFHQw47SHR
kfn+Oxkj/K73FM66dEYtBIidwvvLrkrMVp9YqdVM5PbM6rKirU7HzN+AOBE9NhGi
aIHWiTtFKUj3uYZmmVlJbKQpDc0s17CjqVMRQj4+EXOtyZEVIKt71kBfpxzE85fG
QZTQjoIgz9Og+7ZGV/c5bGcj4KxlL76U7i/NijT9VBPUCgASGyGpCYkPv0SYjDSs
gdWq+Hls+jc4/P8TalD3d1zmVutoTwR8KyZgorF1bBNSvh8BimbswAzD9N//iF4b
8OTaIqVvi5fjTapewWj1W2k+pO06Gjr+LDmUpzdNgc5eb/AIR4O1I9SAfmLC/u0b
EiB3eR3ueV/ybiGa3Ti1PXcZTItyvtuuIuAPWa9Mgxfbclo0pLXKtccNRvmqkDS8
5RaUbvbZ+Wf6u6vbfiIEe7v5lEnJ0SEH7v81xtlFJ45z9k2wv9RDNWbaLhu3VTV1
vgxz+Nqt1bWpldnSBKa3gsj9k/bwRgxnHAIX1l3HEGdhX3Kvc15FmaB5PUxkr3D9
/nu/6dg3YxOx8g8YeMJiQ98SoMJtZSVMkFk0DVJh3f17v3203fTDRt8Z/rh1XkSJ
ev38lBTSGVFUQYEIOiTF1Ye7lglBMw5PEYIRpT5cSXsy8H5yFSxvq55tlMkwtEgo
+Hlmg09ukHkbockzW86SiwGPcgyHu/TIQ+F/H1CD0XO3fbPdUxzcdEor+IMSJMOR
dBxcOLi8NHpP0Kry+5M2wTXiBBFIJSL1s03fd5xeEiBBEqBhzJUL/UroaZ3aXIJb
qb9zn0bB60pm772e9koIiuuYQdJ5E0LAdqDWdoIuHLXZpocs0A3BV7cHUIUhB8/h
Soa0xiGT6g522Mrsz0abRhUBtQtNViZqCgf88pSZB8WG8DaAMJs8gct4RB5ZO6rl
58OSVEWFJIxpEEfuFJ1zaUMTAYtHbAezJg0Bq8GFfM0nyRExglHnQNli0Nd7K/D5
cR4Q9hmzJtRXnqy0xR4SFXwG6ZPe7bYEQbyDOppFxG8f7srMxzIpoN8nEQsGKFtG
7N2SiTJ2wXxFKhmvzptbt+KP2uaBDMPLsUeuiE/DfmW3iZ3qOxx1KTDYzKXRmedD
5xkLPwxwsXoMgElL7M3CsgHAvoji9Ssq94bFKRvXuBaA+lJVJLHnKOylWTYz3OEo
4U6NcEkR04zbia9d9ez0CMUzBiuz65sNpb4YEfanacEcLH3L+JN4n4KbaFORlcAk
r6o1C66ToP9Mz3tI6G04RTzXHD1p7q2eBVgzzvHCwMMc64MNPLfev64pdER/fKmw
orPSb8c//aP1o9B5aKczG4/9D+ZKBIHMJ6luMkuQntUiLUgG7DaKGDMvH4zgI+gQ
l1bI9uL3YNHrmKShu3QP0mr/hILgrCfM/n8zkLnQcqIOlyjnWJYiFM54nKQabgMZ
UGEzDqpf3rRvXvHRk57SaPPi4hVeC4z+OMKpjOoUU93yvPeof9GDAif9z0n59v59
6Ulf1nhTOCAnwx5gDPe+xEOe20/vePjZDaIscmL8b4ahd+jMAEKpP4e1CyQO63JC
7k0wlKwoUWwc4EhBWd+082dqY1P/K7R2ErO2PTgWdT+X9cMOzLVPO4P3RJFrq6Mq
vAfD/WLDCjDrdVZdjia4gA8kUzfQLL32WziGGgD5rY6uJ8EUXzjgtnXAlWuKEDcL
b+fCrUGQYos6PRCJZbPMRb2ibI0DJ+heEvHDngK0T9xqmNK6ZmmsXkuEiAfy9Bix
cnPV/+K+kYEI4k/FTKnsMEmM8ZVOBt96f5KQWXOviId/7JFTk0og9dAFiTsRjiqn
RLns0p7EWFz+tQnkV/w0+fJtek/kICQJsppOaza/L7JFLitRT2mwDnUiTakCEWGY
N9jiqBGI9j7zyE+Ri8CvlueWf+Qo8LEVkpTwrsHaOAsizHUaYq0fOlTA8QJJzK/C
x92/wRaQpom4sCk+/GM/1o0wnGPSETooVreitbvZHbd7OtGNTtkNKWXAJrplsumy
1F4jn72bMofw/X+dL4+P+aUmISDlAf9xaxrYCvDCjyGvkn35VDG/AdK2SmlcqU5F
vKvB17sVWF9EkhF0fbV+4EL8CqMe4uVvy7xiNV/J99age7jr90YZpHE81IPygxPv
YeTYYvO4p04o8wWZRCmHmjpGB7EYRp/s/iUGIglocWw6Zid7RFiHcrtEuYTulzWk
+HSVtD88RIXRf8RsQLfQUxopJNXEdcw+ecQ86irg4Oh0k2QY6Yv8vfzJsi+njrtY
X0eznQ6ZteY3uOslSAA2b7bFSgp7qd5rSKxPG9M3bnDBvNcmNvS3zva7gUF1/aJY
h/UkYfLF9gJSOPhBJ1xPlUiyIYePKw9bl4gVsQXa1d1UYQSSt39nuYpRvDIFgt+C
gQo/q8qsKHJKii5w3Z4z//WJL+czDh9Shb4pMLayr1zTAJK+TuJUdVqm/3g07whk
uv2f1mTk6NOGkMhR30QwEekVUZHSOT16whzkcBR6wnphjzBlvlDw1y0D0LZLE1uJ
Thk82s1Pj2eUW+0npAha73XWqGr3IsjhojCwR9O5r7KQYqXxXP0yTtY7c2Um+BV3
pp4QD+JC5rRIwIKZAqknNSCmt42gB0UPGxEFrFE2no7GyQcAdMIvpootKGC4DS13
B+JraD6zdgVgchyfTAOGpv82K06rKN+mbJwsS05c9f89kOz9gi0rhlkjZM13O8cT
Xp4F6mFy+m/8pkvKyyX5bZnIg+JeAxHSL8jec9QBqpOjdx7MAQA4gB7wOT9MNrzc
pb+br6Q+t0mcP71fp9JByQbgGDsgz4meSD7cZZyxwiOMUfKVLIT4h3MJsg1rJyxA
RpjjAUau2WwAjTxcxsIjgghsJdF4ZJV8r4oKUPn/I/SjocY8LrooZ1l6dF29U1mi
NU3c1lrVbR7knOQzTRwf8O1CTg6FB1d/bjGDEqW0KpZ1JO7/AQk3ghTx8BISe+8H
XKklqRV9wR/GQ/zBGH4ICvZCx0IimxCXLHDpL0mwErpYv+rIJ6LFMlk6JKKwmCGx
zrUFw7Ij5r7NFpVk4p2WZUYCqMNrh87R4VKhsWUzVtk6G437kfB6OCjvVZ5znVVt
+XZquKqiSYKwKeaAVwunD8/FlY76D+rRCICj+AIl8m/w1ryMlqDdIu+MXiakWpyJ
JsMFRKeFd8RYrqh7ZeBTWVEyLtKtxpYm9pUgIlhhuSpLJfjFoM0cYPDeZ9oMcrhG
EITo8lLSCIgA4cAU55eGSvHrGior8MoOk5wDEeTzbDB55hICEhO7pAHBFVvTuBXt
YDokLGY8ZiSj4S3sipS1506sC53U1kq9dgBwmhNra+wNYM6Oc3EQ5w+E2/udDo36
UeNB6bT7m9xtoTrvNeagbw4Lt/AiFUrqDKX8En/G1Mdx75eZHOpjItei9j56MFsc
pcNXd6eW+OddOCdJXHbJvlYxjyaWeVpwKUl1KqeuXzDOWzUO8/P8tm3sr5YYbDEp
dft410kwsaSWWoP0o+8q+p2q0Tve8GR/KspaEXZ4C8pvQwYSDxzuPuQMl4/9rUt1
GcEZoPSzoB6qQXa0W8QfXNDuekEfxI9Q9FNrNxmXNO2lSEwbKdOKCMB6eqMVLfg1
V48qGl6nOW5upJoJ6s3CjdVxqYMrNYoGEPlwaLi5G8wr7TQwMqh2AlMwasg2Nzrw
U8QW0ADwX2rLK7DYwCqVkIi3yo9z35tlSJ+NeNmDLK6UxDBRVAmzug5zWT5dhQ3W
C8vUGzPzl7ZThO/P2bQ2O7R4rIG9O8Ss63BRV6oXiCMzcZYbU6twm48yl5ppus4c
S33mBaMDaW/iwxsCTKVwDvhkzk1ST6kDJqX9B0iW8gSxg0DLjuBSLpKa7wSyymm7
du6fy6zVg1mU9Agq1NyhWfGuWkJL2AK0/vgWKULghnKDLl8zlxZGcL6hLPnoq2Fl
OyRDNEy6zEaNsb6p74/rx3LhdiZgGhZzGA3BpYLUielQ/LVPs+jobCcG8o439jH9
HmC49ex9r5UZNwrKcJOobSLbvSMaAdgkpnzX627H58AxLBjbQRIp3WloxuQYVu7j
C9RCKEhCdbr+zyW/Ff02HdSJ4vvI1kNL7hCUvHvvN8vp1veRSLYSdgJhnFHavwRn
8FRiuiqB0tCtgdt8yka+WMbY78kXdsuKHsktRhyLwhu6eY8bCogp682KdoBZaPbh
pahk4pe/9LUvcFqH25Wz3gcbMWBY3kmTxxfBESbxbeRaOmVHkTD3dbZwPpJAoylh
F71dDkXSQSmrqM+TPGV8mQYAmy4/RY0zuydndNWfehqEuqrmpcMYvUMdbcLdPisC
9gZsomW62MMGCb/Z6Pby3hEWP7/tiOL2EgN5qb9SqeSC3L/M1tlu7zybnT79wYuq
IAf+X04SHXI7m7qmLQxhwUkSEqBnkdITe69ILKY00z2zvxvdoBFBOxr61yWACqdW
7/oFytyIDBHQP+GNJin3IuuzZJxUnwOLaN4N/zPUNP1/NMpkAmDl9R9vPXJHUzJM
d8CmGWPe6o2DY/S0kjJ/okThozY+XIxLvlWz52WVsSOLvWFmpBs3836nmC8WPCie
lLMCLaltxW1O9qc4Z+7Lwd2oILPqbUj3wYA4mQH+ZSbz3gOYh3gM2wDq+802TkFC
NSc4cl4Q2wAs/t+6AoV77sDEaUzYTAV1QZjzPhV0qjpz61G95WTaqWuBtyi7t02I
rjTu8Og2HqGJ1N6lT5Kr+VH/PyPL81Hd6VFT1PRA1umhaJYMcc26ZGA4lLuNzDGh
Hi5/d99Y10m2gUYPjkug32x81t7j232WZwX0mas56lNGeMQKNMj3ZieIrVu1El/v
ptLe2KPGSR7dFhGNnYsmsGguP5exDbvFb9/jZGibJftI9szTm3d404WL6rnf3/Uz
CdivB7RSbGi+Lc4iiF/3P6N65pPmPExNiIRzVnYi7mA0GSZW2ZRPuKPPlBs8VqRE
Ktga1DnMh3HHs8ZkSTIU8KNoy9mFkfoLzwdCVuUzZYfskFbsq4KgcjLQ0+T6RU05
U62RjghhN+N+ckFhIvU0ooyI/d5l/IUJ3W2+oBQewaB6b4XFy8LAwuZBKli1K9qZ
tKth2W3sNkoeQm6cmQFEr/Mf43K1sIk9IEhZof0TeKje+03csF2DuUXxuBLSjbYJ
8IOmeNPRcSC489fvWxY1xmofTFUt6ztZTQWYlp4x9QpLhcFGBOfNn4+mgosZsdZF
j9r44YWGnIU53MXzoIgUVeKLVna+iW/J1AZEAnVSThUEZulYuJ1TD1q1VPlWhl9h
5/ysCGJ7VIxeOdzb+0GbaZMBubMSmLoLycV+W+OubWO9spDQmmAoqJuSqF6gKjjA
3TLkhjApF4G2ibvTwASPpG5jD7CygN9v1EzhstXbf8hlKlTuY0VDtn4/9opx2ykJ
rivEa/DfYWiwM5NB22pthWbt2BZEtBWNug9W25fBkfBI78RGwr53RaiyNzIy5Uz9
gEIzWkpuHc8LHq6pj3Ad6eLfiwhShj5RhJK65hm75/7IjgcMRVFMewF89MMLNWc1
Y81S+pEsYWT4RjO2F2ytwRpYJMcXc/tOQPUGqvsRQ2NmeUIwWG73KkrmkeDAJt8z
BkbeTrY02k1vl2Q0k3InOachfhxhWLucPOa6O3NoOeYJBnLyrqztnvhR63UHvcgf
SKpfa4CIsuXNsVNyYLuGQWUWt+djiC6585d9lxys/PgVJ518aoqlbS71zdfLFNcX
SeMdepDNcvFPrrCsmNWCVIGJKzss0FKtdzRk5LEK+aRnx1V4FLXecQSV+CeVhi8/
S1NprXE6l5uC/FezcC9b139GnNEaKJjw4nTORBT0yCx/ts4vCIopYkreH6i58KsQ
KU0uC1Q9lFwET/e1xFAywYAmCbpsaGXJVAHWgHFzvY0FTp9x1kTe5fgbh8Je599u
BL8KaMkWUfn7tjtWgkCw9Mx8QIpNr+tWrLZDfTjjhN1rhCEqeEqS/F5i02kYrfFS
TjqKdKHXeiCOyMLcOOWwFIryTJ5olXtKM73Ig4pgIOUxNSffWIETIvE+Tqbsyxn9
2I05QLKf3j4hxkm5sLgeRL2eSi1zLPWqLfw9lTeg31xYpZ0wttIcAhI3DLEhb/Hv
LHWj0JElDVgg63SeMU8kNr92j5gAmpWB4gkvPsDHlu6lSXVefQpLwLa4rm902gBN
2aRRuEjKwNSXVzOO5O/ibddztQIX3jObbSXrMJjJ8h9vE4alUgbqnHKrpCiQwTUy
6qMHOh96s+mLWek+XLpdJHcifXpAKg6KXazU5S+lUStjx6qn2S88/6JhOFlowO+p
sKqVMjjZn4kOwETmQXStloXy/y8QHhPczUeJY4K/U6kJGVB1NG5DlnWN9YW1+G2N
AG38eWUt2DdsG9mz6TN42je/uYnwHWbFeRZt9mr8aiHDUuMux1mvAXmoZVA2MHex
4A8ayopxpOeNn/l1TkW9NKtfEfhWeZy8c/E5gXLVRzsGAOJA93vZKdhxadRc+yCl
iKIOogE+jycNv60//yAkSKFWbLQYBKEvz87FolQ6172vAzsXiyLG0dPe4G0tzUHd
tB7fWjE1PLBU18I6fiEmS8/Zf/kGYtpOSIq+znVWssGCsHd61XYt0pBKE8uBKmZV
uDnqJQf6TPcdeyqc1QP9WT3pcGYGV31IYGSwDNJ0uOI8aWTWzGzv7ZWtSJBLHn07
QiJ63pl8JtKt6XaNWJbeTb5vVrn3sCHSkglM3pJN92G9Bn5iMnTDZGQ72R9Svjyd
Inwq/KCPDOt3G8H2tuF6tM+FvK5rpXAnIesSAI45hEIDnQCKjAjqI+MdRb/AW3ba
Kn7ccagWqfIS9UZFeF6IFsWTcKHd/kBQmyVZtJ9MkXMqHNWwl9DZKIxJdsXwjZKe
LExHf1NCoUowpEOkGPU5KZOKMjPmJQXkYXeIIey6XWJK2F3GMrk3RxxIPrm0tiEv
N6PPmzkcj9h4xu466pCNT0Emvd2CzCdHF87yXAY+eil28+Z1jfKTrsCOD30szg+/
GvA0YmlM+uHnrZYF1spj/q1sQV91CGCD/O5rhWNcn3QwQkqSyxKgH407N+FJyQZn
CV8lVRzWjFdxo5tXRiVYLtruS3tUXSmHFHCzp438NI+F9MP5OQ90tVUC3RkqkD0e
bI8Bsu0baJhEOZtsQcvxwvHbkx11BfkhlS8eMT1nAumXabKmDsCwxJxFlzAwkXhV
uZj2gUAnxcG8P7lT31+4ko0mFikg2UY0NajJ6+e6Dx2LJ3fMVxeCyuLE/F1v2DIR
lNWR6IUdhT2dL1E07FJYlzb98LRiB/UFmHECa+obDspnaX1EHxw9bgKnE8GVuoPo
sTrGykvylEm5YiOLEHPu4D1Lswvq4t+l/9DTTRMpc7sr0hO0iEzQvCkhSLfjh4cF
4yYqxuf7nuD7Ujm7qjI6qXrYA8jHo7UOZohrf0lhnJiQYjmFLgLld7DWWeZWPxiT
+9/WY1UW6FebiRV8Dq4iTFQc53jYyl+P51/3NJwBz6fJtveyA/ySugPKlT9vgdau
egDrTHYI8FHr71EVPNrO1Hf/P17jqlxgtA9nVptt8OIVhjQd2+rxC2mWr+d9Uy1u
eokOEgZnFw99hf2eHZTJkpkAg6MhzO29BxVRSHzuW11LQlUH2A0IFJk4pBRcljRK
iC5qmGQF8sY5qfjJcdQ53ydpSWVYJV6viKWQsU4OLQnqfRIp4txX2ApnlTcVM55/
Brb4A7K+3yzRWWjwMatGbbsz6yVLlqLm/R7QyZf4mGrh5T86oYsRs5T6ryd6qQyi
r9BUrCLB7o61d4vqqnNHUd9ycJa1UCZd4upv6GLdljHFuYUYvyx1b8L4Rep8W+kO
V3cetU2cSh3Dceqnc8jRrDiteBLFP4o49mRGlTSrlDSSLiv9XDMAEovcGk0ct3n5
h9q0gglRAiZoxSDBZQpnGfLsG8+tp6PBBRmQyk18BRO7Hfh+BnTAk11J+zQ0dZl9
6/wSIdPHSbhACQYmsjkpzdfOosvqJ05q5vhZHXBFW+mpdOFodwMTjSgbqWElNfF4
GHYi9oNzl/pGpx1DBVaDZ+gt/GyZO1fTvcRc7dkiVaNFgkz/htWjBD2D0oaSvAFG
1Vo0Zj3KYaWSjzSZYt/rq1YETyZIKohnn7xAncSiHMyfVuX/xKZk+tIlMvz+INso
G21Y3ic7qrYjD2i5IP1YCNgmNwz9vZ2pU+EdyWocIO4HvXYo1D1p7bz0GkPTMqlO
zV6LSOrJXGnlKnJAVNf6A/RJUEPL/YiEiLPUislT/cDfMJCPQfHCMa3hUZvpHQLy
y2nVpE5KjQhkwnzK13L2b4RjqfmVbawkeXUvqxNIIOOqVDVigFP4klgtVx6L7iQ5
N9FO/PM5NOFsXrIFPUp9eiSCYhhjkusNZKfEZzGmx4JcVPGtBPL11SmbCF///a4X
2a5MVu1wk0Mthx6RLVKr3Dy4M7JhkBbEwFsnxQR+uwL4hYJFTP5756P8h5GcR1Nf
q2HN9boGP1UpYQmCcK551lDr2AOtJn7JVewZkDsHWw0FXo4eRY66oz3yhHMgwLa7
Ki3IZdFrvFrUQqf0kwZaio5k0hAHOD7KPuSCvumhdShgPnzAYX4FXn1arcoytX6f
WKhfHX1ELH20nCNwfw/untWcR6/WtsjY5tkPQ4WqpLEV6YK16L0p4cI5HEVZ+pDW
aXrq3yo4lz1Hm8t9XH4gqCYcB3RZ47z6URu+6LUbF+V7885efjZJN4zD2rp9PfCv
bszCmCQYj/gTHR95bihGoFAiwugwEvbAwWX+vYyHHWD7Yr9jd1c3AIjWpG5S3zWz
kJLAS7hpANIMhVgUPG7dCJFxB4+ImZ9oNY/kFGPcP+lNbDkUG0zLOs9ndUS3P66x
bVO6cMw46kvQa2+B/DOq+KbFRzS0amlFSaQ/dlMwa/Ktqwyns5eUIqcy6lJLfHCM
S/LqWmiCbIBkkf94HMUdxcMyfvdAKVT5tL/K54xA459ymM1UB3amBY/RiWmcdr+D
Z72+5vvaeS8ldE3SbKkJ+l5D/FXuxhQEMwuVtaaH65ZZM/a8BndWCL2/XnRSQ/AL
5H6e9GusmCSB8WXsK0RCe42HlgnnMR/o/fpQf8dGOPmx/w7YSBvOPduhuogvmnrx
AYwfTEJ6Pk400ia6492ZXvjAmXvyKaedih5XwVDkcp4P24vfdDwLCFMqMzDHaXc4
PckEJzcOHG8E2Mokfp/f21wTId4RQSism35iF5b/9doYKwj1NH4JWNZrHc2XVYOD
SLksqtxKnnW4pTV8sx+fPwelCflfCm8An9tqRmB0wQP+UhADTcIE/RxOGngtdU3h
+k3FgZ4HzhpdlMoDrchvE3X30FcwfQfNvGzBGEWYM992ewo44H1OCXYCSOiODzUg
7lI+Izp/jHALBCVznVSKcTNSaJSTptSJw3jCK+mAYODhdz3TyysR6fBimPftiggP
wOoM7nkylxRrKY0XyGCgUyH8KhJ3842wre8XqH0eiywkVNAiAc0dfsoBlS/vNuKd
l7Cvrw3w9VrzlzqGqVsP8+MsHfl5LrmW9WN9WiPTkZ4cDGfV1sbMQzWqReA1Cy2D
XyyPxuOanZJdaFFH+/vhaN98RysJH7dgaRnlPhwm8ckai3f4zHYG9ryO5hYIWiF1
1EnVr/YP9e/rT+sxnEuO3r+7OIcN7yDm6njQLpGlvoqKJ0GdILfZWbdss+MTT+FW
C/1QVBUmnmx0EhfySA2ltDAL8aYa965oxrUUiw0+xboQAXbbmLDpNSQoKa44umro
bsLaLRGF7YHc3/vQpb7/NgHfgu96GzJ88DXLjunL2KH6qm+pVQgDgYdnvjInBNnv
XXtBYvclddMWbRr9P3dLcNTRYAw71awF0gfSoXZZxmBniznxYeqiSlvng/GAQBDD
bpX9qhvGhdx3ozBq9e1QfPO5u1i3a32y3ReNTfZN9Be4ntfUtwLgpKKFSn4jwDdd
tBnpJ/4zA+pasqSb1R8L7wiFKmPzhGodaHGnYFouWjARsD8CeHvtn3QlOq905kyo
AH+rDdShtZyagznqbI53nw16BrbfWpndG1I0aejq0N9efZIWg8Rb1/iNdBn1+Rkg
+kqAtELO5nq8CcPsFn5dYRMGjtaEXZvU4mijsp/jw8AKIU2OhkH3exE5/eiQoQBV
QpY5IONObWb4sLmD5yAgGZa5PkxJRnNVDBnORr0n8GdQxdMMSKRgGc9Cfn4UD/St
fhlGLX2CpRdN0Oe70Y/MDovFBRowmU1bEen9k2Sf1yUPLCit6Wqa7H/Wik5X03Jp
kbR11tbC4Abidf7d2E+Q0kH+nb9u8yI6cDp8SZ65G+QJ/1RMrAfw9fGGlL/Uj1Uf
FM50y2DmAmgr+C6LRDRroV/y2SZA5h/u6KAx1WcpqLHiN3fqdvjb1Jk8RG5JJNj1
gvgTrClcPIqMF5WidfmOXyjBYYCBMpzMeB9zDdbZ8bEhKCbJ68I3X0c02zRaGDxo
6ZeH+AFj6bIawSvJsjt9Yv1oSiVEfJV0UxUu9ZuHTLNdU/JvlykSbpqkTlgFTd+E
5A/ckNgP31tV68MyouSic/Yswu7Yxk4nIoyJwN6OACsjQJoNcHFCnWNEbnYAHcW+
DquQKXLDmqgL2LaaIfLMf74b+jGFfFkQL3hz57BcLFwIy+sBoFXCNic7ev2YW01w
RaEEDEC/whtj54OEgClKPC7UCds44H39ZelNPYDOMJE3WdxEfShUR6kXPVFjeBsV
5/dC9KtppqBInyPXPPZ34q0BeZIrI1tZavdrrK8mUMtdf1C0DgsTViAhgALSOHml
B7rTUDXNc8XlnqXuI+d8v97pQK3pCKr+2s2XCm8PchwLuoohhLOkUDcWKBzNZFRG
EC59AuVPShkdQBq+nH4ottnXDskwTburrTsuWzAIIZ2C7Xmrtg0jY9Kr9aWWJTtz
8G2NNz3soZhHsVIssd8D8mspXLIQ9EMQ4VDYLASp/Ky6v3mv8HKd4+Forg1qApKk
nEk3wABdok2WzJI9ymbJjl1+KRdMJE3VDR58aT99/sM4iQv3ZmUNEZ53Ocar3LcZ
ok6aui+l81dDB46arT/iyIJJ9ttaDgz+B/CygQi8dKe8mhIf3G9GR6fI7uJYZJr/
gCJ6fS1pvJKag+Lp6XBmwMMWmcJRnsi8/TzwNlZkefc7PRbfxwFfH9qOP9H6Spy2
7Ra4TuhNvXvzGDm2N/2NLo1umz19D72c7x8YxXoj8/tqgfVSy2PO9LHEAS1vk7qG
7bCZ4/pFDSTuOIOrZUGW4rYG+0PpyVmhF/3KbJw2Jduj4rSbKKYQj2yh2yHVOMOh
S+KUrvlqqk+B/B83Q867OR5ZhZkLZ5fBK/2OLbVDpS8zg9MwXKTV2XJBOLF7ut6Q
soSJDQTeSemU9YRJAzGz1/z9ytKb5Qpa/NAcDrlvTT0C37mPgUoxq9OntTHwMBIg
S3iS7aXoSkk0iAo183J428OuAzbNPs3viSGzs0muNKdibUsmep63z81890/cOpmf
GsWwEJc/PrShLRX8XS4iewwyq6/cLQTfR87wbrJJxU135mspmMVuxvbwr8BvfFWi
j9am5G62FvuhGo/CcGg9ubC5LshdkFmIl/nu0+krY1BIEG3LyOqdaX3PpiPUpbNy
cvbK7mrwMy7WrETWdGe8l3UD/631W5Zw7F1vuRURTCp+ztn2LQTO7avACI2CcrMf
ZffJxfzZLT6J3rjdq6C+eqDpgkp5VRxuUryHbty/z5eWAbLMjMtMWF6pVoJF5Upf
+yB/G73qBOGQyH8S9G3eAiJIGtJexWpx8zM85LZEM7BDshUYDo89ITarDZLHk4dW
PkeTLjS4D+dixVjWfQVqBwvvRbN3I4oA5nekQcag2U39j9ReMAGgNaUU35Zr0OBy
YCs+njQWfqjgqhaUisjSdmWEqg/s/EOcyPRoMmI/lEAJu4+nFrYrx7URqXffZDRD
frFY6quMpF46h6wVdM3ld9Nxsg2OArHOz6PMPoc5RYcmUpqafnwT5UCmMFfn4gO6
1J58k9ipVP0LbHN34tg6L3845XZDBXk1AMBKTaq12fYI0D9OzXtpfSstyEqMT7zB
wurBusXceYgAkO+a3ur9JlczbKEKQECoVzeKtjFEBqOjWvvBVDRt3SCJYoxyF/jT
z+Mswigc2ZCpjheq2pK8kWV7rZei2+tq42j0N3c0co6pWOgcx2b7rqIoK17N7UcN
7piE/kpKHj5PyEJ+/y7mWUPafjKh9S1O7s5X0Tl1sBxXYrzIkdXQFLrDdyVKJWEF
UBta/gwjiBzysjFWs7tAs/bT4veNSFwnjKh/cCzRun6ndftRj8brkAsNRTq+JzYg
QdKDrnthtAtQVK97kKrWv2USTavr1/UK2i8LvSJkTqzAkNfj2cpWnelCVdd00LOR
KWanZJI59ZKUzjrQnVBI0+nBPY8OcbppremWhWhMj4VSE2uiR2q/EcpVT388n8dL
viZu20yE2pFwhC/A8LEayM0yaYuHiBXGXBF2iuQigfaLEf7oDgsdtlOiNWGZGbcm
LvXJNRsCbNAyzVkXq0UdaGOTPcqHSngP45U1IziBbrhBUNJ/gjl+S3ydkKNyuzs0
TAM32DzeQ0/LvmL/Nqzx7BUOzwda6MxmU8/uL+TR29GNQliXuxGvBy0JHoppr82t
XLi24AY8KQYbo2olNAxSuk4a1TZMGL6WOY72cSUbm+OI1oL+CYQgD5XnxO1ylmgo
6dUxBG1Pftt7/gTFH00YMytPhKOMZI7zICmh4+f1IxT5yoNEHmGaWwVxwkDURvZM
ryRiOKAWGZ/LbFKyEv5nOtSXMy/lBDY9zUSsYKeDvC2vbPuB+LENA8PS5aO+gKd/
Dqv4okt3c3LqtLiLKvjSbezmIPSMfcZ9XuuIVhaqwo3CJuP5rzT6+5D9ItgGGGhF
OEIagzTNww7+sq48YhkfDnFQDv8ad8ZamBTZX+iEM8uZt8DgZYczdEzvuCTTIbVc
aIRKnrKL7dCR5WK3wOpYiaise43jgqJStUYZIwXM3EjkTOXfKAfmSr5ikQaWIQkv
PSQy4zdraC1bil1HD2Utc4/hYyqwqC3RR/5F8kYJvFEeGSL3ez9+tAlsxaKJno7+
LdTwEM8s07TbuANtzLXpfncrKhEQTCRotmvbx5POjp5/NwAfL0w0E0SY198XUl2/
1wHPs2A/F+VMVmTVru7zb2IHKa6McwKTdKlCQG+nty8N3HCCTH8iud76b4wwQJII
E+Eo/jvklYTb8K+lM0mjItUH0VMyj8QfxTyNLlLT+wbcb52VLhlSQORKZMeOTZlr
GLdOyG8zAjsThMX5v+rXzXw8ewjp5C4q4W4oB6HjgiNNtvS7maXGySzkfdrr5p2i
byjhcqvNKuvK2upRduwRIimL3X02PPpMzraNUVvHeXHxqWIxLYP2vcwqzrs3e+V8
w4aMe/YHW9vE5FpBuTy87xFqd7K39EIluU2y0A/gGDaDcpVwGFG8GBuc/5sZvssX
ZOck8j9nbdWA6nhlMev2O6rFvxgoLkgi9+FS9YcBEZWOzZUtem3bJbBdPVWHPXn9
krR/5Ub0WVid1E6c71VlHTyZGcsh6xU7jxlGnipPDcBDjWkN5VQ8m1fPhypX/glB
Q5fSpRPu3J+yuNZUzgdIHLXl0UBr6QrovA/hIFapGJDOoEcIoJxNc5o9AGDFOFaa
Nz3aCKqY+k6y3tMjApg4XYd5XwS1kAYh8kHJF4x/aNSWU0Q7Ubf1XzMAtEiSbe9P
MKsdIuiSCu794hbQABqB93D7zaqh+hqYw9TW9YZjDLml1tf+MNvgIDAafpsJv5Ja
CtsoAHy3jR+8jLOYQTOhSMVBh5aUkDfYTeh3v7iYn/QrXMJOPAs3OH46gW1paQdd
g5yUJYgvg5TbmC7pu45uvJhiOxRMu3yw8fdM3mRBIf/GNPQXGi042+sDT7a7fqW2
ir5Uuq4wod6BaSej8SgOT82oQ2VaVxMHtfEZRISGT1IODIbj2ATBcOqduacCbgg2
0RFAa5e1EWFuaGrfTQ6pMLGNnXngf5c9OF136z1/OvakNunLayjptAb7VAyjmdzx
/FWAWWHbYGtiJqOVoR/SDtgJeqORNyTn4bQRRKU2PBUqmoP3ZnO41qALNVHDtf8U
J/851t7eoNXZ1jzyw8Wp5po7OYAAoOGPPin2ndTBoBV4vYyMxDah+pVDfYCdiL2L
cGkp2wk0YgDKvsoC0yfFQLugW+GYa4Sja3yBI9tAU5qNUKcDtvXlJxhx+YlN5Z8V
WYzoauBt8yTDGA4AU5z0alvpRPKHs1EfPCgsSpvwDiBKGGD1kxs5f4wClJW+p03n
sEDkoh12mZK37lPQjhWds53WOBASmj4QwGw8IgtOpX53rOMFFCm7xuyRvATqDU15
EHCdX4XMRHD2/Uk3OcqGki00K8iNA3DcdnpbeDNjhDDO6J+Kt7+AnF6urHIDpMJa
uUMBtVSxGsShv0caoqXT75ASA530FAVO685msc3XKJv4Jv+SLIj3VJNJ+zjHhhwb
6XGCtI4BroIaxFDvoO+XmRjDVdJt7s1ipFp3BJfkfA3eqCGUNLnSFZeEgVV8W32q
dJ1kJjYfJbz8oJGp5KSg1qxeR5oEGEuJU1qoYwZ3+UJXiglrO2aVnMKQCr3zQbSG
CdKezUXeicOloYFyvzlhpkJbmiqCndKAQUWhev8JsUJEtCzWnosmdi+ThBla+aCY
5UeGqbJSHGDtPluQQbwyHbiNC6K20MP685rgRR/sj8DPOUvVHBy0oV7D8B3aLdRi
Bo69kxCnmZIuGPf5rY+OcfKRzzbgjM+G7v3cSiWWQU75G4Qo5F2QzWG194r+dyEI
bNR9H43fg1daZBYUbcCQNbjgTW5u83nuHswtafClP0aNTTohUABHVqmNknk6jbKM
ze4FgGjCclyu7gjGF3B06q1UQDHACj8KvoVkx5ammc2pUMB6TS54Cuh5rCxygjQ+
dprMj3eUTuXc1kKPZjxGD9JOAM6ONlJ34ox/WOMBqAWDkZ+EPBmAvbnbIL7Gz4tu
LrHDEspVpACLBHFEfedka+HQ3baIREOACE+f4QP90UkNOJ0FIjCPyNAKT59M6tbL
woBkJRLyTckV6hekBvIDvaWEb1+nmABtIh4jS6QPMMfoCQqyunayMsCx3quiycdG
myf1csVMFrUbxLgH1g3UL0LPqYraN9Dc+SF+hURW2zRd/ILRMUUeklkOEVEfC72i
aJQ5lYRDVl/+ImnLZVEZxOA6/HTuPVP8NPP/Gqe/mP1Irh8q3y3OKyNvpo8pvbCu
NCccTniAuHjb+Oma95OcqPaNe1gaYZxiKeFPuocMzxUAQqtFUmNNmlpSRO4YMMr4
cZvX2hMvFiTMe4QI6lRoLCldhxNk1az5u4UjcgZMqTB4+pYfpZV57lRUQXQw6MI8
o8BattChJHBmiMnfvUm9V0O6z+c2S2rA3nXVBQ6VCY692SJRejJZp5pm441dsfzX
V8CZEQhx9CMJ/JeYQAv10i7WkhSLLc4KEvfQWC4AF4RLeWCuGfnIKklyZAx/xCUQ
bQevQDboP1NgmXz2Pl5EWl+BOXdJw6rEozv0Jt+C68qD678bM++N9gPV0P3Nh3wl
QskDhuG2c02KweYFtgT5S8tgaLPGMb2Q0Nk3RzB/F0vwwPQSy8ESOHzTnJ0YnJz4
9cvRFoO/BT853ThieMO5hxGymgVW9+UyoM8DqF/jDYftyuoLN6k/pUMU6A+QluJV
FyorK37YQoOLXYRlpNH5f4BjUEVVEUypnIbX4sntWnthSaPnGIU7WqgHd/IogLIZ
7bUjOApa5oXtUVHqxVFEVADUyLfV7ID709t3yE7H/XXUnSuu9ocd0A3DTfy/qjWy
S6qPFoNpohSZuVTgRmScJUniVxKAJ43Zc29h1FZtNEDGwI2MG4n0LmxSrm1VmPs7
q7Z4Ze/ijMRngQYOO9i+VjSR/fEye5emEwV/4GUbGxUCg4afvzraW2FmE0nM/xpA
faVXT0vh+jNl+Oocm7DDBa5Pl8++FQVM7hSbE98XlAJ8kpjN3DZB3gc15/FbCSiW
cl6nK/d7GzNbG54EQriMxiZ2qYC/harsOMjuQ35d8SGhPTl5Qg3VK8wzkp+YoH/s
mMaI3WbRujRrWRabbUi2lqRepaiM3ZqmoSqZuTq9704XYMtxiUaYNdZN87PShhkx
s+kEuC6PPXFC62OJ+7c2IxhnmGbjejCa7K5y3yzT4DuCrTE5nS2d0BolVONxhr+A
5984w7my5xvJBMF9w1hUj3gUmnpqY43m30WW3cT2Ilu1XivHaB9F/kxCq8x/2mcI
F5YLZbxddk8lJuaHaSz4x+jeCqKfnaa2sZ2wrU8JkaEuBCk6x/+ukMr4vv/ZQ4rz
3P8Wz8iFDgfdVKOelyOQW5t9UGnNsAD/jOBGmJAgcO+SYjNZAHFsq4m11jBm91JD
byZgAeXaVqfgBekndS6JJPiKAdPGxRuVJAcBMPzpreZAT97YJ3X7D1gYVcMk00Q2
pxrHnrmo7A47FIpER++H8p6lCVZK7b5lpbCIoU0EhUgEoT3pBz7hctjb67Ctdw2o
VnaWurzsBTgIaegxMLHypm8P6ptxPgo2F6UT68UtO+kWrjMTRemu1t5NcKXMt5Bi
/bg+bvnoxN4K2vk1WZl86xXsrasrk/w76dTsy+GkYiP8CrrbUc4SHOp+knEm+Id3
eeUrdCNUHnthMwb4gskJtH4AilD2FFSrANRxMlhEfav2h0A/zSGhls/QUSAewwcO
CJjz8jZ7cusU8wVRHXLTZfCV2/s5nUtFrGwE8oB+OwUp2ZVByd3okk1YFogq26NY
zjiA8jzNWtFBCwQ5kO9MxF8WO+ySPljJJF/fXmNCIZ1ypiwlyeMwQqFZQpH093gK
NM0NYPmUTUqp9I0VedLgMJ230cGUJznXbJ5BHZfHZIJIDWN9Ug8TJ0hZfLw07sIj
PtLITXB7wHuuJWC7jh6SS/bbefa8Nty6z/wqSb7mLD614FVG2BMWq3OqqMxjeLc3
kQOCwZvFDoaLhXDxPdF9JzKrunaD8W5LOjx4z+Q4PR+BuPL1gYjjbYo3hPUlpUmE
uxGsIhHWFzvZpOopRh7qIgGiIikYRrAwaXyvMK3bOoAI7nygXvBLP9G95x9Xjy6G
0ih6ZRks51BxuuEQyumsAR/apKWbNPoOYcTh59KPvIQ3boH9if6ki80zIhRYD48N
JM3AxGZIroW0byfJy16JRZahpbodNamz4iTptBxgay52NKSqzTy+bIG0jYiJ9Krn
Y6tAIC3Cn5gTCnYrZmF6Zu0ylU0LRQAcQiXqAUPnauicUzhw6SWR+wtGE9PdONPb
MXm8NxWERAPbBwuDW7JHSSj2iCZeJRSHOgL42Jerqu+xNqh5D4eBZfu2Zxcp2uLI
Mbz7lM1EJlvR59PH8uN2wi+wuBsjIynqNvEWNK6VDvdd/6RcnnCqy2PZZrlSJdTM
F8nzZZncX/MuWskm+W5FTHzZ4BWq56ho8L/0bjzCYuENgLe5QkMTfgl216OpIO5z
CXHALuQIVK7dpi1WVOG6EfpsIHUD6Ks1ZfP/3YEocBWxtzRl3AlByQPWnu1xi5wo
T4s+pHne+LZ9p3N/kHLD6wWrg96nlf8+scHMMBBXbKJOsJ7IjVfXaTrHdgEEXm8z
zEHUt7EkHmF7So0D3V/7YFN/GrQvZ+vBeYsYid/GsmrWX2lfyW90nx9LNpeR/ooe
Mg/y3iDTzWZjwYO4KnZspx72tnH2RQVcIuoI3YLVvq91Q71geoTOqeIvkDatEM/M
lD1X8NtQO8l0bb+UQEpGL4Xh7L69OmIngKTwgaasD4htPPzXnU0JTv9U70j/l43/
eFJxrVIVQIetHV8ES7VVXWJ7ZQhCnus32NOIIlfhljXxfvelApo5mHJ11pdIb07B
Bb7fOplVOwoR0atixCP0XcIgCMW39JwRRJQx8M115y/6K4QNwx4MmjUxn4ChvKKx
T0lK5/1W2ZupLSdfJ3W5+ibiiIfWOk/6daarW75jgkqi79jBXJRopay/JdNieGPr
WgzrxUeI7E8K4Oky3k+QgcX3c/YH0LTJf9NfIGGnMxwu3BoqaZSlmjhNo6xscSbR
EKPR0wPY95ZiUhjxDWp81cL3PeTPRZafVlvVNlLQ85IMNV8U3n4fYINTRybUuI9x
/luwQ3Pbj2faDasckxMmgiUPm0hrZuKYUGaI2mTGoSbSma1equLHIhZh9O7+b7R1
49BMCfNRJOq6guT1LlUvTLod3UrVzD0jccTW3GfdxKW/3Aoc7iNH9OOzNvSDmace
rX7n8VbzhyDQu9yIkbPiEp7Rn8Cn58SnJdwm+/5/WF2ptsHJtxRFRW+x4bFLuxHr
0QyGmzYVL9AXr/jepHxHmfO3Txj7a2wYiaIye0ReUyL3rE6XmR95hhm9bjuem16O
gI53zMkZXlZ1K0OcM7gFLXUQ7MEOnQ6/N+0yMH0GvTxGnIUSaXU2nI5wsX1sEARx
Umtf51Q6eXEvaPDvAL8umsz/bQg+4Jp7DJJU5e4FPjSdIZ+ousvDT80ib91tXaCi
llP7BdXio6h3yPl/2FRegfsjTd+5NUIibNBU04xIUWxnWKQPe0mKncBYFIokkBHf
5S6DsF638Pi6DE6INHVEXWqCUwkI7mVhuEg4VFsATXlp/+HLyJaGoTN8n2sof5Px
DjreZQpCy034rZK/OxHAExQkmliCik0s5f0w2grs9KtL6dzTOVao9CeQ4fkh4wVr
3qi2x51q5f08YcjVJL8FkQD/yYh/1bpKLBmlTS5dIin9m6yr0kwi4xmsyivYSzZG
8llR+3kqhMfJpKwXTGI2WDthgkNQgg+KZgr7aK9GL5ex2mwZ3PSE/2RtPYv2csjb
kxYKf16Ib56kPiMJVzSofQueLYF0aBn5LpOdG/EoSrIK5wmBNylkrOBW60NXaULn
JFfe0SqaIQfjvgIvxKj/MgW1KNtdRCkx7Q1JUH6UUJwqLe/mHzPEz9vfdx45sYMl
pQizn5EUw4XXaJsr9F2cifygCjNDUYXlNR4AMc0F9t1WevWVzzazSRySplIqug8A
RuLln+QIjnhfancpTwoomBnQhanyl0Y0bXcCKdyu9VM5Kh4k0ej8CMJx2d1bcdXk
ASy2o277LwfijFnu587ETWvGEVWpcXEnCV9VA71/8zvbzMdzOvGABk/hD7K7Yw6a
q8tcbaDRp3cSeipTdFkWI2WEJD1XAfaNZ6mBQv2gyhYoHNM37gz4XATFpnPyfsTr
HfMqQotCxZ8MHvWMr3tZwciKzDjEKRhmGWNNEwy9W5YI9uJWbZyNkmWk4l7F6UMu
7px4rZyRqZE+Htm7GIJ7Zxn8MjY0y1CJmWaJh63fYVvq8HJlJ31WEvwY0KCA57xc
vULe9tNj/kGzzmQ/blW3YCkeayDN7XIDlJIZJZiOraIGSH8u16AVPPnXVq8Q1rM/
8Qv9dIFCx2nSdS8xAmPJ6ErJVV4pB0y1ej6/8u+5SWAHNz9CNR/6+2yAXZr9za6S
F7zNqJc4g39iAhkUdfjaNPCHsj+JjuU46jyrJkwTPHSkn5nS4fkz+YfCAVS0Hkkx
bCR1usvZD1mngdEIfuraT9XFWYpt1wr7gZBEon4Jqgb+ntIYhtjWm5zbBSXEVvGk
L8DWfQ4c5RX6Ulov3CEYj8WH7Y4aiUi5EoVHrXqW13lSlGX4Du87/agtjQ0hHwjr
8ayzoSlYgY3lw24q20XOpAPdjZ/NjESoJLmMrV6wubcYF+w4QE7lXxmngKNZxhll
940RyxhXBSVSx0sxO/AAAI7R0xqaXb6kDPuP/xyQiJIyhDWBLic5iENsMSP2uDvR
8n2t6/++x958uygb7KMsUURonCXqb8cKpSo3ntPOw0yK/f9OBmpdLgyOBakWmu4+
gQnpzXXltl9RAvojbUBs9dZ8t9jyhUV/6UMkZIvYYpcs5UEeQiUsnXm445s7Amz3
N9tC3WniyxPUUrSTDf/fjjqFmynwk+MxgbWDdAdW9V41goQqaauvbV1tkdO04iKp
akffGFtYF3vIGQcqut0SZxbRoVhgyMV7s/HJYFFef7G/STI8yKLS+4CXJZ93e8Jz
4jIQnI1gGCE7i5543cLOkeWR5XU06e4Nchsmxn/b7v6zhO+iR3ewQVJnoXqCEjfe
fOG/6z/y/W8NXUd+kJhadVjhmJiHem4aO2MvJBXASxJGAW5Qc5FY3R7ZxOsxXxfN
ivzY4Rlxzr7IyJdIXB0W4b3wI+RcICqEcZvZMV8b6Z2PWzH4+jr1g6envUxYN2fY
m1cieDY7bASmrfS7a0IjKscSJZ8TIcUU0zF+5x9blGL5vIFTA08rd2+C4bzfx1l4
bf+KVtIlH6ALRL5w4Z3S/txsglMgE7sXSZ/tOZDAa4QG4pn6ZZZDLIjqDX4dSV5t
PQzVn1EDC82THX9HytN16czPe7DLfdeZsGzKaVbTZb5qI8i4Rcs31xhbIIj9BQ3T
Q/daoK2IlJtnc7ne9yUlKpatF+s2zn/zysvu2ND0FdVhNgTBonORrknqYBcuekQT
vPUa5yMbtQvTOwH9O7oMGoMhh3YJqXvE5p3dr7oYkxYlQfaHL5xbFAgMGOhjkf/H
k7lJWxuCzspkMG6p0NNzOhrxueJnFEXCTIhcs3RMRAAlZAkIYAZtWlK7FoT8O2x4
/1vTmsrSL7mnX0EA4sZLSS6ElyvzBAdbV+nZEZMI5zWwCCa9vQiEyLvhWp6IkbT6
/Qy6TQamxqwKNjMi+mqwDqeuj27Nl8X5DlFsischMyrQGN7NQcpnhx8m17nR+bNh
mmfTIRFaOe3jcGo/8bhVECRooj0zJToqQAJE4N1uiV/T/ZMZteUyZLWfgiLYdhAa
Y9ysj4dLGsSwyBvrVr57IdcSvWBbP3cgTXa+l+vKTfwMg2Yab4X+7tOMYPi3cSxD
+K0GJQPBTopZWF95hTc/1O0d/M8omznC5TZei3JV2Tg4k4bMwkaX3UptE7wdr2Uu
H5qAmaKHpQ1/75RSyunHfwoZr8h2YLzUv/pGpIbIPegTu7ADYFeyY2XPrfs2FppZ
RRHBotpE/gNq/Da3CeGUHkTKbs48OHGZVj/J6GrW0+VrPgtI6TzTY4TP+BYHVgNE
KMzYhALd7iQ2lKpcP0ycY5YnANGQ2ypB7yu55n/kf5HPzf5m4NU8EdQxJvbAOMse
pW31fO/ZU2EW9wSK1H8OMS5Ck4gSytYm3CJbz/48gJQ2i9MiXNl14G7e3SYR5/vS
A2oteIhmA9Kp8yS5skbQE5UyUBtKR4ZWTh2IvIiSYEsUABnuAPOxsI8SSU04LCI8
aiwvlgV1ZyvDDgQxdjaykHJlajowEobixwRoXMOZVj+wiBX81LLVrCkISCMtem/A
M8PrETW7TeZBcGJwgVur185jAEPiQKe6dSAjMUzQRwMbAKH6NKj0gOui0k8xd4kI
1wlCcjqYOYr0zn6GaTytvQrA6wDHDe+DQQvRo3DrxHbz+/OGiOV5OzSOgwOlDOe2
fsdBBDiFAbozikKrVvXYzE/o0HWNjNg+EvfGy1v2M74VNNQWldQz2CxKrSHNgJXy
eBSjj5DYgVV1EN+31+VDl+5LhGwPDSpwlDmGQmKPSBxQVIjXaTRg2l/v1pjnqDrt
bv4TuEHLjhCuL5m9VV0U6Cbu08MAYcVOt1nMbxHgQ4X0WxsXTWRvxAC/XgzFVJFR
2tGWUMdbFwiTNck6ITbymyNNRVc+YyTCExJbHwbknSqcZEoKE6riBvTB2bVB8DGb
w3/4uLqUIukPYJUcw6idJT3G0RKbohWF+4MYzoTvIvpTVUCXB0q0Uvs5JSuIkowH
k6G7SVJ5qLtvSZyP53HWBrv7kbFYrUD04/d2voq2S1vee47jo1MnnAj/RUXEhetW
k9qNugnq+0HJylc/XXnmUvf0Uxu2z8J00erOWtTu1kjvb3aXNZAe8S89/vHlqHb2
bMANuY2+NymfQ6i72RYYFWx54y9sre4GXbjDnExKUAikSP75pqnudzTUwNWkpEpW
kLB3a7DQUoExNbJKEScpFWaAsJqEG7yeU37vxB91oxvvwI+Nn1Bf8wHWzG/PGiJR
BH5aJvvJ1Np3DiXvJMosL0Z1Kd1HW+zGvSzjGI6hXLEk1/AAWCzcRZqXS4LxAkXa
737wmp8JpqW6sqx0neZ9dVaScC056w5beY6WbPQ6d7N1rYA8wIRQVtflwKcDNzhX
GCDrxlCfzY01mW+pCb5iJJCXugMLblInIxJ/ZOS3SNaVy0Z0PwjSX55SuWU6XPe2
o1O2JXinwZekUtiWNp6ZQXtV/rXkW6YcO/xp+sbvJhjDEyR3jBfv621YG0WysdAm
xm7KZERMUF0FRdq9kvZjiXBD8dnH61P+jjr7iLFhuOoYq4/D7fxdukbi2Jn+YMka
1WnqP8dXmbWh/gWH183O3Hm6GQ0nsNAwcV28wxpkTNOyFZBTzunmHGB6BN+/fa2U
mWOviVwxz3PP1oIDQKRLNpZ78K5r5xaYgOBxQxxkvCGOjYnD4P+Nc6Avnys6IxCE
KZyRHMsFQbuIhbg9YVflrpvU401AWEvsCuMHqMzl2X/ps2mJuQnL3kbrs1pH5jsg
nz2kYC5gEp7nKpPuZnF2IkUY7Kgm2C2i7j3LfUkCfoG3YpCg0lsCm170dFJAbWeV
ZNpmeLHWHKwUtFPVQ4lq2S9csqA1IngwEWpSAcSglRiS/L81BfUYVqd5fQ6Y69mj
NLZCplRPlEMIbMZfbkRe4cIMG64giGLqhnH1lNUuCA2lO3uuWG0z79FUK+kf7iGq
6pDPlVoafbaid9Fy9poHA8aYcNrBi+Jczjv1KPh126OYHjEfmLglGh/DKTx1aacr
Jk/wSucDkskcRSWxMC+z7VvT2V9Yn8Ndoys/JaTTfJgNOCrDayBofXlVRjvcYuir
15T+Ez+uP0tfeTFkKv963Xq9XoPDVOhKaIIdcuXehUDpSx3IDml2muU4laO3j/Lr
RZb/gyRPwFaDPOadN5NmQFlnhYjHdDY2cqpEVusXxUINwLNh3pzfHdSCm8WV91Cp
Cazv3oUM9QJs3T6x3WpAfjQ4FWXjSUqeA2rTEKRyEs5+siAGwjh4EQHVyaSQ70sE
B7sG8Re0ppifCoN7gpE+Wz0WYo62szHj24hVfocrlaYTQYYH3oCkRE+9Sj9wHvMC
ANQ6OowcfvItPOz10EFO9S2u3oPx6r5ck5FTMRpFkcYPSXoLtnjUHICgQRoow4On
OLAAW7T5FsY6ms+ZGIrf62NFvpMrn+V7JQjG46Tc/bCca2X0iRFWKCDzHzRlqHXw
ZCr3eRoxwiLi/xMZbaz5fdrhd4dbs0oJAW01lEXJY97mYIgjaOmkHI6Wg6VTBhYJ
JYZ5MbU/UI8OB1UnqNBXi/ouZqCF7PwNUz0cE7YlWoB3v3ioJZsNzvrBb9UvTgRe
pbYR+g8BKnLcLqlZ+KGb265Tp4bwUmDwnNrd4K6lzAwU3wTcmtSj1LhXJFGelQCe
QBDU4m+rDjRrLV+5TfSMUjeNbOsGSagRJCh5YNvo9nS0LtBzW3+CEM4rUF/9glJ0
zQiVlmnOjhaAq42ht80FeO2exdwuKsIZ2J7ouvnYBwKKRWJmn1kVQdXuWV0+CUbJ
+Z0pDKWytpRNx1OcwdQPwEg2jKlZhY5BvBjhM8SLfDJPv7kPGb1Lx7OhhnyvwIG1
ZpdbskiPBAV6mE1d/tdc74Y7ghpJSBvXtILCBQ3OZOLqMILtpRCXZm5OfWNMPVFX
Dqrmks63VRmCT9AIFvZK2B0c+6UD2AQMl2zmDmW6giGJxuX/coLfANu/iNvO74wH
xATca9H7sYbXjqXjCxDjnP33N4BK6IHt5YZO0vYaChQyFjdcp2FiGAq896NJa9pP
LeWYR8IcsHyyMZnxegRNp4E+U+FtgrEjn61Uusi3qQGHBz7WdruILG/oMBtmBrBC
YsIXV859cs91TWh45m0ug4BKSXBdMX6HQqbx8BPlYAFHTs9oFbxsSk8kXB8zXUk4
QJW1lqQVuwC7hj80vs8czYYQjsM7ho8ipa8lOgI68JZ8ykLWkn+vdBqBNtb14fch
YmLarU/M4FFGQ2lK0537+IOxmpgNVPigi+XxxVOPqD5OrQ1A4U29/dL7gqpzSSkl
I+vMQJMLrcEQ0LR6Wpk04MKzwHfKVPZEbhKIjsG+Y19vQRpMrn8RVcMIr52F9gJG
Pi7mKA2/L/8zMLGiuoUyjvDihRdQ37AnB+TAXy45HrFSnjTNGo6FuWS4pFI28TIn
RqKEOoiWcXu2t3x0SXLNKjXy1NYqeQrti+My0MdhUh7llwjNJZQgDFGd9m6iwNsY
QOQGwPY/Mtx39H2NSnqqA0rnse1hl8N39+IwyD32x6UZ8QSD/qLdMKQ1C0Z1/Mke
oKP2CWrJ8qnwh2pK3rbtJ2RMIXe9FyefDIcuzC2HXnv5xcInmvlhgQcA757pyiGb
V/6ntrGw81GZmfUY5+92gCEer/lWfN6j61bLq3dagGt72UQjAvtROTEI8hXGkgJG
emXIhp1S78lHxFdpSeQz5E+nOi7oFlRLj7gTRlT15AjBashQwtbt1uYKFmX7ewRb
/P7CTqQ5+kEpmWh6jn7e3S2YbevxrEmeoKsTrpB/Dmw/WenEp+qEfnUq/jaTk44m
QXMkWUTZR4oKl52TX+xTZWr8P3p+o/e6WMATNGKjVBrr0BY6RLKlwUP1tQu3hGXd
v9U+oaRs2zViKVsWoEu33uOWkd3s6bfyrJBToQUeoxgKbf2ZLCmD4btUS6dKwYfO
ermCXK4iDVFEVDahKdYC3OCcmimbMe6734P6RhkR6hQxaC2Vv9kcS/6+U3v8C3hP
WyfuVW17KwUtYvyv/UKr5vYrI39ytUT6fe1Y8Qk4wzOWL9CEcRnvH0/Y7TIm6T4v
QJSzmGZLGiu1m8Nn1BfIbcpylC3tBbz8oqQNKHbK4pKxEjkXMB35gn3IdTCX0imR
DsWk/PnJ4qYejIhkUsnKcIhd4pGhKU1V+nZoZ6hgjzyuU2obPOutJPwwd3+4pA2w
EREMPycEhE33ZoIg9o8qMsmRPcehrEzZ0Qqr7qtgzY9twknNOnK/+HfHRwoH/j8C
PoXM3xxrWOkyg+MvcRR6lkbdyxtLEbZz6BKw/Kqq8MhVbUOyibjtkpMcpraKT9Qh
eGW/5vYYwzKETM0CnILY1IOFMoPq/YXq+IoRryIEZQrmSm2ztExcCwIYYyznb726
EHu85q+0PH8Y9Q6GPHye54PRZxnHh04mtQeGsazppfuYAmXjOQ5osEFQZEluEiip
c3B8wly/OOiNuVqIyMwgfW+nc1ox48nqSGt5dsrfMVsKEoscLDstasABwwgd+/UR
ij9e5pAGdIz0YruMvL4UQyqPZDQFhtMYVYcqf8i/hIZH0bMlmhNYQtwkmH04vXPE
FB3cmvu9cB5VxUEftOsv4HqRbyveOnFLj5FbFW/ecBF4rxNS6b2d8b9mIMXNHYIm
I8MEJRmK6T9sNE5mteFtRMv1RJtzNz/H1Wj2Bm0B9PTh/1jqMEr2CfnR9rW/J7jN
hFTp7ghANvqpWg5wOZKJILJhctyBv7QxHb1dWP1pc5qzagCDkVVrojPT/PqW9LLV
3kWhVCec5VO/eew/abXxHymMSlSkH0mvXb2XKiE+pdi7wJI0NobAuphcwHJkMGKJ
8XYzXwrbzF2FI4ym/e3/XYeV50E10S1D55Ap7JLIOnzC/JgpQWL1UP3LkMvskeKO
+XvHoYBgHvBRAfIGznrbjBv7S5LJX8PxApRmloRq4xw+eBl+aFwzFJchGp7fxjIu
sbj4fzKa7HEjcfIEElk8q+LR/pZdERiY2sLpUx1uZSdBXulIvGe2qRutS0dMOfVG
6SvBtBYdLO9L1FMxlkl0RLTajFmVXI8KbNskZNgWK3qJ0ZVoavc7qlk3XFwmSFup
iXnQr0p63IWM3ggafQh0fCY85V3367Kl+26UmZ8tfChBtq3hRqAkW6LKGNxPe11R
ClNfX2F4Mf59pOV6KWIqgm9IHqn43IviSh/eX001/Qy5k0hWxCAf4VX8AvwMQMnM
Tg7nLyIsq3KblLzUtc1TjiFnnOaaPn+8j6xiAbmfr/2rRuWT+WiyMXmhbN9FTS8Q
Bl92aaUWTFkEiYQ6ceU8PnDXFDg7DLTDTa8+JUq1AhnHqNWkP8Bcvh9ppZygJaCt
wIploLGQpFc2EjdBCuL6WRJGuW54DwfHIrZACH8D6Uz1lqRXb2VHy+3TbXbDn5at
WKjkLfTt6HUcYbIpHHXt3yCZsfpRH9qzbUYlotqdgnfcpvPPPBco79zCfjWummZ0
NwHthtUGLqOyW8F6cU6MA/czg+w7QkyaO2qvnPjuRQ2A1rK5cUqFbPadZNVgThh0
rCZTyFEGAm97GAAEMhO1B1hiBOjEXxWuEvryLo6qF1loP2cbxf7QJ4yJxrWvxDxr
A922KDMAMHEdv0NdjABpH80yvdBgLX+DDbl5m9yeaJtcvJZ0ja8Btepiok7bKgpl
tgLR+HeIl/lAC3x7f6njMJhoCfLO0Je1YC9Rn3TRBeqw8xnBN1KvpL5UU8m08XRA
Aiw8v3B3POol06Fc/SWlYmSJ9PZmDe1a1p8lKR0aS8dBRQGZfd5TzklDikSJLG9/
LnV8VS9w2LJjRlX1lrH+e7jupxirnyZop8SfVvrT1H7me4QbVDtE3XCYY5Be5R5W
m+vUH+cQ5jLaMGA7UEzQdYL44wYa018kCwgCAeDjWJ2/+CEQcoP+T6g2vpVouEkT
QOzif7bwPkqILbIeVMSYFent7m0ED3qcGbTBybgDlZkrYzd/cIVjGCmPH7EDNEHp
RJCdegR3PGAkMw8b+rjw3lIMF0GnSWOkRRlGLQMBjjGo2iyit2Y5z/WNEQoFIqOe
9qY/sHqEPt1Kw2fPal4kN/t4Nkcr+FgqHdw8khCR3mt8VYTO57aGA0RDOX3xJtuT
kZxKJ1Xnc6meXwPUKBZ/LPIypP21dW3krNMkbEQ8ajFvoq6GZvxJ7z0FnkPocMDa
midxMXcBU+uMT9EjLNtPqwSTQvjs2mCQWTkAkRIV6ql+KsYpW6jQZ5JZA4oVdEvZ
KKwQo5yudPCKK5eE14/0+g6Y6KyeIqbxYP/fpEBu0wH7nrAGVmUXG+Q2mhYI4jkq
k4vu48aLdeAXzZvfWKn0+pCO7z7sFoaukbvKGuGpPAZcEeAv8a5M5C62AQpT1exq
9kS6maptSXQo7qcTstwqlVb3ZK4XOlbDBy7C2G6AnYKOhF0r/4ZsvlWNTsEvkeND
CgF3ZWtfw8H0PSi19NPI15LyR8dbOmX7MJ98wEdt2/KtkbmA3X9UKcM75VBBjc7b
8ui2EVsDtDkgwSe3Mgu43vj+mg8/eb8N1wlZf5RJ4uqzH2pRFrYXtybrOvTko+JV
GzRUqLiW6tgI86iKWWX+QrzNIwseRwsfoNRwEtwjbCpwoNPji4pYpykrFdtyIhud
Ta4XfTQnA05zB1bGmvKnccZaqqaiUHhzvt87FH3K9NRBV+v6EI/dtNzQrdiI4Gz4
PmVT9+EvvUb+lJLTJ5CWUWyJOzQKvcD0hSrQtCpeVb91bCPIR/XLqbW7Z9n9JOPo
GrnQkZIDOEMOVE6DOJUAIxqeCAlTZNzcvBV+G3nEB+kRVYFfMz8/9P09qEmRjAUO
OkQDFovzXsYVUMf0/+JlSshhxzncon09m4fBYQXHrCJe0uhnsESakhsZ/OH1uwCd
u72EJQ1iroWmCR4CVei0+LW/URuydVPfvBw6RtFEY4VLiu3WsZKYLp8dO95yciII
E5oZriCbkGHa2m1/51+NXe/IvKxB0kxb632eEvJgl9wymFFKshkfTzziHuRIeJhm
oW0IPGxY/o7V2NN/WqclYsXxM87UZTWW6bO0qANjnVMqqk45Dk11dwzfDb6itMnF
gw86B8gRliNCM4ZqN5OA0HJcM9NZkS3YUkaiXC63VBgltFoCbv81C2j/rTmfptG+
v3ILS3rB53NzEIPhv2+L3GEOaszj++QL+pVrHS20M3Xk7iuSCvhHLnB/DJcY+Vy0
9CRjuFEjXsG/nliyr0xRVi5F1g6LaFVlVKutdIgXZ3X8wFpEFPm1oErHzSet0P2x
/dhS/D5v7HB2Y6DMpSnQfngrO767m+29MFYcbbxppsjgrO1d6TXqrKr5ZKELBbC4
moCSQkU4oA+Onch0J4u4BwaDatMvlveFmJdgt1m/I2KCLrrTfVPCTQ2qpptffPil
KSv2J/VrqLG2LDhuNFWPfSL9cwkItXi4gk4nseV33wuHgg1F7XWeadApUfG92J4W
mEXbXBAQtXIvEZW+3usfw+bLgw4EBn1uKnZTrqjr5eakShndrg2SfaqoUC/HbHQO
GJn7oXzkF2Ux967DefMX2mCx8lVwph8AH0IUBxOeKIN8Y/jeXTAv71j1ACrgJQuU
N96f+lzIDlE3a90xWkQVZ/3Vmpt8mmpo42Yh62DV35ClWZ4ekRot8rOoGXx1GNTl
Nr/vli8oLMnGnFvHcKc0azSFxf6og5ZRRkxbMaB7XxKTIUGo7EL1lLC75yvvGeQT
Y3coWqHWDadj+zDjY6GSe/F3q8jEK36qaYM5U6AFd0sbuh8vbG36uHmRa/0r9XDp
EEkm3HGklhM3d+L6+l/8IWU06zK3XAPJz9k3VRXBb0sF6ixHnHtGtjAiYmhhTd0g
7dc/gicBCMCxPCrajrUxp4MGT1yAkMrHA+2J0BTuPEFwaYTGpb3CwghazhYOOkPi
Ya3L/PX1gcpgIi27NZkIHtro7ZQ1WEgW6/SrTeujBqv6x2YRlUXyB3rRMbcA3Zsg
GfR2HAjyC/lHsR70q4/N7osDX9TcryomzQwlh711UkFwijdVe9Wg5cmsMVubRdkj
r0AvFoEEbwTlPbZvC0zvQP0fZWYcNIh5KgHoxC51EswmiLWKRUWZrnJ983itCi9z
DFSRemQdtU9Fy0c+f/9gKZgskHGHYQn3S7ss4kyilifUEVrQfJpLE1SRTGlxw4VA
4HkWZbNQ0QK3l6QnVTKtxDzHhSC+mYZKhe/2vswUAMwmylVoBZpFdtPmBO1Ye/r7
xmCQXLQbnA16d0Qrf4WWlkK0ky4L8DoHbdeT77MPIEq3GKu8+vAX09R2SKbAjk3B
wSB1SrGVyz+2/RsNVLqVmT35Eux/hV1DXFxFlK/FJsc1QwUcLsmvuosQK2FSVxke
XKNcqFqx22mmYEiIjhUfYj5XE2Q+FWG5QVw02ng5K3QQl1PYhlhPF127LzZziLI5
g3c9Zdl0wNaMLypSc3pACVwZt4mdbAu8znHWCj+harhLAaOeMem2MCAYkHKNs4Yd
RWw4eEYsT8LxqRa7PbaLuMPzNa5f/GaP0Gem4g9a4W/sRHriezpc7Ef4jkKaBqTQ
/FsQCNdiiXmT5JimMFa88h3Riqmw733eiO31G+hlCqCAg4UNEoTDt9qxlTZv2dkI
YLHP01jaaihRx1CSLVRoHgWYM3C8x61zROifO+Nu8GAEs42HXYVISrR2N94TSahx
e8dOu/zjulZZbNzlrNs0vSb5KEiIqujAuG5VsqeI+oL2ZU8RVRdoWfM38hyfo+3K
Wt+VBBDBSFQ8D81nVzQOXzOrsU30vfLD6tDAWhrYnCJoBwyUxaGmgxMOBggXiwAc
/8gUp/BhAzWMc3L9yFuCX2vM8NVamizUoyK0n0kbzwhAVWyoiyJftcj1gTm2h8pg
fn17SwgSazdrV9/UjaD0ZSrVyPbZRf3+7KIdzR8/3ToUj7ImTPBkyrbwp2rnZGst
OKRgGh8RORDbISaLl+O22zReBaZHdph3UxIuW5Umlm70MbdFFHYv7eGSCEtdXxmd
FH6VylgDKZTOLkXse+65xGDhgf8VEH/RodjFXgedBM8meztezM34nRVjbQQ5y4E+
DYqj1GgI5ZdyAyjdBTNqf/bX1hkllXqaNU9xYy4NA2n/EBSh93WkkB8CFg7bcV6d
wjoFQy1k15N3k/NX9vQxBoIGYT9yeD/WVhHO/N6G37kHsl8fyP1FWGB5y0CGzJ03
upi6z8cAHyEL1hHdSaP4q8xk57IDS+prK9/V6DscgU+dbL/296a4IRQ34ETzyr7b
HL838G/x6GQlTeJRlQksWmWioQDlwKfeVCcyN5yKHtAgeWElfocV3sPl+MApoTH+
Sj+2l+TFcVIVbVGRd0Nz6FaSNWBlvLv67pSZxcsEvC8vDfUvlXaWXRv0OULyoesl
+IgEShq1yigNRCEznqCWjBDrEDvnAhTLNj4I1Xo+vDd7GOgaICzNQdyadlfFctit
P7ZGs6PtrYxSIYtWaLIb09v2DB4KB4iEktFpDKq4QFpdxzlhFuOdsHhNftwsG+r2
5ud+S8CcNqDLTm868KpzYBCvoW0MjmYpjkJ62Wd/wuN2tx44Q5Z349yop9xeDqZQ
Fm27qaYdAFnO8ckffL8pCjty0yh5Q7iMlEp3qVVBfLWLBsc6eTXRCN4gTd2WlL+A
/aT6vbe9TMnlM2waDI7JYCZAYgawfDH4mIkx9zY4/pVPTpnNn6wF2fsNvoqx1ciV
lkffnCQo1HxTGMYhQgKtrtLwwZrJOyBpoRn3r32nGFfbHdD2aIe81vXXX7ZRcvvJ
oLpVG9iQ7ceTDwUo8tS/Ng/F3o9XluOWC+AsfsYFPvfQSaUSg//GjiSr9mAa5YNl
nruch4bKdFuF00n7I1l/ZNmYV5NNPg768ERqv1N7ijF6fJUjBb3q4gpCGhd7t38h
GRETaSPRORIaiutP3esAFpyjsY+hDC48f2ZNedpQ/otGGeyy04S7xRmLN9czxjYa
0LlY5h9v0Z3TyWdBJlGMei/TVtiW8uOKHJf+TkKJXsafiHoaJq/kGkm/MaeA1kbz
s1iTwEf29rtxub74dfx/BdllflrGh0NpgL61qaKn32alKYHEr5X4DVCiI+ShNsUs
NDOtyW/FrflKcPLGjfDk/eYnC5dWldoDS/N05oKn6V3cGaJkHGGxWo+M4cwTsfaR
upkr6qvlcLonVL/gGF/Rvxn3fgbgTVea17xx2jJ6Jf1OUbYZbDiH3TGoHSYmFhP6
A8XpFjGzkvVmVsmKznLU65v+8P+SrmD45kRgiGROGNImNN88gmgQMkv4fSecQdOc
G7Szt2ZNba91miqDfHjZ7PhS3FpD1TtHa8UB+kWqouReojpBAz+mJNCeOclTrGuB
NUVqh38AxIxOHihaUroV+AbsRuMMOSBuOX45GYzvV0ugj/UwJIk7KFoOEn5KwKGz
S8O+suksXBS1vVR+y0/xLjC0oWlGdB7Vuu2XF7S6gGml7+mNSBZD3BmQNuWZamHL
5DETBKHpZbMO//Sym0SxzxU2+UXfxt0Zsp2FKx7vQJgE0nr+YNflSo/V9LiyhuzP
1Z1UzrbwCqysg/X1NHlh5+Zh7EkfhVlXuhUH3l4wP9hpL1V1VXj/jWzcIngPy/46
fWCEVZhCYh1Zj/S+OTp3PIKvfgyDIUewpxVv0MRUfCc4tIBBH3qshcW4OaqdpHgf
0ZqQdbga13IvJD1KJFAsDaxVW1wP9JWRrWqppocCRb6JnZwk8YS9WAtrn2Bs/q0s
syk/ixelEdeVwUuqShHI9noyQ4A8yWZgEXCAJtc5dU2Vy3LPw/RF7dpiTHepLoUy
8N2gYxgsEeOkVy0EKWOok01CqYOJa56DfZnUvUmVJsWKyjXTNDqs+oZV+mClpdfa
KHGfcQ2rNhM0HT8zh7YWy3bqrjiPAboonzUbPkw+zLrHzH/3hbz829dDb9JBWiF9
ekLsSEra/+NkEBpdvoBjEdGutZMf6Z50k54YLznD7N+KfOtnFizNtFKJ8w/CfcoA
6mjbdgnC5z4NcBIti0bFQp5gorQqCJkFd6NTr8rfyK5X2azdC4fiH/cE8LNyodfe
L/yo/ug459viEGUh3+DKO37Q6iR2tnzTWWfqe9pV8mOXvwP5kRl8jQK12AG+rlZk
tkks3tw+Tp8DjMssNYb1VLCVmZ1rLysZSslu3UW+i3sNk1/G9mZppCBWwzK8Q50z
iEWSsGJ2KTjXlrj39P6piQUhlA/ik/EATOW9ynLhsCLOsAOE0CS9kBYbkWbUwz68
w9sP7BngFNe7iPjHZn7YBRGyXkUl5WjM0XyrRsE1BtcysAkWVY3INuk4DN0dylii
44OMMotrtBIlWCqux+B+kSxBej2NSHy/1nqVYLTi1BRU9TQvCSIeNJHhK2pzXrdb
bGbP4FyE37AOxGGlfs32jc7PA+vKDP/wNY3uypqlMHbJ5OWXqEtWFd8UyRIWoUlz
nH/x4b0s9NrfgGr3TxOMO3VtvBjtgY+Nl4K5SXpEDbfpaHT9I8RQgWLeKo50UNvI
dYRKLXR9IKxWk1cjxeYl6SSIVupsLqgqeA/djrFWrehO2+04ZE3LMZ2kqy3m/YmD
7SjKb+OOQ6mQVdmFFVdar3pYvPPC8XIRKdUn3P24jDVYJEaeY4rNPuWjU9iunw80
Ewcxoqb+sVw//AH61m8nDCSbt8MevCXCltXBiUT+HiHde13pN2VXi1bzeBEf1k8Z
XtXxve9olSL8AvlFbozhIV/m/pa7EhK3VKEMMRS8vVnVhgESfeALLS/tPiS1E4+H
93RFq2ChmekTftZvdxPcWr4JevDOqh56RH7C1b4b1/cYuXo8JhAQJ3EUY1tYVTmt
jn+OeQOqQc4mIMcaFgkckhaT/9qCmh2rMFWj3E7SVhR+8g0Ad6o+WLQJDwCLsvIv
/LrPyihQM4tH7ZHe8SRu2D44e1MYqkT6yoHjffCm/6LZEJm3uU/FK/0/ahEFITKC
YdaPevKxgDhv20pUlvGo8uCF2oAwsa652fB8r4QF2M66rgMj9IhrSC9RCRHFbsSb
2OeNCZV6yBSyZ1WeU2mWr1gSpFhzktw4DfL+59A7f8y2W0hv6dIeBcMNUpm/JZpC
+P2wah18zkPlBoQxcuv+x2ZvicsgeNCTpu+XC6I/k6RtNGsv3OLQL8eh6sXOalgR
Ku/+nhtquJVNYqTQctt/Vw8M69gm7FDnn70V8pJjXG/up4Ls9C2OaflyitLlfSdm
heVZhx9148HjPK6zgkZHGVPWF3QCJnSvyPDHVJH1yLGq5ZjsT0UgsuYwYnLF4Sbk
cou/a5+6tlyzk39KO5hxJGKJ1vKK+HMcHBlpmnYbuqqf/14Qd3/HwSpYBrlbeCQf
QHFtzdR+Ozb1AgjwN5uLkebbzLFmo6VvO8O80llCNKf/Kc9+ksxcDJMuuEScV/Pb
N+5tT9qIWl/LYGyq06zQ4r/c7HNWL4OGbcNvtvTaYqnkUbX6qOY8sQTDHzreGyYB
8w8QEEzd0cjYJwzn5MAuOSS5jEHo8Xl4F3zyhNXOMIT7H1ozhFajj13nAe/naizZ
ujHa6AjzyeQ3K/FeKeBYe1d4q4irjbWHN52hcJiGthT1TlGvWUnapKB84p/awDSC
Gr4gRmctulS6Y5Kso8xJ36qQLh6+zR8nsdYhORj++xGmaU+s+HnDNX1COhx8W/HT
HM6lWxPf9UNcQ5zTFp5fET7rrkU7CysjRp8PetoojA5YBlS/kCDYJOZWX8fk/eXX
562AcdkSs2mrlPybie85Yb8k4JnYMXg33BvwgLWy0VsIyEyqmkKwadREIvYJ3lrs
Vf91VHu3XYmV/4+meBc7j8mfXovBqH4D2XXkXf+UXRULz0KGkcAm8rdWTIuw4HCk
Xqd5FyAf9ALJ31RfwXfjATqgQdyxi0DE4qsSwh8QHWSV2MJjZHtS+DVBTTkl1Glm
do8ET3twTouWdl5bi6FK60KM0M6qrNFk20vmYStXweJxjUTN+OQU8FlimjYWdqIb
93HVe2sKqDv2RI/7+OcKEks9IVrUcODCurSm+pyhxdt4yrAOsQ4ODYYj6gjbr3jV
gI8ppnMbq9AmIEUeyUo8uHOeKhvlkdHUUzu5XuJWhjAaAr9oYkG+Te4r7+WDD6a2
m/lX2JeU6x13OXeXouzGMziZHBfgj0JpnezvEXhXleakVHU9xGlSE2MgMRJnAxOQ
J/nhWzonsJXwIb/EKHQYfMg1x8iuB1JA5DJsLvN3ejiRieMl4xgZCTuqvgj9EZrd
/W90bMXiludX6+/t7tAtnGXT7KiOeWcocaC1IKbK/ScGbGFIWut/NwWBn0cWERXP
8xdwr7W4tFJejbJYpqeQq9pUFn0LsdsG969LWUDPHhET/LFqsmJ2CCwJFT8DcKGd
wC4zXEW5ESkH5BjESkQpEiRz62Ets/uEo2qgZ/kU92JdC/Bbq0IOf+SUXGzcViA3
69Vz5GHl9sYp7euI1kQ9KbQwtTN0qcn6BuYtKfVEmGe4ZcXvJh76p0e7Iaz5fDzj
3vTQl831OjRkctB7OgpfXbWK3VKlLzyYGHoIhH4tjDjOlt6vKibJzmUnngMpmh15
4XXE1M57kEj97J/xImta+evqj1SBWOhu7SgLLpy1ETdhMimkGFdCI+ZNU0Aa1ztq
GywYf9Droo3xBnCgU2tdCl5mI7QE1SFj7BMiMqqizDYOQbpZsF2HAzM83Sp9BhAu
EmuE4TAnPZospAmN+fxV6PDs7HkYOuEQ7TPPBzLyfTYr9VKj2cQXHNU6Tm7t897G
AHMhFkEpEl4wW/BedrEFdXkSdZrcR0OY2zck6VwIQ8VOj/PeDhM4uccKq1gHhsVb
oOAp620YGBqc9ZadOXRZfkJAO9HxY/jgCLBb7n1RcpiTPaqGAtwKtWe09+L2weon
kUdQfKYEBhZcU8rTQpSb7J16sesWSe0tcSyNneY7EHJkyDCO36w+ZYmO6XdhXXRZ
4HRmaour2ACa6x/Zn/OEkw5xJw3/3yaXvVBDM/5SdhvXNKYmyguAyISe23eDHGex
cI7G/AOdSJiSxxnKHYmDESR2zsgFDkCHZfdXCcO2XM+EuDEQnAOm+tNlJEaiT2Zi
sLcimMfDtLUeEqJmvhb7rcHHLZCIeGDqLJ8K1u85FAOlRvCMgxeKcIX1Z5dJkblj
Dg/TDIyiOCaE0jbH5ePUVlFArDLa3mm1fmUAy5v6oJc4bl51D2807Y0W+mtJ/3cX
IiYU7u4zvewk1ZFxlNDWmi3q24DHM+plIZzPIaJydWVPJ38lHmDZk/9K4p57oc6U
D4IK3tqu/ZQD74WGNq4LPD/PqL1BRmmhJIFeHkhanG1wIf4+qrssu/tvWPlCOYjT
1tn2F/zSXV4pCtibwTR+PCua9x2t/1hCZec2NXxgauLy0zt3F4ZFpAJFVAjhqEcp
wX3iUj7+BNebOExIgAGCEQPDLfUzkORAaR93n0kgxgRuhlwKo0V//F6hZDOySzKp
RUQ5Z7sBJHl2WzaqMs6lpqnuF5v6UYoGemUQr8Vao69AAsc0EZUuBZeLfK26CSRF
L5mfEgbMvN84n+EBR4/Ig4aA48Msu1hTBsxQmoU4XdvU4YnlsT6qxvYWjOUMXYu3
KrjMgk3UKaN4AEgpgkMC3JWJd+GOGspPU+FIvItCEO1IdNGUyiADG1xcrD7Iw1Qi
KJTEtKCXThtaPQOQ0/mCQaFegOtQzA1KdeaU25SgYpvh1ThyvRrpqaEN9gWATWdA
Wz6RV9eMzt/JpoKICInFcNieqs3G7SWbSjxrAGPBzJ8LLwq91nS2vobt2o4nQK4e
bEYVkEJVeY+bWN6khZ1AWZ05ZOFj5Ev1zwYFbBGkSaZCuL0xCrBcsrpYt2Bolkh7
XTtKaSgodbdYEy71dgZwJ+Xm3URfeo5s/0b1Mo0wlKzTnDpG2b3lx+tXPf/fFoyl
3EchVNkUle4C1U1/2fc8hv6mRSGjyPzwq02QEk7KtL4p7/gdYUSAY8hF9SSHWVx0
T/lVhkcmZaZN79ltRXgZ0prbMjSFfPXvwPWjqbl6O4gJnuXxSffSr8/TSywfgrUA
lfwXxrsCMBbctoH5S6Ma2M3jrko/VsOVUIJuLQDhpoVsxths7WB9whSbJElihkrh
awxhQniR84r9UJv/AKJpUXl4OtYsLfUhTxPi74gRH7PlSwzqk+zZEi6mX1Ti7fMf
FjCXY5/jtuJYnTV4Hl07xAQ4OEXXrbIWyTjvKr6011TzeXfVK++s0M4YxnZvU+DU
u3nhgy8USEm6mdjTnWuI0yYP10vYBj9LX+dWlWPRmr7huoe0XrksfMqa0NJCBN9Y
dDqyF2LH2XeuSGF8Q3WoF96sVXcB5AZd5XYkg8kB2MDc04UQxZN1Wfg3kd7ChfOI
W+UcHGeFzohTpbp2mg1Vx8je3wH2z6Xjyt8EJADISuC2FpgJzVFJARHcJF26nc5c
MVZBmm/1Q/s+exqPfT2QJJs2s1BTDsOpMGvEnxloeLmVjbo3YFWwkzyKZFqM+gFP
07fI4FM/4jqe+I+Z0ZrOafts6WAHnffDaewpq9biItkbArqQ1scLRUXYrEx5kcpf
WbfQlB+g9fOO7bKjSXHJdsHhm8CzMV39uoB64ylbZX1qSjFEFZXYmbpJLSs/SEu2
1ikoIaLHXvwM/NzhWRr0oMTKsHUhhRIOqWAapRHZbB4ND7BVziKUyWJUHKmi5mJo
I06atxmFmFDG2iiVi0P/V3itXBSoJD62019LsHJfrMk+w/rPu7nNA9DcoWAHUj4l
x9AToz+ihdUJbxhCbTkszbxaL2CuABwReJQ6mu513Uv+Q0OtAia0v41xHx4MAZ+w
P9KErVkBGdX5naqpr2DXtd1VBw737YlbjpofR7/WSrso54JoepxKassAyrFipPT1
58CW7KWwiOsAllwPiQg2/ou1kcRC8V99yGx2l8OiUvic/9AsUMSFm8rAuTKJAkDu
HOj7jcBMSVl4lHtxUmbR3ENI+Hc3KAvI+OrvmmhRb7UeCJ4vZNJeq1JvHlMr5Wnp
6kILRwOaB75kC8xC/WSa8Vl9TO2dB1WQaN+bsLaLuKK/PiXoMXxrGDsQ6NLnFyr4
LpP/tHpIkZBmTiwauGag2uSCSMdEG+MvOrln1irODCx3J49xAYqytaPwueAb7ejn
5ZZWm8X63wvMHdZMyNqwJIzK1p6IrZGXBDSCufk3dJoThbibAlNmOUHSz8ln68mp
3aGM8J8rwe7GMChENhEyTQoIPS/ATT/BMWzklLMFwI3NM6c+y/t9i/sUEpOIHht6
dFKt9NmPRbFwT8fM66s2mw2HjvTbwoQ9XcQ1sW9QKmXq292pgL6APGx56ikdeJjN
gzO/hfbvRZ+9+LP34sIDeC4FgxLlspLCTJ6O+S33WhKamnv3SCT7W0c8kFMyF9nH
bMXk0aMZCpXiOHh9gt+bka+Lhw5sKb6lswYZYyv7z/eIzwAMQ16BYFjXht+5uVFZ
pn6HfKmMHM2QtRpND80EKtYiyRTQl+ukzQ8MgL5wZP03tDm4qopRun78Q1v/WMK2
F4twQ6QZa+ya+e4Jkw5MHLWrp6AASC7wSsDiFHr2Nyw1D1Ze+fLy7FJgc2UT8i5h
Bl6A9MIFSTDVVn0LZMonbo2mhmbVirchl4Hv7AADEn077qTwUZiSFJGEhD5mH8o7
qX7AfyhznbV2Q8mgrrERKm8Gap183M/u0BITtXvyiHjXamE+JNbHeuLDlUIKRr2W
tdGfyl8yBbdOtwPNagbE+QwGINmWHHnMQOSWqnUt9lj9z5aSMRjClroxcdtWyRsm
gjyuk2EG9oCD6mQ5s3HQvQjqOnAVfpDRslAZN4P6yIm8Ci5hauZYLaGVt+qbPiDE
HIf6XN8oI5TUGl9fuJy0DipBqSwPaBYmt94xFaw4c6TxKfHjODGk1ZD5YYvRdc+0
UAd4TZfea3DS6TAYj2kkv6tTB+gQT/th+i4El9ikWjTuWgBLZFqbs7VK18muz0/d
6+ogYf12Xcp822u4CoCBhCT1reut3YswtRURJXDbaXpQMg57AOd3bGpVXxAzwG7R
Kjnev1YTz6GzpScJ9GZxNLncPfezMIypxQSsP3NHF6ZARApZykELrSy62lTmgtjY
iYOy5iZ20pqJaajnGwuNFBvPfwpVQRrErT3rKKkPKkP0qlVrXZgMx0k7dPk9kNaj
DqarckJyCohoWdB0Rx8Ma6QV3Acfz5KpunxodAP9cigIjokiGEnFiZd7Fjacaz1J
77UJI7e2OoUiMrHmzQ6J4nlxuH9ZMbkSECERv6CuNxgATDLcuXFXTxofkwgIEr6U
mckMs91FiYMrIFPxETNizGp0UDNjzl0Kon0GCLqtkyGgZzJW6yH3Wzv0hLVhDlg1
O92evtYWmqNG9f9KJkHBsaCp1WZ/35u36/gBG9ETpSY/SnpR38de1dNCHykMcGWN
hISeQo+Y8nxrWr7gvcAz41XZYc23grWvfqpW1sijJMhfNrJRfFz6sTBNwuA4m5ia
+BT0GCY+6fLSe33dTEHu68aOiPr+yrRUuCa51Mzn3WmhZvmsUJ7JXD6snFLhYdQL
+uYfWipbRRsnxLqGagj10zqlq/s/UvwMfvu0VASsNwEOto3nItPOIc/J442YsEf0
aCsRXy7bjAjcJHKmsPscy30zM1BJ6E91xB7lMOjEjmX4pbhm8khJ6N3JC7shjEnh
zoczb1mHnb9vfVvoi6M1nhfe2W9FC5aW8Vr6vED9QO9QvGLahw/Om8Ile8BAEBvY
UZWRxlI+Benborl+EOa7EqBSgiNt/pkzYTxW2RF/9VASd9/WG4mx5z4oANQ/ZcKp
ryFxbwMU/pc5htjAKKNNdu21tj8o8MO98eJkDj4D1tLHl1BHK0eDC3xzHbFbhzMA
83RcbGh7iUeHPSdSBIwys95oQLHwiHNm9Dl/WmsouZV5EpjI6jr5QF+3oaZEhNIx
dGkn/Bq//4UucHK7BoZYLZptkIv4oGsDhFs7sEq9aIfk7Vgo9rS6ANJT4wheB+V9
G6LBiJB5Uo1Xu9xxk/cgcV+As4EpVHsCQvo9sOdRuLogtDMmAXbPdRHGbhEfiesQ
fAYRV4LMezp4x69iHmZNrrQqrvyy1zcRr0Tzf2tczv9wT3sst0BpfIzi1/48zrbs
iNgpSZrXzSEav6PskzMZpx9vpgH8GEqK9meTr1jb8he2yAWav2xiXvX0y7clspYZ
Qa+flvSyYLbqKjDmezlCjuxbdH+TMr4DOPFi3LwiJTHRok2Igzwcbb9gGBx9QESM
e5YfNYbBMk0yOZt9YK6rECng3y0P0BXo6ImVI3nl+NisqHlkRca7fJIf92zf5sgr
DHtvp4dJfDxoat1WgrKWSOak1dF+O0YWuSWWvAI3vgsn+jiKIfk/wfc1Jhyd7tuf
I6YkDlwddsCO8VjaRwdRkQrFf49Ztc5Nq+G00DlzGDjyYSon6oS2eUKFmIMmCHIC
RcIFFzzTwpt0kOPgb5R5wyn1RbYZRzfG/1QrHvUIHH37Pq7zE+E+n+mpJdJQsCM6
CcOwP8q5nrTSMWoaa0L74Fwqy7rsoAcgSnCOZ++BQONf0odC1m6yGRcaP83eNfOq
MI21FZLzMdN5GuvtqBXunpWPq9UG8fTAjgYsHtwbGDMuNs9NsHDHwWJc+KxmJxOs
q1UBH/PseHVCdm+okIX5JYbNX7P8OFQfElQmDnhIUA1j8RbbqyLZFSYf//KYKw0m
0LlAP2YtLf/O+7ZPezsJxjEb/0eSoqya7F4zPQpax8j/8WbTdce+xQkh7vQGUpuf
l1umNo9LJNSULurb6DNHhKyIKonrMVEYo3N8XjcgUIRd2QYU1R/CJbZkWJFyaZuA
uHU1K6kuqbF/ytrRvYaF7sTNaPSUFxbHlTJKlXBAaneprSAs5ABOgIhJfOqLGKYT
FdNH4KRHntknaDVwXbRM3JPJoimvyL2ZjA0voJdy9D+HImYslMQprl0jzPAHNBUu
wGG0Q1695DJRJEZ+XzkLFEOCnAtLCL8Mx/Sen8FR/V3Rrb5TO8eBJuSsamOCva/Q
UurKrZCxr9IuBDwO1gSiwm5JjRb2N50PpU2ZfSVFIg8RIpTCBSYlcgV6CumGLwT9
HAR5/SoNTLXKNVAlFE/RP9HJZt8iQGKQMn4Zrn6b15WyXtMvPydKV/kH/6IeCU40
YrPI/oO004XN7cYoyVD5aBVYDOiEaCvL7YwJqRwtSLg0yVT1uNs5aQNcXOWAggW4
xb1Ma51HFHCkiO5UG2myBGHkejMCfmLs1nMOg386a1UKErrKcCuWnn9fNpbnhQIm
UwyV+RbrTm2da1wQimLG1FsqCccoiBLFg1AWHCQl9M4G3Sgpz8+2apf4po/7e4U4
BmUMTDX/ugmFs83Fbi6/Wyl/vKnLS28FtfBrxMUUAiZr3HcIivTRt39dg+fXda73
GtI/ccBrdq4EGDDopU0hO3XVplrjsaJMd+RhACiIpD/yUkOO5b3kMabOuGlnUB7q
ECUNznggtGBqC8uxfvkxSCUhv3TrSmFzC2Wi4yr363C3ihHUI1PBa8ntoTjwLFmA
IrTczZ7TX1IvhAlsvaKExHzEZBqFveE8GBMoQqZJ7hnyRV4yUHCnVTe7tsjL9ZfJ
CKyXxLKzpmDb4hDQ+vc55nQlH3gBBTzoWzwPo9vk3xD4lS6+RK/getdmyyTJnSY/
p3NXHr43DrFp54TijUnjlYZCTcJuzywQlSDEd5hYad6W9dIbN2S0e9SPQnunYGcl
gvYJnIEMQP22wWJwj/MCAAvgTBm8pSOSNpWsC8Y09PatzPpn/ygYOSDVn85O9Fu1
61qiqHXxI1Spoeg/jg6PsZLuiS2vhmVxYD4onvpy7wvMC/gf7kQue9PFN5QlWRw4
v7+L8/hS/u8lz0CHtMc+uhp6weN3DVnSVD+17PgyplqrnUaGfdpSCca6T72wOUka
QAjs9e8iF+YS8hfUfhgDcLCNEDdlFkZUz+dl9wVYLaODuUkhbK2FzKAG89XZHwdb
Z8ImwrhoGWCk58ve4jpszKz0scDPVAtSjHrDhCJeR61LRBhJw5fnGgo7xNp8hQhx
RGdb6J5+ME0wqHJY5U4NKaRO1p47h2qRz9Yl11lDJRbgYtu73EemI9DwHTe+oVNU
OTgmD58BG4KtkZKrccF4tsvfn/nmmwZSPN5WYWgXYqIGDqxR91Vy2tIM0zdqnlCJ
xxJzjwPb13Jji4I2/fhhbMsC+arBawkvNkJODR66NyheXcoes7BFYFizeQb1szFA
qQXN8XQ1KMl3LAIeFZRuYf+yHpJWdbzxcyoJED1JiPctmReUZS3lTGXBwMAo1GKX
VcwKI5oJDHoxjDSpeQL2B9X2DPrd8Y4lf3HwvaAjIhBZbr5yUTT5WuHGLAaIHSaa
IoPGQ5m4aon5TraT5Hj5JPYeemsLV4MjrTGepJc9XXU7FOnjwltIYVsfD4UK7p3u
Yj1+vL84yFtBEU0Zm5CQALx52Wf/9pWyVdgC23JctxcTQ49VZix4wTXtWdhJdL+v
4/nxHfQD9VUw052u5GGD0tF5k/4Xvi3K6TCT3T060EmJTjCWivPp2IRb4DH/OAcj
7DJimcQIUTZ50eCQ8VMVIMkDERA9dRoxk22yX33rynBebPo5v9m3redHxDE0dTq7
ZbI4U7OMoGxLJpaYEdr/M0lQI3wE1XQeYuAtCLZbF4VWl3eqiuvFRP7bPgwUplZA
kjH6E0tmxJtmaZcemI4srPD6CGtB2ZIY47V7WA+49gS1Yr5iMs5umr4Fp8xL/VGY
KlKBq7vtOTqkZtc6Spp5Arc8XRWbPBihv2Fs0s0qpFHMTG+XFN+/USJAW1rPbdsA
VROGRSdaJDyiIHIYC0ibJZhpMjfvyJJt+S3Ni9lMv+S+VspQat1TCG3v36txuqAY
hJCNzQI/E/yLz89Re2YXySUCJJOX8FS2iyRLtkg29BbV38BW8YJ9rS8O8v/APCOt
oNbZ+nda1zgbYFwohiUmC/8LGiLweLeER/Eew7D79GxlIsGXrN2uM28ljcJCX8Ld
EK55ahQef0lD7nTIxu9lZREEU0BFofP9fJEpivHw5YXb/qMQ2JPsSZBXBgJ6hCwk
yGkP3Ire0tnT2v+huCqOAenMX8a8zZ1cFlZV9Okka0U5e2rKdbqkGE8gNMyjFM7O
iVvcYAt8zvYWoDwwVANJ6TE/YMvqw19cVRP1Xk8/UIZ5IsUHewS7P2YEEcvv+Ndq
d7e3M0dFtTNGJOv2aQW+eNozkv0IOUB09/L312GZdUzddFkCXPmU1r7S8ZLH8uDE
DrETCH+ny1B4c0rL0P/r98GfYG/i+EWSGiwc5t2XbTVifejh0Ui1AAwTnbDnDDX0
MNJAdh7mKtYvLpgzRBPf3dPCSDcKT0M0TRbjE2i7HVeV/8yJ5R5iDL3WqvdpmB6k
1f3246PSfnEWit54ZcUp82fwLqbuS5+NIUk/Q4ygSuuWPykqPnFc3At0DxkcEpSg
F3mY3DCbta+djc4LikeexiosvD9teiacYTSGRVh+g5ZmOpNi4KL2ALx1O67LK9L3
9sGBneazWtBCgdHjZmyuuxL89zixEFyAAcuGJO7/1squ2LCGd4jgyvOgoIe2B5P0
+028sy5mBcgoyiStdnw8E1e/Ts0zqGTuzbf7nVTRCnUS9zfLcLKKcqmcjxeAi9aO
reshTvSRNYEZVgvNdFh9FFRu8guciWkKWWHYIGN+WdIKTnkS4Nqc26QY7JiTMi4K
k1Y0x4Hl1c8cQd+vJPCadjWP+2+CCLs21oOrHwJDugEWtU3+Y7lrMF/05Gx2JWJU
rJq/zYKi7vFlOqFJaVwZBREtpEdxc2A96TeO+jUJXgpXbazwBzDIdKvzdUVwmyqe
Wz78F5zR653xR+UL0ja+tRrpLBn89TIHNTWyqaT3YFxliNm+ARltdZdvPplziFKI
TBMG20HkuR/k1lc8Pi9ZLGpFCru+ey7lJwmMYfew9a4i8EWIY/qEMNaHEtrWPk+H
kTvRwyW2VQ77jP8VW+/tcxO5BWNq4tnHv3F4LISiQIv+0lu/S4a8+kRmfYmVvzcJ
X0VpUxUGghpwSTOhM+o6YvLZRoO7cbof+Sqv5T3B3Hf3sACsNpNnli/nTlm1oelO
6QJMcRqAvDWMaAcgT80YKCCnkb2fbBlnmar99e1+XLq60rSorCkaOzk+kc15UkA8
xqLfcgivmnWHJbSVuh2I5KHZxglJfDpVTfi91a6BhEkJcib7FSlZKqXdZZNacwVT
qa9h/WAyvXAnWu+IcltzAam5/eHcs7lLUuxOyohShReOCiHgSo0VIZoEXdOQNLH8
eZ145u745jKajxVEzecLTa3MVIskiomOwX7p4JKKUv8AmSVc/CL58GQSeMTy6GR3
ZCVgrGSoPDxloBW+oCCqnSN9hgPljZTK6nsFFk8QrXCyoTCPRWdt/ybhg6H6SzTQ
bJEZjRCihS1P9LfLaYHDyYyHM3T/HosGS7VcTFimGhMq0brcnhPYcIrza/t5r2ka
1WV/3qMPcIVQLBaLQulki6/uWKqX5BXzM/HTHspozvf0yEQKNF8MuiV15AZnU/Y/
PLSTUNXEqzZq3mOR9Pbx9EEEcE4dj+NVFWHpiB52TlQZdKsWkqoHd6D/kZ8qWd7q
TYJ1In+Y4HeAdz3vyH3XFROLTh1JKD0MDaXwkWUPKOPH4TtxfQZCNnIzkLzqbVLN
i1u5Jro48eXy8n9SiIwkENmrR5LkOn9E64GlA/TX0tEpFk4EL9E2yHL/vSl5Hk7K
AtBhwJ8yWts8fgSOGTGbQ8Vex0dHB6MOsrXsd9zYzQxgOjFXkFXXEOGANY+w/0Yk
nWen93O/zfvIpBDvATLm9KGDv0ERaKqekVDjRF9lGq7TnDRbP3nntTXbi12OQrT3
HtuVD1vOHhrmEk+lTbxtY9dKe/2b8a9uwjyd0/Z5udmD2ojl2r5PGcDwxNAIx537
ZGWxMdNsdYsBt7RwJ+Gh46dHDe5xmDxustWn6yWeM+JEVWB/d+GfchQYx8Om4O7F
Z+y4DTZh6Af3aBb6NCXQ2TiCWXcMTR35jOjkbBhf854BK48KFRyG3rA5rqqiI/9F
qyVQTAkBTW95iVCUFygWVCeVq0qI8J4/v55udsv++WCcCICKLS7Na04krXRWWz0R
J/mPKT432rke/xQqBT/Zi/HzBhpssJMMyY1tfSoxs1FTUlEefCpppw8GzG/zg5hi
nqSdfPBXweazWlKvBYMD1xN29toETTq0Eyi0mhLP8H6EtpsJ+hHAqwrTZ3ekxS4h
8mg5WnWCZbiEFgRrir+jq9LSv0+y8T21TQo7M8AGOOBbiV0l8LK81NxPjzeeCT6x
tkHSMaVu1BUHrZizabPs7XyWsyN73WN4pgNCYU3+2jkL+4dMwEeEhDV4iDzO1k0K
OsInAfKTrh1eLewC/3GN05VKCncbcqVEw97nCHYsJzcg9nb6hXoKE5gL31Eczk6u
sGSIOMdemUYpHNQ8rmMlwk1ilfaxlVr7/swPplrqLcJgQ3BkBFAfEOpyT7rh99fi
YyAI/SRxDibtIcocLAoDJNE75x81BNN07AIM1U6XAtEc1DbPOgvPa5iu+H4rrYGZ
PFEbOzc9FbkfbDgJtIqcY6ZVHXVfyUKJx4QvaHHyalLwWmizLADxe4S/wRzRuGk9
Fm97EPDnB153Mfr3fSMofxbY25DiwP8DoGNcp0dSRR3VgOAFMInSXxicEqPH6UYT
+3/N0Yz1b9OrlQZfK653V2j3pTMSuqNArhzNAP2Pjy4KuXjdsR5CmiNHP650X39F
n+F0RriFZ8aSRyI9ZGEBH1G+v6+Lq3cswsDrdfsyHn7OAPh4iXuNFQ5sJ7xGGab3
1LgRDqUNQ9VVRzvcDKo2Qc5CASbVK500ZYjToN7aZq8REG1G9kHyXi+wiN2+D9Zb
3Kx2zlfDhkg630RHpCusS/Hb9QZm5QcZDUgi6Dgx+8MdqrMCyr0hfw7TG0cS0wkj
4nHA8hyX6cloPhCZLglbU0pznj4L1+DMBmMQ8S6WmtntE1YHT7i2LWf/nHGrbHvm
XmzaO1CNaOlBFMDUTA1bqJE/H458UL81wGZhaziDsrxxSfZ9WmNV+le56AOYi3Eg
ci8n5G8TvfgfoGmsDl0lrEh7nRhRqXt+7QBptgjnllxMG5dU7mLYfWf0dgRy+SIZ
oQnqtD4/pKA/I0qcbQbH0CuuzfZt1puhEqGBpMQnPg9KwN8hUz1x5BgwqWfKkSQa
02luTBJOVJk4jSvEhvlWDh63/8m9ytSRRVC8Xi2XM5eQpiV2qnzua8bgSZDdr9s0
9SLikFqOrLhLLXb1+cv1j8gXYe3Wj1DHuBQs1fCfvrpz+DdRjQvGKHP2bKhgEZEy
jVdiSVNnOUbX6zQbY7VZt/Nh5tKUDHyy6RQxNp9QpvgxPKm8K3kcJOAtgGePkKbd
KYBNRBRF1mmbQftux+gMm5ehTgfKqpt7S77llb62meyOaSSD78jDM0hpcyK12bKU
Rj5At9qN2fTIYivMBhSQwtTpO6yxv14e4i+sRAaKp0O97ffMZMtTY7EedGgTaYRo
m4FnVoJlY8nlRv4IQPbJME9NToLhO9GUFeD6kcFN5NedfZy8b2v4loyJRXoCYn+U
B2xziANs3MULSbFhUhmT6mj0IBwNGFQd67hr9m49Nn7qmZLQXNGK/3wmwR5H2gSJ
Z3hLX6iVka3g4pGnh9DVyZoQP+qoZNKRKss2QwC/aInhYY48iIdgtkcTr/FH29S9
TWLpV8Wi5rTeGhvRZydM7FFT9B5Lg6Yl+clDLWFAUCzhkJ5Q7N4TaQRYGg1IZlfw
AJsk3cmZgtod/Ora+QvOVi1rjj3m/Ch9rXkQ6e9QibzO66qcxCOUjzbmGtV/g0Uv
ajRG9sdL8S8dR968YizN8kvoEbW2jM6LdmmK5afu6QtQzCvs6Xrhinqev18Vnzdj
cC5tcKlAYzm0bWZ8GiJmMRxHMAxZ/TcaejxYK3FwnD+bFbgrcTLZ5wWZcps3FH4+
i0iE++3dF5ymMCPXzH5Z6M+RgM2zjhKajnLD/75Iyh/88hgbXH7I5eVLIFV2rUke
exma6ke1lhKMjD7DVmSbkiWRjr2ICWLzjlEdI/6LFMdYX26dwEQ5gqTG4HDbXOPz
iGPYkPRJUqEw8GpVOk2/Ywbe7M56ofVN+cgixXMVKQcUWj3E+syEr8k0xDZFZ+ce
wi9/ZlgVv8309y+3MGJsG3f+1+B7pf/H8bKNGWDxsxDQuD+9TcHcZQ35Dpl2hvaW
YqH8Jmme/HUpsoH3mm2PxoZXMEygjXf0WkozUTtrqK3y2SxQAMB65DPNPyuBfBjN
FQ5U27BJtba5RZm+lo4S0tQwPOkUs1RhoHYBOV5Xb2C1laUgBaaCJE69JL9vlz1d
lKtT2w9nI1po/D5kZgNtsnL+e08q9vrGpGrpn8Gvoqx9xRDWtypcFRTsQL7iwTIU
RqFCZY8puMAXONGIVgfg3snvgV7/uVyFEXZNYGBvvi1LQ/ydLaqj+mS9c4gxXeYc
7IZNr+l5oUzkiA8KpodlxnRDY1PfxsWUhfPU+YJcLBpf87rKt4EKMLetgky+NePf
DRZfKuxyntf54SHLBaNsYaK5xrqTVjYYMRgk/SX0Zkm8kLolVg4J7viR78j5H+wa
ovGs5PIzZJRxN21h4AIKFQbP7r92QHek5/MrbWyG6hD/BqjW1sTQEfXTtro+KAyD
ra3iNhX9+/MMDXd+FZJGa160YU5OcqFi2GDeEeFbR2i4PRsdU4G8/QYCnYhQLjlP
bmeqPF4dOFI9J+TYOXIp/N62dcXA6QulCm93EKp0gwzAJo3tJ8sez2V+s6PCgaSl
RY205M/8mWecKY4LyD0U5+zBV0/crZQT2AKTSxw1jqDkqh1VKO6l+bq+7RcXhf/6
a2uTgKa4b4tBM95NxES/7k1FWOFHtr/kzSXsjCwCEAwK4Sj5QMoOKkMpeAB9TRmR
CExLANVOsAUlOaC66fCgjRGOb73gBTmziwVHKHRRnUPfFblGSFEkHz8i/qi9qT4e
/NVzNFHakLKkiOll0u1vdu33/XtR8I5sUkBf/uycDbSSmFPicI2zbYXk4Q8GeClC
tNdu6ZgFKDKLKp8NLgPu609627UelqrEX5hZp1FUqUzSmAaBtb7IapjRyMLQWSNy
ffsJod8/3GGRkP5MooOzzRyAXCbDJonyUfNw3NUeBKyF1ZQu7LX0dD5zlHz382Ex
uEYPk/sh8TyEmOD1vtsxDFYuTrNw295OZ99Lhkl4cHNutimQ0XaB+k6V53UQeyyh
++csSsRkGTCGaKQuFbGWPDnh0lXq00M+3xrbcZphS1F9rP+NuPlVFdijKMkaiP/9
mpnuAdvq4eCDXE5HENrG7VHhIrLkC5BvtRKTCfz5tmsNZyr52mvLTjEkzAg7yp4w
M5CNvJ+kP/z6kgNVlpSo7mtAp4V6DIaIbHjrjE8kBI2vhiWBOIyUBx+f5IeBl8Im
eWTMwEy9a03W96Nx6HCHI4Oi/U0l2x6uC4fqmWRdyrIcFaUo4VIU+2LOBMYsoNs7
CWr70n0J6Mg5FYhaVc2B+aq614OJ1G6I4VgYmcX8THUNW6vy57ywCbK8KDscxt0M
s9RUXOgVbjchvPzIeXSGSEADBT91rNfLaudthuHkFJuMxbqlGfcG5BJtJSP2jFsT
SdTKw/89ts7IUB316oMhJKZ/XgHaWCw/btBDXda0cnOkVMcvgtEXm6AuD39JIiIS
AuwIG0W7cm/Ru7N7M32khYQzrnDg2qmgXD2vQ/0+9GYrVRTwPIDp/lVEH4HbPMdC
eH19RI+x3wnqrde15cuzGQtb53zm6kd5Gsidq6v+awEwUsaAwbTdEBOftvj96g93
vsAqPAEjzxeGbVue+dhFvWn7g4Us1GrjPfjPq7mFvE/7jAMlbfKGF0sr/C43T4Xq
ZEYoEoBYFKH3NCQ1eRH9bGFpsmmw+oy08M2nH24RPlX5XjUqRQ7D89W/IyDt/JAO
WPhxRMxTz8Ir+x3ruiEYu4D2fRV8I/yg/cV70j5sqzv5wTVbYgTdbdifpgRxeZPv
Rlspa4vb7NU/OVb5OgQx/aaJnhBsmf4BI6Jax5SdrFItJzPyii+qrA2VfBZYSc8C
WUD6vqb4IyLMDu33S0pFvhujPcOLyIeLyl8IfK/nHGjTN1yrYoU7aS9rNWd0FQif
EqgciWLnq7LbQoP4vN6NoIHTFdqfhLr3kJqcEuZeU5/rC4f3EAchu1fQYLCg6gqk
+cXZzKqDvp+CaEaha9HeNaEJQBOnCc3jl3T6wca4sf3t090dahCqqKm9iQJEpg8N
bTVOoqmAWzQNB7fMhWuLLE6e4nHK5LOVQkDGswc9sWI4Y08NzdySkmejk6SvMYsG
aW0IEXzRf9oJGHo6YQIwk8eIgQ+tVOhS0mtbulLEhy3rymiF4UXNHnI922zbEB91
4IBjypGXwlC2RUIRYwmibiH2IEIBDUQP8c7jINiBeRWIGa9V//d8DOMojXhktXU1
BeAcm8C7vlzBDf+XZtYqbBXhEdr19Why8OSvwaiPChUfI9GSJKHo7Seyh3/8o/Nx
hl5bBjGRkVT+lO12/9wHCyFh6RpAQcQhw25GokocrWY/x8p0aHLJNtyu0EsHTRpp
ogirSHwHZi9ysM0lRR64gg0OsCCRRKfzoMuMYxPVW0adnjor98r9TKtCOcOJA9RB
P/WNqsac354a3QhlL1vIHW2Kfx31mHxYJLebNH/rCgmjJcTK+yHhYaVdm45jB+Fe
Nbm/wWuhe/uRTTDMtYjV+Ditpn2CbF95eHnvQG22TyJ+xLAsE89sy8+pUCOU6P3j
V02m+cWyQFwumAfcy84niEK0ql8gKlKqn9dj18+OR1VdjhPhSUEbaeqGLRtcooQv
+iWYXmxk9nobpP6uAWENdbebcrTPoCVGcSw2CO0EH5T/3CgHCitMPibp8p+sZYNF
QTpZSx1KBdzQDhNSQHA+hJiuTurRvjgUlEwRlt18kT4NVGx6Z/WHWXPoU4Eck/QQ
fSZPIDCha5Qu6l5J3lYTCGRlbjBwgK+2s8M1EoJxuLhIdRMgHBmMVc4q7fiWGEBW
`pragma protect end_protected    
`pragma protect begin_protected    
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
L2PxRyH8PEh2QaZKRzDM4qpzI52dqHAs6+mYndoqb6WHCFIGk1zb2HVpi4iQe0j/
/6TFViETjpA7PQCIHmOEYGrdwQQQZs/uuGGLUoHjkZ2aQQ8RBrHIofjs9omi5/KA
sHz1WY8628Un3hSlc6LQ3flaU4tGoOAPRn7yuh/hWC8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 67358     )
t4KxJI9feigEfkhmBPhaqnlsc67NWjAI1EwHGJSEmFamiTfqN4tC4AbNrLNnrWVL
iluRggnYd/UW7rkDszeUnWbaVlG0oFt6mmyFB5vmiTXYKCGx1uYG4sTdYIxZfoQh
CSb8Zz7ngVGKvRM06dVLUh7+0ChEXh40PZxaCOdaXbAoacuWj/7tRSIfpNGrF1Ui
RpIop0j8qYNZ7ynQFGaN7zpR3oLWIH0X/w6l3jj6zEscgLa7oR6H4x9iBSY7JfU8
yMbviIeb813Wi/zN9Xcr+dmRw90fK7bjgORDQO8r3UH9BysNZJdatoTOW5AN0CgL
`pragma protect end_protected    
//vcs_vip_protect
`pragma protect begin_protected    
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
gfmzYGkkkIshyxAUqdnWz9qQhPM4kKdcZf+x8E5Qhvh2KYS7BrYT9wQcClVk1rHU
Yg22B+92gotK+MHLJw8V5x5B2tPS0LqPmS3/NF5ioCHxjUlsLQ7yAZotNujlWqdD
41pUL/HiUT9rrFya5d1KxqvIzWFhO2UqdkhWqpl64As=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 86796     )
txw5zEUoPl1Frly3O34jyHdHvNSg6zLDxKHOKRRFZeawhx3KKaZmvU8K2QaZI4Zd
a6Got7DizVJzrf0I4UGGtiy9fmCrzBV2qq8bKujELmpyZ4gHf29x/4pZWc/oGLNJ
5hwFACLi0lHOEcA4g6RBDylLHs08w8Dn/3GXORnPSEAsCYr9I4A2DXCrA0YnS5w1
YIw/o+TLTPIE8DGl0mOPOMcG1qqo8PH9AK34BUjj7rwW9tKVc9PsRKaJ4T3NTkVE
jjCvDyMroqPZbz8Ye0YH3PucH6vATQ8/HvRUkEJwP2Tg8dNgXzvb73vf3A5+bh0O
tJHF9/9dJQtLX98RPsrgjSiJXqpqXJ7kpChOxGJQooG8Z2+kVOw2pLVf+j8MHwLB
JYE3lJfbKzsLqy2mCqWE6mgOIC7jPnWY9eI6UufGQ2HbYTmgqeek5gbUJt+ygOE1
rD5SsLqsbhGx0QjO8du9zRfOv5Z2SiZm4/RuS/KodUIs70RjeD8LEe5aWzfzihQe
nvFl0gNN/WXAgqjrt/+K825Mv71yqojR0rNczKqSthoeX7k2ZRn1gmlfqg4etyJQ
VHVEpkY+ni+MW1dqz3gKRvE0PyZjnzJpWvjc8LOb6XtwYsUbuHAao0sa2Y0ZB+CY
fQ45Y5Xx4fde6vglmWjX3KYlrPXXl9k9WzXe+r22XGQVP7OkJPy6ShaLKFkJcYjx
QJSqAU01uAmAWW4DgszTkQJ6D3FoRxb5ak/LNePRtdf31NJ6OzcglDiApt8DsmCJ
35vo1fSvf1WDDlGRJL7Y+R4xySOejY2hhf8/126Ukml71tK4apBQ8s5lxZLjQ0n8
ZnF6IeNnLTb5QfJMBiRNu+MNXHLwG4MTaV0XFP+jfLKfAJlEboHJvB7ZqP6tN24w
C1668OnLmk34UCRjFPyod1a58hfjK+yqbYhqBuXlXjfTP0aANI+v4Zq8c2PQ4tPi
vEBmCKqt9RiIxLbcPIMLLAitDOFbeXoi+qQ1TVmfaCdntKZcjcP4o3POSiqJ7Ri1
dEAYkhpyn2fb0u69A2aieB3LjmR+7B9bCgzbX91jowwNI3a9MVRKMm3Gj6z7nBu2
BVBSDv4WewvzSV1bUVu/k5j69UObRate0I1aG19P4CGNgDKmP/MAmPSBWEXCsJ5E
o+EhUqwOtjO9nkcXHhQ898ZYhGQ20iWefOycQcCr+nJeL6kp+oYJgY0i2jPWMR9j
HcZmf7vZpf8Wh5r3+4xUZmBqdL1WpS5p0pRfyD5YsoHjoFJLh6hQCo4GfL7AXUYr
AUbMKBpK0V+n7LB1/S+zRTStn+C7BdFMK/rrKVJmZA1UWH84fYu+myF7GCOfpdKj
aUQLfQeMkKsXd/qXDU+J1vv/0ZfLlb3DmvYs0O/AXQhjnEqQWCgzw9IH2rYcnxEE
T3CkIRpjJ6FJGz3Vq6syvJuK+Hdr9HOR9PGyy/DoF91cnnzzspB16YBrc28uDopJ
ZyjilBMGT2y8AEPD2CmoMzkpI8ZmN+G5MRf0pm5CCg1SPtg6LAV6S8Ve+VSHIP8e
sfPqfndKHtg/quzvHpGWaDKQbsf5ih6lh5V+EXXegIJ75hC+Te5NO7kzSi6fAi7H
V6t9UrnPX7+9eY42pJM0HVAW04QsRNvf50IBgduTlUQGUXFswK2qzvzvJfwEzrEo
nPfij9xtTaORxoK2DV9D3Z7ydq3OxtsedQQZkta9mrlFdv2Hsuurx/rCctkeD3oU
8F/rLAzDrOvL5Zy0vdhsLhI087ky/p+twkA64TshMuUlJ9UoraaaC//sVSoq40oi
/FI0mFE4hwBBw7aR6WG7Z5sH+uBXaHsr/dewlfsJ4bKCDXzQ2967VtO4BkWhOh4N
NTkeyWUF6xzR7X3qDegRWUpkhrJ7MNi92ss//BKYP/m9E27OYJHlY5XP8R6eHVKg
rkIFB4uNAS2QfULEGU2knlYLW2fk3hg6DXsd2itoYHMBHEiLAlMQvLv41tfa64i3
2M2nv7Km0OL4dlz2LBbYJgyXEJJzx89Zjc8Mo5AYIQosccRWgAC7Mr+C8CuPte4i
bzaWki5mYiydDK+XuTDglPSFql8+yfPzz1iN6eQ1LjfdUpPtFVFNdRlXzz1hccm5
TJMa0lFoHvxtRYn+y7/LEC8rJ8Slflz5PD99xtO/GuZ1ITgY8uEPpXJ2M33ocT4D
0tjTyWvFunun35uyclXOf31/LczevOB+mAly+N1xX+umI0M8IfQCVhDeOwTL76dU
nqsvda5bClfuBqe0OkH33A+WQxQ76gLvUWGM8o3hgkx0jaVn4CKIJIALVavpiETX
9yge4dUNDEm8TEI7EcxPL8kewYTVJoO4kZI9zbjL4Q/WNqEOgoTkSBdzgGLeRWlB
Qn0EJ+vS+CK21KTLH2oRPlAjRZCxPcj+Nz4RBDPh2zKXPTHXD0PRLpVm51O1MZ/B
bA0Etecuuw1QhrRPGiqPbCzc8KBgS6c+wasMR51rFMBgf8J7CM3B/Intly9Eu79P
W2Tdb0pkTxJQ4rGQiKl7svPEdQ19OqjdkyIts34Dc8mE5AJRyAoWd6etmo2QkiIA
0DCUsvl6TmJLY5WFzHRXKJKyI69mmg7FL2O5Yb6z8ra1gmJmhHmAQKP3QXyl8Vwg
+Y3REC0L4BBki2lV6jcOLkHQk+2A6ZnpdCcXDSpNCpybO/2c16P7hOx1mzUojJRW
ylXT+3xK/vVuGMUmoGMAASizuVIkjlSx+W6mFfACSTO7Jr/lIY15mO++AyhC8ea/
V7cWYId7WkUeeH+KN0cYBd0ZGANG7RJs+TihdaQGJ4snCGhlUprpy899gxVcUvC/
730j4xhvSfmbN+YUvr4fUe4k9NZ+KiDE9a+L+kHb//akOkOVypu1xNxX23ke2POU
balbW/SGxEs7oLu7SEp+sObFu1TCdHb5QSo4iVm/JoUh78S2Ni8Twn0oN+061mu+
wKEEGlUWU2m8Pkp1b8teDj1f8rEpT6AI93pn6HpN2wSkOfwiOIzE407C4lcYP5x7
XnRME0yxclJBz4+4DezKbSUO7lSU8JyeXr+tPQ7HrIOLwaG4r5ax5sVhfwodP5Da
z78oLPmZYgc9CUQk4zCicUs4t1m5F5b86J8LLJGMd7dd4I6nf3azwA0TSaKbv9is
0BU+wd12ebjpIH/k/cf3zJrz2mfvQu0TFS+0RyQbQkjO0/85JMk0fjEMrX+ECXrz
+0gIl/J6J5ihcgJlRWOvQu5cgFa2rJ9aREdoH/hQYKwEFaZPOjN/2SEgjG70QlY5
O+8FOxuRrpwquhiIRt6YTtzELoIMquabFFG8wqGn+LT9SWvM4u8cpkiZfRnQYQss
tbhS2jH0nLbewG1OIZQfPSCc2RXHF6NcmzQ9eAXqAa+R6sp5HIYxgrDb13cn4oeb
ZP2okjJ05BH0Kjm204+Zeh3cf1LQq/zvMhI/QCNZFICfWARj1JK9zE8HqzJm0y8p
YmEJmTOVnWEanx7SDB/8I0BENjPxd89efjdfyF6unqTERNbJWTLcw5Zcjm2nmCCk
e0fg6ozBJ21/UakWHpfCJXux1hQV6UHE7p96ZSbD33zP7mIm+pJGaraFbUxVPMJl
kragimkNdcrUVExUfHrNgL10r1P9wgrFwbwGE15CtOJm+Cs1FoOP9sbNzXJI/3RY
f4elxONdP3Ofiy/x/UO8WsI0jAjm/dkhdRjHJEYaU1U/462U7XlFzstqqBRvC9/q
v69Wng6kqTjyerg6yaYxuHo5Xu4tx46/fxirqfp1dx2OZDEgpNuDRfGrrCgvXMmH
VYjueN31avtj9p7tynFToFStpuPKfPWt7qCwEATFVq64Jl5Bq+zDDwuo4AyJ98tf
RNS4Wwb5334Q+LovK6p8MYQo4JaOBbmUA5X0a4fAvQnrDQPXAhvwO/ExGk0xT0C3
Uyv5GhyJvYdMdYLK/TsRxf3tEBDjaQaryKYtQKaVm38jyieAhiXlbX8mnU4+FtKT
57Y1WYPUF4B85WXChjYb3iH1DCzGftGphHJvH9nOCMsjYrufblhsC/OcG64e0jAE
Fg57TCL1XIrI/vqHrr3iQTRlyA7gAVUnjYdOGRrbBgOPW7CAwXR4D1ERfD3j+Cem
U7330cjGBgxzPMAfF5ohob08RvgNYXlc2aYYt/5PrxxESR3QUuOyTYHlKdPzgOj7
8gTey+FnJ5kov5mHlg+TDOB9WzoKaLeDwS4bjs+1JNtjKZtDcUw/8w/SlajECbsO
PGiy5xVpxdWD7MjIiamWB8komFJmbhQBxkGmEFTpYbOuNJs5dXQw8vJkBXaGXqmO
EsemQK9WIqQMG+eX06K7RBeLEUkB2YLhY4qOZ+Ul0jK7jF1fzchnCwOxOJ6YkvSJ
jWiTy7Oyv+C93JjoOHLUWohbUNYzHyiBAmUoS/PBFMaHfWBsvxfMJ9EgvDUQiY2I
YbVSbz+Osf9zL9ARmjmYjVJtb/FxRoHwlrfij/CSfQTObC9kVSiFRg+IVL1V8l14
ACcM1DqDaz3ZiuGXMsO45WxL468GsXjVRFd7+ZHRDQu1vElYIruaVOekS+kM0VwD
P5yzWE/xj7TUcpMg4kzM5DzEFjRsHmUBRVP8VsOoaivJopflEY/uRAW8ZfvwORrv
zzUnL8ZKGLfkqYl4VsAh4EYdmjpcjA/TshV1MoC+RIJcOUWruKsXGdheAS2spw4N
uP9ZWkABK+o8aiYozOp8U9SapiRUufxthe379AWrv0TYPjNqX1A4CiVwRRsP8opr
02lyhx52i+2P51psLg2A9Y/F4MJzlSU1vP+3QWHl5VeRRsWDKSOYG2T5Mq+k7HqX
LRjZVOooN5V/loeOb6Kq1NJ9LF4UezD+Ixud9FT548FPwYN5MnAEg66AJBPTl8DP
JLa4n63sN8g2QnmqitM9BxTcmLZ25cpXXgDh/UxUDjgvwqP6d6ZMDmphrmupQxqA
hJ0F0iU4SBXyVuhwe2+mKJNz4HgSpIdESOyADmMcdnauU8+FeNNjoZHCwMCeu9lQ
zp86axH0VSxEqncbcOKUilr6eaTEiftccE8jfNYmjp24ZbnmmUSaJlcdGArkw45W
YpJLEP6kLpGC+ipZuXhGp8O4eCvsTRwHTRuWRVEBsmF61VUf6EkY1DdmsBqozBUt
jM1gybv8BHxLajZ2GOeY9fc43SqsTPfVu/5816L1F3NqAI4Ijd7RxioRiSo3G2Fi
79WxS63SvWh2ilsLEo/McQHi7YmaUygyMNGv1ob+yanPSsJCBEwFDNuFGGhDBbPF
N4btnQmVAlsiIXQzJPMH7a07ICdZM9XxdIlp9aZ8Taf8ilHi6F76pmxlteYOk/Kl
fgnZO8f6FHax7655NhkfYLOJO40Xg3qenN2Ax8KX9mNzBsUC1anggRCF1oMjGNQW
tTAyeWwsCRM+jtn8GeRRnj2RB7n0FtTeGsDi1lSlcft7BpjChSQvF6FwxC2kFHIm
ARyHi6ozfmVFaBNHm+geQn8yQqaimIq7aaygG2fzxWzKoFRU78Vz3RIhnouF6YEB
i5J86Rql79rKVIOF8RcszIRBN3IUD3lZa4nG0L9FI9YvMpC7yYdEVob11GtHNVU0
5LOTkz7tvTgNliM9bOUCroF0lg9dC0H6pBjc4UwQa7S1SAmcVdaSxO8UigO7rYkN
AXECk5aPZAwCzulsM8+3t+bSSagZlL9m61QL6u3ZFX1Hp84xbLigXXXsf5Jfkgi/
/8s/j7s/wruBgdAkfDbcyy4kOVQokCwCB6XZNrGWBmpYhFsDEEzZGx+PKs8Iv2XP
AZRr9PiI9fP1QhKhlnMATFkTN5v8zA/Hqvt5R1Op3DSUmu4tTh3/jP3CUq+3KATA
DauGmcws2diKZcAGvCaNbW/sHy/H4V9UKi6gwX0IPfLPKaMqY+vavxoRoJUew+Rz
XlOBHrFbu/prw2igEGjkliBKinfOnqOadCZgIcHwhak1SXG06z1AQzuL1t3p/nuO
sCwZA4D27YOF20z8U+096cM3QWp2nPsS/XrJ2laCAdjNNEEn9b3eyXfl4pVZ+5Qu
oSDG161c9s8hd1o93XLVnwOCsEVgblpYmEVX7T291Hg+adiPTLEWQdVqKfzZa8e8
/xMGDUCtflcdJQdu7xlJumyU1cnmsSM0AjmbiUCWDYqqmJktYzNAudWhDrwAF51J
/98kQUOx3t/k1A8pgs+tR0/8NWK5WSy8dn42uJxBgIsHocZPZHZuV7CpzCZEGOnt
nz5Rfl4e0+J0A3yi2tB+EPQxeKKMyRIn2kiYfTaUgU7g9RGl2FcuQJmOpEt2qqTj
CrOKR6okGwE7b8ta8gmUs/9VC7t4PNCv5SiFg3j5AbJhD6FnT/VOj+8XXaIwyz7S
9px6/62bpkB8NorGlvu9vvx1dtSyUBKuHhkpau7Z+A+5GCLmfBDl2qS500GVlJmv
Hpn6Pm7b7Ka43cY1UQY4oOjwG67qpgIZKucz7tIhz6kpVpLnsWsMiJgnw78EK8V/
YL9Bc+iJe1mh11QWocrYRM/h3D37qpayxAstG3wHy2TExHitUyIaqwfZQwBBlrbm
2VmDWpF6dHYgu8vjAJDuih5Tf039juuAwKmKzZWpBUb4j5fvbg42O1XHNL4WZW/d
2pAs+ohFui31XQBCTj7BAbhP00dDcRr33pK+UZ9mCuwBvZdi5u1iwJI7bF+B501d
NlMJNd/2zWaRjy/xC7Cl2YEddNJ+yyAxz4+k9jhuZUvGSNACyaidwkJkQd5k+H3i
8XIXp/jAtRv0HrmWfXgvS+PdiMcpx+Em1Fb4eyKt6662G0JToOro3fpw4KDJDrvb
noaDragH99qqfHq/zZvJCDi2gJyokf9q9QOwVmq1kNbA2IvKuVRhIdzp8e4gIWpx
YzTM0KbaVLYD0QSs2METYlCTje/bfREeqBE0zxUO8z+nH5QyfZ38lGeHmk0FmAzu
g8bJ0vRdvOwXGF77BDRK847cwMwH1VzzMg8lKyHgYlsnnTI1skL8/prF+CawUXTp
9ByPNnMdeGzGd0idne/kdUjTtkXtw0gX3WOGhFQh2b/wiP8rM5vN4rKzb6xYnxbs
1nyFX/TaigG29B/ITyLDKWq50EutzHvxCpkrlX3OgPsOQ96eplIQkNWWjSFG+qBK
aBvdOAdb7oYFHob0rERWPhHjcEgYWr8aIPVfK9EDXjutUSgbcnKASQ2ijJIf4CK7
hIVsbH2hyL7amYhanFhLty8Ko2/Wu2u559cWdV43TNFbBfCbR0tc+XR+dz2RG6Sh
Bhb02H8e6p7R75FeLcSSj8v1HZVmPI2fWd1DXAb0qz1dISpRYaj+FQfZviI0eKwB
R9Vaz87IFuSrv4giuXHueDdYkDFfMNpcKqgjd8e0QEbIbg0UwN1/ph8GANp53mSx
/WZy/a66khh/cZ90WoZjoD8A5sw2W3l0oDi5rxMM+nXNSgB/qSYoVYfRSVB9OeMm
50UDKY5nqv3/X/HnvuKW3KL0FZumqk1B9DzrOsUJLgfVFg2AtM00wA9ijGYfRFBi
VpxYrkTTVh5FNO+CVen6TqUSUdqw/tDZXaCOpVMtt55696YCXV8c+BzGICsD0IWa
TcZ62cxUYfPlmev1neHmqpML+HBUwx/+R3YYrpIeZ7zFc5jI7eFoHjePBNcTyA3M
iNt+WDTUe2dd/+b6gsqzo5KemwTc/fxNQ2mOLlenO9lZRHMoZNkcqNmGl22eI/Vq
NrZkbSUEnv4gukMLklKlTeDl0wvXm8+91t3nlR0kfnUiuHRI+RihHCJ6ngpXM1Yl
Me3y9675GkQz8MSHbtmMNDjNRLYtZ4Yrvk/jBbi+iF0hk9QL0Jyw2HCIcTxXEWRQ
JE8NC3MX1i5myyh/7BGO0LLr2Hmb80tFyLlMAtQzTB3uoldxrIw6QtYm784jm+dW
7BONUL9KyQx7PzvR5mfLYMfSCJayI7OIzf7u/NZOge8LQSZU8nVvcrtgRkoTzWVE
4hfCJXcgXjG4qPsQccwWGBc1YP+QCOL1ORKgEqGP7dy/GzPqoUYlEbl+SO7MSt3J
HHTGsx+0Q2l/IFcx/Akvx//pcyveDnI6g+rDO6wXbNiEmI2cjKmHVmYfMJ3obbj3
xoFO6D5r+QzCl1hu1yFBiGG7SOWeKigTVgXYfRkGBKvaVt7BFLrqJNJN/cS0W7LD
dXOSz7MwSO9ZEnXleAhfATAsmy/cVb0swR0QNzhtVEuYhYLk6oBz7rz7h2F1gQD/
2oSg7ttXgHJpVWF9VW+rEfJsXLrHLCW2ewS+366N0ya+QemYkSCCaTazwHZ9qQzg
hBSoIkqNp8/lk5khst+FkwZdNz4NpVzpl1O9GOYF8hAnnKlW4Wo6uiz+nagp3j80
UtdXqj5M+FmKwzSGJUVIYCY8ypKPgfhLrcll9lxg4bprdeSvf43ccNt+unoAjQqR
tMHIhTPOokcoyvHPTqGqjFcisqq67+Zuiw+autAgsnPiuJr49JaVjRyzlZiN9c0s
s8qr8zJJGGAIolr4dr/DGNAqrhDGfHDZCOxGGw3621u9zggRI0AZD3e6fgW8frAB
+QNC4JQNQK2k87kcrh/0KzTFG8ceg+XNoucklIk3fVSSQW/d/yF44lulV7TcTyFY
9KR1lJdMkQ4Bt6awujKyrETGkmBdafU1Pv/ij+B57uuE+SPL0WhU6cCvu85yvY/t
utawhvC4t8wzoIHz7lSd3nqKLrm47T546Uvo/iVsTIHCISB7EvNaOQJvUjKYfK7K
rUSuudzMY/o8LV07WNQtTrUO9hFwrcWQ3bEuJ3XGoJruF7NO0sjNuHxyBNybmyAq
RW+NDVC6v5Wc/gFxkU3KPMPkTbnjKrOMLqnUdNHVM+15SO8B/WFRBJLgvEk+FOvG
omoe5K2ur1+nLmbMVMo1CBZLQc7yQsIlM0Oy9g1TTLYuSKnTnCk8kkkB5X9mstud
YOFAzbrPEPa04X+/BB445DOYmXLKkqIEU6mx205N9PwLHOSpa2X/pgQvWL6jrEHY
oqdC3v9FcQLjc8KiKI5Psa/QizsFkRRc2dxtkOFt4A4mQX2zvAvG3/CYlTfTmhZV
98ypJQe1qr2DEOyWFhUeiHKJ18Fy1JS0ulyDdczDgBihNnnlAxTufPjo470c9fJd
9n9I2ZWcVm4vTUCKtLaERV47i6ntkKXacqIzAygNnSjO938/XL9iLur+rMhxZA1h
AhH+eFAouOTNkHld5w2CAm3pWPuwJJZsYIccICVECPRO5+OIL9jVSd9ddyfYid9N
ke3Co5+jCcVZcvBnd0/j1XhNCc0V6uARRU7RiebAGBem1FnOEHhqFW1L9Bb9wB4V
VHXOS8QHnztvRrAeeD1+ruglqmxSsdqFz0KoC+8XdjqP5msRKN3Pm59FyNvkJH6e
uSrkmLY+QclzxYq/6nK+qNmD/wV0j0jWap1pAhrifvSr5PXjzJhi60rntOabHpgv
rF5u9EhupsbsrwmqWXykdQdPCZsBMFJj7sIa+YUS/A7x7TM3t3hFoYkH1z0Fp1tY
+WU0u5Nh+wlmB/zMeF+BsIQrBGGoaBFoGVsDKbGe3yWLUcSCW0H51pLe3ryZWsUu
DXKVp5XH1bzTtEKXwvBCJt5aeSRoHepmna90x+YailuUWlrHNBXBymVy6R/5IR8F
R4o4peAeJmjHGFGiv8jJHbtf5XDlVy2XXH7DjN5Nl5YrZntXlKg7deYt3YqsE+OM
2NevBtlOJOxp+vNFG8yx/eTMjN90JJQ8NwywvnoR7i7iRBbIahwUypkOjaq9XlG2
iA771nahaKF6Wv/URahlHv+RoNoGt/YrIKrHQQr4RWsZd7QaFCx2GESGtfbwTy7d
Sr45uX1RB95LCi4E8BPgO8e1fw+rH6T+hcWS6L3KsiAWaOJ6BEZSSOszqRn2wTeu
aGAXb1H7/xErPp9P3zS5W9eo2QUN+43CwSTWk1weD+8rbP+5WHRjBQGaxRE7sLbJ
/2QkB10ra55wayWb9pAzaMAT89bjEI1XzLfZ0A0O4LgXZvv2/RkcBQ8ciIC4jHDM
IHjzaTjBEUmDC2glIsDwcay/Wus5gxgbmD9/TUOglLnItLIGjQE0s8rp76TlANpO
eZl9ZZem5yzPppzeHQaYsy1X59rPPaYBTngE9WwF8Zx/dTt3kfrYK/nE73vMyrfW
bfX25CCN+8PRCoXc44ZD5vqzMX9Jle6p6SwznsYpAltY8eUMSJtJj4UIOlQM18CM
8m2PSnUgF6PrCpop+j/C+PHD63pfhVLkloxdHqdx6iKqFqRI4TDgNBv31LFix0gN
XSgHFhOhwG4LeNQZV16jESEIN2dd8/GlovNr6B1I/nNAIRP6FatDVPy65QLVXkwp
Sn1dv31RNAi5t9eZF3E6IrD2oXeh6NmlTRRFNTc8pd9/w5ftYiI32xlS9F+5A40a
rWTaEXbHPfHrC924ls0qhtywMVfNw5CVBp8h8fUYGMMbFD9gCZdvqCE1i88ilgvQ
PMs+58QiPon8xEGAnucLNdJVQiAlf9Zf1Y57uCfjkDe2ervuNf2xe+FaXnamYf53
Mcb+rI/AA7z9LvUybHKf2g4VRGIHVoZ4RZuKZZftXEhyjW4fLABUeOwTVmAbuTR8
XjClUHkmnjCupvl4Ncffk2ekeeUEsIiY/GhGtq5BHH8x2Ti+4Fe/AITT8LTvD+e0
EMGWoU9fbrHKsOrdcWzxRZyjdliTfHvoUow5KNx2xuLwMicHIbnZZcFMwpy8FEbR
Xyz6UeyYXqiQo7eeeDHaePZ0tP9QhnHVSpyMYRFsoRysD/uerm2nv938O79tIk8a
rPXgnpzKf1uab/HcbMDLpy9UK4gVanVP2P554FMJAxWT0aQbwWBqqT4iFXQ3xkxj
NcPpJ1XIWRm34/paOXgE7/3dGu098gMspzJ1m6zY3DpJKCGMwr4r7Sik7/otkbMU
4sEyriq0P5mv+2zZ6yxo4UP0RHxRwuN4GWDmwnFqom+pZH79rMvbqgQm2oy7tSnW
UOJ4/HfB1lxE8B1iSohz/Y86EF3mVCBei5y4XGqCH6YcnIBwoRM1O2GNoNKmVghs
+oT2fTXVPYZ9bM/L99CeRJBPhMmqGry8/beNFsr+hkwD8v7dTpxCUUuUJKXKrDzc
GvnaX2VyVOWd7khHh70H526wBogX2u5iJ5ZGwHwLj9gJ20vszMrKhqhV359/ZsQD
UecLPx8RqYYuptBgrKDyNyu3oYXyVNhMZfR6TVjgTW/ExFrM6SExOPXQ68NQwYLJ
/NGBJ3uGnfJY+bB+D5EEqPudCob6V3UoaCN2b2QJDCqxAI4ag/NjmeVyWmip/HTf
XoakQpfqbkuWlgVvcXTyZbTExP4t6W7pFzwwFed5abpubc+2+RsmGIDsIuKq8MKO
GemrcAacbst80IH6J0cagoR3Pr1zLa1wHocwU7nhQOhYhJLoSBFoLTN4r6UAIKdz
uzfoiWo84SxfafarwYAG6nK5na/p69vwbcH2WOZpyc7Wnj7yS7g7lV8Aege1/dnZ
pKEnAjVkD/CB2gwrcVlJ34D4ttnZr/69SC6wzdGAHR+00/W4XV4VeUhcFExVo4L4
VOQsgAfDxz+UZ2+rDZjAH5QE8vgC4Gdc6ZzHHE9Qlv0qvB6TANPGeyHT/pLwPdYM
ypW2cmEDaKAmbbjTOWDTNAN+uOcHXK1mCnGubvyR+JEeFSIaKcx16180SKY4EpXN
fdVsspVW4H44e0dFMjHlG0sScswIJjox/8Q0nwAYr53jLcSm5TuOy6cj7XgKYxEo
bR5hLas0NjBN8BPvK8A1kHBOCtKIslG5iEJ9lf0Mk1ElN+A0SkXvOIjNNny1r9NH
oclo5+ViYnnJkUDYU/cSZP4HyIl9fn4zXuLEmx97MYaTBOPask3ixtFChhrh0Fdq
3q74Wzf0yDiI9OWZN4pYY46ctv9nuOEEO+wqD2Xy+mzZxxKbOGUSbWIIQTN0cjj+
J9wvZ7nQCV7cuRuUQR/hXEQCiN7GtJ9FG9z4tBtgMZia76FRRGX/whvQR4HMIKfG
zKi2aTV3Bcefp8doChCQtfNOwTw9HAC2L0BEkmFMfrQqog3rMd0psHJiGv3kotsQ
zmMve22DlRj+4HQznrhIAxtZkfxbz+YnfzpLEHA7X5BMAs3+Q14/FUCc7uArsn/o
JWNGtysLPGHLRTvykNMkbnGAHUK8d4PfbwXbeL59ucRrbsu66ZnsuG9nP9VXtrWr
qj7JKLEnSBw+VQ8AUNf+cYgroy11RY2Y+okZVfrQeMvoHsl59MBkmLAfTHSlEZdN
kB+CuqZMFGsv6lue7BexjQQ7Bx8psx9vojhHgGWB3L5bviyadpQV24kqv8yHL8tV
rHXOZS5OzRhNfo/p0hZgZNIiemfOQB6Pbuaw+xL05jnhpDAmaHhERr2O9rH0qz56
eXEiwvdLqZMG/ytLs1URsbaA+L/5RKPHYDo0S3GI4vhodO0YPk6+uASUiDNFQqll
uGpNil9BDc+pdcpRHZiAuzUlxog/kcHM7d8JdbZPas9I7q1tirK73pb2f3G+aeeb
wTun7+gOSD4wBpVLOmIxCB/RN8bvC4qYL22Vmq6XBGxmzEN3y4J/+TOOT9HAfi55
ia930FQUT7wIB/fARhm22N7I1iqHlr+QcSXIRCI6zGgJy0N7PkQDuK50ZwpjwPEb
nZ4qwFAJc8yXQ4Bnx97XYeNG2gZ3/IPRs5d1v9kGwuBnb5CQoJe1fB1adsWX123n
kqC6tdUg1BRB7J8mvOUqgW6WM4aONe81sEff8ZIUqlFyRh2vBljhEsdRUOMcyIFg
ZnUjXukKQ/ofW5XCH5cBMqkYn9UlnG1/8e5xtwsQuO5Wcp9KGdyWR8EUf0sXKHFo
9JIoZbCPogS23hh7MTZtNorm/3AJ+e5uUUbOWBOqGW3bSAAJIbAtlp3CbenM0IYY
cY4d6HLvigei589Bja9kapS2CGgOl34tXSYikAQe9O5a3b1V1saJkWeMnKrKckVQ
LgNonOxF/zHSfp1Wl4gAudQ6TS64uLBn9UgbEwsacS2jBiOjebFA8MGgpdb4jfXS
sOMP+2wPvMxaLbNpZUIiDt82goDJgct1CX3Uyr2TLuNDb1qV7hgBxZUU4jXJoZIx
RxbxfYdkOU8Uh/G5ewG8T0SZofnxYIkZ9JsnJZyKLTePmQv5ZyJ1hoH6edKgeidh
3a5/b5zvuIYCpac6366tby/g5j6zX5CR8pfIItfvAS6Rs2hPZgpX749X08q1aAXu
f2n8BAPu9A931GcWVGaXnLNwIXg/8O3tJYxddtH2coUsR6pKfwBEsPu+zRMJAIM3
/jglUTmmrD7rHXVug11NkHU1lbBPXQqB0aJohjjYpwiaeRJ5hMEMZpMAHSrOI9N3
0Opqdh9xo0jIDvYG8asypQoD4cdU+9JuCq9z/JogWawhDxSKOWMDJxsb+gR4+iBh
qSi5dxP0hNuPc4EPrpqDRu/DJyiI9mst0ZkHGpTTAs3tyGvdlElVjPk7OmYsNvAQ
4J88cyYcmXZx9dOnD3dpUMMBHAIPbOBxQILMtouxL8N5599eE6pXsM75RsWqd8v3
449xdHTr7mn1pRclDC4SVClv1Qfd0FeOdd61HvwAoBH4yB242IWY36yeF0gBk+Gg
WRMBWpMN1ur33G+CfNwdXaR62UxwJg/RggUrVOoOQG8WZdTLw7/fvoTOSreYe6iz
TSkk6CIr4F57Zq2Qg1qEFpESEv8AULIggPL9KDHkQLBZNFRL2cRGoblZOC7v+5ed
WvoQq1q9lutE80M2NT5PmcMvbDu6W0Nruip3NnLual3pshBNp4HIWlmUe20x7Wb9
N51tLL6FMjk0GGXSFzR0HETd3dgSZP5MnKTxfGi8NG5DvnNDZ3cMQ/c3kCxB7+U9
uowMb5ZgDgY5pVSRDZNbowOmMfn/y9ci/D8/aArf+ED33y/2zrY7RHLgDOmrNixX
Ze6y0WDsm2VqJvNHE1hR/DA31KfqvrTDXDrISLS0HImuvm1OSIckIm+AYCIVWgXm
cP/eo5DfnJwsxgtGpLa3sMCxL8IYfSapgDhznwrym7+LyojDLtJR59XpOpqArvLk
4L+CxORRhxPfdVQ6DdfghRkIj/QxBU3myxVTXu1CyB+Stvq0fe1tE4GrhzVQj5CC
TgDMX/cYLvY9RwqmcHC8zJ1sdWN8NPO8KdtrgBSEJZa43W4yUYzwm4HjTOicAKU2
SyCqvqwIpC+up/OP3fKLBAJRdA3anA4BdU8l/tKVuTDAyYtS7rzAP87l74a++Cwb
DIy5PweiRaHlT+PuSUMCEy7mQ3r6NojL15CwifMiBCiiuSYICw3XDNpMKmiMgatS
hcPnMSHYtrGjwq2iDkzIUuXdy8IRDn/L6Hs71p5wAlzhgZIxMaHGevvZusyNryVF
X75Womcp/jzvb5ti47qy7j59gxS9nSlPI0i6GVM+KIS/Lrlzhx/O9pWKR1kDK6si
SkLk/loH5xNP0DxWfpOgjkADvB8M/N9ofmWTtXV85TJzE7f1P00byYco8bM3SkMN
MgUXpIwxecdb2z9EMy5SBsmVsnW+nZD5MOwHWfwqADqzGwVjvpXqvShX+xMFqS15
jm1Xz6wGQzIq9NjdKejA+9X6wKmCfHrmsr30BKW2kAS/fvsdXvVn7KvxUCZhvLLn
DsdgUOJF9nkriV/S2lCbnS3CftlutX8kJlmVgq4xBfWtsVXbFUL4d37yFPkOZarz
14ENU6eaxG4a0l9FnLtw6MiwXjUHlCW6GveI09iL9q2L0+ZEV+ydQ8yq6Yt/yZYv
noCdEG8sw4l/RT6ngrLKzJu521wCJFxzwDHPISNalaO+4KxlyA72YnUXJs7irysd
ESejmo/zohwjLIWDIx8KMp4hsWXu4L6GIHiJF/OgRhNVow+h/62klGPsz0SwFa7I
7gQ1fibxaqn2tRwFr7qKFoRSN0yXmUbkeTkUD3AObXR4uzlUR37uvOpe8mRXxs1Z
JeSzYEKtetgSiqkLvD+RqAYsuPc5skIcTSODjyX4KkXOVccCccmTkaYXDOYsblYC
R03amwh1iU2uaU+BZPywOEhMH8munsVEGglU/PSS8DXHID0d5Ra+AA5gHaXSK9pc
eOXdrEUZTEFLwVjXzCUvanYAs8XlGCJ6bCluH+5h8E0fC+S18xSaOb2pLZFhOlNe
7nPLajO2nBMNkSuv+XXJnmD/iwZ8gGsluG99+Nctrw4PijS1rQh9Yf2h0TaoZIJg
4WvvUt0P22iov74DS0C1ZCsLVZeU+UhDbUydk5PB/pvvnIh0ZtErBm1Uijj+h0Ne
tsymX8ptx4KMQOgUWIVXi73XYBQZOBDYolLHJMleGvt2+l1u0eTbbUZKlbQ6sHln
Zu9FrenTOdY/yjHQ20sii9cT9AsoyjH2yciSF9WUss0w6D7PWkzrTEYqBc10/tZo
6XpQlHDsJ65vjnZwt6O+lz+txZQxtBN1I0NlMz5QgRwZ1IFs/3HbGdBLEy745OTw
J2xmagy3+1m6BekEtakI7T2VJFCzlvLWnbd5tLp0WEfssbUg7X1OLqx92NyiP6m/
lzf6CNSjuK0Ynrr0x2hzfvXukmvVW7W7PkJNSIek5ikr+Os8WTQmROR9pdVcbaU9
kWc35+FW+lXIKNVdZMBPXhFvZ2flRXteRA9tNt/m2VwpPy4qfv3LwezBh/aLHYVE
5QODUIv16OdHa6rouh/lvIu9KmrWyy6KIk3VkCDDUIwR6iJNz5l2MD/CjC16zEab
sGRgCrIYVCpqSI5VGAGZ2+PXRWwgsh8krkM7rPThC5K0aZMLbi3UaGE6G55n40Q4
tlvaFpcWfsOS/j0KIXiVib0j4ead9TqAWr9/i9CdmJbHkiwD0muD81qqViSv3aGL
ChkiVjSB0hFCRpT46MwRhPytc+4of8CL7WLERwcRWcE7/aOLqB+0XqrePIGtIr6E
8jHQVg5RBYctP8kb5WyXKeDG17g31RStqkxesOp6iO0YFe4BAprEPCkv30w8tI43
dOHs1G3+Fq77flZXnTRVROMLNCf1FuKsZydsGHAkPtVpmtscLCeTBmFvEQX384rn
l6DAOF6Q8WzhrQLzJcmn9KbwOfVc8VOAnisHoF1zI+ZNtfri9vylPIl40JsgjSU+
GV7VH5zMVg9yzbbLUScjzaAJZGqbotkO/8eV6PUsPuigM+k2UmlLSPRkuKTN2Z0e
ws++gX0WuQF8kTZf3ch87ACb53T3BfMTd0i7FT26Q+k7R2fryMryHG8WsSV4Fs9D
zmIwCnt7WRAOVFHrx2l9iXth7EHI0qkmQ04BJ6e/BJtGX/2wiDpRnJguwhD6xyeL
rll3F/clG4vBRqScSAbhxJ9fWxmZGixD8pOETIDBkfUCKvLk07ADGuUDYpqMKPaI
E+A0cTi6YvZ3OMkJZUUi0ZShmyxuJR0DqiJ77LP7I2egg/eHGKc1NJr56CjT+HQ3
2qoryxm/s3wXR3UiZjrXDSEUMxcBKA0pWd9s4ooqqA5CPLskDAUWjIIppUZ31rAh
eD6V8M7tN4JV0XQ6/UDligpLi+qhSf85HE4MNkhhIndsKBsDRou3nqhikc8ao42P
0aEWR2YiJ+0iq0ehD4HdjOE6gubz8W6PUZ1DrMUyJRcnMhYqQYuPWTVK0j6WuhAY
jANeviAVZkx45rQF++FwQyYkoLsr/ubQkrL8HYJr2U2ltCl33nE1KgWEAtde3cVF
oSUCfajdDxS9fVsAtWXHVnCaG4vvhXM0G5xd+F+9yV/tcpLTiEui7qtCwkKsdh5R
kNsWjZiIxFkCi3qBWspQ/3YVUinFA5JKZCuynv1SyuEiJqH4m21DY09aewIwFlXC
EcLtR8YMR99ggQqbGZ8VVEGBk7M0u92IXGNidfUmQ4xB3Dwu4qVp/qjRVf2nkajc
xbkp3lI2BvALP93ge7AxwbRde6+X7k023ciUXGA3Wlink7M7aBWc8QUaOeukhRc/
9cuI8FlSpG33YTWH+nZAFh8nqHHFEEysEGv1ze5nZYqIl8qM6hZm9twrI69ur8LS
/QyValyitUjNVJrVsnHdKxNW2t7S+SYMYGZPnChTfP3xUe9RGdND4UTDyeCYdHbJ
/mgBlwaDyyh18gRrwp/vmE3CNH/yK14q1SaXJTbdMZBNgQWJ2yWT3CbRurD1wvs+
qrCrrxmh69mZVjGc1DNpy7rMEa8iMDCgy/1a/8wRk0vrKILZ8C6LDD+D8Cb44/ro
ix0NLGg53aB2Gw8R3pbtmIPR3JiN1vNc+t0nxvC4HRSdUDejCjEr/ZKMDcBOO4ga
x6fH/kbLo2jIL+TpK103Pxt0cyclShXekWjdqAyT0JRFnFJ3aA4rtxl8FG5Mt399
ECI4k1BZ+kopab8HuuYS/r2XCTJrBB5LGJsn3JK9FcsXoiKKLIgGi5oIOCzVcbz9
mIJK4YaGTvG+HECqm0kYfD/w5GIqj1bxuoFnF9l0svtiow/1kAZFbYxp9L/K5f6U
ZgQ0qAiw/7sUoWUHh7gt+P0dQnbaj3kX9smORjcB4bQwMCE/f3dbMJo5ZgCo4ate
I56Wk0UvFdxlqus1khvY8/q/coXya2cSAj70M90Zyvpp3ROvAvCepB/cznLtzGJe
tKTUvVmWpPOqfY534YtyO4okmf45//y5mp6pnGCchZGXHEtXBbIxL6N4fcp6XQyV
ucjPD3Q619rRX0nxlDbteX+2OP3n6VoViwB8/R4bMBX1ipDy1ZfqYPS3YZS9X8Nx
qdqIVC1EANrnbF0/SoHA5jrIj94swYQ6HA6I4ztWdV/+QVTEd44bcBQUssVo18D2
FoWa85WndvoYd+1az5D0hbi4J1PzLodccyVcHzk3han4QBURpjrynCXIjxQJby+d
REtH7VKTIQHizey1p5dhN6acoRGkzXE6n2S4Xr1upKx1C5JTRnsb2XdlLKPXbYEc
fy5AvBBAwEIqlZ7DA0lCFWRgVdX47k+CzR/8TK4oJUTZmnJAFQodMCVVd37/Ayys
pvDIjIbh2OzDx9DIlCipir5JQh2ANA6tpNgMml9hf+zHWuZRilPl47wn2Vv/tt2w
XAAFK8+deJCUfHFiy+KQG7FBeLUT9TEJZ7B8Y4S2NbUqefe4mq0WRDvBpQTyYgLK
qw5cdMOuE7u9qLq9/90BkDh/e59BNWe2IMerp5tJuPvjnyBa9P22JcLb625LuxSA
KJqZm0BUpTL0voEp/BzPQMY8/UT1Z7+bH9VRaps+GRV6XZPu7SBWfotJH+3eQijx
YiBnOx3C9wlv+1GQdsRqa8V9if1b9VpSNyqzBdrwkr/U4in/ig4yjz7kGg3o3eTp
H9MWZsNPf7SPfirppwoIDvchcuIN/8Rt7iz/wTnXwabQYXJO5gO8UnxaeOop77fc
MozH1w+tXk3g7rDX5AD/qMy3oHGJCtIpydOVxklCgwtyU1L5MiGf6489lLNbU9YV
92hXqDnrBmHJ40gWktp63br2592gCFO6QE1KlNiI2OSVE/qGF4zrfQuFS9aFkoWw
/wuJXSZ4sOSxAPWFEfgNyGd7BGKBk/cRCccheQXI665td8ww6ESFggIA78C9Dwsp
hZPgFVqYw2CTd8qRtNtmnXj56XVMlDOzKZfUP1oKfxogyOvJfxwCBESJ+xWnTtoE
tiNxnzkdg+QusJaypAtHPazGLsAlfkUa4dacPyfa+KUKRq52MgK/6gHkNy22nJga
LgFy270haK3hiOb8izwbtVw7dWzGOwRw+EzwRMLIhGCwtbZAQ1C3vQVpJb85XAmR
BwLvL/b8JpL5hMzMgREegDc5Fx0AJQujGOfMw1paA8eXyLdcnqjV4QgIYblZcC5p
0ByGCMDH/jz9ssy6qPcjemUAsDnhaos01YG63Kaj2aEdbAWEC1QjyNtTh1f4CVO6
46+NbINPliFD2bC+5qlXhzTSuzqI4ri/wqDi+X3sfjTCijnMPGy1zuyzdR5gucvG
nKrKm1w8Td8AW5K5PHi7TObPjzDlVFRZRKxmYuFfC1DWz8zP9EKmMYkzal8etMM+
MfQj8G3mAMD9R+k02Ht97MWMuLW7IlCSNHu18RNPcHkEy37HHza1L1tBedW8mnDw
swbHkGgKhURFAyAKcgR4wHE1vPrbZ3KIzeRW/YRB67z57BC5E1F/YJw9kwZ7nOfX
PS6D67Rl+0wEEMCQCA2SnQQByMHgf4tKx/o6EzN4vWiyz1X6MOqDOUnzwOSO3VbS
msTPJjtg18/t2O39+xlFAMKGCWCx49Ue4SvVlSzQuV/EEsAbeR7yUHI04KMw523f
ct5KXnGNX41Nmcrw32bOm6ELzeAOnTc3j49PIzQO7Nv3Qnoo6vzdRWR2dWO954aJ
E9ytTlE6nf6jeK3dAadtC0VC3lt1cQfv4ukrG8dtVH4FPAPKg57HT6Ync9N9gWKg
JY81FmRzWKUQIYC+FwLXHdv7B1t9W6nwSMOL6hbvwXP3S0vpeBukSLBoGsRGWMSI
uB6om74iIZJy+AGT2FeF0fknbmTNDfh3XGv87HctjyfVam0UakQpZB/DHAihPggo
8PiYJXoCXUwzmegaQPp7Wa8YcNJ2qyZvBZsrl/yS+8iM5Z3UtrSKfnSHfC9BBSaz
Lp0ZeMcvOX8KiwaJM0KggRpv6plQCUbhFLWSRiSGXS/rHoKT1+EfWYE8ZYt6CS+x
92q0NHP2qjwFrI0fy2+NnlM3I6lONCnEBKyDpruKdbQbYgte4lYD+YWJKR+8MuzF
kJ0wgVWuNUBLxBvSulfqrWu3nrcC8rTw0WWGQXYCvTCxc4FBdKPtQlJnvH6svjOa
JxTUAFKrazXC37HPaTMNXK9bVUle8+XJnHpYN3CJNc4jwUmGNnuUl50gcJiCsypK
bHETA2w8Csfaz8sTBlRPROJlEzN2IOUtdMPrqSdewYZjv0+vM1DdsgQAHL+CnZgR
E+qKq3eyqN4XEZOSenU+30DoTYUrYsvRCUjspjnPKbS3zIHILhNAfaiRvBrhzLCD
zwr1KWvnJmzLcNZLyXT7yd6VYrK1EAiKebMeyiBNenHGZXTQT2orEzyWcYjHrevg
0e5BXLCUGKRd4ESyFPYbY8kFT6lNXTD9+6x90irvmKlH/x9IiH6lbUYK5I0w4Qk6
EpTo1hzM7LCEJ2yJqncyEqQbXpAvJO5PJS6we+VtoskTdVJZh2t0TS/tHrot1FNh
NxD/6J8+oLIYTZftwXdaxD6PlziP2sfI5r0O7L5LceEGR4EAC5rMbyzfKSJ+Rx92
E+RXODZqK2ehW9QqZiw1/BDaCtP3K4YYY7CPm+GSdKVSDrRVXEahkERyAV5HUFPI
/ZqyNNDHSM54zPv1ALB/LwXoDHI+9PtWRhlh8TzfVCfVvwJoudGkCBH8GIWOUcgT
2erBYM51Gad+IBNtr8nXYxnTKdRCjU4HpSO9+R1HzPuzNE5LkyPPBDUPCAZF8FfC
s6zxBEdy3YwO/KpbEeK2wTiDSRt0y75h4kOtDAu5pQYHBlw1x/0/FBnZeVdCGBa/
FTN1mMM+VDokKqpko0QkHnzGKeb6dEEj4N633a+G7uE6AEkGu9jRcrMJ57qV9uIs
Y7KsPsAPenbI56WHXnjz5qFsRCko02SRPcIdSSdlaxnEfMXjVtXlUrLN+QlVAtlf
LAwk3xiTUFYZDbdsiZ0XpS6mrBBWM5e3TCNITFSZlHpv+/MAEh/YnnpdqY17jRyz
qUhOE6LdyE7I8JH9Lf1puIaiCCsviTVVvokjwn9NmRNMTyIpU+P3S5Mt0bPqbQ6R
UwjGLjm2+mHuBry2Ai3iwZ+RGHMQcdHE6FD6z/yiizjnP9E8X7vo0Vxoyue+3896
GMqO0SxzzHAKZUaSpzNPvj10HR/GHkjiR5WK+8f6GA+ImLZUL2Gg0hkILvyHJTqa
+ZDAIzjAMkUQtckwBMnuRGRh0pdwUzw1zmrsbJaPaqeAzWNcypOZ4emZy2xcfeiQ
edIW9OfXVXhALouPVWnLWNv/NeGgnwSb8jQqrFaD3LdR20vROjUHN91oC44GJ6Qa
3NhzmYtk2+6XBxptVPgRrjcxp7dpBWcERRbnJiSqQMhyKH43JydNpmVs33bLtV1j
jQC8viIkBgBDxfHMhfMPu6fbYWaKNiQsicJGvav4SWP6OPL5Gfe9LwUMamSRm2cu
eRvVX8+Z7SVXpUYwmXoRMKmAqyKhg5yA0B77u7yaWltiW8SQAKmL5WCiXO7kXM63
WBEnb2YeRUyUtlk01We5X2WnreBZDTqA1FCWzok4voNN4NvmrCoCHMDr37qGGeSp
d0joyfTLnnZZBOo8hqFGRsEqAT9ZCbn6Xyc7Olc4NFIcQMMQwYzLqAeVd/k/zoLo
eZc3Yd/GszOHHfVIhzE+L1QfrCpaD2D6qU9jc+gYjTwLpnbufQimHVRbbUMOhcZK
H4EMGHefwesy7lWQ77wscUQSSqbv3XGtgJ30faWAgbysuuWnny1c6EnnkXRpzQeV
HXbMBnUWci+9MHzyeX+Ms4CYgTY+JsF2bn8CUGR9ko98Zo225bD0LT4kbxCDePz1
mM7nHzU8ePNCx5M2xdk/anJvxTEejo9JdfVxcqzCE0dcX/TRzuT6kXGm4cx1y+G+
Shm5hNkfM+/PBOKPNkTGm3oyVnUbwFAIYxnwcBhVIMCyqiU+nUZqzmcAQ3BPbV4f
An0GtNnfGtFvMJhy7cDUy2KnyG/8bg2SbD70kcNP4Q2Zj3JnP+6x1n7znv7C0YUE
9VQFi0MFwxW+DioKDu07biD4AJ8El3IONuBYQG0NO76XWaffG84fWZyE81h8W9AL
XZ0EdlOkAfUBxbwEcepAyv+HKTgMK2QMZmdL8vJdKNKagybs1dnQL/xnN5N8u9pZ
epdWvUb0C0G08hOTxNgG3VMu+6chrTso9rfKmnlbAj1OE8oNkUDNWoZz1PDRxE92
mjX7o3XqHHIamla1C8vbCTDX3kjLVJT+Dnl8JI5Pswt8DyDxoYUET4AGpYggVUTM
UDyi8BMEztmp0fZxZxf5UvTOXeo4JcOPsMVwn89lTClpSzd4jQTRWMiW4/D9/DS2
7u/kj8U618iV+dDa+Sxv6auamOhxIdsp7xQe0n+6aa98SNl4dnEg7VTEez/6LhmH
BgT+Vek4PauxobnLBZKUn1hYgAQc/CCX4L93S2hfnLdpsADLdsmqUm759jgAdoxs
LNuBceIZG6gcOEVekjJF/pNOQxc1WX3x693+1oRscIqmk31dIRfJ2XbYT36yfC5D
UqHnDyRbihKNc80DF2tErIhJuBOnBBsWwhr60rUlE1ace1TWDp786GZzCPwPYrgF
SCtsuFuu1/mMl6v59RksfLkyhZ8Nrl/kwaptwMDvWws4hOxZaeEjg6TjaFADkfc6
4Q5lppKkxqQwTud0sSIzI2d0lzHf3pB1SC5SOqDM1bMp7fdPLwelcTpI/2jardj+
GP55XNeuP3IrAepv+ThM0pQIeP1YvySzSHunDRAmuvb/2t/2o+9RnvAeqiPj43eP
i4djCM1jnuE2qJhPPb2cDdVhKRyUCuHLyyGAOaHgnMljBtnU9mxuLu6RNeAZ4XmX
Z7t/p8kDvZr0WyWgHXtTOV46qzANMU3m/fOIF/BPjaghTZ63RxxfJhgEs37IV2CM
98ojUzRQ6MTtjcKt6m7L0XYJgkmIqVK0cmjFltOGfSD3rUZM6MkS4tGl+i+O2FHD
itVQYeZ2HCqyr387qksOzRRd3Y6dcv9kBioESCt/NidMOXAyon2ggdfpMXRuxhyO
RvNHaxLinkIc3j80NA+da85OPcGaarpM++RzzpBBJc86dXYYWM1BunayAa2JTxhu
xuQnRJqkjODKPKp0doWwp8tYjFbWAI0CcbBEURvp7JyymO+YnZXS57OX3YelTWN4
TrUYDcnq3kHJaWRpmyQNauK5PKeh6HDJbg/YTDxe4YFkmfUV8cxuqSygQe4IQswb
iTLJvadVbgutAZ1yg+rZAZypIUj3l5GOkJGjwd6xqGz0zfzMJcMs7TujS3njn9Pq
+51VZ27ga1Un9qCls+sTVFSw2k1JDfm8AjWt8KBzGVHfELARQ28V/wEUjZonT3aL
BVOnprPUdXYbwVE7a59ebignWwClvEkhK5eovTG5ULCcWkoEclNzJ94jkRn7NeR3
FPG/Dv9QTJoqs/MCi54cAFntEUeVxI38b0DLxerjfsydrqNC3jGsak5xY0UzM8Cy
ZZhDsZTeWdFe1zJ31GXv+abKIJN5KqGJBD8i0d3VAzM5j5LFz+nw8SkDgHmIuXcf
+jbmy+tEgDDo5h8/+3+cQHk2y28scsBThMC8HqfJO9K0wyneu4tGuMLyw1XzWxV+
BZHTbFZZVHxt5hTklkw1fD4F61HPIHm6/93riYahj83ebdc3cQFVJUKL0J8Q/ZmP
e2u+HrFb30i+90jW/FipMvTY/j/S2v8iBb8Q4lDZYubzqnXOvud+bfF4GYhHNl1N
KTUzL8tTahr/9ueO87WL2f8dlM7x+rkUp5UXxFDt3BwrSG+3Z5dmQS9T2hKkXbYR
56iUM4GbId3Sc5PiQFFVGtDas/86bs9ZjoyX3GWAgXtUZBWr/usDJ69vn6RNs/8k
jO3TX89DJzauUm57f2dZsr3zSuYy40plGMz4/s9OxwLxbzu4vz6rJg3VegTf5Nh6
ccT+o2xlccDs+NIqJ+DLvFTZZfpOw82jL7Mw2uPcvXSaiLyUUBssn6EMRMYidcXI
CXMRA4qAp8N7TlHavGFaDjtuKptiY8RfIwee8PelWiH7SvCWNzve3+z7PpBftCPn
bWKeSuqEH3gQAjrD/oeuectycowPVGfNeJNvlDjXZWQMNr1jUdekpR0tOSrCChjO
BJaXQyI+WKa95LkPwRS5GJswyvZ3hlmE0LWozIirAB84RMdqgNuBTEF144BNZ6Ri
L0t8e9JNZbJeGsjTy7lMbcuoyKPqjL8WzUgdzYWwTqU+Bsq2pRdY/Tm1Vp3YdGqf
wC2fVBGZqqmBCbK4bwyXn0VXu3a34oEQ/HcRUxw+nQSZyENcnLPS3jY98GImDRvq
AzKa1HHSfTf8YR2NSYf6JmLUjBZUg5QxFLDknFMsOJA+zpLkhI2lyrNG4gHy/w3t
l+7eKj+pCnvCV7DdURq92WP5SRPtcAQpRXOMGp/t2a7edUkBOZmaQqaFJoJIXsXb
CLM3sleJTME77dDwGtijep77/0KvNjrTy5nXKJKeTkMA21u5gipbRWiR2avwUwrb
GyMJawZeYhDMnI0fa/nNfNexHPw9UZEiPTfHH4NFZB4Zt1+ABlgSU6jElRAYq6Cl
hmiJnpk3cXR2GhTknPG5b2c1RM6LKt8tbNfsQU/j+2Z6TG8WUbzDGBBIeMuwvv1o
cEFdGiE4PmG/pCSqn1wr4/iXKjMV9wjQiRUYbNlHxI24uhjbIzKfmhA53yO/WWBg
/BMet9m7ZV3l198/jUx8N2Zlmls1aJW4QJaANhurwHBKd9AnKxMLU6uoAyIjTnj6
UuNX07bw7BIiwF/mv+7Oro3d5VHIg8zp5ecj5NBHtBj9G0+XeEqnuWk2K0C4+4wd
JcuuYLgdjfHRBcJ5nSU6ffnFUfYJiljqTHceWPIh91v+p9ZYfgd+cGUaMN/1ncZM
ZdUvF1uyeJLRwxoSA/wuQo/H58q92YwZIiZkjn3Kf39gzLtZ7f6Yk2wYFB5feVza
/jxmp/Ay08SUjG4ff6JcC/Difn9Clmw+XAw1t0xMEB+wqki+LDHAvLQHRhs49lLn
dBP00gz9Ly91ho9iLZBa5IqEt0jiAGSxhhhUnPaBFuT427Rk2zYA5BTfAtfzOzNb
dl4YJSdd636k9udEOEwwSbIWP0M4YJfBsIPP/J22uLU3FoaMUtWTP65xf5XzH0AB
z8gMIOxrp7OHufVpjWc4j6xMb3V50DvRXP8/LTYwtDg9OIETalP163RZNi73s55I
fURBsPUJ+qtX2pfHqGSLluCClhesLhxTRmp0DbDc8PgPboOD/m8FTNYVi0QL2FIE
Zn3kkUYp017TDBhDUrt9TZUeiURoput8//Xvr+Zdl9TrMuqz5+0B1XddnyVEGh7w
UjfqlWwQXnBwj1ojgEYuLqBG1FrxOrdOvB2dJZSysZ/4RslRpGKfWibbhJYhZdsO
KfgphScHinf4KKTX2ZaIa/5hec+w+Wbv1P13+24FFXwHdHjGTdkUEQ75GDbGR2RY
p5OS35i7+ZKZrXI5oGrqvQQrWd2NPf9mwYqIkcfNOMIN4WHqRbDJmNtjbgwmN8vD
HUNHELk47WCrXfZgNpevrKTnipuBcRXAi8hQYIgegg3FwEwCLHGbum8f8u1b2UQY
JhaKB2gdp3JAgxzNe3my14UmvWzGl5Uh3WZ+iZE6LPUXeYiXje7j2asB54hXFTLI
plAL3VaZsTnqe2OWVtu/FfmRl4TnoXLD5FWOfpEOrZCBig2B9NgoZ34PCOWC/Ca2
HCMprXJjgzeN9UU1RL80QA7a1MQBfvY1MlsJ9WTkMFtGdXDwIHnh8rXMKeuSwlhi
WD2NsbxB/mtshll9Fu8chpA1pxGiMU3b7ukEqh8vMSZKMn+9EULbZmNZVyWy8HNi
bmW2ykTparCHZECxYT1BmJYK7DZF0wWUkGZ+rd0uIeyG6IMGyBLygc4Lu7Pc1pYO
3sLlYR1CjEZcUrHO05nIjw/2lMXnhN5IJqOZ2svdF7OgcuVMYGGD3RHvwXobr5D2
5DVEkGyeGGyUPT2p+KlFx13D671puAs7FO9fX3oCGyHZGfZmeB3h5alklkFNItox
ErGvMe2r1X7MiCrBVrtDcsUe8NZ7IkTMh7hvVNg/9n6Z9nWrKSp/JZs4AULoKtJi
yeTWykncghifZ5Mzi0sc2mwdmjvvQzWdnyZusMyllW83/nYh21Mx6aVdB+MpIpPC
TmXZuMYKbtK2yrY8gwGcB0r6vXXy9luNHOtGDBMNiXUSd86Y2ZEUvrxAHWn1HyV+
QAF/TGaOsF+eciV+KF09CLM9ToogEhuuWdF6OD+V4ogic1U7CJB+vQxRXU71BIcM
`pragma protect end_protected

`endif
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
YGwoO7ncUsCqhS4vLNlvATlsygBrygK0QibhGBDLrEjxdp8UZX8vGzU74OUvTazK
e5d7iJYeBY20ca1qd8EfMsWEOyMoVhqDtdpGiL7NoTATJ09srbXFZWAONAk0cojd
/trbyKR/rI2bjghZN20d9bGDqNGnJ5sJdE4/7Vi+718=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 86879     )
K084BW6nnH5nMVdXsW6c8DtiE+JGY0K0+ylmjbIJOwM/BO45JbCu+FwB2yatlPlD
HH0GCZpRqHw48mVkI0jlS6CtZLkiVzARCar/In6NZxS1ffoRDfoA5nEWp7k1xOpi
`pragma protect end_protected
