
`ifndef GUARD_SVT_AHB_SLAVE_AGENT_SV
  `define GUARD_SVT_AHB_SLAVE_AGENT_SV

// =============================================================================
/** The svt_ahb_slave_agent encapsulates sequencer, driver, and slave monitor.
 * The svt_ahb_slave_agent can be configured to operate in active mode and
 * passive mode. The user can provide AHB sequences to the sequencer. The
 * svt_ahb_slave_agent is configured using slave configuration
 * #svt_ahb_slave_configuration. The slave configuration should be provided to
 * the svt_ahb_slave_agent in the build phase of the test. In the slave agent,
 * the slave monitor samples the AHB port signals. When a new transaction is
 * detected, slave monitor provides a response request transaction to the slave
 * sequencer. The slave response sequence within the sequencer programs the
 * appropriate slave response. The updated response transaction is then
 * provided by the slave sequencer to the slave driver. The slave driver in
 * turn drives the response on the AHB bus.  The driver and slave monitor
 * components within svt_ahb_slave_agent call callback methods at various
 * phases of execution of the AHB transaction. After the AHB transaction on the
 * bus is complete, the completed sequence item is provided to the analysis
 * port of slave monitor in both active and passive mode, which can be used by
 * the testbench.
 */
class svt_ahb_slave_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_slave_if svt_ahb_slave_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB svt_ahb_slave virtual interface */
  svt_ahb_slave_vif vif;

  /** AHB Slave Driver */
  svt_ahb_slave driver;

  /** AHB Slave Monitor */
  svt_ahb_slave_monitor monitor; 

  /** AHB svt_ahb_slave Sequencer */
  svt_ahb_slave_sequencer sequencer;

  /** A reference to the slave memory set if the svt_ahb_slave_memory_sequence sequence is used */ 
  svt_mem ahb_slave_mem;

`ifdef SVT_UVM_TECHNOLOGY
 /** AMBA-PV blocking AHB response transaction socket interface */
  uvm_tlm_b_initiator_socket#(uvm_tlm_generic_payload) resp_socket;
`endif

  /** AXI External Slave Index */ 
  int ahb_external_port_id = -1;

  /** AXI External Slave Agent Configuration */ 
  svt_ahb_slave_configuration ahb_external_port_cfg; 

  /** Callback which implements transaction reporting and tracing */
  svt_ahb_slave_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

/** @cond PRIVATE */
  /** AHB slave transaction coverage callback handle*/
  svt_ahb_slave_monitor_def_cov_callback svt_ahb_slave_trans_cov_cb;
  
  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_slave_configuration cfg_snapshot;

  /** AHB Slave Monitor Callback Instance for System Checker */
  svt_ahb_slave_monitor_system_checker_callback system_checker_cb;
  
  /** AHB master Signal coverage callbacks */
  svt_ahb_slave_monitor_def_toggle_cov_callback#(virtual svt_ahb_slave_if.svt_ahb_monitor_modport) svt_ahb_slave_toggle_cov_cb;
  svt_ahb_slave_monitor_def_state_cov_callback#(virtual svt_ahb_slave_if.svt_ahb_monitor_modport)  svt_ahb_slave_state_cov_cb;

  /** Callback which implements XML generation for ahb slave for Protocol Analyzer */
  svt_ahb_slave_monitor_pa_writer_callback slave_xml_writer_cb;
  
  /** Writer used in callbacks to generate XML/FSDB output for pa */
  protected svt_xml_writer xml_writer = null;

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_ahb_slave_configuration cfg; 

  /** Address mapper for this slave component */
  local svt_ahb_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils_begin(svt_ahb_slave_agent)
  `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void build();
  `endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
  `endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for slave_if  
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
  `ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
  `elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
  `endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);
  /** @endcond */

  /** Puts the write transaction data to memory, if response type is OKAY */
  extern virtual task put_write_transaction_data_to_mem(svt_ahb_slave_transaction xact);

  /** Gets the read transactions data from memory.*/
  extern virtual task get_read_data_from_mem_to_transaction(svt_ahb_slave_transaction xact);

  /** 
   * Retruns the report on performance metrics as a string
   * @return A string with the performance report
   */
  extern function string get_performance_report();

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_ahb_mem_address_mapper get_mem_address_mapper();
/** @endcond */

  extern function svt_mem_backdoor_base get_mem_backdoor();
 
 /** 
   * Gets the name of this agent
   */
  extern function string get_requester_name();
 
  /**
   * Set the external port id and port configuration
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_ahb_slave_configuration port_cfg);

  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);

endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
xZrdaHmK2ZZCBNQ3fh6KOy/kPXjV2KVpUdeJ5++2WStu3Vr4ReF8sr55zodnjPSP
tfnU9OumZRYdPM07QXJHv4XsDAqB/O4I6LHyMvmGIWGb/BqzqL5SHeqIEG+X+t/X
h2oz+5bmqrVJl4aEKjgk0Z3YQORlo4iW0Ty27FU0qlzHmYSUWrHz9w==
//pragma protect end_key_block
//pragma protect digest_block
Iuz8q0XiBjVmKRg7Y4Oht8kgfy4=
//pragma protect end_digest_block
//pragma protect data_block
RjYWpMNoyhoK1OA0uHkreKN8y7WufahzTaINkeZYoULiOhTyXg+tMdH/mcLYOf61
YwXEBw6U6WO0lFGrDYChq0RIeqIVPWamaBi/w8fDmVDToCcnIpguiHSeWDGSYCyz
c6kM+NS5XWvACv0S1z9xpbDsn/wIcyjctQTHX21uo3GNVNFbsokDZ6IdnqY6CJZO
2qG2iHUrcmq6FQGQYnm0MLmqS21ATrwNBNsbH/ruVz9pIUqbhBvtENcLjRjFJoaQ
YY4p+MWbVBfhUTgMOscG5w9Y3uUM+gczqAgLomWaiqj9bvnkvQUtyce4odBW1jWf
fkUbBJyHQWOibrJzudYW68LlJAK768CKKU+rOwC2x5BRAmFGeSSF2FJK46FIB5Mh
xB06i6yQCfc5ZIHaj5yZ2yBgbQiXyxNLlaIKzmKCQaIqub2+5fHdPeY36JhFctC3
gOiJU+TNOp0kJQ7spIdZquT5n2vE6xcphDOQUYtjrVI5k5I6oocONl2+9qWqTbBP
eWxzEqXFI1UENuyrpstLRLNbPggekhtZ1azQySqOWe6yOjpLo72qC07fowH+WK6q
9k3IfMU1HeWD4SyqQIVxQZb55vyqHvl5/GghtESGVQv6a31hNtdZKXZfwmHlVyRR
97R6QjN9kwFO7s+sUPtLIgcB4n23nGGKAoiOjV6GgS8=
//pragma protect end_data_block
//pragma protect digest_block
8sEr/CLjOJIwILds9/yodApai7g=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0eihmmkRmkNpj5hL7NJtM3eC2SakZlKqNi7p7Q2NKr4ivNxymZa3o55Q7AUEMzBZ
knUmklGl28CsafKlIFZvhOCPb/UVycppw+uoBexK9xfWrS1hFIZ3xwflUwxHmOSW
KoDk4X+LPqPRow8xeIvmwBAV9fkLi8PBc2S62zb5KsYkRvybZwkTaw==
//pragma protect end_key_block
//pragma protect digest_block
YeV07rRlmnZ3OabSH65cGxFkdzE=
//pragma protect end_digest_block
//pragma protect data_block
J04GOos4gYezImuriOJXLwQtuumFyhxy4HfP7o20fy170ZeMYc7r6EH0I0dO7Ivx
9acmargoeZQquXyFbpyjUx8KlgsOS7morC1pIknA1nC4lf97aLlZNddsHzOoduPi
bY7pW6H3pMWMQjWGdRp12dCPqlp8X3M4XczoZhN9VqmG6+EnsV0yhybqJFrkhMS9
hhaRke+ewmKzASS5jeuDkGqlGP/imw8zHyZjL5OLuGxjdzKNZBGABXHAxk3ORVyJ
jpPh7P8PevzhdeKPK7qD8HAe3qEkxjAJZ3v+di/ix6cA1o3Du+J/bnF5o3wirXZT
/jad5YJwD4hEvkvS5TLV9HmbIe1FokE8lrLRTjW+SaZNSCruMS2q87FJV0ZB9RAx
LQ0ocUiht8gsccdQJlHyKDkDI8EcZdSxe2Zd6Apts9WAw2AkjUejWFCZowj+G0D6
bjyXJgxIbYyzsT5kdv64f7niBDvvQsdZtALqGaNO5afDvbF7j/Pwdj/+RHW8tWgI
VVL6FLhOjsoHkHDS1+ZFPt9RFPwn0hSGd4GvNniqa9RE2cGNTzbpve9lKX6M/l3S
x2b8G6YKr5LkcdgZxPt/oFPiqK1OboRWQ8arhJtLWXoqUoxk0aMT1k2RKVCrSWsu
+saeNHIM5y7DcJpIMcDNCuAq0Br8Z3jWCVohKOel3vz1FJ0JgTJOGrjefBeIpBpA
lKLQ709uCr1E4knmTCkcCpuflXneBnaPlmmUMioOBvIQywh4vL8Ao9dOw1lEHEWU
vzQ2tCwePW9fWbzPCQzk96gvIIUF34e9KCQPHZ7uX85TTVamgDNj7nXHe3u1MNcF
3kn+x7n/xGnfdjOf+1yuOlEmbO/+q3flPKOM5FhPlp9Uzt8QBp2Y6JjcJ4K8WP41
b3dfoh/40xCRxyWFVM5GX/TY4nQqwNDon8GuTzXD1/9VsdYw4kvV3h1UJkhjfsks
M/qIS+8/iPA9qB8wW+UxL5M3cNWQWmvNl816IlhpmtFTHr4jPbuv9CjwNSVkdmzD
ttIV96i7rZUBA0qLUF2HXwTiWlY5q8SEJPYuXYCOwuivOf+GnmN9+l6uXixniL1a
7c31U4TgCkCXk8hBTTNwuvwGNL1LpcmYLgaaOG74HN2iZisMSS1Vp5/MsOgLrzHI
kHkbkj6uerTcwWmpUBq3MJRgfaKUwgwULtWnnhO2p6xHQ1xAy8PEl1tVfT92Mjms
rRs2iavzgF3e/PGABlirwGODMpgNJsgth0aWexgFvfy91vpjRmDpD7N47Q8D97qo
ssuQQ7KG4ODdCuPImsIwV30gbaYtepYZ8YEGzb0qICI3iofOA5OWmMrWLgy9B7ws
0dtGny5zvS9evgg9Wh0E1mcdQ5FJeYMfIRHFNpuTI98slEAozJEexIZRLP0nWdm/
OZSp9/2Jeuuil07uDNaxgjpCr7DtFXG6ZTTCr5GVByKjakMDh4WfKXotXBjL63eg
BUaFMGvHDvVYbrl+E9D88sovO0FItqTntg+W4/bnusGYNwKtpiTfCWUW3nWwNbEs
PJcWa3wzlcFWsGDrw1Lmt90yrO/NBDKb+7jm+65zlAYUcdU7VL3akerKjAKDyhP9
ACNJNLCCn5ZHXvcctOFmqzCAyb9WIE6cRDWRwhnfkCzE0ROiK1pPkN5VCR+8kjLP
Y8+G8gShxkDqFcdCfU1JKfhHeCwnqb1oR+/dkYaP3CAd+uByumLUPoR9Zbt7krAd
RkUef68Udu3+skmrBe8SIVWmU9blalpNLlOk+jw41IRSoN/TtcdSUr4qHQ1zaCj5
eb0R+I9ru1HQp6smzaYyQe0bzUYDKht41WJdG2BcsW4VFwOkOVM2TGYVoFI5QK0z
o6N6QPiYvcv6J3fKJMJE1fd3GHkL5gh+lVwEK3H2cB/Fx4y1i8CLlRTchGZpYz3X
NTDIejUA2gukXw2RmRwNBHS5ZXjWnO2QrFZJPCIzsl9raQexTZDgB/NDhWGPwuNM
6FKHK+unsjFYXudT4eshabBSlDiqsndOUfVrMawhalCtle8WiO5bhikBy5VwecGF
PmiCp9ISYXx0lA+k7FW9mhMxqhQKvd1mKIezFWDjsf0kkpJUi4gYNsgKQcZuD0uy
83n1K+3lwwp3bxhTrZ6iJ89/5y9VIKi5BFDrYyR2CSVJQHzGZMCsmCW/Eoo6+4dE
2y5cEQJWfqLlmCwZLd/P0pfEGIxr0ZDFSjlbKN743ZF8Gm36wV/qXneuy9nbMKH9
cmv83bLtwmKd4kt1l6ibeyJNmzhggpueBzcYeyjLjHq41e87G4cP1Md8jnjMSNMZ
Ix5subItwSGjH1f2ZDJmBpk7iSBTviUlQSE1p9i81IxbQk/INXh5zluOLXUkqn3j
8HuTUUbIQBcCk/uLsr2y6CyZp7bTQoQAzQjCVl4ZhsbDd+N2MhyvN9FFS6vG+FTR
IlWYQFqleWzPLbrq6P+INrlFB6Ga8OC6DH/1AhvwXlQ5wez3cZVdBmWnyRX9iiso
g2HqvxT6TB0pmc5Y5IwaKL8yH5Svm/9cndhmLedEzXgp3RJkqckSioRUvpa2qpFp
quvelDMy3lFdtOhZTn44JsVm4nGPuxS+vXUH7FD/az5EXbQkN3fZEo9sgtEvUncc
BMo7KzoapMrTHw0knLgmGL6nwZ4awcRkmd8lbOtXWz9IHRP5Y0kyKdUNNx7uvkPE
YE/2X7/AoStnA1kQXdQqggvMH5twbM1tiGusVPBW3K46xpUkjmvTB3yD/rvjtxWV
yQWBOqPscDZBwsIiJqzU5+J7siZdycc85RUSrUZ25Ltz7LUD6F1GDPUrBW+ld2Qp
05KV/Pu8AH0SUuYCjgEV3Oad7Cuzu7PaipInIl7/9mwtnKstynkQg0lqWqYRqcHw
aMWYouwAiZaUF5gr0lTRp86J2AKUqE6CcPGq9nABGSAP2InioqAo25UIdzzLdp5c
EspT8xbNvgkpJdjj+zErjPCbb5A9bjJLm22DYDvJYt8yDkj77Yk7zXDl4/AwcW5m
7mUxagYN85/qyQf08m/NTZi0w8ZtzGUtr9Ul6cRpqyHIr7Ed2DXpkDXpakh1ALet
WNd98apAnVuyTKEU79mpSL729yd24IwYldAXwJRPWJeTl69rsiOrH6jP1tcsRxqx
84847ddY+cJUxjsFIllb07zxE1oTKsP+UHN4PApgklMRdUP8R2qvVj2xXgeg/WUK
oCZFpsgUoyryCwu/BYhZ3QlHq0tTrWRTkulJNSQ9EaoA5BfsKZRi2jYOeQR9D9v4
lUgOYew7OYkrS5k07Z+dKJBQ6+nfG/qrTPVq1zBLcB8KAKBe/GiO4OpccvmdRFNZ
0vlJBS5t5kc9eMFAad8U0PrGbWL4SbV+WiJLana0dQcz5mVIRi2VqcWtIYY97sKe
/IsaO34xoY0ialMvP4qGlVdOzZQOrFnkOKcfFKSbCARxcjE2PzAA/puy3bIpX78U
Xlbol38wMQqXOYOovnKh3b5+RQL92v435+ljCma+sAoqo1ko8wAztHJQQAOVVXZe
1jp3x8WoZ2bwgZSXVO0hYmItN69hdm2zhOJ7WDqTzAa1h/sw6syk0TDTf4JcYr/X
mMGaciUtrOXtCzXh8EulrrrY2UB2k/S7F4xLnDa/6xQAzH7NZx4aqRoH+Tx+LuX7
RgsZzVd0k2pJlNj+tfFLaQK/Y/JKuE6efY7aLeQBvZC8oEwv2dLuAUUIhwaezawZ
HZqp1pqlf/0fGB+OIXREaOrTjJKszbyPbxhGW+4RqWYjnMDKUNAWUGJBSOZOodjA
fBBcG81FlHr2T2sJxy5shl1NFr1zJy2+7C69OgA08we0Zf/MfHmvamzb4Mh2Ttmp
U3YhL1J7dWrkuoA/GBh3V3Lnz+zindyQ1xHzUCHWKD8rNmHI2n2IC4M+0Y6/otff
0jeC1DV8eo7rqSn8HIg6CGBcjDO+Wgj00xdTygJD1gIhEvKu78kYGYxED/5NcRlh
TH5ugllwNZ9JKji8tv5WDwD0ShpIVORDlwAw4BagL8GSUjYaaIwyInfQ6NJwzGFQ
6to1rUaY2+V6VoZemsvT5B+TFZuvhMf8YM6lnDwd44Qjw0jC/Sy8OvqdLhHBCBpI
m31xhvJvCEy4r1EWvHMX2Z+5Oxuu4rtlqPNBH4vUXxpqqyJ461QYwTVLGgFLixe+
i3tLOvkhJs3I39oa7Tb1sS+k7unfry3ovibPX4ZezBq3OWCWTywUcTnxUXBUXg8D
8qym3+Z++0av4BgMa1Do0uDU0LSUlvh+cDJ9G/aB4QKvJNCiqVSU9kPv5LzqWe5h
Ur1j63c1omgOWkkDYziiLzxlcFmDJGue9MhNW5Onx149OD4n3Vo9Y9xHk+LK+Aua
Tly8bT9pPILXW29IekTHbLgmw1yepjV35EXrbjGNY675gmwYsb4Gw7qwFWKIHdFv
po251sxnwxPUSzy6Af7L6m/88nkP4W2brZXeKW1lRmxoJz1xgyQCurQxN5E1SJrG
MVTsfuDJCssbYuLzF7hxv5rkzGztMIYEVSaLs1SoXXbcJIm8TYJWM4fejBU11p3o
szXwcwA/+ps/wQ7LVKs8p8YbMylmoiPgf189f/Fd6K4imOEY7RBZrCX0tjljFhhW
z6CQ3mHL/7Sgp5PtLf1BqnfMh+qtkWuWAccKsNtbvefPZjJgw7ek5+yWWpxcrnpC
dBUZSjDLF3uSk43wbi7e7fbB7Boa16CS5eFRJuJfATFW9xAL25S0YBl4paRqaN9M
d4BozMqUfVTqDkM853+m5WH0K456zCvbAROytj5sC3IoJZvmOUQXp0DOk/p2QRLS
IsG271XZAFkUQZ82UrElZGAXYqBxEZgL+W8PtuZT/QqdL0RXCiM7ckUfc07BR2e9
r3wLoFs+XzYhOKEeQ2/3dZChEegOZbqHKZhzfHvWyi+nvQHOXfz8AqNAgG9TC9ro
t6Ef+1sxOqlSU9vI9iPu7CIaspxHp051InJz+zdXKETtN0fMefMxCFop2vwRM6SB
pTGRkOi7Bos3gQrMr/8TWNc6EWiHHNQkFNtSpYE4pcOZkmGMO4wNFkoXud9ExHJv
YaJWE7ygtsdB14EDkXEHwlMZj1AyEcUGzgfVrKgoMAHkfTXxdexPKzGnuX0Ll6PL
emJbgJM7lSsLReKHYPadkVu6H25qPUP8HMRAsCQWGg6t/ugqL1UI0LQ81UUcraQB
ZrRdn4CFoyU6Wgy+Qe87jjQsir/k05skGbNWQyOJhh+ESCvhSxsR6/x9NX6naIUW
3YGxZDeAJ6l0yrPuwgPMsIWYO+ETSdxm0bdxKwGXkHfvTNit4Wr/RwdFtqcRs1+7
qf5Y7GTHE5UthD85k+ckfYVATm7phYSOEilVsA569WvWgK/sm4iEL+w3ikeXvPeb
w5oibf2FXl34onYvwN9j9Eok8lVzAJoYht+3OIi5CYJx50X4g+evwSFWfRpfQ4YZ
O1bUQz3LHe3oAXi4iMlII4KFuM1hIXBNIF04iLr3t5x36g6Gd6DWF1wubKdEr8CE
vLPEygzs2pfyXBIYnwOqEJXs8D4D0sxPfdJVtx4uUmCjeHEd9jws74TifQGB3Vjv
/cx6U/6WBB37TjjjqgCJCDNwy+fG/BVaYeka+B6wqRMpyd/++UnGlXq3clnp0Kku
bV9nKjnmSKvcoVdnxqXD4m9itoOVNT7+SrLdW5xy0mA3O2cgogG4Q4k2crMFMoYC
eAvU2+1nW4vgg067LBfTifYI9AXIVLQY7RH8R1MIk0LGBmVXwQk3YoOn9r+mreY4
Qh+AUD6COys1m7T57NcFY+7c3qlNVfNncuWd9Fa11pN/UKnvwWWYoWAM1Fjg8TKJ
j8p91sPpLJo9jfuhZJDHsBi3myLG1cxo15YZ4IKB7upcRQ6L7t8fDxZHQ2UY8utR
ZVPOcBvXrKOpgFMSZbIoOntbiebmAQyDE8staMLp6a7uPSmlAlrDIBoSOPZDzq5K
f4JvbnZwZ58Zy6pmntYapOMuJdyzYD1bdtFD1zzHoKV+QuaSPIQLyIK+rpoidxRA
d9JfJOB1DvDimGIOVK33kDzE0ok9//fsdKNiidm9PgTGTPfI8zaXNdvZNUWlQvqA
u6huA2X/ECmHFBYGAiN1bKz2129ycXdSsC267wky+jMy8MUNUHegdO3HQ/kXZ/rT
tk+6+RtQ9hFWDx/IZAXPXRWVaplWYH1YhnCASxI9Cyf4pn6ZN3cac5og7ZHre7PK
9E2uwQk92obwIZiLu1GW0z4sTFIIqzbys9gKtNsFZ6CeQNOsmecYsVmXVIatrPgD
lx6l6mbYRoWzP3/J7bN5/nlbYAX/ThXIBFJPgQhLFRAJdQpD4PqNa4jPCpjpgqzm
Ob87THcjVJYFBmKRJ21pPONZEGncjLNjQ60hDGPt2+X/M/stINsHF/StgRXwnl0g
5l9Gxts8yx1pS6NI+oO6ssLzHHFh1kTtdoOcTguF4K2nL41If8cCH5uq9whjwNxh
1JdYxhBQKQsM2AqGsFj+VGBEURPLX11NTV1h2thBi4WHib0/Dx8GvIuEttSA76iU
RyHE5uV0bjUEph3pIbRoJLvbjzI8CvOGMX80oRDU8fEjSX8T5vd2K6h164SYNjIs
Qs/Epb/R9wBTHgH3PhVloThNT/lSjIlZ9fd74XCa2xVfMMacG/6PTwFB/6p0H65F
p6pdf/tL1cQXGy3qVVZQ9DWkDAuE5VwPDdvKc4/bBvb6vBsNFfE7aSOCfpLgnbdk
vua9dD6MjRDy5AgBBbO7UUUE8TI0yt6thMRdaSjGkx9QGl3jYC2ark3/F/H3XQ0M
U5/ldd3TER1p8oLumu00NLv9brueLY3wxoLMOjTCVq0cgs0t9MF1P5xOsGv8BHhq
20B7bGDnZncnHVki0kMdJYid9683WXjjSsSK1HsGLCzHiW4dWs0khEy2gD0zoJ/A
DIoayDn6Haqq/pspSkfncL3IwgIkLrtHyjqnEVNTZeOX+JaUpYZSpEs39Y8JDvOI
vF0+QTYTGLoClw4v2StNT3ndOmaqL9xxKYMb+fptK8Y1rlqkKZryFuGp2jz1hHLt
7EQzG2zfnPHGqh+hoe2+vCBky7Dr96izUa5NM9hsCAh0Xb+oI/tDRW1t9Ju/cZhQ
OpWjMFdeOu+seTmTLz+ouzRGKYrr5jwI8IHFL2ewy0wVt5yHClir5FS7KFOM2zuX
Acwcr0yeg1B/ZabOcf3rMW7fbuncZm+yheOd0Ohy07nV449w3cBvzODDQWpN390c
3YGZrG3qQynuomJngmQhPn1xoLoJ5b8Rj3oYfbA9uuAKXk0MIjiZt76g1xKIZBNJ
YpPbC7w8jBMxApBaNYoc10w3mXwXpKW1sFZvvoY4ohJcRJqACtl2q7XIRqajvQWd
QIUQIIHYTvSzn8QysaFqYT2cgpfh6SiB5aeiA37/1OlNiZRaYTa4vXK7XeChM6/q
EVknJQwPVJ0giTVs2/91K+/BGm/17AeROtQsbpe66hVEVmo+Mb4/SEhlbI6w1Nk+
IM3DNy1cqjmPClFvzA4wDTbGav0CcBqqPV86kaqPRCQfJURHxSy7R88vHu8SDK/n
1F//QKH7JsghdKKGIhTuuXPMt7r+ueCBJ78TbSnZjqqk3v7qO5/8VSgxainBaqpD
uh9iAjRCifNdbn3Z9xDv1gV6GPHbUSw6YWHCnpHe946X6o6yIdZWPqZqOEUbdShS
xVP5Bbp4fggBlBEH+eRZa7qZONSKxwmxqK3Cz+ZIrQA/jHCyr0V9+4BlAtfT0jjU
O/RQITnDzUNKWRTNGUnNG0af6GYCI9mU771pe+FE7VKIVXNfMQMfECA+5kXGhdh1
/y2EQvCSWqWmyeFTZc+RdMuKj+0cdXdxpU63FSsCiLmlWBmybEl3BNBxOSQwko6N
6uhSfzTbGKzwoclJISclP1GJfgfzS74sU51O5Jtuz+Jx7cflXAb8PJ5HdVZrI0IS
tRkOFTjPsWR59vhhj5yjebil+BM+v2/bSW7aO9ociefTUgEQxPwh32YVYFdOY3jP
AkpBMMqnrpsnRswkx3LTaPujtCufueOEF0SUP6s7z4wBlQ4LWXrOxrMbY4/unAmR
QZD0ccm8ovEVqPc/7t4YAgkhcRcEfk3m0CxeNkAq/3nIfRAJsFijm2ZixlInhMr/
sB2jX83bWh67iZcnA4J9P+LCqBi0zkN1kUGyK51mG723Ldl6qJb7QeVtn7EK1lJf
IXZoBFXI1MjZys9vijMEsdTht1BAeOCbwQRsMvrHEQk+XYjO23XhsGC7t6/2KU23
jtgT97ZaXw3zu/zv6nT9p5w/vWPC+SWl6U/uY8XtbR5zbIwBicdKxZGzll7wl1wF
PUOshFiEMr05uHvzUBOSV3XMdCq4yQMmJTkhdlfuoYSqQTzHgzQY/s7w+/tZMLZP
A1puscjvFf5kiY3uNWqW1kuuSThPYkVB8mTB2ouNhjuGGYixf9tnQVD/AUzqvx4/
urJpXeUG/j9uYs4j5zoCiP0brdl02tKNn55+yuTUsAt5AS3J5biFF/UHHtl9J0Fn
1x8W5p2I/DiOhQtW8QZYqqewKQmNFaW1IKhukMGGFONEs3oNO6VymMuXW4Wnc77z
Qb7ucBq/KBuOpV04ggLSe4ZCizNVyPhCpi3jZcvH1eCe9OfG/vDeSZXUvPKxYB/C
9BMoPYu8vzTleBa00buQIzTCwxfEBxzBY1jKJ+0ieP1NAnONaeEG96/h0egMRewY
vmoSdJKE7oDD1TPZefALgK74Ljs+vO+blY4KN5dWophyTK4cYAPfdW3XKVfwUZz3
bfG++/9AQxt1j0QSQWVISbaTbpgno/doa3uxNFg/cThE5ff1YxdGRuYwsxAERiWK
s1MGDc85oj0uYNLm3ks3h1/G0+ZH/vqMh1L/M9LaxGx/wCsYBG3eg6hrAQ795tQZ
AB0zbTbOJ8+eMp4BZdmHzIx8KWue9Di2BULi86UTuSUEVBU9yIn5BqWFrdRO3qOk
iOYChHyzqPrvnESvmlAyWJ7q0f6lCk0D8c82RfjrdvbOknyZmEKMZidcEqi0iLmm
wFq7SPHDlP6bYP5uMob9VatqShrLRbGZ6fBPZrzigUfT+P8v7DvBej7luTeXPYcZ
1hC2vNOqTiOOw1WRXRwA1q/F4iIojCf5AGSVFfjj4RkjuroKwBknUCLV5szAqfy3
IUM0KqW1HojLbn3bDtvzqkRTFX9WOLaP6BAjUWwBeBwGP1U4OeHeOS5K/e2OlZna
gu48ZxJS5uAcf6Bu1CnzHkVIZemYz5aEAsx6Yh4rUXwEHhI+Z/3VQhg7bpYuh2d9
Bdc66At/1D9JKNYOb4HjcJ1S3XJPkK2uaHpEDXC5IXpM0Me9ly/Ze2u6cFhnrXb0
hreRFiBOLBKoxA9SS9v3OC5LUNa95Repvi2kaXAgkBCg+D/YEMXwED5Ds+MRnh0E
5Q6Q6QWdF+ljnHr49xPgWwEee7DTLesF3zzvkuxVSvwXGggWeeUl97VdzfvJLuEq
bkJ0pS2j3rW2Wo0/YT763lLl23qonVJp2aNwocEdN3unn4ddJLCqWasmUr9ChL1C
/qvt7i1EmC6GXxJdaQrJl0yOHm7zVAbN6Ct5PaNYApP+tmqH73GDeRIkzgTv76Xn
+AYLuuhNIPj5QlQm9T78IankTJSHTodwq0uOQZTTd9hsMyomkzwN/G4w8Dbb6Ynt
NGiY8E6krMruU+rYyiabpXaBuA9lZzsV4+4hgBVVFydIC3NbJ7s113xzZ+hW2xHg
bDPdp0dVKxy+5XglUUoa6OwXeA2thDz7UTkSibiZFLmX+ZWIZoBIfIqXUc4BRjOQ
w5Dv2Wy/l+2vEvfV7j/rE58Tug1CUued7H8Jf3rcSmLvEA/EOGP/jdDJ4AEAV3hv
/bF+HONZoZfjeVrj8lxNLMPoSoCbBnH5CA2PJonNPuGL5KxbYdlv4n6wbk/wGey3
LD3VxqovL4T7yW00/kk0Ub/EQBbbR2b/zaYpe7Ow+Q8xQJlCqRlA+/7/YrPZpWVL
9jSOuWH/cSIXMVXyZFVCtve0je/IYTBkdmUdPG2dR3VazJil+CO2TJ4M9Ppa4i57
WeYR8+aL+fvT/sZSxEoPlvDRFpsLc3Yb7E3OVA+uXhC685NgLRYORv76pHB30lD6
Qex0QdOrgMLyhlKuF7rbuVyDPExz+AkLrg7DYat/SPY0NYki23SiSe/9m6EfvbQL
rveCmDs4zVjJ/bVkETHXAr2nBkgxSOUwdNGNav/Lam4LiwaEC5dhK4qafJ5QgwVq
OdME0ORf8UFm+rsmUGVraS5fMfI9Dz0Crvc0HMVgWyqegSm5tBeyejV/314/HsCM
p3WAMgmAs90iaKjt+W+RJYq75d4bVGvQGQO5W+AEDyYssDBjV1s/JqUA2AsXkqyV
4gVwhIi2Jtf3KKl0ZzEq8+9pXF3xAShL0PzghNu/CaGoIR9S6SO+ySZd50Y2OOqg
8dU4D7xdmKOVNlNBqrWZnaeeJiVjaH1edyf3Ns7Mpm0fcwJeZKphHHdTnz95ANw/
8hBgOMVV2VzTPCRYyc+ozAuxDfjciV3phKy4vOOuUsvXqGJAOx4jeWOMf5pWgbED
LuvRdycHgpk8lVBudiDqYv+hbTLNgTvmg9QrBOP/tKq7I9DGvQBdxlExfFvnpeqG
jOqd/ITUvJ3z1deNMhgybnpR861L8t+gvjRzw5bGRV7Ir9psVjJAMCkF8JYjXPhE
yT5LQO4X3dPklqDCFInpokcbhhTTmEw4EkMaiKXU+FwVXnmJeVfLvaf7mo29aYgg
+IE3s+wab6fJiDJLLn1QJL5CmqtF77hhHiblSF0yxgaZGnJvWMxSb4/EMEhzp1Zm
+iq88dBOzjkbgDTVkRu48GLe0Rt2uyOgd7DILxkNj+3eatiQXeMjQrN+dptjVUEU
MevENyTggVsTcHc//+GTcc8M2loAlD0bMvPTSgcExKlYcLA6qpNEsH498iKkMVHW
BOrQ/cgfaJxEqEhhzG/z33L7hrh7defpLRBhVgMIR/xcBbtkYZsq2ClKNM3Dpoy2
/+Un2nlXIsE1hLTMh1ROCNXFkYUNa7aI5Frd+TuO38IWQJU0ec89e5NTl82YOVcL
WBChSsfX105+7MNBNWGAjUmVbzSa0rS4cfXxEHWxfYiSg9hgUTSE6MzCcbdqSIvT
9kTKeQOAeKQJcRkD6pdhgVKxh71EHm4L0yBnTsbWfB3UmuH0BDCHchXfE/XskY+g
FNpjOIILnYHCEMRXEDHclflDAJD9L1zEV0yfZl69CX+vcbgItOMDVsnMSp7/NpI7
NjJDI1bHlM3ButtYcHWXUDfopZQUOfTfiG/h3YY0IdTC9N4ghZnxCb8v4u84/fQD
d91mDfDRp2VY/aH5hJNOhgcY6r1O7I/mQGn9BMv8vhgxcwH6qQ02S2EiUBMto2kI
Vs8DCbRzNGgZnXqzm/6Z5y+KrqwpC2utvRaxZwVn4AxBNY044v5CK87IWHUtfiza
H3a9byX5RvFTezXEU7DZwQjNs8FIQ/VJ5XxxOboJPyII8z5yPWk0AAp2gqj9Volu
mGPrALRVDEYF0OP6O/qwoRPwAsPTcHrYa316pVTRmd2+PLQQoDQE5q3ThPqWW7A0
7Vigpxe73E3JtVrYMm28wtgLM5rS8UfN1fP4Kl8mKenEujVitcnf1VLRZMSfK1Xd
39enXicfo5IG4MFANi34uqLfsw0DYag86BSYXqS+IBzZovjEiXZQs4sqRseVGkmE
YhNltvoqD/8eF+TN/2ZnRbt1d04vkMh0MdHBhvUH07D6qHB20H3p5CrIiZghoigz
Ov1z4T/gquX70ljySTUv9bFCCoPxIpoFCi80C75imRdaOuOA/qykay6yzk2eHpgf
zgbfOh7wpk+xNKoZd/dAC4gMKqcXYMldJBeDXCi/aDI8fhnDkL8GAXjNRNycoeuO
5J7xrmp3Wb7bshlxPVY4FM8D7IR170LaT25W4ZzW8+JZ8Xkp+v1zEj2sH70u7886
+I4VDy9gZDhf5QvD4X6RhpmflLrK5Yt52bUu/Lu4sJmyMCkPzE1krYaAdYlaBPl/
doa+IRhiLczI2QPiYoPQAxmftiHCfoi6BnuNAoGPNtxsobcPM/Vv2/ku/cCedUAL
hai97q9mESszvVY/6eLdSQLfyidqsxx2iD+x/SX6Qu1vmTeta03sCd3sLIrvn53G
Za5/jCXlr74BTrTifYVngvteZgRDzpRMuA8w+bKrd9dD97b89Sdq8yQU6i3l45uX
P7wkrwdCqnZGWdGYgejgu3Wv1sxnVtEUZI61Mlmkvf33vJFCqs4UGF1T1KQgFhRa
yrpomfv4Qib0xxrqmO1QERST0MpHIan4wl16kgZS8NOeL8SxqPI0MCsw/3QzqG6L
wjYCSdd9ijjdleugFjhJNGsbfHrRh9XIcVZeVqY2kGflul4tL39Gqr7+OXLbLjdH
riSUdTpJKS7QUiHnl/wBBvcFtuifx8s+hcvyFZqdDzp55YKnkKPr/ph6AwmD7KfG
zKNDxQruWtbF7ywCHjKjzW1p4Sd0aTS+xbMRJqC7w8Ylw4RSHZSQlNhmXjCvNA5o
LCKOaeq1WSkwRYJTmpwAECWB70gwS9wbDa4Q5ae+iYlwH31qw3X53z3ZlO1Rjhr4
G1ejuvr/3AZRaQJYciMipJKTHVBvolrH/+u8oCu0q//cuGwnWfmhZjhxQhRAmYOA
wUFus4iY4cwXXMh2K8WETcpAA1mLOcbAd2Ca6yS/hqPdwf9+v8enIVonsCiu+esF
PIuEu//XdR8zAU77hLTnove0GVNeIloJKKXGwE5Yi/SOkXLlmDPzGao+juVjx6KR
MIgE+50lIG6dCq8rIfjZigB9Gz0BHEJIoz8qBoTW0HtTyU89AFJOBgubdUUI0Fwx
3H4YfybVdPqxXJcHQAEZtdbpAN/PEeO+0lHv35x7lInEhmIVasIa05l3YY+Pp4zW
arHgWCvjGSLu4Nv52UFry2J1T78HzCeaeX8f0Hb+EGyUCR5AOsRs7Leto7/6232M
sVOWO1IrHtt1eX3FSYAi1lUCSr2dObJy9ShclTgrhdsZKtpCutbDIpkMR0iW4Odh
ZYh8euD7Cpqa8wCsOtiyTpMnMTqilto7fLeAoiZCumvi8ceDQ8M4z/6J25tVcYs6
qJUG9r2l6f7YM26FszgtDyY9+7pa9hm+PqQVEhEjlhIA4s07X/uBGZB9kK9ao6hG
CZuHvWt82zt1QAaWrpYrameFGROcJyuTenCIiqN/x/562+GyTz2ad6D6jMzK7sy2
1q8pi/BdrqlViZrdkjqDzFilvEEm+Sm02dHaaYxqHGNZNA4gv64cFpGpFXctoQUl
KfCT3L5TrcM22tjixDbGA8Nb//8BTugJGxuH3z4z7eOkB1HummYlfFPj3xoZWeYE
FN25VrYNYcsDzmKXsltYgzETeynPojnzgDXUIyVGtvqm/5G+Yi5EvIE/GG5bJRXv
F9S2Ca3VsHaVKpgzguiw9cH8gh8g/tOru5b+61gnXge/eXUshb6Wa1nZ5ledNgJo
kHlEo8/SnHGc723RHwf8U42jugsRXP/JSdmjcXYNf9y2RdUFxCuh+/Zzlljkvxvd
vtH3cVaamtYJ7NOP6nfRsgfZUvKKQGPF9JslI4jjJR3kgA6l79JzPzxW2Lyjexbj
XaOyEdZeJmKQkWgwPYTeKer5QaPriv4DftMdFjlU0w08b2A+tDmdUerzyH6gLB/k
QT3qI4Lutu7MCKJiYPb9H2yeSnOS+pQWtEZtb7GWkx3di3Qh+uWrefteiReHIC/e
EJS7TY2rzrcMoZlsgedUOB9OmReSxTP4qZ8pquEzfI46lSVfy2xhlpV2SzecejcX
zSi9uiTmXkaJFxfCMr+4vEWzttmtDejYZZtMqWFUFc0tlFIUdInlmI2i3aBUAWW4
Rvpi/fwM1cTKoAq31fLvvsDK+KMiSqcbXycvucNcwIEAzfWs5CE1D0uSBxZp7/vn
sEoZCTEx2Osq1LQWUQenUmwtGRqMVAnHKQzPIdK46mTtTACtQX5CPUxIxq4fQ+Fg
NPJe2MvGGylMT+Sxn3lhsPoW2VvaqU89cPswmpVFI5y2xJBzA/QcXhZvBq686xU1
owRYvjd5knc5tIxq2Xu+855hjhd8bPuZ9Z0nhhtWKM1V6uKV8LybFSsHfonzxO6Y
4Z1on3h8uY+b2OxnXOz0vtlBw8VBGGm+LG6zlA7EUSNZ2FA5dGs4lBnzpNZZ2zgC
etWebGECd+WPJDRSShx2YxUdZB9k4mfNzcpn5eywxw3DpwSk99pTAI4AxQmHVZSQ
I0Gtrc8b8+iXapOlOXN3AKZv1pWVZlwn+xtU1+K76XJLqefOYwwOW73ZJd8OzNiw
DNmJUCE669aqPKnmwnRty8D29keiuda32Y5qcCV7rXT/Uj/kAyGBEyqLI3NDDRum
9gfjVS/sCKSy2KcU82GZ3Z5gr/GKuLdwAEUbGImUb7w1SWygn5lsAE0xL77z3OOW
jEa2aTnnYbgFW/d9nIFj0y5YkbmX7GnNaiIDtqktFIV4xjoSuba8xng+Ouzd35s0
g7BojWvxf83UoJASWxzziKub1cuz9y1E3kpRbXLWwRnxbZdQ0XBTB7vljR88/Gl+
xJOJOoUBuaOGSYCGOG5Cv5gCMA/6Bgn99pshFTkU6Gp3XTY5MOo2k9vpSu6cWLyk
xSoJcYpd5p9LkYqPKVideXereQKmH+847rwXaEYgN9axNfyGcdHS1AP/xAPY8L5u
vSQsoQN9Ce+xGMtyDeebSU6siZOJXj9AgLYbh31z+MvRk6hS0CgrbdJrgTNQ4YTh
jN+eBVPqMSHu7UucR+uHPXdOlSnfaPDm1rj7jXjYoCMrfhvdpJsqPTeWW4l0Ft3a
Vn04qcPTxEF81Ay8+Aa6qiKF284ZY7gTbuoRW3QgqesnEgYwZfJQJIyU7ipXjgAQ
M2oe3NrwLLejOQX0TkTncFtFxwce4vOw8mnUh3fBWgvuCnSxrUTGZHSBxpMEw2+n
gm58sPalqBUUIoz1lqzOQZIR0LZifvMVy3E8l5gzt7vKVEZSvTBnqfbsS+Clct8e
L6wXOFfUur6FWmojG8PjMXqygbkq1pIbObN2ef59ehuDX8nA0VGH7dyoEumBYo9c
6GPYOaX5pZM2+QhTpf+rM3ZAgagtDgGVNx3VbriOJFZRFV2QOw/Pod3on7t55SIm
LaKrVHEfwJvxtphtWM5CuNHcl0b6Xb+cRCJxg4gYt2y2ops2bh4lyKWV01T0QAT3
Emrc2TxYzsmja6W0YdvHwuJE0Ia1IHxk1GX+a5Wm/Ga2E/d45AxzZg6m4WW3Gn5w
R10s+q7uKETys1j8WZyrN5ZjgyyY5upUP9C6bKfUFZOrrEbDnwTLH2nFsKAIj16f
AJvdkJH0Nx5A3ffY2LwXHggnrVcVl25coRXPe+w9NKf+2y2iS3pZdejZgaYjF7i2
/bxGe34kF1VjPg/SLYX08SsZ3XZxM/0TO14FVADaiNyxLP6WpqeTvBM58ku8ZwTn
+ZiPiRm1s0xzMLSLqRjolsUsLEm3OgHJU6IHBvUmg3If6gd8nwdgRvPet7Ke79dc
jZ3INhWcFXjXAIf4PcaafRrlLfZ1T/T/U3zO5X9Cmsxmpmuj1vw56nPcY1AY3jie
3OEbRRIdMYYUl13BhrvJmG+I+39sbLi49xWyYnFqGjLzuggTiptauljYebRgjQtJ
AjZ4wLk5Fagty4oUHGTglPaed+YNq37XULBOLHmYdnOXGY+PJrKU9FmAv1Kg/ZU0
Z7x8sjBK42VQXhFB/Kp6aMkYiPhW6t6c3V+l/YkWHEqwC88D8F50uKPdTsKSpSID
hIWxUdghGZZLr04HHybZMFXBoy7OECTQZsEvkaUGk+o1cdi975JWxbY/Mauf1sRH
j79b+nller8M3QJWhsvKYbqprdhf0X4iUEI++J7X1xdHOpMpE18e6bL4AVdKdQfZ
qWQkaHzCq6LmwyogLGlUB8CV3+zMoaES1dV4G1hl0upcr+tmyBash29XrdnhXGE7
uTKibMMSlSk7AP8t+i33zilzGuGIAoXY8RNgJaZ2g+t1XJlJaDLzE+nfrczKZZE3
r7T6j3mAVAWeaOwYfxg+hXtUtkD+pFIo/Nk4L046J/FkiktEcWDANzlEDDJZrTWo
FiWIv7TXU/Dveig2+xCzmRHqcHR2zGTn+APqqVX62dJgU5XMQmBihdDQ5U2D1b8W
kJHjLeZHDxdXlvAS/Y3PgiSe+8fu05jld55azUi1wP1VY8fyBMVsPpFr/Ghi0J+A
NwXAdFBugLPVbtUzkHX7Ohl4m+nDbQbmeaxXwh3oq8sOKWKcE7/jD3BoZNqv2N+r
G643l2qDoisqaxB8h5EsSvSHwtgoWuI0kU/pQJhWYDfc5E7WmFw/N1dESyji/kit
mr6ixY0Ev6X76XHvsMMThSQZu6MV+RobmADESLJr04CzxdMPw52Oen40FRFwoIHP
Ket/l7LjFRP0DolWCJILnK9OIQY7zioPOVWVsx/g3ASkcT/S8lyv7aXKSavlhfxi
RsrFkBf2asZZ+9L8Z8QqRfViCMqdnC1kJJvBY+x/icE/CleXyua+f82y7mIp2UlZ
kM5eKXawOfbGq3H9rvkazs6A+MSWAzBtkXNM3SBNC97RUNDEDvfQUq2z1mH0swPA
S8VxaTMrU7M7+JJwsmPCXgAD+moXuld6oa35KtzfZ9GLKMdUYRCzGRKo2u0KG/g/
i4tOSv/wt5jHK3Nr+aqXuQeaZnEs+vvK3LqJ4dct8Xc1wXPR4HIqY9d70BcrlIgK
Nszl27qMH0vLLVgZeZCKKeiHKNGYk6lHNNdMlAC6i25qsdUvPaXk591Fwlp5keqY
ow5EeWY3bqOhEBkqM/+jfaF49JNBZ1OZzFN8qJx2GoZjQrGVF3GzSuSERicUdP6x
C+/Cv2V1qZPngSdQG5ma6Z8IfThsLKf3zW4u5/w4SyUyRLHkBZj3+e5gthonp48E
Uzf0yl4FPULBpADDzwSctoekTneeNRQ4EG/nOabmrcfNNiZmzmKCtkjs5t4r6P1y
ejhFCuluELDZy4AAA8QJb+3rkuoJiEolQEeSgwAQbUf82xzKJAzdn9JQFykD/KUy
eEOcMSa0k09Vt9zCLzv2z10RyLgS4UHHsb+SVure1MjNrsqJIbAAlq/0Qx5TIRq3
8wxc4VYxX1EAJS64Sb0WUIuhi4Pc1cPR7cSngar0tbiVaMZsHuiaoTd2eEWqcYva
W3IrIVNrDGEnd4udnCNl3EbuTDBqy8+ICRTABo16FI+qgCnx1mjuRSuEmL1rdcIN
k3COvmFfxAeOpmJjE4hASvHRGW9+uzF1ugLNSh41KvPkeyqsqE8QnsE+WRr/sdD0
+rn5uNygf/TkxqCNqxNUX/mbk2ChTj6M53SJxDkFyYOw/FkC4uRyu+Yy649KrFJM
y3x7G3q+vy5Qbb3Yjmhd86qFZI2Ahl/ath3XiCU5lYhecxnoaIrvS422zj1Nn8C0
BhfOEVxkYor0WJrXggGLFE8SLe2xPNsTGwu6nrFS0gTHZpHHlKRdM53t+TH0KC0r
tD3BxPfNjKK1PX7L4BszMoyqezgg9MMm///JpiYM0FU/MY9cBaECc3n92jF45+oV
j8m3bDVbuNlO4GEUWFjSv8GL3bgZjzT066OJFel45I+jFQExMbaHq5G6j7gImE3Y
7dseir2HAZINaiEitGHkvH06Vp2Ov1cw4+MtoBP0bYj6bmB4EAh0XRXWFPIWMBgt
H5E99i2lPf0ESNeAGeAGeBDKK3l9+pVFSEZB39BEmqW8VfR/x2/PwsFLtX29Yj/S
zy9jb0b6BTxDiqdcSF3nypJCftHysQinOp02tWR9XwCagTKVuL5dSeKRMV4ZTK4t
zI48KUJZfvEbvFlpJEjO90GL0io1Ob8CVt7QCFCeIYGTV15vr1hIBW+FvQka1D0b
UhvAtHFreqs42cqAs515eNGHxgPJjOv2BRSj3nrhWxNrm05VUsR0ircgegG5Tp7/
nsGK8zpuHrepqbETXyI0XtzXt656jw2Ccw/Nd9FKXnxizUfvTYKDAZ8D3oerfe/K
ZovjOiJr3j2TCpNU3tM01dCbOgZAfnBe9wmLfteG7vkOtDG/ejYrX458Qxsapy5X
sctGJvXGLto3qKURUWa3YCN4WP7Qwu9YNsFGr1srGPGHqIqri20YhFHd1bJzHZWq
UMbUUiSSDtHd5fOUkU1jHGMu0T+FLXB3Rx8qJyCgwHgYgMwrMgZV3oSx9GHjS8K5
ccQS0VUvsy2pDmzVInsKmL9mNbqKGgFBfPZjxocbBJbIco2CgEMXIc5tk1m22iQo
0hGOrU7ySBuXq0zGsWF9Nh3z9zaVEYD4mej7uei6nom7xWNw8SiJYECeFIku2NH3
Wf6SDZq8dFVbT1HNLtLV2CZEU3/z8EUhbTCEuDzCQwDGjICwUSG589RdruWm95ZN
arD8Qod6TfwTX73qyd6WbU83vd1Y9uxeukfp4vqF+4leWlInHZlzKOoxNvsgACnd
kxBHme55VUDoGXjpahJs0hHfxDgtSUuC61LTlupOFoKEtnE2hDa/uchw7EC8zIve
h+Te2QZvHfg9DLu9JSvefsiNUpIHlYXou2a/aa1VZesmmm99H3g7J5B7DbQrApf4
AYo5I0afVc8SW8b0tUGkp141Yv8kgZuMeXpHWtwQSGqueaFo4Xkselj2crqPPnOh
MupVYSgaGLYOCJgp+UvAXOK98FgSSjoAgERtqPYOB9Jpwv8I9XG72TgeFB7NeXM/
tpewUImf8bPu7bpECUBgf0EVIYbGlsjCycVLeYr0Mw0Q8ddM9uMkPAJ8vViJvQ2u
C/xrivWgZfDMSYPX703MnuCbp7bDzz/g5HU9Nyg5AWw5TGJkYAtDxL099a0dpZRE
QsXlzTPY4uqfadQXFYeyxOw4NdliIPcn8RCsrNwqg3yrLryTvh8uKZxwwHW8GqZk
fBNb2oab9ynIh85pCULvAOLKTQ/9bnPRuvHW+Z1YsW7fTvQbfa1VsJ54dv8tIYDV
5kNZYhqJpTQjCR9sZKXZkzTNfkHJp1UVpp8AusrBFFupsgHnLuK+SikbUk7GMrSF
PpSoNzdO7bP54ZjEaN8obk0ZL7sxffyHB5li8vdszTeRBpziOB4vrcbjJQl523gp
++rhk19m3BdLVSbgFQgrz8bsR7OmNpu762wsE8ffbzf+4gvA46F3Y3gTUIKNMamc
o2wGYNbea79Gtcg76HIPC0QVGOTjIemFPcI86bk3mczbh7/epZySN3ypjC38BEln
CxcK9JZIGErf5m8NM6hI6vptpPPvSHO91p9y/+n2jq4qGRZZR0lQYy/oEXLm/f25
FJBbOhqxCpSdikYtINilID9OO+IHM2VHDHwuWoDKI6ddrU/iCOjTzwFW5oJUVRTY
I9BsAyeFspNDmUiArF7GhNH2qWOl2adHGtnPie9kTYb1tDbkJhhpfkOyTX9FLKHp
XJEsd1BMq0QyIskjOw/kEymVcUiRlpA3guNqtTIVruMxC3bRaytwQ3qzwA0IDyib
8+CwyFTlGAJqkEJJkn7gNVXOH+oyERm6Z6nBNu1Fm8k3HhGL9d13D8XwiBFM7KCn
mQS4v6DgK4hwkJ447cxzGZOiKLrDn9dGiYhBLYzr/YyJxkvsB4EO4jC4/xXWUiYH
ZiRCxgjKhH5JMAy1qT15cLgI4SiZm6beY/dQkLR7oWGERdgoZ1IQd6yotNdgOU4d
uReL9IfZCcUlW1vpQsvwhFDwwRcJ3CI2+IiQnnAW26jwjcx29R/uk24JEdwsObT2
gJVWwxdPtSe50B5zB5CBo4BZwOtVhZWf35SzTPLODnc01b65g605wq4ah8KUEWiH
Y6cY4k2FqN9ukvnTagv5KsMG0u8CR56r55HbPC0TpIKubAPyuUD3bm54s3tfyWrG
UkuSaI7+MfLO4tkvU0u9H9CqNMwB+tm6Im9PMVSBiZh+kfWp9VNWwaUcGjHXAxQs
78CP1Otsibx7HuI1GwLCkp1LEZMkzHl35mjHaEuHdZngonMEtUHIGoVanZAh1/et
jSAtQwIwrcwqAXWk0FlfR936/PsE1nvlgRnWzi/NdJDw2TmvqXW4d+Z81IGmqIm+
SVa3irCplNJKY0txY7VE03AavJSV21lyXKTWoE99fKy7Was/acaWeD0F497LNREt
qRm/g4toUawkXtlgIvJY0x3bvG3B1nxEhkaIvtvZRthgs1ieio/cwqmaaweBJL1F
CWjl7HnqshmDlh5fe3tG/YzeKQzw6riWeB5F7msA2RSV/Ov3XPTQMCkruqtFG1Cb
1mrFh8Iqf9Vg5zlezHr0nS1OYQg1AshACTKJpsySXrYLW/ggV6OMaHYz/QucMKpQ
Fl7zUnjc1+AzPiZhYINFFvIz1Kfp+VF4E1DRYAIyzdUQ1nTgN/GsiBuH+FFgjyZR
xM9UsxpErKuX9Po1a5rgz+BYKXSQRMHE98Mj1Jvk7Ht4O8y83PcGXhxzcNaIOnge
Du+9RHqdeJjka9R/QyhogWB1N/AaC15BAzatd+KwKic77XdITs1x6JxKWtGGz2lK
1etk+H1qACQFO8TMdpp/YMNx7utCZFnXdmVZwMnclBYwKYI1r6riTHeB7VHgZZR2
1Bf5dSr4H5k63j5AcYQ57sURPodVEwEeYXdbxcK59dAkEiCV+8YbltAYssMOuxR7
TaX67B+jZX5XtMC6SNLp8nVrBJSEbUfJV2YCiOm89drHEdS/iUT9TIOvFHgB5HPq
0xNeE+AjOSyxpNf7mtuAnT0jKtXHF4bGxmcwP2KikO9jKND8awQ2vO9ZmsQHhQQm
Ml2C1RuYsZRnYCy1mEhz4M9fopZVs9ZrIe0qBnvGaOvLrhn5zraWNiWvoOo787C0
Nr6f3cAdConIuda0MzoiRpGBjfKXy9mE+BzchUA/os9rPAf2X+AxPOlwrGufhdHw
L0nYtH6p+a2+ypVrViqQ57x5o+MjYBssSOs63MvwnqAFbec6TBgOqiVWkoFQSClD
DKK+iMDbQUjsbtJ/UJ3+dCzVoMRQvJwXyyaHB8AIzzYRyiBXKkXXdhY+ocuijhBs
SbyojU5ij6R+5JeoqTpq4gOMHcz07BFJ8AHtGw+U1roFH4svSfGOreuNvBAebujy
c3639O2W+XgPu3ZQ1G8fmYX6+itN3T8R1tjPanFc8kIXuhL9S71Ttb1vPr6jm9eE
3ifaydigm/R/YdlUwb1UExgPaqPaBuusieSRI3esGToyrqUXotJBueUVm234xtmu
1vLn9Mg9+KKVK3NT45a1W7DW+jL1qoxxKHGURNiZO37BLMg8kXDfKYDkKEqCbd2w
IGY+kzQYlgaM01aXTb0T4gv/gHYJxtew47dOyePOf72KboFjU3PHUkWQlh6IB050
zky0Be6uQlyolLSDC/3S+FwvF8DdJbmeBP59JgR5pxIclZ5uP5EFfFs2YIPRmL92
FGAqOyWjnly4fUQHtAUsHV0GybgnaKMcFjFn7G8mucjqriikojC8EC9VMCumMcIZ
Cq5r5iDaMFdXL9TfMkPKIK0+bG0gevjir0z65kSPG+jrMhlereUddPIAccyiHyl5
u1uBzMRjsz6T9F8+RgGhsX702Md6hU0xlsDqhs0czwYm5UlW7EfJ4Ho8ZwahE8Mo
rfCRtEk/dJOD1ndf/W7ncw/pIoU133ttZfME/UMx2QAvvgQPYYjg5/a4fxpoMdvO
Js5hYfN9mQCiwUMu29x7M9umd+t+gTgFX4DwUAqxKZl4R3o7xbDYgajI6wukA6zy
lxsYlLEwQHHoBaDVAx5tWdgGOXG50a/N/fvTTO5dJ9Iam3hnVTu4EizQt2zGZNW6
syKNkGnvdftLwl0oz3vZTS+lJoOSNWl3nuFTXBWU7kXX1TUdjFKruY/71btKjKNt
xd/vkOq+aSmq+czoqT5N54WBHmi7fb0VMZ0SWK7YmEq7WZQERKmondQIo9WZsHnl
LKxSectsZDZGB/Dkg6MDqjo0tr8gmFRAviAm7HNBG3WDaSnUQTKrfzmVJZu/C4Au
ijlHlHrtHfXVtchVXwpyoSzTK9w+3q1Sahw2PBQ1uMONevUwHRRu9UXKW9NtgOZf
T4ccthixBZuWZc5Ji61uFrG0oVFqCD/b7XookCbiUSlkJlbmgEwLAx+MmiBxZ8Vk
c7Weg2SCB0cRW0nPa/fScY9mu6xO+PAD3fdZsC4gB0NcWkBNnlblWX2rC4XNHGdC
mb7wFu80z4HRjl5LqjHdQWyxKFESS5q3LOJqgUBuc6ZpydUP9fRcbToKT6t0hges
TPyK2F4v9gzag1qbW1z5hDPl4RHylBp57TQSFt2hmNLFRGecqHw2BrOzjOPplqA9
vIY8LB8SeI72fV/kLWikTdcHqySIGxzuUgGUd1x1HSGHt/AHtPJ91Q2pPVgypPPV
DgnJdRUnjwE9FIRzRTM+wvvxKeArI9yOCdyTDoZro3u0qOtgcM99Ss8u2CULRhPh
RPw5aAc1UDWYTVrF+GUMTdZM5myN1VzKAODZ4Lnmfu0B+NS08d56cEOUQCdSTHqs
Ol+HS7o3EWlT4m08YCuvQ834+MeOwSGc6YBfIJytUWQGFXbkPAoiyQaJCRbx1u4X
9B+mcuFS0/uKln2iar1NscWibWVxTbQb8ZpHvjUqUGbOwD1+uoHwqEQ5Kx9P1YgT
nWVkH9bA07dUMy6r8w5PToerN1VTsO/xkos4SQhzmcS4t8Ait29zDaPrhX9VHfAR
QV47YuNWKJ7/5PgLGkn5DGwKB4040IgxOosPV2NQTo2VjRsiDvf5mcN2HkDGkOGy
nE/mnHeOReQvVmXqrYag0TI7ya+4wQrJ5NEFghSBFIqudxX5jxm0vHf4oKPMiu1/
IVQB2yoaNjWRSqU5scPfSU5KvKnZH3OsoqA0BmLOFHoO52T7O8gDgvP6OACpxEdJ
MJql/m+xtae+sBjL0RcylSqMo0+ZVeiyTo/jnRWHt/Js6xLtnZZnHXF5GUNKjntU
GdZrjWPDuyS4OROd9nppMXl2ChnmqtHFbsqniLudriGkTeKSlwmgWckx7GT8bwat
NG/48eveuSyQJC1pWESzdEkUJSZtD2vt4FkEyQv0dR1LUPjOKdV7qwkVj8yXD3tB
K6Y3Hg1TM1Fgdkj/sSHxe8S63NPb72IGheq/7an0NR3MmbNKZr9ONw0O1wXxROG3
7JBNUKVwDARHIpEy4iRgWr9GfLL4lLdQiWbWHSJigBM5pcy5gxs4LZ5HKh+KTJgr
W4nmQf/Md6bak3VKnQ/snErIqA9WjL+WmFvXb0N9egJ6o4uK+9znjBwFcscSQeu4
H4YExtiTbKPE5EuehGBkupCQT85R1mHI328PmzrEOTrI2ZfQK9+05fylp+pa/2s2
O+8JyeR2aL5W9/ugPUG9n7YOWn+/Q4yzqrlVx4AJhb/SyU0p8ouwIpjgQ8z1PzNA
Mvkq3W+xPWc6EM7R5vZHaJ31M2I60FuBlWaCWid0xHMSpWgiSc24ZwZEosuOZ+wV
QkrQwqrrMGOxMNqUg5ra/J6suW9ZOELcqtInt2C8C6ijuPIapCxeiaMvqXury5fI
Cb4rwAQLfiBGmXfsI4GqqUUxC6+UTsUMjH2MA8osQx05IgOZgQKD/jIqthnXrTnU
mYZpxiWMxQglSCnUbUDAi1Iahu3d55zfwoXfvct7Ab/3bZWYFx3yIFpbUn7gGN0M
1Q1zPv35NKly880qtC141513viNC1FyMpFaC1dejpvBlAYM1ABOSMZcINmxh9cs6
sTMRQ6IBYi5VxwGquv8EXik0HwJc1HH2QoKIzLjFLkoPLREDEiQtRiJv6eZ8TJpf
wXpZkTVPGBuwcihi8K8VFj3xsh4f1wbAHxJNCcTF2/Rsw8E4y8/A1fXhpouPhHrd
pptG5Q+eeKjStWDWIVfeRbBU697fILS2QBPFEQo5/UdmrR4EZrYpFYr33xXBy+wv
7BXdhFPjOZdC4cPNi/boyBHsD/y5smfGKyDMD68wpQgyBL510mtoDmRy2YqwxKZg
WXei9A0TSS7T0/KDpKuYgnjt0bLOO4LD58Jo/c/gy8Bl4j0WHMdVo2qqBf1evkFP
nTBf0Wfp11uqFK2DLxlc2Ss4wrt7NbqZH/JArfP9a5JSJ/GVU4kmemvXH2kad0pQ
SfiLhVbsnxt56R6Vzasxl2ixSA4uu8dKsX1f4TDXTHOI9ptUEGTD+b+C+V4TNvPI
yWrDdy29p87Q+kEYsK+PYB5c4NNdlz9BJyqYkZbjMVmxR66XSq3HWxXyVU0f3niC
PRjAKc+iLLWegXEm5TAB4PuzGZLbZSNCda6o1luWIqx589/EiR7/JGyz87QunNzI
Y0HQhiK4rV0zxy86WY1UKf6ew7XCODnMgab1FM1o+irpc1gn+/m56/QN4lz1u+Ta
pCd9xKxbHrCIfc/ZlDsvwRzB6UBBYDIwsf8QMpYKtYvq5wQEptOsDJS4zRTVMyoS
0+6GD5Yfom62hjGgy+o5TpfHDdaOkLWrRRWPAH+GGHLwvkujuFlB9RGRlnbj0uIt
S4TLjEX3ZTcwyhWbcHpTUp0g1yVJVc5oQfyU2GZ0h2zGICI/hpWNmjU0LMdGmnHe
BQKi5M3MOsJV+l41GhWx81GPe5zpihnFEn5uWRo4uGcdzV/YZQmCxaVJiXAgItPQ
6/dPl6Ixkj/R5KuDcizPHlq1ZuETHll4flMng3r8cJqIlcRonOoatvMrnqO3laOo
9dGAxz1KvvhB4+8PwBidhWYjcH81V8kKbP9GuEUPvT6p3woDQJtbwgym2l7JW0tl
6+9zHKbLkp13rNDoDcijsEMZ7+88mouEeWjzUQ1E74WAZCOIypd0AUSjbfIF1IVY
jRTGGvf4rgeAsC8dELauzvonPQky2oKbupS1TqpZJFurDv1b1qNbIRzNU0Dv/t8/
JE0R4lah+mPt2F64vF5DPfJdngmamoxUMmGfTnA9RTIBVlKySiDp7imSUM78hbMR
dmAkw/NJ/f+0fLAHO8xthWJVbonykBcUBjc5/5H9WROuRaUWZf/X2zR8jdp9crLg
ItdAD4QyHfq3QqH9GvzItycEq5nnDbV9KTVnt/0Za7jCLk6YMmD8OB+8BGp8ywuN
ncix4kmRtC8MiTrPPJnu/M/xp56OIS2i31Ls2EpFC93n3zcxRSgzXx0w3EnCZDZD
FsZk4HB5Z+B4ZqjNKtZJqO5TDanwxpOV9KmerWXSVQv/fFHNSMReLdeKRsSmh8Lp
ms+zH4ymU/KQd/wrgy/epzy6eEhStNOO4pMZZWkwPYbuJ/6/M/v0gLdadHS0jkak
1I+1U24nFRNtmIFyrxk7oFvR3/KWDumbnmDc+QWuiD22796uDn9ugklqi917BgOD
7vcNV72KNFk9mi9NXYNiTk4jhwVWJz7q2fdLsyzOR1HBc67Mz3K42rk6GPzAwASP
wjqTc2YRU4FvsypMCBq+p8oihhFlN6kO5vKtkc7xNTAjI4PAMdiAFIemOJQZl1qI
QtdNCfu4hV3fQGeTsgjmGmf0pr4qiCHEt+A8GwwVPIUuCVt6muDwo/ocdMpGNioc
w4/ffvB0/EKWSG2r5Ph8+T9orv9Td7yqqyoR11r4wGxs1XgIfDZ7rMgy9RdS/g8Z
7i8GF2u8OQJMRH7MmwoV5XNbZW+k1Bqy2ng4hpT5GSMn3Qdj44SNahr4lEwc9+ME
DyM5zxBy2OlFKqm19kr0zWsfjFdmhgMVv7LE9to3unsA7q2DxiyCAymhLeRnBxFK
ILdAF2OEGTb/AI9SEzBYNtJpxd0Zkh+GLCYwPJAKRjFl0tCDM5isHFr/bp6LfSyz
9gWcJsy7S2TQg9Jy4aB79H6pGDbAomTv+XIPbNZ5rDkQJxTnnoFhnEu4kNC45sIy
uUHdHEd4oRT/FCsxIbrblNof403u+LK5j3RezzJ0Bz5Zil8NNaHre9p0Mhtw4kpC
30KmGXlEYEjy4ciBg3FHwXIYIHiddj3RA/xuIEF1Pamds06/INpnggvkuzGf7Ceg
YIejij1jorR2eOpAmFe+G60Dr1T/V8AbqmQv6p1uS48/xVF4TKmmp60VLAQ8Iekb
ZmfFOJsJ+uogZJY4oZ+vSWEhy6cs1v/WjId0nHWdGhLNnBOgcxtzLsQC2XMhl2Ew
roYRQ48S3zQiAersiMyUnEelDkpLZMKG0zY3HL0WMhqFTU2yhzsKxKHQjTLehaF2
MuNm+BzAniLlYw+eF12+R7Jemi87VWkH3NLyq3iWKU3mPqkGaH38yekQdLkMp94L
9tO8gh1gJXXv9zw97DvqC9DQ3sWtnhMz1qwENPw+ssjFHmdJULgNaUzWgRDKHhYN
GqQ1iAu+TKfIVcmY7zaALStFHIsXPRJnfLKoA+YEJcEoRAGj207QVA6pttYWUHWo
hHjzL7IE7Nf6IA6sAn9tB37ZqoWL82V496eho8fLYDTnwdqdMHc2Hf9laQUEqZii
g32h5z3DBcw+8RzdYWOISqQlDsyUqNu90SztFZqZc4/HMf5awUxIkbsXt82Jekt0
LulTUG3XyThev+FLt8czvdSozBfB7OH66/hNerdUhwmvNCXRSm/pooU4okyGQXX4
ny1htzA+E/fjVX3FotiwAW1bclJCMkbYRgIMttEsMRj88L1vkK1BZA8If0qCqDdt
szTF4LaQhFL1PEHMelOStN5lUCnIMbe9nCqhLzfBrY/rFWcl62EXxCtjvjuMlbNT
xLKBuLWDryBRiRuCaJKJYyE0TmswonzNq5QPmiOAwid6ZzWwflYpN0JS9mm7AOgI
saIBdyZlV7Q5v0WBrYkZmhy/1vgZEsmSqlECfGWv/8fViG5E7qA/0ZBIOszoemXk
5nIl9mbnRTXnJegTdikjPHOIFCEq0qm+wRVv5gitohWw17cjcstd2wT9XuJhrZUz
o816Hk51b9Opj3Hpd3N1dQvLhi3WtrdPEtt9lE3JNrIduavannIgRx8eqQ1VXIod
ye1dUtbkiKn2CazNuLfgAOYWGcOOhO1HLe/0Zoq3NWIESm2MbuURDQcA8+orYE1+
akq3CzC6oP8Y3L03lNXFFitN+Ky0yTQbeXYNfbih9QuDvSnKN/FLWx5yWZmbvDU7
j5z5B68GHANdS+c+XUKBMiPMNNQW14umKTkvemZHyQYL6327JS1sC+3+t8MJw8Kh
wO6DEip0NxCXXBTRH+hqrJ6zoiqcWyb/4nYoqC01izENu9H67Y0oex5YaqolNMUY
VZslBx50q2FD6BeEsV65KnQVb67RTa2Bbj17l4mRy22BnMG2J0Oyirnd/Z0p1EOj
hI5pcf7D0WmLNHlXBU6FNOfdiHkOGP3Zlo2O48PCLuBqSe74Fuqass1cCYhq9h2p
kmXwfkoh9jpJ5h4dsFKj3NPj/OOnMGmmpUPws3SfaFm5EzfkVBmBq9abLKDDyhuw
HqPHTgfKDytC6Dty13R9GwIq6he6T8jS0VCZ0GscB951Tjqk4BK+Mk+XWgdzHKzJ
mpN8S8zJKHUXdQQFqlS7XRyJkWM60+pRWV7CrxG6lKitwblWAClqLiROsGCSEi4Q
+58yfg68afD7UHECZfdXm8S8uA+fChm2oy0MTxDsMS8mcpFkBd9zrQngMCfl5+Kd
WsSepOmEoUR0o7Z5D+DjdXkjEEKp7ErV6TegtJBH9ViTbHxLEq1t4tx7bkCdku+w
Q48C+icfwZv15cO8oG0xsacV8P+laitzvhSaMErETGqx8EOu//ebqpKAW7rgn1rd
6il06IU5u1Kk2U1Pca1lh8/EPcehcQiZA+gHgDFe2C7dIzZDSkFAFx4Hh88d5SH6
TUchBGQ/5gNdtYzWYIPiXMIINUaPZ3GtSorVsdNgShUWiCs2f14p3yT3ZlByJoMA
T8LQdAVgq+3vIgx6LrAzSFepl4qGxMVhvHfQXW1jJuBcEAtHutPwNwv/NVLWOD1a
PrMZfR/D81M7+yto3Le4Ch2eoEtRpzl5sNz3WAk/+NrB4LxjsI7uoCl78Hn8rJLk
/q3p8ypGsy007i/7jgAtmm4P2kgSUH4ocaLoCJKjCBY+bny7ABZdQhuWqtDWAhNG
tvEwXeRR+8xA/OVPCZYew151D02YO02UtgLulBeEfvU+QxSXcLoLLE311RKaJDxf
eCml2Zw4mJxfrnJrGJsTYHc6BcTbDFbg1sT6HzZWuv8eZNE9y2AhApER1LsXs7XF
qKRWLo2P2siRV2tGI9V0f6kGgD4b+1mKlsbPJTTZswo5fZfnlb9tHARcMzknmY9K
QJtrKSzdyD+l0tJXSealtKnz3XhtXk0bSNR2Vqckob+tiSNsokd96metyIxEpQqh
94zpyL7wEdegYe6Ev5crOnwEtMupaVDWXPHJHGY0P0sl949fVF2aQyQK3BEiwD3g
DBy83X5vWHKeJ0gwCUqPG5C/ffkQsjcZf+IqddmMqglY6/+/w/WRKrGbUaQ+yMfr
E1mqKVJCWvh5/EHP6VRkMtPAg5VnCLJVMoSri54HFPtYKaFR25CsaNnrRIWxyBEB
nuAkLRqhDii5lHiUv0nNRzCiz4umTi8wN6AJ9adD57rrqoutcS3zvMVey6FU/hBJ
n5OlmfqFsFCjOJd22hEX3rkFGDE1tk6jwtRkac/twGjPVm7Cg0gtr7uu6rmnlwQI
73e3QnOYGC2ztzKnySO6vrddz8oI2s/ptMU0Y5PilHKTZ22ILITwW2DOSUEPjw2o
A3TcntcYx4KjmwDwqONJy9NiRzclE8C8/O8sK2a7pewShcIL87oc9neWwEgh1Dds
gLf32Ku97mmaLDCIStrZrvnIFKAeOaariH+jvr6z5OPmAdSFWvEFtjLuKAaDKU13
ETz/GFQbsJIljohGD4xt0KEdya7PRuLPiGGgwhLlcSFlM0WF1pGvGtLHBVN4ikrc
lOMfKrr77kBtizvWXQx9cXXgsuq+NLsu+5iUe6y33TZgP/wAk0cONd6QpS+msm0A
gCC8ax3wnil1CA29beFtgGTMGszyb71xgMgaOFek0+9M5BYkcb2PJ5QBNDXE4G2H
q0rRzm94HcJNUIsMuLyRbbaqrhxx7DVZc+NCZySSl+wjQTEAVDUYUgcE2iyunrhI
9mFsD4njbCoRQ/kzcVsDV0l61rOP52hlm671kPKi67R02d0uT9KYKl+GvTFls7Af
9NOa6IYCGX/r1one1DsOK7zCV2FB7wCCupmDiiXWUTUGmKTbg1fLd3Y3POjsVY51
sm6QZuNPX/gMn6H2M229etnOGh7RyMOWg7cGN8GvdYGBXw/uAc1NueOoKpk2vjLn
ziAKxGcTGsy+MjAlUXo/WvoeqORnWXPa4OY6LGINpdX04YvM/H4cxJ26RdIrKNsP
1lX4+EIupKLDneGBirDoHvgd/A1cu4ETyJHdNrpqvPVUG8mMV+Q6wIsKQte4J9NQ
dLFqjcniFBNzim7Cure9MaRjbxL2NcGtQE9j5+4d+VqsON0gC02+vRS1e1aB5kVW
zicWtqhCTFfG6OpvAoaGIERX2GN6h21Amx3cTdt68XbRacbzvA3n9eJ5UWwPkT4P
nxy7h1buiPxi1vh5gfhnwUJnfzMvJMpk510Ti2ffpy9MuBQzHZjZyzM8L738Inmw
JSogsPMlBN/VC6y0MgTmXRswQtTAvhsKxYQmZp+lJfkCbqAjmXE9FKTIGF4jeXEl
JkLNzfWj8om074dbNkUqhAeJKpvHhZ2BnJI5bpllM8UROQ2OlgksMBc9nJUH0bJ5
sAWoEPXpGldxZBW7Vlu8uDY/NQPYm7TyU8l122VH6jtHW8vH6wnpRDzZinw+z+BH
vpaeIZOqUwKkN4ybmwjpP3QLghHA6+MfRrQogdFIq3LriiDZM+FSqeaPxXlMAPNB
iLS3sn+b5ak7v5cs7E4xF8RZ9szjCS2uWLhy6xGIlT23ZgkWD0UsISyWcIBQcvvf
E0gucjwDYkvBXESIvg8i3TOoGu+RWe/yVNCuBLDQv0BvovOmN2Q9TrosN8AXOX6F
EDCg579rodPpVsFOruJ9Xs4RRm2B8d67r7ilaqDpk28n00evTSAjlOFA+/uaXpL4
fwzWiYlxiUeJoyBQyx/sx3uxc6+kuRJ4F/Es57r17FTf6Wp7BoJeXUEW9hLt8W3m
/83Qrjq+U3o0EJniJSigyMJ3GtYJM+gT/RZcdKn63NaXGF4OeKdDdb/7HHZYKceW
7lCnBuJHowoqTTD1BJ6mFNUYpTVLCIOjSxqlqidA9bBxiKGtbd1Gw0aT7T/F6tmr
gBQUOQYMMWfNbdSpYrKLiwhUUA3LabilVkeWAkNtaugVIZ271b9JTvl315HYCcB9
bQwrWr/EFS5bIskd1KNYqXsG7Z62zQcvppxNksop2F2a5odZyZU3jVQ2hpnxuDip
Ed83b6IlbSNydD86gEG3rwdAahU04l9i3LypkW+xcOG4jNQT6IoJrGBnzzs/j0Wu
0CpSPuMuDB+Zlq1d5xRjNVvi39aWHUDvjsarhXRUMIJHfFt0pk6fhg5wd0zy7aMV
n8b0bLmY08Yk9RxWt4Hka9Ie/tDiQYSR5PYtpZUPeZV3w+u9YtfuWSgkkVrhot9r
n9iiYwUMurS2ZGid4h+bOpedoUT/5LGojJZBn2hNAYN62V9jGEvMSSBBMcHlBd4H
g5nLwH618iVDaBPc5NdYHzZXijKUzIULxllSmXyd/j9DzHJ+NLPJs1g3KrNsP2cm
MelWbIyCJZCcszrw1zzxrn6oxlmemX/jc9fnjvO/D8SQP9x2D5U+Uxg0FYvI7Gld
lWc7GNQrNAXHZs56EA03TS03hIPTaoG1qiNp7qRhqSe2DLR+diJvaKyHOyODpBMU
AGm0fR+NzqMe+MglLVQDh9glvuukG1Z1Cbvde21tWJrjx3GVWGBdPcRSQd0k+8bY
CQ1Nl/MV1XAOr4F0W0h/0MKvyzvfAy/+atiezlgsb1wepLfv4W04UNcVqXty4CP0
yNKGzDqTSZtzmxXXEGFx8tASjYfoKLPAPFB2bYK7yDe4+f6mKfiV9iVqbEKOoLGd
i/L1Ch+fzwbOFqd9bNmtXutePr5J79+wgT1uI1O66Yts+8a7T2/hMp98s9bzd8+d
OiXGkjFP93+bA8UfMIKZ8nKg6sE9O95O9Ym57tVNSOHr4C2RfwL4LPC9YerfdMgf
c89UMRjVhvY8X4FImUikhp6t3afW764/8/cf/8o4QhkIuJ6KGFWYT3981nVD3KXK
LLIblZnZyr17JkljF/nwOsYTrWvzB3Ixt8vNMcC1LDiYPeWBM7PCWcH0ar4QoL3U
Dnd4+qhZky3UJ2sJ2tZr54zYCvucn7DOjqm2HT0KecY6XiVwkzMHKCzSmNXPH6vl
fY2sqZkeNBwy+v+OwIMcSXfyFdx94PnGVYe/eOQ1wd1IbIEzm9e6etC/p0rxkVWI
ttO4aeiO383XDzUzJsXp5vxqnyy42n9g8diYtA/4btS2gGk6WPdyUlEdUvUCZbsW
numO5Hj6iEcGswYEv7CV958d28XDZrewgVY/6IVZP+S3Uc6FUXUgyh6/udS1Wxg+
XAu7LAyTht+Q2Q373/OF+GVIecdRe9KyUFUPdp/Yn550urX6AN2yn4HSvAg1MePK
/W4cdBzTxoFavuWJZxObm1hIsC6VjZkD7+QwcSJH6Il5TGMeFedBr54aKVTtMpG5
jYHWWwCeOkpAvVF9Qc6QI9t0sy0ZljB1AypHTbr3LH+dpB+hN5CyC+UFf/YD7FX3
Qwe4JqXqkg7z8f6IL/cOgkk5bONpa7W+WZYfgtcB0/u3oa9o8ul4nrSpNi+IkrAo
iQeZNGvj3EfUJYgVQfvSPvxdeid6MmfSf4XmPcyeHSBM+HQIZuKWTrxOMf9EP+/R
RF8pAMl6S+C3Tei2hzdzhOt0bg5mK/jggbV2N6vIlhXQrQL5iqCMhhjgEV9Jtx+U
VIoKDbAmBEqKs9h8WyOltns54tSTPNWrjLxR83b0mTNhQZlS+DQ3B3YcY/BeNTZC
m03a6HZm7q7UhHQxyvQ9hWW1vtKeZ0TcC/F76qs5Ss4mch8k3VRG5VOrjBcYUM18
jUUqK+pIf2jSn6M6gusEaNKW9xybusTAtNTwJICdhP6Dai9C0QcOJ106yJ9RVxR4
r0RL3C+a3Ukmh1NIhmzhEzCzPg26V807UQS6KXfCDxxgl20/F1fwLEy6hHT98Ibk
OE4lKnvfrfk8+Gdg17HHtf0+7Busc/rnZaG7mjHP1Rt8UCFJC1g2/v1hXLwqv9CL
rDRoxygP7cErTFRhv28ab/0tp/aTSvkNfPVP6QGhxjun8DGzf1ln5oHHO2EcOAyq
KKXTSboPfZdkq7C2eibOCninnxmVRUxYCkuwYTxJIp9rzh/dwAR1Gvq5Z0Ay2dL/
xO4cERjOEIQhgpVxts59cBxts9EMYXDdLGN0N3GIhz2QAkmgVVfttnZsLdx+RSaO
qetTybf7VgC1icPZDb2sT2FaHY+hK99/iiHP4uT5qWfcd8z/WRALwR0nDuGm5Uxm
JCCCSZyj2noNY3BoyQR44St1XWDzccZI+jWbHVLpZChNO2UJLgRQsqcpkCVp+jH7
c0I+rlvKKpMrs9762SIhfRwpiRdOzmpUu36/XVpUaUrOsJzEhGoYjDtjliETGeNK
fCGCwpNm01cxuVIay6AblILrONHdq5HypMOb6kkU+CiCNw+MXBaklVFU4Z00PuIl
KZqXyfbihVSCo6VmviNl6hqTrpQT4L1wug3ok/PPSWWo6XLuhKE8wOFL8k4+JcHD
VOcn93rCTzMDAOOeKEOqGUkixvuOSoZ1oNbw+9fTuK3GgTsNdEU102VHfDH9l0ML
5AU9kgxkiXx7XH/eQ0x7N1cpZRlWTdIwSB4XE3pOeRFkF/YE4RkQ/GVfIpRXP3gv
wslZxaPhBVhT9xofeOESorVOsGGr0Yhvopg9+IXxDSbT68fN5vWyIUseiSfK7Njc
S4msqKBXV3jX4xcZ3XH6C30SH2OWnrUK0BTgR0y4IxLnR7d1mjQA0CmaQuqx6e8x
hWemT7n6VW1mAXui3GoHs4ruv0HY01iUuS7mXzUB+01yO0RVrxK7dQ3B2yE6xEY0
qSHtvOYJz6CMpG5IXoF4OOpDR+zFtGGLc26UoPKXp0VdmlPbj4hWy/WbEpB15gxy
W4BbG6+IdpDBR3tHIlgBTVFYmNQEw4dOOkBSgSF6sRoUFBi8PL72OJvcM9LC+Ue4
9UdakzTaeqtmipnDY/Ed7Czn3nxTh3SN0J5wgUVaz1G63Fn9kSQwDt9JE7u4U127
7HvVHtZyEvxVwQzHvRsyZXnUjM+Gdj8fw7ZvDMnHgOAab+8y6R5cLrB4scYvLvjg
IOVQl17B6vTeb/o7qEydFeHjDL3lc8n6w1e/Vgq4TAvjDUl8G93Zw+79eJmMbXV7
QXtnKdhDTkb9HQK+mPupt6SVOBdHXi8UbSVR/gNOKIlUl6Hp514MiKSBorh2sXVu
OoSCUy7A0cdJwSjC4XEvZfjSWGlTTZHtTy7xvEV23HExQl3x+ajX66nS1KxGxTHK
bAhupnQELXzNqzUnworpoZ/S9OHdRTn1H+FKh0ayCyJep0YvmfVW4mNiqcrYChR5
FEicD+4MBFqz/Kb/UkhxUKBvZO6tGDI4VuZkpuvNQI2HRN84TxXvpX7m0SpYJcY8
rxobmLCWHCyTw28kL3EFXCAbxVkoI6DlmBbqPfSSxCreh+q23gNnqDBkkEzR3BdQ
MgyM8ikWYUX4j56XZ1f3+rroS+nDQkktS64sNM3cj8XqKYpAmwO/arUrvBBwcqA9
2ywblTqm9mbGWW2FHd/tDbmKL3s1G5+JpdSE6Ln0kyYOjtGWafp8yP7STCOENWet
8Im0YJwSvGmBV3V3Q/mLaN2LUvo40/3UaEQ6kNy/qxSFzuy0SUg+chEHeBnS6VgT
Gn0f+hNYSLa/LoYM5wvDXTS48C4HlQDbU1YK8MiAEfzhCWIUcsTfDGuEspr0efId
kiqpFI+ppAq8mKehzSlsMPt4KQvOgV5wV7WA5eChRpCN5BYLyGPpVsCAaiwJwqL+
QRH91pLUcP2uudmiFofEHKPLEeeEOHZl7S4g1CyddcfWepyVpkt0dzmrikeKY7WG
KfaN85/bqRnzRr44KmI7T5NUwOrKDpFAyIpCQgT/ovrYJeoTVidnPMTZrEv2yy7O
VcwOh8eYQL/F3LBRzgoV+RfkXgNIf7XawlNbyKTnKW6GbKiBl1fN/6G7wFebmt8d
t1VUwDcC4RU9hbFWJ0RYoGqcT6ESEkSSGpsPTv4FvRc4YFpXE9n6HCEifDHz+NSz
JIg0nfYScBfpsK+iXtrX1hxH6oDkLUDn6SPdCSfKAzh0WLQn2qQbG5llc9drqtoQ
vUWXr2NurxIFhJthUnvlDX2y1HnEA8RRt06vElgTTEZ9pesHo+qvNlDxoGaRJi4Q
DA9oJYVJYPPJMx6OnvZN4TRAYJ9mCe4h/7D5a7te9oQIl6XbuGl8ZeHEisJqDcPI
ybOFx6bpJlnCls8yug9CrPubIJyJLmv0TNpm/nO4+uBUQy1wQIzHg878qyQrVbQP
Eqh01Xk4KHjOythtzeOtFRoOl+FsciZXlIAt8UG6+mVNaDJrdy9dMYR3PE1VFp0O
m0HLnDIptv39mdytN2iPNNNHlEtESR9nkwqzKsb/sA8Giw6VikJpusHtpzjuhlTI
Dk8zeoYWjssFoGP4O4sp+JVKvgMfPEMctRH00mRxORvM5cVzO8rhzFsFELLgJOiD
dnn8NWhaKNhbjWNOQnCYDjP7Bm0L+/5qERjpp9+V828dvJeRpghnsGL2PzuidSCo
EvIPJuULoiOQG8SYO5tyuBT1SZ9F5qT1sm+9x+ONboedI34tkkBPHIdxJ6KCqDki
QKrKbG74CISZBJo5N2Ek3dWFdqAIvdGUy4jbrdp7wMG0HBWjJv2sZ+3ln0tzA43x
fdqlcVgICtAnXf293YqWStsSzKDbm1zrxWgxa3HfTdhP7WvNw0ccMTe+ESOHeevV
fRxm+nQoqybv7V1X8Xqf9G0wGx30/KjzhFZPvkTC/QLYxpXIIJazFE0eDCQm6tDG
piITQAEKmmAzB2pFmPnJczb3kTRng1GXjSaCUBlLOF5/SlTxIYVf4Csee6KXXlcu
lkrfkbCJbMCH1FvDcr3NeHiOWwzDyeL3flN+VWcvPc7tQJQ+ddjvqsRslH5vF7qs
kT6Fmx/LWf4FhByJDqm1oBPGE9qa2qisYBYJj8f3Nn8qEAL3T1gjWlyjWv+nF0ox
585DhJXbcJW8rSkeONJKIuR0gaErUvFy5BWxQO2TeAjhpgUAqcr6PAC5XMt0mERz
qRhG+MKPG5qOVuVr6RkTNyH0Qcm81kkfFi7YlANuoN2iB8QJjlyVeeIlqf5mOTJO
/9BgWOVf8huMUoRrlkcAZ8dcqoSndGn0lAhBKN61clCofC5TLCBCcH54G7t1gHbP
tNnizbTW+Vxe+b18cs93rxmxlnYFEFsq6KI5brm0D2GVRLy5QTARb8/tGm+YYU8n
eubI/kB1FiXFzP4UHetyPKGRXlvbaLnwIPn3mnmIKgAkgt+2XxP0oIUrrCEzMBp0
eto1H3IHC6TsAbGQd4X1zolAcYLJIbu68CI3CKm5rFQQk3KGwW0TVScZKtIQCSL2
or5p/gow587Vx069pCyjphOw2eykoTYcWT1RXDCnn5o1IwZcXyMiUfaMj5XCd05/
+jzH/PtYEyHj6Njqpk5SmtcXc9ew0NlQOnOGabkRlEM6fy/2BziEtxPEGkEAbKk/
Mp4f96qyo4IzXF0kUrT01zOIJKDcbo6EsfrmCwQO6OixWJxlJvNtke4VHSZ16BMu
9gPZ4CnnluQbHn62kMLP2ZyDzztxbygYRmw0wJl8S1WnFWobLejdVaidlWhhFKtb
NsiSK+puwMP4oe9XgsWe7ky5EVrm7HYZoPxgQPEVNj9090XdOcNmFefkGH+3kuBJ
39Sr28wGEft/DEkX/FsmZuwTS5Pcqc+c0XHA2ViX5qQFhz78O9QTDcTqM2V0zB3i
iiy60IlByniAqLEmElGrJImLvj4JWp+FgZval6nI7nXsexOgc4ZWaD5SoLW75BWU
IXnsIogFvDn/y+RUyWwJ1TKeTh3jwFcS1CiybBcXCIDPmusH33aUEC30p/ySbFEF
hovK0MWPkL6ycNoTbaHgKBi+bKyvblA/CtSfmKw/jQpZcwUN41popn8Unv+yGTR+
HbPVJhSbL3EKaLzBhmsyM9FFgI0jaq3bGxbiPgyMIh3cZYJKIrqBCmkud9DGBFG8
6uYoigabfiO8bEUzHIsi6IyNukDQojTYf4Z/NJ5Ohm8gcknoUDjF6Oc6FHJjZ6Gx
OQtkEkeNpafvYqSjXq7MYJP3UONcCoFCUhz0x1IG5Ui6UC7+ji6eFhr2uVM+7Nfk
+jn0ZtquqWC8d8afz5KpQiPDPyGtVTd+TIcgOFVcCkNaSOXrC5DBMNIVBCeC2Tr6
/IXLfeoXAHSwOz8BhnMn5KQ8vq4i4f8vqK4mnGEbnjZ/OnpsZcmOmkab2qNb6JKw
z91rPEtxPwgunG5uhX6cQPnZc4iO+ldgd+Ak/2cc5oda27EAW0HdyfEnr3bSTpZW
+985XnttP0Dg8hba7+8cQRqiY5FqZhyP84EJ49abo1JEAr8WtMzaSc2P6vEBXKLs
B8ng/9NhBLI263dJQK+gwRuBzhcgFWNZGxUqaewcfqMJRf6mnVorgpcm+1ITH549
NF8SAy3If1Q96tYq2Le1l+iPSyrOR+HFZmulD3RWCwl/rOw/8wPG0VE6vq3Fip9h
yFdYzgOiUJF3RhvUHOX6Z2e79Q1rS6Cz3nOmFcI77ctwoyZsHffTCr1nHDorDqqI
821z3llW13HBJs4w8NrbEnf//2BXcZMhtQrto3E4fzqLaTKT7cCBrixXKQevAn2f
BsBeyPeTf8vtuWca5Afu5KNRAEQ3OovTN89FVXx7sVI95G3mTuvP/Og/6et02+8W
QniXfXg1o3gKt4PTwwenfeirdZ346OSAUgcIpz6VnA4gxWWjJ0/HnCnA2HxmSKG+
mGO/h8MOQYIPQCmGt5gKe7fQ3a3myn/Y6uFWMgZvhoV3xUirfGvqbHLaHEY4fk5G
bS0KYVi0c/JFUbheSdzYOQbIUXTeFSc7vkZZRdX30K/qx+c52kqQ/9R224k3DCEo
mW5SMvJ0gNE4MT4m2AAc+25V9zFw+d3umbdrjyQ5RxVgQKWy0Qp18r9ybpi56tya
bIJJYOcXYT5VdFM3utOeJNAhftnEwzEtjt1B2HzfzOEobDFP9pSFHlwQbi+uLtZd
4Q/Wd6Mrw1Q/5xelfIqrR2C0ro00VnSly31hUJjr5vVwe+seo2hLRofC+3MK59/k
5XEFmf2OIuIVsEh5I43ThAii2RLsQSMnglXfHthDEYokSyLKpoIe7LELBA7/fsCQ
eIxA7w4QS0I2sWBNf3Jgo5ADyPNc8ZXfxVPZYgggTcCsB8Y3EVucjTNy4g+yc+k8
yfkexuLW2sUHzaZ+byi2YQDZ5cCV+KGEBfz4Z7ntylD2bHDZDByaGP7im5qnhe+0
pxrTnvMEJDUCQvXeQnchNB9je4p5yzo+fdeK1EvTVADOdRH3am38pfuW5Yx7mNex
QaJQEkFza0K6varyJbo+TXPHm4EffaupVCPb7TZ5pRdrtw/RZ1QwsSzX1m0ZBBVh
SZTyurSKt7/8LKcuVdu761qDXwTbSZQjhZ+4GiAzANZ2trrTF2aVUa3pCwPbNt24
WQHMB9boUGLYDFHB3gOn4UvN8rYCZ5nUp4lm3YhaGax0mociVOHy/rxAMWCychdC
Wbk0t1J+sy2zPaMSYcG2K69wIJ2FoFlMbaQWNO4W2OrQEHyIIVd1GeU3w2g0ShmZ
TEajUCtRDAa3V4EN0LnO4BomHXp3BDQeZ86nneR50aKLWFshRbuvRdsVxZNuiioh
FrebgkXkF8OHsuWwyoQuEhCiwIfkNwvOf1c+rgLeJdNIJBMbqN0gzip2pWtsYXmt
vQkftjyeXZRfqB1mYZzDvWEVXmV9Fb4KxwSf91s/akJg7uJj+PEbZzlBjRpvsfBU
F/9rR/EaSuNkACZWl1c2G+kQ3sck+FGPa3147QWLBcZI73aK5u5MyBEzdrv9N9Lz
4+PJntHKvlslzwduAFhqapXAtNTvnzO2/5EjiY6Sd/O3s5q4E1YC7koNqhzz+GOW
dPwt02N9sduGJp2e8lP5vqT/zxtoUVlwoSdULTBSaRBEMFP2/wUHNmkDvghCXdG4
Jq4RRwCOxYb444xunUVbj55df71/KRRV29MoRyXr2+qDjLdlo77Pk7AWHsWzrtVC
Wq9oXOXjXjj+FkVSAnInI/83GcgcWFcroFZvBouosjVs0hlDcDrnoiGSla7KNXuf
NgOA1K5y+BfvL1YbjCRs+U2onyrrkvGBdYGIkiaIEAX7RmlzVoLMS1yMV4k6OOPX
RLuXiS/Wj+J8qMpjLf3uHnQcf93WSknRQ/Av8aWKEK+l+mep7PX+I9DKZKZL1jkk
D+T9GMz+mAffjU2KZRUHoFmoaESCFxSsxuONDSqstGC3UMWxT0P1c18E7+Qrb4Po
WvPR8DvlQqSIYQLzGiOCsS7CDTkJQw99tHT18lTVaVxsbp2dVAUWF9fmYDS9kNSX
zNNoLGFTYsVWT1qLXaGdLHWcdbiSQCaLYxacPrRwOsGE/KE82fgbxwmoRUYedEPd
m+vQ87aRNmPZ63GE7YlzU3XzB1Xo9OwkldBbaMtYhIYXnh+vNdryr3kMs1pSonXZ
CmczswA0x04YbEeeBubRFBZNPr/ATBGb+VSIqUdk457FNkE6aptGOfdNMOR8vPn5
F7s8gpoNqilTw/2j9v140AKg1Urp2vb8FMeHOF4b9Hx+g+lSq4kjE54JAWI4JopP
ETlleQvHBCJZ/Mlt1ImQT5pJRKL/B5a7TejSsJpLhQ+HN9pxfCz1Ojh4hFec96So
PofHjb82tnho/oYG4zglrdQsAZK9K7JCX9cTl+7UHR0XHk93zlivsUCoFDibYKzq
KqGdxzrjgOIwReAQeM/QiSJp/uNtYN+loRNfwNI2+tj0pWx6QMGEfk1YdkVmuJLB
DJjeAi8Tv+QmRguRGkqHBehOgxRmaipd8Uth/CuDuCc=
//pragma protect end_data_block
//pragma protect digest_block
0TMBYlaJGEGVXqBcZTecWq1/w54=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DhSjbLqGkx9oySlh1iX/VNbModukUpZHxvwoeKEYFDQ7hwyWmkCczpSgWH8zVVxO
q/dn+CXtaHfqk3VnRLB5VBmh0W7UVKbnT5sUWMNhINpVbbursNpOw/vL15l0h0J8
N/Q/UnU29EnxzKcOT+5NdULLJHYeW/9KNaE2qKWPcktetpdtov2W4w==
//pragma protect end_key_block
//pragma protect digest_block
/ymmBCt/7EwHn1+6G9iTirY6LBk=
//pragma protect end_digest_block
//pragma protect data_block
e5uvugnipy/z+jtTmFOFklehJWa1JVpKKuP/KqNcL1JXyJqALvcMRHRf6Es4ps2Q
1vlThOr3JWwXRRjT69kvqOUbAbNkliPyC781AX0ylBaKuXL/mHza0FLdbu/Am5bV
ESEMNdTEyQfSMz3EG1CcxS6vyzyjWDHVJxQlzzC7s8ROnFI5yPCupaLga6wpzJjR
3yQbqeyooyYYvKm6prx26q/nZYjyiNYM+bn2HW2RwpuwErAgW4bjczMlnRphZ1SW
D1Rct4cjbeh22yqrCy7SJ2m8wIqV8zQpJLfOPYyBeFxE7onvGnvoLJEZWpQ1gEzA
acI1k8gzqFttAuO5FXt+FW1o84SO+9f0rpzHW1i3SmllW8BCeRLAvMcCHU3/tC2r
jlDSjtY3UvCFMtACPH1P5w==
//pragma protect end_data_block
//pragma protect digest_block
5sklou08Jh5Runq1GICAUU+b4hs=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5C0tyWOa00PkHu1VtXdF/n0V8qpIPVmDKim7jiEBuvYHac9pzOZuX6hnKfjCsGVy
CyiY4Dy4yApZEVaEdRbL/l+qV3Xtn7zjKG3rV9qv5RShEiLh2FIchEcLpBfVacoU
I9ZWjTBZOspk7sF8moEjzaLxXNfYPvAUplrFMLnyMV3uWup2S1YUAQ==
//pragma protect end_key_block
//pragma protect digest_block
SEJGxPQFT8IaMCE9acrPCkw5MSw=
//pragma protect end_digest_block
//pragma protect data_block
UsuDT2ffuvl1kTv8d1Hj4h2IqkYx22ykeeMaQ3Xdnnac+qUkb0JC0aszdwoDEGc9
U9fT/KG4rSWEDuhAvcbiUvmeKQABFV0vzD9bDzRIHj0J9iLQnIE77ruRlVLBnwAT
C3aHg418jviGiiwLGC7JiwJ36K9NCwbcDpBKegk6iMl6TO7wdZsuLqxnxbii7CCa
e8AXspTBecdeT2Z8Uxu02Wz/mPfLdl8/MwddEawk4oTa9+U9NbH/6oueza54koWX
rNN/OPQwZ4c42hOhQcuEdho2EJ99lSiUL0QTwhUmtNWDKg+aJEYccjaKUQlia2Dm
diklyylgWLTFbg+zLqP/83UZVsq5j1m2t6QsVDC0e4LrMNZ733a7OBAFAW6FA9Op
xPq0eRYwpSqiVtofb1Zvyn77zMkixQfLhApxhLZTtT8QJvFjzPlQIyTUI/g9D6NO
GqEPxHRnNKdlo7tbmXCGul3XEO4ZgJdnFcNuAMzq93Jz8zBvOwtGLxqYOibNiUyT
a3wiZR6AGecDK4GuBatmk5l9wUQb+3CcYZix0CH8FrmYt8LKxuZny3HgWIGYrX8I
t1jMYO5FAyUnVLW0jr41Uc9+PUmsORGpCElyNOPLfo2GGjtg65+e8GHYmTihZeu7
+ZDvCac4oa/oHFs/vQRXRuhIme3Rc5HxaAD1zhuBcmSmoThDZkidspF0a4dbRHmx
sLOyyr+j25Dy9sX6TSBeEsapAQqyCZUeXJjQ/JWbPZUF1vFpp+kYwLtWZ0vGBpJE
l61NwyjKX73Lijrss+fxA4BIgeKF3tuFfovLO2/0TsM2i4LL9Uu2MjuXTTuMDmBY
+uFgCpmjtghFwTI81fRCwlQLIuUkEDycmK2CowTqlen1nA/BN2ZlpnGsHexeyYKm
1XzWJLPNl80VjOpHmK3HD4TLMCAdklthf27BcdYF7Hlk9hsY7q9RgGVp6ytZHQIB
HcYOAcpRtMwNwkrg1bcjEU4lnnhJ6snWbsbsBi2iTy3F30Bn8NZJxE48cCuIsbQC
3hqv6pgXQhshNM6d++oEG3wiV/qT+7+cO8GRMbziKX0jfJmB/Jp0Lg54Bcuvh3Hy
pZ8wyMgzp2Vm6r6/8arb15xf+gI6spvKFOYEa92KdMHPI7Zv4WPt2l6nLLsc3AYW
jF2MlNflNb/YBhvKU5Fvq206f+Gn8nI3F+jPm8wF0l/3SMtFPuEJucyR+GOYbyZr
Ni5QK8vAwyLjXkSixPg5M+haN9g5IwRdtooK3CAnjppZPk/+gPFll5skMh2hvi0h
ef1blm1TQmefeHt0HzGS0AZWTS5Y8qYEjDJ49KrdhxLGJVpd32F6EOYvx2ZPlUap
VW7O+JFVMvlIdhCFrx7WA+BMeZUUAv1/JAzn6+YlS9Tr78lLIaVRoD4Rdu89K10l
OHg8ZBdq8fyhbpNsL0T8KZycJ0921RL1xMBfcx43Cf0RY2NMRXHrKuDuJyVsJvyT
q9Ov64c6F52W/pdD9YdvH6mvXbnAuctCt+u6DlEYXR1jHVar9IRsC9miepIEtaen
ORU08r+Bf+0KRd3FouCTj1yx8/K1ujurCyMzpZVOZPauS3fa8HM18TR2010k8+/C
QzCkTJa7o3bOsmbVJTmtAdOuWiG9oShlYVTSwbMvRj8nKEjGXPGiTrs01I7eJ1Ri
4TY7yb66bm3udpT9WDrfA2ZT9xduAuLY1DD2oDGFt604DaDfRfXfj5eo3jTbIdWw
z/sRaYYIWqd0VaSyC31YhCn7fX4onQL6HOZnhGD1GPoRMfW/6qug+GyJZq05mZSz
sjJHnEBgQJSBz4V4TEkS8OU/huyrbOohdWnn0F/Z2i3mR8ehYSnu3G9V6MrQMKBP
sTlGsBsm/VoSNFTKfYKZSCDzv7vI0gGl4jpx9Qjp3g6OV+J/2cEh9pKzZC/USle/
ZqYQ4h41IA6Iak6LAIhMCCQwSoXDOAfU1soK3mju8aRm9vttpzwnSggzUXAljdfC
8/NWkkxa2Sbyoml4vDzdoj0tpjfNrrOhVW1w9wBuCIJGnzQlOaYRHtGdjJIzdNm0
4mjaHC4LSsnuD0HVdrvp7xbrSmX3zogSXsnfx4uS2oaQ+A6//W2Ro66ALU7gnFQn
Ku4HwHa91221UPsyHGiPLsP9KNUNR1szL5wxTqOhtUx2gSuKDPzWcsxkGpvNqBAR
ynRCWnSpizJHQjdGKiukd/btw2ObWFiEKMbSZZ+litKMXzb5WLLRhXMJ6OUX8b5m
aTTxAGZ5swgGJ+lXmN2HEVwh7BL3vz/vM+igv3yIdZmHumQrczRz3chdxa6Ij340
2u8rYbEMvXv02q0PuBlPoz2tC4Ha4ZnUpOMXgsoWjE0bnYemT+UGd6wgJQoH/j26
ZeFO8vHIL4Uyhhr+nTXzgOD4YN3M1rnLCZJdJDInEnb1HIpJrdwMFC8SfAbgcECy
I1T17CrvR3qoyPCVvcJdSw==
//pragma protect end_data_block
//pragma protect digest_block
pAZw4zwFUHnVVP54RAUtt3d3Rjw=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_SLAVE_AGENT_SV

