
`ifndef GUARD_SVT_AXI_SYSTEM_MONITOR_OVM_SV
`define GUARD_SVT_AXI_SYSTEM_MONITOR_OVM_SV

typedef class svt_axi_system_monitor;
typedef class svt_axi_system_monitor_callback;
typedef class svt_axi_system_monitor_transaction_xml_callback;
typedef svt_callbacks#(svt_axi_system_monitor,svt_axi_system_monitor_callback) svt_axi_system_monitor_callback_pool;
// =============================================================================
/**
 * This class is OVM Monitor that implements an AXI system_checker component.
 * The system monitor observes transactions across the ports of a 
 * single interconnect and performs checks between the transactions of 
 * these ports. It does not perform port level checks which are done by the 
 * checkers of each master/slave agent connected to a port. In ACE, the 
 * system monitor correlates coherent transactions and the corresponding 
 * snoop transactions to perform checks. The checks in the system monitor 
 * are geared towards checking the proper working of an interconnect DUT. 
 * The current version of the system monitor requires that cache line sizes 
 * (svt_axi_port_configuration::cache_line_size) of the various master ports are the same.
 */
class svt_axi_system_monitor extends svt_monitor;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  /**
   * Port through which checker gets transactions initiated from master to IC
   */
  ovm_blocking_get_port#(svt_axi_transaction) mstr_to_ic_get_port;

  /**
   * Port through which checker gets transactions initiated from master to IC
   * These transactions are sampled from the scheduler within the Interconnect
   */
  ovm_blocking_get_port#(svt_axi_transaction) mstr_to_ic_scheduler_get_port;

  /**
   * Port through which checker gets transactions initiated from IC to slave 
   */
  ovm_blocking_get_port#(svt_axi_transaction) ic_to_slave_get_port;

  /**
   * Port through which checker gets snoop transactions initiated by interconnect 
   */
  ovm_blocking_get_port#(svt_axi_snoop_transaction) snoop_xact_get_port;


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Common features of AXI system_checker components */
  protected svt_axi_system_monitor_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_system_configuration cfg_snapshot;


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_axi_system_configuration cfg;

  /** A semaphore that helps to determine if add_to_active is currently blocked */ 
  local semaphore add_to_active_sema = new(1);

  /** Writer used to generate XML output for PA support. */
  local svt_xml_writer xml_writer = null;

  /** Callback that implements transaction XML generation. */
  local svt_axi_system_monitor_transaction_xml_callback system_xml_gen_cb;

  `ifdef CCI400_CHECKS_ENABLED
  // flag to avoid multiple process getting spawned to sample cci400 reset pin configuration
  local static bit cci400_cfg_updated_on_reset_done = 0;
  `endif

  // ****************************************************************************
  // OVM Field Macros
  // ****************************************************************************

  `ovm_component_utils(svt_axi_system_monitor)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new monitor instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name = "svt_axi_system_monitor", ovm_component parent = null);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
  extern virtual function void build();

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   */
  extern function void connect();

  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads that get transactions from
   * ports and monitors them. 
   */
  extern virtual task run();
  
  //----------------------------------------------------------------------------
  /** Extract Phase */
  extern function void extract();

  /**
    * Report phase
    * Reports cache vs memory consistency
    */
  extern virtual function void report();

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

/** @cond PRIVATE */
  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by master.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_master_to_ic(svt_phase phase);

  // ---------------------------------------------------------------------------
   /** 
   * Method that manages transactions initiated by master and are sampled from
   * the interconnect's scheduler port.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_master_to_ic_from_ic_scheduler(svt_phase phase);

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages transactions initiated by interconnect to slave.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_xact_from_ic_to_slave(svt_phase phase);

  // ---------------------------------------------------------------------------
  /** 
   * Method that manages snoop transactions initiated by interconnect.
   *
   * @param phase Phase reference from the phase that this method is started from
   */
  extern protected task consume_snoop_xact(svt_phase phase);

  // ---------------------------------------------------------------------------
  /** Sets up exclusive access monitors */
  extern virtual function void set_exclusive_access_monitors();

  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_xact</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_xact_cb_exec(svt_axi_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_slave_xact(svt_axi_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_slave_xact</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_slave_xact_cb_exec(svt_axi_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void pre_process_snoop_xact(svt_axi_snoop_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>pre_process_snoop_xact</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task pre_process_snoop_xact_cb_exec(svt_axi_snoop_transaction xact, ref bit drop);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_axi_system_monitor_common common);

  /** Gets the system transaction corresponding to the given transaction */
  extern task get_axi_system_transaction(svt_axi_transaction xact,
                                         bit delete_post_get,
                                         output svt_axi_system_transaction sys_xact); 

  // Checks correctness of data for transactions that access multiple cache lines
  extern task check_cross_cache_line_data_consistency(svt_axi_transaction xact,svt_axi_system_transaction sys_xact,bit[7:0] mem_data[]);


/** @endcond */
  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------
  /** 
    * Called when a new transaction initiated by a master is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_master_transaction_received(svt_axi_transaction xact);

  /** 
    * Called when a new snoop transaction initiated by an interconnect is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_snoop_transaction_received(svt_axi_snoop_transaction xact);

  /** 
    * Called to override the expected snoop addresses in system transaction.
    * @param sys_xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void snoop_transaction_user_addr(svt_axi_system_transaction sys_xact);

  /** 
    * Called when a new transaction initiated by an interconnect to a slave is observed on the port 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_slave_transaction_received(svt_axi_transaction xact);
  
  /** 
    * Called when a new transaction initiated by a master is observed on the system 
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual protected function void new_system_transaction_started(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);

  /** 
    * Called whenever system monitor tries to associate a master and slave transaction.
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association Indicates whether the xact should participate in transaction association or not.
    */
  extern virtual protected function void pre_master_slave_association(svt_axi_transaction slave_xact, output bit drop_association );
  
  /** 
    * Called before system monitor prints all system transactions,
    * using this callback user can remove the unmatched slave transactions present in
    * the sys_xact_assoc_queue.
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact Indicates whether sys_xact can be printed are not.
    */
  extern virtual protected function void pre_unmapped_xact_summary_report(svt_axi_system_transaction sys_xact,output bit print_xact);

  /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void pre_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual function void get_dynamic_coherent_to_snoop_xact_type_match(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts  A queue of all associated snoop transactions
    */
  extern virtual protected function void post_coherent_and_snoop_transaction_association(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
  extern virtual protected function void post_system_xact_association_with_snoop(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
   extern virtual protected function void override_slave_routing_info(svt_axi_system_transaction sys_xact);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_check_execute(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual protected function void pre_system_check_execute(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);

   /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual protected function void interconnect_generated_dirty_data_write_detected(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual protected function void master_xact_fully_associated_to_slave_xacts(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * In some cases the attributes of master transaction are required to calculate the slave address. 
   * So this callback can be used to assign this xact to xact present in the system configuaration. <br>
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations(svt_axi_transaction xact);

  /** @cond PRIVATE */
  /**
    * Called after a transaction initiated by a master is received by
    * the system monitor 
    * This method issues the <i>new_master_transaction_received</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_master_transaction_received_cb_exec(svt_axi_transaction xact);

  /**
    * Called after a snoop transaction initiated by an interconnect is received by
    * the system monitor 
    * This method issues the <i>new_snoop_transaction_received</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_snoop_transaction_received_cb_exec(svt_axi_snoop_transaction xact);


  /**
    * Called to override the expected snoop addresses in system transaction.
    * This method issues the <i>snoop_transaction_user_addr</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    * @param sys_xact A reference to the data descriptor object of interest.
    *
    */
    extern virtual task snoop_transaction_user_addr_cb_exec(svt_axi_system_transaction sys_xact);

  /**
    * Called after a transaction initiated by an interconnect to slave is received by
    * the system monitor 
    * This method issues the <i>new_slave_transaction_received</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_slave_transaction_received_cb_exec(svt_axi_transaction xact);
  
  /**
    * Called after a transaction initiated by an master is received by
    * the system monitor 
    * This method issues the <i>new_system_transaction_started</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param xact A reference to the data descriptor object of interest.
    */
  extern virtual task new_system_transaction_started_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction xact);
 
  /**
    * Called before a transaction is associated to the master transaction by the system monitor
    * This method issues the <i>pre_master_slave_association</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param slave_xact A reference to the data descriptor object of interest.
    * @param drop_association If 0, the transaction can be associated to master transaction. If 1 transaction should not participate in association.
    */  
  extern virtual task pre_master_slave_association_cb_exec(svt_axi_transaction slave_xact, output bit drop_association );
 
  /**
    * Called before method print_unmapped_xact_summary in system monitor
    * This method issues the <i>pre_unmapped_xact_summary_report</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the data descriptor object of interest.
    * @param print_xact if 1, sys_xact will be printed. If 0, sys_xact will not be printed considering that transaction is not matched
    */  
  extern virtual function void pre_unmapped_xact_summary_report_cb_exec(svt_axi_system_transaction sys_xact,output bit print_xact); 
  
 /** 
    * Called before the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>pre_coherent_and_snoop_transaction_association</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */

  extern virtual task pre_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact);

    /**
    * Called whenever system monitor needs to match the type of snoop transaction to coherent transaction. 
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    * @param snoop_xact A reference to the snoop transaction which is being evaluated to associate with coherent_xact.
    * @param is_coherent_to_snoop_type_match Indicates if the type of the snoop transaction corresponds to that of the coherent transaction. This variable has a default value based on the following:
    * If set_snoop_type_for_coherent_transaction has been called on sys_xact, then the default value is sys_xact.dynamic_snoop_type
    * If set_snoop_type_for_coherent_transaction has not been called on
    * sys_xact, then the default value is based on the static mapping provided
    * through SVT_AXI_RECOMMENDED_SNOOP_XACT (if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * set) or SVT_AXI_LEGAL_SNOOP_MAPPING(if
    * svt_axi_system_configuration::use_recommended_coherent_to_snoop_map is
    * not set)
    */
  extern virtual task get_dynamic_coherent_to_snoop_xact_type_match_cb_exec(svt_axi_transaction coherent_xact,svt_axi_system_transaction sys_xact,svt_axi_snoop_transaction snoop_xact,ref bit is_coherent_to_snoop_type_match);

 /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_coherent_and_snoop_transaction_association</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param coherent_xact A reference to the coherent data descriptor object of interest.
    * @param snoop_xacts   A queue of snoop transactions associated with this coherent xact.
    */

  extern virtual task post_coherent_and_snoop_transaction_association_cb_exec(svt_axi_transaction coherent_xact,svt_axi_snoop_transaction snoop_xacts[$]);

  /** 
    * Called after the system monitor associates snoop transactions to
    * a coherent transaction 
    * This method issues the <i>post_system_xact_association_with_snoop</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */

  extern virtual task post_system_xact_association_with_snoop_cb_exec(svt_axi_system_transaction sys_xact);

  /** 
    * Called to override the value of is_register_addr_space in system transaction before it is being used in
    * system monitor 
    * This method issues the <i>override_slave_routing_info</i> callback using the
    * `ovm_do_callbacks macro. Overriding implementations in extended classes must
    * ensure that the callbacks get executed correctly.
    *
    * @param sys_xact A reference to the system transaction descriptor object of interest.
    */
    extern virtual function void override_slave_routing_info_cb_exec(svt_axi_system_transaction sys_xact);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * This method issues the <i>pre_check_execute</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_check_execute_cb_exec(svt_err_check_stats check,svt_axi_transaction xact,ref bit execute_check);

 /** 
   * Called before a check is executed by the system monitor.
   * Currently supported only for data_integrity_check
   * 
   * This method issues the <i>pre_system_check_execute</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param check A reference to the check that will be executed
   *
   * @param sys_xact A reference to the system transaction object of interest.
   * 
   * @param slave_xact A reference to the slave transaction object of interest, if applicable
   *
   * @param execute_check A bit that indicates if the check must be performed.
   */
  extern virtual task pre_system_check_execute_cb_exec(svt_err_check_stats check,svt_axi_system_transaction sys_xact,svt_axi_transaction slave_xact,ref bit execute_check);

  /**
   * Called after the system monitor detects that a write transaction
   * initiated by the interconnect corresponds to a write of dirty data returned
   * by a snoop transaction
   * This method issues the
   * <i>interconnect_generated_dirty_data_write_detected</i> callback using the
   * `ovm_do_callbacks macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param sys_xact A reference to the system transaction descriptor object of interest.
   * @param slave_xact A reference to the slave transaction descriptor object which was detected as a dirty data write.
   */
  extern virtual task interconnect_generated_dirty_data_write_detected_cb_exec(svt_axi_system_transaction sys_xact, svt_axi_transaction slave_xact);

 /**
   * Called after the system monitor correlates all the bytes of a master
   * transaction to corresponding slave transactions
   * This method issues the <i>master_xact_fully_associated_to_slave_xacts</i>
   * callback using the `ovm_do_callbacks macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param sys_xact A reference to the system transaction descriptor object of intereset
   */
  extern virtual task master_xact_fully_associated_to_slave_xacts_cb_exec(svt_axi_system_transaction sys_xact);

 /**
   * Called before the system monitor calculates the slave address using svt_axi_system_configuration::get_dest_global_addr_from_master_addr()
   * and svt_axi_system_configuration::get_dest_slave_addr_from_global_addr() methods of system configuration class where master transaction address
   * is needed. <br>
   * This method issues the <i>pre_routing_calculations</i>
   * callback using the `ovm_do_callbacks macro
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   * @param xact A reference to the axi transaction descriptor object of intereset.
   */
  extern virtual function void pre_routing_calculations_cb_exec(svt_axi_transaction xact);

 /**
   * Called before the system monitor adds a transaction to the queue.  The
   * user has the option to indicate that the original transaction must be
   * dropped and split into multiple transactions by setting
   * split_original_xact. Transactions are split at the boundary specified in
   * svt_axi_port_configuration::byte_boundary_for_master_xact_split
   * @param xact A reference to the axi transaction descriptor object of intereset.
   * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
   */
  extern virtual function void pre_add_to_input_xact_queue_cb_exec(svt_axi_transaction xact, ref bit split_original_xact);

  /**
    * Called after the system monitor splits a master transaction. The transaction
    * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
    * Once split, the user can modify the split transactions through this callback
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_xacts Queue of split transactions 
    */
  extern virtual function void post_xact_split_cb_exec(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
    * Called after the system monitor splits a master transaction. The transaction
    * is split based on the input received through pre_add_to_input_xact_queue_cb_exec callback. 
    * Once split, the user can modify the split transactions through this callback
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_xacts Queue of split transactions 
    */
  extern virtual function void post_xact_split(svt_axi_transaction xact, svt_axi_transaction split_xacts[$]);

  /**
    * Called before the system monitor adds a transaction to the queue.  The
    * user has the option to indicate that the original transaction must be
    * dropped and split into multiple transactions by setting
    * split_original_xact. Transactions are split at the boundary specified in
    * svt_axi_port_configuration::byte_boundary_for_master_xact_split
    * @param xact A reference to the axi transaction descriptor object of intereset.
    * @param split_original_xact Indicates if the original transaction must be split into multiple transactions before adding to queue
    */
  extern virtual function void pre_add_to_input_xact_queue(svt_axi_transaction xact, ref bit split_original_xact);

  /**
   * Returns the contents of the L3 cache line at the given address.
   * If there is no entry corresponding to this address
   * returns 0, else it returns 1.
   *
   * @param addr The address associated with the cache line that needs
   * needs to be read. Please note that if the address specified is unaligned to
   * cache line size, an aligned address is computed internally, before doing
   * the operation.
   *
   * @param index Assigned with the index of the cache line associated
   * with the given address.
   *
   * @param data Assigned with the data stored in the cache line associated
   * with the given address.
   * 
   * @param is_unique Returns 1 if the cache line for given address is
   * not shared with any other cache, else returns 0.
   *
   * @param is_clean Returns 1 if the cache line for the given address is
   * updated relative to main memory, else returns 0.
   *
   * @param age Assigned with the age of the cache line associated with
   * the given address 
   *
   * @return If the read is successful, that is, if the given address 
   * has an associated entry in the cache 1 is returned, else returns 0. 
   */
  extern virtual function bit  l3_read(input  bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                       output int index,
                                       output bit [7:0] data[],
                                       output bit is_unique,
                                       output bit is_clean,
                                       output longint age
                                      );

  /**
   * This function writes into the L3 cache via backdoor. Backdoor accesses are
   * direct accesses to the L3 cache in the VIP by the user in the testbench.
   * 
   * If the index is a positive value, the addr, data, status and age information is written in
   * the particular index. Any existing information will be overwritten. If the
   * value of index is passed as -1, the data will be written into any available
   * index based on the cache structure. If there is no available index, data is
   * not written and a failed status (0) is returned.
   *
   * @param addr The main memory address to which the cache line is to be
   * associated. Please note that if the address specified is unaligned to cache
   * line size, an aligned address is computed internally, before doing the
   * operation. 
   * 
   * @param data The data to be written into this cache line. 
   *
   * @param byteen (Optional) The byte-enables to be applied to this write. A 1 in a
   * given bit position enables the byte in the data corresponding to that bit
   * position.
   * 
   * @param is_unique (Optional) The shared status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @param is_clean (Optional) The clean status to be stored in the cache line. If
   * not passed, the status of the line is not changed/updated.
   *
   * @return 1 if the backdoor write was successful, or 0 if it was not successful.
   */
  extern virtual function bit  l3_allocate(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr,
                                  bit [7:0] data[],
                                  bit byteen[],
                                  int is_unique,
                                  int is_clean
                                 );

  /**
    * Invalidates the L3 cache line entry for a given addr. This method removes the
    * cache line from the L3 cache for the given address.
    *
    * @param addr The address that needs to be invalidated.
    *
    * @return Returns 1 if the operation is successful, that is, if
    * there is a corresponding entry. Else, returns 0.
    */
  extern virtual function bit  l3_deallocate(bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);

  /** Clears the contents of the L3 cache.  */
  extern virtual function void l3_flush();

  /** Invalidates snoop filter for specified address 
    * @param flush_all Flushes all entries in snoop filter
    * @param addr Address which needs to be invalidated 
    * @param snoop_type of the transaction used to invalidate snoop filter entry
    */
  extern virtual task invalidate_snoop_filter(bit flush_all, bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr=0, svt_axi_snoop_transaction::snoop_xact_type_enum snoop_type=svt_axi_snoop_transaction::CLEANINVALID);

  /** @endcond */


endclass

`protected
_N3M+-;aH=fBR\PV(H0&_eB?RKP^RW<D\TE)_?OFJ@_2N4:=:c0\4)X:Xb9AAc5Z
/>9F,6;,b^1.ac(^@N0?a_aOT)g<bGT&2aG7OD;[U8Y&.O0;5\CT9TAAg6e)T5ab
/7\9XOH^GEV/_g9c.SAJS=:V]?]/Bf[T;N[&d(YQRF6_^\7,-SBL&\+<aO10aLGR
Z]F@gD0Mf&OKb8aRCK&\ACI\E0aFG]X<=1W>&,)[K-K=#Ub4Xd<8M2HY4DH)a&,I
;FP-+:COS?5B@MEQ.D@-3+]BE_A-)S0>@2@Kc9-JeLW-aI?&586=a1(I;@a]3EG,
[;2gZ\,aKC:?USW=[,[7E,\:/)&SQ1NU8BY9CE224.,2g27/=aU#D0:SM_(a5QH]
D<34gV/Y9TLRUO.=3G/1X\dJ9]]83Ke3>&JBJPP4E^WQ5MIOL9/B&CUKKP1L855c
Y8/#aTgK+FB5KW8VMUI2L16UIC0B=IIN,WbN54S;+]<<[FbIS86>_O+9AN>a;_ST
LbL)@9H\X_ZHfAKSGMO=@?[)AXdAJOd.aD\7WE[7@64,1IGQ7V;E^M@bM)c.^3?X
6/L,]8L(Z:+_F7X,C34[J8=6=5SHJ2AH4@R2=_/ZPbQ5BP[bM4,&GG5V=Kd=FZaP
\(g^45N)C+]<dRaFbgPG.H&U;f<_DcGC,1.RE[U6)L(d^c(O+0+9Q]XMbVRA:=OB
3CYcP6BRF??XRI9R_FY[,D./b+@?#T7EM,5U)1&^.^G>eXBNbg+f,A6f(f7WCE#I
7)+N3@SNPW&f[N>QW>;g2A@[/6O/ZV.[])R9.//ca==_M.P^.RJ88(A:R?<N_B=M
QPgP#\OMWCM-=WX.BJ,(]g1=JOQ=eGgJ-e?#6_\0adZ_E$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
LKD1AG7L@=H33NIY1,a;3.a046R-Y__\21X-JHS9K:WV/S<UXfAJ,(81G>:&/P?b
A^SBfSGg?c4ZI<e6X;dZVb:bc0[;ICIIL0COMP_.5U>d^^SWW6C4+733BKY^ITg8
XGY;._<IH-L[60JcQR7BUFZKBfdZUW@/IV9f;YTYA8,WW#/WU2S.YSIbX^N&0#gB
Q2CK&E=K^2;YGW[E?a#OfMIY#LY^H-b8DKVc=X:<,HDDVLeW<UPbJ_c_]D2UdM57
f;]+LaD(cX^E(;/SXI5;06MQBMD2QTJ._9Ue>>V6JSUB)Kd8-_#KNL(O_N8=?[))
M6U7X8YPO-Rf.]_L9=\d^Je6;YVV6H/VCCPEZT.9>>;R7SLJZ5Y<F<-9Pg3\eWR3
6?LD#RW)BgTgg9A?/+)B,fD6\.ec+&2E/SMT0ICF?K.YPdTR=I3c;>UVd+-(1Z/4
V;PPbT@HaGDdUW00F<36B,bdR/G9Ra^W,=.8X9A1&NYdK\B@ML8FWTL9[6T=Z?Gc
\TYcd[FAJ2-(HWI7fM-R5:5Cf;]/aH=Z.WY?ddY6e_J[<dKH70[T:A)(4?fVY?#+
8HQJ(B1Q#eWBTFfK9HNJMOI_Z]XL?_6YQZXKW?_7]QX:YcP9ZR5<F1f\SYLZG6XA
e3QMC0fDSQBY6TYQS:89\?c1deWA9EMS5g#Kd+H99EWQ3^>-d0bM7_G&A^F7ATEX
95DeQ:8V/+Y=][EDC+5:<XE5NPeOVJ0<;DFF6#^#bdG6(;C&I.L/M\IDMAZ0#1?b
:_0RPQX,f7@f<d:3H^KD#7Ua^)Q1WEC5U.W74P2Y:RH)&@BdXf;KK?STC(X1_6M-
8&bV<F3R:][BET)K8Z9Z0:?&KZ1EF_C:C^KL^><3I:f;]6GTKJ#C#(FAOIf]L0E>
0)<.d?AY?R,FHfI(V7=[D^W0I-5#T_#U?F5O##7YXM^d_J4McaaJ56M=HD2?YU<.
+KM_.,<JQG&>DW48TSTg9XF9bZg9IJbP(YgJ]SXC<R^e@LFM4,SW,&N^DF=J9/+:
(6+<]3IK7?Ya&VXfT3TG^IZZ445OIA9XJT04#Be6\<>C=/Uc-6A;PN6>#9T3)C]?
Q.D^AI.0JYGYI;&IJ]G[bXSF-<Na;QK:N6O9Y@ROWTM4D,E//c9QJGPLbKPeT,DD
:<]X+gQZMX@g2</[0=1G1&.[)MR@)-QMM=Z,J6\fdK9f9]f&/6;YTfS=9N(ACBR;
;\HeR/UQ\W:BYY4<\QVC30H<QNI2K@BGC^YeaR/^>(XSTP;;2G).U(/_77Yg0#ED
?AMU72>EEcgS_6Bad=LGbeJL_FUEB_7PaJWdC)fT>dGg4KV,Db:[PLOR.(3L^>OW
5dYRQ;#V9G.V5OM=9cA68?gI_IXbN@G6g<N[71OA^N=<_?C[MPg<?-75#W[2U,25
/ZV7bK:eTAHM.OCWXXEWJZ048GQ_bV<J>fG8(a2&C2+/Z<<35\;^;JU8/388F_eV
;HH^UIU&EBNG\@C3Cca2CAMPUVD4VV?0B^9;A]_FV>UC1<JNQY=BOBI>:W5_/_7b
RSQ94U#\VK0=WbVXOUe7QN03=@9M<52TKGW42C7Y;SPZ(-0_C4O+VMf+1OI=+13V
:I@34,g:666/^1)HRefd4-b@4NLLJV2(6D_Y?5V@Y^.4(cd(a2B8H)Rd1)\^ccNS
Qg>Q2Y3=WU4E-UGPI;#7#3fB.8./cSQAUW+T?ZVLFUg,>:X^)\:<U;SSeG24c3/?
/RAg99gO,g2YG;c^IDAK<e71.(F](H7[@eDM]:&#,+3LA4F[HX9NFf?WeU(9.PY;
4BN6/:IU9d?S0cLP&cZ..g437g^)45CGD-9TB+;25RQ-ME+<7N]9(C<-_KdKN,K0
X(K;BRd/ITH2^@cd016+D#6?GK>d6b-VO0)SE@T.NY\YaVG?b:FZe;cg;\7N_10R
WO;JO]=aZfSA5^7C<LVW=5a5BZ#JH:7L>5QUac-UUK4-+7K1ZI[fcICY:/;2ZTKE
?5&6E:UDLM]0[>E;-?;Sg>C.=D/3V;?.Qa6B_MGJ2JY8-X:DUf<Rf_2FCSB7aZRg
-ILJ5Xg]JG_.0<c[JfT0YSLXWJQX,c+cZaP8d2(F5]9UeYIY)KS=FQYM,Q7K=Pca
;K?\a+]^:436VVgQd0BVB\Q.8\@7B9_C^Z+<UE\@Se+I>4\&38(2J5Q5.fbUY?a)
@DU[V\CX6A43SP@a@VSOX6If@gWG3I\JUR<eT.^/T^6]Ff65CW.7BLRTJG[TWFd2
b(?[[Q9MRHM@I(VVVHI6U>5.6Y)T7f5;28e<X85DAeNP=KE&6Ib(+,:0;G?\(&X9
e=1]?I(AO[F-3,YL;PO28f]Ia?W6)-6aGcK2>/U1M&N5a95)1(J=DEO\QR+1M9\Q
CFdU>2W;]f2@;XSbcd18MSAa<H/0^=OCP-&\.b6E0aS)@d5f1;.H<3#P4N@5Zg#U
Z7^28G:5K)#72,1]D#R2(V@fF6H/[WdVNfZF@5S8;VB>S>L]^##E=;<]B7VU_6^<
W^)SEcF[<Z:WMK4GTWIPMD.FS(<AM+.X.e4Ac[7,VD@HF=dS;_G8f+M]0a3##/1=
WJM35bf:fQN7?9c#OFZQCa-9:^-O-3<eZKbQZQEBQ[]+F9/c5A+[e7-)4P(eEECN
]HP?L@M+AfM[6/,3>/:>TVd]P]@40eJG:LRJ#-[ZA\G4&ee_CA),9<egC3bK.BXL
5=^QZ6=8K&YaRAbN4bKY]5A\Ugc?J?[AHA^0Pb6UQCPG7RM;\_g/-3_9ME+;L=QR
OT,A6H9D;L=XX;6?)NFaV?6.:X?SfMW)\9<TBb\gQZSa4Z0-[b[POZI<6;622?bE
<19fVG#c)Oa6(V#&?[Z@Xe?3e:,S8HeX<)/W^;848S5TH8D<[)69S#UF>KEef<5Z
L=AZ+#<_d1BeGJ78R_2bGQ7TN3R]1a@^.ONd=IZcL-(X\L.]7a.I\QG\S>;.YIKF
29DR3&_YdfD(\W?YM3cSM?_/1SH\,bQ;R#5P<4QL?T^:X^&F3dVQ8+ZM)0\5:-ZK
1(0>T3a>SV5WX,@MIC?3=)Cg0g/[26?.5,d\-R6Mb)ZJLWUHE)C(B>A.MfdcLADX
O12Mb@CG,\/27@,RKBBV#E;)Bd]G8,-:81bZ>@(>O2#(g5M__ZXP?bbU#APC?1eY
&5>PFH@<(gONJ/eX#2Lf5Ggg]R<fY9YL<[^7-R/K6\-96,W_9AaP3]:T+-^<cBZc
AJg_PMG+?@f>5056VHF)7NO7/NJS^JH^Y)U<N)><aDH<K_(WZAC0PQJ]K11gH2d9
\?fR67@Ea0P:DHZ8^B#3:Y2C1ef<@WLD1(0NZM0[g\WYG_1Te98e[E>DH0feG)L>
5JBCRSb0:9eQcN/ZHe-4W/?R?O,>WQ@UY/?IRb4ZT[U(F(+RGGXQN7,[2&&YSE06
8W@dcfV64(>4\L41NGIK98Qe,FSL[aRUf0Xc3U/H.0MYBLHQ=0CJ^:1H5b[NRX,=
@2^N3JE&EYQfLCf.(JT9;F<M-4PC3BA@B>>2,3A]0VCbF-K1[>4V^T<2J([bR#N5
Y#f4@9=(YLdG)4KCX]NP8I1bDTgE9N&EP=^T[cRfJ^5-O2RHUf_c5J^RESS@?#^L
+LUA3[-D7Ic#3::)&)La0R8[4[;_gPN<\a_PV.0K^:S-2^ZD^YVaKfVC.fL0Q-)e
aPS0DdPS-7BB&fSCB]9&[@>BE(A+7c0agW>PT(<Xee+L1_cgX9+;Of-9f\_M(#UL
(X+)@+\,gG.WN&<;=N).gc-,?68V:YN/QFKD;geg38S>/3bXR.CE056MY):ILU@(
\+YN?B:)<daK<]NPZS\5W+IR@MSQPKPCZQF3aCI=/-69Y),PDYY^dQ];?:WBVYP)
;R#9YE2e5FE\<HAHLS7<(LFS8.Jcf@3SZ,2LA=6Q&9XVUf4LdU/.Q9K.^gN+^/b3
E-;7#@,WDcg>,7WVg18J[Oc^8<d=HHY.HPE;;1P6V@,3G<,FS9MN30<X;,_@ZAFF
1dQ-O]?8>V6_A\P;C8V]TH>:Y7,LF9bcJ0;)0IZW<R6f9g3J-,@2<:/KKA7:1=.2
)S4+c1KC?P/W_,X3#1ULX^1=H9RRZ;MBReKgUJRNSb4/J--M9I@\KY)>YH)<R;Z:
IDYPe+TDKO,/BO?-;MdRLO5&M+V<,Vb;1&ZJKd&W=>EQ/:1_2\[+SXL83I.RQ1\:
65:H1.;4C#BTQY]RfKR?e+>UJ/D>4845NL_1LM2Y]6L))IMKd:3cT:I#732Z=La:
XB0Z8T-0SO)OJS5DSB.L\JMX.WEeAcB^:N@Y5;FIG998.8G67=6R:,:;9MXOG)Sd
&4P3R1,[e;E3F;\+/W4\G&c3O\Z235NSCYQ^g&=8a8=/-0ZOGD:^]97J_W2?>NVJ
)H,L2^)I&)Y@afOb++.GFI9(Ic]CE=8NIE##9QX33dK/7b92#MA78L;QNX_A-CE0
MLH90YT5<#S^4T&Z9K?6=C5P-0Q3<O7bP?=4S]0NA0L#&7X8G98XQ;QQcIPRKRPP
1_H+d)Nb[RNQFC_&[?+,HYB>^90g3#K:Y-B/,K(Rg(FL_UNc&_<#US?^a/_X^#M0
(8bdF[g)H23&X]&W^IO8E>8&;1#T?A,]SN]UVT8CES1NeeQ<?03cgUJQ=3IT]Le+
57Vadc,d.JS85]K/Lc.7.2+J685>BYI<T2fSg@N3<N=>Db_]&;KQ[OY.1Qc+\75A
-X#04a-X5eV_00CEMC2;=4?,?1LAEH>4c>/8f1G)OR+9^.3F_:2#IRY\QgR;IS3.
64UDeLZ<DEV:),aN=.E+=Q^b(^aU?MFB2[6.B49IN&Y^ISB\H)OHE;/,T7geWLJ\
><D=Kc)d-ZQ,[F7Ub:,2=I[Oe/UAQYe81\O=9ZCO#>:TGG:<;=#6,aM>.e6.<Y^e
eV+?KdLDG?W]aP3b8f3N>]a_T/+DB-IGDQ49&K(4\W\SV8Y?9KLC;\)<;cJ&83gH
S2_.3W8NS+FE].05.5A\G#8a@[=DVa+<ZU.E1?#Q^HAb7E29_SaEXeU(9OZ6KWd3
2=CeHMC?M_9UP3f80JV;?;0H28S,_UV6RTa0d<OG7M;-B(85W]D\=L@R7VJN7_1]
EgIe@:U1O0UbQCMPfSVWgKWO?WB^[L?OaNaH1?1]-Re,XZX]C9FQBK/]/;gHIMf/
SC?LZ66+HR+X<Sb?-5HNK0fQ@R4a1@/7NQF#4f](]KV_P#d7VMeIL:a7-OI#-Yg=
OJcL4R+97P7L7I,eJ(FATMOF9<SO?H7JL16)5f?O,UNbE&g66P4RJN]QXI>)&f2;
L0@2Q,@J>.H.VT@UUT9G@.cZ3#7XA9^,ZbTV[H=\0Y5/\PdP&;)K+DeVS<:=1A16
&8gc@R@VVT=Vb#NEQP;.CBIRGGYFV[7VBFUL@d#]SIb^U)<dFbFN-20V920#.b/J
]0M#)eV9(Y+/P\YaFHHJ(>.;/_SQS;C<-H/3<AYR346a<+gKGCWAEaHc:cdJH1_9
YYZQ3O:eSg(7(:9a^aW]+<D00,<YKaU7C9B(B<NLM62dF9OHQ+Bg06TeO]UH6K2)
:ISCSLQ\(f:a[>S:_)F[D27IDa[DL=LBJV-O;+MIOAeCfCc(0:LE2F4:IBYO6ZTX
]1ZC0f/4C@90c1A[F25JXJKWN_U)gbW1GR:XAW/Wc(+,e(Kf<ECXBagBA4T8+9\>
cg&f861([^HIBU^WX++\3/7,8PV1J,/<8#?>R5C_)3RH?+^S+89V]\JX5(I<,<IB
6f:O94]Aa9dbW/89/#g6dXP22?586fU8PKF^3SU9e2A_.N8LO1ZB0(,=YK0VZ+2#
,P1;Z+A^H@VCeI+_?B#Rbc746BFcGH.33g+S00QHfdaT1V::aXACKUU)1/IOGES:
-&O@J#F8IO0T96651]/3,(_?FQNSF362LPHTE_adfg1\Re+R1)>[5TH^P,PH/W\Y
M5JJ\?,\>78#U28<^3Y]?bB+1?C)KH718+@UQ#HW1ePQOb]Q6I]7K?OB)4-Z/,63
GT(ZT.e_SM)dD-9@+9))(T:f:A)S/2?44[gILC\N]VWaLcBFU?6WH]M7<V1WGYE6
@:UOKeYT_Fed^/2U#@>dDU#U>0cWF:_,\/8fd]FS,:L1b;.c;aV5(b&JGW.WTYZ[
UHHFc6c/?:5F9];YbC;,E>0.#ZWa4cUGc=0/b0W^2b-4[<T]4@>d-]OaK3G;.Y2E
(.OI&M&b)S5&7REDd(8V0G;FHe16bVPSbXF/cNFO]+[SQVZbO0;99SY@+E#95eMJ
X+b<B+cg-AX07E?0.G6462WX/269HU>VZ,#P,800@0\DM/V.F8d+EO+=0c4^gF1J
P71d\E1S0S.NQW6R(#g1]^I><?^)T.ZSZ5dV2>Y=R+bIFW1S&QRWMBKK2GbFUL(g
I4AJ#,E#aK[T8b+?7+Rg7+#Gb2D^ef\QK4/R?Z4^6\U[C)XQ/[^RbUOc]6>D=3/_
\;7\UO1c=g<ATCc?_e_Fa?McKegXH[W=N5C_f._?f_cQ_#D;I=GST+_QS<[@F#5<
,e5b50K5:<TeIb.bF=1?ZLP:N?aI2UYJE;CfGFfbO+09#2I/]^)UfU9(2d1TL^.D
QfHAIU#SWCeUX_#NMU.>XJ?U+,5LN//A_eWOO<S@8-A8<TV6P5d-WWL;0\6://,+
a(^@Q(C/^3F<;H?cSg]RK+34b+@6C<ZG95HY(]O>+F_EMEFWGcI2<,9SG.>J3Cgd
+=590BB<CPTJ1#\0W6e#&PG42d90@,AJ^&(1#)#CW0Nb0-c?Yc@:\&6,0;5V5I15
Ig-;f]Q.D5].g:?-ZD,OC=T<:7/52f(SbP\L-6R.bKb(bBJMZ:(MfLY,S.I/9b^&
dQ1.T0YB/JO:57B)9:<X7gC9=@N#NQ#][Ge)DCe27]-#\6GLEUGAFV]@]GM]A)Wb
Me7QWVBTCELHX^^J#A@Qa(&[aH@>=ZQ;Q2V(V(6<3W8CBI=aA/E2dbT;-RN(bL]H
>da<<Q>1S9b0RQBNIFKF=AU_\D,4NEAC>gfe1AYV[A8:O62MgeAW/Y(OBJ06.6cV
9+B.//[34,<c>08_OC65.O9.acgJFF9]\EaQf]XeeAJ9<M(CJEF[5fb2FS1.U@(.
GU45dLV(&UJ2dSRA9B]L@OXBBIMbIb]-Z0DMB?_e8VP?AKGgXNI8Le&DaDU3YB/E
6QU+9JS\&A5EFZ6]_OSLSe2QSK57.UT+/T\F:cgS:Qg2IC&@\V=YK@]eSL9-^U=W
9K:[F.LF,Oad[)1/67cIIIBd2&>@[QMUQ[bSFS,:^;V(1/b)P5cWM?IdW[?cY1a2
ZQ[#QNY&bS[Z\3+&^^_/@[EYREVI2RG6@VbVE_U7C?g83ZN5.IH[Zd]?NV,-RAH0
J6U6R&-WUANX3=NV3fJ3g;[=7\Ucc7SEKfB;eXG7](2fCNcR_:L8FEJ:<-5dO-1K
a?<H0b<Xe4,L-ca1U+_FOW.F9;cJ-,BCJAe=+g3B1=<X63dfIbK]J.DB8MOVB]NZ
V9\AI52]KA3GIT&J99LL?Yg,\)6-+g1McVD:SA=<5X7&_^+H+C&A0HM,Y^Ec:8A^
MUNS;\;MffS9P0@XcMMKeG9#H;.S4I_ScOISC,68Pb7NJeJCJJ>B7Uc95UWC-?2)
VU6Z;J/aX@IYIJg:4IRGT4?O]OD5CHS[H.J#C?2)I#5AKMOUX\c,S4<T2CF]@cX7
d9=FY=gGAY+[M=c:SDY^E5_2e9(DNEAD9dWXXW<^ad]^?5B:UVSZ\Ke0?/+-S-eC
fE88IC+1=Z@P1:XRgfWbG]^dd?eabY[V<;)S-G@,2b,U),+?1W1@OIOMDQ5BG:Q;
SM[P^FdFb2MI1eg78^M+R6<d_/[B8d]>4c;D.O8cgS7M>_\Nb7OLRA.gU.0YFM^#
=W/,^GA_W8)cM0ab=.HO(>dK.c-4CA>8gAVE51cK[7K&8Y_BH:>5R<C&CM-N=W8M
OSOHa:K<2N4=)Q-#RY.0<84H7S7_=P,Z]L3J17)I?QVMG-6A;,N#?_D-V3g@ZQRN
&0SE(1GS#I^c=Pd.Y:eI#9IC;IR>E7b3ag\E6P1&GKLg@VD8LJR8?_ZDFHAK2_2P
07Z],daVO_M5Xg:aT6CZ[_d2J^UV25&?0[DA]/JW+Hb3LA-=GMH9^PG/[R-b<&\g
aeKcZbJBD/3K66O)0,X92;cW\)0cV_g4#8SI&.2_POXQ1Q>+8J_[QT=H6f+eIG4d
J&S#Z?I&D]?e]^F+P=RB?U<;c<4f(\X4TGD:g_9TQ@QBU@Na>YKKdX:\&?9I>RPc
+@ZJH9U/41A,g#=?V[@OAc1cJ6&EIL@LFQQ+^S5P^&Q=FOST#,:gc(5gY7(XaKDX
M8[A=+&LMcL^\EH=F?CYV@BL:EK4X,VECRA1E[L]&_A1P.Dedb2MI/eF,a[+b:#-
1TDSZ68(\5(<&7=Z^QUUV1:Z)F2I:gXW:J4L73[_H9afFK;]b8SR.CM(I)f4@74W
CWY:DQS/\#5B9=]8MRM2:I9E-Z4K0:LK1CFPW@#9JOXW7P(fP2WaHU=Z[UXJe27b
\[XM2K.EgC?:(5KMX,L\;=3QQ^dbQQ<.1O:=8)-9H&Xa=ES]R3f_XE>2d.[#JE+K
TM)W(R_f88:+-<D_G@=2Je2Z=?Y_bcBdLI2226(Y2K^I]d7cTQPD8(OUYTC#5&9C
dBC)J<NFC-.bSR/ZJVZ3aNU8[=9)\=f0).-\ILULPS3\U]aLTA8IXBI?\__83@+6
V?D9R=31aAbQZ0-4I9<(/b\^A/AG/T;:fMBG_d?53K0C[N\4I:STcOQQ6J1:>;JG
X^FeZQ@0-UcNK=/H:28\X:<7O(.F3=/e^#&P7gE3)((VGT85NGa^,KS9:=T;6SD.
<3#MP_ZAc<eAL=f:QPK-Z\)e&bUALO20S,HO3c-8?SX\LEe6eX[N/c#a7RdIV_aX
R8?)A(\-g6_;RKHgY1\(cC)+Zac\&N4RBBQ>3T(S4b(@.&\LWU3(J?/,[,D5HK:#
aD^C4/L8]g\K->>2-K2K3b@SC2:>VT?SOWDNf1/dY7<RL49-g\;g]Mc,M&FD6KAO
6>7-^TI6g/g(HGS(]NGGFU+QC(b5BOJb#JB4;A:g4B3K&7;e.6ca5/,cQgQ6QX.)
+MLZ)1YPFQVL\&_0,3bCNbF-68C3;4FE\4cS3T69>JE-WGBT.^W.=42UUQ>2N/HP
\QY6bXLKA<C;39H\J,+\84[Q6OMA3?BQ)U@:4GbP<5;-eU9X;CVg<0[ETe]R-gF>
[cLaAP?:C]WM1A=^RgP41S^R5KV6CECeZL_?A)I)GZd,:AbNcR/59J0^Xg+a]>D1
<CWd16_1;GW</OK8I=SR4+RZ42YeI-^59JY4FH_1;L))-?4Q0Kf(8bP<J^5g,N0J
SXUY(VYJW<DG_[5E+]5P;c^O7e18?a^JQ6(J1^fZZAD(fC,^V8;\bMAT]?4CaIfD
K2cegIPNIgcaBdEAG+ZJI1-VYHHSAAcdXAbbcIG1997DTD/aT5D2Md@SD-DH(e2\
0Q4Y9MN(C8e[>EB+B#/I==g]F/Ug<W4(YOIW:dg07&(-TY_bI^(X80Je78e>fg_1
<KC6_cUP#+W?2.[K>TDT@ag;@Z>75M,FZ)TLV2WfSbV=IgPMT>M0X,(gMR;..1C9
W(:C)5Y5;@7X7N-2fWB0O,.+K8d.G6O>^GWI,5\D[:)@EG[M.58/?614+[=L]Qef
=W;<K:-eKGN#QQg?S960?RJE->+&MLAD#.S65WE1?GJ[1JZEH8_.O(S0Y_b]fIG@
YV8GZNe^U\@MZ&2ORB:B3GcSBBb#>NFa_/X>4X;JIUg2fe:.Z/b9?4X10KY?YC+1
d>/aRYE:0Og4;.C?>ARHPE\07ZB_OT;fXEC2ce\b5;W@/:2ZOMC9WU3\G#aa\C+M
=KVD,P>\+b6-Q889UBcFeHFUB2.@g0&P>>:638WQU.5<7SA>9-g]g(5eH&TPHdfb
NbP19\-bb?F13S77f5KQ@35TB,#;EABIX8?7\9=<T6VU@RU.^)[d^I@e#65b)A:c
f4e2E813DY)SP,CIIK\/<^Z_M5MacT03<MC_(AQ-8/e1>7(]bC(M9;gHEV.(,0c@
9NO<Pa1.f-<Sd64M&:-0]X?aBcNKS)RaNBI3(aEHLM\Y8d^81WSB5R>KI,.YSFVS
JT0V&,]&\]EGC.(BC&J0JaaUFfL>&0S-dP@a=<a;<F]2.GGM>:]a-X??L]=UFFgT
.99e=aTd3QLK6NXEEQ3^HBQWFEOMBZ(?B1Q@KEQ=Qa,LTg50gFL0L&M2W1Q4bR[N
TaLO9UKV1Af>5=)ea3B4_534C.Z44&S]Zb)(g,[17TC/=.U-bT=@<1-2Z&7f22A9
G)&c9ZbfCU_d#5O]4a[]X]C=@R(e<;R5THfSZ0Cb/S>T.\?AKQAV[+ZZ,DT7NX2b
GcXDfY/]-YH7SJd0J4TZAWGeb82ac2O#K.88U240Z.FK^3Z^@&S[VUSV2U=N3@/W
?MP,,YYNMcM68EE1d@f]-@B./E9F]K<#61JVd9TK62SI>EFQR_D1KR:UBKf:+.bc
[D]1(;Q]@#VbUZ(/_f,g2b1S]Jd&K(C?7e\Ka:T64M8BO6Bb6+=&QgJV=I?+VY:g
Jf;P]\M,Cc<8\1e_.G4^Ca)/U,MJ@975]/),]W:N3MC4J1=c^-;]Q8J@(b022SV@
)L46Ad(eBf:01G\4)33SZJ62#PaS=f&2V?\IDQf<Q@9DR89I6(SY7aHKWfOQBgNP
3_9g58VD5NTLb>ZSLd<JB7#2;B-T10YI;:DBE04A7b;),7Jc)Y8(eRAZ;9/DEDL9
N=be_dK\(ec[@CG;D4L+Nc\P6W[-EcDeJI1F-_37DMDVSUaC1=M[]X19Zf:f]?RT
6,@25f)LRO8QZJ16bHHa1Wd_A/H(=9,e>8bH101\bcPTQgCI=Xf.7#c;SR@Z3>J^
WJ=TRDc.Z&5dXgJ3F1ZT6.^(R^->#=@R[,7K4(0(gRQ>N]7EY\C:7<TWIY[(N#R&
c.J;5-.-AJ<]VLV&,0I)W[7R+>0U)R@4-HD:KYZ]U1(T2VG6g39C5OI0X67;,1?B
4W=U+-V)dEFCG#+be]C=AC#B]CM5:-HYNd6d5BSd4OY_7#RXD4Df;VNNO.59@^L,
3M4K&4J2\6eBY/]Jb<YYYF=aJWW^5-N;S@CMZAI5g12B9c(NGggYLQ.?F,5JgKI.
G]BO56Lbbf,RY&G[K?:F]M0VY)PX4Z4WLCIEK09C55=U(+5)H03?Wb^fIDY87DQA
EW4[GG:^#dX?.WU/Of].Pc7VR+E#2Y^g6)3I0DQ8)BX4;]g2/Mce^RRC2:HOVAZ=
fG)d\-U<34/-_UMD0W^+#LRdeFH=SOTZ@U93W.]3V33?^3,G;aX2IBTX9+9+]U9D
A4<0C0.2Y3#9d40\;-<E173]B))_[TJ)#.+b.aAE9B+>28N75S@d_6AAPFd:2S#]
L2+g,#CABJaC]6Tc[QU3dM:M(UMKT6X_H]Y;Ec&E25Q>RC7R=R9?dICHeJWTf,c:
Fa<F=1W)8MLEL+X6.@e+90=FPRQ36d8L9ZE:eADc5_9MR5d-(P=b1-g6;RM9L>/9
O7CbQe9-cO;>DbNUOKRLe);fLM7G?OR3LSGRI3U9?@MK50[V+9de1M0-H@b)M[5)
SB0M4V[8L,KgHd0(9L]:@8F-XUPL#A:J^WFCJff@J#X:\C=M3#Q8X0cQ<VP3aG70
4?/-9.66&J<aM=^SaGA;O5CTf0WH9MJcc+-<)PUVOBAB?IXPKCd&[C7KA/.ML<MO
&8<9E3,c4F6]D2WJRF++Q_E54b<+6C5MGT9Z437.1/NR7dM:a>TL)UD@=+/N5HCL
WgH+G>S;S.>E4;<>8.cJ)]\DT81VJ+aRVE=Z7G^WSDcET&IY&O^^3eJdMf0)@U[9
U<BE1T+[eSW\DEUG^g)abeQ;fV2[M^TZRTIH9CI-LH0LN]@),&XD2+LH[cEX;:f)
<+L9UacfJ/FKbST4E8+QTZYXNN[>SISZ1)8dCZbAe\T7,_F]2/W>;0EXT)7(SL,#
0LT(D[eO=TDSGbU[>:\T4aGBJ\;@IPD0Rgb9?fT1V/\DUf)9L:\5^MJa:,IQ9YPP
981EE0R<?)b5TLR40VMVTY:cY\66E6,e^,BF\Y_;4ZZ&G&D:CYY[^)ZbF9WO@1\#
++):QRR8(BJfg0)I4Z&ZU9UPF]8QL-DP3X/&C1VB25cOIS+HN4H6VL#a6R&DKJD.
3_b2.[;5.C#H]>20)WCW&B+BAdQO.cF[0#S2&9]R&5=EM=CL>])3^fc#ad+1GG9Z
GT7[R5e,bNBUaT9Y_V-;H+[,aBF;]CJ;J2N8WJ,\QT:5[H=P59P?JfB:I38R108I
7E2JJce.9T4#?P1Q_\,@:b(-_D3UJ1>\PKP)7(ed2d_SY\<Mcb8F:AWZ5/3P2+U>
Be89C8V[f03&R9\-6,1<NGIJ^9T#U>\VT37bNV3eEU1Pg9<1/CdV3M.VZ9eQ=/C3
)4&dc:/<O2eHFNN.eXd1@4JcJX5Ie,BXE#.+,O(#]FL>-?1SAUA4\;@EG.MEeg9X
/a\YXV@4@J2CVQf\M)@R86K]\3aT6LG\bF7LVMCgdJJ):P<da1&9E.QA@&-]<;:K
-[e6JDKU+e47_0K3+5Wc@aa:L4+4B3ST(WLDHWeS>):P=C6R?fUZD0a1&5&1.#X[
FV3;NGLR\a8TO8+fF2&=GZ]<IcTA@BBe1R@:BZGd;[JE=Rc+KLPcUFR(]b_22BgG
?DCQWC->J)^/>_PTSSLD>Ae&_,#SYKgb-+cF=e[f2@7758S\3HBH0NH9@TBSfc\U
.H,RWHI.@MP<?#9-dRf&9]YO>g@E72F:I_(AF\Q,B9?Na;_M[U.?@NfZ:0(DR96M
X0O49OOATQE\cTXVc2?E7,<ZE\:[S,1_ZG^1:NLRR0d:DAQ0,<8-F1+F-af-(EN;
:aRbE7V(WL]LWY+7-\3:=<@-(/CALJ;f;YKGL.<S2YM-<4F@RTdY3=<C7QJ.Q[]A
(]KT73+M1aH[73<P-1?Pc1]8)#.BPP#4Y,IKCNgHO:,Ye<E/d[(9E04WdK4R[?^D
&J7_^/7_gAf>KU36M<=G4TDKMY+2c-cQ_B7JaM_&-JGQ.^5)SM9/D^2Q@D3@_R9-
#<37FN+-[\_)c6-OM3X@HRGD\a02_3D-J;cT>;:R9O)+G/GI?8R^1\CF3f]FUFT(
>G(9gL4.Wg0.:7[+;6B^fTI0Pc>S3aGOSEKMEUg+,-=\U@Rf+FI0G7Y&\P187@1)
YDRM-+e\6a9^.C7B#/V=:)H^ACeM:IDA)RIcBS#H?<:Ie5YLF,W<8\X1DQU\L&0&
,?FA&-S,#eKP5JMW12^P7Lc#)-/.:Z)fE3&:#U(c:6U=:cdMVM5EGcd?(?9C7GGU
U-JP2=F\(1F=E/EK.FKG^]_2,S&+YCU6T5ZAWaY/[[MBN/aU)RU5c20:E6FeU8UY
C+GZE[1YEOd)6dG<6F>DaPdd#/@^7KI5f^76\/QR:1CcGSVOTe5YcF@IT,^Z-4(Y
+]GY6S._S48W/aI>_Q]Dd3\CNK\\.Z@0WA3-LH\T4M30)<^#HIe1_[5;6_9N.ZF>
>1S7QWXE^gVbQE^=XD^&/3Q.:cQLLL59aRRVNX9969\H]EU?GJ\)cFb\LW#4MG\T
ag4a)AKd#PFUS-D]5ALFfg3]J4?SL.5Pe1Q19+BQ7FF.X.2bC:7D-XL?Pb>dUQ3a
3#M][9_CROK]I..8FYBD),Tf6PK=5H.O@b;QVB&QOF?ZM-V9cU-P-)0g&\&F(VP/
9@WL<JW?IV6A@Ueg3\WBJ2/3R=DdIdZ^[(PSd+c2.:AJ1U-590^:bROOSHe_;0ZI
g?O;B?BgUBT<6:fY\]E^,)dbPf+Kb\R?]_-,1U33T2VLF?K]+0>,5a:J7cP@NSNa
R>^?RS;d4HZ_J@&O]J].9>.KBgS=+&eV^=e?WNU>,T4^2fN](@[UVTIRZ7MIa=XS
-]GJ][7f:F->7=2NZH2]2\A#b2-[6>AG\.A->Jg==[C+I5VI#b&\IN&-fU<EL#Z/
OMI426?NDSTKF=UgM7a4>E7(N+IM_7?.8+HYP)):gD4;fDIO5T2H3+4\J\V^aYD4
+,6H.T3,N3P6Y,,@(EC9GYGOUZ^\5\37;ACG^4&>&UbA8QQ>)&Ie>OKT]Wc:U/Gf
R6AR8+b:,&BBHC#e/U-Zd)L2c#+(;E7^KLK@(0=D,Q7H.P^7O\VHJ(2ZLN_4\d[P
,P-ZULOQXR(/fc:^OOA+dU[T<Q6J6.?^KB?Z5U-@cYPTc2L[L8[5a+A1>P,e4V#K
2gI0B#&G?AKG&XSG,5R88;YJ88M>_Taa=9//caU^1)d@(C.ZVRXOA>1a\_Q4,)-<
(I7;<8gP-9b_=AT4F.9F]1)S7aTdIKTCMAH+_RZ/KS]0>,TW&c,8.g>55GQZdafa
VIG2QY(<_U]9YV1+4=#/@M54b0OBHc_,#?V5UFQ1-ATeHccP-T3=2\gORdM3(B6f
[0BL?XLL6aU7I@Ha&:]K+0QADH6-GW/0TcI3\P&d).,F_;6c(c#5TYR)58&B<B#Q
RRb4:]^aJ(4D/W-(#C7K4(d;1QJEOfBSa]3Hd1/4)96P_OQTZU3WVcU8OLE(0.fd
]99W-I#[8R#,NEXUMfDSOT0X_NfJ58Iaa1_@fW)5X/&73,=M<JfX[0\cYP>BP<4Z
RX?UE?b1B7Fc_c?MSU<Y/X_BXQ.+@Y(U.dfaK@/UZPX\M2RT9GD/N<\TU8QG\P5(
Od+-cJf>19L^_E+-LH6GA4.YLV>455F365^JI4?\[.DGE+H5We>UXcE#5U[U1f^>
#G3fc9I[A^1Rad&>_@3gMJTE(A7RN?OgN;<>:85G6<W0?GAe\AW9,-U:g\CU7D4a
+Z]d?-L#eg/8fS,L7DAUTR2AXefJ[KP_8PI&O]6U,EgdIbCJN>Q\G#5M=G<FMVU>
4HLAV:4:F&+9Hea@Q=S4Pg:fR-/.+FM:O_1[772XC3&ge2(HbY#\Y_]YM>M^C6,D
C@+?=.@D0>bAS1>RcUZED+b7;)9L+bD//:ZX&-+:G,5+RVA41;E5M;=]>TODO86P
ZV,Le=HgPCOSLACY53[X2CC9G6dG[7CLP1/RRK3IV@9,@46]D8ME:MPWB(,+?:+:
/\^G56GB/Uc_DXJ<O8WGY<22PAQC1Z<W2=d30VO#(cY4;9EWSeZ]:10OaDG/_->8
c@M>Q(WEeg^Db=^_S>BVJ(E8fJ810+EAQ(VB;QAODS4g;bWP+R\.D+2WfH2c:=Nd
A.P0Q>cdfP#E-.aOXRLfU\++b9;G\/agE<39:K4FG_+Z(bIC2VQEP4J6BQ-:2/>X
_dQ#FZd=9#F=>I.OOe^OK7=MM(Z=,Nd7+3&IEXN45d^FX(Z51LZfS?17W&-[@(6I
RgDFd9\BZ;[^YK)4c2H4-KP3bS05Q,L[[1b;?UUL)_I=Y5W2)>L84\b<RM-TCZ8G
OJ;U4M),:7Be[GW.LO^P#3EH8G0;FS=6gaVHFWdbT6X7J:Q0D;fSRTQ)I2b)(Q\+
3-B?MGcH.[R0S9#W?[@JZ&TRZ\0O,E^(&Z,f]Q(<4VE3&UVE:AIFJ1ca9B>CPe<U
PD^ON/DGeJZ#B/8RNY94)D[_)VO]?V@/ZDZLW&He>?6:7W5VR84B#Q\f8Z=1f\UF
\b@NH_N7BB1/I9T.BKRIQWUG([g=bVgEgSX8[/BI)ge,-E7@G._7cT_d6bg&TE9g
&_\e90KFK:T?-XZ)H(W8:I./>4W3AW67]A5)Y79SaZR/_eKMAc&SP1EP)<A7?FK.
EeOL^&fZ0]DWIS-8,C\Jb]?VdUYD&a3=;[=[2PeIR4CRM3@>3:RE\e<;86W;9<M;
_R6cUg#Z2O_VS)>S:.ga,(>e;cbaXJM]3)[I_QXg7(YH)a?d1#4fI.]J2RORY#>f
H\O4a2RSB.VZI7]U7?56W])Y.Sbc[g>++7;[Y?ZCM1b13\ZY=aG-;LCW;=(T[EI-
[?aJ+VULcT9ENMBA>BVUYb26.Md8N+#;Y;g9-L;cF#Q>aRNRNX_E96/XWM_&DE+/
D,SB+KH6J51C\7;?7;+E75\DcMK,Q&G+15ZcBFU=^;,I]bXdU<_?^.\Y423B;267
85+e=SY4(\<I?-PZ98U>@#T,.f5P_aO1gEYO<ac(JIa,DJEWSQ@Ba6A]69LW#(1#
(;CN#3ZS4APdMY<fTd@c0[;@aNaSZEG.R1IaB7UY0QBLIPNRaR)492F.JSd[Y7/=
FFN5KQ<P3&CJ><-N<5,d.gJSGX(?7OUaH6d34J;OJA_YT^HB\6#>NPI9X2&X#Xb>
=c#H_^JMDFf.L@C>W9gY#K9cGAM8DZU(Fc@G+F=SXKWbgW8\8JZT5P<89TA3H)f[
Q(?)AHge&WL7b7SD\@?A?.@=Hb<X@3TKPR_2OZ@^]D,9#Q=gR#VbV9[R<g/K=HO_
?OM&)O3WY)eB[4RF40;P[4cHK^DH+K/H7G?4L@=G2,&(&/<K6H0[AG-+M[/KLYX4
DAMd4>C^R7_a0Ae2&G?/N+;=,1W(?+GHGYNYECU^2MF0GS&HWI5eO5Y=SH6=e1>1
(/&RCWe?W6L9>^;3FcV/Y(+NIIWgcK1578<=:9KV\fW3@78X>5bP>W+<-3aR6RQ3
I9TUB,P@#EfF#gOC_,FN^(fg?/ZY=R28ZH>UK>OM)+#44J6F_Y,=J+X(XLK8\L\W
KfUJ/?VJVHb#++(7VBMAMN(;R:Z,Ub^NW-26PAbAg+M0T6BL9S&d7EQ)5N>(\e=K
M>.I,d>>-@d?@FOJETE_R0OFA7(IZ+W&f..2Kc]11ACR-/bWdL9ATXXCWFKDE4DY
=-Q<_5L#>T9F5_W:>@@1bEKC9V_]VO\=(2(DXPC)J.aU^_58Md.3d1@g]g?OJ[QM
Wd253+]g+e72)SCdZ#AeC>d,PSdZb+EC1R=KB0.eAQ1bSdHBA:6MTSLAE^X\:28O
YK[(>X\RX/2V9aCG-2QITN-5Y4MO3O7f>&-+;L5-.f@Cd7Bf9&XE]aG^3[.b2<fX
T@^V]=OXg<B]92=<]X]5VB?3dbZJQABCU.29=FPIY:A5,)=\K)@3)7c,U6>JH-7T
AVD8OI+4:PPF6J:W12&PJ_EAVPQ3UPRaML2b4_>NaeURDW@;aX?FNBNBZPeT9J4G
&?dSFD/\E(;J@/PY-PX=WgWX/O0dV+87D8f8,G[-U7;J&&_YC[c#O:WW\]W4>T\1
]EFXgE?R:P8#6Ha8&)KKAf\5g[RV?2#4;E3TX3WcgFA^1VgUK8Q_Q,Z&<:7P4O:3
-[MA?U[3SW&&R=,Ye[VRSb:@FaaTZ\5T8?KT_FKZ>QMc-4-If>&X6L@M#QcWSKVL
-=8Bc3Pd9/U2-bXU9>Z,N1QfYG7V->PLIQMM?:LSR??#=6A\@/;g-:3GP)B2Za6f
c7[S0IXNcL]+I2/DU.Y+Db_JMERXTD.LEZ?J)M>8_YJT)7HcIT4TGdDSE-ET^X2?
XD3\Z(^BAAN;:KCRg]B)M,TLHf<\C),GRVH-,d8OAYJ>KeJ#Sff2+KQT1d)YG,M,
.IacF5R7e3[Rf?90)P,4\\.N)K6K2ZZX:c+6]G;+?]4DXBDID65\Q:SKGZ(PL]Id
YfVgYeJH;K2(7P@[Ada4Da3D35]90RQe?6<a\BA5I/\R0KaAgL1TF(EW<.5g.K7O
:(a][_.TL6d153,ZSd>Zd:]-RL)4XcYEWN7]DDXPG>6-deg6Dd>D(MgGG@d0CIg=
P9_</-#_4]DXR:N;<,2C7XB_ad&C6PS5LTe69(0[UB?AX=g4-Z>-H?g,S6U8c/3\
3O<eWOE+TYWUR#GTO<EffV2II(#[_D]]^(fR#CGb=CL8CP8D[S5K8C=1=g?D0K(R
JE#7@::JBBVGPP)Aad77CQa.gNBWA5F]6RPIMCfQ+7TNS2L^Y0HfM1@>7PA<1a#0
<EM.#N3a_Q(eS3@0C)]^MRJT9JT7&HO-GPOMVEF7P7B/?BL09^<I+<S8,Je;[c(f
9T]GP^eH_,TV4F2)<Q02W3d5UJ6_^2@FdPMf>Z<63.7X)Jc,<,C>AUYJ,F,8W\)?
@DHK?7&)cU5PUQ_0HMW<MYZ6QJF^&(CJSDB-<42\dOEeb\?f@E/,AGGV+^;FV\Xf
8,L8>8(dd6SN(f)b+&F7f.7,RaY2P2N?eQ??U[T>BFZX52(.c7I<;b?9gJcHeYM8
Ua:J.B&@KQT\Ib8O,#YQ7ef.@C=7E/.5Q6FXcILaRNG(8MX&2Y,\;&=(BAW.eY4A
0F^F0B5J^?)g:J7F6]NU<=T]>W9&=^K1K\P[@<gFZ&bb#A/;KVg=g:9+CNX+Q6KI
Df190X3#+&\9L0MRIf7V,?QD5=(ZGZ^.4d-&QT>1g+cdJ_>E>99R&0)8#40,JJdb
?C;]GgdSI;V/0N6+Ia=gbO7G[:?O&5;S4;XA1(_P[^Uf+7Z52f9?6V@d>9Z+>]\1
[a-T>G529EL+<Y@F@9X0F7/GT7=D3Y3;PFI8.0YLDeU91#gb#J(H]<G+QV\d&KJ1
VaO.IF\8OPXfb5J@>>3c&RfP#N>bH@e;B@I+85OS<UXQKY54:AaAQYc82>4aQ:_E
,(Zfb>XUaK<G&/fc/N:X[?Nf..bP4L<8CE-_]#@:dcfDKZ<66L_BS;a3.--->;D@
]D\7gB/RZ=P-0:U.egDY/L&fHb)8.IHD),Ka#JG?D8Gd;=;QDPX@_DLL6M8\1_f(
ZHQ)L)#22g]SCM:Y4HLFO@R.^E7dbU3C=5+^CZF(T^VC^\VYgaf(?@SA98=\\?.7
U.Z=6;90)dY;3>Q<2BAUZ,.SfXX@O0TXV):EVd1b,:Rd+,B-R5XIacK7^e8aPEHW
aR,NI6J:W[e>^e5WCcdDXCAHa?BQK#d@H3(U/b,>V?]fR5O&4WSZ3:M.U9-<DLE5
2V]_Q)K[KTd;f@Fg^FObSJO]3\GU.e9)\^gN(/NVI0e\N>-T&+NGL3PGLY:BY6/0
+9<=T)K]cOQ1W\I-8^5U,2,G;:Jd>ZKW[>MVO,@:)(NdO<&[M#7Mg&@N.8/?&cU7
@]2/YG^J31D6fc>4_WUK6QAYMYaDdKV+1(eQTSMOZbbgE04E9aTbe9YH,KHe7ZBH
fESINF@aG80Y6H@>C.NF.MG,5&NUJcE,1ac<,,CSRR=ASFV]51;)VXKJ22TJE(P;
5GEfA0cX>a),PELE.EPMQ[BEMV8&b6W&+5,J0FdWgFJ>cA2d&E9PQ\[FbV-@&f^S
,D^^B37:2]+R>1a7GJLU@g]+X4e-TOQA5U=fP4+[55_;OfHOHHZ[8+0[M\<WL/3C
N;3E-ZHC[?0YY/-GW,1V+)f2c3S7ENB&.AA>ZF[ELW8^=0a7EEK<ALe,c.b(OS=,
O(8;?Oc-\^(;ZQ;YbC^/7D]a1J>DcbJ>CE(N[[e)c;2.B;,H1817))\cLL;0-#4F
G&bgb9B5B.b?Z928E/N2NIT(a/;)A/HaR=bY6ZMZ@;>[)bGBK(4CUF?JfcKF#GL2
8c]2@4fULCVL^4YeXQ>bc=ID6_:Z[PGE9(#3)Y[ZT?\TO5DFMI#=(<GA2>VO5_2X
XYC[6Pg:DSA.#.0,ML,bI6XDZFF</AfNJ2IG;:H0C5geUefcbM>MG5UXJG>ZIP@(
[,UA+TZ^Zc)D-8>--YF1fA&U^)STH-)ULNVPdKX:7D+O18C-1C:^\>A+gH&522=F
Ka:+IB[QY.QXTR65^?L^QS<MVF?);20P<\(<,IZB8TY=F>,-4/gc.1@TLU>bJV_<
NTT(a(-9U2?Q5(2^K0^WabEC2X9ZQP\1;^4Y](eV3cN;]C\&NQ_0?^]DB?\e^JZe
<0PR5.8^3W&f[d[MKdPLBXOU.JZ/42gIC8A;H6b2[[YGP2e#eH)AeeeF>K<e6NQ0
4\KaQ1L_IS(:[:6ITJc.8\9WGAOXF>^Q<1,O_^B:a-6&6:8VSb6?JAB];c?L\?,;
EZ+[B2EZO5OC/Y_UZ3C]4V;8@UgAFGJ)UXG.?gGX[#G#F2aR:,RKG^MQJ4#=72XR
6D8M((1[5NKI)6?_AIQJMAfLO[^0fKa(0M6Yd@WT<fCg.S;9U<611XRNN)7-3>-4
IU0Y)Z?JW2c5,UJ1;AOY^3DZ9<F]O\&,[+Q\DDU>+T\S6dFIVN)DXIFAF]A\)J@0
T40c8\2bE7ZI@VFfA+4PgP:TF9RF)3<]AW,CJC6PZ#0DCDe2XTa5[4/>.S/CJU^d
[3<2WKUe9P#;UT0&eDO3+N5e9A7\3_VRC_F2_\7b/C<e/Z,eH:@GcgAU2G[DeH#W
([;2?08\_bR5(g:CA2QJA0JJ=RHIVZ9.NO]Q^UE^C3D\2V?6J)A2YFBQ5.[^8/[C
UeZd2Q-fW?:K_VXc\,<AFdCI&1M\c[AR@(2/UFDF&eF?eaZ54T>ED)PfQTHC61+.
D0VD/Q-9=d_(AS=H0VQJKcD8P-AHC009X0_D2=Ab>U1c+&e:ed<?<GY-Y#fU=8;O
B]a9?aZ/MS/KPJGcH./cI[Z4,fQg6J(dFb7g61>=7.]JAX5K29^P^2d[U,\1+.66
7TTf9DB/<_&#833>_89/WE](=-b048O,6H8<fg601U&0M(QHdU?_I<FfdX:V9D6E
U?b__3GV0JYG5[4Y20XS.I8,\Y1#]b->>XYCV_U\\RgMc84&7,@TG9@J+X3LODTQ
DV7?E=X4S(3;<_US3&6gLZSRHg1&KffKSZ2e3F80Kd\R\GLERO(L>fF8D+H,gQ#3
=5VP3?ASXdQ89HU>gd#U05:ULL;9_dVWeXe)R3X?Z0D60c0XbEE<(0?476Q&K.Sf
<a#=._c1:C^CU&?6;M,SA563eX-(-Qf?d2[3g;V4cE0EZF>5)WAE0;8/V],I;3f7
O(RW:\Xf\^B#2)@I?P?B#YZE6^=9_BOPM=OWZD2?[A6TQV]PB49T/#A:FLQBRNYQ
J.J<Qca(^eX6#&U#V,aO+CB@23cfcg3O2]50C-=Jd,,(EG5OI0SS60MKM#Ye8NO.
9_=,<O=bd^?M98Le)be@d<HbWTFa;#@VgVZ=+SWd><N]K:NK0=H]f,W:-D-OQJ9a
\-T.e(#4T55P(?:2Q>8))CL8SgDJF8J5Z=;AI@CN)d/[_SC7ZP]/L4RGUP_9O)W_
^@=W[]eRJcPQW:,>OSDfQEY:@KSSTIC3WEZ45U:f=]?@CAGX5.?dGS;8PZY>5/gM
Qd4M):UUA.b#N,/bHeZAH0?e]>CO+;JS7N-:VF5^ZKcM7.5+RV4C656_@bQ4>)B^
/CK60?8+ab6\,2W--VOBN@fS15?[dY,EcG,V^_B-)dMFELR19bgYd)>_OWQ^#ee^
gEeC(g8=9fWaP=)_,=/SS0?;_]_5,c,-@b+AE<U2K:B@6<14ASLFg&1AW6f4Z<C]
M6CI9V51D.JJP7^(9XPDe7087b]8g>g/-dBMa.1K>_]&#d7)\XMJ-.YEQPMI5&04
>WE+af]BDbY&DOGC,\L31.FRH4aBB;O=+8&V[/Dc#b?IM7Y5OdAX),RWYbf;47Mc
,4b7&8]9@ATaY1d8gJ#5+cCT]^Y^^U=c91S[+IX=3-VJaI-,<84bC986X+O,9,ZX
Y2SLEE1XOb-5>XVQ7FM48c5=0Ga##V(]]GaMdT44LdO910Y=/13^R+f_#V:NTZA=
:J;XW^V>_ISBXc7MIB[(<K1?03;_](<c#ONWF8WV#G(0V2-&[-Y+;O_E0]M=W8@,
-Oe4+6Y.eUNF[#)[?H6<VFE-g3&3^YF?e1M5TC?9E.,M6EgBF]IR<VJ/SV5eCPPc
X/CM\3EeC&00\a:3Y#ffWN2K9e#B(HVdZ=2<OPK57+_KV^A7&Jf68dO9aCad-0ZO
X9D>=NY(0?TKX#SaO7AS=8^I&B,Z[e?HB]>[]fM7,4./A=[+BY8PQA.?_N>KdULR
W#]<cEQbD(C=c398c1aPb(JTE-:C\,D#,=KV>4AKXTc>DUJWO20TDMG17K@1cL8V
b]MH=;X<>]UCL;SC^Wd&S(6IJ13\)ZW@Z7#6fKPPG8(V.(NOcSUL&]G9=8Z=e/e)
gL\:XP4>-69fa+Qd4fT6g9T]ARD>337TYO,)+gQ>))@>\<]b4?;=\@d+A?316GDf
QVf@ENcE#SSa&eG(Z.HB\#cgbUACdZUVA\(:^CI[Ga0bF8J8<>1LO(g>LdKYcBQ+
(PZ7]GUG:P1Z6f.)1FP@^A]AgLCW]]F-KBEXT+T5,7W+e1<-\36L[U)?g_95YG1I
L28-:?6-H?)J[@cE@bR7TJbD_HOEB)Y(Z6LI4S8REPGDb4&<N7=Rb-LT14I(He15
A..18^533>G:[=D](,>))8>B?2P-?1\HHM/KQE0&F17F1:^P4)#_gZ1I:6XD<FD]
89H+:Z)@Q_?CALCVS[7DPCQ)\DH(35bfNOV8cTPE#_Ee-ag?7Z]);A3KBX2]_5f]
C0&?E,L]eFe9(GXDJZ#]&LS[=MN/eM5W/5MIfgd)IRICXQ^#6Z>=SD@LLZES)bS:
6IG?0=]C1N9B1./aeGZ5Ib3^cHe:A[e-fBQCf[D8,><;ROf<90YO8_52K=NKDO9\
T+JH4@ZU[VOPP+f++)C8H]c(04-AP9e>[4N5Z.#(0bF#\NFGH_CV=5_=1B_>[.D3
Fc;8/3cf0=#3MSGeC+/>YGUF_Wg&:-1.GM9,a?<d>OR&K<503I&F@[GWOfC9[1g,
DN^[,>0.[S&^G>=QX(W;IL(+)J0)b?Eg((_0bQJ=^/S,6AUK+/6/5]].LRT2N^^=
40\P0?VZ-UP@#RfFP#_gH)^]\PbMR0TF6T1c-g;6gf.+T\\Ia]V;L^5SB^5Y:(/,
Q_FM113V:I]+=(@W3WRe->HQ-A9+L9&ZF;J)c.ZD+Xc06F]eS>]]76LKHG0VH]fG
BA#S_#U]8FQC(H(XFWEQ+.f\#_?PZWT;(\4RCe)@>J8AEKQ<TE4==GKW92a?N/bO
He_G[TOIbP-31Bd3d-CZ-M8BH>GOZ>SdRCNGPPeS,=]M15]17\,2a/1M-0GQJgd[
E^-+4ZS8.X,Ac^QQY5WFCe1GeM8-2Ie^:dVcgSVW?U^;0P;EB,JK_K.9GgR[Jdg.
7P<W:&Hg^BWF.J7ObN)+E?,7EE(T3R\b5&W50bMDOO4T4()eD<,F4:4RPG2NMM3a
F@KV#03TM^0,dTRec+9[gWRT5^&IW?.JeG_;Z@Yf;SM</.Nd[?D,Eg,TN]-JOME.
M4^E\C5#3g0/GCO9D.#QMRIF9eT<6,Ye0USM?QV]ZWII@8O9KR64<<=HROYB7_,J
dWe_^OQK/LL3<W]gEc<]<M9)Zaa/5B(If@.^7X9(>(1VR73C?K:-@(29cL/,>FJF
c-M#;B.;_S#>]3O2L6#I>-H+]PJT)]N-d&YU->2Z..g8KP@FBe0K-K4U#5F0?6=W
<R7(Y,aQDT1DcRDFN&3d@gA@KPHNg8+M(A]YW8MYV1.eb<)O=fE3,LJ0,BVDA>SY
8?Q]fH?[1&Wd2W)9GRN?>UOHBbS^3SH:6O64X4[IEgS7;3fH>3F?/TdL=M08LV4b
C5?#.B7:Y?^DbA\Y5T+D&SY:YJN(>S/)57U.4(AK2>/<L#AGH:)=OaTPLa-V+0dE
b+GF_dHF@]0YH/=aBT>&8.BRUcF2#A=ATKbPWc3@2H--#O5Q&AaXEU/K6^S>C@25
5A@FM]Z84FYc;1O7T&?6B313R3-;fH@J]&6O&d4RW&>&E4#HC-)aNH=#)D-.EVNO
&>E704K0+GEG+=L#U6PHCT8cCZMG6@.II)@JGY[;Aa&XXB4O<4SQLM-[_3\[][=R
RH-Wb1DR@C/-g+[Z+c1M1[G8L+^@UMPCSQX-I]f;KW232-_7<C-0[<3L[YN>3@ZW
<N-.BG4GYQ3>[#E,0>J.#?3/XUZ^+E=3MH,8J?f+#ZIDY#.ZY].ac^HX+=DeQNWF
GYJ)N\=g=Cg--KCRRWe#HK^2)V8)EK?_W8=,I/^55a^BA0V>Bd)<S41<N8Y[[=M7
0/8b](S._1EZ9F-;E:;)FF=0ZKEYR-DZABQ/I_I;CL6K0Yd)AD+>^,6^c+)3&H&X
a>b]4+V(TRYg9/+\0gBT0fM90TWe[3)5fM[)WEWTW;34()F:=B<DJ/G(\cCQLZWd
?#9bd_-.N^6EL>2#]f;gTBCNN?BUV/CC\QdEb<<R->1E3OB&OdBC?888JJ[.f1/#
A?T7YJ]\6ZG4P7-B,FW/\&T-#E/YbfAD1A4CO-9OQZH(U]:6T#981gRCgTDKd6BV
[1R?2;c)NRG8LJ=MMV?c;J6/Z)#-^PMBfB#bJ9=D8,7/[PYRR61?8[-[+3Q1MP)O
XJ8#4O3<VI,(ca+[]2RZZXIb76N>O\5[Y@4:4^I6&JJ2H)ZBOBMC][LN=.-OV7]X
-@P,@V\/]I:Zf(L#g/;2HY?:_(;H@c-5GC#S.ILP.64@D>:4_<JP/R=7T?D8<^\Z
cM5f[]9K:7>9EB/[HA)K<>I9eM/DUP_,S.J1g@.R^AC)C4MCALJX5f,:@9dcPdfU
d7;QJ.QK_O>>1>MX]Q5EdF.6/Fd4BH[W\TcC^PL:d<C@0>-^USJ@=[c_U.,84G.&
V;1R9)&#]eL0)dZL@_\ZI4]M3S-3A(SIHE^HG.^G?fS)bZ37AP--NfR]U1-Q.]TE
S^9DN?/9-6.fWM.#&e=Web(&\0@f;T]UO?<J&aR;5JJ)Pe<?M?B2Y8I5#XSd8,Qb
Q.63J-Ic::C(V7U;R@MVX;+NDWKW?2a&)P809?&K3/9SBLc>=[(.aAOfgDLU?eUK
/XfJP7@0O\5V]BX;&89=&GG]adTc_:ITgF8S:F?X.P5F7&BO_];]:_)R\#MRHGVR
-D04W]N3<&H:9+_3HRDKO6+dce#c[F1X)I3.],],]<fCeK3R_[BgPGNYJ]Mb&#__
>8DH6H?_40\G3:SPd.#cJZ29Hf;6E=<WeI&,/QPg40]^7MMLY]=gVN059,EGd56<
3T-,-L2&6Na-40.NAK>Xdg0\H/&2W+590WdW5Y.Q&Z7F;_J\^OC-A#)LUdD#fEQO
J8T29=OcZc-DB93aD#@?PV_X@:TfY;H,I30+VeW]CK_c]R)YFJTGU8@5DM.JY:W\
JF77QZ2-QCDA[4C)?O):a]:S3H4a=@5Tg#1@:ZcaQ@JWO],RbLL:,TE^04SNYX=>
;Z>[1Z/J17.U_MF[7X&PIX>Q7EA;CS@B&f@51:-UH9;AV_)-(V0+,3;+[QW1?1-S
=4S[TY#D5\MVK_?aSH)B;E\.9@KUW+>)[e+D?g/.&DR+Cb:HLdbC0:STd[NS2#ea
Yb6L4Q#QgB2VF>/R)\2Y[P0AT53>F<W(0W7Z._R2dL^97;C&LY<KOaIP?]c;ZD_[
1cFW]>\MGSG.UfCb@U+FB(dMJTbVFab>C6gYZ55F#:.)d7.WbDI&Fb[C=S@)XQ2I
>I3V5CZ+-=ba<-@-?40LUOIeDPe1=6daA[0R1CaZ_Ag\P)VcY,Og.A-S?@.GZH:W
c6Ebe)><O3a;IVR?.aaWaFS]-W3.4J/\&6c]@7<27^;&A@AOJLNR^ef:,#dL;&&N
#N@YWG#981g/6J61NfQg->=?\J)a\Z720]1&1QS39]Y(1^(GRf10YT97HCBK_d^A
1@J\C_\17?5>TcSB:E3CJ4Pg,=bYX+=HN=8GTPOX+J=fNP?5dW/\(?\<GCY:,Nf@
L\<>OR4G6:S:LeF9Ea\N^Jf>Efd(&N]3aND1#MJX+:a8dF4C1/UAVf#;WJfc0@(<
4PT9DcaXYa40CSa24<94EQa,eb1Q)::RBU@ND=A4SG<dgI>-0e=XAcD-5\6gV-HO
P)54;7.3,OM+-/U)(A+TJ_\Y4dN3\6/A?.25C>E-=MP&IB)GM831bRZM?(Ag-_)<
(V&W8.1da342@aU:E2/S?^43YAK4d9=b.E,^[b<O#DR:&:YW+/57KFd>QY_-RW9O
:I3a6^WK\17<WDdM8eN6>99)?4((U6=I)(9#f;8L2FXf[#H/-6V>QTeLKZ_\2RUe
,.IHCeC23b1T._9R2(&_fJ7=Me(R^Na@\W2#G_Zc<@@&eeQg5-J1]Gb&5Q@K:7N@
;-f(RZX[9U1YC1B2gYNdWYFFA,TO)fSJKK33H_<1)c84.),^#\BYZ_+X8Q?.(79A
dLZTO_?1a2#a;e)I(A7CYA/cb?W;ODZ,<f[&1D@7;CB(2d^KLM8.7^1G;70Y&fP?
625>ObJ(=bFFF6OE38-Wg0DO\22Ne-/4DYT9&S:/-84N?2g=Z\26H-CObC5XOX(d
_UW-J_X>CCE:#5R9ADQ84,S@[f]A>\\6IFX_1])5c5H@eCM[dJP)d6?#3TO^HM<&
:H>,IQ7=<H))4d;XMXP98LVU55WE<983:J(gJ_A.fDL6:SZ^@,[3C8\/]56P]]@E
K.X-b[I?1=Y\6I^?[&PH4W\52AK=NX_LTKJBC)?S<#e/+]V+JQcWZ]Nd@NSTBXPU
.T_E3HL@0,aJS>.,PKJf_DBJEZX1\C.&ULO/85\YcC/e9WPPJV,(B\YM=8Y8Xg=<
c:)8EIQJL:1]\fT[A9WO;/]IU&Q=51C1/&C6#_\]b^#UB,K=O_Y2&D75]+AAfSAd
aA/OGVAF@eP=VDGI=S=4ZA+WS@2I/?3@&_Cc.^ZQ:0ICG-SZ[&N-A:2J3/7[2OAA
(9.UB=;H#1:f>LeHI2Q:2+JeP88#JGFKa7(5;0)Xc7N<4K\BeFI8JDBDE#Q6AdN=
S(ZDcEH<0P-V5ZC+e^?7U6YN<7e__1C3BW:eGIKVE1O?-&dZT;F9M/5_<AI8T-;.
QKe4a[DX#TWbI2b<[8,=Ja)#,_C?4ML\FEZ(6#10(7O_-gQN00(OgJD>^bCHI8JL
D+H55ZYT+(\CQDceeNa]VSQ9K(_Q5=PP-[>KTD#P4?,J2KEF9:.MOa#-eC\ATF.e
D,DKYgF@P2O-.b;(\RV(=1N+WY7OY#G/R/(3b6[GSH4>:;HJ]X(6QWQOfONWM29d
H9&^gbHRa/\RA5W-U>P3SC<VR#e\e,Ye0:9fS(UW6_/K&e&\W-1Z.Y5&=O;C94:1
X[e[<&KL)Z6[;bf.[Mg\VS#HWI3_aNW7,#=)8A\]X1TBP_KAFFKLNB_L;4^g=@2Q
^8(.?]GEQ^UeEE\=BT>X-0>[@>#d);/J+^=6/66?W&,Y@R58BO0Y@HF:.;BD,Hg+
+X?SA2gR+g49EKY(^IUI\DA&W/1IDN=Me2K.3eZOg^?]4ZSbNMX@dH-Y&3d.feF(
0NY^\(2E/,,d4dH7:(EB6#5FE#JJI.;dSZ:W);,QQCdRAR:\aY04A,)900DCEd:?
32BSOM[Z[;egV(-1M#,f_7_H2<K6>&>MC?U<aN@;d[fd1)R18NW@B/-4^eeDJFKE
Yf0,@ff),^^7RI+&f5a#1TgdSU+YX&@e8?.C(1ecD>;ET.A2&#7Ue(-?05K?f>@f
5G&-+Y#L((GQTXSXXV,CF8VBbA7J?>dAccL#Z]PE;[=7#?:+&(^I=Hg;eJF[K+cR
G+&0M,37?>/]RDPd3[-(6dXP/VA\Nc)g,J:85J]AOP=0ICaY:E^R0X02#g8&36fJ
+PG,3+M;5@55/V^?K7>BOg>[MaBBRbP6LXZ.>Gf]0;I/[C2IG95\/[6N<AEQCY&1
S;N.NNE=Q=E#;Z0cDQ9B@=R>P<SU2gE38BUCPa[B/d;AD^1S,G;,fR&6c4O2JHJO
E<b52OB\K16f=2BALJDVQQdX+e)]A=Q,<]e;;Y-&aHSLXA+=536<9F5d3>/Y]R/#
YA^c/J<ZXf?1.U15\.G/Pa<3H(/_IAZ711UN1=-f,LY+KG+0?IP+XNJ>(1Hb[:HR
;XJQ^22f@cU6_.=R2.L\-&;1M&5@ZFU(<EDJSH4NA<:D6V8LE&2_5UV_b.EIL,eW
<4XESVZRA.JMaFG6Rf@TOT2g[+3->RLdG\#U&^2:RMLEc/:AY/I7R>96OHfObRI8
Q.5aVN^&+?>;b9PM0bXfcJ+EGRE._/21P/>\(OIBYB=/bG\#S];1)Tg3T];+N&V[
G6=I(#cE#X;,c^FM//<dU,6H6>O?PP(FdIa1LQJ&Mg7dP3/HPbO>3?-,(d8NAK08
2O(bg,:KU&E-M;T:BXd:_GVGY]D^@0Bg52-/8U>^:S_VS1E#:f;X)<3dBf<9/7@^
F3;LNZQ76\X3;e[0(+)9GDX#P\X4FE\B<F/<N38(CH-^9#.P>;Y+YTL,KAS+UX:G
O(:@63g9e(1QQ8TROW>XDe2JPb3P(H(MMCFNT4ZR_aQ9?337(,;c-;7].SV#K/5g
2^c_H757QPOCgQ:.O[OSLXE)G#D,=7S0F=?J8O(@7&/BIBgM]EFO/f6e)^[eQL./
=c?bMR,9M,WW0VU27+&d@<;VEJNb=RO09E-1K)KOCR]gVI>e<9(NK1/7@@cU8HM9
(-&E[]W&SGJYc=4E<:f8QLKY=N4<X+N4aGbR\O>G2+E(19,I>N+TW:S@OJ)2S8S8
c,/.__A5J)6Z-F0I5gS#U9V+Mcg(=FUO:&)2#ec.aS>N2\/>CY[:U\K(C90G=,cB
6AR?:DM.>N>TL.ff+\Sg)c^S=I+IJTY=a.U_7B<K<Hc=W.DK##^/^I>d7JfaD#]\
_\_#[Y^BE][#[Td;U.A:A..@72HNQQ0TW4B?448XeXdZT=UFS,&O6QYMeMM16L;K
H3KOY/L4JF)UTAM]^Y8>C?aWc,B+&\\\UKW-HVBP7/LXdW#(4^:Y(V+G_]Y(CX&d
#MX.8f&.6HE:L1BbT6H^MWLX8O++Sg(@#L?(dSO+/A);7X=JP0.\-=D(RBEFDN;8
[S7,3AV[DWV2EKaJeVBJKH6W7,dUbL.Y6E8a\d/cJ#<>H^dcO:2N.B@K?g#F=?N,
JE<Q,HcB69)Z/6-JXWLFF(1PM7Sa.[..L:7PH@P=VD.F\WAQ+]<D-W6[_AHD?815
?HX^XOA&/;6M&M0.5E<&+@^?L30bc@3#]WM:N?)2,E@.4&WVB_[0R6)OC<3]#-S1
Y4b]G__FP-XLgD3A&^EPL-f@CK/<Hc[bPT/,IfY^I:#3H?/[Z=D6#O;X61d,=\AY
29NQG4.Y9N\.FW_7bAbBENd3X,5f\4Yeb+J7a/<CB^B;aHZI0]FN-\cQ_K]g@\0@
J=P+WK4;&Dd(-=T\b#8>:86P;-FgA98@U?4RI1fN9>7YM<(=;5bbd\g-,Y;B:TY=
#<aZ.eJX;7N073d?-5J]OF:I8YF9>J?.a-7935N4gfHQAd6:J?bgU2PcOgcE,6<[
S?(bQ;F&BCO69Ce@cSe\VAF^b=NcOVb[X]7HAQC:M/[V,[<WI,EJ7:C4-gf-38[4
77T1^I23H6e1]@95IG<Kae-fVJ_-LdN.a#eRGaU23X-8;g^/^@__d1G>#.egDVKK
I[O7G3CcC.4JX4bHe-dST=6eT(b70]/f5)HNV>)&8D_Q40-S?Hda5(H<#.0MNF<M
+Uc)BKWQ+KS2?J+YEcW>O)6PPI_g0.ZGA6)_.GCY\M(EEL4610e8.4O,-JJ\A-U2
F[dfE]:C@2Ab]S[d?-gS>][/#L@([ee++b/)6\Ue+/fZgO#N<W54-FSa.B?E-=TC
9@(6Q)d8UV./7#cVV,2Z,WJ2C0L9[>>9A+)^D30ZAag-aAW6AXAM&M#Z??;.&_IJ
fK)\[-,/Ua-?-/^CG5EHM12f(/1&ZORMPM4PNU/D,CM]7=Bd]1H2H]K\1E3O4ZId
H4D23?:+e.21_bH,KY5A;@F-fTK681QIV0\e3aYGREb@VK3<[X<?G<Cg4,-M(PUf
_Q_;:7J13Pb@4],Z4fLX?(6Y<><1;)Z;=a@?3UN:Y^02[bDQd1NMBS+S+7fX#MgF
QWK74_bQ[[O1CF^I5Qg0)TIKALF43K9MX]PSL(7_f;0YJBg#>(DgK+aRT/LAXb5R
S_Q3VC-#[L40@DFRH=).K7S:e@K&Z\?],M5TgQ>-Zd/M?gV+cE(&gNfTEBIPZ:^0
bIJ783ZRO:dV@feT7E9:S?WX,^W>2ET_42:T4UB1f;)1C\1;SA:>--HLAf6Hg\P,
Z5\fD(;/W>?-bQ3)&A2;=JV[L^;1Z[:T^Ma-\I39(.3Q#U+[eR+,5-?QS?WfU785
(O?9)FVO@G#V?=5+PAZdUb=:(NP?&7ER2XX6(-D1BN43?KDK/6908gWPeJLFK7],
:),TQR1:a.B.^fXcR[[AWR&8^&MU9NJF[c@]67e32=dMTMPC?10/LO@8L[g2[?Ec
XJ0PG_bNcST\W;f^752@#&Q2R(fMZ=-P78::f)A\c\Hc.DMeR\K^7&3<OZAG#&L@
Tf:gLXZ2b[L-UEMf+4W+Fb]KB/7Xc96&A(V31(d._2S5c/D:@EJb0Rd#<gQ>fOM7
J/)6gFC&K3>6]\GWEHSE#/GQR_69&>\_SA,gXT[F:\X#RD657_NGEALNK_2VW+.e
a.0@P[TT)[91ANHdXD/[g&YRD@)DfBe[e?0:OYR<cW,Y-:4EX\B/2O_0L>18)6NK
=@KaKHVVA/_GFY=KYc\-2TNK#5_]8Ib-_0+D7:bg>C;?BL#2XC,=?A#)b8G(&THf
OV28QW]\Z1dEU(MGBYD+)7bTNRSG/?\V0R?H-&1cG(J?\6f\;@+[\V?4Q;>XDA[e
&GIZ]P@]M[Pc4_1#[LT[,_/SVf7G,NRJgaY4T2/#I1d-.ZX@E7/Ob;2b_&9;,A;#
T49XZ3:P<Hgc@fA94eaC\N;)K^a&#-?gYGE5I4@VFDYPcGBgL]VaU[5[P-NSNc8f
BgBF8]GCKbQ:HUQUOYNE_a7Y:0RZC=#[VY6>X:ba1.,=XJ_Ee1EFAX=3UT+g[1Y@
>aJE(<X7A-8AF-:=d/AN)2CVAN+5P?YIbV2GLMGDQEU@cZb>M\Y7OV@L<^Z-dEF3
[?<&b33ZVK_bMM;\PTdd=,9^G916NFb:E7f^#[cV#?gPI[,egK__,]#Bf/cc&3T.
0;#bUIR:[,&K7<J?U84-J96(((OCD)^V=T^]FeC3]\5dHL9GMA9U:LV;aDV,D0e;
Rc.2ET<Q7@Y+#8]0Se42dPGDRc+,S0;PWB+@gQ0OBa&\ZGV[Z_VUW_SB[Z8?K1d[
dbGGGg^f)VWXgS<Z,01QIXH>^#Se_0L[FD-4WXRCBG_S3ecd:(&b;LMA_)#)^ZaL
Z0_>-2B1)(C,F+?</CQJdC,2\+bTe,:\QY?;:4EJ8Y&A;I?3(55c:g#8\W>M[b^[
;TAG>S?B,ER\e^c6:9#2,RHE2KR@98=g7SI=HMG?1fJ9K/^eN@OH_MgcLR8+Mcf#
b(N@dM;:XHNH12c:Df@3RW@5#TOH.3g-cQga;1W,/ZX(NENd(2/>8JR8N[W?H:SO
.74<gL99)<7;SA<_C\SBT]X:]C.Ef)f[;EMVe2?GE@_a_.cDP^>YVdA&0daJOHU+
5P_UeK<(EfgRCId>d>@AfCaRf9E+RV;83Y.PK1T54:2<,=;RBAND\AXbf((A9;b4
PLUV9_-@0fe3W:H@<EOCH[XY#&(T>e+>TVL+d8_^e=HJ/-\C0;-?;,;fe?TFbBEH
>>eTHaN&#.<+[>PEf)@M[VBN=<GMEP7b<+XKN#a+OL5?N+&N.0A^I(,J]4SY4G4b
2BT2_5?N^-:Cf(AKSOWE-^7(N)2[S8S^NLVC=8HfOT[RB<^=MU2FH,VNCV1d0]a4
20E3O@?SZ@M.HX4EFQ5?UTa\G6:[e??NF-YBcCQFWJ0:;:(PM4YJb/,4DCd297VW
8T7SDIQ=Ba(L^D;#I;D_)^W-BL5f[04PI)O(L0.(QV/TZMa\G_&W\O5EYbgDfZ.D
f1Nf^N>46(f7NDXb:X::C&FWI+Vb,YLQ#5BS7/gK3U+DfZV_5U8@f>DAR:P0(7D>
>RE?)G]SbRH:6C\Vd&L[g>.()&UBA5;bADaC^D,IBE(ZXFe2+bWVK?O&?0/62e<H
3LfE.8P^=4U:Z2Ec=?VGee]/<5/)T_@^WUKBR88Y_H2;Of?g&@7dgd0fL\6K.:)M
CCW)b24-1N;5D^-RSf3EA\][KD:Jb5g?>A_GG:>T4TWPFZF[[[@Jd-7_-.H(f[DT
O:If+YI:bCQA(aFG(2c<,Y<RFOXfG0@+930f8fNU)+&;COQPe<X_+U=R9^.5UZP?
S.OgNF56&J(d_#B#B9B_+OY0EJ+X3;>F;fc,LdeG35EKG[QgJ6#RF3FH>cWS;(6#
:.A:(<FMXb4TAEU#K._)#ANAYE&N(T,0XOSdc2g64UZTSP[RKEV(@.G4IJbga=\>
^,)CKf<_[FdPVP5V_L^#^]Xgg@-L-0@].[Z@,a8@N8KE#I8ESP72YRBUZ;=fS<C]
_^bWO<RXCY(3L<B,;;C<\UK>19_^E##-b92M=a/X-Ed<U@c_0\S2dAYg;(b3<P2W
L[=W<@EMME2]8^dc)+Q5=<)1(;EYX>:7I?A--;fF=6.OfF=?.7J+0b/Ca1:DfR^4
H:308g#O_QF(DQKJ4a4^^(gSPKeL>K<-T&6I_>=Sb@908<2[?EW@D&cRb/5,2WR0
P]R8<=WL_=(,UBg1H3BZ/PQW-He,N)K;&KPfQ,g4L0=O?=AB@eGZBL-0#2^P?U>b
PfcNJf3ZRLS]0e2W8SU1gLD;.(?&S82]?[aRGG(]Ra1#XT<1;:2b<CgL1VX9Q.Cb
VQTD)e-[WFKb3H,JDNWCSM<=-KXF#5@T0b3J<AEWaRU]KR?32VcF6T/g9&+74.BO
^-(Y;8N_g3R@[=>1F\D_\g#,^f0e\OY^K?b.R&J\75_O7\>@]NQ?@RB+E++A4/N@
BKEMK_;9=,=P-;_OQR[1,agS?NO?E.\.+ZJV^,0QZ9fCVTDW_4CYgOag]<?47J#G
TZ,&9H&VF8Ra4#;]-05LE8U@>a<&Vg5[]BX[MP7FE0B+JPOAQ6bdE)H39L&cC+7(
E8;M.??Y@Y1O@G@beSYA(F?J#fB7.gHMWL(R3=-SfMN+L@B95T4/cO@W4dXL\a80
X^5]c[GQL=5<X;(6GNDQJKIfgDY,SUN@dSP[^]dbK7H-d^7^<OVXa1>R.)]Bf=DT
d]3I9>WGQQ5<A>B,ZE+.EP\&M#WD?/N<CFcN+:TQEUP-/,F6I_:#E2=@+5TDe0D_
cCHe.SWHIU+RQA)c&WWQL&\7T)5H+e53XFZ2]#1@/7Ngf>=.._[?RIP4<CA;O\EE
_[N>3aSSc8c2H+V026Md699@;A]f+a=;?]T7-7aWgH?/A;AUKa)Z4g:D_^U&/(6+
EQB-<ZF22_LVZ,-N<6>L461>=e?]DI4.T6/F@6g=[]Q<ac4=PeQ+V?JEA7<BZ:ZU
FGB4&3/7L^7V6b#<DHd]F43/28B<?F@Ic34KE+(/aL)GTX9g=8&>WE;;V3P@dS?/
X<;c40g^XRY+_POSa0d^-^eS+_6TgVU]--\BIK/N\D;F0-0\]H+3I??J6a<\>U?.
(50dN)C1ROWNR4_cHKTVed:[0fJBc]]AU@UHD7=X=\IA?H7\3De5V(FE=CZVSd,6
P?P6K/.OLVRJ.NTE9\,K6/I-dHH^+]N=(.:T+>OYC:B5EA^g9Z;BS?E,MO;6MZXg
+FG9Q+O:&a3V)EcV30\H(6gHg^3;1)6MRdUGECL7XIb]cOa@5H=d=YV@4#<Xdb8S
YJRUcVPe:IQ#D(MQ&)g#f(Z+ZWb-ac72-Z]b1P]S@S&\CREA5G.MIcIAI1)aS]4L
gb>7@,K(DDVeeXKb]<5ZXCYLGg6eQ4Y(:QK6)9B_b)/9B&KaUaa[T.T94UbOc^OJ
R^9:C65=RY>f:^9D2H.YX;0GNeae=M<8T^U8ROd4]8STQ6\5_B7/6:9>fCD+]0QN
HX,[(&HU#&<S7)+^ZZF&Y&E5\Z#9&f.N&Pc-T1Y@\K.A3.5+11>dE:eGUE6Q^ba=
IA<(=dU1AYJ>L>Jf)cVL1I(4&^JdQXCQWUPYV5Q3:H0<cU7PW.\;+1@^WK?8fcg\
^(ZD7ALeP:1MP13LAD]0[T@W6H,Y0dS(ID_b;^Y;(ZJL-e&3OOOdbQQTBWGaT,RM
6N?A50.?#F[P@A_a=1GV&)a>WI8_CR)]KE\:WIb(1&ZaOeLe3@Cg.N+:3fRg)ZAJ
.b6C^XA=^\Je=V@b/S?UG(1=]FVcIcQ-dfRF>\W##8g3OU)eLT\N^0eOOV@N++<#
O,K[6,4-.FL..R]6dU.,6&C2&H8D?^WGV\#SY;&_LG++;GW7Y&BM,eW^20+LI3fG
T6T,0Df^.J(=@F2RHG?aE_V1Cb)b@ED(fD6GL67eYg@(P^/]K_@gU&.OSMeY.E4N
TcR)#9>#a7XG;GS^a\N8N9/((^\VgLUOH>ZNeX6b2WLR7>0-,5g8gfU/Se?=A(A)
<bO44OV50cgI7B@f_)LGLdR\__aWUa1[\)LLH92B(>aKTE?0QIb4,]1V<)@R,)53
97M-:GTQ#D4<.F@>E\GY^S>[.0PCEKb33&G66,8QW_g8bA._d?:K^WN8R3/(<;B^
84],.9/b5ZSFF6&KC.+0bOd&05?(,\K_DQXd,=2[M.+?([LQB9f<5d\T.7SV?e\a
R:^D2F12KeU]Nc[-79]S&:\4O#<1<TI1X91aM-MS0WB&DIQc]f1TeZ(1IMAGgd\0
[,Gf>ZLRE,QIWYVfFC_MdbCUP_>Q+9CXWQP)2UcK6I0?@QLXJ@#?<=>]O<V#,I+Z
^QE9JbUOW68eEKHbb7Ee4d2;I[Xc:.JEC@cad@GVcI9;6]2,H9:E3584@;7XR4\U
U:;5=,?(E?+)d(I:d4QEWEG//.4W21TaaB1T0f]?We?F>.B/N1UZ[2==C?:9fN)c
BFRF#+,MYA4PFYbWJ2_U71E<V(=)R=UR+5b(b-6J?bEK[_-P^BV)__3g_+;#-K=:
?OC<(+G1QIdB(6.Z1;Gb5>_9M/?d+YKd/HW:EULT&R]MGL&[&..)]0.56KU1?BfY
\[UP#):;WEcK/<Ag+&dUI0bV205(46aZfDL13,gN(:-c>L[g@g<^/O.R4YZ._FXd
0X[aEW#2g;R[#bTWWA4G,_Hf\fe#AfA?,\.G-=-VEV@C[82?5fFgN+cI9I/g>FJE
Z_T,U,PI129E;_G(/g@[90<g@;4R_4aM6DDW^(Odc#/FcS\bSAfT<]>0[:=</R97
\XM+[K6H_N#DQ7T4a1Y#7f][47c6a(J4BbHYFfYPH&0@5>#fe\a:9@MbNUD[<WHV
4a2a[&.B]EY3GY6]8A=9ZP&(gSV#:Q+#dVOVQP\0#5&#OgMcgPL:S#KE/^HAG&IK
G[P]6DM)Ub1)V@G;1Y@FG(8(>cZN_4HK,22@#2LMN4<_2Y.a@?7;Kc;1:YQ^CI)e
L@Sg4&GKb]71C//Hg#TXTd2)/@J:eZM#R#\)M0eI10KIK1.CcOL7La[d53N\+^+b
X4.?I=;3g?cN^B>N/,X6060aX.NV1RLPF^.-94gV47b]ZI7aV0RD75\^P6:?+?^R
D0_d68Oa38;PZ^G>41@O?Wc5EVJa?)01#2[:OI]@cQe9?PA9KgCDY5PG/8D^F.65
9)VdL)AS_gZ/,(_AQ^U8,UA1g\?457_K/9T&S^Q@X[V1fDA=TWIX@8HNNB6Zac;?
&L@gR<[,2L71]1cL#)\(9[BBQ+2?P40gR..:N9K+;RAKF6;X:XRFf33FJ)L;+.;P
5HSa<<H6S_28RYYW>Dbb_YIPWHZ@3ZDT-?90EVX;DJ74[[BO3=QVF38\6;g?V=3?
1e-Be[fQN/<_9e-SIaIR86]>;R9#[[I,fJE5e2-FXRUdc^85=TI@-ZB(-UBH;RdT
>H.MM&;9(;9;,])G6U\8I6>U+L_&)EVMYE[DV52fg2/M0SV^+ffaS,0ZLBeWQX@R
3^DGT5fW^8M&4E719=8-N=YS_0bQ/K-c1^YEaeb>B#;K@E/#>Ic>@/C-@e7,dX?J
Z:0c-AGf/5d_^E-e&<OT.ADBA/P^6G6>2ULTL<[Z)@P,OUFO/E,LH::K2Q9PX8QZ
F5Ya7?DdU7X\&ZM7GcW7=0/&->X[/@PED+=65eE+]<RSOK-eC>f[4a6ddU[\Ig)Z
Ba9Z/Ed\;NU[Q/eI7fYVGR;\[4057#]3(S/H#F8d?I(=R>9>>AbYdR1e]M,@S\6.
OB)^ELb/HQPC[>F;()3WU0@Kbg>g7HA642PgC@T68L0Z@D73)7H&d=KET0:NfbHI
cQO6R@NC]HH<9/<QC\-G3dcRD&<aeCFPZ[[E2fP6V[e^WR3D(HW1#-XZN&2;RB;g
=D4Y7DS6.O;S@P1I>Z/a9KQNIW-N6Yg7I6\;Nf_E.@N+I?S0AYa+gOcf#0?D5O.?
UG=PM:Y<a:_Jc13TEZ8LV-0]JbZOY@gLbR95\R.414gf6a<:?LB,>>DCQ,(S8f>/
(1S[0D?\,=aJDbEQ@eV4FJad8W]K_VPELg:\cO2g?FF6@TZdK799[5?OLE[W+]X5
DB7-9RQG&6Pa2><OWa3D2e]Y/)&A3)KCYgfN_P/]BT^3/.BY5K;J^)e>C7.P0C,9
S>(AE:X(7/aePde]aFTR(&+_+#Vf6^bY6A;7BO6PXH[7XM^0PS[O#;]9+J&N2Z_S
I]JIL_/ODIHD4[+8T)-L5Z<11&ZVaB?[gO81)6f.KT=XfQdM4?0GHFFAOV7Y,;/;
&H5H-F5M.HA=J31]]LFI(ZS13R+8G,BTI<+))JHX.EgbN_c0Sba+]KPTK_5M0XL[
(1ZQ5VM=,PD^AT]PgN-HI-,2L@]9EA_2U=8/CK9\&-?E<b/IeON3f^N5\Dc6)aQZ
>Z>M2JP<&1SQ]b#+^VQ?K2\2f6_QO)Y:T7YGMV4eADF@PA1e1BLTHJ8WF4f.aG_]
OF0/,Z4ad&42(C+Y)TGIKT&IUef<c@dc\ABVYWHTTc-#;=F_V+@dA30J-RF.2NB7
F8Hc=,aK;Y9?VR;,DUe?@fBDQMS[,?DC<<(NM79Q&;8^,135MB(TN+a:.6ffcf3E
Y5VdH@5LSI#T20?XYc2M\M;eF/O[JJcC^7-R7BG[>[]N:73=9R^=^(^N_:VP=(6E
MZceO#S+ZZJ3QR#K-c-ag[e(9aHBKQ+eSZ^e@&2>F1Q#CLa&c,\8U^_(7HReHB3g
Gc.D7-CSX4f3..JTUMP].&PW=PW+.f9F]]1CP4(gQ44X#1c_CTRJ7Wb8g#BGS(Fa
DJ[VK6V:4X8=^W>R+-<[OB;>L_6=f^1a:I.;P:7P<MIL;AV\V@4_L[K]EK)SHI/(
eIf=SL)^&5b69Q?.-@9MVb]1HPK?GG]\]P0VEW3QDF6f3WIF?fB45I\OWL@K===d
V0.>=JQ5^S&([TET>Y&6Y6[Oc^V(-(>b)LeCeB:&\FWg8^[H#A#LBE<V3.:>P)6Z
2-g[DOM0L\RbL#dcE=DIT9HW6+X##9Hb^G[d\APe[Y9;Y8MP3?9f;&a?O]9gC51/
6F?(S?>TRI(OH]6@#IU@b=YP1C]N,WI-L?e3CGTL9fA,_@Y\]1>P8b-Bg?H1>]UF
:Q)#+eQ9e&LCV3IDW-+fW:D.c(<d6_&(@gOD//S._6V7,,,@Z(&W6[OY@7+]692>
@K1003#QY=Ic,V5P6OdRTPfSgB4+Ug+SDRPU_R-&M#_+M?@TX5<6PIV^f>>BH)Uf
SUMf/.e19/g5Y#;4=JQ[[VTR>;D(.D=eH)_/(K,V)JfGbd>?:CgEKZ(JX0DM3R\O
/)-FY@K1L[-?<3WAWbOZ):FINSQZ[X^FSSV^0@8I=[1g.+&A&4McSBEGC0f23NG@
OCBE3&fP8RfQE0D<?HDB72?>L_J(B7PUK3Z81FZ:OFZ#]F@dF][a.=#(b1?5X8aL
&QE;BeS5T24I(fgMUPCY=NC@2X>I5gb>d\;NL1H.AQ5a6_gJW[;_;]464#DVPSW@
9V1d>\Ba()QXK:QZ,QDZ.YD\?_ceeP5AgJKWGaUZeMXLL6)=5_?Ga>FY;G>&WfcP
>Q[C:6^X^U2HK\2G3#O[BYa@.=@R)>f:5^Sc/PGebf\aL382SFR):W]3P8U;;>/R
\F:?F+R41a-Q#1:Y+./:fEQe:4b\?)\10/G,eGJ?aA+cVd]PJLA,a7fBU0L+/7U7
<YM_GCUE-,eS;41@FFdeE&B&1GM9A^:IZ]SG\+0Ed_S2.@<UEDELGcL:ae47?_gN
LO,R[NEfG-P[AE)D3/5/@)6F8aLTeQ_+6I:YA)DQBb&CU\I_?JG6CP<-H^9[:c2C
\5YaT)S6\e.O.6HVI03g1c1PU>79VR3.bZU=OILO^Q5g>V(.?Ua-W)1Rd\<bJB+D
c&>XNJ\>.1PaQE@[2>?V3;7V9bM4IVZ5GRdI7cS1K^NK5TdgGKa-N)efC4)FFPDTR$
`endprotected


`endif // GUARD_SVT_AXI_SYSTEM_MONITOR_OVM_SV


