`ifndef TB_MACROS__SVH
`define TB_MACROS__SVH

    import uvm_pkg :: *;
    `include "uvm_macros.svh"
    `define DMA_WIDTH 64

`endif 
