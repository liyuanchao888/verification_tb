
`ifndef GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV
`define GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV

/**
 *  Slave monitor callback class contains the callback methods called by the
 *  slave monitor component.
 */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_slave_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_slave_monitor_callback extends svt_callback;
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_slave_monitor_callback");
`endif

  //----------------------------------------------------------------------------
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
LxUSvFCdI5t6SdHzY3Y7f2DffbYzk9pFPK+La7zWMOF6rtECZ4XR4BOJKKBJWuaK
EPr1D0+FFhPM1GQ7mXYqIXWHwCy5BarAQep8BdSNuBAHncjJsBGVHDXb28rh5vn5
iWAXmybp66PUpeGU5juPEs/hmFLvHQiENyZFObX2f3E=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 7641      )
oulPUMuXBcVRVj2IaofCjAX/EEfss1VbowPFJUlAxbE7yjM+LtKOW6wfdc0kscUB
/dTTfpUgn5Z7cZMs8zpyRd8egsvxb2ygQAPv8zZpTwk9Hy8+fTPW1lqrWbkRjizc
yPP0cIUCBdILJElgcLX9U7Axd4Prquazgwc5oAcwT6f6r7XL2KWt6e/eWoekXeWp
h+EqD0FKYJE72lZXLitCGLBRKUOKbASOR0mpGvPI8C8gWg+04+flWftcjnKtjKQy
z5FeuHO7M1a+6cFUffStFhylhK20VyC14msgjnN+aIwmfVU0Ubv6rGPAsYL/+lFr
S1X/JeETiYOm6Uzz1B/DNmSf12cq07tPpUJg7aNffQB8CGEMGJCzQ34+PsEKbaCA
gJe6h8vPKsp4/ML+S09XRajlZjSSOxYL0SE4Mis+DAXod3HGszxZ5U/BWercNkVR
gIAEvR/zZm7bzquqKn1KCF/He+eo9H4GRPS0Le4FqYrfbbWvfx8WRlbNBr8/6ndN
PwtQPHpH7sGkrjFW6yamiNZVBOM4Pdy+C0P3sA1ZkmoXBOTTVMYsqKjL7nPq1dIp
q+Jle2kmJStu0fGcdI+Zr9rpVAbI/ODhubnV4JDU5afYrFSdhF6oEkpMsZmd+/wU
ILl7dxJQYlUurP+LxFJsH2pIcLiCX2izwrj7D7Evf8UDL9l2OflRP/BLhrYP5bMP
cPiOSXYubQrTYaVpvxtNe5jyHkgweH4CG8abGwlXYW8bdIpRYz9Gv+IvOrjkqbOz
FfTnUik6XNemhXUnSVuGNVsDpL5wzDRrD7dR0dck9PW4ZboFhlcxw+P9DDcm3URP
pfXwEW63HxQrg5Y4Kkb3wl5UaX6g80BSkoqUHwmp/3crRRVqN31KNaTTgJLfqT9W
rWxNQABBgpC86XQaxPJf6Yg5zLQdDdIyPOjOoukmCzSvnkza+j69jbQmlqV+8LyK
HtPEnqzPNorPhhWXKiybkhI5sINs261Arap3meCQCItEcsSR4l7Tm/NdLZU2t9kB
el2XGnwgl6sjeHdujugr1CJ/yIRywo5g/KgLY3JjUlD+k3jMNV2pISNq118c2jDm
FlWOjCJ5iM09s3y8NApqGQzXK007zg5p+aicfChAw6XNp5UfG9Gl/9qsBdzF4qSZ
00fphDXv6vKIGwN1ACUmo/EghNtYCBMqqFcaQjUZ5/rVn0iKrjsMqDgCdWDI8KeR
odFmro4qSZwhaEH/m2FKIVm3m/N6fL9+2YuJ902Z3UikWJ7y1B4ENvx7ycoNWARL
szwKYTWen25gj81wBSDcF0r0QQbWs/fHkAr53xpBB1Gm4ct+6CRbIG2TzfBPzydp
YS9mcIZl/ZzswrbyLefOuTDzCCfvbhCFH9tUdtvznu749ymv+aDyRkPSiEnKfcRI
uZUWmoqdWSORcxJTIHvjut4f+D/JeZcQN1Ev5DdluPrE9q/ZYrgP5/AaLuxuokBN
J47AhqD4Bo7PdbFtp3JnouIhCNWm8e+6N2iNX0PU5VaQeHNkgiyLl7Dl2h2IeOnP
3JZffkHRCOQlgWVFp0RAtIRK3z9hZEgo5vqxYYmObjd7jjB4CpzQUZRtBQ5YpZQD
tmFnL/cgP6Y0svrMARLceI1UC3/XsjzbzvaC0SNgSAl9Y5Hj1Re/9bP4vIGE3HkC
y2FL/X1FrrzKfubYbTlhLOKa+gYl8stiArCOXSHcpmLJh0HLHpaqH1OFyIPIo6lI
ZzllLRa5JDiMAtpko+Z0PXzwvWFz18IQvzHIm45VXurjwQ2yWnu6TQqGl3/Q7Ngz
Rpn+6RDoRs+Br3P3ulbL7YvbzUalOKaMtWPGrDGFiYxk4ca4uJC8Bj4GvgAQTmP7
jbnrpG9dN054t/5GxTPzQOw79yYV2WEK/sTS4WOIhvBlko7Se5GCBjMbydh8qH/A
TQMx5BvTTY+2wFNlPoG7QaeDXEC+45QLbR3dClX7Gemd1T5mrB9kH3kDGQblXSj0
3AhJRASnJVcpFdgqMT4HhhKffm+yGQQsfAJb19bqyzM5Spc1Z+nKgaCY/u4mfMSg
neRNv7J74EOV47qVfITOonJCTWBWLLNiSnsTjvSG7lGE/1GLg3Yi/IFWj+7Bg0Uw
QXXz5/PDLANSSPcSn8UVi/gQQ6ZawiYtfX+RNHpu7DRekQLMClj3RjlhATkryoMZ
3hx06Dg5PFB5OVW0LPhPADTeOR+xenJirbi1PwKcqFe84Uz898nHux1lKP6uTMO9
/wJADjIVxVfbgDoiqNMHPlyDKfaLAPilPlEQkqeQzf0R8zxG/JvwRGOOBiGEZJ5p
CKMUUjiWZyYOnr16Xn3K34u5shZ7cN9D4ud7mU5pHZHHiJYC/63SHHqnZS/Exe8R
WHDGU/Lu32kFvB+JgUpr4oryNsFhNQcLxqYkqNrJicLA8MpZyvBA0PQxSItU9bdZ
U+RH57Z2mepGO2XXOV29AskH2imxmBxnERuT3ioytO66/iQtjwVuEQkqQsCA7tmu
/y1WnBM97YYE6iqmlkO6db+IDMiwyhbkbRCmk1j5pbmdJ2Q+yGTkKy8GTaHQlvrY
OGHiI8EyeCjZjtf23FFpeLUQM/v01wCQqRUAR4DosSsMtH8HWsFFMtSdPc1qoOto
LM/ixZhntyghWdxUpnbNeM5y+YxgEtCKd5YoCfwohV8RHKByvmAgPDeo2cfoGpAN
z6ghwSl+CTBVTIVfPGQQWHYNlMfGgFSgmJzeD0EnSzIrzjiLO6pwXmUvt31dnloQ
L1BG4WhVp6ylOOAxeJ4J3T6i5/UrFaXEtenPQIYB7KEeWhVdUDz0Ub/gDzZscPYb
IH7nxrEoDv3y1PmjFZeg4THbL+X0Y12szIf30OQEUxJq6e3eDXbtUobQD6D0dssA
KF0FF7suhsmFPh18XFKrQs10RgXqATuXmHnqQ28M9oSmzQjZuNsYU9ru1tKkGivp
Bdp5LcPyAGYpULYcmeYzhHDVvYOPY02K4PONk5tsR8cuh8vEac2Zojf0zUtHvyql
uF949Indl+xAUyqcPCIIlMu2k0V0qn5ZP24doqSmu6apYDGHq2J4h3bPjQod73Hy
lEBA0rv4VWc/ULOq6TqQTufIVXP5G3A+cTXQbx6r1906hg/i0KTx1pIUE12n4UGG
fNFDOd4pVfRO82wdrqYmHYhK/r9EBSfaCtg/VzfjUo0J77xSKmXhC7mAuaoQazKN
eXkB+raCgtVTDYGqi+/uDbwUSYqWpjDG9FvRGmCjY4IPCcDanUv+WlxdFALJkhF7
0n6QUwKTk+HzjDkCaJBg94HkATzX+iAKr2WDTcl196dHTHY8I/K3LdP3okVfGSL7
CO47TF2GDnkkXz/9+86QcLxteF3c4V9B/w83S1MYGNccI6O2F07tUK3otyHan+xF
Wu+nViM/1dlvjgVftflgdWCEnqhWoUyoaMOZ7aPr41QWH6akAkZ+y8NDwTgyrdZA
q4Rf8JVxYwz1F0Y0bQU36DUYwpsU2CQq90HM3hEQNtCZ96QuTu7/bYINCsMeQRtB
nNdZCUd/P5jG6NA9vjoHwHNudcSOUaK1VNpd6PL5oE/h2np74Luv2kwKv6sOH+gz
Cxmz5rzEpYnwRO0Ko9g3yK9mMtekivkcoudmLWzKDTsAwVCi61lc5faDdF+BB6Bz
a0kxV1wQwPvYjBuDWJlGxBuBBNt2bL8eWnuakbQHNIfPGkKcx1ZFxUz2rngoWBvA
Ksbsb4h+N8Zsxa9c4b2e3J2hxDEXwn/w4gTRmMNh5D92C6PqyjKYm8hS+3EckNz4
56cqcWWTAcSiXXeb9iBNXGakU8eS43rTwvY+CtL6+7Ud6Y70oD2IGfZySiXFs1+0
csyLmNeUW74bx7q1ITUX1rnmMaVwDim8eAhtnzP9zFyfDN+W/ACBdq928KafZav9
W3iO/+oJ6OkWduY5NZ4EfLzvt63fjxmSQSMJ3j8dbBYkcQik7wQx9gMICeITm3sJ
+TSZW+9sZbJrEu6tlXvZoR8YNJsTSKPg+u5qpuoWoeIJjDGn3q1PZpCJzcBP2avg
EfudIcr5hriPlsq854Yyuz1P4OqJWNennPiJIM9jxQ1OUvbI/GsRfOADs2fjljOa
4CqOY7CanFid7Fbpb6Bd5m/SbwMd+ka3XP5qkvgjlWmwOIKBrLNqWwYHhNxUzygE
wxiw7jANTedYx/TMhyhmoXA0YVIv/XV04o6qSzHfNKPDw434RXQcftUnnH74U/gv
Fc0/FFx+68NqUAMku3y5xQBlBqLdEvPEg85FB93i+V0mGMQW4W9Fvi8yGQCGCQzt
Mpby9bNbM7kQAuVv8C6nLcVwWs37RF0lGJR0u9vWqvglC1HqcGf66In0pPQiuIrM
u1Iamgz0ielL/CpON38TGxCj5ZpLUFRX7+91DV7UyIae7IkubIwKnS8HO8OZ2Q08
qCY5ZfT5vj+HFy2q0kp87xfjXnjif/Mvq64tKg6NyeiV3b7oS4Z6u3XBCHCpj6Yk
sxgCaK57utqMh26qIvw35RJZ32aaAfb1/PZqLfSrW4nOG+RiL1TLA8FPF057AX7o
Wq9Z9W3/K5Ed9sERDxap15rZuP8IoIlQ5EejPY5Ou2PFGVA8+AzOxFkCqTJkLo2c
GlIrw+Quhvg4fqhAkdt9DYrdZ+Epg142zl1wa2+CKL8rvaINsExFrkCrpcpeVKdp
IyY+UQB7oB0+X/U+H2+/urGoGCd/FIDtK18Hr2HouxDtRdV0TXZlRuTOQnfs105g
KqVhqNa2Dw1oVyCnKbiv6/VLYfe5TeqQQVCcA/01/siSWBZHQvqT5ZlW9bBThteh
jZUwc0fGr/5dBaZRL6Geno4gM0rDVQDy7u9UuTNweQxs74Rqw214EYE+WwwTMZor
sRSPgxJuDVSVteFbkLmofN+FQY25XLqvwm2kbqZ80NlvXtScShWbwpgQCV+6grNj
AyMvF49WGlarUe+bO8NS0R7u+3ohhlHU32/H0JqnVZe5k8g+Hjib1bzDBxYYdqX6
FDZ7ufDrdmWI/6V2ZGMYpEevUHLfiIx8aohKMaA5bmXtaAmupMQ70g3zwHBq98/3
xrslQ0Mh/JiUUAuqcaXCyHnpxNyAMceAUk5GF4nheLer/+0gPOx6woP2pl2iDUg1
PUeQRFNQPB3AXfK6woqg6kDOg5alEc1iXPUjq6S4Lub+haQVZmuN3ZJU+NuwFXx9
5uOZrJU901hIIo/rQ3g5mxdPM5+DGc7W6btSrnee3IDco3fa8yeQvAz9uWv7hL88
gAylLY5buL4ThWrq2ybV7ryj2peAHPe1nkGqanSqpX+/HA8x3bMKEvMqLok9oEgZ
q4s1bamjk906x6I/EzdklXEkrmECI9Cg8v9e5czdF7Qk/Er2mUP4JlJMrPP0MndC
+sq4FpDCdya6lYCe8cDcJTbq83da+j65TtLouObWMfHv5mJlW2/Zv/zHLVK6ITpy
m4KeJKB6n7EcPl9rlkshLExQK+xycXwUT5zGfWIBc06LJUm00hOG1B3iuwssvbuw
f4Qv7gK6AMZdv76KzmZ0P3YK+ymTZAW4Y0VDF4R6K1ZFPqtMSuO8i1eZd0xFHitL
/f1z5+c+1Oz7ZqmBsN2Aoke14Bi0FW2ci7ISn7amBScmT0DEUQBgHw/ANAo/hhhk
+EK6BXjpANZpyiuecV0rwwVPcEZDeA1k+UW1QJ+BzIJTDoBMGG/wnP2EbDXfpS+y
1SOZOm4JplvIBn7wg5tZbh2KthgxP4I4R2i/pPFj38qAk33EH/DB1i92e+yt5HNS
k4KGN1s0rRHNoBa0v0TQs7YRl4J42T7lVNPZc7JkAkSqH6FwpRkIIeB3iVglLncR
3MGYaWSAgd6CSw+/2C/Me6w3iF58uKEFYWmm4raW4prZGEZseZSPXDpcbbskoDjj
IJqFyNQVqGJNR7BL+b7cVg6z8w7AmyFcimoS1FGncvjwf0fkpyGyAifE1raV2rxn
qvSBHpT4S2kzcLDtLd4u8/jXkmvFtG5wUi8d7fLBcd1/T6oyINHfyKSDU5oZyGHQ
t3CHPr8+E+zgfKuOu0/fNLFkmNmBRpubEWVyQu7g8MlftBFH2JwpsYt+S1NFdEb+
A6/KG8hmBiHtZCM3GfEx0PJNYWNixPq4yONQiUZOjkZSppV7X0x2+qS/R21Z8rGi
l8gHYn7EqBMzO1Da3cbAcI2ohy0z075r0dduFavjIfa0GeHQAXtugyKb32AHutJ7
3WZIkvGDc24rIJkAv98zibJmWp3dg3NAKJYtNHJWsJLBjYGYE7Jwoasfrkbyuw7u
saOAH8VtoxDj4sovKV+ETJLVU3pf/EpDKKlTRH0W3VIB0cuWmOtqyMIw246XCORF
drriZhh0ooSd9CDjNbJW0+wG6sQfYbcJf6s4vJNfAHh6zQMaJRW3VT0X96aWg6JO
a2MV9hNkkdthZBd8u6FXH/PRCxrg8ZWEwKt1JoDR1WKtyUehscf9x9f6l1GKZ5n0
u9Q4ZM7iDtduO2dmRTsPLY2eprYTTgw2QU/KlhpWj5uoCvo9cAA1gmuozxMVN4lJ
H7Jcw7rDGIZ1H6jDE740Uz2er0hTX123UIyxEcFKMZ3x3UqQhdE0e34OCHP8pQHZ
5Z1pEFpheiNDc0lRXNmsN4sIaPMvZ1jzSBVD+oT63Z9qxdRu687+AySWbVMBB95X
p3K/L2R/xjiKfVzyWSNgV5cADa/CZX35jbR21BwsEC5QIeJT9j8Ksu+RytA+OuxV
V3nfix9X7GsXWnsN4Wq8SbRstFgijE7Oo1cG3cQhRcXiTvumWeL+jTz58VwtR3Cw
tp+WPiJ27+x7PZdnKrrRYkswSEdMijyR7PrIij28OP8OC9eogsD/rUfM0wLr2keq
X1Ugn8ZifptO1UcWJ6FMbAC9kIadml4jXN3322QpABEkKKcLMeGvuln7oXf5STl7
9VJeI1hWzRGb3y7pXK8NUXm0xp4edlN69dfjVFceL5150SJSeQ6mRkvc7YBvO5mS
TbLCex/bRsZjAxInY1ZVqoXqQ2FkU5GP+mIBTP0XJAThF1Sx618siyRuPl3oWfLM
ak99L6WtAnGha/TaouqeiUpa558GpwblAyTmOLgZjqAZ/pp43r1z7CJZi3knTlcN
vR4mwxrHEsRPPxrVMW7OkrK3KCnzFGYJPplAd8yuEkwt5DPGpBIQz1UuFHyph4vq
V5KHbiAtElTlkRoOS+L04ZZQSN4PthN4K/quWQRoaxJZwvRvaIObHyCIlFLaGlZK
Scy3GbfnmzwANMRR9gQQp+9KcKyPJmP9YtM11LVhWAj4sybvGaAhYPE5BHhvwglQ
3PWlYShkZgC8gYFVLcewDecBk3kWJw5dnRA5XiR6onFD8JewYnvIk1pIiPvvPqC/
4al5ihqfPnLka/p5LZsDu2nsR6fOxdRRDrXgPhWGQkb+OwxEXVGvyCu7MdYPRKSe
aFb8yV84RZotQcLV4mlseOsUb96WJ3rijGnIpn2ZhWJJF2Aa9NHVpN4kcWL7MneD
SXJoVvoZYxwRqesF/dY8b8szqlEwoqWpABgdSbM4+IfXC3GFKVzJYWOxxYbJywuH
sG3YbePFGwRyq81wuM1aeCWUj2ySUTPxlazkaEiHh5rqvHShwAf3bpP6QfeboHPp
iLdIvZFNfhzy4OeZ9YcEtPFfP3SRCnLhSD07DEfoxZlr9V17EhxYWEC68G1a1Asa
VlI7gNz7fq1TIe6l9TLtnlnYeXQFKYD7qU6yViU9HSh8p4DBIi0G8VkRSWizT3AW
umAq4x7yl9553/GSai/85Z5L/XKVWI3UewlTBD3i3qEte/lVH+ELSN+WUpN1bAzw
GyGeNvpiRj/5Y28+NlS82UiJi/Lwjk+bXywWWEXn2Oi/Goo4dayQwiObhKYqcul5
tLiHNsVW0P5whrtcDjkBtCaPqab+ZQVarP0U/Kvi4UjwZThgqbHBF0FikceoVr7a
LQxJTIKs5d4NSd0al6j28CAEQfx7wkEHd+XegZin5D6H77QwrmPsoUvmO39IbvRa
IJXlu/z+nljNz0SNC1eW+J5mVywoQJBNus3bYCKubsPiUgwPSAolTiQSxMz5NoRu
D8Bj2pHIq55TmzL7b7jbmCcTHvCdIzPqr1KJU4EqsE5ebzI3ToUdS+hZKOQGmCSm
aq7pzrWI/3j9yEmNHuBT2tERxBqbXordNShMYBOyxuv+6VTWkNbl5/g9cS/SPtmH
p21N62hm3ldXO3fBcntDrL9OIlGFHCBfJvIGVqq8jutaYPErT50ulRJ5bZt+JUtx
TjTWS8nB98xNmNBwO7hIDoXcoo42WDBysgHkh1wpAzu58VJ9Qv2ht/49TfnbfHaM
kTubhZvuJ5lZMRAAtYc/ekXzumR/JOFjt1CJoMYCIJlpsPhDxh+15A/qxi6lnXUy
MFkq/FuCt9UKKDnRmka4D3w069MXt7XjiJt+dq00xtKj4cagb3HjemX3rclW1DWK
PoqP2hrE2xIPyYnlX0vLbiy+dr5Sx0582Kz9q6myXascnrkCenkwWlDfkf199ypK
kyUrx9BjAmrAhIamnkruLWDZ1VrH0D/l3zVIONaaO9ALWLYlPkdCY3EdK4FEUAz1
DIT6sYGLv+s6KK6jH4SQchJIRW2ICCXdeSvp4YM7O9J1OtFP4j78Lhsz9NhCcC63
u1ZXPUbLyKBgI8nDG7RhH3e2jTghVMN2R5SYalwr3MTfGz9F+3XcZklZBgQAGHBt
jnyVABWdfvXpMHtbplpF5Gr8+8mhANye4kMhvodT7e6YfVH56nvU3I83xzuJgw+3
m3S1kiGPX/BWCU20FSqQq8VcXvctjHksvwAeqR6SO3qVeZWph3MM8U4b1srrxn8D
49RpGEtbDue5XG5QSaSIwlXpfI8/KaZvyQ2hvzQbueyJ2RI8nNxQyOptrWdbqrJz
QxIMBo3Y4hYqUu3c9Q04eArwKAeqz53vKBYbaMt2r2G+uALtuBdxInwrHsicNSes
FcvweJK+quxLyDKsJnLv9+xy20EW+dqYsHGuu4x3M6K5XQRX+xn5TW1v3uydph/C
lHJ7Yq5lpaMK+F7nY2nD9s9Uv/TZkJBOMYm6XU/4abP3By1AuDUFQKc6cArQ4tDy
Wz92DKO7QtGYyIPOUZKn9nYtMuUo8oDBC9lHG7heY8pxurvDhq8xjKe9zTgl8cli
71H6j2vPYBo9bOl2L4hUuMUrQc26B0hMsj3CkTjryz0V4jJ/1Kp1BO7dg98aB5Yu
IxFyiIfJv+CpqD/9+8mbL9MW3izUH0XyuytL6+dKHguOZhxmlj5r+W6+jROyGdhp
5//eLDILIFfAsSoW2rxzQkYoq1SEp5ZX/A1InRHB9fvYyose5URJuo6D4HjVsVDh
4teJne2qeMjKb7c+vLQLPehO8cm8Z9Zp6MJU+dLER7VB68VW3sPh/jkIvgXRxW24
vOf6r/6V9k5xh8Gg4a882TsGluNyOo3Btxxqs4YVpRwfSApHbyVxbUDpAJ5Tn9Er
sZRoxa7D5ZmcLowo3OUfjyNJTZoFXQxgnCuk+u/JVWX+yX1JAFLZBmBKl8JciKHe
pE8ywJ1rUiBtgZxwOkF3PkIjxH+m8ogjxSfJ1O5CpMtu4MwuizU2wirrHDQo5Lyr
8plICYXm2kzS0B5q0ovUtebe2hDlO9RdJUqnmgntWtI2S1bbhHTF99wCs045FcC6
5oKY3s0tJ6+BFCByZ0GjWcmrQ06n2+8eLnZI1tvgrN2WG1rYKuvTaIikOx3dQ4nc
nzOamGhD9ffomp0oHdciWcPGZRNJHnHk25u3AGX/WLcelY+FHRI9CSu7zb94HnH8
ifFJzPNSfKBPYBosRK8hMak+P/ijBxjcC3IkurTnVxw0rW1vTEDwV4tt7MAaIGM6
4jDwqnUwuthw4hd6iCNwINZK8wZ/a40LnTSPEgCJeoF9RxpsstVC6lRTvP1Ki5PF
+G1vx/ORbxmFZImGN1w/thlK2OCDN962FIW612QflqpEEBLBDx1MOkGtAfgEDDnJ
qmJQvNnJPGqnOixbewiizZNZhQJyTwO2BuAvIYLAB3SG5CWVl69UIoVroUOKksQv
OI5tp+O+fVoWmAAiBcodFIAtLtJ1/TaDu5URQ3u2KBaMlpO6NREE9DPvS+srOWX0
fiSFbfukzhG0Jt4MNl0uSjGw4XRvcjuUAhfL20R6mQOvH06IIMlhZLAgc9TQw9+E
G4PkLkPXCRzhoA8Ni/REKw==
`pragma protect end_protected
endclass

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KO40rMDdpTtokwbJbOW/iTLURxfoHeRgSPWj8SLcCfTN0aPIsE2CBxQ6LYQYxahW
THsv/zRhSmFHuNZFl9Vs6OmCWZ9YA0TRGJl5plHXbMSUBV5dUmXlZk3ZZCAjfpBJ
Y7vX2nzi1TDxG6znSXpgxOsKYKqYQZr+7O1VIXOyHmg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8040      )
Z1LMjeEZaTUvTdEQW9DEWKja4Z24+GHB5d2McmqCuBMSkmhkV1xC4XwNjcjB5Du1
pNbQFtBsAPShCjs6na2ZHaWmINCN6mfyYQ84pFnohsF5WGtX98evsLcX2eNl0pi2
sby5dxzaal1foteXIHc4boVzdshim65Ww7xENlEHT/GS4er29pXd2cY6kUvjRUpm
9Wt7I/afQJ47kS3lsHwb2irpEaiozJXY4kgNxCnHspeDgVCnXscZ1aQuO9s0JGnl
JDRk3OXpZLNvJbLFzHD2xoqFvhsh7fxVox51ncppeFdH4V3fk6VVJvy0bAh4qRaU
uVYFs+n1/6xbnJM3NLF2pD3arogxmf4NsWEJqeJAzlCIuFrgFv+7zU8ADHTz6YHZ
M8fpI+dly36VsFVHE0kgK8VNgaTC2uODES+rq6nS3z47DrffAdSPIO4UI+R8p2Jc
0g0i5NFSzYvQdLQAqO1ivjXgR8VALYN2JEKh9jmPXUDnWF6+eQSIUaTPcFWMUdtT
yQpk3/cGot8KQmnvsPkINQ==
`pragma protect end_protected

`endif // GUARD_SVT_AHB_SLAVE_MONITOR_CALLBACK_UVM_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
RWip+boicUA3o7jxNMBz9FeUBM5MHtCwvnADOtBG4lR+Aiqtt1pzu722LpQQYLYw
RmRW4Vya8w6nNALi6Xzf/t4qyu0uCLDSHwtizYwAlxV6D1c6K11S4oKSzpRSRf9X
Wpwd36nTxuB92i/QRqzRAu6O8wqSxXqBx0lI608g5uM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 8123      )
iFemlVan5bHFE8CR+PmM8IJ0HmTGUgR3iRANyqeayu8dsEyo8UpZnifypibqCQVl
o3oBXBn17DIAyAiAOZFfaDVtzlAT41IKyFwI/YyEg+Fut7svSuagnXGEwNVhWtpC
`pragma protect end_protected
