
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bj5gL2BNH2b/GcPI5+1zZn5biz5V1BoPNfPlptUNBCt2CmTlYUSl8rJgHhe8b77U
WPn8F4xH2b1m/nXFtJTk6O6C/G0/q+xNrtw2eGNbZ+YUlN6804VhNM0Ag6pPndH3
/v86GB591obk8M/xdYSDou1kBenD67Agu6wqEsaG+q0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14126     )
nk0uvHg7lgtccj6TfytDAgXkaGNmRR1caPQzxfdf206ojqgRa6/dnTTCRa9ecpQw
ah3fAgUKYqSYeYPZ1uh3ci/rKqxHTibNsn/UafceoD9DPO47dMKcuxJc2L1OhFLR
9gARcKs8uYlfGwLnjkUrrn//Vd5HdOED0g4L2RU1s9gH4DriNUJR1UU3CdwYKkPo
idSRj9RXd7DrXQcce2/9K72zoqh6iBcRdPJj1kRhMLiPJKUaWWlY7hjlUcqYTBCj
EZrX21Hs2kgctS3K9EUAeZspkEz/ro3taRENU/2ecDZF240z81ZHc+axpUG/JMYo
itdrBcpPjkVIa3cVuTRq+Kqg0HqwX3GDbE5H49X2lGRYDkpH7xvO5JkHG6JOjoma
61lT1rxHpk2SwvBGzpuuTs/S1OHm8Y6xVKXZ3IkyDuuDP+CwFAs+QzIuxfS9cY0U
wx9Mf3MUS05QN9sp0E2XfbDcfF/sknNp5mS0xCHQwnBh9wOojBB6lLobdn1XT4D7
SlGbZF8YygEOHkfd8dCFceinayACHyStjZsybOqNVh1aiOOm5zDKVpJ5sDQg5QIX
UegaEErWSc50rT9vot7bWvzyckaDgOUzzkj/u/PLUTja6IO2YNTRuKrNNR97vTmT
nipGo+5Jx2bwtYldJQemPQva4w9kqAHCjdqy0emI1q+FnijZTmpnFBAro+O0a19x
Kzpmz94L2a6QZK0IrzanDQ21s/GQ2BtQdu+dmMTChWVgikqhLVm0FqRKT8pWYH42
c4wT3ICMMhA13ekx+iSgtVum+P28ZqkcP795BZua0MNjh6yCm1xU8iQF++oehSkx
iDA9V5Zz/s3w7XMCTis5HLox2isDfH7+k9x+dLJKDVtEO+ios91gmbwxG8uLmXQV
/IPfezZxPJkSPNELIdO87SKcuRuR6sc57ReTXLuvRMsI49U+bo6/Pfar/LVZRIn/
QzeP/zanliMvEPLUDnXnqLDtPgfXvDD7N4Wt6OvRFaO5ojvfOcNcXLsIhwdmQQmN
xwzibI/cqxjeB/UeR3uWF3+4Da/9fCQOGqnmv3CxZxirsg5xYi4gAc8euY2rpV9a
3zw/0t4+OcRPXM6kVpuBiSrQ6NmEtN98leg3lB+3WuTSX1kxi8NJ8npE9ZA0rjzk
rr1/uhUMHYRM3m2U5aaTM1H8koCrde/QJUyG7752zWiJY4adfk9nCve4Xi0amUpQ
PaMFR3xKd2FwN8/CedxqNfFreL1gXa2X+5H4u6V0AUD4G07rfjQ5w/m7lqiv06V4
7Ckq2923omg1HxmeL1f0EPpuI/OHGByZGr0evBeRdjCumEmQWvP4nCH0WZ6Bs7/1
ciAUvfD45m7ywDZhfGHDUfAmxJinjS9Rpcb9spfPyZlLFJipsVOF+S5OZosQgvYR
nBypjAdJpbJw0QJpqECj0RFO3A1hN+PV9r+Wh8j4DSbCXz+NVmaQiDnbyVwPP11Q
ZALc+viC7FOo83u+dLazbQtSqN8RpH3xNjhHGcN77vOM0TwFll1haUy3Xns+Botd
U5CrFIFVNT2KrrnG86peB1cFlV1BwzFkX6N8tXH2BShRmfuV6O2p4ajPoeCX8IgM
bDvpDgAOAPA7VaECLnLiJpxNbFV7S9mvnxZhJYKJZJNbB6xtcpBS+o4t1VaRIgb3
oSGWqq8f+X5m4qjtL7NH5c4jgSQOe204x8fmzteChDM6EPXIQ/f+VOh5+rjQjBou
1JHH+RqSZFOBA/dKmM+6aZceSg0NJyWn7YZMzd9yXK8D95dFUAWTRD9hMS0p+PGj
mOyB8BpmEE7tBc5dEkLGAmUrfoI8J63yBu4kFIZCqHA3TOEQCn/rBXL2oHBPyJYQ
g1oNl3hXgKqD35t37AcKkcpmhDQorpWcZBRd1DXJju98+JGINZv6+61m5N1chdyS
xyhcu02vvtVdxxTgB4f64UaOzE2dz7TTbyRRHB5M59UXRDY5OrctkhkV9o4MjzTT
+nCJs7wqGxwD3yMDp8Q6doccv2NSkb9ykzE3OQFSNkBzdpHGS8WEgGwwLbFNYXiJ
GY4tq/SFPFTCiRuOe1RpKAOb4JZXoPby3m5tY4bmYLdZQtI2vHPc3kiKI3hG4dV2
QkvLTd7klMtoK73g5JZBCKQ00iNq2zywUFyfmovtc+Yn6SEGfNRMRa7m48P6EOUp
VU6bJiy8e1j8BrFWqU9TZHcKZJNU3n0MpHSTOx0oy54oszyqHX+RqLk1ZKTPaiMz
YOvbUYN+dFqmwfQYRi6/IlxnKVJTYsl4UovkBIjkhSh6Sry32o8McigzR+FZ0Xgv
Q4ny1iB7aLNAY0IwlACMARUC3vSi1525+9Kcpa5bsv3aUfGgVQ3KYdSSI/RHHTgw
kYaiSUlvxb6hmkaUQ9eU+UiZ0H5EiuaW1qXoqNBeqeabvSpRlcEj7s5OeqexXAPC
fohGqppd4D9anyKcInkRVADZNH5GILzGrQIdgdxdp2XpjTCNPAHmFDTJg/VXcS2y
cfyHncIy9VsJYVqCNc+7TLXzId6rwuyM/Hfc6Yfr12pZwu3YnnrwL2ypd0pckiva
s+iL7mvxrF5SFprpI9pDVBpNCwLTQRaHRADYH1vllFWnU5gEO2MAuCE5kldL7eLq
TRmIjKMeX9WmJmRZLhGx9pfMrXlV0l60ajEWtYtfhguhko9VZ29jX0OJscix+dxH
P+BxLehGCIP09EnF8jbifaxNrwi7S3sRJXilFGgB8+pTEi23nsN1zUPP9kBdEi9o
TzztSixm+Y3smj0rK7Wk969shdFyyhyKXEJIhZE+D2O2hSLHAJShOO3tLLGtta8Y
9qJuOvxeNYHca/6J6IHkmatfRMqs+dtG3shF5+3ztrsnCaG407zvKbdB+LnVQimA
vlHSIEB14ZWQohOojYIEa/aSzB0yoPKv3mDurlO4ODXq/WXwLQv9SqVr7v17sGh+
uaGZAcdXCb/1pZN/cjTS9lxF9rvL6oXqj1yLdnHAT6bcLm5gO3ZhDRj7bMVPtdtz
wPdVVxS0b1OsmL2s00ujl9QqEEvzOyIvEuM3wS+YEWK77pV471uMyrY/Gvt7pB/S
7h8NjPXl9MeIU01p2Oi30PLtDsmrKBR7suYWLbAivu2taAKLq65+kP+NTmQ31loy
ZCEb7aHAQeR0S2EQyzCK0OCg/r+GanA+aAXExk8aEqESLjv8wEykBuNszW06lwLM
MJC9+gjtyC84yIrrVsdY2N6CmnXWKYCd7kC8XhYIsKybiUBiJJvaiaagJ9XJ6oN3
sFauPNcjNDM+nvQVmkqfULeTDReh8dcw8n6lVT7wuqzblTSSn5IyeUzDV2DcFkio
pXDtL8xNEmQTocaDajDN338LbEijIACIVrsaro2fhsZCJdeJERL1TmlF14SrBNHR
OonydnljN6DnuPffNyE7wWuo+UzjgqVF8+r90E/wzpcVfsfzqWb5oiKGwWfajFfU
htUEk3tHJDIDBhLal15JsnWCdzS3Ess+XwW86ua0GfEPTwV2vOBv48Afkri41GZg
oESsKrID3o1iiNvBmXxF/qdA8hdokg7agnFyS8U2M9h0JjVVvM9GMFgxJOC4h72H
0UPUCqAOKCv8lHUauYwIxEoBnRxaFDTO8+OwtrHkLYTcWi4ny8Iyv3liDyfhCJvy
PCbYzkkBvlI2CJgQFP0zJ0yVMMACz1JOCd1glibu7/H+h1YlfBzc1lqI21YOuRjk
mzI3ZRKw0eWhPJerv/zVFpRzJMUWKVmRtoFp+SzgCvl8f2zOoaT+65w8Rb/s38Pw
m2fBE7nKjeN6xJ6QItmdpTXhh3ahHJXE9gMp2XlEVTLP4SA/TrfkHZQQAPWBnx6/
0kIKhplbef+Q1PpEvvGi9cpkWp5h5JhlEMazdaiffcXO4qhyo6C9tvPHCazGWSY8
8JWqe2ud0B16GNMpi81qHyUUD4bAHUf5wu0nYSe+llULVXyXCgwjYc9YH9g9rwKI
Bk9szM5entlf9a0MW7Rk9oLNkd7ti3wC0GACl/ArpQXOjJvg0LyC2nMA5eJjWwe8
uTv8hMH3zFwUFjrb2pdRVzI1YpJp943l+8EoyY8gmr1S6JdCjcylkhKoU8s8kWAu
E4U2qNYPfpJS/zrjUv/cF7B5Tb9ENurxMNHirAUjY4sGf+ykslR9VTndfstuaz8X
/hRAryz+4SkPb+1nBW2dDYJtRQPMdarsJe83QLdDuIJmBDU9g+RJeblGJHc5gH39
aHqBTIPO6WYFlxl5cHWUEyDPrrXhZ41NrZ5zEOXJdmx3wuExFRw/ixJF5Aq/u5z4
xCxL1j1DnR27JlKCfagASFF9G0OSRvcE8VHAz+wt1z6IQAvNlHLL6SjCG8sBs2I8
xK757x4SUt+c5PETkj6h7jG9oh4wlCSF8KdGs6GYOBhOIKaRiYCylWea0z9A2WSg
wstBeKdchw2FUWfTkHkm6+v3AE4xdEUBBoLdexes8mtestp00kyay5Igf+AFaYa8
js+uLR10znfS/YjreqX0gulA61o5yD4OK7ykC/FmBj0CWhEAN53LdLYK1xjDqxYa
SWZVbmV6YsfZ2FCn6Xfze3dU3I0NVZcmylY3DsF1geAt7KhN7saKv8P5Rx6DRQWA
iL8CZwKoZZ4NtdvdvtWqQEqoaZhSi5FISYJjrjt39ZCY7MMp1caS1xXBxpfRA1qP
dwdYCmZOjLE9QFWhd9yhOZcKXhYuSjzfTWopaJyDnB+9M5efyU9km5Xhx9m5rPlZ
xArZapjd+e/Iv0OGuDu0EdqRhQKBkLV0Cse2EwSE3c9kwrLhHrYTSDEK0G6uekRO
oSykVZWVCODHPBogGGl28LPFMIzwaDtShAHcAvxE37YFDoOHoAZdtWUaQ3ucgR35
7Ru67GhHjdoglrvW7cjc1zt7cGJqb8+EAafEUAD3AmE6K4wsttPZP8UDmslih1cv
SmZ/htsrAfesAwP9nj+cE5oT2+Qno+lAZ2UTqbNUWlD+KXqPnk73Cv8kpeI5wtkQ
4dXG1cYcJHA0cs+8IlgOJpyX3xq7uS2KhTag5M7AjTMfGy+x561YekXAZjJLfL/Q
zjksLeFFBzbAdQse3HN+J8UGzzgZJ2yXZz2iBMBJYxgCMEU4NGF9wJlPFagkRjJ2
EvcD2h5Z/GzizO41LY4i0gwB9D6YutVhUlSpsN2XkRuaaQGkueJkhhlRrSxB96op
ZcQMhFeUQpny1pAKoD3covlI6fsDE8XwYC4/iwGYVs14SehpzHQ/CTTfyrKGeVaK
m01rU/QW4V7pJX8X6Rg8W0aQ570651Op4AJRo/mvRoWcoiIBBeIVAmXel5X/AExk
sMSr3o9geWxQh6B+FSqv7xyp6RhG84tYjtt2L8RlbTANlFRuMaAh2efJdqfi50e5
Rw3GJMDMmN6b0lk9ZlM5RvfuTyrLfItAGFlr4Oy15ELPv2Wf/ZcvVhFIBVrP8jd8
KwiZQwCFfTQBxQZ2sSD6BmqUv+imoJLPjYwx4kaAeMlSyQduthNRlTKFewN2A8IU
R9Px94abqo+2AN4d8JuTpg4Ck/Tkkxaqj6TsQ6FfSRqmMtrDIhLeVOAJS9vBaf9W
jrWDpjQWgcXoMmHWU7YPI2X/CNBEt/lkUUNoTnBn/4XP4TSIWPRszMflc2rQfB9q
swYpNbJ0GC+BvKWrI+uF9E2CxfkPtAb6APr0NIM/8H2BQwVqKXHpVqVyzhguj9oJ
dPLIkfbpcK9OvxxZqSHYGVEOsSewGmnfNaD2XJOa2TMn3JHGP0TGEEH5W/RPXz9H
MEfQl7AiB9glLV18bv1rOZIopkyh+1XK9vfIrpTAZ9dGbvJ5Dlm8Kv2/MeUZJAaj
6THaGdcLFVMAeYek2SQlbQOfMBXF4y2N7nKyUPW5J7P9h2Q7SfqacN9LLRUh5Uc1
pbyhnDdKYunFQnRLOYx9Nmlp6IDCNfOrrny+Nm1BXrvgcThkckQIpC6kh8IYlfUB
MYg66NwOIU0pOWGDBuDCg1NlDMmyPwWOJ27vTpGEq08FBjgiqUCV+XlPkuMc0p2j
J/eDCmGpQV+FTwz/5u7IhYSfcuWt0ZSZIwVTlATcQ+FjmjY1hnNI+Pdc0R0kWTn+
H1LpNP/ueeN/KaxwMWgXl+RVDfuj0yOk2IfAxsjlleAGu7qvivej2zQ4o5U0ZUPK
08Bzk0i2xfXk7lMXjxYiGqtdbc9rN//Zcb7OEIdSClrU5cXsCd3MMgN+MV+/fLYZ
vfiIxvl4OWwecxhLkZDMxO6PAMFoNoNgxgLjYRps//KX8iGBdy01FjsbJk9/s+vT
ROfQ/LTFipvJpbQEA5aSLLuAPr7n0Ptz6Tmj+0aHMLsen68fwD77lqabPJz0hLZK
gWM8axG7PwpzOGcRv4SGUvrJdbF9KDDPWftkez5apknml0TzImI/jq1PmmDGjtFV
fHU1yHNkaSKiKwJVCdphU7s5cL35j/eGobdS9GYuCyK5lRMbRkNj1/Ql0I2P5Mi6
twfJquvgTVyhZt9DAvt7CCg+kQMiWj6/or3tzqoI6IJLgxWSUyEdiDeb/QU3GwXN
pXtz7o3BwUvLHdSLHKYBODbpi58bBWjAkOVeUhmTiKGd4RQI1N0w8kHbJSeHK8Hi
DdhvVM8qs98I0g5PTx/MYdtjZ/ifRPMztwgdbolH197lfhZFyvAdbevtMgemYg41
nvrzskVrGEp6gfOTnAvEpkxPScSbRWaft7FoiV31OI+ny2w4ZD0B2XaUm6q+tqnU
5IO5TkBdawezI/0/RrhK/NRg3KWDxjxDArU01v/5kQsFByDE3zC2jJQmn4i9Uy4o
AH2gZD6Sds6bSvdEaAzssZGq0mA3kmCMlfrcRPhq2+b2l5jkvIZERuVK4xtnpl3c
stLNd+faN646BQ+D76xwhreG6IW6B65f/vcOR9mnS7GxalNDCZQ0ek+72iKn37Xl
V9Xs7qtLHedgIdtjM9wNCaJrh/mxdc7D2n0ndUfnj/ANTt9QwIUN8aff156tgGgo
VJUxasBmFJ8+775emk+5yQLjglJuauDXpNRhxsd6ER2NZVFVbKs0uMciqfK8xaU2
aDT62fwJCF0Igh8esxm4nrtUZkrMionJbZ4etPymEiPot3vqHXjbLcEVC1+kr3IY
COTodqSX2fqDOTxB9eQAYdvH43BUwlKvtl+6tailRDekM/NQvQrf0Sj1aujQ0cWU
XDpL+y8/TOBKyYUae9BNyID4y0nPi9sebhEbdEn/fwLLoRy3iDHaxm26DRPVzuQ8
d2M5PNPwG29zuOOCttfXxKivhjp4a4gfNDDncLiroNSLtZvondTUq5yIEWIobJId
OR15JJRBb5aP5xPLhmSFDSUC2Ip2qQZJQ2UML8wD4obh7q1lxGhLHGbVfxeHsPJK
D1OpvObpzTiqy4M3Hyk4/jsYHr+YCMSZ97UkoPo2zGOa1AAyB3a9G9ziS8uf48DD
pxPhrPqWWobKshkgDi7A+4vyd0jnKH/pVt9vlfhHWyPFMO0yX3Mek7IGQHK/RzqB
lUneSsXvdVSpSzGCEJdS9o/icZrliITbUTd07Aux7Iw+dm+I/d1CfgS3wO+Dvkhj
fiGkmdp859FbqrPyGUEW2oDz13D4FIVMZQoP8yCw7Gn9/iq0Ye7vmHugNUfNOJ4+
XDiX2HzyHd9k/ifUEWpnvU+c5sl3jMzEviqc2US9oFWZz4kvL9GiHtVJtyd3qOP9
VC12+b+C2PCmC7qp7b6RiMr8/v/LugCLj7bdeqDXuBVC/CmVMv9oJGrhRFeXK8/N
4Lx0Vi+0/pZ3zmTRPWX1N3HSX0EXIjBbhZ+KR2LljyM5XXuVMkgNbbYl6NLut/R+
L5aHYjyx8ycW+NZYp6GcFW6ovWENtg793KUhsWX2FYS74lG3/jHFyhSwvz55SJUR
NoAVQLwWPOiXj7mwTfKKZ1iPnbBoqIMs61bXb4jGoeNxaH+IrjyaaMDERGL8iJpV
WXl2b+/rPKSK5mducaOZEe7digiNw4ZkM7Hk0N7Asn6QklFLynMwLnLdYHJBhnJq
xImBtCoDMtRVnfpo2G13pmbaw3tcO8ET4OYQo0wSiVvPoRovlU4m1ERcAuBkOnkp
SaGwpRDJNBqPGu0croOGdgSyGnAO1KEobsVc1nnHDG50Kh10vs2R1idkx8r1xi1l
SPqo0dDyf/U0qPh9js5+ufqSy/F8PAxzp623T/57wlmpiGK9Zxu2xshwE5Ku6pOn
/ak/vH1yNoZs/ilECsLIMQPtQxbQHwL6Q139ysxkpAOCDXHxzY/QUytD1ADnYEek
FApKxOc6xekKKVY3HTN1rdlOe/fdWagtoVLseBUX+A/XJIeLAIw+rMlz0AjAoW/8
MNVS/lF6lIq5ixNdF9BebGPKTIoDf5ATx0Xp022ykbInnpH82NPJhfn/XWaMonJf
nhvaUH+tzwpw2hetTYZ1cX3/N79d0lMz7iqu25l0ul+WWpAp3Zs5Y2uKgvnV2l0b
bHbmNztaUaSqSwOSq6lIjgroYsKiPfrLsYbpr/EG04cdOfhnAhafiy+DLTcfnyqB
RIHl1f23LXcMAy0t3W0zcvlSoJ7a0KwGu0XEwfrMVpALEOPuKHwOwEwZKyvzDIkq
TtNCohHPYpixX7ltYtRUbQBYFBHSf9hlmi5nvBr9ia9pk15WKAW7UzhOvT1KgKvC
EZQ5fKP+uOvQtu5UZ9gcw6FshfoKw22VSD3i3r8JRqR3WDQ9BNd0seGzSN/OqafT
OPHYNsnEC+UV1ZE7WJiSc/uNNNaRVboKT0b2x3LAZ4cUo0A580eE6r/60yJKFAcc
u5olM/xcmO6nOZzhQt5Ih/RkvUjYAmQL0t3CIcv9oI/jE95hOMI7TYT729Ce2cAa
ev1JMyRaFcfLzm0o9dkTGHsED0cJFo4uPmPckNI8sJ+jkcwMmf7CNwLDFySpJYF/
kEiSeie9pTspiZwyZqp7BIxfJ8BxLEqfTyPvHoN7QiQSeaRaHGffoRBuwdtBy0ts
X/naXcrWoFQTIlExboByoGWv4djpoc7wuxpE8mo0+uXYY3IEAtNU13gSR/6Tsvz9
HkAuiblDUQzIKqBpczx8k5XZhcrLAkabfMcv9+P2ZhwfwLn1LCRRrM5jSmDaGlJv
RPoUMDJ9fJtGPlcIwct5938QMT2x42kUsjP41+AtDEy+WLCQ0ERfsY1DZ3v4Y4ir
kjiXPq8lTc2lseDxdy70Q02IYAlnKbTAOFrkhlr0qq2CnIx1Z4J5bsllg2ocRZDX
uGcg1QEBYli08CkhS1A0eE6Q3mYS+nQcz9N88d5Vg2X93HL5wB7UuZT7VFHkzRCW
zAhfzNjHDQga1a9UQTywOaPbGDV1KhUUkQ1sN5j8EWI4Ju7hDCf941HM3ljEx20p
VsIx/9KRit34QWHXgy8MoLUtFPAeox72bX9BO9sfIn5nzBE3T36ligwVhw21SQ86
eZJVp/Vp9Nakqs0dZAVsLuZF/xS3lRXQ8IjfEo0kY2LmadVwZOiKCBDBAy4zepjM
77szgEx4h25dFOittOh12hJx6T9i+rCCDjFvlyhNinjUWA/nDwjBWUfQfAMzSWxK
Opjx3ZJD/Mdx/XuhIRRROC1ROF/PlLEO6ZyfxMxpcl/jWLsBNmQyeuoahxT+E3Dd
T1OT0Om3rU0ZizHQaYtr+yrwOtgwqnOojD2GzZCtWzc2wcay/41WrSFptwR/Y8sb
Y17TPyC14KqVOfGSqREt29vWOItaeY2AF90BHf2wIB+dHLer6EK8Vw5jPICgjBij
w0s4KJmha4Rid2PBgjc8YOYqBhdjD/H9CCLJEFguHQc2m+QM4BO0njXrPydx8+19
wLFL4Hjqd90Ms4fsqGGmUZRGmr8UDjLgdSYeK47aB4cwIFTUbv3v2jwMQgMxyuDk
EN9usMJWGnXX8UOmHhWVfdAJ7dQ+y2QFjSwf2n+g6Gj6gAFPHNJ7tL+7XMlU2EAU
ykE3cUg+APTYLZOVcb17cHQndJhApiwAgA/xWqeSr9q0gEuykh5EBSdnyoVT+bxX
PK9pVdb4O4DWWmRgT9ApXIjsfR0L9HBgAANwnTTDpJ/q4+G6EMtVoPp8pTjmwEL4
lsyZ3Ep2gl7PK3SBEoe0fFChs5WDdfdk1jpdKbUUrzA0HE6x4W7PSG5kRGz85/pj
2+hUoq+hXDQu7XHVIlns9nS5AS8IM6ic6xOrushEQURMERLXkpgu0/da+DYKHvin
F0ijbXD7lqqPe2PHBiBaXxVlnKwl+gLUFbgIzlpZwNXfuXq6HVz9jZCbWHQfObsn
+MiFgXjtc0AQXwYZLyUJ/G/2TmrCURq6pf810u9WTeoOviwgts8HX6ChPvrZq3hL
jM7jbiBcs7wd8maXRzWemrw/0AXVYZQCb5clIRyE77ouxx3J9IEueaVC/+7w8fYw
gRl3EPgKQubobnG6YQCgZdXkoZ66NAf3KcWJj0WMK07+PTZInhbjSq/+k/T7hl1M
NT8F8iFBC3yVrtQAWdd1FdQbu5rO5hiwE6SDWFN1nk0K83LeQKp4aYdsQGIAZ1lT
UCXHliIwfHNro4CCNY4e3Y7MNFEhvOcd2v8sNZVIr4L91qWT2T+FnfJ9bHXZm4IW
pMYYBvhEkYwU+RRtwfzlwhIXYdBaRaQs6hHWhd/i8R3Y/z63UCKXu87AqxdfQfd4
ejR24H8gWGJkZUgUGqhjwXRSnvFxRtjcym3wkl5N6uVbGTEH7pTZsxNnQxyf2tmm
+CdbAWNSWZTkRalBosYgno+bJIUvitYgS4mfGph+WPgVpoKk4PgaC3uDO83ND0ne
tr5+YsdFWfLRv+EFaGtTfI8mGCWiR50Bq4Eyd6O23i+XX2VXkyWjxZJ4fMcDI+/H
5aLIG6CVlwvxbNUWkRa9xOTHfYe1UdZZo8kGn6xPNQ6S2yXGGspvyN8cdBLo+2nc
XX4iPkI/kK1qUcgR5xVVgsmbINx+zjPmGe2xRytUCtUW6Il83iGpLhNkkA9d6YK4
G+zCDDJ2xPVESuy6oq/LKf9fcoO8rCLDeZTpbCHd9Wnsj4ICSEbHYNwql87rY6Wp
9q9ahIdoADzzcWCCqvBMEDDWT5piHqODjWnW8SN7v7z6rJIJg6wEZ0YnfSIA3m3/
g7A7MUoV3sCqkjWe7buL8hp6MByQt0+CGbdfDZIPCaHMFzL/j5prUP0dH/2AXtVp
hptJeekJ41X7TjQLvYXXGm8U7rXoMvR26LtkL0HI6hYfOOs6ublwacAD83ki0voG
lWOkO7yXDDMbGCn+RTmK0QdDYKbJi1wW5r52++7kA+yKFBdbSCPT+TB5FULMJnzX
JdjL2J6z5Vk0lXTOz7XYRtLoHYKIuOn3TYsK6VbHI1eluIu+3xWJkva4tWG3WHGp
XcIhRW/p76Htz7a3VDRh7F5EuC4n0CRdShUKCTmXfxGfCSIOF9DzwPQuAhy6y5hd
1iH1QsxIpbKvQ3+dC1AdWHGQGDSCDVdtblF18QVdcnk+7iVihBMBO3W7jP6MWAFh
AhNTnu/LWbUdGTxEwjSmP/xnan1IhtZsmQXtzwZTgEn1ZCfBF6HO83c688fz+wJo
o/hXfGQBopaYg70AvXZF9Wfpn/esgLyd+qNyjPZz51mDg4sCaWdZChwnLlbFoR8K
OU92APjvUvVdgoirJtChYEsZVExA9SkYzWDDIKmYk144cD994N0oSbiVNZHbWmco
3q55DsfoY9Y5X3P1tTejsIAvHianCYue/jW1COYdH/+kTU77a44QtCTnLtxVaxSr
GWuRR7rhbye+lN+Fm0MIYmrfLubdpp24OoKU46E7pEAkRKwK9XBW+ZZ1t0QCKvqT
8CWMn32yleqZ/YHtCbrlr73SZ6c26GmHsNurA8ysjMz+RHiyB+nDOrPrlQ1/XaM3
FCef6RUHV4axUBUoLr/tuk4BGIeoT/09cgGY0mf3XfpEkufk3GHAmhyX4d9jk+gD
WZC0eWxvB6/H/OEOQecwNJJYWfV35Nzv6lU/1aMwQmo7ACGnoWJXV2ppmC6UGZj6
+rkYd1QkKHctvKt3i9gaeScaxDbtuQl8DoTU8/4uteBrNLvSKCH8SErPbErqXOb/
tiYHg3qOoHd5nmyxMxpAy/3klP4iJO4LAAkYXy2GOIKOPKBbv5BKkxP/PWgje0Qw
12ltwvX6qOnJYNU6ksec3Bi32yupEvVLEM4RtSECnv7cwS8fGN4tIufVWcNATPwX
kodyH+fBDEWAopfErA7bWQuqCLdWZkIgeztxejB0jtBAezVaYpetJYZellkkkpnK
s1ZmQcmb0LyPOPQGBNXRj6VxNLFjji+ytV378Fm+V0EOs7vwm5zWw6KgJtNwSAfB
989oPrCY2TwaQxq0vC82f3zuocqikO2guWjUyD1SPaXkK8RWZwWwcMw3/tkOhg24
FnlY94Z4wW3S0bj3WXreaMEpZuHVodjk+Kthfj3c0wAXOqxOEgCp2UNH6FRh4AYz
PBXUcnUh4PWs4/1PUjZKSS9zTUqFLAfi9H3HsiJEDH2HINc5kyLqm6hNPA2h0uaX
O0VBz2D+dTJeLXmh4KTxqBVYnqOC012ilMVqjijuvHPtvJMZA9yXbdk/o95E8y6S
AHS12qycmHwXkLZNbMBm9VFQ3LsAvup1idpBKEklo01jK5/M2nVsKCcK4jWoPRw1
XUGjCm1XE3elTFXNccKqkPPv0+De91LM1/W9ySYFGAGfc2MfHuIjFeTFm02RYE+7
Z+/KdJdaunnnWxtnpt4itAov/Ik9E92PtLukPJSxmELbUhrIAMcXAzBcdWR+1BVK
wE/lMvFyde25E/dwrCEVWa6A2lJra9cRlgFjQY4fEyjKw4uYYXBeHYGtkK7zzk0X
CArqfBBOXqtt1wI5oLXsfdCPP2OoPXuQFyZL/aQHaCk6HZrdGnLTey+WxBlcWeXO
PnCYOpBinqSouCm/zsn50LBHd7mNUxSQ1jucfCYZkXsxNub/HXufa8zSVBDv0EtR
H1XT+Lh+eiJh4OV+1zb7tZD2ev9B25ZPFgOlUySqonkdir60Eke3jhaHquKhaIM6
kgcLBWqoNRuioHjo40YmiMRIsNM0IJS7aVeV9Y3GfGvPMR/GDBmeoWevS5JXo5qS
BlDz/xt8QCsJwvwf5KlsrUfK0TupMUoz3HLBytUlli0ipzdokrOuPaXr9176YVmz
TWzQvS8+BeRjLtVqmJqVFyAO2uUiGW5Mexwz0I6EHUQQ2zFC/kr6XjqMG0qyE60M
6QY8qWtPF3qXA8CB8WGRhuqmm+v/jKzhIIRZVHloTs4fVBYQe7ZeynAHRf+b/M/x
vny07Be6B/y2wC9GwwofIJgqBmUjIqpTA7K8w0EBoZDfuf/p+M7KDJN8AZA+sR+1
/ikFcM5s5Yh4bc+n0vP1PVJ8b3YhsPo0LaaKs3LF/r2FAuLWOCjkyTHILkRNkgbQ
Hchcu0vhnH8Uf1ELQDxOsyDTs9/V6E9DRw/+drssjSR0ky7BswyiagAFvOH7kupy
vG69cWyp7HY5U24HSXc6RLn4owA4cRHeIquPby5zQdoUoJ6sDvGF4/lLezjVZdPS
ZRSx44FuM0kHiM7O6ZzK8ifGcgTxfzmYFIDpliBDicURjxHVouLqrdYeO8TaCg5F
cC+GQqPnvQPJscytaunlywBsrB59R3n6udmm9+mvgLpEZn2cq5qgYJfZEJ+dmQ0r
LkA974uSg4KfagHZwgMsW8QxHCWwjUWK1nBi6/eKPrKShh1F0L+04zrzpBMKiQWg
gqv+QHIDEY2qJgpM0WvVRXPvuObtDbpz86mIdTx10Jef6Dpu8CBQyah4SUVoUEHN
CkrISXwZZkrd6z7Anp85yCJq7i31yAGEk/UWozbksQRcUO+yxI5gUQe3gppYQjqC
k7viizhHFZerntEJWLnvzyP9d7XW39BZieBSd2Vij4Ur4grXEH7WwokSSaaMobyz
al6fu6Z3cX5FjDys+J3bnMlLJGhS3hcCK3/wKknkfChfW5n4CPxM/AxGG6VRiqjU
R2iDODAr5+g4Mefa1Zk1hnnafGSu5hypP3ttv03cfr3MC1Rtc+Ax9JIDTC2hVYVH
vjA3S6+glCKBFtnARh55rz63mA82HXNtl3T90ztbw5XyeoL8pgfSxFLY3lrtDm21
KzxsuM1+ryA0HZ/kIhD3EyPjdAPe6jxnOCy7jVUk1Lv/bR6vynMJrfOfLkT+R0nA
1tHKKuzIUm+f+pfZErH+Gqvi+00vVxPSI5rYDNPCPjOPHdtlm6WbAeP4y4ecf6xe
0A07VthDcrHE8f8GXc5pJ7ggUZavzoyXO2ZDNMO+BIoxqQgflhM9HHp5fvxSEZpF
Ks0+uA1fh2ihfBZFlQixGp+z2u8hQkcILV/Ni6kNuyHh+wK4OrtSH2melvM3PIWn
E0JHIZAg30jiI3kI8A52T5T913CUOkrYxWHEimWRqpToXd0KUxvSS5yCxNWdUQtx
IQ20iBli1qMdF4lijfoPVfaRImDLP/ymgIpTTAmwfO1LzGeH0+14N8zVDwx7VHiC
NzkYulSOliczPHW/by/ldNSwv/MePpaVzD4eFbPrqN+lHw8xzgVFyHaDsVLgI/6y
xd7fzniAJMWpehmRYrM/+ECfnrufCPKYt2E0GCMISS+EhRZO4+xA0LpqvYCqUXvi
2W14f8GalM9x63sAgb+VVzadpmNBIrmDDjotkEcypYhAuZmv4XPc2u1gVoe92pHL
zOxn+/gzmZo7goJ3X1o/1fjLPBnYlOQ+I6N/22VApx+X6YC0W+wlQFCfTAlqIcCp
pfg6U42pgp/FllomoAxbiKsS2CXJ+pmZgGTEeo6pEIEvUtXTO4b0N1RZ4D4ALRTx
1Lazmbs1RmW6Q42we3DQk6W9KNDdtmjPBkuo+vYbo0Eu4Gg0HQ7La9xjDAe2lUDh
lDEnClQ7jL9V16fZXrtQ0u040Vc9IysFXJk7LkycU/lISn1ctkMhZCQgSuyeAO2s
opo33TQj3AfOefhGwquQR0+W4utfCAenj/aHaSUYfOLbx9XBPEtxEqT1ZyWrpqUO
rdYKaJJPJhQGwdFNHC0IVSXxK4Z5qVmOoEBsH2wjjV2C+6kg/+4bjDSjMotHzvNL
SX7Yde2PZrZlGVpyrmFVc1UnhLizvHCfRS3Au/la4XYuKQp6p3lCK2DspPPs2DQ3
mX6ogqTA+fHOwheigo/wPgqNoIlkoB4BEJgNTChOrj/Cd43WuGizi1Qxx3fOg9ow
Xg5eDk+34gWvy9/BEhJ804W8xcCX3136Hnga2S4/weABkkKOB7oUtBXMOQkHLCR9
t6GFPRseswc6s0RxhMMjEwk+9Ug1Xdi+zAru8BShDFUWvuVeOVZGHctgkJJXxY22
Pypf1JUDjAfZOhONxv1VYca0ycHenK/n0EHhR0LXHlJo9kUIQDKThbZIwm9oEjwY
gNZRll2ayOJ/05P1cpND/3B5D8+tuTdW3ospga2D051YncIi3AeXyl/r3ybqufXb
ERxZe2n3GkqIBYQSiDaWvP6iMB1GFs0OUtUVE7dPDWkZop+Avobf1f7Y3TITnGZh
luS4n+Odxez4/L0DRx/VPN5Z6bLhfgB8CT010dE4YhOTMOzUKo9m2zwrC2sFIs3t
+iJAxWBMPvT1xmJvT1U1bXbw1Cwpv7QjWFqvZ4QW4RFCP1wuyDLRuWTph7ua3Flf
50l43WxmP+1+3agZuhVnnrsyOOZtyZRPFO+iufxfAXqOhK7WE7/lhNgJFIxYo0Bh
ISj93TvYHhA9eNm4bYg8PVglhSomMg36S3e/RgW1286nrYr0YuLV34+nphKOCtF+
dHO7bNuHf2NDJF5KRx3vu9UbQktcsFSFuiBdAsX8GaeldMPsECB9t+yp2EaVnrOE
AC1GzGWkkUMi25UXSjJ3SbGcYgmesCwTjle1bKs0I2zqwphUx+4BfELm+MIwigun
cm5YZ69VRC0C9fDMWql3c0+EgQo3qstXrxpq0u9HprKnAO7k3OewX9samWNmuUYt
82kyGUYgjtxU5zj5LxRVbbJ0UDkyhqFhH5LLwuNQANEccz3dfH+y0CDzsCVA9z/c
X+9kOUPs5/0xLqX4bnJlyQOwgiURU+piXyxOEECR31S+pp+ldwhHWq5vqWssGiyb
o/PAfEwiW5HOLW59Sl0k1oKjQH5PWrPKtSQPGl5r2ekPrMR2vXmMuvgMJBKVJ7xO
Dru+Jq9B2KBjsVPxFlv7q9ZIwqh9ra0jythRM7ghCoHBwGiZox2ynhhKoolp1M9l
VVmt8Yy302OP/hiVK3QwQo/n4PKB2eyY3pOaSiIllcYqHdWtZEzGxyoGnH8wnELP
B3r0o3fXvnpuWB1pxqxnb/6T3cPh0t/R+k4yyeNXR/JRI/PgS93Nfese/oo5serd
sSeu9l+Q7adG4SAculCOB90NCQuJOQ6A/olmI3RxDIiCZcL2iauFQziyvOXHJKlS
bLuIFuTxGI8Q1VW+LDGcYtMMKpP9tdvqCuwZdDFvM2SNwVJlSBUBJufhkbidSlrS
ckym+kVQ+iSbXeYFK9ohr9vT5NuRS8K5mhthN2oetZQnk/DBOb2zp4bCyZOBgyWD
uL2LaniddyjV183ucHEJEzzIf3VIBFwL7/n7PhcXdyF2yHN0X3zO5oKieDOrNzHP
PPmtCvF0cn+CzJu1DsCOeTf1EQ0NzffwNvWDJ9XKDmKydSpNZN1oY9sVwi4lW55Q
U/6qeibwSadL5yofpax1zuB20eEDj6OBBhMM9mmVtVVvdk2yQzBGgoDKnLG6RRoF
DwwxeCnq4HmS8AU4VQzXXmkyO0M2VfseA9rytfmfC9HStQ6taRqH7CClkOp780mL
w78tVgFeUaNj2QU9noSwZPNzHms7UoRDQFJBY+/pa1hooCYMmGTy7ARa71i2j/QC
R+3sFcaOqTM0a/XWiu67IEKVwwh2yY78SXiaeelq9110s5QcC4D1SZJCLz5NoZjx
pmvGigUy2Y8dGt/1ft/DYW0eD4eAzYxSoBJEqYQGeMW9kSG3ccw6pZ5qv6/+YMxU
KcFIm09dPfYUsU+QbUAV6lPtuWf6uOSjSBx6Yk58oVxqsfv9re8jDYeIdA76Q0ye
0bUpFsOERfBR7O2ZOmdlV7LS6r2b+ykV8OAOU4cDdYRxjfZ04aKBheG03bsG57Rc
1bujBuN9e7LYOC30KMQ2zFRX0IBeKKzC7kQp4yZXesMnb35EfigmGaRNvOa1FHtm
sS9ffbLfwMSyxD/bTQ3INffj0sv2yAzUfs5Z94yqqFWXIGXRpFNnMP3vtxf1pfpb
+iktfVzvS9Q+T68OrFVbyPRz0XS0aFPWrkKaHuSYXrzSuNsLHG0rPeaoylO7c/JH
lduyxIhHA9E4LmmR8eh1bLfTSrc9onBLMrX84StyRl9+wQU90DaVG99ah0DNY7F8
5dJemow8EXFGUkvMvCi+1NrP8d36m6TsKorwXoLYgDu3VglYMpvpCZAoK9fXsmYy
7Si0LgR0UjNB8stcmRGmfzglrUQsKvXuXcpQQZEzSZXh6zMhxV+Q0d3Z0at2CR4X
7oAfWFONmmjaoBcwokDcJv4DUUFef+E/nDvK5eT/XRaD1wHg3tsAZ3WrXeCtfXW4
Pnwi3PPf4mTLLGm2qZoviTtuPencqfl5v2obgqa0faw4+eH20nazJMnbRwpi8TUu
3F9q39gCRz0JQ/D+l776LUxmHteeGqDj/RU6ZAwqcROIfmOCvnnZHSvyEKS6hsZL
Cxv6dOXHrKXlBs8Ygd2NcJSbl4NJ8kPyel3rYzpahSRhQ769SPtXG3ZHsgjZY1+C
RS5PJ984rj8cTpVVraXYWXhdXlX2I0fKil4O6h2quapStXPGPMj3EJSeo/dkukAS
hQ4+M9ZUcXATn40W0qGFLAxKKThLmafQQCXYFNBNGkPWK2kQszbcKHdbanWbiyWj
UAUB7fVt/yXVVHJnlTJEZ9Aja1XgLR/ju9Q6IOMuwZUsW6augsqXgYzRwQe2A6u7
F8tE6AfXuvAN60bGoh4HxxtMRl+5L30+Jo7U3+xKSLJ/bYi5HrTMMQA9iSBK3utP
zwFigHI7gbXU0eyPrVUTunr/srZnJzGbyvi8w1lyxw2H0FRYb5uFQdhCq/gN1puq
rR+Q8Gra52mB8evFCesgeF0+tzMBTFY5HIcv4VKhdaPWLfQgxYndZToa1fU8WNgu
VstYaK5MfDtOkDishGQ6OApyRNFdrv0PQ7e1G1RiWXPI7WfLc5t4gdnrHlGJc7vL
2b2URnwR+6vSUON2GcSuyXsVJ2RLD/PL0S+hUzblhxlUA29nxVfNfDtKigwujhlX
9Lfou1xbAYDmYO1nhCIhgQx/XXNmob+JdGJZoaifJPA+9tq3L1wXPzqL/tky7P+e
cOqBhCRxt6r94GiU6pv1IveWPRs67yIbrhFsIMWO2mBjKBc6VmyIswwo4Kbj05ot
I9/MD+SyCQSD9r9KOsjxYwfI+++V4U9aiqmYPSfWWnml/DsM1n5i6sGgnfAyZq9b
OXcvsbOkBXeePgX2/zZqBIX11WYaLUO1nmt+nXqpMzhrKYxKe2hrUnpK4DL39DoL
KPNgNwHNP9RCJjN59nUXTiEJdU1HV1/yS1AERCl8irCAxz1fpyoFJ1fdNBJlnwvp
8du70R5gV9vpQwnBPvyNbKxh51LEgX3uwayZCtnuJjD55k0i0xh1SiTpULxQmi/J
CX/o2MmUFo+YTmT1LsXfXeqQLBPAmBLN9drnIv+dObvTyJtRXuIMHWkXTcayOzLh
M7cRNfCUV2n2uKk8g2UHAFaanwjVMKIbLwXyuGQ9mp0+0G4Q69KOI3scrUUYHJOB
DB/CYIVOyZDOYeeDEY5Z+OvC8sFkbUUrYWh4o+aCtiRZ/jCBkE/BUlpYslbJGgp5
PINw7G7Wt6k56PvfcYKW+Q==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
ClsywOUfN5SMZtW5hpEMMK1+kF6OLELed3xUreqHjQJ5+zDfCRg+gv9RsWxn4iqu
OS7crnG27ZnFjHqS77wKSyN//w/VvEKjvNvU303BkGRvrEiRICKF7NoJ88uwfyp2
LZ3CUPKCOGrQZ/L0Mr83IY6nlo2xq1+dha1QoFP1YMw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 14209     )
IgtIIggwgFxqRS5Gt5ptVRWGxq5lZsZWTRHPspEgVoJg2vsi+qeau3aHSCJChvhB
OVTjb8/2r25hL7lfJHZUdvZ6I2o1EIlAflnEelgRxdq2xJhLSUgyZDnmMeK2GkHl
`pragma protect end_protected
