
`protected
Ca/R<JLdA9_T,<GXg?O/dFZOd)7>K9./c[-@Y\]4_-B5=N^dX5e&7)U7L/-^X5LQ
c(f+6HQL\#>gX+X1E.+S=E-9U-e8M.Yg&GOVYCA4G_d^NYEbSF53-[X(0^Q2I;^-
g^+/G>G(?D<K-4#OM52/SNV&\OX.+-C=?$
`endprotected
`include "svt_axi_defines.svi"
`protected
-cJ:>NXS^<()LPD]:\JQc#RM03=gDbTUG2ZXV((;7PXML\=4<H59()]WY8Q99bIc
?T(N8Y\0)^ZUC;?d0VPQ\@U7RfCIUg29^[O^&QX&HQ-cSI?U]>aDX/E/E9<XGI^+
<<N,:;:J+b>ZR7LSTXI4,=S)a)Sd6Q/MO()cI@a9_M@=\AMIMQg\Qe\eEIAGb@/9
MW,D]2b>/c<GdeRBS]f+U<5[WJMDd2fU\>J;=-@RY_bZ[LEI;Q<23SUaNSXO<(J0
A\>#&V.,9S6YY]aTY-_D]3>K?VS\Pbb7[YM)KM;>Jf>F\Y^4N3E#;L@^FD6ZB.f:
Mf5a^MF@_0b&_Pc7bU=>@DF#[@:T5SJ7B>L_6(FRJ:&65+A30X77P2=>-0TNa3=R
@S+Wf5@(U=V5G\EJ2ea#Y-6>e2Z^@c1PDRP^MXE#YG#I]Oa64cVHR-ZI<).g/F#6
=.=&7X6Vg-9S7:EJB^1adaU\?2=GPM]IMe,)XSI_@XS>Z4<)VXIKZV/##>(QfFHN
TYV4^.V)#51LIW2^/ZQSF6fHJgbS?M1RDd53I)d0EME\ca3;V4F6I-_:Y)V5bWR4
L&b86ade^3ROg0:RUI]dScV/QR.C)AZ5(g7O7THF:D?=8_N5J>#&:\3@J[^LVLe/
SAE]TAS>c/VQ&><b@aW\PE#H;T9GN4c)HDbSGcJ4AQe-Q&Y<-b)5aLD]H?8LR9Tf
0:d^HG=DXUE_F5]?;NW)K[FNN8f/1Z=8X4UX4Nf5X6N(9S(N00c<+>g9fLMdL;IR
Q]1-b+fF;W(Y-d]R0^#cK;P2TG_(2&b(fGJD(6/+#+@JH0c>YgE_.(SRXK4<5K0#
)=,V8JWdW&5#O9A+Cb2OfGaN3#bWAZR1>QaL@b_)d3YdL(dWOOZJA,1PP0GWHc_g
)>&,?&aQWc:@VOV1&e?-e:HVG&;U.Dc[=+H6FK^3EPXHd&^d(3Na\J\]35C&IH>c
=VA7#a3;104O:9\C20GYI?&Z4FdR]G@V6E0C9UX:\8&2W/OG?\_@:/Qd<=@RM\bb
MX;8^?<dHD&<?-P8IbZbaV9Q-N)V[>RQ?Q(6C(Ne6@5W(>I^O?cZ5QOJX.,3+&,F
IG?6F?8_G8MQf/=a1eJ:aOYV0SRM0LW.E=4fD-G1O(_NRG:)&2QH.\R)4bWPf7+1
3JFGW:F>#QHY_^]W?=T&I+7VVYdMLD88D1U#ZU#6\K]ZA1RXHKaX</0GTVGUCY,;
IX#UP_a\6Ib5?bg?[:dW?H&9GO/=SC+c<SR0b1CD/.d-A<BEF[Q?KXaO&6>@S9(D
BK+&2?^6P.&e2DcX=@S2;^;HP7F#M[21PJ^/9&_U#b84.(e8#N@O=1&L)?GaB)c<
[e3TU6g;-TIfKJB;2g,D@#aS.MATab-C+NRQMXcI6LgA^Fg]?ZX<5cTUEVJbHO7_
CgPF-EUG;\83G.f?X<O^?a69])JHfR>0f(^?d]E>1_4gQX[9bLa0=RS+DW:gSGPe
Q?QTPgXX6AJ:=S7MYL@51d/0HY/P>++5Ea(]S^E&gUNJE,OTaMU]3W&C<8[JB4(@
KKGf5MK.c5Xe[DAO1g]><cLNY)?S:HS0]&RI14=W8],>Z2[;>,Qb]KYN&?)07LcU
MVG9ZcB]U=56B,Qc&]Le)dE>C+dD89YV_F?Eb+=GQ971c55=9UY:ZUIVL5PSRC<K
5<+EbJe3QZ6EV5K,L6Cc-ZX4A43+RD@C@g5PgeaYOKg?UE#0e],eBHNfagXg.OQ8
?XX<SA,ZAAPQ76^MS@Q/\18,-467)R8A1RR;\9\DE]ID1.F4cZR<<(.EYX?^<&/B
L;H6E82c7IGNY;EC\cGN+EDU+fOJ_FSa2)2a<A70FCF5P#FRf6GR\7@e#3/Pa^,\
RgFATc5@GXaFU_[^WXDY]R2Fe5)#9ZU=b9]TAd()^G_^f+]Ya^^(C]aA[ZKg1DW]
NGP+FF[VEeT/P_,Y1VdZ(ZL#]R)_[<PMB,.\d/E13:31];SZ_1:S1(AR:,a:>^P(
I@FSJIZa&#JaGH0>=U(D5Vb;)_#>XSW.-#YD@4_OW;SXea)fHCV.Y2R<6-IR&RYJ
[VRWbUS;NZ6)5<fAa-UbUMIf8Y#EA3?@;IPX#:9HDBMPK4Nd0S?-K::cBe>Ic3<R
>@Mee/&f_E&K(H./POL?17O>R;,_RG#RNU5<A3R&R1[5#CQ3H_,W6(c:XK8_[(BO
AREAO]TPPPG,K4NT:HUJ=Aca[Y:cg>^8+eBHc84;RM@KY_\QDU^/)MX#OCf-^#WX
,#IGAS7Q<2)R;&TdX<>_Y+:_9,S^.N(CERZ#O:QRD1OT..c)OfS1TPO.G?RKg#=I
55OdfbO.1AP1AY<:fLT9&7#DPdPb&P+#87a&BS\YYW4#DSB&D;L\S4F([1XE<XIC
e:cR4G71JB3D9EKa3d&4>7R[>;\13J#eUV93-F..C8?MeH@INJ@0bC?5<BGDZB,.
TfePaeZ]\e&223Z-MND47EI\>4^^a-+\5e^R,^47VF:?5@3)U7(L&dHDMNVZYX6N
I[d\QaJC/0&S>0W5J/:JW@V64@6>J#cX&+CeY<4bSd\L^BO:RK1D&H8a4<#AdJIa
M3e@(+R5+LP\7#70_9Ab10@HDag+9bRC:Q3g7aXgNaJbZZ\J9R:Y=OG?9K[TeUQ>
:dTC)eG7/b9T5e6#>.a>I2]3#N([6U-HLWcV(G.E=//9GN<.?:#((:Z_b#W&84e(
(Qde,2.cVT7Y:5#H;?JQe-0Y03R=90FGV,bNFOIdYZ/Q8JEY3Te2S(a-FHZ:::27
&I/:=O&gO@SV4,K+A1+^?+HE=\>@BC0)CgY+H0Y]XLAFf8U21(>8UX4K;#52]f5\
O[<26?Q0RK)_><d/U<A?Qd7J\Vb#P9QCDC4X>Z:0E@TQ.6gA]Y>5#/=([X^A.Ma4
ZCN3Z,(57EeP:K-/&R#eHPa9[a-SYfJcHPT&8;=#&-G]1bf93UJY2-N/>#a&WYV9
G-)CBSc,dNUYMP4H6XegGC:.P600@:.VX8E)G=5U?Y-_ZR@Z&Z]gAD-cDQ,G?)O?
]Oa:XK3=Ycc?7X1bcE6,4OT=Y[/YK(\HYKU_XYBEgLB#5SJ0b4^bH>d#B=YE3)>;
@U,g]fD1f.OWWZ/YU/14J[-dPLMW2@0)^P1T/dBR:P8;@E)3NV&<3A(dNC.=b\-3
/PFP0UK[d>A6J4+W5OC81+<UDc4MSRfNWbJIP;SL99<,NWI6<\B]:7_GJ4N#>dSC
=8L:W4GOc#]1D-9K.7?,85\fB=;9,eBZ@e\)TTI\:b9ZXgcdL9,^Xc;S0YdQ2R,9
6]T9L:=N_]MQdU8BPK_OADAF&\4+]]#<#V@=e/,5E6#9PC?M\/,5:++f97(Be:C(
^[Q_O[>K3JW?X[->9Y<5-NWD.,T+,3).U7[@Q68gPG6;7QU-HTV?Y\SMeSdV@UUC
G9HD21:B;[b[@8d,4g/@Xe<Q/B/WQfeK]e(2fOC1&-?=U1g)72(NK=GLBT.L>)b+
,=^5QGE(]UKM5]WF:&K2A\2&/3/#K.P?@.?c^MS[T232KUe2)5&Bb55?F9RR/)/)
[^MA,BGE^UI-ZM;JS3S<.D4/U0DL\9ZD&5OJ7;[MeM<V_;[c=NFQcO>C<V0.X&J?
XSTXC5=S]K]E6a>(94D]UT3Y+@I4aPOH_KU&,J_Y@c4911Vg>eILR5WD0+:3;+&a
#-eHffDf(Ma\6JFUV;abbQ5)0de/V]5/[J&[^_@A(Ed22LC;)c4DZV0HN;2+).aP
KQ:2aF10^_-G[JV^FfWG_ZL,\EP+^gg[95CAFG5Wb8+I9=.P4)P,X4b-&dEe_C#,
@,73SED3<E,-?/2Z1dfP>+RH+EC5K2GT/DI(JD@GD5JN9G(UG3/6-]=D,e:TfLa8
a8Z=U6(98AR.G^2#XV#;NJ6?FeG?S^.1E).eQQ<K\]gUA):=&Y6IaUC.X@5X+,[+
15SK[X75Cf)fI)#ZD\)Y7SY#?8MbEd^RGPAVU&(5I<IVJ;8X^.-5IbS7:(H1>JEN
84M-aW@G\7CJ;3)W^5fdC78)V_?dM4c8I[DO+H,bWB@<L(5eWV_Dd<Q_7dU>;eb/
LC^&&Ic.JR(AP#3c+_fLWQ](6M[P8=QFeaR_85:)[&3d>^VR9A\fC.7Ng_f4g=+F
\5SXGQ0cCF@dIL^I1H/dV8OdM,&-DR5=fNc@\.<DBKTU3g,&0afNT^GLG+AQ7<8H
O0+c&M;?/Y[QAM2@ff_;6L.S)MYeL/9=EBa0I>>V<Y\0caMd[@D@@DCML9(Z.P_5
bG2M9W+@2NI>Yg=X9B@YND+N5YC<=EeG8BO>4fdaV2J-\-a(>3,2;PZK-<L(K1:)
O&C19eX45TY\:G^5NJ^Z\@69H]UNZSQ]2e8a[B<HFCg\g@Aa7>)VFLYeKGPZ8-+G
R+#Q.ST(e0.4JFNC^77Sb.>N(:.J2e>[gdP8Mg1Y#NJe<;Za\dW^W,XdNf2d]/_[
O#e]]B&-R>\)/6YH@A7H();LNf6aJTY=TdA:/TGB803\dO>MJDY39=/A2XVJT_9U
9N0HCNR5&J0.+^S=7fY[;Ng(K^PQ,B=Z)Kf1-GV0K+dO^4JdZ^[@F8<1(1M6LN\Q
)Y_+J)@8&agH1DHc4X/93TPZ/eU;-2E8)>^<D8=Ub7L);@:\gM,D;g(.>@WWg8<X
+Hb;H8Z5)>#FS@@c4]-CQI^?,-Q4)f8:HQfIK2D#OQ^Q#0G^\+)SBD8]T?+(N8XS
U0&X^-bO-Xa#Ia\/-?M;7A(^MT\d_QVPYT9C5Z/2MR7AaMPd-A\=WX:JB@F.NU92
A+8BBdN_N+).DX)R;@=QVO#[;X@5P\SMKg5?S,;MP:a62@_g;JNH&bUa3@I8W>;Q
GJ[8LI)-5YJQe>S2^0C&aEKX<MHFP>K1&E-MA\M1F--@F#?V6DWO[UCeM3+&?,E=
=2Na83@RCMT1HfWJ)M?OZfGPOLS,gF:8beS:,-]3X0H&EI.G9J<1-Sg#TCSd2,gc
]G_39O-1R,--3)+<1Se.FU)DHeJPE\fF@MF9EBR7QL1c5bD)>bNO&)#ZdOV77-f#
fD9IaX<X)VP?gJ5PJJe^2-^@UMJ8PU?[BR-2QdO0190(QK//3TLWEdLg](BVBd0Y
TcX;#MbSFMC3EE\Ke+c@Z@^S-f6EO<S)E-H3ZO,b?DH#2FH/1:&)1MLKP]<;,<\L
7[4F,],PA0IRN1/X,e0=-,O/QAOg7@Jb@+@V#9KB?-WeYB=c)S^IPA,&^cF2]FJC
10[MIb6a>;B#=DSD[XTP2X6[^@()ccR;,UQ.QI-ZbE5=L<g1cg(f\4TL-<L[c\J;
LV<O5(F35N5;LT_d1UG>[9(5EFH2C6bacK33b&Wd4@;/EXT,<]B(;8KEF+)(=6KC
-GJeb=MD7-A@fS2dJAMf@b2N^G_^J3RJ2T;-_/YKI[c>-)2V+.\QFED?V.-[@_-X
MJV41,O\Jb@eH&3Q+\Rd:@(<cBS1[)N<YM_(4@+=_-\C9dG_ONV9d\AB=6@]08c:
7KG0-LR#_,)&HP#;8^X-GYZ0AAJeK]>BK=QS&@F;0I0599R=d63BL_8c)FA0T(J]
^]H&H?PDbBB&\L2#b9#^E&Cc(+:EDN&#L?eF7=6e-4<CF@aN/S4?dIU,b)]^OZFY
g]ZWKT<6gI&VOa0W(JcDVdDdYUBT/R1@R38NW/XdD^L=8^_^TF<]>GgQ34g>SK90
/0f-2;/\CFA^EJF\Q0_4^;0^#-Nb#,cdWQ4SZN@VYf43NNga@0MI3D;XgHb8)#4=
N-^ba1K@HW@I<<fWINZU.5@A3aB.P^[1+OgO&C&LZF,?c]@-1QfcRZVNcdZeU1A0
5BKT@FCV#J_D)JM<J/\M_VM=U@66:8UQB[Zc\,XDF\&LM;JRV7ASMCeKe/5TL>Af
>FKG)3ML^KIDG^&VeYgS\=PQ4_==@9+ETNd2\1e7CEQJ&[([(Vf:L[Lf_M4<2C0-
M=C@GDHV4;Wbgd[QOS,=1IScJJMB[LYJ7=)LB_g40T\:)cGW\6/@TX9GI4QFRf[K
6+D_=^UD84gX;?[Iabd9?Y=3H99)I/BKeMA_N)9M70D9.ZaD.1PMTNeI^,Q:7LX\
.6S=/HCM-g,7=9@AL<J9=Y)a#K[(fV,.Q?;&\eSJUXCL.4>5d1&,Z<^SF-W,VR70
EK58V,b^:c.M#M_HZ2A/Z487:P11g,.9(\PDg>15<>306ZVR+a?Xe8=2?:ILXcaK
S/>5?G=?PBA:SBV0NeF(Q_&J,V8-WXYb>FA,4TS5L2E;K?99JSaB<S.3BcY(/)L+
1UF,NN^2?LN8X=A^WEQG5TU&R4F9:f,_5b[cE<GXA3Y4.2)?c9+UARKFAaYd8fIL
YbTK:8HOR7bY<7)0\4S,8)Ue[U^9EbA]>&&7YICIF&:+7LB8^;<;+geY<H5PCaX&
d_U69T2[^_D\[3;\JeZYP575;aX8gA9#++F4L&VYD1N@_.E_)(&aVM:/L/bL@b#P
c,GOJ_ANZZ:NHH1L7d^GPAKPA4#Q\3[G[[]:dV>9R=+UcY?&GO\>P_UBT:L1I)OJ
0_Y(HWWQ9_P,[QJW;(V2=?fN[cWQgKD94(K>^#L480V@YN]=?2aDc4H_AXOfTDYJ
256Pf@#c9V[MRFbLa3S_<J+D&@@[-f4>PXNPMb9U0II>OCO2O#@VM53)5E@,<;>X
JL^6WH4<IIf/DIcX#BIM4b?D[?_<3e?,P&>bCL_>;@/PR(=UeR:^-V9e\J4,HRAZ
X.>7E+X6#V=2d5#M;]W@)XC>M&/9bW)[(N1U+)2eM0-?RdG>&5a(;LS2g.@(UYY_
&bC5K88LJ=K=K&VMSgAT(DGbcCA7&V--)RQQQ9J43\00EK=]L^>LQ@X5(7J1QYSa
#F49cc9>#,Bg+&J776J->b_5IPC5>\(fc#dVT6F+ZH>X[Zc^&H&f8P<L7Z&ECV+1
:HPVAY\MIX4cObTRQX#EV3-WQ6^8+<7O?]>/aLQ9WP^+E;]S?R)Q2]OSC6\J#CG:
K(L5CCPDQ;Q:84YFY4RZ;NY@Z>YDQY>4^\)^4Zg9O4:>_);CZPEEM/W?O[I3B(+I
F<?C22-RgX[@9OXPRA#daYdU=aJFf]TU/SRIG0>@8CNFVb1>;6\6R.3&VD..f):1
5.OGWfd#1CNAGBC1XPbMg,;15G7-3Y)P#NC^:&.^7d/23IVb^2I?)F&F/5f-JIB?
UR[J_BMcGB<+_\W,<Y)-RG0N7V>X)6OYgd:36.fcf/+Pb\FCfdE+e6/08W2M59\?
+0<VRYA[HDX:I7bJ3<<>,:J:12D]?7=&N6SM?THS/(U/>S\RJSbL#Q3DL9FM+PZ2
T37aEc7:_6G^#GP,TV_,F+927L[JF9I<[0[V\IBQV2Wc2fC08ETU/Ud=,0ObMB2f
X)UIM2+/eR^gFI/Y:E/cW?EDHMaWABORM=09W970B.;\JB<C(K/^[OHEQ(GB,;DL
UQ.L2PND,1S9ABSHbc2L7W9e3]C^5(&4SC:aIbX)63L:bGO)6c39WK9+9\YfZ#d0
39cX5)f,Y2ER0NX7C#:+GQc_EYb7d3PI7\5?d6]JA2E4KS+Pa@\d3G+ZDY7Q\.01
CDRXP<>VedJRaf<GO=;[5.8#6-bHM+1<)])CK3a&.\.]HEa=WLf?BQ6NS2Fg.DTD
OXedF?224_<(:[4@,K:U3/PS+PfaN0fVfHM-LU/ES9),;L8MPBUdIY_M,EdCX[H&
8B<AX@UUNU05QdGS<R?^BVKGIW7X;Qa5F3DU&9EVADB(4^8VUdd=R-7JY,:,e,cJ
C-(c=#:HXOHf8:TY.@]^T9O],Ob3B\T=@,Z3G5248U\F&QO.>=a&H1O&LL-TaS/F
^g@b4Z?4)3V_L-(DWQ(,)b]JJBFa+?-,57.:8AS1V0SO6L,EOb@gXM8b2cPD#<P[
P-UG#;H-&)97#AU\T&J[XPUbS.^Y)WB7;VQ+DC5_1/?c]PPV94<6;KLbb//\UH?;
]O^.GL<:U:T:K63A=U,:,1]I6-Z@<0]B.e3XU8GXTb=+d>&]e]#_&a0JQ#a#a#1F
.>J-LTAcJZ?NfCT(2.JKO,(0FWP]ZWM27,=Y=6+UNS&_PO]^bE45\I)5IS2AUgO0
[[#Nb?<,64]2FHZ&/[W)MCbDRIW-08Qb+JV?Sdb3,=#4#AE#,]LQ3.,+BMW4=eD[
1He2=/#&,4@.@M9b,2\]O_B-fM&:2,=+R4.N84>2f[QEAFcNN6J?QdG[\/f=3P&T
=7--Y(#T#_GK1[dZ0-V)_+f?dK&NfYA.OSLA4RJfRPMG)P^g1;CHbQ2cT8S<CaAM
H9390bdFF<[MM/Dc6&_aICB<dHYPG,9;A#OHUC1-_AW5I-?[W?(O3^1G0CbCZHG8
SVEL61J_LceRKe=HBd7;OFUONN2L]MI[@^<T#3]D^A(KNT^LU3DY7F@8,Y1JQM?g
N;dQ]@Eb(T#e#B72ddJFP6&GS0?[cUE5CE\G:89)R9]_Y9#MX_S(^dI=[d1^/T&D
ca8JYDSQAT\0HB21\BN;G1^>\G.(2+:1/f8QWRgJZ19#e[;OUG8B7:?9RZ.UTIgP
ZGP)+J,/C9g0CK4b2#X=9VGY];]>6[E(09W]49UebK#aGS]:V+52<?<?@+[)1,UF
IX4d/aGW?bDE122,+\SUX+YELPI?E&7.Y)CcA29W\G]&KY@UPCe>[X0<8&3^0=-X
]H/01TXTd3YEW]Hg7^e-ZAb_KIe^9&&-c_#+cG?\P^W.,&?4KaZK<)UR[2EW5,&5
UfUZ9MVBFTH8PT&gX<EKMV]>-a-eYKMSMQS=_&#Tg#g7&=6&T>\f2(EG+Cd>cJIT
5g)6bU_1RTR1:+NRTK:FJHRKFC(OM,H(/\+RW=PFA4Q5?A@NEC>D^P23A/SHJa:@
8:/_,]L69/_TJV1gffDZPN\_6/&<I4_NV0f-fRHVZHBR6Q2CO[Q?be?2c3O8&R]F
cc+3eB^WSXd-P2V\.KHJb[9/(6GQYD3:d@+=7Md(O0F[0,R@.b,+c6,;Y4QQ52D0
O^5Se[e&#O(=RK1(d&GYb8D4c)QP^XRP0H8NJ94gEI\/?Aa\[3B.7>/SKH.0f)#N
KA&3R8<B@6@Q1KX1@W9DA&:H:FF07/LN5W4[aKIP_8/#g2K:C]e9T+^G;POWURe_
=/>2abJc+6Y>Y]W:bXd01ZLaT,2XdKYNfR/FU6WMI]7X]&B,a#9X#31\>[(#DIeX
.e+149S4,<Ub\fg)3U,e)Y)M:ef4Z:a[+8KI/5WRW?E70ZB;.74-c0X<PS.Y8,#X
,CW/21S_6=?-M-B;@F6>g7O.bW.70aJ5ce,NDS5X@--6?G1<GL909JG/#N?,bF]D
BA5fVbK#FaN,9Tb<O0\JH#_H&E[U)D2-<5?;#W=<Q^]Z,&GF<MD:.ZY73WM#YgX+
;D#UEV;&FGVgE/0Wb--(M(;TAJ)(U1CT(ZF>-5:48GHC]].eebIRK,EQW0-6aY7W
3D+R#TB)9Z[fHaNYd38P[H9:TO=-35\Tg?HS.d#A@59ITHVWCR\@2G&<D]c8/JW2
-<BA253LQbe\2B<#.ZXD1B#^DJRA(2&;a=IfY];Ua1b[(@K;3=-A.Y-_/XfPPNe;
95D,,<9d70R8Y-gUd@VN3E(&c)ff[O((2NPHfCPdXU(BH7GcN7)3P0ST/;+YSLTc
eSEbA:F5I4#7:^MJH=KO_eM/BV>a4@=CHXXA;HEd,Q<^HMeeG)>):0XPXfaLeZ?@
7VBQK+[#[(BS9&g6cAJQ2CVgCEW?Q3HAA]]=<N=RLK?CETW<:QXDXTD,8K45OQ-7
JaJ2YO))S(/17eO#[858BAL\c/U)6PaCA-[XI5=MdJL4BOdc]gcR1eBB>4.?@4=>
/?9^\Db^#&^8cGV3E/TSA]=B\MXC/-WcF:Ba6_DB9AOd>PE?cT2U@CJ<C=(Ie)PL
[CbS/9QP3=A1IR#+EgS5BYY2DXK-YA1bKY::+I^LQ;>?C1dI?7DHT)#5Q[;>1Kg]
1a,g^dR:U7]#9A/aR[[M+e(D^_@?,V5c&=:a0KD,#bZVH)P.YE)2F((7G4GXDW5/
>//7CA_0gbR:fG2?Z&#ZUT#d=Xe9L48b82;X<XXX4=.XM^f)7aA?M+cKC<VeL&8E
[FJ_EPGBacC2YW;<[63R+44_9Bd9_0KN/SKd-A,6^eL:/F),.?W^N]4WIVIGFNVL
5;eW;95Tb_Y=G#DKGH-;B([>2<##4aJM,Q93Q=[BKRb>G?DDd>S:F+L.)]FZ7a@-
0VM9\3;&d&Z(J18/R;9dN3=&@UG42cD4-]D4D.F.(7D;VHZW<=(0OV>NF_F0,@:7
Af[?75Q=)PWK8/@^d2)GP9=\bF+;\d480-NH+b5W+/Wf?V7=ROgV9D\d^@@gfRb+
<fBd\[[&NT[&>UNRI2a[_9CK6fR3PUab_Y(&d:_?VHAC)1[1^5g:9H24.0;TH<,c
HQbXe5AR:IHY13N9NW7gfg38V3K,N^V#&7P\_?(4K3b);CNH)g7(JC?<XX5>B?7T
4-4H.X6ee&/P9cHZ6YgPR2[.VF:AJ&<T4A(833-=77I8@#1FF.-Z/:0a+1-7&6U:
#E\=S2?9#<U9[@2FN#Q)7&cR75DPWEFP:4K@S_K?6-Z;OG?IK2,>BLX20EfMb&8<
G;U>:?HaP_4;aWd<FN(KH8#(8e<fFgU3[FD^9/DUW1N=,F:MR=EVZFIRcT9+HYBO
=56IOF.&,3]V&PN9R#;JJ4HQW_A5IBS7BA87EbgFYC1_NDI7g3^U6c^Y0]COccZI
V#J_]7Q;SW6C.XRAA;>/2,;Z).5B0=._cCW&-,5b48AeL@:DGR#UFPML=IYeg3^D
(XM>K6_cNQ-RBb52J2fP([;:CT;3#(+9,1F1eY987<,M)gf@8\4+3_3eeLFL0HUQ
9Jc3E\?f#3<>+N^81DAR@S+e+QV48PWb:>;OPC,-c7OY/3;1EC89=AM#DA4]X)[8
9.#>PXdN=P@L6I(_L;6e1K9;cLMe8VV3e_dMgQG>5[:#BAT);/HX7bEAIN10^d#@
TV2Qe5ZIeU_?O\4(?C)@/EeR^J\g#/?+fNfdPL43A[<_GQOVT.>JV/(6Eb-.V.SC
C;SFZ,(0Me2.5H,RD/>>0YccGI0CNPEg;(Z7_K@_WD;OHb\WP-O+OIU<C9C/8P7c
,JL#S<OLF-Ag9,[3D?M4(TH7UT?aTX@3OW)_/<e3:SfZ9fZ9EOQIf[TMW0&.]W)@
;b@f.f5CfJ29/>YPO/fP_c>,=9;=JMVLb8)[dDX7Ua0.^X(2JER068(Lc\\.]>H0
&DC;-&TU^XJ\.D4=&KMN3-fG:Bd[#Ae9_&GPNCE+S#44]AJIR1);#cgcb]\16^^S
a@5]I_U:YDFe0fg<bd-YP1GR[<V.1T5Z7?Jb5(Od_K@/II<I4X(e5CWW)c1KO#[J
g5,aS/K]ea]ALQD-D82Y[-ZT2LY2_/^Y+I=O9888C?CB3J-91B6)d1:25,J[A;62
]:ITPL[C5/-(:74(b77&fP3L5XFQ/?:OR):6P=QQZ9(2.CdKU8c;/O[Q@=U[]Q8&
9K7#QDVBg@eF?Y]]9VGR(;SN=/bT6<NWWG?)MZ9fL4+4CRV>X._RGTLL&UN93\&?
KC(K8GLUO?7Xg#Eg-HdK(G90T\EV8fTE,3#-0abL>WSLB?AYTYBE442>IU4VBYgO
4W5;=Q91R1Mec&OR)X)=PXDQG/KH:>@]Z45G7ZV0WB\g^=()g8CG0-QM,-T[C#OK
^=NSgYg=HaK+CIHggd:We4ATL>CJNF]#F1UT;1Yc&[Z3YIg=>7aYODN7&@G6@-;H
XG[&gZF&Eg+P159\.\cJG:R,X=LRXCRAKK0H]5KY8S_a2DaU9G[:=f&&-^+H3--D
K1ZAbWHbCfFNA:^B+_5OT=.HIE9BIaeeKVYR]a4K,B=DBe\86EQDeI^f5KcKWZ:1
#5UES-YCT9^WN1Y4JG8NRQ&6;fBK]L>QXTVSC:Y-I-\BO-@(JD15+^FK/F2e_QV7
Y)O>]:QfE:3(G6@S?0d9J++<cZZ^0+2/d(02edXO78Cd)O;7(-/g)[7If=+RN:cB
-Jdd:;?3;Xbcb1);>?MH7^+VD+J?d40DY\Df?KMX?.B^YJZTUGB[^6A-Q(^a2)@P
g4eF[46#/A<7+:JI-e\W?2QWGVEc);EfV[Ee69J,LHgY/=G5c-B[Ec[E3]0OYTg_
7:0+LHBX7gMJd&\R;V&g58LI,Qb2L?OI1\/WJAK^@EZ>9IEBdQ4E,N0Ld4fQ42e2
f[1/CeIe_27#+@@URQ-U?IOV1BR@M_A_Ve<@#>J.I(5c_U8PL;2MIZB260dbI^6M
?A(^NPP0(f5>6Wb@Ec<S;9SS,f(aLW5UGRf_GEeO=79<_aL#a&6UcGH<,IeAYNI.
\g<Nb.5([K)S:^J17W2gGE=1aB\&B1?YG?4@aC,^QRd+RG.-W:fPHA^0A29\3gQ+
KHU(46\c7f[\C5KAHIfF:@&>?:]9^O65b7S@:S,WJVK^AKA]bZKAe,@<;.?V?-T0
,9\C-;+Fg=>3]5N@g+A9/OXJB04@@YT]LXa@&G#5TBMP@EQYVBAHK6O6.2C\Wg6X
#N:WTU#e)PXX<C(7SBOd59O1;XZgd700EDK4cEA_;AP+JOH<_0<T;Z3Ea\^^.W<M
Kc<)f4gWOO\P^-4DAcW?B_,S#ReQ^D4-cK-C8()(+GfcZ^dCFaE++eZEGI=;TcDH
/&GY;WDa&<T[)S,d2IIF2/9=49AQWH.FJb^7LUaB9aC=_,_cedG7=ZVJFYVBBR_K
@.43@dX_?YIH\+C;>MfaU7fS-4QAJ3O^4:=>J)DVJ62MB-e#4bBWfM\>0aIGT^Lg
4MH549KUOg#[=NC1eT:-)>YG)&e9e,FdOBfdKe^cWK2L.92--#N78YfRZPG02HKZ
JB_dI@?NH7EYO40LO/8P9(a<RT,Z3ea7TWZPgWg=MF)3Yf:gOeHHI=-f4MM?#VK:
HD,&V35T,K6?23gY#H;E;IGdM4+P4.A]85C85J0G22b,N=EgL<A4,DMNU?gJ[S_4
dG,4_OVY9,?C8B4=L>-DE]Ua7NBVMa.+(B@>9SJH3^gX];:g=7=@6,)&<R>O0eE6
?MZKU5O>U=KLC:2;+NE^+)_S]&?Ze:BVWC;488]c+[M/SO2ZYL(Je:<8_b@3fW2d
<N6_E/Sg^/<bHM86B7L)C#EF8QS[3);+b&7eJKM];U/&/HY>]fQJMeX,gJZ9?f(E
1O\@5,BeUZAZR<I;^7]M69]?5IP[IPSP6_f/-,d33L)XaG:Y.ODC6_NHbMGF.CW#
>-N[5FR(3b(VcI7fM09AI0-L<;])A<2L6_3Y9faf?56+79;]Ag7>1O#.?HRZ^5->
AfB-QY<46&I=HJ^3Z+7S5Q^X,#_;Te#WadL,YdR,MIKY0(fD_<?=DI\+C+99:P34
&<[KWS?#8XXI>1A0:.U?CU#B\?J^eAH,ND5Gd2D_EX]0a4-P:^,1ZaQPg7ab]:L?
^g6+HD[b&SMC5^8^GX\7VSDG.FT:<4QeJ8]IV6FVc/I+e,@1A-^Z;[UEWd;S_Ig3
-0#KJ1.a5R/GWF])Y]I;KBSGDT\W]M2+\O9b=:5YV)&LgT8<50FC-A-3NfG]W46#
bK+d6<a[1:?+e;(HRWfEOe:\c>?XZZU8:KVV+dPPfGQ@@\:QO]PF0=(7\f<H9+L6
EA)_W-\g@QO-=dS7?dGgDUM5AP;^8<dfHDNS7<N&DfcF\6=Nd<VdO\]+g?.dfH_<
MLF+HDfeR).aa/URZBZN4XM57$
`endprotected

