
`ifndef GUARD_SVT_AXI_MASTER_TRANSACTION_SV
`define GUARD_SVT_AXI_MASTER_TRANSACTION_SV

`include "svt_axi_defines.svi"

typedef class svt_axi_port_configuration;

/**
    The master transaction class extends from the AXI transaction base class
    svt_axi_transaction. The master transaction class contains the constraints
    for master specific members in the base transaction class. At the end of
    each transaction, the master VIP component provides object of type
    svt_axi_master_transaction from its analysis ports, in active and passive
    mode.
 */
class svt_axi_master_transaction extends svt_axi_transaction; 

 /** @cond PRIVATE */

/** @endcond */

  `ifdef SVT_AXI_QVN_ENABLE

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use for each token request.
   * Each entry of this array will be used as QOS value for token requests made in chronological order
   * for first token request it will use qvn_qos_value_queue[0], for second request qvn_qos_value_queue[1]
   * and so on. Each QOS value is bounded within [0:\`SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   * NOTE: size of "qvn_qos_value_queue[]" array size is set to "(qvn_num_addr_token_request+1)" so that,
   * at least one QOS value is available when transaction is not configured to request any token and master
   * driver has to make a token request.
   */
  rand int qvn_qos_value_queue[];

  /**
   * @groupname qvn_parameters
   * QVN allows a master to change QOS value it has driven on the bus, while it is waiting for grant
   * from slave after requesting a token to send a transaction to an AXI channel. However, this change
   * has to be in an increasing order i.e. changed value should be higher than previous value.
   *
   * "qvn_num_qos_upgrade" specifies maximum how many QOS value upgrade master will perform while waiting
   * for a token request grant for sufficiently long time. This means, if master requests a token and it 
   * is granted soon then there may not be any QOS upgrade. If it is granted with some delay, then master
   * may perform few QOS upgrade. If token request is not granted for a very long time then master may
   * perform maximum number of QOS upgrade specified by "qvn_num_qos_upgrade". Once these many QOS upgrade
   * is made then onwards it will not change QOS value at all, even if token request is still waiting for
   * grant from its associated slave.
   *
   * SVT_AXI_MAX_QVN_NUM_QOS_UPGRADE can be used to customize usable QOS values. Default: [4'h0 : 4'hF]
   *
   */
  rand int qvn_num_qos_upgrade = 1;

  /**
   * @groupname qvn_parameters
   * Specifies QOS values that master will use to upgrade any value it has driven on QOS signal for
   * first token request. To clarify, when master sends first token request for current transaction,
   * it will drive QOS signal with qvn_qos_value_queue[0] value. If number of QOS upgrade specified in 
   * "qvn_num_qos_upgrade" is greater than 0 then it checks how long it has waited for token request grant.
   * If it waited for at least corresponding qos_upgrade_delay then master will upgrade its QOS value, 
   * already driven on the bus, to the first entry of qvn_qos_upgrade_value_queue[0]. 
   * If it so happens that master is still waiting for token request grant and it reaches next QOS upgrade
   * delay specified, then at that time it will use next entry i.e. qvn_qos_upgrade_value_queue[1] to upgrade
   * QOS again and this process will repeat until token request is granted by slave or number of QOS upgrade
   * is reached to qvn_num_qos_upgrade value, whichever is earlier.
   *
   * NOTE: Master doesn't support upgrading QOS for tokens requested in advance i.e. it upgrades QOS only
   * for first token request made for each transaction it sends to read or write address channel.
   * Each QOS value is bounded within [0:SVT_AXI_MAX_QVN_QOS_VALUE]
   *
   */
  rand int qvn_qos_upgrade_value_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how long a master should wait after sending a token request, before it can upgrade QOS value.
   * Example: When master sends token request, it will drive QOS signals with qvn_qos_value_queue[0] value.
   * If number of QOS upgrade specified in "qvn_num_qos_upgrade" is greater than 0 and it already waited for
   * number of clock cycles (i/f clock) specified in "qvn_qos_upgrade_delay_queue[0]" then in next clock cycle
   * master will upgrade QOS value taken from "qvn_qos_upgrade_value_queue[0]".
   * Similarly, if master is still waiting for token request to be granted by slave then it will use next
   * entry in "qvn_qos_upgrade_delay_queue[]" to decide when to perform next QOS upgrade and it will repeat 
   * the process until it has upgraded QOS for maximum number of times as specified in "qvn_num_qos_upgrade"
   * or token request is granted by slave, whichever is earlier.
   *
   * NOTE: size of "qvn_qos_upgrade_delay_queue[]" array should be equal to "qvn_num_qos_upgrade". 
   *       each "qvn_qos_upgrade_delay_queue[]" array entry value should be a non-zero positive number
   * SVT_AXI_MAX_QVN_QOS_UPGRADE_DELAY_RANGE allows these delay values to be easily customized.
   * Default: maximum allowed delay range is set as [2:32] clock cycles
   */
  rand int qvn_qos_upgrade_delay_queue[];

  /**
   * @groupname qvn_parameters
   * Specifies how many address channel tokens driver will request while sending this current transaction
   * to appropriate read or write axi channel. Even though QVN protocol requires one token to be requested
   * to send one transaction on address channel, Master can however create a transaction (xact) with more
   * tokens to be requested, in order to pipeline token request and reduce overhead of token grant delay.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       address token as transaction dependency i.e. if no token is available then it starts sending
   *       current transaction as soon as 1 token is granted while requesting rest of the specified tokens
   *       in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_ADDR_TOKEN_REQUEST define.
   * Default value is set to 16
   *
   */
  rand int qvn_num_addr_token_request = 1;

  /**
   * @groupname qvn_parameters
   * Specifies how many data channel tokens driver will request while sending write data of current transaction.
   * QVN protocol requires one token to be requested to send one beat of data on write data channel, so Master 
   * should set its value at least equal to burst_length. However more tokens can also be requested, in order to
   * pipeline token request and reduce overhead of token grant delay for furture transactions.
   * Master can also set this parameter to be Zero ("0") indicating that it already has enough token and
   * no need to request more.
   *
   * NOTE: Even though driver requests as many tokens as specified by this parameter, it will use only 1
   *       data token for payload dependency i.e. if no token is available then it starts transferring
   *       one data-beat as soon as 1 token is granted while requesting rest of the specified tokens in parallel. 
   *
   * Maximum allowed value can be customized through SVT_AXI_MAX_QVN_NUM_DATA_TOKEN_REQUEST define.
   * Default value is set to 544
   *
   */
  rand int qvn_num_data_token_request = 1;

  `endif


  `ifdef SVT_VMM_TECHNOLOGY
    `vmm_typename(svt_axi_master_transaction)
  `endif

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Random Index that chooses which particular start and end address entry from nonshareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned nonshareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from innershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned innershareable_addr_range_index ;
  /** Random Index that chooses which particular start and end address entry from outershareable address arrays
    * defined in port configuration must be used for randomizing "addr" - transaction address.
    */
  local rand int unsigned outershareable_addr_range_index ;

  /** Indicates which domain-address-range has been used to randomize or assign address for this transaction.
    * [0] => '1' represents address belongs to INNERSHAREABLE domain
    * [1] => '1' represents address belongs to OUTERSHAREABLE domain
    * [2] => '1' represents address belongs to NONSHAREABLE domain
    */
  local bit [2:0] addr_based_domain_mode = 0;

  `ifdef SVT_VMM_TECHNOLOGY
    local static vmm_log shared_log = new("svt_axi_master_transaction", "class" );
  `endif

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

  // **************************************************************************
  //       Valid Ranges Constraints
  // **************************************************************************

  /*
    Mainly covers the valid ranges with signals are not enabled for AXI4. Covers
    the state of options signals during AXI4 Lite
  */
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FzIOdusA0aFzKTeF03OJVsd/Jn/XHRPLRRiotDzrlTJKZDvQxQDFPTLyFLDdANCG
WGpm5ORv3ER6VlxL0O0Wn9vCdz6xU0Q4xz0ytrw8lUQqptl+7nNTfOYTdSCniy3j
/3y8jB9Bzp248vxp/InT8NyOGwz7VxdM3RZmp7yhLRI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 328       )
ojEftJ+36o5TWeSmBtpe19VIILobJ7l7AzNSk02y+s05RCDSr3EKH4nUovK4qc3a
Vbe5T9lIwDrUGAuqJAugymRKI7W0pZIPIXBfGo++bfz9AXvLyjwlh1JjYouXOxWb
AAxx0ZM/B63bTNrnSVsD/SOFndiA21GKP0N1XbMqxNQ0nqnIxdaX2sRu+MVJMoEA
7WyoKMenbgLV4qDIH/laj3+ORJyC2xrYjQyhCFLzyHdXyK5nkl6OAeNvUxK50OWJ
QFm52PWli3/IiJGlWC5G0IYb1mN6+pr6nzU7JatZL0DyiTdJSx/vA3l2v3We5Z1e
Kibejg/4cqd8yzLDDncvXQ1ddBOZZWEwWzl4gYfTb9ZR+c5TxxBHQpehxZUL848H
mgf7c9ZAK6q/DzQR9eIZ0VG/GwCmwa+CXdwS3j31iJ86RtUbvO9z0jMeNc5JTi1f
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
KXdESDs8V/GTsQ6qE6Q1TCJM/+7AbqqqxPMUpN9RUSlhvDI6bi7lYjFiY2IbpcUK
GLQWJ1OIFE5oNSCixTzg95/1kB2FOhnh1yTLJlIaucerIXs1IUdShtqOU06PERVV
ArHVUwr6q/UUTL9rO6y5riYEH4iBNDxmzFyxGkFax5U=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 63246     )
XIoK5ZrQ7f8UlDag03sHFA/MPkwW4t7zoWdtb7iRqwaqbmY7SCVkKD23zRX+g2Pn
DMvqL2WxXR0juPfmhlAsRc1ohxeehVU1zwhn+YkDRWEVrJ/PZjljiWPFJipk9r2W
jTcdXkJwSjUJCW9B17g2HoiYUQ70aRedOV/xpeT2Vwnica2beprLWq/hg9TkIMW/
w+Nv2+CmLwV2AnryP1fle79j8PzSXF/t903PlmRBCsFC2x++zelGzIZnMGXv/d+l
DBEF/Bn0UVKzk+Uhkb2RbHwjn6flhcMM1DF/eZRg7+hL0UYx82MeSt1ZOQcsur5S
tf1gtXkurSQEsDoAKBxGotGVkfZb8oAT3OYObmCScGYcWbfS+YgMKeZr6AZk5CCw
XJnvg3u0N056WgiA54MMWGtV5j+KaPJdfSfyZiq3P46FJkriSl6M5flzVQ+fTDKf
gQ8rsISFO/0M4BqvlRxgu3446jUBJbwhb62XQqXdvP6Hngy8kuyMjzgzN372lh/5
LZ1ibX5CDJT2vDzKk2muIMWJZzo0Jvzzs5c2n1wF59ITzNRUf1Z8OBCpHaJmvsX4
OZi3etrQc7HXzaQyVHx/s9+tf+sjYeBbvYe6A/cWZFHPKN//SPBsAIxX+0uNInpA
abAVJ6rVV5dux+78IIR9VbJ3xXHfSdRMA+HA3TdG7NHoh/7R+s0FaK56eTM7WwlI
rowsrQO8BaU6d/Wwhf1b9jxGiCKz4yGUMI5zTlnUJc7PPjKBZNaTIsqjG+M/fB0q
Vl0IsZIeYyWFTp+U26I8b24Vg8lgELDWJ6SsPY3ToRazesmtgnLtlfXeUxC7wTAX
QPGpz1eadsGaS//G9XN9eev/RyxMZAP8+Qzf7Z+CuR0N4VkPv8dOmWtRJFp0gT+H
f83lmyIU3aa9W6fUOW1sdv73M1/0wAkvRpQEbjyG8P2NC3Hdjql/iA7VR0Slt/ax
OOfzOyhq0WgeGi791NF8yn0ZDgmKrDMPSOroncbIbCSh8/Ssy6d6B1tr7bYNTu2c
TeeTLrKdsk6NudJgY2rDPiZ7J9NUFoxr/TPhMIdtqaYn+ayqSpgaRHwr/rpzbnzT
my2np+6umvB3bodLwubWlmCb5Ou3ZbywaqG8EEGad4vQzq+iuille4HQXdQYloX9
pHZN1HMYvnYFm4eOMRWyFA4+OvN7cwQXhtku+1pfxEdwxoihLFRhS6lpT0kFJnPU
EzHShILvSXIVqCCkNLbyfXraM0sPYhJmrXoB7AK40WbNULdcs698khoRxgCx3q8C
BOdjS4d8pvFG98o9B97GyGhjfFxQG0TzUKlBmUXFsbo9zKQohUNUEgSki1Ea3msi
JjmWqJeP9Zn3vd+Vq2JRE+5Oct4t9BJBeVrjlQtTIw/2fxdL8OnCamZuFPtJtXKo
E4Tz4vffhowri9H5XYuzo6XOiFFWiH18GgS8ns2LU8G2vMsBfr/6wIN+UXa7wOq5
FCLJQ2VLs/LD1USzIQ1y3TShFBJJCZU8VxFSP0vyPNmY/65V/4czkfbTPdOd4ZZ5
zE7zDqHERgf1vOCPGe4K9SNyrdJ/xtDBUoXqOzji+hE6fwAtsm2u103TS7C3q5Fi
V9J6CL7+mQb1b36ciPNScH9OT6euYEdnKveALBTOKdmPBEs8QaKtRyU8BEaHsQa8
g6Mpi8l3dx0yXdhOeO5m5rItGfzt3fWzn/33psc3vqYzl2SuqNrYa4ufiw8981ec
1gSXhJqYU2omqc87dAS8zTsEIpfqDqpzQAgFVplVTpwjF4HlUTKpdyl+8AcKw6Dy
vKHbz8M1vlo1jQNX0FYM7PUhYA9ASeRzVc+b/PBGUM7OFmfg817hCuNVsxC0Ui2v
BzzWUSS589Au18u57H/HQ56EwzJN/+ukUgj1B7tBlvCG7orYCTOjy0bGJ+TTys9A
2XkFyB8JjygpeC85lU6ED30UOLkSpP5GpxU718ZQX29zMVPpg9AOfszn9VezCcOl
zkBClo8AFLKBnnB8jw/RuKepCsTAorP9SgfqsVv2GDq1kDRKE9Tru79x5vVtxULI
DTy9l01i8LLvnyWnZVytA5KqaZUmTtUsfFUiVnMLrWC9Tigj5Nswt1muwo0PY0ca
kzs6bcqH/gBwlMFYBB6ojYBuOm2FVXPCnEkWgBGlArBnXdjBEMd/n+b9DS2phscQ
Lx8ZWleCYEpm8Gt5Jh2lYwxsNeFkQ18eMnfhiMgQmulOI/iJvBW3jU9U0V99HU1G
/6Jsg1Q/X2sXNGxfMQXtJIp/UIXJ6+4GcGleB3amouPh5+AQ3TpM3c5YGCSRHPF4
+AUjR1BOCRPGGjAg48eO+8B1T7RI7wVHv58CmP8e1aB2X3FFgQOzVzLtxnTDpPCk
G2e0rMMvw2z677rm95ndpEdN1Zm2XRPyoBwjcV+m9yNJs7qf/EUjZSGZZQMgEsOs
gKugMbuUqtPnn6gx53o6ps17+fAJZ2FPyqTVSuLTXQAoNLHOtt6MUQGBQScNdQ/d
aYRD/zrY5MqNOKgoegDIYzhBdptkQ/cKf+qLMyfEEoM+xQPBRxyY0mKVRwTc47/e
nh1sVvA5cfkZCcZxOX7RbXysFSa+29KEGXkzIFgX5FFBO2tAJJWx+VOX0o0N3qZR
RET5NrRDoNs2Mp4EX4XXugpp2XdMQ6NNMtWDfs7xwGN5tqBbyaDxKI8jf2gxPxFo
hdRYDnHg85avKQ37Y3lVXf/cfK2BZsw3fcXLfTEX3BBVIMirYg46ywLlgTx/vRmZ
tUEydBR3zj6qiGWGH1yp3DkLr0pbGjB4ehcz2mGUbgAlMb/T70bFLPjyOjbypJEW
KpTW2/UnDwkn1cUXH7IIY6Kfrlf0MWLz38kKPXN4Q8/HV2StIFfY4Tw3LXvpPKtr
lCBHY7t++W66ceJM2Eum1+i3n3JpcgXfenIodDALa6JB1nxx3S27E/aNc1S4cpBm
zVtO8Hfv5rPgbyjJ/34quupDy5H4PS+7Al2C9KPlz6cBi3OnxtSAknP714QgB6vt
CJK2WqoB0DduFUoWdg/x1c8CxC6sVsXBk+xgW0xR5L75y/IEuZGPHd4rsrSGkbuP
tUvXrDw8FSByUD61bHPQKSRXQMSPH063+eJj4hJcqtWktWVW8mtCrIMwN84PBnjA
UDR95v7XtOfR+LLPixtiS5Jk2Osy+M1hK9jbXyIQ78nP6Yzc3PeIxSQz3FrPw1ff
3HUctHzs3s2JP6nAHSfWOtojLERt0eN7M8QFH46Q91VLaOV+HJni1aowx1bExbe7
infTAwJKucyw5tnvypdqoR5mbIA8l00d1t1gwHvCRLknD0XYbtJWOSuBJOK3nLRS
3HxTNxxoV9W68aSNKF5GRzejmKOcLfxIFT8MH11riWSzlCS/15CmNEeT6zspGWCR
5csYay06lZaHaesZ5rNe9kPmrvI5+k5NqFP7jAXpNcHefUKHS7dj/KDOl0DRjOi9
wfbs8aOP4uOVNXp5CBsmIBX8yAqwvl+F/99mwiCN1iMsWNbroI2XODM4DGTvnUtG
r4tS2kU3AyRoWQcAPTd+982TA5UT0jIsI27JMvuFyyMahGs1VEg16r5tFOthp9SS
mepB1hMpvbro4FMBnichAlSJURyf93RYKZ2E1DpHsg3U97Yui+68Y8OTKx+gg5EF
a5pynzsTx9CvlOv9FR3vEOU08DSYDYT+SX+oJQs3Y332pFjDiKxan7XW7u9a4SIA
UCOPnk77L7IynPl/RR88j4EJB9tL0ROtRifHGbQlN++zZhQq59hLhqaiNLuKortf
iDaJ/SR+5GFl/VxtBCMsaQVz6wlHOeAK6BsPKAO/X1r5w9ao3XKoEP6pnj/uEUV6
6v5A1cvRKVmN4efkHw3qarvYKeoSTHbZyJntHJYwjrRxUA47NtGYXDCYoRgBQtFg
veQStQa5uSlQ/A/zmIRnAUbwnUd6UxD6L0sFsepmDdl7rx6p0+9GaqHbx5dDkB1A
zvmEmAFdmVwYt65Fk+HPa/W9FZ+1YbNonKdnQKmGUs1aSQdDzULaJJZQbkweDv3w
yJeI6hvinZcxG6QPU+fkXJhE/rQ0r4KHX+yhtTyJ6oOpU/lDn2QWOxBlfb6EwuSB
ofGSCDD2p9PSWAWChSH5LkVJNliy238NuzVMDyWEALKrbcPuTwFygzUXDvxcw6NQ
Pg5rDgUCueVTKJofwNvhbfHDxF/rl3XPkj7wv3qtp+2hn24vs6M6BKdar9Nl2vGo
LzKqZVsoRXqDr0seNeYz9VmKJkyFSFs7UaUVFzwb2HlpdDTUmVkMi2wtrcQpJOwH
w8ncOGe7F5j2uWaGKwoIe3LE83/EVCV5XZucvZBXbtgCgfi+VJVr8L694oFKv4lv
wLw3Dv1wBcbGETivCUEhdrKUNasvByuH73bwWU+GOWyZCyLtVmgshNVXQrHCLTZx
SnlFOeT79nvoxT7XVHl+PipXkfAt+eHANPk1e6YxnA0xNpTRlZ8zI3qwu19CpjCo
fdDK9Nq7dyqGj8kVZq9ho3+FGCeCvVIKnfW73bqTWR86tXh2im13shfatMXMaZG2
I1qwz8C2IHkBmgAeypGutrLCrpxiYGfFiq8FjMRpPFzUzixAmxdSYuh5QzCJRaCh
jhMyR6jFCUN82g5na3T2rESC9/VpvDNNIdYhTkkT++hV/8jImWbw0vSkdjtYh1f7
0gr5HQ54TxExm2dvgSC3bzRYqAQSGjGHSQDPbURah1N1+ew6c1hKFAl4FgbsSx9G
lsqptk/tRVBDjqwjFQmb9wrVHvle9+vsLdhRRWKOpmvHDtpl8Khy9jRk3Dy0C6O+
6aEuDAmvdjPTEJDc1PkH+YJU2MaaiGkiSMlXBvNLe1keUeMWvZkeGmy7vbvHSRgp
h+XeNi7MFryP3DkX0FyyLjLJd8AdULmuwHk8XpATxVtW/C9bWfeuxEW2diaag+Cv
A0DxTwpJ+tiq3rs2wTx3X3X8UQpv9jUVxTIPTcBaALQL414u93v9YJn7C4UW+qb2
kB60oTRx54iP/5zKxW9/fcp9jPs08vPpnGBoyXmofx/DROsDXZrRefkBJjQrPnYF
XVWJV1+xAhqoQL7G1fiGes71UE2FIFKsupFK2LRlJiUaEM2tvCcejeAVD53X6jaH
wCEHMR93Ac5P/NQJ3g9Xa5zGTtSl1A9kXLq1dK8XqSnRsGWopjp/xacAN3Jlgkb+
iWnZ7e69CIPMJmW3NgJgx36Hrzz+Iv4wEmd8IY9h4OpMWZ0LNJiwZ6WBY+aBNZsM
H4saSAtdknLWQ6iIHXzh1bs7CI2g/gbvRpdfifuGrpBTXA8CDgeNyg1Y/cz4vAaZ
UJH8aF0QwsBtEPiLCoOeTqO7Udw/Yh8gZ0jljiWHoPgpXAT1a7zldAmYFMRhlOLp
wspOBlz3hjwWzoXotLawkdjFVD+CU4zauthrHFMbp+w3dt0/s+M/mpoW0wHZVCwO
GIUCNayhBeV8RdvDEN2RnFiBKdxdsuG5qJk17qL+/G/0JkLr2Oumxbs1u/Hs2OTN
2csEexnCFXhcgYtr5rav12BvNkZafnWmGjYF8HoxFmslyqRzm3ewqKtNJrC2Gwi9
x09c/AhwLjRSBYaeQEQukzKFh54h3wDMeAkxp0W6c12fFN2i78cHJvlSWNG5VrZ7
51ujkXwQpKG8Iz/8jJaqkHcuu9lGd+FbcNJQFle9/k8mjPA6ilzwG98jsXB8OMjD
8cgbIPhmOJRR2Gj5kFL4hbIGqCD5Wqov9EyvOJDqWM4QzQqPcwDti5/kAOXRBe92
yJTdWHZph++nDKbW7GEI7bCDVBx855PLDmX13IWx0cQxcRc1GbnAj6VbuDQXSrzl
dtLQ+44M0P3gZsVFamXKX09oW0x0xbGxA9BznKt0K/aO5c04zQ8mYu1UyEwfhFXQ
/6MI6i05+gtO21Xd0HUfHV7OgltRK/2yrZk9+adkUmcSL0/rXbPaj+KuwOtorlFJ
79VSmq+YPNxa3oOtBsNDGvuq0+GOwxzkSR6yVP6wgMo+4ZP/lg+yBUYOFNOSma96
JzOJdI236fXQ9aq4snbseWxEzA0TPrx7WhQvTtP/2MUiXt6Z6M4XQqaYXynG0k+n
GQCvEOpqQ+zBlFXajwEDyDS3aIJwU3+Agcu0iBw1n5JQIusV+A5yVRyppJUZ5+DH
HJXkG0VyS7Ox9CJJa248mWJoBBPUK7HRghsFALmyMG93uQ2B0YuEMlYC4SH0wEMo
8zBa76w8rJucXiRzFJilbKe/hF0GLXYVtDQ6YfJus/zkyP/65D7cr1S8ixPtIlcP
cc1V3/2xVqfowP5W2cn+aDHJ6StTVqzqYT4Kl8N/cmdVA7DopMnpYpjCUhE4GBfB
nA8VWAKvbU787aRIp+qXWCt8/b68x8sn9wKIsjeG9Pkgs1v2msEkyGyYlnK8sxex
BBTQC5dDCdHz/e+CQf5gxOyYQbEQ0XP1NL2UK0YYTnC4Nunu2ZkkT/kE8ye8zKsX
OBdTUCm9xBY/z99lOv6PpLsgiyZZI2HlRW23fsjNt8AHMLd4hlwO1v4mMViRWlb0
cKURW1ePelBZn1lmh+13cRFUydAJm96o+5AeLzZ7nJrL3m3AGF4dt20d2VVgIlBy
W4iaOUqR/v3gPE9fwdJPdATc+vaTXr7MVz9ufcx/qKB1fW8E9JxVlak+GltckJAZ
PR8bVWLHIBpitsz+OfHLrKbwsoTHZv1LDPICnBgPrVQkjvKiW0hj0KBkw8fiTQiC
XN74gehCJYVnbXW9253jVQAWf2zzcx/FELOd3XgCtnRbDJvEzB5F0OS2ch2agzO9
8QFLMeeD23Y1y41ziNr0oTF5SCi5HWBrwf1/d3VctNLYT8ZgE0AXp7UTvWCH367E
AL6xCkZtTSA/ybg7W3YDMTiOWKKLNTCKUShTyIgT0rpA5fNzD56PBJhpfg2P+gFi
XV6lfWpX7F7YdipAvKoxU+3O9w3a+c7iE0uoaubbVUIJRmaggnfqyz/8hpbz9bYP
E0+wZwG5YSP7ArMyohOp4SZhjwD1ttLy8shGzhqAISPsRxYomnwpt5fRuP4/kHX/
L4kX08EfKLzh4jzffHwpvikRvZwNXYzDyCKnz7nVJq5QNOmFt0ON1zrsxb8j0Kg2
ChcpzW21hpt8Ft6MaEICo864o/jsFu9veVYjzBYbjL2HQAt9PXW7XqA3RW7c1P/L
VBgw4X4Umcem6UxIDi2xU9aZQEO4LQS6LRHwUuorZE6HwqqaBk9J4x9/6bZq6cUu
fPJAXprHYO47vdK92hxc/a+r1WUypIrT+oWFoZMLPeAHdcN4Lu4UiQaZbjvSQY0C
sW1golG06GQqR4Ahx3tcVpEZvBx7WdLUIsLT5SyO596s5eu2/mM3XKl3Fh02pzRd
1bxmp1pnHXl0udWhG036R8JSRugnWGd5EZVNyv+vJfxjfPJGBC9VpaMd+V/XATu8
/+ly7XPeZiFV3fEVs7LJAsZeu/PMHEfBvZWkGkKEine6OyOdpW/oMnR4La66Z626
/D036mZdgmsUXy1tX0nC9j6cEqVaSrbsN7XUTJDpZnyw2wy8uekR4F4nF58OR2SR
VZA7k6kZPDWhzcUJdE6CNCK316koeSA4SgTIKr0O54XJjrfCcFl3+dWI2mJquyVM
3/LhSBLs+h0blkgu0I9DGjQiBr6FR3zBoUczIryvHEjxY1YqO+uYK2z9rcfz7YLk
IZMMqmFuN8nLUEHHJkvuIwVw812mh1glj21s8ikWEh5KNOyYxzmzd4maij6VCMZE
od4p84TU/fsuDQ+RWrtDKqpyHndNbDmaP3oJZYGP4GfTCirALxi4t4qL8LQCa+ef
xPh0KjP4JmvTFGqzGQR7upcwNfnvETbeeohOXuQWTj80n14t7O/ZB1hT0/6h67lA
XeyPVykDU1vwHc8yhO2CiawLPie0Uj383qpikEWJGDxeH0W7bm9WOphuu561WIHP
vH/NnRnRp9Hr1tBlmE5fM3cbfbydh7KPgaeGeAW6H3A3w6AmYnPkjtauRVCFpJ2i
uq8ORbnwjyXXADlzYRrfI38qHnHPSYZqCCCZMRhmVyN2LxzuP7caHbOknlOxYDvy
Yo2xHLD/TIZkfVz5Bg3l9c+ZhaLcwbIV16hd9oxXrUBlZNMzfOOLO8UlPKREkiKL
AY7XAx6xgoqcUjJlfhaL1IVC9SRgZgQ+77Xk16A7NovxXKe9c2vuOmwMlI/YUmaJ
rvnebZb/+5oRS5pa5i9/xC9GQtaeVyaABigCmXbgeEdBwV23zzyldent1mqGlyRB
XWkjOZcnk4vkBQpUr4LUR6sa3GAwW5hA+Jw+1v01p8MtRCCf+DjJCLyYnSuUq3JT
IqOj+n2i+dLiK9kyYWbvETJ/4agEWS5mCbhFjknovuPFjAvzEBYwhof0XWELrOpL
EY/snrEbXyMLw6Cr1TCyVKx2yd1Z8d3sAyKAeewkYX+O6BetRsiamuIj3peyKWrU
yMbrJipemceK5Hb1UCrakK99ddjQRBT/eT9hrih3aUL3tSIx3/jcON93IsOkoh2r
b8FgPdbjdr+IuMYogpEijSgtadyKJIHmGV4iyPY0T+p7YDPPnAy16he2EMzbfAc2
gIipvE33PecCa8aqpi63bwdQmCQgfRTOq3TdZBKeSA84jjeleZH9JobNt/sAfFE5
zRtDS/550R1tvVydEepz6iPYeABr56YeczJsYyu6afnuP66mf9OeCg8WOAbtQE5p
RzmwA/gshhsJtGaHRmn0vIRRYvFqvRVwH0hpJty/TuYgSC26E3edDWy73Z5rphDi
YWxJS/yYCm6pRGn1qkRsmC4YqhAy/cFRBNJTs5lFPwhhY0It+zW4eoTomaTIqj3B
uwKaqLpWPwEb3LIE0tBKXMTRmVO9q9OvV5UIqiWCUDNBf83gRrZcIyNHjnaurGyG
GH+fO+1kjjTI6YfvChmK8D+OudKSvSsGlH/QE0YAk1sOr61jHBcfo0L/5Q4QZANb
e38xEsqEFvDlWea82oxL+DmUS79FQ+knCfiwHV35Z06cuaYmdmLqrhco+Zszry8o
rDjqhLgkPkJQrixCpJXoijuLALF3eHXixFrm8OgJvGUcOtOzMcLnl2PGfuXxbjap
RUPabyXUjDRgB9JLoPIJ7CdiWTARPkqV1k397Ed0tKeL+BxwUqDkRDWXsUNcEUk8
ZvapBe5yyRuxjaxFkKONLb2efA3oy652q/xGtRm7FGZcUFW+eZ4HZ5mvzOlfP+uy
QzPRUkB7b9kSfcAMrgqr1E5KbY5HwOLfgDptq3sdF464LDY2WXeMNECoyDSpuUV7
AkZ33kBoyCcbJbWCNlaO41m1KNHw7qSLGNEc3n1a14DO607ckEH7V54HSGr9v75d
qWV7uwYk/buw80OzWXFb9fjkV7+g9PX+XDu0pJ3b9tmES4XauppdrX2SDXo+qVZn
bx+w1BdpE2F/veiltXl99hLC6dmJCy8BTu4UbhUxeL3EczE7ieyR8yyn0pmX+OUC
vvhEJtUQJOkQIk0ShBU/+UZRq/NE5Mrn7doQTuN7AJc6tJERcOUhurFYRf9/+Sq4
9h+DvPmb0T26AnXEFXt9+GOIfjueAHZoLB2qvX9HIOV3X85YVj093gVqczTdvsnB
/jsKwEjmRFhoe1srI7teOQ5N3fF0mds78FTfeTcucVtpK8H9VfJbJ9wvhJ2K8qli
kcUJaGh3V/t6pOsY5bC0CRJY4lsjefYv0X0Hwj9x8nyJbYJXr4E9N2IWxTExRMKn
cTVT1s4fdUBeMUFmpQNm/6cN5ytxpg7BVBBFSPhii8qHr1Pm6Th2wi89RCKl4BHA
mZg9EXKvT+ykzcQKCoV8ZDRI+wWdOpQ7pzDaZE4UvbWcFlgUdYReLVMbQWs9kp63
wD1eIKB7E5Y1wSv9jfVt5Vr19NW0AS0sshsG4NcjjVl+AXRlazC0qejkijz8xZYz
Gif7VzC/Igfls/jY8RNAK9bQ2YNsCgs5l2NGM72SHDi7o2+nm0U/nagtG1c6FNVC
RvgHSYCC0BE/qjtSJPXNXaQko7BfsvdVPuXnyWyGzuqXEuAu1UsFQ2k25MhBjQ1/
1aiGij2+uEy2qPWOUysDJi4DwD2xOFeMKA3UI+rXS346W43AnO7cwLLiVtcivspo
5eAsYtePsDPirUvHp4n7zH2CBcNY0/+1xEbd/T2s4mJZQiah8GORVVa5TFNPWUjJ
4x1/H2x8vD7z1hXEERbZdIsEGqY+3Q3QQsF1Xr1cCGF75TpVkpQk+uWcmfk90vnL
88sYszKIEwlexA/MtXH+AI0Si7VcSoRwkLGM3fJ5YtBSsHBUwIiRx8N4mUpVdzt1
8iLuDbxbdAd1IaN2kf233wiwNeGXa9BUJX6sd0Jpy91zZbEolSPMiUe4XOMJkvdA
6VqgBlXzvetSzkNUSTBLoU7CMXQgWlRV8oK9ekPhXktFMTNOtBDbCQYO27NEE9Kj
Y6+kFhCJfKiB04NKQRXXYpa3OvyxvE1G+O5kPlVdGSbE0x3ByEcB5WrGjh9P8H9N
df9aNvNCyv4vHcXAC0BZ6mrA0NgBCeo3nCFGwUNJTk1DtrDK16oQmnDwkgdiqVbN
1UnQA+L5BQOYl9eHjXE+JsHbA/3S4xUR/hP1cOUeG3b/NJzsFJiCHYnh3xeEyb/h
AzjlJDYnKBlZPg2MEyjsx8t9cmX/jvocHzHkp0vCbbJjfKEJYQYhvtuZMNGmB46I
vP/7U2aLpjPB/sx20UaOGgAwzwZcjl3cxUZ/RP/xmLXhRerFO4hCLDpUdFE15cWw
naGfaruvJwduCSwteFWLK58iOuHL7QyVpURFkeqzBU8i5IfgMnySOihaztrrfrnM
g1yQ80aKfWKYSGAb6LrMnd17AUDa9lwnxmqCUXpzBovrY41GEIWkd0SY/iwgFzO5
2qmknbs7oHcEqaCwT+tOzMl34yazTfbB+67umB5FRoSBJF8eXrSrnu8MJuGUJ1v1
68OdSq3WnOYdgwJ+XuOlDfhUk2rHygbd2phrbSRPdOB9wL5f6u9p7xtUJyIbDdnY
kPdIisHpEbKpiknsJQdEj9IRqUY0RcFUw5hStEGO6xaRbCmKi0LpA/ZN6nUEFAQw
u52rHr7Wq1H4KNhqd+wEKx3sb86ipxGESWn0zzy81XhFY36PMGV9lcy3JrzlXxqO
eRES0cxfv0msEgy65+O9/jkdWBbfNJHsUtPVmkE9cKS630jkBJmz9v0/sNxgxk/F
WCUNAqUUCShJ87fcAoN70OU+XzA2bzKkXni3NluC96xRsECm+nV7QvIyed8RTOtw
SsS2tlZ8ILMTArVUwkcID9uAn01YubT/J8SnLV3n1BRVoKclJbSpY1MRztN/AMsh
VsMonBQN97RwpjErTSrFcedn87t0qSSzxeGJzU1edxtTquL64EE42P43l0A9PudK
Y+wqLPXC4p408OSkoG5WFzNi+NUROLkLZDd6Lc3mMhJd1IFcnB84UeZWYezespHV
zaOwmFY/PQAQpve3ow25GvIqsyhz2Oft6nbQm0CF14hLLNBv0+sLLxAJvK97XhAG
vf7Awx1ij2gp0cteroRq9LGisCGgEhkCXzh1Lwn1o7dhrckN9caqo3uPL5XcWafi
bdYY30LtSWaj0GFsGnSL/b6LvVFCIRPlduRWUheya+RhUZ8OYzPlv+Swfeibalyo
TPmpQ7rB0YigCl/MOfRrUGiqpRkF2+1k+htcrXhwI8h+p5EohDJt9kZnqHA4M/XF
u5+kXVQBVITEebpnoJ+akdKBqoG7F6nfKNPJ79c9ifbTP6C6s8Pi51KgdBAJCGum
Px2q1nPYFPxydPssx8wB9zNQaMdT3qc3WjOBOJojMki2/Lo/6C3VMtn43xbbYGqs
ZU5ulW3Tt9+N/11yLQyVyUBZ6wwXcUT8xV0RnQFhMyXqXO7Xnzztt/GF9bfkRPyE
d8WcG2tNJ9M4w8/tOUommQ62yFTTJMnzJbyKLl9w3LnJote5ncLZVCjNV+46iRqE
OMztRSbUuVA9sis4t/IUGqsIZNcP6DH3rZ7XLSgumlEOu9AL6FImaZORJIchSazH
fF4//8y3aqOj4dJ0UvEZxScWso/Eu5IenNHBG7kZ2pvm+zV+Mr3pGwx81+jD94Cf
GOz6QgaXO1kJWLdvly7FHDtwOJ3SUM+jJ8aMwcdUAUhp2eGH7BK255agFb/UEPe5
pt6/tqfQORFYOReeMoul3YijEUOtWc6ANC9dnFzvch2q6cBC2Fre3BY6OArdhnHK
9myyq8FQPcIxj5QS5i/urW/qxTIQbY1P5JODYxnV2PjWxA/LLqEuvAULhSJHKNdM
UkrdrjUbE78ZVV0TRQu86pPftqWwvvsEfb5+3a5usWYXR2m7gnXRt5ArTb6sVKHQ
NrqnBK7vjuU80HL5jnU0BVqh8IXe0LqoFx8pmQMJDhIi7KnRJgCBAB/6PKIQzUg9
7H5m4OizLEp/TgWNVx+u8iYCYNfBiaCpXor3yNbAPB5LioA+4O+US9rAq9JkLzr1
q5WYLc4koiJSyc2JNYtK1tCtQr7KJXnwyfZy23pfyVw94D4Us4Mklw4Z7MIN4xOw
IqOyXgbyleFYuC+81HPXWARP7QYzdOcRRBYfYtizeFQyEmuI/BGsCNjGnXIwvqbo
eovUJLW1Q2rozzjLfNBjuVubEARrIfqYr8Kh17MQ6V2KG14rNboKvL+RAwb0UP7k
h5QUUjVaTNcZZRUXIoiVdBOk9kW+QjYUmWpRTS1VskX2l36XvNG1xedP7rm6eigm
mDRFPKadJpojsOsGjyQNIjzJ5hu4zHoaErXC42q3JE2sRfxKHPD3pts4P8GkVWWO
PV2eHXefgwpz6VPoXiN/mHGA6on98IhPklsnTdy3HBL0uef//DH/7xVPCQ23NVi0
/hw9pTyDe2n+sBwpJgkDXEE0w7ZM9RzZ4jfXZ0IUS27n7mNYYrUB+JDwc75Dujb1
RgW7UOqBrK43wzXvaar+u9R50UtSy9r+4W4QbxJRsqD2eeNjPPcATzNfY2QRw802
mCsVtBGmUb3M49SdOJYxP8VjE74siMl8k83/dzBr8+G7uStLDBD4UH9wVGLcdLn5
8FR/rl/pug78DPfsMfII17+xQlNITBDB7jso5goSRABoGWgtcABkiIALvfmMLDFr
cGwlxFGF+MtvRkXdkHBjXlp+zbA/2bnX875joMktEbMfKXhJFGQPzKOV0cux9QYW
267BO5g0cB8YeeLdb7kbSe0qxpKwJKy8+rJhcG5STyO7FtOuWnR+xnltLYbduDqI
on1HUdqaQ5l20gxx5sJSZps7z3CpNn/QyLjSRqR1Ul9n0T5zan11suVE4EQl+lYi
siSBitPiTLHoLUPk45YXuX3xT0dGaNYsq2IyT8mwDv/wj5L4azJWgNay6tkjkD7m
iCG/z6rAo7CJ/peikW0IYmqO6Yi+dV5uljt8wxuk93ny8WFR8c/UJr3ya3ZMclWo
NPm+bLXB/4IkAZMsB4SqrzhAEodmjCAhnuO8UQjpfvJeXsBxnWXCTO7Il0JPF4pK
3X0tSvIkBardYOR/OOwoeYPGtww6d9qsuetXONrh25eUI6HJqxbsj1TtSLqFKGCI
yZqk17mmbfraaiGmD9FZhysd0gtOw+F8mejxbBCWs88Ny++IQKhcNZuBdgMjEbRR
GlXMb2LijVBvAEceHgHu+gWiOqAY4V20UAjBTDFgYec0SQafZB71tNdKIMDDreK6
l7zeG4dU2heUi82VvDt8hsYDkymgzwMTru7OZtlhutjXCXxZWuhuWG6k+x1LEIob
Aq3xQnYNOaUr5cB3nmtVX2alFGLdO7IaZhlMx7y9uwVOF7cAW2IjyFgSjzTBzyr6
/46mnBsKZf8OQV5ZDitiqLJwfX9ldFFNKHXBc6pOhLvlYZQ/pPbmZljJMet3rNh6
zxWUK76gu9XlTYKIXew1g1rcAWlLo1VO+JwpUJ/EZj+ZeTP/RQGif2zQP2niBR7D
j7IKYH5zo1M9PPJZV8dEWiHrDJNh+HD8BWzBDCuhsxfvYMBHHPQdh5OnWpy8GDYK
NFWFtcwMQYQ5GpqgZFJOtvcji/mwRfrY1eiJJFHQC6N6fvzIMwndcQuo4xMI3YMk
vu/eXFjPqoGgUsuoJY7tbyyzAkXmeWM2/v59xy6q06w8ly9cRU4i3p8H5oCuKLH1
iJHsu1+9Bmou/Cd720Xm6vd6umF7iKgqLOe3YZMHOXK3WkFuO82D9mMgT0fmYKFo
IAtT1e4/Wy+6mgpeybenhZW4lxeJ2OCnPOM6gNuPNXvJDF6RTmbHeq78x80Ut23A
cT0SoHXKqdCBsfvQMbpx9WRS5NhZsZ7fteVVs0UUzIEwOCcxlbk2WMEflLJBzpmy
PV3UqrbUM0yfXPM41fJ1dBH+Arjau+rDMSFEgcpTRhq558e8fZD1hc+XONMO3O32
5P+osCjrWW54GBQnAs0Ry3REsU1bCFhRSdM7hYVLsGIZjhZIbVOyth01Ir5XyuIg
aV4BP7HbkfhoEk7b+nWmLW49YvCDXpceOVtvDCBknIgs0wnwQsEaNMbN17mOTdKb
4up+U2cX9L0j+fnA2DT3YI01+3rQFDNlCfaZ11r9rzGs8dry9bqETCRCbklIFkFa
Y08Y0f3tyzqpk+oSJPN/fy3OfJ39wY2fwOCS7ybYGns4G/9vdqlIy4IjXuTGNk34
xffRR2W8uPIMgRxEYo0Ip6wNOCPm9u+/VQ7gYZtdqDAd37YoToumdH2pnC7X2qJK
HQOUXU87LoL9dtR0GuGeX15v3qCgPnX3KNnZ4YIvXcOggQfAh8DbNdhms1VFikwJ
MJxiY03VJncmtNECruIfl9Nl8MhcqdQUYm8dktzWdqWEXIAZvHGwRMHvF9VFKzgr
UkwxtxDLIeFKdzKQia7au52l4qmhQBIgtZFifP8jFyaTWA73wA4jXrdVWlMlm262
ZLygBKIJGO455au3Kv7mD7pul+emis3a7mQqc9/bOJH4FS5DfJUQtUT5cd3ELuoY
PnpZ7xl6D9JNWjmyP4EF068Ya39eeW1EqJJ1JAMJc96bbzaA5TU9MxR0PUu/BLRO
MyURrKvzTndTmjncP7+Q9vBW1Td9w1fEWdXqyjNzDkPdFQSHvWBOO3XgSXGW8ln4
8hpvmXVBqyf7D/N2LmolUz2C8nZOsV+BHtpD2oBzw+7g5hoJMaGL1OvFtYPTcHGW
TvI+LFTIb3bGfHlAVbyiFzZgxYCwW5jDifaDwBrIVY4xo8RyS6MJw87lVzTreq2D
Y3Yg5d/JqRDmU5D/7Loy1fNGIZG1E12yDdJh3g9pMTjCXwzMoquEikjViR4pgVHG
japv8XgWG2tYKBC0rUF90SktCZUvfJ5dOmpIe7mGdiVgexTAEd64FW4iCP10E5OE
6ZaQjfpr6p+MFmYrp64uVMLPHkZaFnL11CcGtiGgJVE0re0PCcp3x/M3jQ44wsbK
MdMf0DwOGj3ALIDeUnrNKOntYnoLrp/iF78dmsc45+kXFfdRXM4SkFIYwUf4x7Jt
ABYnTWoxou5hONDtIES352QuwtWa51mFeXoOBYqZvGPy6vb+qHcfETRRXDXf3JAR
yfb6+3glwhR7vippJky/B1zpW+qi3m6OcJ6hofYvOVAOU+JuBHuQz4XTorXoHYL7
OA3LM+LNzGS4/8QOJhjfx2RW1rxYH6s/eKEEIolSewtKXTi8PQSSXqPTf/mYu/I9
Celaqe+7Mzl2dqYdXoUaFJIT8g6j8jcRaiUYkNHUH4H2kLR3Rk0KvM+br3cwNn9f
19oofbAMon3L0+HDs1iDcm+jzwyAlpF6CSm2ZJvonPuixQzOR6U5O+IwWxr3TByR
kVMKp3irCADbbuaeA+CVfRgcGKV9YsSzWwdurMJ8fWVYvHhDhhmca9DNmh4HCY5U
FVDCX7xAJJJgLb/aHkpcH8VZVqE6YVS2QshJvbPTxUFVGWdThTX1E7LXoKY4yMHZ
66D2ZV2uc9EQErLYSefYwmX8nrL+6vTM9QdQPxT/x1cWDEzQiPnc26Pb4nLnJEI7
rzEB6RgkqSrBIlrqMTIwLt1+JsZabPkPasq4g63Jy3/SYeDEo015X0jvqs24lPZ/
OOEJf7XYmHQPit0fsQemk25hDoGVfpUT6flOo2H4rdoQyQcnPYQZYyWnJFwYUOJ+
hFgeJn9FGvei+mpsco9Vm0/YbPBOzvmwxJQKnT7QbQEvsfKIIfVxk618Mx+6Hq+m
jzdDKmUnQk5JDO2/1MwD81yCYgPKEtxOfCqFDUAyvVjXFI05ROqUXVK/1j2JYynZ
QHX8w0LoNoYSWeXvJbJ/yRkXXZeTEpeP8k01pm9xXdP8ZVu3g1lSPmt/i2E6epyg
zcE6+rCjgpCsrNokAso8rXx7heYUsL5LfRoSIefv55z9faZwdDF3eR58GaZYiqDF
9pQyt7KAuPOm658+qCtFMDYhpYpXd3twMOGwRbImqMR/0M4y0JAQXrjvUXcjMm1k
TY7oKcZ9r+74t6EwzZmRvgpA0VkKeu/X9dJiN/wL61tEh52RYo6XkYnPAzKkJ0iR
lanD5fGRhwepjc2W4rmszrbaM861SBMBx3b4P7fCKQMqbU1F2AFmh/YsiJRUV63a
6iz1W5+kRsnNL0yTCIByTBCOOh+YAD5I6k7vnprHwe3M45vWkGa0ziTKiTq8MWzU
zmtrteWqmWfgOMbCooRjVdw2b2g6EjhuS6CA/ibEUJqSQMqIuU36lJ4dTX1VCkW/
yCoqrT5KCYjqIadykyHq4+Ucy/yZtn2iijNw3OfR2MdjxISisoOHXjLxkmn5F6Fu
9yvz2VJODC8KSCmP1T0zGlqKUST+miXyefdfwvftVDlk3rdPWn8Oys7B0xtfdfg6
cMDPoyBmr5L8wuT5s45abSvAJSTkElnv2B9Z40UIbbgVmjwljkSAB210QYV0kfqe
UuhlD+K7PvsjjIg4xLx5EQLfLse7nUPmok7dKjft/Jq2cnH955xMHWeV7IKVzNMI
laAi0q7fwSGZZgK22YLiIJX5EkL4GNDn1JroJdFgjahPPWR01e+3J2ZUfTV6MAHi
EzbXAeRBIaSATDr7foaFWCwSF+mgvP2RUDpcjw+ymeQW0kFJiHmVEmMHDQCBU+kB
NLcYSBDwc1aF0KHGlDQ3r5SLsNVY2+m3e+vdkcTWfrewfguAkJw9ewo06xLKOcuD
kxyRxE8hsiQQZRVgtoCnNRRuqPi+MPXe7Nf2VvsdaY/2Su/No6vGVzUO389t1uYl
1S6qbrp21GJsOCQ3yTgOK3lFPEEBR8ZKmigwuvPk59y6tZDcO6PW4WPi9k7w3gre
Nyn4MPA7tmcTgWci2ziLRRSjGqzyktFWDWbn0ftM6sKRNubVQ+fMNTOJdM6o/KlD
glYjzPTGyBxLNM58IfcN7fN7EzCQTLA9TRIe585otqba9/xl6TG4OfTeit4l1EuX
ekfi8rzxYjxxHe9/fJnOYzLL+i4O18CLRDYrnm0MOOyk7ZdWfmm5MdJoCRCT9hIY
OAoeCv1ie5laLHGhVPYOVIT9yf9L+2tZqCL7cf8LcSdEm8CpTWoQjmXTa8TLN3yX
8Xk8WbvRVe8xpx3P4pTPKkfw1gTwwQ15oaG/Lk82umo6R3IX1nCbalmNlRKvFui5
6wt2CKP5oGUvpGVxODhHqHU9sVwv9xsGFA4V2y+YzFWNp6hcfSxOTD6LDkuMRtPO
b/KZMOxR3WOqS/PlGfXdf4pdmr4mLsVfsoUcv7Ez1wAEHu5Vq1wKnE3kpeMLJI8g
5E5iWfevmNWGpmG+P6Ngh9Y/r7W+0nhwvRarVwMtaE2eISQ/PkmBCA8ctWeczYAu
Tp6eJovL2M/XcBLkfdeGJzXWR0Tfs8k9NWNMJnOOUl1pB3RagrFIM+CcaZDf45mW
3q3Ey0PI5FZLBAsu9FypZXki8DX70AQcUaK6OEnO/Dv/9SdENKlAjkHqZdZNmE47
YdeH878cIt6LkVZpOHS+SI5tWUJoJ/Fs11gk9V6/ogyFO8X58bI9Se58uz+2eT8h
lE7WcYL5ntM2moXEXluL+TnIyO57VcCBjVaQ5ohZa0x75sj4pmL7gVIRL66j+zGD
YsuDUxrlJMNsuNZSMAyIk73TcG/qUCChIBhBHDrZ0e2mknt6HAsl3tlv/482bBQj
LCxtwAkb1aWx9pwW7esYc11V8C2Wo5+7P9KHDQxb2zUhFFWjzV9odZuAwgXTw3jc
0cZZ2pViORFgPvT51x4XBzkDurOOBmfDvi4Hp9INEQemPEdZ1S0hoj0EgFtO/Y/S
tlzvQmZDtl5mC86uoFK8yWcsR0CPobI5qjKTgRzXUkS7Hgv09Es5sSzFQVhL+ToY
y3iQxm6iEIYJQAOiBYmznN7PE7+HS6PKR07d4Rn9crUfAvu4Wft+1b/qJKTLkXBW
dxBJD7KiAZlMm4CWAp4kYO39ORvLizZGHMiYm9/yaJn2e98IODVqu8iMqrlXP2Cu
1o56HCSXyozvX4kzFC65Vu76zfg3N6BdeTOSHqCyWeugIw8IKEjWsQn3fb4slLNA
/rgVggD1yvVXN2yHg/ui8+QXjr1nZv9ube7kOEHMM+uR6P3c+vIgfgGCZRQkhB4J
k/yqfj3E3C1kAPtYoNPs7ifBcXvcwwXDU2IX709mmMsOd4UINvgJUpFkRl6dnAzC
1sZCs+ZXVy0I+Gk/SQEg4Mlb8JZEFSIkDnk8zBHGgnyq6LujX25hVdsOZSw4bSZp
5Cdkjqzy540T8X2kg880uyb4C+p44cyqoxdzkRkHWo2FQNii+pdTOzZ5lJOCPOHY
5eqCP0O1SvrZpPLISpj0ylxMpB2zhxTJ96hhe+XTXVmHu/flmUNv89srNV5VWMMU
nNsXk3Bhqh8dCEWNLr39SA5U/TH9mNvMY2Mg5CPCjA6ANx5oSwfc07ahQe2Y53wz
XIg1hUdI1mbmxreuzDSq/uPivrVdLcdadQf+nxICEMs1iR0Uca0aYrf0N1RoljhT
LNZbms0v76af5Byihsd2pOjbhi5Ty7vKE4dOUUFD6npCD+/YVF6dOM7rGFUkpRFp
mLmlehlq/L3YdBQckaRAircrO7NNJAlD3z1u/Q7Wt1Wk9ATUDVawGjcJ1FcULKOK
4AY+8tWXeJRyQahYtLrUrjQ+DDyYIRqOURD57lxXkOSBlU2TOQoyMOnDr5s1eANu
1whQ+8GWNXVajFRyB/c8PBKX9J8MELcAALpLbQu93ct5DeGeZgi6cE2JaoLxYfq1
7lhp9l+c+3IX2nM4FsZsU8zOejf8iM4ViTm7KQxzJ6NrZCn3wezPWq9kihnQaOJ4
gP4+Q5lWfyO69YoFQhHhtzC5RxX5Upgrn9ALt5XjqB2tfkQbBQlTEhxgqa/pgh75
aR6ShUlR5aP2nc6pGBVJaJLYAaAwgKqN/U0KUj7fGeesL/RrEVygA4mUtW24mtfp
iT2SCQxWX2O9aXW7tAcz9ojXBqqb7XTAnx9UDs0o7qoqPvj1gsYl//2Ohqcy8NdZ
GicSHUp/zw8+/o79roUyk61wS4xy40VTm2XPwoHUbyp7Gy/6n9UCQk2mHZ3fCDyR
EfcozQfGGC0tkCLb30MpcvG+R2eF8wHqbpc0tQ0t8JOzQDvb5QnTdJ9UiP5DnYnJ
kLcH7Je8RLwqaEqa4mhV8zmszGaUTyGsqt7ia3Qx+LPEUf/MG6sBDA/HABRzQQXo
WPjQ0PRedvEIqJZPSSvxKH02FQbi4WFV7jd066C1x4Jkx9tw8USAYmwbgObD99C9
ARRUbKP/kTHm1vvy5NSnwyv3CVHFuAlXG9VsDpxR2HIElDe6KPBEVoQa7+ht+hPZ
2ysPCY7R3v9fqaYbb19QJSc1n4Iz6XlXDGtx7d0/QccJDAZUux2DNVr/UZIp4pZG
ooe82zKTtWw+V7erg5bxFWjlTJtCiwYqgCc9kkp2+naXaiuWphmRi31LF6/wQnEq
6S5bilDhjcgqohF9pM397d8WuYU1lz7zNxuqAOVTS+7Oqzm8+Wx9qh8kK7BF6OP7
OrEhX+7xdCM33FsPfb6cPUau/dTjQK4wWvSRJbIgRmAl1DFnYv9AgmEMaV5QuvGc
iXGZPH0dsJJ1dOa5NkljOwn4y2IpXrFQtmLvPyXVuGJSOMG/MZ4JZm42f7XaJhOW
hLCuD2BTkB6oaOExlmGqJAml/GlAVV9FhJJP1Zu+Xx0yGonKO2S4A1Pm1ku9RKmI
cOka4384Hj72xfH5uO39smMje+Bs3v9ajsfASc5dwlJr6QqDBmuJaf9F0fuIMxAB
K7hfSNRbxcYiE48AeDhDOn+YVAyFaUK3EWlQK19OUrj4z/pEFhOnl9lfWpZC4qxT
OAJfo2UPlE/0n8HxWeUI2UJqT4H3mi3P/kCERi4kK1NdILUcjlrYUEw92h5VlfcL
o0sdvK86sCHdRC/17yHIJ5Phg01wCsY0gDiE4w/YPIt6cPQiktF/KuRq7BMTxrzB
kKXTaTSLFNpavEqQxOArVjDblwxRma8QvcVTZAEqai2D+OITOfNu+X6E5aChEXAe
AVX/eHGDK6OAuSCq4D75h9Q45x8hoZsv+/YyVMzvRhXx9BH1fQwpRfM+xn/FoQBv
hTa26lIRsB6Lls9KROVH3MyJSlPw9D/li+nLBP1nnDS1KBUT4WQnX+psRXZfBYzZ
d0icMx5dOzo4g1ZrWOKgurrUw69VXDNxt3bn4zfdVwgPucUSfW97kDXI2jBUj/RC
cw+scTnffPCU4BSnGTLNRqIf7PXADuD50qayH5aEAPC4VilqWJ9VLGYj9XIMQIbH
KPdmm2eNZes4V7T9326pvK6uF4wcu3N8coc8F64whCfweFWKNzUnfV66pIDf6v1X
RpKILgtYDYhZyAJDmwEIIXitzb2bqtKD/YrIyFoHmJEY9CIGBU9MTf2wOw78iuKj
sDDn4nuXipMbP5G/LKx+6VBeyjXuPW4cobY+pKrB6T2WDI40AzAaTO1wFFqBcDzU
ILYP2XRU123w7OpUFnc/84yIPZWZf1jfxgOkVhH07efWhm83meh2xrvurq/QUwIy
cS3N5zqCX6kSGp+6OFaLiKzRvrwlQkEyfwoyzrZMn+HAqnH9NjtW8wk8S04e2qtz
fVX9nYqBmgiYShwWdxC+aoJFN2AG5vDMZw+DRgm5JMp2HsjwbAI6w92URQmaenIp
MAzaZVEKQK6oiMK/45KVsqf1giiaxby2a752uKjXUt4gOh9p4hs871xkd9ftGXTJ
Z365di15KtH1hGUB4dzHqpDTUyPsd1xffwT4AlMeQpT4Ieum8yk93b72SdXnn5/J
ReuT52/3S8Drj/ttm74EaxWNRlIN+llA8G8PWk41gIkE28pQUTUwQDzDXZJq2GlI
L9/iwC2iai+Mc2aBa2sSPRJKaWf73Whf3Pn1yJ7cVAkp4FbM6jYEJpXg2EsnAmkV
7cGSVdsAyXZ+DNFcBdG0XUNuDSHSrBR+tOgiJ2shT/Ze0RZ8ZNlmL2Y5w89k9mkL
wPfcEEcRycQok97K0ATQIyfZ4gg4MX0vg1ZERMTCLKKhujM0D7tUSMm2YdPmKMoD
8edoReOIS15P0lFAPyC/unRSdzTPFRLWdLbe0VG9ET5o+pSXLHjn7obydNqJ2PU9
JiCuGd/usNF6oIIVDEKWKYiL+MjTA1sZEwculaNsikDOmo2lzspm7oAGWKIkqXy8
5YeHvW97iNExcIisviZHNsVxp2lZhv6rv7sIsuulJRPGthwkrb+9WNOKCOaohkXo
+zfVgxyJGeX7aaVYnPQGi4VTSKiN7U0wDklRyyjZaToADsyYHs/9B+H8K5NNTKPU
uIYGPd8AziVplALFd2VkHFI7sYMGDVbxCklDJZVxI/SGT89qWmmdZUSoSPEJEzPk
XixVm5ipjgD+3jBSeEn0OB+bwIoUtYcvcHpHIqbSnvqVko1oxGV6w5mv0dXknV3h
rfeE6M97Yhs+ZIi3eQ/LSh2jRa2mhISLzuLwIKpX07fmX8SUplWK9I3pF7QgZQlj
lL6AmGcmqDu25Efnxpx/Vq2Xi9Go6PiISAHHJAqDqmco47eMnJh/Uzx1PJwRwob5
R9scy9s4qXgcrN0cH2icGwRAfKNVphdNgh3V7RgLgIR+kl2r5ns1FRYh9zkrdf7q
Mdi7cZQ1XiwPPQaWMQ1pwjAEd/i5O/PqQ3yBbP0tDUGS4G9kWx1Vd8GKUCbrMnMF
hKVlkq8SUKtFHphbrS5NdSParLtvBP7qTXWiPCI462+gSedQLcVCOaB55o51DWjI
7TwY3Gt+mxD4yBPuUrUFs/rNN8clj9Si6IqvKDL7KkQRWdaF+smQZlAtzOhLHmIN
0w2fQF1qH6tH7ieOlrdEWdXj28KEDEXBswK78FXtdV5UaID2pT3OWa4wLl+WxVsM
ZqzAjr9JNwDZkbe3ZL3HAcpAww1/JU3dUzGcn8k2vyojOoia1tJ2sBws5THyK7rJ
6jSFLFt3KEtQ/aFSijUnGjvd0HM+35y8qR5SLmsrJxPJUXMETWrhLzR9aQx7fSae
9L0hO/7r1s/zsRzeW9+EQi3mTe7OWXtyZ/7Kk4UCKBRIio9Kw2cH+WdUh3j6d7wf
eb4gs39vugTGFcM9oIXzRsZfza0DTttfFgugBUVpBcsFDn6jvKYBcb1Z8WaHqF+q
Zl4H93gJPa6KG9f9u56xJWvQAJCBGJF2tdpEhItxHUlVZYxJ7NoEa/4rEeRdbO47
cVbyVNo+E1xeVHz04PoVNqbFIs92VSLygj7zniWAiI5yWZJfdj9H1JU9YJbQxwGi
oDRmSFqgzskIq1ylNhDwC4P6CNX+nBdyb+AcHe1spfrn/HgW9jI2QSQqyyHzP348
h0k1ccQviLVL7LcHE6wBsV9TMzW1cTOWld0uTSjJSCOYMEJ6X4Pd7SzID6HF5Ivq
z+HOJejj3NjN3ix+fS3WL84GLi4AlhSXURVUAnz4TpSILaJvB2igCywEen8mZuk1
kzDjaRr37Hq/Gs4a4gWHarVJm6eLkwckhbWMK60FRpbakAwjIAQ2jKLd0INezvRu
qwG28Shs+AwKv/OvcxQAd/VXr4UXiyNSG52Hqd0HikdX/pWYh3U7o8EOCbYJLd63
BQOUzb0Asig8uXb533hqVjxCkL+BWBixuc52lmIWXHck/qBs5OSMCGDnT2wQd73e
wN1lbOr6kMaI16u3buhn9tay5ALGyu9oIezypzPZtfnPCdw5gYVhZqn0Zvd57nf0
7qUNxxlMlOTIhJNe9PH+s1YVCHxtM48JKUhpjkT3kkMs+yxgKijUaG7sCOo0jQjh
sN3lEDVgMqy739xNzu9MeW4ApBCyFYyK8wHfM3azu1joA3C5qWO9y0W76b2vULvh
sHIKcyYiEd6+5Ppw95CHLagjv/23gB+4G0BQStzI+XNOCHVrCEXaxk+M51lokPFg
EqY8LMXOdi2DBAi3yZIRMvVlXaoXvJSaZ4afEORG4wtYkYbzVlXA8KFAnx6I5HeV
jBKqdcKWYZA8CRDiPgZq3vcEazvQM/Svlr6sU4MjTFYEZsTS4zrIJIYaKLuxO3SM
IVrd6eGX++NPXwNV1kFJ5oqugFBasDmbbzKC1rnodt6cie5IWuIa0WBey2L2K9+E
yzohrvjFwfDzLUrzhpp6qksvRsK4IeICXBGAVxeyB7U86mYWQJPK9jP0IagSETu5
A9MUKlCicHHWVDqklW0/vxthXZeAwXGJmGn7javpT+P/tqmFhxZGKl8UTYrHyYuG
2QAxarTdQ03vktG+nVJwfnSrTV2G5bJGPFQqJwnTEoTVz/BE438rQtCzH2Z7BnpJ
w/U5kzxca2+m+GjRxXC7ldTwL1ojVNEuDIZgd5aQgo/NdKrp4GjWygBGQqZIAxCK
hQxfdd9/iXfFeDw4kWn6tz3KvUyfQYlmqzWY8msjHsTa+ju9xcendP9EwoJWw2a8
u5uCAwBoFfdSQhr9IPAbDLyAL7iC7GAAIxeFOEsHsr3mOdrwnHs0QprOv3UmVn10
3ino+eM5DJLocZLHhU+ZLZrdTYBN7KS1V/VzB+Hh871TPVS6W76WhZqeBKlNwAbI
SQxkv+rQYjYzgYQek8pMc09IHW5NglLLsfAQ9l2X2tQqOJBLzTVx2gsrhh1JUHtD
d2PS1gnUUI5japPDcvZhZNBTanNA+36bLefAMwllOO7QqnPk5ukVaLQcao4KegmS
zftijEa5T16NlyQtGG1CLE9QXsUQ9QRHx6kJbXQs92MyLGa4t2RrCnJdmVydrFlE
o3Lhx014SKkYN3fKBGcwllKppvsIe+L6gZzYI1N7wPdixp+RIm8oaW6AbM/Yc4ir
ap4lnUyKgRhCId7DLjYSwQrfXJkueif0uHpUa3Yo0C7fCokU1GKmId5BnbSLCWyW
vWsomBIIFpSfVkUV0Hw7SPhKXmUzHfNJobBUGAg+opdnRkrEspHIXfhuuJ8xmciX
V8g1GF75rcjhMCOtF7F/PiqKnI9pW1dtZYZWN9rcCZsYgi9N8Yw3wjkwmw4ahViM
OkzEL3zQdNrX5BlHPVYtqhvpMbQ3FjH4NkmvKqYJ34NeU5D60j351f/x7C2KyfJd
H3eFsP8cEAlMKEA1c7DtAYyW6cHZrT0Czf+9n+Jo/Rw6ka7H3ryA0FWpscmwqdDX
kBe3ov4u1987mWbPIL6DlnlsrPVRtJGUC+RVak/ofiHFvbn6TaqpKc14INFnQAhA
wa4x9PVIBqXVOlO9Vj/Na1GVHXjE4pa/QJUxedSPlHCkGBKZU0kCWuAHzf4UE86Q
33TO2Amb5V7+Z2uYMe21HoJHjBaNh5IujR7ektbwEwjKycwUVroLKka09Fed8xbX
BJjhRWUAhoA7aLAJFWmtzDx9oMBPb0oRM9oKhK73j8whqz7rMnoAr8RNhadHN+qh
/MDAT2CpoNTzxtkR5dPzq+aoPgKC80KlB9/o3oxbwDURF00pVVNXA8vJmZBtrLPH
6JsK+u0TOqIdHGCDX6Voa4q70+kJMqZDRjAo6ps8wuxfUV1Ys3dh2+sOurbwn8nq
U0W1gUng4ttHKj16OfZc/WGhpeOvF4Y2eGeS5EAy2Ety8H60pJKtajSx1G4AHEL+
xik4eIhMUjKc3jJ4w07Y0rSzbGvWfnYEw60PRBM2klIW+9tsA9+v7rFaTKJ7eQmw
aNxtKv+a4OAmQt8pyaxKe+cQG8vAp65ocwTaTn+NHFiiRdvSBfJ39DOwBbezucna
4FhTrMxCm2bx+nwLaZ9lUEMq2/AggLMD+j0UwTHQGKzteByeZKmDlxL+ceTQTH0D
tHxGkfomhMl4NhhwX5Y86+CCsHlrOUS3mjJZhzDi9PijN+4caZUH0auFCjmyfo92
BInkMnBw+7YaNKaqBJjJ3UY7sL76wBMtivSzXifu7MBwo11I1jhTXQOZUMmmrGiT
p4nlaAGz/HwjTvCXJ79SIFkamQ6/G1XmxzsinWo9AUOVFmNWAOspE2BNyOwsAuQD
YraRjGHXapq39KhZpFKZjiqReMwA4swmtSL9wpld5i30sfAUcC30myW2koj23oEd
o6QUPr6DftHY/BgN+QZLl2JBtDOUbyCxpcPrpCbmA+b+lqGkUsGFQmAMiAdo74Eb
uSCJKVFVj6N9QBMM3sYXTSNQxewnL8LwxbB5DmtQOpE8R8hwAlrvlLvyuHRa0s0w
7+OBKk4zPwgUYyiNRwi9W8cAx0+1qZsVwcMu2JxhXoJLy+81DlQ+/YY7R8FXcjty
Nvkx63CCxQteWKUWA5Gx811xOsF3mCajtZNpBUI5sVoIRjPc6UeZL3mEeOB69pKP
GGxzFF7bmkfvpmVbz2IVZncBONZ20cRd+C4gDUZM0e+f/6A3oozjyI4c70HH0ll5
+nU29Gw4UTR/vIoGBjXlq89JRRuKBhTcvGqhigZgcIT7TiOrvC0oeXxp5YtNos5a
anL6mshwNSwRpSboD9sVWSIVowVNPnaS1oafuaxAX0JHVdMa1khgGg0NUxKXTbv5
urA0db3T985rPGfa0ZiVYH/dlAzDOc+IpFbn6S8Y/YrnbsFtRZak7xBR3CJBabDV
dmawtOIC0jnNkQtRFfgNM6Xpde2qFaNMFpAsApoXuuiLQorGiNwNTOFq2PEqQa2G
CUCKj13otUVoXCMumnHQxDNZ8IFMfAh9uEEqhFIRvgQuBj7wBrbTLiQaiyranCKZ
q6cjBcKbu9ECnnojwHVNLeb4DcVHKCxHCyBflb5bhpZwZvne4DIrUsAY+RSaF3wM
7tfT3mUO8YxTx5UlXoGGfvGx45HRPzeZjj/TMh8hqMv9cDIxtOh2T+QBva2VXd23
d5g+W+NczZXtPPC8IbS8Jg0uI95q7iFChqkwm2em5S0cx4zCDi66iZyCqnN5Zo2Z
b9kNVCtDoLS3tgG5bricz4fScDCwq4WmawRA1jPI7GPzMgOcA3DN/AOspC6GDw00
23eslxkgNTqdiDWTLgn0ON9D2LxTH35/l6VuVlszdJtAhtfPak3UH4qwVjN9ezY3
944NvD+UjiOVq9D+bJg7PcNiznzuAGoA6TgFOifVy1oSIgHXLRjDsAmgjhfqCQ51
8XEq8fUcVtoJudYQq/SUzcndjiSTCfkwUJwBHyz78sApnV2JLj7pq01XK6B3zmdq
jrXfWSJPugiBdKBPE4cXmmv506yjeus3Ok2c4U/jOT9+tfyoIPTAIMuSrYfslgLU
nMQums1hZ/m9Bsj+rY16e5A7MY548VHlayU5an0BDKTDRrkZfzf8rzV3nQ/cBLYb
0kgBl8/1exFiAI5fJrNmREL2OMGN5gYdaUVdBlvjMDuAO0SdXnEkUJlzYYx372gt
g4CL8nprHlTZMSG97fA/fZVhxT0tgXjYntqAMh8eqQej6k4y+g4LMMXbV6w8I9Ha
t7HAwYbRHKRmnXw5PXCTpTR7DHHoQl+X4JDGj6teIipo4ZCeQKhybf7ZuUTSnVdT
p/6qnp8E1p5hUrws6D+UCQG7zTR/WnoLwuoSS3Aw9p4H8ZC9oTQebtAQ6R+mr206
F1UmmIePSkt6O+TxQd6DkUXkomu0vNQKCM6KgbwcvqkWntuz4MgMScZhRaNcLab1
b3Bf5FajXQOWzbHbru4w9LY5yZF4WBT5uSgwtOf/Hps1r0Vx7luYO0po4L4gU1Vl
ibn2WnOPaLfgWagyyFcZVS7RJnBffPhy33ubAjO15Kztsm3YoXStVZ7xHbWoE0Lm
LTWRNHJu0CsZp+URgjscYvTcV5DoOMMdZvVxSXahXFSZs9Mu/+3DUFSenwxRGoJn
15lYcKjDuVR7K7BbCEG/4LCg5kBON1ASWK6Jzn6WaT/zh8JVWWFGEAFis5Q6I4/M
SPg0IDeo9cV7fQRDkXJ2tk4RJABoaPFG3CyQAAk8qYGmIgHlz05tz5mXjmd57X8Q
aAtq1051cCFt/hPJj6sb5Z9Lbma+y/TiIO5/m+HxhT0vfQU8nkJyKSriHsbsyCEh
ZhWvhWnv03nKqlZPIviGt3b6lRWNcDiokSYKqmtL9AInqiuyE56SLffuNOdld9FQ
3p5St7a5BCUlbEX3gPaFwFH77kSo2Tqg+TJtaTK8y6T+l6wVH+8ChI9h4bpUZ21I
iz2uLuXGNB+Tz8nHB1tWx+KqhxElMu7i/fD4I66kTDRE9Y0nAM16xmhfq9QG7wVB
2wAv0UKqKcp6njRkJoXHWnuZLA0eCdcCuir0T796Xy999fqew9Eo5vCDI417KRPk
xtgiBoawU+hlrFZuQb6VHaQOOUqMtZyUdEvqusv5StTKv3Dscleoz+5oD9FhUCBw
1lV5QzoKCWCnncapWsgr34RsIuU5fu6t6QY/P4zkYaWCT7auko4zsyM/7fy7UVup
A6mAZObMDZjNnSvAPwLVAA/SrE1a6FvQlP/eTo1R06fVGoXLr9Xg/1GYvewB84vm
4cuUliqGdV03t53KJMe3k6U2uS02awB3owWVuSjxjwzlTTFD3I9eaFOvwzJ3hg43
ERXm2TaYeSjve+heC1Bzc524eeMVj+EiztTgRReg1pEXSai4K/CKbcbrAVoBB8r3
Ul7hUYOqTByNCBdkUuUt0N+gQQm8IWf4DImLynvS9irEcOT6cxgZHDbeIX020Qko
cLMR0IRBYrvdMPJZZbJYNUi33VRyHKAZVEzjkyLUrVCbB+D4Rkkm4D88OYWuw3S9
GoWQjAIFOqF5avqiYYkjhGf3u7yCJicPiGDl9xcgX4BCxZJYzgBHTqFiTP2T4vSP
9oATQW4bRF7zXVqQ6UQ4YteNnG8JneBpQM7B7/Xwo1nM1wo3psvae0jFQ8tgW8ig
b67JsEmTnleGJhWTD8NxqfPEe/sOrZDT1Ye0qkzwMExZ7Vkx7fqmC+hOpuA297EG
qXoasHog1B4GFuMXkM07yEwWh7tQgjd1WCM1ZwltHFzu/19E3snLE7uBiaJ22q9d
zJxZk6GywhNxbsRBXxDcv13mlGHxbKyDUNvpAfKyoGeuPCiWB8bRwmu1czmzIDMp
3Q566W8TSOWEeBYCTGoHXlGS8LPmeQf7d16HfNvc6TezSn259207A6fk5usX94TR
2lTZczUwIKUjaiewuQekLKg46UJkrImVxW40K4RW27OESbkg6aH6p0q839lC8w4q
Ve+1y4IA7EM7xauIlzCF0QSjL9wvvZxMsw2zBFrteQYRzWqWgzLMOCsf6WE8ORhT
JFWw0e6Crf7dGRovMNJhoFr/ijN91vV4Vp47H1SRLPm0gMNzyQdI9hS/4bH0yOcT
+53SWpnUgCs8f7A7MVyX5JhS64o8pnub9ryIrdCt2IqUvaOVQl9b/5Kkv3xIymFy
mUaxdLhkeCZY/SZA0NiEf+P8fpL/HsZG5Ic+vE80uO35nz4bqyF7LcrrIdPUKymu
sgfFrcVdIwCJhk3w7XECb4KqrtjGJKHcTUGXKsYd+gKPdsaIYH0xmVXP6TQSqGEy
rJsOnsTPJzBw0tbkNxCY3OFNhWFR/2UcpOSHjGtuOgH7FfVGbfh6RF8OtBhZ8U+7
Fd5ikzftW6x3KEdU2O7FXMDT90HSPGhoWERKpFh7nGsbjQZIVAtomh132awRelde
ZZPG2jpfCmTvTinas3cOo+hYkJanHZ7+7AKtbZdDUAnSG9cJZExi040vGVdEsInb
LyFR7O400giGXfYYl4zKsyOVoE1LyHz07+5hQY6SqpLE7ZNmwFdy+zybO0kfB/DO
oAQP2ABQRJGapEd02CNpMjZidoMaiq6HDljtifQ5B4S0RKHZEcCxdnqE9Gk1ygqf
kg94Sda7sWXATH3ZIrY/Sy92ne1njCIzI+x7Zg1Ey/wLOzAMixDAyFpVaakLWTPZ
8QAAfF+sX1I4P4se5JjwDDKU/h19sHOO29y7MJ8rtPiSshQ+R10iIQjTSJQVMIEm
qJUkZlgneB09lnMBGA/VYm6qJompsiPmnV0nnQ0i3WnG5xc6S0qU6hX6I0wKevGq
jMJd88stKRunTHpHsU3hbBHhvSYu8TMW+veSXmCm2Lhb+RaTAd19NtiR5SGGNzvs
mjnS6CpaxF7YCTfLtdyl1t3OoRqL4x9qBKPDQ8ngG6xcpQu0YLnStaidIfxLRf49
rDsQPDB7mEkMNGiPwBPuX5ABzplWiNzACgwR4HVsVnL7I1oEC9Jift3WA8STAgbI
VDBMlCJZcUUtA4GC4B/H3ZzMS72gUy1iY8Wq3LGnoi4EJdgf4UDcZR8vfnt2BGAD
zV8MbB+ODFY/hNYa3huqqTiAMF4bUmdhruxWEu3aSQzHfv6Xl8KZSHk57m1n77JK
c/N7hdCoovkmI7Ge15eyv+XeGhq1lKmLEG9LK3aoFfAon+c62YliNS92T3J1Iaja
Qr3yd4BiyZboMuNmV5kPd7kVw6z07S7dSMjrvyqeD2ej02tqmsoKG1/T6Z+hSuv+
eTq5YuGvW62F0Rn/SO8CtPJ52mQT8AjEkI3wYX+8o9lbknvD0NfTZtJOn5pScISj
X4zxOVO8gASfJMPAKnrmkMMGzVuq2OKPQUWzfU7Qgh5UXqIc46Als7b2F5slu1aF
XWEhB1ooYwQx5dgf7b/QE5J0Rg5tXsP/EyDHxmTp0zPfayuqsp5SBzxcXrvBl06P
gsjDj/N92Sxotpxx0OZ2JEf3Pbvx8/mEe554JvZp/w91pv5FMk+cq7+rYTFZzmjE
jkd6zjRck38ZQtuhu/FYGzSsqT9qNz72w0dKKuDCZD1Kwc3/r8GcS2uWME34AWcQ
eNnLoHbjIC/5ze+mGQ5VSbu8Fofcg9JxPyFp9S6Nmwux2q9/Rmyoxt0J/JTBfBaI
5wrJ43dv1Rl2BHo0ln2Pp5clHnVB/0SNP2VK8ZRg2gnlzMu0WPbSjgdWyBm5Y+Wb
JBzXM8LEc1rOBTEUSG73Vn+YFd3iQjTOl0V1OWozJOQTxwifLJAJSS63cqRWqJGZ
J2LIRJu7BCxyb8QsDxVzGUY9ON5IJUCyVjsh4CabbGhC9lvMcIGSBcZSEXvz8dlq
a19e8g97x5onfcAiJbP0D1qutps5TwEvn9k+GVFDU27hy+px/k1ScvVgzyMLlrT7
bNpdKFfY7v4ZLW+jk3xpVBDjDVkvhhD3kyYErSwRfvgipBhatBGtPJjsjhplx58P
dCrxJKvdlW+LoQaZ0We49/uY3zS21oIUhKFLTZEdzI49hXmdNFS0AYsb08obQ9Ao
2FhNK1mbuZ581oH+yzrgOkrLfTVrd3fcLHxcejHxiD968EY2NFbD+WxYc8rY8l9h
Mh/mFMKL1gC8LO15liNPBQmTCQhpZJxt540n4UV3loRlh6d8ATH918AAVsjn8GIy
EbAaoLDncNjCN2WeA7hJ3ZFXt6OswxlGcIpHhp1rPBVeavNiqFZ0CPZIn8J6tOSq
yVsu+AIvk+bN41o5zRGYELlon5h5js6eewwoUJWM8dhZgpCVjK7KBWbwGQh5FVDz
xzsy87+Tj3OAKgBgMzNkBgqk6U7v2ZnTPm8XrwfIQvIGad7UrhgDE/TfwUZpad+r
0RMIDb+eOKIRZdQbdNspeeZac8bzIRh8M0WKFf+S0D7Z6DuwTRlShus7CWO1Y2u2
WW3Oo7zxJFSrvP4z+0MV8fLv1bkIWjs0OVfcBIBcu1xJLLhP7QfaLqenlsOsYwvQ
E7TGv5GanW4+hY2lbVOcs8ebGvvZ9LHYD7zBEfpQ3sayjawKKD3tFMu4ZFWjkjnQ
CWLmE5vJcs5sAmnepea7atti5qXrxx7QoImWLFZsSvkIpJIedR8mqmr4+X9OWfta
vKTtf1jjCNMONeFOJk0r0yDFeZw4XtIcOg0aLOjKRkJAEWMVJX/iGH5F5nk8yU+C
8EzyU3TFmyEY6G6g1j/pCkNLQ81VTeq+iDanKufMhJQ+HDVX3lIVpYaosJCvXRfX
tV9NaMCmZxefZGYQ3VnuB06L+v7JwkJ++sM5foxmYQvxhYbaaFsxk6TNEUwuJ0kT
R+7XZokxJPwTD1ctyIUZ/FyDEHgOFyEyZWVdrHTbas1prClyd/jNbl3PcCAuA6JC
sKrrheMEHCqlUgJSKM+GbnvsYtp7Lzm0bPZaFdXr7oTqPAmF6iPpcMHgUp+7Zvut
PGip1+J6N8loOwX7NNv6xA5gC2VSPpAdSm5gD7aTTHrmANJdduHrBcDtWi+Bp1Ee
cyKuWDAogukTVT0SE6dDV64njgNp/MGMgM7BQQcBVKd8ejMFui/COZyWdcscZb1m
dORY8qn09/y3aj5hMDEHPlbgLKxOTUzueVXAA/cB1c03Vpqjs4sP2yJ9A0DaeRD3
XMByv22dUXssP/UgSYicAALWcnRKPTt2+K3PbfRPrwJF3QG+3gd7nw4Vew3ojzM3
tgt1p0rFdQ++kQDyWSFXjAOlOGUeg4G/nbEaLJyFEcqphOAI2Oq7rGZYUgWvv6Rs
GyoFOWg1YIZfITYhsD1vxgHq4GnO49DfYA8DDYduhw3AsJ4eRMPQk1xWechl+ZGo
FBinsBFgjJyve+XDTzdYejM7xXeHulBbLMPoVo4wgUboj6jyrBSqDqYndxAR5fo2
3u0/QHxjLmhwDNDWmbLFNfhD6Z/li6x/CeDVQKS7WM02TIl4opzvjRNhIdQHDQRy
LpftB8DKE9I2aZ3txVHGCLJphWYyfzTBMhjVdIJIH+M+fqSWdM04EfhLqv4+4NZb
Y3akH1aHSrle+bDGIy/sUPMVtzqotgjAzUtbALlrnBjZ9uZFkREOjNCQ/qn5ECDu
bcWTAJyLZzab3EdNaJdkX+YNcrWhpxNPNwvArbjAqSa4koUrqZ+TcYcyye0N9j4N
IK7Q3VDvx/npyRGd03yQoCVC4fELh5bWryZmTlBToUPxP1VXuj3/gJkxXcXNan7E
91H2qaHfMhm3CSLEyJsiyDsfqhmX5SBhU063mAlFM+a0wewvNKCO7QAo+HiTITLm
iyBwoM6lwfdxt6c3p3/sq+cEkxdYR47xVuEueCwFkwsANdWiLM5xD0o+kKz6jqfd
w3iJzYNhvmtUNdGQ1vR4/tW6JjEQRx5Mx2KtH33hGLNVWLbJZMc7ajJVoOakFroQ
3S6VoGZlGZfBOLADS/eN4GFqJyNd3C9ljxOTW1Va3J/Nqe3el5D+4gz1GaJnzD2d
liWF3pVxS7Uilql0hgYGfGEwNoT3M41BiLl61gGNggCAqc7ipxZJS97y6Mt0dsVW
WksbcQmSKiUM2OJ/OstrfQOqZWCooqCmm16skJLpcORQ3oLwAe1+9yiUZqqdwECW
Ez5otoMBIW8PGhXmBvYZAw5UnGoAE/aixOFOT2CVTtHWsGmsa5YnncL0Gr1K4JxG
5kD5oCA54/AaUvHLcwACNSxvinK3XyPPwGAl3KkDAAMuBSqxuZVuLqb9huLSrP9F
JWtX0WGIFPEpcYkkJMVhCZZ910uzdNYVvzCA+WPEGsg6hpwZi/+8+McaNeHx2J3V
KDJ9bWbbT9rHiD11XR/+sdS/a6xzIQgDYUNkRFv10Ji2zSBlexg02LcNW4hgeaIH
4b2a1ShqJUImj7U2xKEeCYv1tU9KpckD0XImWw2VgEnyBTtB3LpsWRkkieJf6RN2
1nwLRobT5oJBVjQ8O9oHm7PkxPBYBb4YsX1jXrilpABVQCJ7TcJc8e4PGRlzmGh7
vL348KMltK47BjgpLQW9IhKfQPHw/LlSj2MbkFM1RLNEe8ghytsW5Dc2O02AedhP
ovpp+uMIS1U4BWiSTf3131RsAYFSFJdYxmdlcksZQLGyUu6Dp9mzI2ScDVxNOFYN
ZZz5NK1w3WCVFk0LgbVIssT5zQubnkLN1JSBLsRseAJMJyNO0kV1MKxysxx44y1j
uHPDzm1B65sNMeO3BjQ8Es+YNYANrdUYGA4NF5d2gylPTi5v3DCoFefX/6EXdI6Y
2MMoPNm4gEDL/p4PtFpEDw0v2CDSB/IlgZCPFHBpBJymuLa5BmW2EHUQZPtGJzdJ
uKV+zv6G3YsylFYaJ3lrmy1oSm0u2rv0n5HXup9GxECPelYBF9vvv1Oo7htVacjc
2WMrupDslcfMw/HGG0MjvZ/Au98oOPGgb9pESzLDpytVUfNlJrsV6JLag4env6sH
0bLeG+BOJ0uMxvCDgY9z5+4aVqaVF5znLzB7cpCAw0x/aId80lJXLJkStDwagKWi
9LNl8kmVNeCP7OQ0CsUglVJCdzPXi61AaZitQ/skt2IyRHmhesO/tRy4lu4ihLNa
4v9Uk0oXsRssB9Hb4zUlD3VcEKOFzDwWlU2J1kMwG9oELDgR/Hus2NKfnZApCBMb
fUkVptwY9aYtpBVGpOGp13/AUXrbe/T144fF9o++MUclcSAqMQx/wNk0RMxfht+V
cy1fmFN8kzKwpneWTFTp7wVMz0D2yZ1Cwk2M9r3RTQSoHSL53Xz92SA0XSGIWngj
zo6m1GDhwnz6X6MIheC1hIyEuHe1mMGcJy6jjcChAnbwKB64DI+1JKgMhDZiGcP8
vb9+1O+0STBNGe9tXLsbjOkjO81hN0ie058pO7sP5iLNE/5srLNq+cT6ViqoF9jT
oeYgNMza/oSHGoqSrxFo71P41fju8+3oMs4uwUA4cmLYlLAhw5+Ksi1jRxzZx9ra
WyJUHRh3IUwen0bdwuVygA17juAPHAIBE/VqTGyrWdk5mXMCqDMz2DuNgo7T3/NL
3htc+VfuiovsDKsCNgVbUJVDjV1tPSL2l9dzi/p9/VoWz4lED+Dy/vA8JsK6FtMm
ZlXrWRuAQpmhrl6yzKsC6eHchZWyXgTCeS67ZM2Odrm+/3xrEmnP7zhTqQJ8SvKb
izcTJmEQStCLZUe08DeJnjY/ubLxVzpqxTkZIXYf7sZuR45s4iLI9GhdxwZeus+a
YwY21aWkQkq14DsDONNo2lLDPkalqH76anWQ+sXZCxP6l0Y4zlziB8pveAeA33/h
weupcQE3VG4PixtmLLTdFNG+wBouYV03+P/NOd9mJgmr4+DKTUCAY3wzcJ6sPgz3
wWA3jxYw4hyAP+NhqKlciK9EbaTIJbWIPhMjtl44FS5wxeAy3bB5UEU1Tpy2LkIm
3Y8rTIA76J05R2BBffwzfayVT8xiqGEk0ZdrpLKL2XsTSQGnObqhh3EaUzzng+Zx
QqvdY7fIUUo9QC7neroFqsBKppUrGrZXif6mTksn47rZY496oQaxDtxgj+gcc7v0
qRVFdYndd4UPzZOXFsVdzIoAadWH475cQ2OdI5Hq05JUC/EbkIRDheRPPmhph393
UaCMu6Wv/M7M0pL3GPiSkwSGF9T8Bq8zK5xYozM8YKbKfmE89Qz9I+15KmySjUB1
BcBjz42O7e5p0l5TnYxzM8/gxT3PMU4SMqSo6L681hjTWRVleRoyW2CcNsanhr7V
WwQYFkCqz4GeIU28dxZJEIgvy3rRfg4DOaYJF5SBQIZ6g/B+lUq7VmnARHFo1IzP
tZIYHtp6HZ0PN/bSVBYX2zRuoEsMI7Apkl1HKEWw/NEmB4qqu2mRr4zfapNkGWwD
eCcJpG+ObM+TRXrXrvyFy1HNj12fMT+gqNW0oHPVjZevZ7wNHemEBakoBnrCNTwj
x3i+BVd5TuI55R/DNJqlFeNvQgvVg41yXRFJsexAjzqJy99izwuXfZSywHWFWNip
edafVLp1Q/JKayFLOx1Sn9AL5oJMRcnFXgkSM0YuOKZjF0uNctw2a3QbFZLIFYv6
hpeBWoKj4bo3awk//iuZ161NJgkSbWjh9472flTyRHnKYQ60cPMFyBVwNoHr7JW6
u8GWzI1A3RjsqzKuEiVOZdGR9xBy4vX46fdmYRT0TxFX/VtWtNGWVXCy90bDAl5/
DtlwBAFKXRmtg64lnV5646DLRVuN13ZPUJegxSxIgAP8Nd8iJVKDMwtZ1PCWFa76
MlhgaEHjpnPBBFRwYqvLZh++dBRsrKXGc2mcJ8Z41jDdsd1dpgGToJGju03+u/FJ
O1LE6QB51fDrIR4PR9/sOS4HzTsst8ZSRCjP+ZLrUKUlHbogM7PibnRvR4QV0XDG
rmTFLRS6v9cFCbmAxTELbafbDQ2w4qM3VPlfjcfJ/zugSmePPxKINDypxAWSZqNt
BhHXEZhczwbTSXVegpjW8z3yLJjbF4BpoI5ZbRKPNLX83NQmcrFlIN1rilYPCCH4
OP36grflMvm5lnUCVH3jDzervsAEaAVASp9Zx7GKianWCexskPjsEAJmU58rf/Xe
4R50+VBL0y82tb79+iJl2IEbLqbRQzb9CV01TdSPtXWt+FPg9GyhUkJRdz0FkUze
TAxD3Djn/BscgyWK70W4nbZN/7g117LO++eeqLvYWZ8bLheaST1krwv211n8oKJ6
4TE50iPjWMbcQqPCH7ZNGAWxQhIhPmbvQT+5jBzl8cv+z+aGiMV8y2XTu9KP+nfh
h+XkFS2POwJPR21mvdjPQfeNt3x/DOCwyQr9TNFivz3tU3TnQng4m/Zg67RVxZ2B
e8wTAAgOUmpOMS+AZlxCcemRhbc+M4YLm/OrytWBkq+ctHAh2bexE/etS7uCQqVU
hLUFzgQGLLG0AMZcpTNH0L0RA2qGEb5sYliZuqKCcxKDxtVTXgV99J4PfqZWZnd4
hjDGYInShiJlzoq3KgIqTL6hTBysPT3/c4Vtl8b7A0pRWP24lVe6dzv/zEzZkgCT
C5fT7V0bw2xAiLYxTg5pz2/KUa0jak7ucDqCBayE2ghJx9dGbGzVpYLVp22Jrz7w
sU+pD/g8P9eCiFWPqB0mKJ98sSryYTa9JLC0lKfPv4GaFqXb2eBzJVtU2FyIifgy
AuWlNx6OWRJ+o3ExpUEH4vEULL+f3Iif7rdKd4jwFzoZI/fY6TzkMqCX3Q3cA3+3
i+i+ptMD42WupocuMvHr1j0NDvi+UqyLZIiirF4f6NEH8jhOZbohs6WdXnJptCpC
wQ5hjSC5nmc56tdEKmzg0cSNGpazoYPPf7kZ9O9xsHIMPsCgWRSmm2G+HGchTGS2
RGxg54MGVQIS+UZ1AEEB1p8ttdzVB3fmMoKVSPlT9sGoQzg32oEA+Mwb0w0yDZOr
f5gFdPPGi3ocil1S7Or/WvoIDmTrF89/K8pRqHFh55PRnei6GsXywK15RRd1gn21
54EgJ4pYYXhWV2BBuoU1x7Bv7w/JCyshEKcVjcsRYGpuNPy1gxkmiYwoTDONec5E
3A9dWC1uZPw1e+Oo7nlGJB7hFKnHMu+ViozY7LjLChEhkZ6v+0GQsvjkc4bPcjJ5
RH42EULxR7qa2bRjq5vRCd6ez5eDhk4uUuvQuM/ZF27n4eCMXqP57rk3b4mIIMz3
g3cy7bQsH9t/dLj5grsGD36u9lCECNXMczcqDr0B194k9b5O4clWBSPVMG4wZWEy
XcwSkRCXJZx6QNGTSuiL2tMUU1NcPWaayEbi6XI/Bpt05JDvDy7JLCTHaK6ULv4b
XNB2NFbgjv+Az4aNlhJluZQ1OBEhzxF+ml3vpfSdyrX14HLVaR4zhQPqrxaJsF9H
mxXERBmtp+end6VnVjQBbbbBGZL+KhoO+oGpeGu0jchJM7Frb0zuiibZo6e/v9B1
CQaY/POjfpzgFMUKYbP7dPvYFFm2Zuf63iq0mV+/UJtzU80KAGL8iRaEhsj2dn7e
px3TRFiyKUks6zKebiq5VyOCMrwvzhWT22EWsYCoGzgd0VzmRt43P9K8quhAr1Wu
LmaiBfhx2tLmkcd7KVmSA3S6Id+7H9juavSQYRQSzRDPIr6+GZ7PUnfUb2G4f6Bu
2Jytg9Y5b8MJI7IKbm1ppyBYc/5re10T0yHbxilhVG8f0gK5H9miV+FYAJjPp7yg
dWDCjOlGLIoXd+8oPyx0Qwx9ahsWcWeeGmjMyGhgsYz7oFDiB7iEJcVgjDbhB/cT
+R55jIjbzwN0+Y1QpWqz22sNwIkwNSKJvrg8tY42PWP1ieWpIumSFG+6FFjrinpH
eRyDIP59XWdbTzPHH1007um/61UofxC7cYAJM4bETgEel8LiNfwgrdeVeEghaUGC
WdU4NduOf+X2nytyW9YB3gSfXpqGihnpdQk6EZ5ck3HjhRgF20PD/Ri1wYzW7TsT
z/d8UPk1og+wBKngyC6DEvbGPtexNxgPfDj3eUADwHt6nk1I12RVshAPWCzjesl3
dt56wdaYf2L4u+t6FL9nAqGudXG2Uyy+oy/mrWef1fVBmbRB54KEpgX1nZNmQBOf
2pzEO4S7zcZeqTkvEMDc8XtPNN1nL1mZ/EjE7oCOCFDNroFWfVp8giLm+BpiAsh5
6QxB0No8cu7IrIwIuJMX2BZqfx5xWlFDcZo5p3ViXMJk1AeLbSH7fyELmiZWloAa
/Y+PeZJ12IRpN4FRvX50ymmm2R/puxMSk5QmJDjCX16AlRkn+kvPXYza5RVsszro
YY4N10SsK28OoLdEzBPj1S3sx5lDwYEZJMnzD8Tyu4sZyZz3CHqkyhuOC2qt8vQN
T7utRdnTYA7+mIFN5gom1f0HIecXnjbzPlpNcEM2kQb0KJdByyrymTlKagjFY7uh
cV+sIkaAUaibYFi6f4B1dGwDT0TZoHGRTKWAKkbPFi+E79pk/OgLLLVVI+M65+2M
n/xVp1qH4EbiDUjuWyso1edWCPAFfSN/VJmeViwaXp5y6GV4ifpzkfiHjt6TEAsM
S0R76ZCmZUUIvR+V0UhlgcbqEs2DfymYb6vcRu/EJAojCZqmUJ2KkS1NBZGtlXyj
A1Vq9Spy9G4/UyycbXTTxHOCAx+1kSGDT1GSgDeHcVJka62w7DpGN+qt+C7ovrsd
zsN8qG/MpYsrtIhN19886gao31ug7W2V33uOmdgSaFPI5wABuOiS9guwkRE3BsHm
hNwl5ik+MgZ9XN012Fe+dHNDG9/O66BmaGEELQM2lU5Z3kSGYbNzE3vkFwzsJB1c
kYZxLNcdQbPz+YpKbqoMBPxor7uNae4rAdMOSpS0fYQ30H7J8X8Z4w2Tca9SQncb
eDiAVo7VmuCBeeg6iR+EFFSGHbf6XyEC1+RVRg4+eSIpcIQ+ARqEd91D+q9WwJXO
JL+4s/D6EXE2Ww2O0yGslXbOPvIanCB93fgai9fwRQENoK6rSBuAeEtQSLNAPG5R
o7rPXzlXagxFyx9H0Pi58D41hIpdNREhn8cC2VwSy54xgNcnWw/H9D4Wz3CDQ0qN
3x1aNRZnnznPGzesuhM1h6LSbs/ZyXnfkXd1eATjsU/haRM2x8m76Vu3C55G17Ha
jQG/myqpQOH+ZQbvmlxuEo7rX0afB8Kixfgwwoo94I9MzClgMYYtosOZH0+FEXVF
beNtGdHHpftbrqc68xd7tRXlMgrbeZal8eiTsHaqO4p0pLTFvw1BF/t/xVjuGNXN
uaKD3V9f138QcULXUzkzqepXWXMk1n2EPZLdSgoD3FWrGwcjeuxaTqU1PJ5ln61c
Cr1IxGA2wE6xLU3PqwKuGawMkI6d0odYuEWYOJC5X8VIDraYZ4ggsTdUS/MYxYBS
tLpE4YLhKwvRIT7ZhZ1mM1iV+i+xFBy8mZCyz93JMwVRB4npJ7zG5ONzOVHaZU4c
ZEx98ISAJ6TPMUpru0+o4vuCh8Nh2TJW7g/dpk/oly49RdV+DSBkr4n/he7IEVjD
iIArsTCwYzgr3RX84ydP5KSBZI7Wwt3Uvj1jlu5rD77XFPkqc9iY0GdRikbO2Cn0
35giQNRLyzvNxtUWpYr+nLWJfy7tpzRCaN2LoiSAGh2ne+pzX0Xfsu8g+eGVFjuv
NDRU+HxlOm0shu/dVKTdOn/N7BbZQUt4AW2PgGfOrQnK0+m7a3EudPnfQVs6dt3j
ypgFHeD0JXOuJQB8PobwhyLB0GkViUbQlbMrlNiJkTjxYCubMAeSaOVRDOCWTJHo
cOfxIeiHSXX2aZWy0ACaK5fU6UW1HlUQThSyrN5lQYA33IS06CplPKXpNIYqEWLy
KeX8ZeO2zIB16xxo6gz++lwuhhZcijLyVag0eYaGFjGU40iaXPAcxnZCj8mgI+UT
z4NHXSsbJKXavTaiGdRtrU7ubvGPtfviugEoooeSfxcNZ39xjo+nYGiSznJpJoZY
EiTJezt6YAw6nwITOWnlBUV2F7Xlj6DsKf5kwntc5Vsx3iZ+GOy3XfEAsjIm5YtJ
woW/B/LkgU4LBmLPkUboc0V9qrLlUET29ZWXQ1uElXfnBdLpeIXSUehm73ZkhFss
NNK6abY7RGTqdp/oFKTXh+9y066yS3OcO6KZzWCnwhTYeD1V/Cdj4XO4fdQJD+PY
HrCa8aSvuBccpv6HGVCy0xtNXLo+reXtiyXaTIMkDP4yZGt8ipafpTFFPx9+Xnzn
48EgjNU0M6S8kA0v0ZXAShkQ20vvS0BDACA6eh4uq0C66fPVECmB4MJ9+Vgn2e2a
+rU/mk3m6gLjrgdDUB2Bz37Bva0l+Ug+hMfGQ+Iq5mhucyuSIYcLHgBzmAlqq7AO
S7Q2sePBzbtkFOCsRJcSgqDyF1B+niI5jLk2vpRjzQEiFCEC5XGXALxaN8/EvxB1
+AjeLkyxJHoq7665kkgf8dHYwgP9pedpWCzH4qvGwlfeSsjEyMoQ2F6Q7xFqQUfK
/arx2T9OSppjWztyB1IE6XlKCHCPGlo9PbqNZT9hkK9khlYpvV5LaouQJwIBFOyL
EzOLgXmYP7i4w6ARLT5PrVc5yP2bJkDl3oPOAsLIRoFwUY3i+0sOU3nWvPN3vDvM
kCa/QrYrFvKaKTpRkUqDsOO/f8V/wJYa2niqTyRt0aY6F3kDMTKZisb5/JxXfQGV
/d/O/JRruywa2ElEqVVsbFvYbklTWiwTQFLujxA9fzpQr2Y7v8XJ1VGiVd+dkSpN
HwTCvcPilbzpxCsjg6dlHW7OGuW/KVC21oCBmfGAR3yCIlQ4GpsOdpIPqYrBUkJk
IuUQZXD+37xxdy8sjnL5mO1w51tG4focoTk5GQea910T2ahNDUPtSp1xLBvkklHv
ie5vtN6kvW/rla2uG/Cy1nRGKW5o1Y/8VQayH2Cp65iUjzdkFMqzejKSIAxQiwHj
TH1WeRj9XE3YDPfYFCMHkPgOLAbwkLciy/4qBH1Lb5g13MSO8GZQvgdAaf7Pg2cq
DiWJcuhFe9zGzr9DPxoYU40OeKi0XVpqRsfZ/tIcsOHrJgLdzrJiQTOS6ss/jD7n
vYiqjtUP89J+bl9FuvFj5HnwQaMybxe7qT7c2rS2kluDFrbgLJYk2qyiPZ9hB/H0
JEaVfbPo8gqMngJTOpssznYq/bejWvyMX1ukWASBJunMguizOk6K/9ATJhdASDOe
YCHg+dm8tQToEHOwkFtgAPOvSh37osZlhfMW3XNZK5rxlDr3xk4NCMvOtRcWQh/P
PoqjGJSdfhJ26s+eCq8LuQGfTU3fMmA5HgOD7BqfL/bfa02p0RbF8Wzle1xY8Fdp
A+ummi3o7jiLQV+F2yYrC11oIDIHSrybXttbhMxCIa/NXu1bUAfUfyEy6RC+U32O
qzFJ1w/tfuMTuwVbscZZIIOFKm8I52Ytr/U4wMZKLXSt63/IOc5PXMzEHJ90WTt3
gMX53ilFKiQR112ysrT5Rzh3A0P4v06+1e/K8VpmRldy/SBPbbQOlUzK10Hrns12
n7jkBNDWr3+RVzp5lEbqexPgncwES4JpOPcziIgUbnsFCAof4xn30r0UqC2S2+1K
GlBe8mGhWyLyWmGKqWsli6FynzEhEgSI+BxrxcdphnAk0/VP8KawYscMS7BQdPuC
1S3i5lGv7vra/e0FbL173fE9vRbeJ+T0yJN28iPGdeJrIdlFsfjppLx6lUQh01TY
uiRzmaVKdfH9t2Hwa0rp70O3UoQ8hgpIoGaK6qvsA+QNkuyEqjBJ2mzdnH+hkAgd
r4V0eYbyfDrJgDBJP0mkOeEr5touOpIZy/+C4kH1LCup3zc5M8Yg/zNaJrniiZa/
Rb+QplsjJMWnF7R7uX5B9VHBQINP5jmR4Rjuwcr9uqiyQV2tRvOXRpvzNg6XNIUn
RCFywHizvmfzPHozvVuXcfrtxY6YKvnLDps9KRHtYzmXhZtC/t+oq5sL9cIrT91B
++7T8X0WxNzunq4+6OPG3/1NLGKZcT1sDM7n06jkBAfqIhVuHrDQfLraUW52yEws
Olhl9KE6y4U24MXZ9o7dItygCpZ1apT09wRXoCTb1XJhfmC8JJ2Vgaht1pbuEWfu
eC9PZaDy+EpRAev9BqiBuPzyQmbSWxatjWnSZ0RrePWW1Tx2GO3z98ks+mBvsn/Z
X8xs7NgHgUZFTj2OKfS9KVlS7ZpyObsm9lzSf88owDe5CZaydjYCzAFHYMI6uWex
LFJJeEG305j2pY3WBFF6sh9L+VV86SQdEnlGDtX02VKKeIt1ym23KYRlGq5c7jHp
u+xahrLaaQVJbtnx2h6ycbx87mKe2Z3Q0ls/6cYxYmrk+5VOEUjJCpVMOO026u7n
cP8yR7ST4k79zW4X2hbet5FCIPdvn+q+BnXA7/jFm3nzNncRT2R6EAZ6A+p5rj7m
HXjOyxxdIvkv4ul3ayNlt/lUs5xGNmHzEMHwXfLmszg5G8/4al3GWZ1RfJV5Q8kx
nDtl93yhG/Apo77tgcOP4HIgYEq1BhCF+mrAB2crxjG9Y/1u3IMGhLeHXeYlfTdG
VwHU0Ur5xpI2xTWlpFHSVmUmi5ceIPAb+/L3rIR7/+yhnI5ySvNIqSoVS9MomVLf
MJ8ofWmM+u05oGWkBFeH0KrSeGNCLhCHlso4eFJz25nz1jSCOtvbuk3TEhd/lajd
vs4hWvAUJEGASYma9s20FwB4jMIvqcC7VgB40/RXmbGpjXAPGXRHhcZQRNg6ZAJW
RDDgmioEuUDFjm//2TLn9bIQA0S6fRFRlOD5qfFON1tXQHbwkciAF+fSZDnjM7QN
yfBMbjcJju6Dw8rIzNnPR2Uvy547PG7YI7/k7irZVs2Wfz8bq2PwXQLOKe/EFsvW
PAR9spYHEspQueQXPRVzaYyW1f7m4kf+haCgALht6FlVlbPHdwesH1j4Fky8pPXT
Ii/+kNGXw1iLA95dbWJE3Nlnt60twdIlumxxdQL6z9koT67qxwKhE/W7Zshf6zDu
95G8Skv2koX7UnsIxrQD6ASh4GCxU4pn7WAl9xVA1cpy8Z4zzjlRb0LmKunWLwVU
j+zGJuckJhHMSwsLqhLcSUNtVOgQ+B+aUZOoyomIzrV8MQ+ITCBbpVeeWZVzYW9z
pJhNFJ3sU+gGJxKBvn5F4xZHk8Pjf9n6jeD2phPEGaqmGl0hkXOgNmFYza6JUyrZ
x7yfQj/qTcdq6yfyisOVUoDdMPmNVCn0QKX4wnPpebXRPTKBMP1K8VrLyTwOCnbm
lWvizaCDELVM2NP/I/+XMWO8zZUoalXopzk+Oze3UnxSJO4wS/5ZDFI4wvYIiljC
6TTardY32YD0w61mx0P3qv9IwiwajqM5zlaL2nIuehPn2UYmPIaF6xs0JuZtHxMP
jXMuCEJVY4wpSTPiuoCOEfviri+WluVyuDAgNp8VWuYJZf/sNnf3Hs2kK2w6EBI3
wPMua3a/KjYkB1rNIQcgG60FrH13F/NZYjwX36b+pvJTNdwqbFDN8I5x7AGwB933
4CgolyNntcpCB0apsVqlPLQiNuXUkwfomGs6oKmPNWyYkj/rRjO9iSbYpWF51WHB
WH+PHhBHL1NoaSI/BihSJxtwhp+UunkFJhPj91ohHu4M0Cf3nncSk1b4SjPwgxHe
D7XK9fcd8awVVS3FArHdIX18EfV/jaFGufhHn1Xp7RyhgOenAqmhHnbDVTP9CyzL
4CA7xlSe+kv1UnH49oV21onTdqaUljRzudWOUNojGqePPVe1JAZdoQjIapZJaNu6
wSIlutT0zW5L/REFC6ZhSUqHJSJ4AszjHQ0EUMS8lqF20rus0tWzBddxIA4QxdDm
H5TYmBUtZhyEanjq1CFD7uHftO+1iCiQl7KSkwm3FbDwNt9g2cOEfTzxgMNmtoLK
PkU2wJZwc7cRBRJpV9O+iBD7TyUbrhHaD+Z2qey6CvI2rwB8knSI0Jpd8f2V63iE
cN7IULU9kRRFDPb1tfTWAdzmUO93noJ0vx+4ktFXt6BrQeFq0dHiPcupeKGbldm/
Wx89SHUCOZ98/PVSJ4X9vw5dTur8xNWeVVuSHEyzmBBBmzOCscNRu4Ikw2pwSxDm
Ki/pLq/y83XLV4eBddDRlCVSjVAI+zD7LPg36wAOt5vJB/VuLq5MpKHAaURDzNua
kEccZs7l3b+IwBcr48RB2lPpLJF7Sq5kZUY3OhpgFxJyGReWd/vFYja+JObNOE1R
gyuwcGxwDGb6lw4/593wKPmmU54bvbQRLQ6XBuQMUQQ2LEnTZfLTvmTchhRdNzHt
OJGdd2xJWgmireunhO0aNphIpB7x0JoN3y1mJcV7H302WmxVzQfndlVAT33cgJci
pAFCN0XYXHDxfkpGcCqqqYPr01iqPBp164Rb4YR0aCIRxQwLnTMVQFv1VMy0zs+e
kkfEtgqSnPvbtpdEiPoHPrPqtZpHh5ZkjeT2Vlytx9zDus0I5l4s+8MNXErfNMa9
aSDYY7LGELy/+3gOXqUaf+RC/HHcqiEMw0McbuRYUz/sSCgaZbcvzsfZZ+ntIHEd
HMCgWJhGru2/765Y+Gdgbg7nrWEqq0gkOiKt5dJT8P3guXiDJ6ayyp6qBWgXJh7L
MEto2uOhsU9m+YBkmSdscSKDQldea8YSjcY2tt9pqxp+scFdj9lNFpgvNY5r1TN5
Vyy4y56J8VX7OwRVq1/vWM3f23mD84E/6LGYJwn8I2QNn1vFEzPobfnhVpiLzPzi
xqrWuURnyF1SguNz1ekE/jvTGHCez5b7GqblWWD48ccTr83MrcGwDf41cKwD38kp
wRF7puuVyMxRXG3fnbJ6Vm/5YOqR0FzGgDDUNlyWkdfIa5AOR2fPU74Ri0NmyMR7
F35MkZ+rsPV0lyZmg2KmabPdKAHf5T8pGLSSNAUPsF4McqjmjEElSMCIyokoMLss
pQyK5vKmzq3SHK7zgOz3SavXoxDJOCsLYmOgRD6TP905CK8lLMCjypNP5Udhz9o/
U7p7ME6PFqZ2i56I/E0I4ZjS9TQKbdBdldEJmng5qH0cigTiCVhnTPYW3TOdseo9
e8B1VPbmprNxPEPTT3Oke8Ces0H2UsiibxoUkXTtXlkdzKTx8w21pPDajjK4AWFp
cHYISv62K/N/bQtGL2nE38VXLtJE0JqQWZsG+FtJ+P5fbhVkv8JTmcZA1oKPFF+G
CoHYUAHeAEbcwBgaKo6wN7XZEYruWIavhMUPwWiQIAhSMrEle+yKHFpHpkzJKIqE
aVRbXTSZHKaTmPaXenS1a3QVpJL69ORDDS8HVETss+so9oCkMMpE5JAZf7tsJ9nr
xwuZ7Lr7STxTbNP4i3dc8XWPs3RAFtmofFJROah54Qf3HM00GWqEHyUpx1oxeHlv
pVwWVJly5On9UeskeleibnIkFwVdvFZ2rwO56wa5xkVCqKa5SKX2oy67zOed1ZXC
6R4z0D92I/t4tXK32haVtSHGgsKY4E6XJqsHbsf02GgoBQcl/mJAsOP59CGqpjXb
daX8/lmbLghcNRN3N78mRduZshI81DRuS9bKWO2BSJ/EixDuKms9klo8h70465+K
xpS0cimczeT+BJv4YA1RBMzUc9y9GnspSaMOimVTEqxQAAMKOHjNGa4rPTDaTkiI
N6JXSn7i3lGA+WDxTdMjpbUaKMT5tlnzf8wQbFQ2xbnjxYdnWyCAeaY24mS+D1Rs
HPO2rtSspUjAHkI9ecXiymI0LH74ZHMOAMdVnohFuYhhaI0DI+KbPXPv8Cnm9IL+
0nc2FSpwliY2hnnutnsTbelSuvBaThKyQfxtlnb68s3HjNw63tyALA+YPVCZG2jY
6BUhwCyoACv0DgmibEJn7JQ7vAu8JBUeliNQ6O4MjAO++tIj239Pvojp1F4fvpzN
lntL2KJnXck8Z1yfjG2b2cQ0LKQwzsgIehdUkFMErqDRTP8gxDST9391mb24siZ2
o4nfQ5Nv+Fc+LDvqgbhYAn6xbauzX2dqJdPZ6fz25d60BdZhGrhSEu5O6110afeM
Nqz3D5vXSKye8H6rDRzPvSzdhosd1ZtP9MD3BPM9dTlfYPABu+NDR1JEzrVVcO2i
I+Fvx8QMat5YKFt3ZHQ3kOoUE6zSNmaFJRR2ZdJfMfQVkV42pAAC5Fmtjz7I+w1G
JIJg/w59p47Tb/75wUcGQw0GZ9XEYEXCtItRtk4u9C/5cr1mOgU/SKu+rLmqUAWF
IspYxklHn13qUhVC11/WydfaPJAkOI/956BO5HjmdZJMjfTVski06a2CG85E5Rpk
s2um3nq9vtLtUNRnaU181PNyGdgLO69je94oNyfu47TUeW7/EZw7KZh2o6jmEwfq
lUL1TtdYXz3k9exYUqQirGX15Hs0SzjnlMoTl/fWQ2RyO7+tLA2iFcBs1GumOPUM
gDU/VDMnOZxjMMKahD6uKJuw46IwEk2t2KDqtxHCbFCoRpJ3bX/2T/l+qA+WKUnj
BHc+amqaBN9hKE+ah5hgt7dS53Ohn4DVDeO2ByBMR5V5e/iisu7Aq5wQ5l5h5Sxd
hsKn+8AmTV2SZkiF2WTWswnTYSp1bKmCWl8yaSoezm+UBw2Hsu+kZVj8HzZDnXbU
/np8+YuqmXvWcSOHzwAS+becN/dz/AXW2oez0yb3kS/N/T3Vm8a19/ZfKtj+seNp
07+Qq5buGFTd2/RnPG0ykz9e/XX+vyuTDTi4JhPfznat6Ksxv7VUM/4MJl2jBdPM
dQ5igX3WqbkqEPG3eusOZPXx+TiTiZV3henXqYKgrSNCwU0k8TLzpKDkrv7F4tO7
DDEp2O1TAzbX2a/P4efvWpNSq3EsbNKdv0JrRtgPoZjdNSXBtavEHpV3uZIn0Nel
+sJmtctMygsBDCLCgaOV2uZVYVqXVa19CVN/4ZR0e3iAnp34e/dwiRiSx1bURJCd
MXpEIYIZnnQimST54lLSpFyqAk98rJu2Oamh4TSbrK29+vnYeK7iudqfgFlZLrzK
IbkU1qLzOjULVpAzbClPCGbImeT0TcC+JWYLtgzBSVibCvHbI9TLIL59Q6VHfZiy
tBGxnjqQSBEGuRwcyS9fSRUHx5AYVJyzKV+xfCh4+pDUfi6V8n2qM4EezYunSWaB
+midBQ/+7PwYU3sbXdRGya1/LqOWCeCXgM4HqYEKx5pyeAfo6BUjtnzXQlu3msAK
PACA/iMWwG1RdTSPr9vdF4cwNwyZBFvzQfxRKLx97L0KvMB1hRYNW99Tmvo7T93g
yOKccpkWAjku6DM7ZMtgS4/mGoxqU20jT8OvT6qTBCeqP0adFvjeOtz6RFNPTXiI
2G4qW1hNceEeDnGyYz43Vg2b4IxMcrAgdWH76hiJnF2i72ERwZ0H3QMEc8YJUgn7
60soZfIDG2NwspDdzjLPZ36oy7pGZteubFuJbFyyrnCmqk6Nq30/FPMjRkch3Efs
8xaUbnG3BW4lLS2kzDV4XqwgNUCxPqQwmJIvEQaweZXSu6XuygUtIYltgrdUQKSD
U6M0pCwXRJ2CQCWMpYJNYXlwuSf8cpFO5TFSvrHoeVj0MEANsICShf9e+wqIN6xQ
DvzXLdXO9z9uJXzRoWXpfGe91rFUY3khTvRjgBs5z2eD3h4YdAzHGZS6LfEBanG8
i99V7tzrE/ugLkAs7ug5+17eI0rRgZL+u+6VdfmJsck64Te4JlNbEQO0fsGxTogL
DFrYWEKVJNjB+P5enDWhFPuF60wpmCMSuD+Y86IN+cI0B1yHaPCIRIZbV6bTRdvt
DRaLGioRlyL2pDfF3JeM4HrZcdk96jmQ8o0/o0pQss20+8DIovEY+AkuIVGBGQzq
2HcPnYeKmCCUbtLy33SiPRNIuwRt+yJ+NghdlVLdncxibPtzM35lSc3eTxrISbHU
K632s2Mra7mmTCABl5QmStQBc0MlWeQxFRkv7rGya5wJp5C5UCANYgisuAXzhfSs
z87y8swazi8qqoagb/I3y5cYZ96Yl0SdyXb8QiWLtikoV+lduuGLsV5IHzWZVwIr
iwxLJyq6IHbD5mRvD345JaBmUvtZC8YKBSoVQm7Xv/51WSXS/3qPKXo/JODqNrn6
78FjodmUOdrRMdnWZlgwAV4N1aZmRrJSRN8oEIqM/Y455EixkS1ADV4l4j3biqZv
5/+NrhCAC0NC/41ghbw+gYYO+flHxVfYZAHcDykti3QTcxG5I3flstnnTyZaF+QL
jKVnxQx/F/rTtZaJfyH5O+kuucE+dvIOy19aQn8VepARxRwipv70kDoGF2VwaIso
9u1Iz0Fu2f0ZQ3MROmfhl/Xb+cZzHsA4kqTWXI0ud6THWMmLnsem4MqH4H4KbGQ/
56SSPsmTIG5kQrN+nqzeU6J3LmMlrR0qRJ2JvaI0u0Smlv0o1qfRho9Y3P09Au5c
T+0aYOuyKIs68YugikTOmDIV6JSVb251DqFOAJmACg/rtaQadEYX1Esc8+sry2Xf
QNRzl/80eYQzj0vVJZXe9aClmWlPZcKHuuN2kfN9w9K6YGNoZ8OSvo8caYR+qGWq
HolTHYu+dyPvvtN2NvTXeXHxu5MlYVYUnrZavGIkYD7kMhrZZHdzI4y4DRCHlyoO
gjxlOpBTg/Orf6CJ8R3DVeDpwOEcUHq68X/Hdo42sbIWDYQra/QwzAHDz/RCarVP
4xlh+xcNyBYq66KQxFHWr/QTMT5avFwS1t4XvAYhctjkGVGxagY71uFBWbdSQxAG
paUaqKKFTW9iZT5H13I4i2QE64H6xEVmX0O1VDOZ3IGUB+WFQkhhfaI2aG3lYW9Q
3TyEv7vUNKtasC7tjwHWk9uho9PteW/ut/C13xVhuhrIDXScHFnxjYWtI6+sRIf0
YbvJq4fG3GJkkeXjOxMA2zRJfcLAH18TJ56vQrZR9Dt4bXWL47tm9qpNz7Bb7MoC
nlhMwfriTvbPIoZwzbdpFyVMrGNpQhl/YocOiHmjwUnXFm/9Qb4gyEy8N4+9t4o9
XuoqTpRSts9nQUj+hidTiCvZDv8E5hE88/N0NhWR9GhYDOJKw3dPicBzw4Z92xDZ
iGPNTLPkk0xzzOUBQPkanXPnJ0CSwPdaUzcjyLw0CYyFYCaP9gYW1H6tEbI81LBD
5P4BsveJed6+mkEH98i3ZdzP3GuN4WWMrS+AsUcltSIbY3vO//d6/9Cw27U0O/5b
lptQ0HPS1qgQggr6R2n1JJfBuDdNgHrNqsO5oVYaCq9K3Ezb7XjrV6BYFzrv+d/R
/Db/h6gSEAKC07DJqEoSa1Jmnr2LAvDBnEL3em6cr64AGvZCiRnr5tjIOr4FmiXJ
jQzRxQJzULHtnGaIHnWSgBEYXH0w2TdxrnfudDe8gxlQxrxMe4ouQNQ/I5XxN6nE
R3I5e6cGO0uH6+/VXx5V4WF2DGJAck6RaWYkFkpYWGloKqRoE2Nju95zUREy7smF
yAWbYm+lK9+zvb5aT6dtm9fU+ZU1cLCk8DA26BL4kT30jaT/UoeCvHoO0q7RSHqp
JjeJk10d10e2YgaqKcCdn5sKlF6AzZgwAh3KhM0TbJfpY+UQGnHPUGRMbnU1IZoP
dUCAm8d8GNJifAIFVm9Jk36hWQBqBaQnQESSfr7u7YIjK0fAEwKHLgyO9BpJzAhJ
HENiLGa1gwanlhDWsZ642E/UGLVdT9kwpvvepDSGg3j6y+NHGagyePiakNJG4O3W
fYJQetQ7Py2MnVq1Q8kgHWovAVwDDbZM5BQP8sZeHqcgoaB/grkMDlyKnwTF42rR
3VRz+I5752aVxvhOg+Q2IkKY67Wj+6PSppc3tl6b7bZdT+dkSU0TkUx09gDfI+Rd
4wBe/heCPWshVagV3VlBuOPikJZcn6Y3YjaoubJn5KKtALBBJ0ruRPulwKcnDiuD
tT+6F/jYUiOVXiD74ripBhB3pzUQm9xSJVf9bnQVQbrGUmSCU2FsBpVbna4WOhnz
j9bPgTP1gSJdw3BcivD9nLGOZephDSXYD6YQZK3dlunUIkwopudpVyMeOhYXyZH8
j1Y9QQmz2k01uhcO3Ujkt9y2Dq1L8Tpgm6fVvSrJmy8yhjFIkiXu5Ds+ZMMk6qC0
vKvEY//X+jO7k0UKHx7BjQx5LepDXcwHSJKEkcQkchwSXcnAayUIFMhkOUYnG3dz
dzJoD76ESCfKc5lTze9c60IKhQsbEen1wUeoSUR7XSxThZ7T/TJ6Q+FnodvvKH8q
DiFzdE2+POCTZyIfiy5sl5vyWe7pbTR77bGyDI4cHPc0PXHnCKDJ9ErhDqkBxa3C
1qIzqwt3BYFE6FzlNPAbofJJi8wXgJG+as8uYcMbwTQaFzo8NTZ8HC3tZ/6H8hND
0HQ7M+2cA0FKevAd8BzlXKrbU6Nj6g2E9kjGd50XMDHEQjL534lV0Vl5dBhf79V7
fFdOBCeL6bOANTD21YP6FA1qBYm98HPZY3AGf5Cf2WA3C8odo7QqKpvpMICDfjRA
xmzzq35mXXrNAIM1R4K6LnRsmDflXBFpzwPbu+KD5LHDx4I5J8QirPOPT0Xb9EEc
tdCC5XsMVErnA34BFJPs1BgopcqjDOqvdiFU5v/jDgxU2e97DI371FXIBJ3inw1O
GPerTF0xESensrOOfs3ejmq/v6CWxlGi1kpYscRhIr91PvFM382zIe4BrlIfeE45
gnYUeRaWGjLUssDhPz4R6fe4YnxvDvHnEM35F0awX5eeV6/1mCAirC1G04suc20o
aTBSzVf/yBWHzoJ6dSTgGx3FYpzypCc6dv3WFQyKvXh4JMlUc6hNN6uysmR6dXcT
Q23kly6A+saeT81X4YCiXQ3YVcqc8tISGS0oSSQhkN6rmAvphQB+9te3s8t86e5L
jBHUVz1HQA42EwphH1Uw3JAdXyBEjVKd909uKDeBr3am6H2Qom2U7imNPcSJczyp
R7RCQx13wlCTRAOCdi8B4Ou49HS4iV69y5u9S96EIs8STKMNgi6sGsgjCclbjs/s
AmJstFPYP/vzc9ixL9Z/n64ny6zdDB9MHeRmfsFTG0izTj4iPbesIMlKqSgHK8po
WAGD1d5Ls3E0dGSU8sebMO/uyo3Wp8J6U0NWUERazTayrYjzfZWkwHNkwqi3vueL
O2gqZjg2zMj9P4BiKZy9OhbaGg/dqhtYYyHeBcnHchZI7siMWgtH3P3BbmHJBCsa
Ytz03o4sK8AHOHvVV9UQ/JKXP7X/ir379XOnxT/3T1tU90ZLzO9ErcV+K/uPzvmx
B9IK7r4kszYC8OfcZsBfKIOU4Zz9GX9vhBqfvPryQ/ljrUEd4WAaGqTtjuP9uaQR
sPGLwkrCguTbolyDBupRt+1t6XMbNuMBZH+p0twHT/QV4EJHmNjF9VgodlGd/+Mb
e0zlnpBsXB86zf7e5uo5C5fmiPnbIv7SsahIGffwQFo4kqIy8dAjZXVYEBIGG+Cj
iv2qQwH8sYYFJbfnoIl65F/DtVIEBY2GhVUU0RkSNLWQG2Q70d2XekZlrTg8tEBp
z/y1W6b+njz2orDXS21/LCVGnYaHDU5h4/BlIQNk2ZBlZMtQrzb4Oha4DTQg2icJ
fJwHPe+pbvyzuTiGnhOWWqCkH060tA8YAWyJ1Ub6znzgmQqgustcWXsp+R6VyBdQ
+OgjJWCnnuuvwHJ7sE3U9ip+6pQqOiBwdbdZwTG6Rndqklw96rQp5o8YN+WDIMwc
lVp2yxTJUTZ55Hx53ceHpeUA+rJKwgMQf4VWIv9uc1sXEHiElb6WpwDFS6a/OFbC
wS7xQ3OTRGwah9iV8oMpZO1pVrCHDq45vqKYcCSWy+/+wRQ/GpZ/6RQM5P2DA40W
oT/N5sdd1rcNlXqiNaE2gHvhKMGfnvQJX9b73Dm5Rg6cgAJQ70leg6qFSgmKABZb
Z9H2FOOE13CrbJyPCLX3nLlstuRE6cLifgDaglrVLeQAfYrnXxB1eX0n6QVJGrC3
XT/wUsB/OXleNuHeBAjdFtLvJXGp0AwsGYGhwdmM4rp6NCzn7YaiqBxocDEvqCI/
sWExLPWOI1B3FBYGNlTqncJGQD8I2v1Ql8mQNhcOURG00du5+QfhWooxhaFOwRcN
O9DHTdx8siG1enAsY+xxBOCoIsMMJszEXwLynxUXBjnyAdF4WCIrrf73VJtlAjXf
t6RLNXfd8sEZCWNFeTYrOufG8Yaw9mCKTyHlmR17Ypdw7HwBk4ObAZw8gnn3y9fi
Vl87+GspfpMrvXIIW08q/Mrzb4qW1saDcPqV6bcu4uApLHxirSj3QnmyV5gAoy9M
yyO50MuLnZbm/SYPDUtOV4SqMqrJFxoEO8mH6Y7U5soIoRAFX3F8mRJwRukHQeAy
5mgNDatFQ0APImWqd+6uxlP0HJXHIMkS1qv4E8ZB54s0BpC3EO4nk4JSa4ZyHB/7
+m1AN3HwlDqBDYwb/16givel1dDPjamnz/yO68ZSKmmYCfEK8XYxO5oKTXcMPkRi
N8ttMGaiONv3IExSFR5vaK5VOpZOrcwmRDOsNXmpKRM1FHj59GU98Dd7fxxeriQe
qCFuZeA5uylg+AwoSNGY+3TIjjemc5Tqr8qH4sS6J34LiO5RZDRdLF5/wrislqRK
lIS7Ick0F1fR9PPYDeUgs5XHaBTs/5/3HwquNwnsudAdyNUwwrgvLm4WhwgHJG/d
4kvO4+g86rbMFG4QHrp0HF0685NgHXtRhgskIvAtd8cQZ5SGxU85Kq4Rk2A0c8FJ
FyyczOQnOXHpnmPZ7ZAt9vrG11o6XTWzsRp2FXLiMUP3Yo6iS1D/22pS3+KxgzCP
mNYk5k7hnQg3BQ4uECgUREV9o2IxaQwdkHpXFrm8BGNhvVuaKqrjFkBWuaL9pCEQ
EeCFvVlqkCnWwHxBQrdzIyvNBj3uVfVXRA8cuG3K5AzVh7kh6xd8M107FzjI2h69
gSgeulU5Qgx6RQQ9EGCVPEkE2PRRUYe0ZStnX7kRTUKqAQlpF1XyUDp5/Vxuc4wt
3oAVuVyw9Cyy534XY/LaOr8p2baxLsZpTSKh9tOA+lk3A0WsvuV2kPYEnGo0D0Mr
ZamQdmcSSGeKWr3kdzWSU7GBRZQIUzcgjcWtN0hgJTlBVzkp9faDM/nPQO9H8gXq
+ieRV1bCPSL5/0pPebLRyZfShvBxruMqLp8N8pYAb273MGk3UoU2Q8OzjtR/V6pR
hs6ml7oiQFPPYGmlChw1iSwJnx7oCe/MWRgIif/8vXBFv/262Gd/hnNyvQCufwkV
XDwsZW5WVHQRnxPUkOnrxTPM50uVxDiVM7XRnYdMK+Sgmpag8fkkYK2STKZ41VPN
AQhfuwBkAOY34T5xiQyz/b2allZTGyv4IKEGoggodA0RY2Waj0BHCqwQAu0X4ynE
U1JubBJaT68kPm8947eyl1Pj2PczeKk6d5jWJLFjf28bdmpSO3/dv+SDVNEcOYVZ
7/gPCmaY443UORzcEKMoHEXlFKYolGw/7XtDQ9dfAp8TV9GZL/zbe+WKhVNumsOZ
TjcBfTQcVxBUK0RFhGNGFo/vLj3A3j4ds6IEHttEFo31i0LjDlCRrPMQtfuqLhpI
9MW/H7ktGEGlrKT7+NTLmp94JrfgFxGNcXkC3V2g9AGA6oVlUBFXaHEV+e0wYSit
Ax/KPtkhe3nE1/ewgMgNh8BtcbkQYTOQMSSDuOVMHAYyH/yYQSfSrOKo3nSG/LA2
JQaVX/6Q/2R+kU0t1+OnnLcN3H8PEOBfa81k6FkVjcaZl/bEV6hIPm4eqsT7JiV0
zlZmkv85icWKIAbiK1NywxNmyEQzpZCjj/eGx6ZIJn2TvDFLP5xTlkITOzOHPFqT
xnyJYwUJ5RrJnx3WnFiiiuS9FT7Xa7Gt1XIC8pJP2eDOmZUj0v1LIzxDQDMKVIwl
RDo3uBwKSqIfaXdlIVtGkW3xr7GOHv+zmQUYUSgEA98mF5lBQUKe0qxsQXLEXOL/
B00+xZRPLn68MFXbjdLiI6M0UfpR5vATuGm2QyUTCEXY5COJO07C2T6ZBdzEzMsG
htvlmcTZrp2dhasIBbxMdOqZ/O9gjkwxCgMVIR0driSmG8r+/Ab3poWcNp/fpK/s
KF6XHWtcU1mL8q/eLC42QLCYH5yTMZFoPRe828pfEf0EHUuayMRrkHUfNavtYfxJ
fDz267HoI+0NRSn5C/x81iW22ASrl59L9HPOMxQTxI3+p58bFpZqsb2LBHbt9Bwq
VFQ++jYt9eip53HG+8lGZALYXUs8wGf2wEFqk7GWDkDlmdApvyd6tpJA0vCkK7aM
U+ZvhRTpS0v6SGQB17yPDZTGszHLiA3qq8fMLroIK6ZPrLzQttBErf4lpL7ZT9mA
rj/CzJxe5n9UtFifjksTOvGXG57bAD8kapSO/+s1HEusVaJO0P6v70pTGmIoHCUe
wxy7q15bFpNF6Fp8kuzAIH0JDZA2Z27LX2D0mGuWMGc+ITXqzcQ7BKKwjCJeTHAy
CKYLJj9lFvrTLAWMidBWmMmF9aX/Hitl0Z39eKOCg69rFGT8zvNSFvqapa/ZEo3+
f7wVUMfZHvygjytzalw4fCLmaj7E4DRIJ/nFKGphst85OXJHhs2pO78Yv4Knm3da
Q8btnv0WObMNKfooBuDQDu+bzL4ss3Ic6pUhoEiv8nupWZVSo7NZo/bo3NHZREPD
2aavU9vDXzvjfFxReAOxxDYbfwUv0rjWwNT9FKuxpxsHneVmeZ8UtpUPem4s8V+g
wzB3/fLSG/3rMbB9VZIc/edWGLacrBpjAVSXHIuNd0SGvACji2HMYaVsEXNYI5sl
Jj5/fnnluNvzX6UDT01VCoCapMY0FeuE9id7jN5TpIhYyC/yqQwj6tp2V1N9NnD0
wQVeTQQQ7iPz3IYRzfGa/ibsCo0M2ty8j03e/97+B9L66Y0fBYWF5D/aYK3S0SXu
tccta+nMxzTj0h7CmGUGLdYsyKqiUnsYmiUqLoFXfPfdvoBVINry3wtb32EeInLc
ZeUR9LYRQjaZb8hLAP/pCep9BcTQwsxvB3BXapcabxyyIXaR0pasm/4/aNFT7QGd
8EYN7WicBOSwoC9bwZjBtWusT8MEhpDBldXuD77ndUHQhNUy4WrEIj9+deM2ATUX
Kc8zcc99fsV94AgyAdCPmh4WA/d38NR3mMzwcy9JKy8d0vZpedQ84eFct5aW90Bq
bAO8B3xgjrWnpot4YdE4YZHWJpzkirgdvb2dasz2TDuDpXH7UQOtHHE7GFbBWSRZ
BTdveI4wbwo+QPVnUj4ASXU1kIsrLaLje/x/xB3DAgtdPHxj7D8J6/3RmMKV6NMy
E21q/jKqDmujq95mXH7aLF0HGs7S1rb+50sivid58q59Na4n5ZEIne3anfiNhk7r
nWxJhLf4YwhafnVy164M+N++ZBWfaonqA01UfYENoZ6RJmFpon+4az7iVJBDevKD
O5dT+CfjAGbjYj0n48bSFqZGfYIAoDZyJFsSKUmYz42kXdsdE57nYktipUwRLlVj
fcaVFce16IA/rMSOhNRIbeNShDiYFXMPy/Nr7AXik6+M6k///wEGgGsRdlE2kqpI
YJID9vtG6XB1pWevI54WKPXuAeOxHalucP9IOnd2d602EgCXmyDFB5PGcibKs9Q4
gUpwMJaoRq8bWWEPZHvtJJO2pOGcM+6uOjKCzVBjgFX4hodY0F5/IGBlvem5skBW
TuGiqnRHgvVGrpk2PaUDhWwM0eRgAfjHYhKlxhejBOypVMJDQpvEiVsXwvhXsYKo
wYa30edhabGoe2AaPfI81tmg/sMKluOR/jXEixD+go6SeKI398F9YsjsINOMcHOr
6/4vbgvq4sA6VzKxsy5pAGlPS+49aq8ag+vL+HeUlver7VQlWKFmtB5yuEZ18koW
Xtrb0LujvIJN0z1gwHJT2T3eDNVr0kLOTawc76cgwRywPbmI8vdkjVp55Za/JHSC
xnzCd/1N8bBPZhOgsddj3KjQc0WnbaLjIkox9m8k994pHJaelyh3Zd7VdjX0pMCa
Sjl/huT4cH8amugzIeEpg9C+Oa4ru0XZUQwy4Q8V77cuQPCYXt/TQ2jx6eSi1NCo
+NoaVEdmP3H6AtLoR/2IeCQg8HCJbUa3IpXWgT3Dg+NXQ2PaJLMQHzSKz1K5K+p5
BmS0Qix0NyaCqm3gf4E4dTl2u6lJpCTJ0oYVFI4LKyvncjtI6JCQh04Z4aOc97J9
11F+30sragp5fJS7py89TRq8IOiwTYX+1+rInyZmQRegw1/g74mtYsjfMrCWFvG8
pYK2/0ANr4feUHEcqUzwbWNKIqSG9gcJ6YU+2aOWPWym1E3oNT/07bwoJLk2xxgZ
adATHLvuJeBb6AEUyG62Cc+rr5JK89yiJvHmE8l9X6ISvyaXH0c857MtPbJuzwot
Wzizq7hKggmLWmwApurEhAnswlWJGuQm1d4lKIqC4r1Y+9+tXdfPQF4HGe+djFMz
sTH3TWeJY64zo9BAyTBLQff9QrP3kmnNOVRiIBRmXYNorcLANPLn7VxODmvtL+v1
Cvhl6ku3+3vR4THVhiVt/+U4TI9SumhmUazSNGgQQVyZZ511F+ToGNLHaXI+YIjn
ikqj/yhD4WfeIlRTrODMIaP3NQpBXS2tR1FaTZ4uu3mFFdjfNUmGq4790ULIXFFs
wR0zKRvBkhLwmo0ZKQvNdW7JUQ4fpLbo1Y6PuvdYiz6BszQCDXNsrMYCxaDPTlfg
hvuKTG5PPVs0+tURMlBNpsrDmTha4HyVG26ZVKNnxE41Ddx9uuvIyRCQkgKFQ36U
QFdUWDJhsqz0fvzdvX9AWkdJSnZuLRWAusH+0UJsbQ3utjVX+W63BT1a4EOVDXtM
ZNXs+ojGCj5ne3TZkCOuRN5MV4rZbYyziE223S85NQm9E6PZZz1ilz6eEe+UdQi6
VRc4UMDGKDvwz3z4BYgvV7Hjy5KaNOKOdXLythMakjm2e/iYi/8MS2NZ4/+wBi1A
ICCJl5awII8e6u6vuTCzeiNB1r57FjRnmYYZ0HdJ9oZt9jY6lmFcSxzp+NwfBzJW
4lEulcV3tYNI9y38ec4niVaRAtVa1G4bZNzrgAEvhwNNdSdrftDgI7UBnhXFHA03
AmI7OXipKN1IIWrbDJk2Gw7WGzUVhJ7vqRgkfIF4cx95Fv7f3Erh82/GxSzMmrR2
BMIpzPLPNcTfncg50aHnSrlzGWfHjQqCRG4O/qALpwlyQTMA/0MQqzpyW0M2khxq
AYbkvk+4xFRDZQ7Dtts7y/dDJKtdyFjfbxfiaRqLvKHERKxTJMyQUTKmSsjgrJAZ
b9XHRmZeU2vnIdlmN0DOt6g4NdVHKHWkNuZDlt+GqvunCPBggpOhGeI3NM8jqpy6
yeiEP5ZTc3XtIWgDXa40OD0kVZYkBajvlkweZtFzGKXHlaGtPCUawuQLl7VheK66
bsqPXRnn3DD+xM5k+/P5DAdmrxOj7ZvxugXbFVK/CEu+HQUzpTF23m/Hu39KRfdA
SkU7DIaY+FZDFIYykQxvYUd0f25YPSzyfPKpgIaw57HtFolHuWlYtIPHkx7BwwN0
RojLAU0LUZs7wPmwrso2YHX+GzSakaGGUr6BIaAHbXvVIGRRzMuZF0HTcmz52ncI
gPq255Knppz4F+eDE1yHQGKiZ3CN7+LbQIWBrDSe9VM3eVNLbxB27VVnYEnigiZV
LXx6qJYsvUeYuNsAil/7sK3ySUgSrM7vhFU/FLxfNUszzK5P9ALU3qSR9PVKgfBq
ZqY3Uo7cGfm/K2g1BUawupVqo+sEBNCZHvUrNyluzSS1muP2sgnBguLk0UQ9pZeL
L4zbSTqbqxlS2tfGi7cDh4un/ArhofKjaiVkaSqs3ubXIzCvm66hXu/lhQJRcpd/
sDnVY0F/PC9sj06eik4uUp3CWNVHZ7F7t9uJo3ZH/k/RPrM6DkNOin2UKKypLIu5
+mWYDXBL7Z/XehHtS8/UP3sZtBAqe8MuBUWD6qAXGIyrpIdifw4MQB2NEDxqlPX2
SmWL/hzC4e6xktX83tN2oULI7EjET9V3ywJxFg5IHRZzW7F7wkppkkpEvRBjMs83
WXJWmEiAZwJwR6Hpj6y86mhsmLMfojgg3UslNBAmb6ROkEoDgD48kITErd3X//aF
UzBcCmxXlmCFDkOd0D1rRg/kHSujqcf0vRLpxAntxj+cmNqTppxiheTULA+ZGgMh
yzB0XvOuwmGuKX+74/4gPPgdvCweKKIRVOERDsnAsiNNtjABSqXTiTXGejgnfPCA
dqhlcEdfBsR/nxbre0N3hLRiDK4uE/qKr1iC/6nWw9Veqy5LmtZFmuca3zapLEUI
5s5n1X1gAAQJRA6RDql3O8tpDZB/JL0VHJ9PGMLBP1z4jHGLJ6ls5UeuhxNqyqpC
iXRTIgNOTcKcFF+e4HYEnpFFCAWXRKf23H0FlrxIa0DbyqBmJ2BEAQwtapoMG7p6
yj4heLM/qi87UesnQE2iVsdP1GuPg3EC5MbCSwsu3w4ZbneelUYbEGqC/RjyiqOt
TTUV20dzBnI15lqbfc8tqyn8/pkmHFSKhgYxtOG5d0LDKmxLWfid6UzUr3pfrqga
HLk4Hpyuv18+8WU5uFFpnalg5Km6EAQNYHeCdQad0uNwv9PVEozypIIKSvUdpokY
CXWmwRhPu88cSo301kXBNtAKyTC5KestxUdilWYzS1aL1cnEOOj7oqQHCcp7RZrq
BTs7txl1mFIEGOe3Ks4YoDloUiyIrNzQBzoQoqL8nrRd4DNXaTm2uXO0PslQHeIB
+cGCHoUBYJNufPtmVtKNDZlPUZrhgtoklh2zQ50yGtKXvSozYXgru25aBhlMlPGc
8WGIjyXJzPRMvSQ9Cd4w5ZiKLyFRLph6CBpcFgIDbAfPuuxUj6HEvxfsZGD6mE50
Kw5tnD/1sRVecYFo+xsZ53KHKQKOG18jGTQhWw3n8QE3ZJrsqa3zqQBuQM85oDMO
WT26POTMYbct759SMtoZ0ciPeSIFCvF+4/1oI26hN2lWvDgLn7G9qD+s+Ot8SWMe
EQd+gHoba+noIgg/zKQNA/NCt2bSkG4gSP/M7ixsC1Z5jyqXkV8i0nwraY93nww+
EqMT669O0/jl+f0wLew674z7mIxwvRVMFUt0ybVJlxugmwPvOul/6DjsbtfTmH69
74KV3Vg38PCk+YYj1OdqxAfMmBqvgyNvD+sX5lCoYxgAFKUkam2zqL6LJKGac3Um
jLTkOiSWmS7E3xSSjuhKTZtQjRcNrtVRcMK72fVd5uUflJMk6ujqGShxEzaIOBfp
+LntUpldJrLdFgGI1HmxBuufQ4uvKJrKV15ouIOsY/ikByJzdrdMTTeThwuJlw93
88+veKOjDA+dbpS3lXZsyr91R0m6PGcxgDQKOL7llUMDUvGIh6HOLDB0neI8QMlU
WCw0imo3ftCSSWZYEj3+dWfdWn9uvxLGEzEN2L2NcU3CRFTQqev9fZvIP8wwOGkY
IuH3GBz2KRCSKuqkX0SLK2Jl6ozQS9m39/5qR1FQQxEowQWx5S2oDXJz6JKWMrEJ
naqvQ1/g6iUEjBegakj9JAirRRrGZkVU2fthc4DbF429XtxISvJVTqLkjxQrdXY2
iPEE7DuOsUQxzKdO+0yE8MQM6xakzdsYwr4+qQuPTTSmJnHYWhmhMYCldl49wGT6
7ta1Rlvfr/7ZtFY4jRDmK20yiRAcgYTISzUBzV5r1zT8Xw3om5LhcgQHiM9v9hLI
32tnMZe5MmcqF5y4/PAQG4utgHKYXq8aLX37CaEPbAhGiFLtLBdBn0vdt6RGyyne
LJdnAqN05/nFEG6XT3FyIEgFsDjsBXa15K591eFVyzE54N0P2ylYGjq8t6RFHQX3
4mMd7soGE09KWpew9Ce1gphrau9U6hTRjbvhh8jqcMrA9g30EEo59YeHumpJ7YlO
JODWUOty4bmrcoFiKVJPaGQin778INjnMr9fqicvaBeAFS72sdYwlypA1T0ldUFM
BsFjaFueTslLTFuRT+goS+wGxHzrsmCfC2RBOoLjzoFm0nPEvth8+BBUuT0r4UmQ
r93t83ZntA6P5eIo4S4IqLcqEW9EPUFYGiBdllUsLDQB/CKWzdA0YpZ46g/CuqxS
0eIM1Bm70RYW6589ER6vJZuAIvMjnOSD4LAB6o0m4pGJsV6MBLVqSYD/uD3jij56
q49VJbmY2xYbgEvIvuc54tr4Kle1RIfJFbQNBA1MWUbIm2a7TMEF7mb4sNsRBFiq
muE7RdNVmLxOpaUGndFHecIONr3KvonyiVE26OiNk/nLYYM7n8rag6XRf7dQvrIz
rduQnA+SdGNEdjeGGbhgRer7b82VMkiQ90IBvhDoPztHfXDNFt5JRyqJDyak80MG
iRAM36Y6MMjuByFUmrOXl8pDgHW45g6oz8gV8BfMNYjzePjQrfIOrjBUc0Z4yr+b
E7VByoD84pCzs+e+0ex0dE7Bp7wtWhIRjCijAN5iX397u/0Zxs/FErstziCmTp0y
+QsJQwVDmG0VdFDj1xahWWxEH+DyvYIuwGbJDQ8vfTDMw0knb4vgJo0TyRKuKAMF
oVakon06OWZ2l+WjvM2heEua9iSGXgZyrlsTpkjnrDISbF8eVCOO/1WqVDiEu3kV
2/5xqNLLR/jw9dYzmDctY1BYA9L50fJERD5ogl/PiDacDBpn8zVqYzVx8gpBuV4Y
Bn8DisPJMordwdtawAquFcq57icKDGiZQlLtvugZtIgpNic2Hz96U2u5D+nXtEm1
jhtM2yjgkHZzY0znvVgac3QNBL+LXWfVR2WaBby848Dl+jHtalm1tDhBlTuqWZOl
O1Z4BJ2oyrQGy2NOskQHP0ldBo8HdtZ+F3/tluK06NT+Ot9UEuALhWq4C42cqYFB
FGjwedrqCUVQgojWl3Ppv0USh/YufSbt+9fXu7Zsem1nRMzXR+elEvR17+LaCCLR
8IBbkx4dgcamadC6aKwbNq8LEdoXH0eQXKTpeNul6Fl28wKTRrmDPXg2roezpFWD
omrM8RNoEib6tfj5LdneonHtqr3lJOZZCKx/2+cV7K6DAMQmIGLHWUWQ+PN5svX/
bBwjP/+rky7Af/ish09z/X866etk9inNwbl+gBmkdudkoZRxdd0rktMLzV7uVSKA
3NqJZcAwZK9MrWDvVDJaPRiKZJvWSnn22GYTQrnnrxfXAmEsihCu49mg4N1UGh9d
+EQHlDwSf6asd6Kt1XrQ4Jifmym9RXTU3LVnWquhdFk+g5dUN7G7KuUEc+jdL2+z
By8XGl/CRbzWLFHHEdb8s4wBhL3PL/l+iztppndHV1qnuRWlhyiY8a5z+7adhXX4
ViwRcyhbO1MgYADOO3WncGNfvN0eZOpUC2nWX9dGHTEGWoU6hTColNyXmK73kZtQ
nn9SupxNa/OyNPHDQHzJ6ixnu6NxpOsCNMbQRxvj48nNh1saaccDvgjvo/SvXc9Q
LMCcfaMkQhMrGBh5VkLOFD4uxGetUFzT5brcF2U2Wr/V3TeksrivkiYBOnTIjFq7
80Xh0hZQF87PHCRqZb/tEF/fWBj504opuA5m00LRq9Tg3hJGf0+tSHXmbwNO4AeD
uXzB8fdG3Y3lh56pnXa9U3ZA2F+s/esZ/6klSmMumUIbRrk5erVLdrwAkdEag+O9
9Im+Y7ms0kAbuhX+PqZ93uiTgb2Au6bImJASuvqFAXxNKnETOnHtT+248mOwjoQW
mKLoaXKTOsIiKGyvP6W8Or8r8vCBQXhUMfxdP6kxqTaoaK6GRYUwuCjG4hT3fpDU
+iEHXiBb9nNlRnc5SwiEKmjSW8I/j1rO9JONbZR59g39OBwVxM35IR+8GwiMv/iW
TfkZz8XuT+rZ29CGGLsms8AZ2BH3d1lsqkjGbPQS7MqpbxzIqod1X2J08AhW08CF
RNcq83cT2DNZKRYxBRgRgafzf1Om9KmE4Bctz/4dvdi59Sy9e6/21d5+MRdWvfNE
5OSxwjhUvYKRabkH7myp7ef7coCMAlF3MVB+AgQV6bmY9f5EpeRG5sWuwubCbF3t
hx7exhTuIJr8xMQj7x5XEbMPKVCd8i0mAdySi0QL70sk8y/GkX6cvDktjWT+qoTZ
fNmPal32O16fkCQSfJjP/nMGhJsVnMtZ8MQ/8oIRxZk4ZBPZQ8FDIdgrTvRM18iL
tN+gTKp0WQsi/t1K2shSfoq5cue1gnXt3nMOW7ImuH6A3PAbH8Pw6t6/UGFqJbBH
rJUSsh8StH48oU0+Xvsa0V3PcnNRF1eL9ROg2K38QaJL+nliyny+avzj7MdIkmHn
wceJC7UIAuLnyxtb3ebLW5rHvnLcA+/Pgq1Ix/UhFZodZbbL7xQ9Qwr57CgB82fJ
PcrSInLXQvZqraoide19WXSYA7Bh18cobjN0yIDz1kO5QXguIXhkeePBfpEQU4NP
VjXeJKsqMW0O/1ZxKxN3U8jhip+vPyQ1vbnhPgI4Tb84tjGHhLakmb6QyLjzAgbh
Rgz+KFFsRcCAYgumltFEgWdIFn/abVCpA3KxYtKpr8hDhQc52yHnFuRIPiwUMAeM
Zqm+cpRSmUPGzLD0KDZLES2Oh3xLgxe2W3cDKDHlYW2h5T8L4ht2YH4EdE13MjmG
Nd/iH9SAqgrRVJyuVlitPL69q3xBhEgpGgC5sWzYeqjchffmiFLBRbYjeVmFMeby
H8I+dMtCbFtBROf8uBBjyQMDbNsyGSrizPI8JRX2fwofEH1P/8gzlwvN98tEtMpK
aq9lWmDvEMAFlx/n8lvJrYKRgSWhKBUpsqnO5WlYwkkF7wH6zdPevsF6FiW0Fsn/
04hfgooRvTLn8x5x7a5ylWqp0kTGaCcqYQY7QnG1mkt0/6SNbyT6t+w7Id6ehyuX
im6dzi5nrwRhyDFYgI6WxLhOklw5YTJwjMOL3hYqdAxySjnrQlPlpmsFsW+QJu0W
4BH4VTO+8zghlaRPGYQBqgs8YsdJ4z5C+LOg4PWbcx2mM5pbEAcDBamiS5cLa+1A
87A0j2W2cgKemB0hks11JoSeILv9i+4cp9wu4XUJpDv32++zmOSD/77nJZACnTkp
3jAb9H/PWCeePbXmMrjPoyPO6yW2A0v1FOIcRJ5RaXy5eR0X0I0U9xINfd4Jngxk
W8QCWOBpl6ynNMmf9M/F1X7v1wzNOF8lHSSiioUBFCwbFZiYp2NbJX6yJVD+DPaJ
3+358vpu9R0aI6LQoNxeTEJaKGAsy6F7nqgOzw9S6niEjkD/s7a1IYyrXBqofwZO
ue/dH0PcsUYON/jru+G7CDn2tTsnix3+PofDqc/rzzrJ5sztHfl1MkYe9g0Peu9S
CHozNUQ+CWLOWDFYbrZKwMuIbp66fgyk9C5MBUrZMC4/SrIFCyDx+R/2ZO+QVpM1
CVokGoj81HsMSXMwEaeSt1qe0gvJvEaKr+pn9oWmGp/qE289fPfhk6O98Jpl6bD+
LmbMX//QxgPFd21cDLM01v6uP2ftoksnLrtthACqjjqhsVw+R4CRWNwey5L/nMAr
ojg0u4ddw9XpeBfBvvJQoSCPgxXG08lUYQwi4wpwgQkTTxWBmbChLKiWSK8smQXY
onh9fT/fDXP0k5ZXIp/sCpHqU05+ZfV2bhu527z1G+UQwcLtaKx3LIbyw505UROQ
xF1sjI6DC43RQYgaz60PbW+PZTh3nuPtDtA3hZRqm9UcxO5Z+gfAsPhU2J4S3Ciy
+VllU0vXxAfxOLHxrBXMQwQunYVS2nL37xEufbRYAfl+jV/Irt1dscfpbNPycM65
siC3hHAUA+WO4y06G3thry+jH/zCj0JSQGK3GAqGzy5W2JrPFYvLWfwA42wUfGmm
c2lbMl9gHYHcPfutXuuCmMSWQGbM39fijqJh3p9QC8/4XgH50Rut7DgTSmZV75hP
RzoVUEs4uEE4kGVFQ2+bUY0SD1ocAFMkol3RxHUwjDriqx9oyp7rDAXPA16G4AMF
Dw//NEWfgiau5PxztSZdzm0JmOmxgW/RSsk5Tt1gmvhlXNfzB7q76hjFvvC4hycU
aPtMDKvlHDBwWckzS7zj1ZC6RiQWBYApN65xtWuHmiXdWOn6NVAx1eI0yEmW7smt
oFT2suTvfJCsD3dCWTfr+UC8M7p6clypJXoxoKOCTBVPq255zIvj9FpfI6az6zMb
qEFY3/SkEk53EejeQ8mK85POHw9jrsU4NCjajNeAyzLcTTRE6WQd5Yc18QQiC9ry
ZNwYitTgbGJVUk9DrJAdSqo26Avc6otrb5iw2qn6qBLMTpv6da7d7955yt2+oBWy
gb8vW2Pi8yK4zk1k2sihRoE3jWtyVEGA7hyimt6uOKgANgiHQO4dolUH4Pzy/Q8i
LQDMYOCNXrW+CLrLcQIOy4/qMC8nR2LZJqe4qo/eLJT0DmzfPMNOIY8rKOWRZ7Tc
CXS/BOjOrUNYJIs1xeXYQlNMt5C+WDOZC7LvE9g0XAfRkcX1msLm3Ce4ZzBP6iev
0VmkT+03436r5isYemiT/R8HMPKQ1b5H3g7SN375Iyfs9vlvfb0Z7iQJYQ8OxxTU
mf9qh5efgldoGsYm6phpeD3ubUmixD07WkDo5GHx4ndYoXSmHAeXk0fC6Hvo7pEg
Es5NOhDuxtgimea9gV+57BidlY6qQoxbtI404c76b0TxczhiNzWxq2VExJqvJAdZ
YDBRPEOWCL8pcBHTmK7TMQUB5H9ULyEKsneVlzcMmQKuEBFG3Gsvxdglz02qoHMY
yTtqfHkGLqGG47s7Q7F9OkgrsvqhN/jPhDU4mu3udKO6vZsDisAZ8Aqht/6KXVsa
d3R7C9/Zwglq95ZR8Sg09fpuc6eGCU7gKIYv3FIP2G8in5a7dn/3KJ2uAthyCkhS
Cwq2cpq5bOnRBtwGar41CMvsoZYIVH0M9HALxko79QKjUzBRiXDaOHwi6iLgHBoN
U7r1hlqai3jzxvfCL0w96TUJ0ReAckUkZw1lNxElzR7mY8NAetln4xnHc1Nznwyq
OVtZzZ3LqyR0fR8GId8jfuZJpuGv8mcmE7s7cEwQprN2dvZByyFiczO7mJuNQw+Z
ucYqUOa7PT31bt7xvnuDFD0A8v9Fir17o/nJmESk9BvJ3NPGGtKfpRMrvgcjyf5o
qB1YNQ0vWiek9HIrGKPaE59Hj2HTFCNkdoepu1lUL4ZrZoHWYFmRFrNqmmyn3mc9
4EO1FrFVwrghaLJYIoTWwPxX+ZNW5ORJKPwxZ+3gAM1MF9FgA/Fa7BbCTCjDptMn
zQrWUCvMB1Wwd+J0MJTZyax6OcVyzmQNVGeuzedNiBdlFpUpj81FTZJX9oLk2+fg
R0by6u9wAiVFztuR6hdH5V+wfZQ7UNhX5zjCsOPemO+92iqDp6O38w4k97HMvTFe
FMChiFJUwhHQ4yt3EC8uxI2DgORn0LBJmKJ1wsE0SzV9eqmY5LieEsuuv5bxEW57
FZMxDGnEgL96txzXtg8vXpKykH3nIP2HODBAtKJQRRMDLmckE+JAyybjr2OpBVz/
cOyR/Xufp2HLH+gSHl+0fUUmxW7OGzQMNVFfM5XDMXy2MgNQ5XLSNVTZFg32jQPR
OI7eOGcWL4pXRQBsZpLvsiTl76L54kKwTjgNI3O45GB5m3yCATarBt3QURO8CFZL
8DzEF7oGhCJyD3FJGh8yLqxttHXr8qxhqL4olZap0gYQAPRw+4s+MmBmEJcTrtpt
KavmEAjrj4pxILHUC5QvK4XyeJ1P5mHD6gcJQnbwrspxL8wzX/U4GSNnizW46Njo
3Il1vLK90XqInoKx5TgKP72l0DQTBAqNnoNBxuPmOeqUrwjIa5O4m2YJc+0Tx7VN
GBzeCEbDfet1PssvHfileAGDCvu7BSUB5gZ2bQzgH8larSIpi9/OQN56feU1NjYb
BMC4KQRnqlCbX4/bxLYJpdUvh3SVGGOf47ouCNy0qwAOd2WGh5DSRF6CKMJmEcsW
wz2mi37KileMatvcNTKXbPKqtfuOQkMYkIp79RhQngYNEWTZb756iSqZFEsdgPxd
AswHv6vbJBk7gVyvmH5HTJ50y3r/xRHq0TZbXEpf4ImaNouGjMQs2GTW5ZV82/Fq
ZQDLtDjDMgo8bJwIbQYBlscuIk5AAFYnF4qbcAfDYMJXhmlVyjmqxZEiyApm4gOg
3pH2P/3d3UJrscJ4Km79YNF+lbWjEdrxccVGq+R3gVQSfWD1fDP4qyhwbceU0HEj
u6bYo6J/6RVgJyiHfnaOcvVYmGcadwUQfgDhddvd9yWNW75BTniRuw82IFUQbr0v
HcoKnI41Q4fohX1X2ix8GMRxrSyYZdlLZR9GCH9om77znHLoHPWpbsvvNQ+eTGtY
KFaDvXo6/msvz6+jGJLWtknl6J61GK6M+kL5xUDhnuvGbGPdv+0DyamNLM4zCDNn
bNUFccNKejx5fAGJAHDk8ACzNmYZYJCTQwz6oIDIVQQivSeKpJOaaEG4pkxt2/KU
CyCw2pZUCSWivJTqlp3rjFKWsS3pKnH4O65orcJ4UTXd2bJhR72F1AY7bGdX8n8C
ZGoPyothJAvUI5EoUhKt0Y2HvtN+khQUakfdMXrnUnv5dPEZL12gP2GWM4RL2PQm
6uw9fbhg6mjz4JUXOeSLK7bzLJN9SzEkDR076EUKvQ84kZ/KMbpY3ZpSr43PD4uE
/HxqbreTaoNMWEyiZNxTRpydU2l0pq267Ze3KOHiq754HrGIQlSjN5cnDEwwZczo
OtjC+jqPXv9Y6VjyYI3SfI1TYkF+M7eKJKJLN6aGgHuznZCFSDQ97CVrd0Cue+VZ
/JdJ1ci6yoZXACbYH1V3jsSKYJpTtMTvNGJ/ArXxP60yOfKoHYAooosB4lHZWX/l
f6tkwdnDx5DQFwZBotn7QaMDXB2HQ6nEo+wh+ncRAM7V/V0PVwejBVffN0oJmeZh
xe4IGbJDg0ef3Jzt+7KWKgOh1IeQGMvIJeYqxM9wIhi8N7v9592wTpcfxeeUxq+r
a1e0N9GP6r9hxJ9JWGWyU5tRb29DK9zWcCEZ0ezMFGOQ3lB3CF3nbt7a4NdkSf4z
JoPPh+Z03qE/oFxdpup1uLedFhfdp9Eup+5VyTCQQIPFrKt0dhNIujUGTtMyb1sy
jKHZNgU5TzxwkLVM+7piN3X0TpnYpjSOGSadIYY5yeLbLAAIU8YRjzdK97CXjWK6
BLmQ7uz2Vzsb2IXj9d7uHYZOGt0rRnYu6FD0QhOZxVceN3MInfYlvr4E7OF5kvRJ
JmkU1wRXr/IQTsDl89knBVRBXAs4BuGgX7op3VR+C4yCXJOMPqPkW5cFma4kgWO3
XUcVm8wckcWlmeYs74FUqqILQ21DQQGA23rD4jTO8ZzqMveh4FdwY/Rh6PbbjF/u
8xhiLcgSmDXKm65uMLl61/rakWmaCr/oYiZ5YrdrLGBjE2ODglC5PmmyA3CXjacn
Gu2JH4Xf4LqQfU62TmvGMrGNi8fDlQO/vHp+aCBo2sTygjdW4KKZ6Va5tefEhHNv
Ip40DOtmui2gY9UnZDqX2Mj2S027AOpIVaCO1NUXTLNqXbmS0jFFfWuE1xFeL5nG
HHOZGzHjQzmwcN6+DHtQxGwpX6iWPyfOdn2fkdSJ67SpoMoEGKmEu3Vf8hKrGRz0
UE510SxVQH3OOQQTTi6EWOPDCD1zAyiPrp+K7bQdeMwB3Bsd9yh6juAPuU8K83Hw
bGSGX8XZU0sD7Yy0Nh/yEmVcJUoxlSscCaTdf5Sq48UkIm1b3NdFLaJ9VHmV6T5i
luLtuOfmeyI5VXKBojFgW7kf5KcPL8b38bIRjQkrANA6Tj1U/t8p0yr7uUrjYQFj
S/rxL2VdzQcyAgVpzGxVHhRtFWYeFfstUI8Ac4NMLpQvGxNZudQzaksTk0oy1vQa
S1ndHb2DL6Q4zIE3je0qaHNJq9mN9/HJcVRYgQVhCBAa5qHZiFytG1EitdBLLs4g
WL+pQ/43AoSstRgyabin00uWxMVaOZA1qeOk3EqgF4zqzkCdTTkgm4HrkOiplguD
VIe+dRBFtG0vEgOftg4NgjtEeBgBNjWY5aKT2LxvpItD4eSdGFJ1C4WjnzzzezZx
ACGmbONFHajCyxFqpe9n+Mrc3ml77fJxIGlhOtbZd1larSlhdjU4TsCmrGCenuhn
pyXFy9Ndr2HDWJBEMV5tuZEURqks5MT/M+Qj3gdCbgaME7gBYykybmMBaVTgdAmg
8josMojrCbm2hoRif89QK3UwzpLHxPB6qLWf4pK0dPRcfKHkPxcReHn/RFFaOaIe
PDloIjWEZqs3g5164HWyEJ7WP5DsiF9jfoqrtrZ8a6nxEtdqCBDs63R4PiWtru8J
34u/ufKvRfV1MmCTqnSAofM6LaH+ltNlpQ/WwhkqsO5sbpgmbC8LqbDve3aMAeiD
xJjZTbT6s77pdrTk5tIhkQFlRX/8ov5kimNZcnYbZ7M5/cRRf0MulQrxtGggLrTY
dMKsEhngeopsWEzgn0RRg6LAwTVlAEdxsA6r7/nD7GXoSbuVhFgAYaTZovBqQvhZ
kM2yUBOQ0j0FDxL+bI8yMO0ihAcBU/xk9/ApUecAJo5vpAgsZJX70XRusOlEnhT+
gsaq0VTYdGy4JlG5V73z/xoxTx2oj1Ircuydns5mfAH60lmh30ZDtn3kxkgakJbV
84PttmbYXeqrHWOmcHmTLkYC9R3xNLCsnHclOlPtkTpn1kNc3kjIgvXk9PNaUJ1v
dbff1Ba13wSuCtC6F82YYfTPlRPAYEecblZatml8DVCm9XDKrlR1FBA6rq3ukgRj
1levtuf+XHj3rRWjQ0Eczj96Dtyw0OL7mdaMnK2kTp5GSL7EW+eEsrvUFKuqOvPS
1g3p95ivMDca3k1HNaV9Cj4MTTZtQkJC/RJhRoM6PDotg0IcY9X8Ey8MMFw6Wdtc
FJvGMb6cdyt83+P4cr2nsZYuXpVGkzNLxfKgrkTyu7AGIZdftYFqj7WxYeaKdUah
XGrNnB42uOVDiMXTbshSxzKYp7EOgRU0ds5Qr8z2RkgR34CIoqcJ85Xf8JXf4Ycf
4pcbqJwSnoPyDQhKYqs99JfpzbcyKswqf0LqaJ/oDki/4T+LuBvd1Fkm0S8xQq+p
y8bzrJgEdX2P7Bh9pILWGYxSGWr+hBE9BV7rgln5FYREFKiyGoJp8M4grRwQ0kgL
Q1/jMA9NhMxC599Mo0Y5bpF9YNOEi5rAMroT/jjI0Om+orzKj5cEpeLOrLZP7SNZ
J+er8YmBnYMxJmEP3/MNoJzhjDFMe/rP71zW68b13k5f638qeyDTeqlTyNCnl1ME
XjWJmgckLmMR5tyPzPENTaICT/daUSeHT67rgZg+mnTvWV5T66XhWRsbu9Z/BGvS
WebjTWaqSK2oAJntj/82sbbSspu5dxIaibA/pQ81/CtUtOdyI4othp1D0N5MIw8F
Pvrqj2kmuGI04LhSyCF30X+qhgtYKN2GK7Z835HmSi0Lfem8fDl2ytQGKWTqqqjp
cpqwvORRBTc7D5AiF504Zee7mL6OJ5RGtODTvNEnvfIq+0jWtzUyPW9YTcoH0ge4
H+Tdzhlob0bXBrCWa5oeKw2Cq7xyNkcpgcs8+gW37an6OkrYKzD1PS37F22dqdRr
qJxyOFoN8cv1LK4KqM5N3Szzri7iD/aa6AI+y7lRnfAT8AWpd48zER6FUYqv7PJH
cRQJF+FRyCGAuM+Ib241WBmSVlcxLyxb44yMia8t6GVnuEhXITYUdF/tMPJ7JWGk
flA3CBXQ3uTV5O6GuULiIFE9/jwnWw0ZVLzfZYCV//dfcCKEuv5WpB8gFy5y6k2L
rH9+kZn/dMNfIl/v40GsYQPekk+cPubDq2nCnIzvw1ZSy0jOfjxxgjzx9mLgS96k
g6uExoarTTNK3ekHxoF9U9A+6hFw7kTu4RkMjIskQJcCJ4yOnOPPejatIgYcIfR1
H8hcImU+BKYvfSeaQf1JlO7+lcXgueNjbiWlnX0CjCe2yVTC+Tjx1zAlCkCpHRCc
7yZjaa+tgXwry02aZNzB8uDGsc//CGa3znclrL8AZrxw680gYV14onkEOW6JDhKl
rYq/otZWGLH62XgoqTW268OCOlJXrqB4ZJxXNCh8p/+h+GxNGiiKp4bRjVVyqS4K
Js68dMp78omDmZpsO3Htblr5NVk0g8uT/sNJZ33DP0oQtKdjwYNQC2qTjuiZzfCF
kj6Nd5WQAPhncwQZ7tvRr65tB97WmWU4iKm0pJmGOvTIODjeZesymJKC5EiPo2Xl
sdw2X22a/vn88A4lNc2hc3OKl90qvDovvKy3vMx0b4oFBFWM7MxRBVLNheX1Cb6o
UyhVOz1RfFgHa/X+vT4pis0IMmG3qL3z0NYBIuvHysoDxSCfMvNr+q0vkTX8B3zC
m/3j2QjcmuhcX+k9rpybziFj/gtoWw3LcSME+FWgB3VAkLdi4C7qkxwd1ZaUytDL
3GFlgLG616aJ137Au6bWSrZKF22yEB1P6WT0Ng5ISrq9IHUOvkKsKcbad7nnjwh6
hYdveXrSBP1ktlbcbX8tF1RD9DTBL+nqQtbUUQ+24TufwC8MJlb3g34MfMPi6I6N
quzvNaTxcqXl9JTmhcU9LsSgnckKrKoB2R75/Icx56Zf1luWhaoveajZg8zAhgvY
3moX20ScOB+IgV2GYYRkZ6c3lYw292pTwO/Fag2NCbzRbOWIzHXvRsgRvSJsmNmy
K3R28Gw1er3ZGxHIC263dsY/R6c8Sa7ww0JSxiBGFV8rv8dv+u2mk24Fergromnl
7w9tVyz1tslAvw9rbDr6P3cYz6mEn2luR9gShdjSigtxp0O7VR7TNBrvKKcGQHBq
Du/VIMGyWWmSAP/mjbTDHlOXHIhUM6cqNvd6XbAsv6+dbIoUKQRB77nMBXZYsVRB
KUs4vkPrQd74qbf9TF4dYz3+5wI+UN+FnoYCyBtgRELfEPcxATn5yWbNUk33YNVh
SdTVN8HCcon5emU3k0abh09CBKccGX23N6dJ//gt0/NxLK5RiuehZpIH9Xo85oqz
GLnn0rsQTNVrXMniysY5uQu17bT+3RbURJe/Tb4d6k/Z0EVdbf5ghKshmc6aEcNs
cPjsCYNSo8xCWVOHSfzhAQvYK3AhnCR+znxNCJ/TrxkbHOyLQM7oe77EUnuqqzDz
/wnp4HtYy3AzQUbO+9nnqtIBhhpFqC23JTABHy05N1LLwh5AeGXX80G2+jeelc9f
7W/7baogVS1jn65PwNCSzyGJndfgdFnnhGatVBYGQksexKHPfiKortzu7VBps3Xg
JXgJp5QbalXC/NZRqan5iTxLeM5Xq1WCc4+brAZ3v1bDs9nwt/1Ve1qBN0GzD2ri
B828lH71k0leUbGQk0QINMm3ZMvGeYnmPWCD2Z20V6XtwiYsmXnrLwPcL4lPnj5R
oD19rmmKTo1iySusK0xo5KMne38vZ3EqCCorKYVbuv8ZtEw8mPs7c8v6SnvHPytn
T1ZZAQfYO6LDahelpRkf7e3pRDU8CXx0XBXT3N8Jg1rVlJSjjwyQgBheTNM0llcx
F/5mm8cc8AJHMIxLxGx9T9kTrqYDGZy1j4B2gUUmtcg9ZIJzC9fJrPSC0o1AXPOT
bdWcv0ehXPRBEFXP8L8gz6xvqbdOHqG9FNAIdoO38NlOB4FmDe6EhNGIbm3XqSb8
FxPohT2kKuTB2u/ekgUG52U5JBxtoT5oZWyEnmzQtLqxDN69tbkRoLDfIQYJgTTw
IKgmrari0hZq/Ff4p+x3bwLTbjdh+IRwtW9kWEDKXs20VyaVNSJ9eQgm1JCARtE1
1uPj1osBH+wcK45AgSKaLIm1nfl2bohwYoG3jJEgy7xWlpIO2zPjpczhF960dIZb
h4vxPbdVUFZeeWvExd99s6CfoDw8DAioZ5nXN103eLfkD3VsmoktqryLlSO6lo1J
b6po1kDt8y9c5wBinNQOYGQsOkPAOwtYzZPScy1CkOgComyhDQSFfV3YXy+U8Rjz
QMNqA8IA4JrV/ptPPnRGRP87hsrfdGnAqlt8f10qpbN2WTrIpp+REm7HGyGIkeZk
1gRX2f15p/iWmwimHwjHLPRGC09X8K/rYf5jOAhLe/byUtVDACtmmIYwllykaWpp
V0dW1UE5h6DAPDrMPPixrg1GQ7NsW45ctB+oQqK3IPGIV7xJw7/yW8CDmg3vK6gV
IMXTIolf6Xi497xMG5ZlYyJEaFQjWhjwh8VqsldEb9ouNuP+jU1HGgrNX/j+nk8k
xJUha1ki6a65HBYNiBMxlE/Fx5tS9fna72MDpDprRbMacq3yVX0alfaOvnCa72NV
++iqqgZekAg9LxNgshjtLj9+7HdFJypMn1n2WHzwnX/GZYNfzTlHSxdDxaw/71Gn
XG1qkrA++SsY/D5lFZqgxJSAIqPpxPENsxBtSGkJ/YpaVD5RY4yTCehfWEfZG4RP
BiYsTsSMHn2V99CxWjJViY99o6U+nF0LkmXjO/WW3UlD94C5QZpQSREEEji6Kti3
7vH60feqfQBzNdaE8blV4dkAAgIpT22x4juOhOygwGYUMgc3Ns2qQSlWbvhMBHCC
H1/dFaUzxyYjFbI9QG6lnP6G5bH5NIdluoA19ZKyFKloNExYq1/mJgNe7a9n8MTL
thT2g5VGA8KfFPqiNSczYdV74RElFxpNyRXSLhIItjFWDjYdu4ZxCyRgo4NUZ0bw
T7duG87D9esxuuZR9xczg1hoT1ICwJcO2Ng1Slsji2ombZJKgODe9t8GRHrhPJeA
ZYUkj1buDv54G6dYlqavDeCBwnCULaP8Hctm3OAroLr6+PkC+MACuylywFTXkSy4
xX1qz1E5QQIBwCU7+dyJEln4xcUORImqqI3BhMBSG2CuoqH5spZ71WHiMe3e1u7J
mmMmQMPPoP5ccm3yy8BKcQ/Kzh3LQ2Myn6rQZMtH4tbHODn3Kbk3cnlNpOjrveCg
FtIFs0ecfPRccnbnOtauv1wbdZ1HpDgEwAGbsI6dasNKTFjjdmFU/S672wb3F2i+
fCoGbRP70OyaRokTwQQnu6RNS4IUBotd9Q6OsG57qVtAjGNbC7veKjuqUKRXr9GC
/QCx4FLTvEEwH710UL9rMtj4nqTirK/tKWxbi6ePnRuQFq6D2XNEzmMBoARZBqRD
hahaqkBORSXNdK3C53vNIc7C5oBjhbGlcIEqK5VIUhMP7G5Dj3hjf0WyOCaALW9p
QQ9NMhJfT+Ivx1jPRM/Ha6DFSklihP9IC2sus+Ex6r5kynwgA2CEertIFJ1+R5n4
+JCH3Q3JmBs7F6cYkj6BNyWiByIzimuewlK7hTLF57/uA2GWepNa+M95/7UfkbYM
n2sW+Z63S2pCHpfgzdY9sfZCGWkWD5d0jPcqI1jdtjrAo4vUY+Wt8V5+NwgGg2HB
TW/CPS9n6//1aUfeXgkiHbi7eAelP7fNKgDIyHQztg3dbQavtatstp+FcQ/Tt7r4
tcl8ajXMy0QNg4rrR76ZKO9O+UomCXUNywYFsnosODYAckuDMrdTOTgH0TZVimU2
XFgzuiPRpty+rAygbHBFE2Jn5tUcu48slIra/TKcJkginM5kAcg7HMnkfDwPbw92
OedQmmV10IzYI7AIDKQrvoVLoms3fzilsT7/ykjDJeEmdzYhcJNJNXnJ5cFPN/27
rGv2RQRvBKyyZ5ZwkhTWEXt+vMrOQZzuBmPeJjFrgLF7tNLqfhe6E1FaTVQAmAkL
APuopRs6LLOUPP6DmT7Ll6h4IzFV0ja9If6WgHHd7oSL1nRW95XgdNQD64O6F9A+
YxDNUlSACsZrWCY+yUI/dpeb7xw+bvlSsgZK8YAGstrhhMhNZX/PZrWau527J2Ai
u1ZuWkTZ/hRNT0DAzC0isMqJ7KvZNGGJx86WsI9uJXPkUVr79omEoxF6zXq/n7yX
O5w4M5IYij1o0JiIGFruKptfbmkq/jhe7OrVzWaJPoaMACiuGcv6ydvqvRJPlFE4
aElHvsVDj5X8fMluDLzcD1kdqAbO/uEw16GFNWX+ja9/yTykvVksmPVyzWqUklXf
ocPLtJB7WD1/8z7aqdq6FGWUcSPk0JZAyI4xJL4SX0p/1TFgTEDBn4qOkgYn56HB
C90dibnqIXgfluJrfWRt5R5sDiFF75SCpZA6mjcJ8LNVb+bH6zCS0zU+LMFkJL/O
FZZSk9YKugHa5n6T427/WqrlAIBEG53ahQFgSnchLS78Ht1uv5VcCvkf1Nt6yP9I
cqSX1FCkZ3CNq7zOhzizF+vlqneuyFnnig+r3e5CUW5b7vQFsxNsyaqLFhNc2jLQ
7fgYKBph6jKsCzARV5zhUagmQDtSnR59+v10/Y9XwUvIdOZkykcZqd27oksLEho/
wEYMIqtgnevflI46LZO/Zk2jBseBlBjrNGv9dP7HZS5UKhMr1xfARD5pfmsCknkK
ecPbkSEHOyrxQB5YQTUMOVQA08TXB206bd+/ROS2YPbqyshBTB8xb5oJ7xhENsfp
twR11qLLTigHQEnMthcSmxsEm6fbEJ0MivOOKJa/sZziXQwJpaDaIe1Hrux0FaQ+
0ttMkUhHg7yR1QmXIpYYH/XG9uCEBtVVEaBdbUmqgtyKmgXbgVaAylvvJ6P7CmDD
dlxaE9NHl2gFTtXpOb8ZIuy50DJiXdDO6zsu9Z3UjHdHzchBQrdRUf4xkDmxYQzx
SqqH8lboynOVnP6xS5Jny3YKGk2SGywNzyRNOKNMdhH+Z3zu3syA0YCZFgFiqvTk
gu5lb3+JVXVh9zJkMojo8mDunbRqHzUDDtCu3UwkwrDqkS4DM8YVPchleJ15nQwe
KquGlE906umIu1QxY44x2PbtNTEUv9cYjYhDuX8G/jdHctjHCvZMxL5auW3Mntrh
nFX96LjY5ohX7fUT5x8mzxACrvDV2Yw2YJEw4buVThSA1ywnaMBnOqUyOzk1W8Cz
Md2Y5Txe/NeKVK6AJEGZGqtX9IQ/zEQ6aVAn8OP2hJ2XfVuLNtlI+ftvPAWDd9+j
OEoVScfHKoh8dframa4J1M1sOMfPzCrVFsiqcMIgawf658U+P8tVIFd9yp5VGULy
xqSxNgcqyT8HsRDB3nvRUvtR3mpxz93FDXE7KI2OEwdhXZ487CLfsJ8BYieTpZpC
9lEHnP4irbr1L03ML80YJ8/YpFZMTHO71SPVDvnDfLSnBSs1N6Jz26avRLRT+pf6
eohoaKrxf40hpyV9qEP7larYLFqlbwwvUj7gt+s8GJBL5QWIiiXZ6Wp0wQY/hHFl
3qJvSHOtYnSIT4SUHpPWkweYqjl8eLp5racFKyOLMSZmg7JhkyLV2XgYv1Ettn2e
VzoD94/w71Sv12sDeI87WKrcHX+YNjfpUjE7OVaQqGqdmIPJCpQFDMWY/KKZsLQN
78jzfCvhQlDAz3oFPQFy3AycE8Oodmv9BAN3eHqe+fq78HnKYSk52lA4h38FJDY1
nkauF+vTOXQmJ2xFLMvrYxUE1aU/TdYvlzV0RvwJFtfrk04yhn1xaBfh3KFFuLC6
297BOdth5Zb+plMh0x30F4vmXWAvwDl238MNdyeSFRTHMda/cIEi4FQj8yDCnZn/
R+DF7UY5vLem7kRKBbyEpUZIvN+b7uMd12CNgBlqDuKPA+3/+K/p/mL3qw9ohaVY
hVVCn/l1poKdFMOopc3r6ePormTRsvPxbucJjG4awWGKeAEYFrfhP3PuWS0JYAI8
tUMe26XQJQF14rCKN2zsg7AJz+SY5WZ0e8W0wNGrpctgMBaROh451OmyiAbdSQeE
2COnIaoaHcKZry2eRdUs4C0FKzuhmx4CDWJdNLc8yEl4KWYEAFzJu1bPqbKk25h0
pyfCYRZ8VSn907ocb/88o/Utwt8OJHoZZ/gWWR1AP+wzFkDR/959ODG4dfIiEbUx
2Y/4AAIQ2UF8P3dYa4CF8OouS/U72LgSADY/JymICLP8PczRub4f3VTW4uu2Ojr9
e47wvRdj/ALwl39+ZXWEslGIRbbOsT8Jpyo3Oftg19CCKx7MMyABdvtaNE3OzMsw
Jbb3TR1un8pj+sfM2zJp+gaCpKKJtZeLjpmM6yrlFrxeNVcweYQApZqNB5z5W/n+
uMEiArNEtCRwj+BjwHv0qgARFuDj33dY1D2+cVVB3lFYHwsVsygXEDwB5a5CheG2
F9gI81013NxvQQVl4R8Mq120+5AZJ6oio1paBPVXw8ixHx3ykjTt4kunSth7Riaq
yfP/j0bP72GcbHOS1Uf0YalC7fl6NLGd/EU+lpwSn2Xd4D6oYlVlXCZXSYALXPG9
3a4glVc9v/1DubSa7eK5+9iB4fbnG5ZddlcwmI4XsHRKu+Knovrq6H3jIXqly8w0
rzVMfujVSkDCPKmdaSPPpUkSX/ggKquI2V8wBr/aOjb9gC9caWwU4YydV1tejuJ3
kL+CFzahEdLmNEtOVxeNc3OtttwxsgJMH/IxqzVb5EKNBuS0OrSfsDXpcHMyt9SW
m/reJ0WHc/jJoZlneDJ940T0eum+zGTfWcWzLoUyKutEa6MH8nvltMCnSwRPQeC1
yhS9YAElEb4wxUZm55w0lEeTiWF/ncZFRhx4c0V7Zir/oS5TlzIUonLlceCOLhVw
EnAL/loQyItEs3DbVi9bs4ygN6ytp6BvR3J4y0OzTG/+t6bKUhRog7GCMEv2VUYm
PD/Sju0UUV7vus/BuJRrK+Woa0cQnZKpU+nOBiY1zubZgO8H4ccqrNvk1AC3CRPA
oAwzU/Zlow1dPxHOMyidcBVvDH1htKFjJNnQx8UeZ624Q3Ghbyu2bYSpLWdlnTAD
gZ/H3u9oYiyXUB0N+0fvwk2U1tF8ysi/BimWwG5LhuGIO3esqJorGoe21LKQjfOZ
AhyELLCYEiEUBMgfXCgTEe+Ym2kxrI6I8sCDdqcWszsGnBd8nBbziCpFNg47eiAM
Z98ea/wYgm2d/Ap41IO3oHgEqc2EEHc+BLrD3bk4Syg/GXRDJ1d0Yl/rG7MBi3us
jm7E4KQRM3eKuohPBL+ayPvCS6lXb2Q1+/cAwnn1FH3DivjqU8vtC870oiQ55Uxs
imaRD9ctmJO5vbpWEs/qglev893yQnsOK7dQRPCUkMBhVNlzBWZEoVrAAPbDRcmb
znVPLAvS1a6fdxN3uSi8I41/58e6vklg443etkabIDQ5PR/WQPrGaUAb1VXcaShr
iP/Z/p5wSUZ0hmcdYsg699hlR84KxMlUlNFT/6yW1G3AwF9TTWTqxxRwbRlJ6pCh
vT41dlkc3J4JtmnPTyBi9fliC9OCXD2YxPl0GfYhydlLhi9Feih3qFcPpPkEzl8n
eEhSVf6SCNhgccoV8LIknLGSey3+fDEX7vY6ms74mbeOvkPsTtmGbviUaECwNoJy
tk+b2Ykg+51SUna8g3X8TFo/iQ3QvOXYvjHphscgRdUmnrk228Kz5fHwqlSE6YsW
+na6c4qS5uJxY+1YJCLs0CTZO8rnwc+f7IhwiNFpGXaOZ+TCKkA44ANiAGv/WMGv
7cbByl0WgNXxvT1luTONjQLII7ZG8DZ3TrjcbqZn4ArUu1lWB/bx7fBrMgZ9rGql
UYpyw2Ov1sQ7/ShyleR1HUwfXk5dlLjPg0OpYvFC/AZpnnuCb0q2EM0acyD3hbGZ
RWZabRrdnn8DOca1NsfmkTwja75ZvdhH5n5qgTEHNiJAY8fmXHA1HPBFA13gEBIk
wR6+gV9uxNyn/mkS3/ZXDjCehbZTUT/B4E2FoA5RPO/0y+5wH0WCdxRci+CN5mdb
MDc/y8xiaZs5plb0krA+JCtb01diHUhTtIDgjTn/dDCouMwYupp9XMQr+Ca1Zw66
m7mygKpxjCPz5br+9jpttG9r1xVioopEEdHNs5FbdOnJ2lFQCYPW+WRCiERPdiNB
+++m76TmwNuw6a7uZ+a5HZzGwGmsbBnRRBmOwnzMhzGl5AxMb6SbM0Fi7WQHx0gF
B0/tWRyQey7VsUkEkpJpGauQGq6j5/sww8d5Y5ASPrGU0XcgQPcjWQ2eNBo+bBax
0leBmBDrvmA1NzjjwEkwsDymoPSQtZz6nivgj/22pTBUoml718qMu1sjFMVniky3
UCIJTs9aApKTMg6UqUqh9uPSRY9+EIkKEyvGRrRlzgzPBhIqddrYrti40JzEkVpR
3DwwK2uwMsTURt9pDqx7Q6Uj1TV9Q31iI4jRdaPoJeg+fqKwDQbqibGfU/weZGUI
1Fd7KwpFiYDrpgrVh7vuAE2dBOKsOhfbgAIRLBcpSZj1R6wufYyx/51LgGy2oRbm
+9qq6oHaBtEX20DiadckkYO6CDo9HEUdr5+q5Mu2C3nESJaTpe2HW0lxvOn8/ebx
ARbVFiDgroHAswtcDwPLpe4ZKYhfvyPuyq0HnHuOpVIdEjcppd1hfxCLWJqS9K6H
Q2LTDVGqHXwkVO7nELMMjq3kg5OCWTz3jzjeJu0DeKn0dx163t1qEe3AMNSxxBXK
89wYWdExvki3l0gUI/pCD7/uufIvKBuboGvzE4vIQAuxghaNDPS2RD41vDkfrH7T
bpBHXmXVTJYSosidO1QVPgyQf8iNXXrD6oH13j/e/vUOOoOmiNZtP611KBwfdCye
SijERcOSe3AOrMU7MhtJT9JuF4TwWjBA5zkQYKdlF49dFl2M2baRFyZfsCECI7Wy
Pe26vK4H3lZHLfiABrNHIWIwL0JImC2o+2894kwZQ4g9sjhH7wzzdjjrtKBidkrE
/qid1GUHRHdLp7r8TYVmfYohy69brvntvUUQdEmizo3RtPw5k0IdlxEWe/OOJuJ5
QyE/n+U2h0UC28/GTDAwinpw6EnlFFitz3fK1bNhIiFKfCCaUqBHVm6USEoqae71
gDbztnVO/OcH4oFqK2OXUnwekMsxijig3I5Bw7PiIctfT9wkye29knK8iYPFay+K
iFArdNL82AFnegI1AFSLqYudbEXLm2JYFmHpqQaM9DyJQZs407d1k8bVCtgfmz7n
SQr7HejSSqypIICUGpcYoYIXGvvdyD1WJAu1NGgR0NOQMbRKx0Y+3MRuzJVddVHX
SHYiy3tjLOkxthpC75tshhWImqtvaudMuUkdSxpEaCAFRpPxdAMwXTaiEI1ojfat
ou6ONNjciRj9jqCrBuiZSEsbKkWYtJu4eI6Lw2niHk0MO/XOYrw3Ms+TetwWQ0ZF
elme/qgN+BwqKjDCMH8/aHQRjnH2uUjpEtTjPZ+2VWzVN85hPH/KtdH3kXwkfz0B
ATdXL5erCwDFswsRlv0Tj37E+jF6t27euwDMxH7Mfw4Sde6jHehyCzGrk4ns5ENt
dxuskdU3stZ9rmr8W+5BxFmFMov8Ilpp8aEZackDXk2LW/VmUYYxb3YNdbQiXV9c
Mni6Q/tHSN7E2+hDAPUv2IAY0FJ/DYwX9+TcNMlpf8sg8FfcNl2PpiLeXDO4HEl2
bjRPPtEvJ8sj6ScUOfkdxBXer8TuNvWa0nlumTyJNX+rOP3LT5Wu3Adlz0dkFDK3
N9+eZgWw9z+kEtBSX7soudJIJSp93MlctU9rrUJuQY6+ZjzIX4ie9E7aIOmNCVgC
j9Wxvl2eFdTsPSorUuUl4pk2S85V1jPxhCsQJi6vYdKU6kWAeZCciS5Ks2FqE5RH
5KacdrxpRCLgUZnNy8Xk1WSrlv81bmrUEe1xcSTNYTZpEUr+1fivnOonElsC3bPz
mMm/0ITIDQZ91cu9aA3NtaaH/WAIMJUeVOUfAP9rL6/9VdNN5uYI9RmZ8ZewKamp
g4RpLT4C0rGxch/0kw8/r6mWXYjSubdJimTdQ9cwYCJRyvizvB4nLMOK4D6K4Xhu
bwEUaRFJ50/P0U5SyergSoZLVX+OfWg/En0kDrss0CvntJep0Jx8jJU7aYGgQ0FJ
d2Sq+yatohmVcrBn1zheqQaFk3wKI1e62F18O4sV971rPd+hNCFUTmHY/iFiIZlB
S5D/UHJ3+QmvQDTxIKGTUf4DzDFpx2FZFQVMifuoX94t3KXAMywbxz2kCx+Mr9AK
xxadGu33QSHJyreaETZzBhzBxJSXI3CSdM9HNb3YIy3K/7S+CBsUS/XIAxxXBwUm
PHNM9QUhFUhoAwnVRvLrPlFP+BS+FFyVly8f8G1cto7/oX61rcRrTsit5NPLsIiC
TtW6xxyLaJ7PTANfF+MPQcwZpKTbWH0sbXDQJpeslbZrH/2CakJ/nYo4sX6TWQKh
MXQQy4s3wFzUww0N4jAQxc9SkA+XbgtPYRXsC9mzd0+A3PWsbivEjiQrLTmV6haf
yizOzpBp/Am9rVqyEkaobTPYNDJGdDKe5Ko0rezGKWSCi6ePU6BoGRhku+Xlm+Df
HY/TIZyx5Hv6dNt3dMzY+3CGnLai3EO5DFLym2eUZ9NdGCNVXwYfs0Let8sL/UQ/
3tR98plAURaEdydg1932Yh0ivtWq6geMNbxc3ZLpbdcBQelB4MYwkejKjq0mm5HU
OAVnyeoiGP5u65iETdoHefeG7kzeTL6s83r1BGqs8Omc/OS3DgTOeUgnPR9HXCLX
KaLIxrgXw/Fe0bljOhmvrqx08mBvzIGpkAyJAF2RSwzeoYZYZs5/3/uAhCj7HYxl
bygqiWs7DcYaX45uCwZtM0xGkUP2P8P5tPoapub1XVoWWZg7eOyqF2OXd2z6dw0V
l7JKoJSE0AAlw0gVZ5lr2x0Tu6A0R/ry83JBFjxzTCmyoRztkcOSi9PBBH0jUOfy
TN0VZBtpH1diin5mXMZQJ3wRJFXqwrOZHMn1ex2Qk+LHqHA+/LIla5wnXAduES66
0undIB3qkp3rgXbwkx9bR8W2O2qHuqk5UhaMDK89wjOJEm3Ia1WvmEF/UwD917JV
JI9J770knQEAV6RWgVTpAu5OG4bTfSX33QPFYNnCtsCe7bqzgAUl9NvSSvuaRCt5
6m+rBiuuy7wBYyFgpv826kNBgmc2GQ0uBqDQYOjHUpQq1R/6I0oqBzZ2kW2308pq
Dazd5d6vu0CEhtz8dolmFlkYs4NMjd9fxAAdwc2oQML/Vo9UKYiUjtv3qHVoXzln
h5LvMjHTQThowazW3gUlqDp26qLhzWrWLaJTt2bixwfwfmxz5chvHyFAHltR8bJw
sqPlg3yqIKkLOTUSeVVltdalaiA4ZbPMi7xx6V3BWhMPXKjYLY8223rxgRJSVxow
fw1GIToeSy23SMxTTipPkiYEumxmUYqinOqZAcJ/U79q2sL1ZwWhNuB6L4zlNJmq
Aw79fBRBjKtiTG9MNOUuqmAMeCLF5+fH2/djSlnhmspbajntwnp21/JMUAmNmUzw
ZA8H/FjEUES3ZXH8JNDgHfXLO00vcqKYpPwGXe7B55m0LftKijkMkUvyZ6tvp2yf
Y0n6e1CHt0aCxtTLjrypuPxuQvx0v+bACh/YNBOAEUD+M2yytvCrLXJQlun6P8S1
EsjOg67hO4HGuyy9J3fKtSo4FWQaXvKjZ2ICnGqdR9fEbfkaG9a5tdcC7phsR0Qp
ByqBrDDRBE1Z5RkSJbUVylbbnt4GAK1z0fB7ptxsa2REfMp0eW2Z1H3t4pDCqLqY
EtIgy2i/jWqtUvsJVLfMrp7m9S1YS08J74Jrr2EyhsLzgxSrDIRpInsri7rBwIZC
4BictaAHwDeOUNECNTrWj0x0SAJSJ1xTnFrUrK6AQ6qPk8v7lOR8S0bigXc9iCdv
utt2MnyBAgxt80guyvJjcXLJgs7rzO8xM3ojPW4Ajmr6y8W0hd2baORPwZ/GY+U9
NkNDAQHcb9pBCW6MhemSK7KYOOzfV/J/yZk9WNlrVQZrCDk6gB9u2m63x2Huj+tz
XiQmYZCRVnP9lvhfDLLWENAMvAiLkBBWKWjhK9x5TcuDdLnrsX52goAIsyR8ygV1
dC+CoRYJf9alzQvmsBzY5iqvd0VzNP89moa4btgOxDkzp3CH+HauEH+Q0vRbq5+4
LSQarcCMPCM/0HXlGF08omNiao99FwgVE39oRw3vkCA/CGgqk6Aqtm9LTXdR+QsS
cRKuqSGvcTeEIlqwxsCdkIv2T/juDcRp6szf0CoDdarZr9dwX6H5kwHaVwQOwahY
kEl4SdjQ3AANJIJ5DRjm9r7lFpPz3MkUb50nwkeVLuuEr+hMLgDabx94RBjUhmju
XKzoVQN6+F3hwulyCFV/EzMMwts2ys3GoYHKC8NrGJYMQ5UNVfe9H2kYWiliuOHO
YmnSxLqEs09OEGQLcO0Awf0RE0ZKfSCHdRZ3+R3ycxrceBA6nvnRWvSxdwG0ch1f
+1a9vIq5YwUIDzMgptiggRJdMjFIKiqLYsUBOokLhR8vmtn/gkWIU38bkOri0pym
t+w1ve5DU0sh7KwIm+JgbOobOrY9/y2H/oVs1yRby7Q4FWgfvDSHTv82L0RxiybX
g6Scp3ScOrsDf1G6bJsd2IGGvLyLUNanNjFJ3vsOxkXYD3jK0YXpVIzb9X/mqNBu
wrNl4SvGYewQz3u44T3W4TYzM2CItlIxq4rYkE9vTbjEfQry7WXt1VU7JSSwX93F
P+QL9AiN3QXwghCFPjeScfJ4TM8OIxoJRs6FgRmsaALDitf+L8XWPOLqW31RcgVG
WmErREZpLbsxdMPtMZJ1ENYtG7VEwywLy3v77/iyiDgx5RBRrZoNhhByGScrrb4F
MMp3lzSvicAvZ1sZbPqrPl6JPgkkSkSXjtjHsGsrafEwNX91C+t/thowQXH50Wmn
IB/dpjmyMp7UVHKcyQYFGtgZAyE9q7GlNyPGTnF0mD2ejODCpsdUbCzfz7cVe5F7
Ycvn6h+gjXouG+If0CzyPHcTb/QKpLH/rRjKVws1STC8MLz4JBMtwA8DT0vAkPYh
Bvn+WnT7XfxIKBHPKXcTwzVslfcVSWxmXrfJSBgLnhCwY57oCCrumtKr7la9cebM
Vztf3bc0gQwbbiXygS91yJC+O3VEGxwKGIksw3YG0Rpz/titW+CpLROrjOs/FuHx
6xfcEd+7aq70R3wo9nXycYOfpdWHorb7/8skOZ1aQopSrIIRbuFJDTxOJVrRm+RS
kOPb9dGglJMlC1/Tqp+lXQ156PpY8DAPIoxHzn/4Z2hFReZG8UtFrJSQIWk4kSpz
6VDie1pu/O6WSC44ZJk7pHuD0OJVFjcmyt/LL4/HIFkX7feWwmR6K9evQZ8mLq9g
trrgeicqc9ka0+akkiyISKIv+sXAMem4pgHpiWjC/Pzqi80ZmQfSgxjrdtPHVJZG
jkpEdpyhHPnbwuhtMxp+tm69/DXfnsn+KVmyZm4lbxlix0AmiJxrfokxn8h2SGxT
5pcrxfjFR6oHswUeulodDAmf9ldHp6nksEaY6hpmwJD4rLQSlT1ERj85Y+Y1BP2b
7XHGoW2bJLVzdyhhnHRxwckeAyP0f3t8zGvlAzJ9o/IUY9QXtL8UZEgH5Y/oCHPv
x9oXgZM4kULeqEnhLasJzj2C46/hrdmok8lTWF6oOHCssdUl7TJuQWpYVyILfTil
eWZPnWo0kQoMMB4c8ZTPV2Bs3Y+T4iNZ4P7NLwesD9Iis6CpBJSQvh9ELsHrTt8b
7jUctvCG2mTlldqcUsheOMMz/TLaLPJYgw0MzEovOx5x8Va/nelaG+yFjN82dOTk
PvXIMp/PsgJ2G59L0G/vQ/oZ4emdhS0wyr0N85lGnQUWFKx3GGImeVTo3i1mQnG4
qQx3qiERSIR0Kt7j1DxZnuoIjp/VZZGg717mFXSLeVEGW78VoF8CkCFJnGxg4Wup
cGlKvKBE8OWJjnCnmOV5JOSQBx6dmE42c3Z2lg9zw/l2toMHAAwfYj+6Dn4f2zb0
bi5sVmt4+FMoyN7iLE2LCowqVe4bgrf2nKfhsQw9CmF8lx9tn9pctGWicWJHG4NA
fwjlhGtBLEGF2dLvY3VJMSHPLOQDjtr5gHPbMnOsrGtQqLKZyrpQQvuAe3HCkBYC
SPD8fMn+PEyq9FmAN2V/4ltlzlQMgozqZw7ILgrpCDq2xWHLL2+UVPmGXlERP6J+
+yWmDI62xH9MuMCmgtaymdY9fy3Rq929ogyxcmFtDG09Ntw8K9M1w+N+rQtg4Erh
s3yl+t3B/FaCNUmQ5IhuhynBKC1VWNeIU4LTBGJwwYJfMEeQ1Ytnx6M3kmj4ZhGa
32jTwVW1grtGs8OFUV/AZwNs4MRYq53S1wYN/YyUXUBoX+oO5AhA5Ztg4X40D/fU
jWXL0KpdzCCUbLkUum6OEAY6ZDdfFsKsgQvg532Di7Pq+5bEFbFZhXokXILs3wux
AMJObEvoowa8i4QGQQwdzGFV4bfkRSSHDEfHceabHJiWJoiOrxT9x46yinKAKODi
xBPshA3OvcbErT3cnyjGGxhIVm/DOD/I57yfOoMjg1B7VyprtBsVQfkk3h1aAL5h
so0HD5JJTCRSnd+Xysz3Yra9TSy1K7IgDI0WVmwdyTeWo4uqbn/hup5xRVABIUnC
5FLsmNDh6nV9L2OVFy6THr05A4tlcKovOtkexl5uuKqgnBaEKRcpYSp4m6lDBBbM
VbZts21UX8njyveXYYJscA00BINco14WZ3QKHMldXjhZ3V72FyvK9qPADH1I6TSi
mYZVEPglIyZJyIZobjo7Pz43bS95mR0R7hISPef3tTUII6/1OSP/B3hRg47TqXqy
`pragma protect end_protected  

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
EA5ba4H+Dmw6lnQjLXkIW80ISamgsSu2xvICtixLJws3DzJn9SMetYGPfK5/T2Cq
JjcNOScb3JwME1+cJG1M0hsydbXQvHldXuYXuftK4AkUmktgYEt3IZxtVrym/zrA
xxcdJXiMZQASHKskcOiiTuCZYlg2hodl2BA+HQiqAbM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 63519     )
LcjukkkCWOgTKc2zga1CRIws/jllhHWOxwSFcpRGtFQLrQhCZ4eF0waAiq5hn1k0
2/16jLt5LIcU2/BO4fDSlXlC3U9+3tCzR5MWBT1L97+RalQzlW04ZaX9c43985t2
arWuosZ3nwdJF9V6nOfY1d8jU9r7UM5RJ5Oox/EhF8An3peHnnIc9Es1VEg/g6Bz
ZQN/3lbp2NRkSZ3AVVdLs2l9qY/svR1814/q6B7LStY5P/lzXYQifWdF6CZ601jC
nOygtqxkRSD0jHqWJP8lvwFESCVp7/ykpHFafkiF0VI/a6EBLBA1EiE+XvDdghSE
Rg2H1kHDaARV2oVVhe2kPM5UP9iYsPV3tuV8bsD6eFAcBT6NJq4ml13e9lZ/n90H
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
D/XbWmzCEQMZvVjy7PHhJDcS/+bw2dg0zMM3t0EzT9QbkuheuJjJ3tB1Wu5lrRQF
LNS/3NyocN8B1ckJ9a5JW0ezu3y0wCRKNrrR4MdHs1+lTF8I3UPL4bo0GtgM73UR
bxJoRl0w4qAy+ajwaCDLsauxFONi+sHnQt8q0jUNSTg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 90052     )
thNmxAWzhuBFAXFe67UvKqtK4TBpeZnGi2vf/m/IP0n7i8PFLu8Ykv25UtQuJv/M
/+Z7VR23V9IY3VBEr/rddobpMyacyvMJu5r0NGapx0x0d/1U6m21IJ7aOspG8Xmu
AZypn+WBYnNUDGLc1PqntL+CE4hIMYnKc444LONAUaWqDWREyOIn81P+BxWCC0ni
7CV0bKzk2JeKELtQggkgfTvoq2AWVqkkCzB5aOoBca8WokAhfxBAWawcGLNC9udo
ucVyVTuFOdVFTxkA24Mef/J0wCrgWyP96G/sAhg7lp2ajEI3WJ4UJAJf6kGx8SMO
lv4q9oGefglfJEVS7nEmH6JOv+GWAcVOk3J6OP/qhZD/vlLNIdxLwL/vOeHwA0Is
SQAyMtrFRzPEWvNLFiXrlEBk/9P9ELodwCC0in/rt1u91iDqRKz+irbKN3Jhs0qa
dnLYRoIJ5q3EZPHqnnewm/8JyCL7UeP+kRY6yM1d5U+85NoAYEoGBM0vIUkL9pK7
dRElBQHJ1fnPE3VafZN5As3sQ8Twxq/D6gecPOYQlhPqRCvHYNrFh9ulEmBzZuJi
nQ05WlnaYIVhewl+qyP3d2HSnz6e3/dKk/VOvji81mvQ7H7+GFPD/XgRn32Y6tGH
AOAeGsxYE9VvxcyxnfX9t5HWRUwFWM3QiHXSXUoZx0DfACz7ljif/A5sAjkMKjCS
W7OxQpaY7clSKo0CCHMi1aCqGuLp3f0PygsghQFnj385iRYCQEui8efYAnq5LAFR
f0eWVZO+BBHtCxvk/oclq+Pds5mgCw1G4OV4RIF5rXBQtQJoqgcXOoBP/bMhtP4t
ExYe2cqhBgcQL0zYHpdDcHd2JVC4EMQzu4PC6GqsdkT816Rr3QhEXToEBDETeZEF
O1IdSUrsLTj0yFuYhziWFOB+865boMdU+oSA5GFsPPwnTeZlc3dsqXFuhFWnqqjZ
6F/qpsMZemj7TMcrJVX1C+z1RvwLuR0CiiWmob+MJWgd1yTF2vRN4+DvPeuUpulv
p6NrCHjiMHGM0201n664M9/zMccLGU0Xvh1CHDJJTirXwqwrJ8AAFWJWJSFHaX4L
JO/8W5dMG9y/9Lo5yTgAttKS8ygbiancrcqBNQuHlsKOG5xUAbcePOHj7iNErqaQ
kWnyO2U/Yp7IokPEghfY8F4+ECPAov2iIhZfBg4l4rb2vLqxFWKoqapMJoXhUvlb
cxa3N0moOxgtFyM5St0D8mh99BCl2yWnR/SiaJ+vepV1wp/F0XoPOeXm/i6CadJ8
X3u8w/5+RAgwMZvOAVx5N4QPpF3vtlydAOS/0VKkFA3KSYmlOKewDETrZzxmS505
+hmbOZqfHUoxIwEPr1rD8EukTnCAHu+3U7rHMjfFLwPZv9cBlGFXFymTaj7EjAMK
lireF8IDoweidvj7UuHwseRr5/gwxFN0Sac81sb7rG6qgiJYHxfjoz+Syk0Ep5ck
dZznrjtGHQuBBacdZ7MuJG0QQHXal/OUDKh0W7bs75Gmy79BXOiT+2R6eSoXj+AW
mR/+gC5pGz3hZsy+wKN4D/o44o2QvUUOJLNT8iVRjB9tHQw7fZmF9dh6WAuYcGwr
Ov9nK8MzdBE4n9GHweZYqq20lsqssfvrVvBKx7ACDMPfUJSEnfBWt44caulZPTxD
IleReSGSuc/6n5ho2GQw5Ogh/ySZCQzhrcwUTJ+Obp1/MdIOkPno2isdzswaXBI/
PrN7ZeQsriOa4eDn2eKgEwR3JmnyhiviquOytrpwbBTgdAw9Gcs8MfkI+JN9kxmQ
J1WRNBETfm/jZoGe1MJr7GbRwMQKxMvZ3fdepzVmy+K1PUL5feoBc/nb/0PNss3W
vJr6x1JE7sW5DyeqmKycIq98atkbCMMe2SXgtj9FZvhRi9CVDzu96Zpw5FGbFGs9
VjlzCm3Qoh6247qhpZhhYpDA5zyPngV17UlZkOpzYr8CjoWabrZvYBWp8kmgZ0L3
0bxZ8pK8KqcXEtLvtVTjvjN5hAb1jyfKosW6GUAtDISL0dQ0A4WYPpijwf+lK3yp
U3E+5IxkeQi8aUzA4tyuB0XwuA/VUUZOxM1kym9o9P+pxvHLgfxrAAi+b28E6Pmi
KE+HzpL7KecJiyBg5svqzJOevyxpYwHaozbgoFHas6eNYI2kE1S2405Nb9eNIEcA
K2+VvMzAxu1sMN595aika78aOwWSBULCKlwr8hKkdVLYdYl9rxAxhZ3UsNAuCDra
DxljEO1FkOPeaX7jLMUCOuxI0rwYjuSLCSAjZ5tlz4hG8ooM+yiXWYt5i1ASpwod
moeUAZtGGOMJhv55XEohgpvSbzM5tdue9kq+SC1HGf4rOgWWq2fb/raSE4CM+auG
7NKeMeNaQz/6EOK36CYD6b0YHR5k3GjSMdB3RwHOwtxHpDUuzeBTciH1CnyK9FkW
6zuSXGKaxCeH8QKjnVqd8DMou9O+NeNc/Ud7XjKqm3JAB0WEPmpYgY+64oPO1Ut+
O70W4FGhJBRf3U9QtmSsAQXUmP59+wqNTNJEgfvohwYa4gudO4seZKsj2z607U9Q
bN3h9X1lEYmJ3IXsmp7WBV1xyFtWuFyJHNx0JBz7yJz6rx8focuHbUSczHePcdyQ
BaRirP6kPAdkNtKztT2au1htpsfZRtsfRHgIVcuS/h2wTIsX92629q3AgsXHXjrX
Ejgku1ksEv5T00RSfdbr/APa8nqTRscULoe7ShsnbYnrTXFiMrC2zlxXozAJyzH0
QcuXUTt/uLa4zkxNLX7Vm49SO/+kaCBZmjWJ2nlzs3GkR7XWcQuI5efNrNqYG77Z
ReM8gGYhE/Qo0YO6QYt4h7ixOJV5H6ff0ik0n0Cb3QRzQxiEHQAujxhxEQ9dGrhe
PMCGwpFeLyCw/FGn8Zc1/tTFOsPhEC5ycEjVrioTvveKHgGnBcQg4oLTqxGRoX8h
BmR/f7OG+WS5DpR+RHwekoImwc8iKmwzp/QvzOwF1lIfuUjY217e3HxF8DjbnOSL
Kv3PFD67WAqv1fXTlT7qffJBMZNPCO/1RRmqxmoHogS8O0JH4n2mrFDRXrRHPwle
44F4DANkKsXDVtufTKjacg/voZxQ5V54yUQ9VfPGgqoJJF+1KsApXMrgvoGE58qH
OletYZDblA+vCOxO+UCp7WpAFv+o1qSJy2UVuHYUzp+NRz+IM+tXenwgwnQbSPk+
ETccBDIUvFIQqlFFMkL9xinxmlHZU3tfM4F7nCfmwknaH8T8+/LGilrPxeuPQuuV
xAbB3SRjDt8pvK/ud1GJH0ryZfNeBleSzjF8zdR+0+1sAHW0gB+AaDNhCJ1WtvJs
H7cQqXmO5CBikKlRvH7BkHL58ckX7TxGr5NA4i2DFRkziZCWdPI5zg/BZdY1G7VC
mzUxONlyskAVagXmN2MPI/w874RxVcD0jNRHb1AWYybonhrieSUAPfKB6dlbjN9E
v60CrA4wHLBJGjHTci3NspfliPT84Ekq0PrhZxB6IGv17nCNqBebA6kCmLcOi+LY
Zl1MtjLnSOh46/dh9Hq5K8gjlO4NbeSZ44HW+dPjOgARzOANWc2egsT5WOaYbfPo
/UhKb4c4somzE+L2CW3qXPKkZg4Okj44NGti9lgKloLU03giiqoURfezcBKWCRyC
WNibSYkv2l0cxAJ7q6Li2hWmp/UAp7sle8l39g7pFll4hqlarCuAeO9wnQGmCSFp
2zg88vCraeF8kKUcqRc+a4P5RQS5gQobpakNcg/NRJMTLsEiXkX2Povlv1odaw5N
f/AYYgBAcrvkD5vyspel7HqseDN+OTdo+AVaCgcYv0RTui7diX/R0rw78hbhI83u
K09I1F+kuPAbGptLuaFXSkfmTKgo5bfMb2D27h0LHNBq/pJdMFaoS/BxuljAfBX+
1K7Bi8NRJ9N0vf6oHUogncYcybQ0PnzobYQC+dWs6a5WLxrBmhdxXGLnCHeULp11
mPAdFfgFvmWmjJQqwwJGVKJ5zfniFmH4I0A27C1DixtZbnvhoDtYJEQJq9Vcsrzd
VpimDdtptgtXVSvCRnoZuyc8CMtJTOfMiSZqXjHBU6J2a044eaLNVJYIacZsg7lq
iYDv/h/KGKEnVKrVjYi6DVOb6admwR6+FF01FxZvJEnk8PNv6LlBuabQwffeUz3G
QYrVhJ4O5yHnvIeKLuk9PNDBKptRUJyHDaeuhMT2Tf48CeRR3kwAc9FNEcGCfWhF
BpZWPRZ3JV1xYGohexKjddjHkIPehsCXKmPEIZq9btMIolcroNmiMbn+tNyrUFrb
uNimBawaDiHKHCjbarvy/6aZO1vSTTdqlgHXJjjXeAPnSytgnnb5rLTcsJl3T1Bq
53YrjWuXx0TanFwDxo6kXQ8qLGs77eiLM2YmoqYrmC/PyVwvOZmloOdx/4jFjpo3
y6RaO7B5FWXQLT+UdhZ7OxqIsVyzJPTZkYhxjzafrb4jxZvNjlumN4kPLpRWQb3I
u7LaSwQIU3J7wG94pFxA+Kdl5qL12Wrr04heZ9cOTQuixgYikByH+4JE2mwxdr0b
Akk2tREH4uEIK+4BySaNoSeopsEkghA17kDBM9qDDqwcUEssQxl4/5zZcM/bVx3L
u0UsghUAue8ZCUUOnnvFaDPlez2E6cC2VzfPJLMvMVYbFCeEzKvN2u/vOUTEdUKN
TBgFwlBjfBPXdhAHksLTtwBgPBSgypNpXoVHRGzv+hWbK2ZVOT78jCSRdMKx1qMh
AZ49GerdZI2azxzvmiGw6396hcqz6fYfxcGxEcFANdCwh7qbjjL4iwBXQmn1y7Jw
j0GUkMJ10OivXYCv/hOZz0ptdrhsz9zawbzpsiZYnBqT85VJO/8syhtBbXIkeXMz
nerAd3WXyl8aH6vxaMMc/+l+IivzqUpSoWN1axxuthJL7NXq4/xnh8YK2UyaFvc7
zImsiObaNsZvHU+EaEtk+oYCbA0M0S85oVFUjHUlLF41ZZnza7hndQAPSWtL5aP7
TSZXrh3METfzh2H3i74n7w5pfhbJB2btg0F/DKX6F/+zN+LcNt7v/7/LqMFOa3Bx
ARpls5bhp6Mz6Ojs7Pxx+rB4pCJeoiUL2/cy77sXr7RGn8jHM/MFdNG9oknAIsUk
S1FwIpC/e7EOdlyHlrkQwpbt3M4WIhGXaTH9NZyxGHxYsSQZO0mxik4g5y6ej+mF
7UdpL+M47MTzl7VZJ16aEwaT8yw+BC3X/e2Th5ir9cs1RFVhLkPsFDwMm6RGDK2r
c+Dy9LpxtH1owGucZzkKGBoyfKbxvXWxbrPpHuqVCzGGF8RQWx5jbL++a0UKsAAl
h6EhoAZgFgjyn3V8Tp46P+YaaUboXmN5gSj0JPyjRrhtxsIiwb9IlGIxBlCMpKDV
LiSZzOnHTpAoMK+BJJoKk8edfuNfOfOGpno238qYL0Muy6aZTu5eVlFmkwnp+fPM
fSuOTk3ksoj6jLXbVB2VQjMPt1vHPQR1Kbo/caacORp62VZZtN4zTpbfPTfy2J12
pY0q6W0EbluVUMH9ykzoYDLFwU1So4Cudke4SH87Al+IVRcowMbSJhmVQ3hpOYY9
h14v9M3EPrP0z+Stsv4GEGgendqIdE6xNDaOe+ZCwMYRJPdmxR1T8fhbOJG+cdzc
mA/4ai1xPS1d1DIxHRxZ7Ep2GQDOUXUL62zvFamAJ4QEgbAeZgT+DSKlIYwyRBuh
pM4IVJ1fC+bmyKF1laSc3ocC4UIXkmd/KEqe7yNgCWoZ+21q5GWvOfWM7wGSw9tz
w1Oez6ktv2C6FUn6NuzTT6+BmbSChUe3aOazipJD0gXy545TCSv/dIeMeV72xtal
ep6XhvGW2o3W3rDtYmx18qLIWFz9QYg5pSL1fIJgjv9CTwFC3CG4JV/ZUf3YFej2
NaWZEbodh106zrOFrwm3yDolj7F7URA9aeU1LSCaDwJOUjDHD7wR4a7aShX4Afzf
lbRW7ue4rOlnCXb6wghmtaWYVTmD1rBINArfU72Um8JrPAlHYgjGwGTvL1SmXKTD
yP3FcB4jUSg54TbxP+2Z4K94WyI5yMl3GMURHqIMmZibyFjn3uc473SM832ncIIt
YPNIZbkvQac3JlGT49UfdcB7on/ehWDNAm6PfBW8ZAoR3QaUAmvlis+0avyN+b8j
27C0gvfUSITdXiKKKC/ncJqRisb4wGtkC9oL2ZCqM6Gap2osse6RF9CigvkWJvbO
rtJNnVoRNV5KZYnkqN/JJxYwIS2QoaxOYQvYquhufLF1OzAe/oHZxs7vcVRdL3CU
vyQpIN2k6dgUoM1q6ktly0OvYdLbXPuG1PfL2bisyeimj35CNhanMMQejX1k7xhk
g6J4MQcFplDkrcc3qHffPUtZbVYJ8jMgofkRoOtId4phecbxGp+5qALpGJccIfBh
1vYBpA8dGKH2P5tRIXOLYJJBBMQ8i10rSWKR0Dmlueee/WNllw1aonmgeJ8a9Vlh
/VPbqDtr/h8Y4lpDbEhuX2pTX2UZ1HV+d3mk72RLXekey4k3UU5MwtDX8l8962UI
GU+TUGGuMXjWLBimzBxPcFGGIlwQ9flIYkXbpUO/6xUs9z+8XjS/ygLFepfmxeg7
JxAIJs0T+jODJgrG4XmGg9d42tLkpmWBLpjmk0+0YAlO1sMuMWr+paj5bz2wGTvp
aIgYP3oYB0lzsFR7SkazcHkPFsz5OsJWH+oeMyIhTDcZtQgyr3lpjUK8L2KEWWtH
jUSKVeihchpe7gVU7qYB00h3zhrmPj4SsWM9vXGGQuAG9jb3Xnwh5wvrR+Tly7ll
9nD5eiRZw4w3KZ94PoOg5gnbprRYxnVWamGrk5JJG/hI6AdUBdf4JJdNZ5uHzG/P
tOZkNyIwxWjOc/lbLZVuJqwag15HGTSv+OFIzGfMZFQvZFjcmMHqftYYh1ONIqSb
d6pkvIjtN/aL2PXlgWKH9L/Zuw3iQeWdUWggVL5dx8fRheaSD7W25sIppZ3VfG6z
6cI3DCBoGrrekwUlfNKuNf3sZ/frqhvGdr5GWol5NHMw1zJ7gXfvFZ62dMaURlAA
vkf61i3noKDjkWs5FoHNZtGPmFAjlm56QElA3YgYTDNvctDBvWv/H1p51xh04Y0c
3L6pd+AXRol/g3uAeQY3HxH/OtW50Z+AHXdUm58K/99TSJjMOnDdtVwMrCY/zZhA
InnP+qyk0r0fLZjXpwNHc8lrTj4RTjZqH9VoBgDxws4hcteGqYEKVVrHx0LRAVEU
Fs9wl1d/hpwcvdg1+pk4Y1A009W7Ro+6ZOTD32l73Tb5DmfGflmzyWUOATB2qITU
VC8j4cyH/hzJSmtNzPYjxZXPCHGGMAuGn1UoFGaZCS6Ye/t9IXl+7Zg+HFxGtGSZ
vguJIKdbXkZ+fPChwYRFaqGITP5jgk41nK2VUP2+j5gswwLuEFPIzpaYNnv3sEIW
yc3BVM+KRl1LGOMqVq2epImZ9nhq+63/mvBuMF/Ksj/bRBWkdX/Oe1o1MuGPgTKe
Bk8sT/9/Jm06CCaepHK16zhKlgRHIJ4oNFbll12gU4WbTWdMdHNtz6ey97suk8iy
J+jvHwRlpg0U+bXuqxTPOPfrQ+0IgZQUrhHLeLPboVg9bPQIM1h9PVRV5yxh32lg
32tMv5Jpuw3iarHbwxAAb4M4gHzDxjHLf0BidqmyzRa7Gzw/sZBAehRSQocP0BEi
857Sx35rpqgZJxCM8NZhxHqYRglDoxAJciWlkbIl1zHS3ocibR2tlSRXdF9+tWSr
QzWtxwm0G8PQcUVEZ4PgCWdt87YsXIOcc5VNkauEr5YdFdiTfxWJXGQP1lu9gPFc
pBMpFt9vhsrpVzkyY+IPXJLxcPlzrtybQgwKOISRIPwgdLI/YqiNqWNIHsiyUNPa
f6Idz3AqGjmG0mqDQL4Q9eoWM5uP+6qEXHdA54GVxR+ZeFcnOOpYAFHehVTsUKP7
8vw5pNWJY4aPS3ndH0q4eClmTsfq76hFMcjPGgeeaNXtaT91+8q0bYyihl8GHz9G
4L9zI9Y/j9dWp2OEa/f/qftTg4t6Al/u0Xn4FQmSpK8TAPghrMw5MTuUSNdvkhcE
2Ms3MYijjYLFR3eNfBTHxPBD1HRrN/LrJWwIlLTmvI82+bYed4pZfRtAPmH7k159
da6btmuU25SXtn/IT1tqBwy0jJubITqpwDJ0uW5zLV0BSdMUrdTvHclQzg/aeBcd
F0FOO/bGmhJ8/DrLtOB8JDlDOYbDVicZupPGuNbyfJUIShoFmhYuH3Szse4ta2I/
FMcvkjrfvUb1fThdGHBQVSQu2wvS7nv7TK/iJGp3iauWSAegQGbzRbF5t8mASdR1
rSLjaXg+slEjOKWWrrRIhA6KlcfAP2hbQjoJF3y1RE5YjvEg/5h8PzARtp/bp4as
iuazoHPCDjX8EEbaP/rU9cJWeNrv49aWjZBS1ZG9J8sGAf8iMv+wt4U0rMYq3gNi
4ux6vcWNWK95uyuBybjWkN9vLFiyi1bcLiegx2pirDEyOCl+FCri+ICtVLIBHQem
d1DDLj5jQXLrY/KSBTOfXANNNpWk7oitbO3wGQUcTIqi2GlahtXXDeramd8RK9eP
dD/ppZho76k2oNG32tocC5t4Y6DMCiOR70rcnR3Kngp+dVheHSs60COXf04os5yE
d7A+bHdoNDzMueUhjs5bF7H9b+Ij7xin8hwOQlAj7csYHQS3O4gMQJ2QcdIUT+LO
wXzvrZYO1/DdZFZbKtpQ2bk/uTlrb+CcISOqIyuFu/TJoedbrS+AnY4SbqyK9NN1
KOD36qPYFSDMeCoV9Xhuw1Pf/x7nzezvx+b9ZILLB+rPOfR43GGBkmw17/vuQ4Av
wksNvokZoENMduVHA3DsSdCvStS7FdLVfo6Fi3KxlvHciEu4RL8dE4b8giQaJs5U
ZXklbnyajmF/utk6wCSJ8zyq/WwdrdHdIFpO/oL1TP6CUyrqkuwyjo1Z4LQR0KFR
BfLGBXaaVx89eJKmxgsRuNUCLOMIYzSb0N6apkf9q3aUIEYBdEx8mVvZ/t5AdXwT
z3oBK0wpLGlpOPg/uz2CQyOuDuMsxyAKLCBTKwQZxr2MA4WoqzFBlrkZTl99MKYz
o7ZC3hYyUyhSXxnIZQWKUdk3p3i8s6/akYKrVQNRnKDAIK8euTE5RPd9t8KIXU0a
/tlTfV+6/9VOda3x5sDD1La+/QbInyTUGZedHDUzK5PzRR2o7DtDNfXpyii8O+EB
aZIMzcwO7ne0hM8EZybz1/E5SaZbutm6I9ULLhVBi/38jhXjAA64JLGdU+tF/l0R
JCTG1a3RVRJVMiReISfvbPu1KkQoHSUBv3GfOgMNlEVQ2l2pWSYFYuGs/2OiwhMJ
d+mUP6xEqTKF1wzeqm8V/czAc84OS04z61AaJ9pb0z6eZdNFasEzrxFQ8AXDlCWF
WABn6MCq1QmgPr28iadkl1QetKOZlZahX4/4vozzUOWrcC//tvve3Z6PL3d5QRkd
/xb7cf9uFNByV+C2g7YSMQZsGdUr2fVwFAOupvVNHJzQLkHUcSJ99+9wEgoT01QA
aU+k/Q12kdA6GjN1rfGGbK5FDDImxuCVnYgYUFNwd+DlovgH9w06iHJeYf0inxDo
PjTJNquu1Jbv9H1os5PrnK+YyLq8yLdRsCT/d8mI3lm8eNcUpOm7qkyvz7EvUFw7
NXxs58z8mkb+4XNLzyL5+6XyRZfrXsMHvABjhd4cI7wjintbdxuaw8Efd+d44yEp
OrQrV05GEAK4KoDRfopiw1f/UmSeB3jHfmawIh0v/e0k38lPA0puS2n9KAare9An
0u3iBMriGWoWZ1Nm/yM3mLDAamNcOelKry1FAognRUva2AEamwWJE0AmOUISdvya
t76vwXcap2yflhhz4lIRu89kjnXlLlsnNkxomB3iUCNnv/h7ZvMYVcZ7UuunDEgs
gtzpTCRPSZp1f6vHsHCo61awVJew1S+QwxuvEFKu0HFRwle6OhVB1Dgjk90nSE8g
ub7rZb3z3WgpHE7NAZLRsndTh0YN6SV6MHRlFWeK85B9t16cIf918rFkdwDIBMRc
/hPaAjTYOJKwXLK5trob0dRypxI8886U7d/A3UkIx8Yd+3A3/7m3ZmeUC/Aajjec
5P2XB7N1O8a7d0TJXqcIhSZIOd0P6rVSHaFP1YURB+aJ2lBdnJF4JK2w2kPCGyjJ
2ETKXd2SLM7QMfru0N/G1GZDwT5nFBvkmUscthLD19uS9GzJJN2VRghFqfkXjxET
GATccUkH4XgrlsKfJ+scdm0n4DoVJiLIdvuC91GVdC/6SUL4aGGQKtusXC+08f9x
mffMX8r/AUOdHWR72Yfh18WJDXtPIV6ogOPq2r160cwHyKaEGEUgRyIDrMVdxfEq
uZPT5IbEoW+VouiHx/LcBVRqTDAdQ/2v/p56h66a5Xs0XujwZa98T24SBkNf/Q9H
H0T/qYk9ko9PG4v1ZGS1UK4AgUH7hCW6hi+YXHRXnozdnXGKMzZq0f0mbdkRzf5k
PTME8hcNYEpEq2f84IG2Ao/8Bf60d4dA7smojCD0XPl2n2TFbDab5+y+HbznMLPU
xFsrbf8CrP1zFRZ68aIuq6XyWL+VwhQbtOx+c88OHcgXujAG5t0SJLVLBj3Ln0qO
IMZsarZgucEjctl3iwmn2MW5H+TY3EBJNODqUVzFNrS1AwWjDPV/GQdgAEzFHIA3
dPyI5+qK4VGVoOcpvgtlttWnFch5jzEpR1HPmGz+jwkOU2gXiSIiuXjmoIxyuJh1
urdDhyudehPRb2QAgjZCRLiYaVRRADfJ+ySDMH6HSkz6h0Z5kYN5MxtOV/Dj8bD6
iSTaWttqcGvVCi8Z4rbynw+cJnjL7ORc9W2lFD/EzXiqjCTT5HMAk8kUmcT1VbEB
nTebUfWQOH6VnidK1YBvsuaX6YX8zSrGIQauTtZ76Jpp0i6tgJGTuNeKJENM4hF4
13NQzujpHij7bb/MBAt/ghG8xqcfHyr5s4g81uIWEKeutzovdhfxXoJBPIDrZWDF
i9sezVfJaSD3d5ukLutkoj+5tRa+GRpKyf5rkYYkoEanIqnPx4QSJHGn66EdVFq3
gYOjYvnUxmLHUkEaIg+tr8aTO2Gi7Cc5DqmRPgnDI/VV7cCK4k4YREXY6b5rRG0Z
lQoEeBUzFFy+hBUoS+zEsBLv8Nml+LHrUJu0cH4tJOhs1RsoQXnmB58L8eudmb8a
xLrFtkw1IanS0FAc/oF++/nyou+05H7AQ+RkEngC353j7iqvgDyGXN9JR7o66gtQ
vYQV3+TvvyGlAOsE0dzkoa9DO5aooTU8Konvls/I+pu43j6eaEjbgFX3RklTzJwq
yUk4IZ01c01wr4DG5YVWsenChBUGQ8+pzVgDeb7wmUf/6/qwRoWQs2liag2S0x32
rODSa4nKEmL4k2fPdMuMpTQoQApDuFicZS0eND4xp5gBYIpveEFP//mKsCRJ/d8G
zOyLK/FvBDykdclEkhw33P5HhyIEq0+lE8VB3GqafjQrtIaEXJ9mHlpbJYZJIqZq
4mV+9KGHz78xh1zf108d4rNXkMMO/O763vbinUOgLDBm+Tq6R59ONTL7QUHeEDzG
T3Y1xdbrPNDnTmS7yh5eRGyulyuzxGpT3p6UcLpIAcBKer92ITS9dz9TzGUvNS3I
nMwd0f3DjEeEYwkDzk6dXjwR++Zaj+aFiXlGBtSYQFDXOoC+eDpBZ+VbFRtxIPqg
wrdQpBHoj2oIKiktgNfE/gS7XzMkz9/+y5APIfGD+vvA4ORLzfAn9tROKzJXj3Po
7rogn2r8Gkn1g1Y79oQ1ZZWWmkqerZaaQQEc4K8+B/4t6VW/Vjk2er3W4XPPvz+v
u6saIybKjTXwNvUjNamLat2GTFz/j4BrCyoIUfyVDBZLxaMoyJism5YamT9aG+YX
ZlpvH1t2B+0BQlUtCFMydxCDvdI5Cwdwy3QMSNBJEQHyCiAR9tLt6I4eer8KlWXg
TXysf3DyZ9i3T7YxF7OPZhBZPwTti8FWW80QmV4jRnBX5J/YYOBLUsqMs0FvRmC7
pa4QnqglEG5qmvYtt9UEjYrwcvU8o03hvSQxJuNCuwVEgfmnzjkmcisuPuswv4RH
VsPm8vCVvsHv79SPCFON3UYyuk0SWXJF/PguZ7nxBPevQeWzxFq2ZRXNgkgESMi1
nEEg1L5yOD0lSzogBpG2tzaao128qTVoh1QhtW3V7uAfvNT1PuLilxFU8F1FHGs8
VwJdRa9d7tmzXcDAnbduOnV/eU+2IOKXHjjufcu9WPAOyt4USK8xbZVMHPF/EnZB
qTGUaqV6nhXFe7peYfQ4D7sBI2dfaD4aa23aeuNaqbBdd0NlHDnIT3xLRuwC0Z9m
OReTKO9gWE6ntuOmbjEQf9y66Ak3XpQhrGtk/nHC8CKG+dg6rFGDUqVEKtCIvKUi
jtn7o21rKUb1l/7eACBA9kxr0QqVT93XMNmKk2YfEOWSWZkgGLfnNpGIYSfpvvXI
YmYmQnnJT27HclpnjbZ+JYNZ92mvb0quw/plqWCWOZC987rK0tjulqHOR3h54H/u
ghw2fRJuuNmIwUWhRBo5hcwBCBX5Mu7pcmpJ2oNDzolgc+83nbvtEN3xGfjIvEer
KeADCknfJWtm5QIiThbMIN9SO072vYKmYKtTh48KvOZ3lDPAnecdTVU+seM/16gV
61OvqQxFuO2ZpC+yTlJ4JNl6pBIVoB5bttVCp3dGWVUJk9/xfENlMEzwespll87G
wYmRUQsrAZv2UZSj9DUXpEoVCmBpd6CcmsAA+CcqmS61FrE99SKA2vkLldvdxbHb
8HlvyZcnqjGz0yqxU3LIlCv2h98QL1NLHLKRR7F0wHko5uktZR25VdIEcbA7D4kI
wcQnlWewztRgkcU5jx1lQHgH0tbOm3EY/f09NH91rtYbOtW0QFgwApPyARAgcI/r
VajXpMxycqaXN75WeixEYRRWzmkbbMhdJ1C9xtScOUT3hINU82vRUsW2/H4oesYs
SeV5LePn/uTscFLfIfiZBYXwVPhx6jzIBt60670WgP+AS0Fh8gfXve/HwjoLZ68y
VCDL7E65UKghh/IHfEo4viKuXwLQfndUeo24o+2V0w5LYCkoXqQGF6mfd+a3UwcY
vfDSM0vwzYRglCsvobxP8U1iPROQOC22MzQCRWROWUwAxVNw1GQNXVne9IuLjx91
3Fr+gwTqO+D/M2XZit5l44RL5LbrsG61rKO/DFTwxeASopPyE6Kjyt3vI1PrWOwd
HB1LU1h6LN/DhEYfEQFHWomysomFSRNMUj4HPB/90Cs2EbIyvzRHhROp5rNM4wCQ
iM5vPDhPXYDpJrjSYDbzed5tGduyWYvOLywYO2NquAjL1bCgmAQ6kw6DaDXPZ83w
IgcJqAr5q4aexwfCWFe3HU8OgIXO4oR41YH5VvSR1SI5xHgUOFknh/roGypdQWhN
ZVaeEc1iuFU00MDlnN4v57TYIIy4VkOoM4F9VG3Sy5SrsPXPEch960r2Rxvm1CNV
onj7+6ddBmiF+RBWtdFAcLAmIW/5Y8LIddA5bt/gdIPlxmzYlSRKmvOmjnIg7HNQ
iG7vJiVL9G0D5pqi2up192yz8XdjzcyG7kmhJH+vFH0P7nbRvGYuIvI9a719By32
Bm7ulFvA2PxpRib7nyJsSjXIBnhpv1ayUI8PReoP3iSPnL5bA0FSGgm0v2bumF2D
u+C860DCfdBSKMKB8PpI2nIa6BGDYfm1iH4paPPQgpGhMhhDppbSb/cYtry59LDL
etpuRThuMW3CLjDba913nHRFcmtWXK2PgLu27a+sx47qb93Aq3xvif9IwcaIkik2
PLe6/x0Qw0DoANYZMItlt7tVjWtmedhMC3fOmDcfM9EGKfWmcFKUC0RHk4KF88Yu
Pvynq5AfZPTdRthvU1U/L4fbqAtKZPTVQn8GvX3EsU5XCxHA/r+aJ9STuWAJjN+d
YqS6tC3/yJqFdIK/e0e/YPHOpMWNZw7VxMBWdjBi8on5PfcmV+NzEowNgX4rGOOs
qMaQ+wendiZWeMqNn3PsuMG+jpDI/ZpGS8xRHmv5mYXwKqTrXb108L9v0Dc7L8Ti
9utct8GJEUf+gb8VYEVvANX1YXETkHnOLTg0Jb4r5pegEQ8NX4mtmL4l1I5gtZKc
Bs1hRkaZeUCfLi641oNVm46GSxMiWrDcup8XQ/aj5DFmK/eS6DehI7tyt08et8LM
9Y03eCn9NFs4MQq2x7YoUs20zmJCFizfPUuBmkU+vx3PBfu4Uuh6+s96CPmoydJQ
r0vxmKd2M7CFjELgZMeweRv1ZffZPadDYFXBeGRYxcBi4ojBsHPWWzzH7axwpwtb
JlXhIlgspGWV38XTk011pMLhYkyz30UBL9KSNbPWpITqK97nXWXY+7ng+65K9jtO
a2U8zAFIXu/JniCu/72SIUTgJkpj1yFFlqEmeLP1AtUy+4fy/gSH6rf562zY+/yj
ZioTBkQeZYqNDLFZ5AgOqPvsnRgvEa/TZsjq59mmiQIMLwr/A0VdfBwy5ttclkTp
Me3gUX+O8ip2hh/jKACNPH1+ZDwtubv32U0c377WK8n9XE9d4jytUINN4l6TEYoW
MrIVtnLn/s3NJfqyx45x1oZZ93Iv9cXR4njtz7bb3BwEwQTGfGI6Cf0xrpbEsTdp
0x6BquzHnAW31f7+pXiS3CIX4yU8PiZEui5AahdzOgF/xUwC3TpnuiQaiDs2hN8U
EWx0+ILHpW8Qi9xBAFea7iyaLuYS+ve/eWH7Q9RvaaKF37k0TGO/fnIU4QuKIdAB
eBy1MVMOUFp+hPBshtk3GMuYQ5yxkpUaf+ZwCcn9OZqb6MV1d8s8ThXVbf5kltfL
XzOmJRkp3kTuAcPxkwn6S1IIVJ8/wHuDqlu3UWR7vfXGUVp8q1+kbYebH58KDWhG
NPpHQS7qEoKAzn+vQE+yCMnhum9qN3ExDhjFG2PUpAe/LV9WzGckst4rsXEIQtnx
3psR1g8PAePMQGUqKEj2UuBnapA2BltDT3TEjiDWsYLJX2vK673OgkKFtNectT+t
MKe49Rs+PuT5IwTL1LKAp+RQ/Im8ms8w7npSBJajZi687pRsd45Y1y3Ri15dSPc+
bglaAbm2CibMuHU17tLYQG1cU9X/S+Jl9sWSltltsMYKkndOKD20xwylib+sqmM2
Hg2rg0qBxIF7zyixZTI6Lxl9xB/BZ8IIb4Hp3ruMnGFFapx1FzSxDr8AbjZESlDv
V5JWi5tK8bw6vGolYiaf2i9vfpHGc4BmweTQb2OMv91HXE+1ir5S2sqg7+GZiNMC
P54lJ3DWBsf7cUPlziAS/7aEwOitE/C3N23sExyz7G2LpJ0/zZWjHTOREpLGgNza
7FfLZ6u8wotpJq2xpE98iMy+KWVdl5LlXsvGw1XwBHFC5dHhCJUOA2wTuAK3WMtE
tg4v5o5U6WMFoH1pMmzkcVZVFw7xm8gQJ5Qc55F4ko5PE6BvREtAzMMps0EjJgMz
DcFkMEaDvnF3BgSCUnRZnQNNpDkPlsd3dtKyVLtZXzvJKFkpXLaOp+UwmxzM6iqk
1uuwtbodxMMf3c06OHY6ACo0UqDDJB9NZO4Vej5ngowORMPoOAllNIszuzWxKqSZ
bgq5yuERjqTttDv5DXa9tksdav99ndJJkPFAt7gyBUopJyB32lORf4EWlOam8mIH
GrQOH8hHqiBzAgRM6NCj4FIMckr1Ouf8n5W3ANVnl/wlJFoCtV+A3fEguK5hmtZo
qKR0ISikdHY5SBpj974Gzp+ek/SmlAhFEcQAG5mL4SxMQy7iyEUMXZ8dgLfb5Lts
xnHlRkzxANgFqpPhwhfZqifI1rmC2MvKBS2v4l7Gj8WZJTpKNzrrvevQMbxSfAgJ
dulfHdrJdjpY3sxoFeOPS1mLl9steULIbRnBXKGbt+zdK4UvxW6e3dXdjpYPTR1I
HZLTuzjBqoSceHipkgq0zC0lmFYDN58vu6O+x3pgGWM5iG1Lffb7+NGOyPEIhJAF
q/DEk3MqgABc8d5PFjrloQM8yOc8hEXsBP9PljVRO6UEmouVdGm9yaENS2gdnLZk
6H95gs83i7ToN5YKqxNgOuSqkZkPhIExZyHhHy5tf+Mt3vZTQnCQ3U4lUu6T8c4Z
gRrrHaWz9G0d2t7hQCdQxclxhJrJJrsPA9CZR4rVwoR0B26tkLhBVJGsM17+9Jbh
CaMMKm9rpihXI/U8D3Gf49KtLkVln2/rr17SmgMVJlrltssAGE2gtqLsZyYq0V1E
VscoHbj1/gzHpIaQukxfJA5ajbxPZX+EY0i5UmqnXCSrLNMyn0zwnzXn0luzoBmc
y25ngaLkTY1ShFGEHL1WbbaaZhHca0ydykRF4d7/UV6xaz1RiWUa+U+gn0dlIHHK
qHGDDdD5YbBgfIjGcC3KDAiN2CCdCaZCpsqq3kBFgrQ77LTmP3PEumUhhYu/ewYj
BN3K07zLBpKxvxWs1qLKQ3Je/IXtacu0rAAPBm6Xrm6GqRLVh3sfIYq9mF05ZqeQ
dH3b7gKe670GuMfIL4RIZWlN55ol/uLWz1E51tcu0QBR/zH2VwPSkLuoEmkGsZNp
V+/zFmlGojG0JiOqwQ8/dLM5DwDUalS2Ca14JCJ6oOhm5thOr3+7EN7UXiD7Vf0N
oA042YEqYOpVerwdXWnJiOzcsEYIXQFeRF20uxtMYICdCwpH/0eSOeDPDQ6abdzG
6aqaP1JhOimxXV1ZfHRmMAY9E2eeWI4PqHkkADoXXGBZL+oe+QhKbTPhy16wR2Al
iKFT6uYEn7hduvIa8AbGsE7Zs3Ksft2Wa7YzFWnFYhQPHXVAizui38b09vAsY+rP
zyRMVZVOV+Q+94Pv9jx65jBgSuxtWa59DKR3XFi+OR1zjUO19FGFR1GCuepf1vBs
ahGaBRilFyVC8Tx3YYqP5Bu812CrAzPnT7psXkqqizI1pk443LSki5uBT+T9uPkY
+DkOLJ9cSTn3xgxSN2V5g/5TtkGvT532UXh4m371T73/AgFzfRkpjrMirfkzlOUt
XqitmvKLfjTXZ6zZTtSx79AwUpOEKOVw/gB7STVYmfniFFPwVxEaDH5nS5sEyJp3
FNtS4fb4eWvCG0Mk8ne93NUDlg31Z5b+HzrdzVveA7iLUXlj8peZJHUxpjI9rOVx
vVV6jBiq2arWvH+OxfBQ7YvJAX0Gqfnt+oobOBBKDthL8jUnFcXLaD81IgWeqGbx
o6XX+XOFWsLy4QzpQOtiE+ODZRy6eW2NWJLxhaNY+7kkRQ2GwnPApO8r1gfyUS17
IKCEr3yPm2EAERZ3xuph5/VEj4c0EaDmsyK5v1iqcLJ+mPFizn9HWvl5z+yEX4IF
d7Qpk3sY5ILMVum6zgRp2UhSG82HgeJtVe2SBbDLRcED3oLMTtdaxOrQvm90AjSc
mf8ZdUpkQKe9aTzfsdvcRowoJqiNyt6MIdL5JGK6DZbARl6uhlVITI/5m5q3z9/D
oWZ6VMys4heIoHOWOU5i7xOs0DGFSoFWWU/Q8iGGDK1QjHk8fBX8NELp1nE0Vsqq
UDMgtRT9Y7JZyfEL18ccEyYQxM2geKHx4VFDBXV/9KfKbbEyhX4ZfsbKGCqm1el2
LGrgkYy3DCx6XgcAdAkSZvsCQCa33Twsb8CXEBT0Z2kXYiLkuigeYpDsI+Mw+MV1
MHDie1Tc7b2+FYoo54TUDQUaZkhJNxbyopDH6qhIFUa6IKeuFpyd8nk3nHbjenP1
qkiy5zEKF18beOtofuJF73HKIdH6AjpdeIqjABVQYxic7++wQfZq7e2JyGoN1nt1
5uVKE2vbDM6X4c7bgaa2UlFn+BOwAopuN3dCnhvKT5XXrKok3+U2ZGr0Qyby3COv
Bu2ZwuzyTPQln+TPv6IhUV7AwbDMciaAkgkzLUvYkQoWRsJkJ4cOEpNj84Wts79h
6Th+zDJKnhu9d9nhRYOC8oD3OFlVPyJom1XFXdpyhT1wuuIDqGMG4CNb3kcRPAfY
bMvv03lMod2062FZy8q7961NV5ZBCJ6CqTD1oy8m19Omo5qar6bHfRrYbL/aOPqM
ihjPqNNk2uIPl0hR5wTuNNMZS9eiqQ+fMyx6z9T0uJOlDOJiupWzLK/JGFloJlzT
ZiMOfpSQLaUREIBATAK7Bk9PTMzoIvDzX4IZB1NXtMjQ8oG0IKAU89GtjB57yQel
rWHibFGx66rLReV25lprQinSYBJOfC50f4CqcmJC7hYUXLozgxXdB/7v77EZopvd
wogIoKb1lRQ5Cq5JYx6eaPPbkNAUTMPQ87DirhJkxKy2nzTy1ZW0Z8wfWCV1bkfF
OiJSgkCiz4U/86qg50N3D60Pc/eVL52XFcuBqEPx9j0FjBs8O71ZileTwu4XnpxX
29LRSkOyIEqciUcuTeVmIVSGWSLICCmVWGNGzv7GoiTjyKmPrZRVHHG/8CSNUsbJ
kC8siAPds3uGMDaoNF6AK/X+z+NdiHPRh4t1gEQsg4BRReLKIIUSWh0stZ9gQlnA
MgS3ZpDVxZHEu9cfgvaFWthuIzj363ttO/f3BtWJfFgsxqsnGIAvePqB1gXNGGt9
USgZN4sFHAB0BMm0xQi0aeZcMGBOBjrmZscw6bqfnf4OkSS3agUfLQ+2mCty+SWQ
RX2Cis5Zy8ou7g9BWlCtAoweIL1oki8XJX4OTDgw2U6IotU3Ba2LlqAZQQIZgbfg
+Skg4vssB/TyRcVYTetkWo1wz/nyo+f6Zt1bQg0OLeTWoPZiIjNPtDI/IQUQ8w9+
H3ZnFRO9sdsSSPZCRt8+V5jPn92SeAU6ZIpAgrUEdyw5bBpneOipfcAhAWYQo/VH
DflUkt8SlIySwoJPkf0GqeEuosMS3CFK1GQUjOU4e9Md5G5pfp/CxfbESkw+cxZ0
Yg6SHLRdzfgWAWrBPyK1UlJrqzKZUIG6KgpQ1gGoNVwjFM7TPuPjSKketGsxqeF+
hmxDt47Q+S3PaqvyncUcSFxTcwJ42F0UngqjqJDLMwHs4vDPqpckmQXCsCUemt7y
CPcyeX9FnB7NRR54uMyO2DkYMjsrDe/seyHyLNx7PxVJ2E90FcVC8irLTnuTSEXo
q3oOX0LSvABFapxvYhkqRW+bh7fUHiGbIVKDkRm42tc2PiLU031Jg7AfR2HPEogH
+kDEfSVF3TiEUE7IcKYxc+TB+fMzEwMytNj0olsz/B44Px3VlUjVmI3tjrSebcFb
L60RlnedUnKizUZU1+/Y8HtfsncGEqIHfxPRjlznPoysmiYbDx4K9r7zFJcvx/c+
+KOwvMQ0LMxNb1CUildapAjisbAlB78RRGWiX3mAJwo8iynS/kY5mFRXaAiJmLXU
urHd+rk1Z9kAyi9KJjF2pncK0DuRS4N+YMqHKGLOoLuwegRxVyENhd6j7VljRHcv
6vEU4VZ9LTuc7wW6JNV3lsxxdHjrYu2rVohD4chQfQxIF6KHd6eyW1GmbrEg4hCY
TxxacyGtH7dRcqCYaTPFA8D4n/sN9XED4uLUlZi44nwOjjyyaL+yZHtm0JHV54zR
Qv9ieaTfVuy/2276qCk2bABAzaBiB1m3bXL9Pi9j2Pn18OkxicYGkWKeQIw7+n7z
wQqNeyUbxQ6M1bQO1635yN3fkyQRbN3emxoI78e1ND1NGio0FTY99G+AOLMWU1AS
fOeHROl8jpxp9MXAbtbPTBVGZqmozBLr5HhsEklb/thMXFmrSKZaBdzRQhS8H4Ko
DKn3eLN+IG4A+xkLMIhnrHw5yY5WWNUrXHTSKGAnqHGOAxyom3V/LPnAVBnsxuA6
4TpWbkfi8XYwe0pCXQlDnQaQx724uas9aXwH2Rdo/MqlD6qmkA9EOfhycBal/oqA
DYVUlR+5WWoEsBi4QuQHeAZTJDfAyxRN0jA9MVMkJl+jyTY3PFJ/XUNEmGEMIe+o
W2B4y7F8JyB87oTawVlxjCJXXbOAijppaUPRNoM7yK0KbpUhqgrQ+dh6LU7imCge
R9jnTB4JR0l/MFuoSwWUPefoWexOM+MdtiNzVUFOimko5HlbtlOPze54TR1cI+vR
/ywiskYHFezzL4WfZP8/G5al1g1Uro6DhEiFidkBP/h1g9ukTG29QubRj+Ien2SX
Ce/EIEiEr535LayXecCCDx2NAvIMHpk6ceQNsMmpSsylrM6GnbgCt+nawW18QYgv
gs/2WZze6JaecPoyX5BdEWUqzu2S1jFtr2+EzSlE3P4Wrm9g5or17R0CfeXYKBqz
CzcAbY/IFIPdXeNkjkUTcJCIVLyt1iXj6Tp7+Sm0Cdm1RcE8AxJ8vKXo5eugCfQ7
b6QTfrO3L8I32kueR5fHSczw000i2lzTMkW5BVCoBFsXrjiM5lp9TvVXksk3qHpl
fS+KjFkDZGGBNvc+Z6W2VdEMX9pHDcd9iORww1giYZ2V6XVkOVSYLr8HXaoBaUIf
hLe5F4VphuYB0OWmnc9shQ5/Z5y0H76bSu902SgOLPn5WNjXPOY4B/F/hGr3T0ZU
JWD3pu0aMm3/jyIZ6DXKtsC93by7OvTBOgSH+uLsiTbHSNshfTrrCRniq/6DZGYn
+gpYxftor3SOWXWcvFhVNsk3dRcmBqPgEm1LczJb9lqcHFCJmx6ArZANVOnIOZUK
o2QqBEAUKY2CvHttJQsFx84r9x6RSj/Nv73fTX1fVgGGh7IVwMstPpQ3F146C9QX
8SulErnZ+VTKTplYTwjZ0hSFeUMbPuPEtiXgZhCwnlTQT3+zFc6QDC2UpJWRtnCC
DP8i4Kq0N9ZFjtLEfcIgcwMxjzgnJJLU1P0g/RSKosunWhgmYKXpQrkohnju+9uP
7GNmIEyGtO2IKimyZWkdZtnca0szbRD1rVMY2Ld4fxQjP4qbyu5RS1pS6L/3gfO4
IGsUpee3v3kXoM4vc9Z5bPsGO6YS9h2UmpZHW9qxAuKHeo1BalKxjF5rCrDsCUhp
sgow6erPUJxCxPgK2w9gJIESZgFXkbwye0jNHyAGeajfzgENH3ufWKj8FkFo62WI
oT66R+hegRjzlHTX3R+Bbj74LnRI4mnUUrSJ/m5B2pubGz1PbK+TQlLhXjbs0/fF
NaQynyM6nJuKopTJL2t+U/aVeCrb5uBLJu/YEyU46+hSuNhkDOjB28uVpiXb81Yy
wi8uEmUxCxfw8zzkM6hiMbIgxm1G1WkSm24HO1F0DBoLq9Of3No4gHag0GJZYDir
IB755wjmlzo5/XrSZPLzkRzy7h0f0igJKnKddEVIhZKqnKHAPke69PSHCFXT3v25
d0bMxPwzQPS61y51WhN6ij3w5LUzQg4cjhEiYharx6HRyI8bIfYMlHR9Lw37LH+i
+OTR5ZVgetip6bcDCQHLffc2b73aSOY2CZG3XnWfxbSP27c4PGaE/buXR6o7lsjm
++G86sk3dxt+GH4kRfZqofI699R7H6qVuk5AANyz4LrTQu73qR6/IO9myebVZ9ei
6SEzPnco7iBztdciwT/VyQiZrt2y1iJ1deEmAvoacPyW7iU80zqMdeEJTVVUah7D
q7Q5tjvP4Rkl5CJp8uxxx1mJaTfLxhdOurBmJsNrvJ5+ho2qh4KCsQr6llzOE2Pg
OU0OTZ8DwzPD7IYVj1fK7ZBnL4N/8q2rbuWmLBvcg4K6E0QKNFSOQNqKA+6DWVu7
tbvpPiWHcyeaKHFgqtlgFMlCk/01uaz2P2MTTWH46l7MO7RMkG4a6CexSAMcFCxP
uhXfvwIshqjlRtJL5saSk8p7BDuLsCGCp9KfW9go21aRxftr4duL9dNFdD5mxZ9Y
yF6QpOvPlHkYv7yZDQ96XUkcz0g0lG2pfwJKA1Rlj9/Fux4V8SUq1euYUkEKMJTT
3Ek1ifZ0TaicTwFH5CEtMwnZv+gedOovdhDHe8LxVbNbspgKafZfDhAUCJuUvAqZ
2wpxWh1Awg5Ro0XzUZsc8FWBQ6e0IOy/zzhjoe1GhtsmgUT522WAXAAMYIdlHLBg
2UQ6MEgGsHiBlk/sB5p9uiqC2ng2T5AfR9qMV5+QZHVoLc2xf4P6jMBt+4mIu+vM
Wf8JOvJNXjqQ27Tf+GLr5SAshuQxG/XI+7/mE+98uTZW1TingjADQ/+bGqxKD7I4
ILRQ63w/wB+SwKihMdAWwsRwrZ1uWb+P0MTRPpp00f621GMuybJHYRPry/B+WeBL
wXJ5EGd96MSjl7YMLjBRODEXl1tTZiBjgR6rxpvchmJZBZfTk+250ch8k2r7rgX7
mAXAmURiE71ddUANi/2NyiHNClU8eEQEXX6YE0l1g/Vz25qt9yfnl7dBPhC2KL40
i2TwIyx1kQADR78Rr6DqSr2ELx2eEbypqlrySCpZMi++XIc56N8v8DujK7sr8iUq
eIZPXFEUODsORF6R+APkSqaqJq2/WHfFmUEN1a81oZkxLgTTn6159rgkNjJetpo/
YXRrAZW9Xz25bo+R2pmzBCeQOSFdxxd02e/OpEtaAvrSMrotSQY8p/Xg5liov6G6
7j9oN7p8aJWqGbI9xFFHznN9ciyZyE0L5M8LZVOtnocmGYt4xa4mFR3C2pWprtWB
KMNUh3v1RmUjhtYwQCIllXfMtheleyO8w3RGEdVAmZd9kMRNDDW638KumjVyIDcO
vhf4dkGo5K3Mk+fAgsJX/W2kuO1haEAZ7ZhQsrc6ZjFBETqO4J2EgAkDJHKaKxoO
YeE9zZ+jIsMKrESO5DuZsnq7P/hMtUjJA8MGfJVUO9EDUeMKjIhqYILgLxq5Q1f+
yICkYshzGQqlD8AGcLLkwLaEQ7SmgPo4SGzPBB1CphyGCHBIzhBoUQ4OFZojCcDr
mMvXkpRYmr+wIJRTQQ7zS2T/3mUy7cgnLohVHuo5UKBT+sIiWG3yX9U+aaOMa1wo
O8v9IlUM69rfC8wLWiY6v4rDSdpzjUJK+mJTgOPzsqDXyjeQYohdRvHEQnN82pVp
eXAfTV+5GftNHquRxE2KT44PIg8pkTSEdDSDdMM7Z86b/HefGoDk7ZYsWGn3M/p+
IkElHyrYjkrBjQ4YFNQMgkPDTLCF2lKu9LdIFm8bx6j5V0Gx/UyjdFxms6kjT1fn
KTnURYZtxY3knsURqpZCDeGXrcxzHlo0RkaO/iSQDG2Drv3w/9FYDOF16tKrMgUS
oEsIZVu4l4DoX88dmip1hKDfhViNYhFUKEN4G2u1E6UR7KMVIf89HxcVvHxYazM5
bspCAgCRAcedchCCCGLImT+SzBPDYYTT7ZifOqmSP8k3Ioa7MmrarNybZSxCKmDD
DDEGpP5M+CDgfyd4Ah1IBZHzt0SUinbJIM8kRehqjDkuD0nh1tRxGVbn2vlDfHqr
BYTPd17BtTLyeJfGUWIDQlSQB2Ozo4OGQ8MFxQTp3IdPkxaupVw3dCqkgDcs9SgN
jI6Kopqu6BRWshHGxBWO5tL5lMoelXQEC4mmgcqivAL4Fp7vblvysT0M03YrkRSd
rj+X+lqn6/QbVvyJBQOgr2vJC9Ok7X6RNNtANEDu2Z3i9o/c89ipM/v/odKH6Wsg
t1BeCRTUhjxin5nCv17S6KFY4l6YoO5fJvfHm2kjA+LPFxbG6eoDfxd/7a9UzRxa
lAMsLBSCSnCnhh9TXBjHdgToSpLMKzRopPkz1Bxla6E5mHhEVVbOefxNpEB5/Y/o
liPhmpny8MOADmPn9cnPOaen/GhCWtOH0Y8scYdtThCEf6dyN7n59pHctXBTSO7n
iTWqZmmPUHNonNa2PNFY7gyTuia2eyBikma4RI98tBMGJkpA0n/6A8XwVHrxt2hB
irP/7T1aR7PTUe9XdY7zF+dd0ePRnlCV0jcZcvlnm42UM0BEYFbCVUCvdS/GejcC
2skT3IFweLG2X+fGJ+yzqzesK2ynmRW41VGC+9Y0jHwjRzmvO6xepIDqGBjU3V95
UP5Wemo6vWaFThDEwNNxXYtWEbity/QEpPFjfgXztYIs46DaqXEiKMxhypk+SFvS
W1Ks9F1OYaH1woLFl+N6AuKY8tVeRPhpRix2avOjeRGK2o1bRl+WbgIaNO5narhb
NToZAT5xAcgSbhD2Kte/l6qhO1Pp2UPM8tmEFDhBElURGt15UkUWo49hIws4Cbl2
0Ajdd13ZO0dE/MPynDSgw6lyNcC99fjXFH6ciz07qxcMWCSLMuHN7JzEnTxs632d
OYUgPyWNpals6jv78FnDhPZtmkS6YLshffJC5PtzS1P1Z/o9/BySTn+lpGwVYAjr
JRgsOS4aA48/1ux/OVfmMfP1rjaxZPMb6f/RKaCTYglMvx8by7QJFBrW6dJdwOF7
rNPa63E8kuVCoAc1I+NMQ22JxLgLFxc5OQS3UxP0ZbzSlF7HmW56w9jwx6w76EAu
iFNgVI93LS9QjAVBjZAb+/ZjXZcl2yDkoDvlbpe0CgZrQBNSEg26hkK1pEsZO8K6
T3xUcLGts/FPOOp/xovNqMl9ae7kHafNCuhglZqhGsxb+pvPj2/5ayhp0PY1q7bA
vW3u0WCZqo0W0O4D9fwrslBk9vgkKD2bWpWoie0R8BYPRyh0lUwGToUncp8chRh1
u9QaPUq8IqGrS5eAYf56DxPCMNZeCk7Mo1XGKb4lWUoecMy4ODWApyWoch0l8j+K
8M+avD39m7KY64bXxh4GeggSaGthNqNXT+dlCLsTC1iXNip9fzh7uWPOsG5BXGJK
cp/s5XpFR4hVo0LA8ymLHTRhGQFT+DwDMv3Wh0zWui5VDIDgxv0eFyRuU+wQ97Nd
nKnSA6224KPYQZLaHw2eqfSLraengLT891SlPRi8dhwGr7XcsAqcGm75Cf+0bM+n
wPG2ng7bNv+E39zR+YSh1HfLHYQOOUq421SjNuOlznIcl3e6b4d0PgqawxHGQYDT
PQnvFBEA8l6aZjGzQhrXX98sHPl8RhlVL6OjaOJYBJbNQsOkCCKKYP9Qc6hh/ZIo
3phmXCKj/DuPgzYz8udjhMg1PKPi9UcnnPDN3emfrj4NzKxk+vvxfVa0T0/jX1ch
dcE4hcaBTdXS96wdNDGO7zqmpZzC19+e1AHuiSl9QIDAApsBEmNVQ2l8nmBCVpmH
qqLRPewEpEpW0F1olX8kmlTHRIU+e7m/Fsq6e4d9IN6j8KVURK4Q2FD68VCsKpfe
bjUNWRLDeGZcJIUaxiqG3oMSK/GlUH6qYoBE9LZsg4F98ieJLf6X2LZJKheoE1L4
E+0463yN5XsIpTziKZJl8NwYMR5E4266B3ArtW7QICFI27NaE28Ug/ZDlYHc2vMA
1nbYZ831MnPqHiKfASlHYTj4RNVZSiPQygeWN3xAOjuXnDDsVxN7gbYdt5ThoYAU
Yds5CVrqjKzEaA4Cwn2Dyv4naKG0asPmpQ1KOR3am119aoAfBDtOPoQos31lUBNT
DQSwCfq95UqPTJSQJg+ED9dsPRYtTto1NRH1lXDexuNb/AqlVGlZb/w3RIPGxpFG
vo+whWnYSXTLQOZvFRByLnbGcfbBVOkfV+xtsJVfukig0widYhpFk1grAbR9nxhh
0wGL3x3Fs+P1ffcqcKSgYXMxKEZWQ68SVCl+bmOtuBL7HfbY4Hs023OxMDYOyeKz
WtQwzuWQHwR3WIhL3jDWoReOauphywVG0B4wt5k40/JV5TmveWsArgkuTMD70fSb
mOgEq5T1T4KX9WOogmk4ZqtKfl0w2YxnMdC5jIuYzcqBkEaLXvD8Mf79Cx6uKQex
REKYZy1tF6RyScnP63oFQOKRSPYLMhveIRMFdMrFSiIe0h+ivXUdmcOOyBcp9XAc
szjEJIAhHKYtgujuOrbWSHx+I/tDR1k7a19NcxFHCyQj+4iCT8tUmybbT8w2FDEA
Yji4ki0X8EgT4XPj9bmBLiK9mcyJ+f4mgl0pkL0FSy7uAfIOTYKiBQSkNiQoQRzY
8nPdLLk62S39t92RLC5Elf1pZ5bofcfltCFwufS/P2kT4a+oVzfF/sm62yJn5eNw
Q0mTokAK0TA7fhlwP/eD9SJj9PmDObZNS2xDJaHCXn0K3G6xNYXNIwNmLWq1QZIe
cY97lJ0uezUvF6Fbr8sFo7NaaymgYmkOBSLco4RIUY1NBezIfZ+DZQ1LtWpKro7U
AOpXApWIH+I552L2zwcy2MWS9LRGI8v9MBuzkpfy84kG5Zyfg5LlqCkriwJUDrPz
hUZ7DypG6p1eaqTKmbh5JpxMUrBYDx0VPtP+vB07OTEG43sai6+BZ3SOYvUo5/Au
DR16dv+XNUPpYAHE7OhEfwOozCiqehh9YRyLTpn0/b4vRzIMxwVJDjwLEKhbAj91
g4bbUf2Da//Pd5EZe8zeMNr4LcLr/xfTe9KrJcUnTzcELI7sZKboeeE8xtpKYY4d
ldhL8tZTMUKt7IE/91+ah08s+Hlii5sZstYHT8Y3HoZZyrus916uln9ktWsBPKlj
NFdbGQ2Pbp4OlG3QIWut6JSmgAgDGIPqIQ/9afOI4lEkzE/fwRmW4CJcybf7yc6U
Xxg9fU6D3lv/KQbzYy18+Wof05RiRG/+56Y+jzKhptjYf4MQIWwiH1aTJH8eUmJM
QNNDTNmEa4l/UtnCzp8MfYu1e6dt76+BLLL3UABHZP/8O/3UhovGYCwT2LcNqNsE
8lhY1+ZVBU8AeJVAc0jfkuYZRmRgFoK4GsrA5kRs+h2X5DsPmHGa4dnELi5SrDHj
5ge8pZfYR22kAMeYVKPLqadopLXzj0zMEBfTpvQ/rNvDyCRzJ0b0At0JFMdiwWwx
FjDBEG23yS2SFBeKHJX2znqmysb09a6wOl2qqdhD1THQ+9AME8u3TiokrSoBAO+r
bdMI0dtfGkra1o1b5wOLyHvBui+ZwwMX+WND1h3SzV5ihE9ez9E72OIv4NLP9LZm
dBk/LYqK/vBq/X2glawoWbmpwO5AmW2aeLggBDfsX8SXKOLiSbddAVvJ7mcblOjG
X9O2xqDM759rMV92BawheHbjdQ7pdPkUj6BOzHKcLBf499YRaJy+MPkOivRui03w
nhNcasmVZiviqaPSZX4D7/6r7H1a6DXRZIMfwRFgiXyH+yqljubhNPnVhXBIL3EE
0f39iiCBEyCA6WIZW4/zYIlo11npCSi2lRGPUQOZ9F6h4qbO5hkwKsevjYTfmjFI
iYMFU7P0e3G9xTXUUFq0cXpw1ZicTmddsGZtalXEfNo9adBIUPZWWmnjlVs5h2ep
o7oO5ikRN3rrQLLAcY8WtRRFEUacMnrNNDoLOpNsZ3nqAsiMP9PkkRfDyb5HvgHt
DAFH1HB2po0DaIOKC63Y9+koRr/mjbkx4kDj5EN13CsEsO3hNp/2N1/7lEhJe9gH
MiE+4JjO+TWeew8AL3RMCB+UgqrZ4YPfA3opFXPamXYqa6fIkh8KQRmgB3LIVLD5
jc2yhzdeJYScAHs7bDMcA9gwyf8XLLd9d4yx6hVY4DTUtRcmitOpwNliEO8P5N5e
xVMkYJ9Lo4T0ltwqgcX36GYNOZDFPS+rluYDWqg7kYbkHBi34cCxaBpSMNui1EIB
ijGL1gJoQERtyr4/YO2hzpIZXCNM1vXdMGrrgVV0L/BtSYGsgih9VXP3SggcURtO
xNaAH11yA6XUmrigO/WbGRGDNlTXemIfF/aPTgmPvUF3cPwLTpCzjzGKPjbmUJTJ
Xy6r0bbrbJysPf6Us0fjqoo068q076QDTd6A4yFDP3burVOaPeT0dIISORzMgWSz
tjTe9RgQk3eyvjRtOdfmXTz5ZQlZaRMp5KEXeyT2MjlD+jBrcL/lR94Q6FpOVM3Q
9xwHsXo0hdaFKDGHJob3aosXx+D00az9IsQ5JO7Ap9fhvhIWFiXB8LeEpif4ySiP
u9E6NjHJDar9osvKGM4k1dpoiWuwW0o7dxbaZ88uP27sVA/1sLPwaj40F3LRTX/d
9JkL3YWmXTSGuIPUi+pZ0mkWW1bQsy0epurlckZix6LzUT0PY/KS/OprPtqm9ToU
ZNHsYrenP7XDYsrVtvVgAHM0foHDGhd0jd2UhmXnTNLOn7iwlg1vpy7gmRYPpW+F
jeIw34MgOoXE9YUO8/v/2QSUBVraa3l+LMerhC0i2P8MYu6x46fX+bqrKoHZglGo
R6oyFIfeGAHOclRYm+nfjr9PxJ0UsTz+leTG+rjLZe7CTTJ9XIhHwSMw3eBmt9NQ
GPh8l6XF+b1fwasltxbrr5U7xzRwsn7SC/+Ooes4lnD4XElLyHlG49zUcNEgHFIi
I1RwDLm3YCiNRhBbBbydkl8/b2aByiZBtlFOvbJYc9yLbg9nxT2coApQe7u6Q5YF
bmEWsTFab+VTvLLdsQ09Tyb/9vUBLK8MKu7vp4oVr3xbsjt4fDerMKXqnyOEHuIP
PSrexFVT5YaQaBXFsmcbd3YAB46m+CMIlB6La34Ko0IhWnRLcMI6/S79ID5Qb3JP
PUSL5hxMY+OQ0sgNtGD02hmEW9OB5S7E3FffwZFlBTZ4EMSeC1zx7uIu5dOXUoL9
C/EbZGFkdRzJ4wJIqLnf9uPiPNqGDdetehF2na/UCaeem79OfeWgSzD49WofEVI6
pKG/R74t8cyWilqNo9Mo87trwqMOcjEu68KlHCHTxieLqoG3aFhBnm7eJbC4vLZ9
MeBaVpOKeZxmb2qMY36nIqwa/L0/uYgeBBqX/mXonp+3qIzodfFu9Inn5vOs688F
YyRHbkI34hTozxcafiqCB0XeUonREcgEQ31X2MjRzR5PsOQUf1emVZds4AMdOsR/
HtXripVg/dv8E+o3v35gIzxrMq+zAnbm4ifVSpgMswY194dvqDc5MC2Boeb/JW/j
4OS4Wf10QKAPIJ4V1Lk8msU5gB/Fb0XdSchCNcqcbA+j1VtsT4HudOA/xD6Q4eZI
odbcQMomGJ0mwQof43je4G8+ufQtJq1t+teFsqmzoh8+6TyojTQSexCBqZdOfiDl
HgyEIoo1hhy6m1VAzVRzqR3Bf1RPceDWUUwm+xWGcHoLNm23itE7hsBi5zDcUabs
eOBwTMx86M6NY4UccU2r/ccKSEN34XSvRNC0SMGEbVd4EkOmBdzIoOQof09KWxRk
KhbKmJYyiOaO2PFUIVZ/6KEpr0tcCrPbDZg84OboIjVkM+u7othWKiVA1WUFNcYX
AmFbTh+qUI6nUz2T6DiHZ5GYABV+LO7pUs9zCjBA3j/o6CLpO2DUnpUU0ARsgP/S
R4QFo2aXEBr5JgBmNnqYWhAd0pfe0SFeKZRfXiPs+C5NgZtdDk0pPc3tK1Ox6nov
/IFsYGCStqm0xb0OL7x2kb1hWMnml4F0usMa5WmGxDvw411PrjTcXAEI0wnTKTCc
4ut6v2yri8ycw1Li/021oTGMB1oZrHeHGRgP3w2RvVLSoCZWveENisOMJOeqpDYq
D63/iUgiBcBJjLdRxKosTbrGpsUfIVwdGv3Fuc9drjsqgAvgWFuKFragPbdpo5mK
Fg68mJAlAtlxe+yhCfd1qHprrBMCaO8mTYOgTc+3d0PvWFSXa7Nw0dJq/XxXbMz+
l5k5FFeaUEIaDzOQS33mSax3TN5mLaI9+oqiE6bJiahUvfbnagSWRGWkRWBhUdFi
hZj1txVRHJf20SMXg7Cw2PCJ+TdEzVwTNCWH/qJv9/VCNLc6wd1ka8JYs6nnni1L
N95NKuxTnw4XVjZKSuJxKakbwRgssZRJDINR2iF+0QRciBbAvl25SCzzllFYG9Xz
HmVjvMJBZMR1xu0KZkV/x+BpVlStKtcduzhfnwPofbn3bl6Q/j+J8VRbq/lZstKf
QhLiZ+S5mUx9u6drzLUYlYuHXWmzZf/f5yOE9fv+jxbEPyt6wCR0YWlIGm+suAvc
1NbjZXSj4d9We01PyK9gKJ/ZbIwIbxFC8B1R5Z7OAMfsqv2iGMIZvUr8SVZAfG9w
Hzl/alVQIQF87nNit9IqdgWe8RYDoxCeBm/cp0TC5KZ3TxENz58zwxnsTkFbEJ3a
lrOBCpJVmrctpyyvk2OjNp2Srq4mPtybNv/muG5jPFHsY2Du8gLZvUVgf3CELkJk
5z1YcwK8q97as04mQ2MUAYg//BzJqudF8WvVNfNR9O7Xtzv9tv1BWkmd79vo6tAE
vcoheogL32Es95912HMQapbflk/gKY4r8yaQj9CmW38j3kUY9ANtTGw1vCn/G/MX
CCxm85ei18Ckjfwjyo2ku0qXyFmdjqpXtmwuri1yDbDyii6Ihq3zuUzFSIKsRgXV
MCJbAmDL+fLUsl9PoAi3XL0Hop9PjTjBycl77IXgpb/CsFDxbzAhfhNvldHQwUTH
St0hNXslk1/fW6jjbAg28/8IZKQs74L6/9fFSTVc7G6hhYHsxf+nSMKHeVt4XrVu
KwHHPFlJjyyi8HPgscAqN8enLXFAkO3bCkT1qDhxnlnpp0lpxLAlRqdvQPkQrQiz
hOnQRhNCri+/bBCbvwa5TUUI2CSMQkx0d1F+h0FWVOpK/3hha3c/0/8riD7xOgkB
tD2erGHx/9OCa0YB8YMiSsGZmNkO5g2E8c1rslIflLINkFP5vmMB8q3rW6l5+Cmb
e3xFJHI33BgrH9oAxmyyis16xNaQypYtiUuEYXs51JcviXwwzd5/X0iP+MksdItL
XFLxnDtHUF4H5gS/kx3nuDEDQwmuqaY5UKF0/3PNEDohhaRcptgT3e5JfXsM6DN0
74LfKDefDJU37OmRd0zETRTkQLfmOS4uJywb4be96rYPzuLl4lOZZ0tRRATK0GFq
jVXIDY6bo9EotjnaGvF2vkF4l3sHj2KpAy2vT04b2pq2UyIjqIkVPZz5qq5vugEg
2hHDTDA/WWZlAAEnU4FqPhI4zRsUx64mQr0ruL5nMc+jdodkAs2rCJ+7NYgNB7X6
E2fXgtsxcznn/YlW6mkCB+mOqRK38tSxJAlkV7X64wr7nX7WJBf4YW48Jf9IqW+U
loq5h4I+ydBYMS0Wk/bTwIPzS3fEmEpkaRSV8/uN7dZ/kdZCT4TfHSzxaQmO78Nz
icUJ/jVDlgdY+7tt3fF0NxHBEDJEcTFuWzw8Jcy64mdcP6E4ZBa//Y19OXYTJ5iU
eMHbfisaFCp74BZPJDrBndOtSDDLzW+bIll3qEnldkUcbHUf1yTL2oHmQojfDm4a
+0lls6PFJ5ABDWk25aGRDR4f9RkavMzmDkQGqcals3V+m36td71Ttj1N0T7twYBA
krmdqf3OkXGvRn55mtJU2V7kP8M5rEzWK7yVzgDtG/0s5iM2K0CwTEiYzN6OGqEt
WItbj1IJa2IDpWJ76nVtrjn/CbTYWXK29/CVJ5vHkyBWz4Hns78WMAxYAM7XVZGJ
pixbWd4RvYGeBVvJjPpc7kEI5qk5GxyCUZwbj00tb9YgK+UIYMYVk1f/XDV5fFQ9
Jv7mNBVCEsQyUJubTgPWKfj47wSf7aY5oTy/tzu2QxO2NgSs/FvNdYJsHawuygNM
IYE+DKV+9JnoFR4nbmODoyHqadXcWx0pL8+N4+IrL3qfk+FIPvibaYuzWoL1mrrY
fP/hefKe1/ktqD+5XOsMFpEhs/l2GznTr4d2wHG4mGtGLJVCclnvfQpmQuFQsimi
wOlqCXhOr/RUxOrYJHf0gJF4Y8cGfQAraqRv4RYu0VIMLu4jvBItZx1Uw02x3FMJ
4cLwxlDg2RIT6QXDT/LK8x4hVFZEbDWNpj8HJnHzHJI36+91xFMH0S97sbQFGtIS
H8bXAMs+q+0EB+bNbs1pP2hjHD2cki1jD9p8jVIWK61QHdEUKL1vD/Uj6A5kHdbc
JxNss8iFCKtvdfcmXIJCJFCtLJd531hEjt7wSVucXMA02llDJfTBftt2Ww3gUkLG
5TwgJLHi3TmaaRdy0I0RlVSmLjrOBFL05BenyoxuR47zeleOXLonPGp4ziiyTB9B
0cpIBnXdkDp6t6H7FUxLpJkqPKsyB7cGlZd2Qo+ecvoVcuwuL6dV0DH/RqgTkojV
iWytuWweJizjMIhvYrloJjFDyHyu64qSSK+dO0Z972MLk4BdSFPDSDcCuid/1zv4
g5pSH5ZHsf7axsF4eYlbSsgXldNkx3x9aVckZQw238b53VYGBHBR3oEHBWNt2XYC
7MVfuDutUQlhJglmzEVmrSEJGUQr6yA4lUry8vE5obQfzEpJgzarpd9WyLMCvqx8
LhK99qFc4aCZJL2JydBapQhNDy4CCMp1TiYDjKYe50f1Pf2kisH7fFUQzFqgFf1S
OSSsZFUL2zLy4yoqNFgLtDBlrm81r4izTfEHAL/x5KZj8ldvbkMbkGN9X1OPujwT
0+CTzAOW4BnPr3CF8BAgw6cM4tN735TyssVODvm2rSIKmhPTcQe0m8CGxZ5x2fQf
dvTX99dQad7uwAXtQa+Q6ploP7ljJriWc2nsTgX3uLRxkD65wqo777/8Qwvk49yj
9eebaWcqFLlwc3+b6O7ZEck+gFpGgqeCAqMYIQ+eu+fsaW9Dby30ps9/N816PpGw
HmLZpO90UfzjSFVVPLVSl5dT/h4+qmyWgX6NXuRfUv9DnFvAdzAzVRAOP7sta7BE
mWAq245c1/nrCI52wZtWPGVQrK1WEGwgN09l5nWqFvo/SbVk8wpa0ckFjcZyN4kk
063jif73XMljL5l5tkD9d0GplT7O7a8Q9sE1kHQI9E2dz/PCImEYY7nA6o6MiV4e
f7hfeeSVWCIYN6ceoMhOQE9h09GRrsIcnivTUIqUQ2sGSVZ8FyT3yNH0NtdNCVmn
3FDMi9pCibfEg6jG2awHyqbAxYKfsSELA9xU17WP7bwSmrJz6mATj2dU8hsrTIvz
dmZCP9pUQ0ak1DOVOyDrcjIbMR5wbpXbRq+QVkUIOJ5Hz8cbiqjYaLB83IF1XDpE
d/4AO+JJsjICXiBIfzdgJX07WujH+L4Mdyjoj8cAMrWdIfIwrkfT02xUpkVvrtj8
9WI9Aw2+1Pr0ROouszYGPx/3UgZjQOu3dcStGCULPaW82YGkKfJAVSJZQvfQGm/l
7f4J9CtrOFba4EYGFAmce1t577NsySuztFQrOiaTBu/U42k4zvZdXWlb+Is3IZUj
9nZXKJPqmZ5fX8I1ljBTDlor0uXB2Krn3x7DLBSNAsVlhG1otlsajOk35AXI2L92
srHTT2vXADVt9Mt+FsSTSy/87WCsM3oTvbeIgBjcqatJpo79iRvRzck0ylkBoRS1
wmcSL/pvXj9jfqQu0fewkayjDbELzWvHFmQGwwJ5/AtpkQKtV206mm5ZPwPpEhTY
TqQJtqZRNUdJul+FDercXchKq5zXRJFp+4qF2AxWLhHk/XWkeO1W6zDXs2uiIvOa
WEDhRG8nhkV6WaEF8AGs55cgsYHXq58WyXncRfuby5+qXcNbn9tzTMqIIi7Q1v2X
L6YOdXvRs3EL3KAJYRXYblw3C6C7xM+ZImjtYQ2gikZ6ZR+urchEHS/uwoBhvXUO
/gh1jZMlCwowAFFOkoQV/gSksbmoQGK+NRT+1kTilgYEkP7qr4kqiQ9hBweVZ6d9
LXQh/gBfftOAS8DtghWYoaKvkrB7WsgEaHhv1BLrFB1/8MiFedw7SHFbp8ARjT2L
vO5XZIKCJ7hqO+Bws0VQpR9O7nBzuKkUCYmzLzxo/+OVFUlMCUclFaTsin05VIxj
LC/eJVdbx/Imx92XoDb0gxOZCPEuSXXQ8fPy/HYb5C2gO5ZjTgERyNNzTP08pri4
EHi1iurtkODgXOXWIagl/Lgj4LcyzYBfuGHpa/b3GRo34rh7FIiMxk0RxVI4QGB9
r8w+tLJz33/VCAnHXjQnXgmSzlIWHJhOSSYEMlVS6g2gY5Zdf7s+xPQG9svzWFoQ
QQTCijqZ6ie+GbVMuvv12+UqSPtQsjHmZftKVBgpmClgl9C9tSYYvckLMDBtjZ99
ks7z8eRGcgFf15iVuv0FwYqgrQngpUk/mkEMD2YobTbT+lgZkBZriGLB/Cg7ftoI
rKlKDsIa+mOyOCeavPWpZOaioDJT/sK3dGtFmF5F6QlyC8wJ3Tervu8DnKzmaQe8
4k71+JKsiAo6fsjr/fv2wBwXJJHEG08dkpKo0vji7X8JRID0rZop4y4zO0x7tRa+
cVwmSjpWOjTOLLjWpeklPfp5a934Q8X59fPgxCdT1xMCpu+m/6LFHPa7dfvcn09j
9ZxCOxwk4FPGxrSMy5BaK8TP0iHY7/0xVPUq1EKwXeAdDmG1OgJVm5Cb+U/tIZYO
gKi4geXtwKdtTqMkSLH0ZiXMJ0KuGqCfr6vHWX0TPLiIDJ+fb/KUOfJaCbDJhcUa
XS+X4JwjFRIxX6tfknKboPDzE0Vcqu0yEMB16gr9461MTysR7Ry33esZ71NQBem5
0FHWZoF3J3XF0AeunQBtosRLwLnxSu3pAu0yuVXdbJAMIHukXPRdjlwFIIPaRC2Y
LMrkwetEahSXUYJeUzL8MZTaOSFBbtS7PXRrvDFKqlvJdRXzAlsKX8XZJ72sk+LK
LsdIUOnosio41tQ1/CVWLi9DNz6v/9P0n/cfiuo7kr/EqrJ6TvNU5wEBZ9CXke75
qKvGjDp8Q0UrFsPwGDZ/j+HFMEaPeKfPRVEOn5JLbLy8ibLHt+YRh5SH3p9t91Sc
2PHvyWQMIjlfn5C/VfCzEgwwut1TJKyC3owVb1yAF+mYCUAwsyT18mTMEFs1xDmQ
WK+6MDIfawF4/7I6IPApTm1ZzupXxez8iVnBCrMXgn2xj8Hg/lwIDNmwx9Ld0aWL
paFidPoan0qw4h36J6X9NpgAYXZfcrnrm68gftIPkTwhBI3fjjgdx3AdORm2EI/W
R7+9njhwCjUOMcbzLjKDCzkbSCSE7MrApVYKiyotnsuBb2jhGt8Q+KbSenswVyMN
xh4L44yAg9nrMxt2xNPeZFkNbCbvXU9Iepy//K/GppqAlcR/wwLfdRRMTTXqT9Fm
gBHx6UGjo8KTO8n8J8LIVDsAwPJxjmpMPA0GlsjSROhC9Cci5nD/37EC89dEAQgY
WNTVxW1IkJceC6B6fR1fjl5IwKN8gWqOr3/YLKAQ0NSybpDuL7oSLqZrE22sk5Jw
Fwb1ZbzR2mmxvZi0MXV0ekzZ2Nv74ErNwGOkC1/CBSiZxIBitA1wXIXGI85UW2iv
c9gE8HMk3nPcIGPGr6qlZ3c6WfdfkjhMrHPSTNqsNaEZHI0Q4OJHpmY7lH1qK7ZK
ICUvXq06kteG35xZdtEtp9nD681jLEAsbFoe+ijSmcSspwnBOYtE9mJraWk0rmpP
TQiTARWqAgkCzCxFEnKpXllDwywzvX0k/FWyBjfrTpP99bN6YqN1+/T5KElVNJ2h
/zMy7xkz8pWVzcYINWXgeUzVPTex9QaJsCqhvNWIrJ3JGC8FQhXByAlhdQ26WEAA
gk1kdepe65mZ83Ylkwqs4k/rtYSmFKO2GJq36HvWZeabJAMMeUJFBHRkvvs/vOcC
CZFVqDkuwjSGcxQSoXpNq5AZSFztY18fd3K5Ts+K1SyooJdTK4In3r61y/rZFy2B
`pragma protect end_protected


`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_master_transaction", svt_axi_port_configuration port_cfg_handle = null);

`else
  `svt_vmm_data_new(svt_axi_master_transaction)
    extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************
  `svt_data_member_begin(svt_axi_master_transaction)
      `svt_data_member_end(svt_axi_master_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();
`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  //----------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare ( `SVT_DATA_BASE_TYPE to, output string diff, input int kind = -1 );
`endif

`ifdef SVT_VMM_TECHNOLOGY

  //----------------------------------------------------------------------------
  /**
   * Allocates a new object of type svt_axi_master_transaction.
   */
  extern virtual function vmm_data do_allocate ();
   
  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);
  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0] bytes[], input int unsigned  offset = 0, input int len = -1, input int kind = -1);
`endif // SVT_UVM_TECHNOLOGY


  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);

// ---------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
  extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
  extern virtual function svt_pattern allocate_xml_pattern();

//---------------------------------------------------------------------------------

  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
 extern virtual function svt_pattern do_allocate_pattern ();
  
  /** 
   * Does a basic validation of this transaction object 
   */
  extern virtual function bit do_is_valid (bit silent = 0, int kind = RELEVANT);
//-------------------------------------------------------------------------------

  `ifdef SVT_AXI_QVN_ENABLE
  /**
    * Returns index of qos_upgrade_delay queue which matches with
    * current cycle number provided. If it doesn't match then this
    * function returns -1, indicating current cycle is not suitable
    * to upgrade QOS value. 
    * If there is a match that means current cycle is suitable to
    * upgrade QOS value.
    */
  //extern virtual function int qvn_qos_upgrade_index(int cycle_num);

  `endif

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Wtwj/Mv816ki8DADc7GtBdznwRj4li4XF5pJR7u28wBfWyvOFY72xSC+KiR9C5vq
rTf6ZreGtJeuv8K4BGfAo9dfoO4prjIBE4mU0u+8DsTSp9K4abg69XqdFTuBqKU8
aONxjlIu3OJgm2X8iuryBgawWMSYPZvSNgXmY4+EIzU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 90172     )
mEAd/LVmzCZG9axMAk44hADYM3WIBKBIBZtVq7MwchmHfbLmPVg6Sgu6otzW0aL7
Bxel09zDbJQGGZp+ssLiqnahtd/9zWxWDN0/Xps7+TCB0Gfxk7RYwaQ7KcEx+C9W
c4wtEkI+F2QqAt0ZJbo7CX8OU/DOPTGidzedysOWk3Y=
`pragma protect end_protected
`ifdef SVT_VMM_TECHNOLOGY
     `vmm_class_factory(svt_axi_master_transaction)      
`endif   
endclass

/**
Utility methods definition of  svt_axi_master_transaction class
*/


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
V1ObQ5cPBs+r76VkuWqZPafwCI0r1ObDxd8Q7eID+GlqQTEFGCG+Ps3LV/6+VR/C
mdcUXv8hR0+UkB+NRmBvqlhqclpUbbIFqH1iqjsrMgHO/yO1Fc6oYHJTHQFAdslv
vO+au7Yc4g5v8x0tfbHzqep3Pt/pk0xbPqW1GEFbBD8=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 91965     )
8cQfDWU53quNL+pP3klnj2preiONsHBgUFdowCdlJxU+xYulBbOcb4AUo/ijpS4y
iDCaygYzaWbsWWJh838EIukJiOejV6N59/wSujooddRfGOwTgX0EriVtHu/gN504
R1WRch8f9ZFuArKJ9plZqY7Gp+Y5ed86iyuuDZZ3Tw2xiyzME/KEFz/QPVw/JA6K
5GPnOesncnciz4xK8P7JlH/mDLHnDP98DxecEmurjxRWlrTXYVss8nT3tKEE2BSp
SwV5aDHhHxsOX+6hkB0aOaG3tk+DHw1Qgv1sOetzARIBo27CpRLaDlo3DAA8gBUT
w8n4eWcmeE/hL3r6CdO3j9/RUZrN7wPDuPwUxWiwgPfl8qcTzgrkyFfAfs3HeOfn
Dl5W3mwgPOHPaG1JAVJRkSm9LTUT3QdM1AfXgGYBvTJqWMwcy8thhaEaCf9lSIQS
RMZJs7pggkyuK5kaVvJC13lQge+IF2PotqTfx7pMpCUpyoyCY790COB/kS4BWWUu
/hlPYBfjU25GyGJKk5KfQI33nEbDFC08z/PNHeTB8wg0vjsHdWE2j0OvfvYRvfIg
dez9HkRvG9/zp+Jzw6tkGPPrwp2BUrjOhvQEkE9qQJiRbx4GMNGlsbSlmGv8yeaQ
rdgm/TmTeEDtnpKcZtgoguPJCj6l0Iic2iXasulMINnhzpkgnlc0Mzmhtlm99+Pv
zxbtDPiXlYaxv5KgFK6kZaBBg2XHf9/jmk3zdnkQ/4DYUYyp2ud8+K6vcUziuMxy
xDX2GSaaFtU65EBNBJQn2/8ip/5+0DjT6ZMwZWYyTxuuIz8jccEiu2FlJ0o3bFmH
ZlDKCqsDsbQ4V37HS2a04q2nw6yT8K9JcLU9QTLmMdBF2KUlFZNIvUwPkZPkFApt
PzDC79HAaX5d8vGbYiATb9bfgSvPpvIAQ2v9ZKsGz6/LhSM/mvu+GX91V6r+clNl
xxC1HQ/c0pr/to3be958n9lECuYldiPK58pqUfYdtLHP1GKj+0VPlhyqxh4zPirD
TZlcaD8awyPQFnGSSxcEPONJusryTPcQLugfV/0ltwv6OnZ2kTfQeKtIrSGnnmH2
w2Wzbw5NTRuvaWgul6+9DjW/4s10o81tIwd6qo0t7l5Z8DgqsqPdmejJhdqoyqBe
F7SSk/Q08iNqSb+a/OmeMqAAhjzg6r2mFR+NFc8x9C1qkye8CaWFn72NdBb0kn52
XzyYyqwVfNq2zn8H71YTYNqRf5SvRfi0dhR4YOOSlvnp3x3JBw+ggwx73Gjj7qv6
t+nLiZsSKiZCa7J3SrXAtL92G4Y4wGohkoq6SFO0bKM9XKnUfmD45P20z35IWroh
Pun3jVZwuJQP9m1jnN97Wk3fL3qu0DJRBG4itWMpHMnYE/rwX21fWT14jaCrfDRO
xxNgF/ssC6Q5lhIwDe3dT4N68TeGJAC3PqsUyhHLFvJVnsmBxQG3twNl3yn8MrVz
X9QVlJohbv9nqiSIvgOyngiJcrDwK49y/SJxxg4Kan0fqiWQKWQQqrYAgIV7BqMA
qf632iefW36d+2Goa9nDO5Ar6gkFwNyT1Y60VOwGXgEl/oczdTc70iCigMfYe10y
vyfpar+g0xrphOZBNl3KfNKYKrhSFZlZcLUjgMgDvevdmb9vn9aqp3Kch1iZyc1S
4NwIw3HLPuelrNRb0KRMGxVd+BGw5pWC5nnhSmt4KkY5kpHAu005sQryonWPYa8+
wTr8HPT5/32gQCAcG1CvU/0VYEg5nbUwDmQTy42AsPQ5B5QzJ4fG9zK2pkvjWcxe
bu57NpDLCijeG7rOVMDuNPAsUIFx4T1YodebfgpnFQSDzENgKIspTT/CZXcI+0SI
xPSM7Hym/BDHk40mcTvfmrMQsU+9VRQSu/W+5d3ZQfqCfyDhtah7Ekl9QlidAyso
M3oCSQST28+WAvo7q5gnhwGoBCTMefscqV3i9HMB64xoS35QgBI3W0EJRSZv6xzc
DMS9bodWlV3LjQiv+Wcu3Xw0DiiwyaM8g7yBJd1qCUgpuJ7wd1BN+rCvhVJmlSuJ
slErMIUxYvb3kt/tYWvjHc8W7nAl7L+QkCI/YTrXopK+kNZE+6CoccvMNH56KoQV
Zwt/h4w1IEwDIr+Tdww6zzqJcMUFb0j211SDGfdemd9VSRi0tex4qZi6xE2sbAZg
VlRRiGOJZbZpov4BtsXTlgW0aCjmNMn8dNYCBEKCSfD/2sMeuYSGCR6z0w8L03/7
MyIA/oK9EiFUDshwb/GW9Iq36SBdWghGN0awzlnFXI0fRXvcqyeVPbk+xdryHiSq
yuJ144aOnll0n3blE3T5XDD+rXrOtHamI2PR6yuz5s48bZRGYSMn9tD82VHVEuCO
wwlws/cAWhIS/hUVRxkGNbK08JYmlgXTy7wOiOXdtgo=
`pragma protect end_protected

function void svt_axi_master_transaction::pre_randomize ();
`pragma protect begin_protected    
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
kkT3dXt+4fYKWhYNhBNvxfdz2fxrbLKDmmRfDV0CeT+5RPYCjqe46O0HBWsW6nS/
2GzvgiRzNzJLDSJ5ojI+TlPR+HnoZFEg24LcOywMf2SifAJ6G+90JNGFNx11Nxle
dV7ACuqjjZA7C19L/Be5SphM3kh1Zei73pQaF5sS0lk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 94442     )
HIwSWinddZaB26woC7xt//4hdIhpXeD8tzTMysShpKLpCeJeimARZvQhArKBSrdt
aVoK1Z9C2HogP4uK9wTep9GQbhtF+kAMuaPIym+wqRmf5eRDy4sffP0dvsG2PiQ0
JlEjbRGW+ZHJCizSecUHocDMWogwtIHIfx1SBE6ie1iWh86gIcpzB/pjvQf9cTxq
Tr/gk7zNZ+JX4NKrp3GL+msiokQtpJAQddCID6noRdYyNQ1dek/VlUfvL4udMWT5
h4mBb4hC16SpLASiDqxXdQ7UyQ/QXp3kFmh6rBfD2clu/JfJLe9/mZWcJTWUHx9C
F92R06HSwoD9LJczTtBL/srXVdOz2DM7LtDsiNsYz8+x44FsB4dSDcLnDGkzZ+vb
fPrM8AsW5NLGW4ha49qxTX6VSMLrO1nEAPDhpW/WS8Bktr9bnXycPUty/3+Fiutv
ucmEwlFcRp3FWOMZu+6IVobTwumFIjAGEqgx5hM9i7t+kyH/13IOx97HxAy7Fd6h
JxUqjHTwio8r7SmJB9V3BqbjEM1JeOiUsbIDRYX6IFpfxkHn87RSsdrqUl0djBgC
689meTZjE5Jghjd4uXA4X+KmiSXxTd8plVP1rW0+8QiIg1gkqRT8bNQEcABrUpNz
23yeVQL9rDL0lE4uZx1IKVUXVhDF9uhQE9e1Du5JqLInaUAsNxcJiflu2XzNzCxh
4terreLBzjApkWsvwmCL2m29PBR60JrQRh7CNNvtVZIEmtRH2KsSC6kqlgOrIZAF
/9/ww1bj9PDx/2+XAeLjzT0EApu4FSaTayNrpzFhUmVr0gRTsnSN/kurrHlkugmP
JOmEvRFcFl0k151Xcz1o/vpdomeOpAvzqigIr5tiusJLOxIOt+GkQPLd9lS1r3fJ
T6XGh6nQgUu2oJda3R2U2U5rhC86LSin9Oq9elCqQV6MyT0RIfpn4kTYp4QGbG6Z
AVM1XI45KRAoBEcjuT7tL6e1RBwablvC1oC+mPy+AcNFSv3Cj06OuiJLvrDTrHZv
3Qo289FOuCLeFd+6aTDYjw2VbAKORo+KhJ2JgatNXcmQ9GDtMUOXIBVVSpKoSou+
fOtW+hXjvBUtvzyVtK5+7EplQ1H9uTyUMx7ALATYpsJyAtpzYnDRL7RhW0tsIKrg
zLnxKFHuvfvgCOKLZzAmxXV0zGLe0Yxy6aymWKBFgF/B1MhD7vegwPs+S3P2XpfH
XIf9zELQxSp/aqesrK0nsujuaWYMRxAb+knC9H8n227v5O4NSBFCTwKpcO8md0jJ
GlD+kPtgZIasxT19QltfQYSqUBdupChcC5XDvQ69SXE3cQqAEHUG5S0g635aC5r3
qZK1l14vU3Co0RbH20UxUnxMlMwwQB1EWz9ewWoTd9anQZs3kn9LZiK6dlv+AJI7
LPdsrWSDoPoz72r2JJOoirUYRk0pMxwtkuWRWITa/jTRmhHk33shUr2cxJYzPnqG
YrTcMZ0Wagzlp2M3MJMDrIfKdPKX8keI6n+uEBWuMxJHUKSCiSWTKvIS8zJvxTUG
xltVIT1SkSYBh65i2AIBvydTm7eO5JzTDspvqa8b1mF2IeeODf0P8H/xsJ7m17nS
wdikN1hWx71cXVHUrrTZfL9FP/uO0E5ICtnRQ66aBwqd+m7l7vup/JpEUqZ1lFl0
da9v1Oqf/0Pn8zBUobsQJInUtuVn3x+MOG64JoyoEh/fwBvE8vB74jPWAy4XntYx
ClkT2M47AXLe6Za/zUDTyGBuj3N/NeNmQE6g9EcABehvx5l9LuQtnRwfQlFm/sY/
PIJRAjwcC8LJfWTToXxUrtUUsOYN7lvE3G8aKufZ14uWwNBDFR+tx3hLwdjkOZxq
euPyFKkZXKMM/uzwURnTZcVTkmgUP4g5YTwyq6jMHN8es6QVbfaCd3X7VLwfHf4R
MAC4hlN/AmPPReq8uExI1vK4Of2yyfq2krzFdNt8AYAU+y3qLNfxSQ8owhC0+GrP
9/RyOTTUpZJkqLmJp9SyrrVUgKdUuR4SpFRw1qHY58y3F45V3GSk2LY4r4Z5+sso
qf6yC6mszgAiyjfQoU8rR1ColifPtjpthalAdzRNW5IQko3cB/SaYCqdjT4+7jys
mIX/x3uUV9mOa8gRqN6j/DyFruyyJj+dId8XDBn6hr7b8oOVoNXEgn8xJ0nPgCOO
81qyQvYVWzMJbRJV9Wslyra+yXLW0PN+CbvS1J8+3oaA9Pd7xhcmxoWFzLneMzFf
Os2g59N2anll1aaj4tGkQaRYzC+E2R5LGBPSTscKsqo51DPIA8goNpUgDntpSxq/
1TBs2SZBHqQMvc/y0PyTHzN1y1FcsIH/BgG7/EgWGvMCty7gAj6Q1pDVfDVq0g5/
YfYzM61Mxj/PGYYw4qjYAT4KxYUOsg3Uhcg9R5w5JcmRuZsprVEoqsCoc9GcniAa
rHD/mJUTlnWttn3mEtgOscLieYHh2NV2CscYhC+GQBBuoSrYpaf7K/nAjr9vaxam
OvBGe6Drbq/wh44hgLTq0nNV7f0Ev3XtG5AKIw7T/tivmvlBUVEtsS7qkhwQxjNI
acXboElxcaoOdWy5py0ykO7LAl6n0h9KuZuI4vAjc3b+4xNHrG3x3eM+rOyaNlYc
hWcf0Y3Tds81VKeGbVfc9XUfYzUDatkMwKXRsEiTy2BgIUSncJUCeG2FQIjlP2Ti
S1diU26Cj42SjHC3RxVMHzQZCLqVInK+DikMyqoP37t2L6Yz4Aon2FFakfnLonOg
irCfwTqKlXvS9EkrMJMpHk1nbYZ0wWYerizNGbFMS4RjqN0oaPxS0L8zsj54TBX0
1jxSBMk+TogzBse3J182Zxqd82XgF3sGHVNtO1bMqhwK43Xri964s946FG0s+BXH
inqQJYXMwaB8awHgzTnM8IfreawMPyud3eFU1Eyde4XdUzwSPYTKRMEkLHBRA6qq
a5CIsymIf1MonKdl1MmTCWCbGThUvaTUaP9tsMcYJI565antMiZOeyCvSS3fasdW
V8hf+6VreFCQnlael1gMCQWHixhMxnRPVnaeUOsmZK+UDt02gZuw16sdS/tCAvq9
vC5j7s/lMpUNP0aA7WM7GWe/aEYNS6z/e02CCYuKIlxTFy4UU/tgwG3mTulwGWpl
rjx3TVUCLaEjCE8njtAXGw6ezedfR+PSZ03MgrEDsH5U3HKlCXtutIQ3nv2LOXBM
BlBmFiiSaLNQ3RFq9Sve2SU3m7YtiAeGTACqnQP9sNK/RZVuwuEG2BiGTWE+xLdE
Vm6Pels5ToB1U1mUZ1GZPRuxVIT6VkhzneYIjEszkG8=
`pragma protect end_protected
endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_master_transaction::post_randomize ();
  int log_base_2_total_bytes;
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
i3GDOCbgzGH3k7lrBjROoz/Ziysci7qmf8lUSQFirYcIZNzrn9ZhsdfCRrcWSWZB
zEqYbLfdH4KxHvblpLsDXsfh3wkGj3dxzqeeYKREBW1oJcf4G8p2x6WPBR3ymQk1
opxzn4WuBb4IdKjbMqTuTBOSYfmAYaosEg0M7ih+HqU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 95190     )
jUXd5qvAkgSeB0WAzTTrrY9QgVVH4dOoYdK24dVyAT4qkeQE4LLrRwA/O8BCtJuS
6foWop7S+Evi43ghHhL4AP94lR+geIWfXDCC4kJibfwUIq4UcRa/GxNz4oSbvzbN
qJ/tWwTL7bJkux9gHFURvw8bLJMzDZjsng1Xu51nJCy6GSTdELkngE6SKBQ+fS5N
NC0wOix/efiTUlkvD7VRzO/L1qTUlvVHuDUQY+/fM5jep28UpPI7s4u2l+wWvkOz
KnY/nrXXDPJO3fXmYxC/dP/3Hd2p8nU0CsukZLtVHcJINFQXKvj25nY0OcPZlPcK
wp73kXADKrPgZZsyDqzvI67tYTYhJ8mcGMjTxwhp6upB/PrZwxgeHPoDLPipN3sG
tHmTG/RE7zrAWGRcsb5CsggDavu6mTdHAnm5W0Oa2p5GLFhxcuo3d0ngPi2dTTzO
flXOk1zCCFMC1op0bRUTiJaV5UpyH+7Ekz5mKNht5+IgfuA5q6Omku7obmgHSc6e
mk3fFg11Ck4E8lNUuFwtIG6uBc2cSuYs64jtznYjnPuyhhD136aJJL5kUmUt9lcL
s/BLJLiz3hBczVD2B15QyhMqQFYvi9OpNOxWDaHJB+h5dctg6NbkJrphIu3p0KS8
DRYYah9IZDv+y1lcz5qsGDk81azM40Tyu5nH9hqxG8Ln70mhb7NF7nvN5ikU6lzi
5EA7Nt3IEhg9Aky7VlA4lhbMdC7f1MSKaZN1gQvmNCiBEmYH+qyq/MMgXdKhcfY6
VPJg18HPq/egm1mwcWGZdT1jvP/Ybiouj+gPTC3Jfc5ogqqFprLxgOarE0wf0Hgq
O96qnnev/F2LfIpYlEF6t3PSxm//h+aaSSasWTx1Hm7aM9/SAjakwKBQ/FjrunPJ
sSGI2dLdMzbJj6I4Go54DIUfXmz/49R7RboYxwo+Avv3aefwCpWUhMTD8csHwRby
ehSdy8X7njzlNeoAWunj1t9x5L7tffgOASwzGcClPpI=
`pragma protect end_protected
endfunction: post_randomize

//vcs_vip_protect
`pragma protect begin_protected  
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
Uqth1eZB6pdKN5kA98h8/EPGymjEFLu+C+smIYBCW46Tv5Qkj+4gfARPKtEdixn4
3KrtT5RfzMFkpM2fXq0Q/9JO+0OL4kE44DGhD10Icbf4tA9aeeLfBAEp7UHVXf/w
BJQkFwpr1nFaPeCJmBE1Z7FTXZmgjFY5OKBrguM27oU=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 95817     )
gL5qylf+YblV1C8WqXsvwmbms6AOQYN9CMRFmb0PeCPN9a6BKbLsaz+NXBe5xZvi
SOQ+1Pbk7+K0v6v5XvsqFO1e6rGmjRLn6oXukj/qSkHLZlR1Hc9iQ9nJNF1vv7dS
oW6/rk6iJQKbDb2r3gtjuZF7oLXaEbEqVHHD5Py4gjXo5Y7q7G9dq9JXms98JdsT
uKh4EN5RauwpmZ+jaStH4N6y/TmS8K1PBzSnX8Bpt3SaiXkuRJ0/u8HTU4HL0jhQ
9EC9KUjWx2g8taUGMGYsVucnncpqESSYPuPz9ov4rZ7XAxnQx4BjwlutDs3Yc+zP
1bQ9WnUeyWCotCqOShLd42AcarosoqD+g7A+21TAljICxow1Tayd9XH6ykDUZTAI
KUZyQy/oFgEDttlhM4fwq/gXcqzvOJURJ4Ji8NYKWmef1wSAB4zJJeWidUhHT+ao
DSCYC+1gjZxexGafGEYBANhNfVF93t6Vl+8Y8sgm9Kl/hyzDhgjGVpuC1aj9y2F5
fPgL5Vc+EcV11v7ewljfKFN39f5lFXLgFLmISJkjvjrbhmHjYuugz+X1e+dBcdhL
kDiVkOEh5/4uzc5jhFszh2uVkAH8B6oSEOMd4nLXIEArR8UeJT8kXgCX4Wxh584j
AbYpSSvJwVup19xJ8bgdLBrtxF6gqatcZ3mZ0+px0qskp1S8VJHmA7aH738QTYMo
uRjlBysgVGkxAe8iYbya7jb9LJH6IC5ZfQhli78i14pGTGSg+aGkgUTaCg7ZdvnW
TSRgWa19pjOUu9jhjF+1a3TkUyI0E1ZrlfVGgxZjhNDKhND1Tm08ZEl4HPR7Hchm
Dy227JXTATqCiCV12+ewFw==
`pragma protect end_protected  
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
b/ueELBN+YX+MNOQ6myKEf5kxeMxQeHr+Qmvgf6+gICPq13TLszHio24d5xnkRJg
OX5zmbQ+RJ0StcPtfboma1/9uaKwJZy8w3AxoK4PohKipW56b/QoLD6F00w08sW5
2X3Am5NTBPG+G9TVbG39Wh0pMtllvcaUApw/o/vbINI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 95917     )
PEuD6MqPpfA5Sw36ZNxDpo3J7/fakVux5zbgsQk7YBYd63Xe3kl5cZFmK+7XUhCt
qcwo8X2PY45xdL5mLG2CvrPeQQCjmHcBnbTHCEIQABgCDhv4s6hl9+zPGEaf11Oq
lkHvjmvT/xknMD8mgW1Xig==
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
AkMsRfdPlQY8HVr+gxBxGZi3K8qw7MMkBxLztRUZgRmfYxNnGKPphwbr7Uj7Jd2l
ZX6J04gjpmXCM7aFlQDxLmeBh2HrSoZh+N3DwcOnkn8wqUyWCFJlV0oYCrvHILek
1VE0ls9jOChN7/n8MfLf3bsw0B0xhL2BmLPRZQL/0lE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 122795    )
HFagyMEE55OxVe2A8xeFDo5dv3rNRlJf0Ki/f1GsmS0cSDk39ChstnSHZwx9x1rE
TBwTbEyAGr/4uS0KRwxRvjFu+Ckj+rAaL8YXTjDy3xfmcyujgJ+8XnugfR3IMSc2
Cd76nIrAi0nLdOe2GKcBv9S0CBQAjEqeMHYZSTcxprEUhwuNi6NU9TGV8HLUOqiU
5uLdD7YsyA33J61W8I4s/yy9DuvgIzndMXwo6HyRHoFKd+4CllV5IhyXYA2GcXqp
ugv4t/JIMDSjbwK3+fzKj8HsJVa5oiVRCletoBSYrXlwxX5UswTgJVYUzJPDo3Jt
pNB2HVAZ+DpSlD+kLFR6THyF8VnK3UBoua/QHn93sTVBd0RmFhtK2YZ/0JPkTAxJ
Zcxdscs0CRxa3NQLQDPYzvf2w8+EjtjycSL1SsTSFxX2++SvsrfS8iEKZ/e/xfPJ
UL7xK4bI7ZtfyL4wg5ccDNo/behk47tsSasQ1ePGga/KajCUNdb0PVNGIuOcLTBT
tY7wvBnzcvBMGqKVmfTT2JvJ7s5ng02UU+sSZkHvpOnFmfx54ek1AgfWBIkWFZih
aCHbcZL74TY4/NoZo6mLSs6frMjYdXg+3D9FwLjRf+U7FAsQzksTHR0KpG6TvMho
E0VlVWrcFpFWgMx+jEGjoA31MLLZkSn2804j7REXproMk8yYjRMoE2jgtEkwOmxE
1YMSvWAnkcNHsVk+I5DVF8CcyKwyz5Z/EkNb9wUdwxAh+i32w/Py3K/lGOpMI7R8
g61/vGsaf+oVWxYLyH2zicexGtvruzgCwx59AjedzmScLCoP24F0TJkh2+xI15wB
RqT5qcjtL3zlyswX5qOmElBJA95IXR8DBmrTO1HzZnCjy6mhohNwxsVNk4fvAG52
QUeFeZRx31Zh0DYC9Yt9zSvbeoYzU18qWHvScfDg/js8qsDHWykvHgbE/bHUUd7c
Jzi+namFS4wAuzE4eMdBHVbD2NZ0irQY1nYDfIRl9pGffONAG4jVoNq9/WIp91Lr
ryb8dtb3uQ6vpuINvO4DRYqw05Nq9abJ2yITw6mZKi09zJvrvpm4JoMOx5wSuPqH
3cjK0LXZHrJUnJri8jn//AeiMgqu8N6cvsbycv6JT8FYwmB7MuG4OmiaBBZpJkap
czDaYA1hCUcB0lZEiIm66qtP31WIYOSpuarkZQcTxwyRTzjkXFTHJCW3vyfhJ2sP
1PD6xEyapJjZMrLwPam58Fp7sIB3J7giniKW08s56rEyacleJISTC0nBk7rxn8rZ
qPRwcSuiz01Su6YJY/Wfy8cXa32V+htc6xRUQujJuhiwnMYDGWWMTZZhsGfe92Zu
tHKyCEqgfzJms+3+EAqBHHJXcWIZPaS5EgFCJNgNFif6bjFj2nZLi42P5se5EpAt
cdE23UZLag6nRBcxmzCJRTAtHVy0qpTmCX+NSFL5FV/6mx8coo9Iy2W1JL0MU1P0
w0Na1CP43keg1lbIDZDwp5Z6lwK8vFkaSXNh8tbyJYma2yrX4aXOBsnKkNkX2fS5
Zrn4EEHQ1oyUCyR4863xGVCVfHB8LI5Ly/5bVP6oBJeNBP0EBMoyU/aLkc0iHz+P
nfoCuUk8OnpvVKPEInGf/m3baJ/ulzkbQ0V+gsZ5hvAy8rRYly1SMLYoyXWCsemd
9bP5kN5JH8tnU4I2Uw3CXtDRnJEcZD8AAmLaMdzotFTwz0i2okc+NygCgyMN60AA
X7FcTB9Hy80tEngmwZ0tdz5Sv1x2viI6QkxEGvDkb4aRYGYabtDTyGoAMz33TJwA
iqGqFO9sz788MAs+v8HIStUvuoHCMiYbsyTVgbnSHsToROcAT+IFDAg5VtSylNrD
13q9UN0afARWSfCWlIHFnW3KjvAuMTt6lNodKWwvOCZ/cWhSbZcjkIWlnhsAKqFK
3/6iPVmLFe8k1Hq9g+gXtvrl9emigW3Zng7lItijc7SzuaUyseR/7DP/JGRPGV9k
fFrG1rHQEN9nrmYQA1VUvnbPnb2fN57sWdfaEKqvSM/ZqcM4USttbYK/P/sZKUKN
x7FaYWVCdigoquqWa1H7ysmWURS7NL53o1MpF+qe/1REuE6aLpZKx/x7OJXH/uAm
Exb+zyxb7iUlg7JNOFnlgeLuymULCoOXAXT2ClNSiB+bycZH3js2sDL1irt2PT/G
sjNezFt7NbJJrlcxdEF6pFNR8rpN3DRm2aMOsL4sjncwrMdks6Sy9tY3CYp5a0Ca
vF2BqyfDO9xmiiV5L+DniNKhwbmvz3ujt6NmJZ2rcxroEM4c6DRV7qi43BIXLnvK
dvF9XgR1s4SIMK9DIOmoRDXH9tz2l7MCauE3XwLg9gYsZ+GLm9zbl0wNnlIl8cWw
2Gv/pNjbAO4sfacHkZ7LYXd/i+PUJTq8xaeN3/qHMNWUhPbUmelT/TwTr/bShefk
vmiWPV8tjVo5FQn2MKKe5sp359/0xfVJS9CuHEc83cHYVcv4/NNZ4erH5cIaR9Wv
bHL/BZknfj7gvzy/H95bpwX47kFEa9u8p4iD7k2krtaDNkNemnqpE7LMWs2KrJMK
oieJLNtAs+7e3vnEc9fbZQ1BupyPU2oOUc0k9/9ob1PrAdb60nnEcvdz0wHlYpiq
kddDAAxITfssBl/aAPm/TqmFFOKfClbIC+c54bp7kQwAkbtiDG1EaTSD9ydKmc18
svn4v+efI6e8Wt7QW3U1EG6qIIKMDha0hpop2GvijWF5Jk3o5gax1zBbhK8WVEAl
ElBzPjAdjzgcTLCEOmY2Ux1ngO7zYguMf0qc8z4+PX1zqKzX+9bwsHwqMiD5Pm2F
l5CcmMp4xskyB6ZnQT8RLhUSDeFhMA+AEBucItpuvxFDBOG22T8Q2ScI8kqEB/Iw
iU0aDt0ZLkqNSCu8GzZyexeGtHf8bTCfjqE1NzkaDqIO4SXGzsNCh6Qd4Pwevpm2
XfdZZ1f1EplV5ON9B3zrc84/pkhDmSMcz3FDSFB/iuo3WO+rTNA+amhnfk4STrA0
ppoJMq+dgpQ/4TteqcvHSTHQncVPJasv6lcBuhB/gw/tQs38t662+328KWkwc2ZM
f+Xm3Nxl7zAH8UDmq/2Gj/yEXsmkMsIh/tFGLia5qNYRDt662g8AskTbhSAFkg/e
COh+Ys5aVdkJQ3VNCrYm05+FZ1tyJ7eLQ7+7M0gZWwLGIVuXKolkoUFHHacw584y
sQTzU5V7OJw/b0t/3Y/S6w+PV/UmH0Xo1U4ryCPblJTPBAzrFOLfFMudRMwrSCnL
kITrg91Ujc5Qvu5EP4ogoaDWHOQtsppXdQWnP2uoNEkPSp3QGitR7UwNf8j32Sj3
QLFdMGAYJiGP61zwEyPG2yxCQwT+rO0MlL0AgVrABSHPan8KrB7NJmQpwBOhLFm4
RRp3M1Q5J1GEYLO4RXz0ilbVmQK4+xxJDHvAuXFfu670dPJCACu7+0YXZCqufnhk
k1NlJSpmYyB3NQhHwR/NIV83pbH4uG/gbX/P2INftU4rR29/BYHqisN3VisBDi/v
BqDlSGjXVgPcI7GdMIPyuzIkJDLKcPSOpd8jpF2LGusNarEFqP3vQr9ePCX2ILgh
Itb+bysuUFb5k9JBsBRSKAkITguKSvJT9ces63IGMIljjrGmD3iRC77krEeoukml
9oZyejKhAEtviRE19len7b4EI/sVDFQjdLTPhK9XXX4NkdEgBjakDhqGpzB7pZI1
dT2E6GupmhFIkl6Qqc90V6ZKOeUG7Z0CGsiAmt6z1kS27+un1vRYnvRyGNyyi9oM
Zi752Iljwwa/GN4ztSqGNd/PR3ylw11Yvyi+qWeaAJ6dkLiBp6bJ/QdIyecr+KhC
k5ind2gC3Y1PviDwt5tQvIGfmpX2Hd3klmCw026qySF6BT9sYlQO63ijQKSDowr3
k3CqUBkc9wCIaYTYUlkDs6MhwFYIXY7oS5xxfwAOu6ZVBF4rdkp3ectI3NZb8k3i
Ux8wdBcbFAKE+vtvOZUzsJRYxpw9FAmUPCyZ03yYgLr3c4gjXZaf6ioRphmFXI1D
N+6Rd9zy1im6N9hmIoqqVb0qxjzNurLjLdzupujGrYhJU0l0An7CWKvi5Zs6UGWy
MZz8flBwlp3hH9dVLbasPvn2XZXsaxy7tZswGNQTmXlzGC/l/0Jpc/FQg1HuPL5g
Z9OB1IaHu1qkz5J3GQsNIfpo846FxGYWUy+gPRCczAgwW6QpCtwKDsWZtqTVpdwL
EeG7eg8gUoE1Er8AMy45TY5Rk+JxlL2l3x9wahmWOcteHoz9AHfo6MhpdosLCdvy
uDF37uX6CRve2k6l0mA6YKtjPdig13EMeoqiUnFThFTdR50CWe/Vrb03FqsMPJvm
1+dUfwbjGztskTUJgV7mwYHon2G7wnufkXe9mvQghTVv0hYeY/EyJIdg0H+PT2bC
/FzyPPO18IcRWUx2aBQTextTSKL3wwnGVp1GAw9NOuMQ2UFBU05vcNpsmLuvvHTy
8L5ssDQcnYgN5LfbvtQ15tH8bywv2/+0Wqvy4kTElPFbKvO8k5lrEMHsXYaKvAur
gtZTwzWEkiTMN3DA30/k9j0ovcnv5KwElUjelCV9iZIzZam2tJXWoYD0JuvGanz8
AcOfJmLCIZq3VEuh0H8DV68RorkAviOoCCGdfnPYVY/udWj99zLDAWG8Dq0S9KGZ
Kq7fuqBz/H022rSy1J64nZOAPHdiOIoHie9iLaXY/ucETRQ4kADnVEcI5DuNkUJC
+qmKCGCR8hh8DmoR+J6PtKW/lomo4rO8MV5mxEEqDpz7hugl99vCkcHkPIxL4Coe
kLoDA9n7u6r2sco0cnTt+rIJ0x2bZezAt6tumH39qLSJ9b0BUACwI5iXu9/bQf6E
zJj3hIqWORTwj24rD1TLUCm/BKezHdadibD4SZx8Hld7W0NG68+ViANQ9uUilsRW
1QgoY8BF38SsZ5FA/U8PKYz9Y4R5RVtv0iFHTW8uqmqVQjlAvs9gMxicLNxPT5Ja
P7eG4YnRjhpiITEcPkr0AKdhrl+P1i+9wXyEBocjDxpQOSc9Yj4kC66YFA9GakA1
ByZwbYP1+6lcQrNAiCAzNoLVUjOykgcl+/ZOJFIh+q68rwt8kXgbH4eotxufC4GD
bkRfr4WHulrmx+464rXSHQklNLYUBlFzbiUTkDAaG/VduCtxZA/n3tbmxNT/SY48
h84lTXzXDporM2eQWs6se+5kGgo9rQuVmQgoP1VyIakkpmFxsc7/RUVwQ+F1IMHC
AENB8IZR9EqS/o27dHU25D0yhYSR8p7FjEwt+HMwsHPiWyF5k0r7KOE3gm8QGHsy
Gss9NPvyPlxZg2L2P8f1XxFCbP0cS3Bc1P8ZXeykeB5tAgKKdne7BPrPzGD73rmf
YL5ovK2v5JuoL/h4TqxvhjB88Zbfd31PCl2TL7M/r+PnfmJHbqN2HW6Ln5PtEUUl
SfHgbhEM8+ljP2a2l2h+CkUKtfzdkc9AVCU0kS+srpbyJ15/GRz7UTZWsgJe8dxC
y/PVB1Dloyxq2sgQoFdycflzMuDb3cFF4fAhOqmyiLx5prps3DuyZ1OQcsGtxSyW
xjV5WiMrwnVC2c4UQmTx8zljpoad71Dqr+mecdrXaHkyCcdPr22czt4sqU1yZ+Kv
x8V5ZBz+kgA73yyZLbG/YiypXnV7+RN9yk5wArQAdicEOFHPWN08aGiBY9KxrkIR
KnO26LWDUckmIP0fDj/nCl9ro5fYlpGw7SF9WJn36wZAHiDYSLyFkMSqQRnBU7by
6kW7ej4pbUScOWYIlx9mcPYC4qdTuwuCJZ7aQ22aUJh/4kMuGHDT9kHzvf6RoNwu
YC6GAg0yTFzhRmN3ImwC4vDOlpL9KwTXOuzJmDmqzwYA0p/TYZk8YBlkRlgpHky6
AVRoV1TyXfYQWy5en1lFoHWo71va5AtcnSmWH+1XE9ADvBjhUhw9cwNgEZKEHOPu
RP4q1jkI06+gntOhXO7s/5TBcBFbkwGZnVdtWiJ+xUStfXq18xCgyZq1e2oE3rR0
PGv+3EVeNXIB40dO9yoKf1ssKgb1b+9aFuCYsL6ZBNMo25oIEeXhgcB7OgPeWT3T
EL6z1DUmsS6/RLWKDnLxIESQUeh0tueOLusxWjxIpKJq7xeL4go9Du+66HS/kQrP
7G1TZHdmnMTXOjepUt/beS+Ctb+rn9PbAAAZ/QCC6i10d/bDA1DIV1dl1FYq4FrF
oGVxufYmjdDDyNZynFAl1FRMUIYuf7j5AxomMpalmGxhamxCUQEjdjm3i1awI8mw
E+ZotpEGDS86bXzhUFmPsYvouKY7XoxKhbXoD39haMqgl9/Unua2AM3saKjsaMTG
jwDPoOed1toeYF0l1N7yrqhjTGz6pb0mTwz/Wocv/bWm7h9i1cjIZ74ixCpg6ufC
aQGkGB+isicxway+LOqgwlvDRFGNAJa95Q0wyDovCRfWu5tTRBKuaAANGcsKS6Xe
4XVam1zFHCUlYbgfCBaY0hNyQF9uieHJqq83ooqwZvVQuLXUR9TsESTOUA7mgFqq
199gJ93vfzyLaSBywrrVbw9ru21GJNNfACyOfi0XM/8hix+Psj6sH+0loBKrOBet
iQLT1kXf1A3ENGTZ7EJNkdH3nhyKU2vualqwxdfQUuj+Wu4DTWGcHrZi9ls8Jf+b
ufN4Qy68ZdA1lrUvwlVHaRfsQqJxzXuTXRwLZ5miagUffdOBPgoKxXyfT3uEYsBj
sHWmBd1xAy/HA+tHI98y7BtC7gtyEk9I2aEycwYNuTpB0/OPfQEXjhC6uXPO3pL1
jB4fNWCuBXaneO5Ypgpq9KOejl+208GqgQKtFapL4OdMlkJnv+KcaqQ5cBOzcSyH
qVHqfn63du+0wkz5TKCGovWgYzvSSKGAqxfsKZf+qsvF+fIv+x0tloG5/6BdGHD7
91AXGd/dWAoZp4FdOEq7Y59z89A/q6JAeyFIWsAvgQ5dK+e7jRczPqobC9OfnzIB
W8Wv3rGC60C2oKAFre4IvyHeXjeVZ0FJPMJ7YQ/zwu7kESPbCsK7PriVV4/Z16Mj
ZGFfh8ty+ZXTy1A1gbIqDAl0ZxwEaRniqKStM6/Z/x75isYCJ5qDu9MTplyaLEKa
JZwPkrqqyrVfMaUGZ8vjNSFgCGMAWfwYYMNHUc98WiaqZMW4FJPzn8+xUWMxdRke
t9k68JfP9DXn3Y90t6FHgW0k8flbj1wFa0+cgLuAErMF3rwhQwqDUD2HoSp5qZCo
vMsLiqiLurnrEnukg/grwPjO7kUuC4kd9tipfJ+twal1Z3A9a3RK8U7Neg5nSdKV
VOCw58RNbSwB1vdChF/EOM/FAdUrzgq1gkp8mv/GZFugjsuVAO5x1khu6CQV8qPX
IIj7S7yW9liVLBJVo7sPPUsLbN6oYRBI1s/fmudhPBZCvFmhTQRvUFKwlt60jR4J
LrrhSfj8Jxm+R02tTVsM9vG7ZzrwU8mLa/19ECRpP+jldp/gZ8oplv6IixhcHbTN
lqnUAFwNHyP1wB0rC28aka9PvPpNkunQ+iXgvovGpTvtQD6KR+0jTIqppSzmyLdG
IlvI9YMUBmQT0dC4kcKjTOHxmFBoOjLDAakdcUr985Cd5WX1tx+dNXyRiOwYxFSY
lQIfuhJXDEfqvZEBsWISfTLPJdCj8TPabgD/zFKomnQgmpoznaQiDmhVpvLQwBDN
dq65r+YuV+sovDyesobWQfxC4SeIRwbFwglbY7Uq24MG7IrkUrnRmmbW9PofhCuI
f/4vH9vHYqdx+NqQHeXGqq/b49jBuxT7mBSs9RTuM0uvj7XaOOcQYaip9V3VrWYC
JyJBgUdIstnjtTbPfsxjdjnNfHixEfR45aulYD4ju/2WQsy6g/xyc3GM18MqYNK+
fCGdxzLT4KKYUKJlsps0PtICfGUc2oGAFJa3xSND8oI6lILX+LVmcmiIB6MXJ5q0
I7bsPgNN6+AtF3ItBRnoyN8ZHhRxhqnpWYBpNQ0kjhEUCimQHXbXlDBeW+NMfFNU
/Mt2nKgehA4tr6NeIPA5cppSaof8LiQUqCJg5B4D4wbeUWdtAg0njhCiqdfrDNVd
MxZZfGYVNZe3wiZHtO5+4c+SyWu7heR0VwArNNpzKGA0mHe2JEgsAVNSyeJ/vAFG
8QX9h7p1CzvUapXi7myOJJjWlgZjuodJUi3HIsGvD9d+us838mmtvn0hfqvqKZZR
LkJfP0NRlDgGubzcHoULViFVhuY1tEhlBXDRc31FjlEJkjSJJHvuhsv6M7dwEsws
yx976SFgzAcRmcf+XZBwQpP/ycfeGeHJPBGdM/7x6BDrzBZ7eQUPtEa42iVOs3L2
6GVIboL5ze8qLYVnw6iRAzcuRdpPp0/t/5OCZmkZYBje+EYsMjyznpQRcjjBhk7S
quaUoO4sZbtFxeqGAwoHfHNS7PTbCIOe85P+hRKczkAFRQ/TXZGXMHgFVo8nA1Wg
xUz1u9Rf9+/6n4nZS8ED2cVxpQGKVx1YdpomenMDekSXG+fSOFFGdMDfZKrkA7GD
bqewSDhVkfdzKHJK6ix+J1WvBypvApXxLAdZ9ac2Wuw8RkVVMMk/xNAiHy/bxoo6
Avv3WwzhfDXdZC+fB5yshXzI8+pXtBMk+I32NLs451HMnUO2c8mZ77jFuyblUjcd
XzDfVHBqC+9QD7bEcB2tyOpBzQ6+zbF7Y7NQ1AmLRnIf8NHRz7MSiFyaNBALp8dR
oB5wJc0S1JC3lLGD8fJ4CbGVbdPE9pXAJf1jKCdBqpjiabpfeyWueh/e7W+GeweV
QbpKM0iibq/+XAgnOv5dkuXWeqi0O/0ILXdtSsPGHJ0kwG3D+U2dQQsHpmbaoENl
R5dDsr5uPLs7HHSb+kkcPBd7XjYO+zWW7jrMXESwJEjtew1Sfz8uWST/luqAZLnu
0K3sORW40Vq/6IE47/oDzCrJdd/4KUmTYoU4akzJEABs3zL4WMfm0uMkm7xESE8/
py0liETbiLsNIqKntqtDu0AmndTK3GgRhO8hZl7We7kWM1Hx0JxE2bMVRYQ4G48W
FkiRvBetiTAfMTAlmglYrfk19o+GNp9xNuCPLX90woR4vZfE0U8jPH/mDmbrpJSN
NkjqFBTm2HL1HdYOjhuMSApZBvygO+tOf8Ng5AtD3W5UU0VHofl/1pZFhSIrVYQm
8vQXG31LuOvWzuGf1IGJr8ZSgr30oMStTiWK0zw6B26uNKr2NG5oDAwlYYPQU4JP
lsXuG2p3R1+ETpmzHBw1Ob+WUmkyOXKhCCgViWZnMIFn7ZL14mcvOLCDD9yTuwJi
Bp2d9Eh4RQlGmApbLN4/kwKTnqsE/K5J7/dJTzDtY0S5iyJT0A/F2cZSsec7fI3b
ZkNHwjgC8rN1gEQDdMO+y0wAQYkAj6e4eZWtYLx4gHcycyYshkSj/gT9tv/zhYbH
hH2nErx9PxXmSI1xjrXXlrT/uxbBLm4jU3xM5uc2AYifCRicA8Q8S5TprQPLvbCT
S+p9LphuLNDAoD5k+vY1vpEOIwg0J7M6WUoD+GBR+ozttFHj5ij3DbccZTF5dC5T
xZ2K06Vgqfy2P35vfnO7/dsLBA/ni+ygqM4xT5GodqrPBUospWKlrL7YPav4GdTh
XKpDFocLV0tz7awgvoAnJfR7PPjMJ786gfZAV0lhFUk0Tadr/NFJM7TdJqR9A93K
OYInNYq295TpgPESj6Yfmfus5Jf56k5Bq3sB7D5ObkY4KwGkgTEseUBRTTcHlEbs
5XTmgaQOUaLwZHhzjGQbo6Tl0kWbJCawlcAqmPN2jPNpLVC0ELVN8C43PtEOop/Y
1bGIvx/gbh+nsY2kvINo1e3hwLC3/dmw0eqHFupjyiifOKkLyDrkDJUD1/JF8sCu
xfH3Zu9AsCqTYQ6TjLYJCjeRRrAUn/dgOhOrA1MtQzU6NqL5yA7nfcRGn6/NDWbM
Chc1QPLcTu1VzENPY9ct4X5E5vGAWpmbegIasDnxeFYv2AUztvUU7DeYw7maM1fd
DsGc99uXbIzCZ0CvL6d3OdZiie7DVAmdHhfNYn3AM7EQTdr2QLhULLmXIHMtEfDa
f4vffaIcreXGUH9psPgqFJ9CzPS5GfURftH2AOx9SppE5bUxhxw7cyw/QIDq1/71
/wrynfkCs0cD11WrAHikltrSOLo2tuxz7vu8jHyBn1Gg0PRcvrpYZALkaPSQsPG0
+Fv2pPl1uobjWKkLK86BAmYB3EEfuhpuNr/4vSxC9WUxn7XceyuJKSyIVkxM9An3
Pc9Eeu6GjfjqA5IyFIAtAK4QT5kM80YedVzD/ij1bc21qd3d3O7VT/8Cmve8rUrg
g/13+UZd6Oy0QmPNRGxaeW0/z0myLgWQV2/SKVP9Q/BlLiLcSgQFmCpEqGayTUvl
8FaXvAc1TNgpGd4eq1hJwJ4o9LobgZFa1xlbmTE6P/0NZ3HzIeROLogcxekWbsyb
OZ4UUx9UDrijiMumtNidqHAAHjFW60niBcGAKTYMDyM3TQMZPilMXPkGgyGpGMRH
RcrByVHp8h7xpO6qYOdh/yMLKTUsRu8oGbKm8XcC4QlkDjcu+kd+sTIvw60PnlHB
Dneoa+Ap1TMU5ejfABcy7zDyjwNTRWQWpULL2PQhT/Iwk5aLkK+x7/qx0G/OUKKe
s7PMViVqc+E44vQSzqG3NZT0lNWZenhciPYzwwq1ViZkUqkwLSKfFNggu2HDB96o
4CWej7fqUYgAWFaXHLMPhU8j7uYgYrRvSQ32oUa5QCLlqHaizLsxfIHAIYmfYwbu
aPl0uzSz66kBWhtdXFzQ+ojMo6ZW5+P+NZQst2eHLCYSX+03jXooCf3tPJdjSvAd
LaKQOdP/Vja7/IqI2WsGRppbPAw9lEv8OpRjbMgh2RH2ZWWcDYDrdhefgjHtL38d
1Mngkarq8BlwKEQDXYjUGUk7cgx3BGIYYGxZmF1iyCE4n5r0s9IGcy0www9sQOyT
FP++quXAAKwWZhjlcbFxEVLrrr3MZRu+z21C75ay8g/7KNS2rdFneXvIvvDoRR1K
yUZI7p8IZNoj/UevFsyyIfKbOf7NKx9OgHz8SssTVQaOPnPfO94E9LEWc/dOPoad
2iAhL7YeXMmVkJ8nzb7FZ82T+m+QHn1dEUlj25RuyU+NS0F/2oLYmL+VF1OLJw6j
rtHBsiwEL8aVRx75GuCtxkpt0fPYs28dQAzul2HuFR7YN7IJI2UsJ/w7TOT9hu6P
/9JPHZJsxlc5+XOmfxIj9L6+QSLPkPXyUwTm+seLBoDgz+5CxFPqpUz42Ok68j0W
MSuTHssCYyQ+lZ2EGBIijQBrRZt03wEUMHqp75MQ0HtHF7MYyuELo832jCGzAiDb
mMTtp6GzvicVXGWe4zTCxe3591Cx8ZE/mW/S0D/o42dgKwpbNpoqJBo7DQE5aL48
9uskz5WOa0YJaBH8A/w2H/YvbIbI4j72F6SB2Yu7lDDDSM2PsRNcP5S4kbHAvhd8
vqJvw0nYxPTRqMxE8VgzFkN2sv8k/zeRrWzzk5dZ1WrQLxSHvTE4sAzqHl+9+as6
GZYYgNcdJyiWWx+eaFco8ILlDj/C8ljTkgeAE0H9zvmrG9zHLuvpNb7MscSGibyl
mOWveun8BsdGEUXepmkcBQQS8momLTRWrrkj1PvUEwGmPoZGdWTFmS0Q69os86uY
hn1swYnCOo7QqMT1afL0B0Og8Clahhcd8b3s0g3ZhUjwgEnHX4ID6BqJ6W8D1wbs
gzdgw+RMOqKog6RxJ4G6MML2rSM0uytLQsCWA5aMboOgm17xzpDMQkHXm4LrCANw
DFLzm5C10HYOLHa+8OmP+pLetKTWuxa+0QYDej93qWqtlolMDX/Xcnb/mjDdpXVe
PYXk+/r49JhQ276OMMqTUnfa74LGr/TtDtDItIS+6xf7zmEtYTHv+IBNg1QZQbOB
RnoxeIPL2N8l54BwMVzSKYuWzgkOjTzI4m4Zjih47m7JUcYugyBRO8tJO9XbJyfU
2brxySc84w6l4Wjni12A7kVfziMgcIucSrM4FAtudrDwPY57SvYrX/hC2vSVabK3
FSagQzCMW4T1g9yhv+5M6JBmaNb825Aodgi7RO5lG4U701GP3fsy3YXeJq3uBIZQ
KcvsYiq9XFnskwtfk1cMMkk0KKcZakCyLXuiXUx8YozaFLA01rahbF369+PCg7cw
vIdKsWjkp7kkSdRXa6K9tsdXMxJxP4+H2w2axpZeSAJzqTKKZGmCIrk3fyplmeKk
BtfEWFxKo9yvjncfyxcTXOfEHKRY3lrSoyqrJdT8iDNqMFCs0G2e/vWD3L9OwIyq
XAQTYYZ2CganjQNqUMfNDm7b+VfI+H/30Yslics0vHV7+Vbn23+U7FZVSO2SQqgB
0R50lArW6v37v1FD16LXRFzb5EBijFN/BLfcgzJnDQhKbqBGHzvRw5EKaOvU3cFj
9L5cFqZ3JY/LgowocwgzSGm0jhDKJTE8gtPEs4w/Xk+n3djHAEUj4Kxp7t+kLRta
knGi8bMOjn6I5kcpnKRsKAzJxIZfLx2cwFTcrq/F+ASZ9xlaHZF0+LorQBmOmhmL
/t6keaRBPdWviY/A0OnKwNfPsRQqlSJL7EV0uRvKM/8V2e0gOwj59JeToSTX9ysX
okCosBXSYqRFzaeearCugInyu90B+Ynarqd1qqpgKK2DDjI7xw6UwpTo0rc6ufbc
lceIPsE3DMn1BrtPgpSi/rMRXJpMB8lNaCSIXKDowZ0wYQ4IPyO9sQN9ULEBY1w0
asfLtJujc7BsOvBM1NY1L3U1IITxv9ZaB5bl8aPF5WbScvD33TTX2VlAyhxaZR6E
PW5HGxRirc1jP/Kr6YiBYPt5LUvrpftmqyQwHBfMSNP6whDV5EBUwbNl/RHTijZy
yEbLW6FprhLZxJSCuToaIkA/sUjW62gxD4w7noOvMo1ioMrtZBh52+93iF92j7PQ
T1WQijZ7S565BD80BO9q1tbldLPrKXVmDeMBLCgR/8LtovNxHyMnLiYxtEiRLYsS
q0xTEcSNy9XUChgFU9yqQXSf3MNDQ4qmwSggljUQXu6j+cZzWWMA6LPBnC85ITnC
txyoewlf3BgEXVjVKu3dErD3gZIPh0wSsrHQaL0DWa8gqku/ExHRa57FWdJGwG3x
+sItxuhu3GL25iuKvBnBaEsFLYflGju3/bX81LjlVlcrskzJ74bQ1DF7rRVU5GLi
bczi6opPqliZSnrt12BCroqNILZVC/JU58/fQEa1aG/LdX+8wOcOj1T9G6YJEDQy
NQp8u30zvhFM8WZI3Qz+jr7P+T/ptz/qhEIe67TcQ68PsLYsueik8Q4YgGY0uN1R
HVTWzzGZa5/CWLVWAeirjBSOP6SckCCX0xyEkleG3wLJWvEE94tpKYWGI08sqJ7y
OPU7cPUzgQEWAR8KruXjXIhaehdQnwFqI5R7daFExohnGJMl6K5ZvsRAuRj9JYvW
SVkc5gZ3PhnhobgGWaIHfWWif3deNeIZCpnHbftN4qKycDOpIuGVxT2yVAFzE7gw
r/dqJrXSev6lDd09Om9gI4M5q5vAX0GhvTmJTKfI2R71AkRJv5Ba/OWJUJvj1HGT
tZvu9EeKGrc6rNUyQKlDvk4XX9eg1+xipN4vtXSs2TywSI0sGtOTBJKDOtt5D7yR
/qxeYQFydp+C2QdhYoyB2/kosxYMgqj3ByzqZOqBw0yAltKHGiNHQxropCjvbczk
8+9KvfhmLb2aWsd/9OvDsn+jFVDdVXFo/oMxMm/6pSpMbaTC+NH1mBgd9ze9zrak
DkJdNRl2uMG/sohneoTbljzLCuIqyd6eviKHqtv3VqTEYrIGffBY74zFy6/A/1KY
9L4v+J/ROWg4ZTVvPXFx2mAvtAN3f0lZI97D+hT+HWalHQPn7hFIzCHWhBV63nI2
B/vfhwSuU+sX3UqZaGgg1cHYMHwL8HFtjuNUA0MKgf18ieffM3FubEMS7bj1zMjI
2i/jn77wy2dgGxQkRS4767kJZnAa0DYg+ljtn7dmVTa2y8AAPgPPR6hF/y24lf/c
lLUd/W0K3YRuRoYRnWfiM5iosLyoHK7SL7w7WUDE7rt03d+X1zcnkIfTXum3a5lD
baYHYI3P3IoDcUlZAKzJLWBNBRNQiKZfUm915sr5/tu1srRTKZrUH6NH2nlEztc3
OTOMgwI23K5+ZFQ1ATEZ5uESTwVrDZaEn8ZD8rqzQHQcCeypcTdzpSI8GTqJj2d9
E3lasQwIt/Tg5emsha9oQEO/EMANvKtsSvwsQkayCe92ZtXhplhS1PRyJhckfp86
8e3UlkKhrvpBZADWfYYKtZkWcIjeDPz68kSUKLqVoBeFkgKN1rrQ9jHtFwk9t/ii
5aGLCh5Vi6spM3KuCG6Uabhs260/KHxh8PK7qlbo60N9NhSUQ5Nc3UfQOznX9YsH
qaGg7PT+MoJvWxAjz0KZbuwxCuSsbJiPuIkTp4D8Hjqb6RsVuOiOm3zZIMZ9/qqQ
5zNfa/46YUaXB7JFaqfrEbhwJOkXiBhuYuNjEVuLXEcdfoPcz2zHoPrwGt5WMSF4
yub4a4dTH/691kq63ZhYMEPs9Kexq+eOG7kYif+ADL0J6MhLTCvAd+vmk9WnfosG
s3PrEaavwKr5Yg9prJ2H/pKkU/oSPeCS626Fwu58J6kLz9/I/aaH6s3PbQN47Mh4
Ujx6Lhsufv0sdceTlRGY+XPa3k+S5VnJUrOzt6QyS/kLZzz+/57Fxosp4nAlOPoG
lawO86eqd5Tx00oCjwCk23uoKoik/SFhCo2X9q0+LRTaFZvsaPw9KH6NjL8WKRAH
zJW1+yVkmQZYqk07BzHxGFIkOI99ju28gkNGkc0cFctS/lCZQadS5uOOrrLUWSfU
9aKp8/rD56s+NsftXp57qpRp6MWMzo4zM6Ee9tVYYmbhZ2mBUbr4DExZBq+rurSM
bd+pXTayrDX+SKv4KfUtiGv0AQPOs+Ro0+1MEYdPc1H06W6dqYcbd3fWH37ZOZrZ
/xSi1ShxvQ293dAhXlJ+b28O1dLqr9p2LLOzswdVMwTn3NtNI8W23QDD0x9gkWmU
XgUN2T/HrJSSR5qycHLX+JQbnHbe2/1sZV8R/mmtHNJ/tLf7TSRHHXdFBAvuckei
Gehh7AGA2xujI8rdshek3ux6+Dpa1FYOvghn6wMkxwwGTpzl4zZzggr9iFaUbc9v
kKoFxyHzzjVaOILuSP/nI3WlxW7mtOheHrZkZhBdG+g1wjmLYQz+8CJ+Y4zDeSbU
5bXcG+4eSn3WrsPEo7ffJcBPC4aVnJoEYYOGbShFEKaf+VSvHX89faovMngV+6ph
FZbjq8aPPv8bF1oiqPBIM07iIcSqMSO4Rmw5/lN1Wt6YgN2YLB27ArsUkG1rQU80
FICQYeTEOhuEngbkLYUGGkGu+j2PhdmsGV/NItmLQqOCdm3oYgQm6NkdWnf7YIG9
VxK3cFSllbg+Hh6SBoWg/1lBxDhLhW9NYNhU+Hq+jOmsgZGAVZiCMxW2WeRxSJCV
vgg2+ICTaIR8I37bLIw1f6kz22R8JnwxiEdgbxJ1ycgIaxJfHarDC8Vsz1hzBLfs
kATgzjQVgChcDZG4ry4UloJD9ps8Uke2y+81mm2PWef7j6ckJ9obxwT8uuUcaX92
FvsdhNr3Hs/FqhaDuRxtcrs8QDcKHq7MsNAXXm1teHIB33h2n8aK0T+xHtTHyoO+
f7gekCmzFDSMqh5MSoyoYkif6V9zoif0s5zNgVTHmy5rU2Tsc2cxOMA4Rn+WqntU
snuCy0fhGXHTeHOJrhY1QmOpnUsTP50TcIaY3CuUHSVtID0cUavIlACdZMrRU1Ve
JEXb4RKEGmMSjY1aevA2ea3Im/GY/FHUfd23zJOZ3PfQ1nflUuqsswe5dVROAutR
D4Iuz28TeeFYoJk8VhvS1uo+EIlsi0rlG/XgwhHjcs1hb/hwS1SOMCOeIlhwK6CR
NedAgllBFXU6p2uwS3N7F/aWZ363gGliuG5doHfXAMvVk4HmC6IHxVolwTFcFlkm
3EMObk/34zHeAmYjoeEKzwZnn6sU9N5nxx1WoJbwgpLqW/cNGBzSq0W5tOJuJxO7
z9dN/n8HzZkNfwzVOBqoJuoCLT4WSfRM2z5kNMNDBNPHKKupWB6g4N6c2EVCQ3/b
d87JKq9vb9QU/drN69UROCrOCJ+Efq3HNMSFICYVLDiCZD6HUnNJIctLAcee215M
zSVd7Y7d+d8t+WGdtlfDlSNcWukjJCnyeT4oGbtLijKYM7hdhh5vnFz4BCdfKhmc
0DeHuzxnvdBxJzbIlVwiYUVNTF4wFoF9gGT4VHslF8mB/BtELzhcv4biREYMBoK5
wyrt1budds+83PJ96xFEhr6Vno/d9mW81F3ehxLFBrcNXwqmtoJ4to7wkKi5BH3Y
wZ+LiKXkyeNmg/ARWKhnz+I/610UW519Jtm0mUKY2hDoUxCIlW5/HOo06Gaw6/46
L4RV5n8CHBKUGbH4ODr8f1/DYZ4M8neV60/yafPS/G2prG3AEWM0F4NDXxsKpNEp
wr+/2+VT5soWh0yUJi+DHTtZANOR3ywlbcBsuJRf+7NSTuZhTJcWN2Bg2M0HI86k
HAoC21zHIQ2e1OmrXYhkgr5BctlF8QxuEthiKSo3aY66kxa9WkRq4bzhufERk9UT
e5m71ccPStQ8eevJrkiYUoWARC/Ak8Ggol9cUkJqog06ch73IF4d720cnAZbh8Qo
IoIuQODxENhzTR/PzsSjnb3uAs9j7kgRp4uGFb+FvgOMhSxcJDh6RPA0frNgX+iX
nTWy5HY1S4n29XFt69YB2ABRaqoPiji54jM1cWSBMpKAR4ERHlxhDbnu7W8tO8Ag
ectb2F+eSJ2+11zRaUVSt7zaYYpU35DlqdZpAdvZsLw26cRoY7/SCfLSKrw35tl5
ZOFeoy6HAOPOT8D7ZSlPbXi+8R/KTri3wMc911Pev9IqXlQ3T7JJgx1jUZRemT3V
E43l7qSAuzk/5GVGgdI1RnSp0wdE1HjFA6JiVYzbTCfLrTVZ3U5OC6FPdav/aDAm
+GIlyD33OHB/3MSFFOJhSWqUMQGg/NSCdP+9H7s7gBX+r7ZzmAn7fAvrW56OpqKu
MyafCSjdQ03Epi0pQvIF762rFTFRcFO0VHKCs/BN1b9EdlL8gfxG1mCmOl4wUNdD
uU7aKAd9Uj8d/YABsHmU1Z3nKvAtIzwG6gm8XiW/r/WqfBqxMH2w0/np11hWPs5k
M7hwxSiWU6ain9Iw45cSsTivdCuYsPlaOB847eoen2sEsNZLeumFzNCjpUb1kH9h
EAJfPylzvDzaFgi4mCNqJo0M+oYpJCLXP7pR7YpQL/NqgfbaBnxDGlS8QaIkPJib
hB9p2mp8SRbdchhgGJHa4WhPcLh01bFl323DznKW6TsCtQP4xJLIfbMtnF2JkR4m
wrn2wEzvF0yEmEesXD8X/2VVpuX67vAyCbDnnOxC4uSy4p4hQGE5okzg6IDgiTEB
mVLTOMyKjUhzgw4IPIxmOONsjNsspDoJXxSLj6TKdIlRAttE2zke8ZxZTTdGX+LQ
4osvqYALlYMZaC5w5TBL0g0Diyj7/U7WS6XwJnW+40A+exBe8GuCeCLAyUnIgwYL
GVOEQGP85tCzy8C7EzJMD3xo1Zox5g+AQKNJhWG9p3d5gIx6b0ly8S3m4NWimmod
OTFQ4NC7nVbSdLQAuRYjgsROTmKKeleqyqrdA4S/Yne3ygoX6GyvExrZwCEETxCq
8YOkhr+NcZXL2/YkoyTtzNrepl5+/xeDsF7NeXMJdimyG6QV8jmN7HYxD8hqODsW
GeT5Alk2JFkyV7ONGURqpUEhUHULIdYlAIjT/Gh0TeGqQBrhMOLxzsET/OD4L9zk
y9j5tI01uUeYbZy3gB2O+jEnIx/YmudtEOS3Nv9ckuPLTGNph+dbjyerYHxRa0gc
gvGqtvpJWhk1+cLrub3BQQZBKuZ1t3tVtxVsajlkaVL+dysEkbjti1iItbg1GoU6
RhPx0O6GjSPBKwmzzyr4EG6mTD2ntYhqF66BBduB6af6jXUuxjRd8pTSks3mgB47
3oaYPTqH+WYHRnW2rT0EDQmFYfMs7JWIgnVRzcnv9nEV5tfgqiywR0Hcv9bWpBu/
CapeWjBJwBPAB6la7sU3U3/ivbGeLBlwDxSdTJOT5K0dCqYCjGOtu5Bfcicrb4/T
sFSZEZPSpHQ/25ieZ1nPf2UhGwsL1usUCeb/Jo48jvfSCsTCKIee4BiH+2AcOT3b
fL+7wc+Fyk4O+aaADNuUaOAqNW0wWTzGEHehxrDkFRQeIKIpaOIqtBgGrX2kx+fQ
j5+iC9/bhqo5JY306ow3l53wIgHxLdBasgeh1BGzOe+Bw8zYP7tUfJ7PaMGIDk4F
GVKJTZgWo71AQCHqVHcqynRSMFvlebhrHIcIU/IH0jr9nbNDgOd2/52yf5Pvek2u
SQVYE29fjqmqjGxVDM6gswaDKyWbSD7zqTYnsULvegR2roZfw5bsLlFyVBMjjQIV
Q2MH3TF0roWHDh4rrG3xLOyRzJCycoTi62F+A2HOop/HPNcNTMsoYEQPCxuoEPGC
UAqkDc/rtaiRqbPwh+t6h0the4mmoquIw9N8qP/K8NDPy4udd7VLViXOl8fPQqRh
BIt4PUK5QMtuPRcuwKMJ8XP/qCC+otbgKIf+SxUxHw5PjXikJtObAndICYFtD1cz
L5tpQjHeIlktD2zR2gYtMdgtL/Dsd07w5LbG0784br6Hp+6rr4ahQLyRpKcsMz4X
xs6oWLKoOWytZTvMmpaSJEG+Kgz8pZsynPX/8sxQwDtRQ2Tovj+IlGNssE1GIsje
QDSik5jb5/knLRSdt7q/mdCqK+PDvosgFc9PHHyFKOLidQ9stSXV2NlX05E3Xsx7
W/j62OAYIvofC4YGVQ6yWlCZsWjBXkzhR0+vrYuBhbcpsVXQ5FYoaDVmj8P7+ZCj
cqoTyS0thsD4MYZQTL8q8bw4Uni1QPsrhxKep5WpUjJDRJZOL7di1UIxRPZM//SP
vGAyLnyoDoCLXLBZacdzDsRqY3hHp4KP3uBPdHm3lNFjz7r9go52UvT/9e8tI/qU
+zqL+zMreNoATARtuFGRlD/QxIsjjNGgDKV2ff3SIOc0C8Td+I91t20jr/1GYfhQ
+HlvHFfthBF1kOnoNrzZSda6C46Y8oc+mCe7i5aIL6wr3gNoxdpFK6slLJbvljYs
MKtup3ceqmzAE0lpKCMIkA/WLbUAtPvU5T4m3IjYV1FZIPnHoRAomCxaIZmj0aed
GhuqBJPu/yevm3IFGwGvyGu67CHyTJJ96EINRsjo9Up62OF28J9o3ABcjsxSAPs9
1LMmZK/lHbNeHhYQ64ntBqiuHw+5Owcfwzn0ojHJPd7p0C7aDpijaiSZvV9p3yI9
ZJtwWpuDCg4sSWGDnqJWVbZ43M6jGFH0P7IUF1T575XRRj7ac2iQ+B+IOpJoyTPp
lJFuoRD5HcGr77ok50DrkI+T0uB+Nj/eXD5K31dwKSYqMuzAOXcGMlzm6X0rUh0j
TYPYTBZ6CnikWHadq710AfbcSJ/IJy5VAg7MDA3IwafOSqB3f+Fcg8v3y9dMqrAA
QixnaB9oDIBAVkLVOFPQ7TNodWs5J1D01bP1zRUn+2s3G1p8RluYVA5v+zZXEuOC
5pBu5smzWnliqWgNgOL7gbxAqnIQthF3FpQRYKiTxBtW5tllvKILbcgKgQVuKPU9
xxPt+VNuhQeCPpHrDjiBchphjVcaTumldozRdvjwX5TiTqqxVhy4p51Njco9vVtO
Z0/pCRz4RHVtQPA0dlb2mLJ4hkxsO7D+otrAzuVC09UOFOcyHfPmO3t5TFe/aMuP
4ES0XuQWTl9aDWG1bRt+NZVtsBjSbcu8iyBAY48f274/W/wHqLZeIzZfhsMDhJCL
pWe9UfArU1+BiFyHoYsJ3l+J6VwT3HGAIYxq4GaHikMWIw86PKNh42ZTnvL+/gs/
VzaioMjTuQdp7+aDpwEzUzNdhOABMT/GwfkFIClerQ1JGBq6vkTjHPMf40M9D7My
Aq39B7t2CGY2QOlafDEc2N8sTx+b13g71pDeprzYOQVolebEB1ALCbEa6uumKGDp
wHG9QQvqU2xG7QOBKix0MszL7FLHGWfvkxjGe7qoHf/+7/EuMwDVSJLC0YwofQUm
Cr7ZWu3qIlm3srXblEk2ShPLilY8CcRKT0CrtbXRWPbf3usgPCP+K/FX5MulkQ1F
cFuXX2ASKOubk1x0gjG9zT6NJKEAjzDPMkATYVokrljhvsTkc7ICMwb1JsIpjaEy
132PWjU+Y//ENpmeiAStdGretHitJrbvD6wrTJeVCiUZrioaKtIIBLr2na7RlinC
9in7JuLaKSY/vhf086fDEenIywH/+Bk5kmuoCr7AuV9geRQZJbt30wnovztKkbgZ
uDsiiPKMmfPYSN/lGR/eq/tCAJVlhXih3MxrWJD0PHKHGqpNn0ob9wfC7LGH5pnp
85bXvDWTetSjtXdI82rLz2uKqZJHCTAb7j3YpHFVuK84PLQDdUD8UAL2kVfL4a9L
vvGAPiMJ85jv+zzqQHoTBI0ouibRLCONusOznyShBo7xV0czrVJHLCCZYuBx8pXm
bqrdQ4SSa5jgwAyE1+9sT1uIKVE64s/EWZtPHBuHNKu+josOuQi8hxoYwwZDcAXC
h4IMhTUAtok1oCHdX9JI87ZYzzNVOwsIUGYDhRQNbg1gXg/X1skpzZvKf1HdfN7/
u0B8DiSGR4f9BowSOsK7GQizou15tw/oqvbKcNd0v2JO8VAMMg3pdlWnRQ8aa/Eq
H9qGVrr6XPoJSZBm2JeJk7UJiFrf7IlZqPvXGRz5f+4bECGkw+RWU5uNIW+NMn6z
reNj/7K+lziCNJigllMcNfRJrppHI2mofZcVlnop1V2mabw7Lpg3rW66HDMWrjxZ
lBsZtQWG+U/vJ6mS30MX93siE2ntE19+5Ciu0VrpFzdI64FESttN5fbp6gAgUaKz
xXl6XimKinEj7wJiMGtwkhZ2ZAwhgAnLEgYbO3ylPhRW6qscLQ8iU61MjwRu8gbI
qO5bVf/x1FV2UUmk+HJZQhPlzO+02NATKU2Dz/owX+BokX+/Ctjx8xlbg0MR4XuO
QxGtxRwtjQxrpOiKIsjbqSjxDyP16iNmazInCNmUu8iNsDp/nzfm4+gWHevqwmlt
NHER3wvMFw7bZZQvYgAf+BrlLUh5Jwa3/cR/WDOgW0Us9TX4epZ4uIk0O9poJuZx
vlQAkU34qPhOq2+6CqgAur+LbwFpEgczQlVRgvxxq8iKOM/XobDUWCrlMnoJT24G
A7ubpssISseuiMiT+5wlpLniOTjQ4D2RK4OyhNwE+sklGPDPsS698nQHkf43U3rS
NK+2Is5loFUl6Jj6hVJiaXusIg9eZ230zqlfbITdssqfg4soeHIVzcWlhe4NyA8X
ImXsv+ZF5o+o1simjEkBSsODv9KN6Ip2XBXcjf7aSod2hz3qgvg8gy2leV2xY1NX
0wyF2S//Mbk8wtfqYJLfkApB+gbA9dLKeW0v4mpHk+IR7HiwFds70WNYpstuGgKZ
yULsA/2wTZsJLVsQcUeK52R02grFURRVfop5evvawVSKYx7EsjtrDrSFhqg5qRlV
OOosdmDYVVvF8gLQ2uRZ7nP0H//uAhV7gt9svTIBGwrFqBehqGycPNv6SWm1+qRb
AoB7M4ug06+7Rt/JwAcF8Iw3JCWBOaFJrlkiTKYvNVBtzXgtw8ttldntyY6SYOYQ
shmr83i1464KumUpWT7bMOKBmkL4HJg14aRuuNuY1g7KVutWfVBAOXU8oF9lu++a
kWtTLdezTiksQKkQzln8Z2kco+I23LqQD+TOAG2lWZuH87FTfBKeT1WPlmod7ApU
7Leiy+1S8mGqbmj70wC8nAyVk3tREwdjnHcikCF5JolzUPbLSUqvOMt4L9GdN+BU
JRNUoZdArw5kUm8iDcuO8tVzuyf1UrxRXbCAwM2h8+J/NYitLVZEx85KC+JgjmOG
zET0pdN3cVnf8QOg1veQk6aJhmwr+GXtC8h5+8MUUvnF+fu0EE3RSW4X5VeEmAwx
CWULtKFkgtdwZ8tW8PNBR3y1QCdTCaWPnbyvEq5yRsssUL2UY4nXZVUcs3Bw3iSX
YwcymkOBf1vnWcPr7FYn3VrfNSUA/r7tltEKmxHNtBZLKJ0o7vG4eNTwUa5DToTX
flVuFQ0J+xz3x57AtRTm1guIXieBeR2op1Qa8Flkckai461SbODshLtOEFfZxteO
LWZKGNLvEZhqWXbnyO5ehJJmFM7vbT38O/Gi3kHFX4291+3xz1uYi4LYje9mU6rY
F4Wcgftn7644fZhvK8s07i75QTtM57zf/Kve8ihJZ08RlXusbZqWJAzA8SMdalQ1
JkjKIW8YOjUjQoKolspOMTNmLSjum9kGQSilNfFrtFyLWxksX+j5yTC2Kr4hKXmO
9WvWc0K+wOEgB1ek4jhBrdR3lDuMcm5Q6OlHpzxhjxHhzotGeOmWrgYpvsYCt6zw
zyYOBPkon6gvcXKAhIS3lmpgSIAesuVN05ccl91Kazg1Hw147V6Qca7mSqRsSNo3
NtTIYrOJp7+VVEqg+57njxxlrWT4yQd059Ve1oonlBWEFAUOteg2TCnE2Z89BMml
HXuXDaW8G5c0hiWmv0cQis/56UIZk8DjYYOZc4gc9mb3YZEnileikX7ENX2s7Xqf
VSr4YESwrjPpy0B3kTJJROi0MSUY5fx87mmFi6OXaMgNTCvagKwmhLNLcsmoTAFL
2NceACQL16fMYmN9CPq/x4QEzhJqjF3hijJABT0ra7TgNQi/XAFrUD77ErOjaJ1v
EOL+4OpdDDHmitxfazWH/TLp4KNVWUN2flWZwbMqz2IdcSEfT2dGPbkWB1nmfEWG
/WWCcXOV5Oqq+/ssQw6HNMvDVU25FAbcMu9f9uk9J1awinxYMbspDpb3rbsgazfh
jertlbxE8lDEfbEjn+/cPKjwtdXyrFanzlQSD22r9f+vfWJV4v7/MZFzPjtnB4qR
92OS4guI39DpFE4gw0VefXmgI78WMMYOXj36Ccoiv47F1fH3gAgyGfVKeQv9pTQy
mnyw4MHCqee19uSxaftTPuUs6hdrWSXbl+1eSiG0Sapxg18H9/ai1QaN+wjt4sP6
8mcY2C2+ctWqArNAcu8HcB9uKMJN6WlOlqNYF5Z5rVxlhcUKMSLtM6twwKaM+gy1
7/3XONZc4nbB9+nWFcRslnZoajwBYA+3pLCAosLPYXj4JhutJAT+ZlX4i9mChvdt
+DUheP7hiu8abB0f40hCk8Gwmo70Nr+5aj05DINEfDi4SQsqsoQ9dCwqxe5gGoub
4u7py3MDpQhIgki1nRguIdmW72CaAdnw8Z0g/fnLLkqgmlR6Ip0JSzSxMvmIo54E
1MBXRkjY986Xgeb+fgTKcoXfGFSl0bthQ7iAWSrH2+wMcl3ekpOBmFeLeu5cgAuF
L3FZUNT4gpoK5/o57b2loGQ1pWR3rmqZrn0W1pfO0qzlz4T95WuuWJQMpY9CLHIw
zvRU/ZMkSRsSS0EngH7BPEe95DhJbOGAbh9akRSRXvnn7nIkvg5dBERguFJZ3MIC
RwRGC+6BgEi9ZgWLpRXU0pnSbjW0bbgcW7HF5T/wkDnU9sDta4kxrhLDNfPB0u8o
sKCEPjlblY6RTkfT302K7sNl7DIkrmwsKJLP988QZDdsFKZKsWCDHQIISr58+on2
+H6urXeTOlKzhwxHsqyWcRLeQDCPGBCjnaqd6K/7DZykmgZyUcuCjykUfxGYWvoO
6hW0Zyo5nW9JrLWDx1Lq2XQlIYY2O8E7+r85zSUvLXdqM+dLKmhqGf10NKHgf9N+
hJU3SG3Roe9DQ50jOdgcHfNdppZqxQfC9n+mcjeBdadggEzxj0fJtZcem9fKZpli
LKN8Nu8aUjBm9VEl3fiC24zqzXurEVvOMIIUROZEsNYD/vGQspCuRyFIbadzw48/
4nDIHIgZaIS0liUeBHyQkBr66AKQVLCdaHgmfh+STBeKyluVVAUlTweaRas3Q8hG
ZrbDWROAI/5AFA5zGyQwa4xEVpieK7kgZUKKm7glOJB3GMQw+S+JFWK6Oc6wkyvh
QnjXFmspUlcokEgWrL8G1Lf85eX7KqjMF2KRuNZ2CdIncSgH+Ldf7Zfe98DgRe6h
jE1ofFE+qsn9be1pfpZVCodk3XK3F6WTM6X4O0hqcgAGeR7C+tYtrdXCm6clry+i
bJFrUZiaDoJN4DsoR3S3lr6crEeSVl7E24BI+IgJnt8mGD+k0NuQeYLhs3U4wvYl
xdlRI+IwxiuSnAcKm5pDTgZ/1NAo4YKCd/4lo81kuEbeEsoZFEM6e43hq/goea6z
COq1EykS91sMywna8taFJC/+BpvmGEscC/jwfheOyLu4/xVDvmgeVPi9Hzx9lTEn
p4Tfo1CoECW8ZKwm9SwABGaRKfhDWPge6ac0fNbWTYtoJM6S5j/fidV0bC9hYCcD
OOmfwScTWsCByJjHx8dwYLC0DaqzFBlbIH4AiWIVuETH1IYTWEW7MzsFxp4lBxGw
rEKeV+rgXc7ot1gmh6Go2voscxsajtz4cDnf9eiza+vpsmk7zSX5515/zV/+Ly2C
6NlmqDDLZcaIri0A23p/d8nbdwM6VWfd2CaMeolaw3L05a90aQ6zaoFuzPBPeygW
WKmfs3NKOJdPhPvNsdjF39N7Z/RxcS0Jg2Zxh9ih0DZ4KK0I8BFgKYOzlbVZthoE
vwcOIi1y39ukIJJ8bcw1gQUQbxU+NnESTVd2kQvHnW6XZW1s8rLydqRJbowoW9Hd
jFnVP6kfpTHd4/yFBJAbeFHG7Vj3HfzxT8Cxh9KtfXU8l98nlNY7KGV1jzqK63TK
UdLee1XWnSmjpiraPSy4lM4UUwr45FiGvf3mWTKBOerTSpattK/o3NG1wK8iVDLv
yXlDb2EvAJo/PXmhLliuLyOO8RQB/7XT132rb9CtxOi3w3p0VDF6/RUgP07Ior+x
/28zLsswMEICvMkyvdurH4H4+ldpJEXMBNrndOXO3YjA9zH8oxmh7Fg9RPhZmdcU
eJtT9ZJRCoCjMwnDS8+qdqZo2cVRoennEmr4OztwEz/XvPL7eiSgA2/Zid1+GZq6
HYtkw4dAbs27B7W2fBe+XXtxMB81Oqe5njgMKUdQd7+18Ao/Z0WY9TYMKLLJQEP6
12PclN+/cXL3LwjbjIWgB2PoxHpMemqHJlXSAenqeZP6jSceDp+9zqm2xfDnDt6o
Sqmp5NFlEu7Y8wfz7fhEkUWkqx7RWSCBmfx842J6OYaxx6WHUSoGnhngC7EbSXn8
kaOT+lPNREnrOEkL7xIoU0MCTyZk6F74IHaLCZmX+wrJwBUXxriIsFnoQ13w4ovQ
enX3C8dcRMZNIk+7G0pzWVTZvz6s0k28asURzipSR2hNa9wKfA+DAKwx37qqH6iB
xloJrVXuFaGlVXAzpyZ8IOIKEiFnoSyNtqeVCkwWlagAUApeBGYQUVjyMq9/aOZo
hbJ3F0YIrLD95XDghIIP1hlpwOK0bUOIfP7OTlMkNfF5FWAJTpcjL5PaX8hkTka7
rI3qBSPz1Fv5mATmJU+2NogqWlfYdkQIuqQvU1VhM03LZx/JumZ9zLmTtHmXzJgR
k4MTN5cxk/ii8wRDkBKzVgM4G2veq19XkskvCkn4py9VLmponi4pE4w/Xsc5awyI
ntI7JFvbQSHCsdKxA6jGyp7ju0mNHaD6rGu7ZIkYNHPA6EEL5loLAZbhzU4vNHKF
4bM507vEROm/xiinHAcfyrqMt8Bj671Do+5YuPAz0aHPHeNPuoETkfFmKC197krV
knbT8VvisW0fHy80rxjLLyc6jDTIKxMRl3DY6Kcn/v2pAlQDIQuKGZzbbFw9FFOU
6XV99rYCu7naUiAEIBgaO1O8vTtkzKoUEY2MeE/2af758knR0PKDe8b/6WRjsKwS
1IXBd65K0kSo5HwoUp1Wj4Wu5E6MIsnwb6uqpzCNgGUDGRH1b3PUM9FsYGIWpONT
SJ9P6P58Wdvxlb7SCXYXlIWMj/SDUKGxvdxML9xBlZFtaYmPQlWY2A8S2EUdd8M1
mCqE0lz2hvdZKH6NF1AuuJVd4a81t7zcFL2VpkeBtkf1hdOJKGlNNWRRMhOhx1xR
26ir5ZbjqMmN6Z7NCupbFHKnf2CUfBqmnX+GXaohi+ClmOAMTcumZll0+lJInYJo
mFq2eLFsjt2TOSuCjK5rQwh0zbgN+iPbitvvoGbeNoWXYLC+rZiboGhmED6XK+eW
scIXnnK3k0XNyrcD0BkbV7mIjZ5yN3QhhUfvqAIH0Y5JvsGGnfbt6VGST06vXQp6
z1ouDoZGsgbCwJUapnw3mIHrz4pZ9lsQ7bS6BSFe4tNe7KwQlUMORhRFi0ewMykd
Q3jqd6q7wdXoF+PBXks7HjCjgzy/0t3mwxiC0iEImFDdRhBJtHR7nDsSL+pHqpHU
nZTq9Pogrrf+9cnuqpVVVmPOJNCMYLdRf6VsSbZZTnjmjo+ViGYPYmV+eQvpoTyl
ulfnPJ9KQHTKY13yzlWPF7kpoVB3gY2SVjyOH8jMZMQPNQJEBeaNSViSiSXyg1x9
vw2AOMEwSPW+tcJxGrCvLfXOP6U9eKS7c2WNRLoFWNTJq2V59CRfmLQE816CE4eI
HRxjK6HUFVxcCLyIXifmA4IAJcrzJPbBOaG5RI3UVgvVz0ONnRQKCJYtsMy7ncP5
GvZIpeb9IZw3eJGoa88Bhp+GyxDlrsLnUb6msxI1Pj5a8ehFRiR/kkcqHRRG+ijU
d7PI/hdqd8gQw3LueLBvGqnfHKNKBHk6g1b8s1oqO6qjLgyz8+W4LtHABgm3wqcC
nRzsBWDZx21CUDQWE8mHW1rsNUFKRb7rgJs6CnuQprHPCM4nGGQDBd73g0T1HOE7
lBv5PAw3bWKTmu0BDrJ5cg4xGRNppOe5/m8N3U7NmUe7KnT5fyLhQZfctttzPM/m
nissZlKhy888WHj/gc9OIFOWWm2ynJ2WERH5unBZDBM9QmhdXQ7Im+4PW0KNK3Li
ebCTGuanvmUnuZz+9TfqguKjvVqvC8FW+Jk/HbA6/9qLQRASd5L+ZXgdCQG89e8w
SlQvFdlIl39r7WJnmhjSwww9Tf2M7owjhrM0nGqxH4AMrEwmDuSOA35KlESrYmBn
HaO2o2XJIAO+DY3PrA3T+muIkIymbHQgQVwaaEAX/dr3NEAt9tOAdYCxqgEG4G0V
xFQsXnUIGqiFGWYmOAqABiIHKlHgBfig9aW7UcHY+2aVWY3SmT9VMR7G+0XgfJmU
Awk1HUWghYiohLmgVCkI86xl916nz9YqDOwbZcDO42pqVMnY7dY4OXUGlNMfBVsu
pkrfMYNrvC2zGgWxpw1+NzijO4FXwtlY43dpcOmcg7bVshNpQI9P0d+jQ6kAcT22
xEuDJAh3w05yItzaLfHm4QgIUmkp9KmiJMDFkeBXqS7SKE3KXSExzYC1K5fv5jPh
Ubgj4KWrZpLuyc4VbuRJ4s8jcbXCV1vLDpoBHxaKfH5DauTLmPMHqkbf48v8spc2
bG47qTofPl+XD/CaSVDNY6lcmAJQMWx3jUKs1Cxxj5sD9nTfQzUPoLDu7l2nEHc8
E3j69BXngFBvfM1Il0EAa/LJtoeZIRZstlqvZcYkZPcFOW7i1J7wbynsAittZQDO
cPst9IEvi5ChoaXW/n0SXADKgtM61iGQWegRQTp8JEcDrYD1QXtv/LSjD90WBCvN
y0VQpHcjC5785yzkz55bKGBGzQqQNpkbMGVVwnK8d7L9nzMvzVC6WDhmGTZzyLsm
4YPskXTDCDBHT6paOgfccVDToRLB4bJSRCidjozP4ifxNX0V+ak39ae6DeLW0Rss
lNmsCGcBbndWGV80r9ApN3wK4f90ACDvXJE6dWiAxAuOwDzjCVsDSZeRQXA8Lm9X
5dV+s1zXh/a9sxYxre1KK6srgoTmwWug//lSlNBs5bNEjAMwSHSyPEJKqFplbOAs
xTzDNypvo1+hp3YNGcALrViPpq1Qppn0AT59Gv1T62D+zSNnWNDWO/XVoikZbGZ3
Rfadkg6iEAA6njaI+wUH4BVYx2WAoagvXI7Z801cJtCNapBjTUQ9hRyhsqFXUVg5
7ZBRB8ZoZhW8o1ycf86sD8Mqr0TnI23vAkQ9fVndVRZNymERiOd1lbBFhqKXfgCm
lG9marwf1SIvJqd4LTBklhyFpLTt6lf6msdOnJyBa/Ai2PTAYgGi2eVU/q9OryZ9
vaGndwinpdXc8vq5qnutC4rw9SnM7PqaacYpEF5Xk5FkittoEO4yn6+/cVmQCHDL
8aFj08jPzt7jZbwk44Q/jkL9KoXdjMQ6zmx9Sa1Nhdc2CPde5onYYhbIxT+6rUag
4U/QoZU2qLkttTp1yeCHxTauPQKLJkL60DRsFVJu+FMOqFnOKQa9xSSWjJviNPeW
tSHdmdVLuTSgSBWn/HIHdr4ZFSDWCCJ+a73LBYO0NqjRSDCVNJLMQ1Em+Lp8iuJQ
WhYehgSdr1LgyVR4HVZRGg7fMOqZxrNzicbAItwfiw5THRjHyFWm1Wt1W4P5WMum
u5/bA7g8r3FFcfIVbiFAUfEKFDVdwe+5dxyTBI+J+cr9gbtK593w/1m9GlxhuWDC
jh8QSK8zY/0Qn+7i7USQpfAzxE0/j8osV+urT8QiHU09T0cZjAWSkuOkQnU29KVs
QNmilPb7I7aC9b5Nxa2/n+7tvFo+z+hnABWIJaJqQO8YwPxR5CPd8MvxMxFUwtn2
/e2HNvbFOQYWMvvg929XFGeKMiE5yfGm46owy2wrtVUXUkjMslOAmizAPxds21jB
eNacc1mKmHI95FSytnDMNrSnJ9rSD/GUTwU6JNmafCcEn+RLgHTOe2r+uv9FBsXY
E18Tzxk0IE5LnGQV0Vmlz1TWId9sjbIBfFvGNCEU/vQPfNZxS7BhrLAKsLY2HhCE
Rz37MOzcVszkzx9FDTnXpevzese6GQyeXti5Y0E+RUwfXBi65f+D+JZtoYKfMR/W
l9lIQJ5pMRvEgaUG2Ae50r7AGJ1dOHfWUl/Nt1N6Sdn5fJeHV17XiJpkQQ45HBTc
F3mlNuYfULKCJ13k1CRUkoH+jf3onAs4Gs3Pu6gZHFy5Wv+PxMyu4WWZNVLZuEuX
ToVG23+BFX3xf7E6W594KzCQNGuAgEMFttFY4B2ELplzm3Cpbc/YQ9dzp16LPkfX
itrBBkyKa0EOSnlfbj43mXKWZgP2Ki/yd0JIMtoC9GCA1jeNQ1YZAgsnn//1bzqX
9okeGuPNBERdB8wEQROX0vS5/GeFL6Ca/igHO32AiAc4XzyuDwtw8MH7uHtLJjOD
j8wdrQtZJ1afRLWibbDVnsgDVnx1RmA2qj6GAKaRDZdfge3/6XNoS2qiIhvC4zFD
Ktq2cmCbuYuPjvCFuflKLxSWtlTgcOqOlpNbmM1mtzn+XVMUtD6jx9PcFjIPOhxr
pwwGSD1ELhS/ndLiYu83utwcYv+yYcREGQyAizRlYV+zMjDgqAWA1cDd/X9tpO1/
kRAXDMMPeRJ5CW3Ugj53+jGjFIuLQEE67o7qivKkm4KGgdvGyrHBcQBXq7FHqy2b
mxw0jJiWQ3+PoVkx/rW6Iru1a0xeEOKYva4uBojsOUCzzG7598nIU1CCGnzcUu5o
1ebzmuhfPW1ssvPaGhPgbwGR5jwexA5/WY3C56VLweBnxK5sQuDN3dowPt5q8J4o
+h0qH0zbGebma93B6VDgBqUpAGC/U5hdHE4YcviDRf5ASd6pTb+VD1/M11yXVGHo
GUcnu/R4A1AVZBouqEi3WcmQufzKA6idCOI1ZHxeZ/oof7sNoLYa3292qBPwaMTr
nxQfXZEvD3AKvNXY2U5MzlwugqA8LHGlOk+VbFvs2NR8egIyUnskHkKTY0M+dZzQ
7veU12dEaDr4XmFxgw5QVor+8FbFggiRIvORLsLSSx6ihw4UNeJ/lHl8m4QKgz2y
aNB1TOnBVj3Vv/xncV7Da5QOtRhsQWrS5n+zNXJWcksjfAoLPZ+oe87FcpUccB2V
JFb9nDAEMc4TndTTkOzhCKz2PovcMwq6aufAuCfEMv9rsrcRNNURfjE5lQbupocE
sZRssvLlUjJXtxcN7maL8J1IIaCRvTnNY9OcgIdlaQMggw6w9IraUcD7497SQDz0
V97Y9aPNJWvVEPt7EIZ8eptj8E/H/NBAxovhrbB3oa1hTi2InbbnKNqSa/NZPWbb
KXXxYgr14OwWW0eobKhN1A/E7vekrl6t+kpTnUPw9u3qyY6SM/PVPfOVy0YDkxQS
NYWUYD5fVyqT0NwEf/uuP0ZKOzk2ae4X59dB5XYOTQ+5OKWmoRfEzXNSA0iHLME1
UE6OYua3+CinJD31JmVNj8kK+Ag6gc7YppE5cOtdSuarKaktNFrMaRFxzKX7gOoj
u4pc/BlVe/1wDXZ22cSJKREtEBkGKPDsRAEVB16ce0TCLGT2tK0dZGpCbEhVw46P
Sj1W9LmP41kdWI4to+eIuSmWhOMuFWazyXRvPeu2R2LMpZyY56HF5Oy6U2otWw9Q
VDkQV1C3KUJ7Y1Sej8HFayVpmnc6mxZwBjk0ELFwTa4gS+WhDvPNS5MqN/t8mF2g
AOSgRg/4MdVtrt2VYeQDscx8l2swTnOGCS2qxjUlQu5ihQwXSroMgCnv5/oM5lE1
pSz3EKSA8yh44GtdvFTwviVsWtpj4+vkp99qqJWxzSw98TQgOwXYOqCRyQR2W8JP
BtvOd+jRAIE8bZ5y+XT0gNK/BFwuqGYyL31VGd5Kyl2vaxu9kio3tUddPIkOf3OT
Hb7Q4doZYhJIbuwfckL+a4cMp/UpIZW3RXAjXPtMEC2iCsWS0iC2/D99y8VztMnx
n4G3ozLK2YByCEY5H7QtqhiXJ5sSiUx86BY7j/xbnsYn9sVl63CK0pbdW1kZChdg
7g18VjfxlP1i5Td9raEVTXf9K01+59iG30yz8jz67XW0IPcX8z+HOxm2uTAxDkB5
EbOSF4ahe1XgcUsczYwwd1xI8EAVXlZtegqyBcGBbP7tP79swA5HRHuD2MXdd9BC
7nApYbXo2yMbwdRd34u9hFKSVkM8ibRu7QjqdgbTjJ15OHPnmotnAyB+8g3Y8HJY
xpwAmsuJACEP4nzi4eeTbX8QwIU9LbQBGrOvCSpq7/t/WgL+Mxri0ZdfZjZi3P8v
CTKw6uqyZ5AYay6r8TPW5GL9ArlL7zNXno18cmK3EMODGHmDdlSU5F7KSTzjlXct
W6+JSOWfbr4VPkWKAVqU1K3BuM9TrjXlQ0lia2oXHLG+spwsXYgg2opih5qQsN+D
pp6xkDASHlwjDzN5Jan9CszK7asC1pWGJztIzPa49X73HwoDe6ZVhzFs8L0e3lqK
q1VSSEXhNy0lObWJnOsOzgZdZXFY5XbL2/bxeV8TDsQEPs3BP67BKJo7Joff/Ryq
GeEIetASr4KGL0xEhxlW/PEfB37/TLW0opPm7T429INR5hSzvP/n5afgToteDuUM
C+HM+N1vja8vHLe21c67r8YZKVxvtWCMZlD+wMXnMR/MdSW3cyR+mhzGgAZ3rLeV
p+FIb3xm0IWC5PciQJnvqDM8/41wI9bpD4zcXdzkozChJIl3Y+cHPSqiMkbzRQsk
IKtB2oDYu/h/Ft0eTP11+sjlEQfusuAW164uC8tn0mkSI+jnsITGImLY3vNdsKZr
7dAUw/NWIxj/GKUW8KQ1psig1ckzw13RYX85ZE0pikEF5bYZ95FX8vIS1at50tKb
PCLbDp83qD31Nc6xP+hPg47ZnCZJzkrVsEuQA0H3Xcw7xrqhy+mSYqe8Z3RP9gv9
7eEqLKTbsAKmnvGv9vCjdqJ7Un5kh9ck0EQcLWdEgeQCCW0MyllOytnpv+0oqVrI
GDfsHDsgQt4bUcI1WCdYPH9Ioaz6LrOO0Prp6MxOKH5abhnb5IA5DeN+S3Ei9dsa
n6S582TZUgOIsSLkGqih6BGQxd+thsm0d1ywoikDPG4+GGJa5bkPlWiCbQcBZw0e
2vBLS20ucGrcXr5Wqi9TNozwf4GKvVOof+HYcuYaKw6ewLgyMiaWT1XEfFO3r9RG
ziMfJEXRMjUnW86kajqHmAuk2wFqraxwzKAVMMqnm9n2JCIk/WvWbwuDK7bIEIWP
bnfqZoI7rYVJI2A8E8ui9YqbsHA+4Lqbi2WxrhnD1GAXPE62Cbj1ppTsPAJjqjby
h+/KDucmyZV5ahOOjXEarD7NwhfiLTRr7bi0R+d7mWdq8Vsuq+K8tnG+WefrNjZw
LkgN/nIu6Za89gc7aPwqdIls2rKBvqg2l4tP7bMeZ1Xr3wTARMQ7E6eZpQo65OR8
5LIzA0URZ6hmWmkOjwRKCIo/lcmYVb3/98o3CFzq7y9AqS+z8m2STONUrga8rsUo
3UbA7/uCPrv1icIQQBCfmSeX51ZN5Xjf+OMINP7mfrvprdiQj5y/INRK5Onm3SLm
kF4jq838ISTCiyZu88lYaLyduhvhAlFCaGRF8fUJC0J4qXtFbY/ncOcKrXXnwicP
fvkarR8Zy1oPnE6j5f83Nlr5V56ISgLF7LcWMuQXL1k/ZCpkKdCikKa7yMftyaDA
DLGsMSmcm7t1rv9tDDysNa4ZqWhEh7tZURgkgTwJYvyEquR1O1KvGuNsp9HblzWL
zjuah5qvqbRbLFl4ez0A8v803sStIA+fDp1ilBqn1ioveoC0HfkzRmvbaL9tTe1f
QdLhTcsSPcLnij2GffssHUFbS2ZCpe7wzKW2VJ6Y0kDsy1G7bwSJJg6xzQ9Q/uBx
cOpwvlSqhtjWsV1FM3TNnUjo3k9BRNYcWF/AFTaxq4eZlfN+cc0CSQ/ogG1Wzn3g
qdMHaXIi1R92t/O0P+fuXQbLM8OCjMRU0j7eGDNQF9IB9NG1IyDUFSdEqdgeHiZD
PfD6dUY2IgQX0jAFBvV1yBqIcyEn8bhzMIOUMR8Z1uGvJW1Cgrcq+LwwwRzt2pd1
pLw6ZrStYEBptfEZnD8RUDBKT+pPO1oC3CicFyBFb/1wQ/yiG763qx+y2yjmLQ8j
3MINx+L+DPRzKOrZKmT78pNDv0f9lB9Pgs1iPPKZrH8z6K3lPbP8IJ45l1PvMYOH
mvFpmYVRQUgHYAMZCmgPEmsvjDW43nsRfdbs54F4VbCQhR+D5nN+zWgIGiXBPLNZ
6kxFZizQLBkpPCr2hBk5Q32FXXPGx/16FNhmN1ub7E6AlDV727/sMLhb3KF7RI/u
b0NVva5qeOP5mmk1td07q3MCXtRRJGMr7UFtKap586ynbDUNz7eKbtf8aseMnspb
VIXdWAsacWoG7OOL7kggYifZdJDC16y9QIsex67Kt3NYxpcne/liJfRsFQneS9dD
HOLGq15D+/NmxSR1iUrWUNRdnZ4oAmVbmJV7WDY5e3vFFA26ZRF5X0O638Kg738+
/esbHiADP8F6pTLD5Pi4xQxDem7Mw7GkCSdbuRJZYqTpgvgo4AqTZtndmcZkKv+m
1KwiVULr/Fy0ZCeJzr9//hcEeEI2U25wk4vqxMSXAS+QS+0CPNGHf8Z9zsYDVIYX
/ksNNpG8Y20k7CuXuQ08gU8XpnfRtlpGYIa0ltjfErefCnD/KsD5o5lEOu8qpK54
V2DUWmufIjJ71D8OcpVro4a1khGJt8JNfKTYwxMdvV1CqQk8DncsLkkRNEWZvS/J
LvxG8MW3nzxZUYKV2bIlKN5E8BU4ApfJTySKcyMNkzi4IabEXGpLud6GR2fnXkIv
b/3pvBlFj5/F5LF5wIJt5hINXXVe3iCsw3hW6dbo6+Z3tkr3QCvi8Qx36kDBZxFs
ail7JSMI7Fb/P6u0A3owZ1m8/CWLzejDEBSfxxfreKa6GuYgqowuYhmu2BP+bmhu
4AbvxbPWxywbRKGI9wWJmztLSGoBnLhL+/K79QR2Jaiiz2f4GGDcfgyr/zw6uxsJ
Qli/wOfT1DgvtMjxO4u+MXmG+qhbJh4YVa4I8j0ggwILGCldpDact3axv9rF9vHs
1HEX5FEjZZOhE3S/PDXgr3W2+RiXXXPBsEn2H2bExJfrL22OcTjzk99cTdP2lQFE
aSE3XKiG5ki40YJoQjOAaIMicmrVgFdZRxHQS+jkggyvze1ukgZfigcm8uxRmO4D
X4yk2jpJn9/AcexqwhcNUKEf5jadCd2svV3dNLQLCkEBfla5KXjxI7dt1hzW77+2
EKxWqK5E12KbbYibVJQ9cOm3P8PkHOuXKbyru/h2bV8DsgpPONiKOdR9ZNXH2oP9
6ksaKtFe7IQGUYHkudkfp5to2mxTgAO02IjOB91mwOamF3vgnjcHlSH07URaNOD1
wLjT06GH5KsNifKfI9RGRhm9EOsnKZtD20a8ec33m1InycTfX83fDkUI6qtfHvhl
1meaTuO6r5wrqqbT3+zqOGawipJI9zbDhBfudFTINupfhuNn5f9iuhffcVrDMPAH
6QNDBFviWjGPqZ24mFpXk3xq36qYRmGzLaqaOa23pV+gRtBHDUXqZ3pTExz/WbNQ
UH/FlD/LYzYFeEg42ClCA6RLLCVp3zc2RiPdoFSsfLkjqCBD9XI/EEghAeQHtucc
OiKZplIHTLWv5Uigt3uRrKYL2AQJfzE7SYb6FgVVUCfEln7hm3NdhC4aM4qsL23R
X8WaV1yJVM5qREfTUwsEo+gJrLt6gQFkuCanX5LPH44YkikBWROXIQ6il9BAmtx4
IFT2zMWP0IqBJagyqR/xBBNTyNCG7gJItzqyxUwEgZP1XOG3e+S6MsS/h4/UbM4n
hs7WgqDgILP/KQATmVIrz4HKlpBWSd2TIvw9+dJymZ5mA4HxBQMrwGpzd/DdpwW7
XYyB4z/Ypf4E1KFEuvhhx+X3BWMz76iPkzy3B7+AerVT+Gv1rp9opv38SuUuJTvN
hRmpOUC2zzcuQ3OvIIS/q8S3rwt8YWr6NrNTMxSY7u5ffJefy54e+mjsckBzwCBC
psdkc/d7n5V+gRYVkWk1U9b2bt/ddpVrsi46qXDXY1E6RLGnHDPobobNAS/WZfhQ
ksb51ApNaGuNLGmeUMHJoliGJImHsBHJm6MJUZvS3wkI4n2NoELDJvci/JswKE12
JPXQ8KffsjGv6YZKxji89W/HwwUAkoBUUV/DBA5pD+SJrP+YVVd91a1lBgaTuGKt
HZwYRtRkTMdrS5RH5LL/Q5xKz1SlUpUahQRHkSNoyRFpIF/9oeZeYXdT42oYRW8g
BnffjAASoImszPrt5+qL5gjLw2dvDlzsApJwqKHSyuZPJb4IF/lQyIELpiFfkorl
0DkkTLENwkrv5gXUACC2CwhcZDsbH/Odlu+vh+9X/6+MQRLFbHOVu1u5xxIdcNFR
ns/iFf5Otr0DxfUgsjG6ccAwrgW1jKlF3NfbArAcTttWR3lvVby5PqhTaPupEHW7
Ld8olkTC8GHqPWYq2f2q8597B7XKFVK0I1dmsfWl6ZIG8WgaLZi/iyzWnKdFpLow
MVx3Ej3MTfhRHnpTssl4gFpRoo+yPBVSxLI4B+hE+xD20G7QoWV0uOISRyUegaph
xyb3tiyWHulDKh6jxOL8ZOw5zS0AojTRrJ9+MsrGhYK/1VS8OLVBCN535gaRtJkZ
LaCZFYysNac0KUo+iciAeOyZozJ4tZigN3GQgFXjygho3/5Rj42na2MEk3T0MKda
RyDWtNJTScuWsRDpn2iHOpx9ujbSK/YXHGc0T3701nidM3i0kxCwXQatQ9W7UhbT
4Hv/J83YzmryqeGgbIXy7lvuzGvNmXEciEwY/uFCMd8+Mp9JCPmvyeJASgDFGQfC
`pragma protect end_protected              
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
lEWs5Tw7LvJK+sVt8gmTpKfiASXEbj0fwkv2Y5nfI6v/N/K+oig2u4qhHFCYPUgO
T/MaKNZ2ZWNF10Tk8gjlN01rIdQgGysXlGH8Eo41njfpO3HAboXKcreKktfldS52
x/OD66Zvc6zPH9Iwrk5ngX3d7IQWO+c/H3ZOUy2utXo=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 122934    )
xY5w4rKGezo/rSdRqUUJC1zpYkY+i/XPvvqbUAtE7fWPhNxVVe8RHbR9nPSUl5jg
SJy14SiJEWUhF9CpjJ4j9SQLLsR9U4uN10hndzxW9D1qDjP1Ux5dLuPPhJEQvTLP
Cl/ZenSQuu+jVUYsrBOfv3QzZxE37LwPuzkvjW/RVuhW6sg1Yz9aaT7c+bnPQRbc
`pragma protect end_protected
//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
FItBIMFu0EXZM/xPex+StdgJyWBj2DZVng7qjeqwDTSs6HwtBOYLyD59pC+k3Gde
nJrBo56MMw3P/GXG/V4CLEqw/doK7YH3DyG6zzhJzb5ocggQH7Jtw/TZN6dLHH1c
AsRNNw19NA2QXxulCDVVAuZFQTuhndT7B1imPqxgz7Y=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 134862    )
CV5EMZfnbYR3Dtu4Mgn4ubiktjSS9TykR4P0HyZMMGjIfBefPVg/oUpS2yxhP+lq
LCgOmJF/jkkamz1dKAKEtQL5IWOJKAFUBYHBdMOdhRaGhwcC3ZKdr7WgVH5+Ni2M
y3T1siixMU088EHfGk+4KYoXidUO3hyjY5awWcVoWZ8db4sTOg7reiwTOKFX4rKU
AKrq/dxE4377iw0VJJNjwP2gZ4GvY1KXD3tcwOMr2CeG0gPrwwQIkX2aJCF9DHpJ
7GhgeEwL/tp/O7xUWA8Ma6NSYULgrJ5kcglOd3pYjgS/rMIznjPtX7bLQFOiN9e3
93BuNk2spNXh4DfqSS/LmnN75ID70B3qF1guqwVcK/IdMd2vzELQWqVjUrDJSh/M
tMj2EVwkXtxSKw2PazR7cRiNffzg7ge0EXZIKYzJb4MLUqXLPCN1O2dk9ScmpLIH
lxcTycWPzNxT2wnu7U1o6/frPeTuyGZhVk8U1wUeK6134209fAk51tobhBfZAg76
1qO+Za+7egcRl6muUx+mA8QDTUnHgje2F+d1Dscr38e8Xiod1f2b7uSH3oQmBqSG
OEHklSTUG1rd2NwRGianpHakal3Vtcv0YlcCmY5JYeBPTs85+XhPC1cDel1OMNj3
8qQch11qg1s4GfayYWFknBsWXIFQg3LDPrYjHq5c1YUJYj1YBThPSv6w/M9MOT/C
QN3naLgjeLdq4wFFp4+GdRNQq9DVX5seQZrrE5Z2ySfC+aMcU3IctIDQ1fVvUtk4
aJ/hnMXHCjuZAI23ujhkg7ttLh9KtUy1QflBeZ7EMM2pCHDpzstbs/ee73o4DCZr
qpQvWWHssxHywdSPnvBzRQ1eayucIZgeYT8qwVptB0DVjyBDq7ysBLNJmlv1Ltbw
/DEGQSJA47L1X6wHDbTo0cZppqYIRtxkaWupdVVTiehsTeKctlDfPgPfrEsMp7yW
JskDcXg42X+hD8i4X3LzFu1Lylzfs2UaLNiuH3lplMg8owFZYZkFW3/aH4B6GH4q
NwH0s11zMpEzwjKZc/eHFRCI18m4TVUG6qjwwabG9Qv1HUiRhHuwX3xXRDODvpLk
ulfNlpgJMKIc+KSGrTMZOZpQGRJkJCouXHy9LXqRxFWbrzaMqNrWTu1lv/cwOadz
WR1warHNIIY7tKA+i3zit36R6Adu+DH2bOBnlA7IznFvZ9Yx3S/Jr8syL8VFtoi0
kvq6J+8cpnW0jzoFJOs5949yAzkSGkm8SOdHduUbeBzAz7H8/IPYTAHv5M8E4Go/
7Sf9v8qt1oIiyx8K8aw8hUTnivLPYlO98+YulHx+RCzSrC/H5X5F7383lDy0guFw
I1UIuJotFgYigWPqfDKTHx1LIEQfXUTOYgtdR59q9aCH6l6zIuWmYMM7b3OsaBMP
HbmQ0TwwWEMr0A9WbzRjeHGrpyat/Dfhz6bjp/RHzEmS+Spz+pRsIKeZlQVSgbfh
uunhKxDVY25qdkqwqThp8xpnkkMxUKVJJo9P8YVO6A9kYz2L4U0JVwsQUn7E4M53
2RZbf+oVxG6dM8CrlyF8tHyPG2E0BjnaToVAOvPMFJOwAwxS5xcWI62WxTSdsq1L
co+8nSOwLOJU5Yl+DD3aoa+QBVaDXteulVgJxbWz+Raa8C+fL//aXGMeIOCRvA4f
8ck2Ud2CFlvGsOUMsOvrfz4uoyQWxAmYd4BOwJxAjvtoSEXkNJt3IyQd6rAkrFpN
RG7d5OVoyTF4ekM3w727CHm7/GfXGx+QVHhQkIztHHfLqzKGsCc2wF1kcpTglAdv
vhBvLou8tLtaPt1ZUuVFmRJSObt2Uwy0sZ5/+YwhkG4aCVxbdEGkdqQ7WRXcsvNB
YdkS089tpKKJrAaQ9sWQyGwYzcu19qczjy+rXKtMBpnI8Cli2Ia1AJzRjTMWbxrG
vKILlXGueTW1MCiB504IJDlBi7i19y/aYnbgW2fFGlAGEbZWH0bi3JV0mf5MCbWk
j1kbh+blkcKft2A4lLpaW4p+EfvWTnOYVNp+SYbQwwQRqrYsNMFsz5/P0zXuW4ru
Vxg/Z5WvKKVcTqvJiMA4sHbb83l6ChiBy3r1EHwQdg/HcoqB8MAkrc6+708LNNE2
rfPT39bpKb+lXuTI5FUiRcoU1t8D1F3zDyGpjTQ9qHVT5CBvWEdYd0USrfdt1aBg
UYftx+N/br2w6CMa52Zm+tPUW1mLsUuB53liR68GBS9KGKdoaF/vliL91hdNcJTx
QKx9P2VBPr4f68IJJTKGn3t63Yj/Mn8PPCGO5Yy/wyIvfPsTbkOZaHEj+XGIGeWc
1jJXRVjebxbYwyiyurOwJY9E8QniztiwOTCHN6y+zEiMpUwcov8CWcgfFxF5LyWv
NJLdt2YW1eEhgkioa8yAacI+E5TDZAQRiIO2RGQJnBHTJcmefnBuPeyDfEjcxmv+
hVjLYLFMNE2CwxS5hNOwk6+hlqbTZWLKKbRwCPvbWsi8F6ggHfnLMMmqPnS0omTW
o2LGN8Gl4bGiKxz2GqRGYTSuY63u2/tsPzanprobFTGEmkINGAiv1kTnE+z1wJAy
CYhN8mP1esTxyt4zcX2gB2CNdd4OGYcxwnerUAIQzE9gH1jZPeZK+Ceri+CePbxX
0jWSZCPMjuBKCC2Nr2fd3uz7pEe6oae0vHHkl8lpDHZ29+nL2lD8pB96mAxUHUmB
GWPM4rjV90pciXrLZwatIZiY7pQu+LSrx3pYd2BHESiJkJa6nhHTI9MeayeI9FsI
XsUogzTStUieJ5aeYUSq1O/e17Kj0Fndc4yum/a4b27lgjtMxJtwg59v6aS9h68n
gviRj96unYfocVQUx2UNxou4iWXMy20VJsjotqciVQqmGWpiIKIZ+NIi0FDNdc4H
A+cF50Mmppv4WzJMaZa5dGubK7LAqOs6oVOlzsHK6lmVBvepqBsEJ7EFZdApPPf6
LrhbnhDouyO9jmDsZSd2Z9ohBrH9c8zI02blZEmcv16s6yjBad61jlBz0/FCdFj+
4iKW7PzbjXvv+ngcVxFzbk4JhsUI5TOcTTSCy4MF5QhgSdNcuVmddPXoQ6UML7Cq
mAlcuUb0dRO/KrqVYB1eSYSXCbR3FUCBTLXFe/Wguk5OPMi4B1MG9b51ZTOmMJoN
OGSACo8HcLEDGz7iktCDXBeQIk4fEm6Tq4HhBPWKPAwxtcaDWpE703RkVX2OnZcJ
De0AkPXgd8f3+1VcFFlm9FUzVp8MfRbmTXrDXvLnlUVPhNRelYsz/dARPVyyx9UW
0Kf3rR+v3M3xyUM6kO/7Uzy6+E7q5Bvvy5mRphj6IW7V0fduhIFCROnib8H820R7
0pmIX6jQO4Ydi5/noVT2T/pxbdlp0GbStHaA3tQPEOjG2F3qO+3PlAEGDGtcZmsH
7YF+fjEXUdmC7UW9YcLyQiBNzcE6A/cwLLQu5uUMh0Ghxra0g3n9aM3ZZZ9AVGGD
4NuADC1nmZ3hd/kKMDLBm85Vt3gk9x3j30G7HssRBfOGUKioKRDcb61+5D2a7Wv3
CGPQwWwzvKplXYO8Hiqf2Ct3Iv7ESFzMKqEZDIjVifNrxBP6emL6wjwcTdB2uuiP
48DjvJsaONEj6zp5fYQFARPUGxLDcJMzjsEoRS/tT9eLFPEQ2rgKlaerX5oNesJF
t8h/EzpHBbVrzeHB1WUlolzMFe0pCFty9Zu+ViPFHAmXqpO6wFAxhB2pTTaeiPQi
IXf2xoYWKfJdlmcoEQNl530pMRht42NY6J8G7YFveHRa6nZ246lic18mmUm4aW+5
3YRCSvGn60WDImnSuO8MGlhySvEgzVqbuFUwA5QQjl72ydpSEjSIQzctxukA57U1
6L6Z0iAY4YrCEZlJnqXvI1nzb0aHkkYWGSxxiQfuek3hYC7kSBXRe0BH01qnB70v
YXCrRJbnufsVxukBPLvfrYVkmKePhJsLujTYbSZ2gQ3uvzyJ8uIuLBpDX0U/lVnn
lEDtU4gTkeSPiyv4iOD/c0V4A7CcSCHJNB2yPoy/MRezKIEVYRyW2UrupaRy14GD
i8NGI6G3I1TmjzkbPAHlJZWolIP4+RbWH1zCi995XYcpc13ylrRNx0KJzm266wu+
4i5o29o5UjAVC2vAV4ufKFxKVRhgz8SkLwIvh701YWTor97ASDoputPTEH1F49Qz
M3LYPcmU/fh/66+inPJ4e4Q/sj+CcwBVYJ2Pr1lNo28UtvAckxbqKVshH6r1SJT3
0YoN+CbiSA1qEp+fK5nSyMrtrqOlGEUodNlplM2bI6W7/LnULfy0Xs0GUiTWSwzP
OtleSW7eyatJjLp2wY8saJfdHf0ILodmNKW39FqdZkC+hRSAPEFGCTSJl+qoubmv
qGFFYTyZYPeuLovyE5iVyXi7BiwHNoQ2f7AvEF0whQ4YPpGICusJPCwLOPcU3lyA
XcqNDyFvj2nEDp7ljB0n7Sj52DrjbPmoY9nf2hGWRs+hmvh8Ob55VsDbJ/JAW5kO
RyHeSSO8uNWh2IRkhES2lgSND7KkgbAVRQRJC8wpZeKj7hysy/9IGS7Ixj5CErxZ
GsZDXNCCV1gTioyrMZInYLJF6WR/NuZxSxk1WJmf4hYvgsZN/dAyq782+3uDRB+m
pM+8ZEBNfu8bGbZrpnwAgu6F5tZ2OYTez19dvLO30mcbIYjrPswWTDH5l5tIsDr1
ksJIzJrGV1sy+XB73kvBPYSxwhtBboTf1oqyUs3IkjUSr4Lduu5OQ1WJrcMegrq8
IZTao5KFnD/QGbJjjKLmfaRCRVuuPYgpk9qrMgVWmYpEyNeeaVm1Dtv36579diUD
uOl5C43TLdAewnTlyc7oFE6WYIB6VY5I1kXOZVfXNwzO6WUnlCSAna8zcQdKhuqC
bmeg67BrCHDYX6HaguMn6PSZN2D1KFZ8zBuvRPb0J4e1L+OOovL5CPT4W7jB1xcT
jUu2TiKzbTaZpzeu1vTGaMXU26qX/Yj+UHhumXC0aOvu4br2m6JkENd/iV2lCvSQ
GwtvVjfhMZzMto9GCvFvjDnEJ3TweEQxkD6jHJy3OwkA6TnBEQP0zfvBM4LN6PT/
rorgOCxueK5aTIpAtHpM5YikONLVDvFhLPeZI+Cu9sOszyxY7quSFwGjHKFAZ9ML
1bJFW0RGKI9/mPlcsJhiXfxPNDMy6lz1af1bGIMNPC7JW7WT6BPSV/nVl3clrkMa
1n+4tcWj2mln+aZfXcRi8FmEuYo0gF5tBJHOcZaEIyXzs9P1GWsFwBBb8pGy6nsJ
PZVWGqBdYyqAkuWhkUWz+1c6mO1K0j1+2G8Qs48KhJtN9m1NB+Lg4qKsyFm0WOvp
I5bRdzLFVnw/4NTmZFL+VIECX7uiswhjD0sy3/ta94+L99o61K/9I4mA5aDVTTH7
l0YkO0mC6Bu+uNpYiu6PYK9gpMee3KKnclWp9bswkQCeb0ffq2gMzt8B0h9qBN9A
yogDV/KjEiyF0QWRrGUURIhZM7oI0s3Y0/YoCDbSx3D4mhTisFw1x9WC6ocM5cDD
BZv4LP9e6a7ZnP5JnsFNEah3dRtm7EXknkQuNrFgYMJvEUbEx5V1awjAAxhFXe+y
OF03/TmpdAkhi0WgLVsPpSfNcSDj9tQ//A4EPYsU0DT0p9xo/RuZs8pV7MRr5md5
vZbpxM9U0m4ABZY5jDZcGFualP8OLV6hk9WorbZESCoguu3noqSDyy3RMQiD9s+x
08By8C7/RfSrGO9evUA7WjksYFCa5jp3S10wmGf/ovNM1H1ZM+RBu/jQtR6nx/Va
E4Se3xW9/n8G1bGLIoOuubqkQJ7TjZ2JJDDzrykHtLAfmd79lluenoeP0cEsRgly
Jj02eAf4TuLr2HnsOenuzwn7T0Lo5QG4lf0vWgjGlYP5/kbbL+F5zUCcmiZECog0
+IcppEYJf1raYUOu2Xac2ZEkkzdeOKjfTfamGUf8WzsYIW8NBZR9Jow4DDoXOU5F
cnll2IwjM1NF4KcQ/qFKTQxwFKoQHd5gaqweKhCw/CejLvQNLZ4s7K8MPyOFeaLk
NFL5I+atkXbgEdxSV/Y3laLLp7lzjlO+vLFE9gaVZnK4KMDv8UrIoXYlP2FznNGh
Jo/H+IPl75DMNXVFksNZgG4IuZA8sRXbyptptfclUSqQeTGguNtvNifnIkOszetB
4BWu8BF+oyzJIoPfr8ufjIT0orAs49XjgYMNtv6lWBdsL9N6JJXwrx+ocItWQSZN
iB84cc8EDvQTesuYTmOkBsrzRayVq9Nhw+krFQm54hnEQiLPNbewV9idD0iErTDC
2YT2Bkl23Vt1yPYHzLnodi4kyCnfudgIFWjlkojSVkoDnzg3vIovVHDq86Ds5oAC
8DDGjdWO7+4YKBzJv2rCLf/4ANR7Oc5KjHStMXmL0oBAk7kzd8OCsI0+5aRd0BZ0
08yQfwan81R5hTTmMr7oyJh1t8hzSule8OefBL4nRWPBf+wBZhiKnUJQPRW/b+on
kwSfkRhfzswv4c7EHUiyyBhclASgPSxMQ4KzrrrK45F0TKGIltZ8j08vBJczvoti
SNdJLcIpOzwNwe2S60Qfd89mG46oRqIeyLVBKYC5PudiOZ7fvTAMsk1Tanxfx2RS
ctc4xE60j2YQ+PczPcChUBs6Dxjq+NXjP4NL30iWrsmTB4AocSJ/SiT7w5ExTSRe
UcOeks00zh0Z+gW0qImI5eDLJK9LeROGsUxVxtDfNB2atbERri6w1KyV6Nyn3+yk
j1Nu//KEr2b/UA2vEzH6zL7UClMlZ7cEPLNmbW6igyKE/zpeAYXYnz53sk1PjCiS
phGvgc9HFCRRNKJhVdUSGWXOEmT0QJ6E5BpqR6LBVeWg+6cvMcvvRWBwNpgmlbSC
uJc9NI3iJE5a7gu5PDQzq6J9TNu9o+42D4byF8+F/IfmvcQng3V4blRc8oVYRBMA
tDOP05EOr1mF/sR2kaqz5pPEoRD4LCLEjOYFN3MfNj+VCiEXQjOL3jZcJnBNjCgn
pCoTBjqyI6DGgYVNksKeD3FDKOncgHw7JNGdWwGv6AThYl5dU/R9w9zonVgxSe0z
zh/vU3NDb1xgsfP6xIh/KLSHGrFK9p+Xfr2mCrvU0D9vDWDTQRkvQlOxHf+GLUHy
avl+VRLL/kJUM6C1TEaNaNBMSSTBEqsiAeFpjM0UA90myPuTB7U3hPQbgaZufPbb
CF9XGGuaClegk3rdLXxvQH5Yl0htr61EFiMLGnlLqWyc10AiQQnoUFBuz27e02Qe
qcLTTSH+o6c/fPAFtSogzWeIxQJpUiS54OiKJwuepZwmEYSjUMLJsommIKzRRheS
3MnFjKxUeCfbaFJ3gJgMsFzKSgjUAr0wN7tLfl9LcCz77PjEBOIMtZulBKlJ3Cyj
dJjjTOpa/oup7G+YpWN3fxoYKRAZ4GnSqAO0Fvxh/RYmkBwCWCs3Nd+xQL9QGcMy
oD/8bAxaPnT0ztb97/mrOqQyBbHdOOZ2fR6YS6aAWcavgpaJw5ezgE0MyCf3+1xd
F2T4yWSI2iLWBjbPr6CyvsdTvI0R5PLmOA4TZD+fZo7y37gEu5FuAhyNkuHoMcIh
CBjHM0sPsjZU5U+WfXYt1Bf5B3tpDMxTxqp1Pf6sGfNXdJiiEJyiVRsGxifmWzWf
xeoHvXzJByGtW4Z/mQaOMSS6tRkSHfhyPDZNophHQRsrlHuW55t9go9T/hcZwNkA
kH3kzXiEE44RfEM+SMTjXHBdugJNXzM/7LDJgUddm0zVUKCot11uVTvh2HAQdRZT
t/uB1bLLWBI2XqwyjSx5Ywxz9b5s9iE4+N4zJM9cG2cFT1l+y/sOKnPEsR5TY67x
IaARAFBjNl5DgszBYToKsWCLVO6Dy7AL0cxf4wRdiFb5eA49o/Mor/zXU1pYYcNj
GxN/X9SAQFtR6DTDZhlEExSFOmx0kUlen5Rt/1mEPMSXPeJjHLWUmQFRNPXSxdS6
ldIlGbNoTnlmomatgwekexFJ3DFD0ScpoOqbsitqRHTFA8xoa0SyfjKX7O1+IqyD
YxPT0/N5z8a2iRH2zOTqSJBJ1yTrbGpch3I5cf8Q8FlzzPNLSneY6sjynp+g1+yB
IcITxTMEO8nl+CDsN5HdLxr+eUGHkjRe86XNf/sQn3Iftk+h3ztB1KnWBBZAC3fb
Xc/vQ8+7qVwRo4Rous0/LbmS9+5dcFDnyXNGYn/LD2M5kYm2vFrw7d7bBqNLsGVZ
oslF7vHAp42PnyGFjSZFUbhEYbCSFR8b0WalV0JAHlRozqyDuEhMW1zBs1JtUOQb
99RCNxWqN63SxE1OdRgat7Jr3aqMtTKhd6N/hapX4Uho+WWYMxKgDVlBNPPrLNSO
YjM3SbYgaCjmJYW/DI7Ji9PBBJLEBg6cKjZ52pqLPxTX7C6LFX58+mCOIl6LIz1S
X2TS1GO7Lpc4F4/hb1gaUOpkwHeyIx5Wf1rwJZAQxbDT8saSiPRGbyT/6/oETLMY
k3KSPp0YhCvVdcomnnORA3JYUCHSOYoOzTHIMxWTED3kjTImNYaP04t/YxZ95ZTl
ItaYTRzKoL6zcVIcojrJ7Xy4n0NNvT+kfqLXAYIgRtEdkTIXj0UGmwJZYMAXEyWD
/jjZfBryO7mhQlUPwi+kuyUldA4Uqbcm9sENkxOy64zNziK4ZE0odOhutkMP5xYQ
loP9UTkoBIf4lg+D5J5KFEfWiKbr57s7wSUCN7OgfAKrfzl0ZFpc9/y0d7K4ZN+v
Jwncd95SqHO7Bf0DpDZHlNA182o+/Jni8ObTopoatIKBLU9REMeirmrCmvnS/RrF
99VDFZC5qj5Bt+EIFLCMWStXJyeqBQlJF1N+73MkYfI521joK+h3J/k7aV9+C/SL
Jqyj8V9ijHQ8zOwwdTA9qaRogsxk73kX4vAKTvCA/L78GHY0trSBMOQqhWm4OS4T
Q5PKUm0ngKyDYB6pCB8ZHHn+5kQq/BKUnQPhey9ccyBmxLgFUfehXIkFxYJOsFhd
NLPMGPG9PUrADZSR3B13h3NGPeJYBjp2/pP9/dd94QxsfGyskBT6P2XQy7ZqWwK0
htUWXrBiAKZCXUrjbZCeRA7f/HMfqTgMU1PeURCBsu+BRQMvDIfw2Eksg5Mj5UP3
1qxXcMBH26yIqE4ZkM/E+XFHJgpfgXK8OwtxBGQIL7vsYDW7y2jY8z19WXZNl5rE
rswQJzKWMb2g521uno6TPY5p9BdSoyKd5zp87KdluiziBObS76BIPhJUhgBHrlOt
lZLvr5rHqMxs6Z+r13iDAR9BnqhX7c82GYsCIoeo9UAg6KLFFZxOMrB0Qzmt0yDn
WooZwpAWk8N1Kf34x5+RlNmAOpLMosWFZC+zvkM6KTcAYuLngi7M1rlFSAdPPKCD
GjyF5ponS5jQBRl+WUspGZy9eeBmwcq7Oith3FN/IDe808fgnu6TGcxMt/XLao9n
jMjgVDi3Gc3sa+KI4/AUmvMTpS+LbMZny7Jde+9/x2AdkYQKQaShSozb15xqw405
5iyKa5zRtRx/vvo4yT/fUEXOwXkCpL1gIJivViO3M6hmEQQh84IqpQedxjoiPuHn
PvGrtNh/N5NNHoYTZ7aPd/BIvFq+/u2jQ/wrrUVuiLxMnWIxMMNYfSgYa8nqu8uK
y67FemTdelgGYHFEhUYI8Rflae2FPcCSSw3xAdqzAploK5EaKLL0CSCct842e2Up
vzrWh+JtStQMWa4yajZ8uL80+/EJJCOWn9hR0f63kolCgN2beXkt8X8C0mbk+BxM
3Olcxlp4SlhkMYXW3wvg2ITcShSP5HM59999kDw66c4qVtk92ujoynINozY+rUvY
YbsgGmJyIEE4KMtFjTYNqMlZRtyjMNZb7EsstEQGzX3orHHjmJbeSLLYgknJkWfW
9ZaKBybRzhQMKsOtRBrjZs5mgfQ2qkJ0AKoXeOCFpsqS1WjF9TQPvAIgMMu7UDyK
eUQZfBNLJcn3YOz1gPGfxtPEOfCnoTjryPqZWyAUjwEDyPdhTUO3v2POUvcMsBjA
p9+2tKr+RgCfGaLAGBJOaypVZNMsyiSV03fJFnRp6U+AbKJRIFO3nujPA8QKYW+z
o/ysWL59NlhO31pf9hS5vVxbh5Za2d7Fg6hlTmRK2vLvEaQfOzbra+6uf3aVrEah
PNAUUmaBxf3fIq7IODeCYw6PRfUgI3sExYKl2dQVaofaZzbxMBM6GGKExsRhhvSE
vaaN68dT2sZvqUyMMp8LINu2B0HM+XN1wkIQHbrZVVhLp8QVNR0F6YWPHzEFG6D1
MRThbgh0esQGZ8e1jJ87Usgoz1zms8I+ABPngr9vsYrKE7NnGVQQEoZxtrFHnM8X
/RGxXCj0x0flZ4p6OWcKUoMMfVYuPzVL79JL3vdp2I9bHNiblp6tPAYId0Uj+6iB
j68Xul1VHeSfCecorG6ug1T6iLNbd8HcQ0VxHFagX77lcHLt1K6cfbLn+UkVc1Dk
T+1fdPWqaX/NrKxL1vsllJtpw424dius+PGyP02aCb7Pb9h6UFjrUTepskQQHcdN
SqPYG3IJb2NcCdyiIJ5kJXIVTe/j6Adc8Eq+Huf2X5zA9gkhM2+Xj6GljXY/JOB1
jSlQccBOp1QGgNMGrYJkB8Jm7ODTnVT/OlScXQoq9JnFqCAa3QEDMjm9woHj5mIT
5J1tWn6hJSRMtXsABOt8t4saPw04LMFZzaByFUBMlV4femlKcjyC+1k89xcK+N9z
EHvb3McMPrxCAkHjsdIujjRKHCFnWcOUE6D6Kwegwk+lyI4TfTJvR5Mz99O4uBKk
lzqll+dfDujRUQAJgrCfMrdgXT3nCFoweBTFmUgr7nkO4kmyUeFLEgXoBBK3LFfa
rT7OlVG+6JP0ZlXUtlRlawj62dCkpwlnB2+IRJC+xqYUMfvNN22+4vhkNRS1FhdC
Ftb8T5TOcc2yTtrsbKxsN9eEHj0tezN5myZ6tzaobxULKGgLM8fNqSCWfxT6nYD6
K7Gkr1yFXOfjzPPTxmG+fv5va0k5e0a2bmur611jkfKxmyVecKXmPpp/AI9eonwq
V6Si5WNP6X/TTdVFAO/13NYmFSm/WsvcETqsONE/f4uLsyb0pcNIDcKuRD6FUm4l
yUsjFmOHbbawZvaXOdsKFzzFc572Kri+8DxZfD0+FOLsiwXtLF4wCmN/ofr8Vv7g
fy6ay0Fa95JvoQhFqFjzfbJlXx2VYQzRzHqfWqe3zyXYh5yMUY/ePYV9pWq9NEBL
fXMcKhKsOVcr3rMxx4D14P1oV0Wr5CTdZ63VIDccVSKBJsRtFv0wNW7UKgSe5qLj
1OCRgHsVQy0NkRgP3e8JaWeRHQFT2ygurGDO+R1RyR3PK7eusiuUImqEYc4ZHfdt
w+ZSiToitF+ea66Yg8MmcjSAUA01C85FYNJhPHur6+OGIhMQhaEmWcbMCn2VjqCL
luMN6PQQ/B4zt9YA+VEVw88Rt5i8/KVL5eVBQrKh7Sqo24V0VsaQcbXSzlkPwCeY
e6b0xdXe1vzJTSdufnHyJjit8TWLrGkKbKUki6XSBsZXQiu7K1i2GrjGUM4oxKPm
rmDc9vQ8jWKCFzXfohqHqXXTOrQ3nWric9xyr9Dorqg6gHriyX8D3zk9oE1mRHwq
TN917OfgXIty3+Mfiu+HQz/SAHjix+5Q/yRDAAKgtc86C78JyeP53gt7r1WfdH6H
Tt0VZ6OyPlZQL4JWusotPdFy5mDsYs9f4RHF5VcVzmFWxitzcYbYrAbUzI+K3MtZ
PJbk4Wz17wQlZJXuwP4iH+TKOorO8iunEwIgT7RfAxJwOniBFTm7EReDXhTSrX2T
VHMCtBmBjUhnbVQGq1N8ymav18W9btmWkBBzYrKQq9ig+yfFx2tQu9yzl43umAd3
n3prdlwFFY2I4JKObgGiKC94yi+OMuKo7XxkYT03C+HZz575JhNdAffzDuRzDHmQ
iFM8N3sc6OIyINCBZKwMJKajg11w8My+9spO2xV5xtC/Z8utCEWK0P5nHRv1nrYN
7zrxWuHLbd3cF6iYWVC9D8GUlxppSM80MfiShwwbWAefVVP61h6Ra46PAVKDZkcd
ZvBdYDE1PHYkjmAeBTRlleHAacWzPw7jCcx06+7uKQnkmHlyuaghjf/h2Oo5R4Qi
nsAsLV4yKpc0qv+jBLlSnAbo4jbKf61sc/SyeldAWWKrq7XM3J2paRFHLIMwLRKE
UVCOmM0B6tbct13EsREgutlNFcju2kBW134i8eIPN3KScO0VZwzhj6DBplliypLG
t/sp0sdSQaO2xWsc04oHN8KWJRJmWJhLBxdgc/h0URCpXYvLuQHXVoNp72yTqczU
I2P5rUJ/rhDhSilqbgfAfuVFC99m+JhsTbzgZs7MBqO7vJoCMtlepeRcoNQOZgio
3nV1I/lYU6sxExLCkhOpiIp/NLDWATpirkztle6SlOijiu7txYgXKwKGCzeeBsdy
vLNgSKK5rLCo10lDNi3I0Hdkhg6Ye73XkeCLDV48qNfZQX5fvIJXp5w9Faf/txmB
RNXRnDy1x7hJVM8Rew62bQgo78bXFji6gJsCK6xAij/WL4PIvsuLVZJXFNitaO2/
6GNYT+Ca8lzLXukbCuavy7Z/RBTxiA0xDxffgDc4w83Irp2FP2PdRnVhjLEkpsn7
oh5JymbOUmm6EIM0lTyT+3HYA6nqgs7cEMXQslLdFQLP3Dcyxb/CmuDWOUM7Sb0C
myrTEtpaNT8dx11jY+99Zq/8HMD8x9KMATh8ZzoFm8ozZKnufWsYvSjEVn9i05au
ZmhIkHTwF2d08fuUmxkeWjiVqrS32evN6azqoCaej7YTFZoKmg4ruqqZL/ZLULYE
2AvNmTrpmNwvwTejrzbb4kDycI8uCh5FndjkKQ5D0Bs0n45gauZzpj2bxUgx3RjP
jtZL0rrJY7ChKEyBLxQ7Kj65592kYb49P80LCSDtkaqrDGGc/BdL1nHmPxX4QUX/
b090AOQdwc5FVBovinE4iFTnWwTDNt3zurxKjb3RlhMlwYRkBPeFrPdI94FcVTkQ
edF+5ImACoL/U9/8pXEPbI1pmYBfDQo3VfLu6hSs5FBLhtFLWn4tgGW+DTEPQxpB
MB+BwmkFOE/jwUVJezPJtXZSHylAsSL8uRBSaqH3+vP4wG3LK+3T9GC2Be0KqfZk
XOiXaUv8GKrZqoWecohEDHH3j6cBD/AupSICUSCOLVVgbsIO50/spJn6J01qhJ96
p+CWkWVkYVm33Ur9vP07M+3D7OjEhXgUMVCTsG+S9XR9O3NOgPcKtDhqMHqnfqLG
HIxZg06i6LYj9qgQhLI+X4kKTALM54waj2g1ju+6tZXUCB6YbFT/G4t0HnMtzNzQ
mICANKBS2fHKWrDPj6N6ss3tVid7xWc35qRVr5LTe9j3Basts/VmDPLp5cvBiFYK
jX/SWftdkky+MCf6fT3z3yPiLIveEGlZN4euktycdiwfn7F9otW9VZ64sVMWtF9C
/AOGV4NmkjY7n4SF4hpgZOykwVXmnimspKZX7j1H4R7TW+XeCO/wXCEts1qJbFeD
iVYSfdvQZTcS+fECtTjXbB2NGCbIzqt6W2n/Ax93naWIorGjpbQGB58cnnRY1nsT
KLD4sCD3QyZXkZM+eAetuPCwN7a4H4KMLsNJpBV1RF/LNmjBiP1PjEARrpdhtz1H
5ZjelCe1YJE2J+ESn210mrpTp7Ud/HqtwY9ikM0vZ9MW6wbIpnFcIk3/+8cWuzVu
W5mvz4BZ9LmLjnn8ZOmCuX9hf3DcWlgHjZDzhOFCe6NhnlTlGICnQtBxycq8nBTv
gg4lhe7GQJ8fp2kR3lBtW3h3claTLGdC44yCs5mR1CpVcOjGBLT+Uxl011XQ6hGz
eVjlsfJCOY7/pU38SZIcEoBgNyKCJ4Y3ptxUDr4EuexaUUqnrbw6AtEBYB8wnviu
JzGbo44WxyYHL3S3jOcexmHrYd0KmOYHBMlBjIDs4pK+WmM0egdS7jn1YqC+cU0q
u59GTfAp/NFtks/fxiIz36nbRR+egl1b0gbWpT4rCT9hyFEyO+ZuXNAUeUuits9q
tCi0saOI1j1Ta9P/MzZ9QqNP5bZi4356504clxMCPOSWE1kvxGjHxc2m3hyqzhXJ
iAUs8LAZ3dqwcvTQH6lXtepahKEigTG4/BdBbcSgbME6hTM4ZIQ36jU3M1salDpy
WSMzn+ZbTkJdREuYNpXlOJSDtX215z3uv0rcX7RdsNxeOfrAtmP1so1tJR8kGQea
o8y7EzvKBufjci+LeZng32DM0RNANkLDGGBIseH/EG5H69H++iTQut703tnopBP0
gcewRy6QWL8gvNxd6u3zQ0I97Z7kiq7+UoiRi9eYN5/HDxd7kT92EcLVObwhhH1+
xXGimpj65tglDBFPGi3Er6ABqZa5mZnR82HxkoTJSy0XMcGU7hRvnrI9SF0JEUPF
Ko8teAPQ8dW3eBAP3JoN3pfeU2kCs1iBI89fA61+e+m1eOHI4KL+QFV2nyFwxLoo
hbSjnoOG22VqnH1cMklBx8xN7ccnAzZpbaSqrJXqNXA26i406q17MvWBdrShDW6r
uOARz1Xk93cBIR6app6TDMgTP/6xCoOEdPNlvtjuLVUWwBY5QCi54N6wQTqD8ydK
1KvrJWwzllwI2N2bUtXetTI6EAmyVh2FW6ETS6XCFxKufBvlSxWeES9zmJyrOqY9
GqcIx/ekBt0uSQ/Q2H+ucRv58S/boT38QEYf2KfpE4nNhDdZxMmTGZAP8zQd4TzB
a6XyEBuTsLGVWfTF+IrgigavlRUOFRlbXJhKUUeJ0BzAqYprxekX0MbYqtvVG5Go
ReMRrZMsea0bMG2EeVbhNY8YDYlUMhwep9qCHYJ9vkLr6wphZGlnajz4f7w1MCjA
RMEhh+gigpiuB+361D03T4bcBUNbWWbfR+r1bXsPOy8hN0lftdi+JuF4x7eoCT5J
vkRGn71txTaGUudRJo0YUhlAWlyRrq9EAotsQsH1aN+ID6qz9MKr9H4wIkXJsKYb
75Zb4a2vu4xLYY2cL1Q2VRY7LNnjziKLyweWX0sL4aGdugaDckoEhivePBVPwLGy
ZNXCacrf47G0y8VmeYfHsmZ+FVtYMw2n+nu1tfLNzz9ZvNldb5A1sqAWfkL//F0z
GGS0mIxz4OA7r64TVizlzMjrAwaqCdq/miV/fXczPj790ZoYcbGhzaXLH43xRsjZ
z8FKudP+0ZHYPa0EVkALBxc7eP21QDiwTF53CtbM91CvMhJr2t1j+shKzQZIT9Gk
5qAXWqD2wDJPMZhGm/Z7d7FbTKida9vwqvLkGMK2+PIvuXhzmHajVwUdWgaIFrfM
/sVhAIl8jSvGiTIq7w1CJy3eelGk25+ac6L0hakkCxmPHU3qDcFEx5KLRGkSC5em
537/FN8nSB9Fzpt8CDPyEM9HQCG6Mh2R+FmYaJviw6fo4hM5PpqQZuaYOUwgDbXT
SF1n/wFFcFBTfcp57xWNG1MMVTPsW96JGK23LXi004EBbrFXTIXqfExKMLn/SzHT
k0sDpMqV6bme4Lho7s0wMqx9rDTGoWag5HG6Y+Jsm5cerHX9m8jDhfH0tAL+227M
5BYvQYW1243bYz2phrlFxyg9Fc5Z58sF5IZ+jupViaQ3x6/k7n0ME0iXHfK4aci0
Zb9Ftf93xw0hvrhGQZIsFnqRJatNUVvzA/Qeyfl+uliXbYrCOQL78qkO1HPG+0Py
vTJT1ptcg8aA+p/ILgv4fxt1/8vXTIMaCNNqypctaZGT3l+8WeKGv7muJZ4nrdcr
hjdVQiPhos4eAjHbwQT5N5IRSW73GoP/AEGxKYPBJLppWV2QhSrbxcWOYebb+biA
Q4pkyveaA2ZtzbQZ/sxyhQEUDFb8N+GuwnT8dqxXqmnqeHiDG7OrnI68/PeuRehO
ePozqBTh8I+YdlnrdXrFu99XA1sD6+0AYQ9PGsyKY+0=
`pragma protect end_protected      
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
cduISWl/kHL+TlxDja6AXe5Wb7PicPaWryegAaSx7zQX8SunxQL/gMcA2HDkdUuk
N70oQZjX3dbmrsFkjR2E84fHDUjaic/KJS+EXM43cWRF5RTbvB1JVGRQeusgXoej
z0MB1JDBTxHvKfku/EeXOL9lqie4/i5mJzcvd7UV5Tc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 135439    )
KRZ6duTuXSxHIaAxEOE6avafBs55JZrrO12iwT7Tn6gvRh0f2KA0wA3VRhWchD0D
Z5pnDg1bjODmlvw2x4w5JSYzcJWGqW9OAlryuuo1bmuXBsbF6Cv7B4R5mchRJa1a
qKD9lFiF7ZjRTIGqI8eXs13OsuWpHF6LYq75c9VMhjbor8DSTjXBQ51aAGeg9NWG
ZUBYhuPTGVt3wzvHglzzBLqUiz9BjaalPzKR4JQJ5u8bVd/QmdwL+O5Gx+zeqK4j
FgW9G4pkXBuxCakhYsEmu9m2JPzhN33lsinB5kS1W+ed5xqCw5ADd9cGn269JLZT
2+161InkL7KB32dh4IYrptoDH410LOY0IbTzv/3PJetnDBATnUEwJGYVhD75hfn4
hE5IYHLMUa3D9oau4vDoLpTCX6M4oWttGEyGbSs+b4fWBtWdWAWVXBGm/HKBrTYi
N1metk1C2GaNFNwwOui2CjwhhlflXqt1Zhz0RdPCFoGZ00o+9x0S5+Fhk4TmcIT/
GwpZu3zSMvvf/CYs1hDwsLcnxlf7Gfjg/9r2xt3kQ0MYWlVolcSXRyedcLejVmKs
vTyZPXzOMQLTKCpBsKTXL8tIiD3RaLtMmFtdujkLTMnsLlhF+eUbzx1zRSeQzBoL
SRTJBMyfvX3lzE/UTEn8weZBPSnSLBdGo7JakMCGAIaN7JFbSx5UOFYdT+KAbNDd
mFbSsd8EgiWc0FS6iz4HCztPx+HUzuNT8ly2WB9aYXllBc8WiGPVryKKu+YRIJoZ
5xSk9CMoWoNNSJ4HrFbqGQ==
`pragma protect end_protected
//vcs_vip_protect      
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
IoUIzR6658JQYyQ1GDbFFTGdolRfNUAOprqaMBNEQdss4hcrCYETq8oMvJjByCLA
+ahsX8FALKpt36SZm2gAMhcxnURnZaMmCA+O1vG+ULaBJQMC7HdnyozCu+YxqPGk
40lKkvzchcLrALtwhCDzfuMvv+Dkys9HTpSzkQ4qIQg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 162525    )
vioGS5rVtKMRnuWNd1tm27DMKF93hgyEeXV1Lhv4lUTxN/cFQ/HfHD3G3yMzZ5UU
yV5DigAvGEGVPDKV0RDRRo1WgbG3184HqrRLC63dVLHwvQ+LDumgg7W0/FXpbShg
LtX8CqyXJ7bKNebW68IicMy6U/X2LuQI/ojNyCJRlSaf7ZzOdHPMEJVMnC6unH1o
9NVkzC9hW0xo1v7O+rhkyiJIUuyTWcJAOnTE0frQULxrizpJgdjjBv65KcScxm92
ETqncr07kaa/d7D+PqSVwYzbq0kpY/4mKsMQ7Bevh2dNo8lfVt9rPrfod8wHhxy1
oqJB7t/1bmj+1uj/MQImXTSCbFhIvOSXaSa4t9YjspLpBbfhay7c7oPjQsG6w00o
ZAZTYCzAl7eoH9SHQxXeiyTHXU/nE0dj6N4j9o+ETs2dliFanLEvN8eX8dyKOOA9
iSCbxIsFQ5YS6/s2gNKxXjCl+09VzgnVZJ6d/FtpU1zPzSAqYFJg6BkMa6EGweqJ
7BwhWU/K6gX9EFZLpcDa98Q6O2mdRcaB/5GdF2/Dt9s76SFXL36h0uOgcCrVcXqW
kRpesTl6GgJwdHgfO+gXPwDimRj6zYBY9s94dBkMu+/9s5OYWdkb0X81TvhxvmXy
dshLagyX8c9gg4njV+ckVALt/9kXd/LdXmSdw1+cyy5el+t52JrWkqjAXbmkzNwz
pzVWX5iFXA863s4wPisi2HIIiISXiMK0szPPq3wiiSscDCPgc6D+UCq6aRgT4ROI
SSEIX9Kf73Pumb6TE5dS8NkmyWrumuoI4ljvaVo9+YPBshqCrW6DxZ2iTOkl0ISf
d6FWlxQreojLxnQvBmB6+dp4Um0Zy9tb/WkPNTSreQt1N5jic3ERkvMY9rSeySPZ
yW6iN1Kq7VvQu+y5kkwEBKbNrjjyNj1psrFVBdMwB6nftpODARWts+HBfxnUCo1P
I3d2Jqo/o1YhGrpqTlyx67UWIVlV6UD62tAf36qQihibZFGboORA0SoExLJRs8nK
+YWD/dd8BWh1GzBa4q10pvsrX4HdrPB+0lAbF1c5xCXpDhcDxspgOlgUjCtt8Q13
Ij1h4Fvs3OFAvLgFXVV2XjTdIcr4hFRMld1UHhmNcqjvYfHeFw4r9mIs8IzpomSB
AgHSkQLpIqgZTO6+PCx+Zvz1CouZCrf8oJp43OX3sCpqdI0HP9lzEinno8GvZheL
Uu3QAuHsfxU0HwUn4G9mf5UUhyKfEc1XfbZOndwLotZ6/LMFX9mz5DZBPMYVz+Sg
0qpjNMsRCvI0lb9zJwyJ0mSTsiKMN9ujwEEiRxpe2V3eqj4jdugPrWTmB7SaPBR4
4ZI80idGljpPqM6cYjLdmV6cgyppAOf2dmS2jQiHjrdzEvcx7pvAXKW7CCDny+l2
1/OpbNm4ZQDVmbm0Fd+DjU6m8VnrI+lxcwoTY7YHhf1EXCWtNZleSqwr9tLiCQ1E
e0Bds0RgJki7AuvQAONAJQCPfdNKEs5Br1tu1hLifN1778fzJLCUnnvIDl9p6PCN
WemHf2wMJ+LaM9JKHUhNm741K/f4qC6RpCU9qmImR3Wv4F24fN442QZWUZuzBbPd
FdbiLGtS8p6GDZfXFCKv2h2rgU0dZbeZ5gWAwlhkF/78NrlJNq1CDLqL/xxD33rA
pwA9JYDAJIk1Bxs+vRhYmdeMX0uWP7VXvxdwENK10xvCri7mx9lHIrUr7w/m88AW
MMd9o9htTHe2LcCGZNBS34FlZj6Hn2ECEIqW9BNno5sZ/muGGYYQlavx6qKU02iy
0Uk1etT0XUTmxBcnZllg9qrp7SDFc9LDXYMPrRp3oFMP4l1twpGeF2BY3wTiwcEp
YmWf5Iv35uWkZ7CwmxtVHaLozRz7LKnXFdpiurDzWWLRkjTsilmqMWdSYghd8RId
xNxORCiv3unaSA7x3cMHHnabQT8F8LTnhseU4CY648LbUZ45qElS16cK/sYvIa3C
N+kTITDgBsqaDuxJID0TNVwHrH3Zd1CGnxymdyR8n75bOBHR/mqdV7IyfZqNZnwG
WUPry7d7rPzbUFecBiyayw8txrNHUiJFV96fe9H64OPBgkF+VHbH4M/xNCWwE40S
8QFHOr7vnCzZAT04rJTzVSc2CAVm/KWrJpMzgYyQe72L9ixWVRcMKU47g8Q2n8BM
P6cb/O00WiD+vs2YL4SWGeyYFutJqW1k5Zd8+NKoBpi6Q7ppX4NqZM3p3Inj8Ldh
FYSNS8btKGcJGj6u5+L2JzMdRI7LmE927eJ0vUPv6+pvtZnBSI8OUm/luhV7OcNh
tHYqG2EIsz+eJPgTIkza9Ap4IappX9WitY2mGbZZvNkbaIeY6szZEjk4K/DcKdEy
hj6njW/2aRl0VGBMZHInUAlTrm+HJV2fl9mmJXX89+uHwfJ50RSdXBPo9ROX/vev
e8Z22Ba3RAwILGUDwTCy+XIz4lT3zMnIQfOvPoTKZ+BdySvvnqtqmVZmzmEtMmqN
/j1galcNIuO6Vp+y+oxn53vng38qPsF8xPR/oJ6Ebv0NRpZzyGtQQYSElzyn9vB5
6NpT/4DDjgcI26PmfSERDKxkS5yFKLqRoIkIvs9TR0Emhd1bUxzMaN5+IJOXzQ7i
7LvDPsfWqaVuRIIOsyt9wttApwnXL+K5lDGY7nA6SuECWOQPEvyFlS3z8QGG10Ns
3W1io+6x7Jm9JSsKfaDXPvgu6fwv8fxoUxjCKsqBa+5mP90wwSfeTZVtlFq2Fimb
UNpxMl0umANO91sfNejyUcGHh3klUUgrjf+7tTSqlZ16Tsgk5dPbbrE+NnGyES1m
cZB7R3LBfHvsIoMyQRcVUoS+QutcWeW/H9byOTlX1GnllF6bcsF1jvcRKoMCUnJ6
wFbxpHPzy1dYShR32v21+wxD6SEIeeUcPouZuYIUe95g39fx8mWp1nP8k472cDtp
cR+orpW07O2iO0SXakN3tw7zkmlgldv6YkivR+OlKwUj72y8V1gjxtsgDRNwU0QZ
yn+kl6J9PVQx41u6+yyUWY7Vtl9aazxYszHg1FXGWzorf7dh0qDAMYeYqdWpDDTe
7MkAMFXLxuwpeRrCm68CGK8z2DLP9UfXs7uJFp6WmhUCrwA66Vj01LshmHomnbWZ
Kwot5C4gpPQu6vFzvM2AwNGjAhJwvaAxKRQX2ENxGVrVMO72NEBjf+iWVSDDmFUk
tnOQWmABkGdnCGBrnZIT8tizk/GGq8rECr3DYUwIXJnwwNv1XrCTqShGtfgjDfT2
CH3w4FCfKjeEudGxebBKTcRBIQ/MPpbEAeGDEjN9zV5NuaKzr/OOHIYExJ2F6rG7
94uzmowDMfSfLn+2weokHVKLpeq2HFQtVMhwYRT6zue4LTMuQg5jWnephR/isTCx
FQmItCG8oraflcKXvtvElK44Dn0hym8WAEDQjXccUc6ohUdeGXcTpAC8uBvfG4zA
HhgojnnX9lIdqg+2I4K1OTSjtk86fnDw38eFjlELxXXuL6RSd3TReypxnRtuJb1Z
wh2h+P48JP8LQfDRlumkfhAmB/yanYOQNcaEXD3otGNmldSRgJc8aGFgni+G1GmW
2FX7+fdiPUJzV24gTPHCgBKmFz+H1t6FtWRiLYyLfbcjTFnIki1JPrqWNHNbvVx8
PpoxHvpcmql5m8weryrfbDWYedWxH0q99Wbu59hN6oVmMZ27LDWH4ZjUl+Dj69Pg
UlR/TJ9pqdD6/MUiL6XoVLdEXky33KlwlBLaiyaGs2AWSu171oXuEUmP7dhdjdd4
KM5mANH6S+ZHdd2sW8iE+qwRZ+bxw3DRhHKSrlgaGnYqun/YjbqbCA+bzcs5ysDJ
SvTJImyO6oSBOgLGMFOSQdsFNX3h6Ip2BoGoBDa38cOSY4wp9Y9thswfMKR5IQvR
1Ku5D+nyjWEh7y4wkplQNJEquT86kOudmQk72TDpV3+H45aZ+YSgppFh4ZGUSO+M
O4+KKdRlkw6Aq8yAA9oMSP3o982iCIuOXodDKj/dLTk4vUfitKv2dI8PAptexA43
Db0OqKTo9xvnIkwk+e3aTBpRak+nnu7zjlPbyop2fxXdAEUBNsE3Ojixi/gQ9Wmu
Rn6agqIR7Uexc7yl6lrf0kauaFIHmTu8XnBYwfR8DKbqOWQXJPl0715GsGmjhRlH
L5AsjLEzsjROggGqDB/EFw00KavsyMDKKVLSk8o136u4xXg/NYk7KmU6To6L9eyr
P6GnJ5b877cHQoBe4C3qHRe3fSaZ/596sqIz0V7azXNnuA6uvaSvjKGb3XvAWED6
CCbWqTtSSBk6Bgf3WKBssZs3L6qbY3NmCXoYiZnG7t09tCMx/pqfFUX2c5y5Ph4/
4ij0WTMp4gGI5q/iAJN9M7XqEDRUWgAjwb96zuq6W9ayuvsMamrXEzIk/PqHYVXW
hLP7RAcjbWxRLfWjrdwvZEeESVEFWRbclYcLLJ/5wH43HEYESJtXWPjnTi9Qmqof
Sjb+/JvOL1yUCOr5EKSKrdh2REQ8GN7sqPWUHspCanDZT/4GDZ5uC2hiucvOoT38
pflz56jRTn1DHP+LzgEKLDH2jnDdhuuXYa804uuYQrCrGS0HPSDUXoTYaKITNPCw
qAjYhkfGq9f/qOvQUdZMjQB2KEsnVdjtrLiWfeYYcDVt5Z/fguVNnXwmQIPyqEXf
uKxn1xJ/8OZJiaUOpuM2TZQuMgT7ETbJrko8WKKhEcGn2yXy3wXbiFEwqhYbvCKc
81jb21lnUx3b3RJqipLNRyZh1VjNf0A875XJj0FoVNY7v00wIFljLiWCKC/dgjx/
bmWX6FodMiniezEpK+CgJxVbf4i92BHOEYCNMyonmSY1qde6u4LeHMKfO357Driw
w5S3/EwxRGlUdWSmsYJp9dbiS+xC2RIkxaAu8UPjMazGCVfkXpjK5JoXREIVQTmS
irV7Bd17EoPv07T6JwvqqcYVeTHDiSiUXhVitmko7PlVEdOq4V+Zc2cTCcQDd5s5
VblFReBjVeuU7nwE0yvaZHeP6TRqxBi0wBv5UDuFBIn2b5ez2Jdf3THmsTvaU/KF
GkJ1+a88Cp/HRg9N3ZQYUuwO5MIVJb0flyMLxte6R9xD0TMXqRrZB5onk8RNRmTr
P6rY+9PgxoMQm9o6HuPqLMjQJhFE54Ft3irF7wwhwu+sYx+MH9cw7cPmAhjoU+lp
7rkM1ELWLwT9mbZ4bD4KbMcN/985NVyh2APQ/UHBLjEjWqcbcdb8aeuR6FA+Xcfp
8bgeKO2uZFzfiA/+4vvWGtvX7Bsg8RoEBvaaxCZ9p/XgPyfxSdoJf8j8JYHZmFp8
yd3QXODt0mgixtvkVWgIvceNqfXH556wSAW3xsnaL9MXRRNXkBykTqXtb7oC67U/
r9jKxa3wT33HmWtCnmW8oOuFi6lna4i7tcigVLc26MxjtH2NGAWMkW+YyiWwM4Uy
PZ9CbLEvukNAgckGabzSPJzpClCAjmiAGU2EZOoD/sKu/JJvX4QqkCIwJageoh3d
r+PdNNSOYKx65fxWiX13pWR8PIn+zsFd3bCaqahq64uFrHpw/qL1q0L4VUi/Mq+X
vU49JKoKQMJU7hrGWli4QxYDgmQjUQNIVO5qLSFJSMsUnHKM5NbVHo29E3s92v+0
PXKmb0nglAwmTX/9N/BbLCWsNpTY0KAWDekSe+iB59DbQgzBiKbwoNTyLOsPFA1R
hdkeE068BE7h5SrIlYe7YlY+kCYTfS6SwCO9l7IbWXN5efx8dPe+xcp0m+CYwRz4
uF4m9q0OEI42D//q6DO3K6a7Nk2iXF/O6m9SgN4XUzGDzfxQhrdjPm0GHZOFozRd
vxUBJ24Q3fd5yMJC6F/qb/nIdoADC9Hlt5Lpu1XYDhCPQs9DUqn0dOiAd7moaJuJ
BaSw63jqRnZIHfWO+cg3X5+8EaYI5I2/t0Hrc4lY5t3+b4qLiG+SRDvw4enXYuX3
KmkxCky64+Y5V0RU8KnnJZsSG4hKDHkje1Y8oMS7Yg/uhEQUiVeZNU9yghique0Z
nXFsdbkSFjVp03IhZYgKyH9uURJHtVG7+E1UhtGSSnnZqHd2+DJPQGV3yfwoTzAX
NngfIKzjZSZaLFdLRCp75es+GudkfHqCnCavcvI6gU4CVokHg24+yLfJnnyigPTd
6SuDuKRcra6vCs5IiXikK2zFYvx3c7pEsX9aIFq3ZapkKqMct351R14D3j5coqxb
RDrWBgkDo0ZMS6laSbtR+EUNDxJXmSmKUFx/u3TfIbmnXpMOfMtTrG+WY80G+dTJ
mAIgQFTgaxHpIGlLamebdBAzN2DZEWHXS6CI6bhmehNBewc9DoNTNgMeKeNBfXIN
1xcHvMeSLkVshq9vYumZ4rWlcVMvzWD3fTheVkz1fbof9USR+FfRovIWM5qkmZDT
xQBUd4vR8sVA0IPer7/v7mta3bKSrVx+NPsK6gY+jGEB+DzqWrno7E/H41zZ2lCN
Ce922ztMv3b5TEDX4PsQhBX1ciQla9DLRtzJKH4QtEE9kyHyewKK7mG4lYI6SD0I
Du8DIF7JKg7pmSRZOE2fy7StfIZ+Io1PFdGQtQXUESO9+unJ77Yv1OETAWP6odAN
4Va46PT9C4znLsw+xGF2jPgiyB0o3+l7gYadpIyWv0awkpDy4yiuKNtLQfWvgAA4
TZy4lulUEVC7GHcBNFfyzg/J5uwJN74e+2Z+xxk041No7gzedvk+iLYoKZACJ0+G
wY1C7wrkQ7dZrhlb84EVq3qLGIB/offPV3hKJiGlJhewaAkCvq6ba22xLVuV/x5n
g+AW+GLt1ur/5Jf2P0pjDvmK6jJKlByonMFEzufu0fHBYLdk5xwYe+BtZcFlDseU
ytrdwQYJ2PlSvSCxa03gL7wtIJOwHvKjUud2WwjRCWhoSa1fy9fvNUxRrLffrARg
V/fHvudV4H59LN7LJR0x9qpUfAf5pWmhhozVlNrOsXVTWHe3Y+Ye+Pamd8edi8V1
DnvO82dETuvLvSnq7xn0qlDzhnnhkF+wRxZ0arSmaj+gFVLAZd/s3gkx3qpinLkZ
vP1oSI/bXoIMPO52Hj96BC9Jg7AuLF8CFZ/tU6HS/t0a3+86PiNa/hRs6V9XXTov
rd66huHNYPb0yIQ/1wRwpefVlClhh0IO1l/tZ9ZGYH0dVYmL89RNYUT1g7q2R9U2
QZH1yk6QTDyHJi3ZmGoQfHEJsZBVqQNT8BE5KFHQI7LvIZWtEjqVNQsR2XSh1EJY
XWeM5rKofzyEf0CPHtWDxMOoB/bWNVw7RsQyzOQSFTKGxuaRi5hvOu5kT+X8MwDP
wl2ithEsBMd3IFvtjRc1M1F0sG9Zb4+2Lldga4kyypoZ8pltQCLCqWzxsRs9NICP
9Hvbkykqy2W874Eg0sPUHRLlQ18+J9csaETl1LPJxQBcqcHwXf989MxTTcj893Mg
Dl5kklIP//EKwiMBo/KcsnO4cI7TVzehQq8USzDkVXu1+3iJf7lXLo5C7vtdi6jl
lGOhzTyqcPiFu8Hn158PAhb++syx9uIjg0jRjWoCq5OHwf/2Ep9P+WmwsXMxJEaI
3bbw7itj4jawjpUIufDUuQdQENLznHrq3CPXo4sAgpS0kelbVNBQ2/6UWMo549mO
9Ts+KoneXan5Cjy7rg5CeF6lgFHwtklqy4v4Y8uAPI14PuMZ2dNzX4fXJErL/LWU
0Mvz2lstR9Hw8XrWRnlEVe/a5tMSe+bHxSuJ2wO4dXyeFIo9NAA+x31NPYOc8yam
zF00Awxq0XxyRs5RQKWq5kj9hjX7keiM1Q9EEKP6aFEsaKe60f/I2zJYqCZZVWFQ
zxUZmfah6coobQ7r7pJZQ8thcPNbYhQVcGzMKlwpYViCB1pPqYVYCwheWNLEcecf
OgM0KVqapLCcr/ZyEZ/dpnAVeuSMeArYPJjloHXDh7bTKTW1mx1UW85ttZ8xYuWE
kO2AcvEC18aXD+iheeIVCP2T/G7mzec3ipGz7vpR/JVmmlqTfzU85JPHPQ+1a2Jb
6PvHlSHd8iO/6xrvzzZA+vh8y1I0n65hnNUTbBJH5BBZJAs7rw5dGTgGBeZcnqVQ
OztqUWlWRHPwV6Et8YNrteiMQjAQq2vm9xtB3NvjPp0P6LDqdIApdxCWr59S1jIV
ogwFmACJR2KDYo7EL0XBjLoewWAoKcxdBY1fk51nd9HJZMM7BCTYOCM8he/zqYHp
efrl12VahHHRue1Z0BaCDGW0vXPzqskNGzVZBCETMlZNKSLkhcncfCGpl+K4QVVd
KNC0DRqbidljVjvSYTs6QrGHODvmgDn14+7PFMDMCodUZoySibnFp16HmLGiL3x1
T4+mG6CHb9xEKgLaFWqSr2qrfBVURRAgILUSZwzaCdcpLyvB+KwZtFV7QttUWpxO
j/axzRKxybOZwoMr1crvJgDo/ErmGc8FruVhcX4Y/Zjpsvq7Vb3ebzTmA9PPc3DV
u3fBb0vwspMEEYfJwpMVmQ1+rdoz7g9oVn2J5gy/R3M0gEeuGHK7VHlGZZT0ti7q
p5ADccGuWrPI3oKZrd9P8P2t3VTrqkzz/qQyGimpinhQaL2u2EzWieynkPUpUGEr
h+yXsPGN2q/+Tnzjme1M5dkK8KnmetcQCU3uizZlkzelPd9ZH+5z7UoSbAc/kR9h
XW7MgIw00fEepBpmZiKKvkFfGnuDDFjcwoggxsu2qyjbFP1guA03BwhpcCFQAqQH
BTGsCIsqyUBkxZZ4lK+gPSWXkkT/R0sXobtV199iRUToVKEjcPmv7P34wgqHsyHW
6AoWNC3lqk5KKW5eJQgm1mrGEwRufbkJ8hUK1KzY4DJ30xOVw1Zor/+7L04ePF8T
JVhqLMjlXVAn6gdxn3tGRLGEpycfC5BnhN9NMimfTM4Y9Un8Z0T5aaVglsno04UI
C2goS5ZeqswUc5dazvGe1Wg4IiPkd/r1I/2MarkEZoa2f63agDi4Ij6VCrVcw5qf
/FwJkYdEPMvuHFYMQED3WIYfo/GzZEJddYyMkYbmRbNqt71gHxnEgzowgoM3g6Uq
8JBg99SjDmF6tjQumG3UR+BHUpUCDQn+G835c0H+NORlXkz3SrFq4sdCbg0fec0L
JcweYrMgveQ5sTM9l8pXW/VPSycWbsgUD++ONx5xzhZQ7Co4ZYh2aNfl5pgJfxmQ
GubGyFrfszLEq66NpIG+ipu1xqBOPb8C/xmxLAHlQhHiWM0fQfUQIyjO7gkviGxD
wjr7ywjlxm2JhrzcaPhavF46ZBn8YsMDCy7CXNgc/S4wc4r5P64BRcX97jQWF7CF
n+tNOdFy+F+UoBUkFknxNm0kbdSDTGaCctlxwhA4IpH521xTDzXC4NcCtrEvTfq+
VfYrsQmtaW+StfhrdLAwK2Sg2W/xViqEC1DMTudvLfIxJ6ZjszpLhU5bihgZf3QH
Njk1wIIjmD1FoW1T8JgTaoKcol6ibDR5Bc4AzbD+a4kL3uFpISlKRVQyyBstcMXM
k/T55DGYbec98toh91ZsEsCTO5gMG6OJ8k9QP1mXywvI+GrK7SJ00Opw8ocmOO+c
gAR5RNb2QK8OPwuDaJ721Oou5Owjq5kHnK/d588vwJlZkeZUbmYNASCdiVwmlkEd
bzkd5Q2gK0uqG1ZBJjiPdwRlGuUxNcQo5/CkLvfem3jwcVc7BhcZv1BcX3qLyhDh
5Mv/ebsjwF7MawVh7ryzh5BoIDjosPWT09M+c2rjKhLynEe8QKNl2hTmES6TcZ5b
eOpbbK0CQPB7lax007Iw1XR5W9E75Ly/5DCDCliPjhbJh8Vvqe4rmRckxwjhXKMn
nUf8EL1wVUPLX4q0f7xoDrl1RHlDBj5ZKtqwOgR7RQyskrJrX7zVl0kQuPlitAve
B36AfckR01GSAE+4QaIA6FlBthxvYbXquiRCtgrXL9aBMK9KGCxxfRgVl+ZRrBfb
GtK+TawDVebRnh2esxnIsJFApfOdoa6Br9VV+nKMeRVIV7h4DPN6gE2zXM4kSfaz
Y3ivfPJuhRktr2LHPTzs/yF7MzpJkI2gKdhHHOzlh14gvEyZugXZXzBv25fZaYsS
+eEDUCkyAVZl2vVBpk1AoPhFC91tQDmPwG9yK8G+vFegBLEtD1LCFezfnRHgMgTr
a9ygD46AlrWZC4miy0wXxydQrCXa05LXcpn33j0myzLY5xsyOf+/a80EjvEYikhS
jvD/X+MqLGufh7otbnFZ2Z+loia3svOvPKGVhSQqXOyeuBjEAvzYwj+3f09BQdOB
nFBw9t3W6mMzILqTH+JKjq/jzn2drZnZdCD6GTsjbyOqL5Sa0Xp8DWByBMurDUGd
z3oCm+foyFg/5lY4ABIjDY9ByLsivA6rEZE9jSY8SpnqHNE4mzjeNIjt5HB0tdqw
p4NUKZylYnHxIYYXjJn9IvDtFqYBk8C6sS/dlS5ynqA4PzL8RKRye7SxsV8X8vly
kC8r6IZqenthIwtxMq+TwWNPVIW1+8QFn916m4xhIrJbWwW6akTYG/ltbc0cOXQk
fSwnxmDF2CtRijQqAYnEN3jU9/zkU4BRRueYT6d47/X/47GCznxNQohNvBlw8bAE
qhbzgykQK52CaJq9AA7jG84dzcC//Rt3ozTV/G3JQgRkvWIKQI64dlYI+K8dDqqF
cKstIN778pqa6SRIMoTk5TZI+pdmatp5MPWHJjEB0xehcuduaRMwI3Lmu8YZj2Qw
BqfxCrx310xsIm1YL/CYbYSl1K8iu8KGSVoyyglfA1iX4ryX4fD4MwKjM5MCmpsj
d//6s44EJBYbpvkzNWHNY1e/0ba3aM02V0zQ0fyXwUWOMB5OKJDp1beB7srYXvWi
Btu3uwTA1C+ng4xyZCkSVF4n0Adqwf5eAH9jnlZe1X3CKlmuSLfoa99iAl+HHsEy
a+TaskAVOIToVUoubTiqXAy3aKkHi8o5M4+M7LJuM/kBNW3Eh5rdWvV6ecHAc2E6
oDybzcGKmSd3RbkVhpXi6uU6JCvVedAhfJcb0NTKFGMGFt3VUxHGvAaijUaOQftC
iPBaBmUD6yuD6+dAIowe67K9nonS8RRaxxIT4aLKUp7H63441Oxw4+R36ryKJPH7
+o/m/I5PzTsp/O07i3WPYtYo5BwsxlCe1gnWCi2uddTAUyiLemNexqTbPZPS8AMg
5ouAwE53+5oNS1lD5P5b4JJXAv/R+ybJ+M3Nhr36ZNpkRmA4y7gbGbzcEtUyK48Y
cxM9J9NVKLFWy85QM4kV4TFvV3g7PCXg3yE/2DErAdSxcGD4Cx4FvppQFRGbYWiK
sl5qdwqQLS3f+G1Ldzj7ClFFMVzO7jq3iF6c6T/uf7ZnWZH/L1NkN4iTYByVDjyR
AB7PbzmopJNtMlfDzYRKJr5CC6m09zPP2hX1xWlg0AoDXUVE0SYGPfUDpKALQpPB
CGnD7Pkc0l7OZ9qKqmLaoNYd6Ukc2rczpp9DdkbWwCB7+1OA9n6V/rb60Gfjg5Sb
RQ0FgTTMNv7h8ZxmP3JDKv+rvRKG4UrD27BLGhBpzHLv3kXw7ykGk3JNwuoIw45X
k16mlp2MnzUwhqubeMd5QyuFbckcJPtTvjl43uGBdXD271p38duVJt69iusKyZ24
xDrFB89z2DIBsSlPsorDtHfC530JTUEmPW9Jo9UR+OCaxPDfLMf+fzi/JgPX2OkG
rtXWtzye1a3nU1AVJ8m5olnYdk6EnVYpz/V6Dhzd165kqe3I4sYxEGu+uu8BDR0M
urRo+0p75yrx0f6iZREbk7ThshkqR2b7ozRKVXrDmURLIKb3WjxBfbTzs+vsSR+f
oD+sFS0jllCcZsP//q74Y0q8SeU/m2n3cNekvkRmlztyTaUaE1byYFVvn1KsV/KX
m4HfxLd7O4gD6LMBM8Iif1AssG63aV/7evPVA0JJLW68nkRNmbUAeurvKbECXRgx
no4tiwIzfbe6TLLURXvjogXl0OJdrtfolmnIWSaFBTF+hORNbFsZ67cYWzyz9299
08LUpqWhIR6gpfnz4HvsJ6IBWAi80GjHR4/yN9EISMN9gAPvsaAEFzkwKyEI0ehR
pBY4bMOR3ZG2XnZzLhI8UytRXYkq2Wt57Y54K/LdhnJAToRapb/zjWm0fmVjsMff
wQh3AA4NbEw/yiU6ByJZr/Cw6atEU1u4l57D54PZa17Tc7ZfiWzxdD8sncdRE+P1
6ZHEbk8+zTYb9mh4PyDeu/4+n5ocigb3HL3mIDGUUXO7pH7OtqGybL4vdHjrPOFQ
3wxIwrbw8AqOb1wLWI7xnaaJP0vuM89Kf+MLZFH4yRS00g/EqUoLHWjXbS6C7prh
/ZNuus1vF/OEqFkGwoLIXjjXCNKW1b5Ee1x12LpGSSA7NU+Bh0mHWiyIQZCpc6+u
0lV8MMcHxTqAa+jrWNzfAbbECcq9b/hxvS5ArxpJK0OJ19V4Yi9LUfKKl1S/Rthf
Auwx326QMY75cAcaPhkAJXtvWcriNMpp/E9MAzk0wzsbM6lcju2GdJv1Vn/DCG6D
cLbzUEN4czS22qhPW5ICn9s9T4trI47E5faoB0mrfRfyN6EMxqaISp4BX5jDOdog
+dtEDADn5kLE/kmaDSG4tqhPPvroXJpdpe0EsxD5F+gUS6pJUDKofI/Oy9a0vsRM
sZqUYA5Bz+ZoD8prk1JxQQMlZ66lF+WXkkEG5KD6nh7ZqYtcXlur3qsP4y2YPOh+
NUu/puCCsa2wE/jz2qv6xZ/EqRVrKH6OBpvW8CB4/7texNMXK5RSu5FK8kCzmRVD
SnA0T14m8mNe5I9RIL1WuGOP3Ow08bw9MP90uHP5X85BvyYfgvYSh0p/NWbxon7d
jDYDKoeKjJlhklXKSAPKmmRyhzUPluqNpi6aKnnjdyOUlBVZ9v4jQSlOFwpuCjs+
rq/a2r1guBc2805MQVMU9mH5wNTyOrHWpSxdQ3gUgVa8ayqKiNIN1vnh9Yhsi+fg
pkTLdG91Ggz227WMgVwLjYroBS7q6+bQjfWZtHC+XlRdNLCW9q83d+miqJB+Gbz5
DdL4UVQo4v6Xhot/GxL4oNnvu2yIrlXgHxaAv90edVVIl39Jp3gk5K+RbDLDT60e
fsiL9vc2ZrKrb/orveWy8n0GJObxarljE9ZV0ap+/51jbFUS/+bf+FJN/vqVxgmd
X99tjisa83FPDIHZ5rmC9ZCXQeYJRDh75JuDINKpr19VKJM5V002NdWN5r2tDWbK
4jLjJIp/uY9vq/4Q+Wj1IzBZmHDC75tSoG3mtvWV0N8umZzlLvDgcfNO0/BwXR8Z
zc6tegmyO1NEa8fbr4aICMlIVQeNX/L5xPHMx481V/FMRBqf4OxbbbTyEwIdq3Z/
1+rPOxn/iehjOvbs+6R9rUz2IQX8gCV/gE7SrbWhnt6vAUE+FfOsUsZ2Q3nrSjqB
2t2mmhUi5WnOplQ9UnLSEXucR4C5kkKldq2hzWUBdkrOuez45bpGEkkItyEkfhCD
MK7/RgaSgyTco7CFP7QT39rrSTCaUlYE6ajhRS6jSUYag3s5LGXSI5tKcg5VqeW2
3nxp15orpcEqkI4yZwP9GxI8aND/0FVo76JC99HvIKr+iuR3pxGMr/eE2AIPjSMd
wqgzvBLYXKzaTDqj4cdpnUdO1Q2Gl4k9AXaoZGnrjDqLwKFidXX6+Djl/h1YtdZF
O3Go8hrzK3rR+lJFOxSfhkEWiLWHJyaeCgMXn6e7imBywIDidBMox3QP4vUvJ3nY
lcoceBEQvtrkCUY8qUPNkTNFC0qvLs5Ky+ZnMb2abAt1N+dPOiltqvaCbeT3nI9d
h1j0Zc3wUmii7H98Qpsm1niPuqFH25o/LdT9w+Hu95K/HEygCXOI4kKGkJebcjs6
gpTMyYJ0TPt236/wi7yPbdlvz3qMfrrkn7dP2H3/OV70QmahYUlcpxBXKyH+MYWB
WkEI5Dl8n8Ng2tt1A9Bnee6CmsR1c6TEmlWhLxcKifQIHfqzaEkgQ5ddvuRhR7BP
YewJ5TT/8/u1dRZuYPZcxhHLN7w2bSaXxQU5aGh7Y96mSoym5BzNhq9zV9EwbBRm
d/plkTAyhCVVT/vfB8RnquJLq9LxDXDs/RqY6DzbFrx4cYzbbiFFghj/J25EF4RT
1itIavGQlmhMAPhpEhDaAA8TntgjQEadmklsDwuB+fAB2+4kYRT6MBQl3wtX0LUJ
nyUYcdVsidOmbGKG3DV6V7kd+Cg1IpJGA9zjedyZvWfUlbSS+iUBq12m0T+jvSxT
HhqpRVfLhdQM2ZkAq84uX2Al9I/laCrPwo7DcF/k1aj5DtLzFxVZMTtCGZW2LEr0
1gscJ3MW6JXApomFI4+y/sOGADDeAhUWLlqVMSVBC9atABrwb4XYmVUKqHWwugXz
Z7SN2yWO6vRXNEQF/xCSWjgE2vpI7kvQbGbGR0suMj5ZgLWE7M+QOcKDsBOTW668
MMhmIVVEH5XVUPIPTwLvqwl3vkTSe+ETLwvUsOgznGCukh8J4/S2Sp7UN/iLlUOn
O8ZJ9uDyJxVunleosfuJSPqyiOekzlynB8emMNpBjhFqK8Cv5Klc7J0u/CorXEr8
UIwby8NFy+hMr1rgKwqW1gaorZJ07EZmQWR20O0dkkDisX1xofQHUeXL8N7Bixd7
HWzj0PC12Tw4inYZjtd4wUIURB/gAzHTJnkyG5nvM/EXOhmuOdiXHTP8ePCc0Y3W
ArePsaD8KIi+G6eQOwvcrypwgN+YVpztw+SrIOdYw3zzbJ96HdIP48C8MXb3hdEB
oItUm+iFXRcMeuAwiMlyL1aF0MlBMFamz+NtrPOAAO29W0Ukz8LkaWPHhk/QrJak
6hffso3q+mLX1BwhKjZ93X6k2Yuj5KwQgVOZD8K6SVppbViz0/SSSxBwKS07xd++
xNmbSQ6gibQ1KfX9VHUdkMnnXfzvpFgL7hFX/YR5uDuek+xcyWYLS4ILL2k8pVKt
qbrjPN2/j54SNPpOR8UoFcR8nqUmoSb6RFy1SZaY2mh8fEPOv+AeUjD5IXEu3r6C
72tFRdu3yG3n8sJ5gD3n9d8A3PjIiN/YB6uieNZKykFmsewXoqvUgg/iGBwMzNkR
89MJU6QWIofYTF8qBJquYYty5Cjw8eapKn4Scn38aIHe+MjlUnEwvTqJs051omhL
bfhX3uQRICw7lL9QjiuwYVDAbC2Rh73zzA/X61oRiBWX4XNUap86h9MmcLA1AGeG
NfayM1L3p2cVXBHd0CyzZj5qH9FSsIcV9v6X1Ub+VMWXmsUYN22/hETXo+EWWHIZ
oLqHtfGl9mirZw45v+ECAq+G+zWiD3f4UBmLgYC9dTrPniMamQ072AxWn2nXAl1u
VR/uVlBYliMHt2JZR6ax4+6of12l29yKn0jmXBHnQUAbQspiuAtjXBzkoowm+ujl
kgB1c56sxZgb1hewio2A7FTUGeFU/0VonbJmd04JUfkFvvUGTNAExu2IaOLNXlqD
3PutfKdnFA5KFb9oT636tHMeHUvzVVJsa+1AIC5HhAFiY66wy5/KoD6Ov/8Q2o4q
EweQuS3PfI77g4BlBXzOR30rJnUXzdYP3r0jTbGkcqY/Ufw1qBZiy4DRkLf80NTB
IazwB1Q8BakqFBMJ/xebMNyR7ai76m1tG7Pb8qihApSGj1SQ8hB9L84QcgJhtYPv
ACQdawr4mHdQD5C5LHCHWcMX8+JpZtaiWMC+aJwq8MyMp927DDmr/T/2R0WuLqKU
EIxrxFDA3EG5pBx4NIR72YxIvdUHUuX7UCwR8ZEVqDTT/yx+1jZ6NUPQ73SGHDi1
yoierdpUymeKsU5sgL3d5cORHNAjTY59jM7Vsu1zs7vVX1KQh9OEyN0aW2SAsSXf
yNW8K6Fn4kowvefgwm2SL+R6eW4qOYTfpQ/qHGqUaNjIqSwRDlk3/WFyqLK+h45W
diXQ1m5TSTwcUF4zsNS0vVbqGuIbNZXPM5LAAtpGdgH9Lc5o1wqyITPlQddMETXP
nPWtUjIeZZJByR5woGxYC1/W3J3dKQyjvJ0513OjD7wPnlJhudvQqb5Q92LOlzts
uefLjldixJuIDVlrWtYBOa0dBv5P526EXplqc93RjSIGfWCNM5LYOYvZ/igbubOY
a2H95I8j0HBW44sICXgt2jevqWAlUhVYaEQgzMjt1l4IwLjrvah3/jVKPXGXaUsk
aCQryntzjJu0SUhKddKHdVs4T79vfWXQkM3iueLpytB0ElAqi8/KMvLDcB4ADG7O
Znv697CeAbbgLmFhBKT2Mv9WaKI3c7hrOTGoKcP41oqcaBl346FNKFr763TBirga
50T5mDzrYvaeIawJmXghH90IW7Qy5EyrnbIv6YstiRELKDN3DNX2zsS4fh5cICSL
Bh6C0Igk6j4T0uiQymEEo2LFxUmHOOi3wiKv2P44HJPFrunCI1lsgYZzrueGnfnV
jC2izGazCMgQ4h/RZPvZZWxd0kicJ9CZgSOLB3in1JpupxF7Ip0Hd08Ej5YRb6Uy
YMgi1wBbnGLMy/rHl+dqULg3p0kR1J8yMzjicV4pCTW+606m1mtIWGiiImXu0qUM
ehInNuLpRINjjzPjgeBzSc1MMRZ0zdmk7fduzymwhxrl7nAZxZ8BHnd/wivYQvkG
u/XvPx/vkX4j1FnbgrKQmL2LJrzsma4G3WHGR8aYCFeoBmRV/J22GIa73lXJVCwY
MdK51TkBj+8ueCE2yyTT4XVMCtFYTpJtGIa0XLBF0lt1jDAKAo4P+TFrs9D6WSmb
f2Y2pd6MLT3+cYlQFrctLpKC72CagVta9auX55CeOyVM7u+r5ghUwuI45LzeURSS
C4NkG8mqsK+YbvZWtO3uGKs556rK8vKWEF9utWquA5gtT/30L0kZiA7I1yz3Aeuz
k5vVdJ6qy2u6xyjkoIPwTONAGs+ehKQOcQbJHHC3hB1Ku1JHG+d1ynbDg93X/JFi
4BRYB19v/SmdomzwZoYBcMZPoxSDoqsmxIqmz52T6MynqcG0IvzPrC4pTbVagoJV
qHvfrTgjz7gbJZWRs0yltwdNFsJHGm4K6qzb5ui1kLPHIcZnL8AXN3ajP3LZHcdF
/uT1oVg2CZVDWHr5tIuHc7dpjlMN4ZLQ3ertQjTGRm0Y1LupXkvER5VqGi3V+bzh
wb5KbRllOhLb7duZ6zLjbUykGBApUtGo/PnaZJMkwQ4wujSO5KnIm94cF4TS3ti5
/fAnQ+mzvX2jvlwreksXLAyJoRdJGhAgVlAQcI10+2NZhvZWWsyYVL7Lhk3CMqaO
vlXOud5xzSVd34tamfIBzHsL2DckNPZy1nc3kHbBA86SrN7KB+XjEm2c8dT1ibD/
qrV2A4GIOQod221lGkF8vsy52ceu7A0Nk3R9q9sbefpwS0OfMq1udXeKNLBW8/EU
OJlz3T8gtlWJSykt8SjpNITdqn/3Z9diCO3O3Ojrvc0UVepILxxH43aKPghezN7X
M4dEasuVQH0glOVFOioFnsMk66Edooi8LWBykghXkpk93IGNyLFGn/ksj4L6fQNq
cpL+A9zpeff0N6lrowjyZNVi3ON9G7VkANp00kFYA1uAZg3A0diNnIRtInc18ZPI
bFLeSiiK5CHhmCQ9v+7VufhJIU6/VpWcu8rWNBnhxrh1x08mKaloEuCGdEJhSlAB
R0Xe0aSNC9T8gWjA3PO93oLJqqiT9RlWknLSSL1qXm1H3ah2HR+j06nGYkMlsOcM
TTfGodm8+y6ZBnfN9RJXO6WzReBhd7DEq3D5KSzyDtVyolg6Uym9sHRIsE/MdDrf
m0KjS/BMStIrQ25JBdELjiH/9zg735YGQcTbrDadi2jn8+cgyGr/qwNg1vY1BRpp
UOpvZLDOQYTopnKrbGpJGhoDWzTwjrLpXtMWQmOj5Jnh6aoET4Tcg2R2cfenxSaJ
deOsmFeGlptRf9npEH8oDg2A61aSorPvM+RzyeR8OAMJXR2HW+r6OXlMk5HVA4fL
BR7zAAd99kOYKe7yD6DFg9ddF2/3mjLLOUDpA6tX1gCHo/7RmyoVwfFbG2lLBINc
nRji8s61Zn0H+y2nNSNZOYAF4pztCEdK4tRX77JKjuFpvnb6CwjkanOn8Vo0IXMG
C7GtIp2XzIkJVxuBZydrqF8+wrIJo6wbW+0fN1bbds/eON8ig/AZrEiaXx5nMgSU
QFE3rkEdgcRHjU25dwUfcT3ms4ejvWD32xz3WdLl8HXZ7Cdn8+7JYX/wGMPzmRop
eDHSyoZlJymnxEkJHErlGoc43aPGLz59pyi9KFMrBlvP9+DJUmQih2xoC4k+emy7
OB4iv3tK5+6v/vtQKceYfXhEu3Rrcyz9C2BZkqlWc+qidItqjXK27oIvom1Bs29C
7MkqmBvT82ZfBv640686FWyRs+Vu4MWw0sfUaFS0YJ/dnFIqsA7xL7ycgHcImT1f
5oz5Nh5gxQyUrSgk1hp2+QbBisyo97kfx048MzefIpRrBRQ+bxWHYwZltObTt3th
7trSpuf57f93I99IS56eNUK5CxWBgVfcPg4lVFMwX1PxyNYiS1bzds7TizeXF9hp
hjjlyD15LiOs8IuoP+8Iw1SAZugDcz9c7XRX0K9O3LAfwalw65kCZDtnLY6AYJj+
25leFTl+dXRqhG4ojinWG8MZz8CwRh7xydcZAA9rhcnbjguSQ03B5fusAnqmyvbz
KwCe6gOm9DPqCfKuIHyfwJtlai5pxSquB4Kx6P75YK88tRX8GUB+AZOAaSDpo7we
HfKlABZZA2o3W664Kerm+/PUhF/cZSVz7Sjv2X+xoxktgunpLR++xyfqOOKjQXaF
crkIk7hm8zkamfRtfvij3vtv0iGEbXXB8a6NLUvZkiS3TRuQ6rmBrNyjrODw+Pxd
WmfiRJ507oasgdIFl4A3+MtzfDZx2r6R76JLIsExphzU/0tvawfZwMLREoM0aeaJ
m7W+jFQqz875DENNO1hxTJpuNo3j2LQ6LHn6ZtjEYge/jdl5CnOfH3pf5WpIHk+d
sAes7XspIZ+ePFK1I9lJX1171eC2DNRn3xCHC2kKGay28RRSaE7WZmzg65ybfFEL
dE1nBDvYyVRv17sdlw2oFw8cHz52dIPC1Bp8F3l4SQo6B/57e4wJNrmkCbG9lYtM
I0pmb3RdPAyqZObtMxKm6FzwqGUrGgP0oc7mnEtml+LmCPHFR8JQfO1c0H6SOs+H
hEYtcDOY7NEXASC/z/X5x3gm0q5gD/PkkBwtO2i3vDInd9LbwrJicGQRga3R7uOn
Q5IecD43rSOPMjz0GjIV1SzJTd9fS6hpI6Z2gbqlhXebUgVzGv+Zy13Urt+JPi3w
VIMme6xhyZAABc0jo93WXlUMLEFBHTzvfZ+CaLIT00dUAgNkGPey9cZDYCgVrFXB
auBouThXCIUJXCqUFy15jhuT7vMozHbYXvE0y2P04zhxqaIHYitPg9D2zSQLn36u
U/0bLVWDjuHpxOZjFzHi5no1gy6MvUAeCPDGWyrTWje85U39bc9ovfY693KB3phL
fqrhQcPD0BnZ/zAOM1F3CD9reHEGDNQQHhXIAJUEK1xj4KyoGp96HcfmeCUrmA1/
LDEHhypAfuLQpkKNXnAJ7jLeXG4HwBkYJeZ0kVJu7LE/WAf8/H7mr4/2HxX/axaG
7V4CusTjLXCLMIM+qrqeAZLofdUV2nQ1fCMkSp3pq+GCMaVCexq7qomz9vfpStR7
GK2EEHvFEwJn1dFOsjEjNdBdcpB5cwED0CeGOwjie7WwkxZTn+18AAkV/8wsnaWw
6ZcQmxUFrGMLJIJBBI6P83mD/qzE47tRf5czvCKk2rhnWC488n+1C2GnyjfYgmM4
dfS4QSx8I8gQEK1l6YgTccpal0cxXCsK55GpVFkahzzyYvqr/GLhCcylir9h7O7e
5HuN2h0EusNPqIKDZliDoa7+ym34qN84E0qfwngCesP1rXikxofu0vs6WNxSHQ2T
XaAcSrJOzRcRwGHj0DdgYX9eNgidnbYCs1TpTjhoHisaoHlFNmk7q+973V0XCTga
t8N3ufv01FBwPh76bY7Zleo0thoZA7KLrB+s7N728sm/kuuOKuRdR8IkUk3KECmy
VvK1d2azB6YKMpGQZ04SVf/N2db3HU2Mhum1UMg7vGxSz+SQL5DwbqWoF1tNWHeF
x3m8+UmtsJm50LcczdttmYfKyoLt/QX1jzGzcJvHJ3JskJhklgjKGinuvBJnhVS9
4w11d5m/I0vegvJMK+nCGn9O5XTIt7RUV8g4sEO+SShdkKEiTF28HEHlayRM09B3
KY6aH+eHVlU56m7d6NYVp20m/itin/gIWpizoeMAK67X0cWK0I1tIXZ8+a5iqFZ9
GEp4uxVIFdJ4hu59mQOeMb7KJVXLe/2zjmvXmryPCcZqAmAwDsvhyW3zLkiOtYnF
n+1ygwH9oPc8PHhg6H/M6HOsmHxYvvQ0REeI5oeShV2vT5EPMegFsiEJq5wEdGm4
nuxKwyUDTZcJxFCfIeaEaxHTAJl4r/5yf6DELUIQU+tTfCFPD5+iNbuLN4GixZsE
OCvweWrHLMn492crHRw8rkgUeUe6rgWL6twXXth/0AasrQnW/JuOmCykLA5rrSiZ
D219+Z/2D6x6jKMMKvr9OQH2/OnQPSxnH0d1n7TmIPPJGU6I7Y4sYJmlohBvY24J
mi4X9qAqpQSKkXKhpcW08R0/yVTyVc6galgeNH6lYfXv9jLR8ui8ZxoOP3wto1ql
uifTSG7SEVxpR44sJUtx7XPySclMC4LxFj4z7D5rhLJdloNUSdA+ne4GI6J4bKl+
zHLvQK+EBPrQagSS1NDZLnhlbxdW4shCrvQziFec2fLzcMDyec/GQ2HjXG7QcBE1
uu6uaTFm49rFbh5uGAxJqd5eUkCxeaeATubvtYrE40YNRdVfJiM/2Wv8hKZi+QNK
30NU62fdF+EGXijPqad8kfsn066GMYkWQ+OaY2OYSiTPr3TRvcxUs3ptidChwY/1
vPgykklX1tTrT74QruAZR3vmBZpnCGq+l2zrff9xxMffUB1zZKnAHAEIe6PlRnSR
XK8qyqK0Hb0QoPU2q3wUhRxELMouyGoiFucwrHiciadkeozOnZ+J5dThpGD91Ftf
E2HNGMR74KBEmnBrzmUf025/WxmNjGDlg4cOmI4wOWAfkYdC5qHo1b40oEp1SNRH
PrL9kEkqHbzmQYfeL4Q2XwTMXRPchlZGkCyd2pIwp9BkOqvvV/x0/sisd1NEVogk
lMklmiWMVteilQysmKyCFzE6/LBIPLMXHENn+W23OCX3QKm4FDTN1Mxym8KnJywy
nIX6UBB5euTfkfr2b3INw/d+9VGHCmcAXtBkv6MGWoBWHl/VHG/6V3XCnxBdBe79
q9/w9IfKsvQTGzk8cZx0amJ3OnfJkGvuE/v6zIbiJf12itd49em6ORHg7scGbMKG
tSEYjuwY26ebOdEJfkVt7mGkc2ISNsaA0V/fl7Abl25s/+hi8rlr3NWSbkBR4ZdU
63PMUObCV075CNNDIXvqk98oMMmNfo08cJMElBTIQeXUBkkJu3iWPWN+kG45T87l
ZDdBW1gxvPpnfoA3gTyL2voPOfdLsDDseBuqhFfHu6Fv5OIyBaYolYHbaTiESvZW
aVy9oURuEAJ4bW1RTHIoaw5kQYKwdv7F6uM7qeUwiu0AAVSXGxxblL/nMiCr69Lw
kmP3Q3BIX5k4i6AhTsn29Rp7LCUDR6iOenr27RRqWhjr6bur5qzq7Vk6GePqJj01
TqUpxlq7/SVpsPTo33BHQLiP5fCz/ehRgF21JIsuq0QCkPlidB3HW3vuBVnY0F8e
g3CSXCNaVt8wJdmiMPhZVWIJFnTPb1U7RnhL1nycORYWNvj0OT5mhgEoNQslnWP1
iqCa+vSknlUZYasnZe87ateXJSf52tsrofhXrSELQxJMY2jHtEysL/p+lhu6OEjm
DgTVl9aycrPKehfQ1/GSaiI8rAct8tEUErEuzIzBRWXuj7CRO50KkJ3C6k6itgyX
yTy0+Fk47WmuJLdyYTSILouw0w1yzYQ0Yb3LmZq7dXb9nHGxmJSOjmgm0mqIy1+C
HEZMab1I7MnM/kwrwDPsBel7Fxqubb6xV3WANWb8Q40c/T2LgAhIt9ib02qEsdr/
1lYERn1Et8j+oSEvsxJ+B48T8kz/Y9GLkXhZkaBPOKSfQWaqQ5GFtylHND1YO54y
wSmvcZI0CCTTUxUsBNgwD8mEvWgFGZK21mXSBPxOD3bDfezxZ5Y6L7crswEI1KHb
YBxof2C0qZ/3fWW7gD1d5qmNlIl3PskIJO6y2AXYR6MK74O2vPWd3hnRZd3KrEfU
Uy5mIqRnydEbeNBTnOlkIkEPLedCUmHKETHhAnVlm03ULljY72APrLEfBDNA2Db+
cfi5z6gtTbxnUjYcRIQHPc7nnhGZqYJ9wV7rxSp7TQoDkVkdfBoo4/e9P4freJPf
JCNWb1ADpzIFA85Tawl2Pv3KEp38+nRpa0Ybty1IGPJX1LBAso3U00KFriTZMycD
9Yeunt0YB5cEC9Wr9eGyAe0+NJMi4LXK2evlJQCaRMrA1h714jI6y3UF1CCQfxNn
rLpX1zGXFVdTcPIw11ogTyk+l4+Z+IXaPuBuYKHi508NfsZ0iX+RzpjTXUGERWWk
c+MRpnJOp/p0AeJZSvNUfP1niUNVfjDCnB7ci74/Rdh+j89g5OSsBl1AcynOsrrv
0+Xr9nFrrbIEfwMP8hwjt6Gol7azRcAtPTiwGyDVtxgkGRmQ9UJtatxA/xtZifd2
uCUQGOqJDVXcrcEGIrnoWqRIPqktOZeG91qXeXCCIl8MhN2gdbTNFAAGkgeuNRQ0
V69uGSWiOAh5QNbRy3SixnHnCSLMkc5wDt5/ukTiJtPz+sMAlKGuWDRPKHiJg5Th
bmOlguhHqrrOLhUKwrlBkJyP4BJNPpTnGN7C9AZ0KPPOCnqQZ3oWulek0e43Z3bd
Kk/SfbaeS5YPYm7eGm4n4u7uPdKKjaigyP7SPWhUbk9yszTJJjo3TACCYphSsNFo
YGokdzUQKyx6qdcLxHJTwmrixJQqqx5QTPF/M5rN+HpcMHqZ/qVrS7OriIgfq6UL
YQmxmuXoZKdE/LveZj1FPpk4J33P2ksNBWgFmIxK2qBtwLr5+d3mBslyc0pzr3b5
OuUv+JWhS4xJ+kYi4+oh2ztMv6IFYLxPJ3zxyujlwj4swpW+U9T5hfLclYX34P+a
qORLeKs3ygYAQQtKA4uEotIn8TGKRXAQWiem+cDic/L/BTnw4V4QDHvxf7YGUU+7
cyiAErjQCJTmhTPSMs5MojtfrYPuSei6zCh0XZTIPP3jW/CZeDV+uPc+PDbZZgWj
/T5l5EP98AHUfVu8Xr2GOc/641BsVB25wal0adUpOtR2Rw7+tVEvS5jd5WW96yGx
AN1QaYlOVfU8oGYQxVbjgUXf1+P6+cmHqSM6oDaqmhLoxK9Uq5qwj191Amk+rqki
nqqLJpJUzD/IPzLUYIaFW8R7HbID7WyBKpwSFRm6QZTvIDw946ffqim9Tw5diVJm
JNix+BRjRuZnosPAF0zwkue3/5wU+qDhaKgj72+5b9tdfZroQxLzvG7IOCkX6Y3m
IMSOeBTuNDQTXcGDWBH9Ygg0LeLaQWWk7x6SJYQv6+qTYFa7LJYQaPdXU1p112wb
8GWAuQbSP2tEsfUkiBJ/iiuUAH7PwKjD5nqb9/bwYE8hHB2S+VM17pQkNLfNG/7N
6SeZPHvOi5rlpyFRYqJ9e42KaOD51FzYmTgFBJGI1Gmx5fSKY1sP6j4UZttTg73x
zF8yvVgQcDd9k7jAL8r+QS6ZJIgYNhZY2l6dhFqMlLNsefRGmyjjVWXD5hRTDv4P
XlEdwic4fiZzXWH1grKsy3L7K5sGBkYAUKDCPBUS8DZc4FlndAAKIEOSLP6PnIh4
lPsqvpfN3Uw6CYJiOPAKVgZzGV9Q1u40EbVLaM+sXbLj3Ao1rMTO8uPDoRHrTmlG
iX796eJGVQ+z93DLWpqCgRtKrSfy5mk9nNit1IQlpid2eSyBm4+VKn9Pl9CeSeDV
aSzgQM3K9WLT44CMGCFJY+4Q7lhqeCTZO1NqdmH5yDdQVpfXtsDjPFiIyaYP4r8/
TP0ez0jn1wN89WrXEHuTzxN+53PQK0n+mVVb/ZgnaZYou+AyZenHFZ4mcX7IISgz
DW5TQhwlQAmNLmcaFhG8/Sm27qVGApXcvqgYUItOekPSdr7zeDQRqT8Mz7y46Tt9
4VtrZ9GcLPVhiZtkemm9vyI0f17lgzFgZnBLacZrIOt7iphMX7npdjQquuvAmHIG
6yFps5ElT2t1kmlzC77+Sc88CNXlHjlQ9wRn5evWnHXYubbISwwRvk0gouyXvJJ2
c/c4mYnjZfYihIrCtztTqGaykf3xywa1bNTjGz6ptBPjbxBb12peuRBOdpvyvtfA
F2UaUaHWmdOK0WWT7CEyLe1Mz/GBArVmzGcHPxT/foMryBc2tpcXpqRMn7RRCSDU
P150XLy3eUJTIucYQCfKxhaYKTkR2e55DYvPPCB8LDMfFVc4EiZAo0QD0VzOGrs+
IQX/Un/lpFTjCBBb/Uy/KbJWsXrGwsFVFvJAHgiSD/z2+0czDRM5q99byv4YCD04
B6fpaZVfK0a+A76P2qy9iOyTjWwwjZlyHglf4kqbBpgQ9f9Qp0c5xX1OebSQSfjB
jKqR8WrexQPOF/n52vMG7TJ9d+Wq8+gjuZ75er0Z01g0TWe2cqMTgVkY35d661of
gKNQ4kcF7O5ie3WPPHl3W6dT8qrsR+WrrR2GvSSN/4x7HCcm+rK/ZZ94YtBG1u4A
eURPFoZxlp0+L4cYr2ICymJK4UNhZbsKSkVjOBDa9jOBngEQpwtS3kmfArkBiGUq
BgVa/Q/a0jqImV4AL3KhtDNf+0pVzilpsVa0sW7cWhZ6c5MP/J5V1azZ0d+I/Htx
Oxj08UwA9ojzDq+C9Jl9r0Py3USXBlyZomqW2fPe4QJwddQRqfVtN4dgSoBBuF/O
J1S+Lk57IkXei7LiDFMLo0cqr/WTQDU/Bxy5YS17fDFpkpoYjPDxZTAS5jDR3FOP
kw0bY50NSEvRYChsqoqSG43eytYqnCTtGW+NoC6g+/TS+TWnYW6W6HSEM4bauapP
3mUVERZKYfvjJCS8Gg5Qt57OxtshFfojMW3+Vnhl16Dp/2JZrDxt7lY2huDQGf61
dDDGkol0PstVtLClhaPZStTUe5EQGZbxhcdnzjCaGxWN8v9DmPy8i2ZiLw/i8ko7
OYr/PiaROfW9nswKeWFVXHkrFKg/VZ/Zq4tRaK2bomPLZLkk2LvtcXxXYlSNvYaA
5TXj+vx0YNAzgr/yCszqVtGY2pyXr6oWHsK64QxX3MnuSPVsPmeJknBF2wHYsxsv
DiSiaDCvljW8cL7i82Bqqo+GVykjYLaXQ5ZLW5RGcJeKSXdrjTH6/IfSGlSVbNgz
g5E8lbKG00k0MrOdYlusiLMLMBQqyk7g/AhQDSPQZq0Oeegejw/9kvw3/0z3cKK8
ZK1CrI3wiWI9fcSfco56xUa27jccvKxQZ8o6BCLbo75/ex9vS6v0QMyP+uK3jW1P
+XzY1Yz5HzrfxvMWTA3hfMA1I5bZObH0iH7n2rB19ouSeKRaUYhdQ9FJ91Bg1uUs
EA8e532FyHWERsQGbYVwWldEkIwox7rFPUnEJPIiuSUlLeoePnj/P7cjzZBHcBZs
sNdaqehy2Ni4TEZMGbh6q4AJ+9y302WuUwTLGnpU2Em4fzliX9P+WQha++FiiwAL
hgycX4NJwcrlv0ihymvy5abU6gTkJQh5CA7tgQkMuJyps35IGYp98hqglPOQaToM
yHpTrItpt56VJ3/N2dgwCTsP1W6um/vbbfgFXl7RXwBP/B3nq3uwIILwiHbLDG5f
xKBV6Ck/GI/AUwBzbJnYuN/NwEeCZt+fWJv0d4kSJXdLZaLYR97yCj6YHd15ZT6k
aKGAW587IeMrZNgyWd/YEqCQB/skNhA2Kbu9KSQhkQ/9y3TYJQrRZwZiE3PrvFUL
jUcNH96hnNd2Q8gqiH/4trk+/nyJu2vgfLFVEMjFzgkvQ9ladPt6IffHqiYillCg
7fSJmrHoG00qCwAOqsZzAa/qtdmBHBnnURWZU/sryA8/5pzE86j49N1AttkxNvBm
Tv1PimtTssx6b9bfc79plhRbvdn3S6Tb6em9so4O56UJnc7Z2RGl3eduP2otGnV7
AJ3pE9cb7HkI+4tH7WIhdWZwYVZStZlhzRMbjRyqmJITwT7YUfkLUnnUQAqOJ0cy
Ft8XDQmnwCT7tqq+yMa/C2kJbk26dRg5az3jzExdatY990/H6AZ7VzMiwB+yPaIu
S9uko/bcNc4fsxT/ZNs/JC75IoRq9l2QE5wgeIbM47Nd1NSuY6vfdFQX70quhQQd
pkvWZtoOvlUOfiZt3JiwzQGTMpNUUWIzBU37pMlXW/XAlamUNXxRUN+E63VqfyHP
SanhmeWYnF2r9l+w/qP7Gbg4+SbpjjANU01m/bUC6H5JXvRqoFIJyuQZ3+yW1Ksj
QYZzOXOeCPN3KViCZMqZpkDVVs4tkiM06rDZgBKIk4HaeKl+LeMrZIt41iF5Odog
1dHoWgo89RcvkLMh0Q0GDczcZ2IDqox4eg44mVZYNNFihRgK42JH/pYQ9UMxXbq9
M1f1QG2TejN2+xfOPd7lfugPmRA8vLlBUBIX58VUa196xmzfqLlgwui7e+o9kkMv
CjP0MxND6URkZKK1ek6GJWVCuxp3DWcnGd2vZL1WFlYjHdaRz98A9FbUsNAAqojv
17APLFwouRouedrCvsgZXUkOpBuu0T7fzqUgelP4XgklKxJFsjtfZhMl9HCfaN9I
6S/Jvr6lvJpPdGoXpheY6hxW4bMTtDnjTto+a4aRRCirNqUG8Uqo2dq3vEUmL6VF
FhDcITFD+4b29h37G1jJvxFzOalXMNn9+EtKOQOaX+At2xOmSK+iAzPzJVXFWnPx
B+6M9Srd0PE9x7UrmRkb/hipN+LW12LArvv12qRBF7gmAsak4fulZYfx+d/ugBs9
g/l5wQOnF7oRoQZxPlCyo6kUpE2Jp95eBzTQwpKejHdsIrzqln440XsKuSszLPKF
perDPQt+qUDM9K3AAExWjD7IsraaafgUTqVXIoyzEaGTeYHzXfdCQ5IfBMbe2iW2
SnVCdjGdwoLv1v4A+03H/14Kb0Goc4c0eery4TQU6eNOuzq+FrNrmRYShfp3c+s1
MgInwoRGcY7+yD+qLeKoT8X+lwY9+hyuZ2YiuoZcsKA05aWZRGFKrkrQsBHabsi8
rX+lCqjOcx/rTb1HJK7lhLTCxITd1ac8ENyJ+fiNgxBtYJLvIRBQyBtAxdbmUery
6YbZNFL21dG7iRHf1N8cTLQrDEs+MBC/04pEUKDqPRnkBhth2VhCdq7LYaFNkBQG
tr0cgx+hWlhFfMAhSfGY/raUoco8V8r9WfAuZeQD6Q6g1vM2lcDsLCSDsHRRDiKa
0dWBnkg0gdQEwc5GO8N1EgyRWVJPF/XD+uvD8c7mImAYCOiGHJSGoRxAUj/MV+vl
2JUF3Z4YkFYOtYuzOP6jYs8kJpT/gMGrDpoBWLQHqpGxf6BK8twPXcSN7INIyCQC
gEqulqzc4JOiOcpM16RJ/VctE39vkIHg+Skb1TSYYhVKAdZ8Bq35qt7308UyS7+1
rFFFsXjdKCwQhVhSbuUGzoGCv2JmTyVV/FW7wwGbFnC24ba3TqQUM33cDqLhaRPX
P0A2xa+BKyYDHIVWDD656wZOmkzsnSASPqfNVqzmXQ6UUo04Mc/31//Mf3C728Y0
Z5l+OJIvLIJBVBKprwisLLhrERGSofGFozu3FaRLp7RbaKtKjyddbNjejByReUpL
PCI2Bga5QddBFEfQlAfaRssbDBJ65o0IIqRLvJMumByORtX7iDiDb00WaIrh70HE
kwhaS5xNSo1kts4I6u1yCKi+9iwASW9Jh+28M37s7949MpolsCO++Sp1cieMKkcN
xVA0Een8cgkCrfKItOPTeYY60+cAzkpPmAb1W6y/0K5Y1vfTD+WH7yPjY6zxek9/
OZl+8S8pnfYxAog7pT1UfakAOMPStOgocMTgdvtJTaJVw3DFZUMmcEAK0TFIS/us
9joMhcBTnbH6NaZW1+3BmYetXWcCqceQZcSb+DKzRj9rrsLuZykrD4lHxP6KNfiX
nYFtFhFOWB4Z6+Ix1NHWGj99Y9C43tjz8rot0GI26nKi2aILwqFnBJzRHh+ZLTR6
gzd8Mcb7t2+d36m/QkXixWEbgJzdUjGiScMFxRqVKfChySp2XxtivQW5ClU5Ae1E
6/0xymKSY2kZalfs1c5nXgbd61hYkZCMFpeAUR5WmnG4aBiFneyJiC9zSYv6bKTr
L7a8snplncG7Xazb3v6eHSlS+RRNu5xJKcPH/3D+NKrpz/DRSD1/64YBDsNyGHr5
0RQlgG5TXvD6N8Y/CUvLFs1m8p0jsIoNw7t1/kJODL/lfQxld99m0WZFF2+oEPda
As9kZGLVr4FjRaNFLRpvP9IaV7oHOJ0Y52uLTMiTwEdE6u/iJIvTdeMUJS3EhRGn
dDG3xuWkt23lfCRMmE2UEY3SgwZQmJPqvM1qFz37XBn7QcHZTS8Mi6TrQgTg/7t4
J3113FCtccQLrBDrZCzsiV/DyrRcZmvmRQgq3K3lmfxMdc/hm1Ljy91UzCpchCqG
NEqZp74oJSId1SmMkZb3dXdErXdNzMeCHDUutI9qTByaT+jZsVpWkLxOxARNYcfJ
u4ysVRPGZKQBUMEvFp8l0a7gDFJaD/RcxJL1SxZCho+lRVWZndKAvQI7m5Xp4U6H
IC5eSmKLIBYlh9cIssYYKBlacRUyqleWBKDMifTvULyYo7Q2V4L2QRvjQ/z7sCTf
kfwJymDJ29thQDWRjry5DEefB/jCsoTCwnyt8RAeahPsR+M+MMn3cBPvXQHhDEVo
9auvcGSt5+UbRlFx2tuBosqTnQKYxZopIbKRF3qr0HfYR/s6wlSajzMPMIxwjNQH
R4zunAmIftf8+iMT9ufiPwNO5HiwZOb0LiHmh+wnW91McCAzk69pHez2laJMQqCz
abPprceEzbP1BkCUsSPJGKFprf6A+NVCxZ4CNVhCAY5MBq/slbZE04aKBu3PsyXM
k7VKk01mpiFLgHIHLilwHTjCft8s5yd1HbRxgIPdszMtJRwwYRGopNBYl3oqNBlm
DHoCa2CwurlF7idHutS6HBq/qhvBXjjNat7VR/UyUO7I/WflqEyWpfb1NS2W8Hrn
mkrb3Q0a909P/C+V+T0JbGWXA9dbq+zAvz5QSgY8EDIvtLjIPyYfjYMwQv9OZhi4
weTh9obJXg9pLR5prXefyujLcg9kP6/U/kl9mYgbtBnl8lEvfefCEvEqUaxw9k8V
fP7CBnuwX1YoKIP0GnlCnH9Nceu3IehaRwgY4cwVBO/XSGgm+LgrLB+IXUZLbATL
00k7PhwK6xmqjf29UiRw+VBk+a/oT2e3VSGwrvy43kyWJNPiI9XFfW1xAAh0WYP/
YANHoXTyCo77DY2XTiILW1KNrIzKKsu1ibGugPAkp2WNje2RNS+8+ixmylZnQfI2
C9ClZMdFRZNSxzj1dCPN3vAdRlVqdvQ8bh7+p9zCU+HVn0U3nfXhcIprFvW94Bto
cSXd+TaC6V/jJbNetfT+mABo879fvTj+5OuUKHKHpioCZ9WijKyf3sK7pr786alI
I8pAIzPIDNqx4vxkpsshNtKJhd/xbBitEfeRWver7MmzpMxyQNs2VpDwXAqaLtr+
JNQHXxcDVmY05d2ONbi164j3SWt/K4tCaKY7WYZId+Qj00MHuvALjST+wDov1Yoe
aPMeQnJyowvDNS6VhnG3XKfpDi6nQ2hPY3kwtCWi7PfgO3Enk5l8RYr8htTFUySH
EX31n3/a1mKhEnLOfr0uMXJb36ec0CxVcSTeX+J0fgmVHCthwKEaJM6uZzgqt2hI
+OlWaw8JUH6NntBixAOGZf2ptEOi9jeU1b3VT8HtsGAEyRhz/0hQUvVeXPhaJHG3
ASlFD575QL8KQEtx1GR5ab/qfCfuW6JvA2Q3BlHkUKJ+Fgwutdswo+0pTlU7ftXf
SmnXb5CYFRchki0LrQfDzxVyJ5Ho5RU3UzYuv7j3OcLbVTv/m3W1CV/QjpDRVLHa
YcSpQfSulwD/k9RmWOoFPpdC6lgZWaeF3pHoNn47wgdi5ft5nE+RDtOeAenxUH9c
8pEFMBwxGwrnJTpxm9nxxklhQ6aUw5GQPGLQtn43fFYGN1vsMvQa97O55FisoLZz
mdz+wkfGRGLsNuzBlldW9lFRvQtCixhSrVgZUhKM1h58st0/Jmev5ZQFKHblK8Oy
Q5FubFNJ+Q8cOK8XFGx9/7feEw7VTfM8eBCE/4yuibUfoCxbQKr5D8aVQuSbmSsJ
x8hNt5IfGhTNYvOIZAza8VEG7AV6cU/EvGVXfql1ERFNKeCK2aTlTJ4a5rev8IuW
53oRfxDhirtSDpB2A4Sm80sdSnbcg9UW0vIMCan8cQaWrXk5PIuL9GqxKIity3qU
SOIKYhFGY8N1EgprYRAKENnpgWNO9VPr+MClT9qR8TlWs3cA3Ihe8kDqGSE7dvDl
sC937IYKQgmmzVq6nOmqjA7F0ucdfbRkajsINhWbMCLSuTdo15mYMK2kbZShjSfa
mmoPhG+dKwikFJzR+8omo3flb8uZchfhzGYzIuK4+fFVMHLW/Lwt2WWBMxDpmvQr
GZcHs6s8yE+eJVDb/qM4sLpssMN2avHiUdi8mAEjtZUem89badI+Jd5xJsP8+hxA
NrTWohROB3Ollc4gja6htCxCkTCmAJ4AZR61pcXX4UKvPQesO0ZVZbEbqJDGUS7t
8UbOu+sa960hmAY0vfPueyV+Leq8hOsKmLRVpiXbjVoawvvqrIFDPKiJbUOfVKlD
HprQuqo5rVTQBpEMWq7ApvaS99tT6CAdy/biyXifxaE9cj+YfJ5lWaIzW6iF87Q8
iaHDE8vSUIs8m8S5YaV9enFqZxRzD73VoSETrI0NRkOpJoi8K5MlT7lr56ma14GS
ZjjMuxiIC0vJNBnWLSI24xVN2Q26nY5iNdmBSefAqZkP7DdT1YEF7r8VqEIhQr2k
EWyroO/v5Nw5b3vCrYLwTSojd7cofi1pGEHjGzLVa4d4orCxMI7Ve9DaqUT0mi9x
81h/IebqZtYW34vwxihsM3o1qgUlNqkR7dFg5ZWkAYt27VisvBcuRCulqM2Z1Tzy
8GKtPeQrIMiwUhKhYXlESVWrc3mzQJiTprhw87jNWGjfCnD+XBK8xsSuQjcu+56f
cc2yAYJQucAMSdGDZJ1aAAzhSEl6CXe1vSRqhlkUs7GHFO4r2QoEWk+AvYElBuJf
81GEKXh87P7Z1HJ0igl4CWVOcAi8oSvpYqkFjYWi0Z9mvVkFEGhNUBuzcFhNjE4x
iBTUc3Wpp9ZF5s10qX4cbScuykTWJ9MBEJ162i/nQ0mjUVfeT7X3WJ8CkeidKLQf
HUO6XgCmqW915RLlWUsImZ5byEqUV2jqF5iWzeB6nRstmico5mAdOaxKMMx1rJ8A
K1VR6k+n6EegJGHcmvBzbJGfUEHITFt+42ggHBeTEvhoou6Nq0ywZjQc5m2eH2b5
6DSKj17XimRDFkkwSe8bBalOzNkgOwDuoH/tGj4YenAxv8PsxA9/G/auyrfsdz23
RELypPTkcwcMlPob+ql8pNlQE5iu8bUm6TDn7nw/VMOVePqFNa3W3jDpugOKcPh9
pa/uXlpDAbf+byjnlc1xvGJs1MtPpehJ6UBalpeXe0Zv12dF2t+5ZF+J93OONhTQ
dLbFzur9qTP1UiywkGTFB5rSYauAu0BMbHhuGO45sKYPFamLUnyNMf3NGY6ROzq5
R0mPTN5yujQ6OulJ4q+3VM6rPUFZ4M1gml2wnnoqTc4WXbo52BPc4OE6NmBIhLR2
2Rp0XqTdi/F/eiWu4DZPMIN1Bv2pjqSBZkFcGYjukk4EsawBqyI1MQQZjPRWFB43
rarAJvH16DVrBHLq/Dnm0/e2D7YNgyZDYleLL2GyGq2M2gWp7R1wJnLtt8Uh1gI8
DMJP5R/rdSkx3SEgnvsH7/x6Hv3w5EGBzErgNT6bQ6UeITt/XIBD2g/n0t1G6unb
pF0phFNqeMI69EPOtlxmVRTPRL8o14og/8ask2ImmQmmnX1egmnNoRVjdZBW+EEF
iJu6lG3g0LOvoGwtTyeP/lYp0rjC6ih/VEDffgYvsBxu3/24qNht9N+iHznfXgto
VaaDrMhAc4btEmjan9j7CFEz8rv4xDCDOsc27it5i3lIGXd9TQ/mP4pAyla1eX96
BLFIqMs/y8eIPhdoZJhFc0BpfvRzxMGKvUb44AxzRIInFbvZjkDnInZ4Ruq/6612
qMyzYoKZb7xnWG357VWTWVhNacKpW8yroh0M1wgwnH0dgleR1g2BDR01v/h+jdYX
L6aYyfxEM7B2l2lkYRBY69CEbY5jz5RoHaBZmXE/37Xy6PZfGpAMR04u/9GmqyuC
clANixpS5n+ZiGYvu2R9RjeQFlqYEjR1349DKVuCysBauVC7yGi9sJg5zYNdy7FI
YY6VP4B5SDMCnzPI+jvtVgWDiBKGL3Ty4q7uMIMYzm4t/aEOtxMdhjrU4e16DNcC
vrFk635K7dFj1QKVZvzuGxQhfWylBIKEELfzl46rs+Dc71rkd1z9gJGz+V+aPQn4
mQKpnoOraRzhBzku28gVODCyHK2fyP3/dPu8MBBWeQp43kMifmjPN9BnYkg8qktj
EjAGKHGZ0U/Yb8U9jraS/Ndtz+bXQN4ONtwjxfiNQhEZ7Tl5ZQZWYr7LzNOsf2CC
FqGyucQtDEn0VDiXL2pTeK5BI2ic0VgjYfggPQeWfDOJ7Frr276dTfr9Mp6dWIUG
ARWWdx+rbJlvbT3tEOU3pHyVbt0Ja284oy77m33WYTC44MK+xXNvjKtikfgzEFjl
teQogsRg5lfxxrjtmKwAniGUZmxLfwIifU7/EZs76ssO8BPUQ4pYIKKgONSXg6MK
kfZ9dEH+LAKg/8I/JT4PmW1CCEiQpOIzg64nc2jh8EbCf/g0Yn6jofWjRtJbt38I
hH4+S0gqPThKQ7vWMkRKB/HjVmJlzTD+23j052Dyk+i5uFfmNCmjJZk0ibxoqWNT
xXBrqG6aAk4oY5ARxgSQ+Q8cpqNfRtLtyhwWjv5HHQZwkhHQ8xKrkASM1Uqor/1s
QAaoqrcb8cPlcumP26qVehEe6bQdIY3EqNFnzyZYrZwPYRBFb8cSPiQvM7aHlJfJ
icAscXbzDGisj6GWr8bsEaQGWZ8A3NKlIyiQR51FhXI3Vz0Of4XhsDIyBVeDvycd
dJ2mP77aPEl++D32mRpiIErBADmXDef+M2cGeqzu0FBII02TgjDtXGkrDovULDBL
dGIbi/juBejq1KlcjeFVcrO+CFwTTsfnVtYXjzKFBnAHZmx1WQAwl/RIRW839UoF
nqx3midVm+NzEaiRB0oPoCkU/pGgsSIXUWdwLaJIVpr3Gk+uZg2T4UaSTlC3pWVD
yE44imiWlgsMVNF1yxS7cAl8Os/N4N2Gy/0CmXsaciRW+wGqVYrt+6rKiSxzYGrq
wUABA/I9eits55+xEyc6Cs9rZO5fwMMRh+qeiAnk8kKgZSDyiyeyVXa/R2rHkVwO
SUqwf29KzhRALXCS5lyv1JmvLLRi4zRuGwlizZrGDtMdwH/9C7tLKvQWhUPiuQ/a
ThZ3WRatAgCthW7VXoAcf9INNcnbpNf7X+n7PqvvSelaoFQllessRmTJSWYKWjXa
A3FXr7DBBOyKiV7Z0dhxwVbcLBf609qdl2sKMibM+Lf4cL2YpxlG+d1EOdW8UYap
pOYxr8V9x/hWFRRj9CENx5xOa87rJ/bHe4sZXrY1vq0wT3wD2Fi97k4BInRBQNVN
11/qZMP2sZY052kqM6gqtSIereK/IS6CI6PWVOnR4+Etyx1ZVc5ORSYqHxGqhqrX
D4FiE1F11AH+TuEhQ6Viuq4MttU0e56vc3Mz1wmjkm+NYktCuMst0OcHggdoLhTq
r/ZUg4qPTNAaA+7/jew+zc0La731Al5gsuiuz+9bx5gHDfai+7n3Sf4xApnd4EZt
00BUlfmTGja1X9DVb0Bl3JfEhDVjfNKjFVwIs1zi0QIOxXPjIijqi1NkrnFsCcD6
0fIoGyJoTwEwsXF5ndTlhcuKNsX5h+vmn3uaKHi8qNXUIZ3mct6iLa27FYzbHTxN
VwFRDwK1IoWvnu7RNGv9CeYOwMwPy7BtzEgIlPIzOT5NMnGJgyGvnP3kK1AFcBVp
Flo8uLl4XKwBEt+HgsWYftDVYraqcL7/4D9x/PSQDc4BMSPYdtQXxz0i8st/HhI1
/+UZrz2yW/Q4Bpsh429nwXfaGQUvE5pCX7DD5GtwgSIel5nGfT+uHy3YOrhAPg4Q
mc0GTQ0q5nyxI2l1ctJyCoZ0C29Y3vOSTVfmcUHRLaWh1FhF76Qc79jI4kpbQOEE
YbV6WvlhP1QPCoF1jdA2ktX4dkPsQIs5SYCCxQ/qQC5jH1XyugohcAqVOaPc9OrD
bUocshahd6aV3e25uXpTwHszLcx7nyJtmmmQE8PbFRQo99kwfluWO/Yz4DW9L1sL
TgwpvFC1pH77egM10AIMiR/GJhR7lANghCqytEXUj9Np53Zda5dh8NZ1G/yis9zL
HhU/NL2EFrBv3/FFugvhCYazk7q7Vn/G4YuD4p0c0CHrZkM/pX7SJX+cuOwFQ9ED
QfdI0RAIiijFGMiyfdRb7mG5urcXkw2BRA8Qni44GoKvz6FYYdK5A0IZ1+u/KpNO
fE/7bR6WgmObJ2U1faOPItdm3jqVKJ4IMnHlsJyDP41ev0JtkDn5yfXAcEjVxTHO
ZOoGN/ZDNPUDwwVKd0RmvVg3CK8QkyKCegDS3rvYaONkbaaLWYpcizjOISwKAiNq
UR5l+t7h5U8UEorr3L3U5abXHqXr5K20heaYy2EPYICaoybYV52+o2L70Pd6KClH
PMm9Mu+4chg44MaRjDqgU4o64Z5yc/ihRrDW86IP410N7GUUON1L+Ch5k/FnwSE/
X41ySNC5vhQiCVvR07Fto59uW+1RPpFgAMreRBtHOvcx0rS4ioGPSuGv4y4QEnS8
L0o7hMimNtPA+6g9fIAfH3sq1szwWLCuBWxUsf0pqcVnKpb2j4HmpJ2vX9UNnrKC
1s0H7L65rtIk88ePsDsOJXxCd1/3ZTVt4d7+291v0xiGhyAM++rzjVtjXPQE5vb6
iY/rwsNEXpTJ6R8nQcPWGeYPIprtrTWY+uN2PIOT1282ODdHHkRf1Jyga+JPsPQ7
xV8q994pSTwo2p3QyrjA8MHofFDs8wYVETfjth98ZkHKNy+wpXkSU3EQ3F4mM9rh
TUp4qd3h1zIamfEJ/MDz+2YKRFjWH8MwxWOk/TGvtCAFg0bXvOtVCdhAC/u9ytXc
dYev8TERtulEj3hgRj699YOxJSyGascd33oaJ/WqlJUklZ9DImbERG/pdUpJ/PBu
uYSwmaVtl7OPxjoztWDKbqNGjXvyyjm/jwsn0ZIHqwUFX+vVLMHXT7vIfIWZEMW5
qvpjKQvoyloImpyc5o3qbXE1TNusJp/34PAXjyAUy0D5mTQQ0S4fYfdAKNFIAI/s
bvvaWZ+I6h8yc2yGPl1qm52zwava6PNR95pqOWRKgO4PTJttP0R7Uh5nlXM1xgvx
qVsAdTBJEMYf5Xb+NAQzPf8BUunDocKHQ/gnWHaukOvhiXVrP4wih5zyo/VTkizv
B5IIAdv8jqDhwMEsudaK64VqlHqh7d3U1QitTb78Zir5IuVYntlm6sAfwe44MqAh
axmLG1G+mmIQJ5bQ08xbtAAhZLmC2J9Gl1g//8WjkYbel2D0BkQOIXf+YwhAN0AL
KHxc8Wpbx1QU9eqEECVFlVmeB+8lIhu8G0eKAcsGagFIh8lEHsFW5m8BVsfjAb7A
tm8yLGeCdJqmQp5tFuxTPsBFgxWwFxm/L6/yPonbfjf3n2pfCGJJBxLAgHqS7yfK
pQYpECLRSks1xVBfL7/2CeIJ5gEdQN/KbtHxniAkEN4ZgNVfz2XJg801SAwOydn3
ZB40SatmasHOCmp4t4DNMQ==
`pragma protect end_protected        
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OMflM87Hn0OKeUKm5nBkDUDBef3o2aPQatFMWNLABdxHREUEsTLg5e/ju8DvsecK
oiJqAuqm+RucbYSKMgJuvBnUdnUgIbZZUP25fLtakg/kiuSVnPI3bjgldagLF02O
6WE9X4I4JBle3OPOXI3fq43RhGah6vcdRgLc0/AKQ2A=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 162964    )
Ijoj1NExmdBWK+bp6RJl2fbx9YZw+jFEXVTiqMic+DAoGGmR7UJKiBUBdAebwFAK
7qpYWq8DBTXDGbPNVJNzXv7EUBl4tsR7zWn/UnyqdBksRC7B6UhBjK/+nYUEoMa0
inB2trt7V59toSBFMXbZ5g87cCQljE5ecMJhSi0CkGUAOHuvixYvrbWpOX3Dai8Z
uVWmuzdK2unOir5PMa5wEH2jNRQgXj5s4TRbADynj8jNoydSOpq8jePHG/sPamh0
rSAZmgi1BOlcvCIF9/wt1ASGOA2kFk4gnE4ef7DdX3TqyMyTvEMr3Pg/z51ylsTD
SdqVQ8QeTKxVEqrbyRCzZBHhPExNdM9bcgpScCFfnBsUPX7JkJxggaO01V6xPHQV
5gVObRdWqVC0ikTwTUA3vCuhucMxdiz9KA4xaU9AOy08QAmcAKLlAz9WMxro3oSc
LzioufGaKwMvQLfdn9tGXdUPY44FSzZS8U+ztR6xFd6DcWZsRTQLsOR7BiMmmEMV
t5r7c+peT2V8UvW85Kfj8oMyLx+OG+3F5Ik9VImLNup73XkWCjgS5HO9Dq5AlqeZ
PmJ7cDz8xGka5fMjbKBPSQ==
`pragma protect end_protected
//vcs_vip_protect      
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
kxfQEhjew4MYseevccQ+nbxw5+cxITa/+9ZEFDGKZD1rx319Iqst4QIag5HCdY2y
tX6NR0OJbf+3YAxpsct4HCUuEcVSgol6vck1uwP2PFLCWE5VACvj2oL2E0af+OCr
1tT7nhZQxLPLo/9GelN/a506sKdZyEr62JIw0rgENWw=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 182406    )
1tRQdHRztPV+srjoVnID+8Bx2lbWf1Q7XzGOMLxL+M7fd5rkciAr1p/+TOYXTGm0
v0Wusa3mEd3q9rW44DhoLrUq3urIIJ+haSFjzJlmi5eNywxArORepMIwQ5wPfzvh
2TXdFAVPe8vlB9FvcwFQ5OqkNZlwKRlzEfZcRv2fuY4ZOIVprI9Hwtp8W50Aonv6
P1YjXIuFTvPyaQHCLkqoCKe3k1ucRRZlxIsSw+T5g9aqYTcIquSDoVN2e2V4sPP1
BTCaUjEt7xwMMhQEe8crH0lKbxvf96GaciF5O20Oa9CzKYHb3odrkM1TYptMjwGJ
wm0g1VZXgtPZgOASboJOT+Oots4d677jom9kGZbjxdhZAJLybRacS4/rLWeoapVK
38JpzYdHJarRPTM40+8F8Vn/bZqHqZzBiGLWPVmEus0w2q3kW1wb/JoESh16Uol8
sfgYOl3hjfT6sdfWLeH4UbhbexEJaOQC/efFNuGepAI+dxLXrnw/K8IxtjtdhzsT
H9jmCkxGxGRtnkUfH/8ua7lJXwYDSwGIgiaB0LT6ZfigfCF+Qg6JCdVJXrJn67OG
BrSDN4E8OuIK8PXAjPz6LFy/R1GAImOzRtMFEesrG+IOX3NR9T3qbWpFxMDEFfkb
qQCEYa10E1uuua3yFv27GJDJu72vbGSgjakKxMqhHxf+CyWaioKdvTVRgzWgCrpa
utHC0DrMQPGwTwKhFk1zi5Q9qhRmiDN/lssUKOfXK5DkdUriJxAL8yfTjMzr/LyS
rTLhK5sYGMaqY5wl1lIlBJ49dWg+nQdl4TVCFJY3Mjz7FVhF7s3ta74D4QlFIXgp
JZApfGBdviG4F2JRl/Lb3lx6Bf4DFV+4zcvD8rleCNBmHr2nJ295gQ5uNNO4p2zn
pnpd+c2DP0cxmane2UPwhR+Av65A7UcUgXLfwYL4EOLPIEpzGXxEHgSTdWMn7wr7
WF5dXo6vRfTyPOx/w6ZzNM1W+ZQrEggmiUYNh4zxhjHna5iYsz5/mUwCr8+P1E1V
bV2k7Uhb7QCsEkBGwFTEP6BGDvUYVfdQH2OfOijAV0aqz/KuuuQPi6cWy/TFXbtQ
s0AEcxDhtmmf1S/iipEnZp1VL+3JXP7ZRgI7AepD1roqiCyOD73LhPgU467gA4FP
SWDkcbIiWFN9dQw2RVjztBh2rmwc0oHsto2pbaAqcHa6/tb+3KZcK3LuXGbG6UO4
vWaXCuWFMYQCJ5JRmkfMCzlDS/2g+3LgnohGBR6Z5xX0w4wj6fDx9yuTCJ0UbUcp
St/MTL2TCr5NGTKucPbAm0peaJT2h3ubDQukS5usKN1i7jgV3u/ydoS8KlcR/pej
2ro6Meo9iI/QF22jxxCCAccXLqZrB6NJo8zxKlgz6o258iTcoi5MHrWyXBCIe9HP
47O5k37ke9coQ79KUHs9VZ0oiadBx0CVtcky8IVyXHvusEsZI4wPCEh5VbTIiPH+
V4fbz+ZSf+J/chVHuKpXvutsmyJ+uhp5fUMZnJlkwTZgiWZoce9VF519PnO+aw6H
JWJlLqb585LQSeLG/Jfo6HMwY6+MiE/lBGflbvbpznJGLMTU5WFwVebQEzErZ8hK
eIBpCz1K2b+Kz6JZCeu3vxazrHM1rAjxv+OF8TfTlb1DNO1zEiysLqus/ckGIJ1Q
VtJKusEq7Je8mdwqqsg4dB+vXc2dz/yh16JwVzmGuFZ7WebQlWSQdxnRwwNuxagd
TaFwsIioQUQuFk0eu7qIqEAe+UaRVsCj+TkyB4WX1QdByUdUF3b4hceLRQYe3aJN
kKiTInhqX6a1sZVPAhpRN1uRGarrJNEaa+n4PteDLpZndnz6bCzGawoYNyVtUbNS
S4P82K+0pFc6XjpA3FvcOSBiMU2EjVZccUT5CfUPBFfxckYEBr0+9cmn69Yy7Huc
EuZ84bdFD05/g0c2C6CmXeRUeTZ5kAZyacquHuHjnPtlp/bsRQYKoy/W24jY0REG
UP5rOxJu3CnAOfq+qMPgj+MUCp3jBuGSB1Rp2J+KTQa4BkeTtG7MIQjs8iabIZZY
j8aqxZzPo1rLw0QNMi0O3eY92Rdw7dMUIr5+IzVGPhhDBvq8GVPPUIM2+NEnya1n
8if5U9ClnB9RPhE3dCWbk+nT/TqKdU1S4PixcWlGkBfPjMcFZeZN44lcxzRgJb0v
AFRBrkVNQzZY8iiQjnS7JV7LpSLl9TYaHIw/X7up+l69LLG9P6jEYolHEgcKKAXy
8BJeRjcktTNVdbeqkQ4j3sFW7DCVy3IJ2bsIAiB0pk/4MIVRrumslZfNNYBrNVvb
+0w7TcdUSrshc5GZq/TRvOCTz7BXTHIdBCxHDdWV7Lu/XJ74/nY8cbtpF0+SFl3R
EvBYaVdApcW453J7dhiziyJZIrZevAweyOujKr5oU3PWZKpugzj1Mu0zSqXcI7Wm
F3gAJb6YtjOtJ8GqorcqjJ/lKNsSAVoBAYyMetQCt0DTzCwBPpRxfTQiZX2kMFU6
OXtcrgX1KBvvnyC7jTraZIUazJEt8UAZ1VnlvUTMsJj5bOh2IHj+EFg078DrMuWJ
QhordAmhWexB4Ts2+31h0pqAeL6zjI7LS0YV2KUXm3N5n2V3GvZdCnaPrMi4d0eM
wig/r3N1WRkoJke/9/lZFoYoFqkvt1wxiAn7FbL+8c6+oah9otgfyCS2wVrZ/Ubu
1Wb/qOOermZ5+5sZgFmIhRzpJWzF3kOWQD3YEjWXXq8C92sAFfN5oFaV3tebqkzu
WsjBOo0QQecobDtBP1Iqt2ZWr7suMbC1RrJZ47jmeer9ib1Ctc9jVfX13NPNa7m0
AM5wtvp7Sy38u18X2nPBPexDF1BPQVkZMevuYjQBle5Oq+ampkTtbwmJz3jhbeAj
2vInMLXqIz52U38AfFPyJCid6E3LLSwY/BxwjEN/uvBeRbG9RmxVvF9xVITO13Vw
BqzN1oyenhBGTjseTcE/8/yd/YxC5mmfWprBpgsUdNXGjexyIkMscCgcf3qFEuj7
5+panKbvjXVfBWnbSO6T95uqzuYlfZIGjUlwAHbTsNL5SJRFYttHnRqAlF9CA69Z
/q1WdPHP2YSLhRBF8HJIUik/aPwcUkqurys9xFE14jGop8YHE6f0M9ft2+Lgc/an
BhrTZbKPktExBYTV5D/811QY13TWiH36EeJSvDcPh7ZlpenYRFbBccEBoZsk764Z
tC+Am+DJx+uelOdEJVLXFx3ScwhqYKbR6p8nSEDAJjo0wuyaK3q0qlnngISIrg4T
6A5En9VeIop3Ud1t/qhaEKyejdEke8nN+DMDtedH6YbuaJpXcfLPAU7zP2XiYGoE
vAZhIuqk/796VO3CXrfWLt7PWcKWAsIQpQAxNApRIarBqQM6RW07aYUB1Nae5Fyr
djmUfwEhny6KeL8VMYN8+DMS8M+B7rxJL0orbum+PFyQEpdW1aXcG25QlUQ619q6
7YD0h5zKJXHjBEtpR6aXpYo1dvQ6mR+9ec+MZpEiPoHkpZar9sffkpSmdZf72Qmf
2ON1SjOo1wiYzzbNNfVjAe9f+5A8JR6ynthsRE365U9fJfLbGWW3t6ZudDulSbnq
tEr586Vee7zzBX5Hh06H7PxY6PJWyHG8uOKMsZdUambmsX62bibwC8iBq45xbSDd
3lAyKsCI5fZ9sy6kKXluU8toe1sOs9WeGiZVSn51Eefu/cBsBBs0XQUMP9oWjQa/
LP4UsLt1Ykk2tNNV2oGBCjIzd4DG0GTRR2jv8DcmCsWE5BX3ASlIN5GxoPmY0r9X
16xNWlcndTbodJgmcPIdeGDq6YMQCHLGQG31rj+Ah0Vcq3HhlJr6otn69n4r81ad
20kCOOV/JnxY+bXzZw/wiWnM9VVDJouVIN9pZq95kOLaGh3omhF0JzZZIzywVomn
6l9IdAT+EMOxJvhOpx4G4j5xRz33Oj/snzoMPJeK4eeO1HfMQAfeL+O7qoE3TDl/
UWUwKNad3Uq17qo8lG2DdTm3Utapa2OMCLxLuc/5ENtS/8qtLKoFOiM6bVM9HVE/
2uc16iOgYcERhmwdBuXg74ZBsBF4Rv9WbLVa0F11z3GGXwchAASCyPrRYnQtyZby
USmJsJp/Wge6i+Umljno8ZJ0eq5dYjzf/KZ45McyzT9pMDIYDxhgQ1dKvdQ53k3j
FwHxlCNCXymifekVj3nBT3Ll5Bi/QvRdoGpVo1WAVn0grLrtMW/JaK8lMik1sBSt
D8wF8DmiExkH8Ki/YM3vEbBxiYHf2bqVh2nW0mUpPOuLpUOmEOhQXwJBpRcPvfHL
LU37AvF4C9W7fwzma2fSgS9IeOtZngMoXuKXon3tjaDVQGCj4ZgBZkC9e+tJrljN
wJq8RjqpUIbaH+dVuZb9dMRiMZQEhT7XpVvbR3v10RcIPj7yB482Thn/YJilR0PZ
It+SzEL5Hsod0RLNHC9xTnB22QwMfskbmv0TeA7YXDkxHxP+7+XuXpGo6AKDzebl
bnNQVVEbsd/qB6ridvIAbPAT5vK/O/H0olM48ZJJAqmprMQcYYA4DlqOnZUpoibB
IccSTHBKF+CEt5q02HPsyWkgmOxqJCOUxftsOi9nDkZi4VUEo2Mllvi+uUjLATpw
TVtZh49xESTfpVV4GpK5UtxkKVQVg28LiVFTmk6K8PwpwGXlUI+XZDl+eoudWlt7
MlcEq17tXb3DzFo0OH3NH2iYvDz7h+BbmN0ShHIPXSYEcf9FxFhS1c/f/KeoBgD5
uxgcxoumLSOT47FAppLqsVKD8J5pN5i4WCUuk/IiXZcIsB780FvcyYZqdYn2Bn5Y
EixCagCbxbwlHgf+vd3ljkQEb1oOIugMh8pwirt83YN+7O2+OfJ6Qm5ozTcmBxgv
oG+AppTDbdyJuaC5buhXu6OZiX/3S7/mTfIydI4MY+rRbyHRapDZdypLgRxRLrpx
09qcLx1rpwYfglBpPBfSAMec7O+fEMPRM2w4yBtEgX0yPEec+IyydjJYgknyhgu5
lpzEPmGL9OhZoq6X3RescB6xx3d4aElmQnal6hVDTCkMQKDFgmoWQTNTKAy8W7JG
9P/I1vLPJj07w/S0TdsjUO3IEvXkZjJyH5M6K6Fe0xkYTsHbMvVCO2HMet8lmRAQ
GT1FvZjfTdRCz8O6dypi2IVojH0SSoHrSqlmc49Euc13O99KMR5kT7ieiUiNwL5K
yX+Ad1johTtNI7jbRbYa6O2U7E9XDjzHxVS5LqiqthqPVhxJfGHVYEfqyvSiRfrY
oiTrY3sbCRc/fJx1NKnyxsXREUdVGntKNBXpVn8U7Q0FYIWcHvMfQowSzG4WmH8g
S4GbIsYxLMu/a78vEvp/HiUrRtedl95m2qZhHpxiQpihwZs/T5N7yG8ObqPKGuGo
ObkKPX25UkhlQhFnuV0S2HEZVeQ8ZmXcfjEJhSwq6vpoOuh8ZGKSB05Jpx/mMJqO
H2U6cmD8SqOsKUFx7sBVjtQ/cvVAjTzLQa9VMh3vgTOCfJshz8JPz3HCySaOHH9G
+ORyqnlv3FVYfQ7Hi0nvw1ENMusHJSbrSRZmd1keApegYvG7MCXWGeasYEAkKTaN
pn43AWfkxlp0sEvwSRyTdm4ypMnUFFcQVtEp4pL5hepKf3r+na+trJN8Q39bL67c
bsPstf3bWXK5GNMpjYwu5SLjlOoFfqA7QwWqpje6zCzYZYQqRKP92TBpyY0pa/bX
03C/tEV57mUt4S06a379tv9enfjcQcpwj1cYqii8l5201KKnThAo8uAq5GW7i4tw
q82jLw7wPsz80dCoLQVrShcBHhOyejoF9KQWJA4Cu6f9mJOW8psgwo2Qf8FTmHHx
hwZSsRtLsFB9sTArnBsuOFCrOu2l/y+SmHiSQjTVjHSe7IMeGpKhbMFESa8E8jkR
JQvbJW6PM43mTQLD/dMOskpu5EDIV4sUncMJMRsQIABgdZuMCjFF29sDl2Be9TcZ
wOI+oBO+ZoDApXMG0NbrfwH2j45idCwrpip7/3E+CadBdHFO+O3cBtDeL/h8wHYe
6fs443yC4PzK3hFc/N5p+XHd0dF1EQEpy3taWIqGCg7cfeEtlQua3Pg8suNpNZAo
GwOImNXnvBbvoIJ0v3tQiTOdywS5FSzJzmMunXzgsMeWhWgZtQn29pY5/QTzHXbE
aMRk3RgQ1FiPaYKkwCTu3oViv3EGmEEMXixMxTum/eZQ6t/HaAFwhZ0O3mR21wUA
pRqFhO8ogSI87FkLOgCvnTmF+Qy8fR0WnwVLcb/8Eun+igVALtwkTrFevMbWzN9Y
pGfIxvGZBHSiUqVHslz5akDlOLlO11iKjVhbKRH9105H/n2KUNdijhxM1tms/Sud
hTiUpQkIjRbPS1fRFBSAxHO33ZQ4K2wolEyp2hTGnpdFeADQHSRjLpFzESHO04Z6
BLufi6RdVlVQ8pd1qf67gVkzAt59dtvaOF3LTwFZ9YBk6Uy3gtpQJAPOCMomV5bO
BYyMxyLG4ldgorTZiOegWIywXNYY9ZTQzthNvorZVDnhBuAdELJHvNgUJFhmX+Ga
UTgYlSlTrgWFa73MrX9qG/0PtHGRIOAPgwxrYQoHWZy/APPT+8QT/fFUrK9VLYm1
Gb6/QDCzjgu5FeHsh4wBZ7f5g1o9Oa2Z9fOujBwy+2IlG9LWfq3QLmXxQMiKCKer
IWdaq+Fjozff7J3XqCL5KyzWbhGQVgZU1KbHApub3x437fwXDPq62eGzzpat3lze
6MGtGfgZCfZIrfGE5BXF4UiqTTqFCQLwcDCUBgNV4gOKIjbCHAnCO2oxMR9LkW4p
x8ZTAOrrVrimBd3PbK+J15zMqz/2auos98figuCCsf5LowN0fKbMO10ZFXt6moSG
jiiHkuyCNW1KhEbJjw4z7AmMw2xy3Upxt3o9vQymU8xiTIGr4duYj2zskdSoDtMD
TydCQAFesI18RERxJRwT3OwH5/tCY2YJNjyIRIhhi56LbvNH32rH9J+8gtTlZP4h
1cdKUDK7o4i6ayZqSmxlxuy2Qqx47Wdg7qF0f6/DVpW1ELT87Hs3KHHJARgW7Vur
/ol7gZMfoWdDShUnC+nk6KlHjvU79f7+NoP+mzVIaoFkLcnUP+vwzZPZR4LfXqzy
dlteiXK4L4bYM1fTr1JxsRKtBBSegfZD/tUaDMgxFWvsDCRU839Rio6ETeFJvxNx
XQ/vkZdXoZVxjlYfF1Gyk/SAmB/k2F4yzVzHzHL6Qv5X2Yoht8ev79jf4s7LDTVT
4+KEKTs3PWadgKSKM5wreod9ngzLfm1qhbKwwe4qoY/Fdp944C3qwM+2FdiRimaT
WGJS6DAmXsJoD1TPCAP9okI+IKQpLMyU0eXm9oYdgbuMubGZIsYNgk1z2KF8PHFL
N/EWTD5B33MtGUj8KxySc0KtCorXEWRT/a0W0oZZk0zRoS3K6IIPHpAAqT3dAp87
pTxWyhMFl+3fx7SYZnYtGX48lT9RA7Plb6zujTNnt0/p5zOBN0GzqSGrj1jiw+dR
+yJqr1fN2qHS8+RKIw0Hy2ojP+abLHWlczVYWJQBKj4Sl4Bz2QADe6KtGOwDMexv
czFi51JHGxhyeMQAq4ymJKucXyqe5+4nYA6BaW7xSYStI3TwYFmaI0Mm0Y4el2YF
uuYGiWSbSLhYwnt3YSsDEwE1ZG8a6g3qm5XbXVAGRurVew9Cb7fQx+WUxirlz6ef
VTrl91ta5eg8sqEinHbWtgHiiNb8KflpnVQpJC6eam8jSi9dCKJ1zKp++f50iQRD
nPUfhTY9kp0qc0/9XUMnYPeAzu7tbyxy7sQuJhZUksouCVlAjD+B8n7VRHoz7Ar+
jNFSIcSHHEQLlRb23PlN9G1Wg2/jdEQD1j7gJtCNxqvla3K3ABCec7Y+qsolBFdY
5gk8xWbBlsMn/R5mQ7w0oWlklIH1/lTJ4S3idiX7LWs+HNv+HdyXc/q79s6rALxZ
Ldw8bVEfwEoYuXEYnN71ddVPDELqKDkglnJaFP40z1NJjQUQJ2fSVEhfZ4rMqzfr
+jNeD/sQoFA9nxc+0gMcdPh1HXkMeJfKTijOVPfZZ4hIE70ajonPUVDCsLmAcufu
TwX2LM0J+4RBJQDmg9EJvgChtw08w9vc+3Sg6GEvoF6d+Be9+ZRT14rpwlLrwdxS
rszuYrO+JXjuCsSGxX3hks2GEFkr6K1guAoi+1tmB7alYXZlJSdiR/5kCO9abaAl
hqIpdY2NCOVZEV3glo9nKKjrFKd1u4KKpebruY3MV/2Rl72kmDDvU8VW9uokNKrZ
uvCYybhMoBoDKU5c1fO0r2/iUZyWoPwlVvZ9bxSgJVTvLvUF43VhZkajHTYkcIpH
5swEt7Qu+ndLPSduBl7ZV3p0mm0iy3wxQ7hE0Zbz9KxrLsdUe17IekqiAcQD91DG
EtVXthPhKCcnYoWa53Me6gunl24xJmlwY4Eoh/CgVh/cACYhi9KSh/3m7Rk0YmUw
soKkn0y4uJ0MkE4s29O+VkxDdSouc1tJbiWbB4aktpT1whTmQxVuEqdhuDKCtFS+
RmxLIGw7IYRtQ5/o9G8VPhZI9zEZao7abGLC0QcN28tYMQelOrX9/f3gXQ8Rh78X
ZrQTRkVwpHBCnWWtXX2NdSBxrQmlGlqqv+2iOJFTbQRsJY1WrRiM9hO97zsD3lFN
W+qzwB3AFd9oploR3MegxPohGd6UgysdLuGm27tR27vewLd/ko18PAxf2zbYDq1s
dyLz43UDxyBDBfIWvxKmjxLjJcbLrCoBv54a5nm7X0uKqaY1RYSqe+j05z8ul/PW
Df8NrQtdNr1+lt+kX4Lm2gouCF2ujq/W7V1hZVG9u903kGw1/HAwqUqK2KucjLZE
6Qp4/1DVMNIOqUC43CJ1Dqw+n3tkZq6nGuwPtuzBbGU2bmYij3wI11uqJYs+SrdR
glxWO5upgCYjN77rfmKMxFY7qiJKkPi29nqMNvVzLzZLgWMOGrumoacv14GKaI6Y
X3TF5CstxYiKzBePHz0vZQJQVLLtZ1MPmlcr6imBbWEpWokRhEu8jqLPFhgK1Skm
1DFYdKlSX2c2pp4k8WeOoqzG1Q4+s8e4dLupvIo3UcPEeKph9Ra35w8q6XWL2FrJ
WCOcq47VMTZhNrsKKK3mwzh1ljFZWz8Cbok9NBg7tTQ7lN9R1BXxO8oaWGnMjX8c
sNTfFIqNIuqpRfSleTuOn1kuwEPzLpXNngt1eHF/lH6gNB1m0b5pFQ1birmT/V8C
e4c5uSF+Gi/gDrlT7dcxVs2lfwdNjjq++EgoL5DlJQXB9Snkv9QoK59G4ZAJ6Z1a
sJvuBYyj1pUG1HPXeALTidS9b19HpNUN9LtQstScBCeY67vgSd5wq0VfHy8kvSqC
TNqyS+hTO+JHrf3/90AbhAnrad+UcLbckK4FVqDGdAUzd3Fj3oT1HtUgdhjpIei/
nxpi6y3FVSNpRILg25Xz12r61V1xgCczY5ACtDv87aWeDA5vFVpmwotA5DxYwjXK
6I5HV5oHVAa6kdSowIJHzRvR09uV7+b7sj8m0WqwExeZgt9QSP48krWu2B9Rddlm
b8t2r65jozUgRPMqnJo8nR6J0mVXbVYmjJJecTESa04/QxbjzBiZGT5ADrmWMQ7w
D8K/wldIaCKBC1/JOXDvMKsRD0lzKfjjHKZsN180pZpJfmHVgJRftuZznYpdEtyY
MTG1VFNDzWWDK91FoEEFAbolMaotpUroEB7IfuZ0rbhtp11PqXE6kmR+MpNFYrAv
v3LOc49BEUWSZF2dDsF/cH1wY20IggL+U2tzq+9UDmGFVXet4rPWTW8niZckkC5V
JD8ImExx5wbLWNKgufsrVOD4+ztTvCDf/74ptCCpz2iF+DNwQu3vylDk7OFeXWM+
sLjuMN7qlpAOr8GVPWuRza5fKeQo4LpaV53So2lZzzJ2NRcIJwbidzIJBXm0hUYI
84iEIjsfw0PV1UWfu95YCJI6CCser3nSwpYtfyshYAaWCHMvHZ9woOySBtSdQut6
7YsMaHhm6XkDbGqj/YYkHieYfy9+m0OBhZdXfFnuWedPuNBdKoWrZXmgWVbX8WSl
BY1gu6964AAIcv/YQFMmB2FD5V7Enk7sKlv6XSWdnZ669AWc2c5nubaD6vOSe8jO
DzV8wvxo2II2oDq5qKpQmN70uBs3ZN7rwI401l8YbVb9LmflrM65ZhPU0W42TSmZ
CfmJfoGEmX9OQQ7EFMLVrp6MuZP+Sv5HhrboTK9qUaYNMv189ccTgoHNul/Msn+Y
Mj2mFgviNYJo2GuzSO2bdk9V+3+jPK3/m9VKShtRU/g4jmFmQkDxEPmzy5TSTkfP
h9GnkmgOEuSIHNlU0tESFU0vo5qgpAzAbkPDZSK9YWuq7bfkfKjcuO56qtLRNo7O
EvBla6sAuR5GnkKF2claOOBsz9s6AvCR8Rn5vid89H6ELKzBpaizYptzagR55X75
dYuuyRFpeiJIOAsLUt45cshStOEXsvgEuQZuchKUnQEXAQerIL5rtvKtvUyF2lnl
4JVaeHpStArwP6Qr5nsOxt08nvYX+5mwKwHuBfQ2kqTl/zR+FbWuFnB88Zsba3l8
N6SkStMFGm1uteszVOhRID/Q9QqFppvfLRdc5wP8vCPu1mLhLV/bt9U7s0BSQn6i
xI8XqQZSr201TiGnb/sZhqAjX2TtXFm+Ykf4jXVLOAtskPERaLAyGbaZ8Uow1K9E
ZjGGUqOKad1Q4O0xw68syzj4hljdUlUrzyiOSVV/z7pqhuKWSFa5exgXzXQ7feVM
QqgOJ7ohuZHzFcF3c5rTsXMq82hNnwMphC9U5B/vXfcDiSq4RZH05d9Vda25xC65
52OHVkZceXer1jQB2SliXOhgQt9llEmsszlpmmyDwUx9iIDIiALjjmEQ08zqf/yv
Fq+6DmH6W70FNtvSnvxPcivVr3c0gkkOt93b7rueaiZGET9sgN4YssVnLCfof82K
L9rda5Wr1wVf1IGyvaASl54mjxhFMMXZDWoHQvvgnqj1Voyto9XRMRFAUeX8o5lW
yf9q0G5k+nx7RWwupzGsMq4wTSkUps3vRuv2I5T74P8LmrhowjXTNEfRRNXREN2b
wJ3g3vdJkz90U40+TMzzeu3FuuEtbR/OSOD7d1A6NJmxW/xrCDa0jcLjl1MPJCap
PBcnHL9myrTonHuZrt45XC+Cz0YNtu3U1owsq6lL8/c6rrQx1W8ygpDLzP8EfjOf
dLnUK8uWRzemh8ZFla7FGtOBaWzvkknFScJIBAv6Ti4saATgXIFg//m12NiUtAYg
PiZSTqzWJeVg5G+qb9q+lpS97LEUbWURfO+2JJxMnIojFkJXBmVTkXiZRhskmsLa
SXihQqVz8g9DbAbVO9pQoWcirAHDmmk0PngvAAVvmworRjL2xZy8EGaxfPyj8kyA
LwXrcraKw/QJef7aclB2Rg79oTVVpy4sLzf4L/abyyt7A3nQ71jzV2SZA7nio5lm
YbBxaB1l+gZg9K9qu0yvfMfN0C7GQ750fNWw1CWSv96xqLrPshdjIvefKnNP97Tz
ltwR2cJ2dFhxHeIfO+4Tks5wiiY3+SDqCPvg8d3uWRYI0CC6iP1OuvdzbZmpOpEX
lMqJKbL0XhOnG2/Pdtq0oWoCrot+3oMzDfRSHZebsfcg+j79tF3EOqq9wCSXd+x1
sPYU6098YvvX4eHTvguyb50D62ZowiORl3TCEQoSlCZgmZzoVD42VoVvLo51ZOHO
B9mk3XuNgaZvE6R5KyIGJN3rQBlwi0jbmhKjIqKFZ611u6fXUZR8InyxdOpU7P4A
auHKIRTTnY9Ya+8biKLS71SVe9Fk4BkUI2MRjqsDxWRmpS/Rq696d4HxzhOWoAmK
RmMbHubXkKSmWQDxm8qPI78WV/B7QTSAnfo7sDJRoofHUv3MdmtU0Ymv6JcZNthB
0GwsMm4FOqYbKJ01eeoSLvr/9SxxY7Ta4nWopfvv2ElwxVmxvMjBH9DZZRi5zY5T
8uqgyyG931VWXMtMOeY+bxd7Dst7//eI7zU/RBQjaTHDuG3gfyCEUybMDt8InYOY
qiiKmrNbAZXn8mMGtUKHaF6SWqpbk6lWbh/DElgHjwjxxNDVfh8BGXflkW71/zmE
fk4eKOzSAm0KRaVb9jHXIGOglrH3kz4L0fuHO/gJR1tx05EcI4OxDz/CLk0DM+nq
a4s0p4UHUtxY7VoY+dfG09y2uqctIogKdTbOkBPEEGmuQEbBRA3gKH1ZATzMt+3S
qx8h2u6QZ1tgWbmuqFz+ChMjO2tERe+ef+uP6tEVPJOWSRmvde0PZExXXb7e2+JP
4OSGbA2P2fMUwtXSDNGDioj8AnFbSO8EVrdkAK8ByvM7heMGtnJHBgYUG3McFIpc
9k9oDEGkhoOg3vOByNNXuhcVXYu7Fa3jk7HOkzq3eBnUumz6fc3AOsWBJ55KFud/
vya8v+HsDJuwQ+GGn808We87TQEqHuCGWSP9mGdM8aotDHftnQJ4I+EgRhIj/CZX
I9FMRJ4YFtm/p8Cht2qfghMgGZ+cNv6KmtViIXWX1XFf8yiFGVSl9/71ngc1EzJ5
D6gTzGJ8UH2kL3uaheLLxoKpxzFVXTO5tIyqOiLBJVh0a16PFQtWZ3cf2W3Cnk2F
C5IjmtDnk8iAux6U3BJPE7mcXmBhSfws5mbgYEEOmoaut1il1sCeZBeEdMhPmgwc
wHBLU/Qihbpk2pqkwo3ynWvbbFXM2iFjt9ZKSh59snaGOIDKyEZT/5vejYGUzsCF
9/LgQiTWDC2e3F79pr+FHovwqRCsS3Avhfi68rULpmML6RFbP+BmnaALp37zpdPu
I3cg5qc7bkEQkMwH0LaJwmJpyZbqiaRoVHYQhafa3QPEGs2tKLPzYJmeztZ8Nrbr
pDbOIjaO/iiQ4FcB9xJzTirojMZPjDTSmZShFHF7vfU1mOTzmPE1KsmaK/0MYg4v
JLEL4mbX4+Q6N7Ts1Bh/G5Va/ZQ5lQSzm+YQa2nUiklXsyvgNf0WvluNl6lzEE8n
BJYBxJXDncx+DOa5xXEL/SmdtCrmvbVLEmIzY4gCxmc7Tbzrbn2rexRDA4Xaktt9
+FpG6yQst2igVZHrOTASBD9usATywLFEzSCAW6tmWYBUHa3Xv6EssRSOLwACMNqG
3ADwlbY6RpSXFGthIy1h/E0VahVtoK3ey7XQgJh+EF4J4YHqoI/2nmE6YW+fvHEr
16X7d4HqqkRMZinu3PP4gf4ofB95Q3DkZkCOhR2w/sFKP404Znq0+4V4JkaWtlvN
N8HvEaZU91wBYosTflzsgppMdOdYHIWlrfemAitYtFoQZ/yXzPgNCaa0SoP4dzso
2LiJbk/SSbfOEkZFVcoEw4BtNaQstyfbzBrwhd5ra5Ha0hVXjXOzesenR8ymqocy
7uML8rFDAASfneU7bgFnzY6pW+NXUoytHaSNm94/luQk9Sy4i6b4JmLky77+UMvj
qz2Qog+w25zfxyICyhM68OR3K1+aZ0v5/3FIuX60/NauNgNe2lC3G84kbGqU7gXS
VGBEVRtV+eEDIEigozgU4SjRBrh0s0wxzhT1PhCwyZvuZcdKprA6xXcuDvt4Hp2o
WwjO0LNWrP3FJp8VmQ8K8FERnYj1BEIVVaTnPbZngjJwWMXx4DCjjqV6eODDSc6z
Ny2xnxjvWq13dpnKsa6dJO+mm0IW3QFRiF2P9ueYr6EjDE/O+tNOh00kvZd0xtPW
C4rFmyUHWs5bl86CwPIAm51w6ocOrQm0c//hk8tZ2vleHicZ29XsBTH01hu4XYn8
R/6jBzUxyar3cOGKvP17p4BucX3J668BaftUM9ChoS3EGZ5uTJxBPPRWXf3t0M14
HsjD0supSkXtpOjLrY+nevV0uoa7qMYNWcZwcF2WO1vEd/LV0aU9DTjE1yEa0CkN
lhGleLO2xt9XDZ6q7QB5g07rZWqsT8F9C7/roYr5xVbWFu5kAEMrh/mwD+pX0AXw
0JtN05BfLLqZzvYHuPDZu6LyqsBqXdlkT5dWq1tTwOvHHGgK6i29OvdSQgr4JMIu
9BmfUOJcCUTfrh8508UtAHfppvO77VRwft9EHRWqApit/R+5vON7HfNFsViMHFS4
W+jodP7OVXdsLTH69g3AHjwEVO8xWR1M2o7T925ZqMrmcWeK/Bct85rly/OFjygE
e2gBRbI84FlxNgPrY3Tl4iElZwyAMSHn/d9jynx4s6mvxqC6J072JR0SAdAS5N7g
0sybLG14iZ+h944zRIDoSLcRyiLUxX0M7c/WCB+LVxRyrDAZB3Sw6eTbKlvlaNXZ
Msyk5TAjR86mmLPTJF2gNalY5Ys1r4yuUlGaqZ1HWAnVJu5Q79Cb/YXdTZwMx4r2
Sf/GzISytDfOgIc4UVNg4GO2pGzBKn7YrInLxyIs0kmWlSFEPd9b9v7bstPIPFdV
Ktlnjxc+mBLWBRpHV9c/NrJGErDfhj25EfnAQBFkcaXSP5rMj8tNn60SLET1B96x
xQ0P89F3/hGIe/SBfvKwcdlOmVRW72uHk1BuCy9j0xvt6S/PWdm/kzjIoAw2scZK
MV8r7/BU14RmxQWMPXCjaxrdwgLqIV2pWjFPRf9LYkYVb++tueHq+5Olcdx67hy9
CJfUiiiwA4SMzu9GDpBi2yCkR5Y9yYk5TiaF8rK+w6JVkI6P8DzIqZTfdj6Q4YJH
zL1Cx3Ml6zI1VR60j5f29+LVBaMQcn8ggxS5OFJ+NmmLjdZBjX5ttNUpOCZ/uq3P
Bq9o9OXIxSCgWryxbLJEjG3l2QiLGfhh/owOHtamvbTISOEW21pcmTJFcuXG/6Ot
H/FWR9m873dVvYPKIUpie0LPwJGcOsLdKC6Y2XTRpl0dBiSIYWJQ1GZL9Ev7Q+M3
XcucCsJOz0ieSCwEjW96pam0A0UfrZ/HJ1oJoxImf61QxC/ewe9CRxIhhaYUwyO+
BoHtcHxBZlANvxmAshOb6besramWyDHYzvJUW/xxjoF9iYmWfJQZlLgtINOzPvTJ
dFnp+nXRakyC9GRTiFKuJQI+yqwf93C+FMbkcwBy1FcbPPAMz4zpf8DXMdPae/I3
8pjbijzmIOTgG7H0lDuIsf7JLR8Fr9cXzXgJT6WJH6fKdi8qhe/45nNNWTtnzAZc
txmysXVFsdFifo5x8wfbM7rmvintoLul93QsXCz8ggJPFS7l9qBQGQZzQWQJ6I0D
fzlNCQlrXC0A5iuI6c8SR49IuF7XtMXO7NjlHP6K+NAu5cRrD9xtkOLazZFlT90y
kGgGW6L/RjM67G7SR43hP7hBtpuYrfZa6aI2iyO2aKZK0UhL6qf7xF2KBw2R81MN
39fWh/YMNQxD+6milnhhxXqMF5KI3B2X/wr9NBCzS7HYSK9GRvoKldCk5ilLMZHi
Ri2aI5SmQvDiwnMqZdMfdDZu8+T0XTa3ycANTIojtaM9hJ8sArLRzwNd6iHeBFM8
iz3n9kQ8JNGOHxYndrveO7jK3xELn4RU5gzRh9lsTCxxO4XrdVpd41UaDyJ5cmBr
oDQZEslSlgYW79w97YsRbJe8TyC+LhqvCCihRwYzYHl607OmZOfqGdsIlCIkmmCp
SxH+rOZk6ECE72lOHrD0Bs5k8skNM8lCSjjc3GUWbIl9RYNMeKJ9KtXtd8GAokJF
MNQxbZYYEBXlnGbkQgSpoRbq4cujbMAOvzFs+qNH3WN80kmeq04YtXrhcE7AxABv
E/R0M6dMWo3/9YfqdPsmVffpsUJSLTmKXQq9QyRORR46ltUWf95DA+ls9He0D9/r
py3fWIAspS3mb04ZbiazPPLbRSAJwFN3fjLrVO/EyrMi4/+rWL1Int4+HZJcTdPb
O0+zzzyOK7qENVaA5gDJl6ntBCaufllB5Chv0w6+yjJg/Nt124+dP7CiG3iLnBAI
U4E7YY1z6Vmh8f2axtvDc9I/yAWnhMH7Ss4WE5vkS/b7VKrDyhw9TjFnAny8PDDi
guvxxVsBByvGHO1LUhYLvZyuCbbKGY00G7A1rSel7m4VUIPlNDLo70o5ClqgD9uM
t+oa475/1ZrlJaIWzHxWJRXbv+Z1Qhb1Zm/3+OxHW/XU5uP9uqIWE7OjHikQSKas
eVvm5D0YYWOflCIgks3Vbdfv0i1JC8n3ukcnKk1yIAkPkhB6AGUHSxslV/GZLTv+
s5bhbwDeVFOiG5u19EL78ubCMYjTx+SzWi7LxEwvOLhHyNW0IlLWIreSbPO8+img
G22QXGS1camHkrtpmhCxPaX9nRpcNMiDIrqlcTOapN7VWp+ivL1sma9+U1WWqYGA
g/jBhElIMVePTVhjbg0td3Cy7dIu50tweoAsn/yyXZ00tMdmZv1WcbMeWPV6QEu+
TSHid4gURRoVIVuVbo41+IvenVn8zEMANmyi+st12qwpAv1uge+HbOCdTtS4DxE1
TtiqtQ2UixShAkmrTyvJmxnnUqhnV/NKqSa9JIdn9+Jftoji83rRTOCC022ipyFg
rOg8wW3AiVpb8schLR8cb4AJZGRO7185GAge5c7VXTMzUZafXOP/qNM1bfPYoDLM
FEPtOz9bMzOrKFJWIpLvOFN6vRTtcgtEXDlJKLMlwtDQaz3ErXqlYbb2jlABOx+p
rwgbywYB6TLW4BtL5/ytdtQPVtmjhF55MVaWdK5HDb8dW0agm8nvhSrrYSxVsnoH
Hhr101Dn5OhBki/fJiGkqXCFV3/v1T5Kt0BgVa/pb29I+bbTRanyi3awagtPBkEx
NS3+yKLndxNilFjv0uT9fZNA1uzkrlcR23CmcACtcBv8/+sCsi8JJ8GQUS2/dfpK
fe8gsworZrzyIuXTQToRg2+mCNZ+MY6CIbfoE3FHCtUGe+wNFq+QWvnvzx+TGnDu
BEoFE7PJrdbvNVbNome0TqdltN4ZUmFnZrO0MIoHU+e5m4f/4R4uuy8YQLTQ6/F/
qv29z5AytS/Gv3iveA/9F4WWUEio0t3vacorWzJKxHuXojHCh4nJjq642J0KaQZZ
VcJREAaLAVMAdKW3kpL8Ei3gvzozgd5mvMUroj4bpHiVm0zzlFIhs8hIglXqWZSl
vdGSGJsuJf8giXo87mh0r8zduVCSuDvELiYPNvJLQLYJ48bgLZI8r4yPNTCtyxH/
xsuduj82x6K+ITTuz766aAVd9tpcU6vGxYP/HO2Wmr1LsCOsZMrK+R3I/sGqUV/4
dEIXBFcDs0EcuTT6G+syTPb/NEGksHDrQffNhult3M4sYeJU7VMLuqXlSDSX8xUV
FVMdpBIF8NMH4q2u6TjvlvtqT/uADlQUIpwZh4o1fQ19Mp43LozvTVQHJQxklfUZ
ydH2j/+/rz2PK9Xjdo/568omPyQ1nIGABXjlCU22L76+B5Ebug5+JjRsb8t0SWxI
cbd0HrKdwUdMEPtDwEnB/DmrWjLGMsB8lin1iTgFA8qYKDBHLT0v4D1whgdD/ay9
TS8ra0l3334+yy/edkK7ZQZs43G+8NLQt/Txusak+9C7/ZlslLWJnfTZ+Qd5UZZO
cIPfDlLAMf0n6c0ueWeLgzv+QcnXC2eO9wfyj3SsHEHf4HWEUEyFuzpEkoRStEmq
xF1UnAXt1YOgfeVIUTz5omPHV+aSHRn0vIaCGQo8829f4/0NneIlELNpyY7VzUZ9
ms0lcZR6gSl3d7tyC+IhDVinfoCzW7snwTiBrerfL9J8qgX11s1O9BNYfiRKZ1aV
lusNyPP+o9We4VqhwTHYsXBxVTKgWehB81gyWU/TaPXxrtnuy2PTsrcCe38wNGeE
Mg/zRVFWZN+mMTzvHpTWEVgCzgeno8nPwtz17X3c9Gh0yh6rwuS74mmJlhcdFe+x
ZEVLfonBSHWV8KKQZ65ihq19ef9HRDnmO4OTqA7z4825cpZhRqy6OItbKIZv3SQM
JqHIaFq5+VjJCph9Q9gR6N4ZN8eUlHnH2PFwPHxKkFMWqjO10kbS6ZAd8jF9LDV4
m8Zjo/kzgFfqS7pRv7xjO9+kUA3YttDp1a7+BhJ19crei9dPNCe15TdZFkkOehAo
F/2T96a6fhsPyzmrpD0gUq2DZie+vGbqRRo+nQgnDKTgSjCZCX89EofgChFFM6dk
8ChBKELScczx3gX9tKOVM6eN51XB8AtP3Cih6L12tX1gcuKMTpSDhyLp6p6Mcprq
sjchMdjrP/HNzUT8s5qo/0DiyqJcgsOz1FKEtKVMxZefu7gmcR4BGrMR5h5qpW+I
gaWbf/HEvSxtf03v50YBo1IELkjXbK1wDR96/+SALqiNz9NAy3C1RN8xQYU6RM6V
6JIesOph9GEl7W/hIlvuU4W7UUuKej1nUTWZ976XeN9ZM54s4X/Y2rcYt/YhTmFq
+KTw5pK7RytQ97eqIri2uPoVnysEwffWnNAzID2nTsWDAyPJtgIAX8ZV54pffRjd
RYUNERpvr6OK0+P9tmTJQPKi0gFHAfGaY/B5dqLXnSUPEzfi1lqUlgq5+Ainwlnt
mmBfBsFijZqYafPFLMYzmjupWcTE74Id3DCkGdIn/konGF3CbuMI4KG5JvTPaE2C
V4jXLkABD/sfCZY5abuzUnTY9MAXPFDiOWlHhNHFYJfP40gwcT90W5+M5+kub0AF
rd2HW/SDKJ8pSM7E6G6o00DdaZwZC9m6ELs+dSZcCLXqkwWt2c/ZCc7KNDPgT5tW
0735oQ/+ssJ0HasCmwRF72dooIc/zOqJ007tbsipy9lHsYwnHnceHPqwpLaWYN4e
R7QsgNrFCb6wsPByq6WuimSOWYQOMCfj0SUn+XZJBmMEIpOIIqKHWMxdVNkWpZHi
YJ1cUf1z6W9QhUiT0ttQfhcoJ9jLonpcq1AmgyChIqB0dE08sqOjSyMwRvrmBAIx
3IBoZq2PtjZ79ggx+KD8vjCEqYxHTAorfZuKoeaFF0VVDErjf612n7w5nJVW7Mzj
2/6ckvNzxyokRY2T74ZrORwgymGWzKYbcTYgzGgAYmaQS+2kW+VxBdxPVltD/DFC
4JxmL7FU3bRXGd4jqhDlomojEvPkg0EHPF2730lq8L0YC1KnCrZdIZNDXBRmyTzX
4Zl5f/FE1Il+8KWUSATpP9gb6qK/Qh8xtxZGdlscoBCYp8obciFFPPk/KBeE5/OQ
wGx3aBcjR+0eTSG6gnPqwhs73HwahfLclIX4upNqueXXCQ10F7Ely7yX4joKvlQp
nt2geCw/NVRUBF48YPM337HuAZe+9rC+U8POmBHdgkTd5wRd2NI7oK9xHC9G9EYc
i8P2uveQc08QNIYkagjLZKQHWCmL4tNWunxXN4892p0I81mmvMiL005Sjh/4qXco
FsIfCiRRbi1xw1i/1d1iix/ANXhI7Pjc13zKJuGhidum4xVC78cfuaCTbqhBal7K
xeQ3/3UZp3Z/gS0OxjhxZH9rTKbdURZ1wBYiWrseFfYCyoP8yNyfLtdtsrfvgevD
Aymmm+nnrXc3ghTtIjDV7hhaFsJIxWrGTsoc/h6c1nCbqQyDEop3A+xx9GbnTsRJ
RcbvjTIPMRts1hObvxqRdcrMOjzUuDolYpKZNfwKmDYE/71bMJ3cDdMipRlGOUYo
3HfDXpWxUjRvWGDjlnIIfJHjcsNa6ENJd6UNDLz19Otl3zX0k5UPpmh2WHMWRhOB
4SEUOmHSmdbgkWiDVckG4NuHY53Mrmuaz1vWeDRVeAo6Jwq+GLUennAX069V2QcB
2xq8IT1zU5zrA9KRYHCUNkHwKCrD/e7g4UcQdpoIHwzgYtRZLm1j27CbDl3ValzO
OSxiNsR70Vm2T+OLTafh/6a/aR49mpsCAWS7AE6BAPRP33CnLKcHkAyWLhl/7hmV
c9epLIHUjdnCZCGHxCesv7P0Sjq5pYbSuW8a7qGqe/x5JONHNpsqlRypxxQa9RvZ
EyH6IW5V95iAD9XzBNWNKmK4TTKDh+dBkF/1g8E+Jn9HINIVvm196JiRIzg08yfo
fo1dQH7H9s36tgWMDtUBw3DNtGFt9Zn8lJl22iwGWgPdpuT6Cm1xjVMY8NoDJszr
FLgP7h3shBuiaJCxZ2/3/h2p/geU6MXJx+UPUxiYj7PapJkDf7HQ01/asmX5H2BW
XlzHllo32mrUUxc1/rUbraVRKq79N29ka5B2hQFx42sCrRdUvUzB7xV8J2ykYjeA
LDkJr6VMtRpaTEldyHyFuLd/E7X/B0DfKuh/XwNlezPnDsIx0o1cVih43bcLqjwX
vfVeF/nvsh13+j97ij3+36FxPFrDRGmmLw2JkUKbM3/VC2OcVMuO5pBLEnQ2wTuD
ifEtGEcM5MHOE63fP+JIbYZFlbqZqZ3OZ6BlbjoEpKT1hY3YmZyHuaR++vQlhXz3
TUBmOx86H5i9KPEqIAnq7Mk1Slh08zDODzSWQ8f1YTF+JL9TqRh7YFiYHdyDdgpD
/CxRJxkJNe/cCo/Vx1vC0L5bNr9XgCnubRHkZN+PmYXo0EA5Hy7/T4M92y04igAk
SlULE9FDdHMmjmg11uPxiW7y08wQzlpK4mA5vBBhDviHSyA7E4nZUYc94ramozlg
sSIfrajulO/UGhaqDo6tBm9hqWUd/iVpKdfiJKeU8rKEZMbyX02+wWSShV0/QQGr
DBf4Io4OQI1bxegnwhPM0H6ca2AyiZitjLaNR847Is59WnkmKZJETwcb/bK4Oj63
5REw2d1wL1UKDH4i49dEA+rdxpTadoIJiMWzA36QSQvSQ/y6ZHaUHkyHZRpn6akP
Xzq+ichchKMixw0YoP2Hdq5aI06Hy1/7xSGKmAs+TW2akwDCxsveN/Y//o0m6F9L
2p17FKJ4M72EtG0bOQtDhx3+33WTbl1wL09Kn0mVUAhjOk6wdeSu4p4x/JpQChUB
nJHCjbDYh+igOaAoE4mmZXzsvY+Z468o1vVnWzP2r+Mmi0C/F/ZjJ/QJenngOAD/
hrItEhQJoi6LMoYT/TSLXnXm04jxMirREOA5/wFoNvT515YM2Nt5HNOk8cP045or
vyHg2FR5fG7G9sOea+qoXykd84KNMA7pt6Y7xvskHl+fYka9eyUJSXYrBVtvL3mn
xWG4QRAySZhC/k1s/PXWy++Ma6WdVXoaj4NMi6euW2ekD9/8+UvvYAX6wypOHtnM
AjKerXcB/tsxju3N7kAQNlYrp4TBsfqR/wCBed4eaJUJ7sk+Zkg/R++3+sMhVpOX
knyERTrkX4/LDoP6uRxzVOGSde1qcNNkNWusIr/ssouhUuT8RJwj7aKyd7FPT/5I
NrRPf8NCprKxAzFtrVIMbAx+v6P6TwuM8R6ZmFCE+9PT5TFzIHbjYpoUGc65d114
9s61kPI31elk6HTXr2GtO1hlGNPfDt8P8QRc6CDnM5DMGW3K31N1E4qyzXcHw/JK
olxXU6bz5OVSj3S+RJS1sC1iB45PTZhRWI5JmyEgeeZGAUN8R20XLaKQva2c7B0W
FEvM1mPn+JLXaqvlN2kW/JBlkvyOXHWS8PCvlNBxBWXCpmU9U8ZZPXcP0NISW8xI
lDI14JcGe0senDaBaOVnzVVtBR/53NKpSD9kG0m4KNTOlFbgzQw5CUbRNMoTseqT
V0VJcLefR0zGR2Q+uDRdqjikqL8p4Yp74qSgbCZ43vP//fbxQVB2kTm84J1+wUMg
PzvW4r7r6p/a0p55Frc6Hgubhh7IuSp1re42Y8AcbX/s+XfLan6zY36Ibzbe6e8h
JRJUj/oS7Odn4LdQc8S5vetJMG7jwPvebNZT5WVCMgteaRFgJT5iPba0hoBrHOrw
C31y8gSFcUlG2rRX6j4VnBWA/40XANUxfE6dP4lEYm0o3RylhbdR9gAsJxUh3/Gu
g5nUXehyXraXeqX0TweVxWqzdQqFhCnDHS/sVVHZx6J5nFbNQHAl5KIFFRrH96sk
G0ld9k/Rir4DDcBbFyaoxUNNRcpsP0UkcRux/KGksqqdgesQkDcY7iZUg5U0kIGF
k7d7ATQ/5Ut2tESnYWxsKFVo1ZTsJwQlHzXHMd+mP9mgWOWzCyahD3LIOkIlPwFK
IwgxOM93fpsCNrBFOKq77gyD1xXVKo/zuQON1T9klhTzT5/+0tg6KP/HJ3hqvrmH
O1uhuqM2SLD+lNF4CpJ8MtTeG/3qwtUldupvBdoK/IE1TpIt2eU2K+xOcFhR1/ak
cGrKSfivbbLsFlhECzVHaiSlAn8NMjEjfv8ewSQ+wjvCGuihnCYsMWdgQ4cVCYgp
bwT0hpMHhebT2fm3/A7lQl8VXRBCXNR2iugkV+dm53WasiURY8XUZ5cOE6zSgXKy
4y0MwnNyWm6skpKo5EgIOVHwEme7GAWdMd3W0wuVP6DU/ZVLcSpKLs08b81zsNrG
b3LAaigu1j2r0akc/eWdqY5tCS2DqaeqWJNpBmqdR0kSdsJvY6G/wYpnp4RU0tyk
fCVoJDSnuUqLxepqLvnFCDX/5yBNPJg/OuoMolLKG7FYQ1310J2B97pdXnQxZz6K
Rr7LnSuflwq86DQKbMyfJUj32JLGUAF5+5+s2bmQh0fUfXaMwOsJ4/F/EDP4cLxz
8XiMh5Xqub+BEVDmSZukCuAuRvsNRxTzFnsqh+TWSUxunPiO7gHeT35kTqy3f9xz
CS3DbNwq5d1+ULIwNzLCHbwJpWpKj3PV5rK6S8gzjS/gtfajzD2DWY1esnni2oj2
onOTMoASB1KrvYJRGRbIFQJg4eM9y7iOCEjUQZMhXn0Z3puFNk4eismUgCWlv+6v
M2X03etMfF+LqlljbEADg3LpkcsJ1ChdxWvHvHaCggh62V3OJmEY8dGfm3zhpiF0
3CVbvwf4kT2ldAy4fRCRY6VOXt8Io4mUvdstxaZnMxGCfyyaNSx7OCRapoRHGOhj
q3+VPzLYwgXE1CLjlGvmFrRlf6fro0Ti0A/5xJsvqGyYOqpluDE/gkLXsvHpPNHh
JQBMA0BrFgDNstF9l/88CoowvCPFmuck6iII0srd0ryhFxv91Jz+m5X2aKulBnjP
TJqRHCi7tcAxLUElQMir/wmknELgqqA8AjtyzNkfhJBhAQf81hwLSYLcIc8DI3It
r1/yCWR22mmqik4Wxkd72FhN68e0j08KF8b5AMlzh8HsZScsriyWWEEptMjL9lJp
S2M2J3LKWvasRrgJE9bbYf5cJ/7Rm9eiaPnRqv+/nansYrmWUzAYS6MymsQYk1mT
tOF1M8LhqfqPAqdld3CerxWsUPRNCX+zE8GgdDWrKyK1yEUV+p0Ov7aMlSjPK+8r
ZAs7p9mWUljtBaWirKun9ijZVymCP12ZlsY1inHiXrSA1fSHTDeMvKIGrTBgnQ/b
HPLshxosqPpAc74AWsUhP/lmXd6/Xq+i0yuAUX7h9nH0Ys5Xdi4bIUeu4QdGsO9s
PZO/nDYjDayfAwpiC5ljc5xX9xdf9iLw7yHJBgsOMPTr1rhvS9ABRtx5hDC5df3q
/6Gj+33v6/V9pGrXzRtvP/J5Aekuf6ml7+SL6pVuB1xGWmWl+AVz8JxEGGgq3Ys/
8rV860sCyUlz4Xs1thukvgjMlIYou3Y9A1zptClQ+i9x6VBArLHPSMcgYMSPpIuU
n7SJnjzN5ZijZ3kZL5SrSkEVzZcguqG+opMunrBhvysstk2UhVktomPMI4M9pxKs
vumevxEFO+u8+lukaLVT6kYszWbBpuInzDHe96JECff4NDjZsbuW2L8vEU0FCuJz
zssZANcLl8+474HMYfk5bwKGbXk3n7OE190kJQj0Zmt7bTatzM13y58Jriv+S5DC
Rj9RyK5xXIuz+a1MrzowDmAVVarm4Dhcy7UHrphqFyR+0yQ/m+8+18MH7WCZAZhS
hmwBQk+vR3glbQUtCEnWFLd8warFM4G3gd/1vRYAVmJP/NlE29ngdSWTCMIW82Mh
4fLEsnMpHKkkAB1fGel7wJQxA5+dQyjeJPsUM7NAHy4eKINyTeuDcp/s32GBlVL7
lMi6x3G9zEchuOta3paJJx8ocWtiMaYVvrHRkUqCFiWJ3kxSvOEQd6rE/EptW2VS
v2o5y8GVkrToH8yyIU6GFDs27h6FPTfD83G7GXqb632rkxfveVLjHsigrV4zkZb/
2k0MPnoCnLGldqQV8nVFW72tjhv3M2W0CF/Rlgj93Y8RP+sQj1Us3Zn5yJO3JC9k
XrVP+EBvue9pBeiAWFOpPuNNbkMvfTzfTPGzKvcspskeRu45DvZDx14UsuZApi5E
xK+fhEd2gIW8NqDnmS9T8CzZ1VT3ugmNBWyrmCa6K4DDosvkQ7xB4Uor2c8d3uJy
uA4bJaNQgKbXGis8woQJAWl6QX2n+qWuCSyKb9PdmOf7gWbaTnWpZHW/R+UfMn/D
w71E9cEJX24YjUkI7qBHBuiILe0JqLOpUADcdloWZ4fExtYIZigSgmz6D6dr1uiO
5swGjmOIWq//rBnpgOR9bB8MoWn1QT8FG8bSjsOOTo66W1E1lYHcrEooX8a7U+LW
G0uQlZD0t8OSPIp2v5oIECWSF0KB5y/3jO1kcyF+xmSdzwrK1WwCqmqORWS4G4ls
VUJVnYeB2oZBJIkXj7HgV1V8lPZn7igtV8GDJoCdkD73O0T8kwIEk2C8FYH+73ek
9h+JmO+lRWO3Nbpj0SIHSQIV5S9Fhnecd6RNwvrCVAC1N+TQd4vdpmznzpwvj+os
75scDrIDUe3eJiytNRXfVS2rZzW0x0ny3fe9G/PhcnevxvCZKYCS0sbnYleFOFoK
QMKHVaFFwm6N8RODPfEHEy70sS6NjwBOtr/h1FgzGiAVfFZfRuiOWtGsI2us7ZYl
BXmFFVHGj4nzmTWeq4HuTHXeNq8r/wMq/VQ59F1T9XLIpXEMBuOufV58RptsLnI7
D196xnR8BzrBCtZznv/aiUiI8svrUkoLnhZ7ZX7CmYOYPczTZFELclguC86B425n
K7eaN+Vt9qo6xEY1rRD+C1pNMHXCMui8p5nEjLJPbRortbWyNVXliw4k5ax4qsT7
K8Wo+q5P/zb/EVpEO3aCqb0w3wul6JgKgV88SKm7V5PYej0ScgwjMYG9n9BEHmo5
nKg/SNTe5+oanpUKoOyO0dj1ivaufkzo5kSXe76sV11+K/tSVHdlyX4QdKOPhSpB
d/F+nMCHyDkFgOPMPsvZfDAvIJgXYdC6Div9qDr3iz9VHkR4E/VAI7Rn+RN8S2d0
NE0bPiE2QUkK4G4fCxteWTLXDG/ZPJDuqE0p6AvvqC2sOWxicd5aV4Xi2mtSTZoJ
NOLCy0T/0kAONIIqbAXcXAPC7/SQ3HQQKyIyRE3fFR2F/xdQ0VyG7mQcDqtolUMC
1ZK47stIcH3vYcYWOPOqSMPmMKCziBp1t6BwOv/I5FSSxVisYmhvPN91oIYraOVl
4yxZ3FVQ2OXy0rQGEyS1hIg869wGzmBwahphW5Fxoti+pmVd2rImZ0GXso6ixxHG
CnbBMaDTQGKu9C33Xutk7bW5N9M5rHVMV5FAQYKSc+S+LJ/hnuOKQHMCiBvoV4+C
7WIJMRNIWeL/wrBvVhgHH2o8HsRkH0cDEBTdvLnmyeH9UoBvf6+4apL/tCyOzJu9
APtYR2yM4Yq/eVi8JaXZShRHQSkwl8sgNaKca86C+uu7ATxCEekSk+b7RJybqU+z
myvJRnRo89LGdhT2BihmfzrQlL7NkA1R0q8T3tL40dQ9ByM2K5/P4FW+zVIBzwLI
C1y5D5cEORNOWV9pUl4aTyFFxeYW0w8Uiu5N83TD9gwE5brCVT34G8hDknC8hyo3
PqXOnmBPJRRJCK+KBm+SicDmZtEeC5PFkehhlcveZL4Tbc64kmeNZl11xI6vNbW6
gufQd/mXKBUG+qNStzgvo4dSnSC/wTpQCLJIVJHzAigsuKOfT5yMZouXo8LEMJjC
ph+6qyPYH5tZcY0c1SmlWBRfGqeUB9JgSSZ77hXz6roNEXEEgrKgG4Wf8sh8eDpo
Bj5VnTBkiHldAQ2xbcBeRKMh4N0uNSGQubzvpTVMEQwHHKdbGHLCUIL0OMKWQlSo
Ij6oRCu4UTgL2Anlth7pcw==
`pragma protect end_protected      

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
CDqhuvWHeQkDjeWbepXIp7gjEmZWBF7NAfn4fAaGPX2BdqwGuRwiIvbqf0zGVONt
zzsZmPIuc12tDXEIOYxc/xToXWQGhk14qN3kLzzm7UUmr4TyDF+ZWzVdWSjAbeLJ
vPEJNeASJzL5Y2FDrrqG5DUf5YgBXlDNPTMgHRCOx6c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 182991    )
61L1KJ+WUXgZQASTN3o9s1HNdzXCZDf+JDTpoF5h45GbMTtarqaxWTu7OAjOP66k
Rrb/wGB1SxNSsk9vqJhnalMXXuRunNKo7ooGnD3bvNZk4GEqQFT3DljMnOVeCkIF
18poVuDCSVa2g+JtXBiM6Yxdsnwvro6xFEFWK3RURHGmbjGfz3fAG3zh06s3rTUg
RX1TDDojCCSmlT+u96GwtC+P0kox+dUSUo22+6ecnO+fm2M8Lnpz0oUoYnXyxAST
99yMUFy+XxhrfnCFBBdTLEoZ2dBASQTJRdq3y3fvKgcjhka35r+WqyhGMG4cLSH1
6RoSRkkCqI+qGnOd5WET0/6FdUi8klveC452RhckLr6j2h4d0N1Yd0Jm1j8tEsl/
x4yQLfg4/+G5v3kovzH/oHQvlTJsbzVOoo8EBraTBefhvX+juLyDPkk/+KStb+Uo
KGkLR3mSHsCb/t+tACq/o9qH6avHsWjjPk/U1BH4nXY4g16YDJTJSWJ4ytR4mUzL
vRHgldr/OIpLNksk2IjIu/h3NFWR2h6E8kKyMCjIGQtJL2WQDhaqHFgqwjc3s4Iv
YG9nZglM8KFXEGQB/l78JR+WauL5Pq6+OSlabf4rbnGgD/irEXdP/NaXPIwY1NMu
m6Iq+XvlYiDvbAaXdCnnm2oYb6Ey+M1WRxc4wpQwtTNagfpEfrUxT8OizJH12poY
Ie4p0VSUhNhwd1IYkxASSXmB/jCn7E6TKGd0eIPRZ8ix/oQTencbzosCMulUJSuS
ww0o4oOUmX3SITDMqhrnqQ==
`pragma protect end_protected
//vcs_vip_protect      
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
JbryXRcVTsPcu6pKTZdZaaohqVtz+6yJ3jTjtcbCwJZBwn2PNiZ9ZGESG/Ch06ZJ
8ZAAVPgGk45dX+D3QVQWBnsmeNFNjGhj2hqc9iKDHQadWu79razP49RL5ZJw2nkW
F2IDZGku207kVVcJn+7EuNJxfH6mpFwCDMwO7gqbcvI=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 183663    )
iRHgLEDd06gFOlF6x0pSOdLTPWc8pF52xXhG16uYJQNH9lruGXeaJesICxw6JhA9
Mo43FQsiURWat7c57QpCpnL8iaelklVEFdiz4MHmNs8LFyAHELGdHm99EClLWxXN
ioNef58IZia7v6imvwm9xKehiLHuPf7r5PBSfEoCKzrj9zbtFyxFI2dusuTzyhqf
nRDVS/1zjOkYWkvD++0dyaehcYj/4SHs7RsR5Qfpry60VJXclSU5rfQ450br/vWa
ZKZVx4h7DSSFLjlPzPO29ybZ7+GmCPaJ53QgBeY2SrAsVoadrFh8A9FP841+GFVx
dqIwKgYQO4hu9j9L9puM5fz6TziJBEnfUsn45QxbjLIJv2GOlm56UyOizR8IVNhX
YXqA+xlSYyv9nYvHejsp0tddK9YcHbNcrtOI6ojNVNephhb+U1HEcKQgxCsQsxbr
47nBZbN5ehVJcC0OoqOHvL3UBRvIOwnytAV3dmGH4qj6r02qeJfLl2ehc2HrA+Fe
7y1km5fwnVvFLKe61L54ILxDUvx0gO1Te7LIXBLbnyevzxbzZIu0A89DjRz0jBPT
NNaZ6zUPWej04OBo0b+ypdCQcpKAX819nl6HpCpXRGMeH9EJz8MKN0by8mHMO/qC
18CwDABq48YQ3S5vHcKH87USv2wKoFjE/PtE/HFzmRPMwev6flCD2GmThMrtAw8c
dnaa1rO+cP4C0dgrF/eznpIcMblRFW4gE3TO8pgB+a9IFzuJlvNECk3jocxC8XXW
H5mOGAKyREaxY1SGYBu0tlhVLt5AcdZe/aFhR8LLcbdwO1Lh5V4OA1uI+YLDYCPa
P10rR3NFP5/X251q/eNHCnVIo809NDFpUKoiR1DQ5+ePvUDV3ue1DaP5VOQLf0JW
/AuGYqPNtprVUSoOrGDFSQ==
`pragma protect end_protected      

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nr8fzOEmbN7c9waW99eTsVHVhZn1g6MCaNgAEfLJd4/jGKFqd/jfBTKp4KW15BiO
C1fWvtoDIBHHQ+VMc9G1UDZL0O7h9Unfz8EXUlRJYADczulTPWT1W5C44RvTdkYd
BLOpumhetGv2ZMltP0h0wmgbNfFpkUVBS40P7bYV5a0=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 184253    )
ShVQTl36chB7ix2uEc5yfPRdbjBzVwnlyKX+GNHOfb/sCMY4EEaKIZUtfy71VkOL
bpJiVFBaArwWvOZvdgryRO3KVUhMyRyohnUYcvwZLvuNEgCMmyOLrwLM7owNTBzn
mTN1rfLg7O4hfJB4N0LyaMLaNRvcUgny8Y/cIyMmLSORKVQp0pZB2ybuuZ+Zgpn6
ISwKwkX5nRMZIKo8UDa//7E8A9QIsSwqwHZjv9pAg1ZumQ41UWMoJVy2ukVyQwyJ
rsj3eFZHHRLoJqS2FCSW6pD4EFvBBVbxAXZ+pwXuUt69HSreLnr8nBbnp1cgHAVT
BPzo3HawLzzRgubJxMcY4Ze7Spt1G2AxJzEwPt3R5uPtgcziNOH/nmd+RrRRBlK2
VjvKImekG+2mEsFsUK+x96Vy8N7bzw20AOGUbG/pVPysQMQvUT0Qcr6ik+5lM2Ja
zqzJTj2Y3qkJf//MlBRi2H4Krt8shzHbrVDz/NQmeLQUGPLeL7+1JCWU7OEswQq1
G0ZbPxoMQ4UTxKEC2713Ktgf/P1fXHxpyU6HLZBw4tltCOsrltC087mEYcU/u3kS
Q9vSoHNNJos7Nv3ficvazcFLktx8OTjpe7/reumTCPrmtwcYyjus4y1nXO11Nox9
uq25+RhDZ4/rMtQLbEJAlicrZi429D0o30KkcAli5JmsnjIIUBtAgQZER49lE6cK
JiU/PtupBuzP5PEGBn7ZLHku3p9PcOmYI+2kLyHM8xi5/eXoJdThEF/hSvBSZk5E
sKSkkugnAjjS/+2KIPgeYw==
`pragma protect end_protected

//vcs_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
DNLxhVykrE6ZZ00Gb4radx2vLJNN07uMN/ojdwovy31ZvQm9vAxE3ENijMKjyJI8
dGY7tkmWb9y4gW9v2GoflItvJNKbbr1v9rdpbBvLbPYqRBwV7mGfCA4v7lsyyCQj
RoGpY14IsuzTtjKGiDuAk40xmF1WmNclzYnr/0Hi+lE=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 224424    )
XHPR/6ovXbRdY1SOUGA9RMbs+OSVFY10TSjUujsjzwMFihCFPVt9vE3oIQXIwM/4
tWBw6zFWIqB15y0TG+d0Wb7GILu/+fzwFa8vZrpsUlGcDe3u6IiqxI1Y6TtAkbqM
b984On3niciyYHrAt67dYLriA+tiDu/Vt6tCpSjPek1iBc06bnGkN/1cltSKDwAB
QISP79IYWOZzmBHr9aIZYtKiFk7hZ0X3ZFRbXw+qYAHkZ1CPOjhN3o8cc/zeoeYX
hNSfFN0eowK/wBoYUUJVZHnjeBODHoPTasFBCsy5J5PUPsM3K40pEOJUoMxNkW0D
7f4FcdxjpxUE4BE6GmJias32sLymDmwR7z2TzKenLB+xmwjzbsj940cWvauGE8Yi
5yrEgxkRjkmjVWBAOPXj8d3VEXvGyg0odcodlP3vChJ+nDQ/a0vo/Woddb6olC47
r+pDcHabjo0VfNR9eJ9ZNHyHIDYS5LYW+mr5f7hzAAq38payqei+VkqfAdEKJulZ
llxuYvN5izaqnrSgW6lMNiHM6BsjFQxqb8fIN6DHtIqrcMC6IstN4+Nf3rs4/I8M
rACSr34OgNGKbICIBDqPUsJxySY0pP/xLvu40ZshuL+5C5YgBckT0FteLGbUbIba
gxlkj95hrmMM6Dfld9ACiYB0s5KB09shtHDB+qujESmT3UCo3XxXiP2ZJdcxPdes
ygOYmJYDzafo40sa2uKZuWjnZkVOaKpwn8we0f3VcFplqQkaX1+Fs3X6cJISwQv5
QW9d42+5Km4WJsrWdQswhihIUXobUmwCd3/3mK0nYO4b39N3Mc6bIvmruC2bK5O5
nMCUQdtxESrla5bmKoA6uh7/aJxIWic36aeKlTXxlS1gEJ9+wosmhvm/n2gTszeg
i5jp3iUodE7eZtxFnzxQHIWh1EYkScqvXPs9taGwAJOccS1f71i1RPt+V7EERJ5y
UIul4wLWxP2Vr0cwf66g4nchP9W6gAKmOsOSmi02fABsg4sOuYYOzdf4kw5liJ1R
59OzGDl8Ppt3cuvEyiabkhyo7tyCBuR64frB8i6K1fhS4KEtW6WH6DH5EwY0NkuE
W3wnvLvp0Wr6LkpRBXnKj03HRbnOa0lc9C1TMUruF1qdofERlep0tGqx5+RfKXRZ
kak91q+JQDgaG6ONivsbxhNXYXmAtupQWgDn4txgXtjK6QCNvMqs6TvVhMLNRVn7
19+yP4vEq1Ehedufy8Tvhl+fUx5iLXArvZXq7tT4ZMy2ch0Lpr+8uN7l7kSoKRRp
iYnqbLT1Zsxj4Am681S3l4w3p33lXiz1CvaX/vNHnFUcgHin/T+ppvF3QEf9YkdY
ZKJYq5+p9B9svn0hPDnN4edPACIHw/09UeKXiCJImAM15iyIHYGy4BDEW28xfCCn
B754vZot4A0oDbTaN+y/vYV9AD23OaG59V1x983ykqXb4SYoTw7b8pW1MVvXNxE6
e0FjJv4QubQB990C5IdRTvWtx103Wudu21oHvj5yfCkqroO2F6ATyISN6NFgAJH0
vjlGFBewAFvpvIrej3iQQ1OV7N0X286jXwtifa+mJvq5r9zpQq4d27w9/WGLfSOp
u1OzpHP6yqKZ9ltab9d0ISWREhMovCnaeCjnJWgUd/wr1uEn/u6a8zJAyuoJeAM9
RereduZkOIU/OR194joU9aSlnjjxVZcO3Boq7CXmPaibzeT+q4TdhS+tXUJhq9c5
dNLTOI6hCDhtNEJiyAVh9ke7EEygf+V58ATAVb/5q4lkmtlG15UW+0FT8Jqh81f2
AbeYCvcGAdP6lA1xLCXbc7ElxSMPLBg/Xw59grURoLNtT8JdzxLusvBgTaCMPzl5
iMhb5YhU1Q3aPVx3yo826La7KXH96iJBF8GCHbm4jwqO3rQeGxH0gTGrc7zR0+hR
d+fjuBokTPZMAi+U7CTCArug9OlO2xiNPaOF9DftxH4LEZ8LNRVKbXnKx5EcNX3G
Y5b+AxGG0yL23SbvC3RMUA3qr9Egwn2FP0J/Gf1wTaP3n0RpmTeCoDEImEmzgFKO
5yCCjUqRCQe/owS15xBleqVgjcjDiLHoBPuC5N9gUkAZV8MxZQIjpvv5vvu5fXIZ
/wla9zVgDzYe0DWLRxVtR99A8RjVhEK8Kj1K/KG4FCDHGx85+2uBQ/VtV+uw2Irw
Ul/Uyt9HoL56GTiUGzN5Urj2UcbZMzWGGxcheyFfNJMPdOAM1xcW99bmIq/ocUut
srgohEToCd8NAcpj7TYsPjZ57vsEAoBe6/Tv5r9nWU5TkZuVvIs3hIHSkJd/aMiH
5g8wClGAZqrmtmYaSKeWfgp9fFDbJg0O+WeOuZQasiBT6NlvnGnRUooEky7AZIim
FnCaz/k8sxmZRbU2WoLT6oOUxQaf2ZTnRfRWmeX7vU6Fh0gHQgRTLR7VftxBsMpN
TEIXXX+RB7ItnE0ett0ZOangW5/MsqxY0yF2SseCLJ87Jo8VY2DLoY+RTuMRQO/A
4Ajc/5xtd/vBny6rfjnPmm9RaZYFHA33dH7nWgNPUDaYb5qX1JXsT4UQX07yjLVO
ktPK8b+myPVLhcykgmIjYmpn1hS1KsFPgg4AQ6XpWW71O8t34tfJmn6gXkCeZmWO
JTc6gF10LBtiMXi9w6gMRnlAfIPcFHldQQ8Zl5rpZsxFQ1N0tYbmEeaMoa3TRoSW
b2ISBEZsBwwJaFrugM/1QejeVv+yaU7refYRQp2HCnbcN03XHftd0lyADWCzgT7v
+VT2M7ZacmNvMrgSED8V5O60PDwzPPyskP/Y8p7VVRobWO8J0hwDRIvqtWv4kCI0
yzMkijvV/UvR5GKVcrG6Am3/sCTU3jrRAwDCM6LgSsrIBlAenSVEu3Id1nhbxs53
euoE/D6svVXroe+EtreDYdhPJw6Qo609dPU0sBZ9ryBaOImRjwAVSB+frLfgVIND
VXSXJwW2eibSmNg2P4u/02kMBhvVCakpW6YjmwkmuerW3SEYOJ65ddKR6vbq/l16
sVqiydHdeKc92E6GtMlQJop0QGK+X6n31NPsytYM/pF00H9jzl2n7/rQ7O4z0Obh
DqD/P6xHBp20/t2qeBwhpo0mkGKBZ9IO36Hfo4J9DBgwQpYRfuMTcTZdq7GcoIye
lqfvOf09yTC0DywmJAVoCym6jAtwQhTA0m6i1I7Z/Db6TTZuvT9SwUytFEMupolj
DT2XM8me3CM8S+CnUcf1V+AXvNd8H/9hvBAsZe6VyOpdrZ6Tky8/oxaPNpexOh62
4MfzmLN1R6GUlIg/JH2fW/ZG0BE0mPGlC3iKIsVbt56Zc58QrJO7aWjcAWxHuXFo
u6GAWJX0SqWhDCNnrG7M+WfvSfXgcPHwWUchiuAOhlXYDpqoNEIeYRrZrv273SDp
OJuKkN+Yzjy8O0YHYth+6X2U1LN6WHaTa+HeV56WAgH2B4xwtQvBxI5ywTbbsZI5
R5BjK1vYOz2drZnetwbasMH587DCt0GYzW3NAPrtFu2r8+w18kDxCrrFfoxWxiHn
G1fhWLxAXg6Bycws4S0eD7TDRB5J+QSzr69xdQBgonsOtLatTVwqMFN8ozg5KvfJ
DGYWSokcbR5cm9FxBNMkvkyNNiRMSY+/KlGoQbcMzJyXHs5Rs6bT++JUgBEdexsB
9JTYN28G8ybi7bzG600GYVeSUTHihc2rLUDLoziZcgzdc6y0+3jB/RRBZOuTfj8n
FrI4Uc/cENr0z0IU8UxWwREcjfpbZey7AyDV7HVdt43Tq7RM+NW2KQ6TA9x1JHmO
J1yfzHRKxZKrvrMqSAXef/bp58H8rgov8GmmhFs9zUk0AR6YhJgYpWayGmniISvt
tbyzFsMvvQF/NOlb3fG+uowZosOgXBAmAb0ODdA1gRGZ/jjImlehDxV/Re0SLZnb
g1nHyYiJo2r/VgPMfp9yw3ZY9H7P49zaFB9uGG72w2WCUXwq2yiC3mOFDHyed3g/
5DOGxSWOpyWrz0X7OmzYR83D81DSGpmwx2fMfZXIn6+xU4ypy7P5cKHQzdE9trYL
jLe7hNiwRN6gFW0lXHCDY+orIMPPDZMUSwN5Ag9EKR9e8n+Jz7fWKSHOdgH6Hikg
Xr+4Y0vvVKpT+Tmkyr/Dp4X6qATPWMWlCrZHV0k22sKoVeDuzuiRP7KgoBRFyt3D
nCT5jujQos9TGY1NQRT7Yh0bAuYzdu9Ew+bvs84Yu9z32NdYq9fLTDsOAwNShkuL
/de1YJkyiI+KYO28jeCT8JRu32X2F1op3EKNyfTjgTwKL56i3m4u8unMintNZ5I4
L983uALrexbpvE3l63uxUYh7JYiZtmET0xjY/in47+b8I8cVhKYa4iuuTrzKFEQo
9CHtBY0lCuawnV3T9WT5xHxZOLRpukF+ABYjERjMVrgMMQ2LPvL6qSp8oBT2wgLx
wj3XQmSJTKAGrEmxjnJKDNd5f8t3JPWR0uInFpaFa+cQTXm3KmSKkn50htxBNLRd
rrlY9Bs+ZAVxodP6HEO2PzGPZtbhQgsEWeIK3arjB2r1blnCjOtUKfWrlb4A1lSB
M8Zyk5Ne8kYyCewmcTEexcqgp5nnxhp6UvrWhCN0FKJq8cei5otPAXXsEXzUIdt7
/LkANyuo8dzBveewBAUH9vIdrY5fnIAB/bDyXzV+bLJwDkGeSIKSKACXph79gjE0
l0JCAdvUQhZKWtRtLrbjczuy0IDhxMfkuEnrBRuDU/9mEb679663H7UUsIKLH47t
g88cRUEtsyVWMAuVNq8ijCV2nYwzGu/6sIZfG/rfoYX83MiAy1D1eYJznswfmNiA
VSjfz4FpW0ODCbQmLcVS7YUhMyjgbNFmxtfHMOc3PRNeEXsg/E9g3QbJxQtJwqN/
g/gX4ePglsmjT7ibWWpPJmmy2ZXGg4tU6MxfNRIaP/eiN5XasUrW94pG/WDQBT34
ceag8DcoJB0kFsSua79jhTvFWq6fbhRRhsQRQ6CBM+OKeDQVX9mt6bUwRPs3Ib5H
ecnMcye+Ez/a5fUB0a8MbXbSUyoh/7VjdADUArXQn/+g35pQnPva2gMaBwg7MLQ9
upzZtWtsJnCsfCvaFNMqVhfRGGazyhC/6fd7eZNiWCukb/CoIumbZCLmyMddx5d5
UCYtYhWZv/WpivEAE8uhkvcMLb80L7ilkLGMZ59FTFBHjUlufvjRHe/bj1rTXgCM
O1wZPzi+bR1lPtVe82CfJPNNmDpcXf2/nFQCKPvHNY6ZCbDo6gPfcQ98iibHtVeR
eiDK0rgbThdX7pls9c8t2+fdo6JF+16Z0dXQm6mSwhFy4p9IfB/dw76MV1cOGnWM
tZJ3o74QWcMB0EO1GPQsIlkaWvfAAfAkemwty7I+tMtMK9GTG6E7U+VEeB3BIbIm
VvYeMjDAbIFnU3uncMDMHFbLZ5jZDRq5SRur+GY1PVCAx0w9irYdJk7m05+By+jm
RqXILhHvEAm8DD2RN8PTE1tYsrHMPxci+IzLZtFYoDag761W8s0kb5tOyr9VFUqX
4v7CfStRD/qljLYdWFNC4nCVn9dN1FdZqfUFwqLwqrzXA8KRn/3cc+/nUgThawqv
XqyfBbuxODI/SwEc/xpb5sZd/MZl2UXXY73tU+D13RpYVW3ysbFIVJOVQwLb39cB
AfdAL9NEuAhnT78ASwQDRWrGC9xG+jWdBdAJ1tR7DDSsFU9ASp7SmJhxq3bMEwQI
GREs9tkWoMAEos2viN7+Lb+NXZfmhPyRxRSrjR8id+4jtcjrrGSIKTrRSzrUHYFg
N2mr1Y2f05hRCCLPOnTbvJ3GkCvrcp/Hq9759jBpbvXzxWOpX1jWYFKr/jK1TU6p
I/rBA2uioa1OQtToFdmu8SJ7bS3olfEWg84Bxhcgk6wLlr5uT1sQUkUxWz59/+do
7z3rjbOOQ8ka5j/IZdDB2sh4LI+G0VrNs9MOMYatdQE4n6XyXZjkD5tHihPXHpwT
51jZWq+O4s5diGZMICzAyRHTpuBPTaJk6tNaZG7xaHdhL6XBHwdIZMdY12paMEPP
K5bhOZIKqMLGQN6sEYmh1SEp4ZCP6miIA9KbwGTCtQhasZlpohWgvgZuA3ORNQUD
Gk2rf8h040Txjx7AjeVgycvyoF87nSqmASppsxginY053bait0VlPqVIIYjlC/wi
QjK5u/7mCMJ4IqiO6eyFItzE0WEY7sVoYdpV82ndipd0d2tHiPJr+t8pUHt6P55i
1a5n1Z/ad20AXH8p4CX4RF6F5Helg+tgp1wv31qW9c3UNak5VGWDiFo2A1dXKI+h
hUrTCgPu7zSkuiE6FjLMRE54rlnNmW6weXm0R4TmZrQJlOpOnA6DlbTSIfa4PFEG
vmEm+uwAMZzgvuegRIPzaGlI9i3acW8T+lNkVbpmjNhFFdsTLA9b3CtpedicYVlt
nhSd/Subj6Z/YeqZ+UOKAGpa44zG9BY78XTDUFpqD4eC8rseKm7FLqT9kPmRVIzL
LRep3RCVqINXG0rFu99nq+Ds5m0tKd0yKXq+SfGWpy33lkzLuxCVMVRh2+XvLivI
mi8dAcbxAl65Zq1fb3+tjHp5+E0jhOwaF485Xe3XFeeSX6a2MNLAC47frBKeLZHO
LT9VtF8im+bTrnoWeezX1xk/QZAt9HJhXGRGjjo1hxzQlDdpJa+T5UQW8ZGOU9Y9
LLZZ8tc4GjTMCby6PROpmPMEW3aasd+KQHMb/Ft6dIWRfyjEnW6iHgrLz0tA7MO9
gSfMmVIRBtSqLDfAwBaoc30bpHlKxxmy8TeWBbHPlgyJWxJj5AKChtxVFeMUFYGw
E6tWlW66qJu1v6qSC98T/SecDh82tr2zhaidFG+aP9jGlVQA2lGbBg2N8WXY5142
gDQZWXufx2hezHvqXm1r1F/nRmO5lDNmkhpz/R2N6YnD/Y3XeYGtrpDBz2RDo0cW
hrz36td5LFysxC2wBI+bFAPrGTnienqnAQTfROoaxz60uMICiGQDq4u0g/5YL9PU
GSONw7+92bRxkd/ytxNqIwTJgmeOZDGD5PXCCKUyNg9Y+oHCb+KeoY61vH2ya9Q+
7t32ucaD5ILtiy0mwLVkKnwwElFq/TD2L6+PpJBifefgK8+TwFWUwJNOL5vImGdo
TVHvQ/fRH/4MnNxig1VtJShbY/44DJ6Yuh3TEZU1uNg7xGWnoMaKQeSMMqVRBrr/
7Mq1g5GbdqfJeiTYayIVG4QX7Erm7cmcJTSbR5P+fYtyMBiimkd6KZMEavexfcFI
qSdpQjqGBFFIa5mwIXcczyiRJy5bf1bMIt3UJb42AONbN73CsUPOgQBNZAMPn8R3
b9glHhOSVekFwmbWA6fVWZSTdGPovsliUCBEdrgrLG4i6bwh3wA340k1pNBwrbrN
0QfdISir8L3Uc3Ovc4s44NfyIT9an6Ohwql6ZH1ZrHxRSv/u3NP1OE9tn585BEH2
oVOptn/JPz9bkT60WuLMNkhsiYkHAp8C/iwSvllALmpGg6ibKehkl6o64mwrc7oK
nm1oARLhMvnQcbVs+CUcMw33nsPDhCcq0BJnKi3WOWAc5ReKbpsQeIhtZVXW2/hZ
krZj9E9ajir2AQ1UqioCACSaEkfnVpxf1xWEI5iPmIC+/5Ev39MzWBuZWTWkzbMM
LxrM+bqaEcOiqKM5C/6NSpvwLVrFZMJ3Sg50P/YnnfqTleVyuzDwS3c7MUYUM88N
tFja7oBaRFHdNhDXaF/QvgScltL5ecviXP5gfgrtMWpm/9Qg+/Xs1ZruFMoSM7fT
gPyd6DkMyYCriNzm9ji7LAHcOGMdWUts4imUlllePrc5dKUVULHHnIUYfDuxn1jW
ghnfOeWLUCxchuheXQFTnSWviapSF4Oy+zCIaXpyIir9WLGf5WdCa7GePU5fYN0f
7fLtfqGh1+Lz0oSP/dQJTI0MUNKavd4JWC5XH6Pun/NxbTGe2QWMS0qOx9ODCxp7
sNqiTpBiIGtgKSh7zNOXRLRdjulQhxDrK1U8dY/aLa5C1S6KVE/Khp83ewq92/eE
4CJym/HxuBic8ZB2S8xxSfQWzl091rb9nrCezpKglxFgsJNE/zhWCOUwAm09CYuP
NwHM8v+nUPzQbzP/JZqsEIjP2ug2S62Ts/sDWO8fRU+EO7Ar+OWEj6KglSrVbm+i
BnCTOcZVCvXxSOJfhOq1OPAToOqV343lzdErIqtwAPteoo0nUdCBXwE7RbV67/9m
tsaM+RLbxMG+Su0/GoPn8g72T84WQHDByoqodAUUO6yHQBqdYEqFXBRrRTx+J+Ia
SxMokyqmW9ZvNRU/dA31Iq+uFCphc4njZc2ofcDJWRyUQiyR9ozv/w8P1yC3PAj+
6V3k+KZCbFUStCV1ajU6zxqLbY8fg1T8Au2OmwQ23UYKAqxc5um8sytMysZJxIPw
EhsDfVi0Me7p7vsKnW03xKvgl4cZxw1nUPMCmZ05ks28kHEtcgw4Y9Y4weAL+wAC
T1IU04xyoj1kbiR+Tti8te3Zf99iYLttwPetNa/WTILj3zRkhoNeY2p1WYhsEDHr
d8/53azvJUZ6tMM2ojRX4j+wveJ4TLUd6hIAMUMW/kjh2r+v7Li8YWY0ZAAKm6Mr
QZABHIgZniPtDRFtrg8GUTKWqa358Km+SrQAiRsFhqsh6WIybQyl2utrTSz6Eajt
GQ+vffJVNI1wVD7hvkESToz+NBvSi6lWOsz8Ct7k6r76Vz10/ik1a8tuIBGtr0po
0XHLbqJDZFKvqWFXgeNYQMtr4MAImzzOf37G4oAH6dX+o4qR5TUgiKGj2ZRZuznh
v71KofNVHPnAB6TUJKvhM2ODn92gXyiDkRoRdw+z61ukd7B6II61c6HfNQar4j+N
8rusJbfOJun/xEucb+gTJoW5qLa67bZdutqo6V+UeyIbN4NgmTSkCh1mqbPGSTWM
ULzn1ESwEeaihwBHVg+RXczw/KXmQcpF9Nb4cpf0CXmJFpZFpyjXP30/3L4EZxYU
Cko8dMtf2/29HsPCWHGGKqqldipc0dKxkXyXi2sU6Fhe/L5zaPO3gVv6G1IkjLLH
yBc8tMPfnucpfVKg5+lhQyYOLFHahJPfPqxtyekLW6w3+fRVuWx8jGvQPUni0m3b
6AAZ5Mi5baPIkAgFMOOkf9TCW1YkmZIbuaWGNJmR4fIYG/ollfFSIV6HFUO6deK7
YX5YAoSYgL7V//LUTzeSXImZVx7dZ9a/utqDXhnzT37bUNyBQmYSEl62crZJEAxE
cbEuuJcYlg/zVdbRSlCk08LIH+J+GjNqJ9/jejfncxp+GcJDmqBtD1F9WVjbKhrf
aBR80aCyOaZ8HZkKkebZVIeixFFqwZQec6b88c+qqSxVWp4V2ZKJAVtxUYdUsIQg
ER9sZkS/YqlBaovWpWAjP1Cu0l4isoFlLzAdeZsYzAuQ62lBsTTc8ghkPhvPVwMS
xjXApUy9eUy6aQo3Q37PefoNTRRlGkhtl2m09LCR2yI88VnQ7r9QzQRT1WDGeEFK
chXzpVJ4pkhZlNuY6vg4IcNel2ZTQTCZs5+XW4a9sk9NEqaAYdVvDGFA2Em93jwT
fKutktYIz2VZxh7rcf40Vlsa31yNvp7MqMYHu4LLNVt7CA52gUKVFYT8OPs6iHL8
QYeAkTkPF8it6xCyd7IzlRYf/6GPpIhN+O8SyyYQQxbvns45msepthe3JthCm7lO
kqalu/vH0wQVTGqR4i3ZO691dxMWqywYby71iq70Fmu2I/r7vDzKxW9cfFjwQOgz
4t0HVBC+tfIR7GItUVWY6yjOqy1J4el9Tygj5YPZHjmPxyKBYPTsnN42L4CJ5GCm
fvktW2GQrUTjv/WSXpxEEGQbtqDhal0P6q4ooerDSbOxa6Ibe2gH0PaqqBiJU1EY
PPa7R0BmN5jB9jK7TA6l7B5m7oUfelEjJVLflHTiAujXwL4BIBY1a6BmUHPtTsMH
2eRMYRSJ4R9zliEspVJOi7MF6BBCej9FbiXXufsL7ksdwE5ecKWRqv65GyNdv7Nn
3AfPYGU/z8MBtI1PEAGE6i+no3PhHLQ3cTRA3dg29ejNP07QmRknVL5jIePqmN4m
8gmSsV3xWNYxbjrjy964wt9q9Q0QOxusSnoSC4dAm2nGkA6MM7FxzINjA5Yg6rT+
lYCec5mI8I3JyVVgQzZRqw/aPnWCkTkloEAtTmNtnmGzA3jsZZKKw9TeDh6XmCOq
Xja0EJUz3ZWxF3h55pD9nzH0UtfJ9UbSEdze4aYkqJrsBqI6DAcGhJOZhsz5/d3T
xQPft6KY3Gca2m8ex2JlzSdiPMidVf4EHuIaaQ804sINFy31jlk1mNf61yEqQQq1
/xwY//9sZqBVWiq/Pv4MoKGnIPgpM4Xm94QBWnHyAulNvp/uLOqXJKpD4u8wRv2l
wGcE36jNQqwKYqRJQoZplEwkV6McM18hJNScAdxBpJHcmdVFE2nWV4oSc4E8L96o
BgG4zOMjgJsK+wKnkh6Q0yCQxU7FfZI5Ak25buoCUGXzC6aYA8ONmricyecOWqJA
5g/hppXH7mZQEARjbSSbzKJ1aPoH4eWJpWrvSAAfoLMHA5fkT6zRiip45VGTiONn
svAPXpAbC6rXPqL+ByTSnswbUjehhQgojywui0vIUegKuvMYD3d9Z35Rat9DSdpl
ovxxTs9ZFBkEo7p0aV9y49a2R7J7jJhVOQ6PeFSbSG+vtjvqXFmCPgsNDa+U7L/q
gF3resjPSR8vENNgvqQt19K8dKME4mlcwZBYLHH06VjLBTPBpL77OP+C4KBB8pP+
wS8AMzEgu1ZcmzklJo9BXj0z3qa6LZMxH0sgMlnQ9zeO9TkN5oSFRkAtDXk1x0tw
szELwfm1eT4TbzbOU9EfWEPr2Kg6+P2zx1ym+x2kXS7dz3/ySdW0ZIzLNEjnMo7F
5i7/Vjz8puZhvl3tmcDYstCbbgoc5brFWI7DeuYxDTYy0MbMimREaqXprhu61pPj
d9O9k4iCx8g93bdu1ZCDJ3gPppu0/H9UUp8PLbqRf822S5lNzj5zOxsFjCOTklZP
3bt30lcf4K5QCEyQbsk/0Xq/aRLH4cUUuzZfLVikQq8+bveyHzGwr5Mw6ZXOAybR
YZaTDfP/8+O+rfI+Iu1qJl4s/xLP7CcUGAP9Ye3w/sauKHZNES8OnHgute5Cdyjy
avYHo0NqWiq5L1v4Kj3OBPJh56ECNSUgdDnT8fcOC97OrchknwUkzyvlhyEUU77B
T9i6MpIKvFiuF/9Sow+n9UOOvL+b9tMmastymFZSeSfaFyRkM+am4+IpANFy0h0W
wGFzt2rrVuveooWYTwqmE8j8uv5q3cnG4ZipeP+DXvBUrSnwEg+JyuRD05ydHwPu
NDNN/7H5D3e++2vlFnEorIPJcPmEUuiRBWBwSJsdAMN279gmmVqjMrz88oHJdStc
qjwK3V1UMgYHzwXFq7jSeVqXxLaBWPR753N4fTfPKBAbnf5S9q7H+HXWh/WpdUKK
dVNAWaKfFBnUaJqqh0aLQDlfftYqxTrfPfm2XhVQGQlGKTo2Bp4K1wvm5SR6NB2a
sh8QSHeqtWYA0mqS1gw0YsTHSOoVZ+rRvdjbO0apZ9VhNYQQ7h3KSotX1E6bGpKt
aXWTR95xRRIRwVnGwY2728IoO9srcZE9o7ClCxUzyT0tTE44xvUCdtmAwhCmG5iv
7cjnz+z1Dop2QVpVlo5Z2PZ1TcI9x4QyzuIFmdKaIuZBAioLjjA7ASF+w0WvDGiH
auySgPoWR+OePT30Drgl+vPPXyCnthkzYmFAiYtx2I9aUCqXRvqEpEDyYMzqH8LP
DLXaTMYKBqMma1eypldaMtJdKEWrm0xQ3JMiLQln4A8aq9QCvGKTLrzc/8GM0a9w
mWFf5btIH2MqimjNVxAekDossUtLuvNhJ9woGN9apjFP5rN6x4x8EfwCd/1Lj9D6
uVbqep9RQDif4NENxrQCsnHwRycmXbT5b70kC520GREgXg9QnHLHZWhbPMijNTxq
dMsXo8tnZWGDGdhW+lt5NMAw7lU3p1oVi6q7tHgP3SUfJbthGEDTTrHOdvwynYP7
Dd8FnEBZIRANORlp/MY/qBsvnVFKLsT3G3S3P9QF4X1hn7UMlerILbJcIlyhXbgn
I8Bp9m6ZwhOYfQeft5e5KmCj4BaciNLhAcEzPuEQxUyIGaNqquv9Js6ZH3VVial+
YQj7NkiX4z6dSLToEvKUgzKDc/aD0i5qE/3IiLhoXDlfGyDrlpay20JgpuxdCXmI
UTtO1CqB0KpEAIhTIzIaGYPp78T0ONeB8UnVCBOpN/ZjVF1IJv/HOnanmSr3AKPx
vNQOuv8pjwfqmnPhswdPgmRumfixgLrrYQP/eruoOQDCgnIRKRfmT7hyjGCpX/78
WjErxcszKikSRwnFrZCAqShHG6obZhA5hRrztJUVABfwKwMoI3fIVaeDST38EBs+
99QmP8H4/FPpoB+58BmPwRsQDGsp5U2eauepV3kK2/IO17pP8gz0swinml3hbWjn
iXzavIvVrzCpfVoI3jlrC9+DpnenBlrNEE0IxtQduZ0BOAHqOIosHV/ppm383hWr
l/E3OWjpOONT+Y5WOKjy4yw5Y03CoVeM/+dzKzvyqopeO/XLyrVljJpaWfN+VTk9
6Rx4p3fc3q2YalHk1SJ6WMOkZG1YYvEdPXg4O7OapmxoyvXo7wNmO/RUZIJy+8QW
Gt9GIfF/91kAMxOO1LhrYJJp4GFcaZ6/a4d0iexesyM41w5ycfxYgZTSry/jKWSY
HEC4R0gIFGmXtkxnWr4ZVlLrptDnfANumxMy4uVEPFYmKKsdXaXy137r/dq8tT7V
RgXKxPD5S/7Rf7XTnp05VPoD9DDXociJdT7nXgSKbscJ9Jm9oc/XbhO5KHI6agJx
/woCSSjoDu3rk+WuCQmawVzsue0AfHgs+sa3f6rNs4rJiHOmJ2Q0h1gAB+XOF34c
EQ5OeKlfXvsEe976PfwhMMD0QAeDHRq2vv4TuWr2veH38nrq2tns7XRz+Ik01Np+
UsIysE2FnfjUTTjwqaKElDcOEspExObWeSjaIpGzleZTwAKmXUwV05aUoVqeE/+W
AGGsRWrhHm8livmufT/vNJM9iJglUKkQYPE6L2Pq4yURxrl5Ch4fOgs/bAu7Kzu9
NOY2rUJl46pyQ5YkbUOWbsryiV/opGHScdBPLaXjDK6FI27f1BHVTb+2ofpjqX+U
/07Y3MxoTZnzY52IS5RAdIyyMw15W9vRnOonrLa/7XBZxQcuzmA3bl7I8svBIFkw
v3ge4M+mGzqM66vI71WbCaS/aGPzoDv5qHanOMKcUYcdeD0wcRCjrlpelOWO45Wl
s48oPL7z0OXBsN4lVTcNDZBfENXXPRBEB2jkC+hE4KEz1RiZZHWApNH2VRbKCTp5
KjegUetu5pSEUz0sH2FRAG2fAkL4PRtRszXmDa8KvRiCgUSIUcn5QVwXwtGo8ROr
HOk25x4DGbPAwBISQCauDgJbM2rv46ZOXCWRBn6NtS9Lg8jl124MfhALBaPj+gST
bxHlhziTX4sHFSQBXxsqitDfi1jvx7i3XYWj+dI5UlbR+i618X7bE4wT01u+FkhU
0w+W4UeQVan7700d3n3jOIysk/g8fEKT05xQqgJX03lp4hLcvQpgG36Qkp038/w6
Q/tc19CrVV046S1BAeqKxMpArq/tKLllOEEBEezWZNc1+ydDfOIchbiJfIxNyWKx
IcUVeGg6FtWN0Z3Nfz19lIKU1WH0dwbovw1+WAlBmsctwKq6pXLQtkkBdrRybJwp
mQzkt2cf86phVaE6FWYMrjZCLwm1LA/cI6r1PA3faHFLbkiyngnDnuNXiunhF+lz
WvNbrNetkYL0EPzW/MIHJEfAlRL/1FYilDDk9eYnSKHMp+pTik9B5totFyC9CQgr
VJO6XUVSELyG5lrHsyf3a8VaNuVET7VoeTGl5NVVZDQKKwySjsPItszYhhBZ5L+f
dGHMMGv+qCJf3Gk20Ozc7cd3ieGxMhaqS2pfF0k50BGjNuASGzbU1Z93+tszsvWT
fPYbCJmaMhYNVPfaXMF5lklBhUz7wI7U6jv2kNn8fNVl9qj4cxxhGJUB1Ct2iWP/
m4yWbPaqpjX1OnrJiElSGmeMqvgjwva22NY+E7zdS88w6K9YE3mujXx0049DkZj+
nE7gx39KLOyZgDk7YOKfREBfSiko3HuiJ+Zh2a778xfWtoZlESF+8eyiCsN2itLl
cr2Hc35g2jl4r8bTZ8Pf5/nKgIDZttGZpjc/tm6tgwM/enbb5+gFouhMl2rRMVeB
+OB/8YLIbT+zmlEeXyA52pxokf4GKtVHA/mvm7kn0Bh3OzaBgJgmT4XMDBRfHKCW
JyfJVICdbNtEdMitj+rPLKhbuLLC8E/gXiC1ZoZE/mSWAMyurLlDE0ayoJG3WF14
YbYip7sbDLfaVojk0PrWXoiUzpzDBVMVAWt+ZBfFmn95yR7GwUlWyF5ggFL0A7nw
gWSVaguSTwbrCgmTUeq7zEkQD9mlkLUr82TJLOpg6LyOXz9I7cLeIantNI1KnMor
gHxji5I1q6R0putfANvfJ0JWFoRfL25FgMquhMaFtmU/nXjactcdOIHyIppthZAz
MQ6OmwgHCgbbHHPnsg8+Uc5yaZ9bI8UCEPtSdGH3aDjMHMtElkE8qKXD530FNWCE
YOrqR1Atx0i83fDaorJ+S67YFXq5DRr4GdwBdOdfU5D1zrb2Q3PbX8Q2jZ8177wt
8FFv/OO5zgVz5303WJJhbMv3ORSI3l+dr79CNUwr8UQ19PFRUwV6zACVcdBmi4Ba
sIgT+fdHj7OVL3YJssyjFDnsqH6oBjGHUfqHG69LSPABf2KZ+riXBGOTYmm7s1Li
Rep41l+EgG9KuaU+DYXnCdsEzGJu7Y6Wi6GgNxWfiIykLtvUKs4noR7YBq8QwH5P
LKRjvaNsTDPNXYpBRNHAkut+uGcR/Q4FY9sIvIWn/JvOLhaB22REAgz0QPuU8ED3
e5+Q8i9nYhkg4P8/Y8SA8YBpfXqAvNar94jDKs6b9wCJKW+dei7b+sYdschgmJHF
VOhhSrb0ECDu1U/sTPQR5E2T5gX6Fgj210kefq9GmTh1af7oEB9xmlpgnfeJNj4Z
c8kmXaRxEsuF/L6fG8m0iwBrQ7SVt9h3wOPLINn8Maayq/FyG9kpDsCc7rEiAdcw
0WsNC0eykqeKbWTedfmlNIJg8d3QKMarMox96uEp2ImOtqep1bclQIyVXcSZRNC7
zhCpKfr3XzSV+fI9vYGb7Qz/B94YDHNmKtBX0T0HQQArs9wCcAK40LeQucch1+sL
n6pPltNv20IW3fSQ2ShbOKPyWgeY77QiyPVTHAanQyu9LjQX92/488ZheGtjgKk9
eOgo2F33quO40CvOtmlvyR9/7ZwP05JHsjONlkqcHdRxUO6SiJEi5inZTZ3Bt9IL
eIOol8Hy/AenHVXh9+pI11yJU5X0l0f2M6dTuttNYSMEuS8qm9+MTlb1zXvkyFfH
sKTxc8kqe0Qn2o2mZbNHyui9i5+jZOrsk+eTUrbKKynVeCm5PtxsoInipMU6sFdA
fQFAwmQRxymxNtz2Eg6oBMjPN5Y0vkW0lhupkIJoOJ03Tc3dY93uyDcszGDsVzQq
zR+xQzjBi6NpmNo1YNoUEKksDq3AULLoNuQL8gnG2XWBZ/Gufxqv4fF7Mh6YUFog
0VCOgYBUMuV19is2ytJDiBdIO9o2kwIJHJr0qmAFP+7guLWmXUHYVxcqxa29MpPX
e/EummDPyphcwni/Of824vWb6SJne01GtAcerMJluTltLXB/buaUUoGphyCev7v/
ZRv6J7hMD8fTyCfbvc2NklRsaF2rdCyopyKEVPXAucYOwcTab/dR53eH0QBYAk6E
3ldqCn/9R/Rck9yRHMMlspkjn2+4wD4qXB6m4dZIqK2j30OTWL5qxSuue/BYWfAe
S8T5+c3sqfNoVyMi82PKLiYoPVAtt/4eYfd+l+0M9YmjLH/2CDgTFGJIQVurX3G0
Bi+ijtwiCl0c8dsvRQUSPJWrK1ZlSRSu9yhDdXkhuNPmf+RGQHQyChob36AZxNtG
iMS6BK/izQqNDJU3l79e6fNmaWnGCgADUvAj7MI2ffJzwnv5uAAvwcw71zNsqtrc
oJyxqfDLwmOibcyyWsnl3PmznOh6l3zI2yoXZexNs8QuizpEi5BlPVkXadAxdWJy
nZ+c71Afk5/9bSB98vZtMkKC9JXDlVVfsCAeRb4tt6pwa+u/gLjIgJ3oAE8cih3h
Z+pJdTIkMMDEdiRdCusYZSrBu+qItfaqXcHRRTVBsMjtDlkbIom/SeJZiwqXsqIj
iRBUnssN1qyPgKXnr3s4h9gyLk3bJ88EfyOMTc2Hl+uGNsbnhA3V2SfBxj2GoGfm
HgjSNeQqTQtHsSHzXwg4wJ1OHlRAj9ZxrGmVyE+jsBnu/heY2UzY2x1ARmoRy2e/
9JqJ/h8/CX8MuZY3Pbw1ot76CqALyack5LItbwcQ9yS77xRps5JRP7/SQ7/DCF9n
cy2UPdvM7rZ2uelZYj9ZZxZEuN9YHsViTZ4La4v+pNZRC/Ie8btSLp2TUqt+NkCo
+iDcVBHJanEjnOYGG2gNVYNQYE6Ecf4fEqjWh3GRO8H1qY7HCWFYrxBKHPMwOIYF
EFikpz0THBTMRntpp05eRuoikLgqA80xJdcBWQ0rvJn97sk3rxJKyzLTSPqYG8r6
j5MM9RzQ25Ec10HjMzKfrIwvs3GDomRIxO9Vp+Yh4Rf4Wc993/0Wii1bxuXBdm7X
sCKQQYuqE+zkXYU7pNgk08oO4NNJ+ecJ22vCl2/fux4fWJZWuQKWS6c8aQDBDVEY
gTLC0Zar7C7EAQsaTv1j5vEPCE97cHuRmxA5UE6AikObJrs0JYjGBFdnter9DpvE
6a1VZM88fRGlfXVo37Np6WX+/GxLyuyPxBYfVrRlaYLIt0gfVjsfSx4UjW6RcE/b
SwdKWlCETLGB8+Q54d9PJ4IPJD7Jpk2w2Yt/n78rqKP7dAhPGLk8WQl3qlrTxiJY
dlSAi4NORkJJThgH3LtX6WahQaEpLRlSWGon5rR+6rEW6qXv0gVIZBMZ2HeU0yam
qTOsFWze8cMrdXj9CYejq/VHxMIXzze7Ih9c5MoU2pm0YvPuhNCVEDr9nNkumZdc
q8GYJsbtLrHQCsqOtmO3v7lk/TCNwoJYf4ZwNWnuV/cGbWD8vSVkANTAooFmgc6j
I4oLfZ3NYz47XKdlfleda9KSXA8a/SDsv7ZcVVbx+TYOEU1URNuw62IUBP2q0VOO
H+rvc+26OL3l6zGlg93KkNwryKJzHcsdRSGKsNI8Mi5qsh3Mj3hl0WTXjpWa8Sib
WY5XmwRV7iufi7DcLVtoBES64KatfNn3kScIhetLN+B2JCMSgZpSKZGcBsJu9FKx
DAo+rpK6oKP5zc4ZMu9Se0EI4leS+cWsWgRodFlLGlb9tzm18qCJzlom02fHgzhR
bFxOFs8e9LJMFQcYSUxQjrH2kseCk/IMPDvjU4HXUuuKR+MRDA0F/lq8HhF1e3CF
IuEwNvPr4Omlczg0eR6D+Ci/44VOj31GHF0OQsK6yByBR6fPNBXh1dAB+b9zCCh5
6ok1L5LcsxC5sV3a0Dq6Zlro/6kZqQc+kFIfFnUAY8AuNvcGU7eBdiu18tCPTz6N
UmQzwJoXcTBXyDW4cHEHLUhlN/5Hdg6Cof4ATcmW07Vn51YApyfGT9DUCZZYsUGG
E5t6gRMfsTqPkpztS2MvDYagaFUmOm5G32UO2kk9sPrX1b9xH0Ez0Y3EM0h1tpkB
uXHg7Bx7Fg9ArM+/wtfB46nWVTe+LBGQBnESJBxmG0WU480YjMVOnI3OvS/ZnIS0
kML0YuyIbmkepJjUTV4GW5jBkNpzAyIuc/iQkC3HQ2vZWS19S0iwzSXlkxfjPXBm
TsRRFXn4sVhlPaSy9ET0/Tp7TGbs1/gmRs6w0tak55kw1VDOEASeBb8c6brWNurb
RJyUdfFfgyPr9UAgbBdB0cn/X4tbAtjm1M5JJWq47kY5IlxNxCLO3Gt+W3l9KuyR
uKz12M9LJEkcrSFnGJySLHMQUu8YO3ZW+pY60FyBDM5iHYT/b34fcEqQ2xuEoGaB
3tHoYVcMZuUbUDn6/0HOkQDGux5Z0Y3EgmGQtkHqn0zW0FPs50LFjbM+dQ9Ly8NQ
sE6dH5Dwio8l7IOf5fGxV/Vp+eA7FYJlLL/fOWVU7dPFs6MRdTI2TJFm9rf26M8S
JN8OxmiHcys+g09Xe4v1CJMHc7OZ9cWzEMoxVWxAG3yhiRi7+zf97PmgNugp7J1b
Z84x5BZXTP2pJGCExFm9g+BULk5/eQLJIdVWdmZXFzA5tObFjp53ErHF9lnZkL9l
Rr+7uCt/R1sTvJLkTE//T2rLJoTfEsEgCeZtQdmNXxAYaHm4HgzYXDj19I8WMV+J
Jat45xmJ6uKgQ4gAXqBTn3zMbVR3P1pQWRq4a7O23S0OnPQJFyAs2rUO4Bbt7A2O
yMTqhV/KTfnEVN17KCNSCj4zq51cmPFKEjObuu/EHaRc9glo86pMxX9m3HemoJfe
V0+d9JSPFkPEi0P45pRuRik7/UxFe2YFZhYYqkjloggocuxtvPoO4/NAxbz22TXX
Fpgt7PxPMuy1Vj0pfe1trtXt4BXz9c75jntw83ZvzrYC4aVH1Vip29YPEzg32J5C
l0hyniW4UBI/3TLKgGGtbKt+xgY2md2kXyOqScxfkg0bMbNW72J4HJHkgi5bWwF6
8f9aYMhi/DM4koLqkl/g1LpxoVmNn851iXeiBSIKt1ngKnRKLDeoMvGBw8MX2H90
fvdU3KbH4OM3TmypumgPGq7OXiu5P5qf/h28XDQIObu9LR32pPTLzuNnmkms9U16
5xaaggO3fS7a8Yv+yKMUU9z4njuPGDn1+ArWMXFEi9QLQ7U2jjYvFglohVaxQSG2
obTxlEXp3POrkKnFFW18LrPjJkPURxl6XHnG4bobFNfRwLuy913mlh3takU0GByo
klEapeDXi45/gydwr1RDBEBVLrXKEHrXmMm3AH7bxT0qcIQuhV1UM0rq0ZzeZVmc
Az1T/ue1UpmtFH38x4QApuEg/sXTMP75DusqYENgSm2gEGsDMZ8d5AWHdbCnEyYc
/g1c5pH9KHYs8OmEgLt1Q0qL/0HUyOMxAk2M7w4rnm4x6J2StjJVi1Ef1ISQPwB0
aZiP+1gA+Kw0wspWoMx/7aGX0R7EVasDV865ikO9AKiQhJ6aWrRmTIraFCrmGIj5
8G1xt+o/wtcibV4bNpcNeJGT8k0KW3JkHCUffl2maUKP5Xae/4nSBDKXOotM4Vpx
NohkW4P6ENh6MZLqZE5K/wqwuIxd16vqZkzxoBcbYUWfrJCKkUH3Ei6ATQ341K7R
Qh9syX6WhAU56Jb/AWuIjOKPZF+ACQE9w9Kd17kuOq/T1hjK6ItCs6qB21C7KFxC
fi4LUV3gTMt2s/F6m0ec9/PWoWGObBnxYqBPFPk+cYpKymUiJau9fC4V0ArvybXq
FXK0sJgIXUpKDir/HRBe0g+hVqo4bzDGdhGId4FdHnPzMJZKfG97EbO1R7rkeyh1
aODxkdGT2Q/4dKRweWyhT0eR0jf6TLlHa6DRGfEyKcX2At4NLZfbQsxGY9lXBcze
tVQEr0YLaI4mhllf+D7hhjygadThuuJLwz9tHkkSfmF5FURDryoJ5t//3fTVA9AA
PiyXOb9pfB179snI/1en/D2S96F4Zj+kapso+Z5v1SMWU5qpWN2yMKUoD4G2HmNP
qZH1ZTcQnfXakWGSliLvcLL+i4sVUcwBITBRkV+Ys/mtuRo3NMzWfK9oYwJSso+l
4/HetAY3WM8USh9L+gBYiIsedQW0X1M5iQwMWSavldgx7DBy5GuWdpWhQhObR63j
VBAoPuxrRhSFEmtCd7emTLBrKI0rRoNCQ1fgDOe9RQFAo8w+IM2C0UoL2NSDe4ky
ROH2GJZS9+QUTLm7fz4Lop2FauIvWURjwCcvb2/W9OeaW0y2QUa/5v4ewXJPI3RT
+E3R7zVNfQLbxUq5MdQ2EYy4kKM+D1gJNt8K2UFq7whbfev8P1oKM01Qd3eveUde
uJnzzbO1orcY81yLyvqyFLnXJ4g4XXiZYFCc4zsAh5KhzhE7Fr7M31tDbZUQIFZP
GYk/9nrqGWAqMz9y87RweYVveEt/GtM0cqJmJZzPTWw1Um6NvJj5skwt2FwD7izn
UAffGMP4zXWt9ivU9gBXFneVTSWScK59tLmYIfMY6qSnz0TFNYNBtaPAAxTvV7j+
coZDoTVFp6SsDG4t2nYKYnXN1NEGWwLmoJJO17cjXcvqvls7RJZ6mFUsQIZqFYuB
L3YBNLmjHp0X7zKMsYGN6VkRU38UlHC8qG5r5zIyfHfpUOm15nEItvH+RQcFEvU7
Bv7bag2vfPfaSUd0Jg+SWH3S6fnX6c7W0zNo5VEvjDehJ6NRGJHki4URYisvnxzn
NtpynAOI2n+javb2/pwRVWxhqG9z/qQS2YvztzkY91+wAx5EKxbBtfsHmFpsD5yz
sYGQqxMrdh4uO904Fti/9Q1vvKPcGGVJI1AuhJF38uCmqhjmxBBcrehUAWYNyQXO
ETqEwSnenwodVwun4LxA45NUDVPTEdw9xGAJQyh+4HIT0hmXWvDlRBatb3FPDAoJ
O2PG7zlkXyDuxlu09MSkdu8L993/68xixv2SC4cWLHDCmXY5emFOMK9Az8klvvM4
iDMSaw4wCL3XCqRoFxtv23W3TGNEf2VmjpDkza/zOs0GPH2CyQooPY5+nNRo5lO0
cEvesmOD+IdLzgQp2qsK2rua4/Xqc5sBAP1kEgdS3R9CvvL+896KtkLjXZZZAaHv
r0lUrLq7vOcLV5F4mPG6tRubtp6HJZup7uk7n+enzUeBdxKhNEeX16sXo8vf4mqX
v408k2qLE1zbVDOg65+tkCSHI16tSmv/hSTIVFsbIOgi0lEYUBBSRwImOKkK3Zu1
20Wtw0vB6FPq9d9lG8CzXyocaFGQdruccLo4bjk6J3hy0u0OilyqYvxlmitzG6oI
GT4gbPeo5a8F+aQlKUYQC5iv7udm9Z+UWqzfjFsBq5cjqbH0324nt4cZEM2itzDz
L6JGyoOgiqWucRJ/0e06VqSwlpzqQSubxy66BcSSmmnxITQE5zkbjwd0XReRT6am
AManAgFCN8MdiXu1rmiNu/zQPUD/ha9L6sQnrFxLEKCVcrfgAdcIuJBoyZFg+6b5
901j/jBe9Tt9gwBS6VBp8G5iaGoulq7VJFUyFmOGhiezhwx3YL/0HMoQ6896PzgZ
kCOR8X+kUofJ5L06yjbtHS1XWgHnwbGHbHn9G4o4k7mc6uR0XHraEv1kfhH+Uv8q
xpS22+Q2wk0QkXElZW6eioTtM8zh6Ep0x9Fpg4ccU+tPaP4bQQtJvmzIwCjQeKh6
ARb7jBmRoJ/ixj3XC1NFKotMQSgg6xVNGi0qTTWPK81zJhYCme9Ju1BftMSgg1pQ
QZ9iWebjL+N6rcp5t3hHIZGwZskEAtRlgyUvcLq56sjdMfRcZyVPySJrvdGOTrGI
u8k+zl3HX3k3PD0+N/93XzZvGzElAr1/PpfH4jP/damnQj1i4M7xkyv/YU4FchVv
pNLtfTr5HEFdh82s3BuxZgX4IhAHiMp+RSPPLIUrGcP/6QQpBJXD7KWU30ZCEGRd
rGW/Sc9VmogLhGjmRRPodkJGOBnGC/zSku5NVDsm1uIdBg+ENdZmf4W2bEtPJLgl
M329t8gWdCkqsqTaF1RaMVyFNixr2szlevSTYRRcP+QX03SrzwDuIR3srq7Fb+Lv
EjyP4yYtLC5v2AiulnWvfI2Ok+72+2Og90vAN0k3gjdYiWIQIpYwIAUX+vZqy/ar
4h0F4E8f+y9bCeoWeiB/tYfAgtUokv3xuCuzVaNvOxiwGBqc/fQSyb/BFbZXvsTq
s8bmBEdoVu99hYZm2Tfc+SwpnOOxZsDLfVm3/tVqnzhZkM+gbxyt8bhF7yfev+vl
qaB2FNT+HuzuNBd1mH7pf5BawqWB3GLTHoORJ5ctgjwLHIhyt9qm27waFof5CFuw
5HBtx3ffaZB4x86YUE/x87GEX/f+wohKDAw0qgbo+nc7yOIdHjMCB/XLAyOwGwkW
584uISoHufGB7qj61ZiIgIR3BTaGtA5kMRRuZf3/G+Ga8Jm+kYordCuItk13cMVZ
8rMnJ+VLsE2qYomyVd9tMHMJ7KcieAX1Jzt0fkYw/yE2fCrSe6O710N5fy07NLrE
kwcAmI3nHA73keW0Jbth7IDkibfdxQQo0bKRa7nGF7J5IbQiDCbRA4obh0WjeFHj
vO7dr9ODowvMar8XiK3DyIhdIaA08A2zUJtNYgYVcYe0/hrulVQ1vWPhwy2hSuWx
FVzlYbIsZGiH7hnBQlMcP45H34k3si400A9wsYHNg3iZ5jigwMgcnUFQbJTlfMXC
4xIZ/zUeiFvl+V2FKsBHZ3nJYMLpR5nV0Caw4iXPjjFdd5mCsjco8HJR0mKEm3Q9
wUOijZUw2wqfoSW1aSiyEkE7/A7Qcb75DadYTSKrRVPn+AYT3V++RaHIQsR0VsgE
6Yniq4V3j9bzB/IHVRQqwTX0Dbcxvts1vqqugOmH137LhLrSlf/ST65pQ5TJfzZw
yZqhtfUCevpLjU56LyZ/qXYnh6hchlqTBc9SKFDAsjDOPfvRKGKpr2/W43isrc7W
YtfE5z0BH/uCEizibMFBDMKqAqBxb+qslVULbj/1as3TiIzWepAvUF+PVj30yqiv
/FpR1OzannLiyl0wIEBXEhrNl4gtmqTUrteSZRjBlNJWpf9dCP26dcnC6iVKp8T+
ldoDnE7rgoxjCq3N1WXln4O/fHlA2r6MsQJX0DEKg231ri3mmcB/a7jaRF5xK2bi
o3Ld17pVazpOqrcbmCect3/OZMh5mSdlM5pDaN+CwN7/lZ5K/b3qniW6OU32eChO
cWvwva6uZZjKTP/uMo13+jqVWdYRKxAC/mkLF4XMwk/SDyc8Za6l0204gVgTH5i8
xf3k7fFNlWVCQhIKkh5IQg4E6yaeQDvheR7T4RvYtILOgLBIYoTqEVQ0aU8NoVOK
iDkf4Mc8d3jlMTpnuKV4l7rgKTm5yA6I8svncf9B1aZPneFHpQEPmG8CIDvFDlE9
9ysorYYO2HqHiqtXcwThhk94LaHdbTDSyh5rmCLY8mjuwH9lYucqCvzAT8hKvsg7
LH09HKKEVPAqBo3/zSSSITvwVOyT3f46QMXLUVYo9Lrs0pX/czZOZ9206zpkI/4k
Wx7aqqvmfAiVIREtst48d0B9AIg5xD+ts4seNV+Y49EnIN0r4AGsZ63d0TuzW105
4tExIxSEHuVZ16W9cXjYiD0DZyYV0CwyAr4Al55gB1zuiYXecYopSZpmV2zF6rU/
NEB2CxJSw7RAa7m4pq2JKZEUjppuFvnrA8CRRCUtvQ77DtFk2LqnRMnChL5c9ln3
hxtUmywl9UT1qQ450qPjCWlXT1lbh6D4XxVYDbQX3AWvZKARVRGqxfuQyEuOBd6x
7zeq1soTpUHFtI+cPfd5hg+cfGH3zy5l+/wI4PWRiU0sf8pW7C8wpvzemcwz30SB
jjNOPAKDB4g6odvsiGt6jt7TgHhyTsGP7zXAuVRm0LeycTe/rvUXr/CagKaXWIkZ
dB8YwbHKGUClk4GC60NZ7+R8wAFUsgKGUdTAMy0HD3xTP7N+d9x0fmBk0M3/HT7l
YZh9BdgwVl/5Ldx57t4vcInruSm8v8Pcxn4cyM3obrUO/RWtUqP/gye70vYkzuRw
7ELIHkcAdwPoyRGregb6sJvhHER1JREghACr8wYXdtkYcWCZ6IMjJP4z/NCPJ2HR
YosjFoyYsCn8VPiyb0iV31D+aRU7iSm/mu0vAziBjcXnb3GnUastoQWKxC7TN1Gs
pehb48theSbkDQfxblEI8X3l8/Bm9mq2AODYH2fvjE0YFXXWly/XbBZz2pS4BwRx
w6OKdyJCg/kFKrLnlEyGH0pITdSZnlDGD3MLxF2U9YEmwiM9EAcbjxf2QvRuBr6w
Rg92dyyRY5O9LrDJ8Ihoo9Bn2wzyB7swTmaLDsdATUHhgCmil600TpMoR8Ym3whd
V11vpJAnk1iJUaZYpJV0z5Z5cRL1XdXbKJW1xBH9jPfnWg7SWNgntAxn5AcxRt4N
0rSYfLFKqrKJrZz0XnENTNOPRbToJwQwL+Xt4HjWku/1kGcj1+mUBzOQMQ2OMtO8
2xTOMneMjvlOD+qxCC2b1l+8YfdI4dPakvWctWjQm/c9knBp4vLS5ngeHsu+8em0
k0zdb8JmvG5tsGCTXL7zFI5XbV6znBuA0R/jFvmgRGRUNIrRbCp0Ea1DN3tFqBoi
tn8MTYPfVAB/nIXY/HEJX3YW6wtNF2SDSBhjrHu9/Y/jqimXiJ9InUrXIw/iLSKV
1VOZX/Eclwl6VKhxcm4a5SdW45J39XdPCg1mFyirXwuc+76CIIvlWbZUpFbPA5Fj
z6enXnXr2QAzVUc+QxdRqYbGiYwFSXka5ebQXQSZzP9+Tkgcl/zpna+oHG0CL4ca
IecxZyhQKvftgdTdn1ym7E9vSaHgcRwsHdQHYQMi6ZR2Op5Qoumazy23RZz2U7s0
0cha85iLdCK967eOU7VdgXvkfXJGPDRvnBW8yN08FgEKHNBeUXhqacz7pDEYn4eo
Hv/t/MZS0cDFufgqlDCYsSK6S6KBr4xC7O9TSRNwSjvJjioztPBnW5OxcyApSOWK
IvecnpY97PLQ5alt7r1HeYr21RkyHrl7XUXsh85OHtAo40bhGeo+la938Bu8Jtsf
xkANy9E7+vKTdg519HyVB9XsVH5FUcTbDFrkslUJNJnrz7B5AO1qNdanJtdHlexS
ioQYUquCwOdNrXHeAEqqMVRUEa7OkCwifGMMwX39X4WeXfyNWW4B3KKflYB7JB6h
mU7fUsoMeYDZcpTl67hZG/xmQ1ZxgDljKasWra1DhtmfSJY+VQ36CPMTQu+hdRre
G9zfz5RXBKyWaxEaq0vwvpQ5jR2kyfRm1J10HRZsElG60b5KMAORfshb8Vpc8PlM
zvOdykGayOjd9LvJU3fpLCr16S72kXasMa7waf6jTK15RWod4DXAoukNg77cwVFo
9+0V7+gTxUyZErt5y4Sx3ts4LmAPFrWeXs0c0QLEvHaZjJmPlSBMDQC8ToCZ1ZzP
Z5iO0/4CdAkY2qM27dXjNXiLw5Ric61dHL31ERJW2Q1MZY/3A9urEpSpdt912tzx
s1RxG89xif5vmft4xJCfSpjAVlXTYFtBrlgaKmX7OcW5NCm6Wq08FF3/RayE+q5y
8Fy9bnY93Zn7bqPtZSJ+M7d1LY6FtQ4clj9GQNTi/3EeWGg9+7YxfDS0oODlGGxR
KuyyFZY0nKdgaLnmSjU9evqPvxQJhE6fBZUz8pKd1Q+17nf/KaFfVC0vZ0FiFxV7
JODYyCIZjYHGbkWJBzPTAh3Ya80ZVpnifmeEUlBpRPJwkPKyP+HatZgKpehMMG2d
VF+Z+l+Ae7QsSAwwLBVAlWnFaIqkm+pPnkwovYsNvJiEdzCiZPNNQM0BfiSBrDV5
XhfEfgGNM1bSyovAggqxYtcPEbCUNU7dypWOjqfFDuuelgSvQpIKAkru+yPcO7CK
ckr2MBLb6COKLnC2crdsTZh47rKXSv3JFpkX4NlgeWsavt1uvI43nKodGeC44DcF
t4Bjr12Z2jRsBdAgyS1NX1HmoD9oIH9xbY9oKeS0ikJ3n2tuszUcKDra/Ag8+QOq
nKwBXcdpnPHkcWMEHcJ4hiRTVX+UH44nxo/r7376FtHnTLeA2/XQ2Vs7jWfhBNL3
Gt5zYgKoBGWYBp8aUHbV/eHLqOvNknwK9PujAElxEsKieOsbX885AiAef9/IcYvh
IIONmZUp2oDTNFJufgMnWJtdZX/BsIzIW1313qRCCLPypMjATXGC0WuYhcc8jY7R
6htyE9CkQkXGF0lrAdGUqh+YFkhbYvDU8Pawsb9xZc50gCSvZnd5wPjTqDcNSZuS
8JO0P6Cl7k5HNhUF/KThatYxs8pG9k4u/n+god37XKfYp8tLJi+iJgC7+v51Gbbe
zWJRbqUvsjYCMMQ5El5hiU24GFF7gR/Iz/5n9bgDGcwtq1a0QiIPY83LAxBKklfn
H9rCs6Drwo+kVH8ZXuglK5yW9p/LqFyDd10cuJLGMGusYcxiT8HbcxeMVG00hte5
nmsf9Ki2Ebk207gTITW4vvtiIjLJpEVPtiUYonBXSIUNvceOogKJ/ZwqUjlU5Vt1
LVf835cYujrvPi7wKcwifJAiumgmJqoy3L7PxW0uAMdBwosJzC0HpbOE8HvF+uby
qh4VlYMbkQpLlgC1DnbQPp/Qdyna6wnqZAtNyz7N/4Nxqoay8fKAZzc5QK7LeRoI
q+eNT9F3X2XPCuMt17Y1ltjAk+ENxYJ442NFpQj1PyOkT/ukAlPhFZjTVG2bra2H
OpMzOjcor3+TksbnClGy+7D6+QyLqJ8dw+AOVkIrIdYfTx6MxEt8BRAwXs6qQ35P
BvvqBI9+DIvlDz8MNNZUVBLVPTFeMSn7DE57hIlubTIdc6ND8GkJFm2ouwOhwkUx
OlYFO0OnGxE4tcnQ9A3x7hSS/REiNSgCtDR5jvRklyfhxVrNqf2rLK0mOpijtiHz
8xYv+/NkHjnMYJqrhHQW3yu/USdHsaG2FlaMC1XizcBClbS0q21T8Zh1fLiEkiJv
aMaWIG8p/aF5zaw1vZXuvWAADSx9whsoEkZFP2iV18Vgi9TgPmlhs7WuabMTSOG0
MLx/vMJJohE8xjIv5Fb63tSnCrzeFaxGZ/Pe3GrQluuv+OJmDiztpZufMamqCMdi
eAsbnfx3OyeCMC4pZWfRCCiMDCfK0R2a1w/nHbB1CfQmu2oW/+pjFUrMo1r0DRM9
lAp/X+EM2RDafAbDbvbGDGM/oJkGA7VKeEL/hrsveQF5CbVzGLZb6AfLfCl6S9yi
PzqlQ61S2r3vG1GnXrQc8UYsDmNii22oJigtcI4KgqmBTN4MJdTxzUKPrkQxHcBg
0qLO6lqcI96skGNbJ4jusZyKt7lJ+XRRQam0VzmSYlSBCfUOZeDuVEavV64ZpTlb
/kY1XOOQaQkV1tPfdNCImji8ZXXZADrWBKBHhKuupsaR5p5esLhLv89Y5+5Uoqz/
yAwFgKTi8acEOvGEFA2tOorsoxGkUqLFqR2faJ4t4UnM0IYXYBnk3NKuOozJTA+l
mHu4tj8tf6GaqpSgmlOpg/HUhd/+KtJNfKwKXsY6rlSZ1YbbxdlJxqZrK5KrNNJj
0Dn6ceOFaxHSdcrryaCw3CXfu5bdqJhPBuWw9atkTC45BRyvIpKCvf9MXf3u9HNF
7ygoXIkF1n+YwhROuokPsdl8x7KIR61BqIf/y+B88HXy4gGDtk9DWzFenmMzCNKI
lYCWjaV77XH8O4sda8H76Q+SIL3KYm4tyyfTWQkqM1pMnav4fxS3eL9n9nX2GYGB
CoIJjXNTuRsW/dUhO8lEY8qvdWTOSATQet30xC6ZfVcgXGQ5182jfWTqlyi0Mfrw
472Q3kMLjKw1cz+xwl7UftJ6pERRHDEuy9bFGcyuShSALhRmWarSiSYDt2wxc6j7
b2JyZplb+C63pSmHo+dIETZdCenHKqexAdk0du+iUJPhMUybZ482ghUW5bMWlmSI
VInydyyE5Sn2NUGqAPEZjGAmSgFCj/qqMVR5wr/s+FQ4lKzTTIrd/dN3IpNkPefA
/tJ9kN0fxxkmPii4G/KclMa/wqsSTXvMpoeAqvtUkA6gVgKzyTing8SMdbjWjKoq
SgJCCeUq8qOrR1NDCI5r3uKURHnf5Ohh20x+ZwPdM0oBubFSswyfYz8Pzz3LEpOa
nALmvvTeE/+j+p2MbU34pGkCGYhtmCF6/+dNSmOeax/sfrpRTlJTqPFsWOuA9JnF
VW06Y6eY1ZxMa6vmPsdWiCpYNRxmRblvChThk3QIu6MLcugWUC6kedH+PeEccO0g
rxn/tBW7f48FdPczqjtLcOfqgX4czLl8UsHrrV7k3kfjFdvD10swymp7+NgsGcGH
jwsM0tm+YSv6O4rgAvbRxkwtCNbrFwad3hygDHO2m5PKy7xIZqOL06/dWPfxV1wK
Sezeb1J1LnB5I+YeTLumZEOW8f7ZDCZdpkLY/++VcaL+Ey+5CHnh/QdJEadPc+0a
UOfF0gnVwj7GoqzHwA0BPQVKWSnWt4FOYytV4p/+N6P4pzR+dapKJc57d33tfxJ4
iLhCnGllzgsnJHmD9MM/pB+HGgtt47uGZxAOoHTy591itW2zH9WVRzeu4PIhLFJe
u2f8okdoiH89F0RIL2w4R5iLP1V2c4ByiL+zV43iRDxYpa7PY5yVLa5wgohF4GnW
52CxdRQMU5SmnHUP46J54TF9e1DX2HSHpsH5erbk7QbJlAjP82q84nFjo8qOihIF
jqU38WrbgC1BnmcbYJ5i48VcMLekWxZnaOMlJCbMVLnPvbXotsK8K22nRpmMjVeD
2HSQfSKm3+K6/CsDUV2KOtqFbX50Gs+8CmWGpmEwYrSCWPNyAWhLE10nNEAy04D0
Ul0Nwv55DJ33/DyOyC9/VrA/Qfar4ACHm2M7TWcFUcoOxGgoEzsOztFmjU+wIDyZ
aesIYzke22psZ4IqwVdazqm3pSm+ojnLNx8oL7w7BytgrpBi+ykArfzBM/hSCtZ0
wF7RW73FfGCwCAuh4xxolGCu1F+oI3WhmWZs4dOzlHFWALGJmbu1gECqNLzsiGOD
8nu3apIT93bjmJv8S6q45yRrdraiZu1FSVDOWT8hjX6C1YBZl9QOe8Y3NPd3cUds
ZdVZRD+rgbzldITIYfRNtMACqZgu/SgC4GjN5MiQ9NM9uuAfA1YDwIAgbfyQ/s+i
O0OWtNzTItiHe6yGNeR6cvEtB6cwQcqiJ37SW2RUt71s6dbB6ghWbFfU8AGaNbm6
KTPLOr7inP0J5pq1dL/roRyemFLejZrP3xH+Fm0kw8CKVcFII2vcc3BzvYxxe4b7
MYaQhkL42WlbvkYAysQ0nGoAC9eiF93fTRNaU9NIrpn0uPd9vR0opO9DgxIgZ5m9
g3jTV0I+zM/z7vRuSiQ8gDfzsTEeoreLGhjsacguRXMRaTqbfyl9cOAeKWGUIr9v
TNJldwvshXpDukqgtRKg80Juc4nEHihqnc6gjiTR9XM6bpA/fz7qqqxU8HgieMj4
S86CSH/tvk68fpIv6Qc39wKJYON+XhHKlTnO4I+iR55tkSihxKkIveugSS9GkVqX
9l8BHVMV+hR86mfKxEojy1ba0zLG7i49U+l2Pf9Yb1dJ76IcwSgaGF/mrclMkof+
WMi/uvX8PUippxiXJZfHilzuGk3hcOMR63mKKZBzqs0BuVTmdoMqmR1ni2O9e72m
q5VJ+1XpKu5TP4AK6j0Hp31f3ox4py5yElfcElLPqd3wJuEqktOMdQ70+gDLfYcT
uYpOSgiLOuZL+rp07dYq0jfKZBQ66Zs2jA5d9suB73qxwjO3C4MY1Z1CFk9yl/2B
9KySxcittyKS5MZ79lrh66Bfqiqsqq7gbEnuzJ13azIx0Sj4W8qFJaYBJzCcBUDi
HweOxle0OEDAPHYgiSSvRAEm5Co/xcXG4RC8SREGslro68r0eZI55qqamWiGPCqn
OKca/752j+e+LMoGOlsqxGj7jwWB2HCTssCUshWa2LpUVefXPHWuYIPgo4P8Vym4
HYk8WOiZ5rid7a+fYFJDV/4vCFDxumVDk7Zi2fi2VDFQ3rp7r8gX6uBbSXctujSt
ZtVcgZOYVevwl5Rs2aN6hYaSJ27njlcPyTjW7vaIIEgOv0gFECt5tGSku3xQjHnI
Dbg3lgwCotOOChlno7IAT+LwzNo/9sY6ZbC+LJzZpa3PTEEhtFE3085CnLOQxfD1
1B525FcMPwmjjfZR7uc1rHjfAjRMQxxncJY0JkNVg1+Bekbn2mQwCdTs34DpA42W
b/aab6Tqqiyj/HBRlfYn4JlP/o8OU1zToOJXzP13y3DJWtXi79SXveS2FLu2GKfA
1fZc7p49e6f/4njMAtGIz34wa2B1+0hafrldz25qmXAzkS0eebpQCEyuMGp98sQS
QrsWDam4z1njDfVH2ZLngZdn1sFAo1RXhZoXJHrlloD+QIfl5fc42BkeQUfkAuYp
+QWuE/G8z7NgrbkCj2h3XFwbG/j+DG6hr2zfq/oe8XgSY+usuoB/tvAuZpFSR7Hf
MAsqujQ0Xb7P+JN+CIaInDVgPov23PczBtyoRM7bG+jNmBTuYNy0qvP2RzdLlFtz
cVx7XPRoNcoPoHPZImKMVcRemAaJQYnnHAlWh/tWbKL6/knSDxBezWfPiyyWsXRG
rmBHlAfu7vnTwOK+tRLQbrzZwJW8Z+qrrCp1oc5zC3vli8aTUqLwgWn/ADCTvYRh
t12oAnQe7kFmQuPRRj5iPRU2AUc8GICbgnDoH0v1YCmK+d0TTyvDYLCMwowQVK2l
m24EkO69MJfGi8ZvSa1r3O5BR96SNGF6vVDJtf1qOQGCQUKGlxTxJ876i9SYNVBX
NZ8fJ8GTzKbScdtgX7QKfC0Ih0EmtmcbOFSvbLfcvgejnQ4O0d3/kO0zgenywSI/
/OZrICvKu4GABVIb3H/hYWjTS8hoTyy1IallbL98433qVkddl/p4pEubWwnlmJmb
fr0vsIvsQzqNTK2WntwW+RI6SHddPHjvvVhDd0b6sV+MoNOOFJw6UBFlUi6NtTie
861YLRWqOLt55DdRYBx0Z//yEKt6brprlTnraqySuKKhp3RyRcM+5c/4vEcZ/+Cu
sut+V1EnO1iahCSmCDtSPWF+eogjicIRT6nTOHDzB82M0bPVhgL9m4t8jDoX3GQ4
z9k72G/15u3WtYCntUftf4DZIDBTKFToV06Pao+Ahir4uNJb664fRCEnfP9Wfsa/
19eKypKiae+sIQTrJj5/1bguxjrBys6RqNfez/3b+FFyeBLfwvEMVELjix3oa/S/
BFygchlv5plAw4yp9ryX1ep4LswtENES9Ytn2+fnolFf47cid6BGu/E+slvsplr8
OZuC5Y1w1D+/7/YykEohS5GvH/mk1gso2P422BQJQUanPcN+JufYr+hpbcBiImz3
SgyuxV47J74z5Ld2kR40fbm9GCdPLvJD8i/n3IR0Cm+2d4sIMA2PjgMoXiGCcD3N
JRfzns+NCJG1tJsSjrgh0Dw3kx90tgzVcpzVoFujY6a9FJRJovzkp1lBaOAE0iNE
CVLVSYjd+mgN/UriRWWhIQoY/ToZWa2O07Wkdhv1omkevvWYL5QpzN5STe5LxuE3
xK3WSm+cJaOAI6B05e/aOOKWdSlFWNB+ZGMaOE/McyRblVcGTg/xq/ViQ4zoCEhz
ZMqmTMo1DDkOtt5eQ7W7XPoPS4b62OqtxK2XjdhY0vMTxUtPru/wmUlZxiM+ou1S
UdXbOK3Dz5CWsWgoaEGOWDzr64EFqMn6FyVX0wKzyOw46UfjjS119fvJq+nMj62+
ZSLdJ+CAe/1OOjbl9+6++db3xTg3CexqlbKaS3POClQLXp7pr+yt6UyGJrJkISKe
YzdqCj33zh7kIyGqu+tXx4OJtrHZaKYOZATCtkdbf2JOzb891hTj/NJnKH5KXEDX
fHtAbh5UEDW8ZVmLtN1+HYhLQ8C44dh9Rpy4E+Kqj19HbCdcvb7PRm5/4rjWL5Q8
nRFWMNTkHH8gdlIAwAJ7TemqtRnc9o3rCYLX6oQ7fS9xR5V0YvQkCtwuZuueLcQo
s8pyjKeOnmMKbAPtP3OURK7JaJKtb655nctyNsT5xMTcXaxyvaaIQqVIvL0gGdI8
s5vtKTeSzkv+SjW8GFnbXCoUGfGE8uPCahPIKqLWEvLKVVWk5C7QBFJT3D018Uwd
L3+/4CsGRyJ0K2+avwX3mfypaoRcW7538wYvJ7RgYfk9UrK0JETD7RIWM2G9AFYd
J56cTe8prQszKBrB58vb1AXcaKdU74oBPBqpFPneRC/9Vo1lMao08dtq0vbRoO+T
OIt6oH8WE9lcNFM0KkQb6pqYQRhcYIjB4dlsNAwIML5alpTgwRIGryUFdAt5km4/
pnunQatcRgOgMQTbaQ8v7O6yUDB6LAf7orrou6RnegTjF6Sazt98QumnDVmc7QmA
gpe0o1+tiYnNG+BKDdrzCpzeQ3fljNnCmGtB/KqegRhDoa02fC8iXd9wpjQtYoT2
FijElpyz4lEtWgGLQHa0fGz15/kTMtXmx/kg7hxieA8aMFvEe5yBZ6tPvJTnP1gT
Py8iKCctPo3kucKJkkNca95mbbGTEFQEnN/Oe84X0WseOcNxlpfW1cUvQ1oWx2Io
U5TixT1JmxiD4cGQdsjkWmKlkxG3nGpy+xR5Q3ZgjvyGBE4HyS9KBixSMALKhwlx
dWNBs2LVxrt40OAZnyRHV1N8n7cdFJdLgN42A6P3i+gYDUsXyq4AILuYV8alQ9KU
vMsWiQHrYOjeOuopgSexYApLOEekqn4rhUZlOh75+TeJvd6wxgixwb8AHuYqrkBV
wYWgWRMN6aOW6yv1hRzp5Tl+ElMLk1R1fpn3q4YbZihi4iE+4VcarPf0CXC/NIjZ
SOlMgei3+zTm/Ar/gJom5KHDFr2K1zum8UTFs+IVxXc4ToAlGXxlw0MjGfUpGRQU
mfjlcHV09HUpttPFA/fZeqrfM5tdylXpbnJAoEYS5D8XSNMFwXJ8ABR0bLZNXYq8
K322hf4U8mFXcu8hThCQU9LZgg/GCKWr5NaiGCZHosL6YGk2bYlqNZlAB1ZH0sfj
Ue1ZQ73PyyhrXVjywDZffcoGUKHXT1GXW/8+FgB1RkvZFdREVaN7ZBSUs5kKiJ+K
XLIsFQC1jj95Wjz22m0hos+iB5SuetgA2xuztu9HA+CFHUnIRPcXLdPCW47EqQ3M
8kg3Uoq58bdQYW/mnWdk7poCUqgvCF22Y9ORc7ja0qeeeqqFUhgz2jkJevBnyPgy
QlhldtJphm/LjCndVIUx6NgqfovOseMmNu7INH4pATlWWfI6CoKHoA7hEMlgWZSK
BalG6htU3nDZ/e3J2nN08Ewwguy7X9enT7HhBsrdIspH8S5Oq010+IPd5Qg/71xG
pavrI+Icf167qhKLi4UsHPXNSzMYlhcrmlFtjapLLQvbLZULmRcOHP85RCwdTOsr
bTy3hWQ0wcAkpz+FHGPh3QVwgNBYFopjH4ZdRGW3zvcuNBe7Ria3nJw+rES8H3Gv
uWEYr7c2UiHRtGiCQ3iQn0EvuDfm1ssuwjAtb8KbnjgvONPeFMR/hdKVnpmDqu4w
Nav6Gc4qa3+TE7/ItHTctB9TsCVfx7WyK3bkVMGP8vI1YJuvJ5fU3KLnntfHcCDR
DcBbhh99lQuVXFA6xG4hTVhj74tH/K+5pOfEuPSe0U+iCooPMRoWO6toIuSecRoc
/RZg9YYO0QfMzsPjpKNV0kCG2Dc9NHqGunhhslrE2KIDoRaFXMjPbwdAvwD7bZ6x
ldh5tNu505AlJAQ5xu37rWwPGf3qezkQAeGmNPGii+xnF2lKObeZK8mmw+1Ymq5O
2aGrkVnG0wdHmPPSLzgywRa2F+BKLhSvkuhjWfibeso1J+m95K9582k6SbRHIypT
LTbB2XSq+uAZkpsHql6/QZnDpfrsXpx9AJkhYcBBHk3WekijXFtsd4TwcWrC+GhP
UQLrikaXhFx1TnGEbe1Ji7PNDUd0UDLpKLvqncYdSf8MAM8RYmwtJmjsYqez9bgE
37bg9cg0/DXC7w8TY7d9pqAULpVr66tMMkeuR/wqjg8nMtghazG1ExQUaqBaTnLA
xTrepOF53BBuGRc6etXujUp8YrHMVm19hlK9A5PZStYB0NQ7VFkLVkO5JEo61/ox
aJuaIHWLr6A+KJ4MyvB3JmPcOpL2ajk4r7OB4BZFyy8VY8SiVls3/tMUJ5gfrs4o
IORSnEWURhckfirmONdaE82Sd1715gnxYAuEaOwo73YNkdG8e8NZ6VRu/suINXbe
hi3rW8UzkaUw8l41CPboKG3RNWT7Bdn1Oi82ack7qE+/SgD1ioDU5SGRKI1VZ0hb
MWpR5X1BsXljl/Pl9LiM6p2Qq4GoMJqmhaPxA6140tc65sSFUmc4rkeCsKoudxWw
KdpQxvGM5KPaj7bOjx0N6VgGCDBWmsiYF0KU7yhklqhgB6j+qA1VWTTnKD0mdPhm
UCLUO6dUk0DJ11iOqXFvT642yS30D3GEhUvlKl1PQxjr0p2Lwp96/HOw+ICFA1zX
IHxyGjwQ/mbZ1rQUGOpc3Dmh848zAWTmBs6xdGvz3IUPituCSUhS4I8UlOwF+I2d
brAB76HLQSzaUQHdIHYaVp2qjKEPK6eVo6JOEfRqxKjqOM673feF37/RF714mudu
YcdRogzPFBCCnfqYm2uJnbl+Iz0Jg2/LJIyBWtruG78lArRquSA1Kq3N5WllBmEa
fMcOcg9I+TeyX3MAD8crexGZUW7HucmBEHN3plxwL1AqPoqUhseBS+SX0QEkQKxC
cJd9XpWrN8KjwNCIAyIG7XUxYs4nVpaCqOTD8ZV5bsraUWH3jUpJw3Mg2N5wdN36
A5JJbdK+25GU2tiwdCG1urr4CzHXxvwvPf0j+V/A5Ktntn7PZiB2zw648/brQJsV
e64j6HQpIBhfOkymjKYDZ71PYJQYkMU1TMPo3MjoHS4WKqFmy+NY4jih994k6+E+
Q3LbwPu7+e5SzviJ1kGap+XVHSrBMqMkysB8Jx5KaoXkLwnPZoo855UejvQhDKN6
vNJXysc98iSqHKb5G6dtCyxAHaNAYpJOpTppdX+7Yxn/6KJOxq8UgqoRuOjQGwWx
8EaWxgpRcAPEQiPbnWTpCIyU+4dm7vc1UHdV/Kw4Tl3be+dzSfR19/21Uyu4ywHd
2QZmk0Y9vDM1OjfwK66lskqj5+82fd34NW6RvpdKGWHEb76e/Jh5jN8cz0w802Gn
qKR/tdEJY0/hNgptFS5qi4KjP8LjTKnYiHwEvEmV4ayK0m7lDNqNd+tN0mrEniK7
Y8+JgtrdUE11oQhi2mK9bWaQ024wFQqcp8GK4Ms5iJfRr9q53G/xtbXshbfX1LmS
LIR3l1t5V5jgaP0GDH4F9nxRINN+Z67M9Ryg7SyQFlG9Ph6/LFRI6NgArPelKiV8
4yeJwfy8WYdHUu2Dxti0CRTg0ncP1ucWJ0pnf/srCxtMWbZadOUAqnlYcgMyt3qh
vY7aBZrtqkVdOeon0NY54Nz26MzuN4aoAEVezueJxRFayEII9vcTGTWB/q4QQWbx
JJHDOeSgmX/UkdFUBJP2AGM6w5Ip5mfSgs45VrVjqbrrb25+R8CD8jgDf7YZiyyf
EXk+fMnvuo1h7EgSjXgqCzXN9WOd9esjAg9tmjsjSgEl3ljGvT9HI6l2hsZfMdpz
kXibW370ZU3fVpdoxH5Myslc8cmIMpD2R+02w0dS4Xw1OSfuamwikrZHlh40P80D
uqtzvKpooRqSLQVdAhfb+AATCNmIu2yBOmNHcF++T/HQoeU5Zr2IR/jfmvsE0u5+
Imnx4pGAog9PghYrLYc0t5WscTORebocvfOeTS8CUYHHmDeK8YSbVYDxxt3lHF0B
nA1tTQSszrkRpIqPUQHMIioFLdLvscP8qFt2/Faq5R1eIyHbMYvV5ap1ok7OhqhM
1iRQDJBuvkZS969ROe87jOanDmX36KaZUvUEQKBne6cnHll4mQ4n6PPeyEjYlqBN
z1dGPZMH8vzH7h/yPXHq3mln8hdJKwgUORhX9Y8jAqomsCDl/9IT8uCP+seg6SxP
4dA0JB5LSqV0SOcsubJe8lmkwNWM/7xppQ0RqvcFmiKh/066FBboFGIJKU7LYBut
qh82Gk5A6fZI/sT8rCXnsjhvTM26ccpyt6PpgJFLgXpdMo0CHob4Ws1BtQgUgGsE
Kg6ZbOkPWmRPI7BJ6DGSaZGNMjXXZx1C3gzpNXxY+A8rDD9hfSMCKVinwwuqq5YS
9gdMDKZ2fI3VA/D5OL16Uc9aW2nR+E7uMuRuwBg+bZfNzkV96T4Kd/O8CjsbxuiN
DXnq/LYMHfh7DeyaGEyHgb5SBHFAWZkz/H6ClQlveF+rfdWonB7MNx7UVhg2z7AS
lDAeRlP+QohOhk44ld5rtF6rew6wLiEi6ISN3r9RaK2oUt22Vd5xOxaCByOpEgu6
L8ct1hRCjc6l/6eTLcmNPVc0UDznY5oNcmBcSuT+k50qF5tnaprcBQ7BwHlza24T
eAh+WRwHnf5FpguJYdiIw7xMytKTHCl0ceFyxfy6PUq1VULghuBSpCYOKIIFIfpd
8Cdz3WYuETWhVwcKEP5TZHksHPQoP+XuabXLxBUCUZEg+r9M5TfJWWwXVh+qD95X
6W+iInCgkagRfBPoU1v2b5TKCrk1TTUGzta9zXlSclFsFx9E8zNQh40KlfIHFhFX
GktgIJymO3+bZtpaXSZEWzd+jn947dvO6X1UGvmNQE/dneO31GdlYRv/uoOwVveS
Xe2CT3e538lQEl5hLr7NhpQRvq+7W6Ss4WmGD75I/6hgUdd+gCjTh2zSe5aBiJed
2eCP6xTMRfr+nZhT6K48ecpHzIGhu74jIaSu5vG+thFU2SWgFjBHjw+zCK0LfsGO
6co6/RXXC9p34cGodqM7Jg/2HR29rLVcvkS5GLVeonxMteeuvz9Sc3Gq4yj+E+2e
41x1tIR+o914NscsBoWZvQ5QigE0GWpkUY1/vOPxxa5lkwWJ3x5HPDfKBN/OL61j
DerXA4OaoH9rOolNMT1I51ixuXVFQ3mz2G12L6V+FA98fOZXEgOja9wgCDrtgqRM
mmD0/gRx55uirpxcqdqb46UrP7cdA9FBoETdhB45bbkiqhS/rc3YFkuGyuK1FNDG
uXNEXWCwg2MVyIsBp0ISi3VEHvaroJ6O8GwYvxeqrojxmiJQF5R28KxOuJfRTm7g
63N781c7msYpSBklVeeNWhFuxkB5rkB88rsqTUHeT6c6Dt8q0n0ROxsFI185yxLS
OhvEk5QTkmIcl8yLBvDWspdp0RjqkxCId4oAv7xeryvchlEP+vq1T+OUNSaOvHJp
/bLwLaRV3hsgnSXWp8uMAId1Qk9mD4a7ACUOD01jkBotL5IW6MM/eStu8d+f1Q76
H5V6/K2XLCcRl7k/Ao7sPprEKVjzdRFbFbFLmZPloKnjH+yj696UZ+tCVFab3w36
fJ7+If7VBTfPTYYkZEiuWE7PeTKd5dODLewSJqpQY8uvA0lSjz55R3Pns9B9C/62
AEMQZjVlu7RpDxRtgw7IZahJ0ZllfdcfGLuxsjC70gp0WiMTuac5UpyDI0sb5/Lx
jnClm/o2cHBGfGdRubArHdTQOQ+hlfHe5vtjbDDZeAtHM/clU6OEu/nELx6Jugbb
oU3lOlcKJFkpN/E9YjrgML2wfB5TTrfDE1YWsYlYXSgSF3/YhyngidL8CAgPeVPN
lFunUF6jz2FaJ62kQJ2cVuT4pu0hNHJAQB7vXqXL6vKsIk7dEYF5xYUL/khB9+gH
zBBk4TX1vGe2mZq2D+MAksUCKCz9vZtsyfreFTtrHYBt9wxalgBmo+T88t3IW0OT
2HKQ2JkB1zV7b8WFw6HG1No3dKsHppLLTrjRd6+53zlgsGr0roqkmlGVg9aT5NP2
wiYKtEQvKQwbFIwUVjHlLpgONFGc6c6vTkqoJ9iNwGOja+zjMifM1yHtbwMlQulN
YXMmKkzomi3Ob9Fw+WM0aB8UcfctuJozzrsjPzOJJ0xKiojAVH55OUab3DEuTBzH
5GziMO3hGXl2UGt2btRWjrHj1p7JDH65C7C5BLUHM896NRSTqfBc7G9I3AmRbNBI
AYdD/Xsu2boi2/y60GW6m4QaKQ1pq42RQT/68Ixmw3tPyNr/jHOZzLrTVAthY90F
Ma3+WwRP+L3fPjtXcdVgbxkShM+VvsrOXN2gxpdrP217qDtZ82fLKwAg4YISJo2H
yeHRM+FQCG9k6WWQSDpdv2S6yfRFiA1ECcLth1Tee7oLx5NC4QkGd66j5LMMBHai
9tA9dia/c63dPftGZekNhpnwO+Z1oCP5Qb3u9h/BfxDrUbE/C1CSsry97q0d7OJg
cwQ8jX4g4ZddXaTSUcAUcFo0xfvwOl4ycySriT7wFTEaPweh09T3BNJRJ9vdhndY
vgkZhFjqyQumR7fLGJitrnPUBReRuA/4u/thJ7rBZLhlBXSAEh2mzSpxSKEjewoK
CiE1MNjgzQRBJxCMANZUhsMQlH4PSfed9E0pMby35Wj5B7p6W15i+FKcgW0MrM5y
3JJBhMUm2eWB3jjR0oOKI4UVnOhBJr6/HXrb5uoGVudD298+umDJcriX5P9BBkqg
xUYKRpg1zaKrFgIdTkwVkROW9fXdiduYSf/bSUoqJQqcxD0EQbp1NtK0gp/xNeef
/9bEOmmxMLE978x9xAqlmCsIekUBZo4gy4tLj29L9iV0qb3ZmPvxzaWt71qiKrxw
Pq+TLj7EKf91Qf62vRQYveqiIFCAtrauGY2m+RNgDH/l+s0v7oHd1iTPK/hWgeBR
aAqtSyJwS0kHmPR5lULo6a8++PTg1sFf3V/VwUM1QqJ09bALvr9jrU1kGXp6ukta
bOF8IFB0HAxycmFgOKFjYmmclryhL/Js8R3cocimBv34LINjiI/SAlhgDv7IChFY
x6p20l/gr3jr2f9WFdBYMlki+95C2kQpzISB0Upmhg8jGken5oUrD+RX6/jvBJei
BSx+uiIbU1qaHdJNmmKT/Sb0oM+DZu5E1sboqmmd52q3F+rXd1X5DtwwOBStsIQJ
oYPugqG9xWhi6zp2AmnWlnYaIiidu+NckHHEFWiWgJOLhQuAXa3XlJRCz/LIPAE9
mxHQTRTCIr7kbPjRuf/HM2HR1LHClyRe7mKAIaw/witMlWi8HFrod/3IJpRpPFGc
Aj3Tym2ZQtwHsS6kobb8k4q36EhrnhjtDB+XylHz0taR/x/T0s94miOHuuLjYIuz
aGw6Afr2l2dZeWixF7qETirTSjHFJwDGKY8e9ZWIXr2DKj7kM445D3YBBsxXis2H
GgcJ1laq9+ddAtOhb4xlNbIeSdZu2g6sw6LwF9PVj/aK7EPXdh+ONneiQ18mieKG
xAkHb2bPqLbpSsslGPcoxdHlLQxe46r9ABb+IpgdrHnwVFRImSibLrwD8Esgu+j4
7+xxLYixEc3LjrwN8nBy1A/T3MRNtkhjTDw/JF77PMzKurJGAa+3Z224Lb2GU6Vp
ICKv8LSo5IRFzrCq9IGEOoWFcn9lGZ1BtCOOsxCCGEDpgxR0tjruhZwI4Zisf4Qh
4uqpygsJx1S43tQPMgVC4RnIonyShZfUllYMauykyzv3TtzG8HWFVg6Lf6Q+kb/y
1DXjgIcnsVFRV/A61Se+elP+3Z6o18znEuBjzITtVeYvsllA8Vats/5tWFMqvPiE
IUVAqXILk36LZa6REA+a+U5b/xatyvWT9Wq9gHXCgC+iz0WXk0PHtuuTHNpgt+h1
0L6CTOATMccl8Ycr4b+eJe6E4EA0WWavLU8DMH5quY9xBtDeFV+uVZdZTSb1un4X
cBqQscA7qRJniHXt0OuhiBv7Juz7MjSKZYntBpzD8Mdq8HmJaZqQYy/aoiqrFvkp
HX+CKfN+x98T0SEXry44P4sZofmsTOLS9L1f/nu3o1TmnCQl4TG5l5v7S0mt6tmV
CbZ9MXLKb1Z3xpHVLN+KH3nzjWb/YKd7YE/hDI4iDuz4s2l4FlrsRML18n0T9PRh
JlwLttWhhX2EZDjevdPuIkNsmOEjBCo7KtrCtOvGGiKPaODt6rpY2YVSRdUVbFdt
+Dx/xhy1xUZO+P4Ahpg/5iMAvbFTxYUapf7mDvxRUJzPmk2e4gVb5WoUjobFCFAN
ot2KCJ1OTasUDFTuLow7H/iaVIwU9nV2Ce63y93HFCabhLzG+JfAid43NLyc/S/I
W9XV0q50xoTo82+V++fZpgWEcBW22u5RUUzOUQZcXHufNeXcI8fc4WE1FjTOclal
UrV6g9iuFZGhxasJ0f5FNWWwHtEfHBVlIqVvzagxcVBbXNLTqfnxS/BH4it6YgD9
oGtgv+B/tT9UgcxdgrSdzJcK0JJEfLMMLqutsuTzqtZamxzWUzjcmduBoKy2S3hx
KWZdik77+w5W+xJ42pgtKiMUOvAQv897J5dv3c31P/kAB1kyboKRuqFaHi/ymNbk
P8COalhqBI/0ZCjAJM4yLCJ/OEmD3kJh7x0/McgDDowBH+gH2QA2dYWQ0asOT7qp
KSP9E2vQdarzbvmeLeAVFOGBsjcgr+8SSWsi+myWO6ON8to5erKieCe3gF4/OBzx
tPUJAmmwdsknSNFJT7iyL24fTWr+YrNmr8LWXuicQPX0QxRUSI6QiK4M4cbgJtM4
zPD55Kj5abbVPn5GIXW1WumCTXS09vUmohCUp4+iagk8lVWDtntVzeYuJIPZMfYZ
ExXKNKlmAqmn5uJCWO/xxSVX/IbwU7jf5bBwrloZW0hQm80EewPt3mbe4enuvnsM
XdAbPsbVEGfPVJanxyP/t+tiKuStfaAiHn8qAO6UCbVjK0LblYdLS5Q6gR5IFpap
UuSp/s/072vUA6IK6y+FlSzZv3dUvQGUtOVkaaEZtlKu78D+Iut7rcOu0AhZQW6g
gCWXY/fqRMg+dNlFjqnWW2YYEGpFcr/o5SENnziZ7hsmJ9U+heOj3JaUL4C4w1g1
hBOur9bUONoAyjmC/idUBlCFaJXld81rhyCgNP/M9KjrXrKC7gUzKXsChpDSRS+O
bE/7bi/P4UmmhaHCSKvAUylcaqBiHpUw7cO8i1mA+0EhB76yP/MJwT9QAyQ/783z
eH0OpBiyG4pgFIDRO9z7ca/s2Vdg89TKCBEmuVgmKCj2QlXzPeMLB7kku/KjucdS
o0b28ni33RQiiN5iFGr7noVWP99J3Aq1Flbhk4111MrtPcx1fapoGTj+z0acx0vz
VrlFrIJDiZzHPmwHlmYYfyfJBaYKSezrpjoAhJCTB5VefWjhuTfrtRGTgBqZhi0F
3lBmgkCkie8A7ouLTWt573xBA1TkYtzentKWJhKlyPTqGgq9rES4W9g20zzpRcGi
r7NEs8Jkut5DjSYquXOAr10E+o0He3ND8ki27aEhB3PGSBGlkVb97YKpcJQAkU20
Ho0Ea74w8Xu6uNbJLwAUJqhXNrMBoIQhepGMih9b6wuW9t2bB+VVXkMAShlKCo4U
+ytnPx8Ik7jEm+bV/uHBev7nlo8jVtJmJn/avIY0DrgDPYIQ4RO5T7H7MRKeMIJZ
YoFt96razp76idTpGs4vntijuu8q9i2zMS0kvwhSr06pNYEQwenpuMpTq2PCAMnC
WUIr3aaQfBxA+WyCDDRBpEMPeKI+Dnze8N8YqrSLjhPPvj+I5jHw2QOUz00Cqnko
N6HaP1sId+ZYeAkRVA3KjOJWc6H0DprACrrHVlJc2jVXfE5IO0z3VnxfZ4apIvZS
Xm9cZQXRejHuxmcaBAe75XaQWfAKFZmzKytD7Q+a8gkcwhIXYsMUTI6IufW8YTdt
1Mk5kKZ7gvJWTwE9KGsV45Ta9QPCGLQNlWSt0fRxtU8eqYVLCm9dO65k/Dgf43ns
7Qjzfp9AgpgmsO/0n7DPJT5jgGf8PN+UXUx4Y2sSlDWxsNheJkf+UTcVjerr2pE2
mA0fEzl4o9roY7odLnAmV/6np8MgS1+br2sg9FqfXH8N3ZpOhgWVl0PFhIDadyO9
ogdWu266NtSvoXJ+TDg4PeccMjDI80jLSFuDZATuZ0juMrBg7+o0bxNnYutLE0bv
E7QLbmkiXlqcxzKhfx5XHPbrDu/ZwbVZPLMlg8gAFFa/qCi26FiTTBDFsXE0zPSH
6iltrkG2KzcFzi+hGz9z5Twh33WYigo3WOzIhrcpzpWBidROHnJHwxr5tVNj6ke6
tRIBt4ZLu6+4zhz/DNe5VvqwcDv7aTcGsgYUHfCr+FXwmCtUoo4qCevlLRb1589M
G5XXcjxP+CJQYbnZXKe6G0I7Vo64SROl2Igxv1I7aIqc5hXXPIZ3YojS5D9lmb1u
40uau168HPS0FVXcvPgDTkjuZgrTK77OUf3GRrnW7GV+3kGPD6TaNgGeNKtEzqdW
ypt7w2jtQUDicxPgkHKgwqiDHyxaIB4BhOoeYtZMPmI1ONlgdJLSVd8HMoUQXHFp
tcFU7orpqXd34KFwIdO0gENCxpM6B5zI/15gTkspPrAJuX5G5lL8Vnyig+JAXsrG
n34aC8GEdz09eZVksr2gOiDzswFX3/pcifKjhGpA4Wuqa3mjtHqhsjH6u5sIQfz0
INZOEFcU2n6i3rp8Btm7uecOMGzW8SaVHrxTUZ71ERVCG4fMvCC06VNFI2U1PBJ3
hKoeyRBpIBSW3tCLzpfdmgpQSNZcTRkL/J/A/nFsa0aoCbzrD3QqqYOjGvWj9e+E
+E3O6DrneO4XFXjGBhuVXM0F3fGPT8c9HQ3R06Im7csx0teJckSfdEyH9ZRoE3PW
braJ5jI7+JvysiJmlKOaZJNqzMSNH/pSJ2V8qXYTJvMQAlc1K8wtvZueAgUDIVKq
m8OLfctF/T8lG6J4CiGNwvSNJAUP6CrJqxzHctd02IAVIeVrn2WU3QX4+YFCJoSl
FvA9gsspJ+l2BDwrMo9HDyDzd+JDrnlk9lBo1N/zWarvsyYytnNu1Mh0isD4LPjp
KMNJq0dPqJ2Qw55j8tCrlRySU5iAgxLnhueUQxA0wf0oIPn0QbRrde/QfZaeovzM
g+CnUi34vHLktnPLtOWYvU1YYmiT52oPKsVhSdgmR5Tekktm0oEc2Rmq17KJOxXc
R1/vSXKSWwEZQbxFfjKGTCpgQkcJpA3Z4TM8abu2fqY9mO/TXajqlTsIxVSGF3+6
E7d2fDdlb++U94YQOygjZGkKeMZuRhzFcSdrWN8A8qvOrkbkKkWLTpRWpUO1GN8E
VmtdQHtlOF/f0L5BT82Z9tF+C8ZCxTOqxH57E0TD0a/U6tu3nJqZs4y7eFDsWtCQ
VkL/4CdRGoMLN55cmrCJMNP5zg/jB7WvmVyddxKKbjRcHb3COCEKLlO4vbYb6Hw/
IVHqg+DJCNwrnvIfw6KVpTPP4Gh0zb07DnJ1oLB2J7DqhXoiigPX1pAqh1UUEpUr
bJxfFiI2cd195VsJPSv3fNpQEfdtjgMDLJ/Nvi2v1F7NuQw3CLz29Lk+3EvklSyv
yIO5NK6Xgrp1USyQGUJzDh9E6ZxuBOtjj2OUFANLVIJJXvLpYO/nH/ur3NwTw13p
ZaHL2kf+PquUzOmTTShC9SlOLlypqMjEAWqzqHXq6N35TFHRVDF2j5tVmEmiU0DG
q7H6X8XbCTUIz7oGrVGB2dyccO+PV7eUCpxCmiswbXH8feSgEx8cXpML4AyalyAP
J2jqEtbpqXZMMHrKVjqP8iwN9oweetLvgDgf4YkTDTOi4Tjfr8MA1T5q7aW9qGv/
7bo1L7nsz8RYs0Z9CzCoAib29MEVMnjZ3iChppA/LXRrnMZ4YuOseuO4lg35O8dc
GQkp8R71n4u1HD5bWVHKvtsBpElfplTnHylwKVTKXNWgxwv4TvIq5xVo3beoWXlp
AWTNhGb0c+qoRQzGiLeLr7Ss6zhqFgKV58CMJJkrJYMRSy+ybIlN0tpzrDeffrLG
JY389lUMuu7bv6E/llSG8x6mWOxugVyotQ4mRivwj6utkvsWuUYBc28hEQRx79tB
yyk/+8YBAUzOevStXzcy1/ffew0FogwkEPTr+oQaAmnHX6s6e72JiTcB4D8y/Dot
OYj6cGdG/FqO6Xn6rHJPSRg+ujce9vhpdcqzacYu4rkX9ML0EFqCTnfGUezgVNfG
0tPDMDFguTRYoyQN72ejCyZX+p2u3JlzRlmgFFaKvNctWky1W7UzJNt3TYM1xu/d
sEAi8xj+buAwe7TATfYUsa83ycy8yhy3HoafvN+V7kAGf3holyRSvHcDr0PxBHgD
ahDMLq47CQoNGklr5A03qkk2h1X8+SS4DNlkQLWVOsI7S9r8bqIpTVBEpJmK1M1b
GjcrEdtIPitUcTE57eTOZaLQ4v9LNewlBfG2ky4XtY44oHXu5Sq9BFHu7X03kXiP
O/75yW+0oeliVQcqnqG0ZajiCnv/NEr0BJHsCzaP4uPzge7b/7tMntS4Rrr8vE07
c7jX4qhaTTo9TJOCiUmdcsdCAPhFH0I/FcQPmqsbwN8yxanRIT1KLq9SNz9LpxsE
ZekL/FkynZfcfdSsXLTa1+CFYXILPlR3PBFc2wJsi7VGzDOTNn1BLEhE//YjsGZL
ScIX2TjW5seyn9A8PBCxpc4hOw17cRKsd3Eu+Po9nlpMCpnxHL/CfDRBTHwZfO8A
yoZO4KK/TwXhaGIJpVAqyBX1+PjoVLe7kgIeqG6siXhrGbx8kiMGuTW4a2hHKEws
NY3+Oj+Q9HRGLxYesIxEHpO/IRI1I++6gu7J7qpo00g8SpyIykqKAOhSZLRNnFS3
9AIEpAnIJth702IL47uqHMqMRnEljMd6czBbmSm2rJPusZ+pDq6pJB4X1YMFq4q7
R/ceZ0hgtOrsvVhnafpyB0Aefmj9rUfU9EYWgRdliAha2LnWxiChfjC967KZ+eHG
5kxX1Ef/YzUBTOpyBrMaSlltK0YJ53Fgsl4j60MwA634p31BhoXfYlDbqP+dhNM1
xu2MB6y4Ht3/MoHCS3hxRb8iQy6+TRWMMEha/Lh3VjLxhANyCIUGujP+u7uneeR0
LGb1Ivd6fipMaDmNWg2q1GfZjSTxLbdrOPbAPRCqQOVxJOfwzeCizUanT6j8b4s7
Q42Oj3wdhzVfw5j1SWJSbXyMtvI9aJi6DPPWKoCP7rjfY41piOcdPywMS07dnOtz
3OhiZk3tps/jJ2YR8xCmjZ1AU5X+rOhtOVcP9c1p+IQt/CVdWnbCQr52+cHQy652
zE5vH0sD02gI0sBlCVwl/1e2HLEuNhOtjoI1c16bh6B1kCH6leomrqHUTKzsQulY
4d6ZTWQ+O9XraZHydyoh93zhbqZ3voosuEuZHCqYZu4fovfN7Pgk+0fndbv6Bgoe
AABsfaSG0SEhuL4lP1+LR6tduKKK053X6WcbOBE4Kn420ZDPR4+ZTudn5VYywDxz
ufRoJplaeCmg/kTo6V7R0cpAhmxx+Cxhm/ET2BzE0kdR2sVeGNL/qQ2r1GUFCIxw
7AAiv4FfX47/m3BQZNqiCJH9H6PaGnf9LAWYXW7enCRpWtZBxrBXIzrAFIzFeIHO
0zkA2ssh1CjyWJNBvY6HqRGlc5MbZ7AU45NvrzCzOVZIos6BhsSknGzgDACyzLZv
UTZhMlzSApZDPuAydF788Np5hFuG3O8pVuaa8Zwcdw+PJxdBLO/gzK49nH03I9UJ
7SOnW5WMXGCfnq02GFHzoRg8J72f1ss/MVaFleIHLvSdX0fUDN4eXEP8Mezr/xKe
wJU0QG9SispB44hea5BTRluTfDK9QB0qmB9ULgK395OLFQ3vGVWYsfR/e9TH6xWc
5cBRjy0F67ZG2xxfJCJZ9OxsuGBeHqYdOmMbhWx2rZPyHUQ63Wb1FtPzuKUTeNVi
U6a+l13Lbjk3t/XzEj2s9qzhUwgnnfik9UYB1FuaepK/vj+2nuoFivdi+03UVrWR
ga9N2Bv9zLvRLZ0MfxYPk50+o794bO3y2Zxduydz85FA4T7wJ298kb0nl3af+w77
LWojRO9Dre8B6PDPR241lN6Py0QYDdkRtWbUFC19eEB4CGg7nc8xUWWEIu9mX3nk
4YSVzrsItl7YA7Bx7fYhHTVmqdE5u7JNwt/VkRJB1I/RIJCAG/AzT9yRM4pqN36c
sqlLk50QwSfHU4eol3/jGI2Z7we7FxyMM9AOHtUbHq1roFNPFw71PnM344oUc4Az
oDPFW43IQz3fV4eY9h3c2VXx0bqvTo3DZssQWQczceCD2depmPZYPRM3+sAw960G
/oFE2LTg2Zk3kj2PvsrS4B2ebzgj+czKMxTAuYE3Nivk1nzW1eDxu/K0hPHIbK4Z
awuV+39PnQyFtFtxHd5J9M3n7swAni1tVAXXOk0r5UpoLZ7xAoXk0hKIczEf0IcP
5q8t/sFwiCsZ1W8rbnOQqaOsotG3urDP/D842aZAoN+ULHYwFrPMfvjbUgo5gW8A
JHusAT5DZBdoj4dbrL0P4dBVUa2nYlk7PLIzi2xpkm7XEs0wv/5u6onTL4W0vrKZ
7cEnen5VsO+KEw/RJbS1zceKFzrQbv/P355uFoZbAfBdlaP0JpbqXmMUmGGl5Na2
Ygxi2CEpUR4HBKJb/g9imuQkOQWDKz08jkp+UuRrhjgvy+B0jZBLS8PVOIEXCGtl
6qZVRocSObaY7Yocwvf67Jg3eCc6l7lhRj6uVOa3XvCcHLlCTQExdBEfEn2MUZxz
1+lADtBwZNfCunVVC9zzL0zsD8TSI5UQBImGPQw7cMzGhq7X5Xq99DD4lwdHNe8C
qQLo+krms8exyASDBpffZyWN5cIs35fU/mytu0RtzvIB0A+di8biD8JjUEHm+08U
DJcof+KaeAIrIxksnRJDq7bF68d0lHSNUhWToPCIKZv8BOQsj1+PkMoIeFvMApyA
Gfb5ow1bDOXEQ/x5ADxoGyKDsyKtZCHxUE+hJgK5t3uGhG0TrxiRZ37Mouai2PEv
2ivZu5Jm5JAw5T38J5x6pjt/C0M8v4asiz6xT7CHjfvC/j65xNhmdFVuRcruhVt2
mDvSoqE4vDtDNvojPOCTyjxkS/MbEpVCAsnTiu6ZdttFELBW4Z7uZgq1OgaRoL6d
MF1PCm0Jc8rmLE3Ty+TshqlqFgagbjNh4iXi7Ass9B6utIURjyejZkkaEF4VPMz2
OI37lXn13aYrbVEM1BCJoYWJWoOgJV/NCAvvJZH92TF4pKCAORgaYqd9FuHpOAl0
jHBmw3d2UUtIITJhb4jB+Utzi4Dv0vqipIajT0GtTfpftaz9OicSiOKBuchKOWuz
FcfJ9tw1dVH3v3GuEK3vVs2SsYTv6ilnIexZ6kCJVyxbhEZOfNWKgDsE9fb63+fL
Velqgn7JUDhysr29wu+W1eYZADGQI6/+ztWBjy/nRpiFfVUNvnada3INssheDBkD
k0hwZzbF8w/EuT9a5sDc3mi5gZtai75vcf9wxcuspcjojYkVRz6qYgahqiuKDhOY
t8a2kHgSXZ0RorQO7O9vgKFhIIWYnAo14vbGA83jCx8WEWbFFfS4SGqg3wst/yMQ
g5jLQwmSr/tqsHE//y+Gr+mZz4ub0M30tDaodri8NsDsMQNKDFJMvm7PdZYctORa
8Of8d+6hswWT9A0JsuIs1ltN+X79XP617NnUX7iVkQzdXIRH2XPDqRsXls+W+NXO
6YhaBeOOQLqGsLhC5U9ttrKAwW9ysNyKMceHo1BVxki/TWidP+88WVCZ7xv+qVMm
5TkJvg2G4uDUXTfs+cdd1JqEPCV8AGvXX+f6yV6CymLCLqc5IoCViTHuuZbYsHdp
sj3c8c3QR7CaCU+sjCwvB++1salXMjy19k8kEvG3MpSa4Lz/FSVbqp/RjbR1BOiL
srTRcSwrMt9NX7yLyn9TRnccUkFcdn6KRMcDKO78czT//Zi1lkEQkQhIU8tHz5gv
JSy1le4zWKFD7/HYiEqL1FsmOf70/juPxKh81kQtHCvPluexVzxuY5oSf1896ZBC
ndM4fQXWOW/7U6HDWfGSN7Qk7pNpYmiMgEj46Bb8Lvr52f8zKKBZD9mtxr+xNuCI
TLMQcFt68mvjsBNdC8lIrN5326Z6CwPa+U6Xo4Pki96JfBFNeM1dZNM6EmB/E7Nj
pXlxircuCy6dKfRbpIquDSxsiQR6qKiJ809ZPDv3t2IpW/20RfS+K4MgXuIzcz/8
hR0D4fbv82lq4xf+2sRu8vL50OyUObmyaZtjIg+00ubM6e0hCjzZKBQ2AnK+iWWC
SG8H6CpCR9t6DBboWV9SBlHCOWQmOc3Jb/RCb8aFgBOHWpaQdfd7oxiRWd8TueJU
1R9ZiU2bm1ae8LayG1qFCNrH+bizEQh6KglpbsuPjkavBfaYtKyWACScdpBMK15e
UvUcMvWm9bgrIBzeFGXl44YD+tWUJLDOCn+3KymW09pLS1j/rMhs7fWqU11XFLAE
cpL9Y4pZeS6N8Ks0F2u9KUFXxWvzptc5IYWNUQKBlWgYwpk3qv4FeCNlpFewHPEO
jfp4ZVFqmGoBH9NfUUc6x6VqQ0W67RHhetZk9Sl9kxeZ9doUJfdDnuBaUcbPHZ2A
KaRZeX9NlGyTOi+NAD95pSiMbtB35M+Uq/mMtV0KsrbUJG1uf0yPmPuPaoF/Vgre
/th1rvHb7jVMnmtR76LW0bu36oYf+o5AO7zh1IOVnUATZ4OGgwYJJBFZjt4+Yzqu
cmBb5dAqLRdfAfdgKp8lDb8e0zPydyWwPybmOhiZmJ7FTLs2wNoTIYx84JTrh1QD
IhdyKtlXu2zLoplYVlPRTJY3RegAIcbWZpUpcHhIIt/r1Li3m/t8zl+Dwui+bS+2
VZi88EOucOAmr/yHP65CUPAQgIjVyySMZubgfSXVvDFfkGRzNBzgmZIHsAq+sygy
ynvPLB8Zjne9c1hDRqS80PSS9CbY6e6BzqagTdYpcWqEbVXWAwU1J+jjF9zs2g+n
Dcx8zp53IXT5Pan3c6vUnCWMUhRcJLU5zm067zeEtWoL3K/6zCkwa4l8PXJVaTAh
vDuefm/w7yOLnyUwn9Qu8tu5lWsV5XfnHp73UJ0fb4aNIyrLp2hku2qnhfQzhq2h
yuUl8Flt+LYCasMmeM2WWeemDARSVC6+jRrHUfDiqH5v05FBh+18F2ocA+sTEBfB
M17S9xJF1tYRyFJ87xiprzA1BZC+lfITSKCneN/7YqRnhQwQeFLDO8RGI7lKrEBy
ZTuowBKaQwO66Sca7QtMnTRfXai8pSwZScC1qwTXGQX8WO3srEYEYStRk/tw/bWy
rMvSAdfTwV8WGmp/8E8/KlFyGw1cCs8uro6aYYSD/IQ/UUngAwLRX5x4ugnx98Fv
82WaC6UpSTv9BRqLuXY7cYOU8LzF5FmZfigZlR+oHnsHcI1WoEL4FhJkcx7p7Kwa
G3xNix1hkxJI0IZBN6746T7lkBSJXxNtmxqPWdJl+KKDl6Tnb8TQ9k7cmNdGdna6
SW7K63mluFbWqJG13+WckqZYATHJbsuL/fQYTsj3g+XdSjTVzJWN2PJmP7VNFnch
Z0Mi+LwyrjDV+HRAghj9d28tlOtgJnkT4FPcrxrsa7fScBfm3oHSso3V8485rIkX
tR1HjhjJI9R9glaZ2zU/2miDw56d1LErn7Ck0VKoZfVMQEO0Skmo8lymxrs76Id+
zwh2TmyG0YGNuBrbncjppjzd7LNnRXmySw1Z9hLMM2XTnDfFNAev2BjekF0L43Pe
pi1TQCHcbyowFjyGYgqQV6JANdIlHMMCPtFt7Y3QNkFSfNeZzdviomo0bB4TdqgC
nwet5G1Wm310NN2ZpCMPkpHwtJAcRovqHUEaiQXRber1rUk2b2I3BJodadLvbZfd
LybKDLPWP2oPzt826QZCxwkTOxMrfuGFWVswtieEBhB48wgK4Ju+VLUYtsZ2CQ8c
9P8aVhDzosgobHgJHawzlkGqXAQfrwC3+yzSDOT02Vjz/zPLU7fhWSR8489zYnAv
4Ix4KitW0CewnjYVF5K+23vkkdf5egha9At7qFp7anA7dgvz7bR7YIpP/pbKCfxF
WAgnTMjZgK7/lQ+KQ0ijKXZviu5v475asueYdf/brr++kI6T2Q0BnxN7PBst94MK
+ur4oPSqdAXuMDq5iXC+OaQ69kHKvn9nR3XgXLTYOwf+Jh1xC8TEFm5q7z4xGBVE
ON/0/PHvPGaUfNS5wA2b113ww5RPZ4otGtW6A9C19BGiOSvVfDdjivVkcp6ltMoI
k8pt9MNWKWqo7i+alC/3DJbRC1UnTJ5c08g4GYU6BenvAiQ9vIY19AM9nC7K+B9H
n6cZlPtS6p3+qHYaL90ghQ3K/gurPFGK1/gMiauo5kKp1A+XR/IiLesNmvmaMmLa
UCRs5U/3MT+MhJNVrFVkhlYh2qFW+jeVdz5Soe/04JHGVML+dqACxWxlDmS0jc3G
c9OyZICns8ozKLDuDtD1S6E0F+urFYH64qL2Xk9pc/Azc2b8xuWuMla9CWbQFm6Q
0cmuQmjF7Bc9gDQPK67Vju0XfEnacpE+l5gLeJph/bu1um54dAp9uuXz3QTpHOpC
MvGv7FX95XqGNx0WaQS64Xh9qLoQQC2K9vgNZ//gntX61UDkEWwctgK3Kgs6esfr
poZxA68NL+B3d13ji0fDry8eOKVWPsTODJkY2fqdQ7A9Xv16mezZZ4lyr708GlkY
knOJqQSiPguGY7VfdFfXojlVbIx+Bsk8t1U+FAdvKjUpkw4WVSHcK2KJ9omrpIAK
FtApEiky4QXOrd8bqBZYeVwExjIL1OlZTLy2WmYK32yeinADxIZYb8g4s/MWHOLz
G25VRKW0LCeSwFZhLQVQwvfxcokQEqcWmSR5RvvM6+e/2h9QaYBep+eud9FfO+wE
jiyPXQzm9wJ7jujJlwqlaDlhH1grm/7291U9ocRUFy3xRmYJ47cAtaaUi2swdfih
non6ekAzGW97gbZ6A+6K/Fw2nH+qNKUYFLUud7LqqmkOvATN7luf+Zk1Aeb5xdEa
F6nyjMcen7f1vqeY32URfa+mI+raqM9GewGLH0xT35ZvZ+ZV2l+/C1PdMC9koLhy
6bIToH7WjanNKuWWetlVJtFt9jmXPZIiTPLP2cuClx4Nr2a5/QZmWK+qIepXvDPH
CcQ8VEI/lYehWp2BN+QfAfG1UaxDu0xbJKPdwL5XamNCRzg71YqG5MiYNdG6r9nM
GxeXi+9z8MbsXt4p/yncz5bC+d0NXRG1Qt4TuA9/Hh4kQNlyqmFFGHdHybA/024M
CQXFZZUD6yik9uWYZQem2ZneoJ//8gAQoVz2jJaz7ZSStcfLe7MY/ZrlWgJV+G6c
nbH06zyBP3df1Y62QW0OapC9V2rmHzpJezmEuQmVWVNRILZlYZpckIsfp7DGN9mO
g6SId+SF561ElHnqIMXsDpNdiKPo/vUIO8CZaOddPJyce/kLUXb1cjNAhJgMnani
rDVlyRzNc+E3bS9IRWR1jjOPukt3pkm+4iGFWXo8Aj0V4FjVN43yyjbaRqr6bFp4
2YSTVkY/gk+htAY4OfIrwZ4zo165eB1QSjV/ikVWT3Xw4BXmcxnbu/N7fHVZNWbP
qqhRaCDZbxiYMVmC32SYtPrTxd+2bU+8Tbckw86YCtevb4Vr6Eyzq7aSDvpKvgz6
vHUrwNvedu1TpuaJj8FLbEVZAuMN+RT5vxvEK7sLsgDd3MGhXrlccZWdVHjLNzpI
2pkcfqg2yGx5+avTPdxfQDfWqc+vkNoWWgcOmyd6ZbEU2HLVAgSZsaiN99j2n64h
wAsl/Rgv0gwjqg/Ott5Te428d78dgQCeMz0/W3t7U6kt0v98CycezbpeN8mfTR7A
Sz61cNMFhgr7kZoxex7S8pEtMLCrvVylASOtJWijqE7c0SlCsEMreiYlpjs6pWlt
VXl4w2i7YHTn01GMjE7rpZFKHW4Wvj3isEkhefq7gEvJ7xIk6Q8P5zYiSlgDvA1Y
xV+1iMfmC+ITVdPM/DyeCWbwayfEp7wreS91Q+y1GfibeNhjEg7+T19bkV6mxKlY
sMs2Fv8d9vpU5syXv9PD83s3aArn7ySHmV++9RDAOGmmHj6xapU1m8yWBnwNzjUb
hC/+8aX7BtvCrOlDuxDRrfbUCr1yjnVfvFPJWxOSpxg9RVnbzsPdrnfaRtpburpo
XzYNSmzJlBLKBz5luWzRifplp7gJ33/Zs+qE2KiPlt8+/lP+dESArqxJP7W2V8UR
MGqTdfEEyzGbNEHOY4aVl/elWqSYOBScPi9lXuWL6xBpGXwplq/D7nOPY5BdIGIp
MeCSjT1NbWQyVzZNkIqc+194+zoTX+uP2N5S/4dEGqR3lKvr4QP+Necr3EK9racy
vkWMYuNhuo5hCSWAm5HPWL6UL0G1qJDTKiHPunYhrrc2Jf4w9pHKbi7KaiZiApug
Zgeki+X2bnbezMLyV4xs5KSpiIxco07xWj0RZuzlxLC8xeMCFT1IDXSM1PMkNbt0
9bD9aVvoWaIi3C939QnzlADGdssHWy/kFMlijF92HIfBTeczRG3mFuRajDLXZNwd
scfR5cKsm5oyUdnyqbo9dMhSkGTg/3Fvr0EE+WZof1AvjOs4k95fw82LseisGutI
Z1JSW8ajZ58ZGPM9Dwszb52Ehs6JjykfppjktWPRGESxxdVgmvHYTzdSAe2OxUgK
LDLVQ3emu8r/zUoSiQ94OSuyriWSZJxUBf5UV2ZSVlzVNg5JDVzyhTxXmQVVCZY7
UDM/X5BvYAnE32OvJ/ed+pt2UWjRVb4GkmaRKwC27ijF3W1j7qwI4wFbMaS4xcin
1fxi7tcsmArSMjVdMcPHTlmWalqO2D9uhpXeiSB3TjKYM9mb6AuTnnjdIW9hwo+/
89/cifguauzOr+H5fPCy4x4QsS5wPK0IJB1kua3z6sDE5NMIi4UFX1Ku5vBa8iTQ
D9Sp5P7Djfad8ypDCd38OgqSpoPUwgOSHueBTwEgkfkNXkyiyD1NZi7jUDFjdmJL
FJYV2gBvFxwmzqCUBR/obqLAX49LKpBNOWatXPdlbVkKK3bmSTf8uQNFq6SxKFr2
hvO3tfRha+5agGfWd19D2BPGTml0rbztWq/cAFiPJYRQqMM6xYD+Jw7qh+lR72wc
F2uedi0nBDIjvZ7MSTANGVlH4jss0i/k9RejLdddyGMYBwIIz9UV5K8a3QivkJgH
cU8NkZCz5BgrnartY0Np2iXBg5AObde0g4OdYSYhO5S6KpYPEnMdGFrGjF+GhEHh
D2iTSyP9B3fma4RYHDtYEXzdmVvmDpDEQ9Gqf8spWx/78u+K5pr8F9tKgcwLLvVO
SqoeuvOcy5MgY+vbpMUFkiuez7MEvnfLpZ4C0rL/9mfhbevxapFwa1sEHTXHoLyc
Qz6wme3GNLqeJmO09oGLi5VnZw4jtlpdqmDw/cXKghWJWMMkyLDgFS9OEl+TREMa
ckHxPNUEqhv1Zv1xmLat8YXGBM8MmAan8WXvlBBDoTpnWZBSW/qOl6J92NKzP/4k
vDZXD2SPyGUvbggsTwxGghhr4/3pj6i2BaZVS0/De1v+COtqEYmY5tHtukp2WRW/
K1VXgern6yZmR/gLxncV/VS5bz+EirL9fq59mkarke+N2eWHRB3jn5Xyi+cgl9VG
oF/V6OXnZZ8T2RdxFqugVsMkuhdFXHW3UxGp9cE8yJxobWSa+W5IOO6Izys7Atfy
47EDbU///wq8qsz6yl5Zgq/wX6TYq40s/uxOZXjDaszrZzuVYK7k9mO7vyzKAHVv
BF3vlDM71QyCNMg+ZfGQcIxDEnvUe8VDv1KV+by+MbhelUAKEmlGdjR/yAS1mZTh
`pragma protect end_protected
     
`ifdef SVT_UVM_TECHNOLOGY
   typedef uvm_tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_OVM_TECHNOLOGY
   typedef tlm_fifo#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
`elsif SVT_VMM_TECHNOLOGY
  typedef vmm_channel_typed#(svt_axi_master_transaction) svt_axi_master_transaction_channel;
  typedef vmm_channel_typed#(`SVT_AXI_MASTER_TRANSACTION_TYPE) svt_axi_master_input_port_type;
  `vmm_atomic_gen(svt_axi_master_transaction, "VMM (Atomic) Generator for svt_axi_master_transaction data objects")
  `vmm_scenario_gen(svt_axi_master_transaction, "VMM (Scenario) Generator for svt_axi_master_transaction data objects")
`endif 

`endif // GUARD_SVT_AXI_MASTER_TRANSACTION_SV
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
pLeDVBzt6eVlBhwzvAeUUkCqMNrHQxxREZ2Qam4dPeU1/PKcRkEWT2EfaTDu0Bbu
hhK41qwPAz+4k9x1sE9WwXBdisvgmQQjKxk8EXAC4zwE5bWMpyzOPI6vv0XcoZxg
RehPbvG/6piAXrpwsl2rlSg6Qmu7A31e3HdfATIn86k=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 224507    )
r5QZaYd9OQjS5TNWvTclZBFNqlWzDmqOSv+zwKfIV+ltmTMRrSR6KiIKX79D4aWe
onk/Yf8an73+Q+lDuItMro0nKn70T4dQNx28m9tdMYfZN4IfwGwcHz05Vp/5Ls5/
`pragma protect end_protected
