
`ifndef GUARD_SVT_AXI_PORT_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV
`define GUARD_SVT_AXI_PORT_MONITOR_DEF_TOGGLE_COV_CALLBACK_SV

`include "svt_axi_defines.svi"
`include `SVT_SOURCE_MAP_MODEL_SRC_SVI(amba_svt,axi_port_monitor_svt,R-2020.12,svt_axi_port_monitor_def_cov_util)
 
/** Toggle coverage is a signal level coverage. Toggle coverage provides
 * baseline information that a system is connected properly, and that higher
 * level coverage or compliance failures are not simply the result of
 * connectivity issues. Toggle coverage answers the question: Did a bit change
 * from a value of 0 to 1 and back from 1 to 0? This type of coverage does not
 * indicate that every value of a multi-bit vector was seen but measures that
 * all the individual bits of a multi-bit vector did toggle. This Coverage
 * Callback class consists covergroup definition and declaration.
 */
class svt_axi_port_monitor_def_toggle_cov_callback#(type MONITOR_MP=virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport) extends svt_axi_port_monitor_def_toggle_cov_data_callbacks#(MONITOR_MP);

  /**
    * CONSTUCTOR: Create a new svt_axi_port_monitor_def_toggle_cov_callback instance.
    */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_axi_port_monitor_def_toggle_cov_callback");
`elsif SVT_OVM_TECHNOLOGY
  extern function new(svt_axi_port_configuration cfg, MONITOR_MP monitor_mp, string name = "svt_axi_port_monitor_def_toggle_cov_callback");
`else
  extern function new(svt_axi_port_configuration cfg, MONITOR_MP monitor_mp);
`endif

endclass

`protected
bI:CV7EXAL(1egSd_5AaC9IG:V)Q#KPD_EK+PaI79&XW#F1Y0\AC1)7^gDC7Y>UX
19S@NIa,G#<MFe/#@;6_X45a)b7[R53A#>d6]dQ[>Jc+#;\N2M[e7O>TefeSR-+N
f:W13&G=eG<H3:.?>LL&L0UYP_/GJRPSM@V]<cZZ[_M]1Cb7^QW_B/58_9EbF)3P
G?07C(7d<K9X>K/J#))O?<&N)5[V-PL;?&)RaXME_)7FePV-,XeTCTEBZ#U=b])^
JL):B.&VB,MFW2A_&@Z99Za@eWK,25dgV[e[8e6gfN4b?2VJFce.Q_,cK(OgM59]
_6//F,\6I#,,J7QP+;8<O1N[M@AQZ6a8?_&?\.fa#T[=7/N5(1<@eaUP0agE-3_e
WbM,/aaZ_OS#0R;-L_&g7<OeKc<g#Gb2_BW)M14AJVC&AP-PFf:F=3@_<4R/<I:K
A(.dGbA&d\&EED9_>R;ObFHX#_g=^@T^4e=166T[,Z)6?6[\MeB>d;KEe;:Ae#K_
93&5<Z7.,FK-I,Xd9YcV;R5WLK1TD^D=HN-H##IQNReYOaM(9ZdPcIUG5g+I?CYO
H45)+SOE;(7.LV&L;&JZgNO>6>-\37(EL?ATWWBF\^OWQ)H@ZN[RUV/XW6S0<W1O
+EV&WeCaY/Y8<Nc,e#]9NP^HY#=>QSPdgfMFc)P\Y/(Q+?F\c-35TL@Ld7/7RBOP
-#0>&g<SSeUZ0\GDgH664bC45+AUG,b8,AegGU<W]4#P1e-@+;>EQ]QAg5Cd@Se4
:4H7&S\LG&XANT+&]>GP#S=V#:cA(E^FK_?FeG9[INQ,4&1Za<L=64g/V1Y&(efT
?=S,N9:NDFLUdP#U]3[KbI)][cB/G+5OJ+P<=>>C;RQ;;O)dcOQ/K=W\[L-;9Q]-
[>da-e2(M7#PVfM\W9[P5I7FI1UCJS=K?P,N\YNcNfEON/WQ@CM+JU.KZWXJ\(>X
&AbU)#486(aY]Pba/Oa^AZ1SW]/LF8YU30MQf4S3+F\,.>cKZYB;SV1>\T/TD__#
VY6,8YT6Y01V,0#\WDT>YZ75LEDA<HeF_]377X>Cc>)+c/0[_2]9^+P,:0;ST-\R
Q&AH8D8dfJaT#MOTN-L>O5[SXJ1]2IX7T75UG]/48[Oa7YN-1Cd66de3G]M4)gEX
N1>&Y-GM1/=^ZI_M2U-J&?^8UMO&IARZ8)=ZLZ.[--P.V^A9P?T,=_8/BJL>PfR:
b(bU8bd+Lc&OK])>Q/)\_WOPT/=N28_C^C2OFKgVVP6GBP<6HP\SgGK>3/d#ZJLD
E5(#MPZ\:UX828>47aR;E;TH]Cb9JdK&JS)_VbG[PV:/VdTBC:;OI+IdII@bcG6c
b_I[:V@46FO[_M#)7V(>cZ/COaXI9?8+gf@T:7B77^eX(E+cE^N8+fDcf#EGO&gb
30KB]c7W-M#C_NJ3aR/V-A=-+WDWd5RBQ_9+.SfA)gS@HRG9-_J]QSQ#B0aN_Z><
?[QVN[-+2/gXXa@L?]HAUU764J6+7c]P\?Dd/0A^HY?DaZELG/N0:dcMMVND]N2,
X87-a#GRZ>,2Q3:=EIO#PgZ?8,D0B&(E?2IJ)Y)E2c&5L-2CdX4^9F)cKMTPM:\]
,\<1MDS@,SXUW8U-@]W:b4Ra/RLWL4N5R8<&DQ=2D4Ef&1^fTDV\]R#-S1De;D&c
Z(^B9W>b_Y0QXR#:Yd/aKcX^R(3Z>3D.HbM&(B:2/QRUgZ.E<LY>RC/H[53Yeb#U
PFGY#]CB@aXN+0IOZ8M+@>edVPgcLFSQP&M:^H;2:&@33LFLF)#AA_W1^ZFREDOa
V\.F5EX5:/6c]eLD(U-S7W#S?:baJ8KAWYRVZS8fT5dT&\BWT2d\FLXZX7:LQ4J.
OPT_=+^</FVa[EH(@V5fU/,f6RWB;-f=Z/a27)&@#-d9]I8-M]+SYC-PFVD,WO]L
PK[d9Q>(Z71+gV=+gVRP=YS-.HeM5B?:TV2:a7B?TaBJ5B)R>ff/=R4eM6CaZE=&
;]2c=]B-QSG@/V6a^8Jbf,\A(</c:aX[Nf[5CaN.07UDEgS:AN7WbeMYL=+,8a=e
U5\M@)f+/VSY73/2K4dXCaXH?]_eM_eDEBE11=RLB/+U\1&F=9=b0896CV:DKgD=
[ZbGEC03.F-1Zf@ZP+@UGfVYcZgUGP,1&>K:@#;0ZP3+_.Fb]64X>N=Y-I,SC+9@
WaFS5CCbXIe7J<5J]dE^V.I,IEI(_HbD^SKJD3/FVHS2V0R#f<VLd>f]-BXDL??G
WMSSB0;E8ga6d0F2g3c56&0J9-A2]MRQfC)[U][He;Z)dWYE1a4VV=;QK3=/VfH^
RYSF6J\9e\<(SCc6&AZHYdE1a]+=/4FLI+F-ZL5S)A]U4;W4;=BVG[XWX7(HBbTd
W)0@CS3;L13b:GOH9g7d8.agS&9d9N[Jf0fd^O2GWLa;b5QSG,3#TS>WZbd#+Y[R
>XI1a#_]-,/)D3G#dH[F5C.6PD4Tcd,d?YSAF9[L187?G-/2g0f_N>:9<e]JI+Ta
e/d=BQ5.\XJLgBNA2^J8C41;&^WP^c[E3+f5TKK/8[<41Y4DI]aO#d45cQOA)Lf)
4RK=FV3+#R+/f,7]35ML4VA(<=]Q:dfDCW^AQAE&ceNd<N.d_[ea9MB<?1#XBU#e
RKQ/_Z6OC;ZYKS13c_?PQ5:0\)DM^e-@V0O5&U-@dX?IHa?PW?&T@C=V&XO171M9
Adc\\2.GFb/@#c:Ja5e@]T#N-@3AW8X/A5+4RSV[D8R\R;WM;<E0V;_N;#_Z:H1b
[NW1H>#3NgQ-/^Ub,@W9O^IdLS3@QNM3]TOU)=9B@N;;7LV3;P]M(&^e7+gQ0f:L
DC&3Adbgb+d,9eaT?NA)GaVF(]P_2J@.dgfF]GQL.RO6WE:L;FXJ:3G1,8ZY[F);
VD]D657KY&B\[2?=MWH\>^L_+NJ;ON49c&])E?Fb1,f+@Tc_,VfXR;;eX)@\O78K
e;UgP9G^@=#5]UYW6P+-KFB6YMF,I,PUG7N0UH:)T5ge[aV)A9ReaDaMcGWH31)R
]K/<f<B?^K)Cb&78N(0d2C);\Pe>VN3NL+PW6c1C;<;BX@O:,+<#SEQ?7J^8[[<\
+)=9G5@8b2N9@@[Y9Z5C);^;N)X2I+L/_Kba8Z+9aOQ0_:CGYV6gT8H&R&WLdU\D
5Af0&HX4>,Da-K2ZZaWfK-47FL/V:+ET>#eE71())(BFW77\?eUcSEM@83J,Wa1P
A6aVJ5[?LQ\/T_cV>/4N6&)9+9G_PM^]2-I<10X06eR06#,E)\_=VRJEQK&FG51.
4+YaEIH.[XD)@ZXM,XB5H)^VI9a+F2Ub,gJJLF8[c.1QcfA:c8^Rf1E_8>SY#>EI
=A>MW7b[F(AEO^&=.C&WC4TC^DU0#@2:Jd).R=K(+ML9aVP];8b]SC6/-HOd43_F
Q6+_-=[FS?-KVBN<=XC0A[>/Z@a]VK2N+,LLMUJ]/e1H:O^_3D2UHD+F\:D1M(6,
(35I9#3=d\?&&J5BN1?()b?5CO\#NSW;>dGYLO:?f>RA78UP0O>FA;c[a=f9BLc-
0g^B+\_@K)CVS6+PV&bPHf#7J69XQF0H(&U9]R/33&_\KdZ.;gT.#[CQ3baXCD1g
R7KDES:)<(5<Z6T;SGg6U)W5,QQ>3^U;A>dcV)eXegQUG3JBDTXa^,^KcUa;U\]#
[.HGJ&fbe;K1J?2eeTgNZGQU&^-Fg+)D((IKA9g#g+OIK(;C]@f8_#@d_#VAT+RY
M?,bE.0CC?4XRX\C(:1?J>@SMeYKVH4,T=1:5.ZX.JZY+9AX&XI/[=EFO:4GGR[7
/VDU.#KV.I&)PZ:?1J33KW-5eVad74,IQQR15BS)Gc>]BMF,V:Xb-6_fD\L,VWEO
/]]QH.+_.;B[UO,#U?MJZY4[DL3?2]Uc^SL#;=<1M>B)K2HAe8-80Qe16>81\)0<
R=X,N,>TB,bd^A=_Q=Vb=](;WVV(COUa;A:G<g=A,1F<EFPTd9OFI7I)#GAc@>R,
cTcLK?4CMY)H19+Ob(/54fX+^ZBQXF+RJ#,(UELS8VWY83U<S0UU(]+^/O\X_HR[
>e[2NVb=+.9E_:.&1OSANfbD?J[;T-GUDH.8,J+Bg[BU8FHJa<#Z/ROU>#@/=??Q
],QdMEX5D?UT@Qa8Za2Fe_)QZ2U:VOGTA+-9WVPcb_87?eFDO#;(]80T,f=56,/1
2.4=_<V>HT&&3/ONLbE]D^Z5#?(X=[PUJd]GE#Td](Q^27C4_0ZQfC7ZgMQW(/-0
\PgE+g10g/]05<ZKY=5dHTI:8NRZEdAUPX5a#@<1[ZP2?7IMR81QN5YDGQD<1/+T
/UZcY7_O7VH[I=L,UV8.gI,&X8DGG[_5,J/^,4+ggMTVZag;,:b:H4.[f::NbHY[
M5L]Z3#L_-Xe6N.eL869@C?O)e^)/bJBHQH.>1b>^2<(?YVZ?><<]FM:X#6d_1PF
JEAQXF:fI@63A,e[-^UB2d,M2&WL\VBb?]8B66_;>AKAP7.fROKSCdO;BF_agA>a
]@S,\6/<L)W#;]7JI9L^S;fG#ZeR&AUaS0J6+HB]WE#I7d<?8JS0W^U-:(K1VYIZ
2-XKO5?CF&EZE/56KBJ>e8I_)aU223]=TA^)b#M7V#].C_,3/+O+L>/Pg?AM1Gb2
,G&P#BP[W[WP9aY\H2(^-D9IBQ0-_/gNcZ5_T=AQAccFCMHUKLb^?9&W]GJ\+E8F
YON0P^#1bTB8:T-&a\;_Qcee73<KB;C/A_fE0O7NYa926AMF]?5JV(3.0VJZb5c_
BL;/V;c^+?(IKd3#<ZML#ZU3T)BHIESe50cb?S)B690fT;R1fH)D2Z;XF80ZXA]7
PMT]F]048?&M?-L1QH[6Y)gCOYB1[0NOc94?7_Lg2ODgA.M:[NOa<\LFC0&067b:
Rc-/8RcVd-+\cM[?e9O9ID7XOU^J_/cfON#>)WI0R&(0X>b7LLP)AT.\(J_5?R^-
LK4S,--FBHR>\NQJ4c.[9EZ4#U\+L.9.J1BT#;dVDUM_AB_AHdVdReXe29HT^\23
9eFQM6=GG0@6^4)XFVQX.]X?4@A^gEXZ?\afU+_N[VF460Y62g&MeWcVaF0^@]6f
CL.JSLaNBX:ZGb3XZA;_6=1b][W(GN66P682Ge3M6b45@8e^bXEA2U>(+E+;bDTP
_f]D)_bXK-(FYZeGR/)adD2#R0K@C:X._ZcKePHI&K=0a1TY3S)?48d&;2,O&/eD
\)V6C.U/U&f<3^:0633C5M>40J[b,(;A[ae-DNM^N6Dc:O=FYH)Gb5dSL_B0^C6(
+1UO0J_DC;8S0J:]:_8f..K;9DU1ZTSR1e,_57HV+E&fUBAX(V^/b[,;E[>c5JMI
aR#Z5^Uf4?B1ES,<GJ&0G<eLG]&[:.#6ZNFMfN,1agC_K?MBC>V,aL;CCPIIY#-V
?C>A5A4H\=AI0VcYQF)B_f<gWeECD-FGJ5?ZWPdP<5C+@YS=4D5<6)Q=;Jc>/_^f
@7bM1<7HUM>8E8C_FD8?I<(dSVdQ#f>X#5F9c,LP1GX0b+1DVIgLVc5_H[2)Qa^I
7A-7Z5;2-/LHJLC<1GIDD7\XcB4@P5P=cD.Oc/>9E68AEXOUNX6U(JeKW.01+@Za
CFU_#TM2)TBU9(,Z6bXQTNBQ-(:Va[1f,,X@A.^a0D#)Vg:8<OBLc<([?)SeZZ?0
J7PV^@^2235<gd7O:>NEZI1Ic)+3A##1:fdSKDE+:/Y&^0M2R(&BN5?C5aO91d0;
VZ&9a280f7EBV(3DG.Y@A3UYEP6fWa@@D,B<3D.\]BFX>9XV^B?Qf1O-R57UU)4[
]U@eC[?94\C<:B+1\U,5QR?0_^(8X)9:@LT3<b3WK_VZ)5@K)8]F&9WRaSAK.6d<
5d=RVF>7X77KXe\O)G8L?_gUf?J87&RSVbVDR.)A4Y.<J#[7I],7:P9N>[C8aM^b
NB\:g;EecP8gaL/5WAf1Bf4aXBE^4A:a/[:YUGHa&]AOGHg0@#g(XH2,bRdS5N@@
b+K>])Af;1XgeKBN#6M/#&@gU;La0,J##]V5H6Q8,U^D4(fI9bMc0V?c?PJ\_JI>
Ug#C.-]0JL1WgY#O0LZWGGWMZO=f?67]Mad>KdbRV&2JNXB>3I+6F>JWL?&J\QV#
d/EPS+0L/-UW:)+>?T9GeCDR9W:5ac4[(]K1T#dfSbX@#Ha/cZ1C=]Fb,RV&O]^;
]C^[HY/]3MD?Qff.:ZV9U\UH&b5NW:.25:Q5(NRFX9e+V:(^=,)QY;;.0)RFBQHC
^R(+V3[DL_TA=aDA^1P:J#G(6WZU>OHa9>^KP03?=G5[d1A3T:NfE#&NSBD7#KP[
OfLH>+N?+7DBHE94)Z?WbMF)Fg_4QJE2JOQ=\J^aL7DF5MX8fH2;JBf,^9Qd0T@f
\.>LHgK?2<I<A;CHE0)]N#/2b9b3_=S9I6@8#G0:TFB0F(JA6f2]Ie)I;4G_:AJg
LJ9Z5Oc&N@U(8@]YJS@[1YJV[<MZbNcZ9?0FK)S-G3F+U[JRaAUA>La;<Y-CZ,.3
X^W=G]2>4_>TCNH/28;9_3,-:->SI^51@<Dgg38BO-cA&:PSOWVCI=\d\,9\_2Ue
<EdG4NVBT.U8ELP?WOMOc@HKVe/4<I#HZ5YND/U=>a@;T_<5F7[AHFC9?+>Oe9Q@
8)3Ca.L6U6Ig8PY/5DR&7OZ\eZX2B\#_B+U3(,J+E(>99Q<a=?HO.&,]=RN4fG9#
)]a+J411ISSSWL^GeVVX17Pb]cP,VA;UL?I&54J0VB0U=gQ>VIHW9D;FfaP+geL/
A9J^ZM5-LK5(JEQ(c8UOAEdDgS/OQ/)(J.7:/ZH1<c>CN6c2>A3_<\a<BR72>1&-
N5B#HHGCG4J@]QY+3D69RS7@?B]N.3D^Jg#E:bF0Q5ReX70C9/Ud;B\g3e+Fe@?[
H^2[]8?)(XWG7a7KWZC]9W<HK&?Y4[,T:G3P<1bOEW^/0?,BO3Fc0D80[fL34X/#
ggPE.AJf.@^,8&]E]8Q/D0.:#b\DG(W7X[a=>8c7GB4a(J1)DV7Te78(\I,=BG_N
b\^/K&>dX6CN^[OUce0JW<KDE2aXNAQ.UWWLaX1OG23KKTVITQ(.+\TDCY.XCUX^
Z+1.;28CeWedSLaB1P+20K0/?4;c\fWRg#PEV4d-\BK)WWB44R\ZH&39S=+a5eIG
)+JeO-WS_6T/0PK&6M]3QXYb.PAbb?HWF<>:TW5TNW:1_6gL00+=_-8:G?BS?fAT
,21ONXYGRM/bYS6SD3V+]4>A3-TJM<:0g5:RaeAB,NS7=MTR=4>T>NIR_]SSL2MZ
LP<QL<0ZFYQYDbG7B,#Rg>0@L4^26.AHeJ9C@Y?VgR_M6fF0_ALg7_#DVD;.&Yc.
>V76T,[K(>+aM]EG@.1HI(K8C_J8-2cS<M#DeLdYBTG0Id#(f653#KVg#c/UK-]A
7((^fJ+^09HEU#CcP_e07BBK=9TaBcWdA&[4e;6Sb4;IN0Ff/TNL5O7/6,+5d\3a
<^U8KN\7Z=8Yd8dAPX,aQ9/?I0g&?#faW9R/1<LLC=H8>EaT>:SJT#CJ46d[88_9
0N-:395(fO?)HTKCgdTOEZ1RCeVPL_Vceeg2_[?/[MH=J#/If3&#/9H)e:TF+RD2
:ACDR.+\ObSFHURA]7O-3b[@dO(+>BS00+/8[CDb5da?T;HT,ZSKZRFPEKYF8P-V
JLDBSD6XQE(5dHS,--(C^EKUA-PRPUCf8F46[Xd)UW.^HKe?.8_WG:GH#CXg+gH_
3H#^L+UP#g/K,&a,::38K@f]FD36X8d?eTA&UL)TL_FQ7D^ZCO&65Q6_2,]P_UNY
faB9QbgS^88RaZFO9G^Wa_VB-32G,:J(INa#XSI&0?5KUTQ91LcBXON\^CCIZK^]
8fc-5F1ebcI8(>9a)@V2T2#/4:-PY?1H8F42X+AAW]-Tc;DYdVB>EO;>G;6.Y:J[
e2IQTKD])E<;<P7+]=DWB5]QW756Tg>^15<K4FY2WF]Z9ab(56IB.,W_;,F54^Q8
>(U3E4CB\b41B?&^X_WDOd-B^[5f[BF4=e[(:(Y?H/K/DH4:EF6cE78I[fL0cI9O
D:5JY+,egb959KM9@&.NA6IW05L&&ZJM^^#fa;7>-5,fZJ.__,4(^aL.EU<^5aX5
44X1(3B+4O/@5d9>HYD]O.2bY8<42N\P5<9(U+8Y,63Q/^P<]3^caD#(@-W\H#Na
fSX2[#E>KaeJ9_D=SRSR5QZ?0SP>[7#2;ZagPE^e;IP+<dLBcRR/(Ia#.]PIHg-L
YR=@6Z8PDT8IYC]?(6WOM1b]268K8+)F_5Q=dFC.\#5/9&AM5JTL020Q_]2cbYT]
1RP[1?7I>_^3^?7,F26EZ\&b.1G.;0X1C0V_P1I+VF3DG[R?1a@cN-)NEXd#:I]#
NQ<=f^7TYB)I99B;]fZaD,9_DTM-X.)Jg.[KgH\<W\=@\[O<;+KcedaDL:2GKFST
8GNO3XeO9EaRN6@eA\Z+K:3)OR9(-6-;,b-^4QN;>EVf32BJ\-W,/7R[fSWE]1bY
P=]O=6QF]-<(=CLR<0#DH=M0TLE?F56HT]1I:=7L&ENXQC_J,TY0<1PVVW_&.#9M
6a;@U7B,Z@E9A74+PEba-QH3)EQY=FLe?E363&A]0gO.g(AP;F2(NEde7R9^;>(/
73&FP]4C?eV/DHFa&<N]A00a+OEAgKHH(e5d)+-A)-I2X.g)DL>cJIF<gV]I&)(V
XE_B2GdT.X#>/@Y(.R5gX.+RI\[C:4MSNZW78_;SO(<50+5D-IWcC/2<R:+b:-gU
PD(6-)b?dWP;\M@PFIUL2?+3:L)&Q^WZ#C6N+^J7cT<7^Ue/fOGPF2YgI+:YceO6
E7=+#^a9?ADQ7WF[^_-J7>6^L-A\\HO>_;a9bcCWM:IBI0eRK+&<LMG-g.J6.AXd
ZfdQ+^cc-fFaf5=<ddD.KaIa]AbL?I6X@D+WOY6Le4a<EWVF+4aRBd#Z;e^Q]ZUD
GHP7N5BT1_=XR#NMXKbQ_WI1cBC2.\OeM3VFR,Y@1+4_=43#)XZ]IEY7AK,D)2XF
ab)K4UJOJG/N],K146<RXbLTOHcgLcgLRYGF:3&gd8d9EV#EA]AM_#?+[@5<U=U&
D,aJ8;K&:9R5gB/LaVT&L-BYR03&c@P#>Z[0LPb=^UfQ\.XF:<g&[</f0Ef:H/Ha
0WA[-M5&G/R:.,UG.QSINW.6/e>LNe:.c.4Tb]ZDgIE_JG?EB2WOdI4Gf9)SL&Lf
a]0(K#FLSf<U>KFeea0M8:4V;S0/fH?[HU_JeV6[G/GZ5(I\C&gYS6,;=OU-H7/c
HQJS<d&K/[FIgVIDY7#dE/7_(P0XK2NEWf6M^SAWXF#L/^R_f7B4ddIgR>UW669e
\K&Y[WP[cb_/6@#c-Kf;8f+:(HSR\+N2<\FefAV2=daVLKg1AL]eL?N0#JZI\B?I
abf82VXHKZ4<YG,&HNP+a#]I?7HBePG&dC7VL7dAZI<+CF9UI6XU(eY+<-_NgI;1
\&g?IO5deCA4)@730M0_DS7&CNWS-P;[\,TGG9fE8P2\We=R].VdG9g1-\<JM^0C
^GI-JB:U-W?DX2UddYf:0aMN)5,0+eFH<CXJ.cTGLMaA0QZ;_d(dU6+TL6a&1bbf
]C]LI>IF,DEgTJI8dW?]e6^X>-KBCf4^B,\KZYWIg+cP.I-P&.26b^6;)MO)>OZ7
eM:ZN2+H-dcG0YO0GYZ/GG&Y^U\=?O-^?+Kb;G_S3@<X8+bI?aN>?M+(H1K\CL]M
d_V^gc5@RcWAIW80^O3=d]NNBH>S3K:PM6FK<0^G#a/a&>_]GX9O\cA5IH1#T[.b
^BZ3X6:N:G_3I7cR<QZ7>81^<?]D]a_=5E<DAUWY:L?(;-NTKE\T7AW<Z2&_X0ZK
ZVGd\_Y9.FXf.#TXCAC7?c&&.>/FI906-Lc6R([#f@1Z]5EaBe)AQ<+C3-WGdW@_
,_C+2S\:PbW@b4S(K?ScOK[5QK@?<PTQ\af=0]ae\D<UQ5R\SGT13.+AgfJ2?EK3
7W8#U2YEd#L^ZHVZOK20B=4Z@T5T-77\Q@L2V]<[\UH5@BAdaG:NU..KK#)O^/_]
b3&(DMR-69JJQ]&&CVB?U?C(@</X^(>E0C&<?ag)DQBCO0\UgAg3)Nf\ORR:[B;M
5bK+9SYP#V]]PO]YRJ>U#N(+A#5>2US6@g[S+T=\Y@@RMfc##gY9ZJ57DQee03fB
eXF=0#J8-OO:Z<c=Y@2J(TIX22QMfCd4c)4_9A8QP^16eE\I:;9gb-MUHgW(F5M1
_(1B#fH#I>IE8T]WL#.YN-8PG40R31[2,ME(&\CTQ2^L<VHA=/GTHA7\b[U])MX[
)d#c1S0NO3See4/L&Xb-JHA\ERNHG#fY,?+0@MGK?JH>9;S[Tf6ZTFXdE?DL32S#
3[fKS\dWJ=>)\MA.AW;-D0#1_TcZ)E,2-M.UAeJPI.\;FO^+#&Af#;?XETKZNJS4
]BKc1I6cb^c^KE:aCg=\FRbcT(]O[P)a-bO4_-/<b+Ua=D)IOb\0+90O58J?4ZOQ
Y\56+SCYEe_IX5NG&&N.(KHH_7(ZS+=;be2.B/]3<;/B-M</Q(LNF1(GTT=LU_d,
GZ,LK-GYCEaCZP81T7e/P0HM2NZ.J39fOfO>TWK9/aAS=5e42JN/UPJ7S-\FYbf,
M64Ie+C)KN6YBRTg\68AP>D414JAF#0XO(P1+19:-@<=Q9S3(G(9H_#MCEWYR:aE
+,9Ef;b:<&&@Bd;12JU)X9W,>-R_?,P16KA5Fb]2I[2@@RI&2?JSXb3QULEg(J[+
31TGQU=,9d1UN7N-8Q6FBOUB//Nc</e[OB?ND4Y^6RbD2,B(YAIU312;<GN\W^_W
CI;O:MC@[7/OC;O;TdO6\XOAHYea+.P;+;b+UO0g9.(B8=Lb4MFS(QZd.YH&BL=D
dAE39G>bWH#9W6A;&P6V#_ef<=gZ;RDP^.dA3US=,\LRM_B68O.gUGZ3:@/fbE^6
ZUAB1ANPb(?;[R)265^[6B,(f1IXA)ef?f)3I8](gXR&RBeMP94OaNFc9AU744OF
CFM_XG?<^,4F,;e+PK@8#=1^5G>bPTe_Q^H3[/(;GRM4&H:G+=f;(>;^XCd0#,R)
MK>HZ?VV6/.>(XcFE:d21aP/VU3,())ELBf<:+J?4P#H.Mca+8dDJVf@9W6[E_N/
1LAHb3/II(e^9e<(MEX@#]4]eb30-+B/75#Pg7]S^)OEY1;NC1K=;:>E&d/Fd))>
TZ<FHYePRO[5E03PNb.V3.^Z77cV)V9,T=[5VUZ>/V,I<[/6O?98U9R@/93EA9XS
G,PC>gKb0)c6+\e(2R]A-8><)G++0c/#gTEENFB#EGcH\NeX\HA+?VM+I)=<,7R9
;XATB9-PUQ^#(3:F1D:LDF\cQ9bW2>&HY]7.a\J9=C.UCFcJ/RFQ^b>NV@Q-?RNL
3:0e0:8<<Z8<NYGRd65E,eUU:_Z@DE+T+^(A(3?T^;#Pb@+D,H(,Of#JC58B;MH8
YUT]>=QU3E4J-VR5E.1WZ])^g4?&CD:\+TdY:ZbL1PJN(AEO57IR>,,?<aDM[URa
:/FU^>\IgK[ZV29A&@K<5g(PG;9&:]<Z2(&H1.NcS2NY4?7U:L[@,Ce[7bE0W#LE
_G=G4?.g#\A47_RNPD#86)YF_K&:HDc2bB?-fGX&8f3#6KJ#2Q];0^&@8B=L0QbO
M]GQ]IGUW0TKI:=WVL]X^8b?B@U++AgePV95T-6(5>B03>A,K>_c@dT&?=5[AT1M
2_=WYX@8=UG<E:QPcOQ:JV2ge)LUNcFaZ,:Z6?NB,<W6Mg=GB>\BI,2XMeN19L7K
OGDTGa?e0E=5^TO6Y@&+W1D0]BQU_Ta8.Z+0(R,d?FNU7__#e#2M#CD?aaLB)<=G
Ja+,K=gIgZTT+^AD4F<cVS0,85-&cUJZZb[d0ODQARVJK0QW_@3>0HD:SI:CGH?G
K^SbH1cWLC=;W:Y=)MN-LM1[NVAD.5(L#,O>=EU@4:\DT#&4ZDdK0].6?6>9VSOC
Q5]c]ccS7.\ge7;BS\ZV[MOeP]gf@,g:gR>S#[EK^D:#(PM;(CYU()[f^8(FBBT=
ZBS=0DKF^Y0+WH?3@S/cIb:5GJ2AA)LM-2^5c[B&ZVX;/=dK4O<#+Zcg=GQYMBAQ
=:1([<3U(@OIMcf(TOZ:]5J=\-DK&<CeX+-c]ACI0@Ge,IfZYf33Uf70\(=X(75b
[W&<XCUC^(ZB>?<?M4#Y9KJ&WS(A[=Q7HA;E^855@?b&TC(>Fc[V[->4=8L,:/ST
aAIM<7WQV&V<cUg>.0KZHUS_=F,c\L<@^FBT^S#/P+?LN4>=PI1gO2S.e_aQUVP,
I#ZDMF9NWOgcAC#(8,-;I[I@R9U4[7EFeMK(&SOb4A;0:RF76F5JfXgJ3@JG?gJ&
,c.85D+dMQ4a^^HA-GAN\#dI8dTNEAVV^FV((3C9^&4bH#37TT7JBG.b?NSWbR2(
-PD535fVc?0K/_A/BCVK.U;5M5@bSIDgPAQG)<KBE0:QL==G,<6W@Z?4T-7BTTKd
C+K=8S#AV/^B1;:?-@>3EgA0=0^Pc@BI[)E-a^)Z0;@B:M1A<TgN]d]O[5(ZcOc(
V0?V[^#Aa(b\\G:-TLW.1>_>b/+1)4:9XIW^?J_^J][:<DN_CF[],GPfPM/e_LI4
MX?fLMba,Q-c2E071c@dc)U>O52RI4dYc@Mf/ROT?\S:L7c0<(N.YA4&LB--U.33
S9A?>fa.],e00c3R-P>M#DQ5AVc&M#M)JXbW@&T5F>;H&E6BbG9COK+I97)FE-[)
;\UU&fZTZJEP[:eKY-,fMS[]\MFgGS#>@$
`endprotected


`endif
