
`ifndef GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV

typedef class svt_ahb_slave;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hrdata is not driven beyond cfg.data_width.
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
amSPcMJhCR1TkDzXTjNYC6Dy93JP4OjWryDR3bHn2FkYWxQaNOFrIqAsU1P331UC
hSB/Alt58XiimLIMeT2pCXmfaApjd3Lu8T464hoxhr6yMejPRLM3XJgIEQ7Zn3AE
sIXUuG0z9VCurDTBgihACL3WVXbvTXkySz59aIzbisg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 367       )
Y5+sC1ynTKtkHiAtIEZG/6t/Klxvf76sLvX/0TjJTwAVT4B3xmE2K9NiHuJYdcfE
Zyx2jHzfStL5IHChDBUSN1Dr1x5LaLnqZPTaE0TRHlN3bckf+NaMZJ6MDJJrY1RW
XQSwYSepUkIEYFIRVhuS84xD3pKEhKvXSJo8KIHXa7rIPBB1F6qBQW+M9z8GlBWl
yvWx7xzgwUU4LnbiIQg8ojH7CqjWeSFk6M64XblIvM+6In3rG1NIKxCLB9vmOYA+
p9Zs8Q9U7+DmzZzgIcpNLGoXuCL8psmGgOKY0rxnV43aKn7UpJOuhtvt2dutR2wB
sgml4f74tX2tSeQYu/ZBj6Qnzw1YfEt+L4dguCY14OmZrCCDeZAuEmcFsa5prjAz
BM2HYlQf8gzdMIBFAfWDCjGsVGD/kNAq4iYKNvBs1rxzU9MXLLibg0vGsq1x/7H0
wA/4UEZPMh1t7iaiTCwIuDbveaSfLW6oF1KaPjJf17c=
`pragma protect end_protected  
 
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_active_common#(type DRIVER_MP = virtual svt_ahb_slave_if.svt_ahb_slave_modport,
                                   type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                   type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);


//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
S074nxUrolE0HspsOSUjtafKyawFlDmRi/Sw2eSMvy6VnuBageMkRZ26FdE5+Meh
LIn4kUotzAAUV1saS3X/4xm3X7G/Q3ifZOY2KRMU/WJlPFp9MneP5UBi+fJRMOka
OcJkHQFyPVJLVe28/5fznL+Y6jfc8InOEc4+236lb7k=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 3939      )
CZjz6rRk71Mj8aKAC0iHruXOvvccIYsevPrsdq3ECfY6XrZF3u+9Hqv1dOoC2fGl
zJdu4lpgr26QlvUlHyyaatuD9SyfpfpJ1q+UNvTxR1PMctuuIE4DykIYUtitZbby
GHl1ZBeOy+E+3HReGzYbCyafylWQ/YZ86AsoZqm5/LCyLLERn9krk8vCHqyORTC9
U0S2lSYWYhe3uQTvZhCB5uyDgVrozznxloOW1E+fFx1NVHLNN9zurA+yBn9vuuKC
vEQghI8kEhsWJYsEXFBMdcIvTr5ZyfNSC3N6jtVc1fBnAFgvJ8kcTjEMQG8QeySD
3R3JdqqBTiyueqa35zdDqBamzySL/Mugv62/SPpWUNg1SqdLpk1rEPXcLZghSdce
PYOCUg1yLjKP1GKz6njzQp0mGrpQONip4gnKj+Zvr3Dq5yY2kajXWV9Xl+zOV2Sb
UkVd5oSwT8ewlfpubcs9L3QcShA2waQZIWXpPuRiM99yRcSGK9MPTWE5g8Wm3bEo
5xzwT7CIeeoNrDOVpVf296lOJLropgJVgK8k/9bKgGRDEjwavkjpOcKbSqc7JvPo
A9GHEaZGLIFngiBrh3F9mbG2tcCdIEJ937d3WP1AgVmRFrmNdFIMW09oQ8xlAgMb
IfojI3OUv47TvJBOpQTjZhSWjHulWUQRwA4uy7xJZKEp56IpN1MvehcoTAhap3mY
N9MpZeiELAjUerrZYhGtIzUOLTY/1Cwz939orCHsIl+WOjqQD4hdgiTqF5X4l1QB
mNvpqisTJgvqpGUSiK2ciqAa6nhh8U+ZJW5xTFnkrtejKkxoSyrnFK9ftzCoI3KL
ks52eThwQ7YX7NM++m2A6HtP08YHcqhpk2tPB8yG/hnivSdr7p5CwbvxADsXeYrv
rtUJYgdOU/HqI0Td/d2D8Sy7uYs4XCy1KHCZnfL/m7jYNBBs1eo+xdlFA3f+t1Vi
Kza8RRZKJQDwHefjKlTBF2vjRUJK7oTBSe2d3EQqMUse4KJO3kYpNlE8mdCZb6oH
os5hqGYyiEMEH48Q+rgPIg9S15jx1355THTZkMc205OrzwMFInHsGpgRpArk1bJX
oVT5PdzMkmLyBIOx+kk0S8Vth8wQWFJCzTBRqGL8QqWBNG0fSJfbXGbU0MeyyO6p
+RKifj/M0mGEh4n3QRdNO46d4l3EaeEHW3FxqPZQ6ylW2+ecQMdaGRx2Pt7EC+BJ
yfFLALexyJlJUqtF9VwW9aSNqdyjWRXkw9AWaJWZuTdQLJDOrJSY7pHjCF+9RMug
N1rdoXsS5mIEqXAdziUKod+XP7/8Vr1Xs09ISg0xiWST8Xl5+PYlwQtCptVUaxqo
jxU7CTODBQTSWkLWT92Y7F9041f9buxmieKku/qI8kFLKxLeoaa7odCqQ4SHqsZa
XzpNtkyGS8tILWpWvkpZH0The1qj+LN8i53wMw5GtixZl3qhmjHjfwmz2X1vdOlY
c1Lv5u3Ub9LRx00ApGb+eiyy7h+eYSYDqE/RpMgCa4baclADHZYDAk8ZTvAcE6i7
2S37N1ESMoKBnvyrknUvNrp7lW7rjfpcWRFXD1eW+DAnQ+i6YA9PujkR7vapwbtA
ATM7y1Pja6q6qYYJN7diXwBOd/XGUu9tQUCcZITrNXmJM+V6lV7NWq1n2T1ah2Qa
56Q8tgl+J2gQ6h6ev1/k/rtF3s7xhRpAh1YHaXdeS4ViUK8P/1AgQatuxWKkVcSB
LkOLJGcewmbj8XRTB7fvgnt574U4lzqlyevvWvDSH5k8zIDrM7+YPYFpSQr6nFhM
VGg86NRksNqRWCRdyjZJBb76S+35JVjUrWZUAWmwB960tNJPYG6CmcRjxsVfZO94
O1nmr4F5wZPvMx7j/8OCD08N/aErv3Y3sYiImtcmP6cXou4ZbO8uIPV0E4KW+Db2
YRxknNzii3KhuXwVnWUVNcSAfFTRSJ4fB668pEcaYH0sMp0ARd7iOd47LaPodlKf
wgTHZMAMKsZOW3hDyJ4E/GC0SvqEB3uExMiwfrBbyDtaiayrvc0hABmYtnaU0bFh
lqTjsycnXTkzslsWO8QdqlMOj/YO+YnBky+V9Oc25X4aoJvwWYEl4T30m607qmZa
HmbX1qQQOI6xFOeZmmLjVvcJ6KskbWuZdrG4mqfijrp5F/o5+waNMdwk5D7j8IJy
1fmOUXoTyebNsqncVitK7sEX3kJAlqUWWU5qGL/9nnEl03SOvhKMwsOGh/RNfrY/
LvVYVBx9bMlhJH9lV8X5xTDO/1i4goKUJd7n3OS0vYmB4k4ivYLb4NLriiinunZU
6lebIw9nckOERkne3SCXQU+fISc72Dc9k/AtFZvXGVgpTBaGwJn3FKSUfY/wfhq+
h+tygMFcWgUS+IgZktokI0TBAk8Mmgozr1b0gmM6Ib4LGzf0FTGAidoRCOm6bUE5
eMx/trbYzHiijpXEPo0nvmSGIw3lt5mxoO/Owdg2yjgIgBPRoMGnTDowfJDKEY2C
uUhSjfXrGesw0w0053kEzYU6gpb8/vj5Sjxhn1z1ObN6NWUGAAE8WzHW7VG7z7WI
k1o6wxvd9CFbVrICSIIQgsvNg179rHwjY0tlcecQRP6BnxiSg80FR8y3Ob3atD23
Ktk8/QkbkOyuoAy4q+BhUEDBsFnMyq9BU3nv5bUBv38CunMI3naQ1WgGsskojsBA
UlBmZAAzZ1M4WsQ8hcvVYpsuXMRjsakXG6d7QAQfu9uRR5mYDB1gnLoLU5dWSsfE
9GPbop1c1gRS9WiuuRYttVzz01PwDrgFYVE5BRT9fXCI2stCYbeNXt23bLkVXkqY
2BP0sHGGRzYUx/zudvCuYfGS/WZd2qSF9oAXhW73RUd1tyydsyqxiP020E5Tv4iN
otKSTMGG1J8PQXfI4tmTG0KDrqgUhBP9y+HJAqF2JZeE5Rini462GDsmF3XHFFND
g7F8WDI3++sTNgbs6BC4oeL6JwFCsxckLfulMhUwVahNSlGjuEqpTgIEc4hY2Wk+
u0WHk62na09gak6SdO+U/+/AZkOa6jlCQMnIfuEim4M2z8nCPt8vq3LSUmL+Ah16
GJ9NIBn3zRFHsrUCjfEI4x4dAbI6vCnKhCfmjGfbkB6Mc0kz6IbZ6lPBdnKL+OV7
gX8x+oOBhN5LFMy5rKECPolfbm6qE9xOY+wbsz4MOM0cHunESe7lma3YR5CGk5S8
kbQ5liN0Vvf8E+tXlnveQ+Iy5MXL84QwydN9oWChw3Loythn/fbT9z6PvNf0h0Yr
JpKURkuYuFLiA21GYHfks686IHNL7ReZ7mS799qDLnrxVSGmvvGOfwHFjMNEBdv7
N9towjFMrqV8pwE3cusavp6OaLOPCjF/54+YrZ9E96Ols44GYRC3IZDz5Q5oEHMb
yAcV5CPU23jEArcgRuuMGbCcTiqPsmOeRcmIrGknwZ564GOja5jMI2G0UrpVnnOs
rAyrgel4Nl1OSqGn/oPbwEG1gvOAmpnUQlwpBeQAuIHd70MTOI+TCawr2yw4dRUl
sqVDEEUV8RkoJwiTdPtepDvCRDdAY9AUzDXPBFsVM/EOQXvLg8fd3sx4hSc7bwAu
NQJd8doNbbqWxFf2V5PcvQpAUF/rOK4Lb6XqdnpsoLl4h1T7vOzlqZffH4/n2IoN
lRsHriThJz4uBgoGrWK4uF5kJMpc++XFZGOs81nE0kU5dxPYQVZ5LrVNHdRdDGVh
3Dp2pdU2y1qfmq+z94//Qo4MJW3YEIe9FWwDsdr+H6qb1y/UWRfiJXofb1o82pa5
vocHkI+50NcI1UgKGvMEaqJWQEBkmwwiaLYtN87Liec0HzvRP9Bw9H1rmXOB9aCc
NzcByhjV5JVA2xVzbhZl67+QImc+KSZ7nZGbIjd/KM1OVi+zarDimJxwx9sOEWD4
452HK8YfTtn4kPyA6XtBtiv0VlXgHwHRGi0a58fLbK09HR6PILnmsxzsWXHPIm+G
SUjtbyNC/bBYVXpUHWol5RIMsv6oVngLQM160B1YrTKDs/HY9k7L9wfVQEUH+Gfd
5BeVC5oIzNCicmq/sqx5UtR8Uw/w6SpwP9ZLeDuh1CF+5hrmk4rblADnMmRa7bFF
8EraqwOuvm+lnM6FAJIWKyBZW+jPbxz8MrRYEXauLkgKr+qJS3uwwbQ72CZsttFp
DhLEmxZqE+f2sq+rdsDgp9njKrF3HxUNDk/Mt2obG70NXhVE+uu2Whh0bXN0Wrs1
tkUJ7e8ma2+xoNxGMFlJYJIKraF7ZCqMaCx06OuGoofAq+n8buQ5ljO89kKu4u0j
Ji6p8C7pJX9wiDOpr7KsuT4y2MWPkJmzHl5Yb8H8WVDlsNRx5H4iKzd4PQzDr3do
KBBrABEsQOCMRPaI/LlEbpose/4EtrD1Wa1BxVPliTK7Zq+h5+mTBWKwxQzgosgv
Drma65nTMLOvBEIOitxnTD/10ydPn8PnkuiAr2uswbMz8hEzyrRQR/XxuJD3ym0e
KdOfNx3wGq69symWmrZ2u7jTscojCmnkQEp9APXhyGzvUuhXzB1EiKwfdNUIiMuK
AB16uCskzG1qDpMAdQ6189lSTwpi3KFXlU2PeO9uHuQzLOxF+rMLoMyK/tt/dfAj
Z1BcnOpN8CCpvPS321whRNBxs9/OYhfOcs7P1ja2Wv+NZ8DjFtmvAo/kkT8wgWCC
dJp4FV6u7zeCiIB0HvUw7a0c+Eas3M0NTRfurX3jwQIW9rr87xSjMOjtR7KJTu0p
3tWemQ4/OSt1y8FZQiZgMiAq267c74im2/WefxAddIM=
`pragma protect end_protected
endclass : svt_ahb_slave_active_common
/** @endcond */

`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
CqfFHQhd12eRl8C//v255QpoICKFJRkzMBxPhndZ+WcGVdKGxLEto56IrO9CFO3K
4XqP/D3AfbKQJ71PNFFqKEHSvdX14G8OVQkOucMwW0y44bFHQE+P/U9kQNt6Oay0
qqte+AcL/zbDzP+hEWQTqzhNkZFZPuF7jLUDtpur6rM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 4492      )
ShRExcKNzoXZj2I1gIdpiBaoBP9XdeN16mmJD/I1zmldxq1FVs5ygDPXdlp7z+US
eoFaEEarZjsrD3D27tH66XFlPdzaYjaV0q4HTkHoPcUEQTAumvuEGuf7HW1eA4U/
bzijD4ll5rW6SNyQ1altG7TG6bnZxoa1p69uLQVzWn+n3JlDE9i3OR1DpzBGqdFS
tDU5a6xfyE6EAnaEx2FG2r6Q1Af9f9qJoLowXjmTi5zMq7P58qO2UQVrmeIlI7rz
reQeVIGrxg84tcJtpmbK9upouk8HJuc/7iIlHF+PqZHmDVtJtzH5WHqFChLpchC1
CLiRmJGT9P2AFWHWCO09eVFvZGpILHCyLhfdpsqvmd63lLzp7TJDm7lkhuQel9Z5
ompjM1l7tD8VtXrLmRX6WC200vULfEu/q9R4/9BBZBMubeTci3TW3WGNDIWOjQQU
AXPxrOUThMvncBZq5pjS5nQnx3tw8HG7/5YjTFxoRRpTvzDsq73eTTym6nlChelT
YGaleDQ7V30SV0Y3ZbOOEL1yfzC4jLtr2Z7jp3B/qVei02rvZ8Ni80a5He1XaYzn
3VHRgcIXAEVPRuZWtjPCUKPiuDm5urEXVOVYXolXBrMAq6ZzDLuQDx5uurj0tMNB
QPUG87LJJ/1fH7wRMpgsy5PhedL1O9qaDWWVFtfXoxMLvY4Qv/Afr36A0fQfW3dh
cyGB1pU2lKyZIVhkcL0XtgVtxQu7tRUGEn6YE0DzDvE=
`pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
YAeqxxj1TkkJuv2DQYjLi3Is96vtW/sMyFPWhiFTx+1SU3i9gjytI1YtonZf9TeA
fBYA1Gif8gkRAduypmHohfamaK+Ej+iQSFis1ve7VYsCnwKYD4VCjPBcH7egVYUb
mYXfe13yYsmFygJ4iJVZQJWEwfelyx8Oo/yb+jqgDRQ=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 5948      )
myoOO1YQMm3vpgPVqigGCuJD2QCx7bNHZCt54Z4NcUmJDfzIg+6WAVjq80UnGOFW
54R/D/fyNZQBv3RgTSN0/xoElbFFVcoXGrObiuw4G4u67dFqndqKJFKidUU8aMjg
Xl3JtTnBl8i9X8kw96gZmTRvlvUTaBnKRTYqwAHCO73YvTnw5KRdOvVpw0kV6De0
ebzlkFE5D5+po3g9ifSG2jTDZ5gjm6b6haMnYsoBigwERA3lo7FL/uzVfdQDxrum
BdgvTtZ6uEfQRc0PR8YV3HYlRKG1TsqgHuvOUApEWNNv0J5sWyJele1dYrwWdlUp
Du82GblttkJFevxyeOfOtHxO06u2KlgtCclVJ75H4/GL1mL+mGkUW+TL7o+Z8BlT
uOXB5YhLzFC/CnbzASsH7uj3Toj4hqgLufuutx6gdec9rpZ5DmZxyil5NcY8hYOD
ggI9IbPUYbnI1i4rT/+8yKcQUongBIXYXCJbJvwiucwzLh+k6SIpt2U2QHgFT4E6
vMtAp4ugc1Uf3o89hqVPD6Ok8sSDE2Ws98eU/7iYM/oAi1oNghYo6sA5nGhnOzrq
kLeL2qtuXGdAoxg1ihidbNjXXpyWEtm+/mm988Z7C+lxcQP+lK+3/5hldKBpQQ09
zO+n755fQSrE3RWpAANXAwJym1LlHUlt2KG+G+mshLR7qObTeh3gZjXYUxzvuMc6
VrYoG4nAh8+iQ0g8lDAuj7OJRmXqht+aGQkQ0EwoMEL+wTF/2+ZDXQOs3BpMbvKK
PWoRxwr75Af7QiTug4CMfPS5FCsBMrrZgqRUsrtEM4dxjBY5EiFOjOQmsKSk+a55
XMiOEheG0GFhKwLi/2W5x8r5A0ZXCe3UYcufp590U66CZ8W0JrMGCR8R5EL8R04D
srEZ52zz72NQF0/p3X+J+3Cwyb6qDMcu7mCL3AkptuHMaduRmN6uALVpSQ0O2dmR
kEjp5FtsDPyvmWtdhePup5r881dQwm0IBsmZcbt1jA/AiUI3DPKhO0puAKxXG5fH
8Us3NQrN6AOUHm7GZMphfgVwauHLVr3QyUL6J60SuPyqejPcbYP/i7SnaIpz7vF3
ZNQttAerqFLYzaDySHwfoc7iSuwiBaIq2T5e85tgsx5AK+/yWgEgcn/ujROp5+4b
vJRit5rXaGd69FbmtIkW4SShqaNjyAgbzlUN12mGHMJWd9Drw+krmr1ABfJvCZ6F
QFohaZmTtI3YFQZ/mZK4PTU3SZ1cDuoytbbdG1JnAxSLpHGS/gHR0ON+vYJk8XiB
kbFdPR3TBoxh/u0Qs3E9+RDGQIKAwQjm3SYR2AF3tV50IYymaKFS6T9ke4OP0prr
8QOpdOe2mOX3K/FmYO4NEFg8Gh91h3qp0nMeI5PNJQ3FHCQej5owZZgyh4MjkFlF
D4O61TRkU52GteHM7VlEvom92jkPo9eMF4RfkxnHknNR4naUFWvPFwik6sD9bRsW
/HZpZBSYJYvYR+cUA3Rd65f8rxiz8139bVTpk21QL3XeMDgfc8iaHGq/9UdDs/u4
6XAltdrYZvykDGHPCJBpLT7Uh7gVFrPgxhLCSZ02+4/CAQ4qaUfnkl9z7n3tl2Co
SHNfZegDYz9G8YWLLMi1X1Iewor2MOcvTFxEADp97dWFxJjomkzStazrwZYH/Mxh
Xvw1KwulpCMznNyk/WcEaAjZy5YRPpcsQsCd5IjAlOYTA68KKIw9VynStS+pbdDw
je+Ph7XWk3/LXZeKiwaPWJOc81WOzxYna93gH6jGvLfr1Z46swfvS2dj/B9RdBeM
z2JSU+Hhpj/l9fm/uJNeaDDBHsD/HPL8bQXniG7l01YCUVbVrFtkEWMQNHcZaO5a
GOxak4/kI8dLEWDnXfgBJ58o7QdV69U22bxySoHtEPKCgMTho3SZTM/US9jrQdDW
es9zZYJ5Ss3Va+lj4a8VB7Amfj8Hw9jNhKHrSjh3Q4I=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
GjWxycvgooqsSNV4JgLUoPdn7SL1XKzLcPcFBTYP8cDtT4LbgbKuWbFjZUIaYcwL
+Q3NZ7/DcrzNHExZqEydgMhVGtoKD19MMT45dRFJVQvAFcV8Xq58xckwE/FumjOK
GviS3VanLXLVMHHb+nVYJLlT4++QVVYs/mEfqxd0uCc=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 6062      )
LdxXQoi2Gv0ktNA2UUqGWu7V0iOoOxDqsSbOGNUXbojfK+6x/PCmjfBQFpVMjWWS
svI60guU1nYwBZczB6Tj86fqQUlmCGuvv/MgNKCMWAR90CQcXiAUqyfmxpcBeO0Y
iEOtRQlp3iiDMgCtbms6MYPxqV239RDb/2wJcfBcgs0=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
WTQ3pCTK0nTpudZOKvVYrnQKgjtHBJ0n5qnSd3xMDX/p8Zbm9ibZc++XuxakcyaJ
ODgNanKvRM4qCsbzEfJFM0U9wtNGiABaTW8PtOcghFuhXaDMjyYZofVNLs8OiFU4
VRHZzYdq3S3zq89dOuNi+R9nfaGDxj7sd4Nf9xgnXRg=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 29583     )
fBOfVoS4KNjuG/uGniVa+QDEpyKNswAxehati46jGkhOhSYR1XiBMkIuC3fXXtPz
ngaQufy45kmeH90El/xe9Eu6khN6G62LSIdqyChhg9M6YXb8RvU+5KIpev96QuMr
30Zj5AUHchvsQtACj7XbHGfjeiofsPli3DE31lMVEomPi9Uz8vioJWZzTZTVQrrz
fCzhUdBoi+iNal3hbANiGouqWs+urVHedSV8Dit4z9m2/V3pkQwP86LDZlqS4Eq5
aDjh6MwFYod5TlQMei4TFJDf43Up1e36+slBGtTA3Y8UD/qsXrv5305cZsfM18Mg
+2YzS1R4QJTZdhOzJgVN8ZnImLYnI+LIdW1qPtJWPBVf+/kCvxkJzrLkyN3QQHjF
jkHCX14/0XhGNJyJ7R8+SQ4OPCwdCVG7E6phD1CGVZV9rfNJN3fzm30Dbl9Mp0R5
sqwlFKDv2AOFQr6UCXXpWQhHoHXV+0rO/lphe1oINzwgybvv98J0xWY74HXsG3oN
74csgd1pXgrW9yDgIi7Lw2XnCnrU251Vyxf34wdJYvh93QOvXzhsGWgCmjWcAaNu
r7FYyWgf5QdcwfrmXc/EXGmNxMTvESRIqk0jLLBQQOUP9jIYPwC2bVNgDZb/m15k
2f5Bt5mL4MDyUR7Zbcd7hyY4EHxVTPvLdZ9Gwa4N5JXWMOFiuEAMfPdsIiYtopOy
4QOBbefXgGHfBpr8GkG8jiGIPM7/fY6EqEEQQQZcezm9UOn8L3JwKorJfhAMJOPq
6Cf16BwwXgDkYjY8e/pxUQEvVNhKyTVANewrDajGJJKH8i5Myk443SfM7moHM6Nv
kMXSd+e/ldUKpgySRXgxMsco9a0wZxkhB9nwkuIqLxRnyj69CEJqx/AOgr+KL85l
PQ+HU7JRcoctQAfmTxupw73BRxa3EzCO8bwCTS0lGh3L4mTyWVJWoLGtv2cMQSWy
vJoM4rqZ9SKoHoXgZUXtYMSYvfMyeJBcUiPAVLdeyuzgVAdB1hZkzu6TtWjoE3kn
VdRvaJpp2W2dY3e7NZO5/IytIyOpZeu6qZKrnaGGVZ1xPKlcv+bYpxidXExe6XQ3
l32zO/EQhTxh/FSKlBSZrjwiTQporDwP7RaIdD8TvVlo/3Auugj45bkY8T3/8PR1
6QUDBoIPh1duOEwDqUwC16r7QM0Q7EKuHJNrEyekuMR2VBYUcZNJW5xnDhoc/fRq
Qf1zQMJnePTMoJozMP+XAzYXzmMCGdS155FKQPlHMfgQ6NQt+tMevVZsUvGKqmSy
n1rPOrMt8T1g7tjcwc3NUBgV5HTljnpUSxZdYoUw5qsDSDhzfXh8sVzhuufCO8RK
e4srCSMRE/TFB1UksIqcPGD6TQLxKSVC1f5i1YLmO25nBEZwjeJbL9tRcxEoSk35
82L44QJ300rSD2xfsb6rVf+r1qyhiUlT9QnKk4zU3xcI9qLsHkBuG1Bbc3X5SJSo
fwXZOUJRsen8ZotJ5zRhFkoCAuX2WU24q7rTgfMTyHv/V/TVTYhrr2GRzJZDsSoD
N4ByJjdGVi3j3/5StAzLhQDS0MdhGHb8dIwJwK6jHT1U/jiyurJw0DfuV8WqXUwz
VqaYSlQ70Dof1faAlkQ6w9h/6jrFSMyIPqvIf6wZ9KEaz5iUfSLztiVnio1KXkGi
H8YPmYBILKuvGtfuK1tUnYfzSIAu0mo2Mc9/qkYwCGKL9u2Fgy+HmkehDAoGbd/F
0gLegJ62Z9W7y/fUUWArHpLogV40fMxpxz6ndJszFN+kX7onLQTSfCDpvfwa8W40
Y4DZuErglx72bNow0Q3yerhrr3/0fPaFwWEodaRdlBozDdApjGfOxI/PYq3+ebDU
lrkbAZ+nXHAb+EgL82L34guNL1UblpdiQPA4IYACGegG68rOLYoz/cgvuRLpoVge
Eq6QSXnApySeCd+lOxiFWKKFXVHZaxoys0id1yc62eGFVVqoOGYJL4y++om/y5Jl
xr1HqOftadiWAG3D6AvlHoFR9WSo3fk5CkKFIkJQrQE3VSlvzms7vsbvT82H1P93
YikAG8iB443buqyvjh7s80WvMSwViuovYXfHPFHzngjykrVRkYA2MRT+JtbgnW6B
gSlhkrOl+GGTyvHqzcj8UPb5+c8GyiMONMfL/R/qYiAE0+Gwib2VvPJsPbPzAvY/
sWmiLyiRSSohh2VoUapsyMpZ/IcBirxPGSTXxMGyYfRgs07VVi/MBauT4Q8+eZfT
p/QqZTqaBzvEY7iLUTpmb1KG2E3eA+c5U8+Yj699RBgpZXfbhu8WiL/8ODE7cjgF
VaicvIWs6HHf99aAHWpkDMUqXfJGJXVMBx5WPCzZUCk7sVfHQmgle6JtmEYfDTth
nFUedeuKgFTXUKEMYatSMPFZ8Z7eG4d7n8aKBKpgHGIpgKVpIW9Vh+gUw9kBZT1Q
MvMwhJ1X/xoi2LqgjmLNsnZBTROuNN2Jyum9GPMiLUtP/SoBkr++FSrQUlfJpHLj
T4KGOAhjmPobsQed48s6MCE6o0i+M/GFP2aojy37+FkEBAFd6FCO0cNhwgKDhFCf
eJP7W8hJtvV872RKZO5/TeiCu6b50GWG1rQiJvIT5/rwyOy2e8dvnOanzieMF6yv
PKJ26yTd3mQmSKC7fjIln2el625cjmfnJQ16VhEVmGccCYMqqc20v+rC4Swb2UL7
sNQjx+MEulJQKz9cMkZVvERUJ9NCCqe+iXPMqSL2/EYAlPIFVg6x1RhdRpbt717f
0nCj51wsc01K8yxqO00CqIah89+Y4t5R+YJp2c/dJtIiR2SDVutAo6upwRQWvzbR
0bS1P/T9cL0K0oGv6s1WJgWxP8GUrMeiLYw8x8zct2CTcS/t6IY8DYtcIbgWACTz
CfJ/RqGQSUN7WeQQ3rGiFRz/UYalq6g1WZJEg5QdVMDdTbLo9v2/A0PW+s8l+Zx3
tf6OOHXUticOJs9xmHw9ijYsPc632UOy+tHSS93lOhQJbPEiZCxu3d9A6wnee/cY
Q/kOsSPEV3+8DLImecxnxcDAfmbhHFqwZ5JReW9sc7OlBSwqkowrCuGQ6WD0hIfC
kFL/au6oc3INYzczq9IkBvW/CqfSsYLu7Hp8RIlQ2j7vQgjc2B2UBoT6w5HoO1Sl
vfsIo1vWP+7QNv1g+SiuQvplejT3bjrlYF9VuTVOJICLswQSAUQvsa6xS602fx4J
Vuv68V8aHOWCz7wOVtn1KstIM0WIc2Jd2cM9ps2hAWuyuCG+KZXNxNrlQPe/xAS0
XF4r9HQHezt2E6N2CesY/A5jBga9JChG4o/ySbBPusSiUsCzqlQvTjykPEgA28T6
jdGb8C20IdZDtgQCUjsJGZsYN3nxZxZjjKOC6WJiKI11/g+J3yN069OJMLQhtaxy
cncYOACvVLczTpJ5NT2DYXj6SvOD9z75NDem2uWeduex8obReJS3cYwrffX2yIGU
vb6nKqS6XgXiwpvi0AsCd1GEAAv/5VjUIChWJ3fgsO6I35Mx8X4E0pt+MrOmGr7p
gCP1bkxLTRUSUrtVDcIBF7Vu3gR4gsmdQGW+LfGH2rFBuURE5dxdnWT6KX6KQP8v
lu3pJdncI1UjpgPYDaQFYX5tG8JHZvoe45hNqe+JrYeVVMv9HxXtKhbCPcNhOmJK
JHSFvz6qY4Rvm6za7ekYVzSbCLLaZe0KZyPKG/pDf4JMsfoLSN+gRJuW1xJ9MxvR
m8stVnlqd/q4xMctafJkgUXs8liWHVd8/yzi8MXHAiNpgmLW49CVpyDu90VM0+ry
PX24VtQbH8RWcmG7Y2YDE76xRFCsLYS/dmtPom/TSsX5WCtHajz+ICnvZVWOsdpf
A1DvqTduv+uAEOivf+NXdq+gG0pjkafHXBXOxYCSUiNtvIQydal+1D+W5mk2SD2h
LAJN/MhhpvUTqql1URDVyofBlHBMQKS9B7jHkQW79DPLQJzFBextzFuEKZg9kFJZ
Zm1i+5k+WT1U9A0tJBVUWIkv0hXaG3PM/R09lI38OoeXn0OL/nX3l7ThQDJS1gnP
JeS158W2f71AGR5PkpqnytLU5qAOmPFsgmIIHZ/B8q4NE2brfAs8FdBNIAW/voHD
ES7wJaZrvSGjwgNGiTXLQFAtf2TDtgBl+vMPz/CqB06Ie4ytJrzm00rfaLrXtcWx
oij13n9hofo/Cn/aKilE+uxlWBuW3oa/oMUCj6B2pfUMPtAQGtxli2IoKOdysflh
gGVmdepjeNFSHdvnsHcTyO0E8kmMoSAzjZ9UQUfTwB3GCYMmsGo7sZBQAyRx4H8d
iV7k1jj43SxQ/IS3IX5GBPF81fR5lp1y6Zv9wYF1Ng0461YQQlxzOahfNTY1Ybty
e5jXIrJRC2t0BBW+ALqNl0G8xWzreDG34tCzVPxP1DtEGOghDp2F3/0+upOFdfZw
f2aBmw+4CQ4y6MVdmc3fsK+HHAx+0bDDGRLt5ElD7izcLVWNNKaRJsuPcyYmbJ1W
mRzDlRKxHCyFT4HjzKzGMkfnChD9eq3hiiAtbx8yofVsI1OnXiPFEiYs3wz1HcVO
oHu5Zpx5fGE/pMySRp5lLBVCtkNxPLKobl3UR1ZrLZcjdiHAoOSlPAP2/G6RCivR
u01Ka3uzbgT4p93JklU/zxEH8c3i5iMqYtIJuZ98GjAKvrIfJ37D1didM3DkJ3JF
rmOoTShFZnHUDHT3OtiFU4a+9WErqoGXlySGQzndUvql5IjDxO5+qC6aQD1l+jFc
RBb8UDxGxiZkI9Nu9qS+SKia8KM0taKtG6YJb2ivAZ7bge3f84mWVoHofUC1EnqW
RcLFJTPFokeFrzuQHBae6QmK2He/YphRKSl6seEWMKC/0hCGQHq8NwnpGGy+uB/o
chMMxfwEgehheYOek/cUTvRFojvEsitVjkfi/33rNddFoYBR3JE5TbvvLItcwDmD
H92GKJXBQPAoKquZcnltVb/IzDDiVOj6DIJVq22sHXNEuK8j0Dmd4IdgYepWKfMs
KV7cCx6cVgLyO/Ciwh34uBnC784N+XxJuhJ00H6uXkY5VCUa/GjLgSphehgIACdY
wOKQYBpfHkA/VcCnPBy/goCCDjz16hb7qVyJp64DE1f8vrx8IYKosVE5dVvcMZa6
pnSGUGP7aBySF/qmNDT2LbV4xGpts1H0vF+vT5FqXSJ18fPlikHuJOA0iEiRSVJa
xqX7zlgXMxxSwOMRtUtx9FuRd5zmax1f1AJLoor2Aln2z7OTDsKP0PbwpMmMZbox
hR9mMhpER8i69Ix3eUCYQMfnCF4YW/8ur5wb0JLLyQ/CukTiEEgkRr4r2LmNg8dT
z16Z169110l4/bKQofBfUNiJnoz3HOYjJHQpkOaCN5oP9nqHlsgvT2oRLe3GqVIF
uho1BMReLCP5kjDv+B+hLiAmt1YzOunr/t6ddX/LyHTDfWad7lq3RQNikEDFQsnJ
L1AREh2YanUPhjX7tfSo4zsW++KAt3A79XnXO8FkmaV7PLDD/wx0zExyJrCK4+GG
TTRfkqfRV4f58bUsOoIp31aY25NMqIQqxCbu9nQMThBh0VAlomPpDVWO6qpvWYjD
16xBKQcFPRtBpifHvB4HvMqtosf6Xzraw6F0sO4RLFB7GlGT/ocsOtbQBUIxaxFN
8UgaOfPHXu5w+VkI0XalJzYPiSGy5D/G7/IEm5z7n1rtMocILakam5yFMq6T2xaA
sS0m6EGQRqihu5GQ67J6Vp3uutJzVCUqnSBSfT298JAcc9+9T479gJbpyE1BRVFw
K32LgQz0Hc9Hehj/6AdA3EyHazRIkT+dQI3Fsu86a9eKAxeUSRmWZ7SX12ba9Bvb
J8TfN6g4QEnhxHqKbaiY2yNT/Fz7A1b0zS1PhsDbL8Jv3MQI/ODAxNgItQRO9sk6
isQxzi8Wnozrd8jHW3SPNbIhUe60aXVO26ApnJchci2v/RklWi8nx8+G/3y7nwo2
r5SK40xuZ4O1B+ePSaBGmL2Ne5mGGo6ByD4+2l7v4jRMR5dhp+kFEchWc7t/Cx8s
4GMCkjq6dZCw0qnEBaclsFwxmL7Ic9mLjHnI2V1Xawz0SQlWbBv6/BC5AdXGWWqH
gu7J/u3UB8WbE78DFDZmDKlq95uupHrEZvJDcq+k4QWI81YRcGbbVhBiCs4uK+iE
Rt1mdYMvIQR5usrjanwMMJRBKow5Rc3asXTwLpkhED1orkoKPscHkS7xrNknI/tW
CscYPGNpDDC6y2J0gDJMp2ndJdKR5GoJw2RtiZOPDxJVvxhdggFz/JLzRE6McPBi
gmugTordAPAXMivvxehZTr40g8QPhLHmX6sE3IVBM4kEYpNhRRC3zVkBdmb5e6W7
pO9qjPUrwbpBHwWtGkZtfqS6AcE4tNuw77Gennan9Ul8cITe4vAglCK7+kKSx8+M
ticABjF+pM+q/sAg/6e/a38o76l3moo7kdnCeF5djHdKUpPJzNJVC3h+JWSjf1yC
1MIxs+yVWzoSvnLuH//YspSp+Yjf8kuVNCtdghNXxmmy15RURYTKKCXdyrrqTrBR
yqET954CMb/SVL2hVeKaSKrujgPcv7aj8B9arIdKGohVrbJKi2RNo01DqXktHND4
6uuy90eZ1EqIL0BqmpdsokAqI+eMSXkbycmooivqsagGY6nB0Z8WWEmTvWYQWvoD
Hl6prZiFUtLVk7v/lbQKsc286a5G90R/cethPCB79BQCT5GRsUCARCh00o+Dv7GH
3PZDkw7YSW/rCLyWgxIVrDFgoMMfTyjvXna/rsyJmwN0/WYlnhzZqWkAfTJfjSjH
LusUFRnLRJ7pia+IBe4+ZNTmQ64yYPlPqawxULZC77JgUDXu0VnxnS054avJouKf
aT0uF6v799eJhhU2b+H1187Ta3yg+Cc0kBD4Wy+fLubAR4Ibruscib/Zw9U+8m7k
+gDJbki7HUobyu7pnXHdwxzqR0kPIfgyPDetm/lvJLKCKPrBwpaa49eTvIHnsUMc
1N9VFqzn8TbjKwcwVPMh8RIimhBanbg0X5tyfjyyvKqoDvvgY3L2OZHvRljSay+v
UtWgCfwENH+GILXPBwslkUpcVcWc+Qdfveagr9IGj7gSH5TObiY1uzTlbe535LEB
Bz922oSTEcvelvVoSL73SqBMT8aBsrg3E1HAxcemcUn2zogjzVVAgDQ4M9GvhnUe
MJDkqM37WekW+o1Fk8h7I6nRFSyefOkBdMxuaJcfwjGmTdPzjAAR3ai2xNLIW1uS
QHMXw7/W973ohxe2dPiTTPn31nnEGUzVHGfqW+K5bOrlbU6tBhuu+fnbx838Kj96
Nz3TQs+fMpfv2lnOUGq0KTL5VCLpR+nvPim+qJfDIYhsI0CwHxrohz8AL9iKGdu7
HPXThJsXxfC8qgEFk+/ZivaQu+tZ0Ch9YzQQXAPNe37/ROg47JsezjAm9R3U9i8Y
FKeP42xd4ZMP+3T/kcJAg2AdYJRGQ0SE/ZNMT8wZ452hJYw+Ya8djZ6aFSjeBK18
eEkc1g0S5Dvk2SDSEtFpWgbTPTN+dCeewFN9QhZmLP4ZewaGld7cmX+o9kWDvZWG
S0tlUWFK0gCXmN++kqhGm/+NsXKZ1c7L0D52Kwz6/8c47+LPEemdkTB7wT2hYo9t
QYyRowrWP/rtQ189RtitNVLtb4wIrNAtGfCtAuEXPDsMfposSqPf4qm5jAYmeOaY
ZQQbbXgm4dF+rGBXjwSiR0KfxSOifDlUXKbhAAZTVZRWJRWudEsv8najljT4QByz
Gsicy4aHbsi6golOtNb17H0NznCQ1a1M3HCFJyn+mG/+yn07TE/nEAqHChKS8H1q
pVjaWNkc6cC4kxiooP4iVGQc8SKqeQJLWNf/yHgH4AJAQD2pbJZlPBGlRmoiEs2m
+0bkPiIHilw6ATMS/LoZbrLsw5oOZdJ5OeM5Gi37vgC4G/umfjEd+Q+o/l7nMTiB
xOysVyNYTNweOcdfOoVaNMcm3YLXSg+oiZUl83gwsRFj/IyBnoHUrukEmh1SZOTA
nxKEv/vsqNwFJteSz/DNQk8Q9U+kXM5U39J0KQD1QXLCEP/ASG3wsQ93sPtLpGte
ajwbbPQx+F1EbAxRY7MPfrjE35rqJqeuvXgPUucXfTsKikMjwM4M6tbEC4X50//n
wLjDOBr6U0QrLLSnImarCY6iJwyEBcbUeO8tPDwNAfelR3EcKotjQ7N5glpvYif2
Up5D+atz7o7MTi9+z9ydtuglHFWsA63PPSEyR7xQKI1pQ6gSQcv59q37fYGXKu0k
Jbds9ZegXvJCHgVMrSG4AQstd83jXem6FXnLtbTgRSuQdo1xg9DYpuNAoGmmnZZS
p4YC0/s04OemfMHRsgWJ1jPsfEGx52DWvFZZYv16sAN8w2JtlUojq5UZHr5UwITh
fxSFvw4qQHt9D+gBSHFL4SjbvL3fxqANsEPSTUU+d0VJNEjMwOo+Z05KT4iy912q
w4wOXBIWfBfq6UXvGkygMk1G+ZVOnRoCGGZDl2q/DsqUD//NkcN+wwS0zNx81LB/
sP9tVWZ5uHNCzidt8xLUj+UEipQjPs9XTeZ/Rvx/GvmAfiSEami0q4rwN8xgE2FI
yhkW+PGwQQ9HFt7dsSyL6xPanLi1IruDBAzG8QT3hJ0zmbHLfshM3Bi06By1vNEC
A0DnSMjdCPSuv1bwJqjKS3zliz8wA7m7Bgqp0EEgJfwPcTck+Ms0DMQMvLxjcGoo
zo6KELUaFf5kTPIpwdNsnPv9NELtaHbco74mGWvUT6mf2NoNc0FFdlIrJ0RiiwD0
BWY+dvIMQN7yCiV1qQlwF7as00U7rx1loQShj2EBr5QyBQAWgSaaMbNHcThR2J4K
GW5lMrv5H7r/X8vzOrU48IrwhsH8YhrcrBE/0PpPDtppoyaRaTAekLBjbTjSVm/1
ST9FL20n06LhElFkZu5RhVXlJdoJ29q8kG6zTLYiBaCaL1MiWDzsplTd9N/68QJz
9FqAtYjl87rfU2t6VZwmtTcq60beb6DdbSiSAYnq7oBak83Jy60Y0jH2jrcuVcAg
WAaBsAU5VYsB2px1gjQyuoeRNPIL+7KIz6cH0ofslY6TZ5YQ8NU6hghHbrA+7g/t
rnKBIAbNykS1FSJjcGBE/FaAl52KntGx/hpkcOkNwlPCuJeGK4GbvE3QnTujgp0P
u15AKKWV/xte8MNMcjU2P5V7ncx4k0Fd7dPn7fVDGY2zdnDBZzalWx+nRCvvAq8S
WFrLrr5bAeoeBsVuBo7EIC9IyjA/5KHKG/irnR2brEnzuKrA6yEQkLdlKC2aC0FU
VNKuZ3AF1uIe7VcahPCALSG1EgA5cYvuOqKkb6SXkHvdbLlGaxUI9TTnAZtmdUh/
5bgG4bIa5XPnEe20VM9XEdM1gAFfUvP4XjsY0mYSeYP2A0hzLgLFsKM+yillDQAL
mF57dUR7qMjAs3PVyMCl1pBw7sJnaDyDlz/NFHi7P7S9mRJzy4EaitG9TQQKzuvf
hiqhLeXRUGmhunkzSDB2zwsSXwFEDj874s2KFKGFTc+hMg5FTfpABUTrKcv1azum
xIvQ0AHHIlVmnMhAxMFFSeeCk8OkitEZfwzsJnrhiQnI+gLL8wlvJsBr7QpfP1T8
109x4/1WajKGpI5E/1ltEiqpxXH1orhcA9UcFWeuptPNW+bFU8pSBdJFO5E/erC6
Hx8ZaVDdtIJ622yAGPD/1Fir2noyUrGgXvCpxwRcj91SthkBEeN0CPb6E/aD+mzc
xMyn973n78/DqZsIJzdZGOuqIPKvRTKMhlppd6eToxWhjRcArZUdiDOfHzxkoBIC
1Amzp/PZXnm7NjAYtdHLZL3hZDGbc8rEN53fP+YqK860+v5WlEU/14vqqrZvKzs4
dvS0AaRDh/ExnjQeqviNkWrURtwrG0y6a0TDM80vXqBwLBIdzgk5xM4gEeVB13Fd
M8wdNxJSKPNEqukNDrEzqMbu0fC+daldactlJDxGn9YSsuFfBlGUvZy5QwaQuO18
a9YzJwPRYMjTj0K+burgtDwgp0QmtLx4gRtid3fM2MlWe6ntTh7/w2AjtgWZGEWN
G87qmSn532YL3OKkobkVh54nxQZyLiUMv0ZzDJiaDmEADMx2ef232dGkLGXViyrN
/6gZk0XGMCnjoU57YwJL3awxNaMgooFRm0q88jgBwyCXTJa8EB+s8PN4jhPy5axl
vVqQ9U8sIluLACfnA5TkTdDjFoux2d2j3cKPsNYX5HdBbO+e1eJaaAUXcwPSYF8P
GsoV8pfsH2ayqs1MOG0tIpIQHlC3ttcQMZ+Jj58LO+bxnw2kRNfp7h3fe4QgIgo8
1mTLswrnKQXw9YT4QJAHJ5yyGSbtAi8RgnlvZmOK8Rb3zBh5ANSG2xoH0zzVdLRM
MnHvttgGAlcw29dem+z0GHHodtm9A1QUJwFsNG9+DxG5zc2ph1P53D1ri0kJCAFC
2glHc6As/VlIrRFiwiEPV+Ta2aHDAb7xn56prnnRVxsBstLFlGoE08CsGNV9eC/s
tQkdLa7bQXXe0RnAeAvzFZOY1aRwOAyhtDAVKP6vmKguNwWQd0Kq4lZrmFY0iBWX
J89TictL68QgGGDn/5iwRlRZTBNVIC7ymskJjPdqMzE7YpIgRIA1jHAVaiDsPsQ+
YuPStJJtpes6lYGC5sxtIiaTxESo+aCvTMGw8dSYywWwL4Oycnxwme+0sak1Ikxd
5P318o4Oej0liv9BWWRYlrNa3gsBXHx+7oJokI6/+trk3ntnW5Ou0TjFikMUwhQj
OkzlPVKV6vV2Mydtw9ElAOenWuHfrF9piOv+rfsV5UDLlu5pcUlJ34gUqjMyCWWX
+9FoR1SvHvBN+G3pl7ByFKPPZ0t8f6WJrz85Szv3X78Eg3vMGvoE8EMu54w5RSRN
WyJjVggBQBZok/pzu8vTNIrh1930xQ8+W31tJ97ty0XnqUJ+UmTSGVZ4oD3G/Wce
Z96WRRpYETNrOtfXCfJzGee0BKr3p1AFC+YNPECuOLG7EkzpSlSNs3I/IztlaP3L
gdn4XuLxmPTE1cBtUS0sq4gr00nebIYvkV6srKrBp07YWz6igXXSXdH1YSvWBL2y
mYMBEKUSoNwcG0URCx0iZ6/Wr4NkwHU0r1srGvdlJMmqrt2XvWYTON+HJ3V6h4DP
8z+uxDVwjoCeDppIqpr9/d0b+aHh2eNTboMZFia5+fTx2VSkwuyEn+g7qAFIBAbB
WhWM2WFqDg8fWw48Z795ZdPMyoI8TMw08O2Ff5dTWM+V2qWoNjnSn/NqKonOxDJU
NsNvUvw2tIJ+nVGJ65eOlJ7zAcF4B8mxI+PksDXP/n22ALdk59sp2jiXGVDof9SG
MDrs9hH9a06mr5at+EIldOotN04nIkOhn1zfhvIGJZUY1wx2ZJQEdKuvu4Z+BKOV
4o2OzwfRXfMMffEwo74t7UGADtBkPiGYoCIPdcYEfxa2cZ5+WA0CEp1+7jNLZjWF
V5ld+RkwVofOw9tD0PGB9LSDhUPd8Wwvz7SJ75EfJsJIeHUmLiEjje4y6bW5K2T0
Py3M/kTqWp4x4WkjeqxsippPTuck39xyCYFhCGWt+usrt/1TAyApjtJfrMQSqEeD
on4X+t87H0WjVbLhp47tfwWKelFzfeBt9XeWM9EA0koKndHeDbblw4Jzs9pnR3AA
yyT/4a8UuNJWEGyOfhtJD9KF7vPhogY/aSZR5wOz5IKm+/qyoUIg3/Sreq2dPPmP
A4ijuwxRQL/U4Qp4u7F131RdAEkh5+HS449SR2kXcjs3HDz8EFFfgIGaUWenaQWq
EDHpOsfJtUTmVqqtkj4/1Qw6hRqmBhQmw7cTZEH2mAUw2+oVytAFE0sO1qWRjPY1
iE7I/4xuVMhKFfALR9klwMmBHtYBN/2QRF6R8oQX4DCJDvrWgnxjz8CJcRTYmeII
Ho9M+mliXgHfOSnTjibQQ8nAVYxQddsG2nalXESHrP10w7rfsYYHdaqrzRsP0PyS
YNzfOxjg18MHVOxG1fzWlN+JX6S76C7P+KKtjzx5/8O8IjzeM1cBSsdc3nctJtBI
Xn6pH6SVAkvnmLJDNJiV2vRxH3dOW33CpB8KoYIOiUX9NthHXM7j3ewP6GZFUDzx
ESwnGdfcK1sL2gw53fW+28BvZoHiXoJkRKB65MP6+2p2ldelCnqf7POzCWunFw2w
MDw0qjOuHn3SNi/kaHQIWc5DXVG7W1d+TNm/bLfJyBmRzMP2nS8iygUl9a9Roqk9
1/0vQZNchUARkqiBMF3qsVpMfdnJB0CjVHqsdudrYxF+//Y1SpAyQ6YLiIsGz21v
K72YSGlRcMpH9nFJ7xR6tJv8ktHFgp81pmyIw4eV57B+obFPQAjhSqr3OkQeWPIn
x2LAQrzJMdJ0l1pHzhem9nbIcjel8nTNLppc7f4BAzD4HuwfiS4vFtcBu+y9igSI
J717rzONxsLa7+X17XdZOImOgrAKaE1HPioMGsjDKAJ5AkFCSS6WWV1nIoVETFXs
SUEC449dGvSp6QhgBRuJfC6LpBPYhOYro80nthJhkprdbMc0GUA2SHOOWtD+TlY/
dIIX+rqwLYlMZotmen4GBUoAhwbl73C1i0O+hM7wYBaOGxQWs0iFe2odsnKladhQ
W/kYm3hatexXsK7wqgFbfIGM+VYi48xiM2s1CE6pNFo7VjwaqeTJA61Bgq/YODB+
wmoqo/kmatItKEeHHfyRbeRTfOQNmMkE9mv4TxiFgyKDl5jEpydSgL46PhRP4hfG
2A/ysOq2g3g7N0RqJdpO47S3ITf+TzKU4PHnDeG9TE85f7HE+oXiK3MasQpeoXgc
jaTUDAHJn9EsUPt0IhdnJLI97sFYZft/6t+EnaP59PaFQCiP2fpv+frVJ4s64s4E
Ld5R27+8sgu8fFXzCqElCOUY8wDkwzyrNiY7+wl7QtOrqGEbu1zcLUwGE5QHOiYT
LLhQuPJeZqDe8CTr1f5yYNxp7JYynvNfXBVzV3MPcDKoR1PLICv0YP/MjDg9c5NZ
YuvgZhEuAiQ6XO9MlDyzL4ozA1YFUIjQZJoNLCxtMfKjTC6cKhy3EbUuODlMQoFI
3nFIHVMCrqWOc5TxkOt8w60rU5shwtpJGYJ958Z5Fkmz674ILDaHSMyu0AG8HPbd
HLzcrCaPfE/UbvWKh+nNDszE1KgVWdjNvFktsAPEJWtqpgmR5b2a+4M39NUp6D5c
O4njjEy1EqhrOzeo3r6Tai12Yibe+gVl/MXvS0k8+S1dE/mOan4UR7Ov4ZV7QPRm
4upW/sONSJsud4IguCOjMOgcF8EwlVamKmN/F1GFanxHjt3at4Dk1Pcu9wJzO3hF
m4y6edo7zaYvrC7KhVbLIeZCC/TTCVmZJ/6UbK0gToCBHaucxk36A+3X2H09Uv57
lE0/hFGe4Hb/sU7lK3LoFi/ZVRCyA+58J/5zRRL8Vo5ev3VMkjX3oggqxuHKoXP9
Fiz+EAK4ErMVQRiFlsfPf+f7ZlCzD+wS733VAMMbVilKXJYa4d3R7ePT8LPQKN+z
dIEpDqShQxqq3358lp+FfH6cVk6Z8hYRkVJLFglFT/I1mRTFcu/IojMexcR0EFDM
sG7oRoGQuF6tp2f0jGsm7hWUPJ7XvNJP2MOwq/j00GnS4mc+J5uWqIUoxTn8SQy6
kVBUJ7VCOa/a/B0cumTz8T2OxD3ePtVgsaRpClI71oO9bry3VQyNRZloBZvVhKm8
on2M7D380/NNX/J1RXrrfJUKpXgNu4+6Q5Hn+mMym+JVIzs/jI4LMOZDoynCkDna
RmEmbeZsARFXraC1qRJn7ZL4zAGTBVQdaf4xuO4AfXxAWADklGnXFB3SySJhb7VR
gvSjol3Jpm+28Vsr4CSNgPlCK4ajQNuP83ZhFr4dKN4RZHyY9E3O37drEVEJxRwG
VhBEOEbk+sYXy07RRIyD6EymUJZnoD4KvIKHq99c8fZIBaGeSlzAd2cTtWyL/uKO
wg7dee2xh8i4pyTGY6O0pUygmP54mWOAhEFw7NxZNgfiav9oy9vg5XIpK1s/QvdE
6ihlbwBqEpG1K+cH/rWTuukpmD8EK8YZsx0ZxcW82JUpGEq9kVULB1clvO7Y4G4r
/jKXUXztv/Kw7JbpnlupKYnw/xbiEKWwcIVg53rawk9L8l76W4BOCV+F+qoQnSYO
UTHeEXP+Irtr/Jh6+7JGr4ZXgEl0Py1Uvd7ptwmIOpQT1XNUgUmDrU88htiT4vfM
6l6zvp0XyhHukqhYpGUdMq1grOHLl2v80xImqAiGcC/l98tCgBGfvYfIVjVyGDue
UAnUBDnSj1cEZnqn/VdXcJ5rGOk/sMvYngUIQ+n8lAKiFOsX9/jj7NPy+uMpkdB8
puhbT/XYQLNd8ijpaaJ7AoigzQt2H6VU8KKc0SIC5RcBYYL644JrMps1rxSwFn80
nzTcUA40VHX6Zbo3hz3c0Wlszi9qYmgMreJ/HrcUW+US12ktaXeP+Rs7q0H77LMb
a4l4tMXa7iG69Xzif8acygrXsmggCUgmoFXqVtNhajSuq9gUh55UTOL1u3j4uio4
zZo5BnSEgBhD+bWKQdHvoJkk60rHhMxzC2q2bfBwtV9X/zpaMMAiuyyFJ4TtoLds
5kP8y3+IDjLrcAd0nD1zdrOIOYvP9LUaRBMxdp54vNC0+/CM4R2mzvc0I0YaDEhC
AEMCD5/RnO54O9+QsUZBw1pAnu2r+Y/wcGMhKKyMalsd/+F8vBTae4lSwa5V0ANS
JnszK1i9OjNhPIc/ruwc/7vKq5merBNJgbJkJOTf8L/51R7gsDLPB2Sxc268xxn8
C8ILmMxQPi4GQi7Fb59tnlqOEvteFWxyfIiOnvbAW+Aquh8enXDZ9O6IM0w+yK0f
kO2wAaHUx3ZH5FcaqkQ4n0YA7xmnLlyBeIESPEgptr56+Z7ZVEgsM0bXqfbmFKX1
KoIEFjz27kpQJP+asl0/t2YctkRjWFEzUy6BoNWUGBa3kidI/1HybiJ1ptI/nWyZ
NIOhxAOlFRtC3lxvBRT2Z4p3BzwIRVo/ECdYXS+Ag2ejvSxa6wMU0PWM5rnBg4W2
/K4q5Kq41/i6bPXaEHEgdh/AIAEJBE/qCcpJtZ8/FmlYMMaMTvVU15g2AVE4As2f
2bOmeS2Ao0n3TX+X40sFwlIrXafBD2MY1DKkOX1/YDZ7kMAioIVBGv6ewFGcwKlL
+ABlsOt8bV4aTsMB5jmX11Y/tlW/SW1A7Xh09ysUtnP2hTvPzTkFaxrJCx5auYHt
BQ2CNom1W7Fh9PK52ie3H5bVJ3gjzinx6Rvihpa6ZcwK2+kWBLncfK3WMiqrvckD
ZtQAouck0LtoKk5QNYcC6x++1Vt0tIWLTuj6o99E/DV58g8DpWVLaldvgzmv5PrA
auX29Ixr4zb81zuy5/g8QVx22GSIo7tvO/QIFSY807QM855DtqznlcWBZ2NhPcuP
mA+kwLPkctnmN/dfldvW5ouRoCiy7q9hAG+r6fFFUszWCN/6V/0IzpIat4Biez/P
TX7OtxqdJrjKk7eHdM1ROUUAljwZKBcLiJxPda5LMkbvfgshLK4CdFzelw0/pT69
q88+gKaiHvvBRKAh2kkCWnAUmDJ0eOS88O1FicGK4HqX5FiX8ZQnwLNtHD5GX9/N
ln7XGRFD52bM8VUt+3YOYMibURNAZi3UgB1zbbwKZmCEI4Ee4odOJxU0F9fb6LgF
WEMfRO9yCwTM4QRd6Q55VWOZOatMX7WHSM8HETs91Dt9eeQdnordAXPb+0oyX3xd
N/R7hs8/jWeLfP1cLjKJA13fnuY/SvA3idet8qHBG9+lndfhjHfZudZ++lphrwRb
lEcESfE3A1pfxDb77T5rEsfgakLQFy6VttTwVgpOVyC/vySoZtC37P9iVgMHHjw/
dTuH7LJ3ti3C9PNWePfCqAsXWEMrjQ9RT1e7mpzgS8x62QkMCdfTGwpLd8H90/oe
4GhWyPml43Cy/SiXoGSfhXHhlxVVXEVEfn2h1H9gtxg4pQdr/UxhCj2i0msW0sEY
pSplGnjKGEHOMcc2aaQ6O8Mf8018rQNn0jOmgd7Xgpk4G5X8D+UTgf5LOE49OtgX
Jew1tzJIYEtcXnPvsTX7RzscRNkHBBTRXtlzzQ9Cdn4msmNzWh8rTn5Y2Zu5Z1s/
HK9A4JdMtUTU4pqfDACfvcrr5u4nDKSiOVPEvvehoqcATOsa2g5+x9eHuJrqxvAQ
E6J0aPEf96cI1vym+cvgYbrfOQ8TJaQnN0Hz6UHlI8aLFWjbYI6a2C/jirzGp0TD
M5fZCLfrOP0rK4dldDzFATJW/bbdYlrHVvI8Z4etKI4fUmXDdl1pHFW6gOAyf+X1
OI1Ys/p3AWv2AwkviroDvf3DW+395RhpuP+j/KofiPAk3pPjwuzx5iGhpnzGOXRN
ioDZGAFV/N6A5mzizqOkTN+iqq8VUzXx84+HJRy0Cke1PfEbbwiHeu/KJ1t5m6jL
8WrDvaxQ9CFIhHuikhxrDhacRTECkVkey0nsTYdqwc2FVYY1K2VCwSQOsSOcgR85
Nhf5aYwZVhrdnYLyia5POd0zNgt5HgKQqcdyCi6jGg3VhEwbkZnws82DiL4euN1t
WiRL45jCgt8k+0NQfCGTyRHKih24l3jPT2y188TncXcDdY5+72FAv5zEa3K5Pu4j
ZXrVE6HrAM2UWRsaxl/jOmk/C6iklJukT021NXhuvYh2y2LqgvRlVEGifb1BGycj
mItBr4IbP70WoQdhiM8PguHBhEe8J3ID6JIK4uLvgPvG32d3yCbc6x8LidD+z3e2
DV0P9cH9YTb55Ctbxqf4+Kr6KpkzfWIDnwIIkFDJTXzhywWCM8rctlxgcJv42Ock
GyGyvjh2Y1peex3TyJ1KeeUgqoMXfrwL0kTTpTAYG9SOKHWbDpET9a6gbM/aKJGm
chgaoHp4l5hAMHALp+evKNvOaseIxg5drimvgvSIvpfnWX3QGVULKtbOmHhijwjs
V0URuFj09+FPwMEk6KoK2Gkl8XQ0Wzwh0u7+4XP7QDkEt7lrgcTQOkstD1ksm9EF
MqoCAyMoQJvR/j8KCjuG9cKkwtKci/TjDvDiH+rEokpJyB8LFQvmQZt6oRBZVRsk
u0juAWnyJn/G09xbR1fIa6eqigii/+UZA0ERYKwKaioVU5K1ABS9IaCcPkuQ3J4b
9+SIB3uJYyUQwwE0250HWLyGzdhaZcOMUj1NvulDg3DwfU1MrQ2KMw0DLMX3tyYE
6ilHwr3VxXreNhWTshB6AT/0GTfZAS1fe9ATAMKaqt4qB8F6GKqgc6xU2lRQLVWp
F1kO03Vm12CyGF8njbY6mGd6G48hf/n2KlU1yCm/VvR0fQRdi6Oviaf4JcRP13sS
NKCBGK146qO4KMe8E7awgYSpLS3p6MDSX7fch+jA4916uzchXNDZNfYazvpnjFC1
bLWS3nhqb6l7s6o/zPvLRHD6+gpEVMLshEJ0Cw3FmAaf5ANu+Tlf5y4sr8cQUJy1
k3uBkZAw2ix/uuBYNpaWD6cg539vmW4JDTsqngX/jFvOkFdmVH0E5RM89snr2wK9
bcl5h//+AVi3EOX4bt/n5rz1SAuG4U432sHspDMb1G5uy59VAasr5PxeGFoQUSPj
Y56WBucTV5T0CCo7HpZX7UJYz+BXNboff5G7LuvMdjbhu1Ot6uuRzCDJQTW5SSch
V6W+zNpOiEH/z9KtLdk+RqM0Aa5DccGbeDXXDiDIHRgtn6uDOejdiRXGmmREitvX
CoSFHt2JjvBN+e/0QG95Kfj0BOTGw/uoVwy0gCtRFqvzOJUjbuXS5+W5xcNhy0iF
36ln4rGuTEtVCRaW8td0c6eKq9y9jCmALe5jFztJ9qSOQ+oEKaGz8tbUqw7aKjec
qp6XOno+TFDPJsh9Z1ynpm8L23KE19sk5pUIvTluwDziqY552sdXLm58ZJhM/jIT
h7Rssuwm1LNwJHKFwc0NVNpoQKKhSqoTqg6bKPrFF+ygkOFw/0tkiaHRKQuWNpb5
ko4q0LrBdyyKdFK+G2/BaFHvv/WBfTUNTwFryzAfmvHKOlYI87kdTd49ypvs1XXD
VV1+DejCJb1M2pFCALOiBIvdZvotmkn3u/QLTrXsAFY036lE5cszLzWYVh+noNuA
EunKkDjvRkKeloNDRy5pW94c+J4e9VwB/9OEDRCbFhUSqVrKObPJFuhcsbOdnkpM
VCRu6RWaSHZtwwrFYykm/2pbGeQOl9XoHRvN8F52rtzt5as9Nlf0Dbhk6I8Pk87g
SST6Z2psrS4qvgRvck5xVnj69JGN/gISSbsFGQsdKOLY9JOlB+hro5Xf3S/A15YH
iJhztVxpWFkkCPkDwQd2kg107ztmfYgd520u9Tpq15179NFI0dw3vhwUtoW6UgXn
W+zt4aP4A+b8kbrQ+1Za1eKR83Fr/V68A/B1mgFWzlPBv2OXr9aCK/K61NhWCRbn
Msn24x3zL7GDbT/N+gRIXZ1R0xka+lZ+2++AEDgGLNRXM7guFcs39BLBrqpRQrzy
7hdEX/e92iGxck7EYYmvDfQc2/9kz/d5hljkhp7hf+VGl2EtEGn26TZy/+0D1WSB
BdBDwiNxxIiWBS3UjI8GGjlvbCcouheIUlYgpYXxPaMEBe+NR8IWtBon3rNXaZLv
DQdj5BhaOIoskvKVK6+ZtCjK0OgAXFf/5JF9W3aDo9ZtStaKoiTIlY4T7QtFJP9p
vU16gc5n53M98mcu3BmfdapAq/uKnoG/uDbaVZdT4HyKeTlDVXwB4ufo9cQb+/m3
30d92bCy5GbqH59/fglwkzqmsmLwXrRZzEXLg5i0JwCl1I+H8RvULMH45pZrvMLs
PKKX4is+l11gkgLsXRWbHJNdN+9lI2jesaklpwW0eqV8npkAm5L75PILpE+9AqyA
/3MwWZy0QBBf+LriZYKBI0Z6x2iSl7NCrXoo6UmQ/jk5dEc3vwFgAcRnw9psGUup
jMiCmC4DjPxB2u8PflvuH3+Wdel8JgBa1WNYOFqQkv8vwMl9FquYYkb/kMkBfnwN
LpukmxnwecprR1Zx9CeTC4fnbjYEuuMD2ds6zcAlQNHxzzY5GTY+QLb/nLof4jrm
bfB1E9NWvz8sO4oJF25sTinTjwh14OYortxGKenZzbknG+KsxF3L0uEom3RxK/bD
WUddsKDANuPk8MQW4U4YVLjfpzT12wUyY7sfvTFrgLB/qBndTBbnOUSeseR7qAz1
IZX3T44GSP2OGmNsixIT76RRJwkNASNYHHpa2s1eEenCytDqFsrSGjzULaMmrSN2
WClmWia0hA6V2hRxHXlZ2yaTVoFOLbgXECMPgYIagHiyHe+orWhoGtOYochPB6o/
Uu7di6D7I8T/qywSnE2pk9M7afTaKLqxhXSe88/MSD+A18xxT891664v/IgvMtkm
pm4Z5B+QdRF+aR4s6hgJY+Mxs3ugiXZQUNEaU1xH0B1WYwJb2//qed+1xMHUX/t6
TgiSNX/Dm2VwcGSSk9AdTqTL1j4pVNIceZwBz0WhBai5WIWsnE/PAO+Dl4MhPQHs
/0S3+3NkMVSu7UnRg/ZuLFnbf0TAJ79gqRDseI1M9UyGM8v3U76dMgMCOIzWhIN2
tFQwT7qZtVX9T9iP8l2XlETd6dgnm2eud2O4cQ//eVVdGHd0QZ3cjXhkZuu1GfOH
B3VQrBMKDW34a9FPk8NUXkn+49zW5UD6V/bmKhFTW2gQEl9WOl5k4qVbFmF00l/5
JknJtMbI361HlEq8d42YOj5YCMqgIYyI/5oFuGq64VNhaKPQ5hSXhMkA9pmJcEEr
+BZaMi+Xxmk5FY7GYPs8ABgQfUKaH1SrIjalhLUlNwtypT7r1cMLsJrYcuz5o4GJ
/uPhxXQ1GIznalk+F4kLtlw4/VNOI2bq8Ll41eLSO3RxnI+zclP79JcJDpEeVy8X
6jll2YGZXEJtGthMWBO9EJ3RK5KmXU3wy/bsx3wORCCLknUSoUW2tJ8dg7v0fFe/
5DFwXKiDgmEd8IEDM6UdXjNIZoDtnz2aJmqEpAPFdUO3anBN3fmJz1mYrsAoGTwJ
45hqaDqa+et/B+7wkO0xYTTWybpu3yraaXjJ3PTRa+xJMcPO+WwrOiz1avAWJykU
TkxNufJ3/PHwxFn68lOPWQTxibWJMyEVrXqG7yvdBw/JYidyMT1mzZUHP/jq5Bjk
9RWHK6QEUa0kYx6StXNtHvOPZtYYgVMzH+s+Vu4MxdX9l5MUlpTO1c/KhOsPZYFj
EWhgkXELOMxIuZzeIK35b6S6XLIrTPRBKTnDWMvKg3ifnyesjTyze4FN6qCBOPQ5
yBorHgwS0zfkBs3blf7V2mhlhVfeZ3X/nprcQT2iiiIOVtDE1RWExfOJbkgdnpsC
7FpgavUrXAxB9G2JIUXBWdqTMwF8d/jTc27o9ghG7gNGfkbpIvb+42A4fPjByajr
lOzi7hFMFOLqR1LbqzKuvPITkQ7lMxusPorLT8g+DW9zFhCYpEnNx3EoyZCRklCh
lYhDkU+rXAD6jTpttKQ6lnDrdWz5/YiSfnmU+h3QYKpy0sew3Jyir2TSNZPR2Zjo
VrZYo7ZZXoYl0DTwWAR346QwkAcw7ZDIFxQLr4N6XhGp20C2k1UFynfDwLZSUp/i
g15DVNOmLep+lVEJfI3igos+cneJ9FVyXk4rG2Yh792kQ6mbfQOmpoj3NB7jcZ8u
fzK2f9D6ZecBeANG7sjw+FhrOuD4pTtuxA2EfkKekQpF1+2UxNJQ9T5eylNnEM9k
2V0JxfY7IJbgwRcOfk/w2VDQJNUqZY8P7TOOEN1xpBuxTiiB8BkUhzAKS0lgd1y1
NdYiVjT7inhqoC+2bENVghXBS932GrIV2Fssp4k/v7jejbPu1mZevE0fzj6HBe/e
MFSwyQq1/0AqcXk5ATvS38dy2IhyA18mrpSba0n2eUcrYZySrrJHQVAZ2yF4xBuu
0bL8oPps3I7pjMuwByqFeS7f4AwihwImrzNVCMCawdh8fBJRCsp3jkeqBhUwGW2C
ND7yevUdYC9HQlLVt/UpDh9X6I6mj0x57roYeOXdQaj+GiNnc39AhZOoVwHyP7YL
mTRg037UdLYwh79zDQlmN0RYYAwlbY96A3Q8gw2FT+QLm0Y87GgJDuiCzF3AUPs6
xPu5BvEzSlxTl6Ey2tcBQ72tly3/zzrt+s2Caqgw7BdfjPziAvJJLIUkzKqjaMMX
8QAZW8y58YIL7oCMqUc4kQUc7xya6Sl3ydSLkmePmDwOjS5N9Cw22F+UZGAhBy3H
PNF82K7BlBfG7yVjEOCBxjisrFguKr3dkt/q6HNcbDoSfj+rN/GoFqTb3DJ6fVeZ
8CgcemnEqjyCH/QYG9MP2clN9lU7cokSdkne5FVSUJpWfjQx1WtzjhwHcWkQGpKC
99VcBRPeauUU0yx3uOX4PDf9TMYiDrH3nOGHFOiegy3wrx1162LPGVdfoC8Mn/f0
a/3tT40dCy8+zQFPLbdS7BuDjRQZ5474sj5UDnQ9HUFQ8U9zaB7+V8H0cJh2J3ak
wYlPGcgY8IKpCzvkqE3+ARcMDXYSBxwDkbD8eDaR9F4plCaD0fLCpMPtJuBiaBA3
/WFTzOaxlqfY7T6hfKLcVeon3TAikwstwO8vtQNWrVEXnP0k/GiwGRN4FFRVEjX7
H4fu8v7+0qP2Xs6V1xtcgkDPuxgnsPQFtG4U6GWaBs0OACMFNuzK9+GXk9cosRj3
Y7siMk2HlzUiS3zNVyECaAQBGmitAeK7n/RdvxNST554G4jZVVNohwjeVk5TrHh+
uMZfRGaVJe8bgWWqOqX685Jjjlr9/3+6qG+KIBgsPlukxy/JCcIlaV4ABj5Ab7f3
X/0BY34xT/k8zhCXKUHoVHBCkbETB9BWWAhKpVLVcwSZAnYZ98PqI7cA1eNn4Jyu
2Oikyu7iNkrZbce/uIBwKeCtJsCnFBeVY1NNmGMvY6yPKBLMuyI4JC61qozQ48Lp
z7xrFel5LvOjJsQOEvLSnVN14hAajT7NrKP04ZDBb0eXyL+7MLdLCws2YUGTucNv
TBoS3oArKNvY4oxWEbTBylng4prcT0WQwns0RURjJKH7wYq3kwiZLIOq28PQ/J38
lpFphoeXZug6t1XNfLl2hVCQqbFIZ+aYq1uejgUDbYv8HDFMajXzxWKSY6b98JEo
iXJ3c1WjnE5OOh9DahHDSg/SwuakEEuz+F3NNJLFS/HiV+7UcmrlAP8mM6Cujc/N
VpxGDbPRIJ5NCcYpzZId0NobMrePcBmZNUS6hCO/qUo1gy9LjoUDxuWw3cDKzmNC
wu8C60qiTTClL7o0NrgU4j6Ftc/1oy3XuHn6iseKf8VMZe1rtxvMum3cNMEsAqMc
Sy+hz7na8eKsesPZKC6PKUApIbiF50UXi6mQ+mMRNZrzUv/lZFarCAmjIp1gCAwl
9klvkkGADQq1CIKctvKRCm+PDpFiZrBo5kBcHVOAjdwk49+sFybIJEVjDGZakste
Z+WPsdyLv53U70Fl0+pT5HH0z0hFtdSsGzMJNryXcgQVKd5WIG0ZuZ/4H2mOa314
E5GKqKs8Q371r/ecxMUMDC5t9pplW4lvJQnPTPoj4ois7jKmnMV1lkYPeJikJ5lk
tRT01qbc6LyAOW1OqdTMzHo2QO+cgDkjEDuDQ9pZVDXTFC8h1To6SzHRWvBvqWvk
Z1UjcWxDRdBXEg6f68U7xvUMFukQc384f2DUccU/m9uIwRlZ0mc3QHj1jUSW7Im6
QtDK7kdpsB/QsOa0dbTrrLVUiIwZCgfZLGXVJEnya31U7CDTQ0WHyRAgmjCGwH9y
OlAxF6ICHRoui9GFG4Ina0iVASu0LaZea8ohZS111PYb2nZZCtSX51yQk46d/ABr
G7fmU1wmjO6d52tNVdZOZ141IatLaGuM7TPjHqjz/ILaeZOfonML5rxY0skjqYF7
vkw9FRZdY1CP8z095SWW/kizGuNTZyOvhHwCvr+SmQnMdjpH2Csljg2um1hX4RcJ
WLPk23+M3rFmxilys6m++x8SBS1d9txgQE+KGuK10mzaef/ilUHNur/BPt2c1gk5
xOVZquW3x2O9hzb5CF4mU6r0Ue95SrDvDyg0gKPcnLDf5p/l1iJZzBpAKl5NMTKU
7q5ypt3vsmGutyIcH0+EB263oZYj9V0WhsgbYVVLfP2Pk7tHo/gYSuOXSYoHWSdb
HmyKaNUUOxNw1OjOG6Lc2EN6oyB4XdUjN+/+TwWbJ47tq/ogbs83Zs/h4Z5qlSSP
mtdVYwgKZgXIWUClHApuFkjSuGnkMVeYP+ENjIPY9d5SEllu2F78wFA1Xrl9fUex
irvfzEk2bVC0r1ifoFu4MBhsVnt08O/CN2gfbaHBqKYlkELm3PWupMuNR4Akolza
9x4O6c0mSzetEY+TLFPtq9E8ayWa33FK1BRzEBruni0ryqsRd4d+QlEzqNpHFJ+J
2Lqz/gKYSsM6WOHMbP45k6OM9c2cqKsfSUruK21cC6NTHBsMbWob4BMB8x+6yJsK
x6w9fQtq2LT2ubAtoLVzjxny/JIMf57QqsIoCDVtiCdvsHjRouWEuv8r9VdofPX8
pc58986pqOLBdy0lZT1Ppizp7tEC8nFG0SKvg9WVY3UiWrh8lO3ikKO4Lk0XRZ0L
YXLCg4i0pH0sBqflbroTfR3kOebOmjzrlcCj0slSrAPjMWU2qVfyBhX4H/ZEn9QG
jkklsC5o5uVkx9ImA3QrNUzWgHMf0So+CG5+Ymgc7qFXvJ/eScyC2DxijrTauHnS
rD4/Yyt0r4X2e6vjYHbrgdY5NDqAr2hQDKgCycNIoJM3o378Cg0SI9DXImJQZFGB
78IY27TkKmDpDdgHZLoW1xN/8q3TPFOf5ZHKMcBabsLvZMvh2RjvkLQmv4WY9Aq2
9OtbJuCKbNMJHYRI6d8ZagDa62Heb8tACTnGxdsHjonGA6bubHaDG7VRsTfP8e9v
UZ+yf2OwV003BQ9rfyj+zE7kwGDuExqXwdW9I4n+/TyCRdGO4iraWmQpWVlWxF/a
zzmbW8SOqd3A105uPmdXucryLZ1gXLG5+02oy1ksQ1wCV1Rt3GQJ0f4ExdL9XlvW
qXBe/rGZz3Gla123BSsS/p0ps7WS6W8dcObetI1v2KBP/zRkZ00nvmRQZn9MX0GG
wpWXT3CdePTb/PLtvRuok1iEGYf0/BnK+SI8fw9BqtSYq+0TBPdjHiK5FDSArVhe
6lWMR2/ltZU03c3iNsG6lIyIvUIchLCJ7x8fnu4/IWOWntsstk9uN7slsPC3IPYf
bxDyJufT321WhT1n70dDqIaeIFn73PGlZpthf3h2K6dBNpuq1CLI0RAsTj3SXkU9
NXOiFasktYukaW3X+sypL7HhO0RUGspk8oLbqJ8yST6goKUKqGcR/hp0NQ4g8f27
Q3nt49kCalb9rcfKmBFbrNvKmjVyBFxOleqCk0zd0jZGThzaA4v24FQ3jTsRwShH
f+ZTgCagQYLGR6xZJyt/1u34JTW/sC/imDfxDu2NjoUv4D8EKcHDGDqkv8182EFJ
IVJ3C0G0dr6/M7aQPl1UDuNNyXs5ZC6SEj3iIkjwjZnIGRoTBqJ/MeYkxx0M6dsU
flGNKHTkuQT+eAUYfnpBDAyvqPsRED2/3ZS7w79ZcGbBH/OzfI2/6xu8nzHBSUgo
hlCdb5iWoWXXSvGz/cM9eIY2I/WvoKzpFiCBJirU5pshhL+RPYdEdGJBGjwjhzEQ
gqg5VQJ3wdeCnRth5vyaWj5YCW8hVfY0d1T14l5oy+VuIXvE7MfLrkuZWSiql+yN
EyuGcnxC3XkTLpZXyKseVV2dTRUe+ZC6N2D5nMRVAfNPf0YK3kUwcOmLDU8XDC8R
EIr5EoeuMVibi1wi5Fl/cMszqCDy9fgTe7hwTW4AB5Yd7uGZ8JHCdw/5IpGV4nc8
PrXQaQY43tjsRTCmssCRjn7gA8NOr0KnGpWOf1q1exsMnYilQYFG0wpjIeabK2An
V9bq0bRXNOgB+01ybqWRQr/zeT/QWzffRxp/hPClSqqk53cRQsNok6lJfIPBZYVD
PxCCSGUko4sSATnybncsLd5mATooFn11qmLdsHeBV6mOOWSLMTji/isEHmfbe3qB
/3IecfvmLBS40NffdGK/KmFdLR3xjVXyaEqmaMutsjGosXWqvPmSHp7ASq9wVPxr
uAk3ZaFhS6WFVEyes0l6iprh8knhPSvFhBLtSMtrnbu4JTzTyn9vCjGp6ms6eto1
C0bRDQglOiIg7KyeZnjmjswMeunwxYhFJZpwGnlQawBusAKbW38R7sDLkljw/xfT
FIuC56O3GL/y3xJ2V9AG+hAXHbWwU3il/DpHyebNeOgMlv19t9VcUBg9PYIZ5xOG
A06+zKMFsac7LA+nYN6D3/C6olg4uVBG/unwOMpiJUmwYGFH2z/55jBdR5wL1BoM
E8QzVma0nMd4HiZ2OnSqXR7U+2OgdK9hFKnIZDgx3a0ScFXeq4bO1l4fz2f/3c0b
8LJ6P5MyLRUzLhamEb631COi8jyIq/WuBFOvcrqeOEDyvRMzufUTqA9wCYlrXU4u
LqDd208bogu09ZFhFIio9AGHQRzQT7+AqiuMbPbPhJRzk5GtCqQ0ZCqxbr0iqnTf
Ec0mAnCz1gzTQuAT9+gdGMNW/ObW0ChRY8v3GuqePRKEW6nLArjFu/90fH3/Ydn/
7HxjkqEzNHB42/7llrmgIFYKm1RspaTOI1PMMJIjLF0tojuCEJj1q1c6fbJKbqbi
D0gEq4CZxC5CjfgISuH8lGWXaJygW3bvqXFXx7genxMn/TH8j/OxhL9jwDSSH/Lf
a8mziw9tAzQewebnD4EaaFtCuEdHAaiWzUw4iS5xVB7RIQMopG6FbTHTXUkFWTwR
B+Cb9H7VguUa4AcAWWUss5olVNUkJwFyENfiqi1yOVZdeN9iOSvhwIEgPRzADs4F
4h4AWiomfzlvAD6rbMfUNL9c8gb7ssrK+0fP16mDItsSpnJ2uzzJyHGcsOQfvBRu
mHvkA8GxAb3AIByxEPPdaJHkKDjk0B9Vc/3I31GBwGintm0OE5yUbKjAPgsrEfAB
XDvWB/2yC4qVJV+dTo0Y0kqkMoh045vLBSPYtlF3CTq0CBBOBW+96oOX1QxlTnjN
uq874LE5uPbJqzDPiw+cPieIa8cTqAoUAJNYy3O4TF/iFauXDymm2gQeVhFn8o3j
y8k9aIsYlVXW5lpJMmrnW/yEZ1pBzW0CRgsIYFmsUj7LfNatR/DqVFkFoJaIVoir
T2apXmqHpse9CjVoAwLsWufOvPxa10U1hXhNgMSdh/65kJnPU7oEa7ILEhVJiLdm
8EmP2c/3TIbM8WJkvjFiV3nR5yajKteCzRGr4CFAKW28unf6UtHD28XolZFYAJ9E
5xYwr8/I0WnJ7a6h10McAcTF+3N7X4nY0faHVXPZHaUCw0Cd3NZBcnWVtpVPvNhQ
YA7AGXudfngyp2SxBTuVIhmbBhfbtj4G7bLtzR1e++F8pqdQqNKmoHtp3XUb6TBu
CQBktoOYBeIhrzvgzJr3CirR0MqH/eeaOih40unftsBXBa9lgJbGkTjzkJmMeNM6
l4pni/K1e6ieu/zZSO/Qj1vRFJ3/tMsGQvl9ktPW8vhgMAdMEcC9wLpKIDuf9nJl
RnlaGIOAFrKeG9KoKCuPxW5CVqxyyc/YUEIvhRM1gYNR6yCKG4tFoN+U6Y5ZSTVu
hBjRo51U5ypKH9qjiVNq3hMxNzYrzHfWSmZcn4ZP2gFQ3mDZLD3ZaGzGykXbsM7g
rivts8KH/l9W6PnHTo/OOvhMfpm4VK+Zf3Xci+X8So7t0GnOh5zMMcQCqPvFXbpM
20UywAA0/VE6HdxNITQntGFJAPQRgHiF5k99Z9//w8oshSRTq1jXkTeZYTcJ7cEs
SQzHK/5oVMDO8vHY12IqG90r6oCay7znoDiUuwPYFr76WWNJPKDPIbzScJcqLlXe
CBO+8uSLucRrdKARgPvnJdnxuzVfZMtpePHAnzqhrwPv+FRhSXMQKdgsGFzvpF6T
crnOlHMduBkqjUS3qfWdnoSjZ4nPTj9Rp3VQD+Zc2WSCNvS3xEiFjsXhtNyIi/E/
nO8/vyl62dHwNEZ4M45tNisnD4X+waMOplB6cF3+V2Q0005BMwZJ0G4j3pPIH5nU
hkQFwhzJCL4o0Mxqkf8jXQt8lzvvfXeSpoKmyC/OMnhFNDV4d0rPhtedO76vsV3K
cojo5p1QIBhu7z82w3Wk/MfgU7CH8KWHo9mr0D8yMyu1ak/S5QyIXiNpsMWTOhla
M02YyhIe6GGFjey9XTM3VXZrE9U/mAOA+lMQHYXwvwpLF4d1AJ0GZDCgyJ8Ma2QV
Lv3rZtYVcoG8bhtS+0gavRTZ+67vOd+OUbAX4+3H36aaXsCVkAAdI7CgpmUs+zZa
9v3yJEaoJc3ZFxd4VnYXQeVKbDo9ox/Fk1YRxLfAk00wpFFdxE7jMEsMuJmedC0Y
NXEl9btyIXKLSb40xv7mVoeA26Eoep/D6+muGZx1FNGQfJyaNwKR2PHRNjNLliqR
vXAKpi23aCnxqa5lXX18XZYCU7ZkbUbR7VHlGc/YAP37dTgscZagmkPDJE3Pubaf
lkx3QLoeAWiyIzC+i+EGtPS0c8Brk8YhfDaSdwOJxESesTgdWDu2omylYyQux0/H
N+t7EzrWwhkaR1rvHFwq12ykvAxyGZg3rJJFzrnP+TQfL5imz721pqp32n82secX
HCL+QdXOFUKAqKSNv6rnxy5t33qIZpOHiHujrQBuaNTQhwWBprstmkOIF2n6T67j
hUCVHjKvHBKFWWcjFZ/RUa3sTyfUy1TS5Kx/OysGUZJHLVo/tw1rd//w+SS94mFl
oYTrBoa81Ry+SDPNowj+uXFDCdRvAPYAxfPGCNaHypKmWU/VOfT9wuIeHg8RXehP
5/Ky7IEg4YgXOg18WPEPSmuKxbGDzvuHclcis6egmIYSNUmJsjQKKJBgYU03Lxrf
kj2syTgvVYxZ1FRKPC4bfcebxhHKedZcknJllZXv50Ge/cdUQd07dBmjnVejvh88
f6+uVw+rDuWJSZ4SWbdcirlFjtQUNYWw06jNCTd8gfnL3MUXohrMh5EeLkKG9DB0
2KneOA+VWgRVqLxyHtVJI06DVbLnpu9y33LUiSYSBXTQ523rCBfoKo0gYcrMc+Kz
O/XuKW/EKl6YcipAi3mygTJsjObVE//wEImVZuwx2G+HOkffo1Q4uZgojhU9q4O0
uNcHLbbS93ip6T88uk+MN2McMPu61VFt7/AgtLpuJUJG0+o8uQqnaKRXMpF6S5zb
q4D7ZdpQ51vmduiBo8FuWQpvcysXU9zpF44I9d/KF/rV1T5F9OIu1p4NNQ5dnM/i
9IHxmhYG8qaT+bcPtO0nMeSwAPQn0TcDt7dIB1hteUnWcvmemJUycRP0DUvLcjIO
10pgyzgYa77c6p6NqM/tCwfPNi96hcn3a4ySMAwHTdF0CHHN0++vBgErrcCLDqXq
issemgU1Oyzv0YXZChN3Ldh7toqc7+/Az9aTFbJwFxRIxZ5Ws1CZ5grHXH+kcm9P
BG05nk6zDavtKIKdBtC/ZNAMHh9VaMmDlJGSAGrxGPU8MbATNk7LqAT4qPpfh8aF
iFsyiAg67MTLABi7whP5B11uQWJ7esZ/BWlpkVzd2ul23cQXN5U7xYOvSJc69dJt
WyG/2k7ya0XkPK9wcO6aWooMLLgvVCWDzZyQATFGMdxSiljDb1lbPOh0Hz03bawz
pX9ciXoDmChb/CtFDcD0PnOMAneJyqoVER/hVn65GEIPQOPE8X1b7gZTAwjavvix
jTbDG08EpV4DFDrO2qMkFApQzxiflPyOa+SFgiR1RbLqI6+hs7A6eTF5ATx5oUID
v85UFpSom6yf5j+r2rhlP8SY5Z+Yba7C72BIw8QJ+wus5lklKgMb5IT6XKTPIAw9
wWSPF8x1hsJSgA0Tzt66c5EokvD8+lixBuI5td+LECtHdHPE/eUBT1RglFXePIXK
bQcTd75+nsntdKI/FbAH31dmy9uhobX03wmhvxfduujhXQ10fgg/MQ6wDYBecLb9
mC+IgZ64Y1hhsHFbfYu3anDAH8fqAiE15/noNrvoTx3U1txc1z9Z7miYjJ8vXC83
vIE8JbA+gY+wLROd0CssJsLJ6yRwl+UiqiXnJtwlbmMhTVVbq+aFGPDxAGb7wNLN
0DFaAsjlbWHdIx2n4r7D5xTCheBu/i2XtPREdtLNfwqwiyRowmv7jGLDjazl0idd
aYb/TyUi+UkInutJ4Gjy41VRZYpbphI7SZ1xkJvKrjMtasYSGMZk9UVSM1HEluVL
oa+5SmYF1eJ+Tpqbm+37rHoKs3dUHXAw3lF0cFZfWiJRs3laF6SlZCy+Tr5NBCkV
/scYveQ7HK11jei7x8Boov+sOv4Dc/zofkTEF/yESCzopFrpmsZ8nvinbnOQcjZ5
ye+uYq0DL0wtxLAhksDN+7CD+TmB2pBkQRDGb2R+Wtgz5eY+9vuTSb41EHk6W956
pReG/PfEUHbVOKdDUYfrH1EfFVk6+XRDhQK0yK5Y0TIpEZ8YRrTwuuOTh3qVazca
MxTZRkzPoRT69PvXLyPOs3MV5sTkrLDac7HtnfzOLSu7WBioORnfNoIFHAdSEGcx
rnU134BnlbjUYhPduxUQ6WALFZ+ZDpCeZlNoOidI+4NsMXtUtguyzjxCYfYoNkJh
4nT5DxVG0uMKtsB+kRV5vNE8QpuQN3IT39TbzZGiNt0kG1OPSZMa5uVO5o1JivZF
cSy5MPDHvFM/OQapu9SgkAtghi/Hv/WD0zgxmV/F6fS7oAUrX907Hn95jYpBm9rf
yCrVSVrr2AkiY8GcVw0iZQ1Db+9l8vEjODX2fmjVYoYpazpyn5IfS+ifwqrSdaNm
1k7mxFetuESfxWjpbdiuNbe4hyiXGi4KZo9YqpAom7v2C4aUaLvi6WUXW9simzS0
u0lCZtvOxYfwNBow+fCdRPa18tgTZn0DfT/HILKxnw87NI+U7g/wPAX4iPTaTE9j
nWsl5V9we9J67BokkpD/TfocKuMa6K3BhFmC7TpAb+DakAh8PBu/VlBOee/Nt+3C
dhjMvst5m4mIKRTfnIcHjymUvpX1Z6gJs1IF1jpoJiO7opk4nCezbw9E6Nc2VMr6
8LvO5rMFLbf9jbFntf0piuR+96KISrhgu9jwjT4jK+6IuX3mP8/3guCcUBQNU1Ku
fVPpdikgsBaEY1DYb+Tlgj5ssnWTSeQcuQEcNfZvODNchqF3Og84IZTx8M0W2NXa
r7ZtZEAWvZHBr4ylgN9K+iF2snAMygBlw9kkE/elg0mK9fY58yBsLgsyfpn+8rcL
ulU4pS7sqDvSmLSWGiKf31BfI6AilLjaDO/od1JOQ1c6U6xfOKT9L3kccxJltxqq
0yg6mYi1QkwjSF+DAx1+bSN0dNLcB0wejj0UaUTP4AME4L9Pyughk7YCfhdLCYQO
PCCGi7SYwhPSQAER0zMtg5FjH0+mQCaabsbtL8WGFgzqXeKVWHSwHtZd1nXW20nE
RjGixH6auIbGYfVqzCFou/2KafarpGU8n6iLrC06L6IGBey+uaBfxPYkVRTdVpSa
29ogH3RdAPLp7Z96uKSnAJ0Fdsimz+cntP+PdJ9rkitUW/8GiZWxvmecozOyViBd
GMAczuTG0m+ZGB2X5iOwcemoIvBmsrb+mgIMpJSqSGbHsqlkC1RZtrUdlv/AYAlT
Ww7dC7MbR9DAdjZa8Zx9xx7GUVRtNjn0bRknm7Tuw3giOhoEhdtJ/Xket2dT61Px
3ENdiUEnWIO6Hm1pLaslO8CZdUtC+OCl8TSgHHnwVQ+B18TzQCRO02ok8+yAZHms
4SBAUQlHQO7K7BgW3bc0f5o8o2/yQNQ3oLjbPCp1ytOrsodTy9ky59cByCXhN4FR
krsV84G9KL+RkJyFFcgFYh3TJf48G3h7ZhzJZ5Tx4V0ziHwHQF4kwz9iaWIRu3ij
ZXPlexb7UZEXLcqIGDVnbIw4KFfVNT+1sufZLqN3RT4n4o5OPPB41xKiOzMcfQey
JQiD0uhDc1Sp0+TdqXwmIgC5sSZ5EgB3AkWUyjk0vuVFVovHi8yf7/q8S9rSGVGo
Ddp3QZK1iQ7kKPsKRa/UPCRXRFXDZZFJ3as+SQy+b0RYE/fKKsAj+o1zxJOC7gcN
kkugPr0kyvoElpBtTNgkudUn3AJvXCoGqxJNKAY4BcHxSxR/faAj1YY6WQT0voFQ
bSmIgpcSnEWtZOKSRyQU6VFINabae4Vfg9X/7niqk3DHVqwPPy2A7Zj6dHjKrkwO
uOIHuCgZ4smv6aPl66RbsxzTncUtht1MeITqH7P5h48ICNbV1SzojXVhBtrU8kBN
nrrcTRh0M1D9M9Nk7OM3HA==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
nZJS9Xxqivm3AsnTdk7mP7/d8OJ8HPzX4ZhUFdaEaikjoETTqSSZ34E1AjN/YEzr
8yXiOFO2+CMVAZu+eXJRac24z4VtPLrFPy+hILmfus5OYsiODLShdmUj5Q7PobEl
BAvHbUvEzBe0sD10y/9KP37frWvc4qe2lQ8mrNsECvk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 30141     )
Rkvx7XOyNq/ZrWHC8drJuwqqOjqgLcvaZ9oonAupkEATCefANlaRuUUq/MjEvszX
5fIyU2mLYDbLEwhf8JQR0iscosGlw7RAGiYFSzVycHiZu8vrg9GADdnLfu6HD6Od
IH5M03wIVM31IvsMFR7wuQNwlPC+r5vS4Xo6/KYbfyDtsuRwS49MTXH+12fquRzV
mzf7OemnMhe3++sd5Ew7Q8Zi2Mf7fUplZ0A3Gug9zWroQ57re4tgQZ0gV17RVcrG
FMxqaj/ZTAB00mWaUFpH+TgA4PaWJ+L2DXtxLuV/CNw4y3j+OKy8cuRdKdY5j78S
ZtJo99+HILe9tkP6mb+UQIS4+NKG32QJ8eSclH8GKhtamZw1BeFDxTQZqucHst8Z
D0m3NRXC8oSQi8sl/2VAG9DKSi+2MLF+yQ1gXB+DGcyUO2+ilCAmKm19zggad4Tk
tAKXN9jzEG5cuuXPqN9f3l4xBcBMvKdpfJkhCd/LZApqwIi6o7jbSZz4h35I5U3P
jWR9dlTE8BVNVgH81fJ0eJHVYq3hw6Vt2g8GktnvJHCJDMOQ/Xx0C8xdhGz+wfvv
7EajiXC/8PqpmLrdgSvk7L1qUZ7qoK0E4OYMbFz8CVpG3o7N+zinEEK/5+2kgHF6
FOh88laigbVLrST6cz2eZMWwmPNRtGFVmaf6jBxDFn6B/zSArgaM+GQZmT31fLKm
2N+gYR3aU3DDWKrj+Vp5gE2DIb/TkIkZD/ingvccBKU=
`pragma protect end_protected

//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
bBj7RE8CA11oxJweBUB5/4KjhCAefeQebnA+7uUAMzo4kmQWIU6N8wmcR0sNw8TZ
MybsNHanripq6+QCht2yAcZGBFfOS4jSBkEWYdF2bexpKGbbWZgollFna4u1HdGY
S1lfZmCi94c9C6UY3QgSDZkvvM+/PuLbCGm9navRlyM=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 39659     )
1wJ2kd6yYpXF42UjKbEY048WtnIdBMbKqidhVQj/CpsYoV7eOTJWekfnxLg18IQq
QQYeipVHqjvHi5gqSC5b58jHL2D/R6qVEnvaFzC9uXNi5tgmV79Wcp84rOxujTw5
P7la5O0Ib3aYKpgCrzNIm/kdg14B4+eQp0FR0PlWMJz1pY8ZUH0/wc7OasEp8RX6
6AFQ3awqzGqHH7IxgL+4t83Aoh9FQ+i/cn0EeLbHdYR6iLKTDa+BeUF+Y/YI0KS3
Ibs6YceNSNehjvVu/gZUdHCDIe3bow/1fm8bI8yUKxxzLJWMKmlilVw/VdR/SRcx
ZvsLUNkAt7s5ddI0um8SugfEr1waQIOuW2DRtw4ZogfsA5RIDC7GP5+NP1hZdXfS
ezp7oLl0DIGyP8Iz+8XP7XjUa4rmyEwy1nwfQJWDjkpuUrVN7BIvht9JIhKi8aPW
qRoxzkHj/GklFceXE/gLa+4xaEbgVRb4lFzlGCfbHoMuTKmplm26uapFeSSvWVhW
ZHS7tE2E4OxXF4mgioTOUsAHnVLMzQV1fVPJ+tAL5ubDFpfBRizJqrrxdnMAJJj9
8TnBdW3U62hDnLDCK9FSzKOibzmOwy4yPrql8FWpsE3Ie4EV7jWMkCWQtYl3QeTk
uaFaRFfuhgRH0fes4/n6k3LqGDuNXXFOFlIZxXsl1YiCb0GkDjSxGaZpP6a5amPb
wNhWlkFHROvQQeNV66RHsw+IYUG3ZCQz1fSHT38bTHGUJCSEKKssA53+pNTE2zcT
yLCXLxwLXCV4dhTw0TlNLGtgwLj9c996yf+UxE6uZIDNg3HNjGto/hhJDE++EcFP
JNezOni/4CJR3zmz6aTm7vY2uukxJbpGYUkJMBdHxQeOS6mduAKYtZFEkxCUMmdP
IErbYFWS7D8wcBPvHPTjC0OvbSLr8w/w1xU4fJR3ML2OMfwKVANda9g8Vt9sTA4W
7IaakQEF6NmwZYO0Qr70LIhbNKC/v7TIKfy/jwd9jq/aAmFyM0CHes0heLdGk2V9
hU5H+AkdVg39yuszlUGqaEaMmrntnok+5/5xvfkjx6xygTDBMV2W558oqUbNRLyc
akA1A3Yf5dRYW53WPOfIDSY1RbpFah1cnYelP0bg1FdxBvwdW7Yf3/dAxWW2mZYV
drNqYhnmHBDrElld/xaiRjSftuJOzmYQ1YG+eNOa7NqS0DBQqPscAPeEJOQiHltm
hJMfXoP8S0yNolVXbZa9D+xENaoV5AXXi3YlRwuSX+68nwsBW1QhyxscYSYlj2+5
hgVbzrewEsQ922780EACxjRW6RHc9i8BEK3zZv24zsYcd+D2PR3f+8lBk/iyApQ/
qaFtD/P6No3LXQsqDgqKoFtOncQ9Q5hqyuSQUuAEI5gMRyTupdSL91hm+4E7qjRY
BL/3MuwLsgN4zTMt4aix4VrXE8KSuhTZlgKKkXX9BkdmqgiHafro9qjMS/m3Ysis
k7DHkJh0LB0N3O0Ghicl/JAa96vOfrKorb+fyBxxJ0xkBhbaAmTvqPw8HQVOK1bh
mn0PV/USE9KF3iSVHYjw72wsSOsNgJvUPmqQtpU/WDoDD9WcrFvnXssA0NCTZbTm
hrzPsJFfZc17hqfm3ozx1zPDHvgTMGpMktIKgMKfdXxJCmEpOOG65aKFo5KNSYX1
dCYYnJ4OKGVb1XBaBmOPLlqvDM3Hk2n+ZRpK18VUJ6Sn2NbSykhBpLwbQM2C1rd1
Ab9VkdtqkfgVkCz5fMqQSwlSohLyGFv4Z8FlwZvYu2j0Pvt4YTX+NoeVIScixn4B
V2deXp37VVoQtMTjaASlvX9jC7oV81mC9FE02Utein3L4miUbEJ2IgqVm6AVH5Xl
EL85YupnzoW+cSsf8QAbZ9Z/TNSGoX05hJJP7rLVUlifALQn2ICiChNd2sRS63t+
oe9COdbH+0wOCAWh/LfoNmX8DpplvyzVja/xKaxJfwptHiBSHaUZfnreC3WNmkux
BrvN9ZbObU3FwBn0P8XG7+9+h9HqvYIg6ITKz28AIA55meLOQm8t2nPEdtmMlIH9
i+i9JOVF8GuEe4hhzt9ldxpsRFkURSy/xhYwnNtjP35s+9gro3E0CNsaI6D5IRtQ
42AIWCufsgAuXrFk8kurnjjSbc/43ssmr8MX1gNjQytq6CidF3hRg7xVwaKFo0k0
DsB3ufX7FY2v4T8zxm2+z9CeFEPJADFJQXbn9/1kIjXPfSRzdvIHsZT598NT7VMJ
mTgcL1NBsARYipAPQEf0r8c/gprJKeGE12oJj5wrX6TGMcTdURJD3ywx+eCiQOxp
meeNcLV2jqzxTuFMCR0chfEKNUT7+kaoqn2r5sdSF7SVay83MdNcyFrHOzIfmEzL
6X3FAbuiE3oefqr1OjkTAFyfUpw9c9b2C40uYu5hEarktMHGH7+HIlLnWfhneqBU
aerUrO99J0K3MN0TyFavbYZFJeZFfvCbOmIJMmSOE2wa4XI/zfBE2TztZqj9MuWI
gZiL6zxGxhfGQ/vs0ph8IKuR0XrrAxAQEv6ixsZjNo3BGciuGZarPXwqsX1SuJdV
ORkaOMmvq8fqx5133QXPz3iUlcfnCNMj+8a1he4ZGV8Hn2u0fZJZ1nfLOipc10Un
0XggSunIw3Z2ngTyUrazz3ZOD4JvgImX5pNFjbwiTZbL7H8T+I307fOqv9Ou1KyL
uDYcHzIxwdPImEx7VtfSs/5uq/MR4aA+knj6WIYNfKlbZX9xDC4/Sn2hCDwZWP63
V20+t7lxYJgYAvKnwivgEZY+XKzCA7HAmwkqCl2esc/lKTEDlL6hCQDY9kaZQLTc
2bEP1Yp4htKogsMhkFKwTvTTSsDRXGphzUaQrGcSs0UREedmLTrNKnt9EM3B8jkE
mVNZHRtoc6RkzHJdR9WDQ08k8tDThPHV3wHlMETC/9X5GYn+IecvIr6RrHxfePq8
gUVJIhCjHTlIu/LBBIL12kEGs13pec5ZLRc4JgmSMVtnwqtYB90Zyi0XbAYhKxTo
5G9LQFmJ0SgiShuEydgZofdFn+0Q5OroMlad8l1sE1NTy2nTm7p6YZ2Wz7McFWwF
QA8mYRuGZc+OskcI17GApdtSuipFjd/n6+AHvD76g60mjEYWR9kB+mCDdNxifuyO
i/WM0JE22cPrlPiscarhJuSoEAt507E3AR+mzPH/LyCdPgYDdpgPwW560aXMRb0F
zs0cMzOJH/FieInWSHUNGPbRelLUJgOGjXQ9ZIcyWOovy+u7tBKeRjvMdrD5IbWW
XfdTlq4Mj7E+VUfBLxNVkD3/t1xQWv9G/v0yqZLUVTnG7Gb4R7vG2nUE+ahtkqNn
SYYrNDpI37c+MPsrrj8QXEX2a6b312X89WXWanGrvLSSmCujRcu2YOJcxFXs/hIX
gY4EkxO4KYfNWRAIqZGWhExhMEL96ckYkMABUPDOnWHdnkdgz1/9e3eJRWoe8v3t
yiA3VJBTiSh8byovTk1v78UR2RR04eR9aAMTCh/futyu4FBu9FlOzU6NoYrwgAuu
DXL6Yk9X+uIVxO0oojWYdJllp9YA7jT+hSIazT7bAHqjhVs6ktr79YKTa9hpao8x
8Vex57rC8XdF9tG/GeIdb/3NvEbjgT0sQmNXTC8jHNM7Mx79pYI4ZhwE3PqmAbgX
KAjR703LnmWeKk8HHEl/9wceOPbCbaMdzn7TM0biyx1oQWclA+1NC/1tkJExGeG1
EdNIBsuLMWtm9nhBpmPKoDGo/il2L3ghJCBhwg4zQGUwp5DE0y7P8GISVEMf1SMs
mS9r3z/tlGVjYk+nTrnG+91UyFAkryIjTOQegB/il6q+YqNnB8owfc4ZQPQEF2U7
eUs2GFbgMZ7P2r46G8HUrganJCP71vTOB/LfBhHyJ4AKSFJAVGNpMnXPxZANaHYJ
xfDHGKvMK9CwOr3iQCKYTcC+GUPvh2nJTzpluKTdfcukn/8v/uvFB/yxuMW/Xapf
XTwFGeEha7t6pI6PYTxe0bOomAWMNnjZr9aKT6UWug7b5X1wSLhEECgK7wSkAUF9
8NzuLnjWCSS2pqoAHBF0QQC4U3EgAU7Vrp8A0Nb95PzFgr07D72PgRxJW502k9L7
leWAwQf8x/8L3WExP0Nj9SKu9kYMa3zRs4N/sm/cKQzWMcnWYVPqB5HmgmqHbBqX
CZ3jRCImoQrVBokrAzpmyLkPY6kd66oZvu8iaqb8/G9RIdqZYPS0838n3d8PJOwC
c6DfBDS8JrGzoPVJN2p6gsvGeR5F+AKUppHcbFIWENJGM+AxaL8ygOzbhltoQnfV
/3BChswo3nrjmD4wxFXkVzFYs5yOH/tgxYRkXLWdy9qzOZ66XTv2LRmFFmGQEu3R
EnXq3zUlU6CQHO5BBQoJ9tTNnhd2zQTy9AYXddpRgdysKhstuMVIZSNtUtK+YEnm
rMGXbThSEY4zvTWh6c79VB2nqQo5q674ao5Gjp3iP0/L2Er8ORosdrI++tf1aMcq
/pQkBWbrapNDxEKxfVQ3VFa1HMSRIQMTU7sdzY98j3o5mgrYIp5POwitffLRawvT
xT3XtYJp/l3J6UDln9i7BVzRDS+MdedFfhwesW5RcDVqtz8BN/JWFHuzTSkdO8BB
zgdoI5mxUR1XlgmCOn8IR4hqVLY12lPAHCgiWpokvG9vMcO9fgSczvUYLFsyIX+V
/alvJpE20VhQuGzXKW5DTXiyU1qUC62njQv9LCYNWxkxi/MIOfBb70o+T40qVNI+
wTUJk9hUT/hL6uH6Mk1wXMlQWENrwoyto9k+H4B4UyUxledZOWwWJFz3PQyeb1Uj
F20wLI6aY0juAWP5nKYhA8Rb/nR3HxL6xE78Pn0XJiUd8YJK8yVDAqW1it3l2eER
OQBkw/CWpgmnxiRjabInJfu2MS8XBBVJPQmd6rmX06p1oNboB8ppKA/kKRUBAmcK
EpQL2dr71lWsTq2jvQutMC4T1WpS+oex4PwpfDNjFyjOlXIP5swCUErKAKg3WxOh
GQ7wbQ3balKbK4JvbUv0Xcr/kYSExQTnBgxg2rTJDGTm5sRlH0TSnquD7y6jca9W
iwoHkgQqKgjThutLcC/ZVJiEHwZsokQjt+uTFeQb9M2KStFaL5OwbcgbVeK6FB6P
Vzp49WW1JnVFHlwFO2djksFC8ZRkcCl8yJ3NlfLfiyzkAxOiPc+G8pbBN5Tyuny4
XpzrJhnI+VezOXWEzESzEjWzrHX/LWrjBOXv+Vdp8u2ZKb8TYl1utFPRi6LAdJlF
DhZyfxie8q7VnBGiDa5F7VaY544CXyiVo5zQZRO/0YlWuZXys2FHmlGr4RhbM0Iy
ed2jSKN70+/kth4Hc6q6MwhL4ZD0BL73OEOYnQsZgrc7XFuyyGMXdItWIk2TIzzv
DgHi3xPDhKwn0UhCsW7MbuiL5g2UlI0f1dMQ6ZwlDUsI2REzR8LaAgVJ/EdEFA+P
M7Kw7JOvX0JD9ZdYqpWwexHwds4yMBgdTyW/49PZ4QHkb+bKw5des64uU4R3d7QE
vmzt5xhbfxtERwJoOXe6WMgqk2jfzCH/c51cvW2cyFhByCCYc8DB6E06OtyflvuD
WGo1FzDVc3ZKgnhpBhOC2y80RUVjtGIVNoOzAx9+2C/E/+Z5vw8w9mDuK0dSP4l2
ldMhIlhJs6ZyRvrF7ErSzJFOnawuvtzVcjJv4JX+K+g9SyLfKTf4HGtTHA8yVMyA
KTCiU/wyBNleMcOOKerLouSYr8ze/kLcJ/fC/DYYRDnoFI/W+fGNPwY+sQbD4ShH
yuUeSet91S/fHluog8aBOX3znjRupcLmTlOcWQkxVISl5p8dBP9Zby/mqbtS21TR
ZqFfa3Hui/pQmiScG25ZlEvfzIC/F0SB3TBcsElXZ//fCLR5mKBTCVD7gdV9SGHN
/vute+Rq2ZC7EzP3KSM5BMHpXg6svUDaTpaz0sK2KKG0NtgUXfb9KOT+PFV0ZmwB
we6G6LcO5Z/ptzGiyilD1gnLO3DpPGJ+ztIZ7PIBYMOtkLwW9bWtN19Sz3kxwiXi
dNuDdUmlYWCAwRvDiwgpb1vcMoXkblhFA+A5k4PQyh4KW0j3YE2hzqruoHbmB052
YZaew3pPCNGgJta8JyUPeOUSWsE3IWo9BOVotAo2vCb8Q2s9NGGyyiwi9E5R7dyb
tzZ+wsEzFT3yBQ6GFalOF9D0uLcUITi9YFH/UI3+jkqbZprsRfEht4Mrf3MuztMY
LkYlg3cKrZEHT7gTqOBs0uo6Br1ZIfI1xu3ZG0VPbTrBMq7vp23Dykn2YteIjszo
rGO/+l169Ca3j9hF+ecIeybtWWDowjc3KgWe3x4ZxzE0KSUmlrdZ8maqvJdjH1fi
dMvSxkNoUTuS1bVPB1GM9JpFBgaOBCihLND7DR4csAb2Eoj90Vqmy0qOD935sO99
h85QJNFXq4MFNx61248Nrv4TMaAheW0/rh17OuhFMoHIWdwI/OyzMIAR5xPkoVLy
Cz4Jz1/QMC4e73xqYxf9zTogEosmAfVkBXxumMXJg4TvYmlgOZIjd9UE+nVFNcJb
x4jrWCrANP8/cpuKkSzI/zvxUKzB7wQ9Jbt7WokSirit28NkeyafhMfDUSlPcb4T
8zZkn7RBknMd1vP6NJjKrAGyQe89G4nUz87QDdlFLypd7C+NlpBHhmfvpHOPRO4w
KUOR8dZQB1tEUku3kSDeX0W0CPQyVlP45LzVgSmy15ZtMTWnIqrhed3/dhPx0WQq
UNVNl87vcdcm4C6p5h7iTVrIPwoQyA+EzOa6TOt1bJoXvJcHcRcMy2wWfHyPpR6W
B6+nk0VNU8GAeVflC3NWWJcpRCEwdcVfDd6twFpGdDXfLkmXMaKNhGT/lxV0QqoH
YZ39fMQMidGLP4Y7CvOfVKPPPwWVxDl5qwpjjXUUx7YlF9CDCoBmOGNmvtnPUSab
+bgeELf0QaRCehP+xPFSwWzUPEkI4c1yO865V0I8TDsF7bTQdwdZf9kShep0/Hxr
OQr7bHEJQUKg2Ao8EpAd8jhvHA9R0AWE/2k7uALSfC16jdXbIBp6cjqM1Ri3n6LH
rmnGlnXMkhOogvxHw2Cb3vbmvB+T+pTSKcuSihdEpqdNEYKnSdHGCz78LyTkqIBk
wmyI4vbVh+eP/lqpEHJ4x481ULTky1txAy+v/M7jaSQuhYuQ68I+W9MV0XrXMkL6
0YHq7W21kmsNs9YCTqWZgnJ66S8rdjcNLNf4kQQEsjzfcHkOzJVJkB1nQBybzXVN
1iyXxQRRUz8L60ttpIeJfaLeZsCDoVSBdDPvo/s8BPRc1nmpgkk8GAx8iU4T1tUo
f3L+dYYIoJQYCG1QnZFgSRICyfkr3dE+4Ge2goL/tCZzqEj6ZBMIpFDzoYUmoeYI
9qyFp+kUlEp+zIcc2r3EUgqNEoRNLFvaIB16OkuvwD8odGVNNnHtSv8yzjXlkKjN
V3Rr8+1JRQpHT1BZQa/4M7kcsKH6VBXeE4tiB4yGaE1i8c0P64LOP9Z5t+85qs4a
NjNdOJVPrHy6Mjhep+qfXni2+DCTs0YlxAo3DzSZck98B2E3IZ4uVgssDavyrw9L
ru+mOJlxvC2C/VG4pX7WUWoAwNp2mLVOZApi/W1dnzCYMqr6rOfDMbL5AMFglW4q
FmItixnlga71V+uUDGSVnzp4oZk69ilj9yuU1/ZnSxABGOQqe2jxwAgvRtDJFCdM
E7p81J6u6AmQHfHTrWpIQeu/NEvnn2Dkghr90XN9aEoD9+LuTk5cBeZqwWf6Ng4C
UIjnkJk1j1yyNByr159IZA7PT5bgPwQ+JNVbrGovoHikkDM52m+isb/lohS/PzDw
qvtSHjCsFLM3gwtBxoGavP1wXAXP+kvglGwnDnL9IwMxxkS4JRNcI/R2Bxl3sW27
RqC/YOosfxVFfpg23y5xU0PYmcL5W9J9uvKFQ7GkdZYGFXiB0HX+QXyo+NzVL84X
wuoMc48DBMR7RFqHPEcNTWl59+ATSudrp4Z584RnQIckXpIkbmVOW/qtTr3a9XL+
gNAbco5lJ2Et3FrnjY+1dFvecc8AKFxCDvs7L1aPwMJ6bKo0ZeYCjDW8G2uclX0Q
boI5LG5uFKodpUrp8RuTt/a2B5+28nipUB7YiB0dvT/2vjaZv2QojpH74XLAeRel
9AeVD3zoQnRRLiP8OIRxl7yT97DoNMtlStzVEOJABTjDK91h4KV0G2MQ3DrdOdKB
v2BbRE6QpM12Rqx4uP1YRJLRcetvydlKq60bMQter7ryYBGDWt6fH2wp1H/JsYrE
LC1BR5tjk68s3aPR+vzVcEdidnc/I0AqXArpNEwi8vGZXaRN2lfS7vQsO4NxIrfd
49s0OWd4zwl2OsVyO1rjOTQA00yOnWc8OCmc/VfnLPCVjpoTnGsjB5N/Mdc+pbeL
nEw9Wuz7bhHzz+AD+Fh/C3/C80DMwKSe+j/PPJtrCX90VuNX2JTBILVYKkyyZnZj
Vtg1gXXiNZKSWF67dV/jtsEFLzL2qO/KGNwYQqZhBetTuob9hPFMixxvlR6ZC3Bo
30bOg+ZXCZ1CLCvEgSW4dIXrfL/Sm6b4Lr0Z6sDi800lguW3y6vrdUgfjcxQEslh
qPWefU5GSg08cDFdPrtgJSJIHSkZq+cy/wAYkX+SokMLNELfjDbm2nUunBgGdOlR
GoAKTjMm2x517mnydKErU4A1D10aqGpeCu+cIliAaBR9g7RVj7z7fdR8lUXmMqjT
wgaJQRUkl04BeAZLyOos22dYM4/zAuLHvD1mSczE2GppHW1a3YefVKriMc42MzUV
CwQJcij3fQZRReMhG46hvJOIUTkbLSj9Hu8Hk+7WBC5sdJ5KppanGjBBpLbmx0PX
FBRCx9Od2uYkKk/fGca+usl44XYUjBoDR0wIngN4r2Nq9IsfDqF9pjihuiynBPnp
qTGdVFtOuKOnC01BgKed6b9GKgc1SvHdHzHLo++NKuEwWvOK7jxtl6231b2EOcsK
ebdgOxYJxH9Ev+2BCAyr3mGoQDKWVW5bEsghTYYLJjDNIzyVzHwIjdnac5lZXYuV
DjYxndeKemnCwXyyQBfus1zCAif3/kuHjl4q4z27q/PzsHbrv5m4BFxnFEH115Qz
lKXsXlaBpwrCWZeHUEsUz/Fgk+/JSVhYhltIf28GsJY7vyQqH2ifSstcY2QTXXPW
hZjmoBUTsnAu8x6oLUu/Z9sjh3IdwIiO4yQRyKDt3K8Wws39fO0WsOP6oIG3f5EH
af2lOMHq5fGJ8TcuVGM+G7Nn1ul3qQJtuKW71hVJ8GltI9p9nwqVUNkTV1HMMdWz
OfKOq6y9pB5zIu/gQWKFFvI/jQGVCAVYFB8bbfejeRqFBr5Uwfu2tEUNov4NmgGY
+hcytkMHyF2vfbkGCYeTOUhOfBAfhu8/oZbfItVhGYi2GxMVbKHQEjVSLpk+YgCH
j3d/qdM+C6Pp0OzJzqAY8dd0IiXTZXKT7eB/NQXOlsJW+h1F7VkeFTXkYUAYZAlC
xGN8QWfcKl6NwuYMLvq75/GXVlXAAe3Wezcht4isRUgA0arkpqbibO79r9l82WVo
RYhZmkdRBcJSDfWWYzC2jWqXv8qwIpS5E9Qxw4WmEWsvjJpnLV/MqySY4uZ8hv/1
c9OqO/7PCf1c4FYqa2z4F+VRUamlhNMTCeqq86gIczU2PTVIyp0ITlMsx7Gn8WXu
YGroftt5NC1/ZQLd75QiYjqieEhptxNlEJeprx+m+58sGNU8AKSxhZ51WtdZasOd
sUGWyA1n91wd0tGHuFTEWteJEYtrpKpyDLi4JVEduKa12up7JJlv4y3Y3OLtJloL
VuRtKfosghRvrsjtP1wr/k6e93Hyv8mUz43UHqlLDjV9cpATWzIolcrofiau3qRa
QDhUxe7crL93qJg1tKRJpcJ0H3L9H8XBlBVLA/KDKN4Ri3xNW+B0J/C4sHb+P0Vh
YdDBhSDC/kLGQ0RZTujrkn/mUBf8pWucwA0j3UdfCnNA6pIAeGFaabMujzDCMYPA
/NByjcjxsH4ag6ylMGgXAAcCiSkTHpZk0TQrsYppP1+f6882xELYB0/Lwukujado
jepu5NxtGFb63rDVhADj7tdhFyaU+BM4fHfe7EIJbhREmHoQr85t7TZZ93/fCr1o
IYorakodYTH5ekGmIs2M5X8PlxT/1PaJ3KP5GwxEjyAwIoFoFLIsQYy3wW1wR1qN
Q8BL20JIHLWbaLLFhrv5UetRpoWflQv8X6jaIwJ2ZCmoUnuwHJvW0t/vXYd84r5Z
/gqvaUklEOFfw5gjcBYo9zijfzho4vSJHQcMcH4/fG1TumKoF344DmhKawNIcA8G
jRzb7NlLSygP3sYonwDnCYFsNxU9yXVMT+/ihcpsBNw4f1TROTrLPsie20pyLaek
GqGUW1v+0M/Aio0B3+TTWFMVqx5NC4aSQURMNCkAKblEqg2dCVAc49E5wXAmELKG
mSjhsC/SvXnt0q0gw+JUGM4IhqfZ18Ph+CgZwGn9pJF4swiH8IpEdWbTA8yB9PgU
sUb9K1P49MezJaJqQS2yVEwLcgqrou0aNSLWCDuUhnaL9yU+U7VFEy45pwKiKAuf
aLBvhzoJsh9+Ci36NJYmKBeq//yC/f72+h1Wjt+r9jBjc+VQh5Bpx8rTd/2AhWe/
WkwWZv7QDyDmcfhDcFDtGjHNkSLmxgVC1dwDKbLeYlSs33OtiQ2FXkdAL6/sgS1x
SdD57Ju9qLUiJzd1x5gRsu893S/z9de/rYOgqPdqzYbW2ceipm3BEEYcvjMk7LrK
oBIA5du1KI4uDwvwlllrpC2ATx0N7d4/ecX0XyBQrDFbDrzJbO5S10uWIn/tUhgT
yDt3HLIiSd22I6rEGKnM2OfS+fv8Vy2htCQzfBB9nKBaAuvrNzrA9zSdUDd8Oqk4
yDIUHUAMiuD4pHhl2pI71vQtUy2t7oh9tHFnZQetyOaDuZZ2SmjckT6tXPe3Ezkn
562Xx2cqyQFhbgPA+7a1nXL2flwbpNYm4ut64UBJ5/Km5HQ5V2f+2gADZRzcUVdV
PLJlAsYLtfrzQPvGYX6A+9Lla0u6a8KGnbYcR21suHHFqJFpPN0MY8EP6NUbHb17
uRfDwPcgU7tIKsMQFnxOzXrB+CPcog7MbtcdLVhXfoFwJGfPRmhTrvjOJMXopZK/
sdKepcyPdIaEVdLCs+s0qJ1ZqUYkcT31CLM15AoCEK7inI3bUT8zOsW3nRLSLgtu
RbLwmNneC5WAzKxBR+BFcaKIJxFsK7Xv7HFgGkmENxGSYEH7S93IYtVydsxPsTQH
b67+YEV8fvzVU15R/v/wS8STO2R0Zaw8JtKCNuqARPZ+jV2MgTKTAWxNxNsqJdVI
l2rWOTK4W1h4gLBuUabKF7lvlcASdPDh33Pt1j86h7CTCR8H/dqTcxYZu152DJWr
8nX480zN/FzuJI3Y34n03wJg/9vLGEWOCvMhyaLUlnsuq8XQcBPwOAqLAelRVFfA
WD259VDttAuftPBkXoOBHVIkebb4ysJmxh7gX+qQv7Z5sXnsm/nFiSdPu8vSMFk4
Jq7tZ6LiodRfr2KVi2tnkVZfTWFdSv31W8O1eLd0qkm0fxW2aHPL/AtgWpQ/RNf2
6D6XU/dMUd35deqovNIdq8gU76HP9XglMQBOkTK2cHMB9fIx0YpEQ42yW8yjsC3H
fjrPV9h2ywFK+ndLUAqdMRw9l+bdcXSXmPW5ROvZHqLIIrNvfKcKmp83oH8lKQHJ
nZ2+ssnov0TFB21lCsUcvZhu4TaY3LMSFiX9A9v4opu3rvWgtFlOtCISYNnBvYkn
D+SvYQAk+JR+99do163t+V/WBrb1vC/DenBdd1oFftbLZg3ajfUIB80AFnyPjOFB
okRZa09VXu4XPgYOqEeUG71dKEyQ6J3c3M6VsWqhS6PXEm4+MS59M37o3IraDVgh
E7hCFKoswnAGZ31wguHtjitMJG2keRZcPLFMOKQx2n///DjbY3NIde+ce8tHo3eZ
i3oEbMy7iO85LyNmM1rlZjeeIATvQHVPRW2TZqA1z7L5SnXcTysnd2MxBcTxzHU4
wVN+YD1HL1Y7pRr7NImrUiep0eN9X/gHCsgWlftuVVwVkLy1HtH6etsJ9zphl26e
9d9G9lVRK0aOa5dJ90q/yWKox5OjOmw8DqCgGHmtQ+cY485unGiEhsoyOSzfEgCN
x6BPKUmmQ80SMd85kYW83v8mFUHRduj810UBFiDeUSZOWHkj6OL3RzEuNVvK1wYJ
inI+UQB3g6HGUlKif3G6y0vG4TeYPelUS+8RbjsfyhGpfoyKwbdct8m8CIUVT7JM
92HLl2r8tB0NW6REjqskIQOTtMMU2vB8+7n79vL7zxnmgQCgTmSt56flA3bBxAen
1JzaTl8PmKJYgba9ExoEofCk6n7ibZuNT7oRk7rIi9WVFw7HfpBn1JwCdKmUFZoa
p98+PAmvZJqmY544lICv1Qwt76noaG6hYXvjkXVbhXi99ItM1bGO303NoAmAqODQ
00hiQ6opvcRq+ojKjRX4aFP1HFFpE5CG7ECGN1A5JpD46NwcyRSrN/2LPYVbUu5o
xk9aET2ki3fYsg3MlWNMf461rJ5msEbGxIVKnTFaeiosqszalS+h5kYmdyaM48V0
2ZmrUPd+k3j6imhOPJJDlEBhCXIwM73RO85MR0fHuCF3/5NKttiZdQ5Xy+5p6RAI
T4S3jRTnj+xC61uEvvCaNg==
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
CRcXB79YKn+Gl9w3I3FWSW7KipdbzwjZdxfIKoyJqNqreLv+dQvj9ZjUriwuizpi
XqudLsdSU+Zr5cCpOx13MtsPqV+Q2AttUEb8K0k4g1rzyKsV58c8wzTGlMqZSPQ5
vOQ6nM+4bVupA8Zs1xEH0NX81jA0h2igS9kvbzBog/I=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 39778     )
tF5bW3TmjqFp3hrkOCb7SQPwGm5RYtqDdlpnyWiXgdy//L5879ULKvx/t6x3dG0x
4eeX3uvPuXNDNJh1hVPSwEMNSOd6B0OF75qeWknxOz5T9h/p8kpdfS+YhTd9FySe
5K3/aWs0WQ//ZTK7aYOhCTRBYT+TfU0MEezI0nRaohM=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
L6VBtgEn9oLB8HG1BhD5exs5PXajYlDEHQ+R1nMG7MaNg8CNBWPs3xUBX6bCDSJn
rWTvVJTjWXvEqyWoz2tJtjELSMW3V9LPK/c3iihFO3RXqLgswzIAsXi0hVVYkxcB
DzL849qKBbXeyxPBzZDPbYZN+5m4506cvLca2Ggc0Kk=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40083     )
ZPJ8uY69Dq3MjlVY/Esb6JdNswBVDuBfGD4tkNE7e9x0YHdq+sWCncYjPJp6Vcjh
Moz9r8E84d99gKEo0+SJUDQcyy/QjfEEeG7LmKPDY1L7RnJ9ezSVzu5JJXxUG7dB
WnHyIPq+Od/8gLuW+u2Y9kUmis2P/Pke555PPKYpCxRjHk9uqEO5WcqST9JB3TaB
7RUoGMJMMBNB7lT8Z8Lhb5S84Zc1fv27Xp60lKWoW/5op+Edvubeacb4jGSZpAeB
yj4afIeczsMJ7P4l01dyC8NEtBbmjuFFC7P5rR2V0dvFZ7EnEjxfnlTmqqi2CM7m
f6sLGCs1olkkvXZ9224y1xa8cBOuKp/+NwU7G9MOZs3Ji8LsUwsqJ///K5rlepUf
ZhqubD77soczv6ERES9ViUDk01sVSMp2xlqSclrKL6I=
`pragma protect end_protected
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
l4VPYu5JwR7fi8nlQjeYYzHlDBraH/Fl+jcBxhBCEz72KWaVytwIlzq28CBEa8Fu
5z0C3tRPw/8bO6Uuuq85Q+3qkUxV/1tWOnQB9n+ZlDUcU1cazEz5ijglG8FExVQF
MygKhM6KZpuw5VvE2YQ7qUE+fdIr0qelOnJvtP6984c=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40201     )
Qkx+3H08t+/RYxE4q9Rzs3BQmuZy+BTh/mEOBNnACe6sHYzHN0a0oN+BN9x3WnIR
q1pEOQAOBajbeKMAtSfV4VW8fDk07IwgGnY0keyfxuAvNV/YTN5Y8G8/GK3KPMyZ
M5M/AGzggdZbeVOvc7FN9+nBdqURoCFqbWdsNgFb+PE=
`pragma protect end_protected
//vcs_lic_vip_protect
`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
OjAw1NJzt99Fhc6WBcxEcuMvIPQGbYLVQUrlwEfOHo6sUDEtsASHYepxprG7qRWl
kH810WQYdriUAd22VbnVAoPq5SlpRw/YdLWPvULY49FBEk8qE8XerABpX8Pvq/Xg
xa+PZ0ZCK9+B6Hiy7VvmKLrhgx+x3zGr8hh78Ann5O4=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40347     )
IZsKnzi0bJqvaBvO5iTw2HkQVK+4bQtSn5p8W+lzGTcN0dOHYZIdm569A1ZwPLoS
itqMsk4W4nIthi7abPAijkcfHt7yBeBGnunzNIqJ/jXrcAyMf6AFq1DYgHBBwW8e
qofPS3NuTYgzFHcOaOh1I/0baVXzTKVqmylA/gU/XP5j73Jz2xyY5Z/ATLsrWZbB
7nxa800sNqZvPD2ii5zMaw==
`pragma protect end_protected

// =============================================================================

`endif // GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV


`pragma protect begin_protected
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.5b"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64")
PJ0J93y2IxSEtxMLHlxWHn1PKxg4hnd27+ASqDvlprFjs1qoocaypu+u665nwzcr
pLuNg/on92N4rfoi7Y+g0aHpcnRv3HPhWYrG9FVatkejCO2oXTLvJ4xUUq+Nh45E
g2yzSp8XOcMvtNaN+3dzzOaSUisXa3kd43IQ/rw+cyY=
`pragma protect data_block encoding = ( enctype = "base64", bytes = 40430     )
+rbrm+1Z85Yjed+ZwgJhDYdRLIhZkaqFthkWcfFCWqxPAZjtn0wakaDZTc4pMBau
U/F59v+LMhNnHYw6Pd07ueUHgYaaw+iNhn51sqqK5Oz57iWyJiOSeQf/DlVEYypB
`pragma protect end_protected
