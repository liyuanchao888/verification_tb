
`ifndef GUARD_SVT_AXI_SLAVE_COMMON_SV
`define GUARD_SVT_AXI_SLAVE_COMMON_SV

typedef class svt_axi_base_slave_common;
typedef class svt_axi_slave;

/** @cond PRIVATE */
`ifndef SVT_AXI_DISABLE_DEBUG_PORTS
class svt_axi_slave_common extends
svt_axi_base_slave_common#(virtual `SVT_AXI_SLAVE_IF.svt_axi_slave_modport,
                       virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport,
                       virtual `SVT_AXI_SLAVE_IF.svt_axi_debug_modport);
`else
class svt_axi_slave_common extends
svt_axi_base_slave_common#(virtual `SVT_AXI_SLAVE_IF.svt_axi_slave_modport,
                       virtual `SVT_AXI_SLAVE_IF.svt_axi_monitor_modport
                       );
`endif

  local int qvn_xact_count = 0;
  local int ar_token_available[int];
  local int aw_token_available[int];
  local int  w_token_available[int];

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter, svt_axi_slave driver);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param driver Class container for the signal interface
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter, svt_axi_slave driver);
`else
  /**
   * CONSTRUCTOR: Create a new common class
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_axi_slave xactor);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Returns the consolidated response for the specified address and control attributes  */
  extern virtual task get_slave_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  // ---------------------------------------------------------------------------
  // EXCLUSIVE ACCESS RELATED METHODS 
  // ---------------------------------------------------------------------------
  
  /** It configures response for exclusive read transaction */
  extern virtual function void configure_exclusive_read_response(ref `SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, 
                                                                 input bit excl_read_error, bit is_overlapped_write=0);
  
  /** It configures response for exclusive write transaction */
  extern virtual function void configure_exclusive_write_response(`SVT_AXI_SLAVE_TRANSACTION_TYPE excl_resp_xact, input bit excl_write_error, string kind="");

  
  /** Waits for exclusive write transaction after exclusive read for each Transaction ID */
  extern virtual task wait_for_exclusive_write(`SVT_AXI_SLAVE_TRANSACTION_TYPE xact);

  `ifdef SVT_AXI_QVN_SLV_ENABLE
  /** initializes QVN signals */
  extern virtual task initialize_qvn_signals();

  extern virtual task process_qvn_reset();
  extern virtual task pre_allocated_token();
  extern virtual task reload_qvn_token_config  (string channel_str, logic [3:0] vnid);   
   
  extern virtual task process_qvn_token_handshake_signals();
  extern virtual task process_qvn_handshake_for_write_addr_token(logic 	     observed_vawvalidvnx,
								 logic 	     observed_vawreadyvnx,
								 logic [3:0] observed_vawqosvnx,
								 logic [3:0] vnid);

  extern virtual task process_qvn_handshake_for_write_data_token(logic 	     observed_vwvalidvnx,
								 logic 	     observed_vwreadyvnx,
								 logic [3:0] vnid);

  extern virtual task process_qvn_handshake_for_read_addr_token(logic 	    observed_varvalidvnx,
								logic 	    observed_varreadyvnx,
								logic [3:0] observed_varqosvnx,
								logic [3:0] vnid);

  extern virtual function bit check_token_availability(string channel_str, logic [3:0] vnid);

  /** Adds a qvn transaction to the internal queue */
  extern virtual task add_to_qvn_active(svt_axi_qvn_transaction qvn_xact,logic [3:0] vnid);
 
  `endif


endclass
/** @endcond */

`protected
KD@,8H0.7fS^89B;7ETZ-W5M&+6S&2V41XH^9Q,H\1fX/UbO]#L(2)e]<_AJAQ/V
5S6E3>=:)O<IdF8NG#2:#.1H2^B@\bTP6,/U(IEFcR?g;?F7?C#]Zf>,dTCBF>.1
OQSV_^L7g=+a^-NUM\Z>YGE?.\9acG<AW&5\:/6M(@0M(P.AE=e[ZWK\)HPa3<R9
Z5O@?aN8QJZ\HHQGQFaAgMC6^LKGc\g2)4/OP2T=<DJLNCC1+#DY5_@e0&#07H1a
J6<77QM4##,d_HGVF20O#=.3=_]G([>X/aQACH@._+:M:g3>WQX=dV-Hc^Y/5\SU
N<;-_/=\b<AX,^EO@f],__eT@Rg)TQ#=^>@[&P(@O@:<?Q7KTeYJd-LX0Z<#ag]O
XWDY(\O>KS@dNa4A\.C._b#U@L;.FP^TJLOD2BA9^A4+B(9E+0#KRC]5X@EL4>+.
[,FT/b#g??#7DBe(\8b,?Y3W1CD^9fQ0,GPA=L(YWCY<)8)RU-;f:73NG-5PET/?
#(;W>BB]AL;Bg37D^&VX(G>M_<8WVW)=a9G[GXb\661=aL-?\ATNE>@XT=4,8.F^
2Rg)#8P<?NL?<8c\ODRYNZ?S<IU#1O?^G<NKCEKTb:1gA2WVO3#6T8OR\W1JX8M-
(S>FcZfdTKB2e+](P5\_WS\.M/O+?dYFTW7K]AZ:MF0IM0+ZE1DCBP.:gQ<UP+7&
H7YN?Ic^?GGLG6080=U,0W_Od?&IZ>,U2S@&dI#2-cfV)@>D>Ec5J[@)J/aV]f\L
\,^E:5d^;FB]UV]Rg(IO2KYFC^3Z:Q&S(TSE,7]g2a;f:;_JH((_#<A#W+Z5-ZFP
>I,_,f,DQ<cc8]WT4cSBMP=\(gSX<@-OgKD&Mc[SLL5WEN[8faA]4^M&[&d2aTMd
,YCR83QP:W[K0=2CGQGZ#_.[MZcE=:+LD+S?Pb4\^#;YP:WU6\]>e2Q/bINIAP[D
6Q\(=&C707/+SD=PU<gM5C^+/JBJ^<[J,4Vf6Rc9fUI[2OO;),R0E0C5=C.?Y)7A
TWFb<&&@bM-)NPY;^32Xg&?5;4SE:<V^,]UQ[\@:f.G=/.^dR,&VCKTJQQX3FTAa
O0gbR@&Q.R\B_3F>.(=M:OP5SO;8E>2[R1SF8\Z+D75c7d.OGJJ(+(N7BBHSC_g&
).\G9cJJcKA=\FeK/:-Xc\OReK4Y0UUfV9AMV)H-\H&1TS=@c(f?Y)\B=&Y-4N]:
#TRGCM4FbATT7/#JY^QD+&#/J5-C^--[4L>TX[bE9>Xcb8aJ0A]TRX>__g^-XY+>
BZg7Bf>R8Kgd,BNL;.IQS?KLKD=B,J\?1G18?W(.?fJYW,g+S2E(d.,=BP#_#J?D
HIA-AegXd6\NQ4[=ZP<#5LeZF+I)a.TJ6U0a9T[Z9?d;BceENgU8XO+3,4LgY+40
+<^[9UHL:Seb@[>DN3<,2L?eFV-b_CFXf3A(2a\;+.8(:FE:FQ]R=^GP[TU.8_+_
54OZg.:OffD7CIU6\E:5WfOH^MMK5RP3gBeI/S0;Y-XE_)R3+M;L5?Qbc97BU&\P
5VR@>.<^28:,HI0Ke2Q+T[#S3XYYS6Y^(EE+=7=RUSF>;#c8C3[L@[ZSAKbOP1=W
\030X-Y&eN8IDTP_@HQ\)&bD#N-BZcOQ=6XC=]TM=U6C_e.;Nf)U^Qg0#C-cJ3@N
X8OU;f(ZX<g574<aAE0F7@GI0_+=b6)79Y_1TE;IEEG7-KMIWQ@<#T#259U50OHL
9,@C#+#47M1[?.IGf7eYTd)L5-Y(\]&\/OJHcT,ON&-\1g?8T3T\@fS:P@U?UU)E
\Q\^/&6D#VR<4.<.8D@aNLc;aSV1b<&)<2/X?VQ_&SH(0XG&@L0dOV2MaI3D;LXc
a8Cf]BBGU_^VJ9C082[DS;L;N4T&5@5E8U]^[JIJIGa5]8bbYW?OTNa3d_F:3a[)
d(:8,f9bQHK+Ye=Q]-R,9a-.3W4J+9=X2Y;1:EB2a4;_1>aQU#(_9G5I;D#_#NgK
X(UM,2YQKW:cQcRQVWag&/0]C,_DLJ-?B\ZcF#M]2\/_<Y6d_5>8aGP_L\+<\XT2
e&c3UZO#51EZ7YG.#Ze)0E8&FZ.<VCU^HZ-#(e9D@O#aa_5\QJ7)4Y+H8aPd^FW=
7-BYU4P@1?[)P-bSJ&4<06UdF2CJ#\CYM.CD3G,B7N2\_@CcP@T<X<]C7RKES[Ta
J]d?5^d5VaU_fY>&^MXH3MeGX)5PY6&<-(gG#H:>7_(+4DDC_GTV/;MASEdQ\g<=
]F5B/?JF)PJD9,LNOOG-VdX#_-FQ6/_JS71QVQU+N8LYUbOJb2.c9]Q7G8-4W@)4
#L\_GRMKLNVVF(_Y)GEC;0YL65#BVP5XK-T/&T#GI1?a8PWNI-a./aaH;1XN4)B]
?)C9)&^8-:S+,&T)<U&TR&)S,YNXS+[<6a?e4@XIY:)=cYLC5KU,W75TFdI.dd4d
VUYAOMYe#fB&1RYS1[2_4=^g:9cgGLO0b8BdDYR0YY]^cK^_Z^^[gKc:Mca:71b<
A-[RSf8QaMa/2U;7J7917O;UZCLX[dBPGAKHH25NYdVPBJ+XX&baKK>>UR<b+6BG
8[UW,APGEa7c4R&R3\Z;7Sa)]@2R^(f<-32ZVOOQ24/=_K4gED&O@.8K-)FU^)OB
&W,a4QETfL20+XG.(UZKd>O::SY=O>C_\&U^7EOK0FdPLeTF6f>EX7f:;OG3G#Q[
IcA]4]FY8F\((2LUKR:NadVBQ60&-E=cU?-K)a]PNO92.3,1U\QX.+;f/P7HE/fB
);_=3PMR0]?YND^>]>aB3V05+0<Z7-G:UaV09QOa/)L^<KbG(afQ;T<cSgd>F?&CW$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
HR9&=_.W3:31YbU5?C]4>G7ERCe2)_J/#T@H&6&Ndc+P>=SOV,G\6(/[J]JO)))^
IX54&[<0+UNe8:gd8>L5[EDTSR?COHc&P&=ZB^/Z<cYTa#90(HTe=@2:/Z<-_K-7
<d0Y<]+c80IH.(a6G2XZLCTg+e8D&HD<d_bda>KC<fNVMSD29U[?b6a<Vfg())(J
]aJ\cPcS^)#gX(A,&E\M=TLddJbYe1bRWgKB_eVW(\\Ge[J?\f_9#OR(1/<&PaKN
@R\B/AKa7C[aWM)3>Q>8E0JMT7=cE@2d2S),H#Y]F4I9b1NTVYY-a)=+d_C/6LCF
I,1c(_P83GP&8)g#M=UMX&X-_ZSEAZ6J.Q]Q29L6J33D2eWIZ,aDECLLEF@,X@]W
8_-DRC7+P#O..+/[2gc[Df2bVdU:R<J_=S)2c:2QM.#SY8c;FG,(8Q:P1-9O1C>R
>N>g-_^C1aPK8?&?7ZA]FTX=1&7G;a(#O-egY1cZ\?TfD-5SKN1XbQZb+(?0FHEf
,3PI+5QBFRZ--/[_T2D@\K\b1]Gc;G_RZDESYM00B6A7?H8=(8g]/RK1B#?e>673
JTSP;7PPJ4AdS[_=MAa7UJeX-3\(_&X&\PB/XMQ[G;VJ@71LT<S+)ZD60T/BJDPY
2F34@GC9NMc)3Ig1;:42:DSM@I#80FV\AZ9<\@N)T[O8MTZVMA;I&903]_&&R_33
R_)#:40E:]#dF?^bg.BNRTSMGb@b7&\U^e_+BV,0^E?@G-7#B0cF?dYUd4/RbU6N
<G58:QM2JH1^]#>ZFa[/afD,2S1#/Ib3BX1X(8>VL8PZ.0-&UG>aMa-A\05SSfc=
-ZYg0EL148.0N-_HYNHeJN,>MJ&&bZ1,0T+f/YL^2B?:PS[?>gX9#:9)4V0>Z@a7
5OAE3KaFC@ZfXY2DC/I@OJMa8+<9UJEU0_73c#&ObI4#OM5</U&Y/A3^fQ;,B)f0
77B]]&)#/(95J43\DQ21<S&?]]:#8E#\]EKT4_+C/+/0SSBT8QU:B,CT/G],_Z\b
cf##6PCM_<B,R@(IeG^K:H3U1RIB.>Q?\SG^0Lf>Q#QTKJO+eVU02_KL(UcLJ60/
Y^\\fHT9W2G1TS0;4:QU&;Tc2Ib>f-4T5G,_Q:92_(Jf2b-<aa\_5Y\-]I4)Q>A_
].KI5c#W]LS[U=UL<K_&4f^505Fa9@1PSX1(#_S5+-2>#2?Z5<RTP:cd2W./UGBW
CVAaV_#d/.\YfaL3[)(,d_c3bDK;6dE2@4F]J+\F6U@S/.D?3931Z>K7X=0Vg\gD
X40UQO4fTW]REB43=-/A(3@F[@Ofc]UaN/B5UJH(EF@N4@)fXa6OK1Y8a2IfBAWP
SF]gV1MH^TIS2M_^S6&8Y#.\RHW)(11[_F3(Sa8/=7><.3^@L5R[0DYI;e+.2Kcd
4GeYM#^Efa0YSf2;0EMSegV]2,5a=Z3=JH>/(98,0+](/4d_QVL6Me_KNce]?+=d
2,LR5XM;F;RQ)R=,>.E2:S#&HU5>>AOWNIeIg2KTU&VQG_Xg<[-ZcX9A@\feS8D]
6ARQd;5@\7G3P/L@NF8cbXBB82MG#-eKF&?c/\G0Ud/M@LWEFXE#2XC&Df[54cN?
V5A&O9eE)U8[aP1UW<V@9UED3;+1F9GWPY#<gN\X.D\(^MLfKSE)CX&S=83O5/0d
M:^0I[UG+:ETeeVg0MYYPGgE67#;6]95d22B^g?&R_N0F2PQ2Za5cE3CUH\#4;dQ
KADTS.^,Hg,fbI#P&03aMeQJCF=T)R2X-7<+9,8U&3U#2QH73d]?cPB&3FT\d7M5
UWF]>:^BJg[PEDLQTD:E3/<7QbMUVddTF#,.<O)P3K_0CgNA)[2.7L+LGI[3_YeK
:AdW]9F5)^8R8^V(SC(8H&@H<(/>YO;,1OQf.QLAd9>[+VQL&.fEF/<+V-(@UeWK
SI59/dEaO#UP0J7(<B34MFH95fE;8[NV[@eNCSY/&[1X-f5..T/Z(DN;P1+3HBBf
c^^EZ3f]@7@G.+C#dKBL)CF+(KLe>Y/e\LHXGR=HR]GTFRD[S@&\U9OgZTOA2GLH
C\KEP3U(^8dSdS;d7afPB<G-F1]WTB3gBT2VW5332J@&TTGgZC=CfH?bBTVWVDZN
_X[>QR4Z@AIG3_N:2<(X#dZ#c[+2K#U:#>JO3K@<gAUN#5[5@L1D9f>/P[FePQG]
ZJbbA_=F]fb@U0><4>CG-CM:2VAVM;QWcJg9NMb)\DJ<5,>Ff3AAEO=QSBYc/dM,
Ab-N+B+<Vd+39aeMb1aVbMH8e6S^#Rf0_@NCcJX&88#J=_@<#;AXZFKF0HRC:gGW
[a9,7=cP<a=BKD>M7W(PAB.EQ[^0JT&TBgAcD.)Z_N1\#CTC8V<YQbT11C7I4d/O
?F_HJZ1@0]fPCP_H39Q^ZBA].L7,4WRLO\e91U1.@ZW2cCT-abM)YD?BVB_VK(f]
X(<(,La;X]3CN8a8DPX9H:W;g4,AVe1SLfC1-Of_3>7bNd<H>KPcY^MN,T+fRN?M
E]>UA\>)f0<[C8BYMfe5E;T[:>P5[@gQT+0&-HHH5cEVX6BZ3#IY-Z46(b)WNgFe
E:Uf,TWd<<?gU4AU7:XX^dO?]=;]\,CU4-[U5+9^@VHWXV,a-&YOML9U?0##a8c[
3egE69DfGCB)TUDE1f81O3c1SWB-ZO],7HWB#6.])fg7d7A4>W>g6&e9;H[0E(D1
W)W&gA-+I2TQ_SKV0L0\VQ3.EKGTbA]-B^W<de;7c1FJSU1YG]b8YaTLe1FVgdJF
OY=C<Da,WGJ>UHP//>\d00X+fd+K-c:N65M/b@d-DW<\69EC13H]GMUB6[c?B=+R
]-a5[=F.0LL##KA.?_fK<GSN0N]X_#<);QC>Id[,.C?;B]7:82P7/@T?g^21QJ@<
cKf7/>GOe38/HOO-4/S&G[;/8[I\8L?=g@DG#Mg#)L:[0F,cAa59+R4AF&7\86>X
4[,:E^@^Z>9;?M@8gG-5I]=;V@&#H5e;bdc6LG0A,93bHS6fNd9)T;/GGc>P4/63
P=\7USAB[&\J(Y&Dc/CU+<dLI&^/+I/@]H8<d:PO(OCE,N&H9X:,d#[G)MV&8c\c
K(V?<#UHS0a[@//,E,JO,a(M?C(4FJ@9<8@Pb.]FV^KW;=bF8V((L:3R(M5]34(@
2:Mf]ZRD56HG+bYN,6SB5ad6LW_XLG<PgBd/7,/EH?FBX-08]<<G61OLcG(2+YXd
YW](KF;U9675+QeA]C/D6T:)23PVg14]P.L>G:(7UG(aMBF=WWK2^c^7gZM>PZ2_
PBLVg3+HRPRDM\RY@V](AU&^<#XAbY\?bM;IE72bXHT2+()N/Yc4<[1NJN3(gABE
=M_.ZM10&+EKbEa3?K#4M,3=K+GUe4[F:)eZTXfcXHP:UJ=@#O:3aJS-V?VRJDP@
&571RY[f3\V]YdMKYQ1fb<@Q=:dCG?SVZ8V/)0VF2I58I<28c(_Bg^#5JbVX1\2c
)VWG@-V2=CG85]40UfB=a[OCR?<;VBdgN9/NQNAeTB<[,-<>K[3NR\[JY5MM>3-7
0<\IJN.8>5Q)^AM4LUS6]Xf/F?Vc8H(ZK)D.d+^TO7U<:a4,6^:#b&M3K#;2&91g
+K2ZYU?C=/KGMRJ)@U7QDR92OP:1(5+PEI^,Ig.E?@&&S\_H-Q&?.L008g?D#]32
aR&U)+>1E7+C.HgT:GR&88N>T^HWA,]U<b[MV[4,-@LegDV;6aX4B4\f6.a5DI]b
:P6:\QafLU@7H268Nfd:Te6IPSUNY-7-EIG:2@-P]YXX&^S,18W5^D6S]b#7L80@
K[Y&W]][IY\8d@2=SB;YSO7P;dQ1O2THLYGZ/)0dgI3QBdK6I,Y(>D;M/DIM3&1T
d://VL?3gU)A,X<G.@8a-FC^R#8<Xd4S/Y5@??:PZ27PF;P=IbT9ZETZVfN4^TXE
-CbU6)9_ee2f&<aAI#Eg4dSX3SUODQV5gXS8O9M+U;ML.K6N33dTLRc#eJ7MTWK1
9OgIbTVFEH21NHfTV-O\4-e/AfOV,<W,(=Ha)>KJ&c4;)-<.SB4H(D)S403;_QB@
&/)WT^=97R]/D_N&b\SfYWW/BL(&-)L,51VO]YYYH][]M0M&1G)NOEHCYB?\39?X
D95[JHY9\Y#65M#Gc7PCX;c_\]_2Me/_bfT[KdG_;6L^9SW?L+aE]I65?DTI2OO8
Z8d\+[6V7MMTYNVg3WU/?Q))H]dET??7@;KT&JW7]XD-<HI+fA5fL)DVH7=;>P.C
0Z&5Jd)KKCR+B#^aHT;1>bW]4Cbb34f745YbFTV16Pb0X&@QRT[]_b3_+8.ZS6OB
e7g3b_^)(5-]@PICHH]JX/^8.W.NP,&V@SZNXN=XI8S^YHAE?FE4^/M]S,I+QE_7
&c_MNQY:IUWD07QH--M4KK[de249;VPCPJ@71<>G6F]Z0[R1PaVSKB4GE\Qd5dEa
/=MT0BV[SQcW07XM8cSS?YaU/?YQ&dYJ-[M1>5b3^,#[WP@[\K&cYP69QaZX@97]
#I3N+de.LHZ=WCOHRH^I&@06/OWR:X1T5GSJ,e2dJ:BgS)a\@1)a\:[H]UM.cKTK
&:Hd.0G]JPg16eb8a+_^FLZ>A1/E3O+XfGV_eeSc[3;<+<VK=(F[75\MC&cYPCbN
A6#Vgf?3I4C;:A&DPY,V=R-6C-&EM>@-;F7f[S&<fEFM,VUfZIC=X,RRN+2L8<UW
@LBCI)I?g.a?30HNGU/:KW2<#(fE^0G>5X\gf&Nd4fZ+RZ9ZI3L-F0FH@KK(aeO>
WU3]/._geZ2?#9#Z:KNBVX8LL4L.cdN.Ge3=(0/5IH^Kfd00X?_A,,T4<_.BKT2=
bL?,^K783I^,HT5]45AM,ZW2aU=QfQV+GKC)X?5M33,A?L.LTAeS?>-JI1U,1#V0
47ADN04/5C9RO?_]WY.-/dR\6.NA_fcMF<O9<U.gL&&@6P&c@JK]B&]UXN#[P8:e
C>#N83c+GVggTT=1g5W0#M5NU)eLLI]KGK;X5[ICAWaNI=8CF&EbC\.-]K&Rg@P<
KMTTeV3d__f]4bW]:EeISZa=O@cL/)SNHC?F#BP.W?KK15\\]f6:>eXH9Wg08O]e
HVCGR5.#)BgDe;CbQC6[8aF4HRLb<H:31]K6Q_:AY4H[)6YP)]8Y1.R@+Qc>>(45
f1/W8IUPP1VJ(\1f,:E#F@>?:>V#<Od\(Fa9OHag0]d0<E^4H@g5&Z2c_@]TCdeb
S<@[6@G2+NDGN<:\:bNQ.L>Z,)?;-C=-=?LOeJKUO1P^-]?Q.Q;>#2dLYKB1/c1W
_bc1ZSS=XMg>+]bO;Wc-U/:HWdFHIYLQFX0f-UA]1BG-ENWC59=]N.g5=M3F\a_W
TeU2,.K[5GV.g5DY[HfG+H.;MRJNM]P4P3e.U\FA[KZ#a4:NWWdBIagYOg/TK#T/
2.PVP]6-:F);.T,gE^6)#XBYVNGQ,II<ZX_D.?.bR)DeTbc[U,_Q9K^eIf7IKU<=
eUY9^Jb6d2;XV<3].Q(?eXfbA+NS?Ie[8(1_68-68G,0.BE[P:b/FaIf^,]B0e&/
5IR@K1+OgdJH3U3e)dE-eJ2e^aLg[H]][]3JEE#+-R0D)Nf+\#P/SH0H6IbTb&aM
9>@A,P3WfM@D8=I[O=#VfQ7E1[M^2Zga)D-&QESQ0IHHU3>?32#<bO_6.NGcYdWN
2&O#<M<L>?eTJ=XY?<dFQ5GLf8YV^ZC)0YT[^+QDEEXT?aB7I^e6D+[H8GMg7,?K
gC<]ZC2I+C;c1SO^1^/,;\;6J/41?4H8KJK5IFLV0A//7>_V.:fQP5_.A@g^W[^/
FOPW=eI56#N=Jf.=1?^ID#V_Z(89gZFccYg?PZE>696OELH3c=LHeOgCV-FfGDc?
g73RTXb_cVHREY;U=GE?]+C]9J@cB-9d#JR(/FC7d)_Cc6=CG\\TV\d68QKY9FWg
Z5RF4Cd;HN))Bf>_7/JJW]PITP]W1HXA3UEY<&AbBT_d[8)BI5<K_gMV125,?MN#
,O9d;,OV1=W\7R6bS,#)Zf>KYLDRb=0bT:E8FR.5:[]-;d=8QI0P8ZN3.AZ[R_gP
OBI[WSY#6:AG[K(Z7fSO,2-eJF+QFGZ6?B]-?6F57MBeP4<gVJb3MO+AJ?URE:X9
bU:cXAM\A49/DUNYQ,.4=^=&M;X98#]OSMNQ1_Lf14;QVFOMcc\V)Le:D],:bI?>
)),Ad3MTf?91QJ:T/6H@e_6bG9NCT]fJU]GI&-Q1T?QaB6,S&>W&))P0-8ge:Ca>
:F&1_R]ONMM;RU+8H),EN;8PK89B0P5#dd>G-e9GCf#X7IFH7>e)/T7G:Hg/^VJE
e^&H[QgQ[dZ=ea<FD4OeXBX+<5E:\AV+C>U7(9&gP+P(IP=U-N48G;.>[<_JP2-b
W)A/a,5g__E=S\]5>#S[g^V)ZMXfI>#9,Jg)Td+?[e]>RTdD#V9Tb;M0P@.ZY,MP
MVeCVK=K6ca<e:(DX2-@QGQ4B^LSHLR\)?OBR80][.7(\A8B?5d)HW584RN23X2S
+89[2N]a6=CDg0[+RDHIDA[gJ2cf?fa0WSD]+THgeNKVV&EQd<_H=C+5)@Q6C33G
cWgAA@2AM9=RYB+A(&:2(^X>aGc-J;RYW;S@4-e=8.<T#V\V&HVR[P65\7_--:RK
PLVb&@,(c89OC2f35ZI<fM>DZ-#Q13G(MC(_GgcN4>G>X,?^8G0L7Yd#34CNNYdY
QLD1G1-:2ge9-F/TJRP=/X\,8Q:b0SB>;N6QANF3^P9Ne5FEF&G/aGUGX-D5fAW/
K#,eV&AE\^^PC[VW0[#bC]DGcWH3[M+G_-K?[Td[8OT98SV,YU^,QF=51+cB05OU
AW&)5(MBY#gcb-A=JAJ^N(3@8PCU4]B7c4@8a^I?P/bQO2\/1c(4#aK7aAPW,BJ-
@B+Y=]Bc]EMB,/LIL&I\ZFaT\],5&84<<D)93,APA:,Z)M#6[&+AD4[KHJfcP7IH
;cC#A/2XbD4?4K\d(eXRa+:JcgGDSA:TDVdY1FC\K&TPFc)H3HDACB65C27L,.\g
D+F/SRN,5@&<CD8/H?4PP;NFWUEDO5FS-@/M#PLTEZE7J893TCB&.H(dAcCA<c,.
YP@PcM4X5e.P+LXWAg1O[(&X:3SATYGI?c]A\)fORgcLa4CE_.g5Hc87BJcA+JO<
^Y3&PNH&0F3,6=6G5(a->GKf/1=Q5CU=ZDH+79_eHP1VA4=V;8_^#SDd[TMcb4.F
596;KT)3K\dH6=SLF&5U1[G20Je)25JFF-2LR_I]bTB+SfIY47fVf9CR2[[C].eF
gff#>1V93+]eI)?[C&)gLL=G[f[8;?^AAM:M].Pfd<,eOJ.X?;XEcMNe)FYbD)ff
]\DAMC1?Vg+AJ\NV+Y&VEXJG]Ud=:Gc[.\@.]D/eFS#???W--\-df^,GFX511+[#
,/SXV-,1[a)Ref044V_>83LPag,R?CTBQO#>=BUF1OHRVX8^MT=c^#W5N4.7f8)f
</cDW8BHeHTK344.fH:5JZ9Z-\:+@&;Z[Q3A6&9QEc;:^cK5Y&AJe8H;UWF,3J&Y
+E0CJ]Y^EKGHJUVNXP5I30^b4E<N]:Me25I5,DOY?WJ;:[.(X=@_V^[&3YQ2NW@-
I#\5J,;(BC55IQ442UIF:3@3QcW<&QNKQA/.aOZ;H@^;-D6ZWbGG/7BgVO&>4])3
I7<>/[@4ZWJFLCJ@^d=BBAY2Uc#V<2TTd,TCJb(5+KEXC4E758J>XN5&](E/>HZ6
Q(4\TUG/.G6&/79R\+?)D;<#I/W\DPBg&7@g&WD0FZ7^bUZ3;ZIH\A5I1?T)gff:
@3=4QPb>G]g1IHV&3M,&D7OCL&.Tg=F4QEH4.D,OMLgYb[PPI:gLEKd)5#(#O]Qg
(XI(:H0K=d5US8(SQ>EU2L+\7.(]QN+9I<TGP4\c^M_C34=f1_-gKS9Hd:+VC.Xe
XVX-d&079Fdg]YW6F=15Pff,c.?5^I3d;AVWe9efbP>S=eL7T<^=^g0;LZD0GD<M
&7UEY/bC@D>:P?CRO4A9dJ\7RI)W#R12NUR#5fg/8<P(@^;T53,e8[R11F;O;63&
XeL@M\F;\@X9JC)4U]&<g>ag\YdJV3@,,H-:34FcJ>]8X3M.(0)XB:;6cVc-7b@5
VGB6VUPJ@NQaYQTQAT80e?ZO1)gKgae4N)KAQ_Y97]=CCNAPf:>b;d,IZSPefN]5
B)<3ge[1f0Z)cJNZYUbDGW?1>ZI0:eaK^)a]EL=V:4aN8XEWf1.RHXY?cTH_DUMd
,CDf2,J+bX9+LM1W2?ZEK0gC<6b8GWFgQ@^AXg@C@^Qf]AVd:egT]37,MU#bg97E
,>?:C9ZQ9B<AJ0@H;&NT/(,3OaI>AbQ1_(O7[@#49Z@U.F@3[/UHc\?88bKINO=1
FVe?ZJW8HS<Bg<ZKUa(&?)N=TG@1_/gM7Yc^RXC>S,EZ4_<960+KU^4##A?VfbN)
?YYZ88A69,RU8f[)E#/Kd&Of(F,QgaA9R[/H.@aDG+ANL\adU:G[X0^@B8/B;33=
+:NV,)F1CIUJg5TL?P9;;V]=e432YI_._YAF^ET@c-^QEB(K82#?&543:VWX4Kc.
[?(Q[dW.Z:aS-\XK_3:E7P#SFIc4E<N^UNeE/X;3HC:#+U37F)3]B0gPXG@DSWMa
Y+LWXd&_9&14[9JUG,f?ND9_daODHHTI;0/A/L==_QSZJZ33@;MS9BBX+gZB3/ZB
:5\VADZ64,KPTd151,6F:1D#YM3V8fRZ@\Y(91KK54;7gNX4G1X>N,E(+GA=/L2F
Xd^-aeA_<0X>:[>6##?P,USMZI=.dTY:d>H)CB?cAJV^74WE7>.(?a2=86RG_S^^
O?/XbLc]g^/@O]E>;ZdKPaXJVXO7;O7/4,V=\+;^-IIa18QQH(HdX-+-RcO-eJDK
B32K5LWMT&OMP)2IFBeKfbU6Kb3>0=,KQ^.Q\.Eg<c5S/9Kd0P^65Q#?=Y-fX8-O
;N@Z\^,NZ<_HZO@GTH755Q_HL3@:^I-CTIXKV[P<[#DIdb4[/g4=G>3,ISX6U9NN
UM1;&.P8VLUd&_J8O5,F)C(aIZH=8\e]b[V2.Ab[e)G[dT05g];?4-=#R]7GabaT
:4Y=;GNYaSDL3HJ&U?#OfaeA/H&1+2SRZ^GPK(7]IJHQ#3=C9T5Tf=DEN_Q+WKC=
=JGYBD7W9N/ebCM0c4(PV_8(SE0UM6Yad,]LSHJe8)MO<b7fVgJ2IEd7@W(GeQf>
W:D=C,3VF5C;QaE/)I^.><WHd(ISgA2<_#;HZ,50\PN9MT\WZ]C(>:P\[+b+[M)6
Q/WTS&5e5e;Z_g^M6/0H\d1eXRg]N^,N^gHC@>C0[IOd(7:I#4/?]5A_689.K[VC
V7X;B6;I2(:6Kg_B&)7=LM<M3^^Nb0+0PP/^-eH0W(IH(R8J6-OIG-;Ag[]>^@(Q
@-C4UPR<2S?154H&#Z,b4?AE[c4HA7&MN9gdG5b<M#.ERR9--J(eQbfW&<Q^GSZM
7U^>WPWY:P1fFP-8,,DDS&HZH[HDGTJ^9RF)02dfS8D5L__BEM6D4&[^Y\dgXNP/
8[WD8Y<D=IJLZb1#PCG_U+(J_B83KU=aAL8CHN)B+J>?UCFX4bU)g709/355V7d;
1-:BcD3+>W@,==0SL^\eNdR5.J8f9^F:QB_()J=A-XT[8eS+eDFH(cNWR83._O?Z
Q(aeTE]RMHK,YTEXS_DG<U)eeg[g\e_[,_1QfH2ZbOa6R&M+1dc9KfTLH+0PP-L/
F8[/SA;X)]Z<FLd2-SG/^(K=#B&]:IP]S>UB;_/M^@B=Sd8<42#@;CW,X5\BR]F?
WI&00VE-(B^_6F60<YTFT;fBbFU1:&W247QIW[,3:/b2+M6(_+HfH^+aQOec:^O<
D48IP[bZ6I+V0<<,Q\dT6WTZ0UINGG,d67-&5/BZI_>EDaQf>+\G&b_@4B+1._DB
YUV4_SdRG5\UVf3&cF=;;NW;GU=AOA:80UNUf9))ZM2_/,g^A1&O]60S==JPU7CY
PU;:&<5CcRH5feCS_Wf4]cZg]c+;[/ET==7CX5?YPPULRV/3>^@7a#,U\G:IcEOH
bM?7g#7_1dR27)INMP0I;S>f(RPW^1V:6_@GK]6#;?8GU>1^9GJ^),M>G58cA8[R
eDd_N-/7PQSY7IPSS@^4].fM&;9Z.;7beXL;0:65DX@C(F1+B+MKKOc9/JHP+461
6&A?d]3<MT[+J9U?MH[;...N6.a8&KUFaS\VcHHJ=5cKZG#SPK=OJ>_+8\;,[,CM
RV/De2Cb+QFaf[5_^FH^0:5=)S-[_14PB9G._GXV9=Ca2Q(86/T2D\(O[Me+)L5@
F,?0MUCJ,&^YMCG/2S&/DE5RU@eQ8a@@MFe6c,LKRO:_A:d(XO[WZE)LPGE7<&AP
K7a<cgFGWRbYfV7<IF5HIG[+:MQa:OdTA#&SLONEU&/V:Yc&gF7eUDT0@&_;6cfE
<g--cTf3[/G2T@)VX<^YQL2(.AR#D:d442\IE5>2+e7E+B71Fgegd]]fJ#XR]A0Y
BCU#8<PTT5D[6H_SW9C_;40BUX\P[Wc6LFJ4FMO?9::QJFJ;Aa?W#T(Kc.Lb4ID4
:S5MK0?SZETMWC6[31O?13;g7HZ15G]gZC,7=H7V\9B2N1EWXKa7L[f^MJ+(7J?(
fHRa-)d5M^34#R0C)SG@-Fc43ZE>UF>S^^/@e]>eWTP>N&?cLI54B((fC]C)SZT.
=BY8[TKS7U,R+V@b0YdVIVCTJ-.<b60OM-5H4XIJC03MQ<4_?\N7VC,TIY@A/>9U
HKbI4gOe0Tf9JbB(C[6-aQY2;B<:L0fX55d^M3NRMEc;Q+Kg^MD?c1W[P4C@TUI9
[L/,\VR08\&E-PTFEC24gW+?PJHe:WdL)8-M_-H6532UOd@=#.WC09?2Nb[QXS:/
ZTV)WO9ZBZ/&:6#^.eQD2)a0+B??;+N6(a#L;E\QGIG6#IIZ0&7.d^^g,?<07G@Q
IE\#HH?C9aDC6f,]])A5J\+XeS7PYYdVZQETgbPRKO5W8C?XY<g)JWF89@XL.(bX
,+5\6_PdI(+]C(;&B0DLcKf38g^1H1gH_,_D(@+ME:_/@5-K/eO4#gQegc;M.[S]
:-ME_.HbN0V<R.EH<NMVFFC[9DdZJ5dd<Y)=U@-LLW?LHWDPVR[D)R>0(AC36RgY
4@gM)M4O:XZR3g5bF#>8CL#a]Q(3/36K#KPbG0H3g2JDa8D-RM[W_]+BHWSfC-6Y
I40B2MYZ-GC,#?NV+OG?g4Oa(=f0.^JGa_g2N[Bd.^?\EH.@YIAcH,M\dCed\1)H
MAZ[BF0.&ZB]gHa_KK@Z;;WPFXfGWFO&X@^HZJcH(M-a&QI)gQU6=5A\<AITXEAX
Ogf)c^T1;C/8cGXX?VbT<eK1/f(CPK^_W<FR-C9Y3+I(798d/@afBA-2L^6UI+5_
D(OMFOOT<+NO&g:>&a3#c6(ef9N4B@.:X4dM:\<<76A165K>N,@U+^+DI_STBC\[
RTSN\NGgRdTI\bM9FDK;X5Mge<DC&8f+TMX@0[8N>XK3:V?3T\F9c.KMH\A6G:B^
VYQET?I4ZNNG#9?_81M)ND_N>BQBRR<4BPXEB&7.b=])UJfI>(MY2d)f\)<O@6F[
-Y6fH6:EKY7&3]1.L#6N0II)6MNPVXUEOf#G>:ZT+A:a+2=6YZS_JHWP-?YIE-O4
Va[5D:)M<MUE^E8>44M5)7+X[M(<RW9GHH5-]UZE4FIJFJ-WN=),74ZTI17HbHbd
bT\:LGK0b#V^=,?2ZWFc7X(eI]#-3-?0IP[R.a3U[6.-3OG4<)9_J@VS525V27X\
H&8J&54CK/7Q/AOI#GdfEYb]A>^G_PQP1Q05GEG>#LdWN/Od?>-/&cV^gYebV(cH
9ga^FC8840:cE6Y3)_4c2.^<Ob\1<+Rg:#5Y]G;MLdT+)CK9-3C]96a(?:3cV&BL
O@F:TH48Wf#RS#1UWAN)83D\[#B>DK=#Y<TA4U1a02\8GOf+WdZJ8RfOYI[_+<7g
/N0OJ+3HEAH@3MRN;;>RVWKNYg2A=6-YR2K>=Y+ag+XS:6B@_2I?+\=:/Ha+,EZ:
VXb@dS4<>M@.VLENc<^[H<,<ED2@75)<.19/JKQ;DMRQTL9V+3?<c7GN<F:>GR5J
BE50YE9\F?229=?V3OQ/US:=4.)/06/.cJ,2g-BFb;NI0^29d0/eU>;.(W-d3.V<
gL+b.9GFU6;g&4Z/A+b\5)#^N_HDIV6\C,cXOOb-\<[5UG5T-?]<K]O40>+Ce?BW
aO+-7X8BGJB[D5f?SRE@^bXgZ#3@#6CAg@WPfG:cP:W]Aa5G\@F\ADPS>1ZZ_M\&
:V3N=;e,M_QQ&^b+CK=<Z1dU;ZdUUY[&?eJG;].[9bZK\X0,X9/QLWQ?T:BVAZCJ
)AP][01Yga?3c.K>IEXPDJB8S,.f_3_>>cB=\C,S5HH;CA=EHU9E6_RNXAFg?5b/
Hf7e9c:BCX_[?OB#d#)B65F-KQ87C,6&.5dUDD53M<,\9KHXO.O/#U;]]1D6.TI=
X1OM^1>TA6Mb(NSgPHI5O>-6^HdeRV]^G#,;\Q912;P@LDH)WU@\_Vg^]>VHBE4e
8Uf35+6[IURVPZWEPG<#RW?DXdWDKO&XR#JX3BO@ddc9WJNN^__\YeO=c9DNJcEF
#S.f>DNCZ/ag9:3@e_CE\QSDTT0HP@Q6CJJ.).50-XfbEYFEJTM)5JI00,Y8E/0f
^PMg.5007#/[DIL.,K,)DR32XDc#IeI=A(a6,&AVe_0LX5FQ1CTP_B/4@.U)=212
d)?&;g(PMH;8b\f<I4/Y[BR)5#RXM=1\58c:6?A878fQMf:S]/KO?03FN^R#Y2ED
2g1)-G>3C]M7B&DZSMOI@e:,X]U8eeU@=&[CV?6U,5bOd(A1XRK#eb^)##g),aQ[
?,8?T(-g@)ILc1e+Z(6PLEX>(MVQT6=E):fdBWRHg)I4.U0Bd5/IXeZ_4O2YVSSE
OJQ&=fgLc5PO6/BV;4Ed9QH:>&#)/,5V1bCA-TC&LUEJKJ6L:PP]:UTCZWT3#XMP
&9bgFSYHB6(aRgQE:Oc3^QE:2aeFe?LX<GS#AR+<R#53T,KUQ-f+4#OR0aW,QLgB
2V23^GB5[I2L)bA3c0C1JE[?QXM>SF:0^^1GOSOT)eNX9YdS80?XdEAM74SB8aT7
2c#U5>#cC(4O/8b81W_7&(=VI4)J/6X]6(#[@H#5Ta<Z>M_8#g,6#aCC4WMC9AE_
W.Z/ZdCe>Ob946FG=3DZ#5<2:OYCQI&EC41g8;FYD1-RSU//UG_)/6&,FC6T3ebN
dId4e/+SMa1C&d3Y.f^gF55Q<?gL0Gg8f6MD-#<8=67_IXD:\X9(gP>Y#:PU-]Bc
b9fHQc@gJe7)JaX4L?V>aAB>?+LbJ.9UT^^:c]5PaO4[:>V7ZPER\2T?YAE@36Hg
Q[_JK>I_OFg+ZMA(;7T3Sf2Hc]D6E>c7)@CVLN^\=RESH/,Z.Z^Z(4C&;^O_OT:0
S/BXdYfVagg1_D@R0RKHF0C=#-VQ]QRO&<_BHf]IXd8fADIIK-M7@+JNTPSOe0?I
,2ADMAT5Hf7]bFEZU?ecD(d=3CX<?_;dKA2<4AHTBUL9I/[6_C5b@_G#<cbXSQEK
P:UbYN_F))-?b=gH1?de\HFeBTB<IQ1GXGLN)(e.8B6@3M?,Oc>/L10(6e46JEKK
?@H1]7bSbUa(&.8I@ZVbF,8G4[3I?O<ML>N\_A/<9f^PJQca>Qg/LHZ>c31(2ZT8
IZ]6)L3X&O-:E9_C\8+>RUI6_e6+0Y2a0T)0U7e)\HD\NBG1&O@cFDS7DTe,#aC6
Y+6FL/OEJ\/\GOTI0HAg+;U\:cF?#B78C7OCW>W4#C(V>c7AJI4^-gGDE36^3WFR
\>^NZ.#d+V,_\GF<H(6@E>[Y>Z]gA.7cd<(2TZ>S6W[5.2Le8(L]AI(=)25A(QG1
K]BKC)BZ)#[e/+[gBDXIKC>\aK8ELYNR,CGXBE)@YJfE)41#>5]>]OD]UU[c(-7A
e)B@20V1L[E_09(1>X.9/2D9(cDE&ALO-E9]5KUcKRN50).8#W,C26;.4D9HXUbc
JcIF]Dca:EF/0K4VI[85_faN4&K_\Ke:,bDV>^K&e-/\bf<M<KG&Z\IKF>,decE8
KgYdc<,A&#ac;ABF#\BYd0,NQOIF)7;1L,g9>7<c#Sc9?WdFD.PX3F:C\0U=GX33
>Z0RXEM3MgZ;2UbW3]M\8.8<;7BdCdc@R/HZf?Y76J&gGe1WSAYRJ7L3L)=E0LGZ
XDQMeMe<d^Bb5g+aH[7,e8M2da[YU4K1c=T[R>I2>5>?>@S0/\YQ@(f^.Fg;J#&F
Q;FRaDG2N&&)B]^gC,)0)eSR47Q;[@;3OOdF:4HE6YNIb-G1U.LM\CV\0HIVaKU6
TZKON0VZGQ,OB0-g9#=06]8M_LOVd6@I2]J#a@([;#;R@F^O>^?[=ae\,4^.H+5H
.Y>Lb2DD1+XddI3;<]f)M]_c287FIN^^H22OB0?6d1;WTR^3AYd8(:,J&)QeX5[Y
LJ>G:1H7O]W^3fBPSKU(.(Y0-a9d5&\RIPQR:#X9e2bOg/S11d)=:VbG0:FeUR==
ZXI)Q7.TdN=Z/2:N+##6YbeN@1DW,AD\=@V[\<)+B5;16&W7TZ(HAHQOBA8S2<V^
SQ/H1B=IC5AeaR:E,.(2?&N8=?0;G_)4V]-,7#)2+CT0<:[\1d=_+PdRF&8A/f(B
FEBLe3H7+Xg(UGL,-W9TQQ&;X6^c_CLNL)2G#ZZ^[d@83:4g5+TAVJ2S;]IEP1&c
.T):M2W=^70g67>4Y\<\gY=/.@45PDT72NW?c:+J.K23K\:TNK;[.F8TU[U@6=6c
K2Q@b^2:ZcN#7M^dFPTK:J5DLTGWA3:>/Wg>C_4c(E#OA9X96S6FNdZ5E1ZX&A1\
CG4L\8^/?.GbUbIZU\FG74#30_BO)<bB3E9QWR92):)IFERWRIB0bbUf?JgTODC/
BJCaB3;1[7#JM>c#X>#VOS4>3XHDD/_H^.1Z-FXcH8EcTI]JGYY:>FHFeC5XbZK2
,.7MJU=(LCX30O/)1-dfHf04F1L]SdA<3W-(Q2F3b]<><#2d6NU(9U?V62O29[Sg
@#;D)9<#?a_V;[K0;a++A(HUd0,a+[(A]fdf=F\NL-JH&17cCcM_AE0<XE_]^,EV
c6\-=G;BgOe,IP>e3AC<Z3]@d&75;.Q.IU8-/?bQfYVa2>aR&e6N-^aANB_48e(N
2;(6eN[#;>bC=#<YSFVLf?TYN[N))_KfX+)&@_EdQCdF-,HF:7RJTeVFdFOY^L;(
>]IcS9+0K])a-0O_<B^-9H-cK+6S[O\8.<JbSNP3ZbOC+X@:85)>cc><H49VeVOM
#9O\^QENgabF#Bb5:FYN^CD)82?B<)b3,XADHA,;QfZPFB]6,5^(;dYN9M[AU,9U
PaJHI1/7A&(baG+5&9cgZXFG]G9CAW]dCH0;14IT8VJ8^FP]?]Vb#K,M<PO-+_-#
5ac)^UUL:5aP,c>I[>cg1)RJ:@7XU;MFe2CK8Gca&b&FDUN_Y#3A@I/2KeF?TgGZ
G1K5UdYN81B1Y-bXEI,94^\EQ1fI8,2_->0SM5JG+SJ/c#3K?3Q[AAN\E=fD9[Y?
gROW]:Y-Rg97QfFRQ.N\9R<>d^P-gTe1#BP)KHE6cH3HVPe/c=K(;4VV7aA^B24=
6BbGJ9<=;PGM01Y,K<-FY0X3@#8.^V.HOg,BS,_IDQWdF9L&5CNPgOK<1[/UH+W9
BEK)\D]Uf/D2)LSPd0#0HPR(E_HNZFD[+D2(SDF-#VO&^M>#U<]/HJ=2.aB:^g^0
6NG36/^,(7@.I+GCcRB>9I@:DEF-ILdZF#G3I1AW-A=>R61-B:fe4N:bNc[:I(a?
eb2:^=UJIbL;:8CS5MeT78O.,N)<&@fAH,O-#aKPbc_FfD#I,:>f.Y.fH\V.7^5_
4V7&>-86+dg?BV/:&IZAC\,KB04;@(H#3?X:]W?V?B3NNZ@7Zg,7;9#,S<0NdO\[
L42FOaBJV)HDVLV#WII5&V?FKd#@J57P..AIZYaWJN+N8&9SHcYN4[.aUJVTYZYQ
2IEK5<3ZgeQ:</eW=U.IQ;[Tc..@UVf4W,Ja#+91?FgCMZC,A@Z7<39R^^9Z@4,:
C>5>AFEgb<[_\T>:Z9b9cSN[c1.O9-TRA#6_O([DE#:RH-,c\PL/_1RcIGMI@QCd
6&RQQ2QW-G_=F-MBaLWGI3FEc-L2L2BcZR^&V6?G(7_#.beW[=X0:[@?=O@92cc3
M<8FJ+4V.E;cR^Kb)N<KAEM7I/>He#d#96AU>S^2>_Yb\KQXQI7:O#)L^=Z^FUSe
RW^Fc8H74JNcZ4D[.KfU(6U+9MINSI0FGaZgCXT--SM[4YG&3_Ed2..UF)^1)84G
C,?YH#>-8>&65I08><#OSQ4S5#efO.DX6_UKCNZR=&K+?(g,,X(BG55/Nc,:3_<.
O/./YFaJW3VG[_-T#HLWYQU[L7,J,Q)Jd5-ZcLY(aU(&AH1[IWg.5aVcD]+Y0+XO
V5&.SS-_TE(>EX?5e1.LdVXC0>HX0FPEP35fa6+Id_E]c@RNeV5/A>3/Y9cJ7a,D
0c:LG(7=NJ_&JSU@1VG;aDc0S6B0C:ZfIDHf0]7B,5<,Q_6U-AAH<a[T36R@UEX5
#EGS&5&+E,Ue8aVQU5cSORM0:B63_ELg.gN:b<3dAGPfYJa]/VG)[E5RVSWH3>5Z
<Q9g2_eAXg=EI9>0E=gSf<HJZS4_9aJ3BfOeOS0=BD.>5NN-R.C\.MHH?5)1EL4:
7@=Z95aL08b=36dSDYO]8;:g3cR_&PW-[XS)LAOGEWZ-Y(KX9>G75/QNMfE>BM@7
\eQ0N@,^:PT1>DGc9eVKB/G:+<KDC7)ZME1:>OW(b,_ESB?IXe,b/[7R&+=H)8gH
WH?^F#>g0:8.)#J(IOJR\O7V+_#bPbYgL[/2DO38WaL]KH-267WRf?@2NFWfA&T3
2/gAa<ZO-9A;ER-:H9Y#(.VYd/?N7#[beV\))>>=<L&RNHP9:+\=;1X\2_<8@I9A
-_8=QAG,daH8EHG2WO=6U>g)Tc;SQKF-U6DX7+UL50WK4ddIA2T,dW(2&eFQ;bD?
d194)YPCS)ZK<O=fVKd85MW(4]>#=E]>O#SA.d.F-;]0DVJg;GEQH8)/-7M,KGOL
308(2c.B[)XH<I=,a>>?^;(:,eSZDUD>)0a<AS]7OD(dCM(19b[fLZ8Y:.?I6-5c
I\g@NAecRfc6<PINS>Q]E)g1/-=2/dL2D22SYGA^]/C\;2I9O\gaH<J4[NMBEH1D
\G1(O,LA]e&.&DG@JX/[g-=1XPKeZ07Dc5Jd7OUM51gXDc.ZIN)c@;,fb4#P/P6U
^:^aSc6E7;0?TWT1]EKF<JXM-@YZg[;9L3N1,+(\MDHA?4G#UCEW0@1N@P>D:(gN
\65E-DMUZK:VS;@-cMd7T9L<=N=L>N+OeZ7UcS<?3KeN\KRQ+0e^L^#AN7SAP+I1
FCf12e)+T:[?G@>SHB;;75>#.,b0RT9(@?9D=M13:B,ZN5]3O;_^Y+]W?R(,.(8=
E\Kf#K)2UZ;2K:39DNL4f?L6e+\9F9,K^O/737?XDDSFQO3G[e+QV<9LEMZZLR8H
GcLCO_NcB(g?>/S4>1M/JT-XI\39?^BGOMKF)BF&=IA;e/8eS+AVV_PQ2VP-YGWV
DV[;HGc,M+)?QcX3LU\H3BRXHJN3>;e^d5(FLP9gB5CaG=+fQBR(I]YXA#:;AJ4R
VLAgR28@J5-=848O4/]c+cVW>&?XQ9I;ZB,:BCcO:14;AM+ZD.)#+A)^g(Jc4;+N
Z#6ZD#>eb?[4)\^NX;GFcICAR?efe[2=L+RAM-1@ab\FR7L1YAQYf=Q13a31cZK@
]E7:C?J#=3U]gX_deBPc(G(O7YF>EK#[//NGUO^1VWb@)e;B9/KdZ4/PB?E\EC]4
U]?Dg:N#V_FH/CE.cGZ_ZO/>8Y)B.a_W?AZ1[6#g;M-6J]U(?.S9),EdXa_(>?.b
]Ib56SN)FG_bD>1HL#c4;U60XZ/3a#gbP-DHG1f\>T/,[#TD?S3\Y-LN_88=E@HI
g<@:F8E;7PU3Ve2ZHR/_TQ_?7B.7eTZ<BHM>PaS)IV4eK<7gQ=B67KIc:S[UMW+O
.A31@Ca\PcO,#)<XKA5WPOE8F_W7BDNaUf<?VQ:[)5HLYNgV&:D@OX=,O8g[)NC>
@V;ZWcMfK]TNF+6_c5?S)BN<INf&5aF2S1@4QQ?&@09Zf:WYO#,d,4ecHQY121S<
O.af;+)I+6#A&SdQ/@W=:;]Y/L-<]/SQ.f7KI#0eTU2fJ>cD0V]P72VXM]MQB7RT
WKNbP,E>eJ=^Q/Hg:DZ59Z<CR;0K3Y/C]P?1HVB+,fQdC.#4X>bPSS7LDc;L8]TH
bH_VY__4;J7Q[2R#g)=e<P=>>H>c/MA/&+>7S?\RC7_P<5^03T28L\=bS5e4AUF#
PT<&;5P9-3#8;E=-8GR:[YRUf5^bb?,GVMG3Q.(61;UP-X#G.\a:fN\<CXY?2]Vf
Ic;gP>[EL5<a8[Q65?DR7GD;LZ+::U\,]5?QZ@ZQDG=.cc]C0&PUN7Y^Q>PaGb\Y
[(RAEfADEV,BAC=7?L>S_WI36&WQc@2;@2<d84f0I,A\(R^>(PRg39/6XCY]0c8a
]65L=U1f#P6ZS07]dD@Z<V<P6DReFJ@I3?MSAIM=;RT\_SMNaBdC-eAS#=K4A@d-
K6QDJ/P??Z/EA4JWKDT/a@D6NZJSb+#:T;JHG;0Yd#CX?_\CbLFIO1,G)@gOU?0U
;)Q_-fJ8,LXC6cU8BI3P&E\XN&VHQ:WN?W:\6J1Uf&3DYVfR6FM?>GJT8[N,&8QJ
^7+f:b.<5EcJPD1MY@,_9eJ7@J)aALUVe18H&DJ(_9)PTd64a^aa3:OQb)RbANJ6
:\#)_\/d4[W8TX+DT?3,Y2A/JDXMXNKFc;PY<?.1_/183NdR\/QUW/JDOJbe2[-5
UY#YHG7&:4S=a@=?8X1+<QWFR.3dTbe&<e2+O<d.Ya3D1+UNCE;U&]RR=#KQ)bL+
S[VDB2g9XTZ<c8eSBfP9Y;Rb:eZ@1;<d45+\5H+1?O5:^[H4aO4QZDV4d#XeSXGP
g_JA_LYTe+WgRV^.2P_6ZD(0XQHg[0a1^a_7VSBX\F2fc[+e[>Dd,G&92+>RQ>.P
UP0L4)8?fg>XeD+-T]f,c[4cDA0F.gF\JNaP.dVVbM5((IbXg\Qab\QWPJ6e4KRP
?0Y;Y2O6/9(Z#b\-JX,b8]ER;U[DB?W_UAQfRf2RFX/Q#=(;)N2\HPbBIScVZ=<K
R)4PDQW9OAg:N8=Q36J-R?27B#C.]@B6_\?6\@W(R9e]N^VENM^4ES7aPL8Zb0e\
)bNPQe3CQJ3IaNU+MFI-6B#3/8#+SL,gb3;V5,>+]U^+c0g(<L1Q39g6M;?De(97
80a(HZ#W7Q7A)0X7Vc.#SbVG>&0RZ[9Ug.&a.N@C)GR0:4(>EFa^3V_HMLP(>d?(
-<O)Y5UQCc)IAP-9f@d2U^7#fZOY-4@2,bLcO-Y4b#J(G4S)2Hg4QB&@3=8N8g3d
M[/4V@gS)SAO2S+A#987aGXKA/R#L^UcDO_8CB_e7HC(SN+H8#1ZV#7c+K6JK9Kg
VSf?&dDYYM+,?#ARHMVMPZ7UBR9d>>g6[SIG)REKX^-U(.Zf1I+g;-(5T&1d\c[2
_dDbf)HEUYS^b5H0eN(W5RN(VY;C:UOf.0D\\[:Lc[J2<Yc74J4W21&FNJ)#VO2;
2+)fCFGNLXLI0e/UA.E=6gd]=@Z1Qcc16N/-.b)NR7EB1PB&:HFHTBdYe5H/1Fc;
#OB)=#bd+.M21>0;Y<WagL4WEW3MX)3VRQM=)4C)Nc,#P[,a))+_&8Qfg;,K_d)S
Q3dV9/#F3JQ,-,--bc2feF/M-14LDgCe7CeG+Cc>=V[ZWP1:/ZGJ=RbU/N/)1)7-
]1gb.//VDEeG(+IA5/,V-b02JBPI#3g,X2+&+R.eQeXS-0.50]E5XJH]8f,K2,/6
@+_/Dc5b[HQ\b;[@MZN6be2A^R9[3WR9EO7Q9#A7>79N^ZG79@<U,<?E7c4-cN)D
<Ob+LZW8;Z[KS0>g]B-)G;/+[CM(.eG+(YDe5.C/1Nb<\_<X))</D3/9^Q?;C1Pe
)=YYB]_=g,7W7#F=&-KZSaP?2(dNI2BEd9dPA32e.4fDF9-T(/9Jb77IL&;[GFQ&
<_I&#,:X[2QbYfd-,X5Z,^GY&]INEUMW2YQR5:MaSHd_[1)SEgK-H:;UV3TO6EO.
f,3S=7:f@GF;g49=d3HOD^;O:#P4@1JWV5B.QGTCXQR8/fHZ.U/09><9_7G+6]1[
Beb8d,TF<Q@>R7[686,)E-9C6^5aE):9<>)X18/CP.0?Q6IK/#bHIBL+UGdFW.?T
g.M.QcKT2BSd]f<4S#(M[+EQ#Yf,:AJaA6JC_4IKa]SF:d(MDe.cIcUC_e.-GK3]
]8DEO2bJU5=GXV_d^H_>B5I[IIX09P98X]G/(Ucb7L+c+gO4XE,S9_NZ<SZ0I=QU
21]5=?7\b,PX8R[UYNUcgfdAgW>gWZ?VLX;M61HYR>83^BgQ.B/3e\H4^I?>T76=
93]WSN_aQ\XV\BWeN@G<Z.^d?>\;QINLC.I[)?^ETWN\+M1:^A7^NF\(VMb3=&;)
-Cg]B8SF5+eEKT+=)?#SdN((TRPF_>F8-g=?,QW@&P1/#.249SO(4]9a54(;5S(T
^0^/5dC[;J2PbTHOgdg;?HOK,E6Wd;&T(gD8LWQB<eb#+T_-\+_c-#8TVI@W]V3@
Gd1e]O,7S^cd21)VA+M6;UJG\aC4;&TKP>E2\#)4PDN]0?f^e,8]b_KC<(Q^@KYF
21f2SaW8;=/<\/69G6O3<0^<Yc)/J<-fTEG)7MbgH3=>YWP6GeSR7S-.b,.MBIE6
G7F>C+)8:@>H#+#_66WcZ5OEEANO#?f\YZ^.&cWS1Z1([#MXbJHde<>TAR)c3FVF
df\WQ-#e.g2d>;Q>WIC^c,#>D\ROHQUX^]9JF+]SN(f]/YH5O&<J1VD=36^L5I&[
:8]?cG_8<Bad7AIMUb1^1>H/5fTQKAUW[O1Z<EF)O44-5-aJT^;2f(XdBA>S6BAE
#HP40IH0PXNDTZ1f_\/K-1gXbYIM=g.,5(X6UC7BLGE4\4N]I+_]KKKM?;UR/K,_
BLX+;P7TH^&P#@I]]YKU5BMUGXZ+7&GI,Tc&8?)e-9.eR6Y)aH7D0V9+FAOR(545
F2B,Wf;(&6]^:U>cCIfAMC4/TCR&+<7NXAP4/=JL8(NNFJSO<U0H[9@1:=G00<@F
_TA^f,V6/D:A4Q0F]^H-QPCe1G5J\/[\>78,XY7X=#.f9eeNaE_aH&3ZXI[N6-TD
-\K4C]N#ES)GIb96K[X6EB3IeDdG[a_U@JKEfFW2)5RN/gEDT441@Q](Y79\YC/7
Y=8-eZeB^#-S@#Uf-L;A,d[;Y_]E&3]&7IA;_@=D,F8ZI&J?7c?#0G\^W(6TFC53
Y06c4#QC0O[LJZeZ3_Z6QK6D\WQL4O:F&(JLJ<=)-caT\_375/6\9f7JIV:-8+gQ
+Zd\O6Te)&(JB[;8S>@.958U8]Q0KKBb.NbV?-VCfafDNJAO/XD&=LBTE95WCS>0
A84^B.7(7K1=8_K3P5P=e1+]-<UL8SCBO+4D-f]Y(QR1,1D990J)fe2d:G5<:#c(
Wc5L?gOPe8YG8O;UJ58H-NRDGc[8b,?/aQ#_OLW46M<[CEKWK[aR?TS+60bS>(D[
</3FL=f7AL6CG=+8E\9MPJ)9Vf]SPO0&;H(#MGEA7e5OJGB_GdB>Of,L=78=T,LL
cD,:;-1IGBA8a4_O:c8YB@<<[1cIM#WJCLW2()SO=R0K:7Md/J9HK8@<H=\g1;._
fM(eeZZW7aMa8_ZA0eNWGE[G+ML0VB.F^3?,D]<agE-77X5-=@8A[a((C7Gb]4?Q
V^dMfdV=-P.T+aDWbB9T#]>a)?:RDKU<MGV3>E^LIN)d5Y#H\=@WSL]_VG2&7QZa
5VIFT1;M2.1JHS:E)Q]CcPK_P\0S@RR/0EBHHZ,=7,EENBef?.[_4:^#Z,:[A+Zg
cT3GL3&RM<\A\<#<1U^RTJFJfFNZ)YSAfb?>M][a=YNddb6-4^<gRUd>\XCV1-/c
<0FU^e7F6F+5Ba6VHHIXdB?-EHg/[E);OOcX8B)OZNN7M7\^f^IWcEXAf\ZH,(V5
5GD8KFO=b5]_JZbf8CT()@R2+L976ASVOSOP@3ZC-^6=JW(3F>+NE=[VSfON:H9M
fgfC^;@7dI:2RS6aP@;/9OZ9#1?)bKU#Q;+.IY[DPLA(39RL7RGZFb0+Z5+=bX08
@>H@,[QB57Cd^4ee.7?Lf)R<Cg#SCf0JR\7d.ND+PPM4+X\RgY\4WaAM#\R[Y^6(
RZ&-d=dI(C(L(-^+O9?0ID1dW&/Y.Yb^:;[0:RcHCc;fE?]LG3fM-V.69S^K6.=7
2X[[+S4O4Qb-f.bgHCY1WcaG-_\</JgIPUe>9;+S#<dXJ99ASU]gMUdA\JO__>D_
8&P#/[F.Ug66PAe)62JHHB5f5c67aB23F>GfTW34ASQ5?g26B=>)4+10M(;PU=6]
9<0#:9Sc;6=Z=R/WCgKAUe_BP_)IQ6YT49BSc(>@0=Z;?M#I?3,GN).#+La0D#[=
J&]RY@4\0eMY#(Ng4.Tb0[W_=NYQ,,636EIL,9(Lg[bdSJ=He+d\(QNL677=cK/E
)6W)T^))?H?6[W=AIAYU?/Ff##@[E5+0=\eGDKeg:D[M<V/[W42WgUP\]-H:,1:M
CB.>;&?#(;6NAA^+,^\]eWK/K:FfY)HD/0L?80Y<,13=-f(X-5E9QOXbE4OO)dJZ
ZC_WFEPF6-<\+ebN2&RZCD)2P:&87#DP3#<=I7HK=.1<4R:80R6#XX,fNdF(]bKY
T1QRWI^8P>(<&Y#\dP1Ra.dSee&8(gQbaM-8QI>a9_3DSH\5Wg:K^+Q4OL(X=SGC
YF<?<F9gcA-Ce:?R,I_b;9RP&G=)5:EZc#?>0TAPdd8+=e3X9aP2H6>db)-bE1dQ
Q?dL3dCQN:2XP5[N#(b_g;;F<fT&LJ/d3dAR=9dYJ/8IANL.=f:CQ1a0]ZOUagMa
K_#3EMa;B5TF^.g@5D5+CJD<\GdAF&_bBA.gUT/9B-)AZ7]^N]3cNF=#Og>7.aHT
3EHWQdLEX,5gE;^9[@0Qgd@6[UP3AD&dB&;DMSd6aa82WY6#XWS/.01,B@K<YB0R
13264>(&F-,1DdSf&0@IANdW0bgQ@G^3?e/?LU_\WMJg&84O[TU[3d;8ID-+fa5Y
V3Y2C;edK\Y^@0HU5b@J^H1=JKeXcEB<->Y#cSXVO[_\H@NgRI][<bV.XDNEHc.4
3c@KcV+c-J>ef2#:(D]C#P0-gD4DSTG<XI-<:HK5BPN/SS0^,&#<IQgcMMZ.W.^L
[)+QGYVJ(AEf_W\Y]PRL<9>;HP1=NETUf:DYHI^QC/G>]HVA#H8SFT+=[RK<QZcG
VI3RKbH#U(_g<2084)I&GC1ef++@/K_Wd9/O_&L24S-Q8I=<-&M5WS7P+W7GK5>4
^I9O[<JTDK;EZ;PfbD7&.Ef6B0_\F.R5]Y44G9F(dHabNBNF09R6?O0BT-\F@4(U
b<eUOfdC-LFOACNL.8KfY^\a]3-g9\SA)QZ5LVHQbT@Z<fX9SPf.e5-&3976D2,L
<[Wb[@+aAKU?B,<N6_=e)f10&[-243]HcNf#Lc6CG-7Ig5GTb4V1eR2ZM>dEW49@
CS\,]K]cVc_OV2BXVN,Bc,3[PE.aMeLH_0d,e+^UVB2g=;752C5YX7H\5a0HU[IQ
<Fe(;H>(A(c\6Od&eE=DBbH(SWc.c17;XdM_7#-Q(gG@JK)e0G[@>EFWO7RA(D?9
0a>e#J3(6_JSD6O3cDVMZYFZ.\_PO^c+H5:WIcf70R[@O)B,9gC&C[XRL7N.\XQP
5W^?H)O\]]eANegHV-0A:#TD=F@7E3@>@#g-R2f1J1Bc=K[<Ld\SE,WNH4EISe,3
K@XDbQR;V8,g:c-H=M>-6DeMFO<Y;b+eFM6ObE4N5?T@QYdA1.>##/<B2;??VGcJ
AEVE0L,&JN=35Yc.6@<]Je9TPg4A:TWb\Vb.Y4S+NKXPN5IEU)\37Z85?Rb6[Pg.
1&Y^&+#6bbT?5IRMNRGXW26.EY^BW?QBf;^G>O0DM&</R=)EM\:K1B9GGM76NDEN
66^XU>FI7^#a]T[_Uad\;J41GAV#b^(3;@aaKR[fEc/1?8J:.O1=>?W_]9LJ.YYB
<dcb0ALX@9:0I#)KY7@(8N?a4I,?O359ed=UNVYW;XO]A9P0QQO?g1NJWFD)S,#b
)3F4YAbRNa1WT4)+>ETgO(3LeFCQ<Q6J^\J#e#>H-J2/P7AM#(1J&#b?bVNU=Z21
aPF0VGN6];I8RU^ae3Ec\G>/@/H9W4TKV17F^4BPUW8<BFOU]HF@L?1aeJ,DX9S&
Y,:O5c#;@B2_+@eY=RRR7^S87-&5F1VJ;)XM:fX[2,O3FFX]S,>3[^f@ADFAc]e2
dMKe>4#g_D?9=KCa@ZE-TY>/a&TXc-\>S2?LZNV86RG2@&H7Y,/7X>:LaA6.^Xe>
+gb[&dWOI8K.OXCJLe+UGE^BZK\1.0KZBA@O@,WTXFL\\.VO>/,8#>+)RU[K>Na)
B6L3R:^?U)C)8LU28eSLV8\:J>W_eM/=Jb<D?2Y<\1U22>>SN7[H#[]:b]UbRb4<
+[;4C=AL__O2^@dY3QK4W^L3^Pf6WT\++[]I]C918TDBQa+O[_R4,L>7,R602+AU
DUF7[?0\Rc5?O4&[(PW=.78bZ[BZUY&_&AQY<1][V36O<BZ/CT6PYF4S7HHSLd@J
XE)g5<T+[1]4c:;7M1#DB4f_Z5dQf,P._U]T6\#fWOdI9QBD&.183SedM_G?<@R_
KNa]FS)^C?6EL_(]9?TZ7_AKM>>L#4[Sg:_(W;>F;a[.85b\V@8GFBB^U>-<][B^
AE^VKHW0OXQc9DD7[OPWO_P[OgYE9Y)gcI#1^8JM?dBP(65Zg0W2Sbe\)WK[7Y4+
g;0_<@?9S9,7aQ7=96I#R-PWbKSbCcHD(>;01?9;>_YK#Z6D1PF5+I@Z0TYGQfT2
/AG+PY0gWRB400UJ98&#-=Ug._J8/-aU:SJC&XUBXRfEGP4WR-^9[^<AHTC;[PI>
G=AI1I.SUd_)\1(A8M8,SCd,AQc&-e&H9NJP7eH77gA6fH&Od4KK4._^K:be[)Y0
UGQVLI&K.,>O[Oa8);E/,WD.a=II/Wb1?Ab#-IF<+Z8c/M2aM26SNb(X?@TgN.dN
++R3GU_@d:E3)#O]Ub-<6#g?F66b,QSGb<B6&>0669QgP)#?\ag99f;KF,1.)HHN
VC&1YP,(]V4FV->)0YS(35ZUdOS:aV<1PC#>]_1]TNKNBZ<G=\_XONCH3)eI:GC5
M\;;I^#faO[(DB/0H+(8U&dfdNdK-VFWOc(OV\gO9dbZ4\;e38W=ZV1egIK>WcJ?
,+K<X9=G-9O3+NEQ0Z8\D-&./4)79=?9O#(]31T1LK([U@,7G-24;W^Z1Cc;TF5T
=f^/80-4GQ7A+5B@]2FIUE-XID?I2Da,4-EaW6V](cXW+?YI;)0W+:<Udd0<HNc4
g67Cb(>8g>>3UO&Y/3E7U?fPT^CG>D1]g6B6T&KCU&7F)1H#M)KF1(feGN7;-]f;
1I5RLT&B;UDEFWHJTe[RD,&X#a\XE=:N=>T[S2U6DOV4FQKK0:3fETaMGQL0VXFM
e<0\9fAIeP8.:E&&SI&+ZZMKA#O??/X,5Fed9DJ[6dIg3?,_/L7\5(g)HX8R[aY_
T)<eeFC9)3:CZTD:)B4.3YKff]0J5JI:^KD0Q=JIPXg8]bIL96;gY>E4A98(SPf7
O70.#JKdg9EG_;2DGI]V_DFC^#Z8+?O(T\Z.bLCP2gNQ+XKWMf4g[AEV>bOVFeN+
\8cA@(:55JD)?4:D2GG3X3N?:]YAR9<+_,7X:J@&RgGRSGBAYg925\#b&K@XaQ@_
4,\2K-GF\[HKeN:f.@JBSMYMg>QYIP,MA:6NAJKX_fSV:S;.0Caf5Y;FR6JA6]/2
-PdO0Ceg1R7G7+;&=9F_,/BA8IXH3M&[(bM^K?&@:La9LT;cPX[,d]0@[TB5/(EI
X).:TO.\VSLY,1QSMV>fa<.4^>GFV,;Y\MV+</26-ROc<+[?/X36FEd@P>gPNO+E
8EEZD7OWbF8\J2@=2+L^<5P,SJDVeA)/I4OY:0N@#)/FH6,)WX=IX(.3GO3PE/O/
fF_[M-1]YTe3dIa3(FbMS:W+e1GVC-M\/3ZVK:9I&0;Q)eBUZD2>#(S#&27_Df;b
c>HIALVWZ[PSc7#66TI_<e-cgPYHWLM+Wb(ZYf:4U[gCDeBcK;HX)5PV@7d+92B-
&H;<VIME<T[P:C3D+7Ff9XUIBg\#4=^76)[&M3>CgT&<-a2RN21SM;((-4eaR\be
_EURF2)5]c?b_^D#S5W&C/QCLH[a^-Y3C9G:ce7WKTS\MV^<S@_Z4[7,Lf(5a;@J
S9fP>JH7@F)P._S4MJW-]AFbR&M&C@c^a[,,Rda-GB0a,,>L]c?>>5dKT7<B]]#>
T8BId_MVe)>W\NCCFaMPT#T8?)D1UN\^.FB)#@d8W:@)6MM6^R88+H\1PM-L-g,U
P^d-6[a:9(T-&T;#Ng)(;2BYa4/2UTY1P&=V6U1c<JPe<6<HEP>G^SW92FP-L<X#
PHM.cd91fSfX:-DU6+.(N09_@&1#HYX9A529e8bOf<d=VHT]V0\H1C]NZN72(^\Q
07[]#V.\Db(\B<=^35-:]UK[f-S\><VC05eN4EF#VHR<+b<R[1^XR3V=fb=ad=D2
6KD2E+<WHSc2FL-CE:A=SD:(C<05T_M:SdS@W8X,cVQ48&@D5[PQ[X+[5>.FU9CU
+ZJN=;#];/UU9VWC?GOc[_3/F-D=O\P)KcUU::9e_7O=V6A/SgJWUCcWBg\ZI8@E
0VSMB_K:02TBK42_9[5^BC>@C3A@d30&6X7T?0@@X>-/<\a4&(VEe-O#aD<W<RRO
[2Q\gBR(e]PA:_=0_H8]2]2<JeWGbO&5FKcK4S<0K_fKTf0HH;^+05&CHAHS41(]
?+?>=]F.M)>QU3MB@#@>aB2g;=4(I4K;L+D^cFMfA1/c:NeU8S?A]O,2\T;Rg#8[
&Xa]6YZ7\&>5@-U#<>J[>GgM6W6A-T8VRTaXd4S=BH?:9WDA.FS0(I]#=5-A/0=@
3@GEPBI9E-/=)9)bO/3V44d\-B495L-XYc>NeIQ#8>AG\U56&MV;?Hf3G55.Kf:G
Dag;69\IWd\C2YZ68W7:.bTM^R5bPfIb#0BP1W@cOMTEb/5^)QMDPT#8<--KRF7#
a+SAYd3eMZ22HO,CId5RePYNC]M^(;dFPD:PMM3[BLM@6=cQ.CBT0HZ[&SK+U_/.
Z\GOX?YW&g,V8HORDM_9Te7E7&;&aP\K&?LO^U3TCBQ<(H#d]_,O+GI6R@J<JZ;<
0Jg<UK&)KHXZD[ZeN+AJ@(-_1FIBB8_MaV-7@g:D>O]WRV8#3SUHPQ?L]R4W0fV_
8]KD]Y9,A/f9?,HgEN17f53CA=dgQ:MWYC6I+S-0NbdFBC@a<<(EK<F_]<G>aO<K
2#dY^QF]U2IQ,^3aB<b36F_5[[f@OfM#.J1.O&[M1?CN:(Fc(@C21G>W([?:#;)?
&Ad2Y9,/_P,@>1NPJd+W?Td.eS_1S.Z^MRX]:b8M^)W;E<=_(DZ<;8KceYWcNII0
=PLFUePfAIa<,J/c59<#c>&G)2Habb/.b9]#@@2-JZdaDO07O0KfE19Yc<97\0-4
O42b]a?d+4W)VQfNKY@5W0K5/G+c>OX\+CS0V5a:^,,95Afg?Y@3(O7\5=Z\VDb3
I7G?0\=L,Gc)#=?V)T##Bg[3KV;=]20IDQ9)eF:Y.26Wfe/QKd30/)]5?H]S_?cc
S.HOM1MGS3/e:aV,#U=G,2,cEM7:>^.eY)(</ZW91;OT8]24#9];4LD7Hc6;W.5Z
dee4DT\Y;)^9.XUD\?QCHfZ]10/[>9JE8_;_f/>A0P+FXKY</D6-WP#G8Y2;HCeC
859.&LYVZO0/T8Ce39WB29EIQ3&6_>=]^CCDJN2W.@;L1)OQ1f5eKHfW7T8KH&HD
M:=O7KYEF88:N>4#O#Hc\LIf<+[]4AT\?[c\+UCZ?G2Q4JDXF25?.8GTA^V_Ge\B
f>6aW_O<TeP(<>NVgJX@XYJ2b9[1(4b]c@L[G\[]=AAd\b/R-:fE\(FWF4]dOGUa
CF1d[;^9]bCJ&2LX3R?.P;I2MQ3M_^&@L:/da>9A+c#7>I0<<+(D7(8aaRM>:Te;
5/C7+O;AgU>e;9^3>gH@3NaL^Af(C]0gcO07L:M.XGS[BM9+=\^(BabHU_JQX-,S
(TJa8^FIKR9&M0BQ<a6UFGe/(T)BSM/&a9W,:_6161];O-=>5=DAd,cFKKYfdTOd
EV[;Rb+Ea,V])(L59#66=VKd\#-)?<86:BA)VG-6>B:/=[(WU4\fV7d^(/Y_I+=S
FLQ#@^8^?M(MQ=Q/FXe=BMX7WJ<P6Q(6&OX/;4TWZ4:LZ&G-P=J@@F7\cN6WgZ1B
Q0/TXTMC\SP\DZd1d2^,O8T>C4-CA9^d.6[#KaK_X:/0C28Z6)e)@^AfT1ZD_dA_
U=X9<RNFD^g\HV\?Uc>c792,/BIW=A.K6:_L[G^;?K=[Q>VVg7Q/6gJb?^@RTM,<
G^[CQRBCcE@/3/J(K4R4/57;\@g38_?9&.<e;T6@@5R=gW,BGaK<J-f<V[4cAR+F
])JBSEOf@42fSVB2QS7Z)3?X9U=9VMDd#:(TAD=f)2cS?9<E:G\O^&3H4]DGPK#U
9.9?#cEacSGKUc/N1BfFO(,>))c290<AG[G#W4;56W;A0_OT8AeQ@ZMf-(HE;5#+
aRC&G.Z:6Jc\>6C<OOJgOT46G]f@2DSE?TK\GWS1=&RJ2OH;HESF633<J](1(Y@^
LJ,87;=ZD-10F[:P5C;VALX506Z9KT,M9WIVC&,&<7:\LT0=b4I(fd6,:FQL(+^&
5aAUG0dBfR-;>cQ>a[6(/#&IgL0B4PA4:baH^IE2<D<U_[.I>CQTW8U8>;5E;AgA
bB4@QZ[GgPM(a4SG^U<0&U-Y[Nf=McI=@V)T6dPSUX.?D=WJcH75_ceY:A7bSF[c
?2BN@9NgI,A_C=;UU]WM[XLOTdF5NdUK)M?Y\XDP.LY\f(81+KgfLJ./ddQQN7[I
QV&e&/5H8EO:+Z&MHV&T;043bHWg?/AKE8Z6+,NWACM]E6SbEB2(6.c<dL8+LZAH
>4I<O.Z7MH/PLIQ_?=#SeE]/e&M5:+ZPR1fS(K<0JfVWO1^<<P_>C+g-2UaE;ddE
IY.(2LO=TZ^2W:5d#.K6V<R<?WOU4T\K9)U-ZHd\]8g+/R^/;UF]4cSC,gC2gfYY
F&L4U7MNEI?>D<c?(g<ILRaO/8;PC65Y2?L]B/@5DIR/;])9BB?573Y;?8]E4EfR
Eg8-OPS#S428\Rgb:A)F8.b.1_[c6:bQ.@?HfD?U>\XO0D;Y]<WZN?-d82ERTO2d
WZ7-DBd@WJf7;/;?<Ma<fbe81dQRKMCCU8aU.0>CC#G@=-e<+,HdJP^S@P)4f:H>
W+]/O=SJ_O^6&<2L,#NTOAWW9,BRIGPN[&S:A>:30P&a-c8UY7/,/a<?[G61[.4B
g</PK^Ec/2[e6;J?].=7aFf9cgS),H8(DO5IDdgH+3;HTY:])]8-P8?eJF<B(J_C
QM3T@NbNEBW>6^b#^:L&X14D:&Fd6Ye3OfDAf5PJXB0f5-;ASg5/>\+Z/W6M>;WX
9I?EA<=3F,1YH.:_dE^QRRMd:,MN:O\#;ZEgUMNP/<3B3YGX79@OeF57AHcRD9(X
;?7b?3851X:8IbR?b8MXJ-DM&>Z#TZF=P+P-f\:X1?Ba/?-W5<eKK]OgcFaa^:\6
_L3^.bZ<3?QC@WE:HZBE<geLC(?\B6;?<^;DCA#Y7MTcB&IW\NLQSHY-=NTNcBX0
gQL.b6I&F;D84JB27(SJ[VKS@EcU4U#34Lg?6edKCW&KGR).XS2DL(;L/SME]ICN
#a>a>GEG&TQN[<ReTZ^f677SeOJB>Z\C^+ZD^EU,H@T>[KAF_1dI;?)f#+PFS]PB
/:-_CfUITB.0,d/^b9GB2>Y(<V[0(+ZIeVJHULGI7+/0G6_O=+8Ge09IH)f-^(1d
)3fV8bf=L4T/7#VX_)-CXH:#F@B^W7ZP)3Eg5g>6)VKfW/WCM(^9KdI2,G_KTEQ7
8B>[Gf9C<g3<#cdVa&4?#\@Kg[<D(<U@W7QXFAFWX\.ABW]9ARgK9@\#9PN5,\VO
4D650eU@Rf:G+2.;8-RIMHa4&Y&3FTP:)G:g@S+3;F/(GD/acOZc2Z,RI=6/Eb2@
(4Y2?O>5d.\YI#[XZ/1Be>Bb)F8342QB:aXK_J<?Veac37WZgA.)=<1@c=cO>Ma.
P,F_?4X]LQL^f3<01M5aU_7&YQaOL@f3_(+Ob:]7DU2G?]_)<9(J^^fQ[fDFW-_M
/SZN;7QN^KQ][Vg248I/P0g13P[T,J&NW/Z#0)Q;X^W8BE_MF+PaA-CEY-2d^M.S
+,9GL<UTc_e_U/A7_<[0e(D.HIJ=6PWRWUXPf7E82VJ#IW166=aDWe2dN6-W,.IV
6c3YQ>&4gU1,a\4HPdPXRf1F;EYA#RKO@PZeST,KD2VPbLZb]&3+8A+4ECC_@^HQ
OT+=ER,_NZ&dI]:3&G4&WO(5g<@EOMOSd)aCe\f[>V\)g:cYP^9-I>X(-LgLH=G<
K;/bCg+b)^ee)G_?g;3[&&g1S1<X#[>>.&<05gS]g5^6+JLTB3Z8..9W,:a\YNUO
NPba8LCaL]^^C,WO<HI2(0ZW1:-T4-LS8_,P@J/@,811C>XGN,HIE7D0@A0be3@N
)eGf3/5T,>^0ea6^W9:UBSSA:4Z6W4]27EPZ,(LX8KbbcU1NZfOW/;gV2GC;8NL6
FAfWe#A\Sf)PSAQ6\ALRIBWRYMD@XgF7bC3>gFEdK/=V;2C7^;BE\IH>Q;[VA5F2
><<DQ2A7&IM.Sb#I?C-;Fg2@]eF=H+,>PfZf(04745@BL&6?16+S=]OC4QKYZ,+N
6=:&bf3#G&]U(e.AH[XA>BaT/.:-De:,?UV6?P1aM&U^1N,L._;FM8=FSd8@2EWa
#E\)&N8G\dKc=UYL:-&JOOPVZ3>a]1C[.]10G<?>8b30IG6>OZWZ(U7L>^EPITPG
L,]N4A&88/dWJ[fFc(Gg2W(6=eaFK^+TIb@dW[&?ECg&U5F:@K.<3QI-GY->88#,
.>9B[\DO.Q;5;14T&K6B)e1cIM/JQR3JM-/0/2JXF4:X?R/b:QHAB6aPD+fM:K(8
=TV_7UFE_g?c93-HcJAf+E7M2eRJc?@9=^Y=c<D/[+Z@KM&CUXO)JR28);+@/a[6
6P-KAVU(c7WYcd2\RH9_08LL[aKY37Z,b8>3/4G6,fN-ffcE:N7081M6Q+A8d1\;
9NS.a^;49N-;#54dZGYB81X:1cF:D^8?b+VJGG\_S\6R4E+;1H(Q=:2G)IHSZI&F
#?g6Xeb3++/Jb-&0S5>^91)0E:/JJ,-M_gbY(#g@QE=F;)T5C[]:=fS-a<fcMg9]
:D>.bK55f4:4/;PW24R@QT7_Y2?6UN1Lc((2:U-V.ZCP6RGDQ5a\.ZHI8OPYOTW[
G36[/?5?N8ZHL7WR6cGV0e6?=Sc8E33>3Z;=Y&P[_3c^9)IE5]\+/d:[K(gc-(a3
P.(P=bfD1dJf5#Z?5/(2XS0>:0VQGJ,A-eg/9QP=[3#5H]R@.d>OCb&H6[JJ;#HI
eZH4):=-:W^#M?d/]4,R_\CO_[O)GVJbC;KWQ\/Q);6a<7.H-BfB]]dag^_5H@c_
8(Yg&S:dU+<I5<&)5@D)J\CeUI\^:gb_eRA>4S8.4OP;>AZ3(5_V)Y33@fUAKJMB
:B?@aZ?2VM1>.93c/G:1E5]H3dCa<1VYd595J4KP<.;#[C;L8E)>6#cL=&:2J15/
V_W-59>-D_Z&@?;+6^9?/VYJfDFJcO3>&1aSWa30NC\g^_C\@gIUcM]06IEQ4R#D
^f^@(P=,534J+EQTAD)Ta+@IW5&7H1&DO,PSC[0(c[U4+@5,T2fL9)dX;.@C[fc,
0IC0WW8]8Z7OH.MP7\;M,c<;HA8.MG)HC1@IXX\.]3(\cU-Od#.bJOVB)<-WA]?D
Td\@;f@DB_9#fLb&KXV9ML+b>N4aPTf,Z^#&6cdX>4gZf,&Lg4P0F4C2[A^<F\9?
7#:6I8)3MZ[40f)89Mc3AOP+#bXdTFBW>G&g,GX:MT2I#:d6E]EbLAR++L@0B9fQ
JNNV<&bg28e0T1;3B4#8S>->[4YC?Bf,)^#IRdD,A2f)JV0MC[+[]Yf08<F;R=Z\
5^T/L.]@(2dBeZR_0>>^a?N]ZJJY2-bHAX[a^BN(#JZ10(<0OC7(OTbXM_JB3bbM
QbTe.(?W\X^19_L+:a-_S>X_+UNGXR]4\dASgNId-ce&QLW1M.,0B\G@?6[Jb)]d
K;5)UE[K._@&#9aN<3,8=OaKO0,3X2&WCfTSaO]?8Yd5]ed]5,AdVD<aZYLX9NQD
4TQ_DD:1,VLBUfLN(@];Z21&JF?2RcPQb#0Q7FYSEXB8N9@dU/ULPE9J\(dFd:2L
7+J:G83Y3=9QPd^EX.JaQ&H&.@1TET5#F3@4;,GC83YMICQZ]4;B.5/-1&5&?&P?
9M5(N+(&XgJ.cEP0cJT5,V=#beE@^Q(CBY0&JA2DGW3C=@VD>R94LcRQ]eeHb&Y7
A@<Vg1e>3ceLR)LQDB@f+A9aHGD4]C6c@C^[68,7CKYcadSB^H_KFTQ2#7gU1N[V
AR];B-[>R=+PBH<Ze@XPW9V=PgU?/gO:F[FL7\X:@.Yd>82Z+I&W#1;-#WFY>g@C
^.S607):6A[.dK[&C,CI;H:2U6_/^,[;8&=\RPPVHaeLJ0c0U1[;C2ae3_\FX-X]
R[AeZaa(;cZ?:Z6Q9S.GcX8=de(&T_fMW,QPKd#9dgGX#4PR_[BKAJCYHE<:1.2(
GKO[b>.6J6M:\;(K\R&M_]Z3+/3&cV91,78A6<KS#a#B-?d4-.RI\0M[W?W<Yag<
RQ,+3O,Xb;H_:JO?@BB4#6<S#5G/@b/A&cb)]CV891>[N=GaG/M/ZZN0&TRaT,41
Yad]0ORR\+^4S96LZCP05V1].R2Q23VQ[TTA/EWPGAUM2.N@MTR?gK/QWC#CIWgC
K1X#1-D1NQ1+bD<.+\a]bT1L@KV.PT0AD^#Mb]G<Z7;V+<@]9M&W6-PGg\@#a:0(
Md18C]_G^c)5+/33CTgX:TMWf4>dVI7</VNfDa=M[C(:Z4;>(QYW?Q.<^d)6@W6T
:-BBc=?VG1XX6cJ36_0_IH&a^-NZ@H28K2G+QVcc/CZYc&G=\(7^>e3?GcUVY#AI
7MS<f@B,7ea@;XZ(=RS:eE&b-G?4A,<R<5gXgY\?Xf1_,bY=4Y+[gZ+c:K715>gD
P8d,+P8If5@aYZ3FaJfVJVRX,(L,,)W-CAZ03)9O\9deC1AG<NDg\84:XWUGZBeL
&W#L<C_&XU=O>6;?G/Y6HTeSb=L99BL.3ZS;Dc+B83e/96c^VXM&(5HA@5-_9aZA
T)6V=]Vb1.UcB69)8B_VOF<#0DL/OVQBO&\;_L-gQ>-XV3Yd(L4+0MP5[(0B3T8g
,F\^@Zd2@Tdb(#SN8>2[QD_Cg0;Vbd(&dFFRbV]a].5_BF;/dW\d1D>W1gH\])..
)e81EPETT\TA6,W_/Y05;0IA8AX77)51)^_QAQ6)c/7L-0_]2.[H#,?U:NN^94Je
GQ2]SMG\edT#Y99_4O5d=348/VU](UIcO,IaZc#1f<TTX:\QMec7I2GJ:eDf_cae
U21>[ZQ9gP#CW5Q7S[eePbAdJKadBgAW/6+9>>3+V(4cGE.Z:/L(Qf&6=K9.,e0/
>)L=]=#1R0;Fd1GZC\PBJ)&;N,9VeOA;DCOD.B#(7K^6fE/VMT,4gQVRY/-4,.B;
&C..(dCO9:2XfQQ[bU]I&35.[JadV-#)d2G#N\(GE:8MfTB.>S&Z6@5K-/bC3=R^
ZUU,AaT6a#Q^311-AK[K?A4K;d(H&UINaf8?G:a>,)8NVKa4>:5S]=U^E+Y^(=.2
>&aW.U&NSa+WL#S=7LK505[8<AS?\^([O3<3M9L\QK:aVW[LbW&g#0T&]:50(KJF
B;A@d0&)-ANCfca#/L[0S(+[2aGJYX:Q1G_H1[\VEeOc9E+@;_G7Q[]V(Q984W,]
J+V&QX=<A2S]5)_bbfR:7b3\3ZeF4Y/ET(^.&M.gFV-/BTKC^U77A&>T[GY\?PP6
D(BGG\/D.@=VT6BWIO\dU>O;;AeZN;RLaZKGNAGW,<AD<AA>Y6W6@><aNf[9#dCJ
_]=GKf)MJO3AU<<JgY1aTS-8F.ab.g>R;aFMX8#:2?7,g0?^TEJWIgL4P9dGZ]]#
YaL6,2Jb/]<72,]TS=b^Q.^,U9TG:\2^.2&(64I?e1&,K=e/N][Q1A+L?RaaefP@
M([=F0MZb=Gac6BIK&Y@-SYJ=\S>EFFU03;)F,,]8FfN51J:+)[J8J-Xe9M<O6^=
PCR[?eA7IdZ16Z_Z<N6fa/]NQV<AH+C;T=.;D1-5E:BY>\AFRKe<e>dE?1,[AD=8
&Lc3;J(Xe.f87d=aU?HH552e-AZ6U4_.6>]/32;3/NR3[9T]CHXQRD>[W#QTDV_#
DUTF[HU<]g>3A9.ce?P5;TKDUQ9S_R1./D&aAeBPJG6MVOC@:1#V_cTTKU&9R]RD
(Be&(GK+VH(\5@F?1ebVg&\EVKYO3[ZAFT4.6T2,IN6DCH/?)1&@5R,Tg)GD?4??
SC&\+a^--UeXTSPW[8Qd8MX6MD:F4;YF#@+P^#JICKEH-AWg;PYB\VdgX#QPH&Z.
T<[@2++L[:CE16<>=E+#CFe]IScACC\E9R-;)W0D>.-.,3ed/>ZL]7R(cdL^:FDg
F:+8)G=+c2M,cd+,Z&H2_V319UYSRU)\g/4^T&-#_?)/gXgG<IE-eT>c],F[HY7a
[M=D6.@gCR?I.#YeE/GG&Ccf.>>DZeYXbe5QMd&Q6EXI7-:,(HH;+Q3,ZSfM,CDd
8D76X;<Q6?2=[^ET5beN#77ASMMS(H6-VcB)?.+\RM]#;5ec&4#5:(=FSPDNA\&[
Y9XM)IY&ZQ8[UKa7OFcUI>Q7<=7P73KW[6LF)#Yc/+>OV=LN4MN6@gOG\X+]5?UI
AYK105cOF+/MA3]3(5B[F07Eg4J)42)#]QB@>cPMHY3R,<Z]f&=4=(,)5FEE1B.5
G1=4de[UX\GF4\,;I2QCWV<:L(4^ZH;O4SaY,MLa(F^dN1cU63H#/-dHX5J;.RW6
34H;dNJFWW[N^ZD11d-KdSA:+RA?;11<9Q)-0BD3;cVOOQfYV=a34fDG-#7SI#]E
LX^9=7EC.bb;NKf3=V4KB:N8I<W2.I+Q0(>UOUCA\[^3b#PCC5)D(DZ/TO89&bgR
KM5&?:PI,<^<I(N:ZEO;G3TFWK1-KAa7IbZ^(/CWL-QTKLI;)<?=A=XN[3KJ9=V]
&44S,,UTeAMeb01?39ZMBK02fK?<_Y5.VXE?BaZOWYHJ0JC.Z[A#8Y3U#B@/g.eO
Fa6#=9>N>^gG=SUVBQ&O;AaW]D.c4G>XKFPXMIJfcgU,S.J8]X>W2eC;&U6H54?7
W4bRcX,\+YC9/]2&K8QS=CJFN<g]T1WI/P1OH?Fc1R/_#DcP8@,RVRB@2=NK4RYL
c/c5c:0MgK?+?cg?THDFP-A2=G.cSR/F[Da&GWWOL6PbM#c5[.KHXSQ4)b6f;>LC
YUXaN6<^SIUb&-IXCH[>HV#Yf-@cS&d>6]cE@I;_0F+CO73>J_e^gb1:19?XU0+)
O>O(aZdGa2XI:F1D)JNFC#fYC<1_4.>;e<;d?51.e;>1N1.W-RQND#D374Z#-4/U
2eaOD#]35C2eHV]Ma;&gUW57_#E_f?[-&6-^:[a(Z>c@b=97IONYJHc+9P)[,N)f
A):;RBX0MJ@LAWH+GN)6Ke1&6TSGMN4MFV2IZ]de)Ig#YACc2ZZD#KS:JL^R3T3Z
X\6Q#@QBJ70bHJ,P8c<):C9eg:ff-WT3dE.>\+WFY^^,]?EKX]B>S=P(E0GTFMX/
Wa&H??RQ?bWJdD=T:cd;S/G&(^Q5+cAS#-1PU_M-6S[Wf/@#G9e5-E<)]B]Wa;QW
:>8TLaBH/D/2LNd>TK>J&ES41]YYL;c3;d4\R=K2E4.aN1=FV>OBAI9SQQ;<;YUR
SNTAZ]R7NF7)[6[EP7SPJe,)b(&0]e^?Q??M@V7L/Rcb(&f,8FFDX\-bP:JM2/\3
V03[M10H9NF?M9WYO5TI-P5RdH(,:^\B9[+(#L]Q7)\K#UNZSR9.).R#B--SZ(RI
E2ONKgA2I@08ZWf5bOcg5XQ=cECF^B>#DTH96-Y)[_W]JT4BRYTaFCZR)]Y2T3ZS
\a(QW8N=&c>8=S2D>7.,VYc<Rf]VG4ed-f\A<?L6fYM3BN0Yf9WD:9SKTX/K8-)G
#RS.5S^[-W&,)S[c8#.PIY]dFQN?aB>eNH,J;#S:Ra:HY5da]2G1<4;RZY1W+K=Z
LU2S)MC4\BB8f=f1OB(OAK:SQHDELPWAF-:I8f:\P&OMBPP+V6Ce#[UIbO?[KG_S
.X>3D6;8SfdG)/QK@3eWKb8S1;J][8TX+F1GLb\YF2_NUc0,AQE>]P2/@XK[?D98
9bF1NS2A6R[PJ(4NMdJ;R2LNX:#:5V)H9d\0[W<d7^#MHaU8OE60D@&a/MS#Z)U)
F_RD[-48U(Y5AXQE?&>4Nc^/Q@@b#Oa48f,8Vg>;=+W9.L=^DF54)X#(DZcf_/^:
90-3b+NP#M)3A:S_9:>Zf?2b4CK2^R:1VJB09dTMdX\P]394<)^7_Z8BG?QX>b?G
[M^KLG)(J[]Q0JY8Z/<GQ=fF]eAT2TUEVggc6O6C#3MAf/5>2Z>)c=ZE]9Y;g<S4
;&;VUd2#UV#b]IJd(D/bYM0TW/>ZB,2O?4]<7QGQM):Y-C;=I>-NHYee+J/ZXW>O
L9:W]fR2C?&8K&OTAQcM=gLBCV7(PK0FQW<I.T2X/7#DA_12AAGHH>3PGfHJL():
MWPAc[cd_Vf<HdB,_,2[O97/Fc+Q.7\I<]:+D=];ZG,)T)Td:H8U+XB4Abg5d3/:
Zfd+;K/H1^3&.:;&dbEgPN)3APL.2aWO<N-U&CP2D^DId3_b[Z#<SS:/+JdV3[YD
dFXPGZdG=a^SU&Z(deGYJM51LRK0ZQ>X;XHG#L9^^<\:1&TWNg1QNWOdcH@ZUcEE
[Ae>eV83gN]I2Ved<=^M]2W>OVb#Q@Zc>PU24#870I>?ICZJ@7@:A+_]\b&QZ;d5
T,W7UVeQTJD9.)/W8eF+3:+cYO9(8S#-BUUXSFJ(\N0EY]Re.UI252+d]C^>V+&#
EQaG/Y99,E:K&Q&,<^GcOB:U,[HC@e?)]-eMU7WA9CI+.O^;VB#W[0WIe^VY_8?g
K+RVK^J-Wf6BRI_EWAKdOQ4VGS-Gd>_2C->6I)KHPO,5_/UH&#NGLX.C<R5bP.GL
.QB=W]\@Df&EK8W5-3b@Na:]]4MX@Q.XAH<YB#BeFK]6^R@T8JBR6R7[ST1[AV]2
;UT+ObNBZ(K=T#VR=O<976:=UDDB9F;S20dP4e1UPIT=^M:aVR[:A]-d#X>c>dF(
>SE4cQ)D5[d19Ug,N8;HK&U/9>MaacD#AGNOYEGE^DWNF<SIdBaa=W\K]=O8^N35
0O0<V^>ZK)>bOcT2+?X=.:O>aV>+c>V+650Pg6UR+Y<,2LP2Qc[[-1e#5Ng7YK,K
I]OaA^N7(T8ULWK,NW7?3aTG_VOPAZ,Y&#;<=36a9,_O3TD64#2B:SNc2b?WaP[9
JeOG2GWW?WWgKKIHMLRe6HV-B6]7aWCcAO,@,TNR_6>Y6+2L^[a8X<RO+7ZaQ]R.
NWO90e&F4A\B3#:c&Z9;4dTPd>=>3b]EB-8?N)3^V2CQG<SL(/)>,,7NU6M8Gg64
IM(^&T+e\dC&7F7b2IebY>XOK.6I]T6[HdG^.bc6LXa-O(5=g8XC.88STYIc;CYD
8GR:L2PW1Z4=JR7_Gc;8PW]9^8#Y[A7C)42Z2P(U]=>]-^SY8+7+Y]1)(CN0.H>d
L<Ab,8?8[>31D>TJgb]3US<JK[K\HA#)0IT[+,,1cHa=c+WT?)_^4K9b?S)PHP@A
WYN>:>40Y\4ET8G/ZF6R/ZO-P7=2&C>.C;c/E(N1KIG^[#A_Uf<5SG2,ERE[]?)<
A<XIF\J(/&ZfU#2dF1BW&8I5DR(Y(0AYFPDNI9a_TcQA5US4]@J(JJ5bbC9Z5P;&
Y=AYDQ&cC.Q,[WW2cQQ>ecb>(Y6:>B1XFg15]+@)bZWN42\BR]<bPNF#FO]5gK0>
9G2G2@Eb>Bg#ZE2.3@E\Gg9V,[N;\20D^F1<@-PKaQJ<<,O99NT)TP>HB9OP:6dc
G;-2.3J.,?cOJKC_CKbdJC94gENaD^P9T&MG4IW3TAM(&35)0,T)(<XS4g[:_[UP
L;6@SRcZfJ??L,04E.XHOPVHPEHH;7]3caJFV+WK\;PR^)98FE/.eQ/#ERTI?F35
&K#6IJaW61SM=6\GUP#9cL:X^gZ28;^CM)4VT5F.0X#\6R/&ZHaB4aVXP+aX/f[Q
]_?R,96.5gZ&#\<4^c_8@8(]b0@YG-66^eB@C7Md2+LYCF)bL@K:-,+H@9,f0NJH
7MMc0G7C(5:]T7b55gMgQ;MDP(c4Y+5\\NbZ\7&bC-&DVegSc)CgV)c[,GEE7GM8
b?2S08+RP^WYYI,_F\^X8(WDL6C>HEda8Z=K:aHCV=+HgJ.?T/bA;CQ?O1)G;MAX
OLbIBJgHOJWK?\7(#0Y9PX.]?:eH#8G=36?E^_4\>bU)fdgF.aeGJX.1JX(B5AV8
.BK+MDf--Pd+8eBI4c76URf7;:L_CD)CYAKRJ\@+X\4?]3?Qb)5Ab[K1K\7RE7\Y
T@1g7Iag8H-@+g^(dNM39>CL3EFb?#;@fY0<8-WQfM,c+T<^JY_9/IUW-5,Y5C54
g[W&)&.EO1].9PT@K+_6D?Z=B[e7O@6a1Od6=YXOI</P6&&;^.MDPXcCIT\0-D72
gg/d>=>:P]43CG>YN0<FH;=OSM#FLUSEBVT99-.]3SU#Z:^)f7)\9e#VXY^6MfB_
6.YT9&14RN1<^bREeE&\f+MBb072<d38Sc\TdBP<Z#>S\,Z5URL_;4NdQAFa,dG:
HD5@62)TH..7FCBJ_15XD1AF-3,,8ZHbMd15Y,U&T0GTYRGO=ENDLTLU\<Q.,9_?
L#\Y<7TUQA&ObY-MFg0@eN,Z([G3[=g?3+79V3&4=C/LJ>3aMLD([3HcfQ>9M#-L
/ICM3QQfHQETgGMMdbNBED(-TU-8I&/.(S@?5Q9=X#3G8Na.fU3T.a:2f0cLQ^HJ
L/QfJ@_(da&9XFH1A4:V?cBd/Q&E[AKN?b;CK\/?U2]HH6e3^.ca<T\&VHPU94.R
#ZH@/8bK-+L,f2].R0PU099A=b759\-+UA\R8CA-5]ENc;R(@1\Z>]SHZ=1DSQJd
(Vf)EY&EFfBNV^[LI];.WNHHag)D.2^XOc(0I1^e5?63F4<\8MWX>G)^>UdMZHJ]
^(=IZe=?&(<fP\F4TJ)JJ_/B9#,[O>4VQ+QXLaMPd#><bG:H1N4)K7MKD&_T7R7J
.>@C[H09<XA.ELD09)=?:5X5246RQ=O79PIMf](152GO41c@T)C1f;2@ebLbO8]Q
[FA)1POQ(RXb7J0W^=>7WCO,S<3]0G,1<&PZVK=AO8W5cO+:)T5V1c(eP#dZP)ZB
@DCGUY1RB=6Gb>XQ8GF.D^gKR<IS>,0[P?<98N;R]#8KR/YgSVA144I5U01<V3KF
;;XKb;Z4DM<)Ec;),UEdO;;;8X&;9/bd?a2&Xg+eGAWUgE\=GS2HZ)E+8CTacZEU
QBXP4Y&OO=7V-,d.a@7L&?R3NH84Ca=/c7=_4RE@&fHHcGS:92Ta9@REfcPC_U&8
9H1YEE?ff.W\b\X=FL()f2H].-N9@K\96c2b@]F\6MGDX[;56c=\G3(F;JZBP8T[
)\HK<.KNe-A1F:JS]_6O)A7NG.L[^+JLVB>DIb83;4E;+6X\e1CCC<7gWgRHN[6=
/V:X]=ZB<1.PRI+^b5fTDPLCE^V3_(;<],e(==7^8f\d++M70./..S6N<G:Yf-[X
Q51bW+J>#dP[]+&LDIC7&@NGPML0JC#D6OgYP,/&NN/0eH1B>dbTWLMP+J]1#[+:
f-&:MOV@Rf[aZ0G&5IJ.JDB#H#-I4;QLI\&^O>/PLH[c+9IC8V\g]]-=GS:@:M4I
Ld>(\=&\^^9b>5-g\8e3H(YVcc1O28\4Y1-LFQ2HGK\NJgW>&HA;?>BBf>XcaSD4
36&9K<\J(0M9]?L+S0KB7(@B5Y]ae5Gf&2#@E5<@+a/YF;1bY.d:+#a=75gOEALa
=<W0)+c>I)IN)RVH5X,Rf-TRW_]QQg9ID5E[436(^D[4gMOKZ,HL70<_,4D+[V2X
538=NZ-P#)IH)@&_^cEEc4IDG8OU<cNYQ\:[G16a?W-)S)DIG2QY:XH1P3WMeVVE
=C^LRdbPO1Nd:&[/EfRS_/U/a[N?.B:OScL2If:d#1cKXS\aJBLH23_SE6dPHSfN
K[;2EX_OCV,EWMK?+OcG0&ccG3.BeMMc9FQMg05:W.5K=FZOE;;cR@FaEPS.AR7V
e6F,43_1J440Qc=_H:6B]NcWgA0\aZJ,4F;S3(C)d(KG(G)1RHTV,PQ)Y>a+B)[&
b#KX7&3UNYd^L1+>2161L)VI-7EO.XK9U9R+U[&cTP;-#^@FB(>](KUTR.6NQVKd
1=PMO-9cFP.Z>.K)aY/(M+T-85eZ_+DP:Q;XRUOFF-BQP>5&9a62;X1?</]7Y-aB
cgY@1KD>Z]UC_Ub^#U#19^J67a^F=ZAa;^#X?a\M9M/7:C\(Y2,/CFJPHA4R#V4D
df\TL3<==1CfdRfeB1-eGP_Xf1AGMQ)#,MA9Ag\FMRVREFQ^HO4+<RB(O7]5gfJ@
D4NVa+&Z?S7A==AE?7gYYc?JS=SWU.THVeJ=QB:fd&A7>F?ADD<V<:116L3B^XW6
ALBE<AGMOfLcaR6UID^<1(fRFIFg-83QR]VOefWC55P6aMX4PWP>fV)0A4W3Cc8Y
#;_ZS#U>9-DG.PcD;90^GS\L,PKA&X5d9NKKAW(6Y7gRZ[K(99B[L#+]JLBHdHM3
Q82JSH.PMUe7(EC>>GZJGJ68K-Y5_;VGJ^9VRC16_@1AM3Ud6dHf1XaWa:E/THfR
D6L>fCIK+)EHVL8RECae(BC,V&>_M\>&FWCE&>NU,,;FW30G</dbegA02GBZYda&
CX=Ke_QdYCK;(fX<SN#Mef,WG8^(7J-U+G^g014V:g14U,aVb9DeDaHVFe+McLUV
LPZ/QHB;XG.RC^/K@\3=+0C[ZK82b<;d)K19;HcJFJR02QJ.[1FIZ0J?bY^3[g=V
,&[-Gc_Va^3e,2ZEaR9N>GV<_/EYR81F_8<&910+N.QGM6,g4XOf1;>)e7;GA@Y=
4ZVA&S?,.I5>4WD-U)6e-PPI0[BW7RAFR,I+SUK\+9a#@?F7P5#a:.FVK=0TVJ&]
8b8aLLBg[g9g.6AacD\[R[88A5VJ<8Vgd7=2WZJHG(NRGL-@9#(BJ@71KPIc>[.-
2GdU(_P>2V_>4]R.)QeRA,FC1K+;VDOB2Kddc(UBAP1c@c^A<,^4^1=3T=b:+)(F
[Yg@dfdIHVPR0)4QP-9=+5WHI//8RbRPcf/I7ZF=KX-4I7ABWK3^LU5Qg#1W7/_A
2TMe2&:([3W^:+NP]JZGS04Z-2<:BJX&5YR+EEN9U=E.X@(1WJ\RcO/3IZ39-R.+
,EO7I0J17L[IE&A38WYdEP,IM-L+fC,5B#..=,EWF<+5A4@=-a_R6YV;H+bD0_::
G+CZf8ZJJaS4?&PU4K>8LDJ^eG:F[C2#IP8M/AGHC_]CETV]V:97+bfLM(FZU_0E
K9?+>YAZbP0\ZQ#O6FD1Xc7R8(NeX(/D^_fZM4I^A)A8CJ9;E[Me8)..N5&MG?Ud
PLgQ9b<G[?.c62G.e+PDg\+cOS#)HMT_fLP_:D:#&?Daf/?EHFIU@(VXEQBf??a&
bY,[9/_IQKG9a)5]UQASE&cXOdTM@03+OY9N5>QUE,K^_TMaC&OAF3KY]BT(NM9X
4+8EPXF8(^.<SN.)#0L5/-)19RKNUBVLIV.gaU]=/NN9^PPeWa[;cg,,-:(QG948
Q^4[eQ(@<+2TIc3422A_:d(d.-+4P5g,f(]&N:3X2Kf^J:7ICF3QG,b;41]EaBed
+RU=VPQ)#H(X+2L#1D<c:5+GODFFeJ=RN_OE>f=B0cWUY,7T2ZX^8&:O8Oe#8[bW
<KE[H?/1XVV@@8ISMK=5cM\)+T1ICUb(UMH;I6J@-P_(]0cIQ,5MMQ-VX\]YXZI\
T+Z^^PG7VH1O2eMJO0YVMg?@Y0b.@=Y95bb#eUOI;.)I&+FSO[>F<DZFSL^V<)0c
FbY,)TV2#M?LJ3DeM3:YFa9;-X4<WH@EI<F_KNRB#LEF]5T2[gLMAOJdZ4ERK#=Q
W><)cVZ@63TU^D=DE>]?>W<S+CV5DQESVa@b[=U6R(La+@cIc2IWRL@8K)S:)L\M
&N)ZLFEORYX^[,^ZC@+=2I&B3>Fg23J#8N^\]IK.B7bDB\&:X5UBE6LG-HI_EP_1
_1&6?Y^L2;=6E7::77@P)[[T^BWF+ZJZ=#)DPHPdX\?VgD\TgSWc5dN[XR;bN8#J
(V.Q4;QI?F<X=&4c)0Z+=d[\Hb[;ZR)_16)0SIaY)LdE,@GX+VeaE6b0@C9UOA+)
\8@8H#bZD6#-\,6g]\</H1F#^/FG0d[VB>?e-^->Rg#4@ceITM<A:OF.;7X6bXN/
R#4\f)0?-;cST#aO6eP4.^7IXM4XE>/JG8[>0bPMV+f?4HNM:Rf&Hb2#8A#@gNA9
A3+eF7TO7S9,P@Sa86+@fg8g\#2]:M0Nc<5WEX]-6dNU)E.YROCT,D=D5+^Zg_;C
[JCNOE2D)?b0E;Bg5OFH?1<IU2]dQ>L3-Z>8GS/gU:2_TIOG4eI,LKacY>^gd8Fb
c;M]V@>=g5FEO_M[T\N9D]?^>_H,K6e?3bO?0L1\NLGZcJb/OPQ/fbb#dI\O>6f,
=O@.I#IX_OSB>K>P^b[4QL[#?H;GC8/>F&C:A+g09O1H4?2)eZPB08dGH&YUQRd\
JDG6LRRec-DO[9be0T6/OP.;bS8>:?f/1c\KRPIRF)+B]9_U;KWZXS5VZe]Q#3Zd
b3HKB#-.CH@Y5Q=YRQ]NO)<P.aZ<^]#+.#JY>)+5f])Ree4.[Yc>L>8+Y@cHOFM/
;?B>W2[71X[K8b6MGLF54GWE>QZACM7@0LX[0)7G4MTdVb-&5#8@8GF;V/DaJe-@
_DES=74?67a:Z_QB<0K.I:Tf0V78_]5MY_O3K,?:8a?Rf)7KZ>5D43Nf1ddJVbVL
VGQ5WO;.L9FFGK;I?KfR98:a^[N91&c)&1IQI,3.JT6aXBOWe)8>&O0I-b@#?6#>
f_6]/eL<F7P4T0ISNf^3a&=0I2R?cS\NGC.-;>WFV.^d_B8V;=/O<3V3\=4TN__C
5.\[b=/PW4M6-8NHU--[ZCJ_R1;.SVGd3.QD1/26:F1OA_#):-bf/>:7&Gf_SENe
dQ5c<IRCD3SA&_]_IER6#f=1.S9V--fD;KG+26:\C^Ca0YQN@QR]ZRY)^XJY]f)8
G)G#\?LUH>TR3F5YJ,UJXe^]74bCI?Q34->_DF?ZF(A_,e.C2=:OVB3I/GFa5OL=
V^G3C43L9gT34-R1P4#.6VIKKXe[,&1,;UK4=1FM],4=DCLHgU0.+P1R^IUT1A#+
JWH6W]BRC,ZECT?QccG(?LLY:DY19#(I[\&6)R6.Q[3Y:TUc[;1MLSAKA[B_gKAg
?/G_LXEWU7T9\Q6^KLDYXOe+ZR^R(6)M[YJT.2/aL6=-/A(4CHGIbP\\]1W<@(2L
QQ9_U^@>B0;;__14J3;f7T(e:#O/7P7V17G6=VIQVd@P8>-B;/V_Y,^3,#&US2c.
<3J05K@7.aY4RgJ&d/EedDTR(X35;E9W)G]N.TAMIK\VD)Z#BNMKBL0]1T938RNb
^LWBD0QY96#Q@MPWJ:d#:=C<&,f@7ZKfS(^XH)HDdN\-J]->04/.4[:,@eR@IUe:
bYBK7eMR#8PSHbC5E@<(UWb1@R0[JD1X2a;)2M87TP6>P.?Z&GTP@^_Y(/X:a5)0
2@gCAId08P?I1/0>>:-A(O7\=S]dF_4.1?,FE@>CW&,A.8K?Y_[dL.<JUV)OQHGT
YW^Y,;<35WL<48R(CeC_A7-_#+2TQ5+8(f9=1O#b2)RRVVf[0(6=HUKa;);g4f7b
db8I5WWY>O(>0L;YFXW8bAd3R3G.5.3_/A3XE]E+4]=.MU,X@C[D)c1OS</=]VCE
c#]@T&4I+^4=R47e8(;O]EKNd4)UAV(f^C-B2cP_L4.MEIZcZg0O6UbgD\?E5?=H
77@E,3@gNSL2X:79#PANW5X.K>\8bY7F-A26[H0.JB&1DT>C>D)G3)F9Ff8_GF.C
F-T,OPad:6_(aW+U.:.2@aI@MM99KT2LfH&g8b=]Y]R?W@e2aO.C/&2<_#RLI+_S
d=FcOELN0eR6R?YM:8W9-,8HgHMN,FY];+7c]+7cVf--L33eG82=P&F/?cTJaCE9
7MdgWR@NcT6&H4E.JVfOWBZ.8Uf:B(>dF?LA;7\)a\g>_RF6a<FU2H7A\C34Q(K7
.+4S8QA_M(?LcEC;G&<WZP(//.L.0(ecMDc<dG(c(TaII:Egag09?#_E)g>+35/E
\9.I0NWS5@]c3+)JLOMG8##RI>.PH)RS\P46fN7cN5a=AOAecQ11MU@RJTWP1PVO
216ReHKK(Mg&SXK8RGJ.^3Z]W>a0>8W&>&7QcCT-IFL_1B=ag^fLI?;fHDGXIA)Y
Te:P;Zg,fPMf<3N/,8UefWFggXe6Jbd/XNf8467M+-1F?PA,QaKA98dGT/c<5a2e
E]\Yb44.<OP&PdI3CI.@fe:JSG&Q4EM>RG&IM:@)L&Sg_Cd^T:4NKcTI93f.-X#E
b/>Qb(XFG8+NG5Z&cf3cOUR-C.W.-@CMVc<+798F1^6;7JU&eV:52a<J8AJP5gQ8
d+3+,;A@>DI6-]X<ga5GdR0(0GV+cI_O6Q5DM;KKAe2YP(W]-]#]0S3;ABP&V@M:
JH;1[460H.A8b3]L]-35X38fd(Q.]9L#/+aE]1&^FNV#?f)(Q)?QVJBGIG7aFDQF
P1(@>bP.db8&OeUIFXeM:&?:BTf=3_JD&bgaB>9#=V=UHEOCgf0)::\S7IIH\1@:
W(\Z..851@@>gS:-L@SRLa3<A(dGJ50>.ECI#c^LKM.,_DJ0N@+<YCRAE/b/H;5&
</-X6PTQ7]K)@Y8YSV-5Q3[NaV:gB)I0BR&@<YBN[RIS7-&1aN_I\6#dK6E[?)EN
M.9)c)COM,LM\PL8(JO_)()IR,c#P909Y6@O+g/7M5<@Ae>/g-)S?U;6W^0.S0,U
eDDCfS>SUK9S20GO9bS7W+OKD6<:?Pg^<6DUQXVN@#.KIJO@>@>dIW#P0HKLW1O4
;WI6d==+FA4NS^2P-H<Z7=B-@(EX3f;:IS<^X48I5cS.,&-3BWWNBJO2b;]17W_U
]475Qf2@?10DYWM(X90H39b[06X\H26&d)fQ;b769RT6QTDJg>7SUf7Fc.3QJL3Z
YgVc2B>c[GH#)0H\G+\:_<B^Te?#I5=U/8EFECFX5:+92=(ReB/5f)93fJ?_6d..
8F2KQ2Z8\D<,DL/NU3S<C:Y>eS[+0MWAWU&Y[,DJ&R#MBe=a<6>//e0gef-,M>F9
O35SLH2N4gNOPMU-5WA1?2G7X)eY.+R6MH.9<,-3?A@9IAP/4-2c@^Q)cOPcgSf)
3#<[ZCaHM?6>=:G5B<QDX][@Zac]XU;<AEB)0Jac]731g<SBP:AJ-XYb>]J.X451
]R5^/5[SO1PB?,]WF1S7g.+;AUAXdHdbZR^=T=\3[64Y/<edYQ4ZNa?9+X&.I2MW
CG^e##e_Z/1[72cJ69^dCHb(9baZM5D/5dGL+Q?A6(=EHQO.c>BF=ME0GX4VY8)a
?XW+84Pd4X^OM#1DA,f-,41g/K(H<c;2eM1ZHg,EB.U2YUC+?_#(0SX>&77/U^Ud
C6b9W0X\N:=S>TK2;^>(GPR^\@F>#ZIA..L<#Q?2#0?fPXNgV;574e7cc(;bS4<A
QTN4]QQ5--9F@XKf,X8241Bc6U[(0+VKGC<LF,4\CXeU];GT^+VCg8)DD)@Z6\N:
0g/\S(6>e>UIQRY&DSA.\((;\EET[2?d,RaLM4g<K\/a;YTV\\YW-gY5Qb3Ha2bL
+()gKY0X/_?O_(KF5[#[RNS,XSJ>60JK#K#KBJ7F9bM7#6PRb[c_9@]e@L06\@Qc
.J(F@YQe/Y(0gS@P3EY]7RWZG3+Hb8@.H;(FY_T+O@Q?24PgU25f/WZcX<(CB4GU
eHDGH+Ng45/fZ9d@BG2F:a(-WN_;]E,43e5ZC<+EU;,K]Dd>@:Kd8L+Q2#U8:TX\
D]&7dR,bZH9eefBN8OZFF?DSYNa1P+;eF\b2&F3P0NXH28B53eJb4Jb@39Q[K0&)
V38UJ/V[_3f?H1YVD&&X#L[-d=&+NOdUF)XRMcN?ED3PR1.Q;<G\FNE<B87)fgKE
FRFW)N0:(B+)5#74K<&J^X2,HH>NC,)-aMRAA>]0AVYH/=X4R(4;cOD&eVG.AH+W
.=I;[W3]=OH[YZ81:S>OZ=F2KaJOR+1,5bYLKf/1/-d73,R;1cDgeeUUQVKL:,PA
IXQTXLEDI4aLLe+@DB12eRWf9DafQ[/a=Kd69V)aW950e<g&X&;e+H75WX:L.)^_
GQA-51\1^:KQI1DKI7EIAeWAL6:KA1CDU?K3DgAQ;(;XMe-N&JQ[TDaCg8/<C9)>
,V+U+fQ=a;7#E>GI<1e^K[fN3_#1f]A2W>D5.JRUS>EBaU.DTNR,5P4O8GBM\8/7
)JD0(Rb-@0DJbB0<>eWeVY3:bD.H[I6eS.5LK<^fNW/;,X(/RRKQM.HW+[JE\:-R
Qg/;6d&+e0PV\BPH.75d[NGD.S_eW_b;SA(Kac.M13@cf[DMgQI?@RQ^AZMF4H5<
:e9Z\UdW^K-31HI?fB./fgA]A/G^=62OfZF^9:BYD)XWNFF[];G@11C,ZD-e2)Le
\XfR52/SN;e8[f8QYVO&?dVM;;]^U>)Q6aZD1&@/4/_g+DT^\G[cWb]P((?T].IQ
KfDK5HgL>^OB_NY?,#26YWfa)P;+>TDH4X&.JI5P8<YeEB6WM1]#\gdQCD<YSPPF
R[KKK]ZFLI[e>3F1R/LGa1.eQT65#d_T+QC9D4OB2YPKL+)YXTgd4IZB>,Gb:LcL
#;J0a82]K2>NLPGBNU/dbL\@/fJf&C1?HSW2gDJQA:38=05]@]VUf0H/Vb>e#6cK
4Kc@f#Q2RW=X^g0>g_7JacbV=J7]YgX/UVX9Xd>6?5&Z&>.bX(>g<,HR=EUAQ[aN
B-Rgg>7<3Wa(J:7:4RZ21ZCT96JP_3&&/@TY3=YdX)FW#Qd4A#3);XQ-SY9D:+/\
J5W?+UG3g[]&2X4,&C9+@Qb(#LdR.4ZT=9056G)D@<D<-_?532\7L=;7fG]-:aDF
C-R3#YO\Gb@7UHC_PVHF2DN(WQGTK\R>5T8f+4c.J3F2TM1b.a+5OBQeX#U#@WbO
EY.22E-OLQI(CCLII-_L-/VOV7^Y7B9Fc(cbA4W@\fDd-S:,#42X#T@#dBC;L7_H
V1MPFSQNLMbAc\3SafNXDO1_>78g/Pc942+Rd@LA[\(M&(9).P3XWV6(Q/(#L)[1
CVVT7V7)c&7WWHR@O9dI&3SV.RbJU#^IK/<L\459Ud,CT-XA[O<BR_YO@N65;dO1
I;(MV6g:K;H7&=1?T_(EAdR;K=&R-Je_[UL;SUC8faB+8#[4O&]f<5EQS?IRg13W
[cX=^,O:B(2Y780DGa[-J.DO-<EF<M,Z=]K3^T5:GED8Z=]_eIHN>_T;PD8\Y/N\
?PU[@][O8<W.Aa6(\67H]2A)N_D)8Rba;.#)V<2b]cE+c,[55:J^04a]bfL9H]Xg
BgUf81BOY,bSca/?4b\&W8)TU4JcQH4CdH9aJdg5:#@+]]S?a[_/TAYM/H[2g,:1
e11Y;>O#F2^-8<NeZbe1XdFI.N/(W/URg,JE&D+?S[Q,c@(I(BPK)AKfd+MZGPS7
>RPBCZP-X:H:-P[D@)eZ/0Deb=7AdCSdJ9VLE3OEWJc(#+[?XNa\6LbX9U0FO56R
&aJTH;TS1d;Q0E<)bJH^618bgGHE[b03G1Q;1KOQ:B=A2#fJL;1O>9O>.7P:3-(L
ZfAA;fReI=ZJIRS^UK>(H>cL>&MT+AI&^+b4Y[;;]6?1XM6HRA2T_b6g,C2DR)gQ
Ca03GI^-f]A:WEHOKgOO;+,1KfDL1bYB>JTJXR==#)Z5H]Zbf]JQ&EUI^R[Da\KO
I\;)HG7Ne;(F+?VNaU<A?Pf-Yd>>TXF]?-:G7)0:7;6RH6=_<W5B4;Zd@.)]fgCU
cKV+a55L/+-J@6A#=^Qe457_\OH#c^8D22c\@LOSYADdS>6Q)WB&079XJ4S1?/dQ
KcVf_N[C0DUJE:>eB?B<dOW7K8H]V@Q9dAMX#<5PJOXI,L8-f5_2?APA;E(FY[;(
AX=dVY/cZ6_#QZ<_[:ROZ+1fa#(]02Y)cG)HQa2aEVZVbA8UaJJO(>>4IA55DgE/
V9-T^#?U7A+dHeLRG>1VAg:(IFPL&g[88&fFI1;R8W,+65R4;VMR<_SE,3C&UG;@
7ELTf-CR<4242E3.^@9,+7HGb0X7R?_a.aFK?FM)IKKB<LA[LC#^[M(>_.Cf:N2+
TRaMG8C6c6C:3,TGN@Z<\E::X5J77Y/IGT[J-Tg8UbPFd?HA_95>Y;fWB3-FU+C#
b(?8U0)KUU3M]OM^LT(bCRTR-0dR-]Zg<,JR((635E=f\[gHC[9^?+0E&Yb?9HI\
/1b5O>HV:eT(M5_ZaAeYS\eeU_J^F?3==NaY.f6M3U<fA&6I4_d=..7=IHY48)D]
D-J_dZSJb,,&DGe1^]7X&aZZ7&X5a=2XHeDfK3PGKH3--4KR7g6AQUGK-=IR:e::
]b+CZ\U6?g/]A)>.6(Q3)3/@f55;VD0L8Q;dbN5GXYb3XM@^<=(_L-AE(,[:?C)3
F;(5#L?\5J@^\-80ae#NY]LPd1ZOJ@8_:<M1OP[N?Z1X:Wg49Wc-Y]EAJB+;ed)(
P)75ebD,\S/5d8#YA+124#ZX2-BCNYVALYMa3>)VLH)3^^17cS[-27UM2aZ=5cP)
VBA2:]J,fb-VX[0^@X>F-6JSK(6DUTCEI2>6DHXDVAWP):_ef8E17MPEb&@O2bE#
Saf7&XL]/U9M9&CT>B70BRbJ4HS]4XIZ>G3V8KICZ0,HZMOJ2^H^\WSR(d3PHU;B
Z<HB_<_b\4?\A\A)XR>FNc#&_&?YBcA-R\I3gYb6LES,c,V.S?/+gB9_LgE_(13\
J#U,a;HQ[+,9#+&3+7:XO8/O4X2>bOfE@&?VSeeZ:6,<>,Pg&.-I];#+efV5E[Hf
-R#O1[MUJ_8O9fgHc>:F)5?gN1CO)RfaPZa&8X.^f:T63&>Q0FUAW2(CK>6[b1cS
b6B.7XaF=7S]8.7c3ZW1?H5aWF&S81.LL)daAd.)1J==aA0Y:4U09ccJP@dPNdB1
=52&\.?M&J>(bEZWg^8U3.bJSa1ZWScV?.)SML;WD.e]gQee5Kg?1+SVTG5M[WF_
\?YBW^A6PGXT0+ULO^<PU#6g44_203V6L,:2/+=)(30ac2=?2(T[>eIGHbD2Y;B=
gDK9=eb+d#)>7-CQ:YgebP/V-R1O<XIAGPTX7UICJ;,f-F]a@9Sgf9-&BHg]Q-GB
[\.5-M3+B18>2aDHR0H5<QXZI1TQW#+:K8;9+E&\;Za_QU0&=,O&+(7L)&Rd]_TV
^D08[2DBJZcK/cg;fH9.N#<:fW&KYXHT?_b:6/?>fHX,Q4I;&(Xc/_LTCa:>\HbY
2]Fc:1;X+;TaLCL<.HOEg)^_7^L-Q0gEH43FM;P>10T2SMFHG&:HB1D8V>aGafF(
T(]H0N@I#I;La/Sa6U9K8f^NSVNgXKCb)<@>TZNG(IP^&6+A1D3Yf5DZd\?Qf7GX
L6N682fa-OM=d_2B36,0ea_O[f?d4WT+]?[&5>A1Sd1EII8b^W6=1Y5#9<]FF57O
X07:e6CQ#d_Wd#7gg;;J[\JaEV=&S1]gcO+(\D)S/+I0+gN2gS?RET?+aX22fZM?
&U>?J^J0O/\UAB-78(MR=-1R+8N3MDXb\80R[\==W1^(JBcNQ\CCNP7<M>2F.gg\
3,5J,#aG=3L3)PeU4L?OXSC/-K7@_Q513gO<3M<N,IZ+7/_ID/Z:4,<PA#GE+L71
AFI1NeUeUVIDb1+.4GSC-QL;M30=D31:K+<?QKJB4@UQ)_E;FbBC;gL<7&V559M[
--F&a#29<gLbD=e4\0G_WR#0#H#(#:U40J(8a)d_78Y6WJ:cW/RP_[ce-F]7BBe^
W1EAea26M+0;K/OCb\N\#H71N7)#(Ae<NVJ6KXOC2A1M(F[IJ+JZ68KB.Y5P9H6A
)M]AO)c[=CW-(1DK\]JC&IAYX/R+,EH1Hb<5?0D)^T67.-LU4W]BM@LA8R]c4NQe
HQGPUb8=_+^7Ic,H<b)PTeV:M7UL(]#<f,F7,IYSV-.D,.;bgCS)8T[/FI[?N_,C
Yd:F:18[a,X;W^c8B[#1&PY9BRe567465JAS2.(9G2(Z0?#X@V:fb7:bO(XB.R=M
,C:E>J@:&RJJ;C4Q<@[DY<AS74J:gN,U0GdfOJ&CY>9/+E)-N[E>0Q4IOC^KfXNg
H9;0P;88?]3V>5EZ+:5D>^g5fTXF1bP_3OMQVfIH\VZE7(/DA)61<)98):Z)PFZY
H-R)/J#4[cc&C@&KP_K+>cgR8KdFD<=47/5SX)>^F\;66[b_[CaB@ZNI0UDNBEZF
H#7S0]0M=3IJ31&@PgN&Q>0G:P2F\[@+IfZ?D(X@Oc?^L<R4O?M^\G]d_7JXW2D(
WATDVU0d>bA5<740O9RN2d+e=>^(Y+_BTeb3W/;=+/gc6=HNJ]/F^Y_7I:)B_1d-
&QJN\\eIWDG:S&bGca7Q4S9_b040d_R<(6NRf9UXVM8@g;F1-R/J;fD[/9KeFgMF
Y@]+/1A5^c&HMYc^UQLcefG]?DC[?:gZcIFQ4Fc@3Td,SS^MZJJFYE:\K.^4]a:a
N)b#?@UN];f-;?[58#JKTg/FCb9ZUCB^T7XY#abQD#9R+ZNd.Ae3(eMN_-=Bc-56
g<;O;PU@EUD_#>[R<@G&JE<LV[bd4GA,UK,5IB-QB2\YPfc_1@M0;5TR#L/aMgQ;
,K&]\&dcAG5d6HMDXH<_CAWPH=>If-Da[.@#WFDb)B/0YJ86CYSRGK(YE\\G208C
3F3:JFO@E8d7eM;9F8Gf?,H\BOTfd<2I2QBF54L3SG/K7=]6)7I_(5CIYBGUFJAc
ARY<NY)J&VgHZUa)&LS([V4?KR>BM#R;0E2/eC<+dSS5^GH\\9Zc[4#[E.^2O5;U
HaFFc2WP=GO74,(5PH1g8;[9:F,U8N?VaE(9L.MK[G:WUWI\9Cbdb[8f2_>[LbV3
?Z/1KeO:bO&XM\4c4W#)7K8CS6c=9VG]?.eL.8B+bH@:SW=L/:F3=;F)2gRUC7ZU
V<VdVE(B)_/?CDWO)dI@Fg&cAIPCZU:eL[@#b8L3.,JRW<=C^OZ3dZQP?MT8^?XG
?CL05f]OH=8QI@Pc>5(H>VbL<5)Af0d=9T6R^VgH](gPe8g<)Z7F6UL>;^VSf=L/
@X=D0SEW9Y;C77HM-g\IG@,H@X.RY)\YdS_B69G0ea#0#;DMU6/>@HK?+>[1HC#a
4TP[K?-YD.]d=VV1eg7UJ@EWO#@d:NIbeZL,&P.]2T:KSNffK;X[cMQZ37+fH+,/
]f+,XI.U08/[f#791K?4:K8B^IG03+Hf&/[QNJ>G0D#P<);bUO9P&Q>EE.Q_&g/I
,_6@RKd8([YS9]0V6-)Sc/(D.9MA44QC:\LN708ID(GGf8R5\N6^,L4e-;EbB^1K
#TSeQ(E.:DW8.V5/K&&V,IcL/\U6g0gT&Z6NK5cPO/cVeO:#T]P97dWGEVVGS:1(
A&3A4IRXa0TV@KTJ&=;?3RHOaK7NVSH62<66ND:EY?,N5d,,2NCWbY-Vd<=GG.<_
09>.HEG(YOC2MVS(Ug6G<T?.;)>Y(SH<CHa8=I,W62cUX?b-@28E#[9H&7g.7bf;
+5OZ&DdC(WO]@N7=,+/:[01G&a\R?=H6F:45HUSE&0.FC;[,)GNRdMGLHP1CR<b3
We.5YH+,CK3<#?QF.A>7(P4U3_H016cG+\]:cU(=?3(8)LY\R>Hce35D8ER_0-K7
Q[8]-+-O/(EX8\J&N;GJR<(6T)\adBT09@>3FK@Kb15048QgFB;U(NK1O1>TN?=4
=gBB/D?=2f)K5VN(MGGe9M4Q__@GGaN7Z23b55[B?F.MP,.(=OdL+Jfcd8UJLNbG
THL>YTH1bK/Jf2P4aOT_F:U/\<XB@.2ILTeJbH=@75VNERX96)/&+1VHB=TVT^/(
_@)bO^9E76]d(O5Pf89BfUO1@K>5KT3)aL)aNYJeL)V+&.T><GOUEB[;17+f,ZRE
fBQPU)YQ_F+)JELbZ38/D^Z;:f&=^C9<<CJ=12P,LEbT<#OG\8B7:d5Pa9HaX<R8
87c;R2H3FB56DV-=32F09NE8dL(8IP,@O75gXM0ELaZ;/;-6#g)18#_@SNK/#_P4
:&X.Y8TgTRE/:)-1da@YaBB1=1D(]@OCS.dd4S&&fJeMPUe<NML/]K<A\ZCgg:-T
&UD<V_L\FE=1Q9S6G@4[(IM,Z\(_+9YXSP?&Q?2E\C9V]U^JQV9R/L@ccPD:8bXb
FVFU)XV:QODV\BK&O,eaM@79)#6M6M/B:3RUN-ZAX.6KM95?YW8),ed[Y)B2<DM4
7Q7@H>T&EOH,Fe_##eGJC3c4W3+4eIWFMeID8A/VW0.-/ELcXM<&P,Jd5H8M::L-
IK)+@=T_T]7DBb<[6C6@X^SF=OCQ?=6DL4[[0edR2RW4,\V\8OL=^)-7.0fM=+-+
LS6D<2^FbWQXXP/9<4[ffbMI;()^@0Ha2]cL_)-W4Kf;F9=+QaHS#Y=LXR-X@.B&
e9C71S)3+<.PDRe?Pd-B7C^QW59O[c&QG#;YfTMg8P^Z[&#XA[,eMVDSeV/65MCb
:^48^OGT=K.MSB1FfF;E7[,BWP5U6M01A8(3\d9GPE(EU6UCVTL6b25B)&.S05J?
T/P0P>96^Jb,KN?Y0)GFfAXdQK,,Z42-S?EJ&9#^@>V?BN]K4M+(9^UDD>?A&e4N
CWc.[3XHKQ(2;6>]]8<_L@?E?U)[g[?BW)1-Y2&/9FF4#-_QZ-fba/T<ZZb.cJ;N
XXbKYQ6:1Q[&ZbWf(N[b_ZOUVFNdI7HW;M=PT_d)@S:RMc:2]?M1N1SP9-bG][RD
,/1D^2GVa=dUfV4\UESfHgEOOT=a1,eRH5W1GTR?A]BbQ_^OEeXH?eJG\+B&4P1?
gK>CVX4fLa,e=M];bWG32I.Z;(P=(Y6W4ZE<(_G_YUGb>,1DE-XV1Q=,_7.P+OXe
1A&RK3(=3\&&Kfa52D]@C&FL4C+2T+;8Fab>?WX&>Nc=V6YXXC0<))I1B8?Zc>T@
:P5[L3@g4_HK;dYQ5B?8Y)I@^d?.L5DL6:RTf3Ca1I]HS4C0Y_4_Q@bLE4GV\M/H
,6Nf;<.1c8,DXZ#TM2WFU7]AE/A;3;aK6\f[X\,ce_aDI>f(XTaH7Z[9;GY7#PTg
L#[OC:FgIGW(2.0eRZ>T]]Z(fa<?PJV^5Fd#XM=bBE_[J&JX@[PgIa3.cWE3A&N7
I.VbQMSR#1f6NNdF?CSQ0>JNL_IGE?Da=FA;ZIP53f?.FFJF6\<VcLER=2XF2.D^
6cI]4Scd^eI5M)5d,R8?8(65<<GO4BR^38(2M(&Nd3@;X-:^S[3+eHcd))G1+Y3F
5OaU8TJJ_3Y()LeFg<Q+Z^1?\#WcQ\fH(QLVX;G2),bAL3<K&J;#_+<3>=M4BA7a
UbY;HV6KH7)D+^VML<X=L?J[Q(_U09FX09Y1>^+\=OOd1EGSW=3gSY2D(a7\>F=R
Y)<XF4&]_SE20XKZO)f>_7/=dEG+?34PUB,IRa7U=/[JbJ(.8fe86]<9fecfcU9.
Caa]Z#K#\NgcH9YF+9c5O>a;0]f,f[DY3QbWM]6)@)(L[JX8>SHcIGgSC(^HFA8c
84FAD5X:D]ZfbCPd(.SeB?S2)K.bVeEMJP]e;T9Ad=O)USH\W]g<F^bQ)L:/1,-6
9K>H66<N3N5HZ;3B1_-+QK+MeJEN5RQYTI0W74ePa1,3_Ha.XB?LLRF4bc1>SJUP
&&@&JbCD]PgB+]:RP2I08KCN->XNgF0+ZSC;1+(/b_c9M,,Q]&SQ7a5K-a?<,>8g
P#)W?6&8-DNE6\S)PXNI02@W8D9SW1S^^>PXL9?A@ZEe1I0[a^c-C,7(+C5W85&b
]:#Fdf^5?AbWZg2Y;UcUU.M#-b0.2GL_=W70)]6DJee9SU1\?baOIHCd,[UU;3YU
F98U6N?0,L;=@Ic)@W68J#FUG,4LC@[;(cWX;<0b>bFe7DJIP)eV8#f#8P=bQD\C
H7;BBUc7#6?W>CO.ER_GFNd_BJ?H^DTEEE4=C38+5Xa9SGgYCQ:JJGBM<GL242=O
K/g9WZ7G^UbLYUd(b\P&7ON#EBHLOM1Ka)b_GLFAL95Q;1+GaJabQ]?Za13F5AL@
CI)-A09f.9EIcM@7E:/40fG^ZUb4QNGI0cNQgA:WKQZ9.=&eD^+[<[ZE:A]-,>S@
-W[,HV#7J?V\4a50_4U^,;a]?D:<<B)KT6)0=gMRcZ#CGLI<d4+#K]e=Ufe^bVD@
\Yf?e2JW@KZ3IULaDM>(b6)cPQc(YA\NfL8Rcd6Y+>=:Q]<K7DE@Z=6MZBae_SV2
1M#,d&D8?H,Y4TJCIKK=4ZVH<XB0PRW@E)=cY;+DF7J][2>(c[gNE2&9@/2b[@0Q
Kg.>:&#E&@<<J;MP[FC^CPVP?7E>I?-T#73\dY,e46&EY62M#9M1JcDLMUMQIcXP
A^#<-=WCb,<.SQ47)0-M,@@2_N(b5#R_,9JdT@UNF#6&YRN4/EUNDcV(OdbO(L^T
^<egc<9)K#fV\&H,>QIJCGO)O&feO76-TBOK31/<^g,1)W@4)YSBTJXa5PaY:USa
^:MJ:a;/dOU9&b2d-HegfgF?MILVG<&L,_U^Je7#UcHD8[#=HL#&/(PEA.<2U2f2
D,P]3NMFFFQQg9OW5S=/8;D\)d()=4L#HS/_93K67(O6_O_WTGI04OdH<KI8#dfD
9]+>J&?E7APg&=\8(XaZT/]O.?+UfQ:b:Ib(C;6U/OIFXRU@M#7Bg8Aa_6DD].,T
8G(7X;#WZ5Y6H4Wg=+<B:fJ@CQH(Mb^;WAG2eLPES0T_bcMc94b#OZdO[NafQRNL
feJ4DVNe+QUD:(P24AeX]9,ISAAP0M553-W\XVV2@HDK_YW,A8>:Za8GW0cZTbbO
R+NQM;49[X>MRQ>.WSCW\SZB_H2NVW]>d=_,e3#O]I:Z<>?O)WT-.N)HVfbK<+0^
4U:3KYOUgD<IYD[D^3F(/CRIJ#MFD#AQJeF&aU597Sf+?]J(ULZ?<g&@+IPV6[6-
0+RK=4K[QCaO,@Q&8(5<Rf;INQ00^XQ;=R_XN+H-K5QWcbB,<(a+GE6cT/L&F?=&
^AES#d756O6aWMa01(9V3,bH35X9XZYA419S4MC0_O7734R<N_74@0EaFJD3\g^F
6AQ,_+48+#4#WS4NCQ.)4G3:]R#\9C8fB[YK4Sf23O6WgaSUW_QR2DO&D.AG2H[0
)ZFZ4>_H#5VUXM6R]C\?(]4g_c.a6d,,G4HGC[>U?5MVJZTBXf1-7LZS][f05/eF
-dDF)+^aO&K;/AO41M9BV^T_<N(g\>84^5<]5S2&B0/GK>>:PZ05?5);KJT-2I<g
:[IZ=,&\.L,H_cSN@,L#5Y<Z#b8OQH-RCd14Sg\C@;WU:>L/;:?H<@3<ZTM^U6V8
N7A2P9-Lg<c?,_0:=]5&?]0bc52a/-fTY^=LI8cR1Y:_DL_<G?^E)^FLOZ?-D=Xc
A@B166H8;<g0]RK-V7OGT9L,I1-aVDIK7D:+NN\7c=5d_:\&X&>I6QcI^A&D1&,4
]#(T\TcY>2^2NQ(WMVD)aaP,A8faagc\a/9OFdXLV@)Hg8RTF=H207XcA6[VA<;a
K.XF=KF-.IW]J=VB:.?HZ5[aWBK:D@F]?+>?MK2@gVR_K)+I<(.)DWMD)2?42QEf
:K+KF19?JO>CBD?(fEO5(TF^CTfIg2,^^9bg+:L/>5F7dSW724TT&V^AETHJ<K3a
IVD/+G],A;DJ+gF).V]/DM?PP2:A?-<)Ee_<dHM>]#,LPc)<&3=/I]DN(QAdU_Z9
D.d:VW2B1CU:MG6+1(K[BG9aWa?,IeX.NA\&K^#ZT\#8bKB<RE2XSZ[JH9+[#KE(
,7B95QEHSK)-1B0084:ePB(487M#GY9Q:$
`endprotected

`endif //  `ifndef GUARD_SVT_AXI_SLAVE_COMMON_SV
