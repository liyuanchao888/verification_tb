
`ifndef GUARD_SVT_AHB_ARBITER_COMMON_SV
`define GUARD_SVT_AHB_ARBITER_COMMON_SV

`include "svt_ahb_defines.svi"

             
typedef class svt_ahb_arbiter;
typedef class svt_ahb_bus_env;


//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
N6JU20VRsFxe+lBQrPnFbgum3MoaHNMi+CAQhIHEmricOk3uXh9ByHV5Ti93Iqm/
o7DrWOCN3owJNDXPFtKSUUe8/Wg7P0T5zUnyiWVjK0ennzV5s+6MfKwNZvoXPe1z
Ka6OxogDR/gqYu+YcwfxHhdIPqsp8b4BmBf9GFfdiVVyA2xcQXuRRA==
//pragma protect end_key_block
//pragma protect digest_block
aEbVxbQBhyFcMhOu+eLF0CCwa4c=
//pragma protect end_digest_block
//pragma protect data_block
0DQA0F12Lgb14ETL9eUMOlnWRcYbNIpxnPWbD3WD3PPiIUEvOdT4KhI9D7c5qmqD
HUc3ee9QaEEo8KS07AHj6EjXoqQD8xM72t5CNoRpoQ0gDtqy+pO5EqoMurZHkotB
XqBk7CyOutQt7RUS458Rg1Er+JXxkadLalBp4+B63ITpodx+p7SYQHCj9iWnC5wl
mn495DrNMu3to1Sxg7iA5Vwc+pWAbT2Wi72MC/f48uP65dG5ZB/IefOEtMxyuqut
vJJhd3UmmGA5/+QpxI4/sAYFc12+SOAjWNZgN+QR+rrjkpZxLjTSiN55Y8g3HVbv
fkxurGyErZUS94aUl1O9cqqL7FEXoGc+gFRbP0xZsn+NRoqwkh2JnyuDlM8O3rNb
y/Y5WFdKdy8i0T0i3KODUblEgYdzsTpTZX7xBaJ6DzjThxeZGwINNQx03iKDio4Q
/regznSrStivKtZNcPP+yf8HIMJ1eV1owwAPA/NtWDfMbZDLPTC/Z57dFP/AuDLk
grcY0BjfOpvR7qJLvyEC08OHuPZgaWcgyJq17TQtLlqj3hCyHDPMSEUvKLB73eCe
47ZcSqEvYbFoEpe5zqgYnJwn5rQf0tcS7KdtRoW4PoppOX5u4qsLjH5XJGrV2waD
tP7VXhA977Po0iPFEf0BKve0AKvpf6oavGB/wtsV+0R4n6hOkUIbl/IzRG+cK0zf
kkWoJItCXFW3wfuucJ1Ck3cHkoLBJhpkMQMVF0VWHA4gytnzOIxEV8YTu2Yq0xhM
jd6Uphq3QFzRapc7ohdidf4XlhwTV4BN8YBRpzQyztQBZ6Z8hYSqi8ggYV1t+0vx
QqgOKTwouzQPVh307BHBmaTTjUrWoYLsu2c88QBS7UwlVW1D6GNrRkRhI+G/Gbm9
g2ZJxEHRRC1i2bpWXP8L6mBEMBveJh9/8E8lDOgNSMn2tp8PJfhib/Poy9pBDrtN
mFdpKbi5+MsX5snH0CFz+8cMM+UDmQCgnijeShsCme9H67MJqdhiYb3hLaWAqwr6
o5084etlnzcqEmY10lbK7/rlH+qLT5eQoV1XAyluCqhwpo1qxkOAF2nt+4+EBPZR
rtEDWq+lv+VE5iZOrCS0pAUrJkBJeONFLxMFBQ3siH6TGibOge4XUE/jAj3iNQh5
xOTXHZJTocoHrxu6cuMPlw06tVy9x2D9bGenN/B0r6Wy3hqcxWrGxoYiCeIyzq76
XiGxEwUm4eJGOvxWzm1ysSrPi0VTwt/CaHy2PFyLffh/nFyE62y799ZzE1lFtX4v
k87m/fONCLBjs3fTkdO2NpizlLy35quFslfaANw7YoPT6TuC2TqYWDb7u8EQ3iRH
vQUqz5xtdkTlJnxvElK4NzqXCvQheBM1loa5Cq2PIn60OgDEkP2CQSBqbb0OE9i9
VibdRs/8e0OM19h+HVbsXTZuL2Fh26Z7UM/nRyBgMmIBbJFXjQ1yUvc3ljI4TXss
F08Oz4K3FGcbREC7vvKbHwc5wx6rSJLdzWKsl/aEIF1hLdX8cIO5PkaHW7VXNTdd
yHcflqQXl6ojeQG2VUi2F39MkCBUyI1alOEWxn5yJYgpHdm5H85zcPBdw6vVK8AR
dFsFSXUOl6ecXqy1Xcb01f//e+iqoSHH++Hv30DhQPexNg79BTmaoS0PN4lkSIO6
iK4T8gRaQpjvr6SUkQsHHXof6iDmVmJRch09HUoaeynVlHTx0qX4W0sHjI3FWV3g
F+fabPUD8ggjwMt+lun35E5IiJi6e6RAO9tgiUkgkXAAXddztv0U3cNNI7yIstPN
Nlqzc6iwWYtVWevoS6YZ/xojrRK616UyKY7LJ/mEr/kmAy9vEBBg83+JcLd5rzXE
522atMaF+yJ+zDUFLMK1O1PEXrGxVXoKv0SfmrsSLFOjGES/grDh/WwKp+vJ3PeA
3Je3fK5Z9emN3osBfJ/dooNeUBDGWv9C6mfKdHorXHyUddm5OeU9JcVO3h0RkDCm
HfT4Pb08kNkazRwxEjbjQMEG7Z9Nw6rfMt4qIUQ00J129R1ZpvYlTCln5/9FR1Hx
wTLyDlNqcVr+y9Md8bdY872xkO2ooAUYYQw8XewONkUwN1qustTSMk7AMtCGsUs5
NnD3sQrVPSeVQWXMInyNrnaj4yi8afPJi2pjFleMrWEPFMs9jxVLPI/yX/f00s4l
CtcOBTRG4svLxSXdf1ZINFWRzPTxd8lGol42E3gVqGfWJjO8kHubEuF1Nglk28ZV
YyRwyJxqRAtfj3CDojTOoCP+mNS9FL9yeWnDjAtiecnclx8J9WX183HhU5RDbrRc
ynO4lXGDLzmmoqPIUgPxFTDrDhynvqbVMWsHrfT6pVxQKYYmQNyCk66tjbcLw/Iw
6nWl/BD2IEN38bKiID+7zps+aYV0khyUVcoP+4wYpe0V+p7A6/eDWS/H4lzTh/8x
+1Fx4+Am57Azfs7H994cPqaouXw2hhUv+hSHfhkP2iQ0v4H8umCP4sxT9JiGnVnp
X97Ow9VFFrzlTcIlu331/SBn1kl/2vVqjLvusjWAxAJD3BsZL3JrL2d9rxWG/wTe
HfJUfEQ+hLn1o7giNvxrVT4o4kA/05FwYnA4otJ4w3QNlQCN33tDcQeBY1nMMlMa
I2pmxlr42x1t4o2sYLk9P+2eykXlIkeKOoaPD7sXkKGzhrvYcRfgktTeR/yQ6zmA
vjGyxCn7xeuDY396nfmgr03UQVTvaERZLOT7c3f+fYIx+1zJLcm/7RTqz4tQQlFt
DfuMwdyCEVdZzrAIjHl/699n+mpn9raYdLm9aYJjdtVVJb86+VMhdh4UALHMA0Zw
yP7UD4ezMN7OlUghXQN9HxB+AyHaGUBXeOxNfKSqnkXwiJer0gqHeIFK5sOEyWzO
d9rBT0wOWaQyJv0x1GTfQOdkIRUyZPeB8V8ZbldYlQxEVyWcLKLsEz/r2P/qONzV
DjY58D39xRO6zgqAM52oHQ3c7tINSkKc9+xg85loG3bTBzwLNdUqmmpRz+4y3GbZ
GuN1gxkonVMzCbwUh4bLfkZ9wJC1S9phq+EKfSRGZf7vVo9mXhgcPMUlUE2DMV7d
NM+lVmB4DGKTLySItLvF/RpjTfO8F4L+kJJce98WeQnaQkBJnf4TBpQgDHXRYC8S
sDkyapoZVQrRJOG5yh97BsfD8KgnjbabUG9Ypo5iJbRHQzXH7U3TzMzbefOrsClH
4fjkq41hzAQl/NBYgT0sdFeD2XfygAkot0g+ZcZAn7dShxqkJ4B8Qc//tOqgJ+i9
dEGYkXG4LkgHTXHqGDiqLPEsf3fwTicEgydGswxcP5js6BgtYQeKcmgw/mK/tsb/
IbhugFOSigi7La2wNusi1S7SI0HvMWFUuQeM3LnGIxyHH+gzBeYqwRCr6Beg97Va
KgV1myvQwiOqnwzgaf2IBuFhtwbDeARS/SgRFrqYObTy53E3AppfIdlhFd8xEpL9
SXpiSWnOSnXHRK+Ver0OQqUE51c52iPsKC34iBizGxFH+yUJzUsRpK6aJx1zaF41
W5cfo7VzDEXNKGI8fT5x1efb8L/WCVigFDAMea8lA2PFkUMgFJ4fZ1AwiSdCdqpp
2uIg43UDBLSTn/h1eifckG3wl6IeRcstExhDw6IXjVgqOOQ0Vve7AW5h6aptge2u
CnRbuu2EVsXrgn2H6wn9DF2NynzxjbRIZASCgDqMzB4wIpbMSpwrO+cHMUXbffC7
Qs5LVUoGMnxNE48Lw8V4OVWMBn241hlg6egkbVpiS2yAZYNZwpF6dFv40svJQToE
leTwTI9M4nG2405pMer2dWevCCDjzEn4GPS2HD2WlycFvMbdhvvbNWHAPsVoLasK
4GeZqG/9MS/aUPnRQLm92viEvvYQIloVTZw/x0eNZ4tgEDPREhWBqKv+Mz8Br5su
gPom7YvC452dbawply+RoRvJNf56TtK58mg1koW6HbHXuwLfHZMGQui2/hyiwDQO
XCiLTNLaiidHkHp/YLvqVWD6+XTCvwaa7FEV1sSEEJ4tacehUPIhuCrID1kJfRXX
HDNc/IfrPiu2GY6ivTlNR5DWnl2KVhAKLwRNM6mmT/X0BsYPKTY1JsB4K4S4x6vZ
+WHBE673KaOSBjiupckqCuJaIln+vK5Y2jg84IfRFmnHYkadIvTpQ70g0QGB8WaA
ncPPiWojcds7PDQIw10qd4nLsM6lHoBVNwnaXV+YgIfmhHWKzp4zWlhlf1pY7PPI
M9Rhnmk8trleYqRgoe15UgAlBd2FD/r88/NveHRqwtFHjEJDk11q63+s2lvS/PWF
0IhbJQLV0qOxaw4VxyLqAXSmL52Z9ZyQnh3IiBAeq1ce9u9i2c5EO4CEzRcH6qfF
A9WXTg9sSU4s3V1U1uTl3F5rGhN2TSuCbeAEgFJFHUu+tnsuzWrAs3SYxwpgsh8r
39EsjqUR9lrcz99mXKtQKVPCT/IMe0gI4wRC7poYbCigM9knTON5wu5fooGho0y2
Y5E/3B19e8U0M85l3CQ8S016YiwoyEM4Carz1tn9Dl4rt6OveL89JBlcl87Xb4ke
UkLjQkEDkTU8+hOwI5FpQbkv0D9t/KKmnmDFYy0dIwR4shoVdXqVtDTPLNjlCb/a
cp9SaQvUpvnFtRb7mMi3JMS1JpPZM7xQCwTyj5H2fq0DC15U78/YEHB4WS0F5CTo
NnYkZ7f8QZSXOlQKRdAWHJpsQFBU3KdzfovRHsfuo/g=
//pragma protect end_data_block
//pragma protect digest_block
icd1EOyY0cZhS82HPcU74nEAy64=
//pragma protect end_digest_block
//pragma protect end_protected

//opening this macro for dvt support
`define SVT_AHB_BUS_MON_MP_CB_SIGNAL(signal_name) \
   ahb_if_bus_mon_mp.ahb_monitor_cb.signal_name``_bus
     
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZM0jnu+duUEWj4bdCbPSCiHcDbQ4ZjdlglXKaDh4tvdFDf0QRMZdIFVABA9obsmz
AD8PK/YVhid7BLhNBgqm+4ZO6l6cY5/RHupumkrCLMkM+1Z4omHGORw2GAH/FTMA
KA4IsT1G7ZIvCd+y0Xy8LsreT7dDn+xYB1rpFTgz/m2vauV1ukD30w==
//pragma protect end_key_block
//pragma protect digest_block
oiEPLR3twjNBx0TnQdmJObOD2Qc=
//pragma protect end_digest_block
//pragma protect data_block
8E2hxIKOKz8o9IpLbNMTvXunbTJfMVN9Zyshq5n91DdPtfELv7q1vo+mUHK3da+Y
9tezoXWqHXxwaAuRa4Il4eJPT9RMOdiLv/8EDO4l2gi3aUARLSlxbCnFFQY8om/A
si4Wi3rIpXYbFH8RG2bV3C0DorP7QItpqeIO/3toe74R87g7r/VPejvP/UCUBVsl
wMsmb+xTHGYeDSIw7GZGKrjjQSeGwzXI0nkuEElxwXS6AicgRUQ+/wSW0DT1gZDf
cUcvBWa4ubeVWMD23g11zD/Bnjr8nim+XNOq0S+erbVZFKbDXvWL0CZElCUOLJ4R
4DFXwFhWAtEq+i9Pv8c2TQDIR1jESBTRAQZL0oaDMGwgimWkvSnHvzEqX9E/P3RF
oGRou88RlyN8+M/HacoBSh2PwsbR8AD51ZHNBETFVzef0oMXR1eWkysvH7qn9BVg
szZHzAum1Dcc5wwMQnytbwnxdbOUODh82hGKuFp4hrhN09YYd8z6T2tcI3o1yZIp
yGSmQAbvcjCYNDE4AnF6RNYEpuaE2B1Mp2fSAu34jPQQzJ8dIpQEwlvi1XmcbgqX
p9dS26oACdtC2qtMQdFbci8EQBHVY08r6sw9UwezfswKNZGsfE0VY6hI8xrlbh5I
R1f0dKi0/v15EGHoRkZ+piCdWJDarncP7oU6Yjn1T//U4sOxBRm0hQ8fLl2sMvwQ
pTSNjq6zuUft12oQX8Z02017FRkOlPGSYfwJxsl55DW1TMm0JOH0/jytudPLH3Jk
F0YC3lHIKFbdsYGhOPKYccLoHntrlEqKL5koQ+cOIFbs4D4gUfD35PV9ih3dcVvY
4Mov2s1oJ6RHK6DmXrDUBGXdqVQNu6XeUOWdEkQr2f3kIbdW3smL9qbzbZwU2gdI
lQutEyNtNjHDEjFkkzXy9fYCt/cgHWUYkwcBGUfKm4fNVXsfnBvopTuXJF+DxeZu
8bL8jJJuwniTisqWYYTTE0dGXHe45pJ71bHWgIYOFDXAjJWV3RakMORpdr4nj91g
S5W3Sr8IsssSb1VxOm+/3VxNzIM+tgOXnk1E2QJV7t2NDHAf6J9bnvHxsK/mj/sZ
4aaxC5ZDO0+Qnf9b+JA3lhsEzYZeZ+CcjkuwuwRVpOFhI6nu/t3Ug22ibcAb9VW1
zgddUAjozmid/9owPVM6Hh29jLjIqEvMerNIatkuZMzHh2SUyC2ZPfwPcEK/LNlJ
gbIeRYGGNWOUkxMea2i0eRVuCMlaNQhPJrVrfTNjCmn3ZkygIcskzpXbrR8TNCEc
rZQFQ5o3fXTRVUj8liPejZhMpap1Ld5RX5ae5JNgIqPMUV6UZ2iQg2ano3Lu5SM+
7+gkpxEC0KGWiLmFa7hkzgKdXkD80wvkVPOHJA3XTGY+N6KtvIPQlVxzYMPwpazX
+HYScDmr1KFOVr2S1tmYrdt5qJcpastlTJV7B84qbrSMEi6fvK6xC9A2esqnSnpl
KxfH8qQgGYLjuTH2wvfgSw9xx34IbwsMlt5Tc/OmnGSK9B/hd9Bsnlb2ukbeFdbH
EhJ16IDsenvehzb6IHer+nkaun6y9+4RXwuqUPHxdQ73usQuv7Q6nfryV9wMMyhF
GdSZHMNg8PeCdQQeanh9m8L1Ck/EjJqd9R8vtZXo0xYkZTTsbPZ8oCglRzWbwUV3
DM1R/mRtNZ+nVrhjPlNMaGI96XQnsxBXYlamkFbTnyl+Webln9I0TphGYWipvJuB
02KsdkY7pwI6+0XOoUwoDMWrZDw6Xx5SNtXVXf0mkDbpR7lwVHr663CRQQjeBXIc
fkjKTFUDQbZXDDlSc5nBsil/5j5fz6qgJ/ZcwMZwD+HJEdpV7OjXMvIpmMwf26Ii
yBlFdhlilikNCbbVyOI7bnv3UBYayxVG8+Xwlwh9NyUW8HGob945/U2p8Tn5w0aD
XAuTHACmB1sAmvesUJcj6ShCn0sjkfI4dgjaDEnRRTbfVofiWV6xHFvPWODjF5id
euf2IN6zSXMely+Une9ydPcamXyS5JS/5T4Erix3jOfnOznoNhhpwIUnJ7L4zJC7
/2ebVaoLoUVO+jrKf+btbrd1GVFeVinKPnk/Nr/Kr2mJCIZPy0dMBSTKptkdCR5X
juIwOAFq4k5+y8NVKCQXFZU5nuBX67bl0okXrleYsHDtRa1aaTGPe0LzEpovHzkw
tRId8b5XjYlfJn35Szf27Cg6mVrLSkVFk+//NcIcJz5XxdQPqpcF24gj/Pr6WSoA
p5P6f9CYqFmG4s12Ukbk2Is/Ri46wZzrZUta3ySgBOK2lLNGnJwostNorRB5KEOC
gzlvaHyV3IYVWoEsVZSRlWdAIQQc5L0lW6zr91jaCyd7Ndeu1wE4h9/XhpL9Hplc
Gg/Z7miNp6qnO18KJkX2kju7RgeneJIjapoJG7hPBygRqdD9lQ0DNT+xhwG2LoCK
Xpg2zN938OKy5BeqXdwT8s2NkNpn50R3gqmpiDQmOrBaHAZl6XDMx+Uau9Mj35MM
H5ItLGiHjSg2SDGzOY9bLh2pXsVVBm93XIHkbPPowZyTQILh4eSTVlfTz6xVlYX8
1HSNdzX29aDeGiROa145YGKC8OncuQk8QT48Zv2ilv7ffBH7VqiNJfXcWXTJDmbL
ExmsB/C6AJpjgvNgIdkSzb6Nqiho1llww6g5kD2OAWwfGrt8nTXu3THNz35mEmt7
3IMKL+vE9maQwQkFlIU5YJRQMH6RrmNtvahY0/8LWpKZzCd/z56M85u9Mq9nPUla
FAt6rNfmA4gkVV0n3IxsbZleSC0OWG239LxnvdzsBAJLgxB0gOckHdeDKBzgZeff
cdLjgQTiKr8j7upqHuqDsaOVfENbEKVu6iGk/x11y/cfHbk37X2vh8bWJPKPrivA
vnQhgvp6kn7JMN18s+qxCPUczTUJRAuKTeWIhPIO1uyycb4RLIaSmmEipl8boX5+
FDWEDG0cIpjoKRjZqEIIJZtD7KL44CupHE7ADDAadySsQ+tJejdWsnCfslhesrBl
ZgtlScL86xQIkJH82TPdUWA240aZVOXX6/CXzUGJ4QLl5TCoomJVT8/HWOQiL0HZ
0IwAt8RHXnxJM2rrJJJD+SRKTVQ7lpeihpVtNmyv12IJqbohuPh/vPeJsptl/aOd
b/OfqyqXEwVwlm9nmDCa0hw8NAa8R05YAwFpZeSfS0Ay832auEMATc8LHi1MIAMI
5nexefT6H3v1yuFLPir7Fu2gruHcLFLCl3MmlxURsSGgpUpLJ61yiy65fiEEAEPr
BkvO1/AvNPGmOE15Ue4GkzIQldRarfidNF6WjFzVaKa6RWfr2faJMaM1RcIwwyRs
pv5IG/5bVapAlwfoPutz0xCK/GNK9sXt8hPxJaKYmqpYz35Z9UAEt34WtI/R2xbq
qoQk7YVvVTvwasTvBNP83U1KzyS6XMz71McB4RmIWJh0HwTQ9ToJjaBI4LCE0hM7
QO1icKuOo9NOaDBg7W95AhfEEFneW3Z8M+YIkBe8nFrgdwvnAaPm+10y6czTSgpW
OT3JAxBbWzWSEWhkR6LmJcpr0SO41ZrxPNCUVe1DWUGlDkyqqzY6cKab1PXetZaz
bEAuRlcSeJ4SqkeUjeydU84iBum38SlFXzH1WpLm2otYqUHYlZEtuqcsk1WqQyDv
D61lyub/1XoqCag2WKzZLNiQXotB3SMFXa9kiVI+UikQDLFRY3PMFA8y+maIYDq7
Z0ledtAbr3snTW+x7xfvmeSE7KNAexR/57Zz7kGUwZHqfzaO+3Ze//WF+imB7idK

//pragma protect end_data_block
//pragma protect digest_block
0JnRa7V+xz8VjetLcBOKPcHqP+A=
//pragma protect end_digest_block
//pragma protect end_protected
  
/** @cond PRIVATE */
  
class svt_ahb_arbiter_common;

`ifndef __SVDOC__
  typedef virtual svt_ahb_if.svt_ahb_bus_modport AHB_IF_BUS_MP;
  typedef virtual svt_ahb_if.svt_ahb_debug_modport AHB_IF_BUS_DBG_MP;
  typedef virtual svt_ahb_if.svt_ahb_monitor_modport AHB_IF_BUS_MON_MP;
  typedef virtual svt_ahb_master_if.svt_ahb_bus_modport AHB_MASTER_IF_BUS_MP;
  typedef virtual svt_ahb_slave_if.svt_ahb_bus_modport AHB_SLAVE_IF_BUS_MP;
  protected AHB_IF_BUS_MP ahb_if_bus_mp;
  protected AHB_IF_BUS_DBG_MP ahb_if_bus_dbg_mp;
  protected AHB_IF_BUS_MON_MP ahb_if_bus_mon_mp;
  protected AHB_MASTER_IF_BUS_MP master_if_bus_mp[*];
  protected AHB_SLAVE_IF_BUS_MP slave_if_bus_mp[*];
`endif  
  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_arbiter arbiter;
  

  /** Report/log object */
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_log log;
`else
  protected `SVT_XVM(report_object) reporter; 
`endif

 /** Handle to the checker class */
//  svt_ahb_checker checks;

 // ****************************************************************************
 // Protected Data Properties
 // ****************************************************************************

 /** VMM Notify Object passed from the driver */ 
`ifdef SVT_VMM_TECHNOLOGY
  protected vmm_notify notify;
`endif

  /**
   * Flag which indicats that the address phase is active.
   */
  protected bit address_phase_active = 0;

  /**
   * Flag which indicats that the data phase is active.
   */
  protected bit data_phase_active;

  /** Event that is triggered when the reset event is detected */
  protected event reset_asserted;
  
  /** Flag that indicates that a reset condition is currently asserted. */
  protected bit reset_active = 1;

  /** Flag that indicates that at least one reset event has been observed. */
  protected bit first_reset_observed = 0;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
0GcKOUTtkzUHjsEdlZOOVf2KWWxwfy+6xXPsfN3kuE5IwTU+uosvmYYjnlYWQnMQ
zOECHOuw6oj85cNfKxQG1WqkvDFrhQaLQqJiweCmsC9BfbA7me9/VoiBE7vwpfgw
JN1N9F17HeAAUO/VyyMAKJRrJXehuWkuPKpb8Hv/rs8AnnxIkPnp8g==
//pragma protect end_key_block
//pragma protect digest_block
fV2u/QJDieV1iPW4YsliXEr8D2k=
//pragma protect end_digest_block
//pragma protect data_block
snt/hrzVs9S6sLuYdF79gb7T/zuVx/icgxxsJQyyIZfUdFWOJWVxcRJh1dI8kCBy
7mUIey9RGRex4Ghh8ivtZ/eEtWYtfx32ZwT7+l55km3qHoJhdT2AhdzBbG5mVbTo
nTCvNqEvLfTIi26DoljLXL0oKiD8FxfLSaGVU+Wv4ZK/1XsgVKQH8n49wH0DfsHw
l5ah0tHUpF2igSdyaXg8hm1lbm6qSAKigxlnakr4PxlWLXeFjVhpVVzBRKisTRfY
tsRk/aFV4iZs7fOnCvzzG8808yLQkDS66bbmA64IPHAkdF0+arXFsLz1SrnLdALD
0J/9gmD/gGJDi2T95GKpzTc2CjFNKvXY5KXV9BzN75rnv35YF+qQXWXD2ndSlFck

//pragma protect end_data_block
//pragma protect digest_block
0qFkZ6QoZPBPBEH28+u3GsNoV2s=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Flag that indicates that the dummy master is granted */
  protected bit dummy_master_granted = 0;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
K3NB1WWq8cYOvczVdIHQiXBIohqc//bg+ScBOq4t6YVE6XJqzvgkYC9u+dnQBxjy
T5bmfOkL9uhZmkrNRy1KHqv/QqqK/VTS5dbJ6TONaR+MXQXeefwUIbUF44W09BW0
g9tIkN4DCRHuVYjtFxkuATcq/kcZq5GFk9CEyto83+YzWJblY5GfrQ==
//pragma protect end_key_block
//pragma protect digest_block
uG+VlHC15lEa7rxYOYUMTpQ9n+w=
//pragma protect end_digest_block
//pragma protect data_block
RoznligiANUsa0YGY/+FONnyAse8BSXV2fcaAHt/dyYVeLbkrLJ97OKzDJqRjI2V
nxRt8wjr5ob3BTX+r58Nnyha5mr1a7475AaqdqrK9CalsNcfrO2e8V28y+n42l4h
KrVqU7QkU7xWmgZkg5bOEVwyUsLCe0HwMLMZywKercZ4vJLamhixiuggGkaCREMX
6f8zcxB/Z0EQr4q+b/oax5EYvq65BL5Ym8jDH1ZBb2j7VoQyo9AkmhsdythyKLYh
x4FqVWbr9xqRk8ehU+mXGZCWGr26VB6sjj2rOujV6hNK6RZKWjtV3+wUtiZAuLVL
WNcAxApwTjIcx962lfb/WNZprBRdQhXuqjUU/578iHE4IhwSq3eFAfBlqcNsQVKd

//pragma protect end_data_block
//pragma protect digest_block
QnnPBM9gQKH+GdDMvjSXsT4eubw=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Flag that indicates that the default master is granted */
  protected bit default_master_granted = 0;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
+ECCs6X4O+WK4FOZwmwDt5hyABvg4htY7XEO+aRiQTagK92ROSA38+5rNA0/4EBy
qGwz0L9J7r6xiDLcmc+udKcKTiOBbkU+92Gp7SSSFc/5049nuo4ppNWWP6MJTE5g
VAnRCHHDz+DiOE/c3lb2Mzub4ik0DRuCUsN2kxCozIBUph8evUXivQ==
//pragma protect end_key_block
//pragma protect digest_block
f7heaOIXjSNJSqVyGMbz++quR8I=
//pragma protect end_digest_block
//pragma protect data_block
GS41FWApu0JnwMKckVxV12hT1Jrm1dvfK9Qlic2CnvX8LYTNGPgrME82QAppsK57
6IpufPT6fdCOhN+/NtI+COxJqeh6g9uqwn6BsuWx+iZsyM96L0x2QIGooMRmhUve
lPrPOJdmYGDulWnR7PRJ2eyZ+qAmpQdgGIbU5rid4A00lBV/i6wibnd4CCRcuaOE
dVmQR7WgfGsAFBCc3c6hmDOGtFitk9gULCXlOJdyLqTEOu8xfYhXAswErl7EryZ6
9Fqdv3f/gRqKSRr15vt93i6JE2lBgb1f9BFJu9VZaXaHTMJPB66bO1G7Na1z3TB1
lGNoFvt8ZGFeK6r7FMP69SdtqrnRkD+Y30slbwSiezRHNIqygcrummiDGjGcrMs2

//pragma protect end_data_block
//pragma protect digest_block
eE4s72RqRM7ICh4cdFajyDNSOl0=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Holds the sampled values of hbusreq from all masters */
  protected bit hbusreq_sampled_value[`SVT_AHB_MAX_NUM_MASTERS];

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SS30A3jfJfy5llO2a8k6BpSh494rJjJfIaHOLNo+/dfW1RdRSsCrga0rEvV0B8h4
rHYVzUqYw2NdiPEc76FpXezVOPo7Dt0IK0YBtOWwqBU9veEIqqyI1IAduu6ZpZ38
Qlov9ajkkQCWSZbQntXPijF9a+SSHZ+sJIn2uMWFKx2d3ZCjE2W0Ig==
//pragma protect end_key_block
//pragma protect digest_block
NZPyjbwH7etCPRLl0sv5tkbnuZ8=
//pragma protect end_digest_block
//pragma protect data_block
dgp8jQdYJDWKyjI+kjiW67MP4gD4UF+dSDiXtvzGXG6lOOaLPWYSD2GHuYkHwUP1
CMvFtV1cKzaMrthSwpcimTfXiUVY7H2AJLKMSEoAd3acrzriVfyrRZNDsdv5CyWS
goskIYphbIXBl/LCVcLRGMSXQDpBM4GBMNNBpam1M0aN1e2Bt3JUQC78CqERaVbn
oQ9UZavtx8T5sbGZuaYDV9riVnGdA7m9JYYKfpIGSS7u/O/ot77aIvkhhJSTAq2R
0rvSq+2CM38znA4TWuvW/DpyNMotYD0gxB4erXyorlSaTEUnS0BSoiBnyLC/f762
nNuN+aDCsD2YYpkDP3oxYhaBBXAv/AVsEQYlzXfKT4jn86Sr97th2JfCW7eNHBxa

//pragma protect end_data_block
//pragma protect digest_block
6PHdiAx1vyeevDadN4TkMywjvII=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Holds the sampled values of hsplit from all slaves */
`ifdef SVT_AHB_MAX_NUM_SLAVES_0  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[1];
`else  
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] hsplit_sampled_value[`SVT_AHB_MAX_NUM_SLAVES];
`endif  

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ifE3E+3HKr3Uqk+gZzQwjesWDDxxyK7NqGC4NAxykNd/CVJCAceVJYoUvLX1Rii4
44K6rGcU+MRsYRA+ZjuhnuXPoZn1sKUYyIa508hgESC9ghNx+bUJgnm+D2niNDCT
HJIzJv8SbqfdW4MXAUjwxBklNyhXUEMquxF2vkfUo+zsXFKlEl7Abw==
//pragma protect end_key_block
//pragma protect digest_block
k1q/5w3qMoMrHR5wTcl08TVU8mU=
//pragma protect end_digest_block
//pragma protect data_block
rT3YJ1Xjy91RaJt60vhXmroOREac1vuvb+5q3qRvWYS4pzI5L6XaCkCIzBuCppLc
cAVy5F2J1Ehkl8/LI8eybSsT+CwzTv7zZAtUcKg2VO1r8WSFek6meKT5ds50u/uo
B3JvG7HuEyK/v6z3uEJzFVD1kZWtNzWXs4HVTExlG28JqfAvUQVboPB1f2qtfuPs
PLWIByonnWHY2bQVH4dLmxSqnAimpTrSU7IUPj5YEYO8AZ/ASAgqd6qeiYF4z1BE
+XAPYfwPcSp3XWmDgagVbRF0Jy6fupxCkistFHsy+FpA94MaEW3+fPK0uwYlpXU6
r+7O2+RKgqsYPRG64t1Uh2MTM6F+ydmHtolF+g7zButT2i0qIloGLUUCE9VdWhCS

//pragma protect end_data_block
//pragma protect digest_block
7/bkjz5bK2Zwvz5aIYFySy8SzIE=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Holds OR'ed value of hsplit from all slaves */
  protected bit [(`SVT_AHB_MAX_NUM_MASTERS-1):0] consolidated_hsplit_sampled_value;
  
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
POMb9Af5lXMalR2zRH9XrKjaa0hShNT5aPrYQnp9tWEgANLZR6o1VDg5nKeg9qTN
23UGYiLspFE41S92gyuz+mKlxhvMM0l5k6mEKRTea2ANbNQq56VCI9Le7zLJBodS
ZoKrko1DCEGqEM90EUxBR1dset+59UVAmyw0Q3WwIIZOAQtuxiwDlA==
//pragma protect end_key_block
//pragma protect digest_block
ozwMAc+/AKQUy0gudMOJTlSCyvE=
//pragma protect end_digest_block
//pragma protect data_block
N0+N0Lt7rCPXWh6V920kPxwacc53J+G6rEp9VwdnqmDpeMprVVh+h5Cz48EYwXXf
jc72xHm3tC4C6q5kz0oDmF6AKR14x1C1zsFaM6t0xaAPNXcTua5hmubOjqeLjCLz
nhjQnsn6LKYh2SaxIAz1RbrUyNmt8busBeIn123psicJFFxvu4wUeMN0TlspulMg
2LQje+2yQY1pChr6O35G75WXwNlZ1tDBgl4/0Kxz3bdU7Vx2ZMoDuHXb9Z5SVUSB
NCKLYT/hMEQixNWPNqJpTfG0gwmy6xjxthswg/Ok0+kFok1S8cwDIc37bUAd+OJ7
TW2hMocl5TGFhLiwruaW3wdPp60NDoQWDgY7MXOD+3k3ogM33sfYD5p67/cC6+Pq

//pragma protect end_data_block
//pragma protect digest_block
b2Ct7CRXRFMRjvKbgOpBGzxP69o=
//pragma protect end_digest_block
//pragma protect end_protected
  /** Holds if a given master has an active split pending so that the master can be out of arbitration */
  protected bit is_split_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds the expired count of the cycles before EBT event for a given master */
  protected int num_expired_ebt_cycles[`SVT_AHB_MAX_NUM_MASTERS];

  /** Holds if a given master has the grant maksed due to an EBT event so that the master needs to be out of arbitration */
  protected bit is_mask_grant_active[`SVT_AHB_MAX_NUM_MASTERS];

  /** Event that indicates that tracking of hsplit from all slaves is done before the arbitration */
  protected event hsplit_tracking_done;
 
  /** Bit that identifies if the transaction is a locked transaction */
  protected bit identified_lock_transaction =0;

  /** Bit that makes sure that dummy master is granted the bus after
   * SPLIT response to locked transaction is seen
   * locked SPLIT. 
   */
  protected bit give_grant_to_dummy_master =0;

  /** Stores the master number performing locked transfer */ 
  protected int master_pending_lock_transfer;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8srcIcDrs+6ZdP/1a8XZbJdrzO64+2V1Osos3CsmjRm2zkMAqh/+hwsFHf+fgFPV
Bqovb5yyaZdaI3q3eNctAvhyiYbziP8KbouORviBVQ/JxqOd5ntNcNl3KKOqOigl
VEgx5rijolByub57KKq93+sDVKL2ownKzd523QeNCe7ku2Hci+WMrg==
//pragma protect end_key_block
//pragma protect digest_block
RY5eW88Ilcd/tJ8Ngatx7JnyMV8=
//pragma protect end_digest_block
//pragma protect data_block
Bfonv5l+/lIuyIDN7+VDyJAy2EKlhnKWwW9gS9mZd95hfPZ8aXptBD9lvwEeN+6V
2ohtJAQa147f72pW14ARTX/1CyVtcrdtzS7X9//IYM4Fjgb6mQRZueJYbi6e7Owc
auxgHCJCFZxW4aO9r2R4RMMjr86jCXTG1RL64UFzRXtnDJGfHHqU9rUw8cOd33E3
KA/XiEWtvVUq6idg1lD7hExTIFarYzicLrbst1ZRBl1BwqcczUM3nE2sMQeFvusU
WFMESshZ9Ga+gLEDDG5oM5oLX4fUTF9OHIFAyeJkDq773LZB0UHLFBJJOgZQcwZS
nZ3nV0GqR/3jiJ2wrvDwaWCrV1uN7rP0ix7+ALyDchsP6FxlqnGmznsZ4x6iO8XH

//pragma protect end_data_block
//pragma protect digest_block
RcEHwoci13JwBuwXl5Za2tyeKcY=
//pragma protect end_digest_block
//pragma protect end_protected
   /** Indicates if currently granted master driven addr, ctrl info is valid*/
  protected bit granted_master_addr_ctrl_info_valid = 1;

  /** Flag to control the muxing of addr, ctrl info */
  protected bit continue_addr_ctrl_muxing = 0;

  /** Flag to control the muxing of write data */
  protected bit continue_write_data_muxing = 0;

  /** Flag that indicates that bus master is identified */
  protected bit identified_bus_master = 0;

  /** Event that is triggered when the posedge of hclk is detected */
  protected event clock_edge_detected;

 // ****************************************************************************
 // Local Data Properties
 // ****************************************************************************
  /** Configuration */
  local svt_ahb_bus_configuration bus_cfg;

  /** BUS info */
  svt_ahb_bus_status bus_status;
  
  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_bus_configuration cfg, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_bus_configuration cfg, `SVT_XVM(report_object) reporter, svt_ahb_arbiter arbiter, svt_ahb_bus_status bus_status);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Monitor the reset signal */
  extern virtual task sample_common_phase_signals();

  /**
   * Method that is called when reset is detected to allow components to clean up
   * internal flags.
   */
  extern virtual task update_on_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();

  /** Method that implements dummy master functionality */
  extern virtual task grant_dummy_master();
   
  /** Method that resets bus info */
  extern virtual task reset_bus_status();
  
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  /** Drive default values to control signals */
  extern virtual task drive_default_control_values();

  /** Identify next bus master */
  extern virtual task identify_bus_master();

  /** Track hsplit from the slaves */
  extern virtual task track_hsplit_from_slaves();
  
  /** Check validity of address, control info from granted master */
  extern virtual task check_validity_of_addr_ctrl_info();

  /** Pass on address, control info from granted master to all slaves */
  extern virtual task multiplex_addr_ctrl_info_to_slaves();
    
  /** Pass on write data from previously granted master to all slaves */
  extern virtual task multiplex_write_data_to_slaves();

  /** Drive default values to data signals */
  extern virtual task drive_default_data_values();

  /** Drive write data to all slaves */
  extern virtual task drive_write_data(logic [1023:0] write_data);  
  
  /** Wait to identify next bus master */
  extern virtual task wait_to_identify_next_bus_master(bit wait_for_hclk_before_proceeding = 1);

  /** Returns the burst length, burst type */
  extern virtual task get_burst_info(output int burst_length, output svt_ahb_transaction::burst_type_enum burst_type);

  /** Tracks the num_mask_grant_cycles_after_ebt for the master that received EBT */
  extern virtual task track_mask_grant_cycles(int master_id);
  
endclass


//----------------------------------------------------------------------------

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZGwxSFR1aM4bz3+g1sorj1H1C9UcAsV34Rq0l8+XkPnlqmAHwp2MwhnX33rQHAzK
tqmv6zu9MG7arGZvJe0+icShBlyUz8VgoNCq/vdZ0fWpfUUG4RstHQmvNKc5oHBb
0QbHAxP75+/MnuoXhr6+WqYqgmeQOWbhQPQxBg3Eh59B05CAd8Dviw==
//pragma protect end_key_block
//pragma protect digest_block
ZZyegbzIYKbU7pl+T63BpMsF1Ig=
//pragma protect end_digest_block
//pragma protect data_block
p5Khto36bNyifyBTi2dT5bhSF1+ugNiwq8tBfiBbn56JxkWkH10hH2lzzFTTjozn
JP1FwK80OX7a6pldPDl1MBbgeckRaImGc+HRDgZJ/OE9qVvVwmVdShC4d3dLd/Kq
UvrlIFIR11++kXlEk6dSOh4kDHXmoKIGt5J/rKiNbui3hDbjRiHt2KLQEJGWgUbJ
tCYR1cRF1oTIcwXljNGP9Vpvb+VNp0346MzAqsYosa+gIoZ3NQvrJ3Z7G54VFmo6
GrC2BWY+pM1an7oi0FBpNY1LUBWPiEljG3+yhFjetDm1tOgC5l10MzSneMws4/AR
0dqFEuS5+HXeIN70DGj64QDGytY1h232fRgB6cRyAOFLeYBTxnYhUhScecWa5dci
US3f8Ec20TV+uQDJGReXgKgm0TApJsLhl7eke5WjKCoGqI6FrslbYQhxD/N/MHKx
Ek3itQmCy6RSGhR2g94lQ32tLBGLBhWwCtGgIIreUut+PevZyfLkhx7RGZpRECKx
rUmADQQaWbWCUY4470mdI5U0h9Gfz49VsUwBXs/APItFHCUHc9hlko8s4lb8keM3
f7+qCPhQ6RiUkK4OlcwEj3F9SCaMjLnR4FYMie0feSZDVOktwC7EVAu3nBbhB7dE
8FSydvCQzFQoge5ggqf4TuY0c3MTMvrJLVprDkAazVtVD9hlX2ItzGHL53qRCo6J
56I3Blf4JpZaLifurDIdAj9ijgt1e8KsZAhRbmvy4lkbZwBs9anwxjYBdusKGYhz
21MQLXx0AXSOVpibvisNlZN6b3Qcu8QrPb0m7I6lT7pn3K5PunjJwWlQ2/uwnDqC
opUSST1JKJ7Za88DYDByBkGcoslxdhtAlTEj5thV9pZPSR3AIV+Kp5B93H7lCzXU
Qfj4k5mAqKrtbmv11Pz1kOrbQ1ALKhAPfhzDvO08Pu5TfAx0tRX4uHWbNjXT/hav
EUPAARNviLaqWAU8qsbIBgldqFqEOl1DOt3MMhdk5+Q=
//pragma protect end_data_block
//pragma protect digest_block
++9c8thTyZEv/CufbF7w3Le2FdE=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NIG7/hY4L1YniXEAJw+gO1gURjw5VfyMq4w8WSDNjS+5OyK++tjrKHCj0VP9hKdj
kZVqMaT/UVqnz3WnMAopwQW2AMOnqFmQU2Q/h0BPKszyyjtiypRdK95PQZ2wp1nj
UiL56N56W69fxoldrSODbOcje+/t45xPJkApqLU/vbMowcTYb/e7xw==
//pragma protect end_key_block
//pragma protect digest_block
ib4c3Js3teS87qRf1murj8aOUcA=
//pragma protect end_digest_block
//pragma protect data_block
HUfbxLUv8iO5gegIg6BmyzkaxWrg1JL4LKiulB0LP5KVJU+Du7nYvU1ZSaqI8TFX
NXahLduJwKyQVD+jbtHPkIbjS8ZIHvCur3W4Mfk4I+40XVwDGvm+kpup6JSybGji
DELuQ+7sEYm1HSdTdRfHjREHzBiMtUkN+Uy6S8uYqNpeNKK/TktNqybVV/u6JaFP
7+QKqNQrhG4OQnmluWsM3UGTXaI33ss3on95Ydj88E1AmCVUhMNV6wrZrKLoZu2j
R3GPFsQnDkejc0BVlDoB5Jxfcw+SaHptrLFgui+fTSS+lHu4YV6oaO0kMlUaTqb1
VDk4GJ9ADo4bv0NLP44hZjLonsbWDMIVLyxZbL3ts5GCHQXFxLPksW9hAuLk1/ID
6xOpGnlob1jSqlWlcTFNJZztEUpZtODswHSPnoy93xf3ZZO4vITpjODBTKGJswlA
467psup6jf0d792ltfAZRaOztxdDrbneAyUdHzd/PutZTjF9GIYb+pfMP00eVtkR
+YuS+/n+zPo1BRmKXZj/5z/H47myAX9n7UIHY5minlCm25VfhAEs5ntKhSEFovtk
dqpZ3ybEgi1cUhygkNV44nn5no8MzNLndQjYpdAlqCfR7vZM2Y0xCQV1FgMfPksg
VzNoxxvOjxhK8FNTiaQuQObCwVEgnzyltL8nxSRxzCj2DxnxZ+OUfkhF8mpAeo17
CbHWKm6BVJhEAwYn2shW3OJ2sUDkJlHO8NKKcf5GUc3bLpyWZrij2P8HDzTak9uR
0d2UCEJcHmQwmaAip7tWMIPM3rR98Lc4WlYnTjzM0rhxV8bapJpxAsF0jQLELNe4
rfVD2h5A8+9VAoozGfOVMRS/3cywhskknnhXbKFAnd2CCX4rHiLs6Ct1oeoi1/u6
YXNSFOZahwm6HTNbIOkkkZPi0uRUWO63agBo7qYFOVQEAcFJuzYH3xpiYgfU2Fdn
t6O9SpHTmoplapXzpF18aJuI3yQuQYbHIdjnHj+ITi1vWPcmz1MyapD1Dro6yG93
VDxm2m0qmHVDxJ7V/M/JN03VGuqlVn6krRJfa2LSs1shpmGZGVseOtgr9Q8nahQ0
T1GBs+AhKEsp+wdC52cvO+M3CWXNt7XwgQiPk9UEwXosKKCQpogCbB6SCXSorGg8
9Q5JDP3wQNqyRNP5DgZ2fAxij8eS03TwSig4iU2ItZpm4YTSTwKIvkLki5euDZ6Q
bAMYhEQmvn4fPxg9tQpPICJm9b02YBOQPKehMuVXd1gXudpb/OPRitR9n/XZ6fR2
Zm9cBwyInbyrzwBeKScvNkB8Zdnm4rYjw/39ESLJPfaSnnjYMLkzwPA5fowdaM66
Z/08PxUmP1HexYenz9eXIrnpSELlfPfei+2fh/aWCzKzt6JshQaReg1ogeACE/xu
wOA6jm37G7SAJnUDukL7vomsVneRjJ12yfmx6TWlj9Dl631tx5SUYZZcWsFP5mnQ
7GwqQbODk2rHwvfmexXQ/ip1gEZqhY8aCiAB9KwpURmF00nbHsQu3RXYqlSxdf7N
S/SORKcT/VfE4+KOGLCMstQDPm++ugKyiyJtEWZjgPWRiTitXNve1HrIrkPh5DzU
Sk/rLs1wu3HIbeNVcYho7aF3BRkVSqANGxB+7PwJyeSYrZyzPgt/muu1X0mxa6ni
nXsxOCfaQh0bhTIgnIrKmKijEATQ1PLe1/11NvLDphv7p4NLZ8x2jffSxBcVmSXf
Rdh4STRWNov/TPuCsoJo+5erSrj7A1lwwj/6HJaAsdSKkJmLm44yvP12s4KfLVVH
NyhPh8BzeUQJVVY0723PCXZaMtQqvgHEOFUbCWTqMwHgbJFEc2ObBnVDELyqMEac
lJKVgfo2RkBdPOe53ZRTYMsRAr+xP3yOcGrdtmmEhFNed7RSceRDkdzpL2XXCNAc
FRjp09EKxAWclscfGtmDuR2Wd3kHeKgjfp0V/E1txIyGR8LTPimmEKgHfgpYYj6/
zNfw0BOsZrNTZH3gD5M1a3FHkGDgy1zprsjCO80znLTNeU0/+mtTwh2ex9P6NmBL
CATqGAvUmh7DtjZt3cXMjH26srSors/FAjz5J7hJ/UBZP46clquC+L6KRFf5296C
m4GpoozT8s6TcAw08KSRet6waKPAqSMyr475UceYbcntM24nu+EzLxEH7WHI7R+o
iDMRNglkrIcZQKIdoLR/OP8ftU8d9rg5zreGLOavqHcuxdo10HDP9HNVZaAl2rif
VimtE+1yPmHGbkH2C6GhrM3bSIa6A3Lf/ls2fhMua9wBVbMQ0DncU48LTxc7A4sC
cIloIjzvn1DS516ALudhKInaZLGp8NPxYsqtR9DHPZ75wtAahkLdwKVb+tAMrZ07
HDwgVAfzsAnmG5EcCdqmmcMcyv2GAumJNkhVDeskAM/xSMhhjw8P45mA2g8ZaIYA
VnuVlU+waKSvuDyN/OF4bL52yjQWi/7bsoO6Uavf9DCPwOt50jpNTt9qafwKffVF
JYO+1vxbGuY/+KrUQ8xD970xAyL4Us5JTi2YabdnZx/YNyN0y4xQgzKU04mgh52C
V9PSs0+j1j7xYov6Q3ciK/xmXgkbKN0eW8OzAMrVOhaP2/f087JN56Ri6Ecoh7cl
rsHVgqhmYHyrDLDxfYplfatO4aGw1PKPeKuw5LHbtrhCaCmANc657wTe69SguoOZ
nGyV1qJC4teDoRpCus68MHI0Gr3Iivmq6Jwv0CF/6ZkyPRD39S9XdUrEgi8uJ+qv
gkOsjT+m8RkhhUb/tltjVr+GaG/fa4XXev9DZxG0CGouA0pLvsmL1l6CMhlZuEUp
LoVidAwj+Y7/gFJQUX9g+C3XYdvAd75rNA7kZX0X9s/jHWTHsI9rbd26L0ovq6tk
BbruyklZHyizTVnlCoy6zfRjPpzVS9i4+UrzTl71+53LRE1VLZUs7csdzBMR6z5t
+kz9u8etHEYjvjpQPjwEouHF/PhC0NsyQjF5JYXlFpw0i0rpxucsY+pt9V6u4QD7
z+SuUDKQovOg8AYbelG5sRpk79711Z+Dbw9/c/6TZ/UX7aEhhRRx9WSgXXRH9Ai6
KEZeSvW2NSo7f1MrNd7OPNee7FyhRRrQdsvu41y5qIV1iw1j++MaciK298Jtp3kW
gTiiGCF6B5AyJlPk5gV+ZrIl364CKnLFy9jXCJ/PeWVkkkWcUVi8qgqY0D6foUvC
IKeVF0sXFg1E50iKqxVuewZLcqWh7dTkXVuABMnBVg5UwlguWkkTekDVL8j9VF/M
/LMtmF1wezZCcIOucF8tQpNxeINXM0t/EDSKcCPdqaoZCbC8HCgN2VO+PSJ+9Va1
G13n+oBWqlHC+VIEJgLeQzOH8NGffHH8SMHDa76vJRsYpHPVA/9PpbAFuz6AfWQJ
riBzQloCl8bMrQ+q/VZktHM+C85KPqr7ZgeIo8dPGdvj0riUCrK7gqTrADveKU4n
6pSZ9FhQSSL9KY05g2NH/PyMzfa4nLObmJOEsLbuMwKnA14M/hQB7R9ygxVBRUKm
kWSe4Boo2yBq31deGD+PQ8/hZli7Y8b9Vmvux2FkjlP/OEtiFxxSSGydeOZyAzbI
54IMr+iNSdGmhAOe5fvSiILqOemvW2Ml0yGikp2Z6yUVtPwTocehoyl27Yoq7q4R
ceRmzH5g/Qv6bAuHst5kvnV+5pBSJVFBmBlmd+3Zaf1McLQ5SAjKkhfxVbmEKs16
wQsq5zjyQix8tKVdHhPpMM4VqveYDM4LxqKCnUfJFAYiGr0voDzr832D9jhlz6Ah
tw+yJ2O9YwwD8WHB5fSMgi/Pt2nyYHcVBHHrgn0R/F4W7hf9cfAHJFAAJx+2U12O
Kl9/VuMo9TyAUpS7cGbk6deIboQz5Ez+ogTzcfKHR3v4yzOQqEg6QS0gcoSxKzin
6I8emaOEqn2NOPD/I+4zkW7r3rRIoOpe8N0+P6+We3spnyjbC2YenVzUAOfwCfkf
F2LI5F5vK3FTsMgFTzP+qothRXs2RHniIRlP/iv/kQwk+Pd2jzAENK5p5Is1m/SF
vYhU73A0p0hjW4TfaDvYivF9pOa25OPCSiQsL3E5Z/HbZBCiJxJ64PfOyD0wuwgw
nEgIoYa9nUWQyL6AoYmj1QtwBqh9YhfziH/FPWojW4foRZIcY7jxjN7vAZ5Uoi+y
cA+k8MUdpjWBksF5CIVaiOjIp3IYHJqlpKVtlQAQdZToLjrMELbMvhkb1bg9JPvZ
b3g8c9HCFHPFB8QXyBC5RzFOmNNtHZ/fJC4nL2gzH0iCUFd/GFDk+wyhrKw7bFjx
UIxi4HRe3dhh3IJegtzL+wL80fDrIp+ssx41FLD9m3yJXh6wAemC0ddDWpQMq9Xe
8QW7N67zFJaTyDjBknQWZ8enGX2ufXzmf+c8QhiSYMm+Wk14bobroDKTCwTbOBKl
bIZpr2+7Px415Spy3SRdLeIAI7JMpx/n0Y48elWhFua+2X9l0/I3AOb0QxghnSNY
0efN2FkXo7/N+93dDdVqz7l1ZMyrJ98yX8RM28GjOYphXPnwIsYIJAdhSGwGWVRt
FZ7//c48VYrFYLJ8aq3E0jE3eMLGwBSkReAgaCyZazArrE2pMajBk08eUbd/kiPJ
x9RC0NE4wp1pYRHYt/xmwj5PC5nE03Dl/V88urMZJ0vt1wMIPjUvD48vQSZk12kF
OdrCt67/NDsis+VVLric4e0kb1vRaw1b+drnoBYIjVGMBDTyogg25CymkpzkFWng
J8MzDvBlILEAaU/ehgbau/1bvxsMPedAo1XXHlk3qf3t81tzFTV6i/nrSNYoQRpd
6XXd7eGto9TNepTbbedU30udoJoX4fXYraFxscTnzXdzad3WeCHgUB7UpxaMdqYz
XV3Z2zXwv9NlWLbZGI1/vo8u2O61JTgvjB0I1fKq9qvwsBIlLs5Rzpx0MKh68k/h
Rm6KkX8f1PXOnQ7HoMVXb+8Lw5CrzB1kB3z1ZusPYpKp1rbuMbDHi+Xxbd1TAo7N
XzfxMdSEwjOaYE9MuO6B5xm46uiEV7QnYdvRD4EzQmulyEb+JqOjtjjW37ubsIah
clyckgKF6k7T1jc2TQLgk9SG88vbgIobEf9fAzMPj5ad4v7tvWRa8VtJv8RKKqUv
he8PCntEeWOLh1Qkn8W8TBqQ9csMi/+QtdNNmnkPVP+ckbF/4j/5gWnNUjh5+PYZ
d4dqeINg0Lu+FoiZXkqLeswVWn/sUbCe8CmSzhfWCIQ90HDKT0XM1yiXZfqJXmNh
b3LeHCauVswLOQbGXkYSfKyXllnmN0MDRX8B55+wyJIVUsLzZZEgc94E56izILHE
NDTp4LWLjO+qJFoqUtFrNPlB9q7I6+q8BBt9reyPC5CxQevN9rk5uPFq23RJTMNV
VRLSuL9HzeevCQ95ynE6H8XrncPr4O0Luf9SMUXYkNvQDQ7DrXqCfYu+uE6PdRFP
WyI8U/lNc4zQh2vuDHuNSfoK12l+4MQEd2x+2eBU/SOtQLZOjokOVpxRnSKs5kFV
aeWAODHLiB/LPX//jqzRARW+xWroShub1C7i7Ugt0asN9jL0PRbhmKVzy0iWfqYz
ZTMnxVxOblGinPs5ym9WsCGEUAE+WGHCjCoSCbpZLkqSBGt/AUZjgPWfqUa2x9RI
zgo6x8rWrygU5teznrH4ms5J5Kx0B35alEJUOaAFEXmRY6Tz2oOxdT92hwDHlzFD
McsMeNneNLnfIDiuYc0o02tjDe75vS0IaCJBYqlW5lS0hsa4B8Z2WVWbsa7RNsSa
BFpgemZZniBJ9vzcu381kDrBG/UG+AD+rMjB7mTvb7RicdJPjfvRGbETvVl3FDZ3
Em1SZxbmyuh+R/biIoLl6hXSLrZCn6FibUvqRlFwhXRlmC0iM5vve6XYIZIiSYEE
BMCVxBObq+TbG0EyvosJWq3vJr2u5Ipj/Zv2m7eSQqGi8IczRuHXEMzhs2275ghy
qIO+gwSqvwhD0cw/Ux2tdRerGIA+F8IbGGxVQ7Wz78n6g49+r0zGAmK3tDKf+nJj
JH4XtwTGHd3IjKx240HZcydt8KIGtvp2UAsuo6XsqleXUM2UhqO4e6tbP14Vkk72
8nv1FUDh5Bs0j0boJi92/xCP9fsvqQbpruDfxnDOsCn2mpLRa+Bix5rAmEaqT5Pw
6irjZrfavX9LosEwq2SnbCQC0t5Lej2+KwzYoGgkqraxzTz5arOwsXPS3kOtHZZG
Zk+opu9uMky3LTvNGHaR1WiVysWr23WdwMB+0S9u6qy4kPW+9DzzJrgz6xT3IlDH
2IcYsMnHsotMk91X4EOxhqGvwAJ8fP7sZrnrY5c/Gca8talaRT1VX4YN5MAO12QU
bX8kK30XLPu+7vp7aCNOnMDHJtm9+WyPahdLIozi33HWKIq/zmjlQb7171rBsee/
J45fm2yeF2sjtsL2yd1+mBXUlgEnxDsSRun2ThYQoKNiuC6Y4XC7BXAoOrVEGuME
XCLrYOA+9HOgsnT/YkumWdE1jAeswA83/oCk+X2LT53JEimDvUamcInXe89+Blwt
dE34LIaaXAiBjapRA9t37VzpXtjhgEcgQrmdQY7uMlTJ2QQsa4iCubodiszqr34v
0cpy7hw//2UwyFViVdelAmDxLDiaucqJLvfHKoGlhAkGgufZj3NL5jgL3wYM93VX
jnlsK0vbJW288/5GWRcKduGMPxf9kVwRpK1T+E1YCIpmw50YtYvkxDCM6+9QX5yB
P5Q/YX2+AcMTkkKDkfc+8F8+7PBnNEyR7+HY4vQYxt9jU/RX/KkgWT1Li0AN8c0m
zTRaNml8ubVHrKZIlVMjzL0a+bLWNc92VbwDcGnlvfkoKY3EnaSe2LYVX6iT9ItL
ekzhKln4+TjDDezonoWFMzoj3no4NLlYCAc8VWQ7l0wOjszfDTjf7s2nuDmM9WXB
yc4jzo/m6xnl8375a2bDSEKiOwo1uwp3obWt/Ws2vZE20SWBbozBMI9aaALbcPvc
KPEzC2UCarwA6R99LdB+InEav9carMo0VuFnHnmAVrQI0RQPBuI/JrQKtgA0Lxd6
C7NPsXUvKDrJsDEZnYFOmu+t4Huw3v5U6OIHLxo9XUZ4xq/4eOpmBWFqyRT6owGA
PV0OrwtzsgnoIWW7QLf9lQH7CTmT//f5XS3yvxBb671kpkrAttqU45nDMEBqmlbC
olHxiSco0g0UQ9cqjt7+JA3TXgy4UUzQBUsdHq4rcT1lo/ZsqBkEIhdqeEtnYHHl
r2oZYXDYkdwjmy+QFWdMSsv77O62Zx0WadNeXH5gTEnW1r5UxdrE7A0fOtl3KIf8
3qwNpqxCe24+eqlfQ18P+3BRSakkwo0+6QO78ebgDzTx4LGLSg+JpUVquukbB37i
Dpy2s4lI8o3sYC7lKURY5kgQiefnZ/0BXMPxn+TXlzLsbUIeU61p4egqTiKLssAe
4DkOH0MFI8nzhF0T/5Ffn8AtEjslCictvNPxRu9GbMsgTkR/L249XyjNGIXdV/Ed
psL9ByKSTORN9yGZcjW4ahhtB+sApuFk0LqKr6193PXlhXg7OGu6rXbwc8puA85q
e+lHEXpeeSNpA8OaIo7GPq5A1w5134eUYrXnBsBHvJVlP10uYTYJ+zcgtGoPwnYB
QmkeY45iJTEyXbNvi2B+lr/vHjfqgMAFBB11hf+n7jpCXVhvbWwtPM1dEdhGwLc8
F1uBBYcuGJla0wXdMHwX3RhePj1O6vkjMAzB8iV0fw89qs+ZcVLIxoM/jFGwUKxi
EGMGjOoqwqouPJNnpcffz5EpYchOFOLGRCCwaY41Px3M1yFN+KQmLtx58Q53karZ
I6agu2fz7sSnEK1sZrXKSMvmXNOftkbKANWRTRQFWZvM2m1gOy+OdvK8olMn+UgR
+kFbEjxwQy4f6bRjxmZpRe33nWWp/fsrA8fiwEw+jcknmuAJc29PqC4yPZwTZ6Fz
rRYbV0eH1wZDq9nLTwbCIwtfeCzyIEdjK+1kZ1eFNRPV/g9ii/rFG6VGm79lyNJY
0rnNgrsR+B+A0ePlXsB1NBNqQAVWKeESZPa8puLkKlrXnNjHhIdsY2c7ezyMVuMC
HJuSwNF5HFlNUb3Qz0PNAb9AF9zbw2wzidWcPi4kI8igKS4a0gJiBUM39Kw8ND+P
Sm9YXQqpS+JYi4xMeUe0LQ0bl1SGLBB3M9F7q9N6HcKK66tfw5c2aFxm0UARIKwm
EUpL2Fp6qmpHkLq8B8E3cYgoc87hZFQCdv3MEd+owlsvPjI4AWHYci9kjpIt4/Gq
bOV7UB/yLeZcla5lyg0P4fXePHb22c41Yn6HxbdlInN9YYQXN5qNBpZbdPU5A0ys
DGqRobvULGo/jGY7EXO/gkp8daYmN7VTXjqwUtwo0Hr9xGs45RIMCoKtQHENFYvs
ZuPCcYOj6kEuewWLpkicEQevIVVHtHJ5+MPCQTZhFzp3Yu0f3uA+eFdiiRnTo3Xg
h6GhcpJKAX67IeDPf7Kj9yYgjwHvdl0BaD93hDsS6exHO8eYL3pHl5DOSzDtLrcT
ZpeMkbHowsifo5zuBuzpWpvsTTfHo5AxJvYbU+cSDy6BF4Qlkzt48BxHbCLAJWQu
+IjnWlPwo4GJOYgR2K3QhUPPlR0YApr32u8SidCs0/mtKQuigVhwMyfp6xUD9LD+
QB1dBYSEG0iYxChcMouUW2aZJs3bsyZbJinxUnqaMnM6sHX2hb15BuLbQKPIhpPR
3ZQts9c91A09m55x3IoJ0VoZCflUx4l0WL9Bc9Dcg8TJS/X0Df20+kgu+r03sm6w
QzqeWQaZdcJlO1532+MPD5Ubr+h0vceGGfMh32WSQ9NSdcHHYN50dyBwuhwVbnv0
vIb6o5kCeGcghZUCpIgYPmFsEviV3T14zOBA0XY+YTZkkoC3Q65m3ecaQQ+KXlBw
KCWMpsgETp3FgQCbf/3etAV7Mx5z0vtNOXeq/raN879MRrNMcLLSbsVw/FS+H5Sv
HQ+NbroZr+ysL3Hsr2uTSOoSCmDDO4DaTwB/ez5QVDRujEtj5K1BOFmp2B4+cQaD
9kBSg/YgrVHC5U1KmiSOL0aLhKa71aXH+Kes4EB1OJ0ZglOdHBYvHeUx8xJlGBsD
3g+YzrDNdNmiFsCRrNv2NoTyhQ2LMA2TqyNsVmI6/X6AWNWX09zUMztEmifhuEuW
AYM3/3eOt89Z/sX+TXZjBkAVC2x34d3lFvVE1zrYptdVGiRXb9dAGtEE9HiAnmrD
wbZmVWvlHxOmVhbAQzsFPD89nLKpGuqa4MA0H32cCG2+LeZ8AztDhwSG9JM+01Xz
QwLszkCyxB7eqy8IizhG9SfupUtTZqY2r/TVIYTPy0hHXX10W8KGbZKS9dJN4Un5
8aXkWujSGbi9bKrjaGg6NrXLaqhEolzd5/X87wVjIjxSpH108uA2LLs4Nvv/X6wr
U2ylZtxoMOSoxLYmYYyYg1jjhPC8NNxMjjJQmxcYVjVX7BeR+T7JTTeVPFS2pVXS
6SVv6oB4LYc+slV7Eesj/RiIs9Mu2FQA2Bzp1lbSU7gbh6XS/Uo+jhSyQulJRzZU
WpzlaAdilwnTKFXoRlaEYJEuqodUWJQakmMnff5H/R57P3MNmzle4TK0G+r+NSOU
UrbIr2RWahHGoAWn0HRgqAifl+RxWunQbwLH+dsqN0GO3GDLdGtXWv9u7jPfWP6x
KX1GGww5zuCz0P8qEvzYpsWp5Mah4YftAKFFd8zGiIKpBxx1pcrHgSE6SPpQ9Okq
3kWJbQbucLLRmGuIySFB9n77AweIvVufE3iCbzwZhMQJDhV3zLw7XOS5c0hg5pgY
SbKimpZjHwz8t1aP0LOKgtrQ/swqV14uj6pdXcl6Zp2VsVyDQQ1T+9s8+1dW1p4K
atJjeDhJINcLrXeadPyx7s0u1WTJ0Tylv1skj1kW/GkI0u7guudHlChsEoFySYeN
KO0VJ0MPrJeWUN79agwFoc426qVj88zXXMo9H2uVvueorGf/XAHQxzO408hE25mu
rl4sFy0C155ewjHJ0UCZhFV/0tNHHSK+mGvfFxocVbz9Y8m8U9pi+HbeeszYja+K
wIg4SA9DKzllNsa2/5xdrGbC3D0jx3BQMim4dGo54apeS7RwbRiu+qXD4cffJr2a
mq8Zi8/gMGB/WK1JwHTIKOW97gBuh7xskEFmiEeNXQIqFCBaDdNzoR5JRyUQPcY/
AIgdh1uFaB3942pXCSvhMVcYaPJDYwRREgpvddTH/TDldZaul7FxB7WXYzpood5m
MM42tSQRJytXQ5vdJfiYhKmE7cfYphqpNA27j7H9PSrA4leu6RTHNXOIV3YawfzA
UjgHXJEPN4EaDsMtGiqWIKg/GcWk1XGKJ7aogneb6x6Xh4UfoQ8hT7kByuz7At+j
rNTUjxVqbo2kVG8te5gPQ7F4g8m7yLM6dweXUQR8DeGA829YaFoBwXcLO03gYtLK
Xkb2jqpGArbYhAs24cETSFSy6ksr7StANjto0ir3VEVvS5QXOtTMaxlHCCuHZGK2
4Vcph3sN257OK+WZ6gUTY4Qv0mSxmUUI8EHXOZR0YABNWn8tei986lLkFWe8eHbz
I50nFaS5zKaDKbxW0GG6cEOOTJGDSezOgsc7KYp1OvZ0P131wL0yqLqTsWYQI7Vo
a8K/I9meiU8oc1Aj75UBGVEQHsF5MqRXPwdvRcd+3gmdHkJtoWiQvposXE2cufCb
gfk+e4W3TAocVSdDNPIJ/+/OyRta1cvgndgbnq90Dhm/JONsHDQyJUus6CLzqk70
icyXOcUHy4MQiSgToMFx4KRQH8sGNL9LM6SmhdjsbYkEtt605+CP+L94luhz6ujo
5lZeg1i+0VL6c5koFzDrI9n9YSji9niN7IaQwM9YaZP6KKOQm9onhZ8wGi9nL6YU
3uKhd+jsLH38LRCFt1NsZMEk2WeKkb6+yv/xkLl2IBYQkJYf7UXfCKXSx14lwWtA
jRm/VkHAMJTfy8nJmwA0u4H/hEgqyuHu8Fy/aulxH3L8J+Df/DtWIPiIMzjG9Bbs
xNSpcARdFQIRSBI63WNg/9tC/MWuiwMAZtnHMk1J4xztOjPLqeDp+rsoMgUL6w0h
sKDkhSVGNzOU//+3Dq469Sq6HRFoDlGI1LEsZDxFAw/iSB69kmnJVFM57TLbveul
Tw8kDhX6mAoTAfeIYVbpFvJmJ4fTRVyLj/pUJKRq4t76qIzl0MyPmwTduB/M7QMv
AVEquVEqrfE2vKS8mOsLbw==
//pragma protect end_data_block
//pragma protect digest_block
uo4oPPb2OiPd+gN9btd4/UMEFJ0=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PH1BXHlHUcIZ3p9zWDARTdopIRzTNyYw03rMUEgziVkHPl74ZDEgBAB5vQobbuWt
yPgK4n1nMOjbS16yddQXh8pZxmuAksO5+4mNfBVNeA27SBWMufEFsQm5SXZu1uOr
UjFnNkJhN/bQ5Duhzs64s/4NDLHHWKWY8NJpWeEjU40QCo+EDEUdTA==
//pragma protect end_key_block
//pragma protect digest_block
ghGSIDH3JJiZk3GYuPFOXRzNhv0=
//pragma protect end_digest_block
//pragma protect data_block
H25Fbrs2SBkHu47ur+dVhM299ZULPyj+byNhsX28aMJfhAPjllzXM0Or8KT1KVwG
9p1IBsf1uhHx/Rmm4hLqaw4OMMIwF5Cs4Jk/YfuTXiuKR6AnvBFqnwyapA4xsrV6
iXurxlfKfq1lIjOc8FAL+i/dledR2YrdJWnoWStzwik6DjRgxvw+Sp/2W7ut3Cmx
964M5+8jMZgkNaKfZpUs0kS4Wak5s9lD9goDHOwnHUAM8FV5+Zq1p1aq4dFvm3Jt
khIiWRRKM/Ww8H1hLSCMVyPAoinY6mBclKsoCsPo5R+yJGT7JGMyWwHYjZIcq6bA
ntKgRJ8of8At6PJ8x0qZIGWF3Dp6+C2yOwcvutihDm0EJup9SLg/Do2DkjjmBzFI
t/6nN1aJn+plyUZKgShHMg==
//pragma protect end_data_block
//pragma protect digest_block
lvQR4z0kI3m/yGU2g0j8VbaBdRQ=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RpcXsLaD+aud8KHreJ0hAlw2SLjXMI9svESIbP1VfjuMqFVM6rxrfvg3Gho9OCRF
mwxVGje3VsnRLtqxqYaR67Nhn0000Aaq9sAtGFJHkmM2Rf8TBoSiuB6KSTJDsihr
Ero1m1AEtaKVBgA6yUwkkEiRQHgqE8KdzzgXuen/eVD3o0A0+3DacQ==
//pragma protect end_key_block
//pragma protect digest_block
/VBVS4EdM/qpkzseX5G4AbIUX9o=
//pragma protect end_digest_block
//pragma protect data_block
Y/eUtt6gDeakgORhF2ePK1I6pIgSEXkHjzhY2FaJ7QvnJZhZy5EY/ArtjsNjOtTA
OnLTSsLCzgAQML9LIGoTumUQ00hHhk5Vxi/ZpxzSNuzeZh0Ck/hX57sFvyDtu8YS
SC+o4Obue3YaoATYiRUnEdR/1TcLqEnZDQHHeFJ7xOrPyy5izMWxqeGe3sfa7tXF
spF8cfhJPeGU9mnLY1nMrSkBzGQMmF48MefI1+W/jUhZlnraiFE1bxSkYeSGtCw1
Bp8BFqXO+NMmn9m/Jk3PZOHXIdMIS02iTpE51cR6SCcZxjUN7zAX6y6qRKSkcpjy
Ne5QSQUAW+1mQayXugSbYv1JbdUdrb0iEsUSfv7VHgdmWmDLJc9XjQCCBU2/xAuz
vmZ9Ycb9mzT+ej70UloLhlCCGIk5ngSSmP+mIhtkBY26WvtaXFAuy0EWj64QfpOA
kpQiJj89dyIYNq8wMW5nFW5d1qP0FjwG6QKHQQaZ2CF//cDIvH58Ggkd5VWHjGwS
SvwTuT9iLmXQn0BVCsvS3KZJpEvMVbUQl6IfsVPy17KR5k9jRGCue8UeeBnBa1dg
iz5yvddaKyjqTVC6aFQ8KEjxVFfmxcyWpbzKMmrNVMPQJoWjoqzdUhKdoKaIwODC
D19Y/WynVp0h1BTFfgiTXGWwBeGQA2eYMdx7+xxele281GYusHjkFbBHa5XC5KMP
/wiaKNmHQMn0Ff7Dh6MHb5oMZpPsmORqnz0nNdTm5aLD+PjGwtj9fYc6DLLHiYGS
vMcN8sCJ6j8hiteiBMWIQI6Ubsm8EjqsdptK6ZjbRccpNgvWtms0EIsyBHKg/9B2
lcUUJyWI7xT1FZa0KjyrAsWKZEIaNj6G0uxoYdma7WhEt84jLLMtF4UD0mEVGqSo
nykfBKuLuTEUt1OSJxNlildg1Te3JRBYe1e94rf5Sp3hZ4ZgiP9mkEkcCeYFcpnd
IJ6AH6ivVvk/eaAO4OJseA7hGVaADqGkFmmP/8mzv+5I3qFCqPfYicI3iWRJrrTG
nXMv4xf3k/EUZ1ou2cYXcJorYQAszcwfyef308hV8urjldtLQQjSuitOd/oC+1k1
TWqDHTrljKEQnOmI5Ax2VrrW9JZEkgg+DJNBAv2UQOxmSp5GTAbvvTeIOOg9UA7p
WE6NHe8GtGBpfhEb16+YqQ==
//pragma protect end_data_block
//pragma protect digest_block
61WGOgMMJU/g/a/MRnoF0eAtY6w=
//pragma protect end_digest_block
//pragma protect end_protected

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
SMI68NPC/0TGzes2W7Si2FeleZkRGg1F4i2vLMwWKPNtwlM2HmNDfk7Fzz5kytst
f+LxOdcMTm2cbMzlmw7XGD1JwAqweBUh1e8di2aoygoa7P9kSWb1XFf1krajk4CA
nUcztfJQmgrn3IWec+abwTzPRSnxtsXbUxuTF48o8T4wHbRVoYMC0A==
//pragma protect end_key_block
//pragma protect digest_block
BCc5BgxOFhoiNMqhaa64Gwgt5Gk=
//pragma protect end_digest_block
//pragma protect data_block
rYkhHKPm8xd06hSAk+COFa8nN36XIrrdHrfjFz9chps4PSiYp0inTC/Js1YqzqCw
OEuftb5Qz9e/81cSe6dO7duejeph7LGHuYJb/FeLKOnrWLyY26keg2l9YODkc5Pr
R+fXlBD53sVoP2yVJiBDTLj7/sjgRcxw/7S3oE3sskxQlanvhiUwWWgOAYCWMuzy
v7o7voOQ9TgWIuhR7gerZWe2zl8kSb6YxtLn6Hw+mN1ZPRxmivdofNoLsFSsiqTm
hw/yef+Qi2Saci7aTfAkCfArQB//jLSrXxJsUucThnzq3H/1iSV5eGH7LWluZYww
OqULJKHXHgc6Zqr84idxg7Sk+jjJ84lou+lzOS1NAks+N7piigosTpU4opJvVnYg
3wVLmzDnQnwsbyC/2dvJXfKDGoaNwtUFDyW04pmzYp6TpnhNRd/Gb72kmAUFT4/I
iPuA0skKm3zB1yijD7qloTNCFo6+NOrZrANpjjkAgfM7EhTfMZsje5M9aXRzK6kY
vje3AK3t0jPbTVm72SpGpgGmYMQq+6xjUMoJY9ogs4djz6vHPW2LUVeUlk0nmHrR

//pragma protect end_data_block
//pragma protect digest_block
UNFIdAi40/SkaShzTy/UvxS0B+0=
//pragma protect end_digest_block
//pragma protect end_protected
        
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
l5sNQQii/ziFqtjOnhVDQT+drOC2voWfFeM3S2LDAjwzsyWwOm6eGich9IOBXZ3u
sFB0D6VEPQeDg3qTWy+ykDOSAdTt9DQtj28VEiCKmdZ0tYLKMQfID6tk/1C89i2D
1AnUahDjS7RWkNydodGSJRduxiNbTmSI4CY1N/qzdsI5UjbtpVl4XA==
//pragma protect end_key_block
//pragma protect digest_block
Kc05DWAYYwKttXDQyoOSY9nsSXQ=
//pragma protect end_digest_block
//pragma protect data_block
YJZwuvvyx8tdBExX6qX+KJ0/G7UMTqOelDlZBpZzXZ1GQJN2GacxEKfgK1lhVh2T
XSjl2SLz0hSDHhH1w1DNnYpFzVz8KgnAUU8u7s/jY7iTRNPRpH6ge4xyebcuG1Ka
dQey2GvrX91AWJb6asWy58Jj+GXBN4RmBn7SZkEfK5XLl7ElmzA0Zc/YppeGel2B
DwE9jk3YxcoObnTqNM+kYdMtbgrnE7Os3k6GIrW2AoWW0c5aJeAKD2lyKA1U2btt
QFXxjyg8FCLuEe50P1+xfVcoM/nzXnwceQ195ySlXEFLQ+wHfrNPH0qsHCMRwxD6
EgRFAJdCmac3/5mvDiiCLK3HywTTUYJaUjqFZzoqe/IkOSCB1b901LVZRnAnSMsb
a90O15ggx3LkA8kk0VWiupSqwbZBT8Z2A5dZvr42EIHKOECsmLIivJQ4W809g0UC
7hhdmIA5AfNKAjQKPowyJbRCcKzYE6sXWWSLLN+u8p8HQPr2/MBGXp1vYoHOfE4Q
AKBDdVCxpHRUDxJher6cEOiOqRPWJkEnqWRbYcz0UGeIORFdi12R/SHNY3nEj5In
O+ImyBxFe5n20vagMVk7lVwtiHeXWGvGFbzzuI3hnoia2RARxPHuQiR7n/zJs6qo
8hkj2jDkIx75oZGma2YJWBGyomE35aKb+p0MfQ8LezVujkr02h8BloV/shJWO7ZT
FMfGFa/K2ZP8Pgjf3EftyCI4u4XnLdSlWWwjYZI+zZoxYzZD6SktY+MiGCQ1/QdB
JxSuniA4du+XucYnggEq0N8N8qMs/xGeQDoyaJKQuLMl9+pWsmGe4fmVN1DjLZEw
tqunK4w9aSPZRXO1dKeoxq0LR44sYdhvKRXViDEUTzBdjQVVG8Slfah+ZP5bDOef
ooOKGLLYHNbgt3DFFN/kq/WZK+LdZLsQAL86zxwjbB2DjyWiOtQjYDIWcsxu/O9d
VAhFdMEbd3Eg9UwU5SY0kc4ZeKBeOMdXbE3EMNmzS/Xk7HWOgzWwALJQ9wN3jrt4
UcTpiCQYkHwm2apRJO2h3+/BNjqy0Rs93EK+rUkct2rIYtro6pjZsC3VEJFIok6G
eaMm3rotjrhBT9hXp+uuma81HVEdoXyte/scOEFBSSQTDmuvOn2zcMioCxNCAgA3
DeWfOvP8cUKCapR86tpTBrlzzrfFS0eTxjEe9TJ4TAyrIz+RyOpQ133s1JfSGcmS
niYQcDeBlpz0K6I/HYV7mPapZ9VLqDAAVYgEZn7VXAMxmpTflPEaAbrFO4H7AKoY
P81LXAz0khfu8Lhs/LzNXHLS/qyrlGlOIQgeJIAWNf8F6pjrk1FWd6/3gFSM0j17
nhuP+YVAEd8/n7hw3DIPnY8bRnKpsJ2PjS5zblUGv3OrE9he9KWiZuKnmbaQIwKb
GLrOqgAGnWOiPl6MTS9mYTLbAcQKZItOIBxJyM9l4Sp74S3MepXOs5azQHgqI+dj
NMBT6Q5m3+Qroa00eboczehs7+3zFSVV7VG4pxJS0+KHz0LdbLof9FyIN7Bjx8We
hDd5dcqFFaLIssWtY7hCoomM1KFqMEoGIMA2u/cmujBO1fl2275wGKaZEyh6qmkK
N7Lq45g9UdzoviT22PyfUZMrSQ9hBr+n3xgIKtSRU3lFt3VY/rfstjx+6oluIpIF
YpMpMF6M5DljYfKRjVY9qbcUzQZoiC/OF2C7+Bxnx4DaX0cUl0628kcYRAUuG763
SG2ElBxa9f+8bI8UOlxt5iZangQgEPGaZTOkQ+Tnv8sV49msLFMBlrbRsdWdXX1T
mrJp1Rs0zeVQvLyQDo1a9vi1DZJlSRep8QI4eKLvI1eWs7tIqkt5vbZGxqHdqb2E
7NVDbG1Q+17/yraxfcjuQBMQdSd5HmKvN6AY68iT3PnXNQVnujrsQr6fUvfux9vK
fVeZANIJMjUylgUdCqoLzSyA4Vj0K4gFIUVue4JylucBJWdb8iQL5htkwnhWCnfO
OXdgLsIYxdcCc3a1e1zK0Ix8pQupvTpr9iZ2mO9vb3vi29cZSfQLJ+JggmIbY2R4
1kCsMShEteMrfC8PTTBI4czbgnwiRNmaSKgYeL7/Zzaj+9Ea24s0+AfF6MBpVWUb
/zecGrqpdry3pvmUDUO2zpa8pe84+dDcrCH9UUwx/1JUACNdfrwh5G5PMj8rOojM
7uRZ1sEsJtZpyjUODyoG9cCop4o77c9ky6fmOtR/ze2sw2SxuMIPtJx3ZUJKbhQ3
OkHYR2LRZ2VViFlV2LOqk+qI9PuQbekVbMaCypbDcPWbL5LFKrpZnl6FErJwIeBo
zazvPkRIS1jtwq3kDIttjTklyJ2GWMXMSd1VhKcqE/ZemLxsGqUF783QJG/+1aAa
fczuI4bpOt8jm+QRqNDz9TNKIdFt6RHl7dU90HUW3jId2r7a1EfBXAW46xm4kBKS
qnzHIAFXzDL12vHsabBN4xdR090MyRkxpTuqk85ciIJWyUShsmQ9xnjGJKgC6c3e
hDT67UeNvjuMiwKbeJGYfPW9wbQtKoWIsuHb3QnxOm2HCZ4/nCUaPL69q49lMF3V
9j4Nw0RTV39J47aRJikIjyFtyAsz1yfnpKiA7RepAEfnE+GL44JVkz6F8fRKBRJC
vsmNcarMd9yYwCCJD0GcRcsvweB3NJoFjn8lzpi/XNcAD5exoyclCFXxVY/8g7qr
2jUx6lmggpFHR3phHhs/TopRVHgufupjSSspuqEod+O8H8KBeQT8cH/40qilSgw/
Mkvs6STqhFIRN0OiPMJHNXGOxgaGMl3tulJpu7OhR2+Rph4VM0PmTY5KLJfhnUgE
Yu1nc7NpRrb1pAhCuQaYPuhyrcdZ/IJRdMj5AexjQ+mjuUTlq6eF7bIMzVPR7Ji6
k7uXrdB6TgA+7G/9PVOPuTJuFZ8h0JH1fbLCUUFnKW0Luqi0BJtbT7dYVmn5eYhe
10dXvsrPsVGsyyEYJmEKguOEPW0GgmuRYYOjqmEWuy3FsrzhRy/2dBGxuCE283YS
kJOiubWNqCGN5Y/LzhNKah1BSvg8edIwnd4nCWSUj+kGBsVW3hn+/faeGdhG66c6
+7mUnvKd2JODiMOpSYB5Iz6XZ3HehOjG6MlilYUmzRtvJBRjNbp8VsqHOvM8n/A3
SsInsMwjPsJIMCTOwhcv/hlsUEPhXFaoJMyK9EJWtADyFrNH9kygfTV+JdUA9jBd
jzwrZeitSbtLWSwEkWMqksQpjuHHurO6WqxbHYIJI5NVLauXBkRWqS0q9Rmf+REU
onG5U44YYHs0/iHBm3B/syFXM1hZg7pyLR6HDBzcTo6IvrcYPEwGavb3dBo/U6r6
Xf9Aex+Q7XWhoZ/hLjD/1suOTdn/9L/v9H7tEwUrmitvG4xSyqO/adYQpBFzdU3Q
nscsZBRbDK//Deqg8Tx1AdjODAi42j2oe9XteuPRESIBiMZAkTb77IuGvDMLsn8W
psvFFO9VmVp9Gqk43SZY2cRy+7ox1cJLlj371O1eG24e6tmOsPwV82vYzFxbz7R0
MeIN59OStsittYIUSq1iK3InBf7w8eWpWMVCH8LP/RQW/CA4fil8ZgS6aXtV32r0
hb3ZSpr+OuMW6Q91EblY1G49asceoGx8uGClRHXwFp5Cw5AR8u1gELR0DfIkVy2p
myyU05xBzROkJbwUNP7jXRmVyCSEllgJxnSHGzplcHpqedHSKHPshEN7d9J5FgUa
jglyfemM+3W6bJpRy7vA7WerR2MgwwQ+NGylI1XJpKyq/9nOAqNq83BHkoW+Ez+I
plCq3/Ve/E5EWgXhxOwcWUxQ3R6N853uaWWt/vuPlKPl/2YzC3CFpuRSeESsKITO
NpHvEQ1FzvstgS7WZTKAAK3WToac3L44gldoeeHlj9MO6uH5c/h2O7Y6l6QH2anm
3tMgwv398+TdrJZzmS2mffYIAYpvtEcncANMI4SZcAZN8l1IRmg7Q0xzHyLKsx4A
jqelw/zF5RdFfDFbRXB61JONZnobKl7MCxe+al1B6+mtmrVGFXoTO/90bx5T6V6T
9PjKNnCy2/n/SQrx7OkTuY4cgyZK+IjgTmC8u1VZWfEvmB/PNz9FUuZryru5Ts4c
AGNPgj4gZPRV9GLWJ3RCsGuOZaFtm4yCuNiZpfDHh7sBr5o/XX4haZZMMrrSlJcq
lXDr4ZXzJFmctGJJwnTvZfEc8/D3VLzDZ/M8nmKJXCN64H5yRA6Ke1fez01Scbs4
xUmpHLaIx/9Tazattq39ybmlW2jyeL/nKH9KWtb5FJ50w4VvIuBItPHv+B274tcd
4BIEvDDKfGm5K9u3R4sByOOoqfDyN192ijS324Cm9dC3Yy97OmLFIHZtglMQfsfd
I5w7ZEmvLlthl1j9zb4UhUlKKNQGMvFEKVzAxHAMCtKnr5Uk1XOI4yo4nWeQd9ff
9vXfEGWbzaCbj/4etnQF93RDOOTy46tdEZ0XQlC3XK9GCmZDRaWUbV0fP10PxuBG
AP7wrDQGXzOvCXt+J/dAHtHRcZ+xFTmQLPtBVWUbnqQrM3CosrOuPXJ9mLtC/S2O
vkoY6902b0IxaO12wLsAk5fmQs03OC7Y/RtiiRMvcQjm5t/YSR957Sf2dfSSB1Ht
THhvA/4qzpb6+LzgwZQmm3QNKJ1Y6WprIzGxV+jF/9hhkaMb0RwKn2MsfTNqqbXc
ciqWJ71RLEmWoGWWs4DxE4jnrLUYrKyt+fEpyk/qQsa2USzoCsETYOZ7rdCrpH0z
GpDVCnuKnDk/wUA7YMwCBCIcmt21dChxd/14R1/j26SBgNcl6FDLudCkfCFq+hKF
8cgv5pAdr1EOK1LifCnDlUtWt4sQ1/65DUX0pEnPp7XK8IDopTkOai97EEgoTjMj
ckFAmgTt3s1SFMOFV5VKke0YrjpVfDNzzrlot0y1xM3mMaqocPuvyZ2fenq3T7bM
vwuLYmue21Wf6RVy9A+A3Ik+oY6KH/VnFMS5gKXj0pDw82w9iOxbyfsnGCFy/Okd
7haqYWsW8bJPFj+mpDbgnDVP1nXA0loSdbJKPx8r/TXzeY/MOQhn1eoEzIVjKzTq
u444vo9gTg+MuiiS5sFw4nzrVOTsIDFb4yvIVt51QCVOm+TVDYF4RHB0mJxbAu5G
CJVjIog1PFCLb3zyr0ctyBQNmeNOVIAoTwDltCXcIHZN54NdgS1WwtmPWgH/huAX
YakUJMgGvWrqw3nA2tt24wii/ndxUoCQOeaf1D93adyH6htzIhlbgzc+SAiKy8n+
K8q5vDHZ9Vn45JmieMsx5uDMHP6r8NT1LamqhfywvvvFBs6MT3A7tMYJWEOlJ5dl
L+GisTesnXyQpDwZJwcaodOK+pvH/wQJx4z1bHdQq6d2KRZtso2xSkQxvtjZPx7X
aSUUHcuvUCGI9vBFr/wHFkhTfEMUWMxAP8R+Ru6e6CpB8Vojs7WEEgA64LQnqAnl
na6SnDDPNKOvML79li6WSyYhabcsRo88TIRaJAjR7tAtho1EkV73PnVYZy7Q68fs
RTrIH9b4OoRk/YrnWnVd+wtdNkWpS8PSxp5Q6h3rFC1wpkeYvwi3nEtXxI3VrH/V
iZE8FxiNQasiailRmKBHr92vMOdk5lVP3nwEgnNEZ6Eh/jw2ru29yk9kqUt2iRdy
9weEZ4Y7nEojueKwMqc888E7zbruDl3oXkJq2eMVNIJfRtHtJhjYRm2qB92hGNAd
GH9x74Gw/83R5XUvFU8dbCSvhXnqhnGkU1Xcq3O1YXgsv80xrVXuiHsZDGYBgoCN
2l8Id+mrDXesFKlxnd92bcVyLot5mrj3MCLvH3p7tmwbyn38oY/j//etdnHePBt8
HQVHrNxxthLhgtuzuw9yd7MUomgzTUqRt+z+8pQLaqQl6AcejUT4E4elMRqyNsg0
7CrsUWJduZeQMnukXdFRsa9XYdq4JQnOVOD+87MZs8PiRSK4YTByOcebbQDsD2u3
g80RFXSgz9mYuyt4WU26d5jWwjN78r56mTtNZ23STc8qeqT62sT6c4KjetH33GYs
EBHLqToM19GOmowG/NcyppvGo75Fc5F68uWPQV+v26kYGjQToTs91U27UMD/RCBB
ZedGy4kVs3hjKx+Tb2uaCAnyfQ78dpv7cr/WapMFuUpIBnUOGDIXuKGD6g0ZjawV
brvt5vkWkeHf7HpVkAm7P28JXqUWn80CfsxsOB05SFD0rcH4GfATdsWg3RJ33LSu
cCyoIFZPT/pX3oX4192aNQy6L3QWWnGVJax+pDK8hqiXqE0naxLrg95aN2hUBBCS
Vdd+tEz26jaAGh6id2+H4EI2hyjI7niJpfwhpC46geWRXQ4MY3TfFhSYeLAtIkNY
uNrVaJpMp9jyu74WGZ7zlI/ODD/ABE3sy5n/HxkZZ44gMDxUFUwstqIJdkdGzQXt
4oW2N8DGvVzzl5VBUPjzdvm1IrLLpDmkNFjeki7pwvQgGFqVnotxHS54hn2AgY3W
4SdExcABY9a4JRNej133vjLPnAsi/9JJBEv3e9DRNZpuCYqOFODXDqhiEG1ZNwUc
JdvJKwqbBlFCKljhWlZJhg==
//pragma protect end_data_block
//pragma protect digest_block
WxDHG5HNtdL4+u9Q7zLEK+kknGE=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8aY+TcTsjtcCMvCGngr7Jg2u+fbw7MUjZcCxBfKrkz/RXTeaVmvZhmswu5sMwP+6
IQWd7qTjWsEh5KizM5diRqqHuYJpTjQCWTA7UTxjygPSeoBfHD7mql2T+O4sfwXC
DZKPLIShu9si6fasshYO/oVsn3C/04yte4jPlHxxLv+kuW3MU1gcrQ==
//pragma protect end_key_block
//pragma protect digest_block
7HjpBiUzIkwXgXSZUD9c1UZQJ1g=
//pragma protect end_digest_block
//pragma protect data_block
Xk4VYDmAPb3wYYHYf5fhBqittsnJ+YqreOdd3tS61+itfniLjdSRX8zRuGOVLZ2D
3CWvnqUMSDmcxxLsiJhdfduJ2kJyK1gMlyV/VQAgonc8Bq+yLU1ICuD9Ue5xjqvT
ENOhtNsq2yygxSsQ+It84ZtbVTGFCRpWNElF+0RSU+Ld58wYjXLvcefCyfAq96Ou
EyH94eEfW/Dd2aLCJKbyJBGreY63Sm3UxhgBfin5g3D8/moDELCCXtWrDo4QnFjN
7Opq0AHKKMJ0Urvq1YCA/jfvylHSeP1XGbcF3GTEvNedoEYaMqHDgM/s0CVU+fns
rHzjDC0d6ZItRZ5y8OyVQmQ2/VxdeOPKyH5wEe9EiWgng4jIQkMFy/n/Ik+akdzt
Hpt4Al+iO2deoVzPu+m7loC2vL1jnorhL2OVEB72oxcKQzkqwEMa4+FJhyfPk38i
vQdyi/oPKUbJlAyXKDUx2xDMh5oMoaQ/ZSgTb0U0Bs9bd+rS8yohpkDYw4HBIs2E
X5abuyeujObS635CYpRrUg==
//pragma protect end_data_block
//pragma protect digest_block
6FNhbGOOF8XJZ8hYjwOI6b3KiD4=
//pragma protect end_digest_block
//pragma protect end_protected
      
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
L2f9hSdpHXk/UHV2pzI89akpzQgJdzLkxVoF06zyjEQSfk5nzqLrlqmg7tVfvQLj
z4AYT27+depeZsOEjvEoyxhZKYmNDdivNh7JNUdmTsu2+JUiptYdOyQvwpskXwyf
FkxiLVnVnAJiQfDFQmkXiGX9vXegItyoccDFla053q2XL0mrNdQ3MQ==
//pragma protect end_key_block
//pragma protect digest_block
XzUqc027UWUwEO2EhBUpa175gPI=
//pragma protect end_digest_block
//pragma protect data_block
SWIbU5MBWjPfadzCBB7FlOPADmn57OoyHsshy450nQko9vguzDyLLXp00tJ2RwR+
ymSeWslXfheUoKh7EU+PtpdMafl/dIAUWtAjA92ewDR6eOGpra7+wk1MYxIJ2Ti9
oETCwOENtcVIfhgwvKvYnOhHpMrATFKpfw7U7AezPVLNIB5r37Ff4QcwTCN5OHfb
PMmjYn+a3Q/pou5ZAw0UY33wg7j3+vuoZcurqYmsuQzI2QpSLjUOFwqBR+1ciILc
osuWDdgJUhpdC5nhc5ny7Zj7wBFxX6/2d6dJSD1oQ3t60OrXq4JT3wTYbeX4ojLD
0eDy8LmqJWqsTL2hadpMHTRPOCJZAKLHnlmoSYKNfkwvxZwnLA5OmLpVOUR8jEYD
i3UYmruvTMmMsjNvoo3i+Q876uhLtNHdW+pGWPujmJJbdouNlhNfUMCtnIMizTC1
3xHJcgrpeyPwCQ0XL77InXzTQW1o9OEi+g2kIRxLeTLTRjrAz42396+aEgNpTheW
8SB419nakHh79N7p6Ny9XqHlaezIO92xxM/WMdw7lCpdzFqpUbtnGKw8RMy/m7Rn
Jq96luaDJ63qPhph80FZSC9Yasa07ScvSiwC+D2gdTnizJ6v/7hMILxnQsb+O95Z
bkSALv/WpzXMMmUjd2VRJkpqpRkGtMWol/rR5DDsX17kJMbRcWgwCRMTn2nYXZ2U
2nglx4TA9xTRDfMTHGEiJuydVW2RdFx35gfWDhPbbObbyyDI/R06xJxlkd+h2Pvl
ifAPl/VkYK7GCHx8JeHHCUdDZJODeAeIL/f5/qzZ2h/FAlRUyXyTP9cSXiDqFNnC
scEZifN9KpvdqFHdXKSF0M3Qj4c7KNCrBh83at/wn1xt2sQNcbWE9tTL6OPgaPuM
w4dAV6kYgeEaHQXV3zDRYUL0zmURi5/nBrtjyb+xpIsF//gNXCPEEPj21NVwIMsH
R9240p/E/hIDURx18QcWrAFVQwccWWAW8QNDUtXDOnBNHSjTU6SdnjhyYjTE4rYw
r2jwlIGbAQFCyTqCP2hd/Je6sZKh17WB9P+woJIJQ57oa8Xz9JhhQMqKRGYsuHks
enwCj9/Z8kssjCbqW/BDpzQ84G1LLyW/YvdkoLqTIlLlh0dL9kJ3hSsJBNm9ekwR
BToa0h+nBglJiBfT2IBKwYlXHvxyqsnD8OXgB1+RKhJ6ubTgtKKmE/hS6Pkrqukd
h2+oVvshA9uYXc+W1eZLXwU71epZvCvqsTwG5yq62tudXYMtsH1zhSBfknnPmis9
XJ2Z9DaAAXriegHyk/Gx5oxDZvDSJtKecCUPZ0437hV2t8Pjikqjmqf3MWuxGxIk
VYbhGM6c87J+g+QRoIUojTqYZczy6Ddh/VTB4qEflQVoyCfDYTewF6Vjqv6uviZL
sfCwKFl1N8CZMEAfbQojNtpm/bsfyFDRHtNr69DQ+5wM0Ahw3n0V0yYe4CU18OXu
FN8ZO8ril1Dlvexd2ZrNCOX9Qn9T62mYYaP/afx4c7HqobDh3U0TfycGdwAD32EP
EZ2I5lwkiFQkfxUH5eDI2h3ZcfF65a/WB5Ss10MXStM1yAOplP2qhcyfYgsTrA4R
pp/UXcCNrAyGEvoluOE/Dj64BgZbm/vYC2eTCKWHcS37jltm8KUiB5zrIwjsYb5a
jjH+nAkfqTiZ6UH7ug5E6BnTmSBPDLDWx48z7GBEJIVK/c6HyH0BF8R7c2NCcBdF
yXbjkRF3RkVziFLWkEj2I0uvUfzfuyrWAcu0JGIkCdrNgZ3RZv+T6hi0VCJO4K8U
ZMsf73HvoRwvlKfGhv4Y2z1a8NXB3J5u+Eib4MS8Rj1T5Ww1cQxkwlZJ4Din+Gmb
2dfLLLgVB57O4YkN1W7Vm/aB3e6/rr4MHU9AjNe0FI4LGvhBuO9a4SCFvWKyRHuf
z4Ec/sT5bNTdVD6LucI4OMA5Ooc+6ZdwLrf3vJAji8EY1Ce5sJYZ3ZCtn3ofBLSv
IzPwpicveuZoQ6W3xpQRmHrNTAVY354IHWjG6FZIKYFnh1TlLc3cZhx0zEfZfk4E
St0Djzbu7mkQNjMfA3lGq2AS9F3QF7xHhrxIImoqM6XoqM81xB5wy31DEoVHSy67
2VeApJ+Drw1UjQ6zkbH+neSTtrSgCH7Cs6YWieElnZJe99wa3QzmxRVR6OPmgnBJ
7fgd+GBtWKqZZtN9zqZjKUtmnqUs7G9OP/QoDRrJlHZiICAvtVjAWfQ4NGzHnmFl
CiCJRtpGgQB0DDbyVzP5iq/h4trS1oblbmuR/liOgGwpX4+BX1rQqbd4it9W7fiN
87j77efBqDWTe0YFBSVe7SrklbXayh6JbID3SQ2oufvrmIc+V5fMRdsvvLeoIedk
k3PMtouHYUQL0X2Y1gX1KpBqTXXPoX07X07u17oU4yADgs5HzhSdxtgdS/g3Obag
hJeoKmRwTKSiJgAswksuvaB+aokcEwgH7Fg9kVVoc/7TU0/ZqYHJV6FV9SwOk89n
vTaMBxVBh3aswpdlTpQ2zEzD53nGgz5yxfJ16wYTcVd0OdqMtfkDcPhp+V6D3wjM
5nXiFGXa3CuXdCvgb5DHvIWjd9eJRv2bnjJQ3sUDgZ9bYyhMAba2XpjkXbwwE+0j
7DlGQ/6Qkk0F8Mi6R6Q83bECPgACZAhX4govFBwuJgqJ51jtX4SgA5Ahcd0mBRYE
X86Q0GKjEXePDN0xGiEA5H5ptOO2tWYjOFfmX6LncQWWK7/5wEPKT/it1yJxBxTh
7cO6x7zSGc03fQyNfxRjp2W5nQhPwdjTigjOKt/N2XUVNrCW0VfitjiEn/n5D3wB
2QkFmY3/mPWAK9JfSpQlhRsjyEtUTmXxrj9c+uQnGFcXewJcPeMUjEo9vPDoBMQ8
ljXk9T/+fu+jV06qgU8l9NP4ukXhF3vLCqn5G3gBWxbZyZm2XlNf7zUJENdKsEMf
LbjS9aRKsXNsb9xqwRZGMwo2ofjVqMYw86D9OYfl7zIySw2w6aLukvSzKjhuKu4m
58DYudl1nKEykZFSMIe+1voHoyi3HoBh8N8nZWVNihEiulNGHX8uIEW4Vr00stks
s581aVvCOTf2SXsr7nzVIsHDK6h8MssvhcJXlrxtOc0QkdP3lY6qJbFrD4Axy6sZ
XM2CI777wmSE9PcVxNG//Xq+BwWeYPbKmyz5b8ooCvRH+iz2ZykrA8MhjrIq2BcP
/4f4fa2klikDXfLsUyjyuD+oQ2/eOIrCsyEIKwdxJv2WaU38lKftcYKSO9eewLQA
E13BKtplmiCKqQh0QUbrLX9/ZPhy7DYsJc30d16YFjhebLN1gO7TXnwRS/JzQB70
PFxB6IxZIjm1AsZSBhl+MlrasS8ZUCQuGNGkIpczIP8Me9g78wXB8Pkg1a7APeHj
pRGlugGDuwY+3B6Q+9ZGOU7orFr7wax0CZUqpTpdTybhdoUVGNWteZhlmg6QoTx2
aZKCjHq7VWgcYwLGMA1bBrgErgNFJ2qmHGT3Q4RhSnyw1GNgvdP0vU3XHxUVL8AD
O/LUhR8IojktEmaopQ86q6Zh6OAY6H5nQWWOu7hXN4JlY6SdasJoR1UGAhZ1OK69
y7o6H9qKBLZjniSfzY54rY9PdEmYcNJ3z2OVCbDKFwxS+J2rZJ4130aUXhUNy8/B
d37sO6Tgo6oWUs4BjECOW8oNMrBv/utOuxULcsN2sBTsLZxqLbjRoiEPh//y56oP
E5iy75zzRXBeC5pBXBDpYE2zCIHnxQlHzNvXuU591zKwrPhR98/8UCr7/jrTsxug
Fe8LOS8cRU85ruZzzxCSIde4Ua1LNvtjD8zu609mg0ZqQp3+6I6h4KEwBbqtogNC
D13Iq6EtyKF/kZnYUwleLcMM13E9JRk9RibMbaavkTeYdyyduYuio5qndEy57gFp
BDkWLS02DAsVttNoGn/bysjIKqMWu/Kt9GDPNRJ+5lkqJYYkCwWksPOT7anp5DzT
vcSaNDEQuQOdgdtQPPViDCn17GFGuvO7gxhs6JLhzvIwtyhm8E8OJKKbyXsB06ed
U4R5w3ned/Kr7IzrDpWu75cyZPaV6SmtG5rwNqcvLYnkLfHedRphYEBrgJb2ypr/
F95SlsLu0b1Cxs4POcMnJlubk74tBtDXZ64U2gl+w2bIzKIS2GwijvK070dyk+kJ
K0uj8j0OXS5ZcpwcEkd/8Vfe2VPPoq852/c7TCdy4yTuYU+u0pydRsXj7LVlOIgy
RSjsko8z3na9mOwQtnbFFja83tyw0BsMbRoE9I6h0vFNDg3peXVn+05FhVRTMlCI
OYtTjf85FEOIpx4I22HMg6drw+CiAgXuqSg2P3Ff/YdBfetIOHRHHM5A/Rdr8f3s
ph4cLKVwDIuyt0FvUPNowyrlo/0weLbY+1Qw2EoiKC4WuseOp2+Gb1nUBFB0Kxig
t66SQX38xQ5flgh7Xj5PwaaNg0mgnxUO1Ro2k4XTBGsoi+xj+mN8OJHfJzcQAiY1
Cbw2H4Uf6+JomCeYvuaWb78guspvMfnyd46OypRS1twu+Bu9anbEiue4r6MtRsLj
bVjvwSKtT+PQl+jqSqUaEx2rKcBr6irwWRXbYiCcW/4VSb7Fp1BLsNOneAMVTJ4a
Rj0P+GSi5U6vJPYwPxKDulzj62ynr2p+IZ0MCeZvsFUYv/Rbsw1Q8gLV39bs5Uot
Mea1vbJKQJCYnALAvhFlAgqpnl7i6gAeo5cAo6N5U++rqQigtK869BaO1ttoU8ud
78JART7oqnQoyNWHAawAsUSLUarfxy0Se1dazX0Ucl5byEGB+6I+zID24tzKNoXL
lIp9svJXGhFekKv00kfo1UXnBoocuvSnKlowXZEhv0bdDDA69XDfLrp0BSS/ylI4
w4fmSKEzKBG2y9eAqBWxjhqvN5HmSb5tGXCchHfZiDrnDaEig8PKCc26FKpt5ZLF
2uEaAUJsAgTMtzUxwOxtTB6Po56xtr4zQdUqWOH9RV1zraq0KUHQSfh8xcyxWbIr
CrOATaoSczmQDb1iwmw2x48/gcRMPhhwFt3LlBcPhzz5hGfz6dOsYm+cZovs6Pjv
YVuIqGiVfS4oTkggNHD3TOva2DB2mRTugPSUpro3JJvj3G7qqRpEQH0CiMAAfKV6
wOUPrW+S1XLHdu15OR0a0V4my6bLb6WZNfCd3+s02JeFvBY/pZ6lOGeFv831wNq9
7TsStwgNuhSEo0BSqddbjF3I2LPXht2+ZwjmvEi39gw4MMxSQ7LwVkKEubPoc3Ei
8DBX6PC/7iGibWC4i0NOeQItUJNXq6iQsbaABjeY7j1F7ZaNjMTEs8jP7dqh48de
9Ncni7xRwFYU+gt7BiVVNnOF9O6wJJQ4kPYaOdZAVRB6zg2cteoETp6y9UHX099A
cBq+DnAkXVcHqj2JDohl0dYKEjIMGrr+saoq69qLYUvYvNN1eAtgiyf96LKyTOjI
RIrCEihV207RUsD3hE/+G52MU6+YN+SarmRdlw3tLV3b4E9ulF/QwBX1JohxG8/F
lp+vzTSFNPI4Rnj/0HH6ooxgNOPbXM8fNLZj3lHJa9QKfp8ynMT35lF/mqhxhhwx
xilKAmPuIfc3bZdDpAcNYi98oFy5hGY3k1E2pHkXUxe67j8IpgepYBc64r7SHj+s
CUWtGTacByMFz1IIvckY3yjApW6YWmYgiB3HYBseU0VhbU8eE8ZMORQWy1r4LSiH
E1fzf6nI2AWCLmfFhcVPHAqaVU4usbiwlXGmWic+VYSzhIPkrWb0KN07gxv5nBbk
wHp15sj+fwbBSrSkt8HpUm4qgD2wdaxNAdNtAe4FJzuAUhOoy7ubWqcDEY6kVq+4
IK0BMVRyrDb2yj9yQUy7Ehac3OtRRZdQakNfiQ6Ba2ozjY+/Sc1i0nJXRkODuIpy
IBl2l5nE+kRQ6NnkgUf/SSrdI1Aa4+3pXklR1oJv07D/nLmlR+5FoUz+eF//xzF7
xSJcPFUU53raFe3VQVjLKZyc2E6eGhhdzXvEM1SGxOKjrI0burdxI21Wv5Zaric4
r2buXtgp2NkpVGMZQgKFkiwnDTLB30P9SkMQvKEfB64P70gQIcYYsYK9BmaNo6u3
C67pTY4UB1j50Vmc/P3VgWBPzLyhIWkjjLjGqG2E5LLKZF6jaKs46gGoO8PMXYn+
+bOAFoMxszT/xVfcgD9zDrXper8Rwdp0T2DRHvrAMIdUH9HRGV9gQY2g20DEbuOO
jGFfYIFhDJMXM8Rke2L7JIaZnX9/Hda3gaGF+9cSADMkRw2Wh1W98TlWXMguILWx
QEizTl31dDHj45MH1/GfpJ+PXsb1zQsjyzuMGxmzu9cA5Ll/QbX3sOj76Ab/jQle
ihfTPXlsn7SH0p1IZQbNF21OzyfQ0oVbCvayR7OJ90sqC/OEqi9SlVRlF9KW7SjW
nIbvFPgumBQReB5YgtEFshr6mYsiEu7Perzq7S+cYjfOF1NwQueCYaZaa/rEC9de
BlL9A4wQ6i6f3RFRWKvhbrjkk1GZ/+7sNYWk+Dn/dvs0IrttT3ljJ3EHoEPApkWx
y2B62jNwgZXT/aV3fZ54iaozhxIGLXh2ZOqMOclWb+RVW68doBE3+qB1UwJAYgv8
JMEkDufn95pK34AxofZKRhfeG9lLhL69XhL/PBavXiSDhoHqxOGijGRwMpfSzZ5W
qOgqnKp4PeJY6x9aUIIihJ09gFYChLsH/KaZma4zUUllKEqforA0H0YabNgS1SMf
+Y2fWYN7NBYCXrQ4gvgy8/DVr1JCLc8W8I+u+5Thl8ce/9kCw6Bm465QkckC+7Of
IicqVSNKoEXNjQ3a6IoU+Up0hhoPOdiSnUoFER9lUHOUfbYHy2lFrd60K8sofS2/
SWb3lHDlpRersUiOhzBQKURyv0kyyT6nlSqRb2n30gYujqyoCLTbc2Etw0wZBU7u
p8katd3wIGd6ChPhMxuY3plNT9iVM9gnVQ/m7UmRmZidUuwBEfF3NWaMiKlK9FSH
uMdwGu+fw8FueLU8YNpmJuxZSNFAMDNMNtutwfV0/h8ehVAVxdd5oZ6ZdZw3uVio
SCv7LgSVxphG0AwPxBUrU4TWbVOgCmtryXZQ0wHYj76v/2iwUIhG21T41TIcWOFM
WX4zqWPqWvZt+ygCUkE3gsV3SK1hFldDN2Ynd79NVA28GDczFgStc9il25QxbSqG
xyu+yC/wI2XFybgCALHQgGT8H7gxINeOR5KrXggSYuWFLyugzfMYGehw68YMyxac
0Z58eO+M1zb97RH6bF61DEGsyLhBLwhaRef0DC1t3thvjEuzRffHkEZeiW3PftPc
yIp0kW8BUmftz0iDajTEyYgt6U3h00KCZ3fVzs2UQ+5X5Bv/dOZb3RMHlisSB1Mk
X0FEeEeaC/xWN+1LQ2+AorX8jdp2wgLP132j6keJ8Ag2qwY2s94NjQNHkOfO2dr0
b9+pnYwyOeF2ndxHkHjtjUlNPRvZ2y5wlpxnDbXWzz944OKJyzyp0qgdqo5566OE
IcnOp4Kk2kDu2QK4KnhmQamHgO8cOBmpGi5UlNJpNjDd6CdtA5fDYKg6RPPt5koY
ozVkLIisAB2q0GIWEAiG6JYfN6TvlXwnxolZYDhl/s8qUtFJLokJo6v2Cyk8Pjny
PsqWY6mMdnvOgeZH3hvSMo32cZ3GmIuenBPJcH1IPxcf9AixQuUhdpaLSH+HgV+4
XWieXgJskedleGfnKYbEBhaZROoi+sYYNo78iAmXOHaMeOtnsN36o4knN7F9a83X
UZuULc8IGrYbdSXyJsLkbIJUf3ei9VdN5RTecyuwP5+2Fxy2D1rcMNRqPjELvmRN
nELtgaMejp2peplUJ80cCaur0OlqwiwzsKuFSuYQCjJBiSRevV/4ql0kNwni4GCD
m7MHL83VE6T9TfjfQiBUQBmXZ1Yf+0shQePiJtLkekGPtn2GKT64qoJWxRPkfxmm
Tp2vzkOKQBI9l0bCHBsUSsN8rE3lYtYFXju8onDltQwJql+ZL3NRtIpHCGCXXAgT
ZQAeCvCdkep5QQQqNjf6EhoZ/EI3uHvkM+l6dk7cwPTda0cBa9Zsi4/UBJf2J80F
56haz66sV9iesL4DV7z+sA6wjw2reGbSaXnjUorle4IDNYeJUEExC0F8Hx9G5/zw
ys04kwIElCgzAGSUeOiIavRZdBKcfb7l/YHKeiBx0DC4HmB/KsiNWFfioiBhBHIq
Pupp5xyaO+mk1aS321JfG9/aQzLNRg1q75pVYLezs1nwN7fk9aEtCDI7BVC3caab
9I320SyXDV+PZmhefyI6b+r4G2emWMECV3KiJesv8R3tspiV6iTa+Dkzrkc1Ornv
5FO3XVrl+vEqfGc90DxIgbnVfC0Szxz/V/JLdQn4qzdRQxHK0KzYkLh0uEdS8E7m
xYFCNf4aqD3lG//WFRSU/brsP/JdJ6+VInhfUHwBFgS610/8F5k6K0U1nB2KWo4N
Ccc7WFf8wmGYWoSaGBVi4CMw3cjAOakSHOnQ99S7W5yWuZZ4l+/j3yvtvxZIIdvD
dlg17R8KT4/TAwUfcY++vMKJaF/DLssMz1eidlf37zgc7pIA0NRXQ4OR1SFI/oFQ
tznD/a1gwk3i4PYE0mVHY/lHozzkqywIjRyFiMHNqurqXaA57oHilp93r6EORQew
BB4G3MxRSBFM+Ea5Wg8F1rYNtkxiC6ifUUdfsTeQIlaZTJsJkylR29jAUSLDghIb
TAYI7YHaSLcstITVKuUxgH2fWlO+tE/vPMIzweoayKI3cIDU4EB4nbDz9Y6b7R+6
P9zrjcbG9/dOYpXKl1qR1HNRcwTJDZW/muEo6eaZSk85s8RwXiGwSNSCBWnKW5ov
HOPRJQtZV0xspoIaKMFMKbQwOsbiUMq8I19HP4nkHICwomkN1MbQb+IAL6JxaVZf
x1G1A019ti7kwghj0MsM3QlYMrTv0Y44iTJJj0F7qTQnwzqFflsfUvHfwqnbC64/
oy3RyOOmiHn+AVDzTkjB6rOo/paqtA18YXrQPUVV/+4k5N6JRqy2yBY3Ts/Ohxcy
sjPZvT2rw9Yj6XBiU7snQwR3LXiBMBiTTlkQajJ8pVtQR358o+zN8Aa8Wrkrick8
fDnlqZIEGw3qKqdXPGbUWPok2QCfsbxa2lTQMZ+HGyerg3cTNDcnRpxbn5sndpXm
NQfWMcijjd0uYTd+4cPxxWZiPFGTaFkQWJJi5LLwDumLgfqd2w1JqZZGtczLz8xI
7nfp+lWE4L4Tn0AdARQwmeKwwGf2DNWJgYPEn+H71TtkrOeuUEm+blnSilh8cVg2
edWL566zGF7bCIdQfqnTVkQTcclHyWv3Gy/cS4kxO5vIJL/QGGdEGWvqNYIOSwNW
zBYqkYMMPLzp6tTw5JqnfQ/0p0qDg/4F5BAIiqfiDeBxn4UaJNlDKSmPL2K/3TKu
RmjNnr23yXROjK8ukWdlXdEivY+faBVyc0+JZo4jcnosYKBlgGE04lrUa8hjG1MH
iKMwpq36fsK6E1UPBNPv1AwHpB+h8EZaK6tkB+CQJ3z8D2dAGHwr5rLowLPTGdKr
ZYeOU0xOC+xLlzEznCYxryF+V0K/3lXJyZr3ii3fG0q5/VtjLmwOSd4X+mrGACls
KIZpTv5tnUn/JUFF9HTfIKNXrocT91KuG4PknT9Z4FcETWfSOXqwnlPCaQGsOrL2
mJuDicSC4Zt59ccp8R5aSCmBtYsVyzVFifG6DgDoi6C+XTn9HEk2A+e/M5oCesPK
2g8B44XbzCvKDODEQ3i3veL25sR6g4kmJQW9jZeBKpkYFfyafBKnMjHQBo85fmeA
MER7Cxcy391YeCsjTfGSl3bsuaR9T9YkJdKgrX84ZY3aWSi6n6h0NmRGCZRP2+CC
AEbdyETMJXKI7x6CAdr7Xa9Ti+0gFaIxwz90E530Dii1ECg5P2KLuXAPAnw+Ub2B
AcFTvtcORDPSGdyQK7woedelbAsMFOBrMoM2Vl1Toe1jni3knZv2XSUPxGdgeodM
7wUtogJeT+ROUSJvWYLBOh9pDoByKv4f7LNKyIpzVaGf5Fi36kjEhpWMXgVGyW1A
lhAWBEi+ehFVgnKQ7xZDQVeVI0c4TwQUSJsaJrBibFdbBrpPAZ7IUSDhJs6Fi/n+
x5hLoSO5Rhk55dCIshoHs4WFdkBLUH44B5wmF376g7hDkG4ZGFhmmWUAgZTZVqnG
RvdJzpbroyg0RWULYrdOfZqCliZGjfzFRaMnyEbSt+ky67IgAyrh3d3si8k/p+5b
xLJYiN5qsOcsiZkCcdgUbSDCDbvyE1pVsV1rnW0suvUL2BEht/z+K5twA7/KeYIe
fdZxB3NHUNfZZpunVEQSB2P16RRSRiLvIViVmS1bpKP9Hqn4I2ERuKutVdqlHP48
j8aavrL7GNQOyHBWQK2mGWL/rc23V8U8RvZf4B0lnd/gXnhGnA+e37jKVxuZQapX
idTnuIJ/jQgGzJ/NRdzc1+/XAZVnj7n+gyLk6/zKp2Jejkzv1uLsBBsBINM7iTdN
qhwbiC9o47RcffK+D794msvlXZJ+ZZWOm5ZVtuKMR39aIILQnWu+0Yg5KAx1bb/q
zY7JXZcFLr6yFthYWvtEFHKUhmpIrs7WmS6ilq9GbJ/59eMJsdEcRzMn/10U5qpV
3N8kXgDhbc+VD/ta+0azD+U2zv8k7uiUa94nt17fVlCq5oTS8lOQDAIxiYiI3KCY
MrC7a4gm/CHsYg/8Cjf2jyv7iahqctsYkIpawkebiRGhcfBRc2gwFmXJEEX95LDt
YQcigyTJ4c5GAyNr3toWOIReeOQr1WShKQN+rTm2+dZ/iKQlOO/Ck10+7YWb58VN
uSIMBuHU20/1/zSwZgng+aZctaUswj3jmfxzEcCoH4EstpTUML5qKdt6RkQar6DT
calXGkG7imJ6x/d8XVpbTRIMIAa3u3OhfP2O/WLSh5jwk205GYZXBtPW4B7v3kVX
t5BtsyJ8TsRVUGKxnbw7yCpOd00bLY82lUSQAVp276a7YkPaLZUk8IRHXAgjlMV7
ekPY5FZeHTb0V+PHS42Gnah2A2OfP7U0PaiibMVbbWgMZFAt5cjFBwup/S9b4PgH
uIYkRPQZzGykwFt7AYYdwUfX8Yd1opOin8TLdlJGWvNkE7vUVPuLjWOcJZLRL9Dm
4/pCpSLbMohhDkLzkuO5dXarIrSn/u4wjxfmlo09CNr3r/FsyaPkG/OscHS73Uhf
IZ9E+YCbOH2LQD42KnHqU5E5Kaa5BbdlNFPViBCIq2iU8R1M7nHX1t5BfB1hvYAC
Q7cpRj0Q0jVerBq3V6vqSkAyaEaRBx1mkD3Hj7AdWPrYy0sv+8hO/SlgAdhiYM2B
LQQ8UISbwp5KETmYhu/HxQYbdOfXVzw3uIiCR9Z17s+w0OqanfB2ohkb/wVv/Sue
rMRcC8k5+Ahdsf3FQC+eW8lTr9PFXYZVoALKNXsQKhv5+3qG/62QfchqUiVmOZga
xLjh1i8Fmt8klViXKB8fMpTGokK4dTqxxGKtSUWIX21l573eX02WN7ps5Ohr6uvb
f2jsHzLkzNZQtbNlXIWv2ABwuL6iuuvVchn6YSaPVKB7sthI1PTn8ioe+O4MjBSG
TuzBsjHsrT4fTkCDofUEk6Ju9xZ0lHcrj2ve/iG0gWTtV/+kKFBNKMCCW56UeNeE
yDwU5wEdcKQxjc6uST4N/AwOFNI0m2rA8B+IFKW43aqo+O9susthvof5nMPuoHFS
GFf7k16lmsQNQ7m46RBAsRssbqGNpT95uqwArY4rnEwsMMqn3wRws9TA2iYIbR7L
TEuR/F7EenMBUeDmqtm8PIjnXom0C47/uACEu8o5d/5Z3feFLNw8OOemEBNe8PjA
f3Ue8fzY5rOwsxGST6tR+rPZjufMPl1KEQ+C+hc1z/2RT2j/QxqT8OKRsFYqsek1
4qhvk74nXY40cLaRnK4dUb406xccvKoBiTf3awSeVYD24EDsAsIrifoIRtq73+Uf
LGbGfE9dggf80lLBqw2SFasL7Xq7Ke5rzbwS3fQnax18SVcGGMZ1s+7FOQd+kqUy
OuVoNYn/iUN7JRtMZHJmyKH8EABiQWa6CD+pmO68xpjD32YJlYyONlSCLMXEJCJm
5zkU94yauRuNw3ShIXNXX17ATTZYKEbCWSnEf8145LksDPjWE0wWw+7S+1oc8tPk
swWV0WPmAYUvT3uUoG+OFf3NDs/eTKnsOK3TjYkfLng8AdCd0mEP0G8TuYQa+jjI
p2Di0vaOLFlXKV0cVixenBvobb39H7y/XsjzhB3bQPiITkdCcuJbj8zUiD/MihXs
mCbj9yPuPiTPal5B5+u8tRmcF66fkRS0X51mijYIyAIzaNo1EGwGrhc8j+yNdXfA
J+AANQLxPoi2JokPo0TKuoz+I1sK+p/3vXIIqvrIlySckZy8Qg3jsywMO/HIZRMr
rUJSWxTJaGz+lmB9gnWaWQ9O8OvZ4HbY1bQN70PGebFRxRi3PDzukes0jYQdq1SS
t567CEKmXdJ4VstHVacaENCIW+ewA9ATphxVeAgoFlwd9MOsKthGt1JHrNhA/8zR
zwA1C7RRXs8u07KYsAzXg4C9zUaOhvlSN3JgYhyTqqTwVv6oxy2ZpvoG/0PLVthD
MlA/4XXMxTwwGyuYO1UbMU4zUXEkP3r3+qvV2COIn3ditu4cWkLAZ4D85hLAiFlJ
pSG4yTOjVUuq+ALBgDSFab48rkvOPpLlR+Wn+F7FiQXSz0NTUTd+mcmrS7HEewfL
gPeqXjgOW6am5LSzIHEXz6Fo57Gyeu/oMxiaerjbYGm+ZaW5oFYLCRuJNGzp/4EL
s4nagnD2QnfGfQyQXo3YDofCgyzyD5LZK+wxRbqR2bgSLkmdpgIG5Xi11yOjJNXP
uxshqz0pnGQd63+X4t+DTJEX83Jm7+IAoxY800e93BC9EzZ+VLhI9g9K4MQMO+P+
7AVa521EEsJEuIc7SO/Xdi0r54aBfwanpZaD4ebPjRtBxK/9uBdfRFgfSJWHLJTK
UuIgBX2AgUAst+ONQYJEcZp3TX8Lp0n83c7dXotdEGSXqRFJa8IipMJQeP+ZULrm
3m770I6ancUQfqcZR0U9dZslVzTjKO4GTWwiMuQY/EwTEykxwxQ74PjDNa9UWsdZ
5NolxMGkznorpFcNUh+OT8rwfFEqEg6I30gm5bmXvABhgvOAottFgG1hHl70WAem
AhfQPqj0Px6mmdafB3W1u2N3Om8SB7XHEpkz1Xs5/Ic1ShQeXyJA+eJyCEdeZCSi
wIk4fZ+yq05WShbuKD001s98Z+JXaXL2Ghav+Rkbk/aQes8LMxbpj7M9oHMN04o8
lU2H49bAM1aIPqHIhakaeGJQXEhYdYaH71pg8dMKe/y0R2xIn1JqhB/17rNIhqNW
Idj3tsUOQ8/+eWQG1hW3KHdqqB+UUmAO55V6V3frsUnLl2NkOuE6efLn2CF5sV+H
ORv3G62XhVAhFuJFqF66g0hLb0S4PWVXH6anNuCVaTaEA+fwbXKruT7d58DSCLlv
jW5crIEcYE98J/f8xKG1wJvoGTsB8jB7Mr00UEIvMuZ+HRSFW9CEdJ9eujMTzh8q
YXquaeEBze4/nuKbZnqIWA/6M7uFHMBfjWyyHPuog4XKshEOty1dppApzHaixCSU
Uin7SUMNTKP3Flh2S+zy6jl+vAg1bc1j8qvSBXM3seuMwjUTV4Ums29oYnIj9CW1
0BOYMnVKZXC4GAWdDbp8CdKzyeBt9R9yOQRxu2pbdk+FRhoT6XXf/w+0tam//00X
RhjFfdW82ICmjzXOrDsDu6Fyx0If4DMQUe5TebnVUtfjhvemAdK005f1cEIxZXPq
CCp8CTRMRNth3bKCaXcvwkHB9ygu+i1lMV45vOtoMLdDhA9+FIPohDHjhzsX/CID
OrhPrnQYgh7X42EPtuBU2vqFntLUByilQ5pj8v8rKlctbeugoxlGtUPHWSYiTljz
KFJhACCG5JayCRLOSI62A1PvBzmhdA29CIb/VXx2FWdTLwQGnJOvalzeIHwa7rCM
IwfIxR/awo57wQ3Y+0aHOvhNU7HBkLjo0Bd+w9sSMp29dMzqfq+0lScHpkhjmmNN
tKi0dMiSNt0R4S8lLbYY8dpuXgBFSRc+cqLJAvIoUdkbtsqL2Rzd+BqWWbbyTX6t
QPwIrUY3uD4oe0lF7PQcf59ercFBiYsH4lKAnvUWxmV7q3QqiJ8nS4/znObNh2lH
tje05sPeNUaDjIdm2yTfkAMo37uLImEPSMrikcF2GyE56M39uv9Z8by06oj/IbHH
F8PQnZvz3EgKk1IuIcvrGHEV6R4BY7FkX4luBYWSDAtN41hqpBs7430WB5JooIv3
tTlNclZAptENvSdvgDqLV3JcRgkHSm2JW+N2VYYf/9lJl08TiqCX5f/6eirG/2iI
Q7GwLiLRX5A/iuiaGemK5K61hiozxbfVx3klxfcIFPTHu21lV6EeO5FATwmepOyL
WurvnFV5PWoGzwVMQ/fchRoKnmInQHWc0frTq1aRkE77E103ZLXsEKL06YMqwei5
7VpgKMJqsqWLbXPWeGfCZJ/0UCaxYrbFsBYBCrvatBsiAYIHxwN//kqCcWEaga2G
qvpuggV5QVUhU9XDebwgJy9Y3Fp5KIbWtxeWzbYAnUiRCgWeNAcKWCqhwy3fnTnr
SVwiBH40050wf3hQfCFoVyH7XMHlTXcZDldDd85zReXFcT2pjhqmy8lITFRLvzss
E8CShYus5SHNW6+TYGmq9Gey+i+OYXzh7QOiTSEsGJh4qidbBE4Hcgda/Ph7t6io
8mNyQNIMaiKCxbZob3xlzje2XV/ed8VZ09CRBmoHFS5z+QDH6wMZPV8t0ljP7scI
SV6dG8/2bfDobX9Hqn8Lbb3x0zUt8BQ9wqFPauqLksGoJFkx+O5dEOR8j4UwuDHB
y37M0JcR1nzZIypyuyuwkE8nZot2UBG5yBDxck1EjSaMfRSSx1gaGAQFNt06ftG0
5fyXnzj4XlTV1zlPAhA3qDulMtkwJbRA2QRaamaBOvDoGe2tirr2OcR9CmQzgVMi
8AhdYg2aNkU+Vnv1N4zhmbjTM33H5XiWawOC/8hz/rJI48AmISFU9jFw0jowrWhe
XPjkokfHbK5TmCY7/miQdCpE6YjE5j9e8/JHOok3wnUUrSv4jo1M26YmFVHGauKy
kuiFVVaYxdgEJlQeSLrxQ8ZZJE1CxSLFhyR4Fu0rEx4S31gmU8QGqza2xK5rtSgW
e0V0Qfluzqr5rwaEnxkmaoNirjiLFM53frcXGKpeJygr4b1PtK1FmM2rbYebxzsd
cWUHFImT393aI+2CUPh0OaHfgnJ/c4kvch3erKdY+OaKvWy/hc/7Kc9LQ+Gy7pIt
ikBbiwKNbRcnBOazTBPUCbN1dSw07XP5krHcpFINdtSKSsvLLJl/Nf/nAyyX1TsU
K+Nq1Iajgcd8xvrKoYo69zRijwoe9fFVSuTzvGC42VDoBKgvrOESY2NppwHdWdDc
LntbyZMSCYJKSeNrEqUnBKwt7ZTPWV/NOMS36xvoIZeKwVVKmfyIIvdOMKyc6GFx
PKqQLTR0sQK4iOFTVjtZU4iZbhzHptBXmdc7+gr5JnhXHp7g+oEyhMDTAyLildyX
nbqpv1HRkudmNYeorjoYLVZHJDikElsX0NUp+9DOh8sGpJqNcfnawWApLKcnRk4D
b3iXC0sLDJM/+dgfMhd8FwvvPCDdBox2P3ENz9dKpMwaTdh1L1+aJnxoACBB0m0k
wM/H9xxBMNaadC+FBoUwOP982OZRATpyTowtLHSOkKyINE+82WHIG2cd40lJcFQS
0L5wkJhEcz1mkZuVktmZ7nvv96nuR04JUOkwSueQ8FFTKFaZB4uqsY2xmxvDV4EI
ERJ7AalQcYpjFSHSlUN8ln0GEbODuAqr3PB66Yd6QXgRcaxSP2k1PAwZzCBOnc2p
k/lNehJ/KysXRKaA2DuVXGuAg/orIW5QSJnBVpuMx/KNY4Augw5EvE3fN76QAFe8
KQ1OeGpBrdcTqw8PZtQ87I68WE5UUJ2A/W1Kc5E3FntkCcmA4y1UE918DiHqKAy1
MWad7TxgftGddfXt+MuxbtTrXBPmQI41rocg6CRTkXG5ZxlMqpS8q9mPjbjJBSNv
18Bg/H4/6smZE5bHkhsY4Prs/d5hSylv4hppc+bKN+nXM85Z8ViM+6Vh5u2JzJr7
ys7Cq8JoLosOv8+FGDqmeWx5LPTEovF5E708ijzbcYxKnoCeeuhf/OcUQIHH/4Ib
yEiJWNqqI3hCI9IcE8UfLY3CpKacQWLUzR94oW1i2io4M0Bcx+rceyOGLUuKi4YP
w2fVksWuuYikpzu0PQ2IrMP/be5p8p/ggX2kM6DTgROHGU4/wf+KTsysjj2qB20R
iv43Qlmiqd49KR3bbYVwf9T/+BTEyX2XEri5Jj83DcRTpXMY6Y7XmS8eRnayzeak
YlTZ3rTsxzch1Yqaop1nGPcz7HYFGycqalQwQVFeo1Aml2O/BAhAcQZZ88//jQan
tJe+bkia16tUq5uMyXc+HGNbHy7rBKWtAUbcvHVHuE+YBLP/7I9cmxXVwb+2cw9X
8LTE5iQ1AezoXN2WC6Py7URyUKMFGg0u0QMZV3RGQVzLfIg4x57IznEV29gnqgLf
VNplfZNgq89M2LxvcyF5wNAh+XKuC1/25d7A1nO72LQMTFjRwUr+M/m7T+wvpjXK
5zXUh6VzhVrypNXOnzbUpRQyQ9zkqy9Ca/Y01i6ma5VYYFX8Ov8kEDopIK+raaYg
6enhftlpttQ4pwCo+F18o6cyId7Ha6EwIZRFNIGVFRnGbonIT+pUDgTM2pHpfYNW
nzwiTw0zY5zFJnpLst9fsRBtdqI5g/NX4uQWu80lsh1GJ9sPqHSONAC0RpZ2IlQ+
r1ucnvQQzbusrWjWOlsO9KSbm1zM33XqtZr5yNZJNxkp2KYE1PBsY/pb4bXybHxq
Z2sh069wEsXozfm/r/LOqm4MUNQ/Eb5JvmczQ/d3HwPQZxHpOSMmmDSt8Ipmd15m
CHikJWcJo6LRHaGWQe9+iyp+lBSA07Xw9eqjZHGnG9t3OnkFYEtR4Y4coTA3hmCd
McjC43MZRdOuIB3caWGoJOm2AcbMWyhIcVqqL36jb7eI5CSSPP0scRjnYcUIkNH8
uMBO9InqFi8ZlLLxsG6e7jUzGZ85zar6Z4bK1QyfIyMUsWjn0buHCMTKwEzdqBQX
+cdXvamRRE7hFc1IGrjihYRcarB1jBgrPTirkzrN3UR24XomP3vj3aR3/wtTgPHR
MRMEJmkpJ+DkdwS0qr7pIGdansUT3v1jc27ql67xIYueq+EYWFnUEdLwSwedLa8h
NMK00/9XENt9wlSa/P67D7hVTGtFAveptdXgFDEE+Rl/qEhCgeAJ2nMr+deqlP/7
8DWsds40oky0AWHxGVb7K7OU7aq1MZJhE1n5TWsjf39tSP5gcR7p/02TBtVBTitl
SNMXuYq2FmqiCLQk/J/gyTlZ34ih5tQvxozqvVFOYEQsZsxIjrWNiXIbBmVpWz7V
bGrQceLiPBb0RnIiu3KdTBY1YLEELqn2cmdURGvj7xfdsU3PDdKkVz0ByTZ3OGHO
RS0nCNR91/Qf9Jeon0QYhiHoOHSjdf76WXBeB1l6TAt0IrNu3ETppmXxD6trRi4/
w3j5/VQF66b5NeIGazUE+VzwbfSSil+db1SPlCNizjH+RWtjC8gwrgku3bhuXv8M
Goy4TJG4em13qQWhafPnB3M1USc4VLVWdX0FKFl1hDNlw4QpMj85fUAZwQJA0IR2
tdhEhWdg+vQnqIruKff+UIFw/ELXTWVqx8BY8JmvEqpHZintubKBlYiStXCPY/2p
cIDjAfP9Kvx3C1p/NL1i6wcCYdoz9+emrcUtm+R7D+rRwgla5srgBjo46fyHa7i1
7v/qzD3leB0KSBMgqfmFRf/z4VgW71f1xcZ6qaXVXWAjbWe4CGHgK1HVnqUki/qi
Im/cgGCPqGuOpzeEaK/Zufrto7W2dG+T6PxYz8Q7DRmnG0Au4lAniLf1SlFqVZJh
58xczkPsVyWOcJKky2ScmYMeZb3RIitFT6k+D3I1inxQpg32D+uy2LDJc7QFYuV7
LseAAZ+sLfZGcNnHmcgVD/Vm7XVj0C+yqGDPEnGYRQu5Qanmw6NrNUSmpw5zX4oi
gnCW2ofHf+ZF9UFh+XZzLsgfM+yxM8ONT9qFlpbGEHTVin2tS1PUOMxxejmSg7nf
hnPFw8PE9wqd2Dby46r1cGEnWd47xg5+Osl3dg9qV4aryi5kOcYpJLCe1bRqjGpx
OgbmH1iAibK8nJi3MvC25N7CUr9QwWUAfnzvI34XQMBDP0GtwMm1j2S3xAbPsC1Q
shuNH9TDdqwiYF9ro42noUCH7nche3fxlQW6lwCpSxwgAMSTj1EQav567d7d8HZt
w92MWzIrfnIXCgylWV+ke7mS/GbRZZVOTIDnBhusPBhIYtrmUEOXpV7JHusQ1XkV
Mxa9YFUb1jUtXKFNKBpjxw81WKDTgpYT79tXb/481AnuYZRDaZGVaf4tDZrF2XI/
IP8no8uzAHmCxDdmYak+93BBsJWUEUImwz9mPhCCbncjTSJjeupBCNlW0+Fn9lbU
4qNyMcLZwLIZw1a/x2hdCRRJtQmw6tLYJaB3zuZGihzYkZ0w/rTw49kSgf+083Lz
VuNfvlqpegeiCOaD/M6XpuI/YAJqs5308onfg9RtqkQ2aw14cQJyWltGMcmobS8G
+0vuWyjC4WJfV5iJ4QKOz/4ZuPMg4a/6zE4l695lYJxXza4T3BgMIPmsRfJwTUhM
cXbwuSFMZIuaZScphkoysr9gsFwChcrlx6ZS+5XH0TP+qrybF0XPVGnFZkWbe1sQ
498k29IfTPh0ZWYZ2pj4B6PjyR7Q3TDzXJ6QbFJKbl3yBTpM6qEyw7AR1mpbuOCB
RqsjINxm+6Y6+zArCRg1yH8pmqPw5BQdohuLJVzUiZBpGt5DnxosFaRYJWwlqZST
15kZjD0DiFd7j/+EjqHRh0QibeVA8EZZRC5qujF4ZtWV7ZvufiPZAlplnW5h0Z4Z
82NiAOUDur759Kt3jP7F9X26YrJ8EkB8E+5l6cz75DrYne8li0Y38kFXTj4pNsSJ
poQjz/fRNBHxIj1Bz3LK7gHPbl+NL0047DwqTmTlO0Fj11jAOZeHEkGQ+R+hYV3c
A4vZOLwlcpp3Qnsj/6diMeEce02F2yicrbLT6Be+JWeKb/8jABxlzJ5/NhrJBEV6
4dqpY9OtoUDt39MHd7ZfHoPHFXyLb9ql9MfBzijHzx6vMppRSeVo8OOYBN4s9gRO
aylF/aczC9UGcOehSDqeK7pBboA+rb3e8QeQmmFZcXsHSauhTLirQ6yZb7NxC4PK
sbwd5ZpodxTLyhUcPOSQUPDl4GI3T92fZe1nr3aiZ12IP8YHHZ1WwkFJRrzITqli
UWpzNDvPivIRyGTVB8t6tYo46P65OIyj8G/i3mgwjE5TjBaYHyoIjfAsC0MNY/0V
5LXubWc0ia0t5dQNKhHvLM51RTQJz+t5m05qukeH1ps02KjxlPHw5Xui3Dh3uwky
Bx1qU5fNBWej7L59HIeu0ObJTI3cKEF+CLXsAt+ccrfNolC3aaYRIK+dQEV7FD96
/DMTnCdC/pjGzkTFJ+zFQ1bsfJz3qL1rA8sbEZfYryVutnhIpWQkZ0U6jGyNPYTV
Lr/D7qLrQ7qbu9B1ucB+Jsh6ANLkaSRDg7EsAlYM9xpxtJ3KgwozQvDDNyZSiJDH
rf+l5MwrfZfS9FUt8jnJLSWIvuV1CoXvfiJPpvJr2F7p2bLZ+x6lNu6PU0qRbAGp
QL2IYch/dummlYKtt9sUVSCLpnHEh82lKP1YW7XVn2lxslLlo2PcCntYRBgGy7sC
ohbTOu/FCGws+geAbEGJ+Org+09hXTXeqXqj8ztSwSuqziiq2juZfNiyHBQaKuf0
ofpFqi1y/dT8PRVqlTRp0sgVIDOBjrp1wjV01GdOWCAnFVw3hyBB3H8TIa0mvQIg
XcfyDD/GATBNstamucBMiQ5/Gj+z2dduoG4IhRLfdoXbp8ON0u+S0zPzNUHuNZL1
gNRjw1lst0HJs9BhNWqZxRk34LO8maphaWJ2QieEoOTOkPcHvjWJkmp8h2mj8N2N
S1midfk1OmQ/+NEnMbSh373fqL4bvFWEoH2pDDcrn+JitPDq8aFchiB2+oxDXVlp
GUO4hMgV7yRN9MYJI1U0UYaFWqbOiFBjyeQCyK/EDRmguHTl+0cKpi41m3LdoFdn
AAUIt6P4b7ZazG+xkh1mir03cGPw/WVCxKB8FfdJGfALqzbao+7MQSoum2Y12hNr
ht8oiuzCKYTODkAvSZPRhhdjXUMgaBHKXzm6c3xT8mtHGszqGqnAhl1/KSaFsCuW
cTdo6QuQBN12uS3nKygcry3cjn3R/5sTsUlgIIxVaELjlL++RjgL0GtEAKpDgpSY
lO+7pJ0u7bdHt1ldW27QPn3sii97awhuUAmXS7VyaOArtnWMIYF9JMoHCXkcffCB
/fRiHi6PtwzAKCva4t98hQYehyjq71e/PsDI/G8VtUPi4YiubOJ+YeROxUDKMzqo
bvvFfhwNH9QClL0eygDrm4gSQw8Xdovr/vKMXOM5TE7oWh37NjdXXHzfMiMYNwCY
k1BsFM1d5VHWYf/x+JqqHYUN8aY09z0PH54gy5Fpk6ZvBrxeCCVQS2WoZZbXSM1z
HdXluBQkZrLwy8Qbo3PwdpqTAE5FD4aJKLQMwYCi5atzMszTYUu5QHqsovlBrgIA
TcUlepzkhsNuB+sNnR+zcTT+fx266dJ/Z6Tl93elGadclJnEXkbZLjetaM2WbFUe
9ANtISmt0gKvs4QHZWx8u2Q/zBAPlSikJB5hwnhNBXiItwo3XN5OAfKJTxf4cicy
IGajWFPXmmnpwS8p0kGlyUYbGnW3ujygxN80wbd0yEM1Ym2QxZLvXzP7xN4JUFKG
BFeuFULhrsOxIacWiHweRr+h26yMojNAWYZ3mE1+Wjiw4s+GPOAR8nV8P4KeNOY7
OW0lpNdrLf1b8uEKTGKSuCQhXVX3shh6z6PIvVX6SpyrPMgGgIV1D/EqLVyiXJ1N
sAjbNlXStG3yOU0/xrLQAd/+UOKMNt4UW/zkUwOMfxwbwKqvNE42dUgD8D5QBoYy
Q8oKGXrPW+8RINJ2tTUQSMHmSoQoiLEIlb7D09b36u0xpv19g1Xcd5ykWFMtF8Mf
m4cxWueDP/cWRprUDWCkr45eBWuMfXB3d2nFuLtTBHRytOvFHysB5bCV63wfH6FM
4oKWazilFqVDrqCvmpBMSwTEoAq16qWh1kFkbbmpf8/UedpBAEsTTsIsxiRZnXZM
rL34RSLyNIW34Ce1Ow7MlfGpxqKLaAdrjUqlNL2s6gXtD4v7wexXrV13h+gDzBpK
TuEEEVgZuNld2/aYoKiOK4qoEkAlPhxKcRGNMcpRK8XGT3QqgBjyfBxf76hy/RUN
2N+gpc9UCAj+keqQ58HQ1fMuN/4i9IWpOobBiejx5Kst0eyX+est1yJfvuvH3STV
qvqgCcoQ98GMLZE5lzmKzPr7/GIWm0GJ5hoKeMwWTNFSd22EqG+CkR0OgUDeaFYO
NuCq1BJ4JzHF0pxUhPhvemgaM64iOSKkZsHoJyEe+MPEuZbQwyevkcE0OzMNybvX
hoW22sQzOKCcqWUU50Ie2uWSUX9WS151tJ3GBOeee342tzE0Zhvp8qQaQIT+WvG7
fHm78/sBRGQN52gWr2fK+tNshCPEsIVBxxCnfaY/+R0rO8U5WA0kLbM9KXDoPvkx
gF5CN+RkUgdVs2O92cw83cX6RbQX75Ry2dp66cuZc5CWbcHVim1HjsiTibvstYJC
O2mScEusBznqjGku2JqRY8TbbcoKfp6/lR0hdc5PAzXTxQrAiaNRurZj+ipY/iC4
gCwhl1GziUoSq8JmBCCcrT9JlNHiFRrBUxahftxO5Tcq7jARbQ2n0lUeXFAYlVCM
DMP7XBJJvvyLD94MC4vnyBD6LXbAtTckfPPdtcnh5+4YgCkSsDpUarM7TMjaTEh+
pl4G2GaXplOecxq88jyRvt4jn3lIbeozlBgUXosRvFmzOXSKv764SVEb0xpQ1cTS
gBeFQ5AdOOXFimsih1algQkXhFN5+IJ9Lx06Hn4KjbhiKfHnvzd4Y/JkadbYm9SH
e5HJzlUhcGNRGDUqRyZXy3mrBeXJo3reDX4KAlfNmi7Jxi6SVVpEEE0kNkIE3rei
GfMhoFMJZnW46gS1XkOpdLqgIA/U8tETRE53qNNTOTd2zBWHlnPNuzeD6AisB9H+
ZpDqihe+tJ/Q75lf2Guyn7UosX7aeLkNCsTXBojDpmtUGBaP4uu/fd5xKHiee9Zm
sh4s+xDgqQptiKhOaqlXeiJ5v676efQKvt4lGxBVfTrntHcjq4Jxoc1SDBsQBL7A
1LLbTUrqfNn8mlrpgqr4FWvsBwpswkRzFbMCft3LRTv8yThxV+E4nh2bCeL0qF91
x0d08LKbCzu9YTSh21LULqrlgF7W3OiZFJUFCwW0Lgi0GPuUxJ8+4SB2Gv2swRKj
+eu1iQQCCydfNUusHNTtTfScD7WyBmGMJ1DKcUr/qNsCiFOoYjdh7/jdINwtJ8Qn
l4c85a9+DcyN9mAUdnp+eH8yULgabQKmweXsOSoLpCryQ9QONWTAb67/Zyfm5UmR
3ZHD88MapwySItIf1VYe2KRzQGjvnLB6L8CbCAeow2w1QnphkfeH7yD6+8+XpDUq
x3xjrQr4O1IzIU9MEHpb6FNinKnY+oj6aAH03QA7XTgdLCc86AFCFHMA7fgFSRvW
UrpYee6pQIkEeWsiG+/JlMCL//YLuh8gSxhr2MPvbB19OARnC4wPiEPBi3B9vPwc
ASFblTDo+1b66e8UVgyDH6nQCC0OUSM5VdQM8FPH/gEsy3gCNS+2mzMq1tq97m3f
C2gNsyL6+mqF/0XFlu9MyL3sy+8N5ycAKfygzXo+YNQ5UNoEHU7ky/1BhS10jRyn
Ndo/zS7T+UO4/KQAzuZJjhLKfPcg7YoAmoLEr2Zpbz5ijRJw9yKycPQlXp+IJGTm
1AMvCFDt4UcuzpsQsHIfZSXNODrqINTJkBzMiNlEbw0N3PJINXY7mpX1qx2FweLP
sM0MyMUDokUTWTHDO9RbD6AQcR1TJIbVuLSXjM6Rog9PTrLLyYv8jxEfwUveySI4
jJPJMi5zjpbwKrzDzCNIfXNYOLFrO4TaHGTwX9doTUDRsEvJ2mSTIXivTKA9BfyK
xdHHUq+D5jP9g3XcekS9FE13eKN1fZc3YjSgdu2Hm5hWR/hg4G9l24ZGC4/7z7Lx
xFALFm2ZLal28sOulz3nFpkXCVdEs2vxqk7155mjtChGu84u8eKWT2Bmud8eFs8N
WolY4VgOQiBk/3reKPd1WeKQj2D1Bw/CPBFXGbk5UUVF1tUJtjIHjxdekNPQ6XvH
xCY+CYBYNztMa8sR+hHPBQS+t/M38tF+H95M0MajiOHj6CjvSAEqtkyoT8MbL3Ro
yFe5va2ZUqgG6vckLBx0QLL7FSkx8+3/TPGeXTiD/cN1eZVfYXGPaRHRlXFodB8b
s5hFwqarIM+ke9S5NM+2Mrx2hZ/NhPIvHoO6SORxVP0xp3vcQkoCvXF+5ZBdQjJH
BFWKCLFMyfTXe7Y0e8O+QbxJNTY5D7JkJgxrmLrfHHgy8/XMOhOKA3YiQplwkbq2
rgJREdMw3lNHA6QAvG5sPHVY4S8oJTYkiABoq4DkOpL5ErXWrn99Kds0ASOxqdu7
E6ENDbdRyXqymMkp+RX+GctYe8HB9LYvPXijTRQdu5rsjfkittpc2NPElYODB5Nz
n0bX9LcQFLcwoqAjBugTQaamnr0UkvoLrWrevTJ4NMj79AQYWi0atDPF96C5mODs
2eTyvH08dkb9Zia6feqXMC+ABhZFi1az1ooeL4CNlvkQV/8vM3UGaVRl7bQKAxIl
WfcqySEEao+ufDkQCB1Io7MN6KQi6dNsQ0YZ9Lgd+GRfLb1P7QuT5Rzzmm774kGa
xUY3ts89Rb9kDdMDFW2PbHhSbxkEksQ//TSxdkxIFEAPgLbjv/hnPfXtPA1yls/o
DWYZS9k/vkchEBZDU0dXdFG6etHXl2BHPCwjEq222ms7mwsOnTRkXMCLRGsqLMZc
8bfGycfqUnOB5Afxr00qNkqzIm7LzEHrvqMIvl0yl5/bYyHCNgJWzzptNTnAOapm
n09PvHERgCUbniaphj9PI4YsoiWsy8okBHbSJs+HdNztVcffIFHRVAidxgVAfXfZ
1phq5Tgjr5Rl7gILiWHrIxjkoUFkjZxAnxBA/BEJuyf+kOhMPQlAuMNSyf2CmlH9
Z32X64bzfHGm6xfZ5IytdgDoPzCnareVTA+CG3rw1aIyusoogSHFB+qKkLSPtNhJ
QWSNgj8tEBQJJ8k9M58OyDFnU4xhS9UMqCPTumtmaN/jKlrWWNmNT81tHinFR1ej
w8J+2JrN+MQOx9SZPQd/lkP5hJtuUfvZ1siVaRVgxXaXMI3R5pNGUqSiZU8FrXQ2
jZMW4upCYC+uFLn7T1Cw721NhSIJNa9RU4DzXMKwDdsA7d39/KhTl7pL1fz+xfFo
oJ6d6NvFPCb3r3wJOZbwkFztPo4TfVDNZ8zWZYhfKNJ9U9/OkvnDqcr735ImIvG/
3UJhClhFlhaYPD1jrD7C4XA6x3q9ASGsRQiinCOxV3arASy4v9/enKiql2nGOmMl
gNsFEWdGIYElq4Qnxg8AXh9Nx9d9qg7jAXp9hrCLCJMdt5QEcxCGjn2vEHyLP9zI
75G9YgHhqvFZX4y62inphqAGH/+dJKvMOdFrL9xHDPbFBcMxVkcIq/lXAImZqrgh
3nEEQgvHdAX4rwV01HSBmvQu2timWQQwJLwpHXlnxaClhPMbD/Tf5mdIsXrEy55U
h9spi6wJOv7fJugtt7nROWPCwU435Kc+dHEMJrEuF400l2s0rbDZRLR/vWYbWrjZ
NgRZEkm9bgyYMiTup2g6K0/hfKooHzRD8qxchHpVYN7Mg1JJLsaotDNsioksa7VB
5oZrvBCiwZhu0EFGvSX5xy+aAQxyZb0E/Fbjxegrg1KPtM9UBG7oSQhfRa3s5quw
dwmYp2px9iK16B74kB71kdQG/b3MBgue63KNqQEgvIRpkXO44XAxqufRNbeI/nn5
sSZvtBqQiSmTePiuwZXKqvE8IU2ECNPdPVFyw5uEaRChuyjcOnN5QHWM4e6DdmYP
gBdBQLYPWzsiBDT/f5bcDQzagIGUBbLpEo5fjBWn00mIRk9eiBRGienM2w3RTqvG
yQA2zi7V5H62fM4bgicpNQGtr1tFfC0KfMvCPw8yfVjINVq3XcJIgIFCiEiwbVOr
goTq7MQjCMxnO1SfyrTetDQI7Ir3GfvMqB7DdZKsdNpM/zevUOZD4AdXkVAuJe4x
t8w4jCuUcmqMbgLzxygKS8QYdVh0Fcoe3YG4ZB0wvN+YWRpu5RUlfCTg8aajJx9m
EuyR2/z4nrMS3iMAF2H7M8xPN836Gj1DO9ZTXfN8EBCRRzw7JgmId7RPKFq8QSaD
4CemiEPn5tEHjsBYaK0mQ1SXLogiBAFNkBB6TqBak6MEAG/7PVWWi9U/7U4Krdyh
dnBms6mvL/9NBiyEXe5MiO7gDIoPN9Uk6rkDm62HJX5dwi7V8MoukfJRMaaJ49Pc
t3NOGHLxXu/MfojTGmLQ7ku797O0OeFwxmU6QXOGQZ0BzyE2cFNYfbW8byzs5Ihk
+1Q0u8+DcaiYPJJdZDe6wahPBhNQoKigcc9a3qGY+tOTUfbx/yqb87I9jmwVHqRR
ghzlEUm/KyI5YU1QHlYXsFKU7IthZOrVtIIUXNHuQTNuGKFYadFjPcE/NPYhYEkx
z7J3TZDakGGKenrfkw3C6lGcrKpUxvMCA+BsBabVCWcvvuxAnulp2S1hb0Iaz2QT
qbtLaVbvvsDrZ7Lc2ftv8InR0ztY6pcz5GZ1MXt7L5iPeEdvZ2IkgmFWgvBZyxX5
PSYbMOXG7WHlkpPUkkfgkt0eoKrVQt2qfc75/KlYJHshTkQv7ctdI/fjKmmPnUrG
oCdlK/xWStLqED26ljwUAe+mnRlb59mY6S9mN/L85u1+SLD0cuXo68S98FINNbKz
D/lpoHSKr+bEhq2/E8uTKh+ieHXlcdGwQisnaRvUTEhHKL9T+bi7nyJa/3V3n/ks
MT7zPW0xzzA7yYJHN5ve5HLz14BLaHYSMbbRQwSI0KTu0zkyik6JdViqTQwnuWMy
+x7hnI6JHCTqmbmDaYCqaGuvm69x5q0gSIHj8hyhoeaVONLPJFIaZQoFhYboCMkM
P4DToCXLji8CBkrqzq9sSxQvxzj4kamAo1KNUkhI1vfIpiU+z9rpB+JPi8woEgS+
ykZrCuIqcb8H3/IzBHazODNKvISVaZPWOtTSCi1o9J8Ieyc118shJwRyqDqqCB5y
C3q4T4JrfbTnUj4FVDxwS4hPi490zviQV8t2qr0tlmdj2h41Br5tuMgI31BCIAib
irJuqAqIjTTI8PLrDx228X92O94FGMy1XihFMekHAM1/SAvXJ6i7csHeBiNNYbDm
QsEuSiTxwr5/RGQtL183VjJxZSor1Iaxh7Bh5i9eujEtDnSGZjlckOyEwD6eeaDR
9/tQCopoiwazTVVfb8JDFWtFokqtc39eRsTzHgQe1k+cTVbRNVRC84axJpPr9UCL
exC1D1dWpQ2k4D7RH91ORJFU31kwG19q9sW/xQuWD5u75W+sotfT1JQ/hHc3EsT3
oSOyfOLCQbimfDga/BdxKIENImErqGBXNNxB1VzYKRmOy3TmRbfUBzXBqTYmBCmd
5OZiHt/YNAlW9/v9xkehQ9i2v5zQJ/nrAcAv7UZSQOIXDnATBHjTiW9L0np/lb0C
gwNpS2pknNdPUPr8N0ACIp5DM9zx9cQetVAv/fPe20Mvs7HRtbM7vsMyRaZBSjps
BkjW+zzHfkn/dQE8+SMwZP65ttPcXkQX5LzAFRUQKRtef+fyy4dgfWowkIz0iHqs
LH7HLMrzfJLk/miFoGO7iVVmRCk7ZxBr9r2wAVHwGNMA5//6XWd/GxBBJVLh+ZDz
T19xF/rRuvmKkULGoWkIburCWDjbWU1TfCI/RC2Wifa+5PkomGsgG7CqnPZb+IET
+AgeihE0UJyZf1nLxKTAlrgIO4LDxi62TXY+5rKi1J2rvLENTTzc1WX8x6AzWn8v
qkAzML1n2GQMkXWdRvXVTaMnlvVKljvwNuDCL2+c9rzuW29zJdvJOgWW8z/KbvQJ
F/A94RzgLJom5SaUZ3xQdtIoN3apISU9wDNxe6y1sFQspwtyykoCdmFzLDJHBjw9
hIXy6CGJe+s7By/XRGY25J4Z0cgIZwx06dzEifO/LrBN5ladhPQAw9eYvxPhtVv0
hM8EJcLbRtoZU3ElI+7lArmRS8mh7O4TosGtCd5DO7nI2QDk2xgrJMK/ioJu7EX3
yLd2HJVkWR7kNWWz+cHadj4HJBlFaEFPM3aVYoXGaq7pIjiQ9eONZQifJRYc3W4g
6Lo2xTgK7or5KQEpNRzPNlvNEYcrAyZV0kg6PvPsUubgxGYZUxc7Y7cbf95rA5Cb
p4yurOkfF4zkBOX2motpdpm8zgJDYJi/3Lae8bsPQL6Z7JjAIreitGdt2sclxmEw
nKoijWPvoi+TTLtBiBVN2cetwTZbxvgBOB/V+I3u5g8PhKCY713ajR5V5c5XcV0K
ahpwPA3CH8OixwPAJ10jAelT/Co0YNbaypaBNO/C9alL3P1WBl4HyuKbzszTA0KM
h1/1jstwv7QTSejFYzKmXMm+BfZ3BlyqvGmBw3G6gM6E6sUzSOUUACa8XRWndFkN
9WLGCz8Oaq6k22bKw5LGVuAOxV0OsYpW1RJVW0cXFT6//jnNpaeAiUQl5VT/zBx8
uTf0OAmBTEVJgQzpKER2onW/K7YXMWkKJvlCjOJzXxnlRDFEpq/UJmdKd8f6PdXc
rjZ2EBhmnA3Vlh+w5QxNz2ADDlREozOoJ/pFBMcSR04GQq/+R8gOwXuR9jYcGs5F
35Jz55rRxLsESxDKJz3bWjS8Xl2UBnHffuFcDPMGn2Y1Y+AXj3XUsLqOVfWghAw+
dWBCJJg/5sL5dRXlW5+ABFPhJmIWrns63fGSejGUNC3ZT1Vkpazim9WBgeonPVSD
ElJ3SGtxSwkzyDW1hxC3bzPsP8yjsZj3DNsNWXXnRTzNVKV6fSzCsNmNxcxlqsS2
BX1nifJJzAMRUK6X0tapOLchYDTtyeUBBidhTm3nmP/ksHGvahEiEX9fhqLoegTa
hf9JgekGF23jQa1aO7pErZ6Aq2xotxB5qNwRjp4J/U0ceIT8b5NtQIfi1HFhzhJx
Lh048ieDWBYgvwy1nxDDSDbSIN+1J5WvfZ608TZltgvEIYnQC+tSK/+tL0SLffm+
JpMTO6revrbpMhMiX4T/QsFxqKqeWalOQ9yWaPBdqc+iEVIgsXvtC6h62qsqhl61
y84RWLdFZmP5sCEAS8jDxcK7ptoFml31bL+CZhbeoSDcubZQ0s59a3OcajF/whm0
lUR/xRUseSezeR7yY1Fu/Q==
//pragma protect end_data_block
//pragma protect digest_block
mQu8NdyHqAKw/sBRTWFlG9+N9w8=
//pragma protect end_digest_block
//pragma protect end_protected
//----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
UUQY2pVHjhE8k3eQaW19dn2C19CbNtOXgFvBPBaflxeZHtv6ABxZH7Z0EdRUwqGs
RqDVxeTPuj5enFRP/hWAUORsr2L2aW3GB7SCvBiJqiLyAJ/O7AfJzXc9/spl4NSq
8c8tkJ+5xMd8HWUdJx+SRCYbgXaHfoB08bXeh7/LJcyrQdKR93gyxA==
//pragma protect end_key_block
//pragma protect digest_block
kyGLwp8Hu2m+K6jj9Kum0g/n3l8=
//pragma protect end_digest_block
//pragma protect data_block
hKQOZU0zRQPMA8m4sIvI6ijTkOm8MLjT6RTz7HmL/GT4gCSeoYAlmnFuJw/cKEAs
HHS4KjgiOeDq2EkXi3PXW5tYEosljR/Txxr7EYE5xv1up+Veq3ikhdgPlfDbGwU7
W1NBcGV+MGXdj0Pd6N1yVE1ZiFhkbP2ZdvlPufiKY7fIUTNudm1toDl1smnJBKkk
YWwEQNDxI2oomhkR4iuE3QR/YioDZ64Hv2qQkoG3ZXH+LgFUEkJde+QMDD4C4+SE
w1xnmKafsmlcSYFmXwFj93g7C5Qwv7OCWg8wWr3Izqe7dU+VFbXIc+CaYCj+TBe5
kX9REEc/l2oI7etDWzlh8IHTuxTKxjEDhNEYGEDosD0slyZU7lNh7ofAQ0+floNS
GskGS9feS7rMfM67gorQH0mAnf78s8VjR7zQKI/XtcoLwaHUiwC7WS+nJMJ3J1o6
OAmh0IJyzvKNB128OS9MQCjqEtxrqcIrjw6hCLXVNuXwaEo4/9TMVvhVIu66QL7u
rG69KnNXhkBpB8KXBip6Sn8WLYATY9EDGnftV8ztd+JhoBvZMKRCS/8PzqlUAWCG
kWgKVFGc5hWRK77VzkxOjkDZSNbVK+9O2EaT8LYgWuu933WuCvt84ECHdsPZZKov
q/GhximjUkq6n6rOg28eF7mAMj2ayHHLw6POf94u2BkGoUyrKfZM+zBAmDcq17T0
IJUX2Y2VkGyPHDD4kpac//ni4GGtkZ9dBdk3d6z8uJbHSx9RTps1w/6yKqcSRnc5
bbtL4eIWA4bZXJmWCvkPRE+b3zFayDUYArUeUj+uMDWD6RpOLmq74JCHqU0dPVT5
vx1j4AW+hQrursMhuQWxbjXtWjNPVUOIfddx5Q9LNfYxgs9qNnfU3+AkEqalovyj
2BIXChHSw4r3tqOXNWy8Tp7fWOzDwFq5JX7XCcJ5of0mTsLZyMo72ZCOymFCx7le
987XHy1f6R3lbP7LrC/jLgMIkKUdYCKueQPJHoCZAevRh/GNq5q48wpS9mC6Z938
X4sOUnvJjwtCOCDYHVofLtpoE0+6iT+ddBShJBVVKC2oUnbTOBM59Zo3vc73Ux4R
B1HWnVUXLsmfVnEj4QXW3O1mstyR2LYGmXFF8Nyxvv/8jx+KGC0efqy1s9ovwkga
OtofOE+ArYjbzvdrsdWVXIiDESPFKDCr2PJO5UPm7O/Ex7feUiiB/8osW+xd5h8c
qTlRQn9AawCuCs6OCnp/4G+7K9LdwpOTc7TTxnp+RUYLFvqDJi7AuTOnEHTgatGZ
vX8SZvKmqWjwj6kyUx/2kSC66osf8Yqvc/co6obVHNWjrP1iTy7VZOwevpaF1Spv
s+RTAE29dVlBkHYYV8LFfeCNPTlOKPCfPuyQI2KyavP21BH1qtykDlepLb0v4vlr
/78XkrpCnSFVuCtSs6X4eH3BJ/9TUDKPLgDXuXNweoDLjFyQa25SeBVS0NazJtHO
dH86JXKEouVIhEuZQ6MZK6MYY9U5i/ZMUS1mpDI7Tyv0VoNU9BrfqdGZtIKclNJY

//pragma protect end_data_block
//pragma protect digest_block
/JHEeLh6IcVRoz7WfvDnKLIkpHM=
//pragma protect end_digest_block
//pragma protect end_protected


//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Y9ui3Iow3IQd7uEKwJ//y9Nx6vvmFFrjiqr8sPFJMIi2VO6Qphj+2ObfncCVqwsJ
BL57WRBXhir/zmZsrKJh2KcGq1u36i2NucLeD9TW3EuYEY1OHsW0br2WGwlVdWom
JNPtadIOp5YA0tbVzJEgNec+Zpi4ChGxhHYWTlT4mH0GZ9ZTH0l3BA==
//pragma protect end_key_block
//pragma protect digest_block
GzeOgJbzbK2l/aiSYa+6LQNxlrs=
//pragma protect end_digest_block
//pragma protect data_block
UuQ1IfqVMZBLO5Fb+NK2i0/sv+x0TAIRXkGS08EcbyeMQrS7AETgTraI/PhcVzUq
rPy5Csrkx2Y5tL/bpkwerk1EaqCBO61xmeMav5zLA8Dk5FQo2GCV3tf3ST/u7058
+EIkD0v+SiWMcbEk7UPOaTiIBA5MttMUKuluNowLn6jaJjmVjcZrm99DRE+7+dEI
oxivxW/+uoSwNf/UbYla8jkW3JUX5g3DiK0PBg3cJ2P0gNgLKiTPgrYYzrcX+EGC
Ep2g9Y3OMlNJggXz+uzgKCEuD8d7CBOqTC404hSRZlUHA4BvyYW3cY9SgZb97sA8
OdHLuaddvzRt1bXnwZ+vgkkW9/3yj5aL9eQkdQGP9uL8jUBpUJIFldPytGzzpAGJ
uoP20pkCYpPKSofZw7ZNgvHErB1r0mNyxMN85HrPKFaxxi46XmymfcECaVvT87Dq
expSUv2DNNFOAjCXN6XCBzquC+m4JtOyQjcIE+tSHw88KvWL2bG4TmI5QdP2dQs+
CiYcJ/BKSyLp1F+4QRqRIWXDy1y1Yy/RgxkHXA4jgXtdiDAnEPxOpP2zSsx2KTi4
h/JPhpAmTzrySW/Y4KxA59ldbZ0mVfct6TDNNrRbQY8wXR6J5qTK+u+e4b3gpMJG
s0v91EaxYuiO5LKJEBbJUeaGfErKGL7yEwOLmeuLEGKYCcfUVjes1LSgeQE+O/Nc
Bq4fYEkGibt+9g9C/LwSC0HjOhgaLPzYEKgrGPFX9Wz+AjqA7hFXCSZw/eUt9u0/
/5rk+Nqm7jxVij7oTUGN81wJiRoHutmFE0NtDlg7HRpE1W2NgwkufIq+3mYTjjuy
o+QoHAtTABh+yPq0ndL3StvSTa77ThFu2pnWt+ww2/XbeweIbgoVnkoTB8ZaQJnE
xCzZFMHezIuF9Fp4+xPZuX+6UD4WshtBCzjSWeWukRAUTQeyxKMOuDevxAt4fPF5
D8xQtcNwFpg2UnECOeqyDjHewN3Af5VLWRnCxnWKGjkP0a240CTQhdClSYOiRdqZ
bZZPrK7z6zaa0zGkZ4HYCjXwSjIuvagYc+UfmAa9lmzOgKULHy7gVBnNlQ+/ZBtA
b27gXAVmbHRUsf1BpkCnFdJCne/02h+98iqymS6ecvY/6V8g3HTMkWpyUFXxPJ6o
PLxArI58nkUtERKAdbC7dGXpcXTtz8k4lMpVbc74F47mCJ9C/xRfZx8KISg47zfB
dK/SPDBLigk94+eEUZd2cF+DZbqqZZTe1ctp2Rpa0dKGq0R7znrIoNbgDjgusRpp
wa4ERf6Mn9kGmzcvRQ692qW+KVxvqefU8xkvSSA50FH3HOmzilZlE552aIJCG1/p
jvqXPrjjOyd7blErPyCwnNzP4vPiY2za61T2wPpI1r1M7GWlFOh+R+74B2xiDuoO
Ky4yyYsQNe1IiccwgrwBttrZNNgstXlJUkuITcEEhVNwRIf1Q1vL/CtecMkqPeTX
k4RCv80L1266iLXlOeqFPBJxTXgMxi/MMmBOPDEpRIrC/MIGjQV/kw+Qz4MnkeV0
idAPqON0q8TXtWuEiD3KW9AtfSRT12jUT+U0imPlKLPzzjXkYeh8COxMndTWUomy
asR/zQG4SUurY68zBDpV3JfekEBGuvaOLjo9iB4xybi7nJB3QNDJ/O27LbYuNohR
JdaRi6/+fYC+VXlB54s1pKQsvurng7R9YIls3r5c8V85s3YLkJXWEPrlxx07Q69o
dKWNSvxeyN3ng+irCSQtetj7RCawHRLqaE6f2iPC8I0cA/6DHLK1MamJBKhquvXK
1HWRxhn5HallhCdiBNhy6HFxc2Em+THbiDa2nDezJPUJYD7uR9Mb4375sQLNnJ94
Bu3JswbD/Kvu9qlak0Hl7a9VKWljk+juHUtpr5PuY2GmWRh8qOv8AZ4rf89QoJ4A
t9/zAR0YY+eN1DGhnHtIZ2JNGbs56RYYrvjyd5g8p+tA/dEqOxrqYtl823RgFTvr
XbPn0J65LXAQXhFD4a7cb2QGrxfs6fgjUnZDg7CePP6wQ7QaqsRjp6rhR9Z+DfGe
5Gy1FgYX2DmN62l6wXUDYolEYwWlNclCu+DGCdOZuO4WeIYba9pr6yt7Ol7p4Ggs
s9LvedMm3vuk8q5CVVUdBWACfkz5A/J4WzcBMYCZFvkv6rPY9ZecY7kROI51xvZV
MAKCR8riZYSrqgKkYKpYirWqnKHlt1824Aq5z2OltFBJ143SnIa2G2i777idf95h
Ub40pmdn25HVGKtsbQNK+NmI8fbWz3dsrJ90JIP6Wk//33oP62fYr+Aqe0aKOic7
dBVxBZQvOUD+MRjEiQqKVYfQ6j0q3WloW6Hhh4lYpz3z9wROWSDmwXPRUXm1Mv+n
kqMz5V4i9Qcz0dTWvQL/v9f4Z2MbIiTzotYwBXMR9DoqN+mCQrni1Cr41HWI3jGY
hKhgQjRUqYv53/Qjxm+4SPYd+LD2kfHZnm/Lj2hBdGhuobFOI26o1/RvnFFpKBx8
xeeKE9HjkTJwG89LUUjLA/m6M9J5bhDwi9gmL/PBF3CZdexaT303nYxZfT0Vb+VJ
FMIomHyeZImHxBW+thLuYFBM6l7z4yL5ozVGs5YSj0L2uvSGXPK1gCUvSOIk/WAw
05o79ahTbc2L9gHKR0u2OzzR9tD+PszeVeWZ+B2JgDDhZk7yEj+TWcRuq+owADsQ
Kvh7/eVxttHx75lNIfFUdsMINWMtRLJuedKwQwHcv+/rCDf+GvXbVQvY7Ccnd5yr
zPshywRwQEDjhmyKn3nO2pdZagctrMmvsbhXilN++uTYmdxx9bs93c5CdH7NMhkz
bwl8JfQNtRfWj0e0M/piQnLzpJ9W6rFTnygjqFWOVZmAPITDLGB3ja+OxMqL3zir
zZlABqEtLViRY8g3l6oq3wfl4fw4Dbf60GNRAVLLb0qVIh0nF0Ioax5bdtxpW0/6
SyOGH8hFuEnqWxbCW0q11ygRPeTwRDQCJZuN0ae3EGTBQXiPH9ikiFPNBVRJyiqU
EdFbLnsbLIijQ8lqxawu4RXQpvQvE8MTQ2AsZ9wdpVVRXQMZ0q4YPhTNzb5reEb7
IWp1sGZfO1Mi24jZVG2vZQXA4D8liI3Y0LZIlmiLFQHpSoBB2sWQjRJUdK+u6i9x
A9kEBEU1A3T8PsvvzFsg5qlwAW5HwGrI83CqMwEVRwdShKXDBStEr3kRxImvVFyT
YMXeEjoA4KRORQMNcprVaBpi/2QlmdIcTKGUsN4x/FbLZW5cK3C3x+rM0jydGRbg
8KA+3/snpd7Wu2ygyC/eTGhZ5EfkbiCXxvGMIdeXk2VkbWxzK1gOb9oEKTIgTH2u
I/APp2dMSaWUUYnw1vIvFK8IHFJKP6fibL7qCUd00mZL8aiGnhm8aDaST1rwEyPQ
tpT6CZtGl/h0DZ/tp5IH2NdYgaZMOLo5mtpNNfDCZOvpmBcImwIgGyihVlay3IlB
opHftxulf7j2X/9mNUCq+5QRj+heht6QLAUNmdVAgEwwLEPF2QV8UoOClwppwkIR
ec81jlYEKDx7aRKVd229G63wZpIzyqE3Jw5RScBO/JmwYrL36lR3jwR+8D/5p4xW
frm/geUem0+lQpTkP9d+Wopyk4g9igSaFRKIFtZmcl3P0e8NUAmTN+gqtcbiFmHu
LGG/n8fBSzujTyjx+mvkw91iXEYme2epufe4G8QJbHSQ7amn2Y5CqUn2WESYsk4e
ZkJXYhuRv0SuIJMoury6sLVTNIyHpbytnqGmiPU0fhhpTGu19ugoS9BUULwyg+fm
Im4e0wJCcQ4q9YW3LyyjHjnGyjZHhIMGHfYuX9YQ4ORTxCrMnIRsyO6+w4hdjAzo
f6c+t8PrVB+hTQ13gc4Nb+zSCJ+RhengKvUV86RfWrnYuVm6G5FCm4UQZ5+QtHLe
pmG1/UC/ziJCnV9YRrpPd202PuIq5IIMyjvNKCbSp3MrxuPVmxWgFDbYIzesRpmy
/hs5scNwpXBc4qfmc7ObWDLTAV/772paG1EbTaUtIraj4OYUbqhvYp0PSB8aZcsx
KkNeC2lYf7JkM2SCKxVtIvqgu9C8cqbcmhA6eawjD3tTWMBoUv2zhiG/M+8QVnUX
73Qp/TItAtq3nLRwsKssDSdCBAd8SlnuiWXHwKLqLshO8/4PgIibzCRsbNUTBrRK
ymCTn7qQ8m16jRzAqBSWjSSYF0enMNyVmUepZqS0vpM5EKydPVrwy2507izu8iBC
0GqcOUfN0oUbWr+Z9HpleiGUv9owkk7s0dA8stBEvB5XdBY/po38ptP9gRnYO3Lc
STus5XeAZ1ZHrtji3wp2BMCcnfpl63+0U7d+3iErI/SS61cdrWLW/KQ0jA83LSjd
t1RC85NJxreVRaECX94rDG5bqWlWR09euuwnhPJZl3NFBdTuBkF1NDLfCJSt/yuf
bGj5W6uzvkFR05SZ2QCB6PsuRCQHFABSwmdhkh5wWPPyP7odU7SnD7Zrr4UZ4T9C
NXoGo9xqYyha9EiIYXYlauMsT9ckFkVMJBKmrCzK6lrtNuRhMgLRdpVdKxp9ryZr
f/JikVSwj+qAc6wmq8vDBF0DTkDJjM3WnS4PRBvbZ/ZlgCac0rcSKu+5Pa/zcYVJ
i0pe+hMJdkvIRxlVEYsjOm0qHc0VJthYqWTAIa9KdCa3L2rzVZ/Iljpu78ZmpMqB
R6rcbDbeCs3P7aceltIcVLsvVddhM5fwshas5LNXOrr3ViZ0oWEwuXlvoxF3AmeB
OkRhi4S/GkHrRcg8PZlXN+mInexeAu1mXIY08Wr+qlBHMnybh1lrit1x/d3OjR4C
F2OQ5j8CPp6QRgtTR+ULxJpMquzBh0uK5aRLTe+/3bCJyxNYCAcXGvbap2PRTHo9
haxZ3WNheTchVRUauYKqyizohKlaTZ8GM4OPOSVkdZ0VeLih2A5xjpASxp6+DOFG
hlBKw9BFtt43RQBzwykxyCuvQnoM97ZK2X0z8W6gTEjhbABjDCQKyCIBBf5fiDKJ
OiuB4xPuhdJ3R52vxJnLED90npfhI546cUiK5zUte9b7hDP/bSd3Yg/6Ua+VnoyH
uaVc7dz18gyM6IWTX5vYnvRAdaD6TjWV210TteTg2gLxXpUg7e/KntC4uI+3GKj3
6xPANm8YWqxCfFG4iiktnZ5529iEMEeRYMOBQ6d23ZGKlgooVDNJgsLB5z67ASVt
aB31lPszqSXsprfhuLZbiUW35RLSNVZh0Ra+t8TNVOh/PMtZV+17iH0W2IqvnNGU
GOd9uTHT98Vz73yea62/ksPT8jz+Tryvzb0XrXf+Vo0Cmsh5z6hGl81pFEGsHjf6
rq+IAVxiRib0eIkOCsz8ObHGtWLXvbCUrDdKF3bUmoRVxVcEei+V90K5eOLhP8KG
VpapOO5xWSGi/pzQOY1ex8s/GOWToABmoCYRPHOohQAsv5WlSl8qMKZiTDdzhAWA
m5QXuQ7ohcPD2UoaDxqNtU8wVBDIJYSp1pXeEeGgHSWxfM7hhxRcFancaB3mSXcp
BVpJJge/90nILJQ5Kq+FXTX6dHR9I+QgscRQKAcXDbo+6QJHnsiN6FbETlfyvNjW
G8rLtLA+EsIwqTek0DhjRaMsPW5ht3pf2IkAz1jXwNZ03RyfdpZpT++tLsfrlNq4
6ZrKT2taUfFbkyf4j39B5vz7XiOiVWxRrbnuwqRwchkfd/B5mH71SzIzTWVhG6qf
W0+5FY2nzpnzgakQix8Wq450Yp7Q3mIHlD8LAomoYgHVkJCUbX8jOTyTNFeXoS44
5cTdFklHDVEDJXwa5mSxBEO3r560ywwX7PnUE2QDMojvsPAZ304l5ikL7pWZo2dV
1Bkl7Eous8U2h75ZoB1pGj2oiOgkA/MRQ9Wcn6h7c8KNWHgB9eU1JiYP0HxKNM5Y
vXgvktVujDmvwCOh4Lq02718V1JSk+gVazNhLNwkrN2NgY9hwpJ3nADVxMp7Ba+p
+sDJGDWvT2BWvLNyshxmMLpnhqa8K0lD7deDlFD3LHZDkm8N/01JWYUvqW/X739g
eGWWmRBUAde8vi317Lk0qzBLMVaTzrNutQQqsHUg0GT1Ve6eSlQ++8hWS9yObAjM
2ghLD/oejKT9TENJSTPelh7tHlzsPhR9tLhFUqSnETmfywM/hgzq+EyJgJPxx9Mf
PzCrHyLWHBzymi71EmIkd7cAE755ds6EiIYjCG6WAmJLmD2ZcdGKEyEky9cx4xQe
4ESlmsNFYXVtXGGOhNLZMl0lx0tS/A1KJfvguU6DUXiKSppJnszjbGvUYuJJwpML
tWi4ffqspwiHfrFPnItBlDI8N4tlBuT9kpYKev9YJT2RTeWdLxZKEs2DmCrRjfJ3
WoXfI7kfsJ63t8RI2tZEAyZJvrd2UNobi5seHsDe7PurNCG1a4ot0JOZxUibL4I5
tlPdFC0HJ/ru1lwAdwS4kQu1gNIplxXaU8rOpvASYmKfYpCnr59SUrkEHRijlqOg
fWKXm7HtNMbt+tJof7lg0XMNY+e+WwDf7v4Pp0mVwHQA5l6K5m3ZpvOgGISBUB1T
NvHcJGPv4XWQs2Y0OSGbHDSupQiRa8XDuxYBCBUn1i91vB05O9gmAc4rFQq7Inwm
bjIeSECmPzbeJaLP6ku3VF3IpalrPVs/ye0hGnWxTZ4vV0pmxviSDBgE0Z7bfPa9
Buek7+aB3/cuXP3QxXggmwLajzMpmtf8f9cOFjbQldrWWFlg2pv3MDen9D2iybqr
AXqA6fV7NafmxEDXS3+Sg93t5t3h+8ja2Ejm1CH7M3OwJvllKO/oB83I2/KmfyaW
3kqg+dX6WI0/wIdllGgMuHVCf9jStp6dUk1dprs4EImlF9fWnS+7HZBQhZ2Ca1DJ
10Jxqpaz2JszWxQDuFeE2beZfWWH2rz/VerdiHrU8ZLJ+UpE7ZQRd9ls595oDulg
o8lyTiJwmbyQCExoqYIt77UT+ZvEoE3VZe7WJTXXPLvj7P0jVcTCZFAqKgmuyZGY
4hGfyFk/4HKpl5zcz3P6A7vOwFFcY6oqGY7PzrzWeT0cmk2t4bp6/vtoy2d2FR4Q
pVaL8hX8Z0xMA3m9UCJpV2ZR6h8Xi//QyXlvrhAgitoGjLGE7yV/wxwL512x4iZW
VfUitj+uvSGnqp51AAt7R1dYrdn81S58nW8W6iQnEEzRYYMTfLmz9JGzFfXrRnNS
/NzXmcNBvCTl0p5uH1Qo4a58RjPWejJK1V8aLN0nGJfRNGYGSOoXaaRCB6cx7j9L
Mj1OQyN72+qDTiHpk01dzXV7KhZf2GnFWiCbBgYhbXtX/09d0fxF8dJ3ArjeqSVd
MtC473FN8e07hvf9EPNqtp1mereDEZiM7EqeRfaYiwO3gRVkxGvVENhCsWEqzChJ
NNd5OMSFiJ5+js0xbq3r+2NcfUNkC73y+NMdQUDVt69eqnagOQYAee5jm3x0fC4B
phjhp0kYMv0JELqvaom3gMbRDHOz3epTBUkLIqxmdUGASiNO02cgqKcAmhZlTWLC
BQ16f8jMtQRX8si2XRzqPzqYdQBtB5WMHFeYhex+HKO3kLnLRHY+DCjvK2qqsj19
TOA22r3ZS0ahpasTxMU6y2ZpL+T8j6njWddRSupPxvzEfE9rPKChjZ7Xt7JFrEsF
u2ExLQ8mKvlKIW2U7moLKsjbnzN57db8nr5yNDgn4Y2AffpwId9EXDow5m7LJ15y
cvIk8rTIh2hTTCmSwp1OW2+s2MIiQU3e4bhHbS2BTE6jbcnSOGBTizMvdWr1BX10
jD6c04On0M0imzDeHX0gyU8xtUCbg1Vtrj4X2sCgwKerMhvLelNReUJaLxfkMMea
QccoQIcaF0YIP6A5l8Y59kG/O8Yp9cnPPNehVfoSbZNutH2lBdo8xdyElB7p4YKH
2ppGTCuu1FCXvrhBx8alcAYQfDT4w4NBhxUlV7bo/dGFKfdsuLjn/5kqVpnv7jFX
vYfNghp7rhnlqBEc//kC6Lp9mxSgPS4ODfhMtxQSIeHRcgSgOupMpITFpCvpXgpH
vzKjqc4IG8J8ClLMS2ndKDKvqCmPNGt6cuulttY7kjyHE7wpmTzfSC+alQYc9v0D
YWaA/eJpCKmCsA0d381FFn/6sk7GT5z3j+B5imJpeh8oIhHvCb/SKQZe6egljSqi
R6YTp67z3jeTYp/H91g1kL+BGL0IxOVPrn0pY8B5C8GZwQUUjpNrqNZai/gjZU05
lS3WXwnEKulVaQOOVqQ2HpqHx2Z7lBmK/LTaQIg+mf2MLdqGt6ajtnlA/mkbjKh4
UhshHvpH3yzEf+f7Y/iMtVy+SI3nN8cU9Ubxx1CnckODzQKu1sLnN1LxBp0KQPvo
SKvsLB0TPogRThxvTjepdrKAJAiYnqpP1SHRl/mx6AjnX9N4YaggdUBOuVM/fpjx
fH+RZeSJknn34rc9T0IzbsdnAuA2fldYNhrcq+ERggIxn/wyDNZXHWpqR25aqy7z
J7GRPxDJRKKK92Uq1NZgPFClsjkYUX2+lXksbi2kOCnCS7rs6wlmEstFaJHKg04O
BxwlZWDOl/2P0G2VoXR+JFPSywXk3wBoevB+5o/SuwJNmMtdQzqUx0cYfxSqCLFp
35E4KxiGn8fCm+b5xaGeTZ6GYqkuOnI7Ydk3lmeqZXbtkwkaaE1MzZjE6E0qBFpi
G8W1URWilbvxAsMWSbxcv3pCh8xjEKYSactS2OBx7gH9kwtLDAa5dRQGO/LKa8II
VcTM6XxG6fQfaI0M4Jks9yFDQJzma+x/D4V4wVbysDMHDmC+3VcIfSYP4be3a6TV
BMyIS4nOSrWRUdNlv3dsU3jw3GIQh6eKaBCwk2J2mjhRhBwv1NiWL7z9otp6euE1
nDeS8a1uIvXRtKv8sNS1M7JIugBnkO8i93+p5OuV74ciynUiJYJJF965qgPcaiBR
/RkoMHLZznRM+7Jo6510mab/Bt58PmDpWRZhB10EG6sn/yJvgNsxSTpEbWkFzCml
IzgIGlhhZfI7Mt2Z/ZoS99CeDv83pILsGnc4Q/DZ0s9MIT0j9rz2dLQog2DsVpj1
blE3PDwHBhyEbp8XNE8ESdNqRdXHGcfHK194/mvim6E9oL6ehGljS8bea81mQLuZ
m10O6SEdKLfTzDRYnwRB4gS6+Z+UDIIyv3CyXdZvXvXdACRhoi9KOfY2uc27RM09
rVlDZIa1TFbyVPivqHX7akWA3CSWR68mn2bn36TTdInuQIcI6LccNNQA+rXxEnLV
TWZ2LlRwzqCgHuPOUPfcmICPuV2UybnrAfy266XKwnhRHjYNZp5Iqsb7+qve1u4d
rt20ixUVDTGCHxo6Rcv63mNS6PADcQd/u/4kKDVAQA4/UtRVFk+54Wp5B+ZfCLja
tV2Cmi9aAzJMUTtu6GQH8PJ2XbLBppDRCMmKWSt5PjkC9USD96UhNlXfKKgNOvZl
t0aXqeeoXZp7eCqMzy4X+aH+BYFVlSkEmXOf2ujo2WACKKHG4Xf/PwaQoCKzMVgb
hVjLU6dRoVtGgp4uMfmKw0t8HsyJG7RxNw9j1J0Iv5hUDvdUGvd3UuFk8T2UBkfF
os1Ta2/xCj7pz2tV43cQ555P2pTa0CasgrJ581uS7BlgCMo7tc3c6Ni11sARwfke
fw0kW2RG1iU+BGIajq7+IQXv5gHnhPy/ug67mGndSpikhMT3h4moXymckET0Rmkg
upcqxX7h2nkxLRMlNq0M+IC68iHtTFOS28MOY8NpqzgYlprxPnQLl+y79Bt7CvK+
mWEYgsPnXJwkD/q+dX+UEMFToNfrD+g5bV20eHuHECiOG+vXF3HuAPUsD3hI8d71
ePP9kSqE96jrGDKzjxlFJCzqNE7xcpHursWFN0g0c45h4kmCiX/uVVdVcNUfWghQ
ixMSDzR44T7f3nI/wxmcHgm9QZ7bC21jgol1B73+M6LuluZz4BavQiH+mVfT2kLi
szHHTeQZWgY2uAuZtLhvFYcaQ8/gVbEnuZY6HoUboQVVYphKcS4pd0SOivJ2y+f0
QDoKz4FhLAP2Wwssy64Z/UpWnFdc9RxAPDw6dmSzig8y1ae4ha5CS7sc2NccAQj3
gJ1SQN039GlRGKQwbBXfcRfIyO6pkUttoBH/6yr0xSn+o88eJgABXqyaBh6BQLoW
H5oVqb6O7GuCjfhJNaju57unEZuD2zxFtbTT71QsNiiETUzwTilG+cp+RLrdp0FL
nzRKUX6vxSGuWvHEhS+AGdi9LrMN1Z+D2qfYz4ShqHKci2+X8f9pvXYOIP9/VEZc
w81Gz3Z4bhxpX/gcCcd9t7ya2n+UhGnUBH1YOeb7eodwbmTc3HKCuLNjskY/T48U
rJNNKvVeF3juaYpeRJfbe0yphjMvxE2tMFKJIii3mrIg0N1stosWPqqKwZGMpcbd
snVHJTssmcI4+Vs9tNMOJtqWjaA1wgw20PXyMzQLCMDx6Yq0IFCh/xbM/PiF2DLE
OT8Clmy/7iph0KWF56C8QfSVWL7GNLA9sF0VDAhvO/XaD93dXQUdRaZzKAzkun1s
WH9KgCtH+BN5oSThScAdy6P39pARlqwjyUMzgDOu/+FG23CWzv+zGoFnnAoO9QQ0
zZxNSZ8xSLkCSQdDdmgzos5DMh/41y1CHDwb27kvccaNlQJYQqMnAAjH0pGbx1Q9
MLJVeyOXCgz27GgyEgJARK2FVXeaK7MvSU483TfdaLzleNChsxobgBaPTrvtWyxE
t11MNGXBhykbtXcZ/9pfcG8CfEAKKSJKAH8hDa0qZZAvIU2MgwHW2F49fETkFkj0
ZkKdpGVPiA7CdOTtJSyyoHusvcY2ZD6d5kG1cmJxS/Hn8b/ykhuWE7A7Z/oeWU1r
MDKdMHHC2NqznUuQVPr1JQRdpG7e1POSVaWDbzHvzJxwqbjkVPbPzYdZ7VvJ9JQL
vhD1c5jKRyhvWy8I+fKzIOrOnzdWNmmMuIxky3Nks5yzH/VLURwj4uhc+J36qaVx
edSqRwfFl88TlUdiY9Vl4qqESspBTZT6pqS9QgJkEnwFESKNr4rU6hbpTjnYPpsN
X3qKnhGrxE1ekMNK7gXTXVBYeyJbAhS/m0z34LzCYmdO9/Ecvy4NQ2VCLrECa6IO
ZAg36I+6HBWLraROFy0m1nEnN7yZfBvOEcNQ0SRMDV6ZP0XNZ/DJKiB0Y26O1BCT
W81ndE/jMDPkN2aOAxqfmNo3P5rV2yOq0PH1ttfOy7Ora1Etl4NjfBsK5W8zwg/X
JpLW2yVJwHJPgg6uamk8Gyi9AuuOnp99Pu30yuyMlRVRbzs68WgwSm0GnEvOccAN
7a4NxZ411+Wtxlc0pTpHZyimzqEIqpvpUnoCtOzPS/t2KmVOHG70vUWvx4rC1wT8
7dk5cQbJ/oBlHlhUl9+aqfUz/p/ETTqGfSEcB1IvY1eqqY21Ot5FFLAr2/KrJ8uE
7GYS2Aln9hSK79qRZep/SQ5qWiJwq4CtSiRkiwJlzxn9txo/D3v/ytLPBPpGZt2W
7Z/VqbU1OPtyqoM1y+ZiQlI5BtEVlDr6HAa6CWJEHzMEPiww2mRCVML4NNwap0ho
YKIb1RW1rI1uGOM88XhyNzDqqP/fxWDponooZxV8RuasNukyy3iWSK3I9lgwc6eS
BBSft9rQnV0QmzCbdIAU8AJsq1Lp5IWxvFC+Y+znePqqbizWenWmjkRvHSO13OzD
Cdxpte4mkEDKPSzyvvGwi7hF/Amx158KpmjIOvLmuujFmzx4KCCEo6MW3rf+PjS4
3/7d918BckjFDIvvQbMr8D3jzAqCln3A9E0NMoqJLfa+cJkqU7ItLpMW9eOj4WNy
Y+ZF0D1KPQ4PQkD6eV2KRZvJj0fz+YYyFbbv3F9TNzqVi6son4KezTVwEgIZJ7P5
90B5s9aZfg4InR1mzquojPkp5gkHQUa/rpf/VTQoiFR7tb121cbZB7RELoZC7fdm
g4FZ8ryhwzRHAJdY/iCvivyTk9pR3ChfqN1PXpbwGI4Z71/+NKoNKS3VIhQGOpH2
zOAC65+NE7h0cbYmotp6D6VxxrBQHg33xAWE41CP1Wv7XdRsOrOjTLC8ludU8h4j
ELmerXD747kjUsuUB8kBb4vSms9wOO7Qg81losHG+iMrZuIB27mEfsvM4tXKvlWT
HAgZuTWn8JIRjNDnfhvG6z0IetIfCsXW1IOjob2utqXrc+R0TuT7UUg2BexSKFGd
RklthqvXCfXcemHOHHiDyF4misyPRoyhNbU2lg8F6OC9dqbsAKAc3Z5XChoovF2b
U6RTi0jH4Heg4+tRhN9xdm/ur+GOS51l2pyYpBtp2kgwItMu59CQY11fOUNlWumO
az4kH84YOolCSOUhNoZ7exWNhA3hFj3XS1GXPwjxq1YZi1rCeOsaCcDNMZHLoZEJ
Iri4OYSPb483Qq6hyC1KywxFqwCtHmpDHX1gt1D41urC032EM9/Von/VRuKZ4xBP
4b8yiFqavxznCmynpt4ZunZl+OxVJfUFFX1dPM1lGKPADizGONje0umODfgsavFu
DJgI4tIiscKuxZO0MXjdNq25ilwKUih0dJGRYbkeNC4nBtAa9oB1lgosS1nfYMnd
XwBqxQwqxaliEhD7Xcs9/uGebt+Ulm9k2x/IsEJmjhJmNijYr1lrvu7rhkjrwOhK
JOTi9QCczR4l23bOHpbNBfjhERM2L43GEoALd6hU/wQPthQrfY3zFkgJve17ssPn
2m7LZQvZ3wVRJRRfFC/Eu2mXq0UprWkUtvqJQxzT8cEL3LXzbXlQe2wT+CbOLRqe
xmWr/G7dDGNYPjivjGGGbfXk1SJujwelHNaEisL/Yzv4JW+sFTRvgguAxSsyyenc
scTqzoGnfEBJ+nflLGGuAxd3QJrnOX/QDS3Y4Ra4z2SFz5tQeALHjkYIJ0TMT4rN
CV6EWLXxpP4hIPdt9Uwj2EGnfILvEKcYuZl5wHVRojLUN7dOGAay/TfC0BEt8kPt
APUbtZPVZamTOls47Tfv8p3g+JxwVLmrNV7T9LEJ3bcPR5Pfqdx9/fCuJEfsed0Y
CpC7G2YhD/tNJ9fD4q36/dedImsSS6tpF+54z/RyFKXQyaMaPet3mc5HPVy0UY2n
rvIhqZbyF0Q5rgPAm6fjKVW1NAhSOpkewWpOyXuBNZ4SF8D4VnfHqIcmW7fT+pfp
B9fG4HFLkxI7NnDtKfZgJ3WPk/utu2mhlsiYwm/zVrwjOdgPCLpoPLbJmot8TbVC
K/GHRbE1skGRtlzd+4ZEXDIUFbbiSQkaCUKyy5qGuJ4paomVv7MsRBGX8XMcGjr+
8h1HicxBeoFge/X2ZrR1CkvYqtD4g4V/tQu3ukxBKhWTEuluUkWFwRGx6lrHknxy
HDssA6GseLWtGnWhXy7J4synI15j/pyTMrwY82tlEFyj5lr2+RRANsZ2OMTEM1PM
DYzLGMIYZGSsBHc8Z39VcpdZqhaJaCInDzP0ak6p2OHQ6yLAvFLfzXjfF36fCla2
t9e2Ni7xQNCTOl855N4cALvFTfyUYFkwYBbDDg9I7Xh623U9bJKCqTXvGhvnhDI6
bMxOAIlSmoa36BXBURnHyjfzqnoLqdLmtEu6wfr7bL0XwOsSQ8iG3hmAoU9iNKfM
OkJMKF7EFnC26g2vTUbYz3ZFMM1JPcDotexYtpQoX94xom1qqHTbUk8WoKMKHgaP
vNoYGJPNOkMH4EGEygtmxc+6anCHcnT1MYsqaEy55Nrkdg5kXRMf39BOL3u+HIXz
7Z+mhx3/Pxd3GO+DBog3erdMXiwmGOnl6pCT+KkbNgdZgLUqOscUjdJtJK5oYbUv
iyg0R6T4xtw7ZpfAfy1IWxYP5CFevpsdSpQAfapgfFy6CvFfRI8mDkiugzhCkdW8
c3//rC1PI3cnO1AYW3ZRYSlgSLLLCB8b+qUcfq9moCG1LuLTBGYeSQxhXINW7TPo
nrkT2MxsgUoROEP1VPJfla4pYP+xpoXT2fNsD94bO993vMJVn+/h1eFqOYrwZ1yI
TE2n29KK49R+DoeDxhqPZt+iaApbgCiiJz0S1wBa8pmT2cpzuCssP8iM/sZz4Bd8
M2+vXvJOVd+fXyPb2+/876JQ7LHxncs5WujdAbgRNJnoy6y2S4qIWCpJON5wzKHy
LxtNdTEOZvqXdobWzgzKSVATlFT6/xjcjZj2WjsLCxnRCHiDkoDX7mdnJnfOoEXG
6AbSg2WfaLmk5U2tNCs6BQcmmFmZPzoXQ20cJOoDKsrlAHR1+VnkmugNnYj7A+B0
7avC86LMDRCo9EGQ/sXN5AczQrdQ4l6WLISy6XO0KR8Y8AMX6Qxkh8vBgqwhSBiN
IfHzqflv51Zjg8e+aW2FYadQPh/c2UmDbgqQrDOojPnl8W+nkKChS/WkF7ck7z9M
dnADE7s2ZO23nRlddwl1tQ/YgiyPWlhyQFxYR7dATUvJ3mULrTK09czGhXd6FCK2
gc6hYUVf0zvsVy95Zxl7rVsdeizf72cQowNlkOqQvS6gi71gmMQ1DibvjYMill/I
xuFxdJYjvnYShyo8csagbTdTVLkCJuehOpq4UE2es7Aj3G6d9e0cIb/YFFOV2rOl
CU+y6hgJfXSKuczB9BYWVsOvkgHVjlkERaxRlHaRpIUFvu/bck5XkkiU0YTQiHOJ
GqN4P9b87NjN4HWSCGs5Vh47GVa8rj3NYwRdO8pWqecjpAp0I2GqF2GX/IpqRtUs
VHOPd9MXmtVhFIUCV3vFYipCGg4rbQtJ0pzc93Qhgd7gworbUQJKHdSVahHg5zOw
0GOiuG1+xthBBuFCvbZxrSGuz0kPpns4k0sCAMm7UxIPh8YEo0Nbu6kJ0n4z0E4x
ws0UK6B0BTD4DFSYg3SNRcIBdYaSW0YUk6kakW4ZAcRD/x+dvkD3SXeQlLbezpHp
z7TcqQR0oX+tbwC0g5VoCRD6sy1qlwK7QPWVBVnqc5mHfd6N/ONCdErvB704ipwf
ew+Qj62VIWXEoXQBLWtSGw2lF+dyKzmQ+/YKpZpUHSh+4+CF3plty9Tk7PcCz/RQ
BTqCeekw/aXeLt3TLlgL7E4idAvtNp4QtVfrT5fYmrPXGw5bz2m7h00NZtIWXBfU
gppbRiUITx13lvGonHg9eAVSGOGyEOcfzi2/vZeL5Y1JP+9LofzB52DVQWEhYdR3
8u35lC/DoShZQEv1hoAYsrB+aCg7csKO7XgA1iUkHbUe8z4vyuQVjp39VL/ZWKrj
JsGqdBT1LVtP+QVQ4SNLf3WAive5oHWQ71H5HTGmJvARzugxQOaoodwaiJZn/7GH
cc6fvnAWf0QHMCyOawYH6rqmKcOJpm26aSsOuWMngyF8A7XXpFnCH5DyQZP0tzd6
Pvi43mOuxtLRk0iAp40vjsKMSe6UqIvfz/aqDNuRTJ7KOwgsRVr0gNiFcxCWaaDZ
YGAlrHxsO7oP5FmdwHKqNmELWbHJuN9+g/Ppx4Ed81r1KDOdDLGzOIf711KW2dcG
vx8OzD5g/HfWLY/1Zk7JebKrQ0kj6ZhHYjewrqBs1ZrMzHLNeuNsrudC5wRUpPXu
8V/2c3vETCwzzE5prcImK+KlhuYJDQk/pdcc6dJtUaEMkEkWVI9F2Q8w0uGQp8IB
asgoKu+6gruVzlTyMM2eE2YYx0qV8qn132VnLQajGNNgP6NE4Df3yB2DymHjDekx
T/i/ndMuqK0dzXXKY8gQl68Zw2i22dAMOuI2cObbo1YL7idLcdEo4kT+gkqVRjKD
trmoNldXiSgh7Hi92oFCYiyXlrWHTN51/GUlFEmQ3rjAsGV2E9E+odaMJ4/j677Q
OhzN16DThcyv2bUraLmtrX+hTrY/+eD9q9I7Om9WumRfCEv6rjJQfZzAWlgxFCXr
lh7xkuWLPltAPPEvTMdBB90d5ErPEsHIiOO9T94J9Z0wTQc2vg9cXa5uLATp9B2E
Kg9T/dXQAo+QAPGiZTZEg00uefAo5UhXWuUXwW94i3mVEz8Vy964rJpuJA8/3Y56
Fiov+4qjzA/eTJzJJobFiP9wgPrt2pZ7gFIFG7OWVxX+KAgnMY05fI9mK3r7lvnN
P9NaiVpbuGIccjnYeKQcfmTOE5RmLKf8XNFOn731dXkMTAL0ROZ+u05XWypdz+or
nf2Lg56zKCve/xpHyf9o5U5pyrRNnVysYWL/dC7cpyUDkmK3uaRKIUOVANW2o52C
Y1N3uv0UnvZOXhxQrgChdr+BCFK0X0c0iYv2QdQRdSFEDBonW8G2iUdlRHefpv1n
V0l+rNKNI2jq9BY1rsIG9GrJJztK6FWmozknzfmsEgyMy0K5kCp4CTKWVacuqrEA
X3ZEvj3NKbd6afq8aTRzkAv2Dod8KeIQSiCezLR2dozvuV+MRf9JymHkQpe32m/K
pzkxSgljj5YG+Sre2YbgUAtckDD87updo/qnZOKFsjuv0RL2Y0vVrmxlJdSkfxy5
LN/nw15PPR9LiRkp/ZNeo0/5/LPUp6n6k7oCt7aODWHAosEigKX1DdjENtb3NV7D
Yv2pHy/3tgMBRHDZpk2cWGp4fuT1Hd3mym4ZWQx58xzTMBTaRPNfeZc8SUV6J91s
OP3k+8XaPPKdaPtOHwjxenk6x1eeeJUwFVimbZRMxaUDoYnwJP/y3dcoNAe4waHK
kVpwX+sX/nOMeOHu7iaCkD4MRgOGjj/KNR4Yc4J0dki4yaobS4/S6HPlTT5I5Rbp
UcXCd9fHTbUo6VX82WEls+8iaMSogH7Ui244iIO9pz2zZBkh7ClYG/XqxPoUb7zI
xN1izTZ+xwGsNS927RDwOGsK+BZc9qISj9G8/O/2nooUxbvjI9bcvV2bm5mFtDFe
M2W8lvaeVY44el/ccDKPiu/c4JG0zsM2uIpVYXfS+xFkzQT9KOo25KC38g8rCUAQ
FiSmZT+nWlk4g/TQn0o3i/BopMy/42gfp1aF+2y28AOCFkZ4nKqTBwVTnBEAGYgz
085p/YTOcSGJFZIYTxVSyIAqekDN0zoIkf1TJ5FhTd016W62einMAs6m3FHtPkgx
B+aTc5XaRblFl735bvTt1AoUNtNtCF5LYxIBUL+vHVaZLhYIpGBbry1S9OxUHGNL
iIWrfHXhG4kpAv/fKpfTliEUU1LiR5a23xjsr9hLFWJ+Adb5XB8qCOJTT9qGzj3X
KqT/5yTvkwzI0uLQbwV7RKYCt9dhiAZmdl5rdoCTbXPG1xenKN8igHbHC12MQO2y
VuoIw71YnRUtMo0unPyhnVDyq8oyhv7p3+OaVDHDY8g71aH22MqtT8+Bkusb/+aZ
WrAKmx9Wch/BsxJpHvN0evcIIXD186i4TsULs00FpVNQBAYzF9y2nXe9QJkfU+7q
dS7pbUhiBlSddkhJ32GWJA4BZoT0HusmDLYeufzu9g4lrzSpjnTPuBnw0QbhkuhB
4viQfSZIO68rRCYQfO4C7BYLgeK8ggwPkGmlwYkvWxyeE3rH20DRkX8wkswbzJd2
KjriOvBjlWi3uMcdsV940p4+8JBG27lJysgacblFyO9f+xnkrGJci73S5sb7zr65
Jk39QNRSp+1wTpVuL/wJ6Yx7jstbfbJbZGL9BqUgBa9HnbqjPM2TiN4Jz26afTUG
MwMdzSlajhjlgF6SwV53leV2+KJXEoN/5TDtR8bqVukCVFTXbi7tvBJSJhInwKqa
o5PuVs+MI+lB/YHSkERG5J/fAmIXRsBN92385burD8tDBrvfCOBB+L0T8crDmXFY
gSM+DUkQq/rwt0imS0sz7K8/2nysg4+GptKMTe/j0hMPbPwGW92S1f5/QZfxcgmC
DkyPxFzfeMwFX4ACUSnkr8Mh7rpx4U9ZzvhMl9j/twzLtpTbQ7fVqOV3JNDbuj89
bO85eF0QeLfAFY895bWKBxCvP/HG/qzdgUucF6DL6IzmdeKES1fujcy+gw5BpD2j
5PmHm+xlDFn90PlCWzyCIM6xXdFg2iBIkWcnRCLhyHudt/lOE8GbR4lc//yEkXZQ
hayGiRaKCyeqBaUn6gyoFQ37gFQfo1zAkquNu2hzL3DDdny/CFZronWxAUYqHBbc
OU6QGDIi0j7tQv6u/j50nImG18cDPlmgJjbOZRAQACU2jW8kzq4UHMgQKL78+4OC
Ti17RQK+FlN5cM6Jqio9u+GJi4UV3IKZHdhetMk9kHRKnXU3daWqjO3gAQkwWF0T
5cCLTvyZ513amR1CZpnDNR5XZhshgkXMHjsCFFzoatpFkxgnwxowMzLpNdgcbBNL
URA8C8rrLWQOgT6aD8sU89LgEIG/5lVYxB7KYlLPYe7X+NloJ5yYgVxRwJyYwevy
J6s/r7Hhrzu2TmWVJqj/jbyCwSwWkCMln1nZQFqOom7X+YMFsSwPF3puSSqRbGyz
2ZZvNjulO9UhsRzTaPY+fduYkqINTF8dEehEwKbuHbW0ElvF0EDlw35GCf48YqW/
8+CK0AOUw8CgHfXAoYQvFAuDHMTPqhtG6hB8s+tOcd0vjOLZ8S7wyRa3nHUVczSt
XfCWGQqaydUcQxS5Gv7mu4e9V8Fvkhqm/3FuQp+2EhnMcy9O7/BEdChZYGzyYfl1
bX0ea7YoFR/X+YUJ40qpqmzgYxijHrMxCVaPh3xQa6qL1W9atFO83Q1MKyrNk0yp
PXeFN1zJx5lT14W9MeZvVa7OkGC5yVevJmKEgS1Y/mqnoOW7RuR2H6az/g5xXN6a
6va91kLQplZ8graCBFzCfUI6RsarKrCL0Nl+Q/grjO8cGx7QkPaXuW5Evh/JtwnV
1325z4RjUqE12B/8uO0HhdQSash9Q5o5Z6BVxNoN8D9Q2i4lH8H08CA5O+4t38KN
aWj+u+mVx0Jvc2NKHTU0Bc8vjNd3pJzT/AGN0wIk7twqyCpAY8GqnUawWClGtfEG
jZxxgr5Aht5Ts21mSAgMjDGupy4edqTDuqN17YubAUghpamWtn0U++07ebIpzwgs
LZM2XHmgDK+1U7NeNcKlAVXJT1dK3UH1MOroqbOEIsMhGe5bteYVfoq7jU+3oGZA
XKh1Jkbd86DE1usHU/u4tJttorkmEXhfnxu52AjWEK7hIcbL1KK1LT5KmRT2a7lX
P5zaQsYdanv/UysIEuI5SK7HYs1WJr6/0Y6JFIAOj23clo2X9UyIS7pwOy0vdDdE
pRa5UtqGZHsaubTqtlXBDlvoHHB/Az11E58TLPtOMdY2j9dKq4TpEHEVqMlbA3x/
01abpGQPExyFca4j5m/esexVvqg/T5mNXog8WMCy0DlwEKZI8F3vW6DNosudyHmO
IrwRpfOi0SKGsgT8U9fRYVf3agDOS+9MsHGSAk4UEZy2DIUHHYdlIKhCyrWVkMbd
Ysunj7fucP3XddygAHbgPeHsCZr80yiDEhhOZcojkGCRlqB3cHeI9jPixxbmxC23
L0MvOiLl1eo8isVE7+HJofU43tzy59Fb5X82Lily4vZ1vgE7I7q+DNhqtTiRkkOl
6HYjihODjtzJT2wEl/sOv63/AgBACJ4Y0B90ESkPN7FskgqEgLjc8dXnPEckPXM4
yPDJSd5Smc6PGjJcUJDjIp2uyJet+f6c0rIkaNLokr+TfslcrVh34Qa2DcZNs08x
+5EPXNnRSxVM2UOCreZnyYi/zO8hWsUMuy5x+IkWw9Z1M2pM9nxodFcN7iMtzGGs
QYmCCK2Kfg0QIEQarMuHI65dPGXbgbBsIyzT0FrlSV/XACcfEG3JSIVaI2I7nfos
4W46KdaVCdc+JUK48sXjWdYOHUkY+91mGAmgJX48BkqTaXLW65Fh/jgj6T7aWwYF
IPE8Evhe34/FwYrF3ZG8lH0ggdmh7eLffP2d9qFjvGWZeNCSFhIS5bT6hjA6ugKu
bH8DczBknjXG5D3RO8Q5Rrk94SZvkSLLXIRmQ+yH1kHc4SGBlpDDXAv6OInHyknI
tWKbN1zfHw9J6JLs/t+IIy3h5jCxAgiWaS5vuqLFcn2vkIv/sUL1loM85nDR62LR
EkAMUXTBWaFTBMnkZ41w0kTEGFIW7nFtRogsaA0QPURoptRzYGDIxmHXdlrDP8g0
YPpezYXpllsvNyCtkiYZmS38hbEYfN8qz5srk5uwOM8xASxHNMNDrVZG8YR8nE7f
EV0hX/ikdgFkgI7LYyuP2F4uhxhDZH5ckmoGz3luscfv9SaJW22niZWYt9ScBAxB
Dc33yMlc3jIUjPpkoqDBoloPnjX4bIBrlJE642O5oHTJWRSIgJXKtw8e2BrtnvOt
akMAHOOol+PLsbJAFWuRN6cAf9FJXJj3jpSyshcYkrlWvFUVAhw2IDWH6mr70clk
CDXmZJyFacmCXTLUz9lPWwcR3Gfd7g+b/gt3waBxv7dJMTBuE1AIEW9S/nhiKg9R
KIPo7dIS2mWBdKDkDmYcRyXJoe0oCoRXWnt4T0dyjHGnmFpXS6Rnpp3K7jwAsPvW
EWZfCDwv+1pjJKTIFms9WSnOhuIX4JgLZ28GK/xvngJL9uFWNNoMFwpmRmcQaLQR
gcke9fkP2o9ueM18vNyE0qK9i4ReLLjpepAfRS3wFotmYRzIe8R72O9hLGeo8DJL
J5BW79QcGZgJEmfTTTyj2KMwZJKI9xbj1p4nalvCx9QHvRaB+gAflDvfMnmvr5TI
V6kyGMIsQ8QMYHZepyTpI2rWVezHt0+gV0UMrn0tbPzlv+hJWfuibsuR7v0ox78a
Fwpgc3Z8NkcVony7tBjGKTqooNr8tdZKM7vPWWC5RBtJRTehm9uFPAdFLGz2VBnV
c7KQdiRpJYPG2DSpDQufFVthNMrzTpL8Dx7qjrgts40FREvgenzRyCCtCtbUpL4t
94cRsCd5f0IV11GMCAyfY9r5GFRFrT/SP6wxy71cRaEsMNGkbt6+xiL/HRX/3dlU
EfMmlAjhUs3p0NIsnDzW4aZzm3SWDoi9+yh+ibM72GUG5fxfFnaFKtseZbkrZMqa
yVcipqP3vAogf3HyZlWvi7RhE/kPmZlZBYc/gCUxrNEe91Zax4829X0jnJKuQg3R
Cxm2unS7OxF0zCq+DkeroSkIHZfflDASQEOvylfnbouBMRqRhcec8GOloJfvwM/J
BdAOrkP+j9jrg9eoLO5vwgX7n3PgHQ2cCDLmcJB+IB82HKBhCFBOhtyUp6ElJiZo
tvkX96qOf6twZXJHVMbNpaJpIz0s0FQ3eUNZBaa5dxpoNw/tLl7o1OD7vu8ymwPA
S4nN8LLPKwAjjsatFIaKmax+1lv9vFXBIulHVUcbU4RUD86echayzUVJLPk27Sye
yGIvScVXPuhl2UBSwJ6AodheQLswuxdKt6verBEth6TEMXKEh8CS/L7aYTACVocs
L8Fi3tHfRvy4XvKZt2mz0mOC5aPWe15I9brszdLsXjD9iMaRDtTFdsDybi7UWh44
cZLpzE9RwOOhzGEm5B5pBgUEpAPV0/WQEdFKBFCX2c+6VUR+c1KHLxGuPPQBrYui
quA24g+0NG+5oGPuhYdJzmxKACkHdhZ99hAFBPy5JR0M/sGwpr5HFUlM8RC+6Vsy
6JG4EUj0lkgg4xgk5RV+UpgJ2yWYgTaNIsSRmqoCPPyaqiqnd6w/1+SWRWISCkZw
FF3jfccQ3LdmzOmwxYYI07GbA9aoo6Q4/9MrhdICuEbSY+/yt5oPRuAUk1/y8S6c
COJ6wFZOmbVhvx+LRUu/Zh6/pz8fqLCZJPhkY5BVMhEQupFGb4iJL5u/dR45xvt9
7A51FfY1BkoiONJaFcKXdMOfDkIso9b4URQSWPluUMgU4pCH9WEIMfy8N8h5MEBF
jT8VEvrawfzfgRkbgfPNsv95zBct26CImg+1BKmWgnYapUaeT02IMZ90XpL+vTeS
RLOLUTnwmjETdWmcbf1v48QztTdtDw3TQNT4AQ4jusOwSyPjvRRfJcjRSRbHuNKk
/lUYTIXGMNV2FbcxwH87i0YNN+G+DCr5o06rw0BTX2hDGsCaxwN+ACdogHyg7DMl
VL3Plp/HmB9rHrzf9oa4qyEiZukxPIOuwIZzZyb0l3xdxRzWLkXVR34IhlO6Lujz
5YsDhVO22HydlWNq+ydUV7DtjSVh0NSjHlQF1CRjBTNqXS+Fl5d7nd0Xlzr+Ja2l
7omQpDTvbR23f9sIG6MEZnxRzgbpjuxssO/6+BLmfxO3ta5RMeCnJXJADxlmyB6M
dCb93YRdCu8rv+fRBDT+JEzBfNzSr67ZuU16bBj2sFHXTx4Drh3neRuLWdmDIq2W
mD4WHSXFj/MS5EarTd61alR1u40Cco9X7nRtvlxI5WkOThFmhdjCwi1pzl3waJMc
VU3mH5bnmDq67OrzIsEig00I17AImqHYqrcMARgDGhTjSeHRsNz0YLuDDpvre3JJ
CP4A5QkL/lXjiDQ8PFZBbNgHGS0lztfQjB3c96aXe9rZu+PwOt6xYKHjkp3lBgMH
o5p+/S+T2vtLgNW07ZSM8nDWd02y8/l3MNQCBjwksqFa3Tcm+cjuvWLo18sJZyAR
fqbBzjTDArHLKGkVHHsHRrXj3UOsrPoCmyuS66AnIm93ruS8VpWrYdvVQmd8wNbS
UxBQwCGMxXjr/wH/BgFGcBsORg3+tcN2npOFwoLz1dcPrwKGpxkyf19HKw5mSVj2
kFbF5+Azn6aJbgjIpdX+WIzjM7NAatu9YM6r6X+mj4/A7htnz+bWH8DD53Gbev7e
BA/rcg0dOccZQ6TiOIAF2S6+/ngEe9Da4tPeXnsY2RcKf3qhDHSRBayjUr3Nm7p7
ylD5V7t5e3IoNrvVAHtmsxsEfijOwX5nMT6ssWBLIhAxFvtCr0sAT5Bw+zcG86Zn
WF0ZG5jB7xu1dAOOq+0VHWws0gQrcWrbg4LUve92ABgww9D9geXosMajeJWL2/aO
5upbNIkmZF0hoPRJHZ5Hgy+rPUqjIa60CYORJE7aThMOsSytOVz5kflGRlKsCnfQ
S9EYyxwwyS9FkHRR0AHxFKnVlF7JsM8Rz0bXr82gdF0sGLAMOPhUDR0oPQtaeHq4
0MaljLECf01cvojWuF5WNNwXIMpg25AKYjYE5/f1p8BW2ZJUoish7GbeLEwr+tAE
W8BZZIidWIKn9/QV9HkyYxYPZLuGsINByF4Q9q8htwyLfLSLsLl4PL2OPC25cmXQ
PM9S4piXpIcy7dPiBhTh3fJZd4SlQj3L11j9VZYGdbJKe9X0PVrNJEGQJ4LW/2pz
kjwp3c0SmV+YTJErHyevk+Sj0LalFAJ+Wz0nYlx41QAsnzenCpbCSXaVhFj7QISd
KBNHsTOM8RAdBtT0y7XKETeq5ajhENwK7QSCMcthbGXWY+gTboUqLHSJDA4T3l14
xlZh6hoDJLcIkUJtQ1K+Plilrn4K/ZRwyTzA05ztD1j/Hb5naa4TCASeLq1wS9WQ
hPZNbL+MAxH4HGZhYk+VA4IP/GXd3Zx1tSXQtF5txSH/2IduSaIwBqRWJryOPEyS
HUXsdJWx/TyAE5ABxVrGtaX1g6GasaNcdhymRqgU02vBm9ZPH6ZGXJI6FsXDS8b/
uahzzLXZMMq1IaGTMxYQ6mhGUm5HRPtgN/yqh8uDRqwDEp+UKJLDKo1ERLSxRFtk
vQt+g8W1Rrj+zBJoNx4hD6kxRz9Ey75xyQjGXGNY0BN2RByiWABB1TdZK/21WKzx
/I5MzkZ2pEmPnFSwZYg7bfiu6shLg5lYvdno4oNBq7B9GfFuCvnO1hn7gt5YLMh5
Dg/Zm7B61egaA5fLJ7R6gxc6R5P/c2Wa0tu9xzlpF4Vsa0xz5WAHGt337/MIlifj
8q7JdFlxbv+04WCKBw261sk31SWyhq3A6maE+75F0BnyQ6MWIN8I4lh3lXlR9fS2
veEP2pfRHb18fljRQb6O+5clMDy7TCChByyT9G2Y9vuoMce0tSHZpj4d7I76cfdl
HIt/UoHii/BGimBm87lPra1MyZnc2IFr5dQpGSwYp3O2BzZ8wZ6WxKaBqMyetLpG
Ao0yo1vMsw5sGZfBXr4BDZi0b6piUTpW6t9L1Q+HjHHbbuDhYphQpnCZAk8K8Gec
tmg5Bqm9we3urnBIlwuXXQTvc0EVE2TdNPVuwXR1fpVRG3FMBHTtEQlp0Ya9Yfuf
PYYzRdnmYEAlIg+YsuWc/5qDe/qDfn7LRE1D6GvrhZdHNitJx/hU8mVQlQgnJOii
3noJx0DYOtT8jSCwJpMPm3uZdRvDY8miVI/EkVPHI/Erviep9EvSRI8POVtFubm7
IlkO9IEnMHPBog0kaBUXrrXxII1XEJIOXDAJl4gVYzvAGOk2XxXhvoAqFp3aUfuR
kgiMKkK1gl0xCu2DYAKIf8QAQD3VLoqt4Uwmo2SUhQdm0t7PKAaGgbNy86G8zg8t
gkrWB1LWReB322BpSxJZ28b7xCB0HOIhVTGbw9rFyFAZp8Z0b2wW+frjpUqTCyFV
ZOOWQ6aLrQvRDtlcsNpU+Awg7JsYK8IB4661KJp35AlNu3e2NyL4bAeyCCzrD+4Y
hU9uuhfmweTwy5EmDCekA9UtPVjjsINWAuNnFtMULVcZOpW/xgLvTvKu/Y+a/Tbo
BGwXKsO5/iqM0lgf7np+Rgr8mWt8MwZzXm9+19cJZ+qJYWFfZakzSnXeGF+FE8nm
eLRbnHKslx7DPriiDHd9/yXEvW2zKGbd1SQQ66WXHLB10bY1ARmK8a+A1gofcMsh
qypHEOQDePy7KXxHqpBf0p/ltbeXeKO5rFKqgYOFspUKiD7YDw3TPDwr/uj2+991
MPhU7euy4tUmTCJWvUwfXIhq6YC0M7OIdZd6ohL7T+mGkhauvnSDd5j4SDXARIJH
hK2CCMf4OKlxvaK1/JTcjsbuRNQxhy1ctCzWtrrkUBo9zpHeO/XhECX5IbJTG75l
NQHpyXor6aYU/HGscMp5D5Xa4ZZjHe0Bzc5NwdFdzzsR/hT2LukxumSa8VYX/p65
IMbGWBtYkoX8zGPGgi3TnwKFfCCXtEbW1i9xjCn/oDdjdScLSiESmh8zJ2Z1RuFB
pXWhMRDW6Pbm4qOwbRWIiWTar2ETTNF/NTauEdvPLGZSUbEWXwG8F3UNYzTgw01k
JhMDzVmiP5vWJL0Iz20c/9yDfH/lNfeKsStxsb3529XQNWHHrJ/UlX1bDXRJaot2
9h8jjYq8F+Z20bxWVcynY3MWRVu8uuUm7sd6NDT9NMluAqfutBlL7WIPdwfZL4/Z
djuww5QSNSvgT4VvtAse+fR5ZdH5hz2epsyEx9rQUM0hZZg1o9PUGzVg494HuUZ7
psd0vCW5UtWpNx91sqHxl60Lui8crt0OBE/IXfb86jG61Wd35wx2TeOSjV6tCELs
fqSbpWhUXOJ4kPixYA7y2Ne0cUQS4up6NKl/Aqxk6PImQdlCwaxWH/fiXxN6bRp5
/opKfYXsAA/qDHGuPeQpe0LdL+2YC0QbTaaS0zTIRBkxPVZtJPy4HskTvlT5k/iU
BpaohvXF0w88LqCaF6dbTQenOVInIcl/paMAjHm82QHYcLoaXlgc283RRdV2APMV
lplix08G6w8na9QxFmn862SrMmHE9uYQUDIyFzRM0zF44FWjeRshcBLjurh3hMu9
sTTx8XX1QlOJPx/uJys7etucD7Np59j8SPlMEQu2Vfhrfr083aXExcmFKQ+Pa+9v
lSfb6LLqlB6PkCGuFno8paUd1YV9MPEeMYud3IbEmgFudYBcJs9yrnyRseYWRUMO
hmJmXFrCp5Gv6Gfqbd1gJ9MNb7V6vGBOR7P4fPPPRde1XumdoDpQwSr2Uj+594nw
7tZ36VTkAvC/cZM2VIIpbeZRpxgxVvXjgKBskqTZjc1R48E8VjRZVltLZkw2vran
K7KtqeCF1w3ZikRQ6s//9qNHqs5w52e+8tOFNV42bvU0x0bbFTd0O9o1NU8NG4ge
lFJnRX8tcHh0VC2Eq1kIDINtSNlVyGcz3vHSwreAhslsGrhps/YkDOmr5uYrt3Nk
Ti4NJJ/ZDmniMxxBt2QnooY3oiu4IetsLs12IM8MxPdfs+ypx9Cx8d+6exztMK/B
HHFc1u+ZZxjFO9XI777Kcv8K++l0lK8Db/HnHhm9iXuk/byuCfauYDweWFBOELuG
2qTSm+VnrzHhN6QJDZZtQk2Dq5P/utjCp+ZgIaPMKD940SrZhpUYjXuLvTSyitgu
A1MoFA2byGrTtscVW7u19IqyxZUx9OC3fIE5PcKKM7esHAB9aoKgiwpDR5rMhMY3
3UltMK3371W2hRNk6YjSb5zXyTj7OxGKiGPnh5synizla5j3Pch83dCaTxF1Y/J8
RxjkvlfktxLsq0g354TCq4t5aWlGV0OxgAJ4jV+KjF5S2XQWF/W44mUSvXNCkGwL
yUfrvPZ13EODe2A8qNi4+d/K6m/jq9pu8k0vcm7+6nm1bUHt43nO4WxynWQ08ZPb
LV51OmY143iW5JziMxSpfhu6iUEA467whckaitP94RRHIRUUluCvWtocPN2syNHH
dgwW13im6HGJBLzYAPcBq0Sr3LmaRxCUqbT6L7e/JEUSmp5fvjxf7lD+lBCT1lOr
RaIoGBIve6/UG9+sQaIuVJzFhFACaQXHB7IIBgHoX0boI2TijCyjdOFBWJRCnNnH
8I9r3wG1aJ2Lumvs7GvmEJics5EzbT+CrmuhiEY39xT+XbmfNqEoeSSg9QMeTvyd
xCACTuukhn0uLRaocYtnf2l44yV4QO2af7JbnbUDqLWkcOrKnFBCm3TZBcNOv+OX
UqqTOnqvmWw3jAA+jqYGlRQvAtNVHi4BYEG3m0xGVWzf0czUrqcqSPHDYoHOCrNJ
25VZF7Ktdj/uVDkSMbuFpc1XDzqDbY2pNZiLcWKserFU22FFbz3401sYTIk701Q/
KXymsHNG5lrOLe84vMImynjjQCcS69xRsbGPvkYU60ssfsGmCdbiqPcwUVVZCDQF
Wug9gxrkqMwddogbv+hN4ahUIDhCtejSgyiKiJ/srGCK01UkOO2PfOPKN7eeOWxB
5rbQMetkhA8RYpXa5w5YwuvG1DOGvO45SUYUMIIgMK2C8toc/gDzN2LM8JJY28rx
zPFSvWq0YpJXI9soLkmpeZJh4l87iSon/AcCU9/KhK8k/FymgUOZRJLNMfRjjg1g
/pz1TSxhmaAqZGbxuS6BlDD1pI6nk3CJgvappjlRp6WbjmudoxzONWfPBjDOYJBs
Z3pgI9RLcArEw1EcxFeW46b0O/wSj+EkgBs8mykdMq7vjCUDHY5EW0T6ng+/PJNK
yDRRVaDu59wwaeBhZaaXfIPSjloPjvnvDjxv78BBEKg5egC7/RQrjyfKEEUlJunW
hkggOPnIx4ER6QZpEmxcbBUvYtiTir3emfY0Z0wbxjsH5VgRtwaoqjKzpBZZFx+3
htMg8GbUFVK1h5w+POfiDRbpox08kmgi2YjG/wTHIPErwC5BaUNt/BVXheDEEQ6w
DvTevDvPWtX4WpweXSIi6IgkQxRIq8N0w3tZuXUn4IFmv/wCPmA2m8vA8QDC6jod
NcF7c8mrCRfnZaf6JLI/ci7ARvEqkaRkZD1ggtLFpzMR7VrTJ93sZqXCrz+sB+b8
IoxjM6qtvmv/RFK0zRx50cCNnE63dz0I29GxWLQK2JuFyO68ZR74/I7saQgYWhLV
L6vA64v2irAzHh0bi6HNGYg+SGWBIi+FJ+PxgVtJcOdGpoSlUoYFl3zLa+3DfIA6
dpU/03f4zgWVMbRmq/93ig5RB/TEzI/lChuPqTbgy4DIVlIXsctruA2JbPq9ga0w
5ww1u9UuNP3GRXQ9rFKMHRf1Jr1VtafDJYWxajwHSeXHQ+QCZuuIshrr7ZwtG+HT
+rfbMHK3fmBorW8hLIKxELUzgubzXNVdv4dlZjl09jLuaIX+/UbzFymiHppxKDvh
WheZ82z2mDySemPbydsxDgIlNrpkmZFY0ENUQs90iB9RUoZbw6nNne7TPWxzpnk1
aZaZ1UU3QvyZ0ZcWsNZScS/cxB8w27dQx7vOejKnsu4H1zSaPx8Fim+3Yn/l/fU5
w9ptpTuSWPiRZtsHlcTBDszNYJ2Ek5q81NvGwQ68+06SwyDm4TDUH0/x/ud2hmS+
64lw87XFhmVDOlak3i3NQBfv5Bv5O1+7k6x2dBHqdF2GeT0H6f0u4GnGlcDsZVzJ
cHnOaVoMohkaYvdjNgr4CJaLtvGwwmeh5JX0BItb1o53x3Rh3AEoUk4p7DIe7gD7
m48Q7/PXC1fE4mwiOwlUd9GYAPS49/Z7LZ9p/SVsBTzvzjRInaErXmK19KaRSy5W
EAnHy/JHAGZ9i8JBLMgB6emvYExg4hrjw+IXe4s+prlqfE2TY0Hczo6z9+HnkhS/
FBoaZs2tBKg6CvwBOlRCw+4axGCBR5QxdG5LwHRegObzNd6EN/6dX0S6waXVxSWq
jyUwIZ1PwyVAXGFxBZd6wfhF9LwZFXiP4zGABOd6dR2ePLZ612Cp04qkZuJ3AwnK
NEFwesXz+VZUY6N2YJR5DaS5/GSRaoD8hRWiwwL2bez1T48e6pa70wLJFofMhNU6
L/H6rY5/xAmSBw7vO19qtiu6Kzd91PnOabtP84YQZydpNvnG40Zc+okC61V8/krv
hZ8+mGAzE5x3LAGjk71cXwzRQV6uHP+KWWC8EjalGtR1Cj8eajOZ5p3+sbX0ki3U
2pvurGIzNkl0OBke/5oKkQT694LUVnPYkysGi7mNvMLRdbOiQNvFKuJF+YX6VJwb
GZwTZWfgX44Ilz7c21bWVx7AoWCnYMrNOHym6iMIb/Mr7/TvkC2oHh+K2ugI004o
NPqHZl052DGjU3gMepO0X0bV/86M5a5BGxjvI50ejpXeDRjbInkdrjkVO9Uq1cMx
EKkJ8sTVwE6jzQopl3xrzOVGTeFd18suli7XSrHWRVORpX20D4Yv4sv17mcSu6rI
eMpo3TgWeH2M2H1zJ83TnipRXFG8lz5E/gqI2desXa4/JkDv78IDLCcCyUHRPPSt
8TSZHP2rAd8WbqPONvWDAlPYegcHMkp/U5ad/ClkNpYfOjxEykHzCYGA6eu5UthP
YHiwUUlySSficVBn5uVetraV6ZwzF0QLbQOL/MvYCo0AhFJw1+dlwacBuKMl5HGU
48qKL9DkuKYeAnkKoVzutDCPnsFUQTJ1mtB3pqMSdOMty5MT4qjkc261TXQqO32F
3DJk2beD23YUaPopPvZzPM7vJkNTw65FpIkQ8zC2O/iBKgySUgKZYubuGJ1/tCqj
B6JV3wGcsjxBoc2A9QYaalmVe5Y9bYVZ5pMQXX9TGaQ3L0UUJukpg3PqT9CapfPD
WEqsLrGK6ZYTC4scBK9b/xdKW87YoGFNqE6q86BzwNI9CaSGcwDIOE3mJyuaJB53
TBWAiq9/cp/pDfXOcGP9tLdOkCzmEjR5utMx85SniZ3nHdlFsBaarW3gW+K9P7fg
6gLT5dJz1AYCflQm1BDXbXh4Nls361U+YFHHgX2QXnDcbALEdMxITnP76umPsp1M
tCvqZWd2lsTF61qz9HE+NEfGc5H06YHwrM5c2UvIwfeIyWKs5QWFisi2I/iHoC+n
RkUhKJ9SmOlO8LQrN4suAqUlEzD5rBoGUoNC6r/KHq5oy4ehfBMElxI0ZhEEi17T
bbcnlivBxVA1sGdzERQYo2uZXGokzLC8rs4eu5cPRPGI8RuUI0+ZMlkLzmaXVWf/
KbfD0iryK+ALAbLqG2WuYNPG/Vhp0g4t8udMGZBXjNFzeRTAUTGZAvvV9KS5021a
BN+lKCaNo2maaSpNHy+3V0uIQftrdn+2CvoDETfU9/VKVs2pyakhRhtlTfsfjijT
7xgGu65V7EKD4MtYzJ1KsiehUkW4PumYtPXeKWdseV9iBU7brOEVzqWbCPCauMQj
rR+hFcc0fjz+I66A98xqIf51k7FWCGZvEVJcb+RRNGvpNqSnDlfz3kfjqD7URZsr
pWF8pLez98T5D5SqK2pAqd9aT99OotCtMXcrKfVO1qIGTsst5L9Kx1LdFAadDQOG
3ZO7b4LrI9bvuZ9DmfI1VJxTOfz4Tbe98pLlD1jdoB2NauCbTg7MNgKI54mXpDOD
kV3vOKtmkOEZyCEZlE2Gur9Tdw0oUWdazz0OYT1lHplGwa9stCt/BIk0iMbOyN3c
3cPzF/KeNnhYaaZCYHgaIpgrMOmjv7GSca0R6hbtjZc4pipPEUstMdGlmp9k/XK8
NqkCZJY7+mMfq2G+jaGgHZ4IP4dypwG2TygMrRmT43HFcc8TdT9RYG/z3XG26c/p
jNNyujfGSlBvH1iFoneCL5tcYJCmkcXMQ/4XU/4yWO87XStWqd6e4KboHuIa12XT
sDgZBQ/qlnmo58T/2IyRsYWWi7DdJbaVYw68we8j8PFOyPyIQfHA0f6hniWC/xR7
fOupLM2CCBc34qTcdlkThkDVWNeTtbXmpwL4+yfZ2JKEu1ehLiwzHC5P2/oK9wHe
TiLm6XdJgYuk6W7zouB8v/CW0lycVae7+qek5YJI8xUfYofd/R1HDfokrLp7cknf
MPrLuQLc1iOLa2WOdoNtTbaFd3FiL5OQeATIPIe3QMX+2gIP91rV276YvS0yZ+KY
13MrCFC/ZpnKTX4ciLD5VN14HghUeUJGdWyqb/pC6FIg0RZ6mcEThUiy9ZagbO5Z
ySXeFrtKjRmQfhtqaI9GD3zHCuHpiMOku1MqdmA79hIKHzw4ufz8bI2Z9aWWhpYD
sw5YMnWTdCEcUT/ijffjgZob14gI/DYEEbgaDksyFdZMDJDeavOFxAKWHsy6XL+S
QbGZ7m8YNMSNmSIysdhOrOCtiJcMX1onRs+zzbw6QswmyBmzPCLDShVj7CleJ2Er
xSRbztiyzb9zsuS61xJayZ/W+D4nVtpuWUvYns3lIXinZ/1xSPfUYPa38Ccgts5O
k0EWrOlgHu7jrvPY1s//aztVADQy/cLUDi2rhi/o9CWxGTmn0j3zsg9u+Y3XTkgB
gOZSI+DI/mBqFjKFrI2ffaxgcHX1uuQyTJ1GW0DTu3HOEEDo9ELU1FlTNYCbJeLi
oIF1oUkcA3JhZs4Oh2PlVBRU7KWZ/BWGwVQxGll+lpgIVIoFRvRyjik5a4h5V4am
+rg9IN/615qN1qtnDTaJ28P3NgiZpMd2ko3+d196pGlpsePtl/VO+AWSuBMb6UlT
La3EYLaynr+wPzoBnPqUYIvk/BIj/HWYdunTzWMeEPrN98ZJpEfHrAJSSRiufgrM
B8YV0mBtlf7cWPDwawbTzCttnDEBm/lBl32SlmYCoHdjw55TRNwoDXRm2vAw3xBl
Ehs6JeAPYELWlXRn3T3HHrl1NPM9T8BzbqiQgO9NlguSGfGa8NaWBDhiObK5dLwX
6Mz8s+8SBp4ZQMuc+BIFyE8YNV/FBzMF8A93//y4q11OOr1HIz2rR9p5al8TjaKK
jfoQZpgTHfEP7lPx5o5KUlYy5T6EFYx3/Qjx1L6F4wtIisF8cDDmAFjU9wymGx6M
35pj2XzvK0Ddr+DJSaTcGT/BmZ9Iki090R8C1zQyTrgUnBDX1JjU4NIfU3bD6IOj
g+3UBdVW2X4E9p0ahr8LNllm1fPT9XREE4xTXvMaAEUcAztVDrfIp6CkL9PEOHLD
EzeV7Rf044vRQOXccY6vorFd7Ee5g7eTJXhtyNqF3lm1qOcpKbrStF3nobnvXO8/
qZv0pl2NB/Y9hOLZ6+1BhqR1411/Q686Tp7bTCMnWs8sFzKa/pFp1BC0sSbeHPfB
Qj+ISJ8/d9xT6FcbD4j9cEOojxcJu1EsM+gwn1irxtbXBeKvWdrQDJlBP7fXjvJx
cN8YvCq0EOLV/3rLYaEfLaVotbN7Gelf3LpEQkwNWcYFC3sDrVgAcOV7563QbJLV
7buDoLFV/3nHRTLct0riJPKF/nt0hmloTGN2APiRzxq99706e1P1j6Ki94SDO20D
Mfi0fFKHR4+xrcQB5SPBfQ==
//pragma protect end_data_block
//pragma protect digest_block
MELS2vsfLHAfybCRW6Vzhk4KN5Q=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

