
`ifndef GUARD_SVT_AHB_BUS_CONFIGURATION_SV
`define GUARD_SVT_AHB_BUS_CONFIGURATION_SV

`include "svt_ahb_defines.svi"

`protected
89;O)\>27ZI93/=2-fATb#HQ<f13fNKX5PVS6ac7C<;b0e9+gKR[/)XY3>V2K)NR
[K;^&WNbKXX_LZSBWD#IIMS=]TYaRdHR3H9LB)KSTQR5@E):_aC0)ObB+))@B<8_
V(c@GU&c;JbI/K,\_I#K))S&baLaUS+__A<&,^6S)17N&FVDCUf2?]4,OPdB5]4e
1>\b,:VMU=@.g<_&TF-/\7IRb^O2-XZ9F4A-A66:(OO;Z<+N\P4d6P@=;;\OHT=5
NA=bf\M92WPW0[@.T8beL-,B3D,;]PJ9]DJ_Og)\==YIaeLg_X[<ea>[Z(1L-((1
Z;F,E(6C?K^CP)B)b#F?XbBD/:E>BG>1\)Q=V9Y3E]W4IYefX9IGK,e-2C]L6)5(
aHX;B+B5U&GHOYX^LFPaPBZSN-1d5)[<-C9=LC_Ee,D>^,@.WEB@@#GJ:H-=0,g_
2EAB1NcDUgaHFO0(=G7/;AdJQ(/OEB0ZFU3(CT+PU?JN4A0F:#O4=C5(Te<0YFL@
0U/8XXF[&4PYJ2HdJ<@NfcVK_2NC_&=PK,XBJ2)V.a##Y)8,,AZPIK[SV@T^f342
.RgT3=F:B_W3?W&PE1S3=0#J-GE,X_+JD0dL_/A2(OBZAb\\EDW#/+P>c.V5SB&#
)8Ke>>X0fJ=S3P42b@XX3H^\a-Q[cSXLZ-.>]MT(&9=Z_QK@>RG,Q5ZbHZ8HEGUO
C#->9O,6[K<;<X9dBM2[3A&PF1K@S/2)3P([]d](OK]U?XI?^?B:.+D6VMI3NHV#
6NI,G&(0e5T(-DVJ8D#WI(>-1I(K)f<KT;fMf/EYe]?/,\9A42&HSH(dUH=fAZ,7
CYc@SfIU4eA+D+<_60\B8S[AN0<NgJgASH6\CN-:SID#dYU7.O5PGTM6P:L1&^Y(
9\8B@fF,4#=63ZD[d1@1(;4#-KRE4\#IS19)cU5-)bDe:7,HMR@D4>4]0=c1Fbe:
EgO]:L7+;/Wg[(9QGbU)LBD6]??e_fVNfSB)&73E497\fO+>V<<2J4W8607:;d+-
Ff6HV?F>IN70S#B?EQM3Q?TY#4Pe.50-Z2O^PKKXEQcfK^>M0#NKQdCW?eTE>&[U
&8?bM\LbFD;f26R.E^[;-Hd.GJ<=E\WCa&T/_Y&MKC9@bO5M-(O@(QGH[J7S:76E
^K=F]8HHII\SG12D[-]QJN.VT,C2._fCIYa_Z5aCY6ZWP&BaE1_+H6],g3ITLRJ(
SPOg;R@W(ceBAD]a\-;)Ya(A-6MfYbJ01ZC:R0B13-8[LO[]Y+L\Dg>HDAN(4,gG
GQ[+SMSGXYLV[-VSYd.4AEDN9&[b;ZU+?8.5[eGUC8=V^)^gdb8FKCBWT7<aOD(&U$
`endprotected


typedef class svt_ahb_system_configuration;
typedef class svt_ahb_configuration;

`ifdef SVT_VMM_TECHNOLOGY
/** @cond PRIVATE */  
`endif
  
/**
 * The base configuration class contains configuration information which is
 * applicable to SVT AHB bus ENV.
 * Some of the important information provided by bus configuration class is:
 * - Number of bus masters
 * - Number of bus slaves
 * - Address width of the bus ENV
 * - Data width of the bus ENV
 * - The AHB virtual interface
 * .
 */
class svt_ahb_bus_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual AHB interface */
`ifndef __SVDOC__
  typedef virtual svt_ahb_if AHB_IF;
`endif // __SVDOC__
 
  /**
    @grouphdr ahb_bus_generic_config Generic configuration parameters
    This group contains generic configuration parameters
    */

  /**
    @grouphdr ahb_bus_signal_width AHB signal width configuration parameters
    This group contains attributes which are used to configure signal width of AHB signals
    */

  /**
    @grouphdr ahb_bus_signal_idle_value Signal idle value configuration parameters
    This group contains attributes which are used to configure idle values of signals
    */

  /**
    @grouphdr ahb_bus_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable coverage and protocol checks
    */

  /**
   @grouphdr ahb_bus_ebt_control EBT control related configuration parameters
   This group contains attributes which are used to enable and control EBT settings 
   */

   /**
   * Enumerated type to specify idle state of signals. 
   */
  typedef enum {
    INACTIVE_LOW_VAL  = `SVT_AHB_INACTIVE_LOW_VAL,  /**< Signal is driven to 0. For multi-bit signals each bit is driven to 0. */ 
    INACTIVE_HIGH_VAL = `SVT_AHB_INACTIVE_HIGH_VAL, /**< Signal is driven to 1. For multi-bit signals each bit is driven to 1. */
    INACTIVE_X_VAL    = `SVT_AHB_INACTIVE_X_VAL,    /**< Signal is driven to X. For multi-bit signals each bit is driven to X. */
    INACTIVE_Z_VAL    = `SVT_AHB_INACTIVE_Z_VAL,    /**< Signal is driven to Z. For multi-bit signals each bit is driven to Z. */
    INACTIVE_RAND_VAL = `SVT_AHB_INACTIVE_RAND_VAL  /**< Signal is driven to a random value. */
  } idle_val_enum;

  /** Enumerated types that identify the type of the AHB interface. */
  typedef enum {
    AHB        = `SVT_AHB_INTERFACE_AHB, /**< Interface is an AHB interface. */
    AHB_LITE   = `SVT_AHB_INTERFACE_AHB_LITE, /**< Interface is an AHB Lite interface. */
    AHB3_LITE  = `SVT_AHB_INTERFACE_AHB3_LITE /**< Interface is an AHB3 Lite interface. */
  } ahb_interface_type_enum;
 
  // ****************************************************************************
  // Public Data
  // ****************************************************************************
  
`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  AHB_IF ahb_bus_if;
`endif

  /** A reference to the system configuration */
   svt_ahb_system_configuration sys_cfg;
  
  /** 
    * @groupname ahb_bus_generic_config
    * A unique ID assigned to the bus ENV corresponding
    * to this bus configuration.
    */ 
  int bus_id;

  /** 
   * @groupname ahb_bus_generic_config
   * The AHB interface type that is being modelled. 
   * Configuration type: Static
   */
  rand ahb_interface_type_enum ahb_interface_type = AHB;

  /**
   * @groupname ahb_bus_signal_idle_value 
   * This configuration parameter controls the values driven on the address bus by the
   * AHB bus ENV when the address bus is inactive.   This helps in detecting any
   * issue in the RTL which is sampling the address bus at an incorrect clock edge. 
   */
   idle_val_enum bus_addr_idle_value = idle_val_enum'(`SVT_AHB_DEFAULT_ADDR_IDLE_VALUE);
  
  /**
   * @groupname ahb_bus_signal_idle_value
   * Used by the AHB bus ENV. This configuration parameter controls the
   * values driven on the:
   * - inactive byte lanes of write data bus by the AHB bus ENV, 
   *   and also when write data bus is inactive.  
   * - inactive byte lanes of read data bus by the AHB slave model, 
   *   and also when read data bus is inactive.
   * .
   * This helps in detecting any issue in the RTL which is sampling the data bus at an 
   * incorrect clock edge.   
   */
 idle_val_enum bus_data_idle_value = idle_val_enum'(`SVT_AHB_DEFAULT_DATA_IDLE_VALUE); 


  /**
   * @groupname ahb_bus_signal_idle_value
   * This configuration parameter controls the values driven on the following AHB
   * control signals
   * - Hburst
   * - Hwrite
   * - Hprot
   * - Hsize
   * - Hlock
   * - Hready
   * - Huser
   * .
   *
   * Following are the different Idle conditions
   * - Normal Idle cycles
   * - Idles during EBT
   * - Idles during reset
   * .
   */
  idle_val_enum bus_control_idle_value = idle_val_enum'(`SVT_AHB_DEFAULT_CONTROL_IDLE_VALUE);

   /**
    * @groupname ahb_extended_mem_type
    *
    * This configuration parameter is applicable when svt_ahb_system_configuration.ahb5=1.
    * This is used to support extended memory types in AHB5.When enabled, this extends 
    * existing hprot interface signal from 4bit to 7bit signal.When disabled, interface signal hprot
    * will be 4bit signal.Applicable for AHB Master/Slave and in both
    * Active/passive mode.
    * 
    */
    bit bus_extended_mem_enable = 0; 

   /**
    * @groupname ahb_signal_secure
    *
    * Slave for which separate secure & non-secure address space is enabled i.e. bit is set to '1', it will accept both secure
    * and non-secure transactions targeted for the same address. However, while updating memory it will use tagged address i.e. 
    * address attribute, in this case security bit, will be appended to the original address as the MSB bits.
    * 
    */
    bit bus_secure_enable = 0;

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname ahb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_bus_masters;

  /** 
    * @groupname ahb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_AHB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_bus_slaves;
  
  /** 
    * @groupname ahb_bus_signal_width
    * Address width of ports of the bus in bits.
    *
    * Configuration type: Static
    */
  rand int bus_addr_width = `SVT_AHB_MAX_ADDR_WIDTH;
  
  /** 
    * @groupname ahb_bus_signal_width
    * Data width of ports of the bus in bits.
    *
    * Configuration type: Static
    */
  rand int bus_data_width = `SVT_AHB_MAX_DATA_WIDTH;

  /** 
  * @groupname ahb_bus_signal_width
  * Defines the width of AHB control sideband signal control_huser for bus.
  * 
  *
  * Configuration type: Static
  */
  rand int bus_control_huser_width = `SVT_AHB_MAX_USER_WIDTH;

  /** 
    * @groupname ahb_bus_generic_config
    * Enables control_huser sideband signal in the bus. control_huser signal can be 
    * used when svt_ahb_bus_configuration::ahb_interface_type is set to AHB or AHB_LITE.
    * Configuration type: Static
    */
  rand bit bus_control_huser_enable = 0; 
  
  /** 
  * @groupname ahb_bus_signal_width
  * Defines the width of AHB data sideband signal data_huser for bus.
  * 
  *
  * Configuration type: Static
  */
  rand int bus_data_huser_width = `SVT_AHB_MAX_USER_WIDTH;

  /** 
    * @groupname ahb_bus_generic_config
    * Enables data_huser sideband signal in the bus. data_huser signal can be 
    * used when svt_ahb_bus_configuration::ahb_interface_type is set to AHB or AHB_LITE.
    * Configuration type: Static
    */
  rand bit bus_data_huser_enable = 0; 

  /**
    * @groupname ahb_bus_coverage_protocol_checks
    * Enables protocol checking. In a disabled state, no protocol
    * violation messages (error or warning) are issued.
    * <b>type:</b> Dynamic 
    */
  bit protocol_checks_enable = 1;

  /**
    * @groupname ahb_bus_ebt_control
    * Enables EBT feature.<br>
    * When set 1, other EBT related attributes svt_ahb_bus_configuration::num_ebt_cycles[] and
    * svt_ahb_bus_configuration::num_mask_grant_cycles_after_ebt[] are used to control the EBT from the bus VIP.<br>
    * When set 0, other EBT related attributes will not be applicable in BUS VIP.<br>
    * However, EBT can still occur when Grant is taken away for the penultimate beat, if BUSY cycles are driven<br>
    * between last two beats of fixed length burst.<br>
    * 
    * Configuration type: Dynamic
    */
  bit ebt_enable = 0;

  /**
    * @groupname ahb_bus_ebt_control
    * Specifies how many bus cycles a given 'master port ID' can own the bus 
    * consecutively before EBT:
    * - Default value is 0.
    * - Value of 0 indicates that the EBT settings are not considered.
    * .
    * Configuration type: Dynamic
    */
  rand int num_ebt_cycles[];

  /**
    * @groupname ahb_bus_ebt_control
    * Specifies post-EBT arbitration masking for a given 'master port ID'. 
    * - Default value is 1.
    * - This cannot be < 1.
    * .
    * Configuration type: Dynamic
    */
  rand int num_mask_grant_cycles_after_ebt[];
  
//vcs_vip_protect
`protected
3-&>X/UNd=S-G7Qg[Ef@?Sb/6F\YFa)IgR>6W\?\TG,B^K100#3J4(Od]S-bY+W[
P;S,gS;ME8(>W<FQb(V^(C,WS8FafIVACY2McO39\9GX:^RL3gT/-HRS?K^?fY^?
@=;9GK@QfI:S@ATO&#G6+U4?I[?M(7R=4+D.XQV]T8GV#1ZE.NSS_Y0ZW(\43H-1
/TB6U32Pb.M+5&2SB3=YLYP7K@<2>PQ(fCD>&4^/TJ=9&DVNGTYOc\(^=[7TX,;E
c^cdX.f5f:a;]TD5+-2JV3dc6W2UPR/NR/b@-3WbF8dcF_:KDf\IAF;P05MOZF6b
aC<]D1HI<E60bU]A4f3I1>^@]6P8MgFe&E0;&d7B>4MXb?^,M3EUE@cITRVRa13,
\[KdTgWL>#f/dGJNXXfN^Y^cg7;Gd=ZF<6,1-&GFMUCg;\RBG/A5:-I<Z5,LBV=U
D2NP@._OM]L</?.Z2W)LSf?E[?/K/9F@>4#LZY<eX0+\e?>A0+<YVUH99/?&6\KN
DNQ\Z@Q,R=A?+DY&5B-R\#HN4R\QYJNT[MH5IL&G10JJ1]IOJ?=Sceg.fD.E4#&E
<H3-W.^>XYCQA#^&&L.d^S3DdNBNa1--M&#@76B\8G(?^:FSB9TfJ+@,&[OTCJ_#
@O2A@g<R<b2[8QO5M15WP;QB=#X,:fC8U@YWDf/V-IdH8Q;-OI>7UIX1DI1fI0D&
O<CVWDa=AgcgQ(HFRC04TG>LU/dK@+\J<@1#O)2-[EOeOL^XCe^.CJ85XO#=,6T6
.U#EGdYB:3YK2MNPI3(NgPR^&/H@>BY(4WfU[1(<XG7=EI3N[(e1@2DK.9U@LDF&
R7W)URN[dG9,1<A9-O)0W,CANPE\R&/U+ZdHVV3Aa0&d[0P@9c87_+1O.YeJ/8R?
#>L6XMG?a->Z#2SQW(TJ,DQ;+N\^LgH#,BH9&4Kd#6C10EE&7F<Y)BLf?>c89?d9
[]/AD>A=KX;OO=SfXdSUHH=QNb2&>O)O9H+5N9J2)[L#UKFTc<-120?[H+3V<<U&
9+H,-/ERe18<g(>,ZQ&D3RLA#+5&fN^9f)-+Z55:d2db&PH7H+\fe5PbeX7D>e,e
:#IaH1DY4fb_Tf@Ca>Z^=b-IA9LKYJN\8Ge-d282eX?YPTUF_[G05XH:X-DK8IZJ
3&@FeYZ(PKB+D?fK6WcTb1J3AROI8@^ECSY#:/f8^L<.<BWP1,#W)Zb8#<<_dD-F
,V+=-#Pg=fH@1cT)Y7(dNQQ@I/F46T5/TDIEeQ0gT4?f?^g4K(J#8CPd/@JMGR<J
#K(O)#>U^X[))<8<0CB7[bJOB1PIA(J\7-f5?;Y:0;H,Udg/:)DZ0L\4g+A5O<BJ
ELS8XHN>IR#5>Lgg67PWA-3>\fR@+Id^5EB#+I?]^aD4.-:Y2;g6V4X>FCH;@+2K
EXL[1aE)0^0T3U^]<Kc96AS_?W]CB;=^SE<B]JPgYUD0=I-Z2)5CH^XeZT7?/5O<
?W/VefV_K6IB:Qg1_2SZc5SgcI77Q+9J-Bg(>BG1S84J8T<+/23&-Ed<#3&De2+H
#[,G9QbggUI2^cA-6+L0;.,B]I;,O;d6]B=6>F)?gGad.aIZ;C4J5P@T\PY-0T7P
<W\1/f<b/,P@/<fYQCW<d6JBV>4d3;;E-6MQ,8(;O(/GE>;8;;/QffY@-bB&d15/
,9[6&ZO62;UeHJJ)+,]_OM]AT^VOJ2ePM&C_-U^#3/dgT6=5N52NSYNL+C2;eIDe
cQ/AI]O[S\Y?a83,=@;3&c-4;7V^B6]/Q:A/18bdeKZGAD1_eM8VQH\:N=7@#<U\
5&)MG0_&WEQ=>FXIZWJ/5LLHWZa4[gf1.fB:gU;aN>YBXe0cZSRI]T+SIET1KY^J
X-:;.Vb3E6e\<;)+eU;3)?1\<D_4O2fQ=T/,e8E#:6bR?]8796eE+(J-P&3eT8,6
@9.L_BYYXR5SL&1F=9gCfESBAV_5-,<?Ng&Ea_V<c)7<F7]9E&+2g>?2g;+?,+]T
IABF5[9C)=<\YL_4EL_,g#1)e?U8T>_INJCc#\D#dW&?U7MV&)KXTEF8(5#V[:aS
F/M?AOK\6\4\aBZ4C>3B/Hf3LXfP?354U/#N9Jf_X+-#XfX-\^<]3aWdSZ4JcY32
7E5W:Y>]0A;51fNG8[8@,6)<MHV=eECIcODf4K2Ba4:RPA+OOa:c_((.(,f5^.=-
#:U#D?gCaX2E,CM1Pa\gF08P7eX\8\;>WUbLIV(GEQ-+c_SS&#5\^dJI2J>\-/_D
MVF:WIZ2_dccIM#K,-f=BC<RXSM/OV0g^.D6131#+Wg;_U9.QDKa=IQ1O<](ZgRW
]WA6<]00K3-1D6AXTGNI:/T31YB<]E+^ZKY+8@Y4PR><PX?GCWBaY^132Q7a^e\Y
fK#/+Q=88M]DUR4B)g;R]0JdB53V+[de79?4P-AVY@XLJE+/;US0BWX?VOAdIFb]
(]L@),.<b10BC>.:Naf=_VYBe:LRT/9e_:T4A^6[NMYg65;f))C(K&ebMB8?e6Pe
cP-1G4^DN=+88R&&/&;UC8D(:B6T46#+Y>Sd@NZ.70M<7>@DdMGBF9NUe@a@R\Ie
JUb&.(G=/2=)G<L5EM1/^(:K(S=g5W)7(]/#4D4#ITIfTS]4E^F<MM+39DIf(7@C
/0X:&RJQ6S1#?&b?-JZGJ/c>G9F0]UF/S8A>7^3/:N:]P3M_FFZN5DUL=5CagbD(
PRS?NF-LZF/b.VGA-@#ALM/NPfF=dS=>\0AD/Y=(]HCQ2>R500<AE,f3+XF=Q6Q2
3(S@O56[9C]<,L:7>DD0;=#)OISRUV\d,+?J1CU;:<:01.9P+F#Ba9)29\\T6@GZ
L/0)IYKbZGbI-dG\Cae68]f\fBb)K)>-&_,5M[2)H?@bb6(J0EUV7^eWQ#@YLPEH
^6-]e_<>_.(aTFaCKSZ,KN>XDC3^QNPDW[YbHB;W9IK3_VQcV6_,D;L^1W:QECbR
3BdQb:V9\SNCW;-AQ1;YN9CO30/N.G^C,>-.g_+\@831KQMCV,5[:/O,=S8]CO?L
J/\;cFbKA;eF8]B34AIU\F,JVVTf^QbS)gPBWW?SEP>OB5,?L)HdZ\P[-X.WB6.E
N7\\H5K]A4RT+&S88T>;=+?5[0DZKZ3Z/BUGFR_=.E.&/deQ[BSRfaXLSeYcgYU0
POU8S9@@ZT_O7^)^ZCNTK.Zde4W,c=Q.T/.;c.T9J(IG(Y?YVU<7_D7AZf@KL=d]
>]N2fBWSXb23W?5g3>G?#dVK573-^/)^2RMaQU6EDWeNUC&?Hg_<(:eQe@gHVJZR
WOX3)NB8ASJFF74I(N[Q^ID87:^IOY6T8G6U^Z5_aXOfaIF.-E7_1_aPcDZ>N?ZP
F?[E-P?fP9PW5OF@cSKAN+2J^L\2PE8fOR9F0+MS7NW)\R=<G_.].-:aG:B<eb[5U$
`endprotected
  

`ifdef SVT_VMM_TECHNOLOGY
`svt_vmm_data_new(svt_ahb_bus_configuration)
  extern function new (vmm_log log = null);
`else
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new configuration instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the configuration
   */
  extern function new (string name = "svt_ahb_bus_configuration");
`endif
    
 // ****************************************************************************
 //   SVT shorthand macros 
 // ****************************************************************************

  `svt_data_member_begin(svt_ahb_bus_configuration)
    `svt_field_object(sys_cfg,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE,`SVT_HOW_REF)
    `svt_field_enum(ahb_interface_type_enum, ahb_interface_type, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_int(bus_id, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(bus_control_huser_enable, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_BIN)
    `svt_field_int(bus_extended_mem_enable, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_BIN)
    `svt_field_int(bus_secure_enable, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_BIN)
    `svt_field_int(bus_data_huser_enable, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_BIN)
    `svt_field_enum(idle_val_enum, bus_addr_idle_value, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_enum(idle_val_enum, bus_data_idle_value, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_enum(idle_val_enum, bus_control_idle_value, `SVT_NOCOPY|`SVT_ALL_ON)
    `svt_field_int(bus_addr_width, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(bus_data_width, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(num_bus_masters, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(num_bus_slaves, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(bus_control_huser_width, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(bus_data_huser_width, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_DEC)
    `svt_field_int(protocol_checks_enable, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_BIN)
    `svt_field_int(ebt_enable, `SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
    `svt_field_array_int(num_ebt_cycles, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_DEC)
    `svt_field_array_int(num_mask_grant_cycles_after_ebt, `SVT_NOCOPY|`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_DEC)
  `svt_data_member_end(svt_ahb_bus_configuration)

  /**
   * Assigns a system interface to this configuration.
   *
   * @param ahb_bus_if Interface for the AHB system
   */
  extern function void set_bus_if(AHB_IF ahb_bus_if);  

  
/** @cond PRIVATE */  
  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();
/** @endcond*/
 
 /**
   * Turns ON or OFF all of the "reasonable" randomize constraints for this
   * class.  Note that "valid_ranges" constraint is not disabled.  This method
   * returns -1 if it fails.    
   */
  extern virtual function int reasonable_constraint_mode(bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Method to turn static config param randomization on/off as a block.
   */
  extern virtual function int static_rand_mode(bit on_off);


/** @cond PRIVATE */  
`ifndef SVT_VMM_TECHNOLOGY
 // ---------------------------------------------------------------------------
 /** Extend the copy routine to copy the virtual interface */
 extern virtual function void do_copy(`SVT_XVM(object) rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);


  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);
 // ---------------------------------------------------------------------------
  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif

  //----------------------------------------------------------------------------
  // Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to);
  //----------------------------------------------------------------------------
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
    * Does basic validation of the object contents.
    */
  extern virtual function bit do_is_valid ( bit silent = 1,int kind = RELEVANT);
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);
  // ---------------------------------------------------------------------------
  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort. 
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

`ifndef SVT_VMM_TECHNOLOGY 
  // ---------------------------------------------------------------------------
  /**
   * This method returns the mahbmum packer bytes value required by the AHB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the AHB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif
/** @endcond*/

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_ahb_bus_configuration)
  `vmm_class_factory(svt_ahb_bus_configuration)
`endif   

endclass

// -----------------------------------------------------------------------------

/**
Utility method definition for the svt_ahb_bus_configuration class

*/

`protected
,S/CeKPA3THf5SK>QG&?4^;5#?cMPQN5[M:8_F=fE:)#@7TGQF@M0)HJ(^gLW5\_
CA:64X0a-\#bVC#F?]:HN0DZHMb7XeQD(1(TFY]2+1ZMKHdF4+=6C6G^?0c@<[U=
M(60:54RH+C&KedXTZH<NdK]_GQA<8fKVC[G^5E;D]VLR,H,R=VW0<Z,5D7F/T9e
BU8.YFO,&?gBY[JCKZb]U?56&-^Ze#bb8#-#f0N/RFR-764bf=H9Ucb>OO6^4@F?
dMS+8AKBJ-ePFA/UTM873=WCD4R#eC8KK1aW/^g&/=_H4R8TY,L<GDe/SH<7AAQ>
Q@FF)H---_gS7FOMX3>L[.[bTEJ8[F#eGD#TA+=C\QGV&S6^I;c]2VM;B&#PIB9=
DMP8_?1N7F5HT-IQ=Jd=D#LVW3,dN-F(g@YLA[6J83AK\^GKHDGTVF?#YBC4f9AA
1I_>B&#5K_D_P#A&9?fQ&H>7^G(X7+?I6P=V0;6XF7/7ZN.g(f5:8,G^HHJf])9U
#OHEebad@MdRb.<4f=^^&C>73$
`endprotected


//vcs_vip_protect
`protected
JH.PdeO;Y&LRRB#f0A2E\K+_bZLT1X-4#9c3g]/g9T&\4SNeRHMP+(+91FCD,cfF
bU3(L@OgJHH[O7;Q8V?H@96]=425La;&>M8;916d+\;4/=A9.GP+.,^JDO]b4=(7
-S>WJd>a.ZGT?&@<UZ.4TC.C=A]5)>8209.+/Wf19>RC_dY_;O6M-[KLc-X?[:3H
YWIb><I8:520+]cU1g7>5B3E0O^G;KCD=UgU+[ca\24dMb5]-cBVcHECeJ\F8U_5
OW.bN7\YO5UP#2(eEXHAbWa5J9>eSXG&J<ZAbIg1-LP-;I81F);AHaI@8868E]UM
3;Y-ISdIbd=g,f/bbO#UfJ7=0CX?@[N7==YV?=GD7=]NLbL>e/)d-fV-R-IY<USY
;4(:dc<^9JGN^SBL_g]<E#FLE2.M7aZ.cP:E^9+3,<D->>1BYA(W-R+LWEF34N8Y
\80Xb,,-=EdINOHCXf);ROFRPW9gLVNU7@22;GM4R(2H6E3&bX6;B&N\.gX[](97
X#H6-SI]5O339YD?e9;g#K;0aWS9+)E\H=8C_RVaSRQK2b]<,bR?>O1V9_E:-7#7
9OGMHY3F(HMUJ2-V;5Sgd_<[8V<N@YCb+[R5^I7=0=(\\FQH,M]?>RSN?P:M451^
[8c(;7=AZa<\KgfW&-38+<G93X-VafW;KT67F,37O9.&,ZDe2HC1>aYH>6F3V@IR
3WH;[LL?U[5@&KB].BPQW0&(=E2TDO]54--eZ(NN+\P7;]gI>[[<-&K4]1PaNTHQ
G-2L3dVX5J5dU&+<\^[V<=:&P+ZGDC7B[6(]S0USA01I529STR+Q(ZQT#MMI:TVT
&1<J9Y5])JW0+LI0:>ZAMG^3Jg:\S3Q1G^1UMcGDW_&ZD+PB^eVDN2F9XN:V:RSH
Q3<\7-c8-3BbXW2(5L8Q@Fb#9-\[<OD\L=RWafPX77CfI001.4D(;<A-\(E&F]Gd
KM=aY?O#O6SSY&a.KM]_bE_JTbSL<#R50:#3AfU.^,Q^N8@;UYE8IAgEMa]?S7YN
cFA]ZgZ<H2K2bCb?KR_5UV,Ncf140FK6/3;K;\A?f=b9-9YJ.0,EGPQ:^&2<39B5
J]CG&V.f.d2A0Q[@f;6>(1@,aU\UMMYbfY4E/C;eFOR9-TP;J<,D0^[LMg7eRgNY
gBRKY[0RgHC-N99WQH>-_0WA<3E&.\6.DR_8;/=4F8#0ZR0:R3PVF@);,V8J&K13
+B^6G+:.20fDNebSf_;.WOG_&ZN:N<Jf^NP<)NO.]^V[<&<KI)X(fNfT[/O7e^G5
d]_67Z)<?ZHIK-L>\Af9[a[T#2Ld68YSfYbbMIHZKL,KYgd0cgD)BT(gZ\T@]NdX
4eS,7OagIa);Md(ScC\F/LPABEDb6:&d)6TO;JR>LFF#L8#0b)J.?8[X8F0;NbOV
J?.dbDfZ<5##Z=.Y+/_R50>,CNE#,>BPe^cPXDgSZ_[7O/,H]eE,\W\^5++N[-#(
TFLB<G.7?ZB5_L)#]X]N.ZWBF,+FIZ:eFBY&2eF[]7gg_[]5T722:EcbDO[PDHZe
4_V8R?:_SN^c2GCCWS4HK5();A8[fa3;3X/T\E=c[eN^Ka?(7,/.8U??[Z9<+\?c
3_]_ce@I/7TaEW<C7)a0J0PB5b^.M(K\b(VSVTV3:;WWIJeKd4d3=(C^X,N4CBMX
(5D)Vc0#=2GU3.;\J+Q6)(M\/QNHMQ4\S]DGET9IML4:?KHCM5T>-:1&OCA/7TT<
-DYg5Q)\8fBfPX1c2,GL[.8ZW7V(TMf?0e&TJd/L/[DVV>TBd/]Z^#BQe9YM+GY7
^b?SO:;F8dFFDecOf];=.1G?FN:KaGI+g=G-R[3RI),@-I>?3,:FTbM1B\#7B1eg
\18T9@99B-OF:CeA=IW,D0b[^1([&(<>H^KWfYN4I[2D@27&QY,PG9NcDX^B&gY6
QgS?Q;b.gF&E[>-<b15S^ab3)bDFL=9&T0]N7c?2bYEe@9A7-#1F=(B;?)NU.3C]
YFZcD3EKEL/I34WEfFLF>A.3ROOW-g)VcJcDWCfBNN-D>)Fg23G8;IQCA3X@AGI#
dK.LE-H9Jf8_Be@,(&U#0;.FX5/aESY-O9^(8ZXN8-]M6(0L]V9V4B::c&41[@/c
THUBX^8525\;@R2T0Y):IU2ODDTQD:-D/7+eB2gQMPd4<d[fAPaYW[\g(+)NW/5Q
9GOPPSbgPdSYB3d28033LM-UgZ)I&S_EF_^_/NAf;\7AcWQ8O-;]+CTKFTC=Sf;5
BHDSO80L,Xa3ER@89bPB(<:Ef<ST=[fV4#a&G:GFHKE\UZ28&dc[f9XWU,^g@<];
#2fU92eb4d(:E;,aPIGYX7O3M?;=CNO=c/WB>@K<N63L]<.9M.B@+WY#1CZXX:^T
P,5P?JMB,Cc(/+-I)08Z\g^c,fd-1]K<7PfSPeO],#I:7TNZR40Q:3LK<JS6[W0>
T8d\N(J\<cg]ZYdc41_XbARW1gVc_P71M68_V]@OB+<&WZ>KcDR@+c5ff@XVK7CJ
-D=H,Gg@PQ.1)e^e&?X8R8RZ.UA4a1-9MEfTYVFW,HT^Z0b3HM3G=I4,].eNS;0O
S,c@3c;?L>N30V&G)DO_f3@Z3T-,T5A?Ub+U;7?KP;c4ddK:WfD[B6R52\DIcJfB
_:8Pb,S7eU16]H.-02?f@O1b#8L^Q.H&O+CJMc)dd7XM:+JGDYS55N^TAURUXGMN
OK>V]NMR#FY382#/A>UL9K\G168TWY[]+G=Ic>JeY84C14A3QT=bQ^LN[/5K.^N<
DCQH/5=9^M&Se,e;U^=:5:CeF?VP-SEQdf5W)7O798<\5-<?_GC3PATFE-]BF+<\
-<_F/((4CQ/V4^HM/.7Ca=1DSEV9WSFc:GPM&[VG[ISgI75L>HB&7g75S?]D69L)
NTc82)f&B:19H<C=4G#0]]eI[L6:WcXF>Dg_9@H44EaKRDZ23[UBC-,+IY>5_[^8
:d.36WOX.9,^af,P?-R,QP7W)#WS^MVbfU8\Q(+5@fU4T1a=UR71^:E?=>cb\HP.
N;g-?S=;:YE?4:JW@A@#Ob:;6KSY8^WQ-Qd\B]U<#CEJ8_D<QgPWK441OSc^4]?:
G3:LMWD9VNM1AZP&4PMF863@7#IKLOM<957edW>46H18JGFKa]CF::\cGUJ<UNU5
\J9Tc=:?#;cab[@c72KfXPWY0VX3?caX+X.ZL#GP0#+<WQ+RgBbQ+8QJXF)U9<OJ
B.MF3SG@d0O.X#,BE0&>[>T,A5QV8M<+)[b?=>^=?HRW0I1F5G.T-F1[#P1<R9M5
46f=EaCB_\]5D+\J[gM.CGI4e0/\@[8SL1R0,XT6DMQ93,C9-1GM..WN\/,(Ae;c
Y3Ca&QI>V9/B?WRWBfHBB2U_Y@X:L\)Cd?V9Q([;AT(CQ^4bA-g\+4<OTT#a:JdQ
DHfY#@TX,WE3P3(b4@C_e5V&AN9:N:Q]KL/].U?O6bVagEJSe&Q2EQ??+_BH).MA
EFfJYJGSDZ0-R)8/O.^[VeHdU=AOPa@T0VR^7QK+YdQL3STOcI5-^KQ8g?L;4I9<
c/_5_W3WK@Q0.K[BZPXK,eGHU,I(ecSVgSF[:<6Yd4CJ=^_&N\Q[IO#/,LCX2U]F
2RF&033-AcIC;Od)_8=NIgRH7JC[V:aPcVYFeG:43fZ=C[9[gU@163JX\35c09MA
EgX5:TH.0\VRH^C--W#dKg3-U>Bb+ELY9GE0.fF0HF^.c8F01@<QT\[S>EDT\.\?
>_>f95PN&A#d8TTa6<RZX)>H]3]Z\L/fZ=G&DQACPa8dY3eRXZ?N];)\YfZ<gHA0
3-M,JQ2R7WR:Q(,U?&9;>U#Sc?@TcbKY\S[5S8/^e489K?Cc>.-1+/.V[<]2aB.S
8]eWVTef.1[F2?-LCCAZW4#]J>,:M-/=aIA42b<,]aWKb=&3(a\AJ36[MA(D46DJ
GFZ>2_GgdNM^BOV(79E[=c?FRBK4ONQ;d]4ZF:@b0_<E5gM5_>[>[bH#U+N&-Z43
NKMC^3c11^,W>f29c97QSQ29B[MJOcGC9=Y)Q(Ra;@@/_\6-?3G>LWQ1,0;@5,]X
YW-F/G94E-JORSV0aNFe[1&:9/V>g20SR[NJ+9?/a_(dL,XF#/bJ9e_[1cf?F;AX
E8IQ(\,6[b>?F=0D-DAC>B0eH:)@9Q.<.RG(=2P1X./1fcR47UM]MLQ+@5I2@H7B
,f:\^<P4c-5N1;5BB[dY4AV42ODJ/=+)^.:([EA#V8I,)<_PR/9=Od#I<8K=HfYJ
79)&#d7JZ6-bfXQD1X9&7@)<IP#Q=00g;1g14#0@PJa91JPOgVBI4.:BN2@fVM:W
8dfaD_FE(:A?\LF4U@[8TR1V,O8HO#IRJ.6EPgMZTX-,A49@+D7&,.S,5KE<K0.J
/@:4@Mg>CRJG]OdZZL=XER1/;NJE1Ma,WdW#S)/_Q0705;JAG-6<<afJAeTCF),Q
26A<.eZ1e9>G\a660O-=K?J3EOPg8:Jf9CIfLd@O-C<.>HZ1LF3D/@MN\_,U^\6^
CbT,EKc/FUBV&J?HGR3cF9g.,5YAUUdT7_&2A9D<-)DP[5JLMAaRZ-_337C1I\6S
H5P:e2+H6QJMPf=,E2417E&fAT,McCRfZBK?5+5(QK.&4Pa(6JMb,LM=aQDWIFT6
0f5f-Z#N)DY=V#Oe5=RD)6)e/&:2#e8NeB+S;DG[c^\8;:9Q&4e^1)0X\&/\dOE=
;=9ec\-44:]45GPOE:;?Q41:0;PDbTL:>299CaZUHKVD[dUIMWA;d[H,CZ6/^M^2
])((_adb:584(9:2#_];B679VfERDN1C7/b2]4X.CN9(K49338RIME#K=0Y9:=7M
SG+NRK1094_B-g#S?=7ADL>4WR.Qe?[Z5M[21&D]91Ad1:Af&=+NF.bE.?3dA:5E
KV)X5U.7#VI6Ga999I\&V<W?B/_A4/5,O?RIMKaWH?;>2.6_YULC:<(3]M0+8;6E
.&E&(:#WGHc)35a1TZC8QS0(1W>=\.1?Y2X=N]d,>R/+^[R]4cUdT@J_a;dBZQ;b
RF0;c+-aGR9:ZCV0A@+8/^Xa9K@X/H&5B;]e1H#W6F+_c+2_d3RD>)d8T6M&T+Ad
cYLO/<R=X=bP@3EK(aHbEK3?=R80=0A&K8151[ME5&Q<GY_Yd537JPGcMV57I.CB
e@&.#GI<CGJ#?WWKYg6-J&D8:QF8VX^@Te2\[GD;F7<LD-(&2Y]fZ^\.K@U\^.6)
]Mb5=QYI?=d9E139:S>b68IAPVP_;g&0&I,1V5U/<)\28cFIBK6HbKFFH_Q=eR+2
#]\a^R(d(QJDaJ^YB0AT7Cc:126@3SC,R5#-3LdKH]ER0bI?08+;4.<Ea_,;K]/;
YSOS60=.P3D_DMU6APZW(O(JH9f&&4LOLY6M8E5/\&[dV,&HeMec673CTWe_RF(^
RM?9BX>DLEf78^HXPVW;[.gQRA;]3+\\:BSM@:a8c@=12P=C2LD@I]45bGWIc]^B
48d.=5gSdGCMF\N9.QBZI<P;f0ZgGZ3fg<7KD(R&2bZ\.XYW)I1Ncd7b8+/Y-KC)
#?@6RBCT@0]J;XX7CA4)R+/O^N-I)Ff0,Q+LK+OXc)QF<A&JE2a\0T.3+)#=954b
>D;W<&&=W)#ggKY?NN;=Jb6+8,D.ffe,:=E##AeCX7?U@4+d?N&Vb@HTf0M_>\d4
/a^=Y>_9HOaPY/R/WEf]B8]9H0<G9V7<Q^:)Id58=<T/b:<-AB..?DKQQ-=@<1Wf
O0E2ICK+gFQ899cEZb9GFBZI#<A>&,aRCcbN)G\2KHI;d.PW5B8e3000I;@NGdcE
5GN>5@KG,c0P.F#c@R^c#eV0N2f6AL4b]^Z^a9=B6AYA^1/E\9.35S60YVJVNA7:
=F#05+c1HCaC_fCF8aSWY4(N7@D0dc<Gbae#D5HYR@d0<GDPS>#^d1Hd>W&A]eUJ
3de/RQVE2@OgW\LL6RI[d\,U];XaI#JFF4Zf1>:N7=/SY5b4eJGD=HP1LbcEDKUG
a2=R48I2[bA:?Ud[X/=aYZdg3&]9YUgH:7=R7(9M;-\4.S)B0bfI)#I4O7/(O:&+
e/SVN80KbLFO-/>ece:J2+[b\BfYE=;TW90e,e#C:E8?KT@T3dZ185^0DASA&dYJ
(>H45T2L.L248gV4B+WEJ(gTTbQE:QJd&J)K.U6/DVM5U4V@GOKNUQe-:Y&MGQbW
d1#ZW#F4FZEX@V#?(^0,SKN+3+8FT4JdgZ85R5?5/.:;<8SaC+_\QbYC.DXgRGPF
&ab]d_7VgR>H\&aP0M5\N@L78H;P)?-1Q?X(bNKGM2-ZKbQMgX6S@-6aPWCD3fHN
f^KcVE[)730NV;TB=95TJNI[-3#=&aaP)G)9-A^1TSO0,e:?B9;]21SU[1@K3=69
0/F^_=@LPL/7g2[GCdKGP3+;\G&ZIYGC_?#-3ER1gegUV9D;.7_7Z&7(ZZ#RQ#c3
<g1?Z23R>2:87QE.AR<E\@7)ZR1WIN+T45]?eO)(1\R\#5YM1a&N.FM??D-DgAc;
E9QZJJ@;=NB-+8G5MVPL?6?U95^VF5FHFMb]KC/9Pd;bF2>X@^GN^G=/1(V/FM70
85J#_7;;RYVWF2fW^R1?^TZ2KU)dO9^#_(#61EY]P2CG6^.CK3A=K:?3_\28-G<3
SS00^.;ceLLbRUcM@f-GU+g3\42TgXUAXKH&N1#W6e_?@7+XQca2P@I)5?MJ(/E@
cP[>gVB53O6X/-C]@Kd8&gN-<4d/XEf5KC@V<QdgR6+18Z0>0f_QW@^BO\N/)JAO
A]Y:#<OOgc614@#N>/&OK=/KV)8Y+:-11GY@,0GZEHL1-&KZX/g7.K(X@FZ<,VM#
fGZA:XNB-HCcL4P&gPEP>_ZP_PYP](cL/UFG9ae2Q<D4_7MG,8G2f4^UTT]BBc3Z
9?.f8Z>IF=N7HVfKc/YE:af+6Z&I(<50:W0AKNHF,^A0=UDeOgVZ/&88>V2cBT/2
(+@S2P&EBYed(1<R/e53:,f0L,?JT<\gTY65]4fPR[+aOgfZa36KI+RE,E(;fQ&H
IBK04QMIZ^R=G\CI04L+?U96:89>0>NHBXX&S@P74S?b#4Y;\EF4g[D9LBVC3C14
/DGC?QK7[+)#PWOCd?7Q0Y^HF)0;EY_AA5bRQ?[JI7EC/Y[RZ)C;^8&TMJPYU)ag
D&)dZ#MN^=g2fQLDT)S0WWO^3CRF1[Q+0.a8@7RG67W@#F;0&&S5I:X9DeAC,1VF
Q7=ZVU/;,ADDU.De\OWbb.==5f27?;LW#;aYfOHTd5,1bHdAd4&VT,VHDC^cd9?I
aR7+3KX8Q16CT6SEe2)W&P&8Ta7;#V24<8:.8L]FVeAc3?#8X+L3E]SLEJb7BN/W
2<bXWH&E2M#[T90g=Q2#_9ZIMY#V]@X#;/1&-Sfb]5e8L,L#SGLMHI=7.(>]M6WZ
E_<H2Q]K]2)S?;VY0L:_CZ<a2aQ05a\M6_A_&MW3?aDRFLJFa3MVd;aRdKe-0M+4
XTBWY]/H=ZMb55g0)60FY\Jg[&R54Dab5VK?HGcMg:Ic0,C2LbKP;OV8E0cU,KXL
+ae<f-FMdO3@94R(aI=\@67<UTAO:GA?3L=_cW;?eS#Wd\VcM,;bcFCF0IRIK.B4
4^b,;.b<1^0=?B<:.K;8:gA@W=L]b]Z=3e(bAL<MVfgVYBZa.J=50<>.7QX(58+9
0cC+cX9>G6/80:aZa;Web.1PN&ba1389RaJZeWd6&3FN#Rce;J_E:XO>^3;OLIT@
e6..8+<T&S4Eb-,P)K=[1+b\]e0QdPQ5I:?(TV@HKV4YNY1O19M4][BI>V07aa&9
MO_QC:I6\O09>GWVcE=)-eIQ^9Lg56220D8#AgP7W9-\EZT9_<0IC(c=L-0:=6g.
:?[9,DTgZ5b>X8b\EHD=WA;ZIc0bPIG9:[0ZY^^AD[&TO[ZEg93\R[-Md6-JHSH#
IeV]<F]?EOWU.\?@-&F\H4<O(?:=9dY5RMg,c<M6T00L,MOIT14B>K&&QZ#eM\&B
#b@-f>N@LK4\1XEA3]H3V[DfX<S=3YM504RM4g4eGH0\P.+9B^,WSLNWafX5#S9:
=YEeU>P:0Q#ENdda80K,OG=[eCFH6e,b85gL[H;K<SCHd1Z:\4V?)A-(a9OFH15d
B\8]\2>&[;,R7T+PcNX.V8,EJ&B_U2cBJA)aMfU\_bMDB@M4DOHUVOHd\(Z7.]CU
_bRHBU:]NI)gb.#5WWDS>N2V))BFKUQ\+.U7X&>U8Te6C321<+(USf2L+<16>2(5
+0EW<@\J(B^RI,L-cb&^BA1T<TPD=T^?_:g76<;e-e+UaUR((CCB[SE[VS_^@:.d
G1YPd^S@0;5?Fe491<_=(_5TJO2-LYBMQ]P-+>ZGB&&5[_1/.0?B3QL#F9LbUMaL
Md0eM:6W0,0F^G3fbR0R(DL?U-7/@&g..@CD),DCfb,8_Y-RY4fMU_9Y(K+3IV/]
\eS6TA:DO;5N[SVFP1JNQ]SO^a7c7Bc_9MH/(D6S+.K_P@\MMdINJfQSFZ@XE-bP
8X#02>5OI#?1(<PCS2&V<IRS3U;B[G,>UI[\S[QU_M&D;[3&X3/IG,WLfDb(_gZ@
2;70Y,4GWcbc+(\(AUMWQN70d9C-(VHD+#<??BW<a]YQ3]+K5/MZ5)<CL#-Q=Y<.
6.#OJP^J3<=L_ZBD]G3[.SPB4&6E0,(&#f6VX^ZTH/[05AMcTNU<Rg-70JVDdc-#
)d.c_a3#WTJTSEN1)e.-9a4,Y4#U3b?534Kc)=SJg=GN>9/&<;:6c1.SbWRX4aK3
8OB6QM3MbLdFQB](4g,N4fM9(L6CPU\)#P(SSAY1R2G/2+M1PV(9\95@MKd0PDW+
)>TH#EN=DNBB5?)V0(GQeS=Gf=MOY:\2-D^1UA^L7]+6?JZLF/_/U84M@?#,D&Z<
<Ic0-?HAB\0FU54QgQMX-4^-Jc)]d/NS]N98)^+_8H<V25\J_H93G#e\:5WMb/_3
0Ofb[&WQ8YH(G9Hf<a<?c3Ke23Q/f#.e23>gg/cL+1N[R3BV\cUSKU[f9SaIb;W.
&=LZNU3Og+J1HR-R[#EbQII#RWC:JI;<VZe_:+aNH65I2-@@_e.43/TFLB465PZF
Q,dcAYYUUM[Y>^B@A+aWFTGY:gDMGA]N7_aA0g6S9F/9a9TXPP08dSH]bI8W#RH)
a/DX<JSY-WO3^TV;c\<T8ZPdCPd6[D8.\0QSf5A97Z]aWW_KM55YK[C:1].YC.dM
eX.Z]3-J@5B,;ZS;>BU3T?Lbfa9>LJW0W<8EaU=6+M()KP]1B+]Y15g>0Q@7_/.B
#EGP)V5g>CT57#.f4F]X9Y2d]T1TGB/.3W=<dYML/geT-0TGX<^,;]@7)=XG:;EX
ODQMOZaS_aBZPLf3>B4SIU+1-ZPE98T2aCGA;YV;?==]2O[cLWJ?aTS<_P_^d31\
dfN6Ia?LMLZYLICXVJ/_4=/4<QfB)>B.EQ0<UL.QSR,F9R8G:6G4f:?]_7Y1HV2I
BHF@2)0N-1+<AFTa6^3a.H+b\gbO/6G>@M\0>FO+5&OI6OMA@>AGAE/^g#/+CL9M
2g6L:23(#M3gcNeGUF\FYH2P0X&F69F4G3U<aYF41P]a[c,)aDbSfEb&,W>LH3e^
6XcV1X=S6B=W/=>8X9:B1U,/KQ(eLDGKZ;U=cbK4AGVFR]36114?1b/NXHK?1PA,
(3d:S252.I[QHa<Fa-\_@7ZCB;f@)4=cCSG3O]C&@NFf#LVTfIa#)dQ<PPE^OAXH
.+V&?#QSGL)Mf)e0G5K+T41#;^D3Z,f^^GR#\(<,>a3E:@VdBc1B^cbWO9R^AYec
525(=,HCZMO11b/#PMAe,?N#/^7?UOPbA,/T8:_Lc2KaHGDc>,GI.D=<g.L\Za(3
O)c3Y#WOY#F]A3&Sc(PgJU4[>Z5_.(S/>/eH(XN.[1cOd4HfI+X85Nb.CJ#<N5NW
[dNO4=5BgF3f=H,YNV#-->HIe_#NOJIYRd?a]?WN4&H)#>aV.9;NQ\JLE+)dfGYI
DX7dNF[1;Mdf3cgCag7)#e.75e<;586UL4WPP4D-\?EATL-VI-Y^]LQ4/N:>L?A,
<SdC:gePRdK)6(0eBO_V5J<])\^;JYRc+d3a0EB<D+T>PAf&TPX.#5J=>AXdEIa@
+.[VI33<^Ie_H))SH#D_<2fR0fe#X7LcFP@72R12.+:D2d.&B;UI.RH6I7^NR_3J
a+&cC^OW6gg?c1Sg([0HdK42[_TM#H5IF#)+0f1DQ;bgKW0&fWN<WJ26bB-D4/dM
7@@[+bGU3KI51+e=O@V+dd1+DgP,T<:F,IM>(.Pa.SO>;<QKgE6;GXQ5DAP-:&NG
@cfS;8,ROR77F\dZa0FIa,&+X)C8d,VbF>NQME5BLM]XNdPA9YDc27>,/AcLX+_3
,\L)ecKN7Y_a=[1dR#VbcJ]RYEA2/)HLRb10K:=6N;^R[R+(BM<N6#a0UKg<YQHQ
Y<;Yf.fV(R(=ZdCS8LK-=H9AY7QTK0\.;6Yg@F4)CWdTbFV\)9.=I973&_e_fVCC
(4^Vc8f(6Lg0+@bO&395-X4Y14R2ad&#:DQZHLV)@#6Lcb;G=5C_Ib&X5G\+=[CL
J^I38.R4PTDYE;4QO/]GPS[THga5c6Y4];5FLGW:ZJ6EW19aW?BKO<<aFFYWSL+F
HbYcaLQ8)U/U[-BBV9F48/)7SC#G8+W^3,UbRQ5:;ceGW)7STKBG]X.XNB[(fPN-
/>f1W+G5<BWcAX8g;EU[^[PD)cU)]HK_[>1cG\^fMHBT)M(97Z:=R3NRD^fF&<IH
b1T,^[UQ,e>=?cc#R:HL&7.1F.5WDc#P4AT@]<8S3JK2MgDSK^+,5F-@fFN0YVP;
>XMbb<<+?MZd(Y(K2J@B^>Q&>]YSSEG4?d??L^NbJ_cI9EZ98c+K-1S2U[^ADHYG
a2Q,_V\M\O,L[cf8eHB(gL.N^D5e_WH4[@Q]_Y->8J@=,95T9MSA,8/gCX@ENfg_
DfeV4/BHH>-6;SEGPB,L4QG-U2@&Y(Y_<c>H#US]T?J?/-]/bCg>X5XQ[MHCK6TL
UY[?=/E9-S[]Y#Q^T7QJI.DeUc6XO+KY@AI&VK>Q#b<<CAE^P72QWb3B<_Q<-J[^
AK-?ZOe,;gA5=d=/_WJaFg#TaVT-JTO(OZU:K[DU>AG]#f,-P:Y(X1YA;C@.[a(^
aP9(F/2<<=)@g215eg<ZbWQ+W#[R;e2,&L)^WR0JAd5a1VcgGZ7HG(gHE^CHR.P4
/bC\DA:<Y,8LY0OD.@BO27Q1UDZ;#TOMXG:^HC3FgT^2=QM\OF9MZ1J)X?R\Vb\-
L2342BR,:MK1c5Ofe5(X^(/;E,5S.?U_Ta;5G_]K<O[FcK4><f/b=:@F+Yg=&SQK
I#3ZW)31TAT-;C7\b?E.0F#cU:&eV+D0TEI3C;_PY,0SYCMX<?>ZHTQF#;DdLW@)
WJ6&=9B=2Y;d-S->#)C,:f77^9H/;RSe;3<I\;@R51JMBJAcNRe6D[-N=cE<&Iab
R)&_GF#OL])3B#d7IeW/URZ1,YRJ5W801,M#D(HHK_(HYbI1D\a-=H5S\&[B7Vd_
EeQb/:-[(K31gK0bdQSZ)XbGKSK62G.b.P>[;-87N_9d/8X7Hd1Z&O2AC\d-LbHg
HS?B_/<T2E]D\UO-b.3<f?LA/1M\TNc^/:OINCg2114BUS:&3UY8/W92UeSgO)S/
.JTA@&1&YF#]M?RA8]&)<C22+a/6D\&NIA^WP;G9cU8aU><NSU]);4,aE]6[;EBI
\d@Na5UCK@9:[V<-P77&P?-#X:.SYR<0K/F@?)V[a<?d)Cb8cf\CDbHR>=O8GP(f
;0eYWJc)?^4aTL0F0O_#8/5<1.bAeZcJ.RVTf^;QO;]MHL8V-T6K#d#&K,+&[C7d
^MgV,F;7,U-4F1V6>eSfRgf9Z=.3EJOD;gM2AfG5T5DAb)VAGN?D?0,>6[e_XEXD
VSS@/F9Qg.6)0?7??fa_b8P-S-\U19A\:SA?^fegO^SGa\c=@a^1HH[ZVE^9gc&Y
7)^73K:/;>:>gU[:E=N<DN<;/OJ:E;XSa:P#6A\PK(H0_DSG0S&+LL[d8OcMAISY
8?3:\-L6FWBTO@_CE:E^+6dXYJ=1IQ\(X\N=3+85MS12eeY8OC5AIF@89>109>Ue
EfUaE[>++,N8X7CL6]Z15;F+R&&C&5MS\Z=?&ETa0c+<8\2D,2^\9aBH48,.7(I-
-QJ?KJX^<:,&OJ5#<PO73\12@+L2Bd>D2Y+A3Z5Z;G&>YD&)^.CR3A=ef@C]_eK>
.&U+<]@7;IJAR>/a69>b5<NUR+TVDO90NS(f+>FLJ8TD(DDB<YaB]WF@^9\EKA)f
5VfP0b8M78=9@NZ[8<+V0L?2WM)fa+1@e)L;PC^24Ib/>d.0D/e^XDT1Qb:RH5e7
+=afZ_9+QE1+S5O18C^0<486fCN>:a64Bg=?ZGDZ&G8,_[X_W<W7S?OK@U=P3D=J
d0ZHfAS_H&Xf0.:B9#Y#WFc8(X]V;OC?TKB]L@cRfE[:ZdW0VZ-T=\TWLZT09I@I
bUJSWET<ZQ]P(2HD=JPQ^>ST(V0W9VZ^JO32g96<H8EC-=e@@Oc[G=aO[^fWZ1Jc
/O\JIF8ZD\HGHBcPfMQV9C5N8)VT+Q5)\f8E;B.&V/0eGO\g-dU7C/?C2G_=f)J0
2<8LS.J:_NHHM<c-S0VbRB++)W;ee]Z]Oa[C&3Y]9\Q9R:U]REE-I1:L&8;2I\JJ
OQGHPUQ49AI2OQOBc+[aYPC_TeA^2UI)_O@8)3PFC=^:Fa1M?cABCXW@.a<ef.8_
5IW<<3L0A<YT?O^X^_cU.4<g2A:<4E\b0BOS>?&X)N+L0HHVZ:aZeUSL:.3:++^a
g9d:&Y^bT_0gM/SC^F[G\+U=0=J71&S(e&#GgA8+JRLg@D=aC@CSJ,d=JH_3HQN1
X).O6^<(A@WZ^.c(L1Mb5E^<:ZTE[?YCR+bC7Y]<^<T_[_=9WbL3YZ4]14LDFDaR
;-[^<)eJTV0)P1WA:,-g.NM[2.<d3Bd4b&c=,6?b@AKM(^N\W\H]Ce4CgUHP#Z.>
+?XZbO=S=##S8PRU2Y<=IRGUQgE,+SY=0POF:Q5CXOCTK[^D5d3U/L,d+T;HM3X=
QR-0\Z^fJZOCeB1>ALKQUC/A:6K#L8cT4Z:U\Q95H@NN<BcRQ\.2(Q?7)^226QMN
<SZ[dL2);18\I;,&SeFXUV+L1>GH91Y5B(V<X>B+b:>9:0DQPEYc;_92?CQRW[4]
7(dXQL9caTFbbO+3FX^M/@e8eg;4-F0O=2?Q5eGUJ98]7aQ=T81^bQce/>C-L-Y7
OaIeTVgQY8N(ff#X8)#JC?9DY>CSDFL,f#-6bJAaJW=eY]I5XdYZ?\)[GcELX<8Z
_K:_=f^1=g41\e&O/=+,_5CV&_a7C@Z39KH+?#J:eIc>#F35\:HH7cUZ3Nb.E2UI
ZI[<Bd&c1)7_8IW7ge9a-81NMU<IfO4f:b9T5A+&@f_gQ3@<8G-MJQ=dC?WL9^e;
RF2T0YA<Ma-M>>S6^Fc3HR=+.A;IQ9/P3]J;bKg<7ZR,b722e2+CdAeRZ2M8,GD0
>KEE#B6N>.7,SAJ>95aS\Z<Q\4(S<,8c#W/VJ=N9N.SYZ.@YIY-T0R+AfK:EA7A7
:&U(4+)TXP<#g5:JHe+UC<\f=EFSYQCWWTdX=_O4d:-#6:SISaM\D:3<QDcOg.Sf
4>:B^^0S5KYJ6d>;<,UNW.gAT+3HVZ&+)T;V4^?d59ON6IacFWF=Z1/C8ZOd8MW;
Y=O>LFFf(SY(f9bS7[:E,L&],3eB=MXN1V6TOBKJNYA@DA?2b6+d&VJ?6/M^RNg5
<Y)3WQ(O[bLOR\/(1ebaXPAWUW^dD9<WXW9KFK>c5UL#/70CJd^S9S__0-)?^>8+
1;g01ZEg<fd]cS2:<8#VK4TR:cX0UXGWMR,?EC6Z3/:C]^bb[Kg=f#-d]50;a]@N
\H[L:N]&ZXE&>60)HR)EQF(DX:-[DXC0g1[Va27E.5ZLW&[]S/13FNg2e^^b9LSP
RAcGaS^b2fM0cPNcUgXURTA8JZaMc(PW1RMT_IZ_.aY1]6C:?V;35/U-8R4^[1K>
J#<@>2;,SE5GTN@8Q?AF^UBC(P)/QV=/LV4L6b;J,;4D,cd9L=VHU7G6C72+f@4+
LPUg7STDQcc:,\E9?(a1Y6U2X\)65-EQ&=N2JN:PP:M(,0_g#><M3f[PG>GMIUMZ
NBaH^CXg03O&1dU&dG_FA8/g8A2,FT_NSFQ3b9<SS=/(__;a]665O()9MQ+DDM)W
E=79AV4=2J7BAI@_d3],F<IHd<<GENC^?a53T?5?_1?I+V+G8c#:38XY5XNI.Sab
F;6EZ==f6.4cK5_2Z+^gD:#&SC6F;f0dPJLMY<)TC/dH=0MR&-ARUK54<+D=<^M&
LaMI8KL5@U5_IfQE()HbQALVTG^=61gFMe^If8d_eC+=O&bg^9IN31c>[>]N)KgQ
/HL]b6Z+0G5J<(=\K4@4e\5?QZX/c^d7e>L_HCKSIZMc).DPc]3T?S,R#M3&\1QT
cCH42/4-Ze/d^&OK]/>f4?0=>6W@[[0;>7TW2D/FO)\J9cG:D1-M/XU.CS\DgZaB
0?;^:Pd<<A?K5=[YGZ:G8[BK0g?PANXPV1@3;1QA.c(NZb\M2YO1(F0BE^(c0P&X
1S9Q/M[bD]WC>R;fg<LCN86]-@S@1FR[B/Ja&-@e;)R-4^(XEPe#V\6]aAR?]M?3
&S>B](c^2:9dLD^L70gAcc;7B1TYDP&DH][24YNG85WR1H=PS7&-<V.RMQF3[QUP
4Y)e(GD9O8&AZ925=2<2(U3.d?0B35^IQ#LD69H+JKCgPfF9JEe[5B]dI:=G8S<4
ADeHX?RWKS/?,C#b7:W<1[DN4J)QD3,[I:3GC+f)+#:I-4@f1Z1HU^d3HgZD]V9c
))K=g;P/M9-PEM[_g>T?K6MdJ#I:6J3VYUY6U-IER^]1P<0NRgOeB]8V)87-7<X]
EH?X/(_^A(W-UKEXRd,(U=3+9OTJJG<#61Kf4+-@f,85G^]Z\:bU:#;\6)3N?S_g
>a?9gYB/\=bWdCX)e]3Kc3:We#c3@;F0TYb2B0CUD1.\QD#O,>])bbJ:8</3aGNM
b/@.8F/2f])g[18Ha?bKf]be&&P#1-3B7@Q>bd\9(-S?7Z_Y?OS5,c-E)5STZALQ
5HWe]Q[;P]UB<H[?T[4TYa[PXIU.#f42_2cQb(AL[de+/T0@;[><FYKe@H6I2]UD
IXKC]#0/MagVeSW8O/8N.:[(KN9:cP23:PKf;3RN/II],W/-9IefWWVW?:BQWSH=
)663OZOQ@SU&(9K>E,L0^E0\&+f,)+4WIZU98B?O=GeLaBA22fVRWJGP6DM4^e7D
HMP-aeM^YH+_#aU++g,>OY5U4#K0[_[#aSFAdBJV.b8=@>?1_^&eM(7-cVB_S(ZJ
d;,:2(C.OOZ@-XA_Y7gDYdbER,b@6e,e03EEB?B66(&g6eS4-X/S([]OOQ)5ET(>
RB1Dce#W2d+/RaNe+aK6+Z7cIFV.I->\;VaN\\?Z/&=H+3R&72NP8)(37C_GZ3@T
Yb&ME[[3dN@F[_95Q]ZBDeAQVaCX_5>?.R,B4K-eAPFaR.)d?FGOccJT58_K]gK;
92+^3,Z=R]b;)5dYID?M8(O3N4eP8B=+#XTIU:[UI\+=@W9<))3_R<)K(eT_O(X7
,B2+@HZGI@1;[Sa@\\2cD&&.H#J.<ce30SY.6Q\CP057,A(fY:@;7RSV?B](9^#J
Q#:6b=6E/bF9AI]JDIS5L082^A-@@H+53WafO:.X);B)gY&(J,FPP9R6VUSSW9.[
RY1G4;NA5XO?43RR6\L?F@UH96L51H8>E<C4.[c?/JL+fJ]8=++&+MT3c)S>,,7E
@G+d);-\.e43<(0XDa/9TN7ZQ-KR9MH<U8egLf,^XN,SA@PX[6eV[#Z=G(0JTP3@
VCf9M=,-Y<fE;J(@PF)]1N9c84a[AdC9cA=aZ9VfS?D^Ld\\c0>dQEa&]7TTfa)V
T80FR\#5T3;[^Z8YL7WU2]\>HGJP\^LMKY??M\GZKeg4b_e)a(X1=5]K>]SFGEOL
>&NBW.a#3;f=&\I3MA.17@a?Jf2c<e58P_;VE16E3bDdS6I#75&[C4G>d65,c]3f
XB@;3/(;N:L(#&PR)Gg_3fE,V[4MK)5(:WA8bG-Q/TYSebH)QVM/141@745<<gK&
K7CE,e8UZ_E(T=]SbUFGe0Q7e7YX<N3VT_S9NP=@,;=eRccY=IFR]^GF^T0;1)T@
7<E@R=_APa&XOUDO<P-=KU[.^(+OPcOSW?0:K(Z:5fg(P:#a,P-XPbUXeX]DTD4:
I<A]^J\PJEOBN.]M?f]0I#5b8F&(XU?NEDdY+Cce-5QMde\QJXN2D1Lgb@?CUcg=
RKWABCP3<,E<W=LCWHCGDW9.ALGLL@VY/HB=]3;&?6?8G4:3YBM<CGVW(+AHNbW)
E1FK+?;d>O@HNNE>>EJ9W&FYg2Y::[1IPP4;b<eEU\0R\=/a<E-FSYb#JQ7(TcL2
YAMD1SX7a,b=E0N@_Ygc&VF2^\NDCS@A5c]59)=)AV]356:FQFTB79XELb&KQZK0
-1KG;3Z6[EAeH(f8JC^XP6Y3<_1]B(XIdNO/N.._LOP[cD97MdKBUb@R?JLcTcFU
5dab[^(OM/A(5GR>b>X-E75UZ]=^9M>9,K[KUC#++(<J=Z\6Qg,_f:g+954EPV#1
]K&6XSO:CU+I:/.Q+\7d,K7bGW>S7ILF0CA8#T4b;F^QH30@J>C:,-CGBFREH#40
fc\-]/5DZHB<.#_S>.S+Xg\;G+2-8OYPR.Q>V>&[ZO#V/+GO/UF>SX,&bRR3f+Q>
@04LNO_H<+>a+2\4f(eZY(g\+C\]=B,MX>FBV#Kd;@2;YOc;&E0fIAMI-DMO#[Z/
H_,9M3fNEV5+=8a1,0+PGSd7^O_+X3Z(8/cPB.M8YaU[aZEAR_#L-&_MXSOaPD49
Fb)W(U3gdXU#7XTS0F(.^^=SADScQ3\OY/YG>D62/>V3JA_\aL0G&QZ4Q31KgEN/
+LZgNJY^#SbQeT^..UUJ#c=6)<BU/MAH+OA4O0dQY([\aOe1H+_Ga_)@ba8KY;FT
LcE[5KUc;_X3CJL6fO(/d(^68eM1^;JeHbZd@4:,fFE\gFAB(eM#G\5XV))]AGL5
Q=5&Q79HM:)J4Z+[:NGdZ?.[FC&aHdd0PHd&8b)Ae-U\54:UFL^^6?I_&0dABL4b
2A96(UMb,C8.PI_WY?Zg4.]]MfJgMDAdQDWT(A7#\-BU?5c7aY&f>b;4>T=gffcR
d=270/+.2fNYVKXKX<D0/5S[ZbED<DF0gM3D2TKV1&B?M-8AgeSNPF,<H4/,a3JJ
S_cM,T:&.M>KV.28N;&:&TJO7>&)=)4g870aIU8O@@g+f:I]a^c_9@785UW4;b-H
^8#a_EFeIS0bA5^5O(XA_PK\>4E]FCSV-,)Q[.]aNfTX.WO&1/[X0=BO/ZO0b2G#
KO;BO(=c?M]RCOK_]aPINa9DRG<P^OXX5OM;B@T#:PM+/\faWg=W+ZBERHBGC#X1
OT=bUR)8FJ>YQ0Z3/aeVgGU_b=BQNM5^^GA2W^7??1WSQ[\/DI0>GX/:PVXK;QIU
XAXJOgV/VB\^(]>5:Z(XR[-31\LE)&JSBX6V-B#S=)dYZ(9S1F3^TdGWcf,7IOAd
MFB]LY&A7KP=H]51I0a<(D[H/RD3I>2KOMeS3T6^=KF-aP3QL:b-Qb&:8)#C)F71
gTR1f[gHJIadV=Gcgfa?#-WTW1XW.BFf9(@Jf6W-ZdKcV?+a\=VJ5=NJ9^@Db2]-
^agc^^Fe_W/QJQeXHb+03EN47I#ge?Y6(1g(];1Z3=NGZcV>5_80&4?3c&FbJ@?9
1:_VEM\OAHAbX>/AN,HR=Xf2_Y;79N@[c_FW1Q5Q4Bd-,BXFFP\@dLbBC[\HaADT
ec2]BbdO_PER3>&L>Rb::db,JR:fPII@2,Lf062ID+KTbcZ[V/G#bGdW]e-:#G(;
^J#[65NK?D.\4R=5Y>_#.1^cD?f\XA.4KbTU-5P@0C/6\09AR,ON\[e:WNa=ZbeH
]PM,Td.8>A<8)aAN-Y.^)]WaPTN/NbK@VP=CbcD7.]=#d@Vd_8>3QM8)L>OC?Ld3
MD91^\YfU&QTKAT:Q)9XW]]I.ZW-+Q7,WG-dF,VU[?3/A#_X?+93cg5S[(gW]Q@A
<J^\HA/J68LAFG,TANId22N(]8Xc/7_X-;:EJ<gYWS;O2H#cI-AJC=GC5A(-S(Y1
\f3ZF1gZac/Na=M:(<K))@1LH#=5[E0EI^[BM@93c-<-.3[@LID6-7^K7+\X5MDO
V(T/IDLEI6X)8JGY#+1cf)S131Y3@2<Tb>3;c7G2XX]gD(F??6.+]4L?6./4;USX
_SVeL.?UJZN1Ab>5Cb)NOCd7:9Z68T#/--.,^D0L2,QNX,BPWQ?e_G,_GV/d>#^<
_SS&I2Pa&4KSLZ9De.2WII+=P(fLH=Q>T.83&+,/d)g&Q;N^[Y0[ICNR&T-3:dXN
A7EK7EO?W;EdS5#c:11+UFEd?U90XH==92M(CCQ?N.ZHQZJ?TEMWI&^?=2XH83]/
UGbD2M?BS10OL>bB:F.UR14)I^^)g5;g[RY#Bc0;;;3974:?dXaXN<P/3<?11@F9
\)OI7-O[=TJe:X]>4^=c[CBW-A8()7_M/HgU0DASYFYH#-_C+.WAKeP@08:cF0dH
NEC2SU9^.Y^>?E?__<X.>H5.]L-.:SK3&>,6P09FIT9#2GBYPDbb&I>2=COMXTa\
fcK4X9H1^J^C<3W=)/Fb/gW8<1R=1;D]Cb:<eFPT@8S^GKb-#95CI+bP6Mc^;AT,
4QPHI)#J4@.PJ:KgG2A#a27;&ICBg9U#f_C\R[(SIUH6#/-X>+fcXcXI=QQ+PH(H
FgcN.8BCST]@KN_K-OZ/U_.?L_Y6Ce0@1dH?<4^bPZ\9UcLK8J2SJ3-@L^&FYVd.
:V59Y.A#U_=,>.ZR&+0P-0eHENG_Q48L#1Vf@D61]:42g-Y>5ga9D&?#c_Y#MC,0
Yc33@dY7W(+B=a/D=c:LBgG?Z:W969]C^ISb_?][=G[:a;@]D.6[J;eeJFZDf57I
G?N,1g\DP+_gH\I=-dXEBU#H(eJORKQ(#F0L&>eXW&B(/AS.UFWK2&d1+T^8<J0>
X:X:#(N,SHP3ecN;VM9&ef+C(>d=R.\CXS0-6H&G,=N[/TDY_Z@XFQ9P?35;Q[@:
(d.;D9/+32[Z]CVP]_^_</8B;WgE@4G1K#=]@LD?89D)UW9+FO1EM:.O5=Zad4T1
3fFZ5L&,>0_[eKg2[^=/BUe4(5GgJbTKFRX4>\<F\OV<_Rga+)ZY]56K7e&D,)]+
f(.NJ3&9Y#<SJN=^E0UITM5fC(g4^JJ@F_,b.1AK,8(_,<1U83E9:V2dZ5N;1A5d
_4M@QS<DI>IGZeU,B3?XR<cIgdNLe)Q_aV&#/aNJ,/7e<RAS(K[T4gc/bdHe4QQS
#O63^WN6\eDFTXgUES^)9Z]TSK[c6+5QOJWg+H^_G(0J0,4UK6/:&S_gcJ)CPf=O
54b(\#9/VN:@bZX9,dT5=2JP-V0Z^\054X0024E30#&/6XUZ>_4Y?I6N?@c)8Q_4
4,(P&f>a91E6f\gP5f470Y?/]:BfK=F+A8AgA12J+URCNT:W1;+IF]JQH;cZ,I>?
&F,YBV^P_?S]d_S/85VdCQZY;]+D34T=[MC53aM4_9/-a;)YK</L6;/FEV=gNcPb
.9^bZQ)8McHX;M,-F_,4VAP42<ZX=<8H>?54d&<0X^8[d/PZJcgL_YfV+NOGPY7H
,BL?L];YdTUB(93?T>a)MQ8]P#TL(L#?7\W<;S&_[I,ad84#ZW<0c?HCQGZ3KLg7
_EQb5fE[Y:.W>KbB;F@RBOf+dYVcdc.<\:d5J&5,JJMJP>S65)/^b)#@AGa4ccgU
eIT]eJ.73?cO=_&8XRT-F88J9]&d=Cga6a+ce8DO6?:AYd>XF>I;N9ZDL1-]e19/
4]CDGI)b:M4a.LS,_f(G1W#Y5ZZ?d@2T.DcLVOa@8M;D(ZR.EgJU:1FfPLA?MM1b
1c/:Q4N5#LPRGS#5KXR^>W6fWD)-f/:@7O./gK_PG&,I#:46F5&VgOVOU/?)P3EJ
?+EZ>c.V,XWI0X/VV<RYJJSb@1JKT^G+SdHfPS^3XP849\S;Zb5LW]M+F58T#B9Z
eaBR@59UO^G9@JQbQ>@g<C>N09.b#f>d#PG4[W,c.e#d0#23fODR84/Z8ZR572aW
?_E>,R1a]NaGU)9B]6#>ULE-_<_?FO4U_3<VKJ1f5Ec\cSW7]a^6V6@>B8Pa7g@Q
P7;FT5;MQ<#VOP>bY)G2(VKfH,Z@Q3a,RO+Y_N8f^+M^c?7^;:a4Q4W=^;Ne)#V_
JQcVVIO[3cQ3MUfCbcFa8B=0da13^[2IAP]33H6&U7T8I4:Vf=<>:NTH,\>4)Ug>
7e\>Z(EID/d9N4@#2a3ZI\Sd+b83P:6,3Q]#/d4)BUQa&MI4@KMM4PHJS.5T=:>N
>73Y-S6bP=HVE1/4^_M\]>);3TL&7eU;N[/&DdNUWR6fU^-8(NGND.KV^A4.>b8\
8YHQ4DF#V4>GE36ZRbRY/Beg(CF9@FdZde,(C8G5O;Z:BGHM88X3Z(1C,,QLK24U
B4?;FdLOd]D_C&HP?RI/;DdD1CCU(X5KN[^[OYBb^QHOL7NE8IUD#ef&F9a:Z5LZ
c;MI[Cd&MW>5XX3dOFQ=/fZW]@?34d6;H&P69+^.Hb?@?0L?gX;5AHd1.VO#]V9\
H;\.A<>)KS+eL\B9:8[C5K<D02C\JJe:9e6M[-)6NSe=8KZ6G=O[eKf3)Uf6_b8O
?5;T4-S3.B._ELDVd5^.a6/.W^TS]4WIFT+cJ1CSFGCV2a2fE8Y=W>B4a(\7Z#KZ
4W&2@)]D8C\?KO-8(+]58[MO[REc9C3.bYHb1#<8d+T/S#,;3=JG23W95FDa]G]F
1BOQADT\#7Sgega9U;#/;.Bg-/&V=8NQ/WQO;-Z]YaWG4aFaQ)]&&gS:\-48PA2J
eL0BH=,K&7XBEOH=Z#R3Y4+#If\c#a=?<G2?O26OPF4.)W_]+2TRHC:1F;]V<G3J
cP.eC(W@/S.O-S_K6F<ePD64TF_e?9d1OQba6PTcda[P+c@6F90WCPY4R\bZTI[W
>-7Q+<9=SX+R.X+=0cZ79?]+Ja/2dJ,OC,KI:U@Db]^D7=5d3b).;OOZK.J4>8Mb
-7_-MS35:0.RDUURBMGUJGX6G:_=JN_YVfL_Dbd4=e6Zb&d<30d.L(6O#5F9;&L0
LJ0]@d49XGg?O9b;ZdG:??faE=g-6c4TgO8PSZe^I13dE1#&JMb@_6b[0TNb)AO_
D]\\^EdSR46]LdMUeAcdVI4A??N2-S?DNCEfWP:)]9@>-+AJD1Y5f;@fFZZ29Z).
a)1Z5(4V2>,P35)^[I@fI=eY#D:QCE=.)@_XSC#f^aX)\XKSNS9>d03Y\-?ScIH7
ZWfb#4f0g4gC8057NXRUgQ9O+-b\/SNRB^9(R2bR.#c5Ab;;#_8/7a)_?Z)2EY83
O_1M<Fd@WW\C)K[O7d[+a>L;FR?,ZMR<-)Y?<+f5?<JKK&#GW8+-(9)<#J5/>bQ.
,DDG_C->TH##=\^g>5L>_4J74G;c/VFCb@0+cUdSc<d2BMO^+UHe^8a.a79T.X-S
ZeLNd>FHgC1aB2b#Je,8Z)NW:bAEOV]C-:3d#D(d2Ne/#7K//edM]Ag6ebgL9_5N
HNA^L>:Db\^8-)^JA#6TcNG9]HQF,-:gCDV]H]/Ub2QO_@]K10CQ<IU96?])QSO6
N(E[cLX.aKGD6(R2)&,6[1?<V4B&=)=_)aHd]]L.E^?:BVB[f3V]g-TIVY+aF&=X
G>QTC>]YTQ>a)1,6,O740&(.T-I,,Q;@gR@_P(Pa;T4>;E6cdRCIIT^K5Q-2XL5G
J5#H.J652<>7V?gF?T@g]Q,WM>_;F1X9Qb<[NH++,+YW,TQXC#^05,[F65f]AfRR
O6BfSaV=1.eV4LcKIG4^gJWb)O.8HUB_3;f8-GXaf7N:.aaJF^@<a/Kc/X3]W?b^
/c.,)E=V7Sf@[_\J257YaQ]VD<?8J)K?Jf++]FE1[9bTc0\.0?IDO,O0.TKDO<FK
J@)T^^)/1\e5ZLV5c4YT>,:4EML4Y<a(Y79+a@R6b#/CM#MWa[1FV^C64R<ADO7a
(Da7=.H@=Y[L@@/FF1A&4V5T+\9V07ZP)=9J/R)3V5L+EXVFKKa.)de/=5W,U[+c
K9UQ71S)CU@0G]CRS-/X?Y24C\;&X./gg9d+A2gX_Z([H_TG7B?a.\HHA9DA.N)D
V^5=#DK;-<OD<L3Z\+9=<3Ga0MI7.B#Z??N6^d5LU(RWL<1c@4;])DLbcMM_+cPU
T91(_@+fJ\L-?51/OM.V:a:>KNf(gAR-aGAY0fO;U+O+.HBfXa7-IH:]F;_EZe8f
1?(5T)^a=OB9C64\bSI7S:aTeYN1:0L6S]T>Y/?]D=C422&7[3eTD?V3(_,g&LYS
V,&#8CVGR.B-NUDHT@9f^X\)UYBe+?O9#0CKM?F^GQBTSB(&VCCe2H0T1fY9Lc;a
WLUN0P#[-dB?=)\&BdPYG7FQDeWH]J6ZU^af-C8<91aF#@CRZC_KR22ZZ-;:6c2N
a;<61,cEFL?_V6aZe+]7F4#SOIU3M7>GQ:_Z):3[?(O//09^R7LGSXd/^^I^^aPR
_43U6ZGU^>39e<5DOd@<+I^>,^8Qbf^#X(0ZBaO[XF\:6SAC/@^WV@@X+-d8FWZ:
aPWK[VR,?TS^?d[<-:dfEfgee:8#Ia/2BcS99KB:I+?M(Fa,NDbSg[LG-G]5\\<g
_M?9DC(:=@L6ZN;EeMGSC3f.C-=.7Gg\O+#R)RMc92P1<=.US\5TSBXXPS2@HN1D
C.^)L&TJ(LO?ZDc<JGOG;b.5?dZ@DZ92?U=Yad(#&dX.Q4?;G,Ka.2+3U7[0,I>&
E-A;0<W>:]Q30BaIC=c;K_VCZ_<=.DUV[:dA&?<C9Tb1^cBYd#;V]Z3^KeE[Efag
Wd#RXNTW<+:AcCSMERT_fW#a7H)-gV4a/.3D6E:I-KB<-<2+_]\_(1^b^Lg(L]4/
JXaT;S[G#(Y)FBWG@d^-8:<BBL3BNF0_5ZLTL+b622NPg._AAC\@Nb#_13AYB107
3W@aMc-XO&71gA-4889B-;Y<OF4&+WfNP&9HJdA^;_9dX+T3>;PISGg/,FO/<5>D
:KPYDf#^NXZ,&#M+7;/ge0/T6[Qf&#D35/5CaK0g:F+aVG,g-I?S;;,.38EGE.Y1
J7<=/PFV[8RH9f]8<WJI>eSAP^cJI(X?aOK=,DU[ODT]9NFcg5M>M\(GI,6+AKC:
B0^OKGN,&O>B&:8dbSf(ZLZ:E,+cN)Z[NM:_&18+]R#V1(g(\;=\&.5>TN#;K0Mg
#&d_>N=M2N@>gEU7^TbWD1<>#\JAV98Ma\RVM\C7:+O,&1Mea&K4)(6V+<@C=f]<
)dOF1JRcY]bOQYg1db(LR3DcYH?J6J\4eRZGGM9XSa:bL^f1BdAT[Q-6d,/,6Pf7
=W38\EW65KL)I4Qa@2>g--;ZJ#_UYP<e<--].FHJfG/S:C&S:-#b1QFM]?B/BdY4
?B4>G.:A;&=g<0U@AVg9PI&>eMSB3@+gPbWJ-&[O,A>-<,)K]?OAFFED),#JAUPL
f#D(6.eX\C9G7^^Za@B:EcRS_K&&REd-JK@+1cN?AF/FGb6V]+025]Ceb&)#7XN7
b<]aP5OG(U;4ZL9XM(=#cYac0LfCe@?B)QL<06_Bd-2QPdTP\;FH@JZNQ)b+(8N0
-&JH1?+7/:aQ<;6?72Z&;SQ<a1FR&?=0GS/MggXXBV0YbgRf?]5&W0,07c>gK2</
GAgNQdLJXKH;/2[7g7e8JHD.6gAM)57.R5a?GEa=\R\EH^aSQXfRM8L[Q3+8H28?
:B;?BW=;17QV@PWTBIeBANa=(T>9[,6<MRC&U0/:?N4]_cM1=@/Sf9O5Q=XH25ET
(U/e^IQPNFJJ(Z0-9Y:P^FZTN)\b.JVIe6Uf9#]B@7RN^WS8\346Qea/GFKEEg-5
J=-LTM\1a_0CHLBNd.=OOd.W<Qg?,JRXbW9-YZI-;MQG5<>#E2FNL]YOg3BA5b-C
(BVdA^RUXcD.TCQ7Q@2COGDKd&9/1ZeQ)KJ@eMKRLVg?C;M.X46R0HH6=a,#CFdN
BHSEDJdI0GJ/6934.-Z?VWEeY,T&d<NaURZ>K-3G[OLY#079gga(J1KZ&LK-)a+X
Je91QMb>6agXSF9SO\eEH@E7?RH.I#g(D\FJ-OFQAba_9QOHA<>]VHGg]F)?1)=a
F0<\\a^60=Tb?g;<aRWS?<:[C?FNTCYE@=_.cGL1K^JL:F4eaG5bCGTFccFIS&+E
6/M+d0,O)LZS,(.T?^Of,)b>0=P4HUC(dZ3XeYd6RSIEa-U2e/-\Pg-P0_=#0CPa
:T)8gY3K_]J>_2+]TEI&ZXS@JN?WD<a_D826UHd1E9>fD^)#W&:7IG6)Rga9P_6e
dU[QM^Z.Q-NN@+18bT.XGH+J+R;.OU=1P?e]Z4<B.Yc4@?)O7GeL6.\-6:3&GDUK
1+4ZX?d7a)fC<.9W010=R5:W08dL+V<0L1/N\6_[8PG3XG2f\g)A\#=H#+dXR2,?
=Q)8,/I_<#YNHG@91<AX@J81H=f=WT8<PYf-GK2K1G,V3a:.7a_P5]S2MLXD?5GR
]P4RUX6\UD>;].#d5-Pe7@<+M/)K.&J/^IU>O(46<5=YLM>Q7EQHZ6]<N8POBWZc
\L7JWf/0@@B9.S?<C/E9dZM&:c?3Od8)(QN17E51f7HG&GbR,#CG_7ZQ4RAAfL&b
95J2@,E/^K8cTTLEgeY]PH9d\L[CSARF:[@1+O(L06S,R[YHM<d^3[c,;aNBH&00
#WRN.?3V=DA[^/D(V9A[KYa?QZcNW[3O=+OW[A6<T=IM=VYQ_7-Y&)cADWYFGJYM
A>3gSAd6^<V/0Lc17#-LeVPQ+PB[9dR<[.MOc+1c(X4LUW@JGUOD8>N1V2gQ0:Q\
#0a^>D:=8bS>F:9T&5CIaY373=ZW#e_.GX8,Rb/EdcL0BBP-@@aJgC.36KcZ&1S6
M]+5H4<L9ZWL)A2?g-a[DVSFSe0UQFc^A3CGJ-:W/S?>LaC&#H9b[g]9gZQ7J\ea
Z:[Nd-=B)^PZ0a4I55KAQ[)3@3]bXb+U+/O@?-]UBK#;e-];dg\fYZ;FA+0:+=L9
MTQS6C1?+gVH:1D#N@Z^+0ULB(=2T&7W9L#C4+Sb\1>ERZD_<96G#-Bb[P97C/5Z
FEXZZQDGQH/gaf;SGf<7GMAg[/K?;\DFJca]2A]C_,A^_?&DIZQ,80FZe_MJOOc^
9O>LV<D[DC[Zc(WF_/U564@S5H7;QSAd>>S:KKK@VSNC:0EQd>3.^(IdLJ0],3[6
;cCOM]7(b>QEB,J;@HXfTKUPH8W?I:gbD7NX>LA\2CF)=+gM<SE+3,AZ?^@.UA/J
7<R##Y9F;+T[V_+?:.Ld2d^?@KVPDY<4c/8)&Te37OaXa=a<)R][_Q<JC8NfP?OU
?eec\J0eYZLcP8=/f+:0;S]GV^P:XYPQ+VSVX(JM6a[D9/=/gf(AC20(@:YeU>T<
#(=7]8X=3WUK6dI/C4VYEV)3O/2H8PdbW>:]#/,A=M7K^JGF25VG=_fBP\Q-OBP9
.<3IQ?C:XB1gdZ-e72I>O6ZfVJ^,HaPZ>Q30C&Z\)^XYJ?9b,Vb(&KM)OOOUVdIg
>;I[33X4912?I9-(Pe3eO6PIEO9bMEA2_>;0;WOTf.Rf^UD6cP38R;d]6XA[9)Rb
@\FD-1d1^<BY0<,+f9-=^a4-QW,+X;7U@7R8I,#B()M]Y-GX[c6eeUA9JTBV]d+G
G?JaJ_b\]J1A-CPM4D30(UZZcf8W0_5MSdKN(^8E>/e_>]L8ARLXNLc0EO+_Z5;b
S@>?Te#UC_/A@d-)7,XX1B@:AI0+Me/F>KR.O68QGgLUWQ8d]<LL9^OH<a<[(O6W
f+ZR-OI4_#RgXOdXNAA]?@dAgM9=0R_M[E6[VZCOYEc#L6[+P7;4D>X=RaL/R_II
=)Bd;-CI4M>[LXS/]G(N?^?UO5K8YF.DC[d9,?-IEUW853aYSNV/R<62dW55?Q.6
_9g?IENf/@<(e@IB>;BQN?IG4T988P^F<ef(F9_]G00#;^<A_(3\A37>(g.7-9cC
G#XY4P;9:EZNZX6&RVPJ0+]IW,-1IC1Q0bbYF[-+H3TDI/^Vfd\e:T+c@>6dY70Y
-M?8NVdd5_#8VP5V,W;ffF8QBDQ.<]U]F,J7^<XE)-aSM@I-f#)(L9f((e#-G/@4
ALaYe&G/25JBPHN^AZA&C5VbdNY#V(_\]0d?S<SD;0.1K^9a-R=9bD(<bFF;[L--
\Yf]11W)G,OQHUCASI5/]S9[;b<b4+g_5fXb7]/B)4\:)SgO-Qa1_6B8-D0=18Q?
?5F4I9DBV8#7A(^+bCDE>-b/;R\RDC1OTfW<0N<NgACd>@GK:#+gA=fSH3R@S)_D
DdGG2KTWKJNG=,CO\Id-IFMTDE9fM5KES[&H02##P\V,S<46(B2C0aXWeU89;9;U
0:@D))SD[b,TTFeO;WD]P?Fc5Lg,Ec3RJ]K+)T.dTfWLLS#.BB>-FP9-Rc<G(B9E
93^L,RNT&ME15gf+J@4I4+Vbd^B6B]UWVZD<G1<:aB->RKK[bbPXI&d4FD#_W7R<
>6#cWDXQFN1DGM7/;Q/C-+#=RU]M0^MKF#_cCWdY2FeGO+C.7MO\&E\ScN_NBM;Q
QaOMOd^G?dRd7c>HD:(S7OG.8RQHd-f[Qf-J__8AV3;/S9HUL#LAFBVHY-91=/G=
KYTD0,^>0VOP@/=d+S4dU6T]c+Dg+EW(d+C_ZG=/H)+eD&T?PVEXeKZI/7=Rc16H
N-)?b;5KM07aNC(ZB]dHMbF]Y?FU+RbgHaO(fC<a8FgbXa\SHO;U&gOL1A\>N82g
f(gY@=G::&A1<LZH>K^fR^Oe\6^5?^IC[R^:]N-U;71\eN_:-Se;MC]f;I4(^_L^
(3HZfZ0IMI;eK)RQ<9@F,=:WI33@Ac-FO7eJ:Y<7RZUdIDDBg0:8_+E5@XC90>9f
JMRBCCN1O=WW-3&;KeFeG^6H(F:b6TeAO9.5g<2Z+)_b=e5fJ1VK/f-;K62LX#+F
3.(QHeM.7VVOe?b+?<QZ(\6@DRPb[c6H<$
`endprotected


`ifdef SVT_VMM_TECHNOLOGY
/** @endcond*/
`endif
  
`endif
