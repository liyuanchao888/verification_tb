
`ifndef GUARD_SVT_AHB_MASTER_UVM_SV
`define GUARD_SVT_AHB_MASTER_UVM_SV

typedef class svt_ahb_master_callback;

`ifdef SVT_UVM_TECHNOLOGY
typedef uvm_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`else
typedef svt_callbacks#(svt_ahb_master,svt_ahb_master_callback) svt_ahb_master_callback_pool;
`endif

// =============================================================================
/** This class is UVM Driver that implements an AHB MASTER component. */
class svt_ahb_master extends svt_driver#(svt_ahb_master_transaction);

`ifdef SVT_UVM_TECHNOLOGY
  `uvm_register_cb(svt_ahb_master, svt_ahb_master_callback)
`endif

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  //vcs_lic_vip_protect
    `protected
)6SCg]OT5/K&(&F&>SfDVJ14gJ+eYeDY)JZB0J(L@ZPEHHWXQ,ZM/(M=]97;\TYE
FLg,>[6Z7F0Z,-QVQgV9#@#b_0cdfED/f/MB1SOT(L.V1LGC.D:9BK8]dT#(OM&R
fCD,0U\@9+1:\@5cf3@JLd^)9daW+Q?B0[:P@M6<MR&6LGET4,Og79g<S&(-aCK1
P(^bMW7TcHJf_E&TP\2O7IV.6Y?d@Hg1fA8@34DVWIf#g3SfP_ER?BB096fMNc=N
GM4W(96f86A1&9,<^<beE?_Z(cE@KP@LW3P9IU5Y0>@_#b[&+@:N/e_Cb&#K@2P]
(L245FKOM7EUT([0M>G.C8J&c]#KB\ZY[X]M?f,SG?eX-73<;\QVCO-BdaGS[B5(
#BUMDUN6ROb=VIR-)VW#W8RA7F<cI/?M0O(/=AZXZNJ,70a?e__DXSFJV2aF@A)0
Z#_:?VZ<0.3FB,T7VBMPTE;J>PLZC[a3>cfEOZJZH4\=Q?BY>/Rb9)5?XWT&d#>-
<A?K]Y>BHFZ;5I-&UEcMOHJJE,6=^-+0-UPOa0R4f/0X=J)SBWI,(82[bP+.^U;(
U0\RA(HR;SL8f]0+Fa(^,(QLbdD1RU6f74.;;4Q>,=H:-L4].X[0gVH8:3gM/O?Q
aS4T/cTOX3GG(TLXdY9LM=[:@KH#=Y-CY._e>DQ2WP4?(KH4[0B57QH8M$
`endprotected

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  
  /** @cond PRIVATE */
  /** Common features of MASTER components */
  protected svt_ahb_master_active_common common;

  /** Configuration object copy to be used in set/get operations. */
  protected svt_ahb_master_configuration cfg_snapshot;
  
  /** @endcond */

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg;

  /** Transaction counter */
  local int xact_count = 0;

  /** Indicates if item_done is invoked. */
  local bit is_item_done = 0;

  /** Indicates if drive_xact is complete. */
  local bit is_drive_xact_complete = 0;
  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE)
  `svt_xvm_component_utils_end


  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * CONSTRUCTOR: Create a new driver instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the common class
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual function void build();
`endif

  // ---------------------------------------------------------------------------
`ifdef SVT_UVM_TECHNOLOGY
  /**
   * End of Elaboration Phase
   * Disables automatic item recording if the feature is available
   */
  extern virtual function void end_of_elaboration_phase (uvm_phase phase);
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Run phase
   * Starts persistent threads like consume_from_seq_item_port()
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif


  
/** @cond PRIVATE */
  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  //----------------------------------------------------------------------------
  /** PRIVATE METHODS */
  // ---------------------------------------------------------------------------
  /** Method which manages seq_item_port */
  extern protected task consume_from_seq_item_port();
  
  /** Method which fetches next transaction from sequencer and preprocess the same. */
  // This method drop the transaction if it crosses the slave address boundary.
  extern virtual task fetch_and_preprocess_xact(output svt_ahb_master_transaction xact, ref bit drop, output bit drop_xact);

  /** Method that is responsible to invoke the master_active_common methods to drive the transaction. */
  extern virtual task drive_transaction(svt_ahb_master_transaction xact, bit invoke_start_transaction);

  /** Method that waits for an event to prefetch next request and then prefetch the next request. */
  extern virtual task wait_to_fetch_next_req(output svt_ahb_master_transaction next_req, ref bit drop_next_req);
  
  // ---------------------------------------------------------------------------
  /** Method to set common */
  extern function void set_common(svt_ahb_master_active_common common);


  //----------------------------------------------------------------------------
  /** OOP CALLBACK METHODS Implemented in this class. */
  //----------------------------------------------------------------------------

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual protected function void post_input_port_get(svt_ahb_master_transaction xact, ref bit drop);

  //----------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   *
   * @param xact A reference to the transaction descriptor object of interest.
   */
  extern virtual protected function void input_port_cov(svt_ahb_master_transaction xact);

  // ---------------------------------------------------------------------------
  /** 
   * Called after getting a transaction from the input tlm port.
   * 
   * This method issues the <i>post_input_port_get</i> callback using the
   * callback macro.
   * 
   * Overriding implementations in extended classes must ensure that the callbacks
   * get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   * 
   * @param drop A bit that is set if this transaction is to be dropped.
   */
  extern virtual task post_input_port_get_cb_exec(svt_ahb_master_transaction xact, ref bit drop);

  // ---------------------------------------------------------------------------
  /**
   * Callback issued to allow the testbench to collect functional coverage
   * information from a transaction received at the input channel which is connected
   * to the generator.
   * 
   * This method issues the <i>input_port_cov</i> callback using the
   * `uvm_do_callbacks macro. Overriding implementations in extended classes must
   * ensure that the callbacks get executed correctly.
   *
   * @param xact A reference to the data descriptor object of interest.
   */
  extern virtual task input_port_cov_cb_exec(svt_ahb_master_transaction xact);

/** @endcond */

//vcs_lic_vip_protect
  `protected
G/]+W;\N\69TB(:TbJ+cYS\UGK&82C:\\WL,e)8\FFI>==Q5SCP2,(L@V5.BC0Y6
;+T2UN6Sc:G8P43g^G,M)5OO\F9MUB)_8Q#SdTB83]KU5G]DO&F=IXL-\BX[>S+W
>&F_I@J?WOS1[0IKW4eA7\NcBJ;4=-QDgRVeMf+[@[E8F+2;TX<12F\_f]PW#S05
P^]1476E&B68>=bSO2ST-]LHMJ55\VUe&3E;Oa\5@Pg5H,V)56E6DE1S)50gdRF8
ZG\_;=C]KPe.]YQC7eC^-8LH6$
`endprotected


endclass

`protected
8+(>(QOfDX#//eF?(XcHG^_EP3U&197M0QDSG&LD&9;NU+JOFceX&);?UI&:Y(a2
TRQc610ReD,LXE(DG0W)]gE,;UEMMH,+1#S:<&98baL:@T\>1bg6JHYcR;+WET9?
J&:VF:S#V;ad7-/,aG(+]SP_bGS;\QfG:0_L>bQ&RMREBF?aS>BKRK56=R<KM1+R
CE9OJ81GcIX5c9M<X]-/gIffB/:9H(YC]LfYae@378A>0AVd9AZ9VK47:<5&HB5f
1f?B=OZd003:[C2X?XJfE_X\/b=[-[2F18bDOS2U7&B:dO&=PbBa(>Ta4?=?0(dQ
:EVC6\RKV.E)JN;0T.cXEHX\7$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
6MH=,#/=(D#IRUf,416Ef_VaP=Y8>6cJ9MDML_CEM(XX(V9[?.,&7(-TLF6c.b-P
F,=@22XW1XC&?Ma5I9ff:a;;)3)5ZX55WYZTc5@\c6g,MfRCdKdBNB_(gCKFOYe7
b,ML+)Gce-QH0Sg=DD3L+Je-QK^IQ4?)38JNMN0BG/523GR^-cc3>#NFXQO#J,^K
6XO&6<DZ(7Sb9;3[f@@0CLG>[e+[L>CK#?ODe:Q3S(d]=J0O<W2YNY^)Y/9])K=8
HDB84AW4)+Zd39@cWF)JQ/G<fV<?RO2\X:dJ.CKWG48-LR.;-@IR+63N?_T32<>R
^01#;7BMF?cb15cU#bL>A].N\JQIFDX&S5[9Nd,^=;ROJH0@PQ(<c/3ObG_LS_&4
PFN0?(+7><K>9D5HUY20,L[dTc^G.,+^fSR+c2_F2ISSZe^8G\GDUK[,]3:b92A6
.K?:?EE/CKRe<O<J81L<N6K=U#-9+SBO?Z__?[@:D#+^V>Wa72eSL]dU0/CZOE>-
\)DV).I)A9F(EcECV+Z-V#V#VZ7X=ge^RPg&Ie8@<Vc[7L;dX=aef.f+K.Gfd9OU
[d&(\+D<a7daQS?D&eb4(2SX.gK?K>N@73.>ORL.O1eF5B,#e9PNZ9D18>^QGL=P
5,BZHQ.6A3=Z8P-KY#B)&W+E]RZ9e^gga.ceN[Y8cQ-9PeIA2Ed,5Gda0I@9R<eX
(IES8QVe&:1D_ZB30_d<B;[=<H;7G&D(U-93&f4TZSMVa;UO0R,J<3Vdd/;<Q0eM
T]VdCWXCB9J83^@07M.P2eMS?>63g)@(P\9#Q[^6Q4Q_)+C_WV3b41dS-V0(QA3M
VX?4W4.\O-)C4267Of1]3Pe6?e]5-<e)5+GRdN4(bB+?g=FQ.4SgFT?2f0/O-dK#
766]-V5SI4>Z#cJ8cIYP/QQ0-\QYL1_?J_L4LK,dQ)^SEfW,[/BF5WRZa2?XJXJ>
3_H.dBe4X.Q6(7RO\D2+T2M=E1\+a&S0_WSWbMe\^+D)eO+U6:K/C02RgJ_KFLYW
1R_KL[3f14OJUdC#5UcI?DdAN9GQ9X6;C9F(0M#N.4bE:ES7IaVQ3_gXX+,::([9
0IKL#X1#0/MP#^11W1].eF+^::.)1:6BNTCV-E#5eeQSc#Bd8U8GO<3.R1]7HILT
c./B=@2],@eTa@a^0)S.aF@cNMMZXD-O:1W\-+XR&d?UbB][YJF+IJ.>\N@Gg3.)
S,X54_(7c5=,8<#RAaJ/dZA^_K8JF;X_2UcaPbd@f7;9SUXe\)#]5fQU3\X)=2KK
;=[@1Y5((084g.N_?:<1UCb]bAO6\^c?>KT=FL[A@^53dR,Td)+Lf__(>Ye8ga@@
a</<J(D0?dD+S8gE\P6U<a[#XGBEW,@;\>-W0>7I\L+Ge73DO\CS5C\<2APAO-X(
E-&->DDXgT,^L/Z0[2G]S?P6-cc@0H>V=GI:I7d>M5QJ3\1M+geM>gX.VEHde#DD
W4H:aafMIGFbg,gg@UXeDa#2KF)6W;8XI>;2g10F5bPA7/^YPB34-Pc-8[>c)^9I
6RQAH9;_)N6M+cNJaX_?BESb(a)O#P.KQA0I[#]F7V40;[KC@LPI7Ma>DbO3UKZK
?BKY6@YZ^51BO)\2[Yd?Db(\JHE(I4D=/\D6:X)[T\I)S4=Y&V93<TJ#S,TP:M4Y
X9FM49J/7c\MHBFUd-FUDYKL4V>H\>)JgQLXZ+KJJZUD0UMgd6BVB5E.1U#VJ4@A
/&NgO8)[#/?O?-7d989K9S5G02Uc#WQ3AUa1H;K6LB7B\A-bLDVO1DW6KWQ;g@^/
:f1a;C1/\gN_Bc@KX)fBb6:#V,^(H_9=I65;WE_FAg1=#=5+NbH@2Dg<?F_RZDS9
e_]gHD97Y+c0@1QV&X>5R;1cM9,+SMFT(799(c?-1>F7_c398Ff4?WDY=3aWbe>G
@L0D>,1_L@)XCFW0#;c_25YF&C9#K>E1>eTM/0_2>TBYC:Oe1?#;C/g8J57KgP;Z
\4G&EH272KKY>P0LW/>P0049f#gcU\8[J)/b-:RL-[YXD_2cK4Tgbc&c5a:ff9C<
MCU7eb)E_71:C,6PILK71E3_a++VF[@?YN-QMO:#/Z.RL,\)80G2C8RA<Y8KV_KK
_+g(REP?Ed6g_DfJ@+]RD<4fJLf.[R;0Q>P]N9fb0HG(.&dB1?CI;W0CO^=#\bKg
1e.7N?[d.e#2JNIS;6G)W/S>5;Q86a&<,<G@C\J)FCDWc<R?Df@CYU,@FYQKH8HW
dE42/&07gbQ3E?[I]A76J4KMSV<_Q.O/(7&=7AH-&D.(7REP:0;)477]=PKDb+K[
Lg,K.7TJdUcWE3EWRL(-.E5D7J8JJDI;KETg:WZ102YPWT4C?N-61b^?\1gG#8cQ
=Q2+Q3=b??K+:dU+NZH]+5b,I+3c3:fU)e9EONY<YW\K-fJVT&+OZF3aDHD;UO&\
CZf6X-_AIQ82QHP6-]57d&.;3fB:(bNC9:N/](\?6U]\Y;5DdLV@(;U3=X0<bI2\
@?bOe_5L]S_-3I&421&f?GT]\F7RG2aXH^/H]:4Q83XT_[Z6PYg0YWY:^)2NHAfF
V7>fG#,))=agY-9KQSK\TaJ&^.+Dc88LDcJAa0:JZbGM/7e?g>a\<@MF)Gb8gg>,
M#G^TQ=Lceee1-&SR:1]G]G4:^[f)O.K(ffZ9)]Dd,PcSa/Fd?K=_+7;1/YN0DL4
^[?QeDDWfH+bQYO3T)_#U,bCO3U3R6):#:4PA@50g-:I1T[Ie]\\@fNfLN=4bU5P
RVQES/A8-bEU:T/1F1G4S0aN91@d.;B2;DR4Td5?S,1]fGT@A;:&IgJN663F9+[6
_984>>[[?@SSZKI[EDPCVD]Ha1f<-BXM7.ZYKJ[OJ#H#Q,N;S&;MF^Xeb&7.+6b<
9=8gM32.19HLVL^4EEBP&;\0T)gaZ?N&Hb266YS8S.(>XX>HcDYQ/H>,(aPQ_:P7
P[Rb6df7aC=GfM]RfKI\Td=GcYNZ4P1&H)N5N91daY3OPc3QF4:e13RDS7/6>Ta;
>C1BP>ABNeQRBKegI+,T^SDP><&TVBMb?5R1c>\0L^7MY0[I\1):7g>P1X6NSX>S
&1UP-B:KgABFM_bS,/Mgd?/^B,GdAFQ>(Cd@f8DM,7LaX5+DA9\>GZ>#caI+LKC?
8\9g#=N6e_[VNTT46-9M1aYTI]FAZa=Fg5L;,LG6@/GG]Y?-P=?B?^.QX:ENGVI;
>M+LFgR+]3H/Ne3HY2CP3P_KQ.ORZ_SIb7LVT[WX?Z8LJNBWUK[MO:2I^fZX:He1
DeY4/TWG?L9Z:]Y0F+F?bfG/1F..[B&G[e=Z/K>e];75+8\_<Xe]D^K=N@0]?Kb)
DdO#<558/OF>\&/NYFSZ/)_NA[\C<OZbJ0@Z@++e1eCZP(0X^AN2\J9-]DW;b_?&
5PI=/?7H>d7PS\T8-5ZIgPT-\d_DW-I(#-VT<+1QFgg&@6Xa<WW/5T#6P9-(+9gS
2+=83V707aITE7@2d)N()0G9F1RNa8N)APZ&E2W>_QN_Z(R05/BDK/X&^>H/BK1W
X_/(;RQ&ac5@D&9<O@KXQEGKWEd.93.EK1.>T=&)c8>8]A=G+OSS#P[=J];90-)2
&fOC^.C\<7-7T/L^,EKaD,Ia+REgY+3/;HX;[+]J;3FIFT21B4Sd60=K#T;H_g,)
.8_1<[>B94^C?Q#a^GN></.IY9(FAaT-Fg,H[@_;TA@QeEVddES@0YK6Z8NJc3dI
><&VdF#](_EI&CBfQ+AI,JRQ?LaI&1Re\b(4-ggg_DQM2?(Yd:FH/7[Q3,ZB77VT
PQ;8+)LA66edXA@c^:7CSWaAc)\,:,g2DQ6=K_/X=HYJaR8XBcQ^J;:I6P8^5-FH
OM.g>^Q.7e>NV-4eQ:=L3V_](:Q>?@<g)QLb<S6((E@MeHXXYUYU(]AI=cAQ9QN>
&E46aUCOeC6-:W_/Z1HZ#0=[>a,P-BbaEa@,PG;bA)WIS7D)/cD1F>IKV3QJ]31#
:^-_FC8-)-4Qg>aW;@WGGGUf5&-8KV(,@g@F;Z0d6Q1g=e0>_1JJR7<,^Pf8S4Gf
a.6E9?73LOKNHfBc+J,bJ5[6+SK\gIZe85>E..QNeP:_I)OX<,\44]+X-KRA1@8_
?1J(f00</KZ=FWHZe7LIVI[9+G378_>TZc#UKG>IXAVMCT2=2K4[0.QQVS(5#\LJ
G(dWfS&a>eaO<CN<,T)_GT:#9>cL+S&dD2#4:M:(BKE]SEe=GQO/5H_@[,W3969Z
XU?,U_?>5DG9=KN37DT.\I5LZ;dMdM,H-d5J.QNCcG<eZ^./NJ1)cW^1_U#W;)[+
F4(8CB_J/<_S=IaNF+-+2<X9\;W73P+7.(LWc/4I<M#X1J/...R:H:U\;=@(YQ2d
U^O#=NH<,c[LNUC#(dEcX>SPNL.&eV7G0c>4LS9XAQ[9BE+M0=2]S=C/bJGQg(;f
MZe20+P0d:.O;E<_(3Y93P,X..d[UW1U&H-FH&J(+4G].ZWV0#E3\Ea1WgO-BKM6
3eVUH.H2\(G9L_X2][:LcF6&8d_g1Q-?2M=W\CZ>.N5YCd74WHPS\;UfSMgY4P[[
6_XPZ6/)gC],),N<6;<#.7&EGN&O,_bN3Vc\dD)]&f>gU?5I]7[T1M.1fg\6eOS.
QA8+BePBU6.(9=GD04&gPdDB+N>6TGa>Ve1+<+,0W.QUW-2O]M,fT(\J&Y_[g+?J
KCdV]-_HN5>+,:+:42UY,GKGJ)aQ8RR5;R=D(.,U;Od>,e@NXS14_U>#_^EGB]D5
EQ<X/0JDb@[?KI:1UF<4Q]D_3Z+Y,FbPX)FTc1^P6d&R]NA:SFN->5_)7M46-7[-
JHFa<;,W^UM9^K05:W75Je5>A]8JVLV(1O7??=;W\a]<^d^-+PG0/5dNZ2>Y/P\4
(F<P7ZY@#(]2+>a],)=A>bE?9B5K:8Qg;N5_^H(f>=FOAa]+@NV&ARb+_eS_@f@g
C?RV_#0.0<@DY,8dEVOTgU&HN\/_[^AJf+5AUagL>+IJF8f<Y7H<E.4,FSLb1:<&
cV=a^fR^B_BO??B\GK]eMJGgF8\RHX/(.MX7?@7&;cR6d??-D4e@]2^eXbFTNfUF
32ZTbcL+EW/^V-]Rf-XeQBA7#S+>S-CcTAI3;^46S@,68BCdbRF?PLOZTOaPXR)4
dW>^1)M6Lb2F;;5?4J81XS57GXMRgCMA8^@L:I=IYR>-d_9aUBa8Y)fS^2O^GL2d
);d9G@5+U7#T+#f0NUg5R_<QIAfBJ@a+E),/QC-<CQe)(^a=E:#(a0aDOL0V0;A8
U-,NZ@#ZCAe/4a2T3ebQTb^^JF4.[Y08F5V2bTK<#+)[OX1?+[(f9aWD6</Md0S6
TJ_c,#AdH0UP1MC#/UF:BLcG>1?Y;?;,FFB9B#dJ1dMb9f;XX=VX23R@+[OW1b^7
@D8eJ#8S5]5BRU,O_UG4R>7MTgU(SCOFV+D6_-]bKgg.>Ng95#](\9#N=.-L+6J&
INP2/XKI-0JC;;dDQ9Q+Z\-Igd6+CA]L;>W--.8;Ba5/]=X;Y@AC^?,HI?LcUTd.
d=AJMZdKa9W.,VHWWdVdVU5NCNIN2F5##;QV&TF]0>KIPHaC]J,P;Fg_,>I];f]S
],DO(EYK_4Uc9&D:#IWNOW2GU_=@VWP8.e^Z<85MIMSKA<^_I>cWY3aT<NIAK(59
b&-?/cXabJ4UEaOE>)[.D4J.JN;O9H=O225;0X06NBScPWY4]b&#(WgX<8=LU.<Q
]KbZFWPX)SSS-,0BX\UBAJBb.DJaG;PeS\fA7-V]c]YdK3NaD]_gLZS^GKaG7P+Z
(8Z?c(7A5EE4OVc#S[a&J-+UW\3_:YUM81:(PGg4E.8,[8B<+KLU(:PX7-SGK(6M
>4W:N3X036J<6/_PH_X)JUa7#,\DZa5)5ZCbU]K]S5PY@@0X=MZ<U(MKT3S\cO77
-[F=F?17HQ>@EV25TW>7aB4&,#5^EAa_VDC&PJBC</D,Kb5Z<?X5T;DDgKPLb+DH
ERLX,S^3-OYH#BQRVMI&aT#OfG#[a3D<?GW^(9MgWZ,PD6\0=_M&fJ+@^7bC:H;S
A.]bc\bRf0JPD&.KTF&GQ0/5d\,,Q8NP,ZWE^9=_?2eKY#Pb9]_=BMWTN60683DJ
.aUd+G?SKGTGY#.0G_LWM8;(<1;K.+3FZ#D(_4f:9DaZ>Qfc3YUWY7Q57d0KL1OM
]-\IfX0]&A,M3+G;-C6R)<Q]0Bf1fgIII--SG9a4K_#9:706X03[):?g/be<E3CW
#eHW=H]U&C2JfdJZ_K^/HYK]DVgINPXdeL,S\//(B7Xf6@P5O,@9=f,;8V=:;248
N=cX6VIM.BIGMa5BS_-<KFWYU/Z9:Ub?BW?Vb35_0(39J&d45-1&#b\H3<0C6fb\
fAX^7\<Yb<?144B^^<0(L0OX#6_[1<QYP-:,a[I[G]/f+8:f6EFgE(QgZ]/)cZ;D
LgO)=+QS;9T7D:&2(8C9aF7D;OYdO:V_X02@?.MB1U^6_[>d;,2#W5)T:?:1G[Zd
d+MOC+9d60b,I0857N_PB>c8[gTF\:JLVLU>\gLN6@[)E@LT+63/K^G[4E)&O+UP
S(-ABH_gcA[<b1ZcH[8>&0Xe#)P-PFNeQ\AG:QA)GI-Sb6OB+S0aG,<KZ&R&/OFV
db752VW2(([<>L<F&]HdWgQ@0(Y^UNM,\#TfCf<IS8R-::2_ENa,OY/K70/@0BZE
)dICBe&YCBG@(=SF7-_IG^,g\.6LcJ<AW#1N72?]<HL^:=DW0A+^_D#A[J];ceN3
_-(/WN[C;OYE8@[5QJeS+WVMD:+\2J?,^GEGF5W#]>L_,V)659?R2:Hf,;9:\V\^
.)--O(d2J,P,A-HIQ\[_1JD@A]RVQWL6@1/8VaO5Q)P-g0INP0]1H4=\4&;<U?@a
_3Da)Xg7?Vc.U\=K<V>>J^>@3<21KUSR8Eb@)TGHL?G?<-;N&KGMKII-QYI-8K&S
cf,D;Q#A<9&ZA\S@+@a7VEH>T[b7<KE#Fd)O3O_VLMK6)a<H<>Mf_/\VRPTL]RW>
=dG@2[WS[_-P7)XBB5LLR.5WW<=1Q:;O6IDf?CEW])Df=&&G6SBUHeU,:eCR#JIE
Ab#T&YDO_[Sb#2DGEA_DXgG1WU^caeB7S,9>XFMN(c&)^[GL[ZLZc72YKR]NdINg
NBa=<[SL^TV\0(XKcgM5A-e.-?V[,d^&EC\QDcR+(@+aT3N7bgcFf^BP]Y,5.d>U
O3K4Q-EO]LeM2a=C9/>;W4QGZ7a5LG\26M?R5JXJ\HAbKZIE7XGg:Q2KFS/Yg;<:
]9K=#EDZ\K4Da#B_TWJ8OV&^Cb,CU#fF0eXeM,6?K<3f9F+PG2UDXKZT/+BX^EMX
4Hg7+<c-5@ZX,WI29ZJcY/35)<5caQ-NW3#)&1?_2Q\RcW3#OfS6-b]?W7\XM9,]
2E[:?f],F#/(Q@U#^/U:8AD(F)[(4EVa/F-C-&:9YJ-=SSdd:KRN>4U:E0<9UG.e
WDP4WJU3a_?5LGZ/N=Id=bg-BN,1X[19N=fO^e0#YTCdZXW3GWc7ZJALf(]B,D_=
0L/7?EVWb:Z0(cESFaaBXO;9<=_Bfg#1S2FWgH&^aE3gU#(O1Fc=aO-0_15+)>--
X5^\3@VB9Q,FG#8gKV,+:I:FC<(aP(FT8<]WSV]eNaACecY;AEb]7bLfAeR]WG2g
&_>_8^I_0]c:.;A1QU=DP.W?5_TcK^Y^JLfK-f8A[TVZXc^Y=1A@SLI;BE0/W0;.
:>-HN9.R[HJYT2.02:e04P0eg<,W:-dc6dALSJHc4WZ,:bE#c1:3.4L7O8YOW-cR
)g0W7;E#S>b&NWX7P;TG8&K60f;REJ<:\;)c/>W[K1CQF<^^&g+[9#ASg];_PRCD
[R46+72Xg&.a>[837>I3TTF[IeBG(8:M.;WKD<R5W@D:.XK]1b;1DT0)1YPfc83:
I.fO3:g+O)#XVd+0,QB>\e@U)]&bEP@K8a-M9@#IH8]&K:Mg[50ePgaW4M0?U^8J
8;#5B@:@OMVQJ,<98VL,]FFXQ[]b/U7_e+=gP.Mc+RRQ?0@6^IdE-?C5d3FO0NE]
/I-PM1PM&Q]L7^AHL[<K)80OXb\099(M<?(YV?0-:Q=/WI\>ag:RYc_;TC;Y+<YA
(P)d[29>PQ/Z>3^^T([2&AeF/E-0@LN_f^2IDgZ_G)9#=f(;c?<b,OHLTU\bH(+X
BT9M-_[R./GW@9eRC4(//W@-2ON3EY,U@2]#Hfc3_CL/C2.#Lc1[+R-E^[ENKP<B
TQNUa_W6RdQ;X(OO+ZEQE)T1VAFa<PL37/V76L-F(JfcS_;7aEP\&4X:OBF0TT9?
ZK4<O]EZ^[ZJP8908=BLSd<#M[+9:\-X3f^KTN@.@OB1/EKb4H];ISBI1&]f[CfD
M2YG=d-//)N2BfDP;.eT]-c[ED2F:\cW<4\U/R^N/>9=GH:.+e&PC3?aW,]M>]7P
C9e96Y[@YHP?\(<TGa<FCLI_@+SH7>#5\a0OU0@AZ6X/8;;1T:de;g\&K8R8^5g)
ca\?cM0<gc&_(4SPaFcP13:f7?3=+5YM#?S+Ye>809DW340;O9(2S\407aBTcfa8
FW;ES]:2R1L/L=_@/^@cdBHBIR14gJ5[O-e@/-dcGb-RLd\TMPQ?a#O-,f5L)>\[
=@AZF-<-8,MFWQWGLPR3:\.?a?_CKHdTKVROcM7WdTg)E.]3C9L(QS:_[&Oc[@M=
_L,VeUMV48d,=1EYV/BN+RQJ4[c0NNN4=MTEG-?:O:F^,?-JZE,.D0N&KXRc)=>0
RZX[(Q,#)b(f144g8I9d8.]U8\bXL9QUBf4@L6<6d)B73fC3aaQJdCd3BYbS\Jc2
Z?a<+d-Ycf?Ia,#Z&X/fH+?I1fDdM-Y]ELc7?Y79a+B-.;#Mb\B3_SQT?Q<WCQce
?M[B=[GdW8Le-?#HfJDTa0O0P&E?36IZ@V,#R>GSJLX;M4Db-UIf[<A;5Rc(Jg:8
FPNF]6a8c(W##L=+C\A1UVR)4Ybf[8CZWR1GSV-SSfUL(#]^UcfWNeB>-F37_YZV
YQDSA5,eS(P>Q4c1AOD?D<-=Z>6,BZ^4N;DA[GZg(cRNC8Wd1]GS,]B(-ND:-5\+
C(Af::e?=\KJJ&d7bQM?>X?-0V6YBL_AR@C:@Z/]L0#[USe7Bc7R5LP),ILe96,D
WSH@AB/ZO^?0UbgL=]N>>M97+[[&OT-VdN]MMM//DX5BW5/5CBT:/.N]0?C0533H
T(R4+8^IQA_1=TI/XfYcE<>MJffN87ZW9D2/eOALUBOC1^-1OIU=W8?@-T3OJG?F
aOQP,Y<bC?YE8Y7K[][?&IC\2PG509U\<7)>gP]caLH+&df+Q3\@6N[08I&C720e
53fMc[eZgS#?J>a#1Z7(+F]=+aBC6BHad&L_VF[T8D+(XHD,g=8a&U6.OP;Bc^ZU
#Qf_K#R=_&=.H#[W;N[;0cZFC+GbfW5VDVEK#Y>)G[T[&T>XT\4bc>SbQEIP?FED
AJbHRPWbRS:+QBKe(6YJ7UWIH/N#f#>Vb>A/,-DBROT5=+gG7#SUZO+e;RC#K[X7
NDYW8J](;=WJ1-T.,b&3X6PS=[#&0HZ<U9H:Bc+V=@P9FbX^7^VW;,#Lf0ABDLE3
/)f2,2+(_I/DC&S@C@:F;0,BBe1/&+PSeJB._4YE,LY801@9HMT9B&E,CN3E5,;V
f;&Q.ZfC/@(fDL[)-4+:DfTd&H[FNU=?OIXW9G/QZ97&3C.(VE/S79<34?FK,R3g
B2CD;VeUfDY5bQ;=Pe(58@.)\Hd.-B8JB=ReZ)a3Q4>VF,-I_D&W8f/,69;E:F5Y
HBH##^I[ad[X9Vb)E^[HMC,g?W2a&\9[/f:Z(CNZ<[7DOa/^-#+1XJ=cCZBG1cD@
Q26NBP_>B5?9.4YR8MA##FG5;56XI-)@fI[Z7R-g2<^\Ob7M406e5Yf[bAbPRB#6
f-IJ46eR2+D>G+]?,gW.\2R).W,AGY1;RSQU,>PJS9=<T5.1PJ;fZ8G+P4VI,,,@
cL02L^fSOdH43[>\?60Z0f;AI553)&N4gRM-\49T6J,J>#b(G.V\/+b3+CB-29ZZ
OZ@E&1LMcB\W&[D\\I0?J@B02ZNH^=WIcERIH0R;1ZWQP[@X7FV@[9YO#H>_;<Me
.#/RP)fUB/VU?\[?I.YJ=FO,Y:44UUR#3A(-Mg&GNaQF:V\9EF_);6\dU8U7ZPaN
8gUdNFcg\L7,HKMY4=:I;:.D.1+;M<ZKNJCCZ,EA[#PGB=2KE?cT5VOJ;3DcT2A)
_-6JMfK>\?^1N[f[#;Y(D-4;,L@Ba_g5gG3\C4ac#0FG1HO.fH95a7F)R@\<V]M8
64Hag,K_5OdML^([USVH(7JE_>,#;:>3YK<d:Y5-.Q6fMb4O];GN1).F@R[g(1/=
-+40O<7d#@6V6fD:H?_F>6H#HNgWK,7GZI-TgJB].Fg3D\>.Kga>ZSQ+[e-T9<X;
7GDc[G9E^=LfA+6X2.&-U&)0G(?\F1WEgbC,WAX.SUDQ^-7=O#dfE:-^Lc1[U?2K
),Na\4bCdJ8a69O]]GG:aY(g?P^;ML_5J_\(M,BZ(R@FFQT;AU=-B@Q8c2_W,IQ^
,4AVe>FJZJQdWG@/.HcQ;I\?b&DN4C5G:QT@RAGNfGfB@;0B5Q?9gZ/N-8GXbPSR
EAYa-dWH5>@HS(Xa7T]8=<J.5;N)>P62UA[RTcb/8f#E^6TIcM9C\L=>M1E+/VI/
V5^>/\(f.b7TdRR_/QA(RS<QZU4bKf62W:V2#9)b1/:4@,Ib0EX5I4>QGJ,VFH[)
a]BP:T-Ve<:ZY)348R&GI.fY/G-7E)@IgC5(QL)eJ(#)YRGMP>M],5O<6P?Bb<6@
gb9]QKW3)/:SBRYdWd:AGQT;ARGcT<B-6(Sb+HC+:A7/a#C)e\_QNU)WVG<bN=[>
[+d05F<TWVSY+RBC6PUE6@9A>Z]K\+_918/F0C[:3)]DMb&O8(:bdHJXH4-X8]5V
O#B_/1,S]OW?)U:+V8_3>bFVOJ33#>Z[5H=DM:;1F8bK?RN>I#1,f-SgS2acTB:V
SCf08J41YAC3.]S2JR#:<IbE]db?d3/EdN39_?S@GKQ6cRC94CZG:gV>.8e8g#=V
eMSMB7gJ3AFW?&F(FHg?F.)?:=_J0ZR#.)6E7]TVS7Z#-JG;Q+1VFdXOgeAQBdQc
PP(.>>dDG]?MI33(d.;BB;a0.;OSJ7RMXVaX:MBbE,BV1[]1B))IYT#b/VC>_\9N
583C=&B7bY>AFP^>.^=BJ=9DEI=\J6aL)g#F18NZ>917SYJ2;5MCfFN\DTEY6gCS
0-O(9L]7GBUg2g]UN.eRMH@E+]&-4>S4>/#Ea94>6>>]/AF8bYc.9@&JQ-T5D:Q[
.g(>fdPR446/OXADV^8ZG1F=;QgPc,PORF#)c=4T176182/X&[B^I^G[\>A2XAF0
T6&0Vg[1/@>WN_caK.d&VSNLBBVA?(a&S^L#F^K^VLBQ]>EL-V:g]WI5+YP=\4Me
^0O/9eQ,IK2=N6gCGT<dNF4-]d_4J7=@@f)-)@LC#TaY[7g5<J@Be+FM>7=+/E1S
0SC^=5Y;VG4D+53eAI)_5_>Vec]Z0X9AZeAQ8;<G80JCD=HSBPCTI1>(8F:3JI;Z
4Y5UPQO,V<]e=OcO68#_FJ@1EYfV052](?F)G_6M^O?FU3--/3bR,@YZ5LW?WcDf
Kb6aPUM=X/:_[;#<IbA6CL)/J=T6=g8^8BK#?)0=6TWc,ERC&CeEXU4a[#gGO;&O
bE99^eCJ5(g/&EH3-P&;-g[]#(TO8gR@C8NMY]\R\bV#[][4e+X113_AMFcfb)^#
SP?Y]/\fT_/QW4?NP,c,\2H?O8R,OD^WXe[PgFT^G1V=f,;6AX@&V5c(E9:[1QNG
\3^N9N>YNL19)X#&KRXARSL/f62^:agbd5=8(J1(SUP#6VB:3[15IA=gG)(KgCNB
.FgM1WIL.P_]/4I;]a8a9V)E]6^-AGJT-.T.KAJR@P&cG&V<3g]LPb90C7KOHd31
a=G#c?]^&[c^bCS=b;O_]e?Re[HCcMSZQPWdH/CQW&C]c#f<Y@]K2gU,cNV]&OXX
&:_>TEM]Be-6gA)0NRd[/\M^g<@4F+2SV(U&8Y)/eedMXE8c.&QVISUCPYW#QJK)
T,,2VeQf1H,.aa.49/02B2:eT/<5L>HEFd;Jgdg7E4.JM[N[Z]DL>1&5J>[0V2f6
IE=cJbSSI=W&e+_KSG4?F.M:bD(.U1Q\C1A,]Q?H\JA5FS-.OX&O<P6U30;?O#)O
WQ5d,\:[?U^Q^PPB1IL6<D:,CbfGab<?K?JdbNZa&1H?Q<g1Q23/Y/g8-;Y;EM5d
dIO?<^G2A_D83cK)KBPFf,QKGN)H&79?^S;1eNa=[;/6\;V2GC5PA^TAPGT&SC<2
eL1dY@ZR(NSWd1Z0[0].+6Z92X?A#NHNL7ecB:8OF_=6A/:7?#^JXE;52E-?)(>(
S[gBV-,gf1ADe#^Y5RH0WU0<DW#-NTWa/(8,1D@V:SAMS&#>ML:9PI6X(GP4;7Q4
c>JL?YLRB;6:]>b/EHKZTS-.(Ke.&&O56,9_&/Rd=Rg,^X+0VM.E>\8X-9b8>-D:
2;)b=44^K9G@?ZC)K@Z<Q0]-(-NLKPMW<X?AAB_^BUTY:KX.Ia(;J6YYXVO&K8X6
?(gEeK)7_KcV\3Q_7G489JU3G03.bMGPQYWgN-6>cgb]T^dL;;.dYGGOag,A0NLf
+<fA9E;E,G#_T=TELLaP[JH.B3OQ>046J9<,G\.fgJfcI@S]7LbRfF9>9ENVE+I(
X3I\FKg(bb>.g@PIaB^#?5YaSQ^#LG69W,M0E7E)MKGV:\#N0\c5(&2;[&c,We#g
W(Q(aY?8+<b92QWa[&\/JIbAZM;D5:A&W-FKcLU&\MccBRDe)+7X;HJ4=6X.&faR
>G=H8c\>DIV\7)TOG_=ZUa>.Z+T\C,ZeVQL-7Y@U8C7]b\W9#VcR/-[&SbIW8f0f
GeQ=BZ?->(6ZBIQ.0KFMT1,IID,c0c>44[6C\ML8+94@TE85Q^58B=4#.+QJ2aET
L&FeYP,<,O7]5HTSKKU=Q6FW>?9gMRU.._B0@#&X[,R;BC/R<K15G.W10gRQ>9gG
56T(_ggWH^f(<6SM(+44CD;b&)D[>QTR,>C5&Z81>K8@fY7fIb--H(T6P9bA7ME&
;-FF(1.MO;B[1<I-?<NP@_)0d:?4C3dQ=>\7MeC0<NNLEW&Y8S\#gd^K(4:&<>B,
M^>BZUOCg5#UZHU:&R4OR#B?^D&@B\,5B_6W?4G4?/:a;NLA\6>T(7V@c\K+)Y__
S->/DT]=TSB.1_M;&dMYHY8N7C??^-+,@Q2/8ZGJ(E)<]0TgH8QQU<,>LP&L^T>#
gL1f;gM>DOJG(@+fT+)_AZO==AL.KW4M01IG;OH80;7#c0I-N&DZ?5.)B^HD6+(6
Nb7b#<[GDM)[B1Wf,1:DB86e<GgDIVNa5c<@aVAfMM/2aSARG#+<b3;(8;5KF5BX
_3L&@:PO2Q0AeLLM_b/3W)W)A8aBfUa=QW-8\WN]&?Q[Q[GGaSJ:VAE+G\Y<,&3f
T;X5BKYRGcG=WF5FZTf[>^gNAe,D)&Z23Pd\Q@aP#A=IFB>A+0eQ;5deXR:C^Ub(
K-/3^P@MG>++#M7M<_daU3HZGb1>5[K>M&EHD?CWHX\M#HW>:[0<=820]M.K.[SE
P=G[4EaUNS\#DS+L1N5U-[0N&)6?;X8X_3CAGTdWVM]J5WQ@3.U6cY_,<=2=&a=M
D_ULf1Y&RDZDRL=\bE:.PPBg#;88fWUND5HN?LfC/Pc3-#&?HcD,OC\TIX=47c+Z
-VE3@aDB(\VQbG?T3FC,:d4Pb?@2SI\=?8##+YYI5LKL=D&@?eG5?VWb@HR?0YXE
B9J1Y=);WV9N@O@5bG2A=_PLN3dU,,^>(NB(</](RQ;6T;:)W+CQbD7;6\(TWK?I
[6.K_B>[8PT/@3Vb05<8V]MB]D.Y0Z)<QcCG8N8U[0P#10#4&[SaY12>>,JWY7Eb
#R,25)beMX1+WJ2R1M_MEY]dgfP+3VbfP[]Af<]CdTR\5;RbX(eQ,IU.JP#8d\?.
#/Y8DLWf<NN([d+HbK/H1,PI_?/Q=Wb:?,HR?/WB5/f4b5&HJ0HRZZ)(BICF\41C
GF4ORf=J;[3:/D?;P4V:>YC8e:(#D2f@YE91D<b2QC..O_@>gK/B;RSU<^8)S5/e
#THT>J8YQV8X#DP-TWONH(eVZ]?K>_)J+3F^T4:/S\0bLRJ:ZcRF)KIPE4),IN&Q
K)>18<K\G&GZVC@YOI2,,B=DYSg0B2A.?[G/[BC@@9[Jb:TfP+V3P6WYJ?D[YGa^
gbPE?cDTB1Z5).V,HK)C6^#ED;@W\[]AJA-_>M>@WcCDP[>>5Af0<:&)0SJT7gTd
\gdfX)/<>3JW40>@Yg=WH3C6/KEd<2KX#e:-(+:L@Ud=:Hc26CA4VFMFP.0+^#3]
gdKS:L;<;<->,179(F\:7IDRaZ<W,X?c2?&W4Z0ZVTNFEVHFRJK=SN<.H;F-=O^5
b43/:ee3F43LLW.T_[a\()\d=&VWCCD7V8(cbANG4W7288SI5-UQ>(aF(^J]S\5X
4_bQM-e;A54C<O1]DZD0M_W41=[Kb\K1N6+dRAWM-K5H(5-#D9F6(E7X)PKRZ+&\
K_H?6,Q<U,W08.cBU]8f\Q?@KZ3cUg_L=WDBa_a&5\F3Wfd3F\C9GfFF)GWW,QQK
X4FCF8\(;H,BA0=K8#QY)->R)c&&)_H:L+VH0Y-O.5&EF@@BUCeJ1I@G)IDYCa[O
(@TJFEaB<RQ3-;?:Q58)X]\E\8[VaT7eR9<0DZD@7R82;-TfL^@@5e#-3QdgDG,V
>SPdWVZ]BZ[Q1V)Z;[&;AYMHP11^[IDa\Qg:A]KNKTL\YGG\SOB=BJ20S3=U[RMN
4KGF7b-E^XBA>gY6(^HV2J0?L:8]]E\<KY\fTJY,-g/(32]55g8=b.;-#6YKP+O.
<TccTV#A[0#c.e\[6UYfWa5B<L=QaF[I3H@N;R64<Jb(@<2].0:V/--J)5CccC.c
AW\/?R#\<6,9X?R5\PfV5K:&Ve[RZ-YdNd9:94]KKXMU<;\I0_5DFB46]:J-M\ER
M4+J\0UH9T2#1L?BRB#c>QODWgGRXN;++MM)S.Ee.)Nd8<))6;06955e\\aSTD?S
GbXTGf:^8bES&758VN.A>E?)GQ8/g6BZ06eFHX81Z6PMK1?FU5R>Y@VO4ER9BcNP
G&ZdK459e-\DJb7T\.04\5g6/EL\O)SJI<O1V[\cZ^TQd1=;VeE<]J7T_#E&96[0
)]/:e#2L/)?3\<:C,I8(0P2;QARTMV\H1Q:P_T1WITa]U-12?1N^E]]B^=.B,0-b
WMSU\2DD+1OCULX#]EWIBDOJ.&/==??^84?KLbbc7<Pf9U0>GQF7_&fN/Q=:aK7V
F8:g6_\MQ@=8BFfA+PEdZ1J\AaH?TNS]WC2@J75#U6I2d(?](RR?Y[NXPa@(V^[4
U>R@]J:)MF)VE&F@Q<W,e:L#ZP#=M4ICeVB33TH5QgD:G2T29@:S&Y<f4eH\gY:P
1;7PWe65XRXaES,LO1LCB[HQO)<]WWUfME&T[C53gY8NX^8ILYR;6<fM-M0[>8^6
IWNOeRN&e6=9^OHU/&Q;C/356QXOHQN(e;8QBc>bII?H0M6VQV_@LJ)FV[J.1Z^N
eZP:>4HV25;@\:-2Fce_6/Ya@^19f3bNDY2U15>,;#(+e+d-UB1EAOOG_-e\Z=D?
?/4(JE96C;[?633V#MBVIg5eILO.,TbWLUNN@SNB58f5LOY@3@d2,9\EO1]L]b3,
Daf^_?I1Z#IdC@W)c\Ob&KC7YZB-#_M0/Cc]1?e4W6Zc)>:8f.JUa\J)<4S?^EaC
)JHL7gd5d:DR)V.7Lc69[QZKIeTN=0cB1A/4;=)+Q=0OUIISd:_Ubb=fYG6Y94VP
?1551+eSACMDBO,\WR>AH=S^Y@_G#6cZgVWY<QF7A=U4<KT._2A4KPfY49#cKa0]
((]Y7gdI3K,2UCd7\bb9e+5:S22SD7BVaKG&#GP>#Q7\ZF#0:)VN1D/+))VU:,6-
/Z(:SBM(-<BI:3+YdUaC1TUbRSIKPVCO<+8&5a,#B,M0(@LS^9X(=7.T0UB3^Q7E
5<@f1/G:?c[ad>=b&+0Y>S<dbgJO9AgRC^]]OIP1cK=-M29+7@D)[f+:X_6P.@+.
:Y2/E>-E[#+7S/^W<L(d^:V#;>,F/G^6;J366J<P/Z_R(GW=NAM764P-,g^b(G-9
<Z<ceO9GC/S-b_U=f?43/RCU]\2;B>E2STAIEZdRS97aM^K(MQ5IIg+c2.#4XR(e
EC,=\08T7C#PHYB/8=)DcPTGN^8RXX)R#3,_5MHSFU/>2MGF4=[ZY;VG3Y9Z)a]C
f@P<;dTde?QECg1Re2cP&.)/,M+W.8<_O^OI,CIF9;LDNI>D3YN:-6RUP7_T#1Y)
42&.L4>dZM2(T/,)56[4f7d(eS4&,7\OD,Q?EWTX@V_R;5K5M^#GGJRTA2(fgVL.
>/KT#_U1@H[]I+@Gb1EXf8K.2)FN,2C)>:NTQ03=R,&CAgYX2P_7(aV0g+g.fR?\
2F637gXbdCPJ;9:.7:<6bHda<VN3Tf008(bV;@Ib7PA3EgV.#^MJ:<6JYa^fS=\(
J=TTg_Pg.M41Ne>9cdB<#_e54/6Y>c,KfX6P\LVO?T?L[5f.[N@)9DC)J\84,2J\
B#;5bT0J9c&25?_8XN.V-;BR&&B4d5>bc.+Z?.0e2]:)a@30X+AR-)4_T1&O;.CV
C9T+QbgGE[P19.5K/>C;B(f-5&603g,Dgd?0VBNcYYAO+b:G2=WHCP&,2NUQGA9L
g-_aWCS)D&DMBG+T;1?O8\fK)=agNP>R&2G;Mg\FUKY]9V#BgH4IJ<F8WPABJ>W:
KE]f>E6M#a>L&#8G_4^]S#Q=:8UVTBDg-F>Y1Yag0;Lafd=E?c30>?ec64M;5_7&
KQ((_0PfNgSU_W\VNM0G3?,R;OS&\N7N[P6W<OF?bVDf#N-6_Y(Fd(PI7Z9;UDTZ
f=H;40.]#J8K4\\CB9+29#;BGLWL=Pd=E3Z]XP\5)g<20KL\O6+B4IQX7K0D_Y4U
[3ccDM)H1B^)fL#-WYNG=Ke]/HRTK^PKH(,BTL/c4.,c\J>H5=gJ7P8FVS9TbeNO
Y9SJ\IC6<]2L-HG2EPg_^+[]O<:g/OgdK[,-YPZ&=d,gE0Y(FaL\f&#_Ug9g72f\
Ia\C)QY7(/)VeeN3.;P9f.5OfDYb@cZ_G7QI6&>K(&QO^DKbW+3:+-LS5&V,eb+H
T-D,Y1+[,E)cD8GTG=5>-.YS:97NV=]O-9RaK6MQ^g^VV&#Ja>@]H5b8)J7.S3Pc
VOAM-9ed;cHLOW.)QZ9F@M/,[+(e<KG[4D?SBC3IV4?47bPDNcM=^fUbY8Z6-JMD
/IT^cC6.6Fd</N5/P/cB2QOb31JB858TCGY)Fb5#T]07eNe6##CUa/M,6&aAbU^E
<1G5a@N,GWPdKb_I#F#\USW30dYBbA?RH55IJE&-XXBU0eV+;=ITV,A#9[>[Vc3L
&B-/e\\GILY]REN^g.B6+\,LL4MH1Q53\U;B[.V;HY9^F/</\Z,P2]=TB(HM+da6
JQ/[[9aK0C+?/60;8afFfCD1Va^H#SIA?Q[6)GFQ:9B8T4b]^)),=-J&gLOg1#T8
gdOLda?2;UTZPQf9C^Y:)8FdS)M8?[\)Wfe.MB+^&0<fg]DM2WHJ)ML>?+RFfG,E
T[.\23;D0&gG4UY>gNYSJRU;.E+>,@H]W?5K<J>?.YIdU.g^dd;2@;Q4F&(.JFYI
)P9dd2FMR&1c]OX=5@&GK-M6LEGc_(_80T?49gK35RBR_FVJeC#M5Uf#^#fKHA;:
0W,.T]fE&Z?L@7XCR)14H:L3?dN8ba<.Rb[FZeLcQTOYQcLF4_H\(^F7-]b@EUZ2
MHB+3N^L/-,eIW#:_G:CbBe0QE7;9Ka)dJ#M+B9A:eYaWfAd0;<2>IQG#XV>UM1Y
Of0R@\5;aIF4RC@ACOI.M9AgLB\3eO3acf@>,L&d^d;&JeUDLgP^Ze:8V)NU6V&)
D0BMX4VQLCLfdK_EN#5VLAC2B-U?@-P>S&X,NFA?AE@:bOJb>4gff60fLSg(/038
5JH>9-VCBE\XA@>S36,\CG&:6H(F^.ASJPG3[b#aFc16A/VU^:4L]F&HTPAX(QPA
dY\>(P.IJdR?bNf@(d[P+OfJCF=0g6&9R1YU?+)QNB<aVZFF;g,2E)IR\RG9,g+e
(\aTW>dSLBA3EY@NQZf03FN_PfX=[2g3V98[?(JLZaTLBN66[>BJ1^=3?2ZTF1NU
#7b8BZ[[;f+Of+gEFe9Y4V,03900#F+0>HI5YdY0B(WYS-P3K=09F_5HgV([NQbA
)GVPIc6UG_XQG73BDP=-RU/[f/LD22&;QMV.EHAb@Od<dad?2+4M,#aY.:04cL\e
Pc7(Cd_/HX9^/dbf9G,UG>&F[<EJKOF\OTJ6f;9ZDb1T2G<B?#\_H,V9&LH692HX
>Q0B3eQ4=e8S(4B[2;2?O@e^NA_H<^;\T&S98S@SB;-IY3E2#U?OXE&@),?cS?<R
gGXeMP#P\=A^5FX]df50UXb>PfWd#Dg^_C-;(7?:21c8&1;EM;:5,W;T;5)FX)B1
LSGE0XZE.Y2BFFd^9RSJDg0U=4]aT#+=)#OH10E89WU94\gLU^:-Y\cd)g),>MF-
=\?@-T<Gd92.2=C)AJ5UE1+S^GcT&DZ9RNXF#+HSD><;O3^B?Xa+HaOEedgQf.8W
LT4/Ce9_>PF4JZeFGFOW-1Y=@UH&5K8gM3M^M?(\fe)g.?Nb&S_MdfO?MX#Z1KX]
DIb,?3Y@^@6cXIE;\+9WN@f>Q(<1HOPN)c[.8aB:9Tf@6NUeK3;d.6SB+_5TEPLC
<64A^0=G#@?W]dT8YA^B?M2fJ/->gO50VJ^;XM^22&4<-&>VX?A9N/5c-L,[5\g\
^?A&(3(&070/E)^aJ9f>?c-\OPNBff\9/=2P@ER1F3V[Y=2&-M([S8^Adf,BW7QJ
:=a,3F[&07a@(#7D.HZMe5OC1&b1P_CB2QN.7ZGHE>TH]Q0.RH.g,eIZH/PRRJFL
f2.&:a>B-FDa[M6S_26J&c@BV&+9YFb-Y=&R_VAR=2aSCP2PXaP+MF)I+C/V[2_H
g93</Hfc988BZJ=8e_LdE>(8CF@O@0N[+Ua&1S<5KA(>\[.BF#V)8?4RA1X&IP.Z
e2TMSZW#4#25XILN&8BO=9R96<RD#b?S]\--KGE+FbPPNd?^#,1\9+)L=3DVXSGL
VQ]?#g/\QP2YeC@:<eaDR4:15O6T@>^Sb+XXG7\J#Q1.;;Wf=NHf=K9_ZZ+T/B:Y
9Rd?9>KO7(N0H7(c@+(/B/Yb-<ZKNP:]=b1&^=H&7gXNQSFBcMTL;,7eYS3_b1]g
_[4[L+(P2O#T,&G9_JNbYEd2_I4N>fC@/a:]&_51H.SIgX/6fX]09T-U_MO#>QOO
W8@#K5Pf#@DCT:FN]Tge_80c1\4LO0Gb&6IU;Y)Z/5IZ=X^(ZS6<<YUb6CJ2+?XX
E0cHLC.LaR][9UJ/]e@YEK:L?7ZR2R;+HSXEA2]3>,G>QWWKCF-)bLb41Y,)+_+>
C:_b+M,N#H)CQ;13\T>E+N<+UNUF#&^)C4:6H-9Sa9J)2.TXWZL6UZ)5WE4g9F]d
HFQC/48P?UHI5Q97[R_/5/43PKW>1<WLUQg#47,5Z#ECQ_KENQQRJC06V\MN@BR5
?b73a>aX8gSXBAM]_7?cDB/WX.)-W0NNeD.A&6NWZc=NB5>+7^+e775CY.6BG]Y(
F@b4@@A\(9WC\Z/T6:T;3(.SI.NSQS^V@UX^H3c?5QLfM;Ae<I^_RZO?g0UCc>&Q
Y3C^XRAc,D58<+YE35Sa;54A]-O6Jf.A=fUO@DI1aQ5WU;e3[#\VAK6/[^0.6CfR
N0<5Ib-N.bFEL)3.8U<-8C40=5=L=51,fE1]L1<)0WR=VF3E^Pe[P=DS=)W?JOKU
Y4HK7W<Y_^Qe]gf7BS96P4UER#cB,KfaA&8H)RfZV6UI[/#11A=BJ/NF#6efJYCM
[V)EQ9F,,gQXC2d4fK8-8+5,9;RM+\e3dC4YYRF//gW\=PdVZU#+K+d@HTB7A#5X
(AG8<[2+_.^)L702RB\@A?0S12PP=IfOC[ODXd\P#4/P<Tg^NHOdM3;A?Gc/1\gU
P?B8Bc31@TXT^<V^eKaHQ]cSZ]0[^a2:8\K+Z_D0K&/ZQAB:2WgL,YOMW7KJC0X\
,H1E#^08R&45Z7fTZg:F\&K58P]IH3O2VVYc20I;/6cK,)22,J@abAg7VEO+9@^)
afU_YQF5HEQ&9OeUgc:f/31DHL^&;\=0_4>ANP3C80C,,BXHKBACD^:5fccdcN:\
YScAaDW;)Y_c]fQ(a4I4d>+;)8A0N5Cd+GN1BWT-75#>V3cN,]#7ISFR6gb>@Kd<
CLg@c/?/R9KOHZcNUbGeT36VY_F>8TPDI\d0]&FO.3<;^.I>AJNBVGVFIKGKS0:P
OcJG6)gXXA5=JD4Z:e-(O_4BR?-?;O;68MJYF()A.0:QYf;R<REC6;N+H4X,0A&N
Va8<J[MGL[9DL])YR1L-G>BY]R&[#MC]^..9>1<gCUB=]--F8\J-0#ZYIRNR8KM^
a@-]RI&_689OXgd48RURZ.I]+;6a9KS)@04)-J>Da6LT;P9_ObF?eH\?<GO)<=dI
74Ob;8@=UL?;./5VPYV^IJ]-K\LZ#GWJ^A6K..H7H;3Z)[beaND^[^/[6+C1_eJA
.1)MK&VG=6U73Cb\=43Ea0.(DLY/S;^FITDN]G.-,T0&[_8(dQFcZ^NS+a=ag4E^
TeEASIH6gHWC-Ma[RBEQH63CX)Q9g?6M[JCLa7O40I)+QM,eHbL1]DPe=L:<FJF[
D4260ME>ZL&HR<M/ZEecSc:-ZRT[HOBZ)[(XbR<OP2_WLSW>FTMN5]c2g,=N<&D1
:]F;1ad0>fH0)X:]5=W/J.,#9O#dN795We^SMb8]T6\9OIOWX##2+c02g4#R85gE
F<]bJ-X0(b>I&Lg3T]Z>\4ATOaB^I-^7O._:-b#+B;[>OR?1a?3Z8YC1P_RA]dR@
.dT+XcT?FY>dR\bKO:A@,-3EKNfIU?ID81a4U(+75MU@9G7dZ4MTIOd5SIM;Qe4-
7dXJ2dH3@bDT+/bXEdc7YCONWVM#-?B#7Z:C89G77W5G1;aKVTb+F14fDN<#MC\e
FZ7Z-&aIZ(Z4O75&M7TGVbBNMBQ<16[D\IZF?6GP\<MOUKOUL@M3VEd41)+#QWON
7^f,<_&d9:F?T7O<NWA8aXKAB0Le(=a?-#69ULCQX#:#-EeX[Je=<SG22\dT5Kc4
,FWX_0V9EFUKR#BKZ1dY5[3\2<O.)S]b@c^/UJPTT--d[7&O?@UU-&GB-5O:2=PY
\(K=<SRR8LSD932ODQQE7-2XG/0^SQf:#_J)<Z20-eV.LTQB+G.P9=-PU6V,+7ZF
WYCa0ScUYNW/[L^F]MGMDQR<Y),M,,MWZ#0]LP\(FNR?d/eQ</eV;=L?@XU1IW<]
U?)\CH0H6c),0e0/QNe37EWP:Y6cP+YW7E1;AGHg#22eWb?@#I]e@V^46[2=e3@+
_,_cBEM_5:8;MPN.>V2+Z&cK9_8719J5>W]a;0JUL)PMZ2@JV.)\Kd=.A/(OcBJ6
,bJ_VRM\gC7GU;\W8[WNSOK[<G>9<M5Sf0Q7)GH8PZ(.>FAC=S;TdMKI#Z+#O\[Z
XE9F)F#-:Q^TM6,7bf:FQQ0KIR,=WN?SeaPV_fMQ;G\/TP25/df4AA:L-g<aTQ6_
,e6@XbVF3,95cP?^/H&Q\_VR4f+80&LCTTTVG<?V4^&3;7IbWT6]3N0ZX)9[R<X\
W6YBP:M6,+O__g5]Wd#B(?aEfXK?40=Z5?e,E1bDXT<CGHG8./_b1J+B]JMZ_@a)
8aHG>cOPDH=@C#X3(>bBDG\/b/=-_;Je162QX;g2YETOV]?-cJ(YX@AXZ@9@XITE
N+TXb#bMZS0GNa\9;>+&2g0[(+P@#P4ON0UMHe8H[#?-G:BfdIY]X0XNEDFbE?L&
e>b.S-L30:HV;DJa/_XD9P..ERZXJ[YIc]<gC6;3G(:JI;45L:,WMO6\1;;Vf.8^
.-3[^B,fYIb=ab3@ML;-&-MU(J_U;=Sb6JY36P387#EAOO#^I:EQ<-55J0]DF)1)
Q=:O[_E1LZE.-G(8/(L4E9E.W;:;Y1R&,@X&I#>_&&U<.ROcHR[@__d>=NbT]GL<
W7GA+bb[)]^@O@7K.B.MDgI/Q6/-N,I_)VS+@aXM(94DaP7:b_A-8?EX2X(>+R_9
XHUHGV1K1G4X2=+I4TN/XH?_9\ZW+OA-MWFdK\>=H/LNX680-9;Z85?9+:>73#.W
8GEX;,4a0;LQT>OVN=XSFB/13Xg2YA[X3@PF0:fd?E=-O4Re\VNH@[-@KVBY&()+
d\OU(;&g2d\\+b/DF2\,/Z2(0a(B3b__0D\[;FKe7K[T?&[)d\4==_2?F8<DPBdd
@VC]Uf:0GeM,,A1V.K7@?7A/FD)Fc<U6K6TLBWES496WD3B,-T]NCJ1B.Y<-@\:2
#2P(U(3S)\WTP[ZWMI\21e.:^7>N_MUG@&2&b+UQ3&9N\6L2fY^,0R3S/c#X6UCB
BeA+JG/d1\_W/01NHG_S42=ZT^/[g+[@C2EBgH3N-7.\@_>;bH1L[6\Fc(fDHT;[
gP].\,fDR=-&C6DUG?<f(9U>4N7UVeYfTK@7A[I<Ea/Td)cSA3fCRaM,,>b#B464
)@];7H:+?QG_C_#4F=+6D#7/^C&f8?H:GVg=>KB+60T>a8?c@YEHJA:RTN5_gS<A
AM41NSaUIg:=D,GCZI3T+N]d4Z^&G8GB_UV=_[SRO:A@;62?X^9F7Q=9;_R^J&(a
R:M3Rb/eT_3+65Vb^IN,#)?B&KEPKWBPJD5DE)LL1L-SWb?3&&LRP/)/GFF_1=PG
&dFd8QN(XX@SRTO+Q6B;bAYL(SQ-T,JM;7N+/RM=AH?-a7551/BM5QA0>.YI&FGJ
26aHF2W0-Ydce>>3\?THJ@W-cX1/T?Vc7[f]N@DdV3).#(-NZ)LMCK9#4KS;QObL
[LP?)J9EWPED-D51LLfId-FI<T-;fT+643N&C+f+M6da6-OUQeIH<f8@-</dfX5<
8\a8CS\ZSL07XMF,5Q00(Z<RdWCM&_59?_=dPV_YT.UCFFHBCeUe.:HE>02^P:Y&
7d-RPX=a=VLI44CXY:W/V^d.V?J:^5BF)12=[B+.J18S7JXF\QJ^T=PFD:&ecF1#
TJCJ3D.]98RadDC_UBP8bFCMS1+L1(#/-S^H>VW[ULST@3M@)(Df9eN6T^a95OOR
PM/K@7JUE>_D,@,U/QaKb3^OgZ.d/(T/FLfBYgFb?(a(U/KS@G\V<^dg)ZYDW,EN
AS77b/&gS7YOFH_@SdAGeceAT^-((F#DL\@M[@T@c51=]aJ<==CQU,S(CgM9>bDd
&T;4P)@e.U[A>R(4c9_/P[5?9XTTdMN]E/86@K-9G.JE9cS#N+YWTba)G(-<<1=f
&XU-MH7DTbC:T)B/)OLb,-S^dW8G:c?Z:(6W3>J(b:0YTD/TOE/(M(1a&A&Oeb,0
5:B595YbO=M[@B)\><E:fPg/=BL,(/JS8(NSU5gg0WKXg?T+.Z&[6g-?CY8Hd(b<
6GV=YH;Bg:NI6]9^<+:K9g)P,(TbYD0_-QL1JZe)KZ^&[?K.f2N/_9?Yfe=b(#\_
\8>KcA&6Le2)^cEa/>[VT53DU-,:_[O>^>9K,[:6CZKQ3NeNe88AVMB^RJA?C.HY
2.A:Z<2A6I0L3&?EcURe;C4cK@ZJ+Z[C6\HQ@.4RE09XGO/[^28KCJ.[\[WZ=5&,
\^bCPFd>Y_5(1IELV/>Ae/_&fG/JPfE,:0/:/6\MXSQ-M.3bT)#J4CVKeQAG,#QW
[GX2CZJ4bWHBc>_QED>DC),_UKTZ()M6XfI[X2?afBU0:K(SBOUgR\\Of+5c2QKZ
B^MEe77=aF(:6@Z\F<B)?RCcS,-17#+07RYf]KPTbA2Pcd[OJAAeQ#H^JVSX1))]
7^VSg9c:g6]^5)]6g;.=#/GbY?B()aLT1PQ0?F[O(A>E\QZ.dPQ=8WGP3#[^M0-;
gAed0,1&])a6/S_Kg+Z(CT/V=8WY6754?]8a6:W#\f+Ua6YL2Q=<?d]QA3#BYHPX
>50Z&&&Q4C2MOZRA=aDFYd)c\E=OAf^bH&b]6S8H2M?QNc]:FV[>+NRIQJA.=3+9
FWR-a]:Y8K^g-Z)09-1891bgNLW??;HHNR4IceK2?6/;UYIU@dP45fY3J+D65eJM
;,-6XHN3B5T6O/Q=6GR507S&5RZ9A3\.3?,4B4>8a^I26UZW=V]2KJMS>GG:eL<P
_JS+a[&Yf2\a\8Z<LOY+Sb83XH5]8B^:75?aE6FFTFYS[T2T7cUU9N9#9Y>-@f+?
0VFD@gY[HYd3-IH7JK((=;A-D8G067SS<V^_IN9-dLC1\+,X2b5/26Wf^<Eg3c25
)H&V.7XfV4>#9bC;Fa#1Me.aK+3gc?JI;4<<<D<JC4VP9I;g7N#0cYPY>NH1(3IJ
^Y;P&)=<DZKC?(8EE5eRZ>.=?a2=L)#SVR_0PX#bG4DaS-G#e5ZB.W8]^QW@Z\7Z
,NJM8SE(F7^-CUSW]K[@,d5eY7^#gW(7dA3>R/_?0P->-d.T-^=1@(\O3D0.)09I
HOG6K:566(9AD+.aVO-BX.D3P<XefU2JY3H?:)7M.ES,\Q/XPXaXM^.T4-a0];V8
Da<aNN5061BY0^A_1X)4@Tbe-8.Y=TT2=D;J,.dN);L\29PN;;WbeXYAFT0U\3D,
?2KK-/T+9WS\NS>aUb#H?R)<R19YH_NQR]V4LL2<=[Lg(;\B0dW_3QO]@\NE_?Yf
0_d/;_]36P@/L<+NI=ZAG=(NTDA3f,_]K-f.W.<\Z+)/Na7L=?WJY77;#3NQ#_QJ
)-3@P99#1<W4]+,fdeZN?+Z2:<@AE9\)>E&EFbG=#=WUEI9GR&9#0@;W2A8?_KS1
[+gXWfN1BG9A5fa1Y&(,Z8__YFQed-.O]8.\?-1,=8ZDa348UR9^8Z<\0<a(O1F(
(-X?6,2R-c_(6ea@2,9A,Ua?3<U&J:YLF=a)fCT:fLHZ6DQW\>M7/eaEa6YG2;a+
I7E?6Pd[#ND@:E_5Fd[/@?[faYd\A2)X36Hf5/g90e:I?&?&.LU7dcGY4XcROB[a
4.]?,^d0GKM0ZdQ9^=N_,8NL&J<6+D1&RWD9XH7NE:4S4@fPOe]-VN4S\[K1A)Tf
L1I/M=.#O::(UNC5IR:>S&_6:DPB4VHc><VSg[>V<e6Ga6/&KI^5=CN7#aAg3B4f
92\L&^:2+N-SO/P)7cEWe8@c&eFA;-8F]I@(PJ@[6840E5ZfA7G_((MXdOCHGF\7
\/(Z]6dMW\e8ZFRC85V,;.;3=64Q;A;3\[_cLFB2_HYEP8(Xa5b7W>-WR20De<J\
g3RB]aPWKG<0?7ObXS7J1,?/4d6.33dIVAVbK2GUW=NS.G?<1?e)JJW6>9e6QQDd
5GK/YfV]@\V\A5QUNGFE]Fb@/J;Y)fJ]XeJXJe9=:gbS<FX[NCfV@XYFC/\#ME.X
3C5Z=H_M[1E1a:QI=WO^d^8)?RX2a6bfB)HJFeb+[7A;W(UAB_<daEE=HaD8f)a=
EBLgF>GATb(,(8Cf;WV]QOAELSd=#)RQY6Y-XG-X)Z;)O/IB6dSO#2GZODae#ES^
e91/:0-&,?:P>EE(Z92XM+B[W4FLIaW2fO,&#(GBNE4/Xd:GE97_O4I,AG(V^a+b
)(<I-cID2eGeL\-R2a\T3^^P+[0bRR<^:gMJTU5Xe?]AZ5Yf55QI,#Q[/cHM0QQ3
4bZ1FD\#K9&b1M0)B[ePM:7QDYWFb.O99).@F4)KB#;)2,FX<33.bgO<^02L1I3[
B.aM;=c:0/#@bOdZd/:?b#Q=b\g4:+.9UG7T@aZd=3E3^=J[aW#1L/-:GUggX4dd
4d\a>Ude:,Y+8>(0#\\g?@2K)3D9\:#STUZ;<H\abVZ^/54<.=CKQPg6>^19D3Mf
-f(PEE\Vf]f4L3V\DT#[C?_fPZ]:&Z5UEOH)Xg8NMd-JW&JIWJ:D<8PM4@914LB8
/=d1B8gC8.TA.gW7E+YSNI9#]0d)f\H=H-QN-Vcf)#aJ//7HcW7R.f&7f#R\+EUZ
Nd?<R:8]_U:Vb>Y[W@/47e#+CMERag>#VMfQ=BV@Q0cQ5Wd>P+J)T8NcZG.X#>TA
)1O<(7GXf<@G_:6DbSK<faHIc_>7D2/WFS0WVdDaZfeZ^&+Seg_R:58+?)_&?5RC
e?+a_2VWc97.5IeKPGGfPUNb1Ea14O?fK-d;#W08/8SE6Nb6e::J3g_PTgV:(9B8
bJUUA1=.NG)HE@3/e>O71S&&9g\@.HaDN21=Xc5CU89<4D8L;gZPUKJ/0:R[##GJ
GGH,\XX)>>MV#Z3F&-P4()M0d?G><YSH3N&6O1ScN^^ed8C_A,8D]gXU>Ab)S<AQ
HR2L?W>Q8&S_.[>Y[;9HDX7I#Fg=DgL8+G7E4_37V^SJLbJ,3>CIK-&12CgKBDK@
&aa>Z5WK>\<:eQ^9F8)J>UKPLS:=DR\3U?<[#N;G6::c@d-@):0N@TE0X<=<H=3+
-\\GMY_WK54VRaY2]I8S5NLTWe@TZSA^6F7d;&1ANQQSPe3N,59]@BKPZ2Q+e\45
eP#\NM)HafJd.e&fRJf)=,2Qc?\C#BP#:<Xbb;GY1P+[:Wf17VL_1dLMT(5]dJD1
?dP_M49(f(/+92-B;:UaH2<7ZR\9N<c4.:40\4C2Q<Y83P)A]c/@7BN6SY)>TYX,
JVG(4>0ZOE[&84>4Zf^dgUGX;[Y.R6DH7XIT_E,O(_J;=>IMdC2@\6N#J&Kb7#9I
ZS5:Q(7;]V_A0Q((/db<S=0_8(NeO?Z)ZCF(S[=U)IF>>5<H]FF[eRgQ>2#+O:+E
F:6>TM?0W=X(0&7A][YU>2I[f)4I\;S,9\7a5R->+?&_[b[&C2YDGEK?JAU)TLb-
4<,g9W]7gQX4ON):c>Q]0==@G\G,aSP8JZQ5(IHP[a1e90=(8^RHgNC\e+P@K\<,
)/R2JbAWANS=#-UBI.:A=)TZPDY)6N=&7-LVA5D:BfE4Ofgg9EPLK(QEVf&:Q)TL
N-8HV:U-CE,&cBf>9OCX[F./8P,^USe)bV8UW:NYaX_A?UbF&/B0PWZ<XFdH3K]W
(=^^HbQ6.B&72Na5\KGP>OYX9H(a#U&?](fe#^TX3W;]O?YMB5aDZ7C^/0FL1FA]
\,9<@/,.+\K([6Ub>^LYJF1TY#_<Y,:8>]SeC.\Y>-)FG_VH;HPW_D,bTCU_@RR?
>V=)F?HcINX14JNG/Z-8]8gFF-G+;@S0INT\(M1L.G\67,T1fXZBXJ3YPPeL4R.N
VGR4EM]B)B83Na&>>L_82Y?C=+a\^9YOADGg9;VH]dGfGYI2\9/;?6-1e6H?1CE9
^Mb:8a@I_NG:Ib;I<NZPc59dPKHU_aaT41)4ESOY@S97#JZ:XNC7?8W<TSU0CAWG
dD+:Q8ecN#J@&V(-<[60EBS0Q&SK2ZX?O4T]c6f8]Vd+6bH,fE@D[daQ:]4[b)=]
7TO3/dM.TJD/Oe=QL,(2YVF\@KH\1?Q=1\PQ:(f8Xa1NfVd>-MY9J4FF+E/EE>f3
3R:@56U)a7C=_A2_6<^O4:IVEg6b+OCGEaR5NPW=g5B4?a#\HK#)@:9E),1FX_8a
[M;U9Z5#NW@^<g<(W22:8;V1D6XOSE7KF?gN&eTTJ8;(X.d:=)DV#[g;\+H,3A@b
4\N@R9([B8LP7I.GX[EDZI0[IF1WJVAADdU2L;+@3-F[L;f48F_abbH5eD.ZJf+@
):6gON=-G8UQ.2QI(DdEXF<8dLa4NOVQdaBPVXd:TQMF+W43_<?)GN2Le_[?e<#E
_>a@W5D-/d6D3NG2>BVS&#=L0B([]A<#,)G;XI0RUJI2H2.g/BKIM6I,V.,#2W4U
F]g_XMDP&eRfP?PGf\=W,5/659I(7AbT5G+TedJ0aeZGD]K7WT5e(,2Cd;5H/6\e
E89(&F+/4>-[N-bD;#F>C25[L#1C<L7[?2>)+?eD;dK##K0_OceYTXe:MBgFOYb_
GaX4fZ;+IZHIcC@NYH+2E-.W#(>;OD[TZI.U&H?5([Q-[XY/SXEN>43bDe)@NM5G
-51LS]FGgZ1>#VPLB>Z0T=4+g[<@;Q<cP7J=+R&N-@H4[TVF@-)):ZgX<H0J3HBg
F+W,_/VM;X7dcZ[[UV3?aR.Q?A#1R.KfV.;g^.9?NM:5GgJD0UCeGSZ_S;gdM+TW
=eWIG<bKJM#NLTa26D(AcO7H+I,#9-5QM]>].WH&S#@_Z+<+Cg+[P[1fF=/^HP(>
>_3VQ(B?K+UWJ2B7.GN<U1I/b4O=@O;OL?\>#^E5.?@_7K76\5WC4L-&R]L\/GI;
<aNPG/K80,B3[G]_d>#6&RF\.DGC+XDJ\@KX&/F,aF,1_C6VGISVQATdU\X5M/0U
Xg?X5^U3)KN<K&FJ7[M/^.:AY)V3?NP6E3H6QM@bJ6#U56X_V(0E&7AL>>VL8VYN
gK+(#VcT@4RRaH4Nac@.WIBHb&5,)3)Ha,aS<9T(Q)RPZ-^PG+E7eA5?,QbWH9Nf
adRIf\Xe?GN7OQ[cd^L]^<LPG)0D79MR96U_]>)[66M9WH9[BW#>FV.af_?7#AeR
3FC>,^7=[R48A0&aP/Z?G(EP?c4ABYgQ-4[P?LNTPMG@_cO<3/,b)e^)8TFLcT\G
@\[C<VYd0UHSQ5.A/g^G,OJg6&EJH+AA/S3>D9T8;3d3,,E#I9L7)&&Qf#I/<e#f
RB_7O&CS)G1WXZGS5F8S=8^We7>Q-3,]>=(d@</<[;:)9H-0P<a>@^7Y4e2Q[B(8
d(BbNXa?bV)Ed?LLe&WOG8^7F9XQY0g)84#JNUR&+DaR4U)T:@J165L7]U3R\#F3
bA6X9:gMd]ZGJ4_^\7-Ub#I2UeUJJ1OM@\+YP585@H:N#K=NPPa]685<gMU<58XD
[VXPAcTX#M<_:aa8@_SRKS(TZ.]H9]L[c9S\5F#SX?ggV@#@(M5<fUb^N,HTBG9J
41.aWdY]79c5&4KGD[(d]W@#fC84b3PN-=3V@[5g:</9A_f7SXVf[H3Z=GZ)^]2)
K+[CP\(]IXT&I;.Z\7<58M4YPX<L^cM]A^O^[a<]QVfW?Ja2Z2A#4E+7L77IV,[Q
WN@CWJ>:))<+OGHW_1W4efB0<a_ULCDIFUQ:^MD]B7-P+]G;PBZP6O1C<:46EI2B
)e^W<#Lg7bVTgE=5E>)aS>GOF3#R?;dYB4C8P6P524+0d8#ZYDfPeU/#8+Y)Ca-C
d/I-_T=X@X<d>LX/N;.:fZ9E?YJ\(=HYOfaO@^I58XLePWE[@TgS#4D9OZ]H7-S\
/S@RNd58A\^4aS[AYS&^f45L4_]AYUQVG&MH[M+=E[UGS<,]F&=PUCGUDK9ZV8gI
E]0-f^d.]GYF^KgaEZG<caA07bE9H99-d+Y1d[;E+SAG<0FL?g61RSR@U<4CggYR
S^P_-Jg4Q9+SX)UOA7QPb)CK0FE]T+FXZ(#.2BK@-1Qg>EMBXK<80&g@Y-DT1YHE
bI@\IHUEBDH)RRR9a^?eHDZHdAYV?-4SZd2?E=U>)Q&Ce>R0-7A56fO2BA:)AbLE
DY(Q=e5eZ3&f;:+(UgH19V8RVFf.f]2,7CSP67P#)QB-_^G7-8V<NcI#YefRe_cE
TKfPPR8SEe/<OH1gZ&EWWg<7=T@d+ZI[TQ=_Y[//;;cGTMXNMC-\=KM#ad<,Xg+_
^C;O<6]H3LT1MLPWDa0]OM6AaQ-9,,Y:feUc2^]V?-e7,W,RQPf:ae]d=14E)1+b
Y_MIT\7LGYG28TZ:M)0P[b.3<]PGQfK@43K#.VaTOP(EM?5cY7/L?^\E>0SJNB</
<;7dM7?U1)S6gCN#TB[Q&Mc4O[\HO0?&+I\=eK_=?&7a2f23MFRf20=GOeJ-YZB7
0(_D93P&&O8#\1@b7fd]^?:IcX?Pe+<YWbe4\XL4eE)d).1MC_;YE^Y=2aW+:9(,
2,,g5)&KAX+PQU-Y;d.(>V.^[,Y8ONH;48]11;#?9\LJLX\U>;#P+^a5J(#8a;)g
)(.@;fUOJK_+56OIP>b&&JK\Xb^3f2^M40ccDYWC.fdM1I-<[Z@MgS1a9B2b]F,+
6D)f1G+/IR[,-F_TZXfc&cdD._A4&fZ)G/RDY;:FC1.-EeB,>\J9)15cZ^VDV=.Q
:\?;:VM8-C+,\K=#^BEc.DR5(3QG&<a&X1>#<(C1FC3O3^ZCb6C01<0?/ZT:9UHD
D\KO4HXFXN4QN<-ae^eB&fZ#ENT^66PU@1FFX^2D7d<#4J5>bLASY#eH<T\eXQ]+
e?4+M[A)ZeCX/QdgCL7:9eead>X&/@X=LAH+CgGI5R3bMY^OY1T8f_67RB=UQ4(L
+Z0cVC^5QN]e[4d]8<Q=L_V(Ecg&WZGV@Pe@)MF/XDI]K@^L45,EZY76H4a,]4U3
FWKeg>/MQWc8[WPF9=)daVaKXDJ6a4+Eg]Y#gPbF.c7H;4\g0<4XbB7I^eBZ7=GI
@TZ.Z6e+eeMXeD[I4f<CQ>G)RK?][0cQ-Q)OAS=KNgF3;-3fdTXTWMV>Wbc-?G];
?#eCe=CB.P?UH]=UAgY@^MZ&>O8GNGL4.dUWNgCKM2/=Y/3YE6\:fcV?8a>?NX6\
G@Y\K58I&R97QP2@?Db/VMQ^G#6+?R83.OfU-#09V_\Ed2^D]IS[6#=B6L-3^5M:
BT?G<>=D79N=d8JRaOE&=1_2AEgVN_AN55DSFGK:20CCML1NX)>Ua\V,J;KLe914
H]Ke3LT=PGfML+>][&-V;ZfF9@^c]cH>3Q5MRH#b4U;fa<eO6/#[P6,WJJCLNY#2
0\<XJ4L>SGB\4]\T]SgEEZf;.KVG2QEZ,R69JP\T\)L>JEBAfQOX@f-/OJ,D3fa4
N(A5\998g7XHRXH>M.?S_\0Q.E7Y]ee5a+=Y;&F-=Fe^dI7)U/8&IQH0W@/c#K:e
2+cC6\N):&#53Jfc/B[/(F=)ZTXCFUW7cgZA+aC#9NL?3KL^Xe,(VJ_N+21cCM>S
Ta>TE(J[1[3?NH2;UI5U59U4X6)V<aNN<BZ7,3I;R&P?cAOgIA:aNNNd]HW]c4[,
9)XDDG?Lc71N<JVdKCdCRegTUe&(O)=ZA&>I6YUeDgCA&840A#&WEYgB&Tdc^]EX
65JfB-UZF3RC9BAP,]&)KQ[65^RP7Y7gS^J_-Z(XG^^#4WRM3+FVc6#0+=H9CCd0
:8XbG@Z[g)c2[B/)GM(gM?^V@^+<4I9TMBa)&JbQJPI^)PfY)9E8KNVVb_[L_<dL
g[PLOg32d._RMgS?b+M)OL[UZ/>gbC@O:V_VX?&>]c6@^7#;YV)2^>]+MC+E?CK.
I-_+)3c8ba.-TP@O9&P)ea<)GSbN<Z#5HCL/MEB/8T9]YB^.3XSC.gg?g#J(KV86
1dMUe0Z+HWVQZQBF(J#_6T82:WY[R5\G]D_B/N@=43=ee]b-AfW1OCBF(R8:H8(K
Mc[[_+]8YV:(;_@<#URH59W_5Ee[HS,\Q\,c8;+C?G6f.Fe0_K@JfaE09K)cRPSZ
a^=[S18KK2RETZ5+8]A@:P7f0R9-ILJ,aP4Vc]aAdI(d[-cF3-(?0ABA>g05#)>W
\X-<97X)=3X0d-HX46(:K?_9aW#66-9-bW1,bVWT&98R4U&V9@<Y#-N)S_ZK<^>2
55N94F4WV:--\0V^#DTEH/,N8MU:>IV&S#(;21[^8=->_b;B6a9TWCW64#&)/U3Y
(\<A@X,4PLFSV\L]<XBNNAQ+7RgBF<CJ+6\c(E]R[J3:,b3f,eW.A,f>X0^0+75Y
4dU+I2?A:2YT8L\Fe;gRIL+_5Z1GgHeF;<Qbb7W46UACV6<]S0&b1d8IPCF?07:e
F3-MBd0E,](aeaJWF#5&Q<KHc6@_QBA==9E3<<&Z).Pbd0.SJ<[K1A5\0:J)9R(L
ZK<G1^>/4KIH#X7TF5(VH/\?c.N_b]UW[5OUe/I7VFI:RVH:8Q]B5fd#(gQI/L)Z
ANc3>\G#>TRW03R[VE,PH_2-EN3+R3+ed]b>7-Pd^BU[,&:>);PJ1JK6D;Y[(N77
a>SKTFDX)1?3<5@#SR\6Y,YD:(L:bdScbT;E=E6ccJc#\\&-#)H?I\O6;=I:9)B,
(:[JaPG<&>EE.?EMXBbRA^PXH&C)C;d7S_f4aCE2[b49<&HL0Fb-Y1O6N$
`endprotected


`endif // GUARD_SVT_AHB_MASTER_UVM_SV





