

`ifndef GUARD_SVT_AXI_TRANSACTION_SV
`define GUARD_SVT_AXI_TRANSACTION_SV

`include "svt_axi_defines.svi"

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
`define SVT_AXI_INTERFACE_TYPE axi_interface_type
`else
`define SVT_AXI_INTERFACE_TYPE port_cfg.axi_interface_type
`endif

`ifndef __SVDOC__
typedef class svt_axi_transaction_exception_list;
typedef class svt_axi_transaction_exception;
`endif
typedef class svt_axi_barrier_pair_transaction;

/*
`define SVT_AXI_COHERENT_READ \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == READNOSNOOP) || \
  (coherent_xact_type == READONCE) || \
  (coherent_xact_type == READSHARED) || \
  (coherent_xact_type == READCLEAN) || \
  (coherent_xact_type == READNOTSHAREDDIRTY) || \
  (coherent_xact_type == READUNIQUE) || \
  (coherent_xact_type == CLEANUNIQUE) || 
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == MAKEINVALID) || \
  (coherent_xact_type == DVMCOMPLETE) || \
  (coherent_xact_type == DVMMESSAGE) || \
  (coherent_xact_type == READBARRIER) \
)

`define SVT_AXI_COHERENT_WRITE \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == WRITENOSNOOP) || \
  (coherent_xact_type == WRITEUNIQUE) || \
  (coherent_xact_type == WRITELINEUNIQUE) || \
  (coherent_xact_type == WRITEBACK) || \
  (coherent_xact_type == WRITECLEAN) || \
  (coherent_xact_type == WRITEBARRIER) || \
  (coherent_xact_type == EVICT) || \
  (coherent_xact_type == WRITEEVICT) \
)
*/

// Transactions which always have 1 beat even if
// burst_length indicates cache line size.
`define SVT_AXI_COHERENT_READ_1_BEAT \
(xact_type == COHERENT) && \
( \
  (coherent_xact_type == CLEANUNIQUE) || \
  (coherent_xact_type == MAKEUNIQUE) || \
  (coherent_xact_type == CLEANSHARED) || \
  (coherent_xact_type == CLEANINVALID) || \
  (coherent_xact_type == CLEANSHAREDPERSIST) || \
  (coherent_xact_type == MAKEINVALID) \
)

`ifdef SVT_UVM_ENABLE_FGP
class svt_axi_thread_specific_svt_pattern_data;
    svt_pattern_data pttrn_contents[$];
    svt_pattern_data port_cfg_exists_pd;
endclass
`endif

/**
    This is the base transaction type which contains all the physical
    attributes of the transaction like address, data, burst type, burst length,
    etc. It also provides the timing information of the transaction to the
    master & slave transactors, that is, delays for valid and ready signals
    with respect to some reference events. 
    
    The svt_axi_transaction also contains a handle to configuration object of
    type #svt_axi_port_configuration, which provides the configuration of the
    port on which this transaction would be applied. The port configuration is
    used during randomizing the transaction.
 */
class svt_axi_transaction extends `SVT_TRANSACTION_TYPE;

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_typename(svt_axi_transaction)
`endif

  /**
    @grouphdr axi3_protocol AXI3 protocol attributes
    This group contains attributes which are relevant to AXI3 protocol.
    */

  /**
    @grouphdr axi4_protocol AXI4 protocol attributes
    This group contains attributes specific to AXI4 protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr axi3_4_delays AXI3 and AXI4 delay attributes
    This group contains attributes which can be used to control delays in AXI3 and AXI4 signals.
    */

  /**
    @grouphdr axi3_4_status AXI3 and AXI4 transaction status attributes
    This group contains attributes which report the status of AXI3 and AXI4 transaction.
    */

  /**
    @grouphdr axi3_4_ace_timing Timing and cycle information
    This group contains attributes which report the Timing and
    cycle information for Valid and Ready signals. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
   * @groupname axi5_protocol protocol attributes
    This group contains attributes which are relevant to AXI5 protocol.
    As of now read data chunking and unique id identifier is added.
   */

  /**
    @grouphdr out_of_order Out Of Order transaction attributes
    This group contains attributes used to generate out of order transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr interleaving Interleaved transaction attributes
    This group contains attributes used to generate interleaved transactions. These attributes are
    relevant to AXI3, AXI4 and ACE protocols.
    */

  /**
    @grouphdr ace_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE protocol. Please also refer to group @groupref axi3_protocol for AXI3 protocol attributes.
    */

  /**
    @grouphdr ace_delays ACE delay attributes
    This group contains members which can be used to control delays in ACE signals. Please also refer to group @groupref axi3_4_delays for AXI3 and AXI4 delay attributes.
    */

  /**
    @grouphdr ace_status ACE transaction status attributes
    This group contains attributes which report the status of ACE transaction. Please also refer to group @groupref axi3_4_status for AXI3 and AXI4 transaction status attributes.
    */

  /**
    @grouphdr ace_l3_cache ACE L3 Cache related attributes
    This group contains attributes which are relevant to L3 Cache usage under ACE protocol. This is applicable only when l3_cache_enable is set to '1' in system_configuration.
    */

  /**
    @grouphdr ace5_protocol ACE protocol attributes
    This group contains attributes which are relevant to ACE5 protocol.
    */

  /**
    @grouphdr axi4_stream_protocol AXI4 Stream protocol attributes
    This group contains attributes which represent AXI4 Stream protocol transaction fields.
    */

  /**
    @grouphdr axi4_stream_delays AXI4 Stream delay attributes
    This group contains attributes which can be used to control delays in AXI4 Stream signals.
    */

  /**
    @grouphdr axi_misc Miscellaneous attributes
    This group contains miscellaneous attributes which do not fall under any of the categories above.
    */
  // ****************************************************************************
  // Enumerated Types
  // ****************************************************************************

  /**
   * Enum to represent transfer sizes
   */
  typedef enum bit [3:0] {
    BURST_SIZE_8BIT    = `SVT_AXI_TRANSACTION_BURST_SIZE_8,
    BURST_SIZE_16BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_16,
    BURST_SIZE_32BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_32,
    BURST_SIZE_64BIT   = `SVT_AXI_TRANSACTION_BURST_SIZE_64,
    BURST_SIZE_128BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_128,
    BURST_SIZE_256BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_256,
    BURST_SIZE_512BIT  = `SVT_AXI_TRANSACTION_BURST_SIZE_512,
    BURST_SIZE_1024BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_1024,
    BURST_SIZE_2048BIT = `SVT_AXI_TRANSACTION_BURST_SIZE_2048
  } burst_size_enum;

  /**
   * Enum to represent burst type in a transaction
   */
  typedef enum bit[1:0]{
    FIXED = `SVT_AXI_TRANSACTION_BURST_FIXED,
    INCR =  `SVT_AXI_TRANSACTION_BURST_INCR,
    WRAP =  `SVT_AXI_TRANSACTION_BURST_WRAP
  } burst_type_enum;

  /**
   *  Enum to represent transaction type
   *  NOTE: IDLE value is currently reserved. Currently not used.
   *  Note: ATOMIC value is used for atomic transactions.
   *  Note: READ_WRITE value is used to represent transmitted_channel for ATOMICLOAD, ATOMICSWAP and ATOMICCOMPARE transactions.
   */
  typedef enum bit [2:0]{
    READ      = `SVT_AXI_TRANSACTION_TYPE_READ,
    WRITE     = `SVT_AXI_TRANSACTION_TYPE_WRITE,
    IDLE      = `SVT_AXI_TRANSACTION_TYPE_IDLE,
    COHERENT  = `SVT_AXI_TRANSACTION_TYPE_COHERENT,
    DATA_STREAM  = `SVT_AXI_TRANSACTION_DATA_STREAM
`ifdef SVT_ACE5_ENABLE
    ,ATOMIC   = `SVT_AXI_TRANSACTION_TYPE_ATOMIC,  /**<: ATOMICSTORE, ATOMICLOAD, ATOMICSWAP, ATOMICCOMPARE */
    READ_WRITE = `SVT_AXI_TRANSACTION_TYPE_READ_WRITE  
`endif
  } xact_type_enum;

  /**
   * Enum to represent phase type in a transaction
   */
  typedef enum bit [2:0]{
    WR_ADDR  = `SVT_AXI_PHASE_TYPE_WR_ADDR,
    WR_DATA  = `SVT_AXI_PHASE_TYPE_WR_DATA,
    WR_RESP  = `SVT_AXI_PHASE_TYPE_WR_RESP,
    RD_ADDR  = `SVT_AXI_PHASE_TYPE_RD_ADDR,
    RD_DATA  = `SVT_AXI_PHASE_TYPE_RD_DATA
  } phase_type_enum;

  /**
   * Enum to represent the coherent transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    READNOSNOOP          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOSNOOP,
    READONCE             = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCE,
    READSHARED           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READSHARED,
    READCLEAN            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READCLEAN,
    READNOTSHAREDDIRTY   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READNOTSHAREDDIRTY,
    READUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READUNIQUE,
    CLEANUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANUNIQUE,
    MAKEUNIQUE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEUNIQUE,
    CLEANSHARED          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHARED,
    CLEANINVALID         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANINVALID,
    MAKEINVALID          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_MAKEINVALID,
    DVMCOMPLETE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMCOMPLETE,
    DVMMESSAGE           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_DVMMESSAGE,
    READBARRIER          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READBARRIER,
    WRITENOSNOOP         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITENOSNOOP,
    WRITEUNIQUE          = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUE,
    WRITELINEUNIQUE      = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITELINEUNIQUE,
    WRITECLEAN           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITECLEAN,
    WRITEBACK            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBACK,
    EVICT                = `SVT_AXI_COHERENT_TRANSACTION_TYPE_EVICT,
    WRITEBARRIER         = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEBARRIER,
    WRITEEVICT           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEEVICT,
    CLEANSHAREDPERSIST   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CLEANSHAREDPERSIST,
    READONCECLEANINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCECLEANINVALID,
    READONCEMAKEINVALID = `SVT_AXI_COHERENT_TRANSACTION_TYPE_READONCEMAKEINVALID
    `ifdef SVT_AXI_CUSTNV_ENV
    , CUSTNV_L3PREFETCH   = `SVT_AXI_CUSTNV_L3PREFETCH
    `endif
`ifdef SVT_ACE5_ENABLE   
    ,WRITEUNIQUEPTLSTASH    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEPTLSTASH, 
    WRITEUNIQUEFULLSTASH   = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEUNIQUEFULLSTASH,
    STASHONCESHARED        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCESHARED,
    STASHONCEUNIQUE        = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHONCEUNIQUE,
    STASHTRANSLATION       = `SVT_AXI_COHERENT_TRANSACTION_TYPE_STASHTRANSLATION,
    CMO                    = `SVT_AXI_COHERENT_TRANSACTION_TYPE_CMO,
    WRITEPTLCMO            = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEPTL_CMO,
    WRITEFULLCMO           = `SVT_AXI_COHERENT_TRANSACTION_TYPE_WRITEFULL_CMO
`endif
  } coherent_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  typedef enum {
   CLEANINVALID_ON_WRITE = `SVT_AXI_CMO_CLEANINVALID_ON_WRITE,
   CLEANSHARED_ON_WRITE = `SVT_AXI_CMO_CLEANSHARED_ON_WRITE,
   CLEANSHAREDPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDPERSIST_ON_WRITE,
   CLEANSHAREDDEEPPERSIST_ON_WRITE = `SVT_AXI_CMO_CLEANSHAREDDEEPPERSIST_ON_WRITE
  } cmo_on_write_xact_type_enum;

typedef enum {
  WRITENOSNPFULL_CLEANSHARED = `SVT_AXI_WRITENOSNPFULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANINVALID = `SVT_AXI_WRITENOSNPFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHARED= `SVT_AXI_WRITENOSNPPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANINVALID= `SVT_AXI_WRITENOSNPPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITENOSNPPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEULL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEFULL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEFULL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHARED= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHARED_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANINVALID= `SVT_AXI_WRITEUNIQUEPTL_CLEANINVALID_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDPERSIST_WRITE_WITH_CMO_XACT_TYPE,
  WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST= `SVT_AXI_WRITEUNIQUEPTL_CLEANSHAREDDEEPPERSIST_WRITE_WITH_CMO_XACT_TYPE
  } write_with_cmo_xact_type_enum;
`endif

  typedef enum bit[2:0] {
    BYTE_STREAM = `SVT_AXI_STREAM_TYPE_BYTE_STREAM,
    CONTINUOUS_ALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_ALIGNED_STREAM,
    CONTINUOUS_UNALIGNED_STREAM = `SVT_AXI_STREAM_TYPE_CONTINUOUS_UNALIGNED_STREAM,
    SPARSE_STREAM = `SVT_AXI_STREAM_TYPE_SPARSE_STREAM,
    USER_STREAM = `SVT_AXI_STREAM_TYPE_USER_STREAM
  } stream_xact_type_enum;

`ifdef SVT_ACE5_ENABLE
  /** Defines the atomic transaction type */
  typedef enum bit[2:0]
    {
     NON_ATOMIC = `SVT_AXI_ATOMIC_TYPE_NON_ATOMIC,   /**<: Value that corresponds to non-atomic transaction type */
     STORE      = `SVT_AXI_ATOMIC_TYPE_STORE,     /**<: xact_type corresponds to one of the Atomic load operations */
     LOAD       = `SVT_AXI_ATOMIC_TYPE_LOAD,    /**<: xact_type corresponds to one of the Atomic store operations */
     SWAP       = `SVT_AXI_ATOMIC_TYPE_SWAP,     /**<: xact_type corresponds to Atomic swap operation */
     COMPARE    = `SVT_AXI_ATOMIC_TYPE_COMPARE   /**<: xact_type corresponds to the Atomic compare operation */
  } atomic_transaction_type_enum;

 typedef enum bit[4:0]
  {
   ATOMICSTORE_ADD        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_ADD,     /**<Atomic transactions AtomicStore Add */
   ATOMICSTORE_CLR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_CLR,     /**<Atomic transactions AtomicStore Clr */
   ATOMICSTORE_EOR        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_EOR,     /**<Atomic transactions AtomicStore Eor */
   ATOMICSTORE_SET        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SET,     /**<Atomic transactions AtomicStore Set */
   ATOMICSTORE_SMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMAX,    /**<Atomic transactions AtomicStore Smax */
   ATOMICSTORE_SMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_SMIN,    /**<Atomic transactions AtomicStore Smin */
   ATOMICSTORE_UMAX       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMAX,    /**<Atomic transactions AtomicStore Umax */
   ATOMICSTORE_UMIN       = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSTORE_UMIN,    /**<Atomic transactions AtomicStore Umin */
   ATOMICLOAD_ADD         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_ADD,      /**<Atomic transactions AtomicLoad Add */
   ATOMICLOAD_CLR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_CLR,      /**<Atomic transactions AtomicLoad Clr */
   ATOMICLOAD_EOR         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_EOR,      /**<Atomic transactions AtomicLoad Eor */
   ATOMICLOAD_SET         = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SET,      /**<Atomic transactions AtomicLoad Set */
   ATOMICLOAD_SMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMAX,     /**<Atomic transactions AtomicLoad Smax */
   ATOMICLOAD_SMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_SMIN,     /**<Atomic transactions AtomicLoad Smin */
   ATOMICLOAD_UMAX        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMAX,     /**<Atomic transactions AtomicLoad Umax */
   ATOMICLOAD_UMIN        = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICLOAD_UMIN,     /**<Atomic transactions AtomicLoad Umin */
   ATOMICSWAP             = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICSWAP,          /**<Atomic transactions AtomicSwap */
   ATOMICCOMPARE          = `SVT_AXI_ATOMIC_XACT_TYPE_ATOMICCOMPARE        /**<Atomic transactions AtomicCompare */ 

  } atomic_xact_op_type_enum;

  /** 
   * Enum to represent the Endianness of the outbound write data sent in Atomic transactions.
   * Following are the possible values:
   * - LITTLE_ENDIAN : Indicates that the outbound Atomic Write data is in the Little Endian format
   * - BIG_ENDIAN    : Indicates that the outbound Atomic Write data is in the Big Endian format
   * .
   */
  typedef enum {
    LITTLE_ENDIAN       =  0,
    BIG_ENDIAN          =  1
  } endian_enum;  

  /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DAT channel.
   * Following are the possible values:
   * - TAG_INVALID  : The tags are not valid.
   * - TAG_TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - TAG_UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - TAG_FETCH_MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory, in 
   * -                      reads the allocation tags will be fetched from memory for read transactions.
   * .
   */
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0]{
    TAG_INVALID  = 0,
    TAG_TRANSFER = 1,
    TAG_UPDATE   = 2,
    TAG_FETCH_MATCH = 3
  } tag_op_enum;


 
/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   *  This field will be populated by the VIP and must not be set by the users.
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
 
  typedef enum bit[(`SVT_AXI_TAGOP_WIDTH-1):0] {
     MATCH_NOT_PERFORMED = 0,
     NO_MATCH_RESULT  = 1,
     FAIL = 2,
     PASS = 3
  } tag_match_resp_enum;  

`endif
 /**
   * Enum to represent four levels of shareability domain for snoop
   * transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE. 
   */
  typedef enum bit [1:0] {
    NONSHAREABLE      = `SVT_AXI_DOMAIN_TYPE_NONSHAREABLE,
    INNERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_INNERSHAREABLE,
    OUTERSHAREABLE    = `SVT_AXI_DOMAIN_TYPE_OUTERSHAREABLE,
    SYSTEMSHAREABLE   = `SVT_AXI_DOMAIN_TYPE_SYSTEMSHAREABLE
  } xact_shareability_domain_enum;

  /**
   * Enum to represent barrier transaction type. Enum to represent four levels
   * of shareability domain for snoop transactions. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum bit [1:0] {
    NORMAL_ACCESS_RESPECT_BARRIER = `SVT_AXI_NORMAL_ACCESS_RESPECT_BARRIER,
    MEMORY_BARRIER                = `SVT_AXI_MEMORY_BARRIER,
    NORMAL_ACCESS_IGNORE_BARRIER  = `SVT_AXI_NORMAL_ACCESS_IGNORE_BARRIER,
    SYNC_BARRIER                  = `SVT_AXI_SYNC_BARRIER
  } barrier_type_enum;

  /**
   * Enum to represent responses for a coherent transaction Additional read
   * response bits that provide information on the completion of a shareable
   * read transaction.  Enum to represent barrier transaction type. Enum to
   * represent four levels of shareability domain for snoop transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */
  typedef enum  bit [1:0] {
    UNIQUE_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_CLEAN, 
    UNIQUE_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_UNIQUE_DIRTY,
    SHARED_CLEAN   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_CLEAN,
    SHARED_DIRTY   = `SVT_AXI_COHERENT_RESP_TYPE_SHARED_DIRTY
  } coherent_resp_type_enum;

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [1:0] {
    NORMAL     = `SVT_AXI_TRANSACTION_NORMAL,
    EXCLUSIVE  = `SVT_AXI_TRANSACTION_EXCLUSIVE,
    LOCKED     = `SVT_AXI_TRANSACTION_LOCKED
  } atomic_type_enum;

  /**
   * Enum to represent the status of coherent exclusive access
   */
  typedef enum {
    EXCL_ACCESS_INITIAL  = `SVT_AXI_COHERENT_EXCL_ACCESS_INITIAL,
    EXCL_ACCESS_PASS     = `SVT_AXI_COHERENT_EXCL_ACCESS_PASS,
    EXCL_ACCESS_FAIL     = `SVT_AXI_COHERENT_EXCL_ACCESS_FAIL 
  } excl_access_status_enum;

  /** 
   * Enum to represent the status of master exclusive monitor, which indicates the cause of failure for a coherent exclusive store
   */ 
  typedef enum {
    EXCL_MON_INVALID  = `SVT_AXI_EXCL_MON_INVALID,
    EXCL_MON_SET      = `SVT_AXI_EXCL_MON_SET,
    EXCL_MON_RESET    = `SVT_AXI_EXCL_MON_RESET
  } excl_mon_status_enum;  

  /**
   * Enum to represent locked type in a transaction
   */

  typedef enum bit [2:0] {
    DATA_SECURE_NORMAL                = `SVT_AXI_DATA_SECURE_NORMAL,               
    DATA_SECURE_PRIVILEGED            = `SVT_AXI_DATA_SECURE_PRIVILEGED,               
    DATA_NON_SECURE_NORMAL            = `SVT_AXI_DATA_NON_SECURE_NORMAL,               
    DATA_NON_SECURE_PRIVILEGED        = `SVT_AXI_DATA_NON_SECURE_PRIVILEGED,           
    INSTRUCTION_SECURE_NORMAL         = `SVT_AXI_INSTRUCTION_SECURE_NORMAL,            
    INSTRUCTION_SECURE_PRIVILEGED     = `SVT_AXI_INSTRUCTION_SECURE_PRIVILEGED,         
    INSTRUCTION_NON_SECURE_NORMAL     = `SVT_AXI_INSTRUCTION_NON_SECURE_NORMAL,        
    INSTRUCTION_NON_SECURE_PRIVILEGED = `SVT_AXI_INSTRUCTION_NON_SECURE_PRIVILEGED    
  } prot_type_enum;

  /**
   * Enum to represent responses in a transaction
   */
  typedef enum bit [1:0] {
    OKAY    = `SVT_AXI_OKAY_RESPONSE,
    EXOKAY  = `SVT_AXI_EXOKAY_RESPONSE,
    SLVERR = `SVT_AXI_SLVERR_RESPONSE,
    DECERR  = `SVT_AXI_DECERR_RESPONSE
  } resp_type_enum;

  typedef enum bit [2:0] {
    INVALID = `SVT_AXI_CACHE_LINE_STATE_INVALID,
    UNIQUECLEAN = `SVT_AXI_CACHE_LINE_STATE_UNIQUECLEAN,
    SHAREDCLEAN = `SVT_AXI_CACHE_LINE_STATE_SHAREDCLEAN,
    UNIQUEDIRTY = `SVT_AXI_CACHE_LINE_STATE_UNIQUEDIRTY,
    SHAREDDIRTY = `SVT_AXI_CACHE_LINE_STATE_SHAREDDIRTY
  } cache_line_state_enum;
 
  /**
   * Enum to represent DVM Message type.
   *
   * The bit representation of this type matches the encoding of the DVM message type field
   * in the AxADDR AMBA4 signal.
   * 
   * Used in the svt_amba_pv_extension class.
   */
  typedef enum bit [2:0] {
    TLB_INVALIDATE                        = 'h0, /**< TLB invalidate */
    BRANCH_PREDICTOR_INVALIDATE           = 'h1, /**< Branch predictor invalidate */
    PHYSICAL_INSTRUCTION_CACHE_INVALIDATE = 'h2, /**< Physical instruction cache invalidate */
    VIRTUAL_INSTRUCTION_CACHE_INVALIDATE  = 'h3, /**< Virtual instruction cache invalidate */
    SYNC                                  = 'h4, /**< Synchronisation message */
    HINT                                  = 'h6  /**< Reserved message type for future Hint messages */
  } dvm_message_enum;

  /**
   * Enum to represent DVM message Guest OS or hypervisor type.
   *
   * The bit representation of this type matches the encoding of the DVM guest OS or 
   * hypervisor field in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    HYPERVISOR_OR_GUEST = 'h0, /**< Transaction applies to hypervisor and all Guest OS*/
    GUEST               = 'h2, /**< Transaction applies to Guest OS */
    HYPERVISOR          = 'h3  /**< Transaction applies to hypervisor */
  } dvm_os_enum;

  /**
   * Enum to represent DVM message security type.
   *
   * The bit representation of this type matches the encoding of the DVM security field
   * in the AxADDR AMBA4 signal.
   */
  typedef enum bit [1:0] {
    AMBA_PV_SECURE_AND_NON_SECURE = 'h0, /**< Transaction applies to Secure and Non-secure */
    AMBA_PV_SECURE_ONLY           = 'h2, /**< Transaction applies to Secure only */
    AMBA_PV_NON_SECURE_ONLY       = 'h3  /**< Transaction applies to Non-secure only */
  } dvm_security_enum;


  /**
   *  Enum for interleave block pattern
   */

  typedef enum {
    EQUAL_BLOCK   = `SVT_AXI_TRANSACTION_INTERLEAVE_EQUAL_BLOCK,
    RANDOM_BLOCK  = `SVT_AXI_TRANASCTION_INTERLEAVE_RANDOM_BLOCK
  } interleave_pattern_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    PREV_ADDR_VALID      =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_VALID_REF,
    PREV_ADDR_HANDSHAKE  =  `SVT_AXI_MASTER_TRANSACTION_PREV_ADDR_HANDSHAKE_REF,
    FIRST_WVALID_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_WVALID_DATA_BEFORE_ADDR,
    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR = `SVT_AXI_MASTER_TRANSACTION_FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR,
    PREV_LAST_DATA_HANDSHAKE = `SVT_AXI_MASTER_TRANSACTION_PREV_LAST_DATA_HANDSHAKE
  } reference_event_for_addr_valid_delay_enum;

  /** 
   *  Enum to represent data delay reference event
   */
  typedef enum {
    WRITE_ADDR_VALID                           = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_VALID_REF,    
    //removed address handshake refrence because  of potential deadlock due to following reason::
    //the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    WRITE_ADDR_HANDSHAKE                       = `SVT_AXI_MASTER_TRANSACTION_WRITE_ADDR_HANDSHAKE_REF,
    PREV_WRITE_DATA_HANDSHAKE                  = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_DATA_HANDSHAKE_REF
  }  reference_event_for_first_wvalid_delay_enum;

  typedef enum {
    PREV_WVALID            = `SVT_AXI_MASTER_TRANSACTION_PREV_WVALID_REF,
    PREV_WRITE_HANDSHAKE   = `SVT_AXI_MASTER_TRANSACTION_PREV_WRITE_HANDSHAKE_REF
  } reference_event_for_next_wvalid_delay_enum;
  
  /** 
   *  Enum to represent tvalid delay reference event
   */
  typedef enum {
    PREV_TVALID_TREADY_HANDSHAKE          = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_TREADY_HANDSHAKE_REF,
    PREV_TVALID                           = `SVT_AXI_MASTER_TRANSACTION_PREV_TVALID_REF
  }  reference_event_for_tvalid_delay_enum;

  typedef enum {
    RVALID               = `SVT_AXI_MASTER_TRANSACTION_RVALID_REF,                                 
    MANUAL_RREADY        = `SVT_AXI_MASTER_TRANSACTION_MANUAL_RREADY_REF       
  } reference_event_for_rready_delay_enum;

  /** 
   *  Enum to represent response delay reference event
   */
  typedef enum {
    BVALID               =   `SVT_AXI_MASTER_TRANSACTION_BVALID_REF
  } reference_event_for_bready_delay_enum;
 
  /** 
   * Enum to represent read acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    LAST_READ_DATA_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_LAST_READ_DATA_HANDSHAKE_REF
  } reference_event_for_rack_delay_enum;
  
  /** 
   * Enum to represent write acknowledgment delay reference event. Applicable
   * when svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  typedef enum {
    WRITE_RESP_HANDSHAKE    = `SVT_AXI_MASTER_TRANSACTION_WRITE_RESP_HANDSHAKE_REF
  } reference_event_for_wack_delay_enum;

  /** 
   *  Enum to represent address delay reference event
   */
  typedef enum {
    ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_ADDR_VALID_REF,
    FIRST_WVALID            = `SVT_AXI_SLAVE_TRANSACTION_FIRST_WVALID_REF
  } reference_event_for_addr_ready_delay_enum;

  /** 
   *  Enum to represent reference event for delay for first rvalid
   */
  typedef enum {
    READ_ADDR_VALID               = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_VALID_REF,    
    READ_ADDR_HANDSHAKE           = `SVT_AXI_SLAVE_TRANSACTION_READ_ADDR_HANDSHAKE_REF
  }  reference_event_for_first_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for second rvalid onwards
   */
  typedef enum {
    PREV_RVALID          = `SVT_AXI_SLAVE_TRANSACTION_PREV_RVALID_REF,
    PREV_READ_HANDSHAKE  = `SVT_AXI_SLAVE_TRANSACTION_PREV_READ_HANDSHAKE_REF
  } reference_event_for_next_rvalid_delay_enum;

  /** 
   *  Enum to represent reference event for delay for wready signal
   */
  typedef enum {
    WVALID               = `SVT_AXI_SLAVE_TRANSACTION_WVALID_REF,                                 
    MANUAL_WREADY        = `SVT_AXI_SLAVE_TRANSACTION_MANUAL_WREADY_REF       
  } reference_event_for_wready_delay_enum;

  /** 
   *  Enum to represent write response delay reference event
   */
  typedef enum {
    LAST_DATA_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_LAST_DATA_HANDSHAKE_REF,
    ADDR_HANDSHAKE = `SVT_AXI_SLAVE_TRANSACTION_ADDR_HANDSHAKE_REF
  } reference_event_for_bvalid_delay_enum;

 
    
   // ****************************************************************************
   // Public Data
   // ****************************************************************************
   /** @groupname axi_misc
     * Variable that holds the object_id of this transaction
     */
   int object_id = -1;
   /** @groupname axi_misc
    * Variables used in generating XML/FSDB for pa writer 
    */
   
   string pa_object_type = "";
   string pa_channel_name ="" ;
   string bus_parent_uid = "";
   string bus_activity_type_name;

   /** @groupname axi_misc
     * The port configuration corresponding to this transaction
     */
   svt_axi_port_configuration port_cfg;
   
   /** 
    * @groupname ace_protocol
    * This member points to a barrier pair transaction
    * associated to this current transaction.  When associated_barrier_xact is
    * null, it indicates that this current transaction is not a post-barrier
    * transaction.  When associated_barrier_xact is non-null, this current
    * transaction will wait for responses from the barrier transactions in
    * associated_barrier_xact, before it can be transmitted.
    *
    * associated_barrier_xact can be set in the callback
    * svt_axi_master_callback::associate_xact_to_barrier_pair. In this
    * callback, user can associate this transaction with a barrier transaction
    * pair.
    *
    * Please refer to User Guide for more details on usage of this member.
    */
   svt_axi_barrier_pair_transaction  associated_barrier_xact;

`ifdef SVT_UVM_TECHNOLOGY
   /**
     * @groupname axi_misc 
     * Applicable only for master in ACTIVE mode.
     * If this transaction was generated from a UVM TLM Generic Payload, this
     * member indicates the GP from which this AXI transaction was generated
     */
   uvm_tlm_generic_payload causal_gp_xact;
`endif

  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------
  /** @cond PRIVATE */
  /** 
    * Object used to hold exceptions for a packet. 
    */
  `ifndef __SVDOC__
  svt_axi_transaction_exception_list exception_list = null; 
  `endif
 /** W riter used in callbacks to generate output for pa or verdi */ 
  protected svt_xml_writer xml_writer = null ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_mask ;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  addr_range;

  protected rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0]  burst_addr_mask ;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_width. Calculated in pre_randomize */

  //protected bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_possible_addr;

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /**
    * Used in system monitor to indicate if all bytes of a slave transaction
    * has been correlated to a corresponding master transaction
    */
  bit  is_slave_xact_correlated = 0;
  
  /**
    * Used in port monitor to indicate resize and aligned data status
    * in data_before_addr transaction.
    */
  bit  is_resize_and_align_data = 0;


  /** 
    * Indicates if data read from memory for a given beat contains X
    * The slave driver uses this information to decide whether to 
    * drive X on data.
    */
  bit read_data_contains_x[];

  /** The maximum possible address based on addr_user_width. Calculated in pre_randomize */
  // protected bit [`SVT_AXI_MAX_ADDR_USER_WIDTH-1:0] max_possible_user_addr;

  /** @endcond */

  /**
   * @groupname axi3_protocol
   * The variable holds the value of  AWID/WID/BID/ARID/RID signals.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ID_WIDTH. Default value of this macro is 8. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ID_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::id_width.
   */
  rand bit [`SVT_AXI_MAX_ID_WIDTH - 1:0] id = 0;

  /**
   * @groupname axi3_protocol
   * The variable represents AWADDR when xact_type is WRITE and  ARADDR when
   * xact_type is READ.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_ADDR_WIDTH. Default value of this macro is 64. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_ADDR_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::addr_width.
   */
  rand bit [`SVT_AXI_MAX_ADDR_WIDTH - 1 : 0] addr = 0;
  
  /**
   * @groupname axi3_protocol
   * Represents the minimum byte address of this transaction. 
   * If tagging is enabled, this will be the minimum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the maximum byte address of this transaction. 
   * If tagging is enabled, this will be the maximum tagged address 
   *  .
   */
  rand bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_byte_addr =0;
  
  /**
   * @groupname axi3_protocol
   * Represents the total byte count of this transaction. 
   *  .
   */
  rand int total_byte_count = 0;
  
  /**
   *  @groupname axi3_protocol
   *  The variable represents the actual length of the burst. For eg.
   *  burst_length = 1 means a burst of length 1.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI3, burst length
   *  of 1 to 16 is supported.
   *
   *  If #svt_axi_port_configuration::axi_interface_type is AXI4, burst length
   *  of 1 to 256 is supported.
   */ 
  rand bit [`SVT_AXI_MAX_BURST_LENGTH_WIDTH: 0] burst_length = 1;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst size of a transaction . The variable holds the value
   *  for AWSIZE/ARSIZE. 
   */
  rand burst_size_enum burst_size = BURST_SIZE_8BIT;

  /**
   *  @groupname axi3_protocol
   *  Represents the burst type of a transaction. The burst type holds the value
   *  for AWBURST/ARBURST. Following are the possible burst types: 
   *  - FIXED
   *  - INCR
   *  - WRAP
   *  .
   */
  rand burst_type_enum burst_type = INCR;

  /**
   * @groupname axi3_protocol
   * Represents the transaction type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * - COHERENT : Represents a COHERENT transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE and
   * COHERENT transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI_ACE.
   */
  rand xact_type_enum xact_type = WRITE;
  
  /**
   * @groupname axi3_protocol
   * Represents the phase type.
   * Following are the possible transaction types:
   * - WRITE    : Represent a WRITE transaction. 
   * - READ     : Represents a READ transaction.
   * .
   *
   * Please note that WRITE and READ transaction type is valid for
   * #svt_axi_port_configuration::axi_interface_type is AXI3/AXI4/AXI4_LITE 
   */
  phase_type_enum phase_type = WR_ADDR;

  /**
   * @groupname axi3_protocol
   * Represents the atomic access of a transaction.  The variable holds the
   * value for AWLOCK/ARLOCK. Following are the possible atomic types:
   * - NORMAL     
   * - EXCLUSIVE  
   * - LOCKED
   * .
   * Please note that atomic type LOCKED is not yet supported.
   */
  rand atomic_type_enum atomic_type = NORMAL;

`ifdef SVT_ACE5_ENABLE
  /**
   * Indicates the endianness of the Outbound Write Data in an Atomic transaction.
   */
  rand endian_enum endian = LITTLE_ENDIAN;
`endif

`ifdef SVT_ACE5_ENABLE
  /**
   * @groupname axi5_protocol
   * Represents the Unique ID indicator Feature.
   * The variable holds the value of AWIDUNQ/BIDUNQ/ARIDUNQ/RIDUNQ signals.<br>
   * The Variable is used to indicate that there are
   * no outstanding transactions going on with the same AWID/BID/ARID/RID respectively
   * and it will remain unique till the transaction is completed.
   * In order to use this feature, user need to pass the user defined macro
   * at compile time +define+SVT_ACE5_ENABLE.
   * Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_ACE5_ENABLE macro is only used to enable this feature and signals.
   * The Signals can be configured and enabled by VIP configuration using
   * parameter svt_axi_port_configuration::unique_id_enable.
   *
   * This functionality is not supported yet.
   */
  rand bit unique_id = 0;
`endif

  /**
   *  @groupname axi3_protocol
   *  Represents the cache support of a transaction. The variable holds the
   *  value for AWCACHE/ARCACHE.
   *
   *  Following values are supported in AXI3 mode:
   *
   *  - SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE            
   *  - SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY           
   *  - SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC                  
   *  - SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_RD_ONLY      
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_WR_ONLY       
   *  - SVT_AXI_3_CACHEABLE_WR_THRU_ALLOC_ON_BOTH_RD_WR    
   *  - SVT_AXI_3_CACHEABLE_WR_BACK_ALLOC_ON_BOTH_RD_WR    
   *  .
   *  
   *  Following values for ARCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_ARCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_ARCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE      
   *  .
   *
   *  Following values for AWCACHE are supported in AXI4 mode:
   *  - SVT_AXI_4_AWCACHE_DEVICE_NON_BUFFERABLE                  
   *  - SVT_AXI_4_AWCACHE_DEVICE_BUFFERABLE                     
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE    
   *  - SVT_AXI_4_AWCACHE_NORMAL_NON_CACHABLE_BUFFERABLE         
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_ALLOCATE           
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_WRITE_ALLOCATE          
   *  - SVT_AXI_4_AWCACHE_WRITE_THROUGH_READ_AND_WRITE_ALLOCATE 
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_NO_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_ALLOCATE                
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_WRITE_ALLOCATE             
   *  - SVT_AXI_4_AWCACHE_WRITE_BACK_READ_AND_WRITE_ALLOCATE    
   *  .
   */

  rand bit [`SVT_AXI_CACHE_WIDTH - 1:0] cache_type = 0;

  /**
   *  @groupname axi3_protocol
   *  Represents the protection support of a transaction. The variable holds the
   *  value for AWPROT/ARPROT. The conventions of the enumeration are:
   *
   *  - NORMAL/PRIVILEGED   : Normal/Priveleged access represented by AWPROT[0]/ARPROT[0]
   *  - SECURE / NON_SECURE : Secure/Non-Secure access represented by AWPROT[1]/ARPROT[1]
   *  - DATA / INSTRUCTION  : Data/Instruction access represented by AWPROT[2]/ARPROT[2]
   *  .
   *
   *  For the above conventions, following are the possible protection types:
   *  - DATA_SECURE_NORMAL                    
   *  - DATA_SECURE_PRIVILEGED                    
   *  - DATA_NON_SECURE_NORMAL                    
   *  - DATA_NON_SECURE_PRIVILEGED                
   *  - INSTRUCTION_SECURE_NORMAL                 
   *  - INSTRUCTION_SECURE_PRIVILEGED              
   *  - INSTRUCTION_NON_SECURE_NORMAL
   *  - INSTRUCTION_NON_SECURE_PRIVILEGED
   *  .
   */

  rand  prot_type_enum prot_type = DATA_SECURE_NORMAL;

  /**
   *  @groupname ace_protocol
   *  Applicable when
   *  svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.  
   *  Users  who need to bypass lookup of cache to determine valid 
   *  initial cache line states can set this property to 1.
   *  In order to randomize this property to 1, the user must switch off 
   *  svt_axi_master_transaction::reasonable_bypass_cache_lookup constraint.
   *  Setting this property will enable transactions to be sent out even
   *  if the initial cache state does not meet requirements set by ACE 
   *  protocol. Please note that coherency is not guaranteed when this 
   *  property is set
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand  bit bypass_cache_lookup = 1'b0;  


  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data[];
`endif

`ifdef SVT_ACE5_ENABLE

 /**
   * @groupname ace5_protocol
   * This variable represents the read data for the atomic load,swap and compare transactions.
   * This data will be driven by the slave on the read data channel.
   * APPLICABLE IN ALL MODES:
   * If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   * data must be stored right-justified by the user. The model will drive the
   * data on the correct lanes.  If svt_axi_port_configuration::wysiwyg_enable
   * is set to 1, the data is  transmitted as programmed by user and is
   * reported as seen on bus. No right-justification is used in this case.<br>
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_DATA_WIDTH. Default value of this macro is 1024. To change the
   * maximum width of this variable, user can change the value of this macro.
   * Define the new value for the macro in file svt_axi_user_defines.svi, and
   * then specify this file to be compiled by the simulator. Also, specify
   * +define+SVT_AXI_INCLUDE_USER_DEFINES on the simulator compilation command
   * line. Please consult User Guide for additional information, and consult VIP
   * example for usage demonstration.<br>
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_data[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the Memory Tag value in the transaction driven on the data channel for transactions.
  * Every 4 bits of Tag correspond to one 16 byte chunk of data.
  * MASTER in active mode:
  *
  * For write transactions this variable specifies tags to be driven on the
  * WTAG bus. 
  * 
  * SLAVE in active mode:
  *
  * For read transactions this variable specifies tags to be driven on the
  * RTAG bus.
  *
  * PASSIVE MODE:
  * This variable stores the tags as seen on WTAG or RTAG bus.
  *
  *
  */
`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`else
  rand bit [`SVT_AXI_MAX_TAG_WIDTH - 1:0] tag[];
`endif

//---------------------------------------------------------------------------------------------

/**
  * @groupname ace5_protocol
  * This field defines the WTAGUPDATE value in the transaction.
  * Only applicable when the Tag value is passed in the transaction and the tagop field in 
  * the transaction is set to Update.
  * Each WTAGUPDATE bit corresponds to 4 bits of WTAG
  */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`else
  rand bit [`SVT_AXI_MAX_TAGUPDATE_WIDTH - 1:0] tag_update[];
`endif

/**
  * @groupname ace5_protocol
  * This field defines the BCOMP value in the transaction.
  * Indicates whether write transaction is observable at the completer endused for persistent CMOs on Write channel.
  * This is used to send the response to a tag Match operation.
  * This is also used for persistent CMOs on Write channel.
  */
 
 rand bit is_write_transaction_observable = 0;
//---------------------------------------------------------------------------------------------
 
 /** 
   * Enum to represent the operation to be performed on the tags present in the corresponding DATA channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
  rand tag_op_enum tag_op = TAG_INVALID ;

  /** 
   * Enum to represent the response sent by the completer on the corresponding Response channel.
   * Following are the possible values:
   * - INVALID  : The tags are not valid.
   * - TRANSFER : The tags are clean. Tag Match does not need to be performed.
   * - UPDATE   : The Allocation Tag values have been updated and are dirty. The tags in memory should be updated.
   * - MATCH    : The Physical Tags in the write must be checked against the Allocation Tag values obtained from memory.
   * .
   */
 rand tag_op_enum response_tag_op = TAG_INVALID;
 
//---------------------------------------------------------------------------------------------

/** 
   * Enum to represent the ‘Resp’ field in the TagMatch response.
   *  This field is only applicable for Write and Atomic transactions with TagOp in the request set to Match (TAG_FETCH_MATCH).
   * Following are the possible values:
   * - MATCH_NOT_PERFORMED  : The tag MATCH operation is not performed by the completer.
   * - NO_MATCH_RESULT  : The tag MATCH operation doesn't have a result.
   * - FAIL  : The tag MATCH operation is failed.
   * - PASS  : The tag MATCH operation is passed.
   * .
   */
   rand tag_match_resp_enum tag_match_resp = MATCH_NOT_PERFORMED ;

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This field defines the partition ID value in MPAM. This corresponds to AxMPAM[9:1] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PARTID_WIDTH - 1:0] mpam_partid;

 /**
   * @groupname ace5_protocol
   * This field defines the Perfromance Monitor Group (PMG) value in MPAM. This corresponds to AxMPAM[10] attribute.
   */
  rand bit [`SVT_AXI_MAX_MPAM_PERFMONGROUP_WIDTH - 1:0] mpam_perfmongroup;

 /**
   * @groupname ace5_protocol
   * This field defines the MPAM_NS value in MPAM. This corresponds to AxMPAM[0] attribute.
   */
  rand bit [`SVT_AXI_MPAM_NS_WIDTH - 1:0] mpam_ns;
//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the data that will be stored in the memory for atomic transactions 
   * after the atomic operation is performed.
   * APPLICABLE IN ALL MODES:
   * The SVT_AXI_MAX_DATA_WIDTH macro is only used to control the maximum width
   * of the signal. The actual width used by VIP is controlled by configuration
   * parameter svt_axi_port_configuration::data_width.
   */
`ifdef SVT_MEM_LOGIC_DATA
  logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`else
  bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_resultant_data[];
`endif


//---------------------------------------------------------------------------------------------

 /**
   * @groupname ace5_protocol
   * This variable represents the swap data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   * 
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_swap_data[];
`endif

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare data value for the atomic compare transactions.
   * This will not be programmed by the user.This is an internal variable and is populated by the AXI SLAVE.
   */

`ifdef SVT_MEM_LOGIC_DATA
  rand logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`else
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_compare_data[];
`endif

`endif

  /**
   * @groupname axi3_protocol
   * MASTER in active mode:
   *
   * For write transactions this variable specifies write data to be driven on the
   * WDATA bus. 
   * 
   * SLAVE in active mode:
   *
   * For read transactions this variable specifies read data to be driven on the
   * RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the write or read data as seen on WDATA or RDATA bus.
   *
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] physical_data[];
`endif

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable is only applicable for atomic transactions.
   * MASTER in active mode:
   * For Atomic LOAD , SWAP and COMPARE transactions specifies read data as seen on the RDATA bus. 
   * 
   * SLAVE in active mode:
   * This variable represents the read data for the atomic load,swap and compare transactions to be driven on the RDATA bus.
   *
   * PASSIVE MODE:
   * This variable stores the read data as seen on RDATA bus.
   *
   */

`ifdef SVT_MEM_LOGIC_DATA
   logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`else
   bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] atomic_read_physical_data[];
`endif

`endif

  /** @cond PRIVATE */
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string data_str = "";

`ifdef SVT_ACE5_ENABLE
  /**
    * The data array in string format. Used by psdisplay_short
    */
  local string atomic_read_data_str = "";
`endif

  /**
    * The wstrb array in string format. Used by psdisplay_short
    */
  local string wstrb_str = "";

  /**
    * The read response array in string format. Used by psdisplay_short
    */
  local string rresp_str = "";

  /**
    * The write response in string format. Used by psdisplay_short
    */
  local string bresp_str = "";

  /**
    * The valid_assertion_time in string format. Used by psdisplay_short
    */
  local string valid_assertion_time = "";
  
  /**
    * The ready_assertion_time in string format. Used by psdisplay_short
    */
  local string ready_assertion_time = "";
  
 /* holds transactions that attempt to access same cacheline at the same time current transaction

   * does and started before current transaction started */
  bit overlapped_xact_started_before[svt_axi_transaction];

  /* holds transactions that attempt to access same cacheline at the same time current transaction
   * does and started after current transaction started */
  bit overlapped_xact_started_after[svt_axi_transaction];
  
  /* Indicates xact complets with out_of_order*/
  bit is_xact_completed_out_of_order = 0;

  /* indicates how many transactions blocked progress of current transaction */
  int num_xacts_blocked_progress_of_curr_xact = 0;

  /* semaphore to access num_xacts_blocked_progress_of_curr_xact */
  semaphore sema_num_xacts_blocked_progress_of_curr_xact = new(1);
  /** @endcond */

  
  /**
   *  @groupname axi3_protocol
   *  Array of Write strobes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  wstrb must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the wstrb is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] wstrb[];

`ifdef SVT_ACE5_ENABLE
 
//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the swap write strobes  value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   * 
   */
  rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_swap_wstrb[];

//---------------------------------------------------------------------------------------------
 /**
   * @groupname ace5_protocol
   * This variable represents the compare write strobes value for the atomic compare transactions.
   * This must not be programmed by the user.This is an internal variable populated by the AXI SLAVE.
   */
   rand bit [`SVT_AXI_WSTRB_WIDTH - 1:0] atomic_compare_wstrb[];

`endif

  /**
   *  @groupname ace5_protocol
   *  Array of poison.It indicates the 
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] poison[];

`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname ace5_protocol
   *  Array of poisonal value driven by the active slave on the read data channel.
   *  This is onlyapplicable for Atomic LOad , Swap and compare transactions.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 0 (default), the
   *  poison must be stored right-justified by the user. The model will drive
   *  these strobes on the correct lanes.
   *  If svt_axi_port_configuration::wysiwyg_enable is set to 1, the poison is  
   *  transmitted as programmed by user and is reported as seen on bus. 
   *  No right-justification is used in this case.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH/64- 1:0] atomic_read_poison[];

`endif


  /**
   *  @groupname axi3_protocol
   *  This variable specifies the response for write transaction. The variable holds the
   *  value for BRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the write response received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The write response programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the write response seen on the bus.
   */

  rand resp_type_enum bresp = OKAY;

  /**
   *  @groupname axi3_protocol
   *  This array variable specifies the response for read transaction. The array holds the
   *  value for RRESP. Following are the possible response types:
   *  - OKAY    
   *  - EXOKAY  
   *  - SLVERR 
   *  - DECERR  
   *  .
   *          
   *  MASTER ACTIVE MODE:
   *
   *  Will Store the read responses received from the slave.
   *
   *  SLAVE ACTIVE MODE:
   *
   *  The read responses programmed by the user.
   *
   *  PASSIVE MODE - MASTER/SLAVE:
   *
   *  Stores the read responses seen on the bus.
   */

  rand resp_type_enum rresp[];

`ifndef SVT_AXI_MULTI_SIM_OVERLAP_ADDR_ISSUE 
  /** 
    * @groupname axi3_protocol
    * If set, the driver checks if this transaction accesses a location
    * addressed by a previous transaction from this port or from some other
    * master. If there are any such previous transactions, this transaction is
    * blocked until all those transactions complete.  Also, the driver does not
    * pull any more transactions until this transaction is unblocked.  If not set,
    * this transaction is not checked for access to a location which was
    * previously accessed by another transaction.  Applicable only when
    * svt_axi_system_configuration::overlap_addr_access_control_enable is set 
    *
    * Applicable for ACTIVE MASTER only
    */ 
  rand bit check_addr_overlap = 1'b0;

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * Suspends a master transaction until this bit is reset. This is checked
    * immediately after a transaction is pulled by the driver from the sequencer
    * after the post_input_port_get callback is issued by the driver. When set,
    * the driver does not pull any more transactions from the
    * sequencer/generator until the bit is reset
    *
    * Applicable for ACTIVE MASTER only
    */
  bit suspend_master_xact = 1'b0;
  /** @endcond */
   
`endif

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * This bit is set by master if a cache line is reserved for the transaction. 
    * Thie field is used by task which unreserves the cache line at the end of 
    * transaction to filtering. This is to ensure only command that reserved 
    * cache line should unreserve cache line.  
    *  
    * Applicable for ACTIVE MASTER only
    */
  bit is_cacheline_reserved = 1'b0;
  /** @endcond */

  /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend response/data
    * for a READ/WRITE/COHERENT transaction until this bit is reset. 
    * This bit is usually set by the testbench when it needs to provide
    * response information to the driver (the slave driver expects the response
    * information in 0 time), but the data to respond with is
    * not yet known.  The testbench can set this bit and put this transaction 
    * back into the input channel of the slave. 
    * The transaction's response/data will not be sent until this bit is reset. 
    * Once the data is available, the testbench can populate response fields 
    * and reset this bit, upon which the slave driver will send the 
    * response/data of this transaction.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_response = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend awready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_awready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_awready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend arready signal 
    * for a READ transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_arready is set to 0
    * svt_axi_transaction::addr_ready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_arready = 0;

 /**
    * @groupname axi3_protocol
    * A bit that indicates that the testbench would like to suspend wready signal 
    * for a WRITE transaction until this bit is reset. 
    * This is applicable only when svt_axi_port_configuration::default_wready is set to 0
    * svt_axi_transaction::wready_delay won't be applicable when this bit is set to 1
    *
    * Applicable for ACTIVE SLAVE only.
    */
  bit suspend_wready = 0;

  /**
    * @groupname ace_protocol
    * Represents the value of AWUNIQUE signal driven/sampled on the interface.
    * Applicable when svt_axi_port_configuration::awunique_enable is set.
    * AWUNIQUE is asserted as per table C3-9 of section C3.1.4 on AWUNIQUE
    * signal. The value in the randomized transaction may be overridden by the
    * driver as per protocol requirements. For transactions where AWUNIQUE may
    * be asserted or deasserted, the randomized value is driven.  
    */
  rand bit is_unique = 0;

  /**
   *  @groupname axi3_4_status
   *  Represents the current status of the read or write address.  Following are the
   *  possible status types.

   * - INITIAL               : Address phase has not yet started on the channel
   * - ACTIVE                : Address valid is asserted but ready is not 
   * - ACCEPT                : Address phase is complete 
   * - ABORTED               : Current transaction is aborted
   * .
   */

  status_enum addr_status = INITIAL;

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum data_status = INITIAL;

`ifdef SVT_ACE5_ENABLE
/**
   *  @groupname axi3_4_status
   *  Represents the status of the read or write data transfer.  Following are
   *  the possible status types.

   *  - INITIAL               : Data has not yet started on the channel
   *  - ACTIVE                : Data valid is asserted but ready is not asserted for the
   *                            current data beat. The current beat is indicated
   *                            by #current_data_beat_num variable
   *  - PARTIAL_ACCEPT        : The current data beat is completed but the next
   *                            data-beat is not started. The next data beat is
   *                            indicated by #current_data_beat_num
   *  - ACCEPT                : Data phase is complete 
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */

  status_enum atomic_read_data_status = INITIAL;
`endif

  /**
   *  @groupname axi3_4_status
   *  Represents the status of the write response transfer.  Following are
   *  the possible status types.
   *  - INITIAL               : Response has not yet started on the channel
   *  - ACTIVE                : BVALID is asserted, but not BREADY
   *  - ACCEPT                : Write response is complete
   *  - ABORTED               : Current transaction is aborted 
   *  .
   */


  status_enum write_resp_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of the read/write acknowledge sent via RACK/WACK for
   * ACE interface. RACK/WACK is asserted for a single cycle.
   * Following are  the possible status types:
   * - INITIAL               : RACK/WACK has not be asserted
   * - ACTIVE                : RACK/WACK is asserted
   * - ACCEPT                : RACK/WACK assertion is completed
   * - ABORTED               : Current transaction is aborted
   * .
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE.
   */

  status_enum ack_status = INITIAL;

  /**
   * @groupname ace_status
   * Represents the status of coherent exclusive access.
   * Following are  the possible status types: 
   * - EXCL_ACCESS_INITIAL   : Initial state of the transaction before it is processed by master 
   * - EXCL_ACCESS_PASS      : ACE exclusive access is successful
   * - EXCL_ACCESS_FAIL      : ACE exclusive access is failed
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description. 
   */
  excl_access_status_enum  excl_access_status = EXCL_ACCESS_INITIAL;
  

  /**
   * @groupname ace_status
   * Represents the status of master exclusive monitor, which indicates the
   * cause of failure for a coherent exclusive store.  It is valid only for
   * exclusive store transaction, that is, CleanUnique. For all other
   * transactions it is set to EXCL_MON_INVALID by default.
   * Following are  the possible status types:
   * - EXCL_MON_INVALID      : Master exclusive monitor does not monitor the exclusive access on the cache line associated with the transaction
   * - EXCL_MON_SET          : Master exclusive monitor is set for exclusive access on the cache line associated with the transaction
   * - EXCL_MON_RESET        : Master exclusive monitor is reset for exclusive access on the cache line associated with the transaction
   * .
   *
   * A combination of #excl_access_status and #excl_mon_status can be used to
   * determine the reason for failure of exclusive store. Please refer to the
   * User Guide for more description.
   */ 
  excl_mon_status_enum   excl_mon_status = EXCL_MON_INVALID;


  /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  current_data_beat_num = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_status
   *    This is a counter which is incremented for every beat. Useful when user
   *    would try to access the transaction class to know its current state.
   *    This represents the beat number for which the status is reflected in
   *    member data_status.
   */
  int  atomic_read_current_data_beat_num = 0;
`endif
  /**
   *  @groupname interleaving
   *  Represents the various interleave pattern for a read and write transaction.
   *  The interleave_pattern gives flexibility to program interleave blocks with
   *  different patterns as mentioned below.
   *
   *  A Block is group of beats within a transaction.
   *
   *  EQUAL_BLOCK         : Drives equal distribution of blocks provided by
   *                        #equal_block_length variable. 
   *
   *  RANDOM_BLOCK        : Drives the blocks programmed in random_interleave_array
   *
   * Please note that currently interleaving based on EQUAL_BLOCK is not
   * supported.
   */
  rand interleave_pattern_enum interleave_pattern = RANDOM_BLOCK;

  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  If the interleave_pattern is set to EQUAL_BLOCK then this variable 
   *  is used to define the block length.
   *  Please note that currently interleaving based on EQUAL_BLOCK is not
   *  supported.
   */

  rand int equal_block_length = 0;

  /** @endcond */

  /**
   *  @groupname interleaving
   *  When the interleave_pattern is set to RANDOM_BLOCK, the user would
   *  program this array with blocks. There are default constraints, which the
   *  user can override and set their own block patterns.
   */
  rand int random_interleave_array[];


  /** @cond PRIVATE */
  /**
   *  @groupname interleaving
   *  This variable will start a new interleave from the current transaction and
   *  informs the model to complete all the transactions prior to this
   *  transaction.
   *
   *  Example 1:
   *  Interleave depth = 2
   * 
   *  Requirement : 
   *  1) Interleave transaction 1- 10 with each other
   *  2) Interleave transactions 11 - 20 with each other
   *
   *  Solution :
   *  1) Program start_new_interleave=0 for transactions 1 - 10 
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Example 2:
   *  Interleave depth = 2
   *
   *  Requirement :
   *  1) Do not Interleave transactions 1 - 10
   *  2) Start Interleaving from transactions 11 - 20
   *
   *  Solution :
   *  1) Program start_new_interleave=1 for transactions 1-10
   *  2) Program start_new_interleave=1 for transaction 11
   *
   *  Please note that this parameter is not currently supported.
   */
  rand bit start_new_interleave = 0;
  /** @endcond */

  /**
   * @groupname interleaving , out_of_order
   * This variable controls enabling of interleaving for the current transaction.
   * 
   * Example:
   * svt_axi_port_configuration::read_data_reordering_depth = 2
   * 
   * Requirement:
   * Unless all beats of transaction 1 are sent out, the beats of 
   * 2nd transactions should not be sent.
   * 
   * Solution:
   * Program the enable_interleave = 0 for both the transaction 1.
   
   */
  rand bit enable_interleave = 0;
  
  /**
    * @groupname axi_protocol
    * When this bit is set , it indicates that this transaction has updated 
    * the AXI Slave memory with write data and other properties.
    */ 
  bit memory_update_complete_for_write =0;

`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * when this bit is set, it indicates that this transaction 
   * performed atomic operation and the result is stored in atomic_resultant_data.
   */
  bit is_atomic_resultant_data_calculated =0;
`endif 

  /**
   * @groupname ace_protocol
   * When this bit is set by user, it indicates that this transaction is
   * a post-barrier transaction and that it needs to wait for responses
   * from the barrier transaction pair indicated in #associated_barrier_xact.
   * #associated_barrier_xact can be set in the callback
   * svt_axi_master_callback::associate_xact_to_barrier_pair. In this callback,
   * user can associate this transaction with a barrier transaction pair.
   *
   * Please refer to User Guide for more description.
   */
  rand bit associate_barrier = 0;

  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions.
   *  In data_before_addr scenario (i.e., when data_before_addr = '1'), addr and data channel related delay considerations are: 
   *  1) For programming address_channel related delay: awvalid_delay and reference_event_for_addr_valid_delay are used.
   *   (for more information, look for the description of these variables).
   *    reference_event_for_addr_valid_delay should be set FIRST_WVALID_DATA_BEFORE_ADDR. 
   *    In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
   *    FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
   *    potential deadlock scenarios in SLAVE DUT where slave DUT waits for awvalid signal
   *    before driving wready signal.
   *  2) For programming data_channel related delay: wvalid_delay[] and reference_event_for_first_wvalid_delay & reference_event_for_next_wvalid_delay are used.
   *    (for more information, look for the description of these variables).
   *      For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
   *      For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
   *    In data_before_addr scenario, reference_event_for_first_wvalid_delay must be PREV_WRITE_DATA_HANDSHAKE, otherwise it will cause failure.
   *  .
   *    
   */
  rand bit data_before_addr = 0;
  
  /**
   *  @groupname axi3_protocol
   *  Indicates that data will start before address for write transactions,
   *  even though data_before_addr is set to 0. This is useful when
   *  awvalid is suspended for write transaction and respective transaction
   *  data is driven before resuming the suspended awvalid signal.
   */
  bit suspend_awvalid_to_data_before_addr = 0;

  /**
    * Indicates if the current data beat of a write transaction has wlast
    * asserted. This is useful when data is received before addr and it is
    * required to determine the last beat. This is a sticky bit  in that
    * it remains set to 1 after the last data beat.
    */ 
  bit is_last_write_data_beat = 0;

   // AXI 4 Variables

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWQOS/ARQOS 
   */
  rand bit[`SVT_AXI_QOS_WIDTH - 1:0] qos = 0;  
  

  /**
   *  @groupname axi4_protocol
   *  The variable holds the value for AWREGION/ARREGION
   */
  rand bit[`SVT_AXI_REGION_WIDTH - 1:0] region = 0;


  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals AWUSER/ARUSER.
   *  Applicable for all interface types. Enabled through port configuration
   *  parameters svt_axi_port_configuration::aruser_enable and
   *  svt_axi_port_configuration::awuser_enable.
   */
  rand bit[`SVT_AXI_MAX_ADDR_USER_WIDTH - 1:0] addr_user = 0;

  /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER. Applicable for all
   *  interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] data_user[];

`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname ace5_protocol
   *  The variable holds the value for signals RUSER.
   *  Applicable only if svt_axi_port_configuration::atomic_transactions_enable is set to1.
   *  Enabled through port configuration parameters
   *  svt_axi_port_configuration::ruser_enable.
   */
  rand bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] atomic_read_data_user[];
`endif

   /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signals WUSER/RUSER as they are driven on the bus
   *  Applicable for all interface types. Enabled through port configuration parameters
   *  svt_axi_port_configuration::wuser_enable and
   *  svt_axi_port_configuration::ruser_enable.
   */
   bit[`SVT_AXI_MAX_DATA_USER_WIDTH - 1:0] physical_data_user[];
 /**
   *  @groupname axi3_protocol
   *  The variable holds the value for signal BUSER. Applicable for all
   *  interface types. Enabled through port configuration parameter
   *  svt_axi_port_configuration::buser_enable.
   */
  rand bit[`SVT_AXI_MAX_BRESP_USER_WIDTH - 1:0] resp_user = 0;
  
  /** 
   * @groupname ace_protocol
   * This variable represents the shareability domain of coherent transactions.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI_ACE or ACE_LITE.
   */
  rand xact_shareability_domain_enum domain_type = NONSHAREABLE;

  /**
   * @groupname ace_protocol
   * This variable represents barrier transaction type. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand barrier_type_enum barrier_type = NORMAL_ACCESS_RESPECT_BARRIER;

  /** 
   * @groupname ace_protocol
   * This variable represents the shareable coherent transaction types. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
   */
  rand coherent_xact_type_enum coherent_xact_type = READNOSNOOP;

`ifdef SVT_ACE5_ENABLE
 /**
  * @groupname ace5_protocol 
  * This variable represents the cmo on the write channel.
  * Applicable when svt_axi_port_configuration::axi_interface_type is set to ACE_LITE.
  */
  rand cmo_on_write_xact_type_enum cmo_on_write_xact_type = CLEANSHARED_ON_WRITE;
`endif

  /** 
   * @groupname ace_protocol
   * Array for the coherent read responses. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   */
  rand coherent_resp_type_enum coh_rresp[];

  /**
    * @groupname ace_status
    * This variable represents the initial cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The initial cache line state of a transaction that is driven on
    * the READ channel is populated just after the reception of the first beat
    * of the response of a transaction.  The initial cache line state of a
    * transaction that is driven on the WRITE channel is populated just before
    * the transaction is started. This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum initial_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the prefinal cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The prefinal cache line state of a transaction is the state of the 
    * cache  just before cache is updated . This variable is updated by the VIP, and is a
    * read-only variable. User is not expected or supposed to modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum  prefinal_cache_line_state = INVALID;

   /*
    * @groupname ace_status
    * This variable represents the initial data in the cache. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE. For transactions driven on the READ channel, this field is 
    * populated just after the reception of the the first beat of the response
    * of the transaction.
    * For transactions driven on the WRITE channel, this is populated just
    * before the transaction is started.
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] initial_cache_line_data[];

  /**
    * @groupname ace_status
    * This variable represents the final cache line state. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or
    * ACE_LITE.  The final cache line state of a transaction is the state of the
    * the line just before the transaction ended. This variable is updated by
    * the VIP, and is a read-only variable. User is not expected or supposed to
    * modify this variable.
    *
    * Applicable for ACTIVE MASTER only.
    */
   cache_line_state_enum final_cache_line_state = INVALID;

  /**
    * @groupname ace_status
    * This variable represents the final cache line data. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * The final cache line data of a transaction is the data of the
    * the line just before the transaction ended. 
    *
    * Applicable for ACTIVE MASTER only.
    */
   bit[7:0] final_cache_line_data[];

  /**
   * @groupname ace_protocol
   * Indicates that the data as given in #cache_write_data in this transaction 
   * needs to be allocated in the cache. Applicable only when transaction type
   * is READUNIQUE or CLEANUNIQUE.
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Applicable for ACTIVE MASTER only.
   */
  rand bit allocate_in_cache;

  /**
   * @groupname ace_protocol
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Represents data that needs to be stored to the cache if the 
   * #allocate_in_cache bit is set for a READUNIQUE/CLEANUNIQUE transaction 
   * or if the transaction is MAKEUNIQUE.
   * Applicable to masters in active mode.
   * Refer section 3.6 of ACE specification.
   * Writes in ACE are performed by removing all other copies
   * of the cache line so that the master that is performing the write has
   * a unique copy at the time of writing. Depending on whether a paritial
   * or full update of a cache line is required a transaction such as
   * READUNIQUE,MAKEUNIQUE or CLEANUNIQUE is sent. Some of these transactions
   * such as READUNIQUE will return data (either from memory or the cache of
   * some other master) and this will be available in the data[] field of this
   * class. Other transactions such as MAKEUNIQUE and CLEANUNIQUE will not
   * return any data. 
   * For a READUNIQUE transaction, if the #allocate_in_cache bit is not set, the
   * data available in data[] is written in cache. If the #allocate_in_cache bit
   * is set the data available in this variable is written to cache. Note however,
   * that this variable is overwritten by the data that is received in data[] prior
   * to writing in the cache. This is done because READUNIQUE is used for partial update 
   * of a cacheline when a master does not have a copy of the cacheline. So a user 
   * can actually populate this variable after a copy of this cacheline is received and 
   * not at the time of randomization.
   * For a CLEANUNIQUE transaction, if the #allocate_in_cache bit is set,
   * the data in this variable is written to cache. 
   * For a MAKEUNIQUE transaction, the data in this variable is always written into
   * the cache.
   * Updating this variable is normally done in the pre_cache_update callback issued 
   * by the master driver after all the responses are received but prior to the 
   * RACK signal being driven.
   * An important aspect of this variable is that this data is not driven
   * on the physical bus.
   * 
   * Applicable for ACTIVE MASTER only.
   */
  rand bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] cache_write_data[];

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if update of cache must be bypassed for this transaction. A
    * typical use model is to set this bit in pre_cache_update callback of the
    * driver based on response received in the transaction. For example, if the
    * response received is SLVERR, user may not want the driver to update the
    * cache.  When using this property, it is the user's responsibility that
    * system coherency is not lost, since cache will not be updated.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit bypass_cache_update = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction ended because the requested data was already
    * available in the cache. This bit is set by the master, no action is taken
    * if the user sets this bit. A transaction with this bit set was not sent out
    * on the bus and therefore other components in the testbench will not detect
    * this transaction. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_cached_data = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
    *
    * Indicates if a coherent transaction was dropped because the start state
    * of the corresponding cache line is not as expected before transmitting the
    * transaction. The expected start states for each of the transaction types
    * are given in section 5 of the ACE specification.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_coherent_xact_dropped = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is a result of a speculative read operation.
    * A speculative read is defined as a read of a cache line that a master already
    * holds in its cache.
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is a speculative read. Modifying the value of this member will
    * not have any effect.
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_speculative_read = 0;

  /** @cond PRIVATE */
  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates whether the memory update at slave end for overlapped write
    * transactions should happen in request order.
    *
    * This is a read-only member, which VIP uses to update slave memory for 
    * overlapped write transactions. It should not be modified by the user.
    * 
    * Applicable for ACTIVE SLAVE only.
    */
  bit update_mem_in_req_order = 0;  

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for WriteUnique and WriteLineUnique
    * not being in progress while a WRITEBACK/WRITECLEAN is in progress is done
    * Applicable when port_interleaving_enable is set in the configuration.
    */
  bit is_wu_wlu_restriction_check_done = 0;

  /**
    * @groupname ace_protocol
    * Indicates whether the required checks for memory update transaction 
    * relative to the cache states are performed just prior to start
    * of this transaction
    */
  bit is_mem_update_pre_xact_xmit_check_done = 0;
  /** @endcond */

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    *
    * Indicates if the transaction is auto generated by the VIP. Transactions
    * are auto-generated when:
    * 1. The cache is full and an entry needs to be evicted from the cache. 
    * 2. User supplies a cache maintenance transaction and the protocol requires
    * that the cache line is first written into memory before sending the cache
    * maintenance transaction. 
    *
    * This is a read-only member, which VIP uses to indicate whether the
    * transaction is auto generated. It should not be modified by the user. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  bit is_auto_generated = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set
    * to AXI_ACE and svt_axi_port_configuration::snoop_response_data_transfer_mode 
    * is set to SNOOP_RESP_DATA_TRANSFER_USING_WB_WC.
    *
    * Indicates if this transaction is a WRITEBACK/WRITECLEAN auto-generated transaction
    * which was generated to transfer snoop data. When 
    * svt_axi_port_configuration::snoop_response_data_transfer_mode is set to 
    * SNOOP_RESP_DATA_TRANSFER_USING_WB_WC, snoop data from a dirty line is transferred
    * using a WRITEBACK/WRITECLEAN transaction instead of the snoop data channel. All
    * transactions which have this variable set will also have  is_auto_generated set.
    */
  bit is_xact_for_snoop_data_transfer = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to a shared state even
    * if the actual state of the line is unique, since it is permissible for
    * a cache line which is in the unique state to be held in the shared state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITH_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE or
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_shared_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE or ACE_LITE.
    * Indicates if the cache line state needs to be forced to an invalid state even
    * if that is not the recommended state, since it is permissible for
    * a cache line which is in a clean state to be held in the invalid state. 
    * Valid only when:
    * svt_axi_port_configuration::cache_line_state_change_type is set to
    * LEGAL_WITHOUT_SNOOP_FILTER_CACHE_LINE_STATE_CHANGE.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_to_invalid_state = 0;

  /**
    * @groupname ace_protocol
    * Applicable when svt_axi_port_configuration::axi_interface_type is set to
    * AXI_ACE or ACE_LITE.  Forces transactions which are not constrained to be
    * of cacheline size by protocol to be of cacheline size. Currently
    * applicable only to READONCE, WRITEUNIQUE, WRITENOSNOOP and READNOSNOOP
    * transactions. Applicable to WRITENOSNOOP and READNOSNOOP only when
    * svt_axi_port_configuration::update_cache_for_non_coherent_xacts is set and
    * svt_axi_port_configuration::axi_interface_type is AXI_ACE.
    * If this bit is set, READONCE and WRITEUNIQUE transactions will be forced
    * to cache line size transactions.
    * This has a dependency on svt_axi_port_configuration::force_xact_to_cache_line_size_interface_type. 
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand bit force_xact_to_cache_line_size = 0;
  
  /**
   * @groupname ace_protocol
   * The variable represents ARVMIDEXT when svt_axi_port_configuration::axi_interface_type 
   * is set to AXI_ACE or ACE_LITE with svt_axi_system_configuration::DVMV8_1 or above.
   * The maximum width of this signal is controlled through macro
   * SVT_AXI_MAX_VMIDEXT_WIDTH. Default value of this macro is 4 based on DVMv8.1 architecture recomendation.
   * 
   */

  rand bit [`SVT_AXI_MAX_VMIDEXT_WIDTH - 1:0] arvmid = 0;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit is_datachk_parity_error = 0;
`ifdef SVT_ACE5_ENABLE
 /**
   * @groupname ace5_protocol
   * This variable stores the data check parity bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_datachk_parity_value[] ;

  /**
   * @groupname ace5_protocol
   * This variable stores the data check parity error bit's with respect to valid data,
   * Each bit of parity check data is calculated from every 8bit of data with 1bit if datachk.
   * By default all bits are set to 'b1, if any parity error is detected the that particular bit is set to 0.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] atomic_read_is_datachk_passed[] ;

  /**
   * @groupname ace5_protocol
   * This variable represents the data check parity error is deducted in a
   * transaction.
   * In a transaction if parity error is deducted, the this bit is set to 1.
   * Applicable when svt_axi_port_configuration::check_type is set to ODD_PARITY_BYTE_DATA.
   */
  rand bit atomic_read_is_datachk_parity_error = 0;

  /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_transaction_type_enum atomic_transaction_type = NON_ATOMIC;

 /**
  * - @groupname ace5_protocol
  * - Field that indicates type of write_with_cmo_xact_type.
  * .
  */

  rand write_with_cmo_xact_type_enum write_with_cmo_xact_type = WRITENOSNPFULL_CLEANSHARED; 

 /**
   * - @groupname ace5_protocol 
   * - Field that indicates type of Atomic transaction.
   * - This is a read-only field for the testbench, and is set by the VIP components
   * .
   */
  rand atomic_xact_op_type_enum atomic_xact_op_type = ATOMICSTORE_ADD;

`endif
 /**
   * @groupname ace5_protocol 
   *This field indicates the value of trace_tag
   */
  rand bit trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of data trace_tag on write data channel and read data channel
   */
  rand bit data_trace_tag =0;

  /**
   * @groupname ace5_protocol
   * This field indicates the value of btrace on write response channel
   */
  rand bit resp_trace_tag =0;

`ifdef SVT_ACE5_ENABLE 
  /** Internal field to store the atomic data trace_tag for inbound data */
  rand bit atomic_read_data_trace_tag;

 /** 
   * @groupname ace5_protocol
   * This field indicates the node ID of the stash target. 
   * Applicable only in stash type transactions.
   */
  rand bit[(`SVT_AXI_STASH_NID_WIDTH-1):0] stash_nid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates the stash_nid field has a valid Stash target value.
   * Applicable only in stash type transactions.
   */
  rand bit stash_nid_valid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  indicates the ID of the logical processor at the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit [(`SVT_AXI_STASH_LPID_WIDTH-1):0] stash_lpid = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the Stash_lpid field value must be 
   * considered as the Stash target.
   * Applicable only in stash type transactions.
   */
  rand bit stash_lpid_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates the ID of the stream.This si used to identify the stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit [(`SVT_AXI_MAX_MMUSID_WIDTH-1):0] stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates wether the stream is secure or non-secure.
   * When set to 1, indicates a secure stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit secure_or_non_secure_stream = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field  is only vaid if sub_stream_id_valid is set to 1.
   * This indicates the ID of the sub stream.
   * Applicable only when untranslated transaction feature is supported.
   */
  rand bit[(`SVT_AXI_MAX_MMUSSID_WIDTH-1):0] sub_stream_id = 0;
  
  /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has an optional substream identifier.
   * When set to 1 , it means that transaction has a substream identifier.
   * This is used in untranslated transaction feature is enabled.
   */
  rand bit sub_stream_id_valid = 0;

 /** 
   * @groupname ace5_protocol
   * This field indicates that the transaction has already undergone PCIE ATS 
   * translation.
   */
  rand bit addr_translated_from_pcie = 0;

`endif

  /**
   *  Represents port ID. Not currently supported.
   */
  int port_id;

  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the cycle information for address valid on read and
   *   write transactions. The simulation clock cycle number when the address
   *   valid is asserted, is captured in this member. This information can be
   *   used for doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */
  int addr_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_valid_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for data valid on read and
   *  write transactions. The simulation clock cycle number when the data
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_valid_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response valid on a write
   *  transaction. The simulation clock cycle number when the write response
   *  valid is asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */
  int write_resp_valid_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation clock cycle number when the address valid
   *  and ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */
  int addr_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int data_ready_assertion_cycle[];
`ifdef SVT_ACE5_ENABLE
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation clock cycle number when the data valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int atomic_read_data_ready_assertion_cycle[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for response ready on a write
   *  transaction. The simulation clock cycle number when the write response valid and
   *  ready both are asserted, is captured in this member. This information can be
   *  used for doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  int write_resp_ready_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *   The simulation time when the master or slave driver receives
   *   the transaction from the sequencer, is captured in this member.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  realtime xact_consumed_by_driver_time;
 /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the cycle information for address wakeup of read or write 
   *  transaction. The simulation clock cycle number when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  int addr_wakeup_assertion_cycle;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address wakeup of read or write
   *  transaction. The simulation time when the address wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real addr_wakeup_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
  real idle_chan_wakeup_toggle_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for wakeup of idle read or write
   *  channel. The simulation time when the wakeup is
   *  deasserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member variable,
   *  user does not need to program this variable.
   */
   real idle_chan_wakeup_toggle_deassertion_time;

 /**
   *   @groupname axi3_4_ace_timing
   *   This variable stores the transaction consumed at driver timing
   *   information. The transaction consumed at driver time to begin time
   *   delay is calculated as the difference between begin_time and
   *   xact_consumed_by_driver_time.
   *   This information can be used for doing performance analysis.
   *   VIP updates the value of this member variable,
   *   user does not need to program this variable.
   */

  real xact_consumed_time_to_begin_time_delay;
  
  /**
   *  @groupname axi3_4_ace_timing
   *   This variable stores the timing information for address valid on read and
   *   write transactions. The simulation time when the address valid is
   *   asserted, is captured in this member. This information can be used for
   *   doing performance analysis. VIP updates the value of this member
   *   variable, user does not need to program this variable.
   */

  real addr_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_valid_assertion_time[];
`ifdef SVT_ACE5_ENABLE
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data valid on read and
   *  write transactions. The simulation time when the data valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_valid_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response valid on  write
   *  transactions. The simulation time when the response valid is
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real write_resp_valid_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for address ready on read and
   *  write transactions. The simulation time number when the address valid and
   *  ready both are asserted i.e. handshake happens, is captured in this member.
   *  This information can be used for doing performance analysis. VIP updates the
   *  value of this member variable, user does not need to program this variable.
   */

  realtime addr_ready_assertion_time;


  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real data_ready_assertion_time[];
`ifdef SVT_ACE5_ENABLE
   /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for data ready on read and
   *  write transactions. The simulation time when the data valid and ready both are
   *  asserted, is captured in this member. This information can be used for
   *  doing performance analysis. VIP updates the value of this member
   *  variable, user does not need to program this variable.
   */

  real atomic_read_data_ready_assertion_time[];
`endif
  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for response ready on  write
   *  transactions. The simulation time when the response valid and ready both are
   *  asserted, is captured in this member. This information can be used for doing
   *  performance analysis. VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */

  real write_resp_ready_assertion_time;

  /**
   *  @groupname axi3_4_ace_timing
   *  This variable stores the timing information for the data channnel blocking ratio.
   *  The blocking cycle for a beat is defined as the number of cycles that
   *  valid was asserted, but corresponding ready was not asserted.
   *  This ratio is derived from data_valid_assertion_cycle and
   *  data_ready_assertion_cycle, calculated as sum of data ready
   *  blocking cycles divided by sum of data valid assertion cycles.
   *  This information can be used for doing performance analysis.
   *  VIP updates the value of this member variable, user
   *  does not need to program this variable.
   */
  real data_chan_blocking_ratio;

  // ****************************************************************************
  // Members relevant to Master Driver and Monitor  
  // ****************************************************************************

  /**
    * @groupname axi3_4_delays
    * This variable defines the number of cycles the AWVALID or ARVALID  signal is
    * delayed. The reference event for this delay is #reference_event_for_addr_valid_delay.
    * Applicable for ACTIVE MASTER only.
    */
  rand int addr_valid_delay = 0;
   
  /**
    * @groupname axi3_4_delays
    * Defines a reference event from which the AWVALID or ARVALID delay
    * should start.  Following are the different reference events:
    *
    * PREV_ADDR_VALID:  
    * Reference event is the previous AWVALID or ARVALID signal 
    *
    * PREV_ADDR_HANDSHAKE:  
    * Reference event is previous read or write Address handshake
    *
    * FIRST_WVALID_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first wvalid of the current transaction.
    *
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR:
    * This is used when #data_before_addr bit is set. The reference event for
    * address valid to occur is the first data handshake of the current transaction.
    *
    * PREV_LAST_DATA_HANDSHAKE:
    * Reference event is previous read or write last data handshake
    * to Address valid assertion.
    *
    * Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios is added in svt_axi_transaction class 
    * to constraint the value of reference_event_for_addr_delay not to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * User may swicth off the constraint reasonable_reference_event_for_addr_delay by setting rand_mode to 0 
    * incase they want reasonable_reference_event_for_addr_delay to take FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR.
    * In data_before_addr scenarios reference_event_for_addr_delay should be set very carefully to
    * FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
    * potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
    * before driving wready signal.
    *
    */
  rand reference_event_for_addr_valid_delay_enum  reference_event_for_addr_valid_delay = PREV_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal assertion
    * before or after ARVALID or AWVALID signal.
    */
  rand int awakeup_assert_delay = 0;
  
  /**
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for AWAKEUP signal deassertion
    * after ARVALID-ARREADY or AWVALID-AWREADY signal handshake.
    */
  rand int awakeup_deassert_delay = 0;

  /** if this bit is set to '0' then AWAKEUP signal will be asserted 
    * before ARVALID with respect to awakeup_assert_delay.
    * if this bit is set to '1' then AWAKEUP signal will be asserted
    * after ARVALID or AWVALID with respect to awakeup_assert_delay.
    */ 
  rand bit assert_awakeup_after_valid = 0;

  /** 
    * @groupname axi3_4_delays
    * Defines the delay in number of cycles for WVALID signal.
    * The reference event for this delay is:
    * - For wvalid_delay[0]        -  #reference_event_for_first_wvalid_delay
    * - For remaining indices of wvalid_delay -  #reference_event_for_next_wvalid_delay
    * .
    * Applicable for ACTIVE MASTER only.
    */
  rand int wvalid_delay[];
   
  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * FALSE, this member defines the RREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_rready_delay
    *
    * If configuration parameter #svt_axi_port_configuration::default_rready is
    * TRUE, this member defines the number of clock cycles for which RREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int rready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which RREADY should be high and low
    * when the read data channel is idle, that is, when RVALID is low. This
    * property helps to toggle the RREADY signal during the idle period between
    * the assertion of RVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all read data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the read_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transaction unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until RVALID is asserted. When RVALID is observed on the interface,
    * this delay is no longer applicable. The delay specified in
    * #rready_delay is applied before this property is used.  Note that toggling
    * RREADY during the idle period may lead to situations where the RREADY
    * signal is already asserted when the RVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_rready is low. Similarly,
    * RREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_rready is high. In both
    * these cases, #rready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_rready_delay[];

  /**
   * @groupname axi4_stream_delays
   * Defines the delay in number of clock cycles for TVALID signal.
   * The reference event for this delay is:  #reference_event_for_tvalid_delay
   * - PREV_TVALID_TREADY_HANDSHAKE : Previous tvalid-tready handshake as the reference event
   * - PREV_TVALID                  : Previous tvalid assertion as the reference event
   * .
   * Applicable for ACTIVE MASTER only.
   */
  rand int tvalid_delay[];

  /**
   * @groupname axi4_stream_delays
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * FALSE, this member defines the TREADY signal delay in number of clock
   * cycles.  The reference event for this delay is
   * #reference_event_for_tready_delay.
   *
   * Please note that #reference_event_for_tready_delay is not supported
   * currently. Absolute value of tready_delay is considered for delay
   * calculation with respect to tvalid signal.
   *
   * If configuration parameter #svt_axi_port_configuration::default_tready is
   * TRUE, this member defines the number of clock cycles for which TREADY
   * signal should be deasserted after each handshake, before pulling it up
   * again to its default value.
   *
   * Applicable for ACTIVE SLAVE only.
   */
  rand int tready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first wvalid signal. The delay
    * must be programmed in wvalid_delay[0]. Following are the different
    * events under this category:
    *
    * WRITE_ADDR_VALID:
    * Reference event for first WVALID is assertion of AWVALID signal
    * 
    * WRITE_ADDR_HANDSHAKE:
    * This event is applicable when write data is transmitted after write
    * address, that is, when #data_before_addr is set to 0. This reference event
    * specifies the write address handshake.
    * 
    * PREV_WRITE_DATA_HANDSHAKE:
    * This event is applicable when write data is transmitted before write
    * address, that is, when #data_before_addr is set to 1. This reference event
    * specifies the previous write data handshake.
    */
    // removed address handshake refrence because  of potential deadlock due to following reason::
    // the slave can wait for AWVALID or WVALID, or both before asserting AWREADY
    //
  rand reference_event_for_first_wvalid_delay_enum reference_event_for_first_wvalid_delay =  WRITE_ADDR_VALID;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_WVALID:
    * Reference event for WVALID delay is assertion of previous wvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts wvalid.
    * 
    * PREV_WRITE_HANDSHAKE:
    * Reference event for WVALID delay is completion of previous data handshake.
    */
  rand reference_event_for_next_wvalid_delay_enum reference_event_for_next_wvalid_delay = PREV_WRITE_HANDSHAKE;

  /**
    *    
    * @groupname axi3_4_delays
    * Defines the reference event for RREADY delay.
    *   
    * RVALID:
    * Reference event for RREADY is assertion of RVALID signal
    * 
    * MANUAL_RREADY: (Not supported currently)
    *
    * This event  allows the user to generate  RREADY patterns, in cycles, as
    * follows:
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The rready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default rready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default rready signal is
    *       driven after toggling
    * 3. The remaining rready_delay element represents no. of cycles to drive
    *    rready
    * 
    * Example 1:
    * For eg.   RREADY  pattern (cycles) =  1110011 and default_rready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_rready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous RREADY value)

    * For eg. cycle pattern  RREADY =  0001100 and default_rready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_rready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous RREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous RREADY value)
    */
  rand reference_event_for_rready_delay_enum reference_event_for_rready_delay = RVALID;

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * FALSE, this member defines the BREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_bready_delay.
    * 
    * If configuration parameter #svt_axi_port_configuration::default_bready is
    * TRUE, this member defines the number of clock cycles for which BREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value.
    *
    * Applicable for ACTIVE MASTER only.
    */
  rand int bready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for master VIP.
    *
    * Indicates the number of cycles for which BREADY should be high and low
    * when the write response channel is idle, that is, when BVALID is low.
    * This property helps to toggle the BREADY signal during the idle period
    * between the assertion of BVALID signal.  The value for this property may
    * be set when the transaction is randomized at the master or in a callback
    * such as svt_axi_port_monitor_callback::write_resp_phase_started. Values
    * provided in even numbered indices indicate the number of clocks for which
    * the ready signal must be driven low and the values in odd numbered
    * indices indicate the number of clocks for which it must driven high.
    * Values in this variable are applicable only until BVALID is asserted.
    * When BVALID is observed on the interface, this delay is no longer
    * applicable. The delay specified in #bready_delay is applied before this
    * attribute is applied.  Note that toggling BREADY during the idle period
    * may lead to situations where the BREADY signal is already asserted when
    * BVALID is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is low. Similarly, BREADY may
    * be low when the corresponding valid is sampled, even though the value of
    * #svt_axi_port_configuration::default_bready is high. In both these cases,
    * #bready_delay is not applicable. The size of this array can be set to any
    * value greater than 0, based on the number of times the user would like
    * the signal to toggle during idle period.
    */
  rand int idle_bready_delay[];


  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BREADY delay.
    *
    * BVALID:
    * Reference event is assertion of BVALID signal
    */
  rand reference_event_for_bready_delay_enum reference_event_for_bready_delay = BVALID;

  /**
    * @groupname axi3_4_delays
    * This members applies to AWREADY signal delay for write transactions, and
    * ARREADY signal delay for read transactions.
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is FALSE, this member
    * defines the AWREADY or ARREADY signal delay in number of clock cycles.
    * The reference event used for this delay is
    * #reference_event_for_addr_ready_delay. 
    *
    * If configuration parameter #svt_axi_port_configuration::default_awready
    * or #svt_axi_port_configuration::default_arready is TRUE, this member
    * defines the number of clock cycles for which AWREADY or ARREADY signal
    * should be deasserted after each handshake, before pulling it up again to
    * its default value.
    *
    * Applicable for ACTIVE SLAVE only.
    */
  rand int addr_ready_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which awready and arready should be
    * high and low when the corresponding address channel is idle, that is,
    * when AWVALID/ARVALID is low. This property helps to toggle the
    * AWREADY/ARREADY signal during the idle period between the assertion of
    * AWVALID/ARVALID signal of this transaction and the next transaction.
    * This value may be assigned during randomization of the transaction object
    * in the slave sequence. Values provided in even numbered indices indicate
    * the number of clocks for which the ready signal must be driven low and
    * the values in odd numbered indices indicate the number of clocks for
    * which it must driven high. Values in this variable are applicable only
    * until the corresponding valid is asserted. When AWVALID/ARVALID is
    * observed on the interface, this delay is no longer applicable and the
    * delay specified in #addr_ready_delay is applied before asserting
    * AWREADY/ARREADY.  Note that toggling AWREADY/ARREADY during the idle
    * period may lead to situations where the AWREADY/ARREADY signal is already
    * asserted when the corresponding valid is sampled, even though the value
    * of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is low. Similarly,
    * AWREADY/ARREADY may be low when the corresponding valid is sampled, even
    * though the value of #svt_axi_port_configuration::default_awready or
    * #svt_axi_port_configuration::default_arready is high. In both these
    * cases, #addr_ready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_addr_ready_delay[];


  /** 
    * @groupname axi3_4_delays
    * Defines reference event for AWREADY or ARREADY delay.
    *
    * ADDR_VALID:
    * Reference event is  assertion of AWVALID or ARVALID signal. This event is
    * not applicable when default value of AWREADY = 1 or default value of
    * ARREADY = 1.
    * FIRST_WVALID:
    * Reference event is  assertion of WVALID signal. This event is
    * not applicable when default value of AWREADY = 1.
    * This event is only applicable for write address channel.
    */
  rand reference_event_for_addr_ready_delay_enum  reference_event_for_addr_ready_delay = ADDR_VALID;

  /** 
    * @groupname axi3_4_delays
    * Defines RVALID delay, in terms of number of clock cycles.
    * The reference event for this delay is:
    * - For rvalid_delay[0]        -  #reference_event_for_first_rvalid_delay
    * - For remaining indices of rvalid_delay -  #reference_event_for_next_rvalid_delay
    * .
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int rvalid_delay[];

  /**
    * @groupname axi3_4_delays
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * FALSE, this member defines the WREADY signal delay in number of clock
    * cycles.  The reference event for this delay is
    * #reference_event_for_wready_delay.
    *
    * If configuration parameter #svt_axi_port_configuration::default_wready is
    * TRUE, this member defines the number of clock cycles for which WREADY
    * signal should be deasserted after each handshake, before pulling it up
    * again to its default value. 
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Applicable when svt_axi_port_configuration::toggle_ready_signals_during_idle_period
    * is set. Applicable for slave VIP.
    *
    * Indicates the number of cycles for which wready should be high and low
    * when the write data channel is idle, that is, when WVALID is low. This
    * property helps to toggle the WREADY signal during the idle period between
    * the assertion of WVALID signal.  Values provided in even numbered indices
    * indicate the number of clocks for which the ready signal must be driven
    * low and the values in odd numbered indices indicate the number of clocks
    * for which it must driven high. Note that the values provided in this
    * variable are applied for all write data beats. If the user requires a
    * different set of delays during the idle period for each beat, the user
    * must use the write_data_phase_started callback to change the values of
    * this property for the corresponding beat. Once changed, the values will
    * be applicable for all subsequent beats of the transactions unless it is
    * is changed for a subsequent beat. Values in this variable are applicable
    * only until WVALID is asserted. When WVALID is observed on the interface,
    * this delay is no longer applicable and the delay specified in
    * #wready_delay is applied before asserting WREADY.  Note that toggling
    * WREADY during the idle period may lead to situations where the WREADY
    * signal is already asserted when the WVALID is sampled, even though the
    * value of #svt_axi_port_configuration::default_wready is low. Similarly,
    * WREADY may be low when the corresponding valid is sampled, even though
    * the value of #svt_axi_port_configuration::default_wready is high. In both
    * these cases, #wready_delay is not applicable. The size of this array can be
    * set to any value greater than 0, based on the number of times the user
    * would like the signal to toggle during idle period.
    */
  rand int idle_wready_delay[];

  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the first rvalid signal. The delay
    * must be programmed in rvalid_delay[0]. Following are the different
    * events under this category:
    *
    * READ_ADDR_VALID:
    * Reference event for first RVALID is assertion of ARVALID signal
    *
    * READ_ADDR_HANDSHAKE:
    * Reference event for first RVALID is completion of read address handshake
    */
  rand reference_event_for_first_rvalid_delay_enum reference_event_for_first_rvalid_delay = READ_ADDR_HANDSHAKE;


  /**
    * @groupname axi3_4_delays
    * Defines the reference events to delay the RVALID signals from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_RVALID :
    * Reference event to delay RVALID is assertion of previous rvalid.  The
    * delay timer starts as soon as previous valid signal is asserted. If
    * previous data handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts rvalid.
    * 
    * PREV_READ_HANDSHAKE :
    * Reference event to delay RVALID is completion of previous read data
    * handshake.
    */

  rand reference_event_for_next_rvalid_delay_enum reference_event_for_next_rvalid_delay = PREV_READ_HANDSHAKE;

  /**
    * @groupname axi3_4_delays
    * Defines the reference events for WREADY delay.
    *   
    * WVALID:
    * Reference event for WREADY is assertion of WVALID signal.
    * 
    * MANUAL_WREADY: (Not supported currently)
    * This event  allows the user to generate  WREADY patterns, in cycles, as
    * follows :
    * 1. The reference event for this delay is the beginning of the Address
    *    handshake.
    * 2. The wready_delay[0]  represents the following
    *    a. A value > 0 is the no. of cycles default wready signal is
    *       driven
    *    b. A value < 0 is the no. of cycles default wready signal is
    *       driven after toggling
    * 3. The remaining wready_delay element represents no. of cycles to drive
    *    wready
    * 
    * Example 1:
    * For eg.   WREADY  pattern (cycles) =  1110011 and default_wready = 1 
    * data_delay[0] = 3  Three cycles high (driving default_wready value) 
    * data_delay[1] = 2  Two cycles low    (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles high   (toggled previous WREADY value)

    * For eg. cycle pattern  WREADY =  0001100 and default_wready = 1 
    * data_delay[0] = -3 Three cycles low (toggled default_wready value) 
    * data_delay[1] = 2  Two cycles high  (toggled previous WREADY value) 
    * data_delay[2] = 2  Two cycles low   (toggled previous WREADY value)
    */

  rand reference_event_for_wready_delay_enum  reference_event_for_wready_delay =  WVALID;

  /**
    * @groupname axi3_4_delays
    * Defines the BVALID delay in terms of number of clock cycles. The reference
    * event for this delay is #reference_event_for_bvalid_delay.
    *
    * Applicable for ACTIVE SLAVE only.
    */

  rand int bvalid_delay = 0;

  /**
    * @groupname axi3_4_delays
    * Defines a reference event for BVALID delay.
    *
    * LAST_DATA_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for last write
    * data.
    * 
    * ADDR_HANDSHAKE:
    * Reference event for BVALID delay is completion of handshake for address phase.
    */  

  rand reference_event_for_bvalid_delay_enum reference_event_for_bvalid_delay = LAST_DATA_HANDSHAKE;

  /**
    * @groupname axi4_stream_delays
    * Defines the reference events for TVALID delay from second beat
    * onwards. Following are the different events under this category:
    *  
    * PREV_TVALID:
    * In this case, assertion of previous tvalid signal is considered  
    * as the reference event for TVALID delay. The delay timer
    * starts as soon as previous tvalid signal is asserted. If previous
    * tvalid-tready handshake does not complete before timer expires, the
    * current transfer waits for the previous handshake to complete, and then
    * immediately asserts tvalid.
    * 
    * PREV_TVALID_TREADY_HANDSHAKE:
    * Reference event for TVALID delay is completion of previous tvalid-tready handshake.
    */
  rand reference_event_for_tvalid_delay_enum reference_event_for_tvalid_delay = PREV_TVALID_TREADY_HANDSHAKE;

  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the RACK delay should start.
   * - LAST_READ_DATA_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_rack_delay_enum reference_event_for_rack_delay = LAST_READ_DATA_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the RACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_rack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int rack_delay = 0;
  
  /** 
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   *
   * Defines the reference event from which the WACK delay should start.
   * - WRITE_RESP_HANDSHAKE: Reference event is last data handshake
   * .
   */
  rand reference_event_for_wack_delay_enum reference_event_for_wack_delay = WRITE_RESP_HANDSHAKE;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the WACK delay in terms of number of clock cycles. The reference
   * event for this delay is #reference_event_for_wack_delay.
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int wack_delay = 0;

  /**
   * @groupname ace_delays
   * Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI_ACE.
   * Defines the delay between reception of DVM Sync and transmission of DVM Complete.
   * Delay for master component in terms of number of clock cycles for generating
   * DVM Complete transaction after receiving a DVM Sync transaction. 
   *
   * Applicable for ACTIVE MASTER only.
   */

  rand int dvm_complete_delay = 0;

  /**
   *  @groupname out_of_order
   *  Sets the reordering priority of the current transaction within the set
   *  of transactions that are allowed access to read data channel based on 
   *  svt_axi_port_configuration::read_data_reordering_depth.
   * 
   *  This member is applicable only when svt_axi_port_configuration::reordering_algorithm
   *  is svt_axi_port_configuration::PRIORITIZED.
   * 
   *  This value indicates the priority of sending the response to current 
   *  transaction compared to remaining transactions within the depth indicated
   *  by svt_axi_port_configuration::read_data_reordering_depth for read transactions or
   *  by svt_axi_port_configuration::write_resp_reordering_depth for write transactions.
   *
   *  Note that the value of this attribute should be within the following range:
   *  [1:svt_axi_port_configuration::read_data_reordering_depth] for read transactions and
   *  [1:svt_axi_port_configuration::write_resp_reordering_depth] for write transactions.
   * 
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘1’ then, the
   *  transactions with highest value for this attribute will get higher priority.
   *
   *  If svt_axi_port_configuration::reordering_priority_high_value is set to ‘0’ then, the
   *  transactions with least value for this attribute will get higher priority.
   *
   *  If there are more than one transactions with same priority, those transaction
   *  will be processed in the same order as they are received.
   * 
   * Applicable for ACTIVE SLAVE only.
   */

  rand int reordering_priority = 1;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of zero delay within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int ZERO_DELAY_wt = 100;

   /**
     * @groupname axi3_4_delays
     * Weight used to control distribution of short delays within transaction generation.
     *
     * This controls the distribution of delays for the 'delay' fields 
     * (e.g., delays for asserting the ready signals).
     */
  int SHORT_DELAY_wt = 500;

  /**
    * @groupname axi3_4_delays
    * Weight used to control distribution of long delays within transaction generation.
    *
    * This controls the distribution of delays for the 'delay' fields 
    * (e.g., delays for asserting the ready signals).
    */
  int LONG_DELAY_wt = 1;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of burst length to 1 within transaction
     * generation.
     *
     * This controls the distribution of the length of the bursts using
     * burst_length field 
     */
  int ZERO_BURST_wt = 100;

   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of short bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int SHORT_BURST_wt = 500;


   /**
     * @groupname axi3_protocol
     * Weight used to control distribution of longer bursts within transaction
     * generation.
     *
     * This controls the distribution of  the length of the bursts using
     * burst_length field 
     */
  int LONG_BURST_wt = 400;


  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

   /**
    * @groupname axi4_stream_protocol
    * Used to drive TDATA signals. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
   rand bit [`SVT_AXI_MAX_TDATA_WIDTH - 1:0] tdata[];

  
  /**
   * @groupname axi4_stream_protocol
   * Used to drive TSTRB signal. The strobes are right aligned and the model
   * will drive strobes on appropriate lanes. The model also takes care of the
   * endianness while driving tstrb. Applicable when
   * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TSTRB_WIDTH - 1:0] tstrb[];

 
  /**
   * @groupname axi4_stream_protocol
   * TKEEP is the byte qualifier that indicates whether the content of the
   * associated byte of TDATA is processed as part of the data stream.
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to
   * AXI4_STREAM.
   */
  rand bit [`SVT_AXI_TKEEP_WIDTH - 1:0] tkeep[];


  /**
    * @groupname axi4_stream_protocol
    * The variable holds the value of  TID signal. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand bit [`SVT_AXI_MAX_TID_WIDTH - 1:0] tid = 0;
  
  /**
    * @groupname axi4_stream_protocol
    * TDEST provides routing information for the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TDEST_WIDTH - 1:0] tdest;
  
  /**
    * @groupname axi4_stream_protocol
    * TUSER is user defined sideband information that can be transmitted
    * alongside the data stream. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */

  rand bit [`SVT_AXI_MAX_TUSER_WIDTH - 1:0] tuser[];

  /**
    * @groupname axi4_stream_protocol
    * Defines the burst length of a AXI4 Stream Packet. Applicable when
    * svt_axi_port_configuration::axi_interface_type is set to AXI4_STREAM.
    */
  rand int stream_burst_length = 1;

  // ****************************************************************************
  // End of STREAM SIGNALS
  // ****************************************************************************
  /**
    * @groupname axi3_protocol
    * A bit that must be set by the user to indicate that this transaction will
    * be sent to the slave driver from the slave sequencer through the
    * delayed_response_request_port of the slave driver. If the transaction is
    * randomized before putting it into the delayed_response_request_port of the
    * slave driver, then this bit must be set by the user. This bit must not be
    * set for a transaction that is sent on the seq_item_port.
    */
  bit is_delayed_response_xact = 0;

  /**
   * @groupname axi_misc
   * Indicates the value of the source master which will be propogated in the ID field
   * of the master and the corresponding slave transaction.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::source_master_id_xmit_to_slaves_type is set to
   * DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES. This property must be set by the
   * user in a system monitor callback issued at the start of a transaction
   */
  bit[`SVT_AXI_DYNAMIC_SOURCE_MASTER_ID_XMIT_TO_SLAVES_WIDTH-1:0] dynamic_source_master_id_xmit_to_slaves = 0;

  /**
   * @groupname axi_misc
   * Indicates that this master transaction is a partial write transaction and this
   * transaction will be split by the interconnect into a full Read transaction
   * followed by partial Write transaction to the corresponding slave.
   * Applicable for users who want to correlate master transactions to slave
   * transactions in the system monitor. This parameter is applicable when
   * svt_axi_port_configuration::partial_write_to_slave_read_and_write_association_enable is set to
   * This property must be set by the user in a system monitor callback issued at the start of a transaction
   */
  bit partial_master_write_split_into_read_modified_write_slave_xact = 0;

  /**
   * @groupname axi_misc
   * Multibit array for different usages.
   * 
	 * If cust_xact_flow[0] is set to '1', indicate that transaction should be drived immediately on the interface.
	 * This is aplicable only for AXI4 STREAM transactions.
	 *
	 * cust_xact_flow[31:1] bits are for future use.
   */
  rand bit[31:0] cust_xact_flow = 0;  

  /** @cond PRIVATE */
  /**
    * @groupname axi3_protocol
    * A bit that is set by the slave driver to indicate that the write response
    * of a transaction has been provided by the user through the
    * delayed_response_request_port of the slave driver.  
    * Applicable only when
    * svt_axi_port_configuration::enable_delayed_response_port is set.
    */
  bit is_delayed_write_response_set = 0;

  /** 
    * @groupname ace_l3_cache
    * Inidcates that current transaction will cause memory update transaction for the associated
    * cacheline if it is  hit in L3 and found to be in dirty state.
    */
  bit clean_l3_data = 0;

  /** 
    * @groupname ace_l3_cache
    * This attribute is supposed to be updated by VIP indicating to the user that memory has been
    * updated for the current transaction with associated cacheline data in L3 cache. This is primarily
    * used along with clean_l3_data i.e. if current transaction is expected to update memory then user
    * can wait for this attribute to be set by VIP if user needs to perform any tasks based on that condition.
    */
  bit mem_updated_with_l3_data = 0;
  /** @endcond */

  `ifdef SVT_ACE5_ENABLE  
  /**
    * @groupname axi5_protocol
    * Defines the chunk enable of a AXI5 to enable read_data_chunking. When enable, slave will send read data
    * in 128bits of chunk in random order. If disabled, slave will send read data without chunking as per AXI5 protocol. Applicable 
    * when svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit archunken = 0;

  /**
    * @groupname axi5_protocol
    * Array of read chunk strobe
    * Each bit of rchunkstrb represents 128bits of read data. Width of the rchunkstrb by default is 
    * `SVT_AXI_MAX_CHUNK_STROBE_WIDTH user can change width using svt_axi_port_configuration::rchunkstrb_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1 : 0] rchunkstrb[];

  /**
    * @groupname axi5_protocol
    * Array of read chunk number
    * Indicates that the data chunk number is being transferred. Width of the rchunknum by default is 
    * `SVT_AXI_MAX_CHUNK_NUM_WIDTH user can change width using svt_axi_port_configuration::rchunknum_width 
    * signal. Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable is set to 1.
    * Not yet implemented. 
    */
  rand bit [`SVT_AXI_MAX_CHUNK_NUM_WIDTH -1 : 0] rchunknum[];

  /**
    * @groupname axi5_protocol
    * Indicates that the data chunk length is being transferred. This signal is for interal use to calculate number  
    * of transafer for chunkinig Applicable when archunken and svt_axi_port_configuration::rdata_chunking_enable 
    * is set to 1.
    * Not yet implemented. 
    */
  rand int chunk_length;

  /**
   * @groupname axi5_protocol
   *    This is a counter which is incremented for every chunk of databeat. Useful when user
   *    would try to access the transaction class to know its current state during chunking.
   *    This represents the chunk databeat transfer number.
   */
  int  current_data_chunk_trf_num = 0;
  `endif  

  // ****************************************************************************
  // STREAM SIGNALS
  // ****************************************************************************

  `ifdef SVT_AXI_QVN_ENABLE
  /**
   * @groupname qvn_parameters
   * Applicable when svt_axi_port_configuration::axi_interface_type is set to AXI3/AXI4/ACE/ACE_LITE
   * Specifies the Virtual Network ID to which token for this transaction will be requested.
   * Same Virtual Network will be used to send current transaction as well. 
   *
   * Active Master will use qvn_vnet_id to determine which VN*VALID* signal needs to be asserted
   * to request for token and all ARVNET_ID or AWVNET_ID and WVNET_ID value will be driven
   * same as qvn_vnet_id
   *
   * Port Monitor will use qvn_vnet_id to indicate from which Virtual Network this particular 
   * transaction has been received.
   *
   */
  rand int qvn_vnet_id = 0;
  `endif

  `ifdef SVT_AXI_CUSTNV_ENV
  /** 
    * configuration register used to provide custom L3 or interconncet based behaviour
    * [0] = '1' indicates writeEvict can start from shared state.
    * [1] = '1' indicates no data has been provided as part of the read response.
    * [2] = '1' indicates current transaction is a block linear request.
    * [3] = '1' indicates current transaction is auto-generated by VIP for an origninal block linear request.
    *           this bit is supposed to get set by VIP. User doesn't need to set this bit.
    *
    * default value of all fields are 0 and it is set by user except bit[3].
    */
  bit[31:0] custnv_reg = 0;
  `endif
  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  local static vmm_log shared_log = new("svt_axi_transaction", "class" );
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
  local svt_axi_port_configuration::axi_port_kind_enum axi_port_kind = svt_axi_port_configuration::AXI_MASTER;

  local svt_axi_port_configuration::axi_interface_type_enum axi_interface_type = svt_axi_port_configuration::AXI3; 
`endif

  /** @cond PRIVATE */
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_data_width_in_bytes = 0;
  
  /** Helper attribute for randomization calculated during pre_randomize */
  protected int data_width_in_bytes = 0;
 
  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH/8 -1 :0] atomic_read_poison_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected bit[`SVT_AXI_MAX_DATA_WIDTH -1 :0] atomic_comp_read_data_mask =0;

  /** Helper attribute for randomization calculated during pre_randomize */
  protected int log_base_2_cache_line_size = 0;

  /** internal flag to track if transaction is part of a multi-part dvm sequence */

  bit is_part_of_multipart_dvm_sequence = 0;

  /** The channel (READ/WRITE) on which this transaction will be transmitted */
  xact_type_enum transmitted_channel = WRITE;

  /** The xact_type when port_cfg is_downstream_coherent = 1 */
  xact_type_enum converted_xact_type = WRITE; 
  /** @endcond */
 
  // ****************************************************************************
  // Local variables only for internal VIP usages
  // ****************************************************************************
  bit [(`CEIL(`SVT_AXI_MAX_ID_WIDTH,8))-1:0] axidchk_parity_value = 0;
  bit [(`CEIL(`SVT_AXI_MAX_ADDR_WIDTH,8))-1:0] axaddrchk_parity_value = 0;
  bit axlenchk_parity_value  = 0;
  bit axctlchk0_parity_value = 0;
  bit axctlchk1_parity_value = 0;
  bit axctlchk2_parity_value = 0;
  bit arctlchk3_parity_value = 0;
  bit [(`CEIL((`SVT_AXI_MAX_DATA_WIDTH/8),8))-1:0]       wstrbchk_parity_value;

  // ****************************************************************************
  // Constraints
  // ****************************************************************************

`protected
XWF4?O>f3A5,F:_?-WR51aQJ8McYR,VO(ZfH8aQG?=D\L?O9MB8^2)VL,:E6XE>_
UfVQ2-[93\I,-$
`endprotected

  
  /** Re-organised constraint blocks based on interface type. This will make
   * it easy to turn-off the constraints based on interface type. It can
   * result in significant run-time improvement. */

  // QVN Constraints Block. These constraints are valid when QVN mode is
  // enabled. 
  constraint qvn_valid_ranges {
`ifdef SVT_AXI_QVN_ENABLE
    solve xact_type before qvn_vnet_id;
    solve coherent_xact_type before qvn_vnet_id;

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
    if(port_cfg.qvn_enable) {
        // -------------------------------------------------------------------------------
        // Each Transaction should pick Virtual Network only from the list of supported VN
        // -------------------------------------------------------------------------------
        qvn_vnet_id inside {[0:`SVT_AXI_QVN_MAX_NUM_VIRTUAL_NETWORK-1]};

        if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) ) {
          foreach(port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_aw_chnl[ix]) -> qvn_vnet_id != ix;
          }
        } else {
          foreach(port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) {
            (!port_cfg.qvn_supported_virtual_network_queue_ar_chnl[ix]) -> qvn_vnet_id != ix;
          }
        }
        // -------------------------------------------------------------------------------
    }
    else {
       qvn_vnet_id == 0;
    }
`endif // SVT_AXI_SVC_NO_CFG_IN_XACT
`endif // SVT_AXI_QVN_ENABLE
  } // qvn_valid_ranges

// These constraints are applicable for Memory tagging feature
 constraint memory_tagging_valid_ranges {
`ifdef SVT_ACE5_ENABLE
 if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER){
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(transmitted_channel == WRITE || transmitted_channel == READ_WRITE) {
     if(port_cfg.mte_support_type == svt_axi_port_configuration::BASIC){
       !tag_op inside {TAG_TRANSFER,TAG_FETCH_MATCH};
       if(xact_type == ATOMIC){
         tag_op == TAG_INVALID;}
    if(xact_type == COHERENT)  {
      if(coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE}){
       tag_op  inside {TAG_INVALID,TAG_UPDATE}; }
      else if (coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
      tag_op ==TAG_INVALID;}
     }
   if(xact_type == WRITE){
     tag_op  inside {TAG_INVALID,TAG_UPDATE};}
   }
   if(port_cfg.mte_support_type == svt_axi_port_configuration::STANDARD){
     tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
      if(xact_type == ATOMIC){
         tag_op inside {TAG_INVALID,TAG_FETCH_MATCH};}
      if(xact_type == COHERENT)  {
        if(coherent_xact_type == WRITENOSNOOP){
          tag_op  inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};}
        else if(coherent_xact_type inside {WRITEUNIQUE,WRITELINEUNIQUE}) {
          tag_op  inside {TAG_INVALID,TAG_UPDATE};}
        else if (coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO}){
          tag_op inside {TAG_INVALID,TAG_TRANSFER,TAG_UPDATE};}
        else if (coherent_xact_type inside{CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION}){
          tag_op == TAG_INVALID;}
         }
       if(xact_type == WRITE){
         tag_op inside {TAG_INVALID,TAG_UPDATE,TAG_TRANSFER,TAG_FETCH_MATCH};
        }
       }
     }
  if(transmitted_channel == READ) {
    tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH};
    if(xact_type == COHERENT)  {
      if(coherent_xact_type == READNOSNOOP){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
      else if (coherent_xact_type == READONCE){
       tag_op  inside {TAG_INVALID,TAG_TRANSFER};}
      else if (coherent_xact_type inside {READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE}){
      tag_op ==TAG_INVALID;}
    }
   if(xact_type == READ){
      tag_op  inside {TAG_INVALID,TAG_TRANSFER,TAG_FETCH_MATCH}; }
  }
  if (tag_op != TAG_INVALID){
  // Transactions must be cacheline sized or smaller
  //For an INCR burst, the last byte in the burst, as determined from the burst length in bytes,
  //(AWSIZE x AWLEN), added to the AWSIZE aligned start address, must be within the same
  //cache line as the first byte in the burst
  //i.e addr_aligned_to_burst_size + bytes_in_transfer < addr_aligned_to_cache_line_size + cache_line_size
      (burst_type == INCR) -> (((addr >> burst_size) << burst_size) + (burst_length << burst_size) <= 
      ((addr >> log_base_2_cache_line_size) << log_base_2_cache_line_size) + port_cfg.cache_line_size);
   // For a WRAP burst, AWSIZE x AWLEN must not exceed the cache line size.
      (burst_type == WRAP) -> ((burst_length << burst_size) <= port_cfg.cache_line_size);

 // For INCR transactions address must be aligned to container size
    if(burst_type == INCR){
     addr == addr >> (burst_length << burst_size) << (burst_length << burst_size);
    }

  // For WRAP transactions address must be aligned to burst_size
    if(burst_type == WRAP){
      addr == addr >> burst_size << burst_size; }

    cache_type[3:2] != 2'b00;
    cache_type[1:0] == 2'b11; 
   }
  if(tag_op == TAG_INVALID){
    foreach(tag[i])
      tag[i] == 0;}

  // Transaction type inside READ,WRITE,COHERENT and ATOMIC  
  xact_type inside {READ,WRITE,COHERENT,ATOMIC};
  if(xact_type == COHERENT){
    coherent_xact_type inside {WRITENOSNOOP,WRITEUNIQUE,WRITELINEUNIQUE,CMO,WRITEUNIQUEPTLSTASH,WRITEUNIQUEFULLSTASH,STASHONCESHARED,STASHONCEUNIQUE,STASHTRANSLATION,WRITEPTLCMO,WRITEFULLCMO,
                                READNOSNOOP,READONCE,READONCEMAKEINVALID,READONCECLEANINVALID,CLEANINVALID,MAKEINVALID,CLEANSHARED,CLEANSHAREDPERSIST,DVMMESSAGE,DVMCOMPLETE};
  }
  }
}
// constraints on response_tag_op only applicable in external port monitor mode
 if(port_cfg.mte_support_type != svt_axi_port_configuration::NOT_SUPPORTED && port_cfg.use_external_port_monitor ==1){
   if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE){
     if(port_cfg.use_external_port_monitor == 1){
       if(transmitted_channel == READ){
         if(tag_op == TAG_INVALID){
          response_tag_op inside {TAG_INVALID,TAG_TRANSFER};}
         else if(tag_op == TAG_TRANSFER){
         response_tag_op == TAG_TRANSFER};
        }
       else if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
         response_tag_op == TAG_INVALID;
       }
     }
     else {
       response_tag_op == TAG_INVALID;
     }
     if(transmitted_channel == READ_WRITE || transmitted_channel == WRITE){
      tag_match_resp inside{ MATCH_NOT_PERFORMED,NO_MATCH_RESULT,FAIL, PASS};
     }
     else if(transmitted_channel == READ){
      tag_match_resp == MATCH_NOT_PERFORMED;
     }
   }
 }
`endif
 }

// These constraints are applicable for MPAM feature
constraint mpam_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if (port_cfg.enable_mpam == svt_axi_port_configuration::MPAM_FALSE && port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER && port_cfg.is_active) {
    mpam_partid == 0;
    mpam_perfmongroup == 0;
    mpam_ns == prot_type[1];
  } 
`endif
}

// These constraints are applicable for Write with CMO transactions 
 constraint write_with_cmo_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE
  if(xact_type == COHERENT && (coherent_xact_type == WRITEPTLCMO || coherent_xact_type == WRITEFULLCMO)){
    domain_type inside {INNERSHAREABLE,OUTERSHAREABLE,NONSHAREABLE};
    atomic_type == NORMAL;
    cache_type[1] == 1;
  }
 if(port_cfg.axi_interface_type != svt_axi_port_configuration::ACE_LITE){
   !(coherent_xact_type inside {CMO,WRITEPTLCMO,WRITEFULLCMO});
  } 
 if(port_cfg.write_plus_cmo_enable != 1){
    !(coherent_xact_type inside {WRITEPTLCMO,WRITEFULLCMO});
  }
 if(port_cfg.cmo_on_write_enable != 1){
   coherent_xact_type != CMO;
 }
`endif
 }
 //These constraints are valid for atomic transactions .
constraint atomic_xacts_valid_ranges {
`ifdef SVT_ACE5_ENABLE 
   if(!port_cfg.axi_interface_type inside{svt_axi_port_configuration::AXI4,svt_axi_port_configuration::ACE_LITE})  {
      xact_type != ATOMIC;}
//   if(port_cfg.check_type != svt_axi_port_configuration::ODD_PARITY_BYTE_DATA){
//      atomic_read_is_datachk_parity_error == 0;}
   if(xact_type ==ATOMIC){
  //  data size should be equal to burst length
     if(port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
      
      if((barrier_type == NORMAL_ACCESS_RESPECT_BARRIER) || (barrier_type == NORMAL_ACCESS_IGNORE_BARRIER)){ 
          if ((domain_type == NONSHAREABLE) || (domain_type == SYSTEMSHAREABLE)){
             coherent_xact_type  == WRITENOSNOOP;}
          else{
             coherent_xact_type  == WRITEUNIQUE;}
        }
        else{
           coherent_xact_type == WRITEBARRIER;}
       if(burst_length > 1 && ! port_cfg.allow_multibeat_atomic_transactions_to_be_less_than_data_width){
         (1 << burst_size) == port_cfg.data_width/8;
       }
       data.size() == burst_length;
       wstrb.size() == burst_length;
       if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] == ((1 << (1 << burst_size)) - 1);
        }
      }
      awakeup_assert_delay ==0;
       if( atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN}){
          atomic_transaction_type == LOAD;
         }
       if(atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN}) {
          atomic_transaction_type == STORE;
        }
       if(atomic_xact_op_type == ATOMICSWAP){
          atomic_transaction_type == SWAP;
        }
       if(atomic_xact_op_type == ATOMICCOMPARE){
         atomic_transaction_type == COMPARE;
         burst_size inside{0,1,2,3,4,5};
         {((1 << burst_size)) * burst_length} inside {2,4,8,16,32};
         if(burst_length << burst_size == 2 && addr[0]==1'b0){ 
           burst_type == INCR;}
         else if(burst_length << burst_size == 4 && addr[1:0]==2'b0) {
            burst_type == INCR;}
         else if(burst_length << burst_size == 8 && addr[2:0]==3'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 16 && addr[3:0]==4'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 32 && addr[4:0]==5'b0) {
           burst_type == INCR;}
         else if(burst_length << burst_size == 2 && addr[0] !=1'b0){
           burst_type == WRAP;}
         else if(burst_length << burst_size == 4 && addr[1:0] !=2'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 8 && addr[2:0] !=3'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 16 && addr[3:0] !=4'b0) {
           burst_type == WRAP;}
         else if(burst_length << burst_size == 32 && addr[4:0] !=5'b0) {
           burst_type == WRAP;}
          } 
        atomic_transaction_type != NON_ATOMIC;
        if(atomic_transaction_type == COMPARE ){
           atomic_swap_data.size() == burst_length;
           atomic_compare_data.size() == burst_length;
           atomic_compare_wstrb.size() == burst_length;
           atomic_swap_wstrb.size() == burst_length;
           foreach(atomic_swap_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_swap_data[index] == atomic_swap_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           foreach(atomic_compare_data[index]) {
             if(port_cfg.wysiwyg_enable ==1'b1){
                atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
            }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_swap_data[index]) {
               atomic_swap_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
           if (!port_cfg.wysiwyg_enable) {
             foreach (atomic_compare_data[index]) {
               atomic_compare_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
             } 
           }
        }
        else {
           atomic_swap_data.size() == 0;
           atomic_compare_data.size() == 0;
           atomic_compare_wstrb.size() ==0;
           atomic_swap_wstrb.size() ==0;
         }
         if(atomic_transaction_type ==LOAD){
           atomic_xact_op_type inside{ATOMICLOAD_ADD,ATOMICLOAD_CLR,ATOMICLOAD_EOR,ATOMICLOAD_SET,ATOMICLOAD_SMAX,ATOMICLOAD_SMIN,ATOMICLOAD_UMAX,ATOMICLOAD_UMIN};}
         else if(atomic_transaction_type ==STORE){
           atomic_xact_op_type inside{ATOMICSTORE_ADD,ATOMICSTORE_CLR,ATOMICSTORE_EOR,ATOMICSTORE_SET,ATOMICSTORE_SMAX,ATOMICSTORE_SMIN,ATOMICSTORE_UMAX,ATOMICSTORE_UMIN};}
         else if(atomic_transaction_type ==SWAP){
           atomic_xact_op_type inside{ATOMICSWAP};}
         else if(atomic_transaction_type ==COMPARE){
           atomic_xact_op_type inside{ATOMICCOMPARE};}

//     Address for atomic transactions must be aligned to the data size
         if(atomic_transaction_type !=COMPARE){
           burst_size inside {0,1,2,3};
           {((1 << burst_size)) * burst_length} inside {1,2,4,8};
           burst_type==INCR;
           if (burst_length << burst_size == 2) {
              addr[0] == 1'b0;
            } 
            else if (burst_length << burst_size == 4) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 8) {
              addr[2:0] == 3'b0;
            } 
          }
//   For an Atomic compare transactions address must be aligned to half of the burst_size
         else if(atomic_transaction_type == COMPARE){
           burst_size inside {0,1,2,3,4,5};
            if(burst_length << burst_size == 4){
              addr[0] == 1'b0;}
            else if (burst_length << burst_size == 8) {
              addr[1:0] == 2'b0;
            } 
            else if (burst_length << burst_size == 16) {
              addr[2:0] == 3'b0;
            } 
           else if(burst_length << burst_size == 32){
              addr[3:0] == 4'b0;
           }
         }

       if(atomic_transaction_type == COMPARE) {
         atomic_swap_wstrb.size() == burst_length;
         atomic_compare_wstrb.size() == burst_length;
         }
       else {
         atomic_swap_wstrb.size() == 0;
         atomic_compare_wstrb.size() == 0;
       }
     if(atomic_transaction_type != COMPARE){
         burst_type == INCR;
         burst_size inside {0,1,2,3};
        }
       else if(atomic_transaction_type == COMPARE){
         burst_type inside{INCR,WRAP};
         burst_size inside{0,1,2,3,4,5};
        }
         if(xact_type ==ATOMIC){
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
         }
    }

  /* 
   * 1) Constraint the atomic_read_data_trace_tag to 1 based on trace_tag value
   */
    if(port_cfg.axi_port_kind == svt_axi_port_configuration:: AXI_SLAVE){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
       if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        atomic_read_data.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
        atomic_read_poison.size() == burst_length;

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}

      }
      if(atomic_transaction_type == COMPARE && xact_type ==ATOMIC){
        if(burst_length > 1){
          atomic_read_data.size() == burst_length/2;
          atomic_read_data_user.size() == burst_length/2;
          atomic_read_poison.size() == burst_length/2;
        }
        else {
          atomic_read_data.size() == 1;
          atomic_read_data_user.size() == 1;
          atomic_read_poison.size() == 1;
        }

        foreach(atomic_read_data[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data[index] == atomic_read_data[index] & atomic_comp_read_data_mask;}
          }

        foreach(atomic_read_data_user[index]) {
           if(port_cfg.wysiwyg_enable ==1'b1){
              atomic_read_data_user[index] == atomic_read_data_user[index] & atomic_comp_read_data_mask;}
          }
 
         if(port_cfg.poison_enable ==1){
           if(port_cfg.data_width>64){
             foreach(atomic_read_poison[index]) {
               if(port_cfg.wysiwyg_enable ==1'b1){
                 atomic_read_poison[index] == atomic_read_poison[index] & atomic_read_poison_mask;}
         }}}

         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data[index]) {
             atomic_read_data[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if (!port_cfg.wysiwyg_enable) {
           foreach (atomic_read_data_user[index]) {
             atomic_read_data_user[index] <= ((1 << (((1 << burst_size)>>1) << 3)) - 1);
           } 
         }
         if(port_cfg.poison_enable ==1){
           if (!port_cfg.wysiwyg_enable) {
             if(burst_size>3){
               foreach (atomic_read_poison[index]) {
                 atomic_read_poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);
               } 
         }}}
        }

      if(trace_tag ==1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        atomic_read_data_trace_tag == 1;
       }
      if(atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC){
        rvalid_delay.size() == burst_length;
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};
            }
       wready_delay.size()==burst_length;
    }

  }
    if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
     }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE} ){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
    
/*     if(xact_type == ATOMIC) {
       if(burst_length > 1){
          1 << burst_size == data_width_in_bytes;}
      }*/
  if(xact_type != ATOMIC)
    {
       atomic_read_data.size() ==0;
       atomic_read_poison.size() ==0;
       atomic_read_data_user.size() ==0;
       atomic_swap_data.size() ==0;
       atomic_compare_data.size() ==0;
       atomic_swap_wstrb.size()==0;
       atomic_compare_wstrb.size()==0;
       atomic_transaction_type == NON_ATOMIC;
    }
   if(xact_type ==ATOMIC){
     atomic_type == NORMAL;
     random_interleave_array.size() == burst_length;
     random_interleave_array[0] == 1;
    }
     xact_type != READ_WRITE;
     converted_xact_type != READ_WRITE;
     transmitted_channel != ATOMIC;
`endif
}

  // ACE/ACE-Lite Constraints Block. These constraints are valid if the
  // interface type is set to ACE or ACE-Lite.

  constraint ace_valid_ranges {

    foreach(data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
    }

`ifdef SVT_ACE5_ENABLE
   if(port_cfg.atomic_transactions_enable ==1'b1 && atomic_transaction_type inside{LOAD,SWAP,COMPARE} && xact_type == ATOMIC) {
      foreach(atomic_read_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data[index] == atomic_read_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

      foreach(atomic_read_data_user[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_read_data_user[index] == atomic_read_data_user[index] & ((1<<(port_cfg.data_width))-1);}
    }

     foreach(atomic_swap_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_swap_data[index] == atomic_swap_data[index] & ((1<<((port_cfg.data_width)))-1);}
    }
      foreach(atomic_compare_data[index]) {
      if(port_cfg.wysiwyg_enable ==1'b1){
        atomic_compare_data[index] == atomic_compare_data[index] & ((1<<(port_cfg.data_width))-1);}
    }

   if(port_cfg.poison_enable ==1 && port_cfg.wysiwyg_enable ==1){
       foreach(atomic_read_poison[index]) {
         if(port_cfg.data_width%64 == 0) {
           atomic_read_poison[index] == atomic_read_poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
           atomic_read_poison[index] == atomic_read_poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
   }}
  }
`endif

 if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
         if(port_cfg.data_width%64 == 0) {
            poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
         else {
            poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
    }}
   }
   
`ifdef SVT_ACE5_ENABLE
// This transaction types are not yet supported  
   !(coherent_xact_type inside {STASHTRANSLATION});
`endif 

`ifdef SVT_AXI_SVC_USE_MODEL
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration :: AXI_ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
   }
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
     if (`SVT_AXI_COHERENT_READ_1_BEAT) { 
       random_interleave_array.size() == 1;
       random_interleave_array[0] == 1;
     }
`ifdef INCA
     if ((slave_xact_type == COHERENT) && (slave_xact_type != DATA_STREAM )) {
        if( 
            (slave_coherent_xact_type == CLEANUNIQUE) || 
            (slave_coherent_xact_type == MAKEUNIQUE) || 
            (slave_coherent_xact_type == CLEANSHARED) ||
            (slave_coherent_xact_type == CLEANSHAREDPERSIST) ||
            (slave_coherent_xact_type == CLEANINVALID) || 
            (slave_coherent_xact_type == MAKEINVALID) 
          ) {
          wready_delay.size() == 1;
          rvalid_delay.size() == 1;
        }
        else {
          wready_delay.size() == burst_length;
          rvalid_delay.size() == burst_length;
        }
     }
`else  
     if ((xact_type == COHERENT) && 
         (xact_type != DATA_STREAM)) {
       if( 
           (coherent_xact_type == CLEANUNIQUE) || 
           (coherent_xact_type == MAKEUNIQUE) || 
           (coherent_xact_type == CLEANSHARED) || 
           (coherent_xact_type == CLEANSHAREDPERSIST) ||
           (coherent_xact_type == CLEANINVALID) || 
           (coherent_xact_type == MAKEINVALID) 
         ) {
         wready_delay.size() == 1;
         rvalid_delay.size() == 1;
       } else {
         wready_delay.size() == burst_length;
         rvalid_delay.size() == burst_length;
       }
     }  
`endif // `ifdef INCA 
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
   } //       if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE || `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE)
`endif //SVT_AXI_SVC_USE_MODEL
 } // ace_valid_ranges

  // AXI4 STREAM Constraints Block. These constraints are valid if the
  // interface type is set to AXI4_STREAM.
  constraint axi4_stream_valid_ranges {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif   
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
        random_interleave_array.size() == stream_burst_length;
        foreach (random_interleave_array[index]) {
          random_interleave_array[index] inside {[1 : stream_burst_length]};
        }   
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM)
   } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE)
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
     if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
`endif
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tid_enable) {
`else
       if (!port_cfg.tid_enable) {
`endif
         tid == 0;
       }
       else {
         tid inside {[0 : ((1 << port_cfg.tid_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdest_enable) {
`else
       if (!port_cfg.tdest_enable) {
`endif
         tdest == 0;
       }
       else {
         tdest inside {[0 : ((1 << port_cfg.tdest_width) -1)]};
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tdata_enable) {
`else
       if (!port_cfg.tdata_enable) {
`endif
         foreach (tdata[index])
           tdata[index] == 0;
       }
       else {
         foreach (tdata[index]) {
             tdata[index] inside {[0 : ((1 << port_cfg.tdata_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tstrb_enable) {
`else
       if (!port_cfg.tstrb_enable) {
`endif
         foreach(tstrb[index])
           tstrb[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tuser_enable) {
`else
       if (!port_cfg.tuser_enable) {
`endif
         foreach(tuser[index])
           tuser[index] == 0;
       }
       else {
         foreach (tuser[index]) {
            tuser[index] inside {[0 : ((1 << port_cfg.tuser_width) -1)]};
          }
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tkeep_enable) {
`else
       if (!port_cfg.tkeep_enable) {
`endif
         foreach(tkeep[index])
           tkeep[index] == 0;
       }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
       if (!tlast_enable) {
`else
       if (!port_cfg.tlast_enable) {
`endif
         stream_burst_length == 1;
       }
     } //AXI4_STREAM
   } //AXI_MASTER    
  } // axi4_stream_valid_ranges  


  // AXI3/AXI4/AXI4 Lite Constraints Block. These constraints are valid if the
  // interface type is set to either AXI3/AXI4/AXI4_Lite. Since these are
  // basic AXI constraints they even hold true in case the interface_type is
  // set to ACE/ACE_Lite.

  constraint axi3_4_valid_ranges {
    /*solve burst_length before random_interleave_array;
    solve stream_burst_length before random_interleave_array;
    solve burst_length before addr;
    solve burst_length before wstrb;

    solve burst_size before wstrb;
    solve burst_length before rresp;
    solve burst_length before coh_rresp;
    solve burst_length before rvalid_delay;
    solve burst_length before wready_delay;
    solve xact_type before rvalid_delay;
    solve xact_type before wready_delay;
    solve coherent_xact_type before rvalid_delay;
    solve coherent_xact_type before wready_delay;
    solve xact_type before rresp;
    solve coherent_xact_type before rresp;
    solve xact_type before coh_rresp;
    solve coherent_xact_type before coh_rresp;
    */

  foreach(data[index]) {
     if(port_cfg.wysiwyg_enable ==1'b1){
       data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
   }

   if(port_cfg.poison_enable ==1){
      foreach(poison[index]) {
        if(port_cfg.wysiwyg_enable ==1'b1){
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
      }
    }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
    burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
`else
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI3)
      burst_length <= `SVT_AXI3_MAX_BURST_LENGTH;
    else
      burst_length <= `SVT_AXI4_MAX_BURST_LENGTH;
`endif //SVT_AXI_SVC_NO_CFG_IN_XACT
      if(port_cfg.ace_version == svt_axi_port_configuration::ACE_VERSION_1_0 && xact_type == COHERENT) {
        !(coherent_xact_type inside{CLEANSHAREDPERSIST,READONCECLEANINVALID,READONCEMAKEINVALID});}

`ifdef SVT_AXI_SVC_USE_MODEL

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_MASTER) {
`endif
      // Constraining the Delay sizes
      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        wvalid_delay.size() == 1;
        rready_delay.size() == 1;
        data.size() == 1;
        if(port_cfg.poison_enable ==1){
        poison.size() == 1;}
      } else if (xact_type != DATA_STREAM) {
        wvalid_delay.size() == burst_length;
        rready_delay.size() == burst_length;
        data.size() == burst_length;
       if(port_cfg.poison_enable ==1){
       poison.size() == burst_length;
      }}

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (port_cfg.toggle_ready_signals_during_idle_period) {
        if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          idle_rready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY_ARR_SIZE]};
          idle_bready_delay.size() == 0;
        } else {
          idle_bready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY_ARR_SIZE]};
          idle_rready_delay.size() == 0; 
        }
      } else {
        idle_rready_delay.size() == 0;
        idle_bready_delay.size() == 0;
      }

     if (!port_cfg.wysiwyg_enable) {
        foreach (data[index]) {
          data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        } 
      }
     foreach(data[index]) {
       if(port_cfg.wysiwyg_enable ==1'b1){
         data[index] == data[index] & ((1<<(port_cfg.data_width))-1);}
      }

    if(port_cfg.poison_enable ==1 && !port_cfg.wysiwyg_enable){
        foreach (poison[index]) {
          if((1 << burst_size)%8 !=0){
            poison[index] <= ((1 << (((1 << burst_size) >> 3)+1)) - 1);}
          else {
             poison[index] <= ((1 << ((1 << burst_size) >> 3)) - 1);}
        } 
      }

   if(port_cfg.poison_enable ==1  && port_cfg.wysiwyg_enable ==1){
      foreach(poison[index]) {
           if(port_cfg.data_width%64 == 0) {
              poison[index] == poison[index] & ((1<<(port_cfg.data_width/64))-1);}
           else {
              poison[index] == poison[index] & (((1<<(port_cfg.data_width/64)+1))-1);}
        }
    }
`endif

      /*
       * 1) Constrain the array size to 0 if xact_type is not READ
       * 2) Constrain the array size to burst length if xact_type is READ
       */    
      if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
        if (`SVT_AXI_COHERENT_READ_1_BEAT) 
          rresp.size() == 1;
        else
          rresp.size() == burst_length; 
      }
`ifdef SVT_ACE5_ENABLE
     else if(xact_type == ATOMIC && atomic_transaction_type inside{LOAD,SWAP} ){
       rresp.size()== burst_length ;
      }
     if(xact_type == ATOMIC && atomic_transaction_type inside{COMPARE}){
       if(burst_length > 1){
         rresp.size()== burst_length/2 ;}
       else {
         rresp.size() ==1;}
     }
`endif      
      else {
        rresp.size() == 0;
      }

      /* 
       *  Constraints for wstrb 
       *  1) Constraint the length of the wstrb from 1 to burst_length for write
         transactions
       *  2) Constraining wstrb to enable all the valid bytelanes depending on transfer
      */
      if (xact_type == WRITE || (`SVT_AXI_COHERENT_WRITE) 
`ifdef SVT_ACE5_ENABLE
|| xact_type ==ATOMIC
`endif    
       ) {
        wstrb.size() == burst_length;
      }
      else
        wstrb.size() == 0;
      /*if (!port_cfg.wysiwyg_enable) {
        foreach (wstrb[index]) {
          wstrb[index] inside {[0: ((1 << (1 << burst_size)) - 1)]};
        }
      }
      */
`ifdef SVT_ACE5_ENABLE
       if(xact_type == ATOMIC){
          data.size() == burst_length;
       }
`endif

      if (`SVT_AXI_COHERENT_READ_1_BEAT) {
        data_user.size() == 1;
      } else if (xact_type == DATA_STREAM) {
        data_user.size() == 0;
      } else {
        data_user.size() == burst_length;
      }
`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
`ifdef SVT_ACE5_ENABLE 
    xact_type inside {READ,WRITE,IDLE,COHERENT,ATOMIC};
`else
    xact_type inside {READ,WRITE,IDLE,COHERENT,DATA_STREAM};
`endif
`endif

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        xact_type != DATA_STREAM;

`ifdef SVT_MULTI_SIM_ENUM_RANDOMIZES_TO_INVALID_VALUE
        atomic_type inside {NORMAL,EXCLUSIVE,LOCKED};
        burst_type inside {FIXED,INCR,WRAP};
`endif

`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT
        /* 
         * The atomic type is not exclusive when exclusive_access_enable is
         * disabled
         */  
        if (port_cfg.exclusive_access_enable == 0) {
          atomic_type != EXCLUSIVE;    
        }
        if (port_cfg.locked_access_enable == 0) {
          atomic_type != LOCKED;    
        }
`endif
        
        
        /** Address is within limits specified by addr_width. */
        addr <= max_possible_addr;
        addr_user <= max_possible_user_addr;

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        id <= ((1 << `SVT_AXI_MAX_ID_WIDTH) - 1);
`else
        if (port_cfg.use_separate_rd_wr_chan_id_width == 0 
`ifdef SVT_ACE5_ENABLE
          || xact_type == ATOMIC
`endif
         ) 
          id <= ((1 << port_cfg.id_width) - 1);
        else if ((xact_type == WRITE) || `SVT_AXI_COHERENT_WRITE)
          id <= ((1 << port_cfg.write_chan_id_width) - 1);
        else 
          id <= ((1 << port_cfg.read_chan_id_width) - 1);
`endif

        /*
         *  When the burst type is not Fixed, it must be ensured that burst does not
         *  exceed 4k range
         */
   
        if(burst_type != FIXED) {
          addr_range == (burst_length * (1 << burst_size));
          `ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
          addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << burst_size);
          `else
          addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << burst_size);
          `endif  
          if (burst_type == WRAP) {
            // Make sure that the max address does not cross addr_width.
            // Need to calculate this from wrap boundary (lowest address)
            // Note that the max byte address is:
            // (burst_length-1)*bytes_in_each_transfer + (bytes_in_each_transfer-1)
            if (burst_length == 2)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+1));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+1));
`endif
            else if (burst_length == 4)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+2));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+2));
`endif
            else if (burst_length == 8)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+3));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+3));
`endif
            else if (burst_length == 16)
`ifdef SVT_MULTI_SIM_CONSTRAINT_SHIFT_CONSTANT_RESULTS_IN_X_OR_Z
              burst_addr_mask == ( `SVT_AXI_MAX_ADDR_WIDTH'hffff_ffff_ffff_ffff << (burst_size+4));
`else
              burst_addr_mask == ( {`SVT_AXI_MAX_ADDR_WIDTH{1'b1}} << (burst_size+4));
`endif

            addr == (addr & addr_mask);
            (addr & burst_addr_mask) + addr_range - 1 <= max_possible_addr; 
            (addr[11:0] & burst_addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
          } else {
            // INCR
            (addr[11:0] & addr_mask) <= (`SVT_AXI_TRANSACTION_4K_ADDR_RANGE - addr_range);
            // Make sure that the max address does not cross addr_width.
            // Use aligned address
            ((addr >> burst_size) << burst_size) + addr_range - 1 <= max_possible_addr;
          }
        } 


        
        // Resetting all the bits greater than data width to 0

        /*foreach (wstrb[index]) {
          if (index < burst_length) {
            wstrb[index] == wstrb[index] & ((1 << port_cfg.data_width/8)-1);
          } 
        }
        */


        addr_valid_delay inside {[0:`SVT_AXI_MAX_ADDR_VALID_DELAY]};
        

        foreach (wvalid_delay[index]) {
          wvalid_delay[index] inside {[0:`SVT_AXI_MAX_WVALID_DELAY]};
        }
        foreach (rready_delay[index]) {
          rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
        }
        foreach (idle_rready_delay[index]) {
          idle_rready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_RREADY_DELAY]};
        }

        /*if (reference_event_for_rready_delay == MANUAL_RREADY) {
          foreach (rready_delay[index]) {
            (index == 0) -> rready_delay[index] inside {[-`SVT_AXI_MAX_RREADY_DELAY : `SVT_AXI_MAX_RREADY_DELAY]};
            (index > 0)  -> rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        } else {
          foreach (rready_delay[index]) {
            rready_delay[index] inside {[0:`SVT_AXI_MAX_RREADY_DELAY]};
          }
        }
        */

        bready_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        foreach (idle_bready_delay[index]) {
          idle_bready_delay[index] inside {[0:`SVT_AXI_MAX_IDLE_BREADY_DELAY]};
        }


        // Data Before Addr Constraints
        if(data_before_addr) {
          reference_event_for_first_wvalid_delay == PREV_WRITE_DATA_HANDSHAKE;
          reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR,FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR};
        }

        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) {

          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } // if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) 

      // For EXCLUSIVE access, the address must be aligned to 
      // the total number of bytes transferred
      if (atomic_type == EXCLUSIVE) {
        (burst_length << burst_size) inside {1,2,4,8,16,32,64,128};

        if (burst_length << burst_size == 2) {
          addr[0] == 1'b0;
        } 
        else if (burst_length << burst_size == 4) {
          addr[1:0] == 2'b0;
        } 
        else if (burst_length << burst_size == 8) {
          addr[2:0] == 3'b0;
        } 
        else if (burst_length << burst_size == 16) {
          addr[3:0] == 4'b0;
        } 
        else if (burst_length << burst_size == 32) {
          addr[4:0] == 5'b0;
        } 
        else if (burst_length << burst_size == 64) {
          addr[5:0] == 6'b0;
        } 
        else if (burst_length << burst_size == 128) {
          addr[6:0] == 7'b0;
        } 
      }

      /* 
       * AXI3 :
       * 1) Burst Size must not exceed the data width
       * 2) Burst Length for WRAP is inside 2,4,8,16
       * 3) Total No. of bytes to be transferred in an exclusive access burst must be a
       *   power of 2.  Max is 128  - Section 6.2.4
       * 4) Burst Length For Idle transactions must be from 1 to Max Idles
       * 5)
      */   

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type == svt_axi_port_configuration :: AXI3) {
`else
      if (port_cfg.axi_interface_type == svt_axi_port_configuration :: AXI3) {
`endif
 
        xact_type != COHERENT;
        burst_size <= log_base_2_data_width_in_bytes;

        if (xact_type == IDLE) {
          burst_length inside {[1:`SVT_AXI_MAX_TRANSACTION_IDLE_CYCLES]}; 
        } else {
          if (burst_type == WRAP) {
`ifdef SVT_ACE5_ENABLE
           if(xact_type == ATOMIC && atomic_transaction_type == COMPARE){
              burst_length inside {1,2,4,8,16,32};}
           else {
              burst_length inside {2,4,8,16};}
`else
             burst_length inside {2,4,8,16};
`endif
          } else {
            burst_length inside {[1:`SVT_AXI3_MAX_BURST_LENGTH]};
          }
        }

        // WA(bit 3) bit must not be high if C bit(bit 1) is low
        (cache_type[1] == 0) -> (cache_type[3] == 0);
        // Reserved values:
        cache_type != 4'b0100;
        cache_type != 4'b0101;
        cache_type != 4'b1000;
        cache_type != 4'b1001;
        cache_type != 4'b1100;
        cache_type != 4'b1101;
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      foreach(data_user[i])
       data_user[i] <= ((1 << `SVT_AXI_MAX_DATA_USER_WIDTH) - 1);
`else
      foreach(data_user[i])
       data_user[i] <= ((1 << port_cfg.data_user_width) - 1);
`endif
   }
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
   if (axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`else
   if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) {
`endif
`ifndef SVT_AXI_SVC_NO_CFG_IN_XACT

`ifdef SVT_ACE5_ENABLE    
   if(port_cfg.atomic_transactions_enable ==1){
      if(!(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         atomic_read_data.size() ==0;
         atomic_read_poison.size() ==0;
         atomic_read_data_user.size() ==0;
        }
      if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
         atomic_read_data.size() <= burst_length;
         atomic_read_poison.size() <= burst_length;
         atomic_read_data_user.size() <= burst_length;
       }
       if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
         if(burst_length > 1){
           atomic_read_data.size() == burst_length/2;
           atomic_read_poison.size() == burst_length/2;
           atomic_read_data_user.size() == burst_length/2;
         }
         else {
           atomic_read_data.size() == 1;
           atomic_read_poison.size() == 1;
           atomic_read_data_user.size() == 1;
         }
        }
      }
   else {
     atomic_read_data.size() ==0;
     atomic_read_data_user.size() ==0;
     atomic_read_poison.size() ==0;
//     atomic_resultant_data.size() ==0;
//     atomic_swap_data.size() ==0;
//     atomic_compare_data.size() ==0;
    }
`endif
      if (port_cfg.enable_delayed_response_port) {
        // Transaction supplied through delayed response port.
        // data.size() can be <= burst_length since data is provided
        // through multiple transactions.
        if (is_delayed_response_xact) {
          if (`SVT_AXI_COHERENT_READ_1_BEAT) {
           if(port_cfg.poison_enable ==1){
            poison.size() == 1;}
            data.size() == 1;
            rresp.size() == 1;
          } else if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
          if(port_cfg.poison_enable ==1){
            poison.size() <= burst_length;}
            data.size() <= burst_length;
            rresp.size() <= burst_length;
            data.size() == rresp.size();
          if(port_cfg.poison_enable ==1){
           poison.size() == rresp.size();}
          }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC ) {
        rresp.size() == burst_length;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;  }
      else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC ) {
        if(burst_length > 1){
        rresp.size() == burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length/2;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length/2;
        atomic_read_data_user.size() <= burst_length/2;
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        }
        else {
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() <= burst_length;
          poison.size() <= burst_length;}
        atomic_read_data.size() <= burst_length;
        atomic_read_data.size() == rresp.size();
        atomic_read_data_user.size() <= burst_length;
        atomic_read_data_user.size() == rresp.size();
        if(port_cfg.poison_enable ==1){
          atomic_read_poison.size() == rresp.size();}        
        data.size() <= burst_length;
        rresp.size() <= burst_length;}
       }
`endif  
       else {
            rresp.size() == 0;
          }  
        // Transaction supplied through seq_item_port but when
        // configured with enable_delayed_response_port. This corresponds
        // to the transaction handle that is returned in 0-time to the driver.
        } else {
          if ((xact_type == READ) || (`SVT_AXI_COHERENT_READ)) {
             data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
             rresp.size() == 0;
          // WRITES
          }
       else {
            rresp.size() == 0;
          }
        }
      } else 
`endif
      {
        if (xact_type == DATA_STREAM) {
          data.size() == 0;
           if(port_cfg.poison_enable ==1){
             poison.size() == 0;}
        } else if (`SVT_AXI_COHERENT_READ_1_BEAT) {
          data.size() == 1;
         if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
          rresp.size() == 1;
          data_user.size() == 1;
        } else if ((xact_type == READ) || `SVT_AXI_COHERENT_READ) {
          data.size() == burst_length;
          if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
          rresp.size() == burst_length;
          data_user.size() == burst_length;
        // WRITES. rresp_size should be 0.
        }
`ifdef SVT_ACE5_ENABLE
      else if(atomic_transaction_type inside{LOAD,SWAP} && xact_type == ATOMIC) {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       else if(atomic_transaction_type inside{COMPARE} && xact_type == ATOMIC) {
        if(burst_length >1){
        rresp.size() == burst_length/2;
        atomic_read_data.size() == burst_length/2;
        atomic_read_poison.size() == burst_length/2;
        atomic_read_data_user.size() == burst_length/2;
        }
       else {
        rresp.size() == burst_length;
        atomic_read_data.size() == burst_length;
        atomic_read_poison.size() == burst_length;
        atomic_read_data_user.size() == burst_length;
       }
       }
       else if(xact_type == ATOMIC && !(atomic_transaction_type inside{LOAD,SWAP,COMPARE})){
         rresp.size() ==0;
         atomic_read_data.size()==0;
         atomic_read_data_user.size()==0;
         atomic_read_poison.size()==0;
      }
`endif  
        else {
          data_user.size() == burst_length;
          data.size() == burst_length;
          rresp.size() == 0;
        }
      }

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      if (axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`else
      if (port_cfg.axi_interface_type != svt_axi_port_configuration::AXI4_STREAM) {
`endif
        if (!(`SVT_AXI_COHERENT_READ_1_BEAT)) { 
          random_interleave_array.size() == burst_length;
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[1 : burst_length]};
          }
        }
      } 

      addr_ready_delay inside {[0:`SVT_AXI_MAX_ADDR_DELAY]};

`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
      resp_user <= ((1 << `SVT_AXI_MAX_BRESP_USER_WIDTH) - 1);
`else
      resp_user <= ((1 << port_cfg.resp_user_width) - 1);
`endif


    // wready_delay[0] can take positive and negative values.
`ifdef INCA
      if ((slave_xact_type != COHERENT) && (slave_xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`else
      if ((xact_type != COHERENT) && (xact_type != DATA_STREAM )) {
        wready_delay.size() == burst_length;
        rvalid_delay.size() == burst_length;
      }
`endif
      if (port_cfg.toggle_ready_signals_during_idle_period)
        idle_addr_ready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY_ARR_SIZE]}; 
      else
        idle_addr_ready_delay.size() == 0;
      if (xact_type == WRITE 
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif           
         || xact_type == COHERENT && 
          (coherent_xact_type == WRITENOSNOOP ||
           coherent_xact_type == WRITELINEUNIQUE ||
           coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
           coherent_xact_type == WRITEBACK   ||
           coherent_xact_type == WRITECLEAN  ||
           coherent_xact_type == WRITEEVICT
          )
         ) {
        if (port_cfg.toggle_ready_signals_during_idle_period)
          idle_wready_delay.size() inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY_ARR_SIZE]}; 
        else
          idle_wready_delay.size() == 0;
      } else {
        idle_wready_delay.size() == 0;
      }
      if (xact_type != DATA_STREAM) {
       if(!port_cfg.axi_slv_channel_buffers_enable)
        foreach (rvalid_delay[idx])
          rvalid_delay[idx] inside {[0:`SVT_AXI_MAX_RVALID_DELAY]};

        if (reference_event_for_wready_delay == MANUAL_WREADY) {
          foreach (wready_delay[idx]) {
            (idx == 0) -> wready_delay[idx] inside {[-`SVT_AXI_MAX_WREADY_DELAY:`SVT_AXI_MAX_WREADY_DELAY]};
            (idx > 0) -> wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          }
        } else {
          foreach (wready_delay[idx])
            wready_delay[idx] inside {[0:`SVT_AXI_MAX_WREADY_DELAY]};
          foreach (idle_wready_delay[idx])
            idle_wready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_WREADY_DELAY]};
          foreach (idle_addr_ready_delay[idx])
            idle_addr_ready_delay[idx] inside {[0:`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY]};
        }
       if(!port_cfg.axi_slv_channel_buffers_enable)
        bvalid_delay inside {[`SVT_AXI_MIN_WRITE_RESP_DELAY:`SVT_AXI_MAX_WRITE_RESP_DELAY]};
        if (xact_type == WRITE  
`ifdef SVT_ACE5_ENABLE
         || xact_type == ATOMIC
`endif      
         ||   xact_type == COHERENT && 
             (coherent_xact_type == WRITENOSNOOP ||
             coherent_xact_type == WRITELINEUNIQUE ||
             coherent_xact_type == WRITEUNIQUE ||
`ifdef SVT_ACE5_ENABLE
             coherent_xact_type == WRITEUNIQUEPTLSTASH ||
             coherent_xact_type == WRITEUNIQUEFULLSTASH ||
`endif
             coherent_xact_type == WRITEBACK   ||
             coherent_xact_type == WRITECLEAN  ||
             coherent_xact_type == WRITEEVICT  ||
             coherent_xact_type == EVICT
            )
           ) {
        // The reordering priority of write responses be within
        // 1 to port_cfg.write_resp_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_WRITE_RESP_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.write_resp_reordering_depth]};
`endif
        }
        else { //if (xact_type == READ) 
        // The reordering priority of read transactions should be within
        // 1 to port_cfg.read_data_reordering_depth.
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        reordering_priority inside {[1:`SVT_AXI_MAX_READ_DATA_REORDERING_DEPTH]};
`else
        reordering_priority inside {[1:port_cfg.read_data_reordering_depth]};
`endif
        }

        // An EXOKAY response makes sense only for an EXLUSIVE type
        // atomic access.
        if (atomic_type != EXCLUSIVE) { 
          foreach (rresp[idx])
            (rresp[idx] != EXOKAY); 
          bresp != EXOKAY; 
        }

        if (
            (xact_type == COHERENT) && 
            ( 
              (coherent_xact_type == CLEANUNIQUE) || 
              (coherent_xact_type == MAKEUNIQUE) || 
              (coherent_xact_type == CLEANSHARED) || 
              (coherent_xact_type == CLEANSHAREDPERSIST) || 
              (coherent_xact_type == CLEANINVALID) || 
              (coherent_xact_type == MAKEINVALID) 
            ) 
           ) {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : 1]};
          }
        } else {
          foreach (random_interleave_array[index]) {
            random_interleave_array[index] inside {[0 : burst_length]};
          }
        }
      }
    } // if (port_cfg.axi_port_kind == svt_axi_port_configuration::AXI_SLAVE) 
`endif //SVT_AXI_SVC_USE_MODEL
  } // axi3_4_valid_ranges 

 
  constraint disable_constraint_first_wvalid_reference_event {
    reference_event_for_first_wvalid_delay dist { WRITE_ADDR_VALID:=50000, WRITE_ADDR_HANDSHAKE:=1, PREV_WRITE_DATA_HANDSHAKE:=50000 };
  }

 constraint valid_poison {
    if(port_cfg.poison_enable == 0){
       poison.size()==0;
    }
   }


`ifdef INCA 
   constraint validpoison {
     if(port_cfg.poison_enable==1 && port_cfg.ace_version==svt_axi_port_configuration::ACE_VERSION_2_0){
        poison.size()==1;
     }
     else {
       poison.size()==0;
     }
    }
`endif

`ifdef SVT_ACE5_ENABLE
    constraint valid_archunken{
	        if(port_cfg.rdata_chunking_enable == 1 && xact_type == READ){
		        if(burst_size >= BURST_SIZE_128BIT){
			        archunken inside {0,1};
                  }
		        else {
			        archunken == 0;
                }
            }
	        else {	
		        archunken == 0;
            }
        }

    constraint reasonable_ranges_while_chunking {
      solve chunk_length before rchunkstrb;
      solve chunk_length before rchunknum;
        if(archunken){
            rchunkstrb.size() == chunk_length;
            rchunknum.size() == chunk_length;
        }
        else {
            rchunkstrb.size() == 0;
            rchunknum.size() == 0;
        }
    }

    constraint reasonable_chunk_len{
      solve burst_length before chunk_length;
      solve burst_size before chunk_length;
      if(archunken){
        if(burst_size < BURST_SIZE_128BIT){
          chunk_length == 0;
        }
        else {
          chunk_length inside {[burst_length:(burst_length<<(burst_size - 4))]};
        }
      }
      else {
        chunk_length == 0;
      }
    }
`endif
 /*Reasonable constraint on reference_event_for_addr_delay in data_before_addr scenarios
 reference_event_for_addr_delay must not be set to FIRST_DATA_HANDSHAKE_DATA_BEFORE_ADDR as this may cause 
 potential deadlock scenarios in ACE SLAVE DUT where slave DUT waits for awvalid signal
 before driving wready signal.
 */
 constraint reasonable_reference_event_for_addr_delay {
   if(data_before_addr){
   reference_event_for_addr_valid_delay inside {FIRST_WVALID_DATA_BEFORE_ADDR};}
 }
    
`ifdef SVT_AXI_SVC_USE_MODEL
  // **************************************************************************
  //       Reasonable  Constraints
  // **************************************************************************

`protected
M^XA?.Qc5-GD&^O,?<cMP)F;e+;W>Y6D5=GaRJd6_@[L5_#GE2T&3)^Bc02=QV3\
HZY0.EHe-FVD-$
`endprotected

  constraint reasonable_burst_length {
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI3_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI3_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI3_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4 ||
        `SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  ACE_LITE) {  
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2: (`SVT_AXI4_MAX_BURST_LENGTH >> 2)] :/ SHORT_BURST_wt,
        [(`SVT_AXI4_MAX_BURST_LENGTH >> 2)+1:`SVT_AXI4_MAX_BURST_LENGTH] :/ LONG_BURST_wt
      };
    }
    if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI_ACE) {
      burst_length dist {
        1 := ZERO_BURST_wt,
        [2:4] :/ SHORT_BURST_wt,
        [5:16] :/ LONG_BURST_wt
      };
    }
  }

  /*
    Reasonable constraint for cache type.
    For exclusive accesses transactions , transactions must not be cached
  */
  constraint reasonable_cache_type
  {
    solve atomic_type before cache_type;
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI3) {   
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_3_NON_CACHEABLE_NON_BUFFERABLE,
                             `SVT_AXI_3_BUFFERABLE_OR_MODIFIABLE_ONLY,
                             `SVT_AXI_3_CACHEABLE_BUT_NO_ALLOC,
                             `SVT_AXI_3_CACHEABLE_BUFFERABLE_BUT_NO_ALLOC};
        }
      } 
      if (`SVT_AXI_INTERFACE_TYPE == svt_axi_port_configuration ::  AXI4) {
        if (atomic_type == EXCLUSIVE) {
          cache_type inside {`SVT_AXI_4_ARCACHE_DEVICE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_DEVICE_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_NON_BUFFERABLE,
                             `SVT_AXI_4_ARCACHE_NORMAL_NON_CACHABLE_BUFFERABLE};
        }
      } 
  }

  /* 
    Reasonable constraint for interleave_pattern
    1) Set the interleave pattern to RANDOM BLOCK for the user to set interleave
    patterns
  */  

  constraint reasonable_interleave_pattern {
    interleave_pattern == RANDOM_BLOCK;
  }

  /* 
    Reasonable constraint for equal block length
    1) Constrain the equal block length to range of 1 to burst_length/2
  */
  
  constraint reasonable_equal_block_length {
    solve interleave_pattern before equal_block_length;
    solve burst_length before equal_block_length;
    if (interleave_pattern ==  EQUAL_BLOCK) {
      if (burst_length > 1) {
        equal_block_length  inside {[1 : (burst_length >> 1)]};
      }
      else {
        equal_block_length == 1;
      }
    }
  }

  constraint reasonable_addr_valid_delay {
   addr_valid_delay dist {
     0 := ZERO_DELAY_wt, 
     [1:(`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
     [((`SVT_AXI_MAX_ADDR_VALID_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_VALID_DELAY] :/ LONG_DELAY_wt
   };
  }


  constraint reasonable_wakeup_assert_deassert_delay {
    awakeup_assert_delay >= `SVT_AXI_MIN_AWAKEUP_ASSERT_DELAY;
    awakeup_assert_delay <  `SVT_AXI_MAX_AWAKEUP_ASSERT_DELAY;
    awakeup_deassert_delay >= `SVT_AXI_MIN_AWAKEUP_DEASSERT_DELAY;
    awakeup_deassert_delay <  `SVT_AXI_MAX_AWAKEUP_DEASSERT_DELAY;
  }

  constraint reasonable_rready_delay {
    /*foreach (rready_delay[idx]) {
      if (reference_event_for_rready_delay == MANUAL_RREADY && idx == 0) {
        rready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_RREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_RREADY_DELAY: -((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {
          rready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] := SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] := LONG_DELAY_wt >> 1
          };
      }
    }
    */
    foreach (rready_delay[idx]) {
      rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  constraint reasonable_idle_rready_delay {
    foreach (idle_rready_delay[idx]) {
      idle_rready_delay[idx] dist {
            0 := ZERO_DELAY_wt,
            [1:(`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
            [((`SVT_AXI_MAX_IDLE_RREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_RREADY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  
  // Enforces a distribution based on the weights.
  constraint reasonable_wvalid_delay {
    foreach (wvalid_delay[idx]) {
      wvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_WVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WVALID_DELAY >> 2)+1):`SVT_AXI_MAX_WVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }


  // Enforces a distribution based on the weights.
  constraint reasonable_bready_delay {
    bready_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  constraint reasonable_idle_bready_delay {
    foreach (idle_bready_delay[i]) 
      idle_bready_delay[i] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_IDLE_BREADY_DELAY>> 2)+1):`SVT_AXI_MAX_IDLE_BREADY_DELAY] :/ LONG_DELAY_wt
    };
  }


  constraint reasonable_tready_delay {
    if (port_cfg.axi_interface_type == svt_axi_port_configuration::AXI4_STREAM) {
      tready_delay.size() == `SVT_AXI_MAX_STREAM_BURST_LENGTH;
      foreach (tready_delay[idx]) {
        tready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_TREADY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_TREADY_DELAY >> 2)+1):`SVT_AXI_MAX_TREADY_DELAY] :/ LONG_DELAY_wt
       };
      }
    } else {
      tready_delay.size() == 0;
    }
  }

  /** 
   * This constraint insures that unimplemented features are avoided during randomization.
   */
  constraint exclude_master_unimplemented_features
  {
    xact_type != IDLE;
    interleave_pattern != EQUAL_BLOCK;
    start_new_interleave == 0;
    reference_event_for_rready_delay != MANUAL_RREADY;
  }

  //--------------------------------------------------------------------------------------
  /**************************** SLAVE CONSTRAINTS ******************************** */
  constraint reasonable_data {
    if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
      if (
           (xact_type == READ) || 
           (
             (xact_type == COHERENT) &&
             (
               coherent_xact_type == READNOSNOOP                     ||
               coherent_xact_type == READONCE                        ||
               coherent_xact_type == READONCECLEANINVALID                        ||
               coherent_xact_type == READONCEMAKEINVALID                        ||
               coherent_xact_type == READSHARED                      ||
               coherent_xact_type == READCLEAN                       ||
               coherent_xact_type == READNOTSHAREDDIRTY              ||
               coherent_xact_type == READUNIQUE          
             )
           )
         ) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
         data.size() == burst_length;
         if(port_cfg.poison_enable ==1){
            poison.size() == burst_length;}
`else
       if (!port_cfg.enable_delayed_response_port) {
           if(port_cfg.poison_enable ==1){
             poison.size() == burst_length;}
           data.size() == burst_length;
       }
`endif
       data_user.size() == burst_length;
        foreach (data[index]) {
             data[index] <= ((1 << ((1 << burst_size) << 3)) - 1);
        }
      }
      // No data associated with these transactions 
      if(`SVT_AXI_COHERENT_READ_1_BEAT) {
`ifdef SVT_AXI_SVC_NO_CFG_IN_XACT
        if(port_cfg.poison_enable ==1){
           poison.size() == 1;}
        data.size() == 1;
`else
       if (!port_cfg.enable_delayed_response_port) {
          if(port_cfg.poison_enable ==1){
             poison.size() == 1;}
          data.size() == 1;
       }
`endif
       data_user.size() == 1;
        foreach (data[index]) {
             data[index] <= 0;
        }
      if(port_cfg.poison_enable ==1){
            foreach (poison[index]) {
             poison[index] <= 0;}
          }
      }
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_wready_delay {
    foreach (wready_delay[idx]) {
      // MANUAL_READY not supported.
      /*if (reference_event_for_wready_delay == MANUAL_WREADY && idx == 0) {
        wready_delay[idx] dist {
         0 := ZERO_DELAY_wt,
         [-(`SVT_AXI_MAX_WREADY_DELAY >> 2):-1] :/ SHORT_DELAY_wt >> 1,
         [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
         [-`SVT_AXI_MAX_WREADY_DELAY: -((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1)] :/ LONG_DELAY_wt >> 1,
         [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt >> 1
        };
      } else {*/ 
        wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_WREADY_DELAY] :/ LONG_DELAY_wt
          };
        //}
      }
    }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_wready_delay {
    foreach (idle_wready_delay[idx]) {
        idle_wready_delay[idx] dist {
          0 := ZERO_DELAY_wt,
          [1:(`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)] :/ SHORT_DELAY_wt >> 1,
          [((`SVT_AXI_MAX_IDLE_WREADY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_WREADY_DELAY] :/ LONG_DELAY_wt
          };
    }
  }
 

  // Enforces a distribution based on the weights.
  constraint reasonable_rvalid_delay {
    foreach (rvalid_delay[idx]) {
      rvalid_delay[idx] dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_RVALID_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_RVALID_DELAY >> 2)+1):`SVT_AXI_MAX_RVALID_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_addr_ready_delay {
    addr_ready_delay dist {
       0 := ZERO_DELAY_wt, 
       [1:(`SVT_AXI_MAX_ADDR_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_ADDR_DELAY >> 2)+1):`SVT_AXI_MAX_ADDR_DELAY] :/ LONG_DELAY_wt
    };
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_idle_addr_ready_delay {
    foreach (idle_addr_ready_delay[idx]) {
      idle_addr_ready_delay[idx] dist {
         0 := ZERO_DELAY_wt, 
         [1:(`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)] :/ SHORT_DELAY_wt,
         [((`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY >> 2)+1):`SVT_AXI_MAX_IDLE_ADDR_READY_DELAY] :/ LONG_DELAY_wt
      };
    }
  }

  // Enforces a distribution based on the weights.
  constraint reasonable_bvalid_delay {
    bvalid_delay dist {
       `SVT_AXI_MIN_WRITE_RESP_DELAY := ZERO_DELAY_wt, 
       [(`SVT_AXI_MIN_WRITE_RESP_DELAY + 1):(`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)] :/ SHORT_DELAY_wt,
       [((`SVT_AXI_MAX_WRITE_RESP_DELAY >> 2)+1):`SVT_AXI_MAX_WRITE_RESP_DELAY] :/ LONG_DELAY_wt
    };
  }

  /**
   * Reasonable constraint for random_interleave_array
   * Constraint the random interleave array from 1 to burstlength
   * If the  array values exceed the burst length, those values will be ignored
   */

   constraint reasonable_random_interleave_array {
     if (`SVT_AXI_INTERFACE_TYPE != svt_axi_port_configuration::AXI4_STREAM) {
       if(`SVT_AXI_COHERENT_READ_1_BEAT) 
         random_interleave_array.size() == 1;
       else
         random_interleave_array.size() == burst_length;

       foreach (random_interleave_array[index]) {
         random_interleave_array[index] inside {[1 : burst_length]};
       }
     } else {
       random_interleave_array.size() == stream_burst_length;
     }
   }

    constraint exclude_slave_unimplemented_features
    {
      interleave_pattern != EQUAL_BLOCK;
      start_new_interleave == 0;
      reference_event_for_wready_delay != MANUAL_WREADY;
    }

`endif

`ifdef SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
  /**
   * External constraint definitions which can be used for test level constraint addition.
   * By default, "test_constraintsX" constraints are not enabled in svt_axi_transaction. A
   * test can enable them by defining the following macro during the compile:
   *   SVT_AXI_TRANSACTION_ENABLE_TEST_CONSTRAINTS
   */
  constraint test_constraints1;
  constraint test_constraints2;
  constraint test_constraints3;
`endif

//reasonable  soft constraint for cust_xact_flow == 0. To support default behavior of cust_xact_flow disabled and overridden by user to enable it automatically whenever inline randomization constraint is added
constraint reasonable_cust_xact_flow {
  soft cust_xact_flow == 0;
} 

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * CONSTUCTOR: Create a new transaction instance, passing the appropriate argument
   * values to the parent class.
   *
   * @param name Instance name of the transaction
   */
  extern function new (string name = "svt_axi_transaction",svt_axi_port_configuration port_cfg_handle = null);
`else
`svt_vmm_data_new(`SVT_TRANSACTION_TYPE)
  extern function new (vmm_log log = null, svt_axi_port_configuration port_cfg_handle = null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) Tests the validity of the configuration
   * 2) calculate the log_2 of master configs data_width   
   */
  extern function void pre_randomize ();

  //----------------------------------------------------------------------------
  /**
   *   post_randomize does the following
   *   1) Aligns the address to no of Bytes for Exclusive Accesses
   */
  extern function void post_randomize ();

  /** returns 1 if status of all relevant phases of current transaction are assigned as ABORTED */
  extern virtual function bit is_aborted(int mode = 0);

  /** returns 1 if current transaction is configured as secure access */
  extern virtual function bit is_secure(bit allow_secure = 1);

  /** Returns 1 if current transaction is of device_type */
  extern virtual function bit is_device_type();

  /** Returns 1 if current transaction is DVM transaction */
  extern virtual function bit is_dvm_xact();

  /** Returns 1 if current transaction is cacheable transaction */
  extern virtual function bit is_cacheable_xact();

  /** Returns 1 if current transaction is allocate transaction */
  extern virtual function bit is_allocate_xact();

  /** Determines if this transaction is a CMO transaction */
  extern function bit is_cmo_xact();


//  /** Returns 1 if current transaction is of device_type or DVM transaction 
//   * Additinally this function will fire an error if device type or DVM transactions 
//   * are issued from not allowed ports 
//   */
//  extern virtual function bit skip_port_interleaving();

  /** waits for transaction to end */
  extern virtual task wait_for_transaction_end();


 /** waits for slave transaction to update the memory*/
  extern virtual task wait_for_write_transaction_to_update_memory();

  /** returns 1 if transaction status shows ended otherwise 0 */
  extern virtual function bit is_transaction_ended();

  /** waits for addr phase to end */
  extern virtual task wait_for_addr_phase_ended ();
  
  /** waits for data phase to end */
  extern virtual task wait_for_data_phase_ended();
  
  /** waits for write resp phase to end */
  extern virtual task wait_for_write_resp_phase_ended();

  /** mark end of transaction */
  extern virtual function void set_end_of_transaction(bit aborted=0);
  

   /**
  * Returns 1 if the specified error_kind is there in transaction, else returns 0 
  */
  extern virtual function bit has_axi_exception(int error_kind); 
  // ****************************************************************************
  //   SVT shorthand macros 
  // ****************************************************************************

  `svt_data_member_begin(svt_axi_transaction)
    `svt_field_object(port_cfg,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK| `SVT_REFERENCE, `SVT_HOW_REF)
    `ifndef INCA
    `svt_field_object      (exception_list,                             `SVT_ALL_ON|`SVT_DEEP|`SVT_NOCOMPARE|`SVT_UVM_NOPACK,  `SVT_HOW_DEEP)
    `endif
    `svt_field_object(associated_barrier_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`ifdef SVT_UVM_TECHNOLOGY
    `svt_field_object(causal_gp_xact,`SVT_ALL_ON|`SVT_NOCOMPARE|`SVT_NOPACK|`SVT_REFERENCE, `SVT_HOW_REF)
`endif

  // ****************************************************************************

  `svt_data_member_end(svt_axi_transaction)


  // ****************************************************************************
  // Methods
  // ****************************************************************************

  //----------------------------------------------------------------------------
  /**
   * Method to turn reasonable constraints on/off as a block.
   */
  extern virtual function int reasonable_constraint_mode (bit on_off);

  //----------------------------------------------------------------------------
  /**
   * Returns the class name for the object used for logging.
   */
  extern function string get_mcd_class_name ();

`ifdef SVT_VMM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
   * Extend the copy method to copy the transaction class fields.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

 `else
  //---------------------------------------------------------------------------
  /**
   * Extend the copy method to take care of the transaction fields and cleanup the exception xact pointers.
   *
   * @param rhs Source object to be copied.
   */
  extern virtual function void do_copy(`SVT_XVM(object) rhs);
`endif
 //----------------------------------------------------------------------------
  /**
   * Extend the svt_post_do_all_do_copy method to cleanup the exception xact pointers.
   * 
   * @param to Destination class for the copy operation
   */
  extern virtual function void svt_post_do_all_do_copy(`SVT_DATA_BASE_TYPE to);
 //----------------------------------------------------------------------------
  /**
   * Calculates whether the transaction is partial or full cacheline access.
   * returns 1, if transaction is full cacheline access. returns 0, if it is a 
   * partial cacheline access.
   * 
   * @param cacheline_size indicates the value of the master cache line size
   */
  extern virtual function bit is_full_cacheline(int cacheline_size);

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(uvm_object rhs, uvm_comparer comparer);
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with rhs..
   *
   * @param rhs Object to be compared against.
   * @param comparer TBD
   */
  extern virtual function bit do_compare(ovm_object rhs, ovm_comparer comparer);
`else
  // ---------------------------------------------------------------------------
  /**
   * Compares the object with to, based on the requested compare kind. Differences are
   * placed in diff.
   *
   * @param to vmm_data object to be compared against.
   * @param diff String indicating the differences between this and to.
   * @param kind This int indicates the type of compare to be attempted. Only supported
   * kind value is svt_data::COMPLETE, which results in comparisons of the non-static
   * data members. All other kind values result in a return value of 1.
   */
  extern virtual function bit do_compare (vmm_data to, output string diff, input int kind = -1);

  //----------------------------------------------------------------------------
  /**                         
   * Returns the size (in bytes) required by the byte_pack operation.
   *
   * @param kind This int indicates the type of byte_size being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in a size calculation based on the
   * non-static fields. All other kind values result in a return value of 0.
   */
  extern virtual function int unsigned byte_size (int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Packs the object into the bytes buffer, beginning at offset, based on the
   * requested byte_pack kind.
   *
   * @param bytes Buffer that will contain the packed bytes at the end of the operation.
   * @param offset Offset into bytes where the packing is to begin.
   * @param kind This int indicates the type of byte_pack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being packed and the return of an integer indicating the number of
   * packed bytes. All other kind values result in no change to the buffer contents, and a
   * return value of 0.
   */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1);

  //----------------------------------------------------------------------------
  /**
   * Unpacks the object from the bytes buffer, beginning at offset, based on
   * the requested byte_unpack kind.
   *
   * @param bytes Buffer containing the bytes to be unpacked.
   * @param offset Offset into bytes where the unpacking is to begin.
   * @param len Number of bytes to be unpacked.
   * @param kind This int indicates the type of byte_unpack being requested. Only supported
   * kind value is svt_data::COMPLETE, which results in all of the
   * non-static fields being unpacked and the return of an integer indicating the number of
   * unpacked bytes. All other kind values result in no change to the exception contents,
   * and a return value of 0.
   */
  extern virtual function int unsigned do_byte_unpack (const ref logic [7:0]
  bytes[], input int unsigned offset = 0, input int len = -1, input int kind = -1);

`endif

  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>read</i> access to public data members of this class.
   */
  extern virtual function bit get_prop_val (string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
   * HDL Support: For <i>write</i> access to public data members of this class.
   */
  extern virtual function bit set_prop_val (string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  /**
   * This method allocates a pattern containing svt_pattern_data instances for
   * all of the primitive data fields in the object. The svt_pattern_data::name
   * is set to the corresponding field name, the svt_pattern_data::value is set
   * to 0.
   *
   * @return An svt_pattern instance containing entries for all of the data fields.
   */
  extern virtual function svt_pattern do_allocate_pattern ();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB.  The pattern is customized to contain only the fields necessary for
   * the application and tranaction type.
   * 
   * Note:
   * As a performance enhancement, property values in the pattern are pre-populated when
   * the pattern is created.  This allows the FSDB writer infrastructure to skip the
   * get_prop_val_via_pattern step.
   *
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern allocate_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when a full tranaction is to be recorded.  Note that not all
   * properties are written.  Instead, only properties needed for debug are added.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_full_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is RADDR, RDATA, WADDR, WDATA, or WRESP.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_filtered_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the PA channel is "STREAM DATA".
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_stream_xml_pattern();

  // ---------------------------------------------------------------------------
  /**
   * Generates an SVT pattern object to represent the properties which are to be
   * written to FSDB when the pa_format_type is set to FSDB_PERF_ANALYSIS.
   * 
   * @return An svt_pattern instance containing entries to be written to FSDB
   */
   extern virtual function svt_pattern populate_perf_analysis_xml_pattern();

  // ----------------------------------------------------------------------------
  /**
   * This method returns PA object which contains the PA header information for XML or FSDB.
   *
   * @param uid Optional string indicating the unique identification value for object. If not 
   * provided uses the 'get_uid()' method  to retrieve the value. 
   * @param typ Optional string indicating the 'type' of the object. If not provided
   * uses the type name for the class.
   * @param parent_uid Optional string indicating the UID of the object's parent. If not provided
   * the method assumes there is no parent.
   * @param channel Optional string indicating an object channel. If not provided
   * the method assumes there is no channel.
   *
   * @return The requested object block description.
   */
   extern virtual function svt_pa_object_data get_pa_obj_data(string uid = "", string typ = "", string parent_uid = "", string channel = "" );

//-----------------------------------------------------------------------------------
/**
  * This method is used to set object_type for bus_activity when
  * bus_activity is getting started on the bus .
  * This method is used by pa writer class in generating XML/FSDB 
  */
  extern function void  set_pa_data(string typ = "" ,string channel  ="");
 
//-----------------------------------------------------------------------------------
  /**
  * This method is used to  delate  object_type for bus_activity when bus _activity 
  * ends on the bus .
  * This methid is used by pa writer class  in generating XML/FSDB 
  */
  extern function void clear_pa_data();
  
//------------------------------------------------------------------------------------
  /** This method is used in setting the unique identification id for the
  * objects of bus activity
  * This method returns  a  string which holds uid of bus activity object
  * This is used by pa writer class in generating XML/FSDB
  */
  extern virtual function string get_uid();

//------------------------------------------------------------------------------------
  /** Sets the configuration property */ 
  extern function void set_cfg(svt_axi_port_configuration cfg);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

`ifdef SVT_ACE5_ENABLE  
  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_write_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);

  /** Gets the current byte lane based on the current data beat, address
    * and burst size
    */ 
  extern function int get_curr_byte_lane_atomic_read_data(int log_base_2_data_width_in_bytes = -1, int beat_num = -1);
`endif
  /** 
    * Populates the partial data and byteen provided into data and byteen
    * that is used to write into a full cacheline
    */
  extern function void populate_partial_data_and_byteen (
                                                         input bit[7:0] data[],
                                                         input bit byteen[],
                                                         output bit[7:0] cache_data[],
                                                         output bit cache_byteen[]
      );

  /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane_for_data_user(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number */
  extern function void get_beat_addr_and_lane(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`ifdef SVT_ACE5_ENABLE
 /** Returns the address and lanes corresponding to the beat number for atomic compare read data*/
  extern function void get_beat_addr_and_lane_atomic_read_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
 /** Returns the address and lanes corresponding to the beat number for atomic compare write data*/
  extern function void get_beat_addr_and_lane_atomic_write_data(input int beat_num, 
                                              output [`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                                              output int lower_byte_lane,
                                              output int upper_byte_lane,
                                              input  bit use_tagged_addr=0);
`endif

  /** Gets the beat number corresponding to an address */
  extern function int get_beat_num_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr, 
                                                          bit use_tagged_addr = 0
                                          );

  /**
   * Returns a string (with no line feeds) that reports the essential contents
   * of the packet generally necessary to uniquely identify that packet.
   *
   * @param prefix (Optional: default = "") The string given in this argument
   * becomes the first item listed in the value returned. It is intended to be
   * used to identify the transactor (or other source) that requested this string.
   * This argument should be limited to 8 characters or less (to accommodate the
   * fixed column widths in the returned string). If more than 8 characters are
   * supplied, only the first 8 characters are used.
   * @param hdr_only (Optional: default = 0) If this argument is supplied, and
   * is '1', the function returns a 3-line table header string, which indicates
   * which packet data appears in the subsequent columns. If this argument is
   * '1', the <b>prefix</b> argument becomes the column label for the first header
   * column (still subject to the 8 character limit).
   */
`ifdef SVT_UVM_ENABLE_FGP
  (* uvm_fgp_lock = "psdisplay_short" *)
`endif
  extern virtual function string psdisplay_short( string prefix = "", bit hdr_only = 0);

  /** 
    * Limits the data to what can be transmitted if the address is
    * unaligned. If the address is unaligned, we need to take care 
    * that data[0] and wstrb[0] are consistent with what can actually 
    * be driven on the bus. 
    * For example, for a 64 bit bus, if the address is 0x7,
    * data can be sent only on 1 byte for the first beat.
    * For a FIXED burst the address is same for all beats, so this
    * operation needs to be done for all beats. For other bursts, only
    * the first address can be unaligned, other beats are aligned
    * addresses
    * @param data_only(Optional: default = 0) If this bit is set the 
    * operation is done only for data. 
    * @param beat_num(Optional: default = -1) Applicable for a FIXED burst.
    * When set to -1, masking is done for all beats, otherwise it is 
    * done only for the selected beat. 
    */
  extern function void mask_data_for_unaligned_addr(bit data_only = 0,int beat_num = -1);
  
  /**
    * Ensures that valid x,z,0,1 all four state datas are calculated with
    * respect to data_mask values. 
    * This function is called under SVT_MEM_LOGIC_DATA macro define only,
    * to make sure while masking valid x and z state data also considered
    * towards masked data.
    */ 
  extern function logic [`SVT_AXI_MAX_DATA_WIDTH - 1:0] mask_data_for_x_z_values (logic [`SVT_AXI_MAX_DATA_WIDTH -1:0] data, bit [`SVT_AXI_MAX_DATA_WIDTH - 1:0] data_mask);
  
  /**
    * Ensures that only valid lanes have wstrb asserted. In wysisyg format
    * the constraints leave data[] and wstrb[] open. This function is called in
    * post_randomize to make sure that wstrb is asserted only for valid lanes
    */ 
  extern function void get_wstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

`ifdef SVT_ACE5_ENABLE
    /**
    * Ensures that only valid lanes have tag_update asserted. In wysisyg format
    * the constraints leave tag[] and tag_update[] open. This function is called in
    * post_randomize to make sure that tag_update is asserted only for valid lanes
    */ 
  extern function void get_tag_update_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Returns the tag_update in the tag_update_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the tag_update is returned such that packed_tag_update[0] 
    * corresponds to the tag_update for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in tag_update_to_pack[] is directly
    * packed to packed_tag_update[]. 
    * @param tag_update_to_pack tag_update to be packed
    * @param packed_tag_update[] Output byte stream with packed tag_update
    */
  extern function void pack_tag_update_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update_to_pack[],
                                          output bit packed_tag_update[]
                                        ); 

  /**
    * Returns the tag in the tag_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either tag[] or cache_write_tag[]
    * fields of this class have been passed as arguments to tag_to_pack[] field.
    * In the case of WRAP bursts the tag is returned such that packed_tag[0] 
    * corresponds to the tag for the wrap boundary. 
    * In the case of INCR bursts, the tag as passed in tag_to_pack[] is directly
    * packed to packed_tag[]. 
    * @param tag_to_pack tag to be packed
    * @param packed_tag[] Output byte stream with packed tag
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_tag_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output logic[3:0] packed_tag[]
                                        ); 
`else
  extern function void pack_tag_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag_to_pack[],
                                          output bit[3:0] packed_tag[]
                                        );
`endif 
 
 
  /** Converts tag from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_right_justified_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from wysiwyg format to right justified format */
  extern function void convert_tag_update_to_right_justified_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);


  /** Converts tag from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_tag_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`else
  extern function void convert_tag_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAG_WIDTH-1:0] tag[]);
`endif


  /** Converts tag_update from right justified format to wysiwyg format */
  extern function void convert_tag_update_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_TAGUPDATE_WIDTH-1:0] tag_update[]);

  /**
    * Ensures that only valid lanes have chunkstrb asserted. In wysisyg format
    * the constraints leave data[] and rchunkstrb[] open. This function is called in
    * post_randomize to make sure that chunkstrb is asserted only for valid lanes
    */ 
  extern function void get_chunkstrb_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_CHUNK_STROBE_WIDTH -1:0] rchunkstrb[]);

`endif

 /**
    * Ensures that only valid lanes have poison asserted. In wysisyg format
    * the constraints leave data[] and poison[] open. This function is called in
    * post_randomize to make sure that poison[] is asserted only for valid lanes
    */ 
  extern function void get_poison_for_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

 /**
   * Simple utility used to convert string property value representation into its
   * equivalent 'bit [1023:0]' property value representation. Extended to support
   * encoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit encode_prop_val(string prop_name, string prop_val_string, ref bit [1023:0] prop_val,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);

  /**
   * Simple utility used to convert 'bit [1023:0]' property value representation
   * into its equivalent string property value representation. Extended to support
   * decoding of enum values.
   *
   * @param prop_name The name of the property being encoded.
   * @param prop_val_string The string describing the value to be encoded.
   * @param prop_val The bit vector encoding of prop_val_string.
   * @param typ Optional field type used to help in the encode effort.
   *
   * @return The enum value corresponding to the desc.
   */
  extern virtual function bit decode_prop_val(string prop_name, bit [1023:0] prop_val, ref string prop_val_string,
                                              input svt_pattern_data::type_enum typ = svt_pattern_data::UNDEF);


  /**
    * Returns the encoding for AWSNOOP/ARSNOOP/ACSNOOP based on the 
    * transaction type
    * @return The encoded value of AWSNOOP/ARSNOOP/ACSNOOP
    */
  extern function bit[`SVT_AXI_ACE_SNOOP_TYPE_WIDTH-1:0] get_encoded_snoop_val();

`ifdef SVT_ACE5_ENABLE
 
  /**
    * Returns the encoding for AWCMO based on the 
    * cmo_on_write_xact_type type
    * @return The encoded value of AWCMO
    */
  extern function bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] get_encoded_awcmo_val();

   /**
    * Decodes the given AWCMO value and returns the transaction type.
    * @param awcmo_val The value on AWCMO
    */
  extern function cmo_on_write_xact_type_enum get_decoded_awcmo_val(bit[`SVT_AXI_ACE_WCMO_WIDTH-1:0] awcmo_val);

  /**
   * Sets Combined Write and CMO type
   */
  extern function void set_combined_writecmo_transaction_type();
  
  /**
   * Indicates whether the current transaction is write cmo or not
   */
  extern function bit is_combined_writecmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_pcmo_xact();

  /**
   * Indicates whether the current transaction is write pcmo or not
   */
  extern function bit is_combined_write_non_pcmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl or writeuniquefull cmo or not
   */
  extern function bit is_combined_writeunique_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnp* cmo or not
   */
  extern function bit is_combined_writenosnp_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniquefull cmo or not
   */
  extern function bit is_combined_writeuniquefull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpfull cmo or not
   */
  extern function bit is_combined_writenosnpfull_cmo_xact();  

  /**
   * Indicates whether the current transaction is writeuniqueptl cmo or not
   */
  extern function bit is_combined_writeuniqueptl_cmo_xact();  

  /**
   * Indicates whether the current transaction is writenosnpptl cmo or not
   */
  extern function bit is_combined_writenosnpptl_cmo_xact();  

`endif

  /**
    * Decodes the given snoop value(ARSNOOP/ACSNOOP) and returns the transaction type.
    * This function can be used for the read address channel and the
    * snoop address channel. 
    * @param snoop_val The value on ARSNOOP/ACSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_read_snoop_val(bit[`SVT_AXI_ACE_RSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Decodes the given snoop value(AWSNOOP) and returns the transaction type.
    * This function can be used for the write address channel. 
    * @param snoop_val The value on AWSNOOP
    */
  extern function coherent_xact_type_enum get_decoded_write_snoop_val(bit[`SVT_AXI_ACE_WSNOOP_WIDTH-1:0] snoop_val);

  /**
    * Returns the channel on which a transaction will be transmitted
    * @return The channel (READ/WRITE) on which this transaction will
    * be transmitted.
    */
  extern function xact_type_enum get_transmitted_channel();
  /**
    * Indicates if this transaction is applicable for updates in
    * the FIFO rate control model 
    * @return Returns 1 if applicable, else returns 0 
    */
  extern function bit is_appplicable_for_fifo_rate_control();

  /**
    * Checks if the coherent transaction is DVM Sync 
    */
  extern function bit is_coherent_dvm_sync();
 
  /**
    * Returns the index (of data or wstrb fields) corresponding 
    * to the wrap boundary
    */ 
  extern function int get_wrap_boundary_idx();

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the index (of atomic_read_data) corresponding 
    * to the wrap boundary for Atomic compare transaction
    */ 
  extern function int get_wrap_boundary_idx_for_atomic_compare_read_data();

`endif

  /** returns lowest address of the transaction. For WRAP type of transaction
    * it indicates starting address after transaction statisfies WRAP condition
    * and wraps over to include lower addresses
    */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_wrap_boundary();

  /** returns burst size aligned address */
  extern function bit [`SVT_AXI_MAX_ADDR_WIDTH - 1:0] get_burst_boundary();

  /**
    * Returns the byte lanes on which data is driven for a given data width
    */
  extern function void get_byte_lanes_for_data_width(
                bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] beat_addr,
                int beat_num,
                int data_width_in_bytes,
                output int lower_byte_lane,
                output int upper_byte_lane
          );
  
  /**
    * Checks if the transaction crosses the 4kb boundary
    */
  extern function bit is_addr_4kb_boundary_cross();

  /**
    * Returns the data in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either data[] or cache_write_data[]
    * fields of this class have been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

`ifdef SVT_ACE5_ENABLE
  /**
    * Returns the data in the atomic_compare_read_data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that atomic_read_data[]
    * field of this class have been passed as arguments to atomic_compare_read_data_to_pack[] field.
    * In the case of WRAP bursts the data is returned such that packed_atomic_compare_read_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data as passed in atomic_compare_read_data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param atomic_compare_read_data_to_pack Data to be packed
    * @param packed_atomic_compare_read_data[] Output byte stream with packed data
    */

`ifdef SVT_MEM_LOGIC_DATA
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output logic[7:0] packed_atomic_compare_read_data_data[]
                                                             ); 
`else  
 extern function void pack_atomic_compare_read_data_to_byte_stream( 
                                                               input bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_compare_read_data_to_pack[],
                                                               output bit[7:0] packed_atomic_compare_read_data[]
                                                             ); 
`endif 

`endif 
  /**
    * Returns the data_user in the data_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that data_user[] 
    * has been passed as arguments to data_to_pack[] field.
    * In the case of WRAP bursts the data_user is returned such that packed_data[0] 
    * corresponds to the data for the wrap boundary. 
    * In the case of INCR bursts, the data_user as passed in data_to_pack[] is directly
    * packed to packed_data[]. 
    * @param data_to_pack Data to be packed
    * @param packed_data[] Output byte stream with packed data
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void pack_data_user_to_byte_stream(
                                          input logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output logic[7:0] packed_data[]
                                        ); 
`else
  extern function void pack_data_user_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data_to_pack[],
                                          output bit[7:0] packed_data[]
                                        );
`endif  

  /**
    * Returns the wstrb in the wstrb_to_pack[] field as a byte stream based on
    * the burst_type. 
    * In the case of WRAP bursts the wstrb is returned such that packed_wstrb[0] 
    * corresponds to the wstrb for the wrap boundary. 
    * In the case of INCR bursts, the wstrb as passed in wstrb_to_pack[] is directly
    * packed to packed_wstrb[]. 
    * @param wstrb_to_pack wstrb to be packed
    * @param packed_wstrb[] Output byte stream with packed wstrb
    */
  extern function void pack_wstrb_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb_to_pack[],
                                          output bit packed_wstrb[]
                                        ); 
   /**
    * Returns the poison in the poison_to_pack[] field as a byte stream based on
    * the burst_type. The assumption is that either poison[] or cache_write_poison[]
    * fields of this class have been passed as arguments to data_to_pack5[] field.
    * In the case of WRAP bursts the data is returned such that packed_poison[0] 
    * corresponds to the poison for the wrap boundary. 
    * In the case of INCR bursts, the poison as passed in poison_to_pack[] is directly
    * packed to packed_poison[]. 
    * @param poison_to_pack poison to be packed
    * @param packed_poison[] Output byte stream with packed poison
    */
  extern function void pack_poison_to_byte_stream(
                                          input bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison_to_pack[],
                                          output bit packed_poison[]
                                        ); 

  /**
    * Unpacks the data in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data is directly unpacked into unpacked_data
    * For a WRAP burst, the data is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif
  
  /**
    * Unpacks the data_user in data_to_unpack[] into utemp_datanpacked_data.
    * For an INCR burst, the data_user is directly unpacked into unpacked_data
    * For a WRAP burst, the data_user is unpacked such that unpacked_data[0] corresponds
    * to the starting address. The assumption here is that data_to_unpack[] has
    * a byte stream whose data_user starts from the address corresponding to the wrap
    * boundary
    * @param data_to_unpack The data to unpack.
    * @param unpacked_data The unpacked data.
    */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void unpack_byte_stream_to_data_user( 
                                            input logic[7:0] data_to_unpack[],
                                            output logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`else
  extern function void unpack_byte_stream_to_data_user( 
                                            input bit[7:0] data_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] unpacked_data[]
                                          ); 
`endif

  /**
    * Unpacks the wstrb in wstrb_to_unpack[] into unpacked_wstrb.
    * For an INCR burst, the wstrb is directly unpacked into unpacked_wstrb
    * For a WRAP burst, the wstrb is unpacked such that unpacked_wstrb[0] corresponds
    * to the starting address. The assumption here is that wstrb_to_unpack[] has
    * a byte stream whose wstrb starts from the address corresponding to the wrap
    * boundary
    * @param wstrb_to_unpack The wstrb to unpack.
    * @param unpacked_wstrb The unpacked wstrb.
    */
  extern function void unpack_byte_stream_to_wstrb( 
                                            input bit wstrb_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] unpacked_wstrb[]
                                          ); 
   /**
    * Unpacks the poison in poison_to_unpack[] into unpacked_poison.
    * For an INCR burst, the poison is directly unpacked into unpacked_poison
    * For a WRAP burst, the poison is unpacked such that unpacked_poison[0] corresponds
    * to the starting address. The assumption here is that poison_to_unpack[] has
    * a byte stream whose poison starts from the address corresponding to the wrap
    * boundary
    * @param poison_to_unpack The poison to unpack.
    * @param unpacked_poison The unpacked poison.
    */
  extern function void unpack_byte_stream_to_poison( 
                                            input bit poison_to_unpack[],
                                            output bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] unpacked_poison[]
                                          ); 
                     
  /**
   * Does a basic validation of this transaction object
   */
  extern virtual function bit do_is_valid (bit silent = 1, int kind = RELEVANT);

  /**
    * Sets the suspend_master_xact property
    */
  extern virtual function void suspend_xact();

  /**
    * Unsets the suspend_master_xact property
    */
  extern virtual function void resume_xact();

  /**
    * Gets the number of beats of data/resp to be sent.
    */
  extern function int get_burst_length(int ignore_exceptions = 0);

`ifdef SVT_ACE5_ENABLE
  /**
    * Gets the number of beats for atomic_read_data in Atomic compare transactions 
    */
   extern function int get_burst_length_for_atomic_compare_read_data(int ignore_exceptions =0);
`endif

  /**
    * Gets the burst_type of a transaction.
    */
  extern function burst_type_enum get_burst_type(int ignore_exceptions = 0);

  /**
    * Gets the burst_size of a transaction.
    */
  extern function burst_size_enum get_burst_size(int ignore_exceptions = 0); 

  /**
   * Gets the minimum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Minimum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_min_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
   * Gets the maximum byte address which is addressed by this transaction
   * 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Maximum byte address addressed by this transaction
   */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_max_byte_address(bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /** 
   * Checks if the given address range overlaps with the address range of this transaction
   * 
   * @param min_addr The minimum address of the address range be checked 
   * @param max_addr The maximum address of the address range be checked 
   * @param convert_to_global_addr Indicates if the min and max address of this
   * transaction must be translated to a global address  before checking for overlap
   * @param use_tagged_addr Indicates whether a tagged address is provided
   * @param convert_to_slave_addr Indicates whether the address should be converted to
   * a slave address
   * @param requester_name Name of the master component from which the transaction originated
   * @return Returns 1 if there is an address overlap, else returns 0.
   */
  extern function bit is_address_overlap(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] min_addr, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_addr, bit convert_to_global_addr = 0, bit use_tagged_addr = 0, bit convert_to_slave_addr = 0, string requester_name = "");

  /**
    * Returns the total number of bytes transferred in this transaction or beat number
    * svt_axi_port_configuration::get_byte_count_from_wstrb_enable set to 0,
    * the byte count is calculated using burst_length and burst_size based on
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * If svt_axi_port_configuration::get_byte_count_from_wstrb_enable
    * is set to 1, the byte count is calculated using wstrb based on 
    * @param beat_num Indicates the beat number for which the byte count is
    * to be calculated. If set to -1, the total number of bytes for the entire
    * transaction is calculated. 
    * @return The total number of bytes transferred in this transaction or beat number
    */
  extern virtual function int get_byte_count(int beat_num = -1);

  /** @cond PRIVATE */
  /** Converts data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif
`ifdef SVT_ACE5_ENABLE
  /** Converts atomic_read_data from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`else
  extern function void convert_atomic_compare_read_data_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] atomic_read_data[]);
`endif
`endif
  /** Converts data_user from wysiwyg format to right justified format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_right_justified_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstb from wysiwyg format to right justified format */
  extern function void convert_wstrb_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from wysiwyg format to right justified format */
  extern function void convert_poison_to_right_justified_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`else
  extern function void convert_data_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] data[]);
`endif

  /** Converts data from right justified format to wysiwyg format */
`ifdef SVT_MEM_LOGIC_DATA
  extern function void convert_data_user_to_wysiwyg_format(ref logic[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`else
  extern function void convert_data_user_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_USER_WIDTH-1:0] data[]);
`endif

  /** Converts wstrb from right justified format to wysiwyg format */
  extern function void convert_wstrb_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/8-1:0] wstrb[]);

  /** Converts poison from right justified format to wysiwyg format */
  extern function void convert_poison_to_wysiwyg_format(ref bit[`SVT_AXI_MAX_DATA_WIDTH/64-1:0] poison[]);

  /** Turns-off randomization for all AXI3/AXI4 parameters */
  extern virtual function void set_axi3_4_randmode(bit on_off=0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    * @param disable_msg_info Disables information regarding message format
    * @return The data as a string. If corresponding wstrb is 0, data is marked as 'xx'
    */
  extern virtual function string get_write_data_string(bit[7:0] xact_data[],bit xact_wstrb[],bit disable_msg_info = 0);

  /**
    * Returns the contents of data as a string. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    */
  extern virtual function string get_read_data_string(bit[7:0] xact_data[]);

  /**
    * Returns the contents of wstrb as a string. 
    * @param  xact_wstrb A bit stream array of the data which can be obtained through
    *              the pack_wstrb_to_byte_stream function
    */
  extern virtual function string get_wstrb_string(bit xact_wstrb[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  xact_wstrb A bit stream array of the wstrb which can be obtained through
    *              the pack_wstrb_to_byte_stream function. If xact_wstrb is 0,
                   corresponding xact_data is not compared 
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_write_data(bit[7:0] xact_data[],bit xact_wstrb[], bit[7:0] ref_data[]);

  /**
    * Compares the contents of two byte streams. 
    * @param  xact_data A byte stream array of the data which can be obtained through
    *              the pack_data_to_byte_stream function
    * @param  ref_data A byte stream array of the reference data to which xact_data must
                   be compared. 
    * @return Returns 1 if the comparison passed, else returns 0.
    */
  extern function bit compare_read_data(bit[7:0] xact_data[],bit[7:0] ref_data[]);

  /**
    * Gets a single response status based on rresp of each beat or bresp.
    * If it is an exclusive access, then this function returns an OKAY response
    * if all beats have a response of EXOKAY, otherwise it returns a SLVERR response
    * For normal transactions, this function returns OKAY only if all beats have
    * a response of OKAY
    * @return Returns the combined response status of all beats 
    */
  extern function resp_type_enum get_response_status();

  /** Returns first data_valid_assertion_time for read channel transaction or write
    * response assertion time for write channel transaction
    */
  extern function real get_response_assertion_time(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** Returns data_valid_assertion_time for the beat number of given address read channel transaction or write
    * response assertion time for write channel transaction.
    */
  extern function real get_response_assertion_time_of_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline, bit tagged_addr = 0, int mode=0);

  /** returns id considering only the bits which are used by exclusive monitor */
  extern function bit[`SVT_AXI_MAX_ID_WIDTH-1:0] excl_id(bit use_partial_id=1);

  /** returns address considering only the bits which are used by exclusive monitor.
    * However, if num_addr_bits_used_in_exclusive_monitor is set to -1 this indicates that, user wants
    * use specified start and end address ranges for each exclusive monitor. In this case,
    * this method will return exclusive monitor index with tagged address attribute i.e. secured/nonsecure
    * bit, as exclusive monitored address. This models the interconnect's behaviour of monitoring
    * different address chunks.
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] excl_addr(bit use_partial_addr=1, bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr=0);

  /** returns address aligned to cacheline size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] cacheline_addr(bit use_tagged_addr=0);

  /** returns address aligned to snoop data width size */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] snoop_aligned_addr();

  /** returns the status corresponding to the status mode value passed */
  extern function status_enum get_status(int status_mode);

  /** Outputs the expected snoop addresses. 
    * If the transaction does not generate a snoop, the function returns 0, else it returns 1.
    * However, if include_non_snooped_xacts is set, the function includes WRITEBACK, WRITECLEAN,
    * EVICT, WRITEEVICT and cache maintenance transactions sent to NON-SHAREABLE region as well.
    */
  extern function bit get_expected_snoop_addr(output bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] expected_snoop_addr[$], input bit use_tagged_addr=0, input bit include_non_snooped_xacts = 0, input int cache_line_size = -1);

  /** Returns 1 if this transaction type generates a snoop, else returns 0 */
  extern function bit has_snoop();

  /** Returns 1 if this transaction is a full cacheline access, else returns 0 */
  extern function bit is_cache_line_access();

  /** Sets the port kind to master or slave */
  extern function void set_port_kind(svt_axi_port_configuration::axi_port_kind_enum axi_port_kind);

  /** Returns address concatenated with tagged attributes which require indipendent address space.
    * for example, if secure access attribute is enabled bye setting num_enabled_tagged_addr_attributes[0] = 1
    * then this bit will be used to provide unique address spaces for secure and non-secure transactions.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Address that needs to be tagged when use_arg_addr is set to '1'
    * @param      use_cacheline_addr Indicates if returned address should be aligned to cache line size
    * @return              Returns address tagged with address attribute of corresponding port
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_tagged_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr = 0, bit use_cacheline_addr=0);

  /** @param  arg_addr Holds Address for which untagged part needs to be obtained
    * @return          Untagged part of Address "arg_addr" will be returned
    */
  extern function bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] get_untagged_addr(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Sets transaction attributes from tagged address.
    * for example, if secure access attribute is enabled then security attribute of current transation can be set from the tagged address
    * passed through argument or current transaction address.
    *
    * @param  use_arg_addr Indicates that address passed through argument "arg_addr" will be used instead of 
    *                      transaction address "addr", when set to '1'. If set to '0' then transaction address
    *                      "this.addr" will be used for tagging.
    * @param      arg_addr Tagged Address from which current transacion attributes need to be set.
    */
 extern task set_tag_from_addr(bit use_arg_addr=0, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] arg_addr);

  /** Function that sets xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set */
  extern function void set_xact_type();

  /** Function returns xact_type as COHERENT if svt_axi_port_configuration::is_downstream_coherent is set 
    * If not set xact_type will not be changed for the particular transaction.
    */
  extern function xact_type_enum get_xact_type();

`ifdef SVT_ACE5_ENABLE
  /** Sets the atomic transaction type */
  extern function void set_atomic_transaction_type();

 /**
    * Returns the encoding for AWATOP based on the 
    * transaction type
    * @return The encoded value of AWATOP
    */
  extern function bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] get_encoded_atomicop_val();

 /**
    * Returns the decoding  for AWATOP based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function atomic_xact_op_type_enum get_decoded_atomicop_val(bit[`SVT_ACE5_ATOMIC_TYPE_WIDTH-1:0] awatop_val);

 /**
    * Returns the decoding  for Endianness based on the 
    * transaction type
    * @return The decoded value of AWATOP
    */
  extern function endian_enum get_decoded_endianness_val(bit endian_val);

  /** Returns the inbound data size for atomic transaction */
  extern function int get_atomic_transaction_inbound_data_size_in_bytes();
  
  extern function bit is_addr_aligned_to_total_outbound_data();

 /** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] get_masked_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[], bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb[]);
  
/** Returns the masked atomicop data based on current atomic xact data_size, input args data and byte_enable */
  extern function void get_masked_atomic_read_data(bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_read_data[],output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data);

  /** Returns the masked atomicop wstrb and  data based on current atomic xact data_size */
  extern function bit [(`SVT_AXI_WSTRB_WIDTH-1):0] get_masked_wstrb(bit [(`SVT_AXI_WSTRB_WIDTH-1):0] wstrb_);

  /** Performs atomic operation at beat level */
  extern function bit perform_atomic_operation(input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] masked_atomic_read_data, 
                                                input bit[(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],
                                                input bit [`SVT_AXI_WSTRB_WIDTH-1:0] wstrb[],
                                                output bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] atomic_resultant_data_
                                                );

 
/** Unpacks data into atomic_swap_data and atomic_compare_data field. This is applicable for ATOMIC_COMPARE transactions only */
   extern function void unpack_data_into_atomic_swap_and_atomic_compare_data(input bit [(`SVT_AXI_MAX_DATA_WIDTH-1):0] data[],int beat_num);


 /** Unpacks atomic_resultant_data into beat_format to do the beat formation */
  extern function void unpack_atomic_resultant_data_into_beat_format (input bit[(`SVT_AXI_MAX_DATA_WIDTH -1):0] atomic_resultant_data_);


/** Performs Atomic xact operation such as ADD etc. */
  extern function void perform_atomic_xact_operation(svt_axi_transaction xact);


 /** unpacks wstrb into atomic_swap_wstrb and atomic_compare_wstrb into field. This is applicable for ATOMIC_COMPARE transactions only */
  extern function void unpack_wstrb_into_atomic_swap_and_atomic_compare_wstrb(input bit [(`SVT_AXI_MAX_DATA_WIDTH/8-1):0] wstrb[],int beat_num);

`endif
  /**
    * Indicates if this transaction has poison for any 64-bit chunk 
    * @return Returns 1 if poison is present, else returns 0
    */
  extern function bit has_poison();

  /** Marks current transaction as part of multipart dvm sequence to avoid irrelevant
    * check being performed on this transaction.
    * Since only first transaction of multipart dvm transaction sequence has control information on LSB[15:0] bits,
    * it is important to set this bit to '1', before randomizing the second or later transaction object so that, 
    * second or later part of multipart dvm sequence can ignore dvm address constraints for control fields.
    */
  extern virtual task set_multipart_dvm_flag (string kind = "");

  /** returns first beat of coherent response of current transacton */
  extern virtual function coherent_resp_type_enum get_coh_resp();

  /** returns '1' if current transaction matches expected transaction type i.e. for coherent transaction
    * if it has matched coherent_xact_type and for non_coherent transaction if it matched xact_type, otherwise it returns '0'
    */
  extern virtual function bit is_type_matched(int rw_type = -1, string typ = "non_dvm_non_barrier");

  /** returns '1' if current transaction will allocate a cacheline but, there are at least one transaction currently active
    *             which will attempt to de-allocate the same cacheline.
    * returns '0' otherwise.
    */
  extern virtual function bit has_overlapped_dealloc_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns '1' if overlapped transaction between read and write channel found else '0' */
  extern virtual function bit has_overlapped_rd_wr_xact(int mode=0, svt_axi_transaction ext_xact=null);

  /** returns calculated parity value for 8bit of data */
  extern virtual function bit parity_bit_from_8bit_data(bit [7:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_16bit_data(bit [15:0] data, bit even_odd_parity = 1);
  extern virtual function bit parity_bit_from_1bit_data(bit data, bit even_odd_parity = 1);
  extern virtual function void parity_for_xact_field(input string xact_signal_name = "", input bit even_odd_parity = 1);

  /** returns calculated data check parity value to data */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/8)-1:0] calculate_parity(bit [`SVT_AXI_MAX_DATA_WIDTH-1:0] data);

 /** returns converted  data check to pison value */
  extern virtual function bit [(`SVT_AXI_MAX_DATA_WIDTH/64)-1:0]convert_datacheck_to_poison(bit [`SVT_AXI_MAX_DATA_WIDTH/8-1:0] is_datachk_passed,bit [`SVT_AXI_MAX_DATA_WIDTH/64-1:0]data_chk_to_poison);

  /** returns '1' if transaction passed through argument i.e. overlapped_xact is found active while
    * current transaction is found active or in other words both are found active at the same time */
  extern virtual function bit is_overlapped_in_time(svt_axi_transaction overlapped_xact);

  /** returns '1' if current transaction will allocate a cacheline else returns '0' */
  extern virtual function bit is_alloc_xact();

  /** returns '1' if current transaction will de-allocate a cacheline else returns '0' */
  extern virtual function bit is_dealloc_xact();

  /** updates num_xacts_blocked_progress_of_curr_xact with number of xacts that blocked progress of current xact */
  extern virtual task update_num_xacts_blocked_progress_of_curr_xact(int num_blocked_xacts=1, int mode=0);

  /** returns '1' if current transaction is not supposed to return data as part of coherent read response */
  extern virtual function bit is_read_response_without_data(int mode=0);

  /** returns '1' if current transaction will allocate a cacheline in L3 else returns '0' */
  extern virtual function bit is_l3_allocate(bit is_exclusive=0, bit is_partial_data=1);

  /** returns '1' if current transaction will de-allocate a cacheline from L3 else returns '0' */
  extern virtual function bit is_l3_deallocate(bit is_partial_data=1);

  /** returns '1' if current transaction is supposed to update memory with L3 data */
  extern virtual function bit is_l3_update_to_mem(bit is_partial_data=1);

  /** returns '1' if current transaction doesn't cover full cacheline */
  extern virtual function bit is_partial_cacheline_data();

  /** Returns number of byte whose wstrb is '1' */
  extern virtual function int get_valid_byte_count();

  /** returns '1' if current transaction is determined to be valid exclusive type */
  extern virtual function bit is_exclusive_access(string mode="", bit shared=1);

  /** Sets the channel on which a transaction will be transmitted */
  extern function void set_transmitted_channel();

  /** Returns '1' if write strobes are driven correctly otherwise, returns '0' */
  extern virtual function bit check_wstrb(bit silent=0);
  /** @endcond */

`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_axi_transaction)
`endif
endclass
/**
Transaction Class Macros definition  and utility methods definition
*/

 `protected
(&DVQEQQe-?\f,]Wd96S#@@=BE(>O8-4AR5?+gdJ.ZH([d1_I/+J0)#a2Y2.^BJF
[.<U\6Z>YgHA2+07X1=30?##FGU).:_MOR>7K_bQJ=II/G5@S4WS.>L2Z1T,NIFU
K1QY,7/KfCeeLMMIRaF)T_H)VJcGQYC]6Pe2QU<DAdZ,+<]?&DV54LH<6UL(ZQ(\
cbR>(KJI800NOM7[VF?K0L&8II0EC7CYA+=1+N9>\;SdP?[,R+RdVcHZF(_0_S-b
INeXF2aAgES47fA?=ZQ/>J(^f2:>\F37KO2bQZM2KI+WKB^T<DeB0E]B&7:YC<8)
XAWNG?+Fb?7KC_YSB>,YAT01NOb6F14C4/J<=L&_GQAK\.#.=H?Y\J(HKG^c=A/g
3&R=73Z5?cDaST8\Bc.Ne/YOA+?[^K+dE;O-T23D#dE.^?>RK;X[TD.KKeY8WSBb
T2WUJ=(M<e()P:F0VAK:=;bF/AfSX)\d<gWc2<STR.TX(:?-Q#N9=;TU=e^5)4;e
KH:L#Q-af)U/#Fd-K0]<^:Q@N#,Xa-_MW#^M8b+BPC&TaW92)).)U9;WH0gSUR.<
[OE[<JTb[a.]5SK3]/7Xfg^<V<;S/FM./,RNIbgN4M+)9CA.#8#cX7gD?5W>/Z@8
KZ:.?DYcaXV5@)U>K#?FcH?LaI@4YZD2N2=9LF_W;(R9TFb>bReF]L/Gg,W,4Y#f
NAgMD@2GMUDB^18W2Re_\.Vg-[L;ae_cSWWU5@7R&[895&.N<RFO(IL/Sd/E_OR]
e@&cCV:=fJ0P[8&)1d]IN/6-bNBaSIN9Y:L./7f3WB6FS1Z#:82fc+V+;/@.XC0:
PTO2VO:B3AZN4<P=I1MF@Y)#;.a=5V7DDW/Z/ZU9WcXWPfVF8\-D__g[La]Q6QQB
[9_WeEJZF^55L0gBH?bV;33eHI#H9WEbSf+d@?/>\M6M9(dBPb2)W[4]E^Q#_5Gd
MJ)D2A@:?Za5AV.VNc<Fe\dJHFU9;4;Q1c#&XD6Ud,\6AX0?7DFSX-D6c?De]dg=
PcPH>X4H9Y>E.I9-U8V]0VC27BS;=I,OUG8cH?#0BW-^-6<@B2b&?YTJ/4G-^(]@
V_S5NA=M@OWKe#A0ggG;BXeY-#)0<RYRed:S/gGK&=SETG:7R.M.OD(cW>2:0Y0W
L1.K#eWIO7FPC94C_\\6]#0)?g,ZT];DM=##FCZ8X#<fL#]RSe[G<8_C;K?S,CNZ
/_TOE).5S=/@F;fB.:GNDCgW?86E8FHa9V_D,OVTe+#,C=JF9HbNe&?02R:GL>D@
.5^2gL]9YT^[RH8N>)TRACA\D_&A(E66D?B6IN:fc3gY][_7]ea.b]CV+bgU9B,e
ZFf@Yg-CgYd.a&9ef#D47FS8Rb43eGHL-[ETJQ1WEWXWfJKf-Xg\0&Oe=3I@(,6V
^TFLcZEeBT8N5gW5)g2^6FcHg]5a507?b[d&SMag/7g6dGf0<VDL+JgR#A,B4=V[
3CGePIM>f2+@e1D8VcaY@bTb@[QB,.HK+QW72]bR-@f<P&#930<3\DF/UI[D-^Q=
Z#?(O:1^9dYfbG2NK5-Q3<;0g98OD2g5D?OI>5Ba@^1cEU4QeDTGS[S;_fSMIGeW
(@?X@KI]]AW/0@NY:[@(;H\1^d5:BD[I5:<4ED79;TO>5&I3]f?:=P_@SOB<ScS5
?cB-RdPL8I4==N3X8^905FMNS<ACKLab1T]Sf=df4BP/c/,CdEZT<:E.CL0c0?ET
)B65_^U];cWN,5DV\2A:P[S-?fDR>f6[eBg;X9N:/4c7=I8#:?C)S^S6Y0XM606+
DS3?5&8Cg[4=P0NUgJ0/WBOK9SfW)C/<J6;RcK@.f#P@ZNZ/X7A9Y992-#eN\#J(
QSYKS94fc0VQ9^=1OM=3PP^M(0S<@FJ<#X53&fd+NQAKGX5gQaRf]NQ_UJSbZ/Md
W/;K<]21ZTe2XLOZ@BP&SG)G_IFFKCAIGIGe3(#SK+]]=MA&N2K&I(DQgE,NM1DM
#3c+@XWC9H;9aADad9.2IK6fcQ#<QEKcFO[gBF1PYVdS)\(AJIeU@E17+aKfL1=@
A];b2A0Y>&:.D2GdSCS8+Q>([_<JA2[3M#g=8GfC@@DCF,&=fYK?d.F@AD&Y/SfW
FIUgbXUO37c9d9)d=S[#@N(HbdH<GO]Q2.2/AC#@?G_J-;a.EV=e095NgBD?(?bE
cF&N_HP.^5\6f7-W(a(&Ia:^6DR@B?H1X\1W,>[V^GS^^\/RIK0XF3(#,[>L^4.Y
@@CE&d6&\(L78@(dWcAfX0>:Z2>Sc#54\_R@D2/CW[Wd<(=(gEQ6S_TE];UH2)K,
NB9-5L)5S2Y5)@^\(^_H/DP<\03Y[0GZZ\/eA@M-4X79#,F/>/80^_[f523@1DU.
&A@fgFGHHg(E\#FH9SMXJ)4<]I2,@gX+=V=JJ;^0.9?W(<+A9LacWPB.JeG),;a#
O\deJA=Sb6&V28(XC/:LLW@D:&f0=.&T6][&WaE5bGCTG22UT@+<]Qa=a]@K+7E1
&NF\W7M/2BA/:.7C/ZbLa?IT3dcHgTL6g87G7ZY4M3K=Qd;A5Y7;R&(7>Md=1X3C
PJS:a2=JEX?VW<e8/;K-/_bZOVS;UT_H6\JOGNK#XF:)9d-4&^cAC\XBgcgd>[.E
N\;E:1:;Y::43MA<Z-R#?6,<FHWfW7UL3WQ[f:F6+^3Y&XIa:(2<5b?<CfURH]09
I@S@BAQ]DO-E4d>76J]T4gBEN#/fKI1?1-YEbG-_gQ38OUe.#=W1@D8YF7(5IfY8
S6<d94G-+,cd]SK/AC?SX[E?/Le?VG[=>E]LHTa;PA1MLeYG?C/[8P@9N0>cS=I=
JTQQ+6-5/B?_4.6\M15d--dF2OCdOagI<:<=XT.Jb-Ga(D=;<CbcYI(8&?R?B.&b
?fDZ,Mb<E^WLQZ/WM#\-I1BLX2c8>1)3cbNF187_ARNBX[1XTJ@R..,NVX>SCYC1
^UE[0C=a2F;0T]HR=59D<Sg\/OGeKVLU]1?J509I-5T2NQ>[A7IEWQ6ce]W7>\56
0[H#/??Yb,U1P?XBcNR5Ke-5U;FYAFP56,5I;JNCTI/Ba+<AN5^#>G?6_e:>ceWK
U<b&UW&_cKFZg8X8@c=4@+H\geBNOGM3#F:0UQYZI.DTf6J\^HaN,VS7P/7E=+C6
UfG-Ca&PGb;LH:0>3J5Z[K=]ZHaH==R2,bMFX#R3_D0Fb)G,P.WF3_A+6(A0]P=1
E>8GTE+9K[7eg5?\Rg5Z#II4<(T0U,MO7g.b=J]-K?[-F>[^&O9CaXc6<8;db8(K
dg+(6QcVMB;dd)97GH6+[2Wg8T,=_8RS_8aC;I2RUEZA2+4](IJJ@7Ka(Tg4WH?g
TQ)>>07dg8GAT,[^S>Y5cRd^X(-5_O(:ZGPKeWR6g]?W,>_4Z^fG<I,JQ&&@+V<3
SF2&X8d51^D=R\;;G&P)G.())1K:QE#XB2J.S?YTB;@21G56eBb#E4G9+Z8.a?48
&5gXM2cT9//VZ2.)1D#OcKNW_9M5VRF1QR5CUGK[MUWK3C)>Vd@]4e/]_IJNgFDT
)M[bCZ#c-6TBELL/1V,QOG9A1&AAf0I4>[Zg6N-WK5d7\\gg\\g\^2c6R6]JYQYX
=PUPCea/_U^Ed1XN<L=R3-dUS+TSdCQ/g4G#GA[BTG+/aZ>]FD^>CS]M_+;c>X7Z
JSPT1P1/+TT5IQ65]NaC5cQ+-a6d/6)UaYX:BCVF4&A5eTMHR48H3M,\g730Q=.b
L?E_=<Dg2XMOW)LX]F#bNa5;/_CTYJ4QOKU6B-A3AI[,V<=bFHd8F)a37fRL]cS-
SfR&0dB)3KB52_:#NCJW\He5]2[L>^=V/0dXbbZOI)XbB(XB.[<,)QDF9P5&+J/a
Y1Cg9XJEX=20QQ<#eB/]OMNLO-,BF(VXM8K=QFQ;aA5dIF+N]I#eOKXL32CCL(IP
?Q6+SV&2e;T_dLe(&3DPN#C,V77F@860LO=.ffW#L8HgNWKM1<4QX+/;<5H[26_I
OTfTLVI]4Dg0&P6NL4bc@&YWR0cF)OW0fZ.E<+OV0a35VKOe9ZQBC97L\]fBOVeQ
7E9X]eZgR#e>#^J5R^9U[B>F\CSDR)OE9RPaG.EW8W,UI=REEb,9_#0HeHW:?eTI
/>d,LcIg]f\LV&&^,.\3DA-&NMRSc)EG8bD8GN\XE^QTVMF\;HM^RdKNYeE(I^G-
ZA+3(FPTba^CT0H)[RLU73/Eb:]C1gP1^dL;OL0IZ<B9b8]BL3>U7IdJC4K5AL8N
Zd8/_@+)WKAIA<4[A@]/c;JV,NE<FM-,g[38YXS&@<RU0OPgV&d>PY:8f\4/7Hf?
[gR8bICgc8-6+L69>-dEA&/R7NN/)/Hd38[1S,B#X;0UH$
`endprotected


function void svt_axi_transaction::pre_randomize ();
`protected
Mc^@JYL.-:MXVP_S02QOIaK91PW-[RYeTJI/)QcQF.1>8^A)T3]<2)PMaHY6O/RW
O[2&/#=6X))@KVE&+UFWFb&U7@(\6:8CNbfD@2WCEVd77\4g#La;,QM;\[MK(A/-
O2CT79Sf>PXW-[Pa6W^dZFPa(dW_6YGZX;?c:gG<Y3Pb7/g(,SdUVg6Q2Oc]5c,C
;d^A&Qbf20)0&[4./f&83NW3gKW>#QR6d\>L7Z(AR5Y2P7KUGaYIdO@S)&-C]Nd3
OcgT]9a0c0d]LbZ+7KfU];bRdfP,A>QVLH-HTFe:7+FRR^(a#&9FOS)4(XAAW?C)
\V2Q<7Q5SC>8,OZb+3O8AXC\<\,[S)5+]S7LI)8VV\,??eEA,1RW2)G#b=B83a:8
b/X52-G0OP;)0L[9W<61@1;5\K#E>V#dYQE@9BYg6B.,=UDdKI@+f)[RgG9-3-74
L^LZ/X,X6XG]IXO53/=X-WK<efUdPQ]?2CA5\<[Lb.=b=YY><:5;&OQ1MJ]CFf<H
1ZAEL+R-S/Ng0Z@[Ya9SbaI9aY<\[4dWIARMLLB8g^OS7712IVYg5D5g28X(G?#N
NBO23#I&@;>e:S\63KK\5_1Q7\5Q/bZU[:N2_a&0[Q/9_-2YDQ2=;MbXOOM5T32D
V5bH,NdQ40Q4YEJ97J_GQ5X?BFD>>OGgM5V=1MIUM?Rc#>Hef/BL/R0CgWFU7^+S
:#RPI/[@P5fFV:#8(OHSH/61B2f?_e24a.NLe3:F_ZTKUZF#=,BP,a4JA7T[;YdF
;K841V<EFX_YT5^;J47_R@T=;)9[G7DZ)QS4e&5d=OF&^0+<Je&6)TN4fH+OJ@:G
P=8UDJ8[c;/DCGb&_N#TSZ8EFf1-@2XaT2ETKHONe[DK83ZV>_];e(U:[cF/B@AL
-3CV[g[SWO-]//K8KJ:P<6NZ&.VE30&&d6?6Yg@7AFc^N]2^>_CR>c6^XHNHDgUJ
BYCL@T=D-A+#F<5@A/EV9eRJQ>V+?-+^C)c02>@GYN6THUbL61(B(3b;\Q#^78IK
^S,4=NU)?DV,WUDgLg?-UCZ)A9J0<fAT+C:?99<12QUT0O>M?\VTgd)cY^E+8JfX
Z63RWF,B8NNAN5,0g12(VP6\feVc=DAW&SA0c2W^178T\_U+J8&UU10@cVYPI>-2
U&WJgc?>=d3P3:593)T.#:WeC@LAWMaGBH6C#Z5NY<>ITK>b7)WY(_L1_U1aAG^c
SFdK]G6@I37=8Je5WS=Sde)DPZ@SaGWbS5[0TJJ2O+O-&fN1gL__aU4TE0=,=S]?
+^06K@2VW3N9RC:M/#Hg?HYH/]g[]3)f,g,4)XQWb&WVB_K[1^.=c[Y^BR6VUHH;
#3da)_[KDN;fZR8K?g8@GV_)bR8KM+)0NYKE7cX+K:7gI)fG@e/)E03]R2b&bE6)
_-SU,:-GS.-_DdMO#)L#6=QXQOTXPbPW31KY^K?fGW>Ma9-;EA#[BS6/K4H5>-7<
_c(17a1DU\8RG-]<TM^Q5>_Yd@#G26Id]]A>eO#B<2d#f>TGP;LX6/&I9J/V;]-T
g0&4bDJF;S+2e&6d6b>[AX?OL\bQ,JCM#3f,f&7/D?[c.GGCfcUK>0<aC<?6S&,6
]_TU.[NGFRMbQD_66X((K2LcOF1_gSX#4TU7)/X+&8A112BXddS3MXCOF&,?)R\P
_+S.+P;aQR#UMfL10V(1+(><]IAPUAFeQdD136^b;/fV7?)N;3B2&SMTU+M3+EX,
74X]4SZS9A+X[gA]ZN.)1;bO86=JO\O<__CT/Y@-PO,:&E#\5E>]YQ_[NR6@LT+4
2A7(M\GcT7[0(WWEf19d4&:KGS;C;#TVX/d?X\N>;NG+7=>d)\1Z2N?_&BI[RZ\d
a.0MKDL@&Y\fSV_X37S<HL+=3O\\FafEgS(+&@;Y2c#TUK5;a4TGEQM7@E72WQF&
U4<O:ECUR^8/c7,AGf#cCeR1_L26O7e+1K>(aX)7>a?Zb><cE#171D[-:1Mb<_#5
^NXO^beH_D0ePPC^XE9PHO,2W&0=WRV4,O4]7/FXe0#-eJ4(VZZ<OIZfe&@:&1JE
?65ae97C7ID\AgQOKM\?VR5Nf=LT0N;8(4T30VdO^+c(+TD+-L8#@X<X],P_W11)
EY#91U4V7b[(@0f&^Pg[GRIe;Bd_W<^Z[0W6I1>LKROc8PFH7JB5Z2a0Q#MVZ<N1
-M:-01/\/Fe(BX[bV6ef[_K,-M\#S=Cg<Xf&B0<@:I;Y#GN7OH-HFC6>IK4+RPMJ
??G6^M<D2C.KX3+cc2e6KOTD#X<4G#>\E_[40VMeZG(G<g:B3J@3#.f0LC4]9UG5
,Rebfa6WB(TA+8U5Ud/_LU?0#<W]PN>Ee/[?>@H#@CO?D[efO2b]?U<gS+4L&QII
EF?22fZ7S/\2W&B\O]N.;G0_Z6MWfLW.;>QD^7H^.?9D,=1/9V?.ae@B4[Q/IU.Z
[5A5S.#WbLNLEQc=\F#1eJIXJD1cL8YVZUD+dKbNAgJbI4&(gJBIM>MT&2=1ITK5
V^:Aa4GaC=:Ec9aeLI>3ZJW-E:5=8)\b>1H=,)BHfHg<GJ-ae^/,G4I+Hb45U(\X
@=6<TAg/-[1^:4;1N=PZZ6gYX>4EMK7R/E(N/7g)1N@_ScZ7/@OBOcHcgFO4S(f2
FI\TUE4M2_N]&Yd192e,\/SC(/MD?>EE)1#@NJ]0#B:KDfKP-+[02d9b1YUS.NVQ
18NR_&7b[5.GOHaJ[Ab=eKg=Y[+[0^A++FLN6))S\E-cWYOD&KVL2aRK8_2gIQJ0
d]eTP>OXX,^A+9Q#8:b;U1Ef0(0<66HD\[VYg0TH0;LMV&>T@D).&ND[XDV<VC-^
-A3-D;8g0gS<JY^6WIc-O^93LVf]C&LE22OGW_HMTf)8UCgO)fMR[VDVGc=Ub22C
X(8D+UMHE7^H9YETUEYOJf,eJ9F3N_[Z8BD8Yg/I)XT@R9CPE<;#DJZ4J)&0WX]3
@G,\T3?^cK+.HVe>62.Z:LTI\.JB^N(LMcHe5?,3gaTFUL+C,#LQFR#O1[T8g#C3
>[(G<TURQ3gUQJ\ZPL&9X:<]Ra&/L?=-d.8^]L[5Qa;B/.A]LC0AKVSf53R7/\^M
D7&8+a<a=X6BOYAJ>eUEEdeVdac42(HH^^4+]ZUaaA8/f0SVH0YD&<Wb(UJ[7]&g
PggNMU8?c#PVI=Vd3F3&.C5^H=b44]R1B&81WO.fcA-)J:_L84cD7/9\RR0ZeP:[
NO+cWGJ^bEX.ERPd._:W:B0VV>UG:3Ee0a@,?V3A0I^7[B:I,D)Yg2gI,Cc?:c[G
dV3dUbS,O\JD(S7FZ=K52AUVP@UYFVKGg;,La\J\)N/ObN)74fH9US:><A?.UXQV
QP-+J=bORN7XR.&ZFX:S]LXONYWKGGB+JC@MS+\Me6739+@gO-<0ME,[]YaQ=3\:
4V5&fE6KK5-HZ#eHXEdQFGLF\U#<>8e+,IeZb.7b7XK1BZcRA[5(>));Nc-@23e;
/+4VX;d94GC/JMcd:WL2:8c78UH78B(E9/@==TA=;FV7b3BV^X&dcF.E?2/Jf[T=
dBK3J?O9_=3+Q72\W154BDf@79@V=52>D8KdNGXT^g>ZJgOdRCDP-T2_UYBK234X
D?=Q#N#Ycd.>J[B=+\]BB>]&FQIYT5KKS)6_IQSE_ZcC7=S;eGf8T7e.<OU>gD7+
UKX=S,B<]^HSSTRD7#JL,cZ/6UU>)TNe28K\g6_#H5gQbMdgNAa4Ne;H\J\P,+Fa
(aJ>A<J)0R[1&^/8^fSD+Y+^T>7B^L^Z_>&.#)e\b(^RG:UNBUD]>5c;b^J5X:PZ
JS=XJfFdGe,F-+27#U#RIgR)TZfdZ0gaK?I84D0Rd[a[SbX1,ZD((VW(LO5/OaE&
OC#W1QF?TJaQ[EBAE\)Y;e-GLgG)41WE5.:)f@TX]7D4;g+9C#S3NT5CS5@;<cG\
@ATM>#@41d<gO=4Q5Z]R@gYPb0Zg&R@1Kf]55R,\2.@BH^:+F3U8bVW;42I^WLV,
FBXBFcX<=WU-<VCggC]-0g_+D@MNB;Hga;7<OTe<3d-[ZIP<FCgCLBN&]QX1g\(6
2^,5+DS^@>UGIG:)>4S,>M<)RSKE5SWN<3_GLRI6#64.=5RL_gALH(P46E46gO2.
S8&0E.@e98E1Jf4JgL7A5b+E,ZbKKfVNf0UXeL\f?.+G?==L1#V[cG(0++Kc)2WT
UFZ_8SADW-1MfS3T25BQ?451@QVQH7>RFL3XaeEWJZ;.?.]QT<=1f24@L<04F_7K
I?PD)aaa,\DH?(?G--71>81D0]VX4Ue9Cf_:]ZQcH,6#[P_.._/@RdU1^GKJU74b
C)-#=2g^),2<TbY-O?aX6^9Vb&ANg(,+f[5N(bN\QI1Ccc,fITE(g,)Lg#C62+FE
3A96@\XAMb8g/)17e,OfR<+O6XQ:W\bK_<@DN?(92a(;+=C+OeSab1I1:6GfI,^7
>AB_I8:d7,cIO/WcJDFENYadQ6I[RKHR):59S2SL=U0-fY;1fJ)2DA]6MG#LaFCB
/>\.>J+8fTH:.-F@[+BG:Y9Y_N1D&GcXNPUSM3J&_=S?7&N#Q?bX\..DR66&?^ef
7Z;VSS\;[c@8G_4@1aER?HC4VJ)<Ib]N?[/ZX.-GZ_,BI#?]&[B(7VYD72a-EJ8/
\O8H,[?8R0+fE5&9b?0(L^L^P/ZbeT=+[>Y49CG46WOK.Kf)<aZIKfeUA/P9XbYQ
N@[gPPU=(f.4CF&=90TYIVE/>T(7;W@OOR\\#fABZTV?8FQ7^Pb,04M72=/5.Qg_
J;#e=b6U\Q&#?7_J?F@VIfY+F9V&]QT@cFg5D@FR,Ccc=YB\d,]Y/0OXO&_,8K+9
eX:]AYg-X]13Y0Bd]bb)gR><:0a47QR<ZWVHHL1Pd)DMBL&_E):AGIN(F/BB.4U@
c5W\\_6LVg0DMb7?,LLXE.1A&=)\cI)^^gQD6(SP-8(TU8G25I(D<^.UbM>EMc\L
L:gH:dR?=>()T=S?=N/).Me#E\[g7#UTY7K60[J:&d-AgDX[9&J5B#1Q\7d#W?>N
^-=JNKfDH]&C5P#2R-:F/4_(dFKOJJQ9621:>Yg5\O[8;53.?CFfERYZI-Q./>,B
+2P-X;V(g;^HRd:ZX7@@GcgOED,,S(@3HXAJ=X</U>OU,,7S6XK86A8#L3O\(eIF
1/WB;=&G,W<d4+8QN1gf1S/7-6?.JB/@>DaT>9?MY?)BG[V@PJH@6A(SWT_ZcW6.
f0NTPgcTQ_S30?CC\P(ad[2[IX3\BV\)]fR3Xa([M?,?,)Q7=b,YJ3Bc)aZWSBA8
/T#UcIH#P,,B&8L6Pa[91IV,.J+bdgNQUT-WB.2^I^g>_1f1<PL[L,Jd0)3@C4KU
fW=E_9W@ETVIIO]C=Zc/T0[@WUS4U:(ZUSA6ATY4U1\3N)A.9+[B3SLfG_=f>dJ_
N:>^C6/,69^Y4[eKffcXcQdU7MH3GbMKOb?H>(U^OP6G+G;aP/7JE_C]NBc889>b
6?c#O,L7,XQNPC2,M(FNbU?a4>)@U^N&(.BK.Q;QKgRN34S._VL4,<.?9G3;BR5b
Y>(Ked(&J2/Z1UL.GG0U=?DBM?PIBU;&[.Q9=b8C)?#>XV+,_^+g9NF5<6I;3KcT
=(52H&Ye4SJc0)L/[<N(fM7KM)e:Oda,BPa=H-?bLIHO/VX0=dJ-daWPW(#7_Y@:
Eb#c-6N5fb;T-S?RH_,&fRM:ZA+]@]WT)6P[FM)5FG26cb=<fAHTcfJXJ<=M)2U=
/CZMZ]?2MfMa13HL5g/R.J]O=DdSKW.c5J)S69+X737XFE0,:@=/21F7T9L.50].
#/H#7XW#L2Oa;7_+YKaGOa=YB:P^?aZKg<4+acGTLE&fcIL&)&;ag&1P.OM4&9MM
dT+)<BT6\1&\>0)^/ZS>]e6(Gf>.gLF()^Pf_0,]4#PI^f?9@/bMAbTUN@=58a]I
O-dF4[b&>Y<SX,\Q:4YX1R=7AG:;g<fW9&bHX3,9fccCD.c\5&_^A-2+AcU7+]VD
T9H1N-d2J2Z?.dJYH></2.Z?WO:,T+(eK;K6]0G9]DKZ\Me22)(HT/WYX:8;9^I1
R?aEd4g_O,-7JDeS.g=#S#52FO7U]1_>e1VK#7_-R>SdC]&)Gfdgd1baS\aH:S0I
L<N)SM(V#=4W?9(=.&HR<CNQZ-@cI@O[.2=UF-S,JZVR06@F:f368e8@K7PG,aZ,
1F)29[L,Z^Ia8M@Q<f.1\fX2b:f9CHNO.P0cf7&c?^=b3b]Z7>1^b>OYQD>ecQ@Z
^IGVP@HH7KBQ55)W<Q:2C(D(+:P;C_>J83CQ,efV,EZ.<\XP3aHdYL0_^f#OY_-e
edEg7Q4-d@4719d91#QPeL:_=W.2P[[gXcd5&+QKOLb.&@H9eKAW);>@T&L>8<.>
R^D&-:S9<\S&-A(+,^dd,+0/KA](T:1&eP:1=f=I5<A#JY_9LYXLWR;@2H./>^d-
)IfGgBRIHLH&>N)D7F&#;e)JX;FeS,47-E70W4\RZU63ME88THPM72[5=Z1+@P,[
C>b9^6A,N<+0;=^\^g_N6.Sfc.5fc>4EBL97R75JaeU-f,ISLW]\I7d&?&_/A]B>
IG0ZP)PLG#L7X//g#.@BMJ]8+]I\P;3O]e>>LK17Z[,J<0YYUgc(gb-4+B_gN?QT
<14-D>.KHSeA?/6JBVT-M<FD7@-#:cf4@22(KUU68O7KF;&&eQfD5VPc(R+:f/LU
6T4]\XO20g&Fa,S>cZNS24Y:9A]89.SE5+G81DQ/,T34:?XKO2OdIBM#.XCH3=3)
_NXB09Y9gF-RL>KP9P/f4WT&Y9K7DTHf:c^f<aV<d.7dH+;;[Zb=D1J_aV[NGb,Y
W65@5aF9I[K9MSW=<.2=<^UKC/NNLK]:RYR;ZU=&Z?5]M_N0;A\gF2fFR2LLRXWR
\3YXR\c6[31XH^>:Q/>VVWFQMOK#;g+c=H)SWW77AEde&dUFG;X]H_UdD+8gN]U3
@0G#\^@\:66WU:-SYF4#9gAFNQ2.C25M&56.GI[I#MU]V&3_aG2[-D.B/gOW:;H8
>KA/<?8/77a_D=gFa^2eC5+,bfd5R;E5=XbD[86E&dBf@W(4=?ZXT0O)ZCUG0Q<5
gAW;KUE(bM^g^0fLC^^.DEX;<NYZFgECbdYc&L<g;M>F.2-S]DM62@:FaQ8BZcFJ
bN[NK[=W_&0VUZ@TCOe)Re.7LCJ-LeK]MJSJE(#e2^76+YV8<+5CX>^gFR#Ic^Cd
3TNC_.USIG_Lg##/&7Xb4NQb;>1fSD9U0.d04?P,.PO7J1]fX0(R,3=.8NfV5\_J
HI.E2XIW/7PJ)a<1c6VA5#;O;W9G:C@cJ7B1,a]X7A<(8E,QMEC7_GKA6F4,7+G[
adaSH7M9J=KG9cK>KO2],/[XJG3EV^.<VV8N:L86)/CQfCS4J,A#/,,WQg3=:5B5
PCRQ\IMJ&e:?9\g=D8UP,2+L>WeZR?<87\d,7f?aT#B27e+Ce@1d^;Td+V8bI5VT
QBA+BS<GeV\>,PWg\H_/8=)cbQ7[KZ8;[PPIQ\)(NAZLW:S]R9/[FNcH98J_V=B_
RIB^(<A#UD#_7+J7E5ZJ>1R9DKDg.0HeCJCW?a^]_7X.D_57)X;]JNMJ#Y]D;0&A
d(e.[aRA0,;67[H:YG0MQ61.@Y,.;_E:A.RQ1_5HMUaXWLaI30[QKf/-25)QId-d
^g@KD.;TG891CX)Rf&C&>.P;KB_4Z1RBWAK+b77X&gfYU+Oa&TSNd(1-\dUW#:?6
\#f;S0@eWIbf-,1[>eQZY+3@RNNe5C.B--a:824a5_559QgYN,<<=1Z&,1M/P=\+
H-KW\8:5L3;R\eYLB6<@@W.dI;7Nb+9d^WQVY/H<?UWC=+J^0OJ:X/gBaFI)_7TK
=C]YU&fda&N=^D(@<_9JPI4?><N<BW+MPC&G,:DBRLVb<AZa\4Db^201]3Y1Ocb8
V,2<I+<-B1Rf1B,@>JTJIA=e_RK^Qb;O,VJ].K6-:cdX@\+,O+aG\OM))E-]NIK;
P+A2JX9J?/<PA64GQXV&60?17?,c@\^ORJ7^fMX48OVR\dYQ23f<bG4],S6]^YbD
:#5\b#.M[I;P2/P.PD.]F?_TOZSBK&#6PZ(7FBGZ5CLa7NeXE/B.:LTAU:3/_eeC
C9<4gZY4H25K.EPDdO/EAL9G,5dPR+4J>Tb-(F=B#10(@N.5XM3F;M8bK_JWf+9T
.F3SSe@&1]G8,KH[R5_8bF1+L7C,-B:NRRY:&^Jc+]NL4.^,17/Fd?0N/H<<fF2g
c;T=:IYQJ<?K=_-/fT2&Hf>GcG2C4=Zc\Y3Fg_LUQ)]GZcN>[&;UeH_4KccZMB,\
Wd&:[/6NL):[,.8\#19M(<:8WGQK[HZRJ@#HLIfKM:cZ3eBd\_7cTVLA.?d6-59G
=^GdYRW\?LX,AGdJYa4:JQW,850T8\9aG]5++X;:L0OD>cXY#D.M#?d6:dWH-[VK
M\:fa,<OFM@B+TGAOX3X+TdQT:aI<6UD;#5B/MXKc:G=T^#C45C<F]F0&CF0g9<C
,P+:ZJ:V(1;a)g&FQAGc,,#)65<6@7T.X01fWPY]6ADES_.>V_:4J(;-fE3&0,F_
cR(YUP=QBR&SRMLc4[cYCE2^3T6d#G8#LI4/0cONT:05/E&>/NFAX=U+#d1JP_XS
O6bVGS<^;M25#;G>Hg;ac9?_a?,+8<+I7C]Ue:[IVT3=R4Jg=+.NO=&2H6NJ0=:?
U>SfB5gY1aPNTNHFgO2C[Yg@.3SePM@](QB-^,F-23XS,3OgWPGCVM(LP]C]F?=@
60SH]BL=8+g)NL,/9[B.A&_<=+7dMFUR^S7L;4)b16]V^>^D(BBK(5W8^aA0<G?<
Z.I/8RS4OWd.B43/D9W>Q8X5ab@CJ[]D?6\=M,/[HCB,Jdc,L]49)].8ZAe-McL7
4>g#&,6@]0=6WKK9TX6fT6VZR6[,)be875^:FVU^/WMA;II(bCT/V_X6I0^I(/LY
>.fFDR9KCY]UGYRXa+ae;ST?ga\EUagADE]-=O-+?PU.TDP(0;9>TXZX\a=]V).[
-Uc2SEM=bPBV?].fAfC?]V&M1_K4ZK@XR_F#]QZ2>\Y4]J5FJ:4W95OTf=^,HUa>
TUg>BKK)./NK:.BeC__T::RL9Uf@TG/6PQ:0bPbC)@<.,AAQ1:=S0Fgd(T9S)bQ,
ZeLKSeXCS3X90\OMH^0cLKE8?/<1eW4W51/1&DTJUG6]c&U)^ATA^WeSHH6BN?B.
[0WH?D1KHeV751_CJL<@5JA[IW\eg/]#Z_M357CfQ1K@>XWCLPf-3V&UFc8<e;Lf
6eXMF=).:3R1U),P(J4QC^OWa&#Z=HS/a3>U+Hf4SOES,dSZ_&a#C\[CS8@BT<O_
eHYR2e7P.6UB9.^T(dE_IU:6Gb_SKNZ2=>@E^84-^2])T@PZfA@4d&E,TF^K8HC@
U?2B\-e7-^>dBaF2@a0_HVC&GTbeW)@.=>630;SG>RL>@[Hd4cD+[-S1LREZbHfP
#FfW_Rd;69AG^4_QgQMbWKSXe+^(ZD<WWV?:R]EG+WLaA?c2)J7Z?H-cc?=@ON3F
-#5N1I8a&THLf4#^4Ze]#P#+I)W4L=@]P7=-/>ORd+&UG:dQ.U4e3,V,?AXQS#U?
a23fKc#HgQ5JY).26)8ZaZ1XGA]W-.Ha2\APNV-17S?6OCA1@da5VBf5=(W7@c;C
aFB6Fd2()e2@6N/0LA4>-66\HTRK?>P)G@V5_TfgC,Ef.E9[V#FV;b>@],WfXI7&
)F\ZY4_ND(KW^0\M46R8KNIS(4CUQg2B>FNfE:.ec9SUF2\30^5Vc<7,>6G7B])1
Z#+SNE(59DK)@O1[g5gT_cUf<Y60HJe_dUg36/PWC7BbDG_L(1[GC)()f99Df+^<
DQM]GY\.D^&HP/Z3=/X8C^9EF+8W^5PURCAGdH0I;F]UM3X[8@MW_\fdND<F1V0B
g\O-OPICaXY\LLUQcBEOYH:_df,3Ve^H9N@8H/1[JK\-9bO\]cbFZ(3435J;K97Q
L:4,QcB=(8Bf1FXIH;d3=Mag\N,::P@0[eX1-J4+aedX&Aed.Z#FKN847893cX)Z
gdXL9EW+bf[XZ?@];LDfOIRUPcZScV(f[bZAYONZc\5^X:RbF0gO))[7YfHZ4D)I
_S6/f&..eKZ4FB[[S2a\=6Z4WDWK^-f.(G[<=g]0@&Z8N6TBM1(1WQPa4SBUfFO>
O;5U6O7HdY:CgFf6,]W.)4M#>,UHL?#4BOY>,gKZcF,@]0F.L:FSZX0+VU1-,e]b
_<KXWT;;50#,EIQ1+FFUa)bNF2H6&?PdX^egO8V-XA1.C^a0]TQD#M1/)7(L9/IB
=EX4DUEQF[U&M=UB1@&K08Bade\R/d?8\DZf&9c\+:\A/WO7_OGf:Gb55IJQW4gX
Vdb#Ic8c<S&Q:cN92D9M1F2f&>R/ZA0NeLYC4OV-Od@99:0Q2W94S5G0XB66:\#Y
8\.(=0/YSW+9,D\RY+C(Y\16d4Bf14;P_D-DGK2DA@2cY>2ZGPSE/Nf2?&144\,E
9d9+@=/7WXE;/+Q\#9YMVD&,KT>2:>fFTb7ZUU.M90^:f?I,;gG+=D)L1#K@1HLX
&>IJZPP#TQ^OTRT<=^be?Mf^JIeP0f?U\]73fQTY4\ET,f?7/C/M:N&&gd&N39A\
-eC/WAX)/9]S\RRZ7Xb,cE)U)?1-d;N8@f]IEggEa8;X1WWA&,+1L-.+^SCPDOE@
H;W1UP_cRg/6bZNFb8^Z4M7^@),SP=MD9,]#Z\e/TQF.1DM=;3P,J1DA9<LQcZIK
0GUT]XaHPO^1Td[K/)P..7bAP:E?=/5=-KJ@6TU?QK<J=fKA^5fVOR?I#gQAA\\L
,O5:DIKGZ]G\+K5C:YR]V/#TX:_F@)=2:P:FPc/2=<<2Ac#T4\^-)#81@]E7TQ2/
f/5UTf/H/CFAM[#NPIR&#(,U3bHC)Re=Ng7>@E1A8V_HZZT3Q.3POKFLfL)dfZD-
g_W)&\dI)WT(^2LJN[:,;(_K?56#f@(G2E3g8Vc0&5b\6/K)\AZO32D=K#,U3VJA
KWXJ+U,4^@#<32?2]RI39QS7]+Q4Y+#GU=7WK1Q[1a;#S(CS(<?L-@+K;64cEfJ,
NH/G,EC<4)C(aZN;^HFGB^W\SeGVa8[D0g#6+X8)>9?9&f;aC0TgX;T=-J9BH05_
N=f25XgbK&(gAL,-fSb+R95&.R3bJZ<90N9_:/MDNfV(:697<2>KIY=FCW:2RMA3
;.@._:G&[-)8e0C0-SP+gDb0;3<Yd;N:W1C+D[c/T.e@K\FXK1\N,H_KMZV-;M,D
Kd.YNDfeGcU:60]_3FI.gQZQd1BZQQM-W,XXe4D^[P&J\YH2)5?=TH(6G4KIT4GV
.SI]-_>IG4(-<@3R@VgXN&&EgHgC.bDfW^;50D\,/e^?U\C-ZA>;)+e9NN-Ec/B]
HXC1:g+T4W5URQd6)(bL&(C#(EHH4bZ:H<ZXbFYGF]+(AA.O-MB:=2K?L7_G)TP/
VIW6ZFJ6?0Sa0E4b#b\V5a3?@P,QWUKT;Sc3a4:7[V+;d,Q[2K)1<3\6S&=H2?>c
@E(=L41OR=I8T1S8-IZ)?LP<B:N[RTYG+Pa5bB^U>,N=M<(g3Y<DNNJ.KA].17,B
[,6_CfSdY7-,^A?<aRF&E7M_S9+0^1RJZ;fdJ?O7=6Yb9Y[PdFaD?CGIaH_E>YQa
@c(OcP=)Q)7I:eJ,Y0H@:<:SReL7;:\E<;O20)]?_3D<1g=c3NLYe1BKbf8>RZB8
#S7dVUe-P#&9/LK>;I>ULBU5X=6]d)Z)8KI:M._cf6(G5\;G+-]B5;Z>E1dIOEJY
KN]&VQB@H_:?7-PM_LeAQGT#B.7RQ;.DVI+FFJ<MH#,84LR@,G<F4b&Id-SPQ6K-
fQ]T^>/G]?1.ZWg8E@,cLI[\B?D,R-+(;CSQ[Od]D8B9./<V/XLc3C#9C3Jg7Ng?
NRg#SI,2FN]0^5?:^d42YdO@S+YWF]]4ASaOME6T[ZWAC[:\Rd5?0J5N,S##[1JY
L5a5]TY6XX^J-BJ7X&5TWbDdaKRf?IGG3A?bF?&YJ;gf3bF8FK@69CBa^OH0:d.3
<]Vb\E.<:\(IU9Q1[;,_R?cIc1W9K>+#QR3--+X7PP7DGFSXSPD3VdCO-G0GOE\a
TVaZbL/eR>NGd3Z:+/U?/M)0>Sd?9/-P:2-V]agUGB?Z2&-B^_V#Y2:_XB9>4_.c
d\V.<ZF<]/FALW\JV#;g6I.V0A>ZVVWI=(LD\)E>ZN<@?J:PNC?-(6IF76H9#bB+
]M(0CWOY2Hb<K?8(D)7/]>#VX/3O634Hf#DW9.UZQe[,?8-I.^029/JObZ>>]+@N
b2G&4fRPG_C&3aM1fNP&FQ2f.JbWed-6=FfcU0[9(WEc^;1@GFY)..9./+]/&fe0
N.0YR?^-1<L3g\).VAHaN>PR9aZ:E_gAI4U30W5MQY4P@8-5WV-1XcQ-_-gO]16S
c.=G:_Gc6P7HbFe>&cG7T@)V9P01J0#8UBQO,Zg_7+24X.fgO#W+3IfYb[d.FLJe
JD#5N@3;4]Z@eTGS.AH\T#WO_4L:\d-##834c-VT)/=dR;YZ=DfICRE-:R&O(/\]
BgeF+R::(D.<HIM#&[.V;1;_TP:9e2^D2M5SWOKA^;(SHOF:g,2+Zgb2DO3O?[g]
)O/P&K=5ZDH;IMB0=JZHH8S8\9_5Xe5T=gd@]aH8H@=CU5#YZ;e=;=<W8f]eN,_f
Y<(927/,g;QF@QM&PU9<G>[LOcc@+)?;/@4ZeM^-.DOB?D/=Ib>4EJ(FS]^,(B?1
)-Qg+eHS=2aKBZ=gXAUgfZ#.Y(==J1D:1fLX]6@6XE@7V:&3AH5I:<=RO_PKa,gE
eCaSeVS7T==94gD11UafE^7>.If)_\GC<H[bd]8cK)YJ@KV03d[@F,d2DRT@LNIe
B-OL7[c?d>-.:793\>#cW#I_=TYcc6)dc-FQM74_9^04Wc9D8aBW1C?1VVS7LTEX
ge;,B-:A>R&8\[?,cMQR6aTXJbd69Q(9\98AcOaKZ=1-]OL^f013-\+XDK6De7UN
=@7c[(9\H,FH\MT,CI[M<f7SVC^5WcZD2LAA#IG_6a60E^Rb(1aaK?<6VGZD(S9_
3O^=L4-Gd/QM/f)#.7W.g,R3LOT&MA^0/F=FCC7?;LQ586bZ;C(^Z.2EYHNWAfM=
d\X-G/AFb+/0#,Ae4^,>9I#<@C0TDS@[(PSQZP@:@@P(6K=5GU]RCeYdgI5[XID=
;--fc<&d/ER<,Se-d/.6-0aE?A_LZ-=@N/L4cZ3eU+X;L]),(N(_2C_cS@C=B>RI
?61_3O&>165gB8K?A>_K9MDF<\OI-Z&,6/\dWJ95>O^/&?HK7]L^RGOBf\C-3.YW
^@MSYCT8gb80T=06=gM5R48(:-_HT7FYEI=+(KO6@Z]/,&=_(]Z_cMXG>;4-Oe?T
1K867,)DX@2>Z0&<+WK3W9K.?[86V0M)XBNFNJ/fS,;(Pc<V;N8Q6MLO(S0E0BAP
RWD7]aF]/(H.4,B^;AGQF7dM]PCeb.7gEDG:I#bH=Y>0gedIZcVf8H6]4N^8UI9M
e47-NMcF+7a<N9\):c9S5Q]L3^5G:)=-2NRM1^H[@+a]6[H_E7fb5H3JU?,H++\\
)ZF6g#8(DOJ7;]>^L]\9J-)d.1A-,-cHAK5[XW<eH_(U/Z@Y6f[ERH=O.;[fIGf_
:GSUdcZ9YZ4?@16EB;&#F5&H6<0,9LHNLKb4dYBaE#2<LJ0YAdLAMLf@PO^IdUV8
D;GY&5,Nf1#B^O:0(fXc+L4P0fODJL4.eV&dIUdf,GWP&1-&c-bDg99XD5M2#L)6
Ab^=OJF4OKCP#^8A]EN2L@gb7N@H?]I(?]L6J+17/OVW[6)8<aNBKS\PA.:^R@9c
N/VUN[/LH<2NQY(D@cW,V_S\&[<2=NQFC@WY@F_RSV2+O,71dd&^P@DLF(&N20Xb
X@P._a+&V@YI)IJ#OSObHXN2H)T3TB-4OgE#31]&JdC87MD-,-2DV.,E(-/FV4aN
;X2P0b_KaD<cPf_;\2([Z]5W\T.;)7[\TR+T@(0#gGU+^D]e;KEH9[9\DKXeDR[0
3R4;S+^\(a&_Xb5<BcFa?+<?\BcV@]V:G]a_LG.23+&UFK5cF:+3UY.H]ZWM,733
<\896XNTKD\G#VIIZ7=PU#&.#,KIg+4C7GPG?.S1)OUP@YLfc=)?4]&,SfbYPOI9
O6\+?OVYZ@X96[A(@eLQS?K3E6aYaW56WD/dI=6,\@CSI5U:99e#9Y_-G7#AX:b=
[&2]/>a.J:VS1TLT8S=N)YA+4CbJ0)/0/C2eMIO2VP?(AQDeGS:41^+<>M:gf#25
ZQH;4\893W?IGS<^feK-FGV.7dGRY])HJKKf[>=VCBVJB/ZbISNf,gWH<Ub^EU9,
4ZM,)K:Tg<2;TJ2D854#2/Y_J6(E-;S6.IP\0)/8\feW=1D\D3RPM</I-Dd,>5fL
BUf)+4_L&\fYKS.1ZRW+-PL@@JcN7U8T_ZM&b.(Qe3VO=D76]T>=T>OaXJOVPKYb
1#;X6O_+0\A6e3KLW&A\WQ&[(@[@GUDge6LD2<UUGWOQgY]#BDEXV6B@VHW@fNDI
6c,,Y@Td_c]GCT7]VK=N)<+c28[)PF\VFOWQBK+c5L/e]/ZRZM8=K[;#1.a4T:^M
:L,)8><;.@?KGQ88GSNeP2[RHSFbIT3#NY#_._4/3#4P:L&YOSJ(:M712KXd=X]M
@[C38V6bgcIK2d]MZBQF<TDdJ?\@D#-\U/#HG<\GcI1784]Wd-.Gb?,3cb>b=9B7
63J;:@7@-f&Te_ZR)G,Nb,(M41dc)EURQ;KGdS;]#-;[KH;QQ&BOaZC2_[9g\Jb@
<#<aP_(,Ib>g6.@.a\4FR0(M2$
`endprotected

endfunction: pre_randomize
// -----------------------------------------------------------------------------
function void svt_axi_transaction::post_randomize ();
  int log_base_2_total_bytes;
`protected
V\-\?B[I&PFXMG.SP/3=MVV,QL\,G:PS>^1EF,8.LZ5D9<I\8IID5)b_2b&)a6XW
UC@N<0LTCZ2CL^O5(W7-9bD#,+e:IH([fa0TB50V0S_=(<A_;=/<Qb]?^HLT_ZU6
&].4N)ZN?c[)/:))WF_\-Y>EH;IR\2+].DT.>3_bQGS779I<\+=DAb/L+bYOMLOB
UKA[&_3;145Z<8CXDJ42N4SQ8XGA<,N0J?D\C1[&;WM?GdUA95(40,CD\<]SSN4[
G#3JW-[RXMRG#NS1@PV-W2P.W5GKY]@UKg+6Rdeg66Xd&SEB5c3.J1fGGRWH/J)A
-e7T\/-b7JF1#0G5HbBZT/O,>T[:[L]aRI+A/4X[[U<T.?X\Id&UA.eM=_HG;&3E
bA(gTgJP.P\_La(H\)FGL/Ia15cf\XD1&dWXQDXK9>1DYD&08[5&e_FHN_K@278;
\.MY,>cV+8#GER)Rd@_+/eQaKfZE:/NL]-P/0f[-7e<<>M=&2KB2;N(<H+X5E>6a
OXAZXV;bK>/]12bXcA=@EI0a,1+VA/[5#PU9SX[MP,O:NdB3:MMDfeU);c&M67;;
>)X;4e.I\D&RION>(70/3O)d)AN5EL5=:T5VQ9a^aF3PI(PFGbOJ#d9>1?VANRI)
N@Z[3D2BcAD.YG?9#)N;f^aEXIa7J]>R.JRH#_S3]8Xg.)&(eP_gS5Y2\]/4gVJ(
VBPaQJ38J[IJ(O.\78eK<3ZK/50XCBd@SR^0_TcHB7<>P66/;033BN1b>;M\)_K]
J>TFag<AbA>\E+@X2YVE8e26S(W]FVPDQ:GRb7d=PZRW1eS=OY[7,P&C6#:12SeS
,@&]1I>@fFI/c+0)H[KP;T_2&eFE&2C]bR+b.LLJ)^S(3G)=5D7:>WU;H1?1aQLa
XNH,2;U?Q,,1KE,e;.a.]BP4X0A<:]PG@[26-Y#+GE-H<BA8f<E+2IQJ10H0:]K&
b3_85KXB[cF@5JbV-;84&2>=B[Fb+P?43b8]&;WGOGZCLJ5#,N2^KGE:Dc9/2PbW
J#-:0(U(ID?dAC2&5^-EEQJ=3b&J=f\B^IU&Gd()f[-(:fF/_6HAeb,3;&\,AO2;
QW]2g]8cI.Q[K:_:3F&DV^a@S^Z[)6&8.E&Ne4Sa)D\.Eb4M1G2ZDEdcIP:^HHgL
c@JNe2BI>+4((6RcJJaOGY[9UT923bbfBG2:<G894@AaYWKf(a2<0T#1QOQ>]KQ>
TdFZ-A6:CPd7T2&@#fNdda5ffAU_==_EZ7>1:L24T1=EfF_.M90RAFc)\V5>0O9T
0g^?D?7W]C)5?B,2&+O8/bVLNIBe##T<HWSO6._d\ITNH?3g9]M/3g;?Gf\BKAbD
8VdILELHE)SC;g1?_W76Q<c[C76PYFR-5LJaBX;H=#Z<R[[aWd[ceO>26FX::VeF
]A;PFM,Uba5DKdFAUbM=(>::7;)6;-1?[:J:?1(6ZC@,D=M:Q)+bf:H\(]gTSR5D
@IE4Kf#Z<W-;Z(:LcI)CL-S/.2C:S=&Sf_R5aH&7/d><CIUFdMga?NH39(FIb.R@
[2?dKfXcO:3-:-bDA::Tb-9I)-FV[9Pge^1IcC&T0]3MWTB_]M8QMM@Q5dbA3)46
>4VL2)E@d^1,XW,6,CAGdF-DX[e#FUJaCGabPd?_JSccR\=GW-0_S2Z3X2K?Z,:e
3ZS(&;QabKB?b/,a>##S2)c5\PS++bHU6e5#+,gE;&S[dAK2eEbTE_d(\C)=)g90
\@S_GAJb:IZ@5IU&B8QC]Ee<bG.22CM8D<Ca=S\Z19RE9W5W,PA(\_&V0SFcY_\:
Cc3>N[e6\3QT&P/9,^FM^.XB7cUHMD)5>1+3GO-Xe>L?aU726a:<E8S+SUZX\WHV
CJVDTLeR4KXC+6I+?]B^PSQD6&2(?C-Q3EO1507]V(aNJT+d)d78#1O7A2@50OCP
.D/>2Of?d;d6b_:d3Y19W@J\BK1U10AH(KH);aH_Ob#3EH&^@W((S#e5>.3L5DN<
DL6?3P^6/d2&AR:^4@a<bCfZ5CT?WCWH5VBIC+Y(.-Z+COb\TD)(7K[Q<dcS.Lce
[:cIP4F><[^SYFbQ]G9ReMN24B=C_3B4QEMIPgO:^7):PO8I<18MSY8[,&5<5__a
K=g>f8PTf6<\P1=KS)cJ(<,NdE)0-PJ/AS;/eF:[R.dZ=+A9,J.(SVbWEI_I;H^T
U(aD)W.]Q4P_1GAU)d85RC:AZ.,J5>b_<YdP+1D.(:(M;9M;>3?d4.E&]_L01@bM
/2W&aLXf.1a5:e.d^dO6.^+_>VQFbcZFGX+N)?-Fc(9CbPTR/])JbCMGGQc<>7&9
1cGU_47+,ML)/55).cVTQJ;T@_&YRMD^[STMN[DU+><8JF+)JJH(;+fQe;=&WDTJ
XgaeKKa(2[@0#N_NKMKV>N1=F\SF0g+L9N89f6Cbc5cJ][7Hg[Q11;Sf0b()2Y(M
>b4EC<GC:Q4HSN,M[EJ9S-ET&a<B:^NF@#HUB;#[]VbH4Y@H7RE5RLLg8_7aV<f4
;?,I28)J]?&YFVI<aFVB::7<CP#U_70NU@UE[>CIKf=R[]TY&4]IWBGf:O;:=KK[
)AYgR(]:OQg052+D<8aWVH@DZ;=)35)D5+PIG7\2WL.NeeVDP;_1(]^WI/cRI>-4
3G6D&Fa>E/L1B@>-95_Vfe[Xd2fS6GH@-+c]JQ-(=ffaFXad_HWM2c6d?S^0bJ-D
G_,-+/\:1Ve7(LBX5G_V=UIc)g_#J@7U9a4[,P^c8N:<-(1RZI]HJ?09F,](_U&f
:U<T:8V\g+Y?UJKeMNWM&0N43NW^\,G0>ZTL3,T_2T[@_M,&#Oe-fZ3E[M[TQ6g5
AP-@=X8:R3I3[=5T:UcCP2G=4K_]aFbV8XSKCP#WAf&L):+=Y(9X+J8c.R4P7#9e
VQ]T8<7WbF/4&PA82c/Ea@HZZgGgOdQ1];?XQ#DDSNMYeZgXEBgFKM.RE?5)WUL(
1<cX[1\MLC3?]:d9)#+aSL?H;T;/D6;TQ66@UFAd;ZI+cR::=7X4?LO[>35#Qf].
a\V\XMb;];C6bb(I5Ua<SHe:3<]7][Dcg@\gg+V:0?IT4-?>?I]2:#,N978NOPL#
29G]9Q^TgYe0L^(R?+a,W(=5a1E7^QJ),IfPTf5S0<NA>M;9Lc;K3;GTLdMdO;HT
DJ.dB.IgDf+H]UDVC\YQMO58+fY#_+&dbLNJALLMe[2AJ,WS\W9de)fHF,:_Cd&(
c#0:e?[80a(O9MBQd8WVa_F,VJO[8+NW,.F\g&#/bcgKK=[bAeD>K.b@X&>C7@5a
81cU>fWKeC0+La#bR:\Sf^B3Jf2&L6VfOQ9\D?;^SVUc06Y_GS269O]9;VIg8&&L
1V-O,Y)G82Q^3/S8(-/(IcIC5WU)JW:)TJNJ4,G@Y#>f\72=T#@MG0#5QbZa.()V
PPfaMK9D1V3DT09,\_F@:Z,WS4,L;738=4VZ4(<43U#^XKZ.(89fPPUZS9Dc53Ka
/OZB_Z>NX?&.:\0=K-BU<^1Y<NCM91WZgPON9=F&6c0<1Z=b-#X/O)[/4HN8)^=Z
UVEY()6)+a[1HKC3=2.#CJTI5FYb_6(A<[L)d<AM?D#LTUUJ;0SK&]SU#X;^[GD9
egIJUY>4g4)0H0]0<H&WKFfR.?L;G9eXWe&?,^b7B)NFE\cKC[:B5^I)gB8-O_YP
QMVf7RGYH>;[E16&cJ/([Ic@KLfbOOHSDRV;VL07baa)JcIW8&@aX<_5]L>P^5[/
.F&L.Xe;/(5CEf@@bP:?A@YCSE\c7UMS4_FJA_+PUYXE98CAcAJC9SRBcD\bX[-E
).#53+)WWU478SE[DH/0DTCG05Sg[6A5:0<@-E50+D6.c/.]W)-452AKPL>Y7)^<
V6K/Y@a\@+YP?I0SecfCC/-6<4bTD1KGHO06ETE<?9;.@b17XQaFXDHg:TeK\]VP
B@^1XGEEfLX@=1T<,aDV@92AJFgaD+.@RbTd#OYJ&.HBf-EU((PZ/H)HA,E_3bK&
H:VeKO)^.cI,.;E.0--BE.@_H<WRZ=83SH2=YD#=V0^[B\d#XRRW(I)aeDLR:HBI
>2.G^\W]8J\4V/Q?/58FbWZ2e]4\bKE0\49,2b9.GLAFKW8Q;fCRJ^gBd7JU<O0&
R/6a?2)c19Q6A9gA0CX@J<>+S,EKgMO>E=2=B5R59WUQFQ+bZ1DeYEe?-F;d^R,E
O1SCX/H+abF)1]bc8,NRd7Y2>0D6-:2Z455OE7@+.Z:aWgg#;NXcODf:..Y2,PLD
5;M#R^+<4O(9]9Y/S[P&_3eVG>0G\_Q:-@_eF(^X.4J--fDMY<^<A<f#,c6f)0NB
0e#5B_4eX1FM(ecGT80X#W6L09Z?<d4Eb;U&>d9)>;S5CS8R6cDNMZDTEXBJ8_<\
X)3W?62c[7L:SSHSf@O+6ObO\[@aSAJ6>=BL9FK2Te5b+OYeE#=>7;YNM@<2SCaW
OTEB9J781^[CAUHdD7(;C4fV)e7-^EAQXWED,1.([:YQ9)6>5L:J^eXd--e14Z>@
8>)?eI:9_IY1\)0D[Rd-Z,[&LA6[daZKVD@TJ0<Lb-&(d7),,^?,&^6;LI[,DG7F
>3XQH;8@4+6^H<U?06.aEI+8VD_,#=G@H9Q/9&951@T15,GKO22/=5PaU\89BC=]
DgR>U1(]d4FG-N/?VefM-H0J3f2eS/S[f09_5_^1_(C]=ZTXeDPPS(09QIOM/XGU
TcS0G<8^^YN<,65cS7.S?5eOX#a9-#[@H6e\f5]+>c##gg#GE9X8;8-=E=@e.PH?
eR&bUb6-:#A@58X9N1<[I3ZG@YL64<RcT5BT0W@La/K/DfgBaL.Wg#@@V0Fg@(bb
dO966<NFRc6b7A#@B;aZN^JW=ee;E;feY>O0?;UX+T=:DX,6g:b-:<geJKYP,[EH
IJ+c;gG6+PUFDd8^<FOF4KUCKXD.bII8?U(6+9WRB3RO;dM-^#a.fVPX)LK.H(c\
P29;_J<bJH8R1e/L25&[>>XB@BaW;[5:<Xgb0/FE7@C)^bC@0;3>H@C^(XZS9,dE
P/P_4YRbMI05<+>@,e#(,]J:DgXf&bY5aDc10+b_5^^gd8E0J##OE1IYQ34)I6E5
7&cJ=6BgAV=Q8,;VJVE28TJ7)[5)\DF-JI[0Cc9fQZFaVG)/KOgb)3&A:EBXd.0>
@S7^SU<EBBKS3?C]#TPD]Y7[;#e23HS^3f&@MVFf--R4&,O^H&[1&,_>dbA;&?fP
F84DU5,e/[aSG8)HWd]<K5@>P<\L>H:2#3cf2,?b_4T2.#FCb767JJS]R5/^0C+R
5:VP<^Q#\F=fgd3GHSd8@;P2P+OH,9>Ag)\XW+KZ6\9]#Ed78B_M<0\EP/W;PIN,
>JPO9TNN2eE1gQBY.6VH\RVcHa,O7R9[R<e^d2[VD8T:29?TXL9,:aD,1S9X1N_3
LA0fQCMH.cZU-C5U0&D9^_KW_#Pa?/SbAd7d7//,Zf01K;AWT4aYe-a;9_F;68<4
XOdOEV0/.WDQb;8;J/c2\XRb]40XbZ5PI)bA<FBZT9+<#ED-JdZb(#cUdBa(.5;Q
)S97;:[^e:VWKXe2W7U-:W-XQU.=ab2#;+6C76&f)Z)=R>R9(If:bV9,E&7:H5+#
81[36U<a=X4(,+CRJ]L+:afDcbTZ=_RS6?FI.W+XffF<-.</<K:VbXCX>,H5]J2R
/G8gWT&eRR#8]9)P-d1+3=#@:>e7+Ke>-HW:cEgS>Ce10QNZ)gSNVA@-2[F7;IFI
P^IK)[3>4;cS?E0Qaf9daa4TfS(FI5.ZS54N?O=gbJ7faa+/=Zc/OPREX&G2e[a\
Sf=Z>6L)PN6+-LDfZTfQFIBGO_bBAH^V3F\MfG@9<?ENegfNYF72DC6_J+;(<gaA
gf30K].b/Me-IFZYD<gS0+dT+5dSQD)U8cB+GZRIE_cLND(N?]?g3Ha2UJJc0+<a
I]U48DR^7A[39g+7\4H\N:0RNY,J,)O6F>[WG-1?UC1R8;6?6g=]PQW\&:LR?+0M
N1@,49[W,4<f?\;_6ME+WAZbbB[]QgH>ANB<][8d;RAQ]=;DJg..PPbN?5>5VQX,
M^f)3bdL^aaX^-D.UBg@CH>V00eFZ8#Y56Y3677J&I?9HSV:S.B/QNY5@H9RdNK3
[7B)CHKfOgVWLf4M&5d5b@I_SJYD\bM.:@Z[O.:1HV>aRUR_FWG;>Y3T8NCd2V7N
cO,3Yf.];^N(N/ddE7^MEd<K6>.U3#M>BL:DDOK(8/O7fdC&M0ceDEXV(>6;5=1I
^cd@<8P^I:E#D86,H3TH<5K[-Nc,5:^.E]MVeAZ__H;5Pgf#6TLGZBSI6eUPR:&,
][+9Jc,1\=Z^N-G7OY_7;O,R\ef_]S.);>U19_EOd&2N4)I9+A:MfMG=:f.S\G/7
G94d)F&4UC:4I8]g>RS_W=PP<0XV^S[>ZWR,NIgEPP(N;_K3A7NYg4+P11P@@EgB
B_H\Q[6A-)S(Q7A)L1.0N(S(c@6YA,H^b]4LQZ,B9\@RP.YIJXeYMcVaF[1A>@]R
[41B#U7C(]W5a(I1&-cX.\U;#-VEg\\Z?JaH[VD>C=(I83O9J+QF;YL\,YSFH7@G
@BX>M>,FC&6R.#?V,()65#Y2-W168(X?[4/36W_c,T)1d,PK@FfY3Z+3U;S,fZ7(
6FSGIT]Y4^XBO5TgbIQ&_#-)DIR9-LO-+fS<E3+-M<U(ZcSDC#K7)G=]P(.BOC>V
2_A\Ffa=-XJ57HLA@YVI>17N_La/:cH-cK>QHEYYS]<Ab##cCO2AT>_RLUY:)&Y0
)YTIG&]VX0cU<3JFP.Q#LS(cQ;V-DE0,)5H9_BWZ/+fYe?E464/400OUHG79FK[3
c[AI(1P=H:&_&;2CK@:UXJC3QP(N2JF>UKgcZeKCE&5T]<J#558e[W8->#302FXU
GG4J&g;LJEb^6;J5V(VK<RF\TCa//c7MYe?UA/RPQHgb.3cb=@Y1g_.6S5/bFR6Z
,8WYf#c&RR3OgWNOG#Z_FaZ,f]db-<BPZd:d@06K</FaTc_;I>:Zec+1IT;\V^X0
;7/>+8?JfBDSQQ/&aYR1[;g)2YL;HP15P1]U:;D@IbX-7L/LG,X^b1b\PAOB6d?5
>JAFOaag_ZL,RX=4P<6(.DSUV)gM;ceg[,+C1=6>;2=bR&1WG+)/U>.@b5X60Dc@
+)SD/]5A62-X(1f1N=?BZba8c/FH1a;/J/9(_FJ6ZbgfZQN,_1)J:(5N)0VKD^B0
eD_\S=97+J2J3XaDMPJRUEfLKgGg8e?FHcTZ5&76]a>/ZM9dR1P8:J?>?:6B6G\R
??H5BD4-ZNZ_#J/K40eIE^/<f6=B5<VMJ8d<c<>A)#R9:<]e[&4\Kb:[5.<+F\SZ
R,Z\f#@VHSD.cX(g>EG.RE\MAZQ+B9d1L4?4YT1Yc(5c/@Y-UG(\X=HC?Na5QWg9
.ER],:=BA.g)S[a?U6,O5M<eY@e1;.\5TeWMcfU<-e90c;B/IUSO^VN8EVIH>=\\
c)=Cb:0.<+OFd=HX<TEf:YfPF0(_8g0g(Z_3[J-2dd^<4H4]=7885Id7A[39HS@K
>(BGNcfWAMJ38X;eLWE(0<Ke28HK4d@U_8WdU7N;(MRX^^Q__^G#H9dQO&+[cEd>
,e28)>/W#K]BJHY5KSd1L/JW7]2VW2e-+92aJPKSF17&Y5;]=>_5_CG6<_X4(Q?Y
F99=La:<;&f[K5OTeCPXWJceX1U<I)X4]GFSGC]gc-^TaKRZMZH8F7YL0I8Mbg>f
#>b1:>2([U8TfGaSW4PSa5&GJdS^Cc/1VH3d/.#F2?dB^WI5/=M4RJfXgbA#-LT#
RNe,^5,AETc]dC0\RN1MFYL\6>/6=\D[b(9_&,[JQ4].[[D\7G^SC[bJcCA/A[aQ
B-SR_.23e9D++B>MA36/^?(7XY,dLA=+<6g0_2533ZFV7[UTDW;V&MXbN&QfK\#^
]<#)@;VL^49:D>+;BgVL=0YJRGNY&Ieg4DN(FCQ&aCCX;g6TX:N#K[e?\^IK#/E=
(-gTb_WVU#Q\CT[Y3c++JB:T&e&^KR/\<Y^@-O#)bJG\X]A&DYK@B?]V4@FW(MFT
D(a84I(QEc@KS,_;RM/(S8,:=d])NI-WZWWO#f.^:K6:(]Ne)[^ENR-NcAR#Q3gF
EM/dQ_)Sf:<^F>4X&aQPVc0XIUF)2PUP5_>E.(8>BLO+(eF3R3.AU1][Zd)=J,W^
&GUdb/K-#E>_1KY22FF8CP8WGWg_;7,:IH4)M]N(_^[/WU/fg]cYg0gWS@I=Y7(H
S&GW@C<cTD-FX8-?a+.4-#REC3X:+KED@)dEOUf3?bXe;@)&d>QPUPZe,T_65B1.
HD:.Z=(FZ-5B#,5Z[.FG3D3#<402&D^477+e2XO-0.\H>d9EDDHFg1&=Y_4a[9,a
a,@&4PVYXO5a;T4-3(A5UY[5/c)9aG:f9&/MFUL#PaW:;.P5QZ=\;CI#4@N;d;JB
HTDfJ(YT)g7:QISM0E1G+dL6)C@.5VG.1FBS3#9aS)eW4E@PO^>U:+EJ?fdL&GWY
U@Z+S5PQ#Xcbe<C^S&MC_7T<X:I-g,=O\]0g<Q32V7.#4#MVJTJLe@92.X(<eM#:
&bO@<X\K9fJ:)FfUaAd(5RJS)W&@4,(8;ULV:aVHOC-7/1_^X>21cKNH+>8^Va&W
HHOPL(N#YKD+G^IdJBbF8]?&8?V70=VS6b1\PB._Z0IY_eNS]]UJ.J#08Hdb3_BQ
=<;Z:,G?71.Te7T80@F.ZYNYW23R8+da,7;YDgHF7SQaT7e8K&X[&R5TV\.Qf/;;
RO9S=#(_V7OL:LDe[6eE2U:FF?ZWg.cIO9+40X#d3&4@N0;N(WO.4c_MCHO&,QOR
>V?,Z+I9D9eAMeQ#9RPJ]4\GLXP?6,^\PX3P@SH?#]]\1A6TSQP^:AgJ?g,d(<.1
#)&FY]4&AbPg0=S:cB0#B:P]dMf8]\L>-ZH//HUPE,+7.gZ?)/R3).J#f]LfO2CH
2__SPGSCG.dU&)NMRYF<gIU7<2a2#1[YKe,+8SZad6>,A](UKcCaL<H>;US3W^/0
0+1dBEVQZ1Y.02&SC4Ad=,VZO9YH)4],7X8/5SgRZb]MKE:I,:P3<;=Y3JfbE:X1
L(4GJ@8(@?IJ[4Q;T:U<(^-\=&CG^YK6)fZ#(J29H\T>V+;=,&;_KUSfE34@RCEC
#[.N_(;LTe/:LJd,P8HBaEJg)LBY)?.\W6Q6V:J-80.6;SR>?I/a<<-_=RZ/-RKS
FD8/Dg)LD@/SaXAA\aSUG/MKSANPKYE-2P+8<=TTUR@gRBI\cd(<=6BV^5X@TZQQ
,Y0Gf(,C,IdV))OTgKOZ)PVL+f(\(F&E]bgE/HNF8PF4^KXRZTSL8QdTJVGc(M>H
aJ8C_Y?3Ed^9Ef_,BRdLK+gZcK?K^KQW+&bYUd40^aIQ5=6,DIR5;Q@I8,58WHgg
X0-W:f,SD/S/CS#JN94PeS##FR2f9@fY>[M4I^UKY^2,FSd.?NgRQ[Y:#[B>Q4M@
Z)dT9)<e\<0/5(4aMa]=aY-XUcOS:Ie+\^133B#6CPB),AV#0LF0BB/W2EQ9OZ\W
^6E-KW3BS3>:48LX1.)RQd3GF+Q;64^D-CgSF>,(#NP^U[K-3;\,>bG>&X[6a<Ra
7JRW+.c.ENYV&.K;R1?8Qf3G7$
`endprotected

endfunction: post_randomize
  
  //vcs_vip_protect
  `protected
QL_0>b_,/B,<\FFLYL93fdJ5K7&Pg(9KS^3M.#B=MN[)\eA)c?ZQ6(J.F4.>/>&_
XGEO[U[&aVg0-@UC=-QHQYU=eF\AOEZ3>9C-HYL>1XQ:(8UMM(UYC.8e&fJ>b<gb
Ab(LA^cK+\PaK:dH8-L5KBdI2@=O^HJ0C3(d=N1f]d<NKf;PVc<,8RZ5LVc_0_24
T[.\F3+e,BK(6@X9]>-bT:94=YWX4S])HbG&<6:44<+SU5[g;?10g;B\O6TS,;cB
8;KR,5Z]9e.HFGNc&&=YH@eNRbG)#Nf0A8f9R&A(F#MGcYR#[SLN1;V/<Hb5G?=,
_^b9#MK^D45KC4[G67f>=11Y,1MST2AX<@2]9RHBK6b]JM85>13#KJ&H1fL9FJR<
.?g&961,69G+<=H+K?8/V>/cJVNX@\cW?2_-B6/X;Z/c@8<P:D025X1SP[Xe0,1M
7A1\/+UYVQX27a887,Kd<NbN-fg(/VISK+OU@WY699/CK^cVDgR,A7O.a1_eA=1B
I5dF5T9L]KQ4O^aK#bM++3;;d?gR/L+baQU7,VM[a177OYF-We426D2=BO4W^NT5
^J-Kd7TKF8f>YM/T01>.E#]9Bg-Z:N]NR:24)N^cKb_@=_=#=-OF0N&c/L:SY46C
/e_V<VIU.M\;T/)9gJ<TE]7HIJKN9TI2EdL>-H&[9g-US>?4cJ[NPER-X=UDXX+f
MZPHW1)JCYG@@>a6IY[_J/PEAb<9g=aF&[c:LOY\a(]UE$
`endprotected

  // -----------------------------------------------------------------------------
  `protected
3aYaV_>ee5Y>D<eW:QLB?:UDGG(H//Q&(4\1OJ22SA(c,^BTE[>U))bVBIK:gb\f
@CWb.<=ST?(9&Oc)fg=:?BUD1$
`endprotected

  //vcs_vip_protect
  `protected
>TQ^+:J[U;\BJ)/L:3H8:M[0Q87V6)(P9WI3&)DgBf+ga]KQ:Q/-1(I>gHS]dX8P
8)_.@X6:)Cg,U\X1V8HGcd0V?:GM5(NYAUP<0WVCRPP;T-A7[\3G6AS_,Yba^,,Z
XWOJA6&KR7KW[.0Jf,CXX9WCdPY/K.,U^VHZb2&Z4:FE_1?e372=<;7a+Y10Y_KZ
+G=5=)\\B1ZFc54&S)U;M1RAM7A;bC1O1V@GT^LGW8&99J#BL2daV=Z_3AXC^E2L
F:I)cXZcH=ZR.B.(8Z3cOCA=A>We5A&.1>QM0a.2f^E/Vf8NR,Ka[SK;2?a^)OfH
NcW;?K<9/58(/=b#6SeB[#U[JC#3Se&cSL)S)J_>^Fc+UH^.&]/3K50HP=Z_C09G
I)\]>&XBa07HM2a;T^_.O-,<7Wa>V=-fg8@2SNLZW:TR=aA]:IG7_O:e(0TZL\J;
fSUE6Z+;/N+<X)DF\;F-;^4RRX0cXQCY4e#2255<?O2\JV&RAIU<OX)).fQ48AF+
759,W()AT(BJ#JX#]E,eeeg\gRJZ-Y2]5##J5B:0M4eBZ?gEaaP=H>_?Q;8bbVdX
2-e3d-A:bVC.:3QKW@\S\cZWgF1A?9S4EV>RWDG.5\;Wf75)^Z5.HFJCcT#PeeA)
bD()K<.,EdY</9^^MbFMC;WG0C90AZ5<-6a\HE2KO;/.5FdR)@?/5H:C@d0].aG)
LH+04cSF@:M([RK?_Q1SPX35;(Y?@TgB:_J;89LFU>]IWAa7A3TQR1O5cHIQ,4Ra
9.A>FBIK94YAa5)7UMKMaIU+Af@9;<8cc6V@T8#74=8&9fJ[4+f3Vc?P)<+#FQVQ
5g#)K6+8Q[+@(W7JC4gLN:,gRI8HBW>G_5^HPJTG>H877964D@Q)^(DX^,8_0TbY
^;]WWg0;e\]I6^/5EE3JOE<O1:]2VDZ4F+V@Y-5L;1KP?\dQ5>]^>:)31d0786D.
^+NT13YY)+):48\Q\Z3//SeIA(;N[][P11QA_QFC9b_D.LX-8?K,_TMM]/N2LG(&
edQf_/&[6JX&bBUE9bGNMgc:+EIb=M:H^d#-0DXYMN2F?HB#GcVcL.S4Y?[bf+AB
NZY@b6];3[P8WSV)8IM(gP-bef-SD1Qf\_UUR>3\/W6VRg0e,V\1f2H:bUR\^N@;
?c(YV8PS_F@4:_.-I=ZH7eWTeFE;bB/NI6Z\7bE9d>+(MaJ]N+5;[g=N.5OL1RM2
c77;/V<U2UT[cPf[Mc@e;Q/ee6<>XU;EC1E5]?B,SH,>:K+XV>dcL33;H_6JMBZ)
-DKRD25Sb[J6EZbZ?dAf<]1)HBYK6[.W8V/:.GPF+J/1?1U:fB9X<#32;378R(QM
LQNaO,ZLX2_))c\0AZ.G&;S3,AIe001@4X6D5OFeZF[eMdOYJ@[(K=I9W9Z/;1DE
39Y955/9fEWR)>d99FIX,Ae<KA;@E]b=\4K[Y7,\]??,B+9YRZQ4fZD1?f2BLcGW
YH<-e:JO@0\O3#e,-S7Ad^U]fPV_2>#[Y[5BBJ1>)O&b9MDV=;CF)-YFgcM(+V[U
FYK:LQY(B<FA0E:+Mb^T:MWM[8B,Q8.(bY5-7@VQ[E@BeTU5b#=ZE]a3-\ZcGNe]
;4^DGS6,R):[JX8TR<V#VR74-K_L4_6G=\.BXDRCKT6-cNY&;G&UPB0,M&,GA6<Y
BB44F,YY3<_VIS1#XccLT/eBNP(.gF+;ME(a4:f.ANE&C,&[L-MX+NEJR5@)1.+C
G01bBfZ<BgY[1\8Y2RU7_E5V^?+d2.5T1N.@1I?X]2PI>G_D&-Id,FJFL1(YcDaQ
d)+&DSU)8^_0QH^2SX,57a=U-\H[SdK=C7a8<\Q7YO&G8:3g;4NEWe12,3KcU4fV
86T(MB+IV&6?_fV_</gSX_M&J;ec=Kc3Y,L-RG5/:SQFN],;1H4S]#Q9+Z]E^596
fQ&5WTYA.K3+JCD&2@<ZMCeNM/3ULHU_7-VdcS[6)#?O_6>NA#0I0I7Y]b/<79\,
B2_4,N+g8_]&@g<OI9SHVD6QD=B[X,3dLP+@fRaF5H@d5@]UD>g9X5G4IS&ZR<U]
.HS3bL#B-J2TCLDebL-c0Q+?O^gF,1QVJ#X>Sa-3eL3F8XC25&HECTH:TCE8KLS0
7IVGBM9;Z5Z-500/9(,8<a.60)/&&HKH^(g_0SHedE.+N=AecD])E@[/YddET+A\
\(]-(FTD5(IUeLQWNC_DD.U]\9L?K?C(0OA,^D3:;KM6&I2eCP0Z:=U5;)f-II59
+4a>6HAVcV_ZZ4HIIO6O6RT3==92EQM>)92?Q-0VH)e_>I,B3XGgJC8&R0MJ\ZHI
MW5bRLAJRaH@Z0H<L)Ma_g70b6b^#,@OQDI9#1#_P8bUcV<KC4+>GRY\4S:&/?dL
MT@W>^M;:+a5/6>QFe=RVG\e@F0T<M0?J@XM,eYVcRN_Z9+][2A0\RW?([^^Bb>-
3[\T&A2CN?Q0D:N5O2W>D9gJC710aENBDgMVg^<@3gOKb2Yg\3c?DJXUc;K/+VH4
-+(]?SQJV/_JQ3;Fb#])K]^gAL>=/,e38K2^Z4=HOF?2AQ-/bcH6F-4>3bGF_g1C
T3gR^.XV@EYKR&WZ8P3HBO[E^TNRegQYUE2POE19:L6Gg4LTe?We^]g&RK#9(P3K
\?ACV^beT;,g6147A_dMG7?[;12aA;#D&F&+1[a\?VULc/fGCTN::gH#?36f(a/9
aNa]1bI6(,^dF3SDP_3WA@faRFYK?W2P\Ic@8fD4.GXP4,e<[4@B;V@_\W4(5Zc6
Q4UD5@CW,6M4Df0GG-DTAZED)-32F7H=aY8(b#^>J>\C_ECE?1A,e6&[@4c;OHeO
+G\?Z^,M[,[EJQ6L_D_R<V[9cGF5B7cbPAf7QAcdc]U46aF]e?-)_#^[J9M-_&Zg
3GX;cU28K@T7aF/8a?SSJ[cZaH9248X>ZN84M]bJ;GBFc<Ed]3]YAM.D=LTSJcUP
A3<4-IO<fWV]e3d6OHO\PN\.:/U3NOY+QUV2^VI3Cec+9W6,?MFcQ[-5<,C(a?:7
U9SH:^E+bSFKPN(f5dc=]9?DN,E(N8B\5(HSc0ESN((L,CM7XBb6IZ]QFPPRN.g?
&7PgU0LX>4_ZdI6>TLV\VDL_Qd-@])]BT3_48G]Z3LbGfgO:H3.HV(RgRQFJ,>[-
5NJ^YTAE#YK[:\=8>RFJ/I?6J?KDXeQf80ZFRK&GGG[3^R#QW.OV7@GTaYT3<5,R
#3V.?,eL;-c]g2E_UY;XE0JF[)L3R6/H;F(2HY[VY#_[3HId(=BLbF)9RK4Y\>(B
^XL#ZCSLgTS>Q(Ogb]=A__.K-ZSWHDMTf1::#C+)H.85bbQ^L_Ed;W2T(^YCV@)9
S@&Y5f50gR(Z(+CU&aYMVX7Kf;/6d4\Lb6W=Zf&MS5RG;f>R4-.3\C/X[E,NTGWA
VO3G?d,/g\E0^/@SdR8aSgM]S,]^>1:L+),/_5[<@/GSH#NM(T#-FFG>fT_fUF]^
JISe)O/;G#bAO(^__O3&TNaS,-6X+.RYGM_00?12JbBZ<a9KUJ&&C:KT:.SSDQ[6
0a::?+F0X:Yf+Y55e<WHI1IN+B0R1M1@[;RPGE12>bd9+4(Y06J55_<Nc^=-VSc:
H8&1+-E<G3F:&+HO@-/F&@9G\:6:bW<PI86,-,dN#U>K/-85[J-6#df,:4/gNA7c
d4F?.JI7\>PE,U1Lg;2ZJE.+GD6f[7XNKU\20F(d3Ng._D@8,Y65QG44e0&:/Z)J
](?,bR1<L3VR5<>.B.EYf_UHY)-(HM=@I>C90<_Q]:D6gU=0<OEUff[NUeXAed[?
SMO^+\J6_L=ZJ1HJU3OBMA([N,5CXZ8X@C+J2/EOA4KPa_OR[f_W7<a=1?19aH(P
=:U:TLad.].1g5QRf.\:/]=EW_LGPUU\#A\W1^7&BR4V>U\=)..5B98d,R>9a8QF
=.,07]S.6)d6Gc,J=I-H,aEE(]-UU\)0;BO)&(8fd92PEbcKK4c&Z6)3LFPG=[&0
CV#:80VZ;LeEd(J(/=e9RPDPdBaZ(IBIUf[<d=dN<T:GT<71Y;0AX6VU>^gJ[?&b
/K+@C_Z]ZL7D.W9BR4aU5K+Z6B20)KT/gZ\bQ3KY-/7^AZPb_?P[KBXCe-C<[6IL
bf]\V]&T3dUR_aXFdb<IW,;g-_?b<HBC.BR51&QeKgC;F6,(Tad>Y9Q?;ZF<-CZ+
N08AZ&BcfK=gK+#XQNC3R-TQbI]agUT-)K[7=^<:g&[,ga:_F_R.0NR8afDcB:-Z
0UWJEV(aE0V9g7=8UFcG=1EVJ<a<LC\I]FEd,O:8O;Z=2339#+AH>\FOC+E+g1_c
<5b,-9M8&6LU3[[cLM5B)_V-E35V^;68CKD?#6(X[_MSe<@)I,&WUZPZBB3_e#HM
DO.@3<Q+&2KNXI^bcScO]aCQ@8JT_5&B6[4N@89R.58^#FJOZ9\>^XRg0XF3M[b9
f5JHb:\NB<@<?GIB/AH?Z5f17ZS^(:G@ZPd6UY/ggQLBA,]d/Q+XSL++\IT-UO9b
56=@3\@?,7UOJ1QTK1CG&Q(>E0@>M30N@7#W(:dW<PZ.=AWZX=O/FN2].I@4Z?&K
I0PKXT5-4XG2+#5IAF@bFYa(U:CNXV7X82;DVP2HE<gf=7SdA3SKd1L_10:_gcY7
Tf9W\JQ>C?GU;_;)@X.dP8&[f<TBb[3(SMK#4-[BHceAQbHH-Wb&C3[D^ePT6F(S
0Y=Ge)J^.1VF^aVOMMB&\5VBKd;f[5,ZC/:4#A?&\fR<A@<PJA\]?)67a</8@861
;8U1NJ90#L_?1JPW7e[)&JJ:Pd++d.NU;0YGQI&N<RVKOc7NU37DT9Z#@>CIbePM
]U,\9-]&VO,?MIFA[/7[^D]OXG-#W\cV]M/e3.cU]&?1U.(JG\OWT)6306Cf4\@J
fG/dJYN#,A-#_@/fT10.W\L&&#ObUfUNI4NHde#NT8dL.cG.gdR3NfX\>6:6404@
1<?.B8_Bf8^LE3PCTKRJE42,);-KO:U-XW7.K&FYESSUC=6D76J6G4/MI,CRM&F2
MRd)REE:ba6X\\S<S<5N(\&DeKXP\PD_0,D^30:<I=+>]A9[<LWCdR\W?C5PgRd]
Q#:Ag^;/06BCXe#98e+\2C4MLa(N)V.T&?6b2Naca&\[S>YR.75(=5[fO)M[.7)5
VK)_S])-S<VKCE#3-a6e/@4-+Nf1NV4])UORX7TG@JR6)^N]S[c(bF>MT3a/<;<8
^?3RKJ9,L>M;\QOQb/;b-gETe1efWF&U)\Z#NJ)98MD-V#Z1d6bS9^.dDe..5[=d
^V;OUPGU,Cc?4,E&PG998)GE_gd]ME:^0gg\=NOa\G_EK&E.0ZC1XbfUQ4gY&<O&
P_Z/<[Q]M9&B^7,dPYc(,VLW-eVVR(I.+I/EJ6c+@)@.EAJG_=[4^=bC1ef.IN>_
@8;eAb;U7d273^#Y0d=b79V3=&=g_a[MGD/Da<85_30g7ASPX(3.[DOOaS.PF##+
.CD^YX-(HHC)XKKG^51HD<&C7US3JeQf=D9;E<@_\VZ(S8-PD7+\C-5:6b]5;/\R
YRb)=;(I:QSH_JS?F)X@(++IdKR;(23DV,MeH5U,eI^:8&5L\J@4M46Q9]CHS(SK
[6d7#FAI]ACY^R)WI]QXEf3dD=QO.Cb_^^DS4@5=bDAa:9cNX7;)WG7c?\;GRc?,
=>DA4AbA>Ye)(JZ9++D1cSE?LIOP)SB.6VDd3=<?&5.Z@==:?2cPPWYHGKPRPAM#
A5W(8gO/S-[&@HZd@@8OUfKT@g+&3T:.?C<+W(^(De;YGYG&+R:YS/RT8QGEI9)/
0Vg-F.-b?(2L7/(#2Y;W;B)YZ7_6WV@PJ&3S-Xf6EL[&Eg-9cffY_#4M8KUVD/J5
8EA(Z@2?f(9S+/-IIb(X[c5Q3PZ(Y)NDI@#M;\[49g>Mf201K,&>5,8>D=eIAa@3
\Z^bU4?:?ZdNE8W./T1EMedNWQLGD(N\&?@D8Y2<#Y?OZ8f/>8LU0TP_S/PUJ9J)
&E;f496YfW?g)97;+75\fIMAN@6)&)3D[VbF32cS-RR]/]5dKFUS=5PX\\=HT=W#
2.FeSVST6RUId6)-#T##P8R7.ePLbe<#0I2/6cFZHA6<DD-f&Fb]cT9FPQ8PM7aI
^V[]&f@N(K1#UbA4<._2bfV]GJaMK=MaQ++-7I><@#V^g-XFc-gV\:==M=9AJTVd
;\+(?e?c1F4VcS)I3;3d9MW,B#>E)?DQK92+F1bE+MU4HNdFLQR.4?R9+[[=e&FV
EVQfF[3:1_<3OT[M^)?c22@)f->[VcI^c-W5,4+^#KO=^O5UIAAYTDU8dafT_HNE
,-I(0_c>g>M(cg26HTKFLJGfD86cF?C#:AV]:MN\N(-\6Z]Y0cOUH;Q(HM-;c2O3
+O5XKa_D8(WVB@I6BP:T/gHfW+MU-_dTGA[;(UV[EcF97e2H+]Q^9?G\Z>f:#f\B
c/9;YJCSWd38Q1La.C/Z.J6SN03E@?,aS<c6^Y_5(b(N^d&/0JH;U_V)O\.8K=@D
(@J/eS)+>bSG48Ced_@B6;E7b2V?YJN-Ef-.:[^?E[]g3HeUg+AY:R;9>cUB.&/T
RN.c&^2B1B[UL48Q@J27]A^ETR(_,>S,\_7aXgH6[-9OCLK0\0;9N0Y<1b1<;OBB
g-gVaI)gA?IK]dGCbXWX(b?J)NA2H]\JX(cg;;;+IGT0bMSW135cI?>B/[(9@/-<
^@P^5_bST1a548)M[/8;J(_E7aTb4.0P0K-S3(gA2:]A-3LO]AVA6:4\TX#C0TT\
S+I:^a_@(8]Cd1Ve8(1ZM(\KZ9A5AJM@GPB7@[cAI0Ue/d0/cdG&?-HcY1fEf.1(
A=XPQGDc3:3GAZ/GBA\HG3CGWEa.:TIg);KfWRCf^[32K,_HTb7Z>e(d5Ma&86&G
KZb4<U/#\2YL_N7^B4W/(EN)8g=;BS:VFPfJ4D<BL)I>9=5fA9<^4a<?E@278VH7
+eHEPV2-d@fE]YX(^DQ7V;HFLS<->U#WRf^F:=;f&VUD&gF4gBOZSDMK.,X,W>M]
NL\/DLfLXUAccZ&?AM>#gV81J=KIBc0<9.>813^C#K)X9ggeI#R2<,?;Mf0Xg7#Z
0<T232Z4WJ;N&bFK^N5I;OTK)\M)\ABU/,/AbTJF28bACD8A)B@,96e?.)e61BG@
_db?M+V&O8I)f;>ROZS?Jg=aYX527D(CRL0QbG4VMSVOS7-L/PLTY;JbP?^?4cDb
(YPR6#?&9F94?a,VA&0=-PZ_;J93;Wg\5gTHP+Y[_+f&Zf8fB@VTgMYBXa[<QA:P
N2+^2T8>/UDNW:WCBCFeLVQQEDRMaVDEM4Z3f^XeCMg.UAO=8LV@3<F/-#b07CQR
)J9JS66RY)HO/FKU]):_X3#B20:DN&#2b\35/>eB5&L.a@#?0&d:]A@eC21/O79d
aYf,O#HdRV5WZ4K_D.IBET]17;X8gWbT,C179dJN4fU[X(<Ce_:f7?.O]E47aO?M
ed?+9NOV5N,=11@B2DK.G/.D?,fg=GDISB>>UV;a;0O>GZ@f.-LECPGfaZdW?>=5
c3B&6T;:6L2LTc6++JfY6B[TUdD<\[F^eBb=-:35]IY)De^,[4,JH=X/a/H;aWF8
QB:)U6W73:ES@)<cIY=XH\6,@Q3E=aa=cFHM0F1S5/=DHdQ3WP24(/>K9f)b.T_/
^P])381J4@FU&^(5Z6)gM:9Fg[+VPGU<G,U4@LR@G#XbLQ6B?D8eO5H6/IGfHP#,
^4Yb\(\80FfVXQ,_]M;b^KP6/CE7G]Y0./(AQeD79&Aa3[6:Z=T6\G&(([:DB/>0
)(1<.(E4=1FS?U.aO84B629ee@X0P8ZSR&MSEOXbB7+\\(<J8@b&MS&DI3I]<B:I
Y>WDX5g&gGHbSJ:FUH\<(:b+^L?fL0X+^<&)caG._bBQCO94.#MgbdX9@aRc.-XM
N83+4424=3H)d/VVCP2Fffb9V87_BQH.Z:Xe9I^O)P4Jd(#)\dICZ)7W6KEJ2:_9
Q\E_a8TO8[J<LME1\Ef-#=#NG]d.:[QPa2FAQ7+\&4Hb7J-/F;8aVAR;/?&K?0aU
_SfIW:SZW5]+6)_OTGTVW)B6IQ8f@HKaa=g0_eJ?>\e2/MN@WZ/JVb;Z+_)H>&X(
ROHUaT8)\;+T0bD6+IY[,4//B3gHUR^c7g6<_d.c8KXLA=ULd@^L]65-1&,bU[\J
@&&HD#@_K0U&94+dR.7W/-cDa5F6K0-T+fd-Y(<.UZUI>\TRO,AQ6G^JPLJ1O#+X
70]J\_<(2-CcGO#5[EU^U6[&f_g##1fYZ2R>(I]&OVV5),U\S9R(#ee[=M:XV1]_
CAfN;64I/)P,V,c=ABTf>(BR9gJ9.f9Q@G:fW8V6D@[<:I/58c_J_E:K;2/AJa>,
-Y[U2G^EL2E_V;#+?:3O-eDG@<eD/@Ga@#SB0._KDDNb;f4[e&4T;4^@8T^Rad#@
F]^=D/aSFQ^UODF9^D0cR0f_9@C@KL7dDN6:V].R=2Q^\7YgQVXEN&30I_P/)P;F
H-)ZF9>4Xbb3ND(5:fT?gUgd#CE_^\\&UGa.]RgAc1HPT#24K-GN.=KJ0BTYY4Ng
,J-e]\gXRO][8a=T0ILNcAX:,<B6CR]c_I8&#J=VNY?RL/Ze8EYSOg_T.2SJ<dBV
3&5?HSNNU1KMTVO2G<aRZ=+AO5C0JMZY--&-Z]FS=g.4BQO/10/VcZVZIf?89PGc
)0Hc.bV,DWF?S?9/L0M<K,C8<dH08W.e,&C#>/2\U\bJfFF>BI(=39DQR:MaJ9@=
cR;C:?Y5<P&9G=5F2e+QAYER_A,OT<G_XDE5C@M-_X)]XN[C0JU[BT;Z<(I_4\SR
?^VU.c[/Z\_O37#]fd4OB.(?g^d:;fOI-(LK<BZPP24\/EQH1MILf2/OZY<FQR]a
SQ]XAe:g_+;7/VNgaJK-9-eQ)A0XEg,cIaaHM\McGb51(+bI4QK-T,KI+YUe@S5]
NQ(Q5L#SgKFK=ZG63bL5KUO\LZ97)&BD=OM/S;XG&4ZYcXCS(XL.@Q.>aI.SD.N_
58_N<bJ)&LT>+,baV5\.2VT7TC(^KVgX>?[dO])K]#Q+1^BBbSW_OgLL;(9aLff<
2(5F;5QLU6PL)QD\WNfQ/Z4A?;9F[/XN5I3gZ4>V2\,DKB,13bZbQK\O9)7Z8Tf)
HU>PdJZC&,C@EU3G#R+GS7+@5AC/D-c2T-:YU.HX<,/5;H[VdOXaC=BCECXW(W0a
/eT=<>_-JE^QgC?Ee#[)7LSaS<TJ-a<Y3P+gQ]MZ&MeR(.8fZf;[U;&L+9ZgDR<D
gf38bWG2?2YQ=4+J-QTgHIadF\PF):I/YEE+,gfBc<X?@IH6IO2YHHY]6aH4+EFd
K>cA/cb9SOf=LTA]M0LP88@;TRUMMP2)&b9edaZ&ZXaUgTR2Zbdb?#CP?a2FM:f&
1^?:?cMZGdeJ=,abKBSF#U]^.U5IJdeOE&d5VAOY25g6>9)^[7XQU_6R[_#XY:#_
)bSe;W_]]KT+G)c4.?S,3IV@U:&XcD,?J#8PfR03P^:DC\g?\Xf.Z9K3M)LYN)f:
TO0>\(Ef4WBY9LK[f0dgfI,:IWG^8^:Z<O(e/A+(P=EY])R4;OSSHVYA@YG02-=R
>T9UT:@3D]WNVK=ZZ([_>0]M,dD=O<NXKa)HVdZ_/HU1\@2;Z(ag=5&I53FOC&G@
X@bUSO_e,a=,0XMR3<8gD9ZVbgWaTH4SZN<W5NSGAd-U0GIaB\:gb7;A/47E>1PG
4bbaT1e6XHPBMV:\9bN:aV/#K9Nd=O+Q(VA0B:X#MHFbM];c]Y-f+I9?Pg6&0.95
FF+-O3MR9+XLU;NgC[=B8B>K2?@I6Pe8S73C/F.\<YEY?Y:T9IH-R(#RD=bg/7NR
BY#UTK?\)LZTgOAK/[_^VcOQCL7Ef\QH._SFd(Ab3)Q446\1:HY=OP<(3g]\-gaT
dI6egF7f&B_X\E?RM8&<A7\6?FU:M(<Acd+8ET.QB@G6Jf,2Q3>=X>-15173gKVc
[aK+QEVf[6:(<L/1;6T^X8&WK#f4OOgI5K9(2\bPeNVGLN10=,:;,-ZdS)+ffJHY
I>P/D^1BU4fQEeEG:K7QcFET,O</@&a_CL<QV1&4.]?9@_BS&5V,6Kf-/QK_51Jb
VX[J5aT(dIFU&3ZDN4F9PJ#UMBR@G]>XSdEg=EB)8ZB@4:bFKCf66F_::#)gKZOY
.GDa-42-P@48>\:>bE\:f<JF;\O[;=Tg>B9aNg<^\#[73;-^Q+Z:HR(E/<WG1#36
X/UKJ&=SHY>ZZU>4.\HQZ7>a[P)H3Z0]FJ(PBNF-@W]EdO^H5BH.[]AeWLX<52L6
&60U;=^DDAPgE=,@]Sa^0d06T)L3]\(HbFT<?Z3OZ8VTcJPTb-HQK]g;5\#1T]7Z
K8=fZ_3\6K&a(B_(VIOQSBK1>YZ2\ZD<[JKAe+T>]d2\PIX23<\0[.Y6_aBa>(OW
I5W.:0D^[DVBC+._LZa>Ma),?N08+L;VNN&Sg0-<,bLU(2VJ4U)b#9FRY]d+6RU3
6LSe3PfCaKb&S5[I<&DaNGIDcYQ:^:b#Q>,Gb,OE<]K.V/d8\#C@fEa^RN(J@57;
WV1Tf-Tcf7.11cR]cKE)dC@\@<-?:Hb[L=[e1\36cX,O+e++QK4:XT;C_LQ#\-MG
S:OUHN,c#GG7^:Ce0ZPNaTD(O(8I5g[C)L6RS3+1;NP<91PJ=]V\-Y>)+KSf?M(>
(Ff;4)]JEOFg2gT5]C^4e<0Y\A7HacKc;Q4EX?68C]HLH]_Xa5HD3E^=J-8(_Bc0
E<3>WC4:D-Y&#1EAARL8.eUU2WZZ:.:ZV7:6bD:07VdQ3OKaNRWGLE/0R?-GcT#=
7HY_?e0R.I7\b;XM76.^C<Y_]cO0>>Bg]IM389g70ETHTG^/MS2[_^CM4ePTe0-c
dU<X:#g-.>&>3dXg3P1J(XU@P?2U+cDY=(4-&UHLS,>dUcB4H+:HVf[UR85/3IZ\
70f@P_Waa]D#KS,6BH2J6RHX1CAe1/^<+.<U.d_.2E&1F4MadT#C:5U.?^NAEW(U
/71e1D4]c&EF<;(I33R#+=LZ0&/^2.ffKeQcR3:N7@E,W4^]8-[aV1B#]K_7G<\Z
1Y7Z5X=f[efN[P/Q\/28K.F)BO@W6g=D4\@#D:]?PbOQAcC;_R-<>5F5NBBQYKc_
]1BI<d/43b-1RJ\1@L-bfcV2^G4H#KTW5KZI6c>.1V89^\M,Jc:K6Y/B=?dfU.@<
fM?PHcEI=b#bC9.)5G?]B0HcHZCRR>fZK9ZN1JQeWaLfAS?g,bUbY(96G<OTHP9S
#H=^FY3a&SFA0IW(FR:\D6C.S4AQ^)+-\H^b(@VW(N8U4-fK0J6eKaRWOED_GOfI
;YDN9=H7Y>3;4c7dCL.+C+OUeM@?==@:Wc,g+a07(g8[WH1^N4cLd=_f3Z^\g#(W
.)8\f(@U;\TOS3IdLJ57GPLWQ_\WR?fR3e^HEP8YJ10OOMeHX+Yc8gbg+8CePWKd
B+,Sd(.^-4F+-d+aXU^I[>/=edCAecWDA-.d&I411EU[:f?2(RG204Q+:S^4_=5O
P=,EW:R]?A4#VP=f;A]QZ_O/^ZeZ.ABVf1W4.-XYNN0?WA#;.G&UJU,9PUKeI(5/
DbcQ1e/_bHJHE?8</9ST><gb<?8fRQ323R&PaOX6<>O,Lf;S;BIAJSIX&f2G)CU5
CaI1;Xe=d?:@1@S5-97-N8T)KF>e;=\L;E9f\<DMX.:.(QWgW2(X.,SZ2WLd[B6G
YRG#E_/MAQ>Td,C5?2=4aDH,.FGP6Rg9-)fXcL3dRWT2Z?Y<O-a^S(REC.7(CU1a
]_f^?9bJP8[EIHC8J09XK<9J53.]XJWV5TL7;F9D1CfG/f0YKIC7\8E5/O7e^a?7
Q(0XcW5>8[MLc7b&f5Yb(R2aRRd-/P>>gL_[_@;d[P#I)T)gUR.3I6J7G[YDUHPd
6QGa49](3g+^51(J9-+&SE4,1(gK,P.O[+XLYZY,&,[KH(&B[7BXHO[cfdf]D.,C
b^/\cE+6^dN<f/@R@AFV9YBA(LEQSAWX@Q^?X.B-a(NX]WC()SZ?=_;D)V@b_R+.
?B.aLLCO&:HIP][V4W(O)+aa\5K65)d+?c#1EF#0++S_<+DF8T66A?_EUg()OBTO
RWBbOI/;Q_C<<Q#fD?59Yg)>bd^5Tabe/XJa6BB.I/D^Q2NV-3XINM6\RgOc-,T?
2>_G:Q_b^HVJQNd<@M#=&aHH<.]eEIb_Y<+8TAYAe6cS<92/_F<B<X<)W_FE5P^?
81fAG5gS?\[D7-?WDR#XEE29G&?--Y+>]53X<d/_HIK1B?gD)(B).c?EW=/&_Bd7
(AEPZ:M7-+__aLYI6OMX39.\5UB<98_6LZ555VJc6(EU+)FO?c<@E&:.\_+A@O?e
TeA<X80VBY>2MPBB1]HBSb^?\O+OdMU1.LAH-5+0=ME_Agd3+[Q6XY5^9Yg#?9=A
CNF@dc7_:#MLEB,DXF5S9E&?CW?;UQ;2NFPHXW9J8a(#DaOgM(LZc=CXK_L7S>[>
\b]6cURf5CKUK0WZaU)G^bb,>Y82<OW>@6@NQ.Q_9UUfaga:G\[G/1+M&5c7.MXT
9ID8R.WS(OLc?+MX)gFJg6c/;E/V_-2PFAe-bWAAFAS?G_\0D)VLEd?47<IHHUJJ
NOFH[4b>^/&Db[Q.K;@eI;N<)Z2MPTgDId@53eF7YX2JW)>.5g/^S[M]-KZXfU.E
/C)K^WRM]_FA++ICQ_:QdDA3K)]HUR2Q&6/#[=Q+:#NW/HSa27W?7,ME\3\5JY.7
#>c+:/#[W]05e8ML./CFeQW&bO@<<(Z^f37eM@@-M<?2>HZ9RGDMd5]4H5RHPZ,2
3fCXN29?Wc]0AVN3a;2P3YG_GEMaC+&MQRQYV\GeG0YQdPVXa.0S>6^cKf#C2OV.
MCWLbg3HJ?#>4_d9.Jd@f1QY<FdM=dNJ;.1ZS_.E/)8=\OJ2V/)fP21OYU,?)B8L
YAKB_4<XS<:XOBfa]V.QcP:<OU[6D,F2W6@/XSN/X18MaZL=,XS1F9c>73SYGX/K
HHP:M&\gaM;7XWQaHGZ&RA_-Q49OI=2N9fd,28db6&aD9P/f4\1f8NGV-H,d=]L<
+[V0U68/7A^/9TSf<E?e9ILI2)Q-D;1(>1W<FWV9DJV@178fX49_a2c]),,^XST-
7/KWRIJ?&dc7M=6,8QG4AEfZZ4D@(YCQPJ-&:+-G>Bgg28\MbY=5+5D9>#@L0cH_
d1:N>)dXFcc_CS0>I([Y;R?[M,/ecFZ9<M3#)(TI3?aeeJIHeJP4XA]:#GQaY7_7
]OZc&8.><&MEa=DE#TRT,]=S)6:5BB#C\JLLFX)YGMcV^f]6I&6^FDcZ+JFK3_Re
E2?Yb-DJG#Z<RB[21E^SH9ER,29D,+HG,=Z_87.Q&<GKa6#<^b&;P<G5GM5ZFK&]
Q#0V.MVf&EF2-KaR1K@a9<?^EPPDL&Y+8JELHMI&R[Q,D4-bcF+d[cN20N.bHTeK
.aYNEXA0WKBH&V@SA?-T.5#K4/G:VABKU?0&YKD5^7>C].f0NG\+SLEcXW51+P+)
gVM3Wf2?NUEQQdb#gJf_>S-0IWFODd,Ag/]NFE1+.H0PBY2T1_E2T>LPV5af@g9]
1<fO1@AJQVdcEc]GC>W8/CG5NTV^0\[EZHG]S0G8N\8MMJ_BXfeRIZ-9GY/Q@U?2
061V4]Y@Lg7Xb3Yb4;3gOZ8TX7\T0P,1<,A=]a+]PKB?/?DL-QgS;T?[G[7JG;:V
+-JQOaFFADQ[F+&62.aT4J=B,(-TcYOS_IMNb[PIGCQK?_>8BCR_g22T^:5b^WQ8
[IZ6.C=5J1\\T06b/-cHNJHVL&W#U7H?eJ@/9EdKUU\.6I-d?=@37B<.a\@3MB#V
=DFR;R6_FP-G,VB9GZ78f265O<O\A]K[3S(LD53G;U[O_QGF7Wde]&\.5K4XPg.K
<&N6[P_^7_6I537LT7]EB6<O=6.Jd):TT^CU3D>(&U4?,Rf@NZ(Y=IPH7JW=PJV0
(;5/3PP\a#Y7_,HO\H,_MB_EZ2:UGE=7+O65X&Y(@=Wc1;IAE,72&cC.I8,U75[6
eeQF7dID]K3=/NMPKgUgdU-2)V/.]0UGB+/U:+Yc1&gKITYF/NCLBfH4F6>IBIb6
2.R0Z(N#775eIK(2ZY&8S8a0A;R-G:2dWA,LW;#X<NK+8VT+Zc_1E1a@^BIFRQdf
X35<?_C4a&P/Y8:L_Cc=W0X))XM4V\IcDHeP8#9cM5G1^6C3/)c7[eH[&PH<baW,
;1Wcd7YDAYPI020ZT/#[2HgLP0EP8O-6GeYeef6)F/&0<]d^/d3G]b(cTc6=Vd2B
UGD-,)&dXZUMB4M75N6Da=H>3>U+X2K^G@J#<6&]R\OT&3Ob:U-f+gdQe+a70c1f
=0adZ_-A?&;UJ#8-SgA82NKa/TE)f8bU7_eRI_J>P)gR6PKHNKL6[3,M5@FVC&U-
,V3TfKSZC3XW\>W-ATUAZ5+aCUE8GdJ6#fI<6RVBZQMM-9G9=NLBR4IMD/2BeEd\
I53=LLVY5;82?QcT+83VTL:L8BA2EL.8fYYf1A?XdGQ+QgfMJWRU7OFEeU_&JIRW
].(/Y&K0=P=?6..J5RE5]S-5LG,-RdLP:CJ[J\:ZO@45+F>[F?Q?J,9e[+DB(>53
9Sb,cQ\(bd#IH,?>[>(3)S.2YIW<[@+2HO5_>.]9ML4-722W2;eCXW1+I:@5aA6T
P=#g^;-<U]Z6_&&#B:52Aa^b[(.cEOIVE;CB4VC&VR/3Z:8\.4E3eN&,LJ5YQf#(
^\SeE\d6PVD:NeIQ5V>)NZ==;)#2@V]\^?c@J\W#C=I+.c@)_I?P(bHP9U[2H:Ob
YDSS4JBK^A\^)9XgH_MX\0X&LJ4Od_270V&[LD7M2+ef#EIW.N1/.DVAae6a,M\f
ff(M6\5C>c8?]a@HT[/ZLfbA=6E0PM4,1X97HYCPH?R?.6A+]e/L-d5)O,5TN:E/
12a[5>AZ[[f-B]XW_=^\/G+2U<#N&dM<)QLAM^:I.0&7-Y=)FW/XC84HX/b517B4
R^L697-e=<.b3C.DLS#PX[eg;Wgg0F3LDG:DbOR8Q_M?4+G\4+P0USM/eKPbLC+D
eQDSMZ/;738-dc@:#Rg[(2N,\eg>DM(8B1L??RJ-WfDg:Ua0e(?E2+7H4KM(B0+/
edVMg&[R,1_XF,)0+Z<F)aQO4HS>UW_MS\<_&JfVU]TLO+9U/Id/2Z]BeId^cO]]
9A1ABe8PU/(=SIDW)20,YdZ64I8.L1D@e.FO^g_dV@P=HN#B3T#_9-@,-80<a1DV
Y8R)_>62WP#5;cC3SM00]EIV,+g]Zd8BT?B@L?:Y77Nd3dLEN7fC_Y>?A28(LT7.
TMg#b2A^/KMXC+EC2(.4c[Q5L\:efD[Z(^<Wf0U&=>@W2T@TYT5Ad3E.4P7@>f<R
W@e<gSKZOQd76A&D)S,3=A/HCB2)BI9ORJgCg=]cLF99(NP0fdGbA(Zd2H>?T@Vf
@^TNa,0SKgEcIEQ3](DN-DfEYQXU3N4WG:E5Da-]eFZ67G)K^F)d#SN4^<8>N8cO
g]bOd#9?@gQ7C)QLQ9&e>VB<+E3?@9([EZc@^9B:1LU_GgH,J3cZ8K=Ce=)C:JgU
JeV\Q8&.I-,\8TF+eZ3@_XK00C7-g_QC3ECR/(Gc59W=-a&43TP[CE8abR:<NM0;
ILW:5e[=79(Xe823Z1188=7J]=0[^gGWBN_Q7+@C[Qc.F::?<;/EdXF\_?X1He&@
BI1Rc&>.7]BZ.63b5K3^Q1HLR5</d9eg[GNCeN204gNO,:Z_V9J)&8V6?bb?A4YB
;4@W9E26[[BR]?12bc@eW:10aAG)Y+MbW7H-g2f4O(;]PF=\SJ]V4S]G1MK5NY:I
/66/5DNREYf;NR5\Gg9^Qbfc#9]c)Y#UE#,U;90\9V#G0A[]?8Dd>&1fW,A61)@P
:&<dZB6#Q=/SR[#0/7>e2D<KG@^]Q_NGMPf80;c7&UA3b^-^XDQW3J3[A[.@N]d&
^&[IJ;/Jf4+O59#OV_X6OM/SJ>;>E8Z2#H;NE0FNE,EV+5HGYZ.MS-^d)F1Y[ZS=
8.^>S4>.H-\.PFFIEM,2FOabU4H@0]7CfH1#LDZ_=+<?#4C4P2,=UB?_9JT;V3/a
-4DgEK.c7SUQ3WEFR-=#/:UAI47d8)]LYAASP;U82&Q1JUVR_0.OJQU[bZ,&:GX]
XAUeSC4K8DRT\eHX0K1B75A#X-LOEZJS86B<2B(TX@b#feJ1<HE?_\5e-Ba__U7:
)03+9a5?9NKSJOQ3?NPFH,N,-VVQP/<K(b\=)K7VY#ICH6cbg-P37&J<YR2?eNDZ
bQ:#gO.AN;A:.d,FX\1TEc/GSR<NQL>?=Q83F/=?f8EeI@KbL&[\g^dM?BZ@=MUB
Z+XdG[Yf5TQ55O2V\bV7+S&F9@f4#KW2gZ^TdA8&-KQAP,+5&VZa]9+.+3BWGd(4
1FVL1Z]JKRaIbH\:7WK5LNY=]^ZR0@Z\XTZCc2C9eeXX@)=gJBKTDD&QcdCe0904
BQ0W2K@S&<\2c.&1A6]4E)_g0d]8?fc/9OXY)1P?QeY#+3^_&P@[]:=aEB9;.,NG
\b+#RZ>XJ=Y/\XPSf/bH#W(#<F;XQ2^T1G?RA:Y8]Z4Z?D4a,ESSWK)[HZUGb_U+
SSD.?:;N/)RAc4+?]M<Z0_6Fa,TQ;.#O@_dRWe6g1#A1YU5KCPY6.@X+Y-4C5#2/
D>FTZO.^cI(@-f?_:\_1\YGe>_>RY6VKY\@RO=ef0)MKJQR4=+(?U=INO)U_RKER
Y/K]][H<e8-c(65,+/f.-S#P+NN;-;)OSUfVUB1UBH7WRQ0^Za.+fZgG;\;9:-)M
VMQPAH/](8]X&g[69Y\FU&^MXD.eC7NVD@L?D.S1(7((eX/TI5YUdQ@5C\IV:.F8
.MP=Z<Ba0T)(BF72&8C3&KUH0GD4T3XDdE[K3AVHC8f?He>V5)JMfLN1EaLS)ZH-
JJTCT(31.J@e;Y):4?_e5:LCcWSDS.RFeA,<B.Ug;8dU+M7+SD0FX41.9GX^MM28
FA+TRJPSde,L)1NG55c/T:@Pef^@_BK>;L<F55=ETF+R>^,?456eZMe2LX4c?[]O
/PVfD1&(P8.b&JTJcD>;479>Bg_NM2U6gMRO^^@(&BKdO58:M_X(.PM@(<1\=Z5_
dPA4W@+M.95JKF@4A+F82MS#A3Z)B;+7X5KL:YE89cC@K?#6=aGP8G:-YPQZEA6(
U,E1=.037)[<Q=+G=V?.Me]K-5?;2f=H\Z=Oe4I/4U+bC4R>9_<9CU@DAZ/31<Z=
J4710gI<\52>P)X,<b=R+01;B-bGe/F#0P\[6CGHAabG\OC5=T_GM@RMDZWDK&a(
JXR/TFB<9]\aLRLCY7M:S@:fY2E<T>7HU@>U7F[[^67E/0#?gDSfX&FSA2_LB1QS
EM1Id.+9UH)S9Q[&.2:1;9a:<,J@^E73OV^5b_7S5V.&EY>DHJ49T46]OB)/TKUK
2J,>(g&QXFZ(I-JLP56C3dg+?JTG=d>;.42bV:FSEP1-+_.>KUT->)V#N3BWAB):
]_0SaR]6UP3aD@8@:f9OBUBg#X6BDNY0-BDXYIJP60MIE]ICg+N0FBN>g/0W/,eO
,/)?JYO1[>1Z64.#U-T-_D8+(,?#8DcW/CB]UOVRgSAUWXLcYWY&8=fA=@U]bUGU
DCIG9?WI&O5:9_KXbZ0KC5-BG;(=,<=U//Ue-<.U=4.Qce7H\J_@Of0T>[-BISKX
2L,?d9H:8T(1JGMEG\NS;)3>HRa63fN:220;ML1//=+/bDVC?HW_CG7SbKIS7#^3
\977D,&.^-MFYde)^>dU(XJbRCCWR(?d;HHJ<#cKWFKIJ0=0\CdC5TGeKGK>Q_(#
aK>Xf)E+&)aKMK3Hc]YHT0MCB+_J?Y0E9W2abM,-MJ0B;eU>WJ]Qg59#1b43_J+/
(A5^A]NG6:CTSJAF-[I,?.Y2-B]<T&@Tg20a\1c3<\,XPbW81/WH98G8Gb.g:)\_
7WI9eW\EGXASaZS4OD43@3)\BP5#X[^M+L@_O9b(L);)fe9ZF1=,(A3Fe:&<Ub5L
d/+\<]FCJ#G5VOaF\1EY2/2ST75HKGNBgaQf:Q#?fS(-7C9^P@EXKUOf9E>7#;E6
H2/AAZ<eW(-4:9L,)^=0JFJV&&db)?HI?CR=4aZ\=R]bR0RN-2I;>1MUZTWe6Y#9
=SR@_CWJKX]&-.eCVJZ^AeBE(?f1@CBDOX:ECRI1Y;C=)e08J)5MVW.AV:=(D-(0
3&?K;bUYW[8f>YeM9_Sa.MDFQfd]EOU8\)<C:PAN77?FWI1_1>WFe;gXGAG35@K=
30BL)(Zg).W\/PPPP0e7Af&+U0gZ.\F:W/2_.ZJJ<=I83\(KJM?dDTC/27dI)_+B
b7/T[^S3F;O=EZL-4T\4e0fQ/R<[PLaLP1EB5M,[8_W\DW0:)D601e;SC4a9)g5S
L\L19=VZ0aV_93aQgZXWC=TMa@)cQ=3ATR<W.-2a7fI:(+,:X;T100<I-Q<XA_39
g1#g<=H4RZUPBd2H3T;cM+\I2[4;>2e0#gR\WbCGN<;\eba@V?d@^]U8d)QR1-3U
HH<UQYJNW#/(c6RR?19d)N8JB(T8\X(XO65)7-8HD+76ZQN<T41U+^3PNPRF,#X.
2M^O,MHA[>-b+E,H(RJ9E9L6#Xda]NS>EZ-;T9AB5>\IUc^UH=CbNDPbPN[LT8-D
^=2E^?_[?WS+e)+Fe)8D97XI0MK6^[37IEK7E843:.8,F_c=dFaC]V/9K]<6F(ON
AL?6fGOL[SE3J96,8[2DST/?XWLLIbdZ1IL=5]M+TO9<H#0S>GJY6Dd[E/.fFSO?
fP-c-E22P/(5WC4QNG3)JLdPD,1df^AOR\,a[&@.@)[aY@O0T/FaM5=F<FJaI82^
VETA<GcY4:b.aW-YR2YIO1T=2@/KRe3JDSN\G2R[0A.WRE@5BbTEg@6dN-gI2)@V
SLJfJAbZ@)aBVQ#@08RK_,B_Pg1McI/WAW-C^>5g/#4<9+?:6Y(=fRJ<0<.YHSdV
LH]S5C69P]AK?f?^PG_Z>;.LHP2RA(1D/;c1PJE]4T2]/Ee:88P]^b@5<\9<M1\C
84XSDdcZS&e4@Fc\5::3^M/YgQCSA=^7,ON52)NBQ)/968PX\Z^-==M:KA,I&Yb/
(V]-@#OfGUSSP^#DgYM@Y9fMeb#FMJgMPU]CG?BGa;I@^39.eWT6Q:f8aDfFV&/e
.)EIE6FOa6=G_0V[78[/a,5?QY6TFF:W(:.]8+GAP(^fdSE)Ra@F[WK^eW=.W=<?
)?[;cN6+f/f5_0?[W8bAVPEYf&TDJVe0=^&#AV7cS9JOO_9:e=GG9[#73S,0;e\;
I2Q.UCYT&?09a:,N]F@c1g&SC6e9c2=EW>)LDO\I_[P#W1cB<<V)fd93>b0Mb4b-
UW^FN)bfKg8Ka_&GV5Nfc67[#=f5G_MI]HAJX?eQM?5DAIdLWNXG1IZ_eeY-?J.S
LfM_fX2)PC)8O+d^-La]NBFZ_C_7Y_8-[=c2[a>UC7/]G^PT&T:7f,GI^BQ&UX()
R;#[GS(RFKZ>2Z5dc?LH0-[Jd[S4Z;]?-]U/0GN2L#=Yc]K):(WU]X&]A)eTQ/Vf
AX;-H-EJ3_[^6Q:&)c0MDXV0L<L(XK6=eFD^2-E4-M6eaLDULd;]8GcFcCAV^b&D
^>[Eb&VC]B\d-1-_7U=&5Z(#;J#KH[&@07\Hb?=ZT]]RKH4,G>.-.aXS[He9gSKe
G+Y6Ud#Mf^F-4&CBP32^F_DF,e?f9O+SZ?Y@H\=OD]NY9JS.7J<Z)N4B92OeEOTF
]d@9.Y?7#W7+1QDGX?J>Nd0K5c_YV3OC][dY3Gc#(W:DZe)[PE&PNZe9O?L<GT6L
E6#C5DMWR@&MB(@X<&H:YQHLBB\I2;;I5P:GD:bgGP(T0?5<0U^eM2=QP=IS2)b1
+6>(C+f,dY>f\0]Q)1+VC1JBR^gG1>ZRFO/8N4DbGA10RK0UI34A.^dY50M4W3_@
DUIY+FP0>-7]&>7;7N\UDP-\:-SIN1=I((M3Z(,c?IdQc.LZ)&IY&^TV)@FZ4a+3
Oe6,TgN:GD17)Z3,&M@B]eEFB)00Gc]((E7J>cJa3FS,=+O.-G3\<_FR#F8/GX_@
/K[XS@U+TK?TeO2)e/J<=ZE/eW_)EQV]Pc_BXJ/N<(4d>WJ=XWM_;-;;5/7@^)XC
d-34J;C6VI0Hf:I&.Y4;=T,LZ.9[QSTY/.9_)^fS/J95A#[aA=6DJXYTcL/#aAb4
Ce<C,=CT8VAJ1UV>]7a2:>LUCKM9Y,J]2Pg&^\6I\HD>O0&:1eEBf9\N3e:1M+N,
T8@T#Z=]?O>ZP@PDf)^9TAD0=B+/SZX\JY)GACcZP.S[0dTcYUJB5,QCJ.45)6f2
.W9R\/9=]Z1DC/@#]M)?_H=3>XY-O/@@?)[/[\+G]OE#_RM[:81<06)bgF^XWCDG
ZQT1L2Pe_UDdEedH(N[.OgX2GB4Ba[ZI]d0CC\9bO>)3;113d1D/CNgKPK4fQQ@_
>P7FZUKDN>=37UbA8_@XL,<UVN_]5DFQWNP&e#?#F(b3J06@0^Wa/EXQUIS[1ELF
YWL&66Hf6,JLV0N2+_;\ZD=+\6U1M\-3Wa[T7--.&OJ[:K<@72dZ>G9(47UHe6(>
[NK]c5f@@XL+(9XM<<Q1GG1E/KF5SNN#B7^I1_GW8a)<=8a^IZ)B\U,0RE0N1O7a
5AI/0bA4=C,g8\LgAW6OI;DN=VX\BWO#dRH3TDJ+(VCG#0^=1X8@&J&R><F[(V&4
4b4a&f07D-:CXd@[2PTcb2U[(E5f5#)B0@ZPL[]CUV?+PL4PTa&\RL_W=7@64)9.
\]/=#VXWc&C1\QB)JO54R0:YaZ=eS>?-Q8YC<4,QW:;\8[Q)=@8\[64aPAVWMcKG
YU,US\bPO25bg=gS#YD[L([5d^Ie]dfg5]5d5;D9DfSE+.g3/#K&aVF(U0H3?g,U
0VF/]7XY^6A)<B>MVgegCP#b;D?SKUeUDVFT;,E)MCRG9>E4-Ge5U;E74,Q>0SD#
CcYZT41_E4;4b+G#L34I]2bJP9DE^XW#(#a2=g5TB;#Sa[GYY6KV6L5HTT_V+9&9
<MOa;&65&_OdS<5S?O=e4c-_4][_<E93>WM^LCF&AMS:JL;g=40DADWcZ>fbK2F9
>2++T;67#TS[#9dL<]:L3R]-M^KK1M,;.-O^3Id9#5KX[d-]573JRZ/#?JHaZ[f3
452L-\JO19EEZHg-_S^Q2RZ::7d?]GK6E;IfQ7IYB6@DeB0NPed+U^B<3<[HUEE-
U_+I3>\Og,f[\IKC>\B3bJ4ZNTg.WGd>IA(1+DN[HW8O<PR;=\I8[YCQ,#NG<FIK
9<\+1N[_;CP;W5[/=2QJBQGSW\U9X,7IG:Yg;\=X/Q29R>CPCSU6f:>Hb5LFP0QX
bfeWF-Ae9a-1:S/JbN0=3(+XHF#S+AbWfH+C&f/[]b,.+9G+4WHd)U_DSTY@9\&d
J_?[S)_841KBPYGY)CTaSd]e6,421TV9/=)b/G.]Yg/21^:1L[E5>V@,e6;QJYTA
BZ0F7YE&NW8b5@e@:GY-U98&LM9WO+#?ISg[X.&8?EKPGZ>HGD)0bK.gXR,/&D74
BT>]^=?.1\G8bTH];Og3IN2+;2>3OB6XCFTLbI0E>.3Q?N=Qg?@Bbf2S2GN49Zeg
c5WQ>S(Jf(6&eE4409:-7A:\&-/E8)&YMLS1:6QC?AH,-U4N<>>X22a6ZW^9;7XV
(P?X-.IDcGOE0OVV[?f1TM[9.f9)JD]_]cfTc;&K2ASdELRG/7H8Q1\a?.)]VL9E
6KZ61.X3,ZbKV)BbfY.DU1M/Lad@)8c+\B92PG355BZUZRQ=;UP0H=,74N)T(:4W
:?EO4/C8[aPJ+^HcZQZCcBF_Zf&:aN:K9f.2Q.;_T--#31VR&XB#76=V97N<.6a8
GdTE,SPe9d?gb)G:EB6#&f_+SXGS2?6JTe5E^:EN\6EAY]@6.YXGF@Va9YQQB\6a
4f5>H5#(-cFI4D+BY\GLdb\[:2-/e&b?T?,ad_WM-CXMA-g2Sd7S+#+4C0<BL^BE
g+4;84[.2>8F6[(^Xb?4=6M8Y4EMZ,NT1/OAZaC34Sd:(=QL:+Q1=TX)]7/N66S_
F[DVO3+UY<?7/,2]IO7UHeeGYb[/&NU3==4b=MZ^-Y?fPfK^;X0XU_HM0#TD()[:
EPOgG6<F)9.H9I@;2&&cL8R-fR+O),=&T=,Z=5Y-&PDQT&=<6HQ0/7JF]ZP^eNWC
;WT@B/VC5e<K[JWC:ZQDN#d@aZe;NQ6LSH]^]4VW@c]FCf\I6)M.6K:.<M4T^TR;
-bRSGDVB=LcK39?7Q3ZM/M]4aWa^O9BOUBNZ7gT2\XAb#>9&A:T=&_aK#M4I1L\L
N<4:RgXee[^O^2DQP)F0AD;[8,4IE/c7_>Y)#/e:NbJ@0gf309e0XfV<<8]?3;^^
Re/-I/LEY0>9]59U(^B4M/AGQ)&NZdg+5379Rd64;5RY<ZL3Y;P(BG3BJD9^ZD@5
T[=WGA6XfLS>1dM34-FFXPbE\4VdV>S>I^]8YD3O735N)X8)\KW5YDcT9RKD(bba
.NCYcN2MAB[.eMQ1==4?K4MQ#M161,M?]/)Jc]-4VHd=XI??5+5,QFW[L]9BA=Kf
+d1RCbQH.+R>d/c?^bL3<-<.Z_2>E39Ca3Be?=a_eI14/;M1;HR/GgA?_6M12T-g
K2fd8>;E[=0@+3fCRgYT&C1Q^;QDC\1c+Q=A8(=Q(U]_1>.8bT]8D]GA]C3MPgCZ
8=9BPME8dXHKf78gA?-8\0F@&CfY/<cE)<C_+7,3R]16F(SE3.6]+P\@>,c=1g8V
&OY#YM2@/R-geI_5AQ1R)9SU7&[KFQ:W<B)d1-0-Kcg@\YZ8&5L&9^K>U-@^VGEQ
7MBa?EYD)5W?M/6eB:V\H,_7:-=1Q/R>1f:-TE8K#b3C]f(c2S_cR_VKX&E>B,Je
1.AfW<IDVb^_/=;WPc9QH/2SY,7WcWa1H]-PW83WK5(W6(=EL0Ye/&08(7@AW#4I
../>A8/-c&2N7b=L@FEW/PF#1GZ\-2V./A4e1cf=?F,4U[U2f/H?2.>UTaG/[?LR
/VX:X[g]f^&R;GeT6P/48,9cVR2T98Y=Y?)3b16bJF9gZ[+]fV+H3SFS?-B)_M6X
;0HYb^81A3;g&WR)#NM3O@<_=WJG370\.cP)&<J]adCN)eJ-=/4PK/WZ-L<9C3Q=
W\7=#?=DQCWN8c/&[:TSDMQN7gUZD@UWbcH+94d])RWW208R/WK5A]V.7(Y5)-P[
d?.@;_2YCaA8452@>g5DX&RK+J)LF7-4GVaP?1;Qd;DJV64H@d95]CC,MIV\b9/E
9e]HBDYGc-_g-c5S6Z?-DG#[I)YTg:Y87[CFKU;P6&=0+2f_R.>QNU/TR3I0>ce7
Q90[AXEB+^^+P^dM\-ZdO92F2O+&0)^Nd&W=\A#^[>:MJ[9#BZ6B.G:\A<]J.?44
JRGYLJA\(;M?S4LC6e1TSa_;]1@(GV7:4,>/]G=.8D=AFP_LCMV&fW)1_aggD\)S
[I[Z0W]^9<41V#&^5bMEN-5)24M#-)D4gF-R:H.L0\<ZRK7<I(D/fJJce^/;A_7+
gL0d+SS:ZP(H^LRCV)+K-g/L;(9J#&GG&\aYE37;C]V?GGP_IPW\XVGE-c,+d\]@
dY1Xb>W.A[43]3=QCM\+1;FEDR.JF0cgaCL=Ab?aDcKaN-A#K0+YRTB5eUEMN8IC
+-MFATNWENKM[6L#>Z/L/N9_MRFWO:OJH+3]N?b?Y-06Q56fZ0/C@E-F4EH9a2O(
P]CBX^VEB39[7R3MY2-L-J7@5-#XbH@@R=aY9ZA=b0W.97/L3@&MXb2LWLSV:?26
D)FG.[2B:X/&)Mcb=-UHOR1bS/X\T@;HH7KL61,96).V6cdTDX.\E)Ac,+>W6^XH
JSQcQc00e=JQD<>Q7YR_>FRCcIgDFGVC+@-9WG&NDO)NR-\^GgB@7&Qc\?)Y&Q/I
@:9EG4_6]PQISK]^3W^VE01@C:,?A[0b&B,(5RK3QDFTM^;NVT@]A3Y#Q4:J/>2D
#AH7TE8?]4fTSSZ[QD-K?2:FX,d<G4V-A/&QW78#fO2UE^+NK?(,^M-6C(\(Q@WS
&II+F#-(YdU#)/1K).1c5MG0UM7eTK,OcDRH^YG4bUO#H>960f/^:1-T0E?:U=&E
IP2^6)9]U=Y8TO-df=T/f&HZ6<Q7Xf1aXA_(9K^DJ2CS_K@(PEK0[I1T[IaEbLI<
V)[0)g#7MdS)I0ZVZ20@.HK@WKdaVa.8F45Rad:gI:G55D:+1;D<f89]e27ET/b?
-<1Eb;BF1=a4_7bce-4PbWd_@8#.FUD>HPA8_d9Q;)4,Q3HBd9f=?K3.X4439c#g
+=F2+RS4cRTZ3Nc4LR7/Pff\I6<OHY9#A@c0\Z:0ec]+G@<3RA][V,0Q^=Q46HI0
-e>4M-9=0a;+5J&W#2,d;)9e?C?8B(B0/XWLe/gS_2=CGK+]UfQ7V4L4O+ZUJ/TU
M&96(C/SE>MKZ#TC;0]ZB6]X5T8^[G/?f1(J,?==MgRY]E+QC7<DH.L0:DUc7Z@a
)#)RbO(7,^V<a^1/T)#g7>TgKA-V+aQ6+N&)A6]8G1d3<PX8\<40\Fc.IYf35\b)
fX(29f[IF:13S&AgNLX2C;,.^K6-OX.1b362?WHJJ2A#<J=&C:A9/[OH)7KPUd:.
2F#E#J>/\e8QC-]Q[N,0G_)+YHS:c?5Z@bP([K&(J1.48_(:f93Vg2P2(K:J;L5e
KJcaFG)XR]K2a^bYgV:(G#b5[(gdQOafU[1H_?QW=SF@13A.U0B=FU,aDgO<\2WI
g^K1=)d8FQ_,CCVd&AE_2g#@)803XS4CR52C@.P=R;TJb1I6(5OSgAS@3cW3^YBR
)F1IS]TILB>2DVcRAgEV@0@EKJ#^\8d([9d(eCc1:(C^(\W,62Ma&<4LPH7XJKDS
2ZJ/HJU]F5FC^9Z+ST2bW8MQXQ^C_XY89915Y-;=>&Y4Ece2X]cbT5PbWae@a/+0
Z/]_;4A;#2[H<?fd5EP4>FF;b^7N02]=Q;7g+5LXH>U;=38Y@G]L6Q(P8.c[<NE,
1=3G(0F:WSC_DBO/PY;H4CB-M?0B5X.A<bg76S_7e-LI;;U_,_g>0L]BH;O^b.#S
@D4^=@Kd3][5<d3M31GKg(I-2b:;dcW&MWV]:G<(8?BR.FLaV5&c.LKS9\8d5Z]L
0/[DTW15EL5U8Y<VJb1dC+150AF;S;3&?G5EG0=eSZ:AIg3(?A^=;ad5[R:KCaF^
U<W1;?,<F28NPQ6)>gW#@;.5b<TdP(GS390NSQ;D0^-:G#CS,57]4KQUL>C,V\&T
b73<93:Db9K_1c=,-d],:E#?7Rf/5#;T4;^U?\#SRF6CbOJ.Z>&5Bb9LCWg^PNM?
,999gL5]J?4YFaP8TVN__Ca4,C0)Db\MO+S_ND@SK)7W2:#g7F/DH[Fed@_a)-U#
(81LS[P[^F-UfZ@ZA8Ef>d33IS2I)fODg.EG=#X+0IH8d>0MX0+55/-62(951(aG
6HU=S5b9ff(XH;/EY]G?7=QY.4OTH&aUB_F582,(2\K\7I\J]b:R<I^>R-]fb8OL
.U=^Qf&6GZ+Edd3]a43DeCD.5=9Ac3)c6)4LaJZgZ#@-)S2,5\g_DB?-#Bcd=d@P
fP@X+:<4HQ3[.9GL9O@Q3P?:G^-(:OISNQ9]&75TX\]70T/]?&/JR]:fJ33J1;Sd
[Z(G=W=WRBHU1f?R:3F;X),eG[@([VTcHT\8BZ)Ff^G10.A31=U)=(WV(I)XZgN?
a[9,PB9E.a=@.V@</WM3]QOI_3;:?WW/WaNcQ;We+/Gd=_4<7Q4&B\\BH)gU+O0?
aM:dW9#06:RgSO/bI&QX.L+J2R:M;ZDKTE5(GIb#c&&8\2)c;&2cC3cBBC^(X>U6
71<#R[#Q;f_97e&\C&M2,[BA+/D,d&EJ>EIRIJeO+U[A<O#.)WMGe4.N8\c]1f],
)^bBHgA(E+D9AN<G4+Q@8E,1.O=M\Z@+X/2c\EO(e5AAa:JX523#f957]\H=66XI
G+2dAM2Z]GQ308.)0[g44e5CAZ_[LF+?T47569BZ+X)K7IK8gT23K:eXPH=e6[0H
KCdOB_>.f&>1fEGILNQT^eD[7c1]f@)/c\FIAdU#=D)C4011O/E@[+\.6\.)JdOR
#Y0)c:A9?PSNROM\>gG<d;800:S8Q+bB=B?3_gR:Z:fX<CB4/dBD#3^;==&ccXbO
81R;-5(8#]e)K1WWFKGTK=AO;g#104&A@;UEU-:Z#Kg.Wb;Cb9D<9.7f-1MSb;,E
1Z/[>e6FB9_X&[-K@&SdU/0bWYD+S9E@F)PII,W=>T,6,&?)V\O0bPM51FAI1OI#
QK7QdL0=I;@GDDX[4a7d;e>g=;8dOa)R@<:58+XR=LT#)7+2?_XE@=d^bd13-LBW
ZW,BHLQVF&.Kg7CL1]#Pc;e&O,L<-00/5QQV7KCG)#H[R5=?gD_X5Z^95a+KQ^LB
_7OT(J@Q?P>CP,2I\):=fc)dd-S&]31@Hf0E;9)MO^1Y((4#JBY8CZ4Q3[K-6b<C
JOW_SbJaBCPLebVS^WM;SXLE=Y=#GQ(EJH>3FERDOf<c0c5])O6ZF6g,D)g)>eCO
O,@C?L\YXY]Z/6]V-OTg+eN7I1[CSR=:)B32+^;c,/DGb-CD;(9=-V46&J>[>PO2
3A:G:+aG2\ISEM54e[+56[;<@VR2//J@]bS6fHA;EWcXGQJ[;#=MS1^X2_52.\5Q
b/=^B]_BVRVb6<0NPLa+IG<eC7O@@/A[6R1WZG2=8,:90P\/D3g;R^AF:3eB4@OM
-ME2-8VI5+X^,@2gAXP5KNCI_1=.1+9d02)&A3:1ZB3<)6UA)23Z(PQ0+UL7BA=Z
4,(MIZ,YYERE0;=Z,L<fc84>V)e(K.MR+P_;3P+-1BZ&@Q[UX7I92EH?@3MIL.9_
.F(A^?-;25T>:N,7CQTU3]SQ^RJdGb#I=Z4^V^L>e>]=[BWVf=:[GDTcL\#C/K]K
O<-9U7Z#)fGa-^Gb5-@XgYH0QDBCI[ED/@7&:>-,Q?dNXIL1gY0ZS).ZF/]D&#c?
=&SMPbADNV[]J<9acHc/8-_H-LCYH>/NWS2][f48CB<3;aGe/Q,AE-1FO63HT5C)
+HfCB),7A\ecL>=72UW;<T&79ST7SGRDI,U1\XaHWW\,62b,ZKg^?H9ZK5<Z8RP@
9(YRA/>L-><d#;BL5URc[3UD6&)BVA62C>#7L[.]/\=CHMgc[HT1,.;Y\)@ISFPS
5^(/LY2]?^G-@N^3LKJ/Fdg>F?JFa0f>)#CS2@:KEa,4dC.=Y/Q&g7N;UN)XAd7&
^M)/P->UTW0XW<#Ud4d3(4VF:Ab&6[c<.E_<10R;<A6HU==Q-<+7eONET1<@D^U\
CT0Xg/:Nf025(-B.eWE?LKTOY6@FV0(4J(6_:QZ44;2XMY3/1bEV4D1CeQ5530BN
H(5:==;R_(ON,4,d2N/=A_Zb(fWY:Q1;ZDHUG/5XZTG-BdZ.=VfNRe&eJ7T=-1ed
?Y+P(DPIRAMSB:[#Z95aW?=ZH^^,OAX\^f?I>&Pg:/T7;E?J?.5BPD^]dIaO3A3c
9#0Q]cSH)P4a\Rad>;V)L?2U61BYE9S\EYW>1KLc^C_0KL,RCHN1./CC))\Xe7U,
:?a^Z)Vd3ORQR,Hf1c[;8MWEQ[OY9G=SNgRZXA:0Z-:XHaEf:#4GeI<S:,>&WUNZ
XJOVXDGY_+9([[?DM9(^D?B:R:\b0W#IJKfbJH&Z=J+UZLEN(D@_,EI^?7b+C,b-
G3b)&-P8F4,EZ\O;;[PZEO,Tc-VD[LTQfE@>_7cS0\b7?N)>8?g9I\V9[R5AgU,I
<YbPY#<:P^#1S[+SbZXD[.X_=@B+F)8Zf2J(7e)+ff0,[3YGB=TP/&Yg@A)T+[.E
3b)P\+(&R4e\6X_eCb2cX+M)JIS.\cY[g(V+I\D72LV2HbNJY.3GbYFT#BTW;SIZ
3DHe#>KK05X.^5;Q6-?H8a>)^218S[Q:g&:&Vb:L[;fV9YXS\?]GW_FPc<F5\A)F
;U.FJ54e</E^PW6UP&]I2GQG()@&NIA\S:@EVHAHS7W^5W4UR9CKBcME9bEY&AU,
dUfA[?2O1VO2?4e@&?B>(8>EeP]USEJIdH\)X.6E3aX2gHQ3OAbN9QI]_(,[^a\Y
,f2-L_)7dBLB^??B+@G\f_,&]ZYD?7BUXXd8PHe+>>.QM(_gN0PM#BY#+1Jf\O_f
P@Lac4Ud?f@e//]WBRVPecUKEgKeLN^L8@K]=V.?P0:KSXWCIF_L_]UF+A6>b3c@
?C1PI)XBWR6T>[Y??,X4;\V2C[.:#^\P+Se_X9A_@7&<B&B]=8^7D;E&d1_)\ZVd
SS@H)ANe6>:&\Q3@fF\U\RQ/^1(5MJ)>D>a3J>_?6b;RJFYX3O?D_,TO6MZ<R6de
I3(?]N#@aZQR;=YC;b35gGb;M#G67I8USSY9(<U4K[,f:dT(]X70e/H?S6L9U@SY
c4@QML(d8F5;e?0X;OfDS^R22/W-7#J-MW^R&^-T;YQY[Q/Q+(S[A;fAJWX=@W.)
fOe=/_-0_/)Y(G+V2W(aOGYP>)GM(a(geCb_HeG8:eWHCS63SE=--.B@UaOFE-/S
)VNK<a,@_<\Z;XJHc45:FK2DcbJg[3GRG(&KGfGD0#=PG(00#a:G7RTWV@;H?&:?
XIbV?&?B68:dM[f/#H5]CZX48Db&00@G]c_(3a2WQH_)2^]/@^6C#9:^3e-T:<_,
99KN=;HER;d@PWM,58143b5CY\02^Of_U&4c7GWPV.T4=gUOSQES/4W:IDN[[T1a
0TdcUMX<GQY:cBPL59R9>(NG6X2dN@-,V//,).0W85D9.\P)/WE;BGYdMR\;#DU1
9_4RQ_96Z7DQPC+]+=E_C9^OFFM)-7KY)I+9NdcN;52-@E-e4:AaTP8X,0g&E<QU
?9FP[\TZfD77A0L\#?:4&/4Q3:KA-]F)6J&RRU=EW=.L/bc,8O\9?C(VJQR,E>AM
.Y4;X15=cGHPX&XH5Dd404F@KZ9^U6B#=X<?W/O.YCb\JKee&cC-Id:gY0C/VPgI
),S6)4<&/<f2QHW7PIWIGY5WYEXZe7(^g,M2T,FY&M0&T5#Q[KLL4ITB/BETOKR(
&c_W_>b>#aSJL&9e/+dL;8PG.P@O4@9e^d]\Q>3ae&5)a:KP[@QTWPRQ342:DF9D
:]G030c&F]8KA1-_SS,aZ0a86<@OUDd#-__=g\d3&#ZGEMb2Xce-0XSV5_?@KK/g
f36FUc+7TKBX@ST.(]5FQY__6?P4AG+46g_-RdTE_ZgV#:B;>\(FI/;_RH#(#S,C
_Oeg;4Q_6,=g0O78VbZ/VeMB/d]4G^PI:+4-LSJ[)eDWdLc4VG.7DeACTD7\3[I8
2X\\GR-7WHGENbfFR32EQU#HT4\bVMA2Z3J6ba-1H6T1C_E[dRbC)9M8@7LRC[EK
PEM9gSWSJ--Zef>@X2<KCNNFDI@Z#T@79Q2?&:3D-EAe].@,6^;]J>&LJ5W?&VRE
[dT31DD\86,OAfR:V@Q^ABaL#eWL,/@fW]C5AL;_HN.S:\#e0U=EVU1UF298EY4R
Y9)aSMJD)#(-b>?=#+\J+S_SbA^WOfZa=g&NCBV().]SWI:A[)JVd4(+:DZ-(PP]
3bH)NfQ-aIE\8/J:OW-A8MXAPHHW7#_Z6Z:Dd<SJ\U9/GdZO[b/5e8.,8@8ZED5b
fd(C;]97QeLf3K4<LcG^^LRge:@(cZP>8?d;B6/A?^9P<7^-S)#F(AX-D[42<&)a
F.FR2K;>0>4\,MO-T4I7]+0>P<<.1XPU-WVa7]+a3#ce8DP.KS-R^9974DU;d)F#
C=c>TKf]e=GN&&>_MXdg-eJG[e=C39:a[1R[/4PbA6/6?,G]4(Y_AC9X+\)Gb8&V
Qa+/\BE+(<NM4Y&=M9&MB/(=)=?F(<\X,V,TbY[JfNGQ3bLR&7:N\6+ede72>F(#
U#@@-^ZOBe&FTQ8E7>5eHdM(\?]K]X]8&H@>cd428RI:&Z^?B2OcV,BRMHBb;[RR
cVY<R9]]a&U):d?5T>=.@Y?_F4Y5K\1C#BWU],@/@AS)cR5#&(f:U&Z)1+PYO\T/
RS@D&6FMY/HD,9RFDQB2@NY3QB3XY+4a69U35D.<_@ZZ4&2M?L<eOU>S=:(SCff+
+/W88KD3,;^8;AJ,OZA\<dG4I?WQW6/&D4f7Ie1U4W+68@BD=X9H>(JC8H,,FS5<
2H&D3\.KfB#1-f4]JF;UZZ#9]:.SNR?U+>]RC-LK_OUgEY-01#CZ8M+;^F@-MPb]
4&0^]+-\ODSO81=TY65>7e#6T__Z0BYUV_]R.S&Eg;-,0g>0KR_#Q>F;,aA&S1=I
E0#3+MTY-Eg9(\B<>#I?/6/c;9I&I&cacSM:Zf\4c]aJR\END<:H1:0NIfWID9B-
WZV>?d8:1C&@(bP3;;Sfg,:(>UO.X(.]T=[UQ^64D+1\+#4\50CEDL4f8e</G;[-
_7L=FQBTTWbPJ3CX_2@__-5&TD?S5gc1C(.#HBV4\9M]#Q9NbL/f\/U&c(T4+K.Y
9#2eHHJ8Ga(WRC&R7TgHMFU)/7;N3#G<Fbf8Le+,5G.;9f>WKBE?V8ffI]3=S9Gc
.V9=VYd/Y@A?S:]g/FeL0,L6J)f)KC&EBIfV3I09^T3H9bUHHZ=V57QV-J=(PS_G
-cDJ?-V&#\&aGGRg#OeCeG3@/2<7CCP^ONO1VTDR[6PR6.(=?RE@;eB;P:WeU?FP
OcB@G6/:3gKH?1bC2^L+cWN4]HTfT<H?-WC>aE+]N<EN8ZC.?3Y6=L-JSF5#c+S9
W2T,ZA/=>b_)@/:QH9\S\Gb:2//&D8/.aFN]HfWe4;MScJ]\;PN=dRCVYEO=e7:a
W==5.O@&539H@K>?UZNbaPYCY7c.L(0QH:cIB\OYJ3BP?2L)>C\;>C,HTaO3+HTV
gE-&,CWGXHZ_N8d;UIUSIHeG(2=Agb4&dJDMLE6.)6Z]RTSDVE\g_8+\K^9@GO>?
e8,\\cC<aA-Q^1CRg)C@JIce]MDCE&Q1OG\T_aPe9,ad,I#P6e#D/EG<T0&JXRaP
VL_U^>R4XYfe9I=RM-FU-3VCGgd:b78RgaF.bB=2OY)PbP^c^_4_;D=WFM3O#R_X
&M>#AI.11)T)B_f7-,HI2e#_ML@fTBSMK21I1TGUaXSYE31DFf[a10_6OL=MdaUF
D?H3ba(2\a)78KWSNIGIX.-B-G8U:ZXRg#bK0MeBPGNA>.^MXX9S<PFQe8TE&8/E
_=NJ<PfF&f5H)R5RL0?8_5E2\EHC\1d[-ZF?dS]Zf)L#Y(O7C.=)P48:V&V#fH,a
WfU_b2;[,H5Z@.\>V3<BP=-6cHYB#a/_LaM/F:V(L1TFMM\ZcT/_:HL,P2GD[A>-
>:@d;[2fVC=_?BU6)=gB^_.R,\Ae_:XgF7JaaRbD>RXE@D9G\>[.WM0/NO48b_&a
VOABPM@<98EC3E6RC7BKdQgfJJ[N8<O/DP@=R6DUN@CW,:V]RYdRO8K&)NC78bUL
)9QUPOa6>7+5_IL[?N.J@X/@<1.gAS-_RP:=JA9NLR=TFAb0]ZQUAW(?9;JLJHN_
\f1fcG1L2X.DD8WD54FBU8,LF;/JaK;6c0)0/YaccDa5H]@R.QL1NAJeR[1/UB^1
MS6cfe-D8K)B<K)<FbR]-Y?+4]^bVBHBNMLSM8)fIOQ?S,38B-ZJ;LQ]5KD5e5;G
[:7[5.AP<Q-,a1B(6,LB1DNfUScD#F&;1K2=8FJHYV5Z_U@0G)=a+KSe^8@YA^1.
I?1?=f13A\H]d3&QDP&U\L)#((FPYM&R=DA&WdBH?5CB,4T-UZ4=\9\-2EeRe3@H
0X>W)WZ_H+T.4K(,gW]Ng??;2bB^JX2VR857Q^_N]\?L9L6WM)KPbgK(1V7D)G2/
EUG&/^b>18>@VWJ4/YB\[a/TP78PeP[(FN/=E=OO@Ma8B><1dScd7af)bL)XFU_C
fb)9Xcg8Hd=X#T<:HO;PIHG-XeJK.ffcW;_>]1P)Yc:OO(],SS2\INN4B#074CK\
8?=<L+dLG.W(S+B9D5PWS.()CMTLA?_Z^<P&6./DX8Pa==c7VF5T?=edOS8HZM,D
#9e#&OWW6;3^XGBTGd+](TA83J)-Z<D43\@gBKOI[)A8M<AD0TYZE3F]GWIR&/I(
eKMP?eT.6Sff/c<53T5C\BPN_DIVJ]d^6&/[@PISRfbR8^&fNLcUb/0^#>4fF<Ae
SBDV@LNJH@OA@CR&.<^]>FCR;?JUe5,bTX7_Tdf3P-IDM18e=R0JXH[X0ff9@3PD
YZLV74>Te5Q4M+3GESL[U99HZ.+18##cG&J^TUEXO>VLJ&d#<Ng=A)^&gO>7LQ@E
dPX^abBRFf1P)5AQ]BUCFG6V[GG_7#b3GT.^SAG+0^3&4(X6<YYZ=^KX0LUQdAXB
C-BGG+XF52WBAE(.cc^E,1LUH[IXQUSac)0[6UW,/?Y)@F#NZcf9W5@.\FgQEXDE
@CHV2&(57Nef&AO2A?g^V\;BVR(?[ac2&_X:c^QX:Cd?,6PREY>27CMVT5&5U0XW
U0Z[ZeV-UE/YX=@[:2>2K_]6OId4GR57YU>Z2::>1UW6c&+Kb4e#\W>+/G0#1:EX
<B>A;g_X_<=Gd&E4>-DL3X4(WD2K0dCQYO01BOa:eX<YUf:E(U<1DbAaC]2F2@F^
\,/c2?Q9]cTRJ?-_Y-M#aE=D&PaWS];D00U]J=\\&:/I6HYJcNZWBB.]g52\9XW)
7=[_UFb?>_8VcSLQe24gR3IQ5SQ1:FddFMPX.\6/+L1d1803,d&T;XBZ4_@gH=2c
7X.MDT?-O_?Fc;AK^V<(I11:&1J:bG6b<faeG;@@[0Z9-8&^_=I67SSO@#H\(4C,
&B5Vf#@>J5c7[W4]FD.-gC0OXO+CAWV@B5U-[)RLWIg;WB?6[7)7D@Y,]9=MX4S\
H&:_UXJ83f[[=[?-baJE/-FKT5WFg3A5(T\]d;g9V=PZD5<9;?D;c.0CP.]0+]SH
T)9(BegC&Ja2@EZM)f@c5(BN=@I4#>0,A?F#Uc<eE\]YXYd)C7]8J/QAR_?ZY&[<
0dK>HJA+2X?[/60-O@;1A>,<Y@0aE+049-8]X<5g\XN@HSKZO;,_(MG4Y]2;VeT[
NB+1BJ;B:O#8&:C&G:+E+U,D5/D5I0ZfBS[KGX7cYGdfd[KYLF8GV@B6d4=.a;2)
dIEV37WR_;/O8V.XffOS8(RFXB754FQ[,N<,F>,3,E\#b749D52FVf&C<XJDNEag
)^Z<8;5Cd^A-MO^,dC:BWcH?\/Rg?K50F.,R;d7++IE3+S2AeL0L)b?6?EfHW.@I
W+a4//WH-3Q2ARMCZ;G_aN@734O?KXE>2QgPRgA8W1L9M#R[T<6ZH78C]+7D^5QI
XKLaK7dJ_4C@_FV3,)dFB[S0QZVV);ecN0A<b;<QS#I2QA?R)@2SFO&0K1f&L#GC
)D=7^>Oagg/=DF(2;]OQAX5a<&GG3FCHPfM^<6B00JE5cGA=f1>ed/f6[-YP/7Z/
F1Xdd63AU/1KC/T>-)F28#@dd<]ERPca4_KK^1Nd3ML2OVUW7I4L>ID;]+K-IW),
+\Je,VXM0BBLb^CU6\/)5^E?K6/CWNY82B\Ja_>cP_T5ID_Ff.CRY@Q(I.DY9g.L
>YBbYZ.FIdR^.eE<KG[__Uc+>A+)f/3MK>eB(f(1QZAPKC0g3;&](2)1>^?N;2BC
0[H+_9Tf:M@E4bNe8J4NZ(29R-<1W07KFT)@:U&_.F/b52AKWDDa,XW(DO9AaFD?
@EIL-V?^)KKeL\9,4&O;@9-,O9P5X2\EOP15X>MO\b/.:YO?RTH&gZ#1SVX\cT3Z
eQ>?OVKM^cB=_b/J+[Maa?]+c\b\L)YLe\dNM7_[_A#U?;g-U;b+C4L90NCX8-QC
G,H(7.BSLade,+P8_2-?K4MFP-_]TQ;SF&)c/YR<d+5P4+0@XH]R3KPd8T2c/3Q[
F+&+gBeQ.f:97[KL<Y;H()@d;,4Z(e:d+U36b+gV;d@(/-CGN?E70MQ46eaD;d],
,CVQ5409gS)6GJ6/<3VdSb5Cf<MIRaJ-_.LAQDZf^];Q8YI+)/3&64QVVN1/5=Nd
RSV<3E5@VG/ZSQN<7U;a0G.+5>g/[#AMQ,YY;4?]Y/TbYFC/V98CD2]RQ:#<SJFQ
[H8^4-e-c2HO4gUG=7Q?6e/>V\XWZ&HAf],Z66G[C9(;16F0fG(f&b2JF80PF,4=
2.9deY1&Bg7?Lc<OF;U2g7P?#B2TJ?DQb?R-cd3fCbR2IYASNWS5VNID4(;;W&-@
d0#N6eFY6^T#^ZBDK>Q@)N/YR.^C.S]&.#DCA/Y>ZX(;QdNC,f2cMNd-Yf5fO-,/
:#a-2S/V5R<f,M0)P,GMH/.b[_/3<6)CU)0K92CVHS?eAOX2[:f8@>FK7dB/23UM
57Wg+O5@7^&V;W:1Uf7EZFe-A4cA[g-cHcJGR8E]M8_USXgS<2O7,-Va_Z+>N?_4
dS/UL-S38G+]fN,/c>f\YS;7-+Zeg8.Ga94@42d,OINA0?_Y&d@W4N]_NBJ=U.QL
L7&4:e(P+A23c\DIPMY-I7CT4Ddcg]I/bC--XD;3)@C2Y63<;TYT-FQ<J(>d:1c&
)fSHMIZEAU17SCX_U9R>\\FU^,]L,(RGWNB\EYYI)SGO>7Y@ZQK1J-5F@_U7d#8O
2[Y.)YJ3<f<Y9:cB4VR/^F^L)fd)=C.NA+(Z([bET.#\XG.#_^Q-bQDbWU[S2I<H
2AH8R_.&VgX;:=AL-bZ22NdSAQQM;I62?E?HGC<eAY^)_;c/#NE[&egg6M7XI8F/
T]LMH\5X&,b2Of,de52RK_Ec&ZT_eP:5HNM?&LJL7D(8DC8A?c4Hb4@=(a7Q=IIV
;596&SP,QI#:?;c5B.SL8Ue-DTb8)36Z_:]F6+P=g<#1S0;1f6XXR,G-?,_LT+;;
cF[9&JA/:0PL00K#+?P/CNWSW^HKE<<QP[Q[UAA?S@AZKgJRCLeaa).U7/9>^S/I
,8(&I1W\XA\Nf59G^3YDd<f=F9-Q+ZB,4Rg,)HWa]-gb+7E]If^Z,RQQV3,F,1cD
dgGbLgf7939f]ASJMF5Yb<g<)&1I,5a?)7TJ:D^(C5Y)RG,DcC_dP9dHU5M7df:V
F9,AbQ+??gW1Ta<WZSfO[^J@cC2(f@@/&cZ2PZ&?C#M\M#_a7f56#;ae81-W,f]7
0.MK;EOCN@.=#CC8#O/NLK5QYT-QMCWY6beJ^S9f_EO#B3)#+9_@:=GVY8#\[C>0
WJOD6.TI3)AKR5/5d#(0PgG>7:\N.:Sdd#,_]S:@I)Dg[8<0NJ/TUMM^GG.2;T1<
\^1aY88BU,UG;<NRgJ:^#K3)2SAX,]_b31=9;&QdG7AbeO0O4IQMW\);YG.76OAP
T<TFgU0->;P8GM#O(fO3L:?b04QMS\0-78+2a1R&+TM;M&8Xf2NAe1OL#CbYEg^G
/IQ-9AL(7B3C6TO6KPCW4]1O_J4OZ-JgLWNGXNL:#AIF9&2LQ/&d()B16VQ&>=)4
JOSGEMLI+NGcLSc(4AcL+)F[M3SOA>1-MW4CYL1QbQaa6f(edH8#U29H9#.K&:=8
BIc[JK[gdT&@81#KX7&)M0S;[b;ZAb]F.Q@DPD7X[&Sd9.bUVEN:Z1R)IX[f8F4@
4eOFT;+dX1]/OKgW6]^[aca>=/[EgT/62,T&cPGLg?5K?4SZRBdH(2AUT;5B3)?,
Y+Wd6UdH-BGgL4HSF9e]d)GN\abU@c)Z9>Q5Q<9CT?866+HR/N&G[dCFaV=38Q3,
MT;Cc1=MFNC#])3-2@\d?#c>TUL&5-B[dV1\T+cTb23dOY9cEF@D9b0586Y&=J6@
\D<NYTP,A;/CM)RG>J#5BJ(UBUNfWKSW28[[T>AJ<eB4a30U)RQR>O=b=?2b9NS&
O8>f<@C\A&Td0#LaG8@^[ZP,\#R12GDRV.J9Xaf^J2cAdG8;J;1K,P#2ZMFL);8V
0a(\=N>#619NBXR?Ga^<7JV:cBC1KJ<=,8?^6[4gL[R3V#([\<M#gU&e[XBP#.8N
]QS.IK/7WE?97d:a/&eP428<OTf^A.#^&W>A5PRXFMI#4J+d&3SNHQM@L&,g3QLM
D<O#1C44Z<:I1((?LDRc=-b/6_I6ZXK?8FYEEHY(1+&I0<X\L;;c6AJ^=-B7&,Y#
Sf(3e\AEf@4>GSM8e-04FJN?YBN#6)Q6[;#/AgU7b.#95]O,HPM3]5#Z#(_+D(S7
A>Q@gbK@JBI?R-&?//E7@V,aW&R88TJcKHTcHJD=cZ8:6f=JNgdWc(.HCXR0(Y=A
DNN3]e,.\4fRcRSHH:&8.A4,:6PO^_E]JR^XG];(FHBZ&A,f)89<d8Pcf<b^7G[c
E-X-S;MS)CUKE&[;SfM?00Q<9EK^:RMF#MDYH&d7bP+H+J.>)MJ\+6MP[b>A[Cb8
M7OI;<?ZKN-BAY0IXZ4@&1DdB=4<5UE0e&,+Y@a(?N20#1Y0@3@M2/O\GYZW3D\e
/_OBd:33bLQ:J>1#N,]NW7T@75ON5LGb1DaH.1WN:IZZL.gM+#/4E]JBZJRL+a(e
E8)LXT95IS6411?g4/@(JEdJ7/CP7c3JGP(gC:>==3W;QdgW/DMRBDAfKNIfHIOU
Uc7EYB(VCB/VWKU2NYNS-IZCI7=fQ0N)X^/OBEXP)XdK,M#=]G=g]FHV#5d2IT0@
&YL:f5KH6U#Z7<94Dg0L::c2[1T;6bb(fE[gf87[U3Ib_d@3A:4f[#+L]13=aQ^,
CgBfKM],B?&=TAZD2OCYY<0ac<fY2/aASb6QS?A)5Z+]d8MDZ0@E6&SKbT?d;7Y6
b38a:_eSZ\L9Q\aNM<gU50YdeP2HGA^Sge@A)bNPNNV:P\?+V=OY.,R.^CN(c]J=
BO,[/#J.)IK_-X>eW)1?@/<OKFKB]ORFPSQ;RI?L6V9g>QU2E[7O[<M_?EHIbCCL
7T8(UPK0Y.;M2e79SW/EPST,g;]H+MG_?K33^:fa1f<XN5455SdTUN\UScABc-a5
eG)0?&D.5N?SbY7V?UN-AgK#@=95-NHB>c]:5)N\[3,E(4Z0VZ,FA.K>e.T[?U-C
62BR,dWdI#(MRT8JHC<)GLQ>[)DP7@_SU3GS,MT/]AXc)VYGC4HGFXG\aMMe(\dB
6B72EAV3d)H?=-O[&0R)R=C^aS,M)/#S51O=7-Q9ONOP7D-:OKXY@,dFL0B&2fRC
/cF,K\^=>gS(,1TH-+KaBFf3_a4cgYL3I&;,ONUYW_.bDA]6d:BE^1K7-/4Q?WP@
20X^WAJO\9NfZT0)I4.]KX-31bHUHeAfR2=<H)0W]-M@\R4cUA24\YD=g+e=TgMG
.-eS8AR\V>5cM(O=gd_H^(d&>_73V0gHJCQ)U]P?RbS?]9S&QOL+fZTUbFDUA:MJ
1\edcY4@I85^2JeRBV5UcG=(HCE_TF>\9VV&QK>gE3X<.S#R]RAK,Z9Ve,9=C:JT
T/G+CI^g[4gKGM4]B8>A)KV_bP2DPe/](TG(fW5FY-;f/^03c=fdL=58\)Fe_PbP
8b;>,(,OP71N]PB.M8:gG7X;W-VXGe<^c-;?7ROgf46.1+/\M<_)]6H:eSF&e8]#
UL4SYN?KHE/7:HV@0cNZB/\:&P6cUY\F6=XS@fL3egN4FJJ\eXHU2e-Y&E=NVUO&
]WfZ,IXg-;KTSe5)WcG/HP^]+;OCGbWLD/I#S:c]&WKT<dWVO^<_8CS<D/V,=FOf
ZCKA8&)L>90\GfB&FQ]<d2N.D#b9JY5b:^,^ce=FJ#SJ3b)[W/ZU0OaOKB](GNXO
@QF\;&Sg;]YGIVXUJdP[^VD1-T?.TK=:BPW]:Vf/XHEAC31bO3H@HZIDV+/-57L@
-1,]@S3M5_e/,)+61^@2^H0aFUIe34A+DT7VTLb&5Rb3VD0]d05K<Oa6M;PAd7Kb
UOfe7=9TRI=ae_<N?8U?bF35b<X3E:egaBdPWc8[.G6&S:1Q+GSV]T4eAHa7eFEb
U=Z-1JE4_2Ubg55\YE+#F80d.SQ3MR)IY0\WC^eG9C2Vcbg7XR]Y++W5PG7.2_:9
4W>:(LNMTV^169VUd5\T,-cCMTIc90[BRWS<2&:?aI#;VJB&d_=.]\;=PAbM6_86
(T+MER67W2dX(F&gPD[__Z\<KFSJY.EJAS8S/E5)G.?Q@9B[.8^;+J4efJR/G\C;
QUaN5=?.KGa\1).&DEMeT/8\)33<9A:XBTM]P7CBKEGZ--SCBaAWKK&)cf2-f+AS
I+/LCN^JIfQ(?6F:SEC]T[,T_MUSX8P4aP?DMSYLfVcND]_IFe=_Y@K<+gH(9EKV
ELQ?HXa8fIO0>M@82YV;9:02?ZRI5D(R.C67GY-=-c;I1?2H0_<7UY(5PNK]<TeW
I27\IU;(GaEE@-&J20aEdgc#0^CITB_e6;BH&,5[I,CH^B>1YZ=9#3NbR7L9;C)P
2cL_O1Z;GF]ZdE<Z9)ZT0&&.NOd,9<M6N0#_EMcAa5D+>E#O?Q7aJc=_^ga&Y(M4
D&TU:2EI5M#6-NS[?_0&(ag],)cd(GE1SXN&]JgT)b7(?N2EPH6e+<T@fH2C8GOK
@Z-:;G(Fg&ZI2NV]bL>D@,^-K0/Db)Be6D(Q:E2HaLC]RgS(eTAMH1OOC2],S/#R
1O\5a61H:Z&eM]EK9dA;_ZU[,XV?)QSLF19M3fb>56A=U>B=SU1\9HT;eYC<XY9e
+9EM<7e=ZQ_RI4^PS>EIHNgcR2ZB@6B4=KOe#9cKA(bUcY2b&,8DGeVQMB&X@-D-
a5ELR]c/8++YZeL,T3F+)Sg97EL<;aQ8](>S20fbX@;e@3KPEQOX2@&E.2aN>[(b
H-+O/^#>)I^A8:K:5X=L^CHAW)bIB6N>H@@JOcC+(8gOSO-5YUe/ge3eXa;b,QZ_
EN/V2J@)e4Q:I1WG[fL[O^EHS/f=G6F786_=e&S0RAWf-RbCf80c6OV57aGN:.YN
NTJ&FFPC3I[._9-[LeK]C.IM:bU#ZJ[R/?MYZ^+eEaEAO,#=#C]\&78.,]K?SDd/
d:30VC/?)AR&g97U,-&<JZ[M&342Rg8:Ad>b8MR-AXf2<IN_MPEZIKENDR^cc2P9
Y##L(O)J0^GCB\<FOZ]90@G94Df^(S<E;>-d7CM2,+IcFc+]3/DLA47Vg,H)>Nd-
H4.;1ETIdb;//?cLHYHC^0688D:&&BFR^-7gPfY1fK(Y<0f#ETFN5/W<7&FNfF>U
IIW_3:aeL5L.D&gBb.Yg75(59C5MI^B..^:Y+IEaE2dNbLSS;U;9D9.6JeVG)]fe
X,9IA(g9U:g/_I)<04/NX4@&_:M9;DIOJb819D0IJcYZSbbE2RC]H\JRC_I+,R@(
(b;@Y?=MQZ;c.JE\2GfF.\1[N(BO[NR:W.(3HVg\<g)D\I>[,]DC3<ac1N-A3M2=
^E/NM&=<;/7:3D7KgTaCR:NSb?^CF=EU-_J<Mc_<\-O@#[Y^33]12VdgaJH+@Xd\
T+NPRY,+_@:@Ud.WEYG>5M?R65)XT2Ke\XJI\75&-#HZBbW2Q-9KE&V<OBO+_f60
bARKJ^2\3?+?=e8QE?Sb4XcgX?cH=P=bb2AELN@JM33E<N;@4GNHX^>:17PBOE07
,NH<1&UEX6=\A)0MHOe7>T3F&:f-fE0G=U^18:C5AE/=#@SC4;NBcP]LVg@Z<K]Y
OVXWMa95,^=?QPLQ#XeBL@/^J_;GZNOC<17YR8BKO18^]X.\#J2PJGfO&#=4^WM8
8QEE^RcF#c]Q?R@Tg7S=LEeTEHQ5V5V],_(X3[30)UL;F7-E^HY2OfRLL+)Z@cQ:
W9J<Y9\4/aYVYLOL1Qe[APS[S-R<>Y-@geDVWM6J2M9CGO^T^O),]DNPBIcJ,gWC
ZH+(NZB#e0a0)TfG^_Va1^4+Z\gOe4UDO6-;dGeS,_/SI2JbA;[=:#&GF8Z\)Q&N
:;GJDCVYT66ZD+F2bbc7EIXa,be(-;9g(MOURA<WC/33H,YG_Y1348Q24>\bV_UX
=R+G&^A/cEA3\T@d#745@;c5S6=^+=6B_-GFFg=PR/BeO^dg@R7>OS=:X7V_^DRE
g1[&#ZHDeT=)P>@(BaXCQUS;Y#e0LH39V0J@=f:#)M[YD)O9K:,(N;bJDQ,_YX)3
b[\9HTAOZ\&FJAD=?/601&Q_QR9:^bP@,_/=E5EK1QLWcGdM5ORTTe]Q[5K5Ne-<
_-()\#fgcL0[K-PCbHVD>Z.LN1Ld?)IJY?L_f\gGZfPKV];>HZ(cK)>-aeG]:[,c
\fQZSf?54D?D46EV@S/aU8EgNQ\L9DXfL@aMJEdFe,B;Qb+1P:(14KCHTF+3U>/W
26_YBQO:b5RJ7\cCg_:S1SO+35PUcb:L6@9OXP3>IS8G[b.,NK]\F&[@X3L2^PLO
[Q:@#VXM1#/38/#8=HWY][D.=B;O[4WV.H16cDKfWW[4J-B].PB@72)7Wg&]/EHR
LPM7Q-Ub^e#NQF6NfN(<3_=K?^72F>VS8^I[[@>/3-Q6F\;9@NeQJ7DD98daE>Q(
KA6@M]RRQIGW,-,[BUSUR?+02U&O\_.aAET^Pg\e)NUSSN4DYK@&+;7I0V<R#aGJ
b9O,J1ECI=2gM^[M4]2YLKQ@1)XG;8Q@dH2XJ8FJ0c<TPBaP((4R#PQI.G[RgN=2
E,,g_3[1&cDKQMRX^:APG5)4e6)I\_?I//cfGFZ?D+[=\Bb&Z8?8eX^>L0CYe6:.
.\]6M?B<e)GWSV8B\D&B)8Bab+2&8:0CR:Uf&R,)](]9(@X@\R6bC;^N;IcEDE=,
d[Q2,96)Y:U1M,ZJE7UTQb?gUL2)bF>[WMKPAeM+BWR4=I4R)3<;FR\<49Y?c_KI
ZEgHQD+;SMS-K>65CP,e^CK\bMM3C9Z=R9/X/4-/C>PN-?:=M0_]QMdB\3VHN(>X
fDS+AeB=<)V2\,])0&W@+F7F.7HJ57V+6e#(EMXg3R1e[P4M65THeLRFW=EZ?[A_
YSI:[661,_BUeW:,KL@T?2MH+PI\H,Y3BUZ[-gU(T9[#B&\<bO2:?]3Sb\KS-<2D
MH7=d,+0,ZTKJZ/RQF;#D1:?]04(Nc4LHN<a8T-,6?d)dc0L7[8IJ:^K@2.Y21O(
;,0Af>L.2N/UaD<OKSM+[<G/L]TSG\Q_KXJ,4S9_9-M>ESR-,UgD>C[B(OX<9RA&
U9dZH51[LJ601)N-9TR-G#<a#;3AQE&8UHLcS(,215;+OEdaaNTN?0BDF?TOCHRf
>Q0E+C8#Dc?R6@WNL^#LHOJC,3a+90DCNb6O4@3)7,6,&a(7NA[11N=KP5<](4/c
XI2M(1fO44[.Sc0GSGXUXA)2(e)Vf_,+TG=I[8+\5POfCQP[X\H/1[9XJ\DV81<2
?ZB)Oc)A.VfPBT6cFZG_OO29\L\9&]#[<QAI,N,(@9?b[Ob[@/2OFO;ERA;,E+JX
/9aab0RfXNO/VaA/+K,^[e74NCB?FHe5([Q>+RdBP.1M\5LEQe]T?0[fM/7=T(G7
_=X#2IINM>O8>dI(&IIDHH8Y+JEQCO_=FQ#8/GI]3BHY.J[YY8WeC2eNYW/C];+_
N:-)#=6WOcTIOR&_-]OE_/0XAOHU3V0A[A_8T245Z=K/RP^.BbBZ]S37E89^d_[_
,_[Pg/9()M\5W8O60=R.T.<2G([=)W<P2YW@9E2<.e?9,4B90ff;_BXJG^F(E#d^
6_X9V=N,G1N)GK4]]cNZ(BeS,D6_\KB,PJHD?&S0a&dd[2])f5BAAW-7<ZS2:O@#
D<0H_CG0+:Bd3^\KD[CQ+&RTcZFb(,ELP]Y&LcQ5N0(^XZdgYB:aB8GGX&G_=X>,
\;VRN0YTfFfMO31IT+VS=.Z5?dMbCY@:B6eGD\X0eU2ZA?-XYG<#(3;.4@JUfV(:
eU[[UD7J\+2CG9=Gf4/<?>TcDWL,B&)81.2D>gCd3KU(_L@Q6W@66M8/#>Pg8Q@T
O7/KNU>AJ.DBGF>\X_eJ3^A(BE+Jf6#([QV1S5LBH6J)I7Xa/V)5b,G#+56OIO&G
ZCO]]SNC]<6cY185K)TIU8(HAd1.YM/X:O0\g-QG_=f8V7PFcIU.SE2R#c@I&8-6
WX7fE]:XIe>T9:GL#I>HUK_/=/FbWN_;SI-+Y[8M_bD(SFgI^_:dV=:J&&,#2a8Z
+gG^eB>B@)>/a;3@FbDC5=3VJ3,)cGWgT+;&0I=\WB;3fY+T](XT[K;K?)6:e8_;
]-,W/JT(9E)@0W+T#KgI#BBe6QPTG/@Oc\@569@)MFLK[.\#46M:[UX)>9?[K-E\
d/H<>W5d#d4,B>VY-XRS.<]aA_E@W@F8K^LLJd9N0RK:gE\b+f7YGO6\NJ655A:W
^;U96(Ng:9YdX/9&_Rbf<-=F1X\SJXYSM5F:2b:^Y3:/-#WKgDT_I<^T#;UMDKJL
NE4,O\0WMPUROHb-4E_W>2WC(R81HH,4/2QQe_ZD]Y;>V;@;a^]O8+eb6-Q1PXDZ
ZZNdM=DB98W3S:afO=(Y1)O5F0PEG>8FZ?(GA\A3>+G<fO&Z<K:>4SWQSF3UYR:e
W62\8R=(B]B:,VfI1^^2JeQAYeL<Oe<Of)\>[A0X@eIXTXHA_AF2);E1[OIf;;+M
Y1V4@:ZQMELTDOT.aT/^_6((f14TMTf/JV,X7dY\W?H@2eO914+5JAAJg35LRSEF
N\;^eKD1HB,0ZG=Web6e^-@^DVYJR;YTC_<QEEHCX#gLZg)M\URLZZ#+1N[&be)F
W)[/V;):@&6cJ^F;ge)DbZ<OPa<]2Jb?+&\B839_L2_K,#QSF:f+>ff,67PB<HZL
P+[<KVScN42Q2WVTS\A;Zc+NH#CF:^.6_c6NI:381E7=GQ3=;>&83BJQ?MVZGO+(
cS+eZN_4,+0KcI,;Q9eZEIg0@1\>Y_1gEPZ?D\,a1CXE<E235:DL<;#,@@;Y@5<,
A=fc^\C9VPQ](,Ib90@BaJUb-\UY\Z>+1gDa[]eReI/+6,A6Og)&aA@eRJT]Wg[f
Q,UXE.2g;0E^,089SIb@FScZT7Hg.g49^F\g?PS[=d8a;UNPTV1X7CSN98f<aU5e
M5+),9dQK<<5,[;7_F2U7,Y-U5[>:aHX<F\\H1Yd_;)P((6M7.EM(LFR.b@@]GaI
)Nb^J:gF.QXWV:[=:ZL)^e(>HQLWYUIJ-0UC(QY,Q3-39]Y8C1I+\?Ccd2]&H/NH
b/+-M69]g)J>d./bCR8PZeRN54X;QY2SDF?O^(ScZdHUgDMTSKQb5;a9MQQU.\cX
)<]LN))Be;c6919=(A+EW=MaYYYLH+e[De?Y[ZW_UYJQP<N;[SCWIE<GD]IN8?[M
gO1J[O@B^0GY62&.?D#_;&4(dbI>L)HK6S]^+6<]F@UO#PZFPXH(Fb3>#ZC];[\L
Fc\d1\G]LaSZb)L(UXa>A3[B,H0TVBJ&RKH97Nc>#<Y_?a<^#aRX0KP#]XVD+[9Q
dDd7:A+ZN9CZ56/b9FBN,VG-O@a_7,CX9:cOF?T[-61+Y.8c0_>PdT^PU6_Ca-5.
+5/=)),&g@0N_#]M);f:,7[(RTd,8Q]L6ZX<H&_U0;#c6L2][.0E,JQ?d1@SX9B7
fF=\f>MeJR>]A:PSgaW>FU@BI7&b#:<C?UA)0HW=@eJB(P_AQH4AHbRK]5OIRY.E
G6_-@<WNcN/?dZ,=^B/7[EWK:+8cZ^?V@NO@GIfR,<YYNV\FM+^H#fbI11P.,08c
cA\gVf=):bO\fRb.X7c8]Sf45B4PQ+d5N45I8(6d]7X+VTLOHVXJ?YOaFABDgB[=
bg)HZ9K:3c?Ff2Ye\UbV:S;+A;7\,+(FgRd]P4\]R/F^W;9)@#(ET#d,39INM9@\
dA;R\XZ\<ILE)O)Pg>1(JBS^7EEW#+d&gT9<&WOJaab)VCBFd=5IB&CecS;8<S&Q
^.e)0(@/?DYJT:cOBVP:.7PHSPa#.?gTR.#D\gG\c,PWK&7[,#E4D08Ze+\=&C3:
D+JfXe#&6CV6a;fWE7XDOR[?QgD\XX6EMfgW85>>N44&F+G^R/SgEg@+NW@D(-0@
.L7T6J2-g03=GfQ_Z5DL7ef59K4?I<Je]UOb8\FYBPMLO+e9?L,>^C7U<-:U9XE[
T+Zg<EM.TVB62g-A)<D3V4L2,Ue?++\W/04[8=NX^a4gP#XEB\BZ\Q^+DOHcbCQC
^F,7:LLF2VEf8-)YG.g715Qd+63^QX&b.C6_L\dY+@[03e.g^UOEG#d(#;e<[H7<
@5;JX)dPgKV4V0Z:#V8-:;[0]RJ&,2LS<R@[V(;.S9f;#B#.<W3ED63X-LX-?_CN
QC>L9/?186<C=]X_NZ>SH\eR<32:YPK[E.>1W[)XZRE/LE;AT<b@T<81^2.#+63&
-]EN?C(SQ:N:2409#RT0UdVV3.gH,bCRAIC6bJNV4>VT:R@:<RbLJQL3;@;[\.=-
cQb9GA2=P29&c3X\6=f[e_M]d\cb@g?B:g)K;3SWZ,DK6SNIe#-37f#&)a8).(=9
e7X]3DYT.KKASBI+)(#O3ePRKdf1H268,0.LO_R&MQ>NbWSJN2)];>O&\a7WI^??
8DM:a_:T/:^V?L#VCJY\Y3ZSQGOG3M:\)=#HP1@[HW:RgPT3IDQ0@&(c#D07[V\5
_g;=aQAMQc5TgHBdT\^0,TXDJ/BaT0WP(df3,S<[_WO^>cW-.c)(01=f7X,d3(5H
R(:DbXH&-_Q,ID583L?X;/&W9gQ^L#M#(B3.0DTYOX?-CCd6-Z6Z-d6:+gH83Cf(
Q#OH(9Wa>W#HBe&GLS3aa^_,[2LO\#dMR&/JMG(E7P?K6V+MOced)HD/[9Y&1+FM
P[cJ=6[^FN6ROCQO]DJW54^H2L0S-e>c_B8ZE642?Gc)2+8LXQ;N,ZJ+3f,V<8_;
J2-@e,K^HSC;2B6bgf].O-(I3eTWK3f6;ONBcV-BB-9S3g2)[-+UEIZJcNT-1e:a
Z,\_04eV7G4f@EZFK>.<<e+Kg8:1d]8KE6YRV48].b:L[O)(d[>]SXY:1PNZ#Z:S
K7Tc8E?[JPC(/C:7U-;\>fI:5QYLd?(eFOJ:CT1:0@#Zg+@:>ZO0ZY#.:Ff@Y:M-
f7=Q.2Kfdb(3#2e(Ya#I>8g<4Zb5S45:X_DVfLA,[:U6c>,:=FEK]_^YN1Z2-;T:
<bA6^-U7R)V=DX+KL<H)cG+g1HR?T0+=ZL+A<[+)KbIA3-fK_=dG=:g37E>H4T>e
/6\b#Z)WO_<]?_YfXXNSg_HED-\b@X<?_1G6Db\U@E<30MI-3C6R_9gRD-0WcP@0
ZJ@N?]:G38gH1L^R^dNR19K^+\ILEC0A^e^-G^FZ,X0[T-YO&1LG<,+Q,3X_LT1,
K&&WS]I-E2P\,.00RKR^90PdL,@g9JV(,3M5DZKc^,9aO:?=I,,(>&eKDP;6=U:U
Z,F<?:D:W:9E3U_.REcLDLNGYc85P]X/1g.64XeAKF)aN1KaS#(2(R70e_Ze<8Z0
QE)YEY4#c7E\V24Y-QQNCK;PL@f4UJ3>2^/,g4+f5E&[Tc\DU0QTD]RH>=c5PPD7
4[O<d<S#cVbaa=6RC^6XC1X.aR<+U-Ic.d-KB4LYC=I<#c\XaWM9)ad@(+eD^\KZ
cM+Ne[AOcg(Fg7]KQdccIXfA&LWR0+3H4[dOM?JOF170Ba:aKC[HDX[(aG4F.@G=
#>(BK)=&QA[OH24+C??d:QR\MC&-dG,PdZZ2#e[cA<A)bVe_CbE.IIB71(M#YHI=
@7aO0KCHZEX3O8cMZ71M@T/3YK9@)8EacKWOWK?Pg&f.2ea,93S.N0-5GK3gT>8V
&P4\_IV(18Q;3.5cF?0Z)X0DMb<OSfd(H_8Z0&Dd<GA?=O(,/=C[\YXQ>A\3JU;[
J?=UP\BSIMRY(?Mc]-1)R@&Sg9#5<MaLN,;MW_KD9(MCfT.LTK^[K]H\@WXd#_&(
E_LTM_YCDb@K^<[\CT^BZ=#H]>,/(?IRQVE\a)Z<3N.(gb,Z=d5X1Dc?[>f7]E]B
d@DNc2J6#PfSV6?YC#VBK^df98f)<X6YO[W-.SSATLT^+)T&3\GNNUMFX\C7YB=D
+Z0_JP\&T2a2gUU;MSDXSYK#+V<cRQG;3>GF2C3D?,7&59&NdgOF^BB=)\;1fE;C
4E/I)3-+&/Zd+P^Q04-8X9Ye+7475J:b^O<01G@4g[:(e._-7gU]?NK,NG-2N?:f
09=LC;3Lc.dBD+26WFJfMIOY@)Vf?FD=Hb#3<<AOePYX,.:G&ZW6^N[KZ[dD@d1\
.8)M7@UedSU(7R0;09:H\DVW16MCD>\6d161US8E7.bK8^Z6N<2^KX@1d6L&X?Y]
_8/7)=+\=4McF-Y?O?ZAM<DYeg5IZWX85-S.JM[(/=&gU+e,W1a>R\6/&(@bS1G1
?Nd.Id9d7IaI^VY&>Ma>;K&Vd.M>9@<gc1H3/WE9-,3BP\:K/K1[66g_PINCBULZ
2@WTFfEXN@S-RMMVLc#L\[+#ZP<bWEdGb7/=4DC3])U-6.N(N9_:,=QV1W99.LO3
6dab-c8cM(U?3@;=7<\&8FR1>H&OS.;D4AV[gZ]OAL6PSQIeHc&[<[[7<6]=b[Aa
MFBUSb&cKI:]C[O/<TTYCN-/AUVBUQ3?5]K3>H)[^(PG6S0cVaZZK6G[gb(&\7OO
)XA9+D6CQ>AeM-8dV)@L<NMWefF9]X:R_OA@:fJL7d78M[WKORV\cH_WQ(FR6LZd
/&,@:BKD\[@,>J:/-_Q)3^<6[0^S,FdHC/?7>(ZADIH:UE3A0gAL3AZP_F^8R8P8
<&,P5WC3ZRac>QOL_7]#BMZ?UeU2IYFC9@D37PT>FR#ab]J#=PWS@?2C64f26@[f
^dQCQR[8G.-Kg_Z@PCd/GQ^:W@a6dGF,D5A(.EJebS^LNaUU\).P8#>f[B(?W@3@
71UQVf06KT=M;:F/Z2Se?AU@QF-E/3V.Y],[-K#X/:A8@g<WQ28?-)=LZcU_+M/N
#AgPYScY([)MXIcVI\5I@]HFM_,A1+(Z/b?<fH)cI/(^T5^RKD:9E6@OUUf]3[dG
A:?3ZG-]GJPC.a<?3[MSNYabMJ5@KKAQO<f)-H#^LdCX9@@P?WHI[M\B\P.5(F-^
(CV^YBBD<C]\M-Y[(-OFebCOML&KY2<EJ;:;NU85C>+<^TaWeKe)F1c2Y3RcY[\X
K]Z&W1JVe2AX\2KR8QB:9C\<MMDKc9eZOF4/SeF8K4g#3(ReO]<CNJIJ>)HO<QYG
]B0;SJV@7&MTJN?HT>?CZCWUZ-\-2A+>?.=)dG9+Z4>2aP-RNG)M#)DPdF@<Yb=N
SRFT&AYQZM.B/QEUE65=NG4ZA_gIee\5Y=MTU),9b?YYS65D;R-M]5IEO>])L=H8
Y:_)]#D&g)F,^;cP&_E6VU7.Q^WL=0KI>cXF^@I3=F-e4gf?+57SC;30.Q0DX@^f
3T\,<E97CTE/(^J+:H9/a7+<E<Hf[]9W+UHcgbQFUNTf&DC/QR<?]?AZ>L+@H3=.
ZCYaXDAeU1+C(W21S=MBaJA[INN=NPMV9MQG]L>H31ZHfH>N6\\25NeR29c+Hg]T
cdB:F-E31ffEE3(]D<3>\d-/JH:c_S/)-O4JO1(FWCJA<XdafA?TC5@V[(W[14O>
g[d]9GDU#F4JP4eWCS7;;.0ZIQ/WdV^QH3?7G?>NAI9_F=3X@LC3f(FU)-+c^DB;
bcTf]fW:(Q?IL2;c?QMM2U6_]#^Y6&4G25Y4_H+HB>YB:NE^VKF.K9b;+I_&QHUL
\:BX1PgT2Cd;AF28GI8gdK/J3;RW(bHT:QJ;9X6PQZ07WFaRS]e9TSWfDJ.ZSWgH
7g+c([0JQE/X2+Nb&F0aB^R#)(52;CV2_0e+E@Eb:;&C.X8b(\5<4O&IBIC;J()(
M0?#PYHSbAAOb2P^(L[<(gHXZK^D=6^NDKD=#<\PLPP#eBQe=/.U[:^\c_)FgTXS
:I<H5H?\?_9bQW<?<B#6<@U0PIPCaf566/GA+:B;:0?L#a3AeB#ZRcKET=T08++d
K@Tg)V:K7TL[<(-IPJ>^fB5Y)-eRU<-5A/&b?Ma9b<fbH@;G.>Q;/,3\1/eO?CdN
/S?Pa=U4be35[Q1Ob1V1IC=_-#3#]:<-8+Q?&O4JUe4AGc72@=:d?;^X7VQ@G5-c
?VdCE_V<[/&B@.dLJ;gX;QC&#X[KcVJ\cJ]UMYILQQW>c/AdFY_J^3cH5g;C-3ZO
Of[ZaROb(W1]^PfT9[d/@[]05GXeMVa>>V@c+dQ:.cVf7MAH\3NMAcGB3E=:BG,\
+5JIfL+TWSY1\Vg]B,TW(#Iba^X6>J][)?>?[ZAGK8cUT:=4X#6NR><)a];WK,SU
#?-cdX/=HZOT#PSP)fT7F.BOffA8D[-/f6R^>Yg8@Z(A[fa<E][=G>g=NQS4-X^1
-G><T+TOSdV?CGY<4Kc+HZEH.CcSdePRfG>/0-Z.+VU27>d9W+/-/WWHZC96XH7/
?6d_:20G=PBD6R<)_T]GSOWA]_8J=\b20@)@+E<]^<I-9Z5Ydfa#K55WTUfQ^+AY
UEJ)>72M3=\9:Je3dZ<5d559Ha,BI\+Z8eTR2Z=_NEG^L)cN0V<&.Yce5BDT&Y@8
,_WEWb?Z-bDSH?V^<8,bUXaRIGB,:_R6+X1#BLbX/^#dI<0.4eFeCI=GHXQ9>K#7
@c+XVdT_aRUcGSI)g:.>@1WNb-1(LKF;&f>>gX\PXJZG9/N<9SOW(2W22MHGfg)H
W8WU_13Y/(Def=TW]?8.KH42PZ096:;4:c@?):VaD6T^W9gZM?2N&9.3(QMVBR.V
O+eHF414(88RIUF0H=YA,GQ2F]/=:^.+edCB8I=ZK4+0FgZ5WPfDU780I?V^<8FZ
N6RGf9KB6/^8aX5OD@RG?U.+/PBD=?DP<5FZ)5/1=NJFSFVS3<H,:f05N1M8/F=Y
\f5E7^DUG_I6dE(.ZY-[9_02\^7Q9dRdP<YP#@e[WOg6WTVNNF_a18@:,)6Tb@.;
9)QZX@?QVBUG2VN)S5ZgZUDYXAL<M[)d9__>ZRXHQVX5bX]\1L;aSQ5ADEVV7?>K
@7ZA.a[:a4_9Qe-@+>\0^_FUTGMK+LS5:46?X2/.IFFWR]XR1A)P.3I7aU7[2[U]
>2;M/f+1DeN:];28:SI0IXAA_>--5)R(#4>P^\IYAFXM&=H@1MN,#Z9>T9Ga_NJ,
O\;/ZHBXeK4VUab4)Nad(Y>P/08a,WKCgSb3J.)5FR\Z@8e?7X03bL=9WO#1KMN.
1><9GN1O-/CS?K\CVF.@4T4NRGgP,f8;L5+6>V(12a&A<B^E/O:.,9<=I3I_YaTV
FQd4SCO5)Vf]5?b(6fM:;W;JUV0E[:67EHHaBPAdYb#NEeOO4J-5KZT6GYE^;^Vc
E3\)fUF5<5X/W<?0d&WE\fT<e=5^\(bfdUA:bb_2LD#N]J,1KL^^=2=+b1b@PA(a
TNaZK[(4VTI;,>CbdbEf_B_;&V@TbCS<G4Fa@c?P>S4g/,Y6[BPX()X.+f)6=g(O
:M#D7W?&bIKOWI&^@/b#_X;-XRbS8aD^C,U][(HK9g<U<d3);,2GS>cIJH5g-aC&
/;O0Jd7Ee47.B74:0EO]>E+/fY(GRe7Qf9092dbfL&eA9aW-U?/U_gb@VL<_7A/[
B@?E:P549\c>9G16EN2BL]b+Jd+PBWYYGYH6->g@5I2VS7/dQM1T4_-:H[T+9S;R
<+:-,>B3QWR(0>>\\;4/>3-MH[?)+=4+7?>+6e)b>\:1>0WD\U:LUd^e3bOUAZ,J
Ag_e-:dV37I+[F<:c_Z)PJcf@1/+T6G[a\]GK0fNKB8/BM]Ud^f)WK+[AP=L\:W9
-]6E[Y9JgEDc)4Q4/f4?=P?d4?C;D.(\XaHOd@ZL9Daf89f92b^7JeK.cZeE^RNO
7./.A+=@D:B#_SH0OfQ66&b\]3AZS+VObJMZA85A,L<J#PHBgNH;V9>1DDVR+VSM
DSP6WELC2.S[@CfQI8/e\Cb.b:\1cASU&AS(/BbJf<Xc<^A[O>G80b1.7)EEF@1V
?P=5B,;.]2\/1<1a@Gg=VU6O6E@+?96K\0BcN<fa[<3M/(,\7>6SM5d>RK&SF#(D
^;EA(J[[L2gC?@)8;=,\AaM^4fQ:bQN0V5+\(D2MN32D.GV5Xa4,9K?>S6X&HVd;
I;34W7LPZHT44_H1WW_WFL\G0Z_>[E<2bUH?#cd0F\(G]@GQGI7F49TI9_DN1RN.
VUgTFRbDRXEYT#VP4+/>_9E#e\1)D,\??Y9OKIZS6(;CHW+KJC91aNcW8;-+MV[_
c]VZbDWR5U-b?[J8O2Qc<J9^FJc:F+BJ4WQ;@cL&+[aY.VHIKEGBC[WKKcT()[MM
,CIR?8Z^.NGFB1?],bX5e[&8Rb.-,7>@K(8fb9(e(YD,f\G?fKg)e#;1&K[LefJb
2I)1R^bb;:FBb;K)SUgEEbJe>^.ES(^WA\IO)>f[^Y2NE@f?+CQ05AdTb=cE#&H6
I@XO6Z<&_1^T.T\(O<^Q>#,+7H1c/O]#a4MQN;FcGWX43>7.F;?D(gUJFRb=g3QP
Cd.Fgg\0+fM5_KREG#Ca[QFZ:=L8RaRVaE+:(4SZZL)NFY-QTC-2.DedX@X=WJc3
/]IVc(YO@90/6[XCDG]2W\?4Z5g-/M9,cHaW;g;S,T/&SIe=4I&])B(0U@.CDRf4
L-C6YB+YLH]#-LgHF/<X&b0N5+ab/?&R90)5+7B;TG>dNI\M>D6KE.@TL1gM>LB3
EBVEQ\gR#2/:USV^I3a8Jeg2b,_BV,W2,T(?dY+C[2Q9\JM\^AbHSV=^ODgE,MA>
g4R9H9#Z,\aW@X-QPe3T&I;=J0<+<&SS4=]Pf,X2df=_2FAHeU1Y:Sb::O)7)[M@
NTZ?(T#9TPL-[,F&;Se_RT^BQS+C&Mf:,ZH@B7.K<M=Y?If8)cAQ#d<B/RC(d+cW
&&YYNDdYX-VOUY=_O1gcQSJ(bBN);DeJ&?8HACCU3=JJ5Y=_.ERHYC_UY:\>R.0a
8X+d)PSM=-@5@_#,C:LEgc8Dd0OC/6W&3>ATKd^g(8/[.@,@eL6;_QA3e])_Ae=c
4_(B-D)3PcUMY[C1e),<X.V1Nb5<S0fI:9<WK@CJ<E78Fb#P31c^g<@=:f;,YX-\
<OH6)T2T[6Qb^,.M17UAU0N;;e;Sa=MQ@@W5Z\3CR7)6.dTKHV&R+X\6QPKWET=;
27(TLM9DQZN:7SH5TJ#J<W:f3IfV.c<LI:KH6,,FLV#+2Ld=(G\>8DCB.8FBc,N:
ND^d#T2Tf4XLTdg+d<SH9TT/65g_c75?K,O_c/F0]A&<.8e]0A\L^-A-Gc_Pg-?g
6Q]bRK>a3(PDH2#A;#?Z5=WJ:5X4K&XJMLVcSId<+UNBYfJ#N30Y.LWGASA4DL\D
d\#89DKHL:.Pf>NFQ8(d2I)1D<=PJUc<FV)<:9,^I,A/_G21VZe>,/[CK^4W4YK3
@MJ0CVWQE;RBE)Ud,H&2H66,cW&^^LgD(H>\aK4\;.&ZU14Nc_dX:K#9A<,3V>P-
:67Fa596(G4B^^WaZ#QC]PdZ6e]:QNLbK^CI0Q/<,^\aC;5=/WZXKY](4aB/G]1)
?</,BeRf]OW1>FOI4+K#37CeZ-I#=cHUZ5R;R:(C77;#FcFT#dT4KcFPMKNV<eag
@+e&++ZA07E@@VC]Tde<92=@_;Ze:.ZHPX_7Te3WB+e&C+eP]eFd8-&V=DJd3=RS
7Kg14:<0HS:6&8XDUb<NZ1O2f^\&Z?&)ST0ZP5BMU[P1/PJS&YC<MY,_YEdB+Lc&
V(_3H;=0NFK&R<]MDVO_W^fMAINJ0g5D(+O((g8RWFR4+deT_?]Z16W^>(QfdVAb
F9aKD+Ka^IUY1:eb67DJOA;3YX-@A.P-@2F#^P+,ca5WYE-)0@U.DL+))ee3M?;^
P/f]=O(^K-^f=M7H&Je;Qb<O6RV;=H24#M=CMJD0^+D4QeOHTFGGN(.AGdX<O16@
?YU#0D+=?QP^bY7:\5H),FeE8GV,U/AHUMD>B97&bE=(.fE)>PUU75#]_VNc?>GA
R<2fd/4L.?Ac>:SPVZBbOEJ\7>dbS[RFf8O:)#WU]Y/HXb()(,Fd]d3&eNZ/QP,e
RZU&9GO\_fN@a&K@6.SO^>SaLG8=L-HbW@)B[RQd+.bZ@)RA&D@#b5S&VV6RMUWF
]?N683aVd97TIB#ZHd=SLbEZf[:fW<F1=A>TSb:Fd@eNE21:Jc/(_&,YAR)\K7QC
].8]dK;R#gG=>9TN#A-f:@I4K<dGGUaA<9bV01bK&QDMQSO#X-CQBMeDCAgG8+KV
2TVL-P6?,D/#V7Q5C+IL0AZ/8K+/ED@^9SM28XTEF;d\ET0_fg8C#AMK+4707:V7
KDRBVEJ\QF8bO])_P1061UXD+\91eW7WYEK)(CgM^8)ST39XJ&3bT#<eLU32H?F.
96cHT/W8EHgc?fe#K[HeNZ=fA]/G#]-HFB594BP+8-<UM/9_gOB_PE]QJ/\_)?S.
O8=K_UHdfH[e+gZ.Zb4F)S95^?LA^dBE02bBIT:F-HZCHF_QMc=-1Ng.^-ZB#FVT
8T(5d/e?ZH#M<LabZ+JU4c?JCRdY43ZR8C-(1[Q<R3IK,_N;4.P?.LK;gSVI=S41
.<A>U++>a+K)CEfR<g,SW0\(X&F:+9CEY4fBc2WIYL0/ITO2[RLd@2NXIK:1<9[E
S]U@T\X(-LfK]P1(V:+K(I]9JKAd<J1Oe.88K.?57WYT5WHZX0[?>d0;I6)@(F2Z
UaAaY^3,Sc05K.^ZKIZ7W(e.?:<2GQVd3HW-;[\;_@RXZ\]74,f\QSV#A_\Y9[G>
7?f41BC:I7C^>A_>#L&E:g]?\#2G+[O:2/a.MLggbC\/Z<VK0NY^WK,_@NU9CJY.
DU36;dQ.J:E6YF8fC\TX]P,X\8fG?I0S[R6+SM5L;(>XYIeEANB6TLLKEf&c6C-)
]G#VQ.3SD0c11#W3EK-&-6,GBE3(3,ZA\7K-OJ<;L_W#[d>3Y?>O([R+?f2B&e3G
45cVJ4]T)]6/5^cRN:@2J_7d.g_]D66(=NEe1Y5R^R_T=/X3=U[R>4I/Ra2H#Qb)
6)[?;B>e>1T9M<<HgG0b?aX>K=+@6S^XS#,]M-.G0OK7?++=^Ee2B+I2M_#:W8d9
D3U)E[\5G0)@6S9D3NMfZ3E6=WWN+F+3UT>+gKeTP\5/cOSg&BW.&F5@aC2Z[?UL
#fbQ3;0aM8O/BEaPc#^5E82(MVS(B@B+aN,I+aM1Bc4,4T<d09/MC/<cXdP167F_
K6]:5.W]E(QT7D+=-VU+BFWRU.B+GXQ)SMEa(+V&B;QS:M#8;CE8O\b.+Qb=a_.)
TPEefcYX^5E;XPV/1+TFWL](4_;:?V[@AbaPQ)DP5=#/ZXWHAe@9/&LQJ@>0=HT^
#2[74Nb)gc/F@E_JdS^>>DYGZPJgZ(6f=\K&-CK3O1S_#<Y4W?0dZ.RVX5_-.,b<
/25&a-I[dE7a/ET(:Z4X1YSJd])3LSf&A1B+M95LH(9aW.KSEd-/11cR.g@SM^3E
<g3905W-SN7AUB-GOaeWXVCDfd26cg7?g)L&;>DC7IDO3Se9SC2bdL[_U^43+F>H
M.=>_;e9I::de98#I<76)G/R[J[&DaC3OEP(38dBUZW\MKB([E&=@GCa#D,VGH^J
g6b-^LIb1.a.J0L&J6W0K8EgX]_8_&N3^^bT6E.f2OH,49O&T+):AS?@YC:))\Q8
K;,M;HMJ+.6I+<8bILKHL#H[O28+^54e(#0:W+16/C?V>Ld=46PQ4TNaIcD9Tb,D
E)>O[[PLU:,FRT4<,KCeSfZKU/J\W##Hf/aa#K?7-)KA==3>>WXNCP_[:KE5:d:&
1@@DQ[5V1G[.E),O]BYG0@>R6a6cY1(7gb?8\U<??Ga^=F;K<eV/6<=LMF4W5]1&
MQbIDMX?XZ)gF>00=cXFDM\5d1aaIcXT7e+ID=0I^YfM7XPTU]:<A,=WSfS]/AEK
8OS/gScMSA5WB>Q/1bLXI\9KPE1N3/>gLVDN)SC-CcgWWWCaTOH;YZdU,S/&QQ<&
c,bITKR0Bc<U8:d4Ya-Oa-3E-1DBVRdI/&80R:fb:WPNPF6971Y.X^\+:/\AC/Z:
M;Y0c\b[<>?fPU0BODA#<L;HM<Z8\/IXFK4M85/2,I_Dfb0;3O1d^K^^^.2]2bVI
GS2ga_Q:);,egH7+MZ\F<aD&PLCC3=e[1e\3OeFNNH1&[WOKXS73DWeL]^>aHc:G
7^S04WVW<(4OX<M3W<SUUcSFMP#-,d-<Z]d=DW768[YSL^OZE)I?afSa1^E+L#NM
E^<H#-]_JQ7WfW@QE<-<NgB=5PLg5@G,fP&OU.9D-PPb^cK;Q_WT[T->W:VLM>BJ
L[V]SPL1d??8+.G\WG1XAD4)C9PL;_MS2a<da:aE\;4@Q#\+MeF2^P)=+_PGU_]7
,_K[]H;ZPPSME+B3YN3+\ZLeC-626N/V[bcQ>d2<3ZF2FA8dPTF#1<QZ6O0=(1XZ
D@YL]7g;X/2/(+Z;bIO9W?HU(^]R;Z6M()dBV4>,6X0;)TCf3L,.6KG[2@b)RDP2
@523T]0[@B?f#M1;6/4;,SI^a]3XbB1ANVT5GFd4cPMC)dNdV5BV#(3TS[UNX8e1
M+Z7)0fgU_/N=J&062bW[eda6.9X7L,HMNZXeaQ/74P/IC>A_DK1Me9=F\,,@4?-
T1N25W_f8=[OX+VF8G-=MO,:#95?,A2+NLc46,_9:)W#aZ\7\(T64P60(S)DeJ,6
KK>63\;dU<HRAQEcI=&X,^;U@M0Sad.Vb_RR5JPL3GG</gc1L&A):MgMFg]NVd)6
0,4\?\bKc&HGUaG:Y75fUR3TNDBceTN<A00&)]ZIOS6#&X7<APPOHRa;AWW@Q<#U
^>3#A8aR:B/;BK5/VTId4cA,?BJO,X@PIQ;LQ-<1S)Ld]7#8W\&0^:+&8gPg-SEY
YId)^3/5Je8;/$
`endprotected

             `protected
7QU_18LXF9>>dA6Y,@5KKP03/:RSBIO5+^/#-S^0b9eGZ8X6cS&N2)cLE):XeKb#
=T3,dPR_KJeGF0GYR&3gG;#5dJ7Ff,]7GJJQ1d@L_=0:[E4;=I3SORIU\CNHc.^)
Ib_bYK,(OWfG*$
`endprotected
        
             //vcs_vip_protect
             `protected
#W@7fY]^:267TF4.YNF\S6L0R>GScSWML8X#L(;Z]#7.@WV?)\eA4(E@<^+]GR9@
W;Ub.P7aQT?IJ?OdQZd-.70_+IJ&3OF=V6C2G(X1g+d3E]MM2gDT_[9+36e6dHHg
>]d6d@J#9aM+6HPO@U@aZ-??S;/+?7_/QFa>Y^CG4UT;@_IYT+2?XB9V)87,#VI0
H?;=W(E8ag>-PBQ+6AG#dYQNTTB:YGI3)14]R.VaG2TU@f?@4H-=/)W)degW1PQ+
HcN=-35d2Z5XYYcb0.<)63be.^4>DR0\JG/X>Rd+4Ed?VYa.C/47TaCBfOeM_4cS
:.ZRRVd65_g1HLA&-Fbeb&)a_e@HBM2SVU/R)MI#\TH1R_])dF6^GeILf#..]31-
BF;>,fNRLT2))18&Q;ZZAR5SdLbR:9SD)7=3FNVgH<5MbG8DJdfZHP#.=PQM&^)@
g^4]HBZ_aP0C64\^@?^BX;Z/d+7DMMc@VX2.S\BK]6bYL9S-MOWYRS,C9ONBV6QG
\#bZfeCM,G4?g)gCZ/YFZW5EOT7LR=H-[MD2d3P2?O0#a]6O4#IbJAI(E>M9#8):
,:S&L0fOWA-1cfOINBe__g4<(Yb+_W9@Y>G)e>[<]8\,/NA[]_&dR+:WHMJ@#<@<
HH^H/aD<@3Cd-H=336,D\=7d;L]?Z[d2+4B55]eOD&YCSS]@e^W\Cf&)g<;\Sa8#
:N4\](T_+7T^c26]R[PgUGIDSdaO)BR/]EX>f]@8R/6\<90N6&gf<4T[N\S>[#;A
E=O0:U0JW<JZ4Ud5_VP)5U\5:6YAaU^fCFf^fOJ7SXYC/;Lf[;bfD6b9T(/?aVHa
:<F[fQQ5eUEHY9.3O?\bKHGdb;egFdV#2J_.[1,HBH3Md3=BN0R+]AUSf_W49Q;E
DS6a3(b1Jb):.fbD;M#>7=)gA[;6VeS1,dL&\4&U=+U]:P?If@@bMGR0?\a4->@_
&+-0Z):_99:&=(VC@IDb-HMgGNA2R.#Xa/:DX<YL\>)EWZebV<F]/40]0,Q<.g7)
57N/J\:<K50UN<=1Xe@Z2eLa?bd2L&g45e^OW(T^M-EL4<N-4L?a1X6K#_-gA0gZ
21Ra77>F-.?0b?EAa_]GZ/N-2HTQ]6Q8VG=FCd7[,fRG#R_)Z[.UZ3@4g)HZTFEI
L]C6V13@\GO9@08FCIZ\-[UcIf1L/D-GF8)eWaKT:b?DIDXJf\Z#b2eR?>1?AEge
X<S.5&\I5YYe)_GJD8[7a/OVY3LCDX;U#XR6S9,BB(TXY]bY@+_9f9/JZ&dU,LIf
NG0-T;1H#PE0=62WQERAM4+]CcB)8-IgPI4DG0A4Lc]RHK3AN+2fTTbTZ030e]IL
4V[^YS6Sd@8T(BJ&9\IAa7M<9]N]@(d\K0SWEFdEWU1/5P2SKC@D7Ib22;Yc4J-S
Y?6VHHI1J0ac#:FCQQW]/OZcX_[Z1U>dO0Y08d?=K7^8(^D.LXAIN55PUAK.SVG.
eD##e^Y9&688UM-A?3W^a0Z^fUcbD>^J0.c\W54NA)?V<gYLJcJ\(S<<b2,A,8V1
E1&V?6EJL5GLg<Z_\QKI)c]=HF=:E?5?>AaEH[OG;0R\:I,Q-W?I\RRC)(]<Pf=.
=Xac]_S9Z[]]IWFc)8>Zf;IR0K>#8\4B>,/^]+gfPU;+AD\>G9[K+91Z<2)Q>J@_
2J0Ngf#JQL03;=#U)Y+1L&gGgO3[>.(CEPJC24IG_J>^:agK@N^5,:-VJ+:UT.D]
PU87d(85J(c4[2\Pe^H.f/96CPe)B_eRCAQ2>B:HbeH>U(2_[N-c4B]#RB:]U/9a
>TbV6MO?6(cP].7N_1a^2f)HQ:8WX_=MSJD/[^6(T:g9@#:C-V<.@>9FB>ddY)c1
FDDE&GFH;67G0f@[)K/^YY?G5bV)1/#gT^V?Q,c94ACZ.@SKK57S_YC1\McC2gbb
\JNWY-H3SSMRV.06K@L/@&Rf@7/(e?4OL8662)UJdOE\NPL#Z7).3-WJJ]Aa1e2U
5\S3UD5_fb#R3IT>@egO7@B;3UAf<27aW2P]X#fHd@MVa>INT9Da2cH^GeXX]-cK
5U5?.?JU<U0/R?.LS>[aIe8V93aQ)TG>W7_K+J@c)XE@UT]dd6ZE5ACL>>L+[RdL
E6YdAB5L=2O9QA)SMUB<#NZI4I2KO,DNVZ2E<_X6QO)Q4]W(AFUe+JDW+^?2ef_>
>)7c#NDO,#)&d.@N6BNB:e+9^??C6:AgXKHccILO&\dI#3C0PE#-#XJ7bc0#d^8#
]ScR::M&^W0[e#.8Z2S[]VK+1;GGSZA[;C-_=_@T#=1YdUdNBa:HDB-:a6(>FUJ0
4K3R?4A&R&(9#(CQ=8_-4Q_FY1?U:;0V#,&g(XUd/6Wa\#[Db/eYX.YMPK(AJX_;
[O/6Oa70E+J^.UJ[<bIRQ1-U[GfXIA_B5M4S(2P_2Kda@]HUYF?3TPD+HPOPA?-Z
5(&B_0RGeT>D/WKS3C6EZRQLda=-J?;+/C&)FJaKY^-f\g,0Tg6a^G)#c/4X>7PC
F85TYY4K3@Db^HW=[L:=<?\;;U4?X--(C10-I4EP?<8f00Ngf0(63/L=@Q&;4B2\
JV,>==<OYbJM\=9#VVEL-:9gJ\4AU8gK5WWS4B\MBe_C0]NGQHB\#;TaDAA_,<AH
IL6SQXgSH?QT/0)\T7GTO9#=6D\\N#7YX&gLRgddW/5P(eQ0LW[1_DO<ZeF=TPeV
VbV@-J(BS,BdJ:ZEcX3+W8__Y5R25Pc(Qd^Uc(;DJA5F.#A+fAaK=[JdQFR\?eNN
WBLHENCMU<.44AQc,:A(KB1,6eH>&V[e9g;J98)X_P)b[fG\5-7@6O(G5T#[Y+:_
>KagXNNb-]>QLROc.8=]01+1^<>C4aJ^ZcD)eS)[7fG3Q#(38S&OJ9DeSZ(LfCJ_
WSH/BNafZCT:9>#>-#3QO-&L3;#YHS>R]H\Qb&3Jc(A)EU[c/a?-XV-TD=86c0Sb
#dJ8K&Ib@5A,(Y[39b/1F(K=2dGHQ1NY>g[bE[C?WBOPQ9(#:&4O#BPH)c=+C[b[
15[aZA<?\3#^;Oc+P\U6RR@7[>XWGJ..E;YNJJ@6/YW[dX\P6#9>FbW3FBFXD:c&
,]g,Za+30>A4]G^TbGQZQ_0f)XO3JFW91WB@:L1G]DMg10_bCIUF5g-.74A6EVH&
N4b&KBdD#:OJX:&8E&0G9K\eWHWI>bDCa+a&(NagaU6PIcY#(6b7CWK>Od8HV(4S
N0F@;C4=XB@D;cOTC&\S8X[NEW1?g9JeR#<8g:D2E3c]DH(D+3+_YNR(BO-\gSMN
&;g3[=VcLA\86RMcGLd)<-#7KU_U+GC>O9G\U0#IU#?:+38]KBf^+HICQ^JNBH?\
O<aV0Td5J36ELP&1L]/c&T:?7=4XN=3aHdbF<=T7PKWg@-2Kg4Q-59>Q^^ZI;[=0
F&[H7MdJ2.dZ=-#1+P/\<@612g05<CE2=AE)SDD=OK[#2^46acMIM:+LRW,aGP.J
O7EFgQSS^;OP^)eXO921YX3fW1,_K]M;0eLWTX)W5.OY\I+B_e1?eCb.4+>/>cCX
6AB2fTKA?g4f1SCO0,(Gd79/C.YR?Z,e-e=F[8(Z\ZS5#/DW[2GJ8O(DD960;Mc3
egTV=4bO<?]([S<acW(d7a&9dPMBF))Y@7+9?AQ@UQ.ccPE0-^J9?eQ#-[AE1(3D
]_aE0I11CbA8(&b4b8C.._I?eC=VANg[a_A;=8=YM_[6,>>U6=,e>Wf1+-^dOC>>
S(f6ZQgES14/\Q733;V2_GHS-XII;dRQ0/UcT-Bg)g&54d)[<f=7L3d[bK?OM)Oe
T(T3HaII_/R[6#T6W_DEK1[)2?M1RW)eBaSD0>E62>f[EEgKJPf]-=.YT4)KPAIg
3JgVU7VcP]bMXKUSKM(X,C:DTEb)Y#8Qb0K0N5H1L(SU+3/1VV3<C\+2U#@dU3]Z
QVF45JG&O[0^L>S;KKa4GCHUD\P3+]WeVS[Z?0B?.++YgR(ZgJV)\8^-<5&^);^C
HJ6B<8(4.B3A=0SAR?5.7WgC1FA.V#S?S2OC;<YIg_<DV&FCSH@cTYVf+S=UA9&>
>-MILD\(IZ,QU,N0Ye>V_M0?fcbZT;E2?+8f9(?.H)B;,WI5E:(FL,(adKbA:6(M
A+\0LRAUURBg(b5M./BTZQ-AQ,U6VA#M;_fSXa]eN@C90a<SG@2B[WO1]@DIA3eK
)OB9R7OJCF/e<[e,9+M?AHA)\=FGAD5LI93DBM_7CM:9Vc(1L(/5/=?N@28(65RU
ga]-=A6_MY?WNQ<?NQBJ.3[]bc<+;:\cP,?;GJZgC]66]E/3AM#?(U1.f)?[<87C
>g+BD_^O<U\XeYK^=/2A(L,:_^3YX69=.#C.G_B1-&#QFIISF&CI5)GXV^W)L#5g
G+@d4#67R\Y@)9E?D?gf>6FD]Z59X3^R#8)b3gE)T+L-(-&JdU)HTGO[(bP-\+:_
eS[[DKG1b0D7OKU&&^>_)+--4X@+T.J&,FL40@RP]?Y/O+?XWFbO\:+^-G,Scd[:
LYdH3,9?DJW0^8dJDbZKF2NLPJHc(/W65,5?;e5W(HVMd)Cd4X:bMJA;Jf=RYY8H
\/Y[QZQYc3T:)c1R=-=H<WK1.JX@QfG0cKBKI0IE4gAA#7ZVNK&A.Q]2>.26KJES
(90#>,@]75@?<DSgJZcA/e]g0Kd+D\Wd>LCNWGR=49#b20?^C&MfL5@4f-7]gO&&
7_RG(f2S/(<UK<35NC,?_c;S?Xe]<.]UW?dPTD6>P:T70&O(Vg,N\.dL=K]=ZQ0G
\P;gceX8W(P[]4SMET&5@4_BF?&WP#cC(N/Y66;=I?AVSOM#O=F=NXD1:LHDKH;g
H>\AT:C)YMQ5N9<CR)SfDKg(cXVPfYX<MdT]C]^@D#_8gaMAdQ_O;A8a+NSK;_O\
[d)1EUaASS7[#?<2/WI198.Ybb.@ZBL1:DK[6>@EF^gC20>,>7D6A+BfIH=D<Y[Q
TTR7&16_ZBRe5=Bg\6&Q[3R_8edaV2^HUV(556641;1Q?SPT[R#J=DLUM]=I5\W:
80J&L?/C.^d2U13f&+V7-cYW3d#NUO.eQ(-U(SCT?3PMPOEXbF1?Je_eC-,,\I1N
>3OI&XW/BR>c)_AS\DX;&RH\fWB=?6cBLV=c-+Q:9L_Ebc[Z5.8=[dLF@LP^O>Z+
Ma/Y;QDdg@[1#T?KESN0,)F=6S9>HBUT8O&8Md_(V?[;&0T=XHaX&@Lb3J&4TCR;
_M7Y^+A]7L]NB10,:DbX2?<QAI0].7(9-/18M5P@9G-d<#?XY[cc+RA)Fg\#\H\G
d[37B2Ye[&c-]_Td@cJ)a(4[&&]7g(M[EG7&f#9\>b?[c=AH=X3N1EG8G@e^e4.e
bJe36?2aMJ)JY3B,?Ta+LEM02N#XdE#<#\Q,?OBVEU??28KU/AR@P;?ZEaU5SY(,
F.FF_\Q7RgQb0@I^c<:-^EFdBXW(XT]c:)X9D[f0(HF75dO@?gG(@gY687Z;d\3E
4/MM-)56K[ZP9R9QBKcL\F-Ua_)S(M]<a@bLJRL(.6U)V@G]c2FBW0<1]R+4WON4
;K5,3/+)NR4ee#_5[97YPE6L52Ab=A_@)8F.3>QSAOK>ZDVI-BR,[?W:IJI^a?;&
IJA&>9Ue.68ZT1TY/)5f1FXXb,gL,RLIGY/.R,\9SF[HA:1EB8Z1LZec1-/c1[&H
2->6+UB=<,EDDN@MJJa@6=@2IEbG6<6C/?Z7F1/,8^eYYQ>V10^Y=2)F+JRRg#+9
S2=A2=OQ7eQ(W[8#-U;AO-X716YA5[2\JS_c@Ee[;[1D(U7N[>&Q[6&H;LCNF1eG
VX2beTYd@6,A5GND+8N.X/UH8V^X.P1CRNA8,eN/WcLJ@Z=g?4Z=bF(-6Vd,g9/;
<P\#PF8+^f1,AdFDA=Sd4f@bRd(C0W?TAgf0)21B4P94?=]0@<MPDDaE[(A7);A?
KP]U),d_a_HN5SNg6TfB-b)TD/18_.?_Ic&_APa9D.[&-Lg]G>O&52R]5D2C:EQO
OD<JT2bY;RV]cP_;:Ad:GJ#^>3bNCNJPE&CCS?+I9NNKb&KfV)#?9aUXg_PTMK7F
P3#](#6?/^5>IZgVTVg=9/N;aQ-UPFXe^TJ&8B.B/7==PQYZ<2fbJeAdF+=^?g5[
506SdN90:g::>0ZF_4#,.(17)F5GO20_]V16&bP>BBT\I325EM3=_H3I(QN1YI<&
g<4+ASHTS-\3,SROMcAO-X,A&V,U)Jg]YCP+U2O[-GW>B88@a&KISKeQPDQdE-O-
H.3I44WEH_[-[U.#/LI(NK?C]96G]?+,ZA(Q.K3f.UGX25_-eEX#L@PWX]^<M2<4
HVQH2c1/(CNJ6R3L8T)#8e(;6[DEC9&BfD:&BV\EG0Le8<aS2].14I6=DGd8Z5e<
)/YQaZe5L:c+Oa_&.27+7B0K.5W@#X38YXDQSLRe6.H;O(U_&Z-3(6JAV?KBZ[1/
HF?KXAg9+XYQK3QOK_a<?M6e3A-KZC[TFIe11S2,Y4B@HQW7JFD9.gDE#;]\K(E4
PfS)#?+17L5.3f]]601g4E01VNBU]N\2;_71CTe;E6[+8RIWbY[-b=+Z>E6VX3Aa
NUNKI\fDJIM?_\,N:3Y#G>E@A?=8+cUg4F,<4aWF_/KLF][:@RA4BYZY3^+K&[:U
>d(2@[UFZ1R>I&(G0a=JcBJT7>T7>0=7A&]GJ,6:+:=HbUJ:U:N06bL7:e=_\B[(
/HUd.MS:-Y:3T5R,]\=f-#F:.G>F@7V[M3SdUKR.5T_LKa-Oc>7>#g@?,M.D4V>@
FUS@eQDK:.V#2VQAL@D]KU@R@0@XJ,X58Na]G/89>Pg?/\?>MfZUW4&7BOVZ7IU8
.?JcbdS1R;B\2K<R.V^6.\8SRP.C_^]/D8eAIg=D94bB.,8-&N_CPLYXEED#CgC-
Db20EVNNT?4M[SWJ_:DgB#6aYI8_;D#O<@TNZ.Z+8(ME8C)H5U+<0NE8>/e-;W9R
1YGI23XILH5#6QK\T;:ML1AaTJXZIAV1#.CRMD-)L2?T+@]d?O]1UP(K?=U28=ZZ
8gJ,_FFe::]KF1E1<f1PX^(TDC./GB4^I<.W\L)6W;)F(Fc18NOQP+^=#=-6L63C
4>?U4],EV(=4O-OQ\;AV\ZQ6R3?Q>(5EF;JP31QHULa_@?_BFI3@MPUd:\E\a\2Q
)IdA21U=AbWEb;14+JAGPW]FG/0O6KeIM@08LR5(aAcQ2:.eeF=-@]8E9BQK_ef[
DeQ)Xa9]2:Q_]6P[M@<;/\[H#:<VLS-;52]D)\e^6RVK@DODT4f\ZS>ePAO:@ZE8
c\#8BF=0Wd>a040&\Gg#Me3aKB<(QGOKd4]8JJ&_=?;fUETG.b_KK=Z5[e>+.2K^
S?7-?:4FaUV1Zcb(;27N_XX&<UTT^,C?(XT7K;G<)&XX3CCS>?f=<S?Q)&eF0]Z4
ABV>Re:V&&1MB,IHK]+&-=E:A.UU<4U5SR7:_(DXcR1dB8Y-=EE>XV@LE[/WZ,K8
\(/bNPRCfBX,7]0cFZa>V6gN?^]5B6@[/^I-GTA:45g^Y@VbOVJ3c^WF+SJ6FbEP
?+WL;T]EVR).EXMT]AHY;B1L92X@\Y2?fOd9.&?SZ-5HF^OSGH_Rb<#:b#R0Y&[W
d,MH))G[M4)22EQ]+,&9:SbWY+FNJ&3^GARU1:_7&F\RI@aFS=R>c>0@DV8+#Zf@
W7IBJMXRS]Y731JG]>+aa15N9c,AI[d<W/?DS\.Y^&Y#Ta-.XN2M-,J^/(=U.VM<
1A>IXgNH[N:ae,I)3@CV+#_>8cS3DEA/e,9TfNN^(OU>N3a+d@g,1=/0:TAM=9##
-Zf/&)-9Kc[V6PW@eG>Z:2Pc;=8]SKOC+@a;J1Z9G09]K=;/;MQ41WWOHM85Q0f+
XPDI+44,VIN\0a)(9JOSZ7#^#Z,AARTU,:2O,>GR2eQ6A#/LXJ@83<Y&6T4V&OIb
YadRRY6X<FJ]ID]SQ&D<50Ec&8X3@/6e&#Q.2B#_.aZ]8THCa,+4P#;b_;)GTT,I
,6L\4gB6(cFB>^+PY15^^E))D0>FKFP5\Z=.W;6R7=((SFTK600<5819QXfdC7VP
#]G:^8g)7E(d(G08K]F?K__g@EKEcKfaI\U3E/5X=bS_8NB+E8DgXb#C7^I22QC7
RWW)OH7Q)6N/9VRH:^^Q#2BL@5]0BJ^QFUGA)B-RK6=6[.Pf?35-_5H9^8K&FO#@
.SQ2<\NF+#W#/e/+]/=C1>TGYC>?;fGOUW6c5VS.^Y99TT,7f0JN_e@HKQaCggQe
XZ3aKN?O\J6[SO\RV#0^FLK+\I<)#H;AIf]VEdQM^L];#d7C8;/A-[cV6a@.F.^J
f:S3\XSJCQF&^[;^<XIHXY0>4=(RaC6M&_NaWW42B_X>?T]XW/:S)2;T5I?DDBf0
3=ZLOS3I8T-W6>>8=FO5Fddf+\J3,P<67J1F(7TbH]KT<g=56XFMFEb,\7K4U=^c
P&9@Z^4TUE+NRAI@[Tg,6_+c:^P4Y4JN&;LCY,2cD8ca1H.YAeYdcN0E],KTY/XW
Z)3?0].&WLBRQH8D/gdWK^7B^g]XGY5[(CMRS5?(;^E&87Yd6JWN?QH)WQ]gR5@7
/OU8,PVVJBO)-B@MPF4W2aHFDg-?,Ic@(=N@B#:ZAYQX/.F]?eRLNY#/dRGV=JF/
\?;:);@.Me@C48Q=9Xb+(U>.W7[/U\EcdI^N+cX[ESaa;=Vd9F9(8e4G#G(OLLC]
_/+#eFPf^)3e6C<9.3e<fT6S694A(__d0=fN=Hg@a]>#fIfA40)?P6aC^GV?(5d(
=Cc_<)cD[KV===XF7_&c(V4YH=QFg?8<B/4]P=)2L0/DcQa8KG5c2-(&/&K?72f4
1S.E4DfcZHC;K4EQC<E>O99VF?.D?ZTZcbbeIXM./9^H/7L6D=?S0<&_g,4_+<0@
;[?O##++:A8=M@d#)d?,Q41)@7Y.YK#W^bMGGFQ>CT([4bKf]O1(;F@207[V;:V,
C68e+@/5MK@\2aI\RQ=dPR0^2O&DP6>b9e,#SIKdQ0-Z66I=?7E]]E?IEb=TAC3D
LcXF3J4>)PA(?FXFEQ/bWDg?c:[>UfD[0(<KVgF\(eQed10P#83gAXgN@U5/?g?c
RcJBJ)(H9@3L\R3f-\VcES,D490+)4d+VP,40U2(M=UD,)H@#6VPe+]DS:VWT50D
=-HF0>U+ZSe8gIG<9/?Zf7#R6KB:&/8C;>dZB2YZJ;VQQgO_.OB-X:=UF+:=]+<d
><5N,WG\_)#C89LbKJ1Kb>W0?_?0),/2ORI5U-TE6\9F5(0F9+?<],.O]4YJ].DS
VW_a>db(9QU:DZcdO1eeY80Q&aad(&WTD>LdVA&L_7bPIY.Z?0&&[(X=3=/g=DJB
4f8UPQY)49D[/@\^LCS:F9U]6-.CD-BMc>A:V@ZgB5-]FL17ccR-@HbMg&UPTZdd
S(UbN@O]00)R10.K-[.G?RLA-TL[8IdA8995e6=,?F0I9G7CSR_-AG&c^N<9Z8Fa
VIO]&\Af()^;RI,^b>Yf/g1J_[5@<__(/>@KKBLeRN4KWQ>2()\NP9>R6P&Sg^5^
EI)Rd0G8?9C^KDW\4=30=I5WdHfY0MOg,-2#U>_[C?UTO:;M=g9U<6?IOB_<M\C)
NQ9\7EaS2@LJF/H)QP>MC0@@6?_YY\27FG9#._K?]NG[UOD&Y_&#.K7fZ<P+GdZR
\(EeT<d+=)RNWR8DNBKSXK1]a#Q(b+Q(LBKcYU<8@M5^^E67[<:VPLHH_[4_(Ha6
,,cA3[\eR\O3X\U6a11Y7CbBDPUcJVe7;cQ-?+_)XOQ2/QBLIZQ^SMaOE6>L:9PW
.gPMV21^Z6S;#Q.4V93eNbSZ#,^BKUa9R^PY.eW;2=4ZBa>U[-7KY2MeBJP1:VH[
d69WB]?0RS:Ka=ZUP7fWNfH5QTc[-Z5_F:8/?29X0V9U^0F_?C4:GYQ?[-;@eIAL
=_J,T7@92Z4(eW2EL)(97(EM[R=gea.P]V8=M_?ZDPc?&JO6BKL;Ee0@?&EJe-@^
.:;eaY@&J>dHb4(bIRT2XI6PIL;9W)ZRGXgKN=R>7((+NNK(^.8f?HUAWU(ABP.W
A<^(9d0QH#-fZ,d8[SeH:L[<5&6;;XI=4+)]dBN;<gS>])KJ+CL(e-K_7A9Aa59U
H^+(EWIc065g.([\3N5OR;T#8+BbbB1_6M.,JZDIZ8S:,1?b]@&>f_BMfPU7JCNA
)BD?72:Z/N,_8I_g+7>\UOB7Y3L:_YCC8NV2IS#HSUfF+>/T/:L\+Z;0GP434VEZ
\[:/87d^>C3_29ZME9W/OKG)0>W:WR&D8G<//Z(&556EFLU^Sf.eITT\ARNTAWGO
CcMQHK8H]5:M?<cA4ISOB+3^G/F]Vf?&9\9M8ObA97@aG1<J3K<754[]?=f_ZM;.
=YA,?\\F+Nf&.Ig,[DR=B6N@IVc.G2Fa^8(KMWU-WHAG&TN0^.\U,O>D+K5<6U:G
Z0^4\@7??NQOLHLdaOD;S;.V8Z^E0O)_H.aFIbI5KeZUdbG2>IDTA:b+H<F]&c=)
^7(=17#B;C?SD80^01.6@UK6bcLPcV[K1-9>9:16YA@Wa;._^]G64NWD#Q-;Nba3
+CPXP]:[HC\.NAf32cWeX5P<P4\XO7;XBT1E+,IRUX\1(P/be3.f]B<L><()#Ga7
>b;0\D^b9H@#D2fD.P&?OLW8-D3]UM2b_2KI;V&]-;1_[Pd=)J\K^\V&L?<ZX?@=
?K=_;#bS&QANC3LAK8R8#@TX]#5c2/M^>S-T7IeB88P6.IUE(,dDQf\)R)/14SA=
Q0/D@=_RY_\Ffg?DRR]Y,A^a2f6]/TA1f\...#5,Gb[6N,,.V,d6c/=HNY;eBJU#
8TGgTIZVO)?VR7SW(._K?e.U,C193TK;g>K_2UNP6a[K6WC>.,_:;[9:_[6,RG#5
&BIV#;g=PA8O0Q)5PKSN7JbOHA\&<OC6K4--<;\VW#]<I&abS1TU&,.](G]Nee(I
DO524\SfO10/(5QW6gb3g:)#\9;^^?MNEC5#;Vbf#&PeSF#64A324@SNS=Qa38Y/
5K?Fa[Ib:J;56I4deBIHBES<_#3>=_</A6;V),SEe_NFDVV7[+f[2]#K0-SSECdZ
TZL?,#?>4[-\AOU62X:g8U,U+5IU6c70YU2_;bf^I/,a.LLHcJOSU9L#bM/[1&Dg
e]9Y9NNT:I)2KB8HX9C3CaSa@LfF)ZA+Cd&:,<c7g63=bSWG]DR52ZA]2Q:<)(2/
Y81R=?Q:M5AR7)AcXL(^?L^IcCRNfKTFb(^J,&E2&/M.-1Ef4f/eR_3e&IO20V/(
P3D;HNS5#.08)K,R5=>AT\FJ#=SW.gH=_&R](/V=f7J2JT@K8R[=8K3S[4=GETY4
f&KfAQU#N?+17@F;JdJ-6_9PTN1+KGFe?_gD?V=+f+?1XcN5LB4d&R@4<UF:IFQI
??<]>=]bGH&XGLO0)I5Jg^YFdD4MEFaB2c0J>2=Q6_B:&e#</0JO@TJ.GZR0=><A
cW-HDDX:<WJ2FJIRB^;AWLAfIgE:B5CO^#5?QF:U114SLR_V+-c32WV)RN&Nc1/]
Y:YeF\RTW?g,X6LE)1e8e7_Ga=3)-9?IC8>RI@??]S\?6]1&)JB?]#&L)ZMPdf&9
TYOY)8T))HbFgA>aDICdP6H0=/Y0_+aHPXHA/8MG3a=@CO?N+ND&P/Q^?=Q#QcM(
:K@NIXb&(J0@WO1^adRU7Ma(G=Q\^F1eReX/2?/7Y#4?.FS2Ie&]<^aPL<[NWEO;
:YW]HgD<PE1B6VQ3d.7PE1G1#Of>1ZW>7.e>8PGEKT9#TYKIG^U6@6\X86MVXC6a
]fc)4(9DN7AW5O]C4Z8GXd[D&_GfZ_NP/fVG=->7bc9\FcBX.N+1Q(T3W&HAeXSY
d3WU9(=+04J?+(d44.NPaf<]0C_:T@9_;6ZQV><<E]fIdQ<)LHC.8>5=bG?TK>K9
-Tf]XI6#[CX[[[N_=F([9?aP7OZ)&/SM.WX=1&.<6f?6_]5QeJ7BUGD>LX<?SGIR
KX1G#W^,G<bL8DNV0JPD#\540.6aBQ@Yd_<;b6\bQI(\W_TQ9/ZH6&;8dd/dF32_
^9HBW@I\M>g,b>Hd1/,)O\b+\X(M;+7B1@0B>439[Yc4B(S++WO+_c8=D]AI?N7)
5Ifbd[=R=E^_)+MM_&dYT.=#]@Q.>X2,KI+bdeI]&=:0?O)Q@E]V/WH/39dWO-[7
2PIb\3d:IgN9-,Q9[)XSW_cLP.N#.aHf;4D=-@dUY_[8?Q+O;dH;GK[BN,fNNNBW
V;5_J4N;)OM@PX)QCOJTCR32O@5Z2F0=DEB()g<;Na5^#\Te9,E#5SF[.I6)C/]9
B\XX5HA/3CGK,6c>((E^29.ZO-57Gc(-M)9OYIOX+2:9?7-.]AJU#>Db+3&N:egU
=)1C5AN[XeM-J<G]Y(RL_#GcG.L^V^>WLgg6^6aX4K@c59=,9?(4-1X-f]U<MFSK
H\OE@KRSJ3@&&WSL/I\D;Z3fg7;CEF@,@-)>NL-,?gD^>;MV6TF4.EJE\QEZ4)OM
TMVD-C,1f\DS(DPa[FfGV7TL+\YA(D3XX_PIV>&<X5VPgeLgOgg8FV89]1?^?1Id
_M2_Y-c:Fd:OD(#G_\AY;>GeT]dN#N-d[]SDG1:P#Q./+LW?afNX;./E[#CL?a:M
AWBZ30Hc.NK<EDKNP?3;N(0IgAD91P,7Q93Z>QH\XW(W4TYFfa-fUf\f(<&L@IJ<
[.f9P6F#2G[;N7^12;>+.fK(M4C<\WFX/286RREPD-5L)^0.3g<,gcL+_?;.EIG@
6)B)0OD(eUI&]#_6cb3_D+N42T5@Y8R9GMDQ1V@d)K2S#gY;dKL:34XgEX3_3]VK
],e\I(S0>/EaH^)JgdHZQHL1QT\G<5:_Z[8/8S5.>IGcDPW2064K:K<=RLV7[;Kf
[QXW?O1c9OX(Lf,>0G3Ha@d78OK3=C@c#Fa=6G\6_6T-+V,\43N7<R3NJdg1DHZe
FUJCR0):0L]YVVeDWI#-2[eHbOXa-OJ5[V)?\E(^::dJbNV2f,,HS2X-_f>GfPC8
(a0OL8A/OVGB9B0BKX<6CWGS-W0d;I[P2;,.F&7KV4XLJB#cGC7\O[U;E3[AO:1N
V/]24JT;I&PZg2XS9@R;(:.?+XD,=E-WB#g)Q(SeUU][4<b^;T]<]Q,0Q)9[)P55
8.WcRW[;_gQ=59ECASQGE^M[CDZS/UcQ:UGK9(CD3f1==@+a7UFRRWcLG>A:4=C_
]HJD/[=O]BV\=?I+Ib2.^3E:5&\P.fd>dLF6WWe14_A[+fK,DZ=FGLUg3#8]<[CO
98:JgAfX8V\&&JG;&:Z/ZYD,bLcC?QDd1K./D8T8_1Z&CDR2Id1J;IOE9fSbfSdb
6,/,\9]KPb:^<L+Y9HWVga1@<Q,)F:Q7Ad&ENGH1b>/:/VA2>\(g3e9=E)FNIJDa
G(E.SKd+^,O?(\0Ue/;[f.9Kb1PZcK#fXRH=O9aV)b1@c.38Y<W599/&#b_-9dVf
+gH[8H=HZ9]UB]I&fU26VMV>Ad74R+Dgb-1fb70<6#?DT]f)BdTeag&TI7X@6Xdc
+:abNOO4g-Y:N;:fC0LH1+[+cD28O1/QEF\/9_&;\8dF,X,6NgWTT9Xd(<F@1(ZC
BT?I_.0<0D1WS51P7,S3I3&gL\=Df=X[X5Z<6XP4d@WVIAUYBF=94_O@6Y@N0:/R
:JI2W39dX59^D?3<8DUFQC]0;&Q/;@JVY,F@)JWXAXVC))]LA@47]b3ENFPMYE12
?a#?F13YA(UHR-J;#/+W3IbSM_1H::aaNCaDG6?8>OfLLDX)C.bQ@&C:[4fO<JIQ
TJ<EI>cYCf7b8OB.&(Q0R)L4.L@?D7Q0Ag[5?^b0d8/+]&\Ac@g9=-&b-4.aE:(Q
\_J-EJ<+36Ia@14&[@\+Nfda,NEYBB8])0:6I0b=N;>)ZHgY?\TN[I0VN>Q]bT=<
-9Y)O8V2/2UD6Ma@8f=/M>COLGY/5eNR/5&GHP>59ddA::D.bJ1g1cb[K6]d1#Q7
bad>OTE\^Pg?B?DCG+>2FH6.#S7?GT9I;PHg9OD3(-EWH2JWUegE,bI3_Ie?MLa.
VKM5NL?0Yg8UY,@SMV.c^B3?Y[J8P4_TecEd?F^XVO4Q+3OPE>aDKLZ7D4TACc2:
E3:VQBOYF:JMSGK\VK1Q,8e&;fK-6Z)gZ0MdL-T74/#)BLDMHLUQ(\R3GcUJ.c_C
E)UO\N;J9:,8&3>(+ZNdSU&:D58>KO+/XKJZLAgIYV)[TSWfX]?T+Td^45BZ\4K2
_OfWd9#7;4J_^+CeZf@D9S92SW)A43[HC6eH_ES#9?/H)W9C4Re8I2_W0AT36La5
WUX\#\WRH-(QV[)=2ddW&/b2^c]c_9TFQZ[dD+MX4YI&3GH(a0Xa;2+5L3P]GUd9
W16OY;gJ>JM^:OMcA&c7MVQHGWFb1-K=GfJMK#H,I@KF5LMP>5cWF+;K4(T,7-F8
^.E:f,&fP)WJ-WOU]TM&b;/0^T595OM86<5.T0QPb2<OQ&dN4>B&;JMAFa?7[V9G
N[Zf:S?,_S[7Y><F7]eW[;OP-f2HUR99H8+)JL4KdCg#I(.e6TDR[4M3UF/#E55C
fTUUA566->.5FSAK&GP1Yf&+J[S6QXgLAb/ZdbM=f+&>b]D&-YHa8da<#MKb)>).
D9.f#Y8?,OU_=;CZ<(7,]Q5cLG:8+)[+B14[[D5/AM[+^)a1,;E^FJ3UfV-Z<6DW
HFg&8D8J7S=M:NRM4?]9W8J6S[C>3ZI7(\)Q/^((Z/0cf8-11Z)agVbKM8ca[\JA
4>05a;S>G3H8)&@&\gg&?U#SB8<T,_WZD26=#gN=)6b+)?b)^,Z20;<0=ATT#V7V
12O83\[&\F3,;@Y]20gE_#dY_&5VLN#b5+109+B=]TaXVR2QNIYeHO#-MI79,3T[
>bR9cHfWcfIc7(:CYG^#N9R?-@(fU)?+(7O(XWQfWY^7eV0PeS;,(VUf=;<Z042L
30[/ENc5-#aeZRNd>+54Na/VJX,98&_S0Nd=b/P2@R#0G.V+O/Z&K#a4P.7;F(Rb
K]]#&>GJgPD\QCL-aOCF8g+HE:3U,K5f4W_Jc?VJV0>[U8F(?Q>b)XVYVUBK1c9>
+6J4<2g8W:X&NLdG6eVP?F5@2OFg(41:B^QQ,_BQ=O<Ac@+>@H@bXdeC>=a9X6a[
-.O1;0?;MYIQK]_^^5=\].^IK,Kb;eZX6LD03XJ,[f)F_\Nc\+;9<6\e1OZ;>JL)
3J<+dO5#C\7O2,_.a./,G63bdM9V1g@/DHZP=;4c.0.I-XGS]>#GaR-2J=2Q69^H
.8S6QW@2dg\.NfCKCOT9BFWEREM10^?9(-]0CM;dJQ0X79aVZcERBF)e@PCOXY<W
ce1[&Z@=\[\b>Q1@2dO2J[)b[eO15K]WT@<\XL/[SXQW4/;(K+;@-7JS71=,W]K?
_OE+Q&Me(cHDK))5B88U5]ADAG,Pb6+[\\^=XZ2H-(d\]7:dP0Q7@Wd+/C8&d+(1
bLGg)/7TbWYO:;dL,c8#\2Sf/56O3U@Z]]cA^;C\b2T:PdTFV7-JS4Z3O++&KafP
O.fX6<:fQHb[5N^SK;\_+&W;O/U<^&#=+#FfEQ,&.OfIB)S:JB8CLf:..9A-D.6g
8MK5/]W.-Y9H/gY(Y^[e/9]4XL#D:(TW/0F]\[gaAdT^:4[1HR=#[)4Y366U@agK
DcdEZJ:YBX>QAQ?WRASP1UdSIU=F/aL\+[3gCXJ6(&C8DXTKJ5TNa8BDWX^M^gaH
P[EB&)<5fc#VTG<M<7K2.T]DAR&f6&.gI@+-?a,C21)]1dDT>E/e/+-(:^CI18L?
^>_UH[:M/A8a+DXGQNb^-DPaA/3g>bX/2\J@2;1Q]UP.7NO_W6(^3VJNQ8FSPZRU
_L]\,(+H0>F)).=+R>GJ5+RE+JLPZN=+H=;VE@,IVFOL-RD6>&6_aI:9(fIO7TMa
f.K^NCZABVY=JPKJM6\&_6N5K)6SK3^-7.K2&,=]f/f)9?E4AHf=JY:8V&gW\?-@
T&Z6eQ+>@=V?gO2KGaGP8M4CC2#ALUIS_)52B.6I:HBgREfIIW;4_?8P\M4VAKLT
;fKD]?UHXHgC<ebKf89O[7E@F5>#cGHWPXGH/25:V5,I@R5Z+W?#f5BF._X>UC.M
II232\P?VecENJ2dIP+?d8:M9LK1E)Y;+1-L4]1[I7MP,A-G7V>Kg369-Yb(WY&)
9UCI^,5>_:,IT@GP5U&#DOUBb.M[+C;GdP5gTI@\PN)gN36LDf:PHQ7ZY/D9&T@O
\e>1P<N)6&PH@U-^B.7/5g:W6V<=Q/XFYcFRLXcF<[^?=HQ<99#H=J2dH:D&1B6f
54P^)IbAT:(UG-_J<#/55&<Vc1I(cP6-.-dVAH/,_c@AA.-Oa+G<4-6JK(D&g^9b
.N>0>M<1;UbB9S3I14?;fMKfF2.2@2(X=;O.0T-3;&K>R,.P)Kc8VcGeLV1gYLVc
U/\;.)?OO2f>[8)>S:-a/_H5U,LLBU7.^RJ(_>c@P:QFHV3EXCed>a+T)=5XTPd@
?ZB-+e0OP&;eOL)TJ/R87HC4ZY.B-/TQ#GJ.=7feA<1H[HZEKYHXFU:;Z=)0ZAcT
R+Y/==1#04#/)@^>G;OUTH+/Z:8(TQfU7#SC;8\@4(V7?1P+eg+X3gg7+W[bcANg
DVREBeV]WV&6ROA>-Q+(8d8,R/LIR,fH7gS:PcB;LdT[.FG[a4RBa?B2,9RV,PIW
V)dc=JQCWU/R/JJQ\;KD]Y8b1/+1C>S5E^45_LX5>afO=.>?GQ/XO5cV>)V5FHP2
JE#;C-ecg#>-35.YP^J@U&?NNM\:;78QC3a<W\8Q)NXD1dG+WMNDf)bU)<D&^Y]B
?cFSeVB>O+XGJQ^EV2gA]M3(@(;Dg(#F0:\]f][JOT(W+^8acP3I_Yg=/KKFf1+P
S\G2XYI&+^aAO2J@7D2[GX9=RgSTQ+<D5&b&_K=:,W863Va=1R5/Fe<c7b@F&P#9
K0c0)SV;,cN5UQA]_@^+_F\^/[g0PcHP[^e@YXSOU-?ITZ9^R.CKaM.,UM5F0X4/
=01XJ[6AOU@J\)K+.g6<8-<1VWQUd#VcV/Z;/K9YTC&1-GPQbE6C^&4A?4Q>6/0(
@LAF79+N^>C-7NZ]#GHb:4-:8M,b\&Bcg>Y]IJ]8Y5dFfg;[ZL=-OS)/>KL7-]-1
e._=9;N]=\8QQ0K(b433fL,P@.19JVA^?]0ML_-_NYMcO54:&dWBc8Kbd&RPKK4,
;IeS3?A5ZJ^EPBNb=NA6(cTGIf2.R:J<U_e9QWEJLaZ3Z9<5F9K>X/[0SKL)6\];
DH:H5.SJZC?]H_R;7Q@+.P/<4+R(Rf&:91FF-fYEXL54S6d<R@J+&_<1D4-#Mg1S
9EL#90CZ5L#E1JacK,f38PVd/EQ2VOdZ)gNURdB(B.^+_aR9Pc2afGJ4)/R3[X:W
NaNI/^KNT#BEUaF9P8UYa6DG_PA^+KT1d(T/)K>H+C4D<WN>01?66XQ&+2UO[<E:
]FZ^\b#\&B+VG[TWIY5S/a-YGGfEJdRggfM&_W+V)+?:,=ZBb/PEcV.YP=e>[+0O
4JaSZg&+aR6Y.\N8#MEU:ZVX+<SI=)^EECg7_+2/eM;/bEM(_Bd,O?@)>89RJ,=,
RNB[-f1MP?d502(6&BH2-Y>P?<LLQ?T0[GT8^>aM5]GZP-4SeI(9:@9[aD&6MUB.
GG6[^DMgF21)Q6;<f]@]3#7JX3Ia];R8=Q-&[NFEB^(O18UT04MaW6c8H)9OS#N,
_>\M=dXM)4D),2a+g0;cNe1P@948(:N=HbAA6KA2=6\+8O@;PU:X?JRfN0RE7H+A
0H+/eT^4HRLdgW@QbgCJ\S7FYN)4fC6^6=cEM9)&e]Ce.dL+IMbX_3M)M13R#\Y[
[/IX1RMeWUHK26\:P0aG+(U6KZ?WATU_N^/]WM)]UZ&[ZVI,DBYX3@V08UN/V6EZ
g,&Of:\@2Fc&;+BSG=NEZHEODBefg-Va<T<M>@V+YRP260?Q#/3G#?>F21?(HMC7
\)7HC)6,CI2Q\[/cF/Aa1_T+b/e1ORg9TMH6I:E[#F8F+aO7(Xe2JXcU>/1H_,4e
EH7Y,O]&O2@feCH65g072bcBgaPGa&g9PQ,;7L)B_dM)3XQ3)bDa/2+aAb<M#>V&
+,X7;PZa+/gJ0f.O+&H]c,E]KOcL)ZWHVT7(BONKH^>Bd:KS57L[dL?g4:],J)S:
B3E^L[]F@9I#9(;[&XB/YZ5]X93(eXRC8[<U(Rg=[/Re/W9-g_5&@=.\-L(2&+4a
S>NfHe6^LN;YK;efW_PWc@Q8ZCN#1OYL>KB2bSN1f7HO(JBP\=#_-Vg;\6.4Z3M5
df^/FaUJ4dLa(0K._8?FReCPH:e[,NYI\gCSC([D;bU?b/OAFYe))Y,<H9].^.ef
1)(&&S]K4e(TUBS)[956LZ_-D8Df#9WV>eQP/J_3\>6MXXbE5:MN0&IK+3(JP<\K
<I==0VURU,HG-PBG\CA7N=Q(^M1deb3+O#G/Ga2cfZZb2N](LZH)?3^M.>efK/=2
Q#,:D[O:YaYR;;eAVP@IG4S^R;fa_BLdH2^#dgaa>7,RMNL8Q7JBS>e)HRCQabIW
@4]>>7L1JN__4IbGO<@EUba.eNS;^8=^R.ZSA69BO#8]A2O3ZL>EfQ5:Z/8\##_F
BZ,+=L+TH)Hb=DP=GJ9YHRDd#];CPY2PNPH&0.0Kc5I7YVA+LI2+c?=^eU6+e5++
ab0/E>a^+d/[2b4^4&&W;Eg:37U/Gf.A,X,HW/GB5F5EH&d2=&NKXYgb/+71-c_9
G=@(DW])ET\15\68Dg.gDbR(>6&Cb4bRcT97KRPb7@G:8g:@M1[?GGWP[=1(33X+
H6gFSfQIA.>&ED5D886P:Jd>0bV?Xg&MB9[f#ZNc5MZ77d2HX\L-SSY55I4Q^^cX
#0?OMMY])BMT:><S+@Z>FF2J7gXB-OBVCdba>_[6TQ2e>05\N5-ZK,4^Lg9=]FSN
+HRc8^F1+1e-YN^a7.YXXTA+(12Z+R5#C&\OI\LXEdEN0L&;AE>MURa<M,<B,0\P
_4R:UTK&.(?2C-][PCdWHXQC-R0^T_4CA[?^ZT(0P4K\9)[(S\g1<&;<9P-CD9?\
OFaEW:82fX1X\;U0FXF1K@4RF-Qa(>#1,2-ZbF0;UGaZeBV6d42G(L#VW2UdW_-F
L@-26,340II>86\EDWaR#/,7^3c#Z(#S@@R(B_/+J9F-A<+^50ZJVb&D.fg6d4PA
JKJADOF:V]8EfeGg4-3e58M=UY97&+:1+LT3:BS9BPVN1Bf\&EOJ<7>&P^#3d4FY
c2>=NE=QeRH3Qc\W#/G+S/=R[TKV+LQ>:A5Qg1f_=79&b\L.FH0FQX#PER#Y?bd3
P?-.f0f]fE^1+Zc]7g3H4+dT_8\?)E)NX)ZJH?938RG@TA=(AGV+/RJQ:[#f-?dZ
PCe2IRF_Ce<ZJ(^#HGX#M\;CCG=5/O7\=9FFXO@gH5OEY)8_).eRD@;LNT?\K=MZ
<BS?BZ\\QPPU1MSX/R&H>8I[bD]9IZ0\13BF7[5UA79A6#5+P)4#933F62_Gg(<1
cb>d/T?H]dCQ.^5=1R4O(>.WB=;(&H9J57fc@1RT_I.A(SP@\,+1<3_N#89(;P:1
FP;KB>A#F/].79HDL3U^F(-8/PT-YgOeVMJK\_ab#^KVd&e(01I5VdS5G@3((#R&
KUEXN])SCZAKU8\.2QVPdb_Rd.bVPE^B0=CP<J@89PFYRJ7K>[3G@G;<,G=TYLH4
(S>Y#RJR@5_?8/2C:QeNQbM;3QF6TMG;T<IZJO0RP(Bb8MMddYJ3YC(,OIYQ[XVZ
CB5-\88V(?#a>47W.[QO[GI:c(K+L0#_Og47VI2KP]+1VeH#RJQ78/IYECNRaTVA
Y&,^A?(F&c1[OG9)];)S^bGJcGQA2A?LE9/V)Y9]M:S(HeH25@Y0fN[_2JRLV6+&
IU\OL4#?NE2:+NfC7P<E,7JVe[W&/=C4d]^I9E_F(5:P9STV,O2:d5HO[)U1g:GC
WbPHdBS+/I):7QIc>]^KC(Z^OZZcXSD\=#>T>_XF?MC^LDEZB^g#O/b-PX=(I2<Y
=8.U5UaXH:=2&HB3_SIL+bT#+FGUb+0]GH(H\1,#BWRUc0YIWc8J]\5\ZZb]HRW@
FGP/TfU)#LK6NILI5Ud#c-RF2K<5W+,=KD(BRALd>8_,e^^U51bD);(R0OS8&W:g
^a5PSDe0,EV:(4LSaR1=5^_V+I2>d)&0baV_8We.,RSS#f4#<U;e2]V?Q5R5LOSZ
JOP5YPVaf(_cK&?e/eA1K#:-7-OYf;M]gA/BcC\N07BX\?+[@O<>5B&fF_FGMRF<
R[4L>\IEe]^6ADg9Vc=L/^BK.1e5Ee^],L)4F,8FVRB#&BXaaNA_)UL-V6PP(8RL
PIEK5f2HEgE4EG+eeN/8+e>gTAe1C9aZDaeM7S;IeSQDR9FfA>6G1XW?Y]OS6Bb>
c7](?R>RT1QJ1HE<CbP/_E3T/:gPJD1G5cMQT0^V.YUOK-ZF;F+#2H\3MDeBGNI;
I+6VZ+Z67MfJ-9:BbQ\[@cUP#-6G_B38:Ca?Y7EIc1&)C]0=43NR=I9],&6Q]e>6
HLPDOZbXZ:/20Q)(J/NOf5Cdc3<Cf=JREL6X@8OCK]da]3=0@H)9[Ag,e-1a\=T7
gX&Eca+ZTND/e^>X<S&_9]GPX/ATZ:4P[W2+2BQB^d2C=^WLIBED:ZJWL1.3W)C;
C:#-BG..>:#XSWB^XRCbD3G1KAgX4?@[NPV)8OJD9]E[3W,-.B/]b^C@BR1G,;@O
@fXVMRW-3-C6Z)+AC2#R53WH:bcV.ZKP1Ye6EZ5O-G4P\K.?K,QF+dKaVTV_J:V8
U/KWBBg&/#X59.=Rb87IYP?/J;F2>DDN[9@>84FAU///U8C\0,U@(T)Y]=gAL+K?
fC;?H<#IW@7_cfW^D;+?KT-[;POQWeNNB>JU?)P=_L-fWaCYc:1^d6g\Q_1_,F8W
_@B^9SL,?CMSZQLGNbWg15;.;(I+a&eD<FHA8([KG#-87U?ZK;c;+a__&Yg9HBQ6
4E.eQe@X5N\K7E)SCXT[F._JUQd(5E-_b?=T)NTNU;6_U1T?F#&++OT9=><N@(MC
R&gGCD6d/2G>5KH(\C6#cIHbc[+BP/^\g[bI\>4(\VcEg&+#_:K>aS[[RSID#&/d
0Y])(V#7;B@(DC.-\49-G;e_[UZL_E57=9d&XGQQdNF/&9VM5#2FYQVQ\<,ff#GB
/<Y[=WL+f5D=T]NA/cK]QZ>]4OULcb.@3a,V8_1?N@,CX.f\>4Zag,T86+2H?85A
QeaNF\)LU\SKWIdbJ=LF8(M(0-NF_FX\<V;(]&ZTG[.dQ+2E>MF^TZB?MW2UfNCV
;C+TG(Oc\^1Kb1FQN&3:/AgC;]/Y>#T/QK[\MY]F#;JBJ3ZZ6eUW4)KK+b_Ue6_g
/8_Z)TW=@D.V-[A1==Ef]+RL+>ZKE4/WI6-3d&fB)6B#+B,\EVX8aZY#V(;)S2?A
0fT/)//d2ZXagXU_]?PA6^=NcJd]9@WP43/^Mf1J<E2KARc]_dJ38;A)=O]XUg<F
]6HNGE&Rd=-WSTBH_JPKaTe#XZ1RV)V3c3Ke@VR^@P2U:L;f-E;e\]E@Y\6I&DI^
eJ_2bE/E^MA28fEWX2[_[=WdfS(Q@I;I^:B<2J\_KKFCOTH?SG8D.,D#]U=cN4]Z
b]^QCd<@M;1W]DT2dU[B#/cA#[V]ag-)2Gg-WVK(&<JJc9GKXYR+DZ_ON0\U+1DR
bS+?QLDg76?f)_b(0K^NQ9b13XE#\7cgCRUdeVT1>cZ&K#1MT>D?V)M\^#Jg+V98
ga9XO^ZS.8K9O13ND)8#88F7EbPfeYEH@Z&eb4c,=FD_SeG6RPH_/4#<LK;]B#ZB
g7W9FCOTHI?[G>NL,^3:G&(9[GFH60WD#WZ8FQgF=Wa,VFJ7](RBAgeK#?Pe(+<g
8cQ63C:/^@+fM_E:1Q3FVC.#/5,;afeH2NDCfT:AM[R,IB,f(:3=gH6T)MCVZBM.
C_6GAG8\cML7TaX>>A#b3HV\A2=(59AS\A:KA.RM7YJ(UQ]8e2W_e/e=Ng.2>\]B
aS?U-)RPD_O.E>-NNNH5DMCK<M-=G=)BF.#TTFFV@GKJVQ_KJG@5_TLbN[W?0MAP
fZT9Z>?X7OAJ],Xbfa4HgV:H+YGSaS=LaJ].eSJA&ScTK82:G72_-_4D=F\.L0;]
a:AA66N5P6E_G_H?&MX?NEcfJd<&V@T;X9K&dUK3I1I_dI9N>2E@c4B,g2O,L8K4
WdBX-NMO>5<3UAZO3c4@.<8QWIZ)>HH=P?F0BFIOD=(A4Y.P@-.[XWD[0eGS780+
aXW=^)NGgG^J)J;50RR3[V)AVYc8K,VA.9?J?]ZRW00_G6^^)ZDCga@,S0X1A&J7
5/(dH^WT05dOJ9:&QQRL;UI=B,BWLT-c9[]8C,)+\f^E^?PZMcNDT@>WOE8/O_#2
R5Z:fJU^QL(Y\14@a=7UA7,\1@K^B=LWHR3R6MQ9PB<DRQdD^AB+1-#^C3^>V;&S
O<I]S2I5^=L#,A\N#C>LNSg9^Xa6)c(6&5PN8LZF47Cc]G1Z:1:N^G-W,#D<c(S]
,,&DQ814+>]9O]b#],YHV>L;5QMaU]FJ)<]L?W/ab(W<OOIVO0CC_)<5MEJ3]dJ?
=SHRF_&[N3I4aW1-e+E.@PTP-VJA)-U:?XS<(A4YBP3CN<aLE=8RC0ZVS_J97-cL
#_8;K+[1VaM.]??.\].<&=IbND8&L-(J&V)bbZb4gH073/dQ>1J:d&,/,M<D:>cL
:fRPUfDJT5eB2PgfUYGgG()B)U/RFHB+F2GV?JHD0C(X0WWbNYI<YM-<6IXX<5:3
&R>(E/C)Ca@VLdc^=e#9V_d7:9J0J>CJ&C.P0^35=MNC&Ec,S4OFeK#AX#E54S+4
ZOSONUOc+:KI(cO,U\U7NJU.IP0(;?W-A_54Z&FJ@Uf0=g,H+3&Id3^cY?1;.5P[
U4ePC8X3A\I6#B.aJSU;Zg=M.7S^VCU0U5>LHG,(O,&4)\+K:GJO[+OS.cPggU[^
#Z4P+W4b4A3^C^W-J7OM)@NFVKOU-/&6A)S/Y@FPA9Q@=:EC=T>gDd?-EYP^dE]M
DXS=N&B9RI]>ZR]HIZP:LX.aP9Z\.f@5>5R^.f14B590eUDa)\P39dSTI0>GM2H5
UWF_G;(G25]]E4ae;FS:gKYVF1OTCL6K42HMg1#DF5aeS9P8(fA4_C:U+cbK?.(&
d.B/#Dg[K64SeYCJ6FDf>LOH&;SGT5cZ#@gOVHE3bMBfJBAZRK)EbE/dE&]1U6PH
-&3b]B182e2Wf\BeD_RHACO8?.@N&3BS-Y7L0ZVU#Q@YZ7/?W]ACPN5B21A7YJW4
LGVR8<P@S^S/F?d^T;EE5DB^^.K_Q_^<.R;3\d-3:.?gb4:=e<W#4gY59S4XE-0Z
OFV#]X/.T1;e9d9^L=282O0C9X#NRY2ZfM1S4H>A0<-:<4@AO#B,VRNW9JAfI<@]
E1_@CSSU24:MdMYBWV:]W;V/ad=L\KQdR_a6;?[;g6Z0WQ;eSO\27PdET@98&^ba
g)e@#S#/+SSCR:.R)KU[Z@<+9F\08)D8?9]3Fe5FcQL(N+D]Mf_:.7]8TRD^S,#d
c@[M7WWEAK/&]PNX#?V4=:Q.&cWKXKJHQ?S+?2d^;ID?#W,g/>[_=B]8Q3]<,C-b
JF.6gOX&T3J\g;<>RUSNRAYC#bR]T;&#0_Z]M\&a9=CLE_(,>7>8:FS2NI&)+JGc
SOSeUCVV\.]F5#cfG>+ALH_[<D.15UF(]X,3],6454IW?->^LC2.4K^;_DaN@AeC
6]P4E75HO)NM+.\OZ4;#U]IUM9D)&&().d.9fI-GRU&GQ]E&(D;c]cF&Sg+YK\R,
O:OE_)11+^)PS]KP6WJ\F)eT3;&YR)#^XL;>e/dDSC-YO,;)eEbIdMN;M#Z?W>_X
U:<)c86+9B=/YB,&&FceA#VZMF1MIbXVSGYA@B]F)BCYCX,D&Z@CRGac[6EXE#]P
Z&EKS@D,6d3E]aYLTXDZ8&Z4e>FE/>IJGC;[[SUAYBSe@+OW_3aBb+,GI)<H#AbR
?SX<C0&+I:@Ecd,WGBR7f=Q36b]S>K@#6/aU/]VePAR:@E0gE0L46OK@WNfKH;G)
O_-J<CCN9CWRG9Y,/fMY>7BZ]8YS+BdIc_JKU^BT]9AQQVT.][WaG-H[)e=V\X(8
O3T]=X[S?YV;b(+RIg464\^C](222H;IB?YCDHKLJ02&S9d@2e_(feKdG,V.g3&:
QDL\HO](INZ,7C)9WYATd)KYL5T1g+U4AX<O?R</UNI=W_eL9/94:#8KN4SDQ.cZ
)gDL;gDKcd5,(LA7E8YeQ,g0,CJASTHC9g_RIXDT#2KGR(K(g3.LcN^R0PNB.9?K
6O7-_9I(JQ0EX08[EP[V+W(3E<c.ZG(^=1Q9=&f>OUAE?&4,aTR&8&4Pe0=8K/F)
9;=F.I6).(fX/[Q]X-_-EBGC1@.OBV)&0RU@OYEV9U)>N+T<gbPZ3TcEN3Zg[9\f
5gGID2&.7g=X81cJL@=A2aZ(_4,0(&WR9?IF>/G=TO_<=&X@ccQ,8/@,5YLO_4.\
C#=eKfG0(A6Ke>#]UR\&QeUaDU(5#e,:#.#d<\IaLZ[IU84McJ^T0f77Z/)=.U>9
>468O]DVBA5[B?gaD,#&CO],XE1[MRE#VIA+1#/0g[4T-H.:A8A8DD-I2I/-NG)Y
]U5Y-TdY?c560bEgVJ.]g]WQY=R+ZgJf?@;7,3YLR)B3-<#3T7R3Tba)/3bEb+P]
&R.]ec^0=1[8aU;3_(@UN@a43T8d4I+b?=D;??I?)b#</HLT=4;U0>7&a[>ZRdW.
AMF_17b>ROM,6\95BTcae\V(Nd]GWY[BQRdULMP<-AbgFV12S9E_8Z4U5&F/abT8
?\dSWA2;(2[F18ZLAAI85Q4Rgb:^^4+#S],F#^T[dBaTFZ7g]_J&1]5-W9D97Ccd
,W5WIA+>Ze_)=DEKH.-FfWdaI7MTcYO5,^C_IR28bQB/^bXG8bcc?H:.C;J(@28&
Sd0XB,P&U9;7[@BE?T3C_2<gX&AgcfL43AHJ0WcIIgQG>I]dT/OHOeU_)\1Ab.-E
=SAI?.aZ#_(9AL[FLCRZ8-cY5IN\B(Mg00Q(HJAVQ&J0:T?6Ld8>]0gb[EATcc>M
QNG&=<ce:5L,cP+DWRf:BS[b3;UEILUFfS[Ua+1+/^DX_=9\P&C1]E6=JcVQ5#fY
\>eU:YK>-2ESf&g(9Uf4]9\Ug,)KPI/XK<5B1:E2K3L9RNMPb?9S.)>2d+5a+;dW
PZ1)8LJ3=:B9NXQ::=(OSBP(ECPTRT]ZCN[)6JE2XY^.)#J@.AAf#TGaWB]C6X]2
?NXO1^EaDG:g9FHdJW)UF1b-CF8WZe9;=L>;];>8.1aSY83c5^@^F?,e+A;IIP9L
QA/C&&RM+c4AR,;.XT]9e,/N^<(Z]aXD[a8\M<4WZNO]YS&DWgWD_Y9KGPQ:6GE=
?-MD.HH;48LW6^&QT,H<c>_^D2#C4eOD;S=;c5)IFcFdLHD/K.a[+UbY+Y0HRJPD
<2Xd&H.(65Y0TM\T+R0^\L@,I-Y7A>1=RPb^<NZG4D)TL]5cG=eJNCKEO-f#4\\Y
B<AEX5S_1;I7IJ+T\@;0f+_-W.WYc)^J+4LKM56:W@gf.bgb&)U[(HQ<LHK6GU2;
VAKaba#KX;)N&(fgFH[e+XWeB&W1?.e.PRE.@?I(1HFd<@FWa-S[:Y0,E<KZ.?#D
3GL/5LURT@^fYYRTLf/\L:;:OW(cTgOAS63@-&;aSR/M_]?&(&H]-\C)2^_H.ePa
8IO>&.;=T8<O]PEY;(3/4\NQ=G)AD>R_U>E3YE:9S?-9V^PgA4;LV5EEJN4g;6f<
WOC\\B_5NeFAK(JC6R-F5&U(IU^HJ(ZF++dAJK5?R9;AP(b9@g)XN4VU3DaCY(a3
/B0c)&&=6J-H7D,FU:]\b?J=#>d)LgdX#0fb]d_K\9T@,#_bO>e0,X<\<8H^d9Re
BcAHd[E20H1^KcX74YJ&@K+#>)A:\b@_I<X@0LQXS5DTPgKTb&S(DA4:/-gNbgED
2Bf\>gR2gB13P:4be(TTYeJAFF.cXEZ6JZ,?XLgGDC]_:85S1RGF)AL=/6N1f?R]
d])L#dfLD^4d?/\f,]P^M#Y>Z=f[+6d6_-6LF/W>^75ANU]4DR,D?#_AL[_6.;2+
Pg@7;3;]TdX5Sb#U^(6_5XeM^g1=]JA<]M(_ce61G<[R6g=?O8._711O8>C.(0^g
cf9R<;f.P^a@Pg+\8CE2>FA^)=/<\fa&+ANb,d[H(EX&04[A[3aU>FASgK8d\,1N
a\2:Q/OAIZV/KX_21JN48(Z62OCXYY/RT<=8I7L+12bT-dEG8]bAQ_e[G:05-.GH
(,4K?KPG:=L:LH#R;Q,.d=bE8gd<HS;FPWL2&_YcHR<F^C3:#^14BG(/8<8>X)^L
eQBBP[&:J+cBWW#RYEaW=+AE4F=[D?DH-?PUY?R#X5;F\aOA&_CN74O+3BKAZ302
TIV3SYbB:eB]B^G[;\+>WJ5U1LAGS&-<)V6P=2A:,17QD3=R?8P?9E>=+.>+02Q/
[e5/0WfQE.,WFHE326ZA8Pa#E,7&\T_>-@gOK375E)/H.OP(=.FXb(ISO0e>fE6a
OeD=b5LY?F4,]9):1a3]dYE]/B6A(;3gbT&+88KYB?D@Ze(P[9aC25F--,Z[XWaP
fV_,1LJ-69]S50J9SB0bSa7>/O;2McK3\Vf&0cD+/R-E]^4+BF9B/-H:6c4NKZ/1
e6O6:G;AVBbK?-<b&L/V04NLT&dQdXED#<3+/I^I3#+XBR5d;P44=)G^3XCL2.Fc
P<]&V&UPVVC^))T@BNdHbB5Ib7[UDC:TJ-EY)3d^81WUc)A=+ZBe=e=gH9U0A]dW
L8+QE^Kbe[8)NA.1:7KWeS_Y#TOg?4&e-N5aFO1U&AD3NDLd/-/RZJ.c98LdM96P
d&fYQM3OZ=bB@.V?#;cbEee[VQQQY&T,b_a3FU4P:K4?M)3&AIBQLFAD/eG74J2#
62Fg6GW48.1]2+ZZ++b&g,bBaeI7Ig4GP1VB4)d2&4QD9J-J1J.H@fWN78W)B3Jd
&]3.4-9(9.8/&\G5f;g):+@9;/N8<._\g3?T4dH:=S((+;>F94VbWD_IX#^a6F^#
@48<H_\3bcXI&CfH5.V124L3PCYWDF_[e:52R&+?LPeF==B>]3DU1FF5J1f\;:]-
C:SW&0G8d0AB9&>FHbZ10NPRYdTc:>LDYMDP2CT:#TAKJ@6-C6CbVDE?K0dZ;PgS
7L&d:8\4]34PMB)L;=0)CDY/De:UPR,cQ+<SO;[3D8M\9G[(Z)?G46^B2ET<)9Z_
=4OJY>09aOaZTAM?Jb_<RBYL@#,3IL7<UBY/D-XLHTDTWZd<YQ8c^5S^::._<e0R
eg.e(ON:2FDWA(YO>(5_6AdfS#OJCU.HU=Z2,d&U8(@SG;&CZaPF=-(E=BDAMIe;
[>U@P#&>NZ)T5I)Y>4FE?QXS=1Xg\GZ4eJTBY/^4>Y49R2:A-QK7Q2K-G?X<Q:a&
[N2^AUX8I->8]C>&@<\:g2D(&IGc\:03fH4HF/IQ8;ATeQT;:^ZBPJ12B#gO_JD_
_eJQ,_[=.Ag8R<RF7I0#<@_/aLcH<GH@8bDR,?_-&=G@U1\/BM;)IE.#3F]5ERT/
5S>;,/&J-O:?Bb7IR&_,^:QUF/+@4/4.]WXAM-EW3=/C]W/bgP4S=<X(2d]:1VP=
BGbSV/<D)O[K-R9EdWAfEXDVWW@^TA-DL&EWIOaO@B>XCIY_C?8[\:bfVgf9)3EO
QNdO^BVU4bFY8M@TVTZP_<;O]P_#KBWPSFL^4BW8&aQ1DWWE9Y.DCV(;g<VfOLNR
2,YI#E28U]RQ]EAdG@5\9RBDLJ?>dM7A,T?FY&P2&QWC5SV^#0H>6H2:J_eTCGG#
=aa331PFZY4I9+9ZfXP6RY/g\[KI5WcZ2N0>#:PWcAX=1,78:QLUe.eL;<2UG_1S
7<9V4Z\9<dPR;3(5235O)L,<[&T0CG9f&1@,Ha@:5NGgR#.8#/ZaGd61<c_bg?eQ
VJJ\N:b>AOVJDHLHD4TV@AB,/FY9ZE[b14NKT-XS48JXGZZa5F=Ufd+I6IMB7,]1
#34dMTC;Ug5:NU15I:[(\c?E?eO_NY,P5,cdM8T#f,\R2I28\O,D=PVMaMJWO:U.
W_/MTXa]T#9/3&\1?G3.U4S[-R27C6a6)&RJ(_IY7PK)SUgd,6&2U8;)KGZD@8ET
JFM#TK+^_0(H][fY?KJ3H+&>R3.6gELU4?FdE4RKfcf&cFE4<\Q#;F_TaWJfR8GO
/F6+aN+\1gAN&/&<J^[R)-2@,PU2<?_EA?f]HVMGf762bVI>FOdQ973IK?^FZ-@f
7;f5KIYbN3]F4&g=Z;+K7@)4cMR<T5=964Tg+T/_[\DM@J82e>7RO<S4]FF?AW8>
C3eg?SFa_4B???[4HTWFZ:]4CVF3K\&d>/8a#JbZU4),XSD5>Z,+<6)]MfDEH#<4
9@^eH701@^1TM8FH&UBd8F0UM)69,;AGCf(^9<_QJTB&\:B7]gU2.G#BG,:CQ+>,
bW1,42M_+SZ/\\<^<1#NR6bBcVKO0_dG_YTD);(e(7C0NE<7AePA-f7;;94M5KcJ
BQeW83<[CCQId]f/]R6@NM^E4g)Zf)VRWe>(PE+1@3D4#O9bN6R+JdSbUV-H:=2U
\;;:OeHg9gG>TX+?+9ddX_G1EHRgP8VNDD(86bGb>W#S(Tg+IO4EW]K=B^5cc<JM
P\fL(_0-;U3TYa2LUD7X0e<6@ZdXH..XQ226-S.0)5gQd<M-G+P+@XC,8A+]Yd#d
H>0:=5:2a@=DeJWG4f3N^@]K36e-^K;.48e,Z#1[eZR16AgaLf8(>7;)?&-R^bQ#
F.YbZ]C8AQ]1Nf>]a5T2W.OKCZR@]86,1f;=&U:+:II;3Xd[YE:T9B,]9RSU?/#4
c]U](YT^AP]O8-L=;=T/HMS,P.\&<cCC?g27aO&8FL7ISDC?,RAWP&@Fbd/PaQUE
Z)Z>RY2I5.D+9/\49(6.IQX@8Q(?H)30LV&R5G:104^eB,M>,aFUY_4-G6^2,UdR
#M#d)Z[OGV.BEQKT0_62&A_Y^Yg7HN5Ea17JV_1P2,GJ@^Uc&;ce5D@9_,J\:E9_
W?D:\5N3a_@>+@\R.]e=N,:I=d\J0M6B:JE6]JcU6:.6H4Qd#M72BMN?AR-BK<0I
Q&,GYb<-&+3a[9>T\<e.[cZO24O[50>Sd-:PL=5a@?U\ADA<5X3J6(3CK(T8JJH3
?>U,@0>[UUH)&.6N?R[R#40e6S?dT=^JeW(3E3@CM.X+R/G3cXY7)A+8)@O<W&Q4
f[1,8S9a@Z>aE:bPXA;XMN^K4F45WM3E,:[(=If?@HgM4LPVf0c347PEa6<)Af&?
Y\eG)F(R9B\G#8?RT(ABd&X235@91&^OWcPXH\ACS)KRK(T^9U+Z;J[S?U8\\E,@
\CQ3A:;=9GgPV0;NHc:32()HFcfO:g;W-aZg5TCCAbL+)([63QX1P()Qd8YSBd,?
b5QKTeRR1[1[3]7820aXe6TVI@M>YSZ(YAR-g@1AP.DcEGT<GHNNZFJHLUFgY&(J
eAL/2f[5XJddd&S)&)g@FAZW0+AOeKRF-^B8UA-2^55)FTeJ5L(6,6?(;<;,D^[<
+?gK)7(Bg+NbR.@@QGZBb]SH?c+\UOJ5VU<@BCPQT-P7NBaLYU2,\K]K7_4P149X
O(5)Ka6/PMD1Q@9M^-,bA4&S_g0;UW+(6SCYYO.)M/&,5RH;[WO4,-\JH9#_RCaS
PL-:]g<D.K\+/=\IOHM9K-D]Tg7TW=JK7aO9PeL^&3#)/G#V__TVb@CJ^HegW-Vd
D5HCSf4cdF62?D1+E-b8@,<8JF./+\YYGJg^/<28#IGPJ1.MFe4-A/E6^.FQF^Ua
]ONF)&-19e._OB,WUON2RB6K@HM^Jc8=)<XWZ/7J15cMUP3&,bLN4AN:eS6&I?Y/
GaZZWB+[16=HLSgP5a(eS]c)4I,+F&HLS-T/_6I;5[fW)294>/AM:#c1#OX&O)gP
XR(WdV?@GS)QHc/AR8XEMX?MW0]\5_?5/I)d4CK\F3_&VA[32U<M0+?&OIEX)CR4
T;d[I(:4&B3A]gA.HNGLg4f,<59\@.^@Q.E(N@)PO>9;O\M8P)?>,4(L[RA<P;<e
bW]c8O]FY1>LU>d(Ob0,c8L1T:&2#2#V+c29aZD_4>;_ee]9J7>K.-R?Sd#N6d;T
@0E:b>6eVX&-#U.?KHBH0fT1/ZWQ:B@f\5MHB>GJ]fe&;D>c:/H3@A41c=5M)F+I
WT0Y0?\d-QOP:,8;d6QY?DUYPSfYL@_&&@W;1LM=fW@b&P#bO(]/CeEf_5A1@DE#
M)=F9,=?,G50Z1DND]a-8T3>3-,;GP=QRV1dB#W/]<A2(9V[&3Z6d+PCJ?e[[2QL
7P2bWKI+X&AQ([AgBdTWFPHJ;@RZ+_0SON^&T?/g,O3:0W[d(\YH8fg^+N8W+@+&
ZfbY]A@J-;)]73eI(F&-X9S[[-I-2=<7FT,;3UDEBa4^#aUFXaJ3a]E.>a^9=@;<
S]2E^.d<TT&?M#WUcdTCGT#R4g?HXT=C6WeZQ88F^e;(B;7BL&FXgVTM7(EH1/<#
&S=&RA7P#@ZMWVIa&.:?a^]4WDbc482Y8SEL+L=0)S)^=0OM=83Hd7_2D#)[Qgc4
4X5NeI-eIgR-HG<,X/\C6/P@J;+7.U;/Qc#V(.OM+XT6?^8LFHE+Y&Ab@a]H\Z5Z
R>]AKW2bVKYRN\LJPS(>aI-?EA;-^&cZ48R-EI#YB9\;V8/PbaBbH;Y:edTI/(fc
>>KI^-aS#fAQW.LURUeYRR[DQ3^,8>=Q:/F.K=S:7V;2g#3acISB@YPX@^^S239M
]efXc--QR2]CWIc._NdOIgAV_7GA@3c&5WJO_&M0Y-3YDXaFN?8DT&FQHUKeN1?/
&=Na2IaL>4XT#R;8B>8Xg98]TXEBXJIB+&RK+MEZ9Fc4;-E,M2c(.N/8TT4(LC.\
#2_F[C,DQWHHI]/.-;;>IHWEV)<J:&VX+J@?T=I#.AY4(<TCRTHWd\)bYd+eg>IH
d(H=<bG+BKZ6Td3@B<(,.Nf)-6>I.Zde[\UA&8.V]d.6;,G(RcWB^AKEP7bH0O8]
-a[g=\,>RR_gU0\YWed8+TA5.7&C4]K7cf+f:&EW<e=HgF-_#R?fDEfE;DIZdY&e
8KNOd1]QUS&.UF/FPFX/H):+2b@Z7SGWJ:1U1;,AYg[WVOLLKN#+K=D>+YgP8X&/
a7D.L^AV_5Z#6ZX_3SK&YOQQ-NdGf]cgF+gb?#ACOE[KFZb@H:&7d\_24;T]/UKC
:O[0_?f/9W].a95=\=#@@0-X9XW@F;S.3TP[(>AdW<=Ec\@SSQ.BDFH+f:022+W]
cU,4JDBFMYdc+gQ1),.b[La@CRdL)dRZ_3L>+dHTe4U2b->U+^ZE7C#FN04>ZEQQ
=f;U>LX1DcPgXN0:QdYV7-&3VE;&IATc^MB>=59b^.(0S:BIdQ@cTHgF&Ab+7]Fc
S7I_V1cHS58M6@Rg-]Ib-+36c=Q)c1+N9<D/\bb=:#DC1I;JN;.QXeG/?,-M3RMU
bS(7MLT:&\L.H:[5K8D<F^7bXa(FA4C4c-UV_F[:V5,M87\XD\KgUNc@YFFFC5_T
5)gA^[3fFDcVWW7O:P_f0R(:@_O?7.Q^LU_Q[7WDW8-CX9MY&U>.+TM&7Ee+M9LT
=c__+?Tg2^2B?7DD[[YI_CPI]/e?Bd_I45Wc472Y9_90YE_/43&B5bB.Z,TS+TT:
+CAMV=O;NY]DH7fY9TU(fa?T1baTbN+(>Z\3QWOSd1;YB8T(/bSfUNU#dEP(YKN0
/b:7,>=fb\]0V\7APc94(a+_,E=H^ZJ)/EfC6aMSR@J,,_94-&df>83cYLYgA:YV
F<6-02e.Q=30;78A-2AF2ASM146.(5^/N+=D8J8=?-7_DJ&;[e?,fSRd=QADO@.#
)dM4CM+=EeDG7\GXKFT\4CLd&PA,&VI>\X+>]AgP?]cBHG,gJaUefb>@b.^,)\+<
g+E]Ge[=:a5a5T#fI/6U>E7fQPW^8e[X2[[dG[+<K5M2>2OC(-.\cIA&E(^EP0;W
AF;EBZLVJ&924T#SX@bSO9(Tf@F@7X;FL4OL<+g.eb((G=MC1N6f;^bb=MFJQHeF
M)LZPX2UH8L&G-]G;+^QVD:[ZD&e9ZH8>^SENA/PVKB)N7.R^-K2MF4\#J;:2e_a
INSREY+G2,\6SY2g<.C:ULP)/_OK50e7+NaMU,491M=I8OH.6Y[:OY^8\@O>>?_:
[5Pb<a8GY\0L+_L8_V;1L>aG,;K@2;b5(?2c7fN(CH-<GLY+O/A+2X>GR[>Je<DB
N1M-.8XN[-]LHS)3-&Gc6/9e.S=Q6-DEB.8K-Q<R17g)[1[P@05EHCNA&3&\17OQ
a6aFU5;cP>&B3cQLRWeKgeF?+#Q5.W1(C#[<UTGCA@@&T&VAHeKQIaJJ+(]5\Ze#
#B)OTN\NQPe\6e>6DF2b[\AcU0]U<;GM^Ee>RgBecK@gP&VR=L__0/JN\RJ]<.L=
E>a^N0,_8[B0&YORa=&MEJ6BMACfeTR@_8eQZUPAI_LDF,V\c<2.aV]]78?-_<1<
.44c1,G@+_Z^@D4F2=Q_R-Gd.T:KO&R;6R+SDSKBg)/D[T[5.5N8\I<fUc0@2=S@
DEY[WFDdJ;C-?8fDH46f9C318DE;YG?FY^8MaUTcSe\Vb(XC/=adGZALA_/UbI0[
cU<+3V?K=H>HI_f;@J2&ZDb5d^G]O]SQ<0QCD\7F;J^YDGWf=]gKVIJN@2#71T:I
K^gf8?V5KD\Z)&7@2DUNF8T-Hb[XMX=?&C<8K>g2B)7VJd4Z1O-<dQ&N-bDISFJ^
^#^3X7WReJP--H;89#<E??>P[G>M/:f\OC;Z8)\A4N)+&5W=X==B6SW.)Rb\=XA#
#S#&eGc#_b&104>Bgf78K[CMP3_\M[IDK_7f6;AfOR_&f8PIY@IY[G0IWW+G_V:T
J@37USR_b91(HGK_45C4Y^,UIE2)@]RS]VfIdGNFb,\3Dgc]NU0)P&-S2Q:DWge:
2UW=[]E=aV=:6-&+D0O&O?1;4]=#Xg:3;)Q2.L_1_7;RQ]gT[2H90PVS,g<&)BK?
0,6R<WQRS,&@0W>EQ;]@8O;O\[:U>#X&C.1>&0+Vf09?aCM2CTW^N)/9TJC8(d1A
>80U<QWOL#-.W&=?D]A7/E@Q[I8LQ<(NFK^a0@8LP]OSg:FTN,gc\VR<_?7K=/^2
E;IAaNR^(&#67L+SJM,1g(Wd;4GM8R/_OP=ff+EP-DCAFd):QT&ed_.1WV)5e[UJ
2c,@Mg&ZK]g?ee.IBD;KT\LIgcLaYP-W9-8#E]LD=a<EF-;LD4L#CW^:+08-7-=\
-T8SX=3AX)22X4,0S#2d<@DIV7FYX0Bc/5N4PYJ4_8IR/#0XP2O9A(EQ/a9.MM>8
g:L?HEQ42^+S.Xd#e73UULTg&bVbSJBgQXGQBB),M1AF3aZ#dLdE/]M)e[;FIR2.
_HeZUAB5[f0B5=4Y;:VAA)^2<)XYF76&(-0XAX8JaNLW>Je<4YMX]B;+Ka&2GU=S
+-967IJZYTReKWaLAe=CM_BIW:Z]R1;CY?DYe\UQSaG=1adZY+?].#(Z8Je2V,)&
9f.7C49gIMB;/]a(W?f:b]#>Z5N+QK>Ye5Df?O/MD?FM_]HJ-2SMUb\OaJe]R(T(
;U8Wd=XD8N7.]^&ULCX4[#A6:=-NP9=VK+c?>/L2&\O7E<ZK,5<YdFJ2f,XP]Hb(
8ZF?ZU:0+K[WQ<B.(UaP&DH]>C>.LK2/d+a6B=7fO==A3?ZD<McEcT)c_\OXR/7S
1]Q6WN1&T0)H\Nb^DY^?I(QdE&L])EHM#S9BTWHA8)8BA&],gg1:f_I)<M2MV+?a
H\a?cT]7<2[e?X0D)1,+BR,5;]0GKW4D;H3e23MMSe/2/1Kb>8<^GJ(R1,@AfIM,
=BLR0CD.6/3U2?-c:5J:6]ZL5K#d0b,&_AV:6(J<JA=?IFT#)d.XY0\&=0QPIC2N
1N/)=MV3HNNf<M;]5Sc#dX#VCI-8YX=#,R]I#+-DHbCVG[84&Ya<Z4FK&=#XBGV3
=?6Sf_IWfJ]H]4;gcW3@>IT6DO^2N^?Q9KadfY7HI&JKCQW.+:LY@5agZU1_[R2f
5<7dFG<(=146?VNgIA-7g<bgGT(]57cW;(X_.]g)&:>(1L:1M3>TUCZL4a4RSK=7
B<c)A@ZT4/Q0BYA2(0;U;AaW67[EP>F@b?(1:M7gH6SF3<[,]9?T^@BF/R)(54&2
/828__.HKZcG^;[@G#K02ae@]J<)B?b34L2##;MF7\5UUHX\QE:JUGWPY+X4]eSa
IYOcb_fM64PGVOec<BW2&<R&7:9+I1XC.IbCR.VQA[?0H)8@gZd0)b?Uf6eBcF0S
Z^9-Cbe?-F7Fgg-.7dN+?N0NT.T=YND9Q?AbA<a?)E\R&]a8()7bg3@NXJ18CQJ?
/\;OSaQ8f+;\(W.Ad)#BBZ(d688gIIW4(gPF0?&7LgI7>\3V8,^_b(R0G31Z#eX?
H2Q)URNN&c/,^1Y4X,ZG\P&VHL,8&75A@A(],aE1EUX3YXgX_M7/4-0Y34D]Y.UK
^=2#K4b;7N@]6[1K5f.VcL\ZKa7g3g7Tg(0g>LQ2I#YTAY,03da=a>9C,9K#E#Q_
>4I2UT1gX6a3BBS<PGU_,K(T;JZg6A56@d[1e+gfbUd/FQ9Ub)fWOCDP99)dM8b1
_<ZeUX&BIW[#0bFA1UUDYP\)JAf7e;d.CN+:NG-P.(TBSedM3=,:((bHVRPYAdd\
F7aN-a#E1G.5,Sf&2ATB;aN?A8Vf1#PZ]GYZ[=ZP4c4bBY9PAWHXX>#J?MU5J(D(
EVZRTBEVaHLffA@1XYV>.9=Q6X7^H)e5A:U)<#:D@5Z)Z46:-/cg/c1=7:]=dIHf
>N4/QQH[9&SOZB>8Q:/cQ91/0eS94<2AB3G[X06W,<c]>[YL6XH+JQQ8183b466K
-f^1\#5<D+&+6@gX-89-_B(@>a?]b6-B>99F1bPG\:66@9abB&;<W/WJgE?;)aIP
=.;<IX)AEIL5SQ26La(9AUU@5A^1,H2VY_bSFCQ;V<?KFN5->UZ(CgTXDE(0_1Od
MVR&^LC8F1U<V(0H/ZD/9=e_a16gO\IX&<0)@YQT_FD?@+dFH\e1:CUKB0C>0RLC
e+?e7-F2/UN(V.26.;4eddL+7fEB#^4-LPU43([QC=b7+)QZW@f]5f6L;6I:A.=X
C9M8T54c>(MgYDRgTa7JREKbTM2SY:ZMB[fK2D)@gOPYAGM-g4XD0S?A44a^IT1\
YFEV7b)dO4C@Db,;R:>NFWc+LHP@MVEM&VH8daOc>@:.W;2C0ESf><d?WCB+)?:[
ZSb)/-]GfS_]PQF6<Z31&/LP\b,9B)#F.[^CP&0]@UQ7ba&QCWf0,M#QTg)-T(IY
FSBUZaOWbM:V;,JC+@0c)K0G8f@]CBI<>^QbO,c@=<PQD##?T,#8+OC?H8S9+0@=
9K-OW6a;dc1,4Z2I?QG<LLRZD#aXJ1=cGQCf;K>630.cBF:g-L7)B&fe.Q:6f3E_
^gAC5P9\\M<;053:8F@aLSF6c_^8=AVJ&NXJHdC3[--..)ZcGGI(/4D]QP&e:f57
LYca4&:cJ6eOZa+@g4@)SE:T0<F^;V:IX7VC1/&/VK8]60VLH<\GH2PD2)U(>Z2Q
RS0fFIUN[67LP,Cg&C^SZ,,4H]2.-;+J37b7W\77)g9?=bNb/S)6IBGcPH.1cbN:
dDZ??5We(@e>3LTV^.39?d5\7,>;]:;>:8WGBa/K^IGWGS1ZW?dI6V-YMY3<gO-_
6O^B<]U/A41BW;a<1RFNC4[L<N7RZSW6S+V(E&<&X1_;Y+-#AGcbg\9\DR@@E;]]
@FS0VI7Y1=6CS3b8:4.c(R4]95E7H+05^_BZ9\T_QF-ELK;Z;U8[bW;]VE(K;cPW
g3;+VKWGg1\R>Le><HJ0cZaK+NX?XCT>2[)]YQe+dH:1>AV-6@e/###Z0\(LDaC&
R<EP9]b6Q\XJP/US3bf6cbTc,CB189<LR7</N\f\[Z/:9.^M^;P=CF;UV]=9<R.0
,XSgfBWV_:Sf;-X&<V^9bWI?CSX@I]Ha4dZOZ\a,O=gE8Hg(OHOS:/95G(O+\[a4
[WfG:JBS,A.[ef(K6c9H+9,VL3]ZGV^MXBB9J7bARTHR9?#X22>7A09NDAU</ZHX
=Y0Y?BM,(J[YXFRggAbMCFf:>UWJg=]c1#S@P-]3aZK)\65cf[A#>(BC^@AY\bE3
^NE7K?5;]b.52\Z1SE6E+7EK)b?;-563g[5>5JSQC,^,0KXM0VZU@4AV1<X8)N[R
/eT18g4SBD/8M9:=O1<Cd3aBe/0[>#^E^GJgE_?.(RLc4OF.E&7f-@8J.b\-V=&.
L@YgJ<>cFa\5QC@3X2fC?#5]eg<Xb:YKFD5F(<]D(^d,5Z^e[3?gW?D?f5[:d.MN
e3[=d#K[BWPCJ:C,)e-F:FZ-7\d9ICf<;)Q-J2OSQ2Fc^LfZ+KE3:_5&QGQBQJTQ
fITLJ^+@_c+4BJ(>a>K@R]\LB>][0@[B,UL>JKK<RB:Z1dTV/c4cBE2B1\U,/7\.
(UX981M8=ZN08YSWc1aG+1B7&O?_4c.c3c_@:^#2gX6#aE9fT-dULU\c8#eJOJT4
Sb4b0S;&bRK2HYFG,dA3L\^_#3fH)eJYK)2<MbDDd+L)#G\J=LcXSgBEEC+IRDR8
5)fQ=dCN>dNRW7,4MSPgD<(:FX=GBA>N9fJ[@:Q=(_I,f.WQI,56@ZKfD7E/RLRW
,VP03cU>K2X+_]3X6gHZ)2L>E)N)/dH;2\Ug7E4THY/46PG6KNgE\WCBGLSa-?R&
eOdf+#R:W++JS(9aL<E2<&9K+6UCgJ(#bG4G&PJH6/NY9?dVAT=K+,KD^\[:O4?]
KDbV/&9c:DB4KgV+g[L=D41D-)BdWBC\M6T67&&N^]DVA5a7C7+TG(@_[g;(@R&f
T50,KdO^4/L30[P1#ccH@^+Wd+YZ;cQe\,OLK3GT=&.HH&O\[^]d-EAPfM=dfBRA
:Wg)Y:A87-e.ZHd(VIV#2H5_X@Rg.>^+g269-OA](Nec[R+#G@0.OL+FS1K@PaH,
M9MP#B?FA>;8c>Tf\6b-W_IX8B@P?ZU&2#b9F\?7)BEIV_b<TQd-]V\O^X<GTR/4
]SZgMMB(&NQVaAQ_&GTW#F6S\DPELd)dH4Cc[cA6\YC(H^3]BU#43BP\=YKeB7f?
FN<UYZ]CBM)[:6W\9fa5A3fH>8Qa]6(IRB2<NUD>X/YICY6I)DS(FFONgL,I:-@0
/X#2C@4Z471Z.[QEc9+(<4P>f@ZXPeg(d9T(g,[(YdeXfa>;<[C<IP5E4LS905WQ
3MMUDgZ@V)H;9gU+LWV1\GQJXX(W=X)0SO@7A)^9aM8)Q6f6F^MIA1AbdS(.U(S<
4G46EC-U2X/_]Z6&U>LL?g>0(2JSX,;^O5ObD+[/e1KT62U75c=6X70?1=fSe>3.
_PR2>[\)FM4fGGZ-2LV(dS?CWB4;.C1JE+^]4S&5S1AbR93Z<.e9;D=TWPP+Q<R/
caP:deR7L&>[RbNe:3GUMHd3Q5Yb2NS3^T6N]=@-V#ZMS52DLMcE3dW790<G?9&J
\2#T.b-BN#1/4K,gccC\0P;E72aVMDX4GHfE_<R&@[LDC/WTd,SZCaO0A^M4aCPC
0DZCL<IQXM<F(5Y(BdY<#TGK;/;&XfQe8CFA[QV.J=,V&=[<2>80L\_?=1TcD+&3
<6-Mf_.^=gSdO2]6L\K6G=O-=9G.P>R?R3+g/2Q<c+23](;05EU)+[S[QA3/T]B>
W0ERL3H-TNAAfQc7[7?V?S<P):e=#f,IB1HggLdScVJT/[-b@@^AQGN2a9PH@7G^
FSbPMY-T(e:U6#aeBB#JF_2KJ->::^Y?T+(KH_-]F#.S1)e3DBfBL0dTMTGg0S,G
Q/HP=);9-+_eE5[a]/6E@M3LC&6@/=?J3UO-R.1C/G?#TRUGR(-3]@>,a.M>2e>N
ZUC8OFK1/Q&LA^,#OJRY0PdRQcI;INRD6beWfF;_=4GNb3.)GK.D4N@7-<.J4#g)
.S<:U7\Q4T\G(M5(6L)SN+?ZJ^7+0,GO2M[[SgLR54aX&BLcP/L9Q7(5TE06D4(0
U0O)Y75RBQ7XG^6LW/VK)LU^:5>.,68M[1(12;Kd,2Rab.GfC>G]V>Kd.)=DZT?F
@+C:/;I:dL6gN:WG>Z=W5SA=B,<R?5-9,1?(7^W7IE]Lg4TEPPEg_D8^/aLWF,WB
FH@71NG-9d&+](YeGP7/:d#5dDYfS_2F_9T+2_#<]fB86(^^&X#_YU0bNJ[V&&5S
>,O7_P@a1:A6)bFCc.A29UV.[_\FfA0fS-=Z/@JJXd3=E;JY0UeWWe0cfaZ04?3E
cTW4-cY&/C.3<2Me=HQG95c,2U\c/><RcH,6C<MQD5K7+-^>:3g=Q0#@G12\/.[e
^/]\A&M)LEF6<U9LOSF>;DSP+@-+TX11=badB#[/^]+GG>5U-W8>@^GL^CfV.R;I
#BWB-[X1=ZHF846?4MM^8A;<8CD,=.GH0:DYSebcE)2OZER94[#RRNEO@e)CdVN6
.)XV#@EWA,5U0KD),_UKB\Q=ID\_8YOED:-3;@Y]/N_>9I\+SfO?Tb+IW9Z1U>CG
&0A7U(X+H:IMVQb9Gg5I/FXJ[VfF]VR[L?0+Y9\_Z\RAb7))#XW+U(16GfHY8gVS
R#THE#>TXcUEC<^>W.2)70bA),=2IO3@VRWQET76NQLBZWHN[NT1>M.Qc80)dD6b
628b+d:caB0Q:&TA8X-]<LGa5F7?KeOU46OSI-[ND_cE^e>2VA]fB.LN\;dNU3ba
.^=7)]7(e3aQSH]g1,SXa5I>GRN3Ug;6WYa>\,?T\BP?g<#&9b2,K<R(M=)D?<[g
.>:H\b)e+>7bgc@8&eN5,BH/I30_g^:fB5VdA\Ne+HfWDUR>Pb5(>ILQH7]KO<1X
=U_:4FaEQB\Y,XFgM,ZKUGb#KM@DDD\((UdZ7L.T9TFT2-UgeJ6C66]GAN-c[0.C
/fNfO)d:]f.Z6<<GSALUNBH?)^A)<3NVHX,b\JI6ag2LIQ,O;#E&+.SE.3T;Y[UY
1dB61.-dUcccU@A[5+B\#.C,>Y.=bE@a&#7D_JI==7F6;[/5(MLWO>F15eW+WCXJ
gc4eC8-0^J#0N@@L(8<_LdNZb\EJX;\T<ea,6<E>XadXa_Y,UDZ@?E_/W8=R9&D9
RAc9HKd#B-QUP7J)d?US[-.R(,UR)9(<^KN;,Z?#bNH?@]-[BAA?bD&[1\a,T<Ng
aZDA_g[/UGDJ9_:B-P>,AOM>7-Y03.D]O[QLQL,7S[gT_Y@-P^DC(77.D&FTV,O1
./3/WCQIQdOR9Y5VR<>:&Y;>8<e:bFH65?-S-7\4?2QaS63Zcd??_(#HVMDf0[>(
\<e2[/MGQ\EKNUJ8/8P8f\9&\bb)?B>9g1]61/T\K8Y[8c2AO0237+e&DH<U6^f:
fcJ[/C5T4eYA/B#NRT@?NCLM^U^eY88IFeaLL3YZD;ZEA0gV+\-7JVI8b0fMXfW:
MU<6J_7.O062SHFBS]N4,ZA[]gc\76ZMZfGPCd5TDWFT=,e,:Q[]RD]XcQ,G]fHO
LWa9,9@PGPddQ/T6bAS7.&bT_V#[aES4X>#Bc#f[+eN#+-Wf^2G]TGCA\b_834,#
26@/1Ee6gZC1T,RS/0S<C>;D3UQAMCbZK3ACFKYR92U;afb9RQ0gSaHN4b,d1^=L
eQ6MNM[27L.CC7HCPg9#_S+H4=;U\WEETef1BLc\2K55M\ZWW\?39:LAA61F3(3K
BSJ8,AS7Da:3/UHZHY@?1Z-I>PdTfA,^W^eW2,<F-XGQG9Le2DKG1V8(>97@P?YT
][Gb2XQ_O7cUJF<]eG-Db62b<IUPdf@HR-6e24T[dPTI<\C9]45+Q#LU,.c4<GD/
bL@e_05P7/V;A(]>O:]c?UM4DL1M26-AUNL#<VFZFZI/PMbg:Kf?>SWIN,aC]/_c
4BK7__5D;CgaeE72L_;LdNc#R)9XM<>:,31[_NS0_J-<.-?QTXDX+GW,XV0H67RD
LX7ef\7:>AaQNCWLLbAJ3U@0c_--]B=<4\LZE:<LQPWO+R)K8Y>bO:=S\cP6b)a@
O4Q.d[#M)E0_H_AH<\=H/;S9)\D<:DIa?2_&GS9?(d^I)8X,>Ca]]O7,<I-TDW3]
5R6<OWF4O&P)(4b55[&(CWT.VHEb^Qc2TO6WZBE7,G)K_TbB:fGaF-Gb3EfW1V77
RP?<BCIN2F-Z\BNI+SEY&UA&@.]GS]6g-,HSbAY_Wg_fNHY+_G9^UF>+&\fIK&U&
N#<CX3;gHMBgP8)(L)J9-+C1/SW:K4YfWK=HP(S:Y-eXa=>9#(Ce]E#1LU&LC>4]
2=RTMV0QBgH4fY.fd5([C7E(R#-R\<532B)6,Wbad1NV++N/VC1J5K&/=EJI)U]F
PMW[AX,Ba0bB@YFHADL60+>\=9&;W#(b0\Nc<TBFF/IH;I.SZU_T[S^>M^]BM6B\
dW?2(#+-.;@VROY=CDgeV.@:0;CWe\B4D<Y8]YWV],,U;:M3=SN7P=_10_UXOL@E
HdP4Se&Z&2[c6AQ@>>\&EDH/N;gOe_fN\^4e.Qf/8fFc.RNZQ2:@DaT<>ROC+9G)
8^cF#,XV0E_@1SS/]-a7GED<KfC:L5J#H?IP]D^5HZ0f]5YYO2,8#Fa:LE3P)Z/&
WM@<-DdT?]G?X=/c&/0d]dE5NWagP2U;<]R:.(=3G<1-LVFLN.QOOU)@bL\6P0+7
HYT,0UC&X@Gf8XG4+gd<O?;fQX1LP+c1,NA/)3D/M.V&7/)=:ZQ:&DKg=[+/[_GR
:?U,:@WWZWYH.>3gPa140)L<&/?b5c0VO6>>Lf.PgXMAg+E^aDbR41eY_448PgfQ
;\d<H>MJD&<_Iea6ZAO^]MO8OU]=/6H]E^QXE(\;dV7=UU:T;>&>DGD).,O<F+OA
4<0T4NUIQYcVda65T=B,fc\3)aSb2S,,CK13TEJ5PZ9ZS&<UY3CLT@-&6#WXc>bS
Jb[Wd.UF[fHKW,0-=35]g^O(QX)B_@cC.>4M<H(E_,;.HX2U@8?:5UPW)O2@5^CT
=6F0N(:\HM.9LY3Q\@KOCHf@]:<6\>HPPWg[TE5dG1SREHK]C0_EeSKI6U5T)OM_
A40PK5UGf7E)K>>N)+g>K<3J\ORPE4a[7\e[_f=4@.)NaBB=7+D.+TdPA@OT#g<)
dfU=L:60SJeCLO.I)Zg@ZQ)0OWc<W__=4#S.=P^bACXKL=CQa#f;_-4@Z::F+@^L
A6;?WU[P^:D[g?b2SBc7]4,8+.Vg1\f<<4AR&TK:C(_<XBUF=Vd[:2:GM#JDR^>A
V-bb3Y>@-_SbW=b1?O-/I-M_]</7+QKKHB;A>/8+[K#?eg:3YF_SgNM;f@G\5.e0
EPc#=_^;-<)<BD-1OX=T5,]ZN\))1]ANB=]TVc+=QM1g:eTbZJD&LPB\WdB:2eUd
)//UK:ff<#CN?O13<@SN.#c3;7WJbWYXH=7M2CBBCCCA#eW>NXI5:Wb#+(f5>XK?
N@[3>?dcR<30[ZXFE^RRO7ecH2Q=N:A_M_1C7/K<d)(+a;A;-UP[+>)1A2Z[&J9D
ec39B55bH&ROS3>V6?FFS+3JE4.]:./-(QR#I,0,IdP_-17ZH3NT#VH;?ea\]&][
VY_&Q[RPNTIb:>10Y\2N1]RZd2172)L9_@c9F5@9><TAI0]3A2GZDOaRYJe<O)F:
0G-ILdgSTN9PID7C3+#__HB(a-#\KX5PbMGNU4K]UR62]2EaI8MQCK;L+NAS;9&-
6FcRd_BOXR942(R_(acJL2A)VUg(;a:VEI.(I+B-W2Y=4:T]O1(=CCA5@L;(AbWE
c5XHDW,(R<U7D;BW62B61bP?B)K@Zee=F.W]c+0R[\RbG/JXfQ00W&8RT9T:SgQR
E^44:5FCN_K6)UA^ce_31d.(T1+.AK:71?CGN#K]@dHS\>CB#KJdSQ6[UOa_7@@b
b==/^-gV9-aK5&A(J.\@R;Z_<4AOc^V9@A/;-B<1(A5[[9@]S1M:E?7A:]<_]<DH
@C-OSP?4Nc+V:T[3,IM/HDQ^]Y<W;+,(gV[.\K9@<:1U25Wa)Y)/+e.<c=4<a35J
8E5F98ETDX&6P]93:dNKGN:GNcB]+N=JHQ=0NO,R-41a>>TXb74L4ZBXTOL\.E8M
O>c_.c4VP/Y.S-SbL0b4g84dA/9.MKdGHBIAO=\W_,+RdIJ90POBC(:=31<=:J36
PM>-fFRb@<Z/XL#1OOZJ>6X2YZ71P3IgW<df/^3;:S?=S[@6c[.AZBVXA1d9U+#O
OIH4d<1f6EMYUR3DQWR[.:e>aPS@Og16L1)ZC<TY]Dd^CIOd=(BaHaOYB&7^]ZC7
9L?<+,B(@J(0aS+QLYKHSAa-J(#7)4C6dYIPBT-^^NLM1Z>.3N5#?:\eD1>aR]a<
3?1ZZ#V2<07HGW&aOV=_D&W[8\)JWe6:b-8Z;PE^g060.e8EM3J5.-1>aVM^39B6
a/XS2+CVRV\D:2\3#C/&DOUNI6:GNV?5M3]<]^g1>5:B&<6_[U)86a8\[7]6b<>^
LgUfZUfC/B&Vc7d9=R\-1/55a_N-Bb9<6_1T(S.H;d5Scc+8>bBJ)TCd-7RMT0?A
<HU@gR)E=)9]c87@=I7RPW,gf.GdIGZK<3Dg64YAT./a6>X?5M\.gINgIb_@11F1
YV@+/89^VH#4X0@KZ;,U.9F<U,]&0;V^a.IU).\04P##ZD/3KJ+P:;K@Z#4\IF.B
L9G#\-KTeY(MG0<+QCFfK6Wf(UI0SDGL<H;cBg-GeO[U322OFd7=XQTdf\CIR7We
JS\feN3A/<CgR_g92\H_OT<;7R)-)aMEWX&1;B?^P_\LUN\YEE,.V[P/6W87W?=A
Y7M2+(I4]O&6F;&54f#d0aXfORNO8\HEad),,0T\\PKD0FGOW<c@0Z0UPGFUU_a7
6<O;B=+.LFEc0MYISAO1aWCK#UTO/,c[2YG^0ZL=V_E\67QHU1=Q2,7KEJI^6S4^
5SJ/8.K;B)0XP:I;Ja22eC^,AB0B#7T^Sc548cTD==d_FU0?(^S@(.gb##TG+3Z3
-\Md#8e9L3#77_W>LEY0]G3=)Vg@K2ONd>CHBa<MHIY##@&<PHZ)gKc<ZMQ;e+(D
;eI)BPXJPA[QLRf<Xc0S&6e#.Z2?#KgRH.#5F4eB17fLO:#41/E0A9=[/<,@AFb.
MIQRa3O0;PV&e@eUT^gY[?:1L)(410X^7O,,\?B42#7.CUFGZ>)1MF@)J)14:SXW
Fc@HESND@.C/[cA9,Y7[0MCJ.+E6b_U?V(1\25KSPG]gML>O6aTPT8H4LcC5:+@f
T2EN<bUd81X6G#eK,<\e2F</(MSBeb#)Ma+ABdCVB9SCBF0(8[FE63;VaJbeWLHC
f7AfXKG7E7U=(-13T)B&MZ/c@-@e(WY)&#5EIU-T>O_6X1D-MFBVDS8EXX7]CS-#
T:d2(H&_.g#cA>H0_/ZMR;5@WEB71LDSH><1[EQF)9[Y+4QHSDL7N1BSg._)(P@S
EaVGF7A82:48H,0I^Q(3d]GUdO]H9GM(YSB8<eJDY^R1;a8W]bc93K2D\:>UR,Na
XS+e=3caPG#NX@C5,4PgfOWI;R/GD5g)Tf1X1\B7BH[EfeWS3QZS8[F/@-(8Q:UV
9f&b1((AegA<T10N8PA^^F4KdFa]9].O4VLV1Db6E&5ONb6Mb>#XJa1XB0IeFAHL
29JF^JR\5gaagA,_-DLbU=VZ(HeJdJN_W#@XDQ0XFIVNRQ/S(;U&Wa[M<__U7gV1
@]c\E^V0R7QbQO@]=MUc.HKb7>f_8#f-Y?g7@9g<DV@1FP##Ce.J=_AR3<9KMe;#
Z24]C=0=&IF@1_VT>&He)L6?6B+76G3&[]VC-b4V\NX9(06AfW6S+IfG6U2<U=EI
JRZ=C6eaFGIQO+,TSTbea9Tdc1:NA+GGI5f#JZ2HKS.3&=?)/(6S,.V9:V9#ae1b
@4-N8<aB1JTVV5.#MS\F,E/:I=3#A03GKPEW9S72d:4HAcO3\H0dG2,RHKd.H0JO
Q+6A3]4:Z6#G^e9KY1COTV(e6DE-+a^:<afUcL42a]/C<9Ze7d[9BHBA3/(;YSc9
;]g311Z)<gc&ZeRDX,?KZcRL>+CPFI5I?&C?&OX[H_X(.T8(HSYNG^9@K0?L&beV
UEW>/@9ZGC:R7JQMNDSQZg5,74H12FFF7#f[L&JF1AMT;d>[+4_dU;NNO_M#++_D
ITdN@)Qag-Qe(--WS3&8ff&WM^LIV-#_5HI8X=K,G9+6(Na?4;E_1X0g3)6UegDH
IIQ^YaY[&b5cX9<>9:gXID5f>,V]4ZTD+LA&0<YTIXTD3f,P05:)-/EJT,7VEK:P
0?>-G@1(S@FQ,4UC=U]^Z6-18GJ\(X0H59>/R)]/H+U8PSNSJ7O4/U[>8H;6@J8]
SEMQ[2=EN0&6PE)>3#@(QT3VY=-<AQN;9X;:7=[<B7Cg(\>b,W>)U<?eEgY]\W@O
3^[2dT(4@1d]T-Pc:X?R(8-QD[If^VN.Y8V.NARD0f;AE:b6X^.@P93]/589E+Y#
F]6LZI@S5gAT,.7#XRRH7\YMFB]264MSRFXDaMJUCaS^3Ma6[A0KN1W_77_BHRd3
G]_OW78c@E_/OH^1I;5>/Eb]b;B,4=_Ee+aU@:6AINN6AK,P[S0dNFG<J<^REB\?
.[eE<@Qg-Og7e:7K,Sf(0.fgY&E^DfHg)QZL@39XA;[L5[4+.P@8M&d<@@D-P<_M
F1-]5)0CC;;M-([F\OLY3GCA34&.<_?eB0KMO\=T<A(J\[(BAe\0CL,/LI:<=CK3
<;6gM]d]Hc-<Tcf(g^#Q-X-^3J=_V4CDY<6Y8Y=Z67L&+.,@\(Z2.HcHJb1#e44N
ZTa]Lc^VIe#Fa,J.,@(Q+QGF]PAN9XJDLd7IIJNPeda?QN-/M(Ma,H^Z7>V[9b-L
U<+=-9(E<0Z6-MTNVB;)ZXEMe+()/O_VEXNK<b@8Pf=@3:eU\^(38b8+XYf\T=FR
39O.U<Z;Q&5E);YgHZJCRE(U?ZF[d3SP:_O/d-c7)FbJAWcFd5HHATJTe;ZUV#R=
;^fJD9CC[_6>)0JAR9IZ3O[GMF,]dIcF?S;:.Q3(?34=#CT37PRd_gd7?FG?:RdJ
C::QV@5N)/#UDG:)SP[3Z8E\PJgVQ</VVe1XU?Dgb=3W)9JS905[Tg71JQNSHc#T
S-5IHPd<Z3VB+8Za#[EQ.F_XW]N^X_53b?>Jf2ZNG@CV]Z+9/.3R0ge/5/_ZZ0)B
CP&Z.\QJ>R;58<)#Hg[TMHJ2=56J_<-M/))_a;<Tc:(:X2Uf0OYC_J.X?O&2@Ib3
O8MO(J@?(@0)H+7_/:SbI/EU25[ePc]/gDN5;O?RE^6I#2AJeJYQ(5UE7+bFE3H:
Y@I@Kb3TeKgX8RZJAO(J.HVH4DRTS;)5(SG?NKM+X&1dK3A[GGWMKf9(e)8_.TNR
;U@74FT4LP1a>8fVCE-b4dV4e]U\AA>9f8TJS4cdL[5Ed(^(Df1CH1K)PG>=<.E)
#)KBU8I/C\YB1,U>T@O@Q9E5?[AebEa7TfI@DF[cWR\]_O:9-#bT^:Z;cM8^fY_9
L</)K0RRFDAYL)HW-T8<dI4J#9L3_H2;C3edfS(KMN>Q;b4<Z1VR;B[/]_]@DK^A
\+())\NeaUg\AK0+]GPN,8L]BGg=D-J&WD4_02Y\a)AI,_Ed::E.>cEEYP&(Ff(&
C;ZX=H)b^@]bf\-5IWNNLK>A722D-)6a]<e2cfKHX\IeK[5MdX+X>5]b-_dT#acD
.Z0ee?L)06UNVVC)/?c-gQ4(A.VSF@/@Pbd5e<Y+E3S&G]@[.?,[DOW1JM8b@A^J
.8@>(#F:9EZd\e/<<2EB;8.3e?G>?dC[GVaMBad[fC^??:H.GB=L]7F#H=]^HYK(
O;8SGNM2,0IH3J9&0@[aRK9O(#-[(JBZY^:JLReF;0G5@9(ef(33)EJT501T\C4E
23,APXVC/W&b/]V&UcLR>K>.>U/2@Eb@;KJU?#X1G?.^FK;.3FC(O:c^\6,HN7fC
7CCOKOBD((GJJ2e/4C1,8Z&W3UA@eeFf5:@[OV+43(7;:Xa&/aYP=.L1,AAS6A9L
F1W9YDd^08&1U:<>.^Y^:cEU4VT4NDR]E#PO_A]91D:>D^5g-N:EWd0YcZe.TW6L
B8V4OPU_96D/H\dObIa9QeV;QbOaAP4Z;Vb>K2J>1H26<7(bb/?(?;RM72E#IHgE
=&HY>=N4^Ib-5ZF0E1L\.JURG#T9>>\[AWGS4;E1MA]O:DbdMHTO1.0-RcOQQQQ4
/EMJH&f(3VJ:)#4@C9GgCEL#OQIda?Kdd65<@)M>D08PFM.7_b_V])a9cWZ_3^aP
F.dd[cc>8L+<N[1[+H49Jf^>>99(e^6>G<(&LHXJ^]+G.dFDa2;Y]A>L?9R4.1_P
@8H;JDY(6@HF&/X9KeDg\\FDd.5V;M&dT_FLb(#@C35aCfZ@3D@&\L3#T.T62[3W
--L7^KEFJKI/C2A:)Kag1@HPS483B9B2-+Z.Q5L&7\ZES[Z2[@K/;T/a+G-/ZN(3
<PBI/8dBBD4[8V_.]]#[.:7cK-f,=-=bY&aCW9+?&=7>Z#,W:bD3K\4:.;\2>[f]
N9[7?5FSC+?f&3M,a@#F[;YD+4M[C(1-gJ,DgATIKDMSWV\:)&@RHY(5&RHH+5,U
)Gc>a,F0>EbdGZ-6KH7K@04K5:eeZK?YEI]DK+)^^\KI(A.&##gD.aH:WW@7\gdB
+b(_^X#/aWaPg([=.D@-GE8\:LPIU6cg>[5Q17V.&5:abA&/.P(gAU#>6S4>)2O_
c=O+5<1>0@:6fHQSW#(cWPb=3(Qa6:GS_f@@c]2^Q<b-E;9FM?b,I:2HdDa=L/Y]
7F]\>WNYCHCYfgIQW6G5+5)KE:5&D-P1#f,,G8R5L(\b=BUUDC(L.QP.:O(KV(4]
?<6^@HX0H,Y8H/W#]H(Ed=Z4@b(dX6W@MUIT\P=f(6;5:A@c-187ccc2^&acVA-5
>7/L<=)=<)7N[&+GTb5V.^->W_9bc?bOaX<>BW6WFDYN6K0fE04f^=56Yb.1&-If
Z.b1:3JM2LRO,9,@@VI@;FKALYO\(8?+?H.bEKF&-5gKg?;VKG/HZKUe[HE?=VU5
8K\THEW.7&VPH0&YeW0e:5HH[.@73dSQ<(7KOZ]3Y2DYK:)X:e-)W)>CEFGdcN6)
(]20W\S-g@d1/N(=J48\.Ce-<fHaM;.LB8F7L(,6H<Ua:Z^GR/T\]0^+4@?5;@V(
KF]1B2JS9G]G/SDadKD0/8e>MJKSW0M>2]1Q#]PM#Ba)M8V11)a2E/D)3NH(2163
bb1c.4g6d/_<A.2M7/.XPeSMD]X=8K19ZCP7fCfaT&@GgTNCT)fV5QR)^D)<cVAM
da8JV#2H,P-gWK4A1CdW)_5f_VTI#Q;Be<8(\G[Cd)ZV,=Y5@?8<777&O?fgB7KZ
:K?e5Ogc8d9dX8VCCUg;-;L_:QC[<E]KY_FcNG,8a;OA^2Ae-eBDI[&0E/@+]6XZ
@D^Wd]H1,PE\J13=.Q2=)dQ^g4PSX0TA)46],;ag&1IV/bYC(N0U-BfDJY>]N3CJ
FGQQD8I)B3?TL8KTB[^?0SZRK.&>FX23QRMLT@@PCcR(PB&08^\B7+K8#gCT>6#W
BVXD6ca(0a.P>(d+If=HX<3a(cG]>S\QfV^D7H\@=7FPVGA(&ee@(1L#B3-P[2\1
3KF\)2W3,(SP4gID]OPYEESR#H&]1O2FEJ]>:eQ>d/.H?W_9G28&8PCgA0HBX:QA
3c(A<)6),.GP\bHYJIe_>2579PRCfE,b)R7DH:,&__;CI);J2@dIBG:3bD8Mb:QP
5N.Ue,gV^-L#FZ>g:KN/K?O58:G:3eB-O^,)Z<bRV?.\b]96R-^CNECIWN[R=+RK
1ZI].c(4Xd\bOOTJ\R4C&Tc..A9:Z[OQP;4?G1JG0_:XD9)4D)9Q?YHDRX2eadQ7
GQ6(#\WHL@@=+a:g(R6=ES3BFUQg2e3X_N]CY7=?_2XSFYQ^g0eA>M1N1=Z;N>]I
,>dSb1Vb.e2PFE(1(^>#--2WE.(e(]HSJg=D;Q<;W:97;\6)3G+=8-eL1R7P4O1D
0gGO486c1aEKVUXe,&=B<_H//d-KY:@:E?S1YR:c40YON=?bH+;QUg)+U+d>SI=Y
=1,0_ERWS5(7J6b&fA\_MDVPMd)EO(cVM8cM;9ga2f:7aT#.5<5R&Y5E\/4RGS,9
[@T\=QZDIQ?[O,Z2(4^4#8eK+X#[3>R37ID3DQUKN:HV)f+UC.9?.(Ge8)gLI_FS
]dUTSVd1X(9d<^c9>P1?OTZ288#K.NMXd36J/\b[Hf(N.5^W#,WKP:/U4JY8b]QV
K5&W9F^&ZcQKeN+MON6]DJY>32baBeG2S/KFe-Pb8eP.JM#ENb06XKSaJLI&V3:_
#>1d34MTSGG1N#&KP+>7E0D9<^I_2O>fO0);EE@b4Mc=PF\4D<-V>LP^AS;TY.Z/
#9+U7^;CXO:_\];T1GG7]JI.D4JEP1:/,7A(#XGgV5BdC]G&57_6b6PNXI:2e^CU
T)NNQM4(?[D=H@e8OI7?Kc&L?1d/.4f&Q0\-FN&SJb+[EV3^CaX1=PQ7G;Y,O2FV
58\P+Z>;97AHPV5FO?)g7_>PLb;O]8+Fd^PZ2H(?.5[()-41?43R52)]5^N_(B#@
I+\\<GO[@_POYUQdfFc9Va-JQ\[KIDD-b,bZ>g)W7]LUAfaDZMZ>;FQfY@JM/.5_
IV\\D?fJKAD#.C&4RW@L<J>AF+3954</c8B@fLe8?:]TD,2GBTUaFF@>QdO0bCZS
STE;0W@8</PI<?/3SK<U<WB,[<a:P[(BWGgWI[R/9WC>QA\Db#Id)N#XB9M;WN)?
a(PI6;R[;UaCOQ20fE^W7b-fe\S4.VU-QfEW8A26E6W4N<F&13_MRXQS69&^][/]
BXNL&ed7/a6-_@XIS:3]Qg\dI^NR3Y(QD2?29YFJK?88702[BFU1,AG@e;HNbBQW
BS[A+=A[VZOG?)3D&+4)08&M4[Vc:Je]U\<B#.Z]>?g8+)_73K33L\4SfcG\7SP>
7UPFD&QUVgHfDg:-KUc+K>\a7LaT>R.T1?&MXAM#BPc2&3)?,/YC;XJ,6:1NL:/]
O^:R>^\VE&4?U@5S1g#&We+S7.>eM=V=g4]e<<4Y^Ta5fAY98X)S^2733H#UVgUc
5U6T#Z]_?aKY.PJ^g]Q][WZ&.]5-)96,dPFB,;AM\KBFH3&B[Pa^G,<?#c?1;2cT
8CT2I#g926UYAETR[Z/AXB6CO<_ZAdPLTXS9:1[EP=T1FUZ9a?@D(;H?S5fDTRRH
6DGFd-OWFC8:];S9MGa.aQ4_QFB/Q])=U9B<@0b(7dV@?H=NMDI+-TdV]g^MXG3F
+S@7GQ_QN9VW;=\d_/BKMB,HF6:cMF/W]JPb;\.L/H+cF86:-EKJ_G0-)Ac6UGH;
^RIbS-UVJMY:?SeO?;XB3UYc,?a75=GUdG&=ASLK.KL_=S,,g#G&0SL5c@??R&^]
g53#f&6RF:f;Z._bg<(YO&d3L^g16=K,/&:(NP5B1#..cKcR\^77#M>I:)3=:DD8
H+:798<</]dA)Wc5K#7BC2BV^0O\6bP-)CU7J6)[Jg_J^BI7QJf\,UML(e=g.>g=
efE6XfEJ45f?H.U>cH(@-S@_,2.[D3VJ/5MI6:&-M5064(H@,C&XI?)Q?a:K6Z37
bg?O&FaNIQ\0:Y22O#2.4K4]D_[I5>YCaBALBMbb3A/b-DeBLTUUG?S6QX,LF-ZH
1DH>/e&bP]gY(_+USZ(GK2>Je)0@4^J^aXO-3Z0M&LV1b5/Q6SE.2BW00@\g4-PL
^CAUM;D5W;HPQJ[aGAUGd#YC,7T&?#DIN&&eRPV7c9?KU4a^f/,,LDRF^C3^<EXN
1AVKRE)P](\GMV#SFUEW^A4^GdQSIUgF24=,Q,?FDV+-Q=:.VFTK<VW7MNOJOWI)
>)M),PC,#@XgIEPV^SdPGU<bcaa=fQBIUY\=\ER_\.5SY1\e?A^H:O-8,2PTPgE:
NXM+ZLNSI6O4JTP]QcY7c^LO<&^/3V,^Ia@-_Aa[HK@M_6D]QAObBeD_]cM<_X)<
g<=(;=82]c)4=)9[ZfO4LCYB,&d<K-(3V.SHY/)PWFX8g)KQ9NB&g@f/J3Lf_#K]
N[AL;U[;FK)2+=::Mb6Z^,5]b)]2J=cQAM#G-N\UG+:DPBB741fLB<?2,+K9/.CD
19b&]?PQ:<9(g7;@[cTG>[2e4f-[>VJ5;SD@?29WNK2S<-]A?J^WY9Od?QJJ#Q5H
_>Nf#EI1+50Z=K;BCJ@MXRE^N96aOHSF+NBWW\HS=/PT/&D&(M?2[K1K9NUQP063
G@Y<3b-#S2:TCX:=/WU[MVe.a7<W,,ddWE8NaP_Q@#P_a\XT9CG4;d@3fHV1IN-P
2P/<\a;(:;R)VXgD_?CJ>aIQ(cXUD9=If&Lg/4bP2;g4,N5)HgU5ZHJ-(7BS\CX-
6Y8_@ZFA.DRQ(D(T/cW@_^(W<9DA,HTb..f49?)SJ0)bV654N?-:_gP8EO0,4KOg
3Ie^5JbKDA_MJ?+(9#Gb6V8?EJL-ZR4V^H\VWQ(SVG^-NDFTU8\J99-a.C<Y:eN-
C:d=aDA?WKR1O\9Ba)5?)<1Vd[da=?.RAU7bMa7)#9?IV\0AVG/+7Y]ZZY/95AT)
QO=T/=2:N7GHBEJA/1L+&X3CI)VJODF&HBB<J:BG[VVADITWYE-eUd#<XWPRI<ZF
KA?NP;P6O2:@4FfaF5M<+f7.G37KULb^G+#f+<I1M<H_K0D6g&1fGdM\]V9AW5,Z
QY3CQCC)#R^\KE_1O6+QO(+=eAI2Ned5F;K>fK3A@S?;R(/-2+P\(2H\&5JGf4<H
Q.[0]HGWVZ:d3.WbMYMd^KN?gZR=3+Jg&Q+_YK&bNCFg.#;?ES=/b3T5K8^5Qde&
6L@/VLPC+Fe6<:[5Na6af/b)-4OaXeB2]K[U74JJ83E-=\g+<MXbKa]_J)+:=@C2
3e_4@>3QdJXcNR>&T^5T.aV31BQ)g1>R^ENVM.Z:G=b6EG6g9\8fUTE/?X:Vb@dB
61g+ZRFX160e17D,Db:JD)J@f1#G1ICT,c-MWE\U&Of-f&C?82M?>U2JD4_bJdZB
/[]aL)R++0?g[<6\[+KWDG[d..d>7M,&&S,BSW]:c8EZ^Xd7DFE3T8WI0[1Vg;Ya
4^56^DEZ@Z:;C6E23UTD#HARb.2FL^8+QE@&&)WHfPg61YJX=2MUQ4=-b:_I1c88
#F2^Q+dDbDNS,S=0W5YH_gVc0L\IGa,16a]@#7(@;0dK=aObBGWH)_Q/;TEQ6:NH
Z#WK1fR;P#Ee75a62??B@cd(47X6^,#/^BOI>eD&+U_.7-O^3+SRg//):=FUWQ>#
S<NaS,=GLcLOY>bV;efa_6ReE?e.8Ie8+[XbUUg?>,;I8dSKW=5R#^,P02/dR.TI
S>;JaG=.7>@F2VL\-ILBaFOFgV+6K/D[:6HRdD43M/aT7#^MSI:ALc]Jae17.LW?
J+SU]I0C,VcDaOMI;7T1.f?XLJ/.J)AfJR)H>L>:9W<dg\>5;0LEc2,L((;3@.?&
.WD0E1H>b?JDCR\Q30U@R,D[X.+884^3I:\<J:SbUW4CfWQIZJ)-GcBTZ#R5f@b#
2G;]e2L_66YELddYE6]f\@.TTKe:O.^Zd68ZDYL&;0^aF^cJ:5.^8GDW5_JdF=5:
-V)?4g/HOLYBOYHO0:7V36fJ0&HY>b4ECBZWb&H?fD55SdVANd=Ba/<bMf8@++Q(
^>LS5>FY/2A&_(fZDQ.e^P#/4U)I@EV1JMA,Xb3&d/B@0=2Cg)E2-14HVTG\gI5D
>V8O:H)AE\-.^FR/,=HH201g9Z&/LWLgMRTQ_F+I7>Y(fH6<[WANf-OJ6/N@ZFg.
[e,Ifa]/U#,a9&XZ^&Z6H3\?F3[@<XOC;IQZ.A4.,;.9I:b>;@V>>^Zgd&6gRN<#
GU<ZG&Fc9@Y-bSRbfN_:4e0M>^_@LG)JAfOH8.da#XIC;@._J._5XU;S:^8\-#0e
)aVE\8(^a2;K/EGDIP_\1]fU^5IQ&9dQ9_<dd1=3B.=OENVUE00ZfQ>Vf6TAF14T
Nd0[bP@S>bGQ<K20-CFP/V6NYW>gLM2Ef;9W_eX7&JJGgaZeHR4\Y6HdYUeC34,M
]]N(?:T5HA5FF2G?JGIHL+dP[gMUa[IL>>__9IHP=1Y9+)O6:Ig>e\&-5T=)V:Y?
)N3=cZ?-d):ZE26\#Ue)4Y6f?GbX21]66R4eG35G\E.=@AbT325OBaI3Z8K]09C0
M(L+XT+X;40a#5N((D6J?aZ+86=11SQfcf#TA)PL>AO=GH1,?9fcC3/c/M:&[Vb4
2W&=-Tb<,c[6=SXDcYFGH4e[EJ,V<KU9@B;/ZFTB:N-B]dH+,P+//:KI>HZB5:UP
/9BZ1M0;fd6^PUDT+/@6A9V801?MV.0<Z:?:3gC,?Td]<?>52T4)XODZ:FSScY&P
KgHMUPPTT32<J_Og=@<a3_QZQ6\87);1R^^:LfWf^T3[Z0Y)#T^=8:cP8Y+cR.)?
-_GA;Z0T(&E:DdP;DFCI#7GJUY@F?OV>_F+fgEW-7H3+d([.E7c<R2B/B7IH0\3L
B0_gG;U.3D?Td#FJUBeOc>7&9G=[P:)N_6QCW4R=T>2]Z)@b[>)7@Z:cW(5Lc()f
E@>8RTA\Pd?ZK0\((65B^B5.P0TF_-X>#MKOA7/]??N@7HdDcYIZWOM4Q[ZL)e3Q
B1BO>RDDI-H<DQOHWgbEE,f[NaP)]N:&)Xg1[=3_&OH=7g6f^>(b8ZKOUX1IMS^[
PW<YgQQB&b=:d_Vf50&C.J>1YLZgJWQH;062?]/6EFd7@d.1UAg-&9aTIQVGRa.=
D.QC8Q5g^_B-_HAg[K86(aC?]R8O(QaCZ8?Edf9WM]Q3=O,\8aO<N<0<caW)841H
Y5,+FR23B=OM@H1F)VVNK5@HZC97f?D/\YbWcZPbK5^;1?7?4\ba-Dg@A7^:g(_+
cKC8[9g/4#0(_0_UC5L2\P;>\UP_&]J_0bTC.:(ZbY]]<G<SXaVb1<ATg]3b2\?4
98e?Fg<EHHGgMd-F]+aS+AXGM/:bNb<R1&3TZU4E)XDK[,Oa[E5W05)-FL(fVA/e
5P1DPfF__g_EdTP[A1JVF>@V^--2aA[G+[f1GMRAb4C0WeA7#HWQO;3E[Q0cWfJY
:R=9TBO<aUOWfH@B85+VBDKYdD0)&^@YB;77=-2_26UASEP,L7[-f^3VRJN.JJeR
dO7SQZ8E)G(&[g#B(7TY5LE1a\M.F8IBVaTN:[\Y[/0FM2,5Q;-P.KGddaN4ISBU
Z8^=TgB&K9GJ@Qca2GGHB6Y)SR3)-DRZ0+I0DD]/Y[0bG(Ra]Y?0-CO5&;W:geJQ
U#f@@4FAMFP/[=P]4^21EJ6S-[-<A81&B(U5cP4OBM-UFa/M<D&VXY_B@Y,<E(0,
LS^[0EK?CI>IgeIa+9)Y6-/#U0)T4?,E\QK]W8)Z[C0874R?eYELBTHUHMNYg84B
N-P)JBJAfTJaU0HZ=D^Wf-6:#9Q=#=\E[P1^0FgV]:.2[Y(ASC-J8>YEeOS/7+We
B\>&:2[XXcPDO#:C]M^AIDX-S\4-@ME2V#(2I[QWZ)>66G^#M;0BD8))e+2Y,?.,
W9,\UMH@=cPJ+f8gNFLVX8FY;<Z^O+Z_60IJ?N?1E_E5BKT-\]g(SM<4-:dQ(P,A
N8L01;6HUQ=eNYO[eM6;Y.]CL41W^-9Bd=EJ</CAED2-RJ&/?4\+K<Jd+5R9Q.:J
SJI8##2fFG\CX6BJY2(2@UaZcE[+VBa^>9[=@.H6WY,P9^5GQ-&7\eN4PJc90c+(
860bS9ad8;PQ_FC1ZDH6;OE5?+<+S?1L?3WFYW_@UK(Qb[A(,SH<O?CQ==<H^U.=
C^0ZN-cb_.Z1]4R76RNgObbDgBJ;=\g/dUfeQ1e0#=J?RTJ:?0V-/a,(DM=DEG;c
40ZUN4Q,#8b>=Gf^d(T]=_\bD?5L0C0NI8Y8Md;^?&&;8;8,c/PEO+W[I37X((Od
O>Z&1.D\LEZ.6f#NIX1T:K5\:43&BHOQH,]g79&1ZQaVc1]IbWg8;Kfd29[K#+fg
A-,[RgOF=ZF;#X>&OB+\/HJCS06Z\Q-b5\,ISF\A=117K&OT0DIY9[?PTDVIgJUC
S69XIDJ/C7JOgJD7K0_,P_I^<B>LJXU5M2Be5:M[6P&d;dgTGI-HDdJ[W&-H&KZB
G^5SfPe@:ZSS;[U_P+-\J1,)7Y<4[N8I&7&5V=MdXIME\&5>W=[]Z;E6Q\JgJDc(
#N3^3Q4_(]JFFAfF<cF^IB-4@g4<LP.d06TRN\=7,GeV.KC2H8WNP]#HO+RT@^-G
HJ8</K;.4U\c+0ZW:G_UeBVGcD/I1H8fT)Y/JS5)KJ3[aJOY&YE&JTV)BdZ?GK[]
Z@NZK7A]N-,7dGDDcT7#fHeI:KJ-ddZT=PDO4Z#Q?&dF0I::>GJ_@d1OHSO5=)<.
UY&R31X2VK#^LO;M68(/abA,?BW2O&MA6HXYI+f?02Y^<?@PF2:RF_-_F=-E\>0J
@.=Z&A-Og)d7W0eLX=(\P)WY8JSBGI@02C_C4fVH-8d86)<00Qca=Y12OAS8(_Z9
,SX5LDCA)gZ7&a/&3aSaf:aFC]I6gV;W[M.dM#9+7X\#?(^UQ=FH/7B#Q6>d.<0#
-R32=C(R#4agc)IY07(TeF,R=AfDIWC@gDf?0.Z:NgY1Zd9YN6dL48\5GcQ7/eZ4
ITdd/8_(V-2)f[-LM-#)1WCQ^=\LS1Z@0&EOY@48\/MO6DE-eX&CM\JHF&WO<f:f
F8W+&)J4c?POH//aR7/MQ.f:E(#YFDFVe7-/MR+QDb,E9647(73#)))\K/SKE28O
.1VH874#.X9?J3=@:F\)FK2_6a\e<4S\L8:>+1F+KOR++)\a2eN&SY71L\][cUN>
RSFF@WTN347DLE([YNC3gc0fX35]O.O^87]DOCNJ]]G&cG.bM+([gNQWG0cC\cQZ
d_:3?d,;EG.;:Q(7])VXUM+fK#^83K:_efMP-WBNQ++]WH4/(&YBYO#):&c4)#,a
T)X0LM?]cP<7#UCVYQeb@ggEbGW1-g0a;[,9-[/_#5,_V6b5U66JPY=9F.UXW^fD
dSQ;A_YYaB37]GN.dDN0ULC=LSOcNZ)VQ7E38Y)P+1C/SU]CaH/;d,/NF#B3d<[I
7I-#^-7IcaZ[(IM6cgTAHb-@3)3]7aU8(?XSFb@99.2\AJcJ&AO5#URI=Q6E,+/;
@X:2:(6]cf)Y8>fWT?3H-g97/<-,19^YT_<#\1GG?[9=(,-;FcXQ&c6_&ID&(T/]
A\FMQHT4:f]?=F:DHBE,A^=WWMMHI/P6O4@K#K#3TP4KMW&G.H8V;@FT#1M\a\KX
SOJ82P1d-b;NU4(c-61V[30:\L8O@#^7_)R?7aPCH([Q]dW2S<3f5H8BW\[aG,5P
QG9DD>3-<OAcfW+:e51SH[7E:AT2=3?,_>(f>?bH<D?V^SZYgM0_PK.8JUfgRHY5
/I1B7+;S<3/NbD72Ka3PEY231AI\:.9R[H4BNcgMQ.NaE/dd<>/U[&(e)dXT.YHb
U_,^3g4_M5Q_-+Xg-O7(RcDN=(J\&6((5J)#b<]J0I)2EYXKWD_G;L4MW/>AC/;e
>O^)?9#0FP(ZcC(CCZZ\e?Ea6@OPBM=BXBT)L>KCfP3+LCPc->N^-2EN<7JS/[3.
GD^[LUGbG_3[ZHOKRM38b3.7eA64fFEM,[58MF8G.Jg.=TgY3[H^DIKdeHA1)e<R
;.af.R.WYR,_HC7+Q\GL9M\6K+L[S)2dR(0ELY.7LHR?g3/>^8aSDH7<Ia7&#Z-J
XDWH3<C7/3Cf@^/T<X+gJ(#9]eK=X3f5+7KL,^.]E+L,SP.561N/b,R<Z=VY[Uf@
U^;LGd]<GF.fPdF#f]+2:eC_=>DFAc#[3B8<@X&9ZNXd0K<[>\bE+=NP_(?@3/0]
)VM#UC_W@Z)WE&L[9Ha4Mb@9BLP<Q2HY9/@a>VH5QC)<aDUSe4O9S+H9dAQ?3>[S
g734dD6DCgTD+X[#V+XDfF3=8/Yfcb41PN:<YBfO8KcdKdPT6cQJU-KJ1EX/Q]2&
HK9Ld_QL?-N<[6.BRgFgG(/]P?8_Ea(QN-ac=WD1ad2[N;+^aW8\^Jf=G2DC2=a;
8N]&SIL@)74Q4Dd3._Df.\;dbV_PQ>&VfC^c0JKD&5a+16+5D=>-AKeg+398^1fg
SbFEI;=F(_N>33\UEY=&g+,Z;R;R<2W-OMfAI?PH+G#dW+A0HK[94Ge(g[WPPY[R
)K.b/)980<PZ6/#<5aO\(\6-5EQ-=LA86fZ6[);]4,#6D,6a&Yg9DGM&VGg:5Lc-
/dD-5Oc6UA(1G>d[<=J[]Wg+^1BebQ+V//abI5.V93g6T=K>=>4/NQNTR]-Xd?:4
#K)R<49+-:3#?,=P.0(9I]eQF(f1b#W_d;C=EA1&_)(+f#D@+,+:JX]5>:BBNX2S
<<QN4=AUF\g/SF^^[Z(F[Nge4N.0-8.9T+<ggMd?)_BB^[NeB^-(3M^6V235:0AZ
6D49^C6DUFU>3ZY(-S?cd]U9#fN.@I.=^F=>^Q2d6?Z(4_TEW21D4cU04?97LbZC
KAVdZ?WXVcT,DJZO336FC/eB<C8&Z6e?@-N6>baRWgIHV)<UD7;>W7\XfN>-DfJT
>A=fT5f=LG<E5-\<B)H,)+6AC@+_5_#IAMP?g01dHZT4)0[Z@O5KBc7_I?EH.<=4
fG\8@7\1E/SL>(VRa#,;1VUKa2cIU4aK+J20.A0<,D;?<7EXY_(?/G<GJH>e;2NL
HZ+83U)RBBC\Gd=WGTfJfe:0-T+M0\JR2Bff:5_IG1c)f4SC&O7VJ#</KH+\1>I[
Q+Vg=KKF9O(,THMf1<0g<cP)aPNOcWg4>)@TUE\cPMIQPO#cgeeWO1ZJLY9O2=_@
f>^Yf+&C>>I=>634Y)1fHH2#)cC,=1g@NBg1>g#2&U@UeJ7^Q3K^1,J\73g2[Aed
5/O=LQUW/HgO;R^<+=(.UI8dM;?^,BA;MZ?a#S-6IS8)AX-WD-3^<>TB0=V\/<7&
N9JFA>-1&:SS.H#[=/a8/CAIA6PTCLZKe9-,d5=6))PB2R[6(HcA<R24QbAK?FO(
(g9D)&3b/8<?:DAM[b\,0CR_afJML(d;DRV^c[cLK4QF^-Dg5[)K;)Xdc)#H#DB8
)aS9:^T9?dF7_eG@R1E15=^/+5Q/DRAbA=W,b8Q\1I<7ZaC:Q\RTa[/_K^S^&=NU
H0E@STGUGRF@GJ5d;Z<fY]QPe4a;IS;Q[eZP7:/\ceKDLR#QOJa;EM6)UU8b3+#Z
7Z)@M)_+b?SVa^M.@:/O?[J)>eH8(V97N@PU_MET9??]SZN9UVfX&f5KQZ4JV#6;
_Ic0_bgTc2]c]YFX/N9BQ9(@Eb9b&(gbO\;/a\THI-I9fY/b+N-fBDcU5F]M6,f8
WV@HaZe0?S2B;)(2(Ng@0;<4Jd@0?1E1-P2_/<<+#]3PEB):U:IT31CQZdICZ\G^
F7-I8H;4IWISAbYd(</,T]4I[&eDd&E2MS3MUfTeOJBJX_.9Z:(c/DK&<=[]70[4
fK>e),,VSc)RRB7(DB\,A?.:F<cMAD-G#>;>:_(T.Y#:48656GYK+8@==SEH[dSa
OfB?YX:DQS-a<e6/ZW<H_a:Uf+C48-@Y]H&:LSY?VL8@VCLcL/BQ5>U>W2Ud93Ld
TFdEXS#92dU^&,Ac5+cF;Y;AgPSR#;E=,8CBV#Z>ID]<W8Ya<^8M(YS[\_gNf)BM
?Fgf>X<A;;?d1@@bF3KAf()(A(J(ZaEO+2:77W7gRIRBQ2P(05>-2XJTKObB:;^g
2c9e>H)6e1aH8,cP]5WE@M.YY&<]12I:f7.Pe2:S8/?ELCYN:13gBe4@0HRB1CZ<
<;c-L\;]:8;a]?_V2K1AU[->0)1e.[#B,Rc3K)OC?.54PS2V1HIUg1DDFSU\]E>N
Te@=E<bAE;7QHRX([)@A?b:6RX==-b,N4I[,B+D61fMY&C;^SOg3@5KXLN.#TfCR
&Z,Ja[.,4W?U4A<-B(D<:7=,)1CE53MEW#PQ@c,:3JQ#DG3NaE+#T.XJa<RVCcP]
HL^X<bHYG:d[\VG:a/HgC+R]5D\H8>JKW_U-#\>;3O&[E[JM7].:fbO]N]04CbAO
0dDM3E.?@N57\^;c&.7+6V]dPN/O)\9R(/,)L&^<Q8YD9.I,8]g]Q<#cT)RB#4Z3
Fc[Vb_B0+01N_Mb6N->+.?/WE.WDZ\=8Y[YcLYC82JSA([9^#(1/ZAN66#cI),GO
W\0/YgKbW;FWYfFGO88)Y?Za5/<HKG/@5eS/YO]NYgX8E\75.0_NOQ+E&,]a8\R.
QX[M&<?->WSSAJd1^EVCJdF.Fc>=O.b/_?KbW<6K>&X1=CO@>4GDXS6<+>\/?9FI
Y1TUX7fb)\51dL3CM@(R:C8/RT[JRegAL(N6V/K9BWEOPe8A[(.TT//NYDIBOG<I
3T/2JUS1Z(4dT+00QD6VRfP(:8_=.Y^8X/\cQ_G6HV2(9(YY68Y]^.4BeT9#6RDF
;(YMM0-b2fBD,P[W,aN-_aJ(cA85-:&46bGeM9&1.GA:CZT_->_cD;X&V0.7_9G/
5[Oc;-G1IZ1=2I2S31&:D9\]5V9L6LMdK3JR7U<G,[Zc7VbgE@O(QefO_.[XA<;d
NQY<^,dJ#>=])JC-SRb#e3+,>#\JTRQRc\TOf?DAS2T+>/8Se9/U#eI[W\Pf./;1
H4EAWC0190&RI>1D6E/:..;HK^=L4Z&<EU#406B=[XQa4I55F:>aO^B=Z(.6[a3H
4>6eT<ORFc@GWSa(^0cd65DE6gCIJ:d=Y0N)Ka0?X6b20@V)V>XMQ5D:7012XD+0
fa>8JW,/T5<Y?W4L)YDL2cQDSE0SKB7FMN)A?ZKPF0=SbWA4BcX<6Xg\Ef5ZC:;N
A=Pc]LZB:3+LTU4&@J5eUg&+3C6#G@O^e0O2Z]Q@;ZNF_e8BW^P:_]39ff8+7f>-
eB_YO;>2W8Q#M0A3]7=+D)Uef_Y7dH.N?YPK_Y#RYR?Q>NU7IZGYWg]DVW,U36,b
BG=,;<b6X[(WY_MI0+XV>O[<cH;b\bJX]e?fE3&C6Y5-(/E<G1&;D2\#UVF79I3=
:>LREX4=0E4?C_CbPT2CKOF@?a@6eOOK?K4TH]5P@(#0D@<UZQ\(;IeP[d<??)84
Cf-gA.:9e:gVe8)=@C_bI\:)8KR54P[O56OFY&c>g8AQ2f/0MFgS(CV;a+5Q4B35
aUPa=;b67)cRB(CU/(PcbcU<MQL0+0;g5BB8I7-VD-\&=R:C&,ODUJTLW#(Z8#c^
WFHLIe7SO7I6:[I+V:L0=E5Y?@RZGC6B9M,(6c_.&@-C,7>):c?XGMVaLK(D45IH
G<Ee7.B7XAC?T2b2/@#=V1OaFbL-+L]VDG1D;bFPIfZTdSB&;[#PP32<IVaZbDZL
Ia4<+_34M?OYEB>\gVb2+9FU0b:9HE39&Iee8A.EIc4@6^ba]Kf+3.YGYZ#@c<+#
LZ>B6]38:8_VR9?@U:eY6=X(0IbII2UNfZV2EU]^MgH0-#VRHc(.Ca:U;TS=>#B.
MOB7ge@a2=bU-.66&<EUXROPMH10:A[GE9Q8M@:3-D-f25&GWTN<]7aKPfU@&(GG
F^WQDXPN.^MJG@)0\L&<^O9K+66U9-.T2-eecL.,(GHV>ABf>Ze];5g:cO3\#dV6
=FBN46?+e0+1e+6))I8:NH71[.:-Y9GbHOB3:155Z[?CBD4,PH6YE74FG_(44NbI
#I<+L30_TJN<T?N_>5QS6/WJK;K=#Y.TO6H0ER^8-JSV+V8McCC/@cMDbcZ>cYTB
;C/(@H9B.]J>d?=^_WPcg\B_BE69[\40L,)c82O9eKJX5O1)&TBY/.bFAQ3C76??
_0eR2)L:5)50L^ZFU7Mc=6=#G)IIPVQKP5MVS_Y:2324V<NK/LZBTF?_9^6ObGBU
-TBQS:Y4W&K/)]8#0=,G[f9cMU_->]-e:ZG&fY5J,(9][V[8Tb1U#GF8c7dS8[a_
Rb#;&cB:-PR8R>VZf,6_D_V_VJJdM^/,I[gKUJ(&<2PELP<L8O+T)e2?KY?0I7,.
DKJ7DU(RA?78JXOPgSK2E>5H]S#d=L_^OfC6CgK&CF4T_V:f,(+97W8,/(V8ISe]
<F[H];6a2.50D3dIB1;FdQZCX-LIbZ2PT2/&aJ8>JC>)ffOaP8;20BO,NB__f_EH
#[b+fT,A#)VN?bN5OPSAaR#U6#57dg09Z]J>K<,2AE>R.\S#^a?2JWOc<(f[/#PY
Fc.=)UB5BCNC1:eBJVD-\,TAN2Sdd@YdN:A&+7<:&Fcb9[)+IGNHYZ6.S&FA-(_M
1ESP[Z&:b,IcJb3[O:#Y>@?CIJg9<7c4c0-1f[Ua1&9OR6g^JPJK(AGF#0=7&e#8
F\4(Y(3BIKF&;bW=D_IC#d85g_bDU[][A:)?E>U^ea/+e(4>gIG\?0YJR@ML.N>7
[^_KM7T/SNR,>G3QfJP@_(C/1\1RSQW8B=+b(bSKQF-_V5L3O>5SVV\_F(\VAHRJ
+J:XBcXJWET:1AQT091+5/W^+J1KSIRYDFE,6>?V0@&@=c#Te@BCJd(JZ+Q84ZX]
e)A3^6>ZQE)W>.d7@2SQbU8FGdPONDB[=5#11]]MB+-R&^[7^=W-8OcWH5eaUE.F
\BF\H/4L@g>HA3M)IAQHX7//_aIBV=(IS@9-R(X<XR7g#6LR0\fDTQIA?I#KM[f^
,8&2-Z=<B#H[2Ve(AOg8XIZR,;dMA,SJABB:+1;D>(>1/8WO>A@)^+;?)cIT#>FV
If.I[W,1.]OEQ^G11)3Y5H#cRMY4TJSM?Z(S6e.?T6NT=0_K:fVa(CcN^&:+BO2a
VeE9;VS>]?g/T-A?8cb#5W,R:[e^CBL2C[=A80FC;9P\7Z)fT&Z6GB-e^KK\@-aQ
L6ZDbY?c503YeSZgY;)U#;^-H[=8I@Le@Q+D:JI17-HNf99A0UF@;?=[J&X5CHG2
=a86Ja_A)KM/7IM0^DKQWaVTWVdeS)^]U.??gXeWT\OOV-FHeAa9\A)YK+93EZFb
ff8e1.b&B:HRT/U>.FW5fdK)bZJG6>cT@36/DM<1,DOJO\AD\cRgWP]:B<Sd@c>R
2OO][J2]:J10_^09MTUS:.Gce2+eNHafS>)LW75CH\/HT3gdA,\WZ1Ea>&=&.C6e
M^->E_bKQNF5[ZE>FLH@3F(P2?A;9B4>8c7O;GcH]GN_;4&<CI@c[<+HSS@MI&)T
UV=>)B7#1K_dI7@TR[]7BgDZ(IA.#f]ZIEGf+H9\/S\#8QO-&YG9?4653d(DDNeg
B(JV\08f019,X]<)/bBF&b9[TWC</SJA]<J_)f_L6ZUg]ICee>)KMT>H1;c[KF8E
5@H+D)]-;#&R<O0ZEbYD+C]=&-W(fJ>P0YIb/A_TccIPC+^93_)X4CE+aTg:(VY+
]JcJ-@EM\Pg[;9M&H)./W)DEb6XWG<JFN[937Qg1:<@fA[4eT9^E9UES.0Y,M/SN
>gG(Ad42Sd,:OYFB_A86[acX>YL=3M#DR>HfE0B]NV8(E,0BJ,Q?\Ca.K_A4g9O1
=[<Y,YQG/UMIO?HF&bFGYP=\4WFHE^Q:0(b;U)R<N+-#Kf@(_&[caYECLN5GN6.G
U>J9GX=RTA.a?>F8cfXGI?CY-^+1)N]F8aeNDUG5J_B((Z4:3C<eNFf5M>=#^N97
S6C&V8F31Y66DVQ(R(NDQ=LX?I_KC&J?;e8bDZ6B^_1J9C1A)Z/IKX#SOb09C:ba
7g@/e2MUB;:_e-.d\DA-,WT6-W_@V#/(I9K)KD\[GQ<1f#eg/Y3:#\QCQQ.#:NVV
X#P([[cOe,YgH).YVH:M-+148bANV9AJRd6Pge9)Ha[WQ[I-C<gCBTG/K:>]WV\6
=H<1f)G(&8e@RBD:0QYObW\;UI/RT<175S:.@?W66E-H\g_/>(g:fY61OV<VC4#[
]81BKK&VJ(A=XLZd=I?C#H^.E<.<M&-VT7M9EVQH.aQabN].^NF.0L_Y+X=M+VE+
151>]VZ8,Z26<.^VT77/P0.;<D6A5.@7R4KSUJ+U-X,9fYNV6F;7BCXN<_WFNLXb
JMa?PC,RgBaLR\/6E:@OT\B5=1SYUG;aMKg5Ud^M+R3?C)7Y=U#<K>1#W6=-7,8^
;:.QF4?HRP)E<1=1-T0Ae>IKA5G0<?\1EfF=24?/+_/gPOEA]+LN<Xc78A2dNY].
4Vf.L4T.:X2=gFNF??<JJGd^3B#9H\AbT2eg8&A6@bC9RUE@c)6S;._B48^<^bQ@
Ha2a&_J.XL;J@7#N1K<9\F&Y-.MaS1_D>gW5Ye.\X/81C.5H#Z^D^]14_E/T[5b\
)UI=,c/JFB\R84=2a7Q5P;X9S=LF13\8MAcL)E_0N1JAbAY2AT+4fQ1;@H/M:,1)
VH5]NQ)E0KDb4;.dA1TCL-@-\Ag43M)_&Hg:CC?^R4bKTK6,e:d&3-RILBV7=9JB
/T.g\.,(;Q@e@U\V#ECc7Ng=&^Bc^f6K,:8gM6AI+@7eVBP,X@K?S=@^Z<ZCBY]I
\2GfBJC)_-<cMT@+gWabVM1A1ROa92E]ZMJU,^Q.TRbJd0(Y&1QSIWQO78.#6^HX
(@IRL^Y0M[P8HR)39NG/B6ICeH_/Nb[.E\>3N+CX+;:3TT_e+]SFH..\V;7C0bD2
H90[-6EL<g)]aG4J4<[b@2U[)?>7agK1#-EF:JON.#fZ[/LK[Cf<S2D8@4U&J=3,
E;3+5RI8NLZM.0,]&0@RV>53].RAX;g9[Y57F=Z3Q+<,(4<07\60_J2JA/59WWGZ
4&N9(L[HNY/XN]:O:4^)+82GS98#?#Y^UR.AY7Y6K/O8KTA-B<M-\52AcP#0+B_E
+F\2bPEW?Y:+)Be\IW5?Q(I7LgcaIENC>30Q.Q4STUEg;XO7JT8-b1-=;L;)3:A:
eSWNW)\-bddX3(=I1MS@D9K&F6(LdFIO]5W:MLI,a4B^=2J+Q#d1>N@-Cb)KEBbS
Z^-\N_GJPV9dPX@P0ZW\I(a9F9=(RY>;8XRUI@S)SHCN(c=4;cO)[gWAKe=EOPX&
WFY\>W]G8UZOIOMd/GS#Ud1;-e(@99SKg)/5NMU&De9?c\P#NE])Ra:X.PJ,N8;c
7E7(3RP[+#2#O)A6G_D-d0AANJ:C41;?E@MgIZTT@&Z9geXKY92N[YZWO+YRac^V
GK5)N-+B:_a\,b>Ke2Be4;G=ff#7S[Z>2e/@a-FN+TU\()8L(XM^Xf=+TMD:FLcV
8F:T:LIDNO@9f5We(HW<:aO@2DW2aGP47a(8<F+Ng+CC)RISSO3NK#B0+A4#<dD7
+<A1_0)N60&GJF+B/BFJX+Ie(#E,0IbcfbUD(=cU9F3cW#F7aIT]1BC:BJ7dOd^4
M>KO2_40IWP-efc&QA]b-^K8T21OGM[<bc(a)EV=MG5CV82eV194H/(g>@Xb[;\X
Y6ND8QKA8#-)PRaV_.V=>deLL]<Z9(e+<#WRFLQ1XBAI7TQ_:=B#9\e6P.gMS>.4
/cC)KY2?(87^47TF/Q[ee2OI.Tcg2aR(Z\[9UJ/G</4f4DLX=P-#Fd@CN[T^Pb#2
>AZ5MZ#&<4A(]#N&9VXTSSXQ8F([8EBUX+^[g6_GATZ=^5RWLQ@d,FSL+]+^8(IW
N0G--I[LO_D0@88=bBR[>aSg<M8fC.0I=aP.BX6MQRF[(GT@S(0d9\Fbg9)4:PY_
1?8=+F<d6dDXd1a=Y4fcUYLMZgOF_E.&S4[Df90c\<(SSM?&CSXI_XMGWf=)N4fd
?;5C:We<T6WeQP@+D74:=f.K[>=&#6WHgaWLEBJ&LTgT>ffA#1^)-g4B=Me.E?:0
C:T^W:XVNL8KXPeCR;D3PTW8F[F4M4^P65E<<AYT)I;e@SOCH1Ca1B,4AO;:K?CX
I2KG8+\A<S^cM6/fK]JG(Z0YA\ASE]K1>:UG=?da;5EOTg?(YO6d7IEf-Mg3(PL>
Bf@41L085L,C]B_R&_:M^c@X8T@#g7N_O:A#,ZfBS&L#\9B:Hdcf[\XG<HNg6e<d
/1RHVXY@TYR;X#R#W=_RH^U,I]fADX]KCJDPQV21:PRE[9_2IUb9O#BC?^<:cWFW
Jc\8FYe&-d9eJ6eeNIe\aa:#^X/.FA9aY#D<7EEgT\8)(\Y-HOd+#a/UK^bK?K:Z
0E[AU[3>&OaZQ0gR1[_Qbd4A@OPLFeL:T:FcQN@9EgD@^/3DKa39aJLH&3VcO84W
ac:F:+NNS&7gJHBI+YB+PW6D]U?S@9/[0ZEdHSKaEU<XNL(AF>8PML@;GH0E6[^c
=FSJ\O)UW&W8K;E:A.^V;)ZCZ<5<:YATOYgITV./;C:2#;QCDX8Q,N8<OB/\1OTA
TON-@;cDc0f^=KNZ+dW>7L?>/\)>4>]P7:Deca3]D\@IOU4Hbgc5S;?Z2fZNR)U[
[-+W5UO/-/1d[;7AA_]8MR>OXD>BP:fdQ0[8BRE?L=b,cSO;?Pe;<UHHK,@,M^W8
I1M7K-3U;?,V[(QfU-QX^<U=ZIE;QaYVD5BXgRU9eaOF1V=ZIR_57g-)C=>aVU5f
>IS[XD(C=)8HAC=08SN\gRd:<CQ?/7/S0;0HM(Ea/LP>C2g7LX7#.:K8_&&G?I6G
937YP-?MX(PdC+(4Z#J,?:&E@Q@a&7Z]:^&\:)][+?HG+CT@_bJ?cQ-<?4E9[(Jd
[?W7S)^/I\>O-P&_\g]A2-^6SdP(MWF@^2c-<XZ]Qc9gHY36+81/;8Q9ZRDC7T^:
fgL)?^4d.\YQ([Zg:374dW28bTAH23)eaS39f;D52)SCDF3f9Qc[_3#[M/NO_fY5
I7_6GZ7DH0H[)LOg&B(V[N[gRefAfSZ4e4&(:6X8>FgKX0a:8YZOA]H&J4ZLH[af
[Qa,:BH/\YQ/SM6fdIO?]b6TU0Q:2T&[=T=(BP5#<)U9F+BW/XB:WO(3?fEC?:KC
R&e),7;N<?RG2,-e<CGB)GXN<1)RbMV9.=J(0GV8^B7AK8N7X9K1/J3#S_(,USJ[
K:OFFT2BbOLZZaVWD2cK6BM@,@VP=\3&AI5W[J@Kf+PO6Y_a2XNd<g_H8(7#YL3M
CSNT(O7@,_&NE=I53_E.EYecI4c75OKJ9JN\U\P56YL=GO?7BH)X/5WS=C_Kg8)(
5O+0C.WQU;/,=0f5aCWd@>U^:>9/B.49IQ514;^Dd4O(>J@V;e/>IKMbfcgW-H>G
eQ-S+R,#Q5c5?H\20<T>;TC0G(A7-(VC@_X1-S=?W+=#_>3R3U=(P^OG+[XU>9;^
a-^)YO0-d=YFA(KU:5O387IHN4_2?AWPAIe6YI_]JQSCRQXV0?BZfS(f]f7#1OdR
-FBJP:K-1cC.,cIXYf?=Re+)#]/c]/S:NRg2\e(^U07-J91-@Ha]4bKHb3;5WYB)
BU?dIHB>5P\.Cf586GY<<ER9R0Sf9/R^)YS2I)?GI5,9:8--^QL[Q4,Ge(db7Sa+
MI>PefKI_6>27TcbbAA>>:+F?CgG/<W,e3G.O5I<VE\&.F.R^gd[>1L_fQK.\T6b
XT[[S-cN\-8<e7E^LDee;<5F&F2\MI=Y6;+]2,Oadb\&FW9g@=\.,;JQ9dJfBWR6
VHMU2Jd[\/EL&R0W2KG?,_4O#W/C9eDND[/VV<+J=53e33[4<M:cgN4^I3f40-,\
N_T0LM1:F+]8YM[)V=<.RUS>9cgV7C=RFg6gD;ZI^f,@8\JaNW_</;4\R?LWDg(I
)OZ8;#O=Sc9(&EQ-E76?(G^PfE+]/YOgG&7gJCD@&_Q^E3W]\dBJ[#M6UFK,2C3Q
B(^Z_13WPe@\./N#X3LH:A=b8ES;^B6Y3Bd-\SC(^a795CA0&^?S]X<8H&^G3R_=
@W_)>W+Q:+\cCW7M@E916-#@].5Eb/:@1J^6S>Z<a9,Z^S=9TEaQ>;5U7-WY9FNg
H1E/^0(#OWJ&8ObfNWb_BdIX0UK+WEAFdPVBTZa-K)M@..g/6<c):<=ASBO)\e^Y
=UP0QXX^f7M?L&A.\+L7ffJT3BH7SQfMA439,2Bd)F15RNIX#[e(5CNTH_ZCM]@;
=A;6O=Aaf#&bYda0?HQ_7&7;+PZ;MUKM+BY/U3F0;MaU@9a&DR02eF5aJP&+V;VT
XT\O)d(U=U_KD.KV,]3K9I]QQ4@,c3GN)]Z=ab-)B17Db#QSGc-O?L&B_:B0D+?B
W^_3YAW+^c+8J?NZ^-9K_d/4RAA(eI7Y^-#]HbKKMbH;/B-A8M&MWfRV6aRb9b<-
g3R?A158&PR\?4\e4c\2)FFPB]<B)=.7Uf;V>>G0/LG8//_9&(F>@TZcdA(R1^^=
6O=2)d=_B(HCI]b37(5W6K(L0\6+e5;ca<cNQ0,+HU]&L<[^g2f+f]:RM^ND4_4Z
/H>NfXCXW]RNIDUC.B,H/KfU+fZLBI>2@^20]5VFDIcC2O0>JJPf>cTQ7W,>d96T
eIe[1W>c?Z2)fG:NL@8=25\@ZC7B-6Xf9K64M6ZP?V8Ldd+0])0;Q&,;&QB9=aB&
?2V6Y[Z9H/]30gA@J@a\4G=de(<IZcKbT?bBZMA8\5<LM1.>5G,@+HRNDfIJ(1J.
Cc^7PDOIVP5g,E]]Q0R3Zb\@9<[+KE(6^H=dXGbL&]e@OO6He4WI(NO.fFO9LO.1
);9YHQW+\OO)P80Tg5N3ON[JWIfb.Wb?W-e\XEQS[d=[6#<T5LU=a\E()8-=PVcD
ZH88JdZ4J_84e(@R^_NGDPR;)R)#D#U+=V>a_-WUP+J,0Wa6YF3)2IK@++Y^TA3I
#.;cSOD0D79Pd<,dE/.U,C9I3#11F0Bf5Wc5VE(200EG4K3__c>8VNG.CQddRH#6
IKINOPg<[Q).]AL?A>bKQQ==;_E^(cP@MT+GXAACL2DIY;>0dXVC3d[e?D\QYX6E
Y>fL>:-9YJf<=+&IBTe@b&V\c6><U:4[:/I(P51LKCOC^(2OAB_>#0@LeETgS]0>
Z7\63ICXX/[LGV?DR0-OTKb1K<K]PKS#IgB71dBdc0T]W0X7aHE\,F,c=I>f6983
F/aM467?04B@Sd5FRNGWdbW=6EKXOD+aQR@MD:ZH9<Lc(f9L5R6LDV28VW3L]Rf>
UAU;CRK:Z]:IX2Q+N+-aN@LT#ZReGJT#I1\S-aU^&@D?^HAg.N8FIQD46?c(>8#Z
QD<S)&\YFR7YV;1^;KYW#H@JK1O?2Q8EGN)bWHRU[E.2T,AdH<0#g-&[Y9#N[F7[
.C\@^;YJ\LT;-=R7.MEdeI4N6]VP-dEVca)1<WKABH,Pb@A&4Y6R/)#\/.AWLMc0
d_=GNfZUd:<^BM<BTIS9Y;J7T3VC5f53\DT<\(C;[-U2IJX?)F4P85PS2L[cdTB>
c:8a@+cQ\]+18V-WU1[:QOCOJ8;@egJU-.LO6^bGL3[VI[-VMH(LN\eE9K_+Y&cL
R?;Xc)12c-BbO/J+@7^c[+eTgc[/5ccJ5)^K9?A=XS/0P_U7WMd<Bf?b.&1dga:X
#c<)8DN@5AI[+O1-=f^cF+B:9>Z=;f=4:;d&]],57\1+I#&R.SWX(1@N-60-+3^<
;a1CW-DUQIERfgW(:[DaW-C>a_2AX2F[<G.X;;ZZP]=HLH0Jgf7=^-16-8H2[YLD
Mf+8c.6RXeM6Y/ca4(M3Z/A:\H1Gg@+1N?McZI1:-aMP=BGOf@MLF]95<_Z:Q9U?
]YD_eLDPT\2NF:;??e/3M(ZE13&9C8<0bBe<?G1^-b<?2^3M]dH5E,:@PI1ZC;BW
FAfFFb/TC&QMN,Q\cR9Q5U_A)A?c5AI30=D@:/Q/U__2)aA2</-XF&Lc+ZEfGQ<L
Z]O6_NQDa4JF5d<]-27P[NG,BbF^R>__N(e5C3C;Z[G9OH9GD3&VIUU)QZ4[Q.&/
U=]3&gY[Y@VNP_\caQP8=7PVLd<+;G;6SGLD&5L..[MegGF6&),;<3G#GXW)P@W/
58YcODP_#_UQ4;9fXJA]Wg7Y1^1862BKV1<04NDLf\4+H<F7V5f#bHZR)abKQ/]P
,-(R,S9E&X;NT@ed.9)3JU,:\Y60CZaVRa6#7)-dT(+(JPYbUdIQg#\>ME>g.9FS
R7dZGGbb6B30ZFC.2(-7e3AWI3dAR4-Q[0gPA^OIeM=1Ld-PM,1M7Q&=PG6Wc@]f
/PE^[3)7WUL\eNQbUcIVESagNL??YZ;YQCV-8)aJ]:M4O@9+(YQR13fEb>gE7O1=
QD[@S0^4;IB@4b4NbYcdYM)@[B7&YEcII5UTg>N.3_UFM8?N>cGbDMfK14;Hf_),
WSbKMA[;;<XgIcc(-.6LJU,#R<WX5WKI-^@Z;[(O+92X-R<(a<E=#Ec/1G6<9;8E
b.0WMGXI0U_4=,0)GXF^E4B+44O^adE8bOSML<beg)0<R4b+LO+I1;DB@:WeO#b5
KI9I)UdE0H8YCT3JY(42<;A/)Z=bDeHV@:=E),[0=T[^E/5:90RdPQH2V::MFE2+
^G&f@#Xb[^48^-Z?VPX&NYCOTOH#6><?Va1U&Y5(Sb.5__?[>gccL<:0.\F<WJ#E
[/A75GI21?&ABSK:JEW\/BLaBOfeN</G/fI8b1FH\eG6PVCSa7P/d;N=1QPE_MHK
N<@F=eSXJSQ\d(1K_&.N4.WPZW:3U3B99KOc3GfC0RQA[MV?1b.^gV91^N5ZBG/C
<LG-_5&^FW&?DZ4T1S=8RN_GEY-5_O/5(,+1?Z^\Y\WYGL/O-FdDF]<[F^Y-892Q
L1=Z/=2(1AXeB5dFGHI\PA/LQX6X0UW)P#T:@T+I32RM4,BW7g:8JTcdcDMA>.d,
&=PL^GcW8OMR4/_a[<=03Z3N?NRX_Rf8OFE6V/:\P6(AG;5PK\87J>KG[,&CWDD+
Hb7Qf_^KA(>eJcCUN43#;b_ZE9)=U-;502OC)W5=5]6c5FAVP0>.H[]O)K<cJCa<
[CRE6Z39+4058:-,VK[ffM/ffaf5^Z=TOBFZ3K?ea7NM,AN)Pd1<,dKM@cFcH+f?
\=#)B[+TOfT=AZZSd4X_&7F\K<N_)2SSa@Kg\8GE6U=MU6N1dIE^?3J1+QAP-fQP
gPVZ(Ug^I?8&-Z<N+2^N-E:E?0?M&gS^a[Ud7()TFSULHTK?2c)FQ=fKAISc5V)5
0.:[aS?Z_dafaa_R0Y7^K]Jc>FL^dT5=]//_YC]U::7]RdZf/A5(O66W3Y+BLL>,
H.Eg7BU5?Q/3,4geU5_V)]ffPc;>YET/Z8]-c4\S\?aU&>\X?a:bM,RQL_[fWRE^
B/9G3^>GPHY4?UaL.TPH;cN+5g4Sba2Z->>39OBbfIS4,+4>FF7Y;_XL2X:(cP#K
a+_[X&f3XIR#98EB<T0HAH#55#+?M?d)=]3OR5fM-=4#8UB^?#C?]XJgJXHa>+N/
X:0(2<U.+XH,:Z\IO][,]L084QC/W/?^/e7LgEW=3(S(^V_S3ZOJL.0T=9+:A3KH
=U+6Ig]8WBc4BC>\Af2e2>&CW\JQ+:Qd@;b<a)Q?#7g>QJ:=/(7AUBX&/7X=+@)=
MD\bg/?,LHgS:Z?\^.P-=B>bP=YLY#<.L1QfTcC(cJf8.5Gg1LFNQT@/RCS[.bUR
1,0V\ac9gG#_(Ug\5?-@18cR0W-Q0^CUd-?=7Z1IQbJN#cN/B8_J@@CPCLOTfcHG
S,:<ET]Z^\ZH]OObe69_GN29F&QO2>6F9_cP3T)E&PTEP]WB>HA;)>70U##FK/=E
E.1Y#B^=ZB1KbAa<+.=6f0K)-a-a5@:0<g2)==T/f[MQ/,4<<P[N/&T]SNSZ0H;b
PE6R)ZWY]\S1\T&@:SG+?A/c:cVF^BNF2SD;M5XF3@9<e[<;gEL[[[,:1<AMLY;[
NMZ,URVZTMGMe9Sff2a+F3J1,Z1RMEA(]Q:6g959J91T3?36bgT[??]g[-4DQc58
>LV^fdE\?A_1/\G@,Mc^Ka).ZF4?a?:3MAg&:04C<gJ_61USQHg>,gEN>)IGYTBX
cD@-OY<IW?W;)79;\9BO0?LH^1OVDZF#OR?g7+)&X\?LJXVcATJT:2=:?4LHM&7Z
N4C;<Q[9GD\IUJII.:KLJS_Y;[e8QUgZ9c9CAVTMAN(cfA-Oc815A53CHGR_>,\f
+I892-.Pc57g#L#8ELeB,104_;@a4TCfLG?+ZDORCSaegKEFK]D>?cBX56AJ3,#5
T[gK(GAKed@DOTJ+a]X=c#dQebN)D(&#,/A3\bJ4?_1G.[#a^1e82ZSE]>9e?UBV
E@5XRLHE4/d\V\A9_OE_8@E(3;?9PXH#_f6YASE4^H/<A14)f[3M)/b0@NEe@)S9
R=edMB?0.8[1FO>TK)NV--ODf4aV&eGU9V&f_1RS0A<XNd>)D^C?fEIQC=5T?V2b
1S,YAGa1],a<@OMZAAXR39+?J+?^_3).WDJbeZSg\9=BJJY/6G:g)1:X>1L#O100
;N.cb65MSXS93/_8)T?f5EWNaIPBQWS.:6e@6Q4(MT=b=aB^0#gG&-VA@-:5913\
R8a+g+[fRN-ELTFI.1Q.(3+K361.T(FSA),YeD<^3:Hea??I<?[&L(;(a[Id3BRL
f(Y71d/&7,@g/2(WBfTQ<J>IORH-C+7S3M<J<Cf1]-/4Z_FTFe)^3ULVLaVA]J0A
S9]C3ZKc-ea>@^+V9LX\_=Ve<NHEc:HPbaN/G0;.<6c1X;57(;>CK0e4[?F>A:10
=)cfGE^ORG[I.W(&c4JN@S)ZCePeS^T?;5Q;_d]a&DYeV3UFK:;V?@;835f\OZ/]
=0g)gb_R7F6ed:@B=QH574I?SXDNf<U1E((1BOL34F12/&9.dD?+(Z8[:WJM]TaP
L5@PVM7TfL-GT2P>f,ZE/T1GS5+;35<b--_1G(_N6e#JC&FAQ.1/:b-OYab42O4;
E=]QM_Fd/aNbXAZ)N2IF7RX(.KSG,20UL86VI(aTTT8Mf2EWF2)I-02:@NWG>09R
3c&,IfcPT_W[O^eE:Z3]aR:].+0C[5_Q)7_KQ2FS&+Y+.#=f,ce7R/9;TbN-eYYg
=02+VEfV=W:G/UV?b#6A<6/BP#^MR6gE&6_6;74d/>).G6R_XR9L[?)<D<6<b,aL
^b=-^)>g+:&25>HIPca#SCEX]HJ8AQ179UYR<@(HGUF/17R??U.?7H7EgM8ZUI<5
EPMb7EA.@>1RR)@-YX7M,G]J/6Vb:EgQ#+IA66;I/-&+9Y;+:2XV:QQV1(@Z0M5P
f)8Wd3YMS&ggEc)&a-Wd7X@6AcW&@(V&P7V3aS9M+B3&I[X/Fc55&Q8N#73NL1[=
E(#+5VPZgfBPVSHM:[2GX8W&^^R-,_7D)14PF(gLZBdC&=M>?d6>f6J88<8WY1M;
=EQSF[I@3S=ef+TF-gZ_<=#H.T=OW;g\G/TQRB;UUZPBCUIf3+89U2J<_S++;/cN
)WKM<]cMdH^I2.a8Z^WPZ>b=LJ0cRSBP4V8B:JBb)(/YfFabe1K_Z\[@R(YDG1^S
,=I+VC@c2O.H6-SBMN_a,_,9C#(C14C9H@Y&/]KLP.U4g0fQ]/^0NKL:\D3LQZ@f
)T-:=_\Na))[0C[dCgc;7UURDLN<QXgQ3)>8e5<VM.EEAaGS+BVL4MD?dYW8KNS1
YW)?/LY()&MfMe@V0G0SA8D\^gYN.L91V)D-#S,?L0UDGZ=g;d^P0F\2H6CX;140
I3_SL+B7GJ@+I9LIJLC-?_S@AdeZ5b01IN<Fa&UJ.5,gWK/<aEVJW,;He6/)3.IA
X.VF?b6)Y/Z7#G3WCF-[edRQ[RNA(_Q;R5DAfJU->gJE&HLX>0][eG#0#Zb^IR=V
):4V3DGL7UUbVJO\9V8A+b-WWa5_S19QD^E2+f^>3L5&Y&N06-K?36M:2<Xe5S7S
1^ab^D1F9MR;GW^8@XJbU&GZX#c)I]-UHF+Q=+@6_O[&08/B5UMd5GTO\\B#+@(4
ZPJ\XgW.PSeTHa_5J_AD:_.e95WRW<S8970+V&_DKYB;;5#Dd>f<;>-+Tc:(XW96
bB50O,221eNL8A(8,KJE2[?eC6b06G#:R9dP;F1W#fEN&)@Q?1IY(1F<,-S1JG[D
D.B-2#14YOKcWc;b)C1JO40d12XKHZ[5864HR.Vd-Ngg_)1PDZ)b^(F<CAc?G8Q#
Abc?@]W\:[4=g5R+O45VA+b&#N&F82?QK42aXA;dYIXJV+7E\@bPU2?A\683_c6K
P1J2cRbUXHa7:656g.1ZMLLBI83b++ZMVEX5,Hee65B\@+OW0+,6IAZ;V7#X]N)a
<B--JNO8^d?MX2_Zb8W&57-9TN.C:ba?X6aE?G5M\e:3T12LA17H9XZL5BK[\GUO
],bfAIXf8g.I+(A4&Y)E45QO1Z/d0/UJOFcfMKFG&^WLQC8]>O[CH7NPb1AUe#\P
d1JX]/\/S9a5b\&-,FaB,L@E:N/4YOGb(/K&[UUNb-N@FAD03ed0b#EWH]=?LQ#4
\6O@Wa[^V9;6cgN,-)X3]N1;W6)3MK:1+J>?WWS\7_bCW0d/Y.g&]H;1^;b_(6A^
).1;3GE)4JVa)>.D>@V/24fQ=46<[?M#<2]5WM9>:^+-^#Q>ELDIeR#Y#d:O=7,c
L_B@6J&FQ\c\Ia,#=#4f^1f:K5VT3[e+#c7g.aB##[4f+YB7SM]Xe]Nd@3+0IJ9N
S)4GENG6&M5285=<Q@SHC<LCF3fD[C,;P>;DW94S7>):ZL@fI\Q692I59()P:92[
&C.S)Y^AVfA\VVe]DI#0.(E0_JS#D>eM;Q^/[O3OIc\OOP.X0JI?bS=#9J=C[7F5
^&(H[6OM9A#=eQHE(3:TVB7#8cUCM_Tg&)_d85CFH0@P_=@:)#bBfPJ93QGc>3A=
5/aF+a/.Hd==-JS42@MC.:OcSO^+?KIgbH<E9VG9UAR0Y-\L.>Q10SR[O6YC?ca<
P))3I8ZCVaJ?KRCC/HKNc&5[>f@+W=)S6V:G?/aM,f-X:C8QQAK)F_T3+#6;_T)C
2+e,N=MM86CK>SCZf<R-GT7L:2&1Gc4ON1-&@&H0V4E[CI;^,(372eB9SNY]ZMMC
=5\AHfdM\TT1.;U8.92/U-eZd;5M2O?b</<cY/)=\3F7>X&/&,GUbY0O+I>-H4Q,
MgU?dQ9V76[\Y\<0J[a39U7U18(S2J@Y>;R:.U?YRPEP?,=21G6W66)TdbP]\>Y0
8Ze(ZH1(@3_M-\]=aR\RL&0bHBSEfLGO4d-HE>NZF(g]Nb2ECBPA;5G.:aX>2aI/
dANO[NC+d[/L=>I_I=F>L8;[?P0@H#+5F[S;K=HaNISeUTV5VYaM#PT?[C?0SD@]
X>SOF\4/gVHI;X75d5AJ)Xa@TV=CJOX:,Y<)(T.OKH?)R#7CO@a<TKR6NN/L@cIY
H9@W1c4JfKIKBG.gR]W@E(+6YbfBC6,P2]UfGa.ZF&,,[X>/dD<VWWS9GC_SBS].
P+X2/1QVda_+2V>g^L7)0QF4d\0dP^C>BKGW([OBU,WU;^<gU&f4GPP#2X=U/3aP
(gb23016R,3X?05W,Bb>DYK3aN7Bb+@3W?,JYFWD8EbK:KcXI-RUb/?=<d:]#,>S
dfGD:2MU488@K[IG5().5]HU,2,&IQ7N8<4>Q:G]Y^TO17GVF^QYC_UC=2;[3996
-;gD(b007+dHCLHOf?@Kd(-SZUc#=./S)=PfVN.1Mf3g?=SEOPWHJ+Tc#1?g]>J\
(V9Q@5SS#B/V3QEK/A=UA^E#EfdE>.(J]BbFeEGX1FR)0&=F5/\UZ8bF#[.+<?<Z
9W4T9.1b_C22\K]6VfQLJQ>/ga-<?,#a>,^4dO&1::[Ba(B^Pdb<:[YSeR3S6UA9
_<W.7O_G5IWd\1/^J\d^[[KQ;B;2gg\?:_S+OLZWZc6O6E208Sf^Ig_&bK+1MM1Y
8RU-^8AL&)VDU]1Q>4c=VOf(>f[8WS-M&9S1f.I0#T9GKD&ZGKe\OV^WN\N#.SH/
G=B(_Y5HRa]D&#:<OA<e32(d1&cc]D\3TT+K\ZS,/2,CN&I^4@)d+(W-4PPFL:2W
S8+bdF0.>GZ06.GCVJ+(\YMNYBDU0PEIbdFEfaV?A/(cS@Z7JAO,8a;W7^X14019
/.LYZ@9)]fHQ_dJ+\3;M8PG8#Z4MU<>B6BJ2X8:0IIKeVEJUN:-<)_<H+;<ZJ0.F
/VA]3gM[769THRAOFIe:/<]=MGF1(K67Mf=U4,84fQ/K<eMaeCDJ0)-Q#[d:e1VJ
6K8G7fNVAQIJU:1=9.<TgR0LRfHN2b@ZZ[)BcgT)K_2g3Pc\+bc5Qc1T@F?=Uee:
N,E/a\\JG^2)O,.:eU6;D;1GSL[93YO^a<DS4+^#V7EE88J_QNWV;;b=MUFe6]>X
8YJD4:274A2;W\T5[eTVATE0HMRe&3T\A:9?C\P#g\G/U[3?03W>;RaY<ZA:OS&B
-F@)\R42,+<#cJ,&Y=]6S4B6dKa+gE[ORFf#&:&KbFRK]Q=TcBK=5g,TDU]+S&fT
ME_)\?g[@@^.UUPJC(7VF7M[R?ERN^;W+J/b9Y<(F6:\^QCDf@8PfB-PKMHZ\6YW
:@JO6T3GY0Y/Ce2TWf>>L;,_a56TDNZDCZ.5gE/V9.C=SX[DWFb+D_2\[Ucg?#IC
^J/OK((-Y77,27CWNG@>44bPDgZUY1/_fe_&[_\C\e#f1E.41_V?[IZ(#Y@A_K)T
@,1(X_Dg03Qa_W0N<JD#a:aa1VfPP,5.2J:D^c4dWX/Za1YYH<EA>d+dRcJ&WcCA
Z47&^^C3b94+W[.)+_=baVJY#DDP2WV,&M3?0L\PRUZH:eBYOcCV.af4[8.R^8g3
0EE9(A/WUgeMZPgG[T\IJF(M^G@aT,c,WA,Ce=ZNI/AN7PKT[IT00+,LdR@K,GQM
?TKV.9A9XE[bHdGTP)C1N20(_Q#g^C[_E]_SRL(R1fWA<_-g_0=./EFGbfVRNKW4
ccEMHCP[Me.cfL]-,;L)K-V&B;Z\SM<\X/I4WYZ_Q/74=d(@b.]61]>[(IH(da_.
<e\cE_aNVF(cB/I11HMP:E<Adg8gM(6/O?C#AFbXKPO>;SV?a^e7AdX<5,7MJ#gb
(c=bV(BQY02bR2-[:@0DgIOBeDB,>NeE^(&UE1GRUPR]e:QSbBAZN2HT&KgA?<dK
Cc=eF+G8gO\G/+_YE::LNM>BDCLPZB_-a1JFTE4B(N(#+/V-K+6g#JZ9;JR91\E[
04?[(<R;\?dLa.U/gAA(fZ-1.TQ1T)-ZTGB-E9ZEK4aG3_[MPHL[_JB2Cb=)XMT;
d>R&)ePIYd.=Y[/4K+Hd/U6Ja&fH>9+@#A@NCR\9aJ31(c857R?0?QGB0KaO@+.Y
,@S\Z@?3H[L+@L^H<[U.7H6;SO8&K;5H)3FAS,gY6>5IN;^Y=E2>XG;8F_4f:\X#
67_2Q?^.@;KL?073J<>N,_NB/Pe3Z=.5>[.g83ZcWMNfUaX2d]e)DEATKLNCFbF6
C=CF1_\;72R==b]._M8_=/dDc:<9[^K.#<RII>I)2IJ/U=]H(72G4fD1dX1?3^/Q
\]C>6b7gc6eeV+];5d?/A6F+fR>T+GgO)Cb)&5YTEaIT80V0]H47-)EQ,faGcNSf
fcf(+PD,bQNgMWG\_Z/[0>ZNL\A2Le?U7L/Q,DXE8QYOeFE&+U;X;5HK<d\H_26(
9M3#G@K]9>R_(?9)?D)B0><M#[[?LD:)R^Y0dERC#NS[9_VCa^A,4,,0:+4#=#+;
;(QCK8=IDDZ9HZ^(3WR<F=,((UE?TMB&d&\>YLV]=Z^M6?X\F3Ef+63VWW7#QSR<
Kg1Z;/FY>-KVY,&]]+Sd7PgU;(4I]2Y@gRTNHU(K4OP6@9eefWG:<SZ+G12D--R6
NJLV.Q3.F(Y.Q\Z)99K#XH)CW#Pe+I),@)=43=A&:6g-Xb^L@ZH/:?Q_gC0^J.eZ
:XQ645WDWE?UQQ]D?+Z?dA^Ucf&FIF/T<Fe?=/)cW9YS>Mb:M1)P<8e[cJ@>UL:_
OcgLFbX]SM/8[?c(ES>\/aBO;=^4.(:DaGdQ,99Kc?a=1COG\:XL+NDNfU#)?.f@
:OcM:3,fg\Be9,4O_R?EV+H78_#:R+&cOG^A=>bJGY)f1:1@RN,.N_/eJ)]56a\B
AJI)O-2:,(JEfd]6:EM8H^7>=AX3WZBIB73VJ/fI,A2Zgf:a4eWcS]L?/gYD1YVe
@P(/00.@=VYb)J+&Mf<I_Tbb2O2-]1f;9&?&d(3FU24QeeC7X.G3-K0ST2J/T3WI
XF5dZ_a,:-]D0ef>IB[HQCB/[_\ODdY8KZ:;X#N\7M:VeBKI(_a>(=KW4@4HdAHR
XV0LG[85G8O>E=H+N&S?:F(1\dV,4A@.]=/RZ?0=PO=QKN_\c7->a8/^L\Y;A=2W
C4aZ?(1+O72HNM-d=#\^5YQdRa+6(8OD,2F6G_CCB50H1V_R.-Ie(+GW\2TRT)7C
>G-LTM?D)?NK1]QRQSU#ZMgI[)K[S[<.FdLP]G@LgV2@X2(geWF+?]YLV&BEa?\+
F^D7U[0=+[-SdZMLb_]0(Rdc1+Z(Xf&L#VG8.-1G_/E_S<TVL3<@b0ZZAF5Tc.b^
=\S):XIN),a6+1<<gCU+TfV]fASHc]ZKO>YS04DQ&SF@3ZS/HdOb@JH\4YU<fU0B
)6e71;U=6L-#0\>_3G-7\#OL#49R;#(:b,X;QAJ0W+37QNSW7Y1RX?P7d&gA#GP,
7?Z]2.dT.Z&QF[UXK+EKJ-;X1eSQR@#GTSU.4RR7WRD];W.SYd-1?0#-1Q<.3BP#
HdVO4EZS1A9^_M<S-Jf4VEgKBD,74dK=KFOJ\RIME-#FLZb(1/bDb7_7T[W]N=LZ
:1)TRV:Y5+40PJ1)c3.)Y.?^:AJf_CXR,ST/4YUWYc6K;_gFI#YD#F>41@(B>Y:g
EYb?>>#]fO0P):SWE>+d2-NSPYKN.8<7(EDT2a^e@a35UD.Z62K3LG<He^NR;4SI
=&?#44;[^,QMOa&1UN)P,:=T&Tc&HSK2bN+@ce^H,&dYZ>K_fGX)[&8KFJaL?31,
0-4V\:R=6=c1+&P?aFA,QQ&>G^Q2N<aTQ32;D;F=P6TX]X8]<_c;P[L)K)F/APc#
;9:X<).10G&Z&DXc78]J6-&]TFD8K)(<;1eNS6R=DR0Jd2.W?05^#YXA:d]NO1_]
(2Mb6S4]JDf,)40?6c-H=GDJOAJ)@]8R-9UR/K,)A20^V75&_(X]gL.-(TTV:BdO
c8V2]5-9D(C85M293BQ+76^8#8^^Qcae0I1bMfa;;P#4I@\aX&b.7YYQf:&a7/d@
(fD)#abY?>=PRXf:W#=;:/S&_ARaD&S=R4=1bd7O\..U)Z.]^-Q&9RDXXY[V]a@H
L;<AEeg(b]aO9XML3^FBX,XXKUR_.AMgGXB[(</#67;?A.\99V;T=3(.5.9c.>V8
1(M-31RL+..+9VUEO@>2#.CbJ_dVeS8(.,gUE8@/ea5PZ8L_U.ceS5<KVcZ)5Z?,
W\V9U(\fX0D0c+<Xd&YDac/\]_?.LULC-?SS(;[Rccb.?;eGVIIK]cJCe(KT&UD2
VdYCY6W+#]YN41OM)1W.CDJG6ZTa2\TQ:c7TBZ(OOL<H2Z1QU6/_]-:LS@;;.[FR
6BH#93W:@2[KGE7bfU.g1>a4=\)_0H0R&TL-&UVS[J\6/P=2gF.0D89#SD@H)bPX
;9RSRdH-<\Of2&#[<aR_#-;Z;7\f+D-QXN4+A<P2c-Y-JfOWPS;,I=\HF?N48.K1
F-;7W@2e#1X#@IYN;U2.7@TE+@1eH7_GC;GM=)AgS7WNaO82D:R\Q)U7TA\U>O=H
>OU-DW3,NSL:.W,FPDNP:GVf#Ib&_bV&KI+@a>&9V]9E>;3.&=YdO8G)Q4J4_d#@
AM(3YK;<b]=S(X?D&\.SbfLJSaV:/(FS,H[10?Y7UL)])TfP\1:RY_[HR;[X>P_H
./83d3deP(_Yd;\S7D4cI@719Hg0KeS?5Jg5,0;/fZ//7aQBW84\?XZ[I+-=e)J:
U3\A2dH-2J+;OW1Z,9?bOE;(6Lb]e&?634]0U_?;d6_Y47C)=53cC1;O4()dPS]f
g1@FJebUa/NNN1+aY15[&9@>aG4,_UN@^8=dJ?EEe7@beJ@1R34)N;A?WZ-C-\KM
\PJ]ZGW6VWD(,FR/c?gU@aF2EYCB,>KQ#FSBU2N8;H.c</^A5PBS?#DbLBX/VLR,
SHOU3@K0UZ?@+;&J_7SI:S<,0G99J_Db7\T(74.dPV;/fHH&=bA<2?eHYKbIXPX3
A5Dd<g#3Ba9PIGEa1eWISc[ED921,V3WU15U<[Ef6O0<T3NEM,\LD(^&8Y^cYO,E
e70Z.<]3B/<7<Jb?HK0R=4b16WN4)SccO^[_)++,8:KQ##8U:5V^NJ-DdQ<>J@Q;
f:7XX><#5,,C>CR\PRD-L7><2&_#=.+5+^GX3Y3NL;ML6ISG6TL.WMA2V8;E-@fd
DK.[[eW+I(N;G3V9JY>\-@=A(7dc,N.+0:\5M+UW5aZ)GUBecJ6U.,YC3<;O25V-
]Z^d@g65d,C^ZSO7.37K1.)#-M::Pc\M+JP&V[U7fKV)5(_8TA:K1bG@.)3b-)MW
>K86&3(NK4>5#/eIGX=6B,D1RITIS)Z7(FN9\9WA-.0=F&]\aJ(H8>KQ4?IbXbBC
_/S^0L64]EMT2CB)&3D(&5P4fI_3FT#W,,+dEWBfIcfW_;SM=A<Q:bVF,(SAE0b3
]eg^_VI0O2H0d8R7V#Cc954\3KD2Fcd1PQC])9eUHN]A#)^X9)L;b[Le6X-NH638
7L>E?]g+O^/EJ8f[O0O+=a<N/=;c\M+-)M5@[e5E-d32#KA]5GY@T=A(J/eXT)bL
_V^cK4X.M,JPDaPH_9<>NeZ_&[MANF/^e:--&U.XW(&-C-_I#@=WW_AOVS^C:\K&
B.@YNQGAEH.He\;QV#D-@F2?PK1?XF.T3fgbZN(\8:,Ug<g[VHY/@8CQQ5eG;?f4
04Zb\N+<_bJ<F.GX,02E<R<\b:;1COU+_VCE4:05@I_g6W<^;547AN&.]@>M3ZE_
.Z\3@)81SaVbWaP<eG279:^>#0\1?Pc><,WC]?6:(9<@I<GgDYe\/dG^B#G[]\-,
-g](#\)_ad9J)K76)H6dA4bdD9?eL7=<36.CR./\>TKaZaZ<>c6AY:.ab4+RYgPT
#AT;AJdJJ5I95YGcaV4Q;XfK-^ZADY8TGNeK/&@2WSCQaN3\K1bPTdZd01MPWa&H
NK?K,3+;a/f-,)JJ-O+JJI&,Ag#dR.TJc;a\?C1-VQA;F1eUYgH2_.]O44ECS5TZ
.UGSaC18[0-NR:ISH5H2V^M]&IJb^LKVNAYYRJ\c6+-<=8^#[T9>(@?#KUS+RB=C
2B#K0X>Z/(AYAZ9RH+e9KJ#>Ff#XXL=CZBP(a7UB^4GD)>5M#3]DcFU9agYK8c]8
/aL\9B_T(+SC[(^4WAK/#@:&_=:5@0(FeZ&@JX?IW&6168#_B;77-AR4^@b/;ad[
^cJ:Gg-D??(UaQ<4^UAHfN7P84M,^CP7;247f\^LV,#fYL01QEMOR\KAW#7_H2K,
I[DS;C;-eFZS_AI,CV#?8Zb;TB>:RFa_T&GRL.FC<B>MQZIVQcYN:aWYOPIMVe75
gg(B,TS&NH.[;4YfYNX</?CS@19H]NPMT:-]6=;)?F\F;I/f&I_2T+SDMX=&dRL6
J;fOQYF+GX8C9<2(4^J0Q.YZUEN+9+38/51;VX8QZMZDK1F?[\Y^X&^C<O3Y>O[?
;98,cBd;R;U=+U52dLN(MC6PV8BHbLQZ#Q:E<3./]5a\X00C,4c46@3H<#f9W7O6
D+&P,NUG/bEO3a_N467fW1Ha<,)/=^7g78=T=<f-FJg)Z:>c:Ta]4[=&LS6W0WSV
=-E[^EB1VE/f08(7)41.0,XT<HQI&U[LgD+.d@\@N^-F4bW4_]f/A-WWK>,PCB^Q
=\4Xf_YDNV98(g,b<30&124MQgO35X@JO#,.)S\H1(P5FOWg2O/P4d6#7:LTCf58
33<BRHd8<Z^=]Z1\H&=JYLNb&\HV6YK:D)3E79,;8NALAS3,#RCN55L94PLDa3VR
P;&+-=2RE-CccB0^1+(>X9+CRfA;,O^GR[O^UV_>#8;22HD9@RU&EQeWD-F^Y<W7
V(FCKI/>CYd0<9S0SU-;Xa=HNfLIKWPf_.\_+4a87C<^0K+(e>@F<3#dE=VWKf@^
[>CE:&T7gB6fNe?STQ#0eZX]M:QE:BQ;#0G/9;LVYbE3?e\KS,1G7XcL=;=S>:1=
Af)1^.04G)U.^IEL_6ca,X\@O=\eI(@V<EJW>4)/1V]YN#HY<8YI@/JEadU7;?E0
#Z.\>/C#ef3V.@?JNgbWa3/A3dZDDI0-6JFfJD:@6ENUSe^5B#f8/-\,)>?7Xc<E
1I=_UH3ZWBV-WV>g\?OE@KOC,SBA@A<ZU8XRFE))\DD9Z;HY0-<bAb6f,ZIGA[0+
9.:bDNeT.SRgUMW>)eLPLAGPfMfI2/P?R:e>2VJ<D86S#:9L@5>ZaQN]>5V9c?d7
9Z32#d1SB/32FU>bX&bZ^\aCN[4KU\.aWfc<VKNg<R-L1b>(2DPP^W8B3OZ5O0],
FI6AgK[[/HSA;\MH--H766B&=M3FOVT#0)]>PL,4f4_THVgE<GbBL8^H\f+_aKG3
CCX&0?_.C=g8YRJ.&,32HPfd9K]&X2=CPDSQMP:=^DbV5O]<ICE]LFC-KSKNP-=:
:2P6ZeFOg4U\G&QH9[01LWU@f8T:Ng?_O0d+&cgbK>AN;]FH\)<@4CX06b0W4Nf[
^U_XHe?V(;Q;Q:5L[R1)GgV.?0:UZ:SRS#Me9fCcIZC#WV3D6^3@WD/GIA-N9.c,
Oe#@PgC(gH0-@3Y.ZV=F49ITCf\)S;XCM[=CBX]X/)XA6TT+=e_<8@K^5^d,G2_.
#T\P77A]KOg\Ld1+>8ee<aD3/cGg&+KB4b)WJ-PT#e4aBeg6d>XH@-:WGPYFU&#&
:H?),41ZU?U/U&#+\<@Ed5^[0@BJQ;]FD9X0,56HaF&N2[4fSg4Z0O=\+4=dB2>P
08gXf0XWg>>-;Y(?gTaG3D4)/5VD/J:;N;WA?5.\W[.N&X\J4:2>dQQF3#-,RCZ#
3=DQX+Q.46B9Q66FEC#P+fOO+<#4>[(01&/c.9P>B3.RDIM<0A]7Ue]]0g;/W4O(
3YW.L)5TK/<f:a-<:Z+D9H2,=S#_e0_./+GIEC?[-f89@50SLMM,1a,=J&.UZ:+X
15B^U>gJfB/1J9e2XZD6+_NgU]U2(g<72281Q.aGA>(\TdF/N,L4Z_ONYOLDTcVE
R@e9J+M)]M^PW(B#\a:0IC54I6@&Cf>8KVG)CC[0FHA5<5KB#d4KO@MIV0@9C?@Q
+3?NJ=^9(,2ZUU[U;6N9?,CK,VV-7])\MZ.C&:_REA9P0V7V;fWEIA^ZA\,U21(4
A:VP.9=&9deb.^IJ&Z[LZH@9J4#-JSCZ?.PYVI<:&(SM>U-G]3,@IWecOCJ\L8ZT
37I&,VVZ><+dBO[3/\)c)#dOcg6RUW._W)4E:_(WY#C\(_Z.aI,?1X(8b=+,Z6=P
1/4JT1\Fd-U2UeNZNG@6-3@.<SE@9bI,Z>Q&7#<cKV-bEDb\SaH3CgeHX3R<NQW,
ZW6G^7U[]VNFRgE\(&EM3T-,3FeB:bS?aPA<5g+:1(_E1FFTOHA4DJSe5/4aW)T;
AH&\fYY=7OJ>IReRNMAG)1EC:KFfVMS;7?YH2NOZ5-3^O(Y0^<(N)9@0M#76)Zb^
?+<_N[H0[H^,M23:e<K_WF/2@&V#F5?bC/BO@_[+FER<gJ[QV]9O,EL[f(LR7R4<
CRLNC.@,]CK07/Z?6;@Y>B9@Db\T:P.@f#MJD)_LH4H_6N27&AM0YAZ6L1(\c@fA
&K=63A-7PaE_D3Y@HeCENTAK2RL1]D+^6C&9\Y,F0&AR/(@L\Ua]#@c8J?NU))@D
?cccQ^aYaeZL^W1UDD>M3gZ>?eeAU=G/\?ad)fc3g)2#V4P8>GCeE>=/>WRQ;EQY
BfE0I_.bZF+>B<1186aDbWNaML4X?XH@e]fM7K2<H<#GB5+NJ#cQ7N<bLA^(2b\4
C?HTbGMc\R]U.JF/_?:T\_f-GAKRV;(gTDFZONN]3IDd?G?eIMLZf+#cP8Dg-]@f
)\BaS:1)TN7+]\bG,Gg^QAc(,Qeb&b,P3d47_I4G<=8@^aMaWHI4JV1XD?,d3bXQ
17?O4TCS\SB)PE/7HHPI+_^?c<>+.R#M]<3c6WT^9&&1SW.VPB_J.Ga-G\\1&3@-
c/,W^^Eg,^aKNB8g8CAF:CcU@IUOEDfL:1UYdCG1.L^-;.PdE##0,G3;D[-/?/,\
aS>QTP?8dD=)G#,I-3G(\b0T4b;WH)(2?G@^^gaTO-T5A^N=2M6_#EV&EDD;(B+E
.4NWg/D./bdbY5_^5Rb+6dQ7)(6gOJ&b9\EG+77/aZ+OW?2[[@^5-D#8QYXB89]E
5D(:gE.D:ZIWgeg?E-?4N_]3;:O14A;&-DYU:9SUO]0X1AX7VR3(Z1fD:_b7)aE)
7]XdHOS9T,\M)@9c3C-ULMBa=#@4IX^E:_L//O[W&2\?:ISGISfg[:B?O]<?T?H0
]:g:OZ+?8&X>A9_NS8eJF46MeC;G>C)U0)1]eYUT#QC4fTd1^:EIN(1HFN<JUfZ7
0f4>C(A0[Q2:V&,NG,QcgVY[X>KHZKb.fMT&V>.d<eX-2IT:WMF:K,gUBC6T8\g#
VW)Q@SX>bFR[/&>L0L,TFXcG3(:]<(I<8T3A9LG9:Q>@3;]-3F2_=&=GL:2_+7^V
G7fCG>A)(XH4M:>MM_/@d]HDI-:MN]OPW_:[.3>4.VO[0,\3KWX]N87OMc,dSS[)
c9,I+O[2dV#0.,b:E\J5e;-3#?Z<__fP\3IDafdSU-:6=ZO3_Q_Sbe]5<,^&LSR\
YDG><6&fYWS59=O:W4Ua<R-.J<]MKG.b-LP67B8XHXf,?@Uf51g4@V+FQ=#Ec>dX
U1XW(DM<AF\c]c#D04/Y++bG]WN1G-UQS>f\(f(2?4_JI2CMRgW2.a>4@UAZG=&Q
T^DZ7SNJ73;K(J8;dN:UCN0T3RHAOKb+5NN&L@&SCYKbgR2(J4@VP\R-A7M@3AXB
Bf=7b_ZYOf5UT1@EIT.aNY3A6XYg#<O?7c)D=2APE:,5.7X4c/)#cRUb;./:fG3]
(1a?YCI4&L29S0@9L8B&A,IQ/^I9DO3G_@HA/Y:K5,90MU-UZU/AGY+==Zcc-5^0
Q([_<\(CGI9B<QY>fA<?)_:E0OI\7J=0=7DHOI,)-9(W@@b/8K3&5)C>9bJaZ?0[
N1>3K+dbJGL>OF?,d24BY/#U4/(a?X+)<#19:0Z=?XJc.6fDN9J-.?PS]YK=>LDM
-T1S[>0V-O0DCY/XXWI851d&ZO;XS&&-Q@11CZS3LD.1ZT[57-^9>=B4X]/S4_;)
dM2.#D6a(N&WbSgUWDb=Se0--S[bT?@FW?Fa\fWMTDUN,Y5d9=I;1Tb2A2aN8;Ib
ARL1a7X2QQ0^ZYO)G][8C5#RP9P1DYWI9\XS7^\_SA?3?g?2/b5@cge(>/PHIB<I
0Cb/DL08(#>;GA5?Lf<&JdBKOA\2-@Zd2WTXbMD3&C)J3[?gC/acFd>KUC@fO9ZI
;([>BX+ZN?e=4g/?@c&?E(Y@_=N7])@5HTe=VGE>2Y/[&X([dE:eG\[#YPNN>OW#
A7QU;Ua9WQBgG>9^HL6;>1VcIR;6.#5ER/Z[&W5.V4\&AfP1D_]2R60[E2Z09+1\
)02Bd<2?O9ATZC<^[6K:1(f]#9(C?X#V@6>:ba?TW@3WKE8OWZ0[,II9B7f8>\gJ
,;\.AaRJ.MgJ(:F,\2):aG8(9K+<caA:.WK\XK.C0N9T@=9[a)HC6)=/X-Z7F1RB
b;]S7PbD6NfZK1/.,/0g@N/:)JeHJD]KMa(XVPg#SX(6@ZPgSVdcd.A9.7T<\U)b
;@QVe3\X:3KL5_M](U8/@6_OK):(XbO^_<bV@N2/RH+Q\gFB.F3E94U;W1G:O(,8
.NH4Lb)d6)>M7>A:>]V)f=a2]GEX[RQND^F<##[g#G6,Z_(<dK[McL3Y]W>FgDF6
gd=C,IH.(@WF;JLNUIA3fg)DK@9cDQ;NTZ&214F]))THG2.:P@NP[9.]G6\J/Z02
E]eA7fRG/Ue?&TCcF6e04B]g_HMDXfQe9aWDbB#2+&T.()LK=eHf>?L?9Z)MadW,
MB+LVMMBgM1/dH&F-#O,/^&3+G5ZF51M95[L]0cAH:J^OO]U9:L7+]A6_Q=#0V#1
0LB#;d>Uf2,g6EefQA7)d<,).]&D,NF/H17W0cP.=X8#5;(G3^?X^_BTR?]U&>3_
L#.E0(9:C&e56G8:NQ->-PKBJYfe,1];e)e3#XBY)1?I1\cGL&+/A,=A@TKUK:6d
:9MY?gMKgWIEF\G&T5UD1&DT8Z17?=,H:K?fc7Vae^77=.0a5/#^8/O8J6[Ug5H>
3A2NE>,I^;).O\GPC(;G80eWg.L1D4Zc#.QTfC#\F>#TZ[&OWO=(eAfd(?L,.;S-
#FP6K:WFS3F&/_/Y&=/73QYBT</9V?3)3@2Mf<T]2_Y0.#.4L;I5?/H[VRB@NdP^
6Z1J1)#TA_=_G3ZB]2/LA[c2O[W@,Q4A[S2,;BeN8.?G?XBB6P0a^#ATZ9[WQbg.
]WDa5[0OSU5MG8;/UDYYbT)_(F:+M[8_W7SIFL,7:HKJ;I)N3@[Z[ON(L<f7FF:K
[LTOVAbZT5L(X-Z1L:/dMN4&>)C]5?6((@8fb:.H8R1OS23.CP:b][JW;f_-32&7
ec;E-E69B/:X,2->-&&G^[XeAR610N]4JbK15[U14RKZ-IC,8RD2IV;.77@I#[0K
_eM58(:V7Sbgg@e=8]/+/4T8H8FP--L:=E0WKVANQ:;bYZW_?07?03#RT-2AD=E4
Ma@YGf\7-[^c\BX9@^4H,4a[9>#dOQFDD>fGF-QUdNZ=;17\Y^-IHUF[/-GLP34O
R=71)0;M7_2_gcDcU&6gdS1H8M_SeR?XbX[K:T/0B:\;>>;H<0XN(3aBDKZ\E3cR
aHe6ee;1=VOMESCZFUA(Y-EFQ8<#+IY,VUNgS]R+b=3<Z53MC+/WX+=,^<8J[>.J
.?Y7)fWFJ&>Cf(I5aVA&SP+7g:SS4I11GI4L2_/[d:W.H&0;cD_^0;)e[&Y/?e\-
/HKYL&_AA>GA?&VY6TM_(JQRM[>MT9T_E(PgAE=OIcUAY6g^eDQ-#5aC+A\DAf7<
UZG@?QKg>/OFKMCE[6YL_N7)7ca#[L;Y&.R>KH5Q_&G0-J>Y0+3MP^/cGM6Y,;gM
XMI+=;/Z8D4L1(P7=)[8X5<[G0d3JCE##/QD+8IN?U@,OIO+([eH7(G@[KBR(@eT
UAKUVLaZ.(1_?a9VUC.@fRO-P;T99-STgN?e<3(JeYDeAAfc3R+)A.@PC[H#T&b<
2dF;<C^M+1&94/f]>HE4SfHQQKZ(ITMdE67Hd4>#HK4bEQ[<fa2gg91O0/JVeH6X
SOXcA4WX^HU5X,bI9G?(5/U^&UdeABM.G7]C/@L=X:ge7_W?<HPe1MPg,eD4db7F
GN5L)<<Z^J.cccbS63ELR/0=+c4C#UIP7aM7L3DT^UQ]Y#cK_0HR-;RaeOH-Fb54
e6G96NF7b.Fd.VT#XYC9>]:O<87dOI+eS)cIWTabaHc.:VPbJ)Q;<Y1T6YX:B#e-
#Ddec^8.QX4O>JT<<A2ZR(P9ODL]P[B/?U8L8&LIgH>KN=gS@5CA=;_X609<SO+N
MLcHF)b:_KZ<[F4/eUK[@EU&<J><CLQg-8)KZ3,1SD39L3N\WXS<5#-B5MQ6+C\8
[;+DNTK^:FNR@(GRfM.#3POB)OGd-_JA+@-BYF@QF#HZaW?-AW+6O.4d^4AYA>44
7Y<ZD4>T5C7?e<,9>fFQ+dBDS9[I?IX:S-N\9V&]G,f&7?Z38^PdIf/>cYQP2.::
L3_7BaGMaXY(&2a&LM2=1=P[K=?0C5PE1Z57RK+cYC8:D/-EK/_6XH#8?V)N8WFB
TSL[PG@K@+:0OVDfbEU]D=R65ecG,fJ_?+CF>+>O4B-_,-@J4b8b>/,-=@Y3=DY0
D:JfCWe1QN>cHU8PM.1RR5g<;,4AJ9;7,V8Xc]H(=D&GIJ>5c+3G/D+\BX94_IP@
H\e2REK>@Q=5ZdaU<=N7BT8[8Q^X>dX,f(O\55QOb>..D6V?H](Q9V4eQ<(4=)e(
+g[<.;gC0L:AQUZCf]-#.\>AH3Z06FeL5UH>deCeY(8dU_EYD_B&>4HYfWMZ0\UB
TC122:S:6KaOTD[@BF@DJXTF567RWALQ]?c#GZVLT;7#7AH=NU)5aTPMV?:=<91^
5S#E7Z0M^J3.W5MM@WK69<L(,W4AHJC51O_+][RbIF,50&20;-S/d>aa[4Y;QWb:
5,X5;a65@Zc9NL[Zg/F[CC00E_d6\8fBf(@#MPXAXYTV>Ce+T&]R7eHe[>,adcAS
aJS5R<W6B09=JBAcdX@NRA<8(@-?2gKOH.G02_CPe5#_[KfF4D9KI(eD;bP3d4FQ
71QdU#Qd)#WBf7fDC&PQg;/DLJF-O-f@?MV^4/g<L7:aT?04?5KXbI-=2M]KEQY6
ZNc4<;6:3-a0]fK^d]FMBRKg)9@Q1C5,#YQZ3D;&1K?Yb9=@)JAT5O5G[?R@E.S@
(Y5G78.G7-2^gac(65+9<KQ-_T//A=XHX<;>&O@9E7@H4>VY)bJb_J6\B?GE7L0]
QTHJAG<]E>[<@4/,T4S\&afB<&bXQOQS7]K@D&;A7e&,/GaHFVPaeGIWCPC?GQ7Z
f0@D<KY6DSe8>1U<1K+PC#&^O7W&9(/Z,geM7\(Id7dK+W<gC9?R6XG0SGacE2W.
6SBIW6TBH@CNC+\/5?.R_e76;@&bOU57W+QBI?,2:(6gf[,69P@OaJae-G,]\bD[
>bd9DgBC\fKQ]IR+#FS4e^BfFI0K/2M2Z@42L4<[LYDN1HIHV7YEHD>102+P5/g#
H<?1URXD&:Z>3c5BOI@1HLZ1KH(_=,NYU#dGO^ba8#T?F@&=1<b[MDb3Kd_BLbPN
5WfC:-Z?&aY-cNO,;O]eb46UB?OU.A+51LKQ/]V#Mbd1#E)8A)HI_G4TQVD5XRY>
dGU/;A\5R6aBAHG.AEC]9BZAX2Fg>Rf^YbE#01CbR]+bMJ+IFD=YRDQMd_)SF_.H
^91ZS;]/RW6.bKgK-=MXJ4J0O288HR-IBS<cKF2649HgNC6&,)7\TFb.:a^S1c[>
#cFZPWP0CaLf>.d@ec>NaM9;&NH:)BZUHH1XV9:gffdSATS/cCg?3CTR=?XMT+M(
0fgNL1gTLZ,6e.E+C<S_,DLXbf(b]1Lg@N91PK8<YEL^YCg4SC^[-:.^02\3XGDC
9/@ZTd,baSY7=/Q<XY_dZ]D3\;+f+X??A8A[:a48(TEcL-Cc<S1)5K\S^IRXGa\5
d_??&84,f?]#;SBC@.M@E/MU?(G;=eVe.0>T\EA(^)Ue&?S.P[7&B@L\-9H:;gGY
53cWe=a8EcSNY0RJQf8J</g7.eS-_3_9&WX8&?5g>W4;DSXE;3b1U4&RQd.f,M\=
cVf7G<c@:K5HOSRQU(]a+@JVSCJ]L_V&4PR3XRM;K(Q)eUg=2SEGO,Tb7[?8>:+0
#c^AM?8>QJ=^.1QH@D2.1^4.Qd/;E\>EJ)fH-VX@2&CfF/(5bgL??4ZbG<YP+dAb
(bGIeFL4FXV.><H)T-Kf<D-RJa(ABcXGAeO(/.#4#C2Z=>[66\H9=28K^.@3O0/X
C./Z86Y(gQGQ-d#C9^+<[UI97O#[:9WZ:/_Ia&J15IZ&^f3cYbbS-D02ff((R7f>
S89G5I;>YO/0P.S;3>Q?2MG58.(@N.IM>7=3;)9gea&XVW2>LIJa1,>>>B==)B_<
N-(f]Y6e=)[O7[]TbVc:FB()T2RAT1_O&9S41LMX4[fg<DP=aZZ\62EHZ_F(7gbK
+2#U)WU-Sce?&bT;+<U#F<R:_eT.geW1ZfQ/&-?@:OB,8P6[EY5QP2GQbg\P-,5,
2Q#<#6)G@GQ7HZ6X+F2UU#b;A)16^-/<b?>QgD2f1(OOK1cRG/J]><f/e]0Ad;7B
/<4C)5E0H+\[3gG=A(MZd16K;SbGI898Q0dOTUD2d/I2J\-2=]-L?_Z5F&B&CaW(
D>+K0[XIWQ:f^SOVUN(d@T/63W2H/CI\.\2UYgO8@fVLQaP?XAT-^8gCN2O;+ZN>
^V7D3<=69]PT[KA(\_@OTbFfB>cWSCE4gJXQ:b2c)g0a=?S4I#-6e3PC].Z<>=EY
gM,LC?Se(f..QWgWG]A:8+;=dJC-6[6&?ccb,eYD0IX)M.+R8bA,^Y\Tg(\MPBaD
6N1L9VJ:DV1cMW2797KZA-SKc.=HF<&RZEL;_L>D>5gHM#b//OJ1Od??8O7YPIFe
K<^<=BIOXcC)0PR:R0#ME-L[4,3>Pe/&=SRbQgR@K8;d.9?9>H5UGTAL+9gLB&.9
1G454;8&&1_/8FZQG8;VC;I<LW(D7/?Y.CeCSU]<AOSXP2/Q(+5SV_35_DcZH]Y4
P/]6B;?>+YQGaQOab2;KHTS=VF-fM=e=06CX(c=YDS=L7C;f15/OA\e8ff-fJ=PU
APH]#H(O8C&f@7e[.)6489^]\O+)#)TB=\F_FGZX^NaDHK>?Z63cX2a]&,]g12#X
>Q+6edB:f.X3A286&GC^KZ+M\AgL=[BJUL__fR7=QdWFZ:f=.,abI;(&[daXFEg6
gO538fCPQ+f?@d]D)Eb4cA0P&YSU]S?bD]f^J@M8dUW;=YNB7^-a<d5H>,Ab]\_a
7HS5T6TR6(\WX]bUWH,STX9Y##O&4f./R\RbfY4>^E\d\&7c.HK06ISPN[;:,:Y<
;a4Z;B2)L)R9+AaAZMTY1##bLe^EAX>O(PAFTMF\4B2U34CPRA<f)?gfFOC:OMUg
I=+5UNNA3WR,Y4:O,_6+<LLZ8?Q3=(F_DB&g,R8cc+F^X.[,>Z/1_VGKK.H(\YQ8
:MYGRf42F@Jc[(W&[2]([[I?H8?MFfA>0^c9&RWGXB7U]a+6?)0Xe6>82Y<TB<\+
-GUeF6Lgc6WBK\CCgA2/--ERR^)&,#WFJaYYP>2,F6(EYd6>.#@;=#:_QOW5dU=6
#8=YVS<;dP7DJ.\-AE-YA:U@?-=Z2@:f\59NW9\Q,dCa;cS/T@6==a.]RIKPXW3S
4K8NRV\+>)@Q-@UX5R;<FZTCUab8.RXaVW11RYHTI&<B0DV@^9P41LF?E3G2>Efa
fNKQV+OD,-d=RcI]<&e+T(<Ng(+Q[:>Va:aK6FC&RN0fMVH^ef&HWE-L=>=>Q@K1
<<35?G->JH0,5CaeR)OJ#/?S;eO?G;=):Cb+TZAFL<g,gZ;\R[[U4^13^?O7;aPG
K<cOQWNW7XJTLa;OA8,05.)Y(/[KB/L6bfaG[PU8U8IAZGR?)1</J:V\.FeJQ8+&
V)?3HQ:7V5Z[:AO3@,1^+dg>Lcf>(M-M0I<RSe\(=0QCbXODZ[^R&UMMGFXMf2>,
UQL56@V&:bI1P:F7@#IVUaQ+c<+,Kc&?[:FHc?628/_0X(.Ze(^/8Zec^,M=+#,2
T1O.&S3KWOP(N(FKgL9V53AWfbe)]_)fPd+[EYG(N.U/5W[e<HFR@MD6DX=-0f.b
#C)&YOZAc[fI?NN-8,Z2R2Z/^WDT#I.>6R[CIT[\^]Y=;cJF@0A[8:@59CcZJ3E:
bc4R#@.[CX5TCba.-WeCTBN<,<DRF=^D[@He0L/gFD+A<@&@f3F6PYR#>LeC+26W
@<L<_2#QWBUQg;,+gg-1#V&LA[8.<\MB3@4eZB)33Z+Y0>97H:=J)4\U3bc68:NI
NaQL<2&A\:g;X0,JgY8I-Y+Z^OYe.OM:6G(](A.cJ)\DEK(]?Paf2-b#<B@4,?0G
d7^OWZ^9MV^0YWZ?WF\6QTGS8V;aXA+eB=DM0+dH,CA;;J8ZZPWK/H^-5E;(eeBD
,G1FODQbDW?WES<f(-=IMEX>f<NVUF>::V]N>#Z(e5X&=(V-\NaPR)-).VEbZK]&
RV:PQT?CGD,:2YH^fc3/>aP,Kc6gU,CIOb+_<P[N+(eUA7\&F>YKV:08EH/DQA@9
52&ITOCOb>R;P;J,4VPeQ,=8]F1)Zg62(DBC/<F[ZUUD(KfEe1IBY^@,MX1Y:3HW
+C^K]PKNT(C4EK3R+Ved>E@3gAdXXA+U;]BFb0_/>R=V]TO<Y?/>5F4d,#IS2885
;M?2.BT(.H&ga@a^^V8=a5QBGV7gLg(TPI^DK,?43^E6+<,B]5LD91bHVQfW1Zb+
b4JE>7PQT1@C8@DfO<eeLMJ,MG0F=U9\CX]]>WI,=I(F8GC2f,_Fc_6CMAL<O)K(
3FP<E+>W-RdM_N7YgP>PNgKMHK#QM.FRdIOFZ]a#I+#W#]c_OB]b_@.U[B;12TbA
(B.)+@49)MO:W9baF\@)MVS9;0aHI7.<>]2ZIRf2.@EU5ESLD\?E;5628E]NZ/[G
JP60:\LSM12@+.W;]?7QB1PCR:.WGbYX[Q8W+7^2<0]#;J5Cd\OZ62ISZB@L@RCG
XJ+=Z44gP<bRMX-0S#V^=4XK8E0B/4gRX5.-S)=W,@,P@?RF@Y?2Qb@E;SFF3dd?
FUgd;.I9Xc7@GUPJ<)1G\[@bY4]F_\99P@>B,?6<#=7.0NdS?@)#[Fb0UacOI3B[
g45Kg?QD5BRE+U[2?LL7(<@.5a[C_4-29J=RWN6=S]?aN<&ZF4^JN2dI>-+I#+CF
F=(?176_BS\\](7W8IZZ,.TY3A(3-Xc=cG950P[_L>-:PT3J,TWOU2L1B.B04A/N
3)./[:C&&b]a0aI3b[P>&Q,-S358Z5>F_J6LJ-.2:P7=gVg\,1aX3#;>:OM35)NL
HF--@0H,KVcP\Yd)M1&]D+HgX1Q+WfRL&?Q,>#&a,7/gJ#?65TF5\_J-D6F1:]Rd
e,4U1cRQZEUfLS+7dHNY2&&c5b[5W>)MT?.EfY;d(>5WXY#-30RK/--D4VaX0B2O
]0^bC^,.c10A6,G<ER7gDT1.Wg[]1A;T(JM>6633V;C)B(=D&KRES-9bZF8;aVL)
.@QIJPOf+-=F3?76_)Oa;QF[EW5#43Hb/Z>IV=ZNdF;KQ[I2H.H=X8.,g5)XC\a=
7WaeAXV;(H9PBE0M@a>G>:(\-fVF61><-Q\4DJ5FHO/P:H&XL]&98N;9d]0fR&8W
@PgEOF=&)A?b85YJ3<KY3VW3:HJ8=5M8e@d,>d3QB@;3(c1R=#YR/J#-^]DGT_.9
/&[^_2/-IAPM@DdL:8TGM26:(O5WW^432Q>CUH-a/\:.0D^&DG,8Y@Q?MF1Y7_ZA
\NDBW=)]V71Z0WX^7_)>^Vc+1cN.497#e,P[fDUMgR:4[3H;]X1D&2&Vg[Oa2/]]
)AH):;KA/0B,/\9K))J^Sd@A<W0#-L6_5IEb0bL6O5f(,\PCS@faV1RfN:<ZWS9.
;&WY5T_5,/6D[Y)5]TU6SC_cP>7.NOf,#FIRA1@+eZD?MRPa-L7gG^A\bX9a&C(]
@]D^TX5Z4Y2dg<Z_ZT9bQ[S&.=^b:P^abO8_GK11MU#Jb[B)e&Xd@?=N:#36]\&]
LZa>9)HB.b\#a.;R7:L#R8bVd>QG)1SAJM9[9HF1AE@7Z;3^T6LM[3d&(dG1J.&=
W?XA,7/,Q,8+8J7b]cCRG&&#=^fQF,#.O=]I&W<7I=I3d]6K;;^M)0F<XSLQfH_Z
N=<6Md;C:OBLYbYHD\/#ea]5.,fZLD9UdXF&^(\Y9PAWQQJZTCf:9NIC5c7TZ/[6
+g4ACZFFDZ.EZ1fY(Z0a@<7^g_Eg8f[2g6aB@PI)4<_b1aM)?Td;J5c#?-2bD\f6
>L5)3H#B#/&-QeH1/(,_NF>(1#B,#(?XL0MUM7+/AF\S3f5J5XFf47)6.BPB;dca
Y#K,0X/\gX3VQ^ERIG2DA_:C>K=>WUbQB:Lf:b4OJORKM>^00?C4e;CTaI^Q(LcO
1W@1._Y9BBE6@^G^S2>Q&(S&I:B(&\V#IWc\NI+>9/WECgBJOHY)SS.c(ZgI<>,D
e:[P\;fI#]&dQMB7,R@+)@06W7@H]2AW4?G;FS16D1CZX?^O.7W4^Z^/;Z5[(^C[
?1>GYX>OH;UFEO1Fe(;?CE<ZH56HA]1]2fbUY),[?L0L<)4D(YXUcg?NG=+E\d=3
R<S3ZV^0&=XfdHJc811A39VT[.0IR=9cW(O^f&;f.6A7U\0G@M[YH+CcV\E)Y)Je
U;/=9V1.3RHg\dZ&M46/NCUUc2<Y7R7=QNNPa6QbES^.dOKOL&0W7W()4dBP:>-^
DB=/Z8e4.FVF=Y=32J;Oa54BEc6?0fI@QT+C6@e6Y2(@>5]/51@Gg>P[J(-26O\,
SBDYQ&&RM^H3Y=0XQcEEON+9ZKSWa=5H7W_#;E?-9V#Vf0\\Q3&:S#(241JQd^4/
B)(eR2-&@DWB\+^3#&+[N6Uf#;3[\7:;2aA@-T7<^5.J]B5A\[5(9(<B>I?E5XSa
S9S+YKQ-[KAVT0T@fLc]Q\dK&aYR1,d73F+.3ZKVcK6f_RYG06e5Xac3cEeMYL/4
PHg-ee-&4]):=Z>W7D<96RJUIB,Q<(N[5GVQ@09@NA5>@dKH>:e&\N>5\#8>e9aT
2(a.GIV6)[cELNP8:SbO?DGF?QI2<Dfe?]TMJd5QATYgZW+CAa,)7-,NLG5b5eQ9
7eZ:2Nb[GO1]462N\bQW7>QDBg:_C;(/>0cC[(X3>D[E11&Yf/-SUFRW2/&^6gA=
>N171bI@@:Y+H],T3T.39\;Z/YU;@BS;N=N44FZ712-R#4#:g;NX^_N#&3QR1]9[
e^&c<63@,A4]QJWb@ZFN=HZS]SNKBZ5/JP,ON5AJ@Cc)_4c4)=d3JNE1MNI2@#89
E8b3-?fISd^Z=JK63&VA#Z#>><,M]VZ1A87R?6eSQAd#BI^EVf-E,44S<YdA7DKN
/UJaCJaI:L<),:?a4E&0?7/:/\[<N?3,g8LRZ5.VLO]5)?QLZ=<ZK\G\.d<_1L1B
Z,:N/^YD/IMUS&B0XP6H-,TN71/b,(05?]Z#1L:])TR_A0DBG8_H&?_^Xb&X-:25
Yb&I;;+_b/EcRAM)DMJ4Cf/0>K:E&/U)2O4F:OX&JRBGcCa1Z(;+bWN7M?(<1UIZ
;#/-O-f)1E_FRC1BgX5H9@M,97-9PX#^bY@Hdb=RM/(.KMEVM?]=Da8,9>X:CcS=
_5)ZeJ6>5;N(H[8[U\UNM,KLVA\;P=0MF\VMM8#?F]>c#L(VN5]L,XWQRN?aI?1]
=fI1@3bP9F/)LISV93P8X]AHcZ2/HN)RP.-=UW6GJa(CK.@[1D#O^7CSY4M47#F+
c?IQQDL4RA255LKAK@FXNd\9e>DdS-C<4D^TMWP:Le.,K4)EJ8^S1S<G1862GIQK
d@Q,PU=).2dIg4KNP(]M7a;3^6(Z1e2LK?9[>UPW)L^QD#XD175dBIf,@,DT?dbF
G\d#E@f.g7f=(PJ:.16Bd3f9GRBTDa.KD>\K\LbUW1]K/W78;L;A+UbRFeTaFKKZ
OTL\[:3dM]7;WXCW/(V)/0EE6a#bagD;22\.(RG9OMcH#95?VJb]aHH[#=+0Z@5=
KF.E1#I3GQbN3IU)^f#F0dW<W99#.@dMb^bQX+WEBH3\X3\?XgLL2@TL;JLfL?70
CD>gXTfbXBB3D6SHUg:^EcI+]cK0+\dc+>4>CK(\^-_5Z-DJVb8KT#9<>H79@Ff)
M@4EHD)_8e[>;H^P<5F=45:?PF[W:3_Ha3=.IS[L(DccQ8eH1N/M1HOO2Jb2PLSd
bU\#MJZD13W#K>b&Af^D#2O[B+HE?L8@Q^cSUHLTg2XJ,I+ZB3[Y<dKXQK/M?2MK
W884\=C;5CCFYRfG6dC&::-)SB:J^^3-gEdb4aPSEGMX4,Y01^Ic<Mb&?A6.<]EZ
T[YTdB)AG8;PU-WT@;]G[?=WEKG@>]dN)(-fXR&0J@8)P;VEN_S]JfS-INRb,DY6
J&#76OS5eOaSb4We=A4X0RJAGBR4=NTJa?^#BTT^+V&&fO4L5S@<]\bNEQ;=.MQ&
cO25_g^<,g(NdG;=G=6QKVU@U+\e^V,2HN]?eb6Y77K]3HW+X4..5-.TDR&M(.;0
Z?(N(@<A]d?\4&S5:7@U+]bd?YE+88[O9[R6NXM2=I=YPE/FVcfF<&6-aCSQ@_#&
@CO5^9gP9J+QWXK)]#3I7R7K@YCT2J7;INIS@^dQ865Ag^..SB(SJRV5W:VcOJ9I
bO7Yd<C\7d)&1BZPg.3+Ie>=1@)-\:+5P1,gIEJ>I-:I@;(K40gC/eL7XRM4[4\#
HFF(D+57&3S2#e3[@XJL3S[ISZVaQb\28/[+#Ac[=eG:JCW5cK=GJM]_Ee45EK1(
YBJ2YcA.P0WM6MRL-</2FFLc/=7>f>(_.\=>NXbbLCV<.O9EEReMJ;W)fKBf#,:Z
5JBFV=1E#H=L+I6SEJ.ULg-e\Yg?]AD>H#PgXSB:G@MS\]\Z980B.?e_,YYFf?Qf
Q,\^GQLKM/8M:a[#YJ19Z51STae0[UQXbV2-W020gHRA6f#L7T&JH0)MTH)a.g3K
R#f1UO)QV7UY[)[3<@?Qc53e=egcX9GfO\dMC##@]\b(E#_-Qd8;3\2],86;RZ&:
(GbBO[-3>_DRB]^Cd@A>J;#.K7bd1O2eXQM;HeMD(E7PC+VNe+ZLKP:[BSJVR_MR
GU55Y;-#X=^(Y8[=KAGP\J43gD6?Y=:WE&MQ&SFV,=??\g.?_UB>0BKL2+H8AJ;.
_PZ;0].P;)<5#LE9^W-:Hb8/Z4#1fCFOW[6P]AgO\2fK/UFG@2JNcO7O=bIN,e=7
/?FCCGNL2EX1L=8WB8ZBX6B95/Q=N081Q1&9(JaR86U-A#_I5DM][cJEQ[K-I@YK
_g1X_S?<;_]?OEPfM+XXZ9=VQgHgA;WPgL8KgJ=]M8dD_W[&?CfD;S7Of=^JN.GV
JET[Da;0>WGC<+6&QG8c61+6S]a4ffeO.P:bUfT&<X2=&JAWXUUVXU_UH@5d;c+E
86f\?Ob+bGQF7:=_CSBM:TP;(:6gfN/W=>.eC>fPMWMU+XOO\+S8]0e[7QYYc,-\
RWOdW2MPgN#R3K^M-M-N]143I)C:aJQQUa>fg&0.J7WeL0NE:-AE(A<KPIR&U)5D
?QE.?IRcG4(M;[_KPR@A6J,24ZG.R;+F=4-\g^W,,U^7I6VS=I]=U\UbDJDTb2GK
21;WZ(YG[JgE(:D;F<dPOH/.\)/0=RW2&.=+?4UCU<HOb2Tf.4O3e/+KMUVA=a(;
>]:?&[4JB8)fRUG.?2+/B(dBLZ^Dd&^SLT)DDGSF:a>DNGg8g84?K-fNS\O@2Y-+
3+B1gH?\N3NY;DY;=9fe]5G];\SgabL^/)eW8+=U:^,WF\/Q>6S_?\^CLDfD>:2H
16)B<>F[/VOESZGH4LWb_O/E(+C#@WJCQWQG@S[,Ve)YBBN>S4P&\ZTGPJMSJF+4
3UQEQaLTONUc59\8G>P5D^HO0_)ZeK9;7dJ;0>QHH]@DbGPa]Q1a9]B\KQYaY#:F
FT+fW<(7C99L(]DG/[P4IKBH;^5DLE4>f)RN)bC[?gaN04=N7;-Z1+@AEO@aDVbK
XU#@aU:HXWY)+/Red602fAP]a>-F>eQ44af3;>Z,8f>IGPLL3Z:Vg4820P+#eLa1
84dc40U7VRXM=<7;);3+PQ?AIJ4Mg<:U0=g:^RLQS>I,2-,:FMQAW0[MHe&AE?<L
V=:AAY#G>a:ScT:2g0.Lb[KIE-BH5DF8L8Q;g2NP5XN\>Lf/?^VBCDPU33=U^L7/
1L2F]>/OJJ[aC94EcS)ZYK<PVL_6g[\78V4WGT2LC9(K?BOF4XRC9J_bOA4#@B^?
R+X+-LSP.X3g:M-<;5Rc-P_TgX;#JMZ)@U8f;S@JAF/_R+/KG.Xa-&YQ^>fKN?.B
9N9P=#><dQS2d4f34XAM1gc:WE9\36C/XQU5/?X[OU?K@H;^UN54\@)fO]T5#3b\
Lb?99gCLDG19PX62+HQIa:\83]HH7L-0Ffa6XT,?T45D>T=H[fMX@aYS67YBD2fa
Y7MW4[0ea]9=_^5L_CEZL5JE;/E56dTI>X[1GQ>8AYMAY:>372U(O_EB7,#P?V[e
C2dO[&,CUFJa_.DOR<=ROZA@H218HV#?;.L:+H28F#Eb,,A2a?S>IIgc#TJ7#RfA
NWY5/;,?KM?BA(@b0TbVPdOJ(NMaB@DR+;E5_5;8(N\VC,g0GLHYDH1&#@)fEL5d
AM1NS@TeJEL7<8=;IYaVIEV\<:X+?961Ng+L#?6K@CBU^9;b;H=<2D-_-@a<OdUY
.H4.Z&OK;I&P818EfFZS7R/F?_J57ggb8bEfTZScf37;e6@7]L^)6J/35<G6^/C,
FgdaWeAZa9#JfPG=@^d#UdP5.)M_]Y<@BU][V46SFZPF?+b=7f[[+K,a4@:)/Bg9
(_Qe3d.8A<?W:)8W)]65c5S=GI@KEcDSSP]>KTS_H#71K_D\5;f^]UMD&)/)V^b4
9YH#ecN(b=+G_e2VP3PRcZdd_A:/:,>bT@DKGX,PG0#RXcBLDA:;aFNJ6T2>(_1(
C1/_)EB?I7888H3OPH#;/DU@.GUa7,WTM[7SaN>@;LS@U)8=WW,PSS,WYV)E1ROg
6@521+;/&EMM]36e9,3R,0.Uf]NC?BN-&DF+gb7eWLfea+f[(#b?Z[R9]],HNXBe
LUX#](R+S1E4+g=V11UE+OKI6YfRL&_+AD8ReQK:B?g7I@;-V0f#MX[YgD.Gd^1b
N_Mbd1\:gbaR/Nf^GTLJDG5@4>&K1C@:/5K8#ERVFW([Fd_d8L0?D;B6L=f#5d-]
:.UcGKfS1+:e(Kd9VL3cfI@6MdC[R:<GJYAaA7;OS_Z-1^.dQM9+\(-MOP.gc>ZO
<DSL&&#ZCDI-BJ&eEcaM\2CU^H=LF,=\cRS6VVU5^]T=R#b5[#F;DDM;HH]OH@1W
2,\BIcXR9D@;YTd5E+WOCI5^@IZ?)bCHWX3FXT+#_S)K?Xb&_=33>HdZ]gSeD>IN
DIDNA0_>&W9AQX?5E2&cF^(^B@M78?G+d@\2-Sa&[V_<9&8_PN,2<_0AX-X=0/=3
?5/]MeXLUc67DVc&O2T@FEB&:ND68++&]DCb@PWEHS^W<C/J.6W2DII>g?e8dYB\
/4adRC@c8OYJA7gaT^OI]7P,FPXg3c?a1MZ=7Vc)>1MeJMMT5&F8Mg<2DL[5c99d
dUFacSbL6fJ@/:<I=5IRR59bPa\0@T[gKM>,N(OQg+:6F5;#I.[6?PG29E5YEd=K
7--A[edM]98D[D7M+DO@&)<HLP[H(];Hf:Gc8R_BV\dXD_7#,;0+(fBd0.:K/=aV
>fI#)EWd26EQ2F+K&&]X(UAa6IQP5&ZG&S<2ZYHEF;^\R:,GC2CP#EC=JM=5N3<S
-C=OKQ,g1(2;6OgIV<LULI49c(72]3@eZV=f)#\\]E,7T<+040FOU[a/U(a3??S9
,e0&M,H2H]Q710U#029-VcDbM0K(@+adH<.?1_Y4O/f2:I41-S^d>N&<9SKTM:VZ
6E>W+:C(K&9H6KANVI^-1_gO4dA9_:[:><UOH-SNL_J,(FO6V(=Z];A2@_TdC</I
T@3gASQ]LNIU]M\6?H8IEd,4e-@1;^54D9K(D.M#4P?NCdE^S/E[bD<a46PC<O1.
(8J2C[^ed=EgKfcaB.#;<R.V;HF_e=G.5SOeQX\#G8TP\Zf./,fF)7;^eW3LSNQ8
V_Ke86[1?_Q1Qf3_WO^(]K0DP9,d;R/6DJ.dDGF=^DL7H:F\QUWN.EgK)Y_NX.9H
1,W</XJ;&6UF]M0eOcVVJNA#=X(f]L(E#OW52f\b-B-,dTYN_V^4^a++=80SdaE7
dY<1X?V3_C45)cL9I<BQ46N76IP#)bSYXbV_;^\OR\bCCGUOWK+^,b->LJ\FLKdZ
ABV?He:>:F\N+^M.\1:A43fbS4Y,b(#_DEDCfUCC)+OO6,DPOaE[OSE:[+WVYcD/
d,7A-[Xf#Y[D^1[U(#&g1ZU8&/;M)b]#5YG#Vg@B9fQ;?HNBBAKS9A.Pg172AB7e
0c-K^ZYA.UO;LM/Lbf/c4/YG=dIES6&(9/_cQg8^1aeZSIdLbQ8EY+LMaMC0;:YO
,aKCM_Z,X(27^U3(_(7:&KNQKM,dA7DcMIF:D\fM0bREcAC??N+ESdRCMQTc@AK^
eC31\A@72N7:EWA-=D@1OKX6FcR?;\g<K,5fB&3aSc+<IZgKDfK<]H&Ra/@fa]=_
\D8/cX/<+NF?XDQV7&-3M.>O&)4Gg\;DD=;g\T-7+6;XK<#R+Wc<?/4O?E6Z<XLT
EJH,^\1V3/HMP(IU^\4&X2XS931^Y9FM23ae2XHUfGQH.@,b5d]W@IDOA(5P6)Lg
,MTPa2?J(V2Q;OdCR(KC8W)03Z?;G&ZeORc7_BEIOH=M0G3-_b3DWEYFg;;C;U]a
#S@XPaUAKNYA-4+\LS>TN\fA[MP+,Y/9GJ>e^4CEW;JRV)ZD:c[,,1_AdBAK)7PW
e8+A6\7Me6a4gJd]V_3ZK&)Yfe_>c4_A(?X:+YXfTUGZZBGJG:8DP@O#cdNK0&0E
?7URP:P+#);O4e]BR6&feASYL2,+PZ@5V)Y+e^35BF=WFT6S_V)32>-+26geR)Vc
.#MWT=]4SV15a#B(VTDNJf?A.&aUUc+[c/d@cC5_O1SZG:aBXZ&5Q&XFf5?1?OSD
0Y;:SWM]?>Nf5cY<Db245V9G2:NS/LK2,/PP\5:C[#D=QG6R0AY5#L&GNP^<FKDe
bE_&<@ZY1<GRgccf<WTGJ-@Kb>CO]MZ<?OaCH.698OZM#J)dE]\#0agACGN+_f9A
-&O;?8;^9#ZbKcZ/2V2^<-=MbJ=Y283>^PBQ0,d2@8T;AV=a+.,DJ5bH6LK11+3Z
0N)M73R/\f[9GT&#]=L,#Ka,D:4RK_O?B@4CT)LcFcSCTZ)Y:69,e1Fd?:<XRaQ]
/G2c/bGZL84a^/aMXWe;JG&/ALO&3/2)fP<5aID9?#)b+SD^9SI&Zd_DD^C3K^d(
153WTDag\F0C?(EfHK2:We&f)\T#X<H[/=eC(1=VWX,We>(P7Z/=^7g5FOgC[LK-
eKg?1XUI/Z:;e\YZKHCLBZ6TfR\W,?0c1)_R00()4:aJWH8+aU0ZCWN83;a-9/MW
6OPgf]&A-:LYe(E[-XK(O9@,A[QRQ3)FC[@W0Y77K:b?d_11ZeZ?E(:gY\)]^E]2
>a5&&59FZdCbF(.K0@ZV7K(H14\bFg<F/H8>3J5-3QRbD&(VYeeBLVLb=f/CLSF^
.=Y.8^#CbUR[N8XbQXdRaf/IDe4)8C1&S92Y@;c/IJY4aBTGg]MP#Z:/<#SP_\^^
2P=Z&aXSeJ7558AU]\\+DWL#AEP;=+8203T\<;Pe//fVUB.TD=P17Q]].HU0PfXP
7NbT912W]_O6ZS2DY^8Z[.56Ha.@[D^F^G2fJYSCEaZ]4(Dc7L@+_:8UR_NF@L#6
_]MMUR^Z]LR3,F1T#D2(X.>:Xf/^Se1L]_LXa-eb)DH8OICZ24.R1=)?=3>;Lc@C
HDTb];M8@bVF=61^IR8T3#_S+DENUbaLC5AB\G52&YG-KTGPe?TYPRN<,=0B5@ca
@#AF<\.1-AIC_V^UX3VQ<,K]ObPOEM7Bd+0;]9R32A,]gHgcOIfa/U:cS>9\E/D(
.1WW=.HAY3:D3O51^1V:cRU8N0AfTTa3Id\NJ??WN?F-L9;MT4fTgYcRI>Z(DVaY
#0B?D;5GI<3(Z2&DF3CNV[@[D7D-GQ[T8gZbT6]O=@>:YE[:^^aXP\-#WHI]4PFQ
-NC/,(P;<=>FRC\NeJFU3Nef.=Y-HB.1ZQH7FT-I+)8_\M+_N8R_2]7Db.U@g_:d
b_bbAcY&HXRC+Y7@eH=J]bU5IN1+WL66g:,+=H7d?\@WH/:RM.QSbc2=M46#Z[RN
7+8:>CgYRKdHe1)Eg5G.X6/9fB_GFZ6]K_U[a3D)ALU9f]>QDR;P_8/LQ0&_S(Rb
<D^;)LTI=HLWPG/EASA>T4.QPaOPKg;MA?b[b4baW3,-P(D.<CY=GK<TVf+bH_91
d@>J#DeR[D3Z.Sb[Edg5/M2#X9SgSeSgD]D@2JZ(ZB_cQdTB;9/>a(Ig#>U89]5&
K>e,9@(J@Id/J4B7+-2A3aNU2=55IC8LZXc?1f[>HVPGeE;g<e6[;2148?J8F^5+
Ba+/S;_8f;X#g&0B+@V\.(0V7_X_\R@eN6PM>YWZ(LJ64@D-)AJcaMF&/JF,=LQO
N?SVI-4@5O]Wf/-^I_<fZ>==G83V&W(F3AE]KA0MNG2&C:&?fKFYNdPgZ_K,a+d1
44C;/;IG1U2I6#1ZV^DD6IE_JO3:?7,g^fJ]/fQ3CWEG,:(:?@-G<.?d32N)f)O\
?SeFV81aYW(,\1Pf9D(/4_abUe5P+dc4g?HR)8HQ8@_DE-^EaX\fQ<UaWdYL]Z&C
JHU-RY[&[4Y0U8\8WVg09#)5Qd3@8e#0[]0^5Uf)[f#Nf>>LI.?JT)E>J=g[-WL]
/4dac#CJgg(:2^0)+9K+MM4Yg7LOJZA@C<14\d7V=3Q>&_RUV=ceE8,IOBS#+2F@
8=^PcE,5L));0^4ee2RPDU[5OSD\Reb<bIf^Ya@bX^-cL2NDa\KT[H@L0;fP[C6,
AA_(Q2RS@;DCR9FA9_[)+-+G2^>XK=H134<f.8UH97\2Rg,5\dL7eET7VD]N]]O[
[YM]3D<07<.M&RfM1AI9TEcfLG[aIXS(AFI5KeF?)?ZG+<::36#/H+=<Zb9ReDJ<
E<H-AQXbe07-c89cAYLFHU03#f?Z11.\1B.DP^]U.J#R9K3D_HJb3)#D\C@YL/<8
1QR@QBCGBN//=@bd#J;Z^5eETKNK:D_F&?36;I)YX5Yg1dE?O@ZFVJF<)FS/+=d.
5[:+^A[<aPCP74:d1_cV(@c6D2^LMJ>S+IE0aW:HMAJLg^dXO8682B41?=#R6MLC
C_N4YGRc209GIMggYGE3)6O6,[Ia=13MJS>BX98<IK6Dg0T,Dg=#M<:O7)b]43#c
eK4(WZIB^.Q>dMR82Gb0:57TU.3V3?;aG[e/=TGSg:E:C=9AeGWI>VAR)+c(f6Ud
Rb,N4JRSaH/TSbcL2eeLGC7P_eR724^(Y[Z/b+(dfX+=PKa9>WeG6UI\Q5CEZd:Z
Q>eS9Ub]+2g+M6(X=TNL[B>aUf&9]?RfZ=^3&GMAHHQP05M[[UPC]+1R>d6<,PIY
2NEE[F6D?VHPJIXK)44SKT79PM7Ta.[XX/XD+(7Q<@&J;7a+aE[30UTW#]&AG8+-
)YK7FEX#)I,9<Fg[A@0>ZI[^2PLbWQW[bCX<>gUd<8G2d1R8Pf(QcWE+,_3&VAA+
0KG/aaTB8=)(T\E2+H@S0#f<R8&LF<PeQO_ANb<Xe8>1]-AQ#ZKc4X,f0]58S:@V
Z-95C7]1-]cRE@HQ]/96LAR@57NF)?(&3PV\,]Vg<&C+MJ(]5R6+6JcKJe.;C5FJ
;_-JRRb]L?LVJ9-P+1FS^>#Z;]<>DXR-EL?Qd&cZY<NYU8]e=PQ<I(AH]Sb7,Q;G
U9YXC2#<;#YdNIN@?SRY&0Na<XC5I_]NZ13OZfQZ(49>d<X)(X6[3Z5>:R-g;.8-
P[gKIE]4OZ5#eA0RO&:(g?c)T3&<cZdD2ZJ56W8Z7IM\b#_U1=1_+;;L&P1?K23g
M).A4DOfI@IBDRf^K@>e3688?9N,A1DF+acIBcd]bfGd00P:CHMR2MXS6+&@If>6
F6V@10;@JJNAaLT4WI7FYTV=+V9OddWNX=RX^:/-CRE:_)bGO\a8?253@VQ9I7)_
^5IeX-b&Bc<U?#/DSVWYd9_YY;JAFS;MEG6cYSdH#;]#,3]W0;EHH@HO4;^(;5C(
9_N5&A@1<I[e3OTKV(c8YD=8A:TYCIdPCS.NM-f7eG(BUVDc-UNVWR;Zgd&IH,,)
R3\4OI+8B+7>f1[6B<bXcH7VE0UB2Qa6YdVG7=c\Z_QK7IR)F&]K=+5(YE-5RIfX
V0+Ud(]cIAB)4Oe-UDY_T=Tb=#AYQWU#;_0:HbRM#<cKLDAMW^:PbD24CX:8GIgE
+d1[=2>aPLJ&7YSRb[CO3YA&:6MJ;[O6EVeW<T7IQ99)IP9^LL1NWTKN:S\)9)ON
52OZ?:)AWF4P^6#cO(D52Nb/23#.@bJ8JI-_?VXD7_?7gU)39RZ)[_==\,YN(2-1
62W0Q^A9bX^DcXH&R1VLU6eMb>[4WOZN-&8D=\9;\Z>095T\7V^++MM?KHWd9e:f
9E9:V5X<T.SKUD]Q-VWb=a+gW7)DcCK03_.1a#L.H5Pg94A^bD3R1VOEA.&>-274
I,+ZX)6)8R9d+C/_R\1?7U?6WX[SZ[b&NDa-GeDLb5\#U-)YM5:+],#]]PKCQ.fe
cEL=)@9UJQ7S;4H]&(FA)Gg4=c)>LQ+-Yc-4-.-3fcBI(>1URdO)aQd+OOMP9+Q9
H^3.,^N,3JSF,QHb;MMD;)&9gD2I(Re6(-SMQS&/6\E/M7aZRV1:dBcd[B,Ee9@4
e(3L)^R(I>\E#Q812[:4U+WIEDZ#gS^9=f=<&#RX73-:@[)5eVX50Q-TOGSV:,eD
9bW8)\>:;&D<T?bV.L:-d,a?ZY_8F><V:fa,3H^869G#N06X^X9d[;O<8D4BB-5Y
UN?ZSV]/>RJ[8Ja2E[c(bgMIRC9RaIF<)&]:>c#&L1Gd<.C@D4<6B]/Q=IfMRS6F
/5?&#O#:a^SQ2bKNUW86-/A+SS<>9F[&F=[#;AM^+)AQ66#YRX1bB=9E/gSA8L+E
Ne]UG[aR6M_\[VHAHSJ@RcZ)9D85+HH1Rc#W9M-VFD)(095G\>^:JK=)12VS,fH3
cH=?71M/ROcP@],W5?Q<;c@@FRO#/1b;GX6+D/dK.S]6P&W#A+@cF;6#S7e-.AGW
U1YD4_bDgaFBEN/TWMXY=CVe.e6Yc&Lg>e2TgM>0<WPA^,#QF<Z4ScU5@_+2<T\;
[OR1BB4YCBLX1/C@?.P.@E7^CW-ZP:0U;=g&V-Y_/TO9_6L_)GO>SM#UH5I?:LW7
6OGW1>W9aO_UaS3?/\b6JHFF]dH@;F])I-c/d-F:ZCWa/0]=SZJe7?eH#[HUZJ.6
:35[Rd=[2NbcQb402+.gS72>LL8g4)&X@Z?#I7\eFd9_#(UCf?d=\DONZWV/.egJ
R,&#@V;4H]KPOW#Kg5HTB)34SBCE58Y()Y(3e;7KHUAA_]b4H0&5:^Y5aNFSNa7W
G+#QPeHKf<2^=.JTcH)T#b]e.7JK_T\C9T1<5fMIY#;5;5RLTP6G99-WW5S?IS5Z
^B@@C=,:1R1:Y@a@^Q,+Z;A5fS@TG/OI+A+WTJ3@:bKLV3=G[>&^E5Kd51e(X,3V
aPFJWM48UA,S.45C3@fF(76/]C&C2U&,RcJVV9+D0@_(>Gf3#@9,ZL_M_THSBdgL
N+a86ZGD(J+?;6:3:e^NSac7>RHSdXSTeDaI1XEA1CV84WU_XCX^[=,4bT82Gf.<
JUd/-b^D^S49f58L0@G7.;E(XBYPSQ#&_U,>_JUF7g<;9Q^;JH^^]/V+^Nc=>(V?
F>P_^a/^[]9Ab7(JD?g)]a)_]fA0XG8+JfPUDbD=SA12<\H\CQ0LXf+/S]aQHPgZ
X4abD8-T:[=>a=FXPH[Lf,7^bN_d:N(gLX6VV@A<JJ7_X_<(:_f5N&Y?fQbT7MT/
7/O(EO?2X-\[e,J;I?3Z7bd?1^H9,:1/;+Qc>#N]^/E]C^:eVNCEJ93CbWeU)a4X
b:N295JKJI&d^KF:e[-;gY:PH3T#e=U#\+P[c&cD-:Z:-:Q)d);)5L]IX_+D[aRP
J9HU4#NJBLJC7JI\/\>_N0bX=?WHXKJdZ9=<Z+YVB:SC@_5<16aTV:7]@J[1;?g6
8KJ@U[0/1V&@;0da@5SUfE1.P77K^>)E0aR?gc)E&3WN=]E.4VP3+,A.[X27d?<A
M5-Yc=)LQZ<_A6]UB9f[.E<PcF[&deLB+1H.<bAZgL;W#9EZW+OZ,2Q9;;8U2QUL
6Z1d?RNVK@#ZX;31M,G5BZ/0-g&NO:FREb=8QNd@.e7Rd6#beb?A#KO&Y)Hga(7^
,TO15G:A01J45CP:_eG[SG@,:(&]ITbENXX_^]=@1BM3_K6M@3=;.ZISb^JVS3)G
,J(#\:(G@+FIaNTVL/U2.4XE?RC=#TB_OWcG/Ed@Ed?;Q2Yb+b9I><IO0#UK0+,g
HG:0-)5F),XN--3G=O9LOO3F4NMHR#3&F/MU5>3G-e,B\7#7U@ad8.SI[JJ_>cK.
f#ZR&W\J@<114VW._c2&B\/X:JE47fHdB>;=LQ&K9+6]40S4J?gL2)2Q]?f5^#N\
NW1G=O\AKO=g2Tg-BVGGIGF5;-:^0N75L/9=(9H(H&YDT<Z9PP^-ZGHLf-(@H46]
P1a2IgHVOYNa6.O[NGVPgFLVF(VOTa_.1+-GeH8?P:LOQ0_c]]FE,1BBV>c.T]43
B&4_a_Q08+8-/Y6MYQ[&aN81/6-(VW3ZaRDCYG]Nfa,FH>TEc(d1.RS3eM1Yda^7
CXEbU2O00?MS2):;c.K91ML6))^YcKV6Te],#[Z),aT3X#D>I/KVJ+J?R,@X=-;F
PK=.W-&@9[g@7=4aDNef#c))4C.:?:;H[f,0RgU+/)]gMM(S:H6G0]J#J273S2[V
:=QQ>5KFJ2=@OaT5]e7M/(.6L0fWgTPXRZV.f:9G85(/G]50JJ2WU8.a[T76>N<;
/:S(TPVC2aHdZ:C97L7X]YLBH#>-YFJ5NI2PV)+>CD)6Za[KA<E\=[JBe+IU?YcF
6IF9TaeM?e]>3HV7;GH3MHAZ1<2;;\RZ@F2[\V_G\\>#9)9V9+U(a/a^fEN&UIN,
E^aKQ8J@c3cY4O]P3e\&ESV>fPOfM=/^O5S6TM<(T13\ER5Zf:RP<2+&W@0=MKC]
-<Tb(9+B30WYI_]#T3e>1T6=ZQ0K@Gd?57a8Q\,I;A)Z:=&DIPP=7Pg<C,4b+05J
2RT1S-B<(-][^]10SZ<C]O]P54edM.]V-_c4(;B(W[PS:I:)8Na_c8@a)SNT._S>
PCE[++WSF+ST1c&#42U+SN7a/[V]#<GQLJ@Yc\C_Z+Y<BTC7)HWU_7+:]TgS,IW(
&IM<c,BFQ8V0M.ZT=G?MZ6^ZQ@(LFJA+NBP8[MAdESW>^@8Hf8E3eA<:/=._BNQ5
8VE6>gWd(a#Sd,\ND-U-a??,YcD?M)eVE[VS06,^.T3ae?64cLKC?KJ)Qa\K(0_N
SO56Og86B7=\TCX/_]C>E.0GP)^:C>5Q<.N[I4JNG/cH0NA5(#3TVHW2[^;?Ae<b
UH)S[Y,P/L9ed]=5g-:,Pgf[EIQGLQ/L?(ILYcD,R]>A=17g<8O\aA1:e:&3PUc&
28He?+H2Sf(EL_XN>.g(KFGgB_AYgW)fA7\g<.Z7@:aIN/MBM99b]G-W(<DRD5X;
7YUNaM+IPK3F0X?V1fd(1WCEe8H>CT6+/@/GZ[fM^9_DUBHVZF.YeAb(E+V].YTX
g,3bdJ<gTY#?0eN96@=DE_KL=T)Q,&(;M?OgJf6IGCVE@bIPAP)^@=A2BX7fc:3-
2(aA4@-^A4Re#N?VCA1=J/#-M1QE[cT2_,)gd,eI;^-&ZZ#0[P2<,1GA+A.4&cJK
((g4VL^/<#>dIUMcfIX\,?:H@B.bR119bS\F05G(KBHc]1L)QW?TW22dgKG_88AV
6=L=Z:M+D8@7=.8EYOC;=a;O#PZ<1f1RdS^R:MMW<RBK:90g>@&=3WgdSFDL0#,C
JdU2,Y5:F.AgdV9KGbNa9,\?WP/gVc2JEVT&D-1bO?&9aaW7SVBQKXD<]dJRM#IU
A>IPKT@=2ef=P7GZVRVO^];9:&1;6+,;/AECP1M/g(_6PW\I8H4A&EL0AY&Z4d#&
E@0(?C<?L/27/T&<_C0.Qd@B&(]LBT)NW69?<<H_>VZc7\DcF?:-b+H4aB[4Z<c8
FU?aD:[[NELI66];C4d\?SF^FZ227,<L>)@eD)Je76LP_40)cFK;6+b\)C68#ZbQ
Z_4=[-UIW6@=)g@WVBFS11&+,SNY;&7PWZ+6Z/a.Na,#IN:-Td==&+MbZ-H-/9E>
;TNO,Z&_>:d=8e:3.VE+1872<)R?e\/R3HbY-A@J,S#G88>/=O4I<.MY-RP1N4cP
NLP9>U0\8XEHA9P:dT2AR_dHJIZ#O+S\?VMb9&+T2OY@Id:/BfgLa25bDe4Og>FX
@^6JSeS0@<;V?BTENU+:MG5?Yc];O5Z#cQ-]/>[N_a_aBDLE.^gK-:TI/&cM#WYB
gddT@a7.GSPKMKS[eQD8\NUM2N:FHa^f:2BT<MT5=Xa1D/>5bU#H51FH,1GP)CZd
XG7bXU8=BX]/?C8PY&.GJd:gK6=QTT5V\RYHG;GK3L^4SW9BP(_3]bJ,+78QTPC=
I+QTME4EaHddd2I(.Y-1S4-aOBD?_D7Jg<YDS<?dB21d.RD7&O1VM@IYWBNCJXWW
?@/@cI.BNg^DC4.RW7,CUWPN=@=5EVa>Ye15AR6KW.QEB+08NBX8^7+Q\cZT]SP_
,JeB;GOG_.2gcW;0X?U3a5;874.D8[5M_F7H-N@_,,_3<56&RWL@70)Ab83Y==SV
7I8^D8Ra@1IUS#<JfQdW/e?V.+:Ee#75T59&Re>;b\IO5U)a<d.:^)&>@=dQ3<:G
RQL16/UN<D>9G(#L(-L4+N\@E6WWJ5;[/512M8CTU4>?fVM)L1-a=-[2+&e9)BPX
])+74-YL,H,DJE_27><5\,X+2Y9-30+gI:\Y-AJV8Q-W1N=c^7P)\MTH(d1d4aUO
36]SE]&Wc#7CHXX#gZ[V#BVM#MMEPM?G:72+?ZaWQ:HM_ca##N@_QY9d+L@66B\_
#_B\A&=].T-bgcP)]W3XUeXC@4cLL(0G;].W@6c\R=EHV83.RY99cYUS:[:[ZDKF
P1/5MQLfMB8DQ3MQPXe;PS689PfJcF+cIS502XYA)2M4<TP>U9Q#L;]#Pa#KAWNe
WM1QBNYX=eWA-U8=YN4PQ5b7OdIVD]J1(JSF<bc0+0OXTOB7N[Kc?)1a\aYD[3_G
aIMM-B42IcRO5U#-XK/9dJgHHdJ7-T1_X.(L?9E(IW:-B)O&9G7UI4e;@@6FfZXP
\[C#?,-W<P^97BFHR9^Z#BY6?P5N]9;Wc&1NAJ?)&MB0&R#,5?NAg[]A=ND5S(fV
N9_EM_=5N>W2W--0=YC0aT7@>MLX82HGN?YZ4^9(,7W:[-<7VJ1UaX:TW>CR7J;B
bb+>#eH(CS&c>UQO.2=f]E^I397EKEWgO1)K0@:(.CL)&,.d6]GK?BAH2>K]6M<[
d5,M_TH)EDVe:R6U[:Vfa/1+[GIOVQ=;e>(RI#F0AO9QXCLH@57L6AC/F=24?fZN
+eM;5Yg^Z\W?OVL#Z#\42A/67NGd2SZg/JSZ0Td2_:f2&F0045QX4OE[6c-gEU_e
)-V<(Y\:2B-;.Z;F,WJWU[[Y6O&bBQ[@LeFe)gF4e]PVY@fTg]A+^18MBa^X:_aP
SQI,0>Q.2^e5VY9+69W8=@A,<7+L]0@.5G=c80AE4D6Z+>.J?^+Y[4VUc=()YHVA
B&b;a2@?X];&JO-3M3RLfX:C^Y&WZ8#G5]5:5Y#-gM)[FLQ9eFY/cB-X6KN<4B<)
[M-eZ08S;H.WKAY.#fIZYX4Q8[1W>UF\<XG<0PWD2:McW9R&Yb1&(I?)-+2>+a@?
R9Bg6&M;FbA>/F_Q.e1eD,(.(Ld<b)#/\BZ[RSP.Cg?;:&P2TF0K)_IEH@6;3]+X
7,7^A;,Y//PG(dg_YF/5\E1N3A)+8[&gW\-.P<Q;>#Q=#Za,=X:O5\HME?@e)]WP
)-b3J9\fM7S^(Jf.V0ad6ed1>c2V:0F6d+LYe8^+RLg:#7a-,-]DaV[3SZXfdOIR
W\2Z^U+>B-f??B+RBB&Q<d=4RegRM[8S:bN:_FS[0#L)e8<?:c&PJ/N(N<>FDQ)S
GgWUXSV03^J=[6d0L.P0)E,:R;#EM/7^R5Q?BeIOBT:9XQV.\R@ZI=G44POgQROY
eRWC>ANW\5;<0/3M^_La0_T+bA.fS,V;4?D3M<gM:f/-Ig2_+&c@Ad47:-9N/MX6
:,[:EgY9A)7eZ6(VFGb0A?(Q/d^c5MJMfR(_P(L0WH-JVYSM1E)@6F[;>MK>T_/;
[71d)Cg^R@<:&6U(c5Ka+5QS7KRd[=CF1K/B5(/b?25<YJ5[a_SA[7#Db#a[>H<=
XQJIX/GfB[dRP@-.f=Af_\>A<5]CMC+DMKf4FIgBg1-//dOX+:_S:IH?./1FXb2Q
,L59T3N+^#?a8/.+a(K>7g/_;MeV9_83>91QBI]3aTJ&O4f&dA).e[PSIaWL&.Y9
(?>W1Q:+>R<54N4BYNUHLcRY7F[J1.U4eEUZQ6=LRN+S5,S;>)ga]/CLR(@[6,C0
A06MW,R5DDXWCP_3Z#a.^feEe-T(8.L@\@M/d&->)eIM_NS_EY1>1E6RD.78W95F
\J=)DfeGH]Ic.C2ge?&7RJ7[GB,WXP[Q\/gUS>N&ZSMN2,5=IL2^,[W(Z-d7<&/D
:LK+600#4/],Z+??HOUAG>d1M15Rc:bHQ],adOPF55#Q>-\]6>CUHY=Pa_/UgY;d
6?:R#=GX=eJCERZ76ZdZ8@:Se/=S:6QDQY]gHP7H0J?ZYG54_CJSAK4Q_AN8@#>4
FWcX?@eL^JJ(S5V\O/]-EXBG:AMb_&)70ZIQ;B17;#.+1UZR,W&U.I2.1,TXb]1(
DQ-J7==@Fff]Q,^CB^V2<FSD_^4(-7C?LCcPB6+IfXA;./&Q=[Uc5#Q#a_L9>OJG
+7(.E4/:Fc:,&;JY7GaCb>,5=_GOXDYYFJ(7YAAQ9RUV5C_NWKd)Z9M:)T)U8_5]
.g(=gOaXK6B,+N^XCEAfQ)+8]#MeH#,\D6+cPJ)6GA;8^WU_7a0Qdc>>)PZZ3I;H
R=Kg(:[OF&fM-,DZ&(>]a6=@=_(+OJL7;c>P#R6JYB12?&6cZ+:e168D+c-bWMHN
2b&:b9V0+1Y6=XDPME_M?F.KEZCAdfD&3a.6D@Q(O4\Ze3\F-3;WbGT#RE45/\V\
/];WeIT2=E\;>QLe2M2F9Xd]K9,.fc8-7b7W@2]8?P<W-?.B:TO4>#M0e@<E?:-V
;bSDe[@cN14URfg/5P9:YfHCCH[&+-5(d9,.5;3(<cT(I>LMe6T\_^LYg>e9(.UB
;5)fV#I_QLCJfe8d3IAW5W:L)Z,[eCLSe1D>cWFd[^b26/2UW^UF.L6SA2NW=>Eg
f.B;TRBeNE+\IRYZQF+:U@S\)Q:+GTDLUC,JP8KaXOY3?N5K_+3XfGc9&K(2:ER@
Od7X[L:#;IHF=<GFV?00D8J#T8N2=VRV,8[8c0Q0I_<GgCC@Ub,2Xe;?87-c@GFU
(8E^,4Og-R;feQ2_53J2dBS]4\M(Y<^DVAX8Od/(TI\+9^ZMP1e;E.cP2b[Z8>J3
6VX81S[9E3e1QXQ:231)cR/(<Z99=8^?^c9ISH1>400&@E4QaS,:F)_VJ6NVe_L_
^7+=Y,R-@^fYE/:/gA#N/TY9LORO=(:eXQJRXe)D?c1Q1>Fa>GaJQJ5=3PYY3;P3
5<@_IcE<6HXFTVCKe^\;7]Y96Y.6.T+MXEX;](<,@UX&:[2PWMN^=eDH9GX89@f@
1S5GNd[^8FMO?g=AgDS06aVC@LS)a_XJKYX7/ZY=87V>A86Z>VF]J^\S^5@1-eRF
2CH,KdF.g.Y<G@1YT,W9W36A?ZQ3<N2dA?7X:>QUWGOV_UQQL>4;T#aSW&C0cbAW
?U]#<U:,64_a9#<gF<F##Og4^CA\:Xc=IfCOYJ@.=Y(HQ,5a<+3<:]HZf3;e\S\=
\JEYVX-Ad1VfQ-_^d)0^;bF=&J4SFIZ)PZ8R1<([@3&3/E>FG7Z,0cO>07B5dF_b
A8\6O:^QcCXV_F/>V;SgWa_UG<eZ6-59@8#T<XF.]H3J>Z4e>LXHcQAL2MBPdTXW
D7b;8MZSAHV,>\(>L_4XL)PIVG[@^_I#a=+JX5AWG>7KRZ?L>\g51,6eKX[4+G59
0gfF()2Md=/6+KBT59N;.[cSL90LWA0&]W,YHHW1_U[b49La&XNU6\b]g>/6S?O6
E6N^S=\OU/^MH.7<\<8#(YS?Udc0&USBO-Z1d9#cgFA^K=f1G=JV]b/UWZ;2[aD^
Vdedf[^=LH0X-:E[]fF,\ULFDa>.MCgL>4SVg@S.(>-)WP-;L]@D28g\,AOCLV+#
H2)Vb3c80b#I\(H@6BW7PD1)gL3?3a-M^\0GB4B?N@KM3LVN934=abEBM+8dW,EJ
>UVeYQ+>))31bF]L>VFc\B,#d,SSHE+.-7O^TK(4-A)bb1LM/Y;K8(BJa-,;HCU7
J8(AQ5F7(3<?&=LaTGJdV=e4+fe<<<e7:R5UMC.3+84A0]M6gTDdH^.YPNQ02([G
_B5S9S5)(gN@.:>GQdVcG7VL/aE.04N[b#[8Y(@cJ#M4F9=7JA=XI2O3VN:+Keg]
K.=FCP?-c?bF0+6S0-d:3:\>J.ECK5&&=)H1M7H,8U-7\WdXZ=d,0[L6Y3HHWe9J
b\6.,&,=;W,F#g;?3.f=HA4d&@gGM];N3Fd;I=MW#fe:T2[8@K4&IAA=J+6:76H9
AD@35L1Za@M#G8bN8M<6A.8W.cZ\/MJ0aFeaUg\[c=+6G3cB#SD18?N@T+24N2,.
LcbN1&_NNeDJI?@g]3E>D9._d,LVdAdZ-/BM@5ab3Q14SRZVOS9Yc&AYd+Q6feA/
J>W8-e+.K[)7&GF,Q58BS6];\&0A8=5AEf\2TAc2,8H2LNO-9Of>-N)7M/N2IRJ^
,Tb=8KGP[b@?I?[[7f5bd03NB]J8?00[4?+KS4_XQOQEGc5&gcTR#GOW?7T.B^?_
:>OA?N\A,BJd(WEH4Z8A)XTZS--9)S@04N,X(9&4T-aGUG3IUC(:L:R27?RXFE:^
1O2-^e:0EOU.6UM=>[7[JW8S@N8(d:N_?cF@M8_HEA[@EPaQ4bD_FL?OQadbIgQV
@+K=([9-]S\J(:R^)Ya4]^9^XS7[(=9PELc=M)XPC7@^+7ZNVL?;V4@W?EF.L:<A
_Rd(Wa7P]>Q4/X?+1].S_2b,b>gN:8<4<A)&2>1L5+_9b[>-M57eQGF=JB6E^,W?
K9C^#,)A@U)gF#\[[J=VgHA0e\d^VECP=YOf>A];a#21UU(:8Ba<Y:N7^)C(U(=T
F_8N8>G=VecFF[4HCC:VZ-_bB>,T.1I4f.[c+QH,L4JR(H/8KTL6X(1;;[PJ?GC\
/I0@,G)ba=TGU]4(+Y],;;E-YbQJHW&KDecC2e5_JB>48_Z:&_BQP?DIU,F/K)O=
66bDTS7G,]QK#274F[8Q\MVHOPaV<cd-VT[95WRV6\bH)B29L^]BM-QPIggUeOZ1
UI#S:R?f)>cg1cAb<?9+RM;L&2ZMYO:]F767Gf(MBe7AHCDK?DS9[YKZgD=\VBGY
cA<&(89_3?H)/8>>DIN;10cG,KCEY&ce,U]+^&3#Ba?91,[^.N7g6;gKD5M[dRdT
cdAG?ba7+JB@[UP7E^4<UY)D/=3U@IB6gAeHQH@&QN-:1YPYec_]V9S7]:Cb6M;4
Kd?G=6fO>&=gO4_)R=QdHaMRFd8B2?3^42<fYGAKOaN:PL?A#S-aJY=PK(VZ+UAX
QIPB9<dHMW^H0AT7eK\JHY3X@SR-F==,J(&A0bP;51K\\/YgQdM/4<7.H40Qa_9-
1#@R)--7#Q/:d8UGAV1HL-Y2g3f<UNd#NZ75NbGe)G5N5H7>O]HFTF\@Z+f:GU)e
:(;1/P09U\F9+:##=B+U89^cZYRVMO9AE8MUZDVTCU@NJS]VZOFK)3MOcf]@Oc9Z
gW)CJa;.#Q?HcM^gH1P]Ic#[TO?>.aD(/F]IgS>>O5FF^N.#OGeD&U^/5[P=FN=(
5_^_,.b#a:Y]Z99g&-\W9M\Zg,4T#dXeZ(J/MKf-/[U0D<](>TQBf0;5T8VgcR9Z
JSB#>1W4E@)dcSJ/Y7U=9TX_C#9a=[&V_V)D#FS<+;/UeV6YPS&\C/J#J6^Y9AU,
8(RbP]d(IOUIAe5970Sg4AP^fV-a@B/ObS)V29f-NZHK1Z[SHR4DA1bGfaQT>XAU
</?(7ND<-b04?.<;O\P)S@9R)(CAbFX:#8-[389WS,@_Kg=<>\9L-SDaCU4K#<N<
T?(Tb49Q?TS=Bd>?.3R)N2]6eJb#3>>b[18V#_[ZYLW@KbUJ14=0&>5gQTL(0K1\
\W;1:?+61a69gM_g]8Ub4@?9>1,c&NI+]GGaf?A5JEX_#Rf,8YT3>TADK3G388<f
FHD7Te(FFMW?-S<9ZQ+]\PNgcVb,G&#]6aJR[_U4CeNO=#=QNHD_B:N^:IT]McA3
]BALAT35:HHaT#cUSU[Xgd:R19HY;^/&(8XG-8Y\@L<VS>a44S[?gM@Jc(Ubg/(D
T14eHOC8_dDDBYGDZ[Hb]5<4VOYL&M6#86[NP,A<N-VLUS40f.:^B<#02(4W.)7]
R(-0VPZ5L46/6]Z9-SV25N1SY);,O,WNI9@6<Oe[8[9:(fQF8:7]YPeP3.bG,F()
CB9-c.;M2H<d:J&JB_A[)gCJTV,31BV7<_C&7=1:V7eJeg\MR0CNZIDLdWOYTd+N
PXAJLNV&DUN(YQD592@?H.)90.RAU7Zb^1GJ]ZTT[>44,C_.R)F/.;<2[g9=dV75
JDYJ)4WV8N#S:,VD>IYF/\&?RT<?1OEQQ?M=#KC[L8TcEA=(KX(6MgaVRCAG80M3
T[5a+F(8EMaHK74.(3,O^Q5234e-Fa1_GHPCKC0PUGSWLMDCZ=_+)F@FATM]58/H
=P<Y(_E@dbU20a]3E;,[K>3@>(^K8OJR2LQa;5=F)8H5I?@cA.F9./J:99_e=^a7
,N.S93114@FW?.TMS@TKL>73I9]f90X1.Y9X(HQJMFAW:M6J<Z>LLSRU-_dg<\b3
H8=;/(^8F,=)B(#?#2YP3+2:DE8Zc-[>B/PNbSEfF^bfGRGIW&7&5(8d\:RdWe5_
@)KY,@8bDbL(<-/Q,a=_S:\AR5//\\@_V>VUVJ-Ud^^WO<dCK6DO<SR51F9+8DYa
TXME4@3>V;5I^3H\_g343CJ[1/#c5b;U,VN_6803e9Q.J6KKK@(-U0.NfN\TbZSe
#+BMV2>S_eDTH9O-V@(Eg>CdF,]B\?cSF\>DE4+>M2WEW-OY6KNWHP\8P\P3W3Q[
_K@c3_MP1]_5&?,@58+<&C/^b694V(O?+8[8L]I/4(dfN(T5PYL_(TV6,=3E\10H
[7>Hd<@_#MZSZ,c#N(1a(7=-bO=N]OPEEc,(WMX/5\QPC5[^89Q@cK&daU<>_Z\g
NAFPN5@E6>^.>,.349e[aMH-XLg<fPH,[QAR\f,]^AXVA^<WH1a/_S,(5:#]e26D
U9VC?<SW3PG,H5FL7[I8?&1EFMVTZF^.W.<1=AKB<8[:6OJIR[g>^,bfP3-6WCOZ
cN,O8NBDSQbe46V0_8[Y5-@&;LI7Se8UcIa421P]?8=,E@EI<YRQ(>:G)E5YPKf-
<8>E\94IT@c<^NPJEIL&M\#8aU@XW5a>[IJB4<eBE.2+dg(F6W]WbEb#?a,eDLCC
SNNSDX7cG<QF7^,BOAGR3^?/.5K3c1#.d0ND4T4\/PM//;NgR-b;YOffBIEH56[X
R-V/K:I#6:(E,6;JX.=\ZX(,R>YP.c.NQP@4())?;A,KUQ2QNDe(I8ZS4_AQPcEA
_6W[IAIea)ISc964VaKX@W/D?EGV;LP.W4.AM^);M0&g?C:-dfJfaG@B5d/bc3d8
ZDDJ?E(,B.JMC1-a[(##f5DNDIVP0>.>/HTa@(,>Nc&P/@V:_&\bOO<f8JgUe>_T
ZX(Q@RR3)FCK\eIdf0U:3QC&d1(OY,Y[4_R:gCBBG([M7QY30,2/7KWKAe_d#+g#
TL<Y?8<g+077COTOU/B[L>d=9PDIB;S^4>>)9bCOb>+NI3IQGTaOG[E\:/P/=dKQ
K[0I9VLS,9>&c=E)68:b[--4/0@\7BJ\4]DZ0ZIa.M-_@Qc5f1)T4e&V<cdP+#B=
O7PSa+Od@MJ074]YVQ/@UU&I5NK,,_+AaT@)2a70ceL^W;WJ6aLTL^1;;.2:d;IC
E+4XR/2a(\,<0W[?c858g1;]G9?0;I6,fZe]7RbRW\JUa[ICf#c@_70C:0)Ga;CT
[U0=#GX5OCG(3=N9Z_9A8;([+#9?,&6d_g[/5[Y6;Ugf-&-=:20BMcB-NOaT,QHT
D5FR=/9BMWd\:8fN=IW5?)B\FNS,55g[<YaY(:5:97;VI)B.OL:9&(T5Y<(Fa/Z5
c6)Lf4O\),cBYF<Pf=B8O&>;^N_?]NI=9>+.PM]ZG@SO61>K/QE^GE@N&fG@#7QX
2,2c5Jd6Q[5^@If2<H-(\bU[RL@^_G/;:TTIXN/FWe/QDAe:EO#;OGL+B[\=OdR1
]f<Wf<U508ZeT3b-JZR;N5d-OI+g2TVdRRbV\-d^b,c(F\LcKH4PLb23=;G@bUE(
bJDWP[fFBZa;LCQ2)N/D12;&Ug(MO<IKNAZF;>K3A4]MF8M,:GgW^=M/.Me2A,fA
>EF:=cdLWQQD1T&@fK>YPcU1[dX00WIgFMfP>O9[cFE@_FQ.;BOZ3+WGLXad>62G
F3S7G6BJ@/Z<>bZ+Af3dA<QA;-_^L1daGRTP[VbTG6KaFFbXN_9H@W#Z@E2&X+Ha
(@<gB[fZ=--HZXMPH7NgQ+Y/aeX5<.?U.C(ULL7SWM-]Lb9H-I]ffTULNDbeG(6e
1_MI\CfCZ&g&QCLHff3_2-ab@8Dc/Dc:cB-ce&U\.>:7e4K2YWcV4GY\F[=+1,cI
J(7;ad#>2FL8TRNP,3=Y6LCNGNdEFUS812X/6OP]0)(D-ZF],UJGWS4SQK?A_IH.
dZO16cN4Y7U=U+P>d.G97U[=EXW>T=I@ae+&BfPX:1\I.1VbTcf,>A)?S5+;GOXC
EATV2T,YDO4Hc>0;A>?X+9HA4N6/g?R)W)_Q&PV?=VIKF44[)GLRdL91:GE?\-<:
EbS-:Kab0f[R[g1&JRZHfAe^)FE7a[L0I(@>fB<<R-Z,CPd1b9L3XMZ]VEXa)T5P
N)[QJ]=#DH+@5bWc5KN:Hd/JPB:P+(4BeVWFCF^+SI15F4LU=_GU2Yab\BDO>Z6f
gf-\=?OgS5\I-TNI[<0;-G7)SEg(R+LG0,B5B;/GI(U6\JN-\0<C^\TIE>2_2ST[
dNSF0PQ/42L\-O-C>16+Gc9^F;REAQG1a+g5\41L/dIU9?+/#X^/GO^dLZeT(;_-
e,QF2\KXB+>HO[8Cfe?Y@J=C0L.WSMQJ_W=#e#b>gDCLQ[@P>=R[SBMZEKY@c?_;
66U34KWITdeg5Ye4Y3P#WJ&7@DL@)-061>F<ANAEP2H(P9Y=g(edR_=8I.=LgI;(
GSaJAQGNg&A:^gaFP7=&&<@MC-@BPG0@?7TK,L(IRCXU^PTWdYOM2YNQ:PD+JY_(
.OFL,0YU]I@#6MD[/\,/G0F.Tc(fXIHN7V&1dAC[^9G.WG^+<W:AF1-?UXg/dB>.
,FPS=[.BB\&CDQ4=E/4WP/9<<&LdK,XUONG>L<^=8.8fdb1WQJW,Y3TWdGPPA3=-
:bV+=(E20AaVd.HN]8J@f,B6,Z/N+4?E<d+e(D]RJR0Wg]X0/<B]dFUDC@6#CLXA
6VX-B3SaUbeB)U)aa2b=N<,^&(N)-6B8+0<EDd3cTN;N_546117+-E,TSAJW^1E8
C?9SeIC(3/G6THd7K-A@1a&--JO@ZYPIXZUICSYg(VF[U)_OVHS.#dA9@F:G#>/S
F=9.=_^X84NeYe[;.e:e#W-@SL708LDT2NXb+O2_d>>ZF?OV@DB[@JU#2KeDC.,P
LF#0N&)(d_-0<;=+Mb0DV?Z/H1)aODHF:SO9:[C/8aW1L[EB^<9\G2.=@EO)Q(-J
,G[D.+5)H5-e:5^+PLMWY#T2#UT875:[b-_(KT;b^,?_OEWK)E[\7(73I)ZGT8[<
2bG=MB\8.OVI@W)+TWD.#_B#5Ya-M-TBA)_\6?f@2CH,2[gEMH?:=I4#JWYVSfST
5V(0F6ZZ\(0YUHS(eQ>EHM0@OcP:d_f8A;KWM,(4Pa3>8QPZbA^#38L^T:<=-/[H
PeM.<4SK)8b1a-G80e:RXB)ggIF1PF0#IJ#4B#gN4/L&R_,9TGX6-PW+51KG)CP_
61/)V2b3=2B\]SV1=6+A-M,JCS;D_GG8cXeX<XU;GN:0RY4eFYS->DZVb(>.NX[=
/PW>1;Q;G.-=SI^AND5RT32=L.XaRMZS]MMg:_9A8eJ1Yd1I-SQ9-30Dg(/9fa3?
)X.e3JNA^<_F(d2NYN81ZBN_eFeA>]A7I\U/?0a)-X?<a<(PPSG#.H(CC(:SMfHc
9@ccQE2PJ[4J81LWT,#(6B3U)cbSUg(7?(6<96_a3>ZFe1>.Zd/dD78HYUT?NUY.
d+=12]X,?A8a(IBaa(X:?SX=,#b7B2.?#5(ZV/0e/ZHPFfBM2B]Z];GH@/ZKH]9X
LIb;0Q6LV[,4:9fK:(d51faL2FVK=<dc9_-&CW_g/=)CY;(+.U,)(HWON#M;V&L/
[R7\:IW::G^+PLd:PPMDL1g.P=@+]4[1(_dX&fHS#D:1gJbNd1C+)(87=E0U0QLX
.bgV.ce^0.N_IOY:Q9PCeSb,_,Za#gc>e7BVfJ_1?JE^Z(Pg\RNX4VSRSZaU.QAX
=dNP02ZZUZY:NUQGI<Lbf(7H[P:&-1<e1KWWT.V]B179a7;D_Og2a:EX1^W9@L40
7ePI7M3;a#(N?SGC&TaNdHF0F,D=]-VUYED[<cJb&:H\0H4e><Q4e(D^VdU2g2?Q
F:H-7F+e8>(Gc0-HW+R7+FQ7VKa#(S.Z[84@I.)3Agb)5QTc0S\=&BPP)a&8(9=+
[8)^24D-0\EfV;AC>>TJ;bHIPO6TXWG\V3(0>-XJPY3J68eI-I6;?JV_ZX45>=9M
MCaI>[Y&d^aM/WfX:.+\9OZ.+[bI?34.6==&4b</^5KHHbK:9;O-J#JH1S\Wd[?V
F1\0#Re[5.7,,\+BdM4Ta091-CNY;>C.AFV.c2,I^L/_OTL4#EWN>VG/TH=EX.ZR
=A;7fH7&F0@CKGf_d2^JFXJP@4(c]Z=(#EL?Y3,IXA0:((J+M4)2M]<)[?[X9#Z&
Z?AQ<ST[05?I)RAdALGYH2b)<g7d5/7B4TVg(/X>VF/P^=X^ZXS.F@?de1]1[PBY
ee4N@(O>b:6W]W9:C+;UAP;W,3f;8fK7-Z.CcE_aR?;P<dG,f>eISWJG7OXT\[>E
+QgXEI.16c&L\V-_-cD=(G7#ggU[8:]7SF?PII+SQSdQH@33;TZNO/>KGE#KQ=/Z
?&PbD@#+_YIDK;ggcE(E84-U/;<C\dVV>/O24bWRJa;DDacCWUL-;NMK+b7^-bCF
aP5A.Z#e);eP6)1>f,3CU11aPSU[FPZO0,F\F.HIfHU3DEJE>Bf@1FCH5VB+Lc:?
V()?dRbQS9&X@O,Pc+:5E(\_FG:3d]Z\a/65U/_GA8J=f/ZRO5\LKJY;AJc4UAA8
_g(cVYRO4HXb&+ge;_fSVC6OG^BD#7G_,2MK-)N.0A,^EgI3IUYBHT^efaLYM-3U
)CM;5T?1;A661gOFTQKENOS1D#9EIHd[ISSC#bHV3C]&(&W<L^6&D@UH]>U/b3:d
/W.EOJ/-T:fD6ON/Y733J1FR(OP/^(3=IY@g9;P[++_aT18_UN2?HG-a5=;]J/N;
0J4Cg1KXJ\_@+a1-^5Kgg8c?LHQGS4XDF=N#=P7Y[cQGWcdCI_eNL-SSHU&10A3+
FWWI,W@eaE:<+Wf4.][?./5F=(]\)7MWEZW)F4)f_V=\S^0GCbF9PP@ZW4LK3&1e
>W3G#d:RDVB98@A;W7NB/5[T7;;4OD\5HK@=.S/aDTY[JG5)U2;ZP]_d=]F?:I6e
C_4?=#L@9K&ACF#3c<cRHNQ?(YM3QTgAX-6X&U.V(J5GRa;Ya(AQ=22PI2YeaaaO
BU^FQ0IKVN)cK@cV[XI-H,_cC,_Z[@B7OTN)Q(\<;@g,0eM8-CYQ?R(D])SA(VPB
H,@G(Q-?\,;3--M,b]G2MXE;UM),Q]9W1RW0\BLH:;^0K_YVK4gYE(^B\(M[YE_>
XJ<,aFBEW75gT26\<[626BFd2&aSMSb>7O4<WY1>fHE-BH6a#3H4BGH/SSG^9ZSf
M&/fS7&Y+X_?W360F::6P7UXe9#R,V_72TRJ,S\E&.5O235Be>&b@_5\9J<.K1QE
Uc7H8#VN?;YLaS-9VJ<VA\C8B8>1+V8-9Y>.FI#^d_.d)7,,\Ae(GK22H@]5#L\A
D3C9aAW^;QMM6#T7?+U]66LN1fCESROTNc;K2bTS]Z(a\f[@:@SV#>&.fC5Sc=2U
&7;d#_Jf5f1V=@c/R0S:1M)a2QdGAa[AW6,a4,8+?X89[H<,D7)O/cO?1F6R64dL
0EP9&F<\@35V>H[H__F+CJ@e6@9XPIA0I?;YLYc?72]K_J9HH?QbPH7^GgIR\JFD
E&XEafX:)Gb_UbZAR-=_R/bd&C_bK1KbD-FYTdf),:@4@<d>CZD-O3.L1GM&PY:&
/fR4P]N9U_Q0TW?E)3^OcV8R:;U>]3>F^OXb>C\G,FI3MG<YIG/e&;NC?N4Q&?3f
WAA#SYHSJH:_Q@PbEA]^D=S+P/GOR)g//?.Y\Ha]Y5-B:X3cX6-)=X5KNYGXZ#_L
FRGR/=BcOAgAUBa38B^,/f]([DIFbXg023L2)3eK.P)6;QZX8ZU&AIc.+d_H)3:1
;b3MX0c1J;d+RUD@C?W]ab-?+1gd>HdZ,J,0Re:>L\(B&cEg5Q:H^QM\KNR>E@a:
11fEV6RGOc?90^16F^Q/,CMSeTTe/_A+D/1f1AVUdC//g?YdF1[XX#GMfO(N965d
#8W(>)SQQ\1[1WXYF__bPL+e>BGXFc)bZK80V/O[9(DFMPYRbDTdMfW0Z]/b(\](
Jc3f6;/8Fa18,.;OV,2\TZ5\GVbV2YdIR\B@IZNdRPF)N(5ggfOJFBOG>(18[MQ-
d[3]YE\7A0:K#<?d1CRdH\><gZMLTd?I^M@&2I55.KYM&9AE@.9#Pg0QDFbEe)@<
eAf>N5/R1&QYM9GA-5PVc>-@O25L<R1(CXX]PTYUVWAeOP.MPD1N(\#5We:&Ka3d
X2c\1E@C5b,:;eWg]2c55A0A:,UBX/aSa_b2W^^CcNJH>G;I:JSOTKUERb40W&Cc
aVD7g=g/0,4WJGBNU)],gQeW8Q=c#B^DR:6K-B;9SI(+5>/QG#)/L>8M2E7fQX-^
]^gRCeF]\A,LFO#Kg6W8O2Sc^6b.CXA+<&9Z7[N?,d6;#<BBK3Q6BaJ;[S_T)>;W
Rb9RBU/I]6f9[Uf>C?K,@N__G+URY1a=Ma0[@YAV[F2+egM0D]W&#T;Z+b.fe4UW
T^_7)CN\=T]_I:[O@+CHU,\;]MB[]+I.C9\2=).V&Z^8eK04cR\UK4IGR[,#:=]P
:_BIN.d.VHR2^X++e#L>-]T2:#>/[.U[4FCE&^5MT5b]K&Pdb_+MLWUHF3gcBga(
KfN3OT&Ee+<D+VeeSBTW<NTKbf4^8d,I^]YUaR#J0E6U/Z>3Y)^B7.Z^@#.<PL<9
aO:INg3GU<aPXJRZ^4:Y&)eA#Dg2XaN3XOG3<DFN+^SNOZfe]3QOI.+M0+3U)KbX
CC;8W:=J0;=1Z_=KHJ6]gS.CRbR0QIDT]>]W((fA,(>;a+>aB\:-_1+\@feP0HJg
>CED)6>EY:\<V/]W9]D(TYa0(VA(D1R&a:CZ+^X/RZ.H:0.I^WMG-LgQEUS(<)-O
O?R<[Sg[YX8)0.]TRKf/[G5X5B8e8&@FJBU0-?Ze(?QW;WMaD#F)HXN8?+G5U>U@
Q&U\G],\_:9Oe:Z^,ZA5KcX,c4/AeD9[g2g^-2<XM)AUJ@:S2IIBKd6LRY)[\&_[
.(dN:T-[@NTB1C?_K:a>XDOR&10KW-L=P(6&N0(>8<SHJT;J;;XcFbE.H++9Z-S)
\aa8aZA_6bSOCGd(^,K7WI=<LI3<)G/+H4GTG1Qg#0;-/X>A?HZ6232>_eB^LS<B
)\FBD=(RcP=?7A87KC/5[2?8-PgY<_E:^4Zag0AC:3cVA#:_5ae8<e688RMdJ3FE
-]^7)_L(D?SDUfDKRL-OgQZ.3@I1R5=9L4-;@O+T>R^OV@c8D^OeQ)7R)@=(=CTU
0Ff067/9W\&1C61R::(@3DSKP8NR/XH1^#X5fMEYIbESeZB#88=4W2&Y]M.>44(K
V_&>@UMT2P>TfMeRb+dC\cBX:5FPF3887RZMA;3;_JW-.&WO5d0:3^3P;460;-WJ
a3gSV=[3^\2e>7YK,P?622a92A3fb-R0Y)HU2+.R^UVC464,:9/;<9R\3.4ZTC4&
J>;YXSP:>P&[S?ROc/]cP\b86_XKF+-\._0UGa;6CH^DA:;.HL9/@aegJJ5aS(E^
LNZ;B7;64)\&g#Ng-S#O\D&aA-Pge??e78>c?>D1QL3];f=4@.=2bGba+1]+5DRN
X8BcR^B\7O70E/0QH0P(V:Be;L1D->0fODHC-a8f2b61BNH:Z.#S#FdS:.bIZ.Yg
OG+]5)RR1TfMX#@B5I0IWPAMZ&19CIQJT7#)B+MWH&CbIO/0SIKQe:)132CEcO)<
R>b8M<W2ZIH3A=K)3+aR4_QDN=IDC#)GP.]M9MX<c6[O3UgU@Qf(<.c9fHXPH)_C
7I@C:^ZEM.dSP_5\1g+^+P;JQ8WgENC2X-68d#RGB+=T+\F3Q:-5I/I#TC3EV=^+
W-36IW6@g2(ERQCe=^QTN,bWc^SG(B+3HW>;KP@-]Y2Y?I0d/VJJ0,aX(LU9,11^
\]FMX8R9VM>g4/A/bCT2cMO3#,C-2@2GU&FU;c/(,g>PfBNA)\ff1+M]71:2#,Y&
d\ID+B4Y]/WIG#DBg2R:6fV=AMf+F_-]\.a#(W#:I-2fbWb&^3Tg9O-]R@LT^Yg=
?;Nf40P27V13F[K27VaKbK[8=EU?WHJCB]+]<cS689=g:&.ab7.E5MPG>:W-_J8R
dU^E7S#c9N0S<GFK.YL,1LA^^AQ3DDS]?RLgMeX^I\0K]4KNNSZ&(I@9RUEaH\JS
)GK5=HRWDNb,O:6U0WAKTE]#^[0(:JI.(PH:DX76G\EDL@VTDB/.)R?Z#J&JSY2M
HBGE>9F915&KQYL-X6,gCDMOaf,;V[:f><V@SWgc\Q_:cF]5_gAL\Q]YVf>K1cDZ
QW)()CI0E),T]W0,BF>ZG3KY<GYJbf3O^-.,(_B]LH3gYA1F?da?K-+\a31.McVb
)5+?P=gMN2]UD11J>;K(;+IY&T@H64eXB1>S#2eFS+VO+a+15#a#?))/E&(I7EK[
OY_.4&D:1>/5I/g:\;8AVN=O9NeILAZM+B]eH1&U#b7;gOX@;J6@NQT/0KY2WZ3M
^>?]\4[/5&?^3)IP:S#ObR_X<TCESJR@BC-b5/,CZ8feL#9A/-8bS,<?_e<DX:BJ
,<@69L5A?3E4NacbC\E;B:SSO>##R;AC&Eb41d#\\4<S7;d#B)EDG@#:/:71(SKQ
.B3&bL2)<MRNfGV.BEV7eHL6V<OR1gbFH9@R0)7@[Lge:^9c/K_[PCb08V[#I+6_
d2+FFVPaZ&0e<dg64/VAaf533LcPbR754O:;T1a8CSNE\M<KE0NR_?-J:EK)\faQ
BM&YSc>@F&RP_NOTNNE2+;WNNR#DFbf);F_-f0N<I)R0]a[45dK,+R8JQH)JRH^@
_R(8S.>39)OT+WdEK]&b8eIYY>CZ7-<CeWQGMQ/.I[C)9ZHR5gG:9U#eMO>T6?RJ
bP?:We6FfAF&0).B+NTEB&D;#^2/?UKcMZI4g/CCg^Efd1CGCfH2-2[)Oe=Wa,IR
aY)6A:T]A8Y[5=(dd?ID=+KB#cb8^T)4e8CA-7\E9X?OY@?>CB8;gXCd#VP?:&SA
_)FMc625U62BJTcPbY&LD;>0<A-4GaW^P;T(g#<C:YYD8Y+fV?8OSKW_3:BU^/A4
5/baYN880=O)Q&G6FAH(M^@g@N&7K_+AI)HeLR+40\HZ4L;F^NU2#\2Z/M>C+@Y8
:D]K](HIIgDP-H06,I+^7F&]^V8c=V>I_WPV_8J,f>WUC^D>WbAY?8J,>9adUWE+
]8+Qg[JCBdRPbZP7H-G;\(a2bc:@_(CcAA[7O,aHcSD0DF22UPfFXI2-]:f_If//
gL5(2e0UQ@\5bYA._Ue^\,W)BNf]:g?+6c=2U>c<UBeAC5MVL0ZCBg4KK;g3L</a
JFI[#^2<FAV_Qe=)d;WXZE^Z04;3/8&=_dO?f2&-OeaR;]#X)=/I&MX/56;@CeGd
#,Of#.NN-d_XKe(VOKaVP0:T0b81g>bI(@Uc7WWCI@,WN(D[dH:&<O4NP;<9=/Z)
2,Ac71BX)WeOQAAR8_&1XK>\&EKL=)Ob&f)G+FT9_dV];Cg8;9A8;@4efaZ:4TU[
4CgGJOLXXE(=,9A9R.MFOg+d09B,8F5&C[&HJMOb5:.W(a1(geYQgfJA0/5gb=R5
TYWD&DB(cYaAdCc?/QTL@T.N_g1.R::&^OYR(##ND[GO__8EKY#Gg:3D@NT.-&\5
Sd,K<LY#8@\E,4:VWP(,:W#gb@DQ_S(I9ODbd;3F?IU1&/<T(F8&[e#-@JYS6e7@
gO2KSaNa(RQ(>AF9GVC/J9/fYEcc/XIYTVJT=K(@E#/<R^f;+])/A:P>BT#0K=&3
aHGX7TfXdPL0.@LQ).b<K>VSgYYNWaQ&L,]DH2M^L>R;<,UGa[\L4edHgXNEQ<_U
<44IbP,;8PaLHVI-B3Cbd;I?&];Y95ERM)Ta@/39^^X())&9]GcCA@[0d1P(?159
?954MN(PdO#eYRLe=5WHK;>_5Vf-dI_&V4,,;+6MSX__-#H\LfV#8WbT#XaL[5b7
3.PP7NQE=CG-9V:RR9R,YbIcO]6\HS-0@L-9H4>P]\;XeP<(W=C=1DcZY#2,K+K1
DAYVZII570T_I[e\):S:,[e6-)YW,2HEYd#NSG755O5/GI7>SY_e_-\[^16;Q,,P
,0(U50FRQ<=aI?2CLOX(a_KCBAQ2#HO1f4.3b2H&FCEe=M2FPbE?fb]^;9+8Q-(M
K([-[-Q3^2\DEOaUS69V;Kb/33eZ8J[dS/?_R_O_-e9J1d-A<dK1VFV[:g=Wf<AB
.OQfb9ba-X2Y=IE^5^4aRTC)B19Q.)c0KIeQ[Aa<NbS(8P_)3TTY:=EX]QMeOL=^
VB&XQGb?cO47MTK.;;],<Aa+>WeQ-@.#4C_G]H-V[O4dVYW,;RZB]HH,c<&,>Q8&
b[SUEW(QX(BAFV&KKec]OeB>T=dZ@gJEJdg?bX:A\)Z3-I#<LA#OAA-GV/LgK3bA
6JRM06V(<0UQ@RC?VS1QeL((V5IMEM+8Y1U5(aIMNXRcDN]SY?HZE+XPd-=/QC)G
J3FZ[ZX7+KW(8P+U?3&c9[c(#R#6c5]<40:?R-0PLORNFK\d\?FB1.ZIOWHfQ@F2
K1_HF<VWI9#/d?WX203KbD4/]H6)-5f5-4b,@I0],3CO6b_+LE0,69>FdZB2fZ./
-K^&&\_^e7N,_R]UJb=XB68L1f.LXKAeMV>09]IYKPeTZ(a5)LFJ@NQ<d:bKU6/?
&X_Y_3=g(I:Ed(6;0(>Z1BH^&T\-Y=(c#I778PO=a&=&LJQY8>DLO9HH5UecDL=P
4K6;-4NBcZH1-a^2ZB>:-FAg7EZ61/eZ.;ESG4\09^F0beee)?NCBTA[8@VI=d2J
eB0\TdMd6QE[+OYW)VMKO+H)VY>:\Mbb)be4<^[G-W]Ub]KeLB:VBXV<S&eYH,:)
X-(#MaI2??&+Z0HWIQ:5IVLLCHBAbgcD-)5N,<8)[=K:5R]S:=A1I(J>XfJHe?+2
dL2NaZ=GP_6SZR<1e,=DF,#X]6M_DUXBf[B1fPa@d=DP>^2Q0&9e:TdEL^DM>T>3
gEV<\78IBO(8-=V@PS9.?-TNWFM+0B/2:acOGLE)-9\EXJgd4DN#RO_SZEYb\DFE
^f]H>V:DB\UTRZJ>6d1IKG]R73?,]+bHfa.MHE+:G//4=NX3S_)39JeA^OS).Q7@
EQT@de:PfSIYf1K1L3Bc_9fSX[)[U(\?S1Hf5+)5M/ZeV^0:VXV,XW3a17U:HSb7
M7O]=_TOK-;0?Z>gABY6]9Q)H@>J1L99Ff-\6c8M^QK;RZAC->.T6#GQS7<5Z<>X
;4[./8.aP[fWYT8V1@02[272VF=^d#KbGWe5c2HXM7J5cRdY/S=eE;;1&WMd-(D;
C=S3N-fF:Od#A17[LK--BeG6cc3//RQ5IMd+8S+IU&P@V8bD;KJ4/dL0ggCg)8R@
,M:.DXbW6..R8gJGf4g:LS5LXF68Z>8_T0#JLfG&U,Z[T5XY#^1VG?GXQ\1L@<>=
/ec3;L[G9IIB#EN\>e+AW,H#2.E#Ne:0U^<G36aX(c?W-NFS:0d>gNdgWe4^E0gb
&GLM(LLNX#O\I/ON@a&f41X8QI8G5#K:#@]Q0P3--gHC5MN=fO9R@W)YB5TRF&Qe
PKA:1W>@LCSf^S[5bg?[(:YZ+gQ5f=1R/FMGF@7OMgU>B&>gT?-fUD6>AV.Y]MJO
,&c;cM\b/->:^U7U8HXY4eKML+.Bc_Ed<Id/][U?KL?N/V&K2)Y.:]<LEaR&2?F5
=fT-HNR6_&MTLDEcf>0SKV/6J7E:aEd8VT)P.FU<2V9SM9:H&gW2K6]?]d]DgeN#
5QO6=0^_;B\>fY>gUQUaGCWX-NaGA.-5Ggb#(TLa^b#QPef)42U_<E_Y^c#;5MY9
eVd?9,^^HS35)Z#aR;_.\N2V3EA<+423.>g?N8,-P7ULF6SR?R^PDL?M;QP,5)d1
f#1W7[2OV.B=HQ.:13/V<KgY@?I,bF.TJR0Z6QFVa^7QQNa3NYb#/TV^(&F4?QJa
N0H0Sa_HbA++JR_#.O=QQ;K@gd]V-R3(/ZCWS\TIZMK4bKMaD8YH6g,XNV)5KG/)
##ZefXFP:?#;ce7Tc/0)gMDXIIc@B0W2P/ME41_X(G5^;4\T]/U:bQ?[/GcX,;5O
fN[F1FaQGSEYcIXO4?AF-FPDBYKY,A086QG-M.-[/U&BfF#K9/<1MaP1bNBMH7_^
,H1-/,g7&\Vc6VF_4>D3,;L>Qbb4G_;a]>)1ad-P>11C7)EYZ^4_0b8fD;8GA.cX
U5<7QQO6+0\4M^3Z<DdIc6YREbT@GVC>1=<O\W4\IgXYDZ:O^b4A-YJ3H]@V2:R(
)>/;N+:Z.@KS2\7L@P,K8(3YXT,U7RDMRCQ&E>d;\J7B\H//3/7WW3N+8eCc.M]&
f_R+-]fNg#3L6Z#A[e4RU/;,)QZf@5#V^?-##b[)]DHK0MLaN,I<Q(/[C3Y?-5A+
F&VFD+@YF_>9PB_MOB67Ob)1\Wd-cgD#SQ)I=&_@ME2[WX_U@-RF,MCWNe\7Ye&T
_C\3IJP9cI8<(XZ[6@H9INc8F^JF0_f#@F4J^@5X2^A7)c]RR65&HO2U;M@8DUR8
Xc-@fYa)(_XfLRc(YE3GGR\7eY:4PF##O+QPQ\gKEW>)A5>1I:^T:&OZA[H+f,3W
\adQ@W(<6:=&@8MBCUc=63:R17J.g#bcBCMbS/L>42c>c@NI+/HRQE;HP:c4<J#R
GD]a&E_RKRL8dR).2ZcZPI-(1Eb?,S1DSQ(YC]CX>]T>L[A3;5LcX3[8/-T4H,S=
McD^e\S[7,VG8+T8-0KKJF:T;:ecF,b-0dI#&dG9V]d\M5SN&+,;AKJZ-F()CJM&
N:dE/Uf9J=&)9+S8.N<=U&+6(a(dX5DE9(X>8f+dfgQ^3(L2>.9OBRLS+XX&]<OL
KYXLP>C)<MRBf^/C#cBg_W-#Ia1e]d35FNV_#^IO1RXdQe0/-J3Gbdg6\?#eUfGG
@O96@E4/eYN8<N/_>Y=NBOb\B6gBbUL-0DL<?JT3+;8KNWIM:#66YA)eZ6>198YP
0MGD,WB<\TY#EE7FXF4a(H49O\DOXCgaC;Gb3A\,>2;c@V,T<GT#P#&O)5RI&dde
M?+FGYF)2++7.E@a(g.Z8/@:M9GFA2a6#\Sf>E6A(d,5@,N1\OY\&H6EHGP&[;Z_
ONH4aeJ4-A+:MQG+f]Xebc2[>)U-]W/56PL>B)79a?.:C5B53M)G<[N,9M4c9d]g
\5[]D/daOI8:PRQ7[0C;B:4a?YWPK5(RQT_a4X.+(gb+4U&T+4bPGD\_]aeQ9=Ae
8OKUgBE:LYea6?VO:Y,.e)9bXTY-QF4L&T/GI6J4/_S^Xb21[A-C5(Q]0-]K\G7#
=AF4bS-32Og_S^eeJgN]K0SUc6c=><S9TCf[3MJfJ.1TO>T)J0aG)g&@NfC]AN@I
ZNeb/^UCQ#[gGaK-FSb1X.F?Xg2,^+TFSCO=@P#DH;G].NZE<c&Ka[HDDG22MLTg
@9Za?I1P??H1;1gf4/0V.?XM<FJS[/b(9Q??Wd#61RdFYXc#BG+6bM1@:@WU),d2
@<.@^=&DEAe)<)+_R07@?f:d@YPGEfQT(8&TRSRW30M>;+5/(X,[0R>bbO@H\9-+
)IKYI/NVFGV@3g^XD\^Y2bKZ[@:SLV45O4<:(:K-@f1<59UNCcW^8\dHZQc&E7^e
Y]H6S42a;,4PG<-+Y_^P.\46=3[Gd(#S\dDHL,0D@748\HD>7>[/XBBcbK/;ff\0
M3K,X_BN6W?aXEZ3QFM4&[6Tb-9@&\eUH^E7ZT1J?_S6E2^GDV=OJ,<78MF&,9U8
8LENDcDY59D#8eX]W<5&/]1ZS8BN+FBZ9\?+B8V[e38[BEQW.4#[RI>PA4[S8;_J
?DD,GJaCeXFF\0Y/DgMBYY=ZJ\R5Kf=NI<NLebe,RgYKUFB;PaFDK<#^<cWe[:/Y
c_ddU^&<0g9)J&]Q?JAR2>=QXF\.D^=0cNC4^aW@2&gE3-C?C3VXb28>(f0e?#?_
[C,8c\E_Q2#M0CN4B/VGC0F3[PE17SdZb.T3T7:<g];5&CQ)e>KB]?@YJ0.4#/M^
WGbgAJ3E,K7@K/Q<R?E3Z8M+0MgLK/HU\(FS0U<:9,,L@IV@EME#S)754bcX#Pg[
d/A7]1gJ9J&)NVAF@ZMNEFFcXGB_7MgOX+<<88H#.I.BHD3e^EA+Y]E@a0MZ<AA8
\b-8?D\96eBI::1V/0=c(U/b#R\<.:9VF0(;(TgP//G6(8g.Q&7+e6RD\eXAgDFf
H8?)&TQQY=\I/#<[U-g#+]E/E.Z(657a<3/MPB+)9/1E,fB?UQ,Y;+1]<W==UM3&
)PPb.25DCG.E8SD0]gL)PDRG1K:<0b@D4PDgEcOTRU9HDB6eaJXEe@55ee,((<C:
J#J^60ORO:P48GUO]1/QfD_+^O\?A1N20UBfO(+[EYUe@JV4)\GR<=9KeLKWG)5K
;^@>b42MLE(]P)1(-I=6F/2/>,#g[eK3X@)GGQ>d1+03b6LR8N^5<bXDA]be9KA_
V+bXbQN3?CI+S5J6B\FV?d,c>bF[9@(SAc-35^?8)CXL.#G/-]EYSKgLWL@e./X#
#[KR7AX(\\&[K,CFMGM-C(QP::80>XN/2JH&AQfM+B,;&KA^;J>I/NX32[(746TK
(dW_7V^E4B-aZ#S&QS,_,>)e6D1;7FMM+X/#LgY@^Ue&AC916ZZK9?d9G@1&R]6)
_WHOHH6<+E_H(QGN&KCOI2a^52][-W@.F8=RNdMH9(/CgaX@Yd+&K+U2GP<J2:CQ
^8@Pa/U:TS^SKXLM?F^(:DVB:G;][^M_CPSV8.>8&&[8DBe1QOLJD(74[T,BdLCH
M2KR2^131J.N[7dPAX+4]EdXH0;XHAeT52AL)T^)Y0@J:R?_:58Z16(:OET6_R<?
8#YO[E\2@bKA_#\=R.8US;Y/^JY7;,d.Y718/Vd#-#.O.@ZF7c#72W-a5R1S2/-7
/e-UK.LP4.Y/g;#1HO=LVHe0GSb]6cgLXT?25YJZQXX9fCcRfUTcPd56[Ce_aY;B
5gHXXd7YNb&VQV;@g=TT?S]3WR[XXbHD=C4^fb#MA]g@1_8D5fVAL0M>dfJ)134Q
W;>FKJ)?9,1FRCPC,V=6@Je<IWW?V>[LYG+@FGF+JI3F/MS90)M<L(8QL?8SIa@+
NNd)>ARUg4Ag<B^bAZcH;+c73aR.A7#H=M-Q.b:dC=JIX:WF:IREL[)DBHC(Y2bC
B_/?e&+OM<\H6J<MH@O?g/#UcJ3DGMC@F&QKcY>IH/5YdQSCGIe3:(;.B<(OYDF:
SQ79B3IG#6TTW]<>gcG.9X;b27ZWCX:BcW[D0MJ\QS7K=HO;VY\HBd=?7&[(@Y4=
+4VR=G:ZG;&0M8;X2=1:1516>DE2CGON=W;JQ8d#RZS+Ge3?L@H;]O2DJ<RPD#B.
f(]NCBN,#DTRGb#L(\1/<7O[\VA=YU-1Bda]D&aD,IV]>R_P4WH5Q_2S>R=X(U=e
P8S1+2((3-B:Y;[aWHEGbU4[#IPe9OFFS@#7aL4_eQ6<(KX_eDWBaO2WZU?^)g8I
,C.Q2)RRKd.H:=[5F&PSe@8GE?>N)fgEVS1;c9[_>fb5F]NN][@P9.17fbd:b&]/
f[^B4-_AUJB>SB_Da&POIKceN?bYH.9:ZKUE?-.4&=a&B]e7_P29SO(OR=:AZ^dI
[DUY4F.]8IFQ=&c?QS].V#;.+4^K[KE>_4V1M35V5<_.DdSdcg,KS5=f59JJF^&>
O4;eEUgg(?N7:#G-^L7??W[KD\(=LR5@<cSa[]AHefPPZ(?dTYOF_QOWf7P./J9[
>55Z>(7A7G-=,FW/UYd?<L05F6TTH_>=@S#;M&ZA95QUGYL7aG7Z+PAO[\GZMFEX
S_EHFVGL1MP69/Se-a=]Ya44Z46a3_E+H(1KP\.e9]KdL,cSG)ZE[ZH@<1e6-/2d
2>O233SM)I<FZB[b_=gLbE.,-1C2TK6Y+,/Y.bQ<d23[dH?;X3,]]>e0d09C<V2R
5?..W(RadPcZWFG4WX8M&[X]PGE77,Nf[O#)-Y4.>FB9FU>gO&7\^@DZ0TW)EJ0S
CA0[0_cU03Pf/6dSPNXa<fYd(9<8&\OUP,e&eL@?M&\CSEN#+-U8G^@aa.Q3aV><
Z82RNI=7f8gATWa^UA-D,23-2GCBSAN7T@<aH8U2,]VLeL:EB-CKR.:-8dcNVQLd
Va600S#dcM[D#YFJ5SI.Oa9fNS&ZTL&&:ZC[ZB3]d/7.DWFD#[,07<#1Q_,X[;=R
Ue.:SE;S##1a&:0Xc9F.O3<+c,U?cOS@P=ICdgS>=IM@J)[)]N](3)X@NJ.CT:9G
[_S11eH_N,Ec&7QRCd#B3(4LBR[8MNVNF-I^\Eb^CIEF#CHLR7#EJJ&f##LD@0?E
Qa_[MA(W1PN.NN5,NJY=8)fWYT=5--21OO__JB<_1\YX\44b>[eB?8FK+RXTNBOG
cN-?e,/0HS5[-R(X/4/ADP30]/&22e5=:07NKN\.<X(F>]-K3XTMeQJC,DWGET/>
;T<Q[NQY0]ZVQCV]<7;#b6Z-1a>;7dXMR-=^=[eHc6LCIIY.e8TFA[A9?XK>ET,#
,CAN?LU+9+C,H.C+SL;I-YGgJEL<B=RfG>/ZPgLI.Ka15O[HG8YU/_>G[\NBG0IW
Z756MXAC9VM7[(aGV;?BMON:@#S8-H]9#fLRA2(a<AcILDD95KgS(dS33,J_<EAY
3e@:G0^[L=@M_U=U\P#TSL<6aC\f?b#?:S4-bJ#,XObGX5_R]D<)KecQXZC520#J
Q>D4IY^&<4Od>#c2:(?e5-S?.QJU&H@Y?:/#U^26_1[67RS4B-O\P+#\0cYPJZG[
@7@ab.3g+[P]SBbVB,:C9/3_P[3#[9M)S#c(.C?KH0>:Z:L].IB+H\Qb+RB&)?eR
VS-O-_AJYXK<ZTdI6KD>aX7(A/4\SUX1)8XRW&Kfd??TPbQ242ccO8XT6G)A>b8[
..e\4/CS8@6-A[IOO4B5R0\LG:;#aR48gYb45c4YO(+60N>,bCf>,^8V_V>M&N3&
X@,52e=U;##QGd\6;AT#WV<_Y&5F@.1.-,\(N)N\FQDVbQNMJ]&Gg^NQc)A.VR)2
4A>JLTAFDeIR6cG8&&W7LY3We]5W]cT>QPZ1@P/JM=BR#f[QZe(-<Zd_E9B2NV\&
U/BSW2:[aPZPCEVMNedg=@a/d)VBE@Q(.F77J?W+.GL8AdQIS?JO[5NODY@&X__W
>7eA&=/+c(O6&1XUP/ZZ3>cH>T.?<3;>8-O[V[8KJ.T?W#4/2E=0J,)\@CO;84GQ
>0;gA#f=6+E/L;a5-\WMbA\?<,+OQVdIY2,f:Z\UeY(bLJ#?7]S1Oe>)B/IKW)EF
4Yb]eCOW-L4e_[AfW+SA[<f]a47/5GYgHQZW?AX,_J16P,ECP6g=8#S=bG2GU]aC
#a6<.11W^ITE2Ld3DJe1AKDbF]IP[=#Je=e0a(L6W:0B/Y-/@V6_OZ,+;_JD<(g3
I(cg71&?+^_&G:\WGW_NTIWULT9(BOEg):\Q]7cb^2<]GRULA7SZ;D=_48<./+Z^
FQU1fOJIGAC0P)P//aH5VeI6/GcUES&^?O)SS8ER=#Vd4(P50_H73S?QR5SZ0W@<
ZeW9,T\-ER9/#K-I7M]eWL(C[L[^Kc6W-H#>1A<S3,81/?X\?@EPc)a>BX9<ZVVa
[9Z1X<7D[4G@(S+W#HSb60>.-Z;_C?-PDDG(]cN9;POg2?E/A69Gd2-3B/Ke[9@9
HE)Rd,8+W,^4;4XCDI4+9,LYSLO=<[0/NH<F>AY\.68_QafXD2.eUa@R^V=0Uf1a
UV9(gb\VgdH#+>#b/_K?NRg^I]Ug+ab<UggV\)Y&,<N_bYNP<N.g;&eY;:Z.e6Wf
:\ZRS=@)(W(O+:N9?aO.U2]WD=<c-_;?Y)43J9>0&WJY],&/-cA1/S3E)KAOB70,
#L2T3_I8&[@&:0=^)T]4M_H/M1AZI;PM.9U;P#47;f7O0<]>Z[^RWM-bC@8)E>)F
/QC\H9ZfMD)CX.H)-PS24F^2d<=&ELeQGSQN&\D]NB6gPL)XYG8/M6&)QTYb8I^c
F[c;@SW]\B,gC0D6Ve,\MWFM>T4O/Q>].cGABF1(U&2]_b:]@X5(?V7\91X&Y?eU
I>WbOYA])<MeO4.DOZF0UR++=?gE&/WHLBaJdDe.7EMME0/H7CYUKSc>#\1_RdZ3
26d8&U\ecRMZ19#DGZC3T)5OD)8c2&83;9#>?e73L91-W6(QQCU>:]=^d#=9fbdf
74A)aS1D@JR7VIS9>e<&8,02;>1+>6UcN^8(@UQB,PR7]=7#L2840#ZAcVfE+W]4
DCb8I;XW[@^JGO:C_IR[&LgWN-eQ)Oe\^:gc?SJN@ARgJA<)fNTAQ]:g:baUg5Cb
9TfU;JJ3K:G<XZ18a(.[P&M(>7(X5N9aN[eY4QK[[=9):gS^[A^:N>g372SAAbfL
QN.d9G]K/D[(Y&SCfX[/4XJ.G-A0N?Pb&#=?b3;AGO[F=Z>B6)K76/AJ@V\QYM52
a?5IH,YG-QFO6>aZ3#3#WAI^GFV8//=b-YQ.)e)g&20LAVSeY5;XUbO3I(G0K2RU
GIB#>^IIf_bbOMY(R48=T;(38(PVI74UB&G@K<QK^A_)W8/J8IUDbLQf+J<6^^XW
VY_X5#?VV3F_fKNLKc+P64.,^^]Z[;_8F(2K-Q#c(\T><-+4NfO<fa;#TPcNGYVZ
X40C:#=PH3H(&J)][D2QCeFN\36/N1+S=@EU55V6K^2\-HWE;P9d)-+0XE^2:M0S
/]EaJBR2(C+FKDT\_-(,H1a?]@+&9[F_S+]>)5Y.fSOQY8@YNf?F0QUO\EU)?0+R
^_G:K=T[\B8,W6P2Ba.=3/WY<b(eH[?^_dP[HX?08L?S9aT\gS<3R>L22dV?#+-e
&3g1D480V1b#)N-2#09V-,9&;]S<XT>S,\(Bf&U/MZOU#8A#Z@[<cf+)Df&Za#9D
4+EF]2XD([2g(a8I4M1BSf>T-cI(gGPYGZBc+Q.Z+_NT>D7f-gBUKKW_)b6+fHS2
d=4#;H9g063-Y-TE>FOZ=ZU\;5JMPRU^4?d3(BK&F#7-.17#8#-\S2BfZ94&/=f@
#/S_QRD+2@UOJ[9ZNA6eQB<>T>6g,JTEU#^>D@[4YRVfI))afZVGSYE^?Z=BAFBA
LJ\-f:)=>T0:K@?61Xa.P24_^bBFRZBcgc?14aZZ:^/7D0&SGNPAL=:Hbe>EaKPH
b1S3A#CV1:;M8)1Nc>Q7PN)06D\(1/NDeY]7e^@<Xg5KH@OYOTB:;<g;HN:ObfJ3
7WATMD1]A:FVaQLd(HKd^c-eD^\\1XF5c#.O<.Z5L,S+;&][EdO.1>gEd3R0YFDS
NgRGPMe^NLH3?0I:J(NeE+.CeXIB:2P=6DZ?Q[HeEgH,;cBKX==(G)+GSX4MIEV[
[egZ=M7CA)b.ZIB0WLV&U_BC765?V>Pg.MBL6]743P-N_bN/e\_9_M@(Iea-1a^(
]L4]GJ@&M>J\,-?Ja9bJN2BZ5f0P>/^4/OP:CI890:TRaED/?=e<K[6RUO/)_MWI
5XE))BX@3#5<BSX09TKHb6@4>2NIf5/[89ZDbMCXOVF.3V.>)I]FZ(A@6KK7>Nb<
^1BVJ9b@@_LWPO[dXMc^J+/?M^[31;G71IG+S1&Ed@Z9&8/LG]FSEG)5BO#UFgOc
HMS>>CYg#]geg5CN_Y&8SOW-fc(1OSGQVYF6\6(=1;I[MF3e[D6/;7ecRDY71Af3
HPf999<:WFZ>g8&8=,LC9<HSZ;)HK6]SP>Cf4#9UAV)Wd<O.PXc^0&fE.6TO]>5F
P7G)0f)K[8^XDcU<Gd>Jcb^\O-RHagTD&MSSJZP?O)b?T5F/2a(5N0IDH3NGKT^g
,J98Y.R\FD.V&.TZO#D5ORRTbVY@.W3WW<5KARGT7dZe@(Q9UN.AN+1N@?/a>4E^
#:A3BZ9N1MJXA+_2ebNOB^:_S6GR075XT9eHT&MKXPSAL)7a+)S2:Ga9?L++3dH1
5:&C9]9B[7ZC&2;JFDH\Y_d:aHfBA)&PK+Z:H/^<2=\]BMb1BRcZ[Ue0B0[G_gN9
F(N>McOFSKCS^[?@TDOd&M)@6W39]bg?@S-2#K,X-LW;Q8FT&+(^H^dTeM&be&H3
G.a6RA,P@He:ZOHXHK[b9-EM2/ZRX885(3+99;YRB/Vd+2#5NcFS8aJ0f].NCR.F
[gO]-bMQH+agc#DB@eALQ#GL9Q,#+Ia)@FI1^3[#V[E,&]<C=?9UJ8P?OQ\5S)gG
I+K9_aM/916[=b^28SUUZ9GH-O]DO[1_WTEX)3dSA^R<c2Df,d)#OOad[X5&C,:(
;P]Q>7LFfU8B@@;Q^7U@&3315JDJI-4@K5QcPd6.cJ,?]./FHK):>U0;eeO2Zd)a
6OZ2_[082gg;@&PTC^2+19Qba@00.d54O)eAF@[3^]6g1da^T)gY4XZ6b#E><@6J
f38SH<-,G[\U3&eI@?6M2eL_3J,f._:0Tdb9)DId09GI#IgNMRI[+.NGBQ?>.U3\
M&UT_8T&3N1aSZ&JCKA73;6M/gcgc#Gb6Ta]=geg<d6V#_M.?.TOQQ((CQUO=e6V
CC;&AH;(&Z:X>(LK]R7c40U/Vd,3+C,CZ4\\ae0KJWQJB9_>=?H[Q/SeB,<:@c_]
&R>O=X>-Oc.fLa9G[5GS_SJ^6C7AW54YD&Z,A6aI[OfGJ6bP3e7F8@>Ec)C:>H7(
UCJN@@NN]fVYV-K^a\Y\7-f?B,Z+#^U1.9;\8;bF1_TR?MgJQaP:@L&^(VYP5(S0
fc]TO@1T<SWZ.EP0aSZ,^46H7c76-N3=bJaU3a/Z]YC[[98+N?K-a#9IT&?M]&=R
J2.7ZF;=,D>b\-FAJc53c?R:_9-UO9g&(ZSWG4IU&J\2M([H<X1TbAd?9=5U9f4f
\R41=L#O2Q@(&56F-bWNd.K^eT,LKZa;.XbH4+)R3I3>SMgC_V^4g.5P9(DRP,)O
]#MC(=+MP2eW&[Z1V]5JXf4MbTbF9@VGd6#/FK0SOB6K-6?HE7L93.P5g0H72@_N
_QSJaI_#BC=VcY?0ND32^>b4(Lg2#DHEOfePI5L3;DCVVI8RA8O81E?PW<Cg>V.8
HI:VMfeDfJCGa@@<A1X/LT<3S0JZ0)c[NIA4&5??RLWOMUP.O4&I2JP&MIdKK/2_
#?eAU1P+31YEba8#&,d&(.70AZ6\>U;[fgN<8[?bVTS#5#BN=)1?7<FR43L;<e7S
_(I3THa8PfY#?e[.ae4VN&G^E3K.Bg^5EgI9(Q[@W.N,NM<K344.Y-3P\+aO7><g
F;[N+E3<aae3./cM-69Hb+1X(Z(]K0=+=K2>&DLB0KW0:?=1b7OaIB+40g?ZOf,(
6gCQDHeg@g4I&@?>^bJP][9^TBQ4[cRR#O<;FM)5^U)8/4=LN;3/:ESNA2>F\,\@
JK5FXdeWgCEPf]QN_N:K,W=a:dWO92M.63e5d2J0)K<e?bZAXIQU#?QLE+KdG63/
g:C9LD-TR:b;Gd>3_ZP<Q-,:XVeRB48@TgeO&OEHVY_YQR9PD(P1;eLfDe>6g34X
=0Ka#5If_VDHEfT/V.R>+g(cX4FBH@cP\BWXc8IT/.\V_LK]JM-MPL3<&>HTgb1N
CXTca(dX/^OQML=[4[\V6,<^cYD7(T=0,W1\Ja[E#E]54VF,@fD0ab?I+>98T=PL
PXcBbU.8>&[J+F4>6ZCBcH>\8&SVQ3LE21(:RZdUe<BYd&\6f_\.XVTA\4_X)/YH
<JNf2Cg?^28<gNg-/LUA<S7HJaY;:^@1QB8[P]_J?=F[HM#BCK_D,-LK+,8,;/dN
B8B7Z+Z)<-:^G@fW?F[,Zf1Y6e9:2/1:.@CL81)#^<A)Z<gDW+GUPg,GKF?GM2^K
gC&)KMHBHG_W.I:]73_/T\aI:C.=6[V6NT=c@F(YFL(O0Z\LH.-K]g.7[VK-1>,(
g12/U@a=1:)YVNS2FZe(91.:8&YXZD9aS:W11HEN;V?ZW\<(MBL&=-M_.bV54XTY
O;f7LK?5L[B/c=T^LAA_dA\GZ-6R#E=EeOM\:VOI^)H?CU-D_>GHgL,e0A79BWL^
K<b0dLWX-I2HIVGRKMRS-Q9NG-Pb8[O_]4^2]-[TAV?4S)5bN\+?d^Pcd,2aVc0H
9_5bT1.BbV+TMWYAfND3Z(<5dOXDcAM#F<0->#bbG-:8X;H>a,/A2QR[=&1\cJD\
,2H]QfPaIB\CS5,N[1R(=</]?F0@ca5EdQPII80aWg#COV9SILB7[-QP/R;I50]K
Z@;C_UeH)K1[]OUXQMM9?C\ZL)b+TV>D2=NEQHV6C(2f<,XO_Y_;d)6eaAA7,@TP
g_fJ3JPaO,GHR7Z_b2:<BGVGD(=,8TYMC-Q@LRP@#\[4L=E-_ZJIKH5_44X6+8#U
JZF=H[fYQ,K&ZCQDM4WM)DG9f\bX4=CP7b6Xb^&G[HYV87M7XQGV:>]f)XYg<60K
]RL9DOPA[0Q;f=,6gES^>N:#+&a2=4)?7L#\G&X4^4?QgBU[Te,Z=8+Kafe,ROV[
^c\4S29.ZS2\.GIEWQ3:L4YM_f)0I-@9Ze3f0D@XG&\36RER@;efM)R_TQ4C;WFb
,O14:Hd-@SUYG/=f--3J2gG::?+0>BMdGdEG&@]\0#LYV,]/_(V?LHb+_>8G8U_5
PN:X08&@4)(<d/:D>+b0Wb;-gGP,[EFKf^2Jd#8X21^[>gY5/61RR;X.I2R+AMgZ
g79)2PM2Zg6LPb4[H:FV5]MJE.>G\,+(5_:WJ1JI4/.De2ccAIf=T:TF;E04eQ#5
aU5K1Q,3F/E<-4c5B65SSeKJ1SJA;c/a2:Y]Ia5/RL[feW#]0#51<0)VE-#_#X&Q
XR4PD\C+[4\fO+4b##P8\##@<,<4^H2HWD8QNEJM-IZ_@KP[FD.GZ:FL/B)?(X52
D>512P_^g^7Rd.JMF]AMJF@F4f0NG^O?O;=-+<\1L<BdLX.L^UP7O]E:8WVOc<)+
=ZH5@I8EHYZ,7@VeI5[KC886gZ4&\/9UX-?A<fBeD^MN\UN:D+NCIC.5Mb#e^b1K
;&+Nb]\WS4[bb/U0R[V15:/B\,BB#2e)Xd/=D#4K?E\QXUd]g7W]W^FVJIL#H)?H
<I@Y_E)-b^)HGdBeBgA>F#:0Q.dLCVdD&38,P0<L6FYf-WBFB&N/Sd18Q^:15?]d
[NZB03bS<26-PN?a/9[T^(GS>-EUPCf:3dS0V@:46B=A7M9J4N=-@6,BS;3b(:=L
?>+cO(=8]cXed=1-[?]\_#F+N#_GSJJ69J=T,>/>WEE=3(UCJVWCYPC_ETB]X[??
_:cTa[4[]d4;;<3;RgL:2Pe:SYb#<D^7,=e<;6=5^,8\5KRH<:&,<eVN[?@I++=:
@(SS[)Y6I7a6)S?_17a,R2G;C)2[1Rd.L1:XC)e@-<.\[cVP59)#JP/G.SQ@S/M)
55TeX.:6R:.XXO/)?.ZKdN<L_[OQEXIN>[3\D2&5AVE93]BTA@OL#]M[YYCe5We+
:Z)f:<B;7Q:<SJ)8,N)).Y38JG7B\6@7LO:OPLa<@a\0(QDf)S3K2WM,1a5g&[cL
d_1D?12A1/\T6<0/)]EOUQ(M1g&>,B7^TaP_#,EE#E(<L4K#?:V4O,:FCAIP2gYV
9G46T@3)D_c[9K8CA2X9OB6&\V.eGQ+H0GMVS_EUL&<DM]RF.AABd,PR8H0QQd8X
0.#)PVDD36=6KP0BO<d\-ZK3d)a-Q-5-]aTLZec2Y0OF<-DVU]0\-T4&O&-2g.g]
GLK[=66)W1IQLNGfF/NZ\#S<dGd5R4gd4][JZTReVZ.[E[Fb(?UGX4W^Z\EF@ZY\
(+?UcaEd#-.Y[<QAQR2GQFCXIgEKafN0TT1M&M>(Y#G<acZ82F/Df0A0.E.[Q[H]
]8Q[#<Y7d0MQNR7PL(+8a/KXR(.d&E#1QNB+#R,BJ_194;P4@0NRO&G+JG7W=H30
gCNUgVOF3/2QO@C9MNVXb:RK)/W1;;(ZV8>A02Jg)g7/b;YdX[Q2]-_M_6N\bc;F
S4LFKf[0<g4I3S\[+&2a<cTNP4bOBU7bCR\#FFAbA<c.>SfQ14fg5\S98D4FZ0J]
@A7Na@[0>W1@N@;C=ED.Kgd68E\X(=#0gK_59Y2<6A.Ae+_UCH&E+R/-fWO_5(ZR
5S8W93=b7_gJ&_L;X,S+NCfZZc#AUG,1G>N9]9K3Q&GC,H+30Y4N5<&ROFC[J01^
d_(c+5^(>><_:8.\+#W:R31gYXFC;FOBW@K[2QGV&MN8_RM2UD;89c=F(Sc1<S?f
Y[\.a4EfV;8=NRKBeb&Q_);\>JIIcagc1g9\8\XW#>1XbVd<_,EEN8-SgCU>L-#>
Y1F9FK<VO9JL78)7Te-?O6G>:X[B]9N6N2+P5Y0[IC1SBYd615Z@N5L,9BaKJ[OU
S;TF(EcZg,KYc#@U-P/DN2Y[@MN&4HfS(^9CgXXYP>1>SD?Y?Z/I,/@]UgI</VVS
=b(Q.97FD#gYA;e46N:1SK/SU\2A7+a]E=,2b=_7.,d;5UTf#C&#KS;eHe0&EVV,
<VDH3PB8O4R31IY.gCB2aA>#FJ,gH]^.52DW2#aHc^#9<&-F:[T.Iag5?O7,V7K?
cZA,0e]&T,;,X;BddZP0&],QL@g=T49cd1I_Nfg+6QSI7[0cQEEU;e6#(M89D2+E
)6aXH^/?_f=4eEeXTB7f+\VZ1g3eWRG#VVSWCD4dC\^YF.Tc7._E-SC?^C)#e7NQ
0+0-/@Q4?8GUHISfJ.RgSE[AC;1J8a4D/ZDP[7:^GM@a&.?CPZB;_3;aE[KS#BC9
GMg3/a9eEgT_Yae-fEI4.@4WNfNb;f18YAZD3GC4&JFK-cHTVPA:/A+7^M:WY_(A
(CU<4@??QP-gT+&\=A>/Wc.dd+8BXT^K0(TaBU,0Q9H-51g-6P^CCU29RCBYdASa
:[g)+AJ>8f)_[dN98[dTcbQ#DEZV>Q8Q?bH+US#>ebS_bL3VBNAO:TdEIeZ7,05]
8O+<H<30RCaYN48=bUNX#I7Nd3D=?UQHf<)9SFP]?c7d^Q+5+Mdf2^,UQSI3X2YM
c>Z-R&R=R2Q:UY\MJQ6S8NaWG[-R-?fbA\=0ZPS3IY:54;eR_3__AN?UdJ8EN]=a
B^WgY[gbVa?\Ld+?_S771UUbADdd?POV;McZ_gT=,ac36&]?-(,fTKEeJN7@7ZUH
MCTVJ.W?MY_PFJ^&K8a3C)#<5]S5D<b5N8[/#KTc70?PT(04E=K.\2)4WDed?PVQ
A6WE1S#,E?[P09gKR\dY(8_Y0B<Og=G\3e_W]4d9Z(.=M.c.T2-L];;:E=aS(RS2
RG03(+Q<(ef@1\,P)e,</EKe7BUC1=UZ9Kb/>bH8EV=)TNT^+@bE;D+>@4cNA6?_
LbL6YWG7g/\IYZf^&b:(.KC,;7<XKJXZAG34YL=EO9dPZX[Vbfb6dRcVU+\@S@M0
6HeU8C/6N+;G#]KK=QaHC,fK8<8<7:KRT#YYQ\8R3-JbE0I5+RM<2B58c@7fY(SN
Vg7G7Y0FV6I0ObJ.C0S4P-TH&?N[Y311NYeTFHC8R?9:6g.RZJ2F2-<Tgg-3b5V[
5(Ag4<:B7UCbIUB3_a\FD)5N?#GA)5K51A)C4A[6<:e.@BJYGd<B@?D=<Pg:MJ)<
;:K;<2c[1EH.;_.8BA/T+2YS1X+;N09=N?<V\VbT>?E-C8O:[3G1T+(7DPTFIIFR
YaC(7CL<)_EN<O\ZI(688B]B5[LN@_RK#3K)TX2b4YaI@QCJ31Lc3D@,+2KdHQRG
If)O/YX@4N-&Y+B;?R9Vb==PIB,0+c8Sa+g58VM5ddRf2X#/>YWY?]VBM;,YE[9&
?4P<]B6?3c0dHQ0a\,Fg9c??G0AK..HPA_Z;V68GVPbI-;(?JAb;))?7&#WbM?Y5
T>DbAgLZ[O3F5#L<f=WSR7L8LW4]EQ=dH=LH#Y(O+;)OaS8D-NN,H.7T,CES+364
EE2=HbEO6FL=C,8S0[LT[1N2H^3<]gZXS\K&XUE\+^)?_H[cS0ePSgQ;Y/dSL00[
&J>Wc-S=OBNYf2S;MOS<]PVCFaW#NaQU,AD^=a4)=f+@.UJ(O4AJT/Oe[NI(:ZY/
aaT#3;BO.eXGOFXTb<#+/_N>APL6WA/[MUga;V)0JV@<68;^37OW^McgYO7:KPJ3
Pa9TD[J0U:<5<_)aN>;cR6OS^N,I4Y65DeH<=&P]+VL94@MA_D]e)ac[^HR2E>,D
<gIVUDK]d1-WadHSDDPe3,5-.H)DM;\c-7PbBN&/0MK;O^RJ0a+/f7LO/1P5>Ic2
1J+)Z40e1L?(eJb-9F[EX.eJbWU)6;5EK:788R\J/:F>8,G#XaKU(Ia/bXBQ1FQd
+>;b\B0?_7fCa_;GB-,WMMQ6&RD(\-<W=/IDK_3^/60Pg)(g9Aa-e\\Lba6P)C_Z
(X979^FB4Z.R;1HA3ATT-T9D(=Q3LD.cd94?UbC3Z9\D;^DG9E&-Q[#bMd<D-8b^
T0:-+9SHe:HNBc=);W46>[S,\=N/W,CEIJV+-<G@P((X._JPLR.DF70JCBIc:C5&
_TdQS,F#)EV8XS5X#]M/FC5(C^.db;,c-3((^Q_?eR42:\.R&-5I)Y<8<YY<Bc+<
Bb7#79_H62G5C#Z,>FQ_=PG3_:g+8G&:be9,@L[/1aW=V@6UaA7D_eZP9aCNN#;/
ReB#dg,=VT?GEAe-Zf4N::^+#d;54TcUA<Ig<,4UXdg),4>2PPNN]9T\#f<cFZAY
Q^H^\?548cXgSQB]/BG[DYY@0f?UU=-=YAd[_UA<TJFb:4_.Y+(5fWMd3@(\+V^/
<G>6)K^07BUPM\b\=QUSA:QG9F+<R<D)U^K;eA>2c;I)-&:H_)bH.a+^FH9-R^))
;=>(\K6W[PDDc\:K^IPg0@Z/I94:?E@HIY1N@:dIeS95;7&B0T+SMP?Q[1C1R)EH
W5SYd<.D.SbG;YdRAFD4FRa\W82=C;]K;C1+KeBEgRQ0aLAO64IBagPXIS58BdY=
U?)YC,DO;)4++\cfLVJT[<<Vd]K6YPcGF.@D3W=&cCIS))XVEU&WdCdGGg.+JLX2
<BY-)A_T<0AgL]>c,TBV:IL<D:Ufd:D-5[EYC)2<G?N/;)<O(<],H.0LJ_S@bMW.
Q.+/AK8SWRI=I,^CPQd/;/\ELJ[;KK0bBQD=-:EDF>L3)[c6PWVNVW\S=W=9<#:-
O.6eV=B/0A;4/[[ETG^S5W\D7&&T-[V4[=[JF]=F]^S3JT+TX9#98J9^J(aH,=O6
Sd4b1eK32)@Y+2cXO_I/a<P0#O];SD539ca=ZI&==gPYP4,IF/@]VMNK?&[P1#7F
TaF7V:LP@e?(RBOS7K>4(OePA2O(W[=WRHKa6TeXVT(6]I5Kg@V,U[/1.d;/[UOG
DT0&(M9Lc(a>P2U7&P>2S)NKU=L,eX677-6N-@IgUV;Y>Y_N(GgH.XO,K-[,QPJ8
+EO;GGX:F_fS7^R9F(257PRL/8a-^,E86_Qc+;cRSd@QRNZgM\O.^g92P++;D2&<
aEB5^/d--accC>+ZJ?.&W^g-<)@OGM>Z4,eXae[T481>CcM8S0J90B^NC)B<H2&)
<_eF4Oc\V82_DG#UG3X?/Qa/\.LC+@Y&fgL#LW9a6L_:<L9BFba?Q3)c)1EIdFW\
M#B0=68D@9fZ8/G-+05c//H<Wa+LMRH1V2I<@?Z2c4[ZR;=?X4ef8QFXR-9AQ(dQ
2-G;WAKHP(:d9[OMM78X4@_;TXEE^)@D&1Z@&Rb:J98EJC?I502V]AB<TC.G2?Ja
5Ue21\?f7&&.(7F9C,e3f7BMVK\ea),K((B:;JaF6-U^]K+f[#E9_M=0VQc@LN:8
[IN:6=]2LL-;[FTDG3fR^<>9OO7+ba-8NY4V@C\_1WT5AK65<N6R_LQW[0M8:,-A
)OCC\#-_RFE1fALG&Yc>Q:3FR]Ff4VK_4_-YeTQ\B-ZI\M#1,#KRdW\[RN=O4[(F
;@#U9fGT;RAdXP:Z,&6[>CIMPEg6;M1/S@[7I<ecOVA1^DFLJCJ;1BLY0]QFf1.<
6WVE,Z9=e/+Y?06<P0AHD4;2[,(L-YLSMgNPSCG5A3f^IZ()QCF-(90YU-0GBg?3
51Q)7#:OM\28-6,KbVR8G(S/T/;G#cg_CO5R]g)VPgJ#BSUCOR<<X.XdIJe3E]0?
37ce@B4KE:]L2H>(@-GfV&\-dS3F9_#)a=0@#D<f9gZG##R>,06;3RPf,>NTQ,9O
e+HTOc]177\GgDLP-e<W(4DdI8RRAP+P#M)ZgE8<+,?GJKZGK5>CS>-bEA88H.aT
eSD:-=HI@(.^8M\8A6gEeQS>^0FCE;S(79<e90IE#>[aO_7OU:;29<^=:>_0+-Y/
8eEa941fH+eU):+46T8]UW4.7D#MaT3N<JB81^A-_E#_<6I5--C2C6T+K#E<=LeZ
b(;8.VEdR,-O\\I4F;CH_N<2LPa:O)LJ9><A4+MW>#FE(+@H0O=.6=&.ZIU8+fQ,
BOKVF6_9aFP]2>.K(bE,5J.OY?\Xg2e2GJ,)3X)FR,;@-2a;F&VLP9;EDTe.gXQT
Pb:F2E9=+I8U=)8fGd<100X:J(M3PJDZX\a[8]]B]PW,4<48+&<+YH8?_+egODVf
6MU(3:aQK]-/+]e>4C_#+]/IZVVUGJd\S<CHWT@&G,#XPOI;<LZ9GgbXU)I\T7N5
8-bL/-(.HWN#IOPYb+R9>^I7Pe^TI(a]QETL?)UGgDBYF+OT97\5EY>E,H;WYWb=
D^f9H?ZCYFO\SY7b)+cgX7TWR^_ZO1a+@dd20GD\X9GJ7A#Nf0>>,SJIAL\O;b8\
J7g6AYV)b,#?D[0fCNS[1c3bDME5dg.K3[\dVGc@0/2H+cC^&M&Z_<cDe8@1UbAQ
Z07@g6bI8^cf#>6#]TB/&XcR0Z?3J<7f(Y_fC&GSZ\X49HbZe3B=E372PNLP&#12
70@Wcad[BNJ07G2B&bT,?P_E]6AWE.WM8Z^5(N:\\:&PT^f>7Q^M@S.cK&=\bV\=
(62W7d7g<U@-R&F_e7RPSEdd+SN&gV=T7^B2+9R)D,,1#8YeM#O7dGR@#eL)/(/c
#(6=3.DXW)\@9)P\WM^a[NN+55>eS0L\bP=:]>_.=a/.Vf:.Yc5:W:,KP4#>EGSJ
H.HbD[>C9F,e:Pb4Pd8\f0eWa19>>R;>HZUa8Z,a0EZ?I[O^-4?6>e;5:<XM]5)0
UUfXbI]X47dgE]Y_4@&d]Tdd-L^1#Q@UEG/g9=#)c:Y[E&KFJYGV(-PL3G<9;W4g
LZaU\30=[.):?Z/[\Y5CbYR>AKA93T]HI63GK0)3[:](e:CI)R3<K3cLIZY-@EQ:
Z,:RKS@#S<)T(cPTXfY:LUPN_J9Ac1Xf1geE1\Z7c<\f,RYF3Y0+]+WZfg//2N5d
D_?@f1H&7MX5;B\+c\e?X5J0\-LGLfZ64WFE&Z&ZJL3+=3d1KS7BTc,1Fd:B8ACg
\WH63Pe>c-c1OX8(XKH??(CK3F0R_9Ta2)PbDG,^Y??4P(LP[)0NPAa&)LEU/39/
DXHdC466NLc4BI945FVE7JPJ[F)G>YXY)@9E@)#7@FS]F)F_W14J&BY8U=O[SRGM
.@?Q9EO4Aa=TH].:YaaD=[&c85;gcM,\Z4]FMCfRaN9]JS\T[<,FXHFWbNC&SL@]
);78;U0-#-Nf_.L+Sg;&U/[XfR4g9DEEb#-2:I^-9Q6T0\CF#J+cEc[WY9cT#4Jg
+5dg,gF0YdH8<E_3O51(U@]4A7DG#IM<S)BdMg3I-MLedBAM8K.[PC=#^,Y5#N/L
/+9T1f]ZQZ&5KEI=YY;aC0P(=6@X[AS1e\SN+SKS(UV6=Ffb>I-f5L0G@IVP3UGH
VX0LA8:6(gT5TNRHA/)7MSXX-X:cE(5^a(B@N+,U85Y1Fa=;GbZ.J^N]JI:^_(6Z
@EGZ8/=dQH=;4)+fdWD=J&BSK/ZNM/,=KgN?AWA_#E8MCM?50,XCS+0X=dH)I4S>
(;bAJ3dBSY9H#?I)9;5Z/dTAg8@US&cW6EG[8=IJF._OP7J(\AKbASNWBZU^_/?-
[YUR2]ARZ,XZ3\_cPY<KHFN5D/[1-)TTAQ\K]>FefXE9cEc>dNY?WXY\UQHB&&.T
.);)S&V.Db76JRT&/:?@Ld8O_U;>;3>P(3O-Y(BT9d>8,8^gAAD2(#N9H.UWBB=2
,V#;J_I[WY<)=Lc^VAb/N99Pa,YA]bc6E?>HLW,e?L,ZgA/ZE#(DW\BfE-42;U[]
OPBa9g9D/&gU0X@6>G0HDGT,\a=#ZSfX59cWIEM5Af02F@?]ZO<Db1H9U:C\^\3V
a].b/]YX0#TD;IYG7W&;?#[[7X3::A/4EMHY^YPXPX[(S7a?BQ^7cKg8gH3=W)a7
:141T(L>aBVKE.2:?g:-,IS=,\DB]H/@;3FUCDI5@G3R=DEe=NL5&Z[JXS9AS_V6
-4262KWd(d<,6PbT5^,XME9.UHCbM?T)+LR5L<]4CPL4c27XL5RSVccX@4D-Va/6
9H>?Je_[32Ga4_)2K+ZG>d[g.&_DYd@E;#+JRVZ]9WHf.8+]1LLc:ZZH2.O_B61;
b9<:03dSAc[&KLH99b#^Gf-Fe.4=P0J2]\S;7f_2_@URYX9]K)G^+Ed:CKI/L0=B
7EXATZOA2C(^Y\82=3<KeKZ_W.52T.QG=dDV(J/GA4V@L#\<Y=W+0W+\5g+fK3:8
<__O1SEJ[:^:^M;gSM;J7aHYDM?C[\,<OHYL<S2L2/&BeI91D7(9=:ZWc>ccTKJ;
,)B/DQ4M[6^7QI@6=fdP^:01,aNP2)52@)&44.+8NNT/M^X27V+GZF37WK<KU9]&
2TK2P>Q;@39^KT@,#?-FUefS_RB</,?:_(#]348IL1[#,Vca?]/\3ga1C:@3@>_g
^DHUGISZR#9QBTD)OU.+G>7#519>03J/&B4Q74?OKa3X>dKc(2)@d<NSZ:ZRg\4K
gORcdCY_,/4FAQ<@_I7/26C<L\bQR9JW9/(##XJSBLT&SbXe?_BM:EP3DW@#W-VG
Y8JM0:2>6BAZA+)a&];<2R@JA9&IE+;E&-9+2&X&T1c9,0^CF2WQZK_9O>,X/b/e
(bc][;#T?+=7LD54fDZGP9DP6,T:@B.HGD2egf<TZR&gXC>?E)NL=NCUS;DMH4b9
dEf,<[O8CF]Z5C&7.M]&9,FHI2@IKf_a^?J\;C=-XHPSVWD/;G]_WJdZ;TB8R(:1
BC[A][FSH/G<PE.+Kb/NcZ[EK>51<Y&6)cVZg7>NM1H39[DYK&8AcF#[Zf?>5B.V
/),.]2_]P17C3P(TP8XSD#.T:0fDP(O<4dg_D9]ML@HFC:&N[&)<LGH(S3]YT;[L
4BHW2aM.Z+C<UNVE9]O(9aN_;VT=,Y\,R<d=(ef;f8+B:X,CePcHNc5^fVeSBUPU
N>1DVTZA-^B_Q^PO6,3,Y01IG,Z#8-<(5/-),f&L>)@8@_HD;YPYeO?UTM</_bS\
:HFCROeIFg4V6:aH:/ZBd^J5SKV)DQIYb[.3G>W^S9FEW=7RI-1,Z+@O+7LZ6dQW
PQ\?W4G[62\>#gBeR.AMe7PUb[1RTR]^b9Y]Wd-HaJ&]IfNIU:LUWdJ6eBUd>,.K
9\#]&NaI+1EEAE&6cX(=FG&)L8.g\IO9;_(95fFQ[U7]+L^g&EDU?JF6.LdST@[U
YD6;5>f<#@g?a-X;Z1O<8F?=eJ6EFYSW/#Y])_0WPSU)ZDVMdgZ976GPb;F-gC3U
6E=G@+Gc/#D;)D@+,I)T:)P0K=?<)9Ie;BS?;(5U>.#=T^;[\21Q<1_-S=4eH912
92QJ@L90C&,S=;1aH29=.>A-1(>#?\eQ\[H\6\d[\R38_[S?S[M-eO+P-+63:FE2
-U32)?S<Z]YgNR,7?+F[#Q+@/0^^FcLE+_)&VRBFffO:KL8b(=+Pf-@e_?ZJd8DB
g\1g4Ne&8Ba]SL\^^]6T-^-U6(7<:C.YW20/6MJT@V\/KP17eE^LWUfL?,8?D+-X
g[3a/+/[U[g@3<bAE7Pb)DW92]GScL2e@a3>62=eU0J.Q=;e:H1DRdF]U&VIUg=A
[Ad2f/6;T7>#CL37+9]gEG6[;Y#aLeI6PO,f<[#I4(9SgIWZK(dY<?b40\^)agdT
eX;BRE?[W0[[0@ONX;UODXP[Z=.QUOZ)TQWfE1.:#>a\2\=OYWZ86&AX.[MaZ#W,
2?M=;>QNVIPBK@YL-AL-S0P],X^;XNSb52TeS6U[GS-M-bbW+K;eX9HB.0R2MB)1
dZ61FHR4aO5E5Ia,7?KSFF:/Ta-5AS(EX9EbZd:c93B@)IRT:?c49aBBF\K^V?AM
L(W8RJGDBS<TcF\L&H.CFDe-?[C)FF3,9+Gb0f8&X+?c5T>OLS1<ePcc+f-@\HA5
H<<H<cg<F9.Kc.CVU0HSH6E2+2=^,?6>fE.V9G^5B2997)bb7\(\]RZVA(c[SYQd
Qd+d=QS64Bf6L]7<W9/C]6(0ES5_f?0]aM)SO?aYP@8GG2T5P#KGSK>19WO#N/KF
-H]2X^1.^71M<OT]AZ<M)(SfR/?eZX6]g8>e\F@E_F+.ZS71Dd#=\S[fAN&#T@;3
\U=7V^QF).#_U6RWX>#]=]<8A<8NP5bf2<)S)E1RCQ?45.KUNP7DI=1?;(;O5f.@
S[;2EaKC<6/HC@DZ4N^=U3e^FQC#OKcWFPMO^:[CE@T9HLA]cR:3RGB+<=Fb,De8
B&USC9:f=,4GM9S@)2dffa2,eGHQS.[6IP<,:\F:9:#6O\67]/>3)=H.;C)eW6&9
^>e:^YU>Vd;&XYPWZ(P?PTD>H@1F?<f\IM>WT6\>[^9O2^RUZZCW2W#>/?QQC=N-
;Efd#2X_d>92&7[SSR?EZQA;2^Y]K3WbBL)ac+X]-#c0YASb8&Md#4P,T)SD[H-_
R/.68,c77f25YC>F@>F6b3bM,O+Z9ODc,N#-87^6DNe=J1Sa2^7^_^B-VEQ0<<=C
=(&e6^.T+[C4]N]/?cWPJR-f7\XXT\)H28OAgLH1M2#_c6T#3GL7;5][D?S@]ETd
B#[N<e/8Y.ab\L0L7:X?YH8O(63Q.=M[^L3K9O6,[1g/[4MON,XE00]RAf/J[L/1
c:;3\(.<QXX4G[B8(VeTg+16;X4LO:,Y8U)G<B57#NQN4IOH_,MQU&/RGC8,c^VL
G3)Uf?1_Cg5]1+ZAI(_-/d#]2-=e]Db^+^K@(SP^/#HBTQ43f7ID/66(&DdH1714
3c.dS2X73<cK+Z0^Og]HLN,X[QJNTB,&<d(RQ+C-#O6Q04ccNAd)QZ=eT:63D:g;
(QGF)]\641<]E0H-^M?^T0==U/ZY2bdI0K1(L=,<K/0)\b2MGZVgJ6YK0cFLV9Z_
KG,M5R#294Kg0#b^(MdR)],W.g3/8CO<0AP\d<BU1#+TSX7TLJM?BV(92:aBb9bP
A&L4E?F?E92>We.3eIY]HX73\N[#dBFVBY2M(>_5Aa/)[.T<W;Ca1^60fK?Ef^>-
C9MC5\V<WT/B@OCK872MWTD[9UX;:Y&T_B>GL=Bb[Kd-71[MIA5+=GI8L=FdWfRG
e)L)^W&XA:8ETJMR#&GR4b#\I+#K6=VQ8&ETd=S+#TFKe9.fGL?8NBUT^ae7N;a3
]D6N__<a6\,;++aR=<&Q0#^&J7LJ(APY6;TV[7>SY\HXD_ZQV-_&<c[0JK\7CW9W
O>2aX:/S4XPH:HfPTdKI9a((_NF/7S8&bgFRe9Q.7b)Bga_RW#_0IRF0SU>PDL#O
5>/Z-Yb9)2C7SK67&3_:I(Eead[3Cf3.B#,]5e?Ad+bZ1#>AA&[#=ZeeS-S9]LG4
R_\X.RQU15U4RU^U,_?8._f7FR+C/cFD8gAgb9;&Nf[D<VPRF9JcH)LZa#AL@XdW
Ua?:ccZL?5CDccKS/TWHBVENT/[<+MK\M[Sf?eP(8:D#a=BB8A.=A0M<K-:PEV/V
O;8c[5XRA7C6\RW70ADN1EQ/)JDR=Y[B@>Q()4HBDP<LD;^>eMF)55^(?b.[JC>0
RCQ[<MKJLQS?^N8;Hg\>LS7A48=75478NS1#GG#8R[+B_7,9D?@?6M.OU#F8P&-H
)[C8Ia::;G9dXNPgbC.::]XJ=XW5]Bc3ICT\DH,N2Y@L?2F\#aF#^4UJ^a2^AD3D
6(57#D?6X]d?:Q6cT-3WQOP[6@_7]A@4=03?7ZTL#+\K:c.Q])K(N^2W[dNLZd:H
U=+8B=:5<gdePS5\2Z[GELE/4[#P>e\^\P1SXI1ES(&7DS]XFL\b.M^O2EfG)P#Y
d0@;XKH)fR7gZ\GD>^GYA>_)>BHOR_&5KYO7(bE[S0Qd2c.1CV-0B==,(I/Y:Vfe
8N?g#GJ9SC8#V=)-K^8\/MS4=1MR:]H8Y(^)J0-)Y;RgQUKOT?#ef^EII/U,,FI?
e.2g0W<1:M_TfZ7PQF_d6CNObMdT8:3<)8_BfDa#.R)H=2>\Ae2:94DI.PG]:M=4
6BF72aW+:0_L958ZG+^gXUTN9a?6WX)2LUR9A\KeZO\fbb^NX&WC#]MD=CZb_bJA
4_Y@ATaTQH8<e@a+=RZ3-MN<>6I_#;feLX0HF,#NgUNBGGFZ[e\LX#W8W=5FE02C
OC)a(U?Y2_Vg/\V<f:,2Nf^N6Nc1^:JTU:Y>,5\\@X5eZ:RF[g?Y\?NGWDU:;5I)
/S7<BG>Z,9e4</c&>\&Fa_<=<.IN7JRU)fCb5bBK[_)(>8He;J0_8@gaB.a^)9@+
RU4B);a=S:d?4[1_B9f7GFC\4FM<;0G<?a#a2,KF5GE<+b2c_HLR<g.X,a/0b7(L
#Hb5SG\0(cJOJWC;8\d7>)#;[LQQ-:\:2M.=E#[@)cNUYL2581ga?N>fZ0Q@;2&I
;Y)M^7)=1VRQ+UL=/ddEJXOa=18[O7fIU<c9-BA8L<@WUUT2FZJ8B9KJ1GKe@7.5
WB]<GNQDB5-TKUCXDQ]E6W-+C1d)2[GFJ,_X@E@BG?Aa^>.3M1cK:G(DCUFN)TP0
IdP7L8,QTZc&Ee8.0#O1][1,]75-R&6=5=H3B[bO#CQVA\EUJT</=DTR-AU@V@\f
>d?9a+eg.\7FPCb]I^0G>XJ(=7DE^<7Q[#UB5SNf+a=5Zd:X,W0dX2Lae@.c04Ng
+C#L42,&LS>?eC2NLQSc_d6H@b2Mgg?AaX587AI>:[\NV4Od-R&]DW#)@1aX#1)[
ADd]@2=X:bVBBNPgJFU3^.)Gd\0CYE0)70QHH50N^?^S[BLUH\2/HG9N35Z^X=D<
9eTF\(T[M6MK7:(;dVf=S52,/2AGCQCAG3K--^(\f5P5+a5L9\SL(e8X\2N5(4[7
VWR@KG2MVA[LO2ULIfL&b94D#=)/bGX<ZbZ0__6)V.&>\<>AXdW2Pe5=J,Da4&:F
HEI-9\8;[V/H;-G32U13#.(7MM39ZeD(ZQ0g@C6H\1^EeVKDQO[[_H&&^D0DgIP@
Ddd=RF4J-8(QQ;eZYF-bA<]/B5afeX/F5Nc7c_18g[[HdZ8VMQaETCF&5c3BNHT?
AEbFPU_FRBGe1V.;;V&)ZQQ>ed:^P;_C8[BBG+dE>c4E60I3VLY_gA(#<&@1+\\)
?cJ+KJR#,6Xb4e)LW:(DgL_A_-@/DF2MfO0K5_@,ZAE=H\7]Tg<.fXF;b<3;U8eN
YTUN97I7/IRX)P(3X>f,)U/TWOd=S8-R4gZA_4V?6)\Z3?W=D)^USQ]K1Uf+H0aW
O7U+2M<b8W=VU[/52CDRK@SHfa#Me#a#)3cRD.N>;6,Vc1,68Wdb\Kf4Rg[MaUR8
0]/0=F/L7&.RSD<GH@M8O6HMZSd/b2R\L6(UG#-B4^AG40cI[:T3-+LV3K+\3(ZG
.Q=Wc-<RQ,_=,Ed&-O.69YFDI+PY3TP8;M9:=TL6@I\BHPa=&6_HTe3&]BO&J,4_
ZL3/eT8J9c3Y4SKATV5>A=dTD<]:_:G@Af6VXBQR+H[]@#?Uf^DP]>,g)O8&7Eb#
SK^J9>D>N6XJ5)MGW[IF][0)P2TLQ6O7HP5^=X.DOBM<:].EG-G>Y:UI_2?8Z.8,
VTYIR>d82_JbG,-G0:HcKIU[Rge/HJX.^Q-bKZ:2AP.//#J,f[(BD4:Y^^O(a9IT
U\_Y#E#IHa087?#F:ag#a?DKQ5@feaAEB2/&XY\Y//V=AYL]L6aXQVabXHTRCBOK
O28W7I6</54e&PX57(6,eP@=I]@T>T9J/:<.P;_\YM[O8_cROH]9S5U#IY^M-]9T
>b]_NP/C^g&X&.:bSe=9DZb5;M\?bfSZ0C<YM^1aaN)4:[7-dEF:WS-J8O/2_9T;
U/4(00;bZaTZMQ)M:)MQ5/bTAYSd)0)/?8DK.10/80.R@#1EB/H3_ZH-AX/Ug&:0
MV^2Vc6,LW;[beITRX+L&VLD#YDT&X\YgS>(KLG;9Q8aT@80)YA1?V^RdA=:JSY,
6&WF@:]X4ZXF)T,(>=X;L\1X\8(^&,J&)]H\Oc)-ae;][d)T<VTVP>E(#R)^HVN,
HRZ^\/5@>^:HG7QN8.:6IGBR_G\TEN84]URM:&&,Z.3?KJ<@+4]VEV:JTdHE?gd5
&P-20ZL5/dUDJ&O7A4I,W72U/aVWXVHVZ@G#U741T7\-A:=7]@Y<fLA1We?f:#]-
:S)__)#X#/=#9?R3YFYaQ>X;4UFZ(&c7HCUMLBY3T)R_^TaU7]Y25C+P6T8E1#\M
d:SO_3AWW&F>K)X99;A:+_bKe0Z+KOMWB4c_NH90:LLU.-8PgL_WT.@;0:ATE?)W
+\)]HPfAC=f:,9SUMU638g/(B]Z.]2,:D2NAB(,[1N(XR(/a4P^a;HV/0/bXa?H@
00KfU\9?F=g]MZ-#.^G9..VRB\Y2O/>P&T:=(=LYc29)RZSKF(J8WI_XbA9a3deT
F=1R8,?.-9<K.ZbYD)^;VXfef\C8(VK8B66d)\]03fdAR3TN_T8.MR]&EYA_]LNI
KYd&A(D8K4NgY,)4XHKMBXd.A_&P6J>U-_L,EVgf/1HAK,[:>)H1M5AT_Gf7V55B
dQODU88a(U=KYO.+Tg[],LC<I;-V<3\ID6OEc(&RY^[]#6dN+Lb=2e.#-)7]S/@4
U8&2gRa&FZ/C18M=??\HBaUXaF7@[B2]Z.7JASc>N0JM,X8G,569Q,LYVE[P)W]&
A&2B,VJ-08S-aI4CIGb[,9f1^/cXU>eQ7E@EKg9=2WgKWeYcO(@N^MgMaKBb0=02
(f^ATD9V7NKHV4\>NR+f+cF-OFP]NdJ1W&<^[A::4+;FeJc?(2J9/-7QXTAK:3b&
P/Gg5]YV?J@XYWB2S1PfYYV,_Q\67UQ[;I4#+?g9XFW<HI?M52b_S&4STH?O4e0>
c_4\ZBfJ;57IE+/TXWCY]eR3f?1U7ba,_37gJ<&f]:21D,BN@;:?@-1S_?<I1J&#
b+@[VT.8d8D=LOMVe?DEXNF/MHa0VdT9+0aK9R-AUfOBgB<Q4ceW_-R2O&5/:3ZI
Sf:YGaHdcgVD691dCZ]T_Z>aD31]f03J59B9^:V(+Q55e-ZSV]D66^E0,/.C#RZ0
#]3:^QK#?HKO2?@(#;7Af/JETMDXH[>#_b5EO,GWS_<b>egLTe4^]bZYHGXXH,L8
g(<OLeEaH1Zf(6R6&:(UNH66?b+VCGLa;f&51M?=,(P_E2MEU/-P,[B@)XfQUJPd
6+OI+MBGDE7DMOJS-7_5Pc5g(?e&fUVVcga9eH_/.2/J?3_:AC/,#EOWBJaW]bAL
B@g8[,L-M;HX<4,IR(Qc1:SD/b[=NVTTf#dCdP\:ZI<E+N&g,=?=>VV>KN>XGEP5
4WB7b&@d@CQC^#?d(N/>PXeVJFdV\SW_J0BB+IgW(,691c)>]@82XM/KG_BO7cdX
53]]ag0?=^UA\fQ;VRD9O9URBLQ(5b#HOY?1Y-=WQJ&?YD/Z;TZ7BJa((FAJFPQ&
;Y5Tgff)b)gS(QUH5?<If>^,Cd8<M).4,]Q(U^/N@39.\M[J):84>,gc?I=K;(R>
MVF_\d6:JJ;>AACK4X^P/,_7Ld@QG6.)V=8Z:E+#GBN_YQb&[f>D6J]CYNW.XX2:
:T2S/NaD_fHGEL(4F4BD((&8&/-gYMF1Qg.#46#\[LG1^JQ^@ALJH)ZDVH_^9=.C
P6_0A-J2]BKVH.bC48fR+A7F6RJTLX=;X]7Z\>QU^.@dP>YZaW2;6dU7]6g8XHa6
:8]c[3VgEP?1U]BFaG&6VLE6\DEc2#)F,,d\VSF/-D4Q8Z1.Y?&dK-^(^Af2L:1\
N[V#?CU-1K<fEVI50<AF(XV[-Gc:34W9=Q(7<H/MdXFWL&f(C8f7B5;I7fNf;(7X
QAebA_f_,E#3eN&D1/K[RG=\XRNUc7DcOA;2^ENT6NHAV2GbXK[Ba)R6aaNQK1-@
d51WAC]<CK=CQ1@TK1[WJf4)V+)G2;_U6I)Y&+)0:1=e9@Q#_Te^1)XQ+X/XA+&<
S2[TgEDF[I];(HbgI68b?g-cT]N/)A:^a?5[Eg.L.XF0(7ON^AX2G]>IZA[PH\@9
NbX&c,0I3BW2OOSBQX&FgSD=@45-KJC<,>]+CAbVEN@(R\NcV4EJU5R[I(0b/Gc?
E5/KS>OeVB.g6U4Ng5(F(;E-<YAKA^SOcKAHYQ(8ME2KTY-R&_JeFY7&<[:&ISIK
I,5HK7E^>X3b)09@XX[(;A4,V,<6B2I36DE+WY.BbGD_Z=_KJC&):Kd.U?G1#V3>
=T0(_a#K<6[D_9IRCR&cH]1I7\9]TJe1^5_PW/XGd/BB@35/OELP+8g:+^2FY^=U
NS?_P&,.>](=?_#9=)]^UGgIZgP@&KD#/,N^@OSLIBW->J@RR;MLgGX7(0b/UR&.
dA6-e/Kb33&F?@<R2C1?(DO3IN2K?E-e8^6R^2HBYWB6/SGN8H(YB<QQ/(5=c#IX
@eMI+LIBgV/aKEA(1AAF=f=EF]11CJ2G[4:(3cVWJ8W&bMT+cQPLTYY-^(S,03Q2
OLS:?/\=?=bHD:PG.6757R0RaOA3PXbCM<C0fZ[#.b@c57;/S+N+LQJObEcf?/d:
QICDJAL&RI<7(aLR@]9-LAP^U\TEc_K7X#?DSfF[K5R4T4CS67-LWLC?1B->3(7M
V5;CTWDK4SGaI?c/SI6OTQEMG794FV\BB:f32K/Q[S&VV4C#&_05+Z>@_+DV6E(+
R[)HB?H+T(&/AR6BBg^Q:8Te]:FHYNVdSK-/NL0@1AfZ?>L-Z7B;d&e98\?>02T\
3Y?YG]?8]=+cIOUJ7XK,c[KCKBADEC5-eZOMBL5^RRQa9DGH],K8R\c>]NIcYJ]X
TFR&@H+?Vb4C<=8-1cP1VVPV&a6e1U\&4HY5F8_dZ=f-Ia:SAQ?3A,)EMGO[\#?Z
>MZY^8M=>A,T>YA,]V/99N4:TdE>KTV)MH?(c@FK@+,7a6e1^T0D(P1ZeEcXL>E@
C+4g3fA[];N)c=/aP7fg\^,acQX[G54@\+(M8c@b(,9HVZVNW2<N[F_)UU-)X7@Z
<d+#e8<5GgZgHZ,K4E4/4;[+QG]6A@_&ORZ,2P<[/BA?Acgf(bR6;dXGL\d2F\P^
ba(5+:O75FJcca6;K2#5QTga&gg6U4Y#4-+66;-S2W8R?R&I.#KaD;YXObO&>N#3
9ZZ_ba)MKg;T\V(0g9-b>/NP@@>.-P<7fd&H;8BfJU5P4F\4HZ-d>4QQEO6L,#gD
V7578)@+bdBg_b(OUZ[dLAf=;DI45a:-ZfIdG21X)F4&cIZgSK2-9:[)Wa6@]Hd=
LRGB&e>(Z5K#;:+.8?fI-^VaGX2GBFTZO@d,PH^K#H(8\@&B#[=bXa9>F3gAM+=E
CeR\D]c=Dd&ReI3F6Q7Oce3L)O827(X;/7W\Db>WU/J7I^]<a8,LC9^&_]+\D9\7
OD+6WL>&HHdDHDYEVX3,(577[5\J4LDYMHaB4X/@8fWT&I93=Cf=4^<:9+Sg)Q6d
:@8]fVZaR#EQ]S<RIHTD4PC/.BB?[[54Z/TK?d_(&DP7R.eV/3,:+Lf+/J^HVgW&
?8C<8MCY#[ZX)R6:>>/\(9(a>9)L0?RA[#P9R:H[51c7EJgH2(]2@>>2F[S_4e7[
Eg+b:6ZRPPcNQ7>@7PWV(AA9fZ:H_)PW?IQ6Sa5VR:GID9TG,\f7JW&f3W6)76.T
I3cNdZ@EVBe0A&R8FX#AJ6YI3Gb-J3-Ie2AePB#eB4LP[)XO30f6&A)=aM,&Jd?7
=C)LbG6UVM7\(O+V5SI_d,&6b2e3eZSeRXF5e?WL;+3Y<1.-^;J)-+9KMMGS4;c;
F^:e\)?)EZ#@4/.[@4ZT9#9\X0NIC3CE/4JbGSD?SG(J\?ABY8,YM^\:?036C;Jd
0V-;#PQ9c1c=EVG^J_Ob[W^.P1Cd;^R6S#OfDXgEA^\5S[M)Ne\47J9U8L6e^URe
cU;_80\,TZY\&(8[PZ+bPVA7T^V18(E:Z66ga,B;Mc^1<<=(1dF47=+<&Z&]?&95
2,Y_M&[M_8WWHW=LAK8GX7WSWZ>A?@,_2#,1O,G]]O:?ZEdRPa_Y5CWf2:)gO7(C
8C_F5@b[@YWgE2:)W-BMG8X0YB/-@>bM?2NY&I6LR2L^\2?]?Lb)Ba@N2VN4LGAY
C0XbY8L_O]U2gPb_Y1>;#f9X^[5HEB]:<(:J=L@)4./&V\M6F_E<EPXL?SF7aWKK
C:Hf1+\I>WS)a<&Uc0RI8)cG#JgQ>:ZP_+M59P@E5dXd]dY.X=RgJKB9OAb5WPFc
fT<.&TgYdM@>,Ea=gK;E)OG)R.#QM5H:5E\(T4+H(LFW1O-_=>MVGY1?&X<Z@gH[
fI62;.Q)fANX.H]bCA,b05SJ2C-I+)S6\aE>S[6-Cg7(NcLW+G,dX&F2:+ZUN7(U
K#Y-C,ISA@IRKS<Q78]fDW[)9B5JTZ=7D;XJ]EO/>b8A1[K+ZPTdJ1\X8V^24;:K
JP9Sd?2g1GA8&F35?L0-a2A@cMLO8DcEE(NGdO,XJf&g:K6?Ie_=9K4?K[L3cWc2
G[U8Y@)[ab]Z,GZ>&NKXT_NA8f\T@4gA)e[S3[&1>g=A60SD&g3-^bKQOMM,IaT#
(UdYWAUO9_<]6@00:16Ug&-]R=g1@,M7BHb]&C-B#AON;N24Tf_C;EMWD,5MY91R
A/W3L+-6OASWL31.&FXLE^#^KbI0Q,Eb[,AB(4=+?B@M>;0@.\7<;78\>L0Kf&UC
THXaeRBaUVVU\9OB<SD1QQ+c\F(d6GEbZ^Z2[R2VMPO,ZI^c:@.^Sc.BNXCf^b3)
KEKAGDZ,.bJg,DGDKP>MR;P9,4^+_:-/TK3&6R,V.24O?R]@TW;>)T)HT/b4a3Z>
.;@PPg<S0#b^X4:+XCPN:28M=L81E7E2W,GEPT._H82>1fUSeGY7TPZNIUD1&005
bOFX;g3b8MbfFNDR(3N(R/@3J4#e(dKS8XD8GED+HJg)B[5E\1J^-KNaL\3)-]7=
MY7edKGg&S:CUbLVaF-A50>RAOB&9>23?d\A@L-2W=[EV.,\H-;9:)ZVBY1gA?M1
DS)^eT,e4JVR.?3b@fV>(8A18[1fYDg/TRb-(2#VHIC&5@Z[AE0HO.=5TCaW4]C=
^YTDd=\=a]>J+NIJJHC;Z.XNQ8CN9cQ8fF_;D@?E9CL(S#I^H=I_-fc7IU<Pe^g.
M7,(U/7fHIZ_+bCB.b,[_5Y:PPA5]fN839]@,e.eeP4?G.5Aag)P^FMJRP0a@0g.
QXg),D:(9AN.W7:<8;UNbJPAR(^CS1ISUN0<;E;Kg0#X4XH0^fMJ=^^HG4BN:211
6:9M4>MZ+ZG[JLYKS]=0aHBg1.4@[769S;NW[,76>edP)QKXD_8(6FRaZA.D^RT8
=(M):G0_CHK\@XGHH^JYCO6E^,=>L]^g;=Q,c\&1P.fU-gW7H[:,<T0F1YNVS?#7
AdL_Y&>=(CK^:7>W\4.UQ>,3AZ?(5Z13-UfOc^7[;e^_KI>.DHeXT>EZEN_WCAdd
/KOL/0=A0d+::()05>OBdAT@7(<_A/FR)[JJ++_5-&Rc6/1##WNK)-K<.@\7D[]a
(BKcLF-G6J2FbM<ZU?&dSWb-eZF#cB<C@XG558\edIW/gX-f&B(CWF(_@[B+&(:L
V[I2F6.2fa&:4D?d?PK>CDeP<,1X;]L=5Q]Z?Af1KPPO(C4AW0L&(_06f,</5,9-
8TI.aCgEg=I4U]-7eI\WK]E8J^^\M7eM\IC,Y:61.HaWM2#[B.\egP+>QIY839B.
TWLcc4>U0J:94cZT[B?NTX<QWHf)52MC4MALF?GHZ2+]V]DNe3&QKb16+0<4/=EB
f@dVOd(>\6P8^274b23g\5Q\XFV?adXMPaW;JN6cf61HdK4UP644F&bH_KINB0GF
6B@ZY;@^];ES<JE9WN545f_IVd)J@4c#1)47a_0FCK#8K8N4SQ>_Z5W(+53cBP.@
)-]+_f(Ec8Y=H#;C,7>)8>LQ/\NI;E]PGeTURQ4:IeXMUWXO-+\0TbS2bPLF5:H8
Ie.:=SWQYO;>FaBM6YXAeWaT3Z<a^778,:90>DTP5YOd\,4=IHDI?J9OE2/XFX)4
gP(GLC@N1,1^2.dP(g[FNTS6&a(U/+MQ>HFb2DD2(aYI?8g4=LJe^H6L#bRCK7[Y
M=/A3K+@,Y&AR&OR:[P5fW\17[DIcR#73&8&<>8VM<UM50<-IdG;WSQBB+a.P0JD
>F9@FD)YFYGIYe-4(_[6fL#,,O&GDRG=ZTWK=Y]:J&((KMB<VBe&1C&<#Y,U+QZ2
8G0H)SNW2E6C:Y9,bBP8J3LAc2ab:;K>8D+-4]5bDH2Y1WO3:(7L]SYQ9LY/=TRB
Ug)2.b\F@1:4gT=@__)&Z5(A@V;,b;6&@d>RDVVQ_+X8a><Q)TR7dQ+)0LagJ#4V
P,Q=5DT7WU::TM[dgH)0Y/-ID\20^).^N2c;-fZ6DO>UP1[\37GOBDB]V?2gHKB+
E2RKPN>RSfP1\1E5.JFf3AVf#;D1Of4[GJ_ILb2)cf@;J5R^;LCdD6V^_#gC_U;2
A],7VMH.Y<=BYT8)L,cY<88c0]@S5?7G0\>SRGD2W1JIAf/:W4>9Yd=PYQIF^3JH
+)W?BfDBOF5#Og33@0#WX+9Y+HH8KV1.g8[6@<H.VX,];L]0?3KO_Y:H9K,P7d=^
;Ce@FTF8VMXb[H&Z_Kf_XK[>L1<\@9Y#d4MSZEB_@bg#18=+6>3<TS(c;\K-][gf
0P,dQ(T+_Y=YcID?<KbZ/g\6)L&2b?>9)U+PX?.V._SgHC89MY?_U4N0YP)LE^AG
-2f)[0eTP8IQE61:W>F<V8^23Ve/K53MYd5W]?XMNPR=;d^d]H/eQ_)GGT):^+/G
f[OdFE4:^687EKVJNPH#BXWDZA:X:W)N.<f3@+Z@1(5TeBO_13L\B4SaXXASAF-c
O1P=Y4FKL=GTPZ,]Sc\(QD(91R=1CE84DJdT\f;RgR)AOC]d5A(ISW3\G1D4COc:
2O+#L>g\>bRT^8],P5-e07GOPM,eDcIVI^A<M7aD^bLH82SUA2+F[I0[]\YU=[<8
PbI.W@bZBFPRH,,C8AUI0UaP5>/CcB1H.@0&_LLO-IKY/]F][\&bNNA0E<a@@XKD
c7:\5+If(:Sc9IINN]R_.><AJ[(<G8C.(Ka2,bKVDTMCFPM5?SQ2M,I]IO_58S?@
ZPQ7dc#,04J?;Z[M14=O:]L)>E)0B\dCG=P;6Vc#9_3g<F_N(B&0-D1GBZ383_LH
cId3:f.-:.,75R+XSg8:caUgB)@QGP;&@[O0g&<0VVV1:-XUAGfVCMWGc.Y76ZM,
d-=C,GZU6>3dAa;eNG2NW7F2g5&c4F/WRC7;8#(\GB^Q:d9b]X+7D(=/&2W\EL;M
0f_/J@cMGQCYU5g&<P[R+7_WB@<ZNUc5(K<FHMX.7&:)K.PF_@NX5TH:DLH8SRR#
O7X>Lg=]3bfX:0J>O./V[ZH3aVQ38J+V87PT@AJ5=WIV3UaF8GBg[W=#c6VIJUUD
ITKPJfLfbVP8:6Y8KeKdSAIBE5GS>4JcHYSf]EFTEY4Z9ff#&IMF2@8^>1b+=gde
,PFP9#U<WE.(0MP;HY.a[-_De:>UGbaS7:BSg)K\U<Nec/.RWPPR1f]58]a8-1+X
ESB4ICdH;/b(Q#1=c?KY-UFa[=XCU<NC=dUbXSD]OKL,2?_,Uf6B@H_gOT.5,SRI
W7>,cMJ21d]@E#JeS0C-<?Y;Uea=\gY;NNI7GHIZ/)95U\.<Wb>[<II+S<\7d@7g
dEgLfQ3I3S\9:cGK_>\1f6OJg]DaaYDd/LO@L0bQg4:R>5Q:FYL67X9AF<#f@8gN
KME_K2=>bH4-5Y(bW_MDU+XJ?b[4K3A(Z52_?N&Z:]2:BBK?5GB))/N=+dM9Ng;<
0XNB(G0\^e>FZ)1Y\I7\)(N6=-AE\]gU8(KC/+Z/eJfMNBL3TfUHUP#:)Xb(#g-O
Id:H.e<VAYZC]T&[+5d#Z?E,VLY(I,+)cH:P^B:(b&S&F_fB01.@U-^-9b.45(1V
[IJWJ@5eI[&N\<P+GH1):1ZOa=^\gVC:cETJ#/-KaK&,MgA+>+_OgANf,82)MRP_
H.c_N-2LUZ:-WDZ6fKbU/#3-.eQXP:(9T8^/;T<S?LYHO@MIXf?QND;OKUaNRR59
b1=(9C50&+M]bHA1MI7:H0M(X&WOBT//&]e9W75cT2aHMMV\a#Se(da,@eCbA<GT
1#8/P&4R_4Z@);;XAOEI4719V&=])..]@VMNa5@b+Ib8Cd65gg.#P1>Sg3<&3FL-
HN])W=POYWN;YC4Vcd/GV;e^VVBdRM&L4^<BeE]9\1,R;WP6R?+#SK4&-4-.M_Xe
P3HV+G5T>dOXf#QL=U4#<45,.OB):#9]aL\ZF)Ab4EJ7L+RNTS\C/V\AQP,6/aBc
O+6ZRMT7V-W\]BK_,c7a&(X]UBUfL(/++gQFa^>>SUBe][]0U=6e^dNEe)3JCWF@
>Ha^TQ+eB:f,X5VO&HB\AI1(7.7AS^LLES0-U#[)_PA4)E.PC^=E.[8TAB@8[6K]
:;L:R-DC4aS+c?Y^Rc2D&eCY-HQIaVf_=6:&N./=3c56fW#B:B^9V)<LA0P9_^PG
9M.+LNbN=3,:F4a-7G&F.^c_[XYRcgM-d;9,)0CJP&\3TJA.G9+XG,aRE9[3;GB+
O3CNd,@AX#;5c68M.;77I^PI;F-9\<EFZ:8PQ201JS2-WF;FZ:<?@N1/1MQ2XO?.
X?VXFEX1.)CDLZ62OV7DP383\9X@1111bR@Qb6B/gJAJ4C3c4=-N-_==gH/cT^O#
5KeaER]\O#45f1B64&./(5O.3(OOP2SRb@)5G/B,d>PXI\UALD+WZ@F_Ed28K_:G
BgH5]Z;COf;-24F9\cE_EMWb=?_26.X;@28_@FKNX^22LUMT&GJBI?BZ):]U4eM@
V=5.X):I:G):(&NZSALLe?I+74d3HX=O+-KY\)JR64[50XKefB:FN;@55=0NWcfC
0A3QOY40@XG+59&S5PEF+11HT:WbJQNgPH[cF]?]K(;Zg(UUCGAX[RGZK7MeK\g&
[T,MR)6RBP:7KRdPCNA#A1R@YdB-561JD)I\;2@W6:0fMRX.#.T.9[?,LeN6g&4Z
]YKaZ47C]HP6a1?cb>U0A?>]32@RI1)EVW>K&Q6[/)TD?g)J1,:IX.2@L]#TZgL+
V&=fc9fLMEFR)0UWAcQ(.EBLfb]M,CA,>7JaE>?<@6,,a_ZB8M.]Vc.@aKXBJG62
Lc302OVBBEDH@O5S^AMZMNSaf9VRDfD>#]SIa@+=R<cMAgdE(YD,68QQa2/AG1S-
42<,-I4]S0_)B2QPBX/6_O#=gVMJ(P#D,BI^^DNXPQXQ/]]42cZG).gRbe^1QK\4
.@0Q)UR_W2A&ZLM651B>AEY2F:Z0R]HR5WS9D?FS^,G1d:Tg6QK9]RNB0EX6[+V:
OFGL8S6c]O5H(M6W0.PKTd+bCYO8]N)Sgc)SMV2R]3EN:c:2?0.A-]?\a(+9<@7Q
Y@W#CJ40_KRI@bZD^^BaZD@1<;fUY9,9)I4O7^6IUD0QdNJ>OUK0b:eYK[N:,S:=
fRIQ-Xc&JCGH[g-V:.NEMc7-KI<2,^;e&C92>.8<T2UP9cRPDT=97b2g:-F:]CF?
<K=A8(4@I^1d#U[58THG@_a)]Y_6?#GKfRY^J.WJ2c9T8<QeDMfD;43JM]4KOdV0
_UX;QGG1<Y@0NPB465&Sa08gM]#GbY+[Z\KLYMITONW2#_D?9Z^OZZZ.]OQO&a7@
?].9;@DNH>YER68EgXCQGH7SLD9Mb&DL@NNIF=F15C&A]gfEIB->Q3AZ53^[,TTd
a]>JN(JO\)AU1G3)UX6_;Rc:\XLcU^76Zb]GD8E/W./fM>=_AfJ]=Z>)He2/5\@/
O=N8c[OD8B<b5;d/2_?&fYeggH?#5Q@-4=6e5ZE8N-M;W0N]1KG.\5O\AU8NP_)<
Z,Kg-X=[(e^TA)Y<BDXL@aC9=N<[ObZcMA;]b(4+Se7A#F9C\CdT8VaCY#2eSGZ#
<caL+T7<HNCCcNZ]4ecG4BWJO8X@;e@S6;U00\5GD2>B_dFEY,9;]Vc[L5;4X(f.
H;2I-Z&IVdc?=7E:A,M/UF:;9L:V]?40C8aX/KPVLS;<\#U,?O&0[de>D4U7VD/S
1EcDJ9(U7Mb,UG^)W9bD@,\7c<V].?12=JcPIS#OKVM\,SAL5;d;DK6F+;-Kc(I0
^3,GE/SNC3]d4d9R]X\RX)B/G:?S]]]b_-GF@gAK&=GfJV#GH;1WEEJK7/\a[HNe
5[B7\\;2<6@6bC3H4Jb5]A(_/G\]8MAP6@b-9fd;0<2<?.fd?-_:+GJ+UN;HO90K
:N0>g>30/T+:U+T(HfE)A8V1X:g)Y[K)?Z,cV?SW<A/?J2TFWQ+YUN6R;cgVe<(F
5Pg\RW798D(..+c\2+F]1FR]CTKgOOQO8B7,f.fQaJ>TA)Y;AQ^P6XBaH53X+,\J
2IE;eVNB1BH0gFM]&f>7>IE,G&)S;FJH_aV^_)60e7FN02&E,]RWB25;f8LF,L1>
IVX\E5SXGOZRCL1Z_[E3;AWN]F:JU&/J4MUaIf0DVXeN8ON#7XY+<T3I8PZ1K=[<
;8@/9=CG@D1Q__a/[8T]5HOK--S71;d^\/<YeX;<#G:I_F;CUX&d(ER,Q0@P]=.(
(R.I[J=30#MQf:bA4S65_@A[b6I^NXA7PPH9cQ>dZ#@CKg@bL#?Z-C-IeFeG@7>c
_\V??dY)1OVR10Cd@g)5L<SA-J_+R=bZ1;bbLI@^3.+&&#dMQd0geS)_^dXO](PH
U\J&O0Z.UP:304Df_F?^Z]6b=.\;5EUQV55>d5C^3:b0[BY_K,OA0/SDOZQf2B](
f=dE39C_;2aLg+R=7I6eO;CS1>]4VEec?Y2JVKL+0H8:OE1JEaAfJb]IHNFBNebf
fU2_^;?C7-L:(FVPX]_D=D0W6N:)RZ>>2EMKcVH,V)eOK6gYa:@CW]fPc20N0L(B
gCa;A6W6A5:;,&_eG_b=I(;V+,gU9D89#8>11<\^9#O8O>7D<7M9?aWU0THb3<(_
^bF&GE^JGU4RFBD\V)OeQL^?AA-:f^K79RH8#dMc9fD;ea4;9e@ST>QU>eG5GX:Q
#K.E+[=Ag&e:^E8Y#W,IM(GBb)(;b2<_^;@3Ee4b<[.Pgf(c&e6Z[=DKIda8R56M
0fdK#[.<.-M5RJ_H3SfSLI>2c2XK87,Y(&HP::H/e/c4-BK16PL=;\g2R8GgO]OS
L2/fDB)BOXIOd=d\(a?Z:]bIDD)ae:T&OHN=V5be&#^^Rb3@ScB=>:f>FCe:>1#3
U05FYPIL21P9FFVY(OD(-D(CMX_Td2GWO?c^G^5,./,/Y?G0d)B+a?),@gDY)-:1
W(1W1M&c=<L<T8P0XGG[MTeW3BC_B1JP_@D2R8N?FUTKgJHDBD.B1WVYB(+4NP@K
TVeI<,4gUBdYXb[],T:Xg&H6,(6;.29/GX9U>dGTQA7bT@R]2<AbSa5]X&_<^G>g
HL&UJIN8Z=J-A0&(dMHH)b@9^2-VA685Ac3M4A/e0a5O]Ha=5HMSG&S_KP4))OVT
52@b,L42@DQ7NYF-g+A9#F9b7K.@>&BQ_57CdbCI7F9XJA78P8&Q<ZQd7;5>/(#V
:4FQ1Q,XCCJ2g0cOEe/&T,=0:FP)J;=DELT<^BJgZa_RP,>dK=Nb4aLOHeS@?96Z
a^)L3R,BaVDWe&-UPddaO#D&#^?(MHf29-J6HYcU:S0F4WR>]3W<@b&FJ,LgOa]A
cc1:bW1L>eF#LRI7d,ZL?GYB,eD=R@gOD^=#_IJ8KSD2(X#.ML_D5TN]Q-_K>0cJ
SF^Z;Te125B[36FPP2:PXVA.c05\ZKN<[2[RK-71;K[Q3Q<&<_;.7g]I<R8R9,&>
Yecaa+W.02/NaJcE&>@U9>aG7M][D(K:a/8f6Z46=\.(,5^&OTLLHCe_8EZ9\;DJ
_8Z6E,9JMgLG=J,&?TH=LQAF-Oa;>WWR([Yg,V=UYU/1/V>+4=RX?eTFWEZ_Y]<I
ddS6I>99]Q[,8<+e&MBfI],N9-1.:,1J.c;GC+-L4@_T8N\]@B/TdWP\83/O2,E2
09.CI0T>17?G8I>(&>KPAYKd4MD@9(#=c\Q,O4J4a@<b?gCPWdX-1HVCZ82Me;8V
2FT]KaKA_DKIP@N]_T+#fPE973OdgBR,HSAB-;Gc(:MZTJ_BQ0[_[7&+9^K+;[LJ
?PcQ:KC8WcU:8E&aW>D_<RMc9<B#Y8a82(4Q6Y3PRZU6@,)Y&?F:/F;&M]#W:VA\
89aa.PKBAVKYcf?__\b;W0X;g<HK:<_C/a.P9=MKcS?BKI.+C,N7(Be+DBdT.U\?
<[\6Q1;=eJ3QM&=)SQFE1U0bIW:U4:HMR+c0\79_+W98cQZZ0+-<-F5ZI7AS8]UL
aFf3RPe2>XZ#R,=G+Z:^&4RP2RKF\?_(dS?7dd,=LU1_<C/:BfMI-/AN5W61T8X3
X,YA&@P^Bb3&(@Y?,JeJ+1-1aW8Yad4G-8(<.EDD-_1DA3NCXTV7-71Y94#DP4C_
#P8_Pg]<0SPbfJ)9Uc#(0/0TVbB=+EHM@)I[^R[1;MOHeKTC;Kb78<<-[;[(fKGe
PFMPR2eLM6=;]QREG?-Z[[TPEZ.CE1<d+L5^#N^,BfZSg47T2)W^6WNYJaa1b72S
ZX0C\EdTLRUC.[6>[UH/AL60d6gREV-;FL#6DK4X\b[-H_B>R3aEPGI:b^;]Q4L?
67a=S6XIRWM0#JCK3eGJE@]3<LDMV1V3XD:XI14QJ<?e(#&44L4#EeS3I(d4J36f
PS4R,gdfEOLL,5Q:6N--HNV7gb1#>0(>[1+NPZWT>E:-H,b(KW-b.ZU6Pd5aH.)>
TVLe_bR)HIgOY;>SQ9P(HAZSLe>#&3Cg/2gPIUcJVK02V^](B,T9+[@QbJI:d&cA
\#4d2HNYN+b3DUBaK.XbPG1YQ8O/L#-W9Z(OT)-fJTYG+4>\[Z,WLK:Bc=RPNZ)4
PM_fP&I,JP6MIa<MC[JCRY3?B^KSb7b>C-DPX\dfZ8T;4^=4W3>Oa5UN&[6gG9+@
AD>((7/a?SO0bI#bN^O-F/F[^HIDEEdAbZ)T^0/\+]^,E^2[ON+W+UPBgU?KW+d2
OI4=H?+106X<H7U>GU=?5]G-dc8gTIZQ]N[\ZBRH1K[MPHSR2@c=;5VV1JZW&9K=
7?7EMU[^K83M8S=J2CS4YH))6\[_eI=V3QU(0ZV/]3e(N>-X#[d^O=1/Q@BBIdH-
@)e_Tf-92E2gE&1:6K.b]Z1eX+bM38Wc3M<.B8Z99]XgFdC@(01,Y82=_QT_,9b+
_3)(ZK-:T@C5W=7,U12@J_DQ<7R(4S79[5(3AOMbDb)[+9Q(=U(<UH&Fe;@aY2cb
]Lg=\P70Q8e_)LLBQ73g>,>B-JT/I=aW9?_IFQ-DZ;[cE1^)b:>SPcY06_6DL_8[
]AKPWbPeH\\6ag#FBg9PTfF=RG,ed>?:>e)>>RBg4);G7,[O7>(9-6L;>8IWX@4;
658J7Pd-g)\bSFFQR9R0FXQ\B,)-))gOdded@>NB_=?G-R4@G:4Pf&Y8==S_V37]
0F:1FY?a2@XY8VRMOR&0E[@&>Ce]Dg:Q[1-VG>@c\Oa(F^J0OcB;TD,^<4b1C3P=
DUf&TF#8BOGD:__&B;3R+(P6Rg)7@U(<5,)F0[R.O\S([H#Uf4^LDFKIIEN\;8N2
W[b#6C3ZPQ3&T-U;,#b]6.@J;b4PBVa/&]7eMWIbHe>d/U.?f08AA\XY/SWMfQ8G
DeMDO,:X&T7R.-MZHE8^(-eN#C@35\#OXPU]94F)?#FNI0Q9.gG4R-acW.;CSZEZ
\CRU>+b;&\Zb,.9Cg?8<a4LY8OY4XR]Z502U)fVF?S9b4@ae?=T\IB^(S<)1?XT[
&#^]2>2G]:ZeAZObAdH=C14,:b8N8@9fZN=-C]X8g)U-:3NS1-[bYC(fY2(3fcVX
NXUf@NVM>_C.[@C&I3W?LX#S2cF6U_c#X?FVGQeNGR&O.Q/a.\N]NBHH+1#87I9J
QVID4Ze+0U7Z5FDG4;G01RCWU>5-AH=4VVQ&4S#90SQN,U2M^RSG4FG^D,Ng:XER
V0IU4&BRKOZ^CH#07]CfVC<M5F_3ZOM\.K+AV+M]M-8YZ<S[WX5BE3R)dZb^:LOQ
Y,Q437(EZV80F^3#]?=BCgec[H-IK+DL;E0J/TX@0XG0@:4_WXMVaUNOX>D0C=a\
;gH4KCN#UP+c][QB)6geWf5^>dd74>SfeE^B6c0U>Z=TE#_+5cV5#_4f70YW40/c
B(Y2VD(YGgJH3;@CH@50T^^@X9P7+7SS35YHIGPG)>8Z#g>\ZXI0T(<2eG9b2C()
f#I\3R^VbP]]9?9d?f,S\\6VZ3C1b<X,:<ABLXRPQ@SPQ4PE:H/:KcZ^KZ[f.SeL
IST?0UM_=cY;2\[=G6fTSB5Rbe6@KeOD52?D#=,ZP2^-+\=-IPE&74XaP<c#S2J-
gF?&QaScATS]cAdG&,e2N,7LH<-#3R;)DfP,,9:>Q0#Af>4DVS_9WS-XLB6Zf/6.
J?N.(_[#),eIYDI<:G?eP&316>fM3(b9P61?DQABQ6.g?/UF]7JTLS_8=U_,@@;8
9SN4a.b2CPO>Cb_,aWI>V9I7;17/,-8^_Y8P&^#1#(-1Z@60UbSQR7_7Q7,[)UR4
e]^SQDC-2-=fa:4_JdM0?e&(G+88/8Y_?a[N+0R60)L.3;@CYcB4&M]8bFOO(CbY
30<Wa/(37&D\S+K3a(G\1;>930ZNY:eQ=JTH?T[<^W&==K4C#=K,OaE.g.6@aA5M
]=U6gU.f^HFP@^RD38)^7AL)dI6&9e7,:)Xg-gP@+f:[MEG7TF9J0LH/<(E6NgEG
H>eZ^>?cJ#G=F7=QbO(/d/&SN^#6#0:.;^e@#W)S4G3^3TfX7PMdS[_c>;2>CN>C
F?4M4Nb[\RNe2EC]A/LE+c5fPAL#WIF3MY^M?<&#3P7TMJX:Q.]cd/[]SJB(KHIW
9/:;3?+Udg(66bUILM]ZbNAHd7570g4fOg^VL\H+UBL#Q@800PN3?.O5E)<RZ&8O
DV6.YNQU<MP/9F.]I3+C-8=:90>\VMUA2e2<I:6[-H[cAHYHU<J;-X0XC)B<VV(g
dW8QP7ET<L+11\6H)JWe-R)X8XQ\.W:DA.,&+NLL_f7,9I5e551&X[IKJFPOXXe1
a<b=CeRB<8FObL[_IX6^TI:BM.V#[U7X>HXM9@WJKgfXZ/F1?22b<E>P#Zf+eEaH
C6NS,A.,(4fR]7]6+beI7@b9/X\8:#Hdc[):eWU5?Q\S-)ac-Td[\PFIe0Y\PQ^3
V4.\8VE:5LOL_?dF:L8/fBJM-eU&+5A)gB6TNFXeU<<V0#;#DMXQ+L&?+&?cdAV/
#@@Z4Kg[/DJXZ^gS(cR_dVfTSWQUD;)\:;^LQ_RA?NRPS:@:HLW=^eQK##D6/dO7
+TgBXD9G7BI]?/>\X-I7A0eM:CRZb/_\GNZ5_TL^D5M8fC#FbHLK.QWN[egSMW2G
O99Y0/D>UbR?e22U79[+@&&:a#b-CGR[I(JDdf&E+c_5J(.G9@HBI3+98EEAdTb1
1bR-P)/?4FO?d)E6O/D5V#U@)C-7HOacZ[9QC3HAX<;2^C,[H.NPM]0_RFID;E1J
3>/]E5OH7(ZI/gBa5QU&^D&/3#GE.F=@#4F-5VJ9+4Q_?KX#WBfd^#K52>IL6LEg
2>fIB@-;\9Q=E^ESZJ4,29fX41&AR+/8F/]NHN3P[]B[ESY0+d>0:XN(F1FNfC?b
@?g<0RDPLQX+3d]LS75LJ0R_XC9K,?B0c93NgV9fUWT3L[2=IW_I3ZD<+b/Xa)6J
,3gK_]EYZ-P#552QGNX=)4S=Gd,aD[2DTTJKcfR&cL;<dI0K0;?+76]X3V5\eEfX
S_H22\4XG]Y=3eeHO0Xfd\b.OPZ2AN5R3X^;/))/g0AdM;59CPR_R9\ZE4P-PDON
AO?^H>/cT<]7dL]P?G=e1OOLU,SG>)]2+B[+cRRN3QKScf;?Lc?O=//c29Gd@N;>
0?V_f[.N@\U(H4F=>LgR_LR@P>0G1GDXVE@?&:QP[CTROZ?:QQ>eA<H_:cQ.+B31
XU-P_Z(e^FM?#T:fS<dbTHb)Y5YN=-;IfA_aW[SJC2/P3X@^bCeM2,4I/Ic^\55P
bR#CbP?^0HB5af/H#e?1c>(TdDbV6#Y##2>Gf(CZe<-UGSI^g5/H-PU5QDcTSO:(
HO,\G>0<34IAE(_06LW,eD(-99),[6eQVF#Z#4MYA21:4YHX4Haa9d66C@Q4J=/e
&A4Kd-Y&6_ZGGcK-1X50-#0P1:H\[P=MSHB2c/,FGWa.Za.@d;+WNIT?@@HHF<H.
R0@T/BMW\4C3g(>DFN&K^e;2PgY_be=J<?F.RL&[Wf@ZZ2[g/?,^>LR1ZU)cf#HR
+C8_d(JPF&<FgbC]FIJQ&5#XY6_M>>E#WWY2VV3)0MA3;:&Xg.SPYg3/)>?MIX_M
_e_:;eZ:VA88ESeL:GT19./5[F120N;.E&Z[>=XPfEYKF(MIYKD5\-cEcLV>.TG:
e4[c0F:aXCHX0[;@:CPa>GW,G5/=RL_Ae>Z0P=TDTf:9aT)Cd1(b4>Zg24#31CY=
T\6,;H?ee4,5a=EM[93^U>gDJ6+W0e64V_6E8=LTB-#5\1bR\:]O;<7F[+fEXN&f
_M\]dGL@ceYYUO]^9@f7793+B;=Gf<3DYbYG0dEX@U8K<<eWQ2L\eLJNLW6b^HC:
Y/ae(@:0,<=c34A[>(-NB;?=C1B\,Qdf/#0T3_#a6OIe<+_R>e^NK7OGRQNNH#6U
VCNDe[cWMTA83_LL1bR&Ea>[N7d?H(HN9;SbcRLM9&b(bI,6XC=LM=FEBWI[G+2,
1XCde/<:(aG/N:R5M;4??f04F77VRW+\0/^OSZ[GR8?XB^M:A2Gg_0N<C<PY)A)_
H:29D@6_aZJ(0JW[[F4O=aJWQU]MLT\4XKEP0dT)CL^JFM7(DVJ/BM?X0C,\1PEV
C4WKe016dKCJYVG]QS6XU9ND2S(,RaEJ?QJ55F_>7Y7U3g_Gg&P-9\cW4UWb.3@:
B(R5&3^CK;fa2BCB[&QO.175I-++G<-_^(?[Dg208YV?BKF:UKBFLD\X?Ab:\&e.
ZQ5_Q3HI8bP89^Y/99HE9DK>4Kb3-7CM<+#D;E>LH=9092O<E47eDfaM^\;88L:L
AA3BIZP8E<,QOGWd^92Y.QD=\&OeG&(eN:-B8<eO8U]R(Z#)8fSf<PR>5<]fC3d?
AIIBeR4=)b=215-_R5eM+IU8T?bX_3LZ[L2?E&.-WAZQ#0([T#5]MEUN^)BHM)V#
<3\[N-YP&BRbFVV1cW=#4(1aEBUTHD(dV7EEN::<=69THfNU0\TJS@.a7fecJ]VZ
C1OO_]LBcY@X3BDJb+4<D^>8KX[d.4QX/1<3UY[J\U)^#(e44b2\V:K7gJ82&1E/
XKeeQ?9,#4(,M[;a8#V\2e&cMUP+@B2K968@T</EA;QMC<02&P_V).]c,HdT8R(P
A5#KcF+IZe,B-M^/gXLS]G[Xd2fM(,\GL,a1:E]5W+]RMAX#1>,3B#A5V6U]CV-H
L=BK6CACEEQ;&/PR=-@3fX,;<)Ie6eG@SA4,5X(>4<TNUgA.#=SVaFM43<@MKKNc
3SYBNC/S]?MgX@:A7C]ReK_V@=9f<6OQDZOF(>J/)[7>M4f0]EZN;5P>4Z72YU_L
0:DS5?TJ2#ED_Gef</W^#/@8U2ae#.64[2L(S65.Za)OPI&SPR(E9I.d(><Xa[RT
CRVFQI(V7R9Ef5/W&cVJL-X&?R#2dGFYBD&N.Q04A\#^9]SE@85J(b9c;g)DS+_S
WS4OF@@MF/UOdN0(J[3.TC+e+E&V-_:;#V]T.Oc/+3_gMgLU0Wb=:]bR5@]X-8Q3
X((=N9\d@bGRCLF0WQ]HU=7-Y)DeOBc0#I]D.QaU3PN#KROJ.&7Yc)Hb0;D3b(^G
O+Jg[0#bB_SX;5IFCJ0;UMX?=F3@R(.P&5aPDNVH>K@=V\0>+<4I+0?#URSgLXQf
+?4A/E+85J_8S(WKY>:BYMA061#4TWMXUCLcNTeW^):RC5<Cb\fZ]MaGTLNMPdZA
Q(T9,JZQ5>SB<g>6BAG&O^B:O(/2YT)HTe;VT@)QH4QOf-:D@\)Ec)=8NT^GW8VP
)^GRB7UQ9a9I-XcG\\AK_B4IO^J<6g+-efef.=P/+1dED:DFYcAWI[K<J5V8dY&W
UOMDI;@G_D@@790.H1@2607gHd[gAODbJS3(SbU58VK,aZ(c@6#?&1gO<Ee1TIM=
QNKL\J)@G80cDJQG_:>D@W@+f6T)AR5\\6cI:R&18HDC\(O5+U[OIC)ff6Sd,A_9
ccC\8/?W^6X9?^gaI&&GCMOE>,42(6.UcGU[57N<RP>P3O>^eZ3LNVAM6V7@<E1P
8380RGC(BFNL:Ig8@LW00CS=)K#)D6PeU])FV0TFgUZH5+-g@;_>(8E2>JHE8Xff
)f4^XPCSIF/JIWXS)&a6B>g6ADZ]/0[FbRb0T00:@N^K26JH8UORQfI]^(.JeSW2
KB)NW&ag[8e7)b]@Y\KCgZ&a2_^fZ&^4H]&X?_A),DWD,IM0UI;Y,_QU:Ca@;QB;
5NZ71V/acg?@<Z6=Q]2A94;,@>_)e3Xd5@.2IW1eBBS>=4Kc8gLT42:6dg0_AVQZ
L:?\(AW8ZOJC3\--XFB47Q&bG46GbMd:F&;9,G]gRZL&Y3-H\AJc@ZY30Q1PBAR?
>gMNT//3Gg:R[ZgSAKSaLUbSWgRZH(LRB)90J4SH<K,R<#KF]5BW]CLVd^JX^2C)
Mf/&Ee99RL;8F>Saa#URR-3UGef\2b/O:LY>af-G09C56(Y=/5g:(I\XK(YSFR=+
6NUUgdM).8gH4NRD\;fFEC2>_1GeD?FD?ED.::63I/;<+,B7gAM16@&7+JS.&Od^
=K=:<b+B<>RILCQe-;3TLQAD6LfI3/Cg]cf<H3fGD-0aW_<KHR736W4dB:[K+\Ug
ON7D)?,_7GZHR&7&FP0F]Kd.gH1RWT[fZaKJ[4Q(XXZIF3eI&>>(U?bRCbU#OA:N
PPb[TOFR<a.KT2CJ32GCdZ&fD@1MZQGE+fMZWX&PL=8NM=@JbGR^Q8,A8>Q?E8<]
_:c+c>]1.c:OGK+VF<5WUNR76[.eV[\e]ICc3[R,/eLgX?TJ40ZHfKdMe.A8d6<2
@2=#>1Z\gGJE1WdX\V@@S@&/KW-WFL+a#6@;Y;Af>c=&M;Efgb^?33?K]_4NBHA@
aAXC68R:fab18V)Zd08ZcDc_[.2U8H\00HeS=\Y#3H_RQ52OYE[J@a.7K[JFU#OS
^N?#+6RaH#<9;?YeOG5ICD)(ZdZO/X4NJ;C]G(4G#C>@08BU11?P[<SeLe_XHOX>
a^1>HO=VPeR2]NMH_K^f=TV,B1VWVG_DCO.0f/>cOb8S4#H&EPELTG.IVS=>+e>\
/1^FK@Zd-JZg,?8]<,M<OgB(f=\NCLOO:]a>6?U.-a)V.U=)9<Z)K-U.\P6Xf&(M
/5gX_NS^/I,KG/bGY#KC]&CEV0WW.FNb_KUfO]fGW=\9PJgXBS2Y(8EWaV+f5(5T
J5^CHHTXQCDZMR_;;T.H6a>HX8bM.:83U?S\TBA?.a@)=5][c0I#@H>++:H8F(>Y
\TO,;dL-VW[_cUf/[2LIOQ/?]8@+gHRH:A?\@;>ST(+T_.2/PCEX-TTJRKa]\Bc6
(?XMUb.V>-NJKJ#/X&FTC9EX@NKZEdNa/NJU.f3_H/7;N-=U?+O0IAST)c6FDPLg
XH3VV7B2/YU-\)L\b&J.RCIFE/5BDdM=LW^4RASA=00E@\ZSQ][[)\WE2Vg<NXAc
#69N/Q95A[YS=P2W7IIEABIFg<b5e3NMVD^6eADH2e3KCdD;]V6=-+2H01I-(9Y@
O=SPS^11HD7+ZC72WbQC;:XfQ1VJMPX&d.dWd1)IMdVSYR>[Me(=4+d/AfB&8IAc
gT4P:5-He6Q5dDDc/)9e]cbG]1DYEYP#:<0I^2_XGK>4U&&(GZ_OOLgb>9<OW0Mc
@H4T#Oe(TGLM)[0AJI/5cSOMZ?4;,Z+ad=\>>aIO.PR3#77N2eQIGOaO#HZ:=&dS
?7BO\6f^\HMg_Da8WaPMbUF#_]F<5gAGO\+:+aNdAf^^4RA-OF#H;f<f2,I4CAU.
a=7UD#g#6#++DFb#3_-);<?A:.N;E865X0O;5-VFFGfXcIWE>\+A>UFT7d-1@?==
78FNMgQZ5/ge+Q3U4b=]QOL8WG?e17E(JKPAbL6W:H)3:Za,\G24;cQAa)_9]b2a
I72(HZ3aX@I,^&IC?c>.SNV0SWTJJ(5Z97(?50e&>SPH_R6e5=[OJDE?@A(YSQHf
bAeD3DW74V?N\]17>Wg,QIF(\T9Y\]:7d84CPg,>N&E&40M_ZEAU&fGFR0c7e_eD
O^Q)CKIV0BA&A#BV7Ae=TO2V.TG=FgMJ@Q52e:7J@>Ha>5<ZY,Q]E6?U\D\a.C]J
Tb+S53L2C>FYQK6gbN<?+PS31X)QECM1-=P++??/e&96Y\,&LBE:LBAdOM93E7L=
54V\T2G5VI+UXQ/d:\-#A65[^-&(7(JSW#+D=c1FAKZ:1X/;\18BS;#MD)]J:H7=
+-K?J\Yc;MNfPNEGIaC.fO,)9@K)(R?Q/gFB0\,<Sc==7BYa-UR-0:aS>RA]EEZ,
O@HF84N]d(a?d=e,NLFL>5Q]Q;,d:&,+cP4[e?DD4QOMA,8AI<+GEGY0=TTWcS5^
[G9VNK)5eJTf-Ef,GE&^0K^\aXZE^RP19X]MQF_]4b.O#WW?>J5WV]A([AXJJF3E
&7&g>SL9W,LITe)UdOXA@/VTdT._P0V7HCBHFK16(>3Q3OT0-+8+2Z7#69K)?P?L
0)1.M)(Q0bLKEZS3,eK4:;4)34TBFOg3f>Q^)^77gaM)MO3A5.TCXLeg1?+I5/<B
9?>O#YK2]KL2?LHZ?Lc_27)I^ID2fMd=DRGDaO^aI]XYWcKGcH\7c+8B.C_&HK\-
WJ),;I]2F,3G,P(_VH5-@BJ/8IF][N)1c4#4#SDUVPRB=3e29I.T@VSG]HKM439T
bYJ@C<dWXBT#La6=6D.GJ&9.Nd??)(=MS([K51^H1Cd?XO-<:RMd5JHNMa^62DYC
G+.8b)P^gDG#<E_cZMP]YAN=&I0QR6ID>V5/;0B^7R2CR=O-/<9E2.bMCFW8,H3L
#/ZH.\e_OO3UE@Q8cgBMP32T09[7X.GX-=KJ>>(#(&N#<;8.TNP<OG23/8U2-7SV
I:c?BH)5-;\D#)GP8f>9O,FLS;;EB))T:,4(Y.QV]:8GJW>[0;;9_f^V=aVXE/][
W08_Z:ac.9XZIK1(6#HKNOb+/,0N]M8H#HaYE[1\LbUaHVS6&D:D9-14;f4H<#5+
5K70fHDQdW0ER;W_]bc&0P=a(H+R,Z@68_#F4L<=L8Q:2S5PeWD+U(WXab2G0GBP
cL.b_3V]COU+OLb[##H20KcAYbSP;8CE[WKc].,YM07YUe2B+H;Fb.V++-XM>G6S
^TO2g=BU1P9LSC^[D#M#dWg]Q]63Y2PMgT(([39]G:]He_aB[bOdVgF:Y?7QIJF[
3/8eb\8]cGF3dYc]IA[cJCHMB6N.9MZ>9HU3-BM>Y=)^/[60)\f0CgD>LYKg5MgB
b64JIDKd+.;M/>BHC6KIU+9e./<?LMQ-?TIBZ+:J7SGB[=Fdb4dLY/ZBV9F2FPB/
J>@e_R/[X85b-#?REZKA#?/\C_Y:P(S-A72<IdUcL3I=#V8O@I,Y,<9.Lb#39f?G
#+W+MRUedQeZUHAd(_b96deM^^QHS)8&+69@HJaA&0K4E\WCUb\7.c6FNPGfK^WS
f<WWPZVZY=[0+(OOBB7c)RdD7S_3,+DID^F9bG;/T#^8M4.9?Yg@b#PIBNN804+0
#4#SX@?GbM3=FAGW6C[EPS1A,[Kg;\g:3OH(b3d#06-g[\T_BVC==0O<USX:O1-[
H&5-bQb/8B-IU+E7^O#BI8<f+=A)#108SISM@8c:(C9?Jf#>QT/7VFcTH-S/>S)6
e^+7,,35@?9RV:OZ..[fPO3NZ,3,W:/_5V;-b-&^F1WeRF>/?&KS^d@(d)?7/^EA
KIN#Tb?S(>g7bF-&@0L_Oe175ce4-B/:J[./S5.<\9BdP:^#M^G1O92J=4JH99S6
CZ-EaU8HgGa?&AcUg_U_C>;Bb>Z-Ka(+C>JXG#N]2B\E7./&,MNW4N(.Od_W.K^6
G;HMT]0Ba_&:3DeD0D:#>_&0Y]GF\GE8S)XVV)YI0+PZ.0R2]gVY7ec7X2-KU&NE
0cTVQCDVWb.9:&3(X,Tf-;/0?B=WFBYYc@^O&8Y\:-]ZbXTBdc4KG>gG,b)[SY_/
V<R#&CBQDBO+cC&KXIdPHPHJ(6XXSDU6Ogf5_cCR<fAf.&J\bBM#>/X@U9U-_4&:
>e1_Ugf4-&_11)5+g;YfMQ^6-#Y;ReUG?NJ49XGQV,8B8UeO:@?FbU)ZE0S=22NH
SNfEG,1,?7YH\Z(Y9KA]GW=-YE2OI;+5S9MO32<Qab8[,(D-bdQg)fH?/];bIUZ:
Y);8f@=3_P-,[GNMQg/dLZ)#804fgF@D@.GV=E5Ge5.a)7L?g<M/e+LDAe^,e((1
PP@0EA1K^62=F1V50Gad9-L/2JaK-41Ec^f.G\@R]551G(+O>_MMT9Na7?Jg0@b6
;-\URgIN-\>MRQ3;/6#0^]@OB81__1.6:b_D3X45MG_P&Y/@:](GBT>FW&dAadR]
Z8ZUgUIGd-/G@f6A_^._fRcSFOTT^H]/E[CETQ:?XOY6PD6eE,d<4:TgF0YX@9g6
S>YV.O\b)Qf]eHK/=dDT2Mc:H,8O_J?f>GVda,C3ZQdVaNXN2a(#5Pb8MHH68g.W
(4,H,-::0]5=CcHWX4eQ^LC>&US@H4/YI7A+Qe[P[\]E3IIO=T^A0,d;JN((/<FL
fb@L/?bR8TJNV;=J;[DTK9Yc5ac?X?2C6P;Ub.X8Sf-R(/I,/+C8[ZH2VCX=EJ]&
a@&LFd2_WDJ<[P_0bYCa[_(D1JXO;B8^9_Sc46+D]1,gNMaN<E>Y/:c^=P./DLaT
XHA.Gd_b?S8KV-A:X->_+0OUI/dMB<_2f]Z81=\A[2X7[+F8+77.@;AD4DD_=_\e
f7BG@>>0MVU?SAgU&.[>51/TaG\\.^MNd#HfGGQeHNbF4K@3+6L0T9PS<9&]IW)Q
QRS1I7LKBdV:SG]36c@aTASGd0PU8RY@.KBOA9cD&],QQ(GR4W]OP0+\-f0U]\0a
D8_8.c)AR9=VE&Q&EaA?ZYRDG9->,VPF=d.Q2^bDBRMfSD949&_:PAFD3e3?<>6c
V2X;V9<R9g?)^@1:3Z>BH=F?Z9@U>B)gc:/X&0S]<>EG?V^eDT?YJ^[&_BX)8<>B
E0(NCZ<XFC)[X-/;[-[7_:]5TMa:N2S=;6I6R[5ZDedL#-,94#GM2P.Zf=>I.d(1
86,_Cd[VGNK\L9^(?QfZ:JUM]N,NQK@eX>PYf/;dAAgXJ03ST=]MZ?UQT]=++P3.
)&=/\__.)B)X,^QQ[,IS4[.b6R\dCf=(OLMbC<cQ2D#W7<@[ERY[Y[[CTI<)8-e2
TDFZOYM/d\B)783EfE@gEYDe<+\?f74^HCZ&ZUYKSE;e.8\;[N5NH)3SUcb9d4:@
COT(0>g;LT?^8Ib;4Q9aF63J</ACF7PZVI2+FAJ<NF(^X;8.30&0M96P=<Fe5S&M
+LK#dK93M&eTR=&H6AO3#4QEC;D2Q?g4R6c3;9I/?TWB4_XZ8bS/[F:HK1H>;>DK
5MB=>ZL,<KHKQ[#.92fIa[H8K^T=+C62A+1aS5]N?a0AT]d6)+_IgVO1.21:]RB_
(P0)@S<@.B2;U]V3.,L4GAcbcIKIaP;/JP<?#[3[W<]5;=7]SRCI5Z3=K+4)AA4-
=]LQ5J)=fEC.bfQCQQ]1d>24d;/5B5861,TH?OXWeX3FY>+<2Pg6d4=ASDS,-1)D
bb=6@=OMTA?_)[D72KcA4ZIg-6)IRJ-Z+.J(SZF&6E[4-\bORDZNg>SXQR[:)/Uc
O^,8NW-&@NdEbfX4gMH7c99S0V15GS?YcV.C;d.LJ;>LV6Zf?(FYF?EfR[L;ef0<
b<R6gET9F(M9:2f9f0L4WSJ?Fb-=1g\FD/d-GZSI=a[):VaCI&G#CQF-K.-&c>_7
W8S#eZL8]A;MUGO_Eg#H51U#S+34<5M#JY:I^?eRN8W7bHSNT6N\[5C^9SR/GT;_
_P1C\K5?:B#gR(+X0;BWELa<1I79MXKB5Cf7PJ#aGddMHLdRUX7bf7Ig#/[EO^fH
N>]J(<KNDfB@C+7g7Yc;a8LLd+.6DW?6OQK^2W6N/d^\ULf,NHdW]Ha#SPUKWLEY
RXBcGL_1DDDS5MQ=S_=UFBCH6WIUV.JYW&(6b]J3_..dH(57Ib?61g_5JVB-U;+#
7[)0Td,>VN[6<F(3M.IB^3\97UO^Y\+?Mcea-F](1J>#/F)_VD:FJ+9S,-^_dH7A
IA:cU8^SHe:8eKfU75.P6c)?6e\O-WIDU3>>IHL.e.)Z5OHfI)P:9\O3MQE-WJ?9
dEf5O+C(WYIVAT9HU\#?XdEMLG)&S)eUIVUV(cS@0gO3dJ@Z,W#/>eO0LZd0[=.6
^I&A/5:S[d8DHU3>18?2KTR0DR;]dZ=0@Q:<_H4FUgCY?aADO)OX]0Q]e;))25H\
W:#@9U6La@XC4,_Lg9OE7Y0)<?)O=EeT^dUJJ13IR2(56V]AFXIN2E/./Z-+0[0c
+)@UEIV&E?JY5&b=;+51<,,cR?b,^<Y.d(@/Y<aL5gHW]=4d]);C4S2Cd:04F:<4
6IF3;Y,c,Y0R;#>Z(c1-8-K=GYIUb8BbWe5M,)&)9b;2db1e7(BNF+(P^H)dNg4b
?,/&@@B0E__5#1]#>?&:UB)eZONbWDYS9?50^]_Z(<B37.VE#DdcPaTBF?Cg4]LD
\P6T<\5g5[ORF_3DJMYb&3I,H7_1eRYKC:A_VTd-Y]=g:?gP.F5\@SXLXN?QYc@0
8f^GO5PKQG,BIUNa]GZ-&2gZK:[<ac2^a75\d/:YQDUG>M(1?PZ/([9_EYQ?6fYU
<+N&a?GU9\cW70b2LD9-1]#6P-F6S0AW33F4CWdbBGF_WB]:EA(=e(#c:5fA#56X
>EabWc#0)[]K?F;1/J:8,7g/9]DGb44+&83Z44bZ/\PZC8T3bR;8NF>.g(;J0b1X
Gb+G.]+GC:.ABb4LE(KeS?=@@OgE=a>6C5#-b[98E\e@L^1JAe0-P_L(=23F@C5F
6Ya011?GbA@S-S/H)FLg7>Wb[9;@HecVFVX?5C50YO3QKJ#fLS;ZBHF?U.FfIS90
[aZFc4PJNW.R+fI91cRbZ559J4cPSI8JfC5EVYb/?cN)JIX#3/1^KMEJBLV:TE<5
ROJY@Zf\\Y29QF#I.H@Z>,XaL2d.9F(1e?P);7?K26Efd[QcF^5H;-A\JD+c[c2L
YV>)bGDSW;SH1(\VPTa)9gQadKM/I@L86Z@KN&E+?),X-SFOSG?K)2(8<M75CHF/
PQaIO&68[S\B0\Db1Y_H?VMDL#0:TNba8+PKbeKbF/Nge&EYWUEL[YJ_XTZL,b[A
-geTG:3,a7>QRA^..PT(?-2C9c;[:EaEYQ]H))YRSaH?FfRZ^9g39=,G43=;^;;Q
b.eTB1I\^ND6d7/^I>&SH+6,5b7_8Ie5ZcDeJRUC0\2(_/d1K\=eG/e\F6HF6^8.
>=cgDN\geQ#g&)=KW[PD;>34c.W&.IKF>RA5N3WIZ[W?6F3<02TJ^45F_bagL9Y-
Be^Y32\Rea6V_f/=1B8IJQ/04LVId[.-aDe7.7T49bg\B6,Yd&7=#KO;BbCeRF=X
,8gTO5Ab@/@A1LWDdLfTf0J,7dF(_c6+fUI4PV0<1g#YK6\JP^<,7UGdN.ZDa_T3
(8@TSZ4_N6<fI3DR-S9JWOd[-9M2JUQB1aC[[0Z;4UL182.50=IEBLTg@b^2da+R
>1N,cHD(H<3Y^91,L4fAeK(3(:aR2[&J(<:>QW04T/4RI_4&(#2[WbP)NbD9W3U9
=&5a9Gf=c=OHE0CXg5[LD/]3JRRUCA2S:)=1#YWB,F[_\+DfDM3R;-_XSJ]feM)?
3F6(NbD>I,98-02;Y[@dJefTc9gR0E7V[^ZV1,;1bPca,0_U/6e\V/90/Qb]?.BZ
JRK4/abg68>@g0M]=cBNP6X4c):fTR?O<,E7W3CY0GQcJ[-5&07_;6Q=AJ2]^-;O
c3<X4-4Wg5\<C]8BMNV>^XHI&K3)gX]LJMXB3Pe=XL+&<&10@57Z]2U8Q03/2HH;
S,\:X[W@A>eYH_4-+L1/;U)G[4@W5MHHeS[DBBZO8C@\)JG-aR9=2CF^QfN/5R4\
T^AGTDO?H1EeSd:JM7Ne0eZ.3S5>4;FL(Qb,D.=Q2GK1:(=d=G^5feWK2XbL-QD3
]?dRe2^=&3D\L==LAU4M46NMA.gaHU+N?a4aO_2<#afWX0J1=aB6NQ\N),TX4W+\
M_dPB2@a])5H&OMWU+88DaVLTI\+[+8I\gJgX4Q^7A2b3a2e/CU@)]Cb+fLc([b6
OdL[9GcT2DL7JLQG9OLDX[c\J\1273IX>-:CC1(Y#(Y2HSQ8feDdP[&Pb\OW/PO(
Nf1A7X5_REE<ZVJ@\:GG6Q@bGQdbY8)I1:R3Hc^^a]EC9DI#.V(,<5+VCEEQB_TY
Ha\5FG7c3JX#>/P4@R+V4.RTQZ3b\6[E,,eU<U@#AL,dQ+O8F9AY,f1FP>VMO#Qe
G/9\7L2.3/2J+>)FRBJJ3B^.?[Ad,EK9X&GXeFT=HR6XT4SEUXK]c\G-5Fe?&_AU
_PDeF/KSK:gS[W;N/W=3cW9Jf1cg]<J0,Z&MU,X3V6V-P.0N_>4?UDA5J_I>eSB7
4,-XL;E7B.P2T-K[->Ude2IOOg)Z,IGaKCe+.F&U_S5FG]73Yf)7EJROYQ)5]/Ig
H#8_+,4Gf]<#0,Nac:_dC.2adB-E<S4[6Qd]FLUP@aK[3T7,\dG@&W2#-V<-1U?7
a=P8WACOA&+5(g7#75M&0NIaJ,9Ne4cK7d4+^=,9#/M9Y)B=@:&+dg5Rce0gd-00
)[g=9Hd41U1_/fd-&LGFY9GPKT<aGWGEZ[V8V]Q]e335L>SNa=.-Df)<dG\eRG=/
c@;bE6.5Kd=5W3f4K:67S;7]:G59\9K38PPfJ28(=)9<8AMgQM;4g88DUV)I<Ff9
fZD4#XWR.PMagbdPbbgI\d6dQYS6T3P-D<e<e<^C:H/4CbERC3+P0SJd1QML7NOb
NYE.A0/K_@\KHf.=Z]2YDfLSNOMKHM#V^+_R]M<b^E[^/O[R\+eU8>ECfc1dCZ,P
&3ZD7)^;9OY,=P^=7aU/)P+dc^Dd[;?HdW+/81.U6]aGT=,798H^41Y2J[KV:<HZ
-PY]&CB3[9D#7K5-#.abCBW1=#6EB;GH,+=,I798)>gDR]\PRGIS)D?N70NV<:BW
-;AbeS9F-]VOgaXX_QM>82A8]G79DU20d,Z-.IJZ#V7PIg/5a8Z>UAXA)1S;@JZN
ee.3OF+BY+a5@UR^<>1FPN;)2PN2FHQDE:GfTH,N_D(9WL3LcY#9096@VEUbT\R=
/LROR1g;#C3bU4gTWG<]J/5d8NLJ6fN/bQ<Z022g<P-M,a.TYN_ZD0-=FYA=..a]
cP41S;IQC9BVc7;g1LX??^Ke-6=@VLNSf7FMg+@EE9c7U/62e<PY,&_K.-LO<PTb
>c]dJ)IbSd5EN=RRBcac=CM0]\c#)TRZO8;GB<b9628W6\DMP)fDeP1S.@Bad>[d
Lf5Na?MedK<1GUeTHJJJJF6>:=g:6)>^S5-_=TT9/S,)N9OcMZGaYF@,JY^J;G^L
NKDRdUCC#.(V;]2IgefY)2#YJ,JJ2E>GVL3SQ:Nbedg93QR[CI6<?A(>bFZ59N58
RTg)GgLd71R@cT3P?GQgT23]0.6)=9MFg[XT)HcXE_/bO[6L2Q.\L@E&e0fAG2+/
d@A#7cc7I3Y;gZGEGcOO5E<a5ZI1JO=4O05()#Y@[GdYJ535NL\^X8AY?4IQfVg5
-)_M@XKBE9X=+MP?5K:TY.d7T16U.eLM]:Zb/CcYS_8G1+=BIbbX9?Y]S[D(<<PE
Z_,QeNJLH+(<4],B-,B)E(ETg,_HL<3O7_c11JX/585L;O&K&]>IIQRAU),G5^K<
E8AA?ZKZ^Q\Ag4c<O5C^cI761X:E#&WKgdI69<,8&NJB@QVL6^.K^[PM&03;;ZQJ
[d3OMP:U2PAXS<PO][G-3X=H8,E0dE5?A;F03d34RaN^<NLc?8IKA/2a.ALYEH5X
^3@SZKUC@eI]8A1eY7M14b4[8+]E_+VdXO3ML9=9#cQP3CfNB>6-FJf0YW.,RA#[
J;ST:;W82(UVOZ(M71C^;c/Bc1cB8b[9E;(c[S@WV=;dA&FM.R+&,eS\6^Lg9RJQ
_&1.Z#?X5)K#[6cg=\&;H:d)Pf_\K^:ddfc26&9Uc4b1U,<OX5X;0[7YJ^Ff8YeO
aUXec(g,UCgd[58O?dCV[BWI)O9H[eNY>I7QJ@K7B-/OfY2)A/(c3G^G#;7FNff2
:g#@9d(6YbA>ePSb4S7/BZ/F)P2V5.H>H51d2<UUDY/DW^<]Q1L.9g,K^)TPV&Oe
\</gPX#;5Dbb:aKM)\R-@;0<(ZeV^/+<Q&AE#MGG7U8EE@#4\^[;ea<FRReA9TU&
O8a@2S/d0L#6d7G+GS3J=c>Z)9aJ&92TL=&[.)3A=U8((VPKVM+6:D<f7]/)GL<1
/TWWIUO(6ME.VN-UIL^]6_ET+F:0I+X8]2U#<-39bGW--A3N<MgU^fBJeP7;De>O
_a;^]QB3V&IM.Q@XBYgBU.aJL8C)]GR/H4OYaXE\LGRX3#?457DRL(ZdJcTHDM68
?Yd)W<Y8R7D9\,<cJDCg[1e)g>O8CC&:U.d5>F:P^3e#VA>0(/4)J=fL))<+BU@;
<FA6QH_-d1F+7]6^M4^9E5JaB#Ra_)1+G0O+BKa8?I.-C:/A=E@7M#]1==d_<ECc
G^7__?U^45bOZ/NL)8ZZX+W>ba_V3MNW0R5)Sc^JEX4f:D+gQ2FU9UWb\eVccScG
2bV]S9SY47HO6BfS8O=Ze04XS_N9_T=:/e\G7cPc-ZJfFG_F-K3;C;VaPQQN(CdY
_&(?BdM/WYBGf89/\Zc<AD\]2T+Jg?E9K>5A8#9^a41>]=aS7B<c.R.=(GELVWTD
Y])1PLM94T8aS758CO/&G&gbWXD@C[TR\aKKFK-O5,R<MTRI.#a9L>:d0=_([^C9
^;LK+5/1Pb<NFU&29:)W_3+NV1C[<[XXHV5@9(T((gQ.\<aA/Z<@?QECc3<[E-1X
=6Pg;&U<^;eS4H.QRT9:+)MD[NOJdLaZ/3:2S@=<W49N1;?^=QaD>D]#aY/d6KV/
O&)]1g7gMd[#I\YeA#SCU))-DG_Ab?1J4^]\<X4IS@;X@OKEM.e-B=d]P3+Q28Zg
HN\8V[W7OC#F;R\[8Nd&&ZMGEFdH+.;J<@gLfX]DDN7AeFTe];Q8M[IS&gFM[[Z?
c[N;]=afFeXW;(O5TN>I7YS4LK0D_?1b1JSSg2>OZ[Cc0>MCB?4D[&#-3NX/d?Qf
)/M\fL+(RPOU9ZGDK\+R<QM5(\,6W<KF](26,;YcU7N=YEVFe:722:0J7Xa\KKBT
1Se]CJg0B7FJ8<A1_2)N@[d>2b^\WTHc6&(MPO50TGLWfHHN7L_-Oed1@I_/:DNT
L#_L6D941^-a+d..61..)d@7b-JfQI^SW-)+9FMJOYYR9b6;GL<0XUW2U>_886@,
-3:D5(R_P)(/03.Y_?;TR?5.R?\^S^,3_JIc9e#SP0&KdQ+IQ^31c[BbF[LT\<bP
MZU-JIeQU+BIL@,f=:E+_ScN.O&PK-(,_M]Z,Z#f1P;/2L4Z_N0XL<PR2,8Z6+(Z
0]V3;5I\^RQEe(G(C>#,&\(+a1AcLU+gdQDJ73OV_fB>17T4<T#C[#TVVQKZbZPR
XS&UL9;S^)bPO+.LK?U-E#f&-NS#67(5Hd]3M=&@bWS@-G<Z=E-]32R&AgfQP0.4
J#7dIZf6Vg,:T\>J0B6K+bG<[8M_.7RU-8fX7g=P?J,A2BeZdL^,8-EGBbE3G]=3
A6=O@?8J_H@Md2194D1Nf&;>Af2d(SgWT;KHBCfZMAbV7UaN-J+gJc.&aWa7LL\;
N4W:5-IfV4f0X0aeCQ/NBa(a7]BU]fLV+LN],4\+3ZK0XWfZSVY78XESc1-2\cU1
S89Y.a,Z/,.-/\8J2Zc[ZV[[4?DJ&#\NNLRMLW(f6/J>bDe>QeJS65CY#D,@4[+5
WY#&_+[Jc5fE+)(_\,/&GF72\^DDX7b_a;>L478<.Y6+OALXBX/f#Y.W#S(N8+?_
9<0FO?TAG:_Y@[Re(g5+/@?ddgV]<(/(QW.M3QcGM8/^>L^GP&/K9\f[E=K=HQg.
^6gAeA5L6]XL?8H6B18]K#T<(CB0PM)#9AABG/C_2Lf>#:CI-Z0_7bA;XX]QJA0H
4?6IZOgf&T\BB>TYO.dHd4I^0KU,f0b[(.:,-QDTaX._\J,1#ZYW\46&aUR97La<
@\dLPWWYeEeK;ZX4fag_?)@=FWUQ3#[7&A)0N]W8.eOA80?&AY#J?@&9<I]4EO_F
&(E161c,/Y6G1WR4XF:HdVSFBUNJE?6^5Z5SPS&bKFdb@6U5B9W1U&\a+6)_6eN9
.;UP98QENIC\a&:WG/)_+PO6[Z,-KaE9=KQ_MRS+Ag2QYJ;ID+a]MA24c2KULUY)
;5W=Xd<g&GU#\cFVCKOF6eL/EL<EB;V;>H_af2/J&WK9;JEE6O?]4=CecM>^:d=&
Ye,Y6FdT5>+V/IE^KJ8.ZBb]Ub4gK8J^5^\JJA7P[+Q.SQB_DMF^54=&VTII\PVD
W_g<f&2dGV@OMB2d^X/J42BG2d(>1UWNaeACb>]7:6/QIIEL@\U<Z9W&cQ2S03c1
5D5f/&[S3Q7bNXT^6Y]I5>I[N(<7S4HQ=+FK:Gb^Gd5XPd<fGE+S)cXMJ4/g5.8(
5]1MK22CbI@;W:,\PPY.G\#g1fYb[?<d#A4QO#YEQI#&TL42+;IT(Q7(D-:LXN9?
+>=3G8>OF&C(22b0.U31MPX,4142)6:5PS4[A,)\d]]VSKWFSVYd9.+9T^>[c>L3
CdVR:(OUG=K9>7WNK(M)fTJ#P0<eaN<VYXBKX>R+fXF(?SZRCQ<bO&_FF_V=J<2=
_@_UEH)cH-O&5[INMD):@Md8g19SQHS=b7(^=^Ue=GQQX-7PE6XV-6EbQ9@UEb3L
+LZ8dN(RG9eFFb+I.C6;HKX[;TaPaKcaZU=Z40=?cGS.<Y+Z^M-6F?Y4DA_(\#WR
Ggg2d#Ff.SgF5X/Z4CQg+Ec&ce(BW4CYaI&O;9@V)]=,;/V&YK37e(5;<QKgXfCc
c+b>+cO-L#I5+Y(<43&]e--[FbU,KWH^O&5VQC;aH3eYQ)6WZLMKJ6/;>KMd,4U;
W+\V+54fN#H[,H+YCIAH;^0X(Yg#dQD8N1WABRe-,)BbHgDV3K>74-U0aL^:FKTf
?@I8bG@\BX8[aea1Z4=A/KJQR1;,,0ADReFB]:QYQE#-QP\BKTA2P=_LJd]?]fK]
aPfY.WRG@Jc<8(g.:6:OM@DcCdE\3HA\6E-AUd2.DQNIYZAD?fX)(7fZ0NCNYOeM
?/Z8P#CO3O0R/Z6L4I,+BTa,T?&<eZFAUF5,K>?=.Qa(-IMdMX7Ie37JJCI16EL6
TBeQ(O6Fd[(F^CEgg@V-fUObER,a@8HOb>5/OE^P/@W[1]#AfSL&F/YIfEbFV4,c
9:/[@D^V\0bgX:I\.62YJP0]>SG&@OE;\FQF]EHYe58V.8#eP-[?HT.K/2L964CV
d(R6EX_R8T++3K7Q5P64QX:(FB<+<-MVUbf9J2B[<&V4?-=W.AU.L&AdGJa7DeV#
>+9:(Zg<6BJ.[CbQXM=OPU;EL0JU-gc#cM<J.=GOFP4(MU8+G@I&df.dD=SC>XIS
PU+>0(g8bWEE121^cREMO4EGCGR:+(4EZ)M&DQ=eL+]>5D]H]=IB-.&2CI5/:\WS
;Q[R</Y^P-Y?eY(66CX/&Y6SR>>g3Y4&DI1Xae?Cd(]L(H6;#6fGV0=+GfbGM4-[
W>E+YgM;BP-:^<^ZbWC.BB@2[(LVddWV-]LKSYOVO,SOG(,(@Q:e3\4T/^@-IfC.
?dF232JK]a<b(Y,M(@VQ7,G0XV<(,\eZNgKVH38H+Y=[0\S]/8N@CeXfe#1TVH0f
UK9J7,H6SMJXQ=Cg1[)cb/LK4];X#D2779OV,QOaPWf];30[(+@9\PSH?;L2)9M5
=7]4.MgfU848VMZ43UdQ-(?7?WHaK5cP2Pb_SbU2@9QGWGaDY7OIFXL=01SM3b.B
4+-J453g-\DM7&AL[3X7<e[@^U=TF[Qd=PTQK.C8W<+680]a-8.\^C.@2C^^FS5M
FcU235Ff0bZK;9UVFdOD?37@ETUe+cE1T>7QW(HE#)XQ\[[]bd([gT#AcK0:/T3V
U-&^.&T/cJ=R[(^-a@aS->c5V0;1EW.X.OXB4Ec^I+L6bg8VSA#DX8=UO/N(M7T(
W6Q<>L1=S6HO^YW0Jg@,O+7CK2d__^+D\(GTTa?PN/fg\G6EHT)A0-EII>HaPS-#
(^&#:>)P6OI@&6\fOe>XT-K??O1Xc@eg4V=40TcUg2]N9]LL(:GVfd9NY=/2+6fd
BF(93A.8:X(>(9K:X:K=,g9[WGFO.QXFT3D58_?YSg8OfG32QG8:+KbK[bC^;1GQ
?>\0<8#PLUGKT0Gadde@\)51;:T75T[e>b=.YS=BgA)aBa76,BF#C4;[\YG22c::
F@L:V6><TaH,];14b##4VDUZ/);BRK)65a[aOdTJB,c?QY)fCY3AYSAgG_H[;<<\
&J\d4N,DPI[d0)&>T3;&fZb@>g&M(@EcH-U,),[ISDW#8YcU<.T--<CNRA)cM@[P
^:X3X?).a,OO82L(YMR[-(\.)BVGcBE.IdeG#E@[#=/\Dg2CM#&fAHZgg9QE+:[-
O=.NRK#fD,28T1>7UTgJMbDaCN0<WfKb.&B/1[V=,_3D81N;178<,QdO3V<==;Qb
7VZ5G,B)FHV1gO&Md(SZ1d,+]3>1\?c0JHS]Wb#HEG+9b9N#]:_LVI696K1E;35\
9dUdI,KBGR+VPETg>AYbb8XFV2F&R/73:c2PR<V^=;S0L&#5.=8P6INV&&OZZ^R)
&TJ^1:Ec_1e7V:W58Q02gSeJ[.EeJ,:#8+1,1REVV.TK<fC@KSI5PXDZRfGg9#eM
,_3bR,G54-f?E/FX7^]O<AF3_aYB@(/bOU=</:fP_9945c73aSGU+^C\#NMV:<JU
<[-;Yd)-.E:I2EeF[PH3H[&2C/0gSYDB#c@C8;]F)A[BQe8K48AI8@[fWQTf8dI_
\I&f0UMMK4CKV0?UZU0U[&-8(CaCH@e=ZaY9eW+AQ:_(.+K)YB.[T=NgYWI^]-JY
\T5IU&L?0VMO,P;\.ED,][O8/f:e4+#&O(d4Cc>P#F?d]=.GfaQKXDBg\#2\CeQ[
>LXCN:N28))8I)>H0?)))>Z/)gF&._a#f-W/P-D\5IRUFWI^0c_F0.OTKDUdP6/L
:,2MH9DJa#]\SZ2WZc58JP/XbRAdEDVReP+&56+^(<\QV<5gF.IQ(<5K[@e;:K7<
HMHCZL9>7&0GA<,9gcNR<JaS<3#0FdT:D@)C/7YOa7-JYF0SBF#POL/9eBCZX-b:
QY4+ZHK8D?B3HTVLH>UUSWX?,&d=LT6Z9:0Vd,:CG,^>Le=,OP=+THCfZF5=0_J\
b?cBd61R1(7+3b)X,gJWW,^[7==5)S@9]OcU&M&>3WG]NN)aP<P9#)=QcQe#\\>N
ELQbHgRS;EGL[TQ,KY=@V)0_\XBLd:UKGA@H^@FXNgXLIW\9;Q4?A=40aQ_c]7c=
^4J7C3HEK_5@.1-#;R8.M8d[-LJYPJD/&GWE,HGE#EY-_#/X6HJ\DeBL0^A2WR6Y
Qb\L^#-W@><f)?4/dbK.dTa5)&L8@+B6dbcZZBK>-E;\4c#PdbJdA[NYHDI#Y+b+
PgbG)@V=Y&V8Tcf0^+27YWAKWL[:#PY(?D?B?dbPPQKI)@-g.GS1C1:DfQP3)bX[
Z6cWVXccA5CY#&>VGUJD21>caC4U>:WBVe[3JC<aEb6Mef8SU@^;39HcQTP2_fK\
g>ETfBTS:M@=bgZc+(E6WEN^X)=XQ#,Hg0Ke2Z=2EDe;R?4&G1f0,DMRIT@R3B9;
_4F:O7D=cdLP(N1=?)fRDN>/#R4E)ULg_?MgDaZ]QIBTdO)&\[NU4((AY(-@fMOa
f/0D(R0A(EVf:\[PO1Xc#7^b@=>_?3b6+DbEcL^3W??)^L1f,bT-+[0)10_U\gfC
4:Ye#\Q.V=dQ6f5H&0V19)SNHWKa;aGY+GME;FN<Nfd7+=5I>6^PSI1,fF&GL&E.
D]/)F4DFUU(.g)?T0TAD_N(0aM47]B4)XU.(N4@;b1PD,H+-OCLI8(F[6W]b;W<F
Q1,aWA37M+4H]>(,e<80@a0[2[&@b3LY;&5Cc.7A/9L1OgCQ[#&LB_UgZ&3<RBKa
=A924/]U5K4g9BQeI#1<^)+TddY/3@8/;+MNJ?5M&LPDDKXWA?aH(5-T9#=W:Wgd
GKGAQ&6_J.884Mb?Z(>ST4/BHaAS#_?I+JX&1X.@/=DU+fR9610DZ5G#f;0E&,6-
DF8c7de0d9a1bEM<QZL^(,M,YHcA)&&8.+aUYa]K@(0#<4IeMK;0_AeKR5D=_KB-
7W[)&1QKTLcfQW33&P-?6>Y1SX.#0]/K#YeL.d_TF),)YN,03<af/54J6DOQgB^E
T5<gDW2]@N]Zf]]N+:<YXG+bEdT/OLW)0HGd@I@ZNeR4\c-74_\U-bQF^(IV58>.
IfR_dd=F\#F;J#b1&fe:c-@X25CaY;.g.c853E+-2ed^SHUd44eD.9e/;MF@FQ_7
GYH#V4V+2ZM@#XB?+2J53&W<<b&]C0X_YW]<UKE.cNSZ>4XfOH^85<deN0?K9Y+4
5dVHNH>TZ@E;N6gL6LW&(459>II]D03C-<^;.:V2JJ2WceVU5&\D,b@L#9^6KV?M
+f@52cQXJg+c9MaD2]=K,=gfLJG\BbQB-]_G8PMMGG2aAZ6^PDCMXW(fR)dQQ&fL
0S)Gf6?N:^5^^7_,:1b]&IB)X&9MFWUJG;KS-#@@/Ace44/4DD52L1T\6/D[JA]-
7BWA\RQ[BQ-W?6W.(DG#X(I_OJL6(g37H-JT>DD_KgWN?E.3LMXVa?NHIL;I0Gb?
af-8:RB\P4)1L63QE+;\((MBF#dAYL1+(1,HAaIcNPM1fOVM@T[P6d<d^:T7?;@.
=&7V4dc]IeV:+DXK42_1\X1d]X+,]G+/]GdBa)NOEW9(X_??.>RJ<ZRCb):=TG6[
?#eI5D]Ob,B39dELZId2_UZM0]<#DU76,0-fa@T&]ZCQSWd7aWIKHI@:R(N\,>_F
URTb/G/gLY>K^+R[J\^>&:S7F[ZEd(?<X0db>A.)bF^_ADVE\2.GdCdP7T9)7aM:
O<AVB&B]QA+^67WTM1_aBKNX=_^dM\J3UaE2:OgbUQ+625C,.GXZ5da\ND9J=Gb)
C??:>+<KC=R4A<?\,eR;8><)OIY2^J4NB.)0AK,[fd:?AXHI551bPQM].c6CITbI
CE8)3>&2Ec>&MLB2M0AI_ZG.V\OOFbU6[W4eXaY3LDHHSGEK<]Fg1a;SEAfVJc--
_;HQ>&+^,g+V51\VOKIHC@d0><0Jed8OAZbC,N7AP&SI=c.3G38\]SgO;2X6_.F6
C1c6GQ_JNHM259g\G:96Gg9&I)JNR7dA8-Q_=RaGT909<A0J-=DUN\&R?Sb0<9NZ
-IERR8[bX6=PUfCFC,U2E8E7BXES4/1-R4e8]]#U(fD=f.^SMK3Od.XBF(7.Hb6_
\#U,H08eC#2[d68265@9Z@7D7AWPD]?/1F1HEHC&#^-05]/5IBB@[LHJ6OY6<EZR
99bN][5L3CdG&8S52.NEY0@CbHFIF,D)K7BBDXQ.)fY>e2F=4@>BD6JbMA5JV<;W
]K5H5D5=++_/VBP/)RSe)]/E=A2TT>Z4N3N-<EE-Kc;N37a5EQIT<W[;f3RHR?MI
O\U@PLAARO7,0RX^>;9;Ga>R/Z,&9N/WC#GMNJ3b25+C23Vg2KUEXJff,=(:R;/[
S+N^Ea3bWEWD8IBD5=[c69R1cQT5L2KfbV5:E(.NHKAN=21_<?3dQ,UH72IHB?C/
eUKU+PW)fZXL/>XI.B1SM0HMERbV@f_E-aUW]\&aZ;&6/HJ^USDPc&EK)L3g0YYQ
6(D_3:)4M;IP974+1P/O.]f6d>2f;9Y-(HA8G.4b&g9RX&KAaOc6?ce1_>OEE2W9
#;90C\5:JT>H3]_1PXaUI?fCU+0SW:^^bL_EJb._OX?FG8I00MQ@.0<;.aC3[<];
0/F[]75b?QMT#8YN?YP657:5gF_,<A<IDQ:?+[_[TS\/S)F9\OgIX^@-[25]2JTC
3C,af>5CWe/\#N(TL[A/>LCIZK#-@-fSK^_a?G?]]#fEY2;[QC?LbOZT9ET?Le]J
+J=<(+NGEB@30V,]_I#3a&cX=_)NK(3W9cD[2198PTfgZEcFLD)B1?57/=>K)9:\
Y7MFVBW=P]<GTO[^G))Rf27#[e2T?cY+EQ12#?7gTQcP<>;&+S09d/JY]@PSFaAN
24H\Q#-VKCR^AXOM<UHg\[X5?A_SXCU[89A5Pc\O.,8F(45;AEK2#V<RN4bK.5M2
dA461QE[bEd95A@S3R\51M:BO97[2]@?9Nbf_gRbPfUN7-A-+U&]62CM_GK6@\@&
TVTS:A,G;8^QVF0-d:;.8B:]#1.GAP\)M:.Q?Z-:1P\FL&N6#:YH/XJ]8&A])R&8
>?1<_M.W^=&Z9]F5U1^dI2ZB9GYR#>.[T_\V9=1:RL[R3]7@,B]1RICE=]9AgcWK
7RM4?[bSPOG2KYc</=^YA^[cKIS3?HbJO&7XY-3f\<7/&C>&_/N?T5F=/cbMH[WD
F=d_Z)[>9LAPB>Z#R?2W?Ze52+):LLJA)Z^?d0cS<.S6C[EI;@T-XM[W&YQ\JOaJ
3AVfC-?P#^b]XX[<\3Y&I:?YM;\O&A:@X=7M1IBM^W?&+#Q;-(A>H3CaJN>X7gY^
Hf8M.+R1_M6bIKfA7d8c@eQCP8?YQ8=TJC6VHg_^g5SCbJf5DB/7JfSZC+G;@HQf
VA_9T+&&A@J^3[CbS7\C.I3d-\F+=VeEG<Zb:]+c]+C-\[fK3<0EXE:ZQA#M0F\/
e@56<c#Zg>-gZf.MX_SSS?\0I56M(,ALfV9fDK@E0HeA3):=]PSOMT:Hf?XcS^3]
6e8V9g5=UbRcGPJ4R^^cF2QKM:40-:Z4&#?bfKe.E_2aX;MF7(6ZMEb).P6EYXTf
gBC2509);dZLXc\C&O;)>)O?=SHC@/AH[g;5VUK^(N+,VCTXR;VNJgRU,-A&aT<U
1aTeXd^d:#ST[f3DCe9+OH3=OE^(&ZW,MDg_d7+O>022Ka:ePCQI<CgUCg2]F#Qf
#T0GQNXc;=@)W6e[4a@M]FVd4XYLT=HcG\]3@NNX.2WG@G1;SO+[KNTa]<TMbLZ+
3FE?^4[G3<(U_X:+WB+>^bIg71eKJ=.>B8_T0LMa1:d;ROALTDPBO]0^_38+6=I@
BZIG0&A4dg2IB?9fU(PbZ]AN/M>Uf-Q<bMRMBIf(?N1R2Y9b(:N?J/c-BEMY^]c6
I<?;)9CE?K/\^G5[W&I48E3\FF=/dF,H,He7(7#Mf(2JA1K([<EB66f&<2IF=67:
(PV[GO&Y0ba<,@KM3DC)H>KO3NaCRF&G3.e<MR4[+=TP<FIIaLE2-Jd6e_?\CfZc
7M448N:1cGT;cfIeUDIU4Jc=\+CFSS/CX)#+ZEZ.g.O,>f)g5&LA20>R[21VNOFb
RGGFZ9+5+YK?CMG1TDAQ,4ZcIbJe53,EU;Xe@EFBDe\9]RF0;):EHK7,&F4U2M.[
9);+J-Yb84EX+[TWdfe1VCKfAD.Z3c>IeOQB_N(1^G+P<P]a)#>IR32Y^^XbEFSC
3&&&\-J7FfI5/9Fc(+)1a_=3\Z4Ag>aD13?^g7XG3O2^_;A7117JHDOK:P2X#,Z[
QA^0T2V-f-AF[]Zg7PASLG4Z,7.+>&e(Ce/GX]>)1-LD&..P,c_9<1d<J,P3)gEN
SBCX9cDY3-c]8XA-XNdV@37>?\?Fe;5-[7]BGND6@U_dc+M=32f-Y]aO0FfagVcR
\cNWV3[#2#-&38f&J[e_g7H2e(<\I2&/CWcOSM.dFcBa/M_VNOY.#Q3X>]W4I--S
[)A16_^[N:^0KV1R5@;4d@1Z[\:O<94JfKT7.9RZ>EZ;\TM^U,Ld2&-YC.H;AGI=
TF0f(\KPL0^]:XJeQ,VaK:_b=XB9ZJ^]1;)\BG7cFg=[J#>ag(.)922dCMPa_[8@
G=E?f+9@e4C0D-=VQ=aHEYccIMT=RP9RC.-?6\0MP812W26b;3Z-YN(WY?8b;Jdb
aF_2I31dS)7E4J<AEaPd?/&UfXgeOdEM:/;?3WcBJ;RM/I-ZE,\P+#,>;72CU\U(
;UEE+dD&?G-P0+L84(ee&]B=c0)]VS6Ja];K=]V8N2<e^gBFFDgOA[IBLA>4Z6V^
GeLG@07UCU(c/=8Fe0d],N4<2dgVdSJIS^/f\CJ>fF7-89R::>UN3TcJ-7JWWf^G
G8JL?_H/EYOSZ><)C;^_\WT@FZM#/eg5eH4cD:NMW)CVE,K_M53R@@6C\Ra-c\+L
c=G6G[d?V5+fL-MdLcWVR.4):DH.eB8@V\=(aKV56E981HHXF[]^=2=M=7+)?bLE
QeA)bTIVK=2=.#O;[ICR)CZTR4;c(T#(<@CKbKN@.M3B>XTO<cLPK9X?MYJ8Oc]R
WCYKAVKGc3C[f\L9(Ef2;)2G-=AK+Q>].:)aT2G5K38FO+=@f@B^:W#X0X0#)S:>
_N1?BE_KRI55(@F+Nc0(?Ob3aT<9=c>I]?0;\YO&6VA.9f)WO/44#(gI-0+5EF8/
WTf(?J?70Z\XI<Kda(e[FF/^RdN(f=L(f.M>L]P6,=,_-W<c]=-C?KM:#;2)(_0O
>=cb,F?#8:@]9NU70OS@;YR.ZAR>Q<FI]E/dPS,bY;Mf=0c,-MMF\)W30E@f.U-R
=5?gC+F_^9bXPVgT=_#U:6>G17+I\Z(\1=N\PCQQILN)F4+HgV]D3SL8fP(3?ZMZ
F-,?Te7S5KJ[RbZ(5VOI6F^<7c-A6@aGDUcFC<OPd@Q9G_YL872K#R,[_/R6M05=
8:H7DgQ3f,I&GN5;8YI-MKB75B\aRY:)L5a94\^L8^Q^RWU)X\^cK>O7:]-4E(DS
3L3QeQH8Qbf(XF@&bLDJY/H\^\1=H7S@8QVdb]UJ?YKU]SAK?.PV2WP,IIC?3=<5
/7?\0:SbY(4(BC1<3+):dLW1BbR\KOF7I1=V(+dLD>ceZ-5Q;L:D@\QRbZO:g\I2
=P2WR4M&1L//@aJ?&_O@0D4SbG#T5=+ZG=&O=RH]ND1TBO8\P)-Ef(]_/XX6gW@#
;1B^G6?c=gf8WbRPQ8B]M&2L;T6684Q:DNY+K&^=cbSM.K6S<R_.\KO-L^;gE8PG
C3PQ(7ILOVD0A<C19CDA>VTZD8BD&T/<N7Sa@fUNg=EDBeF+I(dRS-Wc0K36+IN=
<-14(1<W@<#E)?3]>Ig6CIYFdcB33&fP]Rf@6/,BHHH4<a4@V0I7<+<abU/HCU+>
=?KNUIM,.ff7a]B6U7g>@_]NQ_E5S_R2N7=RU;@GVeLX]AXJ7-&9[WWLH-)<KM]R
/JXZ1T=966V#b4d>Td>Nfe;JITO<^C3OS_=C]/g^DE;WYY3TE4Mcd16./=NBGd>M
gH>[,385ab422,g4ZNV<05&2NC>Z)Y>5TMZN]BM:5RSTY_#a8X&Y=S7,g0?T=<8.
^g08+2&Q\,d)1RGH8f>PB<]8,T+/U+=gMC:SI\@EMGZUQDea+8M9)7.Z&.U\@PQ=
(Lg)?AVOWBg,NM?X4D(+OM&M>>cNUcMP7\8Pa=\VLE^A1YDR37C]X>c?FOB)5c+W
&UUG.A@<9LdJ<(.O:6WVcCFIeLJ.U>2c]b>XNTA>F](U\N#)3)VNGZLG,6AA&7/V
=WV;</C3@,IffXQ#(B4f1](Kb/I(N.@8:TK@7_SSU>_PJ9ZS\I;QYGQZg76&0,2L
7UYg7/.1/4AdLSLIFVP@2=E_&T=TPLaWNZ_@91V?VL:&c72_R,@,;+J#B^&BK<8@
;@;W=1?2dLFH^F@()3?eM</R@Z0U;.WbUXD96^GK9O]/&0\FZL1:8EB>@F2]F,B+
,622HAY]O>:?[OZIZW;&5La=1^-G3@3KOY4=^;L#E>J;YIaC[c\#UTR:?IR7&Ce9
JTTOZ@EDPRL81I_5.L1/2X>_]?13&Lb8,)Q;FV52>_H0VUad/ZPeNT6V,;3Z.XD\
ZB\:4f_ZcO&&IC6BYC?gU]QIJO:5IR<dX^&ERfg+dC)cR9U(;g7=A<TMZGT=PeR#
GK35P3OT>dRD=2N-WERa^fF_bad;RgNRHHM+TgN]cX\9eEN_OS7Z;Q4Z=bD8N8JK
c1M)TV^XJg3TBeGKR@68+&F#<370?O;4I-5=16#Y<PSVEZJ4fKR(,_KF,@?<Cc98
U,&-R9^Q+&6C:F4=]R;J=:QOHG._>/;adNTV5@ZBXX9,AX4a,A-7,#,<JBSQ6d1^
dT\FX[P^0#-,bXC31=)WMd@aA@(\\^Mb^M[NLN+G>^]HN)/95>L2,Q2T[QZ_C/OH
>G&25P_DJZEfGG^0df&7-.dJ-3/W\=OJX6YU\S-9T#G.SSQ5C\QG@/N@L7N4L>U3
SgWg\PUUaL/?^,0D^agB(N>MXEY(R6<\;+IHRbAP<5g-d4f(2OAO]_RQ,<CgI^e1
2]RF_0;FZ8FA2&-4(C9Tb1B8@DB9N-K:/EMFfEKE>-aL_2,=&IK&4(f>..(863(d
3##_>_;Y3IJJ)FSO<>VPS@3]?Z#L;04XdZOFLV@GEP:VaXI4K//&F7QR.aZd#Gb9
:^N#UDHa&&F&K7S#2I7SEF?9STXeHe:X^EANY3X_RHL<(&^5URTC=U-YJBJXdJ.6
O9=N#<MbK63M.JX#XTf?M4LE.aS1VDM6J\b<O2X<#_0OKdSB&7XKd=.@61]Kf;JZ
_S=M9\Mf;3/DG.+RJYJKEN3OZAJ9]GfeK12/HZSNE;a>C6e(a06BDb_;RMaBNRAQ
:XV:,)W,J6+KJ](R<Bg<O?Xd2+X;-)UB9a-R,A_EXH,:P0eCJ5NVNJ62\V/dJ><G
aT5Jbe1B/7e5W)Rg0TAC5<gCI+]J#WCJCO9YfW\,>U=-<)^1?)ANV^aD)3BWfOV9
c]NP5)DS0S4(KE?(HI68B8\BJD=,V)85H?S#GPDMg_f(+[@:I]E+JSF[,T.W/4F6
ZJ6KBc^72Jg]0-Q+KG)(FP9VW.8ENK/P+XBO>(5QZ)9P?4H(9>WcNN7D((;J\[H1
&4bI>2ZVWYQ4UaO3e-4P=Ea:cP+OO6UKYS[C\NOaPT_&b89acR#NT&<[cMIB[JBc
.<D:-55E3SdJZ^M3YBMQ?7d/(ddTgS1f.+JXGU)f.7V?5/J[(de(TFY1?R-G0G9Q
8aC6.B17=P]M2ZH=IX)6J&,W2).,4b@a-.Y9A<UYNB[T?Abe_VNCHXY1KFeC7.b3
5:J(_D-fCF;6cee&O^CEF@M:I0I_AC<@/+)1+Z-=>NI[fO9agZeI5.O@TR_XNR\E
/3_F#.6&X&#]A0?DG9ZMRFa^2SI]6YfY<2ANO\Rag2+N3UIg6JRX.RX(0_4#^V(J
V&9\]FRC&2[BP[QC+K4?@)f5d)#C)0dQ_0GSS2_B=1A)=?YT)T[8/</P22?>Q&\F
(&OVKggVE7WKSF)Q>^>I<bNb;=@3J.L2RHP,]S7/[c7#]_9.9QY(+da?Y^A@bICY
UCBb\JJTFX@TF.g=DJGWN]51,7P]GX];HbIX&STSgd?8I:QZ).Wc</EXf4GTW40B
>QQVSYFdBDFD>9B79M,(/=#[P8Qf-L;?_0,YZTE#FBC3NS+cWLF7f)?J(VQKc7ZO
^0PUY8<)82Bb5D;^UC(Q]>P@Y87/#IE312,\QU/>,I0&,>VB=\2g1)cVa+K&UH;V
^5,0c.8:dDaEe_9O);S^UaOF,?S#a8Cd-#1fUZL-,H\R80&.31c4\:4@@T9;<L,W
-;DGKXc+Q7#Kg#FgV#=?A[\^SZ^a3c<14-MIb5WMJ=+ZUGFKM340Q5SR@WJE(AY8
>.MU.FE<-LZY/)L.SO3FbP=B.,e8+07[L3UCbWRFIN[+EW[g.?HZ1BgHXU5.D6@M
]P>aU?Pef.Jc<Pe8\5A=dTO&Y69f8:0YU/.e[.(Wd&X+ZWI.W]T(f^gD:^4gJ<W&
Z<;]/E,0AA@)ZI^GAE[B1TL#Ke3V5>)EY.=bAR>GR/SHcM\eLYLJN.-ML;,9?Sb=
cKE>(/,e-OK85R]e3B-;fL_3DQD(G.,D2(HJJX&<4d@[2/YDgW_aHLC(:E3VL;G\
5=Qf,BE,]b_T3Y4X-M7-Ng2]3:[6;EZ2dM.\1K8^3N0V0c4b.8&\:)[S;d5_#:L?
YKP2K4L/Y^^K@#V)LMK/JbN8@eU=^7P<=/9X<,<Wf&#+L1.L#G(W;WI\/>:AaKd1
=849Xf/HT_;cPTbF_Nc8O=>@]fgGU^1+KD<S,]EC6_:YA?;<Q[\7^9JI2H-]b26)
W+68Cc[BGV#@/bNLM,bH#4HWZ7ND.Pf3CHNNDeQG^-,Q0@(;0OG)<4e/e<Xb30\^
UW#:]fNQ>7U+KZM8Y1c(EAa&;K<U<,b]@WaUd\W40,,>L0LO78S5F?ACC1T-FTEZ
YBaWV04XE)fEb0dF00BBZF6Q?:F@F38#=38K1Aeb52<RY3]RI=\/T/&@I&2B\2Ec
8c:LbE4GI_H,gYGd@Ta^aT[cDL?I:#a;9960dc\P\g;,O2FPWUHG-8&8(,MAED7T
R;CKG[_2;SE6@+QYSc5MD0OG(J#aFJ@^@H0@<:ZHKa)R@[gGK:\/H67RI&M6OTHM
5c#RLZg[&Z&>5T[6X&^#Q:Y-\SJ_d0cf5aD5T\#Wg:SEFE&&24b/\.Q5GYe8bE6)
3V0AD6/)+,CgcdTMY()^aHR;LR6(NQKT]O[W5/+\E>QdW1[O3\HWU6X,GE,[IQX@
;C71B56VT)6S,\<;>K<4QgTHSHQ1XDEGN/PU;XJ3RCTg91D[N<-QF1_fX,DY7d68
95JBS=IGFP8cDUO9GcY5\7O1d(9^&HQ=dCX[HA;\;:SNX.ZcP+3)[O3d1(J\WXfL
Z(-EE<OYOP]@eaF/F#YE3\bH]V;,Z-AII\4/Oa0^>:<AX+P&-@U>W4:BcXU2L@6O
99B6[J(T+],Neb[MfRDNL>a:TFbHEW]LVLH#EM_0E>0gZ41E>+b=^7QgFU)B&2C+
DC>@Y2D#Z.dH]0,:1agD_X]=SNf?4.NKSE>>H\XRIV9;^-GWU+,#9f#[8]VQ\U+6
aY5eZ[Ie>_BQTW7DEWX(;&66^07f>Q6A]/@D]4J@;3<dA5^>ad_VYgE?We0Se#f5
EWcCZ6:TKL:E9;D(HY6M^_H[>X>@T4CONP7\<Bb_(@A_B6C;5SG>VV?5EeaafFG3
+.ge-F6KN290)#A\RZf&a#2[1D=<F/g:,dP#G1:]+M#F1922XX4c]2bJ=66Ag6)#
^QB?R5,S&^MY0QNCZUL7)],53#45XY^3b5OGG_3g3eDXY9\MaSN;?&EY\Q<eV^,d
J?FH30gB^]4I,4#M\PTVR_TYOIP.TM7+R&^(LDdIX,^3-)GfG4ga5-g;Pc9=)0M]
I:b?2(Cb,eZ3>UOa7f1(GA>_U>M5)@N&.+)g-2gc-QUAX?YEA.7.P55TIXX&FdX?
2V,:JQ[EQ(I?L>5d^_e@8]39fOW2R84,EAD<(PTV.cDZeaVE[.AQAZ?]SI5#SO0W
CL<<^A#(N1cDZ5(<;)(/\R)IZ:10S5P_3-K>C)a-/Q(G#X8dNMJf\T;T9Q,U;A#+
,e#Q=Kf6[O7G8;S+&Q:_g.5Lf4dL)=&^CAdY:=BTKSKW6eGbgXTRTJVc]d0.JZEa
-RUS^d(QOd>YG&4e(^?=J8:<#Z\.OCYQH<OW:Ag#1(=+c[g0fFP92M)_R8I5c[,7
&))96KJ54OaZAG4HR7gT7^eB@)9:Y\0?/HZ77)Q?>2D8K\2)c2THQfbFNgYbA&[Z
5)FCQH=e+d5/6O&12R0ddK@Y++>1)eESca5<T@acPC/6H;/g_#?;V(H2K/34_ZSM
K?FM]@fU(TQW-I5HNRYJfJ87I=/WH<)A8@XW=ddB,TDe3K@,J#<5c\COBZE9b^Z=
?<()7J2EJP-CV>BW#2<M\OcT=8b^40>64(-GfbP,1@^6,UVM[1VFQA7Q:fe/#9HX
R@?.e8+FKJ14?Zc@cF;.:<+QZ^8\EG8C)c>>cSAI244AA3MV.SK/33#X\B-fbLTa
,S<aC/d<Ba3JVPH+eeaWSEE)]aKV::)BgA_dERF,VZd,4C1P[/O=GaEE\9GL5WbV
Cb#^1-<65T1UIgXLg1gC?eQY1K<f<Rb+@607-^WU^TNEcR\+M<.URfaY@dI62Ja0
GYM&./CK:W;^J+J8/);9^^-f0;@;9^I];6-[Y7:5;6&W;]0-QBKD3fDB=dPHP-BC
WZVQ(>&[Q9:1[L]_a#>:EZ4:-1B-E5c##I2:63J^VTNZH>[f(KG(=6b#CTTVK4+E
8FHTW,IY(L,HB73fH_W@N6;H80>2XcV-LB93Te5EAP\WUbG27ES^UBJX>3(fJ/b_
Hb^a@,Ng+&U2CX>U\W-9K>V?^:E9EBINPS6FOE2dRTU<<6-_WC79=53KOg?b(HbB
:)eYN)BVQ2:RQ1D]/4R(-?.^-c]0>BGeg9P@EDd[+(TM@]4<^b,M,551LNKZ2AI^
@<^+ZO9cWYbC=1^gH(W[Cg_Y>UF5YZ>eOM9X:fZB6QKSO&eeL.)8YB3QNV2.W6.-
2G91R?ME9&;)^@O<C(1.1bQQ:/-c716>c?fKRg9[6,UZ/8SV6;Sc:6?U?IW1cd\>
LW,PJ.QST@DP57<IG&Y7K[M>f4_SKOQ;^7HU7WN@cS3XE+R^)J]B7Rf[946gQ;Jb
c6F14H/IU=OB(EKPSb=7[/F?01IG.:E7>Y:,.+0AE^(H]#_@f_E=A>#Q-V)7H5E_
9EKe.1>\\\-2&E-T[OZ>J>KQA6fJIGQ=eb-DUN2I.c)I&gUKgB=1bd&EIX+:@6U+
.Q3#)I5=(?&gO#>8S</\8+9M]+K7W)?/OZOKOgXG_bJd#1FKIQ-dAC^<_)^S2-Y7
2[<CRBUQ8#/aa5OM3^Y(K/7d>K;S]:14C;[WXBa@7LGWVdgb=F8MZTf5A:fONQ)f
#c5;\2b:G[72AM:f\MH(XQ:<UKf:;/?:;GC[A0K=Vg#@J35MJ=AReSd;1@1:P4=e
;LZUH7]5J5T5ee//L5_K8SXMWYB7&eN&-2FTVVU7bKQ@W.^f;2RGgBeBDRM)\(F3
UdaA</771_X#.Zc4D#6\A&^N&QY[TUWY?(A4e#1a+.JAXeeK(<QD9U-UeS[Zc3IW
55CN1FMF)V>ZWO+KL?O]dg7]UfNI1GYE+2,-T(#=e\8]RQ?dPEM?7V+O3UV8=HMC
A:4+@[N&JIJZ2Q;+Mb6XB8DF_),7XYfZ^4YY+6dDZEBJ\;HLR^,RKIN2N^_>Y2Q1
Wdc=GN>9IQ+26#:B4<=WQFeg0YK9dOFfL;c#J.;,),GXMIcK48^gKHVE@d;6D(RD
N7TZf>dKUC^/]9;-]F9,a>cEL[DdZd1)bI(LS&X;G^R)Cf-,aeY^g10RBODZE(,)
H,39KeE<_;d,.[)X5N7Eb?T9S8D>+YJ][f)MQI<gbZ[?F)(A0\)-TFdQ1P@XW-B.
IdH<OLY/f/=Y7E9R>W9QQe.06=J:15\X\Y(VAMKV59I]S[XUce6B#+;/^EM/A&bZ
P<FaRa7YW]D3ZR-ReOJ=[X7YW+(aIUgHg,F6_Oa=JL/QLY[H.e1Ue8O?F5X(/f48
C_\?Wa>#@@@:XHBZMaILMBeAHK56bRK?9Y15-.MRfU.^,:#-,J2>OGOC8bP-9PTP
SDX,#@(c9D7-V(50V^J#81]KRUF<7/WB0Uf25:=TLXf8NdgNWR(UCN84P@c>Z-.I
QJ6<#/Q,PY\&M(?N>/;0,96#9^eO8PEP,65.MT0]Db(B88;g[g>S.H1C4KJgV;Q:
<A9Gb?XWKYf2+?9PEO<P:8ceHWfK.0cg0g2?#,[3-bf\<XB]7=MV:b.M,7>#)RM@
WRM3WC4AVPRK2#5aXA>6G0eSN5dOg(b@cJPT/E>1/4IAO8WfB=Q=?4DCL[DP7-\B
;1AEd,UIdVD7X:;20=TVAdLMIT3.P(\aL.G:^33A\@a\.4F=M9+9dY:676?>7aXK
RFNgMUdFOWJ&BYY7#\+=YH;]4db.39?Cf@VMDDSTZ/BU6[?R@),V2Z^F2FP[45J<
8[10M]X:5Lf;^,WU0cSHU?]=c;4JgL;-Q+W1NYd(BHg1-_6,8_6;F-LHK):<J<Z(
aVJ]NY<J-X/a+@>.b78UP6CXVeW&b;5B2FQ:\WS4WBGCZ/C?4[[f]=P],W:W21C=
^Be0Y=Y8#TUcTW&]R#XT&2#.edd-P3N/R,[=Z&5?da?XGW8Y5U<?MTa2dd?)V(^4
03OXA.TF_\C05QQa=_:0@gedP1Fa03V6NJ&ZOYF0eGR/ZJ,<(.+HWHBQOI5aaSW=
2dLUB8Q@gLJ47e.dI,D/=8B6&MRa7W>KKWF&]&IZG4eX<K4]]786X?eN2MHP4Vf;
.a8g[S.9;FC6FX:7[871&>(^XaXE(=UU/BYg:[+.P1^F.7a<5VM1:_ggc9/7S[>@
I84M>[A&.J.-2-S@E(D7D[Y.:/Z.,dM/#11JIa:PMH.dU0-A7,2[F;UG_Z]6-b.O
8_WbN]WX7aA0/A[(f+e7b==>:U58,d+Y@>PF6c^0/IfK5]^g1_SNSaSB(UdeDI-_
MZDP)5IX3B=67_/EL>:WUDY,[:R+-VgQJYdd_XYU(@aWKAK88AgA_gMda<,F+EXF
CgP7]G[CI=4GRX4187+Q?>BD-?B7IaaPWY<7SQc_@YbIG,[MC,egR)=I]\_PX,gD
5B<=(3Y4]FNd7f=?UDFFgZ#25]4-<W^:W7aWRKNeO>a7eM+IG=PVO9@gTg8EN;L;
/J@#8=^E8M6VBaWI&fRR7IOH6gY6gd08](HI_PP@5P9Q_fH:3.XF:-[TR:80-9c1
(A0?=_]PO3O]6]T::bO;NX8T2Q#.HL9Z]#geYHIG;FMD.IHNb(WP43eRg\\7OaS_
beP0<+X.NKI+.30@>ORb3(9Q>C4WJa>Fc/IP3fA<W:Y&PR84Tg(Bc>S+;\HPO+.K
IX:W7bYU<.H]dI8@XAe/.S;d[[DfY7[5VP=:<;:69];1?gC0G=SMQ\ZZH#Z6Ta/g
-[[6RBPd\1FDA\KHY,/QT#NYK-DAS/&6L8ae?DX\=LV6R(,#O;P96K9J^+GFIR]=
fIRTX-W6Z/,@8aI;E0@F<GE0#F?+@,VI^DgcdZ<#g:5c798d2VdG.0+.VQC<TfIA
a9a/H^^^?U4SWE2EB_ZN7Q43A@X&2[75@Y&?F-IA;70\d:5-BD<>@CGAD#[32>^\
?0RgUaZPZA.IL.YaJ.93>bPWc4S,ND3^IH&JNg,@ZE:ffaKG1#YC8WEG.Ua:_\@4
VO2<F?c5EgLOK<-/I-?6+.aO;=)T;CBZ](O7>[Ka\H&?3UU<Z,\DONOD\FF^cN5R
),:U[:,/^LJLD_g,WF>QK:SNT<Q(ROHZeJZ2c.BZ7@#ad/I5+;7Nd>E[1YHcOR.V
N<dcS9)&.>L6I+&P#]g</3=[B6IYOe0A3_E#LU59SRZSAKc\O:Q.Fe6GR6JWeEP?
[Y=LW/@e(C_C.3=J@6&gb,UK65;GN:-Y1MXW<=BdL-AJ3X5SW7@N1FOb7+UD&WEC
0bg/U/P+^Kf81g(5K)=W318[_IF))F5Q/8_1,E;TeL^;EEC^]TY&MM8IHfZ8TQbd
[TGUVO05AW4f\<Q^f#g82LbD/S+R.UCWE5LH0_^M\:X9^5.<NZL)ab?])H5>(L7[
IR;c+LKCXHfHV59Wf60:@+SQbDN=KN31X\>,K<EPM.4>P-bFSgVfKC/0,NH1GZXA
g^8N64X:TCQ3/M-=J8H5C,QHM6/T>YFEY<fd;V#3<]=Q<IUTND,RW/,8]JT9W<cc
-FXL:O3SWF3Q:>T@R@BUg?e0[.[17K14dYB):]E+b9HN/ODQ,HCR_&B3)7E)/L9e
P>N4NS\>U:E+&@:3A>AJg(MJ.2(ZbRYWK(JPgCOS^1d,3TXGZf#Z;WKgb594CeG8
[2ATA2QB?X#G6\;A8,6=<_HH=eK+63?3/7V7RQ^D/7f8\_HD,=E27b=eF:f^_E,,
@V_?9J(:fX8AB\+O2;I&29C,HSCg;-O#PM[66<?^@]f:/Z15R-QM(]S3-2Z<WI^.
:R_9-\JBO5>O>WRIDMEcE)5[R91)I:/YXFL,\>,NODC_2S<?5L4S:dK[T)8BW.\+
#3<1eF^]8\CcPYWEZ]#<Od,RYE&?K/dKQ4O\]EJdfV[<ME@F=&3WBSDK?=]&@D4Q
]\C82&aP8-6:0Feg[XWeD^.63[_@B/<G12AL<H5E#EB5YW2C9F:U)WPWbK#RN6:=
/:/8e:2FR>#(ad,Xg6U^#XF7fdW/MP(+01_9L2G<>.XO+R6RWLM[3c]NdPPdHdEY
41MW50\0GGg-cP=0VYg(:>H-#+Wc25AY.:RSKEfO(;6Y<,UJJ^C;KbS3\_ZFbGbV
(Z,W6_REb\gPcd<?QSZKC,J1J4]9SY>]P>7AIH[I5WMMS.=9OB6B]Z<6R5;c4\VX
K[CePI9<KVNfeU1a9&24gKN@(85NZDUS[+g4)VbbH07A=:M&JUGgSg)gdNB:gM+<
@6LPa:3=0PW26Q&Ic2E8&N^N+F+<8OCC9BdR;)/3QXYR+0UL&[FfWdE;F=6a(Jd+
C^7&fc[NeC[<[Y^-P-9SZV<SQ/&4+#00c,^GO.\+-cD])Z6MPLI-A5WeV?N+cSTR
6Y51#2]D[X0O5Y&M26V?a&]VQ2e;c]f)e0[LdKG,1Y3=9?2RAGX?#dYP4R;<=Bf-
?J:B[PMCQc[LR:eCaa(,Be^-P7F;J1H\bZS4,0?8JNgN#Mf1,4LZ+AR0Vg_cD9.P
S8E\W0/6FJL?PcR/])JV\=56-;Rb?NcP2&<6;_I)BQa2.dW+I/W8+1&[#]X-P,K\
JVCF<KA&CT8J?LO.3L;]10OLV2<e.e(?_:U[B]QM4B.U;U&V6#([B<:3TWV2^X:L
Q,bd1F)Y3Vf.L<.b2VDMZO_f0<T\2@5-,TJITdGPX-A3acW:M8+^[/:HE5:^@)+S
M41]_F8;Td<0f6=(,e;(QK;_dC.aP\#Nc+Q&PN_6JW;F[]G0^V\EDXXD];ZSGD]P
NL1c_N3O-K#EbVA+P7Qb63T\O+O0IOAOAA_L[F91@6(KUW#9OW]UbJ+W?#W3FXD+
8a.KK-Y+WWM]aM@[e+Z77^(9=)IUc@8#IMcd2)R^,X<@DP)NaUK#<T0WF&;\ZY,>
22CcUDe<.XELF;K&#@K2#cF0F.SI0LSL1R0&Na/T^S7E<;KeNJL@S3>e?/5KcF^Y
65?60577\?FWU:@fGMgLB,/@VeN2ROdJKV:KC9Q3)bD3fO2J&VEBD^#?afe?c&<U
?&=5H09H>(NT_HcLTSH7c9RJRT5NBZM0Ug5:Q.LO(V:)T(=8W6@)TBB/Wg=d6G8;
I^3K3C;H/HHQRK-\L8DV-F<HB-LM+TM.dWHZ:>GN9QAI]>/\.+5)9-4T8LL0/=)L
:6X9;VVFP2[?Z0?YN<S2[Ua1L,_8N7/_I9N_R\DQZ&Za+N(2C5REf?@0gSRT1e4G
AJY=LA5gdC6aEY=Yf73PbBI65GPHJMV#Y5L:bIOQ;;OY<b?\5PX>1A0<=J.9URED
W##W,Z7)HK3C8F>0S]IfBg<]FgKS<6J8R@cI-M[6#g>-1MA.>bY1d<2W:=VeZ_]f
9bH:J^A]3BB6Leg9S[E>Ic5c@G)eIR@5b[&[.EY0Fd/f/TFYA+=5[0fWX#=LE+-&
75R_K):@+&@g9]2)\3.?c1>9fcZ/G#?cFGXJ.5aCKCGRBAaYWRU+_Gb3.J.8/FCZ
c:R:BZMX5K\#;O]SAa-GPK>.gV75(>f&36=KDD[7@D^+=f;>dL,@OfZAH;^^MX4E
IdL4[UIb+f_-;RZ9^FP1f#<[UVC&BIXE6-A]UNE[;HWNc]GB4A#PS>g0f5P7L3YQ
O77+=7/6U,f75Rd@A\1<06>@D)HF+OM,e+X/M00@Y8;.Vc/7(L(bE@.g>AQ^b-2L
Yd&]eV>K^RB4.V>N0PQCH[d,;LOeU=@FaCc2+/&O&Oc;:JI#cGC6e[=F4P/5VY=0
W@8&96<:OaJ1fO9+/J:\P@?b<+#I+,7+TN4?fPP4d59?^2-1&#TPU,8^MU/>3OUG
7C/QR[c,/5&A+2\fWT\_SG.SF/+?H,BG\A&&eOP@?_7[:J9-<](IR3Y(JK;Web>c
]gY.5QNTK)5O)C6C/0NgD+/P@T]>-Q11HL^_\QJ<5;Hd1N6(TGCER4_/^IL7A&0R
.?2Ve37bF58&caJ+4RS&ac@VNMbT_+Z<&:U8/4@=]X1b/^Z<GU@D3F3A;:8SN@&8
e+eE-94A7P8PX.Dd1Tgb+a;fWBM9C,PY.cJ^+ef;_U[e[;,Q2-3JOQHXECRYB\^c
;O=2XGg#7KLI):?7F#KX?PHB&a4Q.a\HN\KHgT_740UE2[,:.+(<T0a,Ab:ST.09
7(g16Fc1L1VJ:dcc0T&1@f;I,[?4N?&MX,O_8c\TcVeN<?[0.Ad(7E2<^C9IK>Ee
f-&QW&_\X@bWN.XJ\\0?MCdg#C8L=2gWI-3[3<E7.38O\)Z]=ag3]GC,H\B(_IBQ
^ON\R-CQ.-^M2;a@;Z2[O.FXU-L2a=Z<[bIT2>3=0\cJ>O6QagB+3K-K[.f\/3eZ
^C@>U[04\-3#IFP,(D9/B(T3OTb&BPW4K28[f>V/JW=SIX2gF8@?)7]80],+)_V/
JP3HBW0\dZQ3J(7d[U@FB1b2:f1YfMA2CbeeDB_SK=NQ1FF8]c:9HO_F\],HW?aE
gV(31RSO8I]VdJeBfT\A=#:.Z)@)YfN/0K2<F7-4Zgd-2(5\6G?=0/)8AE\/Y7WM
[fY@bP)C<;7+QI_,D-aE]b1QFYfA(XF]ZC[5W4L+-E70J_#acV53/L\;UZ=cZFDJ
<^WLgG>L_8.JBXA(QHEX8F;K/NObI#7g.0PAG-6YOaX?af<#<Fg=UL/Wf=(OEE&0
BGIc46+\GSBN0FV+=;+8&c5+5<\]LC0I1Y.EVT-gUd,f3^=3^cT(@fGENf-OV@_G
fX&?bY@OFC]0&K++7<&=H/[_F<5=:P,JXM_E@D)Xg7.?BE>&b\FWg=<gaG&+C+OV
7Sf5_]FP)C]EGYHA.Fb/X,71TA&cZc3M)UfM?fE8UfX+U@7cMKR)_8=a5G&N1P6@
2J64>FE/X>;Ye0WY+D0\<Z7^^(8C-QcWI\X2c/(F/UNLR#CVB_XAF-0+_W<d(E,X
=Z5#=6-.KO&(HYe()5Q9]^1bCF.ONTLe[8>UG\V)DE9Bf@d;fBUPbVfa-G6a4cbN
,ddA6X36cRPX1=d>5A-CMQWVSFH.ET,&2+PcdU0J,2OHO54-2JM29Ncd.@W2CAJb
RDHWGC861]TP_CAa;UL:c:JW5)27X:&1,[YOT34B_B=Zd5bT;f1DKbH(S[YK[;_^
=a=6Q2V54?c<I3cAUd\<GfN-D7_Lge]PZg2,=Y[28bGQ[(D_?gdHFc&b3E[41VMW
--^1M9U:R0Jd0(=R>W8c9#2c_8\YQa9</BHE@7_56dHg-RQN&cOd#8#dSUXMcd^X
Fc6XX\R6IGN(U5feIf]0Y,-_E14g28Hg56N7:M/H-@]EV89Td<Z4IT543B-\./W5
NeaZ6f7V4V8T@^/T+aK7Z3#DLOB+bEV-LXSc=;K],<cW3E>MVV0M#.)[H+9EHSMN
MUAg+bZ36SO4V0VZ?L#eMYF#gKB.Bd-]9e8YB(eFD:gG=De-P.^O:8-[.HafO#>X
dNd9TIPg<23YWQba8D<gHf51..g&Y6:OX01_]4WfBD,6G\^;&S;8MZa<K.eg5&P>
?:-NOFB4)_JJ6LQ0(1a.aS1ZU0\dK-^C[?^E7L]6g2SU;<E2KIWLM9LHE[LT8?Lf
^7/.TF7>PJF9/INJ9PCe6+N030@Y4=?/McW,_FB,2>aFJBX^+T&6&MSTT]LR7f]X
eZ_;M.,@/RL?V3S8>B/8^=-A87b,d]F9A:WE/4RFZ:GIZM/3.K,QI(Ide-[W\ecZ
,Z)2&dG+MOgGBVR=ICX\9LJe6Tb6KNVRUD^-2AL_FI=/2/Q?[F6^5FEKAEK8AC@?
F[1^#.fL[TO;T_N[6_;J<>6cZeIDSc_.+BPE\f:#(/DAPSOSYSK6c+cW:[aP>X@=
N)LALW[OcgIf^:8;=HJ&9QQZSJ9a5].JQH;589BTdB<U8&F]WSd.]X#DT^bTgf_.
Y[TPKM]-J&D6E\V1D[IHeIR_K:H:Y#RV#6.^A0NIK_SWa=8a(E_::4_3(D2cVg@O
c&.LKJJ-+N&AA3eWJGOF&-=3ae^g^+G\1bQB?RT;>;#g-A<66H#,DDeeQ0ML3G<_
D17ae+AY+eBAH^._3&R1D@168)&BM+1g0FXHRN)695@JP;&SI#-43-W1cc0M>8FV
J-,6g\[LFf&E@R&4fc^529/U<PL)bee=[G&ePDZM(adfE5ea\LR4b_7/e8cDIUX0
4Tcg6:&ZUTQ/;ZQQ:Y5[[6gg5NEd3Mg45K>gBPbL;SV7.WQcJ&-f>O4U@&B:E,KX
Cae3A0K+bJHX3XE-C^7;HHR0B4P(E#=TX7BaR6?WL/6e.;9D(G<gKL[a9ISK>]FX
#^0+R9UT=9)F9XP(_^(W]=f3a.^Y^5/5PN)H3>f<:9UE7E=S9gEf^JNf>EG;+S2>
XL28,T)6A@=22e8Q2g+Z+_&,e8aa+0X]U0)Pa0ALXPZ/A(DQ[CWGG:]d0bOR:JME
&-&VD0b9W^94==AY>-7Dcg:W^@C0X_fJS5>3HV;)D7M5(RG701a:a@F.R(S_=7J,
;:H;7[(7\POE3b/NR[=KU5\ZY>KW#?-7c0U7^^9-J-&[LC(AdVJB^VH:-<IF@f2K
[2Sde^0H@&(H]X)A3R.aZOMSCKaB3[7f7Kg,_WAcZ#?[7^5D=a\8g7+TA4VAD53T
#f=.A+,[NQQJPRA8>f1Z;9AK_I8aNL+7HCRWZ_C56I#CWF455Bb#JOQef<T0Ne]2
IX/?<b.e,N&KE(K<Zg\KXUI((E,GF<Z4>E0M43^BHAP.2;@7Gad[FGGJL&_0bcZ?
VaPQ7A>N6&CcE33QB2F7<Z-f)a[^7.NG\;OV]G^M@N8J>OGZD;XAH353QY<JHCd4
>1^ZG?77/3A943]:1=J\QUdR4T\WF#OS-a[0Z\>P.T.a@3[<5Jf]GdQNfSY8+1a?
eN7F8(<B;T?JI\Qc^JV,;/DTbEI<@2Ye.a3]Yd2P/Q]@2eNK\#(BHO.##@]2#1Fd
Y7X7XC77a1HJe5c+eW^C\-.0^gL_UQ2D@WQbW[</OT4_WPJG^Gb-f-RGO2@J&\@8
2aY5:.f0J?7U<H[@I>(:#dPHCZ8N(AS(ee79+>2CWVI).)BX7V.eE@c10_8M<@-P
&dU+2O1SHT]acNI_P]cH.54dJ[1X^]CEY)cKAZXSQF#C45,#=#4ff[XO-W<.D)A\
PZbFaA-<?\??3JLQb_?8E?_^@[(a5A+/;R.SRMfIHgdTU)??gLe2?:P&6H#712\?
]14;.NMS-Vf/dB9c-DK:40[Lg68VRI:A].LD>c12-7YL\[HK)K8Qcac]0A)HLd9V
;aPT[E?a(_#Y4);L(9eZFJB2?^Nc(;:OX<8FC/]1cDfB</K@:)()S.<5J)OG.b>)
a+1D\6_5:B9WZf,M[&T]^d.5HW;GLcaFg:B>6,N8,3WNKC[M9X^V>.;[fEZ2G?@9
Ia5G#g35E>T9@6=,BQQe]^.103I?3]g/fdOe5O7c0-VI,>0SFVMZ,F:#KD5#G_Da
Z=g&+^HFNeZ1?[>-fP.0F_^HK:b[XVa]9#9:LPSeR:D8I3.c46THe:A]G849=Y2R
Ye<,QM9GQ1///C_]I3S=3/_\I.2#V5-RX15.C4YBe9#8^R+6;P._?)N2+55>)&Q\
B97T20P_dMBV^.\V0/JDRQNO9cOdEE->>QI&G:GB/++F:a:72WCOgK7#3UKHV7VB
MK<++8?^48P2#EE.Y6d8#_J41UW9&=JSf[g1;Mc3.9a;[Y:<e=O3YZ8ObCNG8K?;
;_\gd<TJ;N<H:>_8^UL^EM;XRb#cb0SVHW<;SXbGBU?0MQK^#-VYAT+0?TFO(TIE
FN;6DUPIX1IRDTQ0Pa&RWOP0VCB6E(LOR#Z6-;4:[)_Y0))N+4O(;f-/(A0Q&RgN
4OEdY:42J_:E7Wc@5FVPVc)1/V0-FQa;Z8ZDQXg\44,G;@1dPZC]W,(9WND7B&VG
OIFIV.D)]a=<Z35GYOfCPNLE6BY5=[?L<\SK\8K&L\+5QZE+LO;=)].^?C.Y,Mf-
d#=cK#GY;](@cE91HADa>_L=8)-ZNP+HK&XfJ<_1^H46ab]_:QL:^8K)@=V>f<4Y
JLV-d66=>P^TGO86=322=-JE6Ucb5cC#SEA[22Z,K#YcUKP#[)aGL3Q(HbMBI:&e
0.U2XNcJ6(3KH=SaON&&EL]ec[>L?c]6E>?^#DD1OYM5,JbIe.:XKK+6Y_G#.;;1
:^9f3&0f?/_gf,<gF^+[[G1-3<YZ&KJ-R5+T5]YGJGL\Tg(5@14G<Ta>b_(V?aee
4PNHafQ.37,?YL^K3<dbQ->2??.C=BVdV>C3@[?[U[:7.>dNb/0#L>cdaYFZLEGU
[]=K\4c:1bX)E1feFOSfB/bbR>;8:PaI?Y.9+1cM9PcK3MZ3:ZZX86<Ac@I7HXH>
]?gW&bW6;X6RL[W-_;M(YGQ<F/:\R?X<.2I,]1e?5ca.V.PHSc<O+7C=&bHT7=4a
8Y^R>8M@?SL#&\Le^^C7JHHRGHcOATU5N747&V+YJWbf^]:gUBJE;-H.:;81F-=M
8ZE]Ec,e\.[[S2EcFN9=IS<a+EH[K?P6.^LSg?I,/8C<af1/RD)a7_e5.7TO,O@A
5;d+&6?V(FFJ5?F<MH-SW-RfCM55<38#=&7;[@HgLL;:F/7-\F-PfT\0ZA_WTK^@
K@BLRY[B&RYT-#<ETJd05bg&^.&OR^CKCA\(eMOYQNAROA;J[1W<1JCE44=>D&1Q
KZ+=g2BO4K4&S[7^VRRA4(TKQF/HUFCUAXTS;^I17IdH\A/CbNOL:D_/_[4<ee+V
S5V7Y#N+6FfV)71^LgKGR]<BMeY6_+aTM7[[&0^OW<[7[6EASdaKEQBRG>?2V)KJ
Q/_FdFe8_K.NL0/J<@X]^-DU+0/-.;_W#@Sb<,NN>F@<XO9<EEXQ);<Fd^5.Sd;b
RCNPIGTN9A<0CM]5G:O&PBgbX=-EDY1):XU]T5\Kg(<NE,A+AX.0:aM-B61&4fXQ
ZM72K>aM6<Y@&VD20H]F?9X_A1WM@24XM@P;gfF,ScNe,SD3aO<.YRFT66AVAUJ\
E:f3P#VR83G-UB2DD2).2AP5OR]b8X1J+EG+4M[Z8THG#cda_HP9LQ/Q\]f7<(gg
_[968D^FRbKfWL721a1&;K&?+@]#a=a^dHg<2EYTKY3a>.#(N.^fAb8AP#X]WF:&
7V@_<e(\A:eU;9154^26C)46W?V5Tc/aPJ&TJY-24WT8BF,Mfd<@14@0YRRKNBZU
OKT,FaDO4BKX96/9J810#<^-VM[_=T@^2:L&D@9/WWJTNeU8+4-fF&Z=DceGeLR/
<(#D>_ZFU-Y9D?GHe8TW[f#_(EGKFR\Ode_/H5D_72b(0PN+?]g8XWRDgUOYBQY]
gCT6-IC:c.+_f--[MG[9A?L9#Q2Tc[J3<58#)N+Z.A.Cc.g,-/2:.Ob)VSKYa[DY
g-X#<=127_8VPBN10V<O[La\2_19LD.d45?2AQ_Z5[a0fC1]cD_#-MC<JWC(UDQ8
GYC,GLeV-W]B(EHX4:eZ[_C-P/ZK.KEV]7Hb>;LfO?V<YeBO5R>P_L1)aH2Jc]M+
&>6,6EbEc+M.0g7B?LX6P<e#Ge7=/\G=(H_[N@=OYaK9?6dN49RBd8.=1-B_Ta<A
\Xcd6/0:>GgBc2\W&,OX]FU3)CPNE)d,Q)c\eB7E54U9@PV.()XJ@<V,#XI.KY)^
M5.<VCYD(5Vc7@[Z,FFAbZf:-QR\HcBR=:aTHX-:]K#718eKT]RFfD/#EWZP](Ae
FcG@UT<LK5QW/FRXSdDEG+d4U&RdeS02C&(C(X9@LU/6fY?YeMH]?T>K=I1[M/11
6CDU3RTe4^>TEN0ECXd?UOC>]<a]KFVcO=bG7;T@O#[e&M6:>)>BWg&<a2ZM0RY>
3CK54a6bP^FQ;>dR^\/W2RJAHS@6S]QE+cZM<)MI<1(:\7JD7e>W_a;[.1(_A]F>
9d7W/&A#I]ed(XG/QJC^B)SK08\Jb@.5FdKS)X=MR<e226E1]aOf8]6b\Q-#I08A
H@?VD5[e_=R&@gK@Z-=5&O5Mb(]dfBLBHUN5OC;N(TM_Z\c>b:SMfDPP]6+)/V\2
(66XTQFE:L5+gaI#5I]DDc?4#TE+[+:WU99@9#c7FHPXZC1_,,Z?);9H^1MI,_eA
fH[],<<ePR@DZ\+Ia+;?:Z7&\AP[#C/,Z91[Dc5JR_C>VE0W655@Y>S5Q522EJTf
V^9P5=UdA]d2R\=ESRYLO2V7JI/4Y2,WW3EXJPF9,U^1/bUIZ[<YIP70=54WC6S2
A<Z>PP1_SaRg0JQE)/>+TST^O,@)PT:KBBAL@5<V5^A,dbc_TGaed0W?cXQX>,:\
AdKO;g.d@\6_0^-P^fR3<SA?[9P247S8RP0M?3WOLSE1K=ga31c)SDJ:;\F6+A(5
^aV8=X]T&74M\]bbB^4\ME\D=&58UV;:3g/.?7,ZBIGM1]eHY3[GOF7#M^:8/=Y,
eNJcW8I-[Nd)fTO@X\Nd8L)8RZ:(ebge1f]b7#J(+)C,W[Z;/W(G=J7=MK_+@T/g
PWW3KNd&#_IJYJVYW_+R;JI3f\Q<N1)B.=,cOG6C,^M?(V+6M-<PbXF=)XHe)U9M
C^(M_,E^Fa^P0_+GAR36aJ20-,aH]?Xa4Y^aAS<K?_Q-87a?_&>Dg[Se30UCc6Eb
SMJ<2cA7^>A]\RD:b68@10-890<^bZ73#Ie8@TS:F+-1K\f..5LB_2\_11]HSHaC
J-WUHUZTK[G1;APEZB?,7;_CT//N9=8/aGLP2@:PJ1?g:L-CK@NKIG/;;_)_J(>0
(X>ZN8KT>8CBC:/94a>7Q;CbMFOd+ZBZ_fe=[8,7CF)8F=3dZ]VY7b2NR<L7Wgb\
gG^=I&U9XW9(/&@W&agdZfRZ#&YaF9NVSYb4^>:0>C@1[^U:-B0XO]F2YGDKKJfc
=?DA>a#HA^6[.BfF?D,^c[7_,4.f#W)FEC90O6a97V,eW]_CcY]WES.V.C:49c=Z
>EBXc;R&6,N]c>T:ZAZ+gU>K82W,]N8]Jc81;6eBbSRWGL6\PII+(DJc=S6+^18?
G<XM^J0.S0CEW-N+K^E1&+(QHeJ\(6W:JEVG^TF+#O32?5:@8a&5_SXg.EeX.34-
^:T_CZ]W(&3JCWd#HD&IPfD=Vd_S6eXGQ-#<DfeTaH2FBMWfO\TH+W20@VL_V97^
NQ5DcWWb.7X=?G64QVQO7LSGf58;)0X/2B=f<M^]^a7gW8H?a66O3#eR(N[X(6&6
0[9RLa5)V]8^U9GU[EBKI6UE+<\,=)A?EcOSb=H1NaC-3XDQAB0@8R1YL(0c_]/C
2NU[HFYc0+YS#<TaEOVNdHEEZU+=ALID:#c]\4SBW0(Pd1?Oe[D5eOW2AcaKF8Lg
2XLJ_XW,9QT=#0HSBX7G0-5,VMK^EV&F(_M/N#JS^6A[bNP=)W,6KcOS^OBA2TD)
?HA6FU<&K/EWOHE=CH<Ve//1.ON:6Q[QT>F?)QYdH]GMH(^(2;5)?B7+M,MU21VG
K+>)gCd&QAJ_R3SZL)#d@BPJAe1AD6^K7H-CCRR6TJ[^H>8?);B.O]2UPBSd0;5g
06Qb9KZGG_G,U8V/1=P#QJ69O&U_T0_IN0ZKU/TK=FHY,PUX5RVB\b2O2++@g<c1
9V@[4U&3-Mg16HCZd31>:IY;fG#3]/dM=(DEVS26T,<CS[:21LTQA+5W4c.B#4a,
cfJg:IR.7C\I0?NY97L6SI=;7Qea&7fdc]^]JZ=;M<\5]>_GKYK&I7#&?V.P2eGW
EP#7A^Bg9N&LDM8,af+F@,SQ1Z5TTJE:N:a0S8:T+MbHI6If@WVf77O2B#?\b@?;
f2^>b/38;QaW/0aJ]1EW;Ng4T(CaYWDKS7ZHN2@W_,7UV0(O?EZg[_Md[F^FF&N8
9EVAO@M^0<DWcYYG-3#J99=B8Z9T/)]R3&/dBda@5PA7S,I;R]E)5aK<&N0+DY7>
\f:1JSTE3a^/CUU16A1f\VN,9=KS.HKVLaX3.K]J<PP2DO;D&3^5aFN[aO8WQfY1
5&+CGdd0_(4O[_U]O0EN;Tg3g?5b64eLJWQd2(5<E\?[aZfVOb>9HTe[L.((DN^/
SLF@b=L<d0YB0VdO/J#F<8f#b_UIe1WQ]We)BbM;a^e9Y6Qe_DO/X.#G@LHH;acc
,H.,+##E46-:5A(UY\.g&0X(@B+LKM:KVR_UgMIb5:RVWD?4^L,50[SE8QPF-Z&)
\,IOTAg3RB,F]Z3>UG(#gF+8JT==8;:\Jea0936LBHEfaF]GeL0EI27U<Ja?6></
0^;S8>:I]ZDWLP,3&M\YMa6>S&=4]b;.)cg@B&5LO)@LWR<]9CM2c,NN5d34O<X=
G:^J2ege(?#R4IYKf^#L@Bg/84.2W?<Z>8P.56A@F6JOef;c#ER/S;S])<BTg(dW
+\+WPN@:7/9g.MVO30IA>_]5.LS85Y?g@J0Md5ddB,)-NLcPA)6?1D<2==::FO+G
gH,E)?+\(J8^WJ[-=TUH@?TZA1Dd6>5S(eH0VdP87#0@aWffZF_Xa=IQP-&OVdbA
(YA@4(#[(UV;=:d)8.)3>QHRdD,6CYN2@W_:Nb2LJ6F<2ZKa1247G00BONI\B6G.
F2Ia)((CgZ6\=OU:gRD<MH<KYC2WIgS^NaZ3J3CS818_G7M?QKUe8d_,:gHFI5,X
SR2Z_=K_>:bI>T_bK_T+8D\4)?,H8PH+#,ab,<Y?Tb_[AUKRdX;9I;-df,27JaBL
HD2G]eY<2)(g0(K=g/_<3.X0efCS,7MWb^FM<@&EfA,O+M(I-aO/d/e2AOB/\8P^
M[7,B3A_b8]WAPQ8bWF2/(=b-XL&5=W>:Qfda=Q/XBS>5_7OEG_9Z4=Y0<X=@/ad
F_YWK);8?0DJF>IaXT[ZQX?<64>_?ERB2,9E2#?GDcFcU7,J6d:EVC#&6>C2@IHM
[LU1&I-gLegL@UP1U6?8+\QS]b?c?S:Nd=d4\?N1PJUbASdQ1;7_?:O&UU.TNA(,
\2955+?,GZN-1++bgQ3<cRH^.e?HEM1-JCA(g+;O(G_^3+ML9&#.BE.b:203[-AA
?789R&TF_U8QG<^UJUKSY?]K@5[Rf..J<HP+40LLK;QI?EY85OO[J]U6#)C=&56b
()8MA&9WfW5J??W:R8.eQV&LcLHSVR.UT,a5H4NPM]FW-NV?JX,6fXK<_b3@9G#H
bD[/0L907GY<QRb1P,1^P.^f>>]&.4N1UX<Y:NaJ?LgM[#IT-^_3_-6U41GA8QX+
8L]D9<3X6&ec2dS9YM#\&/3NAH<;d?HZ-M=EJdd9\7T[?2.MEGVag2^BYD=?0^]Z
g1T3SO_+8FgMRH@aH]?f[eADNLO3XZ@SQ9e5#0>KRSR,0Z+ZECR4,c<0=f&PRC..
VgR[]d5W3-XE@G4+OXX8K()Y1fgKe\13S8VS]__T&B0FB284M2)=>HXKQRQ9Z-c-
C0056b5UZ7dP6=gdW7PMK]d@RPK_-0+_fN.c;Dc:3f<?7:+_S,KR5JYCTW>.WM)A
)706Z\]UJ3;66IXa#XN:#KdSR6X(+K/FeWHE_)Ta,NTc(3B;>?Z1L&E?Z)XHM<<K
:(/;ZK1HI560WG.T;4c.&STDa^Of=+B=)6?0e;WDY[gUR=[8^)_9//?L2PHCG,CO
K4GIWP_O5(R9YgC9(SYQ3E_)gF+?a/7&MM-P1?GR?&9H=6Z_^UY<L//0CVeSS&>L
gADcJN,J_LUBOAM[&I&cXX1DIN\AGG0(7TgQ><-AdWbaJLP8^MGe>>c4e4c=AED=
CQb?^[AGDR/P5BE94I5.BT2V;\C.7f-FF?^I^.O;8@OgEb\_S37L]O#gRSWIOHM@
AQ=?6D5F[++\6C^>+;/4:]cO=9d./7S\<2,@VE-fM1]6MXBGDf.cT_d:45]A-<_9
V/UOW,Ld@W\W&Na/?gJ8OD,I:^=EC#8:S,+#[N\fDF>K0VfeQ\@<ZgC=8d;+<FH]
K+,Q(K#;(0AUNQTUIP&d#)QI;-ND=6WJ[B-BC;M@=B]E#dZF[T.Q1<5587g/KNa3
KVQfP#?)D]O3^IY#B12.c2B#)N)89-K4D[c4A=bOOg_4OW]2E_Ad/78:)S;5@&=R
\bMI.[Uf-C/9L_-f8&>G6OFaYO;Jb.>P8Y.10V7=6d9]-Yc\?XI5XZI4X?/+E+[d
aAU)f0]1A^0RN6P=HM#>(E+:OHR;H/cK1acKC21&Od4,#/UJ&/7U(]fAD75=,?YH
(NP)E9c>KA_[HXXA5=PB7fA2b)-W4YJVI8(QU80Z+gFTLS-9]021G7QP>6,ZQ^I:
eB.V/ZKP40Y-ZC?T[f8/YR2ZC22NGEP\b;>_6.^Y#e,0:c5#QOXP0(&2AXF-Z+?H
YN_Z&ECe/0DM<.X5CVLF))YDge[XJX_2C^LCDF)41\XD)2eCQfMN7D&2d06F@^IB
@I8?&fK=?,#6c>W?N8&G>KB80f:OKd6U_1-13KY5E\T.+54O7KIR6>U/9]^2O;Pe
b5_R=^gIg.KX@G?BU@\(19X7IZ[\eWRF\6>^=7f/=\4Y_(_.WU&+XN&6=UC,BdWd
,,5@#\XZ)KbD3K9W))<g@@^1S),[/@+_UQc]RO(/,V6,]eNZ4W+-50d,<\<N./W#
.X;7I:)cB@[3]6+^&f?,(4FRR)WPLQV_L7SQ#^>MC7^:6PV#D;ARgdQ>7;,FXJOS
LA<W^=(E-54DX8SRWFNVc?AMMYMZ@U#,g8e03Ec3<=e3UU,B:^TedDR76f+3^CKB
(5A.gcF&0aOPgAf60D09BdURHKg,;>4-8/9>2&Y)JTNEJU\c9FTA=KM>U2ST&4f3
T6)a0=ZbR_BK-[Ua_B(c+L23;G?XZ\LT62+MUX3JMKQcMN^+#df934SOfV2b0A>5
G^<VNB&OT@f)ENMY2NF+;I0_1Yeg+CNEP=cHXI:TD[a:I]C92J60&WI<3a0[,V@9
1]6ge1Q>/f8f:7Rg7NZ^Ke4>TT6^dT8V[0D21-:+]9Uc(AM&FQ7UYO;NV-]_db6C
,3d1VZ[M^;>]bO+LUD?71=Y^3@4FVY<=f)(KY@5)=f#^-g]XT+\ZEHV4D3H,e^T,
CO<G<T&_205U:/;E,gTG5;>1H9;WCV=^e2MPZc)#I7&^D9/_>RcD+OIJ]2D)#>-;
4]);@bU_3JGP@B1BI8\N@]YDFMR70Q[<JM\2#EA?deJLJRE>aY@&TG^2f[8PB33K
5H++<P8)7/^d>)[fO4#P0b@)cK=BF-ZZKW\4R/4#F32A>7YTCB6U?9ff-,_TK49+
?^?8NbW0BOJ4C^0ZT+FE]NHd=Z&BI_B_d9I_J5[Gg:b,CYP#Z7S<W#JV=Y+3;WG6
&a2,U2HG[IT0_<]#?9,)[O3M0.YDBIQ]JK9;bc^A&4TBdO49f+JZL[Sf9/+9<dcb
19,D;/b,L/F2L=4;fQO6>>EVXP0.@PJ7Z(HN/8Jfa:\BHW>Sa+TB;.E2OZDKb6]T
VE\VXT&/VGFI>RR/=eOcMO?:9RYO+<0&JKf<P73X#_&231UQKd@6O,BZA1K,.<bW
>-caOYa3C(#/S)?D0.JQCT+T#I1NZI5I]]0aNN8Y[23X9_<.6K=)[-4P7U8dac)e
<a=>N^W15H_c;<W4^Rd8T8+LG.BS5dFJ.+:b)<[OG0eQ?bWP09H(70JZ6D5]O7Q@
4W;M[3bJZ[:UaYD(5B[CI-Q@I@1;K;/TOD=7[>fYb^b^8ZBUIFCV=&FPZN5b52O1
+F+E2Rb3^6ed&NbEdKM5Jf:E4[B\e8MQ^1UM#UaeL;JK9NDf)B#(#TQZG7gP;NO1
0^I\eJG7);5IP6R3fGV?g88JI9cR?QJFF)A@H.C#01AIeEZNNAY73<gO:7LZA&Z[
CB;801Q4/2F9ZHF7>A1Q;31N2C,Eef=UAFN[&X@g)DMPcQ9eF\[0NWgBSFP)^H5g
0EQD@WO=.Tb:;T[RXVFCIQHYVZZ)&QQ@MOD;S-UY3fMFX\/)FX_TO,?Fea>3IgTc
?5PEPa=+HIK\dG\<&9(0?LI^0/^\b39W,e4?9@(A?bFa#,=/d#7747QcA_>Y27HF
CaJ\1A@1(K?:bg11@KHKV=@f/P4W,[#<VH=O4TCJW#^cN]2(W#(L7;NMQG949A#a
[,#DPFK-#GF:8,:>J2>VY&Bc6L=PEFJ97KIT5AN8gXYEL;B,WQMT3cb_>cc=@d#G
88#fgI1ZIQ=]@;cMIT_91-M_F_KG0G61>6BAVYYI5d9Xb^[(T_/S.Q1D#5[_K=Lb
bS0-+D0IcK04JHHDGM5IIIW_(:aP41EL#_1;Z+&78+A]B5KR)SFN&3&2<=7c:T@T
bfg,_N^W(_M2S+LCL1PIJegCbSD0\PZ3N]T4(1M>NMF?VVM?\dE)6_1&/KEBD\-V
95Jd&@NFd2/?CP.K9G)&VR+TJZe+_&8+Q0g_ZQaO.J@5Pc<T#3J@XdB-Zg>LP>WF
W,97:&H1/3\\KffdW.[98#57)<[.^cXGPV-E.;#9beNKJ&/E0JH0K.dVAbW+fB2f
d&X1I6@<=KaBD_0@Ob7MJ3Y:@2fQ^+:/Ad96AY[?(B+cKeQ-:KNc^/OP<RYgX5:f
U1S:QbBM;U0eWXY2<bW.F82CdF1]KOFOA9I]+dK_D<GM&0H1LB>AL>b6]c[VS.+^
d++MR2aH^]Q-R?AB1VSfaG3QL5_E]4P_,&XCN+EO6&?0BU+=MS6MNVdcMG<(7I3-
e[ZCS@SA#^4K)5#Q0</#DKWA]1A]2eI(9CaG-Af_f]TL^c^>BD+N[2gVCa@2G0,;
0H,)ZXT4Yc7^&EefMEd)129?V4-2c(YPMg4#ID#0VP1Z2P3IKc@VYg0H33N)V,4A
/a=^C>d.(YCO6W(7W\4g5e4?;&[Y-1<K2/()ZQJ6<9He77E@]M--5F-S3)]3SYLF
]+^^)25/I4I+#,:bKQ)&[IaCR)TgTGa\1U6Q[]M^QP5/:11.LPP+F^dgd];@0[6S
MCZWf.1ec+6./AafAFI-gS(QCJa)+D1PcTV=R3H=B+gLP^)>e6]0;\PgXOXJ\d94
?_CY>(\@4e2eWSKH+#:IG08E+6&NNV]]OSZ]B7K\?HWf<=93ZW,M#8@Ie2@+OPe8
Xc^WTL<2>[Z=2@QY/55ac5WW_Y#[I[T=09HZD)@IE[;4HR(e^LcZc8b0dMXJe&IP
2)]LMK(AM>V4_;5-E>_AQF.?P<?>H[:<>f5X:A9_MIUIf9a?S9N7><]F2Y#,6a&N
^[9W;;5dP)EYLXHZ#)]0_Ec14],06;7^WTV()#c@3),<ZFV8YOU4dQ?[+,.G^KEN
I&f7P@/2Mg_LZIH]4YDC>ISLVZ:8,UV/L/2L1U<Z]bF8+>V&E-b.:0E_?<B#P-Gg
;D9RSS]>aIYLEK0cQ_d?1V@<<5?^E-JTX7aHJV@Eb3dHPZ&_OGYU9MWc?TTFAT61
K_XHCNTI&dg,7&3MB,;GJWLQ8/(F>;f:^T+gc7M1VcA\?Z##9Hab+.2+<N4a>XV8
?],VWRU9_)90)?1-8E8C&&][]^2.5ceA.AZBD,=Nf;JA/,T\JJOa^TX58aS74GWG
6<U5=?b:@Z0?HH3/V]fcNLbD#4FUPV<NC0<72B9OLP(EFRW]UW1d0&;F-/DfOI-^
Ub/[X6bU?+<D43c;=0:]K-fYC3;LfBCPeI6D1d98aWA\GQ(eKYEOU---UD>8]R4H
3CcA+^>X(])ObOHW4+<V3(KN1.JdO?Y+-^V07\[fV6A?2@=&1cDf-0](W\f,cAEW
gDLE:&U:A+P[6aMI0d-8;d1+,1HcZ(/^fFEU#J:&]cB-6JTa&3TCM=bc7#[bBXX^
d#015a=He(bP.JfcK()Bg;]5;.a;CWa4OL.ec,Q[Af9./?5Rbb#XVg>Z@R14[DEI
DYcU58Z<,g\[+)7_+G5LR>,c-d_ZG;G@DaDBfV<P+AO=X9#R=,7VPc1-gU:_VYV)
;,NX77@TBZ:OVMg6\gd[9Y?1=L)eMd-K/gCF/MgJ-K+I+BDX1G3UdM:O(V8&3GE>
(T1eIbL^^X[#+3C\&\RV,OV.P3NAd;eX>\Jf:[,P=40KMEb:I4bLTA(Yb><3a&).
(fU+#Y+OaZ.bD.1<L.@>AAc=eZIf(_7?;POf3&D(eS5AWaU19?K^d&0g6J1ZLB#R
1>^e6X1Af-@e1;ZP;cKZ&P(BMe8V[DHOe)J:I7K5)<#KB+2BZL#cZ\B=c[8+DJ]-
TEIWCO9URa3?3:22bG6a6<eeX@0bQZ6LJ,7MJb]V2F[98_:1[JC^^LAS.I[e-Q&X
W/Bg-W&>(B\1=LIc)D&eDR:V3)1USQN(XVL@@W?Q]SXK4gVH+FR]-6VH08PfT.7d
T4F:/_PR@.4T/M?=CKN#38IFI5+LEI\Y?FRV+T=I8c=afCZKG>dB_@6_-J9PO6BG
9(C_M#BH/I8fE<,<MgTKfVZIFYE]QF(-&JATb6Z+=Y-)M:8P@[;OGK(.5D9#Ga8=
4K8VSQ.M6Dc/<]9+RgLO,b^QH.ZMb.KK[^]<FXYK1A\UBeC(BX2IVfWbYMPJ^.Z:
Fc]RJ^6U@3)e67=K[B=-Pc),H\&WQ]5/5)XZZ@fBQYZ;XE;3Q431[5D&2(#3@>CD
7RL[@TUGbITLd5CEEQON&de0DA]TH86WHH=Nf41@QQIA8D-6a[1?;(/<UET8Bc_b
@0<fT/Q+I,a9bG2N.>EGV\YU+f(,e/FVLL#7X.&P;MAE5TWIVZ12]X^3Cd[C)1WW
;=W(7;/G<UK5C=^K09FHI?gTQ30d56^cJTP7/3fLBIWT_O69b6?PJAYU@DO5O+>J
A5@@[[FYQN&ISeE(F<L35<b/FQ<d-,G@2A:2\?[W&YOYH\?F=0STFUSE)-8H@2d#
_4\79,XSE6D+aH@f&Z46>-<3<Wb.9I>MFb(8INL7.a-IRM:,USY-?9C7d;VUCC&Q
A<<C)bcV+ZT@HUL9/aKUJf.WBC2[-K_B=cIe+7I_(GVN#bE/4+6KFV.@7KO44Yc-
ADY(2IWe\(B#)cA8E<..>3eYcgRE=_T:J-.08C<>A#8XYWcLAgDe:F2QDOIbcF,K
-E:SNPSA8FZ/=:F=CBMHC7-@__FR^2ee2HG<H?Md83WKK?.#T3f<1f[W7BS>b(AI
?C9=39>ML:^\B6IE68^XJeV^Yd..))I[W4Aa?B\<RJ?-8+2ZP?KbD]?9^??7=TY^
a2?dN0KN1@=N9SC^Q6e09?@dVOGRKII(d8VI-Jf9e84:)@5EPWSQ4A9EW:>0FB_9
@6WJb0TZSDJ_&Ua^ffXdE4IEFc3Y#A3Wg/NBTUM65^PH<22M<P.1\^d1b#0\Z.&3
5C3ObL??VV@2Aa4H0>2+;8\=K(,@HQE;APX]caEPfQ;=C2C#_SfV>ZgB#cIE@TH)
Yd>R5Z6AXdWP8?e/F^3\EaOD=gGU2a1)0KVcC-)C\\9D[2MFa[(_;61eU9I(be7[
..R1.HN=cVX.H:0/I.b6D5HH4Tg02Qa?0_[I/_JfbX3SPU=8B(MAWb)b1eZRRH=4
W5X3OR,\TfW-T.b5cYc,:fgL;+aC.=:X<Cb0UAa4dT;SVT=Z@/VAYQf2NE3I,&PG
&A[\)C?Y<A+Z?Y<T^gC12eW1F,:ZeY5=B7D9g>N,^265=G04g0c1F##8;+K@1I5e
(J5L2f=[?H;eY&SM;R(OCBe[(NEI.F>JEHLb9=fZ&DZR5-/#A/6)F0>:aX\CZU22
dg(KKX4?OP6S_OM2QYfP.2<Na0.[Ng?,aG<BK2FSYXP/CfJX&E>BYVZ5GE:.(G<)
]a_5T[,PEXV@\8dT]?^ffLE(YL5a]>)I_DH[U.YR.TQV.RI9F</1_(c_+&>CAA]8
?6=XFYcU(J:N4G.e@E.A=EC+JT0/AXP=18MP74/gC_dT8,32K7W(#4<[,b5aE>64
b52DNK_+SD,I,>J2@C.dd=T\;,K]#1R[4&G#+dJK\d9b3T1J88+JC4@A0?A)M.H4
Z_WbK0..ATYdGZHa-0b,;Lc#+Kgbf#D.(O6+BfG?DNY^=-Y:#,[^71:X[afN(Dd(
JB^#SHNY;#bVIE2XH]29Q2BU-[@FZX<a+S.P@XQXcS<Yc09ECc/+)O>BWQM6S)68
SY=>VLO<+TSE]0LHPOeZ4dOQ_AL<TXBUS2ID?OZ<_1.E5Jf=:-9)C/GE/-.D(5=J
5,V;4TIWL&VF7D43^W:)5^9_@_8T]=F&VU-VBW+,EQ30BSY3Ve#@MW6V,@1Lf7\)
Z6fcGI<R5(a_3G7-[1JOT&V5M3J]<AAB_EC58)4,3\QFe:?NSTb#H/KP^=T[+SVL
[\b=d/f/P;Ka:M.VK6RB/309?WU=GG)Eb767DR@RAb=AM2E))bbN?ZFD1)W2-R_7
5@D7SQ[A/(+N-P?PXD(Z;RG9J(SA&)J\+:Y_L/-QAN;+YI@LUG1?)T6a,c;TC2A(
.D(,4OO?Z64T)\_YFab\.TDZT4-RNGM[B^-Ddb,1@A;(F:W#O?X9?.aND+5La(Q_
(1FOH>cc-VB6cbPKJfd[0^UdDa[d(0RMY#5.;Z#/2:H37M0.[UK-/1N?8L(I:eWN
YW3c(c\F3:d\5f@8ZaVWENMb/N/WcHGbN-KA&_GP3?)[X]b6+CCFUY9MZZ&V1S0\
NB]AXFdT\S<;]JXC3D<\[g2NU22,YXa3VJQ^LV3(&OW]#e)&(Y[g(H^5bNPb8&:K
8d,71_FQE&H&/N#YJD@M;YF6GaD,Q)H;>Rf/,[,(@G^J=9.1<&^:\_T(P=X;[CIB
EFc=7c8ZbM:aF07aS.Y(S[c332V;AU[VCESf,/R=]S.EY6=a[Zb3?[V9,B@BGNP.
@f(T7g;_UBI,UI+/9YT&TOUI>B&df8T-Fg4(^>6e#dM.4Df1OK9#/#gLJK4RX0?O
?.e8bDf;W]4ICXJO2=;7CVT\(;d+VN13UOG\HMQaKCKFObHEFJa.g@TQCbY63.:a
e#0=^SC_JGAUQIP37dK,?MU>3_GKDO5BfC[SGDN5OIQM&C,2gBc^=Z2CHI3>Z0(=
?H>L0\L]22aH591BU?a2]P\ZgV8UD4YaR8YV<7[-8>=9;^<YQS+7=\LB91Veg@;K
?;Ze^G#P87CWaGH&GGJ1I-UAR(9g#2d5ZYS7-;SG;0KJJMJ1O1-&5g_+efag8GGP
K>gKJ9-U1-@cGNI<AB1X1K)P18f[g<&O6cE0<FOYR1)-YV@MfAZY9PIBbQDc0=57
08XdA&=P]Y/8VXVg5Ta95f:K1@\>&bN9;D29T#8]Y;g8#3^JA&[0T-Mc2W^FX-\-
\=dT5;Xf7K_-N,b:_aVPF.5V8ORBV20d<D,f2eUX]7D5M8UN.+\Y/C5dKO525->2
QgbFLZ[Md-c2gSc+XY[?VNc6EN+T2TRLYaTJ-PK<7e)_HFC4f+2:86E.eX62M&I>
3UPX-[F5JBHdHO:L@81(FX#7E;90_P@KVJ-4GgcMc8BR-(4e=\Y2,,C?Q>aG05F+
^eF5D;>4J7]W0<8/]-_784\;LOF?Uba<8__+P_6Y&(I+OM5OXR?PfM4ETc5()<Vd
f73JJCbGdSSUIM,EH3be3GDaO\L86])6cM9<)V<SFT:A+CG?S.VI>21I=K7\=QTZ
AC5+gGKPIT]WF_+e\\?6S;H&2/YU@:R;UNZ@[&S9WCCUI(NeM?AQDTC<@D4GZR><
_<#V#TM<&5[Pc7M?1.IE?LBFJF<W?<7@MBMQ<N/3\\L&cLS^,GZ^6QRGeX\(dD\[
IgI)W6&OV]MSb5_STTZgY.V8ZFBQ-2e@RLfGTZ;:a38AFZ_Fe7aIF#eA^VEPX2+-
)L<<G<MDd4Z-+cB@8(EQ>LC_5W>Z9GdQ=cOWLGF_/E3^D=BX?\[Zd-]8cg@R_EYW
dMEQ>>]X,<GPK.HZf/K5CT4UO?#?:#?SC3P)Q57=f<Iec)S8P4a8OSA9G7.1a^H8
Q;4+06O[UAeW<cKIcEgQL4^.)WB)RE+Qc+ZOdPc@H8SL72c40DRd:I<6OC_,&]C5
6XdTF-?gD3QB<O9;BW/:^6f3H7D3)aUaM@8WRTO=1^fIg/CU.4Q3H8(7c_U)CJgd
cSTKD2..L@&(Y/fc&g22J4\[Bd?(@?UWI3eM_GL3]/8L@#f]0EaZbaJ\YU,Q\2Ua
9Z8Qd@V@<f>A>)(-Q>-:#f09<L=CJB_X;DO1BF,Z877WRfXT<+U._?WIF5@S&4[;
[S/fMFaAZ0VMe;\J=5@CO/G5aR1>+-:0]6P+)Fa&e)TfY+<];CXc]gOIH=QOFJ^)
G(Y(DXN0=(TGfYA;?JSKg^?Ha-618M>eOFg>&;8d?JWVg5:1WZ.T&;Z6[UM.Y&>)
R56Yd[Kad2O8&:H<5L(a+ILg=)>2&Z@O\>(H]]?J<]>F&?>R?.N)UeK4IR_ZeW=\
Y0U&3H=83Ke>3dBJD0eaPGTDSf2#eEPVTFf:WBSFe3_RF=TfDRHZ6T2#2@2AcY]9
T99g@7H:TffR9Pa,.)#GG;HOc7TS>_CBV72=CZSGJ6C)TBSBDg(3L0D?E+Z57#2P
HbH.HK\N0[Y:K2-24DT:f6e]?I<.3^H<<Z;g#D18_-S66BB?9@:;D6H3PE\ER#BR
:R(X;F23OP._D7:<>2AIgOIN;5K2S-PIDQ+W;W,0H[G@_CeWAf,)CIG&LX)CD7]S
<CV&,Q,#/^?+<e1&g?;E2S>9)3OA9NXdAd^<J_QP,A^N98+06\XJId>&G.(A4]DD
Kb:A?Fc2\PQf[21H;TU^FB</5SWf:M@SL&baLMP.9Z^^#bUR?c9[.T>\[^WRM[YL
EV.#fc5FM7-3OAF/)P@NWJS\[eF#^.X1AOf?VF^<CS:4/DIA)Za6Se3ABB]K1Q1f
GMf.J[[g5:6NBCOQ1.]c8L_@UaGT.R3Q5^[D_]\g,I/cN.J5+<Z]Q52DI.fTA>FJ
+8H(@P+?9I68G)ZY,Y,C[^H0^DB9HY>;X:]eNC)>?1fP:)YJ:b,]_4D1<&:P:<=N
4,K-?Vc4QcZf3KW&X842CQAIa?>8?25:^Ydb.S2P;g7-+8476\MWOQ1fPTU>EC]E
#KXc22QRH(>@g,^O[LDGe0P#eZ4P>XDH[=Bbd,T0:JTe26>OZ/OIY/FBKUATKSL?
=-(.eJMO2-e6b<WV53MLK^M]H+B:e?8@ER7d&O?-R0K707@3U_O)8W?SXf.dfZ>T
K8I;QUc2.5&P0Xc?R0-X#W20V_JRYH)SG]]9S#Rf=5\B.&+CZZS5F1O3CB,8PL\;
&Y5SE(&\9X5AFD#BR2[4<N/#30OO(,FX34YE&1Qg+WbIB=OPH;T84T(9X)e_O_QZ
CM221bL7.E2:a3X#(C9137B8J]7&96PV9V)6L9:2<V9K]S]C-]K[Rc1La^1[:MHB
Q?@0G.9A?V3S&EKOD@B>B@+[1XOOCKWQLfJ,ZM#RX-?V/W<+I)-ZB7_NTa,J#54#
6TIge^/([L\>KReQ+;c;SD1N5>M.a26I[-K(U#/7[Y@VX48IA<,aTF#\dR^8,3a/
Td)G./_XT.K6&LQ._6<ZYE+_5X0Me7=59e(;7M0Hf[1Z^d0^1W\O<L_Sc[DG+AK_
a#=X.#cP_\M3/?\=Y<6gF@^ge:BVW-]Qc_eFHcJD^5L[>W08]45SHMXETA)aeD4N
#H7&GR@]N-T[Q_bC5<O7+Zg@OJ.,QCW16T=YDf.A-R&L&^F[[)CY]F-e<F[=UHPA
YWdSc&+(b_TWA>&,Jb8QHf)fM;/^PbQd^M_?gaWK+>4+g)93;4MOFN=0O+:[T6bb
/d?N3bVZ7V^#bWIYIWZ2^DQ7D]f=egB[O,L,[CP]&&QIZ.ea4B?>Yd3/#2,>)a)C
42c\#EM.O48F2T2;@+:<ZGIK&Q9LK,S?@JQKALQZ_N6f0_?]N?L-.S;2c]&-&+)O
TWa7FgSd:M4c2[JagY4RVI/_F:.bZ.,@V&M9GRN3Mg<,e(^AFd,Q:TfY1?0QAYIe
9g[.e7;5We,PN,^c3?B^T]7WS,DEbZPGFNaWVSg;4C2,<W<]cIZZ24<T?IBFASS#
d25gFZ1KZ=:47dQNEQ)#JgA3bUX.O+&;K)Z-]KUQ<KB@7fa+HI=D@Qf3MQB&S8]g
aDB&8@N_gVg-#99:=Ld7<)bII9MO0Ug<bB97&F3BBTG[#X)<7;7V-b>I&E&1:[;-
9J-gLQPL#^.=G7g;P+1>3__RdD(3c5+A,B^9(NfO/;1+d#?7,gYJ@,D/6WA6E2Pf
K5Lg11F2.:2Q4Ng\gR=9f^G)c&d^R@55_5[LR+a\U\(PA.5fV94dB5JMDW]UXcAF
\L/Ud/C4H4D57\RY#([U\8^=^4CXQHL3,0b&00(MJ7I,0(9a)XO6WA:LL(^JcPAT
@a5<Y9D^4<<QeRH9K9]LA74LgQL?M0\=)4AXPW,_2H<19DG\OTHLS2(GQG.JOgK^
#c#.AUdL2PTB4,bB?>_,BUC]C5[e-[)J&Q&ZZQf(YCW[^c169=&+8>cS-5J(R7a1
(d^d8DU]a#X.KO-H1@I8-=[616<3DdAPWZWf=?WDF(0>CN,g7Z2RLa=>=4(gg^gU
1LN;+FN?45G6H-NAI\Sdf#/>2R-WVSV/JB5SU/F-_.H.EB)I-Sf5Q@1L6(G#&S,V
[NNPFW^M]M/MOB7]HO/PR6-BFERc0e0M@/<14:G_cWIbEQ@U72P2#F75D_X-ITD>
SL3PM=VFDTU02daf1>>QL:WNQ0=<)2S-GQ.FY@D-E]J<1U;#&Lbb^.:6#J>]T+&[
>S=fXfK6GT54-Y4J\OVU_,2YH,fRHW?-5G&UB&bedGKPDd.)P.6KHcBO?RWJ,&3>
4:SS?-2NO#+&e\.dB_7^Mc_;(V.IdV?Xb+_HM@)F4,SMF+O4,?SL6?fN3#3JOdLU
9QR08_K+OU1@8F0-]6)JPCCEf<f]E?F42WYcMPWSK;]AZaP-4Z:<C#OF][D#L>dD
N\T1(^2;I]VLN;JG)TY7;>S2Of=cG7-)OD&F@MH,<J2<PVQ1gII,6OX476\J[SPd
cU@WXS)ZK;LII#gWAN38\0?-B:=.a4:J<Ge4SJMf2;I;URO50)#IU9F<\6\FWWSA
f.[,?_WWgd+O&\T;_,#gVa((J&7^,HKgDIJ6a/&-(VWNF@fGc>=6V/9VE+]ddf)=
:H?9Ra6M8Bf.KTe?AW>fJZM&;8,+WR\:CG9W9:J3QH.K#BD0KTbCBK]R=+M#/&H:
FBB)XfFB_N2LTV2C1^B\53)];HaQ8=#QKK?:+_df=ZM]ZT6Y5XJ>_\RQ;2PEFJX^
]PV8U:gW]P-;?R=Y<R_5Nf<6]=U,^/KB-X&U_;7<\U@f?b\BHI=O=E/8cDHFQ9E#
KMBT]SdVGJH<cFafWE2XTe[A/JcMT/[N&gH\K10P.aTH+(F?LK^ZcVC=aAO:?5<)
[A@dd[GQE(<5ID;6G.A:&Y8g5C?eYdF9#9F#GN&64JW-)Zf><]#[?PRIb@\(1OOM
A/-2P4d&GM4I;ef)UT9@OM29OT&01ZU&6O@Q<:BHCF/@W^(VY55(Z_WL7)Z_I7[\
W.GXL(1/KDK[/,J1(KP/X=EDO3>>)FH7+a7]]V6(==bR8]D[_d[b=bH2GLFJ?PRH
Cb2a+FI4@KA761I:9MJfUT\O6X#g)00-E]LUZ4PDd>fX#.[P;5<gZ(&VJ3\//]C=
S<V\W\2<YI^eI]PF\L4,21VSKFNK)D\PDJ^UB_@^^0&g<OHf;Z=ZM0FJbH.e-MIg
B;O^S<(Sb);S9D;F.-JMPf_.\UH>,Y9fPA0fHH=?7A=7R(-EAC\6^(Xg6,J,A\c5
6c1^6WBSN7_#?[f[O&[K0JBVJ],B9GQ[7^/_NT:<c-fb-@+][gP5Fc#^6SKeUFFI
;;O_MgTW(A(&-S2=Q=0M4ec@QDSUf8LSE8[BE3N_,/S=R>4fZ3YH]^d5:@:8Z\b(
,.7UYV>=3UZKOa)@PGNY6aY9ND;f11Dd4g:D6)NcAaH5O5YW(6&W05aFCWWT<^YW
bOOC_W#R1U.N?XDUMdLO[.?IJI<TPQGPPa&ORU2d;&DL#+&eV329fM:4:A1B#20[
FfN?USS#2Z:\(dfYb_.b@@E6]_1EZ6W0E-:+/)D/9A<ab]a5YM#:,ee?a/2.<2K;
Q0YIV)XXe0VT,CP\U@)][Y&]KL3BHIeWaDV:)Ka^T3UMTG5<^8?Cd6P-<Z,]1.Z:
8.BbBe:2OMQ=K_)^P\MY6+U.#?8>3O785[M,CL\Z<)Y.JH3-dDSE_E&&4<93LRfF
OBgD>\SQV[CHe:Z?c.JAPGd<8R;g9UcDaEgH]05U4/E&c)PLJ.aESCCGY#(=EUW7
e):S^\E9N=Lb?e[^X@62R9;.^9BaQFV7^fE5EJ6_@e]?9=+C((@9Bb<6SVbgKcL3
):(>]]X&::8[#S57S7F;G7J\#2e07b@L?=9OCUZfdbB@5&KTVG^?Fc30.KB[dE=W
/NXLX)49H>C^7O0D7;:]5Ua46g)(3dVCTT_SC_N1RQ3:g;HHO6FfFH47/GV\WB#+
G3A)1Ig4-D97VK4Hc=&RACFcY])4ee(ScWM_c0K:9DY32^ZGYC(G_)PdK&8ZeB14
I/4<V]YA5X\;a>MJ9,R@)P<4Cf&EJM#bNJ)^-QHQD#f>IT69Xe]M.T;da;+4cI5W
,e6cMY\[\J^TcWJe8]T7]T-359/P3)d+E__+<<;YK@DM1.EPAL<PQ-P3YI/6POIJ
>7W2T)3K9D-;ZNIW,>J@5a,D\V/9>7AG3FWV[[cEUS#4dg7\Y>9N?I-_JVMg:G9^
<+6LUS#/V,P2E63026S<F<#H9]@W_XYWW^.BZ+KPdZ;aa>cJYZHG;IG0<QLg\B5&
JM0>IVL1V^P92[#>)O0Vd6d.X,)dVI,5>g3V4ZI7fT?LDe]R+FRVJS/T@E_M+PNF
Cd>]9aVf^/BN()K/FA&V):9EOO676#(610QX\=D7W)_M-gZcfW]3Cd:)H[?TQ7.8
,->,0/Za/PGZOJ=F+VT^d:4HG8/(5fM>WgX4CVPSKTM83K0@BM-bC<3VE#S9&VV4
U\(HSV4@<JWLX<^9RI.W)UE[ObObMO4O38ZfFf3BTKL:788cJ[>70[F3D5]+T.DA
#M&,KMdcFFDSe&SX3PVge:(##IeLQb1\EBE[CQJ=f48fG_\?Y(=4+8XQY+V065.A
:F&B@g^:Q#<\-YU@-/Qc.@>RDZ=Ba^cX@XVeKY8IEP5W@(>)e5\PeX2_R(C:O[F/
1NHFg82RfYT3=Gd3E:=WOSN?+e4DFX<TS9(PcJJ7I=A\OV>0f^.JfcG0<4JVW3@#
8;#Q??JPW\.Q(f]DC_C;VNb#3Yc0X/P>PHVS(&J.;RCS+6C-G&8X:Oa7R>LQ@?b_
TRH_-g>TG@B[b:M1H]dSA:7>SJ?WM1,C1A)MHNAFeNJ?=85eH)N.]U6H/e[]M0PV
M)SG.>a?C#d8&dW-VU,QYP1McLQWF544/)T4.A7CSSI(eYD-BRXd@BO-2#H?QIZ3
H,[M7][ACc3d^U7.Uc]eZ[ND:JIc-LID9/]4/<?AeT-NRAAS+HO=+QC2.UgWPLBQ
>3+FSJ/DgG<_8):PYQ@a5Cc<;3ScGc2e#L&^g[Y^M1BafM\L&K3R6D3Ic9>[[P/Z
,N1/Q8=Nc=_AGOH#C7g5;GX+]FaENcY(6f\Mg,ecM9\RLJ0KL3JBMFO+MI(@dE:>
+g];Dg47FZBNHbTfL8S2&:I/MD+Qe&c>QTHfZDQ0I<N8V.L7)f\Ua375\N6:Z-DQ
R-P@SC?:Z0V<I<FH30]+=^X^R9adYLAa&]+XTN5Q22b@fMC)Y9J<-:XCYc_ReJLc
0N3J;C?F,cc+34;YNE\B+b01(&#V[eZa<dL3&NRS6@6P=>Y+(FV?fU:I3e2KA[@[
KN:&RDfT2bV9:_4)T]bSD_Ta\dC2CXI03Z++4KJeA(3CP#M]#KK#<Gb7b^^U+9IT
HU.H6M,\Af<^MVWca92UBJT,^K_+0aKc=X1P)4fXIg7)c\=e:;eO9<7ZKZ?e0@2O
7A3#LV;K(#K?N4KT4BKC[B-^UW]OPWV38PN4JS7B2HMRc:5ZTJ)Zc1/KGY\(S>C4
MQdZIQFSGgF<T2@<aZABJF?_A;;;KRb5<CC,NcOC7,HN],3G>P^g(/]]=X;5TgL[
d;ObHI4aGCBf-@+(Pe()NOXfBfQ?[NNH?-WOYaZIL+aG_dGB/],10V=/<QQg>A9L
>-\Z+<_QN^-0Jg8\4S6EBa6/^;S.=<W50e8dc<U:Z00?.9KY96ECRY^Q.@c7;2LS
c)+T,1T6)(\.[IK8\C>5bP2NaAS;A/8g2D8S_6,?UW:e;ZCbd3_HA.LNTBI^X:][
3VdBQ_g\6EK\XQ,C30-?RgF=OV:eJF@^e<-33EeLgV;@T&:e(_WfEQ4+==D&1E.(
5S.K[.,)4B?fAcT)2V0gE-(bcDZQL-RIZ(CDFUf[+\K6C@;##4Xc)UMb,DaY\.UQ
cc([Q\;]ed0K#_+aQ<e-G)H<H/JJRX<WMICX=IY=C9T+VVK[GG/Ff#[?&0UD/dJM
Z3b<2B\@[?-:.P+<4L\LP&d(7S,#9&?:>,8>7fMM95:#KJ_R/AI4?V>&<BI_2B_d
:,9OD,1+67)OZ)2NFY.NGde-bWRHKB(EAIR2&E=WXA?W0P8]\X6\1#cLUM98Pc0M
G=5Ve\T]/;a-g0GAM9f3P@J<B\E@4@D0c.b;/S&QTeI/>O\gAQYB;8E73I\ML6EB
bRGSRd>\2:\+RDZ#ICH:O<.Yd6PSCdXd>DZ(DWef3CFM>(-(,cgX?)a:a,AV(bd=
;(-B@g#Z9D<BW?SbVVFb(068I&2f_JZX,<.bN]JdRZfGH1S-J(\,KOf,]8(3E-aM
3P@c[>/79CJ+CJ#C^)16=,MO;.LC]Ca-KCb5N)cXUf-E3O69Ega]TN)Ie==9QDK0
JeX=e/M,)_T\fYVA1MQ3,CBQ,@YdYLL5],YS/VLI-4ER>(_PRGdZY48V3@>L1(T6
QW+&NVdE@g]c&:\DO]XOgE2-d3+^WG?@b\X2(Ig:0[FcdfE(K^:JSAQKH?X=OME9
TNd-2H&>ZA73DUZ7JM4-VfZe,4=X:.a/39=2-NW7Ya>7U&SNGL2a:/T/AUYF)>fP
J<X+>,(?UUL;#[O^OW11ZQeA+T^)VdWOQbW5AP[]KcDH3KO;+bHZMW?dH+R4[9-_
(_CLZWZc3=SXSKL.;Q<V&MA6)QR)[?,9dA((fb<,G]8=(V[FT/Vc0BfLI((KN-?D
B^[6EQ39#G>;3S8,c(/TU/[,dgLAXVX)Bee^W/c9Q#L^&SA<1R57]ROZI(UN108d
WL-Zd88+LQU2<Z@/d^[PFY?LP4DQ@d@S3cdRSbC9Oe5SDV&.3:=:YV8O.@(ZA[:>
B2\96/6_M=ADgZT?O;afAA0N=@d9^L&c8@>&5V/L6T,;J>^.M2/0/=MCM4C,AX]^
=YfE#&/)[ZOEUH.SOXU;5K1TJ4L,[ITcG@F?F&,0.(TB10/a7-ZUE^OcQ.UXI4gK
)C6D<#/f9+JZY=D9OD&UX4&cB=6PUXQ1[2e&c6;@C3=43WbOHa0#7<7?)]T7P5<6
J\#VJ?K21858N8eN?W:dZ^:H782M+,NcOT5-O(7a(1Xc(E#TKEfEA0X65M[:8H2=
RN<F#:=gd@,#(9WW1:;OJ.;>)G@5-RC2L<H=G=7W<CbWA@710\5\9-DObHW7b3[P
N0-&+W8Z;;9\KR0.WD1;:Y0J/AdO_\E#-4X/SB6VaND^^0,cb)C&>JM#/:ZG&^^B
/268\MQ<eE/RJ\KC@>TedXdRA@V?N;PB+?B_N3>.HYdU3>#F>)Z.,/E:O>^L8/#K
(2>2:IW2HJJ/ZGLFDP>D5eV/LAQH&<e3\\6<(]I1EGJ=SfS4Z88;8_;fOd5eR>GM
\-ZH74G=@cBMU79cI3B+&I68U1[;QACYX;BRS<3QB@e0,HKL)T<[]@=.F,a4TMZK
EN=@d&7D@R;^7f)75-^-=C;-I+/9baVLJ9UfPaW<6:30O-/W.>H6WFP=BT571Z_?
0W=a?@\(KeH6&02>53&^8/=c4b4@I6S;--RS1UN5S?M3GU@RARd;K@c.K;Z^JXY[
3IUUQP28ZKC\N,N4,I^\bC6S_MgC.GI0)-+[fSWS,K?;Ta59=;V=WS7WOYT9>7FC
#F&^0S#J3+(O,<ONeCReRIQY2aRSX-0&,#>NN6R\[DZc9Sd/4g@^a.cGfgQ[,E0Q
>XYCJ_6Z6-faMeS=?TR_;VO3beOQ^_G@fbB9[47WWCf+FCZS3/ETW6R,;<e5U,E@
,A@WZeP9c49)\+S:-Z&<e=c42,Y0@5RN<&KFHU+<HYT#^5DSVGSHQB]eH3e:1K;T
ZJRCB#-cgW[2b]@-ZYYBHJCDLF;LSK53AJ]JH>L922/HWI^R8A.3M-S](-=dLZcR
=0O4Z>^5Z=E4c4e-JR>=2J/+WS3<X_=dYe2#7c.:SeZE6<Z9I[_P3c&3HAV1TVF+
e9X98B\\GW(ZX6I-[Z,\9O3:NN)UZ,-c4^-ae[+V0LP+/#@0:7&eg;abOR9(#P]K
QFLC@g:HTY-SfC_2-Lg2M\f+7G04^;T<^7@4L)M#,ULaG;a5\88,PQ6QgG:=fN>#
@R\O@ZJg@ST(&]2\_98S\,LVTSVF&gbD#^NdD7g.4G-R?;Q.degH6M92)gZU+K)0
>LM@2?Q;JBYg;eb-R<NfFgM+#<C,5(T>G-^9_CXH.I7)4=W@[Q]W;(8aSBHDPTJA
WUH5#ZdA#VYU2gN^g6(8g674=1@\_0A1\R.@&aP.-+VGQ.&\\4FD.>?.?d/e)Xd;
Dd26G4aWCU_3=DG(J?:5:g2AE18C2DP^/F.D(U:)NA+a8cEe_BS&JYE>I3dQ9-ab
#B3(;YCP2LVO4VId=N#08F,QQE?^YAQV_:8D7:J9\EXKV/Y;G^b+^R2D?^?Z8IeL
770.V7<(J=<K(-T#@1,EP+^>=Yc;4;K(,49fF?NN>T;D)+GZ/8P[GY)0U9^1K&7.
8F\Ug&LPDYW882;?TYaS:(b,?e^eY&9eV-=ZGYDbP=:DGfLc?Y_7:J&HBQ8ILX0&
IZfMY4K1f+ZbZSC8b>Gg6NcUKSbM9O=/Z8cC>6<Zb3B/1=C([LY]:g)]Y6>^f;TP
\b\G2L3?1];;M=98<ff&g1[(]^WHHaJd[P.Z<(gF_GR?64&#N\+U1bZ0B8#Ed#12
DJeDO0cH__5]/0F8=0Z](Gdf+,K5-c2>;CbPEOaZE<I0ZO0_G6+@IBT.G2E;U,([
U&TJ@.TZ,g@F\YMUD1V1gN1cJUM]0>/<8RJBGK8d_VY\N.K)7QETeC7.A]5X/_(-
PW0Kb#KH&WfUCSc0XH\985CLW99(AOJ0:\B)H7G^cN8GNQ#6dc,@F4]6g6Q#R_0g
6SH,(:c[f58dNd^>+cEebd(\19K3H5;)P5GEEX#Q?)F)4-,]JF?WDWUE_OL\:>QF
X_aG-89IL6bf65bWg#g-<\bLT>^VRF@=Sc;1CFCV9]X]\51e?LI_5&(G4.fM?Acf
;2[IQ6JX9WGJ1-S?@X;9/0f6fVBO:8:SK7Ec,TcN(5[=G(9(B<:TP9)T)Q>COHVU
\SfXd0CI#C.5WQG/?)aP&>PbFSG:\QAE+1ESEeE\E/G]EGEAP+a<]#G1bd0E9H4>
OIW#>D8XJ40O)+WJa)M569<f=F280g3,T6D&&R0f[6:B+@.-_G[YW9F83H>bgXE\
B?-^bT2_geKca0-7:_J^[;6-f8IF(@;Fgf-Qebb92:0400>-MONd^8)+H?_/?&Nd
M#cFD4B?\K=G\=e<a5=>9G<eG4TJE4SK5ZG8fCdV+W.6G+7/.Od\OMJPIYb,4ZB,
=S^3>I7>>\5.Ief9gab/1[7(279P/T=)S>C1DHJ<V\F#Q:b&B[2g78__ABP_4cA>
6MQHcc9/c71BdS(]Ie]D#Gd10gFKgE;HJW>BOE(^7gU3fD9ZBN1=@7#IL@EdA?TG
&??5#W<:b[]\AQ]+P)dad]eK<@3aI#X/R7?<3@KIS:bYb+];_<./FZU)<fTC.@0;
;gYcJ0,Y[4NH=bHF[/(KBQBBfL\,&9YV=TD(Y/RN)16/4b?bL-fEG)4#]/SN-(cd
?bb8\QP=MFdR=<GCQ(?WMT9ZLUB/BB9(L7HYYA/.7bA,aED5W,(E/RdR#NWYSg&g
M\1M+@RYFNQ>E0J[([KRd6@=40#7WeP98(A>TPfN^cb&^EHFe,O=N3HYcE>_+](6
3:PfNa9BZf@IcHW>8OdO3;LXSI?0a-Me3KL7Z&=K2@8Edc9@PP44-HDMN:>5^]=+
f:P5^;c;A]A9Hg[cW=.OcEg/&Tc._\_WP]F@W@,B=,2=,F<O()@K&A([QH;+R+LG
KFLCC-eaDB,Z;IIcU4,3[R^#ffC;;=fI\PG6BF^,,eeVMBHQgZg:PAVb4=Fg.;@X
-I\W&[bB1\NTS[83,?5EK71B0aL]bMN-.5PXTE4B2N^A[L^40eT4(/e@APR[1A[a
O3X;E(714&^24269Vb\41SbaH9L]O7?VS5(\NCUZZ.Wg85F;Q&]Z-Kg&(:fOQQ,(
HUKPWZ?TD]6?2LN;65g]8F&.G3Jd&G-RSQ/7Y3cAY4O14]3Q+CE:300dY0;(:FcK
0)bWLOD7Ia;+-V,_Sa):NX2CBF2>NPeT4.Q;C-g_HcXR\C2B@a4U\@/JV2[N9H#S
TCQc[Ha+^L2&GZSNYI6U6.8;fO&Nf2GI/X\1gUf8+MV9;)F#&S7X-4.#^Ua:5TUA
42&@#9-QgYTI4PgJE\TVY(e6#T;:[>BFYZ#eO#&HHH#(cG20H0N?U>(/]\2#bB5E
+^+c0/T\V)L.SD/9ULO[0#P]4BeB+U]cXOZ:.81Wfd9ZZ#fZVXeU/@H/_ITQKV]/
b3.ALd43dJ3L.IbTJ-UR_V;#&HU[^e\XEDOI87N4E2BdQM9;HOTI5b]RWFdR]g+E
RW6^06/Q(H)+[a]U;0FE#5adcfVR/&,3L<DIQ_1:A4U-ZVeG4X=BUXQK3LT:(T;T
(CgX\bO_95eId/\VEYPd3+ZaX]ECJK.Z&GbA)>JX=C@#4d2Wd^YUPNe/MX@Y>&e)
-eO-,)@N4?>O8=>e>\SBZ(7f1/JEVD_c7\[g]M(.M796ZH6d./XV&TN)<WBP^9;A
O6&/b<PMLHN3.7FEC#>Q;Hg6U-@<N#7=WSZF8dVA,RAeb9fBW6aEebXU5L^Q,@B5
NWVb)0?<A\HNXMe0(4e@XG5BPe_2Q8:4;)L4@>NOQ18C/Y@UU_@#PWJBU/TRLL05
/U)5TabN/G@P<dUYWb8D/#.-Y=:0)N0J:NXcVVYJ,Q+d]B/,^?[7V^12JGL(MC2:
3+9)T]MR.6BDH\B&5DLVWAB;\Q4Da(K7&PAUC-IFX?P)Q(M8K77V@I>THPYTX02W
4LHH2T3)GV7SBYMB]9<ZgOZ.;.06:3ZTMX&YfFGQ5df?Z/0U]d-:Q8J5ScOQ4fA=
&&&W]G-T_IF[H\A>+TSOFMaHSg>PcX8UC0/-\VQ5O2KGUcP/H3ZMJCGRX8f&@+OS
4a(?fH9E;>^=#C]K;7GeQBCKcDYUS4WQf6W(K2VWdGWE&JLMa9+>?]YJ@80PBbD#
fN#8_0&Y0a91Hb;g6VLe=/1AIA)(gY:@gCSR,;R]HX7G2TM;FI/U?OYI[<2<R\,L
+D@eR@,7)2B4OeK&c72d]VRB3S]--A4@T8[A\JK)/H:VV]ZTK\_R:8+bg&R\X#V2
_B[3LB6\X9C^WIg=?FE6/XUJQW(5Ec>gfDDW3KIM,TWOPUQC>P^?J2/)7\\1Z(8B
0@(F<)?>GI((C19@-BB<CXZ[N]eEI/KI8<B[?F/(,eU+TP&[+#D#aQE[_>Vf6Jf]
#IO)TD>bII,G(.dKTf@^R_\&Q0);P;_QHDJ<Wg6;JUcGP^6#R^3KXS8,NSQ#V.&M
8\W5>@&-)6R=3]SUV3HGa:d[\\S]TIP51a?WLESe_K_2;M)U:->H00Qf]3BXZR9:
ESa49#M:WM=130MVMR57SE3:C[4MX>AEH&5aXM>3.G8#_>X)YZSWV\<_0.d\:VIL
:P-6+2=2/W(L1>0(U?9G55ED954S19?A0HFV_?;a@>/d?)-MAeFP81.Y]4-S6<N-
F=0/C3]P?CW&XU@E>:Tf?,F>J77b;D/D;KTKX2XW.OSBef_G?Q,B11F4\X]:X_:B
4JbM=TB,?AKCJ,\Q.EI2T02BP]3-&@ZK[H=6G4=?0DO?G90N:?C_+\Df)eUT3CF.
WTZAgf71Q76[&=(PeM6,2GBb<IXcN(g5)2&Y&>6@2Kb.8Fg^G[XG4OEE)R@7gYCA
bc9dQ2MNPK=4D&32=HWc3Qd9c?1O23&0MZRW97fM)g^,gXGY/6EU-V#5(dN6<BB-
+dISGCG]5UNd[MSL<;:A)<FU+B;EMVfMK;85&@-=OY;+()II&B23.MJe?I56I_I]
4OX,(,9Y--6-R2_K9YE.:4.4]B)\-AYRPf?(+WH];O\Nb>&Z+31\-1ZgaT2XRH]6
KXOM0g9Gd=:Ib-<>-3XP2OM2Ge2Ra^MGPI_\@?/aE74NK\<8P6DKa-D;C@REZ+6Q
2M:2Q,P4S[VK8c?C?8F?UHIcAMX?H+Y&P.gP0,ZLbH^OIVW,+6^EgL=17PVSKcGN
&K>D,6:0((9[,P(fLWS\J.)ZR\G;HZc@U((_/cg.S#+&d>=-.F[+bX+Ed9fRc.gF
Q48IK;?c:1M>>)@T:H6,R+DFG#MOZ#bMYc1HX5T];70SdaOEC+[Qg[VJAIX,L,Yb
Ee:<JC4?DZ.gO3A7O]OfUUI7dGaI2BEU\d=Re_1Y5Q+bb1O)TIDKD4(3;2,30=-D
S#0)T&#c&H))DR7+QUWgSf_IY^Gae&[-0O8>/fOF7/#>5V@,g.b6S,KW])Qf-IOe
[#QMU5b;A2(]>fWTWK7OX7O50@#-?BT5?INef<SgA]0)=F^13B>CgP<-M/:Z:=M6
:;2XA64I-1.-?gJP;aFXb4>e@^6;UM4bR-R2=4b=MTc&RL^#g/R.MDD)gB#?;:)^
4:/U0WV&_0_RKE<UU-ac7W?6^a4/@e&?LQ@XZ3S7]?EedUGMc@fa5d@J<75^M^QX
Nd4fVLGY51BW[T1(1+QR>+d@->5g9?Z:CX[&I2R)HgHF@1@eL3g0=5Y9.QOX/g-e
AQ+:4ZAVR^YUB#>0]dd@?S6KZ43=aWgRPbA6JE++NF;1/O5M<:<@,W4Y3<QcE/W(
.fU)/FO2D^f.D6=;VfJJeKLR6]<VXT7WaXM:L^;XQOM.Q0\I<.O.GG/82-Z(57_d
H1H<=NPHC9fFL8\/&8P,ZGL?\AeM0ZaDSF&AH4g[.\Q)6fO?B/P@TQ0HH=B1_de<
G?-9<dU,R_>G1N6+J+T,GX&gFKfPGIc2cE@KHIEQ9/5g[OZ_QYPZG-Ub1.0O^gfe
gS3f18(X=GE=0L^&AY01ZUYJ-:VCO:23,M^B8QfXV1Y79c=]R6<9bLWN&YJ>.K@S
O9M?A)__+c,\NPMc1793aUc<0gFE-9d4[6P(B(H1+9W@1Cf3PBULH)T:7f+CZKV@
/BA\Wb.NWP0_22WfdYDJ\:6VC/Q>aXc_6<+U]6C]#db<;SUfI(S4?\+H[;cSF7.Z
J.X;_QW,+ac?d[EQ5K(;VI0@dKM5+g>H7Z;,I0I?JCR&YD6@G]:V]D2P)B0F#PGT
4,4S/a<:=6+Abda?402TfO@/6JVc&MAe9<F);8ea@X;AUbN>Q4;9DK[I3O[.(<;(
TaYLe;51;LM,ZPd]L:1bQ7KW,JC)G74OQc6<K>,b:4/L9YE2?C8V?:BPZI&W<-_@
)4FHcF81+^S1BBdfBU?CG96.3b3e.Bg@KG@@:KC49LcPc_)U[,K:g.--QcY^(PZ4
P&F8_VII6ATa?[J2ITAI\g1?KYU0Q\Q<T?G;f?=,>1,33DTf9#QMUR&XHQ&T\#C.
U20)db7MK0P]3Cd2/1,UfLD)PMH/7U)1:78HT9+RE.>cN5>)O+K^G6S[@E?F[Q:/
R>fLg4I@X-,_Y:^cJ:MFNgYGF1D;)X2/(Q@JHO^PGa;B<KRYf/=.FUB<17D7KL[(
8:?C)7G)a4EfUVGQ]V1MYGVaIZcL,OAJg\XM?I#)[WEC/4dV&,TLC/3OVL:GM0-4
7Qe9N=\@+R\Eg]15558S[]<bfCF61D;-U,T^9S=1TBda8G?7;FF?(69T/0G)]&HZ
O;YP0#ga7^/P6DG/H^KFKJ_H<UYBK4.;.#+,C,cO2N.U>BNZ9SEQ^N05/[&;0CS6
29G-@C2>9Y3SK(3(R7MEZP70-MFRdfRC(I6+dafU-bMW]&aDR5&Y<\Na)B;\agE4
fFO(\OSCBN/-B?dJH+5WGX?,+3]LIGN:X/43T2+0E75O+8f.<2V\O(A47#67@>M#
8K;X>KKf5bU<6=WH=.18C&G56^FK,+J@X/\]_XEH4g@W,E@0OUVF:GF5M\0?[R]b
^7?USC[E\S\dKS\=]gNMcPgGUJ^\NNJJg^>Y[G)[V)9[EGT:1YB,GEW.:;0N>R<[
ae/LQQ68^OA>9U^3H;VYZL27;)Z#)BPcF51/UQ0(V^V-JGM,1SI1_;c7(.5FBROW
=#SLf;G7:#Df&7>K5+d\3]DSCNe[>c,c5D=7a1;W)aG;QQ?[FX:@N1A,[+e4;[.F
4,_##]#:,Pg<(gR;b=@=b_MC804eE7dWMFWR.KO1d--#Z&D/Y?@Cc[+FV(&UDPgH
U,e7M.=TJYG>Cb9PUD,/fcUDFVFTJ10\HZ@D]F[QGV97:^fMFLgC;]9M()7RWUT0
I4\3]QXa&+(HPQDW^aNIB8QN,gLe^:UO@GRO>MJA&WX^06#K;/AD8O#45.C\DI0X
_+3LMTE#f[7aQ54??EI31<O)?B/OOP7J+;90GM5:,fCDXJgP:(NXPR8@3-GZJK_:
+>dV:KIVP+CU1E&:.EH<[]J>.F)MbTb;_4?1XfEXJc&H/KeGHNBFg:6TS@f@YG7#
ODdV]>CZ;>Sd[RYRGWO07G8PB,O@P6.>0=ZITdK:;g8TC5N<Z2MC:fKS\\Ie8#Pb
]RY:;e.02NO=:9gB^F3eR^;5M1b@&C]dP^9^+,=>[,29&(O]cB6=??bM)\PaJ<I-
_>-#GMOHBDT=cfY6:&^]P>A.a<^Xc2Ib]X_ZZ.d0?B:K(fcU#56EM4YP=W6L^;IP
?SUA<_1CZ&87SbcQ]a)Od\dG[,=dL<RAH(&1VS5;;d?7Rb[DL&TVIaAR&\2MS#4Z
<Pd46094W>LZJJ2\#-:IcgcZVSV\+DF6HJ+D_bB2>f3#]26eTG4B88(:-,CG+[9&
(K_c4,6LZ148Dd&>aX+Ab,f[/U(e?=,cGPb@=)+Pa(#O1X76(.dULg2bf0Q)4e_R
=.PX]83.:9)8+9S-/4YS[QL,WR=f/VADH^Je9D-Z4_eOB72aHIX_T,H?M<+S[-AT
aYE8b)GKcJe:I:GJ.U8O2Sg@?2c8_/[5/A20IGHQD,5AGNcLb6VIacG9]8eeL3LQ
,/,^5DY=)XEe&V<SLfO?2(,4X^^4fVF7TBL^4IcV=BcR@@PaQVbg-AKNC@cJT=-:
:3CVQ50c[_NW(I.O+gB<VfM)[egb,6Y/-]cD.VN7)C8AgUS4R4T;B86#Ye)J5T30
cV(]81MQVAe@e6Q)>>GQKO36Q]G)UT(M[7Y<W?UO1H2?7\0:9463YUbSET5/:#c+
[DVGNO0.=1=\C9Ud#&KP;>COCbMLZ8BQ&>)8+@AgNVWO[=4g<S2O+EEbgL4:Xd)S
=RcAMA8>f+G[:6c7Pa@DfFe@^YC7T6CBM_USHdV_T>9<)Y2OZ76:8+DH_;9+YT/N
(b@VK+V&0+MMV)VVKTR>9#4UX>,TVVXD<_ZAQV]4NK1cI)X9,T+5]XK5;;#@P4A?
IZ68)g5AM8A3#&&[NP5X2S@3-6=@H[Q:G[Jg-\HaJT&+).+ZEX>J&/=0V+b#ceAK
Le?TAK<4A8#)d8OK@I?EGFA36c:bee@B5RE<Bf+6FWD(U=BdWW2FbL:cEIKAD>/#
N7,#c@=WH0#gP>21NfK^J>0g;7IFd&S-\2&5WbI5eN1GFOcTWQ7[fN@QK]PB;NFZ
BW18FPPC@WZfGU+&3UcBX)Re9c,.b@UP3Z@+RK[A4E5dDI#(bVLP+2Mf@4ZL.-K-
9f=DH,6fWF7.A_R\[6.DbE>:M2HF7RBGgN7(8CY1G?Sc,LB=))-B@[,]1G-H]X05
<OY-bZX+dTIZUK2VT:bQCUX\G4CB=c3\8/3X2Ab3U(Z7#==)K/bCMNV[+\)COPG7
HJ;20[4#Dab.\])W.:F?.Y+9F3N3MH1XSX;1Y)D[]<,D^SacMQKRZ;aF(?5a>VZb
8\I#F4AO>MVIW5Zef(9T=8XPE>b_&8GRL\EAOFJ#]+Hd9U]K&QM2+,F&9b0#S=EM
@]6O20YXH,?(_f:5ZG,ZYS,NO+N#VaFUQMd.(IG]ccGU-a;F(W=6Dg=F)#QU/F^&
V7O/@KRO])^OdS,+X>,A-I@E><,L/XQW<P0F/8b2#8.EWUG?A0;5IK9G038ag4<S
dMaL4VUEP?dH-^(R6II7,2E\:EBTY;<\P.G.LY3J:IAB+K;:?CMbFH.;E_YZ,/<:
(8(3+#Z).Q\^[M]8\3eWbGbg]PP9&\-TH4^V-ec\,6]a>7[-8W8OB5^;,]RUcVZ&
=:#=9CB\c)_dGdEH4]0eK\bXAZfT?:cGFFQ2CLEd26XJS2KNDL2#-=PH,g>(IA2H
T253G6-[XDTI1dM>.DD<5a?(GOBR3DC]2P1_:&+fB3+<V=_CX1-7DA8O)8f+&YM@
JZDRD964TWI2YJWLWU]gfFY[:?RK1d=_<(Ea[?E8+I8GZ/G=FNeSPgJ@L]_4f:EJ
T#a98+^@Z]Lg,NSBc3=JPQ,D7&0Q6g&V(T5FBaN]0dWB_YIF&>1S[&(HJbN>SVP)
aD&S.:[-Of?FW=6T11=e5B(?A4/=//Y/PWA_GNQT>YWA+U^^+U;-=DA1dI+_B\,C
CEXYA?\ZC4E1/K@VHC10QdOO3W=YHHeL6;C#\O>2=-R@61[OH4M=^)HH[7M]X]<_
),O\H,SU<+KB@=7,BXM_V)4aSM[/H_/5G,OSdYcK70[O4g\g-FH<[dIJ8[da4JH;
8(H80g;XZ?MMM5?HPfF@8[XaQ/<:BT8MK)6>;O2T=J708MX+e_8eLE=S7Sf1MaZ;
G-->^UXcAf)>HD6H.:;\bQ2S74DM6\gRJFU[QORN-4+=VTWQ5[EIXC?^<@H+CU)F
aeDW\3W(gVN#[ZcV@ZV4D,U7^AY?<a\2U6X&N5?;5GPP\W^(fN=>GSG0E1aR.R<Y
OG;>W]G1d1[O>..B;,:0YY?^>(^G#(JSdLg-/.YZY[=^aT&BR\+12N<WBbL+>6PP
+,(cc6Mc^c-X955I_)AK?MH[H,:#3(N3c\+8fIK]CQZ@@c/Y^a8KHNY0>Z=fPKP.
O_<+GER,T8NNN<ET/0+;ZV<1f(CgIW>D?fB?A/T<#[WU)FW]@/3;8#YI\;6F(8;<
Xd1^?M@&^b-ZI1^#ebMBM3]2a7UZ3@Y>e8>UE1d79b3=XZ9d^P[g_^R7#YN;Q<.8
c5J[20-X<gEZ10WM-TL.Z>V&5-<1^HO(C,bPD.A?BSE)[;>02e/-/+PAEHQ4>=WV
ec&d:GDf?O//FO8K,SbQ[8&\+2TMdN2d(57SZM3@X12YK6Md&abK=a+Y:WU>LN[P
C+b=:/9L.1NbVP1H6WW^ee:cXGdPbNWf0,B\Cb+1U:OXPK8]2DEQ7eYQKIf\J9,#
.PFL2e(VGdLR8a?9Z6^)f,W>.(M4N9/9]FbfXDeeK>45(QOV&\U/3J9Cg+R>W1[1
(-CO,;V\;@6JAPVP99?+eb:YSEHZ[?LaNB&AY[EBQ@cg,-I^fGgT-KT,#Mc_J@?g
>VU5L,D]V1P&)O_19R2b&1C4N@&8>R-V154fNOI3,^2S<6NFbTM>]T\>7&#L&_#5
0ZXE5_P>()FBM-Y.,K19X;@L,#_<cO2>PEI[E#2.?[\QQ]T^<J,e4CDC)OET\8&/
M-J6W?=U0VfcE<5()9e+)1)&cIa[>X6>3FGQ:/,=J2c6Q2C<7^EY8[.4g2T91,IH
A+VE6BR#R6JNX=LFBY=4:+(K+]U+:XSHU[ECQ==5?U=#X/_TL.G#617\^HbL6N)W
Uf=cBVFbW?6NeI;/?7H6)VcW@QKg\fY>B./?5,PHX>FS;=J=;7&PNY4R8\fc/K+W
VYC7_e6^12\(B@M):9R_+5gYQ&CSP\,9NOWMJSV20J-;47T25-;86b_VQ=FZSI/-
:RJ18RY3KY_+dY<<CBe0I2CAXVRB)X2e?BY=DE39PYB;7X_6;M@CM9ZB9a6bcBJ8
U[=5A=^Q_?(91\]e+ZFdTCVXA.WeDVAPf>8b65^C;#1#8b:NH86d1gP)9P(S<05_
?BH-/Ncc.6a2@ES_6(Y9dD9-Q<KG5-SSQFT8#C9L8)]CSB0==FQ9a?O5b,U?:R9K
ZYX#XS>MWZ<g/XN&=LWJSdB=13I9BO_]0JX5g4):TDG\GEcS^,?T4JOK>d/aGST#
B#2_&0M0_g5A)5(JO5EI9@LYSaL,@c;gRWM3F?aWNBb?8)-F5Qgc@T)>JYJX<eMM
AA&U1B<=Fce3IMAX7<d0Od?&eE[_P;^/c9>)cX4;UB3N4eOO_[gXFC:<b92#G>7-
K159^GV\<K(W7C++O[\3:(a9d9WOY>PQ\-K<3T<<W<GVZBIEK./>@4.8L/@MbO?7
c,g)feeHHY>@]g27Wad#H7g2M04)NP#.KGX)g?H@d51(;J&Y8#B+?dI,>>aBAL/<
DPX:BQX?)/9;-gF(=1ABYb&D0V6MFB)F3H0e3+=N>71R\a/-5:],+S(PfDa&6^LJ
7.W_O9\7bCY:FH(OQ]0/<g]Pc#c#1eIgdA)I=,;]1A7&:X6e7882QAPL8>D_X^=6
VWPO=&6<-@0Bb=9d:A#)8>_0_,A.<7BJ<96=7E9Q[fM6eAaN?ZX=E7,,Rf^9PaCU
F<-e0.LH#25(b,8.Ld]U_?+#bCVe(gJE;D@X,\)())<__>3)6X0-TNW6fT_3Zd,-
gJ0>b)F\UY@dOW>.?NH0^)H)9#KU(,aFNZWKB[M3fRa29YgJRK^B>8^G,V:+#_d#
fZ)6>N?XJL[\<HKSP-QTJ>W<QFb0LB(CJP2H&E5F5fVI[H0.UfT@XX?;F\5?SC^U
EJS@0c-JM#a^1c1/9a=:HHf4^a?5g9)cR7UObZM5\>3aHV<f5VK654>Hf.=CAb9W
GB11W\aOUf)2EVF5]D8#f>];gVO]cLQZa-b(.U+]+MYNg[N;2FS@0)f@U\>#d3V#
b=QVa82aEAEcK:J/(ZH#g,8Tf:PdWWEFU.UO0)TM=_+]1.0Z2ZR/G1J;,d-WVJOU
eDbM]G4@2UQ^LG//;/1>_9D5/Zf4DV]\:1-B)W?Q-91)5X7Kg>5FP0JXB(TJdOBZ
c2G:Pf[;A^eHW2_+D>GJLDB#D+/;&Wa0+R5#(G#QH\<R?R+J/R^Og/>D<;B[,#+W
?:fV_24ddgdc8GH>;cHV]OQ(FCeYBYI+Ugc4@eHO0CGe\#;JI8Q=7W#EbBFZ5\Q\
6^IX^ZFRc]Q)gXE,(6g6dB1Q&6N,^N6,:X?/OA+\0DY3QQQ3&aa(03-gB=#?ABV9
VC9Z1OMU;dF;Le;5<Q=X-[A?EP>/f-<J+OX:I24\\QGHRHS?aKKD?L50bX2C:ecA
OG>LD.HPO9fH(a7L,#=H[(Z]8GFbL(VU.8BF4OKb56R<T@7/f5Pe[GQYf\(cY\A8
Ed[_b=RW^A#/+0I\?Q,4GGTfTH<(45Z(X-Y[B_\b,(3bTFS#Vc5R<eW:_21.^WVO
aJI_-F+71=#(7QU#-J?5YL>]AFKGd7C@Zd[)OX-;KH82cg-e>c3:4EBLGbOK?B\#
b4f0=(<VDXD[Aegeb16Q:8UNgGI52M0LM9S2L2,>&L;ZL)\.V<+X;C[c;Q.JYZGJ
3,=Q[?3_4OSd]T=cc2dV,<XBe\]LN^:LSeaE[>N^3J]6c?5e+;&=)3Ze5=?JJ-M)
]J9fgG\N_9(L0_2bU9?GSd0fTGXK&Yf=,)K_N#cZAJbaACDaV_Y=1:9>-\_<;HG<
_LC3NI#/_M]+S>Z[@fUHSGJJ1Qd(+b,NUHH(-44]C:Z:&&fBUePCHN.UJ#<Sc-L8
_V#LeD@XABfN0fPcZ<##4Q?Lb_G?b]Y#Z9^_c1X<@=6T1G@:MW?((A^caY/;KfMW
AKYe-><T)[MZSR,VI1c,dO3K-1LIgggF_f.P4AL/11^4HCPf_<QD>X7Q@UQ+5gX5
GSEAWW6g_LIDQ1?ZC^/.Z[&MICK^.15EOB/PEC_0G\B\S:G3^KB#4FRFgZ1cUBV\
6aG@UE[90bUV=Ie1/EWZIV>L=@2--6[FNNIY>S9]WI1?fdNd:eERO4XB+;]eK+Y)
UcIA#O_7ZGAGbOF;G?a>G,SV#)ZPP2&>0cLE#Q\_8(,_:#;6[IAP+:?,(1+92ONO
4SaA60E)DD)D1][A<-DI+S.0_7e#0MdN?]O,#=a39C9b/>D,GWQ;TIdN)a6[[Z-4
KPJG/(H^UXf.,aaL6ODJGA&M0_6YdZDG)4/OU+LD4^e523>H9U_IdXf3D=e,_.@B
8RgQcR3P9NQeNBXZ0G_3+_#G(\+HYIS\VS1(QFUETY139E>^-ddP46a6J),\-&W?
FJ)GF2SJ25dFJ@5.E[;UNYU=;YbXb4N63ea]^aSHQEcg3+@M()=:Wbc./CAc<5(X
E<P-f]de/Y]/D]_?OW@0:G_QFaW@.AG&T+B^X2D]#b\R\8B9fF(Tg^gTZXMg_aM6
4eKa<IHH+IKIH+3D0d8<]ME[OW:;Ga:W)HVRLM\R7a6WNV=.A?;(/MG2HBO=A+I3
QO[\+YO_2>?YRUgg_dCWcP>Mba:>XM,T<F=7_PLG59=;]9YD:PcNQM7Q.\5\e^0g
U^&-,aC#aV9YGJ&B4g@;_ReOE79JN1[^/A7BYEYRd)W\a>eG+[?4.ALb=L[?+;bd
VX\=Z<K\ZKZ\VOO90/TN\\F?SCUN-Ra6C],gY(KZ1]F6E3H_K>N+^N:K\f?@YJ,M
+LW#?OFR=7dUVF5AVef,Z?[?VD8a(W3f+3B9-YQW[_HKe3+NE?#IZI9@#>(1-NDM
90L1JJ?\,_.83Q.\?VD+J;65ccb=28R0I[1/bG4LKJ?-S.3g8GB23c]<0Vg=9eCc
V;NQ2bGMDQ#L+4V:c_E@/H#2-4.&7>XR=\KMWgQ/[c/.\##CKdg1Z7d,XR46MNH&
VbVdO_:)c).c+;N4=9(I?J?aC@6GabVc7O-P6W-4XeK?:.=c7Vd&b)EDLSScL_KC
2?BUT)UTJ22BL0R6S3[(2J7Fd\8,dK8EX_ISGL^2X[(WQCgY8L16Q<SgMbHM#5I[
HK:Q-;T2eJZ<g/C4W(aLRFcO4VaTM:X\dZ]YMC=_2M>JP<;403PW)FRba9;D(08:
-+@2J4=H]X>?06LCe>]Od&B4S0_LLT?-)O(TP]?VI#?&S?/3M.A-^FV,F&:H][5S
\U>CI-9TXXA[O1Q07;@^OC3W^HgT48]HRgVa(]HQ:5RdeIJ5+UaJ51.O:QCH]]ae
,QW6ZE;[0KO-Y<;@/[CMNVR:@+SFX3&g:8U+G5AYc-KbLMFMEg4GX32=<^M>TQM_
8/Rc_5_T#aS9\gaS:U,17TGV/,GRH7?/0,()@1MPX5-5A0]cBA,@SM>N]L@aQ,4?
),GS7>Qa,aL#[1TPAgRRW#PIbgg<IJ9+E7;K8bgIN]f&a<bgLfSVZ[SJXe#fIUac
[H\@IaQ4Af=^.U2fPeY6b.N&&#2.=)2g#[_[,]O/B:Q63I->AeO?A[>87VA]3OYT
04;4c3dGX/-TK1=FJM:U.,WDdFbXgP>)9AI[gb66UZaPTT6M).c-:Cd;46P1[UVV
3Y&B]#1X_VE179adHZI#gQA&4eLG&H=8:?5V((.2GJ7T<N(NMF/=HS7@<(]-eU-K
NIBAT?4TI>;./a]IX45H6MAJEa08M&.1ceM\e0K<PR1:_KBgYG3UY.b^[EA.BN[&
87]C&e>_f<BRKdO^>1-&@]]fYLdU0b)XU3VR\?BP<T7P2?1EU/@3Q;MYFg4e[&>U
.LfQ@+)a9SW>M5YRG80)<+,8BTd2/^Sd3]:.J75]3-&N>E^Z17Y;F<aKfJB(DNQV
B8g_FGeJ^W#[c_PXgTK^KC]18W9U/,IT]QbI5M6QX\370,Y1<U4KC>.7eG]5Q5L-
#MD]?H_#P[caG,483CD?,IIN2LJ6^3W27@6/K;6f<<M>IB[Q&X9X;13Gb^I/W&V<
c_=S9LK,Q993P+DERRC^,7Fa0)MAS6(4W1XY03(fI-QGTAT4f,FdaEF7>OOMA__M
DTM#E.FG7W[)3Dc\+KGKLRCZH@G:5PDaE8N9MLKR_-+8I#JG)M&&G.B8\V=K,=8K
]O]Y1>DJ:a<?M-SePSegb4C#5O<SG/K[FTF5WH/>_:XeGEMVb\e9.L-7;L-ZBD#,
KNdTYH@QFf4YZ,J]/\I_1?HCdNA>SD^Q?.C]LdfN^>F:aGQ:PMKVb.O7KZU-:#&K
KRIJQ.d7ZTUecf<E82V^NgS5/9dFA8.;Na581<W+ZV0&X/3e]TQHIUTGIK2[,K<7
C(c5>#J,9KKR+2NL:U@6fZe=P\JA#&g,f4d59<AOE)a;&QN(>_@TNO&ed30T+R8,
8H2R#[[FM8(>>@#Y0D9<Z00O/GY\)?C(#(+\DM,_\47e.eWAHdUXgT,bHPL17gWa
A\&g0VB:c(OKIGe0B_g(JCC0/(FQBD?76.Q6-[&EULFc@[N/O;Q-6]W2PC9[(/L<
&g=#]L+Ae/\;&Q_6;RbUE:N_H.06N<d43<QKMQG3Da95W^E=a;@^YWI4@1:8.Ud2
]<<K,JeP^L=ODS@XU9;)_]g/V)@-AY@[dA/>3CA1E;c=>6f9F#SR[P-D?#&S#U26
(VRQ]M/MY_KWLT^[M,HENVb[XLYZKZ9+B#B-^1.#8Ga#^eRfUA30X)39(CF)OJ/1
1AGC&AUXc7=]:5<,6<RKF/Q4#ICad.,Ef^\7X/MY6(a+T3S,X&:KQTBa;H5g,,1Q
f5HNJ\F/aNf18]ab?ZdC7KM2bIJI#0eH<NO1RW?LAESA?=SaXLJEXBJ+1=6)TJcS
Y\=H>gF?ZDG6888KC9<]S>P7A#>0G]=F3S^=XFC_Q]@B)@WCS,A8C]#O<08YO,4Z
a\eS0E5bA;GFGbU3e;U5gGS.QG^2[D+ZT@-?Wc13DLHfYY[#H+XdPLV??0:9R9c8
g=g4@NQ5O.ZdQ:\e#:SC4L=6>>YcXI&E3XPL5+OT[32ZR2J8J1[BRLWP0Tg9YgTd
>;F@IdVD6XB\aCFG(YC/d=<L2UDM0d]50>N:&^2GcFa(.>D+XXV[e0PLBQF+;OAS
:;/\DEg,aL>^P)0DKL?]eXe/OJeP]\0(7.ZaFN;9YIM?f^1edZZFEC0X8P53eBC[
-c3;JO1KIA/T;RF>7:\:E44QG2.MA>NGK0#/fM4ePT#c.X&I3+#cZP./-U1Ue+AD
d3BObR3/,fW0-fM==\YgT4)\8/E>#b]2C@A>RDW(^9<C.3<\;-FT@HL6&]e,48#e
>c^B+Ggd+JY0SNGRa8O\W/ZgHXTO;.O]g#ca7]955HY;EJLQQ7aGET=a4O-0cA:[
^^ATO8T4=U)f9Q/eRR?O.4:7Q^bcJ,8#L,F]//cJ3>FgafDf>YZB-DC3.3XPgf#5
I;GAXeU>E/d><3\:9.7VLR9Qb4(H_=5?DMK,>7:,66/I0F9MYDaa&bd);&e9c146
^XU=TAgg8<P#DL;-LGACKU5[1XcEY.0I?7;TEg,K8/#//_W-;I7RPZWeY;Pb]UM3
RFIM8Df>.^P2M7FaUYE_9<EDNg_A9;.9[;P.CV0OHS6V753\cDVD3a\A/;RC6\K5
Z^R(&g=D(5C[[aGc<b[-2/^>KS)53=D3<L=:B&CDdST)-NHE_+]+;<<,^Ie\G5U3
5V4UZNJZ_dYb:S_=_gPB-VBc(>=B?cY)5#6<1^0?A>1WNP)N@Y93-^CJ\)Qe4XB:
B#8SF/La,J;1U7c(OOX3&?D;TV,JId1#FT^Ye)AJ^WS.:P4dIBb>7Y5YB.ba-^UG
I2fA&>5Z[0Y?+ba?M)-E=-].gS1X-X9M\Ga@_I?cH)C>>Nd)C,\83HKY,1SCV8e8
b]gM>XH?e5UC7cP0>?5D2KX@C-<]bL/,VS(/X1e^7XL[>[D_DSU-:-:^P::F-f#N
84+cG_2&RUR0<L2HJG32cKK5fb+>GPBDgI3X@-.HPN>RN1425F(76G#D,WDKMQDE
7]_bcMT&Lb1N?K/a#>;(.=M_LVQHR:\MW3V5:(?]-+0823g9067\>?G9Y2M\TJ9@
I79):.a[B^f_YdC:1TJA_SW3-cPE/e0(2b-LD0:Z+P@(ZY5\7;1V7:;7.1G3?DQN
aJ:;.Ib_>+IUE4[M,gYa0aI(^2L#[(-a54<](\1bPf_+<D=CZ7NR^#bV#0g1?S:Z
W;NgKe/W)_#4BZ:&.L^K2d[63/YQ<YBIeAR4_e_7U\JfddU^[aAPN,fW5e:=?86H
7=A=2ZR+GZ&LF048I.?=D-]6IT>&H2\&-cUA_&4TP.2VXP>-e\/C-X]95Bf7JM6c
(K,/.e;=PM7ZX9@#2ag>]@KNJL]RD2]\>#VISQJ2VWWKL&3eNA=c1.H,PgaZ/LG0
CXg[BO&bfSYK/,5K=eJa0Zc,)cO-H2L3:&[-1L^>(Ja<0V>):S34[42??N^79JD7
F+4f+LLF+eR<aV+@dNTM^S\Q3KSJK1[]>fP<#^4:G<MRWKIB]^S1C=&EVCbF9B\D
GS0/7?V;092H04+T[W_5;bgf1E?B8c1W^6EAEb-B^BH6fV9;;2f+^\d55@Yc0KSd
^/5V+QW\_<J;e]^_1eIUZ.9Q.6WNb_Ub\[T680cSMYLS;5(Y0W^1Xf7>;TO2M]/6
1F>YLEg,42YY3cB:;@I]]KL:FT:WLSNGL+<_VO?BW3,bO:bE>:8>QWN)4dC3CHJ;
VQB(IROS=,:I.#;G/bdf72-BH9:7^7:ALS.N378dJZUM:)@H>;aGW=6>F=XE<O48
UJ3\.Q2Mc9&g]WL9aW8YDCd16YY+[/VLVI^90Tf9&QTC4-[F[f7PQ5Sg\HXBdJE-
FGf2=ef]GW>74.)R1ZJJ)fbeY2FRYF[LSI,9B@1N7+:EE2?f:O?);\1Y\;<=3.1?
e=&1bGH51#3PTT.\C?:U&Ma+fff)g\Ka;bLFA_6ZFf]Z(=:K7:ZdbbH?/T<GUV])
^<+0\/Y:)MR29?]^:\22RE0Ua7PI&/ga#SCSD_1RV?UEV^MMX3gg(Sc+ccYYJ7UF
[NCQa;P_#DPfKa3)9M8V>E1^WM+Ka]<S\abKZVdGQY_NNYB#JWWGR<?I#6&=V1,;
GPSD/P_#N@IK=bON,DfaK^09HeM6(AQ2#<-/L\1_T.AUZEL+.]^R0+A]I]eFU7NT
@\HI&C==JbHgb/6Re?-[G>#]OTLHFa:.<HZ.S[:IOdG5e[K+@\)]/H).0&L0dQ:K
&(b)Y#f<W[QYCI666)-,9^HUP((dHN<5.>JV\VCFfG</>7JN&5C]+=?VPGA;(MFa
\-<Y[.9Y.D:VA=DHe,P7KQ)Wg#Q5ac;_><e,0UXTgAB^9;Y<bX>#Zb//_g4VgagZ
SZ461=XC_dXgA;M-ARM_-+gOFR@9XO2^?cc+V:-8)4>OdUWdfY:R=N42BD(FMg:N
,(0FIOMQZ+M=<I?fceX^e]&PP3GE4R<P;=;B6?\F)U;][+-ZJK6Y5+<d2.FRG[CW
+5>J@R9\-GLPC4d;(K6+YIV68EYFKNXFUd5=96Q)7-GOP3J,5G78,gFPZV[XWX35
C1cS?b1Pe1O_gXJ]=47>e_a=Y>59TS3AY..\,HOeg4=G)[Q:VeaUNb[d[26aV\_Y
/aO/YH73K7Q(EY9YNY=&TA+RPcPfE)FV3^5=C&2gZb;UeR:KH>5+JXba#YFB:S5(
dCFdTV=cLb>Xe\PL=]d+5&fb9@]gCJ1(KG4Cb;=B6?PH=DS7^eHee1Y<,gOaW[N+
Odf\-8+AX4X5FROU2fBK8SKGK:Bd,Sd/U/I36[[3?I]P,D5a8M_J+>K<.FW&)#@0
0>5BD>5=-BJ+dQM?6,#J]P:4cHHOPTFU]L.^)A,KbAF.T+[U<.=PG\(@YaJ#OKA@
JA^Y@,4&YdFOgK(=\-0FCeSZ),(-dJ&1S)&4^;XYC5JJXF=7^eIfZVaYC<gV7@P-
9KX0U/7:SVgJK;.M_6gP_)V9+8/O:BW7+,EE<egD8[.g17-e^@0/7g1J\)CB17-T
#NUQ&C-A;8599E3[_3M7d+:5PU61]g0-#I;GGE>C)VAT,D[5)>RL?ASgLNH<BU8,
8O/B:_UeF>U/F07c,43P]+4BHdOWQ5e4:=[&)_]Y:Z0AfBM?@4FU/E8aP8M_D4>.
T\H&Pb8(;fE(8V+)gY_ZE,<;7[^.[#&U(d)Q3M<K^ad\6WD?/E4HVP#W:@[_?/(:
Yc3^<,14e+c@2.c,R-D^FG7DSLVZ=&BIdaBHBCE>[6,3dTJ23J?./_.A/L9SWJ]J
H-+(HgaZf8bZ:Z[ZH?CP);T@T;^fe\CCS9IebGTBS\+R#MFW[PaWQgC<g1d(?gD6
6TB9NLG?#[\d1.954+2J98C^<g,H)L-1]&2W[?6C/b0YDe)ZIR2):aYRaJ.?-4CR
34C7QUHI4O7?+@Y[ZSaA?1EC>4S7;MYN0cZ+VKb2,<2]>3Q;RPc)L^NH?2.)cNfL
91;P&Sd1WBC:1RLf,YP/EgH#4aC+cND8)4Je2T>?_AAV0-Ja>MKV)R;VeQ]2]G2<
PE\e\):bPOg9gU&Q05#I>6_Q-.]S?Bc/\=P5A]VSdD(I>_e59ea=Qd)U&<BOT_(1
S5L:g\,?e#W<Yf^T>8SY91+&f:d&B2D-GM)0GQ;F^/#Y^IBMP@/RJ-/EXFfd9/&A
^7d<)4DI093@(2JB3:QQ^/0J8QFM>@UUH@(]:,N5(=(D;KHcQ3JfA&]^/F8egDRK
g:BC07ZJ7gBJbaB=]Hf5&]0/I7SQWgZ0)e&I(aK@??+&F\H)5RPOQQEB:9:#R;c,
.AICKTT^dX,7#Tb2K2]E[]IIFUU;\NV^1KW8N7-S/Pg0Z924NL2g6Z,,<f499GY:
^[DZ]Kc[Fa56T)9Pa5/Sa@)I/:F+bVaH\Qf2PFPJN&?AN]]=]AZDJR-^_MgDIeFf
e>IYZb0Y.(CI/QE<aP^7<FTK5FA:RJ(W\5c1g<#V<Z-?AV<-;RTWJU=(:.]^)4^S
_E+[C1L5G6[:R&1S0.P68eJ7_JBOL?PH4J.DW?_bRJB\#YPCaX[::aET+&f4SJL.
C[R2,>N/6;X-#_PE^3JCA/70f]:-]=>eI+eH1[IZc@8JNf@9GPgEI@0R@K/>MZYB
]C<gON@)XP;0NLXIa;6DB:d^P9X+-c=DNLQ0(Z_Dd0)4Kb+JcH;UN9_?L7@3dP#K
e:LN,?IES@<-UWcF^,Qa:&L8.T072OMU8+[;(O5&3V=]A#;#A]Z<STXHFf7#Zc<@
0Q9)@7f_PC+BKXTJV?^b)bVJ0;BR2N8(\SF4+68V#e52F.2R\<?(T:bAd#^KdLH=
#HVM)E/a?-@X0,4?->:=ME=]7V,f_-]#2Rf6O7L<FFSPE=RP[FYdMPK(.RLQ(Hg8
TJIGB>@=,8W](6b,(OAfHa/AAQE+5\f>ZQ4WOHH5)E870FM</6CeRMH/,bZ0f^C#
BMcgXd(#Nc61ZT^XfPKY.>.WVB;e_.a<(g0:ZJ:P5?<8)5U^#==2g^NGN]KSR]-;
&HEc^gS;6acBMEL5f-5N,e)=ge[7.RLEea?@#_EQ\4?6[K7YF<8f=fD1H:B<<e<D
CI/)CXMVYSZ]^bOV-1.\-+:(JTCB>RGNPG@/g#P,YX>1\ZQ9OCWBGf)\P274EFE1
>MZf\<[Z4<DU7=99U+V>]HbIP7:O)]Oc:KZ&L^4dT35ZV,Q>Xb:[>Z:N>2e]A,59
g-;L#fa2?Wgb_A^NS,A<P3SI>F>O=WZW36U)=9AN5#U=PHY3S>3aW].]O\GKH4fS
2R]TXJV]WR5&DUC8@V#6SXQb)6E=8(/4Y]I]1]+9KO]O-(d8ZD&L\IA;HW7K3)5/
[P8133YT36=<B5B7KITd#dWI>,f,8RR3OcLbB:1P6>e183@TJC=\e?R99PO:2Yc2
D@c0_cIITN;8(.3U8IFU_+C\e^Eg,X&P#7^@246SG9E0\O;/GU0C&NWRE&<MY8Hb
B8.9I3^La0?6f>L2CdX1)M^\PWB(?TKZ:e4;G+4N#),#<Ug\0;9YEXNL)_4AIF:7
<W)CI/b.Q2_]?f\AOA/P78\8E@a7NBRP==/Y]E2I>@(U+6FGA.(_gfPC.Xcd.8QI
cGg^<XCT^)g+:)HK&7CS6M22@BA8J04&COQF(1,N\MWG4aF67HX:JJgIMX#9d(8-
?d:5=<6bKa-@EFHPPX^8RQ<dCREf+1)ZIR6[I,eJX_VPA54VTKZf6g]7/X-[G.XP
>Ed3G0(--9F<0G4:&CMSeGWQWeJXZ)aJ\6fg_1MA.DWF&E/MHP12SGcIP3W?#g)I
,DU1W0a[c]Bc<e)2IfTIK0V--F8.A/#Q=_Z+]7-bNV-ES34_1/WWPbfag],]F-F?
Cd3_68QB7WIUfYYPcaGVXC.Tc195<+-cEH:#CeU[FQ4d0;FME\.a74&_A/HHA5g1
ZGFXDEPLKAb[S?O=Ae/-S2\7^MHfB42C?C/;WO07.+8>/KTR1b:L2[1JA(AeY292
f1OC9U^2[H)U+;K(L2;1>N91Yb3)J#[a0\PEgET=DNP<.1\.#Z]L\c_#bQ.N:(A.
X-J<;,EaB572;g80[f;ZWaQZR(KAG7T>HY113;Q@QAXQ8U?)00<3f>,-f69^1SRE
),a7W2K?7WB4T1N/U[CP6.BKf]LP47WJ9#6+e[R;JKa<4YLc)<TV=YD(6\@F/(J[
CLDO;fAa8S/1^S3VC0?#7c9g^6FV\AEfc6-AP0[Y\b.#U0^ZGdL^PSX6E_0PRI>O
9H9@G/8@b6IWRT7U@JW=,8(.XA6V]7>dE7K&eVf9H;8=:f4LU,a.7DeK_>\6>XZd
=7_Na-.Hg1<B<a@W7C:V@d\aP(&X,7;XdW4(<\-b;gaGIE1Y:L@>,Z6<]cX,<0ce
T5g/_TW7EE>]Q[-Rc:OI7H9Z11E#HfTL3]Tg=H4]=f7Z-)e/S)DM]DM:db2eJ-Xc
1NRPRW+]2Q:BI?,G_:Vc?L8=#<\I-;Z@XFbFd64c<NEcJ+=^gFaLJKL4e(>VIe9a
TC0-7g(UJM2c\9?F[A]bBV=:(GM8];Pf#+7c])ED@.[fNfe/dDKe.P5gX&f4YC;J
9P\#-88^G.ZNV(?HEVX<BF<=)Y\#/;AN#2_BG+YW^gKA.#a#K-/R)Z-g)UR.T(E:
d0b:GGB;,SGd]N0g]&&F9;S+S;QaF5T/V(,a#EAN)\VW2_CL16\g776=XN</VR?d
;7OA&=f_PaTLg&16TKVdf/6[Z13[,:FFORLU]LL@Y4.eXC^Ac\PV.Y&>S.0RP36R
(9@.NQc:MYRa;2H.RJg]:a@G2U(Q,>B)LFfD/L#7?6_EQUgDYUaV]H-@Y,V1O[.<
3^aDFEeVA(-B89A+FMUU486geURLXNdbeY)g(2OPcE,2Hg4,@adPM?f1KKN-LL>R
]b-FdY.4WIeeK_G8GLC;QU:[=VGT8@dK4[c^T>#+\8gdJ-6N@[T&Vgf+AaV.6ENe
<QdSB^H7aY&N.NWMVS=#/]_<Z.M(NA47bAEZBVDR<aR[>b7((:OR6735^+_<F12X
PeOHbG+adE2(B-/HFc8DaNR72U4d<UgP[TCG2-^9W[E<CSTG7ec^YP>:#BR]E>F&
;LC78]HL5+^PH5)5Z2TZ]L-dEf./N>;H.K&gDO4-+N-eK:K.<A:2OZ(2.B_)]4Y7
L0G8aa1@1f#3Nd5CbT?&12,+bb8Z5>4=c8@.]VZ[ZP)F6N>DQ7?Pg;MT#)WA[]TT
7)8DI)W=Q4Hf=+b1,:Z#I^)0d;@BN@aBd>@4?M@Y[d(C82D/Y=T##A.?d=]=TfQ;
27&Uce+Vg?OeMdeE0R3R]T<R5[J]>;e.Of[3]Wfb6=PYY]R&]53#@]Z4dLX+c17V
Me=<M53S9NDX&Ce]:7@=OS?PV;;J]H7?[3deWZTWF;2e,QHSY-_\),YZWNZ6WF7G
b48g?8<?(X&5AV#2eAQ2Kg=-=6D\0QRUDd>?4Y=b9a[0/U78N_T[<A]:ZEd._a;d
\0AF_M9SLN_+(<gE<B+W)6]&JCBFgG4D^;6O_GMX5/_C(^gaCdJB+]/UVD=MUK2[
.g<[IC515OLF/N1LbZK9K[SU8^FUD52d=T6eF92(/WPP]TTJ6?7@)6]KP.2(NWW&
gLHJG:?M=9J\8ed4d1f_^/<=;>&@OaVbbE3eW)&219.>56LSc]IQJ6=):EfFRJT6
0W=,34+,62TdB;UEc2BS7X3D-S(/YLBAc3JX<]]\P43N;?;B9Jb2VNHS;a+FYIXM
[9PP->7(H?8NePF)8R6,&67R9+HI40FdgETY<<=MGaa:+3PY_\f(ZYX4g=JS)b0F
X3fJ-\2e0A2G:UFZ+/(NKH++-2VO:T^eB#0M3WIAca9:^K.T0;(c4Fga2cH2+H^8
9YKa[QE44BME6]O7aR)9>J;A5:B;f4?F3GU_U3Xg5[-Vf/AO,MNBL6MXPQ(-IO0I
KX4<JSJ/0LYUaGNMLNcQC3V)2e?_59]:#c(UcO5bI/cB=TDd-:aFABX64eM]=ZK(
U1VBNI^.W\87J)7X\@8V#Eg:H7c3XN8V4E=Z:N#X(((0LR=b28G209?\542YDfa#
>9?5G>UgbcQ<L\Z^Y>_790SIgWED44329@(6DE&/X&H<dL5D,Y)T\87d.>JJ92;d
#S2JE.B#)[@[1N;#=-Y2O8Yc^KJ5<c1^EXYU+&#Ff/>.Md173S(2+;SU&MF-X3UV
eHAMN3A9B1T^\Y77O805S=AIM]YVeD.8+dKc(:XQJY;1:]?RAOcT5K/+L744H@L5
NUR7Gb^B7:/^G+2E^N?eKLE(Ra.3;D\F:N_.\)TPH>Oa(La9ZCEN9RL@ZC<KHD:V
Q;^NfXfD(RQI7?Jf+<Xc//QWXLTZ[d(5(GB6_TOY+3H7I0MA9>@bg,5MZAI7.]^A
O7AgW\0B1H8@^WN&3,&d_UAN69,A6N4e(Uf5YCX]_Q98U^#1\))3Y@JJ^c5AFIaf
6&^Q3\8^XZL_LMT(^g)_V))bG0b3&.P\=:9PfMb_VK7:U#<g?);egIaY;YH15<f&
EO9+V\Q6A_?O91QNKR@,\gJ#=<.d7)&9_=XQ&]N56MP=9Xe(\;#<--]YAC0/,J4J
H?dZ_.6,2GB\&@dOGKDBRR,_dG)a<aD/92<IWTIc.6dKHEOf->6/ce0)Y@aS.7bL
#)D<;BQW<dXfK(-=.0OF=4GZD;(YM,RR+Qe:T<YUfDAg?/Ve2c1/F3G3JITX9.e_
&>SJJgFd+WdDJ3SIM#QY<6K]#..XBaG?+@Y[/NYAG0<04Hg.Q+2&=aKQ=\^R0KUC
HJ+&_QF_W]/+c9G5=EJRS;Z3K<0eO4=GO(:UHR9+RPdd0OcGSZKNcS^5L]A#63f-
C6Fdg4)39)L4N1.^+9_5CeDa)GaW,J+;O\ZQ&Lg<>8PCbg.fZ#(aKDTZFcb&&)3(
Sf#5T55cdTJQ)e,Lg8)-3f)4\@L^.7c)G#0ZCCMd?5d_CD5[CACfD\&&/CFJ&O+^
E#VP@YC+XD::g=RaU(9X1@MME?aLF(5D4Og;8)JMbOHcH@bX^6P?a(5M>[W]gK[;
RL<ba_SVXPE\YNR9IG,-C>=)8Z.RJ)aO4=EFCAb6A&ZPB];:6Ifd9AXU?65g\]E9
dc+E(00g63<0fYV;&SBYV&)R1.c#EZGYUKK1cXfR-:dN(6PX7YGF6.aAXB,/VJ?c
6Y_)0ODEaAe9a)0c;NENbDCCY.D)</Z4O1M]VRS28RG,fbbJ\QKW<X3ZcOd91SbX
[gYF&G[e-5)\V&Y8]b7+_219eW8f;C9S:M;(bXgH_&?A8\HIJ\S#Z#.;F(_SPL@T
(008VM.X.K)L\,ATD/VDBEA/R2K.H)(S[Tc:H>+G^V/cMJBWKJe&\,^K\?f<LQAd
8BPIWJI]4f_0PKdBf_gIJ1G63(P^><^2/fY((?1X<D@67PC-1]O1K),O)E@V8LH2
<\10;Ed;IZ42PB.JS;?:B+aPZe+USM0\P2M6)c/M=S+A34U/)>K,^&UAH9UgE,NP
4\PW&a[(B:bId>9BN>7L;?@<9a<1^VaB>QfLDS)#(F6&:)/AZ6P9#.cM3=#6@/bE
RA#U0RZ6L\T_A8.+)J#7J/E27=dP^P]PMTV[9]-B?]3J^Z\][W11;I]C?bMI,fPU
QDfDcP]S\4Z;NU<,#aY?<Z@4XN,DM6PH0Ncf.W_&f>)9S)=Z:cWW\MeDYVDeIZIW
O9b4T2>b23fYR)7GI_/?B8-T?<4g6+RF]2\FbfSC>R84PW#S;c]M],EPZ>9fF\>Z
U74&?^?1T)4gIR:W#E.JXJ3A>EOND0FRf[8U,7B]S(47[Kc&S+)KHLXE2?2K8MD@
>f3-A96#2]CVWHP6WEDaYN]3b9D-CH.fKE:R67,-^N5g_.0NOX7.KV0(\Z3&0>aY
628c3>bfLfE,+\L;6DT2f[^@e[-R\H6PCQP[5]_O61OGUE5PG&&34C:U<8d7FWSd
IYLH^dX?EF;)L5#E3W./VMeY>X-&8Q;Ze\dIZ2bM@-DJVOUf+X^S<V;-I/TCID5+
;Ub\+^O]7T_&gKFG->Z<dWY8LLe;b/[J8U6LEG_,GAC[P9)fW2\bfOJSb4&]2X,R
EM2cc-\&?W>8)#^:WB\MK9Ig/.<)8>)d#AEJ3-C:W-AGB8.4[dHM#[,cY1.BXfO@
]59GDXEW[PY=<;:M>P&S:)@7(8@@:)7Ld7AB6Lb<1FZ\,8P+/AEg>_\8HZ63K15f
4a3O/N,7X\@bL\cY6O&&JUEI877TK^NRCe#)[(2M3bKU;<>P5a?-MTJK>HLYP:&3
6W6.K.<f(3a<5b.-;VR)]&LZ\-H-#+[d<_2JD9,cY/1X:TfGQN,M-eKd4_Z^,\7;
_1?:SL4OC4RY#,_Y1\PIU;H0:6=O)d0+7++Z3W+HNNPN,Y[&(H9g9da[9<NV=B5&
Zd#cP1Fa[H]PFE5:.D73=_LbKW^_:[AESCPI78S3#6I=V/NE:?+U[cSK,>TY=#gP
R)77_E1,A>2PIN-4];91bTYR-#I1LXSCb9WD@6g&WEVfL<:D:aLf71]:;-RTLMB\
S8gPJ#?<EO/1JBI?U<8f^;DQ#A_/EN.N[N1AO2]P;>O-+6(eJ9<^:fce,aJc)D.V
J?JR/)ZBd#]bNa4?0d5FdXe]IV8Ee0C]W.4DXURFX#)378B,K/OXILTbO7NU5.3e
9?^c:g,Q^\2(?IR9eDLB<GY>bI/I#7()T,#\J6G96#/<V;+K.BO.Id:I6L^T=@.)
44V>-0191?I?6YF)eKVf7]>-LD6RbUVGcbH+;+Q\K[97JQA.c5F3<?P:;ZaL5b_S
Z<UGKD)4b7WC502=V<K_dXO4Sb:Nc^2eAHb&Z/6\?g8^;_3:HT1=VP^#@[bX4dU[
>Z47T>2>e[2UBaNgH<P0+>+S18>P<Ya;&THDF1.8X>?#0Q85ca4aRCB;?,.&)cPJ
)a&@I[\DZWYHNZ2@/R]JaO3=?B/)cI:BN/J6e<4P(G9J]TT)11&UD@=eIETdYLge
^6/1bQ76SWEXT]V:g]R=U]ZK<<a#IG,>[#RQ^Ff3J=^A>7a+d41<ZC<\^?<b>23K
e-9E;^SM(aXDWZZBMGYa;AX?,-_1WeQKN3VG2K=0S#5+MLMGD<3MgXX9^&QXP^O2
?0J@[FY8.0X:M<C)R?4I>9:3T:GR#S\4\FWfc-IX=O_OdV7KT3H\@;<[S14_:A_e
31b[MB2ge+[[XbP0JQ2Z2UW/b@_Z;KTDXFD1P4ZM[I3BCQDUY.OXd6L=EN/21EB]
NeIQegS1:QLTL&8We?aKTQC#69&3UUE<X<6#O)V-3:<>O><d]\-&RMF&K?1;4=/(
gV<-7FQCc)Cc:a[Oa_9W==3bT2[g,L,]8QG?#0YU2M#SDHCG3>GRYgd/^KB_OBD+
/FSEY/&Z_R\8eM/V?gTc7eK/AU?AD/?Qe/P-\-b]QM&KQbS3VV.[Q2=/decgDF#/
L-#V^bK(JJW;JOT]&\W@^B\]>X.5/Qe]T<98B+QU?PYXecKK?<,,WP-:@<\DS]KZ
Zf?5Z4</:1T<=E9P=7)=U)=Hf(_(:035,QB12J/&S;MNSO84JN7G/R+6,M8,.K[@
YI]gBCa&G,W,>]PJeV1OE?M^U-HcEWL.KdH8+/EW>X/WJ<PM3?V;E>+SPH[EVW<,
;[]@a[G4J,33?]\X[:4g<WLD[6D.KA[,T(A3FH9(+?T.dFUZI0b?Je;IJ,^U0SYc
<+U:+MZOT4Wa,g5L_BJSF@aU8ON-2^V8c<D5I?^EdT5&W?)LFA-\/ZI_,SLJ<d6U
fe?GNKRa&B^Gb<&?DaR?;4B2=_2>A4W83_8@O?8b:b.FX4SXeFLHFHZRaCC279f<
Gb>T4E@1:)/GENSUF,[KI1?(O5f8INGHTW0?W.;g-Q/@_918gDON8gbJHfPDWT-R
J1Cb,8GDVL54.f-Lb2f2FNB^.a#HaY_2,B/J6U6MR05=ZQaU-EB7/WfKCZ+<YBLd
IQ3=RZccU=OM#BNKW_=D0fcbf/5CAcQXG5HVA:>fb8dWZ9d,<FVAYV)5W2HW7G@e
3S6Q9FU\f=#:\e#+=4CcMaG[12<06J][,=DeEgLI#Wc.N0A#g;0<1?5>6]XLJH+O
,IgQY^g2<2Fb2(^a(^&=6BDFQ?&M\Na5YNF0#ZPE]@V/TT6Le#P;)e^Kaf:+Y>Z&
IFG55]F;34afVX=..5ZOR]=#(D9T6e#dfAg[c8URfDY;D&KPN4+#EEc<G49(NLdJ
4XJFK?.PK1E.]-Cb+[Kc#//&OFVO+OBMFJ]cIFEc#13Z9aS<<<?a_ea]7E6B=Xb]
OG=P87Q_^4D1)4I4fBf>5D5N#)L7&a.E<L82+TK^TL0+A2@a\J5X7SF6;JSeA-/6
-B4U+)]Z7O)NQU/L?Y.JWA(#]19UZ/.,TGEJ+Q=G<]2RdM-CT/>Vb]dScVS[gg:Q
0gO9T=WBY+\dY<H?>-0E/JTF4INZ3(@MFbA\b.b7a)C]-)S9^O:/.@g]9=#YE,16
W5J3c<8I6UE7K&:\GVUeN4YdK=f+.Q[)F0K]GL44cI(8fSe9=4H:;UXd(FY]DCb^
dHDf0AJDK@648EJ4Gc;\GWT-0?/2J+O#//bD9V<daJ6Vg<e2)UQWB<93I4QB&3_9
aD4_(5G6.+NF7(GadJd6de6U1NDA9,&NTYT(3fT7KLAYUO\9(V09D>V(g=0PM-QQ
b-Wa#GN=73VT5L:CD;e]MeA,Ke[,K#e@fF_K:e1Q0F5#Qd5X(SE]RN1]S:<Z]RQ=
/X=3F+gT&<Ke-4L6X_6Z1.P/JD(1E[\d]9(#+6QYW_VcVZ4:1X7WB5?50M(cDfR8
R5(:dK[S^Ve]_+-3K2Z7TVB__H#.6da.cQBRTBSWJJ\[KP=OM#;;Y\b6L2ZCDX^U
S4cbaR:;[/IR2c/g63Fe6Mc^XV_geT6&2,G,,2?Q7NHE(PO&AEMa_NHH1PcI.g7>
.8Q\>^:Z5V6gfAB=EH>AA,J/X(cVSAI9&#fM/E7C7Z4/IL2\8#U(N@JcbFITd+.<
TNZO-I]0PgcKT<XT7I@YdA+3V8)3cM60T)5?SNDde+3E0gY8599>5N3Tb9(]Mf@>
-_>_e9_SWK+_Y5NV,4Q&[,Q0QgO0;03C7H:8dBbAM#ZO(WU:6HV-<9E,:L_=F73#
/[cM-K-3GQ60:d/#+&SXg8W9W(Tg7]X;MLb/6[abK[V?/LEWA8C;9g+G>-HK,?XE
9N+e54ZLT^g^2J[3/=1-3]4IK-0U-FQC5I:L9#5Q[VJ8^+;H58H2@XSCN[WHSQM-
^&V:cf.T;0>H1@.VNL,.>HfDgLV.d+NYgV[I_Zd=1<\c,=KHBb6UYcfLeW5DL(&U
Se,dQfgNg(/WY8^FcI]f2E1AbTg7-R]V_BYGTJ,@/JQ90E81&L,LFQ-JZ(Qc(agc
95g]AC6IbBIRV[&RH2FY7#KY8H-V9c2)4TJ\S>A6aIOZc/J3ORFf07Q.L-dNgANc
EQXBLKEOTQ).)8W(MP^=86)a75fRQ0K[9L]PY@X.0cc1(WT,;0Q:OgCdF^J8ag3Z
#E[#cfN:XG^XJ]SM<]5.3>9Z#d+MTE:d52TEFY?562XYJJ.,Sae#L(2<Q7O,./fU
Q[XO@;d-HT+Z1^N,@JJ&SN:\3[2L/I#A/@cO1.-Zf#e[EE,QQ9_(-YHIZ4d5Z//g
;22(VOPaPeWZ&3P]:f3e+;64<Tf]8=T_@@6:&+]eLYWd1)8Cd^O3#^-cO&Jc&gDX
4Z3O5][H7H@71\L[8HTB@SMQX=[7d[13-fIgc)bFXH1-<L/D_ZQ^d[3ggX,Y9H1)
N_Yd_M/X&AH3TX/G_-bWQY2Ed_:1HWgH=9d6S[TB+?_C8A)>(d\<V/3>_BSM66AU
3\8B<N.[P5EB:A?_-BL^P#WIA^NJ+26=b0668bS10LS[PQ.3)K6,8f/:3XC1b=E#
8UOUb@HVH1f26aLAK&B5W3RS0;^6I)K(:.eCB@aKZ;__\-:B^/,8S)#9g3<8444D
eC>@:.cc6#L7PfVL7CV7bPQgeQZVOb,248U-7DIEOCRFUCGCI7Y#NSA\#V=IC=Z_
<[A=D\]g<?T;@VM(01\-8(,T>8,2)M5@b>P)F=gDPAI8=QRSG^&X?UO:_@0,+b,Z
5K&@>(\>+I#C;++8cT/09:?6N^ETf^&LKbZ][X9RYV;23eXM3LE[gXS<4,c8D)<G
2RFD/8(,TN/+-8Z<Lb1HRbA8ZQKY(MB9+CDP&DJFIKO^5cC6_.bf/ZK,?\?OdIG8
&,2f-O-#+ZW]I-6b&VWK=3./(8M8VV/WRKeKS##F2/Ga@Ba76I1@:FW@ZMH/7E((
T#]9)N1(:+C-0&^745)?G,A@K47FAK)&aVG#[C.=AYLU2f;U5MA?_>TfdNASAEEP
OM65gR8]>.+\>MN3CXE>[->@fA>=UER]9QIB;M.SDHU2OFMX_4.W1P6,OURXg2\e
^9#K:#UEA,f^U&E/10Z(<W^S7eI^DT]R@^3,A_CA=M&X.#RF(MW:YY&5[We#.MU6
IVR^aKJ:I2a8UB92Bc<#2?E_;5bc&]HB4<^fI#FcJ<d?>L0)3.NXPS:e=GX3&P5;
F#Y8]N#4+L8-L12H-=4VBEHT:<L@6fFRIPV).1B:,g):M56BaI+Ed98V[E1fI@0U
WT,.4X4^4A[IK^>#6ZV_>MFY-X9<XbP-<X^PR<25e1WEI+X.4SOKd._&(TP5cg:Z
U88ULaa841>2RDU,W.c=B[]KTK/(5PA0_#KB3MPUI0#gZgKcAFI>-FIY;_\;=V,+
4J,:egFabR653K8EQAGUHGQM\+3;#TT8=a?W-L<HT]Q6#O25Q?<H<T&4bP_b_1e<
D+XAbU3B2#H1@1[L=,WE7d0:XSA8^DJO4C6AYB.2bCX;&LY2.;a9^;83eU/B:d)?
76f?\WPF9g3&WDM)#7YNUWDd=RS\+a48U>;D6U;7^DY6A9TQ(=#4/>].C:S9E/R0
;0^Y#LA;2+2JW/_2D9eS;0c5_FM1@OF<JD3?P5[N>Qe3@3[N0MWH^PUOd^H,C]3A
-R@<d7._2<&_\ZB9J2L[M&IXc7X#4KeQf?0V(/?8_Qf11.CBZ894\HBfG?\@;f@J
H[.C_Jc<6PU@SE_MCU#HSEHHH.EO[b?(Ja?S&0@5<YK4(YeMB1(gUSQ<.3E7AgLT
M4KPcS0f:IM3ffJb(&WNcGaYM,4?>I;R>BNgYO_AR:<V\/G>Pg<@aBfb)+9GD._d
+^\._IPb?&98[IGC:[/S_?_a1U#:]Oe(YA/Y#cTNa,B<F4a82]I>J<RHCI<CWB:-
9(_V2(^VY/#X5?:bOOTfOKD.FF\a[IT^+)=GN-NBSCVOF9]/;Q,P)J-e,E(+X_5K
8SA-WTF0C7c^N@:H8DDZDG\_X[C6PJVC4<UIKe:2_>M+@BX4eBR(JIg1OFF?C=\d
;c)aP),8XbfKF;_@O<AGd3^O;Ne;Mabc/OG7Vc:BFN>)3DZPb(C&R,63_d0D)B<8
2@?=+eDcd<LCe02#(8Tg6RH:(A>,e&D?-@Y7@<+@R)R(<MEcP7a2]UX37N>HXQ\2
9SKEQGW>.[?JD7]00]/V.b@[@HKZUI;@&U<aT00A?;VY[R8W)9;,=W><)Wd#TLRB
XQUaDcSCa?,\;V@;/#O7B,ZAHMTf6P0cGHc[J30&9DM9+2Q5KeE+Q]]6#aKS:FYN
I0f1VX#&CJUW)AdbV#e-BDYP5=L8T3<]PC.aV1VfB+.C,;bYc59XbOGR3bTf:7R0
=RI[6]W0JTF(^.ZEPX0D5/U&4+dKWMba<D06T-MaU[J?bfb4SLFFeZD2/KTU:86Z
12U_KM@LYKaae0/Gd402gcSK?E@[T#g=b[4.5#0&QZ9[=(:a;VJ[8W.84=A#LYGd
M[RN)3OX<@?4ZC+3\g=JBe4-;IL=1R1d)TBWW^<U@;G16@TeJ-\#CfeWWNTT@X(b
H07C<@Z)7Y7fANDdY@FDF&8>WPWNXc<P78I+c26#)7I<7R16cV_OGFLFG.APe\RE
@T&=bgG[_\].BXB#R19\R8_99Q)C9MFXa;,OQ27,.d.1]V97b#:Kd6J^I0;#M7PW
00=4P1Y\P6WgQ=UA/>1^&3E_>U?aVV<K.MW5@g=ObPY1W39/P]f?be?=_dV9T08D
MX47.DE:M9K:@g1IIJ/XL8/2M)?/bIeKUD?bGM[c.>Kd&MP8Y5e\EQW;Mc95,U77
f<e7NQ.M=QE6KdX)P#PSG85MU0J94VM>Z6X=?MSFc#GeW#_+/LXTA1YUd3>Q;VbY
RUT8W:=<.=@@5?+[?[?22)SEWMfY+BgL6S3:56D<Ud,?I1(QZ+ac1:d.+D?W>09B
Mf17V27[9@C0e_Q@OZW^fM;/FHUHY79)fA.S>aSNgINJ=gP1\S-V)7=+Q)5[X9[N
>3M\IPV?HdT@HMT3Ree.U+2718fRBO>K-SJcRB3,WC#(67VH(?LH//[4N_<Z4OJ8
eRETB9g.(A/E\M2[OAgOe<)P.>03/#Y_D\8G>@N7AM31,WgGSg7BP8[F;08EL+,c
2+:f;=&3031f?;fA41gbfL:d]-:@6>:OJ@-PG46R;HJb@ZT?[[JS;c?f^0OG4WcT
K7+eGSVIBH___4_1e^9Pe=DV/@?6BS>I&TO]-E-]C+2X,)E6B,Edc].VZQO4^3T+
f89LXC4G[fI1;D6B,0W\.P#VVL\&G4a-ZY#FQTY[JAG02f:YBW1<<1g4178#76IO
+N2B1#d.CBIfWY0HHBST1\S:Xge85M0I.=+<CZ=+#c-O>\.,H:SZ4R^O0]XNJ&,S
.OdHDG,(A-gM[ZdTb=(JO37TXDW#UF2aB)NPY9=Td:Y&\-eN?A4JN)<AM48VTbUW
2S@IZA]LE&e1S\VE\QPP08X2=aZaV6gA?2U^Ff/W2-b^M+W:]W_)Vf.V5DS(JGC,
<8NE+7TgaeY)LcBIJ8?/d\cNf/bV@MT2)W8-QWSMdO[?4IL2WZ-G+,VEZG@f[PJG
YQ=+45##CZ@B<,]RJ&@]K<@]RZB)bZ[9dD]]>RP3M7?]3,B-P,[^K\NI7D_d[QVL
Z+M8[LW1)N4dJA:>VUI+O^cNRKdPGNDM7@NRA/N0)N5JZXGc=/5CdCV@@e9Y?.G,
<_;3#5(7g]gT>#>HC/;+gg(#=/b6]M].B<(ZSAM2a6&ET[Y81<0d79BJXV^MR5GE
(C\2Pc@7Q:KXH<<_-7MFRM#W[V9L?/+)Z+G&33C:@#R((U4N.:V/5SYe+bW>9AS#
E0[#6MM_DT;?-eOOV[D9LfBUIH.&.N9@E(A)WGf=R=c[(+[/fWR.aa+L4aP4TG-e
HZPG4CYVbK<=MVMD_GT=4KCJAFJLd1:YX_,D>GX_BS/fUUKGdVUOgC/@OS7,HfV=
AgeOCG)gcCC1_<G69;U\TL/-U09)e@0?MSD]?^6T:Me]#-Z@I\?Z])JNbb><7Qfe
Q@G2H]OA@@U3c:EB#U6#M2#Y4d@ER#dHMRD9H-Ud0e_-T.V>6\EEA^-KRc@^,d[9
C[,EVA(c8@#D/\]AQ:f,6WALC++^KQ:,(.(10.c/e6b-]FY-]Q_K8S[O85IJ1Aeg
#=IG>6?aB_DV;_>fUN6=d7N;-YM^/:aWEeUQV#JP3J1M>;D0-ZW;d-M?712@?9]F
\f>I_02YUSPg57b9[;],_0#GR#F,K4^4](eO303D6JP<d4c:D,4,HDDf^J&XT.)G
<KJYd(a5(^0T#g4Q[IP[b5_IMBIbBaQf>?>.N.F(XA8\<,-&TRZ)=T:)70[_XTW+
2DGSF;dU7UJ35X166B-Jf:7U@@E0YcI9;:_=];KRP:_=bbM:We>S/PZ#PfHA3_&W
>,RdE0E,DF@g19Mf1S0#I7@STEY^bDV6DI6+]3TM=5&4L@YIB&A^GME4=g/7:=#B
@f<5EaH3&UZad#SBHI=bCQE6,PBXS/?DV@3?;eQOZ:,;V;-;\cJ@aP-&>b?e/7&E
GPOgF&51KRZ4KN)g-?UL0dY8KT#-]C2[7CGS4MZEO,VgJ-eJCQ<Q50)?TOIHPEHa
4-AMe,X0_49SGS4+X;SF37>+/\UL\?AAX6=</9G(3T;/2/3+:FKLK)R,#C\RQP4^
0#]A3:]KL4@&NCJ6OEPfgUIF?<4^A)LM3<IR0]KefSA=07C3f+;?ed.D4e+7>/1H
M1OaXS@NS1-;6\,WYR7+<CbE=6OQ>gID+0ZAVLM:N7M<.2Z)EPP4E?>NS,M^]N,=
Gg?5V##E8T(+F@,G,I<fFE<Rg/R@0X-L8]0YU[T[LM_J79-V1gFPSNIG68b#\G^R
:K>_8@7DX?K+.EN4OB@[ebBHdN==E=_)XS[<\#4gVb:;U2J1]DXgDgEeS6Ic[21e
H^cRB@FPE>J;QSU43VIaR\#,)4T?Le+)0N^UI?KdJ&NC-H+_O.M([L5=)6a@9G^X
4+:5eJ3-5]:1e&#_KD2OTc1[aIdf[E;84_.FKN.J=\I]Y);8K_3#N3IM@g2f-?L[
>N5OT/7Jg49eF;G_(TF]8?LgaVU-N_aTe[ZR:W-L_]OUM6#(Q4ZYAM/)CQ0U45_G
,f,=0ZPY^\#>:FD38d&e--Ma6Lb)ZgB(UTe=#Sb&Z<P2+Se4AK;fJM3f#gIY(N7R
N(78,LC@N:VQ6aQ0>SHZCPEO&6@OAePY7S8MCUdZ#Od6@/P[TcRPT9<(Q;4;3U9/
_gd&ZUN4./+]ZB2g\SDZ-A0SfM\535UY<d_XIA&Bg#&IY,\O5af(.T1K(Ha<VX&.
,#1?:VaB+7NaLJR\6_^MC73\DEW8+1]21da4C)QB-X\HT&H<#@34TL:E/>a;@19R
N&_1G4&[_\7[M[TdGWR785B;4BI86,W,_<dW/Vc&2-O_&/=H]O^D&c\.UCD=2==L
[5@D=[+I_=GS7TYFX42X4GF&Vb-GW1V#Md\<a+c7O2aA4F_+JDHZeCA=(X_3g?-H
/b]@ZYagO=bBT]&Z#U(6eXP7=H^M#JK?MJD:H7[R0EU+bI\(=0<_B^g96.GDd+OA
KP?TU1X:DDd:H]9g.)\>W4\gD_X>].HY_##C8cL3f7MFP#,RRd#:.H25QQ^c=+3A
d+c3dOdgQF>&SW8J9aD7ag/X3.=WD<3B^)6)]:.VWMEX,6>Sc^24ZTL=&N(:GB91
3ASg1ZTI^@)2D,L++W6XO6gJ+.J;A/GTVZ720?0<=IF6NBa6b\^H)R^>Ue/+A;P-
VNG1WS26ed4&+_((QG6H9/0GE9g:E-1e61=<\Mbd.A_0b^Q^ZbDA[f;;Df;R/:Y9
&3d7c6R@K:2=5gQ:O+Vb9FM>#.-e2N,,R<7)NU8[cE<9+Q@eag]O?<T[>]Ac7f66
,OQHdGa1/8U10_P41=<UBd^PC6[D1f#\I>PEA9]7MX?\I/;Y=:6;X]VZC9Z[=OT=
=,e>N7>VPA+XR=;E-)ScGJ=]-V8)PeOZ#[IT.@4@&61BH(BID3464QH9;&[B5+b\
0VUM3/?JY&OFF/\C9++g7&XXJg9#^ROIAb^@5C6VRbHVZ]ZS3I[UNXI8H&3B?.C5
fM5O&]KYOLJZSGQeb/dQaO-eM/&gCN^(;&02:Z_ALOcf;/[b_;=BKS(;(1>(U/W_
FJR-/]CR\VI7632[?L=F1&H6+F?^6JZ85;.0[.W?F]HaA@3HJ.&SS\I0)VHf-:+1
SAb#L7c0PPCB3,,)-.;E.OM<.X^G,G&4b.<V30WfbD&5?J((aLa2cUZd>eb<+22I
ODbSDe[98Y<;c^>f)T4ITNACL2J&)6aG?9\\+INa:V)S>;XF9C_-^C;b<L5Q)HV(
OSb:dT9VLMBUUcG,R>,?\JXZ;^<91N?e7]FA\L[YA-0G1Za7E3AfRd@bU:+\POaf
FJ:WQb<<S5Z:D>@0L(@b,PO7L<SS3aO8GQd#e<T9MSO7GW00E8f679aPRSCRMA02
B\5c9I1PfJH+.@@>QKQ4CYH<L:(U9D.[W>U[_N,egg-JD(<-d01VYf>IU81M-)Q-
Q[KB\_(a1QS+_MF@f81_c0(0OGPY=,PM05\8#8O2BS\9A_]K2A9DG_=^+9PR>(.;
5[2?fLe,;D&[33[<C\b[<@P>_;8cJL.SBPfaSb1#1MXe&fCfTEggd(B.gP\KSDYc
Q.?:g?TV7Id[g5,-J>K^2UUbZKA?Qg_]ba\gF@B)->fOdUNSL0+5]V^2TLG;>EXe
G09LEX@)7>g[@:#M0R.D;G[JDTgJaI>5>55d87A&>Q([_:XL]^g<NcB7c5#Uc)c9
eN1Qc)bc6d.c0GCF\^dF1:=K15_;H;/YgLcH#47=W;c)I.5AcUZ0J5aE&A;E=MGG
NF5L<d;@SH:;L^1LU<I@-D84:;<dN@<OP[=G+?FcSf<+d8,QX_&W-&>cK/9Pg@(f
TVK12(;eA=BZC:=#:^Eec4J>#FR)+<S-G[;Cg<N=.(?3#))#G82gPZ\,/GK&3J,7
3VZc/9M)2&S1]8C&JO:3,=TQ6?_V]cM\0@8C6;]-\RD+._MP3Xd8SS]]#JI6PS/_
F4Z9WPaZR4A?+U/\g#T\]Id[Gd1;^2_dUDNZJ:&(Q(TY+bZ48<2Y4eOZ5KW4KXa&
(NaO[KH93&Ua_6D0NA61/]2MM7]F47EaU]R\Zb(\=H1f#0c0BDA^ZUM)J5e&#QW\
beNL(]WVSWXG8VA\gK^WbA-(SM#fT+O4D;W@a-Fc8,9g@]W657O4fE,9f,AX(2J/
U3<RL=5AZ97XBIDWKW2->T0NX7)9YXA&a2ZGGK.X4TRO[;>SR2\KJ=APZ0WC9QD#
/]MHYE)#<gHJKY1Rb,FO=\>++0+Z:g.BP^8YK97W<4C29Md3D2JU1B=O4>0LEF_,
()U\LGgWJQJ3?Tgf3?GgU-]Y5QH>;;B42<&0[\.(VUZ8M:Ad>SSK,YC:b@ZI2L0A
4(XdZ<JfR/Z+23NQVH+=+EB.VN:X9Q^L&.g^ZJ-<f:b__X-T&KgAe1.eG45LM,&(
+R@6H1A:(E>W#)\JU@,R:/gU#2-RHU;<6AF^fY@41+OMeWec3PF1F,/1Sc)Y@F9]
Y9/dH]R7/0_Sg:U@ZaEaW^YVQE7H0&?[EL8<ZbPV/1Tb_6[G:L?8T:>0G_K(?@ef
0:R>(G,Y&.</V06_L9cN([SD?4+7<bYO[Z[[<+NR.1dbR3+3XTQXaEa>#:R4.V6O
QD1L0,)9;?^X+=c58]G7-.KdA5f:RWG)S4\-@A\K=)I7XA]8U>Q[.eL#M.0:L=B^
SG^M)4d_Tf>KG2P0\IAgf&?[SP[?6S3.Y[cX)+[+JQG1d,-_J/)NUd/?QQOXa9T^
Ic(IPS#g&9?DXP_D483O7b_2L6EEI/<#WKgUEES>4VLd0@<<\D)[XQAD[.PBLf4)
S>&EBN#c<,SJ]bG)+LDKB4;T0FZLL[UQ=.\dZ-0.5].A^V=Y=I=W/Og=]a2^67OS
28DP&Z29&[I,RK:FJd.b\4A6=,WR7R8OdLP1BP3;d4D>aI[0&Za\:/#57,#cXAW5
4]H<PJXAHcf>fTMP2A[9@\;KD=ZQ3B?#ad83)F6)#J3IC4CYUaI@>>YL=^9T+9<[
V9X)_X#@B:P_\GXZ<V)AaJ08:N.>91:;+.d<1JDGR.1U@-cdO>XGB;GbRH\N;;DP
aMCLZdAE3(<:YA15=fXKMUO,#;)??=gN5WeQ9-Bf;:(A)10A7^<E//&FREX=QTMU
K[OD4:U-0A@BdZZ98T[HB\a-=gbLYV/:d2d79OUX#[<]ZNJF0aM]QB)Qf6;Q0Ae@
caLgJK4-ecZ.TYF9XYH6T^ZFQf:YS1/gK]^2Q?a((_WSA:b7E7A1TM1=9GFO5K5E
_2)aKXC0>.e>IZ&P/Z.a4<P?Je9GHT8MIE9R#LI+Z<)3&\ZL0MLNJPBVTCKBFHOa
/#O&YM,dKY[dPD,d5:/42NM;5KLJ,e_,755;X5#0;cSMB.bI-fAAf<^S@)K8IMDF
f6VJ#NKeLA>c?7EC&?;YCAH^[EBdIeR^\I2?:-=^@F0?9VV#_fc6R33XN3G.W#Tf
\:F<2EQ[9a,EU9Q.#Ca4K(;+cRXAJ2O5J(=ef8S^@b8XaRC<Q2P@\c/g[.\6G8(K
?YU.G4Z]aR(4EVeKH^NA=a<V90\/+0(,U@&c\(c0+^EC.](<FVIAQ>NfQ2^g;&#:
A4=^Gc5S00BH\X.\=D[UBPe3?9MAI@fJ=F\:XW^VD;H<R\3^V0(bFTD^eTYbC6R=
IN:F())[Rg?:(7dcf2Y#X=(.C95Mc:(#)2EbB6D6&/&AU91DHAeb-O[aZO=1c;dd
6YDTZ582U_)D[IFMf9:TID]]PCNI=E=B:<RHUQ=GB7UP+#K0f[aN6^K\8]<#JOME
NdB<6(bW7@I164X<H027[K=PBgGEGM0:PHb4A[Y-KI9X(9VCAI_Ug)ZfA&AJZRJU
LY8_)5#g]a1A:eR0L#6d?d4OXZ+FV/aCL_^\E1[bPZ[]eB/V2B\ULC7OJ[B8_+K#
\AabAD@<0bdJ?Cb0M0H>b<[\/)A]dC4NSfeX)16Ke0:TL>V6)@H7YB6QN=A4HQW-
c=/0?MGdH#:UVY)MW()&+ULM/R;fT\3IY.Tf4-.\FE:g4Y;869R]eSUg&#dJ4PH_
F]NSI@B,S9,0^/.gP)e#a]edO\&^II4E/)H9UQ=\:C,+JKbdd1Y2?AE0UVYDA^,Y
#63:U/L0V&U#M\d.O2&##JK9d(_45DD7CS[QfR/D@T;8#=#a,6U)=@ZEQW;(G.<=
=JN:.b+e<VN&SUZXM-DcB7?UB9+ZDI^8^,==J<SS/U4>45UH#/1AUK^K.-RTJ&T;
L.J8>OWBGU-?BYNP[\?IHLgV;.6E9Z^b_7DU(485J4GH3OPdaYF#C?Fc@N6--?K\
\G\-a-DFa:6g:8FU8NH;58ED<DKG9&IL/CE0TD,PN?FUKZ4L:7)-eVNT=B,>)M@Q
[dZ;:^[NTJPDUdXHV@W:^5B[CR1DL?D09&^4c7TD91P\A/cA3S#/5J^Vb3T>MU,I
IEE]B1_c<1GOA,M_(K+0_Y/44Te46SWJ[>N77_--5<a-HU>0N=)KJ&0MLC5;3@^J
E^A?HB)+W@XF5G-g?^Lb.9Qd+>d](YE/fU8D7b.aF[g?_.SQf3X5af0AZ&Z[[;(S
JM&_dO5>Sb=Y7J8#1KU)BMP[R(DJM]8gKI;8c#/)<^W3;<JP]Y[\HXJ\(T6^SFYN
CfK:??DcQKF&X7WYQ1.M?7NWO?Y^;N,P]8aVO>8G1]]^;PV6\GffdWaCZ=bNB6F;
#BOKLbYJK\M-#P>57HeIgb=(fN,WZ&MX,L[X=J[FYCP8ac.=I(\X>V1ba_c)3O/J
]&=>JF6>@f[KcVA^_H_N_TCT1b.2),Pegc,HI>O(B^aBR38S?<^30@4-Df&CW==f
D75Sbg-RJ,WfYR4TC_RKVM/6\_f)TXA17?;3[+BGHg1.:33Wb<](95CC1@^^+30a
_S1TMJ>O&bb<d0;/LW=d;4BMW5:[JH/Pf+&B2:2Tf<>PC/b;]X9^OTOTVXdBHY8J
\-;fGCHXfXeS;^9.dY=E?g=XTE[T5O+JB?aXBa+;C2\(BIM],+N&H<e6>Y6G[-DG
AaReZf?+HS7M6CdD[)=(?P)>YW#7HNQefT:)X6cFP9fH0:VA+bXfeN4NFUPY<a?4
IE<M9fF+FfM.>8dbSgg:Zg&+.H6^f,I;X:-g0dAERQYN)8_&^U0IU2/7.^1L4g0?
Z.Je2>1?#G5/(DQPRS6BO]RA)TKYI5@\Q.ObV\H7;5VgT(4KNWg^Vf&=7N^@g.]P
:.<^Ab,a1^L?X[Z]c8.@N[PE?MgfUe/KP^G/XIA+CDFdQAD=3G?G_E9GB/L(a17?
=5W80Kd(V@aZI_b=T53(&1>VafL<bcB:gJ0QIH-PBJ;9/;HgN1a^J3Na7[FLYcW(
_BKeHD)bHLN1gJb,\DAH4-<a\N[a2U#Q9fH8T->Ra#^D9M0QS4CUEGRR?2+[/#,E
Z2+J>]8cCJWG;KYP[^eGBD5AP7dg7[L2H5e,S_-c]b^CD,[T.Bd88?)[9:+T@0a&
faO7BOX&;_QSS]C1Kg&2Q2J?L8EFYY\+#D25W(3V)eVXEI@/9#/GA_8==5_Yf@CE
d8N[JM[008JP8@17gdNET/QRLfbMff.HHJ<B,YVS_V;KaH7?T&B,Y-DRE-8,D9[T
FK48(1BX_8\G?KB659U@5GOJNP+9<)_0?_9CK,(H&PZg@52CDM-UJJed.20#HD?8
:_RZ]6aL[)A9a37c\93QUdQGGKa_7F_Y_37JTM=fEH1J^6e;U&A(F&P802R/<F26
F)SUAgE+7Xa]DfbUMM-J2B6dW3A)CA:ac@@OJCPQSB7ZHHBW_>;R\XI?MCb0HBL\
<+T=]FcJ)R>(Bg(6UfW;<7X[.4P-fA([L_)7&AR>ALKPU<&;T0eBIK;;]:SKbVa]
#CRU9MeW,d4Y):Q)8YHCP(,H./6F7FZUJ1PaX_(Bg@[LdCabY:8?ZeL+E.PPaNWW
LRSb1DFIa1SU3/:#6W=]A&cWL5BEP\R#LR_+H]@^<\:Y^3Tc#\?PS(FJ:-Q/FH]I
8Z?JST5=K1MT-ML30;a;Y>fND5Z-7CZ]8HKX47JFMO@5]@CYTY&KCc]0P64\Dbc\
CTGA^fgM+X:K6dI4JbP4PU)cPaH#56fO0</9?KO;+K;GW);FLQ6+c1Z>_?aY8,^X
MT#/2VS5[K&QPOVC>T2Z:5F_f&HJdF(NfVK7;H,P;YW5MB:#Q@8YQ&(,gN>d0@@F
7bKcM&OVP;EU;M1+<K[JK[PY<Q1d)\f3)KgC#)K1,@Jf2?0.HR,&bQ9gO/M:BX\7
.E-CZ[HGa;D\0(^SG]-H/FYJ>ONRALTZTO#X0[+TINTE#]R.)GfKa5=Zb6Ib86&g
FF<\2HVXMMHP_1-Q8U[EU@6?-379)gA@WXPR^U/X8fdY2>LBe#CaOb3d_]^aBC8T
@4(9RPI-Xc(e/C3e1?bYZ\FdcdcJe?/];-\1\83E[,@OUY(DIXU+g;7W0F9aV6Ca
g<//D>a/FNF@6/&:MT>&ZXE,#KF_c>U>IaD\ENBL&80/0^-W)Q4\0_bfdO:O<V2d
,ET2L[R#P@6Z_^&N4JG9+c9F:UT-CfFX+<a4-e/R9L4UAT\SMC40:F&T^7I(ad6F
KN:=6FWJN1D4VZ<8[)dAOdbJ_SH,Ta2M]X;U?:^W7cDbEUZ^7XY2C\V2#D)c;2D2
&9W#CWdUJVKOK;</Q=KaQ3V>?cfcWUaQ8:f/,^YAP<\BECdERQVU;fI6eO&=,D@8
_8QGN:?R#OaEa8>c=UeNWF<J.Z5Q6#La]WVU</(0I>[XB-N[0,@&ZM;Ee]=8b)3Z
/f1c-9[]RJ15@HE3<2QX6ZccU@D]HJA56L9OE]g-Z+M<BTcZU2AR\.O>fg0c@dL:
JM1/b9T1cO_&G.\_SVg.5:<0=RED41(]?QPGH0b;b7GY\)a,#.BMHb;)b9EAaI7d
MSaPDYA@&fJe3F64G^8)N0ZFJ?_WI5d_aga-XM1c5N4AH@7gSF0Q)XeVAJUXZZcB
SMK#V,I,;:OW3CW6>]c,#BE61Y7g6TW9\1:1(XTDWEaE0G(e&1e:2==I+0,4MV?b
e\N/bOUW?:agU^b7+B]LR2+&/K=a04818I5Y991AgM.02d&=G7Z2=J@AUggf;43[
cWIO-gE4FDNBT-?]AWP55H0LHA922^[&SSOUgfD,1D\Y<eBceUCP>IL\^ZBZe.Fe
T]M^[&S&VUHH^&6B;aY-dOB?:LTEUZ[IJB,[R(.^YBf&e;BDdJYPB<BdNJ1g]-KP
]L_GF/&0-C?_U.=2O)ac4[6=3>4X^WR=HM@X2fK6E;+g[<^1J>_b.Sb4,KSS[QJQ
NB\78ML-9H5Z4_7EB#dbg4DC>VM/(GfABEbV8:4?]QFB^NMB8UT2-29>MK.B1TQB
[A,_=?6LDgdG;Y<>eZ]]=?JX<DBgVN)(Ke-?5DFaKCC?>R,\7=_2QK5H9ef3c:))
X4XWe:cK62Z5G06?[Z[7^Z@#R,bB[73g6TZ>IJV-^]:_V3C;@gb/Y,:gV[SL?@W1
Fg.Adaa/@?71RD4BW6SLbU2Y>=g4Z,SS8_T^2,Z<WGb@Ma6d5_-3YU3T#_;7Y8=C
[CZ?V\U3X^M_I-BC<D&9_9Q<),g69=[d,Z1#(&NgA6\VU8PYJ/_+_9<?WO,?d^_N
HQH.NA)N>1O6[f\(UY_EFP:E0\(edVD6LZSSKQZ_K;]#,JUc\Q;FgNb-T6#EP2)G
8BSCK3AS+3b_OU)U:(,4B5F(D/PXNdPVWEKL3X/#O9NE5f=\+5a;FbZGd(YQF[);
@#(\FSa->D_^=FcdXd/PLOR_gXLS&-RAUB3?E\H;RbQ]_OaF17LTReH3F61KN5CH
._&Ka#J9F[0)47^&EZ/]]K>7Q/B1B&9b3d600,_J8.ST;ca2a&:KW6[Oe9a:\Q=8
RPSU1=^N=@cJ&fDT<aB_Ua^\_;-5\]e03>a,@_AS;cIH+>5O\V;<R;Z,>JE-/E>D
Ta_YQSd49d@aZQAVZ2eFDN5M5(08(.W0X3EG_g35@+:b.Yc02eScZE#ff<P<T#5S
B^eSS.dNdg_UUFDKA;B37CNR#\CNG9FX7-AUF=eLd;]XT]dT7#@J?G9,8\KH7]HD
P#OCfR@0G7.3.J?0eB#;L1:<V&[J.(.,^W)M_>G=7e)81Y4Ld0:0&/3HDCJcVfWL
U.)ATVaU/e/V(9K.TX+,cSZ12KL8P8QOD[Ig.4#D^6af<?a#P[bKM@7+a2:Hf6:;
YBHWELdP5?bN>AR;J?^d_YHd>aC=fMG>3AbbIa1E##H2g(A)5PODV?D6#?L_cN3a
>aUT0QBVNP:+f)45I10fD(Z8b2e14F#/??@4Od/(N6E=EYLST7HZ0=\261Ne_)F[
Ag^NA_Xg[)bU2Y+#2OeBEQ7NFeH4657[N0:P8#Z>J;LK+2Sd_,RQV5ABa8VJFbOQ
3H/NVZ?d3?7c_?IK>>-K:Q[D57FZ>-M].Y_gcS7;b1=>R0[EeOFfe&bA>^LPdH6Z
7_O3,;92@UFSL#_]<R(<dfNU5SZ#AS@WT0P+VE.ADGaeRQgH-Ie>8L>H1^Ve:XX)
a&fD(0QY;?DDLg3)@bIST62-KE]^)We&W;FYQaH0JE,<^E:MQHV31[2,b&9UC\:K
<;4[6L@?.:caAGIae1decK[I1f<G8_/(V9JI(18\5)(LLgY]^M4@d<8b9bb?\Jfc
VD[1[H8BUV@;,)=W71.]?60+DLdY(+4JKHJ,)<_gYEb3]L#Kdf=^I&-@UeJ\BX8C
SW==QcH--1X5Q/HdWB.V@7;Xa1U;G\75[8cU-R3WH:=L(_/D,P7Q1AA-UdD<4WM&
6?635?O+9&a,MQT@L)g9(SMCAR#Ff-YYF.a?7aQ-.V)K^P#<&PGW[//S#AU5N_[T
TR4DPeUZT\1\61<dZfb6&L#T.@3O1P1O_6K2G39Na;?EeURYV.?fefCe?[:8#DW-
f)HC:=c-&=4JPa\eS&#<g29.@)88\GG?M3#cW3Z&NbagI/c>R?&A<;cECWW:8+>f
5HJIB1X0CI:a):H8E9N[gBY4I;K];WgV^Bcf#649FQ+a,.Vf]^?#8ZMPWc(ecS/^
^:?RU9[,[K/^&4(<VcW5/?4>-?11:QTb5^F]O1\3JUGC6N3.:c_)93Q[Ka?FLY;0
-ZbVM+2MgVRg(T_&2:C&&\#THPBZcKXYT-4\6a@+C/H<J->BV3_578Y^Ef4a9eO-
aT^^&)g)Jc#&AXUaM,NW1YEPBW/bBP&aD7,:@-Sc+_TeAe3aRKSC=3c=+>?3fA#B
P9&aDB;]K=9\S,P>V,^Y4@-VGcPEENH.WOg54\,5b/D@SVH<fY<3g2=7LX]K9>-(
6UWAP/+[N\9=[)/M9/D+a<Xf(HbRI_9.;JFMN2E,B3V9I^HfLQE0Ng;_a#SLGBa6
?^XQ6Y<VaQX2Ie8B/1RFBAg?ZUX(3MU5GZ_D2Ne^d7c2FE/g)1#dNd.=.\>\R^bA
7Z2g@ZZMW,#4T(6@5U@-+I(&IGQbggFW;C299X)9E_b,F&bJR@]O0[830DVc^bL)
TD,CL8dg?OCNV9G]6]/TJ)^+6V=ag6@O^;QT3daSI&U+4BL/NU>(<Lf0S.eNO@72
+01>0JS1T^=TfQ(_Q:3gEeTI8>V6)WKMBSU^cK_&Ce_;)D<ZU/P@&AHL>La<gfI:
>ZP\/VY1K]/c4Hd.\1#@g-^=Pa-J3FT5J9bcaO1^adJe-V?aC6fQI2.A-CUP]4\&
?RF]UbXg@G5L@Fb[]1a2#SQN)VNY3OHN=W)ZJOaGg3LJ#RJ3P>H/U1RSO5>a\:gc
+VA@52(Xd+5bLFHSET_@/LQ8.H6MMK9&@+XQ&.;9>^SDTfDY&HN.1EPb+KVGZ7cd
:7d5(,GR=@#IZU]<F8LZR2U.B:\=f^^9W=-A<748-ZBf89#MIcR></;Y]?<@0>HQ
QeE_eN[Kd;fN(BUcQYIg7V&MZC)&^I&W0UX6LEI3O\NWE]gN)3BQR.[]ZTW-_X8e
96J6V+?;SUR/fLH;9>G?&R]SL_@c<W)#]Bd8W[XSRLcg[DV+@NJ;ZNZC>41NK@90
>K1&U0]G]:8JG9Te13M+Q+;LW4:A1X4_g9Y7@V9@Sc?50d_E2?aa\R;gPa[aSXK+
8MXC#?MY8dfWRdA,4-FVF)L/7UR-6WYC6QPH1/[>R2XPSMJd2LJML2feDA(,I2BZ
g5_U_5G+ED:MF.2+O(F?cW+b8XRA00Qfe@GeXBX39fC20TC-Y92gL8995M3;PC65
IJ@\S+bVfc7e^K_TGB[&/@)2_PEHeOJ2ffNe8BFZ>B@C[.2ZX,L4bCO=M]QX>(3g
bg2^cYaeD7aJ014VU;O,1X4ZZCN-M4WRO7GWUH(X&VBFFCbL-R)O[KE\EEWK493U
J/.CUb=G;Z7+TJHKAeVTPdbRTa2H84DA6H3,6+be994S.NR8d)6\BS5@8;;gHgAB
YXFA@[(d7cEW^5\V_(QSIAQ>?dLbE6g[RZ-89/Y1BMW#&d@M0RXS9=[^GL3f7?>R
c^#L(LWTA<.OM0&ZF26C:Q,a-2,aV5M3\V]>+RFP[V6OaMZ;YfW4Z7?\KY=U0^(]
^0GO7STGDPWH[>3>PM-;]#3\-VN1DL(0+=(@XJ)Q@;QKdZB@SBFF.FT[VTIQ=Zca
>JKa1S8O33:>ZPcBV1UEX7]4BQHQ-Y>GRM-#eL<);C[0d46d:,SHA4f/6C]S2&b\
5=^d]:4FK#aObJ7K1^SRe?e4CRFUMc#/d\BK#>LZU#H?AHea>D@>3(:\VVd7)\R1
PRe_18\LSb?L4#],V_DN\&/^Y@/^^PKL=<<5LAX0(:^#R@?+58c@ZA:AB:FXTdKg
0LMEI\5DcLeRC5a[/.&F]M9Nb,T.625.KH<?HE6Y#gYgS)ag[L+LH#L]9[VRe&;(
93KUDEX)2d_/40Xb+M?_EfY1:UCa3fb]1R&fdJ&@II_a=I?.DgVf7ab3?)Wc-C7;
X62cB]LT^^R.D#+DE-EFYYR+PJ_YX#UdY(DT3X]Y=);4N=F<#[(Y-,)PM_1KLUc(
-J0&RX#6HO&,LW_a0c7LQfSW:KG&aLe3Ca35U#V(]?g1_9/e83c)HT:.AC?A\)04
\7)>7ZP06W>[faI[=HbO8ebVN8/f2d\-DY<L;4;c&](;96U/ZG-+3?551S@XMf]e
,9V5.N:GTFb@>-K45#aOI1[2QR[G@-K,=&Kg\YSZ918/0,X8SN=8WLf.V_1SGZa;
[^]SU8CgKN.B28:,/3VCb0\HLUK>gM#3>U--^./H0G#-a(]-R#EX3_PAN<f\=^0X
JA#e,GP0f>dMV6RVAE2GTeHVR2E(N46W.O.AYAOc,K5D@-U?_SGa5d[X+=[B,#,&
)&#H8>\V8<d/:4;)^fP)XAGN8>&A.91a_e;,6dXZWd^I_8<-DXPM1^6+L[EDg(f5
eae^&/LAJC4//2J;bM_1NTc8NgS<T&RV-_(M]eQgVEa>7-Je<.XIMP_<\GBc+;K5
bR#-Xb[E;GG)>;2Z[HT2W^>?2<MG;2(9ga;?]4Z8b6CD&Ib&Y-Y2RZ3IZ+U^O&.9
^PJTP9[R27X)D]>^B^f-M9PYITa]Ze7N_/GTV@RH4-E8/a0J06P=ZM,M_US9F(,O
Y<L0Z&[A1VZN+?@>T-U]#ce^Tb@I+X0TZ-O_)g_1TPU3dND9C:(L+@P>e#W>J>6&
/FWCH5^2BS&^A1/XbB>7(CJ<LW8C]]UgZ;[TZTTEHRL8TRQ5>;)^DJ\S9+E97CF+
Z&a+S32#^Bc9?Db\.WGO@B<C?).fa:B[E2O7PK06:X;QdW414P;D3&(\8C.9-U8T
#5B\E>OI/C#XG1=F-E^6ga.Vgb3GP(DLd^YgRB^EGR,UJ1(Q?8Y6;:P4P:1T-O]I
^Td\?ZV[4cFO7R_E[_Y6H+JJIbA+1L).D)d#c]7O\[E7Cg@OLK6ZA@CXe\3:.4V?
VG?ZT9-]R.)\EE>\OW2)GY7T-N/;:J\,:0LCc-A+8?&4JdB-7,KMN6=RE;b\L:00
+7;M?)(3_+#RaWN\FcT.1&9LE-Q?5PPf@O?0Qg#aNVF:S5;:df3(8(Q#K(7a4SY@
_PRB4-U4>He:K=QC424H_BN#12a7Q[a#3;>B5Z=\f(-)Cbe\TC:>+bd_<TIB):2J
R6UBR)H_JA\^A?VeE-:@e+f=>NRQ>;4e=8[WdBC1O/VfE0CA:HF:&@V=>@OA,C/g
82PP_,W9U>IbTK0@QG:R^LeQY+T[W2]e[@-[928AB+b2UfHT@g(9&EZN;&RR5:==
O[)(<IH#X.d]HDa5Hb5dg9QaXf=^V4-+#.J^6ZO=X?Q:Z63B0#+3gE6X9b.UM/E;
76<V-GGYB.IZ>A->K,R.(JE-771D+^^.]Z,=(4L8-JC@E\(1FeD,?LVd1aOBDE3+
)0GP4IZDA32<==)eAH3eMbV8+]&C2[_ETB+ZeZ^9@JR]S;663IWXQG@5DCPW=FQ>
.f)7@+8,,X[_PIS&B\MX81Z\ac]G-3NAELQ35gZ5c,@7)b<32>]JWM0?635eE;@g
.da&\U:@>OBS#Lg^AD7fe@Y4c&(7D_+0&H78@_J1KZ0RR1,Y.Qg;I<GfCe[#a2HV
6g@QWRZUS1gJJ]Zf6_-CTL2HVWI,?<P4[AgRDe(/feMF3L10<dEg>K0X+(.U<4?^
Y_fYAKK5P/RFI.F09,[C[-#(]Qg?XL,?Y&YR5g-?Zg#P-#XTN#CHfXYVg7O9^/ce
8BY\cfRc=OEfL2g,Q-d)6SLTO=H1P9R_bC-L&YOSY2]J3?I5dcFadc^.Qc&YT_U.
O<fT:<#OEI).Xb/cVT3+eb\B.@O[4.CC(bU+Id__8CS_<7^L0Tdgda_:F7_73f[.
5)7.U5\[g9a.5&MNcU/ZgV/B;6^41V^,[R6ef)CAZ8>,;.2J@dA5P7dCYX/\IeSV
\X&#9>W#HR&DXc(Kbd=:-(dQfE9dU,.ZYQ;3LLB&I8QaRD\YIR7+RVgZ.Q(\R3a?
PLd]b9C\eMI-AS7Y[8.bP0@S_HJC:+O1;GIfU>XTLaQ3K<AKMQHJ=7c=7BV@&(<]
ZM(XE-0MSI/+[\<N>L0GQ0M>8[.)9YDMg)I?U0TW.Vd@;4KR(_ae2P<_fR\4g5MK
8A&EORddZdRF(cFY[2&+68-Q]&VTa3Q-FCTV29^Q(e:02+9\I8/P>]:4>F/9OH:>
Qf+97>NRf:_6:cKY<@N(K?#7bF;Q_a)R.1\4#b9#[f4>dEL<P\;/)+U(IG5c2FTf
KUS:5_@<S=HF1:H[(g=8+R+e<CQAW8=V6CZE2@9>P5@\=+D]e=?^Wc0F,;]4[^+H
M9g,>#(HJF12/VReaRMa,:7Zb#;RJANM4H.Z2;1(5O^=9)bO5SCWfQB44;5OI.]P
QGZ1KaAS[SCGHdB)#H4>]S7BWbfM=/^6I,4F18I\89(6;a(>25@9]8_?D+gCB?DI
PQE>9\\3M#<Z5,UOVa0J-UD]9:=IY&.(M\P-()C6b/47JK74G.BJ;+M)CM<G<])P
A@BFJ-\)Y(#Of;K]RX]#<fLXT[G.@>CC6_2F0VgADf@V]S2dB9e<#]VTD[gB_aO6
WA?,ga:&RO(7[T[\4^CR[CYcY=@LVX.KHR3dC88L^3g+LRIFbfd5cfPN.79H2@<I
5M?L)Y0(B47:UMS/O7b0HBAN\JZQ(963MSB_^/AO.W=(11g5g]JFT#eGE+J>4K\E
8#N(3/>J6ZRU:Bc,P/KNU7L+Xde&RL47g:&/<&&DFd4LVcf7:B5<4gSF^bfZe-A<
S/#N-OfW4D_<Q-c@]9C#@TRQ.dF//NNZf:)Z5gIX6H5V(O^Z,VWV^7R@7,S^?_:=
?Pc?<SC<^1b1==^),^C-8W/08>@FMYW_0YH&AMa&3R=>OJI<e]0a&,[-+HZE8LX#
b@&6?JSN]UMKA]]D#I#0:CZNVGGQ@-&<g=bQ/\CC,..D-#,J+7WIJCfCEP1VLffR
UX@?bOg><e6@^)X]D.^a/(LI[CR2C(E&]P1SX^EF\L\I,fI>\V@+]#OKDV0\-bbe
f^WVU_a4Zag@a6RC;OX\0UbUY2PD^3S&a((?I;g@JN-1:3XV?XGQdCS8/FL^I[)c
<FHZK=Db-E1_a5LV#dF<3[39<0Q;DWR)PdL]H;]]((UcE,IA5dL]1b[F^3O8&fY?
8O3D^,/P([0bf#N4.4)E<Eb+?eDPU+EBD1fJ\ZC#[H+_L#6N@_?CL(IY;GPQf3[(
?IgO.WBDW?ID+D[b41>Y^dO:X\7__=N@A,/f(77e7+N;B1OPc2JRdD(Of_SWC8;R
C>NB;&K^[8a#@(8&VD<g8N4D1G/[Tg[#1;A;+fc#L)cY\\OPCYRI=1:f;4G-7C^?
YZ(2:+Mg[#fa7AASOTd(#Nd3fX&7GS6K-H+6@J7KM=HfKe/cEg0YNG6HJQ?H-b+/
Q(HVcbO6M8NdMAT-3#]QA8SDa&;W)-&=P(K7:G8XDI_Q)MDF<O05U:@8Q1+c:2R^
:CX+N)UI(I4cbUKbB^=P[1@,4&--L-)PMfD7-AC)ee8Y0#c#,_dX5][(R?,Ob;<b
17OF[c0M=,/&F.JF\+9GQePd<53C@8;@1QcWS1NO/AHf?AaI(eR64L\PJD[-(H9:
T1:6AF_>a0&E80-7@cHR@07K&AdYC:)dOO5&XOcI17<(I^-b/.^8P;c2]g26aQX/
I@\45KG+INPE^e&56S@)f43UgMc5KQY)aX&S9SeaMCe?Z1C&6cX@BJa2_CbT7S-E
9Oa]9LCV2D7#Yb+]P.2BLG.fZ5R.9<eD_(K9^[U6&BaC,W&3E8cYG3aY2Le:=[g#
WNL&BL)\Uc<=9Vb<0,;=fSZCZUc/_DR#5Afg<H+=DSJGXO/OFEE<;H>>]^JSZIK,
BP2JecMDFEJ^G6?F-5Y=JT,+T?)U^dZ9Q3<6f3,[V_IOT(31JfYPfFR7-E>ge(b7
S>;L?F&C,L;:UX&-^&gI\>:IUc+P&B_<M?+P[KeAb3RZe:BLBa4]7Y8a6cfO1XWK
EAM.7ND:E5?A_1^Rd=R>9a@W:JLf&U\^PU-DdZa-XMJ=L:dE[P_.MWQW_/6cLLT6
8R<e/7-;#4[?C8E0+;>cQ#[5NPaINAGTK+Pg,9LaOU&Q^=-XDH9_[[)B4R,>N)?g
I;)W=9[APcC]F&WOI(YBL?CMdadK0:#0cR3[K(R+Z?Y>I58a7eFU>PT8R_8[P^_3
6^[aCDW[TQT-H]QbFGLT7f1I<c+1>NRKM@df=F9+E0PDC5DZ>D9^1Ned^C<E,=&E
&2a?D>ME1?d0K.,O-,@FD;RZAMCFCJ,LA1S5/H>15W/::[[_8VDf]^S198?KN:[d
e(O2_0OG[12U(F8eE7&Ag3.R9L]G:(N<AZdA^:c.KH0\M+UY-<dJ3KE8JKJAA/b4
If3dbUC(BHU<Cc>Sd5#3UZ^.2EXE.#7#(FE5^cB6=MMK_GX]c8C.5)+[3JLO=<#.
&:[E^Q<3FT)<@(US-g9<&>A70X\[G7V>1[>>VQ&WOJT&H#M]e>B#BP?TaQ.1A]/]
g^M;I+Q7N,2e:/&0D>ec<4@fY]KWbGZWT7CSFM81C[;;7cD9JNH(^A[V?@D[I<#2
PGL-4NY)?6N@4S^S:b^]3Q,[g[N^VL(+f/0TgXB5+Pa:NWV86DF7TG/L>EfXIIAH
.Wb-#C:XM+QK5D8AM=JW(4P2bG;bD^ePa>9^;Dcf[Y(]Ngd>R^;;_dV^ADB,dA(E
ALAV+3RPfU+bgda[-8BH:7=Oa@cIO?2Ve?0d<gB^aT--=@=YLWec<D/M2W5:];58
_Mf;1MX\@dRb8-2<ETD;-e?VTCN1aWe3&?::XeUT\M(6J\ZR(IVfNdYTY#0Ye+D7
H7;0LVTD_-T6^C:Q.A9#L\\aK;MCW\@9^>d4VO;/>T<=CIJVgW:OdBV9dY(.8G5e
)X/d/E6?gW+._K8LPHeL=(ARGaFaE786P\d11gU]ZFL)5)3#<aKL88>QKJ1.O?,A
D5S-M?Sa>FbG[XM4cJ<?QRX\9<HDVg0@2;Y2-b\>35#6QA_WR)UKgR.\KK,^N)2^
/?cE?XU/OIHbJ&4#A/f2abb4M2.LH4Z^a6YOTKE39dd27WN<#-8:U+=DBB68b^/X
a[6NTOa.STU>b^KAbZg)dX/H]7fOR7b:)C8JX:0L&;N2Q^,c3Z\e=S)5LK/TUCfK
6IR;B;_PY>+\T>4AJF7&=-U#=MAIS3N@V<+MX;JBdJ7Y<)NA0ND<O&R^f03C]H,4
8JV@&gAP:+4RT26RF@4B(;>]<1fB2VJdJU/cPKI@?XR486O.&Y)bUE#=A:DGddf5
R;K4B\AH2B^DVQJaG.YQN762]IB[JACW36ATD[^<d+]aDTY(M,7.D2^B]#085QO&
\/T#]<1OVT/?HWD-/BJO0L?IXS5F[)<-]+a\V\<YH@]XbLU#/7GCdH&HdZ0AZLbf
e^MP:X]Q(NKCPB;F)8dV>=^HF1)9??&c]\2eG2/((eV@A&XdAEL/80-@ge+c_XO)
S3I?@/7#Hc#4CHL:R#-KD(B\L?Le(=IL<M\[+ZJc^-YO,B)[SNE#X1QG)LcY(gSP
[OF+P\7T,,3b2FH=F#17+^/)X.(NeQb^@Qf;.LN2bY;[0dOP</[aG<Y2_+RID))\
1=2f8TbY?V#f3X+9#?\87G_^-fII#E@d9)#dK1W]8\G07K0P_(B/1]T5:#(+U]c,
_^@8]fc/]9_;b7Yacd)S-6WP=fA3(1>G0CPB5R+F:^)LK.g^gT2<B4==NOBWR)2H
QTaUM0(G@^:Z9GZ4GGW>E.^=;9^XcaA4O/G<KXV>?ceR#f3,\4.We^cD79\a^EeE
G4N)I8X?f]-)21_GQ[g7()\;.f/G]c_fE)7>F<CS&8.PV,<R9Q\d(LLMC?F[_TYG
192W<C^>/EYQ+SZ^+OSKc-1F;d4H#OINEP+1=?8JI?IG;0BZ3[[KBIE^Gb1&\EKB
:EN[KLNMJ3?K4)F6KOB5BGF<;?0?<EY:b,Sa9PC@QB>HSI]SRHB=ZJfQ>g8(<6X;
YdHMd:YO/^(RaFOeURd=Z0O96[4B,bU+eGU1:KJ@9+\WeFY96E[K9bMf;@U4#Bbg
KM1Af8H#9BPU:K7S:=9)+?Q3OQFO&/2dSceE8GC>?1VJ.g:8M(W0T88I?N5PM30d
5-bUV):Bd7MY#9(LR)6/O-^5O/+,GU:_>^:b_d4Xd+U]NJ&:/aN2-MHGR8TM(&fC
bR9CcJ2OH;)b4V>&MQXW8&\3PgONJ.#Z^NJ#@=L0G=+>2JZHLFY[7A&fUJ<_bJ:f
Ne(9RLcVZ/&KL]NBg>K?b#DV@FWM.F/bQIgEALAUABfMe8,]P?9H#-KLH>;G@939
^Ee1Q7[FYcW<7JM#DBdfCa>C(^/g39NB8X\?</>:JYC>3(d9f#9GOg8_M<8a.I9V
0/^&Z9P-29_N,#:;a96@L6K+^XePS^e@PS?Y^T9I14fKCV=ED+R+5R\P)O/\_OaX
_YJVCK#WKWBP3FJ6)Q[6AVQRY<RC[1^;N\@(=PWM@Q(N2=fW)K8f\b?E[d?-RUMC
)Oe/SY\5#67GNC#W<[a/dL?UF87-4H@3X=R-8]ac5R@If^]\I#>V\H&U9E9@QMO6
SFBALT6fED(UMVROWFc8ZLV#X.b/+W_a>\6,@T;(.NPW(W@L]TY;X<\6KR(8V@dM
/\+:V==3(U(<D/+b#<Y#S?E6IY+T]>,PZW@4KE)PFMdFX[&5f1TO)S(PSX[A(2Ic
]K+R:(M3\=2E+a>.B;HS2L_TE^)J)f\)7P5]fEfAA&J+J)@DZ.L/KOP2M#XLdc3N
(F<+^P?:&f&D6:LfE:bEWb>\3.<:SU5,\O/J6->L,O)/;4c13MgC?dDPEZfP&6Z,
Ze]<HP;?7K-(f@5Z+Q1C7EZcK](<6&8:0Qb1C&[NDT1KN\0_8HXSg.]PDf\CEdf@
G.c78bdSK?XEXIY_JO259:C^a7TGJ2TE(/Ic(1[Qbe?6Ja:BE/(g(OEG60UI7W/4
K((F):dX;V^DOLJGf/LT?_8HQ08YfDWZ96.Ab&QW]N;5Z8+07..>AAVT]^92eb\9
UPf3[&TJ)7\SV,9Z6MIPC:)T&?E+[N[I.PG\GX5F>.X)6.WU:8;7IU_U?HJAZ09V
BGAEZC>KBU8@UKFfUJ_O&.T6aeS90TaI(LT@Q#;@QG_L-?dUH.JI(a/Rf[5#0@Ae
f33X-;O@,[:.U<AOU<[bDF4OaTI0;FK,M^7?SW52B&QMFc]5d+c[Y;e4.33gL,.7
9QL1:,ZEL9\;Q?.VQ9c(:I0A/_U-bA<@P[4ZHJ4=>V>5_+3g)8PZOB3]Q>[A<9RH
Gf&+P9(YJ?A6:-3C.9X42<@6X1KIY4dQK/8X)F^+)dB_/YKQ:GH.GG\DZH8/I4YP
(Ig@XQ-<ZWQ/S@[S0Q[?7;g4S_9Fgf7.S#Fc:Z\DEXZ@^#KEA9B\_2:U;;D:C^7Q
;\a/;XM\_]/S1Y0I<(e<T=6U1aIG#0bCD<)71;aND3VULM@[aT=:G9C9ODLMREeG
:^&)bRH\1F0Y+WMK1TA>[WCI6gNBHc67&OX9Z0/SaXdVO26cM69&.gc(GWC.]WWK
QLE>JeDX_2ACJb+URI8F2G/T]f(aSZ+:)b,\309^Q.>U4^\R2X+De>&Dc,b=V5fd
,<:g4VOV?@4aW:74fd?feLPHY92YH7S&b\5V)dY.Q@O0,e<CfH\7C4^AHNf-E&PI
cY_[[W1AX\97S=KRJR-Z&)GW0/J2NJGF&1O3;f\W,=c&JRbOFdRTgQdR;YbKMHVe
3SFcfd_8\R+NV7cdUY0?#(M[?fgJdc(65DU?Y<P+LUJYbYG5&SA]S@cR5I[[9PCB
AIbTdXQgZ,c8@R+Nf21[IVX]gMT5,S@D.\0aS51HHE=,7^Qcg0#7UBS&0=PJ<5GZ
\bA5)c?bL.#=<E3+N-]RE[^IQG<8\]-fd4(Yc4B1cTOE(fR5Q?eBga/XQKOO-?_^
?f-g)1AHG]6RWR-bd>.aIa.aRPJ^EN-19f/GX.Zb4YI:0e1RN&Gd(F#GU&DN3f&V
6N,4_T_X:JfFJCfR2W3VIaX^M\M9XU8RE\N+b8]b1U)e:2c_)7@POHfU&-<YT_=c
HE^3WRcMDgSIgb[RZ71OX_McM?IW5b66?8Ab[WV0^>1<6.>+&?bNY_K/=RHb5YY_
VaWV=EUBN<0KQF>MV@(^F7X4[;U)8L,I>9--:9]GJJ528YG[(f,Y0bI6e\d?b7(?
J-88YHWO##FXFFG#)0)9B-=@0@>-G1J/01[9;IOZS>)/@N(0bRbNFK;f:eF_X;(1
=:[.(9eOOM6D]8FZ7>Ze)1U)&1_?(-b=>+INVa)4L&:8_YD)Y]L(MbUXcUE\5-F:
MUdHS4RURa+JTF1&>1BRb@_SZ:JgYXI5D8^fGB3=b)>_&XF>e#JZ5c?g^P,D5+;T
?U28:@,.JM:/MF2XJ^BS@EZ:I+\gJ/I(#MG=7dRaR5+SJ4UO0L8(R=?XEUa6.^4W
E78)<c@6gAN309-4G[JSS,E28fB;c8c,Z3PD)8R2&24K1RZKWI=C9V4aV2NL4:3e
#[aK=WFJT&;H9Q@,T\Lf#)\BFOJUWSYN)e9K)#^<OU7IU38^L7=f@2S,]^c[,EZH
[LK(#]PESU/(TGBP.:?_ZgXXJN,+K\G[=_>V2Tc=@6+=:VdG8[e#[C:E:I1[H_PH
\JXE;)&6Z_;Rd0RJ6,9RQ[Re4>bJ1)bXZ5JcCZ4e3;bYLZ/)D:=^D.);OT?\BgTY
b_\aF-7;R5PM<\+\#(3,@OV:]WLHF<fQg9]fXC0a3PAM#2MZd&4JUO;4+5IbUg;?
O2+g;@d9.[IJ2ce@:Q.5<c(2M,;E./V;5G;:M:@U+FA)bERO<@TdS5,\752Od/^F
f\;>XfJ;9[U>)+HbZE]&W:JLA52//Y5g?a4@N4#=)JN5d/J8ZP@0@Fe+C=+N:[3/
/Od9[D;P,IcO81X.5^I1^VK#[&[4+S3cNC;<PTE7MI)EcVCe,B^VSQ];4-U)CUd0
.;5?[G5eI:I4EG772:/8AaD#\/D.JD^Z.P5E2695=MOKcGMM9GPfQ8LUV#+5d2FZ
,D&1<cOcEB<L=SS?f(SfDPC\W>>)+\F_P>1e^]RO\OMUg3(R\E3KTU7SZ>HQG?C/
SOOFUaYbW1PA5/egPd]<A,Ye?]:PWXAU5&PGV+M:U2E?Lb&+f609G0FPE2::TL7,
28A0WP4UK?d\f9=N9Y/#2:8=]-KB7Vc0LCSe+R>7?4c^U]_]_Q_1Nc3HR0GBMN)#
fMB=E@L@Z5?0+QGTa;KI(Y\UT0\I@b94JOC=CFTU0Ib2g/@]H4M:e6A3CY&F^GCH
D4_:Va\7@-(c+:-(&+f[Y^F(&7fGeLCJA;].:F9E.V:aE4L2N9[<&XaG5@U?S=(X
c=@Ge^2><[1CNJKC@^9CB^efA(H;N,/c[25;aJ?F6@/Cf2XB#EES_,3<fYJ&4G[U
5<F;0([Z5PE;1[FOf;?81egI6((0.4W7_F2d;2W(^?I8??)G;>WBM^B68(@-bLgR
(/LNN&#]SO8HBT8fPS4TL&//[)8cbc66UUgPOdV>=2QOFULRL3M;BB@La-U4SMFA
,gWgQPE\dFM>c//cX3^27>c3Rd5M^DcZC6L,VR+,\7S:G_S;C[,8?,Y9+>_C2].T
#PLaY&]?eCT@#=L(IBIN(URbG[M@J<DU\UVT/_<]6&YID@84NY;)c[ag40Eg^7bJ
3PWHM[0LaTAOfJ7b+4>A_gH;T.7C^)CGT#GBE[YKKR6[6X=J5IS03:AAgZMQLQ&D
>\X1fT96,^>L:C-d78UW0YD0d9EA5AD_X[6D8_aeA_0L@_QZF04cRc8AV-IN#Tgc
C0]ND+LWd&VLTU/)H3CMIA+U:?5?+<O\O-=@FWH=gZB=_SLE/Y@(XBQ#/K9@-5=<
2K\5<EgB9C?a(TXRK&GH5D]]@Xd94U27f-LUZKRA/R&(/8KLMZ:Y,GPLT(>2UBU+
#\0XLX=Xe\-59@NM8^W-/DcO293(.>gc8J2<N;EgJTCB)P>O?9Mc(>?=0aZ(b:WH
>L39SDH1^?Dd^?_Q;M>9K)+:,@?>=M3\=)ScS6R>c#?CW>CTP9B_;\6)UB71MZ99
c7ZZg2d;+YaA1X64G;F6N,R^YJC/daBQaCZ+:.R[a.2RU90IAE1NdB([FP?6/EbZ
52>#7:=L479L0?C&UQ8b\1^>IE5M?U6\2g_E@,F[T)D<;9B^I=bg)F2J.b?FD@Z@
HO9O3ONag=#XE0H63O^Sbb0ZNS4CTA[#28J6B7D68;HGIU6CcE0GG1>d^EJ[b<C:
Qg):f+2g^]5c+D75KEf[gYW1Ig8bK(e0[?74YO95WAKCUG1W9/Q-@VI-EL&)e)SW
]&S#(:f#dT)3f)?QAVB0f1Z<20c/Y4&.&dgb@I#H\:DcX1SQ5B5D:NR+_?]b46A[
E.QQ+3NJ@HU_:]cAE(g&83</8dSMAa#aBN?5,^/RaH-<.9ZR0W8=JDOTL_3,JU\E
HIHC6[(>U^[Ce&&[XDREdH1e1#6FYaUU1[bNAMZ?EK+K7.16JbV/=c+O:Nf0\WTR
@FM+OXXU&/-9UDLaN/.=/AUc:Q5@Uc_=HJ0&LYK&.XQ#f<#-8S;EQ]bcPQ4([\-U
N51PeF3E,\C_Ja:#7^.#b(OCPQW_cJ)EX34_&6c=b91d@V\BE,8?KCG_C:K7P5d)
5L>S:g9MQgC^</?C.C^=7PNCRS>4I9a,UbG&[T?&<eFE(.AdCc\BY-ZK>X\^6Z&c
2\aXM<Za(I6OcC32R\f__S0T0L.aN(2GG10LD-fU2CNVSI&gbc,PAf\V0?a;+WA1
/abC3Q+ZN>Q.Q1Jf,,>La=:6#NeLK>\;=F).)EF)KR@N3&FcEP+eF>IIF;F]+&Tc
HTccI8(TUFOUaM:K8^AGTRW&3cJ=K?)2=ZY=af8KdD1A[6,&#T.3[Uc50VRTEI]^
.M_//P)-9HEA^#5H54NT@]fTG35@(gP/0XVdT>:LgHMWKE;XPW\UIOE4c=e\8O;e
Y?f#&\f+<AUSHEE;YY;U2F?4A298)1,I9A;4=>+ZQ@H,9-06DO=76O8b7GTP3KD8
XPK9W>]Tg39VZ=,eKLJ+\P\_/(:20I5dI@Dg@b)2.]FWD?7WX\8I\PW;1=;d4ZET
FK:41<Ud;,35cA1RBYf.)DV+_214Ob(_-^dGK+.FeG>d?E1ZdB)?Z0YOf)0b2MB?
7F=>1]5Z^D/Q32670^YJaZMYJV#5SGY[6gU\ePJ)PMZI=-6]G0W;I_ED/Uaaf2S6
IB(4@^EFL3@#1&HGO(Z6S08,B:NGM:D\IC8g&I51MQ^Jc/J0@KHRgH6Nf>[aF>/_
W?LB.HTGQgIbNJ0R_.._8AG8HX:_X1<J,#?,UQR[9dage+6a6Q?Y=>K3L,a,[0(.
.cFT@S]+LTD6V,I9aUA1ZVd/]X=c,8&7[Y-SZB#1(94e/g?8^I:?[6U8Y.Z2e^fY
.L4Pg)<=G3g-(+ddHWV1814gM;aO[EZ1UF/OG]XGafR<3BX/SK6\TX>.&O1aRY>6
7HY#;cRe\71KQcRWV1QU<8U5JNa,S3QR<IIEaWXZWNK+LJA)]DE^=M9eFM7,#AfS
BZ]:6LX;=7;AG6YUDb>=;EZ1L=Ice6M-8aO9E]NXNT=CaYIfTbJ[D[I2?M7ZTAB<
9-f+U3Z64N5]e2:.:e<(:W#BB(..@KXCZM0[(2XM&=MX?P43L)(.-AQF72SW#RUY
2bEMPH:\c\^Id#[K&O2]6HJ#4GDP.,X391I4ba&W##.S:(MA8G\>_2X9N^W+[()@
D2^4#.)BQ.<6_AUPQ4+<4</RIV-aO;\Y-#HNV^,;(2CUDB1(&27OE=\f@#?b_H[6
8Yff1X7#U;E:fKO]]IGUO<=)N,dGEZA,2]e=eR5?bAaS#CeSB4cb:W]^E5=G5(eK
55;SXd7P-cF=V2_MCF:adbL@CL6beMD:7dVLTg[4[d1N/^U5DFb]L9^>4X19C\bL
Q)CFO:9_1]GU6F,57ZfW<L)JVKed)OSJ:Y4K1<VLV<AgC9CT6\e(+GSGJ2RXfZG<
c@E[9/45<cEcZ2OK=VJ55DA)+c5]2OSZ[IUC&\_QUV\/)N38G[6E<:),#1+=.WI4
I2K(f2A;;:A]TT.\-[MEc(K2WYe(],gb]L75)IWR2OUPTCJ:dUN_g,LO@K>Z:^ZL
7ZK#>D+=EK7U(V+JfCg0GXUbD&;C-8H#-PFP9EOR;XMSa)U7b.BX2137,YNA<#)g
UFC3V32-Z:E:S34e=bDeE7aO-+b:dO\?gKeI3b:ED)GP_HbK-R[4SXPGUF^b:0<\
&eXA&?VBJI9UU[+SV,[MN\A<YV[K_#,1?A710/G9;M#9>Z2Rc>EEd3c8NZ0AAH8G
5dW,8,ZX9&U51:gC-FRR>9,M90U:,L8TOJ7fNH<P-2:4Ra,6=b\6WUcMaACB8CXf
>_Wa-JDJNI?U.<4EL[9&NX;K>CUM429eEHb#?ZAWQeO7];_=6WQD2(^2BY;>.TY]
JGaXO6SV3VQaAMSE1:VC4X)+dCE1Y>K)OT/8IG;F1>&/.ZQ#0J:&B?HZE4BC-W2+
?5gL976>^&b=+IE##.YEB@b/,,G9>6MPO<P9#;fg4W)DU#QJITaQbR=J#;9WGM4H
&60L[)D34RSLRACG/F^cAXA>H26(?:R@cG^CbeD<Cd9#RDd,-CE8C3?/ZVFf3gN[
LdcfZ85fK(N:KBV=(+ae:?JM4FaIZ@2^S#+G/Tb2?B;Z5QHW1Z_KIRQKF4BeVT<:
5@??;R63OZOTdaR;-6N_8:M:Dfa7C2^Mb1=;Rc&,6)bO^WR7K(De\70dP^B>aEQR
d.b;ER]H-JI@-dNF@@SWA1)70d5=O(7FA]J4gfO)MXFPEPcUE+T18<BWJe3R5DGV
IReB=1cLGV>\,-YM[-A6LIP9fdWZ:T<fS(P]gVb>.F6:g4AN+IVa2P2/A._D^eVK
/OX\LF)L#DCT&9F[X@,O#S0:[CGU4DcLd4cA/VN/?b7OTF,G_g71.:fJ1C7=8D[^
81NJF-gMM3_KOe,-K==fS\/<-?)/Y8G&8V6W;g),_\cJC(B_(O]R&CF4=,@Le]b#
)&9Ka4__e?^A;62UHReDe8-@]3J_U5(.(KJdbIF(VKH<&?O-]@HAee[B6fW4;=,;
[)#g]D,LDXBdJH7eGM3<A^_^=Ua#b:UB_RA^^fAHOEYHLbBUUL.MG5#=]9(X2H8Q
e4SA=QX7fG4,MCW4bLcDR\5B0eL?+@C.T6@>JP\Mb\Jc&XdXM+222ITdge\))==G
5&ZcLF@f&,:IIfS<II6d&(WWK/M#V0:&Va.8f\Z#ge/GND/<+:C/.NdMWWWMFa#U
?90JLc49c?YH((dG8>WODI)VLH?5a-d,T2[eR:gY<XbUTaN4=T;W31I]T,80M4c.
_)XVb-V+[Ef8b6NP]=O5aVO(BK9Q?X>TR/#O1@P[?R/0NZ&4F?2BOM4R-0JO77@B
2c6e&#C1_K4dZMNC+R)G6@GS_2dc4I,=6ZR0+9<KBF1-8_Y5#<gIOP.)BF9KM1;B
f(,gZQ#2Y<I8JNd1NR.?PeU<ZdTIW)UQT2N[A0?N887;:A086QD\G2)gLBZE+c)_
-.f9BfRg=@GU2YH-Q+/-7dEG),C7fcf@DOY?F:Y?7AAYP4:+W.T_;-^&c5?g:\GE
c4[9^PGUP5(F/Z2UDE(0=N4.QO/;b>0<d+7ZAMcZY>URQbIFf6D_YJGg9I8]@H>K
1T>bWVe&aJUIdOKSc=V;)fX8.@P#EKB3Z,M_EZE,S)8b+c/==P2:e;f1bINHB5#.
Sec.G\.8[JK1KZ&L<:4ONRDM3NcSU8:N9=9IXGYHZ)3PRVSd^T+JZOPH<282,HH^
M>:cA@@H[V1.OEL:UZTa]^[SCDG833RI2W,EDCSJH\\L_P&&;37?:b88)2)1cDB1
_F_UR^24U7PX/dIfQdb4H:dY_F[9NT3-YNEJ_\P>Q-=2U+7a;U4A8a#fNGF0K5]/
=]P?Z8,+0UE,VJ(--e\5d^H0^N&LP@;=0?EW4K0^<4D\FJL7:P3,ZWF?05S[]1)R
Pc.2F>[2fbfJUf\G#U7X85f)M1/ZL74OGSLD?faWLPWH[68]KS=a,RbcD2@Q7^.;
(-^cg^8b?7NA@FP&DUBa&N#-bUc75&<K=/(.4:H+7.8_O0bVWO,KJIO/fD&8\AaV
)GQT>@5+A&WK[PK3@[TNAN33BOb7dHJ&eGN81JKf7Z+0ITWJZb0c=RNZ/dV7YZN7
>@4<HN.:.GZDQ[/WJHLQd4@I89=GcQXQXbDB9D:Nf:2OfJ4&IEC7>bFCKGZVU;-.
XXS&WK0Wfe^4b]>#4[H3EeW64AG;MBKBJ6CZ2=-U5SfQ0OF<=,3c:R9:<&5=B2#-
+R]_^((d&8-[cIXEPaGN7J0dAc0_)MK6LLQ+aJ3cAc\TIG29c@)).BVVQa-f\CJ@
f,KQSVd\G0]8>02fJ(,d(gIM+4K)VgOaE2N-_KS9TXY#H=eS:2)0+8;Y\H<(T=Y8
178AN4MJ,2aTJ8NO;Y-->IM9/13</7G?7LBK.:S4A\R^\^>FKOgU+(+Aa\\H]+ME
B(T[]RRd3=fdDZb^W.E&>3e<-Zg9K8P5g+aULabT=BGc>04<66/;B1+A?.5/9V84
KQJ&YV^<:X4E;cSU2c]M_[?c;DcNCB<SUA[1FJaP@VU\25Nd]8dS-?8B:E\9@@BY
#C<I)73\OX2(&@W)NP6^E1/=HUBG(QBK?3.?/C^ZIb34:+O,,^#,/&U^<b)980We
g,AJ++3YdfHF(T^X^>O0IJ1QOf>HCX];.=SJ1\43(F+B3RW46<9[;1Q-N>:/VXS,
U468W5-2L5(QYF[e?3:U?KD_fBe>YK8R?+J4\b36Y4KYF.OJ@K2;eV:5?#1a\0?N
;<fL;N;8[_?V#(_-3H&Wa4gJE#;G,.#PF,SA>3R(dPZKM-4eaL0OCYd)/G?b<X<1
K9<_G4[C1/RYFRV:&K31Q&fY<86A?0[>D,N;X:@),=3eg/1/K:L,KK&Pa@Y15P>M
6I);5/B@&,:WF7J-Q+E+,NO0ST?]^?H0TFF([TF3^_+e[#001Ca7E[IQ/]F1B[#5
=VNDc9)&(,.)>#SDd>dS\;f09d\T3d/[:cMHS5,:AS_HT^>1(:O]^K.2X;SFcSG=
:/;OTg-I0VDeS;OKN.K84>(d\@Ac/5+:EQe#a.(>bX^5aU/FMbWF10Bd9gA0\@8Z
DO+,eU6[bPX?(&#]M+@JbCZDcaQ;WO]UV0M)<J]2[3WADdaWGXb5#[36cCVZ_VeS
Nb\)_fPKS+I96)X:\2D]BWaEbNKSLNAc>9BbVf93EVBfUb-3Nf>_&.XO(@GQ.Z\g
2X>c&Yf);&^XQXdB_,XaFA>L3EUQP:@3]M6g\(X[Jg]+DYZ\OR2C/5NLRPEDc[#O
cWK=UcA>bHO;#c.NW2b;(dg&KA]-[HVB^<D3TA)8@]Pa&GU(C/KWYWU:U;3G^5.=
d;7&D430gDc?;XHE/I#,Q2.bWA>Q:3X\EZeCQRYN\)RDR0O?]U7GC.Y^551:#C7T
QEgKSNM3Sb.NF;=g6WQ_8\e#GTS)?8QfCgOQC\E9D[Q1W#W]]6@BRA@fZ0d>[Ged
5H[LF4&KIYBIcH74bWbI9D(Z6ebF:BH@d3c:.7<PG)N:SCe0A,?L+8G4Z\(C[(0&
bS.&:]73V+d.:,SL/8S2:g<0EA)DSPfdGYT?6#DU:d_&dB5)W(OA/D<F_)S6@@=f
IT6/5Tb(9&IX^@f51YK&4.0U3YK3++F@c>Y++L=U5F?cJ;^_H[?5][()@9C>[N_F
eWMPLVT_[(S_?XU1U)W[\S/A@g?M/^I>(#>ePPN@]./LOB1[6U_<(J2[G@WFg.d[
NRV3dTOG#HC7,aX#PG<@:aEBYA6I\I.)8)d0>,M7aPBccY^a#R4KB@+?\d_@H\[V
EPA(ZLQ&4)/c(CH]\I?fDQUWURc-;4,QN,dc(E3P>>_?]X-Pf3JB/7SMI-LT?K8=
4WH+\U]>;Q0<=.bXW<cb&/+MVf]^4K&N?ENJ_F3VT\MZ1f)0TXH0F/&I3Eg2A<<9
:IFa-8E_[D/RU&=Adea;SC@<\/>^CL.=B8XbM4,F@\^[YaJVNZH3.O8MS8c].?G2
[Q?7MO7fT=TQf<.Rb8=09-g[61GH_.N6IM94RD=J9dP<B,Ce0X1:2MFJXJ?.&EAJ
6G5.CALRL9Q6\1H^F&H@<:+&OKJK9/E@_RFZH<TA73bc,K3PT_5;c]1T1gCB_&(R
)J]^MbB8\\/Id8K-Z(_&^JNKWJH=1ag0GbT1dcJC<06L8T:\I4E?,JB+L)5OPQYQ
^SP@_S)@M<YP)<HU&)=2>)]VGW,.\BRHY&[]N/)ZVD19ZST(\H)QN&f68@(#2C-5
ZF9A4=aVCI@>]I^28KIQB#N-M98PeO(>6Ve^8UL,U4580d<>?M]&5I,N8&3?EPLG
SbLB+=A-])/NS.O\9<U.F[@/Ag]-Pf>FN)aFS;(VW3X-DMN@=S]LW),6@ZQfQfA\
O5/@[L+d</#,2L,K>KcP-2c/0AI\UD]7c_B9,#G6.BJe;4.)OHDOCCD-VI@++ccT
),K9=&d,X@8aID@a:(T]C/7\=]W.W;+5E6RI_^6T>;_Q2P<N.b^JG[^+M@f9aDIZ
K[WZ)E=&XD@0UEd=CW_eJV>E[X(Y;.E6RU+cbCKB=QTE_X<Y=_)cPN^U/M<WWUHK
2;V&9I9F+MOQ;=cAVL48F+10)Fb+CJMD<ac?/eW8X6;g\44Q\+TGZ=LV/&#5=J>B
6;.H<0aI3PVVdC>-b&1#.R>;Y?H\?M;,Sd>aX-S^)QO^f]cHKHa0-72EM]L8BLf,
3Z,U?Jd)FV98A==W720_&eW:S3JQY87&89a.W@P2G#65=U>>[K#<2#D;/F^KK-[=
cb]>ZHQGDAg:23KEWP[]7fTA[BC:OdD\.dBJ^C_&2_THQ#,2?:XbY+7e#UWBWGRL
M4=HA8_aBII55:8FE7V@G5\6H6_ZL-=_bZM[d3_OY5/C+45c=O)UK+,/Q)eU&]\_
S5@a@Q],(_2V7GeIMNb\O[(@BNY<+d]cDE&JW?GQGZ&AX,KgEW/Y<b56W;Dg?W+f
YUP;XLI7-R3^)aXcGDLcQI>.d&P+8\44XC@-<1fN3R(.V\gGL?C#)fLA0Z58AT<A
_&(QYO37C,=YH;dcUIF]VBI,^C@aWNG_;Z&?a^:<:[T<M/c;e348M=CLa.XaZ9^7
K_&T-d#1M7D,)JEOJgHGAd.=+U2^VH(8d;#fNO^/a=UE=_?1LS9CE.-B(MG4<)cI
/S__V&JJg:OS[;A27-+adbBO^P26]I0C<Bf?cU_]X0/,9HTN2[R;d]dT8G=8&9#S
/4;4+?Q:;PUN-VgO,>T)^:;&1Q0e@\MZVBgW2S;gMDRO<H90\g]>;]^IB2K-K1ZI
ATF7e?15,S@VKA&d#9(4]\f/:/-UBX4>=;=C@?+Y=F^RZK,db-TU/_C;:^L8A8Rf
BFAWB=K+3<bcRTOE/Ne=e,^?AX0>aE]@?E_KKKJT4)X#4/ZN5[1c::8]5)NWUY^E
]]D\4M04d2L:\M:;]HB]SN\KIa<[&1g/U#K[J(Aa<D@HBO74LX7[WB:7[G9[31Z^
DX0@O>CLY;OS\:eMW8/3LK1DI84;fD8L^C&@?0991GZe1[gBeD2\M_G_#7:PNO5+
RPN0VEOGd,ZG>8MI=OeV3VOc]V>W8FVW:7.1A#>L8f8^M1KMda#>dRQFWb9OB0(0
2cHI)3/(G=]QOVX+c07U=+YR&9X:K>9UPFR^-eGT+0W=^T21E.@F;dNSXcA=aXL>
f:9V/_]\;H>gYNb3FVcPG\W4d_c5aEF,[;)JWN^EB.]+[O0=QV;H6ObS9_4B5VR[
#eWZdSaDW96@Ab[G14/>9/RFF+4cf.\a,><Z.SXE\e=;=6>X6GD:dMTUEW648Rca
<^0A;D[E_\75e@030;EVBRaL4.3^R7+NN[6_1V4^@d_18V?M@HQNDSO-^HHHZ44Z
bO2<-I6c<_5,J(=8c+&76W4T,AG9;T]MW-\&#SIY@d7bDdS+MEK0HZdPA@PIC:ZC
1eTAPH-;A<=RfWK.C>(L36-?U7XSTP_g#LMSPA^.g3_9gL7-cA_bHKV>0N0E3=8a
G2WF@6HE<M;0?,57SYE_G#@)eM-@/_E&;ScG-)S>DS0X1\eGG2caA\J3?B6)<TC,
J.6#cGY7Q+Wg51M_)QZEeaZeW\0YRRcA0^dLJg=T(=36<N8gOV[:;^<U]U:PgKWJ
b&CI2MAP@MLC^4BWL0),a\@(dJfeYAFfV3UZX23FS3]J@75/;aC[d,TV6<].U2gN
K(:9<Z6X]&dO&>R0/[X]M(^L8#6TF85_D(7>1(JBe.3/70gS--#)#?KZ.\#7J0dW
3J=LD77O-A2Z4fM.55GR-/K@g=;Gd#PE]I=SB^I+8?-g.3Yb4b,^#6O4B.I:4gE;
Q67>]A3B8M9;+:fa.7e58L2XfK\,OGMJIaBb5VVDS)Ua=RM\4I>;4IEe?fE[C<YM
5,PN\\#K8fe6/GD(X\K61VaG;Y_>gCSg7b5Uc#=DD9B.O.B-#&GJf.1=-bU.N9MT
\]@fR:#WI)<^IQH5_^@^MJ,aS.A[B==,=a&D7b#a,a]H-D4KVVK@X2225__VOgZ>
R1EIYfRI1gWR>_Z[X</X=3ZG1BQbH___;Z15T+gYeQGA,N0C+KXEbD]VZ,7,QaW(
FefD.1##Y)X6:P\<9M\dF2,::+BT<Z+0+0-)-1UYOUg_(2VA+2F-[+aKMCUWBMRF
1T-7R(HNa::a1,&,8.dCO#()Q467?d/bcIgUK842#=L\)#B_7.&g#Wa)@1=<HT20
JI:0&7+)FZ?Zf4C.C38_JXL.5YOfL,f^0]+R3fB[gY^I.#c0W<acc:5b(EOG#,\[
5D@B1=9>Q14NV^9[4)9B@:&@.SZ?MKW)W@/Jc]:#C,8E_VHdPOB1M:bb4V58)4Be
^ZEcV4X-7e4&6e]d\6L92,E4S8gU_;DCXBc^._aaFD-\ad28D:&M18F2Z3HIZT.?
O2ZQIMN;/-^)Q77@&7-;<E<WM/BAN9SgO<c..TNNX#@S\d+S\133KZ494^EY0I2K
[9b>>[Wa,2PI()Z<WAg/CNbRHbW6]S7IH_/Y\85G]0da&F94-XeO>6,=B/72IUf6
?R-_@QFe^/#W1Y(<B.3:dX]I.T1YFM)I8UDNWWT)KC1HH5e997M+ae9V1LIfba@R
MGV;fZN8:3YK7)RFCM)=CXGA=56^.TeCX0333:_>#H\Q2)B1BK;<B::9bBW?e.C;
3&:,,F^<aK=-<ZNOWO)6<AgQ>EAW?T2_.bUb\]4.\eTZU;J--8gfNfeRa-gB2:_)
,0J^QI?dX1UD(:,F.+#S/[Ld9;\V9a_WG:3O3_gXR#YMIUKG_b-0=Nc4(S85_I#/
QQ4LL(@S;>T>6/2.)G6_LVVa6DL29a31&1@XTJ>7Xf<Se.VB5PS<P6:_7T[4;@LL
]T>IZKH_8F(RT&2/2YH(#YA^/:;&0,5[A/09:LDbE-UAf[ARKa2f41A.A;CIU61M
T\Q+X+(W34f&GV>5G]VD6Pg2fLQZ/3.eU#VOR+HD#E;M\78?T8I-TWb8bb#cG.S1
2@)b9F(BO_G_X#-FKKbEGgU=PS1,W+.#ab/6g9)L<M0_)B3F/8SW,B+ES8T_gW)J
IW?/W3SED>_7NeL8.4Bc-QWCaV9HDJb#9)EReAb0.1d3MC3Na@0:RILX]_;e)JTT
;P(21TMCM_\/)?VUS.gQDUC;\5d;<6ce\&<;bQCHV/e-F6fd?TO)#f69Z,4IO728
LdR6N<.V:R1#O)ET8V^[(M(5I4.Rc).6F9MN--/>/=g[Z)-M(I2M67e^+./B5e?;
.:_D#VXJ6TDgPR9,3.=++X#]MXM?1N+\g(/F+7]-=ZA>-?QX,U7[,\OdQ4M]eADf
dQ?;9Re(KCF;DP<1dEJV&?U:6NZ6/5HcA/B7.W3F/JO9Y_gW;g4d4>15PE8CHC_d
f9NcY<1HYON/GSB-RDPd2L=cWWSB]Q5:(NcaYa&6+1UdUd.8edUfa(8T,@\4eGbK
1/-68PL1/A8U=f>3=[Ag/\I\Vb;1AdcV[M(UJ&:AWO5S7\&aG=JT9>M<+Xc.d#)5
32.DIF>\JgGR[BePbYKV[&8^<(3&BYK#[EN._I2@a/RF>O^N;SdLBHZWc9]T3U=D
RXPP7_>QU8WgDN&6S#M-g&]c3FdRc<g]=^=g^C3OeSMPR&U70VY?6Aa[\H6D:@0-
>dQPRgV&\1#g?CRZb.A5L(:,;U3,?^N/LAdC2,<6,QWMS4BNG8&-+e\Igf7+G]36
.G0[GRf\U>L@(a3cJ/Z[O+236?=.CRYVd]?eBcFD0H#V-YD7+THAUE6bdX>>O,#S
/UaE-7+&M@\J:>aBBcD0+9XV;:/-.X09)ME3/bBWT09Of)J/>68TQ3KI(ef1eL;9
97?1b#=8[HG4I:Z8S;UMZFf/IE<VA/&S-e(dD5_J=NI2ZNF+6F3-)_ZMBB0:Rd;.
Y[/MJBJKU<C>1g+=JA9cSSJ<?9Yb7N.AYQLHG<TRH<^6>EAPbL:Y1afILgJE,KZ5
,L,-STe9N04@]EKd].abg_4&X84\@S08H.PJ]/ac5:L<SCRSK0D\bVgA-1>-2S]K
B;YYHVM]>F?a0,2T1dTRg<5efZX>4(8X_b^J?Ga_-e[TM7D6;+^S6UR;#JB]9NJa
2_G<JRgADcS1MBQ_fAYCHLHb[LN\3RGeN\63[B]XOD=b@N-ZS/;P.J2#UTI^-?JK
eX;+I:g3McX_X3ANI^4>6.5IbL;OI_DDBTBSEM?0D>D/Oe]G,)O8FT>e+ZQBT4dd
P)I1&CQ&&UGI(,96,A<;>b,L3LITYYL=S=RH:=EWT4J3W&M><S7<fD/X8_L:B6@5
UXS.EeF^M29[78)Z]T?0Y6YW0ZP5B7eA>^RfIgb6Z)=63:ID]EW1Qc^GI;6<VIIL
g7c^):I;U=MJ1<F[>Sbf9G6JR1LafA+A0gX@<<RD)P&FQJ5V:\6Nd#6Nb3ST4>]>
YRHdQ+C@7?Padd_&_CM<@a=X7;0e_d9>W2W2,gT@VU6dW6\b+T)K8QQXX)>a;X>F
)RgfWS4a,T3YXUHE<IK<R=>&c[<IUBW&P.M@<S4PH1]d_5UV]87&NFG2a^NHa;)M
4RRd)GPeN;E0K,EH;&[)Y34G.96-2;Z1(QU-JXAb)#C4MS003=dW:<PC+WVE?;1T
]56,.#)^?4U>70<7a/MJ(2/UFI)(eCHH+;\@U+PKRJ^LE1;C#FO,U?A3EdXXJ709
31X4A5^aVVSF[U[a]O3VZUL^PZ&4#WHM13SL?;9TNJ)VZa2X<P<fMFEFPUOGW=[H
aE])RUHe44.H2SJ[/M;FT<.=8V70,?_#,_gdD/+>2>)M8EFDBQ5U)5-R34R,e7=e
C._.5&ESMA12S#T]L#^/.Z]N9fMGZ77B2b4]@ce4:..L5?ff(GO&<B>[H@.R2):@
=498Y+H67KWMZR4+]@QZcX/K7,CK[a6c?dRBQX(W>:46N;,VG5WUTbGCM4bY1IY5
R)_(eFPG(T3^M[^68[T-Ne<GK;FBIM78^GDNV0^/bXGLC-9#-cWI9P/60=9P&KG.
F+3;bQ8?(D6:C>TD@^0G1D3T2JeX]OOXTd#OgGYADS?aVL^+O9Xa<c?R^<<51112
ZUdYAEQ^bd:dG.-YgdV5-\.Ge]cNL-+QaKWf^7F>,f:&8T.N5H4TXfH(A22&-b9U
\cB,9L94Sb5>KBFM<,=UGb=6.cTDXJ99F?X:bG<AOUdKb376ZaI+8[/)CbZ+[Y9V
1N?O:.+3M&^dR^^5Jg&4=R1(\7^@9K56+FXA-@dTDD/4SIUB2EX[ODaF^5=)P,:7
)B-S[3;8UMa[-^W:&.#)>9<_P2M6DT6B=B/KL#=J<V]D#3gBU0>)X5]0BY^.V:T(
1NH6=.JVN^&O8gPC__D^8M:-;8aZ>/CdIN2H-0V]+M6PRLXO=e17B0FN:Y_0H#LX
_9K0JgSGBX+&3=?AS\,J[)Ve9)U#TMDdY#-AYCSTbN2FW9M7g[H1RJ0S7B1D_RUD
1bU58C(L_.;UI=5CE-/)=\Ba8G<BYVOB/eI-]C7&Df,[g6a59Kc6T50=HcZWd]>g
(C;6SN48\<GUIAYN4cGIZYFd2P-236g8H4N/UE1;YU81C&O92CHFKZTTP1^@f?1H
KC>93bJ+\<gX)=SI@,()PP\3\LXMZL7[)=Y\[T=g]7->S:@[+;E8d.29<]HaaK#P
-ZW3Ke(C9]^)BdF7(59>-KgMN\SQ)6HODG3<gZ7Gb4;P,(_[2G)>N]bIeLZEAGA:
B#-,0NFS=E5L_U.4,.Pe(aU=0@C7VaY>9DZ[NdI?\Ib,Sf<>R;LB)L]/)0(T4#;#
[L854R791]0b<UA@(d]2aeX]CY&a?+YKNB-\;R.9B5+D8RVJ7&YP-I7VE]RWQ.&c
[A@&;L14&CVS\;&W]RT9fe)<-gG4bDDeT>75VVD^GSc<Xb,.:7#006^)eTH:WV;_
SSKC(>bAE^:4@V^eP]G=1?W_40TB>(++ADJ/:_:XB;LW;a(0UHN:\GGTAX,5S396
\FABIG4DdcELR?;9NJ]dS5XNeYJWbcA\PS)/PUefI^Ab\f_4BS=[&YO>E0f.Sb=J
d.,4b+,6b>a5/8&H8OaO@O[^?(X#0C8RYWF#MBa2Pg9?H58[YM\fX=f:A)23,f9H
e5f@d2SC;RK@Z0eROb)U>dfa[ZAS[G827Wc:/,acF<VF_/4FA1B1O9O3Sa86ZPB=
L9gMdBGA\[(_II#a#0B(PI4R28gS+_C>QD2@W+US62F([_bIM16a>e79\SB/;(MI
)&X4XXP-PgSf42E\J_W(JP-(#7P]LV91,:d1HOO4\#O1+XP:AbWg,PI]AW7@UP+I
Bb:<(.1P_cO3PQ>+A^(Nc3XLDNY;,EZS?HG-Q^@3F1?<@\aQ1RO;eF)Z;-&55I(@
TeS8Q\P7,F0DD?UD?7dQZ,d5],a:)UWK5BT841f.N_+FIA5CD50aa/4LV)YY+XS+
2(4W=)OEX&;cE=H@Q5/RMT488@)_B9KM=]K\Y0gGJO94_[I/aW:6]FGGQ#=7(+c\
E>.LF4BL3d\WXU85D\XeQW/GK_&A1J=VR;[#f[7M,.:ade(7ZWS#?9>_SY-F:_F1
2.=gcW2A8ZG9,K6C)7:UNfI=<dZ^E.RLGfa,F@aGWaTDGDK-,G0ec3cK2a@>NK94
bZJX7)X_XD::LM^/Q6BZMP^aDS#^#+ATRb;1B(_G:#ID2433e@+CGPSNL8O)H)^d
(U2@bVfX^gX8VLbO:XWC+^2C234NZ[U]^3XD@f=Z833<==0S/XaAY[#=e4.5O0.+
P;E;-,H-YBN@.:>98]0_Z5.7=<008=aHMTf&;QRgP<d)gH&c=:;0CY=8b?1aB<-<
)6bZ+-&(Z_LS]&AfY>c9]X=?[:@c=g#E:X9fQM[_,W)aP[@Ve?IRae4BU&_ggcDS
G+WPHB&<=WT2-A@Y&B_H8A710F]e&6g1g\CJ(-+,9g8FYAC^Gf)<8FR\3O/RM@TZ
4[bI<E[.T].fQH@0;JQ?M6]32?ZOB;S3Te=TZ?+[DaUP1T?)CZ_JS</U?XT(0a,J
^6_II(Ta&;/FgQP&5@TfC5VH)@K481gR-3g<1R/<O=cd;NYMTNbH(CK5;NDM&R1;
Uc+RQ\D<f-e#D5()Ya@b_]c;239<-U6QJ4G#ca\fM@LfWCb#2[6O:Bdf]3cZ:X;B
.2737MF^&G9.)Z:g6W#V)..-4DHTT:86J^daAfU1H):M+@U6GW#7PCJ^MZ#+&GC:
7dX\2a6c@+J?);S@^&:\:9?8OV?TQY/-N2D0B0T#O[2ZTRMYF5dcL/G53fDbFSF8
@Eg^\99E5BOEP8cK+-P,O;_P2OT)T=+5N5PBU2f5:6aAa,;:0e_WeSc?IYf+YF,#
)8E3\aZ3JW,=aW0fP7.-@9R(0P--V09O(DL39_O(&[J<g@T)eP8GBOc,7_UN3N4?
<ce9?X_SGK]3A,Y@1?40Z8cOS<[JaH2GSX(S[XG)7@=a^F)C^H^b=Y?;cU+;ST@T
X2:JbQ)0N6EAWMg@f--FY_E^@/ADDTadJ]D7JZ2c@A4._L(A7_0D:M2b6\K4ZX=^
7B;3V1OdKV_eWZXDa5.9@L_2BUKAfXZea?_g)B7XZeQ_534<g,_1VfW2a89C)ADV
a2DOgK9Ig^Hg^9A;+-\9;OPeA./[LZ&2,L=>3+#Y002PY@?R_4SB&2SE-EPf4TPC
a#7QI_H]KbQd[4MPH6F.PfeePb4)K=(;fKD[GJDI>GbB3HEFc9+>J_1EB8^\Q+^H
MBBELA^R4^Ba?),cLObWDE=FEVE<HaNC:<K<HG8[2I5^\cC#]f]RY;Z(+fJ3@^0=
FBgX8.B8U8]QKSO;R.f3_5I-<c&6@WWg==e0,.7cR(XL.fVB/(UF_aCg3bSSK_2R
:_XM2_6BS&,H.BH6HXWC)V_)?N9/N.D[Pa2@M-])T52H57gV#E,KVY25)/4KVQ7(
RVL9DF?/4b:0[-##MA9C,;0gPgTL;5<81E?HD,.9@(bRSKa(-0fP\&aEKS:PZ^]G
9g&HPcN9.Z(F1WKH<@9WJaOJYc_9TRg].e#8KdEU?C(<R.fKV]W]H:^^FE&6LFY1
:ceBQFVNQ;+2IP5/c5eV0GTcQ4T1e=,Z/-4.PF:=-:_,LG9[X(Zba3#]D)1]BJ(5
LTHD3>B_.MDE#LaA9DM=,.a\,6@Ifg&_e9dfd/8P(UI]]K\H0g&.gJ(99HM4Of35
D\#_<T]YS_O\C(6A:X@NB+McW9cQF9S3e_A@8@JUIDM+&_Y(<A:/^6YK;E[^-&c)
@UA#39=9I2P<g\cH)CBg>WXI,/3O>/MI2SC[OQ:g(,dIBDH?4c=/](7dG>MLLMK/
dLRW><Kbfb?[-/YfEbR)P\&-20>@M-YTF6/dPL=3CUeJ-]S<>K:@B<L-4,89&BII
2&c<PN?>W2BJ<+[SL(I5V?fUdNJg_13-#(3e=NH<a)+KOcD2aTR3M(-JMTW3BN)F
-1AS0KC.gAFKO-#4eBU(+LI8D(2gVX0,]Vf>E0(F>F.#dQM@TgEZY-#\;]5Zg]BC
G=YOHG=:LaMKIf0ScI[0HY;F#5GUXLg@^Z]&cP2?P+D7g[1RV?>KIKd@@^?fR290
&69GPQD<XA^Hc)4/@S)97D14ee:9;U/>bHU\SQ(0P(M-B)7@T84LQ\=8<d<6>SPF
;9B-U(MAEL+D>IV,[12b3>Qe3WY8fBONK.PWG)a24#+C8T.7]bT;/KC_JaG<8VVF
a)?F+SK;1d+S4M.EV)07a5[69Q:<)5g[[:NRR6/O0JOYC:YPVV5Xg>>[2gVF_e#D
d3;ZK1ETYP;CHWWJL[(UcNJM4TX/\EJWUUJf_S@<:Rfe[U_JH76BTfMA3.Q/6C/V
9RCII\-N\T]F?D>++Y1TR^<=(dgdK0=]0_NQR.,:V9TG:-RD<U=(<)I61[[WaIDc
N?QHPb_/_28dJ[3RR.VgJ_YL.9>ZI6;[g[L+#,[cHYF.^=^+R44D9#:OXa/E\,::
=.(ONBY241/^HeV9NS4cg0+gI:Y5BT8CLCELRFDaXd\B\/:fbQBZGRD;,S8ZV-gF
?6L0gHd;G4ELEDWI7RC?PK=e8ZV^1?_BFF,eZD5eagFf#bE-TC7E\]gT#EUI?.BQ
1gcQB]FPQBU5\>RO#Kd;@EggB,L44SU/.E;O+SJN7?;O5YWSI,.FJP,F1Lb/]1^N
^>8)QaMK8:c-J@LV5fUW1GN3eNdg;O[9)=2:N7FHUcK5K2E<3fX.dYUJ2P^g.BP(
GV[F4:\\3#P]:aF#LA7bBCI:R.;()Hg##^J&8?Z=7YIX5T^c;]DW<92T@Jc3L\5?
7;@O0:0PXcC@O4CLZ>/C:1PH4_#Ndc7/_a+K_fV_JZL=XST/[)A6+eb29+Gfg0Vg
,\2fAFTF@+HV,R+M]F&2(KcI);O.;SS140]N\NZMO[a4Y80ZKBG/L87Ce2I?@LGf
?\Xg0F(.BSNS)))=P1651KTeL=bC+-V2+P3,5PESG9<;&)B:5[^d-);UZU,b1^]R
-g+L;\TO1E/Ie6Y,W6c37^YBE9K/([U9-6=;X2WZTfZ7E24V(L1A,Y_KL\,,NDR=
b)JDC?3WL-8>WXG3)O-79Y^I\GQCHb.F9B;(0^<7->aFDK-]e]EQ;83YPeAFQW4-
]]B6L3IaRaL=e6BC6g&AONH?eAaP(0/dEWefP(4]:QXPEAW)PO5TPeLDFZ0UCB3+
>HB=1JS>c.Z#P>?<RX[eCL:I7YIJQ[fF7aMe[eJBA<g<4[;Ab?;2>a6X]>@N@f=+
\ec<Z)3#UBN86cC7RJ[ePgedHM27W3?SK(^OOI8#2MBSe;AJ?_3,HbaE<R+^g=/P
\5gQE_:K=f?[=P6gPZZR+bI.TW:-Jc&0/[f9TfKS]U74KPdHWCZ2dCHV__#33E72
@;_4fc?#ZI?X7HJ-QfR]&b.cV?]OX.Oa;Z4O^fNEc_>A(?BR&7=]HR=c^aFOJH2O
>P],B_KHfe3^FgL#+#M_UEe-ecE2TW.=c18OAUR0N4]\3WZS(1^fHWBgF1;6<R;f
<B0-04edHWT\(E7/CI#;\C]d+;&U)2d[Q8XSFc1-eIbHcA/fM/Q?DA;28fCbdO)d
]HdH5;1a5Y4g4(2<Ab(7VA68,@7^g5+)OO>0e?DN<QCMGZ8AdeM;a_B.KSbGOVT0
XPaX;7]57;5..Z)/HCHG>1KA,7QCVWOReS4/]5B:WU707(N&R>6E7-G8P?1,C(1I
67b]+IS)<b)e.c9_YeH(\(3gY1U7.a;T+._DRDO^?AS<RBd;9R+K_:Ga#U,/T0SJ
=#)Q>EXZ:PRO4AWO(aY[V8d=(6@[WO:J)TTR.+_b8.^W^^QUF.D1ZZd[RGOE?_ef
LN>3?X5^\KVEOU(^IH_cFPOWL#MSRX.#R.Y?9A:D-1R@Y)PC2A@1EE3&84X#/[a7
H-eR5(ddXAY@b(+]2Y;\L^N,Xb<^JG8dBDP](MY0=;Q,dN\a&2@,P#dA/3efGH16
(DC\A7BQ[?<3ZL1OV+-,FOdD==d8(1\#.e@AM>X2eP36#6;IK;eJ^]KAaeU8)<R=
I3X[e2H.[8CDFJEf=72[PUX:MaE0OO8HK+5f538dHBQ88K,SOVRC7HB@?b\\VE[T
HHKBF0/<<=DI5bF/?P1V_G/.(^I;F@Z-K?<cRI.AEC[EcG-1K:NOK>@#H_<-Y)b3
@c0ZEH9A^Q11HXg164Ae?7E6N8#T]?W6>:F@_?64R,&MgDL6K,GLH7Mf(I@))7(?
g;gd>K@Ie=eJHc=P2K5(CXO^&,VZ5XcgY;CG1bK2/N3K/YKfc+VU?L)M_#_L/gOI
4Na9dGC[=T=&+WEfN3NdC[=))BH)7#(1]FYf,a<bMP_6L>0<C4/10(Y-NcbDW3_-
@?\&)823&4MT^I)OI2PF[P(^L+f3(.\X]ED2;7IZHFbecW<S(2eV<d]4Fg.63M]/
V\>\^GD>(,RXB#):P[a398a=3C/6Fa\4\\(eI:Z7Z4TVZI:RDg.XO18^O/.QE7\7
Y)=61P\GFD[<fFgRfaX=W.<b6-]^_15UgNO1<&1C1,;CP.cK[eZ?31>HN?K;#7:-
2EAWP-Dc89VV.D=UP-:bNS<f[;U>dVH8)??@7fIC?=<K9A_6&)R<ddHV3HMJO:S/
D84TESfd)7_LX<X7)]VR9IXBW<-GfQ4-4FL(:5Q<Q9?S6NSJ\6K.1&f^g;/QN+Z)
U[.6DR.6&WAHI=2N,J3QcTE^EL0DIULe.[+f2\^QP1d#dWXR)BKJE]bOO6HTDD8<
HO(U0W=62eD5A0EQZ=eX9Y@;F&.I?A6>#E5CD[SFGW]VS1V1)=.eL_M.DK,C./>C
Pe@96ULc?M_Rec@gQVSBdVA6QU683D:]6X#R31)#?TW@GK4gHa,@G0UEAEb=K,cb
2c2TV23G?MWPK:+)8SI>\cK\2X&ZZ<=S/C=Q8B4AAB5ON575@4cAV0(\:8Y^LccR
=16YSYBeA0;?eEJEWQQS?:)9;5OS:db;I+B(a,^)OK4]NL/R87=34:S,7VZJPG0M
F7,R2,:/<gIC#4YbU\=@BfYJB1+BVEI8L,d1^Bc.]#7R&CB5HSW64?2a>,KeJ8Wd
1;GYegH^NBN8/0BG[PMN?6.YEF)1)3B7OW/dJVN/g,Jb\0;d46F;DaS7P>>3)LI6
GTL=>c2M3DXf=5\ZK4U:P5E]gVIAC/V^N(f11dP1#VP;cce=Yc#MIHd-4)(Re;Z_
Q3R;&cgWRY?6-4=A0b=OZZEHJ^bEP<[I26I6&<Y<Tg1W<gO;TIJ;L+CHBAV7aX=)
CYKJ2Tfdf7[dB@eIA0(bL8UGf@M/NZNg/7NEU:C<Y>\Pa5cf&=KQ9UDP>SE][>B9
#DQ9bKG@IZ.50MG_d/C3.FWZVc^O?HP,9Qaa>.02.9D_5WW7#_Sf?aW<2DOgeH;G
Dc9R)S9SJ[78]KO)R:6]G=3_OP-2)UJ=[\KCSZaVdB3:6\]:#Z@6ggeIRMBD;FE=
B,eb(K1X5:#bRBC6UDO>=cU9=W@:La.eSYH\/EC7Te2<EY2L;F^=Jf<QgHPWaL=?
^)[DEKbG=0=d>CQL&#\.#NR\b#ALUL1(=_<4XAf,a:@X6NfG0>b3,.&=+3F>=5TY
8bV]=d1d(fe_AS(]B[aTL^)IYXLS-@R3P8.d+:a+1B[3Cf<&.)H1_\gOQM^g5F6^
UVU<=<I+M6<^9<K2be[SFRY>][/YJGfWI3UH1AZ5G?W9:3b4_.)L^I,W[X0V]a/4
.gF1\Ba8J;7_23=BUSbOB5]5],VQAGXXRTUEAI\PF9)Ufg\S/P5V96J,aJ45;Y@9
;6M,UKGW(];T#V.ETXIOeOea5BL(f/FH@FeQ];FT>,e;IfR?L<9[E^?BRfB8dB_X
:d6,Qc2[/;FcW;(/TQ\e^.U[[-9J2/7EQC>1N9:PX9<_P^-9DeCgP\BH@W9NB7S[
bS3PLf9c_]U,YR78,L@>1[W:0D,)ce7aV,cP1KTB6?d1^XA+7\]4R;[>,Va,]NZC
CeMP9\_Y;UGOc^U[bQW[-+#M^S^e]=@F.^,Jd6f.?2XeS1f1)A7a&B:TfgS-^LQ_
b@<^0:QQcV6RA(1WZgD6f87ZGea0>MaZ.0LM8:#cf88PD9^2P_aG2[cd#RUUe1[g
#IMe)V:3?,fH\<&++b#e[=;f;.gZ<5_4?TX(cG[L=]c;F8CEYDRD<?W4P,O4-ZU)
AEAg=9Ng)0@C@F&T87)bZZL/AO_K6N9QB8?TbT<9;5(aS+F5^b.-4c;abR\JD9B,
]PcU9+Od<a/Q9XgSK6N(F<L=9e^>J9LgL:,dCZ(WQ,YW;:P0cGSJ?/K]W9_YTO2L
Ifeg2eC>V[>^))/QOWf?^]b#AC(^GbAI?1)#V[d+LC[4OC,O?[,@OEA92,RN-cF2
B99B_:&TaNBgC<X6^BJE8bU)^]6WY_LJFIfWZI@WICBSOJEU3)FS:K7\MN8@Bg+2
@U+/A#2]\ES6ePAHF#;THX#c5fYY<&MW8-NL+6N<CX=Q6L^/=HFZ1PeX(-a7e#Q#
69;EaNLCQ518PRWg14MJ35Z[>YH5<Y>I>LHbQ,&?JAc)3ePCMY\3-=+YBOb4ED2Z
Y]MH30dZ2;&=AHgddaS+N[cXKG/54E-TFI))IF=;]dSgH;()W/-=O\H?;:A=;7.1
fcVT^dT;ebR&Y=KTMOMRGB&AWdB79NRP.Wf[e3MYgef-4N4:5+:L23Q[LTJCDSfa
fKKeHAPO(#=QYC0I?&LZ9U8<TdK@N8]TM)N.;<DN?LAZ-3F5VfY.g#Y,I;6/42-R
AP6H2)N[8PCWL1L@R-0(\KW\&,CAc:eD4Q@6D0.a-7HS_Q5VMP)4WT##16F58=L<
0J7]8Y8P0C.5I\?UJ51Z]7:5F./_Pb>V?-.N_gL(SgO;637ccFdER>4W5N5\4ZIQ
.1SVXAd&@P6<eHBMg>5^>g@1BCM>BcO[YKA=^cU4+)/&>SED6Y^BZW&\.@6(F5fK
3BeXafT6CYX?fUVg+4]dPC1V6WDN[#dC;[0M)(6b^B2#]8<CY8S&;2T#D7cAb=/6
]&T;XTVYY&E1Mgga4IgHK<a[3BM:^d?TVO\G1Ef\7[.MGgV5AN,QSGR&Odb=-G=\
6^2.MRZc9&O[-]F70bIH[=+5_g>IPBG5N_aeK-F6J&-d19f#4EPH,<II\dfQgJHS
YOd+:W&K.eXaQY[LcSEJEF.W]^YUPKI8,QHXF=SZb=gN2f^c\;aMYbNN(bGYBFW\
J12,+,g=D_:3&BL-O(LL-8]aeg:OJeCX;>URg;cf@63H\2.QeaQaG=?-2R@/6,2@
/f;7;/#@.dSJ\K=MG2>,(+=2;[eKJJb7ad<.CSV,8cfAFU3MKeTZK6-A=8Y&JgM[
SR&&XYZ;.NG\I+Ped:AF64RP02LYWUJcYM4\J.;dP2Mc]F?6+0,Lae@gGLK3QJQb
\UaPg97)W@&#gUS7=-B+W;L+>@\6b1/FT49K4>:V?I=De&ad4&;Hb4^Kf-(Y7.>G
[PURM01=RF^]<S.>49&EVDB<3]_K#.01ZgN45FTK[E6Y.GFd=TLVRB^fdL(<6dQD
.\fbM[Ac(TYEKY&;R0O?3[M;@W[GYD41OQPA^a_?f--@:C>TR\f7c3+2_,IYD+L(
>Td3g6dDXB^&Q(4Ea3G7<ad+3;CO<18=BPD0<b7UCZ=7fTb)5JbN04VSJRc8R7+2
V03();@1W((O1/M.MC9f[b&F30K2H:D:DdNeLT@6B9&cE?22CbRe?38XF)(N[T[@
TbK235U/3(@,7;GSD@8URYb\IL#@H;E<3.8?QU,<,@HK:&);#KS6[39ID#/=1)R;
#+0H76G0>>6:M.>>8(U</OD,]\5.>.;V=&XU=E#9\]FPX46M^;J0aW23FSdf6Pc^
APfCX(@3V11E7&P7S]?<5.OF^;>3[+)e=/;;1<S\CH5(MHUJAZ<=b]E5ZOKG9+d-
MFD9AV);.[M\[K9Hf5>&eQKJS>gHbO89YXcJSCGCa5^adH@)Q+J6eg>2eDeH<FFV
0_8eT>1)d+Y/3-DR-Lea0[XM9,8FI6JZNF]L@LW=d@O0b(+FRQ83OQH/CUdXa&c6
YaSL3DSPJ3gf(),0F<Ic<V?9;Ec=:D5DG+Pd\GIM,1+AEZe&]&VCIBN9PJIWa:18
[/\SW\OcVF1,KWL>&Ee],Zg_]0^&@X,&Y(5V,?MN5a;YFFJfRJM5C.5RUdLD\9R]
#NVE]XIJJH<5^Vc5g#9_b+9C[Y(EfEdW5MaaI1P>LQ2>.KQL8R/BFb#(N\2XdNK0
8LW4R7K#@OTD<E-SHD]1Gc/1.(e8__IXS8G/eWM82_cBX@+fZ=Z70+==9LU.7f>Q
f#&(VC(.?aJ_]0#Z9VL\CT]O?<_>=6J^]6+LS5.)>O.Y(IS,(<6J<F0_9b6KF3I&
\2Zf[N_U9bFRS=1bA]B&CLdJ1UMW_XeRFY]1gJ0&ER]Y7L5SUF\GI@_fKbYY&e(&
M]d^@TfZ\_#>9:S6#U0Q+dC;8<KZS4B-?fZS8./2YLe(MQL-3?.Y(/GT#=\(.M5B
B:eE+^KJe\G0/U-6fBS#QaIIaP)(DR7:N7Z@^9DLPLY]9\0WVe5Bd>M[ae1CGggB
/\AC8W+EB4+N31YeDVY\7O>b&;/)>3#Q4^8A30FC77FC;+AVYWgTa&[aGLa#-;P3
9:OW(D?YT)dcN@F8WaH/4fc<(.YFQTAGJ@T#AC,=?0aEf&G6^@R7=0V0a-]Yb=Hd
N^e[]OB]MWA4/3G,^;G4>E]/:C8JZJNG\O25GG6Rd.U8)g<-?8Qb:b0d@PcX:A+1
J;HRXJ1))ZH1GV6a8,(24\4d/ca2=[FSe#TH@a=2/ZU1,&+H?[=7JLT3HOD-#>Y>
5O5IXVbC#6CR17;IRVA.AFK6Y52J.Oe@5JME\4<JOXR)WE3BU.adDQ-eF?/5d0M)
4bT7Fd-.VdM6geObgHg/1R++7\XGIZ_]HVF5Ld3ZL-+)28E/gX\71\5LG8^NWO_a
8=;De2eU_/a,P_b7f4?)#4-S3,);dD=-.Cd@#6<(-,A).IG7bP3_TPXZb:UCg3=g
+<HX5Ne@-Y_>78528#&H\>bDZ+BCXb/DcBO0>T.TK:a7?97f5Xb&J9cS^8ZI8KXa
cU0;?Q,6+B_&:#^UO;091V:WKV_4UU-C#UEeKWfA1IVVRLe2PeZ]/^V_9-T@-PSV
80C>BV(VA3.E?K[^(2XZRT_LO#f3VZ=a:82=.:e(J4Q.5P/a4,A?7_;2)<c=]RcW
T,5[(>DR=#91M3>FMD<g4ECIO#6c2/[0N<)=2P/Yd/CLYW.GOHUaOWd;UF5:GdYM
W]ID;?E(^9D=\Cd0;gZ:=\:+A&Sa#;WJY]XL)63E(=1ZIQg?RT-YSbF/T/c/R&g(
289_8>)/N-BLWbMd5>833<=V_5]6XQGU4N:C)de8(RL]Rf]8?fIJ>C4[4DbaUCXG
GFKDW)(e4eZcRYTg,EGLY^?],^;E3J+LS4L+JCf1]5\RP[.Y-4UJ#ZIc:(?eO)UU
_]UO/]6.</Q/JVC,TYQP8HPQb5Ta,RKa&(\3D)cWG=HV//?&Ya@/)F,P&CO6R)Q#
FKE:]R?f03.T0;VVXTAT?PgWH^@NcF(>3F@H)D#VMWYWW07DMBbRNO&6S6,8FbWM
0,Q<MMF_U1HTD@^0.5EVF_3;10]-)f^?DWTLH36Ef\WT>9.E5:?.N=JUaLX-/8Za
3AWfCTL,S5:ONc=Y4)eWX9,QZ5Gb+1bDL5:#C&aM\eGQ736c^<Q6EFT_,8/aGY-^
=NV[2dU+<MI=N(e7EEYC+1,KacA[^G@VMOHBUZc@Dc#6a5?ACL1eFEIJ:<EU&fGe
L,[H3&=L)^9AF7[?6Od>A_]<c3E]Z>fK+O=[5JAX20Og@FSELSTK1YbEH@=/J-[8
D;ecZ,DW6LB8Q]LAWW25&DA^X8LSX>A>\1OD(g78MK@O7_R]#J09X/I9SE4VgE.f
&<BBZd5FX2JEX8;N)f,dZ\1#E^MEEU&SRdL=_O.bD,;QB>]E42U+M\TTO\)c.Z;S
&3VF[)+)J1.9g\;EEA@VV?bXD50(F=BT=<_M&+@NaNML3=Cd>eLPB/O9G=/Q(d.5
:WS++/UY7X/E;+P6E?51HU^6+B9e3?1<RL/2_\4Z[2<QE^#)7T&VO(OeT/5-)O<_
aJ]Vd:N&PJ@LO>FT9B_6gCd[GgXI&Oc)OV<,^MAAH4JZ]CRF@;Y]XRIU)7^Y==CR
eNX7W;D=)(9H7Ncd-OZ.L\3EX?T:@,OV@IFa01_+e:(R,G^Bga(=HMQ4=+@\.:G8
3)\+YaJSR=a0gG\8,?)KHR3X@_gD2/2gN_d+d-TCLA\7W2TGMfWN=W2-3ZP>8\@1
5)g^1)RPN3U;2/^V,217Q+RdOS0f=94KMMbfbK9C+89IJ7QI#-a=-De5Y48bS:R]
^g6,,>/](IMANB=U4>RDT2Z\e)Yb4F26bY6J^ae<GWD)1[N_@5IM.:=dOF.&S0ZU
TdG#[bP/:GQ7J)VE=\AUb825=NX=DEB]F+.(d_aI+4<9L5QDU?/A)U?5@EBR_;cS
Z;TfV?J,5/Nc>[UL/QPQ3@WIdMe=0PK1aO^=UNE5D+_c=R8Q(-f)<>Qg.9O&9&3b
D6P&de\P2cVRcN#\>cP9#_>8O_B_9DSB(]7cFC21K3>ROK<C<b;8Od>X.e/I\bI^
:+:86_Gd/ZG,>#7SBLMN8XS:b98NYJ4@E\+R[NI4MJ^aJb-aBgM5gHHYDF.bC3:[
(4;,-&4BT[,V&2<6RV1C5(aa9@a^&&N;.g4QO3++9#\KDcZ+=.SSZ?5P9&J:@PRe
&[SI/IX#(AJcdeA.&(,GVRH646YSE)(aa;5g7LAB>\^E4dOL(CLF)MRL]ffG3TD^
<:I\0ZQgC+<A80eMZ>LKP&]Z63O_+=N(J+QV4bBHNfHfeU\AR^ZUF,PeOg\2/S:e
UQUP5Bg903Ud(3P1+HCSNMH^;N9;9(.V9-7cYI6;]8R6:;QATa<>F\(EY;NLQBE6
/#@TVe-2K<:..E];G>-;1c,GRW^1H1eg+^#,3Led:SV1#V3C85[3A[;)#<>[NZ^4
5NS<3[6/UZbL:J-b^P+YJP_R[;3]I6W#V<G^8Mcc#0[//;\U6AcLY+a1?04_?NOH
X0&]f0@,NI[COgJ\5#=((01)GWcBH+dUXF[(X;-S04M,VbNTbH+EYIOB3E#?SNNW
F_F@cE[(Rg]g#D;g)043R0K^\PfaY:2Vf:LT++TOX/E.HfV0(?Od5Y1/NKffN8]Z
d@^D;aBW=SdIAg\,UW9T]P>JT^<8)20&\IC3fF0Y-@>XWFZ\\f4fW[f_Q2?S(2G/
CP_<I<R5I&8PR4f9RP8\V3FH&cca?RO^]-7^6fP@SaT+;C#@4aaGSET,G.UA[fYF
4f_RWW2@3&+TE3A0TK4WbP>_JLW2#JZgJK-,&U3DaQW+7DZ#3?O?/SJ(Xa@@cQe4
([a#W<2Y6E6ad+-Y\V[W7EScI?3R)2)C;cVdP,gcb:Cf5d?\]c6TMXTYab@TG5>Z
V=KR<>5+]g+LET,7fQ^RWE&+B:Q?d;O/c:c:b1e8KWfH>/dg8HX\2#D4e9OLJ;8X
^TN_#Y@+JD>6?T1f^(QeV8UB@)2\+XQ/&14:cLYRV9AL>7=e5G-BT71fBNOgIJ.G
\ONJR:a5/H9&XNf=KKZ6>ca6fM,I&ETZC#c=Q-SIR#(-J./bQTL1cBY7FM)QR#>(
A0Qa_#3Lg(REJ_2UTOP1;a-]cg7P;MT9Ccf@8R-4&POLGffXC#BAM&M,NKTaQ1R;
NRfI;7H:(Z=_c&/,8JdD)8_#.e[aW^?9-GD94;(ZR=d:bFbVC9>/:J>Z7YB06eT/
Y^We>RV^?>>+@bBgZN[]9PDTNP_UD415MH-f:BP?C(0<9:]&@FQ]8SUD\U6=A])I
M<R^XHL2P?E8R-fabVE?SeKf:?>4OOJ[8G+HT-(LJVB-d0B\GJW3R=]?>dWdRSeO
_>a:\POMHXZAF3)bT^A9T&S)4;9CF-J(,01],7KKe;CH]LCD/D0,P2XBQPIDE)1,
?/(F86AG4X=4B#,ZC;WS=Ic7O072?K<YaZ96F^fE.#Bd<e+48a986F>/:+RKD)),
0dQ90K/ST3;-Z5f\,LB6?>_)QM/3+7N&&7;5?BN#>QVd(GB;aT6[S[X.fAD2P14f
6Y^babIb8R2.<8a78a?:.[#+>KXD,K[14]])-7K<N_3X1d\8\IaV5_R5U?F8L00^
/#[b-fY7GGV?=29c]0:)43)(GcNa5dcdfW.Ad0.SD=9AC<e1>&P1IY#73>>)MD:W
1a5LQU8J#X)49fSP,3^D4XI\?4EaU1fQ-K7(PQCN20]gdFX/-9_0\275/M4-(JD)
HQ;SCV.5CQ=T1(#=(E(@K52L^0+93+RD<MP0JB6-OSf[K931\]X1&99V^J06W^-?
7PLNdIF=C3G(_bZ91(G:9eELN=(TN//OFK5/\I.>dcb.+<7eOAX=[#<740U=KCG\
O/YgL3&7ce=?=>ZK,_\7W/64,5O/L;c>0KJ8,97[LT1\V-H#Vc@HA</I\(L:A-FM
)(H8.4FB6_C=RDNQT1X?AG@4d;I#aHcPb]Y[feFH+://aBafCPN@6=,>5bf^##.^
WN3PJCOI9fbg:9f^>@1)K\ARF>R]B4O#]=^e,DTf)b@fU>[H@A,;f>BYR,WWM)G-
ac,\;9N]/<X:QD1cFC[<cgUETH+.SSPEG&03gUF[8,D()_J35I.(aYI=-T8\@]HS
dfa]1PH83ATVN^aB6R0D=Gg4E^^/A=,)(03DZI34>4OUNU@e8S)QQ/Tb:AA?b086
d5\B:8bCbYQNC6PDNZ0Y:\BCB,.WIRWEdTCfaR-#U]LaK&L>V@FNHCSC+_FCg7.d
<G-;8b:dHc?C2Tf/34e<c[HGM5PL.EM:LDQ\.B/==/bg+bH2,3ZR>=TKULJ,5c#X
5TA97Qd?Y]O=G_D,,ZT_NUQ/333d+f-#<0^eSLRZ03TB9.D2,7+2ga+5Xc2TU5:,
d6f3X?^SUIYIW33<8OREd-[@/C6SZE+WY>(&A0AQNT5L86(LS&4B-3V+,X8=N\:K
PaWFU@)(JFXFN\aV0QM78+=4^dgQRb1e@P?DYP2-BQ&?&#@VeF>BVL)XAZ,O-Q.F
9b#?QM4R,++eG=eb<.C-Wgf3cPSQI/9d6-?LgC/03eMKaQ:MY.L[2YS^OBST0)3F
fbH7\7(/8gc,,]X-4<R.f,:LR9[+A,3V:T\?Y#=3<=d&=QWc3AW#+E_5Kf8_cde-
/J078Y3<UCP>1,T^6/,1X=W@-Ng1>G[9O/f7bB,WO/[e1&S;N_]N>8HC.(&F2M9L
5PE)QR;4H8d;4</5A&4Lg:)7\c]=/aC7,@HMOG4Q>&RL66f]:EV-2U?9:GSFCcA9
B=EQ;364>PLG?R8e2#\+K?\:Ma:^]^GXX&G7JC:Z<G8ZFg<2QB6LF[.-P#PEBSeW
1GU^BVVE&#6U)IV3#N2QaCM4H0RNgO[T^&eR=>U]VDOGW:?Q?<_5;70Dd-]&f1/O
)5:>2C7>XFXD]=;/)HMO=2/,CW5aAf9CK\8fZ+-[6ZCc<IY<#VRZbB)gKCNAKV_O
+9J#;+;(BAU+;?&#E(:Q/2FU?EGg1fQcTX3Ef^(SNV5:/c[0eJMCVAcA<Ua?0IMZ
ZS2U\Z0Y@K[(_DYV#_X>E<HbD?SX.@:Xe3/6T8Zb0>2YF<?PX84b0D.;bd>bZPM#
QHZ[UV,KP)f72g@9)?B:0Dgg,Ea[RUW=LLYQ96K)]2?4ab[+:.EJ<I3X>[BdZ55:
6Y)_K#JK8?SK:Xce5UM-aIgXS7)K^>8G\:,Ed>egNI=QgKIP&VgHZ:7<LG_<X/4/
@DN&DW^B:OX4_2^ATE(PNWV[6/,Te^9_9^,M>Y@]6UH>.>5NT8AU+JZ1P,[;3B5>
Y.T>,+7H<7\A:SI@<V>]K(A1S6\S6DU^:](MI0@\[51Bc4XJ=-_26[#FO<;G7ZVE
Y0?=TJ@c#P1S8<9K1Z8V(+a\d@^4([UfEd3BB8(b#47@(IUR:fK;U7HBJHE<f1)-
YR(8=9ec.+;[_7-V#9Q589_\DNEJL(J-.[2A+L=?d[[D@2e8C5872O^+E#IUSR_N
U+3RM^KIa=KL.E4JK#5/T1J?Y]6@8baM89WFVE[bHG48UXR&;:2I@N?=IBFKTI-f
;XB5509.LS#B#B09af6A(._UTgWLd2M4/aTTR,JVHc??aTV2=0dPL20_O+c/?0VU
IVJ.XG:8[J@WHW=>?aU>&\>0?&767GCTec)[R=@Ob(BdX/a:OVXF,\/A=eV@;N>F
QH5&;1e=LbP\NSK?J,U)=ZgRIP_ZI?/I+XKM7ea&,ObNeV2(7bG+8&VT7=@IK?7S
Re,L[-)L1Eg.0c8D8T+FK+5^&HT7YfU.E7;;1KcbBeDTeJgV>UB,0B#8TB@&F(57
VT7\gfaHeAeA>70SO@ec\W</+A_GT^BcRAA_f?b;N\>IfP\(BZL;@]Y6-TI03[I#
R9GXPYfa=aI1Pg1^&XOeO7D#2-?Q&&K>_B4Ld^Ic8\WI>[CVV:(:V\\H>Y:^^-M[
?W;8^1d,.a\.]b-\X\Vf<\gX;<RM@+N/EB@gW5@Z_KWCG\X/2e)a/,/;+WKM7GV7
0A.g.bD@I20MKc#9071&?e(.4+G)1=.Xf_RWbRg)B=J/M=ZKW-e)ME^N0NFD_;3-
Cf+]7:;Q?W<^W4=Tdcb8_Ed182U1<Y_d]eF21OJ,5<1ENg]+;8QM60O5#J_JaHG7
B+N3+ITB,-&]>V4&gE]A?]e1KU-N6JEC8gV)4gH0GXV<Y=?=Z^IJ&/R&ETHVI[LV
6=>aOUTe(R,:fVUS5RYD:.:+:)E[f#_7@P82WD:]bDM6_IJaaS&Ig.H)KBQV/87U
#PPVF-<\T/9:?B]-AW1XD^>2&4@4E(Y-]O\PaJD,J)<B?fMOWQ<8;g0,8JV<4&XO
R#3f96bE@]:)WY\OW;.+GJ]a2JB=PBNBX[2KD-af@NNF;N.cEBJIe)f/\W4CUS90
_2M<E\Q?V#:f3d]2R:\KF[:_:fI:RbGe\^@6HMJ1<MC),=V(>WUTe?MUNV>756TC
[EKcJ87F=2\7Ag4HcgB.d0H9;X(RO\X(8316YS:UPR0VUTR6Cf7gf/QW@)],B#@g
T+d6MU6O23..;YBAT:Aba-4LD,#QEIN5MM]?cdKLNa8\QJgW9)gGV]7;(O/P?:(C
EIfY;5<>e^>T3A(LJNV](gb+ZSa2SXD00A(+Z.d=3O/C<[dBag&E>dJ+AMM#_e-R
CLffVOQ:&M+SP,e7:>g1DbgcRH2f&LL^,e7B\Z;Q2+YFG0N__d,M+8:)5K1;-RQ)
KXg[NO3/#&dfGFGC@6Nb:L;T&>A/e.)+BAb(gB;IJ6/FFGV=aU:Ibd7GaX(/8b)#
#:X\#EIBga]LS\YF&Bed)64]0Z&=d6:RH:GP\7EERN,57<DWIK;MWQCG4E(1gZ55
GC6B71+>F;0_U<5WWB^(+WBDA4A-gX/MdI4ZCE&,5G__Z9=6H+/IT1&50GA#>?Pb
&7=I9bCO?V&(&+bBcSggJ4ABc>bCePd/T:#:Xba8K.g=I]3H;3G^(V703SH:?eDE
<7[bY?3d_E,E([dIX=RC@AeH9=52TNFZ_eg<J67T54]6RU?NfOD3I=,]NF2.PDfb
Wd]eCY^EYP2D8@QV;fd:;D9(<K#IO159.(_cN/U[f9]3a:6C+,(Z;@a;aVA:@7&3
WQG^=BWa-5EOMYI\13@VcL2a?O7Z+M#\M1<TB)D&8)Ua,)79/cfc2^HV6=-U]L?N
CR[e:.CBA&GQ5@<=McA(^/f4AZ\eI6B8V@JTU_./PR)PKGWQ8<O11[fNF[TgN2_0
Bb5>Y+IO/2<+T-T1_QDFM#6bN6Hd0Nc7^YTPA(5IBH#3.?\dTaH-Q;A:Gc&J0WPW
TC;MLN2T>QN>S_ILT+^<T3<[=8[^Ye[.\a->+O\V2F[P&>gB=FQdE.fR;O#VgZ.g
6CJJEGN\:Y(0JfG7?08^Og0TH0<>e@HMIgGc5.BK+G8,=Qf:X>K?Of<(BSgUMcR1
(+H,#e#G1[f&^OQH<@8.a_gP?Vb@K4>g&(ATV0#JUcW8>/^]YD0+1VNJUZT&(a>V
:G0VB@.6\,WHe4MCE_HOf-&DQ-O_1f7#(YZ7O5?8cWKJgdaa3-M(bQ829gCZR#U-
MOVBZYID;_6cH+N_R;8f]24Cg_G7a2A7\,Lg=RIBeP9.-\M-\=);g(?S[3<0\4\:
d6Kg)Ue-N[-2<8/G.6]VNRT_JI1+P.f]7MCCS#W91M88RJ<N>4Oc.WbW5AAJ8=UX
O[=].;e3;aEM.J[/.ZFHRAUK)K#@]@Ea8>P^L>53dc3YeCBC<COQC^81?XIE[FC[
7BG(AE=(_C5W<dAeGR^a#P=Wc96C/^aDWZMI8^HNBC(7c(8J8AeLeBOcF:G:29B7
]5-HObUf6-BcIN/^Y;=TaBL(dZYe7S&Y[P2_-_&&;YG,:f[=-PY[B0Y:1SaUFIEJ
d)^C_DRbK5\3Ge0MM0eUO/AUHC6SK>\/&/>-<<d]48f9R7bJ.3V]HDLdF8KI,J8D
:VG)W+d7D>g8K(Y5e,Ggc,cHUT;ZG1,=1/130f8J:e>:JJOb]ge8UIQ<9cge37JH
<A7c]bFVIN/:e/),-9>#LBSeT@a;K[PG-HNA^7[PgUJ90..0L+A8&;E=,3@>aV;4
HC5;DF5AA;O5_g3QeV:7)T(,O.T=LWW)39M:IGCS3/=YgZ8,M)fJ[._C(^;@US>0
c-4<8L#FTfLND:WcOfPI_3TW=:#59X2B]SIcR;&+6LEQDB&&\=5X-d0B9W-LNDNf
IRU0c7/:[eST160a\a=@)aFXIJ;Ydc@&H&e?N3A_:G[[e-fI2<BB(+Y]H0b4d64g
A[IQ,-T#AJQ_OV>4Ng^Of,_cO.#b8JRM7<e=5a0CK9b&5]EG>^9#1W(:a6CQQ-L;
Jd0Q)-XV=A>#3ZKI-+0L5ef.(aH\:TH.9;Sf0@1#8;F^d;EJI+DHA.^eB-5eS48&
7^))JdbDR0b\V1/_8f41Je/S5A2J#9?LPNUF6Y#G<1,d&P<GJXfZRA@6[>#AcB+N
)^YJ4,EKMOfNF>Mc6Y2(^&IeWZaf),=2ZD+9:S\TRaSBcK4+LGg2f09A=+X6@,(7
Vf;3;30Eb.Rg7<S9:XL1\N-:f-]C)BYDVFUFL:5N4J)],)&&g3/7@DZg;Xg4aPBN
B0@6H-Vg5a/B_e(3UA(\\IEfQRf\GI3@L]>2OeG&D[c)Y9IcF&a/L@JO[&8E6;BM
@DX)MC(3:cN;c5Lg:QHe:RSd.V<2;TM]M-)&Ca/G)QVEBg/c@AaTae7f6#5HRa(D
#9PU:4D9Y2(/5;4?+SbCW&UIcb<#XcWMXN2NQIL=HX&C:+[);GKe-@HE2@g,a5S+
c9f:dbM>)V=>,c<45g7J6KW8+b_&I42D_CF..0-LO&2)DM/GA,WD[S=(fP@#RR+#
f#D]:1#7SBQZ7@5]86dH8@dT1-F9/>;>X&;c2^9_?W.Sg+-XZ4DRG/HH86CMM<4C
?VX&Tf<+c.U9N9ZM;a;19Y:gB5CG@;BTHJV+&B;^M3XJD1UbP=d&AJ(NT8YY?Z^S
K2GBd?1bDY?&/4?7YGE)aVO(d/PB---ZGYSBK;fU_MQ@63Z;KG5E(G2XX4?dO.9:
HJ#QOaVGT2#>e4E8b<B;eW,WEL\f=N\YTFX5/Ob3P&+OaR\?&I<M?H.DED^gg-@D
W\(E?E?_M3T>._K?XbW5BdC+\^GYCMUN(fe:^LU(IMU5Ya\IA.7Ga9H^MUgENH^Z
-:Q@7@O063=?53VJIVE/Xb1<5WFUW9<ZGaW-OTB,a1\MDXYXEVVTTA;S,eE+^:La
WTMS_EWE=O7g=-4Id\B.O6g]O+U=E0C=:9cfQTU)3AMY5EgVTOd&e4KOC.1UHKe8
?ZaBV9E#W#I1)V(d0V_]C4:Z3])65;<4;31Z0SOOGR++ag0f,L#Wd5G+f9B6&\RY
-7\HGX<.8ULSX3K0N&/VOK[[3A#X(-TK9(T:Z3,;-7e#fB(X&1c5[C]1X4=Z=H8W
+N__2HUDP]Sg(d2>8GRJ:Y=f[G(QX?adUG)f&>+Kgga]JZ;Y</Q,,2?J]8KS&D]M
+8J4(8^.2O)BVPM:>?_V^GBX7LQVRYQG8SX86LA\[fa+Z@de_IM.],Q,e:cTG)(G
Q<E:R=.XF?ZY\OIMBW92LM:e2aT?Z#-@M2;3(R=6I8Je07UOP(X8V=NZ1Ib?TCM<
XQ?XUeG92MgV(4MfcFc(bN4WYJaVAdb#eA;3P_(1QAe=E0Ubb)ge&.1_9Kc16<.M
@F7#C5Q&,(0QW\CK9_JFPaJ=X_Wf5;La3)-B3SI51;YE]WX,(eMcg<5]fZB+^64R
,OcT4#7D+(];;4I6>X#/&ULO>B:3/Be,;FY_,8WB]]D&/]X(E3b3W#^XV1-5DMd=
>Q.K]]9<SNR94Za=Z04a_ORVe5^PS((X[[19UQ95G:YR95KV=J-fJ_>.cH4HcHQ9
\c>TcbJ064-WIFT;:b<FF02D(8fdEG,3=YM93/gE(:NeA/@:f&A6VZJ3TQ&BUC[:
L>@9b-#V7X/\QBa@TaWQ4[EI\PaJ]f5df#(8P1_++8K[]OZ]9_;Xf3)]>+BKI+C1
2bR;6L0=e\CLT4087F+T2D_O+A:ERG(GI6fXWb=F-(O2c\RFTWJBO-b]QC-OVW[>
D=NA04>(;7&SDI+E,W5X?Ff\=8:WA7-.5MH/9Y:A=K7I5JNbI(LWHe3f<Y5;be#N
bZI6F89TP(OfDTU1;(+6Q5,Y0Y/CE89U.6\AP67@00?ac::0XRaF.QF5])X9b3[K
/T_,LG=eE:)M^gS(G.(#V80QPdZDO+62&c1</)ag4:^>P3TSJ&R?]Q5<dJGT)=aA
,EA/)Qf29C3UWX0bc-S]8#^M00^9BDc]fB1\RU7]c^+afe0[F,>+Wa2:]8)6(,8/
MIBYea>:MTA.49Vg1;DQ&E2#BfP&#@<fFUN[EQ.YPe/Wb_c]2&7<44N<-^fc@>I8
8EG45]MgbM)T:JK2SO_K-3.<Wf5\JdO_NV3@3E;8b5:?QKB9O=e1c^5O>0<9Y_f)
U>eGV#I<(7CS7B<6)RCH3cZd&723LNYVaXX9<XC=(J=<&/LJ0B^N,]E;IZ2V6TJ+
?CCZI98GZ1^54Y/V=85TOAN_U?4f@USREQ3U3Y+#Eg.F+?0N/@7&fW)D/?>c?8]\
\>aG2#CgC>)PVV=R3MDFN#24^5g:W&bQ6T5@a04;_g;QXaLSM(>M0Va;Y/_U#]7?
f1S^W[M\LE2PT&C&V2>f.13[\>(0-R[Q_KFH4S\BUG1>XG;OUFTFZHCF8P?78(6Z
4@6NbG\N6e^0^g.0<3VKNcbPaKB\=;4^Q=P7DBF\J7XLNQ=JeJD#R/<UQ67&ab3[
\-]d<UQ6;ZYNCPCSMM3JHZ(GaDZP\\WaX^)XL5dKeL&Se)O88D#=C;\417R^LBXJ
.[5Q9&8fdUK2gcJ=]a=e8;4#9[@dP=Ne^AH.IdBK:K71W9:f^V2M#QDH@J)ON4MH
WG/UR;SB,\Q_U<3.4;E2GXb@\:LA1)-<T4?6>#EQ>3e1B:]B8Y7c\c8Q5QPJ7feY
CL\JMYE5E=eGM5DD#_,5J-geUCgVUbe3N/gY9gV#Zg<)PE&8[S#DUI[2A5_D<?78
[Bf5S..Ka2IX_:9d8B#[b2bDI8c6[TZQ:-Ag2T-\T#b3?IZS1;Y,^I1#?B[ZHBdU
ZJ_WCKK>D2NX&KYBf0HN=6GMC<1@^_gP2R=VS4=+Z]B6)^;fe6(N8#=FBY#\\:,d
_SEQ5:OO9:S/QO<H;C:\C.b;,>d4Y[^0^X/L2T5DZ6e\I5/.-Tf\\)e12Y4MSV>a
6;J+&KcaOPO+Bd3;bE(d0Y5eQR^XX<7(2Ld]4ZdLc/fE@=G8Ub)]I(d^HT3Y39=5
?92ZY0Q-d&NO@GNC[<X=.20P+D[5VCS5EdL]gO;dRV)&L.Nccf#G4PRQCUJV#:aP
2?(feP2][IDOQf,b[J]M1,Q+TZ9QR-^W0CJXOgVF_;3I)TKW6_0CD(O[1^F?M/VD
^cRY(W@IFgJQ1M6MR/HA[Y&dP4b\N/H0F#/H<ZII[=:U\KY78\eW9O6E(H4[N+U2
GRf-.ZB[FE;>;D_CZ0S,^5g@+T4Q@W>ZV_^eU3+>KgXcY]X-HF;XU;@]F-<aEB<1
\4M#QT6g21O&>V6OU:Y-D1).8SPZW<.gLf()g]J&5V-e=EGaME<8H(A0@58[UcN<
(:MY05+M5\OcO_7EGJM9dY9.J[J><7FET)WNJfB_C3J(K8D:/^^5?6:#@GUPKA/G
M_NMVEDYHDH5Wd77P;M9</?1(5?YX)J>^_)#c7.&-AJV[Q>DXfIEI2;H@_1Ub/dQ
#&@?BL8(fEX;^_CGTd@6TMV#F&e;Vdc)^P3DNeJ3^J0VQcZ/L>,0]f[J_4AY_K/<
&:HZH+QgU=_R<bYNK==[[,^b=BB)(2YQJI/]>[)W(6UK)K<][86c.5\E9aHe<?;W
:JQ5\3K&T=@Xde9Z]+0F6B,ATfG#;13OFUE-2=)OX?g(W>Y:44,EK&LAY#FAD4[F
ZeWcU<J8BMQd/25SN1/=GX;7K)V-.+1=_J\&Y^WJDg]^R9ON.6H1f[UIB_7M_+A_
[TS&RZLEB++gU3acZS4SA2bXBS36c\g:?=S9,F#T>JX+3STL^5UE8?\_afQ]K+<O
BZLg[<AVddN#1HW0QVGgB67D#e8:JTK]#F<CcY8O(=c&/KX9I=Q4d0^eT7aKVO92
-#RgcQ=4CFNOe7PMJ>[OYM1VVB-5_HP>)(&0WH\WKDa)Q7O#+#ML+^5>]6(2Da1V
=,Vg92F^EeKG3QWT.+^g-4V_9Y2RA\P\J@Q_(FQUVSD7]0fQF-(:P?RM;^Re+2\e
NA4S1&cFAD&Wd1:HLLT1(/ef/6VQ-N:L>b-[/TG/7-<^)D]30BD@Ae0Id8;?QKeb
,HNV)J\;Oc1L[)gg>XYN0]>Y>XEe_EM[TR@<1JA_OW.=TCcM=\2)d>cS<>9Z8DJ[
S?-.=_cW@UA6:/6f-V#--,-2_M^WW3.#<@R-FZZK]<XgDLLGf1Z=Ge/fEZ&];5.B
12J>ccU-G95H4IF+./D;^;29XP+9b#:#R36XA/0?f\(HUI02e-@5e=,<:CO6MT6U
Rg:X&S4>+dI>L)>;6[JIXYOU7M;_=D.4gXC-6J2dM+_eUKdV919T;])<,a;D8X5g
ACZ2K7ec10D@(B6@8/GM,[M=Y<4=>\bcgC6(bB/_KP^gF-g]<J9E#abV?9geU&/8
eAQ9b&(HW)JQR]T>Z5Z^eDQOY;TA+O7+bS_7SGQM#^\.>QVC-Z3U6U@dS@&9a(6?
g_dT:)b.F<NcYHAYc-5SE,&&A5(1OTOE?fgFGJ\:OQ&77?MPQHUI@U7B;XY2+4S8
A?K<V#UM)F?U<W</,FB^5U7WUXU->XfaRP-5G^S+<B(<\W(U\8BA4B[SeKS[EJY#
,;OabZ2SK9<-^Y@GKb1.7]SL31B&;:dL?ASH7Y[B[/\YQSO?NTG-1.<Z@>HNGJf/
9&O_/T>b]2gSF10RcaTZcA7eH_,^_NdL0,dZW,OZ17Z,N[8KYNdDcV8YOE;T,@Sg
[M[T\Ve4YS:1E-[b+\11A=A6BDS;cSSAW+4;8ZZ.08PG@>e(Fd\fT9E)&>D.F/)X
+<H#?&F2+7WS9)950Y\U73R6,X4\;P?#.U=d\68VSO?\&6+6ED[V,3<<d\/@<#\/
L<e,@Q#CWe[Pb)SDPV3:5Dg#0(@ea^g?ZZ=F80V@)3?SEa&.4ZXd4X\OX3aEIPb>
@+P[Y&A;FKZR\&aSG+fZICc(;;RD+5:O(dY4H9474.SZXV5_YY-9YM.f??DJSa+T
XE6aL0G@E/\U(?I&e,DL[;03XX__R9?2Q.5J4;Y]2K;<7]-X;S&FFX;S-a636c2b
<9J<:XeQ,dcJFBZcgc2^28V-YE-42/AZWQYBO[3]KDV-?Y1^N>(V-)e.3W41#17I
,[(WX\fF)QKPXZ;H&f#H7L=C,eJ9(6[.\H2NY8bO(+O@(JOKPJV[0aQ;7.34I5FJ
7@fIV)ZT,8;B^&@^[)\WD;6YN]PQJdI=4e\dBYFf#AIbW[U](dSf7+:YG(TUa^K\
d9ZX#N1PIA8],TB#Q\f+R_@7U9DTK)0@d+];S,#MbL_fGG=07S<)9)bNfbY2#KKL
T/b1L[=SG+>-]HE-f\:1PR\5cM^Y>HgfIe8;];&AD=ATYO.dIKJMMM?X-VI#S936
38>FC3fHK(OZAUW#OO=NB=a>^MI=.TU]<d6-M?A&OWEF;-MJMWQ@e9,(L_1[Y3,.
dfXgfY;HbdDIA)-VYWbB1G:P@#f9+c&P4K<4@3:=RaLf@]HH/=NT1)MM\7QN88SV
61XWG]D=/R+feM5A00X.5I11XQLUGIH8\H9c)3K&DQ;BS@DTV/45MPLQ9X5A^aD9
SgIb1DfA5F3=,U-;TI1-<&K.4RSe5XG)I[?JMA^d])7)34Q>0I3T&^#_B536]f0P
O6Y_SZf_HGBK]BB09d@a#T6?F.).UQ@g];^cdUb,+1YQY]-Y_J&,XF0&5WM>FHQC
.DU(=W/&IGg/&gLZ@X/5e<@;JQ+>?X,BADK6.-&WI^_LX@eb,1Ve10d#<J5AZQ>_
K:A.)R92KU\cR-:76MK=03d=d)(bJWb(O88+=3S(#FDR^45[1/[Of^;[@B1_ZJB,
Wa5Ab3[E]Z2-QfD2cPEJPBY:?[2Ue87.86C-&<,R)I+.H0^+X/./?AF/UIOEMPRZ
[g=+WJ[eP],HDM0U\C/:(@USE,1,-&LIbQ^>0^0/8RbeX+HG:f>fF_JY8T1Y-3/Y
=L8QF[DAXH]NR\5]QF/=PTPBH.bRNbY3J,0.FI6Y?d@DU[Oee]U.dI8dc3[)&3:J
F(&[-56\80Q_g8RMA+-27_6/I#<[gH_BWf17gSGdbaO)<b9d<1_QgU(#.\QK<O&F
Q36KaK+F@dWQ,S:Of:X@^2E^4^SK+C7/>MVJ-d=O\E?dQEb.^_)6O[fbX;?01@.0
;1@16<[5VRP>g<.3D&?P,RLL&]25:cJ?DVBRPPY.N4\=dAE&YZ;9c</5W_dZ=3R?
4/Y=UULZQ#[UaPT+/HA-4G1YXI(f_IA:4BV#2)gE\G4603JA=T#]X?2Q^T2GeBA/
]\)_D)3P\B9O[)#-^95BG7+0R-LW#@6XF3_FG(I^=GR.;WJKf;;66f7dVCX0R?G2
WB^V40Pf^F#XZY5Q?C1,Ggb#918XX-e)Fg:/LeBb_Z_Y1P.MAGF=BK#)0S>)XGUP
)W5,PV^3AGO/4M=;c+/O9R+0a?S&)Q58+\-H4O1-8a:CVSJb-3d=D4H@Egc6[I7^
f\<LL?;L^]NGJURJ0YIQ?b[K2ZMV9?c@D&T;62a(LAUL.a@JFXeI/J:>T,MRcFcO
7^EJ_IcLQ5OdO.TaFPU[S0W0;A+VXG3CYTgBMYf1YYN5Z(CZC5+f(32B?-SfD.B^
,_7cBFK03-/gfHI+F#&7[-2F5ac16<]fR^N276HdW5C?K)f-047#S&Y&(YQKT.OB
M6W#8;WX6<MgT=SafYG@496[V-0,D?+5QZFJO)<[R,Q;+J@\5f2=93-#fZT8U(DP
4T\H]6T8Z/+5(Z&5NVY,H&LZBdLF33CZ8f?MIGS.b0MNB4LSO#BL,;MbQge(_2W^
7:5Id<F2<N=>.72+6e5UF0AM+\\RXG,_T,DeH:Q@aXgO2EE@;/c2OGE4Xfe@HD@G
YeR??&/(17gWBaTVJS1BZYF&X<Q(d?CIeR=#=,^=,7d(d17d.6Na^AVDX=0&gG>A
]?_B;F6S7QDJ9CT2Q[_Va)+RP\B#]^1_CcEA-QMg1O.6Y.WO5EDD^5e(<M8FX#FK
0aS0#]NODE5RF2ZC\02P)DHL<-.Ag-;F&a@J+eI@G.BGQD=OcHe)S#8fTDE3,82M
WM7&\A;H8c(MNR/Hcg&/+b3(^c#-B..//-EVfX_Q2U5J:;8N/5=.<=YFHaGbA^2D
:3..7PQFFe(;QZ<9^2]8a0YJ2VdCN39RL:=H8^IIYI/]2AbE-&/QFXR06&QSbS<=
DefCG=13f-P=)b3M/g9JTV9&?gC5)7UR[:dKIDILgTcK/C#2?BC4bL.I<b-_PaVB
8OZ.FdOXX=A[S0FD]9#/7eR]P(.MVZcF\0c9MPCbKcW3#YKJQ4T2(CB#8QDKgE^@
P6YNFF00K#VA;MR-HCXb4-abMdMPNc=6BNR4^><G2:[5c,FU0Naa[dc(D5V@O<)C
;0BR(8aA6&eK8FJ^:d-VFB+TTI5F]ZZ3BZ-QFYSTa@F?^/e1EMCS>,4/>)9#HZ9P
W=RU:4MU1aZJCNXe3=2Y\25HF\aC>c4+d(>AOCM&_#G@MD<feJTB=6Kd0FSS2.We
4:G@B\\#]<[Lg>_5)T5[?_b@<3d\=3L[>3\eJ9fZ8-a8IU)cUBbd^U3PdS&d0JcZ
5)A&MgO>IcJ:(I8\:fe/4_J&764BWP9?PQe0=DE,Pa30M_6B=74MTTID<B(Oe@E5
U2eQ^IBOcCMEPD3Q6DM:F4V?Qe0L#WLcI=CV0OWWD?EO1K#G\,E;2[Rc)[AH[@[;
:2AeSb22)TZR77>].T<WK[2SZU\V]2Y12E<eJ2MFK4a#\]L:a#5CNa^GBP=K\&6+
6c&;g3.-M0TTdYA1Ac_VLc3X-FAVSZ_1Td69fZJIM,VKN5](eIF<7TKQ3:bV7-<[
bG-5Q(98cE3T47\@T(;3JO&(8<)c[>5[GB1_g\+N&0E6UW[\@Xfd6\&=_ME7MM<K
Wa:e9M5JO@3-S-4F.EA1.@gUg+HY#ZPIJ2^VV9,#(1W8Xf@MP#JHdU]fCEC:,3_Y
SR)76TNAc=d7/,:#W&HG?&Q^MBa5#W@RFYB6:<-=TE.gbZE(QB:XP:>?,)6DOe27
HNI,)R?H330f9@IT+PMDEC/D:3BV@BaUR2UK1#NBfg1b=I#7<8XF\284JGL..P6C
[^U&DfD?bfX6UWR7)RC,)KE:]95&]=Ie.d[QT,3X0#)O/V[LXR]:,fV,0KHN?7CO
c:U8df)#gUOIW2N&9QCf#g4OD4\e.a;4dQ4gU(27<dW3,?9D04-7eT2-,K(Z.?<)
T#R1HCe0DJ&]\+Ie6EHR0YfS-L9.+X/&?AG@7NJ@FK_S[SJaGBX[O)+XIK+@U3b+
f^[S\c-Q\1&g5_\>RN;(V)LN(0.[G4W#;CN0RgLIOQ4V^0ea<=(M[IM.F:ANK8d@
+LFPZDd/LOZ5BQ/&E0MURVP8GFc^Y?UP+?Od1Z8E>CeR8UUSAc(8L<XdcBK/&8Df
WKHRN,Z4;CB-R,@MUBI)>C4,0(c)TZ(:T)@1[6RXX[LT=^\fg?.W0)LT;&+1E^0C
R/2RgAJF[AfGgA=O6d@#C.X5]g&CbY0NQN+N/HNc>D,2C):458C++X?0D=e_?3IB
&FC4-D=<W.XXM^IYWC4;:A0d_0\g:NET1<:0X(5;,WI8d=b:O8C[:ZB8]L_N/U6I
GX7].Z;J0RNP@=#-(#;@0.5JaQCQ5FdX0.Q:9_HJ/?c:-#Sd-gP?;1?)&aJIcfB.
J-Da@40O#(N,?>H6E9;0/IGE#R<4#+SaJ[.F9:/434]4FQ)]TK47d:SBQRcg\eef
C6;J4#C9H-Y&bc&<0CQbcA9=1.(Ac47>3Sa[CDQ1/ZdZ,4N;#DL[.6NZIYEeY#P:
RbTGQcaDe_093UYd\;61S88@(UK<J\ES-bAG/[L_[\a^ebD4/Wbg,(9bP)PbORWS
BU+#AJ5:ABLe:JA01T[#@IcVcbIa)J]J0<eU>\6U64Q7TWN\VV;]LFA@J@#WZ^Y,
/UV?2H#<+ET18^[A29X8YR.fE5(:BQ2@V/cQRKDfD,4\=bM#A\UBN;I4VA<fEI1S
d-/O&()e&fBET<;JE[cQZc:(;?daGWfU:U1S2?-IG.XJ+;?_#QKNeIYgeZ.):]D@
Q1ODE6^\LgXZZSH7@\[Dd>ZZeQO6@9.IC6g>HJ4K_bPHgSd95U6@VZfC+O^6:b?;
1Z<S/>IP6aRUUV/R1-JSHPeN?3[0dM&N+&g6W3fK2cX@@H+/V8]=4&,FFM^B=)Qf
J1)W629eRTN<3b<>+VB+GKYdTJIc3:e_a=KKJB637#KNRSE3cf3(X+,V4MMPSEb[
>ccXO60dFDdT3FIPN2M-gM9\^CNM@3VJA?KFS[:1TSc,5(cO3BZd0?UQEb^PM,J_
PJfEXO8c/1GKf0Kef>P?(TUdZ74Ed;g;)(=MM#,ZFJMd7,1302T1:V:K35AUgC_Y
_1R:I974E;C(OZMD,T(SR5&C7PV@(A1W2VG3VdD)?__>0A#4^b]O0\FJJTF\=fP6
a+4g-V]AS;Xg_9^.A&-OA6M<4TCEA35+D:#QX9KgO]X--BM_JX0F&T@M0OT:YMfB
fGE0;Tg(:QXfUOSB39ZYU[+)C<QQ5TS_[R+L4DPEaDS<Z3dRY:5A)>@PUMDb[@?P
#ff.9Y0#K26f^TJ]]=IF^-617G.gX?LO6XB/B2Nc-5C<&BAL;?6T;)K,ES^X,W^H
:gd-H-[7FU/0([e,#]K9W^4J:[E64cHe81]@)cP)K)JUQ/QOB]]+FX)/JI8=D0BU
Q.Q,M:<8=<]-0cD:PK<eSM_[Z:>NV#,g(+Q6/SPU,-\<87+af\&)]50]BLF7\7a_
RL_d5(+&Vg\PdJgC1#dWN>N?VE[WRa#9HJe-Nf)C+YS^VJ0ZLH>V@aA=D>(M^=DP
;B3LZ,=HTb0]aDf-cF<b,ed,-DQ0>dN6c\2g/>]O;gd1/2]DPT-OS9GEX&U#89aV
K@]PMd#d^/[)U1ceNO[&SVR4V],5P>4HZ,Y]<S,SSaQVc\7AbP]&/+,\8>8]LWR&
OX.DLQ0SM)5N,9fD4=03f8f<e2_VZP&UP)O53);F#75RV,eC:@DC+?TfNBdP&8cd
VA3\\SQ1F7@,@C<C_:&5(T]-AeG)ZH5XI\[B>I=?&G@+.PVf:J:U4R<T:I,6T8P5
O@/6&2W>4EJWZ3P?RDG>(>92HZT5#?)NQ,FI\<&6<H&2YSJe(V+^XMTd&cX?K:4d
Pf,+9F-AJE^Jbf3K12Q9N,M\\R5cWJZOCUS9(XZ\RKcB#?D_^:EE]1:-gXd:S:DS
5)ee97J#>(9Q1?9YOF7FX_[SZ5gD&(PG\=VT(2..eCWPHRfP&_@TeHfaC:ZY6=2d
G@5=1F#8J#eBFEG6\_^aMS-&7P<T@[COY;I<.AG^^]JA0,gZV8ALTf;QJ3c2HO2O
gSWKfO^<M=TU]7OV#c/VgV.+)d#J+B-E2aCRN<FI)J_F84CeM8e#(\B8XQ2MQS6S
c[-03F-OCB8(^?d&-YPFHgc&D(A:#)F7^]f6@+MKbBaH[+[HUH^A4-5P#Y3<@gTa
-,6/?V+g6bbZN2WX-[QAO;TS.UDeKJ1Z_M4A>1,1Q(OYBY6+)<5U<IPWS;&.)EgB
\:0d23U\C/&<]7)H8.HHRAPSM2c:6]F#S1]UIGIZXeab@31e?=fc-RI3=(C@Qa2^
5I+f]^/3<e?gFM@E^C/PG3gOcVdTN]#UX/7,14Y3cRcNO3-Y^eWLL8eDRYJ\7>IH
S1H;HL4eP9BWE3-X59a6,2]@E20bOPKJ@Ke@c8E_d3<MVgZ,:(>3AB/1V?#_H;M2
H6PgOB,3>W(H3Oea>:8TDM(,AQS=MeS^3ZaP>544g/)>.7d<Oc&?0[>F?L(BM)GC
?b_63d[g@K2-A.ab;f5?-4D0#6#T)T[#S?Qg]If>LDRW.e9>A6gY1R3-WfDeM2=L
&c8V^9^eXH-;>g0W_NJH#Q[L&2KYT&L2O3FL<POf?UGWFKc9@CRfeYDLS@8d>&M0
98V6UBJS(>Uc<#f+Ac=QCI]P:OA9NKge_L<L6_+/V:c9YM;]Md])K_f,]X8bXa+T
U,[T,=N\VNY>-b(98fZL@#IEQ0D?25d<<-T):[L=VKW^/ca<APd8&=-7\SGCWZCJ
60(Z\72,+S^5EDVC9F/9B\JbO_&CgM@4B[J57]((=RXQE3:,RIP9F[WGgKTaYDfd
E7UXB.0b2D2Ea^)G3GF(H1IKDD+N>2cO6-<2S>+E<-BUeP)g<J+/[Of::0Mg)B2X
RXI+\9bS>J;5e.QbH;;/J=0ZLIH(<S1;^E2?D4+,OKATf+3AE93W\eccE8Lb7e#<
F+-75P6?H<-K3-[4PeZdU=QI_/;<gK[LCe34bB+d\BPK+#@LgYQ/88>1H_UCFCf#
PE[>g26=\BUMH[]b@=+7MR<)\gQ\>J,XLK1CH9H3ETT7A1.0IV4QQ)IM.f[cQN-]
0L4[bZWQ@aB0@YO#C&CcA_bfI)]WSIHJQ#,7XI<L+KSc(GA_;&c)==??G<HLLAQb
bFGH=fKH2=ZGXT@bT[HM4[LR/<3HaE:];OO>XL&9=2H?Vf00=UM_\AVH>P\VG<5^
9=BO]Y1ZCXKdJLT[/-9W,\UV38:fFaTDNE4X][O\U4I)U=EcQV0GT72IY.^f(3AD
-&4K(,X8aNRdEX31MRC0a(IVH6XZ_\]HeK=2BWN->L>B[7@cS.#XDU<3X=^gR,TU
S@f=A51\bQT_VT<O7)&4[7CCfB2(R?X>T;KbWd7R5[F/3<4P&-JYe=O-Z[OG/LeI
BQ+b)H@SNIBP,ONF[-.T=RPe_dFfS,KG@;ScB(=,a:N1_>.^3X0GP/VZ](3@V#^B
^X[80CR+cE,:bFQ1Q2b]deb@<V]2e5XL2dO5Y^0+M,gB.a^c1(<-FFIe>+OZ2++F
Be9J2TKd\<OY<J/f1WF<P3Xf]NKRgK;RS&D-;M@]:(LGD+W,T>J.S7fOILHg#-6U
A^S=K1TK#\/C=e^K(=H:<K9&bX&6,X?N(::B@Re9^-f4:YR+e:F?W(_.fCWQ40T-
&5UM/I/I=Vc1G3K1[ee=@dP>\D<7N4X8]/2=DRg7Cg;3cd\,7/A2/&0M0[a&88eG
FQd@9=Q5KK>XPaJa4.CObKH3d>??3QcOa04TD1/94J)NT/+dYU<A/]dKdJP4Y=BU
<9_F7UB_e638R,Sf-/CLZdH3C)FC,KJ;LB&W(:bPZ#FfI90UJ&F^U(61-3Pg=XV1
__F[aDV3A2^1L;cZeF=e=eZfX4=NC,09<^QK9KPb?EX[M+?4N\>2b;\U\N]6g8Ua
=#5,+>XETg#9QHg5^HW^;HR:3.RVD((BIWYcSXa7IbTA4Z;-6J2C-23LK+GXXLZC
_MaFd7XHJD).96?S>,6>7:)8NR,YEK_fIcO=.;_@JJ1-J&&d8SP(#ZCbG)5+Rf^E
B>9d#\^@+#bR78=;4DH,T@67cGRb7C/48&G#;Be<R/KRdDA?RV0ZA/>d/c3Me(I8
AaX325Ja/.3OS]&>#-8S@dAbQLFBb+0dc^9,.5[Z7KWE/>OY.-D+9F@62E>R/+e]
,T1b\D>c^LI9P45I2(/?X[-5d8_e^ASa88K5PTT?U-[H1[7V[fFG>6C&JgP/96>(
-W17>@,B@0TICQ#O(a8YdL3U4^P#XDc-#,]=[]T.aY,C,K.HV6]d<S\fM^e7#=NG
aP(gN>&JGD04b5FgVJ3J33D(728I41MG_.GH[=FAN0DEIDa,.dDAA8M(?[(_:.cM
JTAJKZ\A=,6IKRBTbEDBWOVOT-[DDI+dAKcO;12=LG9L)8+?)+(X;_+89S,DB\GK
/M4Q(aBTQ:#NRF\=C^gWSWdLBQGADDedZA8c+;Z-(c?W.d<3e5S+[Y<b])W-d.<-
POHCXTaNZEDb4BC;N7X@ecK3e[V[RM.GZA=M(?V@X&+5VLI;/CM[^BR_6B2P7aVO
ICZe11^f9K3)[(ZVI#Z,,:;1=&A9R1>d09e[.:M=&2<L-aTe4<dZK1Ug5Sa4Ac9,
DIWIO3L>3BD8DKeD:c\E(U(5I)PL6;ceeJ5c-@Q8X6K.f_b2VKF;2B+.C-d=e@H[
PPX&/NU,FbeZI=;N/^&LPI_2+@Be).MU[J)O?3ZOcS>F:OW[>5DbU@6U/5GW<(b/
4g.XHUXUHYGYX5W-V@5Q\CAQ3LM;f\g)d0S3T+7eJ)4TNd9_.eG<4(:1AELD(Z=c
-J);+4[^9J+-C<6+Nfa=Ye(Q:-4d(4F]eAXJZE_QLPQMT<Ya;IP6>DSV/\11N_Rf
2\e:0D992_2X_/U/K[;3]Z1<&6c>0T?&T/=6cRc-6HK^XYfHZ691Hd:T4Q[Pa/<3
H?9c9EdPDe567E64\W,C2M[b77GcL>f^VQb&G1O.J5?B7__O\AK9?XU_4>)bLQBA
5D(/0?]a5&J-_g?/e@NfPgIB=VSI]ZD[bb+=T=8])c09>#Ig#a6fEATHF&c+WSRW
Aa)>2I(cDPF\>GIg.Va]7f?8ID#O+6\3)K:4O,@484b;DbSQI>IY:E@9BHV197V9
8,,>MB_fJ(d4:fS:b2<f5WZXT?4.G&G1H3+=Q(VY>+)\g&a?LfU#4QN-D2-IBJ/d
@.2NYMACH4O=N-H/107)LLW#a\5b9>5L-3\R^^gL<:AO)9E9@XXKT=17a#&d0>CD
Q6d3>314-cUPL(>PPdUQ-YV9ga;[KM.cBXcDd,e6V)BQ#,X;.C_I[e>S,Y8d/d=<
C[bVA088\XNKG_g77T5^a48>AUBU#BgTE:&\M70d#f]Df9WJW4576+:8Y/cg_gR+
CP)D96RE4-8;+<f]H-32-/b\JdYFCU<(.cNT>&L&INY(.)7).I6Z.]2SKZY?c[Da
9R@\IKL0\>BB4V]QaY;.P4^4N7(M<@L;)9KU1M(6?DY?\NG7DVYEC(,=/Y3?HY)_
O9EOHY8\@@,P&W^7:L0HTJS]P4b9d)0b6UIGX?egC84X,1e-1+:9-M49<8FYM^bN
bcWRTUCEgb>YCCN<,E^C8bPOKTB5#&NBLO:>(/TD(4Pe?aGLY[TX&3@,V&QP-OZ5
PU1D3BfUQaNF:V#1cNc+_WPPVQ&VNgG4REG8c[]65Zcc?R1bH3G-EaYS<RdXga\;
S(bdQe4>M:N:Y[Q6(W;aJ6K7IIVOF=8&-ICN9A1I@(VIKDC4O(]cD0;F71;93>;&
B\L58.<V[NUc=AcU>2L961H_LD1cQc?[.)=Zc>Zd#EL9QJJPH__Qe..dG;bOdAg>
>_@4dYXXg#BY/3,XBg(5MEd?Hc[c)&;PS[aAKd2YW00IL([M7/.A3+>gO=AcOJ\d
R7)JfOB?RD^OgDd^;fgX)JQJ/JD@OXgfLZ7/g(@JPF86P;ZRY+6H#7^+KB2\#3.#
T.43]W65#^MLCLYWB;(I2/6\J5Qf@.RW^17MEI,\8A^DGfP_aZDCK\]^Ge\Cb?#6
0@K_UCB[3aef(5(>cJU:^@-D:<R>U]XH^OWT47EE2=]W85HO]cBLDfYWQH-0BYWO
a^[(L@TNPTE=[/B65c[f]dRW1U/D3KI@WdA<-1?7.GQ#/?;JOf?XW7F945+&],GZ
^X0He@8:IUCU01X?J12<00@5\VM/bAJg>Y&/G5(6_D2?AX_M_C)0LdB79JBdL<0Z
97++a/Q<a[+DbFcYA1@3+?PP].&AK9;]:ETgQ)LH:3d+RLZXF14N;V-I^<c?898#
)c0:,E(WBa<bcR6a&@MAgg5V:9]EYcOU9\3c>&8H3FK[_Yg/DDZf\a<.VeT^[WQP
g7Fdc>1^Y7J.H,1M<.<-4,J;@PS#(^\28&IF=EM26#fF@X(K+)CLOe9Y+-K&M2IC
T^/BA3WfY8bC.XO>,_-WfLLWDW)O2LRAJMLC@+=d4A,@f)CfXUZB+-C_]7TP1B1I
dO3>40)^QJ),S^bd9NY6&UVVb(O6=1N?;ZQBNW,[<U-/]#G_&fX/87C5CM.1D(0Z
MbRRV(2,>ePY2CSb6HVM)Xaf@C<3-KV+YdB\FD=?FPQ0U\J(.X[JG-P<<Q?.g\+]
6V1I:\4T\Y;E=QZ@E:B>3?7<M/A_O2=RZL0EbaZX4EJ:RDK,,AI7PHd-Lg6/LUMT
dg@?M]ee/U&+2Z&0Tb]a02#=A#Uf)>H3e&\4a)8XM[TR+CFLId\f5a,^]CcFDZMY
9g:eTZO5d.V\-(=IPF4Q]#_d#g9):PV702(OQW_3)AU+.gaG:(KfK0gO7[K_MX-6
FOVea4UT7YW^/83.>LU,2P_MNJ&2K<O-_\4bUESM7S\aTZa([K[?T^VT0aaEgB.c
X263Z\Mce@c9WYWC&eaQ(VJ_)^b6:+KQJ;L]=,097:?C@1aGD)D.bWQ7+AC;U9IJ
M-7@N=ePMN@,27BYfDR4MN,PNGFE^)-^Q;&3-PB=g?/Zg,Af@LTY,.]QQ]W+O:bA
(/D8QL6N4)9;,8<Z@QPg)#ZeQ=(,G0D(7P5<MOfC4TN5[D=f;3F</TGA@229@2T#
INJG0Z1X./A^\Nb5(:;#<1_<g#ReJ_KAN>/Gf-Ra[MP<V1A+R6(6HK?H7BaFTGc5
5;OKHGE5>T4N4]TUS#BQ5M[.TSBR>bQdXMD/[GXN@@J5EN@^\ZP1S2)V6.D05SH5
32UG&>&7G_OW#_?Z@Q[^U>0\P;/NS7.cXTe0:9BB=\8(K7B;bBGL)193EO26YRM,
BV.XC0KM19e^CPA<65+(63=DY)YgNQOTTQQd5\_LXIId-)\1D@60K)6(a9JT@4(Z
6R\S<d4]:RD,ZJ@7W\d..9S@B:O=OOb+5Q48C?3E=OaT/A>^ec8Z&P3ZJO^;&@e3
B+GOg[FX4D&D[K7AbL2@;[.L=4H<Q2A)Xe6YQb6RV?^#?]AIBBg86fS7ES6[YSA<
<.H0Ta.?>d338FaJT0GG0E\(X^XHVf=<2.]4ZTgbbP?60730[[C_?#TX@==N\O?8
147F<D9gUHVXGNZ>c96/eOP<57b4NZ+MNZM?WP@OWHZE#R2_HWL8A\ECS^70(OYV
YS@8I-BbMe9?A436&AWK\6b;>ZTC:e/g@(\/SE>48TSKH+7+(L]b:G^RZ7>[E67P
&;8LdK9_c(O=Qa/9^_cFdSD.;ILT.IP7Rd0R\5=Q&GFP,6TdF,ea:g6&RG-<W8@?
[0cI-/\aR4]HJ:_+.CQ:f421S^GP\=1;\1e@Hd-49Q6@(3LRce\]KPM-gB_fL\2b
<)a18g&IJcYN.:@&.+g4I=EFY>.Yf5eOJK;-DT)]25>5SYX4?b?eE8P&F>/f(Xa(
_LSP7Z)(UQ,eBUeHW8IQ)HFc)80eLBL&65eL1.2/_FRQP;55?N,;@9]\&#bZOA.3
e0FFI.52/KZ(69FLfD4GEb2aRfU]48\P-COT)EHH0aQ[4_\eXMGS\^Lc.-&CGYD4
_EP0Neg_[N<&(bS(2WHe(Jc3EN4=_[CbeUO5bX,9?-6Q.D(J#\fC(g0:6d\]1&CQ
HTC]KQVNATD:;9d[++I&7)Z<A=GI2JX:67.S151T\&,MO?=LNKQ\(e,[45Mg?7>N
+YSN2daYQ[@,O,@:?-1\;4b3a>#L_=F\:#+3[.(ScGVG]CH_=K)La\V=0;b]2Z#/
>5B[>&,S\:)L3US6WSRQ#A4>DIR8U.9B\JZP]V<]M^QLgEKS0W\cTT0Ld;]g:B?W
&eI+BRVX+.d)RN0JQ[g,U-A65N\WE;[8dbVN[XG;GP]QS?HVTUJYcUYbO/5->X@]
eQE<Q&;d5=e<D<eJXe)a8QBO@fZK9/]Z^(W-<]@ZM#^aEODAW8,ATXW\@I8X5JK_
aUYD-2ISB4YPJ&A6HDQ+@E2-OR(QA_=eH+;>;gEN/LF=>]Q5g2cT=YRBHV-#Z(>_
U/XZKU]+H<6\:R,GX3>a9]Ke&b28M_4TU+UCdY-W:4K@91/-4(\PNZ&#HES&>>UD
2d<AZ(+d;3?XY-eR<M096:aGR>DJAYC5IEUC0/C]=Z_HJJ/8#YA_<O\3,>YeAZH<
^f@8BJS=c;[T9)6>A+M8UHT;6>)b,>3Fc8V^1J:]U><<JG/@;>cN?6Og_=2T2-:1
V]:-EOB.IJ72-U20Yd.U&44^926gVb8cYH>SHFEdV66Lf,V#NOAKWDaf]76RB;:J
+>#I(8OH+SOJKD]fafT1?)&J==6W,dBV/8PI:L)58Q4QXX7E;97ECJdQ_]:_ZK(B
gC9g@UfMS.&?fIK\Pb\&GB;XQ8GZ1+F?>4N,HfVA[^(TS=2[=F[Y,NMCU4)@K)8b
D&0c:5W7(#cSTC1(2Y[RM;+/)F,SGZ((]^O<7-6EK0^]/31eBb(+/@a>:,Q->eE,
@;DBWS)QM-VA(SYb6(JbFS60=YO=?A6/;E_B]FQ;H9[.:gVF6#cZ-/01N-GUbcML
TaHC_E3^-LLFaI3KJ9&&7=7:DS3/N.aYN@C1?(.50VgKN>bMMC8]AcN1L;gAWVR&
-@;3O^O.+2^>B,:WfEZ>A56/G4,@LU;;BOP:5S3(f#.^0XgC:+OM28Z_O6#DK;dB
X]6[0c&1da4^XAXDPUMMGeM5&)8=J/W^^P:_Y]BRZ8a_I,I^FK_:&L==R9HdAZ,A
@O?dS8>[.OF]<4<6;=[0g>G<>,=?e)-?;:8E]D6Nf3eJ^I_6VWYReb8cN^ZFXNA:
];LWcF#c#)7UJV8e5IN/Z<cZgH5cA3+OFEMK@4/9)XDF55fQ=NU@ZMYO>5I-XST-
B+BG)8PM^N,NJ^B:HD(57b/3Q?@/:Z?eN&JUNJ(:26Y@eW;+\W5AQ:DG8<WK8aJV
06>6#=E,->(d[28bFd;42)D_LO_E7:Y2F>^c2VX^[Q@=GF^.#bL_MJ/ZC6P>@;.3
R-:Hde)S3Y\9G\T=RKbJ_OPE&\&S:RO3\,;;[V,,c^/NGDY8UBWY0W2Z?]^M=>Q8
SZbe4<J-0\fQGKF&N1,1\fdE4##a;U=0FV^5D9RU0KTI6Fef7ZF.0/#YW-U05#H(
,H<ONLSMUVfK2QE,;95c5WK/;Q:c.IN]f[fVfW;U:IFEc47#c6,#@L(<SIQNEQd2
&?2EBZ[?B?aDG)A8LKQMW&RX_\W3+KJA25R50d?b0AGC-0GF8EX]_g^8KNcRO<JL
:(d:O=e785Q7JO@VH8\J[9J[LCFd\E:(\dD6B8V:G_;a^>+MUg.Q8+.075PH;MeJ
V#Ya/)/O\Q((Wcf^IZgCaK\674EOGD(DJb:V.Pe3N-,f31N2c5Kg2AQaBI8M^X_K
@\/2E])<?R/?,e@?FM1Te#:0^YP?=d/W_dL>J4H_E-<aL^(+aH09VSH]_H#<-J:4
fZ.bT+9SKYa1K#09?DPN7(IaOZ3YLD68L:b^4+GIGcU\<YgS@YCX8U0YUf(^eVV1
/FC&KC:fF,.\72cB-Oc9=<8TT:PD<J16NJC#B/Z=^(4DSS:ABRW@7U#ENSJ5a]-3
J9fH00Z5-/R3d)VX/,IbC6gQ9;-^KR-R;Q8P6N(TEDNV<_U/U(b;NGYUgO7/&PDg
-;:Z@7/d9;QFSTL((bJG?#<1E_OdERDMSHO;4U@A>&V#=Gc>9(R<R##^ff.4AK2@
P4;,f2LaW73gVAc_@)bDN.]bZg@>d<HE8?g=H^2B<@H.F<9>SKEJ)G34-?K<U5-K
#f0fQ+g#BG<@PcRN0(3KAMeWI-O-ZDMGD2Z@?@@Ab>Q1IY[^28)=.,4,&:=ABF79
2@Na/?[\/\FOJ[NeZQZgfJBeSVc:#JcZUDe.a,H9M0RQX;]F)UM\T4Q=10V1(c;O
U_X#C;362YNeGUYDZ(@[c/1-eS3LHHWF5PAF6VZ9K>HTMPM#@RfQcfVK8_FQe.e0
ACE<:Nd<WSK][^gV(IMY4ZW2W7H-AC=T^GV&?@SB>(K]-RAM\Z&+)fc9/^)02d#>
39.-?;c-Jd;B.U-g63E:Pd?&.F6JIJ0OSc?J80B?a28fDYAS^W1)].G=]^FBKZQ:
9>\/,gL4<UI00)J2GKXUe7g]&HNcg)KL?^G^aCNIMRW/=#SLO._FGH<A-I.&KQJ;
[3JK9>R0HNc]f,@c@/c@2c,E^=EPOEa3:bZc_5^S)2OEF8U<4,ff@MH8?0R2W,C-
5MT&3KGN\_J1b-4ec/D/FXV=3B)f_M5M+IE\5IG(EQWQWg#5@)Z:(eNMCJZ?-##,
6<cL0?1SNR((a-NdF^X2d.X2WJFKc<T37(6,C1^-JY,/G90:e:HRI]=YPW3\(/S_
KQ,Q]Y0(M7?+a]K7:(?cS69F93VN69f[-;Z(&O<G7?GYb779IDN&5G0-e/J9f8#G
Y7.[[JcEHV^V.@TdZ[NJ7VR=9^T?+@ZUJ1VFD4=T<9CNP(J24ASRe/<G4W:cHL:@
3,\L6Bg<&/.3[T0b2=C^?FR)4,b45C2:bZGCD+e^bIRBY5#AO33eH^)?Q[);^NS?
GV@ZJ.;^R9[F9/Z?bRMU]6L+[-FBILY:X3LT34_KHM9JH_\Sec9V>/JN/MUIeG[\
8Rg.Z-3&UR\T;-5Qf,7N6b5X?GMI;.CL&4LV54)O@1MT>RS(+a?L.S9A4A)#I-^_
e4.U#[=7cc-e&(2#Jf29N.9..A<X>2,1[[(+X6;X/;aV2P;A2PE5(W_[V_HDC@#5
0Rf_,9.1-3R1AcLcHSB:,@,##MHgUN,0#EV]>5W-J58:,G[dOL8QY^WZDSW;cU(U
)4WTb?(>TB_HWE\]TKYY#LK=eDT839T&/PY.\[d<WXQA@c?gBJ-P/g#@I9)dZ[)e
4Xdd-&3;IM0PG-KE2\6/e3_#^\YQ@f30^O<eI<dRE6^V4G]9:7V4/NLb[L32E)OW
X&CWT,64H9\?Cdgf4,/C=Ia+]((2>S2ELYgZJ#0Z@KD@Y+M]?0c8S(JX/bNgcE=&
A];be(X=Qb+=@^g(535H71:C]NZ<[+Qa]cBcSEV1(cVg;WB&,4,6(e;eVUB?=27\
1AJFB^e/5)>J[KYe3RQb;>_RaB>;G?@9AO,L08UL.38?=eRQJ](\:PTJX@91@X1(
@;W)QJ0Dc&8VFLIZ_a0D64W-B&DJ9A=^V&^-71\74XAV^WV];OeZI\PC\ZfI3=Ff
+Mg,Q>)a8[;K75N9-LWQVa(]83;6@eA)Rf&fJKOYdbA7=FN^I6VPMLSGNQVZCH<4
KFSgU^d1?g959F(gg:/:N8bVYCcUDd,<^G0TMA0=dbGFDKC+SY9[^(J6N>YFI[Rb
[[W;VIU?5f?U19Q4K3#CM]_;\Ua@,CJDWa+gcY55&QTJX?6)fb/D9+72ND-e3IN3
c;WK19@2#XeHgXC76XP]O=E9HDcZN.[Z:e8g]HW+ES-C(.b)L0<ZFdf@KL^N@g/1
:@N\6a6J>EaX<J:#PU?f.Gda^-5^(d<)2CYWG1H+R#R-:NEbUFY&7^>Q=\EU@dX[
5(?U1OR<g;S7+_BE9;6FLB-ZdNFI:)15dSQK[?>^A5M5W_140S8(J=a##Q-Ua77G
706&YFPIe#+.[9)>]Ge>9H+^[TY-\JXS;I,c8@bPNHDBQQX4ILR4R06&f)(e>:/K
/+DfE?#Z4_6EBdaTP+db:46,W77GBd00.HLB)R)(g\_.Q:Q3a,2DBOL\[ICVBC/d
Y[7OPZf5(?O+^.9<:^bfY^.>\[OK];79(4d];0eb5]KbR7+bR.CV(?_#&8B(^HZe
X^W@;a\V4NN<d1@T0I[U>P.e_V]K_#]GO<MAW^_39V,>2U1Qg^R+(+Y1@fM2[VGD
6X11DF&-DcXUHQ/B_B9HG(e]aYNMC74:+Z)bK6@U9(BITLZHa]2M\C^WS(E?]6L:
=aMKP9gZ:2<GIH2aGHDL?IN=;)M=,4L56W.=NEWRNXLI-577g[2G9,4_E(@)7E&<
@+46XfX6,<Kg/]R>X@<.(+f<U7gVK^>(Q]T)=F(HUL<a\4U<3/)L&Q+c@Zf[(S+Y
4.QBb;DZ@IK[PgO4@]8U5J?_5cP2fKH5;NPaO.VEWKK\E.;=cS5Ba^g>,OBX2KgY
V;)C^a;74HFQ=Y/C:Z_SJ30>0e_+0Xd]dEb@aEIW/7J?QH:f&<VMPEG1.66#8.XL
TD@^:(I4Ia)FQ)F/1Qg_Cg.3QGV>bPU?6Ff3&&VBeb&=)/0L<L:NK5U[b[M32FEd
Q@\eC19H2)MXO(MM0QWXA@d40SX5?8^6\.6#^/e@GZ3b^:<WI\GB0@+e0&UgSCUW
4N;22_:bdU9UPWON2=+LgZ-S3;dC<F9DI=:#UNg@^9YX=:GW\g_]K9BW4K2CBMN\
YKD33]YP8aOD,S_,M;0gU9.d4OIK)5HLJ]A+#fb;Q+PMA&=\T81F1MTP9RLO<22(
RJV(7C+/]QLJP[[>d2b::?Y7>IP/T7JE#76>60FH,;^LbN(U:^Vc2^><(8dP@e>/
BX])8>P[ObF]HC/G7/fab0EVNHb]d1-K[>]RQY=HP/B#AO(5(bZ&QQ&=RZ);5BE>
<AC<OLc6<bP=3.NLWe/,7KX>,:W^a?2eQ,6bZHTf3;MU^e/;=N/NZ,\Acb(b0VcL
DfIMf+V^Bf;NG&g?+BeGb/^4G^8;]+HID\&S4^Q;-3<3Zf:2SaTX.YB<[S.#+FC_
@^aWUePdA3fA:WFgVNOTW;W<[]eG[Kd<Lg;5AOTBR-Sa@3SNPL+Z3V2(<8<JI0-A
PEOQ:)0-CU3[JH@WOQ+DI-bEQ[E,--<B@W4^Ga>@,]]A@/NSVDa7:>>,EZ-OC-F1
f.RI<4[=Q(DEG]PYR&,.gXK1SZfV0bI/[\.3,1GEdTcAR9]DJ\S+0D\BdI2DR+]d
-<I./+P@aCV2HW-+EK-7[Z8_>5_[CYg+VJ0U-abH]Z>F6;9?\Q?UDc[U2UR=Q6R^
MIDASbYPU>LgNW74S:GL4f#0JLS1,g]49WT7)C-:X])VH.);3O..6#M(U&dQ+;M.
-/J5@B:M5B&WJPgL]9WT=?E8:_II3aMd(90<-)I\1YZ3c3b.A^F?JH1e2gC(WE5#
[RC^R=:(W17&3_aFY3Z+(U&IZ==dag^M-b:&+]Dg).f_=G8WLWg/PaeS(@CLSB1S
Y_McMObA?[>K6H8.M6:JRKSU-U;U7(Cf5e&IWDRISL/Z?B1I-_3\26_cYA:D)H3V
ZNWGS.df9IaL\9fEScJESfZ:cI]E@<>[CeXf(:e8F9c>g(SbdcMH1UD=XD/J(M1S
V4G4PJT21BC<FF&.RL?;b@_18M+;@OD=cR47c6Y,d?b6SF_TUDJEb[egHI4T&?I_
bP^1G2VeaCX<&Z59[SU:gc<I5HY?F^_:2B6)#VC;V^1],HdZNIA]]8S\/06CW.fg
PZ\gQ<^<UYR+B:.R0b)ZHPRRD>[QNX@9\Y\Id,gJ2gX=<9?VFHR38BDa,&QJ41KH
L(-Y7,)ZYU@1Y/UL?g?ZM,8+[R/=989Ie+:8=P5[c^1#MgdT=2)(_@FTID_^_)#U
P0fg).E&0O.FBf3R+\5I.H2WZ+gHP2F-5RcZ^Ic470d7HS\;4g+E4f=9IU<K@^6V
_/D3[_0,:3QT=:e\YP;]+^(,7L+)&(<=a#M6>G\dW5F7-b8:bL;S8;:#cKP&a7\b
H\HAHJI_\_J9Y((T_9=(/6AU)Q7-b.E&-Y&b_7;_\d/XU2+SYXO1]Z[-<\N\/6Bb
/:&U<>Ld?U&4=;2]&?>.JK[]#T+I@FJ2(cN/+77W5\\Q3(^OT[^7_4R<dW2aM&&C
DPG;C/CY],5Mf&cSJY^P-V+Q;)A48_/?.O^XfdK@?C2NLI+30G&WZ?;G3>@?@+&7
3-^73+bU=7bRV,DgV+:7]:>2KQ;#TOT,71eg?P[IcV[.GEQ#Z+.8R:4UJV6BI=8T
Sc4X0^]TTc]IO<c097A.30U+V-]KX_T1UQYIUSG.-ZK^a4C+J^+b)W+3T6\;2D#D
WOa+BW@37,NOX7>;R(A6cCHROW-=)2@>AeAM^L\KA(3<g4SF(Z@E5MUa+ZdWaM8/
-+af-1+BW4K=ITC31]\/YG_dY7=(OEYZebT6SA+M/L5\#8FK)A?_KJDR(@[01NMe
-1dJF2XW@\L1HHIY;F6\7-]cTa9M>7Kd_=5E:DC23S->JcQP8-O,?]?IS^g\>FFH
;SR8_U[4E(Y_1Z?CBYb&HMOSEgX#2f;Ja<AWO(>K4MPA@;#N]B20-1F;/DV=PZ\T
ZO4-RTM6N)ULAVFg#1A)>9cB35LPL.X@c:5g2I6SGB(;6F;DY#E#N8>4M+dU3SX.
R#c.<VcA4Ub^WI@;d^,\?[YfF>(9^YbWT+MHX=(1:T-:ZeaJB-)[>N)8d@KRZ&W7
U8ROd)JIODWgf<J/#(QgKf[=g0AT5@U0^[VeB]0PT2W0MU)d8A5IAG&(8&#D9TOS
KG>\;Z2(b\gJ.^RTaZ,I.J5C)(>KD87>F-A>B+7G;9#JKbdK\_;3[8K4G((dHTO)
I?LfZ:cT;@7(Z1.70)YEdM+)^D0+KAQGdOg4WOZaTIY^K;^A^7^:V]MP:NHFTQSS
IQ9SOFQ:L>c/LRf_7EK>OAKZGARKKVCEH_Z__D;5&EYNFP#MN#<,P50Q9,KRVV(4
T-gOD=88?7+4,M[4(6)QG&TF1PM+K&QPR&YNUWgbTJX+,.Z(V@:M9JX2(C97C8AR
<.13I(R9?KEDP0S0NMQbH3.Y^Hb5^H=d<TBS+@1/YNfM-f\dAT_bE8.1GcGIG.A#
/?f:@A.DGON,^FDU)BJMHYMHCE3PMH\S[IB(22<fe/MP9\]B-8>5(.beL7]IT1&(
#=D^&6e,:eaINE=M]Q-VCCE0U.cg#TX9E5@-CK])CNXdCgbcK@@cUQ^W\<,]Q>UY
<<ULVUCVZ@;_N-95cLQ1I+-1F,+KAM=QAE=7YaT^UfQ:CMF6f\,0-U9NUKZa0Pbc
ca?0CKVOFfMM]TAXeZ)M5E9P098XGEHBU@2C^AL(]=AS.ZYV<(8af@g:KMe2=KE;
=(eI6/YLN(]1R8&C:b^BNV_I(4XH&#5_N_e>A/>/=_:(LV4KEe2/0PR6a:6?W4@=
gBQRCg-Id]G:AP^3f/S4JD;Y_S(7W_,6f^[_^L34&7@(?1febdO<&^L1<1Q)IId/
UC^C9EUTbS537g&756KYO24//>,O#KL9Z0G)-:2Rf4W8?[:b<R7\b6R\TMDE3K;-
MYdPE;LaZ1>4SP]@@,QA-Ge)d2eV_W&D)dLFQeX83]<1U801>1Kb)=09BM[:<2FW
V@]4M^AZTV&\C_1CD/?K^R@aYY)ZeC((Q&<dWH0?Re>eaRU)+#cL&[GRGK]eLSdE
455?>#:2E&MP/b;.(aS[D]R.4E.I(Ygd76^JH5_T.BU4effP#K^R87(4IE3&]V<U
?WR;+)-4<OS0@41@M:HU#AGV91J+</P5-e.FGR0C1HMCM4T:f2Y)H83S\FCTJdH>
TEZF]:eg,>fAg^T]fPRRL9ecCDG4[KEDaW+#GI;RLg-AB]d>P5f1X)&/TJgA_f7W
^BF]LGb-f8J8DM/GUU.&GZG+F+A69d,HAM-1SfP>+[OX8B/+2\a+QP,W1>82\MJ6
VRSQMXIL96:+LfT&2UW&^d(T4E,\J]#I)Kb#fbL7GPea[Bf[W&eGW2J-^5E<SaRS
4C1+@.BA7QdC?_A4LTO1dGgN_,a>-5-QGb0OYa2VKD-W^aXQ4gcR3?D))<)N:_Z/
DM;LEMH)GY0g>8?JO/2ZI_\bA=Gdbb,G4.CG8C/>dPfX,BDW=Y:5_-UNbN]?RV+5
]&1Y,-A=<;d(b5XbHD.MZRDa<81a<]dQD-Y@T0ZY]X@aMRU^7FT#:dT@_G#F#V>)
J;)M>G(;NF4N6eE59I9@-W-&GC852RBTX_00<-VYdf_g_U(7]Uc8^LVQ\#+Ld[_I
P6Y^1H[?;P9g#[(M>E/DDbSAE23_]5b.;dMUL<I_e-7(GYHdeM)^Y\f&6.2g7##C
\<XX7XI.Q(</)99e]1QNO.7]8BIR\P_64:>f1]c&I52JNTEX&ZU4/HN=@Z-D8BBA
62U)]^,[Sd7/-4^]>CJ/V=E5bT?;A/VV<Ifa=Jc>ERB2L_.&?c<CJP_:?9CYb&W#
W7+deXcMLf:-)XN&8/#T3N1+#cW-9cMLTfC+[Fe7-,JaQB&=8-c9E>T2c9;]87-,
+F<8a9G0,CD9MdfBQJ-F#;HFafB_(caP)egbc7JD?fT@VLU@#WB@8]G7ZJ&0BEZ,
QK:a:__.1)7J2G.(-b6RI;6)dKTZ&LWb^[R]75@+D8S<dMTNQ8#d]A^N].<41aZ_
(I8,gL\Dg?F8B^JNeO[_GDMcZ14+[f=^#edU^VK_.<aVWWd_D4g,5gQ6+&:<_,2d
^QL8d18\3;&:0f/XL_Z@#VM[Z.dNB+<;YT3>5M+:>Vd>NLC_=FWa-302ZR<L[dPe
I@8:?N+c;g)UTO,>ab(J1H7P4f?ZLVA]@+OgGZFNUXX8#/)NaJdaCPKPY1>AL5P7
SL+YREVS-D@1[1):9H>RXcE]EMHZbWR^;06Y>D0#G)9Y0H;([W[1S12>03]0eZ+W
)dFS7W&)D25Aaa6=fYHFO>Te^2.FY&OAC)GWcUX:/+_OT,@Na62T?007)VD[?1fD
5c;3/.:A@KO[KH-FLXQ\/QIU4<9.2WLcVPVeX79(4OU.XKK5;A8H0@;9&M5W4GI(
c0P&>5>13TE&eGAVX[Xd)YGQ]&&GU4/PB1AQ8BAY_.RN@^Y>6D<[)MCL4&CP]I2a
5gc7fEF#Pda_D1Q<(g=KOf,aGV<.Q.;PKd.VW3.bYc#-S1#E;SE^A[Q1aK#fX4HQ
<=WD/L;>>Ed0OLdKW4cBXXB9DJgE4&E,Q07WBLM;AXcf72>V1]9Q+@A9cEYGYV[=
cOA.:+MZP@dW=)/>9[TS:TBJ1)3.KGRF9G5PBIN#;bC\W]d^/[GUT=_He9169-[3
<YVV?SO>A93PeU5?e@F3f(83f5<XQ0XNP(fWT@?3d67:VYHD;,\TDRgAVX4Kdg52
CJ?9(_TOB)EaCb;>WG<9HXJ?)69J0fN&O?d.W\BC6<\TBfHJ[)_3:ZM^c/;GR4AO
Cd9S,[G<DH3XXH)9eZN<SL.WIMN6cEB^D<:I<2CF(K5OI/O0dGR_bOHB0-\#X[PF
(e>1;CT-KO48?IP;gd&0gXZ?&ULaU:MM;2bf2<c><2cX(RQ3]#PXg^X:^>#5W5&5
LMKOB.U\_FM[Y4/EcJSDZdRJ:A9R&W95OY80Z;)W3U?CL#:EFRceK=TV=70M_<4d
;(@<]VC:D;B058\\\V)(Z==R,&BB131Gb3&?8LZQGM7BeHYd=>91UcYC]XF..8eV
I370(VFOGC036^Z6&8EK(:2^C+G\>,X_1O7O?3^JG/[d6fM\<Z/9bDbLG3f0I<G-
Q,ZI^&0Qd9]EDf\5e/2O?U7OTPR7_58bTJ]T@OZESTE@_D>61LT5)M0X_OK;G^]S
JT32=+5N@62g0f=\3W(d;CB1(P.4P]f_C2<_]NX3?F3Y.\[^[9R,RI#AN&^<77-(
?fVF)UBEU=2NbT8F+.,1cFU>N;b5fdN1aVD-_E^22M#0&(WL0YOEBC[V++/X^bCS
X>Rc/W#K<J\).[Q9bdaYFaELTe4cfbB-eI.4.<Cd\08A)5FfY;&SP&8P1?(b1#MN
??,7#[5OI>AJ^a\K29K8CIC/B9\:dZ[,.5>H)O4^c?Raf=aL?[Q=-/e1+g;L^P5H
(GbQ)OL.CaMW5I.),SQ7Q<aR@H+&Dd7[Mb-\EHB[G_Vb)_(8-[>US&H=^Q,;d3.(
?PFW6^T]BD]LGT1-_<8Pb/=YPVNfbNeR39^/V4/0#7;(Nd9eEF]U/cSEP6=R_bYK
I@8aAD/_0R2I(]@;5e:4d-?8O\HX1)OB7d30>GN@2+aLX^U@=HI:bEd^1423BKb?
B6)S-#M=P6S<:U07;[E#UMg)5Q35dL9+KC<H)_gCdE:FFf5^-DVWYM@/RgW=SUAT
bGV7cLB2eT]^0Hd.S0XBI^KdSZ6021.dMHGNe+P=H=/K5IeWME>#OYZ3=;8_g]gV
G59(<Y;P/b0>++VYU>a3E.aU3NDWP409(Y[.ED:902M@Rc?T_6@&4&<G813fC2Wc
YaP^>L?LPID@U=gBd1Q@Q?GP]NS3N?2\2EXBT,XN+bS.Q@HG8gAgLYCR+g#HcS30
BB915OUHgW[C;V529c_-DD[Aaf,BW2/=d&7?[8@,RMMZ\JEZ,S.?-S3A.+[W@OS]
.W00a\?CZF[]aOf@+=6,VSa<\f<Te)X.[-dEBJ<Y\(OT(39.a<&_U/ELN\1>9:P(
5)[RQNZYZW]3T9a^U(b.ac/<UA?N@U_ZAQd4&GK6<1>\=?FWN^=U-1Bg9bGY\e6O
c1J_),f.DT@)5EJ;<bPXM3^,018cI>Y1(@H\;N>\GX@_<7OR2.,fLdY)IHNg3>F?
4N?33Xb+/P=CKdZA[gaMN2#bLF8fR&Ga:NdZ53Z]7+NNQA0,UDGe9+=UbG?[E^M;
AZ9f:G,#GOPD4[B;F[#+6.7N<.TZCe.M-aGff61gTcN)3Q+cPHMe-;W]YII#J,3K
Je9M5CN.cN;2c3Z>JB\4;.@La?B_W.d:4FQFa)IgG-:H>5.[7,=?aKO&1a2,8;#2
VG^TfObD1IdB@Qe.4S>T@J:fY]Z]C,Q;QDGC-4RP5[GgJZPS^cFeLDCG3?aIVc;/
O@6[5PP86dEGa&?MB#(f=2E==NIOD2\-2c4P]bN27?c[bf4KTA#F5?=#DF&#]8ZE
61RQGf86C:72QS^ON+B&F,S)70QAU2QXeZAc@WX9XKZYR+Ba&6EMe^HcIY(>-(;1
#4AQTFRZQcbE1fbR55EC1O3EE1LZNSB:[16QHIZ9g2^8=,Ab?9?6)aEQ2/53.26Z
<]bP1;=ZAH:a(RRa^O21;4\X>O1Y#.-0H2JXJ\2_U_+D^eK@dT9J\g91.7b2Z<XJ
A4]7KPHF;1Y76YE=7D7RS0/GP^H=<,[5D^X1F:N84S\ZI)/TP0FW@&@XXd)=I7;1
JaK;N3MG@b<c>LO@H\UAQ3:4MdJ>=1T<)JS@S53OW2<8F1D;5d1]He@;J25QAFaX
+C17(bS0JM9DcJY+>3&F3LX8PD?[H8&O+>/@H)67F9E^^?c=/>G,<&H,E=/I[RWQ
=0JE&Y14;C2S,I@X^C2bIO@3]QG]G#_S3.(6:SLY&>V^Q&Cf8PWZPa>gWV1cXQOe
0;FRI-Fg[7GQ=,d/bE5KM4/LXYYBJ8QF34]R.2\?R?@\]C\3>Y5D?/5T/;=B+L80
G.2=/50^e<EHN:&1A2W1]VJ4-Q7JRW77J#TWg?>S)[(e+5T7,,U\51V?:O1GE><f
:>dVM_SC@<N/SG=fP>IC_KQX>a=-aAP.BQUD@Y^Wb;P<LW7P^LB):KP1X/3,,T,6
VIFf=b[Y6#R/9fI[MQ^88f,>_f1\0&T7eGS(0&TAD^ACcb6Kg<cO789a;,2DL_;.
)^)<<4SFb/F(UT]Wc:,)C#B#c3:bg^U)80.Jf<5Jg@K]#R/Ig=JaK;,[[VEc@0O5
879_e[0V308;Ja\758U;Y=JFHK:P_K)>aQa7CY>d;92b?]dQ3HP59TPU[df--2@(
D\Z^LI-(DgEI9H#0,2dEQ@)KK-I&58@BCdJU_\d+GIOQ_[fM:8>)R0Gb^SeQeK15
(-]C3A7MI?=0Q>c)>Z64ObK]<6HE2FGRJc6@fXg9)/^TT0gH:<[S>V.8?V\+6WWc
^>KA26T=(LMTU^XNRK&UB.E0^CT;;CHTT3SD\d-baNd:.^(-[#QC+YWF:P2RKW:5
?a&WTVP9XYR:1AW3[Z:/4A^23\HOUN@[&LKeGf:)C]=JQ\6#L=7BCe(:;I)JMR;e
Y_?\.91LdbM[<f9@f-1A0N.^_Xg2-d\(-Vd#0WFLJ0aC^P)Bb5>KEQUP,1W@^2f;
_2<>FU1I,2M(978SV.62I0XG+G5T1EY_PTP6Md7g&[7#K/>0:WLHF&JG&8D)JT,d
,,eb@GMXAV@+?4[]K\X6F)a[:CL_Xa=W\d[PWCG01/V=MDL9JaL7>FbT7A+g;d8Y
,DX05g2^J[6GY--+RW>EWGg)SQ1D\7BV.PecX).,-XLQ(cY&aG8;g,[7KP<E6b),
RI#Yge+.+G=<YC]N:PU)Fe<eQRY.V0/HJXY,JXEDfZX=T^8N@YLA&)22KEG;HL8S
Y5:8C+^PX44R+^4C)FJ5CA>G/#Md1JB;^<K4b1(V2IY00A#SV/V9;:MQ+>W?dCQg
C\Z&7B+4/2-.N8BYe(,CMV3UJ=@S119[M2\NN#;].3QcL#6&c+=P)>ZV&BC;3]fY
,@,gGB,,VI:1?FJQP-<GJ&[a@#agYSR8NeR&.TgRBLcB9]KINCBU<8LHRNS/MA;M
[]f.4/dg826(H9.@]7+1FM?_<9&VQC@0D&^)L]dI=8M0KRAE8Zc8O&.BU.LB@AL+
V4>GL]&8+:/TG1[E.X>>NBFR@[OHP+g-JB4-7A1?N(YM[Y92d:\g_ECe>D5e?UN0
7MKS+XC2&c;(J]P=>(PcU1@cOS<A>5GKQF0;6&-&YLKcQ.Y&Eg5F^HO13AQPTY=e
O)1+DXI)]VPXD:M;J1N93L)F@ceb0Z&bQ4Ld&DQ8A(&T^8SFfUbL(<#16K2[D6Te
@^4gI,>C5XLX1e;Dc21\6IRU0/26d6N.&+3<Q]dDLEJJ3a#\K&QAS-[7dU/9)201
bE6Mb^.?3>EAFSC(R5]LV)>)L2TT3_>gK2[XXY&5RE=d,0YT\R5eN8I[+V[OV62A
[Q+gB/10NgFfM=Y1b-@R[f97_b8_,0^NRcOJ0Bf_N(A@d=aK8[]JQ+<.bCSFC9P&
cE@4^9_[SC8+6:ZN_VRM@W]K9G>V.I-C(Ia:LC;@fYG51aaP)^9G3cBD[LK];=e@
FE5R@KO_c8;T:Z/7TW_c=94#Z;3#VY[M\_#098>F+W20K^^^>EF_YON_HSU#A0)@
V/cTC4NP)RgM]G/cDX/WK&=;L,:5\Ye6FI>^12.@0_KU4Y,&+;bFZYK7]dPQ,&6Z
/(42N0#F&R=.;45PU-0M6F[4AA=[5FdXINLa/7DY7XC:6AF>@VV=g^FS@APWcW)\
D7OR1Obf?)F8DN66JDGT.;8G<H@U..0FY76+egQ=-PLC-.I[HJ++-U/_(7-eGTX>
f.cgI-K:+,MFKGT\3[:/_MbGK:^(4W<UJ:7XB\=fPRf?_+OJ]+UQ#-N&_[Ebg\@2
2fB:[#C=R?IH@^N,>>3OE0FU/NgG<Q0>+9/fcXd93gNREEg\J&^FZ2Z,](]\=<gB
4Nc7MXAeD83DZ\PRO)fG5]e>=b-&V2a2D^?+MGeA;Ua),GUOe0D<R,7JXI]:-_+?
bHf9W.M1f4G,5f^D-e9ec5Mf9ZF,S[-dd6;U(7>+^(20/E^CZ+<dL-5(?EPI2W:;
#(N]?8(MDK+78B9+CG3-^PWMP/>FdIT-GW-dEdQI.,X-&\,G^63TJ&L0_O&7JbAG
HK,E8gG.CPL,KQNcSfNNV7ZIX;=WacbcZK+Kg@+R[7afNK@e-YXf+^;DOI63ECDM
eT_O/Z6NVOT;DDZ^].^-\=g;,eS8@<,.S#(e9^]3\6Q\210-U^VI+.:E(PaOX+[[
KHeZ\48F(UHCYNGGI<:bc4d?0L/JC#+GI&HTC,e2;O0F#Q:aZD;:AEZ6RWOaf;7G
&cVQ(NQ?VUXBT7J\.:F.aLTH^O::>43+.9S/X7#_U52aID\1:XFLE#JY#N3f0g4?
IcHHG2.]S:6@YMb,4C@-X=\>g/ZabgPW1^DP_5H3Jb\(II4UH+?b@c&@/GeY9(6I
Fa=.=QcI&LMO^(@f+QS[_?fggaK&cTLdTWW;g)gM8^3<FLgAfQa8]NR:0Kd<G+G^
d<O>6@f<ENO+29aEXPV)T>&9LSd^d7T<:(DCZP-a0cEVNPQOUB32D(Sb,:EK0(7>
+&_<[Xd:(5a3]d1=1>6L@S<M\6_ZB<2].cSD3Qe97g<.<-7/&OJWQT2O#J.&Q4QH
.HR#&OXa[=^7MVbMdaKBObR?ZQN5EY5(&RT8)][LfZL/^,gZAfD\?I8e9/HPX,0G
+0Q<Y+EZ2_9#6SM3Z.@2(KL2)P:;?9C3H>5M5/PUK=S/PGdJ\VS>-KSabaJN&N\I
GR?_7.@I8I]g6Jgb->?4N0L.\0PLeZ?FT0]DAF,=[f++KD;PSDfB@HGWE+CYg\Pe
QUaIId6^-?R<KV9X&<\[_,V&]/EO7SE\=?fL;Q@Jf,U,2S+=5[B<5O/W9;[0/@Da
9ACTQ,-2&MY5.3X2Dg)-_,_]1PdY#9[AR9F&>_]WK0)+:A(&L.7JS0(T1CKEO,S6
)UW=6-YUJ,,);U=>MO0E@,SRN:I63/=G7;>1I6>[,WM71(ea@.O?4<7+U<^IT<>B
6f&g4;JSXM2g]+eWGI5c#9JUe=0]a;8W3+IRC3MD[^N(a/4.FHB)/RY^4a3MB_=1
/f?ITP<VDX4V_0HXEM]-4:.Q7HGTaaHd+\/c1.8[N6?d8<U1\XUfHGJ;DbgC:5D9
,>OVd?c47fK]E>F6:=ZXFO9Z=M-8#9J:T&_;PHK/g8#_U8Kge?SLEE1Nf4.(Y.20
>3MT&(6SLM2U8?cSK)7V>;,U;LAEQ#Md?ZCR9.R(&E1>\8+BPWYc^Y8a6NLZE7>F
.@-QRCBDffUJ^e._b<^5V2WS>HF9.WU9&8H,6E68_/^.5QGU^>fNHIbC1=[BLZNO
665?#bP^T?YZVWSUA82OA(@/LNPgMT=Q>JgXcLf[\;C#+W/gH@EPegPC6)B.g<TW
_=gH4-7&7DYE-,&QQO/FdKJ6W(ACaZVEgEfEcaA?]G>[6_e_34bWM/Y@\;bg--D\
_-;F-/fVBKa]QJ+>&f;]cVK3K,a6XB8IX#Z33H;4SR6O7F,.6=fC3Y4K9HW5L?^Y
fAIg;a0Z^VGb@HY>AZ?5I+G]G6@>3ESVMD4#P1R&N+G4>>>IT4PJ&VNSH-ggX;_S
[6RW4&&d+<0-Y+/MN7gT_-9ZSTMIdQ)5(g_AABWJe@:_J)]]AYKT7H:ebe:4bO2Y
TDB^W2=^81fJN;eE\0BGIgT^0-ZEL@[[RKNE&^8b6?1Yb#(QSVD91/BL3?S/N&09
NU+HD.P4H5COIXPQB;D9bR3,Le+9YcbO0M[Hg9,IQJSP:NcTA3FBLIHK>W=)G\fY
dga(Cc4RadRf+2)=]B5AIdWIZGb7R1]f3LW8WV5:b)YE1LTcGRL>N1^.RG/<JNB:
5W4OQf><P28Y(Ra.GJUd:M>OR<6ETV&/A,K_VL;3L&_Q-H?;KbFT9T7a]/ZL+-XF
6.3-DEg:@T6LE((^KUI_&T?^:P/\[DCe>bM@Ie/\QW45O4Ae^@K[[HY3(DYA71Ee
-6V_Q&3O&W8V;a6#Ic&]IZ9RP^5F89.,)38IMJK@TDZ.V01>U3:J?[#E[RP9CF_W
L98fd97<e\OS72Y#@I&3E8\g>]Q0D8\E3Y)cE+)-LCA&B<=)B&Y-J.Cd1J8](S5N
/>?2Mf)^@K_W#U@GY#Rb8MX.NS;cf3eG^KCaD@NK<E@R]()a3OI9Ocb\_b(TcT<3
cfU2FQ.8eWB<H+0U8:TY>=5e++GT,,1Kga.NRF^S7C[LXB[1Z[[gRV^Q(>6K^]&<
D[HHE=KI/cS<5JY2PX5[K.TgC]&;WeU=TBXS2HULdf-9)c00Yg4cc#)\H(+,VJ\I
FWSe7@-J516b>V-9Ob.BD+139XJUaEBR3e54F_>MA)Ta#7&9#-;7fQ1&R;[.fY7(
7GK>=UXbTLa@gO&>:>D)X6-1H#93I0E#>,V<T,AdLT-D+UL?^eFYU;JgB@\B3N4Z
O^]R<^dY\&#g;=N;7cO&V6a3B8.LRXT+[MFPSRJ\(9JE=9JXNJJ)R9(9cUX1TLEV
U@c[VTS===SOC]@8CeZ#COHb.M[E/+Y\[)3)-I8cSabZNALC\6B)?,U(3(0)O?F-
6f.#gDGB8X^Ag@cFUM_RBDKF?B>JJO/=:F[.f)\^^gD/^0a_2M6Z8:I(B[LI@<#;
T3;MdQ.@4/@3QGbbJI05F1D><gZf9e7J[/bRQ/G57?Yf](F52C49Q;:9N65dT,_f
[]?gSW;3#R?dT:2DNNddSfWE6c&,)+D6FY/S8_:L=GRN/]W?OE[4LE_^e^2FcI;[
+6F.gJ=aC:87P]fVg@)d#O_T\Qb>@fa==X<O2TY->W>(d.^S(Y0&\+PQV&R@S4_@
FN2QRdQ&)J^:g:)T^f9T&X9ebVeL3^Y63F?654M/T?4O>f&Ue9bB?E=4WIb@0eFe
CHV(>?81P1DD7J-I^;#bC_3f^&>RHQXK:D@[b2V@..0S/S<bfa[gTKK#0J@(H^>+
1,Y817fVC-_2\4,4DH_2D+N=-])gd6[_]I746O+(Y;+8=.JKP1c=6BL,(5QJAf)B
/J0UfG_KL:/[XC;O2/&L/<X3&9IZRV@Za74Q]GC0#?aL:GbQO:15Q_H/@S0F)f#F
UNDJ[///L0XCFd,N]daR)<PeWKWF88E7:F.,EP>CHJ^81SL\+II?,,&/T&GQLIB7
a,[K,3c@4I6+1DLI)Hc;&.QU6@^.,K,<18>[B6;Td4M5H>[7&c<gT8d\SQ^)20V#
REE],24TFZSeL-FYWMcIP<bQQ1)^.US30<&=U-)UB2a8QUH:J(2C(<(b+GJ.,C0f
f-D)):A1E2._/[?gPd_XN+af)JKN^USIGf^8^;JI=S[MCI2]R2KgOa<)9CC0@7_?
Q7#)KLEW?2>G\S^Ob)7PNU[&>P]#/4fbecCPKdI\)?1DEU)LM5=fY+dfbT5Q>JSP
[<[S^bg.;gO6XI5cE&=eWX^]IC99:5>g)<a7].aZ:F#0/Ie)8Y_NKPbJT^/Y+?HD
EALOT(fb3/EGXEJP\FHg>2V6He_@(c;&D4^E8Tf)423J_]1]WPTDa\8e_PNfGL/E
f]fA;GA_:I#H:XZ9>@aTPHWEb73T[+9eFZDPA+gSXf9T0&3ZI(36[:YF33E6AK-Z
I2_#(HfQ0N)CcC38(MEU>@=YAL?bg2QOARP/=CY5[XQeT+MSVM7H@J6,U+BG_cC]
G;L.Me5\4;D&K<WM.H1Z\;EB]DOTM\<_.0dK-K9AI>cXF)(30/YN]g_ZYfAa+ND1
C9]W-(H6AZI_:=8CDTf;8ASFgZOb.L1cP.W2.Q5MH03C8EL_;P>:/J4\>C)OKD6.
;2=)<:fL+UNHTESWKc2-G_bS>g/GCG.__,eRb.Fg<AX>G&K:GI_41Bg=Ee^1U+bC
E##cF(5>B<IEP]WccC>+SW]=/XZ[[,I<S^QO7RDXI;fJf\GSOLf&R<f9-SV6A3=T
Yaf73f+V8=R=C)7CV?0[\3K](Md[I(WR2#(<RY,4(b<d;)59fa.2e:?U=/P@E1S_
+^UEIU?e<YfO_54&7::PV0@]:OHTcTOe@P(b1GJ.W1N@1^HfdFLc&P]ggC+K(SRQ
0a+P[LQUU(A0dDYb9XHeSCG[&cKHHcA;^=WfJ[G0A7RGMPe1U?OYA#9?0;aDND05
AIG&0Sa3TH?BE5_MYeO7F05#NcgLX^MBK:Lb^fAGLW9+JP^.T-dNd43c)M9a4F@R
bJQ[(__bUeN-Ha2\MTC3A.H[NNWQH#McM]GJ+Y:;Cc-OOF6aO->WI6BDQLZ0E8#9
-TA;gLa63&^TBa_KRESC,)K,YPC04_HS:<F>H7:c@UNc\g;><52=+P3H[YPGM;Z>
AQA>dIe4EOF=fB;V8E=3-8JI0^+9(BPLNQU9:J(3=d>d^_NQ=2_Hac\Q>c+0S9P8
K&-6a@I0BJN7TEFL<DS6cMA-TP1QWKR_V8baYVdK/)TK=NE1V6E0XROD./8>;XU(
_YK6fYR[4]Y7bG_HI1DWM&M3]KUIe2?642&#7A<g\_(AA?L8L&c5A3]_gAKC\EH]
4+K-H?,Q7;]/A7;6]^O3C(6.S@_)3VT?K8/#7Z1#aZg:LM:dJ7\L\SeR0HN=,=T#
+]@12f5F41?&9g7d.&Qg&J&M)?:.#>GCD#?NICE;49dPDc>B&+^d+Z#_dXYG>g&Y
@aGJR?MQ#B>e>-TH\(Ae_IG1,[fOeI?eL/M2^4:KVQgOF5CaEN[J+/DcV_Z5PZ/N
7]Z]+U?7Jf>Qd4E)/(cXgD:T^W-WJQRQO3H42gI\b-FJDL7b+#N;T#\95@XIU#-9
8[E;-&F0M^ZFa__;[E<G-Y2c,HV;:G,L5G1-E/MXI(M72#]D-0C)5cWHQSO07)R0
&Uc.@K8D8UOGb/+fC,D/ZGUcG.:/I2VfXE^56ef/L;>EfCX-D+8Xc-d\X0KNd?5b
AFe-,362]dOH>_)C&E7U_aZJPR2]F>6.^_HR)^I@0X,RaJ/YK_)IEV/-.H7\GH8\
a6-L2ZMVYJSR-[6LNNV8EWPH:2T9PCL7EeYX3N[cR9DXN3e#\^)MVVMJc[V5QG/E
&-TNY2+feAaZ]NZ@Ld[[+K/RLU<d(0JJ&Qe7(^]WM-BWgJ>]c[@ZZF8^[,:0/2CG
.4RJ>8(c:B?O;)7M:ZIK(2A-/DQ^#N_#KKIeC,2F+B>&Pc(e+A.3Y8A5TBE2Z9^O
UXUC7+aMOFVE68A-DO#a&B5LAO7Ec_+<Q9B0\V3bd<3L<CKdQJ(9gB#>37>8).JU
.feC,RY:I4dF9d&FJGa,&YaF(]BR-JVUU\\]NX]&&9WC/6;PJV/WSWa]#O1MG1C6
I)cKdca1U^(L=>VEN,SQcG7+68#W,bTg=HF&eH#DH3:(Q[eWMB-c?RK97<a&T+A9
E(7WNaRD)UY1/62;9VCF/,M4b#8e5710/;RRL?2N/=gBe.C-S<E=8g-G+\8gd4L8
NWWK<Ua9)5b2D).>3G?Q&Z\,0?)Z[18H0fK?a\;feHM_XQVe[D8SW6S1X@c(F>B9
CYa>QEe\,.3_KB<MSV,\.E9dO[Q<:cF^7O:,Q#Ve&ZC<H@VA#Q=A3f.T^L)N>WQ.
UUS<Y8K5&FO#3&OK\?0JIbA^QH\f?PZbgXNV6Z\-G(4)DLB(7Z#R[,:^bd2g8Lb@
3FUB4_NV<@g#9UEWcFc8(HYZ6KG@)Fc4.5[#R_?>e=PAa<dP)MYZ4\D,[B;gZI10
M;+WC9;TW]2><YLg#.,IV1[KWSR=WfZ_d?S6ABd;AXIJPK>4;,?aA93b;2a5,VH2
WNG,K]1+W?E?&CZf.>0(ePF4DK&4RbBdaZ]R4K7Q+_[-H48U>7DaK,R]YK82W+KM
U)-BX2]>c^9^(g\DIA,IDGW_[,EF=)1C@P-=V//4NcB^GOD,SJ,[LAfP\KX82Ggf
N]RN]52UZFWHHIOUB\NYM=:OT)M?fa?S9a,&\:\UP(V7JM)V.I(ED>[Bg>GB0<A9
4=L,.Ke(QI.:-6/F:.K4B3.:T8;KcCD^6d@Y15=YKef\[E]?d;<cbG31VQZR;EPa
>H+KN;Y(<geA@HaF5@3Z,cc<)N=P/H7P@EC^CdCKDgZ.&6(4+c32.JAE;,@Wf/7M
?e&+#<#MZFPA:V;P3cIP[TF+Ye@:)7aeJbe=3RQ4LP/Db(/CIQFW[&d6Id>XZQY2
ACba<S1UWUN_G4LeIcEO-0ed/B&]Ff1AMVE[\Of.WX_KV;C;\aCCDC-U],MBU[SU
c;953,]1Y#-.#5</-;2eADgK(007NG&=LZ@.2gYZ,Q-_@bU4:.+<WH]+Q=5J\71+
@^AR\/?b4^/NPS<@O.4T]c5WM;?-BLHg3F1aOb+RFE97TQ&/5?@6G_5]5=9#TI4Z
P,4UbW)N\aQHcJSX)Y.D5?99ZC+IZb9B?fQILL)c7U)V-;O^_BL5Q<egg@IKB.;R
Ae>cW3@ga(+.Nab#]N1@\(#fbY&^6+JKNV9MdTP.LW=792_(585<Y;+C,)c7\Y>W
VeC;)(g[V5OAAd&-P<I[/RU=e^PEb4,M:_<U\S.:PEOEb;HgBFO-G])@PZ;1X=/#
>ag7B/7,\<e4LY=HU9edD)<JCF9^3K)WC^DF\@L3=)CU=A<Oe#;a)E6(f9&<)Tb^
SWXST&_/HV-:,.Y1RTY>GTVIG+]VYH6T^JHJL(MF=1I4YJa8FM\^Wd>ff&N90Y)C
B)62;ABQfVg-?2)#3>Ic=ATZ;3]R0B?OQ^+Ng+<dD:=&Jc6eW(LU2[LK6LJ6M@aX
a0KYY]BVE92d;^N_G5_1D^;UA7aH3ZbJ(PN,8]_-WR=E;\,8.X)Z_?dJeP3\G3;N
+\Z,4C+R8F<X8d0=/4?e/I;[HOLJ/.;OW<f5\fePV)B]fc.W6bVJ58V3U)XNYZ=c
BP82dePR<DUD03K^30O&B2J3(K4d+@U@H_2T3,9:dc[53\56?OD6?fEUW@[N@B>&
8-C;8aDRT/cc7_8J<.N2K+eP>LR9(#I<3[cWALC68,ZJA##,Z^:Q]AEe1RPLC6_X
4#X/g7(M_1(DUd]U&J5E<X6cf\f?(]=QWN5c7C=_K;O0=5Xa-IY2_7IFJ]+e;>,M
LBSXYZE8-LS@<+H_aHM20D5DT>2)T4JIeGG0-N-._MKB>(KE]&Kg8>O>dR&KC7BF
4[:e(Re1bO_+)DTE86CfOOKI@cg45=Q8fX=L]-(Q=Y>OWV[X_+6_HVG<^>@+R&MG
?d^H8Nd-DRO3M,\#X<5>[-Za?UMIXI)3WB<:D_2JaD-X2.RVZTT<,fb?,2gaG6&f
IIgKg,L3AgONb22[)daZ#>_V0c4WPGIcI3:SgKSfZM\f.H.DZ8K01c[U9AU,8W_Q
#cV[^<R,+N6\f>E)C0c8UMb-a=FU9A89gfQPP+7.DKe,K0&U^4(PW6+)51S@O0?e
\V0QPCUdg4&G9<JO1#9HOf2I7ZK>M_)F7IeCdU35Acf\YAA=MNK)dBNLaTGUF_7>
d>:S,149@e=.7IX6gVBbO?Y97:L5/RIA:8GMWe]O-Re&X\QPd;SL=ENK\M)1S@RE
c4>S7PG,AECRDHBP9F-W_/HI>[E@PU7U3#E,Lfg?10<-XaUYP_cI?++dN7b;gQC4
>^A?3g;CD;c_Q0W8c9^,A7gJ+e4Z3aC&IS5c>RMG0a(c4K9ZId6W(\_8KS7H(B>c
W0D^dYNW46E@c^_QYQMOg[Z_30W04g-4MM,_JZIX);B\Za8LES]6LE,g,,/11Xcg
O0EK3FOA)Ude?\<^d]?BCJU-VgZ:XbJ1UBf\G\\:CQ,Ia<f/U9fCBeFGJV01_D5;
G?8GBI]6TdCP\&/Z/OHP#J>97V(>B]A+aG[;CIW+E.D&L]+=&F&J68d)1Yc5S0;f
ROX;JE.T3[O=5YZ7.fP9PR825Q[cgeMQBC4(2.R#gNe^c0[P_begLCY\^0a=&P>B
Q.3ea(Q?@XR]K52@]V-HNX24G7Y_1FZa;eJA8&_;?\91+Ec\C)H,54\)JVf/e[#]
<M9\>D_#<])G;,\YcCVGMPZW\:<&dOP:XC&aCH1I#I38KJ0SXdF:R0U#gD0I_,RB
VOG>P):Q;cOGaDE#29?8M/b\<A>P-[LcZW8?]BXd<J527Pa[LC;C#:A@5&/UY2JO
L,WN7+fR&F4c,U@XK=Z=/a@YF]798\?5=FX4g9LVebD5#5#a]M-F(B)]/5-R#PO#
Qe8E=J?ECH&Y,(0@]gD-5-+^#:M72BbRW[TV9.K=]I79/@(S.N,\O@W#d.K)83D)
.9ZGTU(]UQ2^Q)Hf>H,D;AIWER#_HN]E2Q;eZV^SF=>?CZcU^f@0\2KQ\bG^AdJQ
7L5L:T5)UNDa^_94E.P.OA):5IM52VLUDa<c(?OJ7G[#O)ZaJ7+^P#N_/\E02C-L
:)3Sa&\D+##C\c,AZ0>WY/(J)f>^PEf#Ee..ELE9d?A2#XU0)EVK#T2fP.)CgXAf
Y/UUD=BVCYa7OS]FT]ZXV+XbeUA6>B-b6K=J#IRW_.A_;OTf&c3;TaNbC:?aP_,;
VSJH@@=E?DULR,8F)fE<T8a#AQ2629DVCb;NaOW6a7,_P\T28=A>JBW30g7H1,(-
_7U+5#GgbZNQa:3-FDLQN4dHd;g0ETYE9&^1N..X&Wac^F.Pd9WKc@U^S\<K0@Rg
BDANgOL6)9)9e.SFc/eR2BJX?4:e+SS<;X[d\,[X)#B1?BD2O.]Bc&^DIU8K_,bK
T>4IRZK2N]@fGMgdLPQ^7d61WP[eR3Y7=HZ\3N9[Kd^FI#7PJ\a>34gAc#R58JNU
.aH=fC0Fc<2.2<BX@SUY,eW&PWXX3BVe9eG0Z5S2MDg^<;?W3N:N^H&9c_P2>0DP
K<&D\bD5^3<&2,.;4_7Q1KW@bRdP,>]1>@IBWf-?[QLe9<KI)9H[5]B(E/DebX2C
9]>08..WgO/^SH0[3B8+cdC:;+c5SdI[:?T3E0ZS05@PMI&/@P2H-22X.(>;9,XT
COgF#I<a0YP66HfV4D62=B-QXK4E,MC8PCX3,V>#+9]Ie0^E3>]?YC/5X=I&H3.&
gASY(^:VSIf,b#.-RUV,f5D/Re67B_?604&^.7^bEV0XY5-g[DVbQIA]g4H)Pdad
9@06+&@0ZS<dF/QgP,5)2;b.OWF^PR7JR)#<cegDXWXdg\:(B]@:X0?X-W9C#E1f
c9W#&)^Q;/;d2QO&fF(7-#<J[_793&NA4E6J66db\Q4/b(0(HA3#f/F]R-c8,KPH
#6C#c>8?T[7I@;2V(Y;.]CP@VH7L&_=T9WMZ9RKc9K^[1\\.)QXLR-aJfW=:XD;J
?P035;F?L:HYd\dGd]9=]ZF31=.LN8WQ/.X))Z0[W3WDVb7=ERKHaeBa^LXddG\W
8<11A0CWEZEK@5U(M6Y5+Ga:.3#VEXf/-4YX5>\5ggRE^PW\-V[V;Q9EV@eO60<R
PM&b=.)?3-N)MRAQ5E#__b;bebA>3FT7BNFZ)8F-8g10IV[^aDg[#HA:<=QFGMfT
3[CSKNV^5K=OWIQ;PV?5IcOB/,>QRL5IA/RS#dP23K,N=]ab#6KB2=S4S06g:<YO
+1OKG6^0bK]3SJ.dRC,d7_Jb9BRMVMW68>Q+FG+E72QE_(R616(+;R:F<6IMFbK,
&JYF3;d#.V1_Ld@0ZHB;cH>Ud9,XX,WAU7Ya.B^7DJ)HR)XULf2OD5,(]Ae3U][;
<DC6;9>72)-OUH33([cR+[C<K+81@?6(7BTM624W+:Q8;I=(X>aAA>D^],^X&PGB
:.&GO;f[#ZCdb[5Vad0<-^S7X9d&6#fD3dXSDUAE#\M)#Y>]0/CDFDYfL-?\fg@.
DeL9FGFB7;HBfcRC&A3:[/CFEU^I+)DZMTBDAJMRa(I^PIe2c467S@DF0ZF8LQW-
efB0?9QCO1f&FAH3_0aI0.N6Xd_bDOU/DFTb>MV(H7S^(OJNLaA7Y2Ec0N&?XKdb
FW.1#[KQcZ&59M/-C-HCaH.1CGAc,??H]cWH8g3ddY_.4[:8XBg<E-A6_/&/7OXR
c)N7/OH5/ITGCa,U<E4[OGF5dD/8E,G96SH:+[+G.Ad+.TEPBaHYGG(W6[#2>3+g
K?#Y]8O8gB0V/ETA0JJP,G-D\F#AfDB5W=,RZgce+1_3I-THP]Z\4/f3b02gQYI3
[9G8T30G;+_@7]I>+).1J<JeBLDM<=]J?(7afe8VVN27E)2,=QGEZMUF<0?a6__Q
?&JLOMYX[+>>4b#;W6.^K,#E;;fBFQZ8g-TZ8_,2ceIL]0ZS^/<[41D#W3R#.8A2
5OR1_NKGPQJ2V-/Ba@Y][b_]T2IZ<\WE+0[XL;QZTI7b1P64J?E=3JH7&)//8G@7
W@E(IN\N06d\5I/fLVJA+O\I:&90)>\<0(UaJe2C,/TYLX3X?V,-L:1K+M^4?,#_
+FUe=<JY>AE;&W3M_RW]1Kd9KIEdR1DfR<Tf-/+2\d@._V#Xb5]MA6D>fTF)&RA0
[]O46FVe]g0E3G;Fc)LKaP1D23\f^a8fVKQ;dH>\U:>7K>)#Z_.&e#ASGOAa>FSQ
3bU@\IR5\9\A/V@b5-YS8eJZ)G.dR@X[Y&I^<5R7(7YJe@aCF:+T&MB0/Y?>EIPT
0TEZF+OI?M#7\:L5.RU9?Lg7PVGL-0+L1(\dXM_(8((EZc@+\.JGR3:VaB.1aCMB
97RA2RJW3793ZEAM<VDVK.bT/#gEJg,=_+S7_L1QY<cXP\IHW.<O/c)X-ZS^/JLS
>_CX:63C5(W-7QQQXL3GIKKBI410)W_.K>VGRJGJ9IYDBAZWOWU]5g5G0)b^IO(B
^AL;L#[8MA;:GCc]eRJV<Q:1<2CE+=0GEXE8G6e3_G<=gG+19=M\=@5.)W(R:WW2
Bd.N0]9&e\8,^#e356C^6f\]\+&\#Q_5R^B^]9CJMg]96:?6Fc-R;3dQKZYN4EL4
Q62P^J(IMWPd&CVAOB,,8NNI/4SV\_T8T&&-G9\;V3:c+.KB4<b^Ge42F7&\bQFf
)2LFdBc6(eF(DH)Ia^K<>Z6AbXPQ&..KB[;@2VbL/a?<GMBAHX]4-3]N5AH>3(C6
L(#f#]?>D(JbV>L7N86d9JAgAUI<eH._d?MOC)LS^]2C1KYLYMG-S/?<SfaW5BI@
8F(FYe7GR4c&K2OHYXgU08?5R7HeX5fW6HQa->R\,VM?8WGgYc@.eS)Ie2<g=+BM
4;3ETN&d^4eYeSKV#-I770(2,@Q/7WKE4D(d.H_..&0O^.Ad1dHFY=<.I@F46CR[
6dN21+M_bBUgg9G.T_?)2GL&ACTKU+XP)^aX1OITFV&SHZ@OZgW]gK8\:9Ha3C_(
e:@X6fP.9E,9f^dXT8+4J+(fDR<S326e8ZM#EOFYO)JfO[.VVM,JWS4f>(1<-:W^
<WdOPN:5PbU+Y8b:XOZ0\+NMWa&U7<X3F>cdOTa5bPFH\Rd,KC#ac2?]]>;W/g&a
@?O3ca632_\>&-(V?P0DTC<;.AWDG#Q\;FD-cbL_Z?aD:390QD.5A\B;^P:;gB\U
6MVIHV.g5.U;NKQ(-eHB=LS3eU>?U&3f/JQ-a33@2A]bGQ>dF;50</PH,1OH,-^f
@>GM^-SPf)/STMV1X@-V\];1OSDJO_EPQdE-HAP1TDE8;[::7H5PW>-TU[X[e/)c
\Gd@H3Ud.W??U2^LfH4Z/\/L/a32(L.(SC&\]ZcfW6HT7B:deQ8?.CSLWI_EGQOg
WT090&-\9WCFHYMSXLD#?S[?C_f9P#eN5bFFF57RM.-2WS,;WX8(JFU6(;_:^GX;
7\NB?PfBRU^TO?@&3f[>2d/6,,J1>\T51,D&Y>&aKIP?3<AJ?1]gG=JEM0]Z/\Y<
Ng<EEaQ^B3&0[MgF(_-[L+W29K<L4X^++R:;bT/@HZE]dJLf;BI+[5=fdE4Y;C?G
Z,JJQV]OGE,(<6:=b6XJ]JZ?LL+e&011TOa=BO,Ig5c[T0-MH\-U1/@EAd^MWB0+
)SZ#M;MU>&OMg5U+8@dWK)<IBTX:.@81+&P-8BbYL6#a?8NH@I+J/Na=&1#e_&[g
(72Vbd)Ma;)D(I]c_VBMX>K&?V\D>^D^c=3(203(N@_f+2VcF]BW)cA]X_8\eN;:
P;HB?CfaCe4ENFBPNP[^XTLeAI7CSZ9COce+:\A](N2+__Ff]^V+^J>\I64V7.5,
Ub9BR)Q:c3RX50\V8(J5XS?K^9:D.f9R\CD(?>X&T]DM&Ad1fLY_g]3P&-5@7&GW
/M>KT[_baI_Y0WCE<TI^F(,00YbUZcRR0S3FI[J?g_D83.D.B>U11cXJP\DL88C_
.NF>0ZMWN[/Da:YMf8_8JFR;Y6<8GM8JFQ:NQ7T:ILOD/\S#_>J>6:9U9M#D>A[9
CgS-Qd-e7L6bN,]\:@dJe5V/dR?3e>92(.+@L[-f7Y_JC.3VT):F(L7>A4.BB)BI
CH_HbS+cbZ:.9>b@^/g;9X)g@3[265=5dM--9\>-=H@1aX;54fd:AP^&d+9LPI\U
S(E6WN5fROe.26\+^(4WV;=Y3=_+MN2_XMI+1;KO:GO?GGN6<Kb]eI_6f8C0d+ae
&.a@0[19#J3\B@e\7HM<+D(D8_WXND)19Y&D[7W,d(a5L#g?Vg&^dCd@3-7:T+VB
C=2L>2@[?Y+R:NXXV8L.DAU]de#VS0,AKJ@A_7.-0b/.VgfV\@=M7-#[PRKfA-DQ
.CD(1#TLCTGB@)c;.DR9+[c80bWWbb2g4.bV8UQLBCY^YUEKQYT(9OeL2\(13g\c
R\N6IC1a]JGG[,5HTALWeRIIfRE1B0+]UI)&;B#QPPSSZ7_V1gCWPWFb#f\bN7OY
.1NNJPceQ15gTOM1I]?E?(BJL+FMK.#]+(eI2OJd5D>8[&0UQ_]:3K)^H&f[P)H[
EK@0/BXOV>S)\EBHI8DTY3SZ&:OV32S[IAUXb[]LN?IZ@1A1-ZU/(9]);_23_9<X
?DgGcC#C2bHZ3S1X:+J8WN6^Sc6V)/#a=S,_&:XCV:@<4M-Z4cX?Sb+;<](3EN:\
DeOae+AQW\bDJ2P1<O\5Q9;[7\cCIIQFN+=1?LXE]YXGGYA=RA/KJQ-O@N18E4NK
\FgEP7(Z]g;Q;@c+OdY(\G5MHE8Q8_g+5+c5eRd(NT#,OH^19RJ,9:>H1WGT1KYL
7Q1P?2b)N&7(5/-2:>[P2&#L0N3_IF^c\C<Y_b/b^cb(<T;?0M25F5-d(Q=<aPC6
-K0HTC+9]Uf+^SN>+<cS52gQ:0@8>3VY49AXJL-80#ee[253Z6.U.c7&.:3+AZLV
;^T2B,[=1Nac.KIZU&f0Of7,g?05.5TUQ\HCY6[G6\GWF(7O+Y@,#XQ1CT.ANWF#
a0Z8R106aC4g?@X:DVK87^P[aN8=)cc0;C/L/<L)H.+P@K.O5]72D3eK..db.dUJ
DZR]T?c3M8fC9WVfYDN9/V;\4,82cYDQ]#Sdg#f0HWC93/W7T2NHXbX<#ILN7,LV
B(.cD4UGOG&A39CK7<H+N9ORVfUZ?[;,7TXDVH@3#@g,.K^0SgS(P\(I;XY4g1eS
2U(RH_1D4bf[X_M_.dT<BL]AXQbT,QaO:H81fG[<YQFX_QP.-1,02.6GHA##TRPG
BeETV-<Md^U=Pc,UG:)XPaLUU9Z-.0;_7RKL(?HQC)/[2#aVcf;F83_SQZe5PN<Q
fg9UBFF#PHA8,GAXefFN6cI2BZOHY?dW62LQ<,+?SOSf/CM-=MWZ0K]]+>J@O(W/
3\Zd=6DN9/W28O3:4&RJ4/+ZZ;[&H#A6I2+Ac1,A-1TF7AK,D&I1T<,E,aFV#RFP
>OYAKgVFJ[6IfLDAH)OWRU7LK.Gc>QD87b<S(;c:gP\d/7JM]d7N_8DKg6LSYUS;
RS4:TE0^6CGS.gHaN[TKW0HJ,EKS46WNVbQ#=XI7?EFY0O8gNdKV96E12^&).dH?
_Hc[MZ>/+,Nb]@P(9Sc\[1H/(<?ebNH=?ZG)?;6(>LI9&YS2TN9D9G7G-TCb\]/Z
&T#N,<<a(CcQXaRJ@c)L9W1)U9;00&DL0#.TW03OM@(?=.0>7bX;P-bA<9]4FT6Z
F+.?[OV\8=bUHba<J@K-bM.KND@T1bcJL2JK(D(J698cb4U@4\;;.bB1GS.,@7\N
S^.#\MZE)E(R1#+(e>R:HZ&Xf8,?Tf[Z6Ub9+>3:J>OL)S5Pe.7WTVL1F7gQIJ2a
<2J8Z[5fU&:NE=RY3XZ=N1+B750R)#+BEE=T#1<C:+HHF9dEPHM?ZgP[bfW/6GWX
_PGTNRb3DFX7SG_c._bC&&566AWeM&7^]fUIT/b3&[+Z;/KYQ3?IT4,N1,IVOBOZ
ALMF?bF]11\>?7I8H=EBHU]4&E<FaM>11+S>UXJ_6aD)Zeg#EV.\/;<W?KcDaaS;
F=A-E:-b>Y-J;7TYE9+R7fEAI0R=K+D-&9QRYQ:20(U:dGMM<V8L0D[A?L\Pf3dU
];_E\[Cb>#NfNCd^?f_b36<7NQ)JZU[K;,0RdA>7P]=bMLXW0ZRO::7>S0(/@bG0
-3IJM<L\BN:?@>[ZFYeb9RQ1//L;\/>W8RH]\\c(2B8-ZE(B9-A05]dUSO>XZcU?
F0E]\O+;-3@P@U;XR5=X053&?PCf(+@SYFZUJ#?=&/T+Kb4;-BV_29ZTW(?:SWOK
90RM983YKZ>;U13\4(ZW-eN6XCOW@CYf5]#8G7Oe?=1(40)6SCY&U_]e_DV>A>Y-
1/[fHP3/;>-RH&V+dDU&@[O-W8dF>Z\d5(YFADLD0OY5X=f:/5FMO3DPX0/T-XAG
bOKU+PD2S-W7&?)eJRg:^):\>)JJbK1N5@2B=#;f/(BRETKZNXVZ.JH1[gYSK;CK
UF7:T41=HgBVVLA/e_EI:/\.P)AMEa=7X8aL8gcZZ<>-BI^^Se8\M@<Q19XHAb5D
9PVg?Q4(/J,_=D;fNUfU/?)Q<&aH=cD<bWf@T)HU-ZDd0549K#\9_Q8>WYF(BUFd
8-1U24<8BPF@2UB(O3;R3I,>M#3&EX@N4^;]G1L&X6^AL_f;,]1GFeK#UL,;8GEC
)cd5#7Wc354+;1X4a(71DV=#[S@S0I##ZU(^G+O:O5&R2^)H\CD72d5E3TSdX9@+
-1@X9U0XZS;Tee#QAQX)7HW2>5RBF_IY^a76(E+a\LUO=NE#KV^ZcJKSAfLS5D<:
O1ME@GAXY6=M/+10fT_)WBgLT-+S4BJeGE,NKYM8#-8(B>bP46D(TM,c,a>D5?:>
N+f>T9A0DCe@Q,e5(104)]J+VEZ]1bcb9NcdP6JVHMURgQ239(Z&;,\DSE=T?/?B
>7YGV1+fP=67K57f^SY0+_3KAFAS(\6e(+C^?5<da2<aWd<Y(R5Q;ZgJCa_?_515
GHOALAdB\dJa^F-_,ZEeHG)/:6aeU+\U(9>8&O-Ea8a4_XK.Gb?39H>W/&_Cc_L>
P:YDJ\>4CES+fA]7V^8Gff2U5d)R;VOBNdeb;HFFQ2CYaI?&fa;JT5e[@LXZbVR<
IP.S4D643R=>><2+CRDWVb9cFLQYFL37;O1Hc//5,.00aQb4W=_<1E:SbdU4(W8R
>Wf</7>ZeW70EPM,XW.E96CaX,)RKAY>AIW#ZAaJ(Fa^]A.]14:e?9VH#-3)V+7Z
gH.8<7V:>AT3ba^0J[/6TJ--12I7.8G_Dg,Z=X,gEaY8[3D[K)-LV-e?7.DC^_Zb
4-)T5c6MMWC.D.Q:_;6Z@1T5;>cU9;>XPQ>2QT8/361HQ^/1TNR;d6]ODFPKC;XV
4^W9N@>BU7>9O&cB(Z.V0QYO)PVE[PUZYe>b)e4[(d0D[)/,(D5J1b?:]K_Q;<W1
.7\_;d<5aNAdV?SJ4(5XAbOV4[VIabVQIEE;;^?e3OM@.23/17Rb;2D_#UG\g\HN
?L_A&=dadf4[JXf/?;T8<5PN-WdRK\_A5/N[VFc)09VF>WO-@dMAOO(:efe.H#?&
.JN-@d=M/KOAU(c0H[g+;a;5?DJ8)WN>SA38C#O@7V?WEeTHGR#[)O=cZ9=76&J\
7?]\(V_<,H^WP]D+#Yd)192a<4BG</LNe@J(63RVMd?P#&f<1_;&@b1M,b=S@E^+
KJ3ae?M:.TX8[JUK)f<></QT_D:_IF>7QCLMZbW2-=CA?W#.GcDL\N?<^SF+;ce+
\&bDP.EE6S?@VdbJ7+)2YU-Ia@SMW]<;cS,F@3PbG=H(YE=D03XLgX3RGbc1V^>e
Q5N+WL#R3Zd-0]c3V)TJ^)f0+S@Ta=O8P>8C)=NX:N<N:bf?R0PRY,XK3IL[C?QI
FFbR+=&U[ReXW7b7@H0NP&XbT.cR+1#:B0.PCBK:KA(^MLcH_aC@PA?be&]7]NAF
aW=>_3G?Y_(7F4Q#[V&HIK9BJC<39)B5WCNV3INEA/W1L16VF7.-=;Jg2=6]6eLd
^1O9M>X7VQ>4(c?O6F;T-4MeJ8V.\,WT+DW\F#-\09[=K5]M[Y13W)U1,D_6VK29
UE>g=3efI?Ef^K=-QgD+#(QFGB\5_-U.<4g+&)\&-R4<N[@;cBU4_Q],GGTeB[-K
?Ee7:SS2BKYBN&[9QJEPIYHJ^N.O5@<EfYe?-Q,?R-NR+DYQb_Na@.=4^Y4TIg_.
<4?WS6I[W@2F?f2eKcKfA\g1=7+:O4@+AL-b,C.;(?)JVY]95H,M<=4,/[?Z]g0.
-CT-E5d/_MZL?>fQdV3>gKL#3bX6(G-3_7N0INZbE(.Z:1H7#<GC3=D0KR\(60A5
_g>DQ-(#IVW2<c[5G+08TK)V<3UPaBFF@:bKdG#_2SVFH/(Ee7;MO8H=Y<@:fd9>
gPY@,D)f_I,5-gW(:FI:ZTK6bSL^D01^>Z;bX:TYMS8]D,Q41A&eeISc7NbY.V9O
92#fYKPL.G5ZH+a4<5-,OI2BabKF7A)YF8aA&&PPL^>ENB0gVCWS3CCa/Q+^.HPe
N0Q].ZOgY;.;8RgdKb83EL;TX]G<cca200:B>N,4#Fcf>R7^-D-7D]:E9cfFRH2b
Z?M5RK=<SfI?LV0UU_#8F5:4,++J[?H0-P]4Kd+-.U5=LgZ#aMU1YLL0fT)YLcPd
gCM-27]&/:SH5?bB;#cF_-eXX98;3E^J_[KT2b-80SI,0F-?T)+6gK^9b3KVa<MP
\[=H9,_cd3^ME<H\P>5QDO.;JX<1f>TL?+C&O99gYL8<BXP-EN1;ZKMeGa\1T537
[Dd(>#9:Y7I(OF3S/T8=VGcF>V@@?SE4/KB;Q7J882fdI):fIY5F[N8@)[NY?M-\
TBPaQ@fQF^;:Fe/6:S_A<BG#<LFMDB0R,;.Y)OS[;fLd_U1-:RFdL0S.5H<3&5OZ
S6(1a[07_6<0\_SQI:VK&49D>_39>6BJ[L/NN[L;R9+U&S;)c]1Q@5XLJ1/P46[G
NX>85[W2Vf][D^3bJ36=b<\T2&V,WPQ)TDeB5+O.N(-)@90d6\@)FAZNZ_I+.Z&2
:4O2HGD9)]@QF;g@9TE_;>f49KGTDH?+.Z4OGL75Xg<dd-#dNb89AXZ/=Q24ND20
K]^F^-:K>g2A_)766JWL_G<e1<B)1>K4SKP<.][CCGHI@KUbHeJJF8?<IOUbb;-.
88Q]BB]U+DR+-UA8U5:6_U3dWYJga:/9,8c-2J<273@MF-QOK>.fX113M7=+(2+D
/Ca=88_9VW;99VDDLBa+0S]SGL\[e5L[D@Z\L(:I0^3)?F,[#\U(RZB45aFSK,NS
g#+OcFJEZK6:XW?b]c^b6>eg\&cab+2VVB/3WGY76==SeC3Qc.EQB?U.e[=Ha;-O
e2)+S]?V<#ZF[NPG@GJHO7Q99fM0LTb=J_@GCA#K7Ne3/5CR5bV9U?dI&ASSJN@X
C+(V(#8Q5b4_=J+f0WTU]^[VYAZ64&6]XPG?YC2:[SGQHX/=<VYOU,9SC.57M-.?
+N+.^+T>I>I-^ES_1YXQ5Y=a^]7\:F^_=Q(_<572:-6ZE@^Q&+(<TB&:d/=e+7f&
M/L2JH?H,KN0IE,C[_X67EA)WUW0f/65PIRGcZ>[g>e7?;[F;ff98@OJ8B@>EZG9
_E^F7K/DbWU.LJ<3gWGb42L<CYT>B#gN0:[C>[.],(gXS4IB_703S\JDfa7/LfFA
#2I@HW7b@\C5ef2)DLMUFJZ6P=(_g7?KOL[BT/Bf^/.V4bC.(1DNVbE+SFRY.;+W
=CL>-7BdU);SID0-1@MC+S<&U_&f4N_aKcA[(;A+/+C4UD-gJL8@XDU^_8U\JNOG
U]68EPW(_CL_X:ET<UVdaWAFLcN?Z,WK)OMNS2I1P1_#c4FC;NfdH06d/?BO+aCV
M&G[aMVL5AN<g@ET3T3aaIYfX=A/B&)-G=.?WWT@2RVC^@+Gd0d&1^<7?2>)f,3c
:d;]Y9aXAJLQMUNQHL-ReR(Na7HbXF2)/>8EE[0PJfN/GC[T^</WONddS&/aIR/+
O\B_C][-<95g>_HgKAa8T.T.X=V]fM,3X2&Re_P>_QSZV>g96SR7(=[C@PL0>BeQ
_G\?DU[<)c8/:Og]WWS#=D)8V_QdeaS;7._N,-K[f=9c93M.B9QH;R).>^9HfY[L
B#a>_d1+)Ja0a0OW&S//I.8O-Y/a?#YZcX^?8_R^I&><=[9cU@3)U^DEL8Z,EPXU
?HEF#Le/_NB:P4U,SN9CV^SESB[Z27#)UT^+,A-.-a6OV>b&#<.C,;ZNgKG0S2::
)FaXS:c4]5+GO#ERJJcZ.D?LODDRdUC^RTS&9UI4\fSA]#TR8?G[>L^Ug>AM\cg(
Ra?)@gML^L<bYO[--Ug12Q9(C4@+2PcbfcFD=TcD.Gb15DR,D1>,I8:&:)>#J@K]
[FeDXSKdU&fDKP[6/WK@3?)gZY:Y1;IL3/-?WFfQ(VXe#Z?M?WI;4_IBTBI):KHI
W_19fJ_b=EH9bR)9#M(QZI7RYOAETdG>TZG=Ic&VK^\dJ1U]&0(;#2@0Qg^-PL22
WCK-^M@1g^N.J.CA/KQ_DBR]@DV+K--843=V#JLYcO.IO8:KZ7_KBc#7K_ISa-W<
,A>)#/YY&<:PI7_;18H=bVeS5GJ,G1(a16:DLZ[ZW,R]LF<.W?fdFf.TP0UHQ-J1
@^.SKX6ERE/E[c:;1&8+.aCgY9N9<55VN+5#H#R+O<W+Z02g0JL#gb9A8V-cYG<5
>9WPTW0a+(.VgX6O?X&HDHIcK&eaE?KB1?EG\,2:g-_cg]DSbAZ8?.J:TCC&U]J7
\5(.K9f]^?2+1575ga#IFIG9FL<3-eUI5_F1C:SWdVGMS]@e->MMLgVP<KOET.CU
OEG+d(22A\bS^.-Z36c==-K+91K2gaV[6DML--7_f<3gXFMY(CT,7.b;gQ9SR+,D
VVU>K?^8Q2d;\8Lg8G.F9E3HKQ9;:c=c20d:dTdHT<W/5MS1&f?F0LA\M]T,MRPW
3^+IX8@N9F\?8B<f_:d0JdTU]IF1;J??MdS#Y+6D5T\(PG7:U0;WX\6ZE:&\2Q]5
=E5^L5TK.PFD;b0#cE#LB@YA)HaBWe5SU\R[&;=/_<P?4/#OA^-V3[H[ZF&G[b@3
=L;dO;:FZ?V0?V&K)@459;E.5Me,)Y>U^OVa4?IbCYf2-I1ef@JVLY@,SaR\TRM?
Gcf]0(&2c:3<HY1;G9KP9\7=9JQVU#d2gDc\-F<8T(/^:@b+QR:646IF,@9M2.&P
ES\0R8[T.UO5_SKc2,?]_-._D6)JBY<_K[>=G:3RE)F6SM2DSa5S:TE8OL:D4X51
^/S0N4G=ZbX7/(0[A]WP(-0Z86NcJ?=GWc@9:12E8#IUQ4U<CgRc,H.)79e)C9:@
@1.F6C9:XW.@3,1BPQ35aSE5V15_E/W2Wa.fY203UMfRF<-&N54T<;](D.HcQ935
\V5R>2(F:TO8@,,(?cB^)AWdbLc#A,OV&Sb#Hb31GBDU2^;b@KdP+ECU3<5dQ/KP
GS4Xc2+Q=)R,V8@P&gLWBPK=0/\WW(eSPO7Ha=)A;P8L2YP<>Ia;-d37C\OE<9>\
:)a(dFK7YD=Kdb0K&?/6[e>KT(T=gg/_Q)[_JY+MXO7#OHS2)J8Y1(SLB@<TNJZN
dEZHX@11T_Qc]SSO(^IRRc7=:/IW(c]5.\8FFH]/UdDL3L]/D[UFX^@+_#D0L-dK
^/F#&-PJ4\67&M#AacR07COAVT<e&\d([^aR]&&^N)XER-.e81?,b.PN-dY:#0=D
<^TgTCGU)-bJCO3@a?Jg[D<H[].21,L2SFdD0_B]@5OKg]4JMa6.7Ub,H2QN;e0D
>/8;3)?bF3QbQMNT=IMUcA7aEREZ1J]JSJVSf1fPED/e/LQX1Ba72\--PY/V]@=>
O3Q+6C_=1T4=X6?]_MF@CIbfW:3<][cTS/@5^.g+?;9O:H]QG</-XM:&\Q]d\^J-
#[5)]E\#Je+G6VM@:^6[;LF@,+1@QAL@>@PM]SN].N&P/c1a3.3TDgg5IV3b41Yc
DZ&(M1dSKI)]GaZd>#[>-C[_P9<[7K3gWS(R\PW-fg])<(X:J-/RDAL5(eS8B>X2
&Pf>R29c^9HVAT(3?9VA76MMR.[CX_9YJaaT&OJ;8&]I^e42&O6Pd/d)NC0@UQd_
RA&a-a,++4)PWf7FS6A8cV1=UID)Wb=e3WID6=>VYQSbF2^Z^+H^H-/4^[&(Yg2N
6#GBdT/GEWQL@KJ583FRLfJMeEC]5L+P_/JG>#JN6-;0[6MAV5-Y8\+)Hg^cffVB
.GNV5UB8Z;=?6HU6XgTBX+<S#8g2\NYb3BBfS-&=aGCB)+P]G1d+)LIMLa&I2UNL
=IW/A^Q2=P4>,5)6PP>a\]9>dY,8NMGD]McA]d(G?BPJV#YZ+/JfOG31@QW@)e6D
38V<,^ZOGVE):?)PH<:1]9Xde2F_]J.c21QgVBZHa^g94E<dd=Y())a7OM(<cbS,
[]BaR/N3cGKA4O>bbC.SB+WR9NSG<8PN3>-@g96gf0IcTHJ5a:7W-=CR;X0UcO>0
@7a(26fdP)2-A#M?_g(6=e#EO3DM<((VC:dQZ(c33F>8AFAHT__0a4M/.29B7>_S
;(Z0K9Od-#SS67RTM7+2+UY^AN[@7DM\85XNZU1C5@SbbFC)U3AdCE52Af7.g>#J
Q-YFf8Z6WcJYSYJ<#LJB,?=NJPd\;#ZI=LRWTCVbY?4:BS#-_TO-CW;5a8MaeRD>
<Nac\:<DFJJTLg@e3J+\FLTCa[PT=#NEaVgC=JYg1OM_7=_Y&3KF6[]_bZ.]0\RI
-)D4K4N+<IE2&fQH6X8>L\-L-VB=aVR>Q#=_.2L>#J1g+R[_Z:S<0UED.a4[0F>S
/3Cf[G4N6Pae(O2XfV,VNHR&@c]SR71IG=S+0WOZX[UdG7V4GO[-IQ]ef3^AcGZF
X<1V\;Gg^N]KJ+cP\X@dT)W115=b/d,_?VHWA(9B\P+3IO=#O-J4H+0,X4\-7NE/
C<3.CT03b8O7@B5L0L:>FG=D2MV,V;GEU.+4?]g05MT5BD-U?;6S7L];cBK#,#+R
R+RFU99[^KGLQ:SQU8McKBL;_cEL5Q<+_cT1M#OQBQNfW;>HXTQg6<(0gQ3QDVLZ
-^#c9?^VUI]/RFc=.gAC;KTa;YKL;d):H4_@OC2>A]+<A7fAQC.IJ;->M4(&S6]a
^#g,;&QUe&D;2_3>#&Q:-3_&J=D9>a[R3C0e.5(g&TE/XP)U-\2V5RfC9]ZH\6>9
+?<a3Q_/R,+Mf)14+&^9;0F8C.#.]]dgd)Q7?XF4,BZ@INdAJVa_UND=)E=BDG/G
J<,QZA:eAaBG<&Zbf?SaGPI6P.0=2[BT-#+QXWG/1cX7OG-[:bU@AW.:G#B;MQAB
ac3+GUD6DM[SMfAD3&=O-ECU0-1HAJL-4a.GOJB++g;[/?aY)1#K_:8IbWY2DDBP
FC-b^<SOBA,VHag46+(_0gIe6RH&BZJBT(D+4L[TI.U-S<4+E=BX/&2VU2Gg1>ZM
6W.c?133E-I6U_@Vcg;eS/5]b)&cTVgK>&E9EL@E_U9]_.D_#Oa6SBGN=QNU<;08
=RSO3.F1)X[[ac?-Id4#G:a,46,g9U>SRJTBPOYCd)X6A7.44dPSC@6(5)J<;,a.
,c/&=7Hg<D\OAfICBW>:)T@T2OOQ?LA0V41Q3aLT;+2<bYM-#OF(N=,.b3eUcSb2
NK]=aS-fT-DR/N/61C9-I86Wg-MT7P?fOD<;0--+QcKLHe^H2HP)C6e3T\1:XI)/
[bBTFO@NHE=b3]1,E.U[]1,=QGH7OB#V#I)XdH(8KX;[e6CY3\02DB\-M1@/XPHW
.AB+4I\O=[S4ZHG(I=OD:gV)GI];:,Z-JC1J+@ecK/BY695U4K<NQcFUf)?b.Y_@
>8,F:5#O?Ud@VF.PL_Q>.4OO1>dB]L,K1@U:)CGR7VS\fZ3(8Y,:Db<50_Z;;bB-
N^_R0NNW^4Q#Q]Sg:b#[8-PL?WC\>/@a78=O),2.begK2eIS3f8K[OM?gE?;[[NT
aD^=SULOa=UV&ZRYfE4@dNA3^g=)Fa+,5bR.WCDC5bb5#1Z#N/UWI;9DNWC6Wc_;
X+J4&/b/?g;[_.Fb3&W_.JBY[-UI06>V6a9)#cBI@SVMS?+V7=TV5LV[V,Y/Z\U+
6Y@B_1@W0.JNILN(9]f8?>?6@+#C\NIHYNRS/OYUJ?9HcRV@;A@f55gQ>U:XLO#C
06[/H)d0G(MB1f3+9PBLH:MTKX4f>W.>U]X_+4BbEJM.-CAf[U].)5a:42>8T93;
E3&W,KI2,C:TZ9VAKGgfF1eU@PfIRKZA1H]ba=[8+Yga3;P\3\EH@5RGP)H)5e[W
W,CaY@BBV1NSZR+J0A65#b4^0=[BPU]Y35Uga]]K2(0.J\+ESe=,c0I:f\4908,D
;H.8HC.RK,)3OPHIdR&:>]G+RfJ(gZLeL(cbZF,f+YQ59\APB8?GJcNaJ;4E]f(5
A7R0f\\?9#&ETDPYUbQ@L64C:Z]aJ50?gO>(O4?f-KTYHK2EP=1Mb7QQ:,C/NB7F
7NH3RL\T2@.L_9,B\2F;2;Q]VODJHXJ]UP[2@)bDXWH7D=/E9U;/^d.Q[A(+ZN_T
KMOE]VW1[Z)?\5aNT]N237V50^:-8Q6:AgJ4\a^U32Q8C9VTR.\RNN2XON_Wc<:9
8W[cUY>]3Af81.#F1.>Z;GI0EJC0LJ;Fe-R_J@c1O=^JW>0K04I]0F83#=B1a;[>
)dPTf5?IF:QX^<N.+/eX/0=6R3SfAJC6bG\/4(Od.^SEfF1[/AN]C[1Q-1)>:J1N
<a3:IF9[ZC@??&X2YUS5JR9W(V/>e2O(/4.IC^fU?&JD+2RL0VO?Ja)\=F)7#-eN
2.6X@((JC0QS#^8&aG]J2/?)(E+W-/NV17)&1EV).Z.gFaP=.T=fU(NM06>CL9E;
]G1KDee>CYME9;K\&N)T_fA7?CO9GH6/;]@>e>][WC_F[2J@12L)^b\25MP+(+B]
63eg)d]<]J#K1<I.4,QY>Ja]R>EIA#0LS61O;F.X_5#.#)_N62YLVVZDa,IUXe<P
WZ(cR)8:1aL&UKG>]OBJUF[91E-8]]MJadT/V&;L]=NJ4PDET,d-KeB/O>Cd\/2&
=N#._J.MHBCQW[(A8U6?,c;(P+@XUHU6CgMMS[/WUXTC2V2&0(ZI3RNF1Z^#V>YT
6\WXO^6_B6f_5GOYI]L8dY1#WA8=0A3G+4-VCUH(>M/fe.gY?,D=)2dOVb=]4]UP
TH48O<ZgbPLL2#.:<K@/^O=e9^L(SbT11]-W[PUbZd4Q/NR29CGXFI8JdZKB57_H
KF=TDJPUQ5<V,gR]8JC5:HV/=f5SdCcJ8.JO#fJZ4@.+cF#P+.WNLCg02\=?XN0#
KJ.Ig9X?K.8\2AZKa9g80A1U@DYQ;#-V<CFQ5W>?)R)L<B,&Q2B12KUG(1Z7ANfE
E+JgR+5W4F88,9>.8d#>:R#FR#VT9LJKH=ZKX[4><(IH(f/KJ01^1[>Y-+7&Y1Sb
f8;./BIZ_YRRUeV#77I2gRW9d_NfCfLJ77N:]6e=b;LWa:=7c2=CT;4f;CV.OA[Z
XBL;fYVY@Ua@+#;I7+U7I&/F,54FZ<K>4_7cN@#\_2X8O1?EMTF6[#9NS(OC;9:@
I-Jaeg@Xe?7OZ,0QS/?f\f=[?&E;1[aP?K#+;V<B#:\gbQ#L^aR@7],@-+J;Kg^L
C(e^@==S>N_c?&:7EE@SHO>P=FKM+0b=4b3AAGH,eSJEK54bJP4VFRJ<JNKGP49/
(QPQ7L7gP9\4DWY/ORG9a9^32DKY^aSK05QVQ0=^A)TIC2?FOHcYTV0b?CbWE=J5
^[<37dL+c[VY<L<bDRW8)fOUSNFJT3B)Q,1AK<XCaD50M_S)e]CML2Z_Y\@e0V6I
8E0V#\EC53]JXRLL>_=<H[K9M&BT+W[6BOd8E@FMd(1M9B]U:aM50K<0_d^,GP\P
X)#,6Ef11a:38DTWE=G\]1N1X@FHFbWHPGccZagaRJHcRc@+&RV.GY;K(ODf^2BL
49EKMZ8Rf8>P,&J[1;;V)EJWP_I^;@)]e<W0M>cd1g.U;Uc]SYYD<SdACODa71O:
4DQ<+6\</;O=]c1L=:[DXdf\&1XQg+Z=Q9:8]+cVCQO[ER4RMe9H]IU8Q\/E>8c0
ebWf^5.dg#<W,-[@>JU,UI.FVHBY@Sg,[&NECTKK83Z>J9)/Q+FG:(b=EH,A\OJ^
>g(A,8/X:68YWMNE7?YED1-&/(>L=ZY7(L6MAdXXW\C#f=f)7bB(S4EBM..)&_E5
Y?4/>X?[3Y1;LQ8NU4geY^K]96T/3a^GDA^If]F1fHB+V5U;O6VAY>N]GBc\+aR.
eSS6,N:1^9f(8(]Pe1I4(H=CfX,b(_Y=-D902MGWDA-SV&2W5BX#D.Igb-a1La)\
ef##>?g-@)VMR#8<4ZE@Db^Me1H<)B_3+HI@_G4-A_EV@HJV8U0Z+N@?C^J65LT:
c3)/OK,W?&IR_.]-DBRZ,[K3GBgJ\9_#P?/bV4Z45UMUB]c&8,e@UF=f,RK?BUJ_
CEP03/X>L/S/>1&KF5QI?(TZ\\gCNHWZ\^W0gA87ERaf2B<7gF+2558;KeKWZX[5
<W6]8/MU_:W,.fW^,VGT4H<c8;V-YJ)BFd/0)WUG6>_KDX=b65;CL1B:7S(Y3)D[
UT1X0I3PPU/A?@Q;(Ic8CRcfeY\4[E&dTW=RPT;B#gK)T7F,IOO^bCU1c06HJ9_]
d;HfZ;6HYH^;ALK0843.UXC3)g_PN7#=>#S^\gE:DgZ;J29M1+G&SF22B2^5]aF&
J&&?W\,R:@L13JB2WV(\a;EC3X;LA8)77RAHeEB9)<YE/R,)]b20e_YKdGPbZH_c
[[d</@^H2X0\R)W5/4C/?NOJT(06_GH]P3/W@(V_0YTT@Zg;U)U3.BPc5T#KDc>?
cM)@b;c],e#5R0)AgdJ)>Lg1Q.=P]86Z\EWUR4ATR_3&Z6H+K4&)^8,dBbER4^^S
4QdM4&]Rg^7>,KN_^XSRD._NEL&/cWO8>.]fTKLT(NO/OM0K7ee/O5HM;_X9CCPf
^g687E4+K0Q(5T3cM\6>0NBH.EV:582N&>aeP720/RBO>^6^KV4?VW,GO;B,_7(7
8ff<e24a#\3.M3NTM2a)4g+@5Y[UM#+JFYbS^^#IYKDZJ8UdeCZ_I,R6R[B;WQA4
T<0d#Bf\A#7/E6^6=?MgDg^J52/JLa+B82(b?2-5AFDDBUO01/A8dSX2<CVUJZ.:
1.J>=B0-3/D7IW?Nf9=JU115Vb0O:A+Z;D4^g4&0+c7DO0Ue>3\V,MW4,bGYe@L:
<S#(=_<7#bASge?<#704@Y>;PNK[=:A;T]8#cK(QV;.;[0:3XL&?>bHA4T_=3eVZ
M6W<;Q^@.M\.QKN<gO;db5(1e3aP\+;<5S:)Q_7;d\RB(effNGRALU5Y2g,ZO35I
YHb=1;9(JB=J@:(CEQ]/FdSbVI-,_T6QM-JMY>@eeF>;OaD&V>5SX]IF+83<O8D\
R3778@1VUf&<EEQ.-:UR?>L&<_DE6J28eG3_9(4+FV4&M9Ca+/-MT&Y6-JO1=Y]4
2]gYM+F<LS3GZbU+)c1NW-Z&XDdG:<\2Z)N&cXD9\^P7I-fP0\9gNeEaVH\911N,
-ATg52=X/IFLPW]7a_-O7^(;3LL.CaKKGgY1C\[Ug[&VHT0,H0VITBM>RMW@H[:X
N>[U91107O@KHgefP#,ad8FGK=a[(&b1TX]9N5=.TC>WWPC696,@:V8a4?,C13^]
H@W8YKERK6gGaG2\O2PZ?AT@f^g^g&\AHAe&._#7)/b>=KW4Y))[ccX,:EHFSQdS
=GSS&AJb_]UP;Pdae.c8d\Q@;/@X[b/LGYeWK.dGS-=F\DOSU[XUKX\A?B/_W0+F
?Og(?Qge&;e#;A(&b9C?WOL#<G8fOL/5>4]H;Q3C3F91\Fe]d#AZ0PGL\@;\65.E
_,?RgCQE(e/+@)d,283bUFMZ^:(Le+0aN2U7CF@B<AW<-PZDN(0,b0_6X:#9&(GS
AL]OZ(<=3<XBHC(V7EN2dD#)D,0AC+.BP/+-:CI2Y]G,,GHTOe6955.73U01=,&Q
Fe3fC8HF0&89G@R)C&K\)b0F7XY8VQY83eAc[c[e&NLM#P@>g:ONa<#;U2,BUG33
)5::X7,edI+99GG=e?+J5K_.?=MHMeeMFZHK2.=(LQHfA[1K]N4CW<M\R[P-PJI-
e0^A]@g(F5.]GMSM/cWJPE65,cAgMK4K\Ca(-J_&B/fMJ_>dF94S)ae,9DUbW-d_
9+B()-XGTUJb:445--75WYXY]1WE?#7N]?A3<([PRYNdeLQL=,&TN4>3^)2,YN1Q
G;fC139=5ROB,Z):0E\1KV9J7+).7\LR>=4aeb[:g]:U#C_H5Y7RU1N5>KZ8&B@&
Xgf6GL7O9TS7eNR?^K#d,,a=6+N&#6YZ3H(^QNT+@+g^RB4fEN2BJc]O/2B^_>AN
Z\88^=6=[g:Ac?RF[5RJ&J7KcAO[+;;YacME8WcJ/L1]5LFJ]L^VU?b:\Qb5<I?T
7f]F&U(Lg_?g7-1F\VR4U-Y3XMW24L:f=cRYgA6@-C0;]MGMf[E<HGaO^0IUI0+)
C#?_fC]a<LFWN@C:D_aH6WeNO)C41WJ(1(cU])54f_^^+\EU]DLM]V_,57YL1Y4R
,#^f_7_V)Sa;ETO_&HAE^deZ8TZK1,.^?1VX-EN)74>=,Ya&,T1,[>AO)::&aW,D
91GPdXB]7)<MJcYP07b],:SK/Z.WP_e8Q^:_Z=V3R]HJ\WFK[7gZ:@#;/]64[9BE
)-:DBSV\P76C0:5,9,09/^21C[@,O#DN._NfU,9(C&FGBK3g8O61a3Ig1.]0WL#X
c1T=;bKA];fOcN+P,J8Q&6CWHdS]1e.b6/#,&J?/2R7HKVG#KAG>7=5DS<cfRF7S
=&d5_B#deC2cVUb54ZC2M]+GCFV5W-F;MEXe1G-AK7V:bR@(MB>T)L:TO()-N@\d
^6a:E37g?&Pa+(9YJPRE1cGPC6B2K=FZI?Z:4+bNRaHGME#OV\+ggfa5D;5&A-gN
75b@aJKZ1ANS/ZJ\L6,Z:02:1Y+KFSVe>>2FV3a<6+C_S3V?aSaT))TEA[())M]4
aTdVCMTCCIZOL-e+PFG&CG8)T79^,-&cdg-+0MB&MNH;Q>)<6Xg90?-8?<.+&3(-
[K:-VQ?9HgOZ-&?>M1T)a8H]^E6VSg9:aYJ1?APN95PYa=_eL[)ZAUH@PcK1#.1(
<84\-9>EB@@d#eb:JTCN;Q4ce_@f)feK[#T23RH^0[OL)_a&Qb:8_</<CXba#@2V
g9\)+3#.SUd8QMeXFYaK4d-3C<PJc@b4@<&]#+/fQ?D3Z;0W(\:E+V.GN0gCF=gV
46QQfS+YT?RR#b2/C_eTSeRPB2(d]#I_9\F_7Gf@QRaBJ:cG[KU0;]fW3+SQC<,c
FJ13-UM3;5H55#c-a.dW@[_.G23A72\+M7SRe\MRI?FeRD9L.48&HO^GE+gL=MZb
Hd4X5HT2SMK+.A]C,&]f,G2YJK?cf/)SEcS5TH<a\P[RM8L6gO(:RTd-37)\6(O&
bZgL>?:#_:MM5P+[T+N.]@@\XI[HDQ+R7cJ<X]d\+G[H75CUQ:N.g&D=,>RW\Y(.
(SRg\FB-@H^U&Cf1^,2Lb,7g#Vcg3X.H_:QE@G2J^f#>G\#O1#KI^P-D_H@O6FFH
HUE\7,R[421ICV=)DJF-6N[DH2D/@IR-2gJ,LYO.TQIY/+^A(<b^HgIgBVDP6gVT
AD^\#cLV1Rcd5=Wg3_5U/8=>:b/_+5G7JaeJCD7N>Jc\C@U7-\N,^S\Sd?:U,[G9
5@CgJED0f.AG13A,CgPL(MdQ@SCKS5GE8#7Ma.2CcAb1A\+[8H?J2I)db;1RYd7M
.Z@@3dbFXXG2G?>:.9d(cOXQTDC@V\6K-R]7-3dVeCa9@1bS>B43bbN?L7JAaDJY
=#AAD>8BG)R1FP32d93C_M)c_Fg>C]YgTeaUd:6)B]J-=_fXZZ?ERD>N7ZHGI.C&
#@\\fM\f-N_HD(S?^/KHX#OR2fc/,##X?3^5gIPEH[_>3)P>e)g[S32)/J=[9NJ;
:bA:Be#;XN_3J\R<OYe]=;1VYbP]IL/;YCG?7CS+WEd>]=N@=)DeXEaY8)T0C&)P
V7\1Yg3M+RD?VN8f]--e^>.+QMdQE=S6,(71g5d[=b[9JFN-W.MNDP@ZHfVXcG61
.+HF\c#c50]:A0?Wa5(RMB-L?X2bS3N0H&ag5IcFf7.Q#TN1f]Z8D8KSN4f\D8I5
LDf67\VL.f[Z=QJ4SbWd,WIZSD1P\cW=OS36R.XeWA5ba\Y@(KAW#\.?d3=WI\\4
W,EI_6.FY?L\^[XA32>(;MZ=dB@Y>/e2PYV@K&M14Rf:/@M5-=NEE[@/EH<EP;;M
];#K@C_@eO4P<\-SI[1+HV\D<DZ@L.9N.0Q&+>HV\+ZJM:B/bL8B1R[7.S_Y^F7\
Uf@(a25)_[1&8B>1=3>M=Lc=MP.B;44HP=+AGM:7>#W&],RPA-[=B7<fB7\;ac,]
eD]<([Z4#54GY@@eaEfQQUS]K)X;.(Kg.Db&,MgG/23fBWecbDWa,^^)YN4P&ZB,
H)SU(f,ed(2AZ9P?)4aT35KGe;=-TLV&^+M\eU+A#d=@L><DMDF=3NcgTS2S/K14
<^H]WH^ZV\)4]gQ[&A8O=Y0/?A=2]2Y];WDb#G@La.eYU&=6DIdRENg[bYRdBK=(
=B7bG.M2,7]GgHDKZe0F5K7Y.745UXKeJS4(^?RB]6X]?Gc2D&?TW^HE+X9M?NB#
(?:c=YP;.M]8W(&9A5NL?6b7RIJW6L;QX=Q)cJ.QfBU[]QSSU&)E)1>PBF9(Kb7&
4;;DT&N?7A\3b)b4S-bNa#L#4T6f?cMa-S)WgATE6AEdedP)9#Vd<2I7e0e=ETI&
JZW;?bE1-,TB/(9gP_Cd/EKQ=^aC<Z[@&MSGReJR)AMfS[;Gb1ZPPVLDB)0)N2\I
P]=1JcRe8ZKIe>G_R)BPeCB<]]5H-#\P?VL5=[?70#^J.FVOcE1FQ2;CR<U61[T^
aL2AEU_dXV;]1QPI#=I\/7;-VadQ/8/g+\0:Y(_d.G+=;]S6YZ7Hf1VbT&O0=[Mf
gJf8_3)QcAFXB(:KbfVBV1+ZBe+3I5gPL/R(MIDSEXd[;(+W/_UZR=6IR>6La^>:
&_53UKSC#P.O0J2,N-3V7Af2-8P:b&gB^N048P8&)_4:.P0Y-<Ag/b]0/DXMX.S_
gd;ES]Y.(R2KJQ&G:P,4PC:;B?P(Lf.2N(LXeZ(>S/RUJ5UYeDdc#>BF867??1Ug
Wf>?:)>FJB<dZdXBL_S#+]-)Q05HSU4<2N\4^<)9)0b\e\BI7)?e/@7d\I1&K_A9
(-@8-?^M45bdKJH3[AGbL7bg0=g3Y27#<FKZA+WH@T\M@/?#IcX27<;]282JVFP;
<f3e-@E,><(VS8K&f>]Z9dRcg:LXSIE@>6QUX(?OX^GG:cM,;J@RLF&./#XLC6KT
DS(IW4e8,:L9b8eB][(MROW,a9^C)2=JK-_QWgZ2;)WN/8^gU9\40cV3]3Fg5QFV
G26P+dV<UcJ)4X5ZNXeFM4L8-^SQ,Q6b&L<0E<8MYBcd^AU3QO43a+9929?XKVJ6
0.E]8A?7=+#BJ\[0?S71]eH[0BaW5:7[>_FbbKCH<@510cc&3@AO9.)MZWFYVLUH
]DIK6V\/LR-51MQO6/:49<3aHXYD4#(;_(9[Ze2)Mg())B.S([S1D58WN/N4A9gY
2.TTB5d,)Y-a;GJUH8TI48PId#b28JHfZM)g&E)(Ke0:+9YEB/4+A?6?=_W,6KNT
/GJI(F1P:GLfe^<GR_\,:;X293/aA2^I@.8,+W]U-TA5=<<eOPBe<gL8.QbWZHTE
/2E^022Q?#Q3I^TQ#a70b+EAY(20.TcREPZe5XF:K#V57ZF01a[XUX>[B#VEL1T&
GPPa&LPO&MFC[8Z\LbVY<J1Z5\A#BgDU&86BGX6HI(]GC&_B)@P24?_80+PD:K=M
[;698fI^Vd&1K)3.>[#3/G5aB9Ed,\2U:+MEA,\,?I<ULZ,Ka=_(2L+7.F(?F9#V
Oe16d[@[+)ML/5\fPK&J3J=<Ife&))3dXT+3HC#4X<4MN<)d;YI0IR9f8S2\&(XG
D@E<UQH.)+2]&FA5YFfV4YCO.JLS[.0=H^03.YOSFZDQ.DN_5R:U>)6Z?@U?fOHM
65&(^dK;4LKD_E;Z]d3OfL:c02dQMAE9OcdD?8U_RN5LW=S/&G2.9bMcRFY8-V3?
O3cS(V/NH:b(ee;9XAE:W[_D5B]fYdReLXI9fW/4gC8(B.I^KM0Me-/CEY,,QU83
&(#XY8\Y6<E?L4&gVg)K1H,W,;fO7=&\dgA#SZ2]IG<B][^@O85g&dbDaa>/_UKD
DA2PGH0M>):/>8aD9a6e_GbY],S;SX48]Ze+8?NddH([.-?)<\RU0FfDB0OP1M11
Mc].1g^7efCTG/)+B^U?9R).KIDWSB<<U&WMW8R_4YfWH6<:cg:Fc7GM).<5g@QR
e>/OTQa>Pa-)SI\IUH)92_RZ&E1-Q0_;-\_XM4.LU?L#LY66JM&;RaB(EWdN@Y?\
^QOA<>P7;4XWUZ2\eM@37?Zd;N0MY>71KL=g28_(\++):/-^B[;L]MR+CIKF@HQg
O25\CYE7#\YY<VA94d\@QIRY5,e_[5?HIf66HH3/#]GE/fG/cN1CNC:++M[#V5BI
G_bf?QC&3YV[JHK\(QBF,W-d,OU<(,B-Y3C8OY+eI^LBI::RZY3/VBI?^-47X\^J
g&^^Wd9bR-;eWA6cOeH6.&BO;:2;N7AC<\:H5G(.ff-5;)EeE_L^5R8<M,X4cRL^
\1>fKG4^084;]\bQ&Tc=7GR?YQU;T<Z+BH-Rc0e:^QB)f4B;U.W0e0@;@^MTfaAN
.FH+FfdRBIB_cLD^0R3>;8KN>d\P&J2FM&UQ_MX5Vf#XaegUJ+0418AbDQ>ZN8_W
1O_7WQ<.^YHX_.3@OZ<Z>#;F1X875M/UcKMBH@4L=5R-8.ef[ZO1X1UdYU[eHZIT
DNIDQ.B,(F;dJSS1eDKP#<6Z5\=FZEcY]XK81Jd(@?3#;C[C^e+c\5VFS,;98&[Q
>f9Y<>b>=ebUAX#4>EaRVN\4;-,IQ)](Z^C2=_YdN4#O4X7:aOY@:]7DdReP;ZJE
5)DZ4Yc(_.Wb[C&d6:96bZb#>TDG+<ZdT1KVWL4f6S<DGf<F(MaQ2QSIN^V06f9X
S/7<3J>Za8_\1d8WK>88-Y(K[=PR>f#-&+JSJGa/0WVBaF[-N=a+cSeLU8C-KP5=
>U4eDV-.2=PaJ,\;RA][-\8[)daeHDI9?P9(A72Dg&,X:\e>D/NH-AF(GN=PC-.J
QO[+-L+1&fKXU)2#?M^NAJ^MBK7b[/d)SWT\8E>DYHQ0:&5GA1bFE2H;dU_c77Fc
ggM\MeS<0=>@-&0Gb.=,eLa/-a/LHY)c2)\?]7\SNR8cW]&ee,.4AZL7/-;cH.D2
@b<DF^>ATE>/gS/F]\EU)Y9L#1]]X/2A88U=d<BNV,B?MFBc[3#fHHD#JG)J4Z&Z
(b\?dM:804)&YK,+2=(W3\Zea:0@JB2^U3gOH+VU5-\R0HZ:IX37_S0?C:=LS7D[
0XY7IL1PV[5fLURZ0BL3HF:(?1WGU/]E#g]>Q+4@T8LebD72SM,_[^TDF\6/@8JZ
L]9aI/Da(HPZ^Z0Ke-SG-_>>=1PP66DNaLA_>C/eGf08IdUY8:eOX]R]=ISeO@5^
L;&c[XfbV6L2aT?QKf\NbJY0^6_\d(R?@;7@]F[Kda/@ADa6)5QfL0CWQF.e4ZB.
XV=FGFC.=fBcQ3H<.E=IUDaP]IbF\1fV=05b/AK;[[)@e4\:>EFM#YJXQN7=K2T-
:1()_UNaFBA]aX(;3dYUGR,G\\F9I>A@=eXGe<,<X\>A6a@+XC@B3/\626IJN1fb
a5BR\=ESH,0>WO]4f^:8:a,KXMR;g-PK<PXaHRLDe<;1S<,SECRa-LUA,9Id1=XI
b/=X>\GH+#Y9&A[T7-[^7N,;1>M;8Q]eg4K5+2>f/J.Ib_K2T,H]@_\[,QG]Hc;,
aW7.XS-GR??UF1g9]3D;AS8Zc,:&/W[H:GR;#(aNOc+7TTf4JOf&fZ+_@?)6#Z0O
b1IZ-1J<e;#6CZA1=B)R^LEAbXW_eKCGNY0]7.;@C/\(;I8SB&KP7=,/UO>dc[LJ
G(J>_U4H+##RIQG,1X-QfST[EJ1D&R^7C02eNE9&YP3]Z(\\WPO#>LX+eD]RM,aa
dXZ^A?,7..;>;L](Q2/36]\CS.FB1@&5VeRMM>1C7dN/D=Q2(VO)(ga@0A8LH>.H
A_T1WWZE9eC=S6?@E.]Qb<KSZ\a\(8;;J4Y(]+[Z6QS4HF6L)Z;3/J&)H_OGW7D;
b6.bEFJFRZ9[,HH8dZ[T>QGIEb-9eL05M90;)6Y:66BK<O[f8YN#G&^BAcN\6BO@
IV.)1=ED+SO:>BGBUaIG;M;N:5+U1L7b]fRWX>+T[GEH]RW+GL8,K5TAeM]b6dF]
AS.&DQObLaTK.a\K<HHgO/51=c7_WQ@W=:A(7][JZA5J99Z<ZLB>RgDQQN_)e3Q&
=[+Eg0P1e(B?.E-73WTL,OLQ<)c-IRcQ)NC0Y3XZKa,a52Gdf#N]a3J/0EfcV8b(
T@HF6&EDS[dfUVSHPSN)=+6S#c?4G:3+\e8BF5>9]W>H@D>#-;.9(@X<a,</65A<
#DB4PE^G_B79KC6AE)K/[QMb(4N9SQ^(V\=)-U5-_J3TFIf4XEfSBP>2AWN[^=9V
:VA^5&b?-LUG=H88/d<MEAA4I=a>JMYQ&Hd.\>YNHdbZ)VVP.T^QQfBb6fJ/E@4U
=GCHa_)N<bFe=>I9E>8;4eK?=1J@R-1QI1ERa:2X&3UR-6+e7J[90aI,\-Ud0J4X
UIW:8@@c1ZNK2dP7[4eJHY2ZP_L2O660L/^7X)C;7L5.1:JAA)bPJ9D<;S=L2#@H
N9<6_Qa4T>ZcG7?B,>C.JC?J6A=,EMcU@UJ4@ITP=#e/.-_,Xg.)S[PGag46.6YF
F[eB)SO4+G=K,Oaf0bgU_Jb7JYJR-+&)cFM@XDGU1)VQJ)2]8L4a>d1O0f5R/@(.
Ue_[G5^K]_FE#eA^.+c5Y05Y(C:EBN_-)])G(3;=7.+#N^I..+>)J;Fc]Ra.9=L:
@C9:LJ8>a-AQX6B+4?eN5[bWZ&Ub?S3a=bRbK)2Kc>2W-91EP5bD[3I+4IUCX:D3
FI6g^Wd(4dCR_D5\P@K&de=PO]:=Q3MdT[8Q3.a@>]CQH4gD3RX5]CgIfIK)SZBG
GU6OCHU(_>??f7Fc9bUK0M)X-VK[a\45S^4?cVDTQ47R:4GNS@1ACHMe(X^Z\?N-
O=?MU@JT62YUIXR5g]^_ZGL#9=>d/)afIcgUPG7;:_gQ&Z\XKW8+ARdT\6H]U<<Q
_\M;Gf2D/^9d;>90Z1H;c).QY6P6Kc_4X8BQUL8Y)e)bVBGI-&S_LR:.W@,H>@c4
&MI^Kg#O-]]<T=eS2;RDgMHE#DNOL>.CR^(=_BO3QL)_;c<;0>VJ+=Y2Z)Z2O&9b
@/_B=,S:+@>J:N4LGU/K(H-0.,F4.;.G_P_NA(,_?N:GRLS2G;G+\e0J;?Ud\Z84
3Qg]35^)+cfa@KIa([?,C9bd=;bN/-a><T7F:[PBb9-YQ[GeBD0bbLH)/^2P=Z&X
Og?4D5Q(JI2gHd>a6_c7N;aGDDU=,QeY3-KN[(WdL0)EOI&[Ud(Cc+=[Me@^2^N>
dbJb(-/c?2=3N^CgQ-XW[AbKJ+f9\Y_R_6@:^XJO&f(>\&g(-Z#_NW&YA6Q6R-V6
16^>KUKV;W:38,cZ1HET/U>5S0Ke.11\]K0T\(_#=&?6:UeSa9)24R=(4HW?.R3J
AEa2eD/15B\SRYPX]0US?>^W>cAK[dN(@?74+I:5Xa;Ye^g70T]N9SX#^COd_8PN
2?_0?^:e1KVTUF63fC9Y^O62@U&eTcUb8c,&)SOD..e]bg@?]YZ4-d&XX.QF;aP7
1LRL<KbON^CR/;.;\)2_PUE=eVAAXD;(MGO:b&P[3&SBK#SFVRaG[7//EHH;4-J3
A1aNF)^93AUOGD27a^ObFBcPc\?P-)fLC32)3fGD0=^+g11O(]A_XQ1M7T@6I]?=
&<TA=RVKdY7M>6/eg=3B5?G;\dbM2G5b:eZ<dMCY90-&M5U5UOf)P7d/GURg0Ob@
?0I1LC#.6307;-6gVU?)4SdX7>D&\2+PZ#HY@1fH74)R+1dZCSR-3_&)K<].452Q
&^W_eVFb?1&EVSGYM>OU9D\UfU>c?b?a[;4T9.^RgD+F._-3B;GM2M)Y&JXBGBgJ
<C62a4eBU2RB,JgF;7]XJ4V+9>,?6G0ZPH5\T]<17XW:-e;0E@W\SOO@?YKaOc?Y
NDQ+MK1=W,O;-XIC591-,&RT5\DXRS&WQL:;N7NB<]E;eAEFUgY)d)?R)6)89NVe
69#D5f;V1FdO[af<(387;1]=[;F<#-2-O1BH3U-8ZS^/IUY;Y-_]+T\Q)@L1g3C1
/3AfDf6Ab-/#_^.+MU_TGL-fGGAe<:Y&[T+4N?M451Db5/:5(?,.M?P/A5CfB@//
U+7?38e\a;+BWR&S2dGE3HU&e?MMRY&K<=O5QRGX(WSHE8UFXOADI.;:[V?eaG@H
<@,ZU;D6[D=<OY_?+G57L#B)^DLY6N9-ZUaA6eAbbB8_N8=Z.3KSM_W(@&EZ5;>R
(4(,DM3SZ^;QOaJL#HVY1Ngcg4\6+;S(+H9[T&#7-@8VEJeab=[DJ^W8QM[QNH+-
N1Va?/Y;:eA.GE4#N/BNV[7#?;-EA)0I(4.R3(Y+ZEHIa(2GAQQ[61P:Fdac<+MD
30eETFD:\G-OT4e6G[>77BN+NUQDWeTQC4@,?<TQOMS?,T\SS458(?U7BfAaS09A
KVgVVA^1a>>74aW;Zb[F[B,+TOb_6bWb&W7^G\e#\N877S?GaR3IP/Z:8T_\QO4:
ASD>>K=C[#UgRXP_QP/-6b7HW63/A:/SV[FHTD<?:,(7]VRa(M3X6<>H3NYK6de,
,<7TE<:-CZHH(+Ed.U5AS?>ME7cE6096]GY4+HWE;F1aF5fA.SUH_IZ@+<N(bQ5I
1b7T#_92D-ZFSU.[FA&;1g7Ea.D=4@W7NdG99g1\,#9Q@^]:_3e=W/\Z6LZOeFD-
+<=4JGM5b#-bF.3[JZ7RcH7OLeLB+c-3fBC=(cLJTZD.,ga+#E/;5Y4;V)N,+c[E
]8^NJHL0=_FKPU)CbOL,U-6W1/]WG6f_EP[6LJ_>RQ00]L?3513,\Z#KM4/:[WJc
&210/W3W#Y+Ka:+2&;+d:]JOD@-f.IDUO4+O;.9\@?DCS5N_MdcXDKBK?dgELQ]<
QEbc2a4Lg]#(RRXTR2TK4\;Y68_(gFM.dAX;/5EM1\]Ub#,e>Ec4ObM2J\,<-32:
-NVU3Ve8Kd>C>_H6[0g/NMK&DD+].L(I2)2aH;bQ9I#&FV+8)GKRVKJYcDQODVJ9
7SRUZEOBCB5BFR?U+_Xcg9I9.KL^;3,)72D&G1=;4R\;\bTQFA^/ZEWFCcX?J;cO
4@>RMagDB05WE5fC#F4=[b4cRII##X;a3KUYb,FHJ/=UN:dW3gOY:8-13g&&TcI^
CR4XV;e7,dT\?2)5Oe@2>)Q[54]9^;X;5Tc&4S9S2TG/f-NOXEWCL^6IgX[&bJfW
=53#X&+b7_+.Y,eZa=+)+R?,<Rg&-^HT3VBVKEG1?-E^bHO#6O[(/]?]G[>3)HaU
#MfD\/94dO\^RN?IDB+MY09aaPM]<J0[,-/WAK:=0,P3b]:BON_[\/(e4.F/Z2;#
.Z7SL+\[Fg@d=bCTN])Ub4?UD.Z6+?e7bYg<,]aU0)7bPX6;I&5eDA\4OAc?ZQYM
X_CHD,>C=,bfd_HGGdb&=>-M1&=S3fU2)BZI11Y-CO2dbT84I)ZTUCFI[DSASX)4
CJ]L<Y?;@0RPHMcab[eH520Jc&6:SBbD@cdUJXY?T_#&M<^18=_PZOUf<USFW-bE
C4G9Qfgcg2V</Y8=CVQC40CH=cagf5=Y<b]J.W=J+/PCK(R.He336Sf@Df7H&+eW
W(D<^QYN:IaQ0<B(&?+7KP8?))U?5=9CZXG],>W9=6XgL6e-W@[M;M70d>_g0\U-
YSD6XE<Gc;;a/U19@NX(U;?OfY8W;9\-+<Y0V,I,PU1U<<VKVGRcC-X/+6;-P[JD
^C6/g3_VW9@&/f+-90eBL/N:V^RQWL8D.[KH7-\-&>GACNT8S80?AcZ#H_R4XGQ+
1F:=GX/O+Q=Q)P9Q9/O.fM\0,-)OYU+J3@eYAM?VAOgKDH<WK,H)O1g)FWT=Pe0[
Q1=B-S;8;Mg0\+-b0Y.aeW&H>DPgO(aV=E5e[&Z92ZM/0]ggeeWC/:D6U9aX-FW(
NB_4L[<@;0Z.JF?,[95+<K24]8MK4Rf^_PZA0TEb724V()S_cRDEad(:e<A&J]Ib
2:7a0d3.Qb/=]+Q8L#dQO8Ybe&g[0ZZ:;N,a:C,#G6SSGLe#.7Y2a6_]QebeGARb
\YS)+A,V4f,K)-3bT[,PT@5B)GG2F>LFb_4LP(8SKUR2>O<17L0_LTGZ#8&/&S6[
e5/)&;&\1CGCgLK7#]AU0Q-FPHNA7=NQ1/f]C86)gC_c>O5>5c)=WXGF8aJf2fT9
K\RDGa@:AcG3\HbM0aD[9C9SdX&#a[&XH#QZE9W?X;1U55V;GQZ?>?F>U]ZYZD;H
dcdL82Ob-X3HF#\OHB(fE[^aM>?E^C=XIY;AN@I;KXUYNLd-/V#\WI5)/f?fF-T_
>=<6/I:g>H/)[.Ue(F1Se?e>:F[HJ_@T[&JZFXKU;4.Y;HKg,G\T:<.Cc1RE4Hd;
G&;C:W7Mgg15C77.Md+76_bdMT&8F6cH+)UZbU5Y^INO-CZ#N_/M@SACN6BL0+K^
GaSJ7D^<;1e8(0,^UP3&4-BZ&fO:+bTQOLK6^?Vf-fG>[2@dE5AJ,(2@Veae/1XO
3A1RQNIJLPF9;2_<F.O+&EU+9G+N&&9e=_:IMOZ=e3==P>J#IfBI7QPKT3VNOdO=
N.Z@3P7MfL[+A3TZ/_.TOX=bSO+9:I,<T1/IR&2NE@N^04^R]b+9-6c6>N^<LE<:
W&R:(1V1]VQN:]M0T=06O/]>e&bJOVb<,+3PgXed@Y9[#6Tb0TY>RY<5BRWJZ?<W
ATBD8.EXW1+eWS,A8D,)3=SQfVQ;@)^?8]8-^NUS1QIVdBZFe^EWda>VG</b97;X
NHG-B>++2IB?^8GO)HA[&[W]Q9(HOW#+K2eD\U-,.c7KE6a:#EE0I-S_77A8:?QN
BYNB6:[(QE#+G;[?PcY#UfLHfX.E5bUI.3f-(-13H-af00@U<NQTGGb.O8E,UA@G
c_W;LO+N#Eb(NXHDO032eP1;&c:T?5^be]Ed<?\&THI(LYP8D>C-->=cK>d5/NWG
3(GOO&5LcCGOS>92__O5:JgZ/]V._(-,Q36FDFI)7d9C_QQQ3M?8BFO:T9:0Wd7b
He;8JB:)-FP0SZ?0(ObU^_gO0FXUMR(OCZ7DH+\c1:S>b\RCXVW+:W-#=a<OYgL)
<@]JUe\G8#YY9)J=EZPNa=>PUd.BfF)BT,XGg_V5L]^G7GKUE)g+J9W9U_,EMH=S
XG=C0?BI/f.<.=@C.>Ob:@5c97_OG/]9=#.U@I_a8,CC.e&R6R6gI&<B[_#6Z\dX
fEV;NT^KeE(6.fDQ.-C4FR)d#]RXMMXU.d2[S[[RcDHU(@=]f.WJQDO&#/4:,]=5
1Y;;7/8Y&c)JH>4WWEe]-&C:@)6cB7a=_S_#2XLP:GH:[6C-QAV)a][[_]c<_b,G
/IA.Qf20_V<05R=W84QQ:U?CLe(_M?EM)-EAE7-UG(@;.:-#eHLg8S0I4JWKK2e-
NIH+3B,Tbe6d(OdZW4g&V-2-7@WQ2U?K\5eVGe>IT=W5:EK>b@<7^6POD;PR6YNA
,WF;@XU3XR8f?)8,L,FS48E?<@:T4TN>J+VMX@4eO7R0FMI/C;@:TI.V8DF3eNPJ
-=#/6]9P^?FE[KOF9&ec23XK:4PO>=(&A4U6&_9A\7_=UV<1ZE=3&[P=7+8@X1S7
e(5RO].VS47:-dcL#-O-P;\[)bB[B3S;EK:KEY7;[?;3_)[B<,g7,b3@>8E?9#9J
<2ATXDTH4Wdf:[G_YcQbJ>SS3+TeAK;81gD]]QB[g;)7EQM^bCOf;BaIbKE-8X(\
eX6<VYU,5,eYT2#-JbZd^ZeC0J^)?2@=&:7PS/aF---Xa<KJ3L58#JY-F\3ALK^-
BVFfUZ4@ed0e22WZZc(GY/6I&1Cc4X?>aBCCI/#-[T&;X#8<.?2@fVf(L=F>&)6a
_V7X.L@g#[3-OMgKF4,>S[SG:a7=O_CeJGe9T]TVG^;cTgW]YRB]M=PA23.L2_>J
[^36QLY__VM,U,BeQUE+#[HI:,QP]UWIV29G-0Q0@7Sb&18^QER@;0\3WV45\88Q
CfFGQ[A(P/?;6cX;AOJ)<c41\NFVA1ELVaOJV]\+;^74?/JfHK@>8Z6:FV9b0K9W
G6VOg7d9bDAK8]&NYc)KF6OXO0e\VKH@(M01L6(8d3+E,=^Ic-6C2L829dWB&\8e
AaCLg9SSg_QXC^^La44];be<=T:B@^&Q@JR+A_G1OP2MgBa8R\(G>A+P8(2H3G?2
]DW<T(@X4U_,[Nc2DOY\FB1USceN@:X8,/D+,VLRVg.RRc.K9.,&/8dV&92)&bTP
F]B_EYc8f[0NaF^\FdMG=LIAN(E9^<e9Of?4RJ-+U,4aTKc4D?+W#W7JU.</f&Sf
g@UNQ>IF<5J>NBSSGF1&5V.IO7+)ZDFI?G#8T6ICM9[,#PUF?N5&22R@;a<CCB]M
a.^(3b/=>WR+QN.#IFE?;<PVD3LPb)><-V1;db->48R>P_S\_]R1<KGO[WdD^3Jf
S]J.1J>Ed:PIfZIH6<A.3_P@4#V1(R)dU06(+=PJcHQHEZGWC;Vc0NTY7])/YS<G
#WIg;QDA&\ac:cP5Pe?6)Z20;I8N@Z+[A2&EMf<4//EW&UD^QF):&>3AOGQ:b2O9
B5(c0BM91/^:I_<BN6[CR,-eOf.?,-MLNQgcaXD+2Fa\U6.6-X8NC_cLW<>=e;S8
UMQfIQc<[W#d^,CcUK8g)G;<1&>IF&,&g?_/bD_gTKDB_ReLfVFNO3.-;egWC\?U
e:d9QSR.Z59W10I]]\(6OAF7_5(UR4_HEF[X+S2D\KO?a-HIEI85A&D/bV>Kd1B]
75gRD4^_ZB+<S;Fa(>15DH@P-?^==g6>EB7[.f.]+6IfADGKJd.T0BO8^JP#L\-A
dE2M@BF>?6C(d>CUITa+Fb3X[/(?8^N:MW+\JUfVV@\.TUNT9=2)2M-+&9eV),?6
Gg>ICGY2JcXL/9\dP][2)4@8;HgS#X?ZS+E<7N;F>XBU>gU=gLK]]\16_Ld\NN3a
+?BSLR\Ob[Y&F2Q8e7We@c-_fSP+&L-+1(+]\f5R@I58bZceNG2@_UE+MY2&-Z@2
g>SZP3cNd=cVdUKJT1CfOT-f[H+aY1f-6]#5B[fH_(HHZ34-ZI>4,T9+#^XcK91?
M10)_]FDT;QO]BbU>G+WW4^W0FIVS=#+Z:-9]ODCa-0U(2L7U_@b=d[a=E+PL6-?
28.8gdZN_Y:AGRR-WC(.Z+[9T#,f[H0.+bf[_RUaID&4/?/U7Bb1?c+=7Q,].NYZ
5Ad.DgG:Y,<;WGR==5E+6O:S3NgJN:JX=(7Kc3L=-PTU13TX#UIJB.><>D9>d/b6
7#36eOH:9#1ed-^58AL\^JP?72?G6F5O8)#::ac_.>Ceb1:9?XV\8@A-,=[:-Uf6
&c:0:Ceb\gPH6BU167ZR;d,TI&U1N5;A&S,C87<<R.DF>gMB4:]2HN5GGfQ;6^;(
M?P5\O@24<_-8T:ga5JT/AfY.V@1KPb2=GNAE1cYK0a2KLDECQSWG(],>cg4)2+T
N/MM=51[G/F1d4E_B8BLd2/3>0AFB../?,E<AYeR9&<\dbgW2_I9\6NZ(0e^C^??
+TK>M&da2)@:<15^O;c[EW&^ZSd#>=60MFW:fY&MdVe_bcGXA9,9D=fOg4021/:U
S;+2A+Z.<+d#LYW0McK/[X\)-&@MI^a[0fX/Q=BXVA47KgBRcQ;T^UDB5#E.^#bN
A<BN\;0GE_=Y=Xgd@RYXPHV7J./ZDUa0?Bg<Pe#:URdY(M.>&;G6BfMZF<\gU;g[
#S#OF@Ne)&0S3bQL?GYe8ZR\>KA)KN[,:&2R[R&6_(PN]1:+VXG:@EJS93f4YcL^
Y(+IT]Z(L\DRQ4eA0V5)OWg;[UXBa5_fb1J_::;Q;&=&GWQ<R=@LDKfAf>OK)3-K
JV))E.1J#=QNbbFU8fT<:/fQ&VJ0]8?]9->(NJf+[HL87cJ9UPgLe:XG8LbS<Q-c
^9XA&NVbfC^G]>-PPJ@]RYXF#7(\[ed/F5.ED@5GY8N\YJ,CZ:=f8d:\#:Ug7WC#
c_cIJCfQU8Yb+/gJ86;\]./6F)I-U@GVY-FDa./f)SMP8/YW&eGEASbVN.W.\C;=
],aY8VaAQ&<U&Pc\eP?gF65]L2WEaW4_TD=f-2eS<1.9V4(/4D.OXDc,fe6)M[aa
aBPO9K1bVN<EF@_.Z<Ndg/.BAI&?b_#/PIXK,D0/6<BI1L&5&eIM/-NQZOBgA(c#
_ZA<Uc^eb>:1/DJV?UM\]=XUOVC:=NHb>XfVD[E89/N_]U/OL<<K5eY3M.=?ZQHO
.bDM:=XO?>9f];LS?3)V\Ua^Ad386=6RP.&PDB1>)WWddWQfFBR+=#Tf[<aZ>6#5
D<#]Md[8e0XA&,a,a.\g>-(Ig74TE7KU4O#-4P>:c)Ng7E=9V)?a:?E5e^>KKM:O
JRWKIMA-ZOaC/_@JX)KKNB72.NMCFHO6Wd_[H)cM?,TH#X4/-A3(UDg0>#(,1,5)
A6GF?e/f/[3:I5VA40W@S[f3_T0LMgD(XS4B?;T#TZgMEP9J=D5:SY1Y[Wc0X(Og
>A7?@JfYWLHE9b6T.Pg_;]H<BL6dXTP/(0WaVKS;HUCH32)<@SG]MeAHEC[c&LQQ
EV2T]F[I-Eb/TH,9Q7GYH^UR^AHS0g=8BeK7d<5B=#<d_P[b08;VOE&+-2:Q34GO
1bM^0]+&)+4[LHQSO1KO[LICG+<KWIQ3T2;4N(6S[FKU?(+]@+-f+]g]cHC<=_UL
NeXG<LASGLK,[8cB_ZBW[aE^XRR7BNUZBX+<011SeD=-6V@(0865VV4_N.+/2R6?
44LZ1K9?.5aRFYe?.GTXbDc,VZ8H/:N93KKJ:8gK]7_g/58Lb4GO>/J()eKF^e?=
A@D\O2]0L+ZV9?)]N/5-M7N^BG:O48H\^-\IbbA6PbE(WNIIeL5J2XH4^WVCXRX)
YKfX6R]))5HJ4O7;?/.M=LRLgL-@ICHW[>Bb9Z)_,E3]L.=RD];1F82Tc:6OKL0Z
<QJ,4PWE2SI&[TN7B56)8Odd<^S:;>b-cZJ&e<+NUeK6g<8&gA&c&9@D<5ZT90B,
@Y18TbLU@>#e#0>g-5^Z(EABAgfOTTNLbG4@dgcM+,U=D<>+8OeD;QXP.Pe[eK]1
_],Y>FZ1Oc_@MNTM;_[CE4W,LSPT(8YV8OO@E5]9gc2d9WI/dfCR0Tce^M;_F775
QeZDT@>>cTB&5+KWRdX#[&=L&?Va?DQB4d;5<F&>JQ,BF7gP2^KFcdFb)gYJVXQa
WA:gKd;/,=IAUAI@//N&EbB&[VTDZ)DQVRI@(/8,d_5&9dOI1?FDKE#M-.N-::C_
YJ>?5CGHVQB/S,DV=PdY=@GHA/I>;F,4&Vg-#1TJ0VeSRG\@f81,HdV?6/;&a=X^
UPUB9YY@aMOWLcI)]#cIa(P)bE_7cL8X[XJ<G:TA+@N(b7_g@MT:4U;Be=.cA[Ye
U(L]C1X22X3fCe+C0597IZ-HDF#bNIEH?3>71Q1MS458R[f;\Id@g4:DW4g^34JE
_?fK]?RP?88J@_LL_4E+/D\7(+K><<(^9:T5SDOYW>L)>QfH6^WJ-73/IE_UD\P0
(2J&#MdKE1.&M[H?08+LLY/c,]Ld-CAK#<gfO-)8E7T)<-C8#MNZbS:dDf-[.K:Q
(X12Q,)P_@0<a(/7(TK.b=[8T&g;+.;0MV4NQ>BEET#_)T?81+IMG66FL.-WA^)T
fQ,1:;b)VL_X/<Y_dNF2R7[@6MG6X42ZAD;eUaQgd#NM5.7E^&ZX4WOFA,YKW=d(
O@(FKg^HB5I9Q=DHD9@4O:]6d989Y,V><f>;),.2@c3b.I2_6P8gBY^(8Y-,QGDg
-P9ZC[CCeXML=)Q)1Lb-c(@WZXH:f(ET&-B.GH#PXBI,?bHZDY77&[YT?B:Ca8EP
&VaO8KG)d2HMa&[RQ?_OLcb;+1f->7#bDA/Z3]JHI>dNX7b6>MedH@4>Y5[b@e8N
TGKR3Q3;1ScD/AJA4PZ>;XNL^(>\7DbD(2]#\5a;8TC&VQX?Y-bNH(@([=EdGUYK
<)]02QK\(S84?AV1dRLC<gM7)NTaP5#Hea.X2gR&L1F&KEC35U[^XPEGT,f-U+ga
2gG/3F+Q>=0=C8T6Uf?ZD+3fJ7]VO5,A;Q)H5+7c]gNbPN<[eg@4TB?FR^0H3(Z:
<,R][_I8cF/^4?1)ZH?#9>=QQ1-_/3KS<H_105P?fFJUY>gE#ZR]==7>92a-Pb7>
Te;PLb&\_P?WTeEBFO;6>/#Z^S+Ta/3C2M5VXdA]+->T_S+95f[.ddIQL@4@A-J=
D7C^<&<VbL@4.@0L8G<VFf[H(-26WZK@S+3EU0DAF0CV?08DE@M>AS.S,C2&eKA4
JNI\8Uc3Qa\18AB-ZYb-Y2U/fSX;.:SdT9:GRW</YfGME#D)./&DQeA/SJG)bP@<
RGYYcgQ.TGN]WR.&]W82b[d9_&S??+E)LA&Sdg7AB\YgF.79cP)8PQ,>GRX4dG.@
I:+9cYX[V/N#0f(;FI.U?)L,PgR).dIWVf2_SGB4+8L0Q^4YgQFSgVWQT7Q/:?8Z
,9LV(^H=OI3-a[I=H(acU(YR;.AB?3E=V:F-cgO(dL3gGP=L1@N.K&RZ(<&;fc2a
^Y99J(e)K(<N0J:P&19NLCb0,)=A3#6#M0=K(\.f2IT@PP,/gYcB;2/TI<[OLU9)
e3E#[&Z7O#77IMW^E6H-&W?eXT7[0ZA&^RL7F)E>>ZVTE&eGYW@BMNBCMWUU+a0(
OF/O=d8S9M3:#89YCT/(S6fDaBVM0,,BYV_HT]NB4V^?41JKDWXN3.]Q@=8d?/a^
+#=GO-(c3^BUMSF55=(12=T)7XTO@PVWJ8+CGMTF1AFSYX\Of&?Cd>LfZY14@P:?
EIY32OR3IW1c#5]eA9EQA7=C&Vf&XNf6=.?AID1(8X]YDTe1M(G/J;XaaNIA?F#/
gSZ5-9e8I#,Zf/W)6HIBFS]^GJLFc(_M]0-QWT#)[WfQ\WJI/B/,;>f;d0:&4@/<
TWGW59D63FRa#DfCKb/#=&IAcJC?Yf_7[VG=bD^&ZHV[G2T9X>B)F46gB435=G^7
SE@9d2aQSWJW^c-H:4&^6K/L6IWOD3WK7cC\CMOD=V6]SX8BTQ:LWWf-Y&TGP2S:
e48Mf&:5/;&HRQ+N9.8NdG\a=A953eIKGf=)WL78IY:/8b(8N66R.=e?V?.QV\3c
JDBg_)X#K0J1O61,QV.Y/S;@4@9fQS]VDG?,^:bfYY-aYAFK;aW=4H()EDJS]5+S
S?2VZ(OaJL5NG>cG3J6G7eb.)FN;#9X]g_5NE^A4aafV58=I+MJIfR_aH[0g1:Y]
c=92;Z.F84bW;Od0[KDXgZGa.H[g2H=dOM<ada#X@TCK=edW)2_.,_XC0D=g8dE[
1^F-ae)N1<5II6[QWZR+K,R<g?59PZOB&3UbE2(O.EV4:aEc5BC<a<)TAS7A<b?^
^];Zd+Fg,7U>^[FS9Y6\cT_:Gdgc13UdD:MTT339_R-[ND4:8<4WY<-aGPd0f\77
#gI+5F=G&;(U_Y>Z(NUB^T6(A&b3MaM1.I/e20V1L;8U=/>X<E3D1BeWG/;aeUDO
WNG<7cE_aLC=STL47]CQW#-Q)2WcaP)R0V3;7(EX<@ORK=A5:,G&_HbXX:6:&M-b
cZ>FFUA>]M/XY=^V>]7dR=MZ9L9/Xd6&^]VH2AF@RNZ79NXYQ\O7a:a<Z0:ARX>&
;3VFWMF:?-?AUQ+AeET;H06S/PY33&V<b(>8dQY:4NfLOZ6M@-;a]QB\&M]gTG6)
K8I:U&:2_4L;b0f\?bbQX]#13ARLg(H2d_.3Z-,V,VO-,2+)V@Q.:.eP.>0<1)D@
9E6\V?XNA0(0#(JZH#>C\@EBBL4?C:ATWe/G=;Afce_gB8#WX&F.MID1g1>_[4]1
9&8<cGLZ/g9Y5-<fM9>_/O./4V\ZFKRI(623^><OVL<&4?#3RJ<OecC]5^P2YcS9
>:/SUYe<a7)]F3/R#KFNP=^Y2VHN=L-1^?COc>:O0)\QfT0E)^6bLAVEQ>QOTIT4
EcddMg(47,^B/QX@9]NE73&G1DcQHD7_5)Yb<OBe[UK-B>&8aI7-J7d+>T9J.[1/
RT=#&f6&YFB\fg\,MGg&ZRYXg163Y)U7Z@FHd>IV3(7[/779\<>OW])SRBHg/=Hc
P6L#8<TZ3=fEK_d><=/Re9N\0V4A,GRf>UfCV9d8cMZAM>NIYQAgBb@Yc.Z>7daa
A7&@d^?1BdW+]gRY2MEZY;(/<_9_MQ)2;>Gb@M2=?RQ\^3Uc8OGMY3FY94I4KH6b
8-LNB61@UD78>4H&+&IH?gC,B15fG,2EOE9&Q27b5ECTL+\gb@:a8+PXKHLce=OL
^24cCE_a6<cAIT>GWQg0/?c(/P3PG=/QB_TdM&gCLMBg_bR&257aF^BbQ6\,)9I0
Ug@N3aMS+eOY@eCB:\;4dZ\5&C@9ZddETQ7&<GK(P3ASa@M+F-Mb3Z=X1G6bW0Xb
ZI9S364=,=c:6,TJH.aVYE##?-f,Q2-f6:TS6@C.C5S7QH[)0>EV1M+N6NSF\8Q>
G<c)XWLOA/YWW7f6R^MbGR1\)ZF3-ZG=P7&^\E1AHE.>(C9?Y5+P0df>5=Hd/4[T
9O:J8O<XP?K&->-c&RRTR5_HbJ=9C:P4B@8D;)F[P:Q\\H(8b>Ff2=?2TO1[f<Z=
,@Q-7&(9LPZUC.#G51Rg?LB/\]9\X+HC4_FGZNXI8F;NC49H(QHXDZaUM#?ONC4T
?8_-=F;L/Y<a^RJ7_GQGAY--acOQSI28SLQX5VQ6FZY@HG_HY)/fe[9\QP:>,-Gc
a@gJGVLfARKc=^:DV/\2SCF>d8^L:]fFLGI^@UB50de,N?Q<9:a586PN?PE[EL:K
]7(5c5EUC./SD4:AXN-;fSPQ-9);;\c(dLQ2NM:\:I/_;ZH6AB1QBQ_Qc].#FFGN
c+;J4E2QJIM>DG(d\M5]>;:53^&e4GQ#,#,\QI>DBH,,PJIO>NI]NKU_I?Bg_/LS
e>XPP=J>I=+1U+,K0VO,7=/@7K(PKS02TC]#XN>_ced_\[?LbfSgc?<(9GcA?a?_
H#=]07.18.<7H#fR3&cd1-b4F>/,H9>L<AKJ\SgEd.D2a^g9V;c8SgTX0R^RNE)Y
?9Wf7eIBYd2?V3Z)(e0AV[CL.JE\-TI0@6DGTX37cQe24B]ZBaf4W@Wc]=>aGb0K
R6T;cfGJS8</C]O3@d(.Y7^-H\5C=?>1/VRR#\0QQH(=[)8\M:a]&8gAd,1:Q+/b
,.:]JVP)H8,\@H.##=XF;87cL\<,>/(d9F[b[BHMAWOcYG/JZ<UB9BKB.a\:KO;J
UbfGPF1JXYMSd3Dd&3/VJPgHD+B-cR-::7AU[_9+_dGLY7#[OXcg<):B1b@F-#)A
,gUY^cG&JT/NP,LXN79bSVceHcW#K8;/Y&E/5b1CTdV:S7;]P^\:]fQ=e6Qb[CMQ
5F1JIXcT3;bAc&J4HLC=_Va<0(PYa2_dRfTT5W(\N2TFE&7OZ7DXb2N^)MQ@8I0\
^K,g2AOS-@&;)gVK,?:YB#4K[F5,3H09GR15G);O7&C.3@e:TN?O:14.2>09+e\8
.QbbeTC>gI8EKE+^H/[Ma9Ae&W2T\7Hdd8#,PddcO,b]dbHXEL>6C@B\\1f26OGe
Y>7g?63e.NB&:(R7,g(44T,V[egH+b<?;DEeC#:FU-N_U=)6KI&JZ(g@e8=?QV24
=dMCG9+K7e[bL7_RM(#+L=EQ:=F4g0WK_RgLFN29PR4?:3-+(FIF5,&LV<R61d-M
N93-fXEdE-8F>#D8@[4GE+I2\eR7@e,/I>dP<NOLQC9gJM,?AFa4RW2=<&)^]8c&
AEEX+YS<(X-OaGe#-U3V;Z;cX]\ISYPZ)edF,cSN/b<d[9dB;5,-E?9Y4CJac-[C
IMS_<)(:M>?[g<8NGG33+DKS+f^17-bJD)(\NOC83@ee0TRM(X(83?U_=GEM7W(f
O1gReBFC?\2WgcB/JfB)Mb\CYF;&&De/BK3GNS](&]DY4cAMJ/6Q^;-GV)NFcc_J
ce9Z?,BP>Kd)PVWJ=:<5:7(L[E(A(ac.S=[OC[0f.<APfS)L9HX&^+dE\3PFE@0K
/^L&J_)=B]Hd)1,RXO\fZ-^4G=XCI@FBD[X,,KS_bY22Y#W3C&<c)3g06>KZ1VBY
2?RDgS(,4(Ya436=/V<I91?N@AI6M7(8ULX5FEAN:dKe_G:(V?3&:K/<<GB[_:^=
Vda-DAN9&[eRXHeF,2R[F)W8?Q7[/.YV2SSRCLdV_;#.^LKO8.CWR0P;F9N4&+IE
..TLfHRB)V#(RF0),\T>a^_;7B&M.0[1UY,1T46^Q?4[b6+DZ3^/GB0H89@)&1fT
&W_4)d4E.D<KQ8I7AW:NT)])C?E?^KA0#M.-3^TbP\)S-K7_TcG](FY=d(_A]+MD
5aG-Ng8?W(9SGB.J?#U:+7H?\Vg>?N/)NVE1]2CLA1gJ)eC<e7cA<=DE+>?08TSf
]^,A3T6Xe),fA:c/?GF5APYV3_O?>A?YC(3bPP68NYf,.1P_P(SJc834YXTW)EO&
J,>g3_5+C6O;(;4e-<=ML+c+W?f?4e)3&OCQ?MI0RZeD,aB@)T6UH(aL>>C21\(5
.GC(--=]7VL9.=4J&<cO=IC8^cM\dFM3V0b(?FOKTOND^<_cA4cFgCJV[eP(3I21
(f=#:?<=(;V+UC?]BW)10#5UD8CS2.S<?<0JM?K>d.]_F2gRGZ>Z1CcA1;e2gT3c
4Y44c:a=EM]bQJEC<2_eM,&^fG?;gN(R/NPUa;V1Z-,ScX^K>>Y#Y[6;,4Uf]Wdf
0fV9Mc.R]9JeD>>B&0c?I2_2)((?#3?_CT#R^fJNG:=]:)9[-Y:P5I&cI5e=\bZX
(5J(DbE.SOa8O-B-Q)L/VH-N97SIYN.0(B380dEa;<1MbdK>Y56-OZP@ZDXfSJ-Y
Ob^F>VBE5&]Q6PWG0We@:HBX.gNbaX,FT68CJ7aF:-J6<APUN8A_0C)/-f(FE082
LC5\57e_06ZF7\Jg6#bBRL(M24(/;BSEe1\cQf:OAK6d5/:S?AYYSOVfNg(:RJN=
,deWONO42TD-^:ML^Qb?AL##8MPF6G#(=Za;VR2VMG#DYHb>dg+&6cI-FZ,EW5?;
FTGc(#Vf\C)_)EUS+UJ>1NGLFH?[9fZ);MaJRJc7OS,CAgE8e+^N+d+=PdGAWGB3
^FS6;4H8C(55@cI^P+^?fDG3TS]#ASZ-O\BV4P[a:O,XggR^C--5dR7ZBA;,OU=L
R?:K0DfOfN6SX1c#d21Q=feaX=_HC3KXL@],AL8+U3EH)PY9GTYC\gK8T6QLUe6Y
8=C(d[5/F]_>C/Q4X9H2dHB2eO3Q?ZM:;XN\H>.P]Q)5a:TcgdKa5=BFWOb/G;DM
?e6cQX/NPg+<g1@Oe&G<Q?c&0c<]F=(020FZ2)M9^bQ[08\BfBcNdfPWFCBD.N/L
\C]D[]]IST0^dIXe0_G0BF=KW=O2^Y6QMEYS;L[K6E3^Q=2c>#V]fcYXVHIA5]/e
f[&(;BIZ,-YR)O6#P?@(Y]47+SO]R9RfQCef^UTP2Od#,.8KKa4FZ^+fI7PVE+-\
B:W3=EM9a4b9Z47)YCXPa,[cYD[I6)E0?YdPg>;/W)f4.]\,eb9;F,?06DffM50@
JUfFePS[8IM810aCf<?ZE;SNg]QcHbb<&KOEf8K)N6d#7Xd?,?fdBQaVXg0A&Y2?
F6R]b5)7;H@.c)U:#UYYI2dZdXSdCUW@+g_dM@CD_VWRgP^J1PDE]-ZgF0fc^^YV
e>RD97GT4\Q0_K.0@;=@;TM?CRg,FJ(@?QQ8(W.916M[b9BHGJLL#g2eE.2C<P]0
L5+\+#(N]S9D)Y5MS\?>gJ<+g.7TF6W(VeIK8GAbEH).@,5;H:IA6&)N4L-U;fFI
5<HWP1+MA6a<fHg31S2EY,U_b&?F-5)f3-M0bU=bcf/>SS_D8aDIL,QY\ZaNH5FT
V2<+WM[[O=B#e?0\^TB#;#_AB5+@YSAK(F3I(S]Y:D^Qc<b).=BHU<J:LK.CLbU6
Od0A#0.f+8S^03B>D-VCD[H_IRHL#W8Jg]0&AZRMd_#N_;f,SaFN0EG@29#IL,I6
b,aa>X\=O-^+bc@UB.Lc#gGYZ2P2a3X@J1,cEB+24]RR;7ZLRM_#93E[g.O4(@48
-g8ZLC8J:eQd9:H&@dD9bF/1)6)?eb?-A_WF6[5XS&;&5(aXgN?b((FgHB.E^W0#
Y2(>\IILX.Y-BALMad<eN_#C[J:M;2>bba=R-L01RPZf&:WU-7_M(M90[:<S/Yf?
8+^NaILK2?&P4bRIXBV(9SQ.a+5.8^VRe7>e-(+-;2/;#8Cdg,#YV+Ze[X&<6296
_/IV,EVG39ZUJ@Z[Y]0Q3KWV,==U?VH,2(WZ+[(N6f--gc+53FeW\D.SAYa[&A&T
?J7MG0VW6_2W)ULN?N&aOOe3+8VGL,K0dI_-8@>)F^[4;a2\G2B_VXLQ6&=..a=V
^KW9&ZYM\@T6,/4K=<f@PC)AYS0@g,X3Y?f4S15R?2T/g;_@dB,Y+eebF#=#\L6+
_YX[4RP(cd:b1:RbU+ZQ4RXMH\1)QRWTVHLS9.7AXMIRP36;V=(0/KA)0XGgVD7d
K7N<CW#8>JIC8-+ZU-OQ_A./]eCQX.g(P#,B9OW2ee#7FQ,Of=OF+OG7g:2Y.=dB
5g1<W(Je.8A58=d<N\&=b+&eE<TYBOFFN:6K0,K^S\G/14fF>C04QPRRaDP?>KXG
(C2LG7N7d5M88A=BUA7B0a70OIC4U\7G6#XdI]e1@T&F42NG5GG&S\\LdA+R^_Sd
aL2EBAgM7I-3RC2>g<U]HATB6b&L-P:@318dScYbI[5@R-W-aEY>=@#<Y.QJ[3^?
;Y0?:7aV1f_fSVdHeZN[KS,WX)>0@D\@b&/1^?M1#VaP)J+e#<:D6Q&992H5ce^8
^8R8O=aE7C>T4QX;.G>2B8JKR;S/MNRGD9.0&9/I[.RS?95c@15-4)@)[Pf0R=fW
WNEDSQ,HT?JP]fI(:(]AXR45?2D0dCWbDKSS&D/4-1aM\a5DD904BRU)(<X7(++1
VU:K@7UN7N84UM:ICce7(V4UVC5]V/^c/C66Gd63H<GL+LEK,_2YQGe1Gb.J)#KL
CS@FCTaNMSHD[3ef6<[M[N594R]A,\T3]K69Z<;<<W2UDg38.(.#)EZ[X2_^#0K7
L0:aB2+A95:.Q@D7RGSRN;<E)9>;c:]&2T<NOEId(bB;^e-a[MT4;D+I@+=(25e8
UDBRX>HPbg:;71=>QG?FJH08gA3RKP@<6cM[+97ZWK)D:#SSK?G[KZK+TDb(&32[
aRV0L3W/KGPQ+J;QY;ZSf+>NRI(P/aC<(CQ5ZVSF9f391YAUNY:-]NQ_/A&DR1H<
P;[H6T43eTY2-3A;]U8d^:9)&I.TM\UXI=9ObLZB>/2&(MeEG,,#^BJ_DCP0gO.W
+aD]MWBb6aYS?/Y:BD9Vc77H,00?^J&Y,_V^V51Z9V#/>43<JeU#)P\Q)B+G)Z?N
bG:Z#=1c6FQ<_-P08g==8V+WQS>U@RRHM<c++M@T029/H9(:--I?aIbW>Eg/WKZK
G+I=+b,g]0[EKYg&YDSIFD<8;9)/cf@5RVA]CC@0\YQRgW^]Nf61NFbHMKBM_8(K
cO12UTU;c9LP-Ee[MI<(+7<+#<,Q-Vc]O67E7Gcg[=a8@H>^P#<4^7-OPJb(K.GI
CFZT0W]ZLJX,J..gYgUT^0F1(3.#ab/g5R=-=O4S9_UL<XA7;fgF#(ZTW#4-c2H1
+fN]YN)dX@)[(8MS1FQ[.B68HTEEWNb<d&.W6--_@[NJ?1#R.#I7[3/1/FHKAL+W
,X4c=F9ZU-20,YV\..YUe1P,_U?]=XF7K7T4cQ.ZY->]LSJJe[=c.(g,\-&S64L<
9DFHK:Lb=:Ib#?6Q(>7WV#JaPTM<#e4M9W7EeF8)]a9R[OI9EfL<]?<,;UWK=8cH
:#Zd6Ic_VEU&SKB2^Pg4:e__B18J1MW<LT-fgG9Z:YZ&4>5C-(=[<+_RQDY:WOOE
76O/:(N0@5)<=a\(7614_V;95T652eZGP,cMC7=L;LEU&I)9afNLC)V=c+V@cc9]
JE>?<=;IQB271YWWD2gbCR1DB4:MFA>E+fGGY#Va(PW:PAeB[T@\^_@\gcB)X?P[
_g1/c\.WL/9CN9,FKHQ3\S7&J)9RcDPDZM,_(L<6]Ng9c_5UY_.7>GL:DHNX/R[N
HTc\#BYDcH\AQ9cRL,=_86+-_H>cY<S\PD1,FK^:E))-PS3gHD05)]-A+_,YRe)U
Z=LDDOR#VB:[C&_RNZ)O\:,6]/1K/P3K+QA/Z/6GAc8>KZ0CX@e9)8dA50.bY9_&
P,NcMQ7;[@fE47TE&82.H4S0KI29.H,>df_=OB7EW)+T.P/e)S^;17<K2X^]WOT[
@d([1V?7KZQO0M4RDb(&GI7_gec/O#?U#/I=2/T82f,[eAOG_>YN603?E5O>c],O
6L^3&ZZMT+YT@V-OL03eH2YB@9P?=+4;d-T^TYJ<XKQZ1QI)4B7MN1ZY8PRL-aA)
MSc+g6eWX65(@K)JP5O.Zd@CA;),DJ;VH1?3eC.QVf/F0UHB.^?02)3fe/XC;R\L
-:A=YW51P0T(1R;N,);aI?G:\Q8fM9ZLI,g+/c>4\HQVa-5H=B.6eT0\+.\SaU2C
G:M[;^/;cBHP^g+S.M:Z<J]gdUYI,S5d1Y)2:95W3PHc^@FO>[45Xge5LOS-83I(
WIA74a=^GMY0Pf_>)S^EXVU/cL?B8@f#4dL&;f\G1S6bA6=c)XP)f\R#9\FN(I)-
O[<NcZAW)HVO7U<L&UFGGC0caHdP75=/_Kb-;?VJMK-;gfM74eBIC(dAI\W8)PSW
\NXc4QXHV;T?<,b1fYJ4C7>YNL4TJ-IP&1;CIHNJa8?QQ#.QK)BI[6LWR:2e]>PY
+L4ZF-G_>/3RbWb5d4O>gV#fQ_9AZ0[@HJP?3O4,G#?+H4(>-M^X3N(NKONW053]
\+_:GD&TFJ9=U/.5L6fQN#Y@EX4ZVTQ?R2<f<.I+>d?TU98e@=@^ZVMN@.<CO,RI
6V]-J=[#c:<SJde00-.ZUDL[6UQa]GQ7IVXcWY4-UM;,NN<,TX7UcfS)c;cb8521
[XA4\Y7Kb:A>LcK\=#f9;0+.OZ@+e\NVSRIS50L0X\\8Bb_;_^>>=5b6ebZ]7#K@
O#^e<e;Y:.CBD8Mb+.TdC3V8OW1J<c74JQSVe7.Rca?&;3]<^<c]R+c9J.9RX^8B
+?)=OXLX-ALg]E+:e5CE=;+4Me:)Z7Z9bP]f&:UcQQD2@5<RUWFa(:cGSUU3A5I9
cZ,Ag,(PQcT09==6T-\9R7D/#C_J8EWe-]1=XFIYZ.#2^&\5^<\GbgDSE.SCf-ZQ
ZA#0H-dLVF,f47fecIHecdfD4@ALfO4V2MY(WgS[CgB]3gQOFC=MOcf4)c?-Uc7(
K?#DL+f:ERaQ&OfR1Z<TE7V78ZfT_X_bFR1I^<MOHF?=P6+F8N13BMV^NVN<,e6)
=;C#.I9<^8/2>ZZ]:bDH@g[9BVHJbBMB:=5aM6dX@H^8:SS_A0^8Z-(^D]>Z5Q[R
EO;_2]H0TLCC8R>JGEcGJIRS>egW-]Af[I?S^7\1//SU-2E-LIOD^K);4X:IXP2Y
;]Y/g0UX8e=a9a[/8EL(Q<@0<XW2UeM&<O_A0;E#P4@;(g1MHBcIM-T\f:/K#U?O
FL2J,A&V>:PD3a^UWR@=6G(2dP1K49(:Rc;8PJ80Q2I2:GU8MD7V5IUK.^++FSKY
eU8LW5?P>E0Q_C.OaWB<H=<=#GUdB>F;eM6K:XN4,99ZA9cGXB\0R3RNgc:NgDN_
R,+Q#9LQ62=Q0?R#OIS[1Bg^>KA]=/Q0fI/MWX-W::0;?MRXAbNB7_3RP;+7=K<Y
8Z9=#99R@J7.F3LX_0A5X3,#.83,N)M>EFD1/-04ORGeV<^46[>P\DRLFbK_,9Ef
5&NHI8QS/a7CFHH+FE(1)6-EI@QIMZga@>=PLfW2=W[R<G59&IFC-c1AM4Y,OTA9
2Z/fFgKK(SXY@.\cS3/]\,FL2f?N+WW(XE4=?A5:74;R4cP8cgB[-Nc+CbGX<-J.
VeM[,U[F9T)F#egbX=_#1)O6ERG?POUL:<##DH[4ZB@T+A=/YP49;X+cH62eJ8O]
.YYB#81)I]M6cPZ^#[.FX3NcQK263)Xd,_7/D;5Og:2YFZCGP2)S?GX6aYN6M4J<
5.b3/NZ0Y3436:7ORJ2>96N?-RT\9e3]BF256&7Q5MQ6S&KQgNOX_(LV@:P#5&Z6
Z/XOTC7-B_^d7,M3BF?\3TNbe6I).HI<P4a5b3BF)]B@J9L(62O<bE14LUPR^M9F
;TKfHeOO->;bSGG6CcF)W8WaQ]Z)=,@#R]]c[?=Z9DX^JVA5Y17;UHd^K=fcC0]^
1^[O?).f,13QD18fKRd?Ve=-AL3_1fH-?TMP/F8R2A@M4RJ;-;8&cQgdYU^MWJ&g
E9OABHLH,9+2L]/9?<dPa(OJb:\/ceUGD-FR(/g-(([Ae;a=IM2E#bTJIT443,BR
3.AcG)[5T1.IT2S^Z0TEeGa032.\O7<QF[:=2/e0IQ3\3dcUbAVa];3MaYB<f/+&
W5YF0M:/0;43<41<67(2<a6>Og&1Nd.L9-Z443,L_X0K=5JCAMYF42UP\b<>ZQ2(
GZV5\+A#bV-OZOWaJI,IEY4:2,])>N[WGc@Y@A]BY.Wf2_+-5ZP7B^D3MEN_38.J
fI)(fFb]R;:U/GL1&G4<7_dQ<c-(\P7R&O9D9M8d4Q3gaZY:cge_L/B5f0B]TWW1
3>^^WP@T-d9J1+(BEJ,)\YBHL:Yd)\0JPQ)&^[:MO.?,SGCS3:W7=0>Y,8)S:B;:
&&D4VXZTPD#XN1QH)8U;Y?<+eIT&fVgfcg6Qg8dW[#aUU1XLS+.WG+06&R^E#BAV
Q(\0Pf5J+,RU7F?HC/eO?5d48gU3.>3;@F2E<SY>QaT5+X^geT]=2\X)Oa+M:GL3
;4.gUS=8TROPALIIe_M_#18a_dUD0@_1KEV583B=0GHEV?5AG3JWES+f92)aa(]<
P)7)cQ[@C</6,-[@=4F7QNURfUg41I<[@f11=4,L6GZ#2U8K=9JH\YBB#b,2OL#O
)0V]AF4,?RFOU6Z6T-]&[e,IDaLcf8BHaJB,H[RDCd@-SCU(4\]Ve]bc/A=BT;]#
4R&7G]>)NJ_GU:(H:b_LT.T30+8<X,5-\:>Q7J[g<^EDJ>49M3a)MNc#EDAJ6\[K
e.YbbKB@580P)@13^,7PV>1S<P-MR;6:DA;VD#]:,/b\Pf<AS6@^],=W2F5_Je8;
?F0G@>g+JXM/,.ZUbV8YJ7#ebI5L_<#A.CK\4W\N[],&IK+bAVeDU+=Wc#GW)V89
MZ20,I^g=KA?,fDSR)#+N0e=TATF,=^MU:TI;fYBUL8^\LM_)W05D=S&E9B@-V,.
CLE.\TO_(WTBA&#eeRDPUIP4=79c\PA+g>-_A@W#U]1L6O37\;#Y@ZdB=8A5dF,9
KLG/E7)UWCI5]@9Gc;Z,29SH-5(cfF]-E#FR:+W2@3U:9f8+I<5:;-77fg8+04U_
WFR52]geg367=&e[3UN<?HH2^_<\(LV^MIUAVfV_9,;.LJ=B-DG(:YV_fb/5Y1;^
5O29cHIZcV#d9\f],:7&?46@TZ87#5_>ccf.MVXG)=9R@eO_J8fWD#X)S31\[Yc@
]2@>&-F/\W/[O0a.0V@JbdeQQQ;[EX8<3]#X(ZS1CTL=FEP(\(ZKb;0@:?aK?C6:
e,M(UN/4@cIIK9AgN\>aV3XL+7DbI2Q1_HC[aSc??P1/IMEa1;SFf;V<=)6JYL.[
506[-GC:R0?87bO+b](Kd0IK<Nc\dEBJ8)HL._SM)]]^JQ.6?=&O=G7?/H;Z44e0
S>/66[P#VC]+?a@PXUP[(eK/Oc+A<R\&#1Og]GAbMAZ_1GX&2.&B&B(XYGHM#BOH
FbF,YGKF=WYMSJ2O&[K)UEM\e^TYC=\TQ]SYRO^bVI?J_?)K-\HbW3KZc#:ee^Y=
1>WO;_V+a,^fAPS04RJfIMe<HD@IU9:U&)<;42Na>g8d/6CIX29IaVH?Zf[;5e99
UXGXE#HOOB@D6IE5_Qf)IBU;Wf_/#@]A:fI;:+-&.QPG[6IBd?=4<;TE4:?EOOSa
d;9>.bW\#3)P/<H-IMTZ8:BJb1YVNA4J[AW0aI4#T.,54cX,(L00gO@SRZ2U4X3=
B1Q+Fc<3HGXK/I-T5I-V?c;1QD]SJRYQ-@X(L\6DN(:2\U256)N^G^T9U18A.)Z3
F37/?IHME^a.GB/E)4Abf-+UXA=4,14MN5^=7FZT^>??]FCC/KN4P]0B]#a3G+;S
aOHM[4K4c#A:E\eWc(ARF8ML6(bM3&+X=E#-4C;#^3dUaEQIe(S]GRgbT&IL-2_S
BDMC^7;WTB.6e+-V]Y89)c\GXCA@;;RY^&.IA]=RGSMEX;b.):0K/f4:9&[T63Q?
2MPT9If?3FU:Q]PdIe?8=3#a@+:?2:FP>)8EOJIFW_b0PPZH890OEZ3XZb\QdNUf
./I+;<]^],+B36N6[Q#V-#N5YbCG6L+XW6(Z(dPXQFYRK\>a+U#?(CVb:52J);bM
TBgB@6]84/YfF,T:Z2V;L>b6-1=g8VUHfG6M//80S\]f6DN=RfFEAQB&U=H]S<9/
Ff]Pc-+eJQ\67X8Z.67;CGG8=bg/XT?C<XePH\HKDO\[^&58#TM8?T<)+1XV[)E3
KESAK#YbUSK];<WKCd&0(gNUI_[2C:Q>P^\O12I9+_3PN\NVF<)IVcVb&^=A#_QV
gLB6?KN&7U)(>Y2&N/@33g#?^5J\-^GLY#+2KbBNc#bL+[L2+@dY(;9bXSUf:E-J
Cf)D,dJeUg-V+9Y1F:.0BDAYN:B]+03PH>4fL58bBaB:>0UT(N=b><:fHWP/K-8/
6gOB=J9a7eA0@E]KQ=JX&c/#Q7J:VL5RUORG([>6K()b3ed<4gV/dV6GOXT&C_aF
aNX9;>^/F<03Z,YZGY1G>/E7(RP^I,D(3&SZ1--^6e,(Q0(3?;LZU7JHR)1SC2]A
/PQbL:UB/B-=abffJ4bS=60[<I@)f\YV3I>11A#KS844V(XaRN#<67_.gTRMXe;[
/4@8[#\(D?:EA.IK0XMZVa>DeJRIZ>GF61UW4-#U[gNc[N.2g-=NF,aED_.cQYT,
YFTW/S\aQVV0@QO(B,HPT[BG+MeV6L47[W:M3PPCXS]0YCA7J=5CLSdY(A)2#dQ+
1@W]WQ2M6Vc_.FTOc?85V=g,PDDC-10T+@[KMJCaEI\.?f0gH8DEKL_R,.E.19f,
3-SCP-6b=PMZP/Zc3&]>MV\8bU;G(B=./[^H370Y#^][^.YD)K1Aa&DJXA\CVM>0
V7>H\Z)_EB>N8R(0OV-/Q:CF/Z;6Kc>]BCH45:OMffVN#QU:OV(?c<A#9LHTC&@M
Z&X:0Y[3F3O4?0C>Qg#_g.:\4>ZCHMDd8(-gc^6EH^bGFQ]g#TIH(9gFL.&/M1^<
X@5g1e5LLB1UPN-90PJHGd@6=,M63\:D);6C7ZPJ?EeNZIODIfZTA?>4N7)7??ES
HXS;,Sb9UO]O(]?^C8NRBLN_,H5@UaDXa_df)>CHf(e(RV=>YD?X^J+>L>W2BgeN
JF50fX]&e6A=(0;0VMKZAf?(G;P7C,7E,P)DW3]#OQK#7QaP47g.;=Y&IEd/R#S@
GQJR.LRM+;\W?(_?5ZH:;?@EgDaGdGa_.E_DYMI1@UI1L[ZL;;,XSG__Z9?XI>>D
2C,:)3<-b+c6--<^/,?VT.?#eS@.5))fG+Eb5K-G#6Gc8<U-Q^/.fCgSPS_Ng?)V
80F#SXJVE-LNa+P2RGd)S&\b;I?=&@7.DdQU^f9U0TICR_C)CQQOVODWbfKK;>#7
Y[QJLfeTGW8JJP:W?N9(3gg[I.Z,4A-.+];D=F:8:e;WO=2/:F\>TAFO7[&\[2/?
J&[A8?2G=BK@>TUI7V)bP4gWIZ.f(Z]80B\:TYIEe\A^&4=4-0R\XL5;V>SO_\K(
\)9H_2f76=#?Dg@@a(1ZHRLU4:<4:W18-(=A_1V-#7gTA=EPC47f>FULc/3/,W-9
M/FO680MY@4f1Z8eD6O:K7^Gg_53#&Z6c<MZNA2:A]?XJeJZ\fAVc=P:#G9?ZI)/
dd3f&=S65S?0WXU7-Q8&9GbWI[+S=PPTeOG)WRY5bAX98_QO@eOf.E05MD;DcAPD
Y5K-F6/Y,b>#33]/0Jb7QH8NB,SVJ5+75W:+JWe5ON5^AVVJ#O+7GCQ9TOH,T7<:
M=fEAIO(#)5LB6Q>;OI;3R<8UG]XAYD;+-8A64TD<B+@<CI?>Y.P3J.0:M^F1WC6
X&@f7P)Pa,^6aQ,?,@NScT?(X1+GbJ+a>HRU/TL3FI.cAK3:KUdfS\5IT-)#Y+EV
cYT\/:KI0a-E@0JCN)X8RZ2:CYe>Gb_&CWUN72T#.478<IW\KKdOg0F,TBU)RMV&
a2Z4JL:X@-KDZ>^&M(9][W/^L\IB6=:MYP4KRQe)B/H-;=[\VZIfE@\[IMWTI4d>
f([\4[bgP>^dD<UF;E6.60^#=>1dWB,H+HUR:WMJ[DN9LRH8[9f8N?W\P2PU[HgW
JC:(R13Od9QE#-;.SNF#e@c]\Te/&L;./Tb,;-98D/FcHYQ7f0:?0V908J4V24bT
b\19LG_(@KB<WeI)OXQ&5_,R>:Qff\&51MB??;7(S<]<+<beGRXTV09Q#Q77dZ;+
C2\JH-]-d)_2fEMRbN@N<SI9@ZS_-::3IW:A+D-I;U8LS=?4=GG+c:POXN078@a#
0ePIS\J(VXHbE,W0]PdLDV0O9\\?SIA=:#Y&-Z=cc3M?.V.@OGeFQ0gB5HFeV@T?
>A8MFL.#bHCA&faTF=:,8,G<B,eRLC_SXODGQ-(?+e.1[O+=)Y6^WH0c>@\2)(1F
Z:deEM3Jc;LD?3?+9G5))G3gI^WG0O.e&)7J_R=,6?8=&#H_OCW&4W8]2W-EK^(#
V@7Qc(NQ-Kd002G14IZbb=\^RSe;J0T<7KC4DA.VDW;=>[CA);FMC7>[L;T]HWbA
,,93M(CD8Ydb5B(eY_2>#88U-A.FSZNCLLTF/W)TUHQ,R._cJdXd1V4<(.X>8B&d
9#.fJa>YX-TUTcYV_\R]aaaI;^KCKga,Vd7>9f3_4fd.C6I=;b98\acK=7>(G[J<
@2cKcXU>fYCEeRV[K:e7?._fA/KV?J35[DFZ7(YX1ER_aU1RQLAH#a64RUM++KJA
ADbS.U-,_C\d4eb^Cg/MJG_(A)Y:2IS^[\M0e9SXN7-=A#>8P9fKCSe_Df&&5#GT
,fe(E8/J]1@T0N=1=TE<EX\V41=?5@R&<(2)\H1R#f=Re76VAVUcAR65O8b0LD3P
\ZcV/HWR.fGTgMFPKB@5<R-U,V_5(Q?a?<A8G8-0Qba9DCDb(M;=(86;URgW<2R-
OC4):FZ(MT0Q7\c,@35,0P6)3Cg0db&&P18WfPCYb-(YeVbb3(=2K2@UG\,R6bJX
MCMP6MD)Z32I2(d+S^0^GW8;3=<UN#Bc/AeK1[:eec/]#Pb2G:eR(8UQdLPHP(+-
a<gW;UO&6&20\0P,UP=d<d/K)5KVECSI46DAe?0KH-R2ICS[)0M1A61VO[V9<c;N
T1863fM?L,]XET.Z]ZdGCQ+<A3W7FQYLMJ2+Y/1)9M7E1REBB9<T):;DWI(0P<GA
IX^I./..+JD8]Vg<1U=P#101:9c=#)\g@<C^)7V@HSaB8STHa1UAJB\.L]4UEg;Q
EA)06(YG\3ggAfOOZcELBEB]4:QQ;LL0#bGA]FfT;MF3_]6:#\@d]d1NE](_\,,Z
7gV7Mb=b3S@CB0e:NZDMg+L_CVQU=bGXLaPA?b9d[0LSEK;6>?.gCB3fHVXG85T6
;)U#P9ND9PWLA3,QVgN;NV0X)X&A>>3T;\Db]BOTISS+E&Df:H3_=HYIZ6_K[EUC
C5Jc=;,g:HFfP<^B)?XYKD>,WIJ8ADaH?e8\aG=2b\;(96gV0^g[U:;AD]gM8=XM
XHTJc8Y5bT#H:.TRKH;d4GT6OIX81Q,=@=)RT_ISM^G?#]FAJ-##F?&PCU-LND=6
]>8M&:2DDZE1-L1e)F271CKB?LOg]bFO#G\[B3P[34?dF43RNDUX8L/N.YY)99YE
CKR<?:AB4cc[IS^=B4cX=[FX?ZJRgQHJeBI_VM-cO/TAA^TT<)CfH=(GMBB_MM:O
5]78Z[3LK1W6Z4\PH:cfZ5J?XWPX,e-1cBAgMCR4H1C8K1M>V7IcL;0IGPLB_d>W
-\Wf)6[-W54)9=D,;T6H,SPZc.HXVRUN.?1.TIS91+eE0g8>&GeC37[f=1L5,f>^
?UDc&cO:D8c&X-_.cH.[Y]f53Q&WT\EK@3.6I\63+1GQ0&SOe0#0K>LM7@,/<E.?
<:MRf6,HbKS)cJEIUC[\OJeV4dKNP.URLEHSV3T36ZA\;CL-,P?&//-gU.OD\7#A
X_1c3(B]I/D\H@K@A4cKA563XS\9^gMM+E?_&.#Y?WEY1IcTFbHQIH8@8bTZBH4N
6H\)4L/(?360??fQHG<88.@JTagH.^9I9_\:WI>:TMN6gS/B)ISYe/Bb[@QU7^D0
0^EaXNFV_aKCf7XgJUE[A&DZ13/>GDddc678SUd+c6MD#BW8ZVOYV3&)(;Jc6=cR
((MZ?5G/M\O?:a<\/C?RfaS[/<TM0X&XEWW7-f6e#+CQ1LcYaQX5M4/Ea171A#:e
ZY4b-aAg[N=THWCW&EY54(U2]1.[bNN7(QY]J^RDGbVcQg?@(9@X?N)Ef@-07L_Y
ceBAXdMIN#)AWJ:6)AeZW?8ZS1LVQ5da\11O10-#<T#d+b-Xg<a]67/7:EEe4/:M
TJKc[1@)1LCC;SKM6C7K)#@JeKT:(Z5?)N&ZJG^(&<)8adIU_)8>45YU=F^#TE[;
g_A56PLOD?_D_(3bKUO;(HD9Y/XECC_=YGV8>X?U1U&:8H.Y/QQ-KfXBO.-+c<L1
HKC<Z2aX(WY5J&UI5SX5+c^T[T.=K^Z-]d;eZ.9WbOC&9\Va3^KEE86B5:\A@HQA
5dKD.JM=<-LZ7GNLUfeBWX/@?0,E-.&>LQeWX0M7Vb(?/Yc)aJbA.(&Zg+M@//VI
-=0PVT;e[#B7MZ/g@9;<FW^bSBEH)cU;?d8BGTc?))1LH2+Z9gMROD/bAYZDH]=^
,6Z>:FMAIC8OA<40V?dV);d(2+FAR=K0G-R_F?=J5X])41Y23<,CAAVA5DRZdH=)
O3I,U)f</FVK@0K_:4&4+8)LB@OIXW15.9SZ-(57<1=gKSbY-U9KBD-=C2JcU^@)
L4OO,Tf57cT)H8(XZ#,\P/Nd794X+\5=KUV9<_L#QFJ_F8S=PJ2D_>MEDY.Cd(5/
L9U1=+ZPg+CS+&fJ_?N&;d6=9;T\R8F#4J)Gfc@I7K9-QW?gVL(_K@GK_=aR6>a:
?GX]fc+78JI_RT+-W3XN#-C9)c[,3,-5c2]Q)3(2d7XLH)/b5,,(=(WS_<U=>H;X
NAPBP.RB=2\N6\:;agU1Y=QD6G-[P<DL8BS.G&cU5HN0LMeD9C8\aNG@0)e@,G+(
1&M0@JZ-0f;&aF=g>5?eZd0NSa[M1_aYLA^R=M[5&2->G[:f.,Cc]KLM7O[=#bOW
77Yba@V=.)Yb9DC6WgIg(6WL=eBJZD]I;#9D>dIKO7b..X0B7d)/H1/,b\@@0O2-
L>IJ5@F/<P49GGM&[+dJ3d:F7d@bTJbTdWE2(WE+_2BZ>e@X)CE_1>M7[6.UKAY6
TY@\b@#/,g(?HW2fYJU@;Yfe>0>f8MNU.@JC^^_1>@V9YKD#cQ>=ES8-4#KW(M06
\V8g_2MUVR_#;(P+7QT#_L3XJY1H5e7.>@_ZZRWL,W&_T,,CK)LeVTWA@8-e6\21
.K#bgRZV0DcVZ:L5?eQgX7F6&J--bD91e:(1:./:e]OSLY4f]EU20NNS(G^Bc6DL
4&W,^?1B-gD\V8KT-Jg<5R7Z;WP=5(T^&gbDb:PP;1dU:_=cSaT22/-U6PKHW,23
>N_R)_A]ZY:]Cf8@@OO@Da6##P:V@Sf<DYaDX[f(d1-5L[\6bQE7,gY/\[3>aUUO
_SdHI.:62;F60FCcB_A(WVK&-&Me>ed48@;[)>B@8.DK^B?B)PHBJVf6fQgf)R,7
Y?^4E\@8-;[PD0&c)JYGPIYL&+5/AJdfM5fMd)IS]W_Eg)\]M(@3+W.<LcdU27[4
GB\8;/HS&LR+,FA70MPaN&Cc/XSQ<PT.:,<?G0M)XS-G1YUg4_&5V[I5,7E)BaOF
g=d4SIX76OYL6;^B,XXMJ4Tc_IDXGgOdW6\>0XN_OB=+XEG??:;,6^dS_Pa\;XM<
@D0cg3cAM69-4c/@c6&/Q1g3eBMN58Ya)]>DK6?W<afS8LY;_Tfcc=,@.+NdJ:5g
LF9(/HIgTb1Dc8+86AHTZY49(C-KWTgO#d#TMd[d>YD@DOQeC(M.:&H-XE;Odg_Z
S?.>TWN=\+fNH(7>QR0F4LTYg_4f7=:+0LN9_G;.(N7RG2f>QXD@SB<E/d79AC^8
9F4<G_FVE1OC;]BcU@3FBId)H_1WEXMUH<O[/+,+S(H_/N?BJa1HbMC:<X<3AAA#
:f5Jb&9B<&2b2PM-BRdAJW[M72>JCg\W4g/Ia:gFWX4MKG+QTTVcL\OW28,JY+VE
<;R>0L6D1:fTAOY/#E<\^/SA#;V2M\&2T3e)AJQT[55d<L_TRGZ]:?X(X]fLS\_M
JI>M7\46ICYgW^C0c&[0>)K\DAXT,3B[bW(F3E[I]geN/2U\7Q5dGY1Vf52.E4[D
>W:57W:dE8Q@=:F;+]=+=MKDS>._?5efQP=1#0&/M4Y2:POe3U2?gR]=H\=.b&&W
=0\Q1/5.G#7S7>6WN9UG-/4MH-fCHYb7e8P>F@HS^_CN(-K=1754TPR1eR_\gVc1
dVL#:</?aBGTb932e_-(99^VT46UPRXO1f8,SCS18fM96(;MHU\K.Gc;2?PgQ/0=
;8/>4W&M;BR_\fVDKf;UJ6YLQ;7OW^VC4YTU0c+IQ:>Z9GYS+Ud[2,65c>(P.]7[
R<,GXg&UI:O0\Wc_9Of;5#D(dIE@@.K#YA_)X/WE;b^e2]g++Q^b68a)/HJ?N/67
6g@F\f]Z_=,3Ka#P\cB>,A&F0cL3.S-dV+&B0g]8U5+PIN>fWVfI9YbPLWeab76?
HZN_P8fMLPG,/N<E/N<DS6DM8.B5A;a8&-6+XO7bXA52L)cQW)M_.IGRgD><_<5;
O6)2JS+Ba&VSCaKMD(#0</=K\b;\(MI_F)JWN&&WMWLW52N68f]-?;<DfJLTZWDW
_XK1IE<[U?S-T(=GIB77Q)\U38CI0?F5GPIMC?@E-Y+6d>+46a_QUT]RV/71.6G3
Mde4ge-NI6TXL10X\KZAZ?VF-G:^YfF^g^GB6ZW_8C[b,^]S49b]B_-g;71VBbS]
cXFbW[,;OU3U7,8e=g&Wab(\dF6Qa/B/LZJe2V4:X#PR(c_P;#M#CH><&^E3Hg-8
&&+#f..J,-MW3Z;(.1#^a=Z_#R;f,8O;P22QIcC#27N=Qcf9,^K<43AA0M,:Y^dJ
K3PfeVd+G0]bb@EY8?8d19G0ENPaO&Eg3NZA@>7d3U;?+b87G0Q=P:UP<HV8^eQe
DY5Ud@6,Sf2AS(Q>:7EL5GBITL<cE:PfO;6a#E(fBDZG-G+ecI694FDb,UEON[;S
-bUW:45X5#1/Y3X;KH_e7cQ\V.98S1WY^967)ER]]MdJPH9P>-ZLR>c+J&2GQ0WZ
TZI1gVY,/1TDXB.ATR4Ta;_E_4#Q8=FA?+8\18THeMfDGUIO)3U@1<4ORI+?g=Jb
:G)=(gERNAL;Lg5_]05.KB4C3,[T@dGcBSV]YD>:c20J?LF8&Y,/=T&YC_8&Dg,Z
,dETXS#.f7Z_OYWNf.62]QR?/F/^g[aBA?,[TMH&-5X@@3SRT<>??V4RJMX/#3^F
S-HY@,ZV7LD&XG@<=UF=-JL=6?@G0/6@BeO@<OL@-O88/\dYXR5^#O9L5T9c:F.U
.B,&La0=YBV^:2&:IM&?=DPRdcONHG=:a40=be):K^d3[IO<RaIH;+Z?N89Q?50>
]#KF9<]@47Ng/cNd2N2ee=4JR#2O?0RVI]Q6::B)[I>N0FPO+2X^^Y@5/14\1Mc5
SMaNLcC79]_;U_V0FS=/EIS0M1S,Y?G?OV^EU4(V?7e?4AC\)B@Mf&U\O9RY]_6A
IG\N:?;W?gSV^G<W1[@QYH0gcA-\:ANY+,M\ENYN>_2;=E_[&)T=UUU-,_6MgW.?
fdcK.\Rb27YDYX8,/A96X6&0@Q9HafKKGU-(,Da>J+=FTA/VLEKG==((M7:e/Vf?
f?,HQYb>Q.V^\bRIXOGe([CYS&[gfQ?=,;QT@g,S;6V]PM_bY3TQHWLdD)1edV:C
^FI\1YgM7<aM?D)NR&1cYaOXDH#@K=V#AZBGf,GFCRL3F+Z4cCCZ:3b^5#b_8cI;
dJ3I_fZ&2RbC00J?=aCM&LEU0F9LK47<AAC,>eS^Y2@c+[M+K3dQ?^V@9H6XT6GM
W#C^6UgF[/F?<<O;2M\Z]^P6/8CD8c3O\8JDEaf)N>7UfV<_+]Y>,?<@<2C\gG9<
4-HBaA8_XgTI#3)Y^Y8TJ,D6+deNVfX=_]ONPV0I_[^.JcC#0D;T9P.6G04cF-2K
aPF]ZgC+[E,8QbAF<@Bc/UN+#XKKKE-\17SW?=ecSK=ERbO?TK;8[T;<;fb&95GI
IRJMP?b.J)+bG?HY]c)K2.KJXN-b<Q7b\a>C334@B(FH_1c,_:11<WPf):2]@60d
4cc:H?:89KL/N7C86E\5QJS(H@1ZMLcfON]D?=IJ6<26JBBC>/0H/<aPKgf0<D=L
K\?1-V@V?ZSCPVPe7C[O]7/;P2MNJ59Z\ILd]Z9b8:M_X]7Z6I#6/9EO=]ZeLa&7
]9C2C0BW@II93dW<<FKdU1OSA?5>)/E<O;G)59c?G3&1UdG;?M\DeD\98XM7QW/[
aYAdO(F-?A\GH0A4e\HHY#-/Tb\+Y04ZcAe1L=7-U;<_.VNLU8)#bXV,6.KGJgZb
R2V(3^)(R)d\-@SV\_&KCSe.g5BZL40A8>KY)_US+T>:U6[F^Z)OVXaP(2^45G;P
W#-Hc[6Xd9F3.2V;)b7515;)ZMYJ@_0D]a8]+V4[_I\5.3H:4Z?P.+4=9.58f]L&
,@YS)=IR_]Fcb3]\9XMRD89W2C(,P(^=b#T^_EdEV3U&fNO2XW?5M;GYZcIO/eT5
LA3;))bQ+7R/2&E:1d4;YRO7ZWY54J8,O(OQ6>H?V>1W.C:P4dB;HU76,PU#Sd4E
f2B<?IZF\;@0P35C8ODZAc6BV7P9/:R8g[e(ORBP)2J.19SFN=\;[WN_2:QaMH>/
^5AT1F;g15BM4?:83:f>HPUXfV>LGVGX#@J<R-E7243=ELSYC5I<A_V?F[-c/.3R
XGE)FMa:DY#[))O-/9RWQ\+PddMd5]FMVNJ2.6\,@NRW93A5/>C+D=EWbRNJU&X^
_\SZ3[_TF?EX-U59_g?g5\35L6T[+BO;+&0)AC,g0f^=#[H(^QKPJcL;SKQ@/eCf
SID7gS>0<@XG59H&_;BKT[dA<(/MA)3+X&I-]VOHYQD,/R59VV@+[S&L[[OZ7I?#
P(C-;O@1AFPfc+7@_0YJfL+Nf4BM;b;1.&>;R3BLg]06:E&P9c,ET#Jb]PX>V(5E
gM-EG,)O);:-;NDFb\64b:K6E(VA.CdC8>Cc.YeX2LD8<J()XM>,E7FH]+;F/M@L
JeBCBc?5)gVcP\0^#[K;QXg3D+F7_MNL7U&+)+39WbTZYU)(<Fd[[F-g@F&eO1If
TffA0W.f=_B<MY0&K5&3f2U<MJg5M<<P7L<-e<M)G:79F/=I,)0^2>\/0@O.)81F
-);IDG+P2D[<3E^BGB&VEMR?=F4JaD,Q\M)FMfKEM&TX_R^89eeN)fQY./c8Qd>.
g0NSdI@NKMcaE^d4c-?cM7b6D>I6#.0,E2X<OGL37BANS_LL1[,&HV7DdL_O-+O-
2KfbWW#O#(J+G3S_/gA4R_;#V<(\GZH(F1&FNLQD>.>[:ag[[23Edg.A=TEg&6^D
DZ@/I([O8>7TYe0]05F@FTR3&A/XI]\^Q&^8PJ2g]?@^5e\NU_gYH.]?0R@068UB
=89.RSHb16-LdY0HV)E<4#YAZI/6^T?d#K5M9d<__:;VUL,4Z4XFSDaVMfBVZ-KK
)?0E<1YIJ0U5@S=?MU4e.Oa>SX^G:HY@CK]e674KbE6OQJ_&:6-C20N&@BXK6ITe
e-1.S@:D,TALAR8J8;Z-?40PI)IOYCMJWV:H;K(+(c(C7e;Q]^LeGKWW[>)07L#Z
/gQF\,b\bHNgYJG(KBL:O/b\gT86+P+N?J+]eR5.A9REgJ3(,,?5Q[0K@V:RC\\]
aNaEa<+WJc.1?JYOY&W(;U[;Z4>CTBI01;EOQ:^WU\][^-U)<?^(TSXC;3>agKdQ
WRSTaKeTM,g3-^gC3/ZZ[e)A1[PZ63a4Z>Q?]F-2TbJ]VAd8aX.YcVSI0WKde5+e
+TBBMJBEe?>YcgWF^-=Qa0FODVU4PBSZ&EO102+?g]Z50?8B8YT.TT)(,30:?PB1
F@@[<LWO&P+P;PA3]WO[/V:KecFO9)@M.W:a2A4+Y;?_#C#\TKN#\6H8)>4G,&34
-DBASYaG).8?@>V5<@XF>1P4RaBG=WA&2Y[34da&QAU(6AOFa;[S)+NgeA51<gZ-
1aB3XC^,bCW/3R\\^8Pba-#ePDIJ+1=]/CK5N5=:HHY\Q_4SA6WJC2Gb9++2[5U9
F-J18??-HBGd>aP>KP0N)[-cP[HA8:BO[,X[5VBJB;&6C+:4]\]ZWe(RI+6@IZCY
L_3RY7FCER6XL^?E4M?(3K<OM2S/2cOX(F#E(>V2=eXYG97E(Db?ULC5W/2:;H./
)IbWJ)W(_N9QfTYDfceR92UA7K@P6C5:,c:)/W80@V/)20<(VLL+#DZ6CW^be>5X
P^<@F8HTVRfZdgEVLBFDFOAKZQK)8F0cK9eHa_+d;N6da/0ZB6-11&?7C/@_OBJ_
6ME]3(L@:b2KHABHSNA)F=#+L[;+]adOY:BIeO@,4UWJNd508DcF(O@b_d@e1]UG
SE6>,Y@>,EF:YS[6\\T.F^RbOX.YMc;H94LJB;S?7?MEIE)L]Z&>R#M#G35W8FLg
B_gZ/J\+IDUDNUSHM@L?R/5R>9b1K7Y5JQ0#^J/XIGfX+c(4QOC)US65;b?)V-W[
6b?[W-].;?6beZ[J#8DBK[4Z\fb/R>A@Xf/ELL9,IFX7-0f<\O;>/_aINYXC4?fg
(<W>\5&J8XS#Oe^H#-O6bM1e)+Kd[(W:b3#b1fg,R8EETg)4CgXfgEcf#U2R@XA:
dS&L5KPVgUGE74/EKT+ce(UC21GWWA<S[Hb=E&;Te=1/;P7a2<QYcIV50I=>J>[K
[?L-5KG8\-#J=8;d#@5-SRNVH?3U8&fUD(HB_5Ngb(_0Rc37FI/SS.H2WW&X@;fM
F3[fND5/+9XgT)eI+CB69&DH\1Pc(R22K)Q)b@9?>>&g=DKNNd3=-Aa&CO8-/559
R==<L-I0L^SJR]24_>bc:JUVZ]V5MDVd<F:2FK]M;O.1OagF\;AA)\N<\fWU4:[_
<aeIf?#F0F<d?@W)B(Pb5ECD72cEIH=eURcRX]GL[dU87-7(VCIB-1[Q4?(aNeZJ
PPDJ6eFJIbAJ[ECV6.T57,A@=+/TfLHC07SEEYN7JcSb=Y^WAF-,2P.H&2PR:D&a
ZQB=/,Q)<UfcZeV?R@R6T9M.R]J]=T8SU2D86c6UaLLJ46[U<7:EWfNQf9H_\,]]
UUMMW@ZEWW[[ZTDE3U-]SO#D6d)SOGZc)VR1+COKLK0=Gf_H;I^/W,ZA:Q>,W8QZ
G+TARIYRL9eU=GXb&LdHQ<;5RRfISMQ\[07YK\UZN?dAB&ZN64,T-U0+eXGf<ZFA
Cb.#IWH;@T\I5fdM8SA37ZHd6/QPJ)b6A0Pf7,@DA][>7BE)989fEf6\;@C)Z\=Z
&EN7>KTD?\JYGUHO1gWQ3+D..N3IZ9<YY>e_M)L+97_a3CWC7Q3\9S0\NK23:R+2
(GTO,[aWEH@4(fe#004PXM;8\^V-WfF6\^5N[9CWgR8gAfRR#_b/_PcS,agM4I#a
V44Z2@2a[KH2Md<0S?aaFIBH=);O=D.=7KQ[0N^:gS=&Va8/X@77g\-HWO;K[c9,
g[05AHM;?eT>Yf2QHJW6=@92U>X(C-C0.)O?/+J+;Z&@9>Oc>4UY]_]GDa7I1Q</
O#F?V2Y#9IL/R&(G:WMXS(MU8RW#B,.S-IY[?HS[EL);W1#/G:Be_#FK<HeVe1#N
A/A_BNSQ0U#C@a[STI0VKbW>)@a5/GHN>=F24@SccFOZHU<XE_G_<,.aS8GJ;)Q8
:d#/)/35>^134C^B,76_#.@I623[@B@#8T(N37E+N3U?USC>K>1RKM6,1B25FXOZ
6BUZbNIBPI1@]_:.9cQ;)Z+;7K:W:Z[I(TY</FTB;2]b0?@.T=1=\TbVe?59P^B&
c2(/)[KG_-I@Y[Y?\8I^fL#9;dgbO60MU.]20e]#D/8_@+MH[_&0.^<#&Wd6KGf#
eb/(&73IWV_IPF60Xc#Q?N0caOgMZD2_40Q6=Oc^::EV17=QU>aA]ZIJQc,aNg.N
>HELMLP#W6O(D@3#f/?)0B,SU+;RM/NbDbHd__#L5ee(L19+YW.aS6X:ZR+0:GWZ
(#YGZ?FH&CJN#GEDNg<E19X>JfT^0Ic7[>;X,Yb[@<@Lc(NHW+)O7VDVAFf.I1T-
-W+Q=ZLfL@1E2bHM_XLOZA0OKHgaMV59;99W?Y\f[4Fg985VBc?,?DD<.M]g/KeH
8EQE>FR,e.<:#d=7XC641Zc4;JN/a]_9(8K\gK#OW\IL]DAE]HKKW56T1b=8RG^N
a>_XTTHK4VgN8[>,cYVSWY)f6GF1#?B))0O6:WVO2CTPe^NXVV)WPfF=A\N[-0?g
a-)NOYT0MNBfc/+D2TeLg4JB?S;&)aLB(O_G_fffDF#_b1C03LSd2JGcg#,dD[5E
fScL/2JdWI8>ZJc.LHBeH9@#GSdRKX+Q]2PgQZb6(FWBH]7B[XfU:97@DWP[.S@?
Q8?R>G:Ef-J]^aP:A-WH6[f8)AY.F-KPfHXG7Ec[LI5-^WN]EV>/e)]\Xf@7d^_A
M2degBIe,CVg=^G]ULe&KNVC&2-0G-XK^2-5LRBe6:J@US.(57Ig0f^b-=]D^N=H
@,N4ELeAWQL;;GP[6e+S+EKG+-/FX.5_<a@F.PE5OHORH>(S..)88PdgVZD:M^_=
\)Gc<DV.,#/#C@&^M1^J,Be4\OHdHYG[KUER978DYQ4:IIIZ\4)WS>G&RYT+\+:>
/CcY)SQ.9#]Lc-8c?5JdaBG)ZM_,=@AZX2IX=6GV=Hg,HT=A<38Rb<?P+UKCVWS:
@^MR/M]M5@#]Z<Le;#<dc,ZWKACJ(]I02-H6+<W;IcZ?aI;4LG#0HCYW0(&.7./M
cc#\70a,3c2(^?fO+O7;,CYNfF=[(;P]g?W=,-VYZ+#19)8L)#d\^IcTX:aJ<19P
W@[UdSFX,9CQ3/]U_eBI?C:\5>EK3R)_f<7V<#<0;;,_LG\[cbbb81VBb:#cO5I;
6<c)Nd=F\Qc,e2,<HLb-dRJ2f&=RL)AU:,\]b)/G2R>-;J+N?KJ?K>d9g/E;O(ed
+A97,[]\W2J8SB#O)X\dVZFg2_&C]A=Z,K#_^-Sc>Hf\0W1)3S@bTC/@-Fb;-KBJ
>f90e--J=;HV,CT]W.)JZ6.>d&BZYD.I&^T;5+/4(4_X@DSQHMI+A]2[9)_0CNZK
?+4@S==<5UO<eWACLVcTDLX+a+_I,GHcIK.5.<S]J0a7/(MZg?<5E3YUI>dVeQ4[
32H/B#0_?8@[F,HDJa=BBBVN+0[-e>f)>E]W<90<S3Z/URWe&VEMPS2BZHBGBa\:
b6G&.Jc4c(9KICe+d;6R(K?_^X/C7NcFER8VM_;.M+INB6R,PCb_-Nf47D5XY.\(
6KEAW]1W:+&B@Q/_K9=3Q0=(^3;1(&N&[V4#M>a73G=[?KMI==_.=@^dAC)S-?6Y
;f\0(F2HJ<J>+@VY_D6@?0QMRIP(VF&T[]g&6-L>A3R:c)Ua-[_L[g<[_D\A\#].
2@VNZ0V[D1+TZ#2Z]GYZ26?N0>Z1)FfMX^CGR?<Da[gTR6@370L.ZbI0ZJW5@4Md
[fbHD+c[8R=eFVHK8=Gf;b]2?<?++C29eKHY_CHAX1.5ZJ@PJE=b.Y+e:<>,E:e+
gPYXT\#b5f3TNf9U8C@gKD]D,L2C5&<M)g<ZOMH51+5?/LYE;>EOL<G(H-S7@R\P
8MGag_.P7EC:I0QV/SZQ^DAc;aA)gC/=c.[?aCOPGRA;I:3Sd0F?>A]M3X0:R\T[
:<#_PJ@cGY-6J6Hg92,SSHNZ2:Re>BKf@NO(C@FHfH&GLIgb<WLT]TH\2eaa-2,)
3e;8O\OD3+4ZCEZ\:XP/f34AK1GMH9c]K)@fTZV)dNH/(@RLMHQ&A/]:KPO&a[W.
P=VQf?58CMH9&]NAD>#H92Y/WCQ>5C4f2,Z#1Uec\#GS58&a]F[3_&CZaWUfJRWB
3J;,)>)IEQRXROd+#-GNR?BMf)>/e8)0I;GG,15\@J1<_(N-c7@HKaDA=5@LV?Jg
N,,cZ;YHM>=Ab)ZT<QZ_&8K;?]ZgP)\+CN_PZJUfD\:TY2T?a^Yc>9\E7cV?G3N9
3D>fAcZH,4FG23YfeV6aR21M;4K9Z7E?6+6C:PDQ[Jg.E.H24D3eCO<e^FO>cK_Q
^_c\U5]KT,,/K&,GX2:?1_QLI&.O>@\2T>V+ESOZ4#U,ZF)8O[0gXBS9O>=F69?:
Q^OS/,W-G3a(ebH9/04?MaT\b0+Xb_H(;?c=SXJ@Q<P[Y_/]#B5[d2[MV.41S>W3
#JdA2fWCaU^DYF;>X6aUGE&GMSa#HIH@4Re2-6&I6Y=Q^@d6d)-4dLTAV)Ua\3+]
Bg8T4AMcECg-:IG85,20,(L6AfcA[6S(e^UQ;65-63gJ_H=dF)5_\QSV&Z@.W)NQ
4VIegaHKR^CXSCF0BQ;b]>L+Z+_Gca)++))Sf@\W=X3-JN<Q0c>+:P#@NK[96&&.
d\6HF-RUBOaGKbJ7VHd0A4N(1M58M<a.E^LLO0>3;__E8E=7)[G(6Bd7JZ1bTe6(
fK-?+T9#\I]g[3[(SN\BFgQ=W6f_N;_d(Z;G(^3Xa.#T)W+U^9Y;7cYNXCNe,ABN
_8J:fA@;WPZMe\QC^a+OU+WW2W2EcF#[0[K9g,24\OO\EQFO9gQQXcJ/G+aa1g^Q
;L;T(#9AAQeEO;GU#-0C7#^?GJ2>8gGRe+0[fb9,,dH,-EA5U]4XGP0;B4:\>\GK
4>-bVY-FLHGaTO05,WSTMPD@KWg72HOC:;RC7B._5:QZO=B;)5)]:5O_R@/9GH^Z
S58D#<eK>2NXIa62bTN\@^AE[NRf+g[CB(NRfX\WB5@;<(=-_PZ&e>?->:UeFOU_
B++V2V?6,&:0Y)WKERO1EL-(IDT:WKD>/B<WRd5@S4)CFAg^@@cQAVQE9b/UMUB/
g\W8-ABQI3YfIRCL&eZ&KY/VC\FTXN97)]e]BQV(-Wa\<;J<F=QV56\)U/4F7@V7
62>O=S)MZ76&;3d4[QCEW;Gb=.DHZRZ:F+?2SaHH]?gOQ6BZVIH^AaDJSV+,g@c-
7CWc(fUL\4X9)MPNHa4g_-@SE+fNYEX572QO6OK+,C/:V5W_T.R/@G3\&YX7PKG]
?S8P:Eg;D[C]X84:)eC\71<FfdRS68PTF\0&2MI:N(ZL.7:BRWXHc=GJ+dV1ZcPZ
Ob\gJf]Y05LFI>T6QY1J1]+:Z12^<Gc7<7B5<K\78^Z>cM(U=BOPd+K?2VK2J-b0
=)G/)9UB3S4BM/YHDYNERUf9b]=R]AUf1\&#gU76Rb/-6?,(E#PRQ65,A>3?M#=e
F<fUT=HEB\>#CI\d6_<D2EVLX<GdJ5AFVYES)P8eW_L>T;2/?4WMGPb]>&JcIbc5
.C3eT.,6?7&TDJ;:FM\[ZXd)cP^[)cICJ&/.Q4:S^B.+T6g.c&MR6dQ4:MM[M&A(
.@gS)BdYC]RH>BQL5cLWG,9[,AIZ(U=+>94]B6=)RFJ&[VY8Mg-Td4-9-?G1QF\:
89Mf8,.GK2Qg9^e?a\>eIca<.3T@+[Ag/164RXAKVFgK:6cc>XgT,5/)()=O52US
RTUV_60b0/QKXH,+]JMZKPKgQ3Mb5[_Y2E+6+5J]bc78A<6>G@(ZPaTgUHF)>9A-
d8]V1+ecNFa<I&&<-+e0Kgd.Sb90FT&2QRW>D7V[95J&GU6ZH9^)O-)R8b6U_&:P
O##d)A/fb+LU,+9-ID8d(T^=-bS),9O2g<2;R@aOKT3+=V\DAA98PCN6g1bK)^TU
)=8035I:aBC5DPI/?[@<OeQAbB536WUVUY3>_^-L8226\U&;[@/D4N:UPNYV]2AP
#LQ/f30#=8RGCUHTBJ5)#1D7/46K4UFLef^[:93c\2bBV91b4]35AVC7)@.?Z&,[
cLO/>gPIc__A2;&V+14d451Ld^Q#.II&-:73(7cbBFD&cbSJLK#_&8WE\MN=IeK_
[TLXZ(#GfYX7^>NH-^QC@5F?9/)fX)4adf(?cZHe>IRWLWa?c@ZY4^<#Gb_&[(QG
VcSTH7\-(Vgc[a^60&YG7VV6WM+?d];EdR_>,ScEA;,MbKJUP(9gc(,?7eG@0T>U
4IS1;,(aD9UYMWLVPQ;Y27A4N:6RO>#[9L?bL4\7<G9.d+?Ia?d,RI35MI:e;Q1E
@aZM>6+K&E46M(J2_R0C0X599;@EMg)PY+QMgM_[5/BP>JO<...FRQFOdLUHS-1&
C?90a98fa18ZV+S&;CDG9&KCJIVX9&I=5>7L3J9E?f(:;8Q5WH@6Q1Z4DcZ^f]^B
56N;D[[7@Q<6@Y>P3(e2W[d+3/6=-_<5)>YH\WZ<6=:,)K^?g\N/(,-:g3A2JF8E
D3a=/Z[8J1f^ZN8<G\g83.(9Df@<?^D?b(FPVPKa0@Ff(/.NVAcX]RKca\8?^S0K
^6gJ/];EaAK^2]d&:/0?0R#E13L-N>VM3/5+,JF9?3KH/WRY<<1c.N0.PW.9c425
T>\).Z62[/BKORN,,D</e294c,>S.SY:/d</GV9S/PS[cF1<6&WOH/NUM8,9@Y<F
)F6S+6R(ZK.7RX:)NcO]#X.40V44H3E+/eIYHVR.V^=TYDSV<I5T4a_MVag4JJK[
)FSD3TQUY(VDN@8?&,)E90T]e&)CfUEf,(BGD<9N#CYST9.KRf<V35P<7W^\H</L
\4D4g<R:F^?Z/ND#H@N^CSIgCV(0.42=:6_4d^<AU]9LaY#/_4)ROTFB\HOW@&MT
?STd3EKeGeXVTfY,41,M-QWU+S3(C)\6\&8]#=6=^-#CJV1.).0V?5W([e8U].>J
-2F&a,N/VUIXC#WC?=ICa4KAZ8b20@C<J(F=V8.d/6+\Ue[2&LX/.bUAg[/X0J_A
?,T1?G(,:B>1eX#P/HB<-@VT/_AY]6eN6FVLePbK]#<C7C[a3HHV:33#52_^Bc_9
0C9eBYG7d;FUBWXXO23>=-_9.[]@6FB1<D35RG5C)0WA2:S8WGFR#PPKD1:EV)QX
8U\]P\<9=E4U,VFc:J5LZ1AeH&8Db\NHE<3\dG3N>@=M\S;fTOEX/NF@RP+U.A0T
I]R/WI_eZb]TJVPA7+VV5Q=V1L[RcJ?WCZ>SST5AK5b<USG4^bLA.VZ,V@9EefV@
d]Gc\KSQT^8]B0RN;9T&3)2HUg?5(F,/33[-0NK;P=F):e?BFFJ4662>)NK>Q,b_
&.QJBZ5&<fJEW9<+P7^3bCL@dfgI_BOT&@J=M_A\STSV-e_cPUT9F(2?[8]LDVO=
.AZaW0[?X>LL]/38\d(0E]8[g9\#P>ACN2L>Ib97L[+P6bQ4d7AN-aCR:.e13(0a
6eP\Gc5_eC=c6dP.>bE6.3-7RIf<RX32TJ#9X##>?W&WJAK:.7C>9(;2BV7LYgJ+
^>](:41B:<JXS>,#WY]bcEeeYfZ@=)UGP2):7]TN=PGdKQZQ/A2FDOecH0McbQ7[
eBT7NaS(V_@g?IE>53B=CQ,-<T>/3O2d-M23Z_.PaH0NW\,+4?2?gU:Za_</^-X6
8T7@PSURD;#ffX^WH5baL#Z)6g\K.6STZ\,fCJTdLb28.C6QY9/e1]^X?J=(&W@,
?I]d^][E.&c5@]cZU5#U@=P34T@3f@GdEH&&\(?BH;2>9&W1,bdV8(CPa);KW,IX
eRE_P_,-0LgIGdQ?3JW](f>;Z2YL6Ic3b@#Og(+&a[>GbS(FNe6aRQ_PFT/fM:UR
RU/,R^fD/2M9Y<]d1b&6#Y-<Aac9@O?4A.53A]MR<+KYXf=Hf?VN7U/#26Ha>[7?
A0)[YVI81,f7XR_8D-QB8H+<.#-HA_WD<NKLI(ZP7Z3M9WU//BT.ZbbO\E\MUTD4
IgP6ZUT>XP)B^_C27#G(a&?[NbV0-/b<]&HDcT1e_=(O?&BO5X55#&=OIP;UF=_e
[S8bbaDbV66:=OOK4#BIF\B4SaUQE8H(P7[+\/(-NfcZE?]Cb/7/?-)HT83DTgac
JH>T38Y>#((OE7[2#_Vf</gWI_?UG-_VOO\MAa3WW-[UH]ecR1?,P@?O-YdVT[0N
5bJGTJCPWWD>VdC)99?.O9=T1Z.\DZW\&A3Ab_7(4dOKQNe4f_EOb:(WEc6N^1FE
C.NUS=>YeK1(@7[T,JK1:TUWA6NBMU0#X=Ze=[=Kc5SN?84VE\1TCJT7?Ng]@<./
0/:-GQgEJ]8=HI3JXY7dYUJf9efeUM#UBBFQ)3BDN7_:VQ#^@8f=0e+Ef(\3^57C
)Z(7AME3VI@M,P(_/2B[S(^I-:.5UeQ?(2>_+^H-099FR9<4TYZG6Q:+1@0aaU&N
MRe9&C6U@]KR:OB&RTLHe4)H5dG/FK)@G6)JW2NIFYc]_2QU=RdgHKXA34+eL>60
_:QT1[\;F^3X#d,+N,O5;SKZd^?d/H;N\9J;]-\]1YFeOHLG4++f9+Z>4WK0);(W
@SE]Y]-g[1+1.3d_A=dQgXT^G24JF0#_dAMJ<T9b5&YL?P_X^/&a>\P2NL^1?b(a
YZV0U6=FS)Q4Ia_L3SM[M]GWFU7&\\3eeb4gcD/P_91^_G:,fcfU+f5+O+T,4BDH
@>1_)U@FVe[CO8)KF4+CYI)?c:5J6@DN4[3OcIV_Ff?NT9D\KG_^IR(OY<V[\f>1
N/H+]7gH3TE0b^b0DI=D83]VN(CdCQAb<++()M0TEDGA]28bJ\4)BRZ]ASJ),e/I
a6NZHN;Q\FIUKI0OU<fcU^>)PKE5F8[CF(^X@4H_46QcWWfcWe/22YWIH#bM>(;[
<J\#,Je3#BbLCN>A>52X00KO5AVHX\\>8U?\BZGSGFAfJ:d8O3G>5Z>B+8g]#34T
3^4:PA3Ig\W(MgVgK<(@3?K?9_BE4LNH=IZeL<9+J#T+X^?U/a@3>YDZ291_B-S)
CO+LdXG;EcCU?fgdHcO0+Z3e+^Nc?de)XHS<EEJU)_c,8)<?G+eI,;^eIWG.>f/O
L\Y/A&:Z)48T5RYee/NeD:Q.I=L[64G)Y\0FHKHc4,J^^BXO+3b]KIOR9R&^/LNa
/MF7C#U9L+IER>WgO?b4D6-W:F;3Z+a[T[W[&BTO1PH4YdZ0@/W,6-)=[6af1KA_
0=HIS>J[O(&d4QaaVCb+T;G0-2IKDK<<2,UY7#\e[U)T)-SC/N8f9\+W:=N.]LJU
,QBcM19aU=VA=/WfHER_VBb=&d&eK]2E>#bCY9UXTMdd<2B_N76WTW@XJK3VbKF+
>Wee,;HO#,)0Dg.ORVSB4Ee4D,@=Q18e#OIcEW=_H_?M+d\_^(V0XUg&6.7LIXd>
f#B:1W6>X7#QQC&Qba(UZ>EQ+A)IUT#\ad+AY9<DC0cJ8Q2bO,(2?VWCT0R35RF3
#J.(f)b_d[C8Og/8E0/UZ?#W+9U-?WT3\:bZ<?U]4S>K]B/)AL,,=DUU)_H1a-<T
X.WeX4\TTW^[FJC/#?@5&]8/Z&R#gbNH2=#Y9_2CbdPf\W_G)W6f4\^4B?aATf3c
FA=Z[4)HMM:_BS2[)X;)R81aVReF8T8B\3d4D:V(\J>KZD)PU<Y)GM=/.I?@G]P/
U\XFZc,2P@BZ3]HB+&#cRXfSVJF;8NDZ,V+S9_/9A0V7T=F(5aO.(P)[\53NEYTc
:2W,M56/U@<SdT)L0CMP_W5^A6U,DOW[-KgXg)05X>5X@4^BT,6^I8V6A=<^0CD.
-fIIFB0PL),&\4-.(CP?)/Xa3d0@Pb=B@+/dCU4B?]3TC&SAWRW\56d,ZCP_Z5NG
C19(_(0MIXSYJL8PVU;/CB)WRCH2GYO/Lb-Y[8.81F5XF38GBNeWM90]H)ZS5f-\
K,c,Rd_1B<#e4FS#SG2YH,U8GZ2Z9_bNQF67T6,BaUb4IFe1F.g8G_NLCNI,\YM?
b+fEcVTS=M.]?:8TS?IDXLY0fa1fO1#>SZY-U1Tf&+9BY)J94=APQF1K4Q,&F8c<
MSQ-8RQK1TAT_5T[HQN[ASFH1OaSUR@:;g0;?9bG/aK6U#Q2C4e(NZ:8U+5e1(8Y
5\b.ES<WYaLQU.dOSgTNDQ&5<W:(XT+/Q<7\:7OdL\,C4\=<AdRe\NcaT]&E^5@E
fc.e>E54=ZO+KF-S<R>5#GPfYRg5DO#M)cMCK+M+X7[]NWVLBTR>-(4_NO8ZP-&/
.AA5UcC/._F^3,85Pe-L>46TPZ?MP:670J5Z&KU<e[C/2(&X<g]:I=JB_(-NTV[M
3TMAQ5(POaIF)-?\5RY2DE?96S(X>&)WeW2+:;]SK/6(D88(dT&2&P517>)726c^
P<?VQE6@J;3+R+0T7,?<FK\HeW/b/a=16CY?Y+1]T.2RPf(>2N2BUf;D>IC;FUc)
O.NQAF=O[Ic6Ib>V<0,P)3S@Wc8CW8dS-VeSW:_Sg]K8P->7Gg\;d<HY#e]\I#G8
T)IO&6V;S\8409:GX/SB:8-T:Wd1<^cT/CP)GbUdK&T;G6(-NY-MI84&IAKZ1;BL
M:1Wf[#^:#CM(O6(g@><KNE5ZW=b7ZLC?L(Gd_B25:O;c.7.ZBBW(?54D69M+.X0
?6P=MR=JS02_O:8T<8MbWa6XDDW](M9&4\/4TcX@X,26,VK/2>XY\=e;e+WBa3BI
&]Vd/M5B1cCPRfIT)\5Y#JX\FVAZB-=4;X_d<D,95&)M/1^#+dMfK4,b+4J8>fLX
A,X(KBU_DaOcNE#P^<G,V\8I3:U@g7B(\d<[L:V=S^-;RaJZ>?)WE0ETM.&;]fg.
/P9>71Y4gO^C<L#>JGY?>Gg@2U@5O4T9PWd>=H]>.BgZY2UQ0Y(ZFPA90<D&-4#E
0>AJ-?Me3fUg.?DJHOgAADb6=SKX_X5H5KD-]0G=+N0,g(BfTbJIA/fNQS;,,DF(
NGFC.c<_&G7>_=4HOE91D4cL]&UP]A1;K+2UP[d1;T7P[aP=BX>D=UUgAYeP19EI
KHZ.)Kc15_;I3LB:FKO[#NSGL,2I=5?7Zd&,d()&OTUcJcLMN=cTA1LFIXU1P.?a
981fV7A=-#Ub\H=2-bZ6@P&UL20Z/SHW52VQ@DJ:0d+cB8A2T\/I_8bWHc?Z9YSE
5R[@@;K:ZB_@10>a4/<E^G.+&(_dEB3X0ggPgaTTO>PQ7g1CW9])JS>[bf3FMAMB
,eQ/b.A?E24LOILQ?R+>6aZIQ?>5Z?YQ4a?HD2a>/cd+0^TOU0ZFRTP=ZUBB)=@/
#])TX<=7J):e,1C.\@(J.M<+P=#(_]^?/Q_W4T8WB#c,X_[\790WdBd#NbEV;<[d
+M]/.[DUR#HV(5P3=X-OC5P&Q3:DPC6gWW<A:6A,<;^,H&<XXR7J1]?C?bCBI\L-
7[QT/ME81OHH(C#\Jd6_cY9g6.?ce<GdVW/?;N31QWW@PII94Qf)JGb<_VcPE#A&
CU&B6YaFEKa,O[a)a6\NYHa>-O:JF=VT0DgN<A/5IY[/Z8fN0D.H[SR<QMVW(Rd-
#/81V=T5LP(6BO<@)<0f&0=;c89>/&P\aE#+,?/I]3:K6SO5X\-&c:aPI^(+PKbN
+#[<fM;)T@c)9JY#e_#ZHcHAd_<+L70MI0Q@KMD04BK)[.S3<8SNg)NR]+d.=/)@
5e9H_]N&b^536fR51.&c(3IeM6)#8aLJDg?&L^9V._(I_T[8W)^4;W:b8=D>RP\G
AbUL98=b0M&7fX<MY90H:)0A,.aQ7A+#bKI0Q[W00JN<E^IA#JbaUg?B:?=YO=@9
DDK_M].4Z6,IF[Id8[AON9.RW]L5/D;)B[^.<44:^2+LFaYG1(c]TSTDJS5)\[XR
N998ffE[-#F?.JMA<cVI_LfR&F8D<+G)\8:HZ7<^I<L6aNK.>H(V2(ZEK9\H\La4
/_I2U4\gSSUMOWH<PIPY,(D?QCCNYC9&IUNbV)gPa<5d07J^WS84(\>WT5;[5:HJ
U](.;Kgf82&M5US#Q,DJ_Lb2AHV;GZ4M@+[GbD3gM(YUM[,M&:F7[R]+0>-;/QK-
<TRO,TZ;10^9ZY@?J7D&2774E&,EL\U=fY;GD/>9D0RID<L4N0WW[5V<QFAT9Z=L
SYO<VfM<_((0XZ9Q[;)#.5<_7@fS&>3S_&CP6<Y+[NG;3:[YTP31IREIS?5Ra^0Y
)@JdS/dYM_]1)#00@7NAD[^R,c;K/J8:)6Z3]WNcW5:6&=>0/26c\@R4UQUUZeXE
(/T?1<P00L=aR.ATEQ0OP;g^#&Z9<Ed&.^Sa.e;(A=>HObI:cb6_(2=?302[K[/7
GZGWDHca)cY^PfHL?8A86VG/N-7[>A?NgK3C[8cb&V5_[I9T9,0O1;\N]fceSQP5
UfH&UaYbV9VgfeaU&JZ+7K8;[gF?/aCG^>Y4g20#dX.BB3QJRT2XKBQW+YZY9ZXZ
Q>#Cg5WP(]cfYc&)S@0^\66<,H9,GU^E8,LI<>?:#,=\C@6IB:^V=DGT>+,L^>NR
H4&aYK14e475/Bd\d:HMd(K-T8()8PI&7Z>#DW?31(-LEWc@_?G9[4PKg#gKF^7O
3=9/#aZ+?5XVWIIdF)cU)N3Q\37a78U]3ER-Ue:fQ=LZ5,2;/.[A_<5EZ[L@2<<b
a]Y(SZe.0(O6Y53\5ZICf&38@W/-A]\@[H:]#L-(BK5J;AH0,f(6g<1c.=gGLaUI
-]NHI1fIIbZ5GQ<]4YP4DYTVE9RLVF0_4=:I@;2I(?>/Jc08OX+g;TMYQa<?fd[;
]-K\A>)H[N3)PgS\X0L-B-dB>H5PSaFfd4&KTZA4Gd95/EC^48,Tcg]5^bZ)X(;5
F5-e4(#dVWa?&\U7;:HHd3#+a2=2DL]H&72Gb;Y8-/HD0;L+7W(e/3IaXKUg0.5Z
;fY+fVgX,6EDg,E?gL^6aHVC-[](U]^K+0P>&/&eT8:ZLE=-X#=8JY2E8>N^:;aV
.:YM1bI8X<Y;G6)=(@Vg-J;Z1ZZQW)TfPDDWA:K^HER2-U<X#6T)G8FQ/[]5G.NN
;OXA<Z2(>9CAC<MW3I@1\I5KNf81]18<V,6N&DSgXKH2S9>JX#_\NdL1JO.0LB^I
2O4b0DCSXB3Vd/;5#@WaC7V97,IMJ+]a)&McC#/[\46W5:,e9YO5^;(VG[A)Q.(J
V=,]0AceB4?c@Cc_E,],B=-RN3U\SaK<@XPJF15G0B\9M&7X]C/UXJQ?]0UDR87Q
L;g2<?aW4Y-JOg]<aIK/c2GbG=S6L1/J.3(0GT[fJ2+X>_5WRDQO=b(]I/T+V81[
L1A]7?H#f+/S,7PC^=I^3SB]NOE/;)cMg9MVXe6ZZ9Ga_](R6]A_.BPaWF]T3HDX
[U;,g<XW/K2U_T\..Oe7UBS(BWRQ[N=_0)/SKAb6F-F[JR2C_ASb=Bd:NGL5>](K
,?0VF:U1ZN7eR:1Y<E/cRE2HKdFQBgYUT9ZQBO(dCY9K<]/FcPdOe4YFZ2HSWHLg
)?PXD<.J@Q@+-PP+>TeFeE05>H?1d_YDHL,CMHM6PU7[C_-M\KSdNEUWa39QB763
I8=/AP=S0<LLdNODSG-\PWRN9,AO:EJNGefMAXI,XQ^2O&6K:\+EP2\)^_85:4?I
00FZ-ICT41e/Z64)Z3KbO9,4fQUI2HN_6K0Wc163H8&X,T7^W[)K?]2F&@f;^:.4
@C92;]1J-]EE=DQ]-WUV1D:Q]R1#=.J?=U(-#<e,E27^L-#eCM.U8_#HB//f94Q>
K.8KTe5/8I-L#Mf]P7DMb^?2Q-Q;7-G+d3&N#2&5[]Oad)(2,b[[ca0UK8W->O3O
d0N[FX.49&X@ZOO#<.^85)(TYfY:/Sf:=\54GK]QF&/(gHD@AKPP0.@I@3dF2_?S
OX<&@X7YbA8)\62WGJM1b#b0]S0T[(d_;R9Xc?(^?fDcF?b)eKeX::,\[C9Hb,gX
,g1SY._I869=J<N>bED?7KgcP]M:73IEdNX992=)35[(W5\]=8-I=2\/.9\B_7>,
b5]ZX5YEfH_e=d=)R;ePY_3A/Tc/734XZd\[eBCCZ;BE[cgddDI^LHaMD&)6HFBS
SIXbU?9/eM()Yf,6b52;2+dfPJa;R1eBWP,MS/X^U&cA3:[g[N62T6E58QJ)VPb.
(\K:^V8;9FA(+1OLf@P8aV3QY(W&,(6+9CYY/S@G-HdaMFD=Ze>WW90GgUFgW0T2
WK:CT2[A((AaOM1E8<SEc=fCP2bLcRK^Y2(bC3SZ7.dGD>&JO0d=3Z1U>S.<12g9
X3=4881=Cc;)G.I<AXVd4@[eGHB.<D_]E@QOG5AdZ4]NABcO+QIdUKDfRE.f_17Z
_6@\U=S,g)UE3FFL_\Z1;8cdaQ6a6@fbIWf]ST4S-QJ&#S>>@7NQPRXe725QY6_+
FeM<ZDD=S1@R00P+VP10(DH5ALQE,?J]\1<5,U3::61cL.#]QR(U40N-WLcbI850
=20JAXKd]&YeH7^([d+IN\Tf=a2aCTBCV;US@eZIDdUbENK4X>gZ;THWMbVCfIJ\
_+.DS9-4Nf\0N3FJf1)[bUHX?1.bgJ5e@G^-0L8ALO.^JIcSd?d3:FHR4,)LNMB=
]^b_T[0_C;4CT>4)R30c^,dBAJN(=S1G_UVG&>Q]=32-G;:DLA-d)=MbC#?\V-VX
MdH#..Ld<g)O]X>.-H)I__/H)IFM.RE6MFc5ZEN(#1O,\B_IEZ45,e(88(&,NeMc
YU)<3=EdVC0BSZ[:8/2IA,O::E+__D/,cg^IfFTYWYPeT,c\IVRID3S.U)OK?FE6
=)ZAfGP,XH1[A,da1=_bY_a/4c,=A5XE](LDUf2NP4?N_2I9#1d1\<A<Y9XXEBbf
TBC?cE=Z<DSI:D-][Z&d5RFPB_d=@L<Lb@3a#UXeO[/c5g<a^(Z2CP0P5-WCT:/B
=SeS-KB8-0W/=LGQ]E-)_@5&L<EZF>6Ta=S&>TB>HP>]^++>I?W-HI7?HLKI.=Z&
^<a;Z(XWCF.<\=f?9.\.B5T^_?<](OO\..H>eBIADAWBU5EFM;=7g,JZdYUBGWV-
D5f4SP;1V[d;+N0L.&IU<g]AFYc<ZBTF;YUW:23ER]EOb.MM)eI8R60I.f+:707S
BU_Ob-<TT:\e3gRRL_73ZWHN@(Ng)gC#[0(#DPDT8&^-]ZEe:)KbC[\9]YPRY-fW
71_;)0>fcDfV]7;Vb<\TJ=](7@TbWG>E-#?_QI/6d#][J]@Z=:5?c)426/c]BGT0
P9d4+6P.>CIRN/#G?gVcJRVQJ)<L93-dEF>,T/f(BK-@H9,0[?]0Yg+=3d/dcJ:V
H1/QTI)=[b);+<+UI[(R^gJS=2b)Ne3#4C,fd?bY2>^B]Pf0#41gKMN13JKZTQE&
YK<f#QJ-W0/=28IG,G(eJMVa-R9SfF?1CN?I.B5&@\BXI0fKb2?+GeY72IgfP8aK
F[b<I<aZga^\UIS94D7OH>@ae<.EEA7FTA^N]5&3><TVY2L-JN0C6PM\7>4#S+8A
O?g@(b/C^FB=52=_gK[\0L9b)<36Y.P<15XBVe;?2VH,cI;c&?N.O_GT[3JUZ,cb
eP<d&8\bWX&VQ0&6T-8V9WdVSbJ6LT3V1AeSFEHZVd:VGU].&-fN2S1-I0Fg@?]]
c#bB6bG\dO_._Nf3QWTa9/1/MXE6T&L)_DDB?)KS63D&[>Y5A4OCY.K5TJV0:M_6
.B\8FGA;V/_+\53[J0#9I01/2$
`endprotected

      `protected
(2f?EGLdRY+>=bIQ7S@QbOZ+3:<&8E-G][cJ6QMZN)HfcI]#SfVA()VTVD@+6-(]
+;\K2+gDgFJg0Sa>I2c-BcZ+6$
`endprotected

      //vcs_vip_protect
      `protected
aa)fW@07)c81D11V]c3-,<+_]eHS@/<AcZXX8]]X6S>+UBcNK#a2((\AS_WJdc&M
U8T8(LG8>#[;IWgM?UIbb<J15X;7\\85,YffTCa#]#_AX+3/BMF-6Y0?ZMKV(H[C
PN#;Q-E:dAR.S73T_<a#E<@0]KD)@1IDc\LSWR4OH+X4XOL&--W-\[0D7RF]GF]>
WOSa<J,4RF_YQO;&AWJI]f3T,@/ZZX2e3BE:fV3aQeLFLFFW>(J-.g6AH=KUUJMW
7#a(4L&9.A,cI1AI],_)D_](ZS[0/^]<9/c=&/M=+BaB.EgIGZ\)#8dcV[H6;Md7
+:\&=+4b?4Sd=3N1C^LA,(FPfTO4L3D6TdR]1J9&]>WaTPI?]Qa8F?KKe;C9/@d&
Da[#6a0eEd01N5ZZOLd.d<V33bG:D)\[#2Uc>0M-/6\4UIA_<4A#g2IK.6RTR.1g
9IM4(WKdH1AQ^aX05PHQa;H/.4PWcc\4@8-I9CXU;R:-RW&OJLb3.4ePCgWd+?KC
E1WQ&F/JNF#fJ#1:P[K^]2/bWF\3@^3[6^B;2\DA.&Q)=22[\b<=N2VK:26^Ee+L
;HM.dG3>>_GXC366BHcK0C3@QTaQ9)X?9#TL0B9#RQDI+MNQCLdZ>a2Ic,TY8,]O
,8Qd?A+c-4Z5P+/\\]1^Mf#<PeJEb>9Rgf^Va64cJbP3]@=MI]_g=(7WG>[[IG/g
DBd+\4K-3Q1J4f0(:cJ7D#K[+6\6=gV(#==G#.YB+@\1dd(Z80dA_ZY1X_#KbgXI
Jd6G)[-<5X_VgHB>DRc7f&9VbY)bF->:@2bBeF3FFPJ.&TXXFEc_8F6),ROa5ETT
02NF^M7/-6QF^AdD]>-N>Z\SA0,fd+<VY7KRAE8L<5E.Kb_g;,4]W14^a6.)<cR\
+G1C#[,MD2eIWK:N48J1Z;H,WB36a1;#+cA6822:dCaTON]I;dZ9U[3O,HDR^Rc6
7A#7eYMJWLFVY@;@]&MJ8G]M05M73I\0R-;H.YSYYOJH@W>GA@^H,9);7@I52?5f
.)fc#^<&7BIFaf)P=TL2?SELW<K&XNPR]AK\L<HLWICD/E3a5a2G:)fFeN1\1G5I
/+gEQYOJ[=D0J0JFB8OM4+L,Z5N0>a2>E>MRJ:+/U]Te-aaN&d_a)&2];0eF,RC0
IWT?cT+fLe)a@^EG-QPE,25.;gCAW_D/ZRV3ZcE7N?>CF9::df4>URADVJ+56AT_
_?.:a)BQ#NXLSLQ@3d4/T>HJ6O2BA96SG\-X,EN4a)FYVBgFTV-?7gIMb,OG:&5,
H]K/bgSH-20g@X-1RbO(R#^If:aec;.cbI](de-UB-\#23T7]SQ>;P_7UbKTUa?d
+)A&9Td_LD&T6JdLN@)#Kg7V^)<fEbQFCa\60]f?d<T<I\GLN5NKfQ>+I62f#(>T
9T&-J;-S/ba:S8F3^:<bPd]ZN9<(5Xg].PDP_QK4W=4Y2UGFBC_+CGR97^KO>c1f
IH_S2N6&g+W].H(UJ2Q9gb@4?3E+8+0@_g0SC.SU4MGV]^>\/_b#EQJ@M3U2R-)B
:VJ>8GGV+dP6c30FJ)Xe,PIA:UX4D1VURXMS45[=@f;2-[@eU^g#PL5I6D.>\,?F
f\U&#3F.aVWN7<W9a^?:=1)4SB&B]._6M72G\T4FNH+9W)0e0&@_ga?MIF4M:Ce(
>=8+^#4<3&aVRB0ca7-M.&LFJ5PID6LLWC&cLD==.;VB3]OH<9Y89+V<SA;\DSBQ
/)&0E_F7\QSCG.4KKc3Y.I^L78@W_?+b]PHa3Q.UUK5D<Zb[U@>88K=I:KR-(5,1
7JdCO0eGM)YRdI>I5bTH2HJ6?^ee@1,eDFA/[R\Kc@35X])IP??e2V7<[d_C]e?<
5_8SQd<W?\-DNFe-a]=,JId^S5N(GS[X;:)7B0PO4:A.?G7NcFeMVN5]K9?TA7\K
+9(U-L3+VF26g,X)R7RGE1X^CeR/OdVUF^E>=T-AP]\X6Y1@A>_2997N)A_SJWdB
F)-ZF^@_6#BC;8)YBW3KZ1>7WKeF=D93R/PX6AA47/4d:J]H8#KU)GF[A5[2FH=a
[g2L_XeW#TP:IR1daAPU(+]J&S]#fPOcON9d@QVW@L6bIVGK@AD412XEg6,XYH?-
URT1cFd@Xf]T8/)DA/[RSd(ROMfPVg[G@KG:N;GI?J>cB42]PTccH6V#CKAC&QUC
aFT<Zd-aL.(/K)]=F+#&Rc194\=Rc:C^_/c<f[Q3L(&Pb&C#UQV:M-IeQY_#;G3,
94+Y?>,>&dEeaKAS9=3a:ON6>S_e(;G)B@.,3/)aae5bTH=(aVQ))NLYH>;[f^WU
?a3,F.OW/]9-6Z6WYCcbcQE++IB3_#@JMXaVX2VO[K@?#F5&7W:+B7V(#.(44^cZ
aQ2BK952fc^#?M=V.K+?0G]-&DZC-Y,E4[/J,NH47SS]0=O-O3)F),e[6gPcJ\SU
a?cf+\OH]QJI)R)M&0\T-62gOE/QV&,6?bH3&YG\DQM3S7EH)=PG95c9G3ZL[T,:
Q@[]O1D+&P^?]>?MC5g,Kf0R3J?(A<ZP0?aELbcd^MTfVK:Q_90)]?TH8A#H,XL]
-);KEEWJLP=2\P)W^O)_O5_#[K10AD865EM/^&g5)6a[g:6SE7QBJ/)BU@2N,>9R
C5_/JO2D>N(.GBT1\[;R=(-<?e(,;DaB8.:fB\aUS@_@#[VRTK3UL;Y90?[H[geN
d/_<c^U>ZPW6@X6[fN[Dc9NY-/T_^.U]#FbfC/L#?B]&IEF934S7_Hd\UJEN1#?g
[D1HHHZB/.7#JJZTGWD@d@D:;];IL/RS7(UO\5/DbO;NaH0^F+?>MNQdc]Nf4fD<
Z1.;_]DH,Tc1UY,44KYQ_0cIbR8E,]3e6L?Xg/OLN;F0dXW-4>5#A-ddF_PaKC]#
VTa3c(B4+<?=UUV+4]&Td9bR=/SZURKEUDSC;FWO@CSB5eGNH<.]ZGR&[AWe_0MH
3gO&b;MA[a;AO3=e&H[_7U=g=YX^13PI)a3BFU1U=dJ[<(/^S/eZO8_)DS_Y]e+<
1SPSSR)Uf6\RcL[A_A078;VZAf1C5db/,b#2Ggdd>R[]Ee>?R(<)4I[.Z^eQaYcZ
KWUIB-]L#Y01ZK_MTM.6W/AWM7;P.ID/\J7PYH][W3P5f(D6CM3LY<GeWI3-O@+R
S]aB@Da63VY@:G:b.KEONJ[=P.b#.84N\@BOI;PZTLVC4JI63IX.3S/=YW^3TW:L
S)#0N^\Pf+I&UGfFQGFYe5^J]=a4?g(^I<JH4K_E6cHW9@O-;BH/FGP1>_0&)U><
AIF;&+a@7dR9/OUM?X>T7;EAAMAJ.9b7Ofe4.=/HSMJ?T9\_gPFe@\a2.37_dI;<
2X?/?;4g>1HbJa\_J-?EaH_4ZWVF9g]:A_Pa3:]PeU&V?:Oa_>/aZ7Z;Ecb.HYb0
_:QY9LA:OH/UP-(LAC2Q2c@.9dE73dDc=-5JD;CM-BV8P>5UX7:N#WG90?IRc,Z-
)Iag?F0XDWZEPO+77\(4fKLe(RIR4>K,Y:]FNgYR5GF_H17YK2IFX9P5MFg>?+-^
M@1RN;bJcb0WGV)/\f3dRXUd,5\K=6T@)Qc1A.c4d>gU2K+TUQgNZ\1/W\_&7U52
Pb&&c/\0b7YL029^49c#3BWP#OVbTXPAMLW(_]BZ.U](9RN2/\?<<7&LG)T5<,LF
KQ04EM:f[SWZcV8]gY95_bCEW+E.FL1Y[7M1X0>31>f0B-ZEN(C7;AH5P30[,-ZV
FLBLF;81(Ze#/S@b.&3M9]V1C2UQE(W,)^50&Q,BI;IV52KYE?0OT?BUfRG11J[Y
c.&?+#]3Q-//L#c0CeXBQP)T(,84M3_3O+18&73#b@R#DWW2Ze=>9K-Y>EH5WJIM
g<6<^ECf[]0R1P-BG##QA.M@V_3Oa]2Iaa^]LO_2+4&Xc?X4;[4:YQP6UW<3QKSK
Ze/E:Ac2J@e02Z;379G[a;ZCdd.GXI;e(@;E19f,(AC7+g_gTC06_bWg=P6708&@
&):fSf7T221>E)g08(6U27Qb9&]<B]3K0,2B+PfHT&B:Y3_8<U_ca_O&d#GQMZ_6
B2c5L3KcR^b0GG_1M_&F5d\0Y1e&INO9SAH9NCLE(@c0>:Q)>OR-3E4XAK?=eUK>
PZ:?RTI9]S-PaGO_;XXAH9Q&HF/Z1-/:M:9^)DG,W&AE^6G6#8_6R/K&Ag]W]D36
FPNL1F^4?4)WSU[OcHN.M5A3bC(Y[@6J(;+]?#>GBeS2<99^S_^^ED[3YS&WDG<,
Q(RHPd&;U,Q8-7:aU72IZb>/a_(CHSCbC4PR+IaO-<e+Q:W[Y8K(g.6CggET]&>E
/19Z[3BMNSf=\\1SDLe7IM#T\G@V,ECDU_.)^JBWBMGQfXC9B(ZdCA6Z=(TEF+AO
17+XcZ(eY^[0;F+e1I@97^FY,>&-Y[43X5M&W-]OHG(M^8;^(ZeVDef-;J6Fa-Yc
\]2HK8S913G]WARAd#E@_Yf8U/J>P&VN#Ke&_L/OE=XGfH>5ZZKJ5HR+:c)&L^0;
Uc/Vg,.4(/R+Lc?9>Rf-<G(E]V[=(B>-0&c?U(V)8N;fg3#>=?:\&DK?,,HI#e_+
SC-bSVRHHG&74F]bAK3/,<EWZZ\_9?38\XZH&O1:5>=N>=aY,E8TG&=,Pg/H>6/N
F3CDg2D7:S_Bfe=)XAMfAYAPOABH#356)[@VQJcIaWVSY_9U?=NS19/dZWRRWdCA
5#+bd>ZYQ-+FF71Jg0VISCWf.b3AVf3?/VKg<GN5,TA8V-/:dg<QHe3b@VdHKW(d
M#6J]W,/-[L\3&Ug]4#2\/EfXY26dM.6/_&C.S+4[OCa,48[76S6@9Pe@7d_6A6d
\46\DE=D893-2_O=,&)_=##LKOH=CK4&;O4_Q?)eag=N;8KUI:TAQ=.gc3XI#T.6
=ZD_a?RYdD^;E?bK>6;5_Y;X),KANWXG)]/0\)6K_e?1F;WgT)^^U\S.;FeOfAa#
=W-AYIVba-K_[/_;^T90=)/C+672EKRY#+O.eRE,X+dBLJ,fGgMaFd=VTWb\Z@Z]
H:USaa?dXQ:H8c-.CVHFZX0(I.(eFHWg\(g8)Ua)c^ZMKVHbU0[X,?)0:;.2L,2(
+5+dKRRPbNEGOV)ZDecABP>W8g3@W;#)&J26-UPP029&<0dS)?U>-5I(8&f-A.Ka
f=H4;fZW?#@83fHAHZ]^M7G:YdA4@STD#&.9ML:aJB>O9BR>HMG5:74ff\WO:,^0
d3cM9[]NZ#I[?W?__b#8^[[RKI);C,0:-75FCPED8bgW>RVd[IIH@]>aCC?@ZD-Y
B_056_R)WXa#6N.fgESG>XcPc,c0JU8#4H6RGQ;+/ZGV&23ZT=\QM<V]YX&+FgI:
_KNSY@.1.N62HNQN0OP7[JP8+cONNN^B(Ja0aT&;67e09f]0<H\:L]<H,a]<.O<U
/HL_<UF5J<d=+f3f+e@defeG?I/d&?WVW.HEVM-K+J,J-/CM^H02E5BR9c_35QXe
(Y]#PRDR:0DZ&I[IaI[^SNGVGQ5#T8W<M3Bg[4)Nc;-Ic>8O0YQ.L1^>[bB,Wc#J
16X2JF9DO&QXKO)9&IF/R6gP8Ka_/T)N/f8_TK_IK.J0YV52SHETZ&:Z&8fQI\Y.
Q\K3=8I4S51fH-#S,ZV02E>,gTgRL?QQL8BO^M.ZUU_X8_AUQ^HMX,C,-K98-FD_
[&KUB.bX-I64;Z6>[L>+Wb7<-.006O4AFT\<3g=D3G3VO9OS1D.].NJ\5#VIQMcV
<YJe#O4cRHXX8O;SGST>KfFCA/2(ffH,:/g<4Y#9)XB._f41CF/:ZW>YL)9:KHRE
[@:VHI0PX>3>3d)F2)#WQZ9OUQ+AG<?CM@;5cCM1e:#]CS[4-feg7-d7efF7S.Vd
9V2MZNdGZA583bb)RfO\g<SAfe/bg_CgIF^g;[\XV19\g+IF=;15M[PaU)@V9d-E
b0YVKQQL&7A47[f_]fcA_4I-[@9<AY6M/K?d)Y&+33)@&d]Y66<b))>TLYe2-_GM
0-KRIGK09FeTfL&(>K:Z[U2Wc_@TL?#b-BF.,N(B0aBYZ9\/BUc(F^\RE@(+=<)O
7D[?Z(>M,?LG_G@BTD.J8&PVOOO4QU4E]0WKdd>L/8#dd9=+W>H:DU->a8?L&Z,1
(JS-R^fe#db+_EW3=ZF406#C3A(PT#7S;7Vg_(AU#Mb6IE.[[6cXK\KB6Wg5S2]5
&5dKWCT2<KEAP\f<1)TJ[a93(]d]NOLPZATO:>Ad5X=<<_TSEdTH_d5MC&Pg?eE3
=2/:Q.+K48.G0)2\(P@dPgc6L))f-A6b&;JU2F;5A1]aBb^3A@MU66.cBJSH+NcC
/M?8f@bL2Z\Ye72EDSO(L4^J@1N4KXW+,4:GXfc-+/=XX3NcQ@R>dCC;S2B)7CBT
88ZZ>_0;.F=0V0\;\.]ZA&e/,3]A:[<X:N?IISTD);L^_XBGdHN9-<KA#4K>N_d3
I)e2?Db[O4gd4KC_NQS3T/)9O-a,D),M-+DfW:4Z\O6<17\]VA8B:QW)3cN7bSBC
E\4dFfTf\\?F4:8OB+P-eA8</1SBCMWE<89<9G2)P1eGFYY<XFYgI<@0)[Z4G>UN
RcTC_O+6Q36RO)eI8EX(gQ8S86ac^+?VfJD?aG\N6T[Y=@0OQ)OaN(ZAI5ff^W4\
+X48=TLM<dXf-#5S@bbZ-B0(;K[CS[ETFH1P[&g@DFA?9FA>P;#L&NA?ML&&(VZ/
Z#SBYIYNfQ+7NNHS21bX0f,H)?\,<8ZM]91N9A=LFSNCe;>1XcVZYdZVBI38RFE3
RONAWb#@>2\OD@QC9DU[Fe6.G7NLG7(HZ\@_XZ(-RM]3BTZLOHSacURQRE.1?I?W
ZZ^P01/^N&RBEHOP>G=GRXA^I34UL9ZJ@c3>-aT53Vc0A>aPO,.^75/_+([U/&E=
2TCI8U9O8,((98aYE>JT5/20[X240A]3CE[X,O9R>1KWadE]ccT)WA_9fWC.1-RY
AO1.bd6)5gA<MN?P33QT.S7L;L@0?_Aa#;=I_g\<Yba5EdSc<)Yc_3U(7FUfI0;e
bPSS550aeU2;O.Q,3V[&7eHO3L/;]?I2eD9CV.>fF<,(]?AY2b:BK0/S^L3UgNC1
Y@H@3UA^/AG1E5&<#JH]:QX(Pb]J.\.M(M;Y=SMb]H_&cZ[eNWW&-SEceZF1<AL/
&5A3DA@4?C:?0[:9\R?@B<A^^I\04GT2=UaF2Ud0[)?GXcW/F@b0#dfPK@3dZ>,Y
cDCMITE,>5HWF0Z]<)eY);a/\fCLI^JKV@ANAf1Gc-8/+7&Q(.c3HBH/5SZ_?<TS
578Jd,L2BZC95&<4)c8Y5XS0C>&YRNaNQUT[bfaJ/Q(O7c_2eT;f[?-DH&?P^Ua1
6c,?dD1@;)XeCU=4/bS1Tc2-U31V1X@683)]S[3B8>Xe[WMNfHRH(H<,ZZ]@=ZI<
IUJ>Ke80(LE8Z3QgZ+\@R_]M8;)db[D@J?.d.6^O?^dN2e0:7=@NDfe8^>V?WA:f
P](I4\\_ZZNI7-;#:FP?gYaUPY[IM<0H\DY#MHPXfQKMS2TSQJ,;Q2P@0><0BU6(
DbZP4f[KQ-N29WEC\TKVN>R43J9\E(18O+MAR23<WAQ>,=U.aaQaXFL,B+^/\Y_A
+I@1afNLM]cB:YJXO_K.+=<P9-\cZec8O;?Oe#LXaM>ceF49E\<aa#BH9#TX3AEF
NUO5/eE\a]^UYc2W[EDG.Y\=+5WO_TGKBQDQbVW+,UIFEL-^cA0&cT7Mgf(#755J
N?FD_.YWFdH4a_04Tfa<E>DE@??Cf(,c/V_AR,,LM0<VTBC(U_69N3K2W;Z:bPS9
_U46Va]VOG7__N&;Y^KYgD/?bP/JIX0Xa>Ig=#AT3cQZd0)^I3@3RaIdLQ[LK4BG
UM54=CN];9G7K3Ja[H1RBETa6\cB2<:?0?5K?fIP_CLf,+)1(Vb9I<W,Z+eSVU93
DVf,X@g0fK1a2&5aZ\4KGJa?/HFY/_e9NUJ@]eDFaP7cX,ISf>0S=b,C<C+>.S]M
aPZ;KXS_fb]=.TFbZO#KF&IZ0].JgbS^D,N.T.;D[<)+Ba+5D6eE>T4,H[XYMEQ(
.UaU5.^H&JHO,bW55PfDY.W>]]W#8;+#75dU7(-[_PET[Z8@E?>_UMGO[dN2Df7]
+-=.-G/4aVZ[PL)QC78X=^V&?#:D#KD5#?9Z_G+9Y;O1@1OLY7Z&+8P:L#DC+J:0
K=@,MQee.(=@a0fY3eFN0I(4O?A.-Afa>,F\[0+.Ag>Q\eQ0-U5LHd+Lc,#VHFO#
W:ZLD-+B2IEG2UNf?Z4YKK5&[f5&>F>f?@]c@/P85.PX]OZec>gM\H6B48/gG1<T
d-&>=.b#=20M(Ldb(ZK1;#-:[b=;,?N.dTSG8)A-G,T14AH_+aYLa40[Xcc@W_b@
>REZ-C8fAa-7JE+d&K&JOa/#AY2Q(WP=T;Ic.)<F8.A?_7>24&G=JO.#UEc:e&WU
ZK;,(X]F4IKV:(G#N.aL60=O2]2DN40WEJ&.T9(YG/1<9RU9C@cK(C?Eg5Q[JF.C
^fWUS1(<&R&R&@O7V2G8b@_/F7J9#<.Pe=)@]\eV.T5KUN12KfC4eSYL0:OF,V,@
^1,X>?BH,)2TRf5-NESQ?C5C,eX0&M92.d-cX.=;+f,[E7J.BI[/_EUbMMUP;>89
,7@#2^ND_7]KO)ETT);4]VS=8=(BC?6[f88&#8I&[?P56=N<2.;]/d._L#2QeAM6
9QX]eb)T1HZ,UVN8C>\O9B<=INT(+e22]V05LH#CW/=>d1Ec9a-5>I,Y8MX>=AW@
UQ@U&J+^gQ<9:XgX@U&P.7DY97OXY@Y3eBCI_V<(B;7d+gLY.)74&MK,2H@7;D.\
8bLE0AZ1A[&J;KF)2507H_CX7AG;](=X>MCM@]B&5ZRaD?,>Z8GM\OM7HADaDHQ1
&ea=OgGR+ga1]U+&Y>BLGCQ#3)9K[YV2CLfCg#aB9^ad&(\M_f\dABE2>f7.#^d^
bEA\CK=c.OARMM,\TT9=>LF#=CZ6[O<1@Q)YJ/R0-TVT?+f+[;.:4;\@DUPHX8FW
\D]7V.Rf3-U17MTO(@WAR:7XWTdgJLcHd?;PLgNDL-O;G3\PXUYV>6ULZZ7Y,9ac
=LS6]+WfN83S4BGgQG]SNP,^UF)TC>_>R3GYcXIK_\??g3]IGK]-_\31N,+6KQPJ
6614ZUYb[2gcY.Z>2Y3,.,O1\-0f9f)-Y<Pd]?WF^Q3G+FZg1_]/a6\AWHDB8G5&
8X3FKgb=@_F8T/@L4\:dQ1ZR]FXIZP5O2&[eA;Y&:)g:1KR&]8D9B3O/ZYeZ2<7@
dIU0I2d0c?e-F,6W4&6,0&6>CIYWMgNFbaLfL+632:_?O?)/<3E_V88>bU(APcb\
Ng1H?V2Rc7SE4f^U^N.(Q748I2285TOT3\3CV+T3L..,W#^VZ6<H.]/UF=3KJB8Q
cgE?/H7YJDaZG;?dE1O<-Q2()B0K&-bLaV9f[8E6]5NW2KVKaR1#[eX^\4?,J^M0
LAdZ\:.UaQ_\<;QUf>U#L:S7d+)BbW@?0=F5bA+NSM/a5_P@e<a#GCI4&FGX&cBC
9(ZN_#1LNgXH1B7]f:EaDH;:fB?D.[SMed^;[=faQFFS(I_/+\7=V9T@<_d92K?O
^eF#_f(;87X3Ra]<0^9A1=L5J>0^O]Y]FNK\/3DG/+<(_I#7]6d;8,N/OB66-Y7R
?P>0a52:S(<282Y9dX29\>4X-)1gOTKbUF(0YU7+=0840<D../1[4X0UBbeD,8(:
<g9+J6a8T7.?NS#ST8PN=g#T^=#]#=T_BI(E_I-(+4Ke@SHC>5@>T&^:;e00J)=M
\-J9PaZ_-+V40HL8?ZRa<f]J\UVW<2#)MYQ;TGQPTVA6KU.V]d=Xc]J)OQCS&UP(
GND/AcHBTa,)@]I5:/eP&0V=dY5MJD+WF^O30H7b<)XHKA]RP@P#DeY_##\H0\R\
DKgIN(1Z-VI/6DR_bgAa.CU<T[YP6Ed3:,];+^I-BBD_T-J.IZL[b_);;dF^P1@J
&-CgfX/AVG\;)d,6f]&HeJ#A@8RZ&^8\)=e#&27B8[@Y=8A0XA=g2@9CXIDHedFY
5\PK6#4;4(7,X:O^>K5aMPR>2OgPS<CG?MLU7L^9;]\S@U6.)Q^&H)HP.A^27HR;
0fP/K)L&,,?E[/D;JJRaQ<3KJ42&<C4@NI[Y^NVC_G^=IMeGBP&0JW738++PIL/.
(aaQ85J;d6:_e=<YIHI_BH-C&+WOCbY6N+\>S[6A2A1gRISF)/+=)N]?LSTZO8VK
UFaOG]Q]gCaPfe8a-[Y/1<(KF]SEDb\FS]7]AZ44Af[[Z9^Cg[;PfZQIA28&V#Wg
EX=(,,5(2[Ag)9&:aZP=+?BU@&-f7I[DT>?\SL6MO;gDIS^5K8ABB4S??+@^cMI:
M5.BUae,8bB5gAI?YC+8QZ+)]ECOG;TYNY;9E@+7SSF00.;^G,E#Le<\8L<IJ]:(
\\9/?3g#.[d^b))FR9d3&<2f/&BFQ):9F2\_0Z[TG2:dK1BQ?NPM:f4>X@[YT[WK
,@c;FadI,1.CgbFG@C5P2a47I1T7@UgUd)fF_=d2&B2Jd@=3Ua?U@<)@+PZ&Q.d?
_WS78\^f50_Y9^LJ]+&;8\7,df];9E8UbAMaQCBF0QfH(R+B6:<37bNC#+5C2a<_
BTT2#M92Z@.JMQ=?g=)M)]A#AETFV09FAg6&gHI.O[\02ZZA-+A2W@B#]^8/_5UN
]>9ZN73e00S14g1a0VLR.3?3\E0WHL1?W5+-FN@DfT;\5TYA4Zg2dN;2]#N4F?[4
3Y;eLJF?0Jd6LHOVf#GX>CZ>6NDH+_5/]d?_Hc>W66ZM\(CHY[>Sa&J=-Y_KDG;,
J<0bG@BfR[RF,7ZW0R-+=.DN#PZ8SG+OT#a97R.4gcPIAd7,MJb<GICLUgZf4ARQ
ZF9L0N?D<KTdF>cA22EX#1gYO7EL,QD-:cC,6#Ba2^<c_Kf^DE=V+,8A8aV<SA>+
G+94FTMcA\\A@XW+,NC84<+4K_e3)=)9KTAML/#fI1TS1a3dSZWIdSBE4[IgbG<W
U=?5<V3M+.?,Ma1V:?5d/dG:W)?7F7SVU2:H?IGHM^;aYE24?aJ[PdP:-2]VZf-#
dE?E?1DCfKcMM&,<LdK&_20Sd.=OR@)6.-U6DF9S[T38>#5?XP7+RP[3BR1bC.(=
-)UY&39XS]7ZY2[8cBZIYN=9MX?BV.#e@J@7#I#geZ9).FaL9/II>+-:NWQ6TL;(
bPOBc8dUAgH-)M@T_ZH0>(?I>EH7P<H4U[K/>:C-);=5BCFS]?@#:f5F?Q-Z_>(D
eB(UJ42)<D/e(BI_1U94G(DNJV2@I62>4PD-[3_JEdGF))8aHB9]C_._e?JG)#:b
J?G<5L:gB5E?c@bK>(KdR5?gQB[@R+F_,&9R<EQ(H2@:NC^<@?2J#M:gP<ad_b0X
aCY2:-#(;4MKV@b]&.K1g&#SK\3/V1]d/KGUL9>#@M1>YXMPF0?N]1eTPP8X,(Lf
Z4-^M17^TYDPLQbHU9O:,/RDSC\3d&EaSE<M)X3gE<53W_57gF&+1RJJ:8bX&F<W
6HE>E]S&X5FE8^Zb<#IA^^((EM>&\I(3WUT30>8X/\4,1\KgCgP6e^[-Q86bZF<A
3;5WbW:4=eDdX?=H^^1-(F574S3(K[.db0GXIb)6PL#](R06M/fabZ802\ATUb,0
d#+SY\X^U[RO7M)XWSJXd+L@A.[>&G)O2Ia^;U,;#BY\=A457NDYK#WJ3#RPcP8L
VFX^&e\JY#WI]X1fD#^:)=b&Y7ff/,ZE3,b6P+G7OGG9T=^/EFU4O4=;^-[@E^=_
=T1&4f7=/Ud0D^ce9>(GA5<DP512RC)MQQgff[f4=S_c@5CTE09FOW(Zg@)_I42I
@V6V021^S[1e0909WD54@J#/H8^5@C@RTeg\Q5=YLL01Y]=EF&9MP5I=9<FG+4A-
&X8\+FHBNP#N)K]D>c\D2IA:4PKIO(dS#V?)WA3Ff2KL]QKYAJ^90E\dc.BQd43F
&_O0DbF[Y,]>X[D5)W8/:Fa<e6)F9AP/B>b/F,;:ea#-?F-2bUbDeUSLb_@H)3Ub
Y3g6-1NbK1A^65=DHX7#YCFK@e[70&RFQR:0eW@b7gJU6^UXTH_aPC>bB,:PKRGL
W;\?@==A/+Hd#+U<d<=A(F04F&5(+3FH^]IL1P]a94OFH40OX4D05TVC9Ng2.d^:
5]E,2YSDFf0a6-(;/X+T[KdfA3&UP9GWf[d2#&K7;.R;A/.G1S_ZcS1@YeR/;fO@
W:5PQTQ4B9FEgVDH6<TD-f@@AT;+-1<N_,H6;gTQ?V6c-Ofa&R\OGb\BfZ.4DEU?
TQE&@_Lc;RT2V;N4C[0T.+#dU,E1@UT8B=EVb=A]:J4S5K6fVbMRN9HS\cF>;#K]
3P)Fg(_d4X;dCDeMD_)E7,c1#JNL0]_L[fa9X=HH[6.Qd<2.NCU&_f\MS2@(;7f]
aMGOIYT<R^H@d9_LVe&3Z\OV=1E<cX1=T/.bHWb]WQFNcUDG)0e4e_3c8Jb#f503
Z?1E?;@L4P4PLV#g)\BX_PQIBgFX,PgFfUIA@P=/-8c;DNef4QXN<HC5&Z2Y;c1:
?4Vd2NQ:A>KPVbD0]gSRYCQ&T;IMCd2egMe6Mc1E&7E=U-A5S-6:d[T)ZDe5B/<G
&&<PLV+G?/OLR8,Z(+7E64Cf#L^]FKV>O^c?YTf\]V)b1A6V7>GE^L7\[2EVUM0+
N+>M#I7@L7R(1eABgDa3G3HbD@b[EX9803Cdf;Z8[)A3GO7fHYBdXFc\WWVPBg@W
I-C)J8KWYA(O=4eOQCKVBR1QHLYF]FBW1Pa941gJI5+_MCCF=6^GVGaL[:UU9U./
c-#11B-J3V[6[fQ:/0@4\@6RU+7F6[(_9DK5+NPOI+KC1E2c>7/C8J:1)X)[)f]C
A+UcVB<Ye[YHLOKe(@R85R0]OKA674+f.F^I@)#C?S&/RC=CA54-(SC=5>SM8?MU
L^;[9J9YGTCZHZK&G3f88Z>:ICeCQ:+Sc<C<+B->HAeA(,,ODfMddgC-GXa3.X))
?4TM2E5G+3QJf9/L^-@2^8;^<-PMPK7D51=e+cGbSc_C-4/JK+51=PK.N?,C[I+M
=OJd_e/>gSD>cW#AZK57^f71<CD&==SPP=7?]_?P>:HKEC4KX<D3[d)B_\;FTZ@K
A,?JW-MQ_[V&+c+]KQC[cR1]5P)eSUE68RLR9GQNBBcNfTMe,Ac5I@PJO2Od#H/L
O>NCV=b7M<d2HJAgV(Q]-Hgg:,WPKR9TV<PdN\JAb&HY??eE&:83HeUS[C-(-&gR
(Gd?Q&f9QS0\LQ)_(R)^47XdQXQ-=E<_5W8KJf/XQg:NYP)8>\N/F),5PV.IZ1.J
[FG\,Mab(Wd&3B005;aHQQ7cO8)<0+:N4+.RK2Xe+#_=])(8S1^<HJ2IZH8+]?Ba
ed-.U_#FC0049^L;2#aS#+6P,3V8edJ@Uc9.NCGQ09T.C4T(cZN3/>CJ42YQ052c
SCH=A-Rg++UdaCYcZ^,/W25=X#c\-NTD8a)&gKQ?-a.B71H]UTHLFJLae&^HB>R1
dPb:0[6eA\8HXLMZAb6^agNc41PI6,-Y>;KG_2;YCI,[ZJfR8R6Xg_?_M+B@b;M;
B&=;BS31#.,UM;)Q;aKVHeSb/YE+V=7gb@P\Y+f0HDX\QeQd_T@W+.#G@WM)DaYW
9<&g4RRcPGCQ0KAS]9<6V0789D>359APHIeX9D&+a;8]/=PUD7X#XVS?L\#L8Y/F
OC]Y8V+8J+H2fKKWY8?PBL0Z#0MQW]_LG/\GRfYMSNF#Gf(ASL;6de3M8BF^1DRD
<#76[A9a#:UZaG\gP66ReG?&60Z\UD3)/d@b?<QHNQa1aEAg8\&8Nb68M0W=32==
ZJ&b/Y0>NX]Ced(C2RA;UbJ2?JfH158c6XdQ.BI5)GAaOc8N[(.UJe\fUB+LaGVU
M3Q019B)g>g,8\INWP08HIMYd]H0T@e+ebF2=IPD]DHE;Vae<GI2)D4LM5FK67FB
Ca?LZDR(LX./LI&4XHXQ1eVS[Ze^FC0]6;F05V=#9cb2Q_f2QaG63]6[:b3MI</3
5gXN\[4eR5OGO0\FgbfJbLMdD,FI3>(3_/.FaI@GgNOF+XB>K8P1)-^Nc;58TW&f
SX__(Peg;VZ<=)KcT+)ba(Y.QP8>+N#J;e8]XO;O&d#TIKfDZ>)0?Ce;XZPcc14@
>J?#2RZ<^6+>C\7B-[8NAAM-W8<ge[fD://?-/+XE:0WQ3<9L1c;)d1V53AMbc=X
=L=P9,#5K[0gab0&fP+\#bGcE7O0c#/L:M_ENT<dDXSV9E;\)-/D>g8Y<@+2g0T3
0XVF-@X?X109fN]@+AFAX+V0IgN/Q+3N4-F#5\bL]8bRJ55,/UZTdU>T.FG^GRK6
B>+J4bK6ZBW0<3b@R0YPS9C.]I[;gBU2g86BRZNb5+R8]C+F):K;PN;CW.R;<?g8
9;V4-QBA2EdZF6W:TBXSQ)+VFI>1K1@T64,1QF_Gb+;G)_EDB\S)]S_9(g6gHaDB
<Y?L529P2/Mc><3E9fPEe&?EF37(QF-):Wc+C/5#&A;\Mf4caEJg>YOd-X0O8W=a
72\X]Z_CMIAWg;H.-TDHJ14G#UW/H3IfO=b1.>:WKLL:6#YI6.QX-_]?^WdKGebH
PV[:@A^T?5;BA7]g3/=&\P4L4#1S^Sd2XLVV^HZ9&Nd\:e9CDM+PGZH3EO6S=X?A
[5]HdaGAJ#XDD;^RaJGVJ9fe/JVPG)<d+U/_]eH/.7XB^fYAZd<b7RLbNQg]1S+1
K:B90V;2JgL@]B4CX-#:^bHL^e]6bg)<PWDc#EVEbHLMC;969K[fZ(-ec1-_G@Ne
VH;cF59Uab+AN;M03M27CO/=f&:]PQ@8gJ0CL2??M5O3WDG/L71?IK:MdS.[,d]9
367[&RE-;.Z>)HM^QK<g#^Q,97JZR7b=8E:=N+QC2Ie<>QS/(8c5OSgdJ#URYMg7
cFgGd\;]:DV1,[:LVMW/8GINL?LOWHLFc\+g:1]^^Rc^dd^)ZcGKaGNC;@\CGLaJ
[W\fg>O[E<ZA1;YOgLWY_T)YcBDGSd28E=]?dCZ.RSO+=;<-?Y[TJSA-X9^E1L^J
]QZPL+JI.5KWOF@#N(1UP\OAD]<CMS]]K:I/O,fD[ee-@?-.T/5]6QF8UG]EaKVL
P,<FT2DVKF3V^MIF[.=N3-2+.AU^;@97.1C0;N&UW1N@de)RX#);gUD,6DB#SRS]
>U^(/R&QWTbfEW>GO:V3A&)HAd>^+<2g7=/_D#[bfYXQ)>4>b<LE7^6]LNaf@POB
>X-8MQ/#cA-@H#7KebeCSKE;UEI9C93g]f_UcD/cbVY+V_9I(4H_[FY=92=L8\S=
4bSWVC0Le?/D^Ga;;\EbObYYSAIWS]059>-7c;:5W\0]g[:V==CI/\<+a(\+233N
BK7GJ@dD0YM@RQY1)&M\HC1aMMYX8J-W>)f]aO^8F4563Tbd=05S+H(<d3#BaLI&
]VDYc?e/A>C,=BTNJ(16.PaD:)^7K(a;T??ZEXbCRSf1YeK\:55ZR>#\.b.NR^F8
I9&PK2Ve^>Zb1&#Z,F]8;O9N0\W1fdY+cBE(+\_F:0N:GHc:,Pc_0DUD3(&46aVe
Pb.VNb1[\N<g3_A/..1F<?>Xb[88._T7)5GH&[)\2YG?c[ALLaUM1BFH0_D]FgJe
_KL@\ZM+F9U_KV6&1TBRWg5[g1SdXV90aKE5>LFL=b9@[5P[aI2A<ULR)#4=1#U+
70>S1V;eRVO,>XAP5.SI_94W8L=7J?>U.?;O#Z1TS[BGV)/6gH>dcP?L:HPMS)d_
[<?>=J@2L)<d:b&P,SBEBW7L,dL;B(_EOPaEL8fIHJR=]W,U_=_[AIfd^R-a^T3O
1LE=<#A>B:?0^0Fg1+)/Y=FP0eEB-MO5e7NMAf?:9+QME]XL>baFeDCU-\J>F<?,
_Mg1)]g42d[#^)HR6T5F2O]eG2]=aFd7+TSYb\AY5SD3Q:QKTF[P33eID?6+),f>
J?T>1_@];9.)fIS04g@T67eIQ#M0#<D1W+[\PH7RHA:2b@I1_IRUS#M.g#c=[A)?
<[XBS<1B(GQ0J9-Q;Z5gGO4CB24NAO=M/JccS/VOPO6]/8IQ?]-NgS?&???;J)>)
a?7)?BJX(TDg2?^;+Bd1c-LJJYEN\H3T7?]4M3;Sfc?1Xe04>Sf;42eccMBfcYec
4df0C728g46+K_8^\AF2YF=E[JcA;VD1-d1^4,L^EJC^Y;1>Hca1=:&-+;2d:aK;
W-C;Q@=NXZ?H?)4HF7c65#NG_HV4O#>X647_VCbJgFII1V]44&[<.^T6-_?05PPg
b:).>>)HU@J5\B5CF>VG?dHA7,X-QR#F7OMCPN,(M.#M_@HfX=9FcX(^;;aK(W;H
<NUI)^^75,_,9_?M^8g;(93eeI>_(?HT.5=.5@=](.3Y#SE<Pa#Vac328(Lc]XG1
Z4C_?<Ad:QPE[Y,)I,L8GZf><&VR^T@PZd>dA-#JCc2_IgY[#:NOC\dL7RNe+Sfc
MLAfD@ED@KB?5@.XS_]0#+.fQA0>6g4(N+IV2eMSd3f1?^6YcGVOa[_eK(fRTa)C
EGSS8aH?8M5X28N3:>WgO4DJd..T(AX7(Q&fK_9Q(3)S>8BQ,6_e.&e;S6X^db?B
F_\J,,1J9+9S[K@K\>-I8<<[J[;Q@2g=MJ,]Xd^OcgDEA-W^&?\-DBT;-32M(d0&
fU>7/f02^eS8@E])=C:g+f)Pd:1aPC>[:L2M8#>CPZEAcW.0G=NecCIT,<[VbQG6
1XO-RV4[\T-PZA<T?.&>GF2Ge9(f?@(R:81b(6J2]M,M+gA[XNQ:0V7^PJ;-/.>S
M)?)^=3f6^676L0^d9;8@LS6;e)UV)XVL5?8ZY,][W_I,:.UMYSRNccCg_4f&HO2
:.a),:I]((?WD^D-4]MF)0g4)e)EA850)3Y[&NfIg+a.C[7]=WR?844adDf)CZT?
YfO&?_06(-RbLWA]f@Af69_(B]>f-A-]\:K]-+MJS&L<ACJ(R2I&&QcZ>2G?V1UW
O>33gSYW@)PJb_+fY,^#f79Wc22NY?9d,)0&A0CVE3T+P@OKU_d-E\6g(C9D31V[
cN_^e4Za[35?HKJD&]395HR<dJe\3<03GKN]eZX:d6(/P\+EJ^EKW32H2[eP>7bZ
HBb8NBfN<?48LIJ@@6C)#-#.bAOWW\.[++)A2f^W_BA-FTWc.:>Z7YV\#U]b5=S2
-KI8a\a25d(;U^D@.>&1VAdeT.?9f>XJ]G\GS8QJWFZ=NI\Cc8GDXF_6-e4MdLa3
G+/FHeM&SX2OQMd9_Q1W+/FF1VH8fMK0gD7e8M(VTTOT>b5:Y,Y#?9.?4g_\14F6
P7feN&c31e?X_NUM0WT9MA:XA#WR0]VQ7@ND8c>V8fJR@0:_9Rea-3_\;4+V6F=&
KYN()Qg_XP#7^VT1>(.+CL0e@=O;2BbL)R-5:SEE&:C.6MUZ3>&W@A>1aJW5fJ9\
6B@c6)6A4cOXa[KO:7BW;a(5gG:QCJ&-ELPXP)8/8fFE/<IVP5+(W<eJ@E\c/ReO
JTL-65OT36W]FQ(JEE?Ke;dO+UJfU_dKAB9<.cFWJ^BA03gRe56(D3L&UCZ-(?31
:YQJQ.IJ@RcY2</fPeIZcINe4)DSB2+XN7-@@H2QB7<(0<?e3L+TSfTL#2b_7\e]
ZU,6U@1?7BCZF72=8S1e^+6#XDPJF^fdY]NMP8T\AAgXJ-?I&:e@NVP\X/)a1G9+
7GK8bQ_/67[(^9W>Z_BOC?9EL+F-#<_(DKI9SaL#e=3aX6(N13PA+[:aN#-J<H/C
8V):0SUbG3L7/#GbNV;EdV.+6E:)OHf\+gR8A^QI>.DS[69RXb[#^RLbb#3a7Y>+
?R3IO=_JWERE6d#bPB6.Y[FID@;_709_#<aX;Zb/-S6>=0UF@=XNRdO;]+?d)<b:
W;43Y:K^f]N:/+>0ZWO[A+=D^ScJ]+P(S[KZ_d9dIa\6PC<_VdM7QGQ4VIdHQ,[U
>MCMGC[V=7H)^Z3QG9A\Je,991L=a-DEa61Md.7BK\SO2Q->\LTPO\<Ca&NYUf_g
HAMZ<[B(8XM,X5W_cVG+_\+@]J@(P8eKDa5>4:R8M(ET3:<^U<RZa>03_:/\Q+=J
P55;,eRT0YP5@UV.5W1(PUc3g^;4FB7aW6]8(D1&JKH>EV0cC+b-XM1^JA<[TA[3
KG-TRU#A_N&0Y^NJ85)@A8>F83e5]7+4\]b\81cfFTK-L>\>+@0bAH<OERJ3\>]+
?2F(9G/D7O&f\HF&IMUEcb@BJFa4_7^MT=@-FW][?F;,5&>1L@D+:?=<O[06_V+&
QAG.2-#__Ba<_MK@ZPIbHH.@S\1JbXVUR3M<U+9VEW:[RbGBQdVA4U#(J#^+Y\0f
OQ_;;MU@=4Ab/9B-MTA\c^OQAZXNPTZ,2?fPQNe&PIJ-/G<]^\9]P<(H;FQQD,3e
IJRLE1@D<)9aPMPG=\3a4,+KaXPMO3RAUI^A1O/X=g<XU[>AbOf2P?+GP9]DEOM.
,6@O)TR9PL1#Ob&T:EgG->&VRaf=E6.H6.\S)4aWR-V>PY0K_TZU13S74f>,C?fS
,.KTZ2K4UNF=#K]SZ:aLV&cd6<;GBMBN@42EK:)e,@&IgH:<E2R1N-=/&D?>LOBA
3F?0DQ02)Xc[49N(-2#/U:MY>-(WUd3:^N^D6#1J.#N=YDLRI[3U\6VPcNB)IGRX
9:&>3&Bf11b0]/42D9BJ^4)Fd;#TP4e2fVMcRQ=(S?RCAA;WbeaG.FJDK=2Ge&>V
[A\3KVFJC4+.a^\fSXMGcM)#46\6W6cX[,da#?,feA[NU28=+cKR7+U@];_3.:0.
ZL6<-E.X,==#T&MS6?KgH8&_/S/,GV[8U,_M1R<<;#dg;@<Z/fb\V07W8K5/+d_S
J6Df.+=GTgQNDb=eJ3fQEL+5VRCf[I-8+J9=LHfL><5KAQV943^SP80=cDf;#gL[
\Q;+UL,J?CQCeLJETUFV_[2XA#)@)P^TZ?/8.ECDV[T]LX>=TYZ5D,>=WRbQN]7H
=3[BO-KQA:LeBC;=Z#5V,&D<ead4CJS@E4P?562X)Ia2cFeT=X+O+G2Z.EVCWX0T
ZY^/=EUWTUcUU^VX)HaM\M7B^R0KE<HEegZQX-T3DUD6(5KV1X5-P(QYJS\&XEH4
T^&Dc,^K>(;P+SSTX8YeSFLP&5,D.^KUFcD<_>DE=>W3C[:[c+G^4HC]04QTZV^)
<fI^ZS3D\Z3G<7I06.>]RKVd6@GF3gEG=dA_?A7cQ8/I3:VWfXfOU<_8QLV@MBB4
:Sf&DLefH&SMF6d9_g,c)ba[Ae\AS2LY6Ic>,)<HGJ:ZF>@NQ>YV_294Lf8BL5Rg
;VT]&GFZ&-1(E/>/K];-fc&TDACC8,N>QM16ggRXX&-M;.b^_?aM[1Y9E:(87EE^
ZFHH[^.V5gKISRe]OL7+EL]H[^[BYK;8=8Rb,P(6F6Ucb8,M6J=3XR[@9ZN/YfN=
T>a>G)&8Y6ZLB^F7&..<.V2KLR>f7,D:X)+ZJ0LZa_Ja(>Z,b/aPDZB+)fN_ACH8
F^[TRg+NB1f+5eLKZ+FE\+NW4Z0:13<)^C6,C;PBOS7M.14JZ#EFQA_TFRF-&Hb^
-Cda2N9VVMI42e^c5R0-@F__DC+M?_5/5\[)\dTSJ7fT70AG[f\A;KICUe<8:55W
bJ.,2P[Z((:)@L]Y060V[(cU+M:;7)IK>bXf\c>P9A#YH-:aJ8IL#>aD5/fbRWU7
0+YR&ICDf67D[D4G#bF7/_b>L>8M&E]U[Oa&CF]e&Ff>#3N6a-cS=aEF8Db=[2TX
6Kg_LZ-TFUI;@G7,+@_a3XZ_5GYCMILX8/b9&3,QE))4O6PTCeWD(B[I]6S>HY&1
HWVYHeSgdW/Y@O37]\CM(=GJL:Y5bO3D<9#?gL.(L=T<NVO5JC896R&FFX(CPJ&?
7cZW51e]G9DE9FD3PD-fGH9.S#<6d1d<a3g-ZRG[-4;KC+<?a:g\ZNGX&6&^-E6E
H8aB+/)&(=Hb<(?4^B,O=NDb/I::Ga1R]9=<#YV?BMMfIMRMd]>2C?OB)D^^3#(Q
;<V>HN8#c(Jc=2aWMS8N6&^JDEFU5F9)=OH(9Y5N^=AY^J4+UQfL?]3Me=7dcZ)3
PT>M85E2HFN[RMI/_S\D;4C29^0CEP;U<ZREHJ@8+<DGLP9b,<HXJ[f>RZa),?:2
B.TIKQ->::#/eC<KgEEQKJK-]>8/?DIH-+)I;R+(O:AF/4&=7gZdTMA=;.E^]I:S
0?L]TZfA_7.1Y-UQ[g&5;HWV5b<?UXJ/QKH)d(B3=D<3ERe0PT]124]?3&0N\AGd
]\^]5[V;dT#1)YTLWO83b[YW^J>VHUKVU_\\S#Z@R-fX\)JJ,1EN/T[L;AQRG]c#
0FdfN]G1)feXa(UK?06D,#1<HAV74JR-67B9^B_J<JdNF,@0S\6W)^ZZ.:eeEbKZ
^b@37OCMT:GW(8L_V+-DcNHcaH\_]b>>ZS:EaHZ7I&6HFc2<FW,U#T,\T0=T2T@P
JH\F#7[JZ9=.7a+@ZK2f1EU)I@-]a(ZXWPA[FIM7.]MH]+ObWW7,[+FS<B8/5]&V
O+>-2H-+2KKO9\Z_WQ>3@<076.5d?V?fEEPSbaD,J\2gg]=ReVQ3/C_dXCYf9WUV
<;6@A6NT&&U;;/V+@<OHacZ>@C.10H.AO#;U8eXgV88F(2=KQ0O7.+)a]2U82U&;
MgT>CgH5#-E71MZQ:eP,g5Mec=@84-AST#VX672#I6E1N+2QJE2V(\V34R+8&5HJ
716\@BJJ9QH2S3Q,b#+<FUHJRJ,RP()H-ALR22L5K-]09D0@bQ(MFT.VUgT+ZN6S
)2C[@>+URM5<\U^5SJSKF]WXN(6\6N+<>g/FE0??adH9g?UBK?ZB<fB0IcYS#^(#
8/@;Hg9Q6EXaI3CTa]2+4DNgF2<.&aXc@<aQN0E]L#/bDV@ESb&Z>(_gVPU8=;Tc
BfD-MF\KeS-eT):ZPXa)eMc#MCTF^1d42TTK^:3P,R.Z+,PZ>?-OM9a.2eM/e<@4
^5e-DaFF3N0g)\1a6@#E^>2TUdbL2@c>a1_0GJUF1G]=B.),>R3b0..@M7LFdLEM
d/3T(;(^1;d>\S1:A=&P/]U6+U\ad1#-]U66P^?NG4>68G,,G@e^T#2B[S^I\Z3\
YC(YPR\NL:8e:^M,VT,Z.gH9B25+5K.+5W,[FOgbVZ+aD7H7YB?a:MNS?@;(WQ4)
cHAA#U^^f0.+W?2Rfd;dG(Q>R(=bPEId\D4MWEf=7ACT-#\:e5DU8;?=G+U>.0a?
6?ae^/>;E[)=E,c1aDbXWfI[M1]gR&eH>=F)-RI8[4NSMM(INE7@VS?S];(fJV1A
_(66)<]/2;DQ?WZ]4M+/Lg1Q1.>L&Ag1_8OcO)@F_A;F^d5cL#BX?U/)2+F,X>JE
NGTAUU>8dT7&]Wb(4),04_EGB?cf\[QfR]I16LR]@N_Q)W9A1Q]L84H6J/@8F:<F
ZA7IBeS_4daeKAf-HaQK2;K4:4fB-IGN0M74GZ1].)64V[gRAG8VE)/?@>GMPJT+
X@N1b3JZZ8-J31RW5?,3T=K7<527C:=J370BS\Vc/X/6dAfKJ\#]a9LHEZfGd,T5
gI9??+;@.\Y+;5@3_3K(ZZ?J7<@J_E1AOCXRQ4S]fDKNfZKeSe6:P&f&Y)PFeKOG
I^6\>MaQVY6@8Z7DZd4c\2eAJJ,=3+WKQB8Z\(S+:L+R=PL+f)]<BT;a;KQ.C[_Q
@TY-Z#a6#]aZJ=\BWX8W4[3;JKgXa,V4K?=7eSQ+LdRV-&g]K[^^b#OJYF.=3dRL
Pbd7AN8^ccHe9J(g4-,@>YK.6C2>OX)TLX7#IM5KIK_@]J,QfO5)U14YJ2WNE@73
f7e_f#N5R)_[B)5BSB2<QM)X)4@#:0I+IHJV3SZIK;W7a,+16OcG+e^fQF4K(T?9
1Tde,R(Qb=:,d=7^AP6KMR:<+eV(fP(>(NVT4MUVe,:+2XNJS/1[5Y70>;K0K/V@
eXX><7M]_>VCT_(&8+aAZgP?78I)6(^N[]&K=C29#;_d^f&+])C557]I0D[QA@+B
0Lg9)K1f7KNE-M#.UD:,2B+N:KNM33dDaP/gST/fZJ5<g?\797IB1@OCLcI@dg&Z
QGVf>:8092=D0bU(O&:YA,+<e-f(M</Yd/FOD:Qe,9-S@&fgJc\U1EgH-HD2.H3;
(<XICe&VJD;=LR@[C0QGcMR[D<B;79V74I_1c&5#N;^XRc[+KM,<>1<_b.9Q<9fa
R)O)#5AP[bV\#D;P1+1N\RBbE8MYb,,P3V\^=^>+##8fUI>[INXg:f^P7OV,34C4
B:HX9GXC[[bMNCW>9MaA:</_c@Y:I,&1?B9eE#84[2b<Xe+PdEE>@]O9RVQY-:5A
QU<DCI6eSMA\:VW]dIN@PU[ZA<)9C8Q0KZ]X76E7\EW,M1@81QBM=6UW45Z8=#4C
,]@A7)94RU_g0M=F;V1)1X17MGH.J1Yf1Ve_)J^202a;30E^]8P[AdS&DC^;d(I=
95dDA\YYbXZd5eXA9G?[_NKQd9b0Fc_#0YX^UbTVT=@_>^?5\A#V8ZTJ+K0>@.RF
cf3IaIYG_+fVR@dR@a-4cb5(BBa30<P[HD?:D)a?QG5V/6HU.235>C5JD=J-+I73
@3eQ.#&-W^Tg.U/2+;6Mg[bP5CBI#H6?/ZHg3OC-/<gYZ(QZ@d3,^0RW#0cc9R,)
c,,Jd;-0&])182T8eU5dK5<+:XB[e;WHYBMd3VB#3IY)&X]+2X9d-IbBEW7KXJ5Z
-(YcQ-+--7f0=J#LW6F5[W)>O<_eRc71,0bOTRBQ[bT<,>TUE\P<-5eC@L8L-Q@Q
6RQ;8.Q2Tcg_7JI[eV,e9O,>^0CIXZb[GE^a/Y?_XcD//\HM56[>/Z1<A78Gef2O
.I16Z&@aa@]6D75Y?)OYGGY^^.^<:6O[eI?MOa.;&=M/03CaN#1IC37B)E+T^?fJ
TN^TJWe#?LF@VR<.<Y]C3^52C&B\-YJ5TYcQ04V37OC>bFgd?1>Z@?CE+P<X=;U;
K_N#STX1/54g:ADHe\5Y3V.N&K&5FIC&I)+3GM0:eI-PF_dTa)/BI[2X&0ZZfbXb
856H\JDDX(?S7=^37.__&da:8)[ge>#AADNDM[5.eS6STU6gJS]4XP(BL;\VQR^a
74<,geebaPcOM+\QfST]9?[>FYA@)O8de6De).Og(CDCJf?+OR7+M=dNB,0A</9M
Z7-ZK:,)5BU<7LGd>6X/bP#A5[ITIb+=FXQ#[VOVAe+Tc9VK[C31L,.5;C9Qd+Ee
#ScF+:6eFDX3O4..FA4f:Lb37(BSYKH+SJI]T+)MS1?L0I=<;g_^/:\9W5OP1^:W
Wf:<.Q?M^JNHO0<e>,@@4)^bK9FVCV7WK6&?^e.0e:&6_S,Hb#PHQ,+SE?Q/?RI6
JA4)=cRdf?D&&aW=NgZae,A#E&EAFYOaH02LLK>:(C#2I@@D1;\P-4+gRT-L];/_
PPeY1N:Z.E+gb]W_@01QX7TY[/.A]cPCU-d#I?)]=W-MKd&P)adD?edA(g6C-[Sf
5<f4\S/2-4@A+_PA4&<WC2CeFQBgfQQG6(TVa)M8W[RH1M9-;fa(]X^E(Zd8W63M
3N>-^ZX/6=f]_V5MJgc@19,fXG5@&Ne2R2ER1BXZWTM4>If86ETeEE,dM7,YP]S[
O2d9^ec=8X^MO.)gFG47&c\0SB=F4a&FS8)U5+YE53H),&=>7dT4V,[QDF4gX6P3
Y#9Pb,#4BTcd(4?EFP)Y#g/10-=;(eR_D.0b<:CTI00#C2F(:+M0&/4:Tf/GfK\5
&>888MW+LP/\Z5eO[^7DFTI1;,Q?)H_-N\dR+Q6/S[CNc9W,\K))\eWV(A(Q4b0U
YdD)=^#FG5HJ?CdIYfg&_eX<&=QfR^2IL>bGd\T:ZOa_c+=,DR89LSgAS97&KWaW
DB@&MF_b;[XS<]\1a)g@R+P=.J_F=SeDaY:+.8;T=/QHQLB9M7&eN65-Tf2dZ@&]
dZOPC<:WUBDcC_WD>WO#F[8#XN5ZC[KbY-=&4aWW?dGVS:L[T]@bgb9\L_01B?)R
-N9,Qe:+D?YG6<c>5U5G9EY?UB(EJ@_1YJZ4A.I<)^YEb^\#W=</-(f1(D2LD9?Q
.]\]&(9&SDT5Y[JdA02A>L2CUPZN582YeX3f0(Z,-8YXZe)F,I61,^XRH7G.>dE?
Y:+FT+(2I?PC\J#UE>GRB8gJND:>Y<ZacE#Y?:)F#WD(c^IF7(Hb>.+WUc2(#d5Y
FcbD2>5HVXKOR0)[W5cSSafd8(ZL6abDZcZ48K;5H3>6X)+Q7A1]LQ/:P):(,&Wf
GOaU?W=_]H5BR&FcGM+Ye0P9#SIP.KM]4C.924P]1d^KfR^[^6<9)L;dZ\F)(=8D
La&NWY8bH(T;We5_S[02f4KC?3S3aB@I\GZV]Kd,;+#0.911GUP7J>0)Zfg_Ff]g
H&PDT#-1K<5<YZ@;F,59\L#a:@T,]T[#0PObI&]_aCY-XLW00S,E5.6\BFbFIe0]
P(->#e+ccAPTQ(/^H^.EWC)\eAT.ZY5IQ:,VMY7<dX#O//PRA7HIe;EGLHBV353V
I#,DSK5ag2+HP4fcc6N_N4ILY;aJ/+L91)T145/YN4\TMfE.gZ(#4_&U<O^Y\e?H
fdCgBA>#6Fcf&09BPQ.:\=9T7^-I(2Y1]3A=#AJ)Qf4;00\#P^U?.XA?PT:_)KV4
LPe:Ff2?7cKGg^UY@ZN.DMa27+A5L2=/F57#CeAUO\-\E]LcRZa[CLRee20CY.9;
=CTDbIeA>-^[4E;^7R>c4P;(-IU1G];W,eTYW79#d:11Oe83YHce_EXag3/U-NRB
L&JFIRFc-_<Y0Ne?WOb0PSdC\0,](2/KY]3d]?8W,dXQGeZK9,_5\0VTD1Ze^YgJ
Wg+EZEYFU5H#WIRB1R1N/Qc6FE57RRg.R5.HCSJRS?H@IbFD,?81.fU[<9fSS?QK
\10;H@e+\E531WdWF]K,6f+=-W[Eee@P6VMA[;?X;#AC^,&;g-FG?P1--=>E[/(@
]TV^C;#AS=C<ff^KTU,\DIa7,Y/Db&C,RKB-RG/EQ\6C_B,bLEJfVM0(bI]QBG8Z
CGND(g1D_+/.G4Ndc>FGAUF(H/O^:8d^1G7K1@#8:0,TV2^L<01\B-dgE=HP[:B.
,X4YcaNB:N,[GN3N9/AUXYC#@0.C@0BFQ\YZNFOef=RZg)UL8a[1[e;/>7.7=BM7
ZIX1\XDYcW>,3F;N>F0Wd:UXIBaf6:,Z@5G1DX_:He)DYaQDcAS[S9ZM?GLFb6C^
8UNYR<.Y5T)<62b9I].Y>ZU&AGH9YQP)#<86W/NJ]057<1\ED+b50Z-;-:aX-d@>
gCF,+MCKGJ762RXZAB,c?Qc/SgEK4=GfgLd+&gb>GIBD3@E:4GAW6;#D4Ma02(Ac
&AL[=[-T0WU<aV.RXXadBf06dXU00?M)g)c:N5cQKPW?VZ;a@@D<NCB(9L762L25
GM=7,P#L=-^\C#>(?YY8E7#BMJA4c6Z=Kg^?O9P.7C)TNZ\SNO(C&M5_VP::&^.>
A>VCU,X@?SHVORRB1BXCHYA8(>[Z.#JVH#3cOD]Q7-?2DRP[KBC[@=2?F<fRfdWC
SAaX#51R)R3PV18BPJ\JfI6(J?c#c?;#[6>AN^,F46:>=bceH&Z67=>ZLVO++BV?
_]E3eM9(6X;&6+C[Y^71-F>,DK0G2aO=W4g]ZD91&dUW]5RMeYdc:3QUP?ZZeM6J
\N+\<BEO^[WE?<\?YO]ED&<TfPBY+[5(PRg#g8ZS3Q2Q4?FW40IABJAXc[cVQa+W
VQ/U5[U6Ue0K,&5VYLM:P=d1097e&S\W=YgUKLHO\[;C9LLQ@6RGONE/c98FMC3E
N3DIU]3@()X6>.GXT<7,Og,S]D3+96C_:YPM8KE0-X(S7^XJQ)bJ+#P7[9TD;U2>
L(ZRdF;b64H>XYT_9Z6AXTXf#50ML[gA==GYI,8K.URH@N_6D5G2E8>EZ8P6dCO]
?6RWQAWS;&.[ga.D1.4</e+G0W:/d<d2T>S\.MDO?3;/8\WP.;P8X@JYCSHC5;T\
+c.LK//bV/(-IbL_f:,\DH#df7+/&B+;6d_0f7J?fSK)H#3CbJ+/D):-E2&?N:3\
J(d+YU/f0be[12.9E:8Ia=56L(CLb.+QL7Fe,a^2YC-YU&X>EeUG3e-?V,O@YHO5
V:HCP26++M+&Eda#7F2BX=7,)GN^9.)36=bQ,AeUX6d^GZe7\,71;2XFF9YZd:b.
TP;Z5,d3U:CIH3bM,\(Jg5d[=QNM.)L]c.=\TF2/MF,X6fg\C<D@JZ)/YW22J@f+
#A2M>7J=TVKK(Sd,[LaZLFa&?H#TG#C98UZ1]c4^E8#.+24I>H<e_RQa1WOIC5_C
VaL3=15N-X@=R6>b7Af(0ED1OdKYK?8eLZ(7GQF>91(P2&>dI+g<a)4Q:#7IOWGU
N^1g:6L+Ua#S>Dd.X&ZRUE,RdY1?=-T]UPR5?3:F6a#2V1E,WJ[WEY.MfGC=08,F
O2K?MaOPOA.J+=B,V8^/,6JW1,?1I.=K/cD+7ZX5(0T<a@9@)<1Vd_b=<E49OZ(&
&f5?B=I7#5)WSFTFW9;ZGR-;U[X+-ZTUPZGO8=>@^#(E\^O?ZXg)NL?<MS[2-ITK
.Tg(V;0aG>\a<5H]8@a1@+Qc&2^&WU:<Ca+Qd)F_>BIFCZ5B#2>[-SPTdPVX(F7K
EfII.c\Dg(\5S+E7-cAaLXO&(7XS-#fQ^XbYaC>PSP1NHd0-A,:+I<R6KAXUFH(/
aM;eZNbH0\VB_B+X&CI1149Y53J6V#g2Z7P#T]C78@eOM&@#McE,NRHcCJ:XR(D.
_a=Y]Cb.TZc_CU:N6G.PVAE<;>_A-D@gU/M^UY3]NMI?N.0D5WXa<eX2a7K/^JB6
YV6P53GWADX)Y\_:H]N+gg/:D:@>Y=-aDFOV,CW8WECNUa^PGWR<;dTU8YI<-JR2
?fXZ::Bc8.@V7d;2U561)N3X_:VbG_9V3J[>f0AO48Y]I(5;C:SCEddKT/dCf4C8
BTe<,A_W(4WKX@YQI:bK#PV43FZ^N+9Z:K;W&,T(YV8D6TBN@aJVdL,FA3\+fB>/
4J1bK]JgR_?[;Q^W8Y-HM1C0e+XR<JPeK8D7O6,10#G4egDCJS(<1T3474f#U3f:
b27[<TAZW[)@A?1EVWVd;.2S.LNC33Nc1@;f_E+3?GBBc+(C0.=/J#HT4<^0LbI^
9eJ;;,)2UX4W3:&+R(RF/PN@W5?R(NL8@TVP\6S+,(5IgKeTHQZ^1M/&,FJI/@0R
;-UV+(-O)VEDd6W-P?,=0J>-b?;7N0G-X5PQJH46:Ca-JKYN<FHR-[;3RM/EJ45&
&GVFX1SIbcF4Y?DXAF4/1W1C]Nb]BTG;#&_>4E<)e+:[_WWGBQ6;0Te6N@)afb7c
KQ[<<OB&f:TO:g8M75AF(7e)1=D.M/aRV-.GE-(XE2Ec\#W0XQA+-?+4c@JbgP0;
?E?]P]>09+P;dE\N<00\FdBHTZ#YHDgJeZ-=]0E9c(:[N_.c22CJ,5^;Z5@G1_Y.
\:31#<b8,LEVZaG<C=Yc@MFVD#C9c7b)(UHW@TCCL(,0=FZ/\NBXG5EE#5&-cT3Z
-VeZOD1(9Y41bJG#48<<RQ)\S[UP#]2P_R&)KXFe^S8.@WZK)4fFC2/F2gFLA8Nd
\P=<T33TTOUS/EF&d6+LIc<?NZC]ZZ)26LN)MUNLS(e7&EE@A4RX6cb:[S>D#K_@
Le<EHR=ad/a(FUGaB4RK:a7(#0>ET((30>0aW)B+HM)@J/10C&#UGd[dJ9KAN#4=
U<e0.M\dgd0,J:K<X8([XMMIR]HS[VAfaYXW#@Y2TA^>KPM_?^gG8L4H(C/J-@1;
9RP&69KI[/8]OR<86K:>/[0@\/<YL:c>R@RU<S8D^;;^VJ4@K(KQ]GNBUfBH9<TZ
.cR0?b+HLS&DRc[:UXd1<^HH0^0F9@?M4.,QY]DQP^X(0C1W3<cMM0(6E)e+<W0D
]U7a&.1Od41TdV.IeNbVS:P:&A;NZbH7_@ZYMQbOWF7A_K,Ob+T.>b]QZ^3a24V?
&@+?eZF3>-J>.ORB?IY[XKW_..?Z1JNfM8^QLU<6AI(=,I4>.V^>_7e61e,Bb><)
a>e^RB71VLeg]#T253GL#-S6AGIH^^N#QXgBX#dD;UfM>&Db)??gP2dccJ(5+T@N
-,[bE:EfdEPa7[MJO,<f+1@^>Q373^ZS0;?Ega99DF@BPIP0)MV;OO8PQ;GDFEG\
#I;3f?8IXH1069V[-)gHJ1bAHXQ\b&]3BE?+[(IR^PSa.WceG-66_fM\<E[;H>:e
[SM;NfW.3C:6cc^NE=+=Z7;^dX_/\dL(EU\SA_fM/eI9b<./O4[H;_-)T?.dAWeI
4JCH]_6\BOF1ZBLH-cB2I&TO./:1S8gW^4<YP<Xf[.-1>BBCF6(O=J]8SVaI6d0P
Fg.e4)M7^8a=b_?bWI16-7S+P^A/fWQ(Z/<?0NJQ#:C_/NZg5M3:0&aJ1CLBJd@K
5Ud_/=V48CB_,aA]R3TM@b+AD56#R,.bXO<ILW]O7a(VA4(.g?c25?eIaS,]FMHD
[8D.1:D4PXfB>BeAU.#ZI,R73-+a&62[I)-I-#dX?e#1FcB+Z@Cc-;#L_(BSYLe<
H:]HffQ3[g?,X^Qcgca0VA^/NV@JcgaF/5&8MN86g(Q3]f\&J7DW0#C3JOCO(gKY
@dE.&6c#A^Cc1^9-DC/L;]K)V.O=<ZFW)=&0?Dd^D).C2@^EJVIX<.8V[dda(H&O
3FD40S7_(&L\B3Q?/3Ae]2,bA)g8&26,NCAJG5CC7KQKUb_,f0-dWMW3,d0L.3IF
.Q<]FP]1eJ.^Q]ec_P.5_=C8cB1U>R1bU,)<#FQGWTE-e<TbG))P6aaAL5B\L?P,
dG^@VR?Za12)V[LLa&MdgX.Qd;NI3.P4:;/W.&0^+\IKZ=\TI9Lff3E8Uf>NYT0(
,fafAeR=0)RN;U#NG5KdC1?D9<9V,f^]c2+C)<]2\K/MfEL(1UH7^)G?0.7[;L8(
bE+LHQW[MA#\/:JIR#a:N[X\K5WW;/PG^YZ#[F=5ECc(P](:P\&:UV\X7)gXVgB#
ZA^7+9_X+P+g28\R[NDO+S.RL>BQd1NeK6.&,Yc&feB=[R[)Hg^-?D5;7BL)/(OE
UgM?NaV)&QFMIMYF,RONeI&^U^0G,3;)ca=f9CGYL4YX>c8+C1OW4F13HRNO)W-S
H2P9M-W]aJHg_22I&Z?<0(<b^c19QbaJ-ICE8f([b3b=&K/SMNOI#K3#^@]_^>CD
)E9A,]?=X?WP\444DYY5fKc2eA@O8Fd8BAGN3O().BNIJCXUDXPaP>aBc44+>FW-
RYaKSBXITSa69;[f8>(QXP-3aML.]e[/KT;1,2W;GJ2O]>OU6#T(.9^NBbURE4G7
NeT\BcM;8GeU6-Vb2\^DV#7TgDM2KM4/N=O.I<9.].R&V),K2<3LaA-?\V8:(da\
d1RWTEKDLLH#.:@gI,D_F-ceD&M2S8^6VN+gM?CL5#?=GT?LeeMGfD=Tg34KEH0D
cQ_[g9B@SG88UT):5CHZ7Z>SbBD6+R2:PK1O?Ug@NGC##W6OA3>X1>]JF<I@[4?(
gD(\TV@Q=fLDLcJHWe_XZ>&?IOAc)de+4NBL=5)6Pg3-/2c5@K\1YXB+YS:#5P:d
VTOB\08@/4,HW54X7DfIF+GI^f.@ePV=fd0Rffc47]JWBgNFJ:&f@W/ae]]+-C0N
,^?eW<1O8CQ#GT?b6U=-M5FPUQQc&cLc&8K<._NQA4gUIXdR25fQfF@9J^Le<X5[
bN&V@+gNeGW4b[B/]I/,39K-3WD&=KC?B.0fO/AVFT[3MfOa\H(c;RY4Q8;J4RS0
W?e+2-eISeY&P<H])afKF6V.VPJ0c51bFB8-;2S,6_9c=/4&9]O<=QJcbfZ(?7HN
2Q+Kc[_NK#>J]]gY.c.f#]\0EG0UdBM@[?D:9-8+cKYCe:S/;S-(N;8=#;5BQ;WB
WA.6bTef9&I#USb;-RL_TUET4Q1I(B^VJNP53(URd4IBU,C?A?:aa:>><2V]4#GK
\_8OA\U[=YJ24/4,db4c0K9c]NZW^ZgJ(;/[JUd/[1A1R05W1O7OQL>M90J955(H
d[e^94(VCZ<=HTQ3VW-/<YHOH&1KNDWZd&OF2Y]eYE)<,>_:?S7##fJR&.\cCO3U
<#O1UO/40a<?5.11I(OE3QTfPP:bCC6^46+#d?,;F>U+SaSLHR(/G,a85>,<.&&1
dZOU:Y)C#CL^R\MYWd?/R8[))LT<MTTN#]+cV?Xc3d9GR^TQ-6cGK<?b#Hf-LVc3
-H#/Y#gLNF3W?+X>MVB8R0JL>;))Q0X81FRYg,C7^aAbET6^Q=FI>&cMHZRS7./f
:S6L);=;BWM4@?J+0QU\]O3]U(Y(d;Y><1@b9fG=OdL<P,V^K_7EB=FTf8T-+0F:
(Y.J&9S(UP#H:WP1;N.X0SJ(]B/YXVCS9PHW9X9#1/_O0a0ITH_g7<gDNgX]d5dV
P@8gF@@TA_A8;V-0.HK.WOS,(Y[]W:27&\5D>E<+C.F3_T<QA=J7K8=Yd6;)c<[X
acHR?@+eH,6(Te21A?HXaRR)ER]@75J:L\4S6M-0_V3\8A/A,OP2V89/PZ)EEH(A
CK:5Q[O[K/:a36T472Gg9GK#E,(Pc;,fd6;LcF-NH]2RQ=#@c(4M+U&L:?WUFQE9
Z4SRWa[?>6QV=#1,baaJJ:dV:HfE/0=^O-=2PbH+EM)F?Ze3N[&<<dH/MU&EN-KV
<:?b9KB^WR9agSffK#(MIT_S;BUJ87.L9KN</41EJ;XKd+_/3?LZ[:(bCP8.QRS0
W0/&#6L23==\A4^IWABTLQ)Y>SYb)N]/_aC72c^UdW#,8;<E>Y+KR0QPBf84F#HD
HaTfcF6QKb#_)P6&G(b\g9\8;];:AI9HAXGF::W-=.KU+LEDJ<.dG.D>64Lf73-9
ZJ?a><+=747=I6f1=@=Vbg=6-1+EDDBacF<aE_;2;+;0Fb6U@^H9fT.0UU+c1,.H
AD^FV1>CGc\b>B6@ECR>:V:[W1I3#aLM^(dRB:Oe3Dg^UK6]BJQY+BLK?Q+d5[Sf
1W[\0eD63-S?Vd;aSdDW:fH7W+\?X\;6C,&S/eRVMF#.1Ig5HP@:+;d)[]6?N+U_
B2b7M>KgO,?@?Qd@6UYdT[_A[SaOTfQMACQ:A<[Zg&.QPN@U)A5;TGVKa509&#Te
\R7JVcV_ZQf9aF_@+9#,S[&YG1e#RA_8]8L?TPLdU_#Ce>P2I735OdEcHW9?UAKN
S0HZQN4SNF&4g3;Tg0CP)W9H?)XXN[6I.V0OHg05Lgg?K5V@ZI2=(>0KLH75eadc
RC++P?;VA?-=776E6Q\6KCE>bB90M,5=D(LWP_]3:#534RU1[\3]6&GWCE6O-G93
&cZN:cI9&,Zfg0:,Xc>b<+:\TdG._7:9+G(I&dE5,L[^I32V/Wd9f9AEC91@c#[[
E]Q]FaDA:]XEMDA1DHG[7QeGSP4GAXM7UfFM:5C_Qd^a/\T&W0_^5@HV^2HI^7^&
+6T>M\27F,fJ#YP5Y[]4&::1Ja=a\dgaNSI4A7F[#b_g>UJ>CR8;XFV[E96\70KL
&#NZ5SE,ZDGdA7[ZO&K<ZBaR0a.]d:4dDgfKc;Y8H(&UQW^b&cedP],GV^WE[1,e
H,]1R0aeZRIfS.0bGO9LXaaE.[Fg9fH[2SK)TJ.Y94T+-[^Ef,a]J<V(L4MF>#O<
R)1T<[:1+I6XaSW0;WEK\.>VBXL-=Z3BN3dPWD#a<^Wg).7GI7LY+a5MeXcX.[O1
PTLY.0f9WYSH9AH:U<J#MW@D#MS[8GE2CS+QTRaIR]6MZ-]eC9JX?E[T84_d,>:S
U#6Qe/WYWNeb[&HS21COCNVYA<&XSY\[:;H\XGXF3O+5Gc6@e.:@FdX@(;E9-9fD
84T/,.2RFYFgCM2N73P?IbK+eF.#1]#fSg:YCb4K4^-C@Z+V/O/,&\D-08QbT\a[
X\4S_\Pe+N@(O5MRK5ASb/TS_ed;LZQ-T=V4)W:=#>W4B@Rg3C0@>8Q,+g.c@U.7
1;DdWAbbO,K3E^+Wce:Ya&4==ecf1gN/f.08B_9QOgV2BgXC6?>AQ<-W8^#Q_=];
@c6]3\-FDIY2+Q>3<bK5ZK(/.[SYdMGL>dWfP<_IIcS7:VC45:QOSD--U]FM)[W#
@aC\+^+97PZ6=I(0K8^#P)U7D0QO7FH=Za.LH<X?+?R3\-N4A@Z.]N32=Z>M)9gP
J6F>H^D;1JS9M33:G:M=^,:]VAgaRgS>]_50++L2(YLB<#=VE1JYg(J86=@?e&g,
[:Dd22V@AUc@BS6?=-:=_<QYU_[2;W.OEBO2N#39XF.e7eC&::V5KE/_CNJC2Y-<
WL5I:]NT@B\U4@A6aRY9=D-Y:&Q]9#a#;\bQP]N-U-Y00[G+)0R7@?85\+eYFc#_
K8?45MU2/LYdVLO[LaN<2,8[J=/FBVJ6NJWG?CX=XFTF2ZD.I(^2@7.fO#_Q:WT.
4)-ZW0#S3A?#P<d@1MJXI&YOL.MOZ6ee<#\+0Z:BB]eZ4cUa/@.^eL[NZ)?OAdbO
;&Ybc6:[YI>AQ6&,>VaSH89)P-6ae97egaA\Lg_LD10<:BafY18MHJ)Vc_,U3OD^
8E@;<3Y(D41@O86]dfNGaLaN)?^#7U<TZ)\6/5[U(8[WbaA7L#>1KZYY#C5dd;N1
1g:KDJWZ:G2>:7@cKGR>G:V32D/0N:QEMgc)?-T>&eaF2E].L=aJEZL3,g_H1.3A
]U>(Q>9(Qc\UHa8_<DF+9CbMI)O3#C15NaID@>8PgDbZ^QTP5g??&HaS+JYTGFJ<
e78H?Rg#8L\6,;=472Zc0QG^/16]=^GC_.VC&CRO69VAb=TVPAF;\\PMf^QC_cHb
Ic^agA_CKTU>6IB91H@OLXF[XDeI^R@Ud7>X[,-J<GU;.3Y2XGT)IUYeJ+->(1##
RRPUUGZ1>O@AFLQ<L35+PV?B9TENMEQW5@P2(,JO&NS.-CHf)bN;AR.3U_>#Q3_g
Rb:XJ<?^H?\/b\9gX&?XG.192.;\)1-Xf6GQ6RUcYZ+9]T[/IS;J1a[:CXX67J/B
=Z[GK95II3@>G=5M.]O[D+U-5UZZC<X8QOY16<Z/3d_\RT8b[1dC?)IRIFR:UH0K
8e3-U\9IQaH9^-c2N^MK[Tg4gXD1]]_ERd?]P7bEGZBOOAA6dE9LMXf9SEZ;+gQ[
59BaOSaTGa)-7S^P>G[YE>;9(=:<G&^];P5?3,V5R\^Rbb\7[P6AQL0.dI]&^dG\
IU52T8MSM]44]UH?&[L^:MEf/;V)K/SO@,[P.g12Me7)g-(W@a6OD6bgG<STg8QL
T;T9UY1aR]O4<H>gD&HgMUI1?><I,Y;IgGe8(3dcA&__.J5/)#f=)<[C0K?A49V[
>OHKBL8e[4KNd#=B&;IK;MDQT>H2Y5UdH/65U4CP:/E<eN1KAFa250Cc<2T^ER.c
;I@ZX[7?=;W[0MHVB5/L=FQ3@2-7W^4NAV[VZ]U[NY6)2U0G=4X288@\eX80?FEH
5U=[Q0C>4:O\1&a(WSRUa:N1CPFAPKVf&@PE_gAJ]PgEfI9X\T<c90YC)W8P^,DS
/a4a0G>_7[LK]T74\^=aV7F1T1?V3Kg:aUP,W_@6fQC-Q>6S;B9PS(KPOSaXVWU;
19G:f6?GQY@4cIRB,1d71+80\\AQ[EFZ6#.<)295:ab;QETV.B#82aFRN<+Y1TX:
;K@)SbYC3/6>Y_+/A4[bba<AN86=IE,g;+(e^7@/YfIg3)LQ)X&ARE&PTbQTCKI\
&J68_+0c;-X&HARU<PD?dNO@d=?71&b&Q4.LaV+CZE_#03aMFSS,G?&[X>BB.HB5
6^#G_;.c2:I@gZEN?W7S>,P5WOVEB^P6(^MGZAVe\+;ZLD6=M-Dg/[W;a)QZ9M\C
,U0@EZ13g.5P;:J@eU)TKeO)IP=T<IM>3dVYATCA,e<;<UU)Q+a/09-U1;=9HLU[
<KI+R0E?W><F@Q_Y.JT:b@M_/WAg:LP=;NA.E[S-20)4;S;)1&]\C_;;FCRP&e>+
DacW/UPDPHVBA_E7XS3ZL-LWEL3K=#g3377BRNf[M(EcG]SBF\@eBe+@f=3d\X.\
[QL2<.@::E)#g\MX3>a,<@+M:<f_SaOT?KE@N5JQa6dVX18@4+HL#,+U:)^+f7bC
\G::(e?QH(W/&.XRFa@\E0bf&IG.5S>8JJ,5T#C8dU@bQe^Q4_G^&SO=]Zg?FF?a
>M8faIaNTNN23HUd<:0bDC@:2J.CM?;1((4bQVL5Ic=eF&Q]V#dg-Rg^?D7^-3e-
-S.1.L?&0>5c,O7dSD@4cGJMKPc9]^_deOU@8]ed8:X?0RNY-FIVVDd?4.U1<?9E
.-HQa1WBJ\SNZK)AIHAQFQ,fFWLg7)@a&fYZT>:8JDKe&M6A(.E,f0JQ[AO[QdK_
3ec#b6/1Y#f&]30TV2QFVEM^F@^]&?+X@8L@:FeVJXBW24KXPaC_De;);CIQ&Sb_
CEYC,Q2AU,.E,IVU:20b7#@@]HD^KG[B_O,ZWBbcK.?9OC^DPULG0>P^Z5Z4-1Fe
XHF8..b\#W@YN310H<U_L<eM?=)gN7Y9Yb0U>:7C^&6T/gYK;4-;RSbe0^3LIFL>
&>6b<3g?E.@]_;95H;c]O3)c[5-.SNZ7WZNS:\^Q(^BI/Ld#GMW.-6RP:DEYS22e
a)9+RIeKY<@P.(5U9b._<(CRADKfH6,6WQH-EQd@IMgZfX<MIYUPTI0>6d#KU[RY
STR8e^BH0KU@J8c3_G#S@VcAR<^C)?95(aTYG4/[-fb2aQB1KR\JF&bTOQ?OS-TM
XNgJd&DUI9B^?:a8,a<;5,(eB)LV-GO4JW^g#4eRc>5?7R\7:B(0KH2)PYWKfUKD
BeYN5YALIaT0??966_aU:1L1G452/6CLLfa].KU-:I@VHaLU):[QIBH+ZCLGE04Y
Xb;^SSCb;^EGFKRN)#b#_L6VY8A)A+YT@1<a^8\B&OH7#WQ30_A7@6XCT;K5e^EU
Z8.^f=H3I+[9X?P,d3;J^Y0=c:@[6;O7)6+=AYc=(A#6:Wc=e,.L5YCSeeb#c6S\
).#N&8_a38)I4)5g<FMcDRE)cRR9Y/D]&F7f0#9f8JNB7744M@0;C+REFBdXdEAP
K&H+EKKMTR-^.]fB7H6J<AFR2MCRJ72.P6&XcM<S7<T5A]e_dASDN)<],:7#<+5e
)2N>gdB-N&5=g-=+K^QZQCK>JU\>ccDELLJb=6S]0KAQYBN[WHWIH2+WUbPY5>LW
\DT#VG[\(2Y;.74E9UF,4+<=3G+&,5\+U+edPaF+Qg3,5E2Pg=2#UI#->^[c3dE^
GPVC.2Kd;eJ-+P@,B4(,a#S_^C0W0fQ]/+1:X+5ULQE?8\3OOOX>b0IYYa^H2CM]
\H.^=]]E7RQBeWEOML:6_bTI8c1M5fX2TBb(@&GBeK1afP8>b#B?+Jd?@]:4_C8-
BO=WK)[gK4EBPD<Z.7>>DIcN];0(Y:5I#Y^;0[J)UH-XWHND;&3fEU_d4ESb<;3b
5<E2_K_KaPgJGZ\D5^S,:U2cQSTLG2-fc)7X6fM?,@&L\40DM1:I&),&;5:4<,@N
GKc+_f(9Q[:DOa]2K;Wf;6K/\#/_O/TB[cS\BXD3+:B4G5799f_&XB^ZBF)<>M)T
(^5cdKa<2W/g.V8?f0(?6?/93a@NJKbDF+H6E:C)f/U0)^X4H@>R^K?&(N9M6,C8
\VV#E#2Q63[9bG^.1=U>b^B\3GZSR,TD8#2fUIJdY-5Nc+-IGSC2Ja]gH+=e_+Ad
6NC65g.OCSF7:0]1E6@.X#>#^LcACX1AYOaLR?/]P+B?9T8bL02U6.JB3-6F#BW>
Tg51@3Q70+bc?TM.H37>fAPY)ON10cR^M(2182C0H.3+L3##bG2]dFENcVV.C6EK
P[\aPB8HT@5T3#:d-AFb#DPBGaZQOX6[,/XdD)ZX.F#,ObZX7DafV5ES(K)K5&1C
5>SDP-?I/e)>dN6WR+O^+8JRFgW:3849(V2SMb<1MT+(&-(G//Hf@;RX[a)V)=9E
7\\I9]&,I-WVc0fg)U4WTCT.>NK1P-HVO?aDI>KD^_@S[@D(LQU\J8_\Ga.Y<ZB)
a5?:K94K#^SB9SGJ/OS=L+<aLg?Q+\;2&=L;DCH5,AIVaW.-7Fg)(A9)L=FI&I(X
@9S81\0T_CF\aU4Nc&86)gO<XRV#FZ?3:ZS18__O4C?W)RdcgM4]A?]C_CXQ1L@+
&@8?5AfW8U#M5VVY@0Ga\8[A/UdIb5D=,P@_27Wg7C;^H0[@]_eBGYW@.Pc3g/5Z
95]7E_F]M-W342[,(=NES=>06+QZ>=A57T5V.\E<e9=Q]@C]a/(bKbKPB[C?(H8P
YC^G>A;M>XcMI,AbKc8^@&HHYOHCU+V+6DAH_FFGc[dRBH?6\90+8&TE=T#3<>H2
&B@cI=-@BH&6WX,G@=0OZ<NQPY.fZ>ATG&B<g3[:1W4.]BLGdD=&IR,_Q>LCNag_
He5PI66727OQ#O>]O7I_Y\)(f#>E-GW):LOfG,Agg+WR<D:0V2,gWIg^8N_U#cAS
:+LUI>9;gTWTYRAUOgF84<bd)fHCPb\Ca_)HXaTD1TP#989GP5X;aP)V67)@Na-g
DK2GH9&cS6aE+[UXO2X_S6TKJd9&2:0K]=+)Y8dCI)5\(VA7A[bb-E^^P=G:L_TE
;T(>A<K<9c(K1deJP1+G:a]AadHI_b/1)f^1U67GJG@L6Eg67R[6B.3DL(9I_^0[
6N_6A1dEXN76c<LJ(N2?b]b:\0c4=aO]064:\6CHe@A)4FYcV4?R@(IFdTXK@M+L
BGcCd)BVFN_1)G>)&e/F?HYNGV/&OfGC>N0NVZc?SR;a,-4e4LM.?B#;>]1FTR>@
R]@;Y9LJ&A6&SLW:4@OMQCC5]b_QU]V#?0GL1;<(XIF6+gg#:R(d=V.3(BO10IKe
\BM(bI/abf8dNfFGa7G(51gLCE5A#6fK9ef=C0>cWH<V1K0_3KV&JgJ@>747gc]e
P@?3\[De&3HHTZC3EUAWVDdB<:PB&&eE?8N6e7(5a()UA0L?2TfJ66-fI.H&KI+B
/A7;#R2NcfMP]22,A<Y9KcM#74497HHNAgT1BB4C[N6fQ3?VD>eT6]c7Z2PG-D)M
0JJbc)1<O+8V63VO2O7Z#1ff47J-)?6YAd8NB_TJ.Ta9@c@_TK+c<UfdCS+=Z93[
IBUGXc;FK4V#4?3)\IU&dSHg.J(:W5_.=Yc^J+EY/)5#LF7YA_0(Jb..U8M3Jb-#
2Wd+04I5#B\F;=>;YccNObJ]6HS?^ZFU?#,9MF((S?U(RGQd?Z>_^5-7N3[>(C:3
2f-C_2e2PU,A=;-HK>(aR,NI-I>&7@^Oe<DDaHKSC?bbKZM)@G6bJ8Tg5+U1FV8d
<Kg331+#AT)-QQY/DJ@9bU&6U-b[@H.P6WdS\?V(/dETV9((ZZJ^=E<VA>b@K.7a
7ZTJJ4d&YRbJ9\TJeCg..#:7K\15bR,4?.N--RJ>=5)FZURd27T4DTC[@Q??7)<@
0H0MG<4\\0KEf/.M]<acBIJ-e;01VB825<FZa-a/N-=[+[KL32\EXV(KVOLOa9M^
T0D/d1<U\-d9=-ZbbDCX.?J,)G5U;H2RfS)J3S6;9GB]LJ=2b<>8f]04M4O+D))&
;.-FdI/eHL1:ANIY^WK:@;WQcJd)B#gdA;EgC4/bUfMGS5(BV+<^c06@<#cCe4&H
N@],T3;XO=/<>)/>2UIG0JQ^QeJ??@6<&;B28Qe#Xc6,RBIVP0TJ;#JI3]-,#EM:
K>KBR)=Z;gWgP_>;=e&@4J=_cIIWZbfd:5_,>8SdJ\3JXKT72.Z<W=;Fg-2?#1\K
G:GP2bMEBFTRL]F+2=#BAE@3WH(BI/MS\R12DCI>BTK&XW)UR)ETCZ(4@1(1&-f1
PV8).P_(c,YY:HFRZW:VZ&/^BVC38(4#V->@7DcBGQ,6]aV)XDD27^,;M(:;,^V+
.eC3K,T>[-],@6_O&2ZP)(B<,KV5>Af?55W2J=1KbHPG&64PT8f4F#M>MCWY:#-K
TU#K;eDXbSGT(TZ7K00^LO[f6BEA.3EB]5F_6\ae;BCJSEVV108_fYe6dW?#MX4U
4dB]^7Yd=ZPY>_e+)<7PD]f@3O]6E)-VS\,OeLg0)>9-ZEWXLJSSC=e?G_)]ZVT0
5aScZ/fE68)B\)?U8(C)F:6[M-;#(HQB9)>.M?I\+c&[_@J?<)9Y[EO7+9>U4/>[
<1.F&E>/]=XS-:M=<\8bO_<O@UQ6Wb5-QW_;5b&6E>=b9+6.ULV>.-KV;0.<_#:A
?Q+aR5e,f541<-+WF_:W94J4f+:,UC^SL:85_AaJLL6DcLECIUY=&d2Z;OU4G>6S
^9,dY?0=FGE+1[3:bWeY@PB59,5E/(.LG+:fVF/6+#-#_6RKH9QSX#1[75U41JN0
2(DZ,)AWFd/)1bX(.TZg&#5H_E-Ja.e,d9c9)4g:XB^>D_K=a/0NgP8eSf0SKbQg
F7;RIBR5Qf22RgF+L21e<.A;fJb<IG@14FB:=P(L9GC9J)EO@5&+F2P0@4=^B(^P
DULH=16U[Z<>TKM0NSC6>eE;fg4>=DWTbI/V,I7fMd70^XcMKfK7K)6d^c3+:DD0
K)F<W]LMA8;K0cZ531A:1\7W1@;I(C2C0+/6#B;]=10H\3U]dacA_C3NU#C-d?PK
?.BA;^gb::>ef):?Q7D35:^4U^^aN(A@\B29Y@V#@V?Pc]M].eD&R/_LJe(FV0T,
6>#g+U.A94^b3gY]#VESQ=^/R)@c\/UD4B:4-e0#;+4J;4gEU]N6^=37EW<IA4QJ
=-07WHdMYKR7e(V[]2I0TAT5(L@_4:K7&8]IH-C9/7#1S_K-?KNb?2+,\G>90]-V
:#ZUDF(M(EFIQ1THQS-2[2/,CdUB+6WCGfL(>H[#54?N<ENOdTg0LHD\YY6-MU5T
)&RIK>PFU;I(-f.#Y3?QV80(/RA+Sb312<[.T[g3.NC+O?DQbd&)UN8UZ0&,@YQb
.A7WF5e-=GdQf.V7NDSdM\f&e.G5=[,SU:RL\aYIK8bcUdBG>>[KY-(W+PTP8G:-
5?279><c=L@aZ(T.?PW=H>>.SH[09;-2FB:+Bcg8HW,&=Z=F/G=FZ[P0Rc=CS\PO
?7(O(OR?)==F@T3AMM1acD-YO[8^82[_aDXOLO;_[IgE&ca/N62_V@;RFN\5N?PT
;,8-^G8[SBDRb?e4?@<SA/e9WEWG&9/Fb/be4K9fDg83SOdKU:JS-VF&-IC\1fS&
^&/fKC(74G4P4YUdBE9H+F;MV\\&bPeWF]77@FfRF&5MTA)AY&LS^g]FNAMeM]W@
bBD8&eU:E47@_@42^,<aWK#<.3G-@LVWY-2O;7FL:5INGJ8(bC[8YJ&8-C&3:P8D
9]JJ42KBV7Q(.Q@XfeXf@;b8?>4.L27C&Q3=&6[b+JF>>7&-+EV\6\2.<cc7&[[e
O2O/R8\fS^X>Db#?>>a/^EA/?@1-RDR@LPP@D]/^Kc<LIZ/\,OHa_53/KX5XQ;)d
EVUV?8O24fLg[,5D97G\CFY<,E]J9^YH;cG=HO;8Cc&4A9:CI[McaB7Ie;D_Tg-f
(b?YJZAD+APD@-M/<L?/,a:#(B]4;Q&K)P\gPM>BH\42,)NAUNNGF]X^MZR</U([
R6d>])&OV4.QI>VEH9V]6OgecEcO&Qg^/+/g0f?5_++)-9=74,2>cb2MgI=DTDL[
3<dYB6.C<5,C7[AR>E?ILM(.GaC7AKF<Le+ZMV3O0F#TAI7L<?-Ofa)4;@A@Ge3)
POO06X)E3,>T>d>@J]aWR7bU:Z?;4;a/5L8@^V5Z6eQRAXB\9&2JAV.dAgeJX5-J
Q3ce;6G7XeM4gDP[LK9.G7^BK)9]XFW]<GQaC(=e9?/=-/5:[5Tg?Q^0FEOM,[&&
U\?>.02WJBP,3?Rf^:L;d?:J7-a4eS\3M1I]NdbMVXY-1[ZY3AWD:V<H9ID5NIXX
JA(:+32D,J(+SGe7XSHJ<b_\eSABIEG.7-\c)O:3^;6&)-<\eYQ.8Q3=6.?&)=S?
Y/RR;dE.cIU_dJ2a\-R433A6EcEaNDIX]/SYc0-NJf=QOYQH&FML6Vb=3SV@V7P4
LE+LC_dEF05,JX/6ga4CaEAOAcD<e;,JYX;?D\R,Q_]/C-O/5;VFH^&?IG&+_F[9
FI]Vc>W[GW&a;B3TK1Ug)=,I/5MG7Q)C<A>2^1_I#DT2-+.LgHb./KHAXJe7:PD:
)MQ&:/WfS4X)LML8[0VcH;f7dLQ[HF<b2C4L.b-=DBfDLO)UGD,a=.>0H/NR:4/[
P_0V?4I<CI]8SBWVSUL)b.4X]5F_gZDb]@X;4&&ENCY)V)[,0<]#D?P([KOC5<;+
JQ-TcIK<N2US7/g5XF6I<.AFGcURPTb]c.)D7g,G&@GZKaAKL^[)W7GXF_92I:D(
B;N-\c#LeHUf39L8FP;@BL97<;/P^@cV,/@^MZb2(QYN+OU=QIJC3HIg2L:M0PLg
<^M/WZccCYf+?.2F6X=)]f+XXF-A?PW?gON-80ZegLW)4e\95:afH.54E/WS8:3e
U&d=C71^\-5LW+]S.YJR(5ZU_-U]#UNQ3+RY5S4KMUO=Lcac>+C8(Yf5bAc>SAP6
d(;8S,Y4VP?_f18#(66>YCCR,.KHIe6A2X?L(-2cL7/>C=[YIeK2AdB.-/F=d1>F
>^68.<EHR4+<._VSc\IP&[,feP^#N2;>9]I,JO7)OBN4R>fR35YU^\:2ZMCTC>f9
L:ER-9>1E/=OW#a^KSOPH#f>W3caUZc<a/L\OBIMa-aI3;P/@2eF8)4c_Y2f1K/,
6_Y60<5]e,GBL2,M+S[6,232&;6M2N:2&g=Y4>2bAXbbR[8JI8d.cL3fB]]X.;6b
a7QFAVOZK&52MG9Y;ZX.V0BPf^b9-#S;_3LR5#B4,b]2OHX718A&;AWbBZ>cYbZ4
_?85F/^c[8B,VS3cgU]XG0S)_6A9A^LP4XET6J8^?\]H(CVJ&XRW.Mg_\:DbWd[V
a1157IPL7K\BR<XR&.E3?002fM<J96W@JVEG31FHb2FL,>5?JS3\Y10A/T-L?P:P
L&..L7JQg,@gGL,G:FfFb\?]RJfFQ)6W\cMa]KDES=ebC?GLI/H6_R3PRe:(M(Na
1LP[XU^JZFL2#N-(45-21E=,[H-/:b\43K]MHL.?L9?)bd^^U>BeT)Lc&e3OWAZI
PRWV\U;#\U>F8@MPVeBF<H)?5VODP[1NSC3fT<HOI96QcH\b<eKQ)A88eD@(]C:B
U1X_-K6fJKGYe213_?U<APca/(-/=\MIM+GDcSa5f]8FFX+NQ;bdOO.U]YN;58\K
D>DWV+5U_8\&1,<=GH?1\6aegW[:bZJ+_:R\NLZKCT(5AJQ7b2=[G2426.b2e-,c
H2PD)B/E[BX7D#488^74]IQLO(f]NWH#??(/@\/>O^NYZRR?13]+8<]&PDc,>U&5
G\]geVgeH9NH.(,\MXgPS)3>SN>)[W\\Z9?Wc+eNb<DL.05<&MU,DLQANcEIFJFC
Wa^F8AH:)5Z<bMJ.)NTU.Vba#ATVf>V<&PLC=\::cLgBC-LGFUM[AD9TEM[+X6>a
,;Y<=_Se]EYfJ#-/@14M#LOHA-^Q]QU<GafWM9Y^C^Ig&7@4>=#:MGM>ZFZ?bN7(
0VV5Q-5c^+c93,5V&ZJ#P&,DSLPMAAf?dT.-E8D81:CB3W:Y-RR9GYbQO;2B7/D>
6g-V]TUgK16<4C^^4]>[K9BE35edZ9Z/8OTBdb\?KP3=0>>+-<-)IU:ZRYgdQS[,
\.(B(?9)JMaTGW>]g91WTP&?:6+151#W/J:68J.S/E#F8Ce/@6&2L;b\OV,>aaUS
W:-,WW9R8<0a&L1b#HREb?Q)8-3ZIIP&RM0a@PH7NI]=2IQ+P1Wb[<,OY\TAGL;d
@V>X20E.DAT#6fQ)9EbD8^U@MEcgDF-d(M8aBc\XE8>-,/CE&;MgO.5S33-IHW6#
2cT:C62_-ZegH5J4Ye.C+b5Oa1MNM+cg0SGYG-d9CKc?G6G^8.06NKGbZObb5P3<
XMP?WGM&9Cf@,[_e>@]cEZc3e6G\&WL8_JC27Kf?\CG,),Y1/Q?W&C?LH#J1GF^S
DTEX.E[9d?Q(JGRG3B?YWLI4b-/bM10L8H53F9?>H?fQ0W=e?R#QJbK-4Q[BD6Q;
;eWgP3SV<6Q;#E,Y.\)eGPJ(3H7c1):(J8IC_TJ[7I@6c&X.KF9c#;=UUfg?9EDd
WU><RJPEY2493/.5DBe\)K:#c<8;(OeHWOSECL)?\3^VAc-DL7F2.>N[fd\#0L)H
@S9<=,<:;]/W-Ubd4?0#TPdNE-JGX_7TP;eY_1H)f5C.M<QKO2GM=HMFM17NU5K9
,_-ED(B_T:Xa=,&7ZgN@Y@XK[2c6HRUS#AO@e?25M;gLNd^D<?N0(]8:dd4>N5Y4
9>+2f=9c&IHA/7R;)P(P>TL&21<MRRDdT2H8<(O,fV,-V+.Rc6g2\:6BZMbYAgHP
<?IQM151KRf=U92RXdAAeO>/&a74J7/gM0MU5FK/K8QB86N(K[J(GdZ5[S:]daA:
5>S+MYOQ5+e))6G4UPF)&JNNf@W/\<:MaY7X]3RL_;LbgL??S0cM)S1b\OGf0?(@
TUB8:=TO^-==@eI5I8KM)5=4A#cQf3U^DD8;(@8TeA:cF<6]fERYW#@ID^eLZaAI
PbCfb8[J0X;&7^,VdUT8,&I_@gU@HO5c@VUHF>6HAXB;8d;e\K<WIF8N7aa3.e.A
5[QceE>Y_^=&&J=&XA+>@LG+G,ACQFI@XNBO:-7^L2Ha1^>)LbL.,f+eXH9,GWIH
P(\L7;d984<=a,SKE#FW?/,R76J]^46+3U[F@@WCNT:LTU;&9+/N)//0S1)0[W,;
#J^<61JPW_-JP=/Q(f9\H5Z.M5;6+]?HK?;Zf5;:-#WH<HX^9f^2UN>R;/XS_,EZ
F7&T@8ga7TL><GN]3E+LHHJQN&bF,U,(I;Q=3c9O.EZ]SC4#>8gB3@#I=PUgGJ]T
G\R6-O.gZ=>H7bM#1F^S7?I\@ffY&cGF\?JQN51UN#\BU)eP8JH)CPP/V_^)70GK
4,R64=8?T9YbDX+fSU]6<WM0G/EV+?/1[EX&-<R]:T>Aa[2KI;XL3C/Ub@_K>\XJ
KB@L>Z^(&3&RfHYQ>D?H#@fW9(1O]dd]a+:>P0J-#7IeXGE,5^aB@;,2fb++2,7L
@79K+5CEa7X(&[OG,?]G)>(C=/Z-8We5-.2IE)RcX1P(UT1[e4-15WJ0F=7\V;VG
ZIH&cb=_K^G,^TA&S48Sf#+4Y,02JgA8+WXTW73;4:b_HV604?-_M5\LEI<[OZ\b
6F]]QW]O7KJE=gWGaG/ZB:/GfHc7LBJQ>_T:OMU:82[[-YIYSM6FfVV8f.IE?V7f
eN5,e.:0^.SS<BHG?@2PYNE1AVJ#8P@fg5b2/T5c.C>S^4PKJ91]:OVHN)5;9X2/
WBL5P=>N2dfRb<KD=Q9;FZ,[>\fU5<;:d\2]7#Af#3)4#)MeO2Q_GYE7JCfT99[.
^AddZ1^1I/;1bSGP/G]5BH0SE2DL=,=ZJX\CU:MCD^+c7_.L-b[F-IQ?+:aDaMFV
SE>:c0<P<2:f8:#QFK?]?EVK2#0F1_^UaJDS2-,/eS:../W5YBW#bWBSJ/eRVE\W
1-[#LA+<960<G:4,gXfbST0eD<4Z]2a,^0UQa_QZfY).OEQ.<4I1g6V?NIQNV=.V
1U:^P;9YDI.P^2ZSX:4E<Zf;Be-.fE6\S7?-<S751,3:?F4Y7,L>0&[]+(b11gcT
AWg?WRZZ#J><;bACY8^,a(8:@.,V)8666D27&5#&bO_:P&0EEE_X:(f(IF0=..]S
;HY5Cf.G&1-(b/:3/P/.8&WBL6^K]\5<CI]0\FDg_Kd2N_fJAePGca(+]5c-(+?(
:YSDLf/0)X_BPXCK+4/FT&W(+I\g5N7a#VeGT)60A:g6)FWC).QWSC6@\=59GPB;
e^(OL5O7EYPP>dHdaLL/.(>_.&USgFE^]<7cW;a=(WgP=Y<Q56R=86/,_IR_27/S
PeI7Z0V6D[Nb-HLQR0HD4-5BJZP6GT-e4HOI?U,5Z9=^>Zbce8(:-(-NfX4^PAaD
FeNeXXH(-:Y@LdILS(@c.>V1T[23RAeg<(AJgF-/\7/N]Y^#BX(&#;I[U.UYBQd=
+FLdU=2@2M7.W@,4=5TcX?SOR#[Q.N+a.f/&+>=+HcH=X3:TQW7R4_DSDe_/_)I#
\6Z2-3CaUFDbQ<f@Ka(:5^d.<YUN750fN?Z00Qd\<G3=)K1),RVRNgG>+\T0>E72
dO&KJFE,@f7.R-O0V,ZLKCS5A?Bc=Rda.gT@)Sa<MB7/I-Uf,[aX&5e:09<+6S/d
<]+6=GRD,YXY;W/5=OMd00>8^+SI?HJBN/ZOF_T\YKQ(58aIe?>cV@+0[/a+.1,2
:UW8=gAIVIU.(5;4U]2XM9eU28B;902##/g95G\3\Y?10/gZf_M,:6W8)B&,S-(8
F-HFSc/Ga./(a?,QdULOTZ1ADJd<)DgOfC-(8SeE8_DVX04QWB)E&A-gU:dc5H2L
DEZH5(XJe8J>,SRM^ORGN-5^Z2dQ1_2.K/GK#?W#[20LcG@^He^4,+SQ8_GPbTb4
_N(CA@dL-)@:9XKc_.B\GcRYJTVQ1;?a4_AJXcB[++1@bf?^E.@&BVI\MTUd#9?E
39E8+HLO)4D=K:e_Q;[0@.7_QE&IQ2@_g_<NYc/ES93K30VgD2KIN4^/aXDA=&FI
@0J332=3&@/K9^aM5+@5R6Hc&&X1<>;(R+;EXb?04^;XU9]Ib?5TRfF(=4)?;:X.
VUB@#3_YV7\WF4WYT@HCUJ&>RgKZcTR@5g@?00>>NS)g75IH>c80ab):4GX[NRb2
M96N&1S?)7J6a&5L_O8PJIBSX[dNECFB9D3Z5:]?,F)b-/G(D^_F/7QJ\SIb_-bf
-4aPHbR#.&V>c5MEK4-:EgI=2,9J59Q([ZGO8YIBgJA7LE=98#W&NW>fM7[5K>+/
&Ja5R=F:&(bSU=IF(>+&3;eO@\_M73OefHJ(#a9VD?OAA=Q>AO3Age-3O?,:/==B
DfI\E@8SU])8>[>QJP82I?FW[1G>+NKP.K@1\?CL.^b0?QXE4NK7YPJY1XWIAJ\&
<-W0QZ.]/76RI)3-JJ>Y1(K,#2=O2,O5PGLZ7c2G)<:QV6N=Ie3#f#IHOB^3K4BD
D,EEN=FcCKf[R+,Q;+CSeg34G:9KTe?gLCEC.RO:dMgQcgNW,+]OB2eS=C935?S-
W?0=4;/FL6-]9]<AC>c@TXEfM\F1Y/^ga6J@M;H?WJR->29=(;6dS]HD>;C&R^#_
Q_/Y4Wc(JIS.CLA;EDMA#N/79E5]HQ==.NOW^.6(;JZZ<ZQ8PYaN6_CW-RLGG-7W
=G^CJdQ,EEN\B#7P.gV>@@0IbS\3eg#8)2X89-#e76:E<OL4=GX9DcV@6)b?f;<,
ER@V4/^:^]+ZP?)cCbUMDBN.6c(g:]SNF+KVXeDLW=CK:=X&I,Q]?&V-LR;#0Def
:YL55<OSU>&)eG@)SV3OAY3Z-LA^:1g[YWY+@;(e4IQ/eJPN&J;NY2<#L57AOHe#
4Bb1Y3;55/RK_TS+7))(PC7bY>/QSNW04G1W&9H:2LJU5^8CGIbAOZfHEJcJ=USJ
66;;2)V2;HX^L&BUP@1Y@,F\_c_QcHHHU9-H(?#SB]9G;9U&=U4M-MZNBcS_GeD(
+c?Q[f[,9aV(;e-P+a.1<=ED?<.2&YVR1:f&@C[LQAGcPZBH^(BE^QE;ZT;DRX:a
/Qg&:6;,GYZER_7Qb/Q>&>JI<MUX6VBg=[;+\Ya@QJ4=PWNd>XaNCaV2,X=?C9PI
c^-D7fP-@TgT8A3G2BQ(HP&+UWVGP1O1@P=<f&<fB;H(93XZb,YeQ9;e5K[/I)\d
aU=\N&f.Rd(PdA+Q\T;DPDHgb:LDQ_G?X84gW:^(&WRLIY(\++aC?_Q,TceI+7f@
\&CIe#I>5N7GA+SeD=gC)b#6^;^dd;<KfAgWdE:^TQKZUE(R.X8HLLa=Cd<_@>Tf
e3BX[GF(QDO)C-:VY=<&5+4,-cb?.4cf)=7XWQcKYebM_/&EaY;Tc45857C&O[^F
LV?4<6I3ETPG9L0bbZ_OOC^PYIf&XH5OS7HSc<-/E9Z<4LUJ/\B/[cK>FGKHJ+.Q
I:RM(fI2]+6NX6g2+KNG+NJO:L>1TR[Zb@]P8]?P4BWX,DfAH\R?#(J\)E9)=4Y1
;BGD:7AT;U0):IF4804IOB#E-g1]<Q<NDE\fCbT(L-MdTZQPWI@9)-690YZc])&(
2XbSF.YITW[R5]3=(2HAM]L>HM2DL/P#E<9.)H?4_Rc1HRb[dODeVV@Te_d3[IH)
+T7E==K7KFO;0)7b5H_W[37(e5/_]J@6>UOdK&4U(@];6@_-^]CULY)[cdXgVHgN
[PHE19<9b\H_4g=T#B4I.cWG[gVA-Y(WVP5]Fa?+2.aaa02J6G@ZWQE5BIFaR:Z^
;#6aV?]&I@GM4d,I;Q[P&2)1[HfUW3.QI_LI&W7I,]5H&#((D=Wf[S(+^MAZ7e1G
U-S8INCT1-[dU-.\<^H)F1S5KD&?YH.cRU-WcIA,?Ac@^d)@OSJU>BB;UBI/16L6
_)]M)d_\(1(N)(L9I5;6^d9(PD_O_Me]M&JE3d;Gf15UX=fX>1_=4^9\1d(PfVEK
03<492EV8eS2;P>X7aEH1S[+M-<QcYR0Q,LC9&.)JVL&RaFK?KU-8VDNddfQ1a<&
67W/&2?,<EXTa=(dbA9BEAAb[P2#J5BVC00)[1eTPUd.F5O(YZ__16QGVMN5B\L-
32E7<(#M34M>)^^#a<SA&SZS)TB^_g>HI_Xe#^_I5B9M3_R:]ABeO),HEY>UA4[\
AA:,GHXS]S/58Q(OTQC4QO8&QW9G4D6FIX:1+c(DJ/Z_3O?NR3Rf3+0_/de#R\[4
1c:dG36Ge)eQY553+4aU^c1+Ad9.P3+MK:fgOF=P.H]4S&QNR3Y)7[OV91[V6C]@
;bTV^,QI:X3M=(J7H/f::AH0,W)?\L.-K^UfQc339=aC38DKccLR^=,fV\b2RDOQ
e,>EK7H^A\RWd+M\9H:)WW0SMd&/cLLI1K+>/LDYB#O@[RB>#WgNYC3V-D6PI.I4
SZ#,[RL\HAdV>&J-(83ZRQ#V[EAD_9]ZLVf0>G3I]OEOK-+V:]e[G&C=3dBKb@E9
L,VS;BXSGHbOQK[T[&SUa7&]NF4C75V&_8U?DT/V-Ug6R:B2^283?<f/A#+&\&?I
JA9MCZ[A_1T(fA^7D2&aVa3,K3#-Z[\:=N8Tc(;\Jba+LV>G,09fDGaJ+-K0&6V8
A:I/)d]079EE,YSJ20K#fP,_+R<#FBCf9TOTL&PSIQ2Pc6Tf8bVXQZP3F6<YK/R5
JH8gQ-H+=V]JZE6N-5V-c^,TCQ#SQ7-(HGS^\9fF>ceS9gbe.Df9F;+B+H_:2;Ag
.T[#UEOeB\OR\I=SAd\2&Z9I@3JK255.?B<T?-M0O<EM8/Ze=NA-\a]MdZ^=DLDU
>40FKJ2NA<5.SB4X^W&<GJ7)H>N<.5([_A3E/6YK,NB1K;0+CFQPFD4L?W?CFBAC
8^T8cM#VeYQ6UC)VeFX&\6ZRW660&B\WKHXUAX^UaFG46RMS,^W)2f.c:P]D9SR6
JKI&LKR=J#)&2f-AEM7cAOM/P7B:O7E]@Qab=[C,;dV/+=IL@e[5W,O5?(F#eMM6
_BKFM,9?;25W99f8NH4QGG)6EfNTYR5(f?N=HN/B1[ILd+Q670)CUdC]HTg\_2F]
f<&RUT(+/FF(<](YZ^&I#7\&A)NTLK6B)P_H,SWGg_)7XH&OQb=,FM6LXZSZTX1(
dfVU@79MOZYC75gCD(O0AQ98S+(B\g<dIV-YI8f(CPc5;gG7HA(QEV;>#9Wa-]@:
gUV2H8?IdX#dAI/gDe)YF\8=Z;2=2)D7[9L\,Z)H5@6+^>?ES^&=2e?M6&R<MA5B
)Z#=?aL&cMJ@]g,:^T6TE(D,M>)egZX9XU,H(1[S9@X&1UQ2.AdQc=K<X&Z5P&4g
OP3W,JKYEP4R[O6HLCfWU=Mb5X9Da8LR2R0J==?41DS;:3Z(1IBF_&5M<2Vf<W2B
E#g/7P&@M:8O68HU,=7S\FVK1F?X_>7gHD0TeCQ4E;,McZ)?<>d;/8SD;^#HQ#gG
b3e0ZOXF4FFb[ZA]@9/:_)-4FQH>RWOMN+]IXfT?CZ1_-fU:,G/W#e&?.G_IJ=Nd
YQX[f]Cg[W[S63X;Y.#&4_VTeX9Q,7[3SKF/#&6RNEDHTXP;:aeJV[)2(K0\D[HX
&5(;.aUO10HXOEY>F4N+)UY9TC?5?Ve76X^@9#Ff-HEC0,HBA,PA;^T/_/J#P52J
&0WAX=^G1+EeB8g:)AUX\)Q-0;PCZ>KeIB8e2QQ6eNMU?HP/XLC?G]2Q[ZEL^0W>
NK<)\<Z<NCRZ3#^O,]C/[C]3_^>g,#-+FFNfI>Z<V4+c:R=[P-(Q_.c+WBMK@.8[
O-+??/Q6Xdd4<46IEHL1d?WJ6_QCZUE[(EH]9FA8A1]+1bI@-0K/f73_Z^AH1ANa
e]e6B2B[ISPV/3aa4T,20Oc]MTfP_8Z1L]58?Z+gg/GdBG6)6d:;Y)>_:FAFR]#,
M=@A:EXCTCW[&T[202aY9CJe3.3e565)FJE2:=E#cZ0ZG7,=V.bbVbELU)RLAP?f
dCP_.1=;R\SZKH3>DO1E-/gJEKS+[3329D91=\^TB:\>Q+1[g(>#EEPD@H47O,P\
f#d+a6?PD06HY<=,,D7V\,.9LeV/FP12>Y>><Q>LCD4D0DO-1bAHcD>\,e07YYC;
M[A.V5SG^M\9?4BgF<;e>b^/K5VWN?EX-_++KL4:8&bDQ2,]AAN)cIO1GQ&QfS1b
SECG2FbdX50bT;Nb+A--ZWOIM]E1[RJ<#XVV8JeH28TMALOHb/:J)D)6Ag5,-f(6
EV#QUCJ(HJLc5B24_UQA,J3#[F[V29<g5I\2TY<;V:<<^?FNIbPK6PF<^0f:3RM\
aFD=C@F=O)QX/BI=MVMW>_fJaXbgTSAbHb@;gL;S#eP;dJ((KLG=Jf>9d_>:bYB,
e<AGO,Y(b6HX;_+OPGN\eLUN=JR\bDS)KF6e]V<=R<[bL(I-ZSa04K05HHL(2^E7
fFHX&H<@S9XNZ[Pb,(\_S>:7ES:db,GQB+5+GQfeg[7_cW_+Wa1fFA=@CM2Y]b2X
U[UL6GOd=fEP@O[Z(GJZbU[(I-bd7(5&<MA&1JN6+VUNQeB98O5.\4ZRK8BS@e<?
&>.aafIM28+OVTF3N=fUQYJP,_#TOM([gZ8/]6&PK=U#7/7X_G+M(FRB;<0K5H)>
V^QbJQ+\P(-g69\:0Qca)@\ZI;X2Q.X1abIYPS.Z/gEYc-(G0b1@8VK;e9,^]/N/
5gcg>U7^dCYeC?\#Y[U+@0I?_UBUdS+(aZPLI@_GP[2[PTW]IdESJX\C)5XDIG6/
7LO6CfSc2QT60a/#\?Gf5fQ7(M0;&@<)Tf_LORPTH;CO>U.9cg,bY86H\4;9Wf1.
(/\+#:#V=5-3MF/UVgZ8<1S:4b_<a?e:c3+P5DWR&9+WfTTAX&HA):10NUNO/fI.
^/3db1/Y6/LKd=a7\2)N0CU>)8NCBL-PBK]g@J>2A/HUGZPW#+_1-OX&G=bUg>eB
9&Mf,PY&+Y8&F[]5QJ5ABgZ?Q\8-C;Pb+Ob#]:ID>1:-^gHT<\=VJE8=,H5JWeI4
1[&]S&P_F#F<.9c>27b8-[BF]3F,@KXO//T[7FSEG7b=##.N/D:e@E]+MbRIOJ@2
e^TYIfF_6f\c)/)G&7=@]J1f#H14Mf2@f.(Q\-<NV?@U;W3eA,>U,gEAT:<:70A>
O/NU:7CAKZUFUQL/OF@FWfXDNe0Nd7P^Z?ECNA_2P7#_ZJ&O=T-T?3?](L2/^QfE
FOb)DG0B.&bc4Aa)d],0;]XdEI0^7gDcZ7->7#gY1YNeR/T<A=_gPf\.WcPBa(<\
d?S-I4YVI-R092@[dJT+(V\^[^N,=51P8R0,KJ_eS^NAeR9GY\&Ef7M/=Jd0(BJZ
2R<V/QOQ>LGc]EE5^9g0^2?VY:IZS-2N(DFVGfYRB5G_cUE]^GYXES1E+-DE-Z:#
^5\SQVa7KYU?K[MR4GO?-Z^?WeaBVP-F=MWMOPaGUa]YSK&ReHaXH[@M:_6#NSX:
UDbc-WB5+70ee]H53\:8^\d]DfEJ2RX>3O/@^IM,_#6JR,O&E#]A,^\F6^ZA2aUN
B)bT)CGWR#a#>ON;RNF_NQdfdCT47OD10W;A+WcPRcYfE>[ga3g^Q842FU./MG=R
:CCcc/-BY2CcAfWJ/.VQ?S8VFd..SI4#e;Pa1ebYSR75P]@35-/dJZ84b_S[1/PP
H-g3QQJ@]06.-.QebM]dA2SW7+Y7W)W^fJW8P\Y_00AX:F-/,>=-G46AN#Wg2G;\
7O?[Q1a.1UPUE]OEWN0PIK2X.LGFB+c=JY1.[0fJUIHCYa,+2J>:&+]aY+a\0HTA
7RFPULSe6TWg+KO?0VNC2eO[aT.?04aHBL1NH5Q#FI5ae>g6L8(7@DQNN,aGGW2G
BE5=)]Z:a&SVK.g::P0+aNHEION&Z@AHT&M+.W.>KG-a+b#QF05g1DS.U_H<85Fc
J:Ze+B20@=)7I&I365HXS9U/Y6_J<+&WJTBJ@+-NBW_?Q\7.>&?OOU7gOG-W(.Hd
5W&aE6)/ZJ@4X300?^e?L<9YB^P^>H^(fW\_45:3Q1TRANS1I:OL]-I&JbD4b\((
R0c4H31Zd;&R2D#NXK>N#_Q4-?F1&GY>[1Q#)V7-JcPQeXO+=1f-R_H1<K)fL+Qc
/PG,U_gJV5bWRL9T1C&?)C,N5--YIDT7LF;@2Q8YMJ@#WE:.,HG5M-MeU;WD(1.W
-R:cR)NL,LGf&fM[+EKF+VJ6bUXPcMQ2R14L1Q^0.YJ;c9WY&SVL9I#U\b-I--/G
\69D[2f#@]A+_NOP[CCG->-g>,_D4Qf9ZY_<5K]JS;bDdFFJS)A3)]^X6a_E^2E+
RR7FI-6EeeBC>WG-SZG(F^)^,fg4J>VJH8>-6aI&UORMQb.g[,+EB0R#1^aH-@8G
W^WIAI;\9@[Zc<@(N/XM&25TA23Y_ZDVIZ2gHHa;^3E<3])gZATVQQY^XQVBG7[4
OebTX3gT],Z8:A+-Q8WW(f)@58G5/QIgY9M>0VPLL>1#VZH)7:XGN9)df7<_\d>+
E^ZY[\^R:GS6J3Q8)dCZ91eF/f^&?ZMSPHR\^CeQ\H8#aUV@OV@Y9S?^8&G[+0)-
(4LUO9G=6>;BdQ5a/5<H99f?WMO4.+)EJPSR=2#JDW<Y:Rb8OC]aK-97fN)JP+D7
HX<@TZ4Je7,4T,N/<RB^-DaR98KL]E.K?4_7@#O&::5fW;c3_)ESFCdb@d50GW2/
X2LHFARVG8BQSaPH^b1>WeU+b0@f</FG,.9@@.-5CU5KMIM1.J+(Q-)#K0;A6XNM
gI3[5c,FQD_[,>0[?S/YVLE5C[_De0<->\d7X;6<TNJ4Md^1(<0-;#1DL=<S5N-N
.NZ&Y3@YKKI+2[8dP,.Y/)V<<&IYcP_?ZW<;A)-7N(3[1He30SFZW+R>ZGfA#=^N
7LU>[^V<8<cd\SXCGI1=15TE_XAGZWUB;dYB^Q<,#&3T^6W3UE1XXbECDV/.^bcc
B@+-aCMHVbBOK0W/+UK[-(/H.dVT^\=cW+P]R&XAN+Ve@7NHA:A+4L#K6X=aaeU-
4cXJOP=Rd1VI#W.NR5(7>#.9LMIL:-FAXJYe@F<LN]5SX;[GJ.FO1^?O#R(1#W\g
T(TK3d,T1DCCL3U8-:/\[?6fBTVN@IfARBS4]9dKY.1)g\468-9/:3>C&5)IAH5E
((5Q<1;^9)AB0K7U[2&O5F-GL\MaF:-fTZbc5@-3=N,DdU)H<0-C;Ja6//fCV4IO
3@420+QXa)b-PHEY(<3Q7T@H>;SU^aRF5-^=;@d/G_\?gI&G3O)LT<caN:Y_BLZH
D;fSdHL,[agTf,0U<?+f__50,bbb@?_I65eC_FG0,)8-f2ZWS=DaJRY^9PN>#Q0U
05X<@IT#8Y<RLN,6PUN,#WX+C0Y-T-\VeSK+]\0],T4QaT/8dZ0FXE?X->V>e>)]
\3_F:c5=;[7b_7[NWT&W@8PPW3&\e0(53;EcTAX#FdF4<=cH-?XG&H)^@IQb(O-8
7WKbL/W6SI[W.c[9:;P>>.gBOTLca[\^1EbNWMT5ZHM=PH.+VECgcSLZIUC<Y4ag
N2Z=/?M,-YPEHBE:1\AVHETeX^f7HBKG-@-)L8<K#=cG4/cUM3P6<)O(e/Z7HOEF
1J&=9M6T,Z,6_fAYOLPB:eeHfP>M:HO^/e^4)Me5D_1+JOQ7UF+e-c=WAeI]\_QD
XSYQ8(Q^O6&+F+UDMGVE+c9aBgbD(/KDI=EF+@[_A)[g:c?cU>eRW+<dXSP.cf&_
b9E^b+?:X]WQ20WT(7[OQd.R-M6H#K7^8KZD:K3IgfYCDZ2^1)/[C>>SWZD:b4HP
?/:@F1S2gE#+A:)A>B@&Ab.8&U7]\L24:9G,K]_X;GIO(b3^BQEXRaZB]RHe[(.=
1,SX8J00YL^VB=NNHUWH3X6EI1=,Q7^(:d_DL^SEEBQ(:>fBa(D\5TaT([8bN7>,
EOISRf];c[PYOWBW_8QXS&fD+\?TPN&KfdS5M;Tb8=Qa9QB-]FRHI(0YRK@+bUR(
:g<@Ic^JNa9)P6??419=aK>QbH+eJ+]^)RS^_Y=HB+L.f?G/e+.=C=E9]J#/ESS<
^HD:(D&d30RBCfgCGT&f@CE1R1)HVf<eBTeT6>FV^+F@.J03U^bCW78M+N\JGg=6
;5[O(ND1TT>1#TMGdRVT.0LRaP,VRS5_bS);)5H<C=\&?95=_1ef;\0Z0]+_O4S\
.D6Lg[g&fX6.Xg][edfY=8<G1cU5:LD=R@IHQ3LT-<WYH4W2:X&&4O\PFL(?+(Kc
3WR.dLXe<MNF.G+4.PfNBLODP>XT)XS+?>LfSdYXCeB;@E[a/g3M2L.f,3fTKb.^
EC>DKGDRPf67P+)5FR@R+)6IV^\XIBP8]a_2)L/RUGgOEb5?X4+7:?BQ9&RUgS\9
d:.Vd4>3He_Q/5JF5^gL)\+:SM+?A6\3Ae4,Ec7=NL?BZ9-\741f0T0TUQeAA_g&
Q)\.0^f?bF6aPeF7#FWdbU:TY<6SF<&AOVN>V)_/(&YD-I-.>b(_2cP)<IGN&JZ0
RF#QW#;^9dWY,F;:-)_^5Tg5J1A0L0C3#Ub]:VH#8^]#TXNB#e3?Z//3fHA(C/39
20.V/f.b2R#cUbSeZT14IE&W5RVU0,dZBJZTW-CN=09-JZA,YQaa\LBXSM8X&+bV
=FG9/2\WE-6Kfc8J>_O373MgY8V4XB+]>J0\,NaN1f&3I(9^G]@QVE,0_L(-O_(>
3I68C:ZPZB?SNOR&F[HP75(@4\FFMY@U)</M2PZe@46A1RZeC^LHcOR\2KXWMI&N
RP7d?])O88MY\VEPgMeOK#C/AcWHX>]IW(Q2V.WRO(>cPO1O+T?,MR+,9M&CW4,_
4>0@9c;Y4GSNQ6:GdLB)PUA_#Y^3Kc[NK2VYYPO-/\b5@#RdTV7ZZ;@7<f^K-&9R
1>5Q^4X.(TU(e@<UM7a[g,K;f=L-)bb/&Ob:Z[I?1]9IY#OSgM>P#PL7b45Z^.Of
+HebT73\)=+H)-UJ2NAE=]X1d)<K;EF9a#Zg\3<CJ(A7T:X;D#06C):0F0)&&G@&
Rf4cL3ge7O(e<U>&G4+UHKH[gHXQ,>A-=@O:L+=IE6dZ;a4@V#2:S);T2eEUL#4J
G-BNCCHTF<],RZ5R6:[J@:P2OE_IVSWYG60H)f<cHRDc.=d3]GUSRE#IZM7W?VeZ
,b#N2MS/(dKO.;#G?CHQ/fRO?8.C547YZf[1L_<Q9X[B?dP7e1AV_GUATT0g.;B=
?N4CMEVK^Ka\S9=2H=1V&f8T8gKPL05X?T9Q>BC?9YP76U)H>4J84K=V)/VF^KC?
G02;Y;7D_Q\FBXXX1bM0CF[TMdRD^@ceDc0>G=^LN<[Z1Z\\VJ4MW&M1a@]D6M_[
TZZ.03QcP+_YR._>T:VY@d#4]M;Z-dg:O@1^5[NJ4/g/KbK;FICP#4^JHG;JJ,A^
(O:cSL/QE,W1;3cA=b4,X65U4;b(\&=:HL\R@4_SN3-H1P)_JH1[@b167D=[fJF[
\]]<0RNSSTeG7N[OOKI#^X&Ub\?LA<ZUNP&X[UL##_L^S@#7AcWA<V/E=&0;L2@b
GLD9RJW]2TXYT?/LD9NFd.-&&P4c&b;KM3^(MXQH/bGA4H?->I(B2/[33AV?OV96
4/c8B7B++aJb+[P=b_215_X29:<8]K&97d8O>,E[3(0[bJQ6X2UI-+;f>5>WLMN0
8;MH/XM0dS8OW<C)15YE;1B_Ecb60e^N56g1DAHWV#4<Z)PUTYEdLZ1I[:)PW+GJ
,8671,:JH05^NDBS=PXe7LW/[FHBCf:OXRVfgZH6#;?HBf0F@Eb-V.@\#/4?Y/WU
79)P:dOMD#(L2K0?9O)2A7FK:<-DD+aXRQI9,,^R[>;BBCQHIU6[]Ua9BdY8+1<d
D5HedHBIAWH#Q+WQcd:VeNdV5N>.A;5HY)+Qd?4fcMP7LP(g[#M.^8IZGA=4fC2f
/]=6@;4VT9N.U1;ReI&ERfd.BDH>5baca;(K/EOeR0Y9aJ=bQ#>(/=6,)gODf5@,
]=G:[0WV,:>dMWJ,>c2J7VT@[f9@Q\<4/O>@+GMgSDTG7b=0E-@A3E_DJQ,O7<=^
)AUgWeH#;A/P4IU:&8]&AX3\YNaK;2.Q?dNdBL:3g+(c/<J3E^XLa331QfU3eQga
PaPZN;XK;GDCgHI9bLO@[D97Y1Eb.g.0,]6#_5AZ2I^Q9-(@T1^,124-N-6P[<9+
\<>X38R;(97]MfTCDZUC1J4X#0H\XC[/1^5TO,-g\2aQ@3fW2^aB^:K<V?A=A)f3
b6J,:@>.G:VDQ1bV_UALT(HZP];f?BYN6YNQ?\QI[CXH,TDWW^4ME+364_=Oc2(2
6.Jgcc5Y\=_\ceX7UC/]H@<PCLR-GXV::9.3?+-#.X2W4.)3NL(OC8IYc?C7(ZSB
Q8F@6.aJ45PdEAIPKH?35RTU-XKbHQZUFaH=?K->N)\7W(eE3T(H+LJ4?b@+0.[C
>QL4B)3KMOB-JIbF2U6g,gG@O?<VXDSc^3K\)ZR\;;dQL-GVKI6bEE)MAbN(8aTQ
5UNe&Rc[;=,Z)K<g)d-?Vb[&7XG8J/dJ#N]4-&[eg#UX1&>\cS5ge62D^V[<YFES
](gMU/].+7U:X8eKDARO4Dc5RK400;c&9GHC\VOUC:?&K8@=YO)6#=Q958443+-L
?V?fXJ3PNB7L@H8P6)PV?H3[+7(EFH1]?)2D_N0\DHScJNJ?MBSE.Rg(>Y+O:A(U
W+;P+S+_f5]g0/2.@aX+1.26CgXfRZ/@KW:/I:bZ)(+?@E>fB_70eI]D9ZD2,\7R
d:TBVY&K>MMEJ6@Q)L+M[5O_XH-dKee2_fE#K09HFD,+S(WS#UTCOSAY^12-VI8<
R1OPHGaFcYU,9a.HOTW5\Bf,FZa9b9]\2&=@_)>O7FPJdIP^ZDT6Ic/-;5d=D(_9
[O2gZS_\]TbZ</eW>Cd[:ZQ>]E)DC^&4H_dfXR3@&3fPA?:KfeO;]D-]>1+eKGYO
aWT]#/YN64]A.(]XQ652c:=bC=@NGJPNF+=<N3e:R3WQbN(H#0:7>)==-dPaOcH9
U02L;d1K5T_&F>8g_4[7DcH5L1NfPRN=KG963<1CY5Se&=.[fg@BfBXV(F#:c9C#
1[F<S&^KU&RfZB)g:If,<6c_;Eca7:IPe0_7F-ZK>^(X1X&R3_^#E(H0?TW=AFAa
H-S>3+U],_S.#ZI4Y(.S\gFJQI.K@B92e@@V93^,PQLa.^J/4N:D1WY&00P=G-;b
1@0[&DO3\(5D45&TAOD1c?V,9_NIIeMB;-:68BX5L:bG6TScE>6g<D^NI+_@ZPbU
<F4Y5N+/OZ>FQSQdP>DVO-G7@:&JQ;K4;geV?8g>KBd3R7eJ>PK5g0=f0T?90U2V
,3G-M70K)_G7&ZV6N-M?UTI;\d#L><fd&K<ObE]cSXbgG69;9,>gX9DdF75(Xf_:
]H,=fDQB4eWQ/C8b6O7<5-@P@&]S9QHe:KBb=J_F=CQM]+gfe-aX_EfBDg9W]KO.
&CBVIU2H;F,RdM@;]F?+KIbT\.6\FGa?F[6S<Xc)4?DX9T?e2K<[(DV+#U]3/[W^
^a[C76OX^_4754?FT-L9VW8PeW\R7/@_VR+<RSAP6T.J4^?2/Q6+8/ba]P-gXT<R
(?fO3T&P5A<\d=_-c/CI4VC51_AU)B;_326IZ;,ga36VfJ=C1]>VJI=>82D7EHOe
<>ER;P&(PJ+<K?gSWS65TaM]g.^]@EaObe,c)Q?HOEQ#TH&WS_caaA@eMT?(^6HD
BDee_^&c,59^A06Z?SL=34:^UgQ,dK:JZ/d]4T?\QLC6#YUc+;/22J5d^:N<>JLF
L+UHX5aRa/H>&2?cGDQRO=1PZ((,A#9/<(<b)Hc/M<Q@<>=52B\S[H/3VLO1b>C,
[E&8+JU14eXZ6^Y(@gDg_RWY\Ae&KEA>T79GAIa]ge3Cg;@O,^599:T;c6eWY/&f
6WTA_]NKU>#G;OGEI1GXIMcf7,(7(D7O(=1aeTfIeW<ca9S/<PPaAI#.\6(d:Z2@
@+LC#_7L#\V.N,^dY[7Kc<J?b5eQ_b3^fRf<a=00+I[#a##7BQ5NbE@QHZ7XILRE
9@2dD^&IRJWO<KJQ(4^3G-R+C-K(K;1>+/4V7BPY,=83YMC-aQUP:(cH,29V7@A4
#-:Ie[[#(H2]bWX03ebA)?/^K8X=WJ2GQd>V]R:&[_S)7V-,+TN_W_B[S.e&YGba
\C#bbdUC<C6TbQ1\;6_Ff(.fNJD4U=J#LTT_<SU6<X1GVB^(PU5^#8g_g=.AE4HJ
>PXRO\cF4M-_8MPZ.B+b(Oa@D;]XL,AU2_SBf=O89#dE-A+/=,L&/aKNO.^O)EOI
>fR.A^ZLcNVI+D1TAJC9)PI[QWO4L\6GeSc](Xf3MR9OF;C/_SUK\SEJ:&?M+bHS
c;g:=,9aU1+^b/)6N)0[0LNU<0H;5^ULFZ9=bB&D3]>g:Qe]f_b,GacD,3(L(R;M
IU7BU:Id\0JCEM<JSV-GWD]J>ERW306,5&a8,YFP>O(0LEP44gOgQeOLV(H&:^,]
=\L(P/PQNR.2D(c/7U9\OY>>bK>5RdKDJ[E=2WXG.69X.7.YAN33R_aN5_9JMOe_
\&W92TZJR#P[<F:Y#+<U-91gcgRNSB>=(([J]ND]UHP=<0cdeIVJ5&XV1^R=J[53
/\E0X8JYL1E^4/QJI+,Y3]R<;&HR.3gBN5O0c9+CT:]@RUBNOL-eaFc>?6e-gIUW
)R#I^>(OX)524Q^TK/J?.O32g4AOM^</?]95AW[F901P_FNRfWZ^C3Xe)P.YB>g2
eKTE#K)H471\gGYKJI\V.S[cSVULb)8L;BL@N^dA&^)Q4aEW9.d,UUf^fD9NR=#(
1GZe/2O0Ua9^J7J,-YPO-)BN=9TaOP)#]9&55JSgLNf1.@>^g]#c<UJ))<I,QQbO
&LgU]65@W(aK:I#OX&;B/L=]Z^OaWXY#AW?=Qf_9gS1;/.N-a[<A7dW2<.BX&JYg
UB+7cd6BfDED6(P[]a;44+A/?V(]J)J1d?4bAB\G]VUBC/3G2^fW=BEL]Z<#,Pb\
T:fIfQ6Y[S1[d[>\ZWVWYE?WcNFa?Z5G+)J+<HZ2_4L;d;<P-K<E>>fX[&WIL&=M
T,a7E:[PE/5<?dbRQJ5b2]]?0M7EJDLWU,AWK7,HR7Z>gY2ZdF@(,M2T+<9<3K85
N8?bFYaSTG+-@HY5dS5:W4WI<K6,]F&a)+0@WQ0(#JDGR-KAXLHc6OcU#>6ad:A#
[HEQCL2BJf=_-5V,(2Ba.1GL,ZH;2[J-f4E3g-gQ8LG\MfXZ&/^C-1QV_9P]LMBD
1H.#\OEBHXbR<[P7b,OX.#>D6(0C+e#DF?dLYS.6W-:^3?[=#C&=[a#(7MEZGAZ3
XM;4/Q&Fb7Eg3HFKG6V]fP=P]EW#OJ:HbIc9&Z)<F\<fa>7E-7WZH[9D<7U9S_#C
6P.5DA+bOKQd/X3C-NRfM_=)I/I9(<]J69E.cCbHV2;EAF_JOW[d)UF7<&=?0=7<
VU)8cVe0PZ2A7+0X+EG(\0g:<_N.BM&2G64f0X=T&dN?VQD;[]-UNB4Dc/fD[.O2
]@8V_N7FRdN)HU/6Yg5G<8BPe7(T/>\^Y,O(>SfDf-Y-F&7=g.a;?YYGRg&[?A;<
dU12WD_(g8e5)K(O2A8H6FY(aEGgQ,&S5cH(C-H^;La>e#6FHB=8:-2L5b9]SS,?
caEOD1M+fDRcY1_F.2,\YW/-QMZb/UK<U.S-LO[g1Q>>YSWV=QC^U=/,L.0/f;g1
6b)9<XU>N(3@_UHQ[KX9_JG-g]I+U^XWD1[T1P[bF+ee<g[163EE)ZIFM?P;d/UA
KCI:d&/)_R^dcM^3bRKM7d>[f;F:W4@B/6QO_K;:UaVCVIe4#6+RPKB;:g??^]C\
O[HVOGg45]#8d^IgJ\<@RH2,,T(DW/3c+R6WD#cET&W.^V,/Nb6@J+3CYU1B?5g&
)RB\?7bG?9be6^8Y+R]30<8D_SZ4)8<]?5JZ@2&fba&EW0[:=JGKYS349#3_d\PC
7c&Z7<>J(-[<[C<?e2;FT[g;XE9Q4M#fW>]0DCC^4<_/8aeV-f&PKJd2PS,G])]2
:5L,gBT7E6&]K@RD&TY7?6(7J]#G@>N(>(bM2Q;YeCf@Zff9G@+_I(Ka\U40gFQ>
&J180OXMU4GC:]V4(;RC#8BUU@aGg8J[-^[)(QVaF6T)(PReL14T?aIDU<1J)a4J
ZOaXJ:\3ILO_bC#<)2IDUQDDR,;<4QTdYMIcLCAORCX:Jdd.gQN7[/7NZ^GX_IJ<
X7N>M20PE?4GEKGH,M@)JI=a@Ba=0)SYA4:T2Ug_UUd?D/HEJ9SYeeZ]E1aY;:[4
Q:OX2?JRf(:0[,)1HdIN<A.NXfXGHMD1=-_:_gB;2/>BNQ2@.Ce47X_JF4HO_G-;
/P2HPZ=,ZB-RV_=efGRFTZ;@ZMRL;,O]fM7,7>-YY#?PIL(Ua/R+g,,2Y0YVI19]
gD9)AV4#5R^]D.T35=7fFO1?(_;._1-#0ZP:5d1#aBeUbV2E=4SE20:AI/&1FG4A
0UdN@?AL<BS]FN=<7ND-&LT3OGJUc+US/CQ(e<C]0e^b4a6GSg67C,^SA2?V86Q6
]R>-Y;UNFGT4<3dJ60LM/O?@U2GJQARdDX>#R;W?e]f6g^)MU==eM6c88CP-8&,e
>@UCD)^V#U#b8A3V;D)B-207JNgeN==,FNTb&/<WU@Z0__+X,1[Wc3UI.3(fYad0
I&H4RS:(PD_V53&W.e\;LPK3[PD\2)F.a__8VSS;IcT1,+BJ#?_<T6-Wa_KWAH2W
>?C<6IMRLQNF&51MQZF.YX9#ce:FSS:ZKbCFefc6]-NV3/9?)cLUc;.J]=,R__XI
&.NJ(LV<?Z?Pe51B1+,[3IVg1VELGPf6JN>/[.CZ/SSFGX3)^O4b1=KEQ]]8=3NK
CCeV]O-O:#aPBPI,^)\;@8#fP[3(bH]F98I?1Q=+gW3/b^^F1OBH+](4WA2.E-B,
B^_c)7@PD:=/824+8@PH(PAbA&O[c?86I.+5.JHLG:7Bf._\NX^/UUB;P/R/E@(&
\>SPf9=YCGF-)bS53Z]E3CIL0LgBO3_Y/+c:X#L;1Y_E8,,96cC4IL7G,e=>JY-[
eYeA2gL9;Y]2]DYW;AC?fIU6a9;#\0?(a:G@H_]1G5F1:R:6aR>e\NP]aE?K06dH
W7aa#D.C(>U[VBg4e#L@<UbV&f+U=#;))X06AAZ&Ib(5-ZCfg=KSUZ3L-A7ZLT[[
LFOf^afD/HVJPLEP#\=]G(@]eGf6Z;d6(?b#f^Fc(XEOVK3#\P;O5P(.]>NMS0Yc
#068HdZH:=3VA[?f+#](2G0?L[-78<W1COO[MS5a8(6(6]L^=N4RUA6CHDe05b.R
(D_fO5N/Jb+@]&5?K-U;_FcRO8NJM,ZN?@1ed+LP:fCT673+4UB4C^2]#BT,5SeM
+M2GMHZI-)MW)S?W5WJY,DQUVGe5O7_22QY7WMfV4BJ1\N_8S_eFK](&&)dLPC)4
U)ILQ1\FA)<Sf&IMC9&4=V8CQQ+d@ZfF:3_ZYfa6&M77U2ObHG86E8Fe]R:OQ)N4
GKeZFS)F-2(#JcQ9=JD^9YaE)/(#?KW2f/[7S?(+:8SOV-TScOg&U6RGHZS-TT/Q
@RS^D2CbT@b0J_7QO[F-e6&^4>CaQSCF58_D.LbL8dY>T#V83ZCS.cfZ?N(UDbP=
eD.3\#Fdg,-6Yg+@RJ#T<e-<_?[.Y:PY>[LBH5F,T<&&.F4IE=/S=J#@C4L.3T].
/bOHQcc\UD/1<4OZ0N>,g,bgI;>XGa9N:>)eF94\F[26Fg7[Fd^X81.DIYUbY9O6
(2A#W1#\6L.H<8Q(8#<_J=c.aYaQ#4bYD<.B&@PNKbbZNX2E_NDg):NWda\\C:R6
Z@,)2]<P+AOD?6ac/<SgO9W^FW]F,#)H0,KN^;7YA1H^O:eA,cJ,>8735JE.-8HR
#?FTF4J>4EB?[J#=R,#dP;aMGO,<XZTZb,(.cZbg1UM#Lb2aBe(MR353?Ce>B1MD
\);&QYfNA=e_<3RNR0SI6CZgOD5F=Y0T.Hd^gU,R1NCKDI^4=.OJ:[AR+EUUNc&+
>B4W797Kf21;<X3cY<X;ECR0FEc48O;^4M<J=d5.dN^@[>eggdY(N>Q47f8G/0;)
.7eY^f@,I:;GR3(P[ARR]()1[#E17^H8bbUL7^Egcd=P^JBB,.;(Y^4?0^9Q4;(3
-cJ8L&#U0?R/_UQ1F8g8MC3NRL]0)&eJRW75O/dN(I5#Y/SUc)74f7:^f@8D+e8R
YK.<:N)NHVGZTW:YUHP+FW>+P.@.^#-ab3GB[2ZABNcGD&,3H1P77=W\Q2a9e<4G
-KcC7<X_UR\1D_cED@DJgE:fFd7S,(c5@DCY@.C1EaWH.#J\<[S(:+PQ]@,5&IL5
Ue\dAGROee2EP^K5R(J<X?MU2(AV==,1Z)B9]f(VgdV)H8d&QdfTM7.GC.?XUFf6
8=/9MX,7;VRNYKfS<IT?0@&-VGO4=G<03:\H;QD/5]\U;TCW9gDaaP&0e]SEf:RT
W<=U?>4)QJP7<-:c7:487#,bN+eb0WMYYLA+:E_I)2;Mb_;Y]+HAEB?/23F=a6<?
6U5>)R+EaBRL1>OAV6X3g0J-RJa1c4,O5US59[B0R,EI#HE3.f&&W6aPeYPXTQCd
KSTe@cH\5D-^:0EIO&Z0(0W7/4W7PL5=OS2E3MIL@6VeU-X4R6.]YZ2./R,0C\44
6WPd=KY3P&GX7BeRK<Q8DGNXM:B;a[a51:IH<ff.N(D@W616W=?HJ,G+I/E0E(>+
c(&\gO]8A8^D@,B]c@:K&46@6.6MK\0&J0KI(;R&+^cC1eGAXQZdZ08SAL6@]2:,
):]WV[&7,FVVC@KW7BaUL+;RPHYc(>R6P(S.VJVK<-G@L3K0^<O3b^Kc@8E6@8fT
28_H1(N[R&4M/4&9&,1M(\KW6d>?HH:-4,]F]:U^0>P1]V:NH-Vbd8<VKEZH<0aH
37XbJ0J&cNfPD,]C82E5/3JcJgPfR&(fg/U21S4I4^9&[ARLM+c5I4gHLV/>#gg)
N:dGF3UM:R=61^LL)g#=RCc?)]TNL3>S+MBV@<)=AeFJ2^)ZL>-GCIZX?Vd(?6RK
MFMQ;67TJC53N3R<U>ZN_e06H8(L^J1@9&?2:7Ib:T84Y]>5YX+a]^40+;1FBCfC
)->I_a<a0c9Dg.O0dDfPU+GU6MBTM(<QJ0S\V=Wc>9)G6_[7SNDK.M,O@2>#.?C[
7B,:V[Xe:EEK=92TC-\+&afM&MJ(5Ja])F7\[-2)dOOES567TM/.&:.;1=T)U>DQ
=4A5(=X_GO^\>FH/P\?=R3DXbY584&,77J[&W4SLL:1)_8QRZ0UPH>Q&aPHU28U.
cDSI+7_O4]##1&F><IRZYS^fRYJg8/=>O7REIXYLbM&fT_Fgb7##7\&6T.:D//Vc
X8:eQPCeT,+]-\>N(SB3LND5J)[\1>f[_Hb1Y8A&X6?>D?J.C+GQK#LO18K3aC/6
F06U5WM]1MC-Yee+YH45d7bMSd.;TDgT-AP(Of#W/b<8C[U\&#RR^\K=(Q\.a]]I
VaSY<3T58G[,@&8Y_RUS5af0REBBcXG[.)M>9ZQ^(&OGT-IDLeK)e-(FS[G34QHZ
W\=D08bJLBH>;O4?TEA_&@2.1K(DK0_FV<b[),?g:]8bVMG;gV]QK/;G]gaA?,0X
b^UZ)&-KPScdAgBJ47R/09P=^J?(M;E)A4X.<[&^EO5\:VccdN<J&:Ze.S,MNC[B
:d(acEONYE:#\49S[MPU=@d9^NUAS\KPUdT4OF3<KLS9P7-_-gJEYBQAP58e(Kag
Q.,fE4\U4(>L&M]6&8J]<I-cJYK6TL)S)N9IG^L?F=<+BPbL2&=/3SZTU>KZZ,TU
a6\?3#b\HWER&f@LP0/PU@N2-T8,F(/)]+cPTVZ0:@FT9U^3e//O6S6SMbK=[Bd5
)TdVQZC/,BK<Wb30X;H^A,.1>J)O,d1N.B4RF>K:P4TbgR\1^1F_e,.C54]9:V4I
#RY^B_2M9P3?,#T5Y60M/AP?\]CP?O=(-S\?DXV0\3AMFY[S3)4VND8NY=T4O]6V
1?bd_-K#L+aR3.Y^Y@(A5]_8X.CaW^<ROSNN[GMC.gK>PJ2Z=:1._&#Xd&g6fXd+
B3RS1M9^5@#]Yg.=YGRg1W8XBF_OP)G:/VCe8^.ad<Xd)K@;?_>ZcG<_#e(5>N\E
PKX_Wf6888&PJ-5#G7bA],\9J7H-Z+?8.V5.d?)cZI<CC\F#:>\/UO9.FU7&,b/=
P^Ed1?Y&1b@P;+V#2KL7G@(@D(4d>27>_J(K]HG5=I&UE1VA;X]0edK(JJH<RKH#
1OW,WcRHQYH@^D[f>YED#eV@S6BP8M<E9)R\dS=.?CZA-2=SROKR@KY=.NH[@D5M
+C[8Vd[@11ERaG+-MBdKg54dOD7_XO>XMe<F#.T[gOgQ</U1N;UFC][abTd4+_BF
&B+P,TFbLZ29;fP,S>YW0JFRGA+NT>R^9FPX:B006)e_U[FWNg\TOIB2#PB+4VU3
2Y<S,#GF(W0F<=1D;=AU[S0[PI8F6B6QNQ;8YEA_TH0,X+UF)YBK+[U=G)8AfS<=
D,/FO1\2@S46+VC2,@27Z5U\OFgUf8TB83:R@&[G;^Q5Z7ZO3_>1?2I9c;QfH7N8
=fQG4JXf&eF[JLaaXc_>Z=e#aGDc6)cOLMZ6D576#.GD95>aPP.4bNNHa;_>#\<D
H0D[CE5P?M&Z_ZY6+fIQGT__]F8/[Z5VR1Q0f0>+O6Gd#TIQJU.0D.0,Q=YH4UI(
4E6@YKd/35PD?O<bK/9&Z:3\&S:0->@_@491+(O26IT]fWBJ]KMcBd?X>\6\,1,;
3[86,RRd700/O.TV(G?fP=+#f_B&f5KdT6XUeb.faEP1A2/&UEAF4d=4]DR1Mf+T
abIbf2<9(A5:P=1:_8fc=UK(CBXf4]N40XN?(&^6T6d3F0eCOB4GJ?d\T;FC>GY6
#6,d:?VeN=+fSGDS@QJEbQG1HUVL/b:_YQ\g5[Ae+@8O[0]+I9B5/;+:1,K>[&=.
HQ8b&Z36)HaP4;4YUf_R804SPT&g2LUDJ.:Q&@X+6W,@Jc)gK.F)1&#Ig/?;W&LH
PD?]P>LJO47#cdP36DNI8R9bNVXF.5(<Y\a.2#4EN>dN,JX;AWKHOaS3>DYbTbA1
F+CfBa^\Of-G.=BBK=6CBMD3bIAU?>Z_0cB;>1R+NNJGC;T;,GgG\L]AX?#RDF<a
?IFW55M<RNGFHO4GAUX,3950N.;3?1[UX7be&5HZ5S=I1dG5G/ab?/B\.&PYL@^U
>^[=F7[?<g)ERDed]\IB9d630;1H(8KJG21JS[E:&SQSK(R##c7=Ob_9_LX-9(UN
;1O]?Me[IR;@<0;BCKR53JZdSIXOPRYRcf0f<gP9)1/VJSC3d&>Qe:cdJd2=f,18
K1O_Q;b8/,T8KLN4Pg+/P\fd=Dd2V:Gf-?)S0:->[+d/7SJRU<Gfc-gO]P_]<MN7
,MMXHOCHV(XR4aFXE_MT\L,.GdQ;B@^551G0F=D?05IWf2O#2]>9]12V\-DO6;]d
bC_DB:AL#X8Q^,Cb65YNB.g/a)12gQ95\CS\L7PC=e9I3[e@0aM7YE_=VP?O<9\-
Af&1aC4)I:AS/(TTOWN(]IDa?5@(BJKVJfASL69.)#8&]&IXNA0RK=W#@]Zd0KQC
T/<S/H]^^EY]gd;Z-KR,;)6H#D-]80(=N4bZ)?bX#6LIgKKCFQ6gWWEccH&PLK8Y
;JcA8\R66RH#bBd7[RRN+RYaL5f89:9/g?9KSBY0BN-7B)>1_4OU<=<EHZY\\9X_
D^I9?&>C4Z/PX@ISQI8-@;[20c&T27aeZ32KT-#<&N+E/O+G]J8;8DL.(N[PJ+3X
\Mb]^A<N;,f,JMEAQDeVS3^gX>ZNGgT<Rb+BU[?;X\]:8PX4Cc^TUacVQR&;#PF7
d?69P>7XBBgF2_N^9fLI1NDUL\1RY5^d65aPV<.&150@9V@\;CB_GX1T<F[WNY?>
UJA@Bfg/ZIR/]Z#T(X-fGBb18.)&F>1,YT)YRN>ZDa<T38DYXA6\6TUTUMEJORB<
US=LNXUY8??C@?]_11JQ@7a7&,J(ZT@E6>c[[Qf1T2_LK\,dE//5K+7FQDLS^R@D
eSa(C<b&P[ME&&/31c_JI-^X6I-G7U+N@]=_;B3X/4U/RdXPac.HMOfQZfOAT2I4
]C)Nb6-,9I33E:U#I]VIbBVCAeS,SL+BfUHe?.b285V[58d,+.Ga)NcZ6.fQdd#Z
RG6Bd:R9]d0d-;&;+ONCQ2aC<C)_Y/E;..[.43]3O)[1Kb-BIQX=Kb<PZT7fe41c
H&^OY7WQJ1g&c)FTY7HfD?@OJ0_f?+ZK&\fX^AVf8_X=J5)LK:[X\L^;]cRa5UD7
;f..U8bG,eEM#2Qe=7L;ed]eR^>S#BC-d_f0C:>FVcYc+/Zd#XH7U7]B]Ze70R5B
=cR]B[GGD>1?gJ+fKYeYDHX38:g?T?P@0R@VQfbU;NJ(:-aOUaW#0.L<g/Q9eRKE
2&UXg)CF7.V<Jd3;/J=,6+S=;Z/.U46A:<U3?RBZ4K6Lg8ZK#M6=1Z3[4@T_S/A.
+7gZ=U)#E;FQXf.J/++Fd:RKD3#:+#b46YgN)BX-]&O4fC8W#-)K(NKA7,PEC((Q
NB74-@NV4SaGH=@A_AK#B=Y^G<UePXM?dF6<=.^IEG_1/2<EHObG#SBNRad8OKTf
OK?@e+@65C,TFM=/Q?0W9(=B2IfKS;8_4\L,cDU_B]<-Z_&R(60A+<cG8YP_=K8c
0,3H:@--[(CY1&+KQ;,#-0&<eQMQdeX4Dae>RO[?B2+7MT=O4C>=XO/^R5@P(7:F
6TL=T[F8aC)FHa1_3P;LG8OT=^03TcPD)L8PVO)D^N>KLMNbN=gS3UbgBL.@F>E[
6A]NM+CL[GY:LIIK08:TT.11?XfY>KN=+MJJ4c8Da82a^AFgQ:2g<-g7_6&3URN8
XTUaA/GS>4:a[cOEF]]>I<@B1]I>YP,@T5^7.AL^Bc9R[QU>&=&Z6PQID(aE(-.b
/M/16g#]VIZ[]R>_R;:N6Ha<aZ.A?DZccHG+MPC()ML6MS9,[09O,CHd/ObT]@V_
9bRDK&KRZO#Ga#C7[,dBgg9MSN#;4O=E4/eBF06SMLA@+Q,gQN(0;gHS)3K&WCRZ
0#\0]>:T#EZ<>DPDZ5^_T:K\U;&;MRUQ]<R#HRR4cdd8)LJdB3=.M[-1AQ=5^3@X
]N9KY:NV9O^\KC)+#HXT2UVJLHUBHK>^S)RW/aKA9eJ0Y_N&#(7fV<TM=.V>FU8.
).1Kgf>NObKe-e?Q32#44\<GS4)IC&;S<f+.SRa1@FFdARNP9N8fXUR[6gO<7V\X
YYH4&&\-M4-H1L[N[8IK3CK]c+Ne3a2HI@DG:-C-.Z6.QLc[M,+1Q1UOH/[T7[CS
7WZ8)]6gJ<f/QKYT[bA]TZ->N:]C:KY@\OPR,(P)?..WP(65IC5F-=?U;2N6KLM=
W48PYGB7@@E0[BJETW>;6cG#I9A[<KeK-\.Q6Y^aSHNJ+@559-ER/[HZgR8G:af:
aC38.3(@EV1)0OP\PVQJ.10\C7SW/,)L>?4T(3PZ_OZ\(+I^FLQNE=JC\VP\,BZ2
eGLU:;9G(BF?;H4X[a00ID(9-B1^],:A4;R+X4MKea/^0ba](PJeW(M]]#1fA&SF
58Y0QgV8TLUL3G&\5\G)DD+-BB96SD1AK+(E5]HID,J3OCD1B]Y<6a>G0.RK):D0
>(1RYH>L./>838WPIS-U963b9b1CB:7YY;Q^EH(<<8?IMFA>9:<PI<ZU:9(HSEZ7
LH?/Z\;;.#UNQeVMNd<RbEbUJEdK1,=gVRb&FL\\T^ASB(-^9S;Ne[.d3;fe#7c;
a01d2XKIZ.DQc@KD09(16\;T/;V&TgG^BR9B.gRLdXM/W80^Q9HGY8MOFEPH\M?f
W]D/).GPAIHUWBFA/dYCA4]W&E5-R(ZO):?4QR&0>[BP=Eb6(Z,SN:9JMW^W5b(_
,5f8_F3Y+TKAFeF?OA&)YBMV9Da13agX9&A&D4\YVU(VSG]g^f6JGLBEcJf#QF^(
>Ca]bZRYR@R]MIF&@;RHKYQS6HV:dK:8ITBHHUaNZV.+RYEJ3bF^PXBMIf([JcD1
D^^F396.#783(=/;T;J#BRN07P#aF[BML.<32>@2V)/)a\PNH^5<F[TI^FG&@>EJ
CDU(,9[R-?W9bC#?@+_3g#6d-=C8;#Kf.NVVa<+I@gE]37/VKYe52A@FPZ[,:EYA
I=B#,b4eX@8?=g^F9C[7U7PdFSF3P#JX4<gT.NFT+#@>Y^+)?Kf.7.A+BXGe1RT)
5;fb.WW:H=2(>=)fdH_QAc,A^>+a/Q3/&Q#U41WLSZ9N_704d2K25HJ.b,W0_S27
H_?\Ta_8Sf:KfegdY=?1T_EFVf5Va958E0UO8_2#E1@<F27KNbaSBGH1J)ZLH4[V
GEIJ(?L6(1UaUc<./F;PY,JKTY_?(1K;Z;@HKb6F<R_SYbV[Ee_^/eK_Z4aVX;^F
,gHeYFcK3V]bSH.P82gQ0K3IGIMCcMXG)2[:]QEH_9K=Z:[#5,aZD2V>5DF(T0#f
ZX?FD7/>3A+=Q\H#>CYO.0@LeS)(<fX9-:H#D7e6__TD&-#c,LH@gQA=X.G^8,#-
gXbBc;@d+:?Z_0Rfb_^;@P&]S^N?T?03\PeH\WR3M845IQ;<R;(a3dU)@.04&N=2
=Ce,Le#_A3-:9>ULME]EQ^/P&+,\H81J;+7?)X-gY7b6>5gQOKAUHT:Q=FeeO)71
[#/BA]=[=eL1:HPW<V<6c(=U@F+PHc^@A;E&[2RN1+.E5@6,@4P3XWc_Q_(JJNX>
d?0OEEaf?8XA,I_#\9K(;V\S<N;8I=gR[@AH_6FJQW6SO]N63=I&E=GTB_\_K9/(
9Z5K-F(gK<UJeC-?Y.6eZ@Yed_#Gd6DgVB3S0>LLUJJ0PG;4SR#G//)XI@R1DA\0
3GC=6^39.g&Y]S&DTK76C^&-,E/O;=A(<.YL?0#e1JVdDPM&HLE;f,>YHVAb7[I)
:^RU_R(ILX+]Z^F9/J\D];-,FUCGYUCJX(S?C?+WX;MS2dd33[JUW)>3)\Mea3?)
#_>;]?f>J5T7=,UYf2<Q^Y>f&\/eD5EQF&B;6aW/Z\_(]:ZWRZ,VNZ,.+__8;caO
CcIe-C&^0b@SH:ZA^f^0-X0QV:8N>G16[561)S[-\_50XJafN0LV=-BW<9D8P:>B
6TS29.aQ;D,?8aRT)G_W<;AId5+Q#4>RD.]ZQH16SKZ8YWCP:dH,7K_-bAOe/FS[
=YF[YMAC>,XQVVNEa;aFL-7&939YfL+O#E1^-WBIAcgcSB^L26BX[H;#BOb3UY#K
FL?gK)PJY-)M/D-7^g1[=_PL+K-+_?.5edcPGX=+0HJY4;dac([BS#OYS)P8+M@&
W#.H0XV^(=2I.O]/)W:IAf#,;&A]RAJ,RPD7I@X>QYKb90/7E#3?bg=;A1DM/MWe
,g44X2PPg)f1\1(>RKL;UK<6T5@bC<\CG+-M?dYE?9:YQ:.HJ.E7&+bJY7Y0])&2
d>CGWcd#C53:Y&/ENT[3X+;gX)Y;,HI5WCg_GB3eAU.J2JWeQbAJbM3bPdd,GdW?
)QfcSKAVXS9^;AcB.690\&NP,9be/AcaYCW<dGbJS-\[.f=NP&Q2T5&./_+9ECaD
:&^KT?)Z_LEJGY:+<&eWf28>f=SA\/c_/aEDAD70^_2JagJe/9EBc_a<eSL\38&=
b)T;A4.3[Z],5>=,Ma6W];+A8E:-(,[YYAP7ELa#1:FRW)QV?7ACYF6b\/-J/=YU
;^]<:-N1e2>DTYD[A;_D2cV?D@JAJ2EI..\&?[+(JDg]+Of9gOA0Ibe52IWOaVV/
Ie;;cIf].^,(a#>I@Y>).F#(2>]VX=N0/=868VGP]VNMFC#ac,4076fb<OU0XV4D
/K>g(+^ICI_VaP;#]L+Q7(/UXA@;7NG47cS[O]a&2AO?>6<K?VB0Ye378>fNcG_-
8dAGa9Z=f-L<R4YXQ57@?7QaWYH@&LOOF;=CSfHV6;?L;fTbPJSDVBIB^.407+6,
^Hd,NWOJ,C)LJ9L.<fX_4N4O-A8BUA0:fMeRZC?E.39a?Zd_SOWQ:1\^5#V/[HQW
?55&VS25&UW2=DDA+Q?527D(fM1>,cfCWfJ.Ig(9I69UKgX.,9392&\9)cHc[M<1
2PQ+D1]MR6@F6DD_LGfF1.bffQ\fQ)H)\W;/O6N&C@M]4NLB_R1G-@G87aENbSN8
]G_V9JMYR\5_TJ;34.g/R[P@cNL[=ScV>6MJ.5@/N=69OT7]U?4-FGgIA7UHP9BP
(^b]X(b6Deca\17[(5F8G&d,?IJ@MUddTPYdH52P)6fGHA8,Ta1X@UA@2.<-cE?Z
&_\;I4/]_?a8@H;)cISaNAR4>/1D90&[dJAfA-d(J8K+^(;6HR.XGX?HeVL)5Q[=
2O7#5:E[J)]#&>fH7J@,Md/A1>\,D_B(HSd__f&>DK/R_cC]U;AJEWJU<S:Z<_0K
]MS;S7+Q<@M8=g8N_78?\EM;L25(_C17-FLZ2>\;/eAJ9E1E[2(TF,H83Q@ZODX=
a\LGLC@=J?\V2:F_ZH06?R\ZS[U(?d]S^/-#,A/H;Ha++?;V2d<O1@Y[P:GQ>+S;
+a>N)+9TB)agdA?L[J\OT^FM:6Pb:78:^:A[IKeNfdRMES>RY#HI#]3Zd,VD:9AV
&A45N&B6]#\VY1)b^BXHJ[0[GR3M:WYYQaP,N,#7HUWdAM88GMMDX38#F17WSSIZ
L/6D]EGV>UV;C1>+F+:UQAB)^BFZA9)SWKT^2.XddRKB)M;-fd&gA6CGP)-<-_5B
Z@:IRfcDHdIN,NDeA^?;b_Z#-)-D,U0#[C(&IQgO0ZFXQ/TbdR7&HYKBZY:Y^Z[a
Dg.0MM^ALD3_-)PQ@31?EY->HPS35eT[I-KQ8-W3K0/DC4)+K3W7UJ7^F9Eb]Fa?
egdf8UF8a-##1c+T(Z.55NA10;f.+O<IR.g;+;N[fX)aK^9NF7eX&UQRdU+\I)KZ
N[U(6J[R&A0BQ19CDDQO<_&;a@/JL@E;JI1ZB:Z9FUES07DIgP7&L[)f2SD:9#VR
[:85?UC.PNOT]IXQCf_c+-g21):K3-F[\8RTU#JT[][N3FY=BQA,F@[VHdMQ2@6S
VD:2\?.61>)b(2RI3@<5(1D;aK(QK>E62UL[-SDd57?5e,<ADg,UVI(A1>+L13dB
D8]TV&9#?C:g496:aU59+Y6<F[TbJJOB0<fa,Pe?E4H2dQ,\_.YOaX5DHSNU6=C\
gF,I,-9;aEW=FM4^U[feB)fX(WD--(YIQX;.A]19NB&P?&g-IYDXBY?DS1eKHD?;
.XT2+bG6SZM7[[DQLX5=H\7?XRC?)fgYbeba54RGU\856:N_RdU8BT]-GB.G.MGG
=B,]IE5>[c3_RF/3F+B5>+9d1H#d<5g#7PFHN..f1L.dD.VIV3\Q6Q4&d@,5]gc2
9M<cN62\/>FGggFO1\a[1^_T,Q^@H(CDc&M3/7H=PWT_3;#D@:XIO@Q]JGf^)17^
#B3+gS-5^X-gMfI8cc3)4DbAK[2R,O9eOB3.Ze.Gb@&:P6SI(<\7Hac91&,(E2)/
&V3(.S3AP+W9YKYUUHEPW8:F(cAPed(KPA,8aZJ-ad.ZBC,d3F=d[g1?b5RNgF5f
JS7L7]Zg>?]?F.>GJ,6a763adDYP\KC-=A]aae.L5e;F;FM=^@O^b;:BMWYT@<7M
YGV=#FH=FAeRgb)UJEPB_8^C,C>)g7?^fBSZaLXU2E(2[_])=43[@@OQdH<@gBG9
c&@>M0+^<KaP.\)Qg@5gH3TfP4E>]_&WYH>:/dgB,TaJ]81GVXK]:K8V\c#TU[6S
37Xf4I26X/,ae4>4#a6SM4f-X.aG4.@@6AC=]-DfP,-;0]60L>9P4Lg4]>6M43M)
KfET\;WY4c+]<J+;,efee>Z?1\3W;fYQ<e?d4M6JJUUND5TJE>WH5\dg[G^W,,B@
+S2XU-T17R5]CH_<9C@Ha98->-&AC=_<(^c,#ESQ=dYQZ<DXAYgLPLZW>F&:49/T
g5:W+OCeb;I5EGU>\=3<6)LIc:/8U5ccR9ed^R#fHZNeY5W&<1R\GM9^5&N:dKYC
.Ke+RJW<MR-_H4T#4e>La0V2gbV#VV;7b)eUWdR9WGWdOT.5Y1)_(<Q-aO8BJaYP
@12B\VL,5/(f2[_TddgF-C>7LO.g2+@3N/Y=(CZE7M=M/TGfYBQUb2#XA/FJ,U@X
c1a>Z,/d+DFQQS=(gQY=F#P8-/aC&fCVF3V6SIR[1U\a1_M]4M0@Q87.DJgAM_7[
,?\5FDRedXcQ.\J)SED/]a3TQWPRECdI_X<ObAB:.]\b@G]Y3b<NeG=#9cV&6DF:
d)R<#D<DaRT2196dU)_)0bUbg4J0C;=KA;BYH]cSNKNJS06cN>),16-#c,eH2Id.
A)744c8W&@^FR#>;]5@UT3T/E+E_[28:d[1BeaaM&FD@\X3+d=-;]D6J5Z<;;IRd
D1d3P:(.B_4+=QMK,dBdB]?>1@TM-Ua>E]?T(Dbc7@=/.&QG#=/QU]G(W58F6T-4
R///]f+H_,:GLa_P?Z,/)4H,ZDL+#@KRgFgZU[&ZQ0dJ6PW(:1L:GGNVR;X.H.da
=fJOS^6BIO=EO?58=7+:+Y9Bb>XK\dOIa+0WM;[_8H[J(Td1<88L+E<K7c=DEd-(
75:G30TW8=IKF2H60:;NTDg2WK,K26&D62RCLK\N^bTBAZdY#D4@]DdIA@N9395^
J-M>:Ag^f#@D&bS\6U8Y#6F96FB6M>M4/M=F#=EX+[:RD,X-U7e4HY+99C,J=J@@
BaL^;<9LaQ1/7A&<AMZ-Q8K?Z\P00<D#N:L\9b,7a[4^;&.(UK==^g@T9cg@3=<&
^3O[?0_.5Z[VJ\bX=TJJY.e9(^U]@1IF_]=5?[+/g1NFXb:L32ON6R=65+cSGDL_
d#_DdG>.SN9?&/Y5+e:^I_-fe^)+F,R\1[E](.eL)d-N24EXUQ4.7/R2;Wa9d-Nd
NgMd#+I=6?[IUL[P_A_KgDFL2B</FC[e:CD:@5L\^Q)X>B?1EKACBc8g0+d(C;,H
9/311Hga/M(L2XM1XZH2&]B+6T3JZ>=2&K@Z)<AX_IBD_BM8,D3#P5#cDH8@b5cI
d6:gR@:FJKNG77UFR3#DfEFcG^N<O.+c&97OSY#)H;>8U-T)e[8_c=1,-E8+#d[O
<)H4]f.F1@^JF7WaC.#]aA?9Ba(7#652f8IJc@\F2.6SH]GU#-#WYg_QB,V^HB\J
7+(SMC\@WV1WE_eB65;[2H)C+0-K#O1:f5MTUf-4&A/0P;Q@Ob)/+:&56XCQb\Id
G;+ML2f)]QU+\_E>#bTL>d.I86\O<#S27@39\,NF#75A_:UT9]?TDDS&XgJfD=.B
?P<dP<,S6@9S[W-;B#/F?c//@PU;Z]aRGD32-6OY9(Z/K3ASD40_#NJT&=c?.#G5
;3UNS,d;;<2#gLAO1>e_I&aaGP/33PLcdI=-ge2AG;Geg(cS\A(,gL>.+Q?#YFG<
V(a\JM0b.>M.L.D)Q1e4[Xc<YEM6-abe(<8T19ZD_-YJV4E6AE+NS^,.=dVXX^-(
/gKbfRW6Q<DS;[)dEg&N088_BAaJJMg.?]C(NgJ6cY0HYYS<67>KcR_,6L[40<;#
W8Q&:_Q)<UO4bK;J=_GRU&=9ZD\H+SQeEWd>6W4aYL#5WKJR3P/UGSd^_L2X\<M+
6eZ0O&C,,dY#=CO?T1Je\8:e#e;X-O?,H23@4?,FP#?\g.<)TNe_PF5>(DYL>R<U
aQF5861GAP[]9N2J><<C_NH&7/<Mb8TDT58Ac)<OHe4?7/<(cZfFI9[_H?3<0^:L
f4NWFZ79&M:AM[d]NDS\HE:N?Y>:[J<4:5/#;3NL46>5S6fP9b=1QS?JB&DWZgIa
/J8^>SXQ]WF[MG^[3R]?<=]H+.?MVR<)U^YN6+92Q7;#^TUJ\45DQW\d5GBc],=>
,44ea94@S;V3C?X=L1Q>B^J5T?]T08I<ZPR?_4P9&b@N7&KT?NP#8,\?XD1cZ<W6
H-YU#56Y>?&A^U&R.3-bYJOHb=JL0#J)KK_ZCZQA81ACSW_XP@YEa[XF@E]U-Ld\
P[EHGE?.V\U[+,UG8;KF2d+]_D,.e^J#8=_&Ta:dEN??X&C#J<2//\d3b-,]P?/C
&)M6.L>68c^X-U@S<@XR#?,,IORJTCT0WDDO,=-+8,]Hf:d0\+PV1=0/93OD/Q7c
:X>Sa87B=gd(#ae=]Z..?fLNK9;e[f\75DDU=-ZZ\aSC6W3F,B>5_GO&T0RL8b8)
BUR-.FXT&FgKa43P:cQ#f68T+6(d]0H]?#F#eFVSK.J/cP,Q-85&?>eA>W/_JR1g
9aO@([>D0-NKfOIJ6=ZAG&XS)(>V\=f+b275S]/ZVZ@Y1_IbM<3\;IgVgdR+Pe^I
ZEST:<.9.ZWR@;QES?A3E\+3?<QDSbPeC#F60-^e/\5DKJgOTUNRa0__6W_2<^gV
3)]HgAG0FJ6?9+P^.VO#D.78D>K3Ma01ZSg3QH#8&X&JG=&.OLF5\gQDCA9c@AHT
=\b]d)@;4VHR/V&-c7eYQfY90W\475SPCKI6ZZ2=W.4Md,@UHL5M?6,cC#)\K[a8
^DU0^Zae9\=7KDO:W-9b+>#0LAJfZ^BgZG215O&)HTJ9DL8I8c,L[S1fP^>0f3+F
D))ZT4:X#77@KU2,gG5<GaHESK?-fOg.Y(X:6c[R@1(+\VWE7AWba7M[+8B#;aZR
6W0D\4?D6YSf4PS=/fY^;If]3bTEH<<]YO.[.f^8K[,/2=3CIRKD=7R?32f2B2(K
J]>>P6GddI1^(dC:#F6F&e&QDZAfI=YM[aAS?/MDLT:X&=5[?aC@2K_HJ3)1E\;@
UOE/7U-Q>JcFdCO0SX0GHUX(<P5DK,WB2e;@S;5@M#UVGJ[99G,L;#/-^LR0F0eC
N/,0aJe5-=d=X;:C(+AH?VR>)ARPE1V.R)C#^B)fG2e?5dA/8M-[ZMcR]J.;OXT2
A<?&PgN,,D+#W1<J7,@>+Bf;WF9.W9d(L67D;b05&MHWR:d8X\],,+(XbDD7L4Ye
:HdN&/TF5HDNEN5Q\9R0J^)4B?Od#V_WXJEXf58Z7CC[<);T_B8>H<=@_DLVG?9C
fLf+FQgb;)-R0CGA;Q7.@C^2c5S-4,H#IK&<EGHM.Sb^V5<<C\B._ZNZON-c4Z=?
5&8XMEF68K7@a[S-J4c[6f]-HJA<,IQ#5<-e/15^Y,F>gC7?bbVeR[VILdSNT>21
N]-dMY)&I.9[[G2_<,@Wgc^4TcM6JY<+g>54X1dbEHJU#8JC24_M6a2+,ZFERRcI
M51OC\^F8Wgg+D:&#cAbDAQA].VTcBS^MbU&B6K;dSLg/U+1fg+K9fPe]=KRQP8S
;YDdX?W0D7X:6:(;ae3?.>VedK22PU41?QQSERU)e/dHN;YIB##G#BcECC>/:=LI
VSZX)cN(S^)JSP?NXd_=\D?NVV+/NOTD,)W?C<92O+ZB=OSXL3A5WUK:cgg@;T<+
[L(.P&0J5R-A9:1MG>@&<&\DZ2.W].#CO#]Y-ZB;EUQ+0.:CAT&DZNW+YCWUQ#fd
#:[=02=:@+K(-V1X8G#^YE=,8-eJ:?J@0g>?LPfYH8[7>_462K9Q=V#/[(#DRC=D
+bcEJO=A;W9][_Q-cPa>8DF(Ca5KE@;5AJU]#;R6b,Zg04&.21F&\58#287H6Ec0
&e^d\_1N-^,-7W;PX(?/()F,5B.OKXZV0TDQ0L;7NaQINS.0WLW^&0W<;TB?V5[\
\+)\V\UI:XF<?<e^IB]QEHC&MV7@Z1f;BLCAU4V>0[1+NA7LL.@a#?5#B73.Q)F1
[3(\17=QMd@d#)WMd?\gMIJ+V(_M)F1,GNWMT+ZAFQHJgB>a+#Gd7a>#Q-#>.P.Z
:UQ5E61Y/e6:>19NWV4JI9#T-.cZCX;/4@JAO33_f>QLIOY.Jf^(>W?C9VEa\b3O
G4Tc&1XD=c@W:&B20F(O+Z4Ge0,CLgAMO46+VfI_#HeIg1H/Lb#DN6\EYVF6-:L<
&3V1g@&E[2-^b#aJ]O+PI5B\De)),2c4V[5O6N3)SgFD5T_XZ>5U<8R_1PT05=[C
\C:KIIW6:P=H&1cCeI>0N@ZcbD2T4Qb<7VTI#[@XSe3,XgaCDOUECQS&2\be?IB?
FQS^)90Z2AB.:ZBYTS.S#=\\WOc&G2FX[=-C+/,:e[eU5\?Q[S&B4S14LP5Mcd2E
/XAR8e<_gdc9YQ=U-NHR3@M<_H8V]X2.?)?M\ZUV87_H?<)NK^86aYXH?cMZFSJ?
4&I-::,J<:.>K\Gf<gO51?<NeTd0:]03<C+#.Z9.-aaQWQNHXQ80cL2Zb=K,Da]3
07;I2I<eB=^_T[FP+\_WF;EL3,;(T96X_c..>:_,3-PeNa2L]_@=^6/5G.==]\K6
?PTCbCQX/[ES;\8\Z4V-.6JOe@M6(;GA_0[]1VTPf@gMZ)5AM/.E[@4U>7Qdd[,;
:F8Q)FH5-gd?QH;3@b^V.6D>:XX91QV<BD[92ZXTe&)^VQ_c<T&A@@L1-2+,+=45
@4)Y@ZPR5Jd+f]V^E63<IBF^Dc:N(:O]X>U1D\@C@N<9c;G>-A2V\A7<7XC?ND_g
YXQPP.d.I)H<7;E0=Pd^N0e=DFf:\]92f]F?WUMdaWKIBO;.:gAT+(.>6Xb>-[9H
X,Z<?5UC[D=:KB2YSWFA,=NGV/C9FGDD,-CXS0N-g8H4aVf#,Cd6X+P@RPf^Q/P7
@D0GZ7Q(HMQ^8IT-[Db/[[b&e4L==(gNT?[e,3M?c13d-4#45FbCX\\c9IC1dL0-
.+DSTE(0/UCcUDVCBM,K7R/CEDS]JXH#P&fdSc(LMaOKB>YQ6J@@0(4^4dWZ1OW9
J>Z#Rd-#&VGaF6L>KXH&=0L6D+)JQ;UMSaK)2FL]NabU&^0B[I]1O3MJ&/J7=b&.
X/1:PNaM7-PS<N-])X<FC#0WP<LPRHe24&T2)a?-AD=2QR#>+8H_WD,R:Q7a)N5]
-9F4G5<B-4e_?P[V46-U_SZ:a:8BMT>]T+_bAK\618_N._[)T&b^g=-I9MG>HWMM
II^#T0IONG>.FK-Rc\b&D^4?NTBU7:PES<GTOWD:1dg@R\bb>XNHd<K3&;AFUHT6
aeHI]NT\f_J]ZFM0>6]b;eeK#A/H:X\H&>_PJZ3-8MDB4GMg,XKf+_T]@Q>->BE6
<:(WEL.JGE6(>MCCWH[MM/=MYXE5A7DYFc8B;JAae#-=G-_@=/[HPADT[dR-F/S,
c\270aGNN)?.+F(Y\\04KYH<6(EJ0X;T#)M)4e0N3=g((OVY;RYB_DB5KF)Y4N2Q
_6\XKM,D&[J;1+-WLJa72WZJ,-JA;@QeIXMcUE3?@-W-1<:+5L)B#ZNO(_6[M;2#
fXNK5PJ)Wa^>F.W:O.#\YV7A.21,6R^4/=^aa>S=GP]-CX>4C7C-We>NKI7SUWSZ
.U^_E0]/YPZ#HcIfKBDaWI6J;AS[bTOA@36d8DZFH0+XE^M86G30ZbJ0Ub)1:@&b
YD8HV.FH?O^L_WG&D4Af/<E_>9-&:PdP\M17(K-f_F0(O?fO2<D?A@(BPZ1HGL[,
K7)f#&<e@>QcA<M2bgW;OVRMYaNH^-;a4]DL[g:=XO,_3GQ,MBB?Y,>5092.M6ag
W:.e3_<?F[=.UVMQI=Rb86DH:7[0I6@fV?-<Ee^JZfcb8fMYGEE,=[]GOGbXMLA5
?[S2IS:6]@5QK-\UN&#.5dF=Z+NP@^:.G+6GO<,MCYI@M4Z3SBL#MU9ZE(fUe\81
#T[A>a_L@[@-#A5F#R<;c=G2<8SHZHY9=.+C4TR&Z^8N+YHaP^F+ZM:&#NSaZKa,
+THTJ\6D.TKf_WT3R@DVVD4Q.B>Ha][2EaDX>_98E/#-fO31>Z]C]YAVJWNcA4>R
Ua#],aA<U[B9&8<a3ZR_b=X1,,K+F:-M:Fa#1cL5<N2<U5];A1M>VcLCU)1JbL_g
e[@#[+d=8a)XUK--0#gcY_P5S,<WLc<aOMOdJ.IR:#e[Bc-KIeQR.B@bZb(K3\,:
\,a;G-E(6;+7/_]K>+ZKg5VOHU:6g5C803\&8].Z2GX[R/A?X(WWX7I^d#1(ILD_
R,]\9PJ5+1b0?_CY.Y<4@9PW(/O5#7XK<L)g)I2XgP0XB/ESg0+(_Y#R^3a[);a&
1D>SdQ^QK@SPcI^[/\\3-cV[9?^Zd[CY_Z@.Jd>HHMc.L8_3E\5^S03PR-?U2X>T
fEC,L4OPO@<OMQA.0938KHV\OC;?71@]afAUd1I+@S?89:75:#,f9J[SF_^8&/ad
_c]4g9?0K\>V;,.(dQ#0J(NT39M4,=.ME<GO,Z_XSaC651\[\I@)IZ0VHfY4X@=B
aLG]f:U0AQ#SI;O67cCIZ1_&[]SPcV.-EGfAU+S?bZ+.+FO=]?8,@)7Z6f1P6CdM
_>H>DXK6#U7ISQ?I]9&g718,#Xc<40\YBdFU2KbQW2:[[#PK[IRTM<eM?:ODR:UX
<HYDfeX:B:VI/]c-a)S][DK.b+^I\#fYb[T=[#\Vc--AFCY./I6V0-NA\NJdUN6c
7=@&AU+T&E@91-+>5EcW++Db[P8DQ5PI.WPP\eGX@]\_I#DYRT1Q19W8V.74Tc=+
.>4:WNMH4LO^=LZ3ZA].6=9f8VFWc>>HZ:?EZYB?RDg4f\],LZe\LW\(2\(e9XK[
W<6OEH@8.52999LJL&I^]AaLCXNaC&@f+F1GDc6YNG73+:W[eE4,0Z,)Fa1Y@E+4
P4N;U;VH^[L>;@[G&7=g,HUCDGZ9ST2^(JGB\0_NCHP4][&>OWKW1SP;eMZE6W7R
2UdV1,\IZJYgKeIU2-2?;4#K7=aM(.D(U7CA#X:M-/Wg?XQ\CQ.9>f@,\[Fb_\?]
A)ZS(W4.K5eD3@GJ\@P=)R\/\eT^I?G=_,36Lc>UEX>3A?@GU\0)J99TQTMH)S<(
K,R#Y?<,cMaQ^QZ&C)a=Q0MF+0B#EHNE5TP0gT3#AZG7,fXZA,@+\E_&16M&<9=7
#46AD.5KHN+eU0,aP&P4ZT_/:>W\VNL=EWHE))J4U5c0++)WR.eVKb65MO^K6VXc
ebaZM9;fTac//;(<SD>1)@M\eBKI_3<3\)L?Bc@H0]^GNRZ\62cb6.)+4Q@I.T,K
GC8aW/0a5M\bc_TYe-1GJZSZ]RXeMCB4JMg]1g]gGXc0NJM@A0Z3K/^EXHJH5JBY
HLA,8J.0XBC(3++0(/fJG-Y3]\,N32&C<+YD@[O(Qc&I5cPQ;BN?:3N(SZ@M98f,
7f\DEN>c5QIa8K\V8b5Z#F@a.Z7fZ<MRXH:?06AWY=4bcg)1/,bbM:[W_eLGSL7&
3?g6U0]>?>2@@#g^ZQ[LL@G0afT=#Sa8HPD-e?Uf6UV2(A=D?0_9Z]PgZ\^T<F^<
2O]/8CR_A^V;D4(Ac:2UI-e.I#405+JK@EH]?:-c2CJSdXVI0g/^GU.C.7Q6ea7>
CFe,Z2+\D8>L<WJM9^cLHg_X&O9D[8K[(LHe+7/b5](a[1,6?@PBY&ITH?5g@(CP
OC>1;0N;[BA7WM8XA;[g5YeA?>^bAcd>:W9O6WA2#S<::aG614D9U=+M6W^f]\fS
4_eM9cPDaI9;&8(\f^eSD=2^?I^Z<a4\G8NC#X;g?e(76D;A4,g7Z>Q)ggG]4]JN
KG2AQ+P4B(BH&/X#68Q=S]KGO+3Sgd<GCAIO7&.(g<MJ36AZ,RH;>>+/C[A?:ZOL
&b2@Bc3N^O#NA97W[D910D&8[4QK84ZOgCH[X(e(Y3]ZKQ+TT)EMW7W;5TSXFGB@
?LR8??9^-G]E7^dg&NX]L?9V#Fa9fFG-VN^,(#Y\C?Pf++77R=eJ3b?D(2-EX)\6
=+R1[HNe9L6Z7)O#PT^A-6\g#Vg?]BVOW)=Hd403dEQF.9CBC[\\8@<1^/:X0LMJ
RS..LIb\b-DY[Gf#aH_A@Y;BMEBPg/@Kc[d0P3YO_ZSWV7_\.A[GI#<cc=AQEAE:
bG\f0W<1bS\FC[7S=/.Ub5,SMHWRO81-IbQ,DPU@(]_7U>@L1QY=g8;&N-B7#4-\
>R1]\E]d<=J_HK8[U)()34X+4&<_&QN((+T#^I\@M/@V<>@?>VP+[(M8)^>VLNI9
P(M-+O/fLH?^E2TbbIcTK[18F1/&L9JgLRC&fLCO]c[JaDZ8)Nb1TWA_\aB#K]E.
L6FQ]35>^+G4Z6TR&.Q[IaNNY]VPI\^4YRXBIU)^DHP9[<T3B1K?1N.0Se@PcFM0
1)M,?&.YdTJJ-NZCc/J8<?Vaa]?&g#.aYM\?5HOc:;#ZI\4)(@;CD4IY63&&bOI4
967d@NE.8F#d(fdCeXCb.DMWgNAO\(TYcC(1+W?SR^[^L+K;NP0S97)+,?@VRdc.
N&4e5-OJ=QQQUb)9gUF:QNgJ-&Qg9//(DVKe[T)G6?-ZXLD^\3-1gON0/P)N[BUJ
9,HG3Ze\63H+/>=\LA(N6PJ/J]<;W_dY:T/9L^V2J@4K52URK^#7G#8[8\=e05eg
GD0G2([c=#<#,9IMK8(X,,W&GS6_5,USIZ[M^DF0cOT@-Qg_]c\RE2UD.K(E_Q61
dafQLdcOR45^,Q;=[/861@2aNRJ:1NJHOWa8Rc[ND/FJB.8(]RP.0;0,^ML@?1&2
_=f+:Od2COYKCI5\AV:9BU#;39-4g3GUI1+D(.SK_,Na0UTgKMO<c+2DB._C6RBb
^2:ZO]=>X3^8;4R7:NA-<0J>ZZ&_I3_<ZH<a?71KJeH\3]Z&J3/?^D8adDL)BYB_
IV9R=LQ<ICCG]#<2^,S1:\@#EDO:RfX^Z83EN/B.=LAb+Idg15<O((B[D:XfJFKT
2Pg,&L9NZ6-8MW/MTe[:AT>g+0]H3=.7N+f1CK\#KF-cCHY-[C&P2X@KX]B7LDKD
(BNQgaXIS8ORH\b/+@eD@dR@6);AYM-JHDfX9S_YTLWD>.;^=2Q1?(?\?XLf,3=\
&&TIY)=LYET:++bIJS9/(NaFSGD7#D@QIJXCT.DT;>V9.=0O_,U:CX:;NV=\8ac/
\WeB(M/+I,WACY)0(BTPTaO.)X&#TBAF^<Y=U0DQ^7OG-=Z/Ie/(Q0?4K:#;>PUQ
4(d29DW7<;bgGC74=DWE56QP1+Fd&9GR8g>MHg\.R-G?Vd#@d1[bQY8)Z\<RXW.4
DCd/L/:032O?>C#1WALT_ZY5RFN0SaHLHHg3D6S>C)1]L?SIMV(+TKKQSDbfabSM
Q]#++=V?Kg7g:>K=E1O?I\P=HQOWP02;2TB/bG4SWC&,#(NEb-g<&:L+_aF10]9-
W-YSR.ZY)5c[:XBHO8XS63]0]&\O_#:XJ^A)0MT8L^_;?a)8Y<@Hf[2c[CKEPC0_
D@I,6e-16AAT76Kbe)5QWMMg3#ST@D=6DM#Q\KDAa/U9,bD9X@#B,<A6^D0X2LA3
=Q]P2CE&W+OJIee\,5_F.>@NO.?S;L(J#&)MK.72A_b>D;C2LGD^4SeQ_LQ8AF;=
a^IG@dIK0K)XB7e][V()LWG-4G/))FG->cd3^X\g\X#&/KSAId8-6ED/7N2QdDM@
E7@=cY#YH31@PC#L6-4(deH\M>[a4c\Y&0e/T72MHRG8B6);@IeR>4a^fT#:S;G0
O<^G-<8JI@-5UK&IfI]B:5FVY+E<aHMId=:K2g_.d0&W0TbC&[K]O^<KQXgLINYM
O)ddd7fUB7Jbf3QHKPXeW[:cg/3QM@6/aJP^1I.U<2(&Z9O^<PfPGfM#_,P;#-9c
D)(KS.X[T<9/8>]S/cG0.U:@TP0NdSC</g49Q[UHOE:Ze8H/@#@&KRN8NE07K;:H
A/DVHH:7K:E6#L&W&EgJEFbS(&+VJG1U?SaBRX5e\Fbdf-_DWaG2@1/&NcRa8O&A
5H+^dC&1MS1G5XAF1>=_.\Vg?&)I156T<(8O4>cdLKKfD.]5:)4B-Pe3>+:9>Y>Y
O,75T=e4.@KGdPW[ae-ABa,YSN(>Y6NT4DJ@Y3XAX8PMB)Sb(M7_(e=e4>c<f7O)
/cbNAS3]cIW26ZgXN:WgKF]B116:5[2.EX)43N.g@ZQR?]EYTA]0O6&_>8J-TKO4
gCG,&N18W+8Tf)TLfaEbX]egb/40[TA+G^_8>X#)VcK@cFW.<8QUDF,bVV+,V8b&
]_HM8L&066336^#X5JJBI4.CR03LAGL0ZX;Pg<ETU3UTLRG.aO)(,6>@2df_1^<G
&F=/13S>EDOb]>_@]C00)/c@0T46\gb+.+,XT30dC+5gA9W\T<M_U/(@:4<U@bJ[
#BYc68M?YTR\]RN6Ra0fP62G7U6)?[)7P6bd&c(^A6PB:YV?-2LP[d:BF;1aW/6U
KQ4XUU1_3e23G-+L;MPFJ:g^)#JC,e=);7[2;U=OW.NSG06:M(@NaaRZ3cV>@UAG
IcCR2Cc:YAFBW>&X?-.P>9S.]+@)9@4K727O.L6R&U#G;9R_(D(W-2E\&5N-KUeU
.8W6_L@F3;7L00Nc>2Z0cEI#]bC3fIN,:8Q:X;Kba8OI..KT.27\#=J0AP4A0<1c
GYfaQ[e]\3(_KdDIE<-&,YQJeXRRFZ4M3O99HEMQFcc7+a7.e0?.V6AZI>//E,TI
2.65U;X)F@4O3;+Jg918<EEWW41M(.&cV.gZLe6S12-=;Vgf,@LL)e3VZ:;8S],+
8;V[O9;fVP_EIE6)[T8A.8HOe<Bb7T@IR.U8(OMJcXeDNaULf<dO4)Y\gWCAA7LY
W7O+_Od=K<&,9@8&^BODCXM47S#.dX-/;YIY4EgU9?NgSY(59d5&3WXWee>/?cD=
<?7e6MdF6KFKNH(_U?BBa4RY)&(?:4#WDO0)_=bQ@B3Ha7&\L27-GT70.gG@3P3/
fP].(aKXF^RCN+:cT(_Nf-67&::V)b8/D[_EfQd^)B@dATUMJ-d4?J?-[VcQ5\.W
=;b\bfVeeFB@W@ZKT?.&D&G8NX<JC/5-BS?DX7CJRb8ETbZa\0.XH.g63IfKDc^4
^\1R&WD1Rf\);_3I3)C^e&PE=L8S_fa\R7=CfPYg>>-&SP,,FS88Pc-P]5/bB(4?
79KVO2ORN#[dUa>QWR;[F05a<Z]a(;(D0(Nc3)]1a.:I5ePg3BRa;+N>U<\,/HN<
0[XZbAU<^9P.(B#:C=.4bcAJLTaG(?X7,BC7>U?U1O#RYTS(c:GCP)ZO?X,(,_+O
Y+KD?MW=f3.UT7A@=[.65RdHRHfC3<Y8:UN+BU7^X.b6SL112LDJ#e-_2I&1<UN.
9LcW1&V4T0I#(Q8d#>\@F.d+GHHGQ,DKN>>HHb,dF5g:Zg>a9=b=\RTg?b+SN[eb
^\SUcEdbZ/P)O3gDX/_WW5>\UE@XUT.9TUE/TTeU:a?2WEg5?PbF3Q]ab[<DWF@#
d^T3F#^Ae3E1N;7][.1CNWGGg>DRQXgScR)8596de-]O-gW_1EMSP4).;&,H)+8Y
69MC#P-P+<GW540E0[BeWZdGRF>9EZ2ebOb;TE>)>#@?eC+ATBT_C<2WRTHV#Z>S
;5FWWFUP0J^2UM1UM4.Q,64C5([b5aIQbVQ?_K?eB\@IIfII3a,;]>JcXCM44YYY
37\/[bU;;KP[N:WY3b1R\KZIT4/fP9Be;-(,9;/M7b+0>/O1[WZ-790(6-c9R;QL
6Q9PCWTHPPPJR2b].V-fJ+89)@2FYUG0LOLFWC;J\#dF\&Rd491.K,0f#_M9DcK0
:&BX7Jd_BV7[@<7IU9T)M(8@+NJ_5&((].I:K\A6?;Xf@N@.J0;@bB><bG+Xee;M
^VI=BGTAEd<#R^&0+E2ac)KRT[G(TRU?JbF2Vd,0;NT3@I:Y\AA53+eP.[&PfSLX
E_Ja#^H]HPdMPN^HOG??+G]E;>)W[M_6C&NX=JG2@V_fCXW4OA&+-R9FL#d]F(+7
,)20=,>KDZP@MW&Jd@1N:,33Q(+KV.I8V&X=7U;-2T((81(eY#cKN;/ZRSW<QGN5
M]O[[@?L=_.I;9M:]a]fL\-4/UbEd.fZZ#+FKVgRPJ[L>?Zb3R)AeIb35H9OI+0+
>PP1dUH?#)M^\(AN352E.-Ud5c/+/C9MVDO,.WfH8058^5HM/&)6<[Pa1HKV;J>J
MSXB)?GWMJ2JM,:4KMgL#^S,MB.>CV;^cA/;bK@TOM0E\DC50L3N4RC3LWbG9(g,
Q:AJB)gPS5Wa85W.;]g>I9dA<=MS@S_[Z3UId,?7#=U[TU?D#g^9YZXRCbC(O5a?
WUNa:4E3c@.V=,:+:E-K&>b_H(?E1VfA]f[<4.WAEA(#AXe^Z?,7c)]/YPUC\8U8
1RHK-N&4^&&OIeA(K/dMdT]-W0VPacW?MQR&D?#HIO-B75JFf&P74eO-KLdNVZ_2
P/[c(21FKZT/.WOK#L?<\Mb,cG_>PF;)Z<=1Cf5a8@B;&>K:6?#_M&#7E5P#b)L?
(&30d@2VdTKK-W44DW#E1F-T2+C>7B>?d1786E;PM>aJa[a3]GA&IP_DS?FIBTe3
/39NISMV2)P^YPX2^ab07R0?.KIKX)]GO+W89R9[dI\U[4HDeOX4fGS+BgfY9WN,
,UJPUaU_,4E_DZ@9dH8)VI^X5;8]1RbXK#>GFFR<b4?34_fb<cbe835Fe8O^TV]1
JIdRM[eRZb6M<B?^:^&S5B,c7Z)EgBE8[&BZW;P@G;NN_;9CE6H;+bcGPD-@LGR[
))I_<?])0[SMBM5B;)a&H11F4\=./2B2J_HOGXQQRQfI:Ub,^EVY(+W5?a?E:]Qd
gM7Qb7eEO++dd.^bKT&0FQ)QG=/KfK&8dbMb1A8C8BQ,8B>Q0Y((OA-O=:8O].[f
FP^^Zga[R9/HR8IB_AOV&I]^IFfZGa=dY3:K)A3;\KH2F\g=S2Ad3]S+MA3^HLUR
0?^.SVB-&[W38_>YS>=>6[Og;H1T<)ML,c_>?5;fc:<=<N#If5cJP11EAYF-J5Y/
YJ7)T,ZML\TUWG[B:cB<f[(=-M#ZOOHP<Wc_HC7&,4\P9P[eY#Wb3gMg2JQ/(.+A
A:g.IK9.efJ7B@VO1+&f]\EGa9LC;,+25J@XYK.PaYSCPe_>aLeO0>f5(?I1BKE?
5]IeBT-QXabL5QINJg9+DNXT?d/0E;#W[(FGRIJ9=TLB2B/<@U(6/PTY\LV8)6g^
VSHM.XcC],cE#a^Q)]\>3T7O&S\@S^)&8RE0VIGHIALU(]PSZ.Q544G8<M8H)V)V
2X,TU>^Z@EZ?+TMC@_:?-PH_d/74c:=)Le::?3IA=-C#NHeRC])6_0.1&.?a6e5O
F>cf_?BPHdP04LI2d(62QfX&B#9(E<0;aX>7P7V&LK)X&A]S(eDc@@BTTQ24Y?,]
-X6bN>F09H-P>3Q<g0)=;=7\FQZ4MRb;/@\3N<;V\(1FPZR<1BKce\PQJ9&DO,-E
Q]^))F<1\.d[X@>E^O?Z:5E^R2f[TN-52.FU9JVS.b_R&R\PIea<GW[JaLV_.RK6
85JDKY,G3]&da#D0U;]a9:AD9/JQVbaM<3b+&NW86;dJ>)QC^A=#U3(ePQXK0F2N
WcXOPcL[F+GN,?IGU,fD\.5TSF@L@E=.QC)6T;H#LH;_eECAS37=L.J\IcU(b[aN
O.194f?9MM<ePDD,W]b_,E.5/<)YSIff6fKO7:<.^DEPDYbU8D.cgG\gUN]]SI<2
<Bc/;eJ9bfC@4R&9N2c?+_P\Beg9/@?SO8YT>bgFO+>9;5ZRR,0ZS^0Ya1FCW2_\
U>004<cS#ET#bU>3Y@(<S<V>B0+EC=a(9fK@>+RAM^,cR.(Wa2U3fOb\K.C=HeGK
Igf:PFe)K=HA4WfbZ^8<d:-?ZQL5]HfPY7X/J[B0CE+M#[J^E?A2+OSd)ETPAgG[
ZbQOcaR-,<);M78E(_NYA5\KHfYGU7+J19=BV\<Q0A4Q1VND+3_0\QZ:Z2_[d]5M
1fPfRa]7C:G;1aG2>WPNQR:bQBD5+^B[bW.\/<6K,YR&-SI&EfWJd^b52Ub@P2BD
H-L#XX3;-=[/G56DXbCHDL,(N0/Y@8]F1gXcMTIY.6.8N>>T0K;1=F2GV:bJE<\d
a]HCaSKb<5?2VK?<YXPV2)c>]R&Q3466.WMD8VZ4/QIERZbC]b(60#/@F0DbHe.\
c8/.Oec>JNd4OfT\Z]Oa7&+XH+J4BdQ,3:KeWW7X^_M:[ZVFaCVaBVCIN<1EP#?X
T1N-=bWIA.\]db,g7d0e_>FAM03f3U-M(DLf^,4I7-+a@1HQLY6Q9Z0V\4K:)fB,
4Hf-K4C1+#a#XCb@#)CgF62H]f8(H9Z#d1Q=>bJCM9#?X:F>=[BaIZfTJe262:#M
=D?Q_)X<3Y:&W85]8.NRF;C_(/=VPM.c&K_<[A0:R#53LCW5/d&60]PH\D&G(,SL
aE8d62A<UYBZ2EF,XAfDD6bPge(.gg[/d>L\W-<Z0BaB]LAbB<+<AS+Mbg=W<Sbd
fTIUfLG\b6NI,c:QBZ-7L>AW-@2aD3FGb5@9,6B2Z7[W8&J/MgJ3W,\IUHCJAU\S
7f)#=K.(0SDgJb[M8<Y6d.H1OaIUbTZ5\<6J>0QSNATRb/,</4)4B0eH?5fb)0?f
RKYM0&\[=RD+;LRfW+Z-^0[5LbUVO2,QAER07YcT.SU(NF]a3Q;S902_L6],]H,d
D3R^3Z)FD4#gN5dVDJKPD#UAAXZXGCEdV^,K<>D0X+f]ZfdP)HLCgJ\.:9fB[F?Z
3Z;25K#?]QdLXUSW94LC2cE11g419aY8SQYFGN;JNVDZM7&#9DJ=c3FTTAHea@d4
_;H[[7/e8JE<T^#MN;Lfd<?_(68:)Ob(654?71W2T?]#J7e^EL_C]]N,_024X@D_
JDQ(_CJ=;P@Y\#8M_C]-a8?)+RF\CE(<1RDAc\\YU&?Q>P7YD:I3cF3c2LIZEDP_
#;a?&=9d>aJ[GW/1Q4e;c0.Z5^9f^+g5]X]gFad=(7fAg/KEOF?I0SJZU:=U)T](
IV,U6,F7:2ZQ:gcR,^7^RX]8XSF5FT8)1a2f]?X?OI[:\^L(,CF\1^Pg;>99]fB4
MY-g#9FS#g@=F)#Oe@IOG#4DMfUZ9=3bNWX32AJ<JbSAD-ZbBD)@/O<N@6GPT4CU
_5RMDIGdW(SEG]f:V4ceC;;dGTN#Z[HLfU>cC(O.HDUKDfQfD(bTQ26a?M6\>&#-
+LFbOQ(WCfd2D<&KX)U?2<cL@BL>0;6<DHA],8#>126G5T<.+0d.2[S;O^&8W)5&
>9PU,6Z1Tc+/F)LBHJa86.6X3B15:V4?;HdFO-D:+X)3[4eCE]N-7EZ;\#EY1L+g
_U)L6K;c8GTXLTJ98R0gNgJQB:LMS/a(N+H_EgM.BcB#cYP:G5@NN:6aHaf.7cV:
Q?UM>O@PA.DUQ(\&5>C9]B+&G>9SMNK933VY_XF?VBRFgZKF9-&=(E[Uf2d5OU_5
e0GIf40Q91,7ZAJU<b2[4V2^0a[&Jb0GCTZ;4Ug7F2f<)(+AEBGWEX4JK?U.W)84
d(ZIYOY+OD&OcS)9/TMM[b)N.2X7NS0RQI7M):LeHSW6W)EgFT5RcZ[cM&&S^,/#
T/P/9dbE_5ZXEB#?P_[g?SA25>TRR;O5^,([J41]3-IVI/?JD#57LJ+D@VG<O^+P
=T7,\MT7GYSbL18#2Q#LT=8&QAO:bNW.?@d9AL]A2WL^J\4L?\[b763ZFVc#>9&D
>Xa1RcR90?0ECJJEMH6XAP?QE<J<[4:e.#_R)7&d2>)b2#WVgXM@11/S@=]HPD?]
d]T-dfC4W/f>DGU<SIR_7:6B2-H:8V^Y_[]M4X?(^M8TSD4QA_U-E9TB[GY?VUcJ
;R2PXWEdaJH.-dQe\8@-SGCCII2,e&0GNGCU0@c\)89)fJNONTJY0@U=82[DcO&P
=36S7BV6D0DdaM&+4T=3B#,53UOY)I0:a]Ng>[B7EgFgJZZ.+Ze=)-RZP_0PBI=S
fO85JYFS@efZ/(b?YLHAA#,2\M4><2.D+<=O;@5>#O5[f4XJPXMNJ,4ZIWSP<f5C
_,g/_5f\cJITFPgP0F[]db5REI>EGH9EPPg;A[/7C>9@;):W-Zb4<eT2)FA)G4O_
M55[T<)@V#/C/]Q1<RYM.:<@@8.2.VK>Nd7YVdE(X1UeP^NLA?-DD>HD#.:.O,E-
=H,QOT9>Y9JgL]+I/Z&N([Hd4_I/6P40,5X#B=6S293C_;G67dQ7ScEc2U,U5JN_
eP-eHRdcJa7CXO?KI>cAVPCb9a22YCce4C;X<-SU6d^0IW^4W.242<=SSPR]#P+7
-85DT8#cC:SDSQ[.F,M]HATL_NNXJORebN_/D+LT?_HZ9H+_#I5Y8J;SS#1PI^[+
f0_Y:Z;GLd4Q&U9?FJ-(EN]CK+R;1<ffVYKB@_85.;\TIT,YeY/>e:&>3?8R[+23
9->JKJ9DUJWS1E-=c8<BFB5LWY9O.IH#&Se9bTAX<_Pag&7^1,4\/+NW/a=#.S)N
fQ@f4CE.e\:?E#?MX+N<[(;^aV>VECYK\_/#Q]&fJfAD),VDG9d2JW.7,cXe93#N
T_[;+\QQe.\#3UU6_bfEWY0W:4e&Zc4WT5ge((26KdN3H^@Z.NK\XU<B,=/(01,c
b24PSdIR:8VV?E<3SaYS:@b7eB:<DO2,#-SD;2J3SP62@HGL&>6W^B.NN3&=/gLB
1V):;Hd=HPGFWGXJ],XfecER75-(+F]eJfYcbU,g;;9LR308.-1aL@G(]RCZe/aI
#YCDfAUH[H+/TW5Y=L5IP+=]eKKZ8(,FTDVSGME7T8BF^V[3.WR0):(9JZC45GS,
a^FG.:Yf(PH^=/H?QI.GHJ?bgO74>G&,E,[CH7g2_J3=?[_JOF:Ua8#:D9H^PY)K
7]I>(3K^fHH0OJA+1]YC7PU#Hg?Z+YH^Y/09_cVVBf_6Y)TVJ_>CDdIGfZ3d(YS)
-[;OPATOS;&??<BK^GYDb<UL#,UV[faBE:LLKVH,@60AN4OUQTc:<K5K+>=V=^F&
2:TL#JD;^M2&Y,L]\GH8?1-L0C<.?C2fBT(I>/FH_#(=c?CVKTIaZHd,L^Ra/JR\
2P_/]NeEeN+^]B\:\?)T#TN?f0eI);CH5EMALFR1g(I+4R(CZP)?TKVZYF0<DE[c
U&LaENG7^5?^SW-WbMTO#F)RYaQe<Y_6TLR261;S#CD-/6E.b0b[:H+_[>[62_DL
<GJNOf-a1>?H=AcLBN=g@85>_4E9Y6K6H[P@d6bA.1a]J^5dMHYGJabg=;eZXK#>
]aOH>BB]8,:cK]-3-MZe,GbQA4O+;CX@5ScZYR@GW72dC/B0Zc(_:X)FNY)-0Zd>
)7e#C2ed.LeB\;ceRONQ<8_.+HTe7agD9@HG#Mag6^/P8YB\_,^T_J7+^O9YbZND
,G.X2ID)EaI/3bT@6)MMf),M:cgPGe?b[PI]ZXeLbKDNbX\6ef_V_e#O?N#.5]J.
//c0#3O+.1^FRV>Q@A&76eFQ<RIPM:^SW/1U0]b@PO6:J0aUBNd-K/AV,?DTK5G#
6G#+Eb^8+b)1^TO#8BM>24@b[AT6ZgeHE^\TSGW+P8@?09LTV>@fC6^I.a7N3(FC
C<R7X]M+43IMAN8GMaDMAK-&NXbHS5gK<14IZ8S?Rae@<,A&7-2TL3/[VGf9X-6;
3#)33;A4<KD[))-ISDO?EKQ.(38Jd/;OQ&#1gU\J+VMM9OCcJVTS96LW0(V5X-Y2
U(MZ6;-EeWG+DL1=dYgC891+6[>17CX0a;5Y4FQ@J-4<NLD)3C;<LX<2X5cf?>7a
&O<?(SWSGO2D<5.UCT2,UD=.b#@<F2RCKL2V4V@c[]N)?.9)-RML&8?#_BV1a6:7
UgJA5=(R3HX.G30HM^OA#WJ6&g^/];0e9-(E;+CTFdQE]_<)Yb2EFSS-bU(,U-bW
;^93IFM]T5JPYB;C#c@?F?^SeELUQZgbd_f?[=T4caD5LZCFg?Jg]L;C^.(_L)&a
B,Z?N5./P]6eK3&.SWNW<G@;)Bac7?ZEMe./,d1(7c<I)c[A>J,f9(@7Bfa2VO:@
_,DV-EZLPaXZ=L8E+8IA9OI.CG@^XX8\,TaE>\)5ZgST1cDT+4^P/bIe<CgT7Y.=
LJca^_DLD)=-P#_4)<WSWdW])&W=f_3NdJaF_U<D_YA]4(?M5;F;6\NDW=]5(&YH
J]X@-b+K0ZF&cGY2#;5@=.M<(B)U[g)5&4?/dV5;<FH.B^S=G;LaQ=ZNHTQX76O^
GK@.a9\Md0E#+bd=TfXJcP<d4/I51_\ZV+??42b8\-+V6C8f5F8dR:X0TMU&1PPW
-&:JaX-]Z)1gI7X0.+>cLbY/(6=BeSP?E9.<TVKYQ6NPGT73gKW7[DL&F,H-\eSE
?U8H>g&-K;0<0]39KX1WP((4Kbg(I.dSH8G21IYK&T3eS,WWIg\E,=]Y@42.NQN-
Occ3A4Tc1S<KGNSB#08gY#X^?^2)V??5TUGPOY/.eY.,[D8?f9cD;MJ,99<?TJ69
X.BXP5^K=55SR(g16/?L=6P>3EI0T8gDAYZBAKee,Da)K)9E<0b4;=S>0Da>8]Ma
Q1Nd06HbI?eA?PB\2,/LIQf=2O[J&\df-GFdTcQe/^<#IXVaN?fbSag4C_^4./P)
U&KEY&,4QB5B0?g_6>_+_KO&8M7A/a;UTRSC-^77);&?0a0.]dZ)9SO?a<_^<ZT]
&HP:VKBeR))\QK@M7?+<LRdLY-80LAR(-_@,d<GLQ0CL/-+AZbD;REM78W9;V5Hc
_X-[0.69<SU08a8TD1&Y;C>3W:DZP,V/9,b=JA-_RL[dMX;=MZ2TgV4)=aSP:a#U
&W:gdbAQ@IE=eNG0Q>W1P?f+NO9@9J0TH>+-/E&:_LTa49K(GLN1fXB&D;4Y;1WE
[+;BSNM@X(30>:dMEDL+B:f,G]bQA@C,f^G)H[K]3.(N:EE?(B]>T7Wd5fN6:G8Q
&_XV4V[c[6K:>]50AF/6CD785B72>QY,S@gM-7AU:Q/GQ[F;[6<H>ZRLI[R;<M-G
B<AI,\-W8Y\T?]d8+e4g+c8(QP&;?^Z^U=()Q::Nf6SLJ>HMf8U)B5gNL0@5O71>
cO,.E85JKK\O[8-<]a4K+Ka.)\C_:CW\1\W@gPZV0JFCH3d(QW;4g\(K#-C(1_#M
RPZLV3[2]0>VQbHeJ:[<0fE(H3P0H6d8/AY;\SgK>d+P]Tg^;KAFV,Q,.T[&]DN5
)@XJD-&0.&CVJY@WK4IBU;e;T6[??cEa_7:MM(^PQd461PGOMTJdGc];K8/B<_DW
P]dVbB^HO+3CEPY&C0XgJOP_\#4I[;96EGOU#1/d30[=/I(2H<FJUdS]A>c0=ZQJ
SaB2+ME,/X3-92B)2Q0Q.=U6Dc0eJ?]<1#YD#:JCcdJ56XEf-&KK[BC^_)_B5SQ9
e^\&TE2D7_2H(;/)]<DF,<8DOMgZJD\Z-QI.]YBeTMJa+g2C\L/^<7JIZa#(9LF7
/OAVE2Z_ZfJ<[_E9>0ICbO(2eg.T0F6<B>ZaQWY/0aJY3[c0ZTbTJ3:#561/(0^S
C.Pg->_afbg^64G3fHL\bU>OW4CICP=KG_ER0H\2OYSaOSIDQ.)+Z\eJJ\I,^c_1
+U(KKAbY_6OT:=Af03OSU]LRN561#2[GPCED6&H2eIHAOe>D^G>Y(9F,d(RF0@S]
9E3>6?U509e(;B9?M60P8Ab/aK<K.#67H;g^-1LT?Ec^5QbBI2Z0XgV,NYaP.J:U
_95&cdgDY&:d0e-cg[+8R_,dE73D8:4W:=g#Agc)?Pf=;Ad\4dV9cbO08RBEXC,Q
7d#L0GU:RHg]C3e7HKc)KUefYOZ,&4KE7\a[L/P_;8)[]DGN/Xfa&fa608]M20)R
Q3bFA5WXK]L+@&N[;TVC71]/:>-b)Z0M4:T&N1L.-eN]7R.Xc6UdN<L=^LCG<U?d
I6Tc5@HH9DR[)86d1FIbQ)YWJQGE2OB<f7[2M#U7]VX)2(3?D:1ZXJLEQ>I68I#c
WRJ0R/P.JXgO5:K:Q#dMVb.WSgGgRQdNf@g#/eZB(/J.MceX1;#_#;<4/3CKVB>]
\GCU]SUHF=,/NE/-4F]@^^,Ha]GfR34A57>b:?OTH;b4<?P#)B8D?/=a>(CY5H)H
WFg14^<,5Xg4R(fXfa6EC=1TRUWN#4_S6-H:J/#5g(H/Sf+dND9Xe>4H4-@=&JW:
D[(c((f.MCZ&_WIFKQ\dT=#1Yd;Od;JY)TIaXd3DAUYJD(_<,Rag7ZEC0e;Sf_a+
AF&IC)A0>^9WHgac>8>AT#&9J<^A_J,I8?F\Qg1RUO+QMDf7UO5^T?D?5)c_7-Ce
PI>7)#R^NH=Z3,_MeU?-EZAf(f;\6AA7Ge0W>RVRU.7DFZ6eXQBMS?B6Ge>ccN7<
:g7,B1HAF5aX[>WJ1a(E2Z9>J;8^BO\-ORB3ZB-+T7\BV[^_)14#S^UM-C\RDL.4
6,f,9dQR<LQ##]8S5XPG,0>8@Y0F1F1H:2D?IR]C[U]R[QeK,_(W3T1N<#J^YcTM
a:XJ7[d.]1DCP[NICRD^IYRa---//QcUD1F2,>F7MXCPc9N.QKN=S]^,9@&T2f>K
8L@N<#MHLYB9::44J/:/&HUQ]dS&PG>:P<#T)<VW6dKXZ:);70.E3W)b&L]&;;0^
Oe_geLN@ST6^-15-e>RL3L#I_ZHG]Y3JV+2(N:A7;Xa6Q:CK=/cK<O#d,(Z4>M,7
TFA50C]K:)4Q\5]).;_JGfPZE__/B>cU]?T-P_.ZFI.FfS^@Z,[E8@G;PbD)#dFO
[DW]W<J=2XdB;R2C6BI\b()=]S<?RPgH7P<Q_P-HND;R.@54dFB=9KNMDF0Nf+P8
QJVgXBabGZOK/A2LfY++0/.5-ae7#]3;Z65^RG<#)Ic,g7#)Nd.a(KZGBQUR5J4]
;1QB]GU)Fe65/b;4H4Db1-+.&cEeAJA9fFU6O09@PZTVOd(Wd?S:V8RW.a_+5EO-
3?64+/,b8DH;@##Ndg^c8<V2G:-e)_>9CgZD]AE)A]0ID3?UUW&J,U-7:[:V/E#N
+)d\3Xb72,-WPO\&ZE[YP]QWB9BX\CaM561/I5\PeA+VG[U5A>g_O#EeZIIdR[?W
C,C=aDW^>c):\[0S0.c1O[1Od-Z<)S)+HFb:L,;65eZ9.];@(=Y;ECFPZ)+HSdUL
\V#)]e5[2Q.:S_(L@3dET=5bL>84Z1eZW?IN,G)8FTUSd^?8C>O7=a_6LD^&2DL8
c^APNCX=QP9PQEG6V2F?4g\OD5]ScJ6]6_/9]geL=[UB_L(-Ia>][ZM]L=4c&V6F
69Q]SGbHX:W@X8#AGHI4?JPDGA7.Q0aFBWK&C\=BP4M+09VY>Q/^./LO.9K_d#P&
Y#5fGD<6<AYG[&L(,TS#H/B1b(0e1ZOOGK:?WQH&6_C&YTUSE:WV)f4Jg4KC352b
UX?K4Yf<#/9WKLCMCHG-2IS-Q+dI3N>N4RK0O/>YO-WAT9K]\@2W:IH:2<f2(6<Q
&J_fE=:JcPbcJIeFSDNZ;9^2^\NTF;+3\XR7ET7J]c3;.=gEZDYc<7V][5d^YXgV
]W=(B:)SA/M/,8I8NE<T5gMK>Sf[BL6Pd@C881<a<f&NUH6=7WQIX_S1++Q67PSU
X9/]#d_V^\68WH;0<0b)0<]N3VB]?4,ZWgIa2T?J<QFO/S>R7#&-cP?ZL,-Q+G0G
M[]V.d,=B0d08RLON3?caZg1.^e31aL2S(983HL@d)LZUT6DPU1OQ&5KBCZdHCT.
Z?G/1SP6P1(c++4ZLUKYWSF]<47D/^X\B@Z#;;1F:W8_]DPO.QBgQ7E8T0L6fGee
([a=aMV/1T(6MOZD.HC&gRN]65+B5-3Q(Y2:Q=(1O:XB((NF;K?#\EAVKLHg]-Qd
W3dXZPbXP1M(,-3)ec:\BU8WIeYf;Xd7ec;,:/#@A&K,>AMPG^2E++N772:HfFaG
UdeYJ/O9L?CLWA2eX4F6R#?)MF70Y13:)RSaWV>QU#WTa\gY_7NB@Q+GH1bf9DYT
;S+AbLA:c#R8/5g]\@ZAAE/8:)Jd<7Rb^5KIL_W:YC?5\KLL]UG3KQ2+<EZGaXIJ
[0<a5>Q:GY,-9M.4d)TfHQO:/-IOYE(#]7X)&f=\)TT7?-c.W^6c/G4YL8AZ9:OV
/6K,e5.]4f>T]^4,fF[8J2.1M#Z_GO_T&L:?6;c0KeMNT+cOB9\<?P(N9S<J&Z7H
gK;4TQd\4]#/X&c<RQC?E+gNMH2fFaMI.4DOLbI>:a.\YUA4X#IOEWWfdaWX^Ig_
P+=cf<\UEW>:Dd/.B?O6)4NQWD,gULJ7O)NG=A=WN62VX#^_SG=28f@)THVYD7dS
ZTB.04]7[MW3##<aYL)JTQ,XNVJ<B,IAe@)gEF<6(gZHC&\28L5V^d]5IF4BF0FC
JPYd=FLM)ASPCcH\1bBK1KF)2;(;KZHa\SWR@V^DO;VLL#@_JU)E(>eB,J[5ONQ_
?6@LTYW?XCe8Q.ZQ)+^TYOHbK^&V8\QbACVb6+-CYg,]K?11X<Cf_[@_)I(Qd21X
YP5M2CBLC)c?8L,5-\.fZYc:@^Lg338,AL6[1S,=LTA(+^fV2ELZ-U4E#LRLcHK5
UNZ[-F0d,Y(g+SP=:G]39APe)]3Bb10UOSgW=JQg10;U/D1Md8fda\]_)_7ER>b2
aJYIK3A+7^J6>We,3-YHEXM,:cMGDH>+:5E2H2RE]bOQ7F/EO#2_aFG0a]]FRVET
b1G+_O8WGPGDTNeN:d^MA@\=e;FXUKD)g&5,&MR8B-T:O?J6a1Q9EfZJ?a_@^_,D
0/EF7e9YT^U8d[#:[U/.eE4N]C.6+\gF)4fFM^[#(K.RX>_8JdG8[+e[dW>S\H<d
FF1&-/XL[;Z/[^(HC+@QIaa>5^Y.),/VU3C\5&5dg&@8CQFF/@Q@GTV3IaA;GX&1
CcdG59#c;R=E8DWZIULAULc^5L+W2;,_X=&&[7F#U/,3d^TQR=DI9)2VP6IE.I=3
MN2WS@5Rg+c&FKKD\(Z]d;;fKf-Q)Z=8FO^-JN27I@36g;Wc:G&8)7=dVDI/A#@(
H8F3/O)Vee4TV\a+7RgYD=c6/QHYKK1#>Q@YA4@J@\aLV7^^ZUK1ID#W;AM/&-H9
M\=_3ML16X=(;J4BL9[f\@B#]aO^Gc-XN<M2.EG^&PID?KbP]M\?7#8XI5N)Wb=@
ZPK)2L<3VYHa>HZKCf#dZ9JW/Y\A?J(T^-M@9FVeDD7^SK=B80KgYg=(=)Q1O\cF
_>2)D6V36a/8(&X_PW;J7_9YF2H.?EI5>)?/&ffb^=(Q>,(O6[P/_SD>)#UPB5^:
J.2]<8b\\Y,8R;DE./e[J5N\M6+N[A/0Jd2;KeVB@g2)+:NMWUQ.R5A.^>5aR;VS
I5OJ3PW)<c;_d@,[<T3MYNGbCeTLd31FcM8,)fEFQGV;gcbIcHg7^f#2+.UR0SH,
#?UJ.3;5&)E_A<gCfI7,1NPgU&5IMY,.ca:f#]c;?BQY.g6cM)<E4YB6ID-,3_d2
V?W&37dGL7^L&dL:P#.@L@g73S>APgV@g=DPE^f^]eNK)7KS;7_eD#YRVUF?8],&
X9.B&C(P@7QK^XT#U=CQ]_SQ=T)QW]NPgQ^bQ=C5_XEc@U^e0TY\FPS/QR2PcXT6
ZPSZSgP?fFQ]\_IGc7T,dD-S3N2S#W#e]@;N.T\B\@E0L/LNT?BbGc8<D#MeUX#G
8\V?f.\e+=fefZ[eD)f.aCA/JRR?Ef1T/W_-=^f#C;K3B\>ML39e=5.Y<8V(48#K
+X_-?O]FGQE]C<L;YPa>>94_=<^J:<EU6f9,a<PGY9@:U;DJ>:ITc+J?eU=@SUVf
H/(gIVQA3eQ[ZX92Cc\\1)R?-GX@R?()&bV?O_E4R_]Q#W;5E22E9+,#>A7b3OE&
+2^1^OCAZT64SI;##&Y_O6MG#&MWR=W;T>K\?XRTP;#DTR8?-(;I6MgGV?[\WZMe
98Ee#IBK-aH>\;;gO_Z&OROUK,V297K^K,EPLMA&FR;McCAHB.7#Z0FMGYX(9#AE
>X12/SeR[NMZ(--B&f]VLF>^aW65ZW?<KGR4645C3#faG<L7[7+SB,PE(ScUDBJO
2#BGffTTgZfB]+I0b?5;,Red8UYTF00.dI)8US72;;&_(XB;^,F-\gL-B0_d(^SV
gTOZL];GF[XIX0db8>O@+gca2UL0WKW9HFbZX+UNQ4<a.4gd4?@:P5NJ@_S7S&IT
Xg&;gN_d42B@]^56OM78DB<JT^g)JY;V=bSEA0VUOQ9eOXCC-8Ag\gV-cdL94D(]
KB=-K\6H07^US-JJ(T?X>dV833,&[HDZ&[&V&Z39-D]IA/)Ib];BD.@1-IeU\RW(
;+2Qa^#/f(NB(G-FGDgU4N\f6O8K^?JX1d@)[T8DLAEHZHFAM7KA,ce5H#a<2;^^
fEVPcC8+0NfHQRA<-;e@>?P<^Y<6(;F3bEI7ZGH;dN3?QRUY\Fc).U:\G4WEdYL5
@Z&[)0CB6Cg[JM]5V&2-8e^B=V)eO@J1RbB/&PaO0#DEcc0S=YMACgGc&-[C&&JA
GIENWKd2>)J_KQJ=\G/)&?)fB#V0@&5+PD>@[4e,T795gcKO7XNL0K,CU/U,;1V4
W(dgG&L:H=2AC,M85:XS(:O\O0=T;C7.b8YESFMdHMWaC7(C/0KGPUcFZIEU8J#]
d87+gB:UFDd59#AdH84X)W1YUf\JHC5^<6;fDb&UB^#(/;&WWUV0#8TV5?W5XFQ]
[HCEA=>=6]ETEVY.7H8U\L2\2a\?E_K>eGF3C1>WI3-+ZWE>J1<.A>HK-(H31=:F
#H]R+HH[6+I]R@0<FR9(,=UZTbd:L[Tg5>-(3H>I:K[f;.ICd2)YU(e0;#@V2;HN
=>4d[dA(?>^DIa:UBI-.Y4_d8@>(=SUL:;bR-3c9Pa1>D>G>b/PLRcLMH)N^\MDP
G><^cdQN59F(7S&Va,XeCXJ-O1S26cF>TT,F59BK<@U:5aH:+Y&:(3_9e=6:,fH7
W.f1.1+5@0_N8<M1IOE#+aS<<Z^E=/8dB5+KKZ#4?N)-&:U^Ac_:AW<N71eL3R7F
cFLP5+F<,,L7>5[23^7^G+cY[?6-Z4DUfOSM2eBYE]c3O7b,=.37:8YT;K7,abS\
+#74&AUec11X7:f?EIUeJ+bW\7G^-6K)-8Qb;S<>0W6U/OFe6aG-0d@7J=-A[^&K
PZEa+MO7N>-,&-VHWG(A=P.7fN7:Ba.IPKa]CgG2.bNV3HW:_&F3]f=L+/PMC)XO
OaB[g/f]KZ)f1Ce_6G7/8S5R9VI+9;A27dOcK[aD48O<H2KR+/M_A@H]a]&YgX+X
FPW.eXL-V3\]/:JeCWB66KJfX-BgQ@cHZIKD^B:ceC-2d\@<^bAPa_FTcGMW[C[Q
f?U,QF2-R]@>HF;H/0^:XB5gPd_RD2d=gCBDH6X)ZO]D#=W?7+5UC?5RRE4g8VZB
?&ZQF#M9A^G_V=S3UN7L,42+.bQ)9_#.3JPEB55&fW0L]L&3deeg7e[WB&QB;10M
Bc,.C+9X<_X=#6QVVa]c3g@J<)Z#O5/)O=FQdIO]KWL0>A7R.A.Ke-4#3ag;:T1#
E/#83M1d&bR2dGH^(fC63_0PWP/KObaYMZXRB@[R4(D;\[LT>>QYdL@-?SJg2:8N
,.HWgK1/F;9.11V3,@=:581Y^B)NbaD0L4VdIRP)7<UXY8:DN-=I]3\]3F3]<?2_
)CWB_<DTIW3>OP\>LGS][-0/+=dSBYA-_<NU_(?Q3ABHI:ddGNcf9MYI;+Ha_UcH
I2:@@eI#6689-a<_&e75b)8[T9FE[\W+e=PD2gE92:IXSbcd9[1R[X9+f;GHE[f@
E<3)14JDX8<=M@/G&(B>:58O4KNO<d1O-NAe<YS_)N2HSE:#dL8+IJb>)(<fLY5(
gP-7H?:-RM8.+6QVDJW@=1^VIH].a:2X2/].;9bL&(@K(&@.I._:#V4SQ#DQTJZ5
aK8RSD_7>S_aEK:1ae@\A;)AB3]W<ELJXaf@Y;41e928@,/\gegR=A6dICe8@?.2
[OM:A-^DOBK&H&E>7BR=)710DHWY>]c@Z.KLC,;B^W@YBY.=-7S>3&9]R:^;M&0/
&_#LY2O-aHYX(-5WM>>10[\Y+#F)#E:<W3S1:5+/8&LUA=;<-7MJ=I_+.(N57c//
RSV#G=@H,#F2I[[4G99Mf-#.BAKTQ;(O)Y,9:M5YL5/0:0dMON,8IPg+TSW1\]9U
b\A;]Z^[0a\6&XT\0Ca&.0[)7\4D1/T)Yg]98.?VG-?Q&g@GF(H/>/2^dUT]C<g,
FQAPWW_V1(Mf9M6KdWb8g_YCU_M+TB:<(AS[),=,M&LfFKeMN=]SdVK\S+F1S,B?
=(,#5,:GHV5A/J-S>Hc(8@WE5#N=Z_P^\4:0/&\_[@gb+;BE-4)V\(RYN==[4/Tg
BSV_+]&>AQ<^e7SeTS360d3.9E>g4X]:f;HH51]?M]bJ9_S:MgA^,9Xd;?3EWg6]
aJ)Z[W:1;YZK_DI:Z(E-3S)R?RGQTV.W7Q?=&X,(;E:-^S\^J[&.]GNR;#ed8_G^
38;@AQ/X7eF=SBQXe9)O31f=/F<6fRcZ.GA_/<;CQ)+4NJ]XT-LP7+,ZePS^2=Jb
@fUSTQQ\OWT=H-aFgQ9#,@7(/7ST+\^^5c@LHXd?U3;(B>OS4FafaG\^]_B,,O+_
7RJ,-,dFEXfAL]3\g-d<X3WQT3Zg5<3W-MYQX4O;OeNa9;NH5P/-WAZ#ca,OBDK[
_2F/^AXE1_<K,_)UG(PeW>G4N8LAS?I/[N32d>M?K;=&SW-()WUMYYUYQ-RKRZdY
I84c3M8A)bf1IMEJ4c-2&[0CJb6H7N/dLTJ1>+N[=c<2@W57M,A)=,[.M19\&X)&
<FFbJB\XfSB:BF?X[XX<,Y.H[#-+2H=BH8d:1\9CcBd:>IcKP)_0N1fH^XCW8V(6
IG)Q8WDQ#NPQB7,P@4>_>;DQOB@QcEcS#HK5KY]3=Y14HT_VT@RODa=C2S?V#EZ5
ERBTSQRY:@M+;,#^g308Q(/Pfe=-R-fF[[]OMSBLbX^JV[UWeVQD\-.;8AQGb?G[
071(_cV3G90b=dXST7XE:.H\DS0(I]Sd&bR.K=\aG7Za(?F;YVUQbTcK7Pa29/3B
;_JTT@A:GB<]f2M33-aVf<2X;eg#g5M0S68g]ZJ<=8gJCf=1]fe\V)V)aF@f)49B
a9S^SSaV\@D;Q(,U:LJ&K@XTG_0XVg&QLD@e5#&75bO.6b#X>)5BDfg69XJ0);Fd
)U+L4IU_N<>F@Ud_>K.Xd][ER39b:NMb4+@OF:=&O\.A(W28^#J[dgb\8:ZQU:.6
L(S2^H?g7<,&g^55[0SOPA<RW(ba5KbT<6GHG.V/J>1GW+\LdEQPD,,+]0?XLP@4
3VF\1Z4/;2RX:FTG5(68Y7,6d-?cFGU5f;f0c>3MWC60+JJIW4:FdK8P)L<@gE=g
fK-&7>HdQ4,O.1QG?J4/#Y<C[8A-2BS5&N?c/;g;L+Kf.K1gc(/c:+e2&&;X;FUZ
Y5870VHYNS)(f?_822#U/GJCT4KE<NDg5ZJ.\,a?M0cBUPg-Ue)_d.W9;S^,B05V
E3])9ffO1DBPHM1c.W5B4373A=R9],3Ua:7e_.cM(bC2_8Ed+.2?.JHbc5<T&2OO
eU:?XO:bM5LIcX,0_Sc[EGe_?c+OVgUIb+TB<SHMg)e0]),ZO1g7,(FgL^0Y5M9[
VgXbQ=Q^8&QWBfQfV]5c5Jc(KBX>A[]W0U0>5P.<0=CGcRcH-44+K8WdRY,KG(7L
]7#4A\9P7Og-<XU[Sa@-S9NNd3C7;8H@)-]T;cH,.\R5gb&>M0-Y.U^8TS+#B^;4
[:55<K#bP8[gKU>b),O8Y6SGZ]SOV#C&KSKQ[OU+OUd=aWVg;>S9D0..F=/BU1)\
82AN2Ic6N,_c.FFcLd4)X)&ZO#VXMe>97KXGW[4=E6RT)FOS<5_aF.,\a[&/MKJa
Y/a]S535dd0G+7WMM<<g)XQ#aAc.I[FIQ6RP@?3)0EQP.,46+668<S6#9J<4JR13
7QW2JZMcM.VPXP36[d67Zd+5/e52:H3-OBVBH=XI5bJ&)d]]XJI=^NMO/XZIf6GD
D992#B=H4W7-V+Z\BU3bAYOK5V;c+?g/I4?e:PY](X8GNb1_5P-VI/H>DU>2JF:A
/D,KOJ=Pf@@@]KE/-+4L?ZR?)KWg9bPG1HIREW7E0b4,9MNGORZ13ITL-4d:\d>c
LXGQ#e7/I)_Z.X18YU?C[f40eK1DfOS1&)_e=&]5c(\THcJQbL&#/(FNH3P\#P[C
Q2[g&Z@F/:W?3d(b&ULa;aP2E>G5fBWg<R8O4@-O-fL_(Z2K8JaT\4IegK1ML4C:
9H\.37-N.X^,J=;8.@<71]CY@e:ScP)ADLIM2]g[0C5,KCHYUM=/aIQK@4IM,1WN
#OD0)#B[N6US?)_Q\dPM/E]P#f-b2?GScF6HP9cb<5F\YYgO4H[^A5EgP[C6bDD/
NRc1\O)L^?-&S7[4@&gg;8CMS5^7<,1N3g(ffJ=DX=9(O^OP.0-gdMc/B/Y[L7?^
XcGYR_<;PX>MK2QHT;Uc(#4;75L/^P#cWS?;4(PKYTXXKNO0E(BO?JDRSE-G12/1
Y9^F@G32a]0dO]3(JJ9+43.SFW]7+g39gM@+YEN-<;Z&Y&/)0b+ZCIfdIUWBU^^@
1A7Za_/5<;<egaHLO3AJD).S5$
`endprotected
   
                       `protected
,VN#N#L7AGW/MNUcZ>?^B@1bL-2N_<<A:T40C7/2ZZ7=F2^NXb&I))[\8813V.G;
K09(IFAc0F+VL&@<2A.(D84BWY=Aa?eIP2<V:\(3,K3g;P?a,76ZLPS6gXUPKD-R
($
`endprotected

//vcs_vip_protect
`protected
..We-F69.NGd=/[+-9NcWAC97PQE&Wf70K5?3U;^F(J?EgJ01_3S0(fS<478]/PS
=e/A\&T^@ST-HJcNUZN2.TQYGUGc1#Q/8P1AX+F_(a:Q0@S=]AE.ZQKFYeINc=@O
#XZ3SODH8]2G5Ucfd[&XW1I_E^TYQQa683fDK/bHg&?f=4MNJLXPX2+Nb&YPJOF8
OS@P7f_O+@?G#a8G>e??G4[&SI=J_Q^#VLL8\=^QJ[(/E;Af8-7IX_LODX1-GKg;
c?Z@#&(AWP^NUO#35D.P=T2fcW/A1dUf6&a(N.9HDVd+C9U@8@_]NIV]+)#N5UG;
I^H>?DZN9[30(I-4I:G.>gA2=TT59_B4d/Wg>[/&8GN=8BTR5Fa<:.C@@.I/BA,S
37Pg)+</?6)Ga9TE[21WdX6R++2gK.<U/G5cFF+WL6M@DK1)]CBPYX:0R?P\/KV,
X2Ve(9SR]/]H14>aYJ3:S5a.K(GH-.?1T]b_)I9COd^:(+LIJ4:TI93JLCb>WS7W
-YGHa7acE8L[<QWN;GLB[GT]#6+,7RD=;@7:Q[KCKZSfQ&GPdDVO8,bS7YB^L5&?
-^&NP]Z^@AE<7@6KJ]]^O8Y^^JTPf?2&eLE6<fUf18:X@U>2b,T:D]M:e)@,[1,O
2VZbF5ZD/Ne4=W6(,#Lg<VcTD?Q0W]D3EL,HCB53DMS>6H60XE@Jg59fS,5aY:SW
>]I1R+J[1;g;1UIWd+/WDDR_ddV+Oe^<d=g0M7GXWO03K/W#/BM7GLeB@bR78aS4
X2<.<BSJ(bMbC2Tb.>Y&EG<;CFR,YGb2Ad-W5G17<.&NB(^_AH@)HgJbL:bICC7=
;_3OPUIaJ(eQ5D-=KD:D1^=<Z.J(g>P_LdSJe^Y:SU9I_:@c+WU5U&Y>bd34?J:\
0fcT+J@E?gbfH9,9bR1H)&A7a7:USE&E8DM+V,:#fM:VJc\_.Y9/WK3)b<V5eD96
),Ng<Y?,<-9@2J5_]<J5fL,-#5:6E3:OOYMa@@WeaHb5Z2VEQ<d\\^d/)bKG6?Me
0H;3\W:Gc1=XaaFQM\KZ/[:DB8K.&aOD)cR<E>&FdUQe:ed62IO:+T(:AGd(E>eE
X<^OMV[9,2FI-b.Dg0?[[QaHLd=6D(_G,<^FKE1N?2Z7c:TQ&dRX1e(6c7g-_A9Y
UQUId:bCa1C:7MNA8CA_GPe+7;_&fC(HMZQP.RdC)[A8d2J[YeN;]cAX0Y.QN7;=
ZI-Ob8QV@2&\5C(:Nb[\eA8^Z;?4T(]bD_+OMbCfMXF+dKd)5H:e<A]FX/R(7K:^
)c@U4OMe09AA6dZU6:JV2[/=(D>c>]^H9PHeXaR.]Q7d2EB@FT>SM;,\BW\AHV&.
[P+3^cV<DWe?A;V#g^O#4U^[F.9<P2K&c>=ARPW?aSL:YTaEKP@(5H?FF[(bT4J1
3OX&BO<@8Q(AbMf1<AIb\ES>IdbTWE#a^NBbDYf,d/K+P3FTDVN,O82^147SgH4^
I6+cW@8N56,DN3QH5P@JcP.C[&6U&<FMTCOYcNV3;<NGD.\L#KI)aB__D\-?G68(
3-)NK+\Y]9)_)^?7f_&<E72eO46Y&ce(@:;4ab9DW>9VX@:,J(DS)(F>MIKdX;a0
Q,:d,B:6:1_Jg[FH;5=UGfZG4b&e)G#:+V;85N/<^C9/7#1RG-239.-6GQ_PW;KF
MJ5@-2(+\#)=S^GU9TZJVb:_.V>=6EWW@_Y##NK(BJD8&dP+YXZLP((.J5c;c(2H
#86NaC<1dM;FSB3?8]0F@D4e4NTP3P/SKV\80<SXF&4cPQ,:f47=@YTag_Y)=f,.
F2J9M=^9+MAFP:<[,:Y#eKVda@1?f>DX6dc@^3WXb;X?A\M1IIPTX/),_dXI?a0(
];7<3V@[0X:#\^:V@?YAD+>A<d>-=JdQ-1?@CO/0PK&>;(AO_2_#K+>a?/c)\X1L
+XdY>#g^V#+cUIPB2@&MH=dA]_SYIWGLgEYHS3X)IYBET5ccMZ)XED9[a15[>_U-
?f?c?JD@\1d?)_N[D)7<eD9GPWg316FIBS[e@(0dU(+QLDE:=fWEWYb&g=.ZD=;P
=W]8PgIU8aeIbfTB+C2/b:Z)b#BIg?(;dTSa=,U13Je:>5P)9G13<Tg6#edZD1NC
B\Z0VOK.V37J3aE+VS.S+0>>?5_@/IbR62TAB5]V^@M5KbRW37F29+?A]NN&[?LP
P5I.:JR]?^0dI]5?1O-eD7R&+S;?NJE,dI>0RSMKMFGB8&;1>g]1_M4#XUEe/=E>
^(ZOU)AW0]Gg),?7C/6_X:M:fWR<b^E)Q+(S1^Y(39#_IY)WEfIAg&(f4aG[fF,6
=KVJ#TZUK48LT_2WZIf1^E^A(=):<]H0XEB&U0P8)S97R2cX>\cFRPH&D=ePF^FB
^0_^U;FVHW)?EI?;g>ba5WBS^<)C1F:P(H/7?8HGPVCO);M:1UW1:g3-QLQDSEC&
(H]WZV/&Z6+3b4K68B?B3_5]6X/)>5Ug=/f^(d-G;Y>G&ca)e,BfLRGI18DV8H44
SCZ??3I?.+PK9M@VT09eMg[D[<#f>[#)W_9>9M#Q#CIFgK)g1WM-CJ<>=):X3^M-
d3e&NU4P^N2>MQ>218;3KH+Ee:T11GA)\(UKD#XJNM&Pd9/,LJ7?]d29T]1WHB)g
<:O?F7IGb52<E]FW8f#PCC0:?JfLBOA89dG-X(F0PO)D.YPE_9<,8@e]/QNC1Pa2
C8@LVe/Z]AF@1(B#]Jb]UPNBcY5KAZJ3N/(a>/Z7]cP)-AM^:MQ=1eNG62[E:)Q1
UbK,;5B3_(0CDMR[]&0R?Oe0(68L)VS9b#4<:,OTAaO<8:+58bJK2L5EV7K@/:DK
).-9?ARC5#[F/U&[EU(VRKCg-F[/O.5PZB3M\Y+W5>a[2H-?M,B^A2(aA(<f#TC2
d0=7/&@7:RW/O/,;<4ACKd3\@,AO>=KcYgH;1-CfW7JU(BOeY#:WLV5U/TJYX;=Z
:2:.9B1KY?)UdBN4C()]=6KW<2@\,6b6b_#3CMV>7&T+_^Dc^=T9CSAL88G]Y[)g
73N8=U1PS_:dU6=9C3:S(<51cg_:1c:F.:ZS:Rg8QcBQ&J/=/T;Y/c^P:BGCdEIE
;XK<9E&,T36&MLAR,4d7+-5B](,ERU(:44U6VgT]FO<WEYc[/gFa214@9GGI7\BL
/8C:WV,-V;DD6ZSe^-^DZVB;H852#5?(X<+,7O@(10:fPQL4@48WTCC8B)A9:e4O
SW(\g(Z;N+[Ma3^WU#VY#3(a^aL6N,_)8FE&:eFB5^?.R-/R8#Aa+bE34>]O#[=6
6U7:aXgXKGLd@/?b:,+YR/:gD3eRg1Y?aLIfg(\f(L=9ZIZTLJQ=&#>[US.QJ/e8
GJ\O.g+LO7HM_N>eSGDS,1.b+9V^=1FY6/MN@&-Vc)K_fN(;Lc]F0.@1H)FPTWWf
BXO_ZWf.+\48@3DM5?F@ZEQNI+X=[5VNXRA&NB1;1.]&;P-Q,A.X/(IVH.a<D\I8
#X.\RST7;@O4\.0LEdd7ZeU1f1F4+N0CS/6W4+1SfV2NU_AJP#g+A0GD,/DE#^UL
R0W31@H+MQJeLQ5V1E__U)b_<@+a-DM_<gU4aE=W.S.=Q>D&&X5QC(X0C,LWVQ]B
384,@:8-4VdN.G<c9#^J)W^dD=E\Q8CPecN\5]dg/(\C(a[9>F7Z^C1T]D:,J9Y&
.7e0Dc&d5[>Z.V<);V+J]V0]EcAXNG5+MC.T8H:3\]]=9X738RT<=Z279U]B[<Pg
CdR6P_RG<EJHI9XePUHNXU,45cBcR<+JIK[Ta5Yc1JKccI)X<KQL/PM>A-/GB)OM
/d#7(>C:?6](L_dR/+J>.d3,/ZPgg7D/60J9FO@c/_EIL_SKZ2YI7;NJ(35\CgaD
.NeZ#UI<(1^cNXC5YX;LJV\8B==KUbed@EDS3ZIa3_eXLEXM.ZI[H]DJP(;J4)cB
F+25X_8&)/6>-H4+c)+^=/<V+bHQ[902,PfQ=VR.<Ug),:D(bSEQQa=5U,5F3U?d
&eA^>.@#a@Kgg=UMIQ;7-VY3d+]g>b[7?=9>G>;B#56;FN,=eHbI=?LEVd;UWG^7
.3eeKNT>+f.P,fIHL=:FH3X?4]<JQ&<V[5c8fb=JUfI<:AA;G,gD:N30,7H.fCbg
G7T3FUX34LRP^Jf4]/dK<WRKC_]-HW+gd,Uf.(/)G?LI>19-S2Jd\53@F[71,^Ie
_NWX;+0()@QD::LUE?2/-H66/^[(e=+#aFTVMCZ&9-fdB1b,4Qga6Pf)IbH\(T#N
bLOYIIg=_gQbL;f8?]PWHATXd=cQ1[FS>D>_Z[Q;R^>L90E7X;A@6W)M4@AIE1ZU
1IAY?Z=RLGI9>9Q3Q20SSXUaX-#dF=NNBfAG7SZ+?H/QY<^F9UT0&+0/a,BL4<[?
;Zdf.GC,Agf89[8>7^/146Q1Mc+SRG4[.[.ScW[UNNe<K,RYT?OT1SE.[RJKDc_S
Gf5YB:^ZYKg=GZIS#+&2=?.]b_D<NX;<:_C2XF.O^\NK07I#))^UW&dDe+ID=Z6:
Q9-0(MD8EM@d8VNO^_PQ8-+BU;@>aLIK.?#RF>:-)YM9NN:B<+<c77P2@4D[Lbd.
7Lf^9E8(8;ZROWeQIZ22C3K+;9?.J(#LdXTbI;^S:.K8,_0dP,O9KE.7g.bcGGO=
,AWMNS_/VRT1P\<>I>G8#<:f3MGFe.\67.[-ZKMSL19QOcRI9NPQ5c82>6-W5[)>
?W9S1_G4+&3@>E-YY(7a#1,PPC12S^6fIEMaMO>TL^H?N?(WXW3;=df[Ed6J/de?
MXJ7W9c8I6H(Q+6<Z4Y,adR;3YI#TbU@N@ST6UV1A0a-3<(;Ha)]#[N^DBLab^B4
\?K>+a7f0,\HHL6_b+@TeZDKIa/Bd:5KN))5_5.=V7W7MI,4(#^+37:B@89E+Y#]
HUIb/C;fU-0(D?eLfR8>2BT)G]:J;U]YdODAS:JOR?g<5gRR]Y;]R9Te4T,AH_)I
(@:LRa5[.T/4O-E3&K9EebB0&;JIM?Pe.D<H/E=ES8OW@C?:-LeX6):g]<;e4-IO
LX;IGD1TVX6N6I03/Ocd5QaND7_d&N>0\<3f7)_X]3bc#V26#-0RfV2R^eKK4+DA
+9?EaISLF3-E3ba[-LY:e4+dS;6f/QbU^S->32DLZ=,8ZY-+H:X-#HSRX?dJ:d^-
\BQH@@>/9:-._0]EPf\(\=TUWe^SV/XaU6C0/;=S1ZC.W<Z@B7EPL>]V-?)23^WA
[0+,4HT-Re=a-/g..eJdA#;@H_W(Y&=2WY_2=AAf]Z.73FHb[[8&.(HXBDCYOfWf
MCOcD8E0Z<>(Ecd/Rg4UeAI10:2#H21]^aU[)-g_@,LU^><K#_M]@EebdR(g0S[/
:)d.U62T.BMT#,?G_b1VcG(5>aa8>0FZFD_Xf4#?TOV]&gWGMb9BeBZRY,aUB&a9
g7;UaAE@ab1GZH?5\KaHK\V8PN>DHBH>QD&.><MF2WXO3Yecd@,2M4J32^E=Y134
[BL6GLE3BVO8,)4K/GDXT[PPB#XBCHg13HEaW0BfXf>K>aZW3[?1fWI?/BCQ?Q0L
>(;+\bAaUFWDTL\]#FNL=.V(C<:[<5Z\HX;b,J\8ZR,V9;H<_=a^+1FeV,9\E4BX
L#(cP?L3UKLSF_(c=/LF/7H#@0E,=PTgZ>B8EUQ0E#:4,CY5R)4@.8_K>W=II,3I
][d9aS[5NN35<SC)8S,C->P6^K[-EeK-_gFg#/b:A[4.^G37Q\&\5NdY^QeVE=.(
DF-Tb7.:20f25)&/<AVB1Rb+Qd,^?P>a>7KOQ6_CWN#Dd[B^[]/8)WRV)I+(+N8e
.>.KQ(e67,Y5M61F?X?)U;Cf&FO0fWg#TPV.FDV?@>c=EJA2daZCRf6Y43FH51H4
I#NNg_5b1_G.J-)K<QW89VKZSbF>R1<Q5AJU/fV@PO,;>aV/YLR<RX[0^J_/PDR8
gE>=B.DCZ,ZJ^Xf_5aDG4\7NC[OML4LUBg[cILceD9Oe44(W?=XGY/L815:HRADR
[&\?N>E>R]M1E56=:Mb<NF@a54dPF\X/O&E_a(I]UY1b;P.Ja6cZMFKB&H;b6KBV
Z?cK5V&I6WS9/1_+?GX+Z>44.Z6:FQ=;Z1453eeF(RYE2BfEJ#>37BHTOf6R94-?
X,/VK>5LEc\BV&YL3eeU5@4C_[-P+3LH1//(Y;42dN)+.=KJ5=F2G<6/<G>ed[g1
AJ_,VE3R4/,aCR7(&Y@AJ;1+N3Mb7&6+_D@O.3]d-dC&E3&E^Gb^Z,X-T@J7@E59
&@+RQgb])V7#B[U7Q[9H,-YA8C(9VK=U3e]NS5:(Tg++8(LbGTEIBQeS8adTS]0B
R___\gDY\XN20XDT5Q<4ES/bFA99CfXSHPYS1==b]DZLFUZg0J(;)8XdVYZ8,IV=
M1)V0M.]g)Ub>[d3gVP<X]::))J)c))JbgD]X#L3H8&cRaFNR/8\D@-YD;L;WS(O
Q1aJ/:1=A/?1:2WB/FI88/HL+aC5+bUKf1,S1O+R5D+g5a>R_EPMC\N7(#c_c;EA
(N;A\WO03f.5+8DFM-\MOcJ[&VaDCg&_E85C.+65[V>0/9.WJ1OHFY^8+WV;X180
T89^>c>e\Z^I:bg3e#-L:5[DT&9HLX-E\Q?+gTBUN,>#MGA3SWY0,:8D4MEaE6&6
e16WSOI@-S/;:&F1JN<#)YY@^^5T(WZH)FSQ8g7^(SBPaf;:MWT4FDE]<4UCW0X/
UBX6S,H1Q>0&L?&Wgd[5Q.Q5YDfA-97LR=c;EJ]bK(50.-c4#=?G,/ba3H[3O(F-
(FKERY#G2Cf#+?8O-+8-9C\ZYf:,IK;8Lc#KY51>3ZCH4H^3-1&1V?&f8B)9)Fd=
.\8Hc:b(?QH>X3&=_I=X_>g5Y,E9CY9[N@A1;M\3O,LTb?3W:D:J3-gU8Y?&E0g]
4UOg.g>7cU>Cfb\JcVOdg^LQIbD_HJ#@]H2EgPCGO0YB[G=D?O34UaSNN3B#4a-.
dg=9\4<8Tg<=7.V5_R_UY_XeSL#KNb_\MH^0:XB]@Y)\6ZE+Y7A?SE2)OX3T-:\&
U@86/0UCELg2P#-R1750&UK;.V=>16K1W1#DGMbe;gO^@L326>JJHV3bT;AAYSG3
-LK</B+^4^SP9+27:MKb^+:<?2+c6.K+JIRd;c^8RE@40_:/Ze&Kbd6De-K9.,TV
8=+I=UIf,ADE<)2GX^ebQ>=b9=4I;#8O6^:Ha+b=gMS2)^OQYW38MMJH/;+R5]P6
0&gE^)EbG,OPZAgCW33A/+M5<^5,YK/dFO;X,1\C(I>[W.G7>.@>V+Ddb.)<D[&4
SL:W^W^=U?PQ0gFS=:W4b0SOKf,aGX3:R#XUWW_0)D_LQ-cE0URH3.A=+__REaaU
8&^]W>O&7ga4Z>3:,AD:1K79&[H=:\gBASG0dLU8,OD8)Z6U<_WL.V=#VRC\(-BN
+>Wa3e0g_IDPWb0^bX1^(c0Jb&ZG46D^e<U,Q7aLeB-3A<22+.LGT0;WZP=&+R@0
W[(([[87>&[C_^2g>a1UV7fWRPDfC69c\O0>EV7#c-JPLE]+\W2We@^C^d3/U&HV
Q;UD>LEHXGYe,[[2O61X/cE)I.f#K42f9fSQ-7A?]FE+./G:P40)IFEI>32FOX^g
GQK>R0)8&#d;,_D>4K[F4^;OJ.Y=>9fL[GfNg&:+#G\<?/1b[a9K)HBKNDG(UZ/+
:JUL9bE9e@,2.Ie;CM4Yc+O:a\BJ/J0_cI/@^LZW_b@2.PDDZ-QM8=f9#(EO[b8@
;DB>=ZeS4eeWbN#TS.0A=\242HC,X#]7=5XBLb>gQSBSK6H9BC_L_JT[BS#E5f<B
JOFeT@2Ve^QS[JcCGZ(U,6cW>21T@F(<bVL-C-F0K8c/4NBZUC7].09D,cV#:]2L
A\,)VWF1K^H7K3,aLf]]0BII[S[9U<bUD^Cc0&U;YZ]D]QHc#3\QSdJ=+U_,@59]
N@EI+#44^06MII-D\HPM=#:=Ra5ZG[G(4;W-eRCJ+\<;#U0c:G;21))NG:S(#_=I
F?.P<e21N5I1ZEJ(_@gT1=DX1CZf=5a9D]cSF[;2M.PgBNIYV+?(3T8#L+fWa6;[
195(P)=4X.8Q9<2\YT):C#76I#eKLfFfbb.7[f.Y[JSeEdC30Z^XD8\bT:)P6F._
\Y2]AeVcUYV:T4IR1[G/Z_BNG-/_;;T+D_Q&2HDc;5\d1J/(_42/\L>,K(/,UJ(4
37//I/f-99Jf08>eMD[S9\MQ+\_CFN5+d3,08X,b-ER5[gK\=4?/2DQ]O7=.7/f,
UG/-/U.gRV94O)95>D0_]eF7(.;1?,3F)3#&bW\VWE,a9V0O3Gg8]KPdcA1R:-4#
KJ/)<d5J>R6<aCX@b6.>KMO8eN&R0?IYR_H,.0OJMCB_D>ASI^Z:]BA3IT5JMOH;
B9LG1ZCG;Q6754O5DQ6HL;>(OFET4ZQd.C(TG,>\2\fASe)(3@WHIA<K2EN.;OQ\
2Ba/RO?5@+)][LE&Eb[3\DAO0f0DAEOWR>D4B,07_YZS2g_7VR/4GXM56e8<<Aa^
+6NL_J3R&+^(5BOYX5GO=WL2-AKVED,8&L.9K\?FRZD0H^bUUZJ^5a/e9\A86W6P
]M&:IP6e-fCBJ94QVB@D,[Je=3g=)XA&a\QVS\#)63^:;MY-V=TIC6#&=U00)CaB
&U+ga5O=S/)F<ABD=E=&)VcJ.^^87Z>2^e(E>JaG.6-aMMT,gM@TJ)L#?C>>Hc44
HO67+?ec;K/e/PJ[RO&]-H<3a@G4\999DQ9/OK,,[dADLLR3J7,+QSMMD^gBSQML
H)+EB@DSgYUSYVS(1KCO#BDW7_GX5fC;(W&A+T5<)(Tc]8+?I-?B[A12]\@_gW1N
G@:KU#:>BV(LU+MOdCeA6-(I.5W_^bbY_QW<7MLRT^,bbFX\BIL3A)Q_A:gGQMI_
RHA^WDNbU.C\N@TN+S8f[(NYU_YKW-UJ>ROXA+T6;7&3XXe69-R4XXD6-7SO0KLf
?,6F/,\.McX;+fc4;<),O0bL^.)b9R+[Og/a/eVGC[E?CbSA/YfYEM3E_T7>-@X#
1-F/SL&2JBOE:N_AagS&\1=_8DJ)HQ>NdRW.I2AZDC.?/NE.SV6M-LJ8.CGC3-SF
;4U5cL.&=a7=#&OU6;BQ?W?OQ=:gS.P2cT-SH:<ONCK(YA6JE-J+T_O6[7SFHMB1
=@g66:Y3W4.?EaK_]&b?_D]TOU2a0,a6P>96Qd]DS^CbaC6:<J;^FFU#VXV8Ic[_
f(=\B,J1=^R@33+K]gdg<3>fI]Q?(O>G-<RW7e?aTMU8/6?#C]XgdQFEP_\aF16[
2d#J<IcL0OJdfc;^GBN/O@N8G=GMaU&W.T9#5G2:Bca2A42FCa?8++<DA3>:.X5<
/9.b06(1V[MYV06&O2(0<P,->NeUG/YU0F9;/3<4.&Ff=+>UMMB/&WLdGN2>7@KK
_-)7afcD<[3(W=S0H95bKA#e[CV2fN\[c7H-FUU3O]\O:J62/IW6d#I29HaaNTF>
K^Be9&7R1P8fCS/PcH?D6d#G/)_H3_Y43:MD57.314HGdKAN:(PONe\KO,L)(DE;
?HZD[,,cN\#=Y3C:cI^P5)@1@ORc3)0bH;dY2=aNb4(#S1Zcf/>G<7S6<GaL@?5S
K?H9&.g/AQ[#RL/Y1Y>UWIeLaDGA)<5F-6+TK#:=bXCf,&1_@/J&^^9+T_cVAc6g
D#[7d.JM56T5cD@.Ce^I.7-JX.,fL8HK2C^0Uaae--I=?:^MGRMJ7X.]EdEH[f2d
I1gL+gCK54RX@5,-.Z61JeYgDB/6GOc;@]2^0F,bA1HKX1YQ=d5](BdU?ROD>#9E
Q3aS46+,&PW4]cU89>&8d/KIP1>;L/<H._G,b>P,Cf7FJcI9Lf89^0d0aFUYP9H>
g)?#5A2OBdaI1XEA:g[OZ1M3@MC(8fd@MG6HQEV#c046RO0M77<EDCR.T0Q/c^GN
3?c1YGbJ2ZGN^Q=U&]VKG?++/g8;0gCFRZd0>QG?:GAQU96-V,M2KRgRV],>V#P7
2N)38)?aY_1:d[eZS^HSOR#3e-P149U.F)8;H0<A,3[c#SeQ^VPW>fLB(13>VE48
94WYH>/C-V+^6):6>PdAAR2JfbbJf41NO]ZBSJHffgPN1J6Pe^Hc0dZ86B5b87A@
]f7D,BO8O+&H3g(:HH#(;V-DI73e+0K84O>>(>g62dK=g^NA4MTd9)dZ^E9LUGH0
Z4CQB9d9D491M/d06G(^+-g/@[N&HA?EHYC8U+@(_cf+TNe1b..c89NJATYO&S\1
+L)8J1/9YFFX-4&0^3AD23-OL7(^SIV+S-g8450TH@W9Y)0[M+K>?U.1eC00SQ\Q
).X?^SfEbFP]OJf3,Mb8WeA[MOFV]e,(?a\7,5Wg<_d-Y?&B_#S?M755T3ZJQ4dd
?EWcSS]6J]345(A/YWe0QaDSG1N^]UBRKa^)KUc-YJ-F&dC&g]X>YL[8XG150>QD
KO9+9e#0J:2WJ&5DU0J=eTIDIM;RR4bXO_AAcJI@40HT2+:B=W.GSX0f)Z>9J&Sg
0aU)K>\=gKY2\62[gbe8(H,)[T#@89D4:gJ9ED(2E5EQYUUTG7H@FI7(c>^dMddc
2fW)51;GN?O4?<(<.[Q9f<5-SLOZK7C,-eN2[.)42I#\>,^C.Zd.^1f3WCd2DCPZ
/5ZP/L1MgQdSTab1DMYD&/CAd_-S.L-C=VW6eO@GeH7ceX]fA4V]bD)3=b5b#&I/
B<@)\IeV?9#DcZ\ZffJ\b1Be:E#VB:1XLB(_B8e]5YHA1WSV.MKIP2aQKfR]CC#Z
DA.fS0E\-#^U63a[G+JILYgfECS9NU:H1aJIU^X:LKR+?6NT<I,(Z(]^9^fV2S9_
5eOCc#gOe][-TS<T.NJHNJ7@\JKQePJ49a,BFEDG\MO5d2K#W4M1=R^c.0_:N^5Y
9#=1;#AP3U,3#\Ya.D.H6=&/g).aQDOX#_2eL>E^@g(R3_aC<R141LJGcEf.,O4_
((52fO6JL6[2U]>.:?PO9X8)<d?LP]B-4LCMU2ZA?/#Z6U>@EE59/RCPNCG+PZ4)
[:CCYR]R=:g]\LW[WL[97g776c7=ZCH;N.D+#Da[,W7Lf_/JS(ZWf@?9+.(^B(QK
Q=ada7;M)?S:#/I#:d\M\d[@e3a@7^1]#.>7BDLJ]P^0(A#fcII)@P--ZF,CLgP:
7.7E1cPBcF-^L_(3FB:D(R=>1>2(38Ld)@Fbf)V1E6S@^0392cP?#Me@2M]14NM+
[JB25/5B9+_[S)/H^+M7NL,If4a768&7,X,fgG/Rad6PN_J15dAd=JcF0F[6+Q9Z
A5V7O,9?B18aQS2YcPO_;#cB\BU,a;)#_APV1#1DDB)UQ)R6RL45SeRJfZ/0^KMR
\R\.0+T7+>#Eg#_c?,@S07?HVG_Kc<bYc4@<Z.3-C]e+V\;^PGE0Lg=U1EO?J?&Z
g]S/(HCaG?KSC[D04HBOHgB9&#>7TR=HI1Ud4Rd]J/gN<?@6bD5JMBL3FPIV5c-R
Ra#.D]I)21c^#d)dAOO:U9(Q3:CObL[_>F>]#5aaM9B6R((#L;BC(ScDPC::3TRa
+NS33]Zg3V-HV8(E(E^K8db)Q8N(L=(\M3RR>DVBD(^Rd=3VO(=90dLJWL@>HX/@
+_2V0]VcXdB(cQGI-:2OacL>\(aCPPH#c:M6Z^7g42ZG>@D](eZ6_-+8MBbO^V<9
U[\GS/R683()-J:&=XCW<SMaO>8M:(\<Oa)cRG+R>#C)GCJ5dFd=;[7P3c(b>@L0
SBCYJ=#=YHG#)2RE5I@>C_c);F?E#W)9Hc9be#\MR3H:BZSPWV-8PJ,OF\13c#_4
>=a;&4I\E>)6Hb[H>BCO2A\JO^YUIJEGd.+,VgZ+JW6-LO:/S^_SORcMIZgY5A3Y
8C,-94)YQN:B,XSMb]659:B0WVH+#7V3[1R;,P.#@&f]bfH;O+#+cdCMVJ/<RUfX
0/M#WBG06S[5U(_N]4F\J&)AB?TJPL_)/3)9RH_#?K)>UOSb,cUJecD<B(P]VgD4
UXN4g9bOXGF<GB/+<:U?.IV:-U#-8#<JBHWJ^V#8.Xf\B)):3Xd-cMURgZ,Y?&aH
#d=M+SQ,6a/G]ZL=<_B@?A]GFHCfeE5O[881;Fg5N,QUC&A#UE&3-O,AC8V)C5LU
IUP+SN0\-NdJH>R#K45/.E1USU=2F[bK[4;>^D\\>d@M_F.0X1W^7-/Ce5J.BQW<
V\_)C6J05?)0=)>F@EGN510WCK<8GLcU80(N:g1eTd.1O8gV(YEK#,cT^CMdER1W
/eG<PdHg)fbS=^Ha-H][9\X_Z@]38^J=?SOS>O9g-U5f#D2TP68MXfM9]T>/?bM7
,08OK&/]8U9_&I)JUYRGfV;Q=eZ@8aK0:APMfVES65_H[fD[V_JW:4QZEQfNb@X0
_<+8f)fNM_##OXcGEAL_@85=,_DV0E+6Z_J+/1[#Gb?G@(YU]#:B9\..QHCF([+2
SgK.)>b[:88._([4^g#Z984Y3ebWc:.+0./OcB:(=9M5Q&;^-U,AaSCHVMF.R>Mf
G5CSb240//:55+#Q;JCb<Xd@Ne/&G,:GFO)1:M,(S:/\HS3aUA>VfT^ScUBR/JOI
6fI486]4K<GO5=Uec(<9fY@GZY&ZHK(2:ETB(W:eCUTP]#=?X<S(aR=PR]XYWN(I
L\)\d[9c(^[8R>^dF4K_:W&C#IRgXd27G5:&/7/bCAe5N@J.eH0J@ZZ[67J+AJFd
ZWY?IF?g_gHZcdcJ,g[TKB09)]Hd7eU\\b/3f\c-bO6_HZRW@9d+;)OATc_A=#1#
dDcR?Lcg@WA7eOWKD_bTF0TJM)^F]QN:<GFQR/fBgX&GLX.fW1TNf===+9#9WSL1
(/,K_T&8#M.:L5V9aE;+<+(16/(3QF.P0\@@fBb4-00[SER6dC(T.c;CX-K9[SQ_
cDASF96F+RTK3&+Pc4-OQG4F)UE7W98;YEGCd1<Q\b3?Q&U#dFE<D-:;?\K^6MSU
;DC9(-6^>,84O<<\A[aeVUB06+Z.JV#/YefB->^#U7LU7a2X=HQ<FT^(<;93ZgF3
5^c-,KMZK9=FQfbUID/3FIS<4RbdRb+Q94D&Lf-G>&45bH0]4Z438^fEMS/YKB<W
=M:Qf@UA1:11:>Wbe>Q-cFDbFI+C.2f^S6Cb@D2&GM:C9_@+2dCBS)YS_E89]BV-
d<<Dg>]DC;Ra4WaSIL>Y+;K=aVJ0XF#<>V<--\WA1#MCWcL##Qb@8@/)Y_-FU.PT
QfTAELdC2329a1@+QId,A78WOVEYDK;bY[2OG5#-JZBC8g0TKaO>2T>fbU\NO=3)
3UdNWMe:CWI^;,cR5[1a.<(8A[W94UQCUFT5+a_RD\6RgN1.7U.I+?e=H.c]H+e.
@F9U?S<[@B(efMeOJ#_F6G[I+S@Sg4FgQR<K4&#T>_4M+f_IVUU]Od4feZ_7.:f1
bR)C/6BN0P-8E8YO1ROaU:]<TaPB&VD.7+M?)^/A?6-FEA3QQHZ1a6Gg0_2A<(+f
X:dT3GHL<AH8K1\(O2,^.-_[,-cID-.MT\I=KV=R/A+<3+Y@.9J2[4]CA56VU4b5
BFa+b[U]K[0D).9[PBg=d=(aJH9<;TDF6d\XQSNNR3P\(dM9?FFUVSVC0UaIX[UK
?_G^<(B;@#=AEE&51=J2]ZYUMS:176AfK/;Q9)agA)b+XC8.GWG6_gU8)/V1_?4.
62^Tb,C>0g7R(d)/d1B6YF-&([gL6H0ON89Cb&^7:dJIKD(&\ZN-QBI,dXQDa&e2
XbU+8ZHQ/KN>_F8)7OL2L0];<.?_95Cd8P<Sb._RMBBHE_4bJS]=9UM3E.cJAY/:
QO7aFEX4Z=cV37.KJHE3f+AG43)?+SL9D469H4DagZ&\=RO37f_)G)?5T(J-9]H+
b/0RZNX?53(U3S2RCT4>FV2K>BS/1)DQd@FfG=9&Y^.J8Y(.KYUIXY<0GK<QYL_G
J4KFY5<d?We1)SCNUY].+a;2c&KDIQcG&Ib]_NI0dbY<1/]=YVa[+SDgdD@1cOfA
[_&.Vd2JPXZZYBLQ,R/JE&=U,?729)58;@..90]3K_LWe^-XD>UU9]F^VWb,QO6U
DgX_05/O]/aUaU-8U?^fdSR9GN/]16P9+<.866PEMTRc7b?:^c(B0T@@L9;,+]6K
@gb:V.&16]^;<+\X&M1X>Y+-.8H:#QNIS1-G84gM-K2dCa._4O?MECWR(+9MFRHX
f<>\;C([\PY;=3U-,.CZ@JL4A&@e;eB,JJ:B7?Y&D]-\aW9S[6_3/;W+Y_.J^O\,
=ND,F7JAa<QSU)B(a_;,GB[5;L/Q61/CR1a5a42g9((0OYg]e[HJ62@4E3,_S/4g
a;^RE,5N)<+F>GCMZ\WCUT]<]UUf6b=HQ0_@6E/R_<X+A&T]AK>4gM8HVcTDgF+d
b/HgfXA+.YCf/Y2L)K9Kg^db1@O=1UKD:Bf-ZB5FS[#C5,OOead_=9Z?#gZFeaL+
03eZW-JJJ]1G=@(8c9@,+]_+5K120D_(4?W]CQ>JH25bOfEC[He7P0T0GU^UbQ<,
BSJD--)+c5]>@9AdZWWcS.g)PIBU<12ZVDFTVHB2.f-Rg^FRSXeCa9<2@OX?(IZ_
AQ^>-Yd[?:cS6Gf@7eQ&Q#(?TcN[Ff7:G9J_;3SL:BI_.e5@UI>LfWCY&fDL2SFa
B+XM9^#\V\=;?CU6&YR.:<=OJ_AN;:_^==4/EO?4[&(F?77N(MV?gG<7@NB99,6R
/-eWT2L2DMFWDF@IE>(OJ(0)f7]]U88P,]7XX=[VJd:?]Z8X/D]Eb+9-I,UBK(D+
a8:;cF/[@3ZT=7,:V=KMU_D?9-0_?Q6MMIEcJ^Z5T7HK9=g&K78W:\)UQ8Y;@]8J
O?.PJI^64PYPV-\YEZY0K24.Ue?@9T#,^+[b[5]a5S-;[3.^CTcBBf@J-Q#,@KBd
4Nb_A/4Pb-b+2-QXeg,SDcOM,2L7E4[#W;K7gD77^CFD(R]EJIb=>?>:#E=)CJCQ
X:gGQNN#Z1@+F^^]g)#;=IG0)</U3_\[S87/JV.&FeBVL4Y#/Ib\\CDF;6]&L:gg
K/aCP/N5Z48D2EEgH:D1TFZV3?0K-bX7XBQON+dMa86L/A0>X18eGE4<Z0^?fdZg
1Xcc6:]d&743+?+,?a]XbC>.O1L79TNGd-]\-gdPE3V7#;G/S87QO<<<c<&\IB>5
.#aC23FX:b9ZLf,cgX44FLb5VLNde1XT.OGaY1[:Ea7>9H_8#KG@YSH[La]f@GES
MHG8CH3RZ]&HRYf;:62Q<(^:527\[UgO8.BB\8Y#.Edf9L_K[NR0>I_P4&@RNg#V
V>=-IZeZ8K3++0RAEg;XZH2PTL>KeYP[:/,7=5e)2X<1Z[==c]g-V77gWIY..9OO
G.@T6Fa@H<)LbKgIT&a4OA>;SPT9E#7LeP^.M;/S?:UMF[_@aJ#+gGVD2R]P]WG&
d4e1gHHQ7UCBXVTf&I#;\S8_GC-eR5<f4b/#7\FQcD)53]F_\9bRdAJV7VU0fKSX
(:M4/S+(^1WaA>ZdT-^d2I<T_FW8aSCN0=a\.N<G]R0=H7?XaJd2F,IX95/#(D#5
&EF,UW0(7QT5Y.WfB[a9BS@T=_I63de53Z1^fDRXLW(R8a1Q8R=@PVZG@?>H&\g1
GIMO&[dLU+ANOX/)4K,UVQX)3K:eW0T2WMJIBG<:Z3,6A/I&/?,\;M;)L-R3#CJJ
3B7f@^NM<bD8Cc(Ac@gUCc0G<7;GOO<.BK3SCDCS<?P70?(1YK5,<QEW](\B5]N4
F?Be@eFW36aRX=:LSY_0M401C1?@\YP53?VRTT<K2\LPN0E#U&QBWMDIH<M,cbW6
LB,CPL.KHR:a8T;+U,:ME;a1ZY67_0/63#=W:[6W<KOXZN)_dQN<MFa\F?96<caG
:f?&1Z-=a3\;eRa=6C:J)Jb6[/eW3#g3NW-(RKEf-6KV=>c)Z#36WNM<;7G<N+>U
b8&LOc+Q>)]KB5_#g0J?Ma\5:DL)>e)L>W--54C^LCA#;(f0^LI,4f_H.79FRbce
+2Ue8-]E<E@EK=?cO&X3?O>OR&:B.:_/:K)dQ[g(6YOdGMDK5g&7]S>3#g5:FVX]
-Q/<W2d(B,LLIL&+cWET>]D:4Y1T:M<f.PfD9a_]N:+@d,gJD-LTL4]F<:186YV/
&+7Z#>^g8ZJfOa@?ABb5KK)NMOPWW=LQ54]5R5AF;=I#,-Q\[(J^J<[@T)R;K<_Z
0&K6Hd>BCYb,4;fe)+_Gf:e_^XNB^#Feba]H/,W@_<J5G?9S)A\^P1EF8ef.b,K(
[)-59]LXX,cGd[:d0A]I)7>KXM/R8cER-YM,YWe0YN=YYR;,_<MXH:IH/Vd3<[IH
Ud@W6IZ4fXJONWU\NP6dW/e<1>F#:,IKQ4ZO=5Ig3ZPa4<K/3a+(J4SC=G_4e/F<
W()IB>E<T\A:QXNK12>RD;Y2<&aJe^>OG.OBYL.JAU=ZMHd5R@2#^AYZ#<KPIN(J
_Y1)&6XUC,fBDU#^)eF1LU#>LP3)ELb&_K-//N>86[_V,eC3d6RX@Z_]KK^.13=R
N)cDK/VEGA,.HWO?=7-I@B[_bWM7Df;7:X:.FF^?).W)0e/#cH[cE0g)2Y;.KD[0
?UbI[^>[3FU)5WOd-&)e@[2^XHUf8IRNSD]>ZWOR9S87^&N51I?QOP&Q#-f[G:Y&
W-?AJ;69ID_]=)cFV?J;eMcQXDMO^.N5WAQGM^cdPEVDIL6a;D1QWcPB:P/]92[:
,Y7@L;@]Qf0)\>.C&aOL-H]N(IM#</@61Vg_JD&S_b9PR(34W_]X61YU&1L,2fPN
W+d(5E7\QMNY=^Ja5g5/4IS<>E,R5(c/N^Aa@\491BDOCJd7)J)R4K>(O,3VG)OU
H^0\&:>4VM9IggP5-b@RNFMEA\deF@@;?Bg+)E##9JWUD8SO?d#<e/EI(d(Q30&R
9DV;>W#.\=::)c^CZ[A5]MYJgJU;E5A#Yd6H0W:gc^+FZgTJcUd2M?W6:UG13aBG
1AG:8b-/#[O4e]1H:d?.L2Fc(3)9:J8]MW&AXFRG[JB2:R]H:PSc&T?X&aPO3L-^
4BMg-N?Fd0JN-KX#F@5Z&V19JV4E^&<)5/+XRAa-U0;OZ=a+BI-#aCP,1,O)CgNF
ba#Ec(aAd9;A\]XY<6fTc6[?:R2d:CA>A)Ca\4PJ&]>VQ0.?f3cV[\S<C;5O;0@G
e+a\cD&;^P?9HRL4Pf6[3747Ag:<0+GO0AMQS\^K)<CG;eMF^a)46OBScNB09XWD
4LTc^;(/#5K)62<eKG>8gbbQA5(UTO_RRZR>,0g\Y9)A:c8f2-?N842e?Tf8?VOL
D01B^>D40WeUDLK\8(b3.HIdM3SJ>IRP>4fCfT7.X8Mc3PTICGeE\H6)1d3@C.#K
e.D^F3P)E+/?:_L@6TNDV2O-_-e4#;/65-A^VS1d>DELDU&.TO8M:8O^/PZAQZKb
2@BRP8c>\./>4M\<g.B^X1.E]+OXGLJYZ+G2@>=/McecY0;e>6RX6ecKc<HLRBQ6
KSW,;>P3JT6M3\\J\=e^-Z0F.B[9@Qa2\1LX<ND(Ca;RS-??BbJ9<:Tea2H:7&UH
dGeZa#2):-((X<[XaG0I:E7B8O8[RK?BD<J8312=fe/e[TY<]Lf_3#BEZF00^gU-
H:[C0?cI(QX<^O4<8eS+RG]A:2<QE@EX9^EebEW5.W-@T7CL-21DK.Ng;).c/Y]^
cK8MQ>O?2>K;:QZGUe9/LNQIHB)N0;c5(O3SLd];;J(T(GRR\=T\##Pgae^)MW0g
\g)D\BaPPH4(K(YK6D6R9VXVFU0Ya/bP]S3,552LW+\[T;UI&ZL&RG/dcH^E#6QG
I3QZIdM/)^ZX36HR&.2PZ4[G2.U@_XD]Oc54J-\&RM&2Y.@aB]X6W=T4GV/\-L/\
/EUT4J872B=-ULG:;_aP;USDeeZZENAXa)5gQ8E&NQTbXC71VbX^FVE]LZgO:TLN
IJBC1I8ZBN,/\e\HP.8a#.00/7#&3G^=&A21@Q>+6;;OP8b]IgJ0c7&J)A\7Q2BI
P:LP2e1YZM394#E_=M]CO?6[7V#JL#;V;bH^g[&[N_f8\TN)^@&S6;\>F]N-J=2I
E^>eF,88Q/59=20_FaBJ)gI&[(<P</.T4=--\,#;C-J1;Y>CRd2(O[+PJIIPAII6
[UQE/0[@/R6Dcg[]gScaW1g1VS&-Y\_C/9Y^#N<<6&T/PU\</#+BV.0L#,:SYY-.
:&]e[g0Z.WW&fX^PL;dQ^KF\4Ba,]0#SbW]fKaE1[KL:Pe5+fCMQ)?J\0a<0\YX=
+WJ48)_Lc[0J:=5K)Zf-6G8ZZ:I0YDAJQP4[;JW(Q1T95WR_R/;<[(IB^/^(K7[1
\ZM4?GW]^Gg2-Q=XS@D)b30D7,VZP_Feg]a(<8J1;E2Q7D[S8\B,gNLG(3[5Re+3
IO@BgXX)fYSZ.)gWMZI]52#N1Xc3J#R&A@B;A^?.GM/WT;4W&_PPU1VYT)K2OBX8
9[(2TdL/bPf-:JVMLB)baL\=^U)Ya>PAI7X^=aVW)E0CX,Q6eb>DLI2E1>N9A+)g
-Z84>1-.XJFQFI2LL\86S678a+aP>M>aTVX#<7B9fJ5HaUL).HfX7K5-<B9F,LNQ
7)UdW-^[CLS[.I:K=V6W^5IYM@a_d&I6N+E+,/g?;EUQ2&0OI0L>&6T8BS:WP]C=
M_LT6]4E(W--@_WU:;dDf:HaR+Dg<Z[g,3.JUe_5H.c>P2<J9]T:6TYSBVQQaFa>
]K?JaVII.6XOK>PN>=f)-bQURV5VF@H8:]4CN311FG2I0aS4QAN1I=G[K>EODEZB
J/:VWPRW^e@f#D=fE[D2Vg9+&RJ;EV+EJ9gL;,BW0Ac==_4=T\M>D4HF-Jg6G(3-
/L,_Sd55G?0G)b&g<5Z@_9SI0.R9M5(@YO6X9-\K\VeN2V+J&@CC]Pd,agU1U&)W
dKXJ#NH2_^S]?>BRI0U]3a\?,<Y4#<UYCH_H0/Z0HXK[G7&J.)G7&,<=cd,E:;4A
dZ(&\N;YI_NTEe^V4X5097c\R)^5-?Y45WN=11ePI]-5M_7@75E?7ZHPGPSN#EZR
f])f;V,WK83TDgERb4?2b,L;)YF44=@Ye?\G-8@GR(2TLKC^XcJOV,\O93O]]TOc
QC=97b;-][[)OGR.[e(L-=<<W@;_7M#WD3\D5DRKd,&:R#)O>SCS07SG@1A4;Fa#
I\Mc74P(;XPA.Y-[F2B-2Y;B849O,5:#W,UKT_V>b3/faIOC4O&S/I^Y(/J?-DKX
_J@EEBJN;AdB^#[XP\e#:#>72U[bY@8NabLg0X9U]Ga[ZaSRWC>DRO?G//\0ZGN1
BIM2[TV,P7MGf023dKE08U3MEH&E[Y.IXA4D[5I??]\O]C5-1\(IO,/Sg2Q[c])S
UFL\4A9WL8>@H8U>ZN0,bf/QQ,00-VWCRTF#T6]3V>M.,LE.1^L=/-+0H275S[]=
bUY)acX-,bXJ.TPP+M:<aLR^OgL472[^IJ<TXUd/^UX]T5S4S,>5N^fD[;=I^N67
CIE7?6(-CX/3N;0cPRDTNZQE7+T];TX,Y]:5.58^<ZQNJ\&a5>:Ib\L9Q[F/bOOW
0R9#d8de^bMG+,H7;)SE\6HWHTd3J#bP35+A>7(>DRRWJ^IDUK7UGOZAb:MQ/U)J
NYNR?[815^T;PJ7L\0)g0.EW2V-;5]Y^IPV9:SbKe)e=I-U1SC:RfPWG._WFI#-C
FD6gb-1Xd_3,WS5:^;f/I=9-:V^&CgV2/KfYSO&bA)<7,J4M4-&VV]5^[[(_J(#(
O.]<X_b7IOFS)Q3c-dO6JP]6..#PLE6,BL5HR@_).F3+=)c<a9.gaZ[[9&MP<D9J
)I]&CE>OF]f?SgHVOBQJ=R;a)He,c])>812)BWDH&--<E_YY<IC-D^e9RZ<34#Ea
>YC_<52-d9,(IL]J)K?2[3V;_7N83N1WF^Z5F/<A\bB1\L?cD;.d>T&@A,:)2)L_
AX7-TLK\:R\5NEgc-dHW<)dcH(RWVIWa4/aJ<Yc8?=X;Wg&b;TOa-#W5?)YTf,c)
W_c26ZCV=OZ8JZfgIJ_@GBeYZ>,@<)W=<Y9+A9aZ0JH+T.6]]4BOdS7[@M+@PQ]F
Q\f(^3PM7+=-YKaa\_0fFB0V=]H((RQ/_R5^8W3>eCeOU+LU^MXMFZ<)YaG?M)+Y
3\4I?J6R\SRY,C3I1e.-Y]aa]c6Z[_,A.\^W?FX_-+\,?#)724K>+G02TBA1J++=
&Wd@PRQ@3Ee]NUY@H,X4Ca)+ZX[0\5,P+5.W0K:O<Bb9:H:g+PB,IIR_<0P7cNCQ
)O?D>:2MB>(-E0<.GY=47LMH5QJ48#^eG+K]AG[6=+E/,6eV5:S<X:8K;LdC@=;5
Z6.)[1J7P]/K\4]aI=eVECUBcb]d6ZM]<;GKB,f<[MT)NG/GYU82/I-fZE:1SWaO
>5W7YMQ\D],N7#\>eX/AH@9A(#76UM1EL3\64A4R5I1,L7+I/YW5GSWQ/G3SCLa)
JM/L=C[H]_JIFZe[cA\0H@>cW=JU=,RAf[J-7R5AaCUBYPc9OKL/A+YTX9)^PD55
[5210[cKf4XIG+=Y3))E#U&9bFf6-:G6aVL^UN.^PC/HgTgdO9XbG:4LcU??)f-X
#4a)>V:5QeZS08A2RU<#ZM2@ba5H1aB/V:PSN.RL(cHd\6;bB3QQOI]UNC^7g++2
[KFc2.^I?eTZDPSc6)&P0/?<H#,dM6\bT)&)MM:LHSMMA1._Ed,9^>T,SgU9M&MP
JJ;U8.XAB-a6PYG5P2+LIRM/J2;:E)>JV4eV8K(53]Eg\[YL+WU(ba;)0R/Q-]cM
K@e7/\LSJ1?#CUC7K?PIU^fRVe<aYQV1IMd=GTI6^KAVO2/HP8#9WDNBDI8QBYCO
Y\PEX),E,/D7+U_JP#G2VT)0&+_(1Ne;.RXW,Z[gM<-f:[J?7-5d0JRMTXK)7c>U
5,9N+DR-@C_eSZ9Kf5/FD@PMCE9D&e6Z7_H@?WM<8K/7-OYF4\dfZB?DGTG(7&GQ
^4T/]5a6+P6?>C0IMK1EeaAP=0&JEH=)M24,e6eZ+H9&<cG4#UCA7cV-N2A(Zb,-
.G.E-0L,Xa#I1bSIXPV(1OH1QJG1EEP#=#);H=ATQ-[@L[,JTZ4Z&7IL=3@&K^W0
G\VaQW/Hc<HP#+7V[(097faS:c)9?M\_I8fKYN]X7d<G,^:\)f\ZRVIgb\KWT.KK
YZTb7=-)NQ#.D+Q3L?/dDIW7FN>1/&]4M3_Pa7a9L+3U:/2@DWQ,E,V4.I#Ta1TO
2630B6fD4#0.)@@T@..eI;KTLf8d-7O<0CNa#]P.UO/UN#WT6FF[4WQL1aGOU?Bd
SS.FaBQJG1fQ1cE@GTad@Ld/+AA,^,fGN^+5JK0ffV.2(DNXb/,:21E&@?G/+&\H
[W#g:.70&&F+gE=EL8gC4XB6UfH/R=WFZUX[a[KEKb_a/2GX;]\RNEY0=X7BBS6G
[LA3A#>7PVb_SG0]_YN_?@5AH)c2VD#Wd#QO9+;,P[(VfX1bQB9@fAQ[Z0^;4^T.
:,b]:7@TTf-2Q_8A77#2g.e_G&cJ;IdSC)d/.@(Y.4AOG=FF1J?GDG4#aY+9O#/0
FeDY\;.\G)X3NL2eFB1>Z?72@_=a6\ZO-[,c5?Ve\cgQ<?6XaeP.+caALEZOAKM<
3(PD4?e[Cd>@C[_=N?TKFD#3b;Ka_5W[e,6LeS::[TR3]Oc<+\=+fO]XIWa,0J^>
Q9f5fe<ebJW?dMEMIR,Ab>3YHG;_bC?XgD0;J\^LQR(U;abB_HgS.<XdZ.MY7d>3
4(R+.XJP)f5>)51[^>[Q1UeS#I;7ZbN0Nc9Y:Re_4M8V_K4#ABNc.Q]5DK=8DW0I
Yfe4?dL,MB)+ODYFeaEd_T>#T\e#[<JY+MCbd+^PB<^4RAccOHZ#gY\7=Q4QAK->
42MJ_:IX]c8Y#P_#=e8AZ2H=L[C[FM\F?OgU0aV4NO&F80ZH0D6186U-KKYV9[1D
?Qg)WT(@F7&gJ6g9cMDGc\O:A3:6YcaPWT\][\K46:Rb@_-c8//0DKN[=#-4BE:_
g@&/_;?c9?YBYG2La-T4HPN.G[&XT=E?I3+?QF,/LbeN;LcOR??Nb5JD9WU=8<W^
?E7H0AU)U;g@(_B#C:]g)eTaK>aOFaO\FO^E@3T;B74bI/TBcCB<?gcRL]FI_JR<
PDW=3T/B8a7O+,L9FNL1dJDgN7dM^(3,0WGU+2/49:>39Z.N_EA(f7VCbI+D&D<.
<bb4VXMe^E[)5VIO_c)8=.>GaCKA,J&2DEf#1X?PHgc>JdN-=@G(_edbS40(]YNW
;1[V-R5BRTH,0@E9B:&ID@#PH.K-[^f-(b>.&12Q\T,e2bFR@^R)V,?A7WgCU@Xg
IZNeI;R?M:N;S<K/T.\gG>OgPY0/XUG46PM08>IdC7WCGIg43]b88XD[8Q1C0J>d
JX4^5B8D3R[_c2d1B,E3S4N>G(J8#)R#7>dK?c2G2]K+MH6e\,55(L3fV)B:07]X
TR\)PgK-]A(5=JOBF_dVE;>LD1B,U=R?_[GFXP<ae&9NeAJ_R;JQ9J7^04LTOV(Z
G[9EDE3W3bPY].OGR[#0G5MH?PLaWJWdc?W9:_92.#QXM_CT2MCV)=_>?\W62K&&
=4BM9WPMDaJg\N8eL00^8,fR;4a^[#6->/TfQO\]A8I0FVYAZFORKHV[0S@)#gS.
[^:;/6Ee&2A_0;ge<#c8GXY:2X\<>Nd=(98CDKCQeHYCU-0(cd25SEFU\LPDL6e(
_[fYg)1P^X;(TdEHW2f.g@NdE@fME]6,VfYNM<a61DP)MG<>8H+XCBfI]d]/LR^N
O[O5U#Q>OW^F0a_04:FBU?b:d?;8HT[#N?[)Y<3MV1R=X-<8HP#gT])L-/eYGX4H
PA?.8b(@TNYTZN#_Y^2J)<bR5C\<14R>Zc+V6&5U&^(E3&:1)&P@+EDRcZc@_3Ag
6d8IVDQGJKZ#MMb8fA91&H5TUQOg;fb&bbK4E[&;BWV&,&dC-6E1A_S<fRM-cN@>
5,==;D(YU&3N)]g<A<;)>Y;2E;R;=c>:5Q=4gaF-\e.7R_#S(YD:LSPC+NaTTZUE
ffW/\<9Y+D<5<;<^TCg.JW5aYVTLO=HG/:7>R/K>R&c5Ha>aGKLc^;I<@?+UAE6c
/3X.\STGA4W1C,(U>_8d\9/HIW]+SZDV1UR:g3B[DE=e5.B_.JEPI@A#S6A<+RG>
&,;2.,D1TM0?@R<<Ac42TBcLe0]8@/XI48d9DPC@BTf<J=H+\6&5[/,?[?.M5ENM
SLaG679?BLZaYc-O]TZ=d[cK&d\M<ON(1ZSFU]ILO2HXEKZ7EWL-K9_Y91g.&,fG
P3^C27[[6L+:J64\I-^0,+C[?6R@?M0)&@(cf2f<BCc9=65=[\BGA9ab[9cL\e+Q
LRM^9T4^6g.JcA3>1DOV0^#cAg(R^f(GU3+>00eQSI1fQ-_5U@V80g^H,1P,O4(g
ae_WX,DPFQUN\AA;ZXdN&AIaICDM05_+=ZFT-](5H.(=5J@Z,^+IIJ7Z:]UH+LMA
>F_0AZUW>KKVG]P\IK(^E,YBU)8d2\MGb;U&g-M[::]+FfQONQ&58_K6ONe02JRc
e<5gf+aM:\OJ28TZEEF\RJ=e#X\@IF6MaR81(]/6@10P7&MKI7(.&b97EH<He1[:
9BK#=b1DFd69VYbC0STA.WDQV.-\Fd4.G[38GC3M4-904b(N?Fg=-(YS7\cVXMK4
EFA@?_fD:6:;VQNWD-4L6(KB<g[^b@He/Qe4U#S]H^;IQT9U7GNTKO<66[3a/.LR
(NT53.IO5-TcRUa&/R5BYb>B4R7g9NXVT\26H/S^..TEbE=Yba=,&X2SXPC74FC)
?6&<]A>E]Z4ECT(#2O7X?-K2SWVCM40FE@O<N^\MR:&Nc\&0(G9-DXR.@C,9_+SY
UY:BG2IbJ(<<e8Od\J]<d.f?Ya14W^7bXX??A3dBH-fO\LDFPS7B2fOK8<&3RK11
&2CXKQLSg4<a7I(bg2g;DAQ7+e8:3cBDIHI\;:A=YMF#25/RgH@,35:0(JA+_798
FB0]S=-W<Z,]4EJE2e1EZ0&2Ia8c0S&e+23XUG0\5Y?0/-4\+K8P\aIS+F7D_0,I
^WJOO-3a0Hd([=W;a3XYUN^=CF&X42F6/8:=YZCgFO0/<;&1/PF)RUASg3Y&-VV4
D[dN.15E;KVGV[7-IL:6AM)[0_/PQ/=>[N^_Rg=-#TWO,WYE0MTdZVIDPC&;21[2
=FC_LVQJ-G^Ha)UVgTa)JXB9?cC,YH\I:>^THD94M6S]#.)/?C6+E@U.)Y\7a\>8
R?;I7P@aQCUX\Y+c3I]39a&0Z6SK7?A22bP2;GET]8:2dQ\Ea:=&0[#&7;H(5Z:S
RbD^^dMHD2N>P&-3e.Z)7P/MLCHG1SLN+KTaBF2HG-W9JJeMM16/1)JL))JdW-ac
^K7^3KEdb[L<AQgTc=Ue.:]g\AGVPG6@59M3_B@6ZG@I3PF&;@QaS<XgWK0&AA.O
DV0A8S/ffOH]Z&2gcb(,@3)CRcM94^a0JRZT(L1^c[<Z004QB?5WV[295f7(ZF5c
/G69;,&5g]Q6f3IG^[HYH,233L).Qb;bUcED;/-65<f8@O[g>c77#>LXcf\SF:cF
.-ZAf^@KHV;^cf21NV/L<AVRDg[8@>M=4FZ<,Q-J&6C#5V-)(WcO4]>#Q^8V6H.a
)+_gGE8e4_Y.N+I=<H0<eJ\ORc^XFCR1=A2?)UB)ff^Q_\Z/SMP]JZ9(CUA;BQGY
-U)Y]8^K0MDF5G_QN46B<BDbPeN41E#I]c]0LW@>UAK#E0JQ4aOAbe<X1bIHaE;S
CcY\NN:J=&&T?:f)<A+2E7X_TNfMbSQ?P6TB3M)YC-P?69S(=0^J[>17T4KE5NAA
_Bg9HQ;K.CZH@0Yd5IFOVT3G_;U)Be@@:QH)Q3X6)U,G9X2Q88,@SCDW-_.]B?2\
aLE40_,?PL:^A(=JTU&X+HAOVB]+b=_:dA):?:S0S<0(,W[^8b4,0^1af+H.g_eC
X;=;aXX95:VL^+?WUc0W:aDH;NZ_A@1.b9CKEbbBJ=TRMWCD]HRA[QU6Df^+&L4T
d.aG2Ng,YWEL;d?WQSbRN6FFe@L8)(2W=+:@F+G3=4Wa&dVNOL-cE]O6G,a=KQW7
_5FP236,Wg\]+;RFD.8/PAb[J5V.X&B>XF/,O2PBU](F5G]\FYNN4c>U,8fU4;T7
g5N-gbEfPfF5[3_A@M<d^H/62)JDLI:^TDG^58:)>&GWJHD_Q+M@_.6UPR(UTMBa
,V)Ib09D;T6dML:\&0ae0C0U;#A&_,R.+cYJ0K-B7B_J@-cVf4Bbd9;.,5;:b]g<
a\+SeGAX2QDSL>/W&?:_cb>TD5JeJR#\B)ZMYQ&SD:dBY=:E@:ZR>Z1de>MbfO?[
U#.EPVJ_DIP,PD1<R7W@)U3a(73<?E2MD;d+T\RGPSMb+,VJZ4_02XQgF:+)>e,O
LLC@c:][#_^?X\5Wb3(N/@]-FDMU0>7&T2EZE<gC39:c+2ad\bTH&_[WeUEU9<?^
W,8:RP1R(C]>6I_OOg9>U6,W4H&dLE&ER5J7YI(+O6<_e]d5ASV^+H2#FbW@KNO:
)OA<Ba9,(RJE8)<K,V@6fcgY8E0R&e=QE?DAedJ&c>KFT=G.WNbUWg7=.QCMD?D6
MF<X@H)aCe(D;R=27[JaReO9:eaJgVeK+L.HLJ]96bB:S2OgTDQ#/<&Y-=KVC:Cg
6CR)D21O(#g1f@0R6XJ<5aN8\57]@;(#/@4DD]5b]@U,07^^-A5=E]]F@Ba:e+2C
Z2c3bfLVBB84#-De57V38bgcV)KTH0Dce<R^+C(TM/#)JebE2,&f]J0ZB^G/9F&c
SLH4[+B@g6(Nd,G=A2O&:64QMe8A6_JIc_FM=;/BSV[2.#PZ5\#6;DgL:L?>)#(4
T<HB6IJW9<=O74C+S#23TSVQ<W-?Y&1e3dGU7DOILOfM(_^^^cOCTO#B<=Dg@]c)
,S18ANb8@J0[4L2]H>@.#D;]^^&=Yd]6LJg3JF_DN]>58_HM<UPX<+.fFOB2GB81
290W.@_Q_05Le[V]g\1-&1J2SAZD<X=ZM=#<_>9QW>L:,P/&&f_e3ZdIQR4Ab;<J
+,FYB?5cEZg>IK;E@6dW25DMMVR.FS8fdd]+d-75ebM.cH)20_3A[[>GE-H\VW7N
KJIU1AFb8M>P1W7B^X]00cT5Q:=V52-UeDN,fTXSO.R<:H9We#MY0ZZ))2Re1=8B
#Z<5G=>/-M97R.=cL]PGLA\@<S5JLNE0\RXHS9EL[#-9RS_46C#8,NDE68ET_Ge#
>-6YD+_d[fe-<0f):F&N]PD1O(5I-VO=0a21P+?T7Nf<#MV.H?LVd3ZPO9,QJ8BI
dFQLEH>W\4/&S]ZA-<Fe(_U89SWZI>LW@QZ-S-(U7X]^5+&Ug+VIfDb<V.M9<3#A
3LX>ebg[?/C&N[6;^N3?5:gc_ecdfP++7fbY?#Yc,)A+aC<>Yg0YUZ-\+bGf6cK:
SKcE50Z2M:5I)d&@>YW(STI<&=@/DSF)TP+./:X#PI,?a.I.YT5<7fUG\@NZOe.M
?;/WgWF)aU=)FbS3-J]DK8d=@0Zg^+UVM;Z-NcH>6c.FTFENg(2=U/(TF^9[+M7(
V;8I13X?L[.1g2cZZOO<?GN9?&]]E(QSbDG)2/@=R,g:9:)DLD7P\J.I?4<MS4dN
5JR/c39Z7a^[ZXHf.RW&,M;b.\R[:A.OA#T::WP1Q0PG?G=3I5Y9&cDWGR#E=U].
<:OES\.:+-\f9_&YN@5\U]ETd=Cd,LF.VAHV0;8VP@QV@LL6SPZ6.eS:&94PRAQK
;8=BG/@V\UN.T2<>)=-+2BF_DO.[Tg+M:EB1446BN&8]cBaT.g+YU9^K-;WT)?(.
9gUb?>FT25COTUaQ,?e;V,V=Y1?##e8)_QAZ1d4C<ac#a64dK441g^12W>\K8B^H
H[M-Y@F]2@(10+V9DXC6QP1Ag\-/>M513L=:)D)@V>Jg&WMUbGMabAJZ7&^+G59[
ODSJ:OE7VU-\H\b>CASP;FT1cJTK-)MMH?gT:\?P,THS9Bf5>+_d.K_4eE/]gDW?
7bF/@)=d^=QM9NRNPBH-51-.48+aeHG6:,eg&TKECL&CM6O0Z&30U5J-.6#2IEN)
AJf@,PF>)B1;f=H;=@0=J@QS_P4J,):Je:(8)_8+NZL[)NLF2OGdRZA[&FSU;@U&
\W57;?O2V:8N13#=gFg[I=?JAP<VON()1#eE4BU#AQe9=KBd&[DUA1I?QAFPSEJJ
FHP<D2D#4??ES4EM-0#IAN/<4A/JFK><W[J9e(?f@(gAcB41V&MbG-MV)D^[:cKB
I)<PL0>-1YFQ]f:=fd&06IOTfI3A^&1?FTC^6#0D-1B4+8G;@=[ZF[-11V3W;BWe
Hbe@-@1Z.+6/g&2RT,C9d+9TF3PE0XSU1=g4.d_^Y8\X@DNT9V9(W<(X38_OcTU,
_Re\.(>YT=6)S=D<:E5a(Ea;d?W>eT<Mf<F50C_UTVTgI3KTKCd6NAGCMQ_2AG(W
GfHN=<EL9gaMgdXfCL/XEAcOOAXM=f(c&Haf?@X:(5]&LY3F&Y+65WdHQR#CI4d?
H.<F5\:Kg8C[2dg48EC_)/=M2aZA/]<Wb29:Pd.D<9_26C\14dY3eN=?g6cd[\0@
.D)]Y.2D85Ze&B[AT8A_-59B-CFAZ3Z85aQO@9(G[=^3+CV7ETH/,29Ib=6Y4O(c
70G?<d]ebUW@J[GPVQMYc5GKe@/6,>C)&R<2N4#DE)g/H[B&RK-F:G6[F+R61)WV
?<b6#SR5)DL24R/,FFA,5bAN.QV]]g5_.C;b<5TK]d(13<0_0d_bURe;Ja8(bG;0
^E]G&Xcf-I),W0J0eC0[::]U&;MEWe5KU0G.=WN-FaS&+Hb3Q_9D4_G8;<-Kcd^J
U]5d[#g1_9=RZ/D71,3H5aBH2@:b3>:B)=U@PggPdNWg6P)LV#cQA==cY8=](f#A
deI[HB19?;GL\[1c:?6=1^P?#-#B8:W1Ia3WBg,Nc]a]TU&+>ON@W7_0[UWL??]N
AH[2K-::fODP8bA/NNAaCQL:_C=[a#;?>V#:DY\V<,c5HRb9a;(M8TQG,dYf+LY<
GLM_5,3+=,5^M8gd9XdYU)<e;FdGAZc<;05(GV9X@PC4OGJ/K8?EAI.+FUV=DXJG
?S;4YR=0B4ZdFB/51<\0[XbG/T[gUTbBMfQ1^)Ha86A-</X-ZX6968G6CS)/NANR
9)/P,bY_cN793>7EDd,VS?7a.&,<.1D0.12dgXISKaOX=d8c:,W=[1X>(fgJESQ6
(Ya_A1E4A7:Ed9<+eR8Z)V&KTN#R5NBeJ)7\T_22NY^2F:Qc?)O6<PL.#WE\1K=(
=^T2;?8eM:_@CW=4[C.]MG#S=^-[,QgY#P1JX&\NAZ:7I>2TKcSUWOgEJ8Gea[5a
?aFDTV9X?:W<1+?Jg.0&)_,IJ),gXgDS9Y+[&#VAG)P4D&VY<\Pf2fVG5VE-YbFS
c8PUPQHAFTQ^FEYFMY<5HZS:D/8LNKfRJc8f_<\8R>^6@6Na[aKbRegMXNUWJ]8f
#)F:MV?0S.\>b.:JR^+G:V;&NUEb3ZIL9N-=9QWcZWg+^HHVPY8C5[/.e>C4H&99
L<G=8f<\b\3+2)PaV,W8FSJ>W@^XVYGIa_M(H(S4[O\IITV<c4TWP8F.d@cNNIJe
TX_:E.N@CYV107?S]Hd_PK<<=2_2;KVTFZ??^bc>>9N0679H0U4)U[.Q><EJE4b7
A:ULY.MWN5T8YYY1A;U7M0Oa9(&9e=SM+K/]414(M&^HJ8LbFJ^](La3XD1U=Y=@
^DN-IRBJ6GDb^1[Q#L+g=aM\HWcQ#SBg.P>>\>U&UVe.9/P7-YN/3KEGc9](([O+
ZEIQ_YYWaX2Nf_XFJ9THTRBaCIIT7KAMg.b0WB#6&e\H0Uf5CT^3FGN1WbZL(cRY
Z[R1c)b?>I_:,\CD#e?M0G/cC4@9K;0<\1#d&<08\IcVF5S5T^9,X1T#F>3-?+XO
9f_YRccZ#LQ)WcY@D87CDMHDZG#JE[7ee57K/c4\1MW-P0?f>TF]3G[DGFaaK&^e
dUV_,;da5ZDJ8-OfZ-O4#E20g0BR>@Y+;PY4bcF1^I9SaGb2I0S&S55TG)0IaPR^
O)LCJEa1TANL:CL5:d&)(XA1M(aY.EIL+/U<#=A6C>A/4S^fKSUL7YF6;cUOOZEP
T<=dDC_VN--bPYMP871,VYRa98dfERVdCc@&R1fSA=^6>@P@8V^KeD8[4@N^D[<c
B@PK=+[B0V)A68XTN?=U:+=H1F=9d5Q(V+f9cN6._<I&:HLK9)A2d_P>:<B4L7d(
2OM/O^dFF_59bE7UM+ZDHUZT:Lf?GcS2RffK5Y(-]KGgYQ?bIX^D7@HI4,I\Y<R,
A[A^3W#0OQDMHf[6NYc_W=ID>@4X2FaB<#S[G][1P]IbVZ_H38Cee[5eI-FfVW6>
)?WA7IdTN(QYH&Ya&4?<F=I3UE\C^MdG)Oa_TgCK3/[M4?U_B>d9N4M=/L8Nfa<=
&,54^2R6;0gA#))14\08##=E120[E.SD]YQ<YL3[2f/1QW?.^b/adP#-A-#gS9A,
dTB3E0DM]8N>YY;/g0<SFX5)0T]?N_X7M>-J\_,eJf5T-OA)#5&589V/Z7-JY-1Y
2J[:I^IC^&dB3_>X/GR#HRN-g]]+9PJ6X7N27,2.gSCcVOK;KD@HDbNU@aGL<+YD
:7dA=BHC&#K^JEcT6B):GA46,cB74eXG?99-]N+f3NRY4X8B0QEY6?^IfCVRG]T>
OYN/5=E.YFI]:g\69<>.8N7W;Q+][W/Le_4cPD3DO1H-<GP&Z=RKMON8)^QQ?CPU
.W=8<=B(_/IDd925[4.YCEJ&(>OR0@5Wc:^GZZEXYe)fNTL??3UYXM1IN)P+b8L;
MN&&<@EG]9O2UFf.caU:F4&29_XBMF6BbFFF7:R&J#EJ&]f6+\(WU2EAV/]Ja&ZR
-d:=3\37\E=6HUG7UdVB&_SA?(-8fR5b+T_g6/SWTgO7b-Q:+[0FRD4TMe#^I9I4
G+2S]<:+S:]I5,P\?2ULT067RGATb5eBbCQ6aEf19^K4650&_Z^\#08AELY28QX.
6<3AOc(VM7XW+4E=eSY7EDA5<AAXIIS1f.>Sg:B/.e0361bc,=DP?NO5?_>V6RX9
:P](,A_P1SU]eI-MHfa[<Y6I3b>,d6<10+=gRHc:K6-EH6JbEJF,?.bHLNBOU(&1
/,^@J5YE5.TK4YIMSc7KPKU^@&BW,OA^<ECZVBWf&63^,NJ:@WJA5BG7F9Db#;ZT
Rf(;A+#69\ZJK+8BQ\RNF-XG3d5/X9)CW(DCN-:M6ZYG@ISUKU]+g:4eO:d8FP<-
?5-&\X#/^(NGg=Ue50.JB3()-K<)_^cP0D&JY&WF9,KG^SG8Ndg3]&\(<S=ZDXQC
KOUMH3#[Fc]?]]9K2Q/0?)Y02O[QLb</)EPgKb]f<M_G#,LHK8A:9SUD8TYFY)H>
[L7NF;#B:dL73+P3Gd?<J]WC3E<Q5A\[=]A-=-180QL5CB]ZR74ecJH.0O1E\=B5
e9PVPb=Dc&Dc)-(_,_d&@OIIQT9T&?Rc&:E>0C.#D?PeJbPH]S//,Z<b71eXO90J
GB0OX_I9S=SA9>AcPeU4,0BdAV^K<CTN:V4f2PRL_6IFQQC,WIF#R\8K#GNLCf3C
(_B<WAG\JMa#=DG+ILDWCWf9P\7@UCJNW2U2=Z>GX[4<0NAZfW,K[D,7SJ+.3L2I
W4F570#G^K6ZM:_c_&]gO@^0,B+8&1V8>1(PEdK3DO\VB?bMF>5HY\E9(S:@(QCQ
]G=AT3Q_P&CB/7+0-L3(4CB_=V]MM\2gC\2^aN@KD7B;G@A3FNO4B,0@F?VTJ\44
DK3@:7eeM<GCW5IbS.+./LRH#NM7=g(c)5>Q?__GPJWD@)e^Ad+&5574RD&WU2b>
.)1((b^g4IH3ce2B_9=<#bM,3Md&#bW&;EFf3X2;0E.339+[aTC^;ZbGWSVT^#DD
aBEc?HZ)PZXVNR_f=Z8#X4^LU>/E>NQMGHE^g#<2U68,900XGMg4=4JN1fbK/-Y,
^0b_>JIKT_]B-\e\2b)C^&_g^W3a#)FQ0?Y<a#O9P>+:M3G[EFL9ALc7#_b^6@8G
VAQ6G#\Y7C?KZ/>/VF1X/8E&I@>]_NP^5Idc\J]10GDPLa.(4d=TT\6HY(PE;5;D
PS6+L_QaVN#^+dH+RNF)^<#1R1BB,>?eLca-f_E_aK:Jf7,f,0&1V5@ES\M/dS0L
>;afdH@3^=E^S3T++G:F@5I-Z<J7/KQ5e0#ccL99D9Z-XW4.[@=4;D712:JFU56I
ac.4\a(96_#RTcR-T954\@27V)4(PaT7f.6LI>L[7[3TS_<[T__[=M:4G:?+7A@O
PfG,fQSN)?A^#-S+.=_]T]CGS?2\U(3Q0</)_XKZ]FfT^&-5B^&-P0@(3TPDJVR-
UWAP+4TUFV@A^-Y1F4)QAc:WR(=N9HC[1)d9.GK645?QDJP&NDQD35D>X@W\fAK-
PD(TOK)eA3(+>gK1D-OKJKB>V8OG+,;a9JdPNR,]7U;?#H=W])@,R9FV.LEAQ\Z^
+/b#X>Y.QE1BU4A>NCRDWB;;[74g=aKc4#>XX0#(&P,eM;J=L)d-B<Q@X6\:Ugb4
B2L0\Fc2J:#5,Uce&\Z1WJ^e0Df;CQb(fXF16[_]1<W6#5\?eO]>:M7RLKgeP_-,
<2HZ0F8FU+17Q,GZN\35_2Ab.V95@XXD5A@9QF<gR2=221(/?=,He/(Ad[VOUYI-
P@T=A6K@EJXHFaG#[E^-H/P[_D[EaAWS#aYZ=N7V[@)b?(2\B^G\:\\XaBZ#5^cR
1CdbJ&(A@HM@7W>(KR^gI_^BZ?:67U[-Hc,Z39(184,XB_25=[,&IZ&B2=_0UD)J
];4A<_^&OP?TO)DQdDGXWe?EJaY6-(MS1IRB\?FP]YLTM_3c=Fac3)F#I-=BA#a;
]DG[MRgV7_G)d)W>18IHWS\ZU[3LeK#VgaAaU/Lg4DNd#+2fVEb&2\^O(bKS)(#_
]Q^K3c^UQfO#HJfVe<5R2KQX]DB=-;V1UOeEgg.+[=86V.AO[BMYC&ZQI+NTX0Ta
B@@AK2TOF#[/;30@RVZ<6&Ub5C?QgYGbW\Ka9#+JBg3-CB1MgD(@A1bOO&=86V\X
@d-]DU3dEDGI.N4&>DRKdS5_9YG?f8&FXGN[@S#Ba3Z,@FWI:HSTSY2N6&JNK)D;
V_)9dAMdaW?V#5e+U[5b.2g];,21dP<43F]^OGDF?HfBJ(^:+,O:<YD[/b=E0R6d
9[cVF6&I\LRcEa)X5cH?^:D:7g6A)-F9_G@=@UZ\[=0c-+453Ka@eZf7Q-E@FDCK
G8e11VWOS\Z&5MH32[EF+8&Ab]Le6Y]7@2KZ6#U(>bb6[+[b+.-;K_Ke_D-D?[BU
:35MI73).g31P<U<OUcY0.b4X:4+=Y0JR9,,T1RbL4bD_MA<@>\eQD)b4.L/&gc-
HK/6FX.37[5[@0V8<0<D7_^:<A_9,G1)1b/5f9RcJAKbe&>)+4_aBE)&G(N03YW;
3d\SNPX^#5fB5>RJaC3\W9S^+JUPd6Q&7g__T>O.>eRA_X2?MG_MH/[&7WFJWV7\
;c#;^42/W8L/9cZ]F>>N@b(2Ig;<6_X]EN43,@-b9J)J6^Fe@;,I&ZEG?;0-&bO(
B#0#<_4]>TH<8I\[X3D=P,62]G1d\9J/d[NZ&&\C5>OSF]#BK6]_AY+W@>=NZcdZ
aKR.If^Ncf&-MB=7fg_@d[JNI\,H5^7N<bGPX_]@Bd_1V5??gTPHUNd<C@^<]<GE
4KOZRF^QASKR=R_<_fH/Q5HHDO5.0N(7=<USEU:5f0N25VA3dVZ&9M5eJc?V]S#g
QI)4:0;)7[#FUT-a/f(&2__b<^]e]BX(8.E75F_dcO8;YaXR)/A?P0a#7g8?GV3[
HBS#<RDGE?R@\5Qd9UIE]gIBM.ZDZ\^\C3f73>\;@cKFG33:O+feDFX=I5YS3OP(
=R-B)B_K_YgC3R:MTKDJ1L9a_EQeA5e4Cb9cU#8Q0YF:bX]efQ&L1KHSaU5W,2DA
O38K=\JQA?.ed,#_:@A]^W6TMFH6g+-80X65X>aeDY3A7IIMT90XZT?RU4MM>IS]
TMI_^>LV^aBcGJ=.cY73Kf\f2ZI@5/X-G85\RgQJ8]a9)=e1N+A<6)CM];@IYS.O
e:^J_@Dg#b8Q(c/JLJSGGE,aCQG4Xf-#H(A((.gRDJJ7VLS>S6gDW?^?Gf<MN6Fc
<\STDIA,I]>25B8YZ@3?e?)GQ4.KW[7L?:>gXP6bCbM,=&c=V?IP;#VFP[/1^GFT
Z]@bR(;HTDFQfC/35YO9P#RCT/^@>eR3E6L5W=9)=<7ff_;2F#JNB&EdNIV.e9.d
MaS?ZT_EAe_71\)KX>(<#SCU2b16CA#eQ+BPXK=O5GP0a7F2OEfNQfNR[O),N>:d
KHU>WA0SUc(4WNIKCe-a_C8E7,Ob;U,C[3R<4AH-8e/f=5d7WZ;[5G:K85Q;]<9M
A@J/34,B9abD/)\&9cYJ:=Z1?Tf<TRT1>1aKJ=O,KfT]-C;4(V&\f,07IQPW#ZIM
&\dQA;[5F+8Sb=PBN7=HPJ&2\7LYKINI&FD=2QVT)aU>URb(FV5J^:@]K51CS+)5
)9W^\3>T)_B,S:Y^^?,U;MJC4D6;Vb68a=dM6,d83/F2g;b9AgV7I1KZMQP8KQ23
#fX=Z5S@(OW(1S?=)\Q&974-O(;CcVBYDDOYUM5TVQLgN+N^U,cS03:.NK7D?^X:
#fR_=57/-<AE5=0]A&,9T[7Na,8YXZBR\,QJ]d8A^1DbF;09f1ROC5>K)@fPf&V+
W/LfCR/=SYbM<EP#.1C2_U(g9Ud^7d-dU^H7W1X;X,ZgV^.+WQ:F/Ye3Zbd4cg(C
AI910G9;8@WZ52bP;I(P([7PN_7@1(;ONY]WR0)gEbd@;?#3ZdN[C9e3MR1[-:b?
@S/C_(=3e7a6d)QFVTI-+-DJeRLG0=,d&@I8]LP175>N70Q:-A7Rd#dM#@WEWg[G
0e)B,,e5W9OAD94GD,T\]I#0Q<.#[_4A\ZN9Yfe^=C(;NX[/R5&BR0N,&K(?]940
6EXSIbL(dgO8E1=>1T<^-SZReD4R/G+=GN^,,C(N:)+AIZ_bEOWR0O(S@fQ8<33@
U5=@d9_P9;0?&4f552E71OECD1B(>faP(XY3?YDH5C1gF+WY?>_K44TV@:\6HQEH
-Q(:AZb[QQK.PS>]00_=P:VRLTg/ZN)^b07-/<@8\CKW)PH1S1bF6V(D,b];FSX-
R9]\?^DN]=[_1@47E@8B([<eWW=[NI-4181^0Ka^:XI&99N<24f/g5R_UVNRW&Y?
@)>Xd??A(QL0UPGcU#_V<K\BM2(2A=7EAN_G)]&eeMO;OM2IK(6c>V-M[)RaXQ/d
9N/NHR/&g1E\da4dDUSURB4f75BVNAC>LHc<+QeC+O,NJ^WZ8\aCQXgT_UHcZDSQ
,5PJ]+2JCDWS<T<6;FF-][Pdc19Q,;5KE167?XO6ga.YMTbJ;^e>^+5H9.12Pd8C
a6AR>YZ)[V0KI?Q+>eJY_ED,;P2-LF-dKecJS#[IM5&#dGNd;\^fW7UgcQE8Q</H
fE1UIP1THEEaUWTbRd72R.HVV>^VCO0:0#YT/>??BA<TF,=3cd<P_W&S>b]63VPJ
AE=adaXXU@Yg534,ZJZaC3)/@2B/-EE\9JJaY.LG[,U0d2)=PEF>FXZ&@]?\&]9X
[@KO;3CCLO]cHMYL-8R#5Z:P+GN>2L6aXF2a#_O@;;WG1FY,<TY8^aLJ3V5)e[FZ
>I1@C\f,LU8FM1;@Z(8&e/7)=<S:EP=4@H[5]5](8=d08,PASJc0=5MG&aMg2?_,
/6gQ.]H;_:9RH;3+O;+6#YD;/61:HM=.1KaC6U+gKJfB&BQOZH:/V?6f:aVB@D;R
7YX//HYLX,7+&)1(gL4+R]bdG]+5dIYQ@.9MWgJ;(]cB)Z,+a(TA8cR;C-SC6E\J
/+JV]:E)>+Q\PLT=RY\.+#c?Eg(K]?B25d,AX;6>:.@G5R8BRWgAX4@_Sb>7K?I=
e9Gf7cTI(/.<7CTIaSR1/4aB-HJGXDRee@J3aI.1)Cb9-DA[3=eC=))&gBM:_Qe]
N0/PbVb)dHefKKa6:YL7YVDLSVbcFf(LE7LCDdNeF>;A-0ACFHc\Z<;Pf3TI_P0P
R1.ePgV1Af.4SJ<PV4(LSQL>EDYXF?f(6;5dMHI);A3eR/aQccFA.aL,5PWZ\Jc/
9K0QHec5f#^8C&G)5,]/Z<LcX&\e\PMEGF5)dP)B2R)U(YY64NS^>,9B3F14_(<f
TI96SfD86b-EgAD#bA?+JB_e/HdEW4A1J2VBFb@LcVTcc#FH8(V&3RFUV/&e30_4
(0@/0<F7WD>U.N[5cDf-N<QE&0Y5HgPTgZ-=E&QA,6;2f9c=//g4L=?3&EWS\/8_
8@:8_I/R(<[6a6#L9dGPE4b.92WPW&e&GZ6U_f0+?L;GCM\HO^e,G(K#+;P4eb:>
_7<+dYdWeW/&,TU<QJQ:;24IC.8BL<P5-(VL&>4)7QaQ?]@HCN=?dEP;B7==KGfb
U0LN9R=6+\RI(TP.Ef/5bO8gSBG1O_ed-dEL^CXcc_/=;0=Ka#_6F/DN&ce+YWVc
5a=XKd.L&DT@U)9bJ<.7gS[BAU;+EI87ENd23^2@7f_bcENH3/QBK:N.2V#[YX9D
]P2acc=,0A)/G=NV27,^\KeDf:CI&K5N..8.VbT=f.<_311Q.6Z#1Sg]]/8N[3@\
_Je0-51NA)S[(K(N+O:UE-YD1a5]74UL,Pd\>b2;RB)4@P4@&K-ZC5WAVb&R:C99
V]dfD1;/CW8>aK:\>86>0ZKC)Y+g-K+YC06Q]6I4O+[X8N(e]aZW/O,<6a)fJPO0
;b2g1P[QGc-KL2);+CNO+JX+V_BAJD9KH,g:/4UgAF48DM<a;]:.#3?T@dee1O7[
6IE;EPVH\-,E91<#Q3)2LT4NK3U\a]6-WaDC&2&;6P7NN2E0Q?Nbb&HVGO\T_-(#
XZCgO]@5:>?N4B,N#7(U<^BTPR0A.[JU0=gNg(XQ-W=8IQF/N9?BTH&HIg73XV:6
c0]@V/89XSdKKc:3A#;b-@0)>WQ67AgSb]ADf?G5N9J>d[(d42VL\DIY3OXV7cKg
ON?Y.KA1F(bNQE0G<Hf^2()0EYOQ-K/a_\8B)]I3H3Ff-:9S;(-:gcP>TKb8A#9^
-LeMO+YDW7RO=UWJ=TW4((#I-eSXMJfZCAO+f/PID^-,4#YbeZU^@^C>/AE]PHb:
0W]2_]GLHSXaHPU?d.NOC/\97Eb1(R^b8D-HP,60fR=;OT/\3Q[e8&fFMbA.RJ3<
,fD_O?=2>,+[?EP)-AGK^Fd\0\Y(^3F8aMTcCc\J/BQ)>Va30.E.7(F\5<.0D_X@
>T@(\e>^LJ<0D8)<J2?KO>BFOQ0d_,ZXCE\dPgDR?40bFdgR;;ZB-4#HNe:7WCT4
Kf-VJOZWCH=20:&EHbBN(40fY)C=Ng7_3XQa)ZO9V(R5C709WGNf-UJTX]T+\,J)
Yg?DKge)f,QSMa#d^][R0W-,2SXZ.C+\.K9\>-d-F004aA8LYXQF.a7)K<PA;dF+
g<:R)JPO>NZ0[I\_JW77B<8MW<:e&f,LM)e0U[d/Fe\MG<(Y:_:4;Y6_LZ.5=QWa
#HY]Z-7g,?5DB(+C^>C=GPW.>-:cW-QK<+-a3RNO5-AHK#?c^URVg3N?;XVNba>0
3<:/OAd_(S)1@:]_+P;1S:3VLdWT-O_T7WRd_+444]HPb\M.DFE\EOF&e9<8=FM@
<gY][A?ZReO-D)(;(0&VZ@E2]DH8\VVGC7(2S]=R,L.4dN4.#/Yc:.6@e:7Z/7A?
A57\-\5X-DdDW4R_61M\(.RFGQ30VI5PZ@b_Ue>&[O+_YLc;HWS#N\&/CMd\,,,M
/c0=,RQG:Y9QNL.R4YZ80#5b?[aXS2:6&=\CfR&M)<#MF^R1?W\H\JE\^Z2((M7C
)E^O7TOO[DBRN_gY#8X2+#K&QD@U3g+3^]Q3QOY:O(AOVK.X5(ISGA2-Z,(;P3V[
.fYO,Le7HDSf^cP(U0+[A,=5#QWga/Y0-YbDIX003W7bHF6^HL(SWc[9F__DU3:P
3C.?F(f(eBNCUb:E@]XEBNW_[8Z]G,EeO;J\^?X@cf[Gb1PJ03S;AR26AAA,,CWB
GbE&&d>.HMP4c9<;P-8fQ[T=Q[BLO^W)ZB_Y7,P=7XdS4<e\]g,DGb1d[XPHJKS\
LIGF?U1-ZRME\=@B-QSE(=8LdB2Q0(I55ZW:S,/U]M]a-#^W_QW(Pc]>8R[U(XF3
0NcEG^PfG9CFN6+<<I>19)#6/^Q[SRB\E;:eA#)T;1cNc+?fSD+\=G]>CHf9,1,S
6eWa2>TE426(?7]<eLCcd:3e[MT#B5cP>EFMG&(WQG^7D1<V0-<PWZM:gQbY(dbI
=/P:\WRQ>g3C&96TMWZSCK58)P,TI72AFM9/c\YGIBZaC:ZRB<H>[MWVKeGcNYMV
CA_ee0_8Jf=QUF-3Fd,H,G.KQ8Q8/P(1&)E,5g\+f6Y?5DI=d/L./?-;XgA#A/4e
_386PVc1Dd2^aR.,.VH^0DXM.IZgMH;KX;;M(fIOG4SCVacK]dX5RJ#ddAc;cfQM
GTMTR>)L#S1ML:N9F0^X-6D054&@(+b8H4=XJGASgOT2Q_+D/O-aWU\MLC?S7<8>
Bf#@SBWHC1BYT#RAKZ3;HS/f_B_A.d+HIQ)aHX^CJ.]:WA^b<X#0H6J/U=<5QN2=
=]S<1-bQF+><e?1;V>;K6[)cGUC8;g[?X@:&,5H<<00.?T[\f@[BWTL9+YeE&:]W
]T=+Df=cC5,B;MOP6f[5GC[MS^9aNM_:fTaA2L[F^@BcKA]6.\)ZPVE#5F8-#_+c
:S0@=3(0JW50R1H=99CIR-,?a]\PS@4@Ma&5GY2+03\T[W#bHC,-(&79G1D]V25I
Z<?;cWbK;P<[LBQJFb;aZ=6_eE7.>&\44\,CGG\NT;T?/:U&^g3:D:f/_6+>0V1H
c=V7AcO[6SDOeP0a/^?.2-)eX\9dS\O[;E,UO#/W4F)OF[b4FIAX#E^7P2_CQM)C
XDAEUQ9/+B:<1?-1Ec\b-@-[Ad<1M1b1>QK[34XY;C)eJ-f[W\5Kb\R,bH1Nd@L<
:?EFZD[Q?#E[KA_H5&_RR(b-.REcd,0IBU+QYc[52]+\[6HCF(Pg1dAH/YU34=+?
V7c6#0bDW1K\UX^be5DL+TAIYW,]Ve0g,S&_FU)M[8C(bEF2(cc\W).?KBfW<P@6
\J8S_3D]E[cf\5B,AC@E,f_RCSHN[Z_WKY,RJKQG(&faGbE94XfG?KK#:fII].fT
Z20^U/gcE_?,+ffE])b[dDMM:g3&]U/4D1&L(Md3RQK+E>,eXJ)gBN+;<X5fD3E5
D0X/<(UEE;:RH5W5PU5TKW@;>0@e76)KW;D;EDY/d>J9LZb>F79>\QM-Y@.>V.)D
[X@fH^:F5OZK&N40Ma):d\J=^VM5;W/Y5<S_A0W9ZgTb)bG/)0>1d]F98-1f]V_\
W:T,)#Y6R<9(]?11HD?Y<8->>A@OGX]-;AVXA28[U]-g+.BV_e>9ZGc7<0-1W;f<
fWJD&=^MMQe/aUD[+,&aBE&,^:/b[ZS3/^SHFaa<;,aQf)THe6_P5J/K#KbI])e3
<.<_DDI/-OIeDY^d6c_/;.;@cYY+MG74M6=V#aEfDIT;c@a8>fSSX36RCZW__K2A
ZUQ/#ZNHPM?.W\G;Z(=&_/(H6P=M6?FG])T9b:0+/N\gS>4&KXN[I2@d]eZJ-=Td
A8C<F0OgO[?c[^K&CJ,Bd;GcPV=NeE1UFb#D,P-P(6CXB][3395UR?:e35(QPRTb
_b7/XE2aAPD-\1Q1GUIEV_Jf+.Rc26bW).f:?#?V@[=MS\Y=?g/J,\g0\N79VFgV
f.]HfY)M?]5@]ABFH:/_FVUD-3K.Gd0GR31YE,D>W3b/KS=5bPN6K,(\O0>8VP00
S].YE<FF-e)bP)IUQK:4]+I<_BB,];.H6U?N.YCB^S<X:Z.=;5[P<DPcC7_c,719
8YG(3+O?Ja.^LI8)&[[YSaVg]_a38bC(9:/1^@_3;eeUIVIDQMM<-2+#R2GWU^Q4
/>02BZSZBBK>OeJ#8fFI5.Za]S):HVF-36U93[;gN+.dbWS>ePS.#SO=7Sf_Z58-
4#&[:1c#C5,;Lcd&<2?DI2;X@N3A=3MAJadVd:Y5Z[MOJVX.BK08^eS(fT7[)_CS
Q<EGVcK3Pb,U9C^)OYFabJ]9PH_Sc>G#eRBKUPZ-S0#R-gea8/XZ[97SSZIQ93cS
^E>_=N;MK[Z=2cNc<eDMaEcf=f\=ZZO3EV20U^A@M^PVDQ:C]D>SPcI@(XDPGFAU
W,F0)g1E);2<CUC(N@f\4BK&A2MPT^1P>T[Y#9dDKdEP_^K?U)2WNC8IG&?P9RM\
gP?Sa\GV=EMOeT,F@UXd3Pc?W#\&9[c0.Z:I;2)2DKWP>SLTf[&1_G1GS\/4_P.F
2-,@YE_6<Z#1_)2P23=<)c8bGT&<65OGJ@df)c,T=g-b7?Db7#OWe+Gf&Eg:.<SU
]IVa,(Nc;OO_VPe1[PCbab_f#3/Ce62]QA0CEBgK;HEJa-Pfa7X;e=J[L7(3+E&e
&cgEZg,]HXdU:S:S6F)I1aY@>?AffAg7BU_0#HAC^>2<67gIV-:/32QF[_TMc(=&
V+\\XYD/]M_L39aEg=)_HO[^G@62.\LDX\=@#3E@2bT?@R<Qg:=G1A,85X+D<a>8
)b/9BD75;>/4Xd6,5Y9:#H49O]XW\Tb+OgB1GKZ/9397R)OBB6JPdF7W:O(?PB(,
?<BL3\F+FEF4C)APTM]&_?/N?KI6;^A6Wg0#.G:L78S#A:?YJ/A3I7Vb)bH:;,:#
2b\&7YDgKFY<J_+/bLWTc76&78XMTHI7\-b\b813HcXRbaaVK8MY1TUPM]K(EBO<
-M86;IPZ\]QU9fB<5J[fYJ)a+>C_4L=D<a@R95N11:gX>ZfC3^.O9IA7b5B,9JTX
3)2BfF2+7GK8&[QQF+e-IJg[4aZbLB<5/>dYf]K2[#HUL><b@I\&O^1d.f9CaX)9
L,-OGaCa62c:(.#8-E9g:(PH#QG);]:RNIFTc:OL1Y>4\M4GX7:1&Ne3RH6,P/2-
gG\Pb<4B#12S5eWYBYOHCZ/;IgR6>Q[=XPFaP[P0CD_A1FY?E0a<7-C//F,4,O3f
01&R@6CTYM+c,)XZN3a>\6^g>O/CGK+9SFK,IR#VHAP(5YX0-3+(?TDX;G#dP:c#
516=b?J@\c@AO1#9;LQ?VGUePDD+:b/Def@W7UU9C>.#C[[aN_JgVPLg@)VU\-;+
Y:@5)@]PG@V?\948gC_]@_NdD7GeNDXQ;_X\C_6aN9B+8,cA#^].R#J-dT.bYN7[
]fZ9[I:[95^TK7eOIZ\(KR98,>eAHYgBQ:8c.TQ4PZWE=8fQV.f&=T1/UN(KDGE9
2T9f(07=^+afG)2:G_Hf&N0cNd7TQePRRbD(EReNU_[d8-A-7d:&eIQ/&@0+&I.<
?5(D@98)154/A7OV>P8^V/&NJ9Bf5GcC0XVN4dVMfc.MX3FE2T?eVV89.&[ST]+6
-5-NSQ/L78d36.URXD7/4^2[/Oge@J=OY/;e-#6EJB9F9O348H6/M7>[R)YBW:9O
TLDI3L.G7+MU3^KVKc91PB]A=@?&=\ZD@BAcdVVKL7^KcA>EQDG:2=C/51419_[-
U3A9cG[[OI21V5HIG/IKW_S(O1;MR&Ec#B+S_E:B?EGHCZdHc;3^\d6X74F-eBIW
AR)ZMTUE\[)F:?3RV@,c?AIVbY:UeZ38^T;-.SWa77H.()77W?0dPX:UU9IE_H#0
8\__&)abDcfW3)6aTKSNG=-;E<H/]ddF<>e[+-aA=[gP;cFX0]A?O.@2SGZ/O.M8
_NfK#N)c(:<-]=V7/b#0A+c0f[EgGeHDL+Se+>^WWN;-C.RAFDX)[L:O/OHIDIgf
4.2.PLXW;V,Gb8=]a2EBFAM4Y,HG\G9VK/Q)\B(<29;;6\GZ7V07,5L<U7Q1<Ba4
5A&=^adG6bC.^Hf)6N_U9>GD6Ka]ec7(1.@OLEG;[_2QOOH;J.8\#ODMV-L#TV1?
CVMR=e6J=#&TZ[(1J.\MW?eGBSLM]-[F@fWg9\4.]GUBXV0b9=B?E9c,^OO@Ob/f
I]Ia^ECH[BLJ,:8Q[4S+\TXbHdZ\dfZWPC0,.R_b=.^_^dY_9Nd/+[TNH4L9&(e.
4DJ@Fe&\/[02C9OeD)4=Z:KeX@5I)DO)dJ.,@DfaH;g(?R)1fK9A>[_XA5XbW6#b
(^APTUGb]T&SVP(]2-V?V2bgW36I6dN1R\4Vd7T-CZHIb]?^Y]fP2c3bZ4;G]^V6
aV@X<FgG+Xg1S.:AI0/95/2OXHX7@7H(Z:D<C09^gWgA7a]KW1:.Pbc5PJ#7cDDL
8E1?N+<UYA6MfdcB3EMN[TcTSZe((28S]TS15;9FUI4-DEP?G?egQ:VYQ,e6;R\Q
=56IUPM8A+PNX@=#B7J?AUT=2<#AO@P+3CO1^Y\D[YefeFNa8d3#ZI>LAKU,V6gV
TNg>W3)Z+&\_M3f2&2;;UK2^F><c8[fLYQaRFe;.U_NT_8=HR+5Y)MMJ&O\1X[WN
BYY8O@05&OW8&#AVYga@Ia&?JWL/6]g(-0X]COIDXba1La7JTVA8C_Qca0IRQAYe
)<GgBGTbJA.c_8=7>,9&EccT1U=47e\PSI2/,BMN@Q;c3YdV-PEYD=eP;^W6DK3#
bdQ.#-X)Mf&QeU\Y?M7=&7]aK_3BJ0,5eRc,0.S]VFJaa)M1^E)V6;)bSU(@e@GJ
\<>GdJIcD,<KdFIW_[68Me_gTcMFFZF73KD5e(7U+3,BgAb62]6RO>@-dL_ac=:,
7f(g&6g6EeKD#<ag;F:?7,-U?BE3P-60AJT28K6I-6F2:=50CU?;=?X]^0])V7X;
G@,gZ22,Kd+;(@a;671&I;T.;\8aDG<,6GP-(9W[VBWFW#?I7c\MAJ8<Zb<1cK:W
UM9IZV1&:N6XO4FX0Of7B1;EY;>;#:??&QV#K4S3dFZ,^-:aY0d\41?Q0F,KZ6Y+
E]Y.f#cDBfg=F9KI5Q5DcKKDJ[cK,Sg<WTF@DN^0&U0MS_g,,,@4AOVVc;e?XgK(
HE)18F:L5ZYB,(,R\097X8bZeKHCMZDG:B[B#>2[eaYUPT^L9Q1cDEZP;a84&0+f
WZ+94H\9G]5?^Z+RE;_G^QESd/T6.8[d0]XAGFe8.7E6K@G@CN&@df6b_]:^RZQ8
9A>QL]OFF<BY0BXQbK9H3]XB3Q\DH>]M1\,ZC,B/<W6?CM1ASQLe1)?0P@I9,_T/
]I+c2^1>K60<I+G\>?I_7]\^>/3B,A/2YDS@L4-6&23.VP.85ET&<e0J[MDJAD^0
+L?_,YbW,D-7NQU>aR5;3AF3HVH7?IVg+O#J?I<R#;P:A(:UB73O63@T_gfM+8e?
M5J=14VK]<gL,(0B8AR12F[@R_NCUHd-ggFUV=2\/TZEA1P\&<3b4A8e3VMJ6Sd;
eS6@6.gg_E1TgV1FESe;Z6dYA0EXeJ_W\9CcPY@6OS>c.L4c@ST=W#YN6<OaYP7T
,M5MX^9GY.3ZIJ>7B4C3U^C48QJ2LC8[JJ^9U:I:/+X8:4O;W:#DIWf1;7/0L)7/
2)&B#JIJ[6CdWc/fE(fZMfX>T\+_+AB)7M4X^bb2Q@XR2=A:Y\J,I;CHXHV+WRgD
9<.O]?(Z4)A.:1\_J^I[4Bb?HE3I_0JbJCG][>T]bT1g0UWH7WD9>5D2EAM;K()/
_]56g4[P>e0RWVR.IbX2c^9.(#]84e.950&E;.3/S\^[P>D#>MW<RGGH?M7PX>R9
.FV^^RU)Q[@=EAM1LGX11bA--,KdL7+YYK)VC.\3(e2O1<I;AU/&bZ,Mg&:W?gdA
_g3UbT+RF.I&^Qb54T.KRYVT]G_7VC7ZeNSDe5+#XW_G3=]TYc5JaK]X3e)fY.c5
U00>RRY9PGe^6?YB^2Cg&D=Z_V0=_ZU-a-bg<+8FQ39/RMGF[;DT9S2/Z1JM8/XS
_>U8JL(H:5[>TUY\08>f17L]B9;O1URV&QR@f>&1B-IDa1\PbOU<<:,fWIR;L,4.
G=_07SF[YNUd?Hd]H?5bM\\VNg.3UR/(P#Ne2H/=5&)(Wac]dGGAYSIB>\MH,I>M
5YU80c&E6,T^>9JBK>O66Zg^f7FXK[4HKU)EFGY)fXa1ARX_W#HA(@;MLcAAb(70
Na>BXN6I+-5A_L9V9f2./A@HQSe4#@&e/UNeO=T<c<ZebY8f[SdAPCN1SW;?6U)+
D7IX#Y^Q5C.KMP?_/E?(Og+K^LZV7f(P,GJWDL)X@3/F^OfY)3HZ1d:E5\=C-d#g
eYa6\.^WcfJV+H2PJ9,YG;W[6dMW5>d\/6-L0I=M&0TD[N3e;.^&?IT/V&YHb>&;
6PV#7XL30#NGag:FK34/&K?VeOZ(V\HU8_Z[P2f+)YO@>B&D>P3-=OPW\^b;\:PU
;Mge[#58SU)@;U/YHZCf[3VE^YQMD-CGVGGVC5TB,fC@)/&&<JfU5\^638J>]RYQ
6Y3bNg83_cP33Necdc86cWe)9X1>I]1+15;,(X-D>JfIKPZ6:X_Ba,S)dVM&E/G:
K1[GTSV(BcO,<7@4A0OE/>BF_cE;&]?18YHZ3X.b@A7Z769[AS/a82+]00Z-FC]U
[b^Sa8SQ:(N/-69(57E:H3(=4g9KWQQ3E+6P=1EOL#EC5])-d49,d5.gMEG8#_;c
S9W9HbVT=C:Y5;d@4[/5a863,R=+Fc7-LaL+;OB:6(d7#U<b]-UAAT=?5((Q.#8R
W-5b<58OD4.]S/V-,DXPPZ-gIH]Z)8O^><=SSWcE7]W,]@EG/0.HLZS91+0JgU=8
I0)7?I1a[9:gb/+I)?=WB;/Y(7KVfG4)b?RNDbM8Tf<_9]PA>D2#O?#3gB+M(S_3
\9VdAZ)[;[L4(PWVJWADEAM.L544f&/O4;Fe6B47XN#VM?:US4V8+PW>,L4Y,8RD
D\5ZJCS>LY62Be/gf3N]4V#JQ:(]e\W?APTfY+-:c3^b4g)2F-Cb).X;7.-g;S>5
SV4eO2g8>]=LaJJ2e].C_P2.B9.+AJKO^P^@#Y_JXKc<FVB2KLcVF)I8ZJ.&Lf\<
U=W.Fc/#6g@GM_IHea#bXd44<J9I]]U5Jf/E5aA3FcOX<<@dgaVfL]gA^GT_Ea^P
QJ5)33Y(L,\J3ZJNCJ&]2<=Ab+-1Y.Ob<9KFUX<#(:@6dCa3Q<]L\K&V-?&f@JL(
,QE7N.;&R:\E4Z+_F/?K^EWLN5L68#;/\ccT^8=KZUOZCD#e(Z1G472M.:#g+9M6
+d:TN:?;AP\gV,<,B:HMa9).(8fLCHL&cN3WD#_@^M[:7]27]BU^FJdVC>FMG)JD
&..K.Z5g2CCfO5]D_O(?Wc&TM5E8YQ.KKc2(LV,HVa8E.YY2+28AJ4ScRZ&]V;4W
eTU@NFe7VQ:3#cDH0RS7^4,-Q#QKcK_aA=]^eJG>?AR0INBBQC9TG1,(K(1-0_YA
G#)(]O:=_NR6[-O?F7<B]1)ZJ=P?3We,KYFKTafc;<DN12=L[48L;A<HE@A;aM+M
Sc8G9)CG:bE7Q^\G>\;<.J#9c&^(B(2XH1?d@JK:2;DY3-a1-0QI2UNDf1.\O\&>
.<->8SR>Ob9TY:F65BBaGf&.HIP5?3WX92,^WbaBVYS(P?0X-.RfZ38N3I:1d<E/
d9D64GJb(-Td19.311R5XK7ePfP6\#80ZfK/L(5\W],P)]BQPOK5##9_LZO^EVH/
NI,>SA<04cdge<4ZBIY5+Y.O(5&/fH8=B:KOT/7-P/;EE7<3,_IC.N(N2K:(MLZ?
>AE9cURDQ;d#+8][&(4YRR;[MF^C5Ab,;^]a.Y#2S&P[&/87ZN;AJJ6-DL5^O=F/
O\U7DWGZ]OTgS4JV]]a3-WV48JO&?8,=fQg(&F[0S)N6_BV=<WC>3K23U8LZ+T^2
YFaSS\]9_C&PcH<ASd_VaF])Q?M)X6_1?[K#Q;YR;CIMEK,HLLB4VV-<,VeY_B-\
5>K19L&(9E[<NTd>8APCP()=V8&<2==@b:_SI@35V.d36(C0MOEYHUa7#E]:2SV0
2QaRNH<X1DffJ1H,6AUPREB)5SL&CI)E\d.DW^XL56-C3EY[[DLLc3@Kg=b&1a#>
TSc,ESfKA@gSY>ZM2=d-N5[g2):Nc6c)5E^=Y71c-QNP^2&33J,g]1?g?9>.G24d
Eb1>[JZO/K?Y.QX0cVSf/A]Ad;-36UI5TgSf^eUK>(QNYV?OBS,WIO=B&(>L/L.9
L&g(c_E6H+RH\>Z\[5N0b--DZQ<A@a18&]KT&?_H_QH,E>f)M-L/LS]Hf3YX<>6)
DQRZ&cf,Q5aD/UFc3BXMKH)e-._&J9L-,\QXP&V>RQ---GcF/T]4+4ODINWZeJcU
1GT9eU#L1?BLBCO[X.#cdB4=:V3E2[=7XPGO??35XF4QceQ1fD1FeIZR97LfZFX:
@GNNMTgUfIf98^Z3_[0:?P5;MD>TGg01X(gd?3O:^#BQ5ELSNYT)\BK/g]T]K<E\
a06KaL;9WYZ)?LX9fH9=/KDOK1_R&:J3a/B^R,gLd<2XGCQ=1e0bBP)R-1,#71)]
ZSZKcJR+R:=NI9HN06bL&Q&e/<,IRRM,W:dAJbLW0HHQbL\&09P/g3gc\E&#=FTK
<#(E16&FK3N<Yd:/U@(ZE(8]3f=8<52^W)C962+.5G@WLK)#6EPM]NbW3XYJcf5S
ca]PaZ76[.BZGH_?]cI;O;EbIM5XTbe9D_LgYTM2+\-cF7.\7fgO(<59MX=aL;TM
8>9D.58:_GL\<U9]\ZIG_3J0I0IB(:)cA+d11H,4_8O-f5ZfR)7.YGM7T)bT7O=\
YP^R+cIA43]+GP5c2-E.fB]&Dg0Lcf^:5-(^+R47[QE=-&H>G>g#T+[46[:AGg2[
A8VL+7ZXO?=aF9C)g(BL.^/AZZ;UC)d9(E;bcR9g_6?0I._LY\fVMW09bDK\D9]E
J:Y=]GAD;5g746=[GFGa?OZPYc:X3U#/9>4PQAX0W9ef[-X069=0WBda].dcbQ,#
J[e5E@O([e)YMAV;6E7XT_V;=YdMNSYITILI^E:[NgJC#2EV+IC0OG\S(-QH^IXM
]J<KeWN<G73d<]&@HK[-Vd#:Ed3Z=)VMb=3ZYEXU3?<<QW)V>X\>d#RFC_?#M8Dg
@)He+SG]^b&&_[c[71E@<(ZJC9R\IC?T<Y<<+BCE2:E0YVb9C74GM_657-F)[4/I
5-G5=]258gMGa#JP1;e9)=]\c&&8bH<I7J>K9JJdW0cbFQ\FAgR=U:_BP-;cQEBV
,>UR4VPO#02]ION-R\\A#&LKg&Ng)1eMP&[1aL)7O?EB7?McB_eCENI7#d<WTL90
&b&2IF?@8/R(_(DX6/3:-6;7DP9H[XM2[6P-9SbPRVgHL^WMbEEK-]b)O</]Y?R7
94dU#ISPN+1b8,3ZCV2+X@>171&=abU#@<a<=HY9,9:UQIP.AI);YL&0@P17OP37
KCV\3Cd\-[FO7fAD.?caRGB8VRT;.K3/QUSYT8-_Aec,U]Oc2bd4ZTT/RSLD6/H8
,,X14P=JGH0(5WcFa<P73V4#1&6\M2#-JbL3AcQ.-SXQ<\g=EUFJF4fN01T9BMRS
;TR#NB6\WIQ@faY<&8e<AV<:f#YJ6>&X&4g:,;:Q6.<FIeQedHc#,Ld]UH(3S@a+
Je2FY;YH8HM.?F3H.)TLI68c:31A<X5gGe[aB7],D<4OMcHBdd0;,(c.efNU4\F]
M.#gVf#8PMg13<_1+M5D&=SfPGUb0M_SdFcBJHE&3&<6+/#cGPeUTYWW7WFAOQD+
&(:9&]aG+B[2JR1T#aAS3J,&&52S>.=IN8YJ+/VN[Q;P[BT[/:S8(WdI)]?\65@2
eWeS359CEY@[W?<X+:T8.O;9Qc)Qe.TONgX]5&N;Ka0;S23LbYAR<]@#W7.:9DB(
g0P41:Q&K&0Q[FS?G6>cNb:U/?d4WWc3?H#H&dM3^_OR)@]57@.FVA0LaH0]=]WQ
./F#J02U3X-eY56a,BCE>>@0-.0^Od)075D0=SR].V\6ddU3FG-O1TEWaH@X-CTH
^9<29QFG7b_E\;\/J8cS=58F9,W<[#b-AVQaA6Q2UUS8T\XMOBa26/eLd#C<D?0/
R78[&^92+-;OUD@+U]I@TfPP.S:KQOQ+=XdH;&Kf7.D&f434-#.S/cbBIO,SZ=.f
_G0R6:B#&(c;_b(PT\J2ON:eJQ[TEV&5d6g4QY\:D1I\,@B:Dd1H.F[.8JPM.W(D
^dM6<OVfZZ;H^e_SDGZcEUC>5QbL:7;-LgYUX(X24XU0L1>7C_)2&BXCJGaJK[/)
97e[M#cf,S1(GYb>IC#bTL3GRc^M2./]OV-gDL3GM.T7-C4Ua)+AT,[7^)=8#U=,
M);KbIF14KdN#gSFIA;7g/VEPKC4NC[R7bbeMX1O.d(7g#gR;PK\W;f^bCc\a@L:
\OC@,1:9/T>[e57G:gJYK]UIA0Q\=XUgS(8PdgD0<<2]U1=d75@M7N7.JZ:AA\W5
-A>a<VJ-9^WE7A>200^9;ZMY)-VM7UFI+E&=S5MEGHPB<_@O>;;(4_6bPM?F\L1R
SQ]-X-Sd\e9g5B\E,.^M<gCX#]@PS9N_<B]FG?Z9:.L6/I8+V_YYUALLf64.ZP,?
J5A8JdIV/LIAJYP3:;OaRbU4-aNR:9A?b2,0R61LYII/-T07+A-1O;&)J599]c&g
W^?/5a2B#)gODL=<28WOc>[H@_WGFb)ELOc]2dZ3NEZPVdB5H1d3L2W;dUeU]gM0
,0FH)9V8:<C4EZZeN4[Re7K=J.<SO1;<SPCX9X55CVP)4,[_Oa._@ePG<]g<b.Q2
O?EH<Ac=SK9\]<?4)d@N>YH;&IcXCfZId0ES\@N;,5D@,W6#fe>P)YP0bD;<@]9H
]TWMHN<BcL,C1D7c@LVU?XOVNY70>B<:+M\cFJ9FC&SR32ad)-;K7&FB41S:fgNf
/1S<H4ZgHd>&bf<Jb^b\KNSNcN_P.bM]b.;V],d-PD?a5#TcL&38Jdg8J4(2C=U4
<cXF_&K)Z2PbK@0=989A863,P+&1@JF?_)CQ[#451a3#H0_>S:d(V,8:8OT&HbWY
8X4UN6]Xg.S;FGL=EQVSY5Nc?TE]O+16,&f++:_?-LXYPbCQE3S7N)6#f^UFbOKT
HI0KA,5=;.UTa6#Lb+XE8N,\WAC1EeLU.g.]V7<.)/DaHLH_=]Ze[A,[[cXY&RD>
4,7M6dPSN#-@2C1c3e(133V:;gN@K5;Y2=L,T/+HbAXS&dZ\BFFA1C2N/IUDaF7K
6MW6b0AgJ<1de.7?3/,Q)BOU3G&(QeAf.=IMHMN#<d<E;72HRBdB_\6,\\=F8d>C
X.R7T/e9gNRFU4_0:TZ=M]YX=ISWOWV.:1CHT,:]:/V@H@8A[fafCCS?9c:2@Y;^
0g2)@ON2g2gRBAOO7;VM,Pb2#a_2:K<6Mc,\UDdfVZ.8UNb1T3246.,WVSL8Z/.9
[UOdAT/A9(Q^8N/5=&0OCYE:8VA/#8Nf@b0\(M]HBZ-7LTg>I@E\1OD?9[=L-SL>
dX0d&T0GBKDFg@(^@3P(IR2[#=0[O0QITeJX56M)[\([7CYfW\LEWQ4(#:6:aTf/
G=IC]VD0I4)=_;T0aa1M-4>PL3?EKf8dU)]3;Q8&1H(@]f7<[R7LE)FO_M\>(_6P
[.9?K1_5FGggcZRDYAD5WYCRa+#HgG;LO.B27N9,+B2TdQQN34N(X^;\<_Uge)0-
B@8#@KK&(\_Xb9WU=F,(6\WWA3.T751-:f;6#_8&b^?>:7J/TN[\RR94Zb0S8-^R
@)NWY#@.CM0fcN=<@bX;(a5&M^D0;#WD6Xg:I1O<V/@+cF[d75N1fLV8cEMF7RdL
gL@WR[?GL5SUF_:P<2VcD);[+IJX1EG?+bO20<7F.SaU:4KG+JRK[JJS6HRH9).4
=P(_DS^TB+[G,&11APcdgY,8]6Q):K10fU6+Z3ZSdT..=B.5S3:IQ@>3f?,b?E=:
a(a#]9@TaL1]L)-WYMVY.IbLW0#F/e-M8RV&H=T4f?(>;7D\;RVI)37P9JcE<<LW
C./O7E:<c;=^,J+,\@cd]=DTB>QIG>]P5AIA1,1C\a<-ORfRJ9=YBbH_#]<R\44F
XI^]Lf/.GF[^93?MLZ2UOX2>\/\KTfNT/I2J?L9:KRFc(P:K+/8#X6T<AfV[1Ddd
FaA5@Q,XM,]eUFO4?=PXOdI^\8WF-OBf.QSF;bg/-DPJ.4:^C/+;I\0S4#YV3EAA
fE.e1B1G]3+LVa6B9W[1CT=B4OWB]OY,@(GEFe-Zb3?)MB2=;aJ:C+T&CXAdBg##
SG^^BfQZcTKN+c7F?Bc8fHEP,9ePVUO7&[]PF_CHH:.QY6IV(0[&Yc-9))11&,;T
_K)d83UN7BG8K1]4_OQDPAgT_6)f\6:a<?<>5F&2BeDEcD)_<8;P(d9GOB,5KFL&
Z#7JC&b>+LbQA2+/Q9bAP/T#Y27=MJWfc/4ca<=RO>6L/f03HICN1Xc/?Ta=?K4X
J52f+#41RXP\_^>Uf#SgF;3)EF)46XDPOH\5D?bCQ(KS.FCaLUT+6c67PC>_c6R>
[(fKb5,.Gc@=f\7_/Gd(<VJN66?:B95K/Yc;//S+&7>:>TDF).@QgGHOg^4Y.T<\
_9+)g,.,\0+?2T))?R\06;Og[fH47Qc?&;7fUJeO86GB-8EO-XaITf1;d/)VY.<T
8<eGZ0[1?.L]cRG/<]W3/Mg.[B,;?[6-U>>99-&#H7[ZeO6<(X>/U[Q22JAHcM0C
]O/Y4eG&]2#@L+MS<d#1AG?3:L@(1Y[B/APR/&/NS=/f,];P.ZKU?/#3ICc>?,dE
8A\b0PD=H8W;Nd5H7L2)B:_c)(=&<_3QP:L+@TP.,U17cVQ\Q/SSa-)Ff>T/P9=]
;5T&c8401&]K73F.DgB<5PXJ&_N<J>\;P8E9U@YPRD2fHJA0S)5c_JgJL.M@B#e.
=e5^8(K09G?6V[Y.(H]67FF:ZbHP8dTU>,S?Jb@HPD)L?(PA^N_<4Uf&L2G@RFTg
cY0?Y8XGgS@<^:VIC<7MY@T7&6)343B==a,Z/dcG4;H.8OT;##LG6PLV662NH3>b
N;:^MZEHAETOF>f>JfIg6Z5V::FM,A_R,[0)WPY-&ENV]#<)fZb<(U=LF#VY8WFY
H=a4F@d#1SQT]^JZ.6J8JG,Ubg(:2M,:^(YG\^D/YDcO<MN,JQEfeOTPNE:9NcAD
4Xb_<U.D,ABQUcR0B,17(LALAZO-FQ0/DDegGY?acZ>SJb(YG6D]?GI(Y(f7M)^M
0QIN/.A0b2RJX(X5Y_d/b3DaAd[894SD7_X?PK-I[S:2AT&B9a762cF2b.5J3A]P
]YH/?N#5=_d24PT;BTI;LQT6>@a4<a#JQB/?B@FNA_L7VD1a7,(KSJ2Xgg>HW?-H
#/1EE:[)9<B9TYTSSfAgb3ZKS4T::]]=9<P?0T14@4)9NR3V&L\6&d,F@ER;B;.K
9PKP5O@0Y#UbRcf=J<1N-R+5/J8eP=Y/[W-#=BA_2fS_EYX889C>#INf&O[N+U<]
EMVNFBQGNK+9SJ[TIY3ePT+_DOdcd_-4?33AJCY(9?V&Q(=HO^c,N5;>@]3J#/C?
2(QWIE8_K2KQ4d]A9L5&#Bf2/8@./29.g/S^(R#,M#1YdX(SY]PQM.I)(4GN/.d.
aWJ?GfZ0]-ALQV4,+YZ4Vb3)8/\H0EEDRN=OC-;FGL0MF7<ZMU8?M5257T>URO-.
cW0:3IO]V-DcdZ_?gSUH_),U+VMQA,<T^R8Hg9YbD9NA.-IRFP(LOH04_/(gB[_c
2b>?4^1Qa)R@a704A_+?&LV.<TFR8-cFV?(Ha_1M(aD96[,6a36K1)Z[[V9I/-+9
(U>N[_F[>.^FMWER3)0N<SZ85_-a2L/c79ceT0(1TU@Y>de.))>XeDeb()73\d+O
AXBbM\^3;1d5YAOQUXY\I#3c@:0YK.R^J7@;AQII0cTfSU:.gJ[=2H\&3;5/_+I)
Q(3K.1#F94H:;SeG=X^ZVG)>/9da;ffMf6.::P@N?6<_&^f0>?[W>S8-:_4ENW#Z
-9)/U3FJ?_<+F)8M/3UO==<1:4f[<LMe9[&fU]S:e46+NUVK<Y[:GMC?<I9Ka791
3S.WO9&^IVZ,)>H@W8S(Z6^LFZ:YU6bY=?MC?A.ce=2&Q<T87UdAb3)a3<Xf_EW;
E2S>B>Z+#_,Fe@[5SGDcSXYYJ)&+ZXXQZ18aW]2?ES3.bI,4Y<4^,@U,-^dQSO+f
:ZK_M&);+G5-1IKR2L8Ug=63DP82BAY=-2)5BY_WT3ZT3<Z49PB^8EU3NgKQ#2?L
Y7V[?M/H.0A1SWFaVLf\)efY>^VWUA16_fQWW)][PdfPeNW0/,2L.F++,N+cU?(3
NL-O+]Z4YGMIaD?G@(9O-;@dB-AB+P3V_A/gA4=2ecYWSF^2WDe?8EI^V3_bTdX,
THF,=L5O&6EGfQeQJ>7@UZN0/aEaJSAJ^>3c46MC^U-5VbI;>/ADR9?@,25cVa:Z
6LNTH#;cF47J<329=#d.b_(#1:(&ZdXA8CBFR^Z.eJ_5B6=@3\LdRE1c[>d.eE,M
2b>;>HN9NN7cIe6aC0<b5KT/Kd3\(6b\Pbb\QWMaa)VE<?f\66GUS#<X&P)NK=Y3
QYeO7@3&_]XH3F]3#CVZQOcN]5TP-(Y9b_O#.(W7VZ;X0=[D[:J<U0BVDATNH71]
aZW?^KFF2L]&eDe5\WME]-T272_H30(?;(NbL87N[LF>0CcZAA<@T?JKP4]:2PBZ
=4WU_<K6_NEI55Ia_-:9CF(JaR1/O\914EE16^KIaA:+7Z?c7_g(<e-3Hf)-F^6b
PSO8FXB0TEBIH9/4.0.1bQ#S^A(MMW-P@;P?SD4X=S:(F(=-b>:2T1C8cc#>8H+=
SMZ3\IN\N>UbD\Ud17M8AJ\B2C-];H^I?8+779)#<>_[W\#P:(+S(K]2O#2,=.S,
C4e)HAVR=M:LSd3[QFP[ST)-<72)IMAK==b&LAJ\(9:42[2+\DZEZP,SU=Z385bd
P85W.TYFL@WC79;(EB69A2-?W#96<G.S1(RLLQ-[II5E=)+d_+CKDM5[HK60<YFf
\IV)[d_Z?b\eO0X<B_BKXXF75S)VDS(_VDd,E\TI/M3IgVC55Ab:N5\&bF+f11;a
J..3TO\9QLL<:6TF7Z,D:V?Y::MY-&DVCN.cRR&X[O2&R2ET@B]JAb&>e+K&L,MV
AD0CS_[G:ZSZSD7Q+6SGY/TgG,:#XWX7YE+5gOCILa5[RaW^5GEQ&V)=H?fCeMZW
6@.H<f,@Mb2R0LbUOXeMHW(c41#<5?dPG2)JL5_ZY/D1ca+N.QgbIZ>_-?7KBGa<
1fVD7KGIVQ,I&R.PNGP>&?-.NSY=2#@KeVdb8a9#+[R;,aaC8RMY(6BWca8ea)\=
R6>Z+F4,\PVKVB99DK-XGf6M6?&(d</JEeFNZaPN;\&dO\-MA6ZCMcM+Zf-E3#bZ
>GQ@NLO\A\-J@ReW&-1B;)2TN4a;&[90C5GfeS^35+CKNIgBLMeEKKTJVY,YH;LW
.\K6>e+3EgRDBa8M],2b>)OF2#F(,0OW[S2A8S5NEN.QfI93J@&D1]T:&9)2S[#?
g(7J]ZIWJ.#bY27JOVWW[GI,2HOga?^>Z>#?KBK0FQ#8&<=CL>AR)1A@7:T^LfaF
RfMZLIG4W(cN^FSKG8[=Tb3GCc=N\X#:<>E7Yg7SZS:YQH#e\EHbI4QVNFUW<P2?
^D]->\2a30Q5)e(]X3OTCJF,=,>-;c/[Vb88G\&1#[@D>0\HKFC2]^.7M0HC)R[^
O(-G6\H9#+JeR6NP#Ua-5[]dXD;ccgC);b)\7=ZD0U.WVaPE-M\CP0-Dc-XR?7BK
<FD+-T(<c;#;EL-BF-c(5?<F]@XgLK=XH-V9Cg/>B63<MV9MgO0Y20BRZ09)(W2G
-Y]8F)<C._S9&^b)JdBZY-\gY=b\2VcPJd;1GL5Q.EbX>((DN3U-6RVeV0/0^:+7
E3@f#a+@[4,Of6C0:2GTDOVW=)g.^a+NFd7ecdQYXYD,E?gZ--QcM^H,A/HcFM\e
]F4FMUKH^\eO96FSGOeTE=eD+T.G1-XGO205]ERT]?[c<-PH:KJbV&,<Va_7.GY(
W()#92Z[8gUZS.O_7PPIFb2AI[3V2BD7O2:Q?UNAF71B@MY<&90Yc@JM^;674T8X
0N_Q#N>b,=V:2;Oggg\63EgbcJ\]QaZdfG#OeU[GWR^<9<W+FG[8#TA0^)d12@6^
[=bDdRa4<IWB(Y@B(8OAK3dGI#V[O?7(MT/Bd.UQY,.-e199T^;CKG@2c15),KD9
,_ZZHI_E:e8]OV:9LJ_DNBJ9?YGVc3/R(+P.gRQ1TM#UTf#?[GaNOW^.PUZOg3/6
)3X\4EeIMSC]ZOEbM\KA,84XQZQf0+c9ESFg))L2:c(^C+4HKA9^8gJa5J-:19MB
FZ(R4SU6\JPEQ7JS+Q8WbFFDFL_9L&L@9A/XaaR(>/L2D5c?UJWJBKGc#Z&R&&.V
I9G4-@N2/)=#YYV:0)G&,-O]9eg9Y38U<B,JI_(JRag+8fY-+SX[VP^R=8cJ9Sbb
<=L,9_Q6HgP^4bYOA=1=e&\1bOOGcc0;#=S(#GB[.=b2L9a->TB3Xgd4IY-DY_;J
<_AZd,#_FW)/@/FL0N^I\L&(ZUKA=T9=>6Ba4]@dN4KLBbTYE-8KDT,#HdI>2&=2
0a-2B&O/+O541>IN.V/O?D^08d2O)+RWe[Le-J8b+[?^ea4AFe]?fL)G9/^^db-(
]2#3=5;4?f6V@FMR@?7)YLg?6EB?Y#Z8R@D0ebU3f_[U9b>0=Y3[)BC.C9ZG#?B(
GRK:R3K#F[\10D-G>#WW+T+KOQ;dcE1E:-09Z_cF,A=XY2Y)QDY]2d931e2,:A3F
VXHM.fS,=fL)SX+6d+#O5,&fE)\bSX:ROH0Q#NVeCEP2=fVTHIBPdgeTe\cNS:]#
b^_X&J^a.ME<;,2?8A4-Ng9+V\g+PbVg(MA94DJ4gIFQ-[ZP0d#141/fL4CT09ZH
Y9A#-FOSJQO<15HJf/CdDH[:J4C]561g?B148_UF\.01&:R,38K_7K12DYVM<La/
775R;>:D]2=3^J:YBbd]VHND7d]FSZDCZ5WW1&X:cg-53=.1LL#OM7I74GCW?PMT
TC4cB?R<&@V;I-)R+eM#RO^.+55_dfYdT;;BJKRFC<.3I0;fT4TK@]fB8eM6<0,H
NRgfBRFRRR+=df/C]Ae\+E=)[S:fJR+IRHYSZ\((cOT[0FgCK\2Y=9+eUEVEL.-f
G.R5;SPae_K(085V8W.8WZG@5&d__+SLQXE+/c))fgb:GO5478?8.4JdM6+=HJOV
<2E6?YG(YfE/P,.ONF+D,]P@AO@;UN>6=H5_.QbD-K?[)AH\3S:RH2NKb\I8aMd/
e#e\d83Q:9&+M^E2E?^W0H?[c.3T\\)-_S(1-BZ-D7JOHH6Pcc78d[DA>24QeHb]
R.V_QA+R-,BgJ\9PKS[W=^AR3-]?C[Z(+?;7,@&PA0[J30H78Xb&RNB_CJI=Rd;d
?1C##)?@<PA)IYI[a:&(LG(QL<52Z#PHOJJa&^+X<+-B-HAE:;B3&J2Y8QM^^Z1A
L(eS@<,O?J5A\:_V?AKe5eg1dHfD?UW<P<Nb^YdI\2e[:F:@W5DV-?U3f=Q>gHI(
6_FCP[7,J^ZOe.S3,.GXPKD/-NE.]bU,YcU/GKQg#B=C6&gVBYIK&U0FEgK#GbT3
d/.,Q1&N;PH-=6g9BSe7J((():(,f2(TdK1Z93g<DP>SQRBX\:/DKBM>>)4D@I@>
Wd3Z=7E2bRAA0e@Tee1B-6/)#@9TI&CT4d]ULD4K@;c)4RVI_OQ6f@K;45eX#<Ad
=AAM[?Af8N8>0K#;[3eWEQ:dW?+9fTI-c,1C@&.+2PQLR@MbXX@CD^6BgbJ=,9P3
/ANgOZLVH<71@#LD9XKc9793J&3A0AaaQADC(e-L#IJe+LeF7VEVS_L/9ZCCIH9U
OTcCMM27G4ac&(?b6I#bQ=HLX1XC6:6CVRNb9_[;g6g.ML&5OOgdG);R66:86]69
+YeKFORUB3AYOCG,&ab3TW[TU=g8-<Idaa<#U^\7>V(=0=STF[&R@QcAcY=0NPJe
Y=PI(->W_,FC&YBB;d6#9e+G1MW?_J@VcX7T9)GMPV)+L6S;07&,U8VXHJVURM0Y
aP\?OVT0c0WeGCZ+f+IH<IHgE1B3VQ1<aGMM(aX)4H6a7DU-QVI@I[E6MDMaWQX&
KE?N7IX@.aJM2J95M?<Q8)#;C6JU/B.@@7c^(Z#Se^d-SPI]S(T?MPZMH;Xc4PB_
EJb?]>-AY)7M)BIWC:;Wed9-.NE?:FI+Ne[/a.[-1PEb;?QRVa5c:ed^I#B?J2+L
HH,WIe34V8MP:d&IOS,9R\fV+cZbKWQS9,OI1fb_IaP<PPIY@-Y;+@NX3U\WY(Ge
8=9gU1_@)IF#26G5S6KV]8Kd=WU6Xe8DMg?78I3\VMB>O1DMR&a2-Fd/c;d^S.(0
A9&>,C4L<d5FUZ>8WW\BaLA]e,4+(H6,#D&.60-CC80)E^@0ACJG16R-If/E_EDA
8+XCOW/4cbVBg5ae;.BCPC;X1MREVcc3H\Y8>^O:gVP6T2Sc,4KQ=[;;3<+.ae<4
VM=A/,&B4<F?0U</0C\IXb]XL;+-77)?04QU2R@6Se&H7ZK[]B^N^_MPG,=NTf6U
8CUK(f@WbQH\e>V4@>dTC)B\Z^4PU;U.E9O6Y77/Y-O24:TbWc90;]BEN3(f\<E<
]BgM>A,X^-)AVa&\=.?Q4MaIKE5/>LU:&_@1fLR@=-1g#O_=:&43A0NbUOF^aU6,
/_,3=cb]b9XFg>_aHd4QEQb.<1fW(VN;g#6JRX#&_J50[0f\g;PYeL2KfX#CG3HJ
\>\1OH.=8f7>@WY#\7S5Q.<dOB/)ZTbB-[&JW53T[Q9dRN\J;N,6f36cCAbbGZ7F
527?A.WE^\8U<M@SB1CN)H_VTH36I8>3D&ZaEZ>P041HIZ(I2,I986;3W^/16A32
GTO;<BV;eCHSF5G9.24WV4J_=X)]&CF&aQ.(fD(aWM0O9UV.Q/V5GSQ>5H[1O5]P
B^S;1,eGfe_b)K80#aR81gF188#>T0MQ\[5eO[ge&UIPZX<4_dI7/^2EIf\Jd9[)
NUD>_2-V=Gac^VA\HN?28@5_,Eb[KK<gaNY3^8TC_+Y8ITFJ^0c7L,0c7E:PK_UN
6G&;6S4(9[+fH)Cf,eSJ(D,GZ6;S;Z\VAgXD<@eb(OZ1gb2cA^Q\5N^1T-bIb@fY
3YZW&eE8=@<D:2Y\.V8M-#&5A@JM?7W8]G+:]6>Xg?>]9E;U.ULf4aMT14DM&-/U
Kc^^_,AEA=.-APeBV?WB(CI&^>UGeNf[;28JR?3R]@G\/XL.]+[R\,cNQ>_94KEZ
f78ES7I7K0EY+HX[.<SZXYJ1J?>1N.<HTf(7,@^G(#cYDdGNEYC-]U21N+]0V\]1
0E.Le9\a=G[)Q+I\&B?0PUZ4\b1?F_M\#1BAPe=UW6G<2XMXOdLA,=1[g>^9F#5F
C(8?AY[PZ\eaZ-9bO:&9&21ePUV=231#:M(a6I]031d-f9)bN@VaFeNI[CH;3S2A
TG26M+@-0c3CRg,(H[Y&2K4OUTO-:]^A=QFWe8E:.0V7)HEIee,;PA70<KV7d]R=
Q:&PJKTI)O)BH/KeT].//,QYDDc3[4>dT33?H_)WVeG(TLf8C6)27;:#U57;bcZG
\K@C0d>LgV)KEdAUgQSVDga^>=TVDJ+T_AY#\P=a_,gd[Z>4LFGO<H9Y93e.4Wd7
H#>@()X&NQWZXHBLLK.g[.\BE-.26+^aEL?.<<2I#B.\,-9^(5D:OaXe,a^4PG6W
g4WMe11INT[(,3F_?ZFI5OV_@\b:+L[);JcRRM9#5-/&YX[PZDB>MWF-M6Yc;?Ue
8fQ7/@_BO(b&R//P6IUf3d3a9Gc7EK)TH0ZMBN@#92EG#X=SMVONM)4I5Bf(38\P
M7_fKdZFfI#W0Y]>bS_FX(J6_OIB[?Y-e:@GU(\U?A,M[SC13MKC?H[HR&g]Z(Xe
@:3IY4^\d-<?d;,9?9T^,BZ&_=Z;EN)0)_B@8EY_eJ73\)V>GT<fX32M/bc9T?<e
]V4d)#O&-c9:.L=G>7)V9LDU5EG8^2I0Q8]7,cO^;V(:_Q;\Mcf_?/-D9Q7EU-5N
N-)GZ(^?1bX#T9NPA0Uf1TH5Fc^/:+KV3CbeU=dH3eX.>&0=LYBf8;+6P];24bI]
DG7S@9)eeB?+M.;G:LfPI0CeHXV\IJQZ>>\Cc7EA]I=Z9<&;E,)^(QHLAXHff1^V
@F5MH90eXU<4Z-G(-<^SSQJTUfH#P2=Tb//Y/=WJ7c.+=EPL<_D:[?d28+9R<YVF
-3UGGD;<cY9<dETY;\SL?V2-d:EB?f=4&A2VTU?@T4=&+?Y?4DQSf2f-F.WRb@O#
[7W<L27_M6?C.K9CSXB,K6W>48[+:-VB6eAO,<K90\W7&9\X.EIV[;/H>YL+ISYC
Bg6@<PD/Y6VSF>P2gBGY;Lc_];?QMX)PHSMX[,?fMCM=I0Z=Og));<QYg?:Q:STX
I:(KVZ9Y9/g+HB;#J#6)/YL3bAF@e<TUVca3]8)C05&)Z\X8M/8);#/T_E0;#-J@
5-[#-I-]T?P54S<Ige0UU@BOUB:ERLXIPT8=DaG)BPL+;#gb/]d[@8J#-R0LW191
=XcSdfDN)\,,82db,CFW;bJ<DZ5TH80;)<2&PA]8@C[\Ta9O]Jf])eC;U7\2dGWD
D\G:3#93UK0YBI__f?(?RL3b-8+8HD^^M?K\/Q1FC8C+g8Y_D#(^\9M_aaL9_5<U
:e.6Sd\a_(G\[<eJDP9N/E+d;LfCaRSd3,>5LR>Q+?a9QW+c=.Y]:8@H.^MBD;K[
2_Y8\YPXfLfIUPR)Be=.fBIF?,Z1W2W[RU)5;c_G<,/H1YfZOaLT(7(73NceTFC?
TKW@YC@_6,PP#7e<U[YQQ&/AC7:PIdZb=887X4I\0SbOO\S&N?dF<Uc^b7MbJ^_4
_&KWX)QdNYUEQ19SEe+XJ-J/2L,/M=F/8dP#=[.(E?KMGAO1->#3aF7NYd/-c(?L
0Y9aB1&K4.FU:37,-gMU9f-5<=>LbAVbC>ZK7Y#:83.P2cHO0&c]VO/\7;_Pc_=J
)WFW[cB3c3E<,V<YH2R<E7)@fGW.<76;XPY-b5/:dSF=N=E_WT0@:JHe,IX=J950
3A2\,()eUVSE=XVYcd@<eV/N:JS1WJTS9.=[9A5+18G.9f,M[7BB^\?8_ecbVAE1
C]P<dXXU<-?R)98d<.]FX9fI43da:G616V/GI4BI8+dZE;PK#[U+:.<]4A_K=&[[
AX08-)J7F]UMUSG^aXQN:1W#WTdB<3>C2LAe@d5OddLCGL<E?J+Y,e1\9aEcMa2b
,IL]:]..F2TMP9MUUIFT<9#CP1OQ>=SVaC,QRWeH>/Rd:S,&UN):XSa=?4Y&&50^
A^[Y6LG&1>]QMcKF]F+H+N[.bYb(#,.ITISV,WT&4)2IES@>VR[XQFd4:601=SJ-
4ZH.ddBO[H=DIK(K+-&Z>_6KOP7g5+P1PTdgWe3(Z3L6_]9EP92HUb#LZ=6V^eC=
8=-PC^I?]UIaaaceeBFH]IXT3.GH>eVFU>S=/8Y&MPHBaR#R>U,V&4Y.?)__>Tc4
g>&39R0DZ+\:RGb4(,1)/d(BZe?I/4I,(dV^fI@X7C7,MC]K.Wd8HLZT_L?)M(9S
_MVcBMbU)7Y&YYTPAJ8[HXbb9V.SVdJ[/dLU1FY5<:88W,[BLPP(>GD9@5JT#A#;
+aZFgD/P,8U+<P.&YY<dWSc&&2T#Dd/OY\2fg1NPXBOMCU&?8@/4^9Y3F[-.VaE)
DN[NWGU?,F,?J-.6=>F0&[/c_BK&@66TRQ#X@9F9.QBe(HF:T[M_4;>D/d>bBC:=
5N1X++HAd[?BgU63MDRbd6_9H9&C@9_E7-@O?b#b.R=3FO3/U3a72@WMII-HT)e,
\[DIa:+M=GZF+:QH,B^HBUPXECS[.)T#?U+K)HYVOGRc6CfK?RSeQK-ZT.2?@J+L
5f3HQ)4?fH(W@2Ac\^g@WZO@dO30@]^9KVF3<d-UXY=?-I#OZT2GR)[@4_0J/AOP
,NW-205MF0W@eLSI@(.:U,KaC&bDIZ2&Y]@76)ZB?=Q4XB:Y(/\TQcG3:0U8M/6_
J#+S[1L^0BT33Fa+4]8M_NIE.HDBU]8M@W6HMI][8TQFaG:2ZA&)U5K020EHYE?,
3+5MAe^c8);5F:<[C\f)VPJ[U\9-=D2>8:8(?J9DY7c1YS0[?\W29UcK;FR+GN,U
=YQe:-B8^,aO2=5M/29A8=5HL2:LM_b)df#VGfZYOIAO-S&3[9IZZP;gV_9PZ69L
;(3O=f,Z-2-_JbdZIWd0A.5:OK4d>DSXf5+8SUJ<[M+>YRbKO;b4f,0.\H^O:O+<
W2O.?V>S[P^fVJH=K6,J^?3eWXWM@Y<^7Gc,I+))\NPE/N6C51A5&9XddEA>?RAP
4IY6FHMJUNZ)gfLY(\VY0fO@]IZg&YfKV>IX99gE:ag@=@(\1]B7NLb\g5VK,.#O
ga>e4QB](5a3eGC5UG<[90S26Z&Z.0ZC9P.Z#YV]LK:SB]\#Z8AJ+7egP/4]PE\.
(<9S4D/CBeQ9DcL(MONHI\TMA7H=O3;VdZ,?R&FZ:CO>/00B9/#E^EEAQFd/?d;+
[V3#O1N@/acB448ISKC4B<U9EU(KdZ73+>Z>ZQ[C7Qb?()XUEZ7:4;0c&O@7dFJ&
L0:XSGc_9?V09@&_(U4c8O0d;?R[[S7^.]+/NP2D[6#O9gA-(H&&33>)GecDP4XC
SdG5M[2LZRVMO9aBN>:F4\AL^eQT[4^581I_^1&BbRQD.Cag8_f;#F[S5(]]XI_W
BW>EZ7/Q]W0>NcH6TSP..cT8Z#.88O#_S(]-1X.0B_LZZb8#U9,G0916^Daf2H5Y
V-\_&,];<914&(+F5a/6DC?B2ePIEe_/5UeS8F6aY#C+Rc<3WbGDcc^?@ffaL)E[
W8WO1[=7,4J/K=<PgD8Ve_>LKM80dNbON.)A=bHaEKBMN63V2_^B-F<<gN2H+59^
N6U)RF#1__>XbYJ^8c&4a.<70bYXK\3cG:5Jd\&7_P;S#[JJ4&f1Td&5Dd:0Gb@>
dU_1U9/5CbO]>OVRR?,Aa9C1;D^e:EIK?4:V;(S:2D8#F.dJ/6=96DC.UE=Q@P:[
:ZOb[^Jb:GfdF#9^S+8Q946C\fAH(^LUHRGX^)3,E8+8/F<G]>@&TZCUXKR/32:\
CB[7I<O6ER0YU<P4&QPWS+A:/]OSGe-<AV]0+([BP&^4M/8B#W4A>#2N<cQUOG]a
T#MRJ-WL#WV=RWMD0A/.eKHI93.@BfW)[\>U@V=BDGcA6C>=a84#Kg[FYB\WEQA4
OfUG]PEbYJ._.^-G>/1:)LUJ9R:[X[HLU,X4.W4;4-@e+c_97ZNMbKA-a-.BPG-P
fZ]@H_UOa:D5_]-1[D9SX>35[>(8<0GZ\IL1C@MVET11f?(Y4W+5[[ZHdJ=/L?QQ
R8W;GEU\7??d.XSNAC<f6RF?OJ[a:OGBZ1N\g7XS<ceSM+@?XC>UFF9:=-@^/N)O
-^N=QJ^\RTFAG)[JeY#ge?c;)_L]E@g-A+&ZBHH5bN<#aP+IR9\bO44bFUH>#J^f
D(?7g5WHfPZKG/66WX47\_^bRDHP][cYgS8C16Y=Mf-AJ2T/a>=-<W(C]_gKa.77
40LHaTG@590e+X.&S\_MU1UB59+@7^LgEe@05(7K_W.44]c;></Y9.ALA0I#VEL\
6Y/bWgeQ.:e(21<&CF=eJ_4H^&MES\MW^VFMLR#bP8#@:Te?,@4U;TXLeQT_(GHb
>]S^RQ2>W2R+T3G:M@9#1Xf@L8LNS>GZ8WYPVI3=cZebe(Q/0O:eB:HH4D]/^_.[
+XB&(f3HR?]/V=_7WM-VE&2_ceNM_J+?JXG<Y\5?]=7PCKeFL:Y45#3>9/K;-.9.
:bP<2FLJ.7La[TIFeM_&@VXF@D(Q_)a.OMf.e]Y=AV)+DREgbM4e7H:3SEdVbbZB
0?aXKM&I[4[X?6(3C67(#+?D^@gd#O[)[2D.f9CAGdU0TNg:>g#G\=6@8Tb6K&A5
ZE_^7MgD+,.>OM0X8H?f;[0\-ST&//(I>;),c,Bb:e)]2cX@;@>?fH8DFM.LT]4[
bG)4B./74Q<5O_-F[QT8X0Wf7=_cg+VE9RKI+\-)ZcKJ,=E(KS/_a9E-5+;:XPR<
[X-fYAL[D=#f3MUT&Y9XMW:[,E>Fd]f/._gY,:PBVRPe@[K+FAT]QJM0ZO##CF#c
D@KQQ(]0F.cH?,[(=OS-I.1b,J:[=Z8@cE.4ZB5&MZ8Yg;#0KZJ(LT?Q/]EDV,D0
W2@GC5(B,4=Nca/53A<#Ra1:T_#dSJ\?J4<0RDcIbJ?=,]A0cW^K/e6V54/<P\A[
X>H2=W[\I=SU5=&+,?.JZ2UDb1ATB81I9f?M797V87JR=W)0W^eX2^8=.1IGW8f/
QDD4+2);,K+d^..O#eVB9)TeaMA(eZUB9NTGK4GaV4YQL,Mc_67>^I7Y9\LW.ee2
ee?(f[a6P#_KfGK0bZ32..,_fA\IVaR1C^XKO)[IWXcJ1b#W\PVZFEWa)cQ5_NR_
^S(T;6M<L+D(@S-b@\&SX]]R^fOZ3R0[?#8cCEa;\TYXXg/(=2&0@7?@gVVF-VZ:
=6R41QDg+(/Y1=^A1\7@,F->[+E,&W\<&a(9IB^+W^ZT:Ecd)#PCY]CI&J^?K?N?
26P34OgDYEbVGG92-aTKK.cM-CW)L,Z+V;MIK)3Xd27HM=b@N[<0(b9H.-MM-9CC
I5D[PK6JUA:dOP/@2DU80dgM-B_G2B8JLQEfS89)<^H9g\bQB?1?=G1[N4Lf-;JL
Qd0&4H@:RLL^-ODFGP&E1SMZVBCR+;7,I3SV\OMd>=2Q>ALKcbDMH,H4]8_[Sc)Q
XLdd]fCEf:A-TJKgcdK(7XG,YKWD)EY:RaI3\;[ENE+6M#>IMW(-0L[fUO01(N#b
RL=DcYKOD&.V/OdC1W2+J&B#e<^3=JUZ#IBI[A=M_dX44Cb]^FU,dZLK6?>Q2Mg-
b(#SeaI(\##@17ASIZ13=a0D=LQ]:,VVGO621LOd;3gVFWAfN65KcHRPa[19fDFd
G.N)3G5ac,f[A)>A^(5LR7KD#+-dK9[022IEX4O/MSLO]HE+21=c/A&Be+_@Sa4:
eJX/#B]:702+2C89)gc:[8-K/D.PWX<.-.OFYYRE@?b.Y-1&XP^e7<=DKBPGDLBb
4=[2;&Bc[D&NWQS:8HR6^2[b<BV_bd;^bb^\S6^OMbW5EEQUG=T_/8<)>#b>_5X[
5;N(XT5XD5WfMSYB,a.E2#2S(FS/4/+#F9bf[b=5.3GHYX=TD)>2e3:7&c5G7W?3
a#5QEJ8f=A5;(BJMceYEL7ILJ]Pa6ZH_6+=RUHED+^;bXRea8)CAQJ./@&2Z4)]L
K.9=&K2fEG</ZWHgNJ?=UT&YJFT\.))WOR/aUW^3._?&6/M^>c?@?dJ.RQ5[R=J7
;?d1F<CR+.eDN&^b1GFb;-H^g[aYXZQ3??3F_)60F,7cYd]4X#/ZJ>Y06Tg/=C9H
/,6A]CU6Ad1a9TaNUI5P9+dZ>bgQ8fG@YP2dfd+#N+.M9Sba8OCXA-Ug?&@^3Z>/
7-QME:>FZ;D_:\K]5Y9F4ZDE=:G\=TYVH&McO9GF111M:LWXM+3Ed]-[/1CgB^@Q
Ydc-#<O\>Ob8NU=4Ke@\U9I,O_J-_QM.:GAXaLb?9+I[LHDJ6aAK(c5F\TFCDC>B
M8F]fZ<)ef+bKNP0YFZI81B?Ig:TVZY_aE@gZU<c/KR\eE/B4\\1d/L1HW;]1_V-
@>3+&7,9?2].C[:1QG-Y:LCHI6If>S..0&(X5C1=6+@O;<@@OSaMO/ULHQH1Gf_U
<MC@HZ8B,W2LS\<S+9Z:N#2<^eYcA0KE\4@RKZY;).5]U72N)<ET6g?&USMP>g9+
=5YfHGM9b5B5A;TOU._W0HdOAe+_.,[_OCW51Agdb9Q0P/>LQ@YR5b;/1H>&ddHL
E5AS=aaOD_#SRLeE_\TFX7MIA9T97@Df9N&=QZ;I1NPXJL8]Pa4C<4Y>M?../2e<
#&/&X0V^V6^+KS;.@Id-\,0Z/5CJ\XIBU=;CU_6f&N[.NB8LUDKR.Y[Y?H[NNNS8
4cPL)3V;A-dYMHF:9@(F8(>N.GQS&4d_2_IBI^NF6.V6,()-4>Y_Q1UY+5DZa;4K
6O]^Y41g3#?=RDdb62YYU4;(TG^>;8ZP0PHI0,&P\N.04YV@R:AOH?#aPL14E6Z:
/-,R6MUg^1]]\:6OZH>==)<GHgIdKbO?c2N4]BOF[JaJJO.F3P=/#N)OIKX[<[(4
+P)2]eVRbT2395=eIJOTU&7QPYZG5]7IMCeQ.4A48MV\f>d9\8X^X2\W2M..)TM1
HWGNd(Y.?[a<]Mf<.KE#U8)Ke^B(D[KCCYX9RVg_D:QW7:>0S7+?[S#;(Y9?<fJB
f)HC;gT-F;+9W(6.2E==HL,c>VA_CR/VG3QSY3?[;LEQ@@(]@<>C8R@5R3RdbEC<
#P0OcKOXC>62>&5:],^LUB,5F[X>].357KN8G:3S>L#--V<JH-XR.BCM586^2gJf
8Y#MXPNLa_?1e\KU;<?EK+5^#:=@2)^@_4>_gL>DA+QHTH.UMJ)(gYGUd-1CS_N:
<9W;->MS#GW&?<@CU.d449I;G14H]N./^WMO2Cf@R[Q7Ea.2_5D]TB^YeC)M&9b-
FUaC3QN8P/9^C=?YaM<]ATY5V^LW>#H0;^.f#:PW+C&B0FMM]WK6P][IH<I\IBS/
2T_8eVD^?b(6Ge#:#9df=_cTe&_0gcd)M-I:-55??AAJQ&]_(F]@R8^/<:/.0,P3
1f]2PPOT\:^KcQ[D6Wb?GL/8CC8A\]#[4=c0XKbH;8Pd\0+EO4[8(d7\B9G&==U/
[O3fE17:ac07?F/?Z2Y]C7f4Z3V;c>\2d(]H217PZ__0;3/WgV\c9<?-1UG2bc^B
03L/-[dIg[b.,;DBVN+S],)IbX#+28-QXb(Rf@\KbKFFaS=;47R&;7H>E^9]G,Z0
U1&S-VKfG):cG?Wb+9C][(QK.dUU>PY[T()MR<]VGgI&KHRR4#J(XY,0[OPVIN/M
MEY1c,HcJ0U<LKUXc\6IP_.=AbP#FEe_MYTQ5AP3T1838>gSADO??3_;SK:[#:E\
+McTHWX#MEB=cF9)ce=C_W9]:&L,]T8^dNZ-C47C\DfBFFbW:DY&ZB;7(<<XQSFM
#12L5_>;@?QOK+#=12(2Z28^X]TEELJ#C1gB\^_Tc:_;,O4>X2Nf^T..Q4aW(PXH
VF#cFE^,/;#DXKFAb=#e)baK+#1eL.YFacea57S/Ecg]6e2dKGVC6+(d\&3]=a9/
??L=A.U\fS>-)3\IR9M?^Oe2+YQ&6^WRLM](1LXV#D5O9NA9aP\9=93=&f7G;;DG
]G\;PAe?9.)JLe4.a)[[F]+-a]7+G(.S=]K=aWY-58EV[?c#?&#8([^I6(;W?V6B
;3Z6/GS:-ZbN(;D/eGBP_P_P&bY4Db..#[#gdR;@Oec4]?,GJB8.RTTCSfBZWb3O
V.<X8D1QX9b:(V9/@420?3?.WL@P]_/=E9/eE]6+(MHd_0U].NVaCRW+[?,YdB8S
F,-Y6>>LX@B31E6I2B<0Z]GXH[C)aVA(Z^[C7:D9?:+b3A#KR.VgCH@\WQ4aO8;0
TT][9IIdcd7FK5-,g7:J#HOOH&f3U+58[aJFg-(]?;Y:FMaX/)WD.QD#;f:Z/cV2
C1DA[AGH29F4RZK3@:EVYM_\,U[?0Z:d9S]ZF)eE9@/QG13(\XbBW3D94B4Z?XU,
XKIH)9ILOOLAK+AOFQT6^d&bD_CdV/\@gQ.NcHPaBFKV40?FQ;1N]CSH8FCCAf5<
K@Vg<P7HAFFc5<K(#U_ESc3JPCWJ9Z50PP+9&F7)f\U8fW.\G(/5C:MBRG0>>NKZ
Ed=C:TPF71T4LC1,GGNTQK?:NP6g=e]Z(/LdN)e[Q]e8GW:G=NOPXP&7)/9c54@c
0402NZJDO&F\c6fS:bGBT^N+g6N1M_ZJ8Xb?P073YEIa06U?GDc0F<O>HP\H25IR
,XUVM)[#KPEF/FK^?OcN?OJ=KU-LX\#W)BNE+WRH6HE=Z]9VPafXO_RCRDKC+;T_
05Y;-6Ra02L4)\HH<6W,R^-]FLR&].g37YEU>@Ff#d97c_-G2\VHT=5fT(HJ6X5;
8KXRC22_<C:=Q4&#a_?D9636T8K<e4-.M_BW)[88=9E@EGNGCW_[D6M_GO+=e44I
N&a/G2eYEWFCNb\B\8d?-1f.LOSWNa_IGdZ##96eW:0#9Z38f>fbB3@fPS0KfLKC
/[1BF)D\c=Ed,gOHZ#M<2.ZBKHgH#[MQSF2XM]]Tf^O9+)JaA+Q.<1:.J71)YG9g
.de0GOa?IcGFN7\ab;(TW<^43M/]^8H.5QA9?0+gK+.9=GBM)fZP3.fJ4_5gZJ4X
6[/AW3e^MJ&===F5+ZKN&8V4a,e3e.>&M(4=HB6HBI?^F5LdGa<N(XX.f^:QOCA,
:_#6EJATLdCKHQWQ3JJ/?0T-NV#6e-gYXRE2\24;\OWW>ED_?YW9#<UcCWU#XKbP
-7dA-ea>_N,bDYN60(-WPLBUQE6JOfXcM7V2g;Ad:Z[RJK9>L]BB0=3UP4=(a_dN
BBB<M&F#0RL9W-7FEPIa3Z<R&C&,I.4H2U^?eP&(^?61D>Y+6_Y)KQL[Q3XIR&9B
IeN:LEYQG@V[RY5fg08P7dIJLP/ReHF^+Q#?14>e-/A2R#T,MfJL4AMECaD6X:=0
;&CB63Z<,J<Gg@M[c.:&&,YSIQJ;VJaK<IW((T>IFV=0a[3J[?&PKc;QH#)L<ZW>
5NM_@P(RK>85#6R.SaEAVODU4E8,V]@&fVT&;c->5=R8F^Ie+e4\RSBVLML<#Q]0
.&c)4Gd-X=WYH[@Ld7Hd4eLJc[2-Q(#V/&=1)PVTaGW2@-1WPVNGO.NI+d19#+9/
7CFN9#a(2NI;2;QG?=1J_0+UZ+9N&)1__,PD-+7OE8S5698JcQ<VETE?E3OY)>CH
3dND^K>K_>a<K3D5#WN\S46#Z6<?4I];0MZ519E=F(1K^.LA^gUg2N#)WWHbW,d=
e9_,YK;a8&FEP3cI[LF,)b][?Y^W=)(cQ7\R,(A&>L1_^M?JN[AO2beJe#F_4?HP
H62[IA.1<UG)B7O[Y892R;bC+2[O^KJ<\X=U8N:(LE[XV-?ZeDVSYS1\?@VAbd-.
O5;9_^Of?:8CWCVGU.\\(;;CW:T7?(4(<B0=_782,_BAeA>:[9NG0N9FZ4.C_WM(
(?NPE8QH)4efG(aXdU?]/_<GMY&2ScQD-M&F+QDO/:F&be;<:2[>OY6_4M)H.d[K
<SQ+1+/fc5GVQRI/G.8K?^2<;PV0HC42;/>VS<5UC8Oa..J:-UM^UYd]J_SB514I
^bEYG^Z<gZYG5DEICHF;D^1O#9I^[/B.9MG79b\g0#54YP8]\4Y)^cgNK&ILYOS[
Cf,&P3]VVLP7G6^aNS;WAbLP.>cO+8/)M@^/dd##7VMC,,Sc>7=?-D5=]7FQD<S?
,L9b9]V5^R4J7dca8NJ+PN>Q?b2@&:+d-^8)WGP@6Q/B/OT0@E1@T1)J-2:8L-\T
-3>]BB;CU4(#adE^M6QM0JY3S.EEe>\HfeBgZ<S-T&MK>O+L60>T.&,XH>B@c&Uf
4dJ]aG:PHcRRH5&2RB[;1Gc=^5e8fdd&5,RLOHA[_fbKIG96c]bX;X]/>ANLS,TP
D<bU^VAdNO6C+P>-(f-d;\<CA+NB:XO>_6?.80QFF2ARR/)IPIDR/WO??d5d88JD
O<PBV81>E5&e0MI2S=M(,c.]=C1WC]M#8E_#Hc/eF0gPMDQFYKJR_,SSCNV;8JN.
+Gg/J4^6cV;81\Va4Q@M>HY(M/&CEQcZa,3VbWNJEYW7&N:f&\C:^._Jcc.CB[5G
X)ASDKdX5]7#(<-Ke9;3DLH5Af4R+gGA+g@6g[ZS@S)@UUgd?+@[(f5(DHIPg14d
B,A2:M)M&#VTS>dZ\CKHa9>HCb]8(4??Y-::=^VZ0?cg3(O8B5(bJZA5IA\7a,SH
1J#;d[Me9XLXJ,.NdeGE5O4BMO<8\^E+/>Z;g2@R8-)GS-+P/;,5(#T)4[LTKM6Z
FS-#SH3EfdJ7WXXe>#O)PN_F0@bM5SV6cYD1dT<>M1O4]+bL</5H7LMLUO_J2WbR
;CB=>4a##+e@/J.0fG&D^A)U(aO=(CCQXFd=08Lgf^)0TWGg+56K6SMA_.S(\F.f
((Rd:5@2&SE@fXVAD,^g^VC:@8&IN(?@DV^Wb#^5G=CQQ_MbH(L#>@\.PDW5d;B8
UN9RGfAINWLfZL2V7g^?/0)5/#C4aF@]?_J1X^Ob^<a)L+VfRcd+?7a[6I\7=+);
LQX0QNV#I#C+)O[16-VL71\+^M>ZgdOO^UObWM:\S5^VQNaP0Z4EN-,AYA2gY]49
#M1OY3PRA9?H(gD2J?-5[gWHJ+=JBQ^+-.;e0LJAfLa>d,L[-?#P_bS:dE>M1,9O
DPfa9]8Ug0cgRYfV9]ZEd1dZ^QTAb#D;g=0??V\:.3E#^7[Yf[&.b4H>XgIX.SJF
4?J7AMLc>/RN@gAKKFU]c>2,WM/()O@QZP9/896JW(3-XY2CQ=[VPQ6^a?V<)Q,F
cM-34W/[TW<L\Og2?H9D14QE&XU9UN>U+A84E[+G\Z.?Le.;>\a>IL-.I54:>#L\
UL#P59#I:#a.N9V0#,>/^f,OTSD5Y67/A0V=eTOTQCe=f\MCcX=Lf\YR_P-6dP&9
^99Q8;=L?#S2TG#HcK?e#C6?MKS66&Wag]_4L7)K7T#^#GL@OBN#e3UgKX-N-RN9
g#^(<A_d3Je::Z;^-&;__DdVLW]/F+NP+0S=gDWZ-(KfTIfK<F1I3c336-:&2gJF
[CNW[CL@>6T#6T1g]aKU9--;IV/D:)C)cVCEEV&QAbVDP[J,:8ZT46Fc.N:ZLG7_
P-QIfZ-LX1cZRL;@9JG8)Q]\&1^V;WS+cEHE,a>e.LTJg,611U.fDIK_g_T201+1
)=,K>]c,(..,8+;;38e+EL0.Y(XW]OCg<KT=O7bTJ?dd3HY9756X\K+@/;>S/Cb/
QB;3/O,NNH4O2=9a0HHI#Pc=DS6E_a@<TddLX^ae-:V2MV4VN^fC]=BTe)6N?DQ1
bMJ(:f:MB^7&FeO6\\=Y&Ef#TW+BPAY(cFH&PYFegI9DC6#\+9F;AS&N:Q8/g51X
a<Rg?<6W@DE7I?c7NJ<4#(,NC37HS,EO)=fD)dG^\-_]Z^26-L7I=J7@=OEI,0)N
;&H2:T-RU3I+^YO&AZ=##cQ-dMg,G93^BE07M<_3NI<^=8G;&A4<E,4SX@^Xb;@U
64M<e#@d>J@9<f(.MFR>AbO_5A@X,??B?5U?I;0D83dIU[dU[0B>\H19_=2H<,Q;
)Va16PH_6WTI[YFI8&ZA[dDKEN5QT,f<DYd4NJc<T&#]0^.fa&\&D[/f_RWQQ^V)
=Q0dNS/U-LRKKA=_I8^]eYIU-6F3e^d_1@ES-U2[<SMWCT1Q>PMC=12Y4_-/#6/J
B._J]YYILA,7<+[ZdG1Z&))HH[Q)a;QMdXeFKDA^&EcG7c;=?<8F_MZF+RR,Kc.Z
QY[+QHe;DRIfPGXJC5QD_EJHP&@@c[&/4c19Kc4YFZM8#PZHfR.LbUbG>[^4e>@Z
SL+:9.[ccC:0CTAY(/^C(5(_cB):_/VJC_5)Hf@H:L;-L:@MJ:SP\42<HI,+dXR3
TFP_XIG-LY2@I-]9VKLIA;>XebX@J_[=e??;FN([@OR0_&b?gZM8>Lf\4V\@SVUL
.a2XJ\Ac0YM.?3GJ.H3-2g[W120G6YIS6X+FCb;[cXME2)_VYDQRM8>04.#a9P\U
/+,YZJ\V4V:FV<U&K0fW#54#5PN1#6W)7;4GB(TMQc8]TJ\?@c9Q+MU6CJFAFTZ;
C\)CAbd5B:cdDJCd&[IG^G=^WU_H\)aE@)C&=cR#QOQD8<0)NdYK[W:CdH3KMcI5
KAAJ]57&0N0IK]d9:bC=aMHHB6NE=IT510JYGSCP/<eI2<#@d(9AbUe<_)>ZTC6?
=2b>7A,cJaE<eLcZ^X0A,&(_[F-PfF3:(8geSEb8O:cEZ2^3NQST_U?/43XK(,bZ
UW9@-JK8eWV39XUW6()Y\.IP^WRe@9fO[HQbb+WM,fcQ)GgE,LeD]a_LQ-EXO+89
P+_XZ?KA+3fPCK9K[M=_I9D5RIH:@Y6[NYe&&(CHA(-T3QXWJ2J#7&[W4=/7PH84
6GX=3)FH[aLV&abQ2HXgF@2VS51<TRB]@5W5O8E7P;f_:ZG&06OQTX([A&b=@F-/
e2YWNeG:ff.9KeaA3d+8@a0:f>(W#>XX7bQFLb>X#(fE(8BfT0O-Q<7e#-PG23(Z
&890CdLU;edZ;IRNO]bW0VX/)fJ,[X/^JRT5A#THTJ.JOB\.VBf,;cfN<.BL^fd,
^C=e8,\T.fbY:B;E8A+Og6eG>-&/XfAM,QFW+C4<@:US/)g#SN7JR&)2RY;7Yb(_
M8G;-=S<\5NW>D\F7V]e[aZ[WaBTV@Y]c9BEfHBOT3\0Ma/@LHTE@&R((7F&5ZG&
BGHVHgN8dNX/c7+Q9V+cD+PaUEH:^3#f5O./2ITQfKD(O=Q4\Ce&PXQN?=S,>X8T
DC48/bCQO;J&5Z&aW,L2e7)ZU24?C/5<2_>MU#9V3#eQGG7\S61M5PdE-&O>OA-U
^00b7NfeNA[HH_KUKdP83W&SE\[fQYP><&5W=J;N<\ONIX&H->f5755B)\([1JNE
^\@^??WLG?Pf]&](S<GgeGBT,S(3<0-?+]VUEDaQ[?#f@E&,;T/&F3[XBG)B\:)-
5B0R&;KV6+K7LV,cBQ@Y#=aAWJL<Yc)NRX2K^N]/XW&OFRM:Fc+3Q3GC-JcB8Z^.
JL7WA+_]W/+cLEL?aRFTC\(ITH>OM/;=8NV^:Q00(eB+6^+g+;\I#[Y5bI,Vg0=H
)M1f=Kc69H_Z-gA1\BbK8a7/D8<B,4BP<Z<gQEB,+.[WB(O&UPZOHZ2BCP^KPSK)
CRd/^/63_Hd2D]aJ<&c7JQ)[L?2dYd\A<BIH\:V:OS<3:)#^/bIXWgdQ]QXUP2/Y
;<+WZ_;R,fe/UUfg?<>>(U:.FN<+WPHKAP/cW5#a./B/8^HLNZ.:X-\f>:&.FJMS
>E_<F+,-?+XOLAdJX@GSd?aLBg3Z^-W-08Z4^+]b0?QP[6LIc1\eL&CRDCN=.#/)
@A]]BIXQ8C:bb5^0@8g/g_TR521f>E@@+/I45DQ-@d+.>]H8IW?W=@J33=OHaUT]
7XBZJ_U(_-N.B]a5,_fNNF:CE7-E78]1:ZOQE:,Hg3--cb.)EEdC@=YCe;LD?[#E
B^;a8LAR,2;K:0\@TF]>)@/./<a?4f&7BK(U&N&DXK3K].(e^\;D;fVQY18aGY>f
]e83F+_c(9(.3[TKP4a?WJD@P4Ud;4f?R0FML8CV6EFaM/4.(XO::H+LW/X2Y5.e
RU6WR-RAaV#DVJ[)fCQDAP=EPTR835Y:.K?BI7ZO^WWaDR/79DYUL6R&<.PcC-Of
6X?e))]&XR0f_cKMS^&GP-V>^A8S:HR^RTZPSCC7>JGCP/6@SE46TBRM)B:C3UQ.
4TY+Fg91gS)[5=0g+\ZO/7>4b_U^M@LJdH&JI;^P/9:@])[#_P>g6UE[?2OFWO##
NT&Q<3ZHD7e_,#C@7;dW5@?8d\[6BKI7(a1Y(CaSV8ZN6@ZbScK&c1,<\)CB[aI.
7Od6@2S]+8-Lb=H:6U8/gUEF0_\(3SA0W<>^d/S<?\H[Hc-A8,/0P^PHISa-O/OS
5@<:OLL5F[P4VSS^&EFV[K2\TJT_//BeR:+Y724.-IT#X:EY>N_XA8>Y?@CROBCM
<@d2TB^DB;f=J2;VDAY1eT0&V00S]Sb>?P1H-88MKL=S74QKY^>N+4N#RHY]X[J<
OY)GLL+I-:c,269I+69Z@7#)MUBR3C:0gS5)/@;J10T^[PBL@KgX\=X6Z)?J_>@/
WG-9W[@5?_^@<#><OM2AUQd@dH/CC3WLN+&.f9LJEM<-d.^UQR\K)Z(H/+eFX#B/
JCA_;;e)18Qd5bS_J5@V6-.E.8Q=&)gM4QdaSYfWB6_:V\B\P4W-2C3X(Bf80>5[
e\6EG?gFZ.^X1I]80S+EBW/PWOIY@H?<O#-#W7J26?8\gXT\)..>dS+4^S1V;X2E
3aeITY8,7[QZ,O-g(HP]X^2[Ue^H6?NDWHH90P,(>2b.Wfe-/fK2IO)SLZ6<A>Z?
L.NEd&CZ9K<]L6JAARPE#a@SPXQ7.GR0C>PZdSVXYW?8YYN1-T#8+TaYf#=^@\I1
];CTf@^d)LTg^9\;[Z2^TQ7\C4cXg-@Aa_PfedY3/6JE9\GcGPR&g&WX2-5(F:=K
\\:DPAR/=]>Ie8Za(EAaXV&/WP^-0H=YW6Y(J@+/QC)Dfb=+#4E_R;.8C\b_a0Hd
>f7/8(V<_#/+c]Fb23a\WO:ADW^D6LO,d&3Q:2JI.275;Q@,FWa;\2#?8TO:;5O?
ADDgBQZFY0\0BTIZJ_[gI;/[4SgIBNV4?6baZZ0WL6;_V0GJ6WeDS-<2Q8\XNVT]
OM3.Z^eED9Da1Q@4XW0bG0+U#7X>\c=BI(Gd:5LT(CJbJT3<CSYUg2+Q>XL:O4:P
91R[[P^aFM11Q7f.=JAY)\e9\C#<WX3E;GCMAO8bc15:>aB9(,3_;Q3OAP,[dU+B
eM1=aD&#EGX8]0(\;bda89Ce6<NNZ>.Y<3):@VcW#KYRP]1Xd<,Jgg;H[UH]?)CT
O6@GT.>CN^M(RP=Xa1E)^9d1c\2@+=4eVA]>NAadBZEa9IY[DV?]dS6]TKRQN/1C
Z<P@Q5e6B_=aSWf;[7,HMJSN5L@Z>VSNWTZ\PJY58?=T/ZV<:7VS?e5H@2\eT73_
.bO,Lcb&PdgR>4]_-JN4EKcP^X29,U=;MDY>KXM>8YE#^UUH3&W\UBdNY>aQ8^Y^
MSDdc(I-]U.@/-V5?3KGfXL\5Hg>3#:?J1AEGb:DG>XX.75<;8BV5?EPe/_fV+&6
/>>]=a&\IFO4)3500gE0-X9&_KUY30gNe]LJ31]AfE@H4B_H7bBf^aGFHZ=SfY.<
\8]K^]XK:](.Z054d/fX?02]c]1F2)P4-FaZc;eZcaMG.bNe=#D),1BO8=(eTa;)
29=(>R]C_\OR\7[5g6C^OAU,D)g/WEg);>@KF\La@H2Ig7E8.;S9+Z6M(;(]@PcY
S-g.H@F=;R^(9f<d&Fb7U&Gg3e][.HB+04Jcd4XfRFfTFOXSX4HA(RADI17A\O^R
>ZfA2CQU]KIe>^B,EL]&C)9d+]&<7AGZd@M_c[8cXd1OH,97BB[)]W5+DSa]K&-<
I8-3&E]3(@?8(;_W\SWVgJ@=W\8S?TgWUW154#>?^dDEBFA78=NM,W@S9CL8=(3S
fS0Eb5<T+YE1(9UOZ\/@6Z_4bOf-5?5DDJ#CT<1_EUYXOg^>d5YA;7:A[-;7)R57
V)^d[<B(;FI48_]e/fNP7Q<F6Ib23)?.,UGd]Sf4QL:H#Ea+7ER[#DSX4F2R;B#H
8MW&g[JY3.(,4Hfb5D10>B^-LA/S/Fg#XH8UZM6AMU,T_a6(0G[5QSGIU/eB>E3U
/F&N2=e:OTX,?^JIb[GL[^KACdA9[[UIQ,0g9f+6/C:.d_]gMS@<GPZLU&]9b9/I
9\?/O49XL>aH2P+IU6FNGDX,PfW0Y_g:VZ6R_3aARRHe8PJdF:GK3fD)X-J&[9TG
YC3+dgE0E1f.d6X>aJ/8]CLa)0MaTKacS8KF8_DbSTdc>SFR:eD_R([]+7FGWMGF
A2&8PD;.DV\KPSe^W[J)PaL8V)>g;9dSd#3#8[RVM?dON9,)7-(e>1<,V85C[db.
H8g^.Z[I#Wfg/<OBKS784HML>d.Xf(,FWaBGT:YZJ)O+87TbgWJD(5M/3F/Q^A3N
IH,+O2UAH.RbA=-D?N.M[H9=b&0?8K9TQ.HY&:M[6\-^;E2E7c9D7_1.J.CaO2B]
GLaXT+ORPDMfg0^@AT+d\V4VG@>(2):M,aK1^B/#.79@O;LMYHU)<_#M.@+^W3]3
\&e8HP@EaVg80e<EEPg\faOGaPM_4T;MUeP:2#748=EQF10E&<A;\;>H70,H94OI
,b1)Y8?K_H-FTKJPVXFP],YBA8Vd_H;bX[3d(6c?5TWNb9:SXBNK9=FW@0X#-Z7.
&E.1?_d<Q@QY^d(5-&X_-SP321Q.TY=ceAM9XDW\WIQ9H2=E07_.AT23A^TNKgCF
W+(Z39FH6JFL@#FW_QCQ6EMJU8&DB8WeM#4bTNUU;O(;TN\(/6EZSc<)M-&WaPW1
(5-\,7bUJ#CQCHCbbF@,<cL<Z;@7A/W)@A-@V7fSQ5SO8^<gQR8+A7/B^2e2.AA)
C+.F/0=SK@NdDPMM2(<L.aB\Q7.^@^4-R)7)-:HLG6G<HD([^:c0?b+^2JKW>a?f
8H&S7W=0(+8C&;&S-R?U_CAa5O1W6RVD^^6H-cE&5<X3[-BZ<-b1?6X,,;^YDg,I
[26XR2/N7AOOL7&5[D>RR_e\=X96<&OB=S@cD.:]WG7-^2,L)P4bPTT#@IH)QHBe
>YcYGVOc?cP>29+TGYAFNfFL[Y(Q#YJEC_2V;)NS<g41ZbKa>QYQ.0^PJ\CD.J^,
H,TOZ_N)<?ff)0D/?(TFB3E;G]9>PU:[6=)^86dH2PfUb8c:g>AP.fSN?XQeN_&^
-?\^XYP]:)^;@H+4AQ_]]7V_6<G-<?3?I,A2/@YP6/;IE.?K564MSJ)\CT)TX-33
[A09MJTd_g3RUW]PeGeX@,]OQb?TPUU4]JgP/e?FISB)RF9&J?X7.Rf6e3D=J<@f
\.=R7?A::G2L)VD>J6ZRE7>FOCbNA\J^V=Bg;5b##5]&QAF,3BLa(LZF?0NgN<N_
g;6B\]^(:PU--=;R6]GSJG4OaQQERa;G:<aZQX:XWD)1WP^^KVO(G?GgZJPffHIO
#DDP):9H)<M=TTKH69Z6J_^aUSI>BI<-87LA,O45_]fAd.g76L=^_=[^4=4S>;gG
)O.GX]gbSPLKN.ZU,UbK/gX.(JPBX<&Jc3;9,#DL)(6QVb?=2M19]3-5?YNK-,4P
&NMJ?\X8.0Qe<>(MYKYVC&L_gb+V)2&U0<#79Sb+3Lf8WScYO=68N-f[0_N^U2;_
W:R:,45e&WWZKN[KaHOX5e1R.+X@/[5E2EB0O\(##P\F(I^JO<AG+QK4/QNKe/;g
bKUMK=<;^S?0XI77A6?C#?b6S&>+NIN[QX\)5^#@c=Yb.6N@P9VA2XM7bLZ0fEGb
a[7&0LGQ]d&Lf&OgLPb(BS:Y=Ja,>c-)b^9U@Wd)eWXaX-TA@)#MAE20LO:EA+IH
?f=O5I+TO_2CX)-8IU2>g]_0NT7[B_DaMcKQ3]QAA>Y<Zd&7Q@[FCe2JY,H1D@<B
O\;KY6L7Fc7gOHGLTZ//:>bWEQO/W>FMg@(E6UE36b(d:]e)a#c/[dS9U<8Q0GOK
,6DQ=+.<Y49>JQ8Fg;=<Y_E;R)W[SD6#PDF^MbN.<2S\\U?+9H1(L-IF@AT^7-=,
dc^34FFX5[^\>\Bbe4A3UT2YUBB+/4WX>C/XF?V/IS:2M94:gAX,F[M=LfQ3QQe^
1&d,SCI-2(0IG<-=/gXM;f.A>SWa<(,/:#W.Z8ZP1Vg/dU].38W_0XJZMMa##E0\
H>/JKMbF_f4>P.)R\@:&<RD/^9U3@1BdTK77REfU,aN89.?+T25EAX3deJ.D>;DQ
BZaaA3VFLGg6EYF0d/</YfT/(#MW3K@+e4.R3VE\_+^g)8ZN?0:5?F@g)@OS)86V
+cR[/[9MB^/R,gX7OW,1=D7XR#K4?SKJJcc>O@G3f_TUJ;U)Sca+[Z[K^K\Td-f<
agQ@4/YSF)7_Q5FM[_VU9,GVZ,^J\,VOBK/b@]A-H.?^7\QJ.5c)((96>J]\6R\(
Y0f,fI6N75_W#(9>;EQA)]WS..QO_-#(CV+6M>><;O-Vb6UA_ZU4cB@N>b..Z8YL
0d)#<eTcQ?4A,VJcJL=[[.E,c6-89]bYd-H6Ba\f7FWZH@LVR@32M[MVHZ3bN,^&
EJZKTCUM6OMW,X4JV;?Z&J8MePd(P:VT?7\M+A[EKMf1R][,?SA=GI5U&KO,N3FX
bc,(/C0fD.4f0?F<IPfY4QPG(FC7f43G#SLI<\8M?5/=/71=RE5)-e@3:gV7\.b/
6?d66W#,;E9e2R5WRTGZPIg_\aHE5,\FZFf0:HF-a^VP0E;fB-R:CeYV6gf+\B)G
9A,1:>H=79[3K-X:+gaC(3=0bF-Y)]f>c&2]F?0G85Z/F08\#295g&H(5M@?BA;[
3Yd\K2fD[]H4;LKDKOQ0dLT]8Hg<e8=3&EID0dW98;9[d7c:&IdTX-MRL2@eQ)RI
EXZCd,_30HT2XLg#_N&bP/bd&]ZG1U3.a4PO7UO-gb08OAP84\eC]d.aPa^cSN#1
Ne-J<&bK.,-0L\@\C#4916@Y[;Q7gS0W4@H&-SB#M)Y-QQ53ZC9X3;8LJ/1G\K[L
QC=EEa3c(5+&.2d+HW?#[41gA0L;gV<@&e9,<K1^.dPVPESI(fd\KI8Y,7#D,F2b
22Q(f>+2/N)WB^_IFY[?^=5CUD\GW8;R.AIJC#CH/ZgNAY?35^MNU,^;/B^Y;F5G
2aV54E)?)/O.eG@AS1SU-D#@0HD:59TI0HDBY.^?MH8)+/V-E]I9IK3V0YGH1:@,
a@7X05&dHg]Ue(OI_28D3[-T)/]#Z&24bd(TN>1L;,^,IB-4O[G;=WJ=Y0I(,U>M
B)^(XfD__UFD7:G==B98g2\^7/3[1,,VXfcK)e)g1)0T-2ZY]EB]E8CPb>9PI5Y@
N(8.07EY3\5M6DURFJAONASf]Q1Y&_+SOaXIaf]9SM[-2&Y,f]fce5,@]c0T?JGZ
Z3E,Q-^2QZIJ,1FQR\KRKXY\Sc.U#E8aXJ01^NeOC22@<Hf7^\?^9+>g0^D>K)DI
Z34/aLbeMG0JZ.^GKg)>X(0^?4.^I\Vc2dOdP0CCARQT9/W.CODJ[>Q6PT)gY/L]
/[;-b0YVNP6Bb_cH64V^;KHZO55f@.7WZEX_RfG-?6dVVH.\UJH>-QY?e3AR/\#\
e?>E8?=S3Q/;M>9&Q2V]c##,,U+2D0\SHUE[K:YUI9&L6<\2DW0:faRZNL<SH:FF
,+ALYZPY^GFe/FO0+bI[T#I2GP:6?Ja#cN+-V/;\TIde/c3@P&>1]<Q7>bKC3[2U
6EJF4daJ_LTO_0+-#F^=4<UdQY[KG\M<V4,ASG61g5U0)M-7JK@;^X05?&=?W2:G
O&fTN1&<4#;<B9c(DVV)JR@A&Z56;JU.HJ)^>:E4)]LO#Ef\;J?V)e6;2([fAPU;
3cW#CK<ZNT5_YL,D<1bN#YHW3KNB>(T00=(g@(R(GaW=K:dggEU.fM>N^MDP5fSS
EL4,@SAH(GF0/&KMK6<>1H0^d\#++UJaX)RKP(f11C(<;dId6B08HN#AeEZX\U^-
dcT+5I:VGEcNZ4^b<HFRC=NE;3Z-U#BMQf7_XLDaIJ_,^,TO>,cW^N3:L1G3Y227
6IEgUWI9>?8+PcgZXUXXe.aT=@3fY59K>17P5TN276W=P<bUDBL\0aWJZAI2)\\5
a=.:_42OD9IS_RPAD+45YbKe).1Ca8RL5>NX7D.J&Ja-UB1F8HWY^JD8c2)Z+?7f
0865O+/,2L&LXLac;9g#d1+WaS5EUL>4,F01Q4FbaB,(A6H;TDT<XA-FSC]Y-dEg
9QT2Q,H5.\>Z0Wg?aK#CH,?E#XZ:a6FI1Y:E\]gJ6S8H[c)XPF5P(;8&0JJM,:76
,-9Qd,:/UF\>WJd)dJI-L7VUW&PG1@e6b?f-9&NHQ9WPeA]NM.8gI,1e@0]HHfaf
10b9+88[-J_<:[LfL7I@8fd2Y=:57MJY+ZG<.(Y=0Ve4[4[-Jdg?O@)Q(DVec^#M
=/UBERLa8(@b.)-:SQ(Ma)(&WM3CE<.C];JAT(;bJ<fQGP5H8a,8(84Y3>MTP9L4
\\_@N,a4=#0#=6&.8Q&>(Z9c;VR[\SP4:]_6R3]R:^=We)(1J9=fM8F^dSWKY+Ie
-Ac;d_VZ>PcM=2_#QM&\39I:YJE0S.&9)KJ3CRL]=;2X9NS\8V.SGDM1D5J<.H,@
3,6J)M[MbLD,GG\)Ib8HXV&3Q51@?]@\/96\F?.dT_06E\M>(gM7\T,+CD&-+f1Z
b:5N:-IE;^AO5<I6c,dFV3Tb+?RL-4./P.C/\?PU<EP\]Z&>+Ad+Z+5,bVd,XOQY
IfI&#NZI>^a&.^V2,>ZZ0>E)+bT#CF35MD.7]5I/fAK-g?e3QMQ@E&cT9HA.@BSX
46><bHB8)JTX[efX;UKW.G:LTML=]=D1&JE=D^1H2#L:fRKXE)[)=ZU7=f:d-\(#
P(1(]e?D?RgWHI/5MW[H]YD)D;b1)E7J:T4GZY)/=^d1#;\ReXXRY\2Ha]GZ1K=_
8@11RU>I3K+J6Qcd<KPSV#7I?.W2^K2@K5SNJMf<(J#ga1Q?43VLa;Cb/D7\-<fF
a9G,&])-A=.@#eZ=DJ7NRP4C]]ag_>C?0>d85\,@U#5TO9QV7M+PGK+cT50SF9MY
b[J^KWgEDfPA_VZP>_S_G;4H,Kgc&G<;-R[2[K1^#Y_?a#FQA9RZHP\_cff9=eI8
SELfeg&.J]PUE:Z1ba=,#@W?MUYG16MK>&Tg;eIGM-VFP/@;VP-#RE;=<DSM4KLT
.aJYfg:(?U-0&PbEgUCFe+Y@:Sg2XTI6/RPX&EO-SLOX/KQAVDTUYe6Q]Qe\4;N/
5L1=O4[;2ITRGI1PA7;[7PVZ+0>7DVNgA4\3;GScU#Y_5UbCMWPF^]aQ.9V._L-;
>W/LO0;b2QN>(0)[)>>CMAK.LI7\_,#=Z\0Uc)HB(aDC4AYBPR-269MJbGW51[b_
CB+gf:bOfQ7^/c]ICca;/f068A(>^-:^&dF&9R3[g_WB7d)UC;BX;fT?a2U9WD/<
=W[K.QXT@U,T:CV1>_?FQNFXFTBdW8Me-:FN+24\Y[2N+K=]/d3&TRW&D_6c<Q#<
>cZ^8a,gL==cV.adMcaa>8?EVM?U2;ITG&@1?):\gVR.5cGcW<0:^TGC[LW-/OaO
]G_O3_Q8;fN4<[)C7T;K#L8ZB]Q<_Ka=<-DTSN5P,V:0EDAIQ#017&cSJE?S?a.f
&?KA4XO-Z,gLNJI)Fc34a&VJ/8R3EW3G74+?-F[bLY&)W/<;ObeU#GB8dR7E+1dg
(/SIEfa\^J</9Y]2a2A5BG@Oe07/,LbK.O@MA>B^Z)==8YBFLTE5Q_Xa5#6@gW7P
+7\3@W1eM00=Z8HIZTY.<SS[db?c_MWCcOA8UC)]f<a)DQZS/4AB0g2Og>Q_SY[b
AEOIeH_6AW8c2&IAEF,PUG]PVV:(6dW@=<F;g?I5@8&gR;BQL9\/^^+SAY)a7]?O
L0+YZCC5#9S3^a_88Cg#-J1C5PW)/LM\8)N=TF168&-J32JAL5\7WYc[6/6#_7eP
O1/7VaQ+8_-9RW^7BU,B5.,@_;1BH\^KZD1PWSS#\_HAD<S_7EU2Y(bXJTc=+6A0
V7XB.RES+=.7B=GCf1)]5?UfgcM,<J?>5-ZSgD:a54>3\T?f;Z_91@\(1Rb(&U#0
;f=:YS40>+2/^Q&Ng0f@:7VF?@gdgD4B.2#Q6P72[3Z2DV4G,9-+AD3DCV)+=12T
DP]CUgJ?DW4^&@1c\+N&.\W3e004#ag#;NME5E<#^cZ-657F01#X8)\Ve8TZPR8)
Z/#eN7LW0O^b&D[/,QND@M8Y9R7_fI7@:]e7Y36SOEB^UZd1R=OI)5#6F?Yb09V4
>R)dbRGQ4UYKc/T7VA/fUQ00DVZ2-<2-8C9Y.]WTV+[Ra4+?:<TdU?:(,4URCc<N
a<Ne1@YSFd.#DG0#8:QBI=(7O+)XPWVL5NDAJM.E4.)ZED&08RO0b;gFD5\@+:86
OXQ&(cR]8\7UZfgaZH\#M-Ec6RffK=(2B;[RGH,)@UPR]5f&7H;.(QeZT14eN_TZ
=U)JeBd)CA:8#W_#bOP0]SRVQ#N-?)LX2X6QV.]SH/gHD@aE&^_?e5Z&e>1M[TdW
N=>5G4F0dF+M]LF_UPO,4f/\IOWAY14:L4[HKdRcBXSX9B2C/Q3c.<5g^D21JV^?
.Mec&)@a?_20.:cPcRcZ7@bV[\4g0QTM4B3\eRV>5FcgK#PDg41K=F7faF.KE<5W
A-(LT&4C;ELIN&c?:X-YBI:B6NWTSWYP-?,Y_fZNQ8/D.IOU)QL1/HDR<T24;CNW
2VcWaH)HL1d?7a=HS,J+NFfR4>,R_CF_RV@;&aLKIM_Z<N^aFK,JB)KN40<DRF-L
,+(S,V,JPI_=#OO(73H60K:PK?>f^(&R098f#/4C:=303\0d\^=aYL4dUQ\HeHc]
>TDN]BG+[#G0IHfOe>4G2J/;ca1-C;U#&]O;W>7@9/3^96fa&C\O:1dY=]>;)M/W
[_Y.QUI^KCJ-aXC#J-X?Bb+MbbYeK,5\0]@Z]IWcN]HAFHC=6>B^bMJcf>:UG(<N
4.XF6<[Q-23.PJY9cLQ71P,X&a>ZQ]NLKP:+KFE9Z]c9AF]Bf5-TJM/XXW?T;F)W
(Z3-9R3L-E+29_LO,U@dG=;6gUE_C4X9J/D2[QN3-[#<@)TcaWYPS7NM]dDEB@QL
BI<VA^4#]9Bda[]Gb)@[AFf6_EfA=0XD;FgU=d.XM9-W;aR\IAFe1CG:.PY=(9YV
BA49M+OL[7(F=Y(V8;\M1&c#@V<Q3PKM)Y=[=M\e\a?OcV\TEB^,gC0P&\)@):cK
VADDIB[AN8Z#TXL4\NXB:T\);;2aYIH1EW,RJR?:==<gg]1d+0JA?SCc:1[S(^^?
\\F<>d5D_?48F>YX18Q52LJTETPcMc,fAdW)PMGBT4)S?6USR9C6;NaGLQ.9(YGY
WLYLGD8).FTF;#cf/^QUL//+[C,,KFV/?P4G,+=>d]Hf@5.OI71EJ#c@GVN&9<UX
BPXY,TR&_ffC;9;aJ(A3B9_YZ.gT[7VR:X8PC<TB1UKc(ECcT0Z^E5,)5/LL2W_+
2X+HM&eZLPSc/K2S-JP.c-2WXL&K-?K/IF6;89EaaJ]IECVC.Q:;g=aCOaCM371I
-J//fOFUeH9AB3bVBgZN1ZLRaQR;I[I+eNV(M&#2C/c0NN6gc9M/@DTK1b3RZF-?
X/.Q19<^-G8/L4,;8=[+/PTaKTKMbce5We>)=<FWFO[g<c;c,I2-X;6I,FMdP,5/
#9VZ9</fU>_@>Ka(F=@_^5fK@&T^:/,P)?;P?CMeP1ONKO]#7J&/4)NU>&(8Z9G#
YW:fP6R,C[ZX(I,BaGX0JP2#Zbb)_=5=g3M(TJRJMBE2;DL0U=IE4J2,>>SSHZVX
;PbcAdcG2J\7N;Z8G[0;bB.aLF6@M4G]FXCRZ:^CQ8-0D6O0,LW77.f8<=#P?3Mg
88:P^0\:[=G4W42ZP/=e7c3T:[a3PO()_FH&F1-C9;9b;U6BWG2^_)gN192M[?II
NKXDL+)PQ7^=>7>QUE?,f+Rb:04-ddE21EbJBWLG51NX5;41#T:QZ;,M=BL/;?\Z
J#@8N3=MUQ,[Od2M?HA)Q5JZT8F0=+R2+eN4[2CVR_&?>J.-Q3?_2Rd:X@C/4OA0
&<[F2P1QY@&6(f^,Hd&EA)]EHMT9UI:[KK/Af_g7<4=7e-Td)Je[5M@IT&?F[?g[
@XNag]H]gTZO[?TdP.[&R)/<A@cXJJKID/fRN,cK[DG&JY5Q;D\G151KGL8.b[J:
9,IG\T]Cgg5g?eR<8/(Ff-;PONSMA#3QF0E,&A,<SK##9eO;Kg9V@F6RBPP3400:
:c[Lg)#HYV;YJ.IZa3^Z(FDZ>;BPA=dOf;/JN5?#OK\E)BD>Y-FaVbcNIgHB:?YU
3bR+DZ;D\2+CT]R/,9D7MWW=c4I<?UZN0,2=[aKN#g2J9TU;@5&Y<#Zed(aNV)MQ
SS96(90YbXNbUUb9MTc7f90^=.NR6#2LdZR0#4G.OTeEFbU6QCKFZfeSg3^&O6&:
B7NIS[66JMO64gALGLTeO=C^8MbQ\c&Ec-.MJI[]>6f@1I&-_[4LM,AC@;gYJ6UY
+SL-4)>J+?C1YbRIJ:AO1_[=WIF>7=c/Gd3/W+B<(d5CP=fK3dHL(_]RM?;#1N;c
I[e9>U6;cCRS,K_J+fFcGAfS:FJA_b\6LZE5a-Ca_4-5R&1OEWLF/]_C+C2W1/BH
<=Dg/A/P=CP][)J;9](O9?@#S8P<7\cJ9Y[&K\_/8Fa/&JCN54Qe7N5&FL>K7(aR
X3>dWZ9]#_GO&_C3XEU7W/<Mb:>QNQ[IbKWL5]PMUD(J+22KB1)J:#/5gZc1M;gd
9HI,WdNBJ(29:D6fTT&2B>g85&]LHAMTd=c&K+EU=L9?<.:2#J.X]GWdRfF2-[4U
/.[)WbEX1fBa+M+VVYRG&5=g2=]Q@/OP/AQEQdd8X^W^3ZRe8[I0Y)5]KPe[B9>#
10B;6N3L4QA<\/KS#&E)GP0\E@0X2S,MW40A8d=,J-Cab,EV=V<\E.C3#HEBUR.6
/2U[^B67BE3fX6TUP),8&#S^;/FE\)]V-.e89dABOZc-HQaZe.?Cg&HP0_Vg(+LF
Z_,7Sa0[#YI:Q7UQ^:Ec25=M98Q_,QM1Q[XbFCCROcR+H/_0L_]:0:8?\_A#fd-L
fFY<W-[FH?G^2C5#+[4)X0;^&^[f\:Kfa-AH?cFSPFa5S_4X4DG5O=2\;e/\F,NG
efObU6)8/a+c&856A:G410;Uf?2B:I7@b)Z023?PG>S?@c_94,W_^#e)UD9W[6>)
/;ED3Y<)H&/?]fP0;c^))D3(<fgI/Le?e;XZW(I)F>ZMMBS@N/9d(D#K[#B,B]R]
R2&D]#6fT/M@45_X[)c07gX_4;;\e@Pbge--L/WHS,SLDCb-/ORa>Y1;7I:[M_=C
CZ[,2O@L&Wa#/NUf<7/Jf]R^L4A]VT/#a\@JI9B05[BMCU]Z=6T<3SP1-.fZ+?=V
]R>S.M@;Y,PWX[Jc]F1+[KU3.YSQP<CI:.RM#>>=YB.//:J-aBQF<,#Z_#SNQDd;
fG[F111URTgW:DXMIJ/7ZG.VM\P21e<8,A+G+:98>+]AdES4THXcA.L#BcB[-V&X
3CE@:,ggeM]AT5)))<_+R9XbAVY-29eRdI)&0PB08ZD,@_=79afa?.dc,AQE?2Ef
0>/V,6@g+,-W&)H#XF.bQU:P;bM7>]dHN(VHB7?@4#:O+;YGQV9@^gBME,O:-=Z_
93<90P2QSOL#X[&5\4TM\I77>:O4>d?,Bb,Z3[4AaJW/J=X0LV_/W?DLI&LRIPW:
UH-R30@gXD@1):]Qb+WJM_<E>C9UEORH,/A)U^aaV_#A^D)5SH/4e2[1>LED9_>@
_<J)/)VRecE2=GYM+>WC8g&>I?(LH/Y>JfTBP&DdcFBSCJ=aFAS+HL&4.a[a7/>T
CUg4[f:;3Da,8Td/J(>OND)Cf9+L[A6Fad2Y(-9eM\+bD;:[9e\?JYHPIdS1[:(X
HTYE\\7/9<\XbN700ME;X0:9P0G7=K+[F3P,/a<a7_][bW]]][_(>)(6/C2V=)QC
H/F]S_Y5,GCcE>LQWL_\F)GA#L>-?LJ3EeK;Z/[V\VcV?IS4.-J>ED@cQ9,FL6<.
Q^9/29GE/RHZc7)3<,5_(N1;TGF+AcE<;^)(d\b>K3K0f#U@B&J;D=Va)P69XE/&
>JA4]U9E5V7H+3f6HQWQe6aV;+HKfU#HDIce^5\I65>b_1K0/0QQ,(D8R^T7R>DO
I8]YS,Ha(+MaF=?QV-KMNV8d;.7-Ld_>6R0gBHE#BLX-[#ENDf[=;c44Q>XYOJ?_
2_2+UBa1N.U\[gWTHb,5VQ+W\KJHQ=d:=QL#\T_aNG^+CNMLGcLSM6SB&NY_?GBS
26HXUP(].TRT?dbLPZK\a0(^]a5cEfNd74AI(GbS/bL?],Mg+[K>US48;8#.CO:)
0XD@H-^#M_E[#E[2<Pb@8];\()4f-<Z?XMA61+VJ4G]8dEda=H2&MfP:SR]0L<.)
3M[edUQB:#H\RF72:6b3gT)5V_aYbSL<,,8bHC=a)I9YNa83&Q1CcE56df?5<9JE
^+^b;H]GC:F[e_N,X>NI;-K-?)>fZNA7VUdI]]bHY0?7ScId2V:c^E.#__J7TF\W
@^1BG(1gA1-V;PZfEYDZ0<3Qc7fDT2_c<g3MV[]_dVcgBgR:79;;7M#bc7bT9F\D
OB^XD2fdY[DUA^a/>,ZAb3W:AIU8b9<RDfS-f9fb,HE):<dcB@W9]d\)PI1-45PD
.1LN0?fWM]U/4KZ8U5MIg&KE8>Z@R>G)#_YRg[X1PdJ];I0gT:<\^MY&eKFSCa//
_90YO98^^=gZF)W>4@]HA^S4-;LWc2R\6][OXF94B#g309-/AZA]YX7IF;WM>TAG
WIM&R4MMN.^gQd^ARWMGD]M8R0UTU>.03^2VX\)HM&3VLN:VSg5-]X:d5Oba^^X[
MgOG9IM3^\D:08P@5L\@6]1@@YaH2[H@4fG7:WFIIDfCWff3UR<15ZLIQe@E?QT#
WU+,b?Y:f=K/N(IR:?Y?768FP99S+2d=)57aU7<4^c4;,6e[BQ?.4<K>+/Q>PT,D
1,Y7QJ8W)Z)<I&\#LAVI?eYR8^O8]IX#d+[.3T&G.H^V3Xc>)AB32a.K89W3(_,L
f(/=#J#OD^0aQ+=g7<ZN3:T];J6A&=K@VZQP?81LDQHG0EN-B(13Ibg6Uac3O)+W
1M-KHd?APB=52U_H6[U9V+//\R=bc0YD&QUU)Mf91::GF8X3MO;dRNG3e_#U57EV
@QG<>D(+ZaTF=(Ac=7P_L6?\_/4a&Yd(@#B93H5c?XKdSC39P07d<Y=0HcJ)\Zf_
Q,\J8@IQJd0(_#/))cB+_f[B_:WLbQQdV9)[ZaU/5f@gM8:3X[I<TW&Na[LDOP.<
CX,C]-+HG]H=,2EPT?\A(4NHOaBfO+8;)?:1=e/cYLW6Hd5K#[H])gVD@@[</?^=
JNa3,bAC^Ja<^gTL5c8[11<5T&;\CHI)g@.EJ<O<O=MS6X&Af2.Q[Oa]_(J_P27O
8V+L9JNPX01eIdW#&SNNS&)E79f3AT:M4QF-W^MI]aP4(=_Z<)R7<J[fI6BM0V=I
.MfQ6/[7Q8_RKL6XI1Ea8DJ&(:E:,=#f;7))d<?FI?7-RIJ0@J&V81cF6>K\^4+O
[@OG0P\_0F5Zc15_HJXfHXK#Mb\1CU7SD/gOVS+H28UPa\[>6V:F&I[Y3E?.?H3.
1CUY?fDAc:ddb1Cg[g64@QVXC7WG&5-bF^b=dG[WV^.R0<1^ZYZe(H?8TbgGa6@0
8872-cfV@_HHV?R7DLLT6dT(7OS@9L\&Y(J&4+9=D=E:D7FHU]caQ1-0@4)?1T_D
f1.1cbF),gaf]d+IeN,SG@Ue+R]F&fP8XPR^(8T.aZN(J(cfaO=@[38J0:@QI,4=
cV19A+>.D[=QB7a>]C\[BS9^Y21Ua/.K/LT-CH-^Af6:#L+S+]^d-^_IDI0J-A=.
NdF&(QU?62C&\]Z&9d@@FAgQ-aUR6G\+?LfPK5-_,1e#?(e3Z?\@G6.LQ7K\NJ_5
,9XZ6G-I(01_ZR@g]T.4;Y+1FQ_-R)CHRK7<1\5\]/MZSG2SZT;2,)e@B[D\YBBW
aZC1;,7@1T4.QYaVS60GGGa[[-KPQQGI08[NPFUH1ga,G_A0#3e@GMAYZ]A7e9D=
EV:G7DU3_NEI[5(.H>OPD^O?UbA.><HLIOQYJc)LM#HQYe_LHBW>c=-6dfDcM@&A
C#e4RL.aGGX:3S(#9]]BT<0&L?WX<MZVRg,?KOIQg;J-R2O@T1g\gOVb-ZUWCG+g
1L+9f04b\5bb1dIMO6X3X,c;<U.N&475f+KCM/7]NL&e+>#GXUUKSgbA#0N[a+I7
RLATc&8Z6BFZHY+aYT[eNFQ&S]&O6f\@\:83B+E=U=O>7)YRF<)WJ7DP-1@SBOP1
b:HE=/e:4MT:cW\[;>:3/SJ_I@T+)C6EK2\fEQC/:V(L/S3#)55^E-C\H<YA#:Y;
9-_[80D)L-D5NbdR4-)eVJ9NF^T[:(DTRg6UP\-4O/AJGT,OP>bP]cV[MY^L6L:M
YY2\T</A9Gac#@,J:Q9Zf)1U2,&QJ>?.FB4Vce[(1(Y@\@Mcf<#9L[/fM\ZL)I#N
a[XP73;F2Z?.7Y3=@M@Z:I]H6MKd)9MWKZ&[L#JV9^=egBDM6@TOFgF,N7^G.PFZ
c:6NY_B[DZ<MXaa5Y6)L7WSc79=fB5MW6K8Z0C8@(H^GaM-BN3MgKMdH>Gg0RL20
A;/FH&L75S6<&Za0OF+TgfHfX07A7,[I3=A(_+=LZQ>67E^+(R.a-^RFK3ZHBQ45
G2H6K9f.(/VK_#6bOdM\IO1ZP=CRZ+Rg+Y60@4X)&D4UbX?f]f+#A=^K[d9cU29<
VCC_\HB7[7]JN-7RI18[^Z)1?E+g.?XOBZ<(6=Md_GcLZ9L<O[O+0a\-(@YJ=@cJ
ALE.2/D\9QT\3S6dfd?=aBea9gR&]eg@\G\55:+OXQ,/R+cS>cYNIY,RQLZ@?.?L
LHT=eE#J[T3+CL2>>.?>5Z]&Bd-M9FZBXaE#[bHO,3Q_a2=J_cY(/XGRfF\XO(1M
a(L0fM7DL:Ng9M;JgZ=,d)I^6?@3&#YY;-O.-RIf0O4Q^1S-P0,.^eAB))Y/CCB2
]79,f>:QM;I\Wf#?T1T/c+4NfR<GC#(f.5ECdU&OVT^#K>)06cXZ-Ka7;QQHG[e7
RaaKG/DWd^I9#P/<B>:M:T-EL?K@E[GFN6I\A=P]\+22=UQ8+B<9FaWO/Y+_3SR/
W+N0[Y3ag[dXAD_1LY720^F7XB83.VZ0&O#2V+d))BLOe7[FVV)),#Z?J#M:IT9=
(\MZe[d=E#Q/H=6[2:L/U+eA)M;/U]f4gQ@IG0eH>]+5N=f^TJFX5,&Z_UIO1C<V
.<[LL2_\bb1DP@>9aKeC-:3b>,PKY\5Y3^\-9&Z6Z(bAGf<1fNF_?-7Y(C-_;D4Y
6aCNX;\(K;3_E637cb&(d_NdHI7a-FF2;1fBdPC7<,TL)WVJ5SD>J/IM2T^]Wc\P
)E<1B.1SBA.8=NA\TPgR>f8:acgU=L1C0@W.@9UgY3LfCI&X:+dg#6[8VN&VZ/]d
Ea_=g;&?fWZ#GK2Bf;f?Q59O1-&Hb)CA2>PK9>VCWF1Re.EdNXFI\bK>_;a62>3=
2ON49C&0DYdH5/7d--fPS.f.f?EU4cM#G:F604Qg]616H8M?B&72&QcN2[VFAKZA
CFI:\3M[g6[88fKN7L8[N-:,IXb4IDLM_d:SOJ:@ZQ(#N(#3\;/2VRL\6=V.JDdO
SD^_5T+Ud69>HN3&:?)&1V6)9MS7/C]HJMR=?Xcc,+3JGSf+B?36GZMbA7COZ\\L
.e(EXMMM#VIU#8XdNc]5>DE)N5B_I^6ab,[OAZ<Z52NH)X=cQ4K1R>=9CS0IedM6
A+c7/)Sd0@)-3We0]BQ0McH;)N(33YLLcMUMA)<GT+B<HO178NR_Y:;QMTT/D1^=
Of9O3U_e)+<BZWPPS(Q@+:64C27cf/XG2V0U)UJO@Qf+d28X?)D&J3/S):M;+D/3
IMEcMN:e[T5<(^76<@JJ@2)U@&-bO\17-97:OW282)aG7\1ZAPU^caGSH2&-=D]M
G,9+PTYGJ>^K?e[WQdIF^(c1LKYK;cF]#+g).:AeDE1/4e3.;3UDTT^S6eP(P#=C
>+eIV;PI(#<,71e,JRBO[4(?fREUS)bgbVTT=1JaOdg_KVJaNU8H]e/+KH)BT)/W
:g8^M/CcG((D1d=T805ae]^S7+-\=1eKQ6OC)+[D/9E3H//^.3/3QMON(R\U?H,_
/7geW(^3>J=DgW-42cg-BOWbE=b\JC2FASB5I4W)/F;(D=[^\GBd=]?W-5W^V@ME
+e;I96@W>/8^1TcOSa2O9H;VIGb_bfUKXa2Be=62;[R4a/20a,#L8QU/Y7GJDJ1B
11:5e^5/dL^,5^7.>^@>X@a[b9XcCDP\7X,;EL-<HT[[8F67\0c>.W@#R(&?+b?;
=.A83J^S.&GCJ+(^<+?C<,d,4.TV8ZV,)=ODR\4>G?KV[JRA4e4YHZ(EKO6g-+=A
S=#;?V6aYNJgX)41)2(JL>AF8O5&8DN_8GQ[().7DeLNJ92+02gJ1;#JL9[/A=N[
NNZe&Ab/8GPC5Z0P3_XO_,>I5QXTRIV8?AH2L;DVP<0L?>?a8\<eTZbJ1Y>A0a6=
a8bGISde0H.@57&VJ7=bKa(Sfc>;Y8=:?(]R0__F5BBABS4<;R(bPc&KOW/cZUEd
1+N,;cH^S]2I;a.BeMKA9cB:0JGH2)(P@131M\BfQ,5R8<I1Kf,2#>_IbH[IB39A
5,gN5d(Bbge9LR6S6<V)FHZUZ-\OdHU1a1PG#:,WT;G5Rd^F5/_1VH:PL[4K@Q^#
KFP\(3^.&))=Rc9Ld^&2L??]7Z=ebA]\\41=TC_C6-<d\G9S1J(VbFN4>)N[G?G\
/#V[7[&N8F/JFE>Adg(LSb)@6RQX5W+_DUYW(cLSSa@]YTg>YN?6D2<dIIMbH(5)
P],-Me,U@CT]F-?bc/?&=YHb6Y&0W3T>VI<.a3<+G0D6.1:)gJe[G=00<#L(C3-@
;W.UHbNM7,+_K/,?[XKYN,M+7L[3@BgT+Ke<DU;S#:9&3_#&H]d-gC]S0Y0#(U<,
\Mcb5g5#@>-a,I\T38\HEA9Kd9,=,H_1)_Z9EE2CYBRCFOR58ZP#G+<B&d4M:3Vg
f//&NJGH;-\.X=O.2<Nb:7=BW,OYX]HZX]7&S/5(G.a2F7gB#Y0gQI)-XE&#Z@6)
H7W2&Q3f?P1.1C?HFS#)#bU(\HF,@N#ZZ#TKLTI_@WG/>\82P==.89(,c22\bfb<
U6d=:61UDL4PM9E&@K&P]?A(K<6gN8:\<D#.H:>?c4;WLL(8e0dILRA5-aV?R^)J
7^?6YEI\;A.Q?P0Y;;ZCf5LR)BJV)NBFJ/B;-CP].<4dbX#MNb,[H2dY2C7eJ,OT
G0K)8((G;?JU/URMBPgf?5LgB^HYQ=N>>f14f:)_SF()R0@)JI[a4NKF,DVcR2eS
T@f4E:(d_[RWU=D(O9cc&(800L&:=/G?aH3_>ffT(\&G:CT5,R3.K:76?;8^[V1H
WAZ]SI2_KCNJgFC5GS8-g+^c=eT.Q@P:7V0X+?.FQ;Y<I-.aQ8g-7d0,U\I^7=.e
De&@gS9]9&cU#D\eQ1WTX53T_X-1M;J-c69=B&A80\VaQgVZeC(GK3L84F.1-E]Y
-=gG@,d,C?G4GLA[L/Zg9fLd8,_>A#IVT/@)/M\dDIX9)72\M,cLK\LH]E]c&M(+
VTCCJ>=PdAR]?gaO+X?bNV0;2?[7cc?R_6WLS(9,ReL0I(H-B+9aNb5\I8gMXQaE
4G@G9O+LU+;-BYH7V:DdSbHF<aaXPKL811,V(JCMC(T>#6QZ;.-,=N.e1YG@+R&3
QW35]e6;;F-fA=MOM^K7)F.c@2T=<(Fb?WRW)aJ>IS\:Y\-)#Ub2:,^AU[@BV[A5
=+R\B=>^ePQKfKaNXBaY#5;c7AXaT?<V7SaeXGS?#;dK)Cc8d=Xe^XB@f.-H8D0J
X4W/].S^&A+@L7_6-(QN,J^FGOL=H8,,-/YIZ],+#XX&L4+I6>Ra9AS73cBaBbg;
@FTd@e2W;<Y]82=IPbZgHX.=JIQ1=MJ33]XfG8f,ZKQKRXEUBIHCa138NZLYDY:V
7fM+K,9LYYUC_(dAAJN?9VFT+#[EbB(a4E0<Va\YWV@+EBF;S4YbT@)^)0TUg+H4
5g6?M]=6fd?8F4N4Z88#AUafg(B>4L)26GW>F9aF=)b?NS.7@UQB5BKKa?SG2_aQ
_,F6:.7(Z++;6ZOY,4:BZCFD=D^@4PUBMRf51P81UY\LOH##>@N)<9&,?R#\\C7Q
3.G5:g52bJ2+#eXb[b-CUJ5]ecXQZGT#]_eCHW5.3#IA.g1d_P=6I#3ZfeK-879X
7N.5]B+cKgJ?PZUSIcH0+U6<6?g\U,TT_YV/RELK#2:cWG8A@OKP/OP?HB42BcUH
8UO;X^@0GKP^D:[Q0-PXMfUB4Z(MP47ScYM\e;XW3\O5T_O@[/g?U=.\@VAO57</
VYM>fAOC3=MCG,:3F>M/&R;eEb3deM:,G7Fa)NX;Yg@Q#C8EdVM#dB](\6S7^Y=M
+C>=R1P71ZX6/g=@4;HZW6/QbIFg=?WdWIM_AO\8GAR<0=\,LcOJV0LR()87(51G
LRF6V/a2Tb1QK@60DKTQNQ8S?gPQ@=BC^5I)a14fCDFCdH.gLR6c9HIfKLNIW603
E>2[CgGET>NQ0$
`endprotected

  `endif // GUARD_SVT_AXI_TRANSACTION_SV
