
`ifndef GUARD_SVT_AXI_MASTER_AGENT_CMD_SV
`define GUARD_SVT_AXI_MASTER_AGENT_CMD_SV

`protected
aZ4UYS;E3KXD7W0).09;6bYB/_V6-[eAEFUZ-c[;c(,F_+G:#SFf3)_>H)gP4=_B
P^Q-:fLceATH8_?9;\A]0c,]\<^N@L0:bP-)g(:;3W3[;V[(_5GNTJJYeeEW+LPJ
HB&P[?6JY+-4C(Q1-40<WC5L.>S(I@4:FUARHL[FKSUG4WRS19OH5KXaW<C#Y[d(
/8:?/H9bf99NKUQF;FE-5(]]cd+\g_[VKgdCbI-]ID2(&E4/Eb/WQaa0FI2),T7/
K4=P69.fM2Qg7&WbA:X:gI6S<0XQXb;5\L.6c+:,JU3/DdA2=I(#SA@)8UM6=?Sb
T#;NbF]C7F/_.&a+T\f\X,)?,dAZ=c5[g9bB37f0(=3)g?f_XLZbg+.(>HaPV]4P
T171=,(=?,EfaS&G:#d=\8D4+?A5G2f/f,W06dP=AE[>]c\gY=RcYA5K)gNc_VBL
Ja\g\;]OML5;P_L\D#/^5eJWK87):?OOZXN<IUgPQYI/5UBaC<4Nf2,\(O6PSL]K
8R]GQ-#+7&I/3)6\7L8/[0IB/>8RF^L+L479>7eQ]Mbe0gSaW>Ad5YbX)]?XOGeS
^8<\[Q[29>[\H124W2F,Gb01/fBR9W8^H0;<V6(@_(36P>RQg\+Jd^gR8UFPP3aO
FN)(.Vb9=SP.H2>I:FQV55Q-/?J-3L(E[ZYF@HW,4g,D>2,,9(AHD@]LCF;Z7TR\
4<FN1d4XFcd]N:UV-N?Q[?9E9L#7Wg4E#M?,>@TWQSM(YJ-I6\AGR.>b#>-ddEJ,
;-dXUf+2[[GGVL8G,)?Y&>8(^1KcB_.@H;^;6a&<B5]58Y#27ZY@&PVHR220b\V)
V\c78NJJS).O>-Z.UQ/JgZY6]ZXX-EfX]_E\SNZ9GYFI]3G6/9HAT:IFY-JK->f@
@;E-3@:\5[P&IL@]-M?@:?f/6QC->):4+,(RA93fN4#<=CDU>1,K-J;?LZPbNaRA
2f0AA5OQ#:6?0-XS3[Z4</1/)&_=CEJA@0UMCN;4TLC#ScEW=aTOO?YaHDf)Q&b<
ZE7CY12Y_cLW+T^&>3&F625\PP@a5610L:&-N+eNKLd]\Y6_aBDG3^:IGc)6:_&&
cfe:@L;\Y+Yf[--?H7O:S7I6D.46aEEF;93gTXR#>RH[IG5()@^2?&Ga?e(WXOVb
eI01EgC[X-\XZ,0D9^]G?@+cRc+E8BLLM+M=1N4,5NP\+e_]V-,Z&e[ZYI5a(V9;
JeT;CcNO,&8:I[X?Y(-Kg(.Zb?/cK:Je&:9gBb#TY)0/-e:K4\MJ^G+VdW(F@QQB
JUCHIFI&JKCf+a<S@2\7L5a/(4gP@Fe/d/2190Uce=(_>(.f=H>JYEgT3JBQ\Jdc
SKYCT)0@]N31/2,&1LT3d_UQ)Y>IaTRGH5.HF13(WS_))XG:>b=SJ9XFK4S=>^A@
c@R@b/aEd^2P]2LBGN7M.T0Y<<&;+DY9I1B9&CK=W1N58ZWA0fG=SE/1[25EBZ3[
)-SAIVGSVD(=(Z+Ig\_V71g=KAC2\LTZL<Zf3[]X#9V^UA6Y_8.8PMdBG7S+7<@c
,BP&X@:W_Y)IaEY.e##?-WE.fQQ0DG.V5ebR40S1W1S:;OIED2H8]A\JXE,==HOX
>aEQc=:DT;CbY@AA35C-M>>UdPI1YZC-E<WC0dZ5ZeeK[PLK]W.<01\_W59Y2((^
;;[#JA1N=-5&TGJ.C)K.F\7)e>7DXf&]L47V,>),B[/Gd+GA\TB2;9E1&KWARI27
U1^2c@SS#POeDW9Z6D4O]9SEIH-R&Udc;UIKL/93GY?fNS5GP0Y:gM,G_G4X@GDV
aLN0]&D4EXSGJWP?IY@,MU_SJ5?GDbfLOQV5&d7#IFe-eA.&<88<6MVHM]X-+C\5
K?gS=ga@=T2.WKR8gJ7-P<6H01>-V\ZUg=fcgO6<=bfLg2a_B8<+X;39ZF@BA9#.
ce26Bfe@X9<fHE\c)F+@adNfgD5,d-ZW=ZC09\/=71RJIdI1J\YW^E&Z,L)?VCEC
0Y:M;K93<e^bC^e1VQXDFV4XaK<_]Y?-YD,Oc^a52T#de>[d:#;76^5C66V[]TgK
QM=YeN9[#g+Y6c<@?Q#UY3,3dNM5UDI:8+5-/c;dQC\0PK8bX.cEIaMDd#>G6O:-
E7<1fUJ>dF/TG]0#CMP:MFIL@f1D+7R--aMI-CZ3I&9agA<U:63VR1;,\D8JS<f-
Tg,514-Fe&(\^55b2e_HIXVN:NWHg^/?ZMVSJQ(GM:ZS0.HVWU<45YH8.=K:O^8B
X?ELR6LLDffa)?eLU#PYdd^254>a:W37VE^(#],YI^a7B#>(Z/GA,+&I>0cD=ND@
USb3?R&Y/K@.?YVgY^-GeLM1L_C.C\5S6Q><>Q9TAK[F<W[JQ0V28ggMf[+>;\>B
\/,&J;gAV#S:2[ZK[0P_/-#V#[>U5Q<cW773>&[-_Q>U_S9Y>CD,KVeVc)3a-\Ff
(ZT?5fWfDNJB9R\NF072c&20UZ#^WG6;9#AK:3)8]YE?:QKSJc[YcRf#G]V@K^OD
5BB:8DOaVgd[(OGS[/)EQ+C=RcQ7T6+O7@#I.&e^C7gG6a&6DUFWT@WT7+1XbL3H
V(/B+[@b4J4)DYN_MNY2#)f04-(/fF1J[1+b(0eM]:d?aQTXJB9C&8feCOS^/b>:
[ZE#B+[IF6,)^NOUZC<#]b+DISGFMeD=c)&.P2\04OJVe#c)(#fM;A2[Oe.\S80a
<#]_WPJ:EfA&Q2>+bAgX:V[+8d)EQQ9I#3ASA(:4FWgBYMPQb_8767#&G7F9+g89
cU<_D)>f#Xg6X=F4-)RF=Xa?S@IJ-:2&/3\cYS4HKfEFFOQd(8&aC#V<d9d/S)#S
+S8UdUd)@1X_G>KNX7)I;gO=e5[F;.PB_0Gdc#M8@)P\BHVW=f&]PZXSDd#?AU8V
.2L#a+UPWXM<(bc[JMZ+\R@G)NSNVa=H[N.)JRO^KV]B>&=++P&3P__b+<\HXXA#
X?QC_38b0;I#)gQ44KC-VZDE5(b#0E2a2P@8F00N&5&S&&;cG2IOe@MJd;UZM81f
EL9=[aM/];,g5_V1X6Fa^#BJ5:>XAKaTGN7EE9&T,a7:7QJZ?&Kc4DeQPPJ@GUd[
7Q63;,J_AVQ#/\7I7EGX-4>E37)1&0J8H0FG@OGeL3e3ZEB.g7g>-;g,HO2b0[V6
E>CX8U;OO;C66<U,;/3,6\gFf>ed545R@_,H(8B^g:=P6S,#AH4H[4FF[+\HYCA]
R0Pa1Y_??SO)N)T07KcI.+B>O=[YH[EZ=6RfgeU5GX:&3Y):V#8RWNQHPfZ>]g<<
.&[8HeM3BgV/R)7^McM?0F>_UQd-I\W#&6T,Z\E9H3TO[UW#6U7=&Tg#_;1,RfN+
X82>DP_:c?aSbBZc<(X+W0N11ee)&[?(/5P-.Jc?HI\_?2g8?D6U\eb7>;P/g<e\
C=J?<C:B/d:)RA_21KWO&9)Ua,W+:gHR6>]+K7>W<\<gBDa4<.Ad7f>9b59aF@[O
O\9F2a6]K#Fa66M,L?:b2+U+^D&SD>0F)B@LCLP?57g<VN&L0bE6PTY84DGgQdO?
Sa+];<>39I>+<DFZ;?4,FDRWW8-\;(TN+g/bZ6UC]Q5VXY3Uc-JW]U->RX6f,+GO
P9dK?_+/8Vf519;M_[:W)[g_>bUb,C5_+>6H1.AT9NNa5.?GEBfR0L>QU\2#dF4,
1N4@WJQT4O]Ub/eA@\A/)cXa<.ULCXX-:+/dZ->QUcYMEC1:=\<TQSS#B>dT.DW^
FfII;7]_D3ac3)XX-.4a;X92.7DC^G=WG=X(d?>?=FFR;eeW4KFfI,g]I_KYdXP/
aV5d[Wa,Z#&G@(8ZID0EFKgg5B0B,;<#VS<_Z<2Z8;1KMK[JEQU0Q&GJ\SdA@[^[
O5-Z>N/I)PN&ZG:O=\F[N/:0Xg(FP@B@_Xg+H;9@,3#C.[#P3LSVg398X(f/)^/)
(&SH9[=KZITS\-VfdNXW5G.d9&G8@DR\]S6Z.,a<]+)a7YA_;b/ZD(I68V;5?(BH
Re]ab#CTeYGT48]PL&ART5(Xg]aYX9KCLJ0XNWP#F#gNY9FDOWAPX)?_F?TGKQcV
RE?:VSaS<3)\1=]TgP4Y-Y92<EfB]]SVeeKX<QV&e<TB.[G2<SJ:1a2AAfBW/eQY
=FYP+>:?DN=XVa@JeXC81a=2@);d,5;ECOCeZ/8d8@IOI)e?JaYM5f6Ya7)R+BQ=
>-gfP,L9F_]A<83<.^<-CLTc5fQgE:?4S8GMV+(\&IF0S2GId:7^PW=3SOHU7:+-
6:R2O=V\,P+A6@dKa3?_THcaJXa&/_0,U/b7]#[9d9C+^?g<a3g\T+H@7]b[,bM?
661?S8R)?85K@0;7:K)CYBWI9^VW&B7]WD\5Q_C6cKFc>R1._RK(N9NGE\>M]);g
?-(ESBS)gMRRMg:f?Y/EBX&F6d[_7a:V-S1;=2[T-@OIJ^3<SIG157HgRWNI)LWG
Ig\AL>\SA=6L?3E7H3TYFfe77JQY@:_W[:_W_/-J@/GHKJ;XJPRdMN[[8.GD(:WA
]R<<SZT,NN^#8(SG38L9)PE2<RfC\(&:>SM#).=6NG883Ma/OIAJNF?8DWe=dL9D
-],C9Y5cJ167<^6WXf,_@U;VgQF8]_H5&7IYREH_bY@<?@9g^Pf#:;J[dU>bWfAd
BNN2?=.U27(MJS7;W8?YK)R2@Na/]N-<@F;=?2e693/Y11.-L<^V0O0:S9^Le#[f
XWA?CD885J4;_3&KLdMSXH\a>7B,#+6(^T>6\6P>e3O9#NZ/^J-4#0+TAS\b6)c(
S;,dH+VC-AIa6@[[+e]165b;Gc&L_1]^f?FTX42X]aR=M\+Z;.cP7E7KJ0)8).?c
cIPeb^S]\:c>NC0&0VS@&9\<K-#R?M^2;f0F8<Vc>2-b1YX;Kc+d84L.:gfAC6S#
M_0b=Z)#_FXD^IH)ZF6Wd]PG9HHH,SaDR],eDf1].98IVD6)Z>Re+cVV99Q8<?24
PGQ:34f(9KW[P\U7SFZ.c/S3J/DGG9b)[_R_H)[YZ<_A:_;/7Z\.K5#Eb.NgEK+a
M#)X#XK.NUgNPSg,a8Vd;DTgC=[FRRPBOgXG@7?OPg(2<Jf1a=8Nf)3GM4DdbPS]
#(bDg<^dUW4,BXKA9W8b2RAJ3/V3S2\/I807_>/NYKY[=#<Bb+L+R6;6AC>00L?1
VAKXC/P+3C)#O=DW_0=YdBBF?dK6P<<2G2;PdS\J:IJA]Z,2=+,eD2Q)^0aZJeaR
b\L06b&BN6@2X[?5+Z>_[8IDJV1Jd,^0YgBW1a+;a[HLY_GDaBCY=]W?F,+9FYL0
;.SC-Bc@/KU0D&COGae,=a5>17fS[6RD>/]8;g@&V#<Z&M@LDC6(Z5I?6J#0g,+=
X8gGec_]AKe@dIdELeBT^^XPGB6KR1G/#_8dP+FWSdX>@aP]3@5KdNLOR7WOba7]
]QNDX6FV>H&_5]:SLTSSV2LF#_KLCagMJX.>>X;:8@-&HZ_J/CFa6;-F]QIY&[]0
I#&./BG2/3W.^<JARS:2+C6OfbT2R#6:YJdR4Aae5]E06(U#6;QGBZ7@-O&,,VE:
)fg+X,VLW^N]I03Ag0=+#XAE07E/<]QcLdLCf5_>N.Yf3\D584V9Z_RcOgZ#DF:6
R^R9W0e[.F[4cb.8K;T]&6Z=7HP4+a?-KXZ=>cA\bBQC-DUcMRdCY0a/YeW,aU8G
TMTAAc23DYB9_AdbDgL=4Y_1,]Y2)NLS5)D3[E1U+>?7[6)9^UZTZF#2&J&A_.U,
,915YODYE#+@Mb7B0BKCdJfO.CJLd=^)a+E2#.>;1YbfYAd@[.H8.NU2P[-=IA)F
e.ad3X4MMS<+;D,L<3.^c^X[\99M7C6_A>_3Be?O4RSE/\JLV;0,(]g49V,#C:=I
CN0()5T>AU^-KR/D2dKe#,;STD65\(MT\_R-OJN6<?]V<T1&f[C=^/FB(]NW9):W
.#TCDKd1M?7DW^]2JTZ^FaC)M2<Y0;A=<B1/X(C.R[bQ3VYEg4V/@H(6dNZPU/f3
N<N?#aT/GZcU)]F6()7RLX5[C7D;8S?NINPbc4J]VgA7adOGT[NZA0>5?XaNCG.,
X[R6IJBY=QZ+eAJ&P;IcG)U#\M1,B0V)FX6F#[RBNCQ#N1YER3318cELVD4S2^G2
#>4R(CZMRcKWXK(KQY7^Hd3Y9#LL.ZWG-:I-P;aC8H:_0:<.]83dPe9A5FGMHcbZ
Ze(@]LcRR>@)3]1]7F3a:G.#cA_+c//e>UZ/ec_BA>e31KdBd3/I.Q0]V>0Q?O>,
D.)/M9_@S:V.H7[c-Pg\(CRQ>;H#L3aM>E@SH/dd_X+@XJN+]gSF>EQDb,\RLR5Z
W#XcR/&adY[8AeaacYB/59_FC0EA&a>2UcaQWbO_P+<D^J9[FKIRdN3N5WdXWMfd
AaFMKB0]2D]0M4WR^@]@&+cXcAX[J0]V5I4LC1g6PdfbFEC_)M>](YB4.WgfBUH)
TaB=X6bbNOUR-f6L)>e+,4OBB]QQ,]c#?B5R6_=-C4;:Fg3Z]Jg,4^WZ=\cFLT[E
IF#:fD7ZLS[<>AP(XZHg>KDT_E[:caKbVPfLI7EI0Z?(:^[:8a01/bP=+8V0\RP8
IU=T?XIBf9O)^;c5_E]/T,^7ccRB^:cM<cTK7>25b):eWZ/JI>\[3L=LKMH^,?]?
Ad=aI:R0T9CcB_LBPaEL]=QX^#b1)1G)V50HQZKKJc0GFaGI@dQ5VaK<D>73:HeM
)]Uc-L<1_5S_N)fcXRbD7G@0#b0G.?QG0#V.=b97,ZN:X/F,T)+GGPQV+3@1Y<)b
,I>47&>HZI<45dX6+P8\]21d@GB,>5U_V?>:X_-RaKK^([bLH<UII)]Ida\faW1d
#+8U@F8XU,G)@\:X_B)#8[NP6T#G?=,g2NMQ)DNIc)B<YD&ObbcY2T/7_CP@fKIA
;,=Z9Fd:GW9.:6BUIGCLAO)YED:[N[cL8@_XH0@_5:Ef8W56,,T?<=gZ5_0N\f23
cVO(a5Hc=AIfSF?BbI6(=+/A\P1gMI?L8UR)U4Z@f^c_GG:Q6HC1;H7N-VJ(7@\.
4<@ge/2KY,;&0UE2U\<7]IfPSR)XEG)TOg][G(,5)M\^ZZ4,HL;[d+(D?=VgD7ZO
?ZEdIBVS<JB:&-O^O^462.L#Z7K8RK:CA>a,FdJ8fN4^/C:5=f>>&:,3aaHff#fG
9)O5]TE?P<FQ[SfLT(HG5Te;Ne\?QYV>e504Q57g0WWIAbD1MRGBG?X3?S-#]8\7
6dW.GCeZWJ[7=2E\#RgE-EN-;)L3dY>BQ2VaR]2&^Za5PaG&PPb_J-R8HM>Z:]-^
O#W-<(.aN^H5]J(N:d[c(FT^1/QA]-e/)c5G^a[ReY?+ALWA8bA/D[Fd]c9]BBTc
,?BX,&^^EAbH3#F/;WMSABA,B=;21;C-76_O(C[YCaY@G^NM(+G7dd,R+ZaRY<8e
I?BgV=bg;8AOZ\5\W:+[^)5AES,2G2MVQgbPGM^Jb=HQU)]SJQW-5,A,;]S9fCD+
BccZ3,;P-6OBJH]6&7Efe:D2AE.P)Q\(1GRGY(K70a#&GE(K0/aC6GF;\WK&AC)3
C8ce_]2O0Ud?WCE,13J:5KGDQ(SW->H:,QL_bD5P.?^Y?/:CfS4dL8WUJ?.=HM(?
Y3)-;.5.;VX-a1CeSBg]<&UeDe>A=.@0>KP#3UP,&UbGFC_P=F2LX7)EHb?#<4cc
@BPVf4a_d(I@HO#0C1eDQ\F(0_.@14Z;9ZS)L:_0P(^LI^YSNX2IZ?-[3aB[K&X]
BF@O9^/JL<CHF?LUd==7E@+4A[OKM5/B##D.CIgNZ^QTWTAf?cR&P6T1eH);-8/7
8MPQ]53e]dNI6.HX<91W@JM0MTYTA,ZRH1AcP&FcF6E@:b<aD^^Z?>eU7_498##T
R#O@UWcRM_?^SbP00MQ&cT<SM(Sg#U2\DRAg4)()XZL=._JdcHacB,bD[=?A<QIH
T-B5/)[cWc#A_6:H,#P&H[<NaIDW\E9g4B)7889B+9I5/2ZdaZ1UI7KYN/I5H<b1
_<HS1f,a>[LYHN9b&F@B>LBgbHM1Q_F<&W\OfW5.K#]C&I,LI#3=//A>Lf>[-M_L
e&X,\ZAIQ7>2]3fDc=C9NZ+Qf-cCTMOT,^&IRTC6PL5g((dA&-0;\S)BB;TRJ@aQ
K>[3O)(W3S)d=<be00TK+YII][8;F=QZ5L(a?#>7FeL5GGMf1Z,0U5G[;[Z(fdIC
(.Y.Y7H69M<CR6e:=@ae+V:&_EcHe\OgL4P3Z(U9&W(2VQI42I\OI,8+01ERSR=M
Df+-_OROGC2A/-K&\2G=9])UH7U6?:?RLVT+gP:G_M8^<9LGA=#EaV5gaJbgT?L4
C.1J,Dd.)W3[UEFR)C2K;GK@;@8-)NRN3S]:;C5U4N2>W:/2&Q47_2\;;?1W784[
=e>;]JXfF973M7;<O]0+fZRI)^F9TTcC>F:G@-WJ?#J);RYT67>a:[?3H=\_ROb<
7CN2XM[g(PcRPCb38IR68WU&\7?QNS#G+a(3>_,KFA,KZB<\0X;PJe4ME0gF<L_Q
-dIb\Z[H&4c&Y6^BCL._K9GaaeBeYNAWHP/YV1IV3X]^3g>G\KD=-Pb+9#[N-]a_
7F.(OR#^Ga]/;PUJ_a&(<0GA1Yd_Wgg7B@[X(@2Td#9(?B62Q6@7BR,JD@:B&PDP
Tf0a27[<f)8?gYB.4Nf0AW8RZH@,]B+0;GdKQ.S4gD)e[e)NIN?a/?;E.N:ZC#NP
RT>31O]=C^@4L\XZLV-6)R<B62I&\\#:Ug@a^cD,8:d&77PB4g6cGG-((>^dHN+[
AA_Bfb2M>H4?T-+eW24]>]5KWS>H:TLBI9^LL47H@/;M;35W-AEU[YeQW3,1B(:]
TaIQbL6K4PTf0#2-<QW0;S;PS_/<L,,PFY0588;eYKbRX/X.K7PKdV>._;Cf5LWI
bFK^ObL6)GQSPEA+B;0I/VIGg2(>\)dT26PWDW^1I)d#EBb)UQ<-D=b-d#0,/Y45
=46#1c&E:;/J-8RV&K\e/JUW/[d?F-bQ?dE=J;.1OD;G9VbT:(,]McG88,(c\7+L
_(f#VPWN5XLYUJeFCG8cXKQAJZJ;MEW;\+[Qa:((YW_TeG3(:#:DIJIT9IM@cD>D
7YcK6(g@,SH.;826/a6g_U8>26>UL0PS;dM0GY0)3QG#Ke<K]cVf9XP>_[VS:>QE
MPUBaL1GN_UG@I2K+]P79QV5WXX,L8LN3NaOA;WLHS=D-.LT>F7.UgJb&WDP0G#+
KJO,)B=cdXRPAcW3UB5X:OW0LIV8S[D8Zg0L(WA@>X_[V4S->:eOLZCf7F<CS>^)
\b4X0-IHC,Q+dD;^#<E_ZEg(A9E-.OR[We-g:RbgO9:26LcHRfaWFS+:X\F8C&(?
c,C8P5M+W(=^X7@QE,6SKRY+7-RU945=1]A_#\@[5.WP;OH/7E)0B90:_ddDGB/Z
S12OA(ZOTORAD2b=56f8GK&?D12)U3[5+EL=AYT,A.MU4FfIAa[c&CgIEKT82R+K
eAc8LZI\O5)DJ5L:T^S^2>V?M,<2WV^&]=\,=]ce/+H6Nb\?3GPZ><Te-RNGC85S
V&5PYbQ74DO\RgZEB]>(;;<O@0ee?]ZCa+;#?EN??fTK9JQLKC6A/R3(6:Gg([;f
c:TZ?A:C<1M+DHEgTNXHLJQI>/J;0=5gO/gH^_TFeB\URDX#5f]>a]-@3-DU_?NA
MWK4&8PH9,1659Y>#V.)-,2YL(Z-C]2#WL_FXE417g,f&6R<KKg4YMK/XD_NJ3J(
FM2&9WDbYU<\J57f>W@,3\FR8E1S(_/-,6b/c48_aJe;?e0/fdb<A/.0M\(YeYeD
A^/D1O#S35911DRKZa+FgV+1>BUZ(e3M&^.T8^Nf#/e6YV?/@=AI,>=WT5BgcZ?P
(_\@V[>VRU@7D#-\]cdC@^,V?IK0Kfc@YFHFdQW#V6.;FG(1ICC1.O:HPWY2M@SO
_->OcBV5LT-cX@Q)^&<a+<BW6M)FK18@c_JLBbW[>BbUeSYD+-E@?OSDFGSPHR5W
d)-UgO;g1Z<gH+UH:I\HOIF6WO,@AdW24UY.7\=<G5VAM4.3HB\)W\1^cE.@)b<_
[+aP95ZQQgOBH?LPD@N0f@=-HEQJ83;&WZPKc8J_X@ND@)I2^^LE[UN4LF08_5I)
R+bOUGI\1T;BbZ:<V,?fL\(M0_e[aM3CGcK0&b=7a]9Z(TCW/@F65?KZN@FH(=F0
LTV8RWeW-A]=9FUfH(BWV&B8[RYS8P<E0caU.,^H[g@W,>,XFfAEU)^I5aGDR>Wa
.H1=I(=Bg3OJ,#@&\<_G3T:C7_=LA8^H6Gdea&G_Bg_;d[ScJQFc(Y^LRR\DAD>e
RcIPGVRQ/JHPDH?=FQfg/(S)^3))GWc(YScgOT[[7(d=16>3#=-R2T?^?f^#f3#-
30=a.\QG[E?PX=H41OcB[P\N:QVA.fKg+\2S9C-9(6#3MQ@HXaO_]6PWXK2IBBCG
WdL+;@\Db1F#,42HaZ^MCFLT8=6\-E.E5-BC3D&7=^TGB9>W_OPMMU-S8XWCGR[2
X[L:eb#>):YX6ZI#6^X1NY2?^PJ@A^@?UG^:CW\>Q-7\<C@OKc=fMCWT;?=]C^]B
B<U2^K1;.28+.0J_>Z-LSOSgND@D_2TMbQFU^I7?(I4EIe2Ud>3d9>X<a+/[Z926
^fPba[EA+Oa>Y=E+ZR>2.AYZ2[\F_a)eVT^2M+7g-XKe9H@>6B](W&_.VA4F8EPA
36IO+X37^_ADXP;K9aU:Rc&fB>a]bUH\-]JJ._V)C9=DXe4<Y2AaSc9NNF(5<9dN
]2Be8@(T_#I5G.[-SQZbg<-#^AbICK-8Pg7K/;dPYCQYB^;14J__;497OJ(aT/-W
T>P^8XbCG-+0eI5<A,E2,.-W.?a1:Q5[Yc?;+9]\EGXCQeOJ?&,I<A^bWK2&O4DU
X9R;D#ESZ_?6B-:7@>N,_P(6fEfNIOEJS&_YSEOeBZC#)^bL\^H2a7EA_<RAOZ8\
B2,c3]7-FaB3M<77f\\H/_.ZZG.9Of5?__D<SP3Z8_B_#N6PN=dC1/Y#]T6G)GIR
MOQKC4b^U+LK(=QP0T^b<E^g>]f?C98][-^1F?^aKdABO>.0\+]N2AZbN/=aF&Z;
]SRZ>(T>OW-@dR1_g=#H4?:M?KNALUVLFCc7@A:Wg<8/BdTV?fX?;:G59Gg\-AQ;
.L80EeNM/CgLMaZ_a;aO5W_5>/g(1dHd[4K;EI3Bd\IH\>S&GVaL?9X?>YQI;3#;
ZC)&P]Pe)K]a@X2S)29=</6JZ;#6?,]IObEce;UH5:T=,.D?4+894bU]#<Z=C5b=
cggB)9B2KEJ]Q)JJK.bLA1FOWYf-?IMTG<V.C),BB;<g</fS\.(?,0+NW9?^MeWS
PLCdcf>;4LEP#XfTKAb2.>JG+Q<M/G9>QQ3B:=H85FBH4C2)Z9GC[O46Xe7U0Vbe
MMGWV1b(4?=f4aeUN5(<O7V<\Z:K#R&Z(K-L7F?-FSdeK4,]f,D#c7(DR0>0aRT(
<\F]F0;N+OU:F06_YF(/.dSd0-RV:EPbQ71WGX3AS&D0)9B7MCPLC@]K42Z_/I2-
6.V>^LVfB,-LG7I5CAV\>/1<dJ;5UYO.G7I)R&Y)C+8#OP24eS._M(^F&:E5UF6N
VAVJ]\HPP=])MHHIb^KX>#;FX>N1.aSQ5,)?IWTCSY;CV9;1J/)=U6N;1=+U4I>4
(dS/#DD+R_e]O0R@;VTeO@)9Q^\+&)0gETgefJK-2d,Bc)W99cF=8Pa:MZ]09LLT
UO3DMVF#6dX-f]+IUKB2IYILGg/<V:GgL5\H@>STTJB+)(2Q39&^Z9N0#W175;D.
D)L4fIUIK4/aRN5UBL/39EX&52KM5JP6_AfPPcOgXVJ-H1?Kb55/\^eHD[UD7C[0
A3=)3G?/V,],^UV7VNDN^0ALS9U@G)R9a:<X<KVTHV8a#RU8D+@b&HbRWR#f;Bf5
d#J[34?J\fZU8]<JVMUE[;<ac3)+D_NUGN:NQ30F9O/X<TJCA44A,;^7P;Mg^Vbc
/(g2:S:4KgHgfTI5OVRL8a[N^c)f]IG7ZeXYb^bF_.X1D9AD)O^FEK^0=fR4S:V0
e@X_+G,_b#e[&MC/9L]8,I@DJ9PAU-UEZ6W?:)EF]D;&/.eeP?;=O[&a/,]B/=.D
>f0LB\/+6)BG5I2Gg2CD5HNXTH#N2,EfaYET\_]C-0cOc8J]#7]1>@G2EdHd7)[^
A]P1I>-Cd^FbVDVR5@e&6Y7=,ZLV#;gT84&8+7H.1F2K2GU\;Ea)cU(5]\Fb_)\T
0U&Sb]_=N[)YKF(MQ_;M459JVOB0>VPeb:7D)ITeA.PWgP5CQ_@44D(I8Ae=^:<g
dR(4D@B49Lb9VO]V7/a^ac&Z21<YVW7d01]#]_DNWN[=LYG,(H#_:P-BGMJ-EDKF
gaX;1)C-^<)AQgKgUP]Q4AZ).=2?YfgLg\5]6T-JF9;4YIc8M\R>0Ub,1ZU-WC=6
XE^aF[SLADC^D8dOEP_fN6V)^?^_9-cQLcNc_8]e9gXc(=^>J]L)Z7C<B@U?(D)1
+6E__W08A,YG4X3G=GO-[,M/6^aa]W?^ff,RCR5[dF5a(YCe7(7JfJ[QWcOE@YBe
b6TH5Pc4W4H27Ca6BV+3E2?SI@Z4ONMbP)/UObEgKH:@IR59-@#<CV3R+.8?NTIF
EG(VISfUd41DHA=aId/53I5f@QZd1PLN[>=>JYOA387YIcVE@80g^?XML9a;VD;X
.@\&:-ZU\M&Q+gg/P+CG_@J5-+I15:^7W2S]b6SX,4[@NJ-N7Vg;LQ4<AZ,KQ,Oe
-27E.W8+Y^I;YGMI5P&VDS3QS+/L=CUZ(NN\A1FZKFM@QZ3:2dB.--/5)^^O4)D7
[>(2ZZQc\0T>/W(bAZ:R1^&Ka8#7bY4JU=JIeJf&JeZ\REK?;R.5QUPXY/Y5Z>L?
?3K+XAQ3cNL7_D4?b8g?F(+M,S]7SX()aJAaIY<bFNAe,WUUU^6840=bP&dU8]8[
4a,>2R.>\8<JIBPCJbLOKC#fVM.7Y8a_JACaO(b^4C(=/e,#?\^).OOZC&=UPZR^
?d2C=:T,]^R@8@U?8@C<-B_YFM2+(<ZW0A6d&D^2(]-@:O1^+O@K^KV\M8DP/H[T
Aa)0N6K8cQ;f1Z;:[X>3[?TSRCaaR5@:?N>1MW+--:5(,1W9:XCS@aPMF#_3U)PW
cG4[<DVbfM7]P13(?24=G2Xc#H35I+G3>]c/V]cLG,4\A]e+/37cP0]+db,0f?B0
VOdA1KF1[LLO.BD_9ROLP4ZBPbNd4^Lb>d2-=Q+8U;/gPX0KQXaV=F/@W?-^YS-A
??#N\K3FX+2(:abdb1DcO6+^dfVXg-PTHRH90EgD,+M0:0cE)@1LDe8f0[V)R=?e
J[QW^Cg1L[-17cZGb1Lag<E69:DZLY2:eT\),II):;Y(>eUEfP8M(T>]C#8/>LM3
e(S?ag]^KO(QLHOO3R:@>UMC>UG:W=PX&\E:^;b9c_\\2>1X5@<<@L#C@7E:7/J+
Ub+G78O?=2LOU/80(:G/#DZ=Z#bFE(=_8PB)KB33-Y)2]#PQ?NOP4TM:6cG=VCQ<
2)5Q#1gc]b;0.Og.VVID[+P7E[#2ZXc63,B/.[<-9/TdL-YM&72]1YMgGS3[<)S(
9T9DaPW4PW773._T&UV8f[<:?9_\0>D_2.X-#OVeM68?-@F6XaZA]7)9L0O6Y\Ba
&=EMGE=GV_ZO/:Z>J]8]9+-<@)e1SC2&FSM+,W]YHL7OTPW1G\[]>-MM)ONa7LIV
DHO))aYRcCaSKM8<8[H0Ug9C=Ce__SSXO^P)KL]?QC<TBN(9dJ?7):KfeZKLdRU+
ZdN0_4(a[.:[9X]3G1KbW/X28@c:)?KMI0f0I\U:8gA?Q_Oc-T5g:Hd9+?P)H3P[
;(g5Y6;6O3:-D_76<fJS@,d#E]_g7>,K(d2R<?eW\7g,1]FM(A<.52U]>MM32TP9
YPXe4^1(R)M.<LaFdINS;P.DWVZ:@Jf28K@(B(16=6,F92c&OC7e>D>&dYBJ@;DW
XU;\7L2H_@[Ab)c_NOAX<YT^d9FIX;;1eLXE<CDID;T5+eLgDR6dGJd,NQV(=D)N
VEM.,?_<:,)\45bUYXH.RZ.L/RO&)D9E//?K\33E\[<W1ReQIb^^>_2O&7TP9(E.
f@?U[06<bD+:W=-0PY(FAOZ<A7GIRSZ8Sb]RBXG&9a:86(;Y6UU[6:d=)ZM^\O(P
BA..8QOO/#8-+WTX_gSfHI&c>a,Y)T730TY?aQMVd7I(XU^YI#,5A(eaLc^eYa>T
:bQN6#e^e\f\=.ET6f62[1A;d4a^V-@eK-;fS.g[fCb.2?bA,.:HfN3A.@^Oc)7T
BOc:BX<RYX@Ke6@+7M_7>FR01ZTb?8f+e7a],:U7O^H-8@B7.HXUD5P-D6[NRdEJ
F/&Q=#dIQLYJMMaB[eR>K/_g3^gZ9f607[9POWUH,dP.)T^\L):L+1&69f+@]Sf?
9=7)U0\=/dS=)&Y@O/)U[VYJ]DRZU[B9J1N5?O&&gR(U)R.T\7bDQ&=Za0#YBXH<
gCMQ4V,OGA@6YM4#;723I+9O1@aFaHO8+f:)bbRNbPa6g)c?NB#1ZV-I2:0e078>
^H8b&-F8:7bg.d2RO1B911_X:fJeF2?aV];J?^Lb?;YN+c8)d:G&L&)Qe,dS2HUf
d9<aYOHFFSB[E5K>1^Y.PgU_@>NKUJ4/bZH2_0#+e8/_AcUD_Q+28(\#IWG.=@Db
:ET>KG\fGZ(^6K?b\EA^BKU@=Y?dQJI@;&<FcF?c:dO2+/@dB9+5cQ,32#(64)g/
dKOMPLVU&5c.:Yc):12]5B_=I90Od?5[UP]CW8V?]/SDXZ1.B;f&?\DIJNWb>c/Q
=g/Z1cI_E,RG=0Od(.O\(RF(G&H8:,\ZUc>PL>#CA(QR/\4EE@aS@_V+4fPCd^UI
_@H:1g[>.-bJ:<EGE?feU+1d\_)JI4Q=]:)g\YUaYaT3eJA4f#1:_9R?V5UGe2F5
41M]0a0\/d7+a@0E8fZf,U[g<[;^Cb2,EbB+1TS(<-Fd_UWbHMXDI5MYQaJHcfS:
WZ:96C:8\:P/NIccTZ)e+c/J-T/C>_<;bPBH5)EQ>J1_,d(WQ(TWJODO/F.e=ZM_
<AcGKHUFfWg\#0E6eLF_69g4MO:#98@c;K4W=55]bU]KUJQB6D&GPID&=2H6[-Yb
NE8X80(G#7+M#USG->S+Q?;b#>II;TaV.[CZ[#\&?.B]-Q>.ZT6Q0b1ZBS?[9_:2
Zb-ZJM:D]G&2_YM]cAT[_9SEbU]cW.FOg4(6V(85XF-e2/R\1)UP6W\Me],AEE;d
^+E0.UAHe,5;MB@bf-MgI^c7&7X/1A(M,W(<c3#2/,6B+-G/.VgH=\Z;+-fYOc+V
B3\Ng9-UICMH[[\9T9B)=VPQWYa<LE;(\3F0)+=V1af,Sa;W>(\6(T7E5:<SE&)X
#?HU(e+,fJT<dI^+#LdM9:#d5c;3P:cK>:TV^8GP]=28?#IgVL<YSRZ>(e>dV68X
K-QJX^3,K@9DI4gH1U6.CdE9E5]fZE;CRGZT.\QFN.?=_Xf+7;9QSD0c-1GH):L_
FY((2Ec6VTIg)4F5_IJ>[L/N>1IO[K-e=TCD)#KQeV3>5Oc4#9,Y>GT=;G?PSg-4
6eGN)1;>^EY#WTd=J5bUL#&+5JJ^_#3=^#HDF1e]/D5&.\HVTCbX#MOA?2.A;I#f
@#X[gB+4c>_:2:K3G+PDfB\2fV(P?/CM(5G@WD#ec;]AMeTQEPIe8fD=/M<PQL;0
1.5_Q;GKI+X?4Z>JOa7A:b;a>bSO@&Q_]K3:5SJ/W(1gVB5fbI;a/dagLLfF#>DS
[<TS:)D_\#cX,I]Fa/cL>_@:6Sb-<bHdREbJMMM]-^gaZH&8LG9TAGH6&])_4bZ8
]#XX#W)]8Xf/:OGXe\UV6?_OO#4^KW:+RGdeQ8=)@<\8c@Q.-ccgE+\=.2T59Ka&
#H].eeMfE&B:P)dX<4#<WEfGdd?)eZ([PAB:G_cENTXNg=])R(aQG<;M>PdUK@(d
[J=M./FXX4)>,U:ANYM9_92G1X?.E_:PRgC93DEIFd\E1UHE+_?7HJBg/FUFQd6&
+:IOQ)FL=-G@U[fW^^V_631f@K62I&^^3(,c><_V]H;b\RY5GLHVFeX()D42YX=T
f9bE/84K[@P[_(c9a4b^?IRJc.)7E-cP0NG@))&5Y9)LbcR->PNUa+@^=;P0<UXX
42B-b/JO,CC;DBgZJ=5SB^>?KbB9R(T#.=,/NC>Z[e<\0=XU?Xg&^,?8^?[X-=OC
53dbYGC]4g0BSH@0JfGW\KZ+=LX7b^O/?8X8[QOH&F9.Y=S)F[-?VWK+NX)[NJfV
]R8IK4]Y>UJ[?H_-e=:>DDXO-;J47U&ZQg21V[;V(6RSe1Y5MUHU7HO#bF:FF=-]
[1IVK3ZI[J0/L<g0]<?E,+GP2.eUI=VaQ#0e=_L#=b0DO1FZD;&+P@FI-U-V>e1J
e?\eKF?[Wa4&PePJLKV/19ZTEGW8KKJ=L;/8.IRE<2H2W=[HXW72(?XR7PZA#NBI
VA]4X__(&TN_BcM)2b74\60?]5OH>99IIBB1Z&XMYJ.AcYSf8K3JJJT6EVJU]PJ<
dX<,VMLb=;66d3E0]X9,NE;d9TM#EFU&c8D9OG77EVN52S\78-7dB,62:HR:3YJ]
.Wd^#1JAF8E)26O/C@O&H=e&]d02GLCL14aa._)P6MOAAO]aceX2RMK^<&D]^T,b
<95>J-AU389c)WR7W>AOOR]#dQ;ddbD+ZR889/NFc3-.A=88d/?)\6:>E;7I9--4
RgbMcRX)3,V.(R3EIcEF^Z^&/9]9_3,gQ3R6feEVSg#IRceOUPKf2PZYI3^,^e/d
8.?FJ.IY53CVD/?[&bL]S@fO\.XdM8=EB+Zf5&?BP]R71Ia#__Y#Xf?R9XcUJ_94
/BV>XD[_+;E\/KO:B8?&g)fDP>S/Y39HIe5_>NHLO>TV&5CPO2e,+H5ga_WAKeDA
HI/=cDMS6\bLM1FA3fHPgBL.c_c:AJ9P<^KDNY#UC_OL@@S2<ZR70P#Q3(O_RaI=
+U?dW7FHe?;+UQ_J#?gACNgFgE<[Q.DgK/2?_8>I_-PXNZ__X1-WE]f.CbIZ_0Q0
gC7H03CM5=Fc[-Pd7E7+WTWeUGBAEXC/-1;-O7A^&PL25HTD+CQ:e#2UBFG8;5@Q
W1AHCDS6RF?(fR4T2f6Nc^VUM?-^7_6(ZTa8DH.QWcI#,d2HQ(]TI?c&CW.?Ug1d
0d[bC_S-Ye>R[\Y.V1<,5Q]<d(?g/@F7W4+5@LP0ca8P,0KWHeM@ATY7gAE8:cR1
W\F0@d8_/:>QVE7X]bSD,K<\ZaZDEd:V^FXT<1-UQUa_c#2<VP4[#cVCIHY31(KN
A[5M1LZ^3FGOL8MbKWH3ABdRPTI-,VL8R]Z:KMJ^8_O092d9U(.BYBCUFR(Cg(5_
TX-OE<9f>_c0,U3Q7f&F&:VD-^Uf1]]L+aY+P4>#DN,C8T@\5@M)R[J[,-C[=&+3
.&,VSV&&GM1M-50ae:Cba&GYg9?<997MNBG^AP0U25-?gYVGSLcJO^TAN^7VL3BR
[#UQ^Q=(/YIN/5A-773eOEV<H#S)FA#5BBX^>KX,+0<Ng2(I1SU@K]#=K]c6f7Nb
:9.=b5-+KYd_5+X0P8dLM28@]]Z,\8<,-DX-6dY;7O:[VC]07KQ]^&d3bZI_cT9Z
NI,17B)H+08W2d.fW34JT]3[7>bBP0H#6QW-A87HPBVLI)>2b&1S/=g\VU>.<F;P
1=,O#W/;67GO@<W;ON?CfMS2\_E2XJI0X@V=#E>(1OE3DE?=>^^(:2Y?8Xa-J@[)
c^cKgN=+M1E0DD[Z+9V/MB<4AE5d\4fH5b<1F1?M7IT@>IH9E)eNO0;^I/QTE,<f
7Y27e)[-/=4_Wbd7GZO^ZWAKG,T<E?Q_66:/=-;5@;&WAaQQ@[9FTa(Y(RZ&?4;1
8OZW+B=0DI7V9Y@Tg;MFef7b[N8HDG_92<FDJ.J_<D8C26]P:?fUMLO82EHBK#Od
MBMJSc7eMV>94bXFb@H>II[MCIJ6d65SbZfA7KA:^DAWJ#V]<^K>cf\S6JTY_DCM
E+3W\YJ,Le>YQB1ef.:IA]IgP]&aBWY];0IDT@c93H=&R=6+#,&7<\0-?H_G@-JN
NO.P#GLS_GXP2:M-(_\aD)@[0dCJceC@S.gUCBY1+QLU=eX+7.a/@_END,3JgW,S
]1.PD^GcRAA/3M;)/>Vf[1.B&QCS>YH_\O0U^[;81?P<&>DGJWb]>P#X];6LOHRH
?9[F,2DY+BbOL.@;;)/O#4-HT161fK)/VMIPd,_R&g_E9X.(X[AYOdOgBS:Rf\EH
BF()OL^H)IRYEW.?2FDOf]1OTJNdMZgYCZ(<P0a2c:aZG-JP]S^1+5YD54/^0VDW
2H:UU,SC,Q;G^[O89eEAOc3FC-)&WK30-B>.\0@WQ:(;bLV.P75:VVcKI8C0b:UD
=9T/2OF]8dJ>H-]8_93-VL#Y3#cBUQCGAbZ6,>6A/922<O02?HTF<;2#4;YK94QN
-8?SD^G9A,D8&ac3H3eJTGK<I1dVgfKWU)HK0M)Y)C)+\L1ZTZH>.BIQT(1?WVMU
LcSMG6)[Cg..eVDTZa#A8FI_SS0-2G;NH(?JfLH5e^f5P4BSHX1,=KRIKWUISDJ&
0>?U>7GPG<4+WZ)dHEA]L</\L:+X\)(>Z9U3><Q7J+CWSF>0M?gDS:J(FT_C7UQG
f:&7b4#[g,af8Ub[M31e27_2T-U[&IY^90,W^-1.8-8(5fa2VG5@Q\6S2\>0f:fc
.6Ea;65D_#LcG6DEc2a\5QYc(Tc//^UN9bTZ>(K_.c53g<-_bY?WCI(1e0eI&M;?
c+07-R9HHOFZdVHIEc#6:MK>(D/QY3X;YJK29K+,\CL2b<Y13-c#N:\H,E_Q/TC8
R@(OWL]dY=[V(N_I44#9(QNNT.ccA,7\2_/ER+?7,g8@--H6,_-:]WP7J,6RC5Z6
.B(^/YSP^V,f_:a8=,C[9//^ICY+LGg7Vc_/[/YBIC7MKFK2L),ZISLYE>@+/O=>
c6>+E5gVDAP3&a_Hb<JW]^;)]M;UD)=&c=KZ/#5Z^c:&J:I8)f^KCbdFK(E;+@]E
,eR&0GI)?03)E8G+;LIDC9[HYZJFgcPTWDZe3>2PJU5CYNS5-L?9Q\8>eJ/]JOaJ
08:B##cG.+_R,Y8),_;bNE\2FR#,[I_KdSB]-@BMU^5?I\(gZ98FcWKG)7X1KM[L
\0OO3\.=+^#I(MJQ3>\5/LKId84P@:R0gdTW)WS@+VS?]V;NFS#5<D.=O#8G1/:W
=+CeG4cEC:FKa[L6FSG.V#UgW@3fV=g0eKFa_fGQ--54J93f5PU65ZZA=:.<+DQE
77EI#]Ngd0^,Wa3N9GfN9V#_:8WK#/UTB]H2FKE>GF:ccY=K+Q^/7G#,FIYa,JE(
A,\O/W-7B1>9Wf)U6g9SEFTU:\-)eC=E8B;GH14DfL;9\[#NW,-R10=HS#>d2K5,
[)f11PSZYIKT1XP?ROP6Ea\RS2&6=-@0K:0#H:cQ.5]M\YTBBgSH3_I9:]d-SROW
U>C>)Cg\g4)0/VRV?Z;8+IUVO(>@eE6UOJNWK74\MX((QYX6H&@+E3P5GA]0g&fX
-(N(7-=dbHUY.T>>\K=YP=;NZ(^f/QeV:;G_1.]WNH5AeBEVg[8:Zf?D\\I7dF7B
NLX320N:g\@eK1K8L_6X7U.c,dF5SU+PQO43Td+&9g>/OIUS?7?]1b8OG8><#.3e
;.3IV.Ld[.EBcST]]:Sf0b_^.M>KW,7/cQ<;5c>JPg-SBV>\UX0f-a6+VXW5e,A7
P&TZ^1V<^b@eP#eZ[G211S5B])?J\c]\M=EWGW_1CWaCH@4@>XYE2OIC/ab.d#J4
K[)EKMZ_P-#X9L>KAAGGaYZ?2e<.Bd;C3M:gO]&,dQ;eL\<2&Hg4+D16QA\^?Mf8
/Ze0#K>):4SHfZX85XTV]XL;W]QY.F5?.4:P2X\bAcN\Ea/Q#\/0/EPf1Fb5WI;N
9@?UR=VU3M(1c:_D_J1[B,MKF20[7A>PUTO4+&=-8d_Za/X&BO=TUg1.<_&SGW4:
DJ3M[,@f@SHP9GLc-8bZG#4ga18=25C1A]VeCA-5L587W0,cQ],<PC+:3E69<LUM
H/F#-7fI[f3ffE:;361=?NJeN13J&.KQJ+Pd4/1_aP88,192ZQTOX6.J],]/bFf3
)G7##9EQA\^g-5W^/-.Ag@^a2.gJ.?SY)[T5V@C@.L#RUcHD[gRE\gc0Y-WceQ,H
C,UDF;Y48@,d2NA86YB=f360AX3Z_1&+g09T2YR5IV&/Q0FX,,KP</+6Uc,_9eK<
>Tb+H8>b)GX0<99^,]Z[#JAfOPOQE7G@PZH[NFVIWW9Eb=X#H_Z8:RR9c]:3R4/O
d5?+e.Ed;7;6e]UUgb@]P0Z=1@ZM4<e3D[Z=V;_e]&?b/4K#dE/I#N]2VAa&(N/]
]&EdZfM7S]?;H4bAQJd7?ecO7+WARc4HRY4f]Ca6[:V)dFC>,#)833S7fG=G:<1H
JDc]JJHUM\B[]FSK>+BAaN-fQ9CTZEb.:dbT;,3<#T@Nb-_2U:dg=8Xce+#E?7;8
=BZCT46DJg;.&g65<YL4?4HE,L.9Ff]Mf\Tc8<#=NU\C/M[Lc1Z[NJ>6JO(.GLWE
f;ODF&Y)>Y,Q^cDg\^Ac7AFJfJXW3_]QX_^P.:0fAU5O85U-UOD?BB1.g=.MPZJf
PG2E:,9F@E)<45/eP@a&)/@\W2=Zf0aJMVb6bI0Nd>X_C&C<\4&:2SK_J-FDN#dU
Y]>DE\GC\>\VeJL<&cN?F+J[Bd8_M-Y17Md3QD@4gHKd2]d8WFg.W0E+@&L5NNKQ
C&9d\:=G?OG5S><Qg&0L4.CP6^PF.,f4_+QI[J#?58;FJ.e4d3-:S?aA.7.[5,5[
&5;]U?-4ERfOa6O6XV:YVG_gUe.]<\N:AH[PZZRV<gKZ[Z\1W6U&V/Q^1^b_?+1D
gPGcY8SAb=GG4[=\d_0UW,Y-c&b#=[-^:ZPV:g](.b?5bX1Xa7<gLWaCcce[7#VX
+G3YH++&KZg,]@TGO[G+FHODMZ(fCT+QME]FBZ+L089EGfANO+=T-PNR]:PQ733+
=(B;)>Td6MDT<BZ#U]#/PSB;GWV0L&2G-5<4_G;<BU)+YWLa#deBPPN/O9OQ-;#S
)\d9>U1+.e\TdJQDZ:6M8A>2;>TaHZK@STe^@RF8b[/QA^WHAKWT@2=g5RXI[K6a
>g5WA-4Z0G_WVXX([Y(RUHOU3I:CO_2[O7GV7AI-:4E_4\<:@CF.=0TFY1#]KS/;
TUP-9c^C^J9VM4;5YOJbL<bQH#SZ9-VQY[J#,7>5,NPY0J4GHPg,ZE<f)L(,2>d-
>@BI_?1M.U/708\ZM^1=W/K7C_=IX[DKY/8BCE/BJ1@>-d@]2g5)YQCE<?J]#3f>
/1BVZJ_4dE)GI;Gba(G-PS]LKVgZD4dA-/O+,R<OYgcENC,?g=7\](+V-FQA+Q&B
RXdEY=IE_Z,C.O]:)M,#E\>6>bMfFO0<H;(9Gc__L0VfAH4=;)CX?=.+V&C7X#CI
M661.\]9<8c5bM;PGRc-4,#.gQXb?Ib&321#_Bd?IDN+d4<+d9,3^I=-#+Y2]a9Z
[)G0CXBM&D;5G,-J_2/H>P[cHD?QOL,OKV2#A>H2N>PLEZcFgfD:CeB9b]^BcU]U
6HXNT,AP9ZM223IT82eZG[8:aAge\;FT^<DF[N[S-g<&P^A\(NC-F;g&4D&:?IgP
6R;JAe5FC^-7ZW8-I)Q08#5Z;J^BdfI99)P<Z+U]OD,BUUVR&HK_&daP2N-PLB@;
_@]X]RC5M#[L&8ZS91TPKA#3=>R+cYM&83SCSbV?9,@F7S]LL)edV5C@#fB^^(c]
_E)2\QZ@#T9QSQ/;Hc=Y8--SXP:/A/?,Ga,]gF^(9?(GI&]UdVS45C,]@P&F>[-A
W/]JUOWbSM@BRTf75XWCBLZZ_H/X.dM8XOXUB1SH08NOP0Z2M_)?0[LRO=d@OfLO
(/[S>6<N6K4gQV\FD_Ng[LAO,M3c^F-(>=agAJWZ]_[6egHHR+T:;F[a((1G/RGR
SRJ_P/H1V94:Zf1fGI8I<#(V0NAI,+D)Od)J<P?5-QL.22>Je\RbBQNJ[6.Ab2).
P:,JFS/^1>SWJAL=e&8=1ObL]N&fY62([KW-W7C^DaAM1W<V,QN;<_P)H/#]C)AR
aI,X?.=CcVA[U=];KQEPD[CN/+K_A((ZIK\[:(=UFWeAX<4AIZ[N-ATW5NVBce(,
,5?^.F>aeg3^[GB@J+RFe6M(U1C<4BW:H8COI9\35,U6:.B-/;YK]45>_HID2,JS
1H6#/Z=D1bQY^GZ2P),W?ZeKY>aU.V+;P&MD)b8+1<VJ>C?Td6#SZPCSFM7#0-U\
@,I[85aI:TBNPf(V98Zf-WNZAgWXHMLQ;_-@ZI]AD@.)_FHS2,V/,+H[ec_.5A))
U);S&2M(C/fW]RX?#JE;(5U5E[JP\1Q0UPW@\7J#d5U&:90W#Q1K[X<EX(ZZ5K/4
^I4Q/<RG,39LL8UG8YKB#-QV_A[Gg-0-9FPgB;NL07,-L2Z-=YHS)#VXYHBO[/L;
NG:#O&EY.:Q,DaR2F4O)4^DeNA-KWV,&DA^DNKW5W43(3A#K]N?d1a6BcPR]c@U/
^B<Z:G,(TE3[1NWE]C33F-^WJbA_IMRZK7ZEP_5DK<DN&#=c4FaIc]6[T&MK?Tb.
fd=RF(OS#/f\+7fIJZUF1MD.b[U[L3c07B[D>Z65)A,8cQgNa<dFcdGd>J;##PR9
FRVU\S+2(RRABfEGLLKUggH/8\_R+.MF-Le--S(7^;+X^)5adGR6BJ[<[O/JL5=T
,&RO-__5dD4SgOW.=4Q-&DMI>0HaJ13/5@]Q^Qb]DVMOX1QL8G9Pd:8gf@[+D?Rd
5F##56+@W6QgN/RJVG#Q_@TJ&I?1HP/735^T.QQ8:;Pe0BKA=a?]I7)B-F:)H,#8
GYX^)D2NV?+=8Ga0U7,VG3\EAYPYC2S.Fd36QXU9)OZ;^e))CA>cd[-]g]Hfd>>>
W<g)/]=;ITI[O+?^HY7X6CN0=\bVB(8][B)[[#QS#Rc]KeL5@>e-&1@VJ&6d5c:G
?-NVRb.P+6AW#6@Ng9:U:4RfX@GYZJS[PNBG6Je-#&\/g.Ba5PPL9QccTMTPJ78I
1?F;T/565@0AM0>D&&WcIMP]U?T/^/28I\PJ)KK4I4<<e/6KLRKO#Z54cR,9XU\9
9DM[eF]CJ.,)>FJY]:#6_+e3ZM6Ge-Y0eaU,bW;?4Z0(J#9T(L?1KDX4YcYE,=74
BHQfJBWE9Kc;ebg8\Wf0N0ab5>JG/6a:&PB)C58<\;VP?26EfT3K)X&XA)NfCbG4
XD97b?>AMI7aBZFG5=4+[Sdc.JB.R6V7Q\IEUECLG?PZKOS^I<P)V+/DEN7Q:LO^
C-V4He#-H1W8#BZc:-+,#9KI)6XQURPg37185@5#)(ML5Og-2G=JW?<&GG1<ad]-
B69GRI.f:\,ML7C58g^aTO=6U8I0[C?I;K]2XbPg]DSY/F2^3GNPH,;]KAQ4IAQ,
=cE)1FA7IWQ.THS\&N:.aJ?)US@(VT2[M1)C8c9K#^ETC+ERKG)[#]7IR^0(:C50
^K+),CLSUGYW7P2aGgaG&(HO-W@.>M-HWS?&9[XA_FH0CR]D_JFINRI<BIS_[[7Z
[3+CFUJTGK0I3(=]GB[f/).UKf6/U0,CS81IPA)G3>IXJ9^4e&KTGSQ0K_6<]D;=
^&HB=E9e67K8:M5cg)J]c2&GKfBK1+@;]0_D+:Z<GcDZ7Q\e0J^O0Dd0/.,B,NEM
(aQdYNGb,;U9ADI?9B(..DLQEc^H\G8B\4E4K>1/XR@Ab]&-<R,f<TRdIL(;)BW\
8-I>:7\W[V;(Y?Qb_MQ+TT\DF^aeI-e]KXT753TOS&33FV6ZI52CbbA5LHD&FM:I
gZ6##Mbd=I3aCK);:V8W#<AU5TQ^#G+4B4N.+3KS=MMM(gRP#^;7.&.)IaUJ(\I^
[9)/;c)86M<UH0/U:/9SM@5[c6(Ydd100.?YXT&BEP+XT9,9Wb8\WHd=:(,9ADU_
]?fT&MA04H8O#HD&3)FP^W(,QgT]-O,=UNMdAb/3QeMEBFgKD=4Z(O1dW7?02T1g
^<4EC^Yd=gQ3<9I.S:TPCQdfP;OB-OF^JOd1^Nef]T>EL_MD8GU_NR@NOd+a:=A0
/WVZ:-(G:f8.7/,7@#Ld5a,3Q8B^?Xc3N+c]KgdWSO44F:f+5\GbK:NY\6JG^U7-
O7NX]HL?C4P:2@f?E:DZ,2c0J&b=Q->B-WNR1P>(J)8?K(cOHTJ.N3QNFc7CM/Sb
AOOX[)4IYT=FJW@EB3Z]>V[O^c8<=@SFD#RYd.JA\cBK=[&_4/:2e37P[>RY0N9Z
c.>CEL[2;L-IA73&H[BZW_DZ<bW#\YOPDJD]#>5EV\7\M,_:fTQ#W^:/TI1c&MKR
=+@#:P7+D\]1?IL/6]-I&P:3_NPcU\WPNX@Cd5WNP-[=:-E:?:HE/GgTB9,-P_K.
<S;#[DAP7:@XA#8;UFV>9e_gdIT:@GV4S2J5JP(^#+:MX@,MSOHD+C#g0NMTO6c+
Q88_/Of_83S<ZLK0#,)<d+I89-OT:^L3aT9=+LEK::>MddD=>W\-AKc8XBM.WN,/
CKY)IXDRH<=eDHVdeXf[R=>F8=].D/3?)=CA99Y3C4\(_4(&=T)]=dC8^fW=b^U\
))W4V>:VNPG=3KGTcg07@fFLV5[&;UINd3R+X0C2@=<+LD\&>[+f[e9?Ag#:-dE(
PVEb5f3W9Ld5=7cUHP@.;fHMgU400FN7<G8:P]]4P],\;4#@I]]aLDc5W6<gb1M^
ICCWAeN;N=Ig(cTO3f\3#;CcF9Fe=]^33327Vg]ZZ58Bg[4?8&80dSW/DX,0-05;
HC/>cE15>+GW&F8U<M1?F+c^6>Ffa+4ZB65ADHU8&[B_<N^K_F^E]^RBF(17>)eR
&:#N&G<+>,H0@Tb\]TD)C\<^c.cN(>c[1BH).C>2^,75/Xd8O@>M6AIDW>b;eaWG
+b.TI16aF(/#R0_\?J>-EK>/d>S33b0&:ZN5>DQXQE&<\.&BL63Q<g?Y(L3b_c>g
9O;PVg17<B/-B:eNVY<.WWH5d7(_,KWeR^,@+c30^Ud71;Xe@DcE+IU#^H&.KQ]b
bc,6:cgJ2FG0;5K9\1@[J_->X83/NJI\Z+UG-\@FQR/I-LJ)LV@gKW8Z8d&dMSTG
Y)@;a7?EDf_#cMe5\PA@a<V@EL7HPebS]783U^MXK@f[Ig]UM-A-(0#f@Y2E/:U<
:DVUN9HC[8G6Z,gg)UbO8TUQ4ePMceM0c;cJd]4.P:F0R6HOH76<FY,,#X8@O-:X
]\/b])85-Y6AS>7@S6_>_P_<9<]5NLa=U7I:;a0]:&)4a_)IHIZ6-ZYMQS5f:RaI
e_4AbJ06()b2UO#,],;I4]:Y2UVTfd:.bJ:7,+:a\_YQ:c]@+8,LgF6.]b8f(+LO
^BB-SKf95(TXM=H++)HFJAE5Lc<PEF=eRe@93D35ga6--dQL\-)\,P[/WF2?+YK+
K5@f-0-70.#_8dC=3;C53@XCTW(?51fG@LTR;U#6/TT65)L/bM@;XKH]^c.2L1?S
^&4De2-</Q^>CX.;\b13_+JF<2RIS1\Yb@GUUI9#,\P]\B[5BLAN43XGX>Q59N@R
DOCL1/^92RLfT=95-]A/a<MZ1?E//GU(g<<O(0Q&M#<P.)GX#NEUE:9LdY=6<-^B
f6,0/B2X1@Tg\+6\aY4YVHS+/>=Y+-YF:^K_O^QgGe]SM;T1LJf0^aZ?685&F,)P
Y(.WNb3]@KM0,)J6746&S=?>[0bI:SUcRGdBNNNE5E6)a6U>5(eYe,8H;6:;(\OP
J0WeOIV.@aNS<,5fEF+YA+D3.:D[U9R.cN.4Bc2R&H#D.;];KVQ=C9G54P/<F9FV
TC(4JP;bL,:?[CL8Kc&@3.UR+PJ?J_]IL-).ZSDN<)d_&F2e\WGA[Ad[2I5]0_08
4beX;[8C;e0dYMWP-M0NSP3e@LDCRFZMNSc.N0PM+3P?ENKdB]ELeGe5f-=]?@9W
JA^+gRaLY16NB@0P^2&^e[gSCF-7\03Z3Y@^??cC))DU\#4g=+VfbG:2J7aZ1cYJ
68O0Pf9+bA@@X6?GF+&CRJ@(=b:,LOF?D^a,,[a+H]V-]6R#N.3EBFW+([-BOC70
DL&KK;5^6e,]ecH5d#f&OYBF9a7)?AU/4MfE2;FO?I\c1GJN_9Bd<K5(]@(Ub^#b
MS-Yg2aJ^G9PKZA2\@AZZ;e)>F?La&JZ(^,=VgG=cA2,C-9)/Q\611T831eUUW);
\0\(C3>eZ&Cb_;&N+9KfKc009U0eQe#)A7)a[C:O#XK=/]V\B@dA>I;ZEJ^1c>Cg
C/&)M<=&[#]9A:AJSdS,_Oc@6\A=TbBMCa__EZES2><_[F=eB;=RBN.f^^[K@OfS
f+9f3WMWEZU__4_&(V,^B76^(.f4>SW4a8IE\b@V;g]/3BdJ,<A1e86);,9f^,Mc
,edL,51JTcDC2.R]D3&JV/&ZQbZ,+R?A18Y&1C)H9AH=gC-;]/CFV:WIPA0,&[;-
ZRa>f^.:;gEZ9eF)fX\f[81a0]6fNL+P#)W>MWf<<J-+TM.T?/f6_NI:V.C.=>9H
YbEJ/)G^(9\2V:6-/<PAWPDOB[6(,E_2]8^[F/bCZ,P,+C=:;c)UGADdFbSWYbgG
T:,M\IIP5fJaN+3KG^2.#UP-EPT7<@XUe5_+-Z,>9=+.4A\J31c^_b>N+P;<XSS\
]573E4:@FgNH^1_VOc]<U#;^Y]<9ag6=X@@@B\R9VUR)/9&bL,WaM]N[RK?e,V-M
=8.=LLO^K0M;DP?#QfNb^U-_NR8@Zg_3<&6:BTBLgbSD,S8TR)3aPS<db0PM^7I;
.#>/<&D>^VM;:V=:&CcHZO+F]W&T52d(/g58:cCQGfU1J]Ab]:+JY&XAD]&:O/IV
+@D?=W6+fcS40ZD\@3>Q)78LU)\#U:=17/K\G3DUO>>H,LFJ1:D)R:5A[Y#+1L:b
XM?RXYT8Q9YAe+aL]_(JRKZ;Q0]Dd(Ac#;OVSbcLXD^I8Yb;5]W^3Jca]:?QGG08
9.7-b?P\(1&bWJU^bM>=\YJW6>c1Vc<=43,f<9eCL++Q#LXOWI\fMA@<.^:8V=dB
:B;;7.We:D:_+fGUUA;HL6A^RB]RE7;7XRJ+=,X6_X3;XM;5S+4.:-A)].OGfG;I
P4EDfH@WO/TMfO.Z<I5O3X?_MH#G5Y.57RcEO?85_g5.aP:LQcgF+9/RI>;,0FR0
Cc<C_bWdM@.3CAZ-EU8@KU^2CF-NNTHC^-BD65d.S]BHCTUQ/ZF2)2(U)]Uf#S#H
(Wg2;BP=0AFNYe?CS4FDN;</Q8<XY>AX<gSK/[:\YD;S6[cNM=dKJEM<F8_;7;Pa
03ZMMT8Y^&J55Y8;/bS;#5&<?T0)/KI.V(Z]Q.:DDT40g_K/<e<JKYfG=faF8]QD
AGH^LLG5M17+IS#e\_7,I-:JA/eQ&1d@4N^eZ0)O]XUZ0-LR.IT@M@W^C0PO2C\-
9ZR79[Ia96bgZDQ.IVGEJ\^D3MB?I;GZ;9AM^AG+92V7W(+6=#QeBTGbf&WX6KAb
JaW@SZ/.>:Z?d:FE8HHQH?,0>(c>aGc<5e\^(I5-QUC>cV,H9RZ]@^1b/#d=?S36
Q/WW5O@:\FQPO=#MV=IK;e\P:cNLXa5G0^S5>VEbe1+&#(J-5)VV]7=Zc\/-)S1I
AOWA7M==_,b6=4-:.1JY4H#dU&LXJNL_QYC<8Pg,0)dAeXJFDNaZ@8e,<+I(9Zbb
44D4Je4,\PW(0>;T=(S2D7-)g4e#_S+ESdg)ZA0CHZI8O&JFHHWb7)RE8P>G1+[X
UC1^CfB(U#Lc&Y&ZBZ:/UT6a.Z_\_<R>3:#6f?MYG\-:9M@9XIVCF#-O6<_RdQ,B
NC5EJaY=V_)2Y\/TCLZbZVb#bd-6KRCK1Hd0BV29/-QD?EAd[&__3[fSc0^R+4R1
W6;6P\<V_XO7E@]16:<caW64Pa]^O^2(3ZZ@\L->.^?_a4TB,,]&e]21#H-#B^SM
DUA?PXLTX@/d:AJRR5@?:;ZKL2T7\/T8][79W=1)V1E;RHc0++d;HB\D>WQ,O)FO
Hg)b81UaK=M-9Y6Y4\@.[-@W/CcX\gWSV[eA3>QH^89McQU4;_GFIK)2(#IUGYeT
#^T/Z8Hac/NW#<+:]fVO^-&=4VSZRPD_JTMd5YOeWM^W7MN#SUB)).W,\bP@YPT2
[SD7b=XMV_e/.E=.Bf=97F<;TW18LV8C(L4Wa1I43BT6X,ZBV=GK=Rg>+P(KMIf^
:J4cIQ&]K#6c8@e86KT6BTfd@\N0cY<)H_/f/a.[ONZ>AAFQ]G@-a(X)4\@/\S@-
[CG1SEC@^b?S=OBOb^[^XJ\PGU]fF(L<;HTIEBeD,_Sa\Z;#,2R(gZR^T4]D4@T;
^(agbeTW;9Oa,<[UKXBYQFQa?6HeACc(Md3TH]c,FXb[B=-?H3VBZW[_L2HPeO@6
4G&U7Vf5],dGf)L=)&O58/@EPfQQY6\DRNf4<=Xe]eK]SecKbIY#Y:49H:4^24=N
_a9#QCYCcGK2<D988JV>0YO-<U@#>H25:<70U/(/+?D>C.J7J#XA])\2:+^OL>/]
&YHU-cR-?SMW8cV-:^Cb@8I]gX4@B7Yc^H./f99ENHI+ag>.,^]/;N@B/A;4OE9a
)OWMbb?I3Q7DRVB^&P_M9NK3Qed:HZ8<a2YEQ5+/C5A[U<+31ZggL8\V,FYga]9[
W2EDAH&O?.G]a\71)15)Df-&a,aX2UD6)FF7Y@QbFf^VXT^:(F\Z1\O(2^;3ZD&D
cUcJ@Bg.d9KOFG?(:J_7@7PRP)_R(3#([I<2454D>1bMe+eWW/GEH6Va;XOb0IcG
.ZY0>DT)2L;4=McZ&43E:RGQK>[QeT[E)LP?0X417=RF29TGA\(=(3VSS(A&,[eP
0:c.>gRD+eHD=7ZYcU#@Le.BVCS+_f=UJNG23F:SVY&Ue1OPUAMYTK04>0\5#+T+
Q6L5^Pg0ZIG&._F&#.2=KS#96^#IC:WgaXgG0XNF3L]R,bH(eJ58ceGeSE.4OMZS
]8M#I-7V<HG6;#(?0\&>W[)#8VELf#W8W-6>X(XE8.-d]44C0:-86X-eaJbXP(Lc
UDD#MDK\@9b=U.:Z7)f?OK/HEKV6&LAKP)N3>?Q3K41-I+B\8=0P]+[cWY/\dH(b
R<PQ\67GdHVC6FT>VPW&7N\L1^:RS(Wf(G5^.O.;b&8=G&K7d2WUeR\AVV>\Z=+/
fe[3K5]0cgE3N8@E7?TDAF)ab;X3?b?Q,[<Cbe/KU6V?f6a42C^79O2,,/Ye\R[T
L@EV)0BM0>dB;g)]QA6d7?W=U:DYLH0a^JP/=2RFaPJ62R:+?]4La5#Q#W+@_6W9
QY\KJb>/)P>5RJ9NI&^K,dG,9L\>LNQLV:&/KN\\F&6MBW6SFP+?)^8/BTDe4_gI
M5f.B/bJ4c<R1I6>)==+HKK=(+3G=deX9[;L2,YO4fIO&?ZGe&Hg1U,0N-2QUO07
0,(,:.@:>9VT?3UX:NFY3aOIV2T:.S>TBE5]TJR::E(H^](J.O;]KKCUY\(cSXeg
M7#>K:,,]&MN68??PgC6@L3<W71M>W;]cP_YCEL1,a.bHY;EAe-g@WaYO2?DL<-2
M>M_:DR&N-4Y5ef7g,4DQ@.1)_FdS:Z[4.WM[E?EBC>TH8KcA=#=8YL]cB^/(NaX
K><&@Y6&gc@>E11Z5a0],Zc<#B^@/8YB[_(8^7U9f_7I3:(O##cF/_NeB]R2Cd^a
e2aX.5fE7W62?Sde/29)4BM[Ob_\R<>24K:=FJW)VM0deJRA@@(/Kd.13U2W=M@8
<N9IV)8fe+F\DC:LGbQbXH?_<VT&fU_OY+1)QEJH;3YI3.<g.g5W:R&GK/Ig9N.-
&:a@?dP\#?H83aB81)&cNgQ]bZ+7L7RIHONGF<V@.La4-3,8M#0,g8TR(\JT0^Aa
ae79C#e4#G?/]3V,15BMC_NJ\@4O.MD>[#)e:O(?G7fgc46>DC9EDcYPeS\.#CCA
H4Pb2Wd[<Q5H4]d5=>Q/E2V;\(aK3a=@X/.9L-^1RAG6H;[FP<bZcfO@6<,c+<0U
37deFB,9@.O&15UbZF6gCOF;]^^WG71,S5-W>@83B]0MB&L[BU4LO\E,OdG,OeM7
Q@D7V/<QbQIdL10#::RR6HFR8EW+AC2,YL.M>:NQ75S[\J\bQ/7WE6M2K0=46&3A
eE=+KZ4F0^+OI<f@DJ9M,>cWS<90W+cLMBJc19NW0gZgAJNVb<^^35GNeS+?D?\:
c^/8[HDXYX)ZD,82F/I/+)@2+c7\?[EK#Y(>L5Q:PA\HX]GXWcc1?EUde097=\(B
J2;N[[d;ffQV2I@\A#CQcdU1K[7:5]-P-6A.2^5@,=:B0GMM2EU#:3XX=9?;e[])
-KaDHA[JW9aB-B,H+dC:fM3QAQg(=]KA5Q0Y6P&d5/;(eR@Q/G)bW<Jf5<:)W<EI
D;TL\g?B[L.?UePcTF]:I<XL&PBN&Zc?=d#Q0BFF7:5,TE^1U6HbF.ff2]#5\6#=
Z<,N80\+EHada_a/f<0D_GCDTYA,IW(A1M5Z5aMS)\=E,;4@UA\@7.5+&BZdcICa
3+&:?0,5G&\M2ba_6?9UU1-(#;842]O<dG#TJQEK2:&f=A<#AHC&g.=QeOa,K8,#
,@IUMQ[YbW>dUEJWN<c&<NZL>.>-2M51dMD3@N+2K5YNP1G:Dg1D7gE,IY)<@YZ8
(UUXS0?B-VgeBGDTY#=7\bB1e85^FXBSQH[8G_+bJGb3d+dS]&SZJD(8>;BI(Cc5
R>Fd@XF)\6fN:cf>95RL_X?c4/[gAI3:J];OY1;Bc3)65#/WLd>3V<O9:TTGb>6G
,T1\0a^H&M+,XM^cCESM&N/@R@dA,_RC9E4g[YYbN<WXG<X9=ITB^XKZ>dL]>)-)
EJ-JVL3F/<T]1J=>Id/dJBS0EH+d_<I_^EH0dUQRGAR</,OU;C+SU4Kd)I=.dE0&
HY,V-6J_2bU2Jd1D#bB+@&7(K,1:);cF=+@QIb[bYcF;EPER_@=-e;?Z(UJ,^5FM
,DM#W8]KH?JI4YOW^9DAH^:e6&e#/N2AQeHET)19DE<&;3,PWCN;2N[7_0+4=cL[
MT[C]2,2X:I4a^a..3K2FHL]4&^XO<UN2PUfO+XFTF8\;>LcHdaWg5)6SS2G<2Z8
9OKT7J=G8Oa2#L-O^3Q:AGPHfJ9W:WIfa.0WLY8)^NfW2de\dOe@cKKe2ZEB.G3V
:3OGK;Dcf+&YY(56\e2JM/\gRdS,fX51Q0E+O(\PQ^8Y:]LV(9_3&Z<1e\H1IPR3
9CEMJ:S#X<W-gaN@MYEG@_@NCfa-FIG,YWO(Gc.<+47/6fYT3](cIK8/.RL1Y]=/
KOI2c]XRASP:-dfRYG3JRBD=U8K^1@F/_N0.BKZb5WOf#+aFPSaNSUJSg)0TM8;6
ZJe]U_H<(1=94d2QTTD^/^-Z0T?6AV.O#_U=-NQ\M\G5X;X9ae=VUNF@W@]?J#J>
[8;(M=Za3U]33ea]_]QMH/a_1I6E_SDS)A.1FKD5L>[#_:L[(Q#?9S58]f99LXQN
Aa-RRZ3eb=O,EeV@HS(]\/,A\^.J7Z;3B^G+d,_IX&>(@f=?L=MC+BF?8?,0[FQa
IC9_aUSMCT>GDEe,Gcc0cZ[@DXN]ANQCNV\<QQLV3gNFM^TSS4YdQ_d<V=YF.Q<)
>UbR#9#L.?fcD=^,+.&aT1N<J&7C:)&G\A2NC8/IN1I^_dTfD@PLB/a8]8:[?=;@
C6KZ0EPWX:1XQ(Y#@8Q662>^QS??MbQ3I8cROZF1[MM<H\Ee)&P2[J5#^cRdgDV]
H@=G1SIO[;.A/PFGK?RM920YFE,B?>=?a/=e>I21B<TGI=7OVdLVP2A;49]Ed,+Q
b3@ZH&&8KIg_.(6DOO(3d8[W3=[34-SXV:1&T0[,,f,XdH2+5-_GR/O\?]M:Z#=9
H>Ka^_,F4DHG?6IIV4IB19X#UG22Y(([QARc>M2T5_T/\MIZ#TIKd:4([eQCaFJ)
&;M&=57U>C<0NJ-ZI[151?F7O[19LK+O-+_+X\G?;5;<,)effO2<&K80C]aB.@f]
A/1:Mc]UG(IQJ>c0IL[,Zgc;gR^S[:>]I:@BK>XL(WKEA/Re0_5dI\WVV;dW68Z.
8].;_.JE=&eM;:;S[[BX=JS6\aF=[58#_5YdU3R_P4eRbc<Qf4DL-IPc472DVeK[
1ZM)X/IT2UgTFTc5B&,7?e+JM6/M23?b9XVGP23Pb342X5/X+dC9,RAG[B/N8G:8
[2[UAU1FL]aRXFZ(]ST-RU9M^bNZ[W0O/de58(-(+KAX?2d>N5Hc_JVI5<[KZc41
P9XXHWT:G;?Tb[a=B[fZ(2O(b@6PI;T2G&2WfU&/:Dc)dX5ZFB#JL4C[P3PSc45R
XXRef6ZM8@X\=g0Kc&K4:<3VCBOC;:DU6DHC//Pe[=AA5UJJ-IC_G(#c,H&?&K,J
d++KZ[.S>JCZ0K&USI@A-^Keg9?<]2^2XeT^+C58T6K2J7>JH:,C4gWR,acH_.Ce
FYUP#dR9T3RAb\?]-:J8.WbHd0EQJA3-PN#^Y..fK]>8@:F./+2aQ1#b8CBZE\_W
YUe>EN?\9S]AW=P-]]CI;S)+8?Y_)I:Cf#/\(\<g]EUb4R96A;KUW>QH:@ac=F-:
9D4EP9B6_EB:HNS4H7cbGUb<:NYd_,<-GOg#fY+gLa=?TABI)_7R1Og0(=Hc/.2.
R)dCS(?@8OS2dOLc<<0fUKgF6<H.@)S<5BMgRB,JWd0S=]K_SCXD#<eO7(cW80_A
PEUU)@@S&f>S-YZf-SZ3/+-90>?QN+TO_f\J.[cC4CQFRPVP^I01\JR-.3+UKW>2
H6gc4G3Af4IS,$
`endprotected


`endif // GUARD_SVT_AXI_MASTER_AGENT_CMD_SV
