
`ifndef GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV
`define GUARD_SVT_ATB_SYSTEM_CONFIGURATION_SV

`include "svt_atb_defines.svi"

typedef class svt_atb_port_configuration;


/**
    System configuration class contains configuration information which is
    applicable across the entire ATB system. User can specify the system level
    configuration parameters through this class. User needs to provide the
    system configuration to the system subenv from the environment or the
    testcase. The system configuration mainly specifies: 
    - number of master & slave components in the system component
    - port configurations for master and slave components
    - virtual top level ATB interface 
    - address map 
    - timeout values
    .
  */
class svt_atb_system_configuration extends svt_configuration;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  /** Custom type definition for virtual ATB interface */
`ifndef __SVDOC__
  typedef virtual svt_atb_if ATB_IF;
`endif // __SVDOC__


  // ****************************************************************************
  // Public Data
  // ****************************************************************************

`ifndef __SVDOC__
  /** Modport providing the system view of the bus */
  ATB_IF atb_if;
`endif

  /**
    @grouphdr atb_generic_sys_config Generic configuration parameters
    This group contains generic attributes
    */

  /**
    @grouphdr atb_clock Clock
    This group contains attributes related to clock
    */

  /**
    @grouphdr atb_master_slave_config Master and slave port configuration
    This group contains attributes which are used to configure master and slave ports within the system
    */

  /**
    @grouphdr interconnect_config Interconnect model configuration
    This group contains attributes which are used to configure Interconnect model
    */

  /**
    @grouphdr atb_addr_map Address map
    This group contains attributes and methods which are used to configure address map
    */

  /**
    @grouphdr atb_timeout Timeout values for ATB
    This group contains attributes which are used to configure timeout values for ATB signals and transactions
    */

  /**
    @grouphdr ace_timeout Timeout values for ACE
    This group contains attributes which are used to configure timeout values for ACE signals. Please also refer to group @groupref atb_timeout for ATB timeout attributes.
    */

  /**
    @grouphdr atb_system_coverage_protocol_checks Coverage and protocol checks related configuration parameters
    This group contains attributes which are used to enable and disable system level coverage and protocol checks
    */

  /**
    * @groupname atb_generic_sys_config
    * An id that is automatically assigned to this configuration based on the
    * instance number in the svt_atb_system_configuration array in
    * svt_amba_system_cofniguration class.  Applicable when a system is created
    * using svt_amba_system_configuration and there are multiple atb systems 
    * This property must not be assigned by the user
    */ 
  int system_id = 0;

  /** 
    * @groupname atb_clock
    * This parameter indicates whether a common clock should be used
    * for all the components in the system or not.
    * When set, a common clock supplied to the top level interface 
    * is used for all the masters, slaves and interconnect in 
    * the system. This mode is to be used if all components are
    * expected to run at the same frequency.
    * When not set, the user needs to supply a clock for each of the
    * port level interfaces. This mode is useful when some components
    * need to run at a different clock frequency from other
    * components in the system.
    */
  bit common_clock_mode = 1;

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * Enables the Multi-Stream Scenario Generator
   * Configuration type: Static
   */
  bit ms_scenario_gen_enable = 0;

  /** 
   * The number of scenarios that the multi-stream generator should create.
   * Configuration type: Static
   */
  int stop_after_n_scenarios = -1;

  /** 
   * The number of instances that the multi-stream generators should create
   * Configuration type: Static
   */
  int stop_after_n_insts = -1;
`endif

`ifndef SVT_VMM_TECHNOLOGY
  /** 
    * @groupname atb_generic_sys_config
    * Enables raising and dropping of objections in the driver based on the number
    * of outstanding transactions. The VIP will raise an objection when it
    * receives a transaction in the input port of the driver and will drop the
    * objection when the transaction completes. If unset, the driver will not
    * raise any objection and complete control of objections is with the user. By
    * default, the configuration member is set, which means by default, VIP will
    * raise and drop objections.
    */
  bit manage_objections_enable = 1;
`endif

  /** 
    * @groupname interconnect_config
    * Determines if a VIP interconnect should be instantiated
    */
  bit use_interconnect = 0;

  /**
    * @groupname atb_system_coverage_protocol_checks
    * Enables system monitor and system level protocol checks
    */
  bit system_monitor_enable = 0;


`ifdef SVT_UVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to UVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to UVM_HIGH or below.
    */
  bit display_summary_report = 0;
`elsif SVT_OVM_TECHNOLOGY
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to OVM_MEDIUM or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to OVM_HIGH or below.
    */
  bit display_summary_report = 0;
`else
  /**
    * @groupname atb_generic_sys_config
    * Controls display of summary report of transactions by the system monitor
    * Applicable when #system_monitor_enable is set
    *
    * When set, summary report of transactions are printed by the system monitor
    * when verbosity is set to NOTE or below.
    *
    * When unset, summary report of transactions are printed by the system
    * monitor when verbosity is set to DEBUG or below. 
    */
  bit display_summary_report = 0;
`endif


  //----------------------------------------------------------------------------
  /** Randomizable variables */
  // ---------------------------------------------------------------------------

  /** 
    * @groupname atb_master_slave_config
    * Number of masters in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_MASTERS
    * - Configuration type: Static 
    * .
    */
  rand int num_masters;

  /** 
    * @groupname atb_master_slave_config
    * Number of slaves in the system 
    * - Min value: 1
    * - Max value: \`SVT_ATB_MAX_NUM_SLAVES
    * - Configuration type: Static
    * .
    */
  rand int num_slaves;

  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the masters in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_masters.
   */
  rand svt_atb_port_configuration master_cfg[];


  /** 
    * @groupname atb_master_slave_config
    * Array holding the configuration of all the slaves in the system.
    * Size of the array is equal to svt_atb_system_configuration::num_slaves.
    */
  rand svt_atb_port_configuration slave_cfg[];

  /**
    * @groupname interconnect_config
    * Interconnect configuration
    */
  //rand svt_atb_interconnect_configuration ic_cfg;


  /**
   * @groupname atb_timeout
   * Bus inactivity is defined as the time when ATB interface remains idle.
   * A timer is started if such a condition occurs. The timer is incremented
   * by 1 every clock and is reset when there is activity on the interface.
   * If the number of clock cycles exceeds this value, an error is reported.
   * If this value is set to 0, the timer is not started.
   *
   * Configuration type: Dynamic 
   */
  int bus_inactivity_timeout = `SVT_ATB_BUS_INACTIVITY_TIMEOUT;

  /** @cond PRIVATE */


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
 
  /**
   *  Stores the Log base 2(\`SVT_ATB_MAX_NUM_MASTERS),Used in constraints
   */
  protected int log_base_2_max_num_masters = 0;
  /** @endcond */

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZH7+2D9L3j6EXF7VCpAE+nsHEetQdd1Eti4CgoqXvAOmcEKcsUWDG2B1wr4i7UBf
lt+UtyvriPKr1Uy+2HP52drCi8+h+F2NFEsTJJpvIi2+FW399MRVooCVIzu3CP2a
1I3LHEnNrPOkUKlsVCE7FgmHfX/EoAoWElwLkJOqhG79Sb61ilFMNg==
//pragma protect end_key_block
//pragma protect digest_block
Dh2MBxDTPrPlGpBvawALiyHptOo=
//pragma protect end_digest_block
//pragma protect data_block
MF6GbKSK29E0ncUPF1CVTqFr56yQrJE3pMEoMK1FuNOrKIweGY4mRWmIrfUQXvTZ
dz8e7w+T+nyQ18P3qYHrIPoYhAsdfAt6254+QI4k6EbT6urM1qIP2eWa9aqjHrBV
kymf2rP5BpMMp5mM7iKyb0pPt2iQ25XcC+O8fyF2SkgAS3iGKlTkLWqy0Hd6HtM8
LVIl6aP4WXaOysDocw4n4EzFGY9Ncin2f4qAOcGk8i6jabQXfKMCIKSn0MnQt3UI
f7SOebJPP6KAF3SFArU/FSwP+rGQqnru0Hqfk54Qsf64EZMCRMIC8OU3Y/UX4pr1
Vtsi8yNbzbozd2U+MZZfomzW1UQzm0a1p5q7Xr7gTpK3AyX8LVgj+8g3WG4XpSdb
TBxn7iThKpP67Vn1s3clGtxSGBeEVNlE8hdmWFiFwoVoFKYly5XudvUHewWyhvjM
2yWmftcfbXFdicVMdVJYzvKthdI2tfrKtupJ446JUv6HajLUdiIqL06Ndoy82MNv
twttTLgubBFFHEhmBRDZS2rpyWDvBczrtXbAD6noJvt4ypCTLVBgquxyotwbGeoX
dZ6zaRXiGszpRP8pQ4lhJeUzycHJwIac5IabJenEU4AjjRZolT97kdv/eUlMIVsG
8BSbwrjZXfHG/OcDyuyYL6uMKpohUUgz/yA+SHFl1DJBmoBB/8hyUN7Oz/c/iYkq
25jNR/KwNNRapzzGlFBTmWCE+C+WSJ3W3NtIIZZaJAXLaw4sE6h49BYnUgqONU3N
1yS2eyv30v81btc0j44cwWWUT1ANIvQqILVLTFSCHTxxSzPT7KruTwNwFB2RYudJ
CUxqErFL+p1LipHGOpq5LMwEjqbI/zUsoklXNN9HpBu3h25nI8Znt7rnWRBmNTtq
plSAQhSQcehnMcoR7JKOAqDbFYVqsMRH3kZCqD5Fk6YUgAbLdFmT2KA2ZCbJmDya
6mm5Hjc/Ep5obU4M2Y21eRkaPwZJ9qTmp88o6D0Q3+R51j/FC+jIA3TsyJnPDtwj
j5B6Y5CQMkbQkU70BN4vWTg003tWwJvGBMog4F7iEJHHcNk2vZBC1SvKhMMFFDoh
U7XNV0zXHEZ2vE87mpSCLPyY2FYhd6PIiF0khWR0cjn9274eoLDCOsJ/+JfL6cnM
PMkCW2NCEgq2HxypTkHS5ukFsBCqDmT6FKMZXxwULedyAv33ssjJsHXgxlvfdPcc
fCs9sfsDvBdjmhdqSYUol7TJTMjBcDALr45+sb859xE4S5B8ATzZlIkVcUCBT7M9
hO8HiUkuivVctKo9jEBbVJIj9uqHF7Be2zqD0T9vBjR3UiuuPbT6eb7F+ne9tGnP
+0XOu0eM29e4MuFplVA1RLZwxYFnMIpwP85a/Sct+AYvfK9j+CP1HnuctExPpHK5
N2955ILxNf9bEmcO6eTCt+g/kEeu6lkpBByrGVm3oVOAPLWjiJVbmWzuVaykh/Me
YGeBQ9blQFFmncgKS+kpTCFHDtP2aVYjdwOkReI5pScikRwemoKkXYf2T3Qi3g2Y
NCZkLtsds8NBWTWiABpxk0b3wF6WCWa0uCBioEAFO0Uf+sJSeAMKz4hJtoeibiJb
6/ZFx+ggOCxwjHq8Ya/50Frrr8Cjdd7ck3kYj4Gyga8A6IkxWdQV/9d1998sOXoc
AGpq8c4yhCXdS/f9SbaVKNeWUeZONSfycd3XilHVI+2U027VdkLz/YsWwAFVzJMD
ojCgvmjzIE74F/KBnlyxSBXAMhdY9PZHW8Q1TnkIA8tM1B9lG8QFJV2R4kf/5E7X
f9lwq2mv9zFHcHw/ew0weuIpUq5EQGOsg6YjTDSXtAb9BF7x4im5ckU7RcwhHXUg
ktTG1F54JfO0isQJOpA75pUsuVBzz14t2PdDSYqkGlRhZjK3xGBGmdVUXH/jVyuV
YJwbd/0R8JHJ5C5MXii3KmdZN7AzbbcFAREa4y+LcKV+EpIqcrGKKfs8tCIp8uoF
NLeRsfCmgreAKmAq8UNXDkBF0QIpjIgSshR7Z8e62IPT5rAUPFbEtVvAVclgDgt2
5ZcUmr5LFc3wBd311TkJ0o+YzAo+HwMX2GJMUAFRakvT2QUdzgXV8Y+rOT73fKuT
vQnmF4Ev16xmWYF7yS7v+1Od8WsgHceonLMEn29cLGCUDTC32OffNAExjHDr6Mz8
/jlKT5dE8delo//LC/ZOlfazsXwkny8t3EXGy+9Q2u6xjGSaHqZfML22pldKk4fQ
k83vz16uNwOPqQeQCElnEql23wa9wpTyO/jdYWlDMVQN0laKbdE1rAmpB+sgPKA+
vQriOFfBu5An9//cTh2VBJV7dkymRFcXEDWqmoRh0ra6fKi3CdqGtiY98Ma8yIpo
C08O1I8J/jS7Aa/t2agBoPmRp/6GSxsMtn1MbecrE33Gx0AeZiJAOxeRZUAT5aAF
rL5eCNxBD+3w7ErOkrgKJlHUI3nNxTjqpa9+m1arD4Th97HhNVB6u3WOlEXH2y0K
yWxjgiwV61jMwFnZTv2frKCVy6iNggn7JBRlSRf2JaTYwACI98okdujIkEKS81ws
R7g9TTFkMDfVv8kry1Cc03lxA3FuJJn39imdIz7bsFXV4rakXE4mJuZwwm0dX+BL
mrLxjbw3LYTcniUWbBbCWIYyz8YcgHSp66pQWgf9xD+e/j2VRoO/YU/Yxed0jk3i
UeRHJLztN935vTPUupX6Jr3zd5c5nFtLidFApcnk0BO1Ogoa0VAoHpiVUiOE/Kys
Im4PEswXj1qTSvwgVwfZ2fatZZhDYcDDs8QkQHT1yLAzBRvB7qM6gAsFLoWeGuTI
rBJUUXmn+NlCX5Ys1+iAOfVFwCFrBb1C4l6b5dYgq9nrfcseg0XCIGjWbf3c4MXd
MklQp21dPH40GTm9CpF4d3ZsY4rjk+YCPZJ83k/tuHKKEysdfn2YwT3PNCGDIZmY
thte7wjtus5d8/LRga741xj9O9HUb1ieqVlSTJnc09Q=
//pragma protect end_data_block
//pragma protect digest_block
KEQRlit5/7SwBF77b2ejNMdH2No=
//pragma protect end_digest_block
//pragma protect end_protected

`ifdef SVT_UVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`elsif SVT_OVM_TECHNOLOGY
  //----------------------------------------------------------------------------
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param name Instance name of the configuration
    */
  extern function new (string name = "svt_atb_system_configuration", ATB_IF atb_if=null);
`else
  /**
    * CONSTUCTOR: Create a new configuration instance, passing the appropriate
    * argument values to the parent class.
    *
    * @param log Instance name of the log. 
    */
`svt_vmm_data_new(svt_atb_system_configuration)
  extern function new (vmm_log log = null, ATB_IF atb_if=null);
`endif

  //----------------------------------------------------------------------------
  /**
   * pre_randomize does the following
   * 1) calculate the log_2 of \`SVT_ATB_MAX_NUM_MASTERS
   */
  extern function void pre_randomize ();
  // ***************************************************************************
  //   SVT shorthand macros 
  // ***************************************************************************
  `svt_data_member_begin(svt_atb_system_configuration)
    `svt_field_int         (system_id,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (common_clock_mode       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`ifdef SVT_VMM_TECHNOLOGY
    `svt_field_int         (ms_scenario_gen_enable  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_BIN)
    `svt_field_int         (stop_after_n_scenarios  ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
    `svt_field_int         (stop_after_n_insts      ,`SVT_ALL_ON|`SVT_NOCOPY|`SVT_DEC)
`endif
    `svt_field_int         (num_masters             ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (num_slaves              ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (use_interconnect       ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (system_monitor_enable  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_int         (display_summary_report,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
    `svt_field_array_object(master_cfg              ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_array_object(slave_cfg               ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    //`svt_field_object      (ic_cfg                  ,`SVT_NOCOPY|`SVT_DEEP,`SVT_HOW_DEEP)
    `svt_field_int         (bus_inactivity_timeout  ,`SVT_NOCOPY|`SVT_DEC|`SVT_ALL_ON)
`ifndef SVT_VMM_TECHNOLOGY
    `svt_field_int         (manage_objections_enable       ,`SVT_NOCOPY|`SVT_BIN|`SVT_ALL_ON)
`endif
  `svt_data_member_end(svt_atb_system_configuration)

  //----------------------------------------------------------------------------
  /**
    * Returns the class name for the object used for logging.
    */
  extern function string get_mcd_class_name ();

  /** Ensures that if id_width is 0, it is consistent across all ports */
  extern function void post_randomize();
  /**
   * Assigns a system interface to this configuration.
   *
   * @param atb_if Interface for the ATB system
   */
  extern function void set_if(ATB_IF atb_if);
  //----------------------------------------------------------------------------
  /**
    * Allocates the master and slave configurations before a user sets the
    * parameters.  This function is to be called if (and before) the user sets
    * the configuration parameters by setting each parameter individually and
    * not by randomizing the system configuration. 
    */
  extern function void create_sub_cfgs(int num_masters = 1, int num_slaves = 1, int num_ic_master_ports = 0, int num_ic_slave_ports = 0);
  //----------------------------------------------------------------------------

`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the UVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(uvm_object rhs);

`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /** Extend the OVM copy routine to copy the virtual interface */
  extern virtual function void do_copy(ovm_object rhs);

`else
  //----------------------------------------------------------------------------
  /** Extend the VMM copy routine to copy the virtual interface */
  extern virtual function `SVT_DATA_BASE_TYPE do_copy(`SVT_DATA_BASE_TYPE to = null);

  // ---------------------------------------------------------------------------
  /**
    * Compares the object with to, based on the requested compare kind.
    * Differences are placed in diff.
    *
    * @param to vmm_data object to be compared against.  @param diff String
    * indicating the differences between this and to.  @param kind This int
    * indicates the type of compare to be attempted. Only supported kind value
    * is svt_data::COMPLETE, which results in comparisons of the non-static 
    * configuration members. All other kind values result in a return value of 
    * 1.
    */
  extern virtual function bit do_compare(vmm_data to, output string diff, input int kind = -1);

  /**
    * Returns the size (in bytes) required by the byte_pack operation based on
    * the requested byte_size kind.
    *
    * @param kind This int indicates the type of byte_size being requested.
    */
  extern virtual function int unsigned byte_size(int kind = -1);
  
  // ---------------------------------------------------------------------------
  /**
    * Packs the object into the bytes buffer, beginning at offset. based on the
    * requested byte_pack kind
    */
  extern virtual function int unsigned do_byte_pack (ref logic [7:0] bytes[], input int unsigned offset = 0, input int kind = -1 );

  // ---------------------------------------------------------------------------
  /**
    * Unpacks len bytes of the object from the bytes buffer, beginning at
    * offset, based on the requested byte_unpack kind.
    */
  extern virtual function int unsigned do_byte_unpack(const ref logic [7:0] bytes[], input int unsigned    offset = 0, input int len = -1, input int kind = -1);
`endif
  //----------------------------------------------------------------------------
  /** Used to turn static config param randomization on/off as a block. */
  extern virtual function int static_rand_mode ( bit on_off ); 
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the static configuration members of the object. */
  extern virtual function void copy_static_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /** Used to limit a copy to the dynamic configuration members of the object.*/
  extern virtual function void copy_dynamic_data ( `SVT_DATA_BASE_TYPE to );
  //----------------------------------------------------------------------------
  /**
    * Method to turn reasonable constraints on/off as a block.
    */
  extern virtual function int reasonable_constraint_mode ( bit on_off );

  /** Does a basic validation of this configuration object. */
  extern virtual function bit do_is_valid ( bit silent = 1, int kind = RELEVANT);
  // ---------------------------------------------------------------------------

  /** @cond PRIVATE */
  /**
    * HDL Support: For <i>read</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit get_prop_val(string prop_name, ref bit [1023:0] prop_val, input int array_ix, ref `SVT_DATA_TYPE data_obj);
  // ---------------------------------------------------------------------------
  /**
    * HDL Support: For <i>write</i> access to public configuration members of 
    * this class.
    */
  extern virtual function bit set_prop_val(string prop_name, bit [1023:0] prop_val, int array_ix);
  // ---------------------------------------------------------------------------
  `ifdef SVT_AMBA_INTERFACE_METHOD_DISABLE
  /**
   * Function set_master_common_clock_mode allows user to specify whether a master port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_master_common_clock_mode (bit mode, int idx);
  // ---------------------------------------------------------------------------
  /**
   * Function set_slave_common_clock_mode allows user to specify whether a slave port
   * interface should use a common clock, or a port specific clock.
   *
   * @param mode If set to 1, common clock mode is selected. In this case, the
   * common clock signal passed as argument to the interface, is used as clock.
   * This mode is useful when all ATB VIP components need to work on a single
   * clock. This is the default mode of operation. If set to 0, signal atclk is
   * used as clock. This mode is useful when individual ATB VIP components work
   * on a different clock.
   *
   * @param idx This argument specifies the master & slave port index to which
   * this mode needs to be applied. The master & slave port index starts from
   * 0.
   */
  extern function void set_slave_common_clock_mode (bit mode, int idx);
  `endif
  // ---------------------------------------------------------------------------
  /**
    * This method allocates a pattern containing svt_pattern_data instances for
    * all of the primitive configuration fields in the object. The 
    * svt_pattern_data::name is set to the corresponding field name, the 
    * svt_pattern_data::value is set to 0.
    *
    * @return An svt_pattern instance containing entries for all of the 
    * configuration fields.
    */
  extern virtual function svt_pattern allocate_pattern();


`ifdef SVT_UVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against UVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`elsif SVT_OVM_TECHNOLOGY
  // ---------------------------------------------------------------------------
  /**
   * This method returns the maximum packer bytes value required by the ATB SVT
   * suite. This is checked against OVM_MAX_PACKER_BYTES to make sure the specified
   * setting is sufficient for the ATB SVT suite.
   */
  extern virtual function int get_packer_max_bytes_required();
`endif
  /** @endcond */


`ifdef SVT_VMM_TECHNOLOGY
  `vmm_class_factory(svt_atb_system_configuration)
`endif   
endclass

// -----------------------------------------------------------------------------

/** 
System Configuration Class Utility methods definition.
*/
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gGm9OlF7mtFmPJ7CltTHERQSYsrWQO37QMWEOwZ29sLOh5NyE/lJF4+QVhMdFG1P
4yB78HqLtAOIurmy75LiD9O1N7kvfMCvL7JXKfISbZ7sxR351Kw+f+M3YkBb7LlS
OJWn/of8JyIP/TanVUshnI5XTzSrLwzBcio0/I+HrI0F8/H6pMtFvQ==
//pragma protect end_key_block
//pragma protect digest_block
1CmtZs5PyR3sTlTKoBUUZI8AsjA=
//pragma protect end_digest_block
//pragma protect data_block
n/F1J+WvYAJ1F04J7cLjC5hc46L/NfaXym5vBSux+ogWLKxB3csX1jzhApxFxc6r
d2NvRzzhQcq+AJBC2t09BPMH0dJadSX4CKg5xe+H5BtMSPiFojJ51fs1WQdOftXA
eElt0kyrjT6XJFjA0gh+QTU1wvVrq88Li8CRT0nPCUTaVLoZa1ZPClIPqAKTrTRJ
us3bQ6Ea5reWprcWnVRhInScByTG1dUr/9N+HLR6BiHI3qzPKQKXDff0Qnd6pD8a
npD9g+nqj+lD7EPghDW0NNfIjzGOp1F5t2PdOwh9mdKdniwgAaLRl6/jF/MGPeAo
AckZT9PYno9r7ZONdudyj7Oqi+V4fNajUgoDkxnagDy1FxZlewu7+07pX7d1D3Hk
O2YZ1OxZ3HmqDXQAdYSbLB3EKcQjl8vkADCWkfbsFLfpF6H0/LNg4uRGPbCisx0M
P7wieEUPEqnWfIzne5cQV61DNpXT6YsWQooWPmwGPwzayzfqmGgiFlF12WrR8yPc
57z+paiT83xeyc1+O0NqdKtcVezDIEi4mkEAzrpfGEsxe6/Gdj9F6LkqbTp5MUtE
UvP0iyqeCfbS817o3j52CoAc/PNQ0d760Irq1Ue/QPMskc1kSCbSr4FT/ZRctg/7
E3G0WnFjl+AyJJwDmC0ULOBL00ogvTclZQSRwsbRqeKoQo4NEvBXrjNtll2yIxH7
aCMZHdCFLXE8Ny1vezZNbZeJ5DhuYZgPy4gJv1yaM1u/60dCWhajf5StwxUvx9iz
Y5N+Hgc2ULfZ9bwQJeApDhIWi8w9faqCe0x8Gnls40IbeEAfjykaeQv1Aig5VtsC
PE7KGP1FpMi/08O3SwCcrKrec6/54cWmrbpEenHfVWWm6gpF+UR5M3cfUjLALHN9
a13H2VdqZPwDLPcsvE+906AIS9lGXoY6mqvuifWVBxlPovpZ+PuwYzoGoytgCGpO
NHou3y+R6m1aOYhww2sgAsDtNPp4p9e/VYJAiXhN+5x9qJKHAmGoS1lknUL3rvvI
MMs/l3wh0LmS12rz8XTIFaSaTJXdVS0/vaG0cafbmkjfKdh07phKkxL3fJecjoB/
KceEK+mCyt7Ee//1+PMpGkE+pLB4mXTdQQdCPYNiNtbzB5PDNTP/UndLK6ALGW54
jej4BA60F3piv+bcl++Fxn6R0TzpHbZmV8wItoBoXbSmgL0aghODJMR0qxVxpZa0
OjDNTrTIgu07+smIdkDQj3MC3RqkciqUiBn3oT0H4txZI7ORye+is9e4CHSjOyzy
bcamGPGvkyPAlF4ufxqnSk2zQ/HA+6Fk1fKyA93td4gdoH/3e/ibxJvHLPCa2Uam
QDmtNBrycmFfs80SxmzlxQ==
//pragma protect end_data_block
//pragma protect digest_block
rQcSS3V99jLXuaJWgiANGt5L/OE=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_vip_protect

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
BRIMobOjsmlmx4whEkhsEDum7JS0u61JHu6v6w+rP/QsCdTmiswJDjv8aN6OVulU
ht1jHr6PPwzi5dpvo6MXK/R/ZIcrhDNeORmDZYIqY/UQK/IxuVP4eEZ1jpPjygkY
+QPdQUVuJvjH33/64g795/XgVuXt5sphxvWiSkJCRioV1hQTVGFaVA==
//pragma protect end_key_block
//pragma protect digest_block
ecTZLTaHj8uPYKtdePFEED9VYno=
//pragma protect end_digest_block
//pragma protect data_block
ggkjjknQfuyxXqFNWYsDh43e2UQZzAoQE3xeHfVwrdRgIWfOHjGrtkkoex8dX5do
LC2/ximvFudxI9/4eD2214SEp+jlPwyLB7b42naGDcpYsRecQJ2CQImg4aXlzxUQ
2Dw3LIH7xKysJzjrVBhoVFFkuEGbIOI5id09M9VcwLMn7d++PmEIL7nDmMyDp23/
aMkZ5ArLzV7O1qUVRBPqtr8cwUclZLPzUTdCh5QE3ElhMUgBeJLjyDikbKkmhsB+
4Nsi7B/63gQn247wAI3xQpZP4q7TpU+WyxXYTULKGWo2lhdqT3DFHeJKCHaUF2Zv
ZXNgVkFopUCo6CUIQyZY8SrisklVTSHSgynLSwhSqfCbPZ91hQ6JIxR4tqw2u/8W
OOyi15Z7r6WExZbHThi9txEUQrpWBBG1WH+ju97ZBXeA9KcFGa8EESgW0u6RtY6h
Ys8BUagwlDeD+AhZJovD5BGXjJPhUMqLrWWTG/9Vaz+qfcIn8OTap/18fdH5WMP8
Rrdw1LZciFPoa+XY1J3dGnT163Y/kglDxOb6D8tZLq22t05dUYiZyGr7iSTxalY+
40EJUCGEvu2gM5l4Redc5LJhJSw+NLURHfQR36FEH9kzIwl8W+q5NQWquXtgeHAy
EUNq7kJ2JucCyMlzR8KJBvnFQ4ImLGy3Rtz2gyrTzxZJiDP4ber+zb6mSVHzUFD+
9UjAk6eqFXhsHpFzy1qb1CAC7c7q6mE3ks3F3hM+E8nveJelpAohdKd0u8RnAWvw
yfUroBrD8vAJrJecfbRTCJPEJD8WuNqgVaY0V/3xPBrdUJEA1XBwxbeOBtus2eEs
K3Aj/PAHJrjeVjmPIPSmKLSq59wupS1FFu8XPMmGh/dnZ4wRYF6cJ83tKlncbo/b
WFwhgCTZ8wOQYMg/t3B6HN8oG5Ua9YIUxarPzjtsEE/xKbXYRnpkD9gsJqgTTlD/
nEeNQy9k7ScftGhQxM58qQCW+JkooCsG3eTeU3h/9vZ35Q+OsWwqtNYYESr9FmLX
zAv7fJPa2GTHniijk4CPX/hHHUYNJXck/m7aARTveUKtUMVYlWLE2b197vYCHX3c
7OGo2/u58AKl9a0/MPUbF9OmJLPR+yZEqP7ayyVCp9YsBrePEdOEvzTq4/WpXUX+
KRn6Viyv90P0SG8AZeASBbyAgkJg7dyW2TuFbvNGs9iBgYPhvgrYCq+rWs0oFNoE
zfQeiNaBh3fvKF3GignBw8np8zEMhxlDPG2RHwAPizrV8R3va4sgVPt2B+ylBK4z
mEdoiPJ+cC/UDBAtGPIvRgRRu0RL5uehArBIxVNP7agSekk843xoYpDG0Oaed46U
fWwaAvGe/MTRxdE58fJY4v2QK96HFZMej3H80qalq8YGr8adFoHfdWw9femM1CYJ
JUB5zsq1X0ndjEd9GJSaLN3mbfKqQfmDt2PTTngIw/tF+t1UG8BdKgbYEFXGKgVl
AoEmKdIKQ7aTNOLc20PIPkecz1Ay+jRElukycrLRz6ESdsEzlUVG+h4YUqPJnYAb
q99ATzKHYTPSeGuMpivDm2/TtY/SbsN6Ac5b5k0VcIqUP3UQP3NSbz9BC1OOHKUu
1aytSoBdobWmjqJ7KgQhkNNFRKAVan+vZOPlYROaS9i9cyT5dwHX3uF8uiWTSj59
YCCJzi2VSKaTiKekQnjzNmNThGRKfYpb7OOOYTPfiHTrKeH86tfleooKyhkkcx94
yi74THvTyjRCWMcMygWDxZpnhY3QhFIb9R6hRDgPPOXNA8HGvStpYDuA69+XxjlU
o/48ZlQn6xs9JU9WpWMBl0ue/RQFTUcD65La3B5i2WEMbsIJSRt9sIL1qP7plIPp
vDXKhGG7/FkNfCuvCEZ14uiKiho5dDS/VOZ+BlSTccn+54qcUjPQ8izHAE6muXAl
bd6JeX/iJurEUaO6A+PT+PX+5WKCB9ayfn/tr/vCnm1HjhWaOdZxhFa60iIhlUAQ
AtfFm3dvgYGp4dhWVFTR4wFfe/Kz9VLkhnb/7MuvH/7f4MwCBFWUPKii/TwN3p7B
A6bD4KhvSz/MOMwjEOtyGa8kUTFjdGXo3MY6oshBjr6xBCypGiiu8iFliN3Sqc1j
mJfCvMRcknZyFKY8U35PAvNRBYBsEkMTh17Jp/Xt2CqrKV8Mbvp7Fyf8PaRg3iAc
sEsO+U8UUSJcnMSdNd//hoqAMCiaS480RbNBD8PNHugbXiSOp5bMBeJaEjzhHcJ3
d3MI47hujR7ORh4WFWUUgYcOSaUCETUdYkkLvwqJTET/4DftLNEsWxQqt3ngdihI
tPioRAbpVsgNRcsHlAcoxTj3fEc1KwwxVre2gF85UZ9FxdGvZcBJBjGIiM2UVvb5
irUqw/sLd7mgRfUXiNtA2y4M5/cYHuhd2udjmSkgI3zmqPQ1yXIBxdNcjy0QUCce
PnGOUr06qGwoYTONadX428DBhNdLJ2ixDt2DaRdQMqk+CFRhzjvAh1QYkdf5j+jU
fWtH6uZcJenluOBOUaOaYAY1l4YPmOEyPEUhlzL2XKCkWqwDV8nDf0/MKRFsjOX0
P4BKWl7YNgVoCg46Dx1ge4LS5UiMUqnGTCDfR0paIJHOn5OxfKn3Es2/4ebEH1bQ
P82Vi/MZUC6KZZZA4k7a+UWWixyIQ34kIEHV7mNYE0iii+oT5Xqyu0a5sXXAIXvb
hPkSHFqKvmgY7NwbNT33jeJ8Mf9XOsEuM8497WjcpxPmc2GBlk/baxrO+GSxDBGZ
qduKhBZdQvIvqSvGejW5FNYNLJZv1Wc4cqiPf1+rNuS3Cb75ni8EjJMynm77emu+
69eHHEU5mU57UM3GWFB3l7Sh44FBVnUL0jxitt7ofoMuwBEvSL10EeGOQm/gForV
nS9HAslt8XVyZBief0XX7OyWugjB2v91RI5oGxzrv/Dwpih2/PtLN8kN5DnWJwPg
rI9HirgEc7Auc9ER7EimPU9bPJMxBiIxT5zbPKUEG9DMAeIAdewA6AsEGE8BoaGh
y47/5NkasK/k7j/R2JSLI2LgpZfl+Dc5xP0FlnfQHBZxmXx44JVPk3bcGjs53mqk
hJiKYMvsACU1CbVtY1VWSULLHpp53gq3yM3HR8Cu++O5YAIJoexCfJAJ2tYozZxB
A2MyJGZ3qQkRBNNU2Lxct6gQDF9NzhgIw6AldDAsKFr5igHKZD/du4oLM5ABWCgF
V5/tDftEOYrMG6mAc955TZcwh/YkG4DT1KYTQTPNyYVfcOm3fILu+HzBuLxN5srJ
w3RgidUrqymjBUuqvtEycFtIj6/rOKFT2vwCFJE0c17qPW5tN5F+ksWL0UgSoraQ
yxaDDVMezRfeygDxhGT79yNkWdjTD51TTtPd04wjFsV1Qt2JQkWYdWeXqmk8Ezuj
lxz6Wox4Tx5WPLve5agZNLcl6GnixHSKma1S4+lZ5WKOhuNM2YHUfHXz4nNUhsUV
J3aiuTTb7YO5oZyiiLJqO3SmRg58Xnq7jRcx1QKEaCELvsO6ErEekguJMnDj5mDs
y5Pn/a7Bh6qqikFVN5lIxpMOXM13BsASP+1mn/eKNMWgV/1izg3L6gZjCWqbKoxm
3kEcq8BIraq3wEZj5EWha0ftTcPNcdZbqXo/mqx97XyqIZM1pSRNwhfmYzfaO3+p
OXbwDsALr3qZd7VbEGwB+F7UXVI7vseQ1vUhiCu7Ts/6AbtfPJrl+14nc/po3LRp
KaJPzl0gDXS5vK5TFnnGGxAgvJOVgEYnhVeck0b0puv4vpTl/jUd5MZ9WYsrU8b1
KSFbofok7YFEZSS6zBGTUmy7EkpIK2Aq/Fs46sNpA6ENsVNgIFl8PuxTAc/e04R1
TEPUHIyijy2rTRJqb4YcMi+JuL2D+6VZkuTg+cieBpD6p443+PtNS7v33ac209Un
4G0sU7ZAN7N/Vd0rk2ZtpgtLciHGerUzp8tkAxBEkVFqkyJIuRT5IqIDeh60hHNV
rvMNwrBwUTHmHT3fm+OnptCoN9E7QzAcKoWvF1fMsjE4CBkay2v91GRV00Q5dFCn
OXQZxaOWPk2ggL1wACJfqwbpZzjJbU1Ls0zQbQVxl0SYMrEAS5sC4Zxz1BbsjwV8
FobLsIu3o5mE9RTcuqEWOI3zgCkkZjCnp7exlBVLkpCDbE0LZp4nUggWhU6VVT8T
DyZr6eTa/M0qHqr0HCjM/kgFfkorRq8pWbJqPOOH0GM173O6pOv6GnEVm9xgDFd3
fB1rByvhK0AiKnMQ4A5iZO43E4XqvhPtHM1Gz9Ur29NQJS+S/tfMFIhb3XzULFeU
CKTew3ziRPSuIjf3mbxCu4E/gWgEIGpqig9wb0vhpLoHkbaSLDLMquHZfZvQbb/K
gf6nhGoJPR+9+9Hg7Sm000yC7o3XHQ3tL4jsMwgypCBA4OzOScjWOKLgThJPDMR0
C4/jYNTdkii1cPfFtuXXMXVMtNlFOYGCW2nl/4tyoTFFhuNxq8LwB94U0JNLwnrs
4w4fBBIjH95H/SIqbxmoNIVJEbNWeQxOfvM1fZhgD5cxtDGNokQrvSCswGg8r+JS
fkGUNWzjE1jte0VVIlBsliRQUv8a8b4UeB6HEW8xatUGO+1adNsNQR5HfOyBptAW
z1y5STk93PvYt2AGxZ90ULX/n18adon9dTQZ0NqatqxfXh75ZP5XPGUF9OX8Sa/d
EoZDz/9KZRDgrBmB038Q5D7TkveG1UP8ZnibzGZVCYKZbnKpFTRQebsvk6LMt1K0
xB1klXP7ytKpJ+YD7WLSvOsBvlHJmf99BeSbSldNh7rnd+NfwJ4LhjhWgtajTUMP
pVqxhLtvFco89XJbKenxJBkQEWkfoZfzD2spQLjzv4QwlmSkXG0nO1OwXSi5an5K
Q1X1ov1J9jRv5fpqjeow36VrBHFg5Tk15xZvEIUXaY9eBIOc8kUsft7Ic88zc+c+
HRwidcH1r5aUSiv75LJyo13GnVVcRCnze3rIsUHoD1TYP1sx6AU5530OJAb1pBmy
bMM/r62jsr51urSG2sCmbhnXyPoDSJyyJfD54PufICyvB/ztvqjMZqG9+M8LpVcn
xC8XD6JnU9YtF4RXNenexZq79UgGSw0wRpFgJHVRzu+oAQiDaXcVPwdIsqfM0Qnj
HdgTz4o7SpxzfnM2xqL3ve3dfHu9XWlKKlXqdCVVIt1fza9wmRDx9xHHR6F3sPuw
EQzm8HmiDsSLwTa23W0YxokL9k9TkuKu3Six0BwJUKSKEmx+b9ly9nK+IvcXwEHz
EOS4syfO9KEhSqQ44ZIS9BTnKMkM1Hnfv4g3kKIQVSitdmTfEdUlyOKxkfOiUb+9
qQ9ecXYUQqjHeXL0GJLuk8MZNGEca8X4X+Q/GamvzoQvC+7QjlTbXLtNjqOBqUvt
R6AVZtGc+wZkNixMQ2utr0dNxl3rBaQPbVFuR5b7E5Pdm5mr1Oljnjp/m0kmLhBv
6kBqjqVc9Pw0hf5zEfMg63EB1ocoGNlnM8Y0ySHuWAcAiU7kNhjItiGO6/h7RA7U
Lb02AwhAcmb3dqQRw1JH/B80TRjM95BxY+Rz0wWfAg4gT0yYLOZAC49MHH2VpmTL
cbNjJW5BjAf+BYXi7n1UfLxmBCW8yx7wn7jdy8cJfCpwwGJ+yKs766rF7mTW5Dof
aKocq048fSu8LuuzQhgKWgkTvxpr+gZSyxds+oYYl8oqjBac8e26VzoIXkvisXUS
IgLFO/N8JkCcNZybn8v5ITuK353RJTqkmYeEAThNPi3MJCuyCvDtzooS7fwI60FW
reXDc0A9DJR4NrfR+ejcURWbtdvnNACd5RIDj9NDyf4W2hB58lC7VW6E4wEnA7Tg
hvj/3ca97ih+YW6olK7/dsYu+Mr+jFpRSy5W8C/MykJp1D1QG0QVpxZuw0FoKnvl
upvWqDge/+fInLgbjQvjONQVoIlDdMvXCkxXWtB8oY4+IpWdcQUqb2hVtUrV/InW
iL1vQzKfgOGTX2FdyhxhvhAowuMB/5nwA7dmVOjazw8wm+CaXPWrgIuq+5FiTPlo
N7Ro3AWTz2QFochDSOKeTuQm7T2CPfKy0w4rK9A1RZEiwqpRYH5cPFpEhHqHomga
UG+GFklaXxlf4INrW5mTB/o/zHUKymnbN8NYIkmmGiQMjZCjBMoXCeBb5GGnUrtm
DQZkNrSQoZ5bbvfbyUvVTo6skjXi6VdHLAWVZS5/GhH/r0l0LWRW4uTSSsXvSxDs
91gEkowqUI7hhDv0++UA2VZoYcvxSIb5qQA7Jz4PZIewrY0L5DVoFXYVHYI4fZPj
JwHMNGteEFr0QfcgVKWVHFYZ6sSIVNkl9HBjC2sDiqtCa2/BBbFlH41WT8Li0YvQ
ILG47tctRcPrIyCeR0jlr8Lv0RS81w1aqL8QqmgxaBRgScfpUZpWIv/tvaB2rtEp
Zqscv5uhZ82axtzFV8jDVLSiQd6Fgo26INIEIvx5hi3MGvg1tLtvw41YGpRpfOxL
2rAg8yrOuuqaxmfVIjoiLMqltlmluDKXgU9ANMj2dcXAUTl4I4lG5EI+Fxk3tCFr
EPlS1fcWaB+zsSShSCMaslYoTfzyEb86QSwSiIyU6eR1UqciVI8UbYMwlTP2BrA1
EjEqHXUtlCTl8UaUHuZtb6elfl0iOoDu8jQ3K1wptR9J803JHY+Xd6J0eHmrefax
GsLBXarMdNe2dAZro0jeCqy8f2CpBlkUOq6qtixIn/1wrkRAy1McZXhz1VQNwyaC
c74naRUcdN2rrxbA8GRL2XDFVTJHwgu7C5HWhQ/vReiwMQxtrT/wuUo1TkRCqa2y
x81QGlicp7Id0NM596sQ7YetpMezwUgIWcbBef+2Fm8GksdfL3BZCcMyuLx1XWEo
V5949N5S5zrIUnkyi3OrqpgJhxInPuuZPmBb3fX7/5hm3uHxT3dXQYpWBMdHtZNK
V8Nkr5H3LB9g69HCwEUel5C1ZcwQEMltv6vvB3tA+YEZBtmopPZBRzRliLc+jdRw
TmraH/KJfbl5U8UnkliHc3zvmQO3wbNU/qIH3Y5iMWu2L4WBx6UTJmQQjzlkgHcg
zOMAiOmTdj6uYaakgjQ3shbX/ZJ9sullSUFqRHE3zn39YdFLnEuqGHryPFdGCf1l
JPtIxxGZz1xCkyTF8QHC0JRR8npCBsbbVk/mtp0PRpAToZlKvZ6o+EEHPGu4X7Zy
ZeHmgc9m1XNc7bUxNyQq6EuO0oUpRQ1tNLp5wsqn6XXEy1cnAsjMfQmvsGM00ZJq
zJziuaKusmdyByD7Vp0u988Dq4IXvmpUP9NemVEshebuA4/K++nLPQ8a4rO3O3s4
sG54wCBU1lOKbTFe73s+HMCLKdaXARBVeALNOIopJzNEQOJaAthY/lfxTfeX0HLY
XeIFWPnabn9wfh4FIsOdC2mRN/htMNdgU0DI/MT3dERHH8tIE3ihbqxi7r9ws8pA
QaxCJdftz/BXsiwnyt1JIEXO9sPD5V6qrJguMfY4AyFmgQPu12nkLzyGB7nLhwFO
f29T4gqvD7UzYdWPDRNZ0BErepWND3a6vYZQJc9DftVj0LVDImeNyL53FDZiIx30
ARyxnVJgvBIUVIuhk8wI4vD/upGhyPZL4oypBaG3sW7j/togdR/JcD5iApiKYTzS
UEqQeLoxP409QRBu0ctdIaGmO03CSh44Qo9vRNasp1ZjEqJciQmNRW3VIpGOsruv
j/FOX5qNpb4l2dugBs1KpjP8lZTabumqr8GuvQahEnfA6y2Vs7C+spvZSPImE8ig
npdSMfGyetBarcBUkb9FbuoXWDF0expuVJvuJ/tyWg0urjp7daz3Nc2Qyh0E79SF
pCzFPVCsieaSp7BQRt6fY9tlyK+5ZItjCsLNDY+Nr4lniqWDpon2Kie7z97PLRb9
7HDph+uRPLeqlzMqob1pLE6t/CBD/qY2tKI/XTWsHGqPRLXQIAGxg6hvedfVuVFi
QJr54gfh6Eu6tOvhgTTfMlGLjX6uLw3PG/0bf3TfUx2RYrhqVk/uluLZCIIRQQOO
0eBKy8bP8lodjPc/EWFPAziZEXvX3fmaneg4/r+uTzbYx6NAEzekqLDJgUiM7agU
kB4PmJ8R+21P3Uy0lrZujZ1CrIlf6JSo5Uh2ZFeLfzmfrMSrDltZxcYSkn/xXY5l
HNZ8CTfVz2q3cDoOi+5fq6J1jtbC0IZ95J8GoUEiIZflRurN6yMDoZLGMboeu6tp
k944NFUJrQzmk21J9PYl9m0TOEiOuWGsMN10NNs/jj3DFOsdmHMqOM5WpmjPTa7n
xoHrMggmzRdJEG3+k+YTED0x2sXdEj53707ZyNV62scbGnADNP+ICUkipG96e2gi
CpM8LeSRVyKEWqWZrij6LeuQ5+HH4iSttW4TA+g52P8dR0uXaR6sKc+XVByMo/bg
LougHxb50fFg4SXaAReGgZnaYAY6gKJrCoQtycQvGgzEzIF4zBheQMNpNwGDqP4F
WeaJjxcKzWYgRq8l/TBbVqtMT5TlfE6EsEFW/FmBCH8Du0djixsgd9Dkxjtn0jyk
UE1ss94DF7P0tnnj9KuwvwjNQg25p5vFqj4IHycYmzVAB7y7PbBx8cSlP/0QwPMr
1aFiaeCCKnMrffE6cHW9wSPpedrrkFoEla741IS9ou4JJwlPbZnMbSeKBzMFk0vC
QHHI/dA3KqJDFOPrEm43WYyinNwXr6cNVVK0iOP2PtB6xqxk3vKRRw34md1Kf75I
bzAKtJO4Ybb87JOyb0FxS+0Cdy4GgVoyxTjCNWt/exf4e9lk6te2/4qbkHVrL1yp
qzuFjLG1zp5jZieNJ3FlHFTk88YUo4v/H8Lf0ikDdQVW0zYm70zrJIHp4hTcmuic
Z02nS0EyyG1gwY/NdltzapNLXw4Y7fMbyO0/R+5k9RtNwggKvKrpcTIM6ZESwRQZ
u9KkUN2cFgMJsdViQLh0XeB82NbdkgA4wUKubJmRHS1Dgj2ruKTz/WzfaIB2pwY5
U3VzATWSvLPTq5VtbtkqjqPx7ZEfm5wVncbI05VbsQUzGPx0DEsVEIqXnD2SJMjD
KRjYldh88pQS2S+ipqycss7fcFKFVleNb5CTn9cUv8ZGtPHnablYxcriprKVxw7j
+wskGJapIJb/ANgAgY2QXn5MN0baAVnnoaiP5+OTKve0kU7/zYhmSOHan6HAPah6
PnITIpcus+lUzMgrA/8GUPhor7IfhWzPHM2wUNVLpNJd9P16WUZ4H2kTW95SthoH
Ft6ld1+/4H76/O1ZZ5gveP9i+V6McbBPFxYu2MoUPav7zMpjZRCNWweWBV8Uzwkm
CDdWgo0Xtfyk6wLfe4BZNBMlWa9HRDfzPIf1D+GaXSS8+dU+lSH6AAKP7bsXjS6r
PUSsgyA1HXckfVhfYU1FNX8Mj9xVwe0ITAKCHwWFFOQBG4JEJkeTyLDuy6896FsP
MYR/Xt87l/yfCmr7bQCLuugbCyjy0XK1gBXMyEkfoCJ0WslhZWVNJYcVWVnYUEsR
xrt0hNnbh+NlOWI6Tvn7t6orrsU6KW/wlWJ4oOUoseW4oaNY2ThdPsVFH0fxE98C
yZKTTZCxzUGq0/wKhPb2/bmW+vO/9rBpPCaTzZMRY9qMkMesRlWqhlK1YFuvVXNV
DLI41Vp9Q2FCAReQjfEZ4kpLJ8wZ8nVP1Aoz6u+Yi2lNOuP5BLjQGZRIClSx0MJF
nMdxqlWbTxYmgx2vTrhS8Wwa3KnESAZseTPUQHnoU2drTCAw1Hih4Dyt8440MBje
BJ9sruukD3W7uyM6QPLAiLyNyPnj8vs/vchEsWEYnd+c/e3qke6v9sThJ1Yt7Ll0
SwkeIQmOq0lnnIalVIue2djlfXAnyOnocqfIBpByTcCHVYw3ncw2YcqgMLEk9GOw
NTtSqI6oMNepCu0+Y25auVqIK+Wlj0xQAfe7vDnEdIws62zl49Vp8ObP/WVrvwjn
PMy7UJt8wqBZTUZOxrOw0p9GuDtYylPB7xAkCOfF2BrjXvn3G7Xgr6jgQ9zZEHYR
CK2dNIrzdb9kDqKL4BhzZCoGRUczdJRJSHym2D/M66xZRUmRmR0V42RkrQec0O8R
rWo37RpBkSng7zeMTFPIN5oHkbvdRvaEWpk8QE+Ux0hrufSCi93luQAnrmLZe7oY
0q9FeuauJWWlWFdMKgYO+J3GFNYu75Ry5PnTiieyeCMcBhs0dxpDy4mdcC/03MDJ
2BD8RYLcNx0j1W35kaQLfx3e2P2w31iBgIOnfaC3Nfv2QS4cG5qKyxNokKmy2J0J
MufFLk4FgXV9W+QIxZJa3NCIwWVHx3zS4i7/jYFiqdyrExggMHIerbCGt9iGjoWW
/aPm//dxviZ7jJUMNNN6EcbBlWmjMLKay+IaflCnjd8Bd/gnunmE/fZYr2qafAJ1
bnerQLaRjy1uCJkW18w83BxKbAr5f7Jt9nEKu+C0iJnU/KXBmmucYaiUZuuWg9S6
LOcyh4+fNvuGbKmDgInr6GfNgicQf4MbdPADJ06VNKrR5B2+Km95hENWfy3fX1Oc
ozEbfPdac3KC1l7mW53cjMpw4uVwG6E1iP6yPhSRU/GyawBTFoPHMNryFhuhPD4+
sTJwMAw55rP6g5gS8qthE2ZrRZ9mCZHsUGxIfNYjisZhOcPcGn97QZM2P9YYh5wa
rXfvdpqvmQ2qxiGbvA07dOqzZxsUFELxCEgHpYHrRfxlJU+wvfLc5bYMuwpjiMlB
AWjQjyo8PNLg3VZZ8t09+7+srbjcpGtDgtK1C3lZecuuSBH8PZoNP78KVVmLvbO4
OmdvuyRhjd2CCwhPCtkXVcI8S/X7aF4CcVNcNcckPpcgt73yP6bQl8ZNhJ1bjd1k
SKWFczOEjvYRbiCvSxMyZbNUTMAVVp1ntu2zjtPLGhKrWme7rILe2Q5v4E91QvUl
A/vsZ+OENoTncFuN7KU7ClO3RfRocopnzxO7H1szOyZTNIKcaiogQlulxkTyDQqK
DvaHEUJV5r7gmeKfgSd+X/tqr+nMFsLgkyNh4M5LEJ5RWvv6VAS9jvKMaOfH1tyz
foLhVFv3GsHXy2h7cjrTN91eLtqn2JVwm2E8AeTlfIR16njZ5Lmj5PLowHrkTFd0
uXVbRZMMS2Gw8UgoZHE2xNAgJlVn02DeFS5uk5p3VSh+TERuCABKQySWDL61pdsT
1TfPuYjgMufRVOaSDOAFP0Y1kYY05MHgK79YkEBelgsxVuPHb//ovbFezB6BQnxS
c0Z/S3+WZA0sSENaozoHSm+1WE01HiCkHp60vFlkvKsEWfBKC+m7McYHZBqNBo+o
dfoR60Grr2XpXXcuyJeC05QeqRTD3dr31BZg9qwlYJIYnht0s2FUo5dT2nQBo4th
W3TSFWzzqCK4eJeuFmlHdCSTCfDdI48U60vBRERL4avcGKxW2Rsg6k8FJ7E60wHT
xWWaujmvKmelZzbVLvHuyuEEZOQYUD2iGnNzw5YJ5dmzR4VdVKq54pGtx/RnCyvd
gCFSUuCFmdhP3WFPzIiIhSzTWFoCCxXxR59+c9EJuvdnR6uGvT/FYZ5iMVtaUPd3
HJ3vtSLP2zGqQvDdGqItx+0ddBdXojO7OuVgdkQW7FYplfPopMmmKKyGT8Pllc45
EIjG2hM0E9I26NaIAYGM7KhbducsSrjzShFTxR4l1cHa64ltktE2Cfu5MG4oK8EU
EgAXC/kf8DwYT44t5oRhL55HD2cFkwanQTCu5rckG1u61tjo4QEWCvk5gH2yD4az
Ff7BIJl/XsNdfNMmUmUmLfToaTcGsit6zRLTWHJZxlraUeikIVbueGa0Xr+lqwuJ
clWUC7pMmUsrMxZJWJAo93Y5P396QaIkFWpFRHtOPyQIkxQmngx/EhfS5pEPZ5cQ
jRrLYrdcw532HwGGJPXT7GH5P7lxzkCE/CUSbBaHGBq/qLjYKCnMO50l42rBQ5d/
2euvE63wDKWyYeicn9XbqZGoRwFl15EY4CDmB77TmHDTH+RtzPJ39xQRlpIGO4M4
g8+YYAgPSI9cQ718UDjqdu0HsAZQ/PuMtq/0rW62JZLabGUQJrsUwYXxNR+aFLYb
prDaSS+mhyzBABcBJr5GBL+SXCKm0jjo9voQIwZ5XRuwKnjDlDpOyo5wQdi4Y9IL
pR98JUGWmT9kVi1x3myxl7S8ozqQ+riT1CA4REXJHZBEdmWcvbojaBC6Om8LZj3F
191NSqe0xnlnAj0oe1136tqSsDD8tkfwLERrRLRHCmrwy6AjFFjCyDr1tBeYRPHD
8bo8ZmkmLdTtaxng7AkxF+JDqihq06HQrperRZUNvRr0bx0PJ6Sqsdz2yq7nz1mt
+7mk08bLe4WqU7Kn7DvB/x0hNNdNYKNOyC6GuET4281V4dNkVYL7E0hyDYVYoZcl
9/62WNlNpO4Ko7bCppVRYbZrofz5ybWNdk7KT5DizU1gD+QuNDSOW64ZFXldigRF
AIzcUX6hMX3a+y4uel9xphejtHmiEkES29FAGPwxWt3yqS8W/RCmPGtPjlo3/lEs
haCvyylaVk7Sy6dmwv7h4ROrb+uoGRdfA1kPTwZb9AcUYHR6KMLQpvGvpbBaD926
IrQStwz0vXAj7VoKptBiVEtva0198cywe1EFH0MU7FYv9K3HX47DXp0JCbogQaGa
2HNBjjyoN+eZ9W/JzW7oIrKq1ukwHsvZEt4lZKfQ5wgppQIU+Udfw9Fqnv6OrgWi
bDXoLcU/oI0cRYIs5KuLDWXBE5vtrAFTsgAm+Xr3nXms8Bn7r/rPhveoiVs0C0HU
g9MdqixVNjP3kAMSOspotrMYurvRr/WPdix0D+VrMj1Ibges5/JycYQ+80FMu+fB
uUvZqu5DLeUoEsQ1XOh2Y/0nzOhAsdWJ4bWYGyEm4gJsuzXLijP6LmOUOU5nj3ML
8NWw6Gv/A3xk2LQmBX2S98zceklynQvOcf2o3P1JN11e7g63GVCIXGFGfCeTyn1q
K3hpmVyM1h1reEup8xyBwHUZ6UNnc+DrLvjUQXLAshwAn3yjMoh4GnJEpR2SfVcR
LBo6Rp3p2bovsAznpivUXzJBSSlI5IATmyo/9CCeYX+zEizxbYb+837TD0ZBoYKn
DbIeWRlEyXufszIUNCUA/FA6IE3u2t51zZWUx2RdYu1h6BSn+1Ga02qCEo67zIOO
tJrg2McP9FOgC55nuNQGXs1y/BZhPMmjR/6AtqJriS/13zY8lIC8sRgRmiEUhwrf
LTji9dVzvgnFIDE/uD2xVuCmmzEDpm2up+T7PMxCCgBJiyTrLElG3A9o7M1RvWVu
sQ2ce79iwxziZS0uEyou3ZPdWnjNG44GsZ3nn/wnJHM7d4t3WbRjHZRPCVfvlTc+
Umdd0iFJiBeg0xBZp3/rUzv555Bq1Vdya60bMWISy2+hcApANl21RuXfagULE9Mm
Gh8rSCOkZ7+5v2PdWS51Ltm7w38HHNmQ+KyV82vQ+13qyqOt+y7SSEgz8PByfe3D
9oVnpy+00OP8TisWYnQ+xDwnUsb7gDRsrbWWgJsTjMXDZicpL7TPG5KLwxxD2SBS
m46EoEfCixjg+CQhxh47tsuISVdm9wugbBg5bMLqiqLJ6vQZXti6KGPZktn9Kwxs
u9kttV6EHtClqT2Vh1lWHSbEe1mPJmdPSWc1Ytpw0k+yPZFD10os1Sz0TcxrG2X6
coyYrj0oLIdEG5y1pkKTbsfrR7H7teUZJ+mIhzv4rVhAgiIbGss8l/sh/GLKdnLj
LB6iwXWNlznENMGFoK2RlwmRKOuiWBCIbm5gHBZm7EPjJuWRYDmDJtck+xvxTCgm
xKYlHeiOoWlwUF5ErXKG7vBtpoKK7lcGCd6I4qiCl+RzXqQBJHSultA2hOvXoBlK
rXc8m0eqzOtKjz9DUfru88Sb6xSnyMfAAn3bZlIrFqL1zAvqpw6dD7YXo77FRe3V
e1WcBWwCjJKgrmzuHiUj6o+XcTUj6VsXulI3oziud5XozEKm5X86WSoH13kEWMDW
TPt6HqssiEtRxoP1veMASHXHfSKe4z5pYGXkcRx357rf5uk7AacRQk9VnXGfFSNq
MQs5CaCGNtmFUlf5xxPbLgmfMYu8kft9v4AWgoe7NFdk7AegPUeZeqzAEc74gZU/
s00OcHcqWNzOmVEPd5t4SEYi8DkpZi+sJJZRQpOzDGWPrhm8zUNcNrKsVTsE6rcW
VmcBpSbhYXzjLGQPRqhupcrpIHgXWqFNDqm+bPgGWVSuPv2p4JqISCRzhjMnZiWb
kj1plEcr1LLIilZcefcTeeRZeEhllU6S5FIbYiRZ40NkyJ2KwaHCT5YLix4ZpkIz
RC3D5fl1jEmR4KSU/Z9ctjjHCzwyi+1n1Eiapk2vPw9cIiEnEDOIoR71qA0Kr/n8
06LCXmjpkkqCBMPcHbkcf5IwNN8QPwe/NwHVa6uFOAb2I5Z3hjNRXnU1nZ8pJvjb
MQckUJp1pujS5qXbhmQAPnnLmnPHbpuVs86fN2GEqWTLPsSh1tzN/WHzMEjjoNRb
yY3DIsj48AYiZs55bFqbPKZTlrgtW3INVbMvlqSqCGnXP7ea/H0Cwzn3a9MebmiR
wqAocTHOGMFMZQEpF0bRwhY80iEMDVbzPIR8FuJ6tq4A+k9ggyT/yiCgaUflL+EU
aEDNbSznaNypkw3CTmoGP9hSFSeiycfOyhuhJTEjfnCSb1/f11+3jV15FwDUBDNg
TVAf1Nb3Cg8ULhO+ww1as5tmSHK7Fz1pwCk0R00RLgX+r2F2zclzQuUFHarDmIkN
BmjVjBELzY1Qvp6csTn/1LWS4YKSEA8vKu/YCyfCpaZrSJ9NwLTyMDnuqS9gl45C
lUATM0F2WIeehrlh8Z3y8Pqt8jewKgk7C7CujrGAxq67nzpl257+PzvnxskvC8nE
b9TSTlQe2GaGhBwnYxerht6Y2g5NfRZlkFaia3J9ld+69YLaD3ceKmBKFARpg1nd
Y2AjeKpPh5X/e0fY6pJ9XlRVD99Sq3ykfakZliKPnY1NTuFPsgJO3nlnjhWIy0zM
ARTfOPp8TbrYVFn0E9AqgQrHrIAywQTJetbaUbg+Kh0WfpDi2kpMp8IN5ItUHnjN
CPsl5hhxT72WLmLUdvVdabTc2ZutOHQZpp9D+dgWUCkUhpV243CLL6WIEZK0CGq9
DzQhQUCj7+3HwiubLmIrPtZ5MFggn1EutoH67Wc3OQAa6Fgonm9u5Wn0/y1Q2Yw4
TG+o3sU4kI9Icl4rkEetghEHyOBcdsrvVQjCE0gdooeMV+qcBjyKKO+b7tCC4GBs
KFZA42PaXLeZivwN+VCCPSatgGEO3hdQYMETEIZ6OSpX68tHdr7v2xL1Dn7OWEqS
RJ7bbUg0gXb2kFk7R0Z8XGkzHcyoQ4rx1EsnJiYcjBcTTgo8Vz1u/MjRL+0qbCtf
YN1ozETJMv/eIAGw1GIjJgxlKSSrAEppcgXIaf7RbbwaJEp6JIItH7XDfB4jRIhh
SwBOb9ddDZdiquekWXogQhkWgnwSpf8Oi3aQ8fLGo1YXRkFbbJX4U/yCreDqEO5T
j0RbpGFK097lKCTL4lb/uSICkJQom1zsS90bJyJqE6LhRho4qEEvZbnQhKszYDgr
/eErUEJHEHV1tbZbsvbAO59g1Qicv5FgFcbl3Vl1RZzyf0GTp+5PWm/4dtpSVeuB
LE5FEgCtuQ1dJDVTYQyM6Iog1Cx+y9LJX26ywLi7Y2vDiZZJZpHmkfkumvwQ5tRl
7FfQSrJAk3kugYIMYO0oUu+5i/1W8VRRvcoGSsu18ik3f+xGDp686liKo6GSXchj
rzIk5fJ9cYdzDLUt5PXYaDxD3smgW0gvWwKjmtLKT/hXBcfvT6G0Udrfy4lryaeX
GJBYxVVydVZ12Dl0A/CUWMAwcEZB3A2Rt8iO4Yu1zsy7VYL1g3zRfoNpR8gtn3Xm
kZBkLb7+zCUQj6WFL91hXUeyPW1wIATvhFXKogv/ggyhun+Xww8Fvn/HDZr0bW7I
3yPspl/VljlBk54YbXRHvrynJMO0yAuh/o4BkhRcQjTGj+obtYX+bWu3IQHVXnRG
KEL2v+p1XcH/nHoaF84v31gD0l/y5kb55dEiGv7yrcG42VoRkGgwej+WgYwck5cz
DeAIAgtoyZlHZmjN31nzyHXta0miOj/bkm3tMWCg787//WcVzBUu7vAE/fkgLzGa
QFmcQx3TBRx9aRPMPf+OBH+cS1NHnFpdAE49Lc1udcj0CGiToY5m6SI8H5MIKVzW
cTpsZbdrFMyBFqnkTjE583tMZs6L0/emrFgHhme7nrXTdwhJM8J5mt/O1fLjufUW
FxXdfSzK+bb1x0T1I9Y4AD5OZglBFCPOaGoCdfTKB2TURcebRCRGBK9TdtCUh9+b
ewJIZl7JAB900jvkkrhiIN7CnbIdrmAL3AMS0jpXcZk1cd+FgGn1vopwMwVhTiYM
jEIzLOg2F4QN4zCRGWi7JfbSpJNnVS5NA3X63HhATAtfTfg/DwSTt623uQxU4o/y
qqazHiU0QqjC0WHb0HGERbtU5cm+tL+8WDa5dvgn/0Ne6e31ZZtyVBRT3nUfZzlJ
mLaQ0w7lVS3rg/bRBwyNWdFCRL3iHcM9s7NEXUsLkDrtOGbI163woUgLhao5CMPd
1HdPt7tzPQnEmtbbITr3BkZeDeizsHfvULouvoM0uLqHqc+EmhXQcQU3lJVCjcRu
g1r+jTC7INy2Ei7i7dUhQJ6U/ae/0DVpAqB6GJDNxgLDgvXEsqN8JN3X2eYQtIvU
JHzwRwF4utSNEI7uzySX0mg4pOM9O22gEcBClPQg6JT9cfzAcYrKorwPaaZegBBt
+RMpHX1D02E8TjKvl16WoG8QH0hDfQxbAX0fJcdEUl2qXOtaRgFG8GS/HAUAQc7A
7CcopiLm+QrqLq76jJXgsOdmHMGvm+QBAq0iDSDLzOY/cqXGxH7QBsT/sw432MSs
5sB4wXRvVA+/hvyWaxK25ecEvL6yud9sT0bF+fLzOCJdV/gRZ7+lJpxoQZY2MgiD
8m2wM2G3sV0XODlRFry8jkh3lC/+Hs8cywbGjSTCtC2ZHW7xbYsFscqBshFSzwxD
M+y+GjYQJ4/UOgXLUCIAynkKiewq1Y2zP3h6GLfE0J7ivOWUc7eCXc8VgAM5Rmvb
/VyStONLhUYZUmvl+OPdRakTaMYNeovS7903P0uK9nVvGruuAZd5QYURrLn9KzkU
A5dhYfA0jh6+sHIUarGkEzgywdkOVkxu5qNe6C5D0CpnPkayhjHG5QaQQ0vmW8aD
UL0YRg1bViqpoxuAqNZ6jh6bUwfN/NLEtTkI2uVFjhm9ZHy5+hS+EDzU8jLu0vo3
wsQ8I1EA47wib92HC8s5G/mwe/4bZQdKMmZu22/d2zSpWLP4ZgiYasSUOZGMGXSl
i7skMxMuPf8vM6NaZCWCkORuds3GkvMeGboSRNEnh77pVMvBq+jg3c0kqidif0O6
ekeuMcePn7GEus/cMKO18fXl2Y9Lxk+dBHt5xEQGc8e/V1YbDOYq+iuxBHzQp2kH
/+RpS169CtjqiZjPfMaJ/XAQcUoOTJ16wW9PjV/Dp+chS0gGq/We9pIr0YLlOjhD
q/4a4KzRPFcQqyMA6+Tg6mTKG2y36TIAY15sUAfvrQPvcyrmqq7SZn3W0xlT7pwP
gRoiLC3Wmh8gzQUXvKiMw2dKiAqxlOli6caGaBHffrtySj0yOcqinPLo22nbmUdO
pFNDsuvC7C5qSuwL7fXAoFpOt6MYjEX+xlCHPSTQnXGJCYQLMcCq3h1LmyeOEaR0
+MgpgdDFaNSVJ46gQXmzrbt/JXZrgKiIEjPvLaIg7GUzyZQenf4Uyyeuvh4qMCOT
OL9vSgg0lIOvXDeJLj+E7urqbScZKzVfV5I2LF/PpbciB+Tx5anwPggaCekesyEb
IeG0JsZm2KKvJ5UYhWEf2TwS5lyxBivQ1dpAYpcsVC22bMt4M21weG+wOaiP1vVW
9YBRy867gkfpn0waSlu7/7m9B4gRWM/M4cbMzJgCXfOB59vyfPAZ1GX1KxJcKfM3
nPzpvp8+LlypWUF9pRBRQU7YqPZuvVg9KM3Est72CJ2t8n8GdVQwrikVvS4Oid+C
H2XHAVeJ80FZ7NnMPTINPeOqj7dK+/jL7TnMA9Qlumd3jzvGsXUe7PQB3G61obYV
GLqulRrELkPHkEueT8BHq/nac3+YG9GbUFevCBkHAwbQbpE2OL9PoxyBHEVvhIVm
Jz2WlH9p7TVMTinsJGA1wmXsq4Ly7k1iI03T4VmOLq4R5MvktYB0mQ2onA25nrBi
gMuLcUR5vIPPpHJVXqNNVl6q4DyIZ27jPmFiP/uFEmjF0ER0I/4YArGuEK0KRFKi
3pB8PaC4CXAy0XxALiwhKJyLbkRTJihFDdz/o+0xS3N5DnoraXqUJjSQkSiR3BYp
KZ7JkdQMlLyrTgNmoplLB8XN742Hji60gQxwOZgxCzekjmPY5iGylSINLNkbN6ad
7NsOxsy2343s43M4wL7Cao6RmGV2bvxdzETd6Q2NjQ0A4276HwCpOgTgiamBC3xv
nTGKRhZXAHe5tqQJWtts98+Jy8zKTCeNzkmDcNp9lx3rq2/ti1GrLm1N5vg6aKwY
VwK82dbPi6grRzBFEPBN1LLyncTN+XkcBj+dFsIlD5Z77ZALRTjVVszlA+5dRpqe
IrtRAfxARVVKIM2BsuCOgOws8x0BRXS8o7AINqJm5te4WofreMpJMk6Rb8UzuyrY
Lz2LDEvWb8F66QnWNHmucxsNeKfvKyEdWh8iTz5xnOwCbvQKKLYDsWO65uRhZLfe
VWsMlrIGPsiD3znjv6ww+mj8bFII7c3eY7a8XKPE5Gz8Hs+DvAqGDkBSVPeEfER8
fd5HtKryfMGxaEX6PqSgInBAFCYxVsg9cy+VLAJ7rrao5eVSWAnXoZPZ6gD8MOoX
ZTsHPnwqs+FodCZyI33m6iAdxR3aqb5Mg++uAcXC/RJVM6KP+GzbmOAmQxJLMCJA
2fMKJJzsiHr59q2Zf4QW4NTd8PIABCSRY1eWeg8L5eIsuxQzzYptTNOCFMYE08ZH
iffW2NagMwinShqD0ZjjqDgze41Z8tpGc5vCi2ZhDEG/m0iiEZtZQ85V0HXMD7il
K6DU6bAlQecb2XenQIpU5e5gZt1cdrR+hSbF8L2wMtxgtL4Ax7XshAcAkF8n0xRt
UtoEOzkns7a+jXu8JoNqdCIH8BSMnAi+ae8zzTyCDBjNv6ZTtSuMfLqH3kvdVUEe
0ViaRZ7LJEoeEiVyefWLGtiMXKgZE9wepRZXstjawhuN//AkA0zPZOkvdWtcLiss
5LPCtQRyEtL2Z7gBXKT4hLT9KZ7c5wAZXkOJA02jwSEhJ512jSMBrMEcEjvk+svc
fOaqGc2jpi5LP6dOotH/j6KDUM0T6tczAOUV6WAd1Z9Tabn7Dj6ZYgDC0E9g0TRG
I+oBGfA7JQUcW1Bbk4wDw/BKDufJNbZImYqthYJVH9FBrpJjfkPlOGGGoBgUnKXD
ZSYx+WhlbarzY4J8hXZpKzYWjwuVfDhvqR1PnkcB62tQcQ5lxBjgir+lHueAGDCU
O9B6muInzHTmZOqJTC7hyEIhSnQ8+vaNM6VjHab/Pw9frkzVWL1coHFV1XRnVJdg
2TkwPNlahAws5FgXLSElg7tix1zZyaieHalNLa4SBO+ggswZBGH4Hz/I3xMy1KZU
VZMOfwvRacyAOi2WbR3nFweSf5p2eDqjVPR6+GRNIUnkRpYz5jKLiUcLb+9cxO3z
JCP774AuDxMMCfiukOe6DEYMhYxcUWy1KbL4cstWqnHHD+hTDLWV9vYpBThCJ+yl
LpTbk+1v5uOmzpnKPsVrUekCSXZ6aU+4Whe4OAbLfWTBQqUcPLPIM+HQhNgytaVu
w4FMnYp2cJIzX3KsBXm4S10dvD6Nd7g7ZAkuAZiSoS9q/fGwnDubWgYMgliHTf04
6miRsdn6UE5ke6XT3EnTKf04u1cr8aG0q+M+QpUbnesbz19z+kun5qtZDxfAX+M1
fc93JR9F5o5Bw1OIvw7eWJUCN8IsQwKj5LsZTE9R0IXQX0BiVhI1vVyWAImYw11V
dHHldFL95gfRwpRLuWV5ynIoQ6h4vgSzVK54QljYeH+Wk30TgV7ZeSVmemTV//Nm
Vi4Z2pMzmeIr+O52s9Nxs/RK4YJzeOPhEM8UD5QErZWxvyNeMk7U7MLZv/iSfj8s
HfDRwCFMSqd3QjvFxNHTisJH1YQ1eyRXPxjZyuCHrk+0qDm6sO0YpdKRFjTpKedR
W9iz5gHgW41lqDWQhL6FgQXYTp7bwEWbfUi2GuDhYaJ671Sch0K3LCrAuorHo4CI
vfq2eYxjZZHzVK+poRah3iCIroylZB9BOLa3fd8bWATUsPAiVFV4mGisZ5xo1dHE
e4cdqJpCoJN83v8PUPDN4WefYzB3HGulQNT/HFV9d9iHF97wWedoa/5gVBnYi+sr
diHxo3YbvhkqKUHwYBqBNiWtUG66BaSQvTvZggP+eQ+urp0jXRjATeUm8aE/bubh
o7R8Wz+3PRR/8+A8rhvbcahi/vFt1cmyGXeI9EwOp25ai9IK+v+aSZzFWk6wbNSK
DqgG9tS6+NQ9nShcqklMyh3YWikDLxWyqrRBoIrqr+NlgvUsCIYLXqg5B7Tplrwg
rjHCUKcKUf8UdB7kwazDflCJxzW0tzih3qNTDFpGT23/nFgePZw2I+MEnDqlc0P3
toHbD0ElDoOCBKPa/fuiXLfIcpzrzgkuT3gTu6r2Sqx9kvvAvIw2lMFtL08LcNX6
VmPic8nRJEv0HtGsJtZ3ljbbOwjo27L6AFKekrfkjx5aV5kmrgNXKRjMQwVmp4Rp
BhD43r+MG2BgV3+HVNcJ0Km+9y8xOzVZXIzn5LS/iuWNtY6jl/AdF0jjy0St2uQQ
00qAVkqwRI8+7IgP5MHEMMAgEisY+jDok/rkaUJiyDibpg1MrA4ffxHX/7QESG+z
CwifpAXsOA7WOohhLuRGQzoWgZ8sg2QmvApmTydUeLIWXHQkvRhZlrB4MsFCTeqw
3TNtem3qhQLqPPA6zS6JFuNkoKp69gswilWB+/AcAUnYtTxxvZG6SDpeNqd4pJ6n
Gs3lD0RGdzrL6IDJKtWi8zArfTc3Ve4Ip2vEW6umOij28iF6AyLHAprnPKkVP/aI
tZkOy/7NT0gHEYFl4fEy6kJulPo+hO2zMp/aj0q0bkm6++UT+TohI0k3aNo+otoj
nNO4EaTULZnmYwQ2tEM4qi4Ys3CdqP7eq9b05OxC+xd+lxro/zgNfpJDU8PjccsA
teTJpjjbKkjggHE1IhEkpKdIo/HofuOECvQBM4y9nRV1aBtEv12IZnkDALlcqmAh
/vbpxxPcGx2O0m8UB/8OchOb5zr36c1cp1PqZbWAeKsoHsWfu1ZZ/PGZN6ZniYss
zr+Yfz0ooEqewqC5c0iE7B9FACzxlaINUTZ5zgAqvNBpID9S3t29MtpgIpwoWafh
p5xadMT892Hu3xpk6LY14wHCncsVAQVqLMZqRs+lNv4a9NwZNIv/8AxKryP2KwDS
pCAFvgFSFJze4Clb5wm6gAxgeF08/LfYfPVHfwJ4e/b7moxLUueeaAzzNWwSuj/4
XOM/8dLS3b4H0hwsDBEsMiIUdyhrpS6MIFvA0dDI5QGaaLKMz5RbMItE9eeVQkbR
Cx9qkoxsoot/IIzspOxqoYODgbkcKG2VRJkBMsPGK9uxlInCRXTC4uOlMy1OAwFt
Ogk/HFvO5HcC87CjDAXf1cFhelrB8O0S9tTqtghkarbrObu3njXhR6AfDgx312vY
aa9T3gQ1AGR1I4xvXuJsaIB5HBRmlg9GNNQvjI9mtzSSOSSUm/6ZviH0az33ttNr
fJNMpUIECYzj9oW9R9Q/A+Hfm5siQOBQzLDKY74Mcb7XpEqlfjXWV79maIwCFlP8
Iqpxyj7up9VwWyR5YHBJW82ysSjqYJy8W3X7S6tr2YI5V6LH3fsH4V5/GmE3avY1
PjVhPVoIbvUq2YsALBc6xONRlDjfc7AGvp00qfFHDYVEUJBiLhKOu8dw3/abxj9e
4z6x9OHLXU8FGNQx4Sn4RzCOxPRkRFdDyrXgcIW90drhYRzNEnI4KctmGGffRRfn
LqV3fTLTIGbT4eHMcd3dT+2qqaOezySg6fAZ1d8G7AOr92EZGaAz7ekpCgWb/8ii
SZYGrdq/raZ5Nw0IPCjmVGrRWgy5TLUBWfQOoDncgR+z2JGcu9Mc1WU0cSch68++
MA7Ay36eYPFhF6quTeOcBxjXFe6kuyLADaK9HQiZrj47WDhO+w2dl3fpp0b9G7i6
u2VundTpIrrBrRrZ1dImhcBQllLHDHl+w07PZjJgdmO3ylS+0J9NHZvdNTHcz1CI
INcnO2YU6f6aOIhBV1STewoMqjn/F95CGAL0CB2uveAxwFM1TSvFpXqBtGHnSuiA
qVnhDP+2d0vTsEQ8mehA5mr7VNUibJqGc/3Nnupa1gC7UkMghBq1tji+9Zf8nGtZ
FtsmmDGvZxpKH2xmWXB97xO4cgutQEiv8RgYfkuTi5wB/G1xgqPoJHfVQwCURbDK
fBORjREM4A/j+ZpOBqi6M1U2byersAXBRu9Jkn1v/bXNPLh8L5KtPRiWvShmOarg
LowmTrEcUJQFZtSC+gvTOWTE/yfBBNEM4jmV6absax/v4THyZToZqxjMkW900uG5
VxqbLeScAV20KincNT2/uHJc1CQ1W02XbXYvLwx8g54AeXYJg9wLMM4CbnFPy8LN
R3+DyBZCDtUHeke4d1z9mWV8nrjqM1PM34Mk+Nv62cJEXrYxpdYtu9lvn6iAV6eu
8k0771TpaZVyIRvwbblK0or0o+g8cR01oMPtN0LtwCu2z15lpyR3PMBxWJKFryA4
LQVOtqkqgPIPo334dVON2Y2LWDK+hNu5seisydThUTAGvi6bIQMl1TwwocnmRy6D
69JwDrWpADQ401iuVoZPZ0cB9/FqHRCG9Zyh5ZPOB3SehBE++OS7bMZuho5kTe3I
zLG8iBu1zO2klcSCrr5iOHIhSKBHh/0AV2ZzgHz0szHOVC+onzMScu2GkjfRGDm5
UPFjnssu16ILMh3UP8jJSfo8K17OfYza07mxF9vjNQLbhwf8vhYIpAfvOwTNSts4
WWzhh09zW4GHJ1DPdEWNO3/6+W/+ymMA11LSCR33Qb7e5BF4OnVRZrMkb6rV5c81
jsMhfDFEODu3s1O1l3+VxqvnjVUSUWi/90b696crvzUj53RIQ8686DOIf3NseIPk
YsgL1pURBbDGFoxGDskJ0MS1AIWjXrAD4NOixX2GYEmpa3estiYTXJ04SvTh1p3s
BPtJ3r7wqi5zfBhkvrvQknMU+kLs+mc6T/U72KUvRlTgBLXaKuKMgsaoX3R2IalH
27u7eaFG7beN3eqa9jcuIIhasMDG8w8MsDHGINheenZPghKumhIC8jNLjDJmOFJz
lMW+3pMJ+Wxn0pDAvwEIhtfEXT7nR3w0jcbxRm2qgm0KM7PEf3DCLX9WFvNlDBCm
1eZVi5WdrDGSi26ExF+ROvsjqVuhhQ7GhjIaPUlSEEM3FkWCtQKy8GsUfGr+1tyv
i6+x9JdB/av4lebkKiASf07IMY4SmeZNUWEbGyfCA5QPwG87BImFDPgcC88DVbNY
dLz3FebMu1J5xIoJcUCyLPYXdY/E8Wg2uJ+Ci9ED25pWaMMW2iV6eMF5+UQXom1S
fzXaNwlYDscBdGy3hobbdLh2GU2Kn6jYyU7CoAA10YiGx98/swkmiGNR8TOx8YYV
cuH1Gd/ImIGtE8/EQSnESe8jtLQHtbj1XJ6pSTGMAL9XOY7fSV5DcO8sQZ/lseDG
HUftfVkpP0p0+qSZ1xG8JbVr7kk/bNjUjZpm0vuCxjJc/jgKoqSopou152uNZP4G
sV5W9Jo2MOqP70REjuAivsm0jTfwMFoayB++yE/9whg3cJmNnEHgPD5TforbZeNj
915AuPWIuQp16oRNYAFi1kI/o1giwhK21KUvfc9+RIcu1MAQoS+QxBLPyLUCkC5G
rZ/6U4lxe7kbEWvRxM7j9f5gDXXdEDw9ihuXQmXDCz9H3wZT7eOqg/PLNeKmNj9t
IvqYLMAYULYp21MKWtIq/gc/tuSGZ4+pMmjffHalChGU6pIrY+dW9OQau18/WpNI
LHgaXB+h7dLeTBfJWHuPiE1XoOsrYKVMs7hjVEhDXCTklONhBHpIxAu6+bdIAVCy
V2VqyLV/Tm3PN3eV3Rmwqqu4x9+Ui/tEYTEYhQNtVfMXOJOv/YBdGjWjvRG3IqhN
L2296OhoGg53PevSRcc3mKN+kkUxyYd3n6hfV0Q4jKw56NcDADtMHMKTwaC48rr2
qPdR1NgGoyyd6HLwuXjTbUCnyBvXoFsvAW8nRDIwzHR2w7lAAvi1SKaSWFZVT6pm
0gSEgN4Aeau/uOIU09TdYtn1R6L+GSjKHHbKfvEtmKVa38Dz2glk2m4O0eldJvLt
x0Az7SBd1EEECDNBGqKd5zu+d1oQ/dTD/c4cPpQaf1uxoCV2EgB1z9PooKyQmVDL
uzNPCMIGatigEhNHA1X7od7z+vy5U1fzx25qzAiSHd9QLGzeIAcfSNLDodU0MdFA
zJyTm0/tzzOtaqnBM2NuSJ4QZEFK+bWwQS/VPWunhDuQiN9VmruVqjoucP46t4Cx
ktMxctczwWgORJcfOGXtBSU4kN4Yu0qcnBZkY/uHL6Sgg0295nu9ge3MDOQPX5G0
GCtL4bWTB+PWANK15yQcCUW1EJRvjeWwJG88WkGyBPOb3clUmeJl3AEH00SK1uv/
XR85QboH7rlFbaJzpTQCOxCXpwO8X1hx/030QicpymWvBMaBhCzI5JDLeBh50vvl
/57WFxx2IewVPYIYGaepyUAOwfppgpgZ6VErFhmD3esFlzLdy/ziBkJtb+O7gxNH
bgnLhOXgFSqCcbfO37c+bu5E2tN2UW6451fGNS8u5QGiBGlkcgJrGtRFJMiAFBc8
gPWJb3i9ju2WOx/p5IH0pNxYEytXdCiV4T6pxXHsrlqJSGx6nn9uh1n8MWsCfKY0
yzbUILN1YUJW95+xNuoeDg5Etqv25rbW44VxpgyzUXXzWshi4d3O0EAkH7+Kddgj
BJVH6guM0E8LWQtHtOCPNfytDOq1CFdRS+pwxOxWkwzVrQwI7xqis0YMqYQwg+6q
1Kdd6WU+1+KCrOlZAV7eXi5OBzNaxPMlOV3qgRTFfu82LcUByIuGplnzGIFIyDNI
llr1H2l4VTafktAGRf5m748uQ3A0A9RXMe/xAEyGRba2T2Lv+rHu9fvFrV+MRUPd
DeqmFbtk1bnD/xytE3v8vRTrUpbkHdhNdvdzaBJFQVgIP3SLQbO9Jn+6Ti8Nf+7N
OFcVUsA+kJAaL5iSIpBfV7TMTcFV4sktbHAx084+weKE7/zeFYJo9fMDIactbrfv
gRA7T/fJXzlL7sm3lVhj0po8C4qEH3WKsH9I2GIg4bI8Sxj0m5Pvj7tqs5nu4C+i
F08ftvk1tiK2HGGsEcaUdaOd/hIVAFNkKtW59M8P07IDrlSu/CwymphPPwV1/taV
ARTp1T1OGTzOsmCtMRcFxPKrDadMszOUKcgpqU+xBmb9/ExwLIlMp2iSrYM1YHLH
UAqzotHpaggRtfdmQOmXz0E4+4FKrcm7lrhyjReNynWWqAAIntV0uh1CXJrAeSt8
+/devmAETKLoCQI5vjykNqdONoX9UTXiHHwE7r6BczIwLVFXsy9hNyohiE07CYOw
jaMFqg3+PkVv1oiAYIcrqw9RGJqQYB2053f75cseSVWkzqer5x9sayJmH5aKPpGO
EHz7nct1szMxk5oZGc00Qp4D3brZGf0147kkM4+8aZfEjzlR505qKLp6ghWxbRIu
qtffzrLb7qs3LJ3LApK6txDJaUtdbXtDMHowY4+Am+s1RQO/UqgZTgSCDweMz9fa
1pBPOz+Kg9oWz3PYiyCIgRgJ53QiXpX5gw4uHQZ8m9pDpGD3JiivQ2GlmVjIE2Bg
qayOhVszdzrgfUyckr2ev7RnUlgBG+3ldOcyT3VWxRWkAbUmkzdWf9EHr4T6+l7i
tjbj6hHOfD88onc8SORdQCPRPrQIlz4T2gYBCOBJzCEW7uHB1UvQfaaAjyRC5kmA
f6GBGhIBbLyCVQlCiE0GK3OrR3NuTrpdTp9WjDtiv3Yf9kVBm3XYU1Pmwpjig/J/
iZMSrT+BMoAGbJFRMeUbHTKhuVMsl5eZUIvCnxoDBXX1rLFvYoL7q+QRyd2MJpjH
/76LBhes4fDkAT9JnbZOYyzeznGD6Pc/pCzyGHYqD/h0zoljDaJcwEQbjnsyjeth
K+CyAf3DP7TTPnQQRMQY7b2Lb1oogHBRgyK55wOu2qMnc/XA3VSzRsqQPbs3w12v
iiT7feJXoZ288K5L+lPL6Gf/QwwQSdsUN7LpyioU8LPAol5YjiFjDMfa5zGo564P
3KqBglQVmtTWCUd4ZjMUngn9b6K6VGrPB1rc6kWv1QU9MhkcIcgyjJgArHg5nh0W
BkUjYH5bRUmTuhmJS2AFWFH09sspyfC6R05IESuqpuBKeec3VCJBX62p2xfKUHi4
IDL+5Sjd9qYoHIV53qleEgr2qpdkgHG6uG2tc0h02hec5V9BGBN58flMPUk1J59D
QnOg3kVGGLGfoaqlVenbvCPyzlsO9hv/l3JxIfDQPLUtltKi7OUOYRyRzoegrRBI
zUgQR6pAn7HZzZ9DYG2ZMEHV7n0qKoc+c71ITrVsIhV2HTc9kS1HDBKtdTuhdfDX
t5HWfHPLy6EziknNAVVoNd+HGmmXP2++6uQpoD4A67px3A1RNJIezmDqSI6JZx8/
IxEYflwFhgRktOax1GsQvI2jrqcAuSPpaxpHUl7HPj6PIanR/DDkuO6qxnTrvFwI
GPgoBqg4p+xTquvNkmmCmQyd+Yr0gJ0AkslqSx+WiP4AhEYHNa5GjQUzgmR2tENz
Z26uYmzohxuYHQg9S52tojbP3C1M6D1FA0Q+pGW5XstO9/Q6W+Vh63I/XEKFmUqG
iMbTiK+m2z3hRR/c/QQmOELuagV6CVatAUK95qmC0gKMlSXqMUpvczODr7uW7L/S
aFSvQHthQ7XbaeRZSmF+ez6vVJ17VMlhNwkvdFi1xbMNOwXkX6t/thYsIuufCQvb
d/vJvE8EBUmsfHPlfgKSVILpw0RDlN6tjV94LOiMY7XmKj5GgINdeWP4D+R7+9iX
8wHDuGDBJisKgFM4H8rzId6BLtRLogmsyk8dYTAfhhENNCG5aTnnnCZiD81d/r4w
0CrEcSjIElSK1j7UdK5l5PTtxVFRHd+G3BMaukGefV76ULtt/6+1KKy26TbKOQgA
V9N8pXBEf8TOtRfGO8UfHvQOIp3I0g/G08vY6tExo3LxYdrUGRxqDKfQTcY9ziVK
NA6rGZtxMDvh6q2B6EIob0a0BbOBBnVtyTxEq05BR68oiVI2b/tMt+OXUyaTgn2B
Km4xZrhz9wipy6YXHw3s3BBKYLxzpgCrmSWnkp/TrdvItj/dvptcoyh1tu7dsTyO
Q6uUxTq4Z8mU4zbG95SnEtoz+k8LwyOvqQpxAmH0TbAK/PrOwJXlvp+jNhQraHcy
tdDoRl0P8I06Ma8E0bw19oVAjM57L94nVgvwiLN5Yr6l06me1IPmgvA6dHj/uNR1
khm75a7rAjs96L9hzYnbkEbnoxHYHGs4PLbxoQlXj43u3H9w/k66zXvjZy3DlIOl
EAQumUTizY2LtjXJP7AoHP6C/nfgR7IcsJ/bxq9jz0Slla1VPuD5m6iR/KIpUuv8
P6cOQWA/eiJjSbmFVt+YTdrhUzN0e0P41skH3ovYW0yM1bWzGSUOM3k/yRnpwut3
uKYtqjot+b4szPj+wtvQ63XZzoXK+E3YFs9+WEFqQ84fjUxpQ2mpzi+Qlp+cAvCH
iaMAooes9zCacAy9BVHZ+iY/1paszM09M1XVJnHbLSRtzNc6zWKm2/43lYpfbNih
1tUdfNwv1QZdoRgyc7bwKLsZCgRFn2AuT03IoAf4g0SR0a6//E+0qoPwcVD1LX91
H0FyCNIUtUb+0yxDrrTh8VZJdh/e0vsAsmTHOnlJa1SICDtR07PhL2YASOThjnxC
YTn5+cAcjh1Ij/MpAhe+o9TcaJHt/rb0pGMZoyHbfWI4ns5dhwZfAipod0hE3ApN
Sosv1nCGGQgfXbEuiQjv9Ug56WdPWOP6dOkibM0HffM8IBYWtFTf806G/PUIKhed
cq36GV0L2C0XXo/6rfHL3v5Q+fp7SmlAo7y4BrSTaCBKj8o4oR5XJCQLtf9BUd24
cwYMJxJ2dJMBNFgGfIuJ8bP104HXfDhSNOXnNyOWTMnaeourOBKWdPxou7dkovA4
zgovfGMhPwgb0oB95ysd+3CrE/FiSC+uvK0ZciLVbxWphZJtrl0nTPhixuFWxtOc
C8NSVm61BaPQ9sIE1YLNbphJrJPU2GSl/2MGU932ZcZdejnl863f6BrR3sKrd912
UrfiFauZo5UABRyQAKSdB/ePQNGFQB1qWsRoNJSM91p0vigO2gsJ6TqdsRuEYXIs
FLgI4xc3Ni80tVA01d7SIHMSm9MYWRxQDvXSgYbQ0vkOowmZSVkiF+WcEsH1Hqg7
9glJ3xOztGtaXiKLMnfIzLNFRw0Kjd5ceCY+NoL2W+SWWdw4WnrCOFpL+/qt/5tf
KuFVvQPeWHQLIDC5kZe7lo0Uq1tsOL4vKK0enjtBrRojydKqCcT5qAslpmCWtZuA
lphnaWfCBHjrRpGUIiqAI7rkCO+77aOmzSMtXsrNPYt1lZvaEq+xvrw+vRxyg0EK
y1+uCVVdNY1UmwbFoUbeAhc228Hcrvm+hw++LUYOHC6VamErSyDwyyG+tza5hgsK
r7nFA1dTmWufrPzklykz7nenST4z7q/NZpZGYRUFFRqaNzrBsRmNobNJzzLnOQVe
XmQNBpn2dE35mkINkZAgGWWt08nnXPF4P+6QprxaLPSu+BN8pzk4YBUeQ7znW1v5
b8CjBooxOwKK7+pPwtYxv0oSneHoz3QQH9EjXtJEaDMq2F5VjBuI0HefBMN+qeeZ
C8z3QGLE6o+PYbQJGXHBkRRRG6KFfr9UbXsWn5CP/PZk2DLLWLI0v9DXeEObrOmR
JUntpNWkfxJrdTO6rIS8VJp7BAI3U5VEWNEvwe9RtviFdRukxTMMkTlgEHKwvMax
1zi1RzooOgBOj1+GudygQEExPzoE9NsMs5LSg6LfBdpg2xWOPY7Flk/9Zsem04Qn
jqfg8pwBFZ/sxBaRYWlFVYovSYrKKIrfQozNzUrfFHxfdZn0W5BvAYV78D8JtY5V
kyuJtMncKYYAJQEC3yQoCNEIzc/Q/nKwOeQb2IQn75gXnomKYXmwF4dfFLDK65X3
A66BvqfA64vIE3jXcj0aygyFZ+YKg9w1+sEqEwUhFnDbzVHL0ZncGo78wc7QTyYT
CfVH5vfWbxj4YU09x8Qlz6vneQOVzEgvd5SlmOmn1JQsWPYd++/m4fawm7HwMVei
F9ocNF7wJtQl6rdpY5opkcsuVreQI3cH+Lj2N1suMRYEBpHzVY8clRhnRbTSp0wF
V+kYF2x3ZviATjdKSOJJLEx5dYAy+G6OqtwI8B79eTdEHWS4s8vIyZGmV5X3Prri
2/PK2OSJ0i2M5Jl5PSM6XJfBc27sMVuvjXMZWZq3ePp+t+yx1O1dD/tPwdslcCpG
TuIAC39CYWIRXE6E76vnJlXuulhkWTWmdSroe2zNKMux+HC0gpukZI/NP95XDmy8
I73Hv8xlU9QZAu9ohzc3e5GU4L+xis37bZR1GH0RUi0kvqwHm3cl9FcR5p6Yv3Ox
YzIdxjzfL7AEQdM70v9HmKzu4mxVAel+6ijWsf0SClCNPbBi4KijuNVekyJ4ExQQ
RiQmwYreSP+qqi+cA5ISwNAbbdhFkfF9lt/WVLiKZmlDUBckBFw7K1/p7H5XgH5I
AtJtnDt4kzvsc0X7zZ8TaodqF+HhvWx6ocDF73WvNn+eWqK5c4lJT95hVD8+22fx
gs/DrQB81h/E3O0MR3gQYfETCydhQZUPw0ejtyW/3V/Sp0mO3T4Lj2ROlXvsJqN1
B481V7he38fqvVuL8GmZCIOrTA8Ya1xW8q6WD4+UghQ9z3nYl9D3afx6me15JISH
SnfUQpyQJqPFr72faSOwD5Uzp+e2SyZ02B3Z69RtiDyDmqtEG/0KxyLLXFKWxV7e
f5Ytw0VA8oWkmQTSwf04Oq0J9+Kt3WiNO1xgdWaEXquD6F6Hq0vpU0PQ2zi+BIl6
6vOQyiW46h3TCUSJK7X+sSsWMXQmeMCYKRt7hAzWcl4HRDJyRym/q3VewzocNZxh
c+mIxlzl8xqUQ1RAnc8NNJSnerlVNafpnxAsHlK9I0qMf9/tP42U/h/pF4fA4s9E
dgfc+XD/WOH/Q9EwMVy8PDxNFTfcnp8fig3a5nuUoBPwHy1hO7mr+3aA5w3k1gOD
Rp2TtUoXQahHyH3acuUZ1y6HapbNwf4kiGr2hIu4/WzB5vj5gWIAV0hg0t7PtIUH
bFwHvDsYbootjSKkBTMKr/CLzbzqYZzDtVpAKVmZ+XurbecVLDi0Ih9Hdc8fRqll
8fIo/hxAnS8D5SwekKCbYCQk6nkJzAdsTUp3gXgdjGRAgLjDZX+SC3/O1IUL29sN
PFCWhbq4vK9UQEEQNalNZyESBfa15iACO5escWrqC5pfeYARxlGVt6M0UTwxFElK
RstxwULxA+soSA8gCiuiV2AYST/GOrk9Nr0ivRdTsIfvLJJi3cVhzkyPdas5sXQb
tbnPbQxi4hMmo16VftNVzBI3uZvxckucSrD23+frzVMXkdUHyxx5IoQkN9UOrxTm
5ZPw5Qx6UiEheoqv0rd6gMI1YiqTpBGAkhYcjST0BEepqqTT7m1iFmZ/UEuZfvA5
W1f9AxB6mJQRZL9iU3ILxLN8gfSKG6oxY3zgfenldIi4x/kMYarJbhs1Le7z7U1M
4iNX75pkolgxumlQ4GQo0NDVOu3fXkSxdQ08nIMiM55MnmGvJ2IF3iDZBu3Ab899
LoYaee/LIuqCMmxOcSAGS0NaH7hjVNHdx/9iitOJ5rCN1+HKPvD/BBexRnZ7NS/p
7lO5Q/FL4JtjBvH172tisp0u13TNYgnd9wEAhiCOIDNooAVgPVtbgLsJUZwzFE0A
B11eNCpye5YDjLsBhi36FJ51ap2O5wMn9rshYBEKpaMFKaKqVS9vGmM55KLu43yc
fpZ0gtCiSCsbCGxK0ufmSzPWcLdZI/36ib6ZKvGoVPkCF29tNQneRVNTvhcRSLpj
dZa8NqP1quJKfqOm/WsMi5kAV3rYo7qtzm7lOFJrA5pJbRUOET0wjdSLxCxX5fEF
2AUfRNWdDhjlERCENRXaOyTho0OFTDJde4jp+1u9gom6pHZJ6WBNddMbbUSo/Zgv
2nLLyWWgEDg7yfsDJgA7z7sOIeN1I3uKd7TKXPa5LXyBcVZ429cX1HnAzrI0epu2
jkslKaZ/CozTRvDcyvlrwdzt3mMfGzr8Euz9K+II3S6A04k60ju3jHHadRrlKFc8
yvbPNcuJedWpQzzQdcmYneknbai5Afjfel/ty1KXz2Uv4oYJWqpEy0/9T9mHNkOf
X2o1FNEHg9055f2x+Tq4i5zCpAUkDB8blpVJPfHdS5qTb7zcqj9a9txWrZmSusJS
uXdVbg8zQz/HC5j9K8RG4t/G72sDttFpkHc0oD0VAkzdG5AWWeJxj3XDAbwPAUBW
hY7x3bIqDOeqosO2W2OA5VW8kXcH0/MUJvWZ54jaCiG1MTN8bivHmGUj8zWGlUx1
5B8qW6nNH9eH6eB1muYeHKI1gkftqzZVc7SnTuJDF7SdX2pXsIGYbQpswzaF2Zoi
4gyQfZZwhXk8mY7bwGiZefhs9I34uIrTLVoX6/tlKVj3ir4S5zbI83ONjWGeRNDx
aNvBfALFizysopL8gsx20Z8E2ifgdu+xDkVgmGwO1IQGoRSuGKbfW6cfhI7DezU+
9x+wIDmgh8EODN9FuqfShL3wuH+tzB8D4IFXkx2cea8GS155pULC6FVhXqD6Hjrb
Wa4zbVGW0nSAs7+EHQ6Iu9Tj4RKm60dYYkAdbL+r6Zxp1G8qkZP+SkxYLWMHk22d
JC9sN4j8gqIOuYPti1LtQc1iUKDsM/eGAKhj/eNToLYfY35etIZnHTcnk3EdwGlj
adGXTCfMqNqRaXNL2x6ZijrReHOVWs319LEb8gRDcQ6K28JwxKVSRpArsYvDKffB
eH2B4kUnamxZuijHlBY7800EeElTBBTjvP5Tuyc0bxeubK/tphbVgasg69nhkzXn
Ft8s7Xt+WUkXoPrfp5ZZKWLXCfjiCf2ce/rwH+mjEUkjC+Q1kT8LN9y5ff9M0uPy
ce0f8tZ1YWz/lCFEmgqdKAgsb3bKAGbm1VmUST9XaRuCZHD+dfvRW+1lXznawBGo
WI/3Ru0ojrytOv/lDAwDDbVMZt/342Nd1WqX7LCRlfEdIufaNUaP1ZMjBy66i8OE
/QZXRiTEJDVOEQ7nc1l1L31BvHCklHVeQK5/Zr3i03ZAgiNmV5jUiyYzOBZsPSDk
2HlV7kPADg2whCHCkuX9BvFjB+OXcmJ9FXQbcmdnpvkP45PTQgP7SsPu/CBJUCUu
5fSTZ8lXTJ5BlMp9d+Gv/GP6XRZGOX7NLiR/dsdU4lMwiyKAnCEaikwgJaF0ZXK1
4rlj4VLPYtaMEFGb47GOqZDT7FBANqV/Lz8iVqBEoAZazgxJTn2VZDx0RSN5P8cp
OgtHsDR7SHdBxSuP2hJrETtCKq8l0a2bqHWlfZn2TAXaP1liAMNdUgZ7VX+y/M6v
SaCsNlADYuloiIfwXNqTkqsum3+uQLtXPky3vHGFNUmrkkZgfA9XHxhovd/T5ame
y3fam+dRcLn7OE0ZiBEQmQtGnRZTuPaiap4YfoJku1o0YCwpb65ibI1SGSqhRkUy
c2WroLp6h3Ms4gLWR1GuhedAJ2Jb6rA3lk33UrlVPDDfHYGSTo7tfaLHH8jLc35h
ljporpjSFHKbhherjBiOBhejZK1uzaKS8jMCSMu1PdJUZ4QHMUipqr8mkIlaZoRa
2RuM6CJRDk7xOCIco8n2BprZdTdENWXw0tYK2V/hKrqYYWfk9W3DVEYzVbnIDUrZ
+nraB48rXeL8f/+TRUCuDsfZHxfVW99JlOe/z9vZ++cvkYKjJeu/QyCN/4mNlNmP
SYBxXuA3bkvnPWG7v/qbMUhCsexT1OtXh6QlutWh2UELGF0yYZBvt1Z1tcqPh8Fi
GvUR5y6si2eYa5WtbZMn24tkyWKo4b74TEasqgTEFyz2Nt2VvPlVQH/QzpfmJ5Nh
kS76X2fQp3iyj4m1h1t8fdq76l07TdJaXpnj9wyySJwTX+DBSHrSmqUJgSXS0byn
yERbe8IELWyGvq2+j3g5AdajDUQPyjyZMXYay8znpaIVuzRAZCSnZpKvu4UnXaq4
mCK9kI6dE3PDHRDjUpngSR2UuaqbI7CWNkqxJUPweJkigOqutoezLj6rrK7lQ83f
mqxgfOf3tIdCwbJZuZy5Q1knCk4Al2pJNUJNB9fFuR8Nk5FXfbTIA8acveATWO8T
ust1gAQH9cxOrLyH7uqmnhgRTVA+R4AXoj9USC/q65RGd6h3ApggRrcRJvDpPqY/
vUblm4k1lvtJMwduVobWmpC+abXwpwW0+2ujdAPAwClMlsht+qFB0bRwChYU7CAe
3BjPyjJ4VZg/jWw9JRU7aSrfF+5YhjpNRwr75CRniDLdDcMI4e6GOk47165/A2ui
mXFOfmhsy0Wd99/qJOQT9YieRWrJ44gBvfKpg3cT49Mm88/RNHGpHZtLBnn1StSf
iqYq2CkJLRuT4t76l6b5ixi9Rq9h11VMdA3+eRtWuPchTglKnzJ2A3jED48HxXui
7dlg9zqaHSe1ySaElLTr0FfCojnb1cBVmqxoDND+P+y6yPjOsMoFB0QwgS/qJVn0
vYb6H6DEjJktu8POXqV/NdaqXiIRrBMpjn/ORNx1ZUPcDyUm3YhxDPhxes5WGm2w
vIQxraQMzLNdfUgWFpy00ub39WnemPYcm69Xx6cqHG/IoKIg/or8lLgbdp9CdRmm
a8JayFo26cK2KHKrtcs9ePq0xKG/SQV2VwirelR3FvpuhpwJFvGpRwbSyXQLpKWD
UyzvD14F0KZzS2hViKz3Osdee0kYls5SQoAJac7rX1IRkQNJy/jPiIdljtjpykN4
6WZI183wQGSVYDabH5ud8AVPhSQ6GMu2e1zdJyKGt2KZOl19Fie1yrazzmE27KAx
HUT5JTEbpSUar1choDWLyGr+w/RJmHjb3zmoHiWDIu6jjM7K/+9Dg/nf3TGZm5v4
fzy3btEL1OogZ2+87s601FsdGZjBf4cCTss57QeG8XId3kXRfejK2BmzmgVfwci/
atuHs1xBuQ06b/VaE6YbxMUMZNk3QTbQSdpFo7AWseCTenOYrwhCB0WGtPwxyf6K
kUpQ2uvzLQK8sbUNUo4c2pIL1YMwPx0AzfxtSd1AmYLK0hXCGvsrqtVZy3Obms4B
AvaN54xLk8f9Nm7pZxd+vkG9miYFAAhF9qg7aQ1l5SZmUIZx6d01TOvFLm+GklpL
XlM87XiMVcnsLjTdGIlVvkHHPy4qI9FdO2BPC96ilkgHBIww5QHI4vmAUSHhtPY7
CMHBwNhErEGpQ8VJJxpEtFyJpgsYziapJN8EKYOGkV8nwiLZJ5oyTuiGh+HQ+a8w
OhHySf1W0U7fE4HXZ/fYy5ePa+unMkJhHQzRvVb1e88dRnuofxcI1d5fK8j7NGPZ
fnSZldhnylMVxSzjcgy00nSTrYPywsKC/fRNzEMYbN8fdn+mpewN46mVe3n3mgCn
smi6ZSF1sVtph07SdDkRyFhqtybmflDvvd112gG111Bz7S1wFy6LYSKZ5bxUup6l
EE/UiNHUPZh059gcBQHP0OHEq/YKkxj3RDlNc1eJx9RsYGnCafGDGd9YrB4Omwr2
m0WVRbW3iYLmu1Lrv6oCNe4u+9Z1esPB2xgQrAxSmDhArikB8mxcal6vbSTlMU2N
rChanXV4fz+zZjEY4V4sb6MlofCZLblgMyRWrYGOPQhUvsCekTm8rqTkYeKggcWl
75ybQ+OtVbsquQrgvweTF2P9imNHjByQUife7KYEov5HOYlXjqsJjAlIv4+4SB7T
rJwWfwQW9TstcenxjrBNR1DVRqXejzEFFRWYpF6Ic811JY4qGkg2voa659zndlwT
ByRFqx7/0Qsua0JciC4ojhSXAuX4LGbbKGEBJy4rF7ZlQSKSWvi9dI3q9L5YO3Hr
XsHPdY/GUbhm1Ghy8jnZMAJ52AHjnBjEZeWgdavDqlOi2OxboHwlfbWA5MtLV1LF
a5w9g0mcIfLQmCZ9/xKp/f+l0DbShba5wzWxkwowtgTBYtQMkZ6VNbJ/8evic5TP
eyHOSP6dT3B+KzlMmnf0WgcsyvbJ434Dv1uS1zujP0cXHXq8aRdYNkzwjdMMB1qr
txdpUAgX6j8mbYpZ+V07crwlJhx2sB3BEYm0yTnt43snxtW9k1pl/cM+mrmr4KtB
a7q+UCmikt7QTON4KDFAkia0L96J+ud5tjIgMT8FqLCB5urOgnH5TnwbT6NfOO/W
D0PeKACOysn40drcuOq8+J60+J20IsymfTn9TNLKB0j0aVJa9ZA8EVeOHU6g0dt2
hgu8kmZgxgogb5BsXBbD4Hjgl/a1CMam0RvGM1EpZ+6mD0iOAXR9Y80aXL4RdcsV
RNI6TeefCCgIyBJhmMKw7T787lnQEyZiGb6WYrIMIofKLxNyhiDjudaa/gtOnELD
eeOmuMRLxCYRF2YUeiiQG5J3IA3FdT+yNXiuS+U1CWIqHMCz8n42axJA6RJ+GXez
V2fiBQrXRZr3TtQC28dWCoPvwTvJ4iZNPoY8jrl2oxBx1e2cM66yE5jcUjsbSbUe
CL7vEYq/UyYKj8ebbMrcRxgnT/moMMUyuUUCC/JKwNnpFlz7jBARBKgUXpuPzv0P
n/zzis4tw/2/dOi33GBB/Xl0VvOvSqetyboaaObVoCMNbzJgJf/VBGhty68YqSvz
P0bZRYp/e6oqAi1x3tXHndUHVKeqjSCy2jwDGHF1rR3Et1IDyzlhIK3Pa18IFu75
84/s4p4efDbD41hRLCTpZr77WKaLa7sgNeBk1XPn+3r9eHzW/z13wrALkjoV7cv2
jSvRfhVzqL4sngiBH1H1As219MItzDl9pBIdMZsIl1rwgNqM0q5ZoQGPto0h2mZ/
LtkO3pspqHxUYUS4YcuIW5bdmj6UTiPI0q+20VR+uIfbxyNSJ/6qquBpxuRzCRev
C844XYnShOWyTqhGVaQlnmgdc210baifvyW53t52/mtz2x6yNFbk2T5+Moe9m41t
V4gO/zsZR7pgXVkIsbN86yIFGucTGaVU7ew6dBwAiJWmkDNwykbutFNg2WkekhO4
wAIeliCedEG4WjcLvG/uNlcKWV+CRD2Rhe6YMLGf0/z8JwJqm1ilx6qr9v1tAeIH
eQZRY3UJ3GYClZT0lEXmFX/fVSObPToQrRMareHMc1hOa831jqT/3CMJ+brhlXl1
N2PqmZfsHAz3JxaUnG2CvWQUwoVs0kj2zNXt9SWye7+OAhGWEgoMqHK/ltQvo0mb
wE9qhDmykPE+Bw5H4x/SMa9JnTkvfPP2TdSReCVaZqbUasbUpoWqkJIC9D4ZHaNu
r/vpw+HolkjCswIcsFyXTjVrHkJoS39DbPDEm1Kzp9ZkUeUngTSyaQ1ish5svRkN
bEXFSytijwAMbHfx3l/lae8oEtjwPiQo+JF4e0uFPYg6awhDgvONS9pfU+PTciuT
WK5o/7WAJIO3J5exSEZRUaGek5Yx/4KAnUbJSPo83cLtVoFvSRVaC8MynkEASECi
0qhoUz0O8NACDk8xKs+RMxAt3uUQoUaDfBaBnHSYYxWwXcg9otH4kPJ7jXqMo4dG
aCdmSofSLvs/A29psdWSqEcPbYqRg2vu1jUlpWazcxi0JO05NL/IjPPtl3XzQc+g
Udeuy2Ot0rQg7qg9MyEgU5f2SPUcfNEBfODYRLGuTDbcnCIO+OkzuDS8nbI2j/5Z
cSDNKSzPAF2fETCF7NxmviAe4x24X3YRoiNQ2YAEmwEp6j3DLEf5+mmjnn7Lf2T4
hNfMNQinZvswfspAxjXzkWa1BmS8h1gnKdCs1p+xt89EKcL5Tm27eocjsue74T5W
nXyDzj2Le22P5sYalV7PaFMV0KAdypnddDcWbQhTPbU8lQK+sS0/AYu6JJjmG/f6
mkioCQRaXq/2q/nZ59KjmV85thcxU5Z6CjDK0ED0UuFZXu7ijxbn6vODxQU/D5I/
A7HbFIQH74Q6jfOOhLgv6Cv041x6GRTwYSU2ulp8sLXDMtZhrtQsUyYQ2RjwiH0I
5VYe38LXo9OEGiv4TUoVXMzPXgeHcVTJpt6jrKYSnT3x1RKdODUUVpyONn9eT+mD
0JVZHEhuWQvl7lfJiEdPCGFnHpYLk2V+ZpVEaUHS9DbeJ1ovjgrf6Sybj32m3sYd
TwBuTaW9bNGOAZQrtN6Hi2cAh4bhwS/8inLSSf8VpcHpySHDQaV6pbqO0aLrQ21U
+vPvpJ5McbCjV5BJFf3kxEEFQOimGOvfQWr57Zscj/56ncs0ljWYbJN9uEYsFA7r
LzSMLJw6OzdtXHB7MQMSs9zTaj50opjMRimwU0RcclGL1Xz0uogasGDRlN8Ay4Eb
HG75DJyc6dVKlcVWJm9tX9QbNtOgROGq32XsK3Zf+ZoCLLYebxa6MkE9R5eQT/jn
M6diQYB4T+6vOmaOmc4s2MMZ2dnWUCKa5ModcJxjcDRW13DV2q0lIyyaSQndBo1m
mADMgixy+2Wcw0ma88ElWHxxEvi82zJEIRg308RzU2vrFgauXKjn239/puZzdVV7
uHWeIZNyUjFEloYscRU1R/xmQxduXS4LdSlqUhLbaObsxMEZBtxY3AuSaXHBJ268
iiqlOS24S+6AMLrnEQcKIZsaSo9NgKvYw+/cD1+sfoR1OoSFZPOSNOjyeG/1McV3
hKn/OiuBNd4uG0gNuJRk9hX93hQ7H4Tzmy1Ehx0tksuyOKSXYR9YD+iaum8NZZq4
ntMHSoRtX4jCnxOSGsEQ/CRKfVWq69hk2Hc/1qhVrHCu1NmjAm22B5b/xO9D6hgG
LG5znSu1lveaSDqrHDWt8RtMek699XX6N4D2gTjGxD7QNFHRxm/g3FUp9o5s3RGi
pdzeUOpv/GS3LC+TqICgoOITnChRumxUo+gs7s113+LZQB7tAk+/GZBDuaMoIAh7
zOf8vYxmWVh9GC+4H72kO6LuUcux3NdNV32KwZeUMxCc9B35YGS+0WjSrtiuyiD7
Are0YWg1XRcPchqWkeZ+yIJ+ppI87bgKuJWmECQ6GjGpJ2d4bmB+Ka7EImEdibmT
Wmt1EMyiOZvLIgP8jy5/UmMND2CWsJRquQqVUfMgrN7yrBD67sRyEEXen8u2AM5v
AZXxwBRenO0gg1rR7bR2fk5XqrW6pMA2ah9IBgGjrifDhlP6WiJ1z5bjtTWyeYnW
2rSLpwtN6AYj2Qe4ttxOce6soQpPEtfPhM05MeCmZveydOdh8SDYe+mSIK0sVXkq
Vv0bK35ayfz1nuXRbP0rNbWwl39/+cwvQ8BKogfuN6O26RW+wUqYycG7jmHWGs+q
NTFfh3/6bzSeH4vzShS7A4VxCXQQMCWQWseGoEMlW7JixOcXROeBeJih6qSfoSgu
qWuOdD1txCTqdrBqoV0flX/Qu8+onZG5cY7RQv+ZNpLhxxqk6VEInbz4bx8rHbnE
xiZ4Gv+ZOWbAKanQXNCea44d9oRDCYA19wdoOO3sHpZnT+9Z25EFa4KQSsuR//pC
StYpqlfi3BwRTNjeGlEdKTYpY658g9z8YIBTnFh/Z4rQNxcre4ojKjMZ4tMZmxxz
brylgjrMm9wr52k/E11ArfUMQFXJjM/6K9tDVgBJW4/DncsCbHtgqq5BLDAz6/S5
BlotZZ+6IUEo70Ae6CR5WWjFUIo0/rNidlMF4ES34lDidfPVmx8xwuVKfYTTnuVt
9IlZbAcf/KvE/5WAulWs2Xo3gVO/C3AlFGVnMeEgCOUYYrhqwmRELzznhp4QeB7S
zy6EGr48KIw3YP8qFASu1syF8KfrcRYtgqd7T347TYehiw/t28Bo6kQHLaPKasU1
zeeox5HuXcbsiI7VHN8Nl8El8KT5P48WsIjhFG+1Yqb0tb5ENAw1e7mGwg5BulDU
mO/eAG9y00Zfk2HUeJLFlKpoMMa4jb9ak6AH7NTXcnUC4B3b39PnENOaxz7lw5xe
IQa4nvTVEa1f2FbUM/pnNK0MInJbnYItWQ82TXiLPsk/TeQeaSh4TuISK25CybKf
PtGHIbymxYFAF39zEXEbAaLFGYqVO3aH1C+0xBQUOzvDthz7XZoC+zvDv6H+gCic
ZFNUANWYh+znJ3bUHQfE63DNIJ32Xq6jo5sJ22trWcOCl/+evRqiBr+kFb89qtY+
vI+aYaQV2WKa2D0wqMXxG1S1ZJvk8IMvJSJpP2NbehYyXz7P5yByGaKCwosrXWQN
NcxEAu9MC9MtZVpoPg8I0ClWEXucDW6j8agd/tfzaSmm39X63bJFpJw5gRIXwFIU
c0pp8MxceZQCvrwcHpE5rQf5MEL5D1Yf66m05hnmuJCChZG0jrwPxPvB0l10LL7Y
Kw6nUTZzglGMQClaDZQ5rJysIXWlrTz8Ht7weOdqxQi4y+k1uTBXWbdK3EbkDW2o
J6Md9EDEq0LeyJrEoIR8meS47QUjDzObMzVDRyWjfcTIgDyywPoInR3RoCxbTZde
tj+yeWALecAFafy5SKlgQVCldctoV8sfKZmvKGidtXuaGrXA9hdBv9vRZIKk/DTG
ECssOHaK6Z1/P1gifHJMCyyfETA0JgvO3Gr9lFfWEXffbPlBotRHR6L3XBC/nA/M
1zd64JDe2xFCmlCAQKTD8Q9yT0mXt6X9cznot45qDtx/nvwXmjZYLkDeT1AJ2EPZ
ez+5Dr6RIJb3D3ro4F+fZrvqQ1baJhK8ILC5gqu79BQ1h1Z9AeVj4Wzzfs98yyRZ
qRm42PqutIjCjLFunJJ2G79T1D8i60zh9aYZaVuosf3JmVxYDG45Dfj3sBQZC/4Z
0Ff25B8NVX1+O1T3b/Y+6OdObvupiy0JTSsOSA8KCJNitL0TsYl7bfXADOaXO5G8
YCkqr7DFp8WYq91LS/lVxxotL8eryYV5o07SX/aOKpoMGriSc3FwgpvcHTKJXEV4
p9Vl9sHoeQ71pr+mUi67ppSIlyi41H+EfNZ+XSi7+8N9fZ5qYUWXSfQyLH7mdNyH
UAgz1newf6ghZi5LnEemKQjJOBhJeIdwHjLDwBxw37TBqEE9WELyKdE+WfK+SdWJ
KW0pQLqkhIrRtlaFiK+p2nI8mLmjhXTjAEb95ytiU+JMvChBQAJ7RWPYt0ZjJIm1
rRkn4ddHjr9yKg6mBD7R84PxTj0u9Al/Khe6Z0tbCpVjEFF45QicwA8d0wKb3XZp
+SrqolaAmvKL+Mox0io22xvePVhkQVfj2+gnDC+pv5oo9cJjlS302ggEA8po+Uoq
LLuRsezLpEWfE6NCugk1i5im5kVj0HavpL8MnBkfdNixXGcirJdKQmRv/hY5JIAl
W4ClTtlhRTrPYLHu3jlQuq4DuHn7HmsNee/9hQjPVIFWC5Yn3VicZ9MUP+bsayMU
7xA75iXBU4RQjebH5uEtufj7kHTKOeV+pcpU5hoLHE1DY7ee9LlJh5NM81OcH23u
3PKT3ui5wnCi0ziZFrD5RcO5k0vgTtKC+wrvwEhX3EWRTwD8CYwA88Jw/4y/4hdn
WmB67H6x1ZQTZ8cm5psTFV2nKqCr6RLGYmT2vWY/IKCmimjs1ZaQ/ObmUMavcM5v
LxsGl8SEuvYwKQV5w5/btaoeySGw3gCd9WIsPV9hWiGdS0KAzq6Htz0gRfEuJpkt
JmPiZEPOrtUblpomdGacL0WfE/z7MXPvZIvDzaFimEykUSzIwBadx9fOso5aUcZr
K+Gi+TswHuhMPzKeGbyXKuTUhu59pWyTiNE+dQbvfN4G7yi55Yj1lh3IV5dgjKAE
5+IFYgB1GRRfSx9pUTxbPcGb9g3jZIxP2/y4SlUVnqFxyIFe5hAM5gZEqyM2r4li
knKQea8f04e0fh7IJizQ4FzSAPctQj9Q6MXLGIYpmGV2rpn1SxggzhlpI7ydE2Nj
TU0BHL17Sf1+IHnU1J0gKnq/IBchHxqUq2pZlJAOTi3WPLNo+ZunbH77ukN62Lyl
FzdJN0pEUtoVi7dYFLTxvu5IxOB3gi9cApFvPtX0SpwgczoQUZXD+bw9jwdr5Wk8
CcszNPqAsLVV4hEtoFqdbsvt/JBdk3zYiGdkvgBVpNvtyUqJ0SuYG5cXx74JqXKs
t68OJAwsxo/rMI6mhYZ2rZ/b0EW4aehqaRV6/tcoqCz5jA3sWbaHevL/l78n2oAC
cUDOhnuHtm2LfH9/Fs0Gna7DK9m2QxSW0FzeK3R3m0NyHNJcK5ST4wVK8/H809uh
vv/VER25Rdu17rdRbJf6IiXXC8lwC9riZAuC+8+KBUgxp0g3NpyoextGkdigEwRt
mYRkT4GizKfTEJokZULbHq4q/BZxWpdG6ytmAUt3AXSHTtf9UY0EudmvipyMuXbO
9pDELurggFW0vZiyPK2b9gG/HBNeIRy6hBAntpcKbWVdJhZXuHr9yqI+hd6figVV
1Cz+720oFLy2wpA4Hfpr/lbJVJUPG+cIEI17EFopKbGNsqh7lmsRyzo2l92JA9lI
dRGQ39CxPwWJOf7Xs7obyG1/ynpPj9uvY3flI0QIFjH3E7O+e7NNjNUXRYddkpEY
erKcPvffWvfgI9fteon3wmUx4SNZgUhDXBDy0zmZWHJJeSS62NeinbB2AWaZwIvN
urdP4QGop7hACBuzWWqBx9vMuh7hadJoh3CxlPNybt3+nGVmNkC/iUgezxj28Mqd
hFNikimEi+Qf93gY0hHVl7GEV29/ZRrSWVjhAW499R7ZZXSG5BzVKj46ICLA3xup
wYz2ct+2Nflp/xIo+0ErIMepwZON4RDzEa/HpVSt8hHb9Un/1lofUySKryB27TAl
25MnqozwdfF+GJD5A3l3FHt3YBMq8vz343UxvzDAJGmfXopEGw0Tr/X0HseWYabh
GuO+1EQgu1IGk/VyYyZNXlYKoOZZxb4jOfobkZ9ok94m6iJUeCNUWV1pjzrCGH0L
NByIberk5/AnIJvp5HJsqSNoo4aPhrvTHcH6g3NxGc8nPMrC54jv6IppJnuqSNEB
5KMPGOxzDnr/9ZlMV85nfEvv4jMVbxo1R0+7t5j8O3JaWUI7N7+PJztxdI/qp3KO
3nbN1pHcLhYTO0p+uCCjYotkZJKSQcctCVwbK+U1UuST/QMEDWjaw07XtWMRTTHd
YjujBGO2SZxbEZFzJwRVvhU5MYp36qvZz6KXsDCxKow4rmW9uNqXjp+8fzvs7v1b
YyeQCBlahDjFLM4DqwqntyNa6PgPZbT2cIVP7uVPpYtLJPpW5wKrJ1aV2FhEaJPy
PpGF3AMpWpcy/RplMKh0oUeGkduuls2gJK152xgf95vBppI8bk1QkumSYLZtkx0d
gWP8IGiJcuZDeUm0d+0Jt5g/QXZpQ0g5QYGXW+7au+zQdshcHPfdxb9HYtoco0uf
0tX165tTXitMblgduB2e4wtfbbvKuAUveSxJJNdQrCQsLtPLykfktbuBxewDq1Vb
E3x24OGLUZ6CbyBHDiNcdvPoeG697+kRtwROrnjyr9H9WRGvZy+2eZSo1eE6/Q+Q
BWB57WGFJUQtFPl9D5xLW7/EEPAKf1aEFS753guigFex+7tO26EUEM9RcHhCSaOP
KRviI27Qap1+eRCxbCByx5+zfK4Ri5dHpGlS6p8LMw0gzEwzMwISKMp6GXMPtQR5
RFBX+WSs3icw1gthcXXsHq3uw7cWiHekGp2pLAuxAd3JJ0COVsFjUOyCEI85nMQ2
ONLg6XMQ0XzG6nA/zTnWRAn/wKfaxmpIdSAT6AJygj5MF3VEZ9oVEHnViD9sCtLc
1lnPbn2InTTQW5y2V350Tc3ccQEK7sgVeMRqaSprQTIEYe48daXX6nnZLBdKUoL1
4MlhNfGYK8NgAJho5a/14hi28VZ99MNFI0Tq9Yp9iDpQEdxhcZGLlYuAocB7E5xA
B4IAg4NbV7guDGBPCuEK4mPp26PWZyvqQFg/ICOwFWJu865Xg+vWUcScJnXg00pM
nmGQM1zV5OaLDqURorpXaLFt7LPwHicVRG541dMPc0w4SEjoy17yEqvzwzQAf6LE
k2z1DpMC91uWBfvGxTd2JTzNx6+OrwrdAa2a8nl6+vwKm+O1badZ3iEVgwo7n2Ng
WOvD2tnpYZ7FMzbWzE+Zn7EO5C26e20rFwKLTVtEuWdBgAhAW7YDmR8by5pbN12x
ofouVpnkapfObYMDCKbNKM4h7Jnrvd1HiW+0Kkmi3kVqwpw7jha80JbRA7TY4o1I
7Sev9oIUL5dA4Zgd2foKQLz4JG8pQNvdOxQUyQYC1B0v5wtc2qMGaV6iEObznKnl
lkAbzYNK7Q0wkw85Umz5AG6khZq5g9MPKLUxbINKQu8U+hqVPBZ4/hW5UYYlkT4M
ngdSe5xtQaknAJmw7JLiAxqUN1civwIkBc13DQ3RG5hXqjC3ydI/lt9SmAGD5Mjm
E3MhBmOhuNA06YV0OVz0G1cLsIRecpQFFOT8hnY1HnFEFFg7YodSUJI0zu6f3Epq
0ZBfJ1SEgJUZ7mlf7egZj3Z3OeVUo7MR2+Sc5tnHCOlBw78OMxmWXoQEYHvGMq/U
zfIiPT854WYx8xI12w/MDYyYCGf5M2Zp9E+D7mVjsVaCv3HDwRxZ/pkIx3llDt2P
Wy2Mdt7L1eBA19FtNrgv35Vn/ON/SgnMc5w5bUtkuPy0NprF7TLUovQ1B7qRySNn
vxmzvZdWdSRGIRmKmhbE+JO8N+XGLmliGzqg1LcSU4uxVYKbtLVL/MSgTQA2ABKa
x3E9oaL7LrfBILX/60X22aDSnloPcf2KjBoI/IHgn6MsPMwtue7Q9tcJg5+RE1Ol
JHeSWEAxPVrGoa/SiU2EKh+Hm+3HWgW+UlkawhmLx9RLnk4YRBbs6XFvfk7osts4
GkD7nvUNPWKF5CvbKY97xr4MOaVuf7KCFIgJjYeix2AaxuRL4aKp3+XS7Y0a785r
A8FE7R6Rf3f4QIegSFOhQe/XtwtOWCV1FRTCPtsFrnimmUundNasiRVOHna/wf1c
b4veoykndPl3UgJ+7KwO1SlkWffDRIEWMRCtRNjWJi4b0Bnhg7gHuQMRtB5v/yhB
NSHp17t8ue2kR54AvxsxnOBRL+9Kbj+P3GN8DNQidLm1LVXc8nhU+GslycJA9RKZ
jgclY39n5AUUgCQx/Q8Ix9vYpqFv9zkQwbefSaB6hNhh9igZuaE70odXorOtas1k
fiiphAe6L/qCSZN6m2TWh0obzZ9wfG18jX1PGVGAz4UEYmE4kXuBesM5wFfeio+U
jSv2WBo6UdOKaaJ5hGpPyYH+xhDUmwkXj719GrVpENYryaRw6f/MABYlMhC606FI
tEF/9yYTKcJrO6ruh0zv5SPJUO9PbX5nZ3FsiqrF4NDX2oYBRO/J3S/+gql+MMGj
akXSU0HIU0OU0/9HgpHXY3f5NhgjaE8RSL/qfWc4eu2/8dQbgRR/pcCUoezy0bSV
wjTvdeF9bFlxsuOZTghUaajR3EyRujBzltPfh7lxkP+xwpQ+FRuu83+ZPEYimAee
zphbqqDurfL0C9kYi0PxzTe+WPEGRSDacoClREkn8anX9zoahUps20TPkI+ZmPBN
3cA7AZuKmdy6pIdxcivypBXp4kx7y7SibWHaVgXfmdDJsHbCeiaB1z/HfNJsd+Kl
7nXraq89S6dHH5nhVDL8LUnQmi/TK2f4+td+bK+AYzXf/Sd2lmPlBIj0o+9B5U2J
Y3iQwCTY1ZBGqT0RUTwbPKS3fLadqh67M5mPF2+nCGMrDrLc+hgluz/gyL7wYM2A
KIZSrTB/hf8GF4HZzUzVEz6QdUCq42CbRB33x7AE1sPjzJB1KOP/V7HqFmI635Yr
MDLYqHyZnOOTwbYWoFgKHLocULsbxw8CC1FSkQK3f8/WceCflREC1fb/OsmQdSdC
QId8QX7Asqmf4wCFmHwDql5ILd4SWBq3FN6kMFiEw0xzyPQMCnW0FxQVzJSeKw+5
DqBR+mFYik84BJWCM3ayC1uuUvpjeiZJRsA5MsPsSouR7hiLm2p0p/TgMD5LuUCs
VI8kJORKclFiztHameFgwKqV+8EwGgRz2ROO50O7bZvBm1s7Rvqw15iG+iU7Suyx
CzOu3EutIAbMJyKvumArX/N/Ax1xqRVFzYFOwEDk9UuhY5lejWrvR/SCGn+Rh6cd
uYQk5Ny52Y2VsqV+5LMnv9HFlVFUC4+FHtXKInedzJVci7uuFMZ96hhMaCMke43M
CMpZS0nAR03TrhNXujvPqCVCufUZbLAx5wcX0dEqiuIXdc0sPc1GKU2dGK3aEa4r
bhfbc/TKBGXeUSFo9Dc23ShiVJSNWy8EkWwRwxhIYB8F2ByddTRQUn7fKs3MZzrg
/OnPKWPUK+zauH2d9BanZ01I1u5fK74sYqPlQVbC4dvbVwEtvfUyeEXHD51LhJTS
FRKKW2UNgpDD3izFOBEuObywYtNLMYEwbiRyywi+plKdVPUDk+1HoaRp/+sxkii+
rgNrETpr2j+cNogUhh0UxxXWH8RKg4Svy9U2icthroU/xZvq4e8zvWzbADADssDO
w8g7tWcU/9Bx2kkc39/XUqpnd8i4ZVhqdRntMVGEz/5UPi9XEA9OF6QivQkLUjG8
fPmnGK4+iIg5174MHw8b855bekTkD6eueKO9A0/yLBQZQklSf2J1jsXSP9shy95b
POVUAlUQVrrUni91pSX7TrlLIw1s//AecZoGcBKmBqGLdGVx6BoLsHvIjnU2Xw6e
+eVycrwpwldufNNy/UKtZEpYGuaCvgYTWOwlG8oVATVUP16PW9p2nmG+oeYSGrc6
PRwoNPmcWMPtbquzFHF26tYC7anu7i+DRlFBOgfMcxnog90xwO0iCeiJY4NX6ZTz
XrJqg2CFFSIRyJS6+CGpb2IzeFgFlwCuaClkfEYACuuTbTzpQaMqH+B4KnIyTXLB
+ZnVemv7RD7EUBnTyV8InhOQ7ns2DXToqIjdjik8vliO7vnW4sim60V91LStGbfP
wQDAZ9cAZbJ5ndS6NMyz4SJsx8h3bTKPYseE4ztW6lI/C8Dana9SgkbE3oNIvVIr
duGfWxAfM+Asq0uJa2nZlKyTD28sl3waFB+cB4+DZZhUyrge038iW+63vGaZHjbz
LNOeqrpmpcATS6LBM4Cos2+D9WKsDmLeFs3UxkWl58LtXbdiGU9Fgv3Nx3lmWZIz
G+DBos/sSXqu2Kud5R+qx768Bip3p12uKq1JrKvXg77xG2KwJRBLEMeSNaTuK9Ze
W91RLRdonh+FfGZT93yFfso+FVvOecAf3GM2NyL8Y7It1VirkqUQpoLyJ9pcb6AE
YQ8VT5U01qjb0Ktw7IHnTXPQ8ZyHikoOi2UkFp3qsBDJswQx9InFV8b6oo86NYuy
0wIQrLpHdIkuae0sL1KG7mkf8Yw/9P48MADwthTa0OqHcp1xbGpVBduZ4uG3rrlo
ib474UsD5cKNDRonv4/Fxl0SCcVy5pZvA1D1bC9Eou5/6/he5K6o+wJkhtPUnJ9j
W/Ayr7DqCsUcJDl59qWSBfBuLTZ2cRtiUkrzpXIjqGDZYgpPN5dlFOiXtkoVw2YI
tF4CE05HM3RlzuzJd3vkTLBcwuTmb2EsJrS2F/rbmDiZ/7zLTEyoA2iNCon6UgvE
s4vpuxc3kIvacHIJJcFTXC5KBfuS+GatUaQgLXptncsEV0yveQVTRykfNbw/PqHX
2O4zd/zljpVo9BWCTXtDoxmmEXTrZxveEKTHOhZNTYCin9x/Qgjfj6xfO0LGNhC/
tbtDpTEPI/l0c2COACmGxfvxdod2sSWACUmdI5nACnv19fxauyZWAKcH43trI0df
zKEx/03lgcSq7EM/3zhe5lEGTmYAO7Er9Vh7BzLmhAgUZxHZXQQz5ubFOGQicl2t
mF7rYklMT1gnrpNu2R41NvwBilv13+cmS04SKN1SItKE92cpUPjNz2ZqP4lxgR28
ghY5Ch8znZLwP0AakDLeZQTxbKFPha/qeerXgTvaJ1h/OsmZklpcs9e8tYectl1u
qDv5sMDHDCvA8peu2ZcXg055SSgO5TQXBnfir+gVabAZHaz6X9d2CbKVWY9+Jaoj
GR5RzbUuvN0g74irPoOinuigxkCJ8UNpkXO4F2SeVDKP8b37lr6kdH1f9NNnMRLK
Gel66bC1R2Pfwi83g0xwFk75Vo+itZ3m0Xb5ieriYuU5VPe852K+i2yCE6XMNz0V
oQVX/d3ELKfflTuwOh+EXmxuXEBOJrvzGCmBEfxFA0WXIkVCnolEvRtg1UaM3Gne
JThrDnFXqRed51bDQrBrN4NP/u3kQuIHi+FCN+eRgKg6MAOYzV9f+FNQJjApgDRo
faZC/NiETTPMs53vdizjPoIZiJGGAY9O+kWveSg98cfvTnnTvOBDS1c9gZix2OhL
wNWNrPRVNkPHA1P30Z57h2NLxhnCIAM0yangKTk5PfxdIrcia+tdMCRENb7fLY2+
9UypSwcWLadVYiW/M12K28Esjf6Qy/wANliBO/AT1h+ZmYKZaEOkN7Mn5JWZXba2
VJBTZt0LoWONrEl7rnykvLG81jdkAZJeIZzFcSzrH4/qv0mBjKSWu8VDjno8uvHj
Vqwvcm6sr06BA6eQ15WU+4ll1Fo2OudsWNDtlKRJa8J716k/RnMLEGiiM9VN4ZKk
MDOiNy+2CQQ6dPvKQGl0IZtWQSn/ONqJZJIKNrkDGnkdpp82CyAApgzieY0KKAHx
ry+4RpRVTs9FOOijOluJm3Hv5OEszQ+sq5+u+SvUmYT4OA3/e7vnbJJ88ulBOde5
xqXupx6EvL8SoQW0ji5YLycZI0ter0mnjpMHTwHUyOBVOjCNNBWO5uTW8JvHMYfy
j4mZIWkOOVPOqFcT+wBT64aSMvB11Y9IDmoE+7tBohuvqvCTqJ34vDaRwzWl3dVU
+ceKCFjViZ/RhYGLI8E/ZTunEQHHjUQDsqvb5rgRo0ZG+VJFDkBPyyEcfP7uZc10
FSsBC4xAhRiH9rUl+A0zhOIB2WRaGlxaN6mtH09z4uUpkZ8negVTpTvbNZuaS9q2
ZhjusFwfu4MJmolmSrIjLF6h7SHjKEGY5km7ThnmaCg53hwihuO8yczv5qGubGVa
KkPO1KkFTCz/cMPWdkgSkHEsxS3QJAzzHerVXA+5UILi08OndWAB1HobZ6amyPJe
7we67Mbdgb15uftegsRr0gyZCLjcaFGaW0UFsl60Tf2jq1Fd+25GgREWhDV2I6Pl
8emr5ryrnEV7xdf2/D8smt3b8k8qIRTxx21EmWSMbLTuMiDiKlX86hfkxD6473Qc
1dnriWkQJ78vnIosAK0ewlnGc4vmFyl0qxoWzQ/nXXC7lrlewLPqbEqiAdRgUYtd
jxQv0uNLc/I/qMSgviF9z4bvkXhgZFf6jke1nWSicUL8B5X2zcakYErYSJ2pRhxb
I6wBh6vkmIzqw1HI6qzzpbXi7k752H6pmdrKKSj1GVvcU3qMCm/j/PD3Xm2zRCGr
epPQ/+BGFu4LzGZB6fwrHbM6fbQySBC6/Ok9x2LleK5NEMrBr3mT5eTjc+CsC6pO
MF2WQzpl/EFH6RF2s+k6bh7/41qRF8GIK3R7mROA7xAWzrAH6eSR4qnmq7q35f1J
lmH5377udxqrwbyxE0Y81LvuzRHXKzp/t3IVB5Vc9AVvifasS8K3ACClziGabp23
MLhic+e0Ic/XK65oNh2xQr7ykrmZ/osUU0cXU48XprEye7hUupN69foGarf/0VVR
f0tnaoa/lLTWBacTrymmNRwO94jF40HLqFr2dtbf+mDduLipvowRnWhQuAx9zgMm
bPpikMFempIRHhc7Sei6pJiIHZmBOz5/j+kZhito1dxM9kehmK9fN6P8RINdrJ1d
b4GSQ6WDW2PtN1w5xv7Sli4X5NJDKzmO7CgTcpFL1iDJNO+n4GQR3xZvIJWBSQcF
HvCar3PpXyDS1mOAdRiWKC5oGxDp8lKT3LWq4VUsd5dbId/PrUpHrEnPpjf4GqoL
TijXG8MI8MDfll2kbIQExdvyRgLk1zHNWsRztdcu/jLjDf7eQlI08hO6S1qnqHin
nf3UlvV8x83VnlQ9kZxRNBmmPLsi6N0xijGhkIBj5XfkTjIwr2Ge8ezFwmIK3ap3
R6djS+d2Nt947Y66toJoRpoHbd+4u+eZmanuwspI7usF8nhhKm5RvCiNRuyo0LRl
PZL0tgFIWcn3DMu+kMYXmPzhf+eeAIwji/m0SgD/jFRP4ayEc6LptJdKlZB1dxSD
Z9qljswX/napTWMMp1TY3xXo92ynPy93VhgLLJnpa8gjOQmdsDwntFDQBosDK6O4
UvaiFiaaY5OPZaDfJfk1aa03CjKquTJVsmbycyVCQ+Kw7wwqj7+3SHoNUsf77jar
8BfzTTNY8Shwy3FeUglPf5rxX0MJMO2XGtEfnFfxozSEq7eFSsnjprAZZP7hcOJk
z4+/8bFQEVF2OSVzm77N/Sy420dkG1aa0jSi2Y3T97fsZOZeSJ96o87RTQNbcIER
S30QVaeUUAyGrfrN9slit3jlAknety3xjo8C/s7jEDGq78qfyYZ7c/sFrSx2iIrt
K8lu+onoL8qn7QBjxejf3Z+nT9nPAkAdsv4id1EP1FFwz746wLTyZKgaL6jaXDOx
AFdvjxetJVgFJ6JE+0pjgo0EU8wuc37CvULylHzHF2oXs/Wjna9Nx/j9Putfv4Pr
PNL3EKiv4XwCRiEEm0HZTcGZ5mElaPkye9+Y6NLDK3OXRdebG9QwH71M8tgW5ce2
C4b/DaVAtFfdfgVx/WMhr5xjbqaXQ9xqxJ7ivgA4G+I7GO3Cv4fbP8ALwsAZcZUB
+PhiWyMhf8FTrbizVMpAeM0YUHkdglJ2V+eIDBMW+sBAEoy1n8+xkc7aPUQXKGqc
uesSf5ECRHpXbI0zxXeUn5XzOyiij8kAuBxSXGHWPA1T3b4hZGfO2rE3QoogkA1m
hUkd3Tqc/aEwJWBJDunV1o0FG3br28qvFTKX2Vxx7k35OnmNSzq5PGbrcqun9UGA
pXyCnlq9u4mMoGDW5yMEyTBSBhqI7ds1hFwkVEox40f/KwoTarZczuhY0708qgJC
5ZT3ax/EPgdxZCIjlcvXnLVVw4y8y3KSq4sVjylj4j3THNBSEKXOU8KmJULnjXx2
PbJCkM8nPdM/eRa5Pau/4aY7iENInycfid10X+vbXuaBKoOLqjQ3WdoanT8QUT38
6f0Np7rm772a4RG5bCQHafMOiuqa3wS52Qi6j4htw2tnU4zrMaOS4k/QopImcjW+
DCsGlUhCpsabQJvf5MOPdNqgZ30KmDqlm+RSMmkVvVzUD311a2Y+So7/q/z7fiui
T2pW+3I/R+hMSwUAIbcpmiF6hD9iTh1OZaAny6RuAygpAD+WDJHw/onkbtBJofoV
51kJql9bHOU2TcLHkwRhP3wvEnFCzQBWNvljwz+irG2uziQhJYd/vf7x0T0iKLrv
CsMKxRTSvqHr+jKEZ3jd93vVzVd2uuEdOx4DFjXEw0S1dm/gol9m4SZIN7hc7Uqe
VvZ/MAmKNnB7ER8VLm1ujCEqXi6KCeaaykQQnMqvIDSayNk8EX0TbvRm2rpkRxNi
UB5KcmxiNlkvYFtiXKKID2noGLCSXMLa0FOuJ9e3Z/+mD+XZpg+yjRmaMZOTanaC
8v6fVgaAR/Qzsznisot/3uc7l0b4ruqPMdjvjmoxwYgrRK7BPyr3/h/8VsUpdhRA
BpNH4rZRQeTsIMTUhKuRMy0EHSVFTlAnG+2HXPOjHwZ6lZlo+DbnAGmjZ8+pGJlr
CgJB9nnDuOhg90xbQhipCXl0CNMTyrIBQUfzKn9vPrGMk/TE1hNb39Kf/tdvfxrh
9AMXYysMF/pxSvNwztqEdSL3GzkC1VCMozTgo8P6m5EhuMF1CLoQTyEX4fOjYHgz
JpB/Bhn9Yq9s5pl6AYKvG3ayqX5tKPhlzMo7ob047ntm2GigIonSvagvKJHe4ArX
5oZhpvzQHu+wli7NOp5Y0NAzlWP5ZX8oQYjfV2VwBn2phGwGw7W/R+ofbhmfaAqJ
W0Pve33yRneMTENGALGTkjF16NKVIlDTvP+Bjsu44xG4w42myQofL+KSRBHkgtyr
a9lSIkRY9Tiw0KGhyyYVX/Qg5MVmXVgl2lvXXATa2ohAnansMQvZuOUNwI/lTsw5
G+Diz5KayMfTVZ+Ll48s1Tc+/qd0yHnaFiNLDP9d+k52/BuqZYj5/EZd46jF0MQT
ZCsASobtcQSNaAYvI1ZhrEYxuDUxXGNYVqezE/wc2fZIm0iU9siaWkunMSQ+tCtq
Lo9RS7HceihlAEZhXh6g+CX3RpFBCUevxZzFtYEkOqwiEUGBfZkk7GbTW2vh8GSS
P2qVTkXaBz2xNkmW6wKWozSzlB/ULTWQBcwb9gElBgjW88eA6J5P8cxz92ceLmdu
LoWbOWfhvYYJAMrOR5CCP70M7oKQf6CcOCJeHDK5ftslVLsK3Oo+g2zVw3Ffh+/i
1Tyd9bdD+Zish/CkJQENr0mzmElGv7GK4Z1ZEgyES1fGL6waemt/81W27gVhuw+S
6eQxiToB0bNdEfww7Iv5Qt7j0ZGPlz9Gxmk/ANvejf9qYmc76aF1wEjKE8R/e+We
jFOyOAgNnXItTpZfRF0KVVMOKAvBLpRNb23ldtnTOI4HPGf/pCco+ZgK7+OSqapN
PpAPfVkwRJI0lAfUbr8ByIU0gokBCbANuUAaTDm0lZj4bldqeNeBdZnyEhebdzF8
RPGD25p5VzEjHHiLOelyJxdS/4ePQuPmWWwvBnNLS5ke/Tpw4X0hmhlS37GVx2wf
QvENhMBMzTpnKMirkEO7m3pbyuO4q7FsabhGd/crKjvQA8d8gIlD3lxrdRmEFBU/
GfwzCroKav8+tsWpcni3JVwYyYNJ5rVahc6dvvbNGBvYe3qyTboLvNirQhLQ2mzH
3+hpsDb/q51lsJAMCUAFpkQdCDKzxD7SiQxhINRaHeAybvAuTIyvD71x23sZN/Dt
t17jlEdKNjKwMfQJ/D1yfv1rr7hHO1+d7Wpca3u/sOzj0nV1+7zCP34WKRx9M7UR
FrsWFTaW9uoTn0kSEnc9jzNll6mOhVIhfgvvkNQVDdt0HkJyRh3c6rhyzXOlOyfZ
qVrMU+tWDzQftSnj1Q5QYgZGyWBPa1WdZYrCOXcIkIT+FliyFVWC9ZcDm6HWSveS
jPEx+VubcRuV5iwCLX1zpDyS6+MrO5tULIgJ/o7it3kX4YPSMp2NpbHYOXHp/Z6G
01EXxXr6CLP/Qsyafhl2dTd0kD3Q5w1KvqTxRpc/ETFP39hJK+RScPTnOZzKJcOI
icCbQT+Dw8ZOwYhfS742o43cOPBFKW0FA4shzKeyoXIei7v7vc8gqF3+ZhI0rGTM
L1qkutbbzRKVJOPZeOPpfWJme/yuXOyCrTorbPKzvFczxm99lLu4FDOYRpHbJYkQ
e+nwrKuhMMTwISJb8tb1epWSIvYdfdu8OTr/j65LVoC0VPvunCFCzc8HMf+i5Hod
IiIYCfW3SGnyBf/CNpQ2fkMfxuvKZ3bo/gFQfniA0ag2ClnU4h99NN8gx3DTWBuT
HKQYSi82YT8TyhtA9h4k7rKtyjhY/rh9ad97L8AKYNZMTkRfcPztrSdfGJzSU7gZ
xReqe3F0cuL4Wg+OXuH8NNO2JDs+xkr8i0kGlNfVMvE4BE6IDqPk3dUeJSnwuPqI
CYR+G9/WVEO0fXbqR6LXXnnyjAgZuGxg156vhUNIMlPE+0c4dz06QnEw2P4lDxyO
OyLYMsBaOSRqCnw5xOxBRtUYg6J4eisc0OJ5MWEH9SJFaEzw33dz2zdfRX7uxYw9
U7mlYOtBrzBevEMpUFaL4ezoRIPz+6qAgZfCbgn89hN6Q32jI165HclTHacgswJx
HyVcVRhltt1UbRPwOIWG7E50cdXS0F0F0sSgjZIqjxlG+ohbGTHDHYPdOwNMpjik
xT3kY9byjOQUxAqwHt7X2RsAzs9t3q+zqbjRylueoEEVJLdtYsNrRCIoLcSddER0
q0oUu1Vp6mw8dZ3jUEaJI1V8NL4kLZw0n7cA7jLVXEdRNK8d+IpIuSBeixKmlYvG
d5qdyI5hnqeFO+yU6Q8ptRoy3D+Blo7qfIDnI0wwvdXnvUiyPpJeiajCxwDn+N8Q
7OYUiSEOOLMuR44q1P5rSN1C+sTWK1EBQOnco2yfgDQ4OKYdPGy2skE1QyztwMek
nvaofcki/Y6FUsMOfoU+tafhJybKIQNaQNxZ72tucjYYkNmDnWZZGAWWYN4CFFdL
dfQfWPatIlXMjZQuZnE3JOPuS2UMUCoqVxAjcOLJv74oQTGJh5FqPf/1vFqkxU40
pvzHCatPZP2vn69ZlHkbvTWt66u9+uF7fzLF3DUgDv/4F7qNOaiV/Kv6Svu8AYuW
1cGcRkPE86Wm/XQuCzByvYg3EAq9GWT+MWf5eaLLJuzvp2QiDnOeOp6hsyiXwHgs
yqDG+afZCRjDSNIOmaQtNFzuZ5p25Kjex9Do4gKxxYuCTiXji6x0YLYyWOSudjuF
+TehSl8igiCIrVfQIPucYuege0LrR5YtqmUBMKcJw67k5qewqq0Q+f4LcroFAHKt
ptbwpnAEvahwyt6Olg1Nhm6YvOcUtT3Qa2vUbxQhmkdVYREUriFLX3BsPeF2ULH1
6qQ8OQ9mvf3M9cUY2IQfom07ROeamE71dNWEgnJ+nWN/jIFj9VF3ng3vzrlpHhru
nmGHTXziXAe+CFPL7c+22J6KofejaqjgPMbE0dG1olFZPyRPWjD6vywWVB/ZyX11
2/1A1QGLeNuwAEKZOzJAP2ICPXId/0UKwrIkHNQKkL6Ii3XhZUdD7KpsczxEsY8m
Xdidijju4HswFNSBVaB2TwYOFI9aSQM37EqGtqPs8z1rRCQtkWAG4VfL+3cuT1pI
lcja8+RckMuaKuxvpUcM9O7dY2qhfKVCR55X4x9VhdeYPWw8zXTLpNB8l4wqETZG
8an+LgurZZlt3zLZWyOGdG+4aDEgnFhQdA83SwbcN3y6wYa+adVqEB6dzJKFlPtv
Thg7JXfvDlbtytObGv9SaxphGgGq5FxpOY/zwZH99ZJ0W5E3Q6bVfsCF6nxBMGcg
9U3AxUQWEfR5IMm/X/YCApfNfNFOfv5w1rqaQZLmQsbPG/qZrxHDWcLfFuaI9wW0
ce6kpIqCw5ervzbMeR0hKKxGa+2bERYA4bIlBV4+/w+QFWNWuO5Vlv4KHoFxPfgD
+tVtTdixuSFTpRi8Yt6qmC8uLPOOGnHf7+61K7v28eK8/gVA1aR7ssNeJjwzbWav
+RSaBaM5z8XpbPommIv3WV6KwMnzswQNBz0YQSrMwBCAVyAPEfKuFXJRINt8cCce
BGNwSYxCST+mF2NtF3d8VLqoHKAg3D551BA6BrrKmSHx0TV/Huz5TOAjB0Fqb5ca
e1qy1igGslN+kyZGO4qBYVhx6gYZ+phEfBOKSUBmhQvtJaEuxsQUICzx/zxiTB9Z
5DUPvMKM8ruVw/TvPoD6CceUHxykF1X3uDO0+/kAJOxKNUfHo6DRtOiK3a7awHos
9sH0b/YNRNvezwqgCl7+KMRvDvc+Kbio17Fq0kgBAMkr7xdHrvEKI1Lv4iemMaRH
BANpCX1WGpDkyxG9pqhLKj5BQHFkfX9tA2hqbAkg8SjdRsS3VO/AA2l//MurwIRM
5atJLkTA3IGT37rTRxmYKdbAS3GRh/qMsxfCiia/umdTftdjavcP6W2XYnJ5v9h+
MRrpd625ZLS/dfc0NWZvQnCb4HLz79x+pvVhjMWtHRh09kKHxxrGoIEepU9HQF76
8V7KBrFO3GyjJBrSgdKWMCQAqFKYEb7eWJshVYQvZKef+mQXmhxC5qy3jDgX5rZL
rz2ORHjBFr1sPF9gzjNYUOYTtUIoaPb/l4aJDjkxNKmVGq0l9Ev25in5ccjSbPdH
yBL8UaXCWCXPWRskWFM9BTuKpYM51fKntFluzrvJ1cmsMiiOSmf4cHZPdJLhB6qM
9BXOOKv8G4pWR/IeZP8NfEdPWH/fMRfHiKFLvuZGCvGkPVjgHo/6F4f3y5lcc8qO
vOv/gGW0uXJnsu2npnLj48mHCPBnMg5yH65coiHiXFZBm4eZ/4SYJNdG0gaeRL1S
88axbxtjHoYykIwJJmzACX7kfT2U2DdeMQLGt60K3F/v77OZUHer+F1VOtp9hVX7
MFs9UFBkm9AOBhaB0aLSWAWqmqxPYZaHyx6Nh4j2pzp5U1Mq+SyJtdcnooB4Gyxq
wvhgSWs/6ZNNyF/m5sXHYtFjvB6kzP0DGFxULzhstQ+FhqPuw7B1t6rQQFL8XWFM
2inkgNzjG1fdgYlyin8RNyDGiHGYBjeq4prVXbIEN91nYCNPuIyE1rJuLP1hI6oB
EakP1x9k7VrTGoY9Vtusgtqws+cvhpqtptT18owUWfAvHOYO5yWmHtovu/BStBOD
wFun7GeWPQbhJX+wHMU0DZ5AaPM+ippemMkFQHbVrg78bPnamwpG1lJNBs71fRiQ
e81GE6rGsSTD4kTEd9owsfJLS31WV35iB7kNGFn0nBgQLpIHjAlgGbTx+eOiMj2V
tFvTjOsmFEJ3M2I3i/e2sWOBpQ2zmnktgjZBhz8sC8aSqcuvExzyq9EYw8qYqUpH
kexNZRMKPRZSRe0ROTDWQuOzvZcn+LC+NWm1DQj11QJkPA0IDFEYsw1/DeOq2irY
cyjG+LusbiGMvI3QSrNhYhmrvGHTtsbbd9VOW/B1z/lyikdERwm2Vl9tNxmG0ALu
iGGMJLg/51TN9J5RHUsrT1J4+E8ZEYq5xvqLT/S6gpKKRVHz6pOyh48LVe+VicYB
4ecg0Vr0MzeYCZpbKAGCR8V7+Z3ssPgpPNuJ2QwjKXE6NSvtkhnApRFwJALN/79k
GYlKDSTchjlf0j0RjVurm/fPJ3G2loiP7081ULDpM5CcY6Xx1iXGuzB10vwlHKP5
gPZaQNd8r0OInExA2zHVG2F5ojmtnVbpGuvSm30mUAQQb3bD7CiRFu5mmCqOy0ar
M+0Mm86TjkpOID0ynsE6bP0ZXy+S5Go30OljemYc9YGxS93vz0w6c517V54tInk6
b8cCBRBMRBuzv88d7pVNZlmd6EoPYpDbNozFJDr06J+Q7jwkhwR8xQnDESWxCtqY
NCRk62qr9GsSqb33SWKSoQGUkzxaczANoj0gW3JRYkq6JFwXCffvKnLfUvtR2DPD
1TBNdvS3XeWtomnuAhuvX9ruhjjC30Alfyn2Erx1BzaBxbzsN6YX8zVrpNbqC94Q
OEpvEFlZwbF45tEI7VDdMHrRE6c7A0Gg2vc1BsjZDvjHdTrRTWyzp7Erpe1aCNgf
rFD3WHkVnteCmrJHeFVP8m5SSgxTxD2fHM5IsKMDTi+aafyV9tJ55ogwRmMVQMXY
nXbLCUK/ePzwSOJM8Itmd29DAZ7asymqcnHjrjj0SX59Qc5HT++7JrGpj8qBPH6y
gXhuZ9BOJVfGu+LCw9f8lRMGH2cg/1Ms2aQeDJVlapBARWntteC8dtnjlOKWqASj
IPznn4eUrAAWbeuUyC9QbNwXgqoDicjalmycJaH2r2NLLCuYowphGWgxgS1pc9KS
pMG+OzfXneDd+bkf3YGB9YoTZlGwTnmvqB6avzWMX+kYN8t+j9+KAUMFsW6wFymc
MLU/WoudRItne0OsAc+NkCr290pjwHzCYDCXiE2sEiLB0kj0EueG1KUOOWKRAU8c
obinki6JzYqcosqj1tnbOncTZtFtdgAACGJA/DXRfZ8ASPP+G0jHUIHoKkjxgY7b
U0OZw/vEGEQN31AF1jNR6QKFiv9vf0bLVoeRSevgV0Rj/iEFJlv2meQb3R0ScqUm
r61f2wQxu3hKwovH8TmHuRSnU05pIgxfAuSIEFH7qNl/6WhAUcYvXscBbnsBJacW
d4Y/xBPX4tmmPGq2SZSek8zZUI2CUzEGhWd9xB3YAL2LQgXoELDva0WegJAfXJvG
2o53e7azJt8sEwZ/rkPTOAFVCl5ns7dvfPoirFz7XWybULMonZhuUMMkwP1Dy1AO
2g37jepKedPf0byn9KMh/hE+2nYQ4775aPrp/9ES+RUCq00xSyiedTKtHTNXagZw
lalt3xKBKlMsJE4Ds1UjVfipoDpq1vngdEio2Tgvwvnd5rbu9CB+9Ex9OhIQ+AGJ
8fmy0jK3SOyGuEz5DXFm8nVYPzhtvHXRW9lSm0jSgXsqj5Z8RjjaDlG/VoGUkW3o
ioWSsLA+i/zYSyuRIJnJNjUhP29IdlIdQdLY8D9hj8S9/X0Kp69yNHu4hnOGwdJ4
lIvgRRynK6XzAH3eXDKsUsnnlyB3DcyVh8XQPB5OJot3YKYV1iwIUQ7eMBeVXpvO
6IMz8III60BgTftkLKsQnge8GVtynRUt0wagOlQpu0I4uMaE7VYNK7XjquUCK5lY
/IpDMvkXli/iH+EgB/Vh2zFfogn4YkpfYZCU72NnBbh0Z9B8OoFDuc9c7Krk8t/R
jfdNsRcqn8c1Q6mJZgfTJ8Gkl6Wnk6oxjm3jeN/n2mlDcZ5a9vdg4XPukeenyPgn
w+bdA78FnzJ41ihHiDP8sGpNR3dR9gStfSnw2i++PtXY2VslzrHGNJu/UMQ9560o
+EQsZFgiBmb33GJyJeiq/J45ochcbL6Mru2SSOGVC0r8Bc25zWe+c+64F1HhE/7B
OnIvzv8eGMFSjFJrkBfh/ool+MNEpaI6QRBW0I54tqWw0R8xLFPrMfdlHOUUQupQ
+ChmQQtwecP4Vb3dysPib2qSLrMJVJoILpLcYkXCxiJPpxlHfuXzNAfnoj+jKnck
4GqXTtDiEShHjGDCxdKkXNWvj5E2/gLZTRMDY1YFVMemcFGno2fUglEY2xYDuigC
7ckRN3aWnu8OjhUZx40+xaMe4ROcajVUVrYdK5aofMdflIgsEyWrJtaMX14JVDEi
R0hZdbZ/MykPqwfZ04HrINsqbUEbnsVoTCFq8auIns1T3GdBbcDKujAykOpNg6Pf
5ekpNuc4ixLtgg+9iwY6zGhUn1FGu5GvFvspbJe5OC+CaDAKvN28TfXjRlO6bgpz
INFlBSbeonQNQl9Sn10s+xDH9t3Hou9spW9UE74Cz+Ki8OKkaDBz+OmKQyDoqFzp
xWlWguf5flCpcrZvB7enfqAKLc2iu0hF1i3mGj/YdLiP9F9bnkjb1NzPkVA+yyEF
C8Wfucc+GqTQMQxifSrbDvvBt3FtrrzT4lb4IKdQEmCPGLuM+tQTsi+D3KI6ZBDP
l+mTnIngdgetd5cKGEUD4DoWPRx/ZWXfkCnkB7wnMxSd+jma5LrO6l8RQTUrpHZW
RGpZxY/KJd/GjctaYr5a5HWCAxdOe9Tm7djhkR0So3vfw3BUBqRAhKGPcKt+NNjL
xf0h6iIA2zQzTMTcPfWVPvW5QeqD1vwWNI6kGjXbfnsF8xfk6TV2n2lYblOS57YX
u0Jx1N/S8Jc8GMoEgV/iX7ddKzuDqJsCUrizwy8vKKQci69/Jt8w/4o01w2KEzpU
YWVBlZ1DZtQkvK1rmV7q+M+/6+WK/z7SNETQkFiHwsWXjnkTOXt7sCyVKAPfu9Is
865vfnvs5ceIUIjvglHmCSjRfoxotIqEF7HIMTE+j6kRpZEZYJO08Jw9FD5sVcvw
MgZV3WoIwikbhrLDx/L5Dt+lws7s3/GxNPHBH+R2MnWB3yNFSHAHKfDfiaP6VWii
YQ2+edGiDpl/C8672awUhbJLdcWmkgFivRQ3gOjehrHT9NXpsBNvVeshDA8frW7G
Yuv1toDZ1TNhKiy9b915e/Bs49OmAqLF0B3ypqoATsMQm2hoDZ0+VpvvhQ9b0nLw
QWldIubZptO26WyutTXeuT850Fm1+oDJfRpHf3d3weLAT11dNG4rMFFBeAgTTn4q
+WHjCxLaXx3QodkiSPCtQPUii6FjRLJjiD6CBO6ylWWbzS9IsSAAsOIyWPnUhDMg
rlAtOcUbRME9FjSOlweGM7zLpYuhdCAjIGUWYl8gvbfVuhDXHylWgqU8PbNGTaSg
HIkKAg0dKzN133N5ECyNY970Fzpy0VJ56mhi4E/iqCZFQ1jXlQEuOKLwBkn8ZCV7
w2t2Hk+NV7qjep+YI2qf7+bld5nwypxnj0saKJDji/7BSj7PxcJHbKg3k0x2YnPd
d262xvWZfdiQiV4RCDTbLErn2bRAHL9knT+dvondJj/57y6idHN4n69v2SAFAuMC
Rckxi8kpX6Z1gzwpR5+7y6YOt9UyVTHy9uYcW7VmymuW3Bnt3wDx53Ebak02Fta8
qP4qgcGD/TIE2mObLizxx6iFMDw9slfbdWzga+QHw7w1Y+FZR5ZHE0hUpl8wtJMh
OrYgeMhL66fh+lsxxXtm9ssO6DGlme3uCiitKq3RTITLCnZq3HP0V0fJHqEcmZno
4fRoCBpp1Jc4yBwV8HBTrDv0CTPimrJrFDlrbtkQSk0aDXSdUPQ+lv9Ou0c5WQhE
Yjv1FzBdP8qkccUehtYO2v4i3Wfmg3JpMlC3c9WTAv4Cp3jAEFP0fc9BptaIRzkw
E5FzvTDjLypHL9x3g1SbYmLUe9Cu15uhDDDon88K/IBRq/d/dCIzMuEcFmn8hBga
N7sE9pfqLv5VNmrZERqhfE8qNbj6VT0P6d5G5wb/dCleT7CzxGm2h4pPL8Ei8ZKs
+34PDdrzYbxan62mkWwSs13S4qD+Yz9jleoGaPll+dpZRpx8g+1ehQV8v2qni448
y8HTGkGsOBg5Xh9TA5C44Urqgan2nsRbdaV072Rt3RrnJQ8zUJecOKgQzhv3qWax
Nb2YCV9OEBKQMo6MLDjt6bjto/3kKCySNwrBxtp2SUZ7Orw71dU2gHgw0pDgNTNN
uWH4rzPFY9uA0N7Hti4MtmM94bcKYA06t3ohUlhO80mbRS5MIVPsgNdjQRpxgn0U
FQeJO31UebI+G4CPv2DeZoB02sWFIGFpn5XykhYYWOsp7q/KuV/QmSldYfRmzIgC
K6L1vKOqar69GWZ+PgGEzelt/VnCcHEmgYZMgf2/ialz0zHxdsGxaZPawqETNgbI
obKxRHY7KcKDnns6CBo/U1JGeFR2sjPfvPQ6ujuEsdX2SUA8fw0XabYhrcvMlyF2
RPAOcAXe9QARnvGufpeyAEL9794hxyQY9pS6S85vXSVN8SfIB/PCVqM1jgqwv8VU
W4g5a8ocVhisp7AoTVhczEIQExwHV9FdFF+fmc9PF+/Z4YUMZNsOvSKYNDa+5BjU
F570NXgjp2FBH7/5RY6BCmO/UmRQ04zONA3kSGfjIAWzhpUunIiHBmdTYuIRrTur
ZoSWoRDUudyuS7puVA9BiC86HIAC+Y+m+BQHpP1fJNKeKM53jc9Wj7lOf5JsDrer
7ZFINs4/ep0iZ2PAMtbg158tetnk57NyGBCR2u54g0L6znma93ZmOzHezklRlfIJ
HZaZNN3XASwmBCvXY5qzGe/u7uZvkusRhrDrp1Q5IqBbG+XT18KienOpf+mxK+7E
4qPHI7hIlNPX6Z7WDcmURtaz3oSBoG0W8amYNNL7nxWPSSqEAmz+wQy4aS87ZISq
yFgkBO9/A2aKYqEx9byCxpEhKjY0zmjho6p2pNIeSP8C/F8LbrI1shqqMA12PAk0
eWNutBSMNgQcp9zMnj7N/Yco6NRvZOETqOK2SJY55ByFBGZAkmeeeNDsk9cZGsGk
cycRaXGbBmB07gkhXZ2HoKd4b0DOxLMh9UcRzhtc4uSxyb80lcdWcmYIFzkBjxIL
i3HwnJl+CBhOhg512fiUXIfeHbDoGUzxVuEbKG1cYohXJO/rdifMi90oudPjzTje
J9h/V4y9/JBmRdfTVUbuGq5ZTncE4xLrD06RjdhTfzfKcQDRsr9GTA25CmrGeTn5
OSQYzUoB+CCGBiqyO4pxQjTjz1j5hRGaf4b5TvxH2BuhlNh/yIJSDrio9q9hMbCT
vtYu4Brc54Hs18BWga3nGa+7SMLozgCUjB5dWsPJkrwQl2XwN2vp9/fBGtKI72cY
KZS3LZaE9cU3GifcTmIEpZUgUfl4FzeR7d/LGjjmgC2GSqjbfLwxl3f1Gu0257CU
nIvRkImD4IjTOC/tIiZgeYryUysYvAaQ0uH4ymOsIe+FkeE3hhTYDzpJVfROH68e
aCj5TldYpu8UMXdMM69B7Rm1KRhLf+JxsZDjJTRbgkfAcEWARTRgzOMLFcSe1/gp
iJ3SaK7phvDGFzqcn2dH76cQhNbTTory6HqVzws/xq4SURuZSC8ryHRbR2f++Usb
dtdN4+SKrtTVh9MsDeVGUN++Vug/2pNnuVdofRKOfMrdulBUv8zItzdLhcB3hPVe
Apc5OrEyevn/kmIO43LR0J7uo5LPeGwfa+87bVeg/u9EJ9LdSg7pZt9DvI7v4yzt
vh0YSyITwnbapv44lWrVXU27nFJ5YhXyReRyY2Yt9EYcwN2oJcLYSgaD0Qaiw6ir
FUr+VG4h5xECJePoFHP+MQHlqztuBF0jKMXYFAXwASFRibzF0RUyALW/FdS2dfXk
YBv1QvXjH1nceNvsS3zsSnV5MlO5F/p1ffJQq2sj+/6JjMYONIrApS/HOMAr5aP9
RNdIUCefJnS9lg97icaGap/UGg/UNd5WTaDEAw417tlaKcMWh7EWcGAzfAWC3I4a
JMaWvI/fGa8xuVymNrYzsKJ8svXgYD6STBYUzoZkoFQfI0pMJDPgqsVKtyE1fD5m
ZEbmvQf11N6m3KiWt43tMcf5GGzuLpROgadzJ+xVBBtoNvBFlcEi1EfyCB4bpC2o
w/bItFcphMMv8IihxBhabHYyAYqxRIRTpBaqTatOkP/esPEpVTFTQd3atmDDfoPl
EqvpTS4zsM70rsWKk8xivfKu+4jqRIV0CngpRu0+LbEIy+aFq9WCLOgkPVp5rSUV
dIVn0EzoMypdhHvrEU6qbrxwez1ZL8FyiB54WypFSUhwHLWwD4CL6Oz4foNryVo5
DPLdtzCroLVG/56pBuCVtW2LbiI12Kdv2e4AJ7yZZ40bY0CZm4GvijAeu4qdeRLx
tpPQeaYYhTPhbVYe4gqUpg7rBtw0cTFxPCZweW2s4a0jUOEO/GkF6xVlmfPFdiWv
ETv97OwnKHnSCRN+eMimQDPjkqYiJXKsjqJ4OzqKVJaddAhlardAYTLdV5Bz5X4W
hz69IDUjD3JtI+Lzq1gJ0pxIOFoXw4wgZWNt4dYevvGHlJdyhivuuWaUjOC4Elal
/N8GiGHxV2CcArBvJzg5vRkMz63jWYHLGzfMbjC3syPu/J/YyFzBSRjEOTrgbml4
Nsz06f7uJMdgJ7SYHKqPyQGwF8zTKNr265jtMamWslwmr+M3E2xGY43Il/9pTFAI
6QuQiRQKTyBVjaTia9ruqxedmy+2CAO+NMjZNKfI6cqS4BiurXH1MTZGSE3t+rs6
wJl+t8rt9sq4gnFk3OWyd8za+j1M3B/o1+c6GyFkr4JEDZMFuV2l8r6zab9HUatW
/wiXcKdPYh8/yacE/q8+It+iTn1vwuvoui7fAWRxYV7yErXcjO6N3xuTQEeTsLvw
WA+HXaYrirJXQIftWyTbHMy5T5rEZY/sV44I9WmMjN//W2nx/1u5GBczoFUjAnaK
WfCKv2zKDAvngAZwCr0o5anuZqHgEbi8copuK5J7trX/P+w6s7hDmj3nhzGFPcXX
uZNymgd7ZyxThoKstvBwN74qVvWrGlZ1eoLVonzKuHVhAS7hbdrMC9TPS3mnkel/
H0NL1Ija8z9dR7vUyoJH+3iyWDfg5fPzpaW0H1BDw8cifdld+i3zL0YNzrczkoSU
Tqbvd9h1bqUug/ZLXV7y3EgseKIveN2gr4Govg26ai9c8KXG02w3+l+0GEutCaJl
db6HXg7bLFc0a4jXK3L19zisFN1QYPM2CV9AaLVDa/72Im15CGQJdqWGZqhiJ6JG
6jVQ11teeGdyWltdTJSaR9bZdDlsCbUjiPlAhrj1n/Cf5guzGIcdxQiJi35N5F8b
SylPL7+dNMpTfFRJ2DNaqBUsT34EyPJuixHqmBIdmBioPTUQ7eInzME1Zc2p4csm
9b1dUMPjd3VwQLgj2xH/cctbnN0HCKnedn+umNKKNFyDCHNaLxVCCorUlz1z6PxY
ReUKBHaVAmI014ALgUHEXJA+tO15Sse1JrwoUjIQ+bwP+gZBF/iHvYw/RmaZSuYK
/yIISEdQmGB0yZ8jshuv1S0BVNsMpWeN7ui+hbT7NFKKYxvyGeKFkdtru2b2ol4l
IkB3jgFav7VT7l2wglKxkgCK3AnGvvQYIoCsb6KfRcq78spRtB4LwE+JIHR/I6Ux
36WbBaLUk9o+hJ2AGVa0dXdDHXOg5mjicp2Un35IqSlPczc/zZFjJovB+edZLaGe
Duzd3s0z6TTHzwF5YMAuhzGmXELeph63XZ3kMO9VW4QsQClTqEZSYegVAmSRxQ6i
tmfLD9KyAue6mfbiSJ4OzdoIK/YtoIqU3XccNzWkQDvjN+K9N6bXSEl4fTrD6RBH
v4BmXRnHO0BLnPhPe2SrBdme86BzcmvW/smlWCOCILAVAm4uehxEx+9KxQrapKJr
hZCwoZiMFTaCEqZp1Gt5gqrWWxBmv00lh1LTMWTa3+lwhlzi3SN+i85zHoiA18ry
TCTXRRBVInVUsXu2vXUmH+88z1BeAlgCGF5AfNdrIMeZWBq0Hredyf8219j33aBX
d4tBDWAPtOqRaRKf9Kr8jcf3qGsua8TJvpkk9UoaiGN1jqbL5Y2bdlATK9RBSqFd
wUS3CHbLKDn172oM93VQXB9oWORBoiLJ53Bv8o6v8tpV9ORMpGuzqHUfXB2fHIRM
4lfYUZc1MKriYVTExzaheUeuhrkcF6OENLqjylcPkzEBbtui92S8V7vHzBqgG7UX
aKOGvTEtvIbhGGi5uXknviE87ZDjy1Hxp087A+QjhIV/nl7Xu7xUDdqmsjuzQh7Q
CGVX39Lx+qxeOij5UoAYzweGOj9I8XOMy3GxDCXZapoFJ/dI7FcYrE0IoetDUcpO
duSS3tpV5mK3aTJgAqfzGh83zNRROnQ3gwolIveEcyw9pgdVaLdzpby5KqMxCrua
ouSgEH+SLbi+S+OxtounhOVcoC+/F9uEnmSobaVH/n/z9VPkQPxtDudWIsKyaWFZ
0fsglnTqYeH7Hp8OZwgRZZIAuUtFSh71edws6tzTwwKltPi3ArbnX4kkgLWALzrQ
3w3YncdJtnPUrLPMAH6aevG5bRwzNAEuERANJR6bLFt6VIF0AKAy/xsDTBKJ2G3z
QPbVh8C5GEXV5sWhi2cu0frW/lBjAq8cx4zihZiiNiDhGvY7XAQa8oLaV+p81eM1
tykNX2fH7HEbb3GfmdlM5T1c21/950gjgT+Ugar0eYOazjTLKMfZu16StNtXJUKK
hQgIIpe4ThSntAohKAoB9tyi3l3Nc4IjrhpAZE3khVKoZ8p7SZPxiezjdQZKsFiV
0/06mKil1VpxT/MRkAV5sLo2UaETn5Tu98SGst0KdGM92eF72DuCy/qndhoJQLB2
wSV+zbzSGU9NOyU5WlVaT+luRCrbYUedQ6NgewcSDPuYq+4x5oPniybvGwJnAVc7
E9jad4e/HN+EU3CwrG29OjaNCIXuElmgKs6oFyp3B/oKvOuw8V7uCVpyv+XsiJKb
CevMHzHZeyhvpFCnChzMnKn6n2OUk0Ky/MOfw7Uq/uDvV8YI9VMXYP3dKkX8cld8
FryiaitshWzoWfEenY18cweru5Aq8KFHwLERWiH2I8vhaY5fpFOmgMQ4omllyj4q
fIN/a8QzOnILdwu3Ee/2GZ1ZPjLS1iqfjGYJLoLd8c78K6B/cbUYZcksx35TEdG7
74ML3wVi1DO4J/MK56YLLLhoVPnXkLS+AetwL8Kub3FoyG0bx8i0DqoSGpczO+Jf
4c4Vs+jHarOJX+AG085ujnlJiVib/XsrAFTylGE+xfK9C1LzB9u7/eCKHeY2Fc91
L2J0GJdC3KuOuXYfcl1qnfqgDeKrjQ5GjUQvwxE0oG/ryrW6/EFahhml3KTBUlZB
t8LCJYX49rlQ+EZWAB7FyOKjhfoQSJ6kNLT9CVhBLddmdF5/ZhmlbMOC+KbW75C4
ksECvfjTNxDeuIWT9TtzG9stnQM0w/5Njv94BXyYYhneoDRtWc/XVvc1guhQn2Jh
9UNFb8pqkWXhMs/foLLPxgzPwOTaWletV6wij4qIjm/lE7o0i9t7bSjvIgLKgrmu
U4e7yCfWzZhYqbT7p+XJNFRLbxG1p0t9ftxy85YbhTqowPcGMRUcgMA2lUcnM2PS
Z50eII+NOYiq4XUkJfPgxbCBiV/2pmlghy5Zcn7F9TcxbwcPpnH0bbSkTErcR1DT
uM+DYDmstA+DbVUAaDFIiAvOwkTzeKLkkpFD0O/+hRCRwBnkWWBMYUzAbqKvBQAT
yIKPtyK4XJeuio1ZiWq1ujtW81Ux+vpN567yek4w5XrCVBtLg5Kn1+Sil4jUForm
lfuPwQRkuXjtAWQn88irntfx9bgQNRNupkZRM5lLpXzlgeK1xp3yGdtM/cQTT9lw
7wSSQ44h0ZoKjMroWGlVTPWENylPJlMQfGp05L5UBNbHyNRJbBBVVpomflbYMSUf
rEcAWoTzQnrvNIZe79GrrETdZ3bfStdlTyVEGHfEJFicIDiYPp0zifGg9k3sIoKx
CfWUCDRkmeOgyJ6wCTsbK1TtdGk26ochZEzQGHWDZGVvxDfnyiDZFkSkEfZhhprN
xxkUV4vuWr8h2VCJqxyIm/RqrJI2nX1Eq7B0yT1yl8UbYcZkx5kOWevkb7eZhIvx
yVAMB1Md+QEam73N/BwPQzegxu/WTzE8ZEAsQATCeNJsmJw3aqmwI57Yk1tDV43f
kbjBoU+q5Bl8fFBHHRG1QG4Nq3EkeqKxDWD5xIk+F9+AenoYrQ1/r0eXx2OgsHpH
JstlUXczqNj4bnj2OH985CTL64WIMEWUL915G/ed5W65ZvNw/AGN9tlkHa6Ji2iK
CeEs5AxF8+Tt4YeJqyQO6mL0SmP8y2OSsUR4u8+COXjAzWZvbuMAEcTXtRyQtzob
MdLQA1dITqn3l7Q5Y3sKgpe+AYD+pDu4kUy0JBmyB2cWbcB/2ujoxIqrsPSei8zt
QAe4yUuNTMlLTQehA3d/hqL7+FmM3hoHehu/H+im+1UTocfl2+f9xFFSZJoVmrUX
55Ks4AUOsymh30d8od+Z9ps8sa9rXKsXX4bOosQr+3J1MHwB9//OnC9FNB3cep7H
BXEsf0YJ7gRyTnzlRcIrZmLjRWy5D2RgNbgnkGjVtmKtrm6ItfbWuSSQv72SMKTH
rKKniuzWQDoEdGKe9EoLEBdablhtt5RYBDfXV8AL5K8zNXDlmGDb8Axv4jWYYkFV
U96g5LmXtRJMUd4C7kRS8JDE535i0PkEsJd4u0bAlahTfCxtph/pL/JaH0Vgpsv/
ud+HtaBhKPYtYyC5lAXZaqHeXWsgzLSskYKlz/SR/zz+AYXQdL9GqM81udgFW0n+
j0z3Xb16GKzUPNntwLfBH/s7WxKoR+ZXclDpi4vre9eUVn9TXMlUkf0WnU7m3Mgi
dXQcLfTQEwJu6BO9hzsIfckC0ylsp+cQXF7QzFrAQGieOYWcq+JDjmyenGDkVyst
VvahK4HKkSdJQdupwcUnasXwoI3tC1rDazkrcWJytGFNwwaYWJLGTbaVT9MBeou4
RCgCDwEx+hmT32A8DxAyWhfdBSug4z9RhNZfyEVsguiQJG3yi2QdpXd1cmfgMwF9
bhZvzn8zIm1Auf80ER10/P2lKY9kO2gXff7LBm4UdcLMr05lWVp92UtjUtOID5uj
U/qmgyxNxNQfez7TyiTCvY/SoWEiBJ0mIl0PQ9GkYpGxF6oVhUjxQexEu5NcBXjd
sKVHS43Mtc9lLxb4rLfiuzTADM7Za2N2agmLf+k0F3KaXOQcLfvk89/ftGEBkhzM
/EZgNyGwAMcjdyXkCCQvp1INqROQzeq9RjXNvuKBG69P+v5o6HvCVdc/RNgjWGTW
IKuhIGn2fFfjPgLf9k2eBVnLVCyVaqyIglKzL7PHP4x7IQyp76j9elZZs/MB0WCZ
EXY/9CvyLvGjiLuN3h2HNHZ+Ab8E8livsqkitltdKUBpKZBwApP/ggyMEIfZcIu1
7kOPYCkoVcVfj/roRbvU9PeYjVUzZ+T6ydvSYHWEZ1AcK1AnH2dlnyOHX8BrPd8u
yNwyFJ9BcnkeeAR4SrBdBTlvSWoZmuR7Y+0vI/W4Qgmyj0v8wEpFzFk2f4a8qOAj
4W4Sz+9uiuie/cl5kZ6ok6YQARMT/cIIfnNPiGvsmdi2a/GehV39Z9T3kxqkcSct
STP9QLmV6DlUQfioxj8GuIOnaDAKzw3cTquFj95sysRuzK7NI09Z3PvMrxZi8VJH
VAm4kOjkzyyrTBdSQuqpRmWQmXScaeLKeDOzlbzSC0N0KEPi0HVrQC/wG92Jrcf2
X/CsUjTk8btpM8nCnKi6w2ZN0ZUtTo7HJzY3S7GmReQA67AfIfVeqODIob3j17al
Q7SeTXlSk0IJqZvnEv50A8juZRq+XxgJkAUGPXRJKHM59ManSDqCGovwaVdtw5Ds
tvsCKjS2yKBxwnYwJr/Wtf0BtaS3X++62J+QFWECVZMkB7AFC1A2UgXxq/0b1hfu
m8L/c8t/+n1ipDPBwiVp7hJievB01KtpE0JUaltME6UmnMcmJ6sWtw5Z95jz+u0N
sxYrRkPCBxDK0GgOKSDDu0JlMHEWvc2O+eSJk5Ik7Yytlb+3bvu6+ZuYhC/KBKtU
F4rbMhQCGygbRiK+gA6I0EQqPEQXGZyp1K3drA7OG3g9SynF0WrQgwboWr9ay09D
HxhufHUzrJ4QE4lpt6x9o7NPqLSULQ6/k+P5MWRkycBCqev4EgufhSoyqrG+C3QI
xMA0FAcR1oa9wHqyPSENfRw33AG7NAWt2H7mH78wFB5ihHf/H3QQ7N08PBW2Fwax
/qFHKJZ6edhUhZSvGewnBB1GFpF4fHq2nqa9fKdSnl5B26rvjQ1aP51pdTEBrpVp
JiVJ+MwzbGT4/QijCF8clZ8+Ai8p9HsYEtBgHQqVQ9rLjfPN4xIGLXijkG75Qibx
gc2c46bW6rlODbC2u9e1440tGvguBT/8iaPLmQnxMdCX/GZTyr71g1Ak1qITRgdy
9RLawPuR3iS7c/Y7u4o3wCpv5STUdXkBwSASw14Fkd4ISnupB5KQOcEMo77r9zE6
QWLBawJXAXc/DBchNPKgP+snTmaCieXlmnZAlFCYIj0EFBN5GTtbiOZ/8MnLVGTA
Wm93LRSTyFZn3ETZf1XXUZ/GJVSn0clJxqMDxYuOE44Lum16h47xsuN1YpF1/vY1
zgZw3iFRx3VrjiHD5MMYm0p9D+f3xihS2Lc/O+t0ZFrIj9q1t+MVf1POe/QrTHA2
L+mfjFBnAJaaxt96xnkaCxwnaetdl1jPeQWfB39TxE6hs6d/I2PJ1HJMyzw2njI/
g9XfyK3su9bcf5uBdIolKLUQgPU04s2gro3m+PwqgmJRid+PbGwRNBMR7dWxK7FJ
LTWFnGw0QEPse02EzRAFwFl6EVhQgeX8tbcRYB1UFONACQBKUk5TLQxGtTx9XFqm
FU6E37VqyiOjPbPqeT2SVyXO4sF5vENE5Q9l84ZNOwpTt+4ge65gqAvgxQ33ll/Y
Hp6eny/kS8EefuueHs0/CFPVZsOGtFaJNxJkor3ZFYURIFiSAoDqMRD7mNklhvJN
qMrq6U15WBcLjghVlMRWeFSeK1F62Ye1kTsWQDGk3Z6+NHj0nBmTjLrdESePoYaA
eUb6DvdkC/GIc5V1LjLABZIPmekgMrEwwlMKRwvkI3kt2qf8Km/chn5rrVlfNFFG
VRNpqY5nnaQ45L+/ICxg8fJpcRITDYjliGjUwety4WZmfrESU4nkbfj08opaNBWs
x9sr9J7wbrVn/MTN1rUx7j9PwdYlq2fjWCDJxT7DjAW2tOkIWhUEphUD4cqod0gd
FJMfyWT1hwVlT8dv9+Go/5lqE/GPfjXYvola9N6BVr5wCkKjvnUnqgQSciTSU3KB
5R5a8aC/WUDPBguZtEx81OuooCJibWv8FfKBOcObwFWroRxeeS4/CdRhFHnLC9ab
+QVXv2ITcWi3fHzM8hHWTq9n5Yq1CWszzQ42pkb5ZSpIku9SinBbe/87ZgD+wk/i
SyvG+1wVVRS4uIhcYd7hhMYl6AmHtrIZXGxgxJhyqdKYNBoEXMQuy7GqgDkGo0QF
4N9bOp31hPvg+SEYV/VEvfvXQ4QcD4FsBnhhiiGuslYA4IlrdCW0AL3RDznxlQYt
fNFi4pDXPgUZ9MqDLiO2oeVRvrz4YMJOjt6mqER3mdoClvPCEV7TBF2i3Qfocq0A
2vua8RqWJNfjTAay9GeGGq6A+0ZwDg+4a9ANVE0ZZsu7Aa7Brqh1YEZNUbTB4niA
DjD27TGcksLYHJQPio08xiDDqAfaeojofRzd/e1BwOKQ0zjjzxvmaiaFGrSIIlZ6
hT7YpWB3iKm6UPl+2SL9c8OLywPtui7V2ySZDKBdXoIEVuIDu85nQPWWnMS5Ox11
mY+7NVWq9iQTxMCYHvPeqzPY1zbsZ+0St6yNzUyrxrfV3Af9Zi5l2LTvP7EKQa04
LFXdzeuc4MmLP6ZkNurhUjIcRKSzQP1CTHblDLcGiVVI6np0Bcuustypl4Naot27
R9obtMOOE9TqF2/3NvZLQ/90q15ES6EwcjG+LZH08Q0WNC5usnpbJvl3KqWOzTwH
M8R2k4nASqmfBZj5vcj2AUiMvbSe+Ap93QMeoSIBmSDGTvPiDxud6WHAbxj6861M
vWKQG5X8wQgjnNA0s5NGU3cWKfur+QsCEbqYwBHofZapiyO8Mu+GMrN1lNVLpiS1
nFOnWrwWKqenlKe8vEloB2UazgIvR6ETbZI0D/DVud89DHkVb0DeWpeAl8uwfy9b
I9Uf0IPEK9t/5gmGPUXpEfPPOQeTVnmSbK90ff/5ttTVy8oFiB8NGfQaf+z9Bllr
KXmpJPhYb5hzZR5OgwPpCTcPdr16ms4v11+jy09TVW6hTbz/1itXKijcQ1NcPR8q
WdlS7bwWzrjFHAfCNxzQF95+xEJh8RcUpCynpStzc9sgw9SxyBEyRjL6+LraPa7A
lJ7R0nKdRPgyy5gbpGQVRM+Z7b2XUQtbNCahgCOM5iw8JZ3UGMMEwaZVmd/x9USH
0eWZWVkKYku39eeAGcSz+DOcRrwvGT78xCEvGW7/SP7U9qIJ1+bnK25S+WO1ORuG
aMZ584bml2e1/C3ylHybiuCzsifJvHwEGa6tARi3th7lfFgv/8+XpYMszxVaLO7D
FHZEZoDAKdJOX/XSSVgNujjWLsb8jp1yYWaN35VOlYb2w/00pBwca6KZ/FFU2neG
In0Jth2mW//3heKfXD+Uyc57A+CMJYiPio+tvflGWFInKfN3kHLCztJuqkM9UVJ2
JkYa6wWSRsu+igjro0unbI9dGcrlXFiszuZ0Biq1OiFCTvQOgY7ylH7Rn452JXU6
P0VAancKv46zvmo7/zrOBh62OU+Pe/rqPXrzMyjxCevzmRVZMC9nKaXWeu6URU25
URGQtxHDDlo1+1Br+0EGpv99XciWFVEePcisN1xfTPpgMAC6ObwVDTIjjPdC8ipi
kZt4T9IKG/kgBZFuMCojoKcIPsNzMa+oyLHK1OiPSmQa7qvZZkRbvxG0JWCoHBHm
arkVBZ6WnEA3EDCl/FYpnI94HbZFhMHoyZsbBxlCa2XLqwwQpVUK3ABHqmDd78dt
YpP53ThihDulPPxRJYbBbca5R+wLZMUl7JRb/h9DqIXeQ2EXj9s8ti1iNA6mvcJD
eQjO4bL0NVYLtJc7QY5dTYedCyRlajJ88OqxnS/qAp8Ik9kn/4jxQOLobkJlLZpR
0DHeZiQAB3PokrnNfzOcb2rTEPVx9cBc3NSoT2Mt1a8Wk0JFqwPZkY1glH6BRtm5
7Oj/3RPoZVvc+5BDwi/gFl7Yyx4Wrm0sQDykWW/ccdgAdgjUrHMlDupmWPfM7ipS
zmkWtAH1V2/Y57Ap0XeKCv2aMdJegCPG3L7J+8Md1olBwgi1VdxnSbF2jcKJE5IT
DEexuU7aH5Wkto+eQlL/c+WevIE9HYUvUD//izvar+7jfF4INONRNe2dbAU97WQ8
qDldyODCeCmCcy1oZQ841no8YLSTbvck37oysQwbbGIYsEQmytyajgWp7isUE/sv
mvSaUYSwuUnmGQi1ZDjme+hMiQo/L8NJ2YpItjMSfMmiXmZSXUnBRUMVR45NnzB/
XIrV7CoX3xxVbW3xbME7cyqm4+FBqeUTVdw/xCTr0t7eM9Yp4HpahRPBrZpWAgr4
8eGDQSENK12o1ZAaqysFWksX9WSoqEny91PTgMiI3sU9Q/Ev50t1/D7bWd0FPWcQ
7gL99YKKwjvb5WQV2a3gPtSOTeQB7YhyH/0z9qbxxNEl7wSab/Rc3GKmtsbWZoqV
cyFBa3M0erhyFwnVlBbhDLb9wAzcKFHNadIxWD93FVSl1E8u52rcDStz485LwUbM
vDe3ob5nuf9kRzuOvnV0vQ1v5j1m1sykUWt1pRXjWSQ5tyXKB7ltLzDvaMWIeeAz
69KR3vyHPGCT/QePSD2ZR14OqQ2bvUEyaMSHwVrW5eg08i8kcPWTFbKnKgxb6gUK
5LuEXio9oMzGylM7Xo7PHAeLIkx/ldMJcbicgJ54rJNaD02LBiRBGBy/NgjSzSpa
CIw3vxx5n5BvhWRRo1FTHcMcxYlRzxwtoaWbtDefkUrMqs4hmN1QomDkROco1+u2
qgYZFFjFa6DfYRJvh+yzQrKlsYggIgA510g6c6C/fnr1esTkwxdWRK0cIZlZd7aR
pPvi7fLFSA0NA3CA1fAlWKAEq6ZZWq7/bZ88OxwfGjvT95OzlXpMa/T3puCXnTUN
qr93cUwLpxzS9f2ybtZBE3TGbF61tW1Ryzioaw0dKukPuHzK60fwbanuiFcfTqdx
oMV+AeZlk+eYWTGvQ6VWge354XMoNxSO9HLUapNhA/95zQxerp1vFbl+LZmG6q6q
2RRn4eK5a+MNpTCIqGVlsSolvsTUVWOsbKgpEfwTY5vsgKMTmRPh9XU94xAvDyZo
OZ9TStIly62EDH/G4GM6NO94CeFfVkX5k4S3kHXIrhPCYGSyl51geiUkeRCFBLXx
lBRyRzRu71ZLcqdlzhAsb3grb6im3RlihowILQGLjruuGas0QGQUUF8FnGBeKJbi
ztNbkwPpCYNuyuNbLwoR9UrRZoMksa/CMrvFGt9ScubYNAoeruRuhmtEkx6Pg9wX
QmXHFvgULwsFKNiE5EdpKJJg+4pUPIRxb5MgKTLjTq5G+Yd71G+53BvEKhx6iAiB
bet96OcvpkP9z3lYw3iTK70hVYHgmoW79mrGumzdv1pdqMUUrqVBjKO1MXyHvBQ6
OAhc2iMc6J4IV1LulA1I7Dj/gpwnE2l3q1au1GYGHO/tqGQoHuiBUwSksDgSpTM/
IQYpcu0dQYPXiXbH4D/C0QMSe6OORHYummwG2MPrfpnj3ImRgy7NH4zvIx3wZzbn
xwz4z6gBmfnh9FQFOYJaKcRmOruxUWy71Lvvq1OEU6L4z46VJV9nOoAAMouownDA
8VID2+qR3zAJywt3o1QYAOh0pWAPdzkp+pAnP7CJQsKpjwAWpWV3XlfMR/W0+BRA
maTyNimboF1tmE1dKSYxGYrTbAmVg+tVK4fIybVVTpr0GNoQXIUeTj5Pp3yXRTO0
cfom8GcA3njZwSuikRrVGqJmnhGE5pGEwRMLJShvhXzMKxQgRKBnMu8XxByd+cR7
Izf52/NBktccqWPbI9kalitFIiG89lT1kMsEza5EQqNhXGEkmTPSmCxUew/aMAwJ
20BVQovDGuIDhRMaqrrMdDk6XL2HJwJJ5PPq2slqe8T7JsP/oZu56n67pRXB8RqP
ErlNO62hXn30ItrSzXXKJ12kxpPhrJ3yM8UeKt7//wcXn8pnJDIGEljYzSXbNxRu
1PCtu+5jbG2a3NEcStZcJsDyPKGsHCTQhVGmJvOM/ZbKl4joOL29sbswmhXKbMlU
LkovW/UPNHevETJLp7WOOMdJbryXorKujoyiueKEowD8vAs5ejew8IlxF24WXbGb
BuNnsnVt1QjupPvYYolp5ajzD3nF8qeRxBo5UsWtRoIy/3qEiNVyaRmwV5j6Shkv
A3n38JYTJc+kfy4C6OjnBoveNU32JGTHsS49ShCznjaTXwonkCpmDfbWnnsqqlr0
4/RR920Z6OmIgaZuXbn83j0iIAbMmdXeGztbL79Y/uJYI7sTVzOodMB6KWwTq4B1
Vk2I/Hj0H3TaRoO4kIJbGDMIjY/haVDK6L4DMZdMh2g+dO+nXarO49oPB93+MaDx
nvh7IUwlGQem8OkdWPMU4GYHHLVqJdI0tdv3kUqQl6watc6MmZJI/snaGqn0hsxe
Phm4EAN4ECyL1SG7SnzIzU4ciBiucV61Wk5PhXxNkMzP7XLsP0qnmbSh2xVm94AM
CimYyicm0+OAjHbtYE5HlKxiZmXABfW+5sNigKeCMFncbv1RXs2du5cSboMXP2w+
jGTndDWUYfip52CzlbY79LSLtDGYQ/pTyt3n+EiZwfHSrWsnHxXj2Y5jRVJ74yDW
/Vn+aqgl85MOrn/2b/XHC4V4qBSvo/mLt8+J1o3izBRcuAVRp/v0Av807BtlnZyf
2c61nTPNaL140JflunA3Tsc+7n4rPweips9S+GWlXpettDyp3olmefVW8HhgmGo3
hJixTpTPGrbyCVIRP4u0R+QMUIjeJHBh5oyTiju8eM3qXBoblAcsxpw8L7KPa05Q
U0HLTDoz8QBpYuTy7GSS+FpuAfisjeZQCWYpn8dF6atKVeh3OqfoIZaFBfazB2OT
/0u34JBfjgQX4M4sC6vPZ/7rZzKvSYzwTdOuvjIl5nNhKITKaFiq9TEjsKIC+zxz
v2XGLpmOAsdb25CRd7l5psfITPTGr8CEvqE3bcqBYyl4JTqoeiUiRraiR8JsYrwB
RFAVAYH0fFbeYZ5OtbT6TU2av7Z+C+GofusQBCdRI3dgpeajrpHvflWCtgLGei4X
2NpWKvbhu4+Kknsdpor37wcKnbkRW/bvPBC5ofMaw+caWpSTvMxTfLBrY7FptrmT
7ghsqgRdCHxKST+KYc8kLyGys8y1DKT8fqKLo7JJ4VeACKXcDLtNxqKlj7Mv33xl
r8QoiR+o2E6/xs3bjmy6wsWpUKwrTGNm+eUNJdjy6L3Z5LKaw0QxEcTPu7tAfXb7
kAv47ACL69AgXZ0CjQQWESOXodfmVpNn2QRNqNRE1g+6XLDxp6a3UPrreRx3qQTE
autZ8rk7FU1n22ks2TY9nT1732TgUxqRKaTfyRyMNsc7FkzZHH3cIaIhCj9ClRJD
siOA3wyxB7HVB9g/7zEk5vSFhPpXBiGtf7fIL8kco/vtMl+z+en07X8TmDimQddo
MA1Z/TE3GALTTutchjn5S7tgmAe5tNy+yb8G/XL2IofHUsSqbKzoK1jn9wwZXBiP
M9xlOAXTvj0/c6Q8mx7jxVe/ycuExan7BvVWREsf/9w0Fc1+cd0/8eAK8hdOaN/F
k/dZ+ktIJ4PkV7/dbvk/+2UD7LgZCVVq+XsytAwaCHlwpqyUnDEdQA8MojyCt1Kv
Ofoen12mJnviAvrl2UDu8ovRx0QJc38RW2J4O+283VJX2ZjaldQPrqpqpKMcjY9C
KSMS5T75JoPPlkL5kv8sl/8NEMgFpCM8ujRfKEbRYLdPFrtTfombwKum5k0Qmwuk
0l/FiqsuGwX/5yeBhcCcTY6sBMp+4x3eNcXBBGjIjkXB3yDE6InrH1CatV5Zy+yS
fjUyMPrTN6oKenWFZvzt583OGHFFmSUYsk9skOnZMIfDbj/81KhAE6NFAPTIn4CC
tY1SDhtIex5++e73Dd+M5OfPwtt7JhZ0pXBlOCnkZooxAqtnruWs9Sxx2v/X9d5b
LuNIaVHF5VGj64RFGp+WwmH73mZAABGAbqK0gbLTnPH6KBvenjXxLLHkYwL7Wi/j
g3iaGW9VmZYBLwQ/vfnWEDV1Llz1FOONT2Mk1wtdcFiiO9wJpY+pNxIX1mCpmDi4
q1bFzyNHHyBHGkkWTUw81FlXtKMUxtgfGr1RRFNP4axPieQxEU9aFldQ9DSjRg90
yvxAvVZDU+4uYwhhBnUMO9R6D52WRRIMcKQvqRVRyTFyD38p4rlJ+YMxK4fL4hu4
XBMOHQfxt3DyXXJ0kZw/xPvwoAGTBU1liD5rClUPq3QGlAsVzJrVJ8MwL6O+AeoD
+h8tIxUkKO2tVerVrdeq7NKgQV+aGio8X5S11tOxzqp/ouDahTgbMGmy7I78mD23
gKfLksO5J8MrFLZYYc3/hEYQY2b9NR9Np/Lu8GbJb8diSxuD3gFdOeaZ7yQ6jlG3
jrw1eNzvJdSfPIK9cPvDL3GNzwKI7RNak/re7TLfuHAJuazseA34uUot61IwAZEe
YvE0EfW/Ar8HMa9gEjtNA5f8/38YU8X0Uvf5MJkdqGJvnQ/fq4TQiJXaoA8L2sX1
caeLbG9eciL2wUiTdj4NGwoBF4o/OeRPvdRGQ26b/f49GgFIokIVIEi88iLBuGoB
jiqYgb/ii/Uj9k9974Tnqj7tjReFV2OE9yY+p+CM4YvfC9cVYVBimW4g9WVrt+gP
ZjR3mQpPSFqI1u82EWIXrWeqJFvAXrgmbBrb/mpknwFgAu2YOmbTU9uGxcsjxHt+
NgB3XalC6tFNXGjv6s29BdQ9RQKzWiNkS8h9Nr8/x7+Uh93HExxTOgbh2WfJLe70
WDyweY4fkzwd6uFkvTPVoQw7rDsX26fVSQ1hgzcSJ/AGriO9vDUmpeE5Xinw+R8b
cS6lcQrqy0zwFPZH+q2uUZVd1EKNBWlSGZcIHW06uYYpxxyVH7QJuT2UzrRmQLN/
HgERoKxNOIesFYhs6GEkAvr/TvGXeknDkNfKGFgtFM6SgT/Sz/Bgw5EcmCk3rMWY
JXWOUfqTZRMuW+93EVEp/rAbM6uGV3ntp3U9GQc57tGzKBA8HgE87VPRTD0OXD8C
R7PBfGYm5q1lFcsAz71uxYfJ3YcKHhu+Wc28WHjsZL+jef+KfwJwZrQRira95d7w
XlaxJYjLJxN6DqJfDcVhqkRbAeKEEIlQon/1YNkeJjvhfC6GVkGNZwghRxmvJ3Ue
KRAvbrUT5qpFu04suz6Y/VE9D5aBV7EkcCE8aA/gOm7o28lVgF6LZGITmsghpcD8
B1WEcosuCR3cpcW8N/YmBoW9cyn5Dl2vY+lC3klnuIfH+0omhFquaghH+L8alGxj
yYI+tYcjx+se7/hPMiBbF7CAqgIsfp0cc5Y3KGFkrD1sMo2AqR4ZPz2gkwusbobl
nyAdIZjqvgYtc1ftSueoH68F2uQcxBdZubTndv/kjyr8x/qhLZVaqGMwGUhhTSdb
HfbNWNr9E43BEIFa47nNd9APH3tRSwWhh6uKIvlVjom5RxXxJzJMnaeR8P2wb9ea
iNROgu/RxePiH6D7xnydbghrb0GDF61ShJVHIvURfRZCr/LVgW7bvGl/mqFNRv0h
NyPOyyHFdEOLjE8ahWhCaXWbJyPgHCm2r5JpXjuO53PsHD/kCn8RbX5qB9PtP0+i
2CeKNtCHnDECumM6CfX1B92xGBmPY91x0JaMb3sR9Fuk5tVLfCWJku4SnQOJc1Y0
de1/nk2yRrSiWx3nkJzvnDoNRkCBhXbxmDtzcOBfU0SGkD/wuUWf4KEmZXt7oy9R
49AgLGye7bA4Z/dl8dcF9CW+JJqcY1pt8I0W5T29mrHnaM+AUh6tFGl85GXUbotX
vnWfuXgINVb3xenUj70HiFbP53mH5EWuN5+BIR/gcn9RtIcHN+y7fSDHLXhX7PLT
nqul5amQ2g67rlbaJObQN88PhYQAzwpowKJPcCW5nvoMJMGlKciGa61MBTTK84f/
o7/j5E0LagkqLj5XM/KhkWBV1kKz9jujya8RnL0RirVFcPX2XElLneuzLjiMgZnE
AOhYlOJrA0B+Z0tPXp2+O7QVkozcNDMnaYBWLGSBaW7lWvk9pRyFz/0NdLz1M3O7
1yYgqqRK4wfiTCILwHdPKTYAMDPRFGQjVX4FxqsnBkZTdvYKe7r/5NLUxRRdkGsg
02ht6cYz48h6B9mL/X+mC4V3yJdgKjD5e8xuQp2BME93OSDEIxnd1CkbQYzkNddv
7KgDU4VnG3KZTfkZrTcEUJ3Ujm2X8kTfazgRYUApib42+YBeR1F0+duB/cHCu2+F
7TvPItn0Y8Y2w5zIOVXAqQ3Kuy0MjN+MgiwIqdNjoraJT/35SRJTVLEJUqE+f0N8
tYRUkgOQ+S3G6lkiAOHSYT0mY4yT+xiLEH0ryDHHF4TuXodqg95vyPyQvuPCwDZJ
ZOfG8WCP6ljibxWZ9JY/3tPbEV1zr78TcnmTclQFWXNP9V62ZoDIiLOzRv3I0s0R
qzfSIQ9qtaSVsLUHf/W1GxqaDRaTWSbnvtfWaPybYJE878ReLM8UNOUyF+C1Zgdq
23YJsgS/rDftNxT33sEdXU1rPEgt6QC41eAoUbYqLDK5hCpfWrv4WSOAFzsftshR
PF6cyz1pspC/tLT75yk4aVI11JeIG+AnpO+oZNIVdaYm3LiKNMidu0VQaxdVa3Sj
7fGwFTgv1iSdDqgQ4e9dcNOvyqYAepnWPjaZ7s0b5g+yz03fPY8BvuTQPmziuD8P
AS33f6Flcchr4DSz7+zAN9lg+Qlkkysgkd8qC96RHfauP6GUNETtnQrNee83iRWz
e/FrY+iC9ZRq6hzmDcDK4ab0U+3GNRYoTiZnJGCQS5uh3zF+0VqCR+KSwqzq4g9W
K1l+ogk4q4WXd+jFtwy3640jlnlYyU1DJU6ilqeNgmil1Pjz0Re9snhrGpYkEasa
580+nNv+mdl4QVDibdWc/5lPJ6EYLcqqfUZGv2BSMBpcEtSfw2Xw6CNv7bZmqS5L
Z1Ec82HBRpSrGPtq7qD3ZH9cWW1AOeKJwnUuiHjHqF63Vzy7HLTOHXH362E+FVM9
bCbyJbqWB6RqfI3yTWH29fgKQ2Jo0YisAdxYXxvYdoAEvRTKCyIiEn2NjFMdSB+Q
eHT99s9fTOtVGTCDlbOQG0sMPPFUriBx5daNcpbE9glHzVT+chj112Xs9VJ20Ck2
vb9oTNcEM6T7HFBHzYpu7dlVtRHMhUVbVVcZMAUmW1M2eMMe4Y2RK2s46Hr9h++V
zcsAe97SC0pULQt2QN01MW7GTNT7jv4nyoCmKG8FP72gu/dsjfXrGXXFBz2D3RXf
fbv2t9sCMtqnQRVu10AkrQwUzF0mVKaWisluy2lMvEJy/lmPo+IAcPCDRh1N359T
4Dzw7UGu1Je0xVyKbmYExUHd3O9/tklYvcqlh0mv9mzX0YtqSm6DEa0BSB5IUsN0
cJ1Belaw+MDuKleGn59iPE8zbRBaEsQMCtuz3TtfobLwLAVNngHJPwlGsQ0LTjCk
T4hycoX8aZhqCjOJsw1k5jWEYWSkZJ/285wW20hYUxf2RRu2Ug2GWlbWu7OzzVQO
xI17Y8LN3wXyEM0E6tzG7t176XmAjgPZE7i65NOD4oVs8nghRAUCXMgdEoYObS7y
iMw5s6o+BEoTA8RTp4o/3GwTLyHwx9KIiwfEXXK+DIXJbytjcjzomAXY2ykS1syW
kTy4N21xUgwc3xWVW6JHDJcZ2Cvo+GFJol7jw13CbHz2xd/EQlCfGbo91AvFlCzr
QRKUSBEkYNR+uWN74rrDOkxyDFIyGkaJ91pcQeQT6JW4R+w1v3MO0DVI+11RsBWX
iAIkTb+KPqtrUGcdCmvs4JUTQu5Q5ZmoiPL54ldiB0m8LEYDXTHFFJiDYpIPpMxr
vXqy2WWVVTgLTbQBptgNuQ/7wTd6dJdHhx0T0s21lNgbCeM2wLcqduQjaZLo7Tci
+at5bc4FLxhLa08n8CCXGC0Q1RZnuo+p7IBQ1z/pVhYP+JYgEnS9Y49KOZsubTHw
fdQ+A5e6E8BjH5cOcckmmQ86g2EnHPyLvenuk4+5PdB7MzGD1u6K9tFO+wbeZqEy
qn3HpVEAPhPlf2at7Zu/D7oKWgs43n2LVfDHyESLFdBS48qUyJ+NKllsfBfccMhG
YCbnEwKicMCBVdfsSxtgku/XVezHQZKMJNtMbekkHahOawWhXNY6VnrrjENUP/eP
n04AkD1o22Q0Qlnv6fTPVzX+ZDoMZD5/navsjXmE9eH0CpgcR4f/R/eBo+ulPrE9
yu3ioHe7SOPC0kpsCiDOAn1M/1+OaqDP0yJ/mzYfZmJO1xZ3Cmsvzq/r6brTb9Z0
DpMaPSpj0AjJTx+6K0fmc2kdUzOwYx1+1kRqVSJxfcaQVszwzUmGcfX+OTS0P6nf
rUCb9AbI+56pO69liPP2YngJ1/yt68AL3xu2SdiM5ztYYWCoAsZibCCtMdgM0wyP
b32ksWOVN9y7UUANpZj/+OfKyIw+dTxVXbr9ImxB4bSzF7GmIJN7wuiO7nRCgDDn
aRbtQ64LyiuYji1JwNme3NyXsNeXCOMpht4Ir7VmiFFNaY2IBt9QNRpnMyhZeL1M
MO/L825+SDfINKX8CSa8x/Y8vvghBQQMoLsH7zuB1i2Fmwy20xfRqUlw0Sa+dvXc
TcDOmPotGs17EdqnPPGHqSXIMu/PmTD6YHBxUsJSM5eUXxxI20aJZkATiK1lSj74
2uP0mcSbczGsLk422vSAeA0Twdf1KbLZho5aqDSJEn9rbLzwvYmTfOFujZ6iqqMg
k1p6VtyG9SHtgPPoAllUhWt+EwP9S0I1OoFePCGpxhwwNVJE1iHFY8UHpxnYqb3i
dJdXqhldHuLR9eAKQIIjrT4pbX9pQFkof7Bb4JGsJGE8q8hX92TO2wq5oJ2XWkLX
lzJ4VeoEnPnBjhUbpk11UaZOO4jabVaw/MbP3LNo1gDOqUIBqQdYK/r17mgbcckv
tpJiGUll+8xaJHUOk5Nl/WaXnHxb1b1g00ggktb3mj85YG0fUcgZ5uGDCG27aMrG
vKKVOGfZDDvl4rrwEFbMo7ak1jFp1EzZpe9+mdqqwW7PSNxTkuXf2lOi7YJAoLzz
rBvkJHPNFN4ASZShFsS73Nu4nCoXmdSc36zvpZPIyeCL7uhV8lR0CbwBugofC180
UMdQFX8muyjbYbgnkhKKQp3+pQCYmBTH1X/6PV3HVf3CVT5YWFzC3YM4GBwGnhk6
HlVDhD3CsEbhGpo30sJZFzFpElVNA8aplVkzukERdUC64ST5r/rNpJbHIoYdnnOl
R/neCpTjU60xXZ6rGSw3PRwdn6TQQJjrdivSJuP+B7hJXCYrQ6wVsURmvi80IIZp
MaQp5AHeFB4+zcWKTe6nmkkHdABsa/I+bv9eXTdSaZ4RsmWUTfEpebzUpy7OJolI
/x+spcaqyj/yXawW5an75oCYKDiZuJACTZM5hCWPDr0+MOUFdIYh02/MpYXEEmCa
ekCtncFayrX+2Uh77eGmLxX+dRFrf0ukXrt8BCV2RjxltmQUdKLdX3+G1TBsBqAt
b4NMK3DNviRyom9GfuyHzJNOImVo3XN70rrpEnFfYxxLgDEJ65OKP8ONreY/AYca
fPBLbQs3AtpOymggdN0Je2uxe+j533BdTPvZDo4LmNe56Zj5T78rxLiT4JE4mYqa
Cm0Zn4NDfOruSGzG3xTnO6g0aWotsfA0d3ztaJVhL8pqZ5SUutoQ3aDa2PJghL75
Y9WPr+7VBaF+GksOyfap10dVE5q5dQTpRDMkdijavgsnLEkMvUfkCXbqzeoqgIsq
r6h/eeWgu8wOaSb9S4jghz6GCjIQFIYTBaBajmicpUZ6dwXTUZnyjF15qCcb5eph
1SfU+BCBfiYvwwxcNlufe2sI4w2khi3EmGjzt2MbIpK/DDhaEbUZgXq/DIOo5N6J
kGPGjOmjlPCBWE80pqRcpho0JHDvwbbVHKYHKI2eTWmQSV36Kowjmkv00JXD47i9
CY+IHBzK6Lvo2u0RG3yIC0Sp9lWdke7GflEoxEJbt45P3ekbkze0MiIdRB+vUsPg
CHvgc6Db/9H07JnRLWdj5ToOBkVylZWCseaeEQMExlPD0ofDuCcIhjX0giiIGrsb
PLMyR0hRBcKax8NokVUk0SSfZGIztVDB06bz1+elXnAuAOpTNlZJ16MCoETPiAet
hHunUYqD9thAlyNuolNyU6IvaT3Yk1dxS1RVPAwpImZHvl30kUk9FRpn9iRl5+K8
pAu9rrfCwOh2ibl7BPm/a9yJlwonkMYDs2m/k1TmJnnkgQq9ExTlGu2TpjD/Tf71
4V/UFeDNAtk5rReMvQwDv0X5pz/2VD8y5YuFUm3T8rcxDwtbhHs0UkieEx3mFw5H
h0kIF0lZ/91cpNKVCau2httdWNN1tJd2jlK1xxut66jUQQN9s3UW2YFyVNLpEtvK
RTF7EoVg+MW0MvKdMeoqrJsGnSEJ6nQeg8NBBfAcgnO1pmevVvby7/ghOi6HJFPr
eL89xeI6+ny+IfFg3kYC2BSXA3Nxj+29qqiKD0e58fz6j7VTRBHJmtyKePUTxRT9
bHHTljSPjchOkIanx52/rWoXgxMOJk+VnnhZUNqr1qRJjfHgfV7JOJe4OFYQiX4w
DdM9bZv0wMB0sBtxr7u6ARFrLnHAPPS9N0aZV0PJyFMT1pcke5hZYlMpf5cQ4tdH
Iz2JetA3zhq0lLiapTvGkCrG7f3gi/qnxOdD++UWGUTTDiNFq8tPHpzbtHqb0C2h
PRWjWg95ia4iipmf6ho+9CM39Y654oaWYdF+Tb6dKx0DyGnZRk29EmO02wUi+XUs
n63OHaA1hxeO5bnI4crzynsC1qxoyh9lZX2ngki0LAIctdGSUB/V/84k1j9TqdOC
XVGIwlpUHKe77hqYBck96/nGt8O2nUISqwcbCsxd2XwDWpUgHTySo4fBs39RlXiR
WfK5DXbUYZcCxk7IkFK9EW6FHIxjjTgQmpuu+lYcVDwNkErU4ySfXizRF4ayO5+E
7Oox2Sv+xSVJKKMxRPIQlQ7C2NBgrQaUFsjjjD4vUzQefeplvCNC6En0LlFzqNE+
TgYLEGkejhkgk9fdhQewEQ==
//pragma protect end_data_block
//pragma protect digest_block
EATslI0w4fX39XwjIYynA/mNxjU=
//pragma protect end_digest_block
//pragma protect end_protected

`endif
