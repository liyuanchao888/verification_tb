
`ifndef GUARD_SVT_AXI_CACHE_MONITOR_COMMON_SV
`define GUARD_SVT_AXI_CACHE_MONITOR_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_axi_defines.svi"


/** @cond PRIVATE */
`define _SVT_AXI_assign_new_state(cur_state,final_state) \
   svt_axi_passive_cache_line::cur_state : new_state = svt_axi_passive_cache_line::final_state

typedef class svt_axi_passive_cache;
typedef class svt_axi_passive_cache_line;

class svt_axi_cache_monitor_common extends svt_axi_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  svt_axi_port_configuration cfg;

  svt_axi_passive_cache      passive_cache;

  svt_axi_checker            axi_err_check;

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_axi_port_configuration cfg, uvm_report_object reporter);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_axi_port_configuration cfg, ovm_report_object reporter);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_axi_port_configuration cfg, svt_xactor xactor);
`endif
 
  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Updates state of cache line associated with current transaction address at the end of coherent transaction */
  extern virtual function void update_cache_post_coherent(svt_axi_transaction xact);

  /** Updates state of cache line associated with current transaction address at the end of snoop transaction */
  extern virtual function void update_cache_post_snoop(svt_axi_snoop_transaction xact);

  /** Returns current state of associated cache line */
  extern virtual function svt_axi_passive_cache_line::passive_state_enum get_status(svt_axi_passive_cache_line cacheline);

  /** Returns finals state of cache line associated with current transaction address at the end of coherent transaction */
  extern virtual function svt_axi_checker::coherency_error_type_enum
         get_next_state_post_coherent(svt_axi_transaction xact, svt_axi_passive_cache_line cacheline,
                                      output svt_axi_passive_cache_line::passive_state_enum new_state);

  /** Returns finals state of cache line associated with current transaction address at the end of snoop transaction */
  extern virtual function svt_axi_checker::coherency_error_type_enum
         get_next_state_post_snoop(svt_axi_snoop_transaction xact, svt_axi_passive_cache_line cacheline,
                                   output svt_axi_passive_cache_line::passive_state_enum new_state);

  /** Converts passive cacheline state to active coherent transaction cacheline state */
  extern virtual function svt_axi_transaction::cache_line_state_enum get_xact_state(svt_axi_passive_cache_line::passive_state_enum new_state);

  /** Converts passive cacheline state to active snoop transaction cacheline state */
  extern virtual function svt_axi_snoop_transaction::cache_line_state_enum get_snoop_xact_state(svt_axi_passive_cache_line::passive_state_enum new_state);

endclass
/** @endcond */
//----------------------------------------------------------------------------

`protected
-^9&^LJQ.)503JBL&,FRK@0JNG\UYSN8XUfcSD)E(I^6ZDV(A:Y]4)X?>1[\Z[4d
>OgYXe.^TU&7?523A#K\7MJ=N\G#Zb63+G^AT4,4WJ14[@CGdCSaN)>6T1O<@2(6
0@:.g3X5HG]S=I&UNd<+BY+YHE+g?D?f(D361APQ6)VdXUELb-:1(6SSSAMNEZMC
,WW?ZS;[SUE_J,XGf/0eBKE1.=JXHFY(]JH[NA#QQ,,gUdCc^\=W8HC?=G??J^8>
K8e7?,Z;:\X5C]=RR=a?QHdW))?3PgBW@[_Hg\+5,]<G\OO<QACRf7)f:=e=-e96
A#6WCCM=QFa>F.eGG@97G=CEFDgFa&(U\(O8N8U_-CGAL=T1dM+6:S^7X(X\c-d<
g:=B9+24\gOJP8ALgJE(f/_IgTIaHS:_MMLcgIcPOR3#2RX]Qa]#X+f;+DeIgG&5
NV16bI0#]_9VG1_L,[F3LBNW>YNf8Db3/acO:JI>3SC@5[T9YHH.1ZEbaDNG4BH)
F792=F<<J5.4H8&66>GVI2W@e?3F(85#@Z@XaTP1a+C@.f0N0/F6-+2@VBA\XIUF
O.TDU@\cB?K1]ZROG/2F5\VESOQH#+^Xe,59^#HcQb-285G.VgKJ5L;0TT;KE#D.
(3H)\3<KeZ#b62UY8U0#)00-R/4]I=T^U:R7->6@?OS>0I>HH5N:IY#Y?/\#a#LN
Ld4RV:-;-MZ6_/\U<PC]8Kc0c@XNc(beI[_1RV)2B@cD?S9(\2#@X1cd,)AJbPQ\
a0;UOD5XQ0718IBNe\OICD;Ed8R?5-CU,Y<+N,>F9<>./@D@#:[Pc82#S.S??DdS
8@L8S&:7PC9W5&9<7^?Sg^?CK7)O;4@1&B>=YLK9QM^\./]Z^+)9-;e?5e=L?&^1
[gPZ8T@.U1gU0&_4ROg58b^VG;3d#)g5\9+U&0?\?^2e@X,&0OKgHRZ(F,L=M&9C
W;^c&;\L?T#(Q.Y]LYXgX4Ob<NMIU5Q5:)=D3S?VUSMP;PS<Cd[5B2D2^+aJ7Q+,
QK.5daGU:54.>4-EZg\J;D-V;DEcW\<L9e\]1)U+V^_\+_@\09ge7O6J1>P]A0V&W$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
C#^##+@.XPF<(4F<9QfTROQ[2G.+5CS[QY\NCMOXJI?[T<T7F[92-(B7F3+4T^Q^
c\[fbA?(EF#.ac12Gc]_Db:<Kf8VWN1]3QcOG1D7[>-cId/.dcZ_[Q@B\HK+?YY.
VI=2NT([fU2L]@_C,M280OA.\dBASVB-;#DOX=d3FTcS4PT..b\g_XgOcaD^L-#A
@c7e[NEBGB3e,bA>\[Re+RfY?Y5c21(:M2_.&=ZPE/+8PNcYQ9c)AKDZ7DSWNLZI
?ZKO-MFFZ[#.@:^+[1(b59N,Y(^).K4(N0^[.O;_\T/B)0GbKXDe9JD<C69#/MCG
V]4#.8dOK]7DOH0:4I-Qf6./VVb1<NfL^=_=21K&NT.5Ta>1^79?b78A2C/b:,\H
=_.QdB=/adOBf[:BDG.a4DcGDG#&&M+Q]VXO(?=edU<=bGdb#ZNT35CO^(J:dOVC
=9d1WSTZL=[(X&;<E,N2ANMADPS&b=L&[[&/\>XMR-+GCaf3:QL^b:-g8T9P7G]+
X7aC0.XJMIAP_=NF3?I.[5.<^97a8,NgQJ+1c2UJBU8T.V(&W-FaQUa,6HDaE(^;
eYNOS0/?AN+?/Sc.F[C6_EdS9B,+?\XFR]YES<B4N\D(CeR8E9AM3dMG7d968NcK
NA=E49eAfbQ..1+gD\]]@;IL:F?/0_=<P@8a_QRYcDc3.5#J.WVdVQ[TB&#TYU?e
1/L]/@E\Qe]3GaWWHFVIH2QV>&<L=ebP33?I8KNaV6DRaX-.9Y53UaT#-@EI[)>I
dP@1Y/MG)&9GI7XBU#^FUQ@OA(0AfP/fV]@FGUNJQK7MGf.J7Ic/T24^3cSJH@[N
g<dI)d:O[(KbD?P;Pe2>RZVbE/^ZZL]M+,\Z8D,CQA1O>cYCRDMY\[FL-g];MOON
aLJf6J&b74I3:L)__@OY^e;1+&U-&^bNb&7:ZUJ9B8#]JX^e>9)>9f#WDLV&+#K^
CCOJ+eg3+:[^D@c=7S:GNM3AJ6EMf&Vc#g\&SG+.;2)gFM#1)XY^N7e=Ze:?0=H-
3Ua@0Fg.O4<6D(\g42;MfV>@db5d:2//&#;[Ee/9,5/B0LD)a3V;JNZU-gNL7cTN
DNHZ)AS[d=1Afe\8P=P0cLB\I=C5Y4]:Ef&(-O_1,G&UgA140TSF9DWBPQ83YfE?
c39EcMLc/5\d?d\K7gGZ3)Zb?G#>bO2OdJ/4<5#,IZKP=,0b-^YG/P5]a#A^/4RT
8>)^;]@c0]1QAY63+IJ/;JX+_[4@gL&8N1;_N0W@PA16ZV5dDf&g/fNTI_fe+^E>
cWMbK0^)D)(XQE?&JXTKb^a;LTcX==+(Of,g=Y[6^1ZB>B_1P[5#=\9E\2.ZS4TQ
DZ\WEY)#FR,FKC32,LY9MNMDg)BV/C#]0-NZ@caVYJQ7=O]N_H[Sa\G7Uf_;cP)\
-,NRV?E=4:;S9H0/5KC-JN0EK1PDE(D)H1F647,>O_LCfg?fSF.4VdB(dgZ0?V]A
Z)7W&BU3dFGgB5fZ_2GAX&U>>XNF0fNOYH0XAg0/ObJT6-_Y^JRKQd9]f?<VJ\(a
?OBF4[K)YM#LMMbfDRV_FB+=aS=FdIg?BR[bfYIGTN].C.WD>=J>FXUU(.^Kg_:/
,JYN5+B5PaU]fC1^^ZG1^ISG^cCQHg<?H0,K/:924^6ZG@[5d=9:e@aWV39XRGB(
]f,,eO6-VAM[MJ=T:-<[SK\#A7G@/YNbdXbFQ1(8<=.X;Mf446>b0&]O<L>J60_#
.J]4+NBJD@\67eL//MY],S45#PZb-C9>/R7T9RW)a8_.&cU-ZZF7VFcaW=f_@CRK
0O=)H6I>+CH[F21S,0>/FZV#U\;=Y)K#RJfML@B8D.N;.ALF.-J6S[e\FRGUAT=T
BU#6C79<K9R-4P1T(EO5O_]\ENU1>,GJU&<#XLcY2JQf.Aa3R#<:Be)/6JTf):&T
e;?<IKNTJO;^C9.]GEY^=/;W+5]/7E5ZbRb^5&X7ETe[<R(_?gJZ<B)bC]9(+S9L
,O6_]0;C;g]=B6-g>\#aN]]CUQ+QPIK>e1K1,JDRCEEG7O/3G6+X)]MI-XEUd^,J
EK<(W^Q&;OK_aNVFcL9\?cV6BC6O.dIO<gYQIDWH&:M^N/9E\CH1,A^/>g0]ba\J
KA-O)\6_LUI.^N.721^>D,JNJ7&9:De\ccZG=3K+,U\GFV.D:b>2Va(XB3X0&=16
^2a_JY(2H&K^Q>R5)5bIZA9FA1UbC4K/_c[-g3N.A(;#9#/K;Vec3-B;30<K3QBa
BZd.P407+1/]+MSe?V:aWR3F=CD.=E1)DE]EIAae:/UcIJ);J-Ff\I<)\Q5A]DfZ
>:X8f):OJETJR/1HO1\&U9-_aAC\(4,;\4a-[PQYFXU5)ZZ<fOC4EPBO1N#GS,[T
R?43=D3&,HOaQV/]Ca])[/@.M;^LUVB;VYe,2B@QQQ^;76aab()7O(EC>8a6#,,7
Z0M2d1HCS,15IKYI>EJ_XJM7eQ._OD]e@8bDfX)3.FIIcYSTdBMGDgYg0L]a=e_8
:0E2dX\b8ZbY8b10gOecRSZ,&CRUJ/Z)UR(KSfXI6g=]6G0CO5A6KRc@3e6c7.MH
(_@D-LPYV<44/#7N:b4B3+eZ<Z\&U[KfN?d2=CLA49@_;#PPUVgI+V@B,YNR-@(M
?]][9O:NTafOL18X+_H)Fg;(?eaUc1+#3^ee]Q;+T>\Ke6TC-U>:]fFY<7+K4[OM
=H./d9T,OL>V]aMc#gR&DC5F+/C1<5:NbQY1GZD63HdZ;A\IeE#g+_ZO5A>F@2)Z
-SL(J_2G/+P,dBWT9ZAAA:I:d6#44B\g.CD/Ya4]5bgY]c0+#ENHESV>X6G=:4)C
OGST4e295<N#VKJHPTN1UU^J8P>GSB?F1YDV\Lf,g==_Sb6\=5>EcUaF&If2L.P\
7@:069c7=/9#UfCN>YPIW(.T=DM#;9[cRLGD&-d8W@dc/[:SF+#B5bT32\;bK3cd
56KGYAa+YK/;g6Y7&VA_Yd(9H)9gR9T5F5AFf6>=QT.Q#0\8GM,&KF/?[<\aJK(G
LN#P-Mb[Y<TS3+C9)L?:R>0@7e3N1/+B]3TPR>QK+QHQ0P-2&[HT]^WV,b<a-J:E
7P)De9DBb+/JOF9@g2<Ee?ENXc)Ob5G17K)N\]Q\IA=,cXe#1JIb-N8/@.4=dVK-
+D:1VJX]R[Y,?]5:MB7,C(U9@6&)f9fB91cE;D4W2G_6\fJ@T>(G.(Ee)&;1Me0\
&[UEdER4B1QO(ZD@68e<FYM;QKNTKHS45J9J#N/9fC?DJ_=5-.cP#QeAd(+3D>;>
OW75gIT/EVdQ0)Y]QF&A;[(1eGGVRgZVKIV<G\H;^==3d/gJ,2Z8?R_KSCC(ZYdJ
3-[)9#gF0O/6[DH=[R]_<9EM(+HR4AQZe(_CDNCc;-K\,:f[^N0#C=GYJf9aVJZ+
1>PH?)DJSLCFa6He32gc.a9)4SKBQZ3X0#bWMGc0(0ECcA>E_OT\de?&:G3.E<HO
Ca6&1-]EN\0;ab=e1H:823D3G3Z>)>3=(24>WcY?gW#e@MD#8dH8_#)7GT1CCXOP
&4#_GB^WKX]#a54eDCKg1:ggX2Xc9(#TV&S.O&8<CE4\e2]MT#Z#2FPB4N=EWE?4
d6(@1b9QXe<JJH7N<Wf<:W0PTOd=Z-ZGDO5.g&S)fL_KTPdV=#.\K-=VS_A:Y:2B
@M3@J8]dd(2>]BFE6);;9VJ###5UTcC6ZF(:<;038&V9^2]cB<g(JgcJ0]R+EbP<
DV(=,3INGD[=GEeQ>.Q\VW5GX^+QC?&XYL\g=5L,QM8C#M2<aS@7aG?8Dd6W^9_O
YSa8/25JTdPH[?SOV132QG4_8@YH+D8Ic/XDSL-DW-bYfG,/-;@2bNa,#WS.,<)D
7^A&X6PZBJf<HAE9+J+;Y=V-93Y[d-SC0-fEQHdFg&fLF+BFKO^1]K/@XF1:^9UG
aU=fc3-&PFYCA)IG=;4FTH=O).O<B,L^e#ZIaY.006/3a_UARb,e.KeWS;_RO?4;
b@;,E[PMHGJB7-&JW_Y+>0H(VZ@B[[B0FTJfJ<>CW<EL(60:@FU+eM8:[)5WVY]L
Of76;BT1GcS)=#[Caa9MJ2aYa40R3FL7IXG#GG:XBGU32ER)6DU]GWC=/_GNVFCM
T)&NAXa:XeSb&6eIDa6VV\)6BePT-45M)5Q#aH^U)f3,KGZ(3U;L1E-D<c^KefAL
#.d@3LHMZ31O=6B#-gXe4GF<U,DX,UL51c=(Y/Q^f)(UOeAXdLa.[Dg44M_SAc1;
K=fD<C^H(T>M<T=[=.b_afBLT90(7#8_5E3G(g[@+(IQJdZaIGC,A)X1[8PF70BA
DGG^eMIgA+5#,5BG5dda?FMOaTJ4Icf[I5>LeXRa9R)_3E/U(@I6b8.PV#^2OTN7
/2=>[#FCA6M#8)NFJE((V5W=G,TXZVAf[f\3;3JKPe-8AC,76_.?bG6>F771M-5^
f<O3WT;F-=Rc@\DaYE3H,3.cO4e]aYDgBQgZO5EW6Pf2BSQKf7(MD7c2bD8<01.(
&>=SY-L)fBNK?G.L0I&6F7LLHQEc10;Re;+T;a<]3bLTP)WAM<E(KMV8P[RTT@f=
W8Ib#SO(gKGFX/C0\[S>d:d];01&RB\)-M\(BYA>UH^>?>_?.0TaIZJ24+Y?GVSB
@2]7:d]DYZPfB3P4R5F(f9C=d(;U6(]-[^PNY_-PB]7EMbJ;O?=\bD&TB[YMR(,^
:9PJ@ePETVQLIaZ(<:Xd[G]^H\#5Y@2A>Z6]IbX3^5M1,X>X9Q>0X(1gKRPS>3.1
8J->PU?O)>O7C>37CAU:319dcVF9@BT7>[.8=KaV33_6>R<SZC931YPN+RB5::-R
D_YK\c)]e@=7.@VLB]fFIRF@,)&)H^-I,S??H[AIb36NT0]71_bgVUIbM?XaY(3[
[RVgI[_^EbIY0:4B5-RK?<Nb4J2,[EAWgc>\bcTU_YOUS5S[Y291/)dNfM8JW6J:
EAfC&6Y7-1E,\0/6+>C74]b[]ZQ1?eFA6HfcY_],4VASL>E]GEAa8UG:SMbPGb@]
QL)Jc\eEK>G/=E(Q_c0JKGF?BfR6HFXF)IH+6BK,@>CaKD/A]GR-IDYXee5G]OP^
eX3CE:C4<K[7X&3+<Q^ZQDV4H9US_f^-f_EJQFP&BCB/O>_2db[6ggMDeIM+E)d@
QW5;UDHZULb(e@eJ3);I4^P14BN&J)5-QY(G+8V?B&C)<d(-CBRW^?4QdDbV@E(\
3.C)?X+HZ60M,dARA0;3,PM2S[f5<V[0.KFTf(V&_]T641dFgg(G./ONHP_6B>9>
,OH_O_]U\V/DaCB@R8b@3Z?Dd29KeIbaVIL=0T>9[4;caH1(]ZL^]NMAafHE?9G.
Z1Q2).aHXR43G[>dRG0Mf=5\.+[-,F@I)V:[?+).,4=L/?,e]>g/e5-=7_&+GTXK
^@H]S,:/bV^+W:&,P8NP\I?&C8?FS2XMF:c):9<gA#O#UOSF8^Q/O0?D2ZC#/U?8
McV4_abV>ZG0IZ6HLe4)Tg3gJYV.M,Wa&F8T)U(^?^Cg<MQcIC=?#,:YG.D1Qd:A
-IB+[;W2C<E>L&RdE0R(>.,I61EJWV/29<:?^B?G.KTCE:#/6L2C,<CYWK,3;f&?
YMecTg?0,a7HS@PdYMbH?I:BCS?9bDSZ1cISLI+66I9W\?#K2L;d3<S_MaBM(/bW
]8W,@]YI;@-@N.B?bXT?Pd8(55F_d?28IfHV#.1KLd.2Vd<PMf]J72db[0?,HN<T
ce\_7[5ECfUI1R0@PZ;QNFG:=@(MJ+FRd9CGGG=f)X2-EW.2^Z?V15Z@7PKT?-Q&
M6AYF\C><_Md+E53B5-R.60]Kg#A^H:07_e1^J]YZ\NS^/3_?O(W]=_ACX#f3V3E
#E]+97,TD)L+SBJ/@D:0fA?2X4\G,@2aQ5_XI>:@,RdJ<)5ab=FYZHB6.(O\/W=E
Q9g5QD4G;VaHE>HU91&-JO<SVG0160B?0^-SS;I)92H^P8)3e0-0/VP>V3RS2_^0
f2:agJ;8VRQ5C2MOF^M2;3<0U6B9H<IJAIWS]W4=6dU29FZ]\+CG^EB[[BZ#MM/d
Q[N36AF:e4\/BXE^P>,d4cK?S?IfQ9AcFCTfXf_Y8OJ=CIL::T5fB)PHeO85[=+,
#O&74;G16A>f+\>DaIXW\[]\d:(fM]0X)F=C=#([\6/<@TE0Kb(\G,=]bW&V(J2H
6U>QE1TG^\TfXaL^.N@@XIeZB-X=cM?\2^-IV>1;aMZ0X0>=[f=2EYC4XbZ+3^N1
^;EaN(J6D3Q-R1A.A@JEHQ[[QNdG,#?d5Y]:+WMH4X=5F:0T:JQ=5]A9BPJ9?V^1
N,4(fW2&];MeQe?M\V5_H6/:dXW]&gD-HPJ#6Jf<JA?Y>)dN?GO5eZNaR/eB2_D7
_#?C0N/@,]_3SBLSWE[=V?JVfNZc9NU/6\Q-MID/1+Q+e^JB3bA9?C>Ic97EDbaa
:5C0R^=Uecd304()^+DP.L?\_1KaHW:N^:>KbO_3D7bV)Y8PHBHM\L/ceAdg)6Tf
A+6QM5RC>0F/bgH(S+K9FY\IXW_)B5X#/8QB91cK<\4\Kadb2eJ5MaKb7#-(=(=D
\X:FNga#]>Q,PBKTWa0/JRP,RaPF?XC44H4f>ad[II\+PC#f.XVf4OD7K^8QDNT0
1G0Wc-<NI+XX<e#_0e_>_UQ118DB)G9A>B?F&P9;(E?RZ3X5H/JQ.,a<2.Df88]&
)#QaTFW5d-]N#)]9.aV6KeX9K(7:D6T)40PI6XT?9Rc<W(RX?@86VN6Wba289e,?
JTD>OKCQgfAZ?07L?<W,38RRJ:PZ=M@5WEPL..]HaX;+L5P5,<OPOb9NXgcd_0Mb
-.QDfbEb>T[b60G&<#6V=^Z3/5MM0\0FdPMFbUE##Q)8(gWJSdHPfXR5,]8,O(?X
VE#Jf>3GPR?B?aTI-MV4:AW_/0]QF.F)#0?eJGHdZBTXU.EF;AY5>PE6/^TafGUP
_@/W&fUQdT=IL#VEW^-:5^e/R@\9\X&,Y;GT3H\3=0fUUCPfAg(_D6@;F<P](2:&
8T1Nf+GG/_[_&^Ve7NWW+c<257==;U/YV1WZK-KSc/d_2ZOCM2YP0K(O4\KbWN7L
I2cZEY^e9f9\8:=_HP+E-T,E3U68G?_/\?Z;fHC@dWH_VJSeH]^+>\-QUd^#B&;D
Ya44]W0<I9C6<1aC=U]M+T.f7L[6ARM/#Og70d>>],3cZ@aL1R,3a+X<.ZX]0)YZ
GK.6)H+3a:P6[cg.f>\VS&Qa0H,)<W-,fgX(Ag_+;^=V2f_X4\(aO4DD,<=[(Q9,
+E@J1?WeE8<AC?P[4Cd&]^bSO-L;]^G/HNNe&]PX,7S5ARWf.D0^0bYI3Hb=S@(Y
^7#9)H:;M(d22N14Aed(Q02,,JHe3IC611d&4A<,5a]KDT,F/c)-WJ/<e9AdK,dd
\@d:Z:))[6K5B/6\PG\31-.SSW]<,WU6UI)//fRUe/ZH[U?Z:+H]1:T,PPWd_gER
:S-X>=FK2Ldg3OH+YT@;TS^D&(b2F;>YJ\SGAS,2S@U/9c=1(aV4GI[,#X)3GS7:
=0A<_4YAe\:+>S^5#:UEV9?9=&Fcg;fOR;LULJW0f.Y>FNKeJF>)>&WUWH&O;K-Z
-A4gcYafYa##O)A?RELIaZW;\7cb]L7IIf7]PMfGBcR)BMV98_&QNaK<Y^[<4a2T
.L_0=4U8BSBQ9BS<S8aG4=Gc2-P4[<4#_-WY^=@D(1E&N;ZW:#I0U#,;Da(1fbE+
/I@VQeG(6@IIBE2[@#-LM:e3.P2=7f^36G<BJBa3#5@@9X?Dd1;<87#Wg#VX+c8L
O.VF?T)/:#_2YJTEQaSfRQ?4a.NM9MV-PT@L(F[1RcJ=AO[[\(DWZ:5WI<;_0B[6
3)P5Z[MB,YRdXU]\#33>T\M&EHPCb.7+SHX)KGY;CJ[WaTLEG#cQ75gPBUO2[(C+
HQ/27eP(@=ggT+VHQA4Wc8c1a]e)fZ972<L;)5FROI.[eI,A7FFH2SRY]35fJ#M4
eJ@ca1+5OR?QGfY8E..MKAUcCK2d?RdL7Fa\eG,E5#NMX<B3TJT05]QI?.#<[K/H
@-.+V4O/9g0/I7KX)1L8BD/<Oe8_,-c/SY@4]RS_7\O5;A=[6+Mb34^<)8LLEJcZ
fTUeaI.3L[7M?#0^H\OZA&T1&(X9LX,\(37deQa0:JQCCMe8VRXI?V];5c_@G\.X
9U8e?a+eCaB:+F1If@;.SQeN,>R+5./I_TJ:[KU/E)VJTX(Z(a/W12eZd8+Fcd3N
K?OA[S632VU;.UI,/(CXL;(N>W>[KFD6JWC\I1,M9KSCDRN[[::g@C#-KCe5ec:U
E..b>W<b+67@TMg6.<Y#SLdBbN/QM+Ce2[f0?\:)/LZA[@N?4e/J6][T&FAe&b&G
I#TY8P\Y;e#Y]:[cN>+5#Q4(UT<VR/5G?VC(EEJ,)aQ8aT=:0N2N5ZCKDeeNSL+a
,d1-WW3Y;M\X(cWg@.)TQ=\AfBVH=b1BX?d@.HX6L[ZbLOB+V344\L?9Q=;:X-.@
&4c5ZABQL>F2M:<WHS3g97+[Va)JcHeE>]OJ+GD3+cg_4(e550/]_J.Z>7O:NLcg
NfF667\geK5baL@K._SU;_?50>P9E+a5WAb]P5c+]PTLPP=IfU7//WaD,LBN2-Z>
E=UC?\@T-DZCTLVC[[Sgg61<^K<be1aQJ/XWJGfR9O-Z/5R#F#<A?E.f5F</LCCH
V37Zd^VMOFVGI1K)deRH;V\BJBWFJ[]KSTY>TM[:8g8&K;WHY<eB;H-:\e\AbFJS
8B4?7X[H&E7)+2K0>0XVfeY:(=b-e@,@8<YAc2BYXGRGf_FL_T&=dIR96Od)FR+N
4-J6G2?BdSI#MD=806=0W#aILaC\T#^OeL_5bNPFF-Da=3(ZcPREFQE3(-TOQ=_-
&49]-9QZXGEJ,JRP:1##NY<91P:0N#QIMLK-cIO=>0K==.FSKNBM[-Ab(W1UL::C
81S@,\WZ[D;b?-WQU1(,X9=6P?@=/Hag7N#OUMOG/JHNG,cP96/3W-&0=/X[.N\4
M29^CM;V(^ffR:<KB-?2AA?06NZDbLQZW[g@GOJ=Za)((U0^L3K=1ANbcc1)^U]A
SA6KAJ]c650dC9Lg[d=MM&cfRF)GB\,g]75Kb53aa6@ZR85ab3FR<&[5B?0)UcQL
A:]aA0LZF1ab5N3&VM]ML5KGYNbSTWg4(e(Uf-]Z5#ARI]b#PBV38RgVFV4?D;K,
[5gT<X^F,50K4d5?4>#:J7UYNKgA2^R<PZ4gL4,)0)1\&e8)g+b-Le/)5Z1N,X@[
3Z2\1]E)I5I=LBF[Z6G<S<76HE@g74)f10/feeOaBONVX+e[LK-)>]851;YG+>T\
R0dE^3DA4)+-R7HH,FaQ&Q6=F]AS65JN1dGQ(1VcJ.5>0::Yc#:7UK.L/EA)9N6T
]5dL;8dIYGd46\Kg9?:3AT\=C)N47b,@_IP)dKcB97+.;8&dfee\NZ@dMRL;]-G/
Hge4?/J2M_K]Z1#H>W(c9UXbb^fS[;D2+AX0J7V2D^R5g)133D<Jb4+#A:H54PRf
O4QJ68A^,=OcBZ6b[bZZJ(Y[P<#5#ZFP(Gd8/GK2<87+WDT@aGSe>(=?W2)F1fFM
,TGMKOe,8c5\,S>GLMO:+:LT40O;ON35?_S>N3ME=bWeF[0261Qd98((XF;4;cSB
CYXL7.dA3XM^[7ET_0O:g;6g<UCA.X4)\Y+Q6LKcP-OPQS_B;@2\=LfCDO._QDQH
)106@>8BaW28&4FV?J?f&_bV=NK8XT;(>1gaSN:M[QH-YKK2adP.O\3P9VDOQ1&6
egWQY@<.bF-eaG>-d4;6@7b19YB?]S)CXf-(P_e]\WR2G9(e(e@N0S5QgZ:c3-26
N)<GJc+\@35L5AHd2FME#S\--[UM#^B<TIJ9fE)ROa<^1:Dg?6\c;5P)EGV:BdL:
c8eH-&P4IAfRVJe#c7:VeaD=gd6).(e^^d0G^H7=JX#@QU+HN/YTFS&.GJ:a\da?
+9>TC#6XH5-fbA:]-G.MfT<8JCQP[ZeW0L0_gd2O.1UGeeg)#b...&3Q2(2EW;Xd
)[=6:+:aI.C)[Q0)#LO_U^NZ1LJ0.0XB<TK<[5DG3SB6CLT5bHRF:92fZeK/,aAE
=Z5D._W:f&>;agOU4,IYSbH<CfS>e;ad;\CNOCQN)3c[;WYI4Q_e1a9(.\+U(S)O
1a)Z<OXe=,6@MFfd6IV@F>_(AH?E1A\SGK@Ie>-+Fd_&7F8B8[494R#USP)2\K.U
S]4.@O+3;8VJb2VM:<PJM>eWS5gf:1f:GL)^G]/T\Z.2Ngd(Z6)_/g5VI?5-^IP/
4_7W=F[_beD9L5Z?e:-&Rf4&c+6e:M&NWe)87]Sd7@142-=P)-dXYe=c]9fZ:=R7
]S25Y=@HHb5B;5IF_5AWDSZG6/P..4XHZP,6.-DIQ:P=26A#fAMc@&8U>G_Q0F=D
>:M-<^(&J411(37.H@^gL^=6/[IGYP<M9b4F_N.C]SY=cDaZ?X]R0\8Rb?WK=f3D
<[(<9bS0c0__Nf94>9^C=WTV[fEM4=b,G/=]g3TK+2QQ=CgL2N&4d+d@&XH/06S>
JS0H\&=aZD8ZG^QJ6HN09PR??QKU/SW5MAfgG]GXZUC5(EDRe\/C76e4A.\ORTV(
PBPbUeUK/^+C:XXXT,YaG#M/>Na_(c5R\<]CQU=HaZF1WKEg?EE)T4W7Q>>0H^MX
=4[Q0TcUb:O_762FWJO,Va++\f:OAP8;;9P)2N.-E2U@g?g?O0?@9SW=Wgg^.G6E
A@Td6fa@.H2U&Q8PB6]f3J#=f?Lg)841K)_4\.:<HL?]c2XNK^f2IG19[G5ED_BZ
72bD4Z?_cPgJfYZRBL]C.&V+Z3:g^g0dWH6Z>K6O#I[,K0FTF,MTPO\1J?S-6Da+
^D^@RZ3VJ=N]W@=gDF>^?=V<I_.aPN;edW:6d@7-V6,,/\_R\\;gJ-Cd2TZ=9Z&)
S23A7Z<?)-,55&<a6KEW?,?A&L(-,g:6\d=5a5CKS?O/2LPd;YQT8XgQ9-^;#&3Y
Q/=H(Q,Xb=>4O2=,]_F9RPRFI>2WcB-(D^1ZUBC2?<8@80J@1\-P);ag14,18.0b
CHW9c[&RP\C1#]S_ROSYQ<1.(6#,f78YFW_L6+/^?aQLD3_>2f=7+c;QYH\\9SV(
3)91Q:KfV3A9BV,TSBQ7^-7D8ebA6#9QI+JW]<Z6CEC0MDH(\(EGgF@?QgFODO9[
F;XFBQRM^TYd)LbJF&)<3E>TS>\9V,3G=C#dLHRd8g5#;:W@_FP\X\[QQ(30VR;M
^@&,GJaJLcEf=)9AA;=\AK=B=f^G.&XFH^W8/A63Y.V?T>B7e<QVQ?,[=f?-D6JD
8\]a-Sd,1.XF66_PZHeKN>#I6>(9K.AC3TA:^+CB-QF+&0=&Z?bA(d95AUA<VN><
T0IbA&NBFbRgZP,]f4/^)g2#BD35Lc7/Z5gfODQQXP68[9;DY3>[g&Y1ZKWd^4TO
7F0Ec_(BPXG3C6ATg-6LBO;KQ4H9@D/+cg1JM1JafA:E/4=?=Yd^J;-3EX@[F7aU
J/O8([13/H>T^3d?a6</)b]OK>9[>Q:6T=TT;;R<#d68_8S?+PW,@cLP(S7428D1
6GZ8K5I/gS2C=\Y&+IDW9:L,5dFI,;EN/9ZV=>,>CJ?)9ROaAa+5\WL&O+L&EgXD
fX1=.MfH<I_/:5c=]#&4NgRf4]Ha<@HJg:<f_T9?6&I-+#AT5=#P?C]If;N6>bLa
@5<YE303M-O_+[2f,e<Jf8aY(I\]EEfV^[P]@Lf6c4f^J.,E=X2_NS+9_2fa]fMF
#BW0S.1VH+K(QOWQg_335S+YS\41OCbNH-4KUKM-QaI]F@=UeH26P81:7Bd\G\S8
/?^Md[UR@d)TCOBOe9S5b8bZbBN5V_F?-\ZR4)]gb<-c=-G;4V,-ae#De3QbKEU8
25+HF4[RHPf9742#c-H-8S<ZdR:bCc(V/:>#L[e9,KOBCI]V\\I5MC,4[?g]\5FE
VDf,M:/<XZB,.W#_Gc]SV3e,[TMf5JVJAM]gIgB6>bMSG,H/]2/dVTHZ\#-I@26#
R)S^Je84JP\G</^L\.a6=d]=&LD/7+R,?LfQ[FMaH_\0QdCd<DL,=J/_gAc85Q0a
4d:X:)/BT<ALD(AcMaE^5]-B)fZRQ9;g<+?D5&>ZdSS.RWMV-P0<BX&3K/;Q)X=I
K>#>9X(X2O/:Q6&^+B.VK+NcO-CM@dN/N;GXPP-1EPXQT]=L,=]c443Id0=df_QP
CVY[WZ.b[Y50A^@>R#-E2g-9ZZZ].-EgEUWPeR)fSP53:#a3c72=1\.>C)(MA/IY
?5ON-.cQ75bVKJE_<0+3I7TL4P[9A1CF&<PWUA\P#^>9A-?43aF?^FO\:A44),Y[
?]_V1D4dY9)2L)?+LDX:DYHdOfRZWO#I.,\[;]VQ/7d+agDTJ>Wc6\)_J(YH\EJR
#.@I;<0D=;fG<SE0TF(#G9fgZ0/[0dP_K4#:H<WY#=CK7^BC6FMJSRe(KM<efCJW
.\a.I2R(/9BSX+b#[U@a.:P4;)XfEcf[ALPFZfK_g=B2G+^@8>.b&[RHSD_)PN9B
M,IO&.?P\VI\.F_(YYV<0[daN7QV>SCIJ5\,9;V\Z;7M_1\V^[V(9UO,_e^I5Gd)
A]eE9cQKCe1/C+WO>U-[8EA>(LUWc90[X3Q^<MGVV2(=MX1g#YFcGc8+]\Z/Vb<(
?.N8J[S/1=S(fKJDdM53SKJT8Gb]NCD<c8YAa82NDYC..ZAKC)d:3\W9a>L6XUeK
<Y:Fe)E0]I)BX__E9dc<U#b8UX,NWe00<()TG7#J9MAD0c<b2S7\QA?&&.KLG)](
g1]b49\2&TDM367Z:EA#UcEZ(5E&-^/c#?1/1EZY.gUU65.OZdZ#WL5PQY2#B2YY
2;VdFGd]bR42RD:@VZ8QTFYT9I9Q?6Wa]IPXC[N<O<)T-V_YE6\JFZ[NA:3(O4ZC
R_HY4\2M(Z=2^=0cD[(V3#<N&1Nd]A>>C4.?6KI=51TYa]V7IVTfL2^Y:HG-f,3E
a)c+PLPOd&MQ3VADIDbAZc1D#)D#2Ya??>H>a9#R/c6G.U-KH5=2+g\>WVZ/MXU>
CQ(C--<M[--+SQ903HDM\V_P@MV.01c=9QFUHV=8#<K)IbEJ^/J<:+KW,O?7T[?H
?W?D.=1?aEG1246g@bE]c4K3F7CBR=KbZD3WKUZ0?RN+\.=eSNF=\B.7&]DLR(Rf
GD/b2QA:MVN,7R&[8JY,?^XP&5c(??GfNTJQ<-FFI>f#TZCg]UG7beCBX-237cF\
3,^J;Ya<B2/+SOR#?[USZdJbAd#[JZ:A8)R1(.e@G))b?<YZP?K?A1@3./;bN^[\
#eF0gC[A>PO>Pd+X?<]5;QbS:M<2A48WO[HMV]F6ZO_Lc4cL87[A3)R^2)ZF4<:;
)R3f=X#4:_d9gESZ@f[;JZ#:g?;7a\E)Y-R+[MIVYI2VWWc^J/]]C?RcZ?<U)_^3
+9M6D.fc=dE-KCfG?.b/Hg]BJGab0dQgSg;Q3f-F,.eYcSPReP8G,bJ#IAP>TBL9
#T[/\22J)KbY)(;aOY,aX4<@NKPCf>WWg3HDd1E@_]4EfL^Xe5);GNaVLSQ8MHB]
;PR:ZGJR2#VV/MW]K[E9:#2HGg9785G&]1-I(fUH0(D6TZ5X.>XeK?PLb#Nf#6L@
<7JTHe;EMFcEcKLKg4J@,9f4D3#ZF(=e(c5H=C7U9L)&PJMQ&[GMeU(Q,bDfT#a:
<,#CEN/#gB4BQUM1,G9LPbUUL_4.(I,K#>,/^_HE:5MJ.P;?2UNV,2fF2BL,Z<5O
6?TE(8:e1e:WNY&LK-ge&bP3Ke9V4JHY^LWJC@/.NS[T#0@DRNP#K/3IBXXAM,a;
@-;LL+bPTF?b(8KB1Y(G<8AWdRQ9N+<QV)E1;BO50@2T4b&;1+_NKW0/-^1TMSO]
KU^Rc2/I]=V^aNSAH7-3WTU9):b[2UY^#R#f.#\]-8SWc4);UD]B1HMLA[33bge,
6_@O4NM3RS^@e<DX6Ca;@UT)2-AZKO8-W+3+0I#;e]-MF1/2ZD,A1^P]aFWBU9J(
96AG[&-:J7)9?H?G](8&-H86QV13RR0a99=K@_P4Cf#U39BOM(TaGMX(^M34Z.BJ
Z3/;CUc5gP.R[fgKWgVO1OKE;OE[KO.8b?g36616Y6>ATJ5\KN(Q+LHNN2>@Tc/:
+:RPBdb&DYZW+-OO^EFN8:@92/Zb8O-2=]-#2+.FfM)8@@@Z)JCBRdBa-M,VKV#_
E#f?b=/fNDS+UM[8M=g\70\1V=SdK@-H3@]5M7:\__Z;\b<g[YCI?f>L&WWE6VD9
72.01?\VF=0M&0TIcee#+/[8TTKTJPDa/Og0N9KWJ\LR^9TF(>(BcJ_M\BdL@b=)
aETYaL#S4QJ+Qc^;U65.A3b2RC09#J0&S+KR,\EYMM#fS5d\dcD=#c,7Ng,U_E^,
9aS4MU[;VF.[G2X=cIC/-LHHSCX31<O5afeVJ_EZ&B15fH\L\?=gg1efLV&KY>UI
b/714(b:=@8gf3))P4VY1He@NK@O>gH.LWN.-V+FH=R9V6cNadO?DQ+G\7YRe+L8
gM(d&ZCa;B[-[3P&]:H.+(@\Qf,BU6c^.b06G?B7S76OG?E,@IVc&a\M<<68e<a<
M,<61AQ:C:JdGcNd^3Z-?BAXQ<7fg8_7HD>dM7TANZe^&7IB/#+=4Y8E8/7Sa-cP
?f&Q5M)U)RT;78336.E_3?bNbW\-@7g3FcB)K>UH=CD2\MGQPWd:]IJ>4RbP0^##
cSafWY+O]c_0cK+A.9G>L6:_5R4M=b#7=AF.eGeZ8V?IcgTc/9QT#B<?Ze+RQFYX
?KRB^YU0f<e#JK3^d>:,=\PR9-Ra:g\Dg#(?/_[+M#;I++MYU8GWLU]Qfadg\EAb
<&&T:@\4SX]<GfV:<Z].2eF?2:O2-=T_8NN._@c9,S&GC:7NZ7cb&OYW]65+GV62
]<QQMD#K5D(aSaBT\<B[_/_4(SNQd0D0c(=NHBGde:O8,&/A5+A@T67(7VJW[<dD
=]9K7B8/V4H#WL8)X5S?)NM.>6@D)cf_5^+/<AJLIU)GCWWYeJ&G_4Vb,&,\XDV>
)B3d\O7&Df-5=7D54/T+/aEH.L-.MIA:>EHDa<AMDPDcW5F-.Q0?c?OQ:<gc.LMa
>a4IG7)RM@0EeH#M=TTN7O59ET9/L:RC08a@gUW+(S^N&P\I.@&\LQ,d8RBKBMFP
VPL=S+.;eFQO;#?^77T(Wg1=<egVRY\(\OTULQ^gWQ4M_W>U2M3\@+^FYf7Y@DYV
>P&L]Ica&Vb:LZ<OK&:VYNAW;BeY,2:_L0N8AQ+5PC(>U5FgZX2R83>AVL5H&+[:
-4a)DUaeUXSPVU:J8[D:5\:0O;&8<CR8dHN-/ZBT>RXDD],CJ=A6<@YMD>63@Kd?
99UB\JAC7>9bg(LfEcJ][AH:eSK+)66R,(A3@BEY++:\dM6][1,_I@JBD[G_FKV8
R8?4&N)c^K-CT(VWQ/+__eLUB/XafD)XAB50SQdMP)\PB&1;&>ZeUD13/\\E<C_W
Od(.d3CY5O9bbL#I+(;^]^c)LY-7A3U-J>Z(C/0^OaH10IK#1d.0.a\)5+^,<6QR
]2/4X:,98?.3Y[9)X+AN#:/1XV>MXgRDYZL?G:d)8<Mc:5N38P\;#,fXE_W=HU]@
Y,4Dg2^5Z@2BHW5)L:2;3gLU1aZGVR(JgQNcOXJAD>?[U^1e_;G8(>^)HFQ5HOdF
2I.GQ\24KI4/HY752=AS,8HgOIJ+,e6J][<#PcE3Z.e0L\(T1FXV;/MM)LD>ePGg
VL+JC32GNSPJ@+-:\)65<C3()DG5Q3YMD;@b0M\gfc.JA]>D#YaG)N>]NW:;>RW&
GYI/b#e>b?=()PTbA8]Bgf:W\7[T.=?&D=GSM#bOaBWPH82_ODW&9[-0B#e]g\a4
?4,J#@;=HFeC@VAGTQ:GH4U+[([EWKL#.-0+P&D=9gVF.[1a[Q9&Za]7dbG[>#Mg
c.L7A>Jg1017gL,&U;eBBZ)8#eEa]EBJ:XZ:9Jg7@b:4VJ&G7;3YBR&fe]/+;&+D
=a>_1ZWPUS_[@,R.?A-OfIO?ScFA.]2?</0(TWf?PKF>Y)b(g4KS=ET;(5N[IKRd
;>FDW:.GIW6dTQ:TKD948]W,\(a4:gT/K]N+L.B8HZD-g2^+WfO+SU07D7YUXF=&
)]Q+QI5UAVK9/X<NePdQ;V0_V2?[<L#e^/W(#?LQR&V^?X5WaVUb@0ZG7X#3;=R^
AP#@(c[RB41U8G)7]7eD)fRYN3a78FDYVURB2B6QU:aPVIQY4HJfFQP/La4=HV+d
7-VQ?S?@BKBfVTZ/ac+)LEL9dMQbP@F\9adPW_QKG@\c5G8B)Of)C.dIZ4ONVRFH
9?;@@OZN,BK#KZR_=-FAM#<1UWOY-F_7Z?P4\[,596C92PT#?()ZAS+]:CHe;#61
=Q5Gag\bWOP#-&[g^=@3g6#S=/+J;a:e/c_Abge?-V8fLGA4GDfM8C1.XJM2LLLX
^-3D5cWB0@@[C;Df((7>G39\G@2VNE0(._S]34@3D/Yb/7I)>6QJV8F\+bZ.H6.Y
J9-687ZYUS5FO1P58Cg.)QHDI]G3]&Y)TS5gLTK(5f=6&J>15d<^@&>XXfQ-)S-V
L6&6+U_TRSb>>Q^cDbQ/dK=fJ/e/g3AC;.Z?6]WZbN9Gc@8=T[/Ca]Ff6R99J+&8
EB)T<^L\,&QeQg-0-JG032BX^R^\Q476_H0VLWN31FXQPLXXAO^U_3\+<#>eT2VU
241D/a==LgZKB.WM2\c3MRRINb>#O?Ye9.<=aR)4(9MRW)9MWDHQ]0fA,:fF=,IA
4=WZ]HJ50H#K,&1D(g0<Ea\U.@9QDbE=H^B-2BZTE/__aABPG?J;HFG&C387C2=8
YU9][&Q#7aXBCEK6+eL(e?//.)X::6NIGNZ4[<fP4d.QE[M/)8N^T9,K+TINReWD
G(IUgdDQ\](=4cIYHXc4@G\M2[O<_f+>(gN-;P.[OZ);KYf<QT]UOJ7\L<b?0bMP
VHZ91V;f6V_17]BRK+D,)&==>.A.4(W<^E^d+gDXDNcC_Q(I919.eSJPRg2W<([e
_4cFd?4bY&-SW0BT;QfD=08<-F9K3;^JSF1CXXC6Dg-ALgP?E7_fWST\D_(CT_gR
:O<Y6Z=R/-N/OSZ9F@\&&NdG63#57/^(FCW/c/SK2E:OZZO73R1-&69YLRONCTV/
L>;R^UfOGd7eX?YDJg8dAa-NS9OB4MN:E3KSO5]/7e+c2CJ<RNBfg_9@)4YBYAWg
A1KN()YQ#W=\ZTXB5EAC[1CN[&3FYRd4-@cJ.)R+8gg9O3OII\[_8B:#.?c9_72<
Md,11?f7:bc9X5ZD,.CDbe@H4UYYa\cYX[a9>549Af5R_g4Z&e-G0aTbD8:MR@F3
R1O^/-X+M;YAK8NVK2c-<(KMZ;5CQXQPF:Y?fgfF=5P13Q\8D.#5NFLFg3GEM0=e
-+[J(K&G7D,UE;&VQ+NJ;N@EOH]dd2BKBV@AGMPGaMDg[.&W?<,WU80M7I7KV38[
O>_fLC<;NOHDSTNSBKd_D6L;B[L]A1Nb#MF44:L>>Q.cB\5B6TZ1E:,f3=C-^T1V
9OB[([5SQ(S19T+&IOHH)I;e[U:G4fa1U/\PKLH:):Rd4E&4]=O^GRHE]EfW>dcF
F7WYQ7WF2W1PEe,9f;-CX5;XWNAOPO0\(XS[9_)OQOdJfQ&/6W+SE+@2H/MPM?f+
H[,.=d.e0g#)JUSFC<Vb8dV<_?fdMJ^Qc>&,+<8Q/2QC</T\3:L;&>.2V)HAZIO]
c]YO0WGFZ5;9FF&?cBeL6R;)SN2RU0gHF8+1K4)PGR#U/ZHM4V4LO:4G1a]F>4eC
&[)<&T_/U=d26&Y]\102@&eGL?,@1_30]D30F?(92\Ug:&7Zg+(LE@<]8OTH1]A&
S5]ROZ5DK[DV(T,>=_,X_a?/+)6&R9Sf-HIZ.ab>>KZ,8I77K@.PgSVKORQK)=B/
^5TT0_G/UXOR?DNWFfe9FQ4G,#c,:]7LJKXPRgUQ3D)I).da-4GXaZ5fWM5)]dIb
(C2ENZ#P8>:9C;5;g@5I=?JLS]?2c[:U&c)G9](1<=9)(33EHF^\c2QaFDZ7_DH8
@42GeNE+K3f9IH5XS1KU42gZ8=GQHSbaZe[?PX;4;cC9]eT?XcMVLPZLK_6#FZV#
XI?=4-?^H[R9:MKUFFX+bWCHMY?,\Q]5X&8H@<3SKPg/0JaC>:U7dK+b0DO:Bcg<
^J0BL0MGg-E@.\F.gOPdSP(]K.Z&<PVdDd.UIfb;MfU2C#gJ4.R@@=TK_,XU?&&a
PaTZV5K0NW4,_\L330eIES[8C=0<aW7YTaOS3/7Cc.?;S2(W-^2H;(C_F2cI[-Cg
AZ4P0/&.Y+78L6-:G(ZLEO/_O-WI&-J3G8eg=Z2dUGW1;G5@;]CAGB:C<JT(V__G
^WbQSWG_FJ[+9(CQU9e#X_P[B:e\QM32\#bO\\SUL7P>A(&#Q>;U#;[_W_,0[?cV
[b?,9\X=0Y)C8&XGK(HVB//[96V?U\=d/?^J(CI9GK/B5g.JU4AVf-LK6YJ4C.]]
e=FE8MJWHDNH0LOA.L,+Q>26PU0(WPW>.Q)/@Q@GB6)7\19]Rb@=H\7K1DVG]^A^
3(,#a)THJR4LR.G^6(IL3SQ=>)T;-^3&G7Gf^aWDXK4DD,448b1R1cAZ)\1??]#2
<Fg9JUR_7dXCU0^-5XAG]9U.bKU6^3Xf+);]5NQN,TB?fA3I]?KG5cT,6T^OF[Me
^K1LcI#R:gI_g3V:NJ:XVVSHg=KR59;7=&,QTPOC0[L\#)AF17C<@g9e^bNC(g2;
^W[W@#2.ZF9V3DMJ[A,WEJc6ecAD_<d=&DU;0<ZGPMCa54W:HJCY0\E8IV2Z4O:D
7-Ud8f;WN0Y59H1^>TB:c=[DWST\\\I(,:ON+&DE>ObC#/\D1,+>,0),d7@(I0QR
4e#H]7deJD-_[[b&B_95.,dM^S(UZYINNT-MS5)SSZ>Z14&OUV5Og7EA@AF8P;+7
P0Y0R7c7TGV^\48Y(gYP<U@[;@GGK#NDLYRSYVK2#6_Le5>6aHK)=^#K9<2AKT61
;Zg4=KP-cf\4H@.<Uf>=Y4<@7L#_W(3W&d6N599f,85;)0>.M9<9)FK5&&6L,?/]
;MP4###Zcb-Q<GA.K.YbED1LXeYB()ZE>Zg9&:S.1YDKL;RGDFI5U.>MUO4U^UE2
^[[b4;aH^IWZYg>/8R1(2:63221<CYV5TI.P)_HA@c]UOXN>-S7LQOP;NBRS,SDW
68K/:#d1:b&=^Sd=3C0ZTGDB-RX^>OT^NH2cd#3#NS\T]BJFQKE=S.LVVEaG[fU@
A>FBB5#J?@>M;Vge(89c\;81ZXT@LFHb16EZ?^J1a;W-<O/?L:\]^L//[;2Je>AA
EAfE00ce^92)eV?(3UgA9#-GX-TG5(H_e@?N4@7HX<DY-[S#\9_d+]:J>DQ&7Ff1
L,3H@Obf1GQ8NK:)>5U@9^K.V1.,-eaA.&N?QO9+D4&NZ<WW+7EO=IRM,AK^N;Ae
:>_=_g)]/L2;(J3#>DOI>cS\6R,Y^=[XKTNg36_P9->T(R(?3B0&]eLMG2f>_038
O^/=_g]&LaZFC9SR=2]Ca;cc;>[/6-/H-)RA0dOFU&d0K5Gb4T5G;8ICO@&3VP72
I:^(A,-abR=D&4.EI)LO/@&1]]Zb9X?Nb)SQF=L<[cTWAZ:0:f=<0+dcOB8YZ^A=
f.D#[cWaMJA1g,1YD@;?#.KHHJdZ:5=bZeG;\,B;&^XbBUW?HI),Y,3KE^#(9/b>
CI5=gUIFfGd+VgOd[-IaP:c^3+XQ,>bMb0gE915Z)M[0eDTFDMJ<#c_[@RD3?SaR
?B/R@9)8V0YB2KdV).S3H[?8OL&M_]3W\GV,L39=\HLMJMI,fGEb7[KCC<J@OEK@
YG14)^OO=C_+IT+MQ\>T[I79(/7XeBQQR2#&e,WdaN+L/.8ER0>WA_3DYV?&ZMIQ
?cZ5VPN]N2UFA3d(8Ia1R[N3fY+H8#,EbKEKA?WPJ8]>/5)_<f]9YFF19I.?,<)J
8-IKG5DC;C3+NF8\3&W])L=5;T3Pc<?Yf>0ZR-P@8,McWR\McND^6b@H8T;N.bA_
O<P;A9ee@K9L]d2BTLR.#B2.e^HB-<EKN^OZgg\M3g-1gP12f7d@E85R_@9[E-d(
Negb],/D1H>&fA._>Zgc:XZE)M3GPX,f(AZ2353\O,HL-P3?&L_E5=?0C3_[,Id.
M2(_(E.WZFQ>c-9d&:]?,NE&Q8=6f1\7@1=P1c^M2+X9/^OH-?LZ)4U<E-@NNPfc
TeWaYS=R0BOB2+F@W77P<QZdf@Q?SJ8a=.D3PAO1OZ=6(8EPD+Z7?,QbY)2>?R.)
;1A&P#LX[[A6C<0\N,K0.GPO@Z;Lf-MB&2S?@];R@A-N;F^\VC9?FSSJ8M4V+?35
/#XBKa;)PQ(daDe@9@d^.+9&[E4ZZ>D\G)=]QdRgV^:F-Ig^UCT7YB:@P&LKf)D2
5;&[IKBWc@4[U<C\Qa/.Kfbe@UY9,E8P(cL@EDVCOYB)>&IW[^D70)84dII58(#d
.OV4OR+e@)(#b(-Y>\2f-GgV2ZJ<7#46:NO63W>UPWeK\5=)V+2Fda;A-9SI,33&
PNO?W;_5D_Z0Xg-7?-LQ^(GS:@=Q?OX/dES,8A7A&EPKQ3?BP(FWSQ<OU[-U6PaE
JY1[-)T3X5MD1@#@;:+?877[<0eU,@?K>R=AB3J)D]Y[fRJ(=,egaX1XXJVO=8DH
V(<,ZN(S+Ed,6293>37]SOcZ.RU\SgA<@Q8gF>XTB>cS08&e.IW329L>@dXc+&eI
IZ>d:X->96<8SeP9-/U6X)1L?#I#R>KH6<JK/^)BB4PTb8OSXFO?/3X6#7REI&^&
Sc:>VdQ@Y,L7[T@P/FAO4#0M[^7Q+U&:@K>T_>;Uca0cA0)-CUH610;JQ:3[Y2^8
Zg?AUX<;8AfPV[I:#9D<C3f<EM&b>+QTWMe5W)S?.G)Sd+fN/]2J1PQ\V>FF#F,C
/U(:TQTW#F]3_<>CJ(+C(PCdE5?\^#R=^0(TDEEbT&Dd=bHG::^H@7@.JLM#E3Yc
[9HA/O281+B=0ZY8.f2;f83^\V0+EV;::LK/N#]eQW[BO/-K/Q1OS]dB_8O93cHC
^R4JEU,71X)bF;+K#48.e>])6ZfI#OaLW5ETH^1F?,bZC5.16SH+-RebE:C?1AA.
MH\^b1+_Z@^8N&?(/,0=NZG)QTJ?68A2;_eOA\?@4R1H3K0>-2feI_7)g8(-1H;O
DPE[)?KBe\A(#:f@WA^;aIAa,<#NR:/1,gRf]-IKK(9Q&^c4JedEPZdK_@,Z(:fS
(5G;4(,.MRdNLYYYP@g1^6?F8V6XAcUY\N-J-,M0JTRPI?<)2Lf^F.KfgMPS+8.<
+gDRee+_]-QKR,RT>/M2ACO3@eTF6]Z\O\^YJH8\=,T[6fg;I7F-4IHT@[?E1Yc_
d\OVS[<4<TO_g/=_K&E/HUJ=TQD>Ig]>2U/;J8.K>096@0HQK6Fg?.7_,6]6TPMB
(X\9afWa8]5E.a+7;S-bE#&HfRFe0#bQ-Q=G(DXd5_OXDPS^(CIeH_XT47M.,ZFd
?;-JCb#M4:=VKNH6J5fg811]PRcK7^8?2E2[--@Z1BN[4N^4K3d]B3\:U6OINRKf
dMc4?NXe;74NJPO@P84:JAZ-A])>FSYB?.,KI:2C9[<J@R^Rd:P.#/Y@.9P>&ccL
S&Ob/9/3EBU-B^f22D;OM>EQ\&[X(ILeNAe=)J(5cb[5:L]VeK/BKW>8cR#cOE#+
FJ8N21JK(^)BK^^WA:^IdVREG,eV,(:Nb5b;R_a38UAa5R2gD<?feP?Ec7>c\;g^
\:0OTWb>TX,cGUDE[8;T/cVCgS^@;/LR:/Me88Ae3X[MY#MC:=(WaQX1eJEfQDL_
4UPF-NAZfDeW^;_TU<3+I=4RI3@K:_\(KDgRf]^a>>&MLZ/[0Lb,4FZb5^X59eAX
+5NN:WWFd-A5bUeM->CJ=2QRB9CK0WA8CVNbcTROAV^Te&KZ7X29[M]g>&O1fV]U
6[8BHR-]VKF&TS>+/0#21_0G;TIIZ(#4=3MS4aNb<(Ve>=6XPb7D@)E+,7D(5>1d
M85.)4IIAKXa)WRMLY<E5GF[UZg2N2UX+,?E4MR41M)SENJ?,,VM@S6d6@UM5B6G
N_<7WA=#=)CU@b.:/1[:A=/1B-&5[<.5X9d_LTVK/VXO_bFa2_>g:ZB_\Gb+CbUT
d_fXUZc0gLI@>K7SZ0eK38>NJK(+N<?[R#KQXf4)7>\Q;_MQ)FDd[RQMX7R02M(<
B;_RKH:<D^60g:2?c/E;4G.Uc,[)H]]_e3U#)QX,\bD4,[LQ3)A,Ab\eK?gDTLFN
.S7#(693ZMf7QIKY9#3=^/&_b^F8;+1DQcYWdR(+e0b#[U1EN921FXHC;[cWHdTB
/V6EaXgaK;37g(E/?[T7XQJV9+A6Ea\M##,,22#@:f[T=>0+ZM7=KJR8fH73+5K@
PY5YTJQFOTA3DFaWJ5M,=6>Z9&.b)\UN)a+2>R0+RRH0^A_@5bIa7WWD6^Q]2B?^
8HKXZ(,,+[@E+TW8E&6HQR9RBe82_30?Z0\#1U&G80;.=YCF51\SdMZ4>9[Qg2,V
PQ(fJI0P;Q,_U8XX4?)68XWF?gL<[SK]ZU]87g_\#G7AZ.(8HV(&GV67P^_.@MVV
5f3++/Z4BWU9NOD[XVCL2g>V\[EZELB231X6KBU4+NVK1;D#(T>TD.N3444P7-Mg
I-HU#(FMI:>2aJ=?U;7D.6NW)DC:7[DAK]EVbbSW=H=OLP6IQYeOU9fF2\YH?.bU
]Z\gJ7X</eY-^eC,FfX>\]1N;8]e7OMS#g)ggUV:a^^Fd6_d:CZg;_7EHKaFdA(]
1_\0Le.Wc_&1K;6K1CO\=RB6L4c3EbA/)Ra<cS1.S^Pc+0IR9d2fc53RKgQL]fVV
K8-AbH_(Ac;H\fd;;8fE[f97:[R-=5P@Q0G:,&1\E(E>KFW/VY.PR/^F4+YNHJ>G
#MCfXUAZ1SL/WABGPI,<:F@8@[&CLGOCN.d\^5#[/7[O8JU=CXf6L-TM_^XSB7[O
HNTVOW5cHVZ87&b)-98>U+cUfN]_SCZc;]TK@=EDEM?41[d@ba\Y\2;7M&/?RIRD
OP\]-C81<;e(NEg+0P(,:[f8@cIaKRDK&;6gIYTff.a;I>LQR#a;-QHL/3>NOdAG
V3@YR;WX&S3R+Zgf[+aV2JQ^JLR;Z9\S+Q,K[GVgJD(4916]+)bO:d&LANA.5EL<
c8Y)-69&WXJgQ6X&XP:c0d#e6QA/4326R#/6(EgHVU.BeX2+LDTeAH()>1@X4+X8
RbBJQX[K;>L8^e\+L/]T396c./5-ZY_(+P_1@cJ[Rb>,&W2OM^\g#-N<(70>D(-D
\+\DCLcY^,4=-/CPF7Fe9PQIY?F7cTNO-KccQKY+[_Q?1g(9.1T#9IF/LV;G6-O&
XRXJ>R\T7@_X>I^++X=KE4TK?c,eN[TR@(M#]RB]d>3TT=DC6Nad:R8FNU]0<F#U
THK7\DE)&RIUZB511=)Y1<7EH.Z^H#D/g&8LY22dPW)<^-<R]2@<<^gZ+KH^V#R/
SAKAF@##[gLbfB<RG8g(7c:@7gUP.A2(/UR:gTM6;FbZMI,#I20KIeGP6Lb^Q4(U
F1+799:SgV^gA@E3IF69/SP2RZb\/W</B[d1KV:LfaH8A4>I-X\-eNb^Oa/7<&B_
+(dU:T5@6-2V&C=DL+?@&<LFIUQ0LcH-@BIGQ#RR;3Z&6a)L<[O6gfS[3IR#f18^
Q/./_1>^<YWNO-4YN_aXJRUIg/\CDe5G;+PU88eKX]W5Pg7dQTRdMHe(2##-Y#B2
UaX)N6^\ND-O&FMMVcWKFc(WB5IIWI]FH47G/,T^D9.=?>2^1,)0I&fSLB7NLUG:
6-ON24;2VNOFR1<#/24&32-YW>\:,92IcVA1U8XMKL<YMNZ8<5(Y@7\9dMP9M.\;
fLDFKNaLO03?\JB1E,3@abC-5E^9S;J-A+R=JY_gNSgdNGA)TO@N3R;?b]AC.K&a
)MeE=_+=e-6dG8BcZ@IIe7\S_8#8205/(_d:;E+SN+_DSd:\17FHe<g>Ec;2X/FY
:cPTB2f?L6ZVM7#)5(>ID\LcQ)5eNCAD8+MOg-Qa/RJSfF^eN=+8VeKbb9P_;MT.
_[0X6&+GBI8g5Y,?-ZYGJX]EH]YD0eXM;F.J.1JUK[L=03U?ATXcVZ.K1;8+;Md]
,g58H7VA6D[8b2F#E>9HH,&Ie3&V4M?RLG-0GIPAT-?W2KSa@Q:XSNf=VL18MH7b
S,W4+]._5_H)JHT(,&24=K2TA^K<(K0a?>SCHcZcBUSZBF\X\FR#^DB?IN.[N+BK
:4faTX)NNKe<cg.T4@6./39B8GWW&Icg^V[D]T(U=F;f<R#EN(;bB,:OZ#f;^Nd3
L&NYd]OLASQ7.6C]V4<]XEX/D_)W(@A5DIL2</HAA\25S(,L+W4)G^Y3H1@^;OE:
HHZ4SR,6_:3YQg9C?3LP)PdbNY+\4,eI#E)3d@_+Ice6^KNY]CB.f<;D4/FHUY=c
N\05I=+N3=94-#O]#;+-aUL5Y\:\G_LH?QWSaD6aW8@5DeA>b+F257Oe?#aV].bY
fKRI.0S<He/#H;:Qe<3HW-;QK;+2I]61fd9)=8a0K+NGGECBO,4<<B;fNc</bR.<
][a)98ZH_9>K-R03&,VB^8,6_O;fFU6g::=&bRgG#BHRLXMQQf@?4I/FAH7&+C1P
^cOYDM@Pg6a&VeX@Q>R?[b\W:U^S_G6&<K&X=Q&#;Y^#^U^a>29&ZEA^),0^aALf
>3KV>B-RBa&@2G11c^ITf#,DJ>3]+]\g]7AT@Kb7VdT;.0JP?de+[CR_UfCS^24-
0f50W=:Z:fc@_[;c1_89P8,4GeS]@^=1QdB,(dg;Y2^)&_]8SaBOL6E,c@TFQPc:
Yf5];QMV<ICS>GFG5X(O,J)e.X9gNbCd\ILC,gC\KE.P7M1(TE;OO,X#?a^8]E9^
H185V1f@\8M\\2,KFe(@FG]d<+-7;@L]];ge:a;K_N@;?O=\MggT4fQ3L0#1b09:
Q80:Gd#e?^IT\1egEcF5C3TN2156gaNb]0-D(eY1cAc=)W-YI/DbP[HcLR1R(BF8
N4J=:(]<2(IB&EeWcPdE5S]6F-C@#-VJ)J>3@P/Z\-)?WL9W@C?I=0X)-bAMKRSB
69,_3[.:7NI3Od+M7^C[,,,I5[MS_84U>fd,L)aO49JOcAWf3UC/(N.:CQ?X3cII
-38>A(ZeDTNN^SA8:Ygbf;6X\gJ_-[I:-(\+0_]\^?](@_H/\OUIe-0S9Mg:-FO#
:]64D,P>CScNIcfa9.VD\8G,FN2)AcW0K?CP@Q]OR,PTG9,SPf74RJd3HP+&4<8+
2#[IEDUWD,7=.#RQ5dO5//FR@,dKAC\e6bNAJ--CODP/^9>6T.IaY/4+9.A[I@NI
?UG5f<f:[-+[V29_<_)I7<N>U.4ST(b4BCVUI@F?6;Z-V(J7L.PYY)(,LY0d6QJ/
:E-_ZOfgAbPgT1<MF?93W0U,&5b03b,g[W)cT:A)V.?3C+,33V)3^HTbPG+(FLOJ
&[ZXI6/\MI8PJ,ABZE&,MWa^)_C;04_9D;-,ZY=Y9KXLM(NYCC;R)^+C^KBf?6U9
/[GS&V4B?ObTK^=\bcS[+fLPZS&&EU+4UC/6CYX<-EYF9c.U&L+VGLM:AQf4757G
f+f_&]M9U:RaOW?D.d-A]eS^)1D7gDI:.1eg<Vg(QbCQ<Q24[@KCJ)d8g,C+2DLb
92DGU<&Wd:c?:gC]_+(77,,]XI778TaKQ;VZ@Q>XB<0SSQD@S3K-d\VS@^7J2G?/
+^c1g.33[U=:ZH\a9a,fH=@@\4DSURJPXAdfe,CCbQXcCI?eEZaH9CIY;W;7F&J&
(?6@G^G4N[0dC2FcJN8^P((-O#1R[I)b.)LO-Y_aIH#&\=H9e;d,[#&/GAVQC3cI
Y[gW;SJN>bYXW3+4f<>MDGfLV1TXCC(F.c@5d9.&GS<N<W0IR+bdB.X>/ZEf=NIU
6;[3_6RfQ8[H[b/U6@Fd5F;EM_6+UVU8DY#ZVY8<4:>,C?\_C?Se>O7#]dOP,Q.#
T5PGZ&_^;gH,3a_E6ZIFPGd:M+/]8)eH46X7)(9N/DQXgKW[SaDNdL<SW]N>E_;;
?\1,JP4/Ub/0Gd/BV#BI=Sc8G2XHD[.AZV)D]2D)4O(a]fZ;:We?Q-Yg<2B9bVT&
UfZg,^<g>LFLXR9YT6_W:<>]T(CebWE-JY3W-2F(MI,5MVXd^)&JZbM6)QY#,C1O
0OV4X#[Tc\bI2]7TIF@/.BK:LB1=>8N02cUfQRUb]G7KP@Z&_#F;ZR<_#+J+NH-B
DFN6O>ER8YSBTSXXB[L=)N]#cBaUET1]=H>6/?7A8S@;LO.U[3Fc>#>K9M(H(f5;
6bb;TQ4IQWcT#I?<a#93I0Z=EW[8H>+=L,V,3eaEKB2_#>W58eOXFK,\00XZCO[6
/N_FNaDV7\9be))I/dYHOKdQVMA]9.@:ODJW@/_ZYCU-PM6+975>NK^M<5SObCO;
Gg(X-)O9\>.9C0VKO-=f,-P_G2dY=W&BWHSfAZ>6NR5?#WIYfT4ba8B:J</&S]3P
a#_GTBVGbB8gKf7P.DS@TH#H&XZ5]1XRUAV46#f<AEHWfE=]a6\/5:(dGB@UMDTK
YX^Ic2]5M)+dST0[I[Y1)THecc>^/;=dDZL[,fc7^@_5[>L:ZQ==D]QK^Z&,G+G7
L3,^;/V)bJIWXR+Ud/KUB(\Cf1\GN25)Pb&VA1e,1#4gV/[AC=;\@F:8@ZgW3X2,
.1_VD#9\6cf3@aB]2M<0[_f84^O[f;=e:ga<P&X_PIg_SP58)\Wg(E[QIEYWYSLI
&<9-^e\a9R-cV)fXVFTf(F><PB.:2f5/5P=UB-)Q3V9G[a(TR+B4QI+e[>KQ=@07
Z\c<XBa0K[c_5_UR0bdE;ReN8.4GdXB^g]T2H,SE?Vg7(4FL025T#bMEedA<1E&c
cICafUYg./GKEA/D4AR0g[8QgGKdC8>=3WKAL3)b5cO/e[D0M^cIOK[APJCAbDY\
e,@,,IQK7cf)U5M7>?<+gGU\=<O,6cGK(PY.-6^:d[]O^85[\&ZgX2,L2#Xa0&>]
e2c0=8EON.\HMcUY;)?UL965L&LTD8]F7O50?aQg(A<T,SVO+D#BB5A(LCTG&7&_
Yf+[1YBJ92WEI^M.+UW4D>.+J^YFW\3,JfOB3)#DGfZQT>C5,^DN+-(f;<aaec6W
2Y<G:6Z?J#3cG48gF3UKB6-U[O4I4,6LL^cb:)HX5&DU.2BE<Pd32^:WVQ]C#<>0
(DGI=RPROVd+<JW?VWZK7SEU2=?OR/+HWK>T2#XF?7F-I;^/#af8>5E2Y3JCBbLF
U6=cd\\R?bb-@De^;<-gbD12X9\fbMUXK#EG<(Y&_AFe2G(>N7ZY#&^K]+X]+b.K
ZKFcb>/MBB,03OebHReSX=5Uf]?+:]=8G-VdC3a&gd6ZBBeNXXcf0DT_KXI.]LOg
38N.VWY[dT50WNN9g+CE1(VXVIPf?G6D./]XH^PJ.TDNC;V:OPQ>d1&e\+-<SPB8
_#5d.eAYP@+WOSP7N[[ba#2&=.W=K-\DH=:aW@MVRH5-M7ZedGV:(AedD13&R7>,
>YA)JA95GYU9\,bXb6Uf6WB_5c7S[a/1b:(+EV_BEUU[QR_5[bM1Jb_#4P6<;7a:
KQ[6b4@]=))Ra@IU#<:e=K#/N;PE:8>X\[3da9Z>6Fa7:V/5T9;,/J=gYa(4S:5P
d^4_L2I^+ZMR<N=bK=6/OJ_)Y^IL.M@C)OYI6FJ_Sg/c8,4J)Vf@c.BHL?,5(_LT
33df.Y^D@ZE89Rc:geD1_;T[U.-+KP^cUJD2Y:.U6>Xd)9<CO5N8_c#\?\a1N.&O
[D6,48Q6:L#M.QdfC;Ac@d/=K;YOTF0QHb2GR-^,E^g4,FSAfTB>+)89QMf[IW?J
_RH#,V[bY-2L,YWH_-AD(cd<Xa;)=H@cF<PaCGWfHf;7:YSf>Ea,Z\FP6G&<cZ_+
>[-CQ31OPRg:gAbdVFHZ[;AaJcMX&QSI.-I;SZW@MN#:L\13X#]-[\FDOZ&Gg5UY
UZ]^B&)ZR>QL:T65Dc[SeS2N-0gd22dU@.57SP\3,:?eB+g+7@4:AGW1Re#>E>70
^+U5S.OfE;7ZKfN:bY9E0:&^:?9^ALJ0bRR5T5&a638cSN/2O+.ZbcQ6OGSUO=(0
2T^c/CA?^(eRbNbdO.1DgH#(D\Q;(F1g@SV=df(?15],_+S32Tf/\+)4bJ\E-/eC
]2WL[8Q8g/FM1M,ceU6DQK&Y:[RDbJb#8aZEG>aPBLMT>\e;^YL&P2cN?FVJdXdJ
>TWcY\d@gcG_0O\BRF/YDWA#X7E3+NSd?8V^<MUc2Y-Mdc-bA3\&^7Bb=6RX>f5(
__\fT[_Qa#T>?R?ZFCX&I@EfT^U9YbB&MgDPe]T[GR^e=A[7176-a9]3OTWe<?BW
d9E,;gLI0)=?+a^LYX9g)Y3\RJbLU:#F#BSRN2[_^K\gb_P-/C=O;J70W5/5#WcS
R\FDWF&bK78MXP\(P7#A,^?g/Ub+)c_]#g5fE+)<dV2<&C;8]@5DQ&c?>Y<fK6/f
69F<f-Xc#Y4c1V()(?WDYZP,&b;I2BE73M12FB=@TJ3U]K&HSe\A/-dIZE_e3=QQ
BJM8f0e2QF]??,70>RQ3_VKWd)XO9W6g2E7,HgRF\=VAB<3DQDXC#<?R1N2c)&)J
C#C:b@OK+8Q.@+8U\Q&\H\3Tb-B],WJacF?JQ^L.UbBRS+XE8+T4E=VOggJPN3K3
SCeF].,[gENP91REG0^+&+RfG/bfgI.-HL\c0_D<_V+U=6d<V62]gC3G>CUFDQD^
1D^L<[;D?WY4?Ufb19NV-/48/SQS_L\PgUVR)I@GXYMbc?N.[HZd#2QVPEK^_WZN
UCU:da1,ZV\Fc8T:&,5^X/35[gE0\cM:N_#Jeg,7gM:(gW]GJR7E@&-]+0YR[4^+
SLW(\be+d],IN.O[fE;1R#.5::-[RVaP3(84KDABcQRP[6b[KQR8P/Q]@Tf:RgR>
Y)GA+WE)FJN^b#M[IYEe3DL0O^6DN4aJ9H0R::.MG3DP#LMV?R2^JL5+Z3B/IKeR
B3+.@7R2)7^LA9FeJbKD;CUb2ge5g6&.Nf9e(A0=NAX@P6Y_aMH?.0WMGU?E]0,b
)ZJMDLSBX0XSN(g0B,8f0]:J-]bVCZ_8.O.SV0+ZNNbYQUUFKCdM2[0a[)10:/IS
VJFL.Z+e+Lg1TcD7GU):J<W_/0DX&3N#TM=BV8?>M<Gg)E0FR]SISA<5(-21>f(f
I3,16P;XS^_a>>G7TY8-<DGJ_\I:N=03\;0[],+R8bV&:b2eP&fG2d&E+2KaP,++
A@3)X0[.QIMRaM8CfR[OHc;bbc@:RTAU/DZ/Q:33eE7CTaM7e_KdIa>(ZI+<S344
b9X63Tf@=e<\&CJS/?Wc_H@B.V=EY=O;#5\MH5PQ.7EE#9+J#IK[&]E@[.HX]7O;
Q.6A]K01:3?<a+7eI,]EE,D[BSKJ5==J]W;BgS[#&J;M0_KPU&GagW.US@]:b(YW
JA&.agbQ_-Q28H6F41Ue=?_V>9QQcVfI&18fgD00e9W,^RCT6@]?6DL+43fA2^L^
C[5-67;gNeKC@9dH6_WMW>Z_ATQe?8GJ9])aO?L2]9FPe=WH+:+Ld0T6/;e6OPA1
cY#,W:FVOYaESGfMSK4W(Y<,dN5TN)dD>dXPb&-b8.]V\Z@&<(K#Y/_ZQC>XY,5(
4,YZdY[CgcB+=9_VY[W.<]]5=Dg8]@SAVV#MDYGJOD:^P<>gcHG]c7]^aG0,bDc@
eRB.dd4d67g07R;e_JI(F#@4Sg[D5&d\T[bR0]:FM_f83W4]:Z+CDQPVVBfK4ZO[
K5GB4KXRE+YE>8;CI?:0;TC?ag86]I:=YP6;O11Mf+<gaBG3eO?/G[]HG-Z2Na>N
cUf8^T5CL_WK=P9-0d&_PMH&Q<C6I\N3(Tc?/d)Yd?A/HI[LV)b6F6PX>S2eDL6S
#)0>N9dIRBg+(\EG9U^f^;)P-9R(HQ7X<MBT4P:9[]D_3RbGbH]]]G9-L\#gA0^W
/b>M^8&e0>LCU&)ED[R99&^/PFR,GRLYA<dZD0Q(c[5>(]B;TGd7=G;[9E,+agHW
Q2,ggb1Y-b079N=a@AHF(OR^K7N(]Z,3<2&T+X,EN+];0EP;ePWcB0-TH.F6Ba@.
,^6]D,\];TXK=6+#\fM+1]9C_J3?/ZgI=CQG]OfRdC2V-SCafZBGY0bNJV#155DM
<3YZeOc)K-)96EUNC<YaJR\TH2&(MY8IS,)1,;5MZ9J&Oe[FC3<E;\Ob(C=SXO/f
1;1F34Z]e^X)EM8/#1MD[>bVDYY4#@>52B]=GIC7F,A:EPF@0fB_<W:b.4/)\5<:
CT4<e:HI]QPf(GOKAc@:CJB8P^E0aESJN)Q;]?,-4Sb1VH+=1AXcM8_IB5JcaZA2
,2d7O)4VTB)GGWO<I6dX;6ZdAQ.6F/^a>K6ONE#+\FecDZ+G?6,[W?]YDSJH23b,
-#:ZfKT\@PR12JR&(-8GaHHcU2_b&F4f0M<2gI7E,F8WA@=2EP#_\91dR?3<f-gJ
+A46>7ReFCK+,67BSMC66\J)CI@MKLd:MeHI<b9O9C23Xa@KN7FgTM>\6=g4>DAS
K@3@_0U13]DY=?bD&5M:&;U#\g5;WX<;F,\7^VT5(dY_C5IOR:-8[.W;KVFAdGCE
a-+N9?,()[WVg.10+J2YXLG,/f55AbKW#1&[-==E:4;4VK:LW13;A_7Z:LTXF<WB
eJ5H)L^--aM],)K6L>#=FV&AJJ=2/RYXT98EM\(fM,0EB,YU7Z)^c9G3T4_Q5/eX
3^4X60NTC4]UV1]dFUF,^e1HQdb=#_a<RC5U<M<+N[8J3+XQ.M8bX.EMCJSO(&F_
+BS73Jb(cB+fOQB7=)O(82Ce,C;2O\Y1;(7CAZMfU#92e7ZQ2;K@4Y-30.7^)/.N
TCKR]=1QT0K8?DT??2bC)-Ta@0::[0986HJD0de@C=VOL1OTKfR9b8\C731d-A+B
5M5bX]K5Y7;B,X-^gP]4\3a6JJTNf9A?+d#LGSf.M_)IY^[I)g>Yg(X+Y53#V9R&
LO(#&RFK?ES3O4(UHJ_MGZ9f(aBXe#S,QU0@MO+TSfVMUG3L>CX/-S^g;(&WcKR?
;<aET_?(&.Gf3c-^O75M;-@KJJ6d2HIT^O[-:&L=)Jbf-@aT=.S&(eB:4b-TcAX,
ZE&F15aUgJY\@VHUIg#<0E[)^LX-UD[QKZK2LH>]0Z6<T@OSC4PX\S7O[-dK&@1>
0NfPfZ#QL?CTdZ3[BW09#^Y[/>GEVYD/#EQ>-KaVT3CPcV:.--(+dH+PQXV1X_DO
Z?\JWW7)YP+2c[dB7dIdgfbE:d0K)KGDJ&7N4G1g6L+d:IW:9b13GEbF\,cT+/HU
4MCDSfWT\LIB/RS1@]9eFN[+7&D&=WH#B1U:VW9X=;_CfG[Y>2<L,A.6)Be5dW4^
KZX\7J7dGeSSXG@N@,c>7LYC@R3G<=_^3#UYYT6E(e8T1fS1#GcLNZ@2aQXQMQJc
]CC+5[Y;DMV\G@;bf;L<QP#?VA(^/C]a;3gZGR/f7+LI4);TC)f/P8JKWL48\V[O
QJTX.&=Tf&V1X9/M.BCa[&5FK_Q;##eGZXX=9E#^OeBKPP@-/S/fTO[^d5,JQ9>2
f[F51:)f?:_^Z&#&GPT@WK:5(<S(Z3?256<YW<9EU[541-+3F\VUBI1,V^K(Wb=>
T7VfL7IN5TL9?859(+;3bUf6U9O-RQe+;f8]>:,a5@/O=5MAYEU=5&:^WMWTV@S\
DLW9^RdQYQ_/:X;5KY:.64WYJ\a/=L:S.-+W#Le^c;[;#?SM7B4Y;,BPI,Hbgd()
b9[19UQGc<D^>J#(HND.?=U_cd>0T,UW[g>4MZ+JV=Xb1ID_b49TSaQ6e14R-3+L
O<R<?0SA4ZDP(FQ[aZGHID#8O@e5#4\.LV;+@5VZbF9186?98VSVCd68G0?>e+8A
e-)a9cISZYbSPV+5N>U-]3((CIU/CM4)#)Ad-9I=WeN4?g0ZRT+]+-4C+,T&:CX5
@\gd]cSg;A]SaOTTOAV)a8C3&O7,GHUE@V6#S/7B6fMYKXNbcXQECQc/)S_-O=_\
KfY;6L,F[@T/7X7I<Q>7VM-ff[NZ8AP66..fRG<Bg#?V28<dX9[RF[C)H&4UI17Z
T3MRT_H<[5:eW+8Od<U\D=^Za,,I&Cc)U[aQSI^N#@4gcXX;[^>NRbJG+T?HZZJS
a#_@H\bA:CcN]+D/Z8;5I<WeJ>XLUX\I(@Z5fDPgV7cVb.Ia1TD1(bE#273_UdD,
=&QRa&7^WVab3^=@Z5-?.QANLCGNL[+XD:\O?0ZaO]].AB\7#9Sa4D2A=7&=C-(<
6D9EZ1B4__YPL-deVaLN<=ZOXcJbcE[8W15eS1N5Z7J-4eaNSC=CH_AA1ba&d=+0
9TNP@?LcL7+].c4;,SI_4G2^SR26\>0;A]CZCT+#_[,]0C#TU;ge#+3WAgEI[?B[
e#I+2AJOgIR]@LIf.?8GcHYNH5_DEUT0J&I&/QD[MX:<[7YC07aBVd6KCIa(K2E1
(#.IWMI8N9Qe717W#We<WPOBY50RW08/dTJH(ZL_^]7G1H-?[Vb/9>f<R3VWHVSI
[MEV9?..B^GLQ5W=DZC9J&TQF<4YR0PK9F_R,(.D4<Y:>MHb5+DCU:TK(,K.,_YX
\)2HOfH)=D+0aU=,e84gN(0QS.7?SM[KQ6M/@cOa.[DEeC-LXJBC5c@^W,4edG(&
NV+_L.\0:RQfeb(IMFU=ePCPY@B_7;)?E1:WeE)IHd?g5_Z)06?B\^.NgNLSLP.B
1&.M6TgJ:>0aU=ITH4&c+)W?O-9)HbL4<S>_\TA<7Z3>P7LgEH0?\;_0b:JO4WSg
LfSNUNfQ70J)F03Q.]O?4USVRNEMSgWed164TA=0Q190/(T>#\COH@X<(NE<bCAE
9WHMTd;OEN(#Q#1:)3?ABb2;:+5N__E[8_.c6LL+XKgHM4(OUdc<A760(TPE?.EI
45P>)U>XA90ECJS+.&]LT9<[ICfS2aMdLP3=MggFZ^].4Pgge3+T<:/=(5G5N98V
CZZgDO&354aAQc5DMQRVRN3^(eEG-D[J02?8F-DMUKgMb.I&/T0H/AU=_#K;E@SG
MOeQRFS)IBbNNMJA.CVU&dZ,a1W;(d;8.fUU38@^T[_4e(_,ad)=ceRRL1Sa@+\#
.;3gZfZ[J^XCIT^&6ZHM/b0#SLW(UKOV#QgV89d=O#><G9BJd1W[8#H3BP^.g0<G
3MTL>2>M.94JWOff(/<WVN-WK@]EC@7B=$
`endprotected


`protected
83FDR?(-C:ABX,_&U\?eC6Oc?e41PV+LEd5NS0,72eKc2M6cBFH,/)cg;aW>e^df
M@3H;9C:_5@B,$
`endprotected

//vcs_lic_vip_protect
  `protected
(7,b7f7<6PYA:,REN:O1EPFKDGdBNP\<WOU&deKgbbdRaI\;:4HA0(WRd,)896RV
AJ@e@0<IgZ,:Q_ENFPgC;;&,>8(Jc@YAZWSWH_XXNQG>Y<FO;CAOSPPEFf_QCH]2
bEc[L>ZR9(;C=]/gIB(\fQ_;HOW,(07=30?DD:9^dUa^-;Y1OFY\7VFP(S8CYb6D
+>W&B17Ob\443^dd/93bg3QHP3X.+\5T;7#]6/NV#J7A1B<UA77fOW[fB1)O1aHD
UD>@XSN_?eTBf2S^IDd@]b^-,:/O:2T70OW<;/JU]XgER83XUK[6_(AAWPBYC.9[
.JZ.bBe)E(]b4WWX?V.D^,R[@N6]@D+eU7?F^KNSHO4(U/ZS=Z&.0&c(fd\.EYeG
bKQ#6J<.gST[e<M&RLCc>Zd+H>cI-D1UD\B+:Y4-Z5dCQMd3PH_\\c)\(f<]6>_N
f<W-XPRI0[33JafI.+cBSA_74F]FHXPfKO<_/3e\+XWS)N(e2cgMEYaN<X\U[L#3
&A_+.6[=XAPI[ZO++FeFM\-36[]B\7H>W434-3T(9DFeGWUFN)QbN.FJ-Igg\AIa
[]A<0V80D(+BL+4UV4bN7><aWe^6=#fERQ?9I@d/H[NF@O&^fSb/]dF96cT=O;a1
aeO1LW5<==4+42=]Y0?HLgU[BS9d:^I?HfI1[GY9I^WS&,4L;63Y]N?;(]Ib8;9Z
U9,LGA>8Te,8)0-3#2#8:c20e@:OcN(_G313DH)YA-)&g-d0O\SY>DH4,),_d#&c
,2.S_Z3OUGQ:Y>V^LcfINg)HC+C^MH_X=JMVNZ><-e4ag]70&9L>Lg>ZMQ-9bLR[
de)VH0bTc.=7LI3MQ&XdQ@RfZ^a+\#ZP+/VAJE]gZa#Y#HGD>>]]Ba^F#3NQ#ZH&
Cc\&G\J)#,DdVNbSSKc,PTZ1?5Ea^,[2BeX#D)JI246E>C-)XWRK<TUHKW(,FZU>
ER3@XK>BO@IFCGF-3RLZ23OZ=A<fOb0GbPb9@1]I,5MR45YD1dZ_G]H?F/^IQI..
^^)74NEUFJ<M[GZIEGHG[UT9)^#55VDHK/48U?#]2Ud,Hg)\\BZ/;-0_?2-AM-2I
POJ80(-ZX_J_B)_W5==W<\J\d+?ARB6@]0[MB5O.\WVD2UaK7(UYL7/gQ632=b^J
0B=4F+UaD,+G2+IbN<&OR3d(&Z-CM#)@+Y#@LdCN?E1,YJc2_Rc=4Dga?IDGX.<Z
WIAU^/.J[A=L,0SO9Q1b7V8WKKJ/QC)U7?7d=.XRP:XVUEbZTVa@\7-6#Z0G.)3A
O?:fU-NT_@-4<+:f_6/=A)&6&LW#f<?+@WbbR5e]7>35T4da:S058@7=PX8Ma&UX
7Z9OcDU+TM#Q<]adbZEFY2#dM1Ga&2L61eC.T+->-@,[^V6?RFVgJ)O-?YEcK-C.
V-ASgD[dFg#IcTJU;8VA01g9D(]L,fD+QbR8@)038@#YX]RE_Ef>N/^aRVX.JaEZ
1]a\&DQ]B,faTXg&8A3[ST>eNS>NY0X+7]E+DKH+9:HD^Pde#-VT<V<5I4&=9Z05
^fa1MZ<HM;AMfEXXF<21,1R3RF,R^e,<KY>NQ>0BO<.TA.E6\DQQVg)H3.g:c/fg
cQE[gTCU&,1Q(3Nb:)[0GONS+8?b-+[X(HYD[=J1J?F[Z6,T/4-0\7A4cP4/efgf
QS<R).N.>E9.Ma\0=:XJ<GDZGI@@8YMMBB5?@W4?JA4Yb@96.\4G7Y/2B/gQ4GCZ
UU@XT8+e21C&2VfZ031J?b#,EYE&>_N_:]7@X4>:eI??8>_OMS/Y>-\AXRg-9;2c
.fZ0)\IJ^LY7YAP0ECRfI>;2[D>AfQMZ9E?C<2ET]F+#(P-5:de/:KQ@QF:K1OV5
9DD]D#I1eEg0<&8;PN:bZbOZ<A^-E(FIOJQE(BR4TH?T0f4@N5/f9LCEC>P@Pfef
/Z@Q72\Z:I&;7)61(6V?Lc;G-g2-AB.^c)_egd-<QdJa_WM&Y]ICb6/O@HG;SXF1
A(_&<P3g>cgLXNC=.[cNc5?&1U2@@6\&L_L@[#P;:f5M1JX,b4R@^\,EMa\^3;E]
2)4M0=W&f?DY<g_B(<f58WGdNXD0B4Z=4,GZI3<;(86)NgWI=YfMbCD?f9+-6DLd
\:7UM/PdII#J?);VU^a:]LJFT(LJ\De#AKY0YC8_/69,K8;dK71f0\ZXWC[2ID&E
f?[JQIO)@BXbVLA(^gXbU1S]]KXGQb<<.OW)_gC3LWLVG[_RSP\95.V8W2JIPH?b
:1BU;\ZR6KA4S;>E>+TN^Y8KTN5JMUF7#:R[4+FT]QF=(V5X)+F=UU?E]1(Tc&29
V[7&NLg@W-a:HA73QD9^E.XJ2W<2_WfaO92V2_b34P-bC]3^eFYX#e4)<^Y4gD&T
1P3Y(6./f1..Z_fR7IO18gA+(g4e3KYA9g+:=Z+W+]MVMcQ-49c1R,)#H0eT825W
@^LHZJAKGBa@[\NF>]K]NA8c.e.&JLKcPI.LI=P@@bRJ4c2M7_5:L3Z8GZ<4BNSH
OHE1]0XB^\[[0X(;@,JNcZRfZ^<#9aWMB&0K/W<Uf)]?2WK44NJC-6\AfHgOc<_,
@UI8Z@[R@I8VBcRf[/_[CE6U]GUeD:N]PTX5->aRUA1)=cL+>P-WVL2PSA]W:Y]L
=O359@(=OV8<(B9S=1Z^TX#VBa2HAaI#/=WK-OA6HX2OK\-B4V#?\<KK#gNgU-J\
Q0f:?OWQ3P_E,Q8a<<@Z\7HM1,W.5DTdFJ8W1K5a@8a]2W,dUHIReg+C[b2V@J#_
^+2/;0a<I\a^eF52HZ[)34Y_HB./IQ9VLbQV)SGOR/?&0BDK)IH)[)7VWN&4VaK(
B2&J0@(cH0_QBF?Q@D@b0.ARfMb_<&0Q69K.<&9cfZ-=P8E/W0)#gG&LE;SV1JS8
;2c08::<Ng)V;A0F??&LKY+MfCZ_g@(7GA&.8aNc51g5(11<,eCA?(JZRSU+XTX=
B-+<Ee;0-@bLY/704LA[WC04UF]M7,ILZP:GKZ_#9P(g^.:-\LWE2>7(_e[c:O[&
b[K(@cR7c.+<E>F<4R&;(E1TF<6<NJ\PLPS+,]1LZXgIA_.FV\F?/RW^G6[-L:H9
A.8#dIZ45:e_RL6JW0G(/.+5HN?@GTOQIFLKDEHb(0+fbU#DV8RUR)E^,a+L=4S#
Sf5@b:4\a3]C:19^]EOe4]155e.E/OdO\g&Cf6:gDS7XWU_6ZN>)Z#?WSC9=#>3>
3dFV#eK7.H4KLV,&;ScTbb[;LcF.X+/Aa/5Id&IJNGN<.;)@+Z[b[@>N+4D5-2gO
@P(44@UKXL0QWL0D]d+T<C]33bFV9YJR:M\@aT#?8)U5=XUT3M&ab67=7Bc\_^I/
M;gQD@EA]+,HM6:eQcK:T2HcI#WE)Sd?\&;U&KfR#ZSQ4Zf+TWFUee(B4QXH,T7L
X<VgcHa&M:8BRB]\L5\7Q5U]Ye-+LO8TME>PM5)8+KE1@&+U4\3R3^M7.G+bSX-I
7]\CG9ObV[=6<Af.gI;>RV>ObAHX8179^>;_5\ZNFL3_T^W#I92C)0[76R[FRBa[
bV)<+O.cU#^(&?7Zcb;.46=1^?=0Eb,ND,eCT=ba]KdUGL-/[.ge1-.=V_/=VOg4
D[J_L\0J)Mf[/5A]TT^9CV?W<AdJAS70G0>f3O^<S4L(,-Y@5XEc_>/+bX0O(cR7
&?D]\]>4L0-89JH7e//bCOb0UaZ.T:(^T-,VEQH;\3c>\_)S^A\f9CcF8.)\V2TU
3N;b#M4YfK8SX8L/d@TDgI,aB9D(/_:N-=.aA#:PHcCd/(e\5&E]G8fQJQ\?YOCX
.J>0;:I0&SDc+848J.3?K#4.@f=I?WOObbK:Y()JW[C(g6Y;ZSbR4efa[8+HF#AE
?c5c+S_b4ENA_1IUd3_+/)U:54.]Ra5M2@g/S]SV=ZX9SCDGV@DMfb&C]E/PLe<I
\g8;U7,GbWC.K\:[/C7DGGI)&92E6:(@>ObJ@YNVBF6fd#@A,c+2W<fV1TO1fUWa
V@S;U695XOTH^S+O<X^G;T_56L;@5X:]&(HHTK1DZ,]J3I[eZ06fXZ0Bb:3O0c.M
bPB_NNEdV6.Q5Yf88YHf#@:AD^K;<F>[MH@1&PKEUBM?FbNdgTTXeAe9_)95:D#0
]b;;ISGQQFBOKcBgR>dZdb/e^RN<H&)Y\1[-[3OF-;I1/CC/E<-H=W6gWV^#JeU>
M?Y.3g3^=\a5N.34\.,f5cE&3QNUETAc3#U@f1T7R)+;:B?88B_-0V:cEY^7Y8V9
Z(7bcgUO0R#:2+VA1]POZcdF)KC+F,=#.RU\F=R^]Y5ef(]b0:;G_0gN?5fZ4W@T
#^eRC_dYDO@.)89-6&\+KJQFEMSRE_07Kc)L\+CAH?e&E8+XH]+4?4]\EeK;2[cP
g#)O1W=O)X-+0\_?QHH&EDT1/K>8dK(-0TQF<7&GFfS<33&:@MC2N=H4]4S4S_E(
D\-@JY+1C03IZLcgdIaN<[e(O;?R<X+[F(@>M@,RgTCSWHc<&LNDRLO_9SVHQKZ7
&QCNN.@#N..VP)e7f2.e##1XBOY.Mf-1BaHBE2^@+R3Bg6;gUbQ;^E:KL8;UT<SA
:>A2WW7#4N?=N-1I7+I\/Zf_..#EQHYG44=B&/0HSH.^JN9WSJ3f9.abLUVR\]U]
,POX+XfRQK&+>9AK&bM3;BB/b:18L7b<#aTBbL>2ZVY^Z)/D4#3W[#N-0cN:I-(T
Yg2\_C5?C^]-&]U7ZTDgDEAHa@c,aB#KN<O3AZN\X=YYQ<7@>MLJ5MFf&E[0R^T)
HIGGWA.Z]Wa:8A,+aM&-_?/1WDG[YU[N&1[G#YQVOI87^@f^[X0KgX9NBDD7eNJ8
Bb<-JXT8,1cJ\>/57LA_M];cGH^UEI?gE:X#XT=1&UcH4)IV\MZOM\7T93CeE)E?
;N)W&+1;3WQML430_^2X@+:E,JM?FEL::_2f].G;3<.KA5LPca7(Fd+JHd1gS[B^
3&^+#b3b5Y<+K;A9cM4Y&(B+M8.K2#aH_HK7O>aM=a;_YGKf73SfKV)S]RSQfS].
&d+]B8>D(O8gS.OODbb58&#+S5<-H-#&7M)U?G8^<C08Q9aVGEW:(+/6WaFA@[/0
8+6]g^.OH;(]JH?.0VK5,.gHZ^fC782K^X17V(E=M.)dXOGb)B7,=V+E>?/@U?Pf
OKG=][()V>S=#SY;Ve]EM/AKD;&c:35&?g8<cU3J2GJLc6IR6L6LJL^2H]]5WK@b
DX4UUC_<;D7aPT]+gf;X&=O84gT@X\#/0HTBF0?C8.SM6PXdDe49WQF>A504MP+8
VFEOW]f^VB9-a-J(g-,Tf)MFSGF<<D#N:ORKKQ4e?>1([OG(Q+J)Nb=^(T\6=D<K
[?b/@Pd4TEFF\;-PfM/SbeT>95::12PWN\>Ne)YB0abO=H3X:L[IGW[d9a?X6&?\
<KN,]W7B_ZL143R?:(afbDKRFW4J_VOBRJ[e79ePdYNQbDQcXg,(N/dN2b^?PAJ6
Td3SKO#[XcE3)P70F:;:Dbb8,-S>G3,&AOb9YO\B>DG7XdKL8DBgJ4d_;Y9IP.L4
N]?WQe.9eO_-eC\LeBA7N9G]M./.X/Z8R6e4Z2[=e6>7(D:><<TbJ)-82^VKdO2;
(gQ&5B5_XLMZFK0S#\MQQMDKNe#MU7/6Ef)+=GO?EZT(8aWR76e=Bc0M,f)0&F,L
]@=N,EP=LR,)O]c?\6RX0A+ZG4bL.)N,^V\O/>M=C<@F-N1#/>RYbE#\#Z=P@XcB
6+9@==ReO[f>Y@E..^U>@TAI7,97)@^&0dWMAeVTY5PKAF]<PTEP\E@?;g.VDReg
ESF+==5GD1IC8_WOL/\_X=?@<C-7QHf9V:B+3@L:KHLfRT5HEg29?/-<c3<=D&AL
1)8cdaK_/d5X&[B9Y_^OfOA/Y@^1,/X)QEI=Ia&P[@@>&@c[?4S_bAMU>_7SRK(+
,JGeJ(Se@SK/YZ/GgJgA1eHRB8g0?/L?C=E^&Bc/A]cC3.?U;23GBT(EXFB3Y#VO
VCQ#6CW0FeQT8_Z<DW3JR1L]ac0dXZeW#/;-F0GVd@3K+8Q9c9WT(2MFERfCK[@L
KA&U-<C.[H-CUHL3Vb0>,(T4(Db&]\3YBI;UUJ(E&URP3@e\cNN29GYgV_[NPaCS
9?O5Fb]@&\-(Y>,Ba61cD-f>gMQH1Jc]YeK40+;c>KG<g60^UY)<M8^6LaM_b1db
A#RW#G]cXIdPa9WPLb)-^>@]fV)b[UT-D\K<E_e]OS=,#3DN8,E<[J;[R:M^Y<#C
aL45Zd+e)MM:0-9?8&:\&\,58afO)9^5E?8])&@G?4F&ZVJWL6;X(</dCLeJUg]C
&S99?gUd;XY5g^ND6YUAd:e;1BDGcF(UL1?7C_P4,C;?9-M1#ad]8:MXbTT/V=:&
U]>f-8<W<D(Z0WUXeO_[KETT)QBSR2XE/cfE&We/_SYcD.SVBMc4^<PNF9Z;R5+a
cBF18VC,O1e@39MOL(&:f;eL_JG<HGKVX\?1T(e[4IW6PT,97((2cdeR+-(YMD.-
VUSU^/-LK5E[KN8?a+efA0[B[B_Pg-8A@4@e>dIN@CQF7@b0FEJO@-ea.LAP.A,:
RY2HCRJN\P(Z-#aRDS3K5WG:WY96Rgc@e<;d@;R=QD5HOKT@(]?cV4;<MY#g13/W
38]W;4>K.(JON>>>/3H)\&^ec>;KX1&KNB7D+eTfW^DER)G55d;/<G3\HXJ+[]<V
,N@@B7J7(^-/ODNN#]/H/QaE.>9=HS(8=O?X9GW/N?4-G.)=R?,FRY@QCRgNRF>8
A4G9+&A:/(7.67OYL@,[a?g-Cd@\Y&PPOZP.H@@/LBZTVRBDe.g?E/X](Y;JW:3O
6OFTM)ca[L7aD:HE80a/F>GdHd=e7@<#)cDUV_20d78IeR\)=DXb[7.VJ2>(\+@Y
I3Y=R&8f(4A)a<QVPX65D]S-(C1VWI:GHgO@6HIENH<6I(N,47S\W>K-)D#6@];G
dR@UE,5fY1^Y)=55ID6dKU=PM8GPX97AcD[dW_bPeUZGEOE.1cW;6DQg2L]?b+8Q
e&9@^1H?Zc#2f4GHACWY)Z#))/a3O3E[#=(9ZCNL7E_e0#af=K/M;J\WeP1^VD.1
,10\_=)g(e<R19[9##BI[S)O03^[BM02KC^2\fP=5B)50)AGUE+18)K+@;[a-caA
CQYKWFZ1P]V3A4J=250J0Y7>=9.MNbEND^HVQ.<9QLf8Z@E\C3F():DGHb^7eSg@
Dd98dFL0U^2AE>,D-4cJa(OT[b\=FN\A[cQC>G->#f<.N#cWT_a6@BDQBRXfF32;
6K(EebC3b\0Ecb(LK,OC)9N4>+HK07<MfU)C.>\;U=FNa[#[##O1U/5g\QA=-d.)
97#L[0DT2^BP@)@Of4TN=HbN:Igcf,==_aa[A>^dLN:M_4E9)((LG/GT6gD0FfN:
]4g-/UbZ@.BP&dIFTO5?,X,6C&F7D/?2,TdX)D,:(#MY?Z2X1L#;_9S8a./[f&?E
a5CDMV3[]S2[b&^b8a563]cH=GRaY&376=]:<gZXH37/\1X<E@Q&aR)UBfRDe]\W
]aT4I)PMf>MB._F^1T__c>IWADd]Z<=RL9<DdA+Y3VN5U^4\gGQL/9DQ4Wb:KP07
J\S/aFgL.I8AV?A0,a:bP+A,8aVC(I]+.>92=0-I&=VHT-E&E.CPCN)J(cZ@6U@B
DH.(5<EF\@XOO5?E0&Xe:,e+Q]?)5g@g.H^P#345@B?IE1BEACH\EBJ>E(NP#5->
[.O<Z;?4&X:#RdRM\d(>7:D^#I9B_M=JO2KEU<BbN5BBCPAe/bVY?GZ97cXIH9/R
>1A4O?6#PVADXF#/LaY&=3.[[76.+_ID.7>cgbB_JCS,B1<N6:Eg1SB10MO2>.[)
a1]@H/GWbePQ(/:@9U1V=_1D>L,<(2Q&bTKY4f[65>A=3S+AbacaNBK_KC+0R.1X
EASY\D#NZ_(,8G9>d0HH=KeW[LWRZ-0)_G0^&aI0[Q4d,4^XXLOg+B.CJ2;N\7?A
2ZgNZa0HRYYgIAc8e(KTTQAN?,E/.OJ(>V]ZGPfb6+@)LQJaT-(8?]U4[dfRN?LR
:=Q]MI\eMLH#6O9,c)+M(cPBdg3Q@0\73^UDX7CN^TR<I\gIUXTc_J0(M?2K\d#^
^IXCQ.QXXHW(WNeFaV8gfY0aGV2AY<f-P2)B\RUcX/-8B23/PQTYgA[0IX#dc[=>
GG8e&3aM&+=NYcT]OZ1b4?^dL\+geUP.-0NTWEd)3-BJcU#YXM-&KeVK1W]8E?>L
BR3ae,MQMR.W,>5;1=Z@ASULAC&IgU;2WWMJe>Oe37:<ASIM2AF:.ZCa2_MUg(7c
/B-Q]N1Y5K&S/^cJF[[FHBXV(IVOI_@g?L0Pg-G+g2+QeCW55a6dL9\H[>9Ad/D^
Y03?><_^IS6I./a.AA,PC:9C<UMC+;M\@M0X1bIJ&[(7TGZfU+KfPc=76JSFg(f]
SI.aY:=TBQ62ObU>eHKR2RT,Lg^VR4&42ZK#g&#&4Lb72<d+N0E/;DHO5Y1?<?;2
6(WP273cJcGK:YN>e5EJ>-9A;7)(@:TM#&b?#a?@[@Ze5+D^6YGWPd4Gb_/S.>[6
O5d7C^(Q0&O@5DNfSTU,S659P.[Vb81N)d@3bTI(dQB_)]#gU.KT?GWJFOH4.QS#
18=ES@\BN<;c@9/#NgHNeT#N\KE:(K-f8e&[]V]>K)aH40C6D_Z5=K-9Re:68(bS
X=C-@8c7&1KZ41WO\YH]4V7Dba<V4H:@G]O?)S7<_&:e7A)#^BY(KHG08W5]/ZNW
W3-HOb/_(<,4Ue3(\ZD)?.NW33S,X\(F?N0#DeEY1^IA_VVDTdXe)#+R:O/HU8gO
\EQA[5gXA#Ef+aPYL)9LSb2WNQgB.VW4X[>XT_->?GH+7?#YV6@5]&6[5<_;]4\2
4D7X<:^E79HXV(HHEG9+>HOBJ&>.4]NZCNR>OG/[,V;GN=_#X:B1:YXMP3MY00^D
JYD/(d6BGd>EF[WBf\:)3ICdbDEg;fZA1-gB:\:QQVfc6D,90QKQK<_)@(D]JR=>
?GcK-WJV-@&EUA^DcKb8SLV4R&e20fBcL:P[deg+Y+W^7AB0>OH2>N&OD(AHIM+A
D08aNHMA\B_<:e,b3gK[5PA48f/9@;f,d@@#ZXA0W=T=0Ub:5G[R&aO8g7-#L\?d
6.B#R]QEDcCU;RN^A^<M5K.,J+9<&D0AWA4Q)R=W(4(;TY81&NN<]RT6g)X>E\UK
#bD[@09eN\:,)G7g#&Y?^Lc5X@0=YH._gQW)LOLHI;gJ@c0U74/-.6M?M^QI0fL9
ZcgM@=]e+2bW4W19RFY5,M7Nf1eILbF)d&7RMC2e4+b(&NNf_JKeJ07VL+fGBZZb
@E7bYFNa=.;7I6/9aR2bOQ/H8BVBC73.b3(QJGF(^NPf+X0GO@Yb4g#RKA?)&RbE
b:=d(dR:I11A<5G[g(g3I(<SY-A5Q9<5RWB0:4P,M\)cJPH/IN;KR6&-[]]7^GUJ
T\9;/)MAeA_I0Age8OU8&0L-BV28JPOYgP,5@R.JRT6TN<I&:U:&@fP88/B7[_D6
WT\ERf3GdG>R3g]Y.7>MR<I/Pf9KR_:>)cg)G;R=c=/YB)7SI7,9Md=ONO-IE,_1
GF_EeKeQHFDNA5R.FM?4d-9E[.Y.S]e?A3XAcVMXc-G>C]HX]Ta>gT0##]2OJXE:
?3Q9#GLU,1]8_Y[54Xe;T=R]G;:E.^bWRG]6-?541G+QNT_eXL=46OL@a:Qa6@S;
-)Sa6(HW;f<1cXe_.?XFCf9g4CT+4\Y3(8MCC<I@fH,;5_89Z?c;TfV^Bcd(#9Qf
EI,:?U:->/EKOU\Q5YFIW_INJfD\\HZM0L5OA2P;Ue3dT[:9<S66P+ef5_Y(g,0X
.gN\QAOO^&bV)KUJP6f/@F2@)UN-UgQJ&A<+TF/6HQ)8C/17MS5H8dd+USa&>WQ\
Og)&_eY>Fa2XI8[/6&#(2Ca+7b?VaK=S\)/N4Z-Of1.MdDH1HXN>6dZH@b]Y-Eg^
1e^NAV9R[aH)T.Ga2Db:31FN63G#;1R[?;]_;e>J1:&M_T9ZaLE#0g(6\M/#IfIU
RR^UP46ZZY9B7d;3[b\3W-3[R(19U2[\P_g:?1&<8MUQ?OCS2_V:])_WRD.GDZ;G
b7#IGWSZ3DI&C?.T)=X6,5KP(O[6A9)gT=7)=5MX^SRRG37,LY_g)9L0XCJE(D]#
)764=e^>T&.#\7OARF5>J#\_7I?NdM+RZ-^?V[+bdO;KfV#T4Ha/#B[54[T<#0M=
6cF\3<C\HI)CC1BS>X,/_DMXc5IXc5SGK_/1_PbU&A+cg;bZ]b=PJBM5a+ZB[/D@
7]8EH5/T.+V<V+T,5I);+.(YfDH=+ALTbQ\A\<C^aNB#EWIfJ72WdQ8d:70N2-8Y
LE479?97A9R>PHFQ=C(LMJB5fNC5_Z>PD6:D>6,dPG91_2-X1O^3ee9TI#K2YB68
,)NI<N()^aI\9N0NI=;?,5HK[86=_EeAZ[.C6^X5&>2W3]=I1@A^H>ecPDZKJH2G
^7d(f]g[XP<7NP2CM2#5.^8E@8-:FN1P\0SY:&b23N13CKB5+RW?#-ZeN.[I?,aF
,I?e+FH4Q.F_b=K,AT2_R&^NQR3U=c]LEWFeSBe7JJJQ50QB21+:SZ\O9?.(RHT>
WQdL8g8e1/;#D^2>X_][K#QZ+/b@3=K+VVXa36eJaX;7A6ZYS0JMYTUFTbJ7<1@7
a1JQ^J7=)#M-Pc?_T&PcE9\UH&PN+-Bg./L1U<58aYe^IfC/]4Ze)]O7<AdEBKCL
@15Dg]-P>;a><HBg_;2/URNL0S1CG2KH)&B0=26XB0Y9I.CD3U+QfHGK^DI_-5/,
D(NU_E\PCUVF[F#9U3/bc=f<C@RV=&R<9[D]8JB7ELSS<O0fB,b>ga/,XfA+]-g1
NR[C0WB:9O\6cB9GJF4X02QbR<e;2/cG@(:B2ZSd]Q7..L7CG6Q)X8H_e30U2@.@
:6BMKGZY[\\FFZ6c:?aB#.QJ2FFF^Q<>7LP(TCcQM=;W9MdW(X6MN.cACL((E,e0
I98KXMX30R05]4gO^ZBWP9I;\5<,E]HPRM.:F\/VG]H37@M+X6,HVKda]B)HLRY_
TP21.XT+K9\KcOC@.>EQ?V>A>0++R<;R#^Fe&aPAA,fcAI4c:Rg17A+:Ra(9LfJS
AZ/C^#AEBH>F&.)F1YKBP0X787L7@6>Z^BA^NLLVcBc@Sc27DPb5W+<.7F6@@N1c
gfI#7FP>V]&FfP^]X9^:b([Y9T.UJW-9NBO4XOH+TL9^S[9UA>D_A2FZVW+6DVY/
P6K^d\9SD>V</J,aTE5QI6GAU4A@9H;C425ZCaE&@0QO:D1B6/ECdZ3(0F;ZFEX4
AEdJU;SCU.R^1Vg_B664FfNSS>J];RN_b;XDc)],E&4&5/UY6D<50Q3+5=BD[_f2
--=9/4NU2S9a[I3W4aa6be@Y8-M[dHLGRE8bP:L).c+(>S<#&5ON=YDUTM_RQ\_0
f@80AT+I-HGN7=f-091[FeG8HN;C)I6=QP??[E&&BQb&M.]15MI96AE;)I5f97C]
@RMYI?^N\[0;g5DMP-V=2.bR&[Qf<RdZ:_KQSA7#RMOJ0Q/700cP+18Y(E=),JN2
<J3=6+++6+:9SC)X;5W:FOER9<2/2]b<&;4-eab2@+24H6.aeP;_dW8-@:+1OWVI
UC=WP;ZFZ7bYV0J1PC#30L?XF_^a/.>0.\B;=BN&<F0c_b6O[O>4,IWdgPO)T<@>
#P&?ZN:@JJX/1KeggLSXU6L^^]#R:_UZcWI<7ER&U>,Xe>2M@.A\#FQ9L7DD+=^P
P:b,&MN(XWQG/bSRNJ_>aE4IX02UKc_LDH=VHQR2>3K<8^+)6.&L>\[DD=[SJ@BD
VcF3KVEH&>VR&)Te@ED9[90/Dg^-7XI0?4=]4cf0BEVM@P_aD[1fJ?+fd52dg#]U
,dcHb79(2,U()6-KgcQ4#K^Y:SM2]e=\<<>I#E2?S>#&MaIN]cff9^WV]5=9/0HP
)O23K]<ZU,X9O\1@2C7R9Z2K(Yb#M,.(AVN?&=IB(I,M,()[f^V?:T+3M[f=(]&-
ZEM19N&M6d-bf_<K2:NS9R6Ba/RCc0S02c3_E<_\:dAI0Q^<RDW=_STVC>,T+\>0
@8XOY:_0-I,4,_^;V&4L9K9c4cWbC>57[K8L78PL:&64Gf+HW;@N(<9bM78&E]:b
SQV6b/Z7NF^_6(1_,0g9FS0DRYe6+GFD;CAPLaX8<:+.d^0TE.\^K<?EgW5VgI^d
I(ad4_c\&(QJ37\SQg+;O0L1UOY?1-e\WWUQ-1Ja1].?WL/4TfHX--PZ811D.Z04
YdYHY\4ICJY<G-J4AF2BH\)A2e&4La:NMO2B2^YBePAc43SGMdM<f+H^G?U7@gPK
Sa+f]XPAeaW)aBL&a\b49C_gP58:2\Z+=>6W,ge6FEB;FYgQ[eD#W\;,_B04d_aY
8J,QJ)TI?RL2FBF=/6eF5H;AcSHBFN8RZS=(?90,?1/?P?VYJ8c<b0+F(/>[H=de
JFWWK_cKE&MAEdZDU2HXb=b9Zf7:-3&]I[78,O3f82Z;cI7@f<K1WT^gA:]?B\0,
-c//MQ;/S/3g@ad2J#.,A0&[H,GTMMV<\,FTDF>:e.-)ZL>J2FZYJQa]Y?WTeC#5
9A83W)I.\bS&+b#ZaIL-?,;\A3\:_>U_dI<DVc(RZI(SPEc35;cg(8V.F(THB)/;
E-5:\NT^TN3;QX6(^eT2E_d]<egW3IQ?NM[RGOP_b)?J1NEEaZ/OLe5CYH/3YK3^
;>K;;AD5Q>d#+&870Z/X^-:/\ON:<&Wc:NX0bL]>)A<-^2,]3<REdM\RAFX+1?.E
U5::5D(A<CbBC<g_]@E>T#NGFO<PO1[PYdVg7:ZTXH#cNLI6,P,XLHYA=eG_7e0,
+9Z?VT0C2g_aU);RU@2Q_)C,[+YeUaC9H\#f/:I@VC[9<;+,<Q7F6GI&#E08.Y:T
)XHIK;_^V>AP]2C1C0Hd1.O[aUPHTKeKHHZ2+&Y\TcD?.Ce&U:0:,F]X11.L&+_D
bX\#4<Q-,OZY3^X<<?f[RWV.#FE=L[0B1=g;_?d(U@++8fK#:9P^9D-OJ9)UA1>J
BZWX&11B:VD92KRbJU73]M/61];]_5I=bAfH#FYS-FM[[VEOVYYM=##^=HM.;8C?
PW2>eZ<<K9MeXF&-B?A<:K.Q@NB8C85,UMb2YZS)2-HFTYc&R>/8ZVDO&);bA=gc
QQX[(/RLB(0]\L5PH_e[L&O]GZDe]X_BF>&aZ^FS461PH8?Feeb62BGG,7B#\0+c
<42WBG_;gS3c5EKUFV&HZ)(X\7[I6M[^PJT98US?@^d&S.bZ[^.ZbP=-2)M7>0g#
=0S/7U>gCVYRX8(f9eFZ@QGFJZb>H1-8Qdag1GUdY,QXFR3Ld3852P0U>(ER0@<C
TK.]WX]D=d,\WF4gS^UJ2KL\(1RBO:;E&P=B-gHgf#PdCfeP:W3MOKJL-@I,VPZZ
NA^)#b_39809YARDAH9R\;:U>P4d,/8W._c8&b98a=4Ya1/[2<_P+MBV5)70Y8I+
<24)\SRB].g@SG4H6fP[:\3JOU>HG?KKKCHW:(P=B[eH27Jf1XF^C1gB/W?=2a22
:C]I7EbSPN.7=4LWM>&ZJY31+YNN&39;1NKXCXU4:RXYL+:;?J<#d5Hd;J\+eN?6
J#,:]aKIZ_1X8W.;VS#.QIAKPE_.JUXH-9OL-)\7-.dZ4\FBFMG77C(T2_G59,#b
4LB3FV7cML2F9]1PTI8X<eb.UH,F4-9E<B:6O.^V(cZ\]R?T/MQPZ\c1e-22E<)a
Zb9FS3/T?.Wb/a1\QR^DfCWMT3R<UD^G2^_?PW\HM2Od/OR8D,df5X&\cHa;&T4:
cDa=:5XGB7.#E9FJ]?S:ZOcc8a\E\^[2fV.HbMR9MFWbCKUP+5I#=_cL)[2e/7F^
T#@LFOK3\6G?gR4/,[R^M[BH6Z_fDI=W7X90EXO4.I1aL.<+=@ASEa4(.N4:INX\
A\e\Yd.Cd<^,0DcPB^^_I\@dZ+fa5f2<83.Q_3Q34K-I&4/dAL@bP#J+)5S\1;00
KGMc8DV;F;gB;ZL1.#Ha;G9S[bX;?PL1QLdbc.C@M9CL7Q#88:<K_&Vc#B=I>e@-
W7>B9YNO4\VKWAL\,#U=;J_--bS7OZPT(9P5eDWK_/YS^F1OMf@]2W2X]KN)+d=,
:ASX^BPLJ.@>9GG6>LW;82d1A_g0L;Q.H@7)dFA^#^g&BXFdg:S;HYWYT)@,.[S3
SeJR_66f+NL<3^27)=;05b<H2C?:+VD/E2QI#6.dN9FcJ<..3XV4aC?]PT@Lg^;;
X6A@#]B^d(]1a04JA/Y3fWV/GB-B]JM2R1S3L]8_(A&gf\9@;^K@O:<K@/7I#UK?
6GJB_[)^[T6^cW6@2BNaM^OHcf7S\S5#B;/_:UHT[K2:e7+DV2:G&5\:[ZOH?:B(
#Z:/CXNQ0H&3:#bN>d>^)HHZd5U5Q/QZMNa_B1KQVZEEJZOTJg3KE@3.:M5F+b/W
<S\3A_J[&VZ+EN;H93?Q(TT1FV#J8d)>X19B6W>6C63UCL6HRLgBMM<aN5eL?(VB
/@):d]PNXYA8Y)B\)W:,b=J^(Z^0D:GE/3I.FH9DEF#a_6A6TCbd+G5R4&J]Qe7/
J+AG_4R6ecW7(_f];4,4^Q[dG>c;D)_9@e:Y<9&FcgE<2B^Z62K2[#?Y]dPXJ5AV
B]>eV-Oe=4CPg@-M[XC<?I/G_K(HgQ>6Z0)A9e=]\NJZGJf<:3V)>+Kg)]_M0-E6
-NA-OM>H/ZA;2NMLgI(;H\499V4NL<P+M\QC:Se[0LD+2#e:4JW4a&UP5[KV.#P3
J]D]>2Z\e0?MP?Tf1I\dGY;KV7714_O).6,V(\eM_7+Tb9TUMeGEYB1A4#\PdKEM
/@1a<8@O7[PHaNB,TLX@SY4KZCKR/g8[@.F6,S<CA;PQIc+b8=J\?08c65G:?R_(
O=bBPU7EdR],[(IJ<E3Z0^)PLEaU2>L;0G?<c8#?g?<?#=D9@A2_7I_UF(d9<9W=
7/(91YY9K^C7._cJF,YJ=C&W+\=H#>K59<XSS]@#ZKO0.;R,ZGIKZSL[Y+^_5gKD
:=UI2+e)2eIgb4]cP;YDI[J9V.M,4V&C:96]-)RQg1E_,.K8WXCPaXCV(d2BIX-^
DH=?;Cf\(@<89A_P[;4GER6-E2Q]e,T3\[f_acGA:SZO0I^>83AKcFK.J[R6/-b^
CT&EDRJ&1I6@?-7ag=VAPS9];N\1-\A[P5U2^=^#[K1^Ba)YcZVcF.8HE2]K-)W(
e7CH6M\g6ab1U^51c81#8MY1>P<Ce[b0HBW4fCX+.CG4-1)NGJ=g,E-Y[b?d23=F
V136\]ad^ZC;-Z0=A);1;Z<9-MacKR9\)QX#7HN^A]7@[=5=(:Te[\IWGZB>N\R&
AC7YeF<.K+)B<:?LV[^Z6,PI0b^dE8SU2J+?88]4B;EK#1PRO#&H3bZYBE]2Fe<1
S(ZXP;>\AP9ZHU<]3[1.#G+@b[].[HQ@bF10(5bHU=/]+4^2U.I0aLM[;aTKg<8@
5(fO.<MW0#[C^fJ@g#KUf.=R+bXAN+PQIR-+#T8J-=(3[7V6bP5CUUPK>R-+AIN/
LZbZ3#E]e,?]#INPf=I)e7M^T/_T;,A<,4?L3_M,Kd-XKKJS4X?Wa.-7Hf\KcT0N
5L^N=I1571gA7V>.AO\8C;Md3PKYU5:GdDP^)3,b[<L)LIWTa?>&CU-B..G(,1Y<
dXJOgFOJRU@0SdG+=IJT(3H\8S:4/7c7A[#GZVO[R3/G2XP,,H9&Bb9Nd0KTHOA4
5c2:Y.\8A]6X#X=J-SR.??C9e0#g8E\=M/\/K:\b5f6V1SfO;1\2L]+MY?7O9ZCe
BN@]MB7bHRJ=WC[SI/)2YFc.+ICE-/HRA(NZWc\YJ-[9D^WHCIbKe&ObU+fIJAL;
faOdNbR.Y,6X84EGe)9.aIGIIdA?46a)Mdbe\H\FVcVF.dCJHe80FW;.@Z>I48WV
.R6GF@H>?bA^A:=QgXL-<P=NKU>1e_?-J\=a;_QGA(,OO()_73I=[X5(YfKE&I;-
<WWMZ[Z@C_gHB5KE+_ZC^7;7)[;#WJSa/:7XNEA92Q73^3&.;VOJ[a;X6:RYCe=\
/eHK<J/>E1N8J+Wd0I;086^)@c[O=9Dc7g>^c4dJ@3PMM4PG6(#L<T3U[O3M\R]3
fI/-PI.Y]Q;#9I[aWK<[C7f;VbO2b<A<.^S06(J0;HAXJL43CO+Pe3,AeB;g0A.X
C/KaOd?SRDO]4ADI,64<]=_1YWRM:HI__4\fA&OW/[@+?G&SC,3TV35795Z<GIC=
Q=?S_^VUd0FN=OOXd[8)b0_LDO6N+CLf#e2[5J_W0J1&--:QBf8L:0:/SD&U6YB/
F9Z0J8T=0QM,)VW?6LeTYegWI[[6)AaLZ;c@1KF9RZ2^=;#5:LDEc+;Q_9fGPL>N
J1^1^H]BPK:_5NB>^3?+b01S7@XU5-A^);O]M2=T6dDAe/7G2]L/(E:6>49c]fO9
0)DA,6CfDFf3V)HZ7@g73R:G?L0-fXDAX(c)>H(1X=5A/SZ#?H5]F/dDS2_^HO2(
8.Y&FZ@2X+D-T]>a^W8SZ8,?\3-?2G7GXD0YX</TKY=F_D>eHIbgAV94CG<KCM)(
U5]N)cPPe<_\8+>_0[^+Ma5b-2-PeSLME4+G?0E]+K@BZ06e,+fbe<c(CA?3cEab
K=c6PJ9gcX5OfR/g]Z5]N8^bgQ[eE4VEaN:QQ@Ng<YDG\;WTe]XE];C4:&&U<,HG
fU^2I9IdF/a^0?67JOP=Z/&O;f0(I@Bf+<T]2FI1gfCD6);]XSEEe-MFXE=>)WF/
[CAPd7;DL0;MK6)>MF9_SE>Y2.@Z/-7)2+7YCPC9YRV]U=dH(Y1D6S,e\D)2]&aF
7IbX@E7KIF04C[7>.(UcZX7NSDFJ1<R;I)_T_cQL9QT?C-(+]17(TIT..(:X@I<?
&b&X?+L,=Cc@W@\5M+E<#@9:KRFcQd,Vb4SOZaeE=@+6N-D..WfYe/J40ZU1dH.P
BX2I7Z96/:gK@C35N\ZR+.DS.[I=?M9FQOM:G(3#Q?P6=SY9L?,TZcA<V,_8B>V-
MfR(EEX(R,WH&K^TCQ_,/0IXH;b7H&=E7GMF37gA(UX#ILGEOF(A_:.@^Q5ZI8/1
c3K=[NU?)>.ZADO6C;U8X7)ZaF3X5QSfM&,V@aM4VNPIYEQ@X\eN0[I>BLb?6f/f
_56047G82K^dY<J<9PO#\F\#3B-HgI(.R.6BX+]I)U&#Z;#:H-OdF1CSe30Y,3:d
Z)BA^YQ>U2Q@61/TB\aIK9aX&^FTS\LWJ)>\a,f=7@.@=5D#KDT93cGg>4Y8E-()
36DHFG;EI;.+?&^[(Hd?#=K2Hf_8F9(E69@DLRf8G?;CcJ_a0NU1^/.a@>+(T1AN
eW[g3V2W#Q7,<EfB[EEC(@:Q8K1SHN^:K_a=a^?FW2GA+KF;+&S.R^N:393V,1,,
0gXJOJG6bNOTYdd.RWgb(8;Y<fLfRC;B7O4##D[X4?5#bK4ETeSf&#f<??,4+<FO
+I=V]\.3FP@.X)@&7ZRg^)(f,a@]WTHf<(^5AcSeL,QJ_fd+fD5P7UJ=LLg;@:L(
#B(<(KRZ;caSb:+>6)=Oa2<bZ3B@?c^UK5Z)IQ)?:]0fde1P?0^&@?O\WT,A(QQK
C,9JFL;^fXNL>0HH(VQT>,?Qe]F<gg;):@,1(E>A)-/e(VX@^IB=RGbAI3]<C;B-
E?N-3Z6/S5QR\6gY2+/_ID8AW(<<?&+ZY?(QdGLCgE=1f^]?1<Y2\&]]IW1L0YLD
>bAEJV((ZQ4]bUdNY/)7]HUWEGe4U-&@L(HD:f&]8_fD)Q#gKDX2:#CBSK8)QGG.
6a:^_LK81R#2VfV+^g(/ML?NWe=W;[1&.X/KU>3M5>g5<BUV=>UBKg9@]VN<8R[L
CW:8dZ0fDaC6LET)SZgX>&Z24E[f5;VLg^gOIc:LaD@\;_NQSS?4SUBG(TJNVBb=
MD;6cb_)(:?/19\9Y#XU>\H</7WEgPf@TX7)dUgT&UP\.3F?N;JHRNI7eZ//)AO6
b15V(b[2aT#c/\/cYGVP-[I\b6=?I1I=HX#E/)F)-U:0J]-4L3Y(N5^)32QNe?ZA
[QW.&-LcdQ,DS\bXC5cg.^O7AgB+R]>F]VE@NSU2/Q?K-Y[QaEAKLDA.3,)HUD4+
07J-Mb.L^DTE1MZ2K-/?/I>1][(G=H9H+]dfIf^gaK-SJL3DVA^;:R[BO686O1CF
/F89]9MIeMLQd=N]KFH1f2788Q<RIZ\f)De8+.Q7]5<_(RJd+6ce,?KXJ[gH15_a
B^LH-)X?L.S.P=FM7N+.-SaTUYeIcU)7LU.I>.cb7>XA4<F[>AI<,R2FI2F;:?]c
GC(2S>Sc/QJL-QXNU-Fc;Fec_8f\^STQTO:]G=M6gS^@H&JL3\X:6UXb(7g[I-C,
(^&U+(6OK7^49G&X5<5XT^\;gc>2XGB)bL?&YQ2aPUG:BUS<77MY.bX0NO43T58F
cY(;f#LL8C<2]gMO#Z^;PSe6LLYLL4f@]HP_b89OX-)cP>)P?#8^J&V4.P&g#;39
IL0OW2DJc@)_a5)MBX(\WGPfU(3NLILMW3G,.C-P=;0+df]Hd]8VP:U]e_.S-HLW
?.(@HC?/M:-O#d]a<&6<L]Yf.32D?UIE/#4:a/)81aI;]8E,,+d4<XE_631K7I;[
IH/>_DVXWgK#RfANN\905Y8/,DfO/A^#Pc(8X\QW:FUXDcPP9[[Sf-]B3@cGHX&I
Re#4T@U&S;S:g[808c725+Fb>FFBXZ3W>?T4_I[2V?Y^+O9=M9Ye,cV>C.:?/#(W
]CKg0XMTcL2fIHH<5Q)g.4P0[:TEc&3[XW_(a,RX-cT)\-C#@:Pd<(FWU)d/aTLM
4C[[Yd^NAe><LU./D,A9)F>JdB@ER8;5CfPa.NY6ISa#,bSbDRSFe?3X.57<g_:^
15@K?.+Z;#F_;RCe<V,eJ3]V\W?<aDR(A?64ebgSX:AI71./V2E(-,aYabH\GHA]
-^gMA:g4.Ec6^7R&[=W[\f6:Y:[LV@bG4C^E#I&O=.FFQ<K]g&>\)T7cB^U(-FAd
4\GaDKFMXBM#aceD7L],QWcbFI=B/)#:0#ZH)1)LcGFH3HD1R-B0GV?8;?Z4JNGN
UFTc<0[L8P0\Ab(EU<Wbg)GF<-We0eX0Je5+2M(GKS5+UH3=gB]c33I\eP307cbN
[O1MDg^;Yg2+:XKU@I7-\E,^L#VY#^675Ybc:a5_ed^;O7^CC&\I3Sg)]&J.@=,.
;=68[Y?O3.I=1L633UK_W^;:((>G6C+?[WNB=2dHIIagWcac?D([T+=a@3NV9c2W
TgEK(Ta=QI91bW,_T#aAaZB4K-&XCIaaU41Lb</9E3\9F^CK7d;[W/TVJ=WM8=4@
N[BX-S_CE2<_C)g(+/HVU/P,^[S8@L2HUXSg?:M;NS8SXJQPFSQ[S19gBb4G32KE
Z];)P-1#gaP5\[SRUCU.SA@V;/EHTZYFZ?LOcH\00,05=++,,NF]Z0-C#R;(9AE8
A=5<TRJAJd:7\>XD4RWEFHJAB+6F:6U4b-fBM[3;3(W#R,DWFA(]ZAHbFF:I+^NF
;LBQN-/fNJMRR\gXPf(;L[,.]EO>S.G([U)DCBD_YH2[US.5X0Z]WR]6<fA=>-G&
2YJVB^P=CFeP(LE/7J>3K-R>Q57/FCS?I5eSeeRPZYc-F[M]\9_gUYBf1WM-EYga
]0S;]=g+dZM)56-26,a,4QCH;eO90+BS069T&::)L[_T&4)+86(ZWQ9JS(/7#H_X
1=W;ObCP/3]0X8FFP#Nf_>70@L2191<)_>K=E>=ea&N^9<MS<)@:D^C.<3ce_6<D
/Bd75K6A(dK7#:JH,(Q=\;U\KB42QD)(]fN9ZK.YbU-F;08QDOO[2c];>?^P7H+T
6X,?ba=-N=SA)JGWA3H\IIK:LUD,dC;;,NZEQIdd3-+^UO_T0NFD.O6;8]1@:/-f
N+3e-\01\-CY4\[L;[_,K\8Y=UdBW\#=\(deVFF?A:\;LP,c^e?IA)I[DY+DBEC<
Z]V>3Ggg:<NL8[f_,#4cC6eCb<WFWY2S>C#6.F@WFS?U8WG8?JO6F4eN,CR;Q2P.
WTDf;X)]CaYI9&FEa:eO0/3+O+Cd0BfbU[M;9gS</FQJQORBKf);WAbGdgU67VWe
[FgI/(7/]_VSA;CM63>f=@R=Q#/EdDHR@C^2X1SSb;Q3dF+fO8Jd;+B9^TX^=3K5
2R#]AD_QNTUd4d5f7GSG,UEMEcB91C(^faKH6^E<7db2gDd(PWZ\I&UB#)HWUH9V
LC/0cQ0gQEXD8]-P/dA39,g<W:,O<7O;/Z0/PQEI)_9(YG/f488-+6[@U\C;F>WX
C>:SR>G6--?dfQ(IbJ2cBYB(H<31=_>SD^L-OH.3R9ZGBSaNJD0f)aG>W(SH_HEd
G&=V<SUG8-2gL_&fSW7,S<AJ0BOaL2>&g,7gd1#TeO)MV?1bQS:cU<>&M8[EQg4[
/](R>gGXa]),,M05Q8^<FW5XS/,G+]YET]c.8TD]gU4<b:<Ia(:E&bRf@g/HGP+O
N<PX-A2Cd?Yb-.f7a4?M@<JLgRHJ43N9_.6^[<A4eL<EJ=.6V#eWFOJeOOdWUQ@)
ATB1f4IYFZ\>Ggd@@R;^7;;g]BLT2c@2<9cH/c]VUB5L].3.CaI#3I>-\(@]0V-f
282(d1)RC,XV,D.9d7CV:EEXR@8>G[3US4:&:LB\6Kcb8M=^8X[5G8ZeF9URIg^:
[#N#KQI&eHX1##8UZD30JgL.aRR^R>2J:N\L0^=5Wf1OSI^,VKN\O)1^NPMb1/0G
[EcF<&KB+MOK9\UDI<=M-^]1gg5Y=,;L,FJ1W1W7F-ggVS?,5N=bHB,b13c5/Df7
+WP?#-IFLDdSXg4,(<\9,,W[N]b<^?H0cKK8G#[eNZ/;Fg;^?..^.PR4J5W.+X,^
C(=W^eKafBQVBc+AgA1AePfHaTRY-A<(bC6]:BLTA/B-VUK3e\7@N(4&8UJ?.R^2
@Q6[#1caR&7&3N:9,;)F,--.?36c4\S>>W[=)&&;9JY-O;&_7YM1AgE0+H;c(J32
f+PM?ggK8_)d8NLP58[XI<R\#KId?R30(N]S6,5Y[+KM&7)^#Qa;\ATGWR3dQ6<Y
RLJW:&X:>R<L/.e5#=bYU8gV)9Df6].;aZ1?f=7;MQdMR6(&5cA5R#&[:eLFC7K;
aCEX0]9=5A_YgW2T[7.T\Td]35]S.P&;FF_4cRA)Fa15WcHOe6/_^\.LYfZd2g<W
GIM=7b\V+9ZW[O/Q817X[dd.@D)6FaCT<=\:M>E<XX0fc(,YMTX/Lg6g.dAGS4+b
eQ.8^fbW\Z,C-6;;gG/?J2?8;0f^2[?+SIMRR/VF04S7bJDDRQ&a2Qa)D##3M64&
e(W9b+4WJ:-+S0?R0YFb]Ha_gT<g/gIQ5E5H<?K)XFQ2-]+>.cGM#5.Be)C[<N3B
K:(_CEZ#E8-BBU6AJaL>=ER^BTa[5b\fRZNDBVN7E]SM-T9eTZ>DF=(gb-<)S55L
AXSA2.>#:P_0+M<=@N-9^R3&L_g:DBa/c:FDCP93e@B6JHPTK6e\(#3R6C38<,J7
3X<OG2+3Xa]4\W-PVb0C]WeF=EUL+C9CO>?Z_QAA&(4EF917CKV-/3ad8Uf.R-)L
VDH1c,J8Af<N4]e3=]a@>_R>JTX(Zd)HXT0Y=+]A3/0d3Rf1^LROfVEcZ-R8UZMf
aVNa].eV/f?J_LSa6+14?a8C/9TN=D]Y?UZ<?([V[VI8C]K#Zf)E<Ae#^L+de8G?
_>07E),USDJ_b_G1VdHW@@IfQ<.e.40^gE#gGf@IL/QC4DU/cdD>IX(+)M<)[&+]
2F=.D4@+:T^XC53[[gU0PUZHBPJ/29Wc&X;HC]8Ob@[)]P0&7;+JYD99M#-:cJ(K
232Lb.QZXb55@f[URe0bc3<CXU_8/OJ-?@1)NY6EA#_MR2.eNWgE1]6+I4@Q+]X#
RgbA4(XC3?TS_R&D?2AdU6+:)91Kf@:<Ec_N.O\^5?Da_[gPQA6Ia?4a#>>777-0
+:Mf7FMP8=N(^1]VH70.X#QF7W5Y)D=W2[Z9B<B_/8NJP>)X(/(>#\aC#VE@DV],
OCF^WY]?\CaD<ZK)H9[CC&+2EQ/b_<gI5K;IMLX;N.&@gf&7O_FUEc)=T]1)8R]A
NcF4fZ,fB28N17JFJVMRLU5G<_]\>XQATc/KBCE,V-4a&cP\@]-_+;2dfV]FdF76
]3MgR/Fc&??g^Ha(AHe#d0:<<).J&<L=,?)PZNe/Nf6U?P07\:=-L,NeYa&Ha;CV
S19)W5O07E@P9\Cc++fcX+IeDfOXMdb;RWOg85#C^S/UC$
`endprotected


`protected
e?@M;#+S=G[3NF;U^D5)(<88;ZFc\X.SKB2S4Q>>W>)[e\7OT/cN5)/^9<L+9=#;
-,=MaHUI9=N3,$
`endprotected

//vcs_lic_vip_protect
  `protected
[:6Z?&NR6V9f^\D=L2ZBWOYO\\6:7@\@760d:8E[SK2[A0=afc:C.(D&7BM[)\5M
ZX\6\;IaIgEJA1/5X,B/SS+F6fbH^)?/N&e^M?2.7&NZ#[B8+UU^QbHJK7W&;JcX
,]Y\5F:UE3N,#f3Cg,(KcP)F]R=6U3(6a#fgeIFcc5M>E9B4c(-a1aeA89<<CNGb
LKRCNYbV;@Nd]8:53f1_31Q^Y(UXSE]R<[ZW&:gI,FOD2J7&68<c+(FdE\Q):POG
E(&^_Ob.UBS?bBY:-@#@b7\HD3#L\B4I&3B5FM.G]BXV#^?4EQ]RYUgD65e_OBX@
\E?6bNJ?,NKCe.;1<</8F37dg1I^;BQ)43D^G?)9gV:?O.CLJ778Z\ZX;#(21(W3
8L,G/2:\;UV4X?dCg3/^ZPR;e6<fUJHA,f>?eIL/G?JK#^Ee8^MA&HG1?>U(7[#^
:-IWGa,c@g?L/e/;4[Ka6:C]\BOFC,DR;f[N0N,2@GVZ;e0=]8M&0RO62FfSM6;V
>)2S#eR,34E(Y0E)adaG:&5aeLM@5(b^b(18W+NPQ.:Uf/_QRfd7W+g1#7aL78T0
3?)>T_d?4R[GSdF0?5<DD12?f&_^D:-XST[_6)/T7fG8]F^PM:>:L+[;=,7<LA()
H(0]I2=Z^6>QeXUH<M0+A9#9+8OFEMMKAC0QfEL(]-9=0JE8<ES8GP(1Z5B>56W?
/7P[L\UK<TdAY@VDg1?a50<+:6dTc+A2b25V)7db637;;7MS(\T<fMQ?f8b7VK?=
C8c&a:6aA^T,#aL918cYL.E5FM_RNRC7ffV)bCd2e)OLQMN-UDH=c<E:?]\.\4c[
UL30G<^R_3Dc2TK8^fRNJ(I)4+1]TV>:.VgDBC6G>0bf+RO;G2XL:V7>F++@&=<:
5TDWUJ(XEE.EfN(E#I]L@F:f;U@GeRL#[4efBU5?YNCGSC48^B:TgF_R]:e>SR8S
]VQ?bX/Y(_ZM8:ML3:154?5fF77\5\^LMYV)Kg(.62OG6Z-IGb6+TOVb.c[ffH;U
P-4fR0Cc((=1S+\_KQYHBO:9C_D9-Z1U::I9@O4:5;3FS-0LPEVT28,F0775K.T2
D9C+gQSef8]@,J@;FN<G,=;D.QPM,Q[aWTA4X;[\Y<KS8XX8GHB)M;.XcB\3;6JS
T=K]UORR#^^S0;BTYOPSA+e\Ag8Y[2U,)[CgP84D=?KI.0L=/UW^+TBDdbg]9H0/
W@8QfY.4P0#7a].)+J_3NO].NCQR-V;[>eeIF=9Z4F^(+=EdfS6<3IeaK#M&e7-d
_PeWbgZA&@;]>)5Y\>1<,2a0VK-bW^]D^O3^&B>eP_[X?=INWd:&#Fe/Cc)GE7F^
VL(R+-#b\B1DQ<4d1D;?PQA=P?8>/8WLF+[X=Ja+=^V;F.@)7Y>92,M7[FRSa-3[
Cc4YA+PSf3>WcY<A3P0XYV6<5dX6##SE61aa[C0PXZYOX1(6N>gdB+07De/DDG2#
Z_d\L7UJT189H=aGLG^HaB-9L0a1+e<^Q=OT=7G=YVfFN-0Q^b=/eb#7]=--Nc2J
Xa2W-7T<A?]BI,H3(^5gUMJQC,]7/g9KC&&<b>65Ka0[LB;G_N<&&EYTS-U#dE>P
<E(HJY8,AAP(&#6VM9OUMZ104XLMg7NU_2^W\fI=E&U2b^.;0]WT[R.0=TYF;aP2
BMQFS8LN8MaQ?IZW(3?OD9E>]AVP1(cZV<0g[gKITVD8,bQ3+Kc.1FJ<4,5e199X
YQEPOF&=SKaY@OPNT(Pg>1Aa^Cb_7f](=W[?I4cHaZ-@5a#?H_+e^g[YQ\gHD3H3
]<]9_+8Cd,L2A^Q+dEQc0E=(fEQ,b):7^d@>g6_06TD;TYL_P,C[I@C>L+VcNT,C
PaN.S7ffBA2.]W>#NN2HAY6[Rab04JZ)_?UC285@UP1P=NDCDQcLX@KZUT/7E;VF
,5HN-HK_a17G^W-B2+a/Ba_Q=fMZBP6]K1=TdA8ODD-Z?H0OQ[G/XH]0C7IG\I?L
,Z,PTS.A-DY.Q\PCP-d_U;OXNNR,#1D+gZ1&6TUV52:P013c3<CT[+@Q.bKXOH0V
STe-HUR,=6\^,V(9Fb6\D13(U-P6&0;G>FDJ8&2Y.//DVHe&Ff6)-8Pc0;].:,<Z
R8,>[\#E:J7/DOJ-.C[G>If01eSID9W-Xe25LEV]fNfM:=<-gP/SMPM2026b8:(Z
S&(?E^aYX2d)X\;:B#c@RWFIV=TKAf+O#=YWXb]1-Rg@7HOBD5T2f7-,K27OR5XC
E4<N,-Z1HYQ?.d/T=UGE^1LEM4ZF/gMHG+L;=0HaF;A?3#c@X>A2:T,J(_Y>VCff
RG1La]dM&6VB9O(F0fZ;a?=\UHOR^^UT.,N.>8V@?#gFEG4=bV8VHb/U3I3gESeH
#=WH.Kd:.&5^DgRcdI9ZOTIYFKAfMcGX&4H6D1R/=)ZN9<KC95^.Y94PK+A>A@W-
M#/SLd;DJ?#c&-_,.(g=V3d8X<=JO&3aBFA1J[fM(R&YJ/<]25)??KQ^/8XS-->N
3eQNW@<d^^N1WcG3#L0:2-dPL08cV7bR-\[Y.BEPGbMH646D3JI=@>-Nb[\NU>_3
6FOP<QF1P[0P:MN(7FI7bBZ+9A_B\-6_Z+TCg;W\83/U1Q3XBS>U]_6,.\V#Q45V
A+-Td9PHe^R@dXf<;8CcXLRIeG75&7;VMTF(LB,3\[Q6+#.M@6E43B1fRB>gK(HQ
caI(]N,LA&33O?Ad9HgI,3=J@K(6&bQZ3RJ7M)8>a&Rc.;MN\gV2+3.O=)@;JA8D
PKB@/[Z;STcY>NHI</>c_?VQ9^_+MO=d,R=?QQ&W(\^Jg2e-1L8VC>U?<Z7f=fRc
B>6P,@H_Q;5B38<OPQg,.6=;f\V::[HU(AcM0/K(^c@EbL?3E7G9M_P7cH]^WD&7
LML/?;]?.A4^<Dg8aQ^<@#ALeM14>/8.&D3W+?)a9A3J[[I-cfB9Y8\CX,g1.BQ_
DDI08VN\c9VO6aC7#T+QVQY9(\5A-1>RPG7=e00-#5e0BF1S@DI[TP)5B=MKK=##
\b7]S\W:BFR+R&]U<U5aXd7U.36ZN^dc>&#P8JPT1WQ#e,;:LPVA[;3_6&>@6D5C
3;DRWQ\9I1ZE&0^LHd#T+81^-=82Qf-1eD4N_#YT_ZCbDcF&Gc]Y672(a<Q\\.J4
=(>:OI6^:Fa<a8(a&T_A2;I-6[NXV+B2?9^AYgSB^E[O#=ceXJ;28IEbM_V:D:=V
2]O8I])S&-695>@aQ#V3>G]E/VTcLeeMXe(C63H-=_<5LgP1DFAc)dRX=,HH@VP;
(@2a\U3?^O8#f)c&:c;(-M;K&,.Og1ObKJ1EF^dF]F[OGJ=O0BMG+<f[ZA4I0_3T
>dU[X\,;O0^1eKU2P);.6S68AXdV6O;b>RQ;fVD6cLcYca^?G:WYDZ)93&H)BLX+
9^-5_5?HJJ,;J?NV^UOB+f-(NH;),BgI?$
`endprotected


`endif
