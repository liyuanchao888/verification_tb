`ifndef GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_COLLECTION_SV
`define GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_COLLECTION_SV
// ================================================================================
//************************ START OF ACE VIRTUAL SEQUENCES ************************
// ================================================================================

/** Base class from which all ACE basic level sequences will be extended. */
class svt_axi_ace_master_single_port_base_virtual_sequence extends svt_axi_ace_master_base_virtual_sequence;
  
  svt_axi_ace_master_base_sequence  coherent_seq;

 
  /** Represents the master port from which the sequence will be initiated. */ 
  rand int unsigned port_id; 

  /** Represents the length of the sequence. */
  rand int unsigned sequence_length = 10;

  /** Indicates if this sequence is valid on an ACE port */
  protected bit is_seq_valid_on_ace_port = 1;

  /** Indicates if this sequence is valid on an ACE-Lite port */
  protected bit is_seq_valid_on_ace_lite_port = 0;

  /**
    * The start address for the address range for transactions generated by this
    * sequence. Applicable only for extended sequences where it is specified
    * that start_addr can be provided through uvm_config_db. Typically 
    * applicable only for sequential access sequences.
    */
  bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr = 0;


  /** Indicates if start_addr has been passed through uvm_config_db, or is directly set */
  bit status_start_addr = 0;


  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 

  `svt_xvm_object_utils(svt_axi_ace_master_single_port_base_virtual_sequence)

    /** Constrain the sequence length to a reasonable value */
  constraint reasonable_sequence_length {
    sequence_length <= 1000;
  }
   

  function new(string name = "svt_axi_ace_master_single_port_base_virtual_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    bit status;
    super.pre_body();
    raise_phase_objection();

`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "port_id", port_id);
    // If start_addr is already set directly, do not override the status based on whether it was passed
    // through uvm_config_db or not.
    if (!status_start_addr)
      status_start_addr = uvm_config_db#(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0])::get(null, get_full_name(), "start_addr",start_addr);
    
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
    status = m_sequencer.get_config_int({get_type_name(), ".port_id"}, port_id);
    if (!status_start_addr)
      status_start_addr = m_sequencer.get_config_int({get_type_name(), ".start_addr"}, start_addr);
`endif
    `svt_xvm_debug("body", $sformatf("port_id is 'd%0d as a result of %0s.", port_id, status ? "config DB" : "randomization"));
    `svt_xvm_debug("body", $sformatf("start_addr is 'h%0h as a result of %0s.", start_addr, status_start_addr ? "config DB" : "randomization"));
  endtask

 /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

  task send_coherent_transactions(svt_axi_transaction::coherent_xact_type_enum master_xact_type ,bit init_cachelines);
    `svt_xvm_create_on(coherent_seq, p_sequencer.master_sequencer[port_id])    
    coherent_seq.assign_xact_weights(master_xact_type);
    coherent_seq.initialize_cachelines = init_cachelines ;
    void'(coherent_seq.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
    coherent_seq.start(p_sequencer.master_sequencer[port_id]); 
  endtask

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    bit is_port_ace = 0;
    bit is_port_ace_lite = 0;
    `svt_xvm_debug("is_supported",$sformatf("calling is_supported")); 
    if (port_id inside {ace_ports})
      is_port_ace = 1;
    else if (port_id inside {ace_lite_ports})
      is_port_ace_lite = 1;

    if (is_seq_valid_on_ace_port) begin
      if (ace_ports.size()) 
        if (is_port_ace)
          is_supported = 1;
    end
    if (is_seq_valid_on_ace_lite_port) begin
      if (ace_lite_ports.size()) 
        if (is_port_ace_lite)
          is_supported = 1;
    end
    if (!is_supported) begin
      if (is_seq_valid_on_ace_port && is_seq_valid_on_ace_lite_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
      else if (is_seq_valid_on_ace_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::AXI_ACE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
      else if (is_seq_valid_on_ace_lite_port) begin
        `svt_xvm_note("is_supported", $sformatf("port_id('d%0d) is not valid for this sequence. Please ensure  the following: \n\
                                                 svt_axi_port_configuration::axi_interface_type = svt_axi_port_configuration::ACE_LITE\n\
                                                 svt_axi_port_configuration::is_active = 1 \n\
                                                 svt_axi_system_configuration::participating_masters[<master>] = 1", port_id));
      end
    end
    `svt_xvm_debug("is_supported",$sformatf("is_supported = 'd%0d",is_supported)); 
  endfunction

endclass


/** Base class from which all ACE intermediate level sequences will be extended. */

class svt_axi_ace_master_two_port_base_virtual_sequence extends svt_axi_ace_master_base_virtual_sequence;

  /** Represents the length of the sequence. */
  int unsigned sequence_length = 10;

  /** Represents the first master port. */
  rand int unsigned first_port_id;

  /** Represents the second master port. */
  rand int unsigned second_port_id;

  typedef enum {
    FIRST_PORT_ACE_SECOND_PORT_ACE = 0,
    FIRST_PORT_ACE_SECOND_PORT_ACE_LITE = 1,
    FIRST_PORT_ACE_LITE_SECOND_PORT_ACE_LITE = 2,
    FIRST_PORT_ACE_LITE_SECOND_PORT_ACE = 3,
    FIRST_AND_SECOND_PORTS_ARE_ACE_OR_ACE_LITE = 4
  } two_port_interface_types_enum;

  /** The interface types for the first port and second port */
  rand two_port_interface_types_enum two_port_interface_type;

  constraint reasonable_ports {
    first_port_id inside {[0:(cfg.num_masters-1)]};
    second_port_id inside {[0:(cfg.num_masters-1)]};
    first_port_id != second_port_id;
  }

  constraint valid_two_port_inteface_type {
    if (ace_ports.size() == 0) {
      two_port_interface_type != FIRST_PORT_ACE_SECOND_PORT_ACE;
      two_port_interface_type != FIRST_PORT_ACE_SECOND_PORT_ACE_LITE;
      two_port_interface_type != FIRST_PORT_ACE_LITE_SECOND_PORT_ACE;
    }
    if (ace_lite_ports.size() == 0) {
      two_port_interface_type != FIRST_PORT_ACE_SECOND_PORT_ACE_LITE;
      two_port_interface_type != FIRST_PORT_ACE_LITE_SECOND_PORT_ACE_LITE;
      two_port_interface_type != FIRST_PORT_ACE_LITE_SECOND_PORT_ACE;
    }
    if (ace_ports.size() == 1) {
      two_port_interface_type != FIRST_PORT_ACE_SECOND_PORT_ACE;
    }
    if (ace_lite_ports.size() == 1) {
      two_port_interface_type != FIRST_PORT_ACE_LITE_SECOND_PORT_ACE_LITE;
    }
  } 

  constraint valid_port_id_type {
    if (two_port_interface_type == FIRST_PORT_ACE_SECOND_PORT_ACE) {
      first_port_id inside {ace_ports}; 
      second_port_id inside {ace_ports}; 
    } else if (two_port_interface_type == FIRST_PORT_ACE_SECOND_PORT_ACE_LITE) {
      first_port_id inside {ace_ports}; 
      second_port_id inside {ace_lite_ports}; 
    } else if (two_port_interface_type == FIRST_PORT_ACE_LITE_SECOND_PORT_ACE_LITE) {
      first_port_id inside {ace_lite_ports};
      second_port_id inside {ace_lite_ports};
    } else if (two_port_interface_type == FIRST_AND_SECOND_PORTS_ARE_ACE_OR_ACE_LITE) {
      first_port_id inside {ace_ports,ace_lite_ports};
      second_port_id inside {ace_ports,ace_lite_ports};
    } else if (two_port_interface_type == FIRST_PORT_ACE_LITE_SECOND_PORT_ACE) {
      first_port_id inside {ace_lite_ports};
      second_port_id inside {ace_ports};
    }
  }

  function new(string name = "svt_axi_ace_master_two_port_base_virtual_sequence");
    super.new(name);
  endfunction  
  
  virtual task pre_body();
    bit status, status0, status1;
    super.pre_body();
    raise_phase_objection();

`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
    status0 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_id", first_port_id);
    status1 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_id",second_port_id);
`elsif SVT_OVM_TECHNOLOGY
    status0 = svt_config_int_db#(int unsigned)::get(m_sequencer, , {get_type_name(), ".", "first_port_id"},  first_port_id);
    status1 = svt_config_int_db#(int unsigned)::get(m_sequencer, , {get_type_name(), ".", "second_port_id"}, second_port_id);
    status = svt_config_int_db#(int unsigned)::get(m_sequencer, , {get_type_name(), ".", "sequence_length"},  sequence_length);
`endif
    `svt_xvm_debug("body", $sformatf("first_port_id is 'd%0d as a result of %0s.", first_port_id, status0 ? "config DB" : "randomization"));
    `svt_xvm_debug("body", $sformatf("second_port_id is 'd%0d as a result of %0s.", second_port_id, status1 ? "config DB" : "randomization"));
    
  endtask

  /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

endclass


/**
  * Base class from which all virtual sequences for sequential accesses to overlapping addresses are extended
  */
class svt_axi_ace_master_two_port_base_sequential_virtual_sequence extends svt_axi_ace_master_two_port_base_virtual_sequence;

  typedef enum {
    STORE_OPERATION = 0, /** For ACE: MAKEUNIQUE, CLEANUNIQUE, READUNIQUE, WRITEUNIQUE, WRITELINEUNIQUE. For ACE-Lite: WRITEUNIQUE, WRITELINEUNIQUE */
    LOAD_OPERATION = 1,  /** For ACE: READONCE, READSHARED, READCLEAN, READNOTSHAREDDIRTY. For ACE-Lite: READONCE */
    MEMORY_UPDATE = 2,   /** For ACE: WRITEBACK, WRITECLEAN, WRITEEVICT and EVICT. N/A for ACE-Lite */
    CMO = 3              /** Cache Maintenance Operations: MAKEINVALID, CLEANINVALID and CLEANSHARED */
  } xact_category_enum;


  /** The transaction category for the first port */
  rand xact_category_enum first_port_xact_category;
  
  /** The transaction category for the second port */
  rand xact_category_enum second_port_xact_category;


  /** 
    * Indicates if the weights set by user, support the sequence type
    * Set by derived sequences
    */
  bit is_supported_weights = 0;

  /** 
    * Indicates if the combination of first_port_id and second_port_id are such
    * that there is a common inner shareable or outer shareable domain which
    * can be used for sending transactions with overlapping addresses Set by
    * derived sequences
    */
  bit is_supported_domains = 0;

  constraint solve_port_id_order {
    solve first_port_id before second_port_id;
    solve first_port_id before first_port_xact_category;
    solve second_port_id before second_port_xact_category;
    solve two_port_interface_type before first_port_id;
    solve two_port_interface_type before second_port_id;
  }


  constraint reasonable_xact_category {
    foreach(cfg.master_cfg[i]) {
      if (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::ACE_LITE) {
        if (i == first_port_id) {   
          first_port_xact_category != MEMORY_UPDATE;
        } else if (i == second_port_id) {
          second_port_xact_category != MEMORY_UPDATE;
        }
      }
    }
  }

  function new(string name = "svt_axi_ace_master_two_port_base_sequential_virtual_sequence");
    super.new(name);
  endfunction  

  virtual function bit normalize_weights_based_on_interface_type();
    `svt_fatal("normalize_weights_based_on_interface_type", "This function must be implemented in a derived class");
    return 0;
  endfunction

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    is_supported = 1;
    if (!is_supported_weights || !is_supported_domains) begin
      `svt_xvm_note("is_supported", 
      $sformatf("Either the combination of transaction weights or the absence of a common innershareable or outershareable domain between first_port_id('d%0d) and second_port_id('d%0d) makes it impossible to run this sequence",
      first_port_id,second_port_id));
    end
  endfunction

  /** 
    * Sends a dummy transaction to get the starting address of a sequence 
    * @param init_xact_seq The initialisation sequence which needs to be triggered
    * @param port_id The port on which this sequence should be sent
    * @param supports_both_domains Indicates if both innershareable and outershareable domains can be used
    * @param domain_type If supports_both_domains is not set, indicates the domain_type to be used
    * @param master_xact The master transaction which was sent through init_xact_seq
    */
  virtual task send_dummy_sequence_for_xact_template(svt_axi_ace_master_generic_sequence init_xact_seq,
                                                     int port_id,
                                                     bit supports_both_domains,
                                                     svt_axi_transaction::xact_shareability_domain_enum domain_type,
                                                     output svt_axi_master_transaction master_xact
                                                    );
    svt_axi_cacheline_invalidation init_xact_cacheline_invalidation;
    if (!supports_both_domains) begin
      init_xact_seq.use_directed_domain_type = 1;
      init_xact_seq.directed_domain_type = domain_type;
    end
    init_xact_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    void'(init_xact_seq.randomize with {use_directed_addr == 0;
                                  sequence_length==1;
                                  });
    init_xact_seq.start(p_sequencer.master_sequencer[port_id]);
    // Wait for transactions to finish
    init_xact_seq.wait_for_active_xacts_to_end();
    init_xact_seq.output_xact_mailbox.get(master_xact);
    `svt_xvm_create(init_xact_cacheline_invalidation)
    init_xact_cacheline_invalidation.invalidate_port = port_id;
    init_xact_cacheline_invalidation.invalidate_addr = master_xact.addr;
    init_xact_cacheline_invalidation.start(p_sequencer);
  endtask

  /**
    * If ace_domain_ports provided in the argument has only one port, this method populates
    * the port_id of another ACE port
    * @param master_xact The master transaction that was sent through the initialisation sequence in send_dummy_sequence_for_xact_template
    * @param other_innershareable_ace_port An ACE port which is in the same innershareable domain as the port in ace_domain_ports
    * @param other_outershareable_ace_port An ACE port which is in the same outershareable domain as the port in ace_domain_ports
    * @param peer_port_invalidation_length Indicates the number of cachelines to be invalidated from the new port added to the queue in this method
    * @param ace_domain_ports The ACE domain ports from which the initialisation needs to be done
    */
  virtual function void set_initialisation_ports(svt_axi_master_transaction master_xact,
                                                 int other_innershareable_ace_port,int other_outershareable_ace_port, 
                                                 output int peer_port_invalidation_length,
                                                 ref int ace_domain_ports[$]);


    // If size is 1, it is because 1 port is ACE-Lite. 
    if (ace_domain_ports.size() == 1 && (master_xact.domain_type == svt_axi_transaction::INNERSHAREABLE) && (other_innershareable_ace_port != -1)) begin
      ace_domain_ports.push_back(other_innershareable_ace_port);
      // Since this peer port is now different from the actual port from which we want to initiate transactions,
      // there is no requirement to delete cacheline from it. Basically, this port is just an initialisation port.
      peer_port_invalidation_length = 0;
    end
    else if (ace_domain_ports.size() == 1 && (master_xact.domain_type == svt_axi_transaction::OUTERSHAREABLE) && (other_outershareable_ace_port != -1)) begin
      ace_domain_ports.push_back(other_outershareable_ace_port);
      // Since this peer port is now different from the actual port from which we want to initiate transactions,
      // there is no requirement to delete cacheline from it. Basically, this port is just an initialisation port.
      peer_port_invalidation_length = 0;
    end
  endfunction

  /**
    * Initializes caches when addresses are accessed sequentially
    * MAKEUNIQUE transactions are initiated from init_port_id and READSHARED transactions from peer_port_id.
    * Snoop sequence running on init_port_id must ensure that data is always returned and isshared should also be asserted
    * This is to make sure that cachelines in the ports transition to a shared state which is required for sending a CLEANUNIQUE transaction.
    * Other STORE, LOAD and CMO transactions do not have a specific valid cacheline state requirement that CLEANUNIQUE transactions have. 
    * If peer_port_invalidation_length is not 0, as many cache lines from peer_port_id are invalidated
    * invalidation_mode specifies if invalidation must be from start_addr, or from start_addr + (access_length - peer_port_invalidation_length)
    * If invalidation_mode is 0, invalidation will begin from start_addr; if it is 1, it will beging from the latter.
    */
  virtual task execute_cache_initialization_for_generic_sequential_access(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, int access_length, int peer_port_invalidation_length, 
               int init_port_id, int peer_port_id,int invalidation_mode = 0);
    svt_axi_ace_master_generic_sequence cacheline_init_makeunique_seq, cacheline_init_readshared_seq;
    // Send MAKEUNIQUE on init_port_id and READSHARED on peer_port_id.
    // Snoop transactions should always return data and isshared should be asserted, so 
    // tests which use this sequence must set a factory override for the snoop transactions
    // accordingly
    `svt_xvm_create_on(cacheline_init_makeunique_seq, p_sequencer.master_sequencer[init_port_id]) 
    cacheline_init_makeunique_seq.makeunique_wt = 1;
    cacheline_init_makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    cacheline_init_makeunique_seq.status_start_addr = 1;
    cacheline_init_makeunique_seq.start_addr = start_addr;
    void'(cacheline_init_makeunique_seq.randomize with {use_directed_addr == 0;
                                  sequence_length==access_length;
                                  });
    cacheline_init_makeunique_seq.start(p_sequencer.master_sequencer[init_port_id]);
    // Wait for transactions to finish
    cacheline_init_makeunique_seq.wait_for_active_xacts_to_end();

    `svt_xvm_create_on(cacheline_init_readshared_seq, p_sequencer.master_sequencer[peer_port_id]) 
    cacheline_init_readshared_seq.readshared_wt = 1;
    cacheline_init_readshared_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    cacheline_init_readshared_seq.status_start_addr = 1;
    cacheline_init_readshared_seq.start_addr = start_addr;
    void'(cacheline_init_readshared_seq.randomize with {use_directed_addr == 0;
                                  sequence_length==access_length;
                                  });
    cacheline_init_readshared_seq.start(p_sequencer.master_sequencer[peer_port_id]);
    // Wait for transactions to finish
    cacheline_init_readshared_seq.wait_for_active_xacts_to_end();

    if (peer_port_invalidation_length) begin
      int start_loc = 0;
      if (invalidation_mode == 0) 
        start_loc = 0;
      else
        start_loc = access_length - peer_port_invalidation_length;
      for (int i = 0; i < peer_port_invalidation_length; i++) begin
        svt_axi_cacheline_invalidation   cacheline_invalidation;
        bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] _addr;
        _addr = start_addr + (start_loc+i)*cfg.master_cfg[peer_port_id].cache_line_size;
        `svt_xvm_create(cacheline_invalidation)
        cacheline_invalidation.invalidate_port = peer_port_id;
        cacheline_invalidation.invalidate_addr = _addr;
        cacheline_invalidation.start(p_sequencer);
      end  
    end

  endtask

  /**
    * Initializes caches for load access. It basically initializes memory to some valid value.
    * For ACE ports, if use_writelineunique_for_ace is not set, MAKEUNIQUE transactions followed by WRITEBACK transactions are sent
    * If use_writelineunique_for_ace is set or it is an ACE_LITE port, WRITELINEUNIQUE transactions are sent
    */
  virtual task execute_cache_initialization_for_sequential_load_access(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, int access_length, int init_port_id, bit use_writelineunique_for_ace = 1);
    svt_axi_ace_master_generic_sequence cacheline_init_makeunique_seq, cacheline_init_writelineunique_seq;
    svt_axi_basic_writeclean_full_cacheline cacheline_init_writebackfull_seq;

    if (!use_writelineunique_for_ace && 
        cfg.master_cfg[init_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
      `svt_xvm_create_on(cacheline_init_makeunique_seq, p_sequencer.master_sequencer[init_port_id]) 
      cacheline_init_makeunique_seq.makeunique_wt = 1;
      cacheline_init_makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      cacheline_init_makeunique_seq.status_start_addr = 1;
      cacheline_init_makeunique_seq.start_addr = start_addr;
      void'(cacheline_init_makeunique_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==access_length;
                                    });
      cacheline_init_makeunique_seq.start(p_sequencer.master_sequencer[init_port_id]);
      // Wait for transactions to finish
      cacheline_init_makeunique_seq.wait_for_active_xacts_to_end();
      for (int i = 0; i < access_length; i++) begin
        bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] _addr;
        _addr = start_addr + i*cfg.master_cfg[init_port_id].cache_line_size;
        `svt_xvm_create_on(cacheline_init_writebackfull_seq, p_sequencer.master_sequencer[init_port_id])
        cacheline_init_writebackfull_seq.writeback_wt = 1;
        cacheline_init_writebackfull_seq.directed_addr_mailbox.put(_addr);
        void'(cacheline_init_writebackfull_seq.randomize with {use_directed_addr == 1;sequence_length==1;});
        cacheline_init_writebackfull_seq.start(p_sequencer.master_sequencer[init_port_id]);
        cacheline_init_writebackfull_seq.wait_for_active_xacts_to_end();
      end
    end
    else if (use_writelineunique_for_ace || cfg.master_cfg[init_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      `svt_xvm_create_on(cacheline_init_writelineunique_seq, p_sequencer.master_sequencer[init_port_id]) 
      cacheline_init_writelineunique_seq.writelineunique_wt = 1;
      cacheline_init_writelineunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      cacheline_init_writelineunique_seq.status_start_addr = 1;
      cacheline_init_writelineunique_seq.start_addr = start_addr;
      void'(cacheline_init_writelineunique_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==access_length;
                                    });
      cacheline_init_writelineunique_seq.start(p_sequencer.master_sequencer[init_port_id]);
      // Wait for transactions to finish
      cacheline_init_writelineunique_seq.wait_for_active_xacts_to_end();
    end
  endtask

  /**
    * Initializes cache for memory update transactions such as WRITEBACK, WRITECLEAN, WRITEEVICT and EVICT.
    * Done by sending MAKEUNIQUE transactions.
    * If is_clean is set, then the cachelines are cleaned by sending WRITECLEAN transactions. Clean cachelnes
    * are required to send WRITEEVICT and EVICT transactions
    */
  virtual task execute_cache_initialization_for_memory_update(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, int access_length, int init_port_id, bit is_clean = 0);
     svt_axi_ace_master_generic_sequence cacheline_init_makeunique_seq ;
     svt_axi_basic_writeclean_full_cacheline writecleanfull_seq;
     `svt_xvm_create_on(cacheline_init_makeunique_seq, p_sequencer.master_sequencer[init_port_id]) 
     cacheline_init_makeunique_seq.makeunique_wt = 1;
     cacheline_init_makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_makeunique_seq.status_start_addr = 1;
     cacheline_init_makeunique_seq.start_addr = start_addr;
     void'(cacheline_init_makeunique_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==access_length;
                                   });
     cacheline_init_makeunique_seq.start(p_sequencer.master_sequencer[init_port_id]);
     // Wait for transactions to finish
     cacheline_init_makeunique_seq.wait_for_active_xacts_to_end();
     if (is_clean) begin
       for (int i = 0; i < access_length; i++) begin
         bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] _addr;
         _addr = start_addr + i*cfg.master_cfg[init_port_id].cache_line_size;
         `svt_xvm_create_on(writecleanfull_seq, p_sequencer.master_sequencer[init_port_id])
         writecleanfull_seq.writeclean_wt = 1;
         writecleanfull_seq.directed_addr_mailbox.put(_addr);
         void'(writecleanfull_seq.randomize with {use_directed_addr == 1;sequence_length==1;});
         writecleanfull_seq.start(p_sequencer.master_sequencer[init_port_id]);
         writecleanfull_seq.wait_for_active_xacts_to_end();
       end
     end
  endtask
  
  /**
    * Initializes cache for cmo and store transactions such as CLEANSHARED, MAKEUNIQUE, READUNIQUE, CLEANUNIQUE, WRITEUNIQUE and WRITELINEUNIQUE.
    * If store_select is set, initialization for cached store will be done. ie. MAKEUNIQUE, READUNIQUE, CLEANUNIQUE transctions. 
    * If it is low, initialization for non cached store will be done. ie. WRITEUNIQUE, WRITELINEUNIQUE transactions.
    * Cached store initialization is Done by sending MAKEUNIQUE from init_port_id and READSHARED from peer_port_id.
    * Non-cached store initialization is Done by sending MAKEUNIQUE, WRITECLEANFULL from peer_port_id and READCLEAN from init_port_id.
    * For READUNIQUE, initial state must be INVALID, So for those addresses( from start_addr to (start_addr + (initialization_length* size of the cache line)) )
    * readshared transactions are not sent by calculating the readshared_length.
    */
  virtual task execute_cache_initialization_for_cmo_store(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, int access_length, int init_port_id, int peer_port_id,int initialization_length = 0, bit store_select, bit invalidate_mode);
     svt_axi_ace_master_generic_sequence cacheline_init_makeunique_seq,cacheline_init_writecleanfull_seq;
     svt_axi_ace_master_generic_sequence cacheline_init_readclean_seq, cacheline_init_readshared_seq;
     
     int readshared_length, init_port_invalidation_length;
     
     //If store_select is high, 
     if(store_select) begin  
      readshared_length = access_length - initialization_length;
      init_port_invalidation_length = access_length;
      
     `svt_xvm_create_on(cacheline_init_makeunique_seq, p_sequencer.master_sequencer[init_port_id]) 
     cacheline_init_makeunique_seq.makeunique_wt = 1;
     cacheline_init_makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_makeunique_seq.status_start_addr = 1;
     cacheline_init_makeunique_seq.start_addr = start_addr;
     void'(cacheline_init_makeunique_seq.randomize with {use_directed_addr == 0;
                                   sequence_length== access_length;
                                   });
     cacheline_init_makeunique_seq.start(p_sequencer.master_sequencer[init_port_id]);
     // Wait for transactions to finish
     cacheline_init_makeunique_seq.wait_for_active_xacts_to_end();

    
     `svt_xvm_create_on(cacheline_init_readshared_seq, p_sequencer.master_sequencer[peer_port_id]) 
     cacheline_init_readshared_seq.readshared_wt = 1;
     cacheline_init_readshared_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_readshared_seq.status_start_addr = 1;
     cacheline_init_readshared_seq.start_addr = start_addr + (initialization_length*cfg.master_cfg[peer_port_id].cache_line_size);
     void'(cacheline_init_readshared_seq.randomize with {use_directed_addr == 0;
                                  sequence_length== readshared_length;
                                  });
     cacheline_init_readshared_seq.start(p_sequencer.master_sequencer[peer_port_id]);
     cacheline_init_readshared_seq.wait_for_active_xacts_to_end();

     if(invalidate_mode) begin
      for (int i = 0; i < init_port_invalidation_length; i++) begin
        svt_axi_cacheline_invalidation   cacheline_invalidation;
        bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] _addr;
        _addr = start_addr + (i * cfg.master_cfg[init_port_id].cache_line_size); 
        `svt_xvm_create(cacheline_invalidation)
        cacheline_invalidation.invalidate_port = init_port_id;
        cacheline_invalidation.invalidate_addr = _addr;
        cacheline_invalidation.start(p_sequencer);
      end
     end
     end
     //If store_select is low, 
     else begin
     `svt_xvm_create_on(cacheline_init_makeunique_seq, p_sequencer.master_sequencer[peer_port_id]) 
     cacheline_init_makeunique_seq.makeunique_wt = 1;
     cacheline_init_makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_makeunique_seq.status_start_addr = 1;
     cacheline_init_makeunique_seq.start_addr = start_addr;
     void'(cacheline_init_makeunique_seq.randomize with {use_directed_addr == 0;
                                   sequence_length== access_length;
                                   });
     cacheline_init_makeunique_seq.start(p_sequencer.master_sequencer[peer_port_id]);
     // Wait for transactions to finish
     cacheline_init_makeunique_seq.wait_for_active_xacts_to_end();

     `svt_xvm_create_on(cacheline_init_writecleanfull_seq, p_sequencer.master_sequencer[peer_port_id]) 
     cacheline_init_writecleanfull_seq.writeclean_wt = 1;
     cacheline_init_writecleanfull_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_writecleanfull_seq.status_start_addr = 1;
     cacheline_init_writecleanfull_seq.start_addr = start_addr;
     void'(cacheline_init_writecleanfull_seq.randomize with {use_directed_addr == 0;
                                   sequence_length== access_length;
                                   });
     cacheline_init_writecleanfull_seq.start(p_sequencer.master_sequencer[peer_port_id]);
     // Wait for transactions to finish
     cacheline_init_writecleanfull_seq.wait_for_active_xacts_to_end();
    
    `svt_xvm_create_on(cacheline_init_readclean_seq, p_sequencer.master_sequencer[init_port_id]) 
     cacheline_init_readclean_seq.readclean_wt = 1;
     cacheline_init_readclean_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     cacheline_init_readclean_seq.status_start_addr = 1;
     cacheline_init_readclean_seq.start_addr = start_addr;
     void'(cacheline_init_readclean_seq.randomize with {use_directed_addr == 0;
                                  sequence_length== (access_length / 2);
                                  });
      cacheline_init_readclean_seq.start(p_sequencer.master_sequencer[init_port_id]);
      cacheline_init_readclean_seq.wait_for_active_xacts_to_end();
     
     if(invalidate_mode) begin
      for (int i = 0; i < (access_length / 2); i++) begin
        svt_axi_cacheline_invalidation   cacheline_invalidation;
        bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] _addr;
        _addr = start_addr + (i * cfg.master_cfg[init_port_id].cache_line_size);
        `svt_xvm_create(cacheline_invalidation)
        cacheline_invalidation.invalidate_port = init_port_id;
        cacheline_invalidation.invalidate_addr = _addr;
        cacheline_invalidation.start(p_sequencer);
      end
     end
     end
  endtask

    /**
    * Gets the domain type in which both first_port_id and second_port_id are present
    * If both both ports are in a common INNERSHAREABLE and OUTERSHAREABLE domain then
    * supports_both_domains is set. If there is any other ACE port in the same domain
    * as first_port_id and second_port_id, then other_inner_shareable_ace_port and
    * other_outer_shareable_ace_port are correspondingly set.
    */
  function bit get_domain_type_for_two_port_sequence(int first_port_id, int second_port_id,
                                              output bit supports_both_domains,output svt_axi_transaction::xact_shareability_domain_enum domain_type,
                                              output int other_inner_shareable_ace_port, output int other_outer_shareable_ace_port);
    int ports_in_domain[$],_second_port_in_inner_domain[$],_second_port_in_outer_domain[$];
    other_inner_shareable_ace_port = -1;
    other_outer_shareable_ace_port = -1;
    supports_both_domains = 0;
    get_domain_type_for_two_port_sequence = 1;
    // domain_type, num_ports (0 indicates all ports), is_dvm_enabled, is_only_ace, ports_in_domain
    // Get an innershareable domain in which first_port_id is present and check if second_port_id is part of that doamin
    if (get_random_ports_in_domain(svt_axi_transaction::INNERSHAREABLE,0,0,0,ports_in_domain,first_port_id)) begin
      _second_port_in_inner_domain = ports_in_domain.find() with (item == second_port_id);
      foreach (ports_in_domain[i]) begin
        int _port = ports_in_domain[i];
        if ((_port != first_port_id) && (_port != second_port_id) &&
            (cfg.master_cfg[_port].axi_interface_type == svt_axi_port_configuration::AXI_ACE))
          other_inner_shareable_ace_port = _port;
      end
      ports_in_domain.delete();
    end
    // Get an outershareable domain in which first_port_id is present and check if second_port_id is part of that doamin
    if(get_random_ports_in_domain(svt_axi_transaction::OUTERSHAREABLE,0,0,0,ports_in_domain,first_port_id)) begin
      _second_port_in_outer_domain = ports_in_domain.find() with (item == second_port_id);
      foreach (ports_in_domain[i]) begin
        int _port = ports_in_domain[i];
        if ((_port != first_port_id) && (_port != second_port_id) &&
            (cfg.master_cfg[_port].axi_interface_type == svt_axi_port_configuration::AXI_ACE))
          other_outer_shareable_ace_port = _port;
      end
    end

    if (_second_port_in_inner_domain.size() && _second_port_in_outer_domain.size()) 
      supports_both_domains = 1; 
    else if (_second_port_in_inner_domain.size()) 
      domain_type = svt_axi_transaction::INNERSHAREABLE;
    else if (_second_port_in_outer_domain.size()) 
      domain_type = svt_axi_transaction::OUTERSHAREABLE;
    else begin
      get_domain_type_for_two_port_sequence = 0;
      `svt_xvm_error("get_domain_type_for_two_port_sequence", 
      $sformatf("There is no active(svt_axi_port_configuration::is_active), participating (svt_axi_system_configuration::participating_masters) INNERSHAREABLE or OUTERSHAREABLE domain in which first_port_id('d%0d) and second_port_id('d%0d) are present",
      first_port_id, second_port_id));
    end
  endfunction

  /**
    * Start a sequential CLEANUNIQUE access from start_addr
    */
  task start_sequential_cleanunique_access(svt_axi_ace_master_generic_sequence port_cleanunique_seq, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, 
                                           int port_id, int seq_length, bit use_directed_domain_type, 
                                           svt_axi_transaction::xact_shareability_domain_enum directed_domain_type = svt_axi_transaction::INNERSHAREABLE);
    port_cleanunique_seq.cleanunique_wt = 1;
    if (use_directed_domain_type) begin
      port_cleanunique_seq.use_directed_domain_type = 1;
      port_cleanunique_seq.directed_domain_type = directed_domain_type;
    end
    port_cleanunique_seq.status_start_addr = 1;
    port_cleanunique_seq.start_addr = start_addr;
    port_cleanunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    void'(port_cleanunique_seq.randomize with {use_directed_addr == 0;
                                  sequence_length==seq_length;
                                  });
    port_cleanunique_seq.start(p_sequencer.master_sequencer[port_id]);
  endtask

  /**
    * Start a sequential generic access from start_addr.
    */
  task start_generic_sequential_access(svt_axi_ace_master_generic_sequence port_store_seq, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] start_addr, 
                                           int port_id, int seq_length, bit use_directed_domain_type, 
                                           svt_axi_transaction::xact_shareability_domain_enum directed_domain_type = svt_axi_transaction::INNERSHAREABLE);
    if (use_directed_domain_type) begin
      port_store_seq.use_directed_domain_type = 1;
      port_store_seq.directed_domain_type = directed_domain_type;
    end
    port_store_seq.status_start_addr = 1;
    port_store_seq.start_addr = start_addr;
    port_store_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
    void'(port_store_seq.randomize with {use_directed_addr == 0;
                                  sequence_length==seq_length;
                                  });
    port_store_seq.start(p_sequencer.master_sequencer[port_id]);
  endtask
  
endclass

/**
  * Sends a set of concurrent, sequential store accesses from two ports to the
  * same set of overlapping addresses. The store type transactions can be
  * MAKEUNIQUE, READUNIQUE, CLEANUNIQUE, WRITEUNIQUE or WRITELINEUNIQUE based
  * on the interface types of the ports and the weights.  If
  * first_port_cleanunique_wt or second_port_cleanunique_wt is not zero,
  * cachelines are initialised since CLEANUNIQUE can be sent only from a
  * cacheline in shared state.  Only cachelines from which CLEANUNIQUE needs to
  * be sent are initialized. The number of CLEANUNIQUE transactions sent are
  * determined by the formula sequence_length*cleanunique_wt/(sum of weights of
  * all xact types).  Initialisation is done by sending MAKEUNIQUE transactions
  * from one ACE port and READSHARED transactions from another ACE port to the
  * same set of addresses. Snoop transactions for READSHARED type snoop are
  * programmed (in the corresponding tests) to always assert
  * svt_axi_snoop_transaction::snoop_resp_datatransfer and
  * svt_axi_snoop_transaction::snoop_resp_isshared so that a shared state of
  * the cacheline can be acheived in both masters.  Once cachelines are
  * initialised, sequential stores from first_port_id and second_port_id are
  * made.
  */
class svt_axi_ace_master_two_port_overlapping_addr_store_sequential_sequence extends svt_axi_ace_master_two_port_base_sequential_virtual_sequence;
  
  /** 
    * Bypass cache initialisation. CLEANUNIQUE transactions cannot be sent if
    * cache initialisation is bypassed since CLEANUNIQUE transactions require
    * cache to be in shared state
    */
  bit bypass_cache_initialisation = 0;

  /** Weightage for MAKEUNIQUE store transactions for first_port_id */
  int first_port_makeunique_wt = 1;

  /** Weightage for READUNIQUE store transactions for first_port_id */
  int first_port_readunique_wt = 1;

  /** Weightage for CLEANUNIQUE store transactions for first_port_id */
  int first_port_cleanunique_wt = 1;

  /** Weightage for WRITEUNIQUE store transactions for first_port_id */
  int first_port_writeunique_wt = 0;

  /** Weightage for WRITELINEUNIQUE store transactions for first_port_id */
  int first_port_writelineunique_wt = 0;

  /** Weightage for MAKEUNIQUE store transactions for second_port_id */
  int second_port_makeunique_wt = 1;

  /** Weightage for READUNIQUE store transactions for second_port_id */
  int second_port_readunique_wt = 1;

  /** Weightage for CLEANUNIQUE store transactions for second_port_id */
  int second_port_cleanunique_wt = 1;

  /** Weightage for WRITEUNIQUE store transactions for second_port_id */
  int second_port_writeunique_wt = 0;

  /** Weightage for WRITELINEUNIQUE store transactions for second_port_id */
  int second_port_writelineunique_wt = 0;

  constraint reasonable_supported_xact_category {
    first_port_xact_category == STORE_OPERATION;
    second_port_xact_category == STORE_OPERATION;
  } 

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_two_port_overlapping_addr_store_sequential_sequence)
    
  function new(string name = "svt_axi_ace_master_two_port_overlapping_addr_store_sequential_sequence");
    super.new(name);
  endfunction

  virtual task body();
    svt_axi_master_transaction _master_xact;
    svt_axi_ace_master_generic_sequence init_xact_seq;
    svt_axi_ace_master_generic_sequence main_cleanunique_store_seq, peer_cleanunique_store_seq;
    svt_axi_ace_master_generic_sequence main_other_store_seq, peer_other_store_seq;
    int store_port_id, peer_port_id;
    svt_axi_transaction::xact_shareability_domain_enum _domain_type;
    bit supports_both_domains = 0;
    bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] main_store_start_addr, peer_store_start_addr;
    int _makeunique_wt, _cleanunique_wt, _readunique_wt, _writeunique_wt, _writelineunique_wt;
    int initialisation_length, peer_port_invalidation_length, ace_domain_ports[$];
    bit disable_cleanunique_store_access = 0;
    int other_innershareable_ace_port, other_outershareable_ace_port;
    int store_port_cleanunique_length, peer_port_cleanunique_length;
    bit status;
    super.body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_makeunique_wt",first_port_makeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readunique_wt",first_port_readunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleanunique_wt",first_port_cleanunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_writeunique_wt",first_port_writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_writelineunique_wt",first_port_writelineunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_makeunique_wt",second_port_makeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readunique_wt",second_port_readunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_cleanunique_wt",second_port_cleanunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_writeunique_wt",second_port_writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_writelineunique_wt",second_port_writelineunique_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "bypass_cache_initialisation",bypass_cache_initialisation);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_makeunique_wt"}, first_port_makeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readunique_wt"}, first_port_readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleanunique_wt"}, first_port_cleanunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_writeunique_wt"}, first_port_writeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_writelineunique_wt"}, first_port_writelineunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_makeunique_wt"}, second_port_makeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readunique_wt"}, second_port_readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_cleanunique_wt"}, second_port_cleanunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_writeunique_wt"}, second_port_writeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".bypass_cache_initialisation"}, bypass_cache_initialisation);
`endif
    disable_cleanunique_store_access = 1;
    is_supported_weights = normalize_weights_based_on_interface_type();
    is_supported_domains = get_domain_type_for_two_port_sequence(first_port_id,second_port_id,supports_both_domains,_domain_type,other_innershareable_ace_port,other_outershareable_ace_port);
    `svt_xvm_note("body", $sformatf("sequence_length = 'd%0d. first_port_id = 'd%0d. second_port_id = 'd%0d. bypass_cache_initialisation = 'b%0b", 
      sequence_length, first_port_id, second_port_id, bypass_cache_initialisation));
    if (!is_supported(cfg))
      return;
    // If both ports are ACE-Lite, no need for cache initialisation because ACE-Lite does not send CLEANUNIQUE
    if (
         (
           (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) && 
           (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) 
         ) 
       ) begin
      bypass_cache_initialisation = 1;
      `svt_xvm_debug("body", "Bypassing cache initialisation since both first_port_id and second_port_id are ACE_LITE ports");
    end
    // If any of the two ports is ACE_LITE and there are no other ACE ports in the domain of these two ports,
    // then initialisation for cleanunique need not be done because cacheline will not be in shared state.
    else if (
         (
           (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) ||
           (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) 
         ) &&
         ((other_innershareable_ace_port == -1) && (other_outershareable_ace_port == -1))
       ) begin
      bypass_cache_initialisation = 1;
      `svt_xvm_debug("body", "Bypassing cache initialisation since either of first_port_id and second_port_id is an ACE_LITE port and there are no other ACE ports in relevant domain");
    end
    // Set default values for weights in initialised transaction (init_xact_seq)
    _makeunique_wt = first_port_makeunique_wt;
    _cleanunique_wt = first_port_cleanunique_wt;
    _readunique_wt = first_port_readunique_wt;
    _writeunique_wt = first_port_writeunique_wt;
    _writelineunique_wt = first_port_writelineunique_wt;

    // By default put ACE ports in initialisation ports.
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(first_port_id);
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(second_port_id);
    store_port_id = first_port_id;
    peer_port_id = second_port_id;

    if ((cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) && 
        (first_port_xact_category == STORE_OPERATION) && (first_port_cleanunique_wt != 0) && !bypass_cache_initialisation) begin
      store_port_id = first_port_id;
      peer_port_id = second_port_id;
      initialisation_length = sequence_length * first_port_cleanunique_wt/(first_port_makeunique_wt + first_port_cleanunique_wt + first_port_readunique_wt + first_port_writeunique_wt + first_port_writelineunique_wt);
      // The CLEANUNIQUE transaction needs to have overlapped access with READUNIQUE and MAKEUNIQUE as well. So
      // we need cachelines to be in shared state only for those lines from which CLEANUNIQUE is sent. For the 
      // rest of the cachelines, invalidate them, so that we can send READUNIQUE and MAKEUNIQUE.
      peer_port_invalidation_length = initialisation_length * (second_port_makeunique_wt + second_port_readunique_wt + second_port_writeunique_wt + second_port_writelineunique_wt)/(second_port_makeunique_wt + second_port_cleanunique_wt + second_port_readunique_wt + second_port_writeunique_wt + second_port_writelineunique_wt);
      disable_cleanunique_store_access = 0;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. initialisation_length = 'd%0d. peer_port_invalidation_length = 'd%0d", 
      sequence_length, initialisation_length, peer_port_invalidation_length));
    end
    if ((cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) && 
             (second_port_xact_category == STORE_OPERATION) && (second_port_cleanunique_wt != 0) && !bypass_cache_initialisation) begin
      // Override store_port_id if the weightage for cleanunique (which requires initialisation) is 
      // is more for second port.
      if (second_port_cleanunique_wt > first_port_cleanunique_wt) begin
        // The first port is considered the "store port". This is the port from which the most number
        // of CLEANUNIQUE transactions are sent. If the second port is the "store port", then reverse
        // the order in ace_domain_ports so that initialisation takes this into account
        if (ace_domain_ports.size() == 2) begin
          ace_domain_ports.delete();
          ace_domain_ports.push_back(second_port_id);
          ace_domain_ports.push_back(first_port_id);
        end

        store_port_id = second_port_id;
        peer_port_id = first_port_id;
        _makeunique_wt = second_port_makeunique_wt;
        _cleanunique_wt = second_port_cleanunique_wt;
        _readunique_wt = second_port_readunique_wt;
        _writeunique_wt = second_port_writeunique_wt;
        _writelineunique_wt = second_port_writelineunique_wt;
        initialisation_length = sequence_length * second_port_cleanunique_wt/(second_port_makeunique_wt + second_port_cleanunique_wt + second_port_readunique_wt+ second_port_writeunique_wt + second_port_writelineunique_wt);
        peer_port_invalidation_length = initialisation_length * (first_port_makeunique_wt + first_port_readunique_wt+ first_port_writeunique_wt + first_port_writelineunique_wt)/(first_port_makeunique_wt + first_port_cleanunique_wt + first_port_readunique_wt+ first_port_writeunique_wt + first_port_writelineunique_wt);
      `svt_xvm_debug("body", $sformatf("Overridden values based on second_port_id parameters: sequence_length = 'd%0d. initialisation_length = 'd%0d. peer_port_invalidation_length = 'd%0d", 
      sequence_length, initialisation_length, peer_port_invalidation_length));
      end
      disable_cleanunique_store_access = 0;
    end

    // Generate only one transaction so that we get a reference to the starting address
    // which in turn can be used for initialisation.
    `svt_xvm_create_on(init_xact_seq, p_sequencer.master_sequencer[store_port_id]) 
    init_xact_seq.makeunique_wt = _makeunique_wt;
    init_xact_seq.readunique_wt = _readunique_wt;
    init_xact_seq.cleanunique_wt = _cleanunique_wt;
    init_xact_seq.writeunique_wt = _writeunique_wt;
    init_xact_seq.writelineunique_wt = _writelineunique_wt;
    send_dummy_sequence_for_xact_template(init_xact_seq,store_port_id,supports_both_domains,_domain_type,_master_xact);
    if (!bypass_cache_initialisation && !disable_cleanunique_store_access && (initialisation_length != 0) ) begin 
      string _ace_ports_str = "";
      if (ace_domain_ports.size() == 1)
        set_initialisation_ports(_master_xact,other_innershareable_ace_port,other_outershareable_ace_port,peer_port_invalidation_length,ace_domain_ports);
     
      foreach (ace_domain_ports[i]) begin
        _ace_ports_str = $sformatf("'d%0d ", ace_domain_ports[i]);
      end
      `svt_xvm_debug("body", $sformatf("ace_domain_ports: %s", _ace_ports_str));

      if (ace_domain_ports.size() == 1)
        bypass_cache_initialisation = 1;
      else
        execute_cache_initialization_for_generic_sequential_access(_master_xact.cacheline_addr(),initialisation_length,peer_port_invalidation_length,ace_domain_ports[0],ace_domain_ports[1],1);
    end

    // CLEANUNIQUE can be sent only if cache is initialised to some shared
    // state or svt_axi_port_configuration::speculative_read_enable is set.
    if (cfg.master_cfg[store_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      store_port_cleanunique_length = initialisation_length;
    if (cfg.master_cfg[peer_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      peer_port_cleanunique_length = initialisation_length-peer_port_invalidation_length;
    `svt_xvm_debug("body", $sformatf("disable_cleanunique_store_access = 'b%0b. bypass_cache_initialisation = 'b%0b. store_port_cleanunique_length = 'd%0d. peer_port_cleanunique_length = 'd%0d",
    disable_cleanunique_store_access,bypass_cache_initialisation,store_port_cleanunique_length,peer_port_cleanunique_length));
    `svt_xvm_debug("body",$sformatf("start addr = 'h%0x. store_port_id = 'd%0d. peer_port_id = 'd%0d. supports_both_domains = 'b%0b. directed_domain_type = %0s",
    init_xact_seq.start_addr,store_port_id,peer_port_id,supports_both_domains,init_xact_seq.directed_domain_type.name()));
    `svt_xvm_create_on(main_other_store_seq, p_sequencer.master_sequencer[store_port_id]) 
    `svt_xvm_create_on(peer_other_store_seq, p_sequencer.master_sequencer[peer_port_id])

    if (store_port_id == first_port_id) begin
      main_other_store_seq.makeunique_wt = first_port_makeunique_wt; 
      main_other_store_seq.readunique_wt = first_port_readunique_wt; 
      main_other_store_seq.writeunique_wt = first_port_writeunique_wt; 
      main_other_store_seq.writelineunique_wt = first_port_writelineunique_wt; 
      peer_other_store_seq.makeunique_wt = second_port_makeunique_wt; 
      peer_other_store_seq.readunique_wt = second_port_readunique_wt; 
      peer_other_store_seq.writeunique_wt = second_port_writeunique_wt; 
      peer_other_store_seq.writelineunique_wt = second_port_writelineunique_wt; 
    end
    else begin
      main_other_store_seq.makeunique_wt = second_port_makeunique_wt; 
      main_other_store_seq.readunique_wt = second_port_readunique_wt; 
      main_other_store_seq.writeunique_wt = second_port_writeunique_wt; 
      main_other_store_seq.writelineunique_wt = second_port_writelineunique_wt; 
      peer_other_store_seq.makeunique_wt = first_port_makeunique_wt; 
      peer_other_store_seq.readunique_wt = first_port_readunique_wt; 
      peer_other_store_seq.writeunique_wt = first_port_writeunique_wt; 
      peer_other_store_seq.writelineunique_wt = first_port_writelineunique_wt; 
    end
    main_store_start_addr = init_xact_seq.start_addr + store_port_cleanunique_length*cfg.master_cfg[store_port_id].cache_line_size;
    peer_store_start_addr = init_xact_seq.start_addr + peer_port_cleanunique_length*cfg.master_cfg[peer_port_id].cache_line_size;
    `svt_xvm_debug("body", $sformatf("main_store_start_addr = 'h%0x. peer_store_start_addr = 'h%0x",main_store_start_addr,peer_store_start_addr));
    // Initiate CLEANUNIQUE from both ports.
    fork
    begin
      if (
          !disable_cleanunique_store_access && (store_port_cleanunique_length != 0) && (initialisation_length != 0) &&
          (!bypass_cache_initialisation ||
           (cfg.master_cfg[store_port_id].speculative_read_enable)
          )
         ) begin
         `svt_xvm_create_on(main_cleanunique_store_seq, p_sequencer.master_sequencer[store_port_id]) 
          start_sequential_cleanunique_access(main_cleanunique_store_seq,init_xact_seq.start_addr,store_port_id,store_port_cleanunique_length,!supports_both_domains,init_xact_seq.directed_domain_type);
        end
        start_generic_sequential_access(main_other_store_seq,main_store_start_addr,
                                        store_port_id, (sequence_length-initialisation_length),
                                        !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    begin
      if (
          !disable_cleanunique_store_access && (peer_port_cleanunique_length != 0) && (initialisation_length != 0) &&
          (!bypass_cache_initialisation ||
           (cfg.master_cfg[peer_port_id].speculative_read_enable)
          )
         ) begin
        `svt_xvm_create_on(peer_cleanunique_store_seq, p_sequencer.master_sequencer[peer_port_id]) 
        start_sequential_cleanunique_access(peer_cleanunique_store_seq,init_xact_seq.start_addr,peer_port_id,peer_port_cleanunique_length,!supports_both_domains,init_xact_seq.directed_domain_type);
      end
      start_generic_sequential_access(peer_other_store_seq,peer_store_start_addr,
                                      peer_port_id, (sequence_length-peer_port_cleanunique_length),
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    join

    if (main_cleanunique_store_seq != null)
      main_cleanunique_store_seq.wait_for_active_xacts_to_end();
    if (peer_cleanunique_store_seq != null)
      peer_cleanunique_store_seq.wait_for_active_xacts_to_end();
    if (main_other_store_seq != null)
      main_other_store_seq.wait_for_active_xacts_to_end();
    if (peer_other_store_seq != null)
      peer_other_store_seq.wait_for_active_xacts_to_end();

  endtask

  virtual function bit normalize_weights_based_on_interface_type();
    normalize_weights_based_on_interface_type = 1;
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      first_port_makeunique_wt = 0; 
      first_port_readunique_wt = 0;
      first_port_cleanunique_wt = 0;
    end
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      second_port_makeunique_wt = 0; 
      second_port_readunique_wt = 0;
      second_port_cleanunique_wt = 0;
    end
    if ((first_port_makeunique_wt + first_port_readunique_wt + first_port_cleanunique_wt + first_port_writeunique_wt + first_port_writelineunique_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for store transactions in first_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", first_port_id));
    end
    if ((second_port_makeunique_wt + second_port_readunique_wt + second_port_cleanunique_wt + second_port_writeunique_wt + second_port_writelineunique_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for store transactions in second_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", second_port_id));
    end
    if (bypass_cache_initialisation) begin
      first_port_cleanunique_wt = 0;
      second_port_cleanunique_wt = 0;
    end
  endfunction


endclass

/**
  * Sends a set of concurrent, sequential load or cmo accesses from first_port_id and
  * load or cmo accesses from second_port_id based on the interface types of the 
  * ports and the weights selected from corresponding tests to the same set 
  * of overlapping addresses. Load type transactions can be READONCE, READCLEAN, READSHARED
  * or READNOTSHAREDDIRTY. cmo type transactions can be MAKEINVALID, CLEANINVALID
  * and CLEANSHARED. Prior to sending the load transaction an
  * initialisation procedure is invoked based on the following sequence, unless
  * bypass_cache_initialisation is set:
  * - In order that the load transactions return some valid data,
  * incase of ACE port MAKEUNIQUE followed by WRITEBACK are sent to update memory. 
  * incase of ACE_LITE port WRITELINEUNIQUE transactions are sent to update memory.  
  * .
  * After this initialisation, sequential load or sequential cmo from first_port_id and
  * sequential load or sequential cmo from second_port_id are sent concurrently to the same 
  * set of addresses.
  */
class svt_axi_ace_master_two_port_overlapping_addr_load_cmo_sequential_sequence extends svt_axi_ace_master_two_port_base_sequential_virtual_sequence;
  
  /** 
    * Bypass cache initialisation.If set, the initialization for load transactions
    * will not be initiated.
    */
  bit bypass_cache_initialisation = 0;

  /** Weightage for READSHARED load transactions for first_port_id */
  int first_port_readshared_wt = 1;

  /** Weightage for READNOTSHAREDDIRTY load transactions for first_port_id */
  int first_port_readnotshareddirty_wt = 1;

  /** Weightage for READCLEAN load transactions for first_port_id */
  int first_port_readclean_wt = 1;

  /** Weightage for READONCE load transactions for first_port_id */
  int first_port_readonce_wt = 1;
  
  /** Weightage for MAKEINVALID CMO transactions for first_port_id */
  int first_port_makeinvalid_wt = 1;
  
  /** Weightage for CLEANSHARED CMO transactions for first_port_id */
  int first_port_cleanshared_wt = 1;
  
  /** Weightage for CLEANSHAREDPERSIST CMO transactions for first_port_id */
  int first_port_cleansharedpersist_wt = 1;

  /** Weightage for CLEANINVALID CMO transactions for first_port_id */
  int first_port_cleaninvalid_wt = 1;

  /** Weightage for READSHARED load transactions for second_port_id */
  int second_port_readshared_wt = 1;

  /** Weightage for READNOTSHAREDDIRTY load transactions for second_port_id */
  int second_port_readnotshareddirty_wt = 1;

  /** Weightage for READCLEAN load transactions for second_port_id */
  int second_port_readclean_wt = 1;

  /** Weightage for READONCE load transactions for second_port_id */
  int second_port_readonce_wt = 1;
  
  /** Weightage for MAKEINAVLID CMO transactions for second_port_id */
  int second_port_makeinvalid_wt = 1;
  
  /** Weightage for CLEANSHARED CMO transactions for second_port_id */
  int second_port_cleanshared_wt = 1;
  
  /** Weightage for CLEANSHAREDPERSIST CMO transactions for second_port_id */
  int second_port_cleansharedpersist_wt = 1;
  
  /** Weightage for CLEANINVALID CMO transactions for second_port_id */
  int second_port_cleaninvalid_wt = 1;

  constraint reasonable_supported_xact_category {
    first_port_xact_category inside {LOAD_OPERATION,CMO};
    second_port_xact_category inside {LOAD_OPERATION,CMO};
  } 

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_two_port_overlapping_addr_load_cmo_sequential_sequence)
    
  function new(string name = "svt_axi_ace_master_two_port_overlapping_addr_load_cmo_sequential_sequence");
    super.new(name);
  endfunction

  virtual task body();
    svt_axi_master_transaction _master_xact;
    svt_axi_ace_master_generic_sequence init_xact_seq;
    svt_axi_ace_master_generic_sequence first_port_load_seq, second_port_load_seq;
    svt_axi_transaction::xact_shareability_domain_enum _domain_type;
    bit supports_both_domains = 0;
    int initialisation_length, peer_port_invalidation_length, ace_domain_ports[$];
    int other_innershareable_ace_port, other_outershareable_ace_port;
    bit status;
    bit is_supported_xacts = 0;
    super.body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readshared_wt",first_port_readshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readnotshareddirty_wt",first_port_readnotshareddirty_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readclean_wt",first_port_readclean_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readonce_wt",first_port_readonce_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_makeinvalid_wt",first_port_makeinvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleanshared_wt",first_port_cleanshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleansharedpersist_wt",first_port_cleansharedpersist_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleaninvalid_wt",first_port_cleaninvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readshared_wt",second_port_readshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readnotshareddirty_wt",second_port_readnotshareddirty_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readclean_wt",second_port_readclean_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readonce_wt",second_port_readonce_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_makeinvalid_wt",second_port_makeinvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_cleanshared_wt",second_port_cleanshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_cleansharedpersist_wt",second_port_cleansharedpersist_wt);    
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_cleaninvalid_wt",second_port_cleaninvalid_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "bypass_cache_initialisation",bypass_cache_initialisation);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readshared_wt"}, first_port_readshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readnotshareddirty_wt"}, first_port_readnotshareddirty_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readclean_wt"}, first_port_readclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readonce_wt"}, first_port_readonce_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_makeinvalid_wt"}, first_port_makeinvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleanshared_wt"}, first_port_cleanshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleansharedpersist_wt"}, first_port_cleansharedpersist_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleaninvalid_wt"}, first_port_cleaninvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readshared_wt"}, second_port_readshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readnotshareddirty_wt"}, second_port_readnotshareddirty_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readclean_wt"}, second_port_readclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readonce_wt"}, second_port_readonce_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_makeinvalid_wt"}, second_port_makeinvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_cleanshared_wt"}, second_port_cleanshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_cleansharedpersist_wt"}, second_port_cleansharedpersist_wt);    
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_cleaninvalid_wt"}, second_port_cleaninvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".bypass_cache_initialisation"}, bypass_cache_initialisation);
`endif
    is_supported_xacts = normalize_weights_based_on_xact_category();
    is_supported_weights = normalize_weights_based_on_interface_type();
    is_supported_domains = get_domain_type_for_two_port_sequence(first_port_id,second_port_id,supports_both_domains,_domain_type,other_innershareable_ace_port,other_outershareable_ace_port);
    `svt_xvm_note("body", $sformatf("sequence_length = 'd%0d. first_port_id = 'd%0d. second_port_id = 'd%0d. bypass_cache_initialisation = 'b%0b", 
      sequence_length, first_port_id, second_port_id, bypass_cache_initialisation));
    if (!is_supported(cfg))
      return;
    initialisation_length = sequence_length;

    // Generate only one transaction so that we get a reference to the starting address
    // which in turn can be used for initialisation.
    `svt_xvm_create_on(init_xact_seq, p_sequencer.master_sequencer[first_port_id]) 
    init_xact_seq.readshared_wt = first_port_readshared_wt; 
    init_xact_seq.readnotshareddirty_wt = first_port_readnotshareddirty_wt; 
    init_xact_seq.readclean_wt = first_port_readclean_wt; 
    init_xact_seq.readonce_wt = first_port_readonce_wt; 
    init_xact_seq.makeinvalid_wt = first_port_makeinvalid_wt; 
    init_xact_seq.cleanshared_wt = first_port_cleanshared_wt;
    init_xact_seq.cleansharedpersist_wt = first_port_cleansharedpersist_wt;
    init_xact_seq.cleaninvalid_wt = first_port_cleaninvalid_wt;
    init_xact_seq.generate_only_shareable_domain = 1;

    send_dummy_sequence_for_xact_template(init_xact_seq,first_port_id,supports_both_domains,_domain_type,_master_xact);
    `svt_xvm_debug("body",$sformatf("first_port_id='d%0d. second_port_id='d%0d. supports_both_domains='b%0b. domain_type=%s. initialisation_length='d%0d. bypass_cache_initialisation='b%0b",
    first_port_id,second_port_id,supports_both_domains,_domain_type.name(),initialisation_length,bypass_cache_initialisation));
    if (!bypass_cache_initialisation && (initialisation_length != 0) ) begin 
      ace_domain_ports.push_back(first_port_id);
      ace_domain_ports.push_back(second_port_id);
      execute_cache_initialization_for_sequential_load_access(_master_xact.cacheline_addr(), initialisation_length, ace_domain_ports[0]);
    end

    `svt_xvm_create_on(first_port_load_seq, p_sequencer.master_sequencer[first_port_id]) 
    `svt_xvm_create_on(second_port_load_seq, p_sequencer.master_sequencer[second_port_id])

    first_port_load_seq.readshared_wt = first_port_readshared_wt; 
    first_port_load_seq.readnotshareddirty_wt = first_port_readnotshareddirty_wt; 
    first_port_load_seq.readclean_wt = first_port_readclean_wt; 
    first_port_load_seq.readonce_wt = first_port_readonce_wt; 
    first_port_load_seq.makeinvalid_wt = first_port_makeinvalid_wt; 
    first_port_load_seq.cleanshared_wt = first_port_cleanshared_wt;
    first_port_load_seq.cleansharedpersist_wt = first_port_cleansharedpersist_wt;
    first_port_load_seq.cleaninvalid_wt = first_port_cleaninvalid_wt;
    
    second_port_load_seq.readshared_wt = second_port_readshared_wt; 
    second_port_load_seq.readnotshareddirty_wt = second_port_readnotshareddirty_wt; 
    second_port_load_seq.readclean_wt = second_port_readclean_wt; 
    second_port_load_seq.readonce_wt = second_port_readonce_wt; 
    second_port_load_seq.makeinvalid_wt = second_port_makeinvalid_wt; 
    second_port_load_seq.cleanshared_wt = second_port_cleanshared_wt;
    second_port_load_seq.cleansharedpersist_wt = second_port_cleansharedpersist_wt;
    second_port_load_seq.cleaninvalid_wt = second_port_cleaninvalid_wt; 

    fork
    begin
      start_generic_sequential_access(first_port_load_seq,_master_xact.cacheline_addr(),
                                      first_port_id, sequence_length,
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    begin
      start_generic_sequential_access(second_port_load_seq,_master_xact.cacheline_addr(),
                                      second_port_id, sequence_length,
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    join
    first_port_load_seq.wait_for_active_xacts_to_end();
    second_port_load_seq.wait_for_active_xacts_to_end();
  endtask
  
  // This function will normalize the weights according to the transaction 
  // category selected.
  function bit normalize_weights_based_on_xact_category();
    normalize_weights_based_on_xact_category = 1;
    if(first_port_xact_category == LOAD_OPERATION) begin
      first_port_makeinvalid_wt = 0;
      first_port_cleanshared_wt = 0;
      first_port_cleansharedpersist_wt = 0;
      first_port_cleaninvalid_wt = 0;
    end
    else if(first_port_xact_category == CMO) begin
      first_port_readshared_wt = 0;
      first_port_readnotshareddirty_wt = 0;
      first_port_readclean_wt = 0;
      first_port_readonce_wt = 0;
    end

    if(second_port_xact_category == LOAD_OPERATION) begin
      second_port_makeinvalid_wt = 0;
      second_port_cleanshared_wt = 0;
      second_port_cleansharedpersist_wt = 0;
      second_port_cleaninvalid_wt = 0;
    end
    else if(second_port_xact_category == CMO) begin
      second_port_readshared_wt = 0;
      second_port_readnotshareddirty_wt = 0;
      second_port_readclean_wt = 0;
      second_port_readonce_wt = 0;
    end

    if ((first_port_readshared_wt + first_port_readnotshareddirty_wt + first_port_readclean_wt + first_port_readonce_wt + first_port_makeinvalid_wt + first_port_cleanshared_wt + first_port_cleansharedpersist_wt + first_port_cleaninvalid_wt) == 0) begin
      normalize_weights_based_on_xact_category = 0;
      `svt_xvm_error("normalize_weights_based_on_xact_category", $sformatf("The sum of all the valid weights for load & CMO transactions in first_port_id('d%0d) after normalizing for transaction type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent is non-zero", first_port_id));
    end
    if ((second_port_readshared_wt + second_port_readnotshareddirty_wt + second_port_readclean_wt + second_port_readonce_wt + second_port_makeinvalid_wt + second_port_cleanshared_wt + second_port_cleansharedpersist_wt + second_port_cleaninvalid_wt) == 0) begin
      normalize_weights_based_on_xact_category = 0;
      `svt_xvm_error("normalize_weights_based_on_xact_category", $sformatf("The sum of all the valid weights for load & CMO transactions in second_port_id('d%0d) after normalizing for transaction type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent is non-zero", second_port_id));
    end
  endfunction
  
  // This function will normalize the weights according to the interface 
  // type selected.
  virtual function bit normalize_weights_based_on_interface_type();
    normalize_weights_based_on_interface_type = 1;
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      first_port_readshared_wt = 0;
      first_port_readnotshareddirty_wt = 0;
      first_port_readclean_wt = 0;
    end
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      second_port_readshared_wt = 0;
      second_port_readnotshareddirty_wt = 0;
      second_port_readclean_wt = 0;
    end
    if ((first_port_readshared_wt + first_port_readnotshareddirty_wt + first_port_readclean_wt + first_port_readonce_wt + first_port_makeinvalid_wt + first_port_cleanshared_wt + first_port_cleansharedpersist_wt + first_port_cleaninvalid_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for load & CMO transactions in first_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", first_port_id));
    end
    if ((second_port_readshared_wt + second_port_readnotshareddirty_wt + second_port_readclean_wt + second_port_readonce_wt + second_port_makeinvalid_wt + second_port_cleanshared_wt + second_port_cleansharedpersist_wt + second_port_cleaninvalid_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for load & CMO transactions in second_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", second_port_id));
    end
  endfunction
endclass


/**
  * Sends a set of concurrent, sequential store accesses from first_port_id and load
  * accesses from second_port_id to the same set of overlapping addresses. The
  * store type transactions can be MAKEUNIQUE, READUNIQUE, CLEANUNIQUE,
  * WRITEUNIQUE or WRITELINEUNIQUE based on the interface types of the ports
  * and the weights.  Load type transactions can be READONCE, READCLEAN,
  * READSHARED or READNOTSHAREDDIRTY. Prior to sending the store and load transaction
  * an initialisation procedure is invoked based on the following sequence, unless
  * bypass_cache_initialisation is set:
  * - In order that the load transactions return some valid data,
  * WRITELINEUNIQUE transactions are sent to update memory.  
  * .
  * - If first_port_cleanunique_wt is not zero, cachelines are
  * initialised, since CLEANUNIQUE can be sent only from a cacheline in shared
  * state. Only cachelines from which CLEANUNIQUE needs to be sent are
  * initialized. The number of CLEANUNIQUE transactions sent are determined by
  * the formula sequence_length*first_port_cleanunique_wt/(sum of weights of
  * all xact types in first port).  Initialisation is done by sending
  * MAKEUNIQUE transactions from one ACE port and READSHARED transactions from
  * another ACE port to the same set of addresses. Snoop transactions for
  * READSHARED type snoop are programmed (in the corresponding tests) to always
  * assert svt_axi_snoop_transaction::snoop_resp_datatransfer and
  * svt_axi_snoop_transaction::snoop_resp_isshared so that a shared state of
  * the cacheline can be acheived in both masters.  All shared cachelines in
  * second_port_id are invalidated so that the load transactions can be sent on
  * the interface.  
  * .
  * After this initialisation, sequential stores from first_port_id and
  * sequential loads from second_port_id are sent.
  */
class svt_axi_ace_master_two_port_overlapping_addr_store_and_load_sequential_sequence extends svt_axi_ace_master_two_port_base_sequential_virtual_sequence;
  
  /** 
    * Bypass cache initialisation. CLEANUNIQUE transactions cannot be sent if
    * cache initialisation is bypassed since CLEANUNIQUE transactions require
    * cache to be in shared state
    */
  bit bypass_cache_initialisation = 0;

  /** Weightage for MAKEUNIQUE store transactions for first_port_id */
  int first_port_makeunique_wt = 1;

  /** Weightage for READUNIQUE store transactions for first_port_id */
  int first_port_readunique_wt = 1;

  /** Weightage for CLEANUNIQUE store transactions for first_port_id */
  int first_port_cleanunique_wt = 1;

  /** Weightage for WRITEUNIQUE store transactions for first_port_id */
  int first_port_writeunique_wt = 0;

  /** Weightage for WRITELINEUNIQUE store transactions for first_port_id */
  int first_port_writelineunique_wt = 0;

  /** Weightage for READSHARED store transactions for second_port_id */
  int second_port_readshared_wt = 1;

  /** Weightage for READNOTSHAREDDIRTY store transactions for second_port_id */
  int second_port_readnotshareddirty_wt = 1;

  /** Weightage for READCLEAN store transactions for second_port_id */
  int second_port_readclean_wt = 1;

  /** Weightage for READONCE store transactions for second_port_id */
  int second_port_readonce_wt = 1;

  constraint reasonable_supported_xact_category {
    first_port_xact_category == STORE_OPERATION;
    second_port_xact_category == LOAD_OPERATION;
  } 

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_two_port_overlapping_addr_store_and_load_sequential_sequence)
    
  function new(string name = "svt_axi_ace_master_two_port_overlapping_addr_store_and_load_sequential_sequence");
    super.new(name);
  endfunction

  virtual task body();
    svt_axi_master_transaction _master_xact;
    svt_axi_ace_master_generic_sequence init_xact_seq;
    svt_axi_ace_master_generic_sequence first_port_cleanunique_store_seq, first_port_non_cleanunique_store_seq, second_port_load_seq;
    svt_axi_transaction::xact_shareability_domain_enum _domain_type;
    bit supports_both_domains = 0;
    int initialisation_length, peer_port_invalidation_length, ace_domain_ports[$];
    bit disable_cleanunique_store_access = 0;
    int other_innershareable_ace_port, other_outershareable_ace_port;
    int store_port_cleanunique_length;
    bit bypass_cleanunique_cache_initialisation = 0;
    bit status;
    super.body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_makeunique_wt",first_port_makeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_readunique_wt",first_port_readunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleanunique_wt",first_port_cleanunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_writeunique_wt",first_port_writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_writelineunique_wt",first_port_writelineunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readshared_wt",second_port_readshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readnotshareddirty_wt",second_port_readnotshareddirty_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readclean_wt",second_port_readclean_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readonce_wt",second_port_readonce_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "bypass_cache_initialisation",bypass_cache_initialisation);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_makeunique_wt"}, first_port_makeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_readunique_wt"}, first_port_readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleanunique_wt"}, first_port_cleanunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_writeunique_wt"}, first_port_writeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_writelineunique_wt"}, first_port_writelineunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readshared_wt"}, second_port_readshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readnotshareddirty_wt"}, second_port_readnotshareddirty_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readclean_wt"}, second_port_readclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readonce_wt"}, second_port_readonce_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".bypass_cache_initialisation"}, bypass_cache_initialisation);
`endif
    disable_cleanunique_store_access = 1;
    is_supported_weights = normalize_weights_based_on_interface_type();
    is_supported_domains = get_domain_type_for_two_port_sequence(first_port_id,second_port_id,supports_both_domains,_domain_type,other_innershareable_ace_port,other_outershareable_ace_port);
    `svt_xvm_note("body", $sformatf("sequence_length = 'd%0d. first_port_id = 'd%0d. second_port_id = 'd%0d. bypass_cache_initialisation = 'b%0b", 
      sequence_length, first_port_id, second_port_id, bypass_cache_initialisation));
    if (!is_supported(cfg))
      return;
    // By default put ACE ports in initialisation ports.
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(first_port_id);
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(second_port_id);

    // If the first_port_id (on which store accesses are sent) is ACE-Lite, then no need to initialize for CLEANUNIQUE
    // If both ports are ACE-Lite, no need for cache initialisation because ACE-Lite does not send CLEANUNIQUE
    if (
         (first_port_cleanunique_wt == 0) ||
         (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) || 
         (
           (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) && 
           (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) 
         ) 
       ) begin
      bypass_cleanunique_cache_initialisation = 1;
      `svt_xvm_debug("body",$sformatf("Bypassing cache initialisation for CLEANUNIQUE as it is not required. first_port_cleanunique_wt = 'd%0d. first_port_id = 'd%0d. second_port_id = 'd%0d",
      first_port_cleanunique_wt,first_port_id,second_port_id));
    end
    // If second port is ACE_LITE and there are no other ACE ports in the domain of these two ports,
    // then initialisation for cleanunique need not be done because cacheline will not be in shared state.
    else if (
         (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
         ((other_innershareable_ace_port == -1) && (other_outershareable_ace_port == -1))
       ) begin
      bypass_cleanunique_cache_initialisation = 1;
      `svt_xvm_debug("body",$sformatf("Bypassing cache initialisation for CLEANUNIQUE as it is not required. first_port_id = 'd%0d. second_port_id = 'd%0d. other_innershareable_ace_port = 'd%0d. other_outershareable_ace_port = 'd%0d",
      first_port_id,second_port_id,other_innershareable_ace_port,other_outershareable_ace_port));
    end
    if ((bypass_cleanunique_cache_initialisation != 1) &&
        (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) && 
        (first_port_cleanunique_wt != 0)) begin
      initialisation_length = sequence_length * first_port_cleanunique_wt/(first_port_makeunique_wt + first_port_cleanunique_wt + first_port_readunique_wt + first_port_writeunique_wt + first_port_writelineunique_wt);
      // Since the peer port is sending load transactions, all the lines to be invalidated.
      if (cfg.master_cfg[second_port_id].speculative_read_enable == 0)
        peer_port_invalidation_length = initialisation_length; 
      else
        peer_port_invalidation_length = 0; 
      disable_cleanunique_store_access = 0;
    end
    // Generate only one transaction so that we get a reference to the starting address
    // which in turn can be used for initialisation.
    `svt_xvm_create_on(init_xact_seq, p_sequencer.master_sequencer[first_port_id]) 
    init_xact_seq.makeunique_wt = first_port_makeunique_wt;
    init_xact_seq.readunique_wt = first_port_readunique_wt;
    init_xact_seq.cleanunique_wt = first_port_cleanunique_wt;
    init_xact_seq.writeunique_wt = first_port_writeunique_wt;
    init_xact_seq.writelineunique_wt = first_port_writelineunique_wt;
    send_dummy_sequence_for_xact_template(init_xact_seq,first_port_id,supports_both_domains,_domain_type,_master_xact);
    // Send some transactions to initialize memory with valid data
    `svt_xvm_debug("body",$sformatf("first_port_id='d%0d.second_port_id='d%0d.sequence_length='d%0d.initialisation_length='d%0d.peer_port_invalidation_length='d%0d.disable_cleanunique_store_access='b%0b.bypass_cache_initialisation='b%0b.bypass_cleanunique_cache_initialisation='b%0b.start_addr='h%0x",
    first_port_id,second_port_id,sequence_length,initialisation_length,peer_port_invalidation_length,disable_cleanunique_store_access,bypass_cache_initialisation,bypass_cleanunique_cache_initialisation,_master_xact.cacheline_addr()));
    if (!bypass_cache_initialisation) begin
      execute_cache_initialization_for_sequential_load_access(_master_xact.cacheline_addr(), sequence_length, second_port_id);
      if(cfg.master_cfg[first_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE && 
         cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE && (first_port_writeunique_wt == 1  &&  first_port_writelineunique_wt == 1))
        execute_cache_initialization_for_generic_sequential_access(_master_xact.cacheline_addr(),sequence_length,sequence_length,ace_domain_ports[0],ace_domain_ports[1],1);
    end

    if (!bypass_cache_initialisation && !bypass_cleanunique_cache_initialisation && !disable_cleanunique_store_access && (initialisation_length != 0) ) begin 
      string _ace_ports_str;
      if (ace_domain_ports.size() == 1)
        set_initialisation_ports(_master_xact,other_innershareable_ace_port,other_outershareable_ace_port,peer_port_invalidation_length,ace_domain_ports);

      foreach (ace_domain_ports[i]) begin
        _ace_ports_str = $sformatf("'d%0d ", ace_domain_ports[i]);
      end
      `svt_xvm_debug("body", $sformatf("ace_domain_ports: %s", _ace_ports_str));

      if (ace_domain_ports.size() != 2)
        bypass_cache_initialisation = 1;
      else
        execute_cache_initialization_for_generic_sequential_access(_master_xact.cacheline_addr(),initialisation_length,peer_port_invalidation_length,ace_domain_ports[0],ace_domain_ports[1],1);
    end

    // CLEANUNIQUE can be sent only if cache is initialised to some shared
    // state or svt_axi_port_configuration::speculative_read_enable is set.
    fork
    begin
      if (
           !disable_cleanunique_store_access && (initialisation_length != 0) &&
           (!bypass_cache_initialisation ||
            (cfg.master_cfg[first_port_id].speculative_read_enable && cfg.master_cfg[second_port_id].speculative_read_enable)
           )
      )  begin
        store_port_cleanunique_length = initialisation_length;
        `svt_xvm_create_on(first_port_cleanunique_store_seq, p_sequencer.master_sequencer[first_port_id]) 
        start_sequential_cleanunique_access(first_port_cleanunique_store_seq,init_xact_seq.start_addr,first_port_id,store_port_cleanunique_length,!supports_both_domains,init_xact_seq.directed_domain_type);
      end
      else 
        store_port_cleanunique_length = 0;
      `svt_xvm_create_on(first_port_non_cleanunique_store_seq, p_sequencer.master_sequencer[first_port_id]) 
      first_port_non_cleanunique_store_seq.makeunique_wt = first_port_makeunique_wt;
      first_port_non_cleanunique_store_seq.readunique_wt = first_port_readunique_wt;
      first_port_non_cleanunique_store_seq.writeunique_wt = first_port_writeunique_wt;
      first_port_non_cleanunique_store_seq.writelineunique_wt = first_port_writelineunique_wt;
      start_generic_sequential_access(first_port_non_cleanunique_store_seq,(init_xact_seq.start_addr+store_port_cleanunique_length*cfg.master_cfg[first_port_id].cache_line_size),
                                      first_port_id, (sequence_length-store_port_cleanunique_length),
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    begin
      `svt_xvm_create_on(second_port_load_seq, p_sequencer.master_sequencer[second_port_id]) 
      second_port_load_seq.readshared_wt = second_port_readshared_wt; 
      second_port_load_seq.readnotshareddirty_wt = second_port_readnotshareddirty_wt; 
      second_port_load_seq.readclean_wt = second_port_readclean_wt; 
      second_port_load_seq.readonce_wt = second_port_readonce_wt; 
      start_generic_sequential_access(second_port_load_seq,init_xact_seq.start_addr,
                                      second_port_id, sequence_length,
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
    end
    join

    if (first_port_cleanunique_store_seq != null)
      first_port_cleanunique_store_seq.wait_for_active_xacts_to_end();

    if (first_port_non_cleanunique_store_seq != null)
      first_port_non_cleanunique_store_seq.wait_for_active_xacts_to_end();

    if (second_port_load_seq != null)
      second_port_load_seq.wait_for_active_xacts_to_end();

  endtask

  virtual function bit normalize_weights_based_on_interface_type();
    normalize_weights_based_on_interface_type = 1;
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      first_port_makeunique_wt = 0; 
      first_port_readunique_wt = 0;
      first_port_cleanunique_wt = 0;
    end
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      second_port_readshared_wt = 0;
      second_port_readnotshareddirty_wt = 0;
      second_port_readclean_wt = 0;
    end
    if ((first_port_makeunique_wt + first_port_readunique_wt + first_port_cleanunique_wt + first_port_writeunique_wt + first_port_writelineunique_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for store transactions in first_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", first_port_id));
    end
    if ((second_port_readshared_wt + second_port_readnotshareddirty_wt + second_port_readclean_wt + second_port_readonce_wt) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for load transactions in second_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", second_port_id));
    end
    if (bypass_cache_initialisation) begin
      first_port_cleanunique_wt = 0;
    end
  endfunction

endclass

/**
  * Sends a set of concurrent, sequential cmo accesses from first_port_id and store
  * accesses from second_port_id to the same set of overlapping addresses. 
  * CMO type transactions can be MAKEINVALID, CLEANINVALID
  * or CLEANSHARED.The store type transactions can be MAKEUNIQUE, READUNIQUE, CLEANUNIQUE,
  * WRITEUNIQUE or WRITELINEUNIQUE  based on the interface types of the ports and the weights.
  * an initialisation procedure is invoked based on the following sequence, unless
  * Prior to sending the cmo and store transaction bypass_cache_initialisation is set:
  * - In order that the store transactions can be fired from various initial states.  
  * .
  * - If second_port_cleanunique_wt is not zero, cachelines are
  * initialised, since CLEANUNIQUE can be sent only from a cacheline in shared
  * state. Only cachelines from which CLEANUNIQUE needs to be sent are
  * initialized. The number of CLEANUNIQUE transactions sent are determined by
  * the formula sequence_length*first_port_cleanunique_wt/(sum of weights of
  * all xact types in second port).  Initialisation is done by sending
  * MAKEUNIQUE transactions from one ACE port and READSHARED transactions from
  * another ACE port to the same set of addresses. Snoop transactions for
  * READSHARED type snoop are programmed (in the corresponding tests) to always
  * assert svt_axi_snoop_transaction::snoop_resp_datatransfer and
  * svt_axi_snoop_transaction::snoop_resp_isshared so that a shared state of
  * the cacheline can be acheived in both masters.  All shared cachelines in
  * first_port_id are invalidated so that the cmo transactions can be sent on
  * the interface.  
  * .
  * After this initialisation, sequential cmo access from first_port_id and
  * sequential store from second_port_id are sent.
  * .
  * Sometimes if the cmo transactions snoops the second_port firstly and
  * second port transaction is CLEANUNIQUE transaction means, there is a chance of
  * invalidation of the cache line of second_port. By the result of this scenario
  * the second_port may drop the CLEANUNIQUE transactions, Because CLEANUNIQUE
  * cant be sent from INVALID state.
  */
class svt_axi_ace_master_two_port_overlapping_addr_cmo_and_store_sequential_sequence extends svt_axi_ace_master_two_port_base_sequential_virtual_sequence;
  
  /** 
    * Bypass cache initialisation. CLEANUNIQUE transactions cannot be sent if
    * cache initialisation is bypassed since CLEANUNIQUE transactions require
    * cache to be in shared state
    */
  bit bypass_cache_initialisation = 0;

  /** Weightage for MAKEINVALID cmo transactions for first_port_id */
  int first_port_makeinvalid_wt = 1;

  /** Weightage for CLEANINVALID cmo transactions for first_port_id */
  int first_port_cleaninvalid_wt = 1;

  /** Weightage for CLEANSHARED cmo transactions for first_port_id */
  int first_port_cleanshared_wt = 1;
  
  /** Weightage for CLEANSHAREDPERSIST cmo transactions for first_port_id */
  int first_port_cleansharedpersist_wt = 1;

  /** Weightage for MAKEUNIQUE store transactions for second_port_id */
  int second_port_makeunique_wt = 1;

  /** Weightage for READUNIQUE store transactions for second_port_id */
  int second_port_readunique_wt = 1;

  /** Weightage for CLEANUNIQUE store transactions for second_port_id */
  int second_port_cleanunique_wt = 1;

  /** Weightage for WRITEUNIQUE store transactions for second_port_id */
  int second_port_writeunique_wt = 0;

  /** Weightage for WRITELINEUNIQUE store transactions for second_port_id */
  int second_port_writelineunique_wt = 0;

  constraint reasonable_supported_xact_category {
    first_port_xact_category == CMO;
    second_port_xact_category == STORE_OPERATION;
  } 

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_two_port_overlapping_addr_cmo_and_store_sequential_sequence)
    
  function new(string name = "svt_axi_ace_master_two_port_overlapping_addr_cmo_and_store_sequential_sequence");
    super.new(name);
  endfunction

  virtual task body();
    svt_axi_master_transaction _master_xact;
    svt_axi_ace_master_generic_sequence init_xact_seq, first_port_cmo_seq;
    svt_axi_ace_master_generic_sequence second_port_cleanunique_store_seq, second_port_non_cleanunique_store_seq;
    svt_axi_ace_master_generic_sequence second_port_readunique_store_seq;
    svt_axi_transaction::xact_shareability_domain_enum _domain_type;
    bit supports_both_domains = 0;
    int initialisation_length, peer_port_invalidation_length, ace_domain_ports[$];
    bit disable_cleanunique_store_access = 0;
    int other_innershareable_ace_port, other_outershareable_ace_port;
    int store_port_cleanunique_length;
    int store_port_readunique_length;
    bit bypass_cleanunique_cache_initialisation = 0;
    bit bypass_store_initialisation = 0;
    bit store_initialization_select = 0;
    bit status;
    
    super.body();

  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_makeinvalid_wt",first_port_makeinvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleaninvalid_wt",first_port_cleaninvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleanshared_wt",first_port_cleanshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_cleansharedpersist_wt",first_port_cleansharedpersist_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_makeunique_wt",second_port_makeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_readunique_wt",second_port_readunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_cleanunique_wt",second_port_cleanunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_writeunique_wt",second_port_writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_port_writelineunique_wt",second_port_writelineunique_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "bypass_cache_initialisation",bypass_cache_initialisation);

  `elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_makeinvalid_wt"}, first_port_makeinvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleaninvalid_wt"}, first_port_cleaninvalid_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleanshared_wt"}, first_port_cleanshared_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_cleansharedpersist_wt"}, first_port_cleansharedpersist_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_makeunique_wt"}, second_port_makeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_readunique_wt"}, second_port_readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_cleanunique_wt"}, second_port_cleanunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_writeunique_wt"}, second_port_writeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".second_port_writelineunique_wt"}, second_port_writelineunique_wt); 
    status = m_sequencer.get_config_int({get_type_name(), ".bypass_cache_initialisation"}, bypass_cache_initialisation);
  `endif
    disable_cleanunique_store_access = 1;
    is_supported_weights = normalize_weights_based_on_interface_type();
    is_supported_domains = get_domain_type_for_two_port_sequence(first_port_id,second_port_id,supports_both_domains,_domain_type,other_innershareable_ace_port,other_outershareable_ace_port);
    if (!is_supported(cfg))
      return;
    // By default put ACE ports in initialisation ports.
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(first_port_id);
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
      ace_domain_ports.push_back(second_port_id);

    // If the second_port_id (on which store accesses are sent) is ACE-Lite, then no need to initialize for CLEANUNIQUE
    // If both ports are ACE-Lite, no need for cache initialisation because ACE-Lite does not send CLEANUNIQUE
    if (
         (second_port_cleanunique_wt == 0) ||
         (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) || 
         (
           (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) && 
           (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) 
         ) 
       ) begin
      bypass_cleanunique_cache_initialisation = 1;
      `svt_xvm_debug("body",$sformatf("Bypassing cache initialisation for CLEANUNIQUE as it is not required. second_port_cleanunique_wt = 'd%0d. second_port_id = 'd%0d. second_port_id = 'd%0d",  second_port_cleanunique_wt,second_port_id,second_port_id));
    end
    // If second port is ACE_LITE and there are no other ACE ports in the domain of these two ports,
    // then initialisation for cleanunique need not be done because cacheline will not be in shared state.
    else if (
         ((cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
         ((other_innershareable_ace_port == -1) && (other_outershareable_ace_port == -1)))
       ) begin
      bypass_cleanunique_cache_initialisation = 1;
      `svt_xvm_debug("body",$sformatf("Bypassing cache initialisation for CLEANUNIQUE as it is not required. first_port_id = 'd%0d. second_port_id = 'd%0d. other_innershareable_ace_port = 'd%0d. other_outershareable_ace_port = 'd%0d",first_port_id,second_port_id,other_innershareable_ace_port,other_outershareable_ace_port));
    end
    
    //The for initialization of store, MAKEUNIQUE will be sent from first_port_id, If first_port_id is ACE_LITE 
    //then it cant fire MAKEUNIQUE, So the another ACE port selected through the set_initialisation_ports must fire MAKEUNIQUE.
    //If the first_port_id is ACE-Lite and second_port_id is AXI_ACE, then the store_initialization_select must be set to one
    //If both first_port_id and second_port_id are AXI_ACE, then the store_initialization_select must be set to zero
    if (
         (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) && 
         (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) 
      )  begin
      store_initialization_select = 1;
    end
    else if (
         (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) && 
         (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) 
       ) begin
      store_initialization_select = 0;
    end
    // If the second_port_id is ACE-Lite(on which store accesses are sent), then no need to initialize the cache lines  
    else if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE)
      bypass_store_initialisation = 1;
  
    if (
         (bypass_cleanunique_cache_initialisation != 1) &&
         (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) && (second_port_cleanunique_wt != 0)
      ) begin
      initialisation_length = sequence_length * second_port_cleanunique_wt/(second_port_makeunique_wt + second_port_cleanunique_wt + second_port_readunique_wt + second_port_writeunique_wt + second_port_writelineunique_wt);
      peer_port_invalidation_length = 0; 
      disable_cleanunique_store_access = 0;
    end

    // Generate only one transaction so that we get a reference to the starting address
    // which in turn can be used for initialisation.
    `svt_xvm_create_on(init_xact_seq, p_sequencer.master_sequencer[first_port_id]) 
    init_xact_seq.makeinvalid_wt = first_port_makeinvalid_wt;
    init_xact_seq.cleaninvalid_wt = first_port_cleaninvalid_wt;
    init_xact_seq.cleanshared_wt = first_port_cleanshared_wt;
    init_xact_seq.cleansharedpersist_wt = first_port_cleansharedpersist_wt;
    init_xact_seq.generate_only_shareable_domain = 1;
    
    send_dummy_sequence_for_xact_template(init_xact_seq,first_port_id,supports_both_domains,_domain_type,_master_xact);
    // Send some transactions to initialize memory with valid data
    `svt_xvm_debug("body",$sformatf("first_port_id='d%0d.second_port_id='d%0d.sequence_length='d%0d.initialisation_length='d%0d.peer_port_invalidation_length='d%0d.disable_cleanunique_store_access='b%0b.bypass_cache_initialisation='b%0b.bypass_cleanunique_cache_initialisation='b%0b.start_addr='h%0x, supports_both_domains ='d%0d",first_port_id,second_port_id,sequence_length,initialisation_length,peer_port_invalidation_length,disable_cleanunique_store_access,bypass_cache_initialisation,bypass_cleanunique_cache_initialisation,_master_xact.cacheline_addr(),supports_both_domains));
    
    // Initializing the store port cachelines
    if (!bypass_cache_initialisation && !bypass_store_initialisation) begin
      string _ace_ports_str = "";
      
      //selecting one another ace port in the sharable domain, for performing initialization
      if (ace_domain_ports.size() == 1)
        begin
        set_initialisation_ports(_master_xact,other_innershareable_ace_port,other_outershareable_ace_port,peer_port_invalidation_length,ace_domain_ports);
        end

      foreach (ace_domain_ports[i]) begin
        _ace_ports_str = $sformatf("'d%0d ", ace_domain_ports[i]);
      end
      `svt_xvm_debug("body", $sformatf("ace_domain_ports: %s", _ace_ports_str));

      if (ace_domain_ports.size() != 2)
        bypass_cache_initialisation = 1;
      else begin
        //If store_initialization_select is high, then the ace_domain_ports[1] will be sent as the first_port_id and 
        //ace_domain_ports[0] as the peer_port_id, for the inputs of the task execute_cache_initialization_for_cmo_store (Which is going to perform initialization)
        if (store_initialization_select) begin
          //For cached store, the input store_select of the task will be passed as 1 
          if (
               ((second_port_makeunique_wt + second_port_cleanunique_wt + second_port_readunique_wt) != 0) &&
               !bypass_cleanunique_cache_initialisation && !disable_cleanunique_store_access &&
               (initialisation_length != 0) 
            )
          execute_cache_initialization_for_cmo_store(_master_xact.cacheline_addr(), sequence_length, ace_domain_ports[1],ace_domain_ports[0],initialisation_length, 1, 0);
          //For non_cached store, the input store_select of the task will be passed as 0
          else 
          execute_cache_initialization_for_cmo_store(_master_xact.cacheline_addr(), sequence_length, ace_domain_ports[1],ace_domain_ports[0],0,0,0);
        end
        //If store_initialization_select is low, then the ace_domain_ports[0] will be sent as the first_port_id and 
        //ace_domain_ports[1] as the peer_port_id, for the inputs of the task execute_cache_initialization_for_cmo_store
        else begin
          if (
               ((second_port_makeunique_wt + second_port_cleanunique_wt + second_port_readunique_wt) != 0) &&
               !bypass_cleanunique_cache_initialisation && !disable_cleanunique_store_access &&
               (initialisation_length != 0) 
            )
          execute_cache_initialization_for_cmo_store(_master_xact.cacheline_addr(), sequence_length, ace_domain_ports[0],ace_domain_ports[1],initialisation_length, 1, 1);
          else 
          execute_cache_initialization_for_cmo_store(_master_xact.cacheline_addr(), sequence_length, ace_domain_ports[0],ace_domain_ports[1],0,0,1);
        end
      end 
    end

    // CLEANUNIQUE can be sent only if cache is initialised to some shared
    // state or svt_axi_port_configuration::speculative_read_enable is set.
    // CLEANUNIQUE sequence_length, start_addr will be fixed based on the start_addr and initialisation_length of the READUNIQUE access.
    fork
      begin
      `svt_xvm_create_on(first_port_cmo_seq, p_sequencer.master_sequencer[first_port_id]) 
      first_port_cmo_seq.makeinvalid_wt = first_port_makeinvalid_wt; 
      first_port_cmo_seq.cleaninvalid_wt = first_port_cleaninvalid_wt; 
      first_port_cmo_seq.cleanshared_wt = first_port_cleanshared_wt;
      first_port_cmo_seq.cleansharedpersist_wt = first_port_cleansharedpersist_wt;
      start_generic_sequential_access(first_port_cmo_seq,init_xact_seq.start_addr,
                                      first_port_id, sequence_length,
                                      !supports_both_domains,init_xact_seq.directed_domain_type);
      end
      begin
      if (
           (initialisation_length != 0) &&
           (!bypass_cache_initialisation ||
            (cfg.master_cfg[first_port_id].speculative_read_enable && cfg.master_cfg[second_port_id].speculative_read_enable)
           )
      )  begin
         store_port_readunique_length  = initialisation_length;
         `svt_xvm_create_on(second_port_readunique_store_seq, p_sequencer.master_sequencer[second_port_id]) 
         second_port_readunique_store_seq.readunique_wt = second_port_readunique_wt;
         start_generic_sequential_access(second_port_readunique_store_seq, init_xact_seq.start_addr,second_port_id,store_port_readunique_length,!supports_both_domains,init_xact_seq.directed_domain_type);
         if (!disable_cleanunique_store_access)
           begin
           store_port_cleanunique_length = initialisation_length;
           `svt_xvm_create_on(second_port_cleanunique_store_seq, p_sequencer.master_sequencer[second_port_id]) 
           start_sequential_cleanunique_access(second_port_cleanunique_store_seq,(init_xact_seq.start_addr + (store_port_cleanunique_length * cfg.master_cfg[second_port_id].cache_line_size)),second_port_id,store_port_cleanunique_length,!supports_both_domains,init_xact_seq.directed_domain_type);
           end
      end
      else begin
        store_port_cleanunique_length = 0;
        store_port_readunique_length  = 0;
      end

      `svt_xvm_create_on(second_port_non_cleanunique_store_seq, p_sequencer.master_sequencer[second_port_id]) 
      second_port_non_cleanunique_store_seq.makeunique_wt = second_port_makeunique_wt;
      second_port_non_cleanunique_store_seq.writeunique_wt = second_port_writeunique_wt;
      second_port_non_cleanunique_store_seq.writelineunique_wt = second_port_writelineunique_wt;
      start_generic_sequential_access(second_port_non_cleanunique_store_seq,(init_xact_seq.start_addr+((store_port_cleanunique_length + store_port_readunique_length) *cfg.master_cfg[second_port_id].cache_line_size)),second_port_id, (sequence_length-(store_port_cleanunique_length + store_port_readunique_length)),!supports_both_domains,init_xact_seq.directed_domain_type);   
    end 
    join

    if (second_port_cleanunique_store_seq != null)
      second_port_cleanunique_store_seq.wait_for_active_xacts_to_end();

    if (second_port_non_cleanunique_store_seq != null)
      second_port_non_cleanunique_store_seq.wait_for_active_xacts_to_end();

    if (second_port_readunique_store_seq != null)
      second_port_readunique_store_seq.wait_for_active_xacts_to_end();

    if (first_port_cmo_seq != null)
      first_port_cmo_seq.wait_for_active_xacts_to_end();

  endtask

  virtual function bit normalize_weights_based_on_interface_type();
    normalize_weights_based_on_interface_type = 1;
    if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      second_port_makeunique_wt = 0; 
      second_port_readunique_wt = 0;
      second_port_cleanunique_wt = 0; 
    end
    if ((first_port_makeinvalid_wt + first_port_cleaninvalid_wt + first_port_cleanshared_wt + first_port_cleansharedpersist_wt ) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for cmo transactions in first_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", first_port_id));
    end
    if ((second_port_makeunique_wt + second_port_readunique_wt + second_port_cleanunique_wt + second_port_writeunique_wt + second_port_writelineunique_wt ) == 0) begin
      normalize_weights_based_on_interface_type = 0;
      `svt_xvm_error("normalize_weights_based_on_interface_type", $sformatf("The sum of all the valid weights for store transactions in second_port_id('d%0d) after normalizing for interface type is 0. \
                     Please ensure that the weight of at least one transaction which is allowed to be sent on this interface is non-zero", second_port_id));
    end
  endfunction
endclass

/**
  * This sequence is a base class for all barier based sequences. This sequence cannot be run
  * as such, but contains methods which are used by other barrier sequences
  *
  * NOTE: Continuous polling may need adding interval between two consecutive transactions. See
  *       poll_barrier_flag_and_check_post_barrier_contents task for details.
  */
class svt_axi_ace_master_barrier_base_virtual_sequence extends svt_axi_ace_master_base_virtual_sequence;
  
  int unsigned sequence_length = 10;

  rand svt_axi_transaction::xact_shareability_domain_enum domain_type;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_barrier_base_virtual_sequence)
  
  function new(string name = "svt_axi_ace_master_barrier_base_virtual_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    bit status;
    super.pre_body();
    raise_phase_objection();

`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
`endif
  endtask

 /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

  virtual task body();
    super.body();
  endtask: body

  /**
    * Creates a pre barrier sequence to store (write)
    * @param length The number of pre barrier transactions required
    * @param port_id The port_id on which these pre barrier transactions will be executed
    * @param makeunique_wt The weightage for a MAKEUNIQUE transaction
    * @param readunique_wt The weightage for a READUNIQUE transaction
    * @param writelineunique_wt The weightage for a WRITELINEUNIQUE_wt transaction
    * @param writeunique_wt The weightage for a WRITEUNIQUE_wt transaction
    */
  function svt_axi_ace_master_base_sequence create_pre_barrier_store_seq(
                int length,int port_id,
                int makeunique_wt, int readunique_wt, int writelineunique_wt, int writeunique_wt
                );
    svt_axi_ace_master_base_sequence pre_barrier_coherent_seq;
    `svt_xvm_create_on(pre_barrier_coherent_seq, p_sequencer.master_sequencer[port_id])
    pre_barrier_coherent_seq.disable_all_weights();
    pre_barrier_coherent_seq.force_to_cache_line_size = 1;
    pre_barrier_coherent_seq.use_directed_domain_type = 1;
    pre_barrier_coherent_seq.directed_domain_type = domain_type;
    if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
      pre_barrier_coherent_seq.makeunique_wt = 1;
      pre_barrier_coherent_seq.readunique_wt = 1;
      pre_barrier_coherent_seq.writelineunique_wt = 1;
    end
    else if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      pre_barrier_coherent_seq.writelineunique_wt = 1;
      pre_barrier_coherent_seq.writeunique_wt = 1;
    end
    else begin
      // Error
      return (null);
    end
    // Send pre-barrier transactions
    void'(pre_barrier_coherent_seq.randomize with {use_directed_addr == 0;sequence_length==length;});
    create_pre_barrier_store_seq = pre_barrier_coherent_seq;
  endfunction

  /**
    * Creates a post barrier sequence to load (read)
    * @param length The number of pre barrier transactions required
    * @param port_id The port_id on which these pre barrier transactions will be executed
    * @param readonce_wt The weightage for a READONCE transaction
    * @param readshared_wt The weightage for a READSHARED transaction
    * @param readnotshareddirty_wt The weightage for a READNOTSHAREDDIRTY transaction
    * @param readclean_wt The weightage for a READCLEAN transaction
    */
  function svt_axi_ace_master_base_sequence create_pre_barrier_load_seq(
          int length, int port_id, int readonce_wt, int readshared_wt, int readnotshareddirty_wt, int readclean_wt, bit is_directed_addr = 0
                );
    svt_axi_ace_master_base_sequence pre_barrier_load_seq;
    `svt_xvm_create_on(pre_barrier_load_seq, p_sequencer.master_sequencer[port_id])
    pre_barrier_load_seq.disable_all_weights();
    if ((domain_type == svt_axi_transaction::INNERSHAREABLE) ||
        (domain_type == svt_axi_transaction::OUTERSHAREABLE))
      pre_barrier_load_seq.initialize_cachelines = 1;
    pre_barrier_load_seq.use_directed_domain_type = 1;
    pre_barrier_load_seq.directed_domain_type = domain_type;
    if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
      pre_barrier_load_seq.readonce_wt = 1;
      pre_barrier_load_seq.readshared_wt = 1;
      pre_barrier_load_seq.readnotshareddirty_wt = 1;
      pre_barrier_load_seq.readclean_wt = 1;
      pre_barrier_load_seq.readnosnoop_wt = 1;
    end
    else if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      pre_barrier_load_seq.readonce_wt = 1;
      pre_barrier_load_seq.readnosnoop_wt = 1;
    end
    else begin
      // Error
    end
    void'(pre_barrier_load_seq.randomize with {use_directed_addr == is_directed_addr;sequence_length == length;});
    // We want entire cacheline size to be read for all transactions
    pre_barrier_load_seq.force_to_cache_line_size = 1;
    create_pre_barrier_load_seq = pre_barrier_load_seq;
  endfunction

  /**
    * Creates a poast barrier sequence to load (read)
    * @param length The number of pre barrier transactions required
    * @param port_id The port_id on which these pre barrier transactions will be executed
    * @param readonce_wt The weightage for a READONCE transaction
    * @param readshared_wt The weightage for a READSHARED transaction
    * @param readnotshareddirty_wt The weightage for a READNOTSHAREDDIRTY transaction
    * @param readclean_wt The weightage for a READCLEAN transaction
    */
  function svt_axi_ace_master_base_sequence create_post_barrier_load_seq(
          int length, int port_id, int readonce_wt, int readshared_wt, int readnotshareddirty_wt, int readclean_wt
                );
    svt_axi_ace_master_base_sequence post_barrier_read_seq;
    // Read back from memory locations written through pre_barrier_xacts and check results
    `svt_xvm_create_on(post_barrier_read_seq, p_sequencer.master_sequencer[port_id])
    post_barrier_read_seq.disable_all_weights();
    post_barrier_read_seq.initialize_cachelines = 0;
    post_barrier_read_seq.direct_addr_timeout = 1000000;
    post_barrier_read_seq.use_directed_domain_type = 1;
    post_barrier_read_seq.directed_domain_type = domain_type;
    if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
      post_barrier_read_seq.readonce_wt = 1;
      post_barrier_read_seq.readshared_wt = 1;
      post_barrier_read_seq.readnotshareddirty_wt = 1;
      post_barrier_read_seq.readclean_wt = 1;
      post_barrier_read_seq.readnosnoop_wt = 1;
    end
    else if (cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      post_barrier_read_seq.readonce_wt = 1;
      post_barrier_read_seq.readnosnoop_wt = 1;
    end
    else begin
      // Error
    end
    void'(post_barrier_read_seq.randomize with {use_directed_addr == 1;sequence_length == length;});
    // We want entire cacheline size to be read for all transactions
    post_barrier_read_seq.force_to_cache_line_size = 1;
    create_post_barrier_load_seq = post_barrier_read_seq;
  endfunction

  /**
    * Creates a post barrier transaction by associating it with the given
    * write and read barriers. The post barrier transaction is a WRITEUNIQUE
    * transaction that addresses a single byte. 
    * @param port_id The port on which the post barrier must be sent
    * @param write_barrier_xact The WRITE barrier transaction to which to associate
    *        the post barrier
    * @param read_barrier_xact The READ barrier transaction to which to associate
    *        the post barrier
    * @param is_single_byte_flag_xact Indicates if the post barrier should be a transaction
    *        that addresses a single byte. This is currently always single byte irrespective
    *        of what is passed here
    * @param post_barrier_xact The output post_barrier transaction
    */
  task send_post_barrier_xact (int port_id,
                               svt_axi_master_transaction write_barrier_xact,
                               svt_axi_master_transaction read_barrier_xact,
                               bit is_single_byte_flag_xact,
                               output svt_axi_master_transaction post_barrier_xact 
                              );
    svt_axi_ace_barrier_flag_write_xact_sequence post_barrier_seq;
    // Send post barrier transaction
    `svt_xvm_debug("send_post_barrier_xact",$sformatf("Sending post barrier xact on port 'd%0d.",port_id));
    `svt_xvm_create_on(post_barrier_seq, p_sequencer.master_sequencer[port_id])
    void'(post_barrier_seq.randomize() with {flag_domain_type == local::domain_type;});
    post_barrier_seq.assoc_write_barrier_xact = write_barrier_xact;
    post_barrier_seq.assoc_read_barrier_xact = read_barrier_xact;
    post_barrier_seq.is_single_byte_flag_xact = is_single_byte_flag_xact;
    post_barrier_seq.start(p_sequencer.master_sequencer[port_id]);
    post_barrier_xact = post_barrier_seq.output_xact;
  endtask

  /**
    * Sends a barrier sequences that consists of
    * Pre barrier transactions as given in pre_barrier_seq
    * A barrier pair (WRITEBARRIER and READBARRIER)
    * @param pre_barrier_seq Handle to pre barrier sequence
    */
  task send_barrier_sequence(int port_id, 
                             svt_axi_ace_master_base_sequence pre_barrier_seq, 
                             output svt_axi_master_transaction pre_barrier_xacts[$],
                             output svt_axi_ace_barrier_pair_sequence barrier_pair_seq
                             );
    svt_axi_ace_barrier_pair_sequence _barrier_pair_seq;
    `svt_xvm_debug("send_barrier_sequence",$sformatf("Sending barrier sequence on port 'd%0d. num_pre_barrier_xacts = 'd%d",port_id,pre_barrier_seq.sequence_length));
    pre_barrier_seq.start(p_sequencer.master_sequencer[port_id]);
    // Send the barrier pair
    `svt_xvm_create_on(_barrier_pair_seq, p_sequencer.master_sequencer[port_id])
    _barrier_pair_seq.myDomain = this.domain_type;
    _barrier_pair_seq.start(p_sequencer.master_sequencer[port_id]);
    while (pre_barrier_seq.output_xact_mailbox.num()) begin
      svt_axi_master_transaction _master_xact;
      pre_barrier_seq.output_xact_mailbox.get(_master_xact);
      pre_barrier_xacts.push_back(_master_xact);
    end
    barrier_pair_seq = _barrier_pair_seq;
    //wait (`SVT_AXI_XACT_STATUS_ENDED(barrier_flag_write_seq.output_write_xact));
  endtask

  /**
    * This task continuosly reads from port_id, the location written through barrier_flag_xact 
    * When the value returned is equal to the post barrier flag xact, the loop terminates
    * and all locations written through the pre barrier transactions (given in pre_barrier_xacts)
    * are read back using post_barrier_read_seq. The locations read back are checked for data
    * consistency to ensure that all the pre barrier barrier transactions are observed correctly.
    * @param port_id The port from which the flag set through barrier_flag_xact is to be read
    *                The same port_id is used to send post_barrier_read_seq
    * @param post_barrier_read_seq The sequence to be used to read all the location written
    *                through pre_barrier_xacts
    * @param pre_barrier_xacts The pre barrier store transactions that need to be read back 
    * @param barrier_flag_xact The transaction used as a flag to indicate that all the pre-barrier
    *                transactions are observable to any transaction that can observe the flag
    *
    * NOTE: Continuous polling may need adding interval between two consecutive transactions
    *      Interconnect can enter into deadlock condition if master sends continuous transactions
    *      without any gap in between two consecutive transactions targeted to a particular address.
    *      CCI400 has this restriction where if a hazarded address is polled continuously then other
    *      pending transaction issued by other master sent to the same address never gets selected
    *      to proceed further and remains in hang state.
    *      System Configuration parameter ic_num_cycles_interval_for_polling_hazarded_address can be
    *      used to introduce interval in polling in terms of number of cycles.
    */
  task poll_barrier_flag_and_check_post_barrier_contents(int port_id,
                                           svt_axi_ace_master_base_sequence post_barrier_read_seq,
                                           svt_axi_master_transaction pre_barrier_xacts[$],
                                           svt_axi_master_transaction barrier_flag_xact);
    virtual svt_axi_master_if axi_master_if;
    svt_axi_ace_master_base_sequence mem_read_seq;
    svt_axi_master_transaction first_port_master_xact;
    svt_axi_master_transaction post_barrier_read_xacts[$];

    axi_master_if = cfg.axi_if.get_master_if(port_id);

    while (1) begin
      svt_axi_ace_barrier_flag_read_xact_sequence barrier_flag_read_seq;
      bit[7:0] byte_flag_data,observed_byte_flag_data;
      bit[`SVT_AXI_MAX_DATA_WIDTH-1:0] full_flag_data,observed_full_flag_data;
      `svt_xvm_create_on(barrier_flag_read_seq, p_sequencer.master_sequencer[port_id])
      void'(barrier_flag_read_seq.randomize() with {
        flag_addr == barrier_flag_xact.addr;
        flag_domain_type == barrier_flag_xact.domain_type;
      });
      barrier_flag_read_seq.start(p_sequencer.master_sequencer[port_id]);
      `svt_xvm_debug("body", {"Flag transaction",`SVT_AXI_PRINT_PREFIX1(barrier_flag_read_seq.output_read_xact), "sent."})
      wait (`SVT_AXI_XACT_STATUS_ENDED(barrier_flag_read_seq.output_read_xact));
      full_flag_data = barrier_flag_xact.data[0];
      byte_flag_data = full_flag_data[7:0];
      observed_full_flag_data = barrier_flag_read_seq.output_read_xact.data[0];
      observed_byte_flag_data = observed_full_flag_data[7:0];
      if (observed_byte_flag_data == byte_flag_data) begin
        `svt_xvm_debug("body", {"Flag transaction",`SVT_AXI_PRINT_PREFIX1(barrier_flag_read_seq.output_read_xact), "ended, Flag location is successfully read back.",$sformatf("data = 'h%0x",barrier_flag_read_seq.output_read_xact.data[0])})
        break;
      end
      else 
        `svt_xvm_debug("body", {"Flag transaction",`SVT_AXI_PRINT_PREFIX1(barrier_flag_read_seq.output_read_xact), "ended, but flag is not yet set.",$sformatf("flag data = 'h%0x. observed data = 'h%0x",byte_flag_data,observed_byte_flag_data)})

        // Interconnect can enter into deadlock condition if master sends continuous transactions
        // without any gap in between two consecutive transactions targeted to a particular address.
        // CCI400 has this restriction where if a hazarded address is polled continuously then other
        // pending transaction issued by other master sent to the same address never gets selected
        // to proceed further and remains in hang state.
        //
        repeat(cfg.ic_num_cycles_interval_for_polling_hazarded_address) 
          @(axi_master_if.axi_monitor_cb);
          //@(posedge cfg.axi_if.common_aclk);
    end 
    foreach (pre_barrier_xacts[i])
      post_barrier_read_seq.directed_addr_mailbox.put(pre_barrier_xacts[i].addr);
    post_barrier_read_seq.start(p_sequencer.master_sequencer[port_id]);
    post_barrier_read_seq.wait_for_active_xacts_to_end();
    while (post_barrier_read_seq.output_xact_mailbox.num()) begin
      svt_axi_master_transaction _master_xact;
      post_barrier_read_seq.output_xact_mailbox.get(_master_xact);
      post_barrier_read_xacts.push_back(_master_xact);
    end
    check_pre_barrier_and_post_barrier_xact_contents(pre_barrier_xacts,post_barrier_read_xacts);
  endtask

  function void check_pre_barrier_and_post_barrier_xact_contents(svt_axi_master_transaction pre_barrier_xacts[$],
                                                                 svt_axi_master_transaction post_barrier_xacts[$]
                                                                );
    // Check contents of read transactions
    if (post_barrier_xacts.size() != pre_barrier_xacts.size()) begin
      `svt_xvm_error("check_pre_barrier_and_post_barrier_xact_contents",
      $sformatf("Number of memory reads('d%0d) and number of pre_barrier write tarnsactions('d%0d) must be same, but they are not",post_barrier_xacts.size(),pre_barrier_xacts.size()));
    end
    else begin
      foreach (pre_barrier_xacts[i]) begin
        bit[7:0] write_xact_data_stream[],read_xact_byte_stream[]; 
        bit write_xact_wstrb_stream[];
        if (pre_barrier_xacts[i].transmitted_channel == svt_axi_transaction::WRITE) begin
          pre_barrier_xacts[i].pack_data_to_byte_stream(pre_barrier_xacts[i].data,write_xact_data_stream);
          pre_barrier_xacts[i].pack_wstrb_to_byte_stream(pre_barrier_xacts[i].wstrb,write_xact_wstrb_stream);
          if (write_xact_data_stream.size() != write_xact_wstrb_stream.size()) begin
            `svt_error("check_pre_barrier_and_post_barrier_xact_contents",
            $psprintf("The sizes of data and wstrb after packing do not match for xact %0s. Exiting check. data.size() = 'd%0d. wstrb.size() = 'd%0d",
            `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),write_xact_data_stream.size(),write_xact_wstrb_stream.size()));
            break;
          end
        end
        else begin
          pre_barrier_xacts[i].pack_data_to_byte_stream(pre_barrier_xacts[i].cache_write_data,write_xact_data_stream);
        end

        `svt_xvm_debug("check_pre_barrier_and_post_barrier_xact_contents",
        $sformatf("Checking pre_barrier_xacts and corresponding memory reads contents. pre_barrier xact: %0s. mem_read xact: %0s",
        `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),`SVT_AXI_PRINT_PREFIX1(post_barrier_xacts[i])));
        if(((pre_barrier_xacts[i].burst_type  != svt_axi_transaction::WRAP && 
             post_barrier_xacts[i].burst_type != svt_axi_transaction::WRAP) && 
            pre_barrier_xacts[i].addr != post_barrier_xacts[i].addr) ||
           ((pre_barrier_xacts[i].burst_type  == svt_axi_transaction::WRAP ||
             post_barrier_xacts[i].burst_type == svt_axi_transaction::WRAP) &&
            pre_barrier_xacts[i].cacheline_addr() != post_barrier_xacts[i].cacheline_addr()) )begin
          // Error
          `svt_xvm_error("check_pre_barrier_and_post_barrier_xact_contents",
           $sformatf("Expected pre_barrier_xacts and corresponding memory reads to be in same order, but they are not. pre_barrier xact: %0s. mem_read xact: %0s",
           `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),`SVT_AXI_PRINT_PREFIX1(post_barrier_xacts[i])));
        end
        else begin
          post_barrier_xacts[i].pack_data_to_byte_stream(post_barrier_xacts[i].data,read_xact_byte_stream);
        end

        if((pre_barrier_xacts[i].transmitted_channel == svt_axi_transaction::WRITE) &&
           !pre_barrier_xacts[i].compare_write_data(write_xact_data_stream,write_xact_wstrb_stream,read_xact_byte_stream)) begin
          `svt_xvm_error("check_pre_barrier_and_post_barrier_xact_contents",
           $sformatf("Expected contents of pre_barrier_xacts and corresponding memory read to be same, but they are not. pre_barrier xact: %0s. mem_read xact: %0s\npre_barrier_xact data: %0s\nmem read data = %0s",
           `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),`SVT_AXI_PRINT_PREFIX1(post_barrier_xacts[i]),
           pre_barrier_xacts[i].get_write_data_string(write_xact_data_stream,write_xact_wstrb_stream),pre_barrier_xacts[i].get_read_data_string(read_xact_byte_stream)));
        end
        else if((pre_barrier_xacts[i].transmitted_channel != svt_axi_transaction::WRITE) &&
                !pre_barrier_xacts[i].compare_read_data(write_xact_data_stream,read_xact_byte_stream)) begin
          `svt_xvm_error("check_pre_barrier_and_post_barrier_xact_contents",
           $sformatf("Expected contents of pre_barrier_xacts and corresponding memory read to be same, but they are not. pre_barrier xact: %0s. mem_read xact: %0s\npre_barrier_xact data: %0s\nmem read data = %0s",
           `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),`SVT_AXI_PRINT_PREFIX1(post_barrier_xacts[i]),
           pre_barrier_xacts[i].get_read_data_string(write_xact_data_stream),pre_barrier_xacts[i].get_read_data_string(read_xact_byte_stream)));
        end
        else begin
          `svt_xvm_debug("check_pre_barrier_and_post_barrier_xact_contents",
           $sformatf("Contents of pre_barrier_xacts and corresponding memory read are same. pre_barrier xact: %0s. mem_read xact: %0s\npre_barrier_xact data: %0s\nmem read data = %0s",
           `SVT_AXI_PRINT_PREFIX1(pre_barrier_xacts[i]),`SVT_AXI_PRINT_PREFIX1(post_barrier_xacts[i]),
           pre_barrier_xacts[i].get_read_data_string(write_xact_data_stream),pre_barrier_xacts[i].get_read_data_string(read_xact_byte_stream)));
        end
      end 
    end
  endfunction

  virtual function bit is_applicable(svt_configuration cfg);
    return(0);
  endfunction

endclass: svt_axi_ace_master_barrier_base_virtual_sequence 

// **************************************************************************
// ************************* BASIC LEVEL SEQUENCES *******************
// **************************************************************************

/** 
 * This sequence initiates MakeUnique transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  MakeUnique transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending Makeunique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_makeunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 

  `svt_xvm_object_utils(svt_axi_ace_master_makeunique_sequence)
  
  constraint valid_port_type {
    port_id inside {ace_ports};
  } 
  
  function new(string name = "svt_axi_ace_master_makeunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  /**
    * Initializes cachelines and sends makeunique from port "port_id"
    */
  virtual task body();
    
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::MAKEUNIQUE ,1);
      // Wait for MakeUnique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    
    end
  
  endtask: body

endclass: svt_axi_ace_master_makeunique_sequence

/** 
 * This sequence initiates Readshared transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  ReadShared transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending Readshared transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_readshared_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 
 
  `svt_xvm_object_utils(svt_axi_ace_master_readshared_sequence)
  
  constraint valid_port_type {
    port_id inside {ace_ports};
  } 
  
  function new(string name = "svt_axi_ace_master_readshared_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

/**
 * Initializes cachelines and sends readshared from port "port_id"
 */
  virtual task body();
    
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READSHARED ,1);
      // Wait for readshared transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_readshared_sequence

/** 
 * This sequence initiates ReadClean transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  ReadClean transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending ReadClean transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_readclean_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
 
  `svt_xvm_object_utils(svt_axi_ace_master_readclean_sequence)
 
  constraint valid_port_type {
    port_id inside {ace_ports};
  } 
 
  function new(string name = "svt_axi_ace_master_readclean_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
            
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READCLEAN ,1); 
      // Wait for readclean transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_readclean_sequence


/** 
 *  This sequence initiates ReadNoSnoop transaction from the ACE/ACE_LITE
 *  master specified with port_id , which can be a random port or a specific
 *  port configured by the user through uvm_config_db. 
 */

class svt_axi_ace_master_readnosnoop_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readnosnoop_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  } 
  
  function new(string name = "svt_axi_ace_master_readnosnoop_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READNOSNOOP ,0);
      // Wait for readnosnoop transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_readnosnoop_sequence

/** 
  * This sequence initiates ReadOnce transaction from the ACE/ACE-Lite master
  * specified with port_id , which can be a random port or a specific port
  * configured by the user through uvm_config_db.  ReadOnce transactions can be
  * sent only when the svt_axi_port_configuration::axi_interface_type of the
  * master corresponding to port_id is set to
  * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
  * Before sending ReadOnce transactions, cachelines of peer masters are
  * initialized to random, valid states.  Initialisation is done through front
  * door access, by sending specific transactions from the initiating master
  * (corresponding to port_id) and peer masters.  Please look up the
  * documentation of #svt_axi_cacheline_initialization for details.
  */
class svt_axi_ace_master_readonce_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readonce_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports, ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readnosnoop_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READONCE ,1);
      // Wait for readonce transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_readonce_sequence

/** 
 * This sequence initiates ReadNotSharedDirty transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  ReadNotSharedDirty transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending ReadNotSharedDirty transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_readnotshareddirty_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readnotshareddirty_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readnotshareddirty_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
    
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READNOTSHAREDDIRTY ,1);
      // Wait for readnotshareddirty transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body
 
endclass: svt_axi_ace_master_readnotshareddirty_sequence

/** 
 * This sequence initiates ReadUnique transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  ReadUnique transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending ReadUnique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_readunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readunique_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READUNIQUE ,1);
      // Wait for readunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_readunique_sequence

/** 
 * This sequence initiates CleanUnique transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  CleanUnique transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending CleanUnique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_cleanunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_cleanunique_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cleanunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::CLEANUNIQUE ,1);
      // Wait for cleanunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_cleanunique_sequence


/** 
 * This sequence initiates CleanShared transaction from the ACE/ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  CleanShared transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
 * Before sending CleanShared transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_cleanshared_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_cleanshared_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cleanshared_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::CLEANSHARED ,1);  
      // Wait for cleanshared transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_cleanshared_sequence

/** 
 * This sequence initiates CleanSharedPersist transaction from the ACE/ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  CleanSharedPersist transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
 * Before sending CleanSharedPersist transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_cleansharedpersist_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_cleansharedpersist_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cleansharedpersist_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::CLEANSHAREDPERSIST ,1);  
      // Wait for cleansharedpersist transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_cleansharedpersist_sequence

/** 
 * This sequence initiates concurrent random non-dvm transactions from first_port_id and
 * dvm transactions from dvm_port_id. These ports can be a random port or a specifc port 
 * configured by user through uvm_config_db. Based on the interface type of first_port_id, 
 * a transction type as set in first_port_xact_type is sent from first_port_id. 
 * Before sending the transactions, cachelines of peer masters are initialized to random valid states. 
 * Initialisation is done through front door access, by sending specific transactions from the 
 * initiating master (corresponding to first_port_id) and peer masters. Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_concurent_non_dvm_xacts_with_dvm_xacts_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Semephore to control the process between non dvm and multi part dvm transactions */
  protected semaphore read_channel_sema = new(1);

  /** Represents the port for sending non-DVM transactions. 
    * Valid only if send_non_dvm_xact_select is set.
    * first_port_id may be the same as dvm_port_id1 or dvm_port_id2. However,
    * if dvm_port1_multipart_select is set, first_port_id cannot be dvm_port_id1.
    * The same applies to dvm_port2_multipart_select and dvm_port_id2. This is
    * because non-DVM transactions cannot be sent between two multipart DVM
    * transactions
    * This property can be controlled via uvm_config_db. */
  rand int unsigned first_port_id;
  
  /** Represents the first dvm master port. This property can be controlled via uvm_config_db. */
  rand int dvm_port_id1 = -1;

  /** Represents the second dvm master port. This property can be controlled via uvm_config_db. */
  rand int dvm_port_id2 = -1;

  /** Represents the multipart dvm transaction selection for dvm_port_id1. 
    * Note that if the dvm_message_type selected is TLB_INVALIDATE,
    * PHYSICAL_INSTRUCTION_CACHE_INVALIDATE or VIRTUAL_INSTRUCTION_CACHE_INVALIDATE,
    * the randomized values of tlb_operation, physical_instruction_invalidate_operation and
    * virtual_instruction_invalidate_operation determine whether a DVM transaction will be
    * multipart or not. 
    * This property can be controlled via uvm_config_db. */
  rand bit dvm_port1_multipart_select;

  /** Represents the multipart dvm transaction selection for dvm_port_id2. 
    * Note that if the dvm_message_type selected is TLB_INVALIDATE,
    * PHYSICAL_INSTRUCTION_CACHE_INVALIDATE or VIRTUAL_INSTRUCTION_CACHE_INVALIDATE,
    * the randomized values of tlb_operation, physical_instruction_invalidate_operation and
    * virtual_instruction_invalidate_operation determine whether a DVM transaction will be
    * multipart or not. 
    * This property can be controlled via uvm_config_db. */
  rand bit dvm_port2_multipart_select;

  /** Sends non dvm transactions on first_port_id if set to 1, 
    * Sends only dvm messages without non dvm transactions if set to 0.
    * This property can be controlled via uvm_config_db.
    */ 
  rand bit send_non_dvm_xact_from_first_port_select;

  /**
    * Sends non-dvm transactions along with DVM transactions from dvm_port_id1
    * and dvm_port_id2. Only transactions which can be sent out without
    * initializing the cacheline are used. These transactions are WRITENOSNOOP,
    * READNOSNOOP, MAKEUNIQUE, READUNIQUE, READSHARED, READCLEAN,
    * READNOTSHAREDDIRTY, CLEANINVALID, CLEANSHARED, MAKEINVALID, WRITEUNIQUE,
    * WRITELINEUNIQUE.
    */
  rand bit send_non_dvm_xact_from_dvm_port_select;

  /**
    * Applicable when send_non_dvm_xact_from_dvm_port_select is set.
    * Indicates the number of non dvm transactions to be sent after
    * num_dvm_xacts_before_non_dvm_xact number of DVM transactions are sent
    * Once the non-dvm transactions are sent, DVM transactions are represented
    * by num_dvm_xacts_before_non_dvm_xact are sent again. 
    */
  rand int num_non_dvm_xacts_from_dvm_port;

  /**
    * Applicable when send_non_dvm_xact_from_dvm_port_select is set.
    * Indicates the number of DVM transactions to be sent before non-DVM
    * transactions are sent. Once the non-dvm transactions are sent, DVM
    * transactions as represented by the this variable are sent before
    * sending non-DVM transactions. Hence the sequence of 
    * DVM based on num_dvm_xacts_before_non_dvm_xact, non-DVM based on
    * num_non_dvm_xacts_from_dvm_port is repeated.
    */
  rand int num_dvm_xacts_before_non_dvm_xact;

  
  /** Enum to represent DVM Message type. */
  typedef enum bit [2:0] {
    TLB_INVALIDATE                        = 'h0, /**< TLB invalidate */
    BRANCH_PREDICTOR_INVALIDATE           = 'h1, /**< Branch predictor invalidate */
    PHYSICAL_INSTRUCTION_CACHE_INVALIDATE = 'h2, /**< Physical instruction cache invalidate */
    VIRTUAL_INSTRUCTION_CACHE_INVALIDATE  = 'h3, /**< Virtual instruction cache invalidate */
    HINT                                  = 'h6  /**< Hint messages */
  } dvm_message_enum;
 
  /** Enum to represent TLB INVALIDATE sub operation */
  typedef enum bit [11:0] {
    SECURE_TLB_INVALIDATE_ALL                             = 12'hA00, 
    SECURE_TLB_INVALIDATE_BY_VA                           = 12'hA01, 
    SECURE_TLB_INVALIDATE_BY_VA_LEAF_ENTRY                = 12'hA11, 
    SECURE_TLB_INVALIDATE_BY_ASID                         = 12'hA20, 
    SECURE_TLB_INVALIDATE_BY_ASID_VA                      = 12'hA21, 
    SECURE_TLB_INVALIDATE_BY_ASID_VA_LEAF_ENTRY           = 12'hA31, 
    ALL_OS_TLB_INVALIDATE_ALL                             = 12'hB00, 
    GUEST_OS_TLB_INVALIDATE_ALL_STAGE1_INVALIDATION       = 12'hB44, 
    GUEST_OS_TLB_INVALIDATE_ALL_STAGE1_AND_2_INVALIDATION = 12'hB40, 
    GUEST_OS_TLB_INVALIDATE_BY_VA                         = 12'hB41, 
    GUEST_OS_TLB_INVALIDATE_BY_VA_LEAF_ENTRY              = 12'hB51,
    GUEST_OS_TLB_INVALIDATE_BY_ASID                       = 12'hB60, 
    GUEST_OS_TLB_INVALIDATE_BY_ASID_VA                    = 12'hB61, 
    GUEST_OS_TLB_INVALIDATE_BY_ASID_VA_LEAF_ENTRY         = 12'hB71, 
    GUEST_OS_TLB_INVALIDATE_BY_IPA                        = 12'hB49, 
    GUEST_OS_TLB_INVALIDATE_BY_IPA_LEAF_ENTRY             = 12'hB59, 
    HYPERVISOR_TLB_INVALIDATE_ALL                         = 12'hF00, 
    HYPERVISOR_TLB_INVALIDATE_BY_VA                       = 12'hF01, 
    HYPERVISOR_TLB_INVALIDATE_BY_VA_LEAF_ENTRY            = 12'hF11, 
    EL3_TLB_INVALIDATE_BY_VA                              = 12'h601, 
    EL3_TLB_INVALIDATE_BY_VA_LEAF_ENTRY                   = 12'h611, 
    EL3_TLB_INVALIDATE_ALL                                = 12'h600
  } tlb_operations_enum;

  /** Enum to represent PHYSICAL INSTRUCTION INVALIDATE sub operation */
  typedef enum bit [9:0] {
    SECURE_PHYSICAL_INSTRUCTION_INVALIDATE_ALL                  = 10'h200,
    SECURE_PHYSICAL_INSTRUCTION_BY_PA_WITHOUT_VIRTUAL_INDEX     = 10'h201, 
    SECURE_PHYSICAL_INSTRUCTION_BY_PA_WITH_VIRTUAL_INDEX        = 10'h261, 
    NON_SECURE_PHYSICAL_INSTRUCTION_INVALIDATE_ALL              = 10'h300, 
    NON_SECURE_PHYSICAL_INSTRUCTION_BY_PA_WITHOUT_VIRTUAL_INDEX = 10'h301, 
    NON_SECURE_PHYSICAL_INSTRUCTION_BY_PA_WITH_VIRTUAL_INDEX    = 10'h361 
  } physical_instruction_invalidate_operations_enum;

  /** Enum to represent VIRTUAL INSTRUCTION INVALIDATE sub operation */
  typedef enum bit [11:0] {
    VIRTUAL_INSTRUCTION_INVALIDATE_ALL_SECURE_NON_SECURE = 12'h000,
    VIRTUAL_INSTRUCTION_INVALIDATE_ALL_NON_SECURE        = 12'h300,
    VIRTUAL_INSTRUCTION_SECURE_INVALIDATE_BY_ASID_VA     = 12'hA21, 
    VIRTUAL_INSTRUCTION_GUEST_OS_INVALIDATE_ALL          = 12'hB40,
    VIRTUAL_INSTRUCTION_GUEST_OS_INVALIDATE_BY_ASID_VA   = 12'hB61, 
    VIRTUAL_INSTRUCTION_HYPERVISOR_INVALIDATE_BY_VA      = 12'hF01
  } virtual_instruction_invalidate_operations_enum;
  
  /** The tlb_operation represents the tlb sub operation to be sent from test */
  rand tlb_operations_enum tlb_operation;

  /** The physical_instruction_invalidate_operation represents the physical instruction invalidate
    * sub operation to be sent from test 
    */
  rand physical_instruction_invalidate_operations_enum physical_instruction_invalidate_operation;

  /** The virtual_instruction_invalidate_operation represents the virtual instruction invalidate
    * sub operation to be sent from test
    */
  rand virtual_instruction_invalidate_operations_enum virtual_instruction_invalidate_operation;

  /** The dvm_message_type represents the dvm message to be sent from test.
    * This property can be controlled via uvm_config_db. 
    */
  rand dvm_message_enum dvm_message_type;
  
  /** Sends the dvm_message_type as dvm message if set to 1, 
    * Sends the random_dvm_message_type as dvm message if set to 0.
    * This property can be controlled via uvm_config_db.
    */
  bit dvm_message_type_select = 0;


  /** Represents the weights of first part dvm address distribution */
  int unsigned first_part_dvm_addr_bins_wt_min = 25;
  int unsigned first_part_dvm_addr_bins_wt_mid = 33;
  int unsigned first_part_dvm_addr_bins_wt_max = 34;

  /** Represents the weights of second part dvm message type distribution */
  int unsigned second_part_dvm_message_type_wt_min = 10;
  int unsigned second_part_dvm_message_type_wt_mid = 40;
  int unsigned second_part_dvm_message_type_wt_max = 50;

  /** Handles of infinite snoop response sequeunces running on each master */
  `ifdef __SVDOC__
    `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER 128
  `else
  `ifndef SVT_AXI_MAX_NUM_MASTERS_0
    `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER `SVT_AXI_MAX_NUM_MASTERS
  `else
    `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER 1
  `endif
  `endif
  /** Handle of maximum address width supported by each master */
  `ifdef SVT_AXI_MAX_ADDR_WIDTH
    `define _SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH `SVT_AXI_MAX_ADDR_WIDTH
  `endif

  /** Random coherent non-dvm transaction type for first_port_id 
    * This property can be controlled via uvm_config_db.
    */ 
  rand svt_axi_transaction::coherent_xact_type_enum first_port_xact_type;
 
  /**
    * The shareability domain of the DVM transactions to be sent
    */
  rand svt_axi_transaction::xact_shareability_domain_enum domain_type;
 
  /**
    * The dvm os type of the DVM transactions to be sent
    */
  rand svt_axi_transaction::dvm_os_enum dvm_os_select;
  
  /**
    * The dvm security type of the DVM transactions to be sent
    */
  rand svt_axi_transaction::dvm_security_enum dvm_security_select;

  /** Collects the indexes of active, participating masters with svt_axi_port_configuration::dvm_enable set */ 
  int dvm_ace_ports[$], dvm_ace_lite_ports[$];

  
  /** 
    * Handles of infinite DVM complete sequences running on each master. 
    * These wait for a DVM Sync snoop transaction and send DVM complete transactions
    */
  svt_axi_ace_master_dvm_complete_sequence dvm_complete_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER];
  
  svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER];
  `ifdef SVT_UVM_TECHNOLOGY
    uvm_component my_component;
  `elsif SVT_OVM_TECHNOLOGY
    ovm_component my_component;
  `endif
    svt_axi_system_env my_system_env;
    svt_axi_system_configuration sys_cfg;
  
  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::INNERSHAREABLE,
                        svt_axi_transaction::OUTERSHAREABLE};
  }

  constraint reasonable_ports {
    first_port_id inside {[0:(cfg.num_masters-1)]};
  }
  
  /** Enum to represent the first_port_id interface type and dvm_port_id
    * interface type.  
    */
  typedef enum {
    DVM_PORT1_ACE = 0,
    DVM_PORT1_ACE_LITE = 1,
    DVM_PORT1_ACE_DVM_PORT2_ACE = 2,
    DVM_PORT1_ACE_DVM_PORT2_ACE_LITE = 3,
    DVM_PORT1_ACE_LITE_DVM_PORT2_ACE_LITE = 4 
  } two_port_interface_types_enum;
  
  /** Represents the interface types for the first port and dvm port, 
    * selected according to the number of AXI_ACE and ACE_LITE ports collected 
    * through find_dvm_ports function
    */
  rand two_port_interface_types_enum two_port_interface_type;

  constraint valid_two_port_interface_type {
    if (dvm_ace_ports.size() < 2)
      two_port_interface_type != DVM_PORT1_ACE_DVM_PORT2_ACE;
    if (dvm_ace_lite_ports.size() < 2)
      two_port_interface_type !=  DVM_PORT1_ACE_LITE_DVM_PORT2_ACE_LITE;
    if (!dvm_ace_ports.size() || !dvm_ace_lite_ports.size())
      two_port_interface_type != DVM_PORT1_ACE_DVM_PORT2_ACE_LITE;
    if (!dvm_ace_ports.size())
      two_port_interface_type != DVM_PORT1_ACE;
    if (!dvm_ace_lite_ports.size())
      two_port_interface_type != DVM_PORT1_ACE_LITE;
    if (dvm_port1_multipart_select && dvm_port2_multipart_select &&
        (dvm_ace_ports.size() + dvm_ace_lite_ports.size() <= 2))
      send_non_dvm_xact_from_first_port_select == 0;
      
  }
  
  constraint valid_two_port_id_type {
    first_port_id inside {ace_ports,ace_lite_ports};
    if (dvm_port1_multipart_select)
      first_port_id != dvm_port_id1;
    if (dvm_port2_multipart_select)
      first_port_id != dvm_port_id2;
    if (two_port_interface_type == DVM_PORT1_ACE_DVM_PORT2_ACE) {
      dvm_port_id1 inside {dvm_ace_ports}; 
      dvm_port_id2 inside {dvm_ace_ports};
      dvm_port_id1 != dvm_port_id2;
    } else if (two_port_interface_type == DVM_PORT1_ACE_DVM_PORT2_ACE_LITE) {
      dvm_port_id1 inside {dvm_ace_ports}; 
      dvm_port_id2 inside {dvm_ace_lite_ports};
      dvm_port_id1 != dvm_port_id2;
    } else if (two_port_interface_type == DVM_PORT1_ACE_LITE_DVM_PORT2_ACE_LITE) {
      dvm_port_id1 inside {dvm_ace_lite_ports};
      dvm_port_id2 inside {dvm_ace_lite_ports};
      dvm_port_id1 != dvm_port_id2;
    } else if (two_port_interface_type == DVM_PORT1_ACE) {
      dvm_port_id1 inside {dvm_ace_ports};
      dvm_port_id2 == -1;
    } else if (two_port_interface_type == DVM_PORT1_ACE_LITE) {
      dvm_port_id1 inside {dvm_ace_lite_ports};
      dvm_port_id2 == -1;
    }
  }

  constraint reasonable_coherent_xact_type {  
    foreach(cfg.master_cfg[i]) {
      if (i == first_port_id) {   
        if (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
          first_port_xact_type inside {svt_axi_transaction::READONCE,
			      svt_axi_transaction::READCLEAN,
				    svt_axi_transaction::READNOTSHAREDDIRTY,
				    svt_axi_transaction::READSHARED,
				    svt_axi_transaction::READUNIQUE,
				    svt_axi_transaction::MAKEUNIQUE,
				    svt_axi_transaction::CLEANUNIQUE,
				    svt_axi_transaction::CLEANSHARED,
				    svt_axi_transaction::CLEANINVALID,
				    svt_axi_transaction::MAKEINVALID,
				    svt_axi_transaction::WRITEUNIQUE,
				    svt_axi_transaction::WRITELINEUNIQUE};
        }
        else {
          first_port_xact_type inside {svt_axi_transaction::READONCE,
				    svt_axi_transaction::CLEANINVALID,
				    svt_axi_transaction::MAKEINVALID,
				    svt_axi_transaction::CLEANSHARED,
				    svt_axi_transaction::WRITEUNIQUE,
				    svt_axi_transaction::WRITELINEUNIQUE};
        }
      }
    }
  }  
 
  constraint reasonable_num_non_dvm_xacts_from_dvm_port {
    num_non_dvm_xacts_from_dvm_port inside {[1:5]};
  }

  constraint reasonable_num_dvm_xacts_before_non_dvm_xact {
    num_dvm_xacts_before_non_dvm_xact inside {[1:5]};
  }
 

     
  /*constraint reasonable_disable_multipart_dvm {
    if (
         (dvm_port_id1 != -1) && (dvm_port1_multipart_select == 0) ||
         (dvm_port_id2 != -1) && (dvm_port2_multipart_select == 0) 
       ) {
     
    }
  }
  */
  `ifdef SVT_UVM_TECHNOLOGY
    `svt_xvm_object_utils(svt_axi_ace_concurent_non_dvm_xacts_with_dvm_xacts_sequence)
  `elsif SVT_OVM_TECHNOLOGY
    `ovm_object_utils_begin(svt_axi_ace_concurent_non_dvm_xacts_with_dvm_xacts_sequence) 
    `ovm_field_enum(dvm_message_enum,dvm_message_type, OVM_ALL_ON) 
    `ovm_field_enum(svt_axi_transaction::coherent_xact_type_enum,first_port_xact_type, OVM_ALL_ON) 
    `ovm_object_utils_end 
  `endif
  
  function new(string name = "svt_axi_ace_concurent_non_dvm_xacts_with_dvm_xacts_sequence");
    super.new(name);
  endfunction

  function void pre_randomize();
    super.pre_randomize();
    find_dvm_ports(cfg);
  endfunction

  task pre_body();
    bit status,status0,status1,status2, multipart_select;
    bit err_status1, err_status2;
    int dvm_port_id;
    super.pre_body();
  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_port1_multipart_select", dvm_port1_multipart_select);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_port2_multipart_select", dvm_port2_multipart_select);
    status = uvm_config_db#(dvm_message_enum)::get(null, get_full_name(), "dvm_message_type", dvm_message_type);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_message_type_select", dvm_message_type_select);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "send_non_dvm_xact_from_first_port_select", send_non_dvm_xact_from_first_port_select);
    status = uvm_config_db#(svt_axi_transaction::coherent_xact_type_enum)::get(null, get_full_name(), "first_port_xact_type", first_port_xact_type);
    status0 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_id", first_port_id);
    status1 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_port_id1", dvm_port_id1);
    status2 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_port_id2", dvm_port_id2);
    err_status1 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "dvm_port_id", dvm_port_id);
    err_status2 = uvm_config_db#(int unsigned)::get(null, get_full_name(), "multipart_select", multipart_select);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "num_non_dvm_xacts_from_dvm_port", num_non_dvm_xacts_from_dvm_port);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "num_dvm_xacts_before_non_dvm_xact", num_dvm_xacts_before_non_dvm_xact);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_part_dvm_addr_bins_wt_min", first_part_dvm_addr_bins_wt_min);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_part_dvm_addr_bins_wt_mid", first_part_dvm_addr_bins_wt_mid);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_part_dvm_addr_bins_wt_max", first_part_dvm_addr_bins_wt_max);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_min", second_part_dvm_message_type_wt_min);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_mid", second_part_dvm_message_type_wt_mid);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_max", second_part_dvm_message_type_wt_max);
  `elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".dvm_port1_multipart_select"}, dvm_port1_multipart_select);
    status = m_sequencer.get_config_int({get_type_name(), ".dvm_port2_multipart_select"}, dvm_port2_multipart_select);
    `ifdef QUESTA
      status = m_sequencer.get_config_int({get_type_name(),".dvm_message_type"}, int'(dvm_message_type));
      status = m_sequencer.get_config_int({get_type_name(), ".first_port_xact_type"}, int'(first_port_xact_type));
    `else 
      status = m_sequencer.get_config_int({get_type_name(),".dvm_message_type"}, dvm_message_type);
      status = m_sequencer.get_config_int({get_type_name(), ".first_port_xact_type"}, first_port_xact_type);
    `endif
    status = m_sequencer.get_config_int({get_type_name(), ".dvm_message_type_select"}, dvm_message_type_select);
    status = m_sequencer.get_config_int({get_type_name(), ".send_non_dvm_xact_from_first_port_select"}, send_non_dvm_xact_from_first_port_select);    
    status0 = m_sequencer.get_config_int({get_type_name(), ".first_port_id"}, first_port_id);
    status1 = m_sequencer.get_config_int({get_type_name(), ".dvm_port_id1"}, dvm_port_id1);
    status2 = m_sequencer.get_config_int({get_type_name(), ".dvm_port_id2"}, dvm_port_id2);
    err_status1 = m_sequencer.get_config_int({get_type_name(), ".dvm_port_id"}, dvm_port_id);
    err_status2 = m_sequencer.get_config_int({get_type_name(), ".multipart_select"}, multipart_select);
    status = m_sequencer.get_config_int({get_type_name(), ".num_non_dvm_xacts_from_dvm_port"}, num_non_dvm_xacts_from_dvm_port);
    status = m_sequencer.get_config_int({get_type_name(), ".num_dvm_xacts_before_non_dvm_xact"}, num_dvm_xacts_before_non_dvm_xact);
    status = m_sequencer.get_config_int({get_type_name(), ".first_part_dvm_addr_bins_wt_min"}, first_part_dvm_addr_bins_wt_min);
    status = m_sequencer.get_config_int({get_type_name(), ".first_part_dvm_addr_bins_wt_mid"}, first_part_dvm_addr_bins_wt_mid);
    status = m_sequencer.get_config_int({get_type_name(), ".first_part_dvm_addr_bins_wt_max"}, first_part_dvm_addr_bins_wt_max);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_min"}, second_part_dvm_message_type_wt_min);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_mid"}, second_part_dvm_message_type_wt_mid);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_max"}, second_part_dvm_message_type_wt_max);
  `endif
    `svt_xvm_debug("body", $sformatf("first_port_id is 'd%0d as a result of %0s.", first_port_id, status0 ? "config DB" : "randomization"));
    `svt_xvm_debug("body", $sformatf("dvm_port_id1 is 'd%0d as a result of %0s.", dvm_port_id1, status1 ? "config DB" : "randomization"));
    `svt_xvm_debug("body", $sformatf("dvm_port_id2 is 'd%0d as a result of %0s.", dvm_port_id2, status2 ? "config DB" : "randomization"));
    if (err_status1)
      `svt_error("body", "dvm_port_id has been passed through config_db. This is deprecated. Please use dvm_port_id1 and dvm_port_id2");
    if (err_status2)
      `svt_error("body", "multipart_select has been passed through config_db. This is deprecated. Please use dvm_port1_multipart_select and dvm_port2_multipart_select");
  endtask: pre_body

  function void find_dvm_ports(svt_axi_system_configuration cfg);
     foreach(cfg.master_cfg[i]) begin
       if (
             (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
             (cfg.master_cfg[i].dvm_enable == 1) &&
             (cfg.master_cfg[i].is_active) &&
             (cfg.is_participating(i))
          ) begin
         dvm_ace_ports.push_back(i);
         `svt_xvm_note("find_dvm_ports", $sformatf("dvm_ace_ports = 'd%0d",i)); end
     end
     foreach(cfg.master_cfg[i]) begin
       if (
             (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
             (cfg.master_cfg[i].dvm_enable == 1) &&
             (cfg.master_cfg[i].is_active) &&
             (cfg.is_participating(i))
          ) begin
         dvm_ace_lite_ports.push_back(i);
          `svt_xvm_note("find_dvm_ports", $sformatf("dvm_ace_lite_ports = 'd%0d",i)); end
     end
     if (!dvm_ace_ports.size() && !dvm_ace_lite_ports.size()) begin
       `svt_xvm_fatal("find_dvm_ports", "There are no ACE ports or ACE-Lite masters with dvm_enable in the system and therefore this sequence cannot be run. Please ensure that there is atleast one dvm_enable asserted ACE or ACE-Lite master in the system");
     end
  endfunction
  
  virtual function bit transaction_type_check();
    if (send_non_dvm_xact_from_first_port_select) begin
      if (dvm_ace_ports.size() + dvm_ace_lite_ports.size() <= (dvm_port1_multipart_select + dvm_port2_multipart_select))
        `svt_error("transaction_type_check", $sformatf("If send_non_dvm_xact_from_first_port_select is set, the total number of DVM capable masters must be more than that of the masters for which dvm multi-part is being requested. num_dvm_ace_ports = 'd%0d. num_dvm_ace_lite_ports = 'd%0d. dvm_port1_multipart_select = 'b%0b.   dvm_port2_multipart_select = 'b%0b", dvm_ace_ports.size(), dvm_ace_lite_ports.size(), dvm_port1_multipart_select, dvm_port2_multipart_select)); 
    end
    if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE)
      begin
       if (first_port_xact_type != svt_axi_transaction::READONCE &&
				 first_port_xact_type !=    svt_axi_transaction::CLEANSHARED &&
				 first_port_xact_type !=    svt_axi_transaction::CLEANINVALID &&
				 first_port_xact_type !=    svt_axi_transaction::MAKEINVALID &&
				 first_port_xact_type !=    svt_axi_transaction::WRITEUNIQUE &&
				 first_port_xact_type !=    svt_axi_transaction::WRITELINEUNIQUE) begin
         `svt_xvm_warning("transaction_type_check", "Invalid transaction type selected for port type specified, valid transaction should be non-cached load or non-cached store or cmo types which can be sent from ACE_LITE master");
         return 0;
         end
       else 
         return 1;
      end
    else
      return 1;
  endfunction
    
  virtual task send_dvm_sequence(int port_id, int num_of_dvm_xacts, bit [11:0] dvm_sub_operation,bit is_multipart);
    svt_axi_master_transaction tr1, tr2;
    bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  _multi_dvm_first_txn_id;
    dvm_message_enum random_dvm_message_type;
    dvm_message_enum dvm_message_type_arr[5] = {TLB_INVALIDATE, BRANCH_PREDICTOR_INVALIDATE, PHYSICAL_INSTRUCTION_CACHE_INVALIDATE, VIRTUAL_INSTRUCTION_CACHE_INVALIDATE, HINT};
    bit [2:0] dvm_count,send_dvm_message;
    bit [2:0] sync_message = 'h4;
    bit multipart_sync_select = 0;
    int expected_dvm_completes = 0;
    int received_dvm_completes = 0;
    bit _multipart_select;
    int num_dvms_before_sync;
    svt_axi_master_transaction dvm_xacts[$],non_dvm_xacts[$];
    _multipart_select = is_multipart;
    //num_of_dvm_xacts = 500;
    num_dvms_before_sync = $urandom_range(1,5);

    for (int seq_length = 0; seq_length < num_of_dvm_xacts; seq_length++) begin 
      //Condition set sets the random_dvm_message_type as dvm_message_type if it is selected by the user from test
      //else sets any one random value of dvm_message_type_arr.
      if (dvm_message_type_select) begin
        random_dvm_message_type = dvm_message_type;
      end
      else begin
        dvm_message_type_arr.shuffle();
        random_dvm_message_type = dvm_message_type_arr[0]; 
       end
      
      //Condition sets the send_dvm_message as sync_message after certain number of DVM operations.
      if(dvm_count < num_dvms_before_sync)
      begin
        send_dvm_message = random_dvm_message_type;
        dvm_count++;
        if(_multipart_select)
          multipart_sync_select = $urandom_range(0,1);
      end
      else if(dvm_count == num_dvms_before_sync)
      begin
        send_dvm_message = sync_message;
        num_dvms_before_sync = $urandom_range(1,5);
        dvm_count = 0;
        if(_multipart_select)
          multipart_sync_select = 0;
      end

        
      `svt_xvm_note("send_dvm_sequence", $sformatf("dvm_port_id = 'd%0d. random_dvm_message_type : %0s, dvm_message_type : 'd%0d, multipart_select : 'd%0d, num_of_dvm_xacts = 'd%0d,send_dvm_message : 'd%0d, first_port_xact_type = %0s,dvm_message_type_select = 'd%0d,two_port_interface_type = %0s",port_id,random_dvm_message_type.name(),dvm_message_type,_multipart_select,num_of_dvm_xacts,send_dvm_message,first_port_xact_type,dvm_message_type_select,two_port_interface_type.name()));

      `svt_xvm_create_on(tr1, p_sequencer.master_sequencer[port_id])
      tr1.port_cfg = sys_cfg.master_cfg[port_id];
//vcs-vip-protect
`protected
.1?OE.4/B7(Ze&=^?VgD,feWHg_X^(fT/U73?STEf>9H@HeY:aN,4)5,Z2c&MN#g
0(a>YO@<C?cEV<FV13R:A1a>9DD/ePO^AEY-EbJJ-8&FSR2&d[=K)df@__5,AC44
>/bd-:(eG:B?D7>BTb0^QFa>4$
`endprotected

      void'(tr1.randomize() with {
         tr1.addr[14:12] == send_dvm_message;
         if(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH == 64)
           tr1.addr[(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH - 1) : 16] dist {['h0:{16'hFFFF,28'hFFFFFFF}]:/first_part_dvm_addr_bins_wt_max,[{16'h1000,32'h00000000}:{16'h8FFF,32'hFFFFFFFF}]:/first_part_dvm_addr_bins_wt_mid, [{16'h9000,32'h00000000}:{16'hFFFF,32'hFFFFFFFF}]:/first_part_dvm_addr_bins_wt_mid};  
         if(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH == 56)
           tr1.addr[(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH - 1) : 16] dist {['h0:{16'hFFFF,20'hFFFFF}]:/first_part_dvm_addr_bins_wt_max,[{16'h1000,24'h000000}:{16'h8FFF,24'hFFFFFF}]:/first_part_dvm_addr_bins_wt_mid, [{16'h9000,24'h000000}:{16'hFFFF,24'hFFFFFF}]:/first_part_dvm_addr_bins_wt_mid};
         if(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH == 48)
           tr1.addr[(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH - 1) : 16] dist {['h0:'hFFFFFFF]:/first_part_dvm_addr_bins_wt_max,['h10000000:'h8FFFFFFF]:/first_part_dvm_addr_bins_wt_mid, ['h90000000:'hFFFFFFFF]:/first_part_dvm_addr_bins_wt_mid};
         if(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH == 44)
           tr1.addr[(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH - 1) : 16] dist {['h0:'hFFFFFF]:/first_part_dvm_addr_bins_wt_max,['h1000000:'h8FFFFFF]:/first_part_dvm_addr_bins_wt_mid, ['h9000000:'hFFFFFFF]:/first_part_dvm_addr_bins_wt_mid};
         if(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH == 40)
           tr1.addr[(`_SVT_AXI_DVM_SEQ_MAX_ADDR_WIDTH - 1) : 16] dist {['h0:'hFFFFF]:/first_part_dvm_addr_bins_wt_max,['h100000:'h8FFFFF]:/first_part_dvm_addr_bins_wt_mid, ['h900000:'hFFFFFF]:/first_part_dvm_addr_bins_wt_mid};

         if(send_dvm_message != sync_message) {
           if (dvm_message_type == 0 || //TLB_INVALIDATE |
               dvm_message_type == 2 || // PHYSICAL_INSTRUCTION_CACHE_INVALIDATE  
               dvm_message_type == 3 ) // VIRTUAL_INSTRUCTION_CACHE_INVALIDATE 
             tr1.addr[11:0] == dvm_sub_operation[11:0];
           else
             tr1.addr[0] == multipart_sync_select;
         }
         tr1.data_before_addr == 0;
         tr1.xact_type == svt_axi_transaction::COHERENT;
         tr1.coherent_xact_type == svt_axi_transaction::DVMMESSAGE;
         if(tr1.addr[6] == 1) {
           tr1.addr[23:16] dist {['h0:'h3F]:/first_part_dvm_addr_bins_wt_max,['h40:'h7F]:/first_part_dvm_addr_bins_wt_mid,['h80:'hBF]:/first_part_dvm_addr_bins_wt_mid, ['hC0:'hFF]:/first_part_dvm_addr_bins_wt_mid};
         }

      });
      _multi_dvm_first_txn_id = tr1.id;
      multipart_sync_select = tr1.addr[0];

      if(multipart_sync_select && send_non_dvm_xact_from_first_port_select) 
        read_channel_sema.get();
      `svt_xvm_send(tr1)
      dvm_xacts.push_back(tr1);
 
      if(multipart_sync_select) begin
    
        `svt_xvm_create_on(tr2, p_sequencer.master_sequencer[port_id])
         tr2.port_cfg = sys_cfg.master_cfg[port_id];
//vcs-vip-protect
`protected
W5OSS74XZ9?&;d6Vg@KfBg0>2RSH9?)UFC3PFDXG8C2L]QHK;Qc;7)\e5\5I7Z3P
_FgC?0Xd]WdCDST(_[8\/LZQIA;=B2a9T3^>J2fBe?<UAJb[:3EU0DI:/UK-0#1O
2#]9?GT#Fg]b/ZBI+#\2O0ZQ7$
`endprotected

         tr2.set_multipart_dvm_flag();
         void'(tr2.randomize() with {
         tr2.id == _multi_dvm_first_txn_id;
         tr2.addr[0] == 0;
         //tr2.addr[14:12] dist {4:=second_part_dvm_message_type_wt_mid, [0:3]:/second_part_dvm_message_type_wt_max, 6:=second_part_dvm_message_type_wt_min};
         tr2.addr[14:12] == send_dvm_message;
         tr2.data_before_addr == 0;
         tr2.xact_type == svt_axi_transaction::COHERENT;
         tr2.coherent_xact_type == svt_axi_transaction::DVMMESSAGE;

           if(tr2.addr[14:12] == 0){
               dvm_sub_operation == tlb_operation;
               tr2.addr[11:1] == dvm_sub_operation[11:1];
              }
            if(tr2.addr[14:12] == 2){
               dvm_sub_operation == physical_instruction_invalidate_operation;
               tr2.addr[11:1] == dvm_sub_operation[11:1];  }
            if(tr2.addr[14:12] == 3){
               dvm_sub_operation == virtual_instruction_invalidate_operation ;
               tr2.addr[11:1] == dvm_sub_operation[11:1]; }

            });
 
        `svt_xvm_send(tr2)
        dvm_xacts.push_back(tr2);
        if(send_non_dvm_xact_from_first_port_select)
          read_channel_sema.put();
      end
      
      if(send_dvm_message == sync_message)
      begin
        expected_dvm_completes++;
        fork 
        begin
          wait_for_dvm_complete( snoop_resp_seq, port_id );
          received_dvm_completes++;  
        end
        join_none
        tr1.wait_for_transaction_end();
          if(multipart_sync_select)
            tr2.wait_for_transaction_end();
      end

      if (send_non_dvm_xact_from_dvm_port_select && (seq_length > num_dvm_xacts_before_non_dvm_xact) && (seq_length%num_dvm_xacts_before_non_dvm_xact==0)) begin
        for (int j = 0; j < num_non_dvm_xacts_from_dvm_port; j++) begin
          svt_axi_master_transaction non_dvm_tr;
          `svt_xvm_create_on(non_dvm_tr, p_sequencer.master_sequencer[port_id])
          non_dvm_tr.port_cfg = sys_cfg.master_cfg[port_id];
          void'(non_dvm_tr.randomize() with {
             non_dvm_tr.data_before_addr == 0;
             non_dvm_tr.xact_type == svt_axi_transaction::COHERENT;
             non_dvm_tr.coherent_xact_type inside {svt_axi_transaction::WRITENOSNOOP, svt_axi_transaction::READNOSNOOP, svt_axi_transaction::MAKEUNIQUE, svt_axi_transaction::READUNIQUE, svt_axi_transaction::READSHARED, svt_axi_transaction::READNOTSHAREDDIRTY, svt_axi_transaction::READCLEAN, svt_axi_transaction::READONCE, svt_axi_transaction::WRITEUNIQUE, svt_axi_transaction::WRITELINEUNIQUE};
             non_dvm_tr.atomic_type != svt_axi_transaction::EXCLUSIVE;
          });
          `svt_xvm_send(non_dvm_tr)
          non_dvm_xacts.push_back(non_dvm_tr);
        end
      end
    end
    foreach (dvm_xacts[i]) begin
      `svt_xvm_debug("send_dvm_sequence",{`SVT_AXI_PRINT_PREFIX1(dvm_xacts[i]), "Waiting for DVM transaction to end"}); 
      dvm_xacts[i].wait_for_transaction_end();
      `svt_xvm_debug("send_dvm_sequence",{`SVT_AXI_PRINT_PREFIX1(dvm_xacts[i]), "Transaction ended"}); 
    end
    `svt_xvm_debug("send_dvm_sequence",$sformatf("Waiting for total 'd%0d DVM COMPLETE snoops to be received on port 'd%0d. Received 'd%0d so far, waiting for remaining ones",expected_dvm_completes, port_id, received_dvm_completes));
    wait (expected_dvm_completes == received_dvm_completes);
    `svt_xvm_debug("send_dvm_sequence",$sformatf("All pending DVM COMPLETE snoops are received on port 'd%0d", port_id));
    foreach (non_dvm_xacts[i]) begin
      `svt_xvm_debug("send_dvm_sequence",{`SVT_AXI_PRINT_PREFIX1(non_dvm_xacts[i]), "Waiting for non-DVM transaction to end"}); 
      non_dvm_xacts[i].wait_for_transaction_end();
      `svt_xvm_debug("send_dvm_sequence",{`SVT_AXI_PRINT_PREFIX1(non_dvm_xacts[i]), "Transaction ended"}); 
    end
  endtask

  virtual task wait_for_dvm_complete( svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[], int port_id );
    `SVT_DATA_BASE_OBJECT_TYPE ev_xact;
    svt_axi_snoop_transaction snoop_xact;

    `svt_xvm_note("wait_for_dvm_complete",$psprintf("Waiting for DVM COMPLETE on master 'd%0d",port_id));
    `protected
[7-VWedeQgDGYe&8,DE=E[TEC(W=7X\2(UP?/5AJ]]A6/SDWYf+7-)B1^2^N\FP:
eU@:COWD6VQXVR5PR@5>,VgTKFDT6F^2b3[gT_[#+cU2+S_SN9f=SZJM,c_6\K)\
A6>(5Z&bC6DCZG;bPBF)60=(Uf6DYFEF;-ZQSOIN:eOd)O.K^(b9CTJMM$
`endprotected

    if (!$cast(snoop_xact,ev_xact)) begin
      `svt_xvm_fatal("wait_for_dvm_complete","Transaction obtained through EVENT_DVM_COMPLETE_XACT is not of type svt_axi_snoop_transaction");
    end
    else begin
      `svt_xvm_note("wait_for_dvm_complete",$psprintf("Received DVM COMPLETE %0s on master 'd%0d. Waiting for it to complete...",`SVT_AXI_ACE_PRINT_PREFIX(snoop_xact),port_id));
      wait (
             (snoop_xact.snoop_resp_status == svt_axi_snoop_transaction::ACCEPT) ||
             (snoop_xact.snoop_resp_status == svt_axi_snoop_transaction::ABORTED) 
           );
      `svt_xvm_note("wait_for_dvm_complete",$psprintf("Received DVM COMPLETE %0s on master 'd%0d is now complete.",`SVT_AXI_ACE_PRINT_PREFIX(snoop_xact),port_id));
    end
  endtask

  virtual task start_snoop_response_seq_for_dvm(int port_id, svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER] );
    void'(snoop_resp_seq[port_id].randomize());
    `svt_xvm_note("start_snoop_response_seq_for_dvm", $sformatf("Stopping existing snoop sequences on snoop sequencer 'd%0d to start dvm specific sequence of type svt_axi_ace_master_snoop_response_sequence('d%0d) as this virtual sequence requires a snoop sequence of this type",port_id, snoop_resp_seq[port_id]));
    my_system_env.master[port_id].snoop_sequencer.stop_sequences();

    fork begin
      snoop_resp_seq[port_id].start(my_system_env.master[port_id].snoop_sequencer);
    end
    join_none

    if (sys_cfg.master_cfg[port_id].auto_gen_dvm_complete_enable == 0) begin
      dvm_complete_seq[port_id] = new($sformatf("dvm_complete_seq['d%0d]",port_id));
      `svt_xvm_create_on(dvm_complete_seq[port_id], p_sequencer.master_sequencer[port_id])
      dvm_complete_seq[port_id].snoop_resp_seq = snoop_resp_seq[port_id];
      `ifdef SVT_UVM_TECHNOLOGY
      `ifdef SVT_UVM_12_OR_HIGHER 
      dvm_complete_seq[port_id].parent_starting_phase = get_starting_phase();
      `else
      dvm_complete_seq[port_id].parent_starting_phase = starting_phase;
      `endif
      `endif
      void'(dvm_complete_seq[port_id].randomize()); 
      dvm_complete_seq[port_id].start(p_sequencer.master_sequencer[port_id]);
    end
  endtask

  virtual task body();
    bit status;
    int dvm_sequence_length = sequence_length;
    bit [11:0] dvm_sub_operation;
    svt_configuration base_cfg;
    port_id = first_port_id;    
    
    p_sequencer.get_cfg(base_cfg);
    if (!$cast(sys_cfg, base_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_system_configuration class");
    end
    my_component = p_sequencer.get_parent();
    if (!$cast(my_system_env,my_component)) begin
      `svt_xvm_fatal("body", "Expected parent of svt_axi_system_sequencer to be of type svt_axi_system_env, but it is not");
    end
    this.set_response_queue_depth(-1);
    // Mechanism to always disable sending of DVM from two masters concurrently 
`ifdef SVT_AXI_DISABLE_DVM_SEQ_FROM_TWO_PORTS
    dvm_port_id2 = -1;
`endif
    
    if (transaction_type_check())
      begin
      super.body(); 
      `svt_xvm_note("body", "Entered...");
     if (dvm_message_type_select) begin
        if (dvm_message_type == TLB_INVALIDATE)
          dvm_sub_operation = tlb_operation;
        else if (dvm_message_type == PHYSICAL_INSTRUCTION_CACHE_INVALIDATE)
          dvm_sub_operation = physical_instruction_invalidate_operation;
        else if (dvm_message_type == VIRTUAL_INSTRUCTION_CACHE_INVALIDATE)
          dvm_sub_operation = virtual_instruction_invalidate_operation;
        if (dvm_message_type == TLB_INVALIDATE || 
            dvm_message_type ==  PHYSICAL_INSTRUCTION_CACHE_INVALIDATE || 
            dvm_message_type == VIRTUAL_INSTRUCTION_CACHE_INVALIDATE) begin
          dvm_port1_multipart_select = dvm_sub_operation[0];
          dvm_port2_multipart_select = dvm_sub_operation[0];
        end
      end

      foreach (my_system_env.master[i]) begin
        if (
             (sys_cfg.master_cfg[i].is_active == 1) &&
             (
               (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) ||
               (
                 (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
                 sys_cfg.master_cfg[i].dvm_enable
               )
             )
           ) begin
          `svt_xvm_create_on(snoop_resp_seq[i], my_system_env.master[i].snoop_sequencer)
          start_snoop_response_seq_for_dvm(i, snoop_resp_seq);
        end
      end

      /** Get the semaphore to lock the channel until initialisation is complete
        * before sending DVM transactions
        */ 
      if (
           send_non_dvm_xact_from_first_port_select && 
           (dvm_port1_multipart_select || dvm_port2_multipart_select)
         )
        read_channel_sema.get();
      fork
      begin
       if(send_non_dvm_xact_from_first_port_select) begin
         svt_axi_ace_master_base_sequence first_port_seq;
         `svt_xvm_create_on(first_port_seq, p_sequencer.master_sequencer[first_port_id])
         first_port_seq.assign_xact_weights(first_port_xact_type);
         first_port_seq.initialize_cachelines = 1;
         first_port_seq.addr_mode = svt_axi_ace_master_base_sequence::RANDOM_ADDR_MODE;
         first_port_seq.generate_only_shareable_domain = 1;
         void'(first_port_seq.randomize with {use_directed_addr == 0;sequence_length==local::dvm_sequence_length;});  
         if(dvm_port1_multipart_select || dvm_port2_multipart_select) begin
           fork
           begin
             first_port_seq.start(p_sequencer.master_sequencer[first_port_id]);
           end
           begin
             `svt_xvm_debug("body", "Waiting for cacheline initialization to be done"); 
             @first_port_seq.cacheline_init_done;
             `svt_xvm_debug("body", "Cacheline initialization is done"); 
           end
           join
           // Initialization happens across all ports. Keep the semaphore until initialization is done.
           // The port on which these transaction are sent are not same as dvm_port_id1 or dvm_port_id2
           read_channel_sema.put();
           first_port_seq.wait_for_active_xacts_to_end();
         end
         else begin
           first_port_seq.start(p_sequencer.master_sequencer[first_port_id]);
           `svt_xvm_debug("body", "first_port_seq started. Waiting for active transactions to end"); 
           first_port_seq.wait_for_active_xacts_to_end();
           `svt_xvm_debug("body", "Active transactions on first_port_seq have ended");
         end
         `svt_xvm_note("body",$sformatf("All non-DVM transactions on master are now complete on port 'd%0d", first_port_id));
       end
       else
         `svt_xvm_note("body", "Sending only DVM messages because send_non_dvm_xact_from_first_port_select is set to 0"); 
      end
      begin
       send_dvm_sequence(dvm_port_id1,dvm_sequence_length,dvm_sub_operation,dvm_port1_multipart_select);
       `svt_xvm_note("body",$sformatf("All DVM COMPLETE transactions on master are now complete on port 'd%0d", dvm_port_id1));
      end
      begin
       if (dvm_port_id2 != -1) begin
         send_dvm_sequence(dvm_port_id2,dvm_sequence_length,dvm_sub_operation,dvm_port2_multipart_select);
         `svt_xvm_note("body",$sformatf("All DVM COMPLETE transactions on master are now complete on port 'd%0d", dvm_port_id2));
       end
      end
      join
      `svt_xvm_note("body","All DVM COMPLETE snoop transactions on all masters are now complete on all ports");
    end
  endtask : body
endclass : svt_axi_ace_concurent_non_dvm_xacts_with_dvm_xacts_sequence

/** 
 * This sequence initiates CleanInvalid transaction from the ACE/ACE-Lite
 * master specified with port_id , which can be a random port or a specific
 * port configured by the user through uvm_config_db.  CleanInvalid
 * transactions can be sent only when the
 * svt_axi_port_configuration::axi_interface_type of the master corresponding
 * to port_id is set to svt_axi_port_configuration::AXI_ACE or
 * svt_axi_port_configuration::ACE_LITE.  Before sending CleanInvalid
 * transactions, cachelines of peer masters are initialized to random, valid
 * states.  Initialisation is done through front door access, by sending
 * specific transactions from the initiating master (corresponding to port_id)
 * and peer masters.  Please look up the documentation of
 * #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_cleaninvalid_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_cleaninvalid_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cleaninvalid_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::CLEANINVALID ,1);
      // Wait for cleaninvalid transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_cleaninvalid_sequence

/** 
 * This sequence initiates MakeInvalid transaction from the ACE/ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  MakeInvalid transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
 * Before sending MakeInvalid transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_makeinvalid_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_makeinvalid_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_makeinvalid_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::MAKEINVALID ,1);
      // Wait for makeinvalid transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_makeinvalid_sequence


/** This sequence initiates WriteNoSnoop transaction from the ACE/ACE_Lite
 * master specified with port_id , which can be a random port or a specific
 * port configured by the user through uvm_config_db. 
 */
class svt_axi_ace_master_writenosnoop_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writenosnoop_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writenosnoop_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITENOSNOOP ,0);
      // Wait for writenosnoop transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writenosnoop_sequence

 /** 
 * This sequence initiates WriteUnique transaction from the ACE/ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  WriteUnique transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
 * Before sending WriteUnique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeunique_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITEUNIQUE ,1);
      // Wait for writeunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writeunique_sequence

/** 
 * This sequence initiates WriteLineUnique transaction from the ACE/ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  WriteLineUnique transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
 * Before sending WriteLineUnique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writelineunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writelineunique_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports, ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writelineunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITELINEUNIQUE ,1);
      // Wait for writelineunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writelineunique_sequence

`ifdef  SVT_ACE5_ENABLE
 /** 
 * This sequence initiates WriteUniqueptlstash transaction from the ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  writeuniqueptlstash transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::ACE_LITE and svt_axi_port_configuration::ace_version is set
 * to svt_axi_port_configuration::ACE_VERSION_2_0 and svt_axi_port_configuration::cache_stashing_enable
 * is set to 1.
 * Before sending writeuniqueptlstash transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeuniqueptlstash_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeuniqueptlstash_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeuniqueptlstash_sequence");
    super.new(name);
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITEUNIQUEPTLSTASH ,1);
      // Wait for writeuniqueptlstash transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writeuniqueptlstash_sequence
 /** 
 * This sequence initiates stashonceunique transaction from the ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  stashonceunique transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::ACE_LITE and svt_axi_port_configuration::ace_version is set
 * to svt_axi_port_configuration::ACE_VERSION_2_0 and svt_axi_port_configuration::cache_stashing_enable
 * is set to 1.
 * Before sending stashonceunique transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_stashonceunique_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_stashonceunique_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_stashonceunique_sequence");
    super.new(name);
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::STASHONCEUNIQUE ,1);
      // Wait for stashonceunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_stashonceunique_sequence
 /** 
 * This sequence initiates stashonceshared transaction from the ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  stashonceshared transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to
 * svt_axi_port_configuration::ACE_LITE and svt_axi_port_configuration::ace_version is set
 * to svt_axi_port_configuration::ACE_VERSION_2_0 and svt_axi_port_configuration::cache_stashing_enable
 * is set to 1.
 * Before sending stashonceshared transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_stashonceshared_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_stashonceshared_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_stashonceshared_sequence");
    super.new(name);
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::STASHONCESHARED ,1);
      // Wait for stashonceunique transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_stashonceshared_sequence

/** 
 * This sequence initiates writeuniquefullstash transaction from the ACE-Lite master
 * specified with port_id , which can be a random port or a specific port
 * configured by the user through uvm_config_db.  writeuniquefullstash transactions can
 * be sent only when the svt_axi_port_configuration::axi_interface_type of the
 * master corresponding to port_id is set to svt_axi_port_configuration::ACE_LITE and
 * svt_axi_port_configuration::ace_version is set to svt_axi_port_configuration::ACE_VERSION_2_0 and svt_axi_port_configuration::cache_stashing_enable
 * is set to 1.
 * Before sending writeuniquefullstash transactions, cachelines of peer masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeuniquefullstash_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeuniquefullstash_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeuniquefullstash_sequence");
    super.new(name);
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITEUNIQUEFULLSTASH ,1);
      // Wait for writeuniquefullstash transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writeuniquefullstash_sequence
`endif

/** 
 * This sequence initiates WriteBack transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  WriteBack transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending WriteBack transactions, cachelines of masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeback_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeback_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeback_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITEBACK ,1);
      // Wait for writeback transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body

endclass: svt_axi_ace_master_writeback_sequence

/** 
 * This sequence initiates WriteClean transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  WriteClean transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending WriteClean transactions, cachelines of masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeclean_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeclean_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeclean_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITECLEAN ,1);
      // Wait for writeclean transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end
  endtask: body
  
endclass: svt_axi_ace_master_writeclean_sequence

/** 
 * This sequence initiates Evict transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  Evict transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending Evict transactions, cachelines of masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_evict_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_evict_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_evict_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::EVICT ,1);
      // Wait for evict transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_evict_sequence 

/** 
 * This sequence initiates WriteEvict transaction from the ACE master specified
 * with port_id , which can be a random port or a specific port configured by
 * the user through uvm_config_db.  WriteEvict transactions can be sent only
 * when the svt_axi_port_configuration::axi_interface_type of the master
 * corresponding to port_id is set to svt_axi_port_configuration::AXI_ACE.
 * Before sending WriteEvict transactions, cachelines of masters are
 * initialized to random, valid states.  Initialisation is done through front
 * door access, by sending specific transactions from the initiating master
 * (corresponding to port_id) and peer masters.  Please look up the
 * documentation of #svt_axi_cacheline_initialization for details.
 */
class svt_axi_ace_master_writeevict_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  int writeevict_enabled_ports[$];

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeevict_sequence)

  constraint valid_port_type {
    if (writeevict_enabled_ports.size())
      port_id inside {writeevict_enabled_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeevict_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  function void pre_randomize();
    super.pre_randomize();
    if(ace_ports.size() >0) begin
      foreach (ace_ports[i]) begin
        if (cfg.master_cfg[ace_ports[i]].writeevict_enable)
          writeevict_enabled_ports.push_back(ace_ports[i]);
      end
    end
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(sys_cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::WRITEEVICT ,1);
      // Wait for evict transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    svt_axi_system_configuration sys_cfg;
    is_supported = super.is_supported(cfg);
    if (is_supported) begin
      if ((cfg != null) && $cast(sys_cfg,cfg) && sys_cfg.master_cfg[port_id].writeevict_enable) begin
        is_supported = 1;
      end
      else begin
        `svt_xvm_note("body", $sformatf("The sequence cannot be run because svt_axi_port_configuration::writeevict_enable is set to 0 for port_id('d%0d)",port_id)); 
        is_supported = 0;
      end
    end
  endfunction : is_supported 

endclass: svt_axi_ace_master_writeevict_sequence 

/**
  * #- Send a sequence of writenosnoop transactions to consecutive address locations
  * #- Wait for all writenosnoop transactions to complete. <br>
  * #- Send a sequence of readnosnoop transactions to the same set of addresses
  * targetted by the writenosnoop transactions. <br>
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_writenosnoop_readnosnoop_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence writenosnoop_seq, readnosnoop_seq;

  /** Indicates if the read portion of the sequence is to be disabled */
  bit disable_reads = 0;

  /** Indicates if the write portion of the sequence is to be disabled */
  bit disable_writes = 0;

  /** Indicates if blocking mode of sending transactions should be used */
  bit use_blocking_mode = 0;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_writenosnoop_readnosnoop_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writenosnoop_readnosnoop_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(bit)::get(null, get_full_name(), "disable_reads",disable_reads);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "disable_writes",disable_writes);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "use_blocking_mode",use_blocking_mode);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".disable_reads"}, disable_reads);
    status = m_sequencer.get_config_int({get_type_name(), ".disable_writes"}, disable_writes);
    status = m_sequencer.get_config_int({get_type_name(), ".use_blocking_mode"}, use_blocking_mode);
`endif
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
    if (!disable_writes) begin
      `svt_xvm_create_on(writenosnoop_seq, p_sequencer.master_sequencer[port_id]) 
      writenosnoop_seq.writenosnoop_wt = 1;
      writenosnoop_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      void'(writenosnoop_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==local::sequence_length;
                                 });
      if (status_start_addr) begin
        writenosnoop_seq.status_start_addr = 1;
        writenosnoop_seq.start_addr = start_addr;
      end
      writenosnoop_seq.use_blocking_mode = this.use_blocking_mode;
      writenosnoop_seq.start(p_sequencer.master_sequencer[port_id]);
      writenosnoop_seq.wait_for_active_xacts_to_end();
    end
    if (!disable_reads) begin
      `svt_xvm_create_on(readnosnoop_seq, p_sequencer.master_sequencer[port_id]) 
      readnosnoop_seq.readnosnoop_wt = 1;
      if (!disable_writes) begin
        readnosnoop_seq.status_start_addr = 1;
        readnosnoop_seq.start_addr = writenosnoop_seq.start_addr;
      end
      else if (status_start_addr) begin
        readnosnoop_seq.status_start_addr = 1;
        readnosnoop_seq.start_addr = start_addr;
      end
      readnosnoop_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      void'(readnosnoop_seq.randomize with {use_directed_addr == 0;
                                      sequence_length==local::sequence_length;
                                     });
      readnosnoop_seq.use_blocking_mode = this.use_blocking_mode;
      readnosnoop_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      readnosnoop_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of shareable read transactions to consecutive address locations
  * #- Shareable read transactions can be READONCE, READCLEAN, READNOTSHAREDDIRTY, READSHARED
  * or READUNIQUE. The weights for these transactions can be passed through uvm_config_db.
  * The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. If the port is an ACE-Lite port, only READONCE transactions
  * are sent. All transactions sent are cacheline size transactions.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_read_type_shareable_region_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence read_type_seq,writeunique_writelineunique_seq;

  /** Distribution weight for generation of READONCE transactions*/
  int readonce_wt = 1;

  /** Distribution weight for generation of READCLEAN transactions*/
  int readclean_wt = 1;

  /** Distribution weight for generation of READNOTSHAREDDIRTY transactions*/
  int readnotshareddirty_wt = 1;

  /** Distribution weight for generation of READSHARED transactions*/
  int readshared_wt = 1;

  /** Distribution weight for generation of READUNIQUE transactions*/
  int readunique_wt = 1;

  /** Indicates that error was detected and sequence should not be run */
  bit is_error = 0;

  /** Indicates if memory should be initialised using WU/WLU transactions prior to sending read transactions */
  bit init_mem = 0;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_read_type_shareable_region_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports, ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_read_type_shareable_region_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readonce_wt",readonce_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readclean_wt",readclean_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readnotshareddirty_wt",readnotshareddirty_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readshared_wt",readshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readunique_wt",readunique_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "init_mem",init_mem);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".readonce_wt"}, readonce_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readclean_wt"}, readclean_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readnotshareddirty_wt"}, readnotshareddirty_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readshared_wt"}, readshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readunique_wt"}, readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".init_mem"}, init_mem);
`endif
    if (sys_cfg.master_cfg[port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
      if (readonce_wt == 0) begin
        is_error = 1;
        `svt_xvm_note("pre_body", $sformatf("The given port_id('d%0d) is an ACE_LITE interface. readonce_wt must not be 0 based on this as it is the only read transaction that can be sent from an ACE_LITE interface to a shareable region of memory", port_id));
      end
    end
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    // Check for valid port type
    begin
     if (init_mem) begin
       `svt_xvm_create_on(writeunique_writelineunique_seq, p_sequencer.master_sequencer[port_id]) 
       writeunique_writelineunique_seq.writeunique_wt = 1;
       writeunique_writelineunique_seq.writelineunique_wt = 1;
       writeunique_writelineunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
       writeunique_writelineunique_seq.force_to_cache_line_size = 1;
       if (status_start_addr) begin
         writeunique_writelineunique_seq.status_start_addr = 1;
         writeunique_writelineunique_seq.start_addr = start_addr;
       end
       void'(writeunique_writelineunique_seq.randomize with {use_directed_addr == 0;
                                     sequence_length==local::sequence_length;
                                     });
       writeunique_writelineunique_seq.start(p_sequencer.master_sequencer[port_id]);
       // Wait for transactions to finish
       writeunique_writelineunique_seq.wait_for_active_xacts_to_end();
     end

     `svt_xvm_create_on(read_type_seq, p_sequencer.master_sequencer[port_id]) 
     read_type_seq.readonce_wt = this.readonce_wt;
     read_type_seq.readclean_wt = this.readclean_wt;
     read_type_seq.readnotshareddirty_wt = this.readnotshareddirty_wt;
     read_type_seq.readshared_wt = this.readshared_wt;
     read_type_seq.readunique_wt = this.readunique_wt;
     read_type_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     if (init_mem) begin
       read_type_seq.status_start_addr = 1;
       read_type_seq.start_addr = writeunique_writelineunique_seq.start_addr;
     end
     else if (status_start_addr) begin
       // Even when init_mem is zero, sequential address mode needs to be supported
       // However, in this case, the start_addr will be the same as the one supplied
       // through config DB.
       read_type_seq.status_start_addr = 1;
       read_type_seq.start_addr = start_addr;
     end
     void'(read_type_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==local::sequence_length;
                                  });
     read_type_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      read_type_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of WRITEBACK/WRITECLEAN transactions to consecutive address locations
  * #- The weights for these transactions can be passed through uvm_config_db.
  * The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. 
  * #- A sequence of MAKEUNIQUE transactions are sent prior to sending the WRITEBACK transactions
  * so that the cachelines are in Unique Dirty State.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_writeback_writeclean_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence writeback_writeclean_seq, writenosnoop_seq, makeunique_seq;

  /** Indicates if WRITEBACK/WRITECLEAN needs to be initiated 
    * in non shareable region of memory 
    */
  bit is_nonshareable = 0;

  /** Distribution weight for generation of WRITEBACK transactions*/
  int writeback_wt = 1;

  /** Distribution weight for generation of WRITECLEAN transactions*/
  int writeclean_wt = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_writeback_writeclean_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeback_writeclean_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeback_wt",writeback_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeclean_wt",writeclean_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "is_nonshareable",is_nonshareable);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".writeback_wt"}, writeback_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".writeclean_wt"}, writeclean_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".is_nonshareable"}, is_nonshareable);
`endif
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 

    begin
    if (is_nonshareable) begin
      `svt_xvm_create_on(writenosnoop_seq, p_sequencer.master_sequencer[port_id]) 
      writenosnoop_seq.writenosnoop_wt = 1;
      writenosnoop_seq.force_to_cache_line_size = 1;
      writenosnoop_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      writenosnoop_seq.use_directed_domain_type = 1;
      writenosnoop_seq.directed_domain_type = svt_axi_transaction::NONSHAREABLE;
      if (status_start_addr) begin
        writenosnoop_seq.status_start_addr = 1;
        writenosnoop_seq.start_addr = start_addr;
      end
      void'(writenosnoop_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==local::sequence_length;
                                 });
      writenosnoop_seq.start(p_sequencer.master_sequencer[port_id]);
      writenosnoop_seq.wait_for_active_xacts_to_end();

      // Write dirty data into all the sequential addresses.
      for(int i=0;i<(writenosnoop_seq.port_cfg.num_cache_lines);i++) begin
        svt_axi_master_transaction master_xact;
        if (writenosnoop_seq.output_xact_mailbox.try_get(master_xact)) 
          writenosnoop_seq.initialize_cache_via_backdoor(master_xact.addr,1,0);
        else
          break;
      end
    end
    else begin
      `svt_xvm_create_on(makeunique_seq, p_sequencer.master_sequencer[port_id]) 
      makeunique_seq.makeunique_wt = 1;
      makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      void'(makeunique_seq.randomize with {use_directed_addr == 0;
                                     sequence_length==local::sequence_length;
                                    });
      if (status_start_addr) begin
        makeunique_seq.status_start_addr = 1;
        makeunique_seq.start_addr = start_addr;
      end
      makeunique_seq.start(p_sequencer.master_sequencer[port_id]);
      makeunique_seq.wait_for_active_xacts_to_end();
    end
     `svt_xvm_create_on(writeback_writeclean_seq, p_sequencer.master_sequencer[port_id]) 
     writeback_writeclean_seq.writeback_wt = this.writeback_wt;
     writeback_writeclean_seq.writeclean_wt = this.writeclean_wt;
     writeback_writeclean_seq.status_start_addr = 1;
     if (is_nonshareable) 
       writeback_writeclean_seq.start_addr = writenosnoop_seq.start_addr;
     else
       writeback_writeclean_seq.start_addr = makeunique_seq.start_addr;
     if (is_nonshareable) begin
       writeback_writeclean_seq.use_directed_domain_type = 1;
       writeback_writeclean_seq.directed_domain_type = svt_axi_transaction::NONSHAREABLE;
     end
     writeback_writeclean_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     void'(writeback_writeclean_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==local::sequence_length;
                               });
     writeback_writeclean_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      writeback_writeclean_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    svt_axi_system_configuration sys_cfg;
    is_supported = super.is_supported(cfg);
    if (is_supported) begin
      if (is_nonshareable && (cfg != null) && $cast(sys_cfg,cfg) && !sys_cfg.master_cfg[port_id].update_cache_for_non_coherent_xacts) begin
        `svt_xvm_note("is_supported", $sformatf("Sequence cannot be run because svt_axi_port_configuration::update_cache_for_non_coherent_xacts  must be set in the port('d%0d) from which WRITEBACK/WRITECLEAN is to be sent for a non shareable region",port_id));
        is_supported = 0;
      end
    end
  endfunction : is_supported 
endclass

/**
  * #- Send a sequence of CLEANUNIQUE transactions to consecutive address locations
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. 
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_cleanunique_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence cleanunique_seq;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_cleanunique_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cleanunique_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  task pre_body();
    super.pre_body();
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    // Check for valid port type
    begin
      `svt_xvm_create_on(cleanunique_seq, p_sequencer.master_sequencer[port_id]) 
      cleanunique_seq.cleanunique_wt = 1;
      cleanunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      if (status_start_addr) begin
        cleanunique_seq.status_start_addr = 1;
        cleanunique_seq.start_addr = start_addr;
      end
      void'(cleanunique_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                });
      cleanunique_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      cleanunique_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of WRITEUNIQUE/WRITELINEUNIQUE transactions to consecutive address locations
  * #- The weights for these transactions can be passed through uvm_config_db.
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. The port can be ACE or ACE-Lite port.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_writeunique_writelineunique_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence writeunique_writelineunique_seq;

  /** Distribution weight for generation of WRITEUNIQUE transactions*/
  int writeunique_wt = 1;

  /** Distribution weight for generation of WRITELINEUNIQUE transactions*/
  int writelineunique_wt = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_writeunique_writelineunique_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeunique_writelineunique_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeunique_wt",writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writelineunique_wt",writelineunique_wt);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".writeunique_wt"}, writeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".writelineunique_wt"}, writelineunique_wt);
`endif
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    begin
     `svt_xvm_create_on(writeunique_writelineunique_seq, p_sequencer.master_sequencer[port_id]) 
     writeunique_writelineunique_seq.writeunique_wt = this.writeunique_wt;
     writeunique_writelineunique_seq.writelineunique_wt = this.writelineunique_wt;
     writeunique_writelineunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
     writeunique_writelineunique_seq.force_to_cache_line_size = 1;
     if (status_start_addr) begin
       writeunique_writelineunique_seq.status_start_addr = 1;
       writeunique_writelineunique_seq.start_addr = start_addr;
     end
     void'(writeunique_writelineunique_seq.randomize with {use_directed_addr == 0;
                                   sequence_length==local::sequence_length;
                                   });
     writeunique_writelineunique_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      writeunique_writelineunique_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of cache maintenance transactions to consecutive address locations
  * #- Cache maintenance transactions can be MAKEINVALID, CLEANSHARED or CLEANINVALID
  * transactions.
  * #- The weights for these transactions can be passed through uvm_config_db.
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. The port can be ACE or ACE-Lite port.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_cachemaintenance_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence cachemaintenance_seq;

  /** 
    * Indicates if WRITEBACK/WRITECLEAN needs to be initiated 
    * in non shareable region of memory 
    */
  bit is_nonshareable = 0;

  /** Distribution weight for generation of CLEANSHARED transactions*/
  int cleanshared_wt = 1;

  /** Distribution weight for generation of CLEANINVALID transactions*/
  int cleaninvalid_wt = 1;

  /** Distribution weight for generation of MAKEINVALID transactions*/
  int makeinvalid_wt = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_cachemaintenance_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports,ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_cachemaintenance_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleanshared_wt",cleanshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleaninvalid_wt",cleaninvalid_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "makeinvalid_wt",makeinvalid_wt);
    status = uvm_config_db#(bit)::get(null, get_full_name(), "is_nonshareable",is_nonshareable);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".cleanshared_wt"}, cleanshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".cleaninvalid_wt"}, cleaninvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".makeinvalid_wt"}, makeinvalid_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".is_nonshareable"}, is_nonshareable);
`endif
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
    begin
      `svt_xvm_create_on(cachemaintenance_seq, p_sequencer.master_sequencer[port_id]) 
      cachemaintenance_seq.cleanshared_wt = this.cleanshared_wt;
      cachemaintenance_seq.cleaninvalid_wt = this.cleaninvalid_wt;
      cachemaintenance_seq.makeinvalid_wt = this.makeinvalid_wt;
      cachemaintenance_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      if (is_nonshareable) begin
        cachemaintenance_seq.use_directed_domain_type = 1;
        cachemaintenance_seq.directed_domain_type = svt_axi_transaction::NONSHAREABLE;
      end
      if (status_start_addr) begin
        cachemaintenance_seq.status_start_addr = 1;
        cachemaintenance_seq.start_addr = start_addr;
      end
      void'(cachemaintenance_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                     });
      cachemaintenance_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      cachemaintenance_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of MAKEUNIQUE transactions to consecutive address locations
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. The port should be an ACE port.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_makeunique_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence makeunique_seq;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_makeunique_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_makeunique_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  task pre_body();
    super.pre_body();
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    // Check for valid port type
    begin
      `svt_xvm_create_on(makeunique_seq, p_sequencer.master_sequencer[port_id]) 
      makeunique_seq.makeunique_wt = 1;
      makeunique_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      if (status_start_addr) begin
        makeunique_seq.status_start_addr = 1;
        makeunique_seq.start_addr = start_addr;
      end
      void'(makeunique_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                    });
      makeunique_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      makeunique_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/**
  * #- Send a sequence of WRITEEVICT transactions to consecutive address locations
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. The port must be an ACE port and must have 
  * svt_axi_port_configuration::writeevict_enable set.
  * #- A sequence of MAKEUNIQUE and WRITECLEAN transactions are sent prior to
  * sending the WRITEEVICT transactions so that the cachelines are in Unique
  * Clean State.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_writeevict_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  svt_axi_ace_master_writeback_writeclean_sequential_sequence writeclean_sequential_virtual_seq;

  svt_axi_ace_master_base_sequence writeevict_seq;

  int writeevict_enabled_ports[$];

  /** 
    * Indicates if WRITEEVICT needs to be initiated 
    * in non shareable region of memory 
    */
  bit is_nonshareable = 0;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_writeevict_sequential_sequence)

  constraint valid_port_type {
    if (writeevict_enabled_ports.size())
      port_id inside {writeevict_enabled_ports};
  }
  
  function new(string name = "svt_axi_ace_master_writeevict_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(bit)::get(null, get_full_name(), "is_nonshareable",is_nonshareable);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".is_nonshareable"}, is_nonshareable);
`endif
  endtask: pre_body

  function void pre_randomize();
    super.pre_randomize();
    if(ace_ports.size() >0) begin
      foreach (ace_ports[i]) begin
        if (cfg.master_cfg[ace_ports[i]].writeevict_enable)
          writeevict_enabled_ports.push_back(ace_ports[i]);
      end
    end
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(sys_cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end
    else begin
      `svt_xvm_create_on(writeclean_sequential_virtual_seq, p_sequencer) 
      void'(writeclean_sequential_virtual_seq.randomize with { sequence_length==local::sequence_length;
                                    });
      writeclean_sequential_virtual_seq.port_id = this.port_id;
      writeclean_sequential_virtual_seq.writeback_wt = 0;
      writeclean_sequential_virtual_seq.writeclean_wt = 1;
      if (status_start_addr) begin
        writeclean_sequential_virtual_seq.status_start_addr = 1;
        writeclean_sequential_virtual_seq.start_addr = start_addr;
      end
      if (is_nonshareable)
        writeclean_sequential_virtual_seq.is_nonshareable = 1;
      writeclean_sequential_virtual_seq.start(p_sequencer);

      `svt_xvm_create_on(writeevict_seq, p_sequencer.master_sequencer[port_id]) 
      writeevict_seq.writeevict_wt = 1;
      writeevict_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      void'(writeevict_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                    });
      writeevict_seq.status_start_addr = 1;
      writeevict_seq.start_addr = writeclean_sequential_virtual_seq.writeback_writeclean_seq.start_addr;
      writeevict_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      writeevict_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

  virtual function bit is_supported(svt_configuration cfg , bit silent = 0);
    svt_axi_system_configuration sys_cfg;
    is_supported = super.is_supported(cfg);
    if (is_supported) begin
      if ((cfg != null) && $cast(sys_cfg,cfg) && sys_cfg.master_cfg[port_id].writeevict_enable) begin
        if (is_nonshareable) begin
          if (!sys_cfg.master_cfg[port_id].update_cache_for_non_coherent_xacts) begin
            `svt_xvm_note("is_supported", $sformatf("Sequence cannot be run because svt_axi_port_configuration::update_cache_for_non_coherent_xacts  must be set in the port('d%0d) from which WRITEEVICT is to be sent for a non shareable region",port_id));
            is_supported = 0;

          end
        end
      end
      else begin
        `svt_xvm_note("is_supported", $sformatf("The sequence cannot be run because svt_axi_port_configuration::writeevict_enable is set to 0 for port_id('d%0d)",port_id)); 
        is_supported = 0;
      end
    end
  endfunction : is_supported 

endclass: svt_axi_ace_master_writeevict_sequential_sequence

/**
  * #- Send a sequence of EVICT transactions to consecutive address locations
  * #- The port on which the transactions are sent sent are determined by port_id which can
  * be passed via config_db. 
  * #- A sequence of MAKEUNIQUE and WRITECLEAN transactions are sent prior to
  * sending the EVICT transactions so that the cachelines are in Unique
  * Clean State.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_evict_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  svt_axi_ace_master_writeback_writeclean_sequential_sequence writeclean_sequential_virtual_seq;

  svt_axi_ace_master_base_sequence evict_seq;


  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_evict_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports};
  }
  
  function new(string name = "svt_axi_ace_master_evict_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 0;
  endfunction

  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      `svt_xvm_create_on(writeclean_sequential_virtual_seq, p_sequencer) 
      void'(writeclean_sequential_virtual_seq.randomize with { sequence_length==local::sequence_length;
                                    });
      writeclean_sequential_virtual_seq.port_id = this.port_id;
      writeclean_sequential_virtual_seq.writeback_wt = 0;
      writeclean_sequential_virtual_seq.writeclean_wt = 1;
      if (status_start_addr) begin
        writeclean_sequential_virtual_seq.status_start_addr = 1;
        writeclean_sequential_virtual_seq.start_addr = start_addr;
      end
      writeclean_sequential_virtual_seq.start(p_sequencer);

      `svt_xvm_create_on(evict_seq, p_sequencer.master_sequencer[port_id]) 
      evict_seq.evict_wt = 1;
      evict_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      void'(evict_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                               });
      evict_seq.status_start_addr = 1;
      evict_seq.start_addr = writeclean_sequential_virtual_seq.writeback_writeclean_seq.start_addr;
      evict_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      evict_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_evict_sequential_sequence

/** Basic Exclusive access sequeance
  * This Sequence provides ACE Exclusive access at system level and can be used in any AXI_ACE master port to
  * initiate Exclusive access transaction sequence using this.
  *<br>
  * Transaction Sequences Used: Exclusive Load followed by Exclusive store 
  * - Initialize cache lines if initialize_cachelines bit is set 
  * - Issue READCLEAN or READSHARED to load location and wait for the transaction to end
  * - Check the cache line state
  *   - if in Shared state issue CLEANUNIQUE 
  *   - if in Invalid state then restart Exclusive Access
  *   - else do nothing as Master can store directly to the cacheline no need to inform Interconnect
  *   .
  * - Stored data is updated to memory through WRITEBACK transaction
  * .
  *<br>
  * Please note, for generation of exclusive access transactions, svt_axi_port_configuration :: exclusive_access_enable 
  * should be set for the targeted master and svt_axi_port_configuration :: speculative_read_enable should be set to zero
  * for that master as well<br>
  * <br>
  */
class svt_axi_ace_master_exclusive_access_virtual_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

   svt_axi_ace_exclusive_access_sequence exclusive_accesses_seq;
   rand bit                              init_cachelines;
   svt_axi_transaction::burst_size_enum  exclusive_accesses_burst_size;
   rand int ace_exclusive_select = 0;
   
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 

  `svt_xvm_object_utils(svt_axi_ace_master_exclusive_access_virtual_sequence)
  
  constraint valid_port_type {
    port_id inside {ace_ports};
  } 
  
  function new(string name = "svt_axi_ace_master_exclusive_access_virtual_sequence");
    super.new(name);
  endfunction
  
  virtual task pre_body();
    int status = 0;
    super.pre_body();
  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(),"ace_exclusive_select",ace_exclusive_select);
  `elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".ace_exclusive_select"}, ace_exclusive_select);
  `endif
  endtask

  virtual task body();
    int num_masters, num_masters_q[$];
    int axi4_slave, axi4_slave_q[$];
    // Check for valid port type
     if((cfg.master_cfg[port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) &&
	(cfg.master_cfg[port_id].exclusive_access_enable != 1))begin
	`svt_xvm_warning("body", "Invalid port type specified ,valid port should be AXI_ACE type and have exclusive_access_enable set in port configuration"); 
     end 
     else begin
	super.body();
        
        foreach(cfg.master_cfg[i]) begin
          num_masters_q.push_back(i);
        end
        foreach(cfg.slave_cfg[j])
          if(cfg.slave_cfg[j].axi_interface_type == svt_axi_port_configuration::AXI4)
            axi4_slave_q.push_back(j);

        num_masters = num_masters_q.size();
        if(axi4_slave_q.size())
          axi4_slave = 1;

        // directed sequence of exclusive transactions
        directed_exclusive_sequence(0,num_masters,port_id,axi4_slave); // non-ace exclusive transacitons
        directed_exclusive_sequence(1,num_masters,port_id,axi4_slave); // ace exclusive transactions
        //directed_exclusive_sequence2();

	
        `protected
=DGbgS6b=UeDbY9]A;.>IQ7EX3Tc&;O<fCY1/)8Y2;O([X,^<4Bg6)P+R@c1>UL@
,U1=0<\#b)dVZBLKPD^.ZffN&0+TM1I,H/F^F;-fRbK(F]Eb4:I/+fWV,RX-MU/[
JO.YId^=ReRM(E;/L[Le/R@RMCYP5[AG1;fY9T+#H(:1ETIf>;/5;8b<[7_[]#\N
:(D:eE_P4MEI:GKdC&._[aU:CE&J9RR82\Z>SY#ADYX1H$
`endprotected

	  `svt_xvm_fatal("body","Casting burst_size failed");
    	  start_exclusive_accesses(0, //User Random Address 
    	    			   0, //Do Cache Line Initialization 
    				   1, //num_of_attempts to finish exclusive access successfully 
    				   4, // Burst Length
    				   exclusive_accesses_burst_size, //Burst Size
    				   svt_axi_transaction::INCR, //Burst Type
                                   axi4_slave); //To mention is there any AXI4 slave is present
         
     end // else: !if(cfg.master_cfg[port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE)
  endtask: body

  virtual task directed_exclusive_sequence(bit ace_exclusive=0, int num_masters,int ace_port_id,int axi4_slave);
  	bit rand_success;
        int port_offset, port_num, excl_seq_mode, id_width;
        svt_axi_master_transaction load[], store[], _tmp_xact;

        excl_seq_mode = 0;//$urandom_range(1,0);
        port_num = (excl_seq_mode==1) ? 1 : (ace_exclusive) ? 2 : 3;
        port_offset = (ace_exclusive) ? 3 : 0;
	// EXC LOAD
	//---------------
        load = new[num_masters];
        store = new[num_masters];
        foreach(load[ix]) begin
          if(num_masters > 4) begin
            `svt_xvm_create_on(load[ix],p_sequencer.master_sequencer[(ix%port_num)+port_offset])
            load[ix].port_cfg = cfg.master_cfg[(ix%port_num)+port_offset];
          end
          else begin
            `svt_xvm_create_on(load[ix],p_sequencer.master_sequencer[ace_port_id])
            load[ix].port_cfg = cfg.master_cfg[ace_port_id];
          end
          id_width = load[ix].port_cfg.get_id_width();
          rand_success = load[ix].randomize() with { 
                                 id == ix%id_width;
                                 if(num_masters > 4) {
                                   if(ix>0) addr == _tmp_xact.addr;	 
                                 }
		                 atomic_type == svt_axi_transaction::EXCLUSIVE;
		                 xact_type == svt_axi_transaction::COHERENT;
                                 if(ace_exclusive)
		                    coherent_xact_type == svt_axi_transaction::READSHARED;
                                 else
		                    coherent_xact_type == svt_axi_transaction::READNOSNOOP;
                                 // The possible cache_type for AXI4 slaves
                                 // are 0,1,2,3 when atomic_type is exclusive.
                                 // But when transaction is fired form AXI_ACE
                                 // master, then the possible cache_type for
                                 // AXI_ACE master and AXI4 slave is 2.
                                 if(axi4_slave)
                                   cache_type == 2;
          };
          if(!rand_success) begin
            `svt_xvm_error("directed_exclusive_seqence", " randomization failure....");
            return;
          end
          _tmp_xact = load[ix];
          if(num_masters > 4) begin
            `svt_xvm_create_on(store[ix],p_sequencer.master_sequencer[(ix%port_num)+port_offset])
            store[ix].port_cfg = sys_cfg.master_cfg[(ix%port_num)+port_offset];
          end
          else begin
            `svt_xvm_create_on(store[ix],p_sequencer.master_sequencer[ace_port_id])
            store[ix].port_cfg = sys_cfg.master_cfg[ace_port_id];
          end
          rand_success = store[ix].randomize() with { 
		                 id   == _tmp_xact.id;	 
		                 xact_type == svt_axi_transaction::COHERENT;
                                 if(ace_exclusive)
		                    coherent_xact_type == svt_axi_transaction::CLEANUNIQUE;
                                 else
		                    coherent_xact_type == svt_axi_transaction::WRITENOSNOOP;
		                 atomic_type == _tmp_xact.atomic_type; // EXCLUSIVE
		                 domain_type == _tmp_xact.domain_type; // SHAREABLE
		                 // use same control fields as the matching Exclusive read:
                                 addr == _tmp_xact.addr;
		                 burst_size  == _tmp_xact.burst_size;
		                 burst_length== _tmp_xact.burst_length;
		                 burst_type  == _tmp_xact.burst_type;
		                 prot_type   == _tmp_xact.prot_type;
		                 cache_type  == _tmp_xact.cache_type; 
          };
        end
        if(excl_seq_mode != 1) begin
          `svt_xvm_send(load[0])
          `svt_amba_debug("exc_store",$sformatf(" LOAD[0] sent... at %t",$time));
          wait(load[0].addr_status == svt_axi_transaction::ACCEPT);
          get_response(rsp);
          load[0].wait_for_transaction_end();
        end
          `svt_xvm_send(load[1])
          `svt_amba_debug("exc_store",$sformatf(" LOAD[1] sent... at %t",$time));
          wait(load[1].addr_status == svt_axi_transaction::ACCEPT);
          get_response(rsp);
          load[1].wait_for_transaction_end();
          `svt_amba_debug("exc_store",$sformatf(" LOAD[1] completed with rresp=%s... at %t",load[1].rresp[0].name(),$time));
          `svt_xvm_send(store[0])
          `svt_amba_debug("exc_store",$sformatf(" STORE[0] sent... at %t",$time));
          wait(store[0].addr_status == svt_axi_transaction::ACCEPT || store[0].is_coherent_xact_dropped);
          `svt_amba_debug("exc_store",$sformatf(" STORE[0] %s... at %t",store[0].is_coherent_xact_dropped ? "dropped" : "accepted", $time));
          get_response(rsp);
          store[0].wait_for_transaction_end();
          `svt_amba_debug("exc_store",$sformatf(" STORE[0] %s... at %t",store[0].bresp.name(), $time));
          if(num_masters > 4) begin
            `svt_xvm_send(load[2])
            `svt_amba_debug("exc_store",$sformatf(" LOAD[2] sent... at %t",$time));
            wait(load[2].addr_status == svt_axi_transaction::ACCEPT);
            get_response(rsp);
            load[2].wait_for_transaction_end();
            `svt_amba_debug("exc_store",$sformatf(" LOAD[2] completed with rresp=%s... at %t",load[2].rresp[0].name(),$time));
          end
          `svt_xvm_send(store[1])
          `svt_amba_debug("exc_store",$sformatf(" STORE[1] sent... at %t",$time));
          wait(store[1].addr_status == svt_axi_transaction::ACCEPT || store[1].is_coherent_xact_dropped == 1);
          `svt_amba_debug("exc_store",$sformatf(" STORE[1] %s... at %t",store[1].is_coherent_xact_dropped ? "dropped" : "accepted", $time));
          get_response(rsp);
          store[1].wait_for_transaction_end();
          `svt_amba_debug("exc_store",$sformatf(" STORE[1] %s... at %t",store[1].bresp.name(), $time));
          if(store[1].is_coherent_xact_dropped)
             return;
          //RD-3
        if(num_masters > 4) begin
          if(excl_seq_mode != 1) begin
            `svt_xvm_send(load[3])
            `svt_amba_debug("exc_store",$sformatf(" LOAD[3] sent... at %t",$time));
            wait(load[3].addr_status == svt_axi_transaction::ACCEPT);
            get_response(rsp);
            load[3].wait_for_transaction_end();
          end
          `svt_xvm_send(store[2])
          `svt_amba_debug("exc_store",$sformatf(" STORE[2] sent... at %t",$time));
          wait(store[2].addr_status == svt_axi_transaction::ACCEPT || store[2].is_coherent_xact_dropped == 1);
          `svt_amba_debug("exc_store",$sformatf(" STORE[2] %s... at %t",store[2].is_coherent_xact_dropped ? "dropped" : "accepted", $time));
          get_response(rsp);
          store[2].wait_for_transaction_end();
          `svt_amba_debug("exc_store",$sformatf(" STORE[2] %s... at %t",store[2].bresp.name(), $time));
          if(store[2].is_coherent_xact_dropped)
             return;
          `svt_xvm_send(load[4])
          `svt_amba_debug("exc_store",$sformatf(" LOAD[4] sent... at %t",$time));
          wait(load[4].addr_status == svt_axi_transaction::ACCEPT);
          get_response(rsp);
          load[4].wait_for_transaction_end();
          `svt_xvm_send(store[3])
          `svt_amba_debug("exc_store",$sformatf(" STORE[3] sent... at %t",$time));
          wait(store[3].addr_status == svt_axi_transaction::ACCEPT || store[3].is_coherent_xact_dropped == 1);
          `svt_amba_debug("exc_store",$sformatf(" STORE[3] %s... at %t",store[3].is_coherent_xact_dropped ? "dropped" : "accepted", $time));
          get_response(rsp);
          store[3].wait_for_transaction_end();
          `svt_amba_debug("exc_store",$sformatf(" STORE[3] %s... at %t",store[3].bresp.name(), $time));
        end

  endtask 

  virtual task start_exclusive_accesses(bit directed_addr_used ,
				bit init_cachelines, 
				int num_of_attempts,
				bit [`SVT_AXI_MAX_BURST_LENGTH_WIDTH-1:0] burst_length,
				svt_axi_transaction::burst_size_enum      burst_size,
				svt_axi_transaction::burst_type_enum      burst_type,
                                int axi4_slave);

     `svt_xvm_create_on(exclusive_accesses_seq, p_sequencer.master_sequencer[port_id]) 
     exclusive_accesses_seq.initialize_cachelines = init_cachelines; 
     void'(exclusive_accesses_seq.randomize with {
     use_directed_addr             == directed_addr_used;
     sequence_length               == local::sequence_length;
     num_of_exclusive_seq_restart  == num_of_attempts;
     exc_burst_length              == burst_length;
     exc_burst_size                == burst_size;
     exc_burst_type                == burst_type;
     if(axi4_slave)
       exclusive_axi4_slave        == 1;});
     
     //exclusive_accesses_seq is a block sequeance, no need to add explicit wait 
     exclusive_accesses_seq.start(p_sequencer.master_sequencer[port_id]);

     `svt_xvm_debug("start_exclusive_accesses", "exclusive_accesses_seq execution finished");
  endtask

  /*
  virtual task set_tr(ref svt_axi_master_transaction xact, input int port, int txn_id, bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] txn_addr=0, svt_axi_transaction::coherent_xact_type_enum typ, bit atomic, bit secure=1, bit send_xact=1);

    `svt_xvm_create_on(xact,p_sequencer.master_sequencer[port])
    if(!xact.randomize() with { xact_type == svt_axi_transaction::COHERENT;
                                coherent_xact_type == typ;
                                id == txn_id;
                                if(txn_addr > 0)
                                   addr == txn_addr;
                                prot_type[1] == !secure;
                                if(atomic)
                                   atomic_type == svt_axi_transaction::EXCLUSIVE;
                                else
                                   atomic_type == svt_axi_transaction::NORMAL;
                              })
       `svt_fatal("set_tr","couldn't randomize...");

    if(send_xact) begin
      `svt_xvm_send(xact)
      `svt_amba_debug("set_tr",$sformatf(" sent %s ",`SVT_AXI_PRINT_PREFIX1(xact)));
    end
                                
  endtask

  virtual task directed_exclusive_sequence2(bit ace_exclusive=1);
    bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr0;
    svt_axi_master_transaction load[], store[], tr[], _tmp_xact;

    load = new[5];
    store = new[5];
    //addr0 = `DEFAULT_INNER_SHARED_START_ADDR;

    set_tr(load[0],3, 8'h14, 0, svt_axi_transaction::READSHARED, 1);
    load[0].wait_for_transaction_end();
    set_tr(load[1],4, 8'h02, load[0].addr, svt_axi_transaction::READSHARED, 0);
    load[1].wait_for_transaction_end();
    set_tr(store[0],3, 8'h19, load[0].addr, svt_axi_transaction::CLEANUNIQUE, 0);
    store[0].wait_for_transaction_end();
    set_tr(load[2],4, 8'h00, load[0].addr, svt_axi_transaction::READSHARED, 0);
    load[2].wait_for_transaction_end();
    set_tr(store[1],3, 8'h00, load[0].addr, svt_axi_transaction::WRITECLEAN, 0);
    store[1].wait_for_transaction_end();
    if(store[1].final_cache_line_state != svt_axi_transaction::INVALID) begin
       set_tr(store[2],3, 8'h13, load[0].addr, svt_axi_transaction::CLEANUNIQUE, 1);
       store[2].wait_for_transaction_end();
    end
    set_tr(store[3],4, 8'h0c, load[0].addr, svt_axi_transaction::CLEANUNIQUE, 0);
    store[3].wait_for_transaction_end();

  endtask
  */

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end 
    find_ace_ports(sys_cfg);
    if(ace_ports.size() >0)
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_exclusive_access_virtual_sequence

/**
  * Creates system wide random exclusive access sequence on ACE ports.
  * Scenarios which are covered are as follows:
  */
class svt_axi_ace_random_exclusive_access_virtual_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

`ifdef SVT_UVM_TECHNOLOGY
   uvm_component my_component;
`elsif SVT_OVM_TECHNOLOGY
   ovm_component my_component;
`endif
   svt_axi_system_env my_system_env;
   typedef bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr_t;

   svt_axi_master_transaction            excl_seq;
   rand bit                              init_cachelines;
   svt_axi_transaction::burst_size_enum  exclusive_accesses_burst_size;
   
   local addr_t          addr_q[$];
   local int             id_q[$];
   local svt_axi_cache   master_caches[int];
   local svt_axi_smart_queue_2d #(addr_t) local_cache[int];

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer) 

  `svt_xvm_object_utils(svt_axi_ace_random_exclusive_access_virtual_sequence)
  
  constraint valid_port_type {
    port_id inside {ace_ports};
  } 
  
  function new(string name = "svt_axi_ace_random_exclusive_access_virtual_sequence");
    super.new(name);
  endfunction

  virtual task body();
     // Controls sending of Exclusive Store transactions.
     bit no_excl_store_post_reset = 1;
     // Randomly starts and Exclusive sequence with Exclusive Load or
     // Exclusive Store operation.
     bit use_excl_ld_to_start_seq = 1;
     // Keeps the address, id and port_id same as that of previous exclusive
     // access.
     bit use_same_excl_seq_param = 0;
     // If this bit is set then sequence should use overlapping address with
     // active transactions for Exclusive load.
     bit use_overlapped_seq_at_load  = 0;
     // If this bit is set then sequence should use overlapping address with
     // active transactions for Exclusive Store.
     bit use_overlapped_seq_at_store = 0;
     // Port ID and Transaction IDs
     int xact_port_id, xact_id;
     // Transaction address
     addr_t xact_addr;
     // When set skips Exclusive Store transactions
     bit use_skip_exclusive_store = 0;
     bit[23:0] random_scenario_mode = 12'b0000_0011_1_000;
     bit[ 7:0] random_store_mode = 8'b0000_1111;
     // Variable to specify blocking mode being used.
     int blocking_mode=1;

     addr_t  _tmp_addr;
     bit[7:0] _data[], _ctrl;
     int _indx, _port_id, _tmp[$];
     //--------------------------------------

     // Check for valid port type
     if((cfg.master_cfg[port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) &&
	(cfg.master_cfg[port_id].exclusive_access_enable != 1))begin
	`svt_xvm_warning("body", "Invalid port type specified ,valid port should be AXI_ACE type and have exclusive_access_enable set in port configuration"); 
     end 
     else begin
       super.body();
       
       `protected
g+</)_>__/IBPIESR:W]IR&:SB10V5TY)9,TUAX8IY85TG&3d=1f/)#abI1QH?\S
J=dQ(LZ/eeG315@LS0@M]:1]D(V4aT2TIU1-c/E.]Wc>H^NC;;7]&[Y0]&=1@Y+Y
7<c/aCb4SKK&]1CPggJMIXPd^.bO-V4XZM25_-7KQC:K#-+c]f_O)X<8-Nf3A2YE
VZ^>R2MO[gMfd/U;RZ>3X/?VAZK=1<X=L;WH-RPB[?1QRJ^e&)D;g?eP_,,J:[32
1B:cZ(2KVRNI&bYHKTVFX)?V5$
`endprotected

         `svt_xvm_fatal("body","Casting burst_size failed");
       
       get_cache();
       foreach(ace_ports[ix])
         local_cache[ace_ports[ix]] = new;
       
       repeat(5) begin
          //_tmp_addr = $urandom_range(cfg.master_cfg[0].outershareable_start_addr,
                                     //cfg.master_cfg[0].outershareable_end_addr );
          //_tmp_addr = $urandom_range(cfg.slave_addr_ranges[0].start_addr,
          //                           cfg.slave_addr_ranges[0].end_addr );
          _tmp_addr = 0;
          _tmp_addr[5:0] = 0;
          addr_q.push_back( _tmp_addr );
          id_q.push_back( $urandom_range(5,0));
       end
       
       // create exclusive sequence under different scenarios
       // ===================================================
       for(int i=0; i<sequence_length; i++) begin
         `svt_amba_debug("body",$sformatf("random_scenario_mode 'h%h,random_store_mode 'h%h blocking_mode 'd%d",random_scenario_mode, random_store_mode, blocking_mode));

         // start exclusive sequence
         // ------------------------
         if(!use_same_excl_seq_param) begin
            xact_addr = addr_q[$urandom_range(addr_q.size()-1,0)];
            xact_id   =   id_q[$urandom_range(id_q.size()-1,0)];
            xact_port_id = ace_ports[$urandom_range(ace_ports.size()-1,0)];
         end
         `svt_amba_debug("body",$sformatf("Starting addr 'h%h, ID 'd%0d, PORT ID 'd%0d",xact_addr, xact_id, xact_port_id));
         use_excl_ld_to_start_seq = $urandom_range(1,0);
         use_skip_exclusive_store = $urandom_range(1,0);
         if (use_excl_ld_to_start_seq)
           `svt_amba_debug("body","Using EXCLUSIVE LOAD operation to start Exclusive access sequence");
         else begin
           if (!no_excl_store_post_reset)
             `svt_amba_debug("body","Using EXCLUSIVE STORE operation to start Exclusive access sequence");
         end

         if (use_excl_ld_to_start_seq && use_skip_exclusive_store)
           `svt_amba_debug("body","Skipping EXCLUSIVE STORE in the Exclusive access sequence");
         if(no_excl_store_post_reset || use_excl_ld_to_start_seq) begin
       
            no_excl_store_post_reset = 0;
            // Randomly selects READCLEAN or READSHARED transaction for
            // Exclusive Load
            send_xact((($urandom_range(1,0)>0) ? svt_axi_transaction::READSHARED :
                                                 svt_axi_transaction::READCLEAN ),
                      xact_addr, xact_id, xact_port_id, 1,
                      use_overlapped_seq_at_load, blocking_mode, 4'h4, excl_seq );
         end
         else begin
            // Skip Exclusive Store if use_skip_exclusive_store is
            // set.However, do not skip Exclusive Store if it is being used to
            // start Exclusive access sequence.
            if (!use_skip_exclusive_store || !use_excl_ld_to_start_seq) begin
              send_xact(svt_axi_transaction::CLEANUNIQUE,
                      xact_addr, xact_id, xact_port_id, 1,
                      use_overlapped_seq_at_load, blocking_mode, 4'h4, excl_seq );
            end
         end
         // --------------------------------------------------
       
         // start non-exclusive intermediate transaction
         // ------------------------
         `svt_amba_debug("body","Sending intermediate Non-Exclusive transaction");
         send_intermediate_txn(random_scenario_mode);
         // --------------------------------------------------
       
         if(random_store_mode[0]) begin
            _tmp = ace_ports.find(x) with (x != excl_seq.port_cfg.port_id);
            _port_id = (random_store_mode[1] || _tmp.size()==0) ? excl_seq.port_cfg.port_id : _tmp[0];
            _ctrl = {4'h2, 2'b01, random_store_mode[3:2],2'b10};
            // Skip Exclusive Store if use_skip_exclusive_store is
            // set.However, do not skip Exclusive Store if it is being used to
            // start Exclusive access sequence.
            if (!use_skip_exclusive_store || !use_excl_ld_to_start_seq) begin   
              send_xact(svt_axi_transaction::CLEANUNIQUE,
                      excl_seq.addr, excl_seq.id, xact_port_id, 1,
                      use_overlapped_seq_at_store, blocking_mode, _ctrl, excl_seq );
            end        
         end
       
         // randomize scenario
         randomize_scenario_mode(random_scenario_mode, random_store_mode);
         use_same_excl_seq_param = $urandom_range(1,0);
         use_overlapped_seq_at_load = $urandom_range(1,0);
         use_overlapped_seq_at_store = $urandom_range(1,0);
         blocking_mode = $urandom_range(4,1);
         if (use_overlapped_seq_at_load || use_overlapped_seq_at_store)
           `svt_amba_debug("body","Overlapped transaction bit is set");
       end //end: for()
     end // else: !if(cfg...interface.. != ..AXI_ACE)
   endtask: body


  // -----------------------------------------------------------------------------------
  // interim_mode:
  //   [11:8] => txn_type (Load / Store / Invalidate / Write)
  //   [ 7:4] => transaction randomization control [2] = coh_xact_type [1] = addr [0]=id
  //      [3] => continue same port_id used in existing exclusive sequence
  //
  // store_mode:
  //   [5:2] => transaction randomization control [4] = coh_xact_type [3] = addr [2]=id
  //     [1] => use same port as existing exclusive sequence or other port
  //     [0] => skip exclusive store or not
  // -----------------------------------------------------------------------------------
  task randomize_scenario_mode(ref bit[23:0] interim_mode, bit[7:0] store_mode);
    randcase
       60 : interim_mode[11:8] = 0;
       20 : interim_mode[11:8] = 1;
       20 : interim_mode[11:8] = 2;
       20 : interim_mode[11:8] = 3;
    endcase
    
    randcase
       10 : interim_mode[7:4] = 4'b0111;
       20 : interim_mode[7:4] = 4'b0011;
       30 : interim_mode[7:4] = 4'b0001;
       40 : interim_mode[7:4] = 4'b0010;
    endcase
    
    randcase
       10 : interim_mode[3] = 0;
       10 : interim_mode[3] = 1;
    endcase

    // store_mode
    randcase
       10 : store_mode[3:2] = 2'b11;
       //10 : store_mode[3:2] = 2'b10;
       10 : store_mode[3:2] = 2'b01;
       //10 : store_mode[3:2] = 2'b00;
    endcase

    randcase
       20 : store_mode[1] = 0;
       80 : store_mode[1] = 1;
    endcase

    randcase
       30 : store_mode[0] = 0;
       70 : store_mode[0] = 1;
    endcase

    `svt_amba_debug("randomize", $sformatf(" interim_rand_mode='h%0x store_rand_mode='h%0x", interim_mode, store_mode));
  endtask

  task send_intermediate_txn(bit[23:0] mode);
     addr_t _addr;
     int    _id;
     int    _port_id;
     bit[7:0] _ctrl;
     int    _tmp[$];
     svt_axi_master_transaction _tr;
     svt_axi_transaction::coherent_xact_type_enum typ;

     _tmp = ace_ports.find(x) with ( x != excl_seq.port_cfg.port_id );
     _port_id = (mode[3] || _tmp.size()==0) ? excl_seq.port_cfg.port_id : _tmp[0];

     case(mode[11:10])
       0 : // LOAD
           randcase
              25 : typ = svt_axi_transaction::READONCE;
              25 : typ = svt_axi_transaction::READCLEAN;
              25 : typ = svt_axi_transaction::READSHARED;
              25 : typ = svt_axi_transaction::READNOTSHAREDDIRTY;
           endcase
       1 : // STORE
           randcase
              45 : typ = svt_axi_transaction::READUNIQUE;
              10 : typ = svt_axi_transaction::CLEANUNIQUE;
              45 : typ = svt_axi_transaction::MAKEUNIQUE;
           endcase
       2 : // CACHE MAINTENANCE
           randcase
              10 : typ = svt_axi_transaction::CLEANINVALID;
              10 : typ = svt_axi_transaction::CLEANSHARED;
              10 : typ = svt_axi_transaction::MAKEINVALID;
           endcase
       3 : // WRITE
           randcase
              10 : typ = svt_axi_transaction::WRITEUNIQUE;
              10 : typ = svt_axi_transaction::WRITELINEUNIQUE;
           endcase
       default : // CACHE MAINTENANCE
           randcase
              10 : typ = svt_axi_transaction::CLEANINVALID;
              10 : typ = svt_axi_transaction::CLEANSHARED;
              10 : typ = svt_axi_transaction::MAKEINVALID;
           endcase
     endcase

     _ctrl = {4'h1,2'b01, mode[5:4]};

     send_xact(typ, excl_seq.addr, excl_seq.id, _port_id, 0, 0, 1, _ctrl, _tr);
  endtask


  task send_xact(svt_axi_transaction::coherent_xact_type_enum typ,
                 addr_t txn_addr, int txn_id, int port_id, bit exclusive,
                 bit start_overlap_txn=0, int blocking_mode=0, bit[7:0] user_ctrl=0,
                 output svt_axi_master_transaction out_tr);

     int      _indx;
     bit[7:0] _data[];
     bit      _iu,_ic;
     longint  _age;
     bit      is_cl_valid;
     addr_t   _addr;
     svt_axi_master_transaction tr;
     /** queue to hold the transactions initiated from sequence*/
     svt_axi_transaction initiated_xacts_queue[$];
     int expected_responses = 0;
     svt_axi_transaction::coherent_xact_type_enum _typ;

     _typ = typ;

     if(user_ctrl[1] == 0 && local_cache[port_id].sq.size() <= 0) begin
        if(user_ctrl[2]==1 && typ == svt_axi_transaction::CLEANUNIQUE) begin
           if(excl_seq == null)
              _typ = svt_axi_transaction::READSHARED;
           else
              _addr = excl_seq.addr;
        end
        else
           _addr = txn_addr;
     end
     else if(user_ctrl[1] == 0)
        _addr = local_cache[port_id].get_random_entry();

     `svt_xvm_create_on(tr, p_sequencer.master_sequencer[port_id]) 
     //tr.initialize_cachelines = init_cachelines; 
     void'(tr.randomize with {
         if(cfg.master_cfg[port_id].max_num_exclusive_access > 0)
            id < cfg.master_cfg[port_id].max_num_exclusive_access ;
                          addr[5:0]    == 0;
       (user_ctrl[0]) ->  id           == txn_id;
       (user_ctrl[1]) ->  addr         == txn_addr;
       (!user_ctrl[1] && 
        coherent_xact_type == svt_axi_transaction::CLEANUNIQUE) ->  addr == _addr;
       xact_type                       == COHERENT;
       (user_ctrl[2]) ->  coherent_xact_type == _typ;
       (exclusive == 1) -> atomic_type == EXCLUSIVE;
       (exclusive == 0) -> atomic_type == NORMAL;
       (user_ctrl[1:0] == 2'h3 && exclusive) -> burst_length == excl_seq.burst_length;
       (user_ctrl[1:0] == 2'h3 && exclusive) -> burst_type   == excl_seq.burst_type  ;
       (user_ctrl[1:0] == 2'h3 && exclusive) -> burst_size   == excl_seq.burst_size  ;
                                                prot_type[1]    == 0;
       //(user_ctrl[1:0] == 2'h3 && exclusive) -> prot_type == excl_seq.prot_type;
       (user_ctrl[1:0] == 2'h3 && exclusive) -> cache_type == excl_seq.cache_type;
       //exc_burst_length              == burst_length;
       //exc_burst_size                == exclusive_accesses_burst_size;
       //exc_burst_type                == svt_axi_transaction::INCR;
     });
           `svt_xvm_debug("send_xact", {$sformatf("sending %s", tr.atomic_type.name()), `SVT_AXI_PRINT_PREFIX1(tr)} );
  
        // In case start_overlap_txn bit is set, use the same address as that
        // of any of the outstanding transactions from same port id. 
        if (start_overlap_txn) begin
          foreach (initiated_xacts_queue[i]) begin
            if (initiated_xacts_queue[i].port_id == port_id) begin
              tr.addr = initiated_xacts_queue[i].addr;
              `svt_xvm_debug("send_xact", {$sformatf("Updating address for %s since start_overlap_txn bit is set", tr.atomic_type.name()), `SVT_AXI_PRINT_PREFIX1(tr)} );
              break;
            end
          end
        end
        //tr is a block sequeance, no need to add explicit wait 
        `svt_xvm_send(tr);
        if (!tr.is_coherent_xact_dropped)
          initiated_xacts_queue.push_back(tr);
        //tr.start(p_sequencer.master_sequencer[port_id]);
        if(blocking_mode == 1 || blocking_mode == 2 || blocking_mode == 3) begin
           get_response(rsp);
           `svt_xvm_debug("send_xact", {$sformatf("sent %s", tr.atomic_type.name()), `SVT_AXI_PRINT_PREFIX1(tr)} );
        end
        else begin
           fork begin
             get_response(rsp);
            `svt_xvm_debug("send_xact", {$sformatf("sent %s", tr.atomic_type.name()), `SVT_AXI_PRINT_PREFIX1(tr)} );
           end
           join_none
        end
   
        if(blocking_mode == 1 || blocking_mode == 3) begin
           if(tr.transmitted_channel == svt_axi_transaction::READ)
              wait( tr.data_status == svt_axi_transaction::ACCEPT  ||
                    tr.data_status == svt_axi_transaction::ABORTED ||
                    tr.is_coherent_xact_dropped == 1
                  );
        end

     // delete entry from cache image which is no longer in valid state
     // so that, cache image is up-to-date with corresponding master-cache
     //
     foreach(master_caches[p_ix]) begin
       foreach(local_cache[p_ix].sq[ix]) begin
         if(master_caches[p_ix].get_index_for_addr(get_tagged_addr(local_cache[p_ix].sq[ix],p_ix)) < 0)
             local_cache[p_ix].sq.delete(ix);
       end
     end

     is_cl_valid = master_caches[port_id].read_by_addr(tr.get_tagged_addr(),_indx,_data,_iu,_ic,_age);
     if(is_cl_valid) begin
        local_cache[port_id].sq.push_back(tr.addr);
     end

     out_tr = tr;
     `svt_xvm_debug("send_xact", {$sformatf("completed %s stage-'d%0d",tr.atomic_type.name(), user_ctrl[7:4]), `SVT_AXI_PRINT_PREFIX1(tr)} );

  endtask: send_xact

  task get_cache(int indx=-1);
    svt_axi_master_agent              my_agent;
    `SVT_XVM(component)               my_component;
    svt_axi_cache                     my_cache;

    foreach (cfg.master_cfg[i]) begin
      if(indx >= 0 && i != indx) continue;

      if ( cfg.master_cfg[i].is_active &&
           (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
         ) begin
        if (p_sequencer.master_sequencer[i] != null)
          my_component = p_sequencer.master_sequencer[i].get_parent();      
        $cast(my_agent,my_component);
        if (my_agent != null)
          my_cache = my_agent.get_cache();
        master_caches[i] = my_cache;

        //if (my_cache != null) begin
          //`svt_xvm_debug("print_cache",$sformatf("Contents of master cache['d%0d]:",i));
          //my_cache.print();
        //end
      end
    end //foreach
  endtask
  
endclass


// **************************************************************************
// ************************* INTERMEDIATE LEVEL SEQUENCES *******************
// **************************************************************************

/** 
   *  This sequence attempts to create a scenario where an initiating master
   *  (given by first_port_id) receives a snoop to the same cacheline while
   *  transmitting a WRITEBACK, WRITECLEAN, WRITEEVICT or EVICT
   *  (referred to as memory update transactions).  The relative
   *  weights of WRITEBACK,WRITECLEAN,WRITEEVICT or EVICT can be
   *  set by passing writeback_wt,writeclean_wt,writeevict_wt and evict_wt
   *  respectively, through the UVM/OVM configuration infrastructure.
   *  By default, WRITEBACK and WRITECLEAN transactions have a weight of 1
   *  while the other transactions have a weight of 0.
   *  The scenario first initializes cachelines to valid states
   *  before sending memory update transactions.  Based on the kind of
   *  transaction sent, the following initial states are reached after
   *  cacheline initialization.
   *  WRITEBACK,WRITECLEAN: Unique Dirty.
   *  WRITEEVICT, EVICT: Unique Clean. 
   *  .
   *  The coherent transactions that can be sent from second_port_id are
   *  - CMO : MAKEINVALID, CLEANINVALID or CLEANSHARED
   *  STORE : MAKEUNIQUE, CLEANUNIQUE, READUNIQUE, WRITEUNIQUE or WRITELINEUNIQUE
   *  LOAD  : READONCE, READSHARED, READCLEAN or READNOTSHAREDDIRTY.
   *  In case of CLEANUNIQUE the initial state must be shared state.(if cleanunique_wt is 1)
   *  After completing initialisation for memory update, readshared will be sent from 
   *  second_port_id to initialize the states to shared, for the cleanunique addresses.
   *  .
   *  If addr_mode_select is set from test, the sequence will fire memory update 
   *  transactions from first_port_id and coherent transactions from second_port_id
   *  to the same set of sequential addresses at the same time.
   *  If addr_mode_select is low, the sequence will fire memory update 
   *  transactions from first_port_id and coherent transactions from second_port_id
   *  to the same set of random addresses at the same time.
   *  .
   *  The combination of WRITEEVICT and CLEANUNIQUE cant be exercised because
   *  Initial state of WRITEEVICT must be Unique Clean,for CLEANUNIQUE any shared state
   *  so at the same time the states cant be in unique and shared. 
   */
class svt_axi_ace_master_snoop_during_memory_update_sequence extends svt_axi_ace_master_two_port_base_virtual_sequence;

  /** Memory update sequence to be executed on first master port referenced by first_port_id */
  svt_axi_ace_master_base_sequence memory_update_seq_first_port;

  /** Coherent sequence(other than cleanunique) be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence coherent_non_cleanunique_seq_second_port;

  /** Coherent sequence(only cleanunique) be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence coherent_cleanunique_seq_second_port;
  
  /** Random coherent transaction type for second_port_id */
  rand svt_axi_transaction::coherent_xact_type_enum second_port_xact_type;

  /** Distribution weight for generation of WRITEBACK transactions used to update memory from first_port_id 
    * Applicable for both sequential and random address modes 
    */
  int writeback_wt = 1;

  /** Distribution weight for generation of WRITECLEAN transactions used to update memory from first_port_id
    * Applicable for both sequential and random address modes 
    */
  int writeclean_wt = 1;

  /** Distribution weight for generation of WRITEEVICT transactions used to update memory from first_port_id
    * Applicable for both sequential and random address modes 
    */
  int writeevict_wt = 0;

  /** Distribution weight for generation of EVICT transactions used to update memory from first_port_id
    * Applicable for both sequential and random address modes 
    */
  int evict_wt = 0;

  /** Distribution weight for generation of READUNIQUE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int readunique_wt = 0;

  /** Distribution weight for generation of CLEANUNIQUE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int cleanunique_wt = 0;

  /** Distribution weight for generation of MAKEUNIQUE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int makeunique_wt = 0;
 
  /** Distribution weight for generation of WRITEUNIQUE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int writeunique_wt = 0;

  /** Distribution weight for generation of WRITELINEUNIQUE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int writelineunique_wt = 0;

  /** Distribution weight for generation of MAKEINVALID transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int makeinvalid_wt = 0;

  /** Distribution weight for generation of CLEANINVALID transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int cleaninvalid_wt = 0;

  /** Distribution weight for generation of CLEANSHARED transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int cleanshared_wt = 0;

  /** Distribution weight for generation of CLEANSHAREDPERSIST transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int cleansharedpersist_wt = 0;

  /** Distribution weight for generation of READONCE transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int readonce_wt = 0;

  /** Distribution weight for generation of READCLEAN transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int readclean_wt = 0;

  /** Distribution weight for generation of READSHARED transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int readshared_wt = 0;

  /** Distribution weight for generation of READNOTSHAREDDIRTY transactions from second_port_id
    * Applicable only if addr_mode_select is selected as sequential 
    */
  int readnotshareddirty_wt = 0;

  /** If this bit is set to one, transactions are sent to sequential addresses
    * If low, transactions are sent to random addresses
    */
  int addr_mode_select = 0;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_snoop_during_memory_update_sequence)

  constraint solve_port_id_order {
    solve first_port_id before second_port_id;
    solve second_port_id before second_port_xact_type;
  }

  // first_port_id must be AXI_ACE since the transactions supported for first port
  // are WRITEBACK, WRITECLEAN, WRITEEVICT and EVICT
  constraint overlap_addr_valid_port_id_type {
    first_port_id inside {ace_ports}; 
    second_port_id inside {ace_ports,ace_lite_ports}; 
  } 

  constraint reasonable_coherent_xact_type { 
 
    foreach(cfg.master_cfg[i]) {
      if (i == second_port_id) {
        if (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            second_port_xact_type inside {
                                    svt_axi_transaction::READONCE,
			            svt_axi_transaction::READCLEAN,
				    svt_axi_transaction::READNOTSHAREDDIRTY,
				    svt_axi_transaction::READSHARED,
				    svt_axi_transaction::READUNIQUE,
				    svt_axi_transaction::MAKEUNIQUE,
				    svt_axi_transaction::CLEANUNIQUE,
				    svt_axi_transaction::CLEANSHARED,
				    svt_axi_transaction::CLEANSHAREDPERSIST,
                                    svt_axi_transaction::CLEANINVALID,
				    svt_axi_transaction::MAKEINVALID,
				    svt_axi_transaction::WRITEUNIQUE,
				    svt_axi_transaction::WRITELINEUNIQUE};
          }
          else {
            second_port_xact_type inside { svt_axi_transaction::READONCE,
			            svt_axi_transaction::READCLEAN,
				    svt_axi_transaction::READNOTSHAREDDIRTY,
				    svt_axi_transaction::READSHARED,
				    svt_axi_transaction::READUNIQUE,
				    svt_axi_transaction::MAKEUNIQUE,
				    svt_axi_transaction::CLEANUNIQUE,
				    svt_axi_transaction::CLEANSHARED,
                                    svt_axi_transaction::CLEANINVALID,
				    svt_axi_transaction::MAKEINVALID,
				    svt_axi_transaction::WRITEUNIQUE,
				    svt_axi_transaction::WRITELINEUNIQUE};            
          }
        } else {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            second_port_xact_type inside { svt_axi_transaction::READONCE,
				    svt_axi_transaction::CLEANINVALID,
				    svt_axi_transaction::MAKEINVALID,
				    svt_axi_transaction::CLEANSHARED,
				    svt_axi_transaction::CLEANSHAREDPERSIST,
                                    svt_axi_transaction::WRITEUNIQUE,
				    svt_axi_transaction::WRITELINEUNIQUE};
          }
          else {
            second_port_xact_type inside {svt_axi_transaction::READONCE,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::CLEANSHARED,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
        }
      } // (i==second_port_id)
    } // foreach
}

  function new(string name = "svt_axi_ace_master_snoop_during_memory_update_sequence");
    super.new(name);
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeunique_wt",writeunique_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writelineunique_wt",writelineunique_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeback_wt",writeback_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeclean_wt",writeclean_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeevict_wt",writeevict_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "evict_wt",evict_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readunique_wt",readunique_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleanunique_wt",cleanunique_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "makeunique_wt",makeunique_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "makeinvalid_wt",makeinvalid_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleaninvalid_wt",cleaninvalid_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleanshared_wt",cleanshared_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "cleansharedpersist_wt",cleansharedpersist_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readonce_wt",readonce_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readclean_wt",readclean_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readshared_wt",readshared_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readnotshareddirty_wt",readnotshareddirty_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "addr_mode_select",addr_mode_select );
  `elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".writeunique_wt"}, writeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writelineunique_wt"}, writelineunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeback_wt"}, writeback_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeclean_wt"}, writeclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeevict_wt"}, writeevict_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".evict_wt"}, evict_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readunique_wt"}, readunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".cleanunique_wt"}, cleanunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".makeunique_wt"}, makeunique_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".makeinvalid_wt"}, makeinvalid_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".cleaninvalid_wt"}, cleaninvalid_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".cleanshared_wt"}, cleanshared_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".cleansharedpersist_wt"}, cleansharedpersist_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readonce_wt"}, readonce_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readclean_wt"}, readclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readshared_wt"}, readshared_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readnotshareddirty_wt"}, readnotshareddirty_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".addr_mode_select"}, addr_mode_select );
  `endif
  endtask: pre_body
  
  virtual task body();
    int count=0;
    bit start_main_seq = 0;
    int initialization_length;
    int cleanunique_initialization;
    int is_supported_weights;

    is_supported_weights = normalize_weights_based_on_speculative_read();

    //Check for valid port types   
    if((cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) && (cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE)) begin
      `svt_xvm_warning("body", "Invalid port type specified ,second port should be ACE_LITE type if first port is ACE_LITE"); 
    end
    
    else begin
      super.body();
      //If sequential address is selected with cleanunique then the cleanunique_initialization will be made high
      //If it is high then the initialisation for cleanunique will be initiated
      if(addr_mode_select && cleanunique_wt) begin
        initialization_length = sequence_length * cleanunique_wt/(makeunique_wt + cleanunique_wt + readunique_wt + writeunique_wt + writelineunique_wt); 
        cleanunique_initialization = 1;
       end
      else begin
        initialization_length = 0;
        cleanunique_initialization = 0;
      end
      //Send random coherent transactions other than cleanunique which can generate snoop transactions with the same address 
      `svt_xvm_create_on(coherent_non_cleanunique_seq_second_port, p_sequencer.master_sequencer[second_port_id])
       coherent_non_cleanunique_seq_second_port.initialize_cachelines = 0;
       coherent_non_cleanunique_seq_second_port.direct_addr_timeout = 10000;
      //Send random coherent transactions only cleanunique which can generate snoop transactions with the same address
      `svt_xvm_create_on(coherent_cleanunique_seq_second_port, p_sequencer.master_sequencer[second_port_id])
       coherent_cleanunique_seq_second_port.initialize_cachelines = 0;
       coherent_cleanunique_seq_second_port.direct_addr_timeout = 10000;

      if(!addr_mode_select)
        coherent_non_cleanunique_seq_second_port.assign_xact_weights(second_port_xact_type);
      else begin
        coherent_non_cleanunique_seq_second_port.writeunique_wt= this.writeunique_wt;
        coherent_non_cleanunique_seq_second_port.writelineunique_wt= this.writelineunique_wt;
        coherent_non_cleanunique_seq_second_port.readunique_wt= this.readunique_wt;
        coherent_non_cleanunique_seq_second_port.makeunique_wt= this.makeunique_wt;
        coherent_non_cleanunique_seq_second_port.makeinvalid_wt= this.makeinvalid_wt;
        coherent_non_cleanunique_seq_second_port.cleaninvalid_wt= this.cleaninvalid_wt;
        coherent_non_cleanunique_seq_second_port.cleanshared_wt= this.cleanshared_wt;
        coherent_non_cleanunique_seq_second_port.cleansharedpersist_wt= this.cleansharedpersist_wt;
        coherent_non_cleanunique_seq_second_port.readonce_wt= this.readonce_wt;
        coherent_non_cleanunique_seq_second_port.readclean_wt= this.readclean_wt;
        coherent_non_cleanunique_seq_second_port.readshared_wt= this.readshared_wt;
        coherent_non_cleanunique_seq_second_port.readnotshareddirty_wt= this.readnotshareddirty_wt;
        coherent_cleanunique_seq_second_port.cleanunique_wt= this.cleanunique_wt;
      end    
      fork
      begin
       //Initiate memory update transactions from the first_port_id
       `svt_xvm_create_on(memory_update_seq_first_port, p_sequencer.master_sequencer[first_port_id])
        memory_update_seq_first_port.writeback_wt= this.writeback_wt;
        memory_update_seq_first_port.writeclean_wt= this.writeclean_wt;
        memory_update_seq_first_port.writeevict_wt= this.writeevict_wt;
        memory_update_seq_first_port.evict_wt= this.evict_wt;
        if(!addr_mode_select)
          memory_update_seq_first_port.addr_mode = svt_axi_ace_master_base_sequence::RANDOM_ADDR_MODE;
        else 
          memory_update_seq_first_port.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
        memory_update_seq_first_port.generate_only_shareable_domain = 1;
        memory_update_seq_first_port.initialize_cachelines = 1;
        memory_update_seq_first_port.suspend_xact_transmission_post_initialization = 1;
        void'(memory_update_seq_first_port.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});  
        memory_update_seq_first_port.start(p_sequencer.master_sequencer[first_port_id]);
        // Wait for Memory update transactions to finish
        memory_update_seq_first_port.wait_for_active_xacts_to_end();
      end
      begin     
        `svt_xvm_debug("body", "Waiting for cacheline initialization of memory_update_seq_first_port to be done");
        @memory_update_seq_first_port.cacheline_init_done;
        wait(start_main_seq==1);
        if(cleanunique_initialization) begin
          `svt_xvm_debug("body", "post cacheline initialization for cleanunique is done. Starting coherent_cleanunique_seq_second_port sequence...");
          void'(coherent_cleanunique_seq_second_port.randomize with {use_directed_addr == 1;sequence_length== initialization_length;});
          coherent_cleanunique_seq_second_port.start(p_sequencer.master_sequencer[second_port_id]);
          coherent_cleanunique_seq_second_port.wait_for_active_xacts_to_end();
        end
        else
          initialization_length = 0;
          
        void'(coherent_non_cleanunique_seq_second_port.randomize with {use_directed_addr == 1;sequence_length== (local::sequence_length - initialization_length);});
        coherent_non_cleanunique_seq_second_port.start(p_sequencer.master_sequencer[second_port_id]);
        // Wait for coherent transactions to finish
        coherent_non_cleanunique_seq_second_port.wait_for_active_xacts_to_end();
      end
      begin
        svt_axi_master_transaction master_xact;
        svt_axi_cache second_port_cache;
        svt_axi_ace_master_base_sequence cacheline_init_readshared_seq;
        
        if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
          if(!cleanunique_initialization)
            second_port_cache = coherent_non_cleanunique_seq_second_port.get_cache();
          else
            second_port_cache = coherent_cleanunique_seq_second_port.get_cache();
        end

        //Initialising cache lines for cleanunique transactions targetted to random addresses
        if(!cleanunique_initialization) begin
          while (count < sequence_length) begin
           memory_update_seq_first_port.output_xact_mailbox.get(master_xact); 
           coherent_non_cleanunique_seq_second_port.directed_addr_mailbox.put(master_xact.addr);

          if (
               (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
               (second_port_xact_type == svt_axi_transaction::CLEANUNIQUE) && (!addr_mode_select) 
               && !cfg.master_cfg[second_port_id].speculative_read_enable &&
               (second_port_cache != null) 
             )  begin
            `svt_xvm_debug("body", "Sending READSHARED from second_port_id post cache initialisation since second_port_xact_type is a CLEANUNIQUE transaction");
            `svt_xvm_create_on(cacheline_init_readshared_seq, p_sequencer.master_sequencer[second_port_id])
            cacheline_init_readshared_seq.readshared_wt = 1;
            cacheline_init_readshared_seq.directed_addr_mailbox.put(master_xact.addr);
            void'(cacheline_init_readshared_seq.randomize with {use_directed_addr == 1;sequence_length==1;});
            cacheline_init_readshared_seq.start(p_sequencer.master_sequencer[second_port_id]);
            cacheline_init_readshared_seq.wait_for_active_xacts_to_end();
          end              
          count++;
         end
        end
          //Initialising cache lines for cleanunique transactions targetted to sequential addresses
        else begin       
          for(int i=0; i < initialization_length; i++) begin
            memory_update_seq_first_port.output_xact_mailbox.get(master_xact); 
            coherent_cleanunique_seq_second_port.directed_addr_mailbox.put(master_xact.addr);
            if (
                 (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
                 (second_port_cache != null) &&
                 !cfg.master_cfg[second_port_id].speculative_read_enable
              ) begin
              `svt_xvm_debug("body", "Sending READSHARED from second_port_id post cache initialisation since cleanunique_wt is set");
              `svt_xvm_create_on(cacheline_init_readshared_seq, p_sequencer.master_sequencer[second_port_id])
              cacheline_init_readshared_seq.readshared_wt = 1;
              cacheline_init_readshared_seq.directed_addr_mailbox.put(master_xact.addr);
              void'(cacheline_init_readshared_seq.randomize with {use_directed_addr == 1;sequence_length==1;});
              cacheline_init_readshared_seq.start(p_sequencer.master_sequencer[second_port_id]);
              cacheline_init_readshared_seq.wait_for_active_xacts_to_end();
            end                     
          end
          for(int i=0; i < (sequence_length - initialization_length); i++) begin
            memory_update_seq_first_port.output_xact_mailbox.get(master_xact); 
            coherent_non_cleanunique_seq_second_port.directed_addr_mailbox.put(master_xact.addr);
          end  
        end
        `svt_xvm_debug("body", "Received all addresses to be initiated from both ports. Setting start_main_seq to one");
        memory_update_seq_first_port.resume_xact_transmission = 1;
        start_main_seq = 1;
      end
      join
    end
  endtask: body
  
  //Function for normalizing the weight of writeevict when cleanunique and writeevict 
  //combination occurs
  virtual function bit normalize_weights_based_on_speculative_read();
    normalize_weights_based_on_speculative_read = 1;
    if (
         cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE &&
         !cfg.master_cfg[second_port_id].speculative_read_enable &&
         cleanunique_wt) begin
      writeevict_wt = 0; 
    end
    if (
         cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE &&
         !cfg.master_cfg[second_port_id].speculative_read_enable &&
         (second_port_xact_type == svt_axi_transaction::CLEANUNIQUE) && !addr_mode_select) begin
      writeevict_wt = 0; 
    end

    
  endfunction
  
  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if(ace_ports.size() >0)
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_snoop_during_memory_update_sequence

/** 
   *  This sequence attempts to create a scenario where random coherent
   *  transactions targetting the same address are initiated from two different
   *  masters in which one is an ACE master specified with first_port_id and 
   *  another one is an ACE/ACE_LITE master specified through second_port_id.
   *  If second_port_xact_type is svt_axi_transaction::WRITENOSNOOP then the
   *  transactions will not be sent to same addresses as transactions from first_port_id, 
   *  but the transactions will be fired concurrently from the masters.
   *   
   */
class svt_axi_ace_master_overlapping_addr_sequence extends svt_axi_ace_master_two_port_base_virtual_sequence;
  

  /** Coherent sequence be executed on first master port referenced by first_port_id */
  svt_axi_ace_master_base_sequence  coherent_seq_first_port;
 
  /** Coherent sequence be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence coherent_seq_second_port;
  
  /** Random coherent transaction type for coherent_seq_first_port */
  rand svt_axi_transaction::coherent_xact_type_enum first_port_xact_type;

  /** Random coherent transaction type for coherent_seq_second_port */
  rand svt_axi_transaction::coherent_xact_type_enum second_port_xact_type;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_overlapping_addr_sequence)
  
  constraint solve_port_id_order {
    solve first_port_id before second_port_id;
    solve first_port_id before first_port_xact_type;
    solve second_port_id before second_port_xact_type;
  }
  
  // If first_port_id is ACE_LITE, second_port_id needs to be ACE_LITE too.
  constraint overlap_addr_valid_port_id_type {
    first_port_id inside {ace_ports,ace_lite_ports}; 
    if (first_port_id inside {ace_ports})
      second_port_id inside {ace_ports,ace_lite_ports}; 
    else
      second_port_id inside {ace_lite_ports}; 
  } 

  constraint reasonable_coherent_xact_type {
    
    foreach(cfg.master_cfg[i]) {
      if (i == first_port_id) {
        if (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            first_port_xact_type inside {svt_axi_transaction::READONCE,
			        svt_axi_transaction::READCLEAN,
				      svt_axi_transaction::READNOTSHAREDDIRTY,
				      svt_axi_transaction::READSHARED,
				      svt_axi_transaction::READUNIQUE,
				      svt_axi_transaction::CLEANUNIQUE,
				      svt_axi_transaction::MAKEUNIQUE,
				      svt_axi_transaction::CLEANSHARED,
              // ACE 2.0 Transaction Type
				      svt_axi_transaction::CLEANSHAREDPERSIST,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE }; 
          }
          else {
            first_port_xact_type inside {svt_axi_transaction::READONCE,
			        svt_axi_transaction::READCLEAN,
				      svt_axi_transaction::READNOTSHAREDDIRTY,
				      svt_axi_transaction::READSHARED,
				      svt_axi_transaction::READUNIQUE,
				      svt_axi_transaction::CLEANUNIQUE,
				      svt_axi_transaction::MAKEUNIQUE,
				      svt_axi_transaction::CLEANSHARED,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE };            
          }
        } else {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            first_port_xact_type inside {svt_axi_transaction::READONCE,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::CLEANSHARED,
              // ACE 2.0 Transaction Type
				      svt_axi_transaction::CLEANSHAREDPERSIST,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
          else {
            first_port_xact_type inside {svt_axi_transaction::READONCE,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::CLEANSHARED,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
        }
      } // (i==first_port_id)
    } // foreach


    foreach(cfg.master_cfg[i]) {
      if (i == second_port_id) {   
        if (cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            second_port_xact_type inside {svt_axi_transaction::READONCE,
			              svt_axi_transaction::READCLEAN,
				      svt_axi_transaction::READNOTSHAREDDIRTY,
				      svt_axi_transaction::READSHARED,
				      svt_axi_transaction::READUNIQUE,
				      svt_axi_transaction::CLEANUNIQUE,
				      svt_axi_transaction::MAKEUNIQUE,
				      svt_axi_transaction::CLEANSHARED,
              // ACE 2.0 Transaction Type
				      svt_axi_transaction::CLEANSHAREDPERSIST,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
              svt_axi_transaction::WRITEUNIQUE,
              svt_axi_transaction::WRITENOSNOOP,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
          else {
            second_port_xact_type inside {svt_axi_transaction::READONCE,
			              svt_axi_transaction::READCLEAN,
				      svt_axi_transaction::READNOTSHAREDDIRTY,
				      svt_axi_transaction::READSHARED,
				      svt_axi_transaction::READUNIQUE,
				      svt_axi_transaction::CLEANUNIQUE,
				      svt_axi_transaction::MAKEUNIQUE,
				      svt_axi_transaction::CLEANSHARED,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
                                      svt_axi_transaction::WRITEUNIQUE,
                                      svt_axi_transaction::WRITENOSNOOP,
				      svt_axi_transaction::WRITELINEUNIQUE};            
          }
        }
        else {
          if (cfg.master_cfg[i].ace_version == svt_axi_port_configuration::ACE_VERSION_2_0){
            second_port_xact_type inside {svt_axi_transaction::READONCE,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::CLEANSHARED,
              // ACE 2.0 Transaction Type
				      svt_axi_transaction::CLEANSHAREDPERSIST,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
          else {
            second_port_xact_type inside {svt_axi_transaction::READONCE,
				      svt_axi_transaction::CLEANINVALID,
				      svt_axi_transaction::MAKEINVALID,
				      svt_axi_transaction::CLEANSHARED,
				      svt_axi_transaction::WRITEUNIQUE,
				      svt_axi_transaction::WRITELINEUNIQUE};
          }
        }
      } // (i==first_port_id)
    } // foreach
  } // constraint end

  /*constraint reasonable_cleanunique_xact_type {
    // CLEANUNIQUE requires the cacheline state to be in shared state.
    // Cacheline initialisation is done based on first port. So if CLEANUNIQUE
    // needs to be sent, it must be on first_port_id, unless it needs to be sent
    // from both ports
    (first_port_xact_type != svt_axi_transaction::CLEANUNIQUE) -> 
    (second_port_xact_type != svt_axi_transaction::CLEANUNIQUE);
  }
  */
  
  function new(string name = "svt_axi_ace_master_overlapping_addr_sequence");
    super.new(name);
  endfunction

  virtual task body();
    int count=0;
    bit start_main_seq = 0;
    `svt_xvm_note("body",$sformatf("sequence_length='d%0d.first_port_id='d%0d.second_port_id='d%0d.first_port_xact_type=%s.second_port_xact_type=%s",
                  sequence_length,first_port_id,second_port_id,first_port_xact_type.name(),second_port_xact_type.name()));
    //Check for valid port types.

    if((cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
       (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)) begin
      `svt_xvm_warning("body", 
      $sformatf("Invalid ports type specified ,if first_port_id('d%0d) is ACE_LITE, second_port_id('d%0d) should be ACE_LITE as well for this sequence to run correctly.",
      first_port_id,second_port_id));
    end
    else begin
      // CLEANUNIQUE needs shared status, so cachelines should not be invalidated in second_port_id 
      // (initialisation is based on first_port_id and it invalidates random cachelines from
      // peer ports unless this bit is set)
      if (second_port_xact_type == svt_axi_transaction::CLEANUNIQUE)
        bypass_invalidation = 1;
      
      super.body();
      //Initiate random coherent transactions from first_port_id
      `svt_xvm_create_on(coherent_seq_first_port, p_sequencer.master_sequencer[first_port_id])
      coherent_seq_first_port.assign_xact_weights(first_port_xact_type);
      coherent_seq_first_port.initialize_cachelines = 1;

      //Initiate random coherent transactions with same address from second_port_id
      `svt_xvm_create_on(coherent_seq_second_port, p_sequencer.master_sequencer[second_port_id])
      coherent_seq_second_port.assign_xact_weights(second_port_xact_type);
      coherent_seq_second_port.initialize_cachelines = 0;
      coherent_seq_second_port.direct_addr_timeout = 100000;
      fork
      begin
        void'(coherent_seq_first_port.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
        coherent_seq_first_port.suspend_xact_transmission_post_initialization = 1;
        coherent_seq_first_port.start(p_sequencer.master_sequencer[first_port_id]);
        `svt_xvm_debug("body", "coherent_seq_first_port: Waiting for active transactions to end");
        coherent_seq_first_port.wait_for_active_xacts_to_end();
        `svt_xvm_debug("body", "coherent_seq_first_port: All active transactions have ended");
      end
      begin
        void'(coherent_seq_second_port.randomize with {use_directed_addr == 1;sequence_length==local::sequence_length;});
        `svt_xvm_debug("body", "coherent_seq_second_port: Waiting for coherent_seq_first_port.cacheline_init_done");
        @coherent_seq_first_port.cacheline_init_done;
        `svt_xvm_debug("body", "coherent_seq_second_port: Waiting for start_main_seq to be set");
        wait(start_main_seq==1);
        coherent_seq_second_port.start(p_sequencer.master_sequencer[second_port_id]);
        `svt_xvm_debug("body", "coherent_seq_second_port: Waiting for active transactions to end");
        coherent_seq_second_port.wait_for_active_xacts_to_end();
        `svt_xvm_debug("body", "coherent_seq_second_port: All active transactions have ended");
      end

      begin
        svt_axi_master_transaction master_xact;
        svt_axi_cache second_port_cache;
        svt_axi_cacheline_invalidation second_port_cacheline_invalidation;
        bit is_unique, is_clean, cache_status;

        if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE)
          second_port_cache = coherent_seq_second_port.get_cache();
        while (count < sequence_length) begin
          coherent_seq_first_port.output_xact_mailbox.get(master_xact); 
          coherent_seq_second_port.directed_addr_mailbox.put(master_xact.addr);
          if (
               (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
               !cfg.master_cfg[second_port_id].speculative_read_enable &&
               (
                 (second_port_xact_type == svt_axi_transaction::READONCE) || 
                 (second_port_xact_type == svt_axi_transaction::READSHARED) || 
                 (second_port_xact_type == svt_axi_transaction::READCLEAN) || 
                 (second_port_xact_type == svt_axi_transaction::READNOTSHAREDDIRTY) || 
                 (second_port_xact_type == svt_axi_transaction::READUNIQUE) 
               ) && 
               (second_port_cache != null) &&
               second_port_cache.get_status(get_tagged_addr(master_xact.addr, second_port_id),is_unique,is_clean)
             ) begin
            `svt_xvm_debug("body", "Invalidating from second_port_id post cache initialisation since second_port_xact_type is a read type transaction");
            `svt_xvm_create(second_port_cacheline_invalidation)
            second_port_cacheline_invalidation.invalidate_port = second_port_id;
            second_port_cacheline_invalidation.invalidate_addr = master_xact.addr;
            second_port_cacheline_invalidation.start(p_sequencer);
          end
          else if (
                    (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) &&
                    (
                      (second_port_xact_type == svt_axi_transaction::WRITEUNIQUE) || 
                      (second_port_xact_type == svt_axi_transaction::WRITELINEUNIQUE) 
                    ) &&
                    (second_port_cache != null) &&
                    second_port_cache.get_status(get_tagged_addr(master_xact.addr, second_port_id),is_unique,is_clean) &&
                    !is_clean
                  ) begin
           svt_axi_basic_writeclean_full_cacheline writecleanfull_seq;
            `svt_xvm_debug("body", "Sending WRITECLEAN from second_port_id post cache initialisation since second_port_xact_type is a WRITEUNIQUE/WRITELINEUNIQUE transaction");
           `svt_xvm_create_on(writecleanfull_seq, p_sequencer.master_sequencer[second_port_id])
           writecleanfull_seq.writeclean_wt = 1;
           writecleanfull_seq.directed_addr_mailbox.put(master_xact.addr);
           void'(writecleanfull_seq.randomize with {use_directed_addr == 1;sequence_length==1;});
           writecleanfull_seq.start(p_sequencer.master_sequencer[second_port_id]);
           writecleanfull_seq.wait_for_active_xacts_to_end();
          end
          count++;
        end
        `svt_xvm_debug("body", "Received all addresses to be initiated from both ports. Setting start_main_seq to one");
        coherent_seq_first_port.resume_xact_transmission = 1;
        start_main_seq = 1;
      end
      join
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size() >0) && ((ace_ports.size()+ace_lite_ports.size()) >1))
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_overlapping_addr_sequence 

/**
  * This sequence sends coherent read transactions while sending coherent write
  * transactions to the same address from another port. In most cases, the
  * interconnect will have to refetch data from the memory, if none of the
  * snoops returned data. This is because the first read may return data that
  * is not being written through the coherent write transaction depending on
  * whether the data reached the slave. Hence a second read will have to be
  * issued to ensure that the latest data is available. The sequence creates a
  * scenario where the interconnect is forced to refetch data from memory 
  */
class svt_axi_ace_master_read_during_coherent_write_sequence extends svt_axi_ace_master_two_port_base_virtual_sequence;

  /** WriteUnique/WriteLineUnique sequence to be executed on first master port referenced by first_port_id */
  svt_axi_ace_master_base_sequence memory_update_seq_first_port;

  /** Coherent sequence be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence coherent_seq_second_port;

  /** Random coherent transaction type for coherent_seq_second_port */
  rand svt_axi_transaction::coherent_xact_type_enum second_port_xact_type;

  rand svt_axi_transaction::xact_shareability_domain_enum domain_type;

  /** Distribution weight for generation of WRITEBACK transactions used to update memory */
  int writeback_wt = 1;

  /** Distribution weight for generation of WRITECLEAN transactions used to update memory*/
  int writeclean_wt = 1;

  /** Distribution weight for generation of WRITEEVICT transactions used to update memory 
    * svt_axi_port_configuration::writeevict_enable must be set in the configuration of the master
    * referred by first_port_id if this value is greater than 0
    */
  int writeevict_wt = 0;

  /** Distribution weight for generation of READONCE transactions */
  int readonce_wt = 1;

  /** Distribution weight for generation of READSHARED transactions */
  int readshared_wt = 1;

  /** Distribution weight for generation of READNOTSHAREDDIRTY transactions */
  int readnotshareddirty_wt = 1;

  /** Distribution weight for generation of READUNIQUE transactions */
  int readunique_wt = 1;

  /** Distribution weight for generation of READUNIQUE transactions */
  int readclean_wt = 1;

 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_read_during_coherent_write_sequence)

  constraint solve_port_id_order {
    solve first_port_id before second_port_id;
    solve second_port_id before second_port_xact_type;
  }

  constraint valid_port_id_type {
    first_port_id inside {ace_ports}; 
    second_port_id inside {ace_ports ,ace_lite_ports}; 
  } 

  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::INNERSHAREABLE,svt_axi_transaction::OUTERSHAREABLE};
  }

  
  function new(string name = "svt_axi_ace_master_read_during_coherent_write_sequence");
    super.new(name);
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeback_wt",writeback_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeclean_wt",writeclean_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeevict_wt",writeevict_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readonce_wt",readonce_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readshared_wt",readshared_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readnotshareddirty_wt",readnotshareddirty_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readunique_wt",readunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "readclean_wt",readclean_wt);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".writeback_wt"}, writeback_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeclean_wt"}, writeclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeevict_wt"}, writeevict_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".readonce_wt"}, readonce_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readshared_wt"}, readshared_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readnotshareddirty_wt"}, readnotshareddirty_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readunique_wt"}, readunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".readclean_wt"}, readclean_wt);
`endif
  endtask: pre_body



  virtual task body();
    
    bit coherent_seq_second_port_done = 0;
    bit memory_update_seq_done = 0;
    //Check for valid port types   
    if (cfg.master_cfg[first_port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) begin
      `svt_xvm_warning("body", "Invalid port type specified for first_port_id,valid port should be AXI_ACE"); 
    end
    else if((cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) && (cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE)) begin
      `svt_xvm_warning("body", "Invalid port type specified for second_port_id ,valid port should be AXI_ACE or ACE_LITE type"); 
    end
    
    else begin
      super.body();

      //Send random coherent transactions which can generate snoop transactions with the same address 
      `svt_xvm_create_on(coherent_seq_second_port, p_sequencer.master_sequencer[second_port_id])
      coherent_seq_second_port.readonce_wt = 1;
      if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::AXI_ACE) begin
        coherent_seq_second_port.readshared_wt = 1;
        coherent_seq_second_port.readnotshareddirty_wt= 1;
        coherent_seq_second_port.readunique_wt = 1;
        coherent_seq_second_port.readclean_wt = 1;
      end
      else begin
        coherent_seq_second_port.readshared_wt = 0;
        coherent_seq_second_port.readnotshareddirty_wt= 0;
        coherent_seq_second_port.readunique_wt = 0;
        coherent_seq_second_port.readclean_wt = 0;
      end
      coherent_seq_second_port.initialize_cachelines = 0;
      coherent_seq_second_port.direct_addr_timeout = 100000;
      for (int xact_count = 0; xact_count < sequence_length; xact_count++) begin : tag_for_loop
        fork
        begin
          //Initiate memory update transactions from the first_port_id
          `svt_xvm_create_on(memory_update_seq_first_port, p_sequencer.master_sequencer[first_port_id])
          memory_update_seq_first_port.writeback_wt= this.writeback_wt;
          memory_update_seq_first_port.writeclean_wt= this.writeclean_wt;
          memory_update_seq_first_port.writeevict_wt= this.writeevict_wt;
          memory_update_seq_first_port.use_directed_domain_type = 1;
          memory_update_seq_first_port.directed_domain_type = this.domain_type;
          memory_update_seq_first_port.initialize_cachelines = 1;
          void'(memory_update_seq_first_port.randomize with {use_directed_addr == 0;sequence_length==1;});
          memory_update_seq_first_port.start(p_sequencer.master_sequencer[first_port_id]);
          // Wait for MakeUnique transactions to finish
          memory_update_seq_first_port.wait_for_active_xacts_to_end();
          memory_update_seq_done = 1;
        end
        begin
          void'(coherent_seq_second_port.randomize with {use_directed_addr == 1;sequence_length==1;});
          `svt_xvm_debug("body", "Waiting for cacheline initialization of memory_update_seq_first_port to be done");
          @memory_update_seq_first_port.cacheline_init_done;
          `svt_xvm_debug("body", "cacheline initialization of memory_update_seq_first_port is done. Starting coherent_seq_second_port sequence...");
          coherent_seq_second_port.start(p_sequencer.master_sequencer[second_port_id]);
          coherent_seq_second_port.wait_for_active_xacts_to_end();
          coherent_seq_second_port_done = 1;
        end
        // Use first_port_id objects to provide directed addresses to other sequences.
        // Note that output_xact_mailbox will start getting filled up only after 
        // cacheline initializations of all lines are complete. 
        begin
          svt_axi_master_transaction master_xact;
          memory_update_seq_first_port.output_xact_mailbox.get(master_xact); 
          `svt_xvm_debug("body", $sformatf("%0s: Waiting for transaction status to be updated before initiating read",`SVT_AXI_PRINT_PREFIX1(master_xact)));
          // For some transactions wait on all data to be sent,
          // and on other for only address to be accepted
          fork
          begin
            fork
            begin
              wait (master_xact.is_coherent_xact_dropped == 1);
            end
            begin
              if (xact_count%2 == 0) begin
                // If all the data beats are not yet accepted, wait for atleast one beat to be accepted
                if (master_xact.data_status != svt_axi_transaction::ACCEPT)
                  wait (master_xact.data_status == svt_axi_transaction::PARTIAL_ACCEPT);
              end
              else
                wait(master_xact.addr_status == svt_axi_transaction::ACCEPT);
            end
            join_any
            disable fork;
            `svt_xvm_debug("body", $sformatf("%0s: transaction status is now updated. Initiating read",`SVT_AXI_PRINT_PREFIX1(master_xact)));
            coherent_seq_second_port.directed_addr_mailbox.put(master_xact.addr);
          end
          join
        end
        join
      end : tag_for_loop
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size() >0) && ((ace_ports.size() + ace_lite_ports.size()) > 1))
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_read_during_coherent_write_sequence

/**
  * This sequence sends cocurrent write transactions from two ports after initializing cache lines
  */
class svt_axi_ace_master_two_master_concurrent_write_sequence extends svt_axi_ace_master_two_port_base_virtual_sequence;

  /** Memory update sequence to be executed on first master port referenced by first_port_id */
  svt_axi_ace_master_base_sequence memory_update_seq_first_port;

  /** Memory update sequence to be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence memory_update_seq_second_port;

  /** Coherent sequence be executed on second master port referenced by second_port_id */
  svt_axi_ace_master_base_sequence coherent_seq_second_port;

  /** Random coherent transaction type for coherent_seq_second_port */
  rand svt_axi_transaction::coherent_xact_type_enum second_port_xact_type;

  /** Domain type of shareable transactions */
  //rand svt_axi_transaction::xact_shareability_domain_enum domain_type;

  /** Distribution weight for generation of WRITENOSNOOP transactions used to update memory */
  int writenosnoop_wt = 1;

  /** Distribution weight for generation of WRITEBACK transactions used to update memory */
  int writeback_wt = 1;

  /** Distribution weight for generation of WRITECLEAN transactions used to update memory*/
  int writeclean_wt = 1;

  /** Distribution weight for generation of WRITEEVICT transactions used to update memory 
    * svt_axi_port_configuration::writeevict_enable must be set in the configuration of the master
    * referred by first_port_id if this value is greater than 0
    */
  int writeevict_wt = 0;

  /** Distribution weight for generation of WRITEUNIQUE transactions used to update memory */
  int writeunique_wt = 1;

  /** Distribution weight for generation of WRITELINEUNIQUE transactions used to update memory */
  int writelineunique_wt = 1;


 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_two_master_concurrent_write_sequence)

  constraint solve_port_id_order {
    solve first_port_id before second_port_id;
    solve second_port_id before second_port_xact_type;
  }

  constraint valid_port_id_type {
    first_port_id inside {ace_ports}; 
    second_port_id inside {ace_ports ,ace_lite_ports}; 
  } 

  function new(string name = "svt_axi_ace_master_two_master_concurrent_write_sequence");
    super.new(name);
  endfunction

  task pre_body();
    bit status = 0;
    super.pre_body();
  `ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeback_wt",writeback_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeclean_wt",writeclean_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeevict_wt",writeevict_wt );
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writenosnoop_wt",writenosnoop_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writeunique_wt",writeunique_wt);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "writelineunique_wt",writelineunique_wt);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".writeback_wt"}, writeback_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeclean_wt"}, writeclean_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writeevict_wt"}, writeevict_wt );
    status = m_sequencer.get_config_int({get_type_name(), ".writenosnoop_wt"}, writenosnoop_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".writeunique_wt"}, writeunique_wt);
    status = m_sequencer.get_config_int({get_type_name(), ".writelineunique_wt"}, writelineunique_wt);
`endif
  endtask: pre_body



  virtual task body();
    
    bit coherent_seq_second_port_done = 0;
    bit memory_update_seq_done = 0;
    int first_port_memory_update_seq_done = 0;
    int second_port_memory_update_seq_done = 0;
    //Check for valid port types   
    if ((cfg.master_cfg[first_port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) && (cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE)) begin
      `svt_xvm_warning("body", "Invalid port type specified for first_port_id,valid port should be AXI_ACE or ACE_LITE type"); 
    end
    else if((cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::AXI_ACE) && (cfg.master_cfg[second_port_id].axi_interface_type != svt_axi_port_configuration::ACE_LITE)) begin
      `svt_xvm_warning("body", "Invalid port type specified for second_port_id ,valid port should be AXI_ACE or ACE_LITE type"); 
    end
    else begin
      super.body();

      //Send random coherent transactions which can generate snoop transactions with the same address 
      `svt_xvm_create_on(memory_update_seq_first_port, p_sequencer.master_sequencer[first_port_id])
      memory_update_seq_first_port.writeunique_wt = this.writeunique_wt;
      memory_update_seq_first_port.writelineunique_wt = this.writelineunique_wt;
      memory_update_seq_first_port.writenosnoop_wt = this.writenosnoop_wt;
      memory_update_seq_first_port.initialize_cachelines = 1;
      memory_update_seq_first_port.suspend_xact_transmission_post_initialization = 1;
      if (cfg.master_cfg[first_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
        memory_update_seq_first_port.writeback_wt = 0;
        memory_update_seq_first_port.writeclean_wt = 0;
        memory_update_seq_first_port.writeevict_wt = 0;
      end

      //Send random coherent transactions which can generate snoop transactions with the same address 
      `svt_xvm_create_on(memory_update_seq_second_port, p_sequencer.master_sequencer[second_port_id])
      memory_update_seq_second_port.writeunique_wt = this.writeunique_wt;
      memory_update_seq_second_port.writelineunique_wt = this.writelineunique_wt;
      memory_update_seq_second_port.writenosnoop_wt = this.writenosnoop_wt;
      memory_update_seq_second_port.initialize_cachelines = 1;
      memory_update_seq_second_port.suspend_xact_transmission_post_initialization = 1;
      if (cfg.master_cfg[second_port_id].axi_interface_type == svt_axi_port_configuration::ACE_LITE) begin
        memory_update_seq_second_port.writeback_wt = 0;
        memory_update_seq_second_port.writeclean_wt = 0;
        memory_update_seq_second_port.writeevict_wt = 0;
      end
      fork
      begin
        void'(memory_update_seq_first_port.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
        memory_update_seq_first_port.start(p_sequencer.master_sequencer[first_port_id]);
        // Wait for MakeUnique transactions to finish
        memory_update_seq_first_port.wait_for_active_xacts_to_end();
        first_port_memory_update_seq_done = 1;
      end
      begin
        void'(memory_update_seq_second_port.randomize with {use_directed_addr == 0;sequence_length==local::sequence_length;});
        memory_update_seq_second_port.start(p_sequencer.master_sequencer[second_port_id]);
        // Wait for MakeUnique transactions to finish
        memory_update_seq_second_port.wait_for_active_xacts_to_end();
        second_port_memory_update_seq_done = 1;
      end
      join_none

      // When cacheline initialization of both ports are done, resume xact transmission.
      // This is so that write transactions will start together on all ports 
      fork
      begin
        @memory_update_seq_first_port.cacheline_init_done;
      end
      begin
        @memory_update_seq_second_port.cacheline_init_done;
      end
      join
      memory_update_seq_first_port.resume_xact_transmission = 1;
      memory_update_seq_second_port.resume_xact_transmission = 1;
      `svt_xvm_debug("body", "Waiting for memory_update_seq_first_port sequence to be done");
      wait(first_port_memory_update_seq_done == 1);
      `svt_xvm_debug("body", "memory_update_seq_first_port is done... waiting for memory_update_seq_second_port sequence to be done");
      wait(second_port_memory_update_seq_done == 1);
      `svt_xvm_debug("body", "coherent_seq_second_port is done... ");
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size() >0) && ((ace_ports.size() + ace_lite_ports.size()) > 1))
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_two_master_concurrent_write_sequence

// =====================================================================================================
// ---------------------------- BARRIER Sequences ---------------------------------------------------------
/**
  * This sequence does the following:
  * Sends a number of pre barrier store transactions based on num_pre_barrier_stores
  * Sends a barrier pair
  * Sends a post barrier flag transaction. Any master that can observe this flag should be
  * able to observe the transactions before the barrier
  * From another port in the same domain, the location written through the flag transaction is 
  * continously read (load). When the value set through the flag transaction is read back, the loop 
  * terminates. The flag transaction is a post-barrier transaction, so if its value is observable, 
  * It then reads back all the locations written through the pre barrier store transactions and 
  * checks that all the data that was written is read back correctly. Thus, this sequence is
  * self-checking. Note that this step is not done if pre_barrier_xact_type is PRE_BARRIER_CACHE_MAINTENANCE 
  * since the data is not available in cache maintenance transactions. Instead, the sequence checks 
  * that when a post-barrier transaction completes all pre-barrier cache maintenance transactions
  * should have completed.
  * The ports on which the pre barrier stores and the loads are sent are randomly chosen
  * based on configuration. The type of store transaction is based on the setting in 
  * pre_barrier_xact_type. Loads can be READSHARED,READONCE,READCLEAN or
  * READNOTSHAREDDIRTY. 
  * Some interesting scenarios that can be exercised using this sequence are.
  * Each of these scenarios is repeated for sequence_length:
  * 1. num_pre_barrier_stores=1,num_observers=1 : A single pre-barrier store
  * followed by a post barrier flag with one observer reading the post barrier
  * flag and later reading the location addressed by pre_barrier store. 
  * 2. num_pre_barrier_stores=1,num_observers>1 : A single pre-barrier store
  * followed by a post barrier flag with many observers reading the post barrier
  * flag and later reading the location addressed by pre_barrier store. 
  * 3. num_pre_barrier_stores>1,num_observers=1 : Many pre-barrier stores
  * followed by a post barrier flag with one observer reading the post barrier
  * flag and later reading the locations addressed by pre_barrier store. 
  * 4. num_pre_barrier_stores>1,num_observers>1 : Many pre-barrier stores
  * followed by a post barrier flag with many observers reading the post barrier
  * flag and later reading the locations addressed by pre_barrier store. 
  *
  * NOTE: Continuous polling may need adding interval between two consecutive transactions. See
  *       poll_barrier_flag_and_check_post_barrier_contents task for details.
  *       This task is part of class svt_axi_ace_master_barrier_base_virtual_sequence
  *       from which current class is derived.
  */
class svt_axi_ace_master_shareable_store_barrier_load_sequence extends svt_axi_ace_master_barrier_base_virtual_sequence;

  typedef enum int {
    PRE_BARRIER_COHERENT_STORE = 0, // MAKEUNIQUE,READUNIQUE,WRITUNIQUE,WRITELINEUNIQUE
    PRE_BARRIER_WRITEBACK_MEMORY_UPDATE = 1, // WRITEBACK
    PRE_BARRIER_WRITECLEAN_MEMORY_UPDATE = 2, //WRITECLEAN
    PRE_BARRIER_CACHE_MAINTENANCE = 3 // CACHE MAINTENANCE (MAKEINVALID, CLEANINVALID, CLEANSHARED)
  } pre_barrier_xact_type_enum;

  /** Represents the master port from which the sequence will be initiated. */ 
  rand int unsigned first_port_id;

  rand int unsigned second_port_id;

  bit status;
  
  /** 
    * Weight for sending MAKEUNIQUE, READUNIQUE, WRITEUNIQUE or WRITELINEUNIQUE  
    * as pre barrier stores
    */
  int pre_barrier_coherent_store_wt = 50;

  /** 
    * Weight for sending MAKEUNIQUE followed by WRITEBACK to same address
    * as pre barrier stores
    */
  int pre_barrier_writeback_memory_update_wt = 15;

  /** 
    * Weight for sending MAKEUNIQUE followed by WRITECLEAN to same address
    * as pre barrier stores
    */
  int pre_barrier_writeclean_memory_update_wt = 15;

  /** 
    * Weight for sending MAKEINVALID, CLEANINVALID and CLEANSHARED 
    * as pre barrier stores
    */
  int pre_barrier_cache_maintenance_wt = 30;

  /** The kind of pre-barrier transactions */
  rand pre_barrier_xact_type_enum pre_barrier_xact_type;

  /** Number of pre-barrier stores to be issued before issuing a barrier and post-barrier transaction */
  rand int num_pre_barrier_stores = 1;

  /** 
    * Number of ports that are observing the pre barrier stores. The location written 
    * through the flag transaction is read from this many ports that fall in the
    * same domain
    */ 
  rand int num_observers = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_shareable_store_barrier_load_sequence)
  
  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::INNERSHAREABLE,
                        svt_axi_transaction::OUTERSHAREABLE};
  }

  constraint reasoanble_pre_barrier_xact_type {
    pre_barrier_xact_type dist {
      PRE_BARRIER_COHERENT_STORE := pre_barrier_coherent_store_wt,
      PRE_BARRIER_WRITEBACK_MEMORY_UPDATE := pre_barrier_writeback_memory_update_wt,
      PRE_BARRIER_WRITECLEAN_MEMORY_UPDATE := pre_barrier_writeclean_memory_update_wt,
      PRE_BARRIER_CACHE_MAINTENANCE := pre_barrier_cache_maintenance_wt 
    };
  }

  /** Greater weightage for sending only one pre barrier xact because
    * there is a greater possibility of things going wrong there */
  constraint reasonable_num_pre_barrier_xacts {
    num_pre_barrier_stores dist {
      1 := 50,[2:10] := 50
    }; 
  }

  constraint reasonable_num_observers {
    num_observers inside {[1:(ace_ports.size()+ace_lite_ports.size()-1)]};
  } 
  
  function new(string name = "svt_axi_ace_master_shareable_store_barrier_load_sequence");
    super.new(name);
  endfunction

  virtual task pre_body();
    super.pre_body();
    raise_phase_objection();

`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "first_port_id", first_port_id);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".first_port_id"}, first_port_id);
`endif
    `svt_xvm_debug("body", $sformatf("first_port_id is 'd%0d as a result of %0s.", first_port_id, status ? "config DB" : "randomization"));
  endtask

  /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

  virtual task body();
    int num_barrier_seq = 0;
    int count; 
    int rand_domain_ports[$],observer_ports[$];
    bit is_only_ace = 0;
    super.body();

    `svt_xvm_debug("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"});
    // WRITEBACK, WRITECLEAN can be sent only from full ACE ports
    if ((pre_barrier_xact_type == PRE_BARRIER_WRITEBACK_MEMORY_UPDATE) || 
        (pre_barrier_xact_type == PRE_BARRIER_WRITECLEAN_MEMORY_UPDATE)) 
      is_only_ace = 1;
    if (!get_random_ports_in_domain(domain_type,(num_observers+1),0,is_only_ace,rand_domain_ports) && !rand_domain_ports.size()) begin
      `svt_xvm_debug("body", 
      $sformatf("There are no two ports for domain_type(%0s). This sequence needs atleast two active ports for the given domain type",domain_type.name()));
    end
    else begin
      int temp_sequence_length;
      // First port is the port from which store is sent. All others are observers.
      foreach (rand_domain_ports[i]) begin
        if ((i == 0) && (status == 0))
          first_port_id = rand_domain_ports[i];
        else begin
          if(status == 0)
          observer_ports.push_back(rand_domain_ports[i]);
          else begin
            if( first_port_id != rand_domain_ports[i])
             observer_ports.push_back(rand_domain_ports[i]);
           end
         end
       end
      temp_sequence_length = sequence_length;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. num_pre_barrier_stores = 'd%0d",sequence_length,num_pre_barrier_stores));
      
      count = 0;
      while (temp_sequence_length > 0) begin
        int _length;
        svt_axi_master_transaction pre_barrier_write_xacts[$], post_barrier_xact;
        svt_axi_ace_barrier_pair_sequence barrier_pair_seq;
        /** Coherent sequence (pre barrier) be executed on first master port referenced by first_port_id */
        svt_axi_ace_master_base_sequence  pre_barrier_coherent_seq;
        count++;
        if (num_pre_barrier_stores < temp_sequence_length)
          _length = num_pre_barrier_stores;
        else
          _length = temp_sequence_length;
        temp_sequence_length -= _length;
        `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. temp_sequence_length = 'd%0d",sequence_length,temp_sequence_length));
        //Initiate random coherent transactions from first_port_id
        // Sends barrier sequence, but does not wait until all transactions are complete
        `svt_xvm_debug("body",$sformatf("Sending barrier sequence 'd%0d",count));
        if (pre_barrier_xact_type == PRE_BARRIER_COHERENT_STORE) begin
          // Create a sequence to send pre-barrier stores. 
          pre_barrier_coherent_seq=create_pre_barrier_store_seq(_length,first_port_id,1,1,1,1);
        end
        else if ((pre_barrier_xact_type == PRE_BARRIER_WRITEBACK_MEMORY_UPDATE) ||
                 (pre_barrier_xact_type == PRE_BARRIER_WRITECLEAN_MEMORY_UPDATE) 
                 ) begin
          svt_axi_ace_master_base_sequence makeunique_seq;
          svt_axi_basic_writeback_full_cacheline writeback_seq;
          svt_axi_basic_writeclean_full_cacheline writeclean_seq;
          // First make some dirty cache lines so that WRITEBACK will go out
          `svt_xvm_create_on(makeunique_seq, p_sequencer.master_sequencer[first_port_id])    
          makeunique_seq.disable_all_weights();
          makeunique_seq.makeunique_wt = 1;
          void'(makeunique_seq.randomize with {use_directed_addr == 0;sequence_length==_length;});
          makeunique_seq.use_directed_domain_type = 1;
          makeunique_seq.directed_domain_type = domain_type;
          makeunique_seq.start(p_sequencer.master_sequencer[first_port_id]); 
          makeunique_seq.wait_for_active_xacts_to_end();
          if (pre_barrier_xact_type == PRE_BARRIER_WRITEBACK_MEMORY_UPDATE) begin
            `svt_xvm_create_on(writeback_seq, p_sequencer.master_sequencer[first_port_id])    
            pre_barrier_coherent_seq = writeback_seq;
          end
          else if (pre_barrier_xact_type == PRE_BARRIER_WRITECLEAN_MEMORY_UPDATE) begin
            `svt_xvm_create_on(writeclean_seq, p_sequencer.master_sequencer[first_port_id])    
            pre_barrier_coherent_seq = writeclean_seq;
          end
          void'(pre_barrier_coherent_seq.randomize with {use_directed_addr == 1;sequence_length==_length;});
          pre_barrier_coherent_seq.direct_addr_timeout = 1000000;
          pre_barrier_coherent_seq.use_directed_domain_type = 1;
          pre_barrier_coherent_seq.directed_domain_type = domain_type;
          while (makeunique_seq.output_xact_mailbox.num()) begin
            svt_axi_master_transaction _master_xact;
            makeunique_seq.output_xact_mailbox.get(_master_xact);
            pre_barrier_coherent_seq.directed_addr_mailbox.put(_master_xact.addr);
          end
        end
        else if (pre_barrier_xact_type == PRE_BARRIER_CACHE_MAINTENANCE)  begin
          svt_axi_ace_master_base_sequence cachemaintenance_seq;
          `svt_xvm_create_on(cachemaintenance_seq, p_sequencer.master_sequencer[first_port_id])    
          cachemaintenance_seq.makeinvalid_wt = 1;
          cachemaintenance_seq.cleaninvalid_wt = 1;
          cachemaintenance_seq.cleanshared_wt = 1;
          cachemaintenance_seq.initialize_cachelines = 1;
          void'(cachemaintenance_seq.randomize with {use_directed_addr == 0;sequence_length==_length;});
          cachemaintenance_seq.use_directed_domain_type = 1;
          cachemaintenance_seq.directed_domain_type = domain_type;
          pre_barrier_coherent_seq = cachemaintenance_seq;
        end
       
        // Send the pre_barrier stores and send a barrier pair after it. 
        send_barrier_sequence(first_port_id,pre_barrier_coherent_seq,pre_barrier_write_xacts,barrier_pair_seq);
        // Send a post barrier 'flag transaction'. This transaction should complete only after response to 
        // barrier is received. The code below then polls for the flag set from another port. 
        send_post_barrier_xact(first_port_id,barrier_pair_seq.write_barrier_xact,barrier_pair_seq.read_barrier_xact,1,post_barrier_xact);
        if (pre_barrier_xact_type != PRE_BARRIER_CACHE_MAINTENANCE) begin
          // Number of loads expected
          num_barrier_seq = num_barrier_seq + observer_ports.size();
          `svt_xvm_debug("body",$sformatf("barrier sequence 'd%0d is sent.num_barrier_seq = 'd%0d",count,num_barrier_seq));
          for (int observer_count = 0; observer_count < observer_ports.size(); observer_count++) begin 
            automatic svt_axi_ace_master_base_sequence post_barrier_read_seq;
            automatic int j = count;
            automatic int _observer_count = observer_count; 
            fork
            begin
              // Create a sequence which will read from all the locations that were written to in the store
              post_barrier_read_seq = create_post_barrier_load_seq(pre_barrier_write_xacts.size(),observer_ports[_observer_count],1,1,1,1);
              // Poll the location written in the 'flag transaction' above and check for the value written
              // in the flag transaction. When the same value as 'flag transaction' is received we know that
              // the post-barrier transaction is complete and therefore all the pre-barrier transactions should
              // be observable. Check that here
              poll_barrier_flag_and_check_post_barrier_contents(observer_ports[_observer_count],post_barrier_read_seq,pre_barrier_write_xacts,post_barrier_xact);
              // As each load is complete, decrement this count
              num_barrier_seq--;
              `svt_xvm_debug("body",$sformatf("Polling and checking on port 'd%0d for barrier sequence 'd%0d is complete. num_barrier_seq = 'd%0d.num_observer_ports = 'd%0d",observer_ports[_observer_count],j,num_barrier_seq,observer_ports.size()));
            end
            join_none
`protected
,MX@^RRf#\_K85,;)E\5JDP49E-KQadBS[FKbC\?,.,\HXfWIN\T4)#TK3>GX?Z/
L+ePMYJ/O.TM8dfI^_WOe[NB-8c7<c;GPcG1E>FcNTN[e5LeUO6OJce3FUBWP<W[R$
`endprotected
            
          end
          `svt_xvm_debug("body","Waiting for all barrier sequences and memory checking to complete");
          wait (num_barrier_seq == 0);
          `svt_xvm_debug("body","All barrier sequences and memory checking are complete");
        end
        // For cache maintenance transactions just check that when the post barrier transaction completes
        // all the pre barrier cache maintenance transactions are complete
        else begin
          `svt_xvm_debug("body",$sformatf("Waiting for post_barrier_xact %0s to end",`SVT_AXI_PRINT_PREFIX1(post_barrier_xact))); 
          wait (`SVT_AXI_XACT_STATUS_ENDED(post_barrier_xact));
          `svt_xvm_debug("body",$sformatf("post_barrier_xact %0s is now ended.Checking if pre barriers are all ended...",`SVT_AXI_PRINT_PREFIX1(post_barrier_xact))); 
          // Check if all cache maintenance transactions are done 
          foreach (pre_barrier_write_xacts[i]) begin
            svt_axi_master_transaction _master_xact;
            _master_xact = pre_barrier_write_xacts[i];
            if (!`SVT_AXI_XACT_STATUS_ENDED(_master_xact)) begin
              `svt_xvm_debug("body",$sformatf("Expected pre barrier transaction %0s to end before post barrier %0s end, but it is not yet ended",`SVT_AXI_PRINT_PREFIX1(_master_xact),`SVT_AXI_PRINT_PREFIX1(post_barrier_xact))); 
            end
          end
        end
      end // for(sequence length)
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size()+ace_lite_ports.size() >1))
      return 1;
    return 0;  
  endfunction : is_applicable

endclass: svt_axi_ace_master_shareable_store_barrier_load_sequence 

/**
  * This sequence does the following:
  * Sends a number of pre barrier write transactions based on num_pre_barrier_stores
  * Sends a barrier pair
  * Sends post barrier read transaction to the same address.
  * Since the reads are post barrier transactions, all the previous writes should be
  * observable to the reads 
  * All write transactions sends are WRITENOSNOOP transaction and read transactions
  * are READNOSNOOP transactions
  */
class svt_axi_ace_master_nonshareable_store_barrier_load_sequence extends svt_axi_ace_master_barrier_base_virtual_sequence;
  
  /** Number of pre-barrier stores to be issued before issuing a barrier and post-barrier transaction */
  rand int num_pre_barrier_stores = 1;

  /** 
    * Number of ports from which the sequence must be executed 
    */ 
  rand int num_ports = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_nonshareable_store_barrier_load_sequence)
  
  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::NONSHAREABLE};
  }

  /** Greater weightage for sending only one pre barrier xact because
    * there is a greater possibility of things going wrong there */
  constraint reasonable_num_pre_barrier_xacts {
    num_pre_barrier_stores dist {
      1 := 50,[2:10] := 50
    }; 
  }

  constraint reasonable_num_ports {
    num_ports inside {[1:(ace_ports.size()+ace_lite_ports.size()-1)]};
  } 
  
  function new(string name = "svt_axi_ace_master_nonshareable_store_barrier_load_sequence");
    super.new(name);
  endfunction

  virtual task send_write_barrier_read_seq(int port_id);
    svt_axi_ace_master_base_sequence  pre_barrier_nonshareable_seq;
    int temp_sequence_length = sequence_length;
    int count = 0;
    int readnosnoop_count = 0;
    `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. num_pre_barrier_stores = 'd%0d",sequence_length,num_pre_barrier_stores));
    
    while (temp_sequence_length > 0) begin
      svt_axi_master_transaction read_xact_queue[$];
      int _length;
      svt_axi_master_transaction pre_barrier_write_xacts[$], post_barrier_xact;
      svt_axi_ace_barrier_pair_sequence barrier_pair_seq;
      /** Coherent sequence (pre barrier) be executed on first master port referenced by port_id */
      count++;
      if (num_pre_barrier_stores < temp_sequence_length)
        _length = num_pre_barrier_stores;
      else
        _length = temp_sequence_length;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. temp_sequence_length = 'd%0d. num of pre barrier stores = 'd%0d. port_num = 'd%0d",sequence_length,temp_sequence_length, num_pre_barrier_stores, port_id));
      //Initiate random coherent transactions from port_id
      // Sends barrier sequence, but does not wait until all transactions are complete
      `svt_xvm_debug("body",$sformatf("Sending barrier sequence 'd%0d. port_num = 'd%0d",count,port_id));
      // Create a sequence to send pre-barrier stores. 
      `svt_xvm_create_on(pre_barrier_nonshareable_seq, p_sequencer.master_sequencer[port_id])
      pre_barrier_nonshareable_seq.disable_all_weights();
      pre_barrier_nonshareable_seq.writenosnoop_wt = 1;
      pre_barrier_nonshareable_seq.use_directed_domain_type = 1;
      pre_barrier_nonshareable_seq.directed_domain_type = this.domain_type;
      // Send pre-barrier transactions
      void'(pre_barrier_nonshareable_seq.randomize with {use_directed_addr == 0;sequence_length==_length;});
      // Send the pre_barrier stores and send a barrier pair after it. 
      send_barrier_sequence(port_id,pre_barrier_nonshareable_seq,pre_barrier_write_xacts,barrier_pair_seq);
      readnosnoop_count = 0;
      if (pre_barrier_write_xacts.size() != _length)
        `svt_error("body",$sformatf("expected 'd%0d pre barrier write transactions, but found only 'd%0d", 
                   _length,pre_barrier_write_xacts.size()));
      while (readnosnoop_count < _length) begin
        svt_axi_master_transaction readnosnoop_xact,_master_xact;
        svt_axi_ace_barrier_readnosnoop_sequence barrier_readnosnoop_seq;
        bit my_associate_barrier, rand_success;
        _master_xact = pre_barrier_write_xacts[readnosnoop_count];
        // Set associate barrier for the first one. The VIP Master does not reorder transactions
        // So if the first readnosnoop can be observed (by setting it as post barrier) all transactions
        // following it should be observable.
        if (readnosnoop_count == 0) 
          my_associate_barrier = 1;
        else
          my_associate_barrier = 0;
        `svt_xvm_debug("body",$sformatf("Sending readnosnoop for pre barrier write transaction %0s",`SVT_AXI_PRINT_PREFIX1(_master_xact)));
        `svt_xvm_create_on(barrier_readnosnoop_seq,p_sequencer.master_sequencer[port_id]);
        barrier_readnosnoop_seq.my_associate_barrier = my_associate_barrier;
        barrier_readnosnoop_seq.write_xact = _master_xact;
        barrier_readnosnoop_seq.use_directed_domain_type = 1;
        barrier_readnosnoop_seq.directed_domain_type = this.domain_type;
        if (my_associate_barrier) begin
          barrier_readnosnoop_seq.assoc_write_barrier_xact = barrier_pair_seq.write_barrier_xact;
          barrier_readnosnoop_seq.assoc_read_barrier_xact = barrier_pair_seq.read_barrier_xact;
        end
        barrier_readnosnoop_seq.start(p_sequencer.master_sequencer[port_id]);
        read_xact_queue.push_back(barrier_readnosnoop_seq.output_read_xact);
        readnosnoop_count++;
      end
      foreach (read_xact_queue[i]) begin
        `svt_xvm_debug("body",$sformatf("Waiting for transaction %0s to end",`SVT_AXI_PRINT_PREFIX1(read_xact_queue[i])));
        wait (`SVT_AXI_XACT_STATUS_ENDED(read_xact_queue[i]));
        `svt_xvm_debug("body",$sformatf("transaction %0s is ended",`SVT_AXI_PRINT_PREFIX1(read_xact_queue[i])));
      end
      check_pre_barrier_and_post_barrier_xact_contents(pre_barrier_write_xacts,read_xact_queue);
      temp_sequence_length -= _length;
    end
  endtask

  virtual task body();
    int num_barrier_seq = 0;
    int first_port_id, second_port_id,count; 
    int rand_domain_ports[$],observer_ports[$];
    super.body();
    `svt_xvm_debug("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"})
    if (!get_random_ports_in_domain(domain_type,num_ports,0,0,rand_domain_ports) && !rand_domain_ports.size()) begin
      `svt_xvm_debug("body", 
      $sformatf("There are no ports for domain_type(%0s). This sequence needs atleast one active port for the given domain type",domain_type.name()));
    end
    else begin
      int num_barrier_seq = 0;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. num_pre_barrier_stores = 'd%0d",sequence_length,num_pre_barrier_stores));
      // First port is the port from which store is sent. All others are observers.
      foreach (rand_domain_ports[i]) begin
        automatic int port_num = rand_domain_ports[i];
        fork
        begin
          send_write_barrier_read_seq(port_num);
          num_barrier_seq++;
        end
        join_none
      end
      // Wait until sequences on all ports are complete
      wait (num_barrier_seq == rand_domain_ports.size());
      `svt_xvm_debug("body","All barrier sequences and memory checking are complete");
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size()+ace_lite_ports.size() >1))
      return 1;
    return 0;  
  endfunction : is_applicable
endclass: svt_axi_ace_master_nonshareable_store_barrier_load_sequence 

/**
  * This sequence does the following:
  * Send a number of transactions to load . The number of transactions sent
  * is based on num_pre_barrier_loads. 
  * Send a barrier pair
  * Send a post barrier transaction that is associated to the barrier pair. This transaction
  * will be send out only after the response to the barrier pair is received
  * When the post barrier transaction ends, check that all pre barrier transactions have also
  * ended. 
  */
class svt_axi_ace_master_load_barrier_sequence extends svt_axi_ace_master_barrier_base_virtual_sequence;
  
  /** Number of pre-barrier stores to be issued before issuing a barrier and post-barrier transaction */
  rand int num_pre_barrier_loads = 1;

  /** 
    * Number of ports from which the sequence needs to be executed 
    */ 
  rand int num_ports = 1;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_load_barrier_sequence)
  
  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::INNERSHAREABLE,
                        svt_axi_transaction::OUTERSHAREABLE,
                        svt_axi_transaction::NONSHAREABLE};
  }

  /** Greater weightage for sending only one pre barrier xact because
    * there is a greater possibility of things going wrong there */
  constraint reasonable_num_pre_barrier_xacts {
    num_pre_barrier_loads dist {
      1 := 50,[2:10] := 50
    }; 
  }

  constraint reasonable_num_observers {
    num_ports inside {[1:(ace_ports.size()+ace_lite_ports.size()-1)]};
  } 
  
  function new(string name = "svt_axi_ace_master_load_barrier_sequence");
    super.new(name);
  endfunction

  virtual task do_load_followed_by_barrier(int port_num);
    int count = 0;
    int temp_sequence_length = sequence_length;
    `svt_xvm_debug("body", $sformatf("Sending pre barrier loads on port 'd%0d", port_num));
    while (temp_sequence_length > 0) begin
      int _length;
      svt_axi_master_transaction pre_barrier_load_xacts[$], post_barrier_xact;
      svt_axi_ace_barrier_pair_sequence barrier_pair_seq;
      /** Coherent sequence (pre barrier) be executed on first master port referenced by port_num */
      svt_axi_ace_master_base_sequence  pre_barrier_coherent_seq;
      count++;
      if (num_pre_barrier_loads < temp_sequence_length)
        _length = num_pre_barrier_loads;
      else
        _length = temp_sequence_length;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. num of pre barrier loads = 'd%0d. port_num = 'd%0d",sequence_length,_length,port_num));
      //Initiate random coherent transactions from port_num 
      // Sends barrier sequence, but does not wait until all transactions are complete
      `svt_xvm_debug("body",$sformatf("Sending barrier sequence 'd%0d. port_num = 'd%0d",count,port_num));
      temp_sequence_length -= _length;
      // Create a sequence to send pre-barrier loads. 
      pre_barrier_coherent_seq=create_pre_barrier_load_seq(_length,port_num,1,1,1,1);
      // Send the pre_barrier loads and send a barrier pair after it. 
      send_barrier_sequence(port_num,pre_barrier_coherent_seq,pre_barrier_load_xacts,barrier_pair_seq);
      // Send a post barrier that associates to the barrier pair sent earlier
      send_post_barrier_xact(port_num,barrier_pair_seq.write_barrier_xact,barrier_pair_seq.read_barrier_xact,0,post_barrier_xact);
      `svt_xvm_debug("body",$sformatf("Waiting for post barrier %0s to end",`SVT_AXI_PRINT_PREFIX1(post_barrier_xact)));
      wait (`SVT_AXI_XACT_STATUS_ENDED(post_barrier_xact));
      `svt_xvm_debug("body",$sformatf("post barrier %0s ended",`SVT_AXI_PRINT_PREFIX1(post_barrier_xact)));
      // Check that all pre barrier loads have ended by the time a response
      // to post barriers is received. According to spec. a barrier ensures
      // that if a port can observe post barrier transactions after the barrier, then 
      // It can observe transactions before the barrier.
      if(post_barrier_xact.barrier_type == svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER) begin
        foreach (pre_barrier_load_xacts[i]) begin
          svt_axi_master_transaction _master_xact;
          _master_xact = pre_barrier_load_xacts[i];
          if(_master_xact.barrier_type == svt_axi_transaction::NORMAL_ACCESS_RESPECT_BARRIER) begin 
            if (!`SVT_AXI_XACT_STATUS_ENDED(_master_xact)) begin
              `svt_xvm_debug("body",$sformatf("Expected pre barrier transaction %0s to end before post barrier %0s end, but it is not yet ended",`SVT_AXI_PRINT_PREFIX1(_master_xact),`SVT_AXI_PRINT_PREFIX1(post_barrier_xact))); 
            end
          end
        end
      end
    end
  endtask

  virtual task body();
    int num_barrier_seq = 0;
    int first_port_id, second_port_id,count; 
    int rand_domain_ports[$],observer_ports[$];
    super.body();
    `svt_xvm_debug("body", {"Executing ", (is_item() ? "item " : "sequence "), get_name(), " (", get_type_name(), ")"})
    if (!get_random_ports_in_domain(domain_type,num_ports,0,0,rand_domain_ports) && !rand_domain_ports.size()) begin
      `svt_xvm_debug("body", 
      $sformatf("There are no ports for domain_type(%0s). This sequence needs atleast one active port for the given domain type",domain_type.name()));
    end
    else begin
      int num_barrier_seq;
      num_barrier_seq = 0;
      `svt_xvm_debug("body", $sformatf("sequence_length = 'd%0d. num_pre_barrier_loads = 'd%0d",sequence_length,num_pre_barrier_loads));
      foreach (rand_domain_ports[i]) begin
        automatic int port_num = rand_domain_ports[i];
        fork
        begin
          do_load_followed_by_barrier(port_num);
          num_barrier_seq++;
        end
        join_none
      end
      // Wait until sequences on all ports are complete
      wait (num_barrier_seq == rand_domain_ports.size());
    end
  endtask: body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);
    if((ace_ports.size()+ace_lite_ports.size() >1))
      return 1;
    return 0;  
  endfunction : is_applicable

endclass: svt_axi_ace_master_load_barrier_sequence 
// ---------------------------- END OF BARRIER Sequences ---------------------------------------------------------

// =====================================================================================================
// ---------------------------- DVM Sequences ---------------------------------------------------------
/**
  * This sequence sends DVM operations followed by a DVM sync from one port or multiple
  * ports of a given domain. Prior to sending DVM operations and DVM sync a few normal transactions
  * as specified in num_pre_dvm_xacts is sent. The above sequence is repeated for sequence_length.
  * The sequence also triggers another sequence that sends DVM Complete transactions from ports that receive DVM Syncs. 
  * The sequence terminates only when DVM completes for each of the DVM syncs sent out
  * from a port are received from the interconnect
  * This sequence is not added to the library (except for documentation) because it kills any
  * snoop response sequences supplied by the testbench to run a dvm specific snoop response. Adding
  * it to the library and running it may cause undesirable results and therefore this sequence must 
  * be run in a separate test
  */
class svt_axi_ace_master_dvm_virtual_sequence extends svt_axi_ace_master_base_virtual_sequence;

  /** Represents the length of the sequence. */
  int unsigned sequence_length = 10;

  typedef enum bit {
    ALL_DVM_MASTERS = 0, // Send DVM from all masters in domain
    ONE_MASTER = 1   // Send DVM from only one master
  } multi_port_type_enum;

  /** Indicates if DVM transactions need to be sent from only one port in a 
    * given domain or from all ports in a domain
    * Currently supports only ONE_MASTER
    */
  rand multi_port_type_enum multi_port_type;

  rand int num_pre_dvm_xacts = 1;

  /**
    * The shareability domain of the DVM transactions to be sent
    */
  rand svt_axi_transaction::xact_shareability_domain_enum domain_type;
  
  /** Represents the weights of second part dvm message type distribution */
  int unsigned second_part_dvm_message_type_wt_min = 10;
  int unsigned second_part_dvm_message_type_wt_mid = 40;
  int unsigned second_part_dvm_message_type_wt_max = 50;
  
  /** Place holder for a sequence to be sent before DVM transactions are initiated */
  svt_axi_ace_master_base_sequence  pre_dvm_seq;

  /** Handles of infinite snoop response sequeunces running on each master */
`ifdef __SVDOC__
  `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER 128
`else
`ifndef SVT_AXI_MAX_NUM_MASTERS_0
  `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER `SVT_AXI_MAX_NUM_MASTERS
`else
  `define _SVT_AXI_DVM_SEQ_MAX_NUM_MASTER 1
`endif
`endif
  svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER];

  /** 
    * Handles of infinite DVM complete sequences running on each master. 
    * These wait for a DVM Sync snoop transaction and send DVM complete transactions
    */
  svt_axi_ace_master_dvm_complete_sequence dvm_complete_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER];

`ifdef SVT_UVM_TECHNOLOGY
    uvm_component my_component;
`elsif SVT_OVM_TECHNOLOGY
    ovm_component my_component;
`endif
    svt_axi_system_env my_system_env;
    svt_axi_system_configuration sys_cfg;

  constraint valid_domain_type {
    domain_type inside {svt_axi_transaction::INNERSHAREABLE,
                        svt_axi_transaction::OUTERSHAREABLE};
  }

  constraint reasonable_num_pre_dvm_xacts {
    num_pre_dvm_xacts > 0;
    num_pre_dvm_xacts < 10;
  }

  `svt_xvm_object_utils(svt_axi_ace_master_dvm_virtual_sequence)

  /** Class Constructor */
  function new (string name = "svt_axi_ace_master_dvm_virtual_sequence");
    super.new(name);
  endfunction : new
  
  virtual task pre_body();
    bit status;
    svt_configuration base_cfg;
    super.pre_body();
    raise_phase_objection();

`ifdef SVT_UVM_TECHNOLOGY
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "sequence_length", sequence_length);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_min", second_part_dvm_message_type_wt_min);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_mid", second_part_dvm_message_type_wt_mid);
    status = uvm_config_db#(int unsigned)::get(null, get_full_name(), "second_part_dvm_message_type_wt_max", second_part_dvm_message_type_wt_max);
`elsif SVT_OVM_TECHNOLOGY
    status = m_sequencer.get_config_int({get_type_name(), ".sequence_length"}, sequence_length);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_min"}, second_part_dvm_message_type_wt_min);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_mid"}, second_part_dvm_message_type_wt_mid);
    status = m_sequencer.get_config_int({get_type_name(), ".second_part_dvm_message_type_wt_max"}, second_part_dvm_message_type_wt_max);
`endif

    p_sequencer.get_cfg(base_cfg);
    if (!$cast(sys_cfg, base_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_system_configuration class");
    end
    my_component = p_sequencer.get_parent();
    if (!$cast(my_system_env,my_component)) begin
      `svt_xvm_fatal("body", "Expected parent of svt_axi_system_sequencer to be of type svt_axi_system_env, but it is not");
    end

  endtask

 /** Drop objection */
  virtual task post_body();
    drop_phase_objection();
  endtask: post_body

  virtual task send_dvm_sequence(int port_id, int num_of_syncs);
    fork
    begin
      for (int sync_num = 0; sync_num < num_of_syncs; sync_num++) begin
        svt_axi_ace_master_base_sequence  pre_dvm_seq;
        svt_axi_ace_master_dvm_base_sequence dvm_operation_seq = new("dvm_operation_seq");
        svt_axi_ace_master_dvm_base_sequence dvm_sync_seq = new("dvm_sync_seq");
        // First send some normal transactions
        `svt_xvm_create_on(pre_dvm_seq, p_sequencer.master_sequencer[port_id])
        pre_dvm_seq.writenosnoop_wt = 1;
        pre_dvm_seq.readnosnoop_wt = 1;
        void'(pre_dvm_seq.randomize with {use_directed_addr == 0;sequence_length==num_pre_dvm_xacts;});
        `svt_xvm_debug("body",$psprintf("Sending pre dvm transactions on master 'd%0d",port_id));
        pre_dvm_seq.start(p_sequencer.master_sequencer[port_id]);
        `svt_xvm_debug("body",$sformatf("Starting DVM TLB Invalidate Operation on master 'd%0d",port_id));
        // First send a TLB Invalidate DVM operation
        `svt_xvm_do_on_with(dvm_operation_seq, p_sequencer.master_sequencer[port_id], 
                                 {seq_xact_type==svt_axi_transaction::DVMMESSAGE;
           			dvm_message_type == 3'b000;}
            	   )
        `svt_xvm_debug("body",$sformatf("Starting DVM Branch Predictor Invalidate Operation on master 'd%0d",port_id));
        // Branch Predictor Invalidate
        `svt_xvm_do_on_with(dvm_operation_seq, p_sequencer.master_sequencer[port_id], 
                                 {seq_xact_type==svt_axi_transaction::DVMMESSAGE;
           			dvm_message_type == 3'b001;}
            	   )
        `svt_xvm_debug("body",$sformatf("Starting DVM Sync on master 'd%0d",port_id));
        // Send a DVM sync to know when the DVM operation is complete
        // in all peer masters.
        `svt_xvm_do_on_with(dvm_sync_seq, p_sequencer.master_sequencer[port_id], 
                                 {seq_xact_type==svt_axi_transaction::DVMMESSAGE;
           			 dvm_message_type == 3'b100;}
            	     )
        `svt_xvm_debug("body",$psprintf("Waiting for all pre dvm transactions on master 'd%0d to end",port_id));
        pre_dvm_seq.wait_for_active_xacts_to_end();
        `svt_xvm_debug("body",$psprintf("All pre dvm transactions on master 'd%0d have ended",port_id));
      end
    end
    // Thread that waits for all the DVM complete transactions to be received
    begin
      // Wait for all the corresponding DVM Completes to be received
      for (int count_dvm_complete = 0; count_dvm_complete < num_of_syncs; count_dvm_complete++) begin
        wait_for_dvm_complete(snoop_resp_seq, port_id);
      end
    end
    join
  endtask

  virtual task wait_for_dvm_complete( svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[], int port_id );
    `SVT_DATA_BASE_OBJECT_TYPE ev_xact;
    svt_axi_snoop_transaction snoop_xact;

    `svt_xvm_debug("wait_for_dvm_complete",$psprintf("Waiting for DVM COMPLETE on master 'd%0d",port_id));
    `protected
89XA;=G)CH>LL)>A4@C\9d<gTbQTdJJLV6Ta?U+RXZ8HL\:FY_ZZ2)25a(JP;[Fb
1W#L[2@8@P9[&1E,IaFb@eV+QXE5.c80\>13MZ?KQP]>(>CdZH#HNQ@2e,]D/<d6
\cKX]A4Z:X#]F+6MG(fSUT+bfMgZCKYg:R5=;8BgD(7fQQd)M(&UNJ@2M$
`endprotected

    if (!$cast(snoop_xact,ev_xact)) begin
      `svt_xvm_fatal("wait_for_dvm_complete","Transaction obtained through EVENT_DVM_COMPLETE_XACT is not of type svt_axi_snoop_transaction");
    end
    else begin
      `svt_xvm_debug("wait_for_dvm_complete",$psprintf("Received DVM COMPLETE %0s on master 'd%0d. Waiting for it to complete...",`SVT_AXI_ACE_PRINT_PREFIX(snoop_xact),port_id));
      wait (
             (snoop_xact.snoop_resp_status == svt_axi_snoop_transaction::ACCEPT) ||
             (snoop_xact.snoop_resp_status == svt_axi_snoop_transaction::ABORTED) 
           );
      `svt_xvm_debug("wait_for_dvm_complete",$psprintf("Received DVM COMPLETE %0s on master 'd%0d is now complete.",`SVT_AXI_ACE_PRINT_PREFIX(snoop_xact),port_id));
    end
  endtask

  virtual task start_snoop_response_seq_for_dvm(int port_id, svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[`_SVT_AXI_DVM_SEQ_MAX_NUM_MASTER] );
    void'(snoop_resp_seq[port_id].randomize());
    `svt_xvm_debug("start_snoop_response_seq_for_dvm", $sformatf("Stopping existing snoop sequences on snoop sequencer 'd%0d to start dvm specific sequence of type svt_axi_ace_master_snoop_response_sequence('d%0d) as this virtual sequence requires a snoop sequence of this type",port_id, snoop_resp_seq[port_id]));
    my_system_env.master[port_id].snoop_sequencer.stop_sequences();
    fork begin
      snoop_resp_seq[port_id].start(my_system_env.master[port_id].snoop_sequencer);
    end
    join_none

    if (sys_cfg.master_cfg[port_id].auto_gen_dvm_complete_enable == 0) begin
      dvm_complete_seq[port_id] = new($sformatf("dvm_complete_seq['d%0d]",port_id));
      `svt_xvm_create_on(dvm_complete_seq[port_id], p_sequencer.master_sequencer[port_id])
      dvm_complete_seq[port_id].snoop_resp_seq = snoop_resp_seq[port_id];
      `ifdef SVT_UVM_TECHNOLOGY
      `ifdef SVT_UVM_12_OR_HIGHER 
      dvm_complete_seq[port_id].parent_starting_phase = get_starting_phase();
      `else
      dvm_complete_seq[port_id].parent_starting_phase = starting_phase;
      `endif
      `endif
      void'(dvm_complete_seq[port_id].randomize()); 
      dvm_complete_seq[port_id].start(p_sequencer.master_sequencer[port_id]);
    end
  endtask

  virtual task body();
    bit status;
    int local_sequence_length;
    int dvm_seq_status[];

    int num_ports;

    int rand_domain_ports[$];
    `svt_xvm_debug("body", "Entered...");
    foreach (my_system_env.master[i]) begin
      if (
           (sys_cfg.master_cfg[i].is_active == 1) &&
           (
             (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) ||
             (
               (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
               sys_cfg.master_cfg[i].dvm_enable
             )
           )
         ) begin
        `svt_xvm_create_on(snoop_resp_seq[i], my_system_env.master[i].snoop_sequencer)
        start_snoop_response_seq_for_dvm(i, snoop_resp_seq);
      end
    end

    // ALL_DVM_MASTERS not supported yet
    /*if (multi_port_type == ALL_DVM_MASTERS)
      num_ports = 0; // All ports
    else 
      num_ports = 1;
*/

    // Enable sending from multiple ports (set second argument to 0)if all ports have auto_gen_dvm_complete_enable.
    // If atleast one port requires that DVM complete seq is run, then enable sending from
    // only 1 port (second argument is set to 1), because this sequence cannot currently handle that.
    if (!get_random_ports_in_domain(domain_type,1,multi_port_type,0,rand_domain_ports) && !rand_domain_ports.size()) begin
      `svt_xvm_error("body", 
      $sformatf("There are no ports for domain_type(%0s).Not executing sequence...",domain_type.name()));
    end
    else begin
      dvm_seq_status = new[rand_domain_ports.size()];
      foreach (dvm_seq_status[i])
        dvm_seq_status[i] = 0;
      foreach (rand_domain_ports[i]) begin
        automatic int my_port_id = rand_domain_ports[i];
        automatic int loop_count = i;
        fork
        begin
          send_dvm_sequence(my_port_id,sequence_length);
          `svt_xvm_debug("body",$psprintf("All DVM COMPLETE transactions on master 'd%0d are now complete. Setting dvm_seq_status['d%0d] to 1",my_port_id,loop_count));
          dvm_seq_status[loop_count] = 1;
        end
        join_none
      end
      `svt_xvm_debug("body",$sformatf("Waiting for all DVM Completes to be received"));
      foreach (dvm_seq_status[x]) 
        wait (dvm_seq_status[x] == 1);
    end
    `svt_xvm_debug("body",$sformatf("All DVM Completes are received. Exiting body..."));
  endtask : body

  virtual function bit is_applicable(svt_configuration cfg);
    svt_axi_system_configuration sys_cfg;
    if(!$cast(sys_cfg, cfg)) begin
      `svt_xvm_fatal("is_applicable", "Unable to cast cfg to svt_axi_system_configuration type");
    end
    find_ace_ports(sys_cfg);

    // Atleast one port should have DVM enabled.
    foreach (ace_ports[i]) begin
      int _port_id = ace_ports[i];
      if (sys_cfg.master_cfg[_port_id].dvm_enable && sys_cfg.master_cfg[_port_id].is_active)
        return 1;
    end
    foreach (ace_lite_ports[i]) begin
      int _port_id = ace_lite_ports[i];
      if (sys_cfg.master_cfg[_port_id].dvm_enable && sys_cfg.master_cfg[_port_id].is_active)
        return 1;
    end
  endfunction : is_applicable
endclass

/** Sends Multi-Part DVM Transaction from randomly selected ports. While sending multipart dvm
  * transactions it also sends dvm transactions from same port along with coherent shareable and
  * non-shareable transactions from same and other ports. Multipart and singlepart DVM transactions
  * are sent simulataneously from one or more randomly selected ports in parallel.
  * Scenarios Covered::
  *   - independent write channel transaction progress along with dvm transactions
  *   - independency of ID usage between write channel transactions and DVM transactions
  *   - independent read channel transaction progress along with dvm transactions
  *   - ID usage restrictions between read channel non-dvm transactions and DVM transactions
  *   - multi-part DVM transactions
  *   - multi-part DVM transactions with second part having DVM Sync and other opcodes
  *   - multi-part DVM Sync transactions with second part having DVM Sync and other opcodes
  *   - time overlapped multi-part dvm and non-multi-part dvm transactions
  *   - time overlapped coherent write, coherent read and multi-part dvm and non-multi-part dvm transactions
  *   .
  */
class svt_axi_ace_master_multipart_dvm_virtual_sequence extends svt_axi_ace_master_dvm_virtual_sequence;
  svt_axi_system_configuration sys_cfg;

  protected semaphore read_channel_sema = new(1);
  protected svt_axi_master_transaction active_write_q[$], active_read_q[$], active_dvm_q[$];
  local int last_dvm_msg_type = 0;
  local bit stop_sending_transactions[$];
  local semaphore send_transaction_sema = new(1);

  `svt_xvm_object_utils(svt_axi_ace_master_multipart_dvm_virtual_sequence)

  /** Class Constructor */
  function new (string name = "svt_axi_ace_master_multipart_dvm_virtual_sequence");
    super.new(name);
  endfunction : new

`protected
AZ]TV>+f8VHZYb\]8LOC@DL-,BP6Z98@^F8aE.+?#(^f@g>E<[[H+)4K.8X14S3U
H[#CHe>-;/O2H:5I;8G[I=d?R:@VFEE96<_]/a](Z.9dCZDXBVP@+(4KJ$
`endprotected

  virtual task send_dvm_sequence(int port_id, int num_of_syncs);
    int      curr_rd_q_size;
    bit[2:0] dvm_message_type;
    bit      _send_multipart_dvm;
    svt_axi_master_transaction tr, tr1, tr2;
    svt_axi_master_transaction _temp_rd_xact_id_q[$];
    bit[`SVT_AXI_MAX_ID_WIDTH-1:0]  _multi_dvm_first_txn_id, id_q[$];
    string   _id_str = "", _id_str2="";

    while(1) begin
      // find if all the unique id(s) used by read channel 
      if(my_system_env.master[port_id].driver.get_ids_used_by_active_master_transactions(id_q,"non_dvm",0)) begin

        // acquire read channel lock so that, other process can't send xact on read channel
        read_channel_sema.get();
        _id_str = " outstanding read ID: ";
        foreach(id_q[ix]) begin
          _id_str = $sformatf("%s 'h%0x",_id_str,id_q[ix]);
        end
  
        randcase
          40 : _send_multipart_dvm = 0;
          60 : _send_multipart_dvm = 1;
        endcase

        if(last_dvm_msg_type != 4 && active_read_q.size() > 0 && _send_multipart_dvm == 0)
           randcase
             20 : dvm_message_type = 6;
             40 : dvm_message_type = $urandom_range(3,0);
             40 : dvm_message_type = 4;
           endcase
        else
           randcase
             20 : dvm_message_type = 6;
             80 : dvm_message_type = $urandom_range(3,0);
           endcase
  
        `svt_xvm_create_on(tr1, p_sequencer.master_sequencer[port_id])
         tr1.port_cfg = sys_cfg.master_cfg[port_id];
//vcs-vip-protect
`protected
ZXB&f[U=e3P[V6A]CMBQR;ecYbP5OR&@5591N>c<9&EYJ;0ZP1TR4)/DHHT]+2gZ
#8NE>H;B5B__1I\#10\N>P3b=,_Z=MYX]#;(X[T+?dYcU_]1:&cFL(@dWY>-R=Z/
(c2^&54^]F1.OM_U)P9eNd3b7$
`endprotected

         void'(tr1.randomize() with {
            if(id_q.size() > 0) { id inside {id_q}; }

            tr1.addr[0] == _send_multipart_dvm;
            tr1.addr[14:12] == dvm_message_type;
        /*    if(tr1.addr[14:12] == 0){
               tr1.addr[11:0] inside {12'hA00,12'hA20,12'hb00,12'hB40,12'hB60,12'hF00,12'h600,12'hB44}; }
            if(tr1.addr[14:12] == 2){
               tr1.addr[11:0] inside {'h200,'h300};}
            if(tr1.addr[14:12] == 3){
               tr1.addr[11:0] inside {12'h300,12'hB40,12'h000};}*/

            tr1.data_before_addr == 0;
            tr1.xact_type == svt_axi_transaction::COHERENT;
            tr1.coherent_xact_type == svt_axi_transaction::DVMMESSAGE;
         });
        _multi_dvm_first_txn_id = tr1.id;
        active_dvm_q.push_back(tr1);
        remove_q_on_xact_end("dvm",tr1);
        `svt_xvm_send(tr1)
        `svt_axi_xxm_debug("send_dvm_sequence",$psprintf("Sent %0s DVM transaction %0s on port 'd%0d. dvm_message_type = 'h%0x and waiting for it to complete (%s) (dvm_id: 'h%0x) [%s]", ((_send_multipart_dvm) ? "first-part of MULTI-PART" : "single"), `SVT_AXI_PRINT_PREFIX1(tr1),port_id,dvm_message_type, _id_str, tr1.id, _id_str2));
        fork
          get_response(rsp);
        join_none
    
        if(_send_multipart_dvm) begin
           tr1.wait_for_transaction_end(); // get_response doesn't work well in some simulator
           // second-part of multipart dvm sequence
           `svt_xvm_create_on(tr2, p_sequencer.master_sequencer[port_id])
            tr2.port_cfg = sys_cfg.master_cfg[port_id];
            tr2.set_multipart_dvm_flag();
            void'(tr2.randomize() with {
               tr2.id == _multi_dvm_first_txn_id;
               tr2.addr[0] == 0;
               tr2.addr[14:12] dist {4:=second_part_dvm_message_type_wt_max, [0:3]:/second_part_dvm_message_type_wt_mid, 6:=second_part_dvm_message_type_wt_min};
       //<DP> DVM checks are failing without these constraints , Need to check if the checker is written properly as second part of dvm does not have any constraints on the address bit<DP>
               /*if(tr2.addr[14:12] == 0){
                 tr2.addr[11:0] inside {12'hA00,12'hA20,12'hb00,12'hB40,12'hB60,12'hF00,12'h600,12'hB44}; }
               if(tr2.addr[14:12] == 2){
                 tr2.addr[11:0] inside {'h200,'h300};}
               if(tr2.addr[14:12] == 3){
                 tr2.addr[11:0] inside {12'h300,12'hB40,12'h000};}*/
               tr2.data_before_addr == 0;
               tr2.xact_type == svt_axi_transaction::COHERENT;
               tr2.coherent_xact_type == svt_axi_transaction::DVMMESSAGE;
            });
           `svt_xvm_send(tr2)
           `svt_axi_xxm_debug("send_dvm_sequence",$psprintf("Sending second-part of MULTI-PART DVM transaction %0s on port 'd%0d. dvm_message_type = 'h%0x",`SVT_AXI_PRINT_PREFIX1(tr2),port_id,dvm_message_type));
           active_dvm_q.push_back(tr2);
           remove_q_on_xact_end("dvm",tr2);
           get_response(rsp);
        end
        // realease read channel lock so that, other process can send xact on read channel
        read_channel_sema.put(); 
  
        if(dvm_message_type == 4) begin
           fork
             wait_for_dvm_complete( snoop_resp_seq, port_id );
           join_none
           tr1.wait_for_transaction_end();
           if(_send_multipart_dvm)
              tr2.wait_for_transaction_end();
        end
        if(_send_multipart_dvm) 
        `svt_axi_xxm_debug("send_dvm_sequence",$psprintf("Sent complete MULTI-PART DVM transaction %0s on port 'd%0d. dvm_message_type = 'h%0x and %s on port 'd%0d",`SVT_AXI_PRINT_PREFIX1(tr1),port_id, dvm_message_type, `SVT_AXI_PRINT_PREFIX1(tr2),port_id));
        last_dvm_msg_type = dvm_message_type;

        // dvm transaction is sent so break the while() loop
        break;
      end // non_dvm ID list
      else begin
        curr_rd_q_size = active_read_q.size();
        if(curr_rd_q_size > 0) begin
           `svt_amba_debug("send_dvm_sequence",$sformatf("no ID available for DVM transaction to send so, waiting for at least one active non-dvm transaction to complete from read channel before checking for ID availability again..."));
           wait(active_read_q.size() < curr_rd_q_size);
           `svt_amba_debug("send_dvm_sequence",$sformatf("active non-dvm transaction completion from read channel detected so, will check for available ID now..."));
        end
      end
    end //while()
  endtask

  // ------------------------------------------------------------------------------
  // This task sends several random transactions.
  // num_txn :: indicates number of transaction that this task will send.
  //            However, if it is set to 0 then no transaction willl be sent.
  //            If it is set to lesser than 0 then transacitons are sent in a free-running loop
  // mode    :: indicates type of transactions that will be sent.
  //            0 => both read and write type, 1 => write only, 2 => read only
  // ------------------------------------------------------------------------------
  virtual task send_transactions(int mode=0, int num_txn=0, int port_index=-1);
    bit [15:0] lfsr;
    int port_id, txn_cnt=0, _temp_id_width, stop_indx;
    bit _enable_outstanding = 0, _send_on_read_channel = 0;
    svt_axi_master_transaction tr, _temp_dvm_xact_id_q[$];

    send_transaction_sema.get();
    stop_indx = stop_sending_transactions.size();
    stop_sending_transactions.push_back(0);
    send_transaction_sema.put();
    while(((num_txn==0) || (txn_cnt < num_txn)) && !stop_sending_transactions[stop_indx]) begin
      _enable_outstanding = 0;
      _send_on_read_channel = (mode==0) ? lfsr[0] : (mode==2) ? 1 : 0;
      port_id = (port_index < 0) ? ace_ports[$urandom_range(ace_ports.size()-1, 0)] : port_index;

      // there is no ID dependency between DVM transacitons and transactions on AW channel
      // however, transaction sent on AR channel shouldn't use ID same as any of the active DVM transactions
      // if no IDs are available because of outstanding dvm transactions then wait for at least one of those
      // transactions to finish
      if(_send_on_read_channel) begin
         read_channel_sema.get();
         _temp_id_width = (sys_cfg.master_cfg[port_id].use_separate_rd_wr_chan_id_width) ? 
                           sys_cfg.master_cfg[port_id].read_chan_id_width : sys_cfg.master_cfg[port_id].id_width;
         _temp_dvm_xact_id_q = active_dvm_q.unique(x) with (x.id);
         // -------------------------------------------------------------
         // if all id(s) that could be used for dvm are not available then 
         // wait for one of those dvm transactions to finish so that, the 
         // transaction ID is returned back for further usage
         // -------------------------------------------------------------
         while(_temp_dvm_xact_id_q.size() >= (1 << _temp_id_width)) begin
           _temp_dvm_xact_id_q[0].wait_for_transaction_end();
           _temp_dvm_xact_id_q = active_dvm_q.unique(x) with (x.id);
         end
      end

      `svt_xvm_create_on(tr, p_sequencer.master_sequencer[port_id])
      void'(tr.randomize() with { 
          solve coherent_xact_type before id;
          tr.data_before_addr == 0;
          tr.xact_type == svt_axi_transaction::COHERENT;
          if(!_send_on_read_channel) {
            tr.coherent_xact_type inside {svt_axi_transaction::WRITEUNIQUE, svt_axi_transaction::WRITENOSNOOP};
          }
          if(_send_on_read_channel) {
            (
             tr.coherent_xact_type == svt_axi_transaction::READUNIQUE ||
             tr.coherent_xact_type == svt_axi_transaction::READONCE   ||
             tr.coherent_xact_type == svt_axi_transaction::READSHARED ||
             tr.coherent_xact_type == svt_axi_transaction::READCLEAN  ||
             tr.coherent_xact_type == svt_axi_transaction::READNOTSHAREDDIRTY  ||
             tr.coherent_xact_type == svt_axi_transaction::MAKEUNIQUE ||
             tr.coherent_xact_type == svt_axi_transaction::CLEANUNIQUE||
             tr.coherent_xact_type == svt_axi_transaction::CLEANSHARED||
             tr.coherent_xact_type == svt_axi_transaction::CLEANINVALID||
             tr.coherent_xact_type == svt_axi_transaction::MAKEINVALID||
             tr.coherent_xact_type == svt_axi_transaction::READNOSNOOP);

             //foreach(active_dvm_q[ix]) 
             //    id != active_dvm_q[ix].id;
          }
        });
        `svt_xvm_send(tr)
        get_response(rsp);
        if(_send_on_read_channel) begin
           active_read_q.push_back(tr);
           remove_q_on_xact_end("non_dvm_read",tr);
           read_channel_sema.put();
        end
        else begin
           active_write_q.push_back(tr);
           remove_q_on_xact_end("write",tr);
        end

        randcase
          80: _enable_outstanding = 1;
          20: _enable_outstanding = 0;
        endcase
        if(!_enable_outstanding)
           tr.wait_for_transaction_end();

`protected
FED71O@d4<aT&Z.N_-/8PeD^;T=WTUg_[0HJXdQI:V0aED,O&PHa()@Z5ZEaJ)C=
1_K(GDYdNF<_\S(<,2a)@g[OJJa+&CLO;$
`endprotected

        lfsr = {lfsr[14:0], (lfsr[15]^lfsr[8])};
        `svt_axi_xxm_debug("send_transactions",$psprintf("sent transaction %0s ",`SVT_AXI_PRINT_PREFIX1(tr)));
    end //end while
    stop_sending_transactions[stop_indx] = 0;
  endtask

  virtual task dvm_complete_process( svt_axi_ace_master_snoop_response_sequence snoop_resp_seq[], int port_id );
  endtask 

  virtual task remove_q_on_xact_end(string mode="", svt_axi_transaction xact);
    int _temp_q[$];
    fork
      begin
        xact.wait_for_transaction_end();

        if(mode == "dvm") begin
           read_channel_sema.get();
           _temp_q = active_dvm_q.find_first_index() with (item == xact);  
           if(_temp_q.size() > 0)
              active_dvm_q.delete(_temp_q[0]);
           else
              `svt_amba_debug("remove_q_on_xact_end",$sformatf("VIP_INTERNAL_ERROR: dvm transaction %s not found in the active_dvm_q queue when completed", `SVT_AXI_PRINT_PREFIX1(xact)));
           read_channel_sema.put();
        end
        else if(mode == "non_dvm_read") begin
           read_channel_sema.get();
           _temp_q = active_read_q.find_first_index() with (item == xact);  
           if(_temp_q.size() > 0)
              active_read_q.delete(_temp_q[0]);
           else
              `svt_amba_debug("remove_q_on_xact_end",$sformatf("VIP_INTERNAL_ERROR: read transaction %s not found in the active_read_q queue when completed", `SVT_AXI_PRINT_PREFIX1(xact)));
           read_channel_sema.put();
        end
        else if(mode == "write") begin
           _temp_q = active_write_q.find_first_index() with (item == xact);  
           if(_temp_q.size() > 0)
              active_write_q.delete(_temp_q[0]);
           else
              `svt_amba_debug("remove_q_on_xact_end",$sformatf("VIP_INTERNAL_ERROR: write transaction %s not found in the active_wrie_q queue when completed", `SVT_AXI_PRINT_PREFIX1(xact)));
        end
      end
    join_none
  endtask

  virtual task body();
    int rand_domain_ports[$];
    svt_configuration base_cfg;

    p_sequencer.get_cfg(base_cfg);
    if (!$cast(sys_cfg, base_cfg)) begin
      `svt_xvm_fatal("body", "Unable to $cast the configuration to a svt_axi_system_configuration class");
    end

    foreach (my_system_env.master[i]) begin
      if ( (sys_cfg.master_cfg[i].is_active == 1) &&
           (sys_cfg.master_cfg[i].auto_gen_dvm_complete_enable == 0) &&
           ( (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::AXI_ACE) ||
             ( (sys_cfg.master_cfg[i].axi_interface_type == svt_axi_port_configuration::ACE_LITE) &&
               sys_cfg.master_cfg[i].dvm_enable
             )
           )
         ) begin
             `svt_xvm_create_on(snoop_resp_seq[i], my_system_env.master[i].snoop_sequencer)
             start_snoop_response_seq_for_dvm(i, snoop_resp_seq);
      end
    end
    set_response_queue_depth(17);

    // send random write transactions
    fork
      send_transactions(1); 
      forever begin get_response(rsp); end
    join_none

      if (!get_random_ports_in_domain(domain_type,1,multi_port_type,0,rand_domain_ports) &&
          !rand_domain_ports.size()) begin
        `svt_xvm_error("body", 
             $sformatf("There are no ports for domain_type(%0s).Not executing sequence...",domain_type.name()));
      end
      else begin
        repeat(sequence_length) begin
          foreach(rand_domain_ports[ix])
            send_dvm_sequence(rand_domain_ports[ix],0);
        end
      end
    // wait for all the dvm transactions to complete
    foreach(active_dvm_q[ix]) begin
      `svt_amba_debug("body",$sformatf(" waiting for end of pending transaction %s", `SVT_AXI_PRINT_PREFIX1(active_dvm_q[ix])));
      active_dvm_q[ix].wait_for_transaction_end();
      `svt_amba_debug("body",$sformatf(" ended pending transaction %s", `SVT_AXI_PRINT_PREFIX1(active_dvm_q[ix])));
    end
    // stop sending more transactions now
    foreach(stop_sending_transactions[ix])
      stop_sending_transactions[ix] = 1;
`protected
:F2:W?B8eA00?(^WGHKCUaQ@d^2f/K>=8</[C504>I,3I+J)TN(K1))\]QI@[,C)
1J6#deT[BO8[MH\?e98;5;Q@7$
`endprotected
    
    foreach(stop_sending_transactions[ix])
      wait(stop_sending_transactions[ix] == 0);

    foreach(active_read_q[ix]) begin
      active_read_q[ix].wait_for_transaction_end();
      `svt_amba_debug("body",$sformatf(" ended pending read transaction %s", `SVT_AXI_PRINT_PREFIX1(active_read_q[ix])));
    end
    foreach(active_write_q[ix]) begin
      active_write_q[ix].wait_for_transaction_end();
      `svt_amba_debug("body",$sformatf(" ended pending write transaction %s", `SVT_AXI_PRINT_PREFIX1(active_write_q[ix])));
    end
    wait(active_write_q.size() == 0 && active_read_q.size() == 0);
  endtask

endclass
// ---------------------------- END OF DVM Sequences ---------------------------------------------------------
// =====================================================================================================
// ---------------------------- ACE 2.0 Sequences ---------------------------------------------------------
/**
  * #- Send a sequence of READONCECLEANINVALID transactions to consecutive address locations
  * #- The port from which the transactions are sent out are determined by port_id which can
  * be passed via config_db. The port should be an ACE-Lite port.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_readoncecleaninvalid_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence readoncecleaninvalid_seq;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_readoncecleaninvalid_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readoncecleaninvalid_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 0;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    super.pre_body();
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    // Check for valid port type
    begin
      `svt_xvm_create_on(readoncecleaninvalid_seq, p_sequencer.master_sequencer[port_id]) 
      readoncecleaninvalid_seq.readoncecleaninvalid_wt = 1;
      readoncecleaninvalid_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      if (status_start_addr) begin
        readoncecleaninvalid_seq.status_start_addr = 1;
        readoncecleaninvalid_seq.start_addr = start_addr;
      end
      void'(readoncecleaninvalid_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                    });
      readoncecleaninvalid_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      readoncecleaninvalid_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass

/** 
  * This sequence initiates ReadOnceCleanInvalid transaction from the ACE/ACE-Lite master
  * specified with port_id , which can be a random port or a specific port
  * configured by the user through uvm_config_db.  ReadOnceCleanInvalid transactions can be
  * sent only when the svt_axi_port_configuration::axi_interface_type of the
  * master corresponding to port_id is set to
  * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
  * Before sending ReadOnceCleanInvalid transactions, cachelines of peer masters are
  * initialized to random, valid states.  Initialisation is done through front
  * door access, by sending specific transactions from the initiating master
  * (corresponding to port_id) and peer masters.  Please look up the
  * documentation of #svt_axi_cacheline_initialization for details.
  */
class svt_axi_ace_master_readoncecleaninvalid_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readoncecleaninvalid_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports, ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readoncecleaninvalid_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction
  
  virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READONCECLEANINVALID ,1);
      // Wait for readoncecleaninvalid transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_readoncecleaninvalid_sequence

/** 
  * This sequence initiates ReadOnceMakeInvalid transaction from the ACE/ACE-Lite master
  * specified with port_id , which can be a random port or a specific port
  * configured by the user through uvm_config_db.  ReadOnceMakeInvalid transactions can be
  * sent only when the svt_axi_port_configuration::axi_interface_type of the
  * master corresponding to port_id is set to
  * svt_axi_port_configuration::AXI_ACE or svt_axi_port_configuration::ACE_LITE.
  * Before sending ReadOnceMakeInvalid transactions, cachelines of peer masters are
  * initialized to random, valid states.  Initialisation is done through front
  * door access, by sending specific transactions from the initiating master
  * (corresponding to port_id) and peer masters.  Please look up the
  * documentation of #svt_axi_cacheline_initialization for details.
  */
class svt_axi_ace_master_readoncemakeinvalid_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;
 
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  `svt_xvm_object_utils(svt_axi_ace_master_readoncemakeinvalid_sequence)

  constraint valid_port_type {
    port_id inside {ace_ports, ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readoncemakeinvalid_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 1;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction
  
    virtual task body();
        
    // Check for valid port type
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
    end 
    else begin
      super.body();
      send_coherent_transactions(svt_axi_transaction::READONCEMAKEINVALID ,1);
      // Wait for readoncemakeinvalid transactions to finish
      coherent_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass: svt_axi_ace_master_readoncemakeinvalid_sequence

/**
  * #- Send a sequence of READONCEMAKEINVALID transactions to consecutive address locations
  * #- The port from which the transactions are sent out are determined by port_id which can
  * be passed via config_db. The port should be an ACE-Lite port.
  * #- The start address of the sequence can be passed through a uvm_config_db for 'start_addr'
  * If no start_addr is passed, the address of the first transaction randomized in the sequence
  * is taken as the start address of the sequence. <br>
  */
class svt_axi_ace_master_readoncemakeinvalid_sequential_sequence extends svt_axi_ace_master_single_port_base_virtual_sequence;

  /** Read sequence */
  svt_axi_ace_master_generic_sequence readoncemakeinvalid_seq;

  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)
  `svt_xvm_object_utils(svt_axi_ace_master_readoncemakeinvalid_sequential_sequence)

  constraint valid_port_type {
    port_id inside {ace_lite_ports};
  }
  
  function new(string name = "svt_axi_ace_master_readoncemakeinvalid_sequential_sequence");
    super.new(name);
    is_seq_valid_on_ace_port = 0;
    is_seq_valid_on_ace_lite_port = 1;
  endfunction

  task pre_body();
    super.pre_body();
  endtask: pre_body

  virtual task body();
    if (!is_supported(cfg)) begin
      `svt_xvm_note("body", "The sequence cannot be run based on the current system configuration"); 
      return;
    end 
        
    // Check for valid port type
    begin
      `svt_xvm_create_on(readoncemakeinvalid_seq, p_sequencer.master_sequencer[port_id]) 
      readoncemakeinvalid_seq.readoncemakeinvalid_wt = 1;
      readoncemakeinvalid_seq.addr_mode = svt_axi_ace_master_base_sequence::SEQUENTIAL_ADDR_MODE;
      if (status_start_addr) begin
        readoncemakeinvalid_seq.status_start_addr = 1;
        readoncemakeinvalid_seq.start_addr = start_addr;
      end
      void'(readoncemakeinvalid_seq.randomize with {use_directed_addr == 0;
                                    sequence_length==local::sequence_length;
                                    });
      readoncemakeinvalid_seq.start(p_sequencer.master_sequencer[port_id]);
      // Wait for transactions to finish
      readoncemakeinvalid_seq.wait_for_active_xacts_to_end();
    end 
  endtask: body

endclass
// ---------------------------- END OF ACE 2.0 Sequences ---------------------------------------------------------

/**
  AXI VIP provides a pre-defined AXI ACE Master sequence library
  svt_axi_ace_master_transaction_sequence_library, which can hold the AXI ACE Master
  sequences. The library by default has no registered sequences. You are
  expected to call
  svt_axi_ace_master_transaction_sequence_library::populate_library() method to
  populate the sequence library with master sequences provided with the VIP. The
  system configuration is provided to the populate_library() method as an
  argument. Based on the system configuration, appropriate sequences are added to
  the sequence library.  You can then load the sequence library in the system sequencer.
  

  The user can also add user-defined sequences to this sequence library using
  appropriate UVM methods.
 */
class svt_axi_ace_master_transaction_sequence_library extends svt_sequence_library;
  `svt_xvm_object_utils(svt_axi_ace_master_transaction_sequence_library)

  //Required to allow new_item() to have access to the parent sequencer
  `svt_xvm_declare_p_sequencer(svt_axi_system_sequencer)

  //Removes all registered sequences from this library
  extern function void remove_all_sequences();

  /**
    Populates the library with all sequences defined in
    svt_axi_ace_master_sequence_collection.sv

    @param cfg User is expected to pass a system configuration to this argument.
    Based on the syste, configuration, this method adds the appropriate sequences
    from the ace master sequence collection to the ace master sequence library.
    */
  extern function int unsigned populate_library(svt_configuration cfg);

  extern function new (string name="svt_axi_ace_master_transaction_sequence_library");

`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task execute(uvm_object_wrapper wrap);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task execute(ovm_object_wrapper wrap);
`endif
endclass

//-----------------------------------------------------------------------
function svt_axi_ace_master_transaction_sequence_library::new (string name="svt_axi_ace_master_transaction_sequence_library");
`protected
#cQ^GgPe]I_O=J;W0W[V()e;--W=/,Q>F_9^;7>948K#L.+,JdV,+)DT\73Ged3D
9,.bBXD<18B@.1+f<01CE=XGKGgfJH,B?$
`endprotected

  init_sequence_library();
endfunction

//-------------------------------------------------------------------------


`ifdef SVT_UVM_TECHNOLOGY
task svt_axi_ace_master_transaction_sequence_library::execute(uvm_object_wrapper wrap);
  int sts;
  uvm_object temp_obj;
  uvm_factory temp_factory;
  uvm_sequence_base seq_or_item;

  temp_factory = uvm_factory::get();

`elsif SVT_OVM_TECHNOLOGY
task svt_axi_ace_master_transaction_sequence_library::execute(ovm_object_wrapper wrap);

  ovm_object temp_obj;
  ovm_factory temp_factory;
  ovm_sequence_base seq_or_item;

  temp_factory = ovm_factory::get();
`endif

    temp_obj = temp_factory.create_object_by_type(wrap,get_full_name(), $sformatf("'d%0d",sequences_executed+1));
    void'($cast(seq_or_item,temp_obj));
    seq_or_item.set_sequencer(p_sequencer);
  `svt_xvm_debug("execute",{"Executing ",(seq_or_item.is_item() ? "item " : "sequence "),seq_or_item.get_name(), " (",seq_or_item.get_type_name(),")"});
  seq_or_item.print_sequence_info = 1;
  if (!seq_or_item.randomize()) begin 
          `svt_xvm_fatal("execute", "Unable to randomize the snoop response");
  end

  seq_or_item.start(p_sequencer);
  //`uvm_rand_send(seq_or_item)
  seqs_distrib[seq_or_item.get_type_name()] = seqs_distrib[seq_or_item.get_type_name()]+1;

  sequences_executed++;

  //super.execute(wrap);
endtask

//-------------------------------------------------------------------------

function void svt_axi_ace_master_transaction_sequence_library::remove_all_sequences();
  sequences.delete();
endfunction

function int unsigned svt_axi_ace_master_transaction_sequence_library::populate_library(svt_configuration cfg);
`protected
g3B5:a,KD(4,ZW@@9(P2-I&=P\c7X5DS/aR\<@OgO[bI=CKdTW?<-)g&92gQ,<GR
2H5R2:e,E@(>G+cY@c1&dS6W2#CPTP^MW?V2FJ##_.2RZ5UT0\ce)_T#UP<LBH0c
182CF@Ib9fL5C?MS_+:</\>?H7ZLN)fC>HKbJYYeJ2Qc,XB(\b.Jeb;0ZJHMSPTJ
KD@4Rg;NT4cGYaWA0^O\>?X]DM:6^WK1)>^X1^.cWQ;8PZAJfAZU@L.bUeI3@^7I
<NB@,ffFRWBcFOJ,#:EMQBU3+YYT,)S]9).N;[gW5#\V0^gTV[eYeE+JM(@^HY#>
,K=S8#H;1/G?&cF+W;[K^^/)HgHca=WZf30=6dWeR&<f?FKZGf>OaE3?;Zc5L.3@
CbeRT7SY.CX8R+[D+Q-,G]U/]ZV<7E60ZS:BLbcE@-e6PQ>?_P)<)&Y#WdAF<BOF
#OB35Q39V/0I7\_:\@V8ZZeEAK5M[)aG#)cSFG:ADIV1,=[EA35B.fb3(P\ab<2c
M0G5D?bMMEF5[?bZFFV85OEYg?1Z&&^b]d</I^4c327cL)<)/-NJ^d8^9)beU,0=
>]Gg>Z4T1/cVTSbIC?B2d;^<A+[HK:J2R_=J4F:ERB7B(V_A(&e6.MPO.48JedUf
_PFW[=HHE[#D-1V7\;(d3T9Y9A@;@3RF.ZMAYWAXSBWYNM1PINcaMTSNP9Y#C76<
#C=ege-56D<a58,^O3WS/68]21)dE<-0BH-=.LcaQY84]Hb&CI8(90H.@A,,RE4]
:e8BeZ8+&]a)?=;((M^4GcW8YQ(@gV]\6=.#6=:B+E&aM\V8aL\L?@M&a(1R5@aA
7H^R4BSHIO=)\^H;)KO>#WK>-FfD;QDUc3XS(EHZF@5C_()<4.a]/5_[EQ>[(-(B
P8Z@:QQH&^?fTRWa.1fSJ<>LGDQTg,c-ZcP>0I3gKEH:UTgJ4E8=^&8.g;JEQ,XB
2Q;20cWGBIG:HQ[YQBIgb^5Gf[0.(N@A\J&eYNg/\T;1:8DG_6=.C@YVKV2b],2c
a?7F/cM(bQJC,Be7SD]^Q[<59Z.]A^RCPLb6JC79#b#?G/4EWaDJD?&]BDO).D#C
<NXN<c=T6&G^=Tg,0@HO,]4]g#H#/E+EaO+d/:T?R,&\J,B?22gSY8a^Y==DRGMI
+O7;Y;NaB(SJ?E^R35?&##[[:3Ucg\FS.DR?TXb5b<63::D9F[O[4W3b1(>J&Z3)
=#<C##U(=+G2E,1KB:g[dZ3#K]BPOO\YU^9D\Q^^;&3J4:IWA3^6MM&,3LIR>3TL
)dY&f7#4BZFJ7NW96gMBU\:)(8Kg3,;S5DYZS)JK&]M7_Y?g>3KND7+V,0VRWT-8
g&aH;EVLRWb9bVO70ELR0CA=RY[QWdLAgNI1R13R88XEZK,-dSgXQJ_G,A\#=@f2
RC?/X_gN.^LRYFc+?/X_6;>4^@#9>9#Z)d[KM,,+<:fKf8/CZS=BRA(Og+?(0P7Z
JY9ILEUQ>fN<_AV(1O0LZMdb&I[ZV;Fb4J#<[OS1cRU43JJFd->d)O6Y)1S-(2D<
+8>SO_T57@fc:KOPdLPP?E5V7+4(E&T8c<_L4\Vgb?-,NRO.f98E,?U56#AN=FUc
:<;3?AV/;U1S<7[DR5[M[M3/&/ZSK<YDg;L;OJ-D/<A7]S.EReRe>UdA2+@Z<4M2
gIOIeRE^QR^9\J<AB3V@56#C5K.eXe9\F>BAG4fB?6SAWO)aNIA@[DE>9PF<cZ\S
<)GMU-3T^.5>K#T/6;IUC[OHIT7Y[376VU<-/6M9N;/cWPGaJR5YD5B+6(98FYBW
[WT7/#=(T<?XJ3&OBA8?AAN\V_@6MD>GL5R3e>a291fN.F3gGgY+&W^]OCOD-FPU
/HME=_cD9I(<(@T3_gUZSM1&@KeKMgE&/f9GZV9]>2BD]P=SJGc,5LG&2(&4X1V<
_Pd&IFSLUTLE_F6g>5Xd38ZZ?U;(OT#YKDUHT9I1_3d.6HL=0.H?(a6E(QS^&WK=
LHWO7dI>&NQVeVO5M/3fab27-J9ENKZ)?+K5L#7MXXC].MIY4G<eM;/L?g1FX2@=
#(_>ZQG;J+C4,-7QIeQ_bV>D8O<95]\&D/1)+Y-MbFf#-@HZ/EWaC]EM_BS:T)=G
H8L9@XWB>/a0.3U[=.[GB(SEX5M)EAf-Q9LB@0O\>I8#]_K<NH/A.2Z_^KFLNP3B
PGTQN60#12)J2R\9&@62B^TKH47X0Pa7CF:O)f0+1bQd3.(NWW@<B<&7\37I:#[Q
2;c:08,76<@<GZ7-Zf1e/;#\Y?R<[[GfM8fIDgU5&23)U239Aeb)d=BLd_]bLT4F
,gE#e.&._S&2,TTDKMfKcZS2RAXS1>9OJFU:B]V=S<E+H<cS/K=YW[?-8Y=6M=87
8?KH8QR5[3N3;4O9a4<F#?a&COJ;]_BUV0U,V=L].Ff>g\E.0:BDH7PB[E#@),=R
OTF[@^gZF@T(bd3B_TOg&/(CMF#V;&G>.S;A\GFIHbV.eKc(;d+J(ePBN$
`endprotected
  
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_exclusive_access_virtual_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_snoop_during_memory_update_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_two_master_concurrent_write_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_read_during_coherent_write_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_overlapping_addr_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_shareable_store_barrier_load_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_nonshareable_store_barrier_load_sequence,populate_library);
  `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_load_barrier_sequence,populate_library);

     // added following sequence in populate library for the purpose of SVDOC ONLY
  `ifdef __SVDOC__
  `ifdef CCI400_CHECKS_ENABLED
    `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_cci400_reg_config_base_virtual_sequence,populate_library);
    `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_cci400_perf_mon_reg_read_sequence,populate_library);
  `endif
    `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_exclusive_access_sequence,populate_library);
     // This sequence is not added to the library (except for documentation) because it kills any
     // snoop response sequences supplied by the testbench to run a dvm specific snoop response. Adding
     // it to the library and running it may cause undesirable results and therefore this sequence must 
     // be run in a separate test
    `SVT_SEQUENCE_LIBRARY_SAFE_ADD_SEQUENCE(svt_axi_ace_master_dvm_virtual_sequence,populate_library);
  `endif

endfunction

`endif // GUARD_SVT_AXI_ACE_MASTER_SEQUENCE_COLLECTION_SV
