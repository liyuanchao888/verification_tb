
`ifndef GUARD_SVT_AXI_IC_SLAVE_AGENT_SV
`define GUARD_SVT_AXI_IC_SLAVE_AGENT_SV

typedef class svt_axi_port_monitor;
typedef class svt_axi_port_monitor_common;
typedef class svt_axi_ic_slave_response_sequence;

// =============================================================================
/**
  * The slave agent encapsulates slave sequencer, slave driver, and port
  * monitor. The slave agent can be configured to operate in active mode and
  * passive mode. The user can provide AXI response sequences to the slave
  * sequencer.  The slave agent is configured using port configuration, which
  * is available in the system configuration. The port configuration should be
  * provided to the slave agent in the build phase of the test.  In the slave
  * agent, the port monitor samples the AXI port signals. When a new
  * transaction is detected, port monitor provides a response request sequence
  * to the slave sequencer. The slave response sequence within the sequencer
  * programs the appropriate slave response. The updated response sequence is
  * then provided by the slave sequencer to the slave driver. The slave driver
  * in turn drives the response on the AXI bus. The slave driver and port
  * monitor components within the slave agent call the callback methods at
  * various phases of execution of the AXI transaction. After the AXI
  * transaction on the bus is complete, the completed sequence item is provided
  * to the analysis port of port monitor, which can be used by the testbench.
  */
class svt_axi_ic_slave_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual `SVT_AXI_MASTER_IF svt_axi_master_vif;

`ifdef SVT_AMBA_ENABLE_C_BASED_MEM
  //Memory core 
  local svt_mem_core mem_core; 
  
  //Default Memory backdoor  
  svt_mem_backdoor backdoor; 
  
   // Memory configuration 
  local svt_mem_configuration mem_cfg; 
`endif  


  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AXI master virtual interface */
  svt_axi_master_vif vif;

  /** AXI Slave Driver */
  svt_axi_slave driver;

  /** AXI Monitor */
  svt_axi_port_monitor monitor;

  /** AXI Slave Sequencer */
  svt_axi_ic_slave_sequencer sequencer;

  /** AXI slave coverage callback handle*/
  svt_axi_port_monitor_def_cov_callback slave_trans_cov_cb;

  /** AXI Signal coverage callbacks */
  svt_axi_port_monitor_def_toggle_cov_callback#(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport) slave_toggle_cov_cb;
  svt_axi_port_monitor_def_state_cov_callback#(virtual `SVT_AXI_MASTER_IF.svt_axi_monitor_modport)  slave_state_cov_cb;

  /** AXI XML Writer for the Protocol Analyzer */
  svt_axi_port_monitor_pa_writer_callbacks slave_xml_writer_cb;

   /** Writer used in callbacks to generate XML/FSDB output for pa */
   protected svt_xml_writer xml_writer = null;

  /** AXI Port Monitor Callback Instance for System Checker */
  svt_axi_port_monitor_system_checker_callback system_checker_cb;

  /** AXI Slave Snoop Sequencer to supply snoop transaction to be driven to the master snoop channel */
  svt_axi_slave_snoop_sequencer snoop_sequencer;

  /** A reference to the slave memory set if the svt_axi_slave_memory_sequence sequence is used */ 
  svt_mem axi_slave_mem;

  /** Reference to FIFOs in the slave. These are configured based on
    * num_fifo_mem and fifo_mem_addresses of the port configuration 
    */
  svt_axi_fifo_mem fifo_mem[];

  /**
   * Implementation port class which makes the snoop requests available 
   * when the interconnect initiates a snoop transaction to this port.
   */
`ifdef SVT_UVM_TECHNOLOGY
  uvm_blocking_peek_imp#(svt_axi_ic_snoop_transaction, svt_axi_ic_slave_agent) snoop_request_imp;
`elsif SVT_OVM_TECHNOLOGY
  ovm_blocking_peek_imp#(svt_axi_ic_snoop_transaction, svt_axi_ic_slave_agent) snoop_request_imp;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /** AMBA-PV blocking AXI response transaction socket interface */
  uvm_tlm_b_initiator_socket#(uvm_tlm_generic_payload) resp_socket;
`endif

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  /** Configuration object copy to be used in set/get operations. */
  protected svt_axi_port_configuration cfg_snapshot;


  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** @cond PRIVATE */
  /** Configuration object for this transactor. */
  local svt_axi_port_configuration cfg;

  /** Common features of AXI Slave monitor Component */
  local svt_axi_slave_monitor_common monitor_common;

  /** Common reference handle for common in active and passive modes */
  local svt_axi_common common;


  /** 
   * A mailbox to hold the snoop transactions created by the
   * interconnect. A snoop sequence could call the peek method
   * of the snoop_request_port. The peek implementation will
   * provide the snoop transactions in this mailbox. 
   */
  local mailbox #(svt_axi_ic_snoop_transaction) snoop_req_mailbox;

  /** slave agent instance name. */
  local string slave_ic_agent_inst_name = "";

  /** AXI External Master Agent Configuration */ 
  svt_axi_port_configuration axi_external_port_cfg;

  /** AXI External Master Index */ 
  int axi_external_port_id = -1;

 typedef bit [(`SVT_AXI_MAX_ADDR_WIDTH-1):0] _addr;

 typedef bit [`SVT_AXI_MAX_ADDR_WIDTH-1:0] max_addr_width_data_type;

  /** Associative array which used to store the write data check parity values. */
  bit [(`SVT_AXI_MAX_DATA_WIDTH/8) - 1 : 0] datachk_partiy_assoc_array[max_addr_width_data_type];
 
  /** Assoc array to hold the value of poison in case of ACE */
    bit[(`SVT_AXI_MAX_DATA_WIDTH/64-1):0] addr_holds_corrupt_data_with_poison_assoc_arr[_addr] ;

  /** @endcond */

  
  // ****************************************************************************
  // UVM Field Macros
  // ****************************************************************************

  `svt_xvm_component_utils(svt_axi_ic_slave_agent)

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function new (string name, uvm_component parent);
`elsif SVT_OVM_TECHNOLOGY
  extern function new (string name, ovm_component parent);
`endif

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Always constructs the #monitor component. Constructs the #driver and #sequencer
   * components if configured as a UVM_ACTIVE component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif
  // ---------------------------------------------------------------------------
  /**
   * end_of_elaboration Phase
   * A local factory is used for all construction within the VIP.
   */
`ifdef SVT_UVM_TECHNOLOGY
 extern function void end_of_elaboration_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
 extern function void end_of_elaboration();
`endif


  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase 
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif
  
  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  /**
   * Implementation of the peek method needed for #snoop_request_imp.
   * This peek method should be called in forever loop, whenever interconnect 
   * initiates a new snoop transaction on this port, the peek method 
   * gives out a snoop transaction object. 
   * Blocks when interconnect does not have any new transaction.
   *
   * @param snoop_xact svt_axi_ic_snoop_transaction output object. 
   *
   */
  extern task peek(output svt_axi_ic_snoop_transaction snoop_xact);

  /**
    * Writes the given snoop transaction into the mailbox used
    * for storing these transactions
    */
  extern task write_to_snoop_mailbox(svt_axi_ic_snoop_transaction snoop_xact);

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /** 
   * Retruns the report on performance metrics as a string
   * @return A string with the performance report
   */
  extern function string get_performance_report();

  extern function int get_fifo_index(bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr);
  extern task put_write_transaction_data_to_mem(svt_axi_transaction xact);
  extern task put_read_transaction_data_to_mem(svt_axi_transaction xact);
  extern task get_read_data_from_mem_to_transaction(svt_axi_transaction xact);
  extern task write_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, bit[7:0] data);
  extern task read_byte(input bit[`SVT_AXI_MAX_ADDR_WIDTH-1:0] addr, output bit[7:0] data);

  /** @cond PRIVATE */
  /** 
   * Returns the name of this agent
   */
  extern function string get_requester_name();
  /** @endcond */
//vcs_lic_vip_protect
  `protected
4.0EJe?[0_(X_C)4)&35e&OJA5O60D=,1=D(GPR(5HOMIOM^HeW,0(11bZ3;Wg4a
=XDRVGP^6S;#ecB,cZD>:=R]44/TC.Xc01,A4AMVJFK:3)6a5IbRG@[[=[(50TJP
]R(AMGBX<6X,3@G3eSK5cLfE\\A1N[9QHb#L^7:<@8;I\_-)bMcI33&9WGAaaT38
+gQRTbK8S,OV5;^&J_CX?2YaU/;.MCMbLG@@5.5W#:KXe7>PA,I\c/TbAD3=8Ja3
_<^.eE/PD_^C2=gR/2f=.:DJ_Xf^IGFWX-3]6C9;gP3SKGJ62UKIGGU[JF,QL2#d
KEJQB1)<F(4:8+GD5g;.>&3d//,Z/8FR4CBZJ;,]SS#[#/.?/01F<+#7KfQUS@/P
&E7EP>R[cWde<]391JO3+b/&[Z)B/X/BJV.g/^ITXL-^Q(=CHONEY#/G2OQY1eeF
KbbTP>.WWXdBSS&+-RPB9AaPg1cSNR8_2BDbaKOFd7V]<L7/=.Z\E^/-]53@cQIR
6e&b63YbC.GB/$
`endprotected


endclass

`protected
PC[Q-EfEQ0@9(YYc=Y93gZ8c6].QddT[L-GeH?F1N900=Zd_NfJO5)48XXfIKcXX
1Ba1<@T(RE6P[&OEQbDQ;AS[]]eXR2ZC,PU\EJ1.KNbXQg)@D,L?]/JB<=HCSaa/
DeGH?[4_[22::2VY;6:KC2BPDPTS_#VJQWBPD=2H@E]TY>U.dNF9Q1baDK@MFU3]
94P-<e8;;=OGGC0ePaKH_Q#1Y(GZ5XG,\8TJR/d&Q^.IFHd/[:DO8X]c;.J<L0DK
O161\6,b)e.2_,Q#Kb61.g4N_FSEOH&LCfe-X&>4#\ZaU1<VAPe5?G7;C??.BEIC
M7ZHHY6.=6EEcbYA<N#1QT2-P(^WPP61GbB.N=3f8<UaM<2^>c>eQ1F8-+B2UN?>
FcY/P&<XPe6T,_O+;TS\.1LY6;1(6bJIOYe[J8-_T#XN,8[&:(3P&eNN>(;GCe9b
3J0:NF1<X3ER,H?7FZWSDQ8JZVdULF8UaX[KO\JXB]eU95MFR;W+;X,NgE=WJ/XI
cSa4(]4\S=A+OcSW16ZR-WcV)5;BAZ?HGg)LW=C>5>0[]g&H-OT+DAUE\1RfCVD+
e<2F5#:H?6K)I@]IG;.XaLSb)bU[XDQ>&]^8\7]DQ1N^O-4.-M<c:?IS^#SI7JWUS$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
H[,LQ&KXB?2)>5eGA=5E#^e0@5KM?TAXVd1VcD,FF4\QS9X(&O+K.(\+F-18MI(6
cVOg3_Y,Z7Q@N97I>:)-/dN?b@&ZO]4O2E>LCFB(-RPfTDFVC)a_OTd1+:1^;W,6
(?T?49;_K)KQg1R\/5R\\(LHH+M^O2I:U/&?3PJHV[#9=S1d;1d7(UY8W\0.FHNJ
D)[Cb<B;IVbBP\IdCH,GL[:KDNBN0]-1JOfBD9dLeB+T:J).1K;bWba2F^bY,e=9
0?G>b,6Q#Wf^>;AL=6V&fS4c?;3H(=K=4&.fF63AW+-gVHUd+P])KO?EIa_J>3JF
E<#U-EdN_bEX3L\C63H(,_2#LHD89,\[Y(bN5\CN8dY\DgY7bSaI;LbR.\Gaf]gG
g,+)\1B+UPDTFJ(dH3fHSOSV_:168c)2G:+H;EL,LA;Y(#-OI>>9U5R,(A<;XQ=g
Z/WF6TRG;&U78W+^egf).-.ZU](QD+bC9Zb7&19I5D8ZO,B7L<NVOKB:gBFZGF((
W76D(#RDV(:QO6F0OY^7bgPRHLJ(S&K&_WbN[Q<4Y[EX]3:L&G0R<,_29gfJ@-8-
F9I#c9L48-Q00QWCP+6U@2d=4X8[<K/+MU7SHJV5gRB-TY5[U+bXbeGdS-Naa6M)
7RU:DFOW,)]DV1Rb_508Scf(P_:@&_Q9AYD[&2--?CeV-L-S-J2<)&.;?Yb;M^D3
MeK9f.eMF9S9.\;3UQ3,-Y5F-De5#b87.C)W/A>DO:M)^XH-a<A.\326b)D8?E51
,[4?NIS-?e3.89LC[-J#3-VP.cC#0G+R8D(G/J)X,HSY408<K21WKB_Fg,Lb?PDD
(aVQ&97:ff-8Pg0+/R;DD9Z84?8P_d5(?ACR=5Z7TT+,)T9EWQCRWH)O^6CZWN7;
D=+T)fNaJLD5<\P=ZM8CHEGLCPZHe2.?8S9?74LYddL\2[8_4CdL+].4WSa+T;(H
I\?3B_#ff^&dM/,^-eU8WBJ:b:JY^,SME.b3U:OJ2TB+_ea+BLLFQP;IeFE)dPaH
L]UPYOg?&]aOBK]+?\Y<J#\I7;1VQMLcDT\gH^b_[C4,L@Y4@X)Mcb9M0fc\f]=V
GDBFXMP5&F391J2GWdH4UB]<YFD?C]9#ADS2&4CeEc/eI6Le_EbNI?]gV5_V+7(d
OOGEL>;>I\FF]L,=c=B<<+?JS>F2E_=X>?<#g.aI4ZL+1b12P?1#-6(1H,(f0M2f
Ne1-Hc;NR69.(L/XUGPO02GEgOFU@8F9:Y.\g-3de&eF5EeG\X\^K0N3&;a\\R/L
9#c,-R:LV3aK&BNP7RV9fL[=g3;_d2N_aD.)bb6-E\<P)g3W9C8G5E@>8L+<=:\)
:R.-AOBGTW5d^.#gGZKO5+SKAPcd-X-K\[eJ,6D2dBTQC/)R=-(IX=-;Ag\bKD8F
#;Y?<M(1aMA4:_\fXcM?]_Y=#H3NGbY5]T?6Vg1T:)6SXe+;\_gZ9LBCLW\KRfJ@
4DSN]\L<+\C:TE_@A([MfN7Y/;#,J=YZ[.g,2;3P<\=\ZXY9#gbWI9MPbG#4E5S(
H@N\e06Bc)gH(7,63]ZNZ=K#(M65547L8&TaQAa2d&4W?RRU)V@C:=+&cZHVUL\&
933V?b^:eTB;ZKe8K4GGA5SdAcY[AE2N+0T09;1JI<a3D:\/A5Q:Z57.#=:\7&7b
G-?g+@F,S.EHQVZULeE,B7+2ab1OJO=-(F:FT^Y2O7,/&14=(C1XcJ[ELe8BU.P^
E.96Ue1N6^VME\74?fL;)]H<cKR0&+YJM+GJ742=a7P:J[Y;?\O4a9Kd:@G:7&g;
[\UUD0L<M:K/A22@GKc>X7E@A3HK:/T_,Cd0eW3G.P[NP>AaOCZDcWA8BP:Reg.2
(1]>E;fBC\;UZ=,TgW;9AAfGTbB++MFTL7QM(90S)]T6>S+?afb5&KWOG(D3;+UD
^?9a(+a67W/A^WH.PfFGQ.5]&;3[I;bRF?G@@C.G3REPPST&d71BV6JA@_W-3Hf(
+EJ97XH5>8C/d7Xf.-UDC,WO(S67KQU#/[=1H)F3/7S[U7HR-K-5MMeeTdYKFZ6)
^SbcR@S2>,JNGLB&JQ830G?Y[^_K4\b_HJb-4dcI]d+d[PW3TcEI6aEIG^c4e[f,
EWK6#DDK-\B0,E0=A\TBBe6dO7=+^(_&<_4Dd6c;3dSBA/XNP@gM@(],?7R/AQ1E
T&5HH33<HY^L:PEIC4^=8(#JH/8FY#LFG3D6(&J;BZP)\[/DS@L:W&M_21N#3FR2
Tc46K98Q8\&::5<@\).CU?>)7^fcY,[LA9Y^0F(eA5a8TPaREb6[:QVA/TZ>gT;:
P-8U/Y.N:F5^[S5POQW_)3T_)3A+4@XX\K<,d/P<O@5@deX<H>>9.[0W](S=IYTN
V([\AaXPNPA>HJF_<RNUdPH-F3FMZQ;F=J\0=)XVSQ)f:]_@#P=4A?D-+-QPIEH\
(RCLSV>/+2:^;_XVLL7#QdQaCQ0QebNSLaLYKYC&AJ@Rd+X3e4M<G=18]B=RMS))
EaW@UEG#+SeT[#ZG^AAIIY^/df/RZEd#V,0FY;SPV^G&5Xc4X;WGG\@B-ZU6b_=-
J^#3R5DVUD4^\6LIbCS.(BD8FBYOWSeH[\K:9#P7Z8KJ_DcYN5,gZJ;5AWHRX>HM
0<3PUI/;K<Q5L48<C):9?=#NK;+Hf5A68YfTGYO.F\;(5@V6A7fLK>W\44>d5-39
;e+AN8>>+1ID\O)3Jg4eN2f5A\#e[)\C(TW;B#L+5Q=g&AN&<SNQY@T>cGg@ag;@
VY[JX^b29K(]M-_ND]8-+bO]FR>_gb]U(^R9.NB4YZP=;,-(?UR@[f&R_N-F,e5a
9R6-VHJ[ZOO(ZV8OOX+[11S?aUe)&DM94&C,0fU^+<H7C@dE17bM.[1gXa8_FDg]
S#J1_I;SNZgJf#4+g1S2+HDO8N.?R]8B..L;8/DXe=34P=facXN_(F97>4Xg75.X
PKL4.I-PN&O7Ve1ecNdJ[O=FJ5I?5YOdP9aKQ04,M_/MICE^@&SITS^V^0<:VWY6
?I#8,9VCCJbT2:S_E:eMBQaXcdeAdTK)_-a-fYdZ[dCT8b[61??)0b4O]E,9R:>6
JLdcBCIJOWDFDENI17#2):#9YXaCfG-Y(@-^2e&e@:ZWd&4/G#(+2Gg_36BYK](E
;Y>S7MW2;M=cIVXHO;a:Vg5TZg-@df_5DJbGaTX(VEEeHVBY<^LG.5Lg&HedO_95
-[4a)6.bFUJ>+0a:-]#,2))N^Fd^IM1A59N0SV,,L+;>FUK3[eE17?O[93L&fF9,
1cdZ3,OST-8]P:ff3D\[QB)9#20<:K0P#82=I8NG+VL#U<;I0SBM=)=K:4&5e4M6
e1JYe,gJQ@TDLQ3<NT+daTIK3Sg39]4RB4W#(VIX[IJgaLIgeW:YEUG[I1UM3HK2
)(aJ&H3<6GbR>5X4?&D<^-/(gJcQCVdJW(.,#3G(TH/E/-+>KA_SE0MQU]5b_KdF
NRN42[#)H]2]SXI\XM;9UK>c0;1/5XcO3bG_VI)N&PGYOF,U&34]HA0+K5.g_D4#
e=9,KX20\fZ6Y3P4;-Z/C,A]AQ,X+d,cOU0CC.Xg<JU<(]?^,&b/RLMdZ;>P>O5C
<)RD>,@;&d,;RG3BP]ESS7De9C6\7Y\2fd:YNGIL5MSH>G_E/,.O]->dM8I#/.8^
W45>]OgVN4D\2EHQSO-43e3XS^&,gQ,FAISZ)<8VWJK]=TK-2H72a703T9:>8[E<
\b885^NU8PU)T>WGQ991:\J?EeL5MN7(\5.a(aX@L-RG:bMI+)YB].6^OD6_8=bU
;1#UDX\<P7J0#Q.<0J>4^X7dJ>U=1A<W\;6MM&e_34S\N9LRHKSL>.3<FBD4?R#:
CV[Aa3VdbLf^E#@)1P7d_WdJcHL4dS\Vg^0N),<OL@+@Gd>F2Q0EdT:GYHZ&>MP4
0)<^Z^;/)OaT]ADD+d]4M[0FW8HYOC1KH][b78GAAec9&DV3_.>&M0U<<400L<@L
IIf5WFI[V.D2VJJ@GSW]OM_^C(Ve=_ELHBNGc=BWH:79Bc:b6P-dfA5e_+?^3W.M
49YTTN4ZE@16DX/,N9\CDK=8XAe,A@U?DY1KBLgG^Td6-e:#509#Z#.F^gOH#[7R
g2V2QQSOD]c:P/1G5W9R[CK#ZUW?aP?Q\6_/AAI@4;Y5(W0A>?^@[^9R9K6EAZA.
WP6V]]4^IaUM=T.VGgR(5,\9\3RZSQ22I8g2HR>DF+XDFN_8\7ad-,Y1[[R6MX+(
3HNVfCM3.MP.OZH4GZXQO5+;\3=IYIa-M.V@MYBGW]3[?I0<BXB,DO\+]4>.+PQX
>?:2&FUCE;YE1?J,^_-L=)Fed0(HDCL76MaG9f[2&9Q_1_A(DK(/]Y5TKf[FPA,X
7+AX\Lf,(5=5/0W>F+S=E,I>gJaDI_H#g)P0MV37I=39V;Z[GD,R\6#MUR71RK:0
VC&2T7Q1RdPBX:@NJaQ/2)G#]?&gg7:^UX.AP&C6>7LIgB4NZOK>W^2UKXee<^9b
d37CUM>JC+(TEO.0[AZMVD_aLC02H9]-DeUMDX=M4+Sb0,L1aNbb;.DLSgR3R>_E
^3(O+Ma-7XPXF<C:1.#NEG?@HNU07ZQ-Se:ba9P[E9@cR?E,15N7(@AWEM?#:4A[
5KQR:.DEP-V5Da?\PMN4+)#56^,MSF5RH0G[C<4#@@+b2+;9)>WJ5/1L9;W4dc4b
ZNHK-aX&MVW@BBC_RTJaPZ,R<09-Lb\U_ZGAfI>1R7Y^_Y?OaGbFYa7?Ug3?>9K0
,KSMd>,.JST;&HAZ4=F39gCT&c8\&>9-TbVY\<g4@=KY/+O/M4Y7=W/,9O&3;O#3
@1J;?KX]1;=^0T703=Ne,32J1b>CSUSJdI(I(SBZ^NG[S#_GV7WbJ0IO-D/QAS85
d#S8JBG8XcC6a82JC:[J,8461JL\X5#=)2^C4&GIb?,d11SC<N+&bcDWF0AX4;SM
S#K23F/90M-=Ecg,aL=EEgO6S<KF6VPS7N79./I1C((5^534T_(^1.\acP7M<UZ>
;I)HLaQ(5:IN)9Zdf^09^+QL1FJ.601Kg0+QH6G67,=G_KI@<(J&D_.\WS\DP;46
KQM4a&Y\T#V\S1[VGCG/e5+M1;TXN]M5Y0_d,9S@6>1:O&UE_&U=HC\Q4ga8C4b/
KY@NXZLV6EYSJ+3YfD,HP33W:?A1>^.DLb^I^>OY7_]g;d/:C35,V-V(AS&KK7MB
]R@^\dHU>.f@>LE)N2,a63Q([c,-WTPYV6[@(6NPOUZ;U</MFD/F)B6e23^]?.QX
8GC37Kc@<\4YB5QD>@HHcg05INC]PH<&U&NeC&c=6e5Lf0C^XAO7,d+L?#.Z&V,W
:,MBU,aBe?26D86SdWO324DGWc)=FH[,-4dJ1Y:+C]McT3CD\54]_\JfOQ^@Q1U&
W4d&\1:R(:XADaf^]BJP;^D-a8a=cRHa=1:NgcRS^D8<,@-=3f^8J#:@/eQ10N[U
B9GX@O6D_D4Xa;/EW52LfIg7-3)T+N<7Q6C6V,LH_+a-0[Nc2E^\Df-J\L.7+M7#
LK?4UXX3HHVKb/DTOGXMY;c1#E7FSg=7RF(:ff7Ffg7A7+9Z^P6]Z.;e\T4B-YR9
F721L9BA#gV.U=Fb7E6K9WW&:.3;Bg+&af5<9EGFN:P&.d]4OPQ8LT4bPe+_;cXJ
YYT(DY^U)F[L0H9W/UXd9YGC?]WE:A](7)79N7@A)-CF<5.c;S[I-83=.<QWPIJL
JS0=T>&fU4<]3f[BB;48_AOT.G@185N]78f^>^eCH)f._a8(36Y#&[JTa\:c82B=
Bg(B6)_I#+N=P]<[J)\d+\;g<0+3+W\I[8_a,L<QJ^TT@e4W_6G:H-LM@ZcJg_f>
31[gYS]&:F,H&S^O?R/_0@Y03SMgAHNPd3;,S=Q(a#_(CH1+.R#0UKAC9GbKg=&.
Nf6[CEcH7RR4,(X-^ZQA,TJ(e5b1UMDf?]cW^X^K(^[ASe#FJ&\VUKMH/LdK;QZQ
GOO9=:/WW-(fM&C(]aEL,Z-&<QY48J1E.\.HJbZ3W:/ebf8E&>_Bgc@NJ0F[KA\>
?Z.)V=MfDf77^>Z5,MFN\/W6NWU[X5d#gUP=\1TLU3/gN7dO_IXQc1Pe]CTVAY;g
[T&+aTMdN@TJJ03F9,P0+b3^YTReK^3[]_>F_gYaUN4f:_B\QL=ZC[[YaSG)ZC=0
R,]EX93B2,^VSd6Q.[)e>ZU>4KEFL[#\>8<7G((F@K.\SKNe_/ZMYU&2W8>K.+P_
eCK(+Q]HJA6P:?CY>?(A-I42acC<NWKXe^3_<GN)<f@NX0+Da]PN/?Q]SHKIU^6^
a4;1;FAfI=IfW]SfF&2LI@Z_L7.N?c:bZJL6F.e?1FcQ)P=3?XJFUS(5gNTFc0V@
a9gP]SUAK.0=@/LgRg+^C&KG0=F3)IA<eIRVe\?b#_4E;>9IQBXCDd6X8)]SP-?X
UEW0AeK,-K#aBg@A)#6g[GE<=b_EcWf(I@;B\O#1^&0g3LW92<ZbGPS<G\XC0EOV
gMI4<[_J]@fTU2SZ,/Q_KWf>f9_)1Z?:B<7UP85&L@^0gPW7d&2<<D=@^Ib<A?O/
GP@c&aJ2:>4d=IQJ))FIA?2Ke(;\[B.HUNX.ef9If^3W==QQ#YC]<YQ6g:>7)2B1
+.O/@#<5_3@Fdd-fKb&1@62KHWBg.XRA1A_NBZFOQYQ06MDf1#@:Y8J&D6(R:egK
>E?O^&4:e623(IRN2TZf;5Cb,_=4]2ZV5-T]<#T.8#e?N:CcEUW+LS6a-,>7]U94
Z2X5-EQaA915fg#@dDC(&JZ>S&O7;8O[8Sf(PfL.^Q/R[/a^=a(7<CdfA)&dJfM0
6(@4Y_?H6KRVe@/3AX7CALX,[^+Z+97/DbFH@M-7Ff=KCfSg@0W2.2_N(198&A1]
_+dYO9X88[Z1gH0^_AA+DOZ-Ab?fbZ1N?[g-_^]7._;2X#67KTU]]G9F@1ADHOB1
3EIbVCXY-90^VVF.L_L]aJDK5^>0:=B4d5G.?7@-DFF,bOY=GaaCXVB,FB6RO]=B
[E/VT6EQI,]]T^b#E9LLB5OSJ_ZW6S3:,8IG<61H5(6JD.1\GOGK3-Ugg2\4;9E-
F-,S?MHT8PG96?J3NAY4UYML=CZDK(8aC9gVPNcf?YDE.<K&JCI/JM0;&G/E354^
U&Q-9U4WIcL@<C@_I:D.ed=(L;;/b&F40R:MOG2f@:E30.S.Kgg1ZNAaOWX@(AIV
:C9\CObTa(E0:B-eU;KJ5?g@8#(LO(A;d4PeHW/Q7KW&&Hd(K:HVcPc,[L1Df3ZT
90.Z<S2RZTL:>GEV]bb2V&-+2fQ(a3K?I?dV;X#f1,;IMbbL@R?@dP.7:Z9(@O3O
AFGc#,CBX-V<(COI246KTBRM\De89>X^fKI(H,9M8\G^0YIOY/F3<dTJBNGEQEG_
;\&9HJ\CaPDdJ-IQLA5Y+C-@G(^8R5[/\RZF=WR(9J#aS&bKY0f@\0F8C7IGDIF5
],S)Mc>(3Y=DQS>egA&5Y=WDUBOG4/D,cdTBA;aOG=8X/1bAMWGG6<3W37L;fB]T
)ETFS)>P^:g71e9e6+.43OO2&&Y2^.Q6Q-U,PSBD;(&E,TL3>GKA=X^)>&2H.M<Y
5I2XM#7\GbI)64aI[2AUcIdE.UL2HCBD4g;VW\cRDUBPC+L,BO=650U3)45+A3BC
4A<dfPa,#]4bU3d31O@\RW,,>E3Mb5+CgXf0<UF9_ZNG(B^e&4KQG3O#eZV5WD>5
(F5c?1R>I\0W\g_eSe8a>XSTSWb+88Q)/@^IcZBe76W]]=CbL;f^Jcg54Ad)F@<f
Y3G:Y#UZ2d_#aY9HZQTeSXXB8>E-8&T4,FQL]Q1>e#dL32J,cQJ(CLK4-(]?,:Bc
MQ(1D]J:G5.@W_7X(1FSa:M47O/7A?^44/)A4V[f;Eg2KH.aT23Ec^IMDDQP@>YQ
12D@fSP34)XeO^[a40DP?#S?,>3NDBQ..LOOF+3M74]9Tgaa,D/QB1CB.X@_0#@[
CX-a;FO2J0T#&McS^,5R@<caJdB9N3;[G\(R8Re6.9e<##gYH&G@(T<)I0VLW+C9
2+99,<^6XO7g)\b[_]GTTL@McFPPFF.4/8TX7ceGZ-(1WA9N<2D(b^[_LVK4U?44
_VYdb,F^7F8Ya\YAF6d/;1YcUUC[9)f2VQ\XM-B_O^Q6?aeT_-f/U#\PODc(1OCF
1<N\>WT)Aa[LcLOM0[O4^J[-.3-C6./gfR3:Db\2]_J,g40-^LI\J)cGeObV9UV)
7[6QJ4O.QK_dVYO?MOI1]_744d7O?KQ<)>FJBNI#bg:O?.(QB?L6Q0/PSe=JdAJ=
e6Cb3VbJK2dK=C3LS.]?.Z=CU>7:?ITG@NC8ZE(HDM3]HI_Q:F1K;_+4_5_3?U:]
9I0U+MECU6M=GL.KcfP\W@@^[?1aHM/12[=d?+?0PU&@(98Db,+U>U7AaT/>MJO7
R;cW#VJI2\7Bc#.W#cbeC:):[[ZW)E2W&;N-gB</bSJBa;]+748CY,NJ\>=6W9)G
XOa&=0-&0(gG_d-b=/KP(HRO00,KaIbM.C9?1gGAVTXP</36AHD)]92@W[b0I./5
Gd3KMNA?O58I.LRUXNLIO8b)S\G.&3)\Y/c/S+db)VGBUGEC425Cc7&,]RQQ0-MM
_f;#XVO<KR,KQ<(cD0e[\1f12gNVH.2O2&W36d_7Q:1R;\=SW0DN(7Aa,5)#A1.L
;(&S#(D?P77L(_2DPP)&X26O36J,F6D1)VIaS[OD_\8AIVTFS<3MR_H_IM\Y>:9W
aZH)aaJ95@^.IWEQ5(0L;eY-1cec.[D(W+6\Z^6+#7478_/6W5@7>@cNC)@BaIKY
g=AWJZfM;>68]38fUg&#.9]Pb&>W&NUTPZ@788=P6]M<D/8IXbO#Wce(85ET=L,3
1ZTRYKPOQ[F69ED-E>0aOB=EJfC#&^<dC(><.ag]<8HcG,b>L5:/_@7_MW&>a8-<
FE>DH7)__SOM8Icb]<PW11OX@)_V@;\R1;YP:.IX9+SeDGOTBP+<]E]<NG/[KXeG
POD,5a1d>_O]I_?;2X(I0^[9ALcT+S,D2cYSAPf-;:/FRL7;7SGKABR3Ng4YVZ#Y
8]JF1FeU2A(Q-VNP?#F/)(U>-be#=()4:9d<E.d>=]4_McR[FbKKV::=&/[-bfWc
FEB.8(Te).?4B(P0JI;.\29b=AbT]<W,_(-6E]L,G(>X6N]&3g6[]#YIO#,S(KRN
HGJG8I7JcWb(G]ge3SY7T[1aDLZUf.>e8\0e2<KZ7QRI:g;QTC)8I;C9^Gg++\B;
6e9ZW#U]<[e+[)g&4M^_?cRBGeMH:b)(Bg=>I;Z(:,Dc]</?S#,^e[KG7QWLLKHZ
HgTH;=eN4Wc+2Hb#TCe@S6448_Y=##)d0GdaAgX35C,Z#SHIMNbK[aE-V2U>8)_U
@3C7fV_eI;3GgEG_dWE/LB=2RYW&YA19>5f0\@#0(4V>26X1=<M<,\U[Vb,G^3_Q
MM?J_#+3ZVRS,[R-gGX6.gKa1>HJK:Ne<\3^(+5ZC>#>1:8+.;EXB_AC<dR<f]Yg
7E>=VAM0d<KZWOTRcMAI_12gE5T:d6T#bS42Z[e_F(S?\U5L25;V+(YTWZ^P;X[J
2/NC.b]G>:.KC))(E8ZB\6@H;?^aV75Y8D(8AXVP/CEf^H1CF#J-GW#bbAff]R:f
+[]bA;?<<<=g;P=I2SLLNf4.b5fCXS;F/U/XY#QBJ/]Ha2@]cVc@:RC7D-K#gMMX
FW1Z]9..bdR7AH^QX4I2D2Y&Sde_2GAD^9:LXc3gW#=W00f>\58LM\UY:gQJ)\#0
YfIZMNg^CW_/DVXTa5KHAU\O>+:ICD((=@VM_P7BUbWT3938IVWFHaC52V63-T^9
a)XMf.89ZUURNXVFN<X.U#:]U<5LHOKI2?1UBITQTA2YSAQU3GRH_M+I^gOg1>5#
.52,>1#WMX+<))3M.E&J\D+(9:U^5aND85#QcSNCHK<JI+KUVZ2ZNVZ<>?Sf9a_-
fe:=N-D4XG9+VI;L+>FEe[9BU&<3R8L9<eR0LFAc)P8L\IU6OdFM5PEIA4(=&0]U
CG<@SYDUN69+>/_38_UCd?+LFB1YdM;BY7g7c2f#-.CUU^N;LB5?aAW_A_68G:3V
7DOCe0bQ.1\@@/+0SKCBW7<0<aZBU@,CR_K>Q?PM8ON@I=F]f>1]e[?c[PUCE6a:
DbN>52bW1Z>(;]]&06g3@b4W^[WA=D2[Q;7^^d3TaBJ6]M8bf-fGI7GYUN9dZ4=,
K9^(BM@1FN22f]M/)/b+XX):S_QF[K53Q6d_fHd0,[N)Va/bU[#T&7+G&eaf-fg4
ODA&G7KECVHg-)Rb;H;,7RQ-c0^J:PaBOILCQ9)OMc1=LB>6QDIW757?_9TY?dW7
\/PTGGeE>83JB;4IH3ZZ6(?#JT.f)U@8g3I6LWBYH\6LHGeD[JO+(QfLV/\D2Gd_
beSVf)MdM.;E41.ALVS5GcQVK4A^S---:TJ65DU#GIU-/<FgT.RaE1U6eYPNZ@dc
KWBIaXea<ZCW9A#C.fXFYH-#[a&_,>O@??>.fcg33N6&6[N7LV6,DUPW&@KaSW-)
ZV<JdG_OJC_J-54F.ERMSIa)]@,1e2S=>K^0NORaU3AO_Hb>TECRFX[5TS5(3+=R
bOBO:W+HEY>QLHVCYSfMNW;:7a)JZgNe=XV&dZ5[J695&S6VL<ePf7P@6\<>V<Z-
RA.EB:F-3PE.SA;T&DE?]1LRCEFO0@B9SXf^ZDM?K\4VD\/5RJ3=(^GBIZME3\6(
g(7.1^[c?:]#VZRDM6XHP-CdRW7MA(2-17@Z,B&WIXMXe^Y<9_c0.4(c\91,B2a7
;K5FQ2QQ,HPKQXZ??JgQ_+H)XO)S#&,D<1f&V4_)-,B)d\N2?@f?\NaZ=76QD+9?
fR1#2RLRF;E2NYd3)KIY>#FE0XX94_>d##?K)Z2BG838TM]Hf&2AG.=eEH,FYcK<
KY5U3JV/=/]NC2<ag_R2@@be0BG>0Y\C;eg)H>53cU&#2-XHe:QH4?Y]4;>R:NcV
/F_,)7NAbI6a4TIdIIN:ZSeU^Y6>cZ#Nc7UV.\@-<F^Z\g4FUbF6fEEYgA6YJIFf
L61YTI]R8(QR>&=AaXKgR-<=Yf<DYC9b6=c#=g6+Ef9-O95@E0b_&e>J<70\H-<E
;f:YHZgbAW,)XccEL>:1bbGf3PTJ[;C?g5V5Z7Q.f5I)[=f9+;^Ub,VZ:/,(ZRLF
T(/;^#TH2WAgI+=ggaQI\ZZI71;=YI<0.,A:H.3+WMA7FaO\]83PJ<B/TJ2(#^4Y
L^YYZNddZ;V_H1>3<d77H9+(GNFY0bI0\b_1BRV:W,dO0DNITT\Z]XZgbOBDUf7E
#2ELOJc0)B8NEEN/O:#H8IT7(@C9@621FUHbe&04QTN[3TH3f;WOM6H1Q[aDO6>3
bZCdfIY<-_cN-Q0J6TVO](:Y/>Z1/-#9)F,T9.L=J&5QB0@B8OGAD1^9<TWT<:Nf
2ddV?,KS@aX-#.T&^?A7I;N?<dMW/4bLRWbRYdS^_3YUN@.a&2[4P0a<9XQ5NL?W
J-S.LM@a-DV_ZT48@MA2gdQ@WKXXK40d715JLUAM^=&/N/9bK\88#b>f>+TEe]93
Uc-AMT=HURG.F.=UgX9(-fg<7(>IU43eDaL1\.O^Cf1.:(Fd,9b\#)F7L7@c6/R2
RN=/O6&Y7L:_NcJOg6H][8++1_AQB,.:^6HJXKeW_LS0Y(@5V>OU-WN6TPE05E:(
c9Mg-UH96d^BX7Y<]RP2\8J](^UZ7PcTe=;gD(FO5cIFf:_X58+0US7R<;O8(=J2
[+J8PNCb(TO_A>>d2T(A<FJa(da@e_X_NIX^T;DaBYL_;8GY7N/-I=Y=b#NK^a9e
8S<;<fZ&fg.gJ]\XCIBO\4/R9S4<\AGOI?#AQZYJ(P9M._AUA741T;9<7_I5)gDe
Df8<YSO^MO2bX4-fZA68eY#3cU.KAV#DXY-&>):0f&PeOC.1HVYH-2H,cHS9#Y_3
YT3bSQA5#)J#^/A]X.#6A(U>Z6C.0:I@TFe3&G6_M@\4+8L7E5dX3gBR+OEbMZV2
_eRTc?<5AVJP#TUOLSSWRdMOJIbPYKX\B<G38^J/C75=:6=a>UKH0D7;P]_gN2A,
?O8G^e+B/\_gV,.eIa:F#TCLK(g@[NR7>&@LbC31[FPQKE#DKY,0W,6>E&I]))ET
KS47DCMR9Vf@BEKTad=8K7V_&C3ANdMX:aRT8CEPBPYf^c9XPb;cAaLDSJcILNO[
dIF?8VTgXfIHg?XP=NJD:5\M#.5aL.\.(P^?2UWYb-2XLX)=TB:<U<NZA4]-)>fB
Df\1;AH]((g?1]H<QN?WEIO=U(H_6JIcaGM6BYF(dF4]Y[53304KKUJ7@:I#PNgO
dT;eZSI=Ic>+IZ,I4MKGQ44:D_g(c\>-/4(#).?TQQBbbVb-&XA/])e3,-IFPE;F
1Y06bUUdQ7WAd</4&=92-XN]15YE^5:bCT@&9CH#PX3D<U6MVDg8A8VGOO,Q-MD>
TS94UE/7Z\bH;^-3K6Q5D9;K6T4d9d9U+YC-#&c9870We-A72R6K5XC-Ne(3+^VC
gZbf1U>CeF8eb4dd^L+2G8@2)<4?&K=S>TNZf(]:W(^W315IbOG8B:WU3IUdXSUc
:O4d8Od0V)ZAbc/)^_dIJ]ge>c5D;OTWb(R;09\)g[DR01)I4R3=<<DGfU<9PPMF
cb&W;b88CVEYFZ)bQF-3?0XMfR[(<XHLNRGFG[-<4@f)c@KeGCV4\>b&0U<G^VG-
T^>2TO]6bbKRTW4:Tb/.]:LX8JYZB1,=]OG1:(5]^ZPNJPb5Q&f4VPaKEY5\d(SO
^^]S]9T>?0<X].[BIPH7P1gE]AG]gg7AO,_b5M.<.ff@J6)_Z0AbfK^I3;AQT^_W
NY>fAAH:_RGFcgC/2#E9<J5b=5C=E_W78gL\F.Xb-F@-;]\INJ(0NP23_[>CDXU:
#\1<0fJ)0]T:gNeCf6SN4MRP@XfIB6.b.gJ7QT98aX?:7c[SVBR+1O;<W4.A<\U,
&f:4#]AOF8GDB5I3;RRS:I\<[NU[0Dg[F\7PZe>H]WdXKY-/&<JU_OAX2fVd<Ke.
MJ5W=[J>7D#MM[Tb?b_UZN>?)KV?^&cQF3aBHTCV0a<L+3d8//[Pd(D_JIP+DM>4
3GB8?TR\8)</27.bb3F-b?]3P0bF.#5GU\L9ad04>J7faDG+=V3O15YTEgOZeN=@
(bXf7b5ZeP95cKdY.7>S/9f.=g65+]6BFG5Y=fgO#I_DP0=/L125:4M__(SFN3.;
.</U:>F-T:TM[VNZ\^fM)Q7FAXESgHdF;UY)gcDK@?<)0<N\UL,I?/.>9BJA,a\1
?K>:bBQ9^b<;.Y#SZXP,&#7AHB.9QA:\CYU+9,@Ca6T;Nee\e7MeY8;4<^4Ad7V2
)RCUZ2:,K1.QSbPCKN\Uc.^R^fB?4-]]7JQM[&YTd3HeFSZ4B39MU[<OXNQ[ION]
X)2#Yd??FBSa>;2/B\H(MASPYM2F-)#;=VQ-[M2e_V9X+C>3f0SYJDI_209#Vg+R
UE+?KY<CCUI8M#)IN2Dc3aR2N0TVg&99^.)TKEc;H.&KaRL,WS9;S48YRXNPdgTN
6&YMeRCIV#SXFefP7GcVT-SBB]T.E-#SW9+UD6?J:J/[RDQA\)F(7IOS0WU\^,WC
@+5B3])34NV:g.2642+#2#5YUA>-(_^@WA9_Y-D/@\EgU7aC&SgKI#@\)>ZG3Pc?
V@96,P.8Yc[gGQ6(#P]L#?8/[B^BJKFV957M<Q)^RIA<JBe1F8;+0I1;E-6LH6A1
KD11/M5SX).PV/4PS6JW2E<gFf7NKH3]ebg5^7L<PT-F.>ffHFGa>\2^PLK64@SZ
,Qcb)&V3V6\D>6g-BN;[>^#0+eS[aF8_^+73-L_EMEXeeOe//R;R0Q<2P/90[-Nb
K4,)Q88Q(=34+&TB?5@=IL8XDJ>6IR9@?2_&7g:T)9+_G_-MTZZV7^#AYZ6)Y-L(
F(K=K69a2Z5WWCD(dG9&b;\5fA=+W,RM4f:,#ZP-D&CCJ^9<=;(#,bHQ3.(J)]FU
KRHX4@5_LT7IFeCZSJ4O4G?(_:cBW)WeFSLW9I[=HNd95K6;U+9N74+,^[KGCefI
9Tg@S2V@2e/RACA]-X,\EfIW04#&5^/I-B2A>6CH#,GUB#JU[?ZM9G9NEVKb-0CE
<P\Z]]2]<6[>Bg]f#]/PJ<2X6?a.IH1bKAVCXBc)D4dN;.YC?RT<aQg_)_.@#)_g
a[1LO?WS8HP=bM^;?A6S48\W,Z0GEL_a8D^YLNb;^A2d3-?D9c3CA,H@R_R[U?ES
Y,gKGae+18?Z>8,SgdW)DJ2Q)g6LBW3X&RZYFD82>G)2,fBTE?W5JG/]XVE<MRYg
&]8b66.)##;82KC/L&Z?#PD648?:(G[@.3d60W>.(-.YUPDCH2CDB9=K?1:]7fME
H^Y<)0,gU.>:;gQ+5FgSf-cgXH8H/I0G[bI^0f]GL7/B(..+8?f?U/cT(<+D;c#X
A6#3g8XAWO4=AB9^#U/D1JNC^)a#LL^gF&#4eJLY:\]<N6LQd]gA33Z,c:L5VM+f
8O\(1VYbC;AR8^e,;e-;&4g[IeJ4fb-&J;T^;=dIT&RdX)4J.COZ8#&5Qed92g?2
;Q6JW_@/84-]Le,-;CPaXg3/GDM:fD^T+aAPI/<S^\ZISMW69NM4b\Ad4;3/Y;&f
3:F<[Z6]#a97T6PVbY,/5M0(56g07?J9U]QBS1ae41[c9Oe,V>&P+=Y<492)_.a#
[6R-8=2[+X<eS,A1&5YG5/_&8W1N,DX.,KaU&dP8U/Bb=(aeLP>Lc._g^7EMQ)eP
W2:eNY^8,.C+(,NYJGHCWRd[0=[:T)aC;D@ISe#YSd]>4Ta)/(.-839g/=N+W/6c
96(_DI4TWNG]74/.>0f_K,_;(D7/6cO^E:1([QN9D5+72?+MVNLfPNW+9HcIYA;>
<-aCfA@#eY#XSY_;I1VXT6=R-Q[XXY)f?Wf7D\D8^PW9QTg.]U.d(\&YeD+Ed]Z)
7V+R>B8L,E@2]IU)FYbD[M,=dJbIFKSW8cZU;)YP43.&]gfB3\0#88+,O6XQP^4E
S.(+EPCL<Ed7_I4.-/+M2?/cU&3@Ue74#N:QJF#_NAa;#S=D+K(W5LEL#EWgREdB
/FX2JcQF/QB3#_a^-/23D0IVXV0=R.9/VLA61DL6-EJQ1<EJ-)=-8]g7UMg^CT?6
W4Qa-05N4PbJ:(^U>S,O?^YK6D:>g-4TDI\)8B@d/GV/_0^F@.c[F^[2b;#J[cXB
[F(ZT&3d4BAG#c^4ME23/#+E,:Y+WPRWe7.6GFXW=,#?5geZN/?66\BL#H0f+Td4
-bGJ-K33gKcK7=f5+Q@)/?-U>?Q,EABJE:;/F=E&()AeQ#FRdY&U].ZdXC;\-GP>
7BVNc\9HPAgYZD&C.+UbA@2T/QXgN(1<^MEf,4,PJ]f^@RdV2;WgLDE>_[(L2U6]
+Ve]DHR8Rb?:fU?E[H9Z5W[I0W?NXB@?KC<-Tg).eQ5b@-[.5S6=M7O[.@BRD\Wa
4ZUgOc<\0aN0=?[<7=f13V\a@gU/J_&cRSZ:aJ-Ga,YeC>@JEQ.Be?(#.M0M72+4
?6T^[&LF,?fJ(=@WX94.=^c>#10T02N6E,T7<+DeBO2Q1OP&0d1\fCb/YV-E/)YW
=)>3=G>TR(<0)O(/M48.Z+MOY<.(27PB92/@Q[ac8S7(,LIdg@1efW:\CSdGfSZ1
/\SMYDK[bK:/5#4J-OI,50HZ7]Y1ZZ8_gZYb(8R6-/9[_g\-bI=-).bbMX8e:&;F
7@a8]e@UIUCB&f,7X3^I.<aQQJ?\W>W^+1ca7=EBYe[eJD\&7:<[)a/@[dEMG7\Y
\#S,9M;=S1+G3U0,C6FQgb2?5?Ug&9W9/1&\Kd4fV^-S?>4+XdYKY_Y?LSRXMQcO
+G/6O<fPU)AcV._0?(5&[N(4CI+LG<aYg<[[2\Y<f)XOB_eR9TVJ.@#Wa4JV8RQZ
DcP\4SJ>3XSDRac5Rc0/P\U3_I&FW:8&#TWJDC+N&\4;ZF/UZTX7JFVbD.Xa9EVN
S&8:US+9@Q#PS<D8SYAED,,TCGSa;<c[YbH:+05<Xc)P_05&&gG-b]+>I&V>C&[b
_C^1PK.-1F>8NBe6?YN=bb76IcRILd;,\JR0SC:dPADSZJKHf54Q]b]P1JDgYL[:
A;G9Y0&f+a_4P9))D7DYTdPY_^T0<U^JIZbG(7O95&20OO7?8R9IH[AGIUM+58Gf
-2JS0a^O5WAO,UILG)S6]\+\6N>;AA4b^,SJ+b2[P?RITeV)[3Q?SX&ac&3TCOXJ
>8cEKO_4+MG12Cg@F7G?aVCML/P^1f5C>NbA3:19eEW>&BVB]Wg/?bX&?FdKI-@/
-OUE3/824><I>6[L/1R#4=?VIQbdR-YZ(;TEO<Z+H&]F]cA0Y28aVUE;K92X\\S1
b8b(CR,G55PN\gG4Gb7..AMTTS;cf-X\EB(V)Yc8Z^QMO4Vef>\5-;3@=;-1<.0c
P]7TBKOfcSeW]<8)gFegPEdda3CKS.R3O=E50[-#2A@]D\3Be,b#e_KVgL?],KH^
N1\#HT/VZ<Teg(.1Z>Z^[?16Ye[bEC40;5aZC88c3</W&-+.E5,cUHAH8f(;eY3@
?B.Dgc8ffP=-=J),=-Z&7fbZ16B#9IU3_Q(G_Q#N?_J7eD)>3gY,Od.-_N^99:EC
@6g+e2\N@Z6Z+A_d+[f,#;d/,cO6ba?MUE32DL;G@(&fF9ZSTS@c.IK2GW9M4UFB
((I1CdZA4Y4X]0M;^)\KX)@8#Tg4g0g1g,dE2;+bNB,;\8>ceEDY04D;C7\2+/S7
RCJU\^?P3@SFXf4<#8\G@-c^;;7fVL];?4cPKO+[5;Zb1gY4[)3NU@IE5L@H222a
AXbdS=#.,,R6H#E+QdOLJOB>f4dN=LQS5>>MF;Vg<:C4(<BfC\bBA66S3f:@KJ+e
:+N^G;7NQ=If[@0Sa?#L\a.P]^0Ug.I[(VOT^GDOTDK4?eKUcG?(]T<4N7[OM8]e
:0012B^Ug-M(W5E.8AC8=HbXK]1HP8EO>U5)GP]2)SY>edHB.F@8??gH/KYUJLdR
)9cF&M]I&\UKc(@1\IW[WJ8PU][-X/5eMcb_I?TW<NeO&U7L44FBEK=0(WB.S]>O
YQJ0a-:2SYS.b?N?eb(9^;LVPfM1YL6(&[((aJT(-UBHHdgg?S5Nf?8=DY)N<[-O
?I+#=H#21-?_14bTVH);QW2.=_(QNMDQ[=.XLI@G-K;=[D_BZ>Y+K^ATR@5S#0<[
<+M(.AU=c5=@Y4IXMOg6fG=/-ReS.QTgSE:IPG?))gV>0AW0:PB6_P+/8J[CURA5
#@2?[&fVW.^PUA56G#5)R^DGg-T7eFUb)[6I.NET90#74gYR,-?6f8NS[2GcO\=[
G/(_Q2gP0/]b1b^Y95:_gRb);Ud5@QWK7/c/-/118C3;[K5d:]G+&_^gSA-7QPV/
_f@,X]EaXW9=:?_&:A0=B,OZ#.]#\2-X]-AP@O+fR5NFN0[PHaKC#IH8ULIG\4cH
B?L:.[\7<G_2R<Xd8@OI863<TENRg\AB8>RP]A^eA4H20\&G6TIV_eKSG>06NeGe
G)e0;gJO(T#SH2>[R2N4.ZZ8N?ef<3/2#DD_;8Q2SF^,&)CG_9.\7B5UKHOXef)W
,a<d)>LR)#UIggGRgeRPCTcb<1+[c\a(b[N&)+Y;)6TB7_S,g3TQ7LgFA2F\Q4JK
CHKg0KH\XK)O?#g2KAXZ],0)gLWT-G:I8+X[:<14?2,7;=+HNZ@3)VCNBEA;a1)H
;8g=4A&^B:,>=?:TK/2+(Z?+;a-2X;UbfVP:CHU9G&=G12<0W>H&.-^_:b/3\7[a
?#2C/.@)0E@C3g/QQ\2=cYR?F]0QgDAacK<DLH8^&6Q[.CJ5M_RV&PV_2RG2GgSf
)B#6<K=1M\K))M+Re.1ZC2\-O64AVM7<2C768e4)B#2b,LTa95b^KXf,-,J5c3Ha
\U:4BSR)6@AeJe<.&f<AO:]:#4T4c#JOR:&,192f&WCc[7.Jf\BQRAB?U=@[NOZR
Q3EOP]UL<AfDJC4K&<6UT;U:#G,7.C1-?E)d?&IaEEP/]R^gI1WW\5Wb0TFV&@KF
<G7a\@\FGR-M)@L(-,0J>D7II0\?/Y6f3AcQ=#=27SI=.R<fH\D^c<cEGEY6C#,K
MK(X;U&]:IUeNaLH@Q4YJ.[6259=E:;G;5#BLMb4\U&&b?;ECKYPH@W;KG;?&.GZ
Q.I5d#&;UB-[DL_VV9,UY&2a8X_#cf^J0>A[(\>d>Db=N+A#W2L4-A)^&Pb_L,8M
,7E,P\,<HYZI;CKVD6fR\W-#@NO><f0/:K=eAL-QaLY:7P.9/M11S84+-B<2I[GL
(M,Va<S3QabRT=AF,PE<?R9PU+LJXgSCF?_8MF34Z[J@DLO9-4PYHebUDWXCZZ_#
=4PVcW+@9c1-;-;-QR9=6VF[[2+K(G+Sbc?cRO,5R)P@XR5K.f[LT.#eA(&dO2#W
L/CM7-M[8daL\R-f)@<+):Na\6=W8K[#L1=QcdD])LXMgC?ROg/bBb)TE^40c#EN
UB9G#TG950c]\g&cWBQN4BZX&6\c;);77-OBW,^)Teb(<fWSC#BIb7W;^JYF0C=-
TI-^(aM,3g.5BL&_NT-T(.982V+e^)4BDC@YBA;g78U_a_KQ4T@[L]4G?Y4J88e\
[=0RY6d?^I-,G,S9:M^(Ve0>Z4C/E<9WKUe2R4@O,Q?D<0/N;JFY)I?K:@KT3H@_
.8JM<f=D=XdGWP.M[I(O2[U\SITa,,aLBEM0SUJK)]JJDDPa=VPcV\RGg>fLEF@G
\7CLb\W^c&4J64/1a.[,C]c59;J+M\CXD?UT8e^P<dL9N]NK:?[.5JQ.>/DB6=B)
WF>H+bfA3aG[J5=TOd&d0O\/_4bPFYbMZK#(F871GQUSg\SKX;^QdaPg_B7^cc2&
JF+E:AB4:af2c_126V;bO))KEB#0UV/>A5<:+88#FNFT]^]\JT61gcO]LaYU#.dN
7..J;MXM[,OA_-f2MPPJ_YIAO6g074+,+G](e9[C?[3Ve@4PCDgN,^g5OVA&D2ZU
cA2?^aR\D^,@,aN5Pdc0R/?&56+7>R[66#&H6HWg,Xc9d2LPH48-g/A8D4_;aKH_
Y?Sf_9V.P@9XWEUCC(e95abIO:D)#9YWO.-0:?g+_I9YX5(AI)SY@D87E/S&40Ud
=FU+V2+^Z7(&YD?[OE_\MWcZ5[4151fdL57a1L]:4\de,:eIeY)A=J_WcU8+I[((
H;.=@/I?U#06ZVQXCGbSTHA\\E[#;3:HJ@Ke0gd+1>H8fB+1MJZSE\-M55(3@D=W
OE,[-]JALFI-[RRV-b/K9X]&HdAeP,-P^TF?VP]9#N)G<22>^=NC,ZgaQdNOcY4e
#BHcFd(4aB#5ZUBNJ:5MBCXO(4:C@<XC2Q@>,[7Vbc<,WGD,A)JYGPUYG4M[N.0)
6=HefEJ+L&7/bW(Q_cdba65cFLD@?TbRZXRdW/IJC-V?:/d)?8W+@?a@2gQV621K
A6O[7+X.b13ePdS;1\>(F=,:@_[I(eS)aDa;H[#8T8WLT[X494KC6:\:23a./FL@
J=A4cGc4GGEDNeYJ?.>>c8dV;Sd=bG8RZNa>LUHgOg&#SNNA^?cA8PE^+/[f\1#_
a3Q.b70fMK3F?Z4U.fM(&K1T_\:D2?\0Pg&b^3:MB9)C7I@d4ER^\J<9Rd>8+LaU
.6R\0]+0#431<P-MF]>>:BL/D/f9JbeN]e73M=3J-gR4PZC4G_N?MI8SfS78/M>W
(C][<P824AG]Td\F045?>5<F\(MVNfe1Y(.NBL;;PR/1Kb+@[=7YQ-F?_J0f1#fY
F#Ra&VgTVE^WcK;3d^?Y\Ce=R[d2^.[+>DQ>,TMbEWMN?W,0(U^7O4SLVY0WGFXE
9-7b?RHXW#GHCU=0RSVPCUAa)KS2+g5._&QT+9gH5TK>+2ZS-HWHDU_)<YNLOJWG
>.5AR:G-1->HJ;2+SIC)F.+OKO1H:E&J6V<@Y+I>)WU95DJc;;Y4VKeW7J05Td,>
B3KdU^L#fH&66.\b/7N&@ec>Z:S]V63C=1I2?F1AT8)@]T;:Z7WGQ1MW\@1N2GWL
MBPA/I@dbbf:+f7B?T0KYC,+>VbA:>Bb3Y9RG68(L56d,M586^3,^ZW=/(fBOD4)
.5]3Nc?2R1U[\-25(0RNRS\?I,LA?BSfW54DEQ(CVfO-fdS3<+aEfYKc1g9KL=fM
Q(]+e2C8(P6IOHR.4#_NCD(Q:T,Yg>P(^8g,H]>&D=5fV_VF1X7D/a1T^L0DS<(g
))D,LML3\IWgUC,B5AL3dN8aaTGcVda668a9;<BIJ;7T\Ac6B(0MYV9bN#^R.9N9
6V#-_1>X2OJ5M4Z\gG)+L+GfcQ7bULHKAHN.[EdLAPX,/YD:#IF6d+BN-N#cK4GT
]T81f:O(K+e+W:R_<W(?SP+?0:]VRAIY9fR,?BU6_=XNf.YfX#>_Y9^:XM]+R23N
&K;^gM#43CMANX9Pe1.&<?M).2a]ZB_CTJ@+WQ,-Q(5C)+,HI7D;^]OIMCU0eTab
];D-=M\2;NC;LD&0Ud5E9H#D<^Y8^V5_@V=P+M;(/V9.SAd;K>cZFP+&Q8aL1LY)
4(,<+e;?:0-a(+N;9@UYF?M?N0[#R/A@)OF\_ROTfM&8(eRW;.?5.>[PM;&EEQF2
0Y43B?R3RQFVCg_K<;NaUNAa3P2JDVZ+RDI/28<^XE<;L<RT-;IR&c^V>C]LE9Te
C2V(+O(LC((G[,7(?7779A?(_P86ZNc_EM0>YFF,E93</IT]D&cJa7+5O?J]X4R@
ME,K=)#[T>N@7YBgA[)VE>\/b69(2)K5d);>YO;9gVW?8T>]e@4@K[9Ya+B3][F[
?=6=Pa[0JR4@R@5I@9#?OGOI2>.WM&BSYCC3@R5Z^+GA0A97+@G_TZX+\3/K8U?J
P:a3f5a,OY5S>6JU0)W<ZY+G(Z@f^9H[=)6]O6-dJ;\0HV[6Fe:3B_Y^c><3_.fA
UZ]J#/QJJA7=UD^=SBN;&Y3#4^6-E(48CT;ELb=Z))9/&,AIWD8f2CLMgT/+/L44
fJ0X<KLLLMa4ceN8[_WNWIKGD-#OKK+5E@&F:O+/M(W1Sda,@Z3EECCKQ]fC4+==
IXb.Z5C#H75@CZ=X@@)JVXe(V4[+aBGf.-I75JV.(^]0U&de>_cgL>\^EMY\B1Q;
eZ]S:=;5b?:#Ua9(C,6H6Y)<@1Z7EeA;>B/6+.4HE[C.I96^M=1U2a[g9>@0B<?b
a8#Mc:_#UTX_SQ-)cUZgfX#RRE70a1JQZVI<^;a?SBfEW?S7Y]XB+6VW9M&[OfV<
gBg8YI.S+R#JNZ0SKA17.#-^VBf</7_V3=M[J7f=5gF.@&.aV_^CQ9N5g,5B.5([
/M5)(=_&CRN,\JXF8[DYg:9WFBH:@=g0e+UBO(#SN@6[[1]_#e#5J4ULE.62@/\D
Xf>\E[/5AdG@=ZSXWeHS43gR=/MUb7)CAF9,G55+^8GD^:<7.^@RL<O-L=MS,Se(
IOGN\4U27^D5A)\WPXR<MeD3+Q^OX=E(;=fQ_D9&8Gb3=0&b8^a04bD4B-07&A<=
/f\0-895NaDW:MJ@MYCUMTY77FeWbFSF@SUQGLSgb_C.f@4>N-ZVaP1X54d=e>E/
=K))eV??DfZ84930@5fWU=PCKf8dcR5SQUed??73T#X#15.;Z;5U;D^O4f0bBac>
]5a_I1XYeOX/=VfK0.WKW7SE_Y-d2F6AW]PK_RJ3S^5G@)KIS&Z&ec#LgW#5YK5+
6E;VT6L02c>c^;&Q-P(N#85d@c(R=&1_]=?13NU>U33>)B/?]:,D-J4-X]U]RgIJ
5c67ZR+]TB5]:,PfQg_5G(&FDA@CSZ6L-7B]CW58X.0C;MX4E:.Oa#J8(44J-E1K
eBEO\X8LUVD3.[3bIL&J/]G2fOW^W49aJ.VIH\fSFW,8&:]S&OKfKga4>]7Q27Y<
E_b4I7_T>d<V(;9L.4/2=c8A.:WT06T&YJIFSQ>SP6/.-X=^E^NKGdPaVLdGUU5A
1SBb\4&5d]bNL9E4@TKFeYL:XQOEX>6e4;(3c\+NN09?(\W)Zf&UERJYC^ROCCea
#G;.H)@A2f)WAJ:(&SRce[PPg3aZBZ>RUe#CN),@#V?-U_W^+e8NGL:KOgfDIBIV
2;g2[:^Yf<\,+.Q_PS^EF\RUT#;7cPAUT/Yd<_f-O[;;1>(/L7NJ+CCaM#g.d[0=
c=\eLK5QPJ]c2Gc^DQ7@4.ZZ.g+U6=@;P=(CbJW3[Y>6[d7OaP-4F7(4#.7F_1/P
SQa<I-/+a5]4)1gJD4W^_W70K7L4F]Q:IX^?7-X.gf<c3VXOT.9fL6?C]N?J:1+@
9#?(:,>Lf6K8Wbg2:Vc;e^RPK_-gVcaTV;Fg[7];7Z/;88e5HN:-=W36H1(3O+#b
6=XN9Le:RM:_Q[HQ[Ke@2.2=bK;>dC.QU=OG3E<GgLEDB7bbXAZddC-U]UUMA-P9
cLef8M4Y?(C8(NJ/2^8:B;7ca2QJO,@<P,WU5TbabCHQ1IXVCFf8_RL3aGVWRCU\
,gU&RD\\W3THVGa_XSY9Q1\C4I(O74f+A(9;FFY?_4K6Cd6N<(dIbeE@=&-@4H]A
COZQHHa54.8D;c5&(&0+7Y0<2=?KFPYIM.79DMK<&MDW1d=_3M.])FAM89gHY>BX
IVa[2V\5ePB1de5G2AFAVZPE2V[:J46J>@?F+QYYN]Pa>:HR_R=Y:?e<TQQ_0_d[
QQ3(?(LOCGED:9B-]KBZ94ESAIRE9<B,GC3XPF?CO&HHBJ7cL<gVeKG52\MTUB\-
+bY#GW?/,7SPBY@aJPYY4d3)57<B;9UDf&Xg,N_>8I]-(MA:.KJ95RCf-@ESa#6I
@Fc^5F678&Q8P>ae]IOD?_LS1ITKR+:Fg1]aDIB(=I,&(6QS.4;c]BDXcUO73&]3
a9Y496XT#6+a1<G;UA6d^>9J[?bf@EU0,f1(fgEeKHf>^7a^5^Of;Q(]JSO(>U6/
V/P,3_/YWJ+<.D9H;Ue0FS\:XDO#JB8MG_9ZKB3O33<KNCR@ESY2;XI_+Z=@[<Rg
/g_Z>(\BY^=Lg?:XI#6OeDZ3,Y.7;,e>ZE44bP:-Lbf-J<a^PX<27g4^M/J:7/H4
;6IG&eK78@5>7\g,I(NO;21H6/4Rb9KOg+U4MV-gXYPg61R/F;A[Y[RSJJB[_A^7
1c3VbC<2Z.BTQQ&G1QB[SB:e724f3W7=L=FB0?GNb5Z1e^A>bDM\>4MNaIUQ+#/<
471HT)CT]31(:X8.McGZ7<6//WVEd?[^0+@EBd3WW:4IO:)HXH19d4g22U4#Q+>[
[9f7;NLK3NCALBEHJ<UZ5HGA\:&_ZaXJbRHA.V;S?8K_UM8<Gb].TfAN01#;UI+S
g6FfM3NO9U6D2fF,S1EL0_&\&FR2+a;,T-TcN@():<I5a#f[e)S/TJ:-4C7.dD/G
\W;P@A>XUY3V6BE-fAVLcT<Y,#]IC2gD#FH60(1J9Z6g?d-W:E_MPdTCN@<8^C_2
^W42,4f7(^:TW[4+71>_AFX3[BL()<O?FO-UV@U&0Y:c]PYS>g\LK?MK97.O@0A8
INI1G3^J3#0e;?8U\cM;UdV@0X.e58^P@_]/,1Te0g?S-BVZ>b7?K]B@P#Z(G<)^
@(/IL>?,@^DH;O[aL=A^K,XV.3Y;+AdC&Q\gc;?7OJJ#ESUD)R0a\_28^7ZE[bL0
_eee]cA2(cUU6WF&06X-eH1^VaabRC6?0V/7MB<b0b3_I>O(]V6Bf?FWJd8B,089
H6M65:].I1<TH;BaR,]Sf5MeM4]L9H&:c]JKcJ^=X94??U2#W/,2RVgHQcELc/9U
#CLQ>Qe<&)4&[[Z[99.aK4=6)3;6=2eK.+RG6Y8gKP?HA972ESdN^KA?LU7a;;,]
[=<HSCfT.RPVMIT.6eN&)H1Zd8CQ^IX(ZTX_<C&4&.ZJ(MU0?&5)=C:EUCF-(+dH
RPWNgWGIIA8+aL9-2/L4JP8Z15GMRE#gf7.BKBcRP8&YVIHPg3/gf(EE8@1d=Ld\
ZU]1\6aBF]>Q#bWWYL@]_OLZ5_?c/9B(gI\MR6^_MFU6D^Pd3DF^-bBS4._R/0/U
M-J96\_(BG+LAHb-K)CV.b@cT<V,,aB2)b^a_0@C7=<d51(UKTT-=aDZU,8N=K1=
<GP9-#J?QTZ@L0FdIO[E6REKP)B4X(:g43>.?^H26O-[F]/3PK-[=8^8-RI=.V0G
&T[QI56(b9)gT:16GL)Q5O@B2e\>7Y1.;BfX);S_G^Eb>TG6Q6dFXQGfE2FT<(ST
QK2B,R\.bXQ;;?b.V/)>8L^f7?a58]YaM+?5V]PJ]J-?D4\:X2>a(Xg=6BU<G,D8
5C4NFgV:&>E_R:g4T-NY[E/XSJB\O0I@P&7@X@dZWb7)YAI[OS_-0d2?_)e)OZ;U
Y2;/2/B>ET>O+AVLdcGR0aPKHa6Hd;2NRXK:A-C]2c17]aG:3ZGV<Paa?8HN+G.4
2C4f/J36_2gX+..G+b#5.Q80bCTJa?;eg#8S\P_38W+QCXH.IZKXQ6KMFL5aN2<R
[7,eAD&E(?U5eQY<OW_LF)CO8caQDP5&ODG@MI>eBS1geUfWRIS#XZf9P+_O+f=>
77198a929PJc&B#FVcJ)a3[@?30,QcT33DE;QQ1+7Vg(@9++0\-OU5_5=:+&],.2
CUSRN;[E=0aN=3O:^O=F>=SC-YM+P1aN^8eN-ZD<W(NY:GFL3:9NIODc1<R0>(^J
)Z-J_;Wg35U4ZZ4(\^J.^MS:d)D+=#KV3:Y[F4TTI0]=A[5G:DSX3fX[fLB4D22(
<L;GYIXOG^13.B^C_QHJe,(;IUR,BM2;_K1(K;(N+KCSR.&JB7B^\8OAC;VZc.\)
ZN=U>Y8/EUL1a>2O)M,Hf1I=H4+a=Ua/cYaU6C?+8H@,)29J4N(F-RBa]DYOW;P#
^FA3TO9/+9:B1)]GH-d@g<6^AS#2+@<=M_-PX0d:,fGL(K+d#f]b9L8@>A[,Rdg_
K[)IVW_db;6/38#_HI^E67DP+9;;Wfa\A-UI165KY@JUV)J9=[L(e-CgJe4Q&RR&
6(JSQ6IXPg@Rc7;7H5)-PGJ^W7g&7Z5:O.Q&C5dE++8?^8YZ)H[gP[_\Mg;G^daR
Cgga@5=+,5]CWHHP/194S;T=9E9c48N08Nb\=<F,A912P400+U@42-3JPZPS2dS]
HNU51a:A&9H[dQ9GLQA5#D8CH_KgbdG60gN,E,b5>,O5TG^R@4a3SA\a62>#M?AY
@ZI?DM8Ue5LE9/HFX^W@K7:Kf+8;W1V7HANYNH7[fC)&cH]LS6NC],K&T3=L6YP[
>&fWT.gJ3-,+_/K@:<:ga?=[K+[K?HDTVG;W8?JWf9\FLf:JRU.E5/UNCNS<\:gM
2?Ic@K::A8<7OJ#b/YF/)94fNT[?RDb?W:Tc.?LCF+#Cg_V#_e/b9+bB5CRRb&cf
)Z,=e#6SgKY01_9ZO#.7PCZ[F]2BI_cO[Debdb5>XR?;<CHdO\1E>#H@PeJYLEB1
:fe8[CDe\8H;[DD<(4&Dg+CHd2SJc1BW_LN3ESR1gT<U.>:W+G<67dP.BO9X\G:R
,1X-g6WL@+H\;ZB_\1ETQ]fC,Aa=L3V&.IK/M_Z>f&ZE[V(GL,/_?7OT9FLba4?d
4HTOV]^fZ9Xc+,@AE/V<?B6=3eH>,aK,LZ)^].<04IB]Vc:Kd85;bb_?9CCL)ZEK
/-bX)24<0:(=\\K>]REe:eGb;3b4V<VXc([MMAH:SP[b]+eNY^b8U6)<gP?T:\(C
(8P?/++2bc_?-V_M1YD&Y(D4?N8fa/ZP),cO&YFCe8,M>O&)[,TUMCLRP1WI/6#Q
;@16U1(8dLY,cX5BFXd=JBLL@_-bL/S(GL<1D@O_OOeKZC9[5:D-:^4<9U7VUfSJ
8+Ba4d81)IXKZ?G/4fGG.@S8J_Z+gB8g:-(->AF)O-.Od6+@:XgDZca+Q?>LE=Z@
M[[B7C\4KHQ6]7(#22HO17c./TfBbT5\_W&?T+Y(G8./KV8TZYK/c))^Tgd+K716
4eI7CL/+^(K;N@UT,)B7Wb,AA\;GZZ+=5-\:gcKR<#@Z(\2((EATUE_/-RGaWJZg
9)8aQ?T@]<,N6&6F1Z?V;;[PY?=RAS_8)@eALWZ]M45W7HRI&Y1D8>&K_#=>60HC
Bf1&(PC60G6(OWZ5HR,)P+,.MASS-BBILPVK.1OHV1BR4,=(DgG:fF^eBDZNSLCS
1.\YgG-]G(eK?3](]NW+=VRF>]24K1/OASU>AP4]WPKVH1W6<BK=S@JX-:DcC\dG
C4Kb-.MbXZU\dGd4>=H5MGM6)FBFbH6F[8@V_]S8TN1-Z-5afR,56JIbKD+&e0A>
7X0H?QdZ_K/dO;cUG7-V1QPOU(IG#a;&@&TUaWG,dH&D8<3,AK=]Ee\AX9)d]1UZ
RXbAfNQA&Ad+B4LY0ZM=eI7?\?c3@(>GV,8/6@>/T62O/Wf5#;/>bU636JA:g]WY
/T:5TL7P_0V_HS+9O-4bgXWANa?EK#HS-L7PM#>?0(Y5,GLW5/4^bO2;3H_4DU?E
:@Sg?#D-@>IcS027.E+X.L[X4EEQ(gD0,)TbFg-0CB5,H=ILd#/EOeD#28@L027^
c@f(FUbVST)__/CT+((ISV^7ZT:aL6/Y]@Pb@X809C#??6EGXH7aB)3_,\-,V-#f
TTb2-NDge<)g\)7-C#&W^c>bRUb5K0EUa=OBaZZ88a3;#V,3?U(4f=C/R;cI1Kd_
-,56(U3POf:<H536e29TcY=Dg8XO?2@g8;2)MK)?#[H5Q-VIT7I_8B#I?e:Uc66+
E8OBU<AdM=NPJ(\DDBDdfZK,2N,)R?W3>I#AB4ReC0NZ>YIT;#4VS7d7RN(Z09:9
e0A=SIHIILJ)HO=H4^MQ5LcHUH^G+O)&WF8S^0@EbPZE-ZTWG;T@ALMN9O>d/b(@
g(T[eBN]J9O<8=JH##C]\C>P_fHM4MWC.M>38Tg4=:S;2e>.J0-Kga8(><BES[+3
3[<#eF4K)#PR:[d&^ICQ+SGWJ,:(/98AH#]^f@3QJXN\@#-f#bQ#GTaF=;V@..4M
^;=E)N4WM(36FMO?4GCNC0#eW0>eN@TJ1e35I-^:<cf>FNOE5CgETXC_/Q31_;69
PU.A#W12>cR?\1eMHc].b_3:Q31BYRSEVd\,.<&3P;C)_7_M)GT4=6=D=[aMR)?8
+a3V(.^&19-3[]7.JA^220N8>M53.dL6FV33GK[5B9V8)6U:O1S1D.&&aM(:?GTB
LT]HTc?028EGKFEETS&OF79OU4KA3)a1)TNf#1V_(LP_P79FQVT[KM[71XT01=Y-
X=ZA.Z5BB@(J[S??c6DZ8.a1CPd7bffYQG?\Q<4NT,;YaT>AFZX3f<1,ZRK?dU7B
\fcdbV,B?dQB5TPQ1b^A0_[.HT=^_?#<(e:HX9_gL:UZaY]/LXBUb52ac0Ng315+
-J93XR3/+MM4]L)5++gY5Oa1NQPU(<fd]N-5:4e>b6(C+]SF<a6C,fDGBO=:(2LJ
[V+Z68_7WfG7&8Eef\eM13fB0;-8C0f[9<.cMJ0)4.A6\^B5M-W;@ZPZN_K+<D)b
2Bee9^#9]=LXX,&f;H/+XF7B(3\Z,1\#7<-T<8,1Z43)SN>9X^+)=60@3WHQ8K&]
[LJ-2ZGEg>[HMZ-\J>7ZaS66@]b\f:MdO&#]-1)@Vc88J,A+UeQNCe?C+\?(QeQ=
6#6Z:[&f&.9a;gS<7H=3X^PJ2?Bg.KG]-VYD;G7H4CCIgC,@KSJVBM;K5ML)MgdU
Sg:UTBM#X9NGZJ<.YYXL4PC<FG:N@GV@R=7fA0<7<(8)A5QCdRZYNg<^@)QS48H?
4U8CaDWT#DEgfXZ<.9960bcFe)bA,>>?V[b6,6]eb,JZBPC7/J88b;C>1QUSU@c5
U./.J?_83=G]]1.8I.14DZ;Y^6?X(3RSA).@3gS-^aR],+2eMT^?3L1,B_RAeU0N
#_K9,F.>e>YBPeT9YJOO(ET9[=KT=UZB5MOg3>ZMaH;?Y9a]O]bEY\JVW--_:(5W
GWEM41XT5>B;;F,]GG?aeH0faK3S61ca1R?\]QbXdU];dLEd9EY5\0&.<ZgD+K8H
aNPD7/IMR#;T<(0,=&aR:Df33ZF5^V&N<SX/_7N;b\Y&^<,&;X^PBg253Zd+Kf77
?6f1cT2VHB]=?5=M?8EE-^[F+AQ><T6&<.CcV=MK<=eCO,6V.HW5=1KRYL:[4^P#
=XT]WGeCEYBA_)d,(A4e7<+(3JS3<X\ZQP5K9N]UQ1C;4E&6JLT,fEg]=2d\68^e
R44AdG,Za5P.(eZ8ELBVHgO/PeU6G?OMNL-1UU5/@/FUaYQ.&)ePcRC\+L?<aO?O
0(5@GV9DUCXPGIN-cGPI)/EZ)XJ?9\[:O:2#C[V=8<GD7EMLBVI)g/f0P[;fCW2d
Z:gGJfgUHZF/g[/4,<H5K1HSWERB?ICLHF+UF)c82DHTQ4T0<Aa1OFC354E9:9L>
f?EP/@CgXVgG@6=7cOQ7:4)#)d>U/@-M_9YC5BfgaUI;0OC_39RUG8<RS7/2cLa#
QK#3U,@[&cR1Yc[(W143RQGb68a-g_V>SNQAZ7C@Q:]<(WbKWWDAJ,?3XbC]?O:-
IEEKb/U4@aR)XLe&8F2)eI64;6O57P1fEH&8.EWRdM\EPZ&7b[5geO-J.&QQ.H+&
>Ye51:ZCf8Y0@V4)E98M<?fY;H2Vc-^PV^^bfE1)P9I62egH;,cab3K&Y8/GcC<1
51OI62,W4ZNf:d;I-VNGf9SL=,aB-Q#&;ELMe+P6<CScI]AI#]@,7a/faRIfN<Y,
KGC]NEL?]5QAf\C\]([24W=PCdeJ7-a306FI@Je=a^=]08M)b@;=X0#@D1b5Y,.Z
73U=[ZZPCZT2Z#WJ=5:=PG96(/O7YI<M(BN4/De\36;-M8&T^EEa0B<1EK1S,Q8;
.)Wd)UW:IC?eHAZOe7AC=_=aJ4(+3&J&HT2263BX)+OJ33AIO1RY=Df3VYI<5>D=
0&1=F24[g(431EDL.Q9,KDTMg(GabF#L4#Ra^T8]^1VA<V=-L)28=c[W:RH#_,Se
9U#8_\W4aW.;Eg_66T75[4>aY<(LX)\6O+S@[gJ.HRE-7A8^VDJLA:f@<I.-==X;
?b5K3&&B0Og&A=eV<^E_(8PA[W[&RJ/<Y]@ZLA,JfNXPC=JcOcf.)?KYKHG[\SF3
?U:)=NAG8YEO_/X#NE2G.QdXT=Q^8PeNZP,(8+#>X+Q]EAD851YZTA[0R@Y3c@E(
V\HdNVD9SQQP3,Z<5=Wa;c7<b&POK,bSGG0T2g9U2AT@8JUf<U9CBI(@C#4?>6c)
[7=d>X.gB5gJ,5JUZL=0-+THbUI(f<5]2RXf9GZG\2\]A2b:;?.PZTSC[YZeZ@RN
Q@?ZI.ZR1<ZUQ21T-f:?gRcO@MBGO8#N6^bbW#(b]WN_+J4g>VZZB6)CFF/G>Q@e
KQ7C8&<DCBH(;&4=E^Z^X)19D?)K^D&61RddG(.^Q6TPf>Y;#aM)dE<DRg@G82Xf
_MF+)J@)Zc,Y6f^R20Ig,07^]YH;Le>NI_I9O7+YS?0YbB@H?dOa&9#d,Y:[9&fJ
c#RMNfQA;,YEAU@^ZGE)(=d0R&[-?9JP59cFH\_C+_CgU^<Q?YN8;KS#L>=0d8[b
X)d+;BSY#W#LSe95GLP6SN<g]LNa1fJaCFfS?fV#<X3UFQC2:Bg6f/AMU@6#CJIR
Z=T8MXP=LN9]L<JEQ)-2eI\:c.#6?5ZLS<Yb9:_U)B(A\_1Z?.>5H[&#T>d#\EZe
eQ@#I(,);:9N0E]\c=.-YK3,PFgT2e+OQ^Y)a0@0:OV@O(DTHI+F>FUJ-U06AD8I
_,eLYfRS]:R>Q.?.:^^O@OPM;9;WN4_SUB(4Ba-VcDJ8g9]P@)\@/G4Zb[VaSKEY
J6G9TEc<-T-=+&B-;ON@5/Hc\TK^6fHb]M]6L7FM3GZ=ME:5[R4X5dc[;ZRFg:/\
P1eC>B@1dP[e)d^JF=OP=T.[&1<</O5_8RFWR/gB_-C#D]>0Ce+<:N+5OgU\eSS[
3O_C/&BX^b(M2[&F#=.VH;Z\753_49QX.ag7Z+?=D^,Ca&VTJJ>DR<1bJUPb0)If
>[eKLSc?+#4b>ILUcQ5)8UfC&7TdA)E4,KEJLO@[^bbM:IZ#c<NHK>O6KU+9,/#0
3[O3,,S#>[E.DR#A1T>9Q#[=GLbgCY=@@>F@a?<OR/@:H[bA<P(7#-?#SFB4DV/I
A>_f_]HR4]=_(KPR_,>LPO&GfSVdYd4:0J+).Q4BHM9P@HPF[,,--DZ8#fG];_:G
d:A\Q9JcUIa#MGYS4^S7QV/)]ZQ]]UeT85_XEK@@CR[O4DJ;I&cR&,_c.4UA0>TJ
W)>6V#5#<6IV5dT@]DVV)T:27\JA6X0##-CYB8J5C.;8S]f7&C,1f1XWH@2g^U=/
MBgOVWAQS(9/Dc4BS#2Nb]Z)S\H^/5=:FPT>;<X@:/.3UDVCI-bcAQFc^D=XYceB
cY+;WLC4(@T2(]7II?eZa=-3bbf+@]aN:RUJaTS3]0g6STE(9:RTaQ;V+4B#OW2Y
>(E,aVdf2X5<dNgE^2c>D_CO1-&+EAG+8Z.COQTA2#::<eaUI8b<c^,R8==>JL@&
?=?1NQ<Y?OQDab,W.CBg#g)(8WdIPe:\C[[fbAgaGEX.X:MeL40[0B8E3LO<UfZV
>+)fgR^3d)EPU4SRA65+fb+Q)\<0,^2=HC?DB?]2b;?]]U.aYQ2U>H^Kg?G1_/=W
5VFB?[He#D8=-Gdb<0=J7ALBI:&fd^Z@=6)>,I=>2CTdY<[a6R@WZ]<+KK;Ya3#F
@f(-RKC)?7UXDVTHbI@F\TTX?gRDI_BYSffB8]bJQB]\<(4ORA\1I2DT6YX/aCS-
DBB3<C./L/gbKKQV5e\SN,#W#JFF&R1U#:#=T&ZS/.)a/L2;;+?f;TS3LQCY3+]Q
>U=I&2V>BAfcMJJL.YBfTcO>\VeMB/<HbHH71;=#/OP0[#KOUZ.cabJ;T[KT:DAK
/.7[BG>QX0I,6TQJPSG;_BB?+bNf#TXI856<O/)f5]MCC(C?_VUHOU#O20)8GTLH
/Hf/Q?(e>,B]Eg6TWBAI>O5eTdd:G;#A7b=AVbM:cJN;\Ya/WA[S]<gZ@,[U;aS:
MH>ZBWPVRSMde)6d2FD,e#O7R7^4]VYd+63H[b?eRa<d4[_GI+e&F;7X6,b[SUf/
c^eGFbYC#CI.aJG&6O5cg#O+eff(W^NG,H1Z4LY36(IM=cQGB-6bd>F&\(b)fF-Q
F@dD9=?&0gM@0BS,bV@TVG91.YD+_d,G<aHK;YY>bW-IA7Vg@DP:#S-<].;REXYF
T?AB:?&VUHL_A06TE;Ed[A[Lb+@IYO7\F;A,eHN-9Cc9C6bH^8XSKNM=>748d&JH
26\H7/(eMYG?bS#]IU8(IWV)LcAE,_0+aYEM\BYY@c<E].)K^(,LLI/f2c5I/]9D
.b-B8?^DUV:TY4cSbK_gU0;g-6Ef_ad>#^>RDHL,^TU\4aW(,;0a[/P.Wf8L]:(G
cI;a&,,Zb]I?aT\L7^FZB7A1-9]I:Tc]M4:F2V4F@^=Y<APWf\#R5)b<\d]?0DK^
d3_B(V]+)24Mc05d=Q2#SG62IHX\4?]6.&#.7T[TS6>AJ::;DVY0M>(bA,\-T4;5
aDMD[c6AOS1Y[KY,dGN]XUe<3CaK(UWbR=71L<P7.&>g9UGE(e&agg/O9U^KQd@@
eWO)Y/,5[@/dL4P=7<-DVee>U#aP((EQ4]O/;IZe]?=aF-O+U#V/1WJ(8P/TD)J/
8Zd:L)MS@TJS[ebab1SE-NYa.Ie/(]HBHCUITXU1ZLW;<)T:&A8eG-#Y.a-@AIIG
\YE.T(HB[@4:HT6cbN6b(PP&+TF1+6W<6d5N>VFNFOT3](K4+UD/B)8E&R@@5>^9
7eG2>&0e[L&gQ(L]NK,MI>@?G_D_4gXA(&0^=>/Z?I.XN^KS#G/:PR0OH495)PfE
W9a&gM[Z)ZE+C(a_X?P?AgJUb9-)g1Zg@MdTH_J)_g6aHgWPHd51^f@>B3,]f4Fd
=;B=9b@0A=&@\AZ44U2C/3+7HE?D0[Y^#CU.AX4#P_:CdZ2<4dgKeR&e=#70-\eI
;2f6CCQ(MR0W:WXN2)GGFK?MS-)\UHQc_L6(329G3Z;59_Sa@(LOK-72c:RKG_C?
KVdIe9fM)C#eU##(5;:9/F(I2./c72ZSW/(g;.ddYg?6X5@=LQ/;:S/F;YG2HBO0
cR3)I-4>PM,\P/E4S;3[+Yb[]BZ,<WJB=C2H5JVP/+2<3ER.[\6GTeMdR=ZeDZgI
:OLPLBRHJ\(-B3K2Q4dG[A,^)(&KPIeDO2HO2&L2,]@T9SN7)dFN=IW>]_)d@H:N
^#?CJ83<Z.SbdC_Y_EN+Z9[+/U;V\NdGX^?N]9<c]67@JG-+CA^Zf+K0_5>RQ]:8
_M)VNeBW_a;]N\WdJbA+>LSOD>)G#3U:;B2VAMT2AObf.V8T4LU\;CUU\7,_.8UO
4UVR7[&GO^;a18CaOP5ES=\#R8Z\<0YPBeb4B4a<=cAJ?SW][g][G_EP=)I8#=-I
e6+/W((0=9_G5Y\00JR?@Hb&CS@Q;d172GQc3LeU5/4W&K[P,ER<18)^-Pb47[0]
04E4;>[c:)6[\e6ac,=ML4(9Dg-0WVWc(]_BIg1+XWV0:H6BC,CEN96#U5eg79AF
D3<XHNZDM5Eg0b?[7]68[]7TIMDH2N4#;RJ[R^X4L?Le5eU?fU]B609NR9E^fQ38
77@TD83U<:.L)68d9\6.8)#+HJNM(8=&R1=;V3;PHJ&d@[#@)O_&:GI/)fdU._5N
0LUb?1:1=?MM,g.\NJSOY)U,^b4c5WMF0KB[6V2YIaG_6+AC)V4GEUA35dM9Pa0a
TW>71@EG-f;506M6bgI;MCA[b9>#A.N>7F.A;ICCV^#SDfT<4K56:9#/.)\Od@2)
>R(54b(dFee.UeVQIU<[+3e,.6/+O4gSP[QY3LO8=)>2Q<4G/a>OSHOTEV#6JH2?
1G?LM0#FRM&Hd2LJZBfP6S/_DH5>Gb1\<VR^A6R^J8N:M(,Y=aW49DgUY)8]6Bg9
;_HKb^3QRFd@:e\gL_-S60Y<#0WVXI[Xa/dc7&OPZ00TFA@>5=TaBR0#=>,N[/\D
g&+7T8&Z\L=A>S(+:/42VEY181/0\gKS@f30@+[X+V,=HdM(T;:J13HK(6FD#-]#
@gRgYb^1dL=I2YfAIaGQIfS#V_=I7J&QM<<VB_YLQVGBSP1cWJa,?&US>X4>NCHe
@(;1)I&>1Rf>[5]OAX3?4]e5B3Wb3a;1H[?0CJX9;d6+D=A\Nba6+ZB7#EMI_?ID
Q/U1(&&^+^\;E7+Q^MHC^Q,JR\Qd[9=E5,?C_M?f=1>J:;=eUdD3@Y(+^=9>P1Le
,NaZcUEf]AO/HQ6L-&b4?6VE#3\NYC5\da3Ia96C,ZOY7f=\J:\\1AAD.JG<C1/5
Q.cYc7V&0C#Z^HP-VcL0#><aRW<N)/4<5-YY@7[f-E:QVc,KPJ0aNYg[0\J_J1e9
EKN5S9]K;&\5U8?H(KZ;45X\a^<9T9_A_=g>^:2>F[6.FH5gD9^O&=RWLGRO6+,P
a:-EOG\5FD5&8^GbJDa+9T#<T@\>b(fS\X(2bC#g4_c)/b915dM=X\-6[OE_^g]M
c^(+fO>R;?4P>2;cDD:POX2/\;IPc)AR:VP^aSK160(BG9OHf4CR9@,77L^c;TOS
1e9Bd,E7D1;NA-]1f#PM2SBC&RdLIc8@KQ0E&LG_5[]WH^F4M6>cE@Uf0K?B+7+I
>Q1&^-S?C[28aARWgYa6.2S&NX-2)cWK]BYT(S#]P\c0UV4T8:Xe]:3>S8Bc.Sbb
J9[1-/QT:XO)#&3MP,?9Y49+O4QV9F,g2Me=\U;FPO=[Q&G6OZC(SGeS#PDVQ:>,
Xe;R+;QHHb3O(H&NWBg5B48YHfaG>ZMY[77bT;V-SJB<<161@FSEgEC=Ye-WOO\T
0IOb35BU7R.;X@H29VJWcDbI7[FJYMXW_X:74SN+-/=;EA9E3#7]fW>a0DU(@;99
;_SQ,QO^8NVg&M:/=Ed#:PQSQ=>#WZ>PZRJD3U4@Z.A8IOfO+-bAd/2KB..Z0#aS
J)b-9)Q,BXWb)?C#B.aT:GOFUM;-Nf.G\):c-bNd]]PP/[GFU_0/RfDR7Xd9;)g0
+cBbJT?]FA\@.?)bZ\1[]M[I[IB<F[<85EAEPKY^,LN&MaAB>UaNb@V&SK;e18Ka
MC48?&BbRT0E<#(<,OHYMCQR]LF\>V)\48M_7(f5gA5Xee-J@^N3<0G4A=44+A6E
VWL;OR-5A75CVZ2[NYSWeD+D[FT1J>B#[O?.S,E=4_gP7]ZM[gOF_8aG>&fA8C##
gL7E0I(_QW<>gf(GK[3-,34=bKU5AZ)0-^M;EP1A0e]e\:;IaIRY8J(XRV.8g8DE
WKI5V0c=EJR0>dR7)1RVIIYBM_]?C)/-E@)^R,OB2R3<N^17eOE+\BZZ3H^a]2e-
W.T?&&BDK(]:I;b6(8&=Y?DM[>[a@J2<YHKS25=OD1V\]Z01CBMQ4)O^<U>4Q3>b
U\AX,eBA,LE<8AFY;VH/\:M]E5.I=,]6Qf:LND,O#N<^677Ef->Q/BbK+E[Z/\aQ
C4).6G2BQ=BW?;@daNcDOIR>A8(,G1/YScSFaMCg6UG?_YZd2K6Y<FLgHD,Hd7H5
+Qgb:0SKH)3d9FfR0+N-aR<=U)ILX?[98S^ZP(AM.NWF<ACQ(IQ929Tg^daF/UcV
QO@Fbg91a^8-Z4AB06e_^K\<M7<BP=N+g--T#5@5bW[DABT_S4[eI@(4Q(ZD/5)8
TS#:f9,33&ISG>^#MHad[Q,J6Z:a4#=JUFT4B<5R]U9H&PF?\1FTRO+W4N4/Xf^^
80X\+>\6@FB+,]7R38,U@I=U_?S5HDGRJ#XI:Z+,(NK(5AO187\>c5-Q[]T@FK+d
eD;_H=;0?\S?PP6^F72f>Z7W+TSddV38C#--EJI&GdPOb\M#;d4><LV/b9e+C_@1
]QeT/][[XX>cLPd)IJYCC,bUQ7IaN>9OYOC=1<Eg=LB7U&0)V.Jb7b8@WO[]P\K1
1H[W2IZ7?^14QS&VVDTX>gSM;WC[+K.JWE:>2_?BS3=F)2Sb8U\X>6Y<NZ9_JU##
;RB_RHTaR=4MW..G66L7Y>YYC<TGfPX)&@Z>#GGL=A])_:R7e_G+SAO1#BNBO<NZ
TQbfS=?<aeYRE;FW)GTK1Oa[[D-<#-K/,>P)B:D^L9J))4ZV+62P;Ig4Y8D4\.A+
0>Q]3Ed_,^CfPRT[FANcA0&0RYbgfGG7)W9N66C71\#C+#GdgTe-1E0\R)-P]&a<
D=/?<:5^O_B,ZJN-:1\OIeC#A3aV=2H&fS,0IP0F0@&L]5A_@<R&gS2LQC9J>g9L
9K7)+Na/,;@AM4JYMf/[VCJ[4AWN:gC[&R45E,@cYA2G;C3df\V-9MOb,R9J(&&<
FD)aEZZL\Xd[G\L.A=2BN@X6Z4aQ4?)V4PZ#P&7Q[22dX:>(UT7RAd2^Vb<RE)]X
<(a:g32<]eE,>;=XGMFU,6@:.e3/Gb0XAZ#LPB2\N+R[\]bDO<-DH\>>KD5ZJA2=
TF>/VCY>(._D_Y20U-]IVJ:^C^]B+LX+eeDJ-7E]XMX-IeX8X?JH06I?MUJZ44G.
:]<;@87BBM8.W,#?^fO679Bb<8eaKXJ+bH)fRG_U5===A/+K?<?ADNfLJ&X?Z/V=
?\\Q?#U6GG>&c0+2V>2/;RF2>@>O:a4RXa#\WL=a+4.JHfR]7YW7TWcgKM#+RSPM
5CFZYaN4LINMRVW_#XJ6C#RF0?D(4.J8HV=Gg:UgCF7,F5_#LbB@,3OQ/Z1@#3]A
#QFDV1[B&)DK8WFDHL03>G?ES\bK([H5;_1U8]^/g34DV,+<3F\4_c?0ULFE\GeN
7MKE;7\F(V>Vg&(c\6T/HcU\<Aca(1#>O&DgD>:I@_8H:,]G0AY4JQ<+dPN2^Z\)
6:MB(NS>g6FCOgI3Jd&=@..BA/8<c^XAKa_-0]P=3bF;?_WJ[HB7;BQbCUJE0IJO
=F?4c?a&GU1feI2;d44J+P4[79U?-:WN3B]fIRV9Y#Zf8Q;F#A>?J[gO4W1/1:6<
5;IZRAUB5X7GZO=BLHCZ=2KF^JY6MA5>E#2W6Va.1B:D(ET_E6702KLeM9JG-4-6
P]=<&HX,71>&#8/Yg^=(YTR9A1Xc<fZ6G,d0F_O]^5^5)7We)ER(bCeg921DXF-K
TM,[6.5=IV\),5DVT5D7J:d]fB@C_H)]&\NJVUW?>0;dV/2gOL+.E[=4&+_BY;PV
<dT@LZ]/8,B;IJA+@D4_JCc?(,8WN)LX[QJ;6HN@)/B^;Sc@4Ja7=PSL=&G_M/\I
9]bQ?C;733:6fQ(4.2e3[2=gFO2R_N+063e#=5fLQaE-8W1/A2G?S+](>4WGe#K5
U>F8C-#JR[/(A^L;/6d3Sf4C3,3+QY<5E=PFLZ_F<WCXPE6&aEC&\\^.)+>4N2)(
gEdVN54VS-H+WG=23JYdZ:\Z+;#S2BN81Yg.gAg1eJ#)2+E2DOT@9(&SQfL-H<XS
#=P?Z=HAcgaE.ge+T,XLM7;#d\1&F2dX,INDbN2S]I)H)[=X,EY4RCZ@C9EcCWKe
FAeR/bXf-KbcEY3ad>)V]\9N;C#US]A3.@egRIHM0@2d,A5OC.N=:O^>1TG1W?/X
-FONQ\(,W),gFDd;X<_a0e+=Ge2<I-gIfT6WV7-L8@7c]]_C(F\J?:>,]Y[\=.@E
Y-c94[9-@<?IM/1NSU;4]3X/Y/58XGVX#9T^5-8=@>LG.U;HDg+4@R\F-[=.H)cV
f^g)0@aE/G=25eBg8Z^Dd6[A7&]TbF0J.?-:<fVdF,ELI?\][V.8V2gMBY?NTHFT
^JAaGAd:5F7P#-X<KYT^5JP_70dY0),FbU^0CYf\^-7gCV<bQCT6#c6?QM>V+8Z[
DWL3@8RbgYBY,I=g;N-BbddbTY2F\LU>#HG-@C_ATBaGdU=3NS-6YO+3P)]K-GC.
NU3D^#ND[C7GYIb2LZ9.\]S&LLfc1]19>:6,f1YV324)eO(1WF>,1B_HgK&YCJ2T
N_YV:S;^1MGXMTBDHdGA2b<\Y#YL\4,V?--PXC?5#3cKDU??B)D&F=SO;Bf&RZXe
=S5N<LI(K]7127gS76#T4Z?MTJA5A4OKL[80CI7L2.Ue.TROMNFaJ))gK8RN8#C?
7I89Je?,./6)^A-6C(<LYE^6>eNBSUTM0R]?1g8SW(.dFNMR;)U[,RcDA(]Nb2V=
C39U/C+&81ZM7&\3g3A3BOMYNNe-:3MJDT,N,&H8X=K7(F?/-dIO?<WC=L97g@68
YI4a=(b7^^fL5FBN&B.;b^<Hd/4_.5S.EKLaC/E=/8Y99V_;-[C7B6/Z-eD2e4E1
3NK1S[&].;OX]K9^RRcB4XKbB@\gd>84E#4[VWPZZOI58Y_?g;WTF74?\)LS9,a=
D_K)FPW;MUB;,A(O2?GMX@GD:BZ_@H9C<XS^)[E1(,N9#X,M1d[O7_R]>T@).68F
=IbJ<BVO#IVHZIdQ7#f,&(K3RI2J+2WZE[,SG9dHJdc5)9YKU@^N9b<K@B-HG7XV
8bVP__0\TF:YLD(4F;2(U.#dITJd:PPN(+J.^66+5V5/N-QFY^^0K0XTYP_;Y[EO
WXZ2J2/KB8(E2a7=K@1+_[M&,MK7f.]E=V+VXbKfL=70Y+RI=Rb4YbE-;Z_)3UU6
;PONC3+bYIV>0./S3aBCB@cN/]7X[9MR^F,M?(O4H_]/TMaQ\g.bC&]NJ&-R(/dW
Vc&gH^;G^URFX([D47P0ZZLFe./cVNG/O&U;Y+0B0<Q9(0d0Q3g:GYe;,;Xe(]_8
[<Q<M<])<H/fD>[U[FGK4=7VD@6LIc@,L-WK6aQ)+,,H<BbD2d36+Ea@B..3eC&g
Lb<[P^+)GK^LM6.Gbb&aOL6D1PV(2_I[T&gTX72G\XM\T<HO4fc9_A?KgZ:(^R\@
/,N;W;3.@-fAR&_Y1AE2QQ(eH9Wf@5c^CFW=>;^QWZ2P@M??4E\UG=(@LPX)\>14
CgB-d.Bc:bEZA@-?A+8BbBAO.TS1ed_=9G8P;_&:+c<C)Of-Q_5+<ag,LD_3A)YK
SF>ZfWY87dVR(GSYAf3Z^X2?5eA9J.ZL/)b:3K,T9U>JagC29AJcDK5WaE092Z#Y
fOPXED,0^:Y<(3-&T8]bNN.DN&E_E31EYBCe1XFHg+CYWaRQLNU]X[P<NUc,Wd/[
5V,/YRe5ZU)4f=J?aI+/RG@JbB7#cOH>IR,4/6^.<O)b,UIAW4LSM4e[:eB@B)C:
0-QQB_T2=fU,[[R(G:8O4JPMQfV&/>B26d.U#Y-:^fDSb1(KLSPa+^,eaJ)0;4f>
g=[/Oa1W5[S<]OX>I4=YX(bBC-&,DI4.f=18I4I](?c&_Q.VB@0R;8D0Y+OWZ6FF
QAJL3IS[KgbRL]?AU,8&.^LT:\+7J5]fNN<D3/DZAf6?e23^5;8==LT50M1/<,7=
&/+95gO\X1e@aA-S>&MHHL=WL/PeCI#DT5c?X&#GcbX6R)aZ+9+M?DfDU\[,@;UX
X7@)(D?4=FGcUQO\-cN0)(bB^,=?<5[NH^4<D5[4Y)W81S/K@-AW]7dMHd\a@JZT
U/GVdV&U#T_Y1K7Wb)_C.FRPS?D>[39VgJI2T0&_J,GbM5#=7XXFgU?Qb;)\b5HY
+=IC4.)L?eA&c4]>?bE[.K=FISD:_O[3:&F:g1S6X[39TF8aY]Eb^C(VIZ&a9=-V
#H.eRb#af<+_33.5M[6?d[T(PST,;+9f/F0[QGGZfM?.)@H,-:V+B;4bW&>MPY.S
Q7V;EONJVWJa##Gb5XUS7JX#f&C-\>T,/R(V+bDM393Z=Bg/NG^DG14#<WbPf4CV
8G58=O5GS17_]&+20==.1fU2We524KDU>Yf8M@>?#A-C_TL45b-8T8AN.15Le687
#L0FG<R1(28eT_;,FP\KU(2<EKZ4_g-N<BZD;KR+TZY?f50UMXZA;&Z2OF<^?[bZ
FA_+cSVU]6B_0&a]WV56=2=[]-fUU8Mg:6M\(JS9W6;JfC[BSNY@[@7[,eBB2\Ba
3E4?.U5_OJb,]E]9fF&Kg)[+=1L:GW=E=)7.UA2T5c+UE\:]ENA3C26;4X\gG1cY
<3A9J12J11aZ9aME,(\g:.V[b39/\BTbE7YL,eARW9N4Rf#@>1@)U7)7@,?fd4FW
^c,eaLXIN)[S&6&e[<,.-2Rg9HYad05f@GPY]W@7#F?(Q[W<I;9>@fLYG;_X4cE+
g<XCCdfS@cP&6:\<RX7_bTCB7X^NF<)XAPcc,T)X(W]E6<8IS/+Ce+Zeg=OE19^:
NZUSA0#H-4+#-)X^N4IT-XN4VRX,>V?Fc[X?P5X.8]U-]F8Y<_[Q0CS=&@3YRc0F
18O?4;]#BD,-M=HcWH.1X,P_??#KZgBD.L4E7@(0]^>=Ea[>0R4[)X\#/e&dJ-H#
8K.,7Y&&&0&X7?cUUC&M6J>7^3=Q:=X:Y2f8YWK1)&3<H(ZLV91E+1TC^-BNTU.8
\-V7Ab./&?FXU1)-D<0M_T\H(\KHKD;FL]LEXUCa]>_RC?RCFDWOD]SPcT+@.PS<
-D,A&#,#D2#,1g#.H&+FBH+gYR=AGJ41&UQF,be8Y02YDgML2FT-_,,e/TLJ>>#:
gB;T?L^eSU1(7;C>eAU.OE)T@R&^0BG_4=[X7RM52_U.P0fQ(^=[ES=5U=,I2?R/
ITV3J>[/>06&;AL8aUO(7d(;\c?=V@dN]T)ZXQP\O.JPB7;P):B[7-XLQ6dWg[9f
)U?gf#1><-]#/FHEA.UL+V^PYEYg\18dOG,P2L-A:(P^SO0/]gUIKGb/[3(?/__2
?/3=TQU6PfXf\_g4FN@P<_g7&K\E@+<Z(Bg;/\TWAWQFF6+13,5gY3@:eHS=<N7&
Rc&KC-2KPF3@39-EV5DK:YdS[MVQBH229e0^eCZ4@E>0Q)3(W\BS5,]N[&1QE<NO
T-2,;C#5M[QPQVO/)J^PL,&b,RgYf@G#Sg;<URWKZU453N?AO@_>5BH12(?I/fS/
O^Z76;#Z@R@#,.@R7H.ZOd^aD(bICE5Z2b2aaeCMcH=[7JL<C<-X#fSd-GI]AQEL
I3\T#[LUf,aU9VFY@RF1c?FS<-K&#-(e^HK-7IPaK,#W+1.<6@[\cH,f4,_GKF8M
Sf/Qf?_)4NG_(1<_)[g=H;ZD#5Q)G+8TbObK9c/NgB[2H4]G?W.IRM9T<D[#V<g,
Jg@L.[]e=WK3A)aL)7fN8,PISe-?/?e]CL\&6GYI[D#Ac.X(b;ZBAc;1#I27S^0+
Q2[:JM,bAT[=/OAReMXQ&#aG8.9d1IPJGPM>=6AU.Z-#4cdQ>SG^AZ4=A<KZDI+d
5>bS6EUT\O<UF+a^NcXBA(TS_AN,/27EE]1JP(6++LZD@;I,NW0+LLCg1?)df8Ye
N/T=,9Sa^b@g&JBbO>@5CKT#_AFAZJ;6\F\:7IO,<D+&D,4-KIZRLH(&IUW2MfeR
L9<Nc4JfJ,J+.RES#C]1CBO9Hd7FBf=FH3be)5Da09Jd>Z?f#X+&C.DN],^]ZG8(
]Xa.g88545#f:(=R&PX)bON0_@8,AAKKX6HFL5HI.-YVX@4;6=P;6AJLe.KV/cZ(
^+e61JYWGQ[+WOaSJ]GULdVe9AY8RWD2<RSGGM+YB]?]JX,-BIOH@2U<5O]+CIY.
a+B7&\UQ4#\WG4^4.[XbdXM](B;IcccWY+^KCJAT_6\8U/N_9G82==#^XG1>c.&-
-<?.^^a86P9E@aY.^gd4RI6NW,UGT^S15]GC@EYF(Q3g7<E_\WU5fd2OIT.\;Z2W
B0(-;,(MUb18#DB4SLU-&c?_95W17KgQ5UK#)Q\IAdV&PQ.eZ#=]1UL[g&4J[cNR
?\<RN0UF]dGKG]65=0bSGB?=&-,IP4JJ2<JZ5a/QJ^D#&UaA&N\NR-F(T,Y)#),2
[:WGc[VI23/Y-N3W.d^bOWX+6=:LUe=>-,3C>YG0-X=a[VTT]=b:56cZ;TM:._ZS
N=DM;&?-f\B-/-6>TdTf>=?K.=1fgOaR&,][,8A:XdA^<Q)(CED^Z2B)PO6LS=Bc
a7IY-T?[#U7#4fM]\JCQ.=JG_GS^Q#@QSF<Q#ID0@&,4c2IG>IONUJOf,K=gE8HC
L1;3ZR+2-c0<Y\;GO&B)+AF558[#5/)X39@JL@X0_f#AcDGcQ=J@R?=;@Z,WH3bU
-4<;WOQ#-L=eG,TM<LSDI07,,dA;-NS/+\2/&d#@[K::[L7K38fKc:XHAO>?a7TJ
T[MNQgN=E(H:2=U_8)O/XO.)VP.=8=U5-7=--YEK<A=:gc\W6@]D[c,7EDK@L]\=
_MZ@f:L73XD69@aa7cYD9.-CMZQ9e)Tf4a10FHNAC\+#=H8AQPe.>6JL[>M@/N>(
V#7M@N,Rg>ND:MG69^W7X+/0JTSG)/I3CF>V-/@Y?#J>-9D0V)ZSMPY#-IP5DD&4
QY0g,S#_bRdM<CeMCd3K_AcB3_eD#W4D.-0,K:7b)HONT_b7.E1;:@Z;@=WF&D;5
3+P:X<;_=I&601aD/_-YE8VJ9E9E^X/YKP2HQ6+K,)FfS,d5a6U/=#UM@5XUO#aN
]71^4OC0-cG=;Zc3e:XNZ:cMT,&:]E=\C\a#G+[gJbg?@Q<a)H(PdJ-:.AL[=LQ2
NdO@)<9:0L;YM]>WS(NA-G<M0P0Wd.0:a:6U>TGCg/W50[=+<c6IOFF6?bc>Z^3>
[W>.F+O;/X7g,eg<R<,N626WeF6^cE#W6F,EC<-BU9S&8?c&++.K#SaWS8A;C_gW
gBRe]1H<SL[:<UI8NF@f^[^/IG8WQbF@STGVdDd6J<Q5=X\f<L,2Ag^cUc4bRg7I
#QGL)HH8S,\.Q[[=;O3Rfb[PE=T391Q5A-\eMCg6geD)L1)X/B(Lbb9\YGG6];N?
ST#;97Y>#;(8R@Z+,aOD@2R0UHB?\&ZKUPEL3,1b+Sc+D,&^UF@J@?aZZ8/C>Z.\
5^P>/CUIV\2S.K&->Xg=be_XbGX;Uad5-M1^:+<9Nd3X/YQX176Zfd@1eV^W(-@M
U<S\0I23]+Z;A6-K@.0e55@CQ7QT7)88RG[9-3(/YWPL1L#)RR56^_@RFSQF(D1M
M#G3]bc4D4fL(YdNAG7E)V40f/g3\99g/,K;R==b1A;[C@;Z>IaO1(Ge3G_PfRNG
<GVeTVPfGZ?aN7Fc3g1588Ca)X&#M2/SRd1RRW)I@,(DL#KDX6@@IYYb&OQ40HLV
e\NIUYIYP]3e;XfWZH;_0P;LLb.+\W\:-VAgI32WYEU7[OE#(IL.GAP5QRTQ9>\N
YOL/]PVBI#.-fI1P\1PC,V0MU\g@e^fVgGZ0[Fa#(9Q4OEYMGc=TgU2P8?e(^cGd
K5QS-@ac20EI-0\BM8>0#T\Z6^.+A-X_G@)BfM=D?.-JB.e[:4E+#ZeBNdJCY=@N
<5(@cF_(A[bb;9a=9E9[,HZF574f2TRBN+)&gEV#EBf>9B^#LLHASbSPRW.<7cBY
Wc.W=;>E.KX8YgG0XF2bNgVKa>-F>?9HLD)BN(C#<E^YRd(e&\gbDeE90MZ2.bLb
6Y8M<2<M#3TK8>E<#.[<ZPCUMNS#=4FFPF5;DW\_AeQO3IDVW,aHSIG)YW.W?<^9
.?:UG<9L>=;TA_WJ420d:fHU\\R,A\,c:RMY4+HD5\HADVS)DRZDdV<b_MW9B@M;
/Z3K<e0AdY&(8F6@\N#[:[-XdQ[O\P7]aDEJ0@H=:I4-DUV?gC-^,UX<<Gg:aG9P
T-Y9Ob8&bMY(76\HCO]?TC9V1QBC_QP^2QDWeQR-=,a+[/Y.VRZGW)^#2DA#H_@g
&c1VKUF;dfY9XeCNHa<1QO5ED:KG,KBJAUDg>@)QF@FM>8F>1\2A&F^@WU8X<g-a
3\f@aT]U+A12T;=&8FF=bKMBE6OA=N@g:.<&b5EBX-I?OT+c_.;>,f:/EgYgUU:I
.eZV+&H;YU=K-HdQ]==IH@?NP]e?Nf8-(Ab6+N(=FJgD\IW6J<#DG@I\1(#PIZN7
58,L<1HJOJ.f_.BE/4@J0c4D(,8:=9IYe^+0,bd<G1Oe(T?Q5bg9W9LI[K)e;_Jb
M<83]e_c#LEF]>ZWP5H\2Cd(#N?.J@K;cX08g,Y;D955[-A2I76L0]7B-1<7MT+)
HdTg429-EbWaN=X#\X4;VcC&[^N2+W1;c?ZI7PTT#16aJ4&QBaV<Z#-D6Cf4LTO1
d&N,DBCf&[<35R&3V[M<Kc6,;0W;](2XP1B,W5,OWVWK)0Ud@,O\7>^^9X4TBZR&
/IaSD;13@RKFeWRK-F/Z;?F];6@95L=dCE4Y;U/RJ5B)gEI3T_PE7EBbE.b?_]#.
H3g3H0bBBMP0G>eFZC&]eGI&U_.gW?g-0A/2:2I5U0LO<HK2<S695X,3&JPfNH;-
L5GCI]OL9J/.\W]@ZAU&Z=J/e[C;])HeS7EVOU(-I39a9BbPQGCB0\_@.e20a_21
W(NDc,OV4OI/QH:VPbbIHA;SP#LZPVc64@=44N4+bHB4?RgPOaW]IeY/L7+#F@9.
[Y@F6Y1>0:)OJeEF@K0&\&_:cdLJ/@ge:X\Fdg-@2g>^-<<dO1NU_2^Qc:Bd;/,W
1c-Z^BDX:d2Jc-[O[HL^341LT1;>3GB?U<]L=[P+FV>NKK\d26Q8>V#2RXT?7-86
R3E/F(/)cdc@Vg<,=<g;:U&8-==T=<,c#F@+747#d7+QY[O8<KPR/.JB#^gH:0/d
H7TZ/U]fX/e&/a25MSaW/C6#P[Y344QPF]\I>6&UFCY4@Bf7McB,EXK,G#C&7Xb@
JA.g^=f.K9CN0U\+N52A1dFT.R2FCVE4?<(1NA1E2L[fT>&AVGJF95V;+F,FK<LL
cEAZ0C7,@,?AeWBS0\#KYeF@_F[-c7;L[<1&[]>J<393CNc^.Qc(JP27-AE(9Q5+
@I]Nd55HHE\Y0Jd(T<TGB2dV>;XAbV;bHID3W2=IRO#HW4;g\d:&\AEBN#ea4W=A
?=JJ841g57>7+)Oa<](I&@B4d<T/2(I^6THANWL+X5@YF4M8WR>WN16K,adR9[5E
,FeaAM[PDd#^fA2/4Z7b96g88,IPc1GA<&aL.BAUJbJDbQB8GM1g+#g])3#_Y-O,
6]g)a_@N@E9J0?8Y9IgFa@T)3HE;&fFHdOcD>Q2@/MLKCH53][N\-O>]U/#b0_D-
NGTX].-RUIWN8[X4C#W>KTL7>&4CRFV)@S.F1N,,BU4)B.T7a#^V3A#M,HDUP]-F
):2Y7+b^R9GNOa2E@[_#-JQT=D[795EI<a+?=,J+2VYbUDGfH,a8P6,,?bdAGX;B
XZ=G,ge>ScWg4e?DNG^::(:Z:0)93IURW:U2TBG@)7\F;,N4]7bTGe4D943?&.fb
52/00O:G^Q26-KP@eeBI(MM?U^8;(EY95Z[,SB(HQ+A4=X&C:1-4N06>7ffD;,D[
^O8X4P#3&QQZMWT-X7P;_V-SG>2;H[ATH:V+d0(:JN;Ld>QZ8V95e4b#_bS97R\#
.S,HIXD).FB.^BYdc0>(+W3]NY5fQ&20/&49,Q4^T/5PTJK(b<.]6dUdc[O@\ZWG
>46.6DZ@^UUJ<?dWH7f[VB,b\+6YBC,#?g<\<NQ8D\Yd9(0]Q3<O_=1RFId2GF,C
;A[@?LE9WN):^CRQ,_[_>ffSTe(U+^]B&2CP1GTQN.<(H+Z#I?@+O<2[Z]<I2Q]F
N[IREI8L.0G2>CTQcc27J=8RHb)E-K4RO2C8/e9Y3FgP+J=X8gAQ)T+bS\(-&;I2
#;_/c:]S7?3cA-<FX^<G2U]\(F7N#4C32M;MZ<[P32\fU<dR]g1T)S2#^=g>6\TH
(N?8\&Cg+J=8SPKPF/C#WZGGCXG[/R1<aAI#aO^AB.#?-T:QU)b/-.)=&e83_JV9
TV<CcD49Z6_+8L@MA_#Y0#SS_OMLF2@_7H7CG8J&D6(N58C,0_N.0<PV5MIM:K7,
g3VV_;_0/8b&A-E^Vd4,LOS4NG40../G7MJQ98+7>V9G9UKQZM_QJ;J&)R08T>OD
bEW]f\_[f-[E</B5Z?C^=HM7#(5)@fDD46,bKbJ4dM,BAOWPE;W2a1^OFH0RWaIc
Wb/AfM6>Z9gPYF#9XW2Y0_,IVB[Fa1eA/d>ZET4aPY[[TG[>>#Y?Z(M.(9A1TEVB
EN>+EFHfV&?CO&<KbFK:(K#IL6f15H480/2+gT#6K;gQC>ACF_dLFHQEJ8FJ[HIE
45M[fBJ[C@53aId\>K6WWNQ(2N.0QK-BHJ+JcI:12f^1K-P3P)I:D]+,AUHQF_f)
\FM).XeLYbJ>Yf(,fW&<<g,6O0>d\:&52G_:6G2R+HKUC@d&4#bGKN1R=YD/B<=[
EV>D<,\,7[)1PB9;fQb96d:(^.OQK,>a\DO>X[[HCT@CM-<b+;E4?<2QS[B32KCM
L@=Ne=ge6^]C1^54:)&MdZ4CSaU=KHIDH.DSX^a]G<OdDYCH7;U1EdH3JgS4VaKT
^^SNJ=fNU.e;EdW?W-+0M;DMZ_6gV:TXf&W-Y+RMV?bb&Ob_W/b;e.deMg[&H8ER
(aT[KH-ED9NH9P)ObD@e;_c9aD&cFO)^4>=S3O2-T?4/gJgE;+;(65J&cg0J@Y<A
,4^-1+59\.&a]M?&=],J>J-E&,7KQWVGZffQb2VSH=I\56=0JFY)M6&f,.;YM[:8
e?\?LP:JJ=7>^B>FSZQ[WN/9:33MG69L;B+g<VVbRda:#W7CUOF2Hc)GGa[+C8c_
-89CgOP1^3K:D35d6gOS.cL)(g]+]P)FCHC-U+@>>&-H5Y90<ZM#5+=ROM41ARQW
BA.DGdgAW(+I3^T#WSJ+MGScE]5CfF\SH5Hb]ad/0SBRH#=:3P_>^1[,5ddPYYYE
U\F/.IU@YIOTdO8_R)XFQB4W25^>K;TH2>-6XS2f1,H14:gA35CJGW>)d=C>E)@_
gN^=KdeNIC:)[(]:<L@,A;Y36d_1Z[3KGYX>3eKX]BNEMA5W(a;VB^)A]T.I#A4<
g[_TBV^g_9XRM.N<6A8R^U+^75G7Ud&c+>.<YZN;],O-R]_,c7;\,dH,c\HUc]N&
_<9IQ>2M^/8dJZa-TH)+W?/CNd4\(C961Y>cC=-&CY7AXHU8LM6J9>K@)U+dgB7-
[^FQFReF?d01eGKcGPE#FN>8]54Q94gZ7N_4BQ//0EL6eO[]N,MCKePDeLSLg4PD
-aB&Ec74[_3[LZYA]0@)g>T>E)8Meg[9fD1Y2R+ZT8GaQGBMG\dI=+A+2e&^@d_O
@dF0IT60,HU\&[M#+K/4Rd01Q^@B@cgfX?JM>_,&:1DJ=8)Qcc3&)KDO398@a<]A
d:KP\1T^KAOODZU@3.B139^FJGW0H<;ZSX.-dW5YX>]4ga4OXgg\BQ3=+I2E?H-A
MA6b3\70d3g=<^9WJ?AZR0,fPbE=NN+[\M(Q6<+5P>&\.W-D1+0F7GQXWI=SWC9d
X8gbF807(:UC3Q2CU1#d#R^IEd4CP&<6a3_[V>G,NgC7?#N\M3[1:C._V;Ke9-+.
dLBAB/@M4TAJ/e<eW,N/LU5O26.7b]C_EA-_1PT,Va71,^A\PW#e5?<>4JN#Vc+1
PcfG3E\Se5VI;5YQFIdb;a,M3;UB\<Nc>_T2HG<CU[Y^FKR@363+DN^]X;K[+WUR
<V#Ma>IU,VP2TIJMYXcE@BP>>;,M;:TM>dc&-H9^YYHB40g__C07<&;2b5L:fGD6
B4YI??&^I\D&QQ1N3)D^b\0-?aQ.DO]NF8VF[?R<\>KRTNJT:?)9K0@fK2WIXM^g
dC^)8-<6cD[ZU[OV]c0#6@f\UgKPV)a#+eBRfI7/cCa1<;5T^LS(fM6-;&Yf0cKH
RBQX#cf(S_dUgda<O7@:FAS1(_K,(G?,H+AB-?9,]LOfC@6WU]Q;5OTJ@eCL:eO/
=SNaB>7(KL/b=5bZ==AN[YVP=Y)66/L9R5,[J=.)a5JKXVceNDF8P99WMcQg3B4Q
EO.PJTCG06P9>Y=+XE,fZ51V8,&e2I9/\<gD=-KeeQg[<9.YHG..J/;DW)Cg7BaH
,gEHa?KdeR<UfgGgRT2@Nc[C@9<YQ&9RZ4SJ]GQPN9SBd\&2eF-DYQ3FU&1QCa,g
UG)^#Y>@Q7.JMK2V^O=EA)eD_F0HF5KF,AA,(T+C/Gc])H0;YRDf_aKKP&g#>0NI
#Q/c]9^g5N2@7ZT6OH#1/b@+b/FaNT3HGZ&\^2^QTP@J#FF6#I/C9f=D>X-TJB;Y
MdB6<ge);17ZY8HeFHM.d.?)^W/0KUK7B7f3cS-beS0:&,5FP5Ld>(Bd2OC^R[)D
N<YTVX(<GW.E#46=DJYC]HB+RE[3U:AJ_]dTBSEZCG7,.(?ZZ(_cQ>cf,^R6NB9Y
8f4=^O3EW(\ZSPVT,Q0OfAD&NKfecKBB)77Q0/Q44FWgT)Oe7LBK/&6?N[0GcC5T
b.Q[(J\X?5IR3V\ON=O]Y.,EIg>G8W?&S\A^G?9g[)QeA;CB)20C/P6]7d>N0+Ac
WN71/F,387VERXI<a#..Oa44RSO3S2b<KF?4P04GZK-:EV<STB;52XNSP@\SX;DV
d;\#L9:&(SYK;=.#=IWY?(.-c(ZLEZYYYOBUOb^8>II6Ccf6P+b=LHg4>?O?:3f;
+>e/dK(G54Z\Q<6G+-<RbWZH492eKb&N@<Z=#VR8<3O6O)6V)=Y3^BBa3bI33c=<
I@243A.a\2;\=2a^?]gW1M>BOAB&C.O5;Vd?)2^eOS6Y]:U\ZE8;YP@KF;WDI=U6
+@CGJ;&b->T([d:E[]F-KB@,T00-gR+Q?5=>DOf(dMH4B@g/eL\78,AN4JC)WJ]2
geR\fQUKT;,N\(<WO4Ud);,+KPDATGR4IV]Z4-\^;fY5\J<;^#4]6NFSDV3(-FB.
@,]58+YR]^6^<C3B[[J1[MC\Ld,V;O=8[JSg-]):-&WIJ0f_H+/4Eg-U]bDN0]Dc
bf^\M4GKPGKG[d^V.a2&+b-]GV)8_ATcYPYa4LWZM8,C.b^,GcY6Q-?R/SeAY>/d
f,T)P:fOD=0Y+JCd;O0Ca4Q[;8.DYb^BI?2\G8,^a6]Zc>Z/[CgY\:M47adb@Ta.
(>9VXI#J^(]cGf4T]2[?&P/^4:05b]QOOFC(CN=TIacf=g&L;:@6QW9^4MM6N;12
RR+>3eCJ<M-bMML,9c2bUX2D-YP9Jf\J.gG#5/FTHFJ>I>#<)&^c8#AASd=QMMH]
X0)B+5VMU<I?B#d>GPHNR\UPD0TM)D??[?30Q>EA,d/cg3>.ZZ,^ATKb=g5O1]9>
aVR6+9ddX8<9D?eO&E3Fg)9cg6S)R\BGP#FgFG[X8e:7/3?,^,Y(B5?5eL0N,3RW
J9;M@XX0#GXbcUWBY)dcB=3O?])].Y0C4D3OBL1WF0JY-<>_/H,6,E4<&(bL0DZ;
7^IYdX+\(QIU8^eg5]8D]4(cf7)=DE3(K+SD0[9cO&eI<:3E=CBE7OS2CY#73O39
)P[>&9=Zg0bPF?2D1^Z7D13-O\I-[;1.B#-<HQJD3R6B[NEcf6]L&7B((Z#WG]&3
H&5NVGQ50SR[YL6:5/(XBY>b90BLWB21)GKD3_,A;B1WMUJYbRWII^TU>H>O1&O<
U2;764K:H?LJf6,DV[5VB5?bBE_87,WRdXe0@&Z_8[:LBQSE+?B53\<6WS[-Re]>
A+4@-I.[PQT[VQTc-45Kg)@HAPOWF@0dG(SN<\&B/(/aO1\+658;6FP:>adIdddQ
Ya9>AHaWf&;?-bbe.2,,:I?S/B3OR9CEgAfBYQ]ATTQSMe@b?1PE3AW7?I/]=Gfc
AHDQG=g^AM:\1SNF(5fK;;,LVZFaaIPX#9BN0]5232.V>9WB)g85<6#JO9P]@5FN
>QP.FXcbFB6QPYYX-\Y?>E(^\JVVVW\L1APKZ<=Sg2..E-E;CV;HP0\dG80&FOXS
.^GV\]_B680@;gA.f66EM-X9#3/N92K@ER7S<8@8,<(J,Z>]bF:[=aBcgbPR-OAP
d[GP7;c)aU4ALd-?7(1IJ5JEcQ2\YgYCN2[\7L.-gYB-:@UC<P8FEH08@^F=cH0(
/9J#(]4EaVB:c1-MSO98UeCWe2RX=936RcFH&9A14D&33R3\((&)Y#Z=E4,8>LLW
<AFVcf\g.S@-WaI\R8dL\Pg&=V8&&dHe58,JRSf)Hf7=03=gX+Q,;4ff30d+^LS4
e)Z)A7be0f]g,QaRb(TPVW\aELfRB0;c1;Q;3G@2QPO8@E4c./g/(GJ\[2XBG/+G
bI(<(F#;SD0(R<KNLT^W]UZ/\JLE#HK&QU8QLYE/,5IQ#@:3C&CbfWJOU9^/N^Sf
=-,eK:c7\=6N\9b(2JPIag))EX>a([[\,0E#+g)=\:\?NbNHEgZH0-2fA_N-@L6B
ANV]YINM)(BK(ZLDPd7QC64?B(W1/0:0.9e=L\45D#,Ke4L0Q_[.LdGL_I^Wa>)Y
OCBdg=#U9:CGODH)R2A)4:))/R\.+dBQ^_Odf@3C7;O=9,?C_)Sc+ERP+I_9XIPS
(KJ0C?efCM7W;7&Q:N^d:RRI)g5VeV]6:d_[4+9+=GTc<N6OTXVGWJeUF)2e(?Y6
a9#[FQHQRLS__2+@accLH1F\,4:DKDX,[V\6V@NJ,=&)2E>X3:C+51]Z4b7#]GeB
c2c(Y(b@Z/f6-)f#_A;D9^34d[<4<.#-:^3N_[R,Q5bGGSQ1Je)bMfAcW#C,F?L;
cSYNY0Y7BAE#@RfO&</dVT+U-26)?]<V6^CA@J8[<:#f9XO[=<ZT0K#X9:3fKNaA
bN+)f)-OZT[H9MJJY8SMPV\QBFAa0#U:3MA/^fV_;A=Rd,.\,>BJ7A^&)(<cUVN)
O<cR&OB=H@9^ETcZNI:)/D4W+&E29dHI89)SS&_]BQ):d\gF@^0(5Tb>?>\9ZfY\
0WIf\40[V]e=cX-\(>>NG1MZdZdXRXc+KA/X<D@&/&[.aJD6/a_-;WVB1<S+==bW
OCgXA]MXPgHEZaE<Y+>Z;fXgEaB@CX.:]YN914L6#CcdO_fYbNEN-RQJT?c>aB/@
LM6@BDJ/X=MTT.UXYNOKW[FE>+:1K1D>+S_<2V,DO4B?VF]VN93&,;W<N].-dNQ:
[DT,U#T6d,f-=5NEN@c4b=1JOG=SMX^R\fQQ19W1.RCeZT-K48N>++<UU_+,U>PN
P6(9,VTE.;Q]\f_8]I?R<e>D61.bH1N2#DMEGF(?A@+8=:B<P=-NS.6;8d7FSUI/
GT=/eUJON(]4d2H04-5SY@338-19(G>PB2&UXMH]U[D<Q.J8G\GeQ-^eZ<T7T9+U
C&<F#&7SK0)EI;[1C6U0&J>Hd^WCaE_XANaL7JR;,E)gD5AM334>Y+OA_A=P:4:<
V.EWW954LO]BB7>)Xb30J]AM\bWC1g=T/&E:)C#/3&e19WNd?^88JO4?caOc;e<7
2Z2/;@Q1U>H#\JH9R<VI14<DGc_Y07?#-XP3)0fA3f?7fd#9[a[-/9&Y3bXW\B2R
=a&TgSO#)f[^WQ1I^:T44Za)F<VZBR_.\@)5B&@6NL5J(J,[fUZP?BF]a1&+O-HI
YFOZ8c#_^[41/JP^#5gU-+_1?Y90DR2P#7Q&I+MY>9c3,)UgI:F0(bX2c.3C55B#
UA/N6]BCb@CPf\&LW>L,?B1WOd/14R#[/IDPSN0R4Z>BE_\P_EH8dRb-fTAb7KOg
WQQD8QW13M:BGeT1PNZ-A?C-B4?;V.U=^C?(6WYg;T<.>E^(<R]HefX4-=U..\/d
PX=S7c0Z-2eg[BF1,0EKaU4.f4HD6?cK8KO);A+E2ZMH0HECQ[RG5/F:KA9ID/VA
)Y4O#8;a=G:&dI)4]Gb:P1MQQ_=&;+=1NEBVG:@B45=&-^1X-aQQ9A_JJQL.g+O.
_SD,Db19ZE[9(3Y&G)eS#0VWC1&6/SZ\.QT76YgRK&MU53F#R6Ea91<PFP&6eYNM
dMN,0[,AC))?V9aFZ=@+_3;O@BR^X374L)-JO.5HCH59W?eH1/,6dFH9<1Z#RfVb
G[>+87Td;5[]CPLD&50#5WOf]8HWd/F)WJ8QA-+ECcJ#R<?UN.L1V-bR4\1/4>A3
2Tc+b)OX-7Qd-2Y86KY4e#8HAC9QA=2N_:TdN3G(3Q-eW29XIa?;;Y[/?X.:aBMd
AS8Qca23Z6@dc(WFY[Z/ZO.H]DOA-W/I:@^X>[UO5:(EcE02a76NY?[@693H3DSe
:3]GN+gdYP1V5\S8D0,eT](8SJZ3gU454.fH2CH4K((RGI+G]Q;2N^Y1_Y_Ba>d5
)MVCDJ_4Da+K)]+9Xg_\d/:EZ4PcH#.YV[ZY3<A?;\[F1QBJ?,a;c.gJ__#4N>?.
c^Qe89>,[1-S+d-?]O740K.<Af^S1e-\>e&5OHKGAe\8<(T-L@?Q#cJdUHB<WYdF
ec8Hf@^eEEVILM#@)N2SbR/36V:NTgV^b==9?W(^-0MS\1>Y<4H_a9N^LYT&&D/3
f:1SW.+YC3Q;[(@cH>@cLfHR/5B(03JOVV3>)X=@U5G@,??1QP,]5YY^I^[;<L/2
2BH\/C43H#d\(1E^_+S8<ZE?VQ)I0@]#89N=7;4/1a?S,UKKV?+(b0D4-9DB@7c)
Y8O@DY[S\]6YCV/@c@#L1fOTV+,Vf4BPgQ<WW,/@U6VGXA@4O\X-9WCJ=2:dXK);
fEC4:9S7fTA4GH+9?(#:@XYY3OgD26OJHXef>HIE^=[Wa1JaEgV6YRL:9FN.A:UB
;Qe#8f__=SP@D7>+BJ[@;gd(FV83#1^LR5((&CT.bPBT\LML@8/\J.^V+G:&DE+X
c8B=83V@ZBZ9G8K[BdEWXR,R59Y\9L,B)M)7.\4<GOFP=DM_,9X^-EVcbJT&8b\+
SW?;Y=E,]d8C@VM;:9>;/dXQc&U>P;8[NYO_2#gG.W8+c&2AICFK_>9M2Z&C,A1g
NQ5_X^_DdZ/R3f<LTDHDR2-KW.TV:;<Ya2>@/@WJA+-gK&W+c)K/4?W[f@8III=2
FN[\&V:8F+]T[ZNPP[?H475EU\=&E\K0##X#NI,/gPQ(]bfeSV2N4dZDeQOa8@.?
M9Z<g^IF-6f^cL+QZR=08=STEF_4DUUK=)E2NAB^A;KRgROc6\2#d(9<>V3#L>&E
P70M-Sdf^9\W;RT9KN)\RB9/.C//>g+&0Ab\(U,NOda7)S)1.PP3N&(JdeX<c7TS
(3W6P:H8_;#,H#Y;R)85U7,^A/V>QebfbGcFg@F<YM)(.D=F=9L<G.ML\W#MfG4H
YM>R&=cHJ7ZBB3Y7/?TQPCN^R[-D\LJ;d#:f3^2?ZM2)8#V&9eMeL?eV#V[YM_2V
F<)I_S@ZI4BX26.FP=KXDDN;?O.]g76C_3fIM#A&R/ReA2[1bI7&(+F^W30[3]\N
TbUB4LMO\4K-&PXR4)D?dJSg8790fEg5V>>g<F6+aef?8C^41:]g-3=.)>[cVL9,
YGX@1KUGdW0/LGT>e7+T+1.CRgTDf;1W80(.YaF;/7HDKOL[2S[O1fWE2Uf+71FB
^MLQC()0>(]2Y)LJb98KfYFIOQ@\MXd_fARI8N1=Y7LYU^d_C>ICY,3[_MBI0^>2
]aBPCTBW2I8K[&X)=cM:)L1HT40EKJU2^-J6N);60LP1\[</[4^Q?>d,0;2[<C8V
,?EG1d=F\\(;JQOMN08-f:&W=>Y5QIT&ZS79<LNTB:PeKK]@@ET:fQJ8W-g8#F)0
#[:(9F=#P#-=fZgb]f1Y(M(3,:JCL68CZGb:@Se#HT@C9\UaA<ALOI0Rd6NO#?f[
V>MY:O9B+/E_7A)I(fS]d;PaUdEX2KX+R=5?@6>MA8VEZ9LbJY:DB-4#2+540CP&
H5+X;e9T?^SJ^,QP>f^_0>:(.);b)#88a:\>8^A#+I2H4]cTg[9b#ffLS.D3)+FW
W9&9>g;g\M<(7-P+f5\_f8(5eVOJU.f829;E+9:HJd@d=Y>&]N_2JD1W5e?[@.6[
+)e)]K1KQffC#Hd;XK]865P5,J^_eKUWC&81b7d/)#/,,T1K]<XcJGL?e3?^GCDG
(Nd>[<M(>G>=dHA3(>T<K^J>6<f&1MN1LPSMbGWUfYDGaAF@_RT)50EE7g</SA-[
T:(_CQfH)W5P9KZ#TN1=gZET&6VR6NB71KKEG\VY):6d78)J))2=e(MOQSV=&/Cc
FC2<CLSWeVAe9_IDI>T\Q]>+W3<H6bE^C=@D@WKE&c95+EPdScO4gK]F6=7LX?(M
7d@DT3QC10CSb[KH<1;53?PQ<B+-&Y6cP1H&)(H&QJQ0cG561O12,(-JMg&7K0U3
4<\2QFT1_DK>JQ3_2.S)#-D-@^(1H_eb30P,.L6B\DMS^4W^,&&G9Qb8LPa7B)MI
XLI#g1/F(^>C4;A=O9WLO[4QbKQbd1B3?X&R9F,;[,R&+K#8VXEUT)@36^-6U7bL
JN5EO\M^AH7[YW1_<g2f/W0-<Y0g/-YfEG0<ETA46@bGc_UR\)M?]7&B?\e;G^&P
>\P(OOPTMBN],+Z4H(bSVHWA_g&J+<,_8TWLeG]U6U\;AM;.0U4:^g;e0]dgK82-
:F<OO7XT@Bcc;02e[9?(@I-=CC.Kd1^Y5YfdL&1IA5LNHIcMSBG&]@0K=.cK^SfZ
_Z[2&8--\VI:WE)?Q;#;QGc;L4LG6Q+g^BM;I>SZ.Ff+gUL;T42g\_+4J=>(RT&\
;^-IPYE\05X/fa4467a>/@e?OF\0F_?+-=A031V=G;&PP+=a;)CXB^-A?^#g1d6.
g@HEN;V];QROX\LgSG?H9bW16QIRM;INF6aaBJ=.:T+bDJ,4^X4eO2H8E,_F[XRf
F6Je3S=S)+ZYV>LVVTV6(^#HL,]]/aL#RcQ-1-PM^/TKe@9M^MVfUD:gKD[XO_\J
)M49<ea6FO5gD]cBZ#7)UR799Hddca6U((FI7.Z+8KN?90C;[TY\XOG:64eRY<0#
H:aNT.Pc,T+X;2W_g86)F7g.a>&B-HMGQJ)>R</S9\WDEM#(1)=eK&ZB6[AXdL.:
GP[^INDbLO+IJ9(^]b\g)A=3N0CZY2fOP[Ja6@(]g3aM=6_L0?=[G3?:,H5:;FKA
)ReA_8).X#L3/X)G^JL,HH[edZEgS>X?5]MKTMMPXN:4[O39-EY@G.a)SddfLW(7
1(/V2b3f9e[&5J0_U)NN7cBaF6Z_DaKS]a4.a9HH3XAK,3Jf98+A4-Te?O]-PB>J
C/O[30Q=;\]Pg]f/7SI5IWBA.]<1,B0YbZ/A]O#W6OP+IZ,FVBC(_(BJDC(=1/:B
gFX<?IK(bA4AEd:&)L?ENK+cfL2e[(YHEN<&\)g810#6f7cO4]a1g=8+5CIL?@?d
^,:]U)cN@S]NHK/HG1)K]V^&b2XH;@[M<X.L-@#68[C.[)Z=PYV/YT&TY:XP9B3;
N(W-9+gT5^g3=cW5B5IEG874e(cJERGKG[G6;CSWV1TWSeWW5(@&fZU>_:LfUdQ(
;:eJEEb,7fH-?_GcS9]/ORT5?Sab>UeZ3,XGYWGXXZL;Q16G?)A19_c5PIb7EGe9
[,0ZNQ&fgZ\;UG]d+NP\2b2J(1/dAVCS\?9W@37O2f2U)5P:F?XIP^OE_?8GH>?&
ASVW82KM;O65\#09UM)=)f4YS\g3@F&3)IW.W(,Q58Ob?\(LNXH>0F>T+Z:b&g\d
<0)0,TG15@TW?GYV6O\?0_MQdTNFQdReV,MR-bW()#5MN]R<eA>8U64IV8?f,fM\
X;eTXR,J(fXWg)@_#.IYPD/B),0/N9-.M#F,DYcD=GDC;Ic#NM#fW8D4W>U(7NM#
gP(=7g/f8:c3()I;F>LHgX^ARL[fZRLN3IBCWRc>D3G<H2,9?J,_cEg8baQ2cH1D
VTID_8+\(RTBFAP@O;Xfd,<>/(6+D\E[X]Ha6Q4;E_b\D/JRZ<GFI4I]E-K^[77M
/1Z\>;ZD-/(?a1bOfN\@>d\Qf9d(^(RMNPM)?HUDIRg/ee<P36XUWRJ_RY7aAUH#
bbg>R@6#11D_2T=G#I+KXKW6I3]M>NC[7VNUTObF1.?9=MCP7?EH(W&JbIa>5SQ4
N@a^8:&^>7L/LX=U]L<gRGgB=?\WdgN.fAf2B2A<V6-fQJ.1cdV8G9DD/V0V=f?,
,A_I=WH[TYK2bg3WVM\1]3)Q1&J1\]V,L_K]T+@GBOX(.DFd4X+<UC^V;<T@Mg7V
gT?dLaT9FM7VabNfXW)]eUG@<>3Y9NO:Z59f-)^Ub^\J[&_Z,[2RS,#)^S4\=Uec
D[Q_5Te+Q5QcU<5gRb5CWO4SQ(+)OfI3FGG\&9A&U2(]UN9V+<4KB+=P_5=6=O5S
_U8#Ha29ME#@)R\D67K1VJ8gegG:J6.(MN#Q#T&?K9c^)Ab;-\)+Y&?MP5&&gTLT
C/OcZ4&b>A4OQ?VRP?C8<^.g(g-bUB:CBdP+Kg[N[+OEeJLN=OQ[^SbABf14dT3H
.SUNe\N.DNIaDOT^TLFR,dcLCWg?[MIfBFfZ(<A&Z]+LU4YYUZJ)1S+R5Ie.+;5c
CT.Z4N-KM@YV#=(f&I8f9DW=/8g<?&9RJ<Y7J0)?]O@EC[09H:5fcfQaFJfS2TJY
]A_FUX36Ga/gA@NddaIF8\/_/I^b,]_-@e;gB92AP)9e.S\gZ)b;U31^V&:/CdFb
-/HFWS)E=\T8OKH)M[d92)8:X@<X7OgHN;c,R/3DSTV:2+DQM/U6(),A1@@7Cd3,
I.)QZK#9:-?M)@B@:LKAe^MSbMDNMB;YD[?V_B6]DNYZET-?E_5,^/;_8:7:ZX4g
eZU0b3I3&bHS5^++79&<c/Y09N9Y8a41(CT.#^5[U^Fg2QT/LF0=9^E3:]e2G)@f
[RLgX@32_X28C&YSU#=d8)L5RG;M;.+UOF@_FB/\dO>Z9K\SYba?.dH4/--38C0N
9,1[aL_0/G+W=/_YG2.,bQ4)]+86.T0UQZ,9eU5FZX/K(aY(VcX&b(fY;gZ&T@/:
<:.gI?EHa.L.FK<\b055bF5C4&JST3YI4-\Y44)/d?R5XRGC2d127D^]B>3@Q0^=
40)5@39+M^@LS&?DZP58c-@MO_UYQ>c1>,R2W3;90=2W43a22BFfGH^P+7<WVUg>
X01g9B51J;5?eZFS-,<3@Q]bAg_AT<^-=LPcBW,CF39_9JbVIKZRRRH,WX\?MUIG
F6d:B7dVON9E[VF3<HZ+:6IU>14c[HRGG61C^ZQIPHaZ+0HLdf+@>Q=(a_XD(C/\
D#S^<P+2_f80C=U,BN92f?@:\Z=g6PS@_M7__11((\^2>T@\ZI=Fa2=.?YR]MfS+
A)-E[J@_47Q1LE1;ZfCZ(,V<FT?91L-FN5S798CZS?aI6TQ5,QP7--M=);^e^D?<
3,#)[:/01Q++#F-K.e_Gc=GML_<AbF8)c0XCAB/eLbC5L>E/ZaR-FWN\d[O,KK)>
BRbO[Y6UL4)CTba]H7BED<cB:H1MeC5E#F\([57Z@32-I3_IfW;G=.CXd:a3)e\G
OPaYC9(G;BPBU#NQa3)eXV]3XIbDE[72.LK[>cdI-a;:K#;J?;Dg.c,0L[4H:39E
=gaU^>E3AI82Tf8L&5PV<TQG4b?900VfeH1f)SEcH)QVbK#E:[9/7A1K)OM41eJR
<dD@IC.4M;aNI68#NV@Ug]@=M-/-(;Zc2GA[9YT?J#f/9gA:,><6]P><?@/C#VZY
Qa;S>8@(PCF\,2X&beC/@CKEKT5D^I6g,F1E&P-ZOdeS@#Vb^H?cOE>&>cCS+V5-
K3(RaM#9,67\3V1TQFHF+Y7KS]9Q-2[KL\GE6&_]>QL+VcJ0(-(2PgJ-5&X5N^B8
Z;^Lc7eR7D7fA>HX=9PYHa7c)CNc,2)>,Z&B-0KM]-eaC7dWbc2G6Bc3MSc+_f)@
&d-8WaE;&P9;F(SU_2K..@e\&EV4Z\K_=R)226N^C55DT<aY_A-O44I;<DWQ/d3\
G:?#5\9&\1UP_6E.0G:;eVN)agEWD+^E5)OSCO]<<ARDC[G]-8YE>5P^1C-MM6Ed
=[EE^S0eHa_A&/<,OV#QTW2#eTJ3T<S:=E+-QR,4g--#fQ+YS6#B4H4TQ\V(Haf&
AQP?d5D+:79,fK.>>gMdRY/JM(,L7E0:#4,J97Gd(T@(&DDS5MVQ0)MJf_]WQb,<
-U0]]&?>ZZ@WQY;M<1(4I^Cf-8fXa-G<+a)YVG;dN9,3L<2G5A\3KAQD43CC3;^+
e4^3GJH\)@V2Lc&cR@N2[1U\/)2b:D6/B45B@YFScB3LGE?UL/YG0,\a,RN@07EI
cf@cTTCWQ.PV99FU<_L_UX6MI->H[]<AF_5<D0?8VXU1a_U31WH+dMRQb.,W);[M
QV4\OD+JeC>NFRPJc>::eGNK&^6YC=O5><>@GI<a=7+,C&HA;32P3#=Ac_cbQ4>B
GWEPFR72?TJfU]J3dKT[IF)?@-()V7)BLf#L_7/gL]8bX&YL:9_W6#?d#O\TX;@T
0[KH^=^+_>Y3<FgJED+cGAbYR4af0Y>Lf1?4U0AePX16JbZ)GZ7Hb>N\VDaE:77,
fF,U\IYaeA.>?WSDX4U(bfPc]3.4W?[a4g,6CgYH2?F1=,6d=ga:)6geJf0J(a>g
/dPT&DbNX9HaW_?1DQ>B)3W,,MCED6d)[UY<c.FBIL[/2647:6YeDDBJ=K#O>60#
B;V0TH#W_TP^a&PDAITg7>).@TZ15]4(\DG^LM?#7((E>^F474WE<IR=4B_&^ZFa
IZU=c?3V\&.S+9HHb;V#XKZO1S#DB^^7?[3@^50CST3QZ]f>R3TY^TMRZaL;HZMX
<EAWA7#_(K12X<^WI6ZS6ZRT9P^S/F)EW?Ga5Gf]Z<F,;a6N<]SZC2M;MeMcA:>b
LPKGU)P3P>&(7aT?L09+8K.?^7gBaA-(6)[J=3XfVdeKI>C&_\)_b<CR7(:a;a-b
(@KcdJ,V.H<XQFa<DB_SZUK[1G7/fIc/K4=]^A4L-;cUaO46;GL4LR[@S+VIT4c6
Q0:M24)X3JAW_\B.?/ZA[S#^FJ/PA@:F.N<Q_Y^a41K6T@2E]5TD\[FL,\WOXeNV
,(Od\SafgG+L1a=87PK4fDPY[/JT0d0A+4__FJGg?&^/<&gJ=LgUMY4e+d3=M3d-
+>W\-9#\^#YO_?BD]SWT+Z>5\Y_;>RLIPP,>I@a[/_3F57?.UCBEg]5>(BU61f>6
.1b,Ta)XZ(-A:D=(?c=]A/P_I^b9JAVOMDAC.QS3+gBEM<2]g9DXDD.)Z+&@^P[X
FGPeS#Oaa7\&87NG&8a&ONbc89G2fY,8[1dd.a8c=VZ[73@U\Y32Z9B4[[)KF[4?
_6+HA9D>R.1KKNeC<:+9A-T#+Q&KcNX,989Cd^g3GB?:^S1Lg^;5a3(MTZ@4PeXK
c)=M:ZVRNDYd(/9bKBVV\W#^>\2]\;FSb](G=T^<L2VUS05aDY4:(C=]<DRMJU_S
TI[IE)^M#_^+(K>CaW=Q-CXOP662Gf_XG/4d8LgP9Q2:F87,f/gI>H)PE&,eKeBD
U(E#9Y].TLP<Yb5ZKc)7aCB.&J)6X88+)Ye(cCUY2b>3[L5_[Y0]#9_fN+S:\I2B
afg&UFLO+V3+^XbGWWEfNKWK@M)R/G6._;daJF_\H8gA7P.F8ZZV7Y;1XI.d^(3@
.0HeI_A<BgFgVPS#/+>1f\_8c0]E9b@(@7#M&bFYC>S/.?8WO?3HGCFLT5DV(&91
E0]#W9/gc:\7WV&AKgS&EO7(1Kf30H+DZBF@HMXe&M/0f(K+FbC-4_NK]&)O+QC:
T0HHDfJ>)C780JXf7[G?;+US47(;.I;F[Jegbc&94<JE:H_L6[cf;G6_2U(]N6<&
H[86QX5H/7B/.+G6J[/Eg\cXcRH3B^ZeTD-cOcP7(;6+3Q.T,767C0JaA_.ZK294
@3aIg-EYJAK_8ZUdYDTNaYVY2:^T[]V-Mg76FFZBOcQ.6)c>;J3Pc\0IcFQI8G89
\g6aK6fQ&)^=_\HDf1g4fSFCS[.Bb3C?SCG6VC3ED6S/4A,C<;KL=]X#ZD)Q?Q#,
b.JK&9fW+31^cO8[M<@RA1,T;EQVG\RSIZ?3[#/DZ_;[]-,0b[>dQG;gCK8bG>.&
#eYRe[-=M_0O#1gUYY>M65C><AeDRL2dAF(82KZ2J@e?_&]AVK;DEG=HDVP#74[d
-=.DOH&4?aEI2\a6T0dF?Ja54Ra/)XWUW;?aPY^.46A(21&,C17>D&@)LbHAJQDK
8Z0=L/)TWd,3F7?S=aWM3W^O,E&WaZ1Q_BEQ-L05de>Je@K[8N;MI\K3(WK^gJBG
_-.K_b@2_^7+J,5A<0a;TZc\BWc]\515c)3a])7?9J]HK]L\)?VQ6L-KEIe\Z]4[
<8(0&1SUCL-a.:0dY59d&cCaQ\^&<LLB],EQV62]_G4X#O:91<&,B5^QBW3<VQXT
@bSE9#R<_:1:9fEP(@?+B599A]U:S5)(CM:cf<TUdU..-bD;)R7[8RLT;LV14^Wf
J#-,?J?CHHIU<Tb^dg]NMcJcO(]WO\]LJ#MB,:FILW+#agW+3MV9,A9d_CMdQ>3&
P2O?I[dX=GQL+2>_I6XI>X_G+F_/f)B-V/ScA6RT>S>[)AW6g=CSI8^6PL9-V1>A
G-3DBN1DY#e1CJ0,>H0[UXGF&(N3)]1(O6F5C9G+e5OHDbDdQRI\WOU-Z1UV\)G>
3@JZ4^8FgEd0HFVSIGEcUJUK1:0Q9.+G&:I]=,5QQDb>D(62OL?RWAfB6gR:R8BY
G&9d,<2G=QN+0LHW\5g=SSV5=8d5_fZXORDe6MJ@44S5c@0BO<N)_,eW;Sg0L3I>
gKB<D.gT>[W_IBTEeYbR]O/,eR5U-H4_0S?S0e+1(@76)NCRG_-cJ/?D)QUeABgO
TS_,_4]V8g)0Q@[AF)\Z5((LRZD29G&MWVZ@NY?BR?06)8fDd-)9\Y#=QRB.L5E\
6H_4[61VX:0UG4&H@BX:&G3=GGe:9]4,U-04&+IHcCNcX(FdP>9XDUWFXgY?S7_Y
)2b)/6B\T]Q4+,P>0-C[^g_bJ83]_.8bM5<aHW1/P@dD(/Y)QX#6^EX3W8L+DHg.
G=fRZgO3-79]E[3>]Oe.O^K/d_=.(Ta1He>(>R4?)T\=Z)Xe:bXDFNeC?-NX\N#^
fIAAP[6_MCJT4Be^(K#5/W\T[M2M-SRGKYS;WUP34UDcTZc>BX8<)C1:35UUOC]E
6WJJH,C2&TWP][V.>4Gb969@ZdS<SNAV+Te?b50S_;.bMSK((,U1RN_0Td#.,&D_
R;,ERZ,L/X<-Z[]@)fdJ>KZ:PB/^fJd:W?Ke;D7NSHX>4.gHG.K,YMCZH<HNcMS4
eU>4cR:#&NU4^[2U#BAc2FW.(X/]a]9@K4J6JC;V+?K7B0)7+_ER)83gc+G)QVV]
7+MP,]MB+QJUS_HKIAGDgB69Q.17TT,)RF\F0W:JM5Ucb30]XSG7(=/0/S;NaSBa
7BfSN3U4(Z/;0V0U:P+NMR,6#Z_TX[AN7FF=S1)Sa]E)c)?YT+a1JRJ+<b#b=Kb;
4#;]DZ54JFVc93.M?eg?<V\UeW1X3)HbaQ3a&bOgEJ#OfgeE4Q4b((2Y<^L6>.ZN
>RWQ1TD1J&DAPWd&Q@ZTgIJKMQRFUT#7.bXWgIE._@URC&_M:dJFW&??)RVZY+\E
g34T0&:5G;8.9MXKeC0Fb9A]YQ&N8aMHOMN]c]eS0EXBGFT>0TY3,Y_?4TZI)SSQ
F_FH@g3T+)Pc=bUP?Y#[Q(>M1TH4N-6GH^2(4O[C3Z,VP2VCS6F;5Z3Q_Vg#_3Kb
EH/GY@365=(U_/PN9KVfH.3C+f,d7.>Eg6\(WQ:KOGdA/MKcLQ0_SB+1+G&=KGfO
IS]+(E(@;GT?5?]HK/c0/eRV4X>21L3CfgXPAX1>8E/,_N0ZJ:0DRQ)NO4:1)RcW
L<V0D38,dBK^NGaQ6<1J+JaFN5KH/0,X4YW_N/Z;X.KJYf)A:3=-I<Idb^&3U7Pe
4fF;P.GI9B9=W4b<3:,5:dZEab[6#bNR[A.9\Wd0_c/E+S71QKDJ?-=BLI8.KB;C
I;fWLND^@;6T7T#62fVM,f&^2#T,\&2WX=-Z1TG)Ne,NG],93fQ^R4@2K)E?\8UC
N]Y09SZ@/d<4f\W&6[4<H_3>S<eQ;dC=D(:8HATE(<KUPEI/_KZ=e<&LRReI9E3@
QKgRXP[U@U)6U<aBe>&EN<57PaHU957fUH^4Fc@:XU;a#YC_8DNe]Z4P^GAZZ?_C
,VS6&:^gBZB#:3K_P0AYSL.EJRN=E;SCZ7+Z_EXQ&;?.8SP.8[\_eBZ9>_;VX_8?
>#@WFgB4YO4JeK.\Ka<I^G4fC7M[EZ68SaNWGPN,1,?I5V(RL9McUVSF\>@=.8P1
M3A&IY_2M)a+d4J972;11OKXNDb;:4::U,Q7;DQgN0I#7;a>?-;E(R7>])fWf(?R
?A/0^:_M+@/>>,HR]K/,DJgaTMNIARX_Pg()e6)<:/g;J.>3R<X97R2(W#O,S8BW
/A9>?HgX4_/d.aH46FeG?#_B.CaK^(YM@45,I[b0JDdTSSM2cO9HZ=Q-0UEYf3^4
4f>+Ua_@.&AIAfTg:NOO6b?9@4#1TURWaFP/<EN/I;DJ]1cOI#DDEV87P>@M,#=?
DDX)/UXb]La[]?KeBY2^\^&SS-?VIAEWe>PN<)-M)6?X?4DSgK3DIcUW+CbB]2d^
Pb_G:+4FDX\0^@PJ&2IOV+@f829/Bd/a6.Q?I>HPg>_7@_gP-[aU[-H+aT8REINQ
4&S>,M,IEd^K.);GDPTUFXI+?,WScIT;.NgV,c([)T3_aI=+35&C?<d_Z=f?(cg3
bRW<6;RcXCU@56?2P/Vb,S:gMG-2YGYV\87D;b\3K[#G#\VE1-B-+G,?[FQP_:S-
#><HYJ9c@e54I7/&]RE?C?TY7Y]_NZ(4afcAQ8J//;HZ@02<XVg\+-BU:[#-O>5d
)4#R41d(P8XADBaF41<XE)>cW)E>/D^0C2AJ[F+]9\G]X:b3X^8ZNUgM69Sa4:dF
EV_>3/0#bGY_L4F>3X,#K:=A:O(;H-L85?]>0Pcbf@3WN5M;2+Oc&GDS8>:dMgO7
ZI625NPJ&UMaM\XZd<g\I(cR4]&>B377AF7<a8K4c<aB(X5e?9F]S[91L2QVQ2:>
V;&4X6X4Mde(fPZcbe<IWP#[>LFFUHKZ0+1\2bLaX>J,AgR[?P=dfNVcXd1Y]^FQ
X4]bWD:R7P],g1<C>:P7D;)X)g&-EU.WDB7F^bf6V]g(14^A#g4)=5,)&Z(BI5Q7
_JUK86BYdX.f)W+YTOA#7NFL4f@2cVAZWJ-1c4FU[/0RaC#Fe(M@7#eXc+_N]35B
IQ3),]DR)^JKaSFP/f:@Qf<_1I@ETUg>-KeTE1D-3LIUMBFQaO.eeIMOQKEb8Vf(
8)(Z7:dJeS:5X,JfVO_DZgKHcEA00^gG/1.&J/H2dNPCg+J9^QEUZE_6:>[Q/XB=
FR\aRDH6]6RDP0/51Cbe?P5@HE92JcJ9K]&I@a),3P_Q-QNb/W\D_e3d2U+LcfQK
XA)CQIN5_2[RI?+9IeS>,AC49bdK[9S+c-IJBeg4gVJ25H]Da=1:K;K@Y5;>41#<
7O.gNcCea?eE)EW-O=:ZE]fI1C,(1b87B-EBBb.&5eFT<e6fI7F95Y4E38]XMRef
:Q1:c3:T2(N,DM]SAC\6BIVfHDgD)]ICLdf).^?TGVCZa<5#ZCb,+#EE/#.T.]H)
W[=[MK_FI5\AXZ5.fYDDQ878/+\.E<4Q.9?E:gY<IIB7PXQPFgbFB&W(?HDH99U8
BdU3/SOaKD.:b>-JJ?YC)-NHFeS\fHO+^_ATBOQPR]Caed12fe6?f=A^;/S\E10F
R-gHY<#J)GGTI#W2^HDb(8[4VTY\&D9/437M(((PKQg2?AG2VNNWXLE1g@UBHA[D
g.1.c2Z9L[2--eJHQdD@_Oe<T15bJe7STaN3F(d7;a\^;3;KBCO-J&<@eH.>YWL?
:3@e&<K-0>20?VeQ1ODH#\6@bFD1VC>XdgEFg(PgKPI/&cP<VU-Y+02[fRH59MF:
9GWCXX7I+@,2cQ+Y8C41P1=dO^a7XK3CR192Q4.5e9AP#8-Be;5_AZEc34)^Oc+]
LYH0ZJ]3dd:a-,#HA^8_@2&R+fI2#R),IFAF&g/4C@]+Fb[]P,>WU:G?1Ia)b,@L
O5XWM)OW=DLT7Cd6X)2I.-V]ITfPd\AJHW8Y()Ld.EIY+c50(V:KHg^9Q@?6C7@N
5eQSf6C>H#g3bVF#9XQKO?_=@3DL:acJQFaPSIN3IQ8VR((A?0)[BH=]D6YRVKR=
,VS+NT5b?XP-^]1EN+(+5c>Na&eeZU\G]1ZC[L-^WCWU_Q9,YIa>ZT>@9@M?W.25
Y)\9@?\V)SZ8:LdWZ-E2\?W]#(YeKP-Sf\1M(<SCSDZQ?6W=1&#&MH]O^:eUX25\
NG/Aa=_ZDF_+;\1M;7X.,M&;+=G<[?R[7?X&6AR=&?P9RNS6<>\Ge-ZG2S<J5WR_
+A5f9()e?De9>TB]bKMLggV-NFb9(BSDF0Z=H>ORTa6YLVYM,1<&SN0e<-7CV6;[
ICNOQQYeLdM:E[3[XTaDC85POG_V988VTVB&21M(Q28X5:XYDd&##P;bIY<0I2S^
dd)^ZSfO&W+f5g\Ae87\EM@WL80JG=\4:2CQC(DBNGS^gb]NbJ8?KBQ;[M?84?4K
ZYE7P)&>R0bM#]\XT<8Ve.HD0?7AP3V<J#LBgXVA[/_A8K)f&,L@cgHc,-11]A7_
6:G)fQdONIZK41]V0LA]QEa/D8Y-:(AN(0QV0b7fQAC10>R-eQY_Sg,NR_;3D9YS
#\?YI72b.F(UH#M=B-,#dGU2IG--D4RM3ePOAV:P&XC=W^YH[TeQ8KPIg;/SWNZ)
07<(^fZZOf?FU^[NQ_a^C2;OO-Z<-5#KD2R@#J_EP\UZE];Z02[9_\Pc[>_\gHdF
:87]D;,(\CB,K?89eFKPV;7aZ[G]f,3/V?Z_NR-df+BKaWM-H8#AA]LTKO=K&6_e
:3GZ-,WN+(>K.>G18QSf1?V#LJVUAW?9F4^OC?D+XYc;L-&0\DOXd,:PLO0K1W2J
B.O7g>P0TKZG9S6](C\K>NAXfJQ@1O&TLd9AY<[Ma6#S@GW1Q.QQ463#=&<^SK8C
>6S1M6[UZ9V>c_gY:RLX-Z]Rd\->T/IPX+HF)<TATJe;Q\F^B6eM#J3?>+-3a/?_
TLbLb)f&NGLb,2V3BSJ_&/@JK(KVUFA#\NK2QfVP8B2bdd>#dZG>A-EWcFeF^PC0
6Td/H(2,BYgJ]DDdbB5;Jf=-dWXN2TC>CF&0eg5?aGAeYBMg.KH#8FK5=ZS@R-R_
0f-F?T:WL3bB?-^gc47S0E&VQ#PFRYdHM8XHU(>;bf9I??Vb7F]2/^:ITA@:1_a[
]KX?Eg9^K6[:1#3;[K+;Qb\0.,ecg[Hc8G2(P4<M#;+NIA3OgRb(;;_81X)L(e#Y
W0^@\AX<X;(#9(,fE<dUN#,H43@ZQ9J6Qga(Zbe1K25a(R>FT3ac7Y9d4:+b>0Z?
S@Ue@?aS_Tb4[IJ@B5cMUP\PAMIH3,X@0cg)N=MaI19SVV&ea/B#4WFOB2].)OYI
,4LEUFBb_6+AEK\Y[W3gIB(g3\AUQD[O:1P3H[_HX>PB#c=2.fL<\gg,5KLE))7W
(dG42;9)D2)BPM0N2)gO[XYFA&7-<:_D>LR4]1gcbS4W]Y]V66e;a<^^LAMe@f>f
H[Q5N-?=7M1.-BV,5,c)5&G5<-+\/Y?gMM2J=JDdB(>1)NX>.;\\SWXc1aUK/.N8
]:QEO_0&L+I3A/ZH<FARDI>fX->6@C)>0,#QaX9Y@(01T@EQV7&Z77gO0<ge5<8X
?fVf<U9<TXXU,HeHRN8gDQHA@:34dgXg-&ScR_TE:^Gf9MgWICN>&&;2B>TL4WZ^
/bDKZ@S1QPKQ16T6T:bA&NF_USd:Y#;_15@7B4#P>gaD^T>B4.DBV=[:0G<e5@&c
W)d5Wb6:[XYH8CKEOAP@eLUB2K@5NW[5;bMX&1BDG.T=>].VTaU^D/0WV(U01<9A
^#>IUc-_;)(:<M(I87<3F1Z2>LY8J#(&^#f(#^?1a3,HF;f4g&[8TJ[B8ODE03Wa
.Ea.[#M4#\(M+dBI6QeL7I9^PT;Kg(SRY-D8O8-&;UcHBg0/S:QW&P.-N5-XMDRT
-HRGZHE@5FOL]U]<0F>Ag-5Na^d66cXDReSfO5C[6P[_c:,53-RQR<-^]TRT;A<a
O#BVPH^61,5/Gc?b.P4F1(6/WZ8Y8SUAX(ZabY8^9SBK=>9>\=:V]V4=Q<g@S=+#
H(@E=4=><eZ[Wg.35Z,TB^BM8MBfMRS,P91W.^g_E,W=EHGBBd.C[ZTS3LTS(WY0
g4UQa@O9Z?XXA;LXP+WaU@8f.TFX[]/#:6a8)WaV.PdAA?UK7E_gQdP^\3N_+E,L
9<OcU0-4dF8E_U80<eH:Q)@=Kf@C;SC4U?(PAUa7K#gX@OP,TN=YXLD[f9Y-QP\V
M)>MQ67K[K._+fW43Ka.IEHA3f@J89.42_\\JgLG;&W=34R9&g)0\5_B3Lc86#DX
d-0b\MWL4A@N#Q[Zc_2[]9K8=Gf>DLbcbL8GMJ4L;Y]S-dc9+YS;WN12a:/bg7KY
9@+Qd?E/g)Y0VMOX[3_b&.]&[/<@/&J-OE(-[cR@]=_#cf7+P&O-B+Y?AGT(C(,:
P.)C?/LCT@XP6&cH=U0S<7/@:P9#SO(0Y?Y[IRG+1F\PP=IXef\;Z1-.HD]/15KK
c-^I>M^;-)f01=CG;Uc5DAadLVNS&cGMGH+eCV@TTPONbBg83OQB,<F00E<0O?O(
OcXK-L7P?C>D2/&R7/#0#,gH[?ZUNWZ[;:P>c0&YIKMIEL2,=^SXaI?RHB@\;2d:
&<UcC.#4ePf8\,caT/\D7bSRL#S\=92QQL>g2\6[=dc&A40[^SZNMU3g.7Od=58<
6IRI@@_>&NLU3fg#-,#_WAcMY(0,ANeac>NDe&G7feJZ8^SCgQEd>6(RS:,Q<:D_
#K)&?Cc);9(X?/c&d@bVMK-G8WGe&^GPEeGEZfE(/][cEO)I\CR_--QS-=Y?P\CG
aY+6/QeT#^],gBKeY45P(S&\b3>3#)KR#^I#KF9)<6PAaBXgQD&dM8VeUZY&]?C:
GUE:L5GWHA@)-&5W^:2PPM4Q0K0+VXW#^6g^ZRZUK53>6>/)M(29fcCb>ccb?M@M
ZdNT<[+Q2)O&>0+]^EFaQUc<@;,Y7Ka(,_ab^N.\;Qd/WVFTYGJU5]YT@P\]@<b)
T\H3?^MJ7,^X_\O2KRX1Se:;>fX2ICbMQdd+>IN-L=+?IM&Ya[<;fC,DB4+M8Q=X
5LKV@N.HV0W8D0bcC<F&RNE860f-P&0Bb7J\Ca.;CcS10J>_cAU3AQBKT,Y#,ZFg
O3^[Q++I,)M97+R9);6c;\e?49PXP#LE^1A]^A#=0K)/C>RQI9)[:+,X]OH/<9D)
;Z(83/aS;[bPCT\ECX.MdRVARMIW-<4ZOK-L,#QG(^[K5S.aHX55)K.1QF<?4[Md
O-#S\BBD66H&+>-eZJ0Q]+DR9I@,B@8BKBY-W6VNLDIY&X44[fL_JF<9CaRdD=cM
NG)dV:C>2:G,Yc(#\\5gLOZ>T,AdbJeEcI9,)VA79^XgaL]_1Q(16b@GXS[5T<S@
B;Ne=KH8=g[?XQ=_?_BeYH3B^?MX[Ze9FRH@[0)Pc++=&G3RDCGA=B4WWH;W(51(
O7N9c5/A?V\YN@7O6\#.I<NC:RV@[HI08+-C+F24R,_0&=A(QFK&.M]B4f6U^S0(
O,?I+&PY;ce115KaO8QT++bY/,0b6Z32?NUFaP<b_Z7Z:0d;-^g?YP@J1Y3Z)@E,
SfBB1>3)#XQK5QJf2,#\N/gXPEF=1Y&c-JW-B(U36/Y>^;K8T3^ca#HGUZ7c-c:U
(33CaX#/U>6ZBBA@dX3?(E)K1NeHN>PAJc/XP;^&L3J=J-=F:7UY98TF]2c#&0fU
f2KJ8,RZFB1M7FBRf53#10A90X&gWQT&eRIS5/9e^R##0D;.W@-egZf=9:+PYDX>
TBRbC@()XW+;)&WQUU-\3G/()19H/T,.)+Ff/8aME?HG/;8IN5N18cA2@dBcJ==H
O[O]^T/;)G?fgbd8Pd5:<F-\2JGaF[AM#0^[G,<aLa#bIag[)F8E=gIV_gU&4=,^
/b&&+K(C;1cdF.:SH+3I7gd\b05,324&@/X[O(UP4b#.;;LHG8NgfUe/+]daRJ9O
1HPZ1QIcO3g]O@ZO?LD99_+SR&Z3BS#42fYKXb=I_E#YG]M/<B#f](@W/I5,aF[f
eXR,+dAW?I/+:fP_F]3G93J;DP)&JLO=DOF\.<(PVB]f2P#Egb#g+Z7BT=(Qa83+
J4.3-H0N/8YF,V2L-cF9fJ[>O_F=GJ;DW,R+8J?_&ESUQ?[2T5)_1/^BE_0?1K@Q
KEfKHFQI?2,1L0Z^cgNOQM<@VIVa<OIAB15Wd@==#0T0>bZFBF+(?260+&KA6J;K
=<CSDD.,aOEE)R83T;c@&F_J&OGdEMaUD>K(e8_L1Y#.JP6-\>[/QQ4VJc-\Y:I-
,Na],D73>c:\<8FX]ZAOL?MWKN:@&_?7:5BD9d4gK&/)g1^YQaI/S:,d>W#Of\g,
PKcf/GgW[WdOU4DNTfJfJ.1LZZX^S(^9;HD2Y9/#).KO_e^,d4K5PHYWN8FG,8eb
;b=2O-/#MY,E9,U?H/KZ<M8V/&Y;0;6X;c+75d4UU\-3Nf<>bF0fFHK9\>[&^g^+
>5H5^Z,,&7D5<a;fQ^DWDOF?[F@^aC1/+Z0]G-^^F;G&@C0&H9-0@Q>A3HF2[Sfd
M@/+<NBY0@<\\F0CO/9;U:J9EHK.<If;3dV&K(VR66YKee>bOcALe(5+AV2/?>D[
Obb^A9EIQ8?\S6?6SA06Oc,3gfeX:QQ2gEU]G@Q<R846Y4H@KTMa8A@Rb_f2^O_[
V&E/JTB+[L[+g46L;d18\O4V34L+g,4GI0A(1T9PbY??=3A]6MX#:B@QeOUMYS#R
\U0MNUWUYSd2&)TQ=PE+c-_:4A=+Z698;<Z)QbR@fcU9Cc_)@1)XN\@RMRW#6=3W
cK(D;KHMC=FRW)PF=>9?E1f\98W=/d23G:dQe>6_:f7DaOfO8\97bS^egUH/DZb6
A8W164Xf]8J(_e2+FL+\>MG-9W]69UZ>>HbS(7[B<0=dPN>4?SI4:6L2._]:82c)
BF,]3c<S?<#.;/b>2V]Y5E#__ON)8PF_VSAc\&&++P>,73AEV@WW(@/DTQ/,S]J4
29Hd(;=6g1M#Z_fJ5^6W44B9F2bZc?(J8Ha-+ZBAc#-YbS^7ZC@2_aZXf([-3\\E
eC()7[IdGL7W0<T<&d81B+_3\>CR7.P^QUY9^\H?1,c(bJR^38-4f6BKI:#GM7:0
9ONg2aJP=.Z_1?GTJ-N6CKR03_(L.^X_ZINUf/2)CdL8^G4g2T\,,N,UM-F.@Z^4
=We;F,2C#[BPY5[f-B/I1,5DDB^QF66I7I;VNdW2(c4a4[Y[-UD#_gcO8<N&&?O-
CQ36N]A,=#3e2/:FS8J6KXK^=bg;Y&O3b;[[>@gE^f8/PAP>B2:6880^C=T+>TM?
aZFS]-Z>:Z(EI=0><6EWP3]/9->?5b9Tg9=e+UD5f[+:f+4)4H(7J]\4]MMQ,PJV
LGROL?SJ6>^2eTE9,1ZbDOV-aO/15e)#W;R)SE;a++68S)bT\W/Q8\T0Y41gYYY>
-6@R[S\_TP?>(B>UXIFfH1GXf,1WNU?2DJE5INF64dD76><Y=D(0OU==#-R//eBb
@G2JCgD^)F19f,\>-bUJ_&aCB4W,M6+2GX1N5M7[EE,,aMQgUDIgIZa9\<[ZGRI,
fQBG0NK,S631,Md=c/>7A7C76K\2<BK7YFb_4.^Eg,1_-(O3ZGeeIeLWS7P3I4C-
X<fQ^>47G7-;@#BHY3Dg]US:N>dg\/a-[e,EdQ2Nd?PA.5ZMI@9a=8((]C,N?,e0
G,,D&D?E4),;eYC^[>\R2]d3.;/NH21&/T;KA52>e4J2&]L50N(:]f4A2\P?Fe,W
/9FZ11C30CSVbT,CV=9B=LGXWG]b/63YSB6W76NUb:&14CQeVFR@_Y5Ye#OY,OI+
?H-8<f6W92#3c/OY(c@];5fc;X\P;3,T]WM0V5Bg9;2T##?-49]/\VUU4YRDcWCL
2?N/L]I<046Lc&49VMXM)G=fJ&)IS&Y^bWb9e;Ig\F>@3]:\KcH75@BB/9?_;XX\
6H.CXa&5dTCaUaC;[^Mc11-e?>N?(e?HbIIQ(0)1LcOW(UScf8=EB1)?0ddTCU2O
/Y/c.WXceUe4;UZ7aUP8W>DOZ&^-V-:;S)37H<>c&Jg4Ob(f01#@1f4WaNFfg\_C
H4OZ/)5:b(H,2FL-)6aOZ01M5eM65JJ3@9\]2c.bgWFJW)cccagf+09W5YHYd)Y1
K#E]IbD;5dG#51d>&3WP]FD#c>85&KG8>&2b6-.ZC)7b,5P^fV)EBD,P+4VQ0+0\
R65Hcf.?]+ac.9:GGGV:_,JIG(7T1TcJ8M)Y1,:cbGOC3fK0EA?9OIBV[=QDH-)C
#N>QA&.dT_.CA.LM&ICfFJX0JA:PTI.EG+\f^OOYNHCJ0^JR44,IX@:TeFfgaT;&
0B\CYJUD1WR[9[,DNLA0/WM:LMHN/gD#ND5fgcPKONRdK/-g1a0S1:e5);G>OC09
C&)Of<<]I=3);+1a2aD=:HULC7g\ZWG>=#bbceSP[J@0@BX7<A_cb-0PP/Rb=T9W
I]RQ=A(=25Q]\>+];[VG6V8N5aCaR^I35AU]df#AX3FO?bF,@MFDY\79L/Y<0TBg
gS00;abMMd-dK#+I);Ne0Z_7A3YZTR>55,(AM&5G=7CJ[H_V+Qf,4Ac&]<JD7J]I
H@MG9D&(UG;f,cFC]d8d]a@TVcc0\3.BRO^P62FLZS1M8[._M+8O7eY6\B.d2#;5
S/d>77/T4#3(US9G7DA]W#]5_/DX>>YXM?e:(abURY,Q4Z,McK8S9CY);Z2HNgc\
<b,B)\2gRZI/(^54)?K&J+KTG.d>>C2AL0+:O[:SJ15KIbaPH21&LQK2bATL7#eZ
;c:6QgbDe5?a8gW(aCNbe=\AV<YLP,Z/H-a=[/DW7-3R>Q-B4CaQV3d4^N],C&CY
A=7PD8[a+SA<L>dIIM)4Z<g@f>RM=#ebWH3gU(NI8_K(_R(,^fGY^?JT[-,P5g2O
OH;7C>\e2Q/dUDS_5b\4_(WLW5NMU]U6#WS5WY.S[]<cb7CO)OR)OF/_CI1>KM&9
aY9aAKCIRGFNe#:K=9.K23WL,4C,fN;1_MWJR5_QO<TI\U_:E;;;7TPX4UVPRMaX
],<X39f(Zb56G8A.UE^49?8Dg/9.C0MP/6<aA/26f;T#AgLfc5H]D(E]3DCgJVd4
A.M1?18L[;BTbBB6V7<HUg3_U6C9^P(67,gDNc&V>L+F?M2e]4HI)]LK:OX?)O^5
;V3U<ZAJ@O\]ZPQ9XZf8XX-:(31D5=YQD_(MK?5KcHN2?D[VZ=fG5^>>[[SP@6ND
]U77.aDF+.gae_O4)\27N9ETL^/\0]Ng)EB9-bD4=(?>gd/X(4C:A]e\H8>6aX(\
H,J1]@2?.:D,MH6S]@VAdUR(7&=/eTIBg98[8,2U^GH]6#,>5+(LF:L[QJD+N6X<
].79Hg5>MYgOX<;\/.2K87E)&a+8?99J?gR#=-_.)D3/S;I&(c?C/2?g6G>)CKGI
7:(M+RQZPDBJ9Y_UPgO6\b8a(_PJ009X_0MV2NC];ALNf#g8YEd&38K3BE@<WML^
;L<]B8I_Ub@0@XJf_.M[EA8AQWR,b>@R68457KC=NbC.1=?X2b]/U16_U[0X2F=,
CDef8Y=@-R?D)?RG/(=;dKWd7.N#=.QF))-L6E3?9&:;,b,a9dHgF&4Z=82dg:-c
]]E;?C(51Z^2#5Q;5AGH6RX59dg@P8N^O1TCO;;0#F6+?HO,BR:U+eTa@eXYe4N@
F/B_7QD:QP>eeJ@=bRP@0R?\3:X(OAe?e#S@-DL<abJ>.ER#+ZGU)8YYSJ-XdM72
/R<fK;a5J\V&,^R.aC/-]X\Wg4F&Wb20_0P;7+VTZM,4M2@RV3N/5D+66[d[(B)=
-R+P3D4/bFFfSZ2\-CUTW[.)dgCN36?I89HGPNd?Y0(?I)0-D7=VD.+3(UB>O0<Y
PVcPcfXU2@2A1/S&5=.Aa]Eg[NI(GP#[?9F\0_ARTS8b5]F8+,92-JP5><URNYL6
MKg;SVC1>O#YNOfU3HFM@W2Wg,M2Fc+Md(OFJ0ADN)1)e(K/@,6;W?DZ.,a@:^,O
5?A\(BT;JVI,=Q/C/BaGJdJ7OF;@W2JX::dM7He_R^_(C=f=E=BS-OQ91HcK]]1C
>LSE&W.[R70.]FI23;\B?:+B82M[GgU@RCQ\<G__gJ:&[f\+[Za)/eg<LF;Q)&Ab
4U[,M-+PaE&<+>2eZQM);GLgJ]@gW?PZgK.FX=5CX]UK1[OBSGa(LCS\42e_dcac
GPE/@&U>LXI>/26aUJJIa+UMOW@c^1)WHebR_5^d/QeaGL2S86bDWCS.W;0de&bI
@\&F2L7-\&-1C6F.Q;TV&<DS[Y(F&SLaK0J+F>Sc3a,@ZHQ::3:=#/AU9\V/fADF
XO-\.fB],d&5;<<MU8+T=YH1eF5/#XX[\2c6;F9_cI0^LC?8=TV)D.PJXG\CXVTg
;XIQ/,J9gA/;4V)FD)V8T>C#S#a(KD;.+/R,\,Y2f@7,g/Zd=(QaN\M(A=X[-aRI
MG:R,ICQLYZ_Z_Pa:3^S<3V530?T^T#44E.b#a=gH4CY#[IN>#&V2OeFDVHX/C3Y
?O\0E\1LAVfB.b4U0DA1U&(_,d0J[<Y_=d7+fY4KS[LATY>ZSBP[;dESB1e/PbC.
3&Q?3d2VQY,0D?S6OAKF?UM=KHA\4OV6HAd;gcOdMS@^PB(aPZT@]+&2HX7JU9<W
@<;+b&7:QD?[G@9,.eDOZ0DB7WFEYRFa/J0fTA&GOg8QW;1]J-F.-WO[MeOMg#KR
^VI]1)Y@ZOe=AGcIM.J(S+GeHH7X.UX&Z6)Va)E8KT.3@7=)V[+G6@]P<YA0SS.\
]WGUIGII8dGf]e.R4^[G^^;KG37A+\5\]Hd=:dV]F^97bLMVb_+1W2B>H86C]eKP
&#L8\J]WVG;I4TRE:&fE)6C>P_JFfZ#cT2Z-9AWdQE-?^=3ACMB?Gf]Y^Ybea[8-
784T1.e-(a&U\DTNf2Ub=d@Bb7^f^+0.cGX<OT5TE2E8Td^7E34)?(-fe<9fICeQ
ZEf4gf,ET,S,L#/P/V2MTROW/.UL:=?4H05:Vb?/3f/7[FOHdSeRY-bb)U7--3c.
a6YW1)=JG4HcO_(-@&S<\DMTe>Bf@L>W4)M;LMGdBU(UMX<)M74=\ZR<2>YK/F-T
I^c\9^]U.QJgY35TWY-2D(00&?f6259X=P8,<Ac1J<5TN:g@[ce_>48cF8d_AH0V
b0N/D@NE;cW3dE2]IKWR2\.L=N-bC+dfFXEB+b<Q/7,#=aTa)7a8aBO]6KXP?J]]
Qg4QTM>E11?-T@#?.+?&2CgD5@?7H2],>HS,_SZ67T46HQBL6#8Qg@H-I9ZCbb4>
B^S#GAa_9WX4P-O=\fd]10\^5D-H/D&?cWI^5MCN4,#?J-7e4b_D6I2-CWAY8;^,
V]N)8P3^MW-bV^;7LA9SQCK.d/9&7)3_@F(;.ON@G8YQ5>#,/f6[<.#G=&A/<aJ9
Gd8P(LS4^SOdU?.5UOAF22XQMM8N89MDX-Fg4BH)9Lb]P>4BV)#AB5DCb&U;U[gI
O[C/+2_NaA2-E)&.X0c>UN5HcU<cUKIT&]M)HQ81_6<bRB2O\2KT00YOD[/_6BSG
9;dc(6M1=:HCg.D8d]4X1d/+e33fGV\dKSD.D9UMb.dGN6ee]^B8HLe58egUZO;/
,@T.FNC[MfcCH@LBH/0bIHT?(=[>;ZbBdc/F36;;&ITI9OL3HCU8[J5aHJ^O@F3D
>1Z,8Y7fa=f+9<HC9B-fF,XLPB#_(>\Q.QY/16XJUZKcIQ7Yd8dE1<_#EL^)-A<P
J.EH[)YbO-BIE-286HNAS,RbGQ2PFXZU\=\Pc=2?U,Ife<d//OA,JS3-UOH?d30.
RE5>\7<S/V7:H5NZ9_Na&D\-Z\+#U1G4E4B=I4H+.:?fZ9]VZ2+>2;eb1gdIfc.c
YTSEOEVS.)9H1f=eBEXY2U\WL4SHc-=1FN:P>/T0X5T:[(/WZ.-DFCIF#aSBb-Y_
abQ0YB8K^MY)L)T:]a/T-X][)SU<_1aN<.L\=&YS)+RQ8d@AEd;(G@)LY?B#2^RL
SB#AMQN4B[=:XD^OYP?>-eBGN#+]TbZcI;?MDZ6YMe2GXNBgK]4?,(g^g/fEfFX+
JXXYAHP@4J1YTC5[.HISK<?cI]@8/5NHa/aI2\PW&O:(fY48L6UBA@45D_RJQcb^
#3fI)+1FH)15H47GFdg.<d[?]&K.\I-F)?5)fG\0&]YV5R+0J<64YLN;^&7HZT;3
#OIUQU\e^bKMFBW,YP@8O,5b111XR9/e0A]\YN342]NUI)8>82)HNN?\[S#ASMPc
b>=_<WX.?e[&PK+:gHTF\,#VICU>d2>GP=f5:ACV@gc)X]^ITegMTD028C:@QM]U
eVX#0Fc5OXHED@=U\\2T;)A/&@+6Y_?Tbb:JRcOdI>V46f:NO6H#^/C=Ib^2R-,&
CC:<0UNdOKLV?WMQ>66L@7S6RU>b_:_3X.,ZbRR&5OS5BeTBc,=[eTEB#<3\6<:2
9[QPN\9H9K(<81])Q2#KEX5DQ&IcT[?@C^CM(U0&]?8aQ@NPY&IE+AM5Q_#^--,2
MYF#1U5LdTIaP+Ha#5I2?)+cB)YI1^FVKWH@4]G2,K7b--?ae.#^;[)#.^VK8]C?
3ga6)dS[a[?;M]2RS-I2e&K[JDCGFF@2?7g.K/0B>K3O[6EPCAN[Q[Ge&79RXaZ4
5Q4/3H7IV\T5(L=,YKf3MWV<T5.;K-b2:]FX#5CA4KEG>#^>4>(TRJ6F/:<B0;U7
BQ37,,69>Y>K;EPBeL\G,UfK#\&.ecWf4:GOD\H6X#3/7WU(S->JXNAaVM;LVFR@
\<eI9=U-)ADUEa4X1HS-Ne1@LIQaFL<^T2U.P,\O0P\1ZYEZ;TS9TB7;feE+IA/8
:Wf]eSEV&OKUcD2fHU=+[?G(f5>1.cYD)b5M7I5_-B.D([:[Af/FYbHX6D6O]IdU
^]G24H.>^A;dY2GgC+L=A<[,VZ8(>9^FG?N6c\QeCC9=7Q[UeOa)dC[U8Q.SK5I3
[JGgbC+YX-Q5OWc@)4Y@7@S65&3eg2aT/W4+b:0W71=K0;0EQ5+1T_.;Gf&C3BH;
C)=3]8aJ74@\GLES0\9MZNGS\Vb<<cc9XC865Od)1MZ4(?A<-OBD]9-FW<PL,E+c
;XEQG&D&YQeTJ;HP=bNcK:a4RE2eSY-.60K(;;++S/Q:^4>]_Q3]NC^(F,R]E0<,
E@Lf>03/9X;FC>]Tc?-3N-P,B8Sf56WIO(SS[+(PeF5FF65QC+c^dD-CW?Tc-g4D
9c_,(-J:e&aZ9>?@F<2:(BK.IBMTALX<V\^VVM/1C8AVIEA,Y3AJ45L2Q5f87>#b
-0E1FQ7QPF;aPA7@U]1M>#XEG/_78:9Y/[dd8QP8^#;XLVFUa\,Y[K+2>P.f3gdc
2QU21cYVQH7S#N-:6/>WS::d,TdC+G_LeU2&V2[]-J\,PbdL:_0,::aX-?+Ed.#d
85&eQX=XYc?05;@21C50VA,+^cPW@,.Na.5a-GUA]@:?b/5[P)?UKP\IFR#ad4W(
fKR2E37X20>PZ)5E^c6BM?I7I,#K&D4\9eTORV9WAM?@=-U_Ub8Y6[U\=g<?4?(@
Z5O1fJ^GKJUNJH,+JdZTKf4.M;cId\.>X>/:SW.Cde/&7+/TX5UO&Y4E&4gL1b):
6:I-NXJ70&KD:+N@52.K;B]:RB:EE9Y3X#+OZ8WCMg#X9=F:\Qdc0B<W6d62IKd\
6fa]K;)7+;SHWL=)?_:<d8S(@4^=9_:I8c]H57GH&Yd)=YXDT;]@b9&0D.aeA+e+
X[NDGgMTDg\2F?DJJ_g@RWJK<N/@@>6Ta(]O/7@?;B;fL\2gE</2S]YM\6V]W5-+
D2O.bV;d1XA2f+T^Q0F62;gdIfIaW9A5AVNEOB+Q-C#-]5_5gR;(1c[4&;OY\?2a
4Q[)=+@D_QL[&;:=6<b)_WC1@R:[^O(3SSe0+6d)/#E2+Z&_R3?<,.PGAKO]-P\+
AC2]-[S7[W2^cZ-eb4=UdRE4?KYG>gg<SPTgC1^fb#A/F(M2QX=acU,?H4UDKCW:
#)N:Q<.[/Z3a39O/6G_G:FGBN77/2,0aZ9)Pc1A.O77,[4aE747=+&=eK:]P)H@F
=Z]/QI4NUc-F]JVN[Wa4cZ>[,fR=F(Z<5\d0SGG(_[EIGV?KSO/aXJG&^YP;0E(X
Sa0-ZI6eGWd;.AGEQbI3cg>LU?226TC7I,XO)[<\0ACOCM?CJBIdMYFEb/A@2A.U
U]J;0#-<N9.?&(ACeBUQD=<O&B@NGZ#05-eH37BS,O..4\&F4Z;8BCM<D9Yd?@9N
,ANQg.+;eb&W6Y^c2(D3fDfHd:.EN?AHC4VP>\=/K>X>@LY(WQSHYPQg&6>0#Q.W
P::eJDA9(_J]ZIN]YAO:.beCZ>fLb+FL0O0[;<3D^56:EP>aN.F457-9<Y#4:3+F
Q=f<&Id#L=6M7</W_5LJRcR]S90cO^WU6/Z#+07HC2#@D]G27[2@-QHC]A40PZ.0
^,^1S0c;TYZ0ZXJCLJ6E2Ha;;Y0RSgWDP:O0>4>K1J6XY7O\a6a5J)&>Xf:c4fH>
D,M9IW3L/G2U)T\<9>If^Xc\.g0).<1Kca-E<d(-SMS;b27TF@UM<]D#8=?I67)O
P[c.VHJa@Cf?X,)SQECPXCUd8.S=:,C&S8AEAbF6G@2D,L0)04H,708E6HH_L9gR
F6c3^_T;4G8]K:#,?=:QIOVE)=VYAB0D(Q):d.H0ZP5X6-Q.Hc0M&>)gg7[<g;#b
PaEWAdH:OEd^Pff)_Cg(TV&c]O3A6;b7#2/g[T;dXDUO@g[_c_8E,A1U),/W5ONB
-TaJ-Z1B+6NHSM)L[YL)MX;2J+^5.,+Rd=G//?<JS]f=R:_>Wf\FSO(g_+&Rd4EV
+7e\aW]9MS1.;/?(^WM/+WD\J8S-W@+Z;E6J-C<AN[N(//C_?+GU42Df]U[2eTHD
I.#4&@/N07-)X2L37M+KMB1:NYBRdb21e;7UgG9JM^O&e3Zg=51#Kb\;J5BGWH4E
8E?X\3:??;a(=PHXR[0\/P?1fRLZ<O>WL<@V9]Y>(8)SE_D22;>,8dQ.Yg.<97\1
40.JU;VaKa=bgeOgBSM8PK,7GRLd[6VO=V\QH7_?0;SK2bBWO)e\>+\EL>LG.bAO
Y>K-3H-&2;Le8@[@W^3/LP_E>7;Z<d@1QMN\<_PE0ZC24(c#A+ZeCLP.Y#g6-JKN
;4UL9=Yb1TcQ22dc:3cL\EUW=:RQQd[)]EA[&Gc1fg/RR_3-&9PFgX]74:=X>+eJ
eBZ\Q7VF9FQ<G<RY<ZNc05H(W5dN\]g[@8;Yc(T^5W66a4McKd^@E399Y4bCQ(UP
bQOPHY5A.eA/\.L-b3BP^bWT1[Y<NW2NBBR7XfAY(+Z[VJVP2N==]R#cG3I1PV4X
(+_7<O=3Y4Q4BfFAU;,XRG7V8Hbgd=YQcIHH8?a<-?,YcCMNdbA&fLYAM=4_9E9^
Fb8d6R]YHGf5Zd^(J_YVL4+)C)[]S8]L?DP\/e?J2ZUXMaddRG@3OO1f(I1^R^Ba
b81H?Y&gH2#]^.cV\LGeGJV9DG-a\;#2H]82M1Q?[0TC=&:;e5GZ)L9DXDPeKAIJ
2KJH7&CQG,7U75]eU>D0aI>daMN/KOXOcG8?)6&0[eWRYd2eIT,NJD&PIEK&UF:[
Af<GQcO&N4DCT6_+M8\,W.;8BAIHbYB)#JTcMf?S0]8EaO]13>907=ZCB/)b^,FO
OGff[@f48L[Z,;Q)2;P9R+c[c__=OW:4A_\XeEIUcD5[>cDcVF8[=F4872:]c6aS
GG.1.:VdJ8LK3MMN&,>TSWM)L&e^<Zg;R<1#5bEGZfEMAM\)B0O=QLE.(EIUVPD]
N(]@&J;6\?L#WXZK;T1VJGP/H7aT[ZE[fH_OQ+_I[/1ec&4G3=8/eW\Ve]a[g([#
aZ7-IP7g;^c>8_/HC/0HGP^fNJ(C(a<GTFEG[@J+C.N5XK1S?S&YOZP@^,3.4(P5
gY5A&Vd??d[74Ra37]@AF_R&@DORUOO]7XE/,8TS,FC\=e4RL&/&2MFEWV5[deW^
H#d>;DRV0Q7@J1UVe_M/.d50&2\=.C[E.M@_+J)d1_#4&.V^^Q_U?.?:AJ&QCG&W
/0Y/(\CS--3a?b:(2S,^aA2IOOSVJ8BbG3d^;B?L24UODWaX[B/KUSB9;0K?1T9U
3+]H=7@WWecM>_=P.VF0e8(\Q-KZH&WRRFGB\f\S@DLPX?CRR<CWTD<L#:D+-317
4FFTRe0[(WbL8YS[F)g4g;[=P6^VgWgJfgFENeOG&QLae2E;+U0N2Q1=M&g?#\:Y
HgYfObXHJ]18K@+B\/bXKH&#4@e<<6FAO\;.gFCXO_B7N4NCA@ZC79?)Y3e_0X=)
MTgaAB]?2a<[83dYc23ZeF)9L^<:_953;^Y)0M+](@9b+4eWCLbg64D/a##CAB>8
M.-A61A8KJ?>XfL#Y_?CQ+9[Y=JL#4)L8RE#LE2K==3X&cbd_TQX6L8=@D-UVUEO
X)SZDc:7/_\O\T,CHPLEI+Q1I4\ML^LQ.=OW:L<.@WZVH-cS.QGQ.N#bYOOFd^T3
?aDT(6J=9P:W-8Z2OQJ2><HHaC@WN63U,JJ0+LR[B=EV>IS5Fd3c7/B(G:3GZ?I0
Pb7>Y;H](KcO>&>8P3]Q=I,^Q]88MfeI8<]R@Qa7b\9EA3[fJgA,UG&F&&:>Q&A5
/cB-&8M.D=^/H977:=#6M,Y<5/V-(&^gCIQESg1^4_-_LG1S9Z(DE@RET\_1-+SF
dg4V?LGRVNfTFO0T)UK>#-MI=BGWfNPW_K.0(NI4f:C#AA5J0cGN9D0^D.@_SC)N
__^H)a7W8>BF3=OC?L]E>_9E\TF45d+F?[3C=6#\gK])H]NGB7(Z#aACQZ89-Ada
CFIS]3MGa8&L-Y@84>8;HeJgU;-&W,6e7_NQ=Z3?8(D=g>GO(JNVLK=N=7L^<_gc
PaPDFY#>d\(NG7E]KCD19M9]]C>L#e&R_b40YCS)0bA#RL\<c-;)FST]gBK/1BRH
9^L]TIGXPD([g1AVa6d_S.I4TL?dOf-G0^6SPc#O[TFR>@;LH[4P3N]ee^EJd9-]
]_O0E^CB4ZNUgbQ6L\C42ZX:bZTB87bY0^5d;+@5JNGgHKPf96A:6[Y2YS/gKJ);
-<0>7V(^[GZ+([(LfCM4V2OTK;<2<5de.V/@DS++ECAc]HD(>\2U[30@.,e>eF.c
H:U=K,E,B7e-(NB(D;F&)DVW<K],@ZOYJ:N+A1c:PM93<=EN:LV-7)SN\<WF(FPf
1W3?+cVg+7J,3a-5E0=fT0S-/Z^Qc[:a:D[<c_(6;aT.fbC9Oc,8(TT-?>I26+D&
WL0#@S]0bS:D)CVfXZ=a4Z0JX.Rb[DbH,APUE?Aa+P=-4:a_WMEACd/BJ92=4Rg\
dJe)KPVU^dVN?X3.N\(._[VagJ,@9<bN6Cb62J1I=eT1d]KS9#XNMd9I^U@[bG2K
7Y3C.@E6H:AC/S;WJA7cK^T(N89GX]-.,T-8Kg(L&@0^U#bDXMMVUE^6CQZ+9dI,
0X:ee]+DDN]=Qg<?NL:5FdB#Gd4&[.H6^BE;eIX?gVUT@T<)74Sb_GS1&-_(]]_6
]7H>J1KYbL]SDOTI.(K-,JaCMfD^Pf4>g7E@[)F._UCRXKM\R##5Bc&>RZb9Q6A@
K.=5B1HV_9a9C,MWYK7:0TM6JF.OIR#O4JXLb-CRL&T.HDU:,&\Ce2:<\=63RC+:
8UbSUCea6YKg)VVLZ=C0#CWPV.?]HXHf6JQY59NN;\b9#MT>cCOKG5:@QSg&8<R\
VG=?Mc5g3J3^50UVK13LF8N)^<?H[1JDZZ6)>?34,FHBI;?9WRF^@.YTB+:_JE92
&:GWS(.:GbP,NL\3KGFG6FYPK5XGdSJ.gR=ZOEXS&]aEWV[TV7(D:>#NA@5Ig.RA
3Ad_EUf=SZ62+TR9P7>eB/0N5K[eT1#dX&/>;3VeI>0M_UL2VFfc<IM.ZY^2F-L&
R9eLeRRAgGd=A;-MT9^1Z283M,=O,2cUIP9-[&C3?OV@aeYI8WS;\U-(4=H]]QBA
#E/bONTU>2F5G1MaR04e5)VC\8#R(AY@BY7E]f=/9\^H_O62^f6OGTeYBKPMF.:B
LXg<X_;G:LYXP-BHWXU9)K_=P61YWgb&9)\,SV&#CD>[4+6N[CPO1)d:,=ER/,ZR
X/M,9#@VZ#X;V./Z5DTe+(+^)-c2G.f/0BL<UbCJb<G.L3F5a&S4?P;^>9JC3B1/
6\e2EDBK0#VW1Vb2IAW5?+>)Z[Y29eFeW^3#^DR6Y(L&Ef>Ub^^_H]6Hd,=T;D]d
U,4>9>f#\?O7IO8a:J5#L&N7dH;YN-9+ITc,&FAbWE)4bGUJ1_VN>c/]&0c56G3F
&1^W6[edV1=8#BVR3DE&UgIU.d#4&ddPIMAf?&([d>[b_GEEIA#CHUTA;FL?f_:^
_FOES>GEDNJ9W[DDAL.>bM9MAC&.-_TH5UIdU_@5/<>XZ<Y-M,cK2c.f>,UPL8Ub
>QVAWcV:6NQ/&^=fG:&b]H;c3CI\5d)?F.fIcBO.+@e3P8@DZ<:cB6.RY7U<4KP8
a1RANKfQ34?^(#3/E:9/9:.4^0.WHaNSB?[P[>E#4@SVP,D/a)d?+cP\B\6;5G-,
3Oa&+)TR<a\NA0,2aT:#56>)f6S?),;/CbeBfO0Md1Y/GJM&F&\7D&O0-[PMS&])
f#PANP<<1c3ANH0cP.Q286M.F1Ad0B(,cJZWM1bRWg=e\)bb@(B.;:bfb+;T7FcH
I(AM_HCbUH-UVFLd9BF9H+/YJ[)MOeZ]+OB0Dg.G:bSI/QgW=bSDJ.^BbCLL)ELY
1S,(&c,^6[8eFOg6U)OL2M-=KCJEA3Z-C4[BOSD^L6(;JZ5>(L-Z7LA:+UM7#cWO
SN.@4\_SZC5RJVU.\)&7ZbbO\><_;gOJ;4-F;\CVeIfL9X.3)J#RR(19WQ^7bP)D
--G2\5Pe=JT^J(6#3C(N]CV>91GGH,R>Q3e\P]AW48=[4<eB@>d<.7U\BO?<1W#J
(@@Y,VWCFBR21c<+YT\V?RPJR^,TO,#BQ7Yd-;8D2O-Y/fWS@X]TZ/8J<&;;YY[b
/\Z1<?3Ff\&e[0M==M-94H=Q,06QQ,=^D0/.7)IJACEEV;LVV=SR^BF>FX/X6P;D
@W2Cc60.Y^?2>/Eb=+FXLcY#A:>a=7CX^[([IHZa&T/02HaVb)X4VdGK8L^JL4D=
4@EAb272=?@<BT\TgXSUI,=;E006c4<5)>4ZW@KJ>[=TIOVG;fAUYV.U?>JePBg1
M8Z+BR9IYJXS2&_M4,@YMe6-;4FHY/9V92:fcW>8]3^a0fD6]46/=X_6WZHIN>C;
^\Oa,_b9,H=O>_;K2Y]T:AWC+NSd2=SH&KK?J&^V&/C,A)]+0CXb0Q7A^Ud_9FO&
]R.9eQ2N:DTA)Jd]\(<=^.BFT^#[c,4-L_+JIe+DU)>Ub>KMQVe0B?JTCZa;bbe)
]ITgB^R.2)-g<&M9^EJDLE87S.GQ]^?fbXR9PJQbRKZK\V=KLK=2?f0ZZ50Hd(I\
D1#TW4=Kc&HV+&P),/<HEH;-2HS=?aFg#IcbQWDBJ^2ZOBNG.6F/X=a/Z>b27YV5
UZ-b<Y&TYTP/(3:F86a75L3Ye:>&@NB9DH&W9;>IN0;#BJ,/cMS@&-P2FI8C>XK:
)@.FPY1CW.F-1V-cgd.CAIM5YOa#2:HW9IQ43cJP=DUUFH+YXHDJTE6Lf#.P]J4K
V(9BX#b0cFMSE=2MDZ+XbUGAReY5OXSb[ba_#HF85?KcR1[HRWSHY4I#J^E[c;b,
SV_T+f9/12=>.N#<[?T1fd?FY<0dYQDc66TXeb^e3C]M^TEeAD)TK^g?28gFQHe7
.ME0)3BE>K[AK9#A-[RYFJ9Q_GA0-3DYVYd0(XPL=#;TQ.YUS4>\fK)\[+/YJ;+J
+ZZ\3]XO\?3,64+.B_a<R.#OM[fDH)5DC(^MIKO?&MO4@d1>0@XLC22OVLP^=45a
@UMG94ACP(23Y7FTC?4U0R)D?V.d_G>_;:LGSgTK0)=0U\O&HBSa5+=2;6I,BAS8
.G/JF.We#7_0;6,7eHL3A=QX0)U3L05FJBHFa,73(-0L2BQfWW@QV0d6()M&7#[J
[ZUZ0aJKca+.X#XG)-bbP+GIF]OME3>AG5fH;&XI3&1/<O+511JLI[[e3R?dYWV0
]0;QN^c\>S\Tf=CE+R5XNAAN1bgbY2&#T0?a4O#OW5R(\&4400F45c+EXWKOf4\G
gK[,NSKN=?-#)E5E,@2K:U-FdZ]S>^5MW]ORV^.<@<H__RU];JN023aYeQeG0C?f
Z:\&R-DU@PL[.GEFWGW2+&;;9&E#A=HB@)]Sf>G3GCAc3:X>fT^RT7([GYE-5W)\
<]XH]YL@W#T_CVD+4HRI;31S2&_D^0=>YWVF:0B,Z;HQWbN(>O#4I06b-Y.8CNeK
3<\4P3O&MYCYE@NMI)S.T,_>UB92f398U6<Hf>T[@VcUF=V.f<g,T+&b)QN;&)N5
c<NOZe5gI0f_^DBA]#,26GFRLKW\d?e#>AJF6Y>BTS9NZU_R8&D1)HFLEFRAfc8\
SbU<@4;?M[I8#UGb#f(E>B^LKbf;O0fM6CgGUSQO;B@OGCeN-,/WAMY?._/?KWa1
Q=ZCac>K9X_D)9[Z1O1JH4U4+LGad#(N#0YT8#Y[+J/QL:?G0;#V4H0g0[6;2+c.
61G@U5RVI:T34KDDI-6Q.b1=Y[@_C3Qd6P-J(,SB4>VcbE#876:IC[/2>L=?[ZDL
[3G@E5OW0G=V^V0CfKVS./2MG1\1O)38I+AI,NGIWM43QK<QSd-FX@J92-0?Z_cP
O+?=]>(.QBX:CH0_/]?4^]-P&5<V2T97^H\/S&^94-/(bZTF_;7PKG+^b<[<T_ZP
@7TBE2>ZDbS..I@9WggD?R\ZEb482N0fF1ZcS98#OOdOD9[#CNN=?(S\KB#(^NL;
?dYd6/K.)D_<^#<CA8]0I>/2C(cOW.4J80-Q^MI#Ue0Q_67[]E\E6UW3fRI:H:c;
PWeIDW4]DW[EHb;0bF6)>S^=cC>be:>)#8W#QPc^]LG&CDDP\Q@GV>PXJRLd6d0(
a7ZSLg^RCD8Fe)RPD4)MXW;-ba)#?ZRF&(P?4^cL#NP[UgP1g_Y@AIHU11bV46DU
1WAef_411]b[>OfO4B=FH2W<5]XcK)=I5+#-/&E^,_)7WX@8#WY?S2<L<-0CIRb^
N0d#[[?U#\&L^V7cZa=LS3Id,RXP-<,/&?O-VZ,>2)W;If]W2[ZeECHDc&E&W1+V
=#.^VX;PL6\U7EPf(39+U<HP<c-+9K?3,=T8N2WWA;SLMNd[G]F(/B2/6EOc4#U<
1Df@@6a_T0LE:PL\.\>g@4R:^&]2?_(UEKSYA7]+bL8RX1P3dL=5ZEE0&D=.T3aG
::P0>,_-46@KX\2T:TZ?c+M(N.>g:(LKE8O_.18YHOMfEfg.U^YLYcOe4?DDQ8Hc
92_8\1D^PL[9&-33UN]A(WWH=]/G5.=83APZaY&b25DH@3KCL6,],N>6fSV@(&NA
3a5C)0Ie2eAMDW]KPe=6O-J#gf&:PV]Pd[=[dH-0G#/__/ZC63AS>E7aAO4&_(=T
XRea5+FY<bFW^-V4<?N#@P&=X/X0//I[dVf_FC5]G2VI5aM_3aEA&K#8<cI\gDP;
E/;4TD7[QCC7PY9E)ZHGcGLFT1)7Z1<#\]dU^R/ON5=J5P5d,8Eg3XZRO).QY(\8
AR=U?/P45Y2K>T1D]1fd2-=31:GOT9@69M5YR>]4Y@HZ<bUJbV#U7U06>IJIGMg4
3(_PR^Ba6)F4X,e3,I-[:GPTZ\/+4XN][,8882Rc3SBT>RB6AZ5gH2<J<,e&.1LV
/PTWe7Od7D;?M(-cZ+EUTY]K]/06@KGBF@S9PJ7W&=gQDdLGB<L)eNUgKMg_Q\T5
X_8?IO.eDAY5GRGWI:33N@]:C8\X0/YO&C?HKbKN1O1O3,22(L8SQB,D0[(7I[Ff
Z)BT7\@02_;X-59f[:eNcNC].9[Y:EGGLWNd,PNS<[g-\&]faCRBRSa]Z,?eKcTV
;/<egK^V[@gGX<1>NJbNL\@ZNGJ:28:Bc8Sfbb7/0_WRf94MTE8dc77Jf_G#:[1a
V4d8cAIc7<,82Uc/I+P0C6[JQ6Ig>),@TKA;RC_.9C9cB4Nb,FMbgTe:CBE+MLGe
d=<4?0/0(@Y.O))I8O;2bN:A-_2JdE)>[:L.5cVWfJYY6dJG868N=PLMH_SZDeBH
YKe^K_@.?_LE[\L+KaDL>@aZQR8b_NV\+a5PYK=/C;AHNFL#E^P[KNWgEH78<65-
[2Z1gQ7YB89aWF;PY,UHf8NNFDZXX_gc43]dO)T>)dQUP-bPGKe#bD>OFP#XUccG
Q/HS^J9/=.R2C,PHc>ARZO.6-.6.7bM=PF0f90R&LOB<?9bA&D#J6VV)-FVeedQJ
BWLYOPcOAa>B3RMC;Db1P)5Qa@U?-L9G0L</J@KP6+aAN0(b5,;8+<,aIEREN\#4
M/I?Q3ZHP?&CD_<Fa(>R#>L=77\L(QQfJ,97NbNM5LS>]F,ECF<Qe)(#VMI@[Qa5
?bd-2OW0SUc<2S9[&aJd;]YKD#VU(a&NEAgHA=F:<6@ZVQJAA55e)SJ0/8H2P^II
>ZS6c/MSAM6Xf/_?+c[NO+e@3G1TU;&/(DJJ3A?K<[B\[2GE-Y9Z<BH2?KM,f+4@
XK1KZ:aO\:0M=PZc)3@a[H#A@GW&WdG@\)^D5XOF?e9bW</6Fed34ge@F6aTC6QD
P5,e4O7W>3R^8<B=E48a80M]Ra@C-S4.N=W:MW1DVdc3<\LKdQ<Y=U2G/8NCV(I9
^2PUBL4.F=#/ZN-FM>XfP#]1d>)0U@#5eQ1T)=K]&e&@?LLCCd/+YQWFBQYb#=a6
a:R-O^=JDY^UOO<LGdNN.0V)+MD=G^)NZEZ_bLNb/>HG1SV\Y@b/1<1X_T>JOV>L
\),cGIV6O8JSL7DD4d-B0[^1MJ8BOAU#T8?NGQVGGMV5S)EIC@HW&123e8FQ.6>Q
g9[eF2-SY\5B6U_P^;Tc,J--]0[HI#f7Q7@2#\@)?G-LIE];8&fZDC]fE,HMR[IN
@YcbSP3f8XM5(C5d#/XTMg:-cVXVb/1Q.2R@<dg(Nc+#SFQBdZW76bE?S_,+E?-4
Ag[]=2R:5=C4-9g/gY1@6T)C^CZGJY;\\LcG>:L,?X]9?FV-GJ3bFBBE_\0M[<GV
.KWQIUYE84e4bc<:E9Q3[-YM=][Nbaf0PZCYfQ-F(LHR]?3A=b0Xa^II#R_=#GIB
^gG4/9aI+fT)R)&+_A,^&]LJUSB\OEdY0O2^LI4-eR,dH@,9c=Y\\U@L9>aW=d6]
f779&C_^8WMcV;G.67/^1X&#&ONB;(#2YIQaR>XCO)6.YI.)FW+;DI;bJ16TN6R,
<Xac<Kcg_+QPELA(2I9cH<P-S[>OD/OR^4ER4YS[#4F)Ya^K.XF9]d=]IQ7b@9W_
F,,5##?);1_d>C2#fF7aOd#Y\1VG;T0>>N[4aZ\ZgY(1V=U;.LdDVcgW?=(c8S4?
efK8)?Z9Oga,1=P[M9<)-KT5H&TLZ\/Pb7U4A,#PM1(We<Z&<8T11L;M>db@1Q#1
T1#^dHdQB@47\\5?H&@Fb?dQ6R^VePG,XOg?faLW+[UYJ3X;PXJI3;RK6GI^T9OL
)MUK0.:;cf\=U?5L^)T1RHWBg\<:&J;KVP:C6ZX;YP>0;WGe^<T@K566+B-NQES2
&@T&3bRZQXRXdO;J5YCXZRW3VSc^8(+b,M>_.Ie\XNe4E&]:YDI]T,#AG_W9U,#)
2LY1,4Zb94PUc=UBG9>L^MWbHR2:g<9#/FIWSOFX^NeC@NCYC4)>OC&4PSMbS.Ag
CgCZ6,M&&F:,UKX@)Q@Pfc<bT_^;Lg+G<LS1c4Q_3YWQO-LK>IZH:==MI(:=CCSW
=;3.N-H<5e;2]\@&7Z8T<[FbdA<.D9S=FVGVC6b9bBKN=eSR245SgD:BA()+@Q3+
D4b+D1Z4N:?+:e:YBA>KO4g]Y]D;T8HY;gLF/\?:D5U1OB<5Q?SV,=,S;\1^>O\9
@:&4#4eRL&1SK1X/bS-_Z;5H7UA5HMWBb]WZAL;_QP6KRS(6C]ABXf=1.O&eMOVa
Fae=:GR&C(KIIU+D;4eU:X);BX>RbY=NXdT5HZ^[7)D6RVda;b^bLG9DCHaI2@O3
M]9]E?].JW-&OMJeV4QNR&?5]FNOG\R<J6_b\=bT05e/E>f-bW\#aJeS<QPEW]1f
1C4)/[2G)gUMVJ-eP-UCg,B5])WVTOND+5S\8\2)BUM:CS328\-e<?E9.0<CeeZ)
?>acG6V-._&@Lb:dM60fE?+1dAIfZgC-[J\]P;&Y:\@E6RBa[S&R:B;faX>1\\aC
/7\+D:WT.&;fd?<0D@VL>PBFJgNUb3I)c;<[EO[\6V7Q.5X3-Ze+4Ad3XF42A8L(
@-XE&eb@X-,IOU&YPOEX9Ne+gEIZ?O(bXBR-/19CZ]d[73fGWU@IMcTaUdM5&/LI
R)+RFN?#/0L[25dF6W?FM;[<8@fVaLV7GKV._^#+/D&_g\<N88M5_WaV,+G5&N=K
42_W(cUcI_Lg_GQ3\85cO1AQbDcFI.R/.SSeC[3b@>3g>-@:A<LOU\0<.c27;1K4
?569=+D6=,?eRd1G)F6&7U?bW1JA)cJH&0Z?+DFY&.>aCa,X[-/TDf?X;E\?GTZ6
X22?gKXEQY&Z78>?F\;5W^O>PTBc9(:e,:W0Q>C)JdG(MFIX01_abQ=2\/]XY)L,
^WWUbM>SaPO:b&JNP_6Q;/Q,8A?72T-ZcO;F^8:C^U+eXDZ9<CDD7UU?Q\&8;b=Z
BKOb;<MCB@#5b(c=U<KaYa8T_ESe4<(a4/Td:eX\-^J>.d]2g(#U1X0TAZ<RG.,]
.-FA=/X)a.1&@TC3Sf3FGY0S:MYZeNAJ#0:-H()?OcZTE;P<+T;Bc6UXe[NB?I3P
.>Ra73PG(O3T^;W,^;S7_L4:\-:CT()@)U?)TA9[ddGQ,AL>8R3TaA52/G]Xd.CY
1ANfecb37FSK.N[FT)6YFaZ)gIO0FD[DJ:d(>.;Y]_+51,C&3(D#a<T(LWGPbMW6
<VX>T0HXM3VU/O#6?:]a=X(LD[NA?Q?QPdADdX;Qc^)8&;QM[_feK^<2a&+:NGA:
D-+gT@W8&aE;TdS.d=JdgUfC<?eY\Xd8K3\dCUORYe:3R+F7P-Xd&PC=eCEgd?P5
3^0XV23,d9]U)>8ZVZ=TR(=g/Z1&_G7gA3f,+U]GF]G(H=#U8^>/Z=(Z65L/N7]H
&\T829+T&X+/fb,fS<Sf#SQ#3HYO:G)U[c]eGW4gB[-:99>.<M1.:fY;CU,=_db.
^/dL[3>&23=@Sg:R38#Rd8c+a\ODJ)Uc^:93SE1)c2,#-8g<YQAC0<F\PH/R]b9<
CE05Vb/)4H/V14J,IGH=V-_U#1)#OYOBY_F-eaK=+7P551]]\FFVWaNd3QFGJ(Z\
cfF<JL[HCEFe>&8(.V1I6+LIDGJW9f)W/4\Ke(M+-P3C191\G7EVUg3fC(Y]]_F:
7^6U.XeVNe:9;SfQ@:I;3DGd5#>#VLWK=M.U&&#0]5.;,B9:NW.ed>;R/#:YQ].Q
c(KOK-eH;3BM:00J+fR\)=5HDPd:RZ>\;a\@CCD1+GNR)G7;]5H7.cVQ2&fd^JY\
-dHgP@L5=4[@#F5Q3NXVcTGT?E.8@QfTa<;]WNEcD7EVW>A9JXd:1.d0LGQ&S(G7
TH@DV?fUb]5TeW\KaG>,;DL0)#(Ob4=f=5,S+B4#+^E8(TbFS3\V0#@-S]VB0Gde
]0YbM:WgYWK_+7TKLVAWDV6DI,[PcT=M_YG#,O^&O)4=Cc00fVW40B=JOR,Db[S(
:W/B)HDYX(?]4Y<#.74(WU_)(AYSM^>E2:b+5gbdTI+eWB4TfKgaA_^8E\/BJIC<
:BY+GLbg8b@_IMd619MO14P^dPIQ#]Q^9)(eC:0Xe.@YZ;EM/C\&GS]MEEd;g0[[
B>HR-\J(&Z&Y7L4[VK:=WM\7Rg9Y]#cJ0O4L#f363]_g3MN9V\(QVWI=NP92NHYQ
edXeG(][2B[[e3ULM[\45A:UQ;)ZABBb.[E&R3Ee_BXEcCFaBF.dJYCREHDIZ67e
L/4,Be@833,W\\08=[=H#Ra-\;:BT4S_&aBXU9E/9caPZd-PgM[B;77>A[(DQ_YW
]N2E5LVK92g>X)[O^5?#WH)[Y_;DKO-Mf57?f5>UFC8(4#F#Z;U_Qd^L;T-55Q8M
QOgW?Y?c2Tg.5;@;70O#31]:MX-W_fC3B?WSJP=@.;0(D$
`endprotected


`endif // GUARD_SVT_AXI_IC_SLAVE_AGENT_SV
