
`ifndef GUARD_SVT_AXI_LP_CHECKER_SV
`define GUARD_SVT_AXI_LP_CHECKER_SV
/**
 * Class declaration of each of the error check stats instances using the 
 * `SVT_ERR_CHECK_STATS_COV_EXTENDED_CLASS_DECL(stats_name) MACRO.
 * 
 * Each call of the MACRO would declare an extended "svt_err_check_stats_cov.sv" class
 * named as "svt_err_check_stats_cov_<stats_name>".
 */

`ifndef SVT_VMM_TECHNOLOGY
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FmVZMLXMmwRFzEVYDohHf2J5+QDO2pbArtrbWpxlNXEsdbCZ/nulYwGB4jNsRlLj
3X8T3dCv4T/pWYwlIv7lKMJce7N0JxbffRzwzdpJj5qTTxMWIGm1x/KSE6NDtscc
v2FmaTV//GW+bJSR5gJ/LI+OGnr5/aCBd6r4NRXj2r78yZBA7iFy8g==
//pragma protect end_key_block
//pragma protect digest_block
8IVu6vFoTPULBEyP8mK9L0aWAD4=
//pragma protect end_digest_block
//pragma protect data_block
3XTAVM5JzAV1eQ/jpx6uCwBH7LkIB0pVydxOFFOFqJrWELruWOi16SiXkUfXMotr
4tkXuvPy/iWDMvowinW0mEN3sihJlIZKl1sqPbT2CBDlL8Lda+3Yb7wH9E/DAer5
czOzXcio/XEf3B2Wi7fE5QUbW39djCCaMgOVqoXEKVXPcshgEjp5HQY/k/PPtV37
vtkKN40s/BUcg4JnCeobtZZDa/zUyIHpamSFIILNrjQ1/vyrKBauNZbYVonHNXtS
59zPKKrSgGRD3k4Z3jDkKfaiuiMPwHAbFV1GmB8Iv+hPjQ9kFkxdfTUrOWosdmX6
Ub3ymwH+U/LTw/Ay0IvpOUPDTDRJ6ziNPVWPCUQyms2Rgmw0ZeMAFgcZseFvePxk
9QgEsnvax7zxbPTpcL6tzyMoEww41fVKOwvzv1GokZbEm20YWAq3DW5XaIkHQNCA
tcchrm6ywCrS4eFK2QywZZZW86FRTAW6hE9aX1q8U3TiL+bnadN6AILWQAB983YG
BIUs3w7Y4mhCQP1Ou6YcQ9Yysxzbyoz272vbfVzv46xIIWjIPCi4H4hySeB7IupZ
xzAV8B4JdD8399xWqVQiMqOV+NDmqNFtai+GvwT+JwucaMOfD8B6lsZ1gQ46JUKp
2SS8E5+o/xkmtkpGWjdGuh30sXMo5EyV8333D7J167xRF7EEUE52Yv/agr0LHcjs
L9njqJvP28MFrcivsOjlfnbEq3mA7sSXR1/1YemLuww5to7paO2Ya/vmMOovyy1c
0yMx1hWlsHlbO1NAY2MN8lTB9QoxyUwfK6Ro+XkhRX3WEepLkImdncrn3Fq0YE/m
EWVSx4TE12JJtDqiQD08p+zUjivnT0G9OsjNl1Rm8VkC0eEmldsN6awwr7PLwz35
POKlQI+uuOxsralCWDsu/pSymrbltOkvYgyhzkjm8MnMJ4CzhVcJ1T+Nv9v/6GTV
3hUj20/7hjvjeiA5rxmhkCMPFdVMtLJ40JQ2evY9FwftgOyU2cA/YJJqFOOJ4Glk
jAs/dEXZa4R9R3w+jL/BcRvmPwkdJvgtNUvBk3bo0P3URRT8vrD1RI4uEZZtEX6H
LFJSPdU818OxjndcsyrP5VCRFDTJUdeEnGlH8HUcfqzz4vUiBT2zvKwGtX5555HZ
F58PEXkue5xBfjieSRMuz2/4i5antzqy0PE2ogh3bRlS7BZC4Wh97pgR05zFcF1k
WtlnTxx6UcW6vOC9hpk8GawBgMBCUVK1B7sEmJZ3+ckahjN1vctIYP1Ja9pr+3mR
UDKN4cx7oom6nYonQdI/C2x0KZ/ZOnWGe4cXjDgvnkuYqVSune6G1pD/bTTvAXYC
PzVNKYC0Lu143gPaR97N1QW0dYPwDY2WjRGxTWZ0KPkq4TdA/J4J29T5EN9RnU/g
sh+ew2obnngBkLTK9R3DMxL7e1xYxJPidZzwb7ON5+rQkk8Rkxw9PnpM/FD3rr4Z
THeioltNydnsYc0oeG3ZCweC6RCUAWZ1Nldq9usu+OT3OF11+x+KK285S06RE47+
n4jlU7Da2HpCgS9ZJSKBBc2awm0rl9vw5A7qHyjtlMj2zPIk5yFMymoeri6Sy90Y
Aot2XZsCYpgawKYe0G1WT71RJiiErt5cA618YEYNq88RV0WJ4ZebCKJ0pcxtJ7cP
FQY82RtwO/YGvOXK889pUfliPVF4mJBbvshjVw6c/epN6rZyIYzWk/T6e/IHmIIS
moW6NnzyIJoy7dXuYha3OzGiLsZPy/upldky4Ot9Cb1S+jgnmAkdY0xI4lfueZja
eCMmQ/7rZogGbYlRkiCzQSE5bpUh/Ag4vcPg00HXn4iVBPuZoZ30ntmCLiVUFVWo
suoXEjqTwMRlxkcRm67yBlz8pFVMBDqlUNtYNKQuoHKU2yUGg996OhyW6gCScoI7
oRelW4SwYvit7MYEhUSWkPE5pcdqsONkKJ/81oo9/bzfuiedKYPsl1FOab6G9oFi
POQHIZfwnE+9AgpSmZC4EOSal8DuUymv2ycudnFD6RTACL2WlPkW3dHOI19X42JZ
g0aRZGZmeKYbwstwfZvZBbLg5mNwPeuimRl4J2HPe4JQzmhapvhAjSSlcMKP6cvF
R6xdoA3CofQG7hm2m5fm1bdszUQTunmXqHInPar7cssoNATosZzaFlOiOoqoCi1J
IWDf72Nip5kFFpPyDmKsZA4FlevL3yWwlr/0CzAeHT8sOfP9d4BJY6ZF1nmYpV+9
hgg1BhXpbVcNFXeflDX5KWdcKVcLQo3qtVh37NS0yFg7ac9WVaiAl8bydt4xWahT
k4nUMhVB1Rr0K5Z2PCxGS8Fh8nniNzi7bjhDEGPpHu0iOJ7Ct60IAq4dv8qVz+3L
XyDVgmys5EA+tbfK7unR2XpkUtia4oDaXS1o8vhnxJwq8CuWlV5LRPaxJODOd45g
6GE4ti6o/Srn58M71/D1sv7/3XSjCNxx/rqL8tugxmySPXjY0rqz443FtpTWFA9k
9gVFWR/wikCSfg9FwY759CAFj7UK4xruPqvEmc3PAULVqXF2gn2XHDevYkwgVv9E
9/RyGAXPmBRoRUY3yjtqN8lynm4CSeunMzRpiz6NcbG/fwRe8UXlGyJKzYkpqXQi
nR8Ags4IK6/gL3g9aMdFJFWUx3WQK12wFlL5qLR7XvkLay/C/qG2hmjYIVVJUqxT
oxeBTSOZTXs+rzAHHoxqzg3Qao/etTMUID5IAQ+D5f75JE0JrKk+qPGv4z6SNOBO
o6gzSqcyUmPw6lgl7X8DKy/yg7W27beZOlJLhs2uox7ddQm0JzcPU8uyCl4Fe8Qm
kGR8rY2Kvu+nfRm8PQCnTDsFzdtec+kImvfPmQSXDsZuv+Vt19T4GwDuJKhXe7j/
EFpco3QJyX8b8FrIo/MUY9kkVFKHxiEeWbam9K07xXrQYkTGZNGWzYN9UjPYB3eS
KZUpB7n47gCmyw7Nx3YVI6o5Tl/CE/+I+actiVuKWrwpQ0jsHUTRxJ43XTXB6Tr3
oAq12FF2NjI40/2++ugyMSlMvXhNbZfJKblJDjazH1DbnjhRA1iGt/Zr0qX2BuuN
DmEdG54zGeP9Xc3sx0Qq1Ub/xC9Wjbu04JuOfRcas2zooXZAqJwgtx8RPeRdCczS
qFTTE7FEKtSb5n05AssQ5Gvuii/5ZZdfHVpimyOmY2y1e2u5ky9Skux48N/VCSXM
UFQOSx+ulCBuXCk4I2Oew0cRxP7eCuoPBDpq9rppEckz1+SD6jzLJk80/SWGUq87
1FfiJfprqhxc6Ap1+6/YqVYDAEmmBbSk1nB2XILDqBPmE+Z9uR4QfnaXAmcMNtEd
8vmKlChEzJ4aDlok2cnxYaS9QRnAX6gEyfAjImC49DToaaMS0CEGwotced0WoMPx

//pragma protect end_data_block
//pragma protect digest_block
2P37aD+hjvub6cFHyhB1jwaqVeI=
//pragma protect end_digest_block
//pragma protect end_protected
`endif

class svt_axi_lp_checker extends svt_err_check;
  local svt_axi_lp_port_configuration cfg;

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
n8eXkN9x0i3Kf04q075OmEPaJ1HXCrS/MtGVMsM30BvF+34+tDBbfPzovgXC35FO
U/FSMqapGZIOPO86oRnlmeLOWq77t+J4jPwdMrL1ykm4jNJnBPeA3+pwQiT7Br3b
flChj7Q260C/eeXQRbRRWwol9hZZx3/VOcQYYFcvuaNpAr6gFg410w==
//pragma protect end_key_block
//pragma protect digest_block
aQ9C9rA83surHrjNjif3kuMTxNM=
//pragma protect end_digest_block
//pragma protect data_block
f6o2fadNUNka2a1YyKAByxi/7JoxHrVVhDMT53BuuwQc2KwBpiQfLLeKe8m/MoX3
5DeBa8Zi1DV+gOvvvajUOFlXevOr8SWljVXpw7qZkwFg74kCFohqWM0J74vH+Ii3
lczkWIxrzzZk78PG5yWOW6vRFmetabYgMhXbOjjYtC3IJNmpFEgF0wLnM1XBjiWa
ShE2Pj6uAQ7K3a6xxV7yVkHjSxVh+0Tx1NffCbntFlhtvEf5DgTHbaYUQjLsCPjF
rWnCvCcmZyElqPijSNf60+YYTqdl8ti6gUrLaYgniolqE8O4Q3jrGqWW4QguTxue
JS0L2d5YvkZ1uq+wxuDTjjYtaqc5KN7UR7V8G7eMbM9chJQENVWTUzsIi/sOZ898

//pragma protect end_data_block
//pragma protect digest_block
X7ic4+8BDAYguyVlL6iscoGvnOQ=
//pragma protect end_digest_block
//pragma protect end_protected
  local string group_name = "";

  local string sub_group_name = "";

  /** String used in macros */
  local string macro_str = "";

  //--------------------------------------------------------------
  /** X/Z on the cactive signal */ 
  svt_err_check_stats signal_valid_cactive_check; 

  
  /** X/Z on the csysreq signal */ 
  svt_err_check_stats signal_valid_csysreq_check; 

  
  /** X/Z on the csysack signal */ 
  svt_err_check_stats signal_valid_csysack_check; 

  
  /** while entering into low power state, csysreq has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysreq_before_cactive_check; 

  
  /** while entering into low power state, csysack has gone low before cactive going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_cactive_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone low, timedout waiting for csysreq to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_timeout_after_cactive_check; 

  
  /** after cactive has gone low, csysack has gone low before csysreq going low */ 
  svt_err_check_stats entry_to_lp_csysack_before_csysreq_check; 

  
  /** while entering into low power state, cactive has gone high without waiting for csysreq and csysack to go low */ 
  svt_err_check_stats entry_to_lp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after csysreq has gone low, timedout waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysack_timeout_after_csysreq_check; 

  
  /** csysreq has gone high without waiting for csysack to go low */ 
  svt_err_check_stats entry_to_lp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysack has gone high before cactive/csysreq going high */ 
  svt_err_check_stats exit_from_lp_csysack_before_cactive_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_check; 

  
  /** after cactive has gone high, timedout waiting for csysreq to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysack has gone high before the csysreq has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_before_csysreq_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysreq, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_prp_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_prp_csysack_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysreq has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_prp_csysreq_stable_till_csysack_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_cactive_check; 

  
  /** after csysreq has gone high, timedout waiting for cactive to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_timeout_after_csysreq_check; 

  
  /** while exiting from low power state, csysack has gone high before the cactive has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_before_cactive_check; 

  
  /** while exiting from low power state, cactive has gone low before the csysack has gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_cactive_stable_till_csysreq_csysack_check; 

  
  /** after cactive, csysreq have gone high, timedout waiting for csysack to go high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysack_timeout_after_cactive_check; 

  
  /** while exiting from low power state, csysreq has gone low before the cactive, csysack have gone high */ 
  svt_err_check_stats exit_from_lp_ctrl_csysreq_stable_till_csysack_check; 

`ifdef SVT_UVM_TECHNOLOGY
  /** UVM report server passed in through the constructor */
  uvm_report_object reporter;
`elsif SVT_OVM_TECHNOLOGY
  /** OVM report server passed in through the constructor */
  ovm_report_object reporter;
`else
  /** VMM message service passed in through the constructor*/ 
  vmm_log  log;
`endif

`ifdef SVT_UVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, uvm_report_object reporter, bit register_enable=1);
`elsif SVT_OVM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new checker instance, passing the appropriate argument
   * 
   * @param reporter OVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, ovm_report_object reporter, bit register_enable=1);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param log VMM log instance used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (string name, svt_axi_lp_port_configuration cfg, vmm_log log = null, bit register_enable=1);
`endif

  /** @cond PRIVATE */
  extern function void set_default_pass_effect(svt_err_check_stats::fail_effect_enum default_pass_effect);
  extern function void execute(svt_err_check_stats check_stats, bit test_pass, string fail_msg="",
                               svt_err_check_stats::fail_effect_enum fail_effect=svt_err_check_stats::ERROR);

  extern function void register_err_checks(bit en = 1'b1);

  /** @endcond */
endclass

//----------------------------------------------------------------
/**
AXI low power port monitor check description
*/

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GwPHCDH2RLjRczsIgMU4fBA4iUsozeDBqSbDAgj49wPmwYwW3a2pet9s3FX4bQuj
bpFRuYtghmH/fHLsm1y6Sei79KouI9TkNZ5b0g9YoZXMQ6fbRKWcgOaHFBo3VZiS
sGr1e0XTTDxyz9M3O/rcIpgN5aVWwuWrZKZU6b19mFpzUZSddoLwww==
//pragma protect end_key_block
//pragma protect digest_block
arT20+Dj7vWlVDctV/dV10XnzgY=
//pragma protect end_digest_block
//pragma protect data_block
QMuHETJlp5+hhxhzyO1OWTFYYMyttRPEH/7P86ec1BQetTEESUHxBjj9WFPDuSjl
b0e8LE5E6Clcbb6IqWH/7tnyVsCTw9T2adH0gyOqp9eZjn2drgNdZIjxbchawnNU
n2FBW9qxQEYzaLGzZrSCJtDJalDZaxhqOLPauYgPGN+Z/q+KlJVX0F5QzBZzU3c5
EoaRMT7h/InW32ZSWIZuodQ8OiCw5Jgkyd3fDAglMG09XBs8fxA2IemqL8MWwwyx
K+n1EdWb+WCgymzKmKqcM4c62iakPfGxG8ajD98YeePG/Bg/BmAQrGetdJeiMZqd
dnIThviFYP+2XnLxGHyNXkHI6JHn/2ZhpZGxNKmBpSHqY4t2Viwd5jzGcnPQLfKR
Q2HqIvNmKEje8B+4gQcOMLqKvJ7fsok6sgL4aGgUSnFW43oc7tdEI0tgDV4xRGuG
RLdAPCk2QMyz423GH79otD8+cB0bYDa0AtTFo+xxbSYvi+8zw5TmCiaC0gCxHi91
+UiHh6wecRHpy8xnXGLYGUTzAZjyQTy+33Hxdy6oxYN+SBrc4ZCgCoCs9+MEMR46
SavyH2XieTtYHGpAEep+haMmAOYO8Yvcy2tE28lqd1FF0ximy1qBzdgf1jGLfrqn
yanqe3TS0McghMQ6jtzbwOc0eZsd2PNqGPOOb7ENExijNW1JhMS2efn9PG/U9HVh
YRwtvbZxOhmEo2onaH866iREvDWnD1j9+FPXciNENJiZzcKnOmj4l+1v0+ZsxjPD
DnVYBOYLdDCaXsNxN5sR+2mcFym0xkIW/fQ2BrSGjCvbX5XEptf2wZx7U9S/jzd3
z2ELYf8DmI9nw87cW+CVsLEvl7wXLecNEU2CbCegOWsekNoF8M3d/O5Z1WaNcyj8
UsqAGGjb4CoOzUgwlSUkIuSZbJVNp+3BbrCnWYA7QJq/jAq7uLYNb8e31ULyheW8
cFVN9x+kvnsXkjIA3FN0Dx+npYU1ajdcXRSTP698E8kl3a0W90cDHwZfCo4iGkd/
p/5daePfD1aDAS2Fcxq/20IzcrAEDDpXMmcJJDauK+16TLONld2gW6AwUV2aXJEJ
aYtFhwiatBI9IwSvptGGoKgtmSJZU6AlARREBTqV3Bw3KKcoJUyugVjZHW6B3CWk
esFSJlTkC4x0T5McHJAldUlWt+q/7BdWZN1hyBTmXaZqMf+ZWjjPXqOiXAnFd7w3
o5/t+YIcf3Dz0Qs0VgZ42y/xhdKdoJJ9UzKkxA+Whjd71qnkXfqRo9Mbt+rUwu3t
MTeXEBzxepp7uPXXvLZt2rqKRqS524arJZa2ihTYKHEre1h5W49GXmod/Et8Q+zq
YAjOlFs2BRVx+iQZvuxw+00D1nSAhjf+JpTwBt6hLHr1dl/Zj6FlQ/NpO7ZOvb6O
GEfS0iLn/XdMO4ba5FL8zd7W5TfV6VBsCxkjtZFw7ne7B55BCqgYSQnsRLSfrXuo
tN0XMkzQy8hm+LwIHQzDLHrrwRI1LTamAqApO1Mo/CHgocuZ6YYicMPEQwR38NJH
fmz6GtUwvfdUuaNh0aoUi6rgTO2Nb3ifHFdCZipdfcTtHwkY2YXdEw+jg41s2YZ2
JFQNyCe38IasJgbkUMghpg9IZwgwF/zFELFh9P96e9zuUjKlheZ77QbbkcowiMbf
Z6k5QlO39xQhYyG3DVPyxhuaNGMoQCwIgJ7/7DKGGXr7eyiP5ZIzvPoOTZZcmZ1X
Jr/PFTnUMRi2K0XWDWszuHRI2HLjzBhw15UzMa50eFUyjufvvfaQa2A87hsmKkXC
c1mw3if0zEG3Ga2PRJBGk7K4urTOenMyZUHERISPI1ujodw8qnmW4LnG8Sbt5We+
A2twGS55hExtkNx8qPHtNPkYcCMAGY3461kvxQeB4JrfUFNVtoMjRZ4bZJ10PsCf
2+EeOTrOMU5gWOxMF/Ki6z8fPxumsSNq42R5w5bChkcqbPjTBuQfWdBe6+nFIvVX
ZrFKuY1kizBPCxlzz4r5JGRX0mxDdWeft62Ria+TeWibiDxMITG8WHGFSGZTNxkJ
yDOmFxSjy1P5wlVrsjiZftNoF18FD6Q6K63RkaQWEJT2mfxPXMLiOsf8Cr9SFFs+
Z2SVbicMfis6ixhisx8XKp655Kszu/Rjc1827fL0Tx71Z/7H8IxHxpCYdzSFVhhv
Z5EaG1ovXvbiLCYFJDvpKh5NtWn7kE9q0WDZklQqlV0HeBE9YZnM/18O6GAPOCdV
O8qhw9p7od9BcT7h0ZYdzYXUN8IKjPA8/hZ8Rsaxaqc=
//pragma protect end_data_block
//pragma protect digest_block
ZhjtQwuGDzLZtA2Ns11It4r0h4I=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
unEVBICkUhsn8mwgoeUMmR3oQC0YYSusTQTh8Ds6lguWNQ0VN6qcFmpwTBPUPOhc
hbsSCk90fdEdhJisb/zAQUE2KbCL6D6yOPjGtTdulxifg1zNtZUP4737ofnMCnsd
PNB2cEFf8mV7XASQ0foXHqRgrO8Al3eWmHl1otwk6NigTdBLylTYtw==
//pragma protect end_key_block
//pragma protect digest_block
XoNd+jAei6MBsOUzpV3ydQ/FtvM=
//pragma protect end_digest_block
//pragma protect data_block
ZdmVMqzSaEg+pS2d9HkBhC2WAyHgUcnRp4X+HsqfyEvBS3U2Fr0by8g2JSwxDVfc
xo3yB6+h9SiCeA/4M0YmbieXsNB9j6VICjv4CyrpGoc02xAmhpDXE55l62O2HEoQ
3pbLWkvzO6xmnS6aAJrciXEAW07XD4ypXe3MK8sTSbkM9tZegMVYesPq0ZTfNDGt
9UA3uSrdBN6l1TFpVmUwkLvQ3U1Gc398jlXHSWLVcvEZwbSd5qpS1OKv/s6TEZQU
MnOtHjoOTFfekFPOCVf6CkjVPbOyuFva7sj2o7dsP3Pf/oa47/HgCC/GAiwoj0Bj
aasMitSBcfAw1DYQNKXhi4O5yORfskQHtFTahid86hnrTVNWCAFl/yDMJNJrqX3U
oPHuKASpaJrWj48zUIQSJOBN7cjgXfgK326T4ivNa9QczuODkb8958YfyXthH3BE
bjeTtV9fLHGvIuRVfU3PallVTKnpfwCdFB1FHkzeVVlPOhsLpH6aPUOQlPdEi47t
3RRx8YlzxokrLrotUcrjhYAshQCV5RCblteFaaqi0k6gS/xcJOqmsVBwViNYTygg
4fQXtX7g7+Gz8AlbNNV+eaJ3bdyZuPmqQKagba1VZA8qkEkxoKhHjcVLt97gO4gB
w3CA/jhBvLxVZnsMPynaPu3Xc6/r06IEK8geKwjCXWt8rKVLgqgXJt0JqUqPoSO/
pTE414LVwh/C9kIbD71HdqgxbIcPJIgzibXjzpCbUHVOG2SgiwpawJdEmfZUHCi5
eLPcmFQ00llLozjNpLzMk9EQZoWcO4vozLRb+vwerz0U4kWLq6RPcUB0qgrXv423
AcNQDomRMZZHFYwi5KOlGg4APr38j5fIjGYqFU24WvVkYWodV/mhX0Bpn5TGW8wJ
ZXFqLSyeY8z0ufpzrRyl1vspblJk8hh9sEj5bjysBNaJjsF6pGTJ0dYM8Nzr4fn/
XPo6UiiFS0sE2mEC0LwpJKs6qLb8mPijqdvo6n5sY/IcY6DgSS97sYsl7rbkBj8h
VYfdfsG/9A4TVFCsfjY6BQhtsn5BUfh6IDGZiLTKD90X8eDljS8h95AbjKpd1g13
6w3Vo0wqKY5e3k+m3xDf3qJSLMIToA/MLNf3ON65AYStwGj8MjhXdP5u/CkFKMB4
ScKJNKojvrZL9/lLt2X26mVlvFeLgyawiP7g6EINrVZ6nfi+Set5CvAxUl0FfbBs
1+kSiNxq8scGOnWFq586TD77IMpfuVzfCwPiP8rrAwklO2eHWJnI/j8ztTHVDIZo
gWo++6nZcNS/T4f6SFb6NJYlokm2Cw/YIv4ExF+dXuocuk4/tkiVmgwfhisRgjCe
wn4GDF8Xb7b14BANyjE91o+lByKC0S4iS+pHD96uf0gwGIF2/2hrvqco4v8cdOo4
nQM4EleBKwz5mRZzh4o4lDnXDUEUnQgIM6wsNBey2/t8CF2VnclteYlTF7Pikrn1
a9SrXIOpoEMLYIi1WWbt9Gs+sKD72wWnPtkJQm3Ofk+eNPzD3zYIfgp6443+t9mg
gF7fZo5Sw6oYdcjr+pX5cRkQEFLCmygXI/HpDSVG+m19QvyqDVKenZDaOgM4m/oU
fbPvKyPhxrraKCE4g7vkGRHBN7JrsC+UzdAeoErIgCCp8+r5nqP51HgdF4/AKtCZ
W+a+xYVKQxRhBygAJakOekf7HnL53yvfBYKUjvsKGWdMiIqyYNc2skGCHp9nFo5f
z5zj93YaZJYc5tQEvTYRHww+jY6dSKIYp0AZDwykdes6zpc8yqKvalYso/g2LZob
sW1ubhy7NtL2r+V1T6s/0Ttuk7YCPlm23K4itNP+jlQHWWo8wGwpD7qJVDeuTpKX
fUxYIyJldEgucnGx/Thh8XNCoFxyz8NrNy6hHj9lV3p99lNuA4vTDj3T3NLY8qVj
jsGp0idlyIGBl9QPEfjhx+QbwvPvaXGRQeo/BGH5bRx1U0L9W+qfu8NwYXXmaJqc
dpUhgXObGaiMTnNRrDNSlnlgSi1GvBF69A9JrJmE9unyGoJ6qNR41dynXwwFLYeK
KqKotn2S7gKq2of0C4iC6jqXp98S/2fgLL/AxxvbuxE3YqhEa/rdjVT8hTGRwD2x
jAZ6ppaZSRVNHRXOV1OgkYeFm6PgylX6T1/O/a4l3cYFya33yplN/cxW434ctwGs
QwdeOY4+7/O/p/SYWAyhkXyZW1mOubpdCwcEm3PRwJUVhdAR6BB4ZVA6dFr43tQ/
RfoytRs4v/qLLEAvZuKaxaYawcyhfclE7FgmjcTcImK98A0UipVIjhHWShzVQI1O
jmxcEviFz2nEDyTLqYPPMHR1+/LWWPTyNBf7cnBfLRcxgOgkUj3XGKcSbtfPytY8
1Fv95fwFAlmBsWjtaLeEz06i2F9rqam1bKP5GB63DAx/akrgn2wHL4pb9bMCCpUu
vIBKMfaOjiYLl9xKJqv4dpugA6YGajWAn8tiujrx6M9h+pW0Zd4sfkvEUZNCVXMn
Wn+ZP1/LkWCeIKdwunntccviTIp6a4dk9FKMNTeN5cDqZHPzU2ZK4UGQgoJA4Dtu
H94nOV/SoKRx9iseKzS3RplMOdlf8LOSOUMklCBI6aRtt/CeEQPQU96R8HXNkC+v
a+LA6U0UVIa8jVxThT+1JDtFgGrx98TfZIV1tqr8m+cUXhHGsoyydNSHRfOlONvl
1i5hbrJRZ0cdoXNhN7wCKBEMluVX5uO4QJ8U0+ZEcCkizMP2GE1Jrq/DOl2CAtMD
kN+0EIsNP86onjMUOrtnYfi4IGVHkJwboTBntLMK4B7NzgGA/tEMMYYi9AxkA8jh
r1rqoXKidkWVNYDKdgNvGHBA8k5Zahc7c2Lgc9IATssTRNsolRDb+KcXMhYuRaKT
6zoMTR6SNLFtYJGISn62OEeB6FdjU+WSkf9HhOMbqtBj9FNXEH3WPCCE490tQkgX
3nQLtKpMvNRYVG1o1hmlnyQ9l/NVPpLCTesqRETub9WmmOb3L8vCA39kKiz5BcKd
QuvvSMIC/y1GcaHQqtX8ZtmKPS3pPZ3Pw4BieW73Gz5QTXW/E+1fFwYt/s9eYIaD
KtzKrwgh31/D1jaJverUNZCmSsueBsO92234904bH7HuhiRFU9Ex+NluaYTRWb0x
rv9V0Wi4N18pCpU+7aOm91vdu9UbYdRP1IbG9X92CyH9JZhAVwqzKrpIZEIYAYS+
tQ/s5Ug5fb3g/0limF4+ijolGuk6XwrvgvMGX+v/7vmpNKCAhMJ3z7uSgUzdRDtO
5iDg+ZzQgqPLoaSlc5DdmujivuFhDjbRYmn6lfgsIxx6f40d6votOOuqd+ON/RuN
b1Aa2wwFemBc+TYBxtdo6wWOMPL3dq4XU0jIVOLPSMGSvtqxmTyxCTLlRNhBdgAx
InHYYru0YUPKW2kF24rHfzgCYb16qoaG4vazYlK27MUgiupi2ZFXC7Q4et97PHBl
OVgeRRzQA+08zE/7vu8FEJlKMWkFZX+z1JpYFIZT/nrw6FhauvMlZFhAKJhnOv9y
wlN6bU07lWntqBKq5Ecbvx4A+G2dHPKJmtW7kouW2pgLniqL9Hruke9k3HV4bTr3
aqBaOyjOA41SmUTG9HkPSXQLZePicvOwicZpso8Qfhwrb/gCrT7Ccd0doGWjgib/
tM+rCyOQDgVRl/o7QJmgEVLX3/jhAQd/IrIuihp8u3qfKO1gPb8wHqa7tZi8rstd
0TYqIYZQhPqpIlAzI2BNuL9vdUp1Gz7INQqp7J4SDZ+740DZ+PR65GpczTr0DhAq
Td+Ccnvt9XfXH/aKf20stpfBuHQmocN7ayvm1etLGgGCR1i8G2Z40NTV7QwpWlEm
dq8ijBgHYVfruCqgJU1RRQb5NXwswzfAS1EJogg3CjHCDOIizzwL8l62UJkBERTw
zJjzuHvnIb9BD3Y4ck0gCXOZrZab/Zd5nH9kSi2GbguvL1Gp2qtEKcOR+R/kfJ3M
Hj1rFWMp520rBkUerq1k0viwwW75ls7OrrEsSVsfGDV29dwYQJ4gl5Jg5DUbCCAt
VaeA4IyO8whVzTR4PXMLyLWyIsw49DDCjL2fJ0GxoDEIMRM6P1VXEzUALTQyczWd
LK3zFa+Src08glMg8akf/SXjGTiwxgFijrAFsih32Tw+iE4UDmPDj0oSP6k56iHs
UqoBUzixzf9oI31Kkjh0hr7Keyt6Qb7PNRQUIGlPpI0aEFyKV6hbf3Qz7lJDqAwv
ky8OwQvfzGl2m2eHBLBI/fBeYrbAkKi/AxKKmiPDdqSa4DrinxQCvGyVACM0AQ4i
Bo1ZhrpBN7EqtyyLjefYMBn9ivYVspUsBMY5lKRilbKJPO6ImL9gT6kbaK8VBGwx
8x7YbZqm2TsJjxz2mzygbxjGXOBkXjAobniVN7B35nqqEOKTsZXXX9nVRc95F1Zd
TcrjH6X7cnr3tXnAuswhC5JNXjkQj30pslAb4KabdqtR5Jf/kQAQQssbcPnQUyy3
QXBTt1HOCheWRD8S6kU7BM/NzJINiKX3gQHIRyBt6mAiUDpH4uP0U4y78H6SkLLe
MqomDAzzc+rw+ZESHBqcyVnu6dTHezAD4/Lt344uHJnR+WjX9Sxj5RqbL5ZfJX+G
VKJqb9AyFM9lVJhkpBYRcC7mQq0S6d5fLsP95GdaPU0Mve2DPqnUjATh2yezUb+/
lXSgU4UNZ7WdE94wmlVW01DYV3c0J8SGIcbmENWGKdKJYJxFou8tdZxqdb4YdwdZ
JzxkVK4hs0NdBiwXRoO8ljqnVS9NFo4hZeLzyYY/+KoeVKa5x2Qfvmkz9YKHaw/Z
coJwEi45E/Oz8REJXudKRYXxXuwlMdLDhALmftDaGsMmiMiPAV3RDuyRBW/0HBpQ
yNeqtZyLgcxr/AbewyHY+weqw9KIPEpiigtKc+MAUqDdxJABRVijiZiZAO4tDx79
gM5NKTayTv8QoSGeJ6iuO6jncHexhQzeGdgRsscRzF1XAOCj9N2ApufmJjhHq/NT
WA+G9Um5TEzhsYJ+GII3r+Y3AVUVVjbgnMyiGPBrlTwNfh2eZJ9lCjRtKO7Vm4lS
Z6kvZA861e4FIVQuyusuDEBT2gVfkMNil4m6sLSo9M54RXpSSR7E1qlTJIXccpYv
jCAVnoOG7XWEwdoZQZYZrcg60YIf0hK8OBRCWZ6lM/YhIhlSdAkGb1dncbbjVSSY
i20Iy2Nqzmnde+hDlXoLhB31BQfqtwSmAKb1z+cONQio/hcWzeGoaFOADqPDB7YY
bdg/TDERWa/zhbTQQ7i/I+YvS1RWqPZtFBF+38l0MtMBvOgR1outVAT+AnigVkHy
F3AsNp7tGi6iueuxzzTSrT56gHtsaOobcQF0E/iCkNGsluTmuzvhMEAKPAM6nQET
thSC2lGXQg7qkxlFWA/zJHgjafJn0smB2JbDrtTulseGz49ldvo85f9Y71f+LZX4
qxHE/CV1RHCVoe/WOm2fmCJkxO7alhsRGar3aQLNOAoq+TE5GGcdB/pENPm56fgi
mz2BNFPHCVpqPji/LsBpNyutf/x1fKraAEBsYzZ/jCKc09K7bcePGKoek6PEPhrF
lRdYyQ1N7oR27HuZCdZgOBnIhILTT6cc1AlY6gtrr2qKau1aWwK/JpH+eZYbiyhA
qmB8nfj0p2b9KaUk3zOqv0QVHJXXKbIyONSh/Er0BZNs4bYAZxVjqMf0krFy5pIf
J8t51F1iGMdDNAwP1fvZKf94zxgqDOmWKCcG4QpXPlqU9bz4uxuXa/zkwnlfCBGV
syvKaJWhdUursHSr0cs4PB4hBVlyg4IVhLSYI9/wH51O3ZLKjVaSLcR+eKH28ixO
Oeuw3sQRe86bG0WFQmxGT+u6jsROMZJBLmysZeKZtAAZDgIZtuptLoCU2CR8hKWr
S9EAV2dF0pJ6zQi0SR+UdQS59t5yjaWF+U7DggVqmxscRE1MzNecfjto2cj8BBs8
y2L3n4x8Rp+Or9yIZyOp9PXsXpMwAZebQVa1vtbPohSuI9iBIBmmhbwfiQ6YSVUj
QRZz+XFu6daxLsK446DhS3MjSAjG9NEqFAQpxkyr9fvD/bBIt8bPPhPv5Sxe+UQz
VjMdKEeRfW/SJ+lZuY0FUNlDVkJxriY1z2yYTjkuX2rsRSUYuW9reM32NB4DSNQt
Dy+0qzESYQsSdiHrTK4tvSsJ8FI4Er6meYB+ENr07R9sYP0XWt340EzgydxND0rp
nhPDFnrnVMvNAMd+VIEPJT69ydf9Iwjb8iA5abVatC/AXof4dxv8TC+ewaiLQQmT
Mk8aRDTz2RfOTpoZhw5ccYq8hjooD4ZEtL3QItmG/InwF9HXImDqLEGcnGFfo27r
Th8XdI8d4zzJtaoJM5tzPN5m/TZgN/23W4TQoVbhyykKDaPivirRt/BliRc3oiKa
4Nn62ulumvVi19SW+axAhE6p2M0n0Ki0Yc1n6iksZ4Pz9/2tXStKF388DyKKILyO
2BWkZlSpJ+NOAgur5IeR3FS7llJpZNAU1PwuKRkne8DE1Hj+xE1jhQGQnKRSR0og
jL7QTgD8jM+2hZ5xwXoboSfDXXXP4dbK0LOrClo5XvEv1eQ9k7s2XHkubBFHv/0h
2geLLm7y0qOSJamXPz2KBZ+tkiK2UkLfWthnLa1SlTIcpbjZ5qJi8c53svzvVIJ5
vcU3pMzC0mYLKL60FVlJB12Wn2UwFFk2Ah9jr3GKTJcy4eK9pbdy8MTbzB9GceoI
53wPJERf9W/K24bxt2O9IeyEfgiSClzXZohVqFJO9C3J6P/4f9n3GYeM2rEwhcZf
ARxDQ9SbshmB9eq75Gh9ai38YMfYTFQmOBMDSganjDt8XY4llBsdCmwU0n+74P3N
6Xxy3B7tzd8+9HGDCxqQ4FLxW1rRB41wkCcTndDgqQ5xrqM1KhsApE0ACLs+K2B8
QUnql/tTFQ7vYsEuMQL6l23I/oYHbKBUmgiNZrP42MktEtQm+T1E1GHBc/Ku58d/
KnnnU2SewSe6U/znN2t5sFt4i1AD1Ne9SgWJ3I2ix1WAVIuUeSDpzd+TkbYKmoSa
U2eGl37t1FtArPPp3WNyKeBlZGloIyQsVM7gTiZDZDdhgI5TqHAvHATrqWRbRPCl
opVxxpqKT7vEyEe8Q/bc4K0DjSdUkK5UI0hoW7K1dyccik7Yyf1fzL+0qyn4D0Yt
5q8zm9D+2WRSHdEX9ixRQbgpKIbabdwpkWHXTHF/e2+ZFxVcbIKjRXfhIM7+g7hp
0/2BeNVgxwlWIHa5G6f24K3tyIESBz/ooE3HRuZaJhXONlBWKvH4zJL0RXA1lKnh
OEbX5pl+zqbUR3Qj3SqoX+z+JXzQsdr3na1Pkelyyd1A0z7gbbfmfDAnLMvZ61Kv
vqob22gcEKzCA/jeZvL6zdC+va6Ye/yLe/Ms8n7P5KiX9yfpjkEyGGhQsEgE4lwE
u45CKwxdUp8KLI17Va+3E9cFS8Rs9zXFPjaDNPIDxnKifaFIflNKxOCWgw/rmv6Z
8rW1CPoBwDnwVimQ9gluU1X5Wn++TEKjWkWMJxvtDNakd8fuQFboulY7LYuLGKBD
BRL3yOxQYzrsSl1E+l8BaiPBiVwI32RI/bWgOBvFMYC6mX/mew9J38+LXv1XsjgA
3zOIoAkVqbWVqWWnuJUgajDDdUZBzt2hztzl6L3Z4i4Bj6rooas8uqNTmza6WRY+
5Kx1/n/9JFFVn+cRizqJG12gZzA1nP26EIXl3mOTBH1Pw2OgH4A3c6cAISBu3cnh
YgrWdjcMjN7qOnNHoGsBjhDgZNGSSKcan+z9LslHAjn56RqoAR4At0v2CTRrc7Sq
Uys/3PsL9WTK7LuEoVhJtToy0aIseLgtShZ2sMroUoSeBPF1nbfGqtAwp/DsCy7I
sNh2QHMXGz02xP36DI4QIHzPrMD8ILelmK7VkJ5SABVnyYyCcwIeyOR9PRaAFSMA
zikl4dGG0f5ACREa2qUm7Q8CzcDcYOgewFVByy++/qtWC7nrMpQ5m9UnDEhweIKc
GJjGVCsXYQWxzAxJZxNczg==
//pragma protect end_data_block
//pragma protect digest_block
jserRP2x65No1EHEWKd2P32SOhI=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

