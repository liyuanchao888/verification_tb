
`ifndef GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
`define GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
/**
  * AHB System monitor callback class contains the callback methods called by the 
  * AHB system monitor component.
  */
`ifdef SVT_VMM_TECHNOLOGY
class svt_ahb_system_monitor_callback extends svt_xactor_callbacks;
`else
class svt_ahb_system_monitor_callback extends svt_callback;  
`endif

  //----------------------------------------------------------------------------
  /** CONSTUCTOR: Create a new callback instance */
`ifdef SVT_VMM_TECHNOLOGY
  extern function new();
`else
  extern function new(string name = "svt_ahb_system_monitor_callback");
`endif

//vcs_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
aaVFhkO3lHsts6a/wUrEwyiBryemQY+1s/OTTA1ugO4NCJIHwnawqX1CfI/bZ+a6
s04W4s2PPyZvIlE2wJZOw9PWi2QTZNUmw6MC+NhiIuY8JnE5RFczhyBtLAaxgAFz
9S1SwgitlaDdbs3unmF9SXZ3aYl+0COGs0Jo86Lz1bYNQXPUP8T+VA==
//pragma protect end_key_block
//pragma protect digest_block
UsKNA2L70ia2wMmqT5XrTgEJHoI=
//pragma protect end_digest_block
//pragma protect data_block
zLdBGEHv0RuezcAj92GqWKfmTpbSYEbv5OMD8bqM5MPZABq61jJX3AmamS18UUzo
AlLYUaQNXdvKvpGemj9DEa8B6BphKVO3SfBLFJ++5OXwSQWaOGbuL6WevgtVmwr7
/s6BD4rqxNOAWt4OVldBJKzAtm4py61qa1vyHucjSCw1nU7lU7bKavqAJiNkWfIh
4c0g/A9TRr5ukvwkXZ9iGSRf7U6uGiMpa3SoqKrEKbHBUTD/XPrO/po7Hw0mja2v
i3aPKDw2PrEsb5lMUVmj9+4uwEc+Q2gCGBl0F/e98IZhd+3SNiCEgmpDT9L2JLet
BP37RqIbVRW6XE3XiKSInh24REBjIecw3yJoIjA7ZXCwqME7zGZPBu+8wT4vDoZh
mmAIKG8r4H8Ir/JUkyCzhVBaOaK/1GJFV4i+Lxjz7vxpOalRV7xG+MCsvYEZ9xAB
GX3rVjsZrKqwV30xxBacTCF9Di/rVyU+lWWsIrFVdDixTgu90cxe0ceCw61hYeBp
12bNwbD24Em/co2CCL3DYzE1VqoBiTgY35BNPQyzTd8w10wveFo7n1KdB8ERAs8o
8CYDn98gTkSUq0kOTxXNNGCxE3/QFpm5PlKV11RyEhhB4cuKFI1ZNzrCKc4AcEiI
QqFj0NCuC9HPcbVCKr4tukeKueHlDqjvUMh+2LG1k05os5RZeXMO2aLFXnqybEIt
gG/lxvrrslbz4VewI+QZY2RQ+SZmJ7z9J0d56J+DULET6q345AYQwBxbtVC8Z9Hs
sV0vw8KMafB9EapShqBqTSno9BkKRIc6up/Kph2sjG/6BrbSx8lbdGiE2lrExtsk
480SEVFo3gn/LIAmi2NTiZE2xOn0B0vmEi9iIPf0Z+28lqh20BNcI6rBtmpUgyaO
L6iRJoKcIrsm39ZeLeJ/zgP+yY2Wy3lkqV4piT+K/sfEogWF69fow1bzyJ89KKsL
i/gsZHrc19NQaR8RmjyGvE8GCHIaKcbSTemC/bW8+Eu+mAw05StpDAHY5VU3MJ1l
TfojkLK0/iK+/Z96UUYo1K6wYyWITqydmKfjJJj7BUR0GgqNe1A8moxvim7HIIkK
TwcTdwLSc71jIQMzmdoY9Q1GXFWUirKtabXMIyP7A2v1z4wn8AUtRfnHlc5eerQ9
4ziYMlZQPXUouqwk+1V2TSfQpfpFY9L0aWMUShNFZUqykCsN47NNwFxnna4fRe8X
Tk7znUfYSbU0LYOQmskNylPI7U6orH9HG8NNW1od/aGkdLiSep8KYpNTXlkEnQ66
a7F3RJwg1lIOYn6xPfHgKydQ0fIwUNpoC5MzsKWNbtn9i386iBV2rmeKbuAL7rdU
LRFyDBwGlnKAfofKFsAkTR1ORHbNClbr57taf3RrdfRGHl+LIjOUY2qKiCe0Suk1
ofCTF0a+UhA9dQAwPxKh0+lflb6YMPjDtLO3wOjBCXJhUgBTDvs/od87ZUE1vovG
IlHe3t6kSTkUgwYiwRM0E9bdA87fErGRyOgsWX+oBW6aJUhENuyPfu/l6o3xxaYt
4p58KVbt1BGGtFdq+xX9sehKN5sUlkjyrX3Ps4OobafhhMTCxEF8gf+fCUDB5cnt
o7KYROz88lSp4pymuhLbWJNC8Z0LSopFGbAQhZpmiUKT8snzFy/2ZWm0xRLyquva
cEJMx/v4Q/Zpnad81fx4lOT1o/RLYoXjKJNvd9Z77DiZHrvN+azN9lxziMPClo0h
nt8bnAIEb9yu4bfDNFG2uvQOBu1V7cXmitn0GLasOHe8W2UW7c70GtxSIuxAJOna
0sU+0Ueey2qUHf/JWonmJ95XDdNdwSMwTCmR1GtNcfD3redI+rEH9pB9Y4+u4TZC
OWfgaqeKOs+rCZwPN7YiUFad/JAYJd2fXrNaRsunltBeqxKajlT3ISTMWBUq3WKB
RcvJOyD7c19NC5dM+ubsUWt/WpLXTPfz2RWuX28QHvLFB2bQTbauNf6o163oYVed
AfGDCn/7Z3mmtYpiDHF2I0/86RSCu0wP/+wof4KNljlx3doR6HirV4adNUM9ZReQ
D+cCI4+wyrekbwiI6gZg07EF+jAU4CbgerrE9jcJN/+gvVBNoHYzLFydhcw25MhK
DBC+4V+kp6m9dQuGqzIox3RAhSDyQsjPzqYjx0p6L6xmS45kK9D0HneOnzDPelZl
hJGM27exaQoy4L/3rYh0BZDzUxQjfKoRlKPLkuZd/oeGAQVKQ0yGMNxX2VNd0K/x
q+eP11ytv+76iV5B8UXh7johpGLPkofsOuy3bycXPqYvXU2rjAxKWZMrvY3z3G6D
jR19pYGGEy9y9w+DfLVmBn3+Tr4R1FIRPl9VfXxPyrjiZwFUyZAcJz6V3YMe86Jp
pd7BZt17aeH0bVw6XVynWi7ISVZSFgfGUnE8Q8PVTmXErMP1Mni9fhqePbrsV0Sd
a8Ei1zpIf/704idvCjfo0gUZEAMKjUpOHLyw0YM+vrsi0LnhbJ7nHhhqhiyWyRMc
gKvwJht31ugjLxVqhl3kV1kaSK7J06VkDjzzGULwGXciJG+1Xlk+YT6heCZERKhc
ZPq5Th8RJS9U9fBsvt/hu+uxgeNumugcmAG2e0P0l4KLvn8S719uAywsRlsBjvCo
BNrgvZRVkw3X918ZwYiwgFatFvglu3QphHv0SMrp8xc6/4iRQE1Xwn5+V9w8KwDe
3byUXGmGHuOxfpO/y9jHpA==
//pragma protect end_data_block
//pragma protect digest_block
yc7gYGrRSWPPHby6RYMHM1jcEk0=
//pragma protect end_digest_block
//pragma protect end_protected
endclass

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
8ea0whVPrTsTJKmsV454XgqsK4dB6UEz2W1hUBlBhTvUFpY4kPfSzbFduspKamI2
QbmbIVVdJt+3eB2JniXH+r0olYfKRHEY6rr9sPeRGO69BRwu2ik06HWEu4EDk58c
GQPwImcLpSiJ2ocWrYxhRYcVLI6W8RR0cQ02GFMSpBKe7WO/a5grdA==
//pragma protect end_key_block
//pragma protect digest_block
i8/iVOsRIO88HzglcuoKP/btIQg=
//pragma protect end_digest_block
//pragma protect data_block
4Cy2iSXfUxvlDDY3A8RSZHFCk4w3NQlQYIFwy/ae3T6GKrYDcNH8eK/wYQ2suuzG
tR0GBeTfXXfq0lZWHNGktp0YmlzUvSio6QHN4zvADdhPKvto04lWDCD6xK4l1svs
Mulck2UzoVClgTicQ0pQo0IscmvUxOZSCHRlZok4nkaCCwsCFulxHsCboXVXG+/W
ACbc9MxyrjULNfzoLsPUIL8gh80KC+324TkwR4g5yCEpAL05ismhfaqB6rco/AxC
eyO/V9hpqe7l1mJfK4jbxeoSVwoNFJX9AMB3BG7wepCQt410x8RyGLg8RH7TLL3J
qdbzapO9dyoAhCFGNUBDD2xFyLqUk/fTGyBXQBFvkQnHCOIsy0Nev64rMzGmQU+4
c38soGaevx1NJ1kSnkyntJ3AZ/PRCusvvvJu70u15NjxamWxqcRaU5yi2TrXqGwp
svDe/SceM1R5E8CD9Fjn6QJ+2A1Shr7OtDTsQoXjGLGzmtlknSipfn2EIa1pnisR
WLpFyvp3hCQju15ANuoeXe+F9BxuN8LEdm9quwJ0311pGcJ9LEgehWNJs3DnBzsG
0JA/BDz1kliawYYSTG27a8q4GW96td93wuZydyZX6qzsD1AhfrdvaHb0YMgrxrjJ
SUw2W7PveRvqfJtP1xFknjwcSz0kgk+qjaxavCn4DNkCAbAD7iiqJstVA0eyJnoA
uW7+aokd1HJojGzZVUidKQXTmZmYZ400drsdPg9kdLCQj+1why2nRxjIefdYsEPX

//pragma protect end_data_block
//pragma protect digest_block
r7cSNMnacnUYCrZUi32oRuJPdk4=
//pragma protect end_digest_block
//pragma protect end_protected

`endif // GUARD_SVT_AHB_SYSTEM_MONITOR_CALLBACK_SV
