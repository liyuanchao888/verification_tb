
`ifndef GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV
`define GUARD_SVT_AHB_MASTER_PASSIVE_COMMON_SV

/** @cond PRIVATE */
class svt_ahb_master_passive_common#(type MONITOR_MP = virtual svt_ahb_master_if.svt_ahb_monitor_modport,
                                     type DEBUG_MP = virtual svt_ahb_master_if.svt_ahb_debug_modport)
  extends svt_ahb_master_common#(MONITOR_MP, DEBUG_MP);

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************

  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Tracking number for address phase transactions */
  local int addr_phase_xact_num = 0;

  /** Tracking number for data phase transactions */
  local int data_phase_xact_num = 0;

  /** Track the previous HLOCK value */
  local bit last_hlock;
  
  /** To track if the hunalign value is changed in middle of a transfer */
  local bit initial_hunalign_value;
  
  /** This flag is used to disable the EBT due to loss of grant check
   under the genuine conditions of the grant getting changed to 
   other master after the bus samples penultimate beat address. */
  local bit   bypass_ebt_check_flag;
  
  /** This flag is used to indicate that EBT occured during address phase */
  local bit   ebt_address_phase_flag;
  
  /** This flag is used to indicate that EBT occured during data phase */
  local bit   ebt_data_phase_flag;
  
  /** This flag is set once the data for the beat for which the EBT occured
   * is fetched */
  local bit   updated_data_for_ebt;
  
  /** This flag is set when complete transaction method is called for the
   * original transaction for which EBT occured */
  local bit   triggered_complete_transaction_for_ebt_xact;

  /** Track whether write data got sampled for current_data_beat_num */
  local bit is_wdata_sampled[];

  /** This member is used to track if htrans is driven to SEQ for current_data_beat_num. */
  local bit updated_htrans_to_seq[];

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   * 
   * @param monitor transactor instance
   */
  extern function new (svt_ahb_master_configuration cfg, svt_ahb_master_monitor monitor);
`else
  /**
   * CONSTRUCTOR: Create a new passive common instance
   * 
   * @param reporter UVM report object used for messaging
   * 
   * @param cfg Required argument used to set (copy data into) cfg.  NOTE: This
   *            should be updated to be specific to the protocol in question.
   */
  extern function new (svt_ahb_master_configuration cfg, `SVT_XVM(report_object) reporter);
`endif
 
  // ---------------------------------------------------------------------------
  /** Initializes signals to default values */
  extern virtual task initialize_signals();

  // ---------------------------------------------------------------------------
  /** Update flags and drive initial signal values when reset is detected */
  extern virtual task update_on_reset();

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the address phase signals */
  extern virtual task sample_passive();

  /**
   * Creates a new transaction and updates with information from the first cycle of the
   * address phase.
   */
  extern virtual function void start_addr_phase();

  /** Terminates the current address phase in preparation for a new transaction */
  extern virtual function void end_addr_phase();

  /** Moves the current address phase transaction to the data phase. */
  extern virtual function void start_data_phase();

  /**
   * Terminates the current data phase in preparation for a new transaction
   * 
   * This method is a task because is calls complete_transaction() which is a task.  The
   * implementation of complete_transaction() is a task in the svt_ahb_master_common, but
   * it doesn't consume time.
   */
  extern virtual task end_data_phase();

  /** Abort the transaction for which the ERROR response is for. */
  extern virtual task process_error_response();
  
  /** Update the trace arrays for SPLIT response. */
  extern virtual task process_split_response();
  
  /** Update the trace arrays for RETRY response. */
  extern virtual task process_retry_response();
  
  /** Update the trace arrays for EBT conditions due to loss of grant. */
  extern virtual task process_ebt_due_to_loss_of_grant();

  /** 
   * Abort any transaction currently in progress. The argument indicates whether this method 
   * should wait for reset de-assertion or not 
   */
  extern virtual task process_reset(bit wait_for_reset_deassertion = 1);

  /**
   * Utility which can be used to determine if the common file is used in a passive
   * context.
   */
  extern virtual function bit is_passive_mode();

  /** handling of rebuild_tracking_xact on active reset: called from update_on_reset() */
  extern virtual task complete_rebuild_track_xact_on_active_reset();
endclass
/** @endcond */
//----------------------------------------------------------------------------

`protected
KK[N=[bWZS3-f27IZ]2?16fe^UIcd;DF^DU9Y7/)H&VA\0DT@?eF,)GN\4=W]JJU
HYIa:L1d8WMc2>,^L/,+cMX6OddL;]RZ8F?#2[#:[9>gR-Y>dR67BQC?[[aZ&H\F
&,X<LeJ&>C;eb13VRW=c56\8<.F[_>SHK\6?+B+>8273:_MCYJ9#2^&R59b&;])]
g)bY3S9(_38eHNCN^^5EO(LLKEWN<#3L=U_Ve6AXF.[[#:H-^B)PCQ&JcXN3e>eK
^OAN5a#67-2,944)aD0bOBNa2/9FT7@KKQ]TOZ)N@;F\7c#f?M5gHE_2=c^^49#\
[4A4>2c/+Q+X93;f_9E4:E,9QS)[U&X8c>CgWR::eV#@N6?IN-]RL#W/B)V4?VO1
UBF8f(]^()7SXY.dB:YE;&8)7#>f-52&GU^J)N/8YW_?fSP:0ATZ4^LQSR_?2^ID
Q8.D8]\_&)^&UQ5V8C>\1RB2XEA;U?IUfe_PO;[(?Yg+AUgEHGE\bZC7a)W71FKM
FI_ANI0Gf=9P/^de[HIMT=?b?ISOVNf@9$
`endprotected
  

//vcs_lic_vip_protect
  `protected
bN5W]L8_B>T?d16E.38[&;)8XZPN<1:-AWFA0F)cV2H?0e#D?7((/(d#I]/0;PA0
eJ8@<W;S0fQUND(4eKV=A5@I.]c[=KFFPD/Fg8J(\b@+417Ef97Cd?KHYWGEJ;^6
A-NbBc]F&2TD5?g<g(RMQ3LO@TfQ#W]+Ec##Q)9aeM=G?4@H\>c5-#DOOX\=Z>[A
GJ-\(X??L+)K;(1&2KWN@MP8ATV[<KXEecQ=7UG76PNX(5.(@M<acR(31BX[WU/:
=.F\#(Yg5_XEDbHZOP-&9IVTOJ0E8:::4O@.gLg+,1^D/b2/1d3F=_Za()X5K>?F
SECP+H^S98M/::Z;9VW7Rf):G5Q[<O).?7NQAOga3J9_;1WP(/fR=9K<9>+F>=@P
KeHaJ<+G;R0R7D1d;MR/Z/(Y^85KX&<2\LC4:g9[:Ef4M33P46M&6&TV_^H,PL1&
9UIMe8_U)_X\eC7M4X2/RWLGQ_/92W890aC8@:G_A=UdWeH6.c4(3J?c.,T&5g1R
cbHWK8-bZ<ac?[D+,+)0VY;60+F3)aS&)7g?@B.+/LJcWd#ZNW-HNE5OY9V^DT\=
[>EG9b=MWS@<B80C4P/P0M1.QA^DQQ@V+SHaVMZf-d0S7OcaX+H]T,5.#IDW+Z#2
O8=;K#_47eHCWSc(dTFRFIAQS=L<A(6Y(F818B5?CN#>fARXL9@=3DfV?AL&4=K9
41&Q->U;&M.ZA=7G=,<#11(J,&)(DC7a)ZgKIB)>D+)<@#NNKc2?1AO8<\PO/.Q?
Fb^GX=I8JX-=.UHg+(^HV?;O0f0;A]/^\GO@-I<P,:ZZ--_U>-=LJ.Qd1>&VUgDP
1\<YZED;4;N5K5(d#5G5bI^/OB+\2R?c6OWg>D^D&,+f>>.#5M@:Fe-+(#-b\a#g
;=.agL\)6VMaN84#XDbWKBB^/BD+db,a5>@ZJ;Sd9K^XBLf?M64af9.H0b3[)=C5
#6QE_;f,@8.(I.7[B3+Q[?(]1I\C^@/0+HN=D,686D.XU&1BH4aY?:cZ<;OR?@<Z
A6/41]Z\[Zb2d4)4MA-S+65Y[XB5GM:\<&D9UF>DBK(eQ=L(g5\[Ha\UWfQ2c\8f
T[Tb<\BH.bN]a0Cf2gI34KZ@BZ0;;+>>0\7IYNI<e.\0##VRc/0&=3E[72(A5bV1
Z<cfMVRU=9G+bS)0c?bL3g]g\IJ)1LD39/fg(^4CQPFX9B?Uc-4UHOc+7,RZXO4F
aDUH^@.SeX1fFU8:UO2g\05_3ddR3Yfc^gG\1>LGb)g8Cc/FF0FV+5F.3F_A05Re
WVKdB1H>aI9J<@>BG=3:W.FZAcWZ5:d?TY0]6AgBc79c8DV\]CVR/<9OQ)X@6CSK
M3;BK);?OI[Y56341gR4F:e<WfKIc(a4FAJ5\6D/.R^SZBBU<^7,D2(?LTTV&AY/
K>\7J;@/U3\5=YU+J59_XR.H4RE@(VKZ@I0/VL;]0e,Vd2:;a-?DO1-N5/:-B?U6
24VR9Rg0+?9A]4,]YI8IB0+&73UZCJ#INAQCO0cQ@KDRQ)5R;F3g)6aW6b^^/Y4e
+?bYCb_ZE^10#/Q:##__;9S/&f1]8Sa\P,KSQbd=XDXS9RGgARY#63YM2]@6f+OJ
Y/gW&BK./>A_:+b20S6<8MT(c<ZQ@g^V[706_bT)AJJ?GXE0MBA7dMdH/8BNF4BG
/=YgDQJAUa^.Zg62W#Y/9O<F_?1Y:9M0>8A<;B)d/2ZO4=2IQZ?Y_GMALAOaU@#S
ROV@ITNA,:N3//;8<;P,-BCJ@c4d.)RfFUg6b>#LN\a<-]<H:J&Z&G?Mf6HCcIfQ
&A\Q>]Sf>;0VR_XDb#Pd7cEW,;-C<3V_/01-ZT7]/f;P/+<4FOcbW_B:RK)\)M\8
#YX4GI&3Q2J=AdPcE<V(Ec/+D2g&M@/F@4_-JW)ca_N3)bf>^,L:ZTBW-+.B\E>(
-(f_@:bSZXU_KD^(,V[STE+VOWa9QeL&):J.gJ=[WSW;b)?5B0g^0/fC)N3T1K+^
)Q+OP+aIPc=,@<^CHBU-4cQdFZ]H0<BOcRT_.#F6Zf@A4V1Z^K+IT03&U.[DA@^P
gI7T_7/:df,;@B2&V9EQ:-#b&R]:5eLDB+/V/c;)XQBR8F2N1L5<[G49]()ECGE+
F]K#<6PW@EWbF[4&bcG4;;\DI-L+NY_(C0>RYc_@RTO;L,L/^=RSE)ECI:c8FHG,
5]U6GW0ZPDJ=F\f,G7gZ7.>V);G:W48dR=SgOd5/a2U:Dd)C@[W)CT0X#,?b,Q+<
2Pef=^aG;g^V&Og:7IV)I@&#H7INe12BNU)TC_;_RWd3]R[#gMPRDW4:?C3\B)13
a.AB>^0Td/=BP(]gaIR[ID6,eLUJ+#KVdW[02)&AK?dcTYbMd(cJX&D4B0a->aHC
e1UXJ39MJFd&-Dca03IDc#A112SfEGZN;^D/:=SHcG&)HB</XBM/PAg1#JF\M[7H
d,A;eT?DLXKL,#KIN5@HA+#-)B#E85S_becHPbTCQ>6SIL-HTP&C)4MGgRCI/9LM
KR=f=4)R\,X0T<76;2ZF-G4U;44=,2//ccGN>(.b3^0]VeHT0693ZW#NLg3Y7:1^
RS@9HH=\L3C\\=6H+eLSMQ1S(<Jdd2:4gCGT3XdWTa,4P?-.]dV?J<F(2R/W<;.>
3+&UGGEIF,93^ebK)+<-&>);)<ATUPX7^aG6fS1V9=.U>b5@Q-fFO/J9?&6PPC=H
;e;SWV)F1&G&I/_@#IUf(4S=K209=0&@bN,>T-6>SH)D7;JAP<B6A6M^<[gJTWRO
T.9YJ0TK?VPS_C.+FcPO45548gL\@6BQ@]D90g6=K1[P(;@V+#)c30Q+&S5Z381F
(KVE2UKGK02M+39e5]BDgSWX^6I@5XY6XMg>K]6,(_ZM029\b.KBW8D\RE,^P><I
+,9@Q[]eQMA2SVB,a03=#6RYXH(FR:#84U5\LJX&B[TbV,\K>/-MP^>_8D[[4Jc1
Oc;/NOY=J9[8??<&51-N0B9@?\D>ag-[L4dgRO#)JT[^.]IB\N^@:SbW0?[3#3Z-
#SX9Eg+9SG7dO5?_ATL)aUX<>SVX7Q/,bP3WPDKK&D[0-QFCU(d#CFPJ9\ObKF<e
_Q.),)X;@G&S1C\8V]O#Y#04>6U4@<1CTII0-_U?YFEBULG2#JcYUZ6FZK3F;[>;
@&9&O1aG>2;GVc@MKYRUH)[adR@?@C@BTV8D[e:\OQY:Mb-OF-5CYTRa:U,N[+L]
_A.RMSgbA+;DHBc>AENB4T0ea:TB?K]aS@@5DT\(@I>+.HH_Q;\;J#FG]NgYOW^T
HH1aOXS=SKEB-Z]]&ID\(U=/GOCKOT@IJ40MP+V:6BHU8:W7<]SAT=,T1U(IJT>:
.IRC+cH:@eKB)dXQ?V=^gaI;bU;gbOD8J=XaKC&(REe4^N)d?8:=Te[[Z4^+Ec^S
K^f/01?1RJU6B[Lf@A+\@,b>??^Z6/8KKQ;fe8YS.c@Z<CdXYB1\aWNMQOKS:FbD
YZ?=gFO6^9<(=gQ?a\5MTG8+X@fJR,>#E86WN-dAcC.S?/:7^aQ.@W3=&3X;-=B,
-dMB7NH<5HAMW1H8&QE75&5:U_E>]ICW8GR.]8PP\+R^N>7EPLKc;LCY<DJN=7-1
@#4;22)?>T,[YB[?2GK0RG3cI<W8<>&5f)DRB;-DZ@(cXZQ1VZ8AK#_I9V&KJ:ZM
)eaEVYC:)ZQZDB3-5E0M_.B#-]8/T=<NZAQ3=3X2T7LPe;<CEfK_@/S17;Qe\9G#
S_+1^;O8T5/:8G+c,2c6Z-LSQe-W>Q]/5g)Y(SR]1GLM[=(Cf3-J,C]gQ1C<1Q#c
cc2dTfDI]L]Yg3:L7MYaBE<+Y;8Q(ONF]VfQJSD62FWA=B68e^HXK#F8+#SEGdAW
6XaO,LK@4PS6UO^=1\A\O:]>2UW[Le<0/@MM9PR;TK3-&SaQfL]fb)6>eFV93<[Y
--3ZeRVW;&XBeH<BJU>7.>aJI?F;>B;67#6F8gNHTOf@aL)AO0(,cK#O3&#EXbDg
K:\ESU0bK0MN1K^Y<BVG07P4D33?7(9e(eILL<T>)IfPFW;C.NUf:N/efUa(4HFI
X+N[#:QN_7gZfB021RAGVfX&()<C;>>fQI]b>eIPO>1:@N?MdU-),Q[Hf(FZJdUH
4P(E?@WZbD\6]C;gc\Vc4G9QfUI3\;I)7M>9^+=S_K\4W)4dVb>CaIf>Z^5SXO&H
,M8/eM,QS5Igg(?.33:;DR[9SL1+<UaEf<8YMHLeB15ZA+g7U-T7:M9?LBYTW=&J
9@@GU0_&9H+GLI4]3;LT4-cP_FX[BP@(DV8[7[7g]I.R-K\QZ?<cIcM+8BbPRb=E
+g:[>L#))G>U0_bQ<#IFHM0eX<NZ:54S0[e03F(/XH#HLI#+CU<6[.&\#DK0A</\
7AES@IQ4\6KdR(Z=^\@+gdf#:=cW.^2(,9-YAVJdMFNRdHX=BW=LH/[[P7])2E]g
8+7FZ]Jf;5g:#GfCEgOEaBXaBA/KcN-H,VV5I=BQ-1<-TI>/>A@>YPY=FW+29:=:
C-f136/2dT_Y(+21ECY6AB[?+[#c3A,[GNEU<2&\Y-:;KC_SYNXIEc5ZI)&gH,8W
@AgG)PeT7P>>_Cf5YDW-VHAUL]1I,0&Z?<F(WKKW5#9_928FY3TOL,_7?9BX6bJ7
[Rc&W.&L=J8BOKdJ,,bB0TBTZUP#ZKdTQKF2)=,RYSEQFH&c#)M7?+,eIYc#V3X<
440;F:EB85DS1_W3I5TeV(6g56XV6VV(RZ80]g-9]6RQD$
`endprotected
  

`protected
(cfg4RJ8__AFe#FH7[P(Nd(c=O)WU9ASQ16Y>9^12A@XKOcY+?@>2)K-//=T8.:U
L-L7=b^GNS&5D44g+:3\eg[JS(KK47,&KD:>/bFGJCa]B4BgMJ3a4fUF5=F@5MNX
2XVYB.Rd:N<7HbX,,R)N>BVE-.^-COT.J3dEb[.HHJ_4O,a\94e2:YfVEM7/&+(;
B[_R\,)Pc/L@-A[.@APS+\-.J,Y3+TU_@$
`endprotected
    

//vcs_lic_vip_protect
  `protected
=50\F]0BUE7=_2K3D<cacO+&]43Td[Z8g##KYLf]U9O^-C)SCW,7/(:R9LMMKD4O
.0F;V8P)]FU/R72g=a87IS3dR9\X[(2H3eJDB^[_#/DV=c\KE#;#A[35BL=QC@JB
\?3>ST&<7Jf,(51PI[L;XQ+\K;3B1H=04c>0L?<<AL9:Rd,#9P;([f,3b&7#G(1-
9TbY#aOK_5=(RcM@T]aLI)bb-RH7)O^0S:>/_Za1BF[VAL071IQ+K3a#a@RL_cg#
P)UA=^)P-,FF+G>OaX:NHED_0@De?dG(RU:g=N^Z?[?/(?5..U:RK?\[Af8RQ0K7
-(bfc74?YU?)W@T#V91N(]53?g2;WOE.&<>NAP2dE#Fa^g-Z#d/LA(?9>E_cB^AC
A@5,8MKMbZP[N2)c)I/W]5G+R)NF=KZN?X^4,>8-<B<=UEaZ6C:XJZ[#2&ZFYQSg
WV,<J.b]&&V\6d<ED6&\+(T=T48NM56a:eQB]SU=e#EY4#.Qa#SK?)?XdI,&_e1.
U_--\COP?:3\ScZA5SF3JFTUVaHV\B+T>=Yf+7X=,@\JIO5ba>fbYRg;?2623a5<
_fKY/;Q6J<I<.8J&c4O_0W;/JKTQD@3JU64Y.\X>K-ZYR0MVKUX>\)I9ZB=T<_[\
ZM,V7DEFgRJ:(ES9F1);^&W01\]D5W+8EU,H@1B7\;I2J_Q7#6=Bc:UGG&L-T\>Q
KNe1G8FbTTeLde)Fgc)YC6LaMMLBa0PHf)=4#AV4TRc299C\ISJ@OGFT[#Y[@T@c
P8\A82)^0.5/SP\(/2Ld]Ff:^THbJJ6=cC_@cPHbM&BD]>d_b94/]L51M,LN^d_8
W<46);I.E\HVF:P,00BYdJ+,;f;Eg9.Z]R[YdV(?O287V\#_P+?)J(U)),<Xa#I]
a-UVEKWKNP^b/2^]C[NSfM-22]^YF#5HKY;9NF3Cca975J3X?f@IK^511J+<a@TL
9BI4)+6RYfNYc6[?Z_](:-OKdR4]#\-R&BMQ]RW,P-RW1=WBZTWY#8bN6Z?HYB##
,]1W6=&(<,@O<+b.K:Tc4\R<4e=;E>GKGL9AeK8;Xc23cR#X9KP,>V/PY,V&?_gH
g;B\UO,Rac>_aH3Sa4=XBQPdaRNgT=7_JEX.d2+2Rfc-=&N4FQUbXNQ.aJ_7G,<c
&4MY<V^>#g<:?5)(<>Q,Jc&_KScUT)g2X;TIUeK;GFVS<=>(L3?&GB_QYO#g4Z,4
Fga_aLQL(-8,LK-NV&G?4S;9L6I3_Y#N^L(a[eQ.2Q,QEG34Bb\Q^0cW\Z-Rb/5F
?L(cDdSYYD4e3]T@=J-1DRd#GL6K#<JK9ef(:YMAQ7c_,beO^L/?AT0#[G^PcS_+
3E)e@Z79BD.]QVH#;MPT<<NP&WJ6MgV599<@9691\_EQa9PL)UgW4R/Jff?/#6_U
O_U]F[B<Q2d,Q,@M7#cdOD;@eA:JL/XQ]##KILg0_EXGA40/X80,=DP\T@H&R#O/
\@,=M\c<<]J=7<W)9,DK@YZc][84H-BD-PY=&1,b0b?.YfEUcC1<3Z[B_1+RWbYc
-F,^dLBM\a?W,()H>Q3Z.K=L+a2C6GeRU?bL1[2BV2]Eb@#)d4c,fBb@Gg^M7V;(
ca;05DR7g-]#_CX9G3GU-^HITSX5c[b](_6f:a?ZVW-I&?_?e8GgD78I<5bM37Ya
bIQ,Z=,?0J3_=]7IJ6F7dFPaAaT@B)ZPX-3cUXSXSIW9&N?48Q.]?0VS0YQ;c5H2
Z7edP3TS3/\D1\K;OILQ6YAR/fA9YEX76Fb8e6(KLR;O;Q1<YF/0J58\HRZQ=-8>
-RPL)2a@@MR5DBLA0,SH@+ZC00I;BcK-.,4dgK2VB<5T2?YJ1&badJ2BHf1=d1+:
VOE/?G5E/<WWgTM:aW.X:]EQUB:U#?CHQWNUK@9f-GEc)EWO3P=aEZ.9=\^5.OcT
;P5[MZ@;Yf-)GO-5-ZS3XU=e<4L7MS=L-0T>WT[+XM^H_+7Q,0NV#/<)?9W>Y)K9
c_TJ12J[;c3C8;=W7aFf2.fMU]C03)N#1Nf:^Y_eGFX^W7<2-F&ULdR@?#M;<IDZ
9+[gM-G>f-WS;cJ2gGJ-62])+e,IDCUTQ)S.XFLCLb\b)^8H@J=B4H<:)/Kc9N]/
,c9?Cb\V(RC[,D54RCK9DP1/bF4@MbT>G,Bb#(<(4fbd:S3c9=;gQ8^Gf5.K3)9)
9NeE?,DLC)4XLIVG&WH63Vb5.3@?ZDKG59FR#c[=5@_^I:CZaOYfC5K<;>KJc#Ed
f3aX#/-X1:HdU.P=Y6C>KEH31>T81[L=<JO[ZUf@<K3+\0\RFXe9^WZcJ1)b[9=>
]KHS]YS6PdCYLES_TJ.B<Pb]505YKFZ#5705eU#2N-a^B24M<J,0U-g=3,Q,GN[T
S-)-b;=6_\MSH0E\?;M?aIZZ-Nf9-)PeY5.DD^^;0-ZS0RU38,L0>7<\4Jf<7E?,
6B\EBUf3Y@:Y,JB+4\Y_E)<]ga]5BF7f5])B7,&8DODc)Ke2L7;LGDSM4@OEc@IG
6IC3eV#9K.ATUPXGCQ2b[/<+79b\>JP3aRJQC5(3IP37B&C-)>G7>;)+3dd&[JQ[
ODH0QKdf;A0RM\/+YI1dM8WTaI,gV&_HPJJ?X-#)>faB5IC.85(_LJTBG7\W;PVB
.HKASKGQfCQU?D)?5YG<RdS>JO9[UHOMag@V68(:a6>=F6&UBf;N=039DNaACXTI
D<g?9(gSK-L]d4HPQ2gAdH_^N>eC9.I[TN<;Z-YSBf:GY2;DQ2QXLa[SI(fA-13b
_:PIW5aFf<9G@#I7Y5W:@:M9P<^@+U9^ZBKe+NW.13_??I8C^d-6T]08USY,?4Y9
>J5d\cM1XS-H50]cOG;X:2P<MPD&X#B4=<^3Q8=07UO.G>e_QbS^@ADa5bG9A)GU
QbDDI#L8G<H8EfS_K/b#W9IA92MBZ?C/<]d6(.M+CK]bAWDfSd>_>P\WdXUIE7G4
#/SH8:U[Nb>VVg_:6K\?c/+CHNfM3H1A_#eS]CTOA:+c\<#Y:8K)90=/d(D/4.\6
^3]P4Z=K=WBf?ZFaXGGgE[IVJ.a6X3NPgZ7<,>;?BJ(?CXK.F_fHVB5R.1C_)DR]
5Kc93Rc-@eV6O69>3A19Y-a\fY;&4/:7M_^0BMFC,AAG4FO.ZEG2bdARDC_#^DNV
4:<B&DDTa^5\RB+/>]NA6QIEKTC-T80IBe1=;6a&gP-Ff5;O0_E<UgW.\bd_]C:a
S(O9baHUGcg.KO,J_,gIUJ5eU;-0M+V;FT]F[F.SQgZQ77BJXT3Zf0E443B8Z?IU
g@OM7e55+FB[ZP=C2b0([<55F#7Sab?CV:D\85T@\S@=dFJFP:+XDgYZ+JSCGD0+
:.W)0W8+Y-Xe\VKV.>NU(cf3CgE5e^N<f3L)#+C@OLf<CM&a0FZGca>:?G@652HZ
+&#5[e;2.7Y1X@U(_?U=f+,#F[25[,cDJ4Cf#,M,\gS4O4gb(fFNNT_LMZ9O,S<O
>5SOSMYU]U804g>e\,<D\8I78,=-7[5)eZ#MM/;JdQNF^)UX6(cB&I<1\<)g#9L:
9RE?4PX^M_;IfE3?D-(33]8+BS5MQe#2)aPBK.R:c2W@PBSbQKMQVHa[M3<H@@<_
E4&Y#LebMBK0f7OBVN;L_FUZB?\P;2,_BIVZe)V=F06-=S3[F4E7OV/5d-_BV)50
9PYC+&N7R4-B?>82,(&FfN=9W2d#13YR>;ODbNcW_8OEZE>5SGCeEad1c\I2[;EO
Pf_0JCX1ZRYC^M3=d0D.U8T^]0#.7DcPf5CU>-_B&C+HNIc&gW)U7H,Gb@N97XQ>
&Z]T4d<5=g3(C^FU_W_2_753<_8e=8X78XZ^8Q[g_=V44_L1FRbe<462]]bY64(Q
G6XH)1[e7(_ZW@ECHg2RRS]WH)(7b<0(I^T/];KO<WB#7?9BZH=FC+.KRNDV^Pca
f>1.gIcYWcAS-^ZU),WFJYREYYdZD]J4@[B@dX6#R2IYeO+])aeC@MQB&Y;gD-&J
MJ(?RNCc6&=\_LNG=K1Y1O5[#Z\7@Z>?KaPN7?d,(#O^A].PgG(+f)T,?7P@C9c+
3IWJ:^F/RY=(6b]1,55:U.\\MbN3,S[A1=;JCe]&6_@,6=R\/ME7G-7E\@^H3I+P
4ZfbJa<+4LHIERHX86]f^RSG=?5BQ9[#E2M]8-d:0G:YL.-02IB0ZCR?CHG-[P#+
(gC36.fS,C_fO=b8^d_,fcB:LUGQR9VcXL<->ZXeV7>-_:Zd@>UfbN&8\,E[F@GF
S\;CLR(\SGQ/.MYO6D,SScBEH37ae7WT=XIW.OZM4;_NU>Xb.F.ZQf?7;XHM^>E_
_3VeJXLaPeJ0.-/D0+YU<PX(GcaCNI=W1<Qe[2,Pe>/=08D3Wa_D2G=<2D,_>1X1
^6L?a2Be@E76+=@Pd(6O2&C8,+C@;KK0b7YR]LdZ.]6CTLV5THfGQ9gc#YRO<)O.
/TgGRK_eB,;4::,IE.7[fV@cW#.+SbCXKeC6_[P.MacccL&aM2C1=E<](LY@:4.=
AOF=f=S1G>8&3[\GZgZ=4S.>8eM5RO)4K;?#AOGZ^V@/YR1V,1]NZ-H7\G;f89HH
[RXe4;B@?DI;KgM6BPM;7Ffd23KG2:,],9e>KU>2EbD&-<L.HSD7Z]WGW\>9_LfC
N#cg>b^6HO0+&T2aKZUYVR_XaCR(NUe.S47BFd]@L<8LBRU6R@BQ39K[E7S)O]GR
]M:SD)C8dF,#8>:gfIX[KRQ)dV^5D@\9[<-Gb>/)G?^?_)\U(0DF.P?DI(L-FAFU
+3@2;(_?+;L5G+\2:@/e<R30\3a=9-c3HJYD?N_FgXK7D)=36#;QQ\6ISPZ.(NJR
?MIFA4G)U?)DOXJFLU#0;dV)HXR-=VKPBA6<\[ZY_5>AP<+]&Z_I>g;(dgV)Nc]H
#:7SF-P\R5/_?@7>96deJN,b<,3EL?405O/2M.],D=Z/(I7>.PWed;cZ3X&._2HR
Y7.f=fEJ4I95>Q\@G>L#-aUe(.8[F4;U?S/C52(Pg-A<&c(>e;<8T(2A4DDSJ1V:
gd(g89Q^8:;g\e>>8X@CHeW0NM.:>DMR-GSK]gHD?^g0Z6bT18YeHFD+^71O=SMR
QOROIS/]4;;O^/d/9Ff&d<2K]GD_O9[1]-BEOK?G5WU25=^OM<VMfeaL@@W^T_;9
TLXXU;):9f4#R5UE&1W&B\4,+WL/Ig_6F2G2O8/:U/O^OdXHLB6&(R85<RbbVbX1
XecT+IfY><[(QJI=W=g_RD,.U9]VgNI;L;J.WX0PT-T=C5->,GIV65?QZ]K\.D_+
T:]6[0H.]RM@F5XQ2,a-E#f<@bQ3H/[7C.-YW\BP63,Y5<dRaHI^0A5V.dFD@DL3
[G0-5+f;2KB)<L[P,gHM>J]_4_Tb/N._c9(VV4dR79CfRCJK?F1aUF7<SZEW1M&C
cU3IVDMJZ1^OSHYT2c1K2HZLAPGd;VMB89CB#ee-0U(R4-#C&95:(::A#V@HRON.
dSWNQA0e=KKS?^c1NOURDc@=KMB20\ZF6,ZJ1NA70JK,=S,]BDaVHgWF)DJ54/-=
?8N/6][_^#WZ;PW2)ad;5Af#YC.#W5b02KUJJ5P-VYd,+L_)(NIDMgPdO7N#&.-A
4g6ga&f30[95[5T7Za9_]WZ0T@cU/@#<^9R@K_7F>UHHW55=]BQf,K:gM44e38\d
=@ZA6_P<b44267<Y>e]eWgBG^&LU=E/bZ(fS.RW,:b1BIFDYUQ4?NORL9KN(H+&Z
D?c1KWKK,>RLQUf<I:g@aO:(6TD3)J:N)@gLA.,WMTLQIL7@23@,KCW0-F=F09Xb
V,UgCZAcg7YH4SFad@<-A8SVf\JNc/>0(PfD4eIMS5_FaagORKAWNI_=]+SI=X/^
\9A/8V[H72Kaf#0LVATNfV4C\UUJ()C;VRPa)6R<Dd9+DLJ_c;C2?1A3eJ[D<]a5
eP^2#F^7#N/MSa<H;<HN<(gHQ2\Z;9P(<)@Y],4[U/SA_@1g:gJHYJ&5cMGS5>;R
aMQ;XGX\5Zdg1UV10NQ/HFYcaS5V_[Q9JM@e[5,Z_ag4@^+(+K@(Maf8^dZ&H;c;
M7,6];O1VWFG\,.]Y+)cP/Fc0=bdYJ@.L-X9T^88d/fLC;a=EYdNf2,8e,7L,^27
8eB+T^gQaH61@X]bdA=LfPYdGHHR&<Q=K<2CS,D&SQ6^MPB[K45^<0C(9F5_2ZcI
GV-7.3@M<WHDD1Z/+#c1JV);BW@Q/FG0R8@=[CWKOD.Qf[_A@]ZP\B+8:KL\bEUa
&G=a.0R+&CC,SEddQ,XNV^,,Oe&DG4L8EYEAO2]Xa2cLA?DZ[K6-M(a0=T,@4))?
?EBa]9/@&6>T6.MF;B)dMc@W9JM(KDF809I]2XAY59&[I:2;GZHYSQ>.[[W:\EP<
Y;G6F5+2#8A+H&HfRA>)UAA]:0)OA7_3_P#f/DX+I9KL3<D2W0YL;(d]K=&61Y5S
#[0>Zb<8_Sff8^fMAZE5I3S]RBfa_gYT&5GAe=.D_WD(,X)gb#O]H#IZc^MR3_=7
JHEC&S?1/K=b7/RDa/,)cR7BX]f&[O5QW.97QFI^KgRe/>J_LRK0@;=O]3cJ+4J:
\D/F@SgZ&aafQSUV#@S@@Y.F(7+EU^W@_;:7M7/,dXJ6>LU,GHJK))NXeFQNP=I-
0ZV7N7T&)P#LI3Fd,]B__G>I5IH[>_VHY9cGJHS>RbU8N2LA0(a)R#]W.9943K.A
_-a,.JS.#c]5Q_,QC5BQa]NOV5A\ISM?RQ0cYAeM0>/K4c^/>bG+<,JK(WM;0=C#
;g-J92,bWI]Cc;^aB,f,^B(.3]3.?FYM,Q4U0c.B5\>N-HGP<.9+#6cT5Dc^7Zb;
3)XU/9]Q_,WgQD0](N<Q9]#4->NH8PU<Q&3U6<E(6KgE1Q@,:RC8EH.1I;:PBE64
?]J:?a653,;Ng<]IU#e^a01G8gbHfLA>PeNHG4_#)N[Bg^^,@e.cd3JNO&45?CHN
#NQ(3U0/2dJ?35fG35=+H?g-H)#VS[(fcCCE(K@W3,=+EgM,]Jb+__<6bSDMU&8B
c@O?X#B>38b9Z8ASH(CD-a)76UAfdQVR\#bOT)N7SO6C&^C9RF0aUR^_AL>3(S>e
\\YYLF1c4NHILd?;\I5cX^\Y^LHV7OBNEF2MEVM;+<#SeHN#G&D1NOD4.[9XCFR1
5PTD_g(2.=:Gcgf(BV-a[<[QWI:8,20]^OcSIT#MbPVdXUJXVHZ+aLE7E4P0+:-#
?^7TI2SOF>5077;0Pg])(+J8[4M2cC\V@OBaQJ2Ea:A\K#GeU0@^ML\MC7AbfcWK
MIHS3/9/>Dg,[VE;K<W>ZSJS8J2LO/fK>3gBbS.:FG2J?B[8I]4dO+b^QS3XO19A
-7^ETI,(/HHdDU&2eB]<IHF^W4<;ZeIc2_KE<BE@.,^70]QKY4WX5^eJ@-4@SK)\
e#1.9[QO7A=>OL\W0XWF#<M)_1^7#Y#FOH)YX-DQ[eC\&&03aE(OZ^._f,\0QbMf
&dYJXf5N#U][HWS;P889@N1IY&MENWYF;^+XEJKXXb(2DW:NHM.AWN>(Mb;cgW#H
1M/8M^Ld>Rb3]L9E,BeMd()X<d+&NG\]]E2&^&fU?-@#].?HWdL5D93WKUZK_+Jb
eW6CT^(9V/2aeSQ@K81G;MM/ZO1R=B->+[1_12XBU-d[4BU&8,9#5.JaYgH/b7QK
<W>cHB94C_KY7B-=/56bK3>?J;)ZYM,7WV(G=0Mb>G6a/cdR24Ge77#(_FM^:.UY
CbAH.(F)PJQO;;g1g<f)I_fa+Y;X2Jb96U\YV&g,JH[/_\SaNId<;+4BI)abM,^]
b.d6Sdeg74/-0P/430)5@-Qd@dMf1e/;c+9#LJKZg0Be\.T@e\N]8:A/VBGC5WeV
36Y;=\(].02+(8II3?,VD7MeIH8+NMaVB<3.F^LV:d[XF=<,/[#1?77.(.P[&UAV
)]3]Q7QUgJV/(P0[C46W16DWe;QWW:O@M9YW.6Y/[A2H526bD&A:Q3AJ)fZ<3ca_
4CV,AD\+?gHPNWTgN)1L)FN06U46(M:5+[@c23ZgAL.7Q=eb9?_O8<_=^CaG9ME\
MI49?g[&g:1eTEe,=6E[VNC3XfBdeO?bG,7A5O?&BT+..<&_+Q47E3[_?K2UZVQA
c6RDKJ[^13C_K[Y3IJc?BY&YcLH)2OcE9TP2[FYFbHDR&;JFJF+\()6^&--&SO=]
,2N+-8I-PR^3<0N5+d-ba8<4DSS&,#bC14@cfAQ.SgGC0dBP2I2VU=aQW@[4T9&7
&_Ba4b5c\87Z3PS#:6We52Z5FE:<eMQ?+[#C@8<0RD.=)0eUFAec@@^Z)V8b#_D#
FK\g)SXa]SZA[5LT<IA--GW+K[@f8fLFY(E)GC11BfTd^T[HQ;\6CE_=_NRf8M0f
fE_;U)D/URAH6,[7^H2QR)5.&PAAMQc?Zb4#S4[CX([1DO/>N@,Uc(Ee^Q6N&F?a
=Q^1TWdHKI&W1-PU0_BCTAOFK_T,]?01;?W6c0RHPOWf?Y,9APTR-=LJES5#@VTD
KDMIbA[TF-IS5W=B+S@O[HXY;:L7Y-IYaE#Hc[CPY4a7YE<d-,40;-9;Cb6;FeaK
E6T(W+cN=A\:K6BK>EXa.2.CbI\5+Iec@T:>6AQ^ZB2Y.-3EG(RLPO;gaHI,W=;+
TT?gW)<JV+&APbI5UT6CCGI2DSW@^)5ac/S]I4@2e/8L[,9HUWe(L+g,A;MFRK;.
AbRX<NH07bDff6b\5,e_4+#b6^FKCc?c:+^^S)77QRUG6>+fI^X7FLN:>:M-Z[0F
6CI:=Z^N<\&7A5\g/29Lb&0CQ4(B,f\LSV0_bNDC_=53I[ZV=#=M^<1fDISPSgT[
TQ[f5.=b[JW/RRcO^gDN0>13N]L-\W6#c^51_G5.0R,C7&:A3IYQ7N4B/H(NPa(-
V?:(P@Kd#fVMd?Y-TPUf85=1>>UK#^-C,aD=\Bdaa4T1OX&ZB3f[(2K<&[LR+G]A
P(Uf4^<MKY&C6UF62)=3+2C=_#<P5e\^:f.7HDBBcA(&3TYaZ>=&T&<\Kbb&c?ER
85([a&J(MMGg7V>Q0)5\f@QYA.NXT65,A?7O+bM)3VZbZN>[gT]\T&@O\73-Y6#X
[R<&CR43R<-c?U_F:VZe(aAN=I.A<=bFgSN3b7WU1ed^.#38+(42+4YHB56=R1(#
8bTMH5#Y1#+eMCF^-DK+;D83>G6X4QBK@4YgA5G/=@3GLBC[bc?>4JOOGY1aU:ML
_8NP>Je;+W]&@RV1ZCDS&.MO.L3S9e,f[,)A\@cT-F\&=f7b(<\aV@_-;YU[?f[B
;9F@:DKS1@gTB0eDI<1F0VbPA45T^f_)+MZG^7+HS1e9Ga87\R^ae+aY9G+ASfHe
I\g^JPF,7CE@+[XX-Nc>D2,=F3V8,U87aOXA3;f#9#86/;&+b?XMX3@CDK0_b:f>
.?TbSU7H=1=fDT-N;/2b5#<eW?]ee&H.9J\)9f:,8&ee3DT/R>NBM)X9dW;SMB^7
J4J-/\R1_K1-<<<@^1+?g7XBDVPd1aA[eT^g=,;\a78ee5LZU0;dD+AF9,NB_KIR
WD,J9APTX96=<c3RR;B,?58eG=::d04(3.8W1C<#^#QDN\G56@M3>)D/Q2IaV9a[
CSJ-37G&C&?b&,4]2O):bIY1MLb\C0869>LJ^+I4YH?R-/XXG.CNC0)MC[MDEHL?
2aYJ,.5A,6_?+9TJEJYQV=\HSWJeTe.^gN&A[;.&TC/VSTAeD4Sf5U:^ZaY)-S7,
T]^Ue8V]AL=1B4O3Z#V]S85Cbe]?Z:&0Ga9BF0KM]1X<BYbGPVZ=;-fK8?[W-&R;
777a)Ea,N(=Q0.8f#=>O>&DLSa&/6YRDD>),EW2G.;U;56WeO)R#YQ\CDUDW;,HE
T_<)Z[107.Ae4CEMHK:^JEGS@L_b]G]--W?W4(J[^Fd57D:7gQHZdW]_H,a1FgF:
??e4L1b4+HJ<GU6YGD5>WRHVRaF\++:=MKg5OeG]OeXG^Q.<@8J_<>U8d0Sg;+Q#
C-@_^:@QR6YM5\F/>\8/-D)CRMQ)KP36e8NTVg\:#EBDZ.,dF^KLZ(a1ac;g/cE#
-H#)gI8],P?\),-ZCgADJ<C0,1?UI+PWXbFaC@V/,X+3f7L6Zdg3ZT0SO3N9]2,1
&b77SY&TP,V>0[2C>+<66QN;-AHbGF[X1UGUQC]7FS^;YTc^DCXc(@(g7H3f#54;
0Hd4R9.7A_D:;RH\Ed=TTE<:HafH?,d+\:2XHaUGI0Eg/=JT&8>8LABLRQ,5[N;9
WL^DBH0PUgbBaP/9X5e\c.eFPb+0SCR;LAc4K8IYD)OT^3=ZKX_MSEOA=J#(1>K9
&48VD3(#fZW^g6<4d3J+),VE;Q;]0G(T\\H1AI[QH)KNMgQI<7/+N>dO,#2&)R6T
?/Cc1O,b+]-SH-A.W#J,>gG\V:#^9IDBPZB).KBSI=^cF+,ZJA@3_K6B_K.e#\GK
#2&X4>XHJB+^PTY4^9QBOaGIPNNHZ<2I@4#_//f^?cK8Cda?QG57c/aaTN&/-dJC
PY][DQ,UTI=d]QT^dI;F>#^C-B:.#,86SA.;a)fNQgd4&c2_P+9)V>a\WeWR(?UP
eFKZ016&UIAYN>dS>P[LL;aIH)]P\=;MMT0.1B=3]d9[c<FbD-D17,31#\+55<d.
:gNHaY.S.>RV4BZ4-J4bX^Ug,4E:_-F5I<S6RT)/_SSM:G:M7Ib+,=gRX;>0(If=
P+..;4O\D4DWKPB;.Y<3?-H^1#R:d=b#27.-7E5,QW7>0gHW+M9CEQBd-:a<60g6
Md0J1Xe&MA7T[R<f.](XQPD-,]bg&8H-)a,92@:4\1P(>.V_P7f,d4X2)+==]3+R
e3d+LFY5(JI8EfPQ\:J[V#R?;[)Y>/W)9PZU\VL5dHJ1<[Q)9NG>R+MSQDbLW4@=
bXTe8&_?]ad43334A:g22\g>^_?(>,D^2--e2#gUF[-9<H_#9[KTJ:&\79WJ=]L:
4FSPO,DZ/31>KP\AC55c=a<ALF1#=T:OYVR:M4Y2OTG=dG[#DEB9V1H_\?4CG6^,
0@;6_G_V_7A]\.M1ZOD-T,&A9BE;N5a1<g66[.1F1E_-EV,IK/=]8_X]A75(ZUJ#
;-H]5/&3IU>CQN8f&Z,3#K.A+UdfgXH_U7@U3Z8E^S-Q6&YC/](E<T_;55DC=Y86
VSU,,8VC[H9A5OF.>?>:)^+QSGbRPGO.VeU@;cUJ@UI5AKg.Q08F&W(ff+W\@S&(
FKABCPTg<a,;E453+3[1e=DPdZYR+041]J^dHIQg5Gc?W(;^ADY:6LAV(7&MVAT.
-A4N6b=-6[#^8P,=AZ#X9(XOV_?E>85G2YCaHY=a+Rc^6fd+:e@&gCc^P@=99M>c
.4-?C--XZBQb(eO.^QMBY&KN#YSL^Q7GcM.PMY]gNOB5Z&W=4#0S2#X@UW><A)W5
a72XW:5#JEK:+P2+UHDNC;9X,N0K&3(&PbILdc>PX4d<EL=5:a&:31N;<..W=d)g
YTTQA72;6XWf/cCH?(?VQ\Q<.dA6,9QE2<2R@-52>./U@,<[,7@O9L3a:a8NMF7#
JK=Ieb:,/977YMK?-TTfg1\OaJW4T5)88,COT-ZT)=4M,0<MRLL@[C1VJ)L.T45G
1feBA(X.Qf#W=_G<E8FZ+?:;EO3PW<U+V-D>dDNTba(.1B9S]9HgJAbQ8CNRgd\9
(eg)?eFA_R0W24M.<I8G>6(fOC#G=F1F;\/(eV\<6=/YRL<UOP4E\_)SaD_K1/4(
V#QC6XL_45QA.K-#/6OL]0:[818B0PIfAa+/B.16<e?EJedU9aB3CF]V5bY)HJE<
a?7ZD]YECa]JASFI-g.YU^UV(8Uc.7>/VeL^#G3Z9XFFZG/D#\f7AafUf.4V]-,/
#[fJf0P_0C:B/.N+5V+^UI3+HN;.=KN+<0WcXPMBW;?95O;dT)@/Q#:RQ:R9>ec=
BRWB5INa=()7U_IXO/TbH\g/acU>:eRY5e\V.A/VA/K06(f9H0E^JL[Mg+SU)H-X
0P::fPHX9;XW-gbfC_H0PV_Y801Y2W?66^LM/ZAA,dZ-^AL)aM\c#2QIdR[H@[?D
f]_2A+Q.IS/(FZF47Af>[Z+(/efdbK56)^3PO9CE=H7B(GMYc4.T+KO:ggI,P+ae
^@^R,I/7#ga-Vg5[.#HH,d13X<)3R7.@]@N/]c(UC7]C5?;EN0R930);O6=:H)UL
8cH376Bb@.YU-NEOc8Lg&[<B_0I0>;5=P#]XXK[#]O(#Z0gU0=A:IaWI)<4;,\@>
&+YcVC;aJ4LX6;-8Y9b<ZF=7:4HIgL>W^KaM^0XRCXBO??H8dH>VIVN=R62cC&]I
\:)@d2DeA(bP\Z5>V/6LL;;DLL,>/:\DEIID^8+K#A@MAcgeV.0:acb.6#O/bb5O
8[0/Ce>D;VU^XQ9;(Y7HZ-^UOZH?aMO-V;?)#1@0[9Hf547<5K(67W&+^GdgO7&N
b_.<@4(],#=#CUF9IQ1Yc>I7RK,D3]COXRg,8MYA;8;_&N?>+>Jdc@K1<<3FT_NB
XFN2Y[1X]6LT]2,41.b+dNTIMR0ED,+#b:7QNFb-A3/)(57;#7D@P/1/g(ObECc=
C8C(FTJd;;TG#[<Y/&+EK7959;3fP-T((dg5D5AB\1\YC_fFX]J(dV3a[P/AB]N\
a(XaJ[f]gSEV-<@bOcU]=/ETf4V=:IT_>7aZ<T#Fc#Yb(3U&YXA>4d44gSL1Zb8Q
FY)1O9Z8&D[\@ST_AF1_KJC8TE/.>E\S;cG)-_)aZ&&3D=8LKLU+\G>3EY\gXc&F
U77;DAV>8FX=B:T22F=7C,G#PNVfXIEYLfY_b+dI[QT,XeJ)H+g\Mf\_?c.#eM]8
@5TC6HHZEJJ?g^N2bC,NH57=?IM]F//MMC=,gAAAHMf&<P:FW07YV-CRI/512OA0
@>\>Pe>X<>?_-S5c)RD[/W09:71+WL)Ag<F6+P\1Z0a(e&^1T#XBe1fD/cfM:UbJ
-bNJ-OV[/^&-I?:H&dI9C@MH9]BfXEBA&F^A?#AS<85?.:UKZT;-\QXg?I,L@_OF
8Fa5N_(24,cZE<68g@]H^(1NWVQPadUEPMZcOBD6/_7<JR>ZU3AQ8<OYQN\5^PU7
:D>^>0;>7?BNRHR2I-K,\FVPe7:a9HOE0(&UX.ZHZ1J6/<(:Ud@gCKA(A5M1U:MV
6JG1H0He>+U8]1B;\41[UTHH\AU^9Q:+)@<PC1V^+^LOMd._]30MR<E,]UX=C:#)
A):<0SRBLcZEQH-M#97LR>G6cfAf9>[2B1IfS5DER4HK89C/Y^7@d)JA<(f:WeYI
EbU_@6eWR[;TK>4;U?6TZ;=)PAZKM5PIbCC<?<0XSRL,]b64#5^@Xa@7+NQbYS?N
0Bb_gN><@]Jge4))RIX)QL3>4\T59YV;A8UTg7gN^eG5<BUI<299U+.^]dC->d7^
GSb2D@<DJ7.f3fReI5<53@T_KM3\^3Hgf>N4OW\T6)W050ZUQEL[R/P)8F(eb)4:
^Y/O&?e03_^2<5NDcg03/],BXgL3<,<e(?/\K8?QFDI>)E5;ZFX,4fN=KR<GaDTV
WK/R:HA>E5D&0K7IQ3e,N6/bfE_J^I00DHd.Z/L63)P4(AWM^#Z,#S@SULKMG81&
N-]bA@fN4Z8QQJG4]0Gb\X&gI<f:Ca^R:<JW>UKCX0=#1=@8ZVZ+O+F<G[1?FGb-
C5K@[.=8JF[aQ[OGc=8gaGeKCgARFY>B>NdS3f(M+_O?5:CA<Ge<#Z&(5Fc>Q9e=
3I\b&@N1A81DBV6UZD:DBZ=LbB6E=(WR5[.4D1^P?KeP7^,@T/WeA>W>KRT+ORO0
RWVg&V3Ye^NQ].8Q+-/Q>\-TY(0?<e^5FU1TX?DW-.,ZD.ET+P+MfC6fd\J)1GJI
WR4]?#&^,K\/2B=F^:.5Q:B@ecQ;1B_HEK1VRKZ68HU>>f[H+LZ&?5JffDCgT:cX
e;Q9LCb<5e&6T0[]\WMUc_bDS?DPKN]=DHY/cEF@8]UCXZGK;:dTMLMe2_X@8LUJ
)VWBW,_0\[W?L0Ug6>E4O:AV&c9L[[QIS3=M,UC5Z:1C)JF?a)0<7cc/Y&1BQH]3
(71<QMUQJ>[?d&?85220b:>U._5GeV5TK^-P\4YU+aY-=BJNG@>b7g=F=5,#HY(]
MeV[<UVO^JdHS;&fXFe?Ta2,4,,MS?]Wc@3T)@Q;?82(NYabO23cP-8KIY]EQ338
^Pd[7D[F#S7<>>B(E/YC##\]=H)]QNQKIA/FL;A,ES(N(;Zb2B6--:DM.>+/4)[]
/YME)^X1<B35_88>?OQ=0+=H;0]KfgN/Y7afG1TV@@:>ZJ8cJa)G7\J>EA4F&aN=
K,-DRDKf/KQ@.OTXO0#AfdSG,+-IGSQ<+D.42PeGeA<ZI<IZN9)9g2;9FSgZ#H3V
WQK1C_dYgdR^F=_ROX<7EH(<8B3^E7KcF3Ed#?W0BT+G21]Dg0VBCYEaICcXX0O-
M<QGJ\4f[>726(e5C_<GKU=O8_aL/?GbU#;IE\]QDL>LIa:R7T3HVXFPd#;30;9X
3.SgNMZD.]ed<3AbCf7-g&6)FPaIQ5F105\5^Lb]a\=0QPbU\>#&8B7_3B<RLMD&
B9R[:.,9[T(9UD,&7WSOEPA^gWCd9-(;]:D<ZJ,0Ug<g1eA/B7G/]Bge6&6AGFdC
9MH)-O#EMCe42RJJCg&PUKT/];)EdZD^c@/Gb5PUJMUD.+VD0g_16DID^2T<d2<F
;7FFUCH;dY1)4]X&a.]R>a+I^O1B#GG>,S9D<8R10P4\W^?6_^gRHa1^fZ3-9]cY
Q0BAcB<.WC-EFPQL3L[Y.Y]/b]c_LK,#Q&CF>^D@Sc4_U+)aI4:[GOG]O]/AX#e9
0<\5S+N5W4::^LD?8=RIEB?\N:]>3,8<cT&?Q:e&+E8+F1V5H3>(.#A5G(.TW8:b
-(YJJ/=CGM25bH.&OP57R-9WE&K;YDCV+eGF2=@22bN>5gbT=?@M:,X3Lf;W,2CT
78W?77(J^ZP2JI787#GZ>>._U2E6SP=cFR8B1OMLFbCZ4cVI34JW5XA^&@-N_OSc
6D>_6&bJI>@cK94RUe)FHQEF^2(0f9aYBXV[-)W=\=^O?Q.<8B/^4#a<2Q,F-JXE
[YcI>)6ZJ?TZ_e:LV8TRKR8S?#=OLdY2c6GAL/S@<3+@R]]ZR(GF/[2T>L;afEgS
b?<Uc]A>4eQD[E./4GFg,-C6(OgG-Y5+3]HVPFE3ZIa7)2M?GH1R:#I9/L7OC+_e
Na=[I9/#9>R]6L6c<;)eML_YE>(KUTL;<P=L)I#[1,W^+SMUWZWUfL,f1CQ9B#^b
Ged76;gM=e8Y33YW).3=\/Q3<+DET\RbJfV)SU\fb,Ug8=]-_>CB)8aJA:MFST8<
2ZBX@Ug&GI;U3I//+BXF?]=K(RVW6&Ua;H9-W=9dMcVJ_\#Ab0,/Ce,C);^,SbB<
_dWeP19MZDEJME::gG,O>2aKW7@E^=/;;PB5A<Z\J8E(ZC/[]F+7SU.K:+]b@BBG
BN&K0E[@c48@U.d,EL7Y.0DTOBSVKD4f87e/WFGAK#>b>6_US-)X:Q>EQ4CV#-[Q
@)#&Z=X1W1EIaRO5&fQS1A4-eN,1GV+_4XB(af#&d2?XG:HSX0I#G:<c3>N)cL@]
MA57bYM[YeecR;U<4&B(CK3)BBQ<]16W)TT+J7WL,Z&MW(([RaN6,EFE&\+>G(d.
[?fc\W8d#dVIf,Ta#H\YO3F=F3E7])eD:2IKH#g_GF&5VL^2DZ;(eVZ@P27W1c_V
6MW;/,CNABc6#9A/X8AdgbS]X)]1(R_M=(OL\[gR#<dAG6?1HG--W?#&Ng1(fd91
IC14,I]ZMB&(JO/<G,]WF]g0X28Zd2KVU[8@HQJ0D<Ud(72+S;Gg#HMDGKVJ]=bP
&R>[Y:1;JdJ3000M-[=f\^?^4:NNHf=A2MT=#9=TIE<;b6B-A\Vg+4,?9A^/<AL>
G;:[-d>;58E15#EgMZ9b=SCXaVCP,(IU5>H8RHSUV(@b]c[M7dLZCeH/X8+1(39(
>SR..XX_YIYH/e,F7&_:/Db6&e28RX&&3]bG-SGR/+]eTC.+01TOO#.G=@F,4+HY
(S1MJcQ15,Z]e1>3:+Z9_bP&ZI;eRU_1H-857=1<3aR]]aH[@#f:LHOCG7CbL8Y_
_K#PdZXXVXQaR.Nb^c5/:^;7.T\)V2N>2e2?S^QdGT<H8?I=F/PNcVA_\d8M=,;2
a:XIIW#a)ZSQNg1(\EVbMZ&/Y40UD<X3YCC?3^^L&2FQ#+Y?1+Y4B4O[B/NH6F3=
0d-\,2&4NP-\_E80P@@ZG8091N5/6BD-.+O&OM5[^04QW;Q91-dJcL\d@.?]1859
<WZ\Ug5->UIK1/=/ca\-eaW<Ab;F0S:?J:]\-R=M7ecZBXEZW>FO_9=g-RRUXKa/
SdTSZ7[4.=9#d78IQ(R.Ob9>_ASAFKO@#911RLO(O]H-V3):1>e>[8ZO&.Cc8gHg
H?S0CQ[J7^2.Q4gU/R=a]U3;+3N_Y:/K7\.C&DJB8/AZ1JDMBMKFI9@eGVA9NW:d
6>^^7PQdL^13U<9AHa3_P;RPT437+(SG[KQ3YU,(d_;aAdLP:^Z#DBeNP5A5WYOS
UVJg.:9I-FggXe;&29\ObSPY5(Z8.#0CR+H:.eW7CRee/#-BKVQMfBYO-T>PJ)0X
HS+dVS2B4/2@]EY2ATC+#K[OY:7)eWa5/Q_NP^.RX15Q2E?S0V].Yg]1He9K?@G:
1;WF8;L.BM1:#3Y]_,Kb<.0J&&SdV#bA_-BV0^cKU<PgZQN&=DMD4;I&;ZWGC-[P
7,g)L-Qc]>TdIY_^8/6XYTHXEH_76)4OZfA)NbB5fL-1>E,/C9g#O7(AcSBfY>>F
MY8d&L5JS[2&LX-58E0(C20IcR#/7;)S:RXeZU\\0(P[@?U2MES;5QBf94DXS(Q]
BD8BG9PN(\XP7>I(CBe\gPK=+]gSfL/a@3\DK<R/QG1d7@7A<B<^OUIa]d<A,,F1
E]A#&3a2D#Ifd5f&f=32g<H_+[6.IdV<(?cd^.=7XcC6O/>8B_.:)A.TB2N4JQUe
&L-4f,>Mg;.OEI3;>N>4(Z+=1HFSTYQPGP3BC?F^K[[7g>6R]X-P^;8b_11Bac#>
DPZR,g^,J1[)Q<?SUO#W9OU^C(EIQNc/Z0?N&:@<6[];G[Sb:N/6DC9W@#9,e\Hf
c8gPW_HL]ZQcKD)S\\6-.Y9aIHDbZ[3QaMf?Me6.^fY8dG3=4[M@OR?+8\V0A#9L
8FOYfP9J)[T=2g:d^,5HO[E\_:e:LX8P>>P9:&bO/]0e?/O^X<)-@[QGC>DCe6_F
+<4T.[&Rf\0fU&4LT7[NcPbFCGO9MPQOG;\V6?c05JT&K)@E>dM-G-a?7.F+OG@U
3?O\H,WcQQKGSK=.(^[a?&?TG:;8Fd2(,[XTHec4a6/gfR(R5:dC89_Lff84DH8-
[><?]V74)+INV45=d2<I-XU^QD;\d8-HG@>eC=,AP,:aBT-@<d22/c?==8S?6>c)
QdM5E>S>^N0WPTQNB+gH:TQgZ?N:QPV)=\-e3;>Ia4BI7gI><A7.)@41ZMM+,DZ9
g2;_4U+.d=H#O=G+d]SJH1W;D>KI[N-[7NF:IJS-6Tg-cDM=\&PV>F_J9(OM7S;S
)3R.Y:C:acPAHb<IM?MCK0gJ#Y0Hge:7K0ea(83:B9\FKYT9:b(Q=aZX?H;@]/.L
J>^#^\e3^M,077ZP.>E.I.O6661(YT@:>>P&Za1aJSFM.f1@gL(O4_]\]a:NO0FJ
Q?LG6BH6E]+0O>LcH@:afOVJTZRIbC^S;9I#HX7)=?)A^b-51GN8>./=40+Pc.,+
d4g5^CcSQ2-=GF+Y?Z93^;X^,U0H>XLS)c,&]_NCBG9HTg4DSG=292#fEdVbVbMe
Hb@G1X8W,YIg_4GIZH/S&bD^2-fD2_DZLa#J2dB1S#BJ8<Ig+E@?)bQ7SOV2/HN5
QG?V6L#Y3+_L=TGJLe]ZK6NY35N,=.aG(f2#&0F:c5=gQ[H1L_:;7QX;gg8()-H+
4W=33X]bA[K9LECVV._]QPU=?=C78A.Jd+:fHWB,=Q\T1>I/+0AZ?Z^6Z1TKJ0P@
KEgcY2KQ_^&d6+0(-N2[>]L/\)b/AdM68gK/X7HI]d:_a2W+\fZ#U/LHUJMW)@[3
C<FAKE=b34U>]/@.>,(f\OaFLKV=_3K#47CfXS8,[8W/7RO6Vg/)--W(<IH2I#3:
;cXF:U;69D)fdI+.UJ3g2C+</#(\OSKP=V>Z9QHZ98AYBA-.N+PBO\A,e4^+B(ac
OH,MT6,:?V9H6L)VL/;?.)):]NU_0deL3eF.G9B0:Fae?cDH?N5f&O6E0[VIWIAa
;eK@_Vg^?]Ze32fUPN)ceLe6=/;7CW1M4<)E?:KJ(-@dI8:AZMKCb78e;.SNd=CC
<0687JW]T]P?42>Wf6^3.X/GAA-(4d3N?W]QIH)=I?G2Z9C;<-H+U]d+GfR6W3\W
56LQd9NaFIKE(W:/RNcQ,T4ZBb0Y<2P_-/FbRY6@454:fde0(,DB9\7=EWd)9bQ.
BNdR0UL;Ua9RY[:D/43:1>6LW9#QbN5=]=6;XTa;M,S.@.NL#>,=IWWUFG3X9+Sa
P;C&9aQ3\\UgA3U(5;aaV&D3@#.4Ccc[=6(;5L:(SC+Oa))f7T4IC[<W]cbfT8Rf
;?#gg8&7[fAd-IA=b\YH,@_JFL\,@\?F@Z4K,Z(dDa?E1ddJ0PUCM[K;4IAHP2^(
BIAdP@d0,HP8ND9GgNG46.O0I)XPW#H-J_FP6LE@N)S#+Xg,1GV-NeVA^PV6[M([
/=d+ZDB:PK?e+\8]b1#XS>C#dJ3D():D@ST;85#dV4+.c_J>]0,>K1<45.^e:W4>
]P\0=KVGdH]a1,O#6AM2;_)(GY]RdDJVgZRa11U1gLCV:a[RLIRgT-:-EN@R@SS]
J3UY7IRWD-5Z&?;@C_7>D[LO_N6gS8EA3YG2#8I@]YAX_U\YY6[DNH^.eQ9dK()U
7EWRO[1Z#]0;^,=:D0CM][8?)g4=Z_;YOEd<d44LQ&]Z4\cF<.I_S_IDeb<<J[6F
K&)Ka0b#^W?\8Jb=eKf?O,WaRICKYV0(5;6_\^/Vb->=;O8+U1HeK,3f?R2_^dgV
EaU@@KIDd]&,.ZQf8JJ7X59[Vd1B1SWcf#1QU3-88B[(\A^CY)aNG0L8N<IBSG(d
,WFF2/L=@V5g/gC&Q?F5QM-5MQT27/R]:OdUa-6SbeAaS_f5B[_2J@8K6CGO?KAR
;\(Re[7+eZ:KA;.aH5P8\fI8Vc,C)5H3=Y@HJ,@CS7E)0/S[a)H)PHb&X/\Tcc=W
^#HPMcRVL>B5.d7?/Q:;3#>WWd;GCGTF+=4ZcBfXe=](1#5K[=;BH<4X5EVJ<XL=
_AKaW(>#>XMgcD/C&:Q)6cd;];K=.D_L0(-Z/6XOb4AFKNU+Sd^/4QF/S1;@9_;B
4Q9TO38]C0=RHeI)#H8LXHQ^-?8Z&VQ&\64=6WF&ba2]PFVg^BR=((KN2CN4gO_&
eOP7M2N9A5G,@0@B?E2dd5T+1\2\D/NQGZUCD9U3TN2X2:A8[K1=]Ug:&.S^>U9)
TEEdHdN2c>CB_9@/1U2R8S[Rc^b?L7AI#&<Z(\Q&@UL:RPd?WaA294#PfcH(.e4-
/abLJc@#684U]>:eE215PDdOJ(AMRdeQK8@MS])\BCUbPfd8b8UU/FM[-aY91_cL
3D,47M)9]/E7OXI;EdM9]Za.@KD98CB5Y./L[]]+[EJ<\CM<?fL&=D=HV+46Lc8.
EIdYE>LHge7WdW[1#CIV((8X&+TI/K)eFRGHZDE\2A).Z^&?,2:<b[LJ>N/<gWF^
,12GQede4K&MV.S,5Y6<\Z1V[MR+_HSZ[F93X4eLO1)W<_Qf]Ca;N#U/?IQS)Z;^
]B17Ka@KLYX+d85KgM(PMG>AM0gB;&0e9GRL/g99IbK)HK(I;&?<XSd09890.e6/
YRSE^^,RSI(9=)L_7&@X0TK;b/BL3(^=eX3@F^ef(EN8JZV(Q2H/A>K0X7bCZ\;4
FNF&XfH,eI\W/Had:[c=7HU.Ag)7FM1HTfR0<(1QCa\E^IS1,[2Adc9B/I:9c9b-
E@AL#WAX\1&PF4TNaW?/DHbC8eA;UL=E/RICJMc8)Sc(L(/ABKfLc\5DJ3=3HEbD
\W+&cff4^_EF.=]HcYbLXG/KC,DIe7>SKYFS)#BL=P,56gQ9;A#g>X0GY;eB?K8V
fD&\L5RO3AEX@0ZDXHD#P4:RJY3MO<?^6//H:MXJ:2:AOFTCDJGD^,W>OW^5YPYH
:O#^RC>GORVN(Z-0Ec5)ZTW9R<,.Y0FJ[/ET-S5MW/W0IUWZP0(<DF#6I^COdO)7
LYGB&UE(<;TP@FBTg=(H#AJS4^5G,L,/;^d,cS/;S<+X/F79/L)(056^(fP5EOB\
1Z.Wf1=;=8,5[GD;=fdD=^:-UZ)f^IPaW3F-CCXa8RMA3)S<c+W:+)JS@RYWIf&Z
3@?a0S?LF#.6+PP&8L7DACeL@Dd^BL?;JeO5/3+Ygc==V5Y;dbFAW/8_KVg?]UJ/
OaA^AZ,d+:[\Y2R]P?<b_9GIBg>TA:)6P268/^V3#_?g.&L5TT24GUBeILA8Ua9R
Zc:OM+>GNgC.VV9NN.Yd9]VG^cELM<,:_D8YX4Z@T3K[[aH?f43e?1V;b<J)bT37
CFDM;3VWRF5U@B^3XHg#V1T?GZb0:B_J,6g[4fV]4M-BVTDA.D1#T^ddD^)KHB#\
YREO_D<CNL0>KTJ3b/@K;F)3=J.f^]gORH]/1/VA62I)@@@^DA?11bQVKR\KX4O:
4)@AbDgeV\G41@9F@eIAb0UXG,RfNCQ<;+g#Y579Ta73E8V#,OeDc<5,B#\1^19G
,P?I?7LCg]+.@3eSUY=CN;SEZVb._I&]WR7_H]&8a#(:,/(^14=Q5O,+<PU&&&bJ
/OR]Wb0XR5CFdRg0JSA,=[WCH;0WI=#1T\J^BP>>/>,;;ANJ,/dV]Y&cge\Oa&fT
;D;@3GfNJ4fMXB.-4S4GQ#+=ESGa975bOEPO\?;;1-@0=Z/F5,/OX^\M2SXdK>Dg
CU+bB\:@HD/(bLPR)8Y]/4,Bf1W/<M8:L&gAG&dC;2c?bcBe0Q_2XCYR6YG&278Z
.QS(1D8>>F=G71J>Qc+ZF0N,F+C91T<0cAO3O)d#MggO>H-PA:dRSWL;FDXHH?-b
I#aOD543;/b5::9+4<Z\:9E9ORS[WYfWEEBc4UDdeFJI3,62/(X_@QR53KLPOF[W
]<L2ZBb6N13,=7__\OTd5Q<TbF70Yg4E;a5>7[T<.I=7c&ASP(P;63OI.0K(f&fV
.N:]L5#a\U;c/aG=YUgI>G)^90(;.WS1>GWb#Z>OVS)GfaP=S/Gd.gCI&19d7,#H
</]MM-bOb[d.?-P.#>XR7e/Vf2F/Q@=;BJ@O&Dd.\a73Z179A)NV2S8MM#N@(5CG
+H]Vc&@LB]R?P,cNfU&?3<L=?f4.[I=,W&aL,PA;VZfEPb^E#I>SGJBU58I6OXAG
]F:EH1MMSdN)Hb(:?;@XFI#<1A,5_GfGg=^IY_IcKE+g@(=GaXXa[BUKKT.K_+V4
&GUW5ZN4HF#&e,Ff3\]V)HMcS?GR5d]]K)+]LTO6@>TS<e4-UMUESDPH^K_B:;[]
@CB_:+C&77)bUY>)FA8c<H+>[>&3N/]-Q54Pa\N]X,XBV\e6+)a2WB7c,F(]KO-E
6eY7ZWKRT3bfP^8(c&P62_?1WJV+36c/&f;#,-Q38#->S22W9DDTFEWa^W1WN]0&
Y5K1(4@4AM7/8gWQ71R]d^\C=&W6](H([;]LF,^c?A?FDI2+]5[2L)P/M<UNTCQd
_P+@ePd?\5:GYLZ;N[80__9_JHSJd^+@9ZF,HRJ/b4GSU[CgOCESJ0Z7^Vd13XHK
&8FSN,4,M^L?QA<:@#47Y0V_d<Re2Y628bIV9IF?F4CYHUJ/,R(.A^/b]5@Q1aCg
61&Ua-_QI,V.7?8ZPd37SIQ/IC>HKLU^O8gT31WUXFD6O<(A+LVJ1aM;[e-1FZI[
c/;E/g,=dC0WKM+DA-9b=OX3DfdP)0H&@@JcH]65[Xe8CTgXO6[./B+faBN8R#KV
OLZW^W;CdO>eYJT_bV#X6H:@+3Hd1d_g&]JH]8Ng8B\_3Q_(4fV)0BA:&B&(,OL6
<DVNNOP)@-HL(@5II:Q5L\5f(X#]\MXN5AEge,&Q=^=<[JD?C,)P6F0N42_]HM<9
VB32/Ua[,g++6-00R&/fNRQe7@M[Ad^#e&@X?W>F[)Z;7R39O6@1eVW[EZH8C_[(
3XM/M_fD][Z)L1][e/Tcg]gQZgS-09<Z,:g7/6_BERPVd,?edI[a/0>0fT&8H^Mg
]Y57EfX9:eA,X@.Y61OFJ4.aNQD11-e9OAWaL\>;W-YF5K-Z>Hc?=f#8Vf[YV)6I
W=QFTWb9_6+I?HJ:L2@W]f)Gb.QK>.YX(YE^W_EG^=:fP6)/O6C;PVI;@W\.+8^L
;d?c[W+AfBZ0_@)?C3f167W<;9fX1RX9X?gJQDIb=;(Q\#^&ZFH.e(1/T0d2O:GR
988-&-Hc-F;4;bEZHgfQD2S[ZNf#6#D0>[4K<035GULc:J,C[Z6&O\<)8;Z=E_I1
+3:[54T):2/-U77-((8Q8(66f=L2f9^K.,X??[[<#SM)d,0c8bI\:ZWD>Z._X,G>
E:R+fRVC[:BfNfY0G.FGZ:IW];]WfPW9H0C=AUI@F8J16>3&9U_RJ+/eSY_-,X<#
2cMLH&QY]][\9J3LR&XOJKI-_Ae[=4/.bd3(e1<4A<\b3?Q5/b[gPW<KJXU&Pd&)
9#BgLT&ccIT61VOVO>8aLfg2A0Q67fgUM./H?&,7fY+DYO9=HA)6,\Q0MR1NQTBB
7QQf55W9\:UAbBK^.=(N>+3/YGT04-A8@=5M#A=)ANV;b+G/616[67P.UJ,^Q,=?
edIXJeK?OLKJ8Ue;?ggZ-G<c)c@VAT-N5]LX\Q9JO6dD&&XfVPWc-DcZB^4d1PYS
4L,fRY@TKfC.QVJN\LRG>8U)R)EM,HXSR7D[dF;0##dAY2a0->2NZc\(/F1gbb@>
[0)7:/6Tb<OB^XAV&HD\AF6QOV-d^;8dQ#B1S)T4)_?243]&@/;J:NJS+S1PW?\6
eR]K(1NS<6Q)4BHd5B5)SfUXECc-TPDKF>P.e8,V87&^C<K(b18]R_M\gA;?BN^K
W_RX@>eN9M)9K6GV<40DM+Q&Kb]HV8e<dOZg3I3=0TaN1O24FW>d0@[_J[+>+^Y(
U81)&)]Hb.Feea&^dTbXFbg&dQ;NM_UXK>]TTM0HJ+c@+@BGJ5YdPDY946,ge)D@
aI2R;V4e^AZNG#V27/8@Z#,21@F/^[.=;fH[SFK5CE0SFXH<\Z7N=?bFJ7N;,Q1g
^@XJTI<JQ?.E7e_8-P;JZ7Y+[c:TMScI7P+PL3R-V^,O0.fNLA>TLd06DZ;?#CYU
+]:J]?:7cgMIcV^H@&eIJ<C[?#-_-I<PScc9@8<HU:28<b]-KN^\FO>8ZK=VB>)^
;4f7gdF/gNAHL2XH>&TXG;Q^-U-C)XZg9/P.=V8]^&[\=A4Y>b5P61Ie3DUXYOI\
CD36ZcaPbS4#g.#((P/R?4;>/CV#:b^BgI=1f<WSc(=0NC-e5bIU>UYWP,Nf_>?,
3C7G=)I_/(G6AJ9H#A9XaV=CRE60YBT[d5?):fI2ePM[1dJN+0GSEMFc/VZ+3@P&
K#Ef\&J(YK.AS>6I?6:_CHYF,c]E.G\Sd:.E;gd2-?-Q9^-DX1IU/W?ETJAfL7a6
0WJe_Ie=]SV58O4>NN>Q-G/&DgT3K^C+MfW?)NHGGY3JN]P=&gK[[cM4L(L\:KX.
J@;(8dMW_fG=4Q21e=UT;8;Qf19UVFITb=/7A65fGUM5>6WHKJPY6-A^T1PSVaY6
4[S3CU)c4E1GI7AAe_GAbSIGQf_UCC+57)c]1fW=;aB-7F8:<Sf^;;fBGeUbe._f
V+.);BY3FLBP&,59LQ,C3d>8/7OY[YY453J;f-._AT-SFM=SE5#?98CGQ+Egba/R
(MKFX3S(b\9U.dV8,9g(B.C_DY7?T2W#E]daf>VP_ebON\4Zd&B?H-R]_CM>a:5e
>Ke?2,]#:9/SO.e<eME;NL.27e04OJK((3F.?V/Y1\\Gf<S_HW;C^)QH?R.#96Nb
_MgR2g1U:WOHBYCP4&:M7[.+9>8ZZ4Y++5gSY?e,QY53#68<83U=VDDPXUGU?#I&
dc6\MTaL=;@\OSU:1f9<da2/272Y1D>H=HA_N)>TaP?=YPR9,F;W2]\Qg0BBJ_D.
K[.G@0O9gDZ4AY,=MP-]QW\CF+>ENNTaIAg_LKHQ7bd>W_dB?]4[5Cd5@7G-A;]\
fD99dAQf164J^6J/8<UV8aNB#-Y-:5U6&BH2ba+dBN.g3EXaXJW)LJH@Pa;MMa8_
A-SY>a9N(-F^fUV:=(?eQ@2T1Y^fPV]T2N/DA@/4WPS-@/TZ=,N?DA5UfLLLR?G>
HbLYF0=]4Y1^D@-/I/@(>2LgV1bZL_Q8>dJ,?6G<=CgBg4:LCBI:9/G#FYTNQc):
O01S[)#PENB<C4/3NBJWP]dBN+>EZb9N+F0-a]NeU>=BYA)[?_R?[\6bYa,IR:2P
b^GD)@?^_Q4;0^.#0:+RJX+.UWePaAc?K0>]cR(T3_f8+,Z^dUK@/R)17gc5]],7
>/cZVNd5Fe2\&fLd@_07dK-a^[KW19VS-G\S,-gZUEWYS@W?<2OLcG.02-Sg-01D
?BK)gI\2YEGGOVVBZa:C&@A=99GgNFHF23?HeD22VF3)dVJLM+90ZNcdN61EZHXH
T;@bK-dW3c=b;OU?7-U7A^U6bYS@Q6@=99W@/;L2D2PCN+K74<MB1B05bE8;G^6>
C7[JIe9^Y-7R)Z7Q:^HX[53/GF>^SC0MH\Z28?_#fO4bfJ-CDMV)U5L,&gbL/TS-
9Q\5f)6:<U)2FYb.+-U+dc32SC3A#cB_;MI_86:K0-SU/EO7TX7<58f==(>&QR/g
=I1AD9+YN[=2,+(?Mb7W8KF_gP\F5LHX9B0+A5E8ERaALROX>L2WW3,\A_XOF.R<
L_GfM4;X2D<.Y_;KC)YMM<eE:],TeY<6NL^PR6\6CI-WDR/QNL,(\JcUL5(/(ZS(
eCB;NX0JB:_]RPUUJ9AX?5B#Q5fJ>ACX^O^?O(G>g-+&:@[_3CaCg)TV,F;U+2KV
11/V=,g(\+Y[;I63_RWAMc_LLJ^8#,\d7g_P5>?@GUPV9\]ED0A#[C^YLS10gUdg
/XK0&e4N&(@JC)M=RI#9=(D3QMR#1(&]3?<26LH>(\bEA)2EW^N&SbA(,Tg9AKDV
W8E,.;UI+;R?ME>d0S_N\e>5;D#3d3:Ta#>U(<[Qg8JP[;T<^Y3bSOV6)KdEHE.7
E0KPf?D^:5Yf<E,YJ1c84@SF_<&T\Aga)C.bC6^B5H1[.E1Ib/XT6e8dOfYbZgMK
+A93eg;+OU8WKAZ8.=5PRVW2UP7/QNbdfBGWHG/BH5b[J_=I#M2J31A[B2[+L#[)
b4/428SLAR.:Hcd>IV(?CH<1D9;ae<c<-gNH+ESg.AVW+[V<=\g5>)XIEgMV)B53
Ja\eY2-bJ?IT9>3.4<^-]L=6RCPQR7AdT6\0TGgI2H9,)C(\c\KZS,H]^[VB8I:d
#84C<a3B4_J3?GAB(@2IJ0Z;[E:D6HE8,HF)bUJ0^8E5ZT-+B1+\?Y(Pb3TTFIf+
cGYJ/)<UcFIDNIeO4OM<:(AUJB0I4T&c#g^+8G<T1a;d><T<WG;),#?(.e=dMGg8
4AD;A<CUD(?0bNO(eE.T?O@LP,@8,-42O3V<^L-5RaUf^X0)>f2e9,L^3cfCaDKE
?ZX-KT3&\\?aeJ[5>.[3V_TN6^6a4g_+9>?G70b-RR?2(8YN-FY<>Z7.^]4V7KZ[
e&4Y-;]Dce\4Sc)cBW.RZ=:HI3.J3+-M?)gQMe+NONc]/T@.WYPa5+B5I)3&1R+\
L9S/bP-:9a6fb<?G;C?-)J&L\T)::#P;W9K..:XV_B.SZI;#+eE6JT@D75AbcAFT
6EBSPQB37T=?N)/#?Z0T4@g#b<B]VN(YFXd;^KANb1e5H&0WRY#3^]ZGWZFN&,;,
C?aWJ2M9Q(8dI:^?YJeE<KC<gQ+Q85LG);K_C--3G2b+21J-C>]IMVd=Z:=;]MZ.
@S2K[(U.8\K(JA;XI(2_Mb>A(;=Q<I;7@/1e6M^0?QD&+)[#ePVeBZ^<C>(7]F_/
?_T6ca(&2RG[AMHb&4F\GH4aO=[bNJ08X0Z9N-2/PXgQ6<IB@]dM?P+;JL,2dO\#
X49CH6O/:&.dC3YS>WBYAV>8)Rgd-@@a:P9ZZbBT5(C86aDV]HUdT:N#c1P/.YXg
<.[_/Xbf,;TP3f);5+,--?[&Q8LLfPecBf+4^g=#H_FJ;0A016eAYSe:RaaE(S7F
SR14:AMWY?GeWa3TUXBI62-3cTe4V?4FCFRQ@N0C^f#_TLXB<Q[2M\>1Ia6VCd>/
\G58:ZRJ]_gMS]0A_[<[Be]4RW7?+Y6&)]7H[O4TPKY#+<<?aLEFfA6P87\EDXZB
TS]a9F2]+dOM]7&,b/[9RLQ;/Y(>G-R;g=/XaLX:V;=KV2@g4UN.V<SI4#9G=;ZN
0,I/[TEGcDdg.<JB/9,fgZ[0/[CF38Yb=CS6E@)70=J?^6?<NTYOd2X(S3-A0G^e
ae]T/VFBVg;9J8N2:O8>6Mb+WH_M&UU.+aeIP@+E--,2R=B4YI\X33aWegEB[3I5
L8)A]6LKe?b0=1)6X7PH8Va121QGHQKD<O)BICf&NEVD0MCQRH[ZQBMFE4/GD=c1
?Zg(>ODTP9U0bc_W4c5)IHLcG-I2Wd^FJ+,/R/2g)G/_FOc=-R,&[]@]5\M0T<+&
a/8X[8Oe,5<]>W-_dFEb)]:0/R]DdB[H[X5cXV8D2ffc+>QO-SVIJ-ZEM4HK[T<g
S#BE>B6c2#S]d5X^S30N@d6I=8UB>&<A[a0Z+S(3<-#A9c6)_V:<V\PR&cGeF\cL
gOB>ed@0WSQ3-<<LAZV&<Cg9#0JQ\8R)79A0MfN&6_PaX)gB=+U1>;=O)7ZZW,e@
c>AQ+XdW(-.f>497a8L++QYM>dSf6IbUZ)TROb:Q;HYf5c?SgWFS#>&L@8I#1V0d
Z2=WeB_6<e6@-NSQ_(X+9L(KL]&[1T&]3X-db1PF.QUM7^1:GGEUK:>G)&G_&CIM
KJAdH<>)g.QVK4Cf+@O)7J)5=PZKe9b)EP2OD.#^DXfZ5eZ)>gA,EZZ_M1g7+PaS
M(GY[369]XD:#LJR9ABa<KW_/SSB<fKEf4;0(S;dR9Y4d]09,C:9]3R&&c7cMXO?
MD[A]+V>e#<,b/<7YW[3[UZLOS&)WaW8C_10&#HR3ZY<YMY;D9;JEMXJa0:1WP0?
NBbUAAIBgW?HaP4(P4c:-J)2G^G+XK+WE3IP;N)O9Bf4R,-S-42Q3ceb<V57]\]P
Sb?DF^H6>M38^R+R5[<d/<:,4/(5SQID9_BNc)&.52NKbCJVd)=@eRJ6+#a;,M5?
\<CP8-2()<g.\2->BQ5ZEfL4W=.8717)//,U-U;8?d<3.->F5)_<,QfgKKHEW8=6
2SH^dUc=SeZ@R)^P-(2;IR+6X;SS:Na>b_:M02_1cF.VD?[Gcb6(I/S).J\D#Fd0
:c<,eKV.5;T:JG>(8O;3YHS,)_HJ[KZCP,I(43JQ.QXBUZ6\OIPNR/C@8UBeAT5U
<OEVP78C/[Pe[_R;VGM5@eb;V@G[BHYHE25)&R5I@.OG>[U\R5P6=a=5aX+RO5V5
fK5YC]d,&OD0YO8>)CDc(M\eO&TR+H11bPN3RX,R@4X6S70KY]=Z+WXR5)9NWIZE
_8VQ<JMT+FUI\EN^HF(<_)YVfQCBWI&@DV^1Q/AO8Cc:@4d_ZN\8:FVORfd,#;gW
-#-2QB,-:&=YJ[\CI,8J(]UGTa<V+C>N#-@E&--LV,Z9BV?@^#T&#g2=MCg(K=&A
bVE=d?bd/ZAYUF<TS-J08H=N1NbdO/?bg?4fO/3[I#X&8?GIOE,3:b@H3d/>/SgW
A]a\6_SN(\>9YUa5[a<8WW]R61EGBPHT->[FXM5OJg)XOXff6BEQYAA4Z,<C&:Ha
d<G-g2^T41d#TC0F/>\#gL0KFb>?7D3?=+.=gf/5R@EW/7YGZNedbC)@bg?#77N2
;P1X0^VF?PY_=EE=4MZ[BMBG)B?94ad[#cdL;a&S<)(D(78D^G/Ac0L?6[:>TQ6+
:1P_b^8VYJN.7\JfR:+DN(eP#S+>bFcg#EaafB4McE_BAfKH^S]H[0.#fA84RU]Y
SeTe;:WOV1^,^4XA6V28;)K&g-6ORH#=eLFU/b-Y6HC(8Z_WMII.WY26Y+]@VEfg
5;KVc1aK,T#bHg),OUUB7F.4@Y@UdGbcN]bUT/LW1+ERGeH@Og?L[Ve&GWG[:COR
GOAdW-I6CUGe+T9@B\QdOe=K;OTSdOUBd=bZ5Y^Wa18N_;]RS2BfI(S2>Z#,BaE.
RU8NEd#e]VP93^9.FB>RaF-e+IX:C;FTHJ+/7K:]6-(,KXXZFO9]Gg]&]WHQVES9
-6,dYNE5)3[[MBW-.Z^7PbP95b>fKb&)C6^U\A_OL1W^f8<<T\bK,c\g@?b@W3U:
^6=d(1Q+JE:#&)C]b07V+_OP#dQeW-\+M3D(JSKVR_b2NOA8^5X.a=()cRVHE>6\
PcK->5DM7a#N([JMVKU5HUJgC/@]>;bJ+2>?3S.I#\2LC91cJ[8?(80DG4BdZ8RE
+874&IW8(DAU(Y1W(?Pd<e7W>?/ad=@\V27Nc+BG/HCVRT(HSAJ.\PKTT(61(aXT
?P1N+SZZWY.(7-2)Y_E.aORcc5)FSLHOQM7@]Baeb0<A?YCAB9_XS75<fb0Kd&.?
)Z25.V:BD=PL)41PI]MTZU4#10KPSd\SK0&0T6OV#A;J4=IS?>H2\L/S_R&_^,bH
U2Wb?FKb+6dJZbCB@B\1\6a3[aLWPE38_(cQ(dI4ZVQ#Wdf@PXRdR&1cI(UC4=6_
D_5C4LI--L851/YVU=YI7:;@26EW)S[FK+S@6P\:/8=G.YbQ/+73UJFW_(W)Q[0;
YHEG#UPJUcD5HfXD5[4ZY]622+PTcF6FU[C@Y=;W=cOZS+<c6#g7/5R.@F7:GNTE
4+R]K0>N:eC,T6=&+?<ABM15U/A_D]4c_<_P?:L6S0?]?>S/&HfV=)32)1@-0eV:
BN\[Ba?c:RRK8f^U[5ASKZX?DTPB_eafb3Hc,FaZ?HcB72KBJ7E(=7cML7N2-P5]
3Nf@SX\N#,1.UG:I5X?DH)B;)VVfSUMAAVHe0Q<86WH+3>E;@:6YIF1TZ5^b+(QV
7J1MDf]eGeRW6(-KEWFH>/I.]IMVMNM6GCfJPU1Cd/\-;/;afM,EgUcB[T)7;^Y2
@e\^K56=3EdL23_YW/&c=TG\L_M<D7dM8>.(a>#_a?1WXLgTUXU+\=f_?Q6Q&DK/
Y-X=O0#B2.N29A7,:2#;)MU^0EWI=8JZ=LI(?DCSHdYIVU1C]E_bbPG#5Q+QTHc8
HZ/0K#R&C)Bd+g\dZO\_O#DUUGfC-8Fbg^+Q3FB&GSdGAGaUYIO._fT@1,+_Y#T#
TJN9<7N[K>0/+\8A\J_T\A3Ydd5Z=9,Wc/;62XCL0])\5@,_1bOaaafLB(EL.d9L
DI[=c5<=Fc)_2^=NN97?3H^V/SK_Nd.FY:H=@T,H9?S;5V@B&P?QDDcG+K@[>R65
,-7?ZQG&<>ORE#,8]67BT9C/F?,#&;ACUD5TUGU1aBX8WH_[+]0QfG0+ME<]Vf_G
<^[N5.fOXQ^?T5KE;egPJ>FcY>]R=QL9&H,M5_^I2/cCgMEN[PbcVH)BC:3RNB1&
VDUTG-ULdV9R.ObJ(1S]\dRZI773UX_640/46>FT>LE9G=]M+DId?>&12g&,\3]T
:S?_^R(@WB24L(9GPP#_QQ3cAFJc-Z[5T@W/];Ga6g(U,c8@22C84a2/<<f][6>T
+:YZYXC(e3NPV7?Xf-IeVLH]Z-^:+^,>A@6/S?)/NK=N<CCBO_NJQ<L&O7[Ng>-^
_-=_Ofb8)NH#O1BH1-O0:DQg)99R(gMCI7S>8>1H&ZEbT2T[<5c89NI2Y7EbC=EU
<94:X0.JY4DD/F9)&cX^8aHMa(NO9XV<]P7B6dZV[XGMH.KP8bA<49F>EFXJ\JcD
DMP;QcCP#5[gCT/b59O\YC4&<:a]S>,,MQ2;;f5g;LXBT2VbU76fH@?I\L);_b2b
)S&5SO\W(_5e,b_BOWb=@;X0[YVMTH(e6+H:QQ8Df;IO#X\a(Q-D-@4Iac8=3=Q5
bO5(\)EY81Y@MV>V?:?e;_30aL&1G=8\dOg;>f:,7RMTIUR)CS#cDLB7R)PV6\0[
E=:3fCHIQC>@]GGD@6V&-dXRLa3GId#@:]+@B;7XSXf/SZ<F-M/@a^\HN\H\4[:\
9++7BdZJ-a#Q6=K_cQPTCg\;b\@.#_#;#eM0HL4E^X(.._#GQVHP76WbS24F8116
[VQ=R7g;JV,6@a2(ePcL3RbF?O2,NS^?_/.</bO:-eZF7K12#U?ETD1_1\954gO>
T#K>#U:f8d@ba=WDD(&SUW(&aPefL,R6f@fRe2P.PXGA^H:(PPS.NgJ)3:,=8/0&
6\\2S\TM0K0V;Kc7:;S\S=(<OXScQ^Z2egM=R&UedKIfT/J9FEd4@#^H#cC>D@c3
[,U:@3YJ?#Ng8KgCS7dVU(a)FJNG)YTL=Sb;[[9BFQW=M80,WR5e@QXB6=-TW;XR
TY3QAb,PbabZb#U?3M51Fd);TfTMP<Y#I[]>14gac+9L@SaF/2+T?0/]<]e)CCeI
NdVg[Pc7\0<&/G=L[Q@Xcf:Dc0Q4M89Z2P#gR>>^0B,/X[#SKEVb5,8dK;G;-F@g
eP?:3+HH:[ZLM(6SH;(XHFWID]JO)F5_7.:(08TE@c6eIGG^+-RI5COf4.GNcb(E
6;P)C/EA+:JMbL)g+fVJ#TRWJ3-19+VQ8Ee/g>DD;cNN\=1^Id:O^,7Vb[6JX&Sb
ce=,(;/#IHK=F;&J^C,bSO1>CeXEQYFf7d[US7aMG)dC9GC\E3Le&(M0g-WQ]N1H
/6[=g^SP^VK>)VU50bD:@-/R3AH63<bQ>HESL\c<UH0HP/]UYH->TYK_2B^3<5H(
XKU_5.OVd.@HXK5e+5+6PHMV3]1Y\JBIUHJO?1d)H<Y<K]#Z6)#_bc+_W]:g6DPH
Ie,M7LSPgFBg\bKE9;#S^S,KM-]Q0FZ\O:OJ7HAg1[N57K^:2c5e#[2_M>M7:5LD
T;^D996@RP9PgW]aA_?LQ38QP)UOg#C(Hg]I7.]-0WCU@@L.M45FTV.IIDIXAN=O
R+G[[72^#;+7OG;I;=+WCO@FYe;8KTNb.LDbc;DNW7S9dWD;/,_DV4LeR-<3EB3b
)X=Q@@:/:X9=T>J:]0X&3Q7QcY6EbSbD1bFdD[<EOeYYdTEOPE9)0QP5(<S[)eb?
/Z@()c_##[>WS=]beE=7OJ>=AT^8&[I>B^NTZ&P&e@dU+JBN-.RYU<QA9B6HZWU9
T@:TAP-99AP5ec6W=fG<YP7+J3M^6?9;d-6EK)@O=2F#DM24SV6B#Y>O4^^316fA
I(:U+0bX2RK1<W(O#.<(6BFG8G4<X#I\U^H37QPP]eVYO67;4WR42&S>gVd&>6QQ
GBLBST2?IZ2/M0aEP1?;Tg7(U58^#KF[[(CF0:ZWAD&L:2Sa7I(96=Z[B5Wb\8O)
<.SLMO-ea@1FPe2IB#>LLR^CPdRR@NK]gWDa99.F&])gf>4?dX02V^OMLEDQPC#V
adc]c,E(8\XEEd(6MO]1dA>7Y;?KR0G#A_/8#BP\\].OJ)KMXT;#efP+.J<8YZV,
GZ_ABAO5:8QA5?0Ca:XP;JF^USg]LPc8S-R?R5BIR<DL3dQK?K2R66NEDL>]<YE,
9>]OB(CBNV?T[0=cU.bR>O,[KH:F@03;Z(W3)f;^7=\<:OW&PBfX)1BX/#]UM1JJ
MS^bO&?1:UBM,g/&C@^Q:&f[RNMJ(<D>[dgH8?HUadU1XXCZZ]LHT0DR\>YR\-?S
5>MH-SN72]-B>\_8#?8B_@<-XHAOe2K0IN;MY=W0X\6I<@I4Y\CZ9D0M37;aeAS(
,A)VDDaa.4@80N^OBYa(+]]-CG0JOXU96_/QVTEY<Pc7MXSNBSE2:C9KPRf(C)QI
>EX=\d-d<&729M?dL#?UX^,P,2.\+g>6^FB/[V2<^b.ZeQ>DeI\H<24YDO?<E4<E
?H//bI6X,QU:Ae?Z+3QOeeC[aH_(F>[aV.0;V=a_8\YaUZ0@3Q#DEFGBX-GQPV(S
\3XJ-0-_@XdUNLa&)CQ>>=ZL?_2M(_=QIXMM7fM1+#a-VYf8)<GZHC/RLMQ8GBa<
+X>;NE4dXHeU?WMVN?#gfE&9DFYdV/KHOC(5JIBV.aZV:PV(.<KBH8UP6eH,YM(b
&]-SX@6@1MB=#TZ^J6(90O?VbV8dG<W:+RODS<VWDP.F+@Z.6.F(CD4JIC(2/^6V
d+aPG^f/WJQR9LQ,eL)57#6Q=[.QK,72Cc-N65\=[IJBVgX0S=CE:?Oc,CSd@NIe
T+N=d\?IU)5_I(B9g+XK5+JAcQdU^./YJA+APS;ESIZ?KURfc06<P[[CS0GE1[LY
18W5YP\NS1;TcgH)D:X.dF8c3^ZD:gaO>68D,/3Q>U6CEF(.)INTH@5O@6&_+[[_
D)Q8G9.)MNKeJDTSA64NC,fXO\F2=VVJ(28X+(.D\(deQ4]dD8:RTcQdP=_&N3eT
gWW1^@cdI_>)0#L:]V_b_/CQ6<P+,V0)TD)PbP1QLc]^)41MW/?FU6(:A#cNGG3/
52ZQ>5B.VSQEN5,#GVd#gC5S(]LM^e#(Z7(=6&WC_PE<5ED:.V<P<3SK6G9.L\&4
7#^K5F1E<VPI1;C,AS;@.Z^6@)<Ad#d+IagdZcP>(gIQ@G9@[A^?J+3F3PYZ>1H2
b>29:M2BFSd<#=P,4@X:YbV=K+TE^-IdM2?9ZXdgOTf@NE-dLO(5@;@Zg/?GB&QW
14=^1)_R8;fCGUS(ZG[6^4YNW-f/X2bQ[EZ.&V@-O@XA1Kfa=+YSW8,_>_F?1/d7
Z3)AMa.D>&&1:WT1ZSNYB50]FZ]?XZY_;VHf]/I_QE[UFZ4@]X#M1Z_RYIZDYRVV
)>c(KT_VQ6bNB3K#82dK9P99):S=O)YW1b5)\H]-2/X7dX&OT@#3<UR-fB7\M_4A
,+N-ZMRB[L0b@O(d7eNfbP,G54Kgg6HcMIQL2dP]PEYa)<U#]-RC.X&?Jd-S/^+&
Q7FLc3HGRAe<\f[KZ[a7:R8@N99/Td:UZ7.?J#^1AXFW<bK>#Y(C)BXg-VE<0O+3
(:g:;0/Wc2>D/()9:<\.AN[>8A(+IL,O,#;N0;P@1@R\IcO/9?9QB\UBMRZNHS:a
5965B[EFFJfKVY_T13?C=M?^H191Q+5S>XXd0(T@A[)D@<.NU=/g7N((61/Aa4&L
@cEGTMC96D_BB9PIfM2]OQC[04#R>=a(>ef9\ZD7>]eQJ:bV-(LU&>IN/KefSZ](
UMMBO(8)?J/(I&Dg7@I6]6?=VZ2eTOJdOMII#VW]TEC)/31g)SbWgP8@3WRbA0H+
.W/Q23.F\A7aB2c_D3S>\],]b>Y96?E.?dcM,0CTKLFY)5Kc6P0]=B4ZfZ-[52W=
]WJ:=[?OHWPfZfRJH\,42-:@.^bBP0Q&Sg8IQaFN#&2C_g>.<LVEGVE@a0GSEK^D
3SRWC-eg7)J?dC1.B:Zg;RZ>BB>[U]^O73&IZME?NUJB[0P25,b+dHAfA4?B\2S<
-H6f9P:3Ve7B)WDRSTFS-99UJQ+e7C.4KGA16O4Q5dR_M3Pe>UTF^#8XgO@bbM31
g#@[ABNU=Z..1\cQb7;]80TAfY#F^Y>F.N=1^/W2@752KB==PE>PbW@1c4Z=7SfV
.DYc?PNKg5(N)[E+G7:F-d4;J//SK/7+_Qc;]E&Ag+GQg3H,gWcBdO930B8F]:X/
BWeHAU0]=N?_AJ3;dX[/\07WU5Z:6&?1LI04N)^]G8<=.-/:J?aZ0+(f/:<^V@U\
Bbe2@)Gg[+Q_D7&0SGB6>?e))78DMa0Y[<4Eg_4#SCKNIS^b6,d(1F.S#XMBP+TT
QaB<KL3#AMFMVX@/2d7A,4>D+)S1/0bBHNE:6[/#\c=]&-_75QQ2C3(=8DIN8M;3
>cMVQ:?:c7)VO)b9KF8-+OOacgC:&,FgGGa./a,7C7d4[OdU.=#fM0F#FV),,bU)
5gU[81.?-)Q,Z6UPP-TN&9?VcCDVWa]]J@SQN?3G9G([HR[5<N(b7Hf[WGJSFW3-
8>IM?dJ@<JK0F7\8Xa#Ib7(_5+@TH2a2-<)W(MKKG(_cbgPXfQ));,]2D5+-#aTY
DM_JZ?\+S=7=ZFE6VG3WQ<Oa++ZZ5(;6@(P._FLX17G#N(M8b6?@d(-TSXQ273JZ
CN8,BgR/MeJZ/;&+J;&M)_ZI<8:HQTY<eE2Y-BG<FJ&S_-IZ4RLdQ8+UE\&EF4fP
9E)43g2H[T?FDGeMIVBF33J]L9)OPK2TT9Af#@&?EBN<P^>?70E+R@3L,ARbXb+L
D(SO&6RJ.@FHBM7e&.A2KDW.9BL?OZ5-cc5YSebM\\[300VUbcC^67dRHE15C8_(
(C_[V&T5J30.cS7WDINA7?CR83K6RKg.3BNG5Y9A<:5^+,F;8@dW>ZgH<GeOSPQa
L^)0S)W,-,C4R=)dd,4V75RRT6V3=?-2@2O[_[DQg[;VHECOZfR^#gb3R9J-^XL;
J183YgW(eVWG39NG;a>L-<Y(@be8FDb;g:e[&,L/J[I9IfJ++&CZT1:.EK3INdD2
.UQKOB\)>7f-=AbH>4@[1(6]/NU:PVKf-1T16SBNWFU:U)FCCeX?gB+K;,FXJ7,#
TDF?+#3\/97YfO]R-==3(E6]WT>AJ3RTN(XG+@c9QJKG7SLfQ/9)I</OC726:TC.
/RA5/SBDGS5/PWEXV,+]ZOQ(.3FZ11\KT?BRB+?G-#@)(OB+3Vg?GB=62&,K]QU?
>^bP)PbLXFXNWM3fJBT;[,Y6KB@7:UG4JY,;&gM+>G8_[Q[IeXPe+N^M@d3U0D5-
SDK^47KJ=>G5,A493F7(@3-G<X_A0>c&H>1Y2AZQZdf2&Q2C:,@gX@K<-^#a)8Rg
;YGTc05<c\b#PQ8G,.+19=/YfJbK<F_GZ#)ZM.H;W5,Ne1()a@9Oc4<cHR2,Fdb^
Qc0(^[:K],PEY[P\&E<Hd>_:_c<:\ZC6;aEV/-#KW44Ga-@^If6-?6C9NWRUQ?2,
]?_SAJ-Q,-;]QE94b9X<g0^^)5?Hf[3;>d[8JY[[,RKP=C##SdAAbT-.NR@GU<V<
B\M;4)0H3CFAB\:-]MRP/6(Vg0&(Ma(AWHM]C=63IL.5_H#O]ADXb9_/D\\d)aP9
\MR4?[SG]ae:/C:5RSSN_B9\BUC@A<I(5\2L.^C:TTH=9?5OB3DHY#Kde3DUJ5)C
P:fL50^DSOIRYTb2[,JRd)H@g&;YR-J_@d)T(<B->6CG\5RRB2Ze5<)[e7f[L^)5
&>]b>ac5,D>00;DWceFeH74?O0KDaZ?TfdQG@eKF?T=_X/c3-D_WP+5;d-8VH#I-
3HO-SCe&>QA@@1N7gA7&)OE9],^2_FM56MQ8U+Da/5._5eKU?aI;T>Ud>a>PJ=T1
IM,RF1_@4]F.&fH)(fM[aMd=Rb38:<P\BA3TYZdUF9H3dM\0K\6.E;9W#2YGca<3
E47X@<f^:I?QR?CYOYB)?VZEPXR&E_>dE_V\;6&aXG34:cgY60<gBFMY;VC/:6B[
JHCZ3gMOG_DSRU1e=OCF?7DCRF6ed@764<:JQ/7MF\W8PM#e28:KV90I_CW74?#K
e9b:YcfSGe00YI-eM,b8[LXB1MNGRC;e<T23eT3(C<XTFF9fRXVd(I<T1N)9C/P7
b=P?IS@b8(1#aFY3:<U^b/X(.&+Z/+9H+,&e0-UZ&4LdG6XG-8cHXA<JA\WDA0Bd
:A101=YFR><ZZSS#N53L:)7L?E_N@M>:FN47IZBB&40D:LV54;PQE8\QZN?S_@e[
2_8f_):e+PS/AOGHT0?C)Y&K3G=?JA558FbU-UG,K9\Q3+^,;V[3@L^:N#ga0Eac
@<V+WR[++?><b:P.,COB=8?=)>=ZO#fAcXA:@6KWIUaH+G+&:AEcS9g=:(\LM(HO
-=[aAINI[[P.RUdWBS;?E144D92]&_\FC.aEFVEC7CAR:UZ&?<>D2-:a=fV7Y_7]
1c]0;EBcE;;[[GB:UW0\f+X4#?W,&bZfO[MX;a^@LU/J@(>b?,^68N,,&L4F)I8>
9Z=;MSZf-5/RWZaIaJM=-]JVGD:)=5_3PE-cDg.ZUe&Q=M\^B<R<[6#4+QYfeN9H
#E5RKPSC:G>;V/<<)f0,53(G))/TX_+[b/+HYF/Y-<U0VK;OIf66&a0A?Z;=?DWA
UeD=8F6L2H)+ENC7@2aG0^6)a;YJ4L6WG^OJcC/LW=6+D2=S;HWY0BMA)1B.K>LB
9.^d.c\F&2HCY3T,0#BFXR>E[EaJ.DY.QL0V,0CEM=&4e-0RI6:QSLX#,^E&\,\(
c9:Tg6a;[VAI3f]+<LXOLS,L_I+;T=C.&]+\g2C1dP^Q#-3B(VW//f:M9[5Zg,;Q
Of)\3NR6>:0(?D^0+/<^d6Y>4H7^A2.WXg>#4L@e0Z8IPSW)IWH6-AW6-6Pf^^G4
[VID],:L>3F;.O4BNee]BQWaWg9_,d9_PcC4Y:\cRRbH[@L?<<bE2U?PA7JVU4bY
a&)-^;_>EZ4K#JYgc+C2G8ZFeI@.3X:gGB&^+(>JDD]aM_)2153a^b3N4U^7D1)K
+-dfV3?PP(&_df#^A\dODDBNR5>&=QYfH/e8?(5Ad12Q+^802#,@dKS6eM,c:G3R
(S;E&1::S+U7ZX7TT(KS5Q8^7>Uaa@2e,:5S.L5dK?bQXNYVMaU;<X_(]-MVLQ_f
[3c>@>.fKC])7ZJZ5DW(RJDY.]RR61SW3c5]8HO28S;B\Z5TC.-L(BV?T1W^;aKX
R#9^E]R^3@1<H;<ZdSSg-)#,1R@;D1SD9P823dI,ALM,AI+4:<M6&3DWGA?R7gG=
\JK^Bb9e9L/WTUECC@f?1L=K.(G_A[SbH+123V,U\\]VNA/V[_/<;#1E&VKc+=R]
=J?A2E9bE^bVe3&3)+V][UO;J,8<WdYa:=^Q,]>[Z\<cYGK6PHJ=/K<VgDF:7dRI
+XFJ&QV9?F56@b&[g)C2R?/2,KD0R?,@KgP[A>;NEO6^PC#NKHO-A4LCEddNV=.G
W6&Bd(ZbfdLLIcO253HRE+QM2;4APcX6Ta?K<,bR1V,&L:Q?Of7<D?MBI.f/<9^b
JQO^D4YLQY1R6;G-94.:4LKWXe0>7@,9JYU[7LI]2@F\KKY_Pg1-J:A9K;H0(,TR
W6P42@UJ-BD0>21<Q1_(M>aV=LVfTaF(1Q\O<X8BafR1UU1F-&^HUBQ>(YAd0#[P
(d.ST)>,U]fFbWE;5Z;fe\gQN2.R.97A3/SPUYW^GVBB8Z>a>.eS/>@d7](04G#R
e]8Y]Z[b:7+0/,UbCZD_WUWTY/LS.)8L^[d\X2FJ0I1>WL3HU,,BH;.B,R4)=Y1&
309e.Ne)V#LCV#-0.G<Q-Y-[5IH2)L_R]\O?6>R4IR#A85XSg=;.<NdF,/62)Ge<
;8cPOTE-QEP&/J\/4[,\XPcFcRaXVE,&44)0bB&c)FX4X]QSd=E6Q2M<H6BdFX00
:.S3MP=M)d2OE]S5KQ54PA(E1#6E>2ID(R/#d\X@VC.XW]-aTb_:-J8^5^.3@E;A
gTR-3L1YT>Wf2MR#)N,/,A(8;)=G1[Ra4+WabB8W#)g77C.1bVcd=<I:2dEL6CI)
)-be6S\N6LcM#A>RECIXXDWD[7E9SWRH1QNT2#Y:KMY7OJ#U94AZePV:I=/KP8.#
.I\1JDI^KR=H>\:9W:3e\E\\/7PXgPPR,9#aCMAfDMCMgN^cSN;2>2\RIISTE2E+
/=0WDL3NeP6405A_860c>:#O)f\GJ7;\5Q@4ZIP7fMRN=IRP>CN1<56;@+N\LUE>
3#UY&A;[M1_d?XP+C&:(=_;A^D7NM8gF9Q.:edPA1C]<Ka7X,/>>OCAPdT?,RU_?
d>ccGX0K@]fX03.M-Y.;<J2Z^-?H9L:#CNNe[\Z9SQ6^d7dDH1.U<a(UXI.C-.Da
@,L&1]E\;HE)2]36EYLfI_1V+a/FT:)J\/dX9C3dQW+>^dIeU^CLcVWHgg2Vg^0A
UUKYb4cZcL8:QC6PZ<d,L4W2=WF1_]]CKaJ.,6;JQg,PKg3@7fXOIf?UK=^RCc@@
GHHTS08OD/>B@#e@_5&SH@TR@cNYP7.;C+WZ^IJ^KY[&^X#>9(SPg<;+RfR51QP/
a+AA<PP?B=4<Q]29Y)=:TE@fVHga;1,SId4KF&V)8-bed0D^6U9RC(OOZa?<V#Ud
TN=H2eY54g._92aBQ=9]Ybc((@.;Z/I5dRX&YVRU3^]LU1(]f&K3YA,ab1J-9F]E
Qe<C7cAXID]1)WH<AYL3RIU4e_-SBR^KT3c8ZU4>ePga90/b);S:71EaT]-4?YfA
ZJLa4)F\3\Yd7T0MLAbIN#8-+#S;)BY=aGT&>/084Pb2f.-/#dTI/4ICZ4aOSCOd
#6=BcS@.]#Tg-=QLEg<GYCII9QDU5B&C1N[<&<V;bZfbEQg=c>ET.^?UPZ)+e;0b
d=Q3eRO>;M_2T<[c;Ag,T_g?/([8><(_[JPQCOb?-CSRI/?XfU]L=g]ddO(,gLM.
a@cP&aZER4)[f.I8QT^-;+M+?dVd9I^OJ9)C>N[TGBFR?g=Q]4;Q+;+T<WYU5d[L
AELQVJe4/V7M_Vg3A>O^S^EEPfSFENaD&[2PRTda:^d]/NF)74[]=HVR(@.^@@,R
UR)6#XA;)D]J4PO(U(^X:?ag3;bO:P1U#:_:6_LK)cEXLWLI/B[[?WI;b_<]M/C#
L?_TgDb\R0GBY1KM<RcSeM6,;5:Ng-S(766N63TZW.BXK_[X[M8LMN;)4PK^XI\L
VDID+)NO2?aYgFWXc1ME)HB)eP+7_^f]bK:]YLZKKS<4#S)CDL7G4>Q(eSJKY=Y,
6\:#\MORe#<A]PUZ?A(e0@1=RY]BQ8JIdIFLOg[Pf+Be)<bDD2YSG]5AM^f0dd(V
g3SXI>@a\\72H(<^Q,^c;Rc-We]Zb0[8B06Ha1K.4JUTF8NM\6EP1eLY[[72@D:\
^?T]HE#XIRF@=[<0>AUF=Y..ZPQ\MW57N3<NF@fJYA\V1Sd6/a.ec+3bM=JI^@H;
(FV#KMZ[#E6PIWf&TE>E[76d//)GaR&1M>1T\E38LAc(J8/[^c:6&=[4:4?-b2>W
@?.WB->R1KB]f,^HdcMV1/O@KF^8U(:aK6&a1/5HLK8DINY5(A3XN+OD0_6R2I_9
R_gL:G.dM=TgQfPNP4^2E9O>3-W15PPE6<J96K-V./5)BbdcQEOaF.V#81ZL]d72
CY5;c<\HecY0S32bX9YEE(QfG6-X&?@0V2R7)22eJATf=SU?W#bR:YfEHO>7Edc6
HB6T0KJB-.d?TP^VJVRHaY/3#&[UH<N04?<8Z:U@g\QZ0g]HIRd+/^ddCLf9[>A;
6TG#gTLfFJcb^I+G:[W6-A29TG=P9=?@BXHMEL0]G3f/acZ0[0C5bM)]D@5.)R,&
@.Yf4M-A3WLaMXKLJ+)4FXWF5=?a\[4Q&7\B4TG&+?T=-C_7_PC)6;UOgES[1I=5
gL16b\Z2IEDZc[g/<I?\bF>]7LOP/4_?AGO+),H^(S8P9V>/CM_:dY,BPa#U:gd\
Q,@^e>543[DdNGb05@.ZW^66g,MD4/OE<C/AL2@S57PG=_eY9.5J.e)3@P@c^8KB
REY/)b?(<S7Q.167#AHRa-^X&\UK1VO)0R1GfYXIXMPF/Z.E&NfKFWIIc+B]N9F(
M[V5VJ)c3[bBFeaX7;7Y0bM9aMOT#F_1E2,VMecc.HeK+4>9H-00W<R:\=-OfIO5
e&XA_GM])P_NJ1Q0bK.31/F&#4Q1<7T-Ga9KPC30<;;8g_9XWV(C+;g-_JI3=gcP
V:K)e(S-aZPK-]RG]VbDWOST(ZLHa/4Hf]Vb+4,2E=Y=T.P8WJ5QWf,SE^49#4IQ
M_.TQ.AO5G:COK>7bBI,)#CH5?IWO0?)]562[/BeW[.1V;<OP=GDT9;1QQ)6P@/c
S)GI.)<&#0E@61BSb12-eJN50&>2P:--c_Vg_S/U7Ha9BV?C,g6Y/IJ66gSb@2:L
4#,fc8\?bR#TG<6\?P7Gg74M7]]TR;<a14]VOBUdW.e@e4AgW)C2XUb5BW8:Fc>(
W-cWZ>I+Rd/H>::(L=I#L^HM7BF/1T@H-OBC3cF1Z6f^_6BP9L9dFXW_AD)K7+?Q
YRCc9J>2?(LR.=5I\gJLP<eg?2AOQN?U[D9))AZ/QZ0:YQg+0@<FZVSJRLZ-P/4(
fQSKI+]C;bM9N&(PW?_,\M_-XV(U4c>(6061E3f7S]acVZfB3DgWG@0aM@4AND)(
CJ5<8\N>A?4C7,@P1P;e>@EAYWERBB,=_)_aRX<b43D^eAIPIG1]?]C#KW64:d(0
]G>d5(9M_<OWCa\D\?M6a(DO[CcBYUHBJVTZ2aTS?NG);9_NZfPX5:.OX_[MP8(,
>HI42&BbaJfGJABF91TY8e<>8K>,>5TC19K_G5NP>@,9X>30,e[a<D\,?[AWPgM5
K5+YLVD>K##2M=R<NR;FNcJB&bR5H6K4E;B1K?.8<_.(\-CKNH4S(LaCPXNBH9,@
^@7G^8BFb3S9NaVaNN?GVCXX[LaA/D<S:0:PG;fcgA@0+&0d=5U8F/_/7.B_&=S2
5OGQd?c+fO48=@c&WR/5ag.^X9E:KVATO39N2SFE)cCE6#KK)H;[RLQ/0=b4aY;g
[CR.SaA\EWe;?7YHZV4c_\)S<H,Ya_^6d@\1BS,+B]+;d1XcRZ7bQf@PTCH#42a+
b\TaLX+K>4JIf8XD;,9:]Wf#?.&E2NLV,X3?ACOFH97gR.[KQV8?fW1=LaI5@W?,
]Z+D=LKSL[#;MGQHAM(HZA1C?#;Z?T=2--Fae)[9_ZHI(E5.YK1,f;eH#[HY0?c=
[YK]&Wf=IUU7OO2F2SS4F<\,:H_M7TO8560<0MaH7J7ZSUf377aZKf-1M;U16W:E
Rg)4LaBbDCT9Rb6aF>R/7DU4_K1G:1;(8g^NX#Q\f#C3@41)Z0?J<P(caGKYgQT.
)QESZ).Sb)9H9D#>d_DG1+I)A@XeH3&bYV1@?d16I+HW9Xb/][,H8bMJC2-Y=#?E
RO\FT?MU,^,AS?KE)3/Hg?Tc5FVYABDJGC260]QZLc9KV+0EaF]GT@)-Je[4W2ZX
00XB3O5Yg67)cSf8,WdZ8/KIL[^)E1?EV.g0Pcd5_bG_Z6P=:=R6_X\^-X[[J-;M
/C^(,=E34gXLbR@KII?@FHVXNR8>J9INc29>0:30=_Y7QWWEL,;4CfR,_XeD0-K/
A1T8>XR](@DQFRcAH+HQ]@43OZ.f:N86WB->[<^g<FJJV?^>6];(g>2RTMVTZWd=
?RA[#;a3;]EgC+CYY@D7^SVD(KHMe[eBbEU(;4\8MN9PKeP,N8V].FE#a6;#^#F&
&F72_7?QGSYOM+CTZ\E#R\Ag#G=6J4=3\#[e2_)9PL7HBfA?Y)?B_JRJ-Y:C^UM<
AH]NfP6VFP:\[M)@Fb9XB//Q-dID?O9L]eL/):&9dB>Gc;/;E9C]g<d[</IMU#VG
QAe>b#>SIDW&ZN3^MGB<L+=L=L8e:8?:fC-?(CW^[)^02U:^US^6Uc)TS8S/&)LF
I2#0QOHAG<S8[-#\:E)HWcfZbf+_5=H2HdAcY:0gJ^_8SC+a]V_X5:cE?2>Be2]f
PB:#FY5-1T_W22+>\7fF,9V29]TW<X^,GD,[KDL_6]IV9>cRS?3=\:QM=CAM;_;@
UH_PWe3)e)Q1:(BO(228KEXNXON7NUB?(6NeR](#4(7ZUP+3)O.WY-c22F=a=6O,
4;gUT)P?A]\8EHJ1&Ig[9S]X63LU_?(FN>()e3Ag^,A:bMAVI1CRQP[cB[Q,:/a0
WFMTE3KbD8)/dKc.g[>T/N&,[0-GODVWSP=DMM08=]]0[OQC[@_/YD3SQI3c=(LJ
U@N(.;U9E3L/+MU+>Nd><9.PJTC__R1S9P?SSOgR:BMNW_<[(]5VJB>E=B0E\1[E
@fJKKQWJ&IaX@/]S#4fK\&55=gO21D@I2I1.0eFMe#9)[19276O+E5H(e@U?fN95
FRF2EbDIQ,[>ZYEU#b8(e\ROOKYd9d4#abA7SJS;^,8\FSbCIPESf3dGME;3KB+-
N\Lg:#I9DF\A0.S,N(2KND\V:_]dX&(4(dF?;F-&[MM[+2dO+^RJUOM9]eD8?0]#
GQ0ZHXbDC2fQ^#6:aCT5RfW#W1)QI+]cW6#Ud0Md?Ze[<-eN\fB-90@WZ#ZEa30W
a&De7g_3,2ZD7BD9e76eEUR:B&a^YS,8bO?L8N86MCaY&GW&2<-+aHC/08>@AZKD
cYaVHADH04&<8B1XY#SVH^VR6-cdZP?3J#_K7F(,NKfb+\Y,:b7+1_P)2-MP-3FU
=T4#G#81f84fgQDS47PUU<e4T#TW?4H;R8WM/bH+WP>:@f\>TSZ[:MSbA;]YTJf2
)A1G,75QI2S5f;F5ZV>3+Q&FUE0>0c?_d#d,&^\6e]PdKQ75(UIAO-XKG7B-\5e9
XeNGWVI&MBNG9F(85B1VJZ_TYedF(g^7O9)C2bX[X3?=[0D3+N87g+#aUL5>Be^7
+gcVJ&bQV,N?YZ_g:)Y&^eL:9OE@LKUaFOUR1^.Nc::^0XdD/A1VL(P?F./@]HNa
SScgMO=+A^.A7NgC7W?,JZ+@V@?D9RfG,;7ZAa2aK7>N80?I&2VCcHQ,T:8fZK](
L+-1JLCLJgdD[VG6a?B;OYF,dO-<;FKF#aaX^50@Fc7<F.\Y.&^Cg)&VO#&W9(BM
Z?/E\DY-]b.gSS3EX68e+a5C,I^/[ERf&)46&SGOf4L<1,L:cZ[&Q.D;1<GFMVOc
&c[1[QbH@aX[ce)_PJO.O7Sf?832K8VR:/OO6(D(6RT#IF5^MY2<Gbg0WOI?6RZP
BS9\I[@_KL[J##fELQ_]>_:FaGAM]S7Dd+-39V[cKIPce)4PB<W.dg;b1;S7OKMf
8D)^bG51(<U7GJbZ;,ZH4Q0Gg/<E@4Ad<UOb,]f&-b[UU\Kb=O[;?J(2X^gCPA.A
GS\@97Be;d5Qgcb-?(b;#=?<DZaW0KWY)Z](;604(9E0_?dR/EF)Wb_#_S#8BR=:
ROP&8<1.QH_J=\I7V.8&+<aQ>eWd=aP2)FH591TAc>F)1XKSPdN.gGS?R5C8eH[Z
;ER7/?)aL=@7G8QPP?EgH?@97K3b275H4CA]+E02<HCQM@3X=_?M30d66ELT94^L
-ZN.VZc20f4D]Z3a#UK:cL&P=R(g4];7aH]RT[N.+UX.,C#-fNT)b#eOff#FCR]#
MO.A^&Y];dQ4bOb9>B_06^).c,25D4U8^=D8@DTaAF1[b?OADLI;#G/]DYQ)^Mca
66##eFWNVgN<=4#_7?RgU47#\R26Xg+478T(A(>G^^)E5H5f>2PC?P&-U@<8A^/F
PLV^O&H)+-HBaaY=F_DcSXVC<O:+I6Jc)^4d?b/DBXRW)75G/g>VEW+D&>;(5T?a
2B]d&P.A0W7U^D(+W-8&3?Q].0=.(dBU/0TN:b[f>D/XXC0<D7UAK>WU6MdW]H=C
b3Z0UNR7&&0A.[#.7D4,<2M)Jf-F5geQMU:Ye<JWX-2QPH?Yae481YE4@URSQYdD
OA5+ID;Q/#\VQSN4UdF8<fg#7(O[6F+A3f):XFUQV=-IW)K3#>BJI]aAWE&:K5LW
72Ra67_J214FA?C^DO>_)Y17dI0@3MUO#K2O)D77&D@,PcaC<J#-VM=-6.?<:,>H
EF_P7Q<SY)@47;>M7<4-I/bgFN#X-A9T;/Y\^5e8\#7d_YS\IKQ<[02c1,#RGHO4
?LJ2X?F,8+(,d-BJ0+.@H47^VKS:.#RITFS_,U&(>DFB=(3CU8\\?80V#8TTY+,0
TC:ZXI#/dTGW-dW:]N]I/6+aUX81^WM[Pe9J^a.e+(0eg&g[:/3<BbVIP]MA],XD
Z@3c7H95TK2:M_dR>(O>V?_MIJf+.&69^11WPS>JIJI&dL^0^^4-(gg>VU7W8g7P
]U@-.a=JgRG,X+?9DV?IUREN)JI]4@)^U<ZGCa)MgU)3J^?1TNa[77BFbF1560/9
P3-LW:F:#CX/ceFdc5[_ZE[+ecc#K^Z^-3IO72MIc/aTO(dV(d]V=2Q6Q,BO:4[D
:]a7>,2FTb+N6MM8=/UOOT4YXZ+\P>U@_?9.U?6>R@2GQ.M6]V2#@MUfQ2c\K4BO
QJ)ES<-F;:bC7G@?\[\X<Ma:/YO?N/(H48;1V=,RSBfBfAS5843>cfg:c#???:T<
R>]Sb2eMVZC&GAFWO61Y-=<2,GM,^<Z)]g^S4<a3MM0C-6dCY7?F?g7c:M<\T,Y&
JYMVPN>P(d7>LOAb/^[5D4,6RXc(5,,WCOf38d^3<&1ffLDXf+20D)Q7G92](4-M
XFEXfKUV8/P-bg_4NR;]8d?f^5(L0EQd34A4bRLd^C?QN\d2dRC&d.ZE1B.>SU;^
N[.=bEK16.c]>]c6;MS=1LNc6S?=1LKaL=bb\.P>JZXGc&I2MeDU5;(8H-6EgHSF
@=W-3IRRQXCCK;=Q0\QCe1MC@Nf-:&bON?9ZQKDN/TbH>^X&[F1(\82^&aDe+MHg
.E7SZU)@VaH:YX#GEINV8-,LL+FT7ZG>Hb<.?2DY_@UF):=ZF](Q?<=7,J(fRIHB
FMWQ36KUMSJf0Qb^BJYTZ7Ub5Pg7S/A-]@M#I;5]J)S(^CZ+\F)U7U;(X6-8KXW0
+2)TdFd^MV;KCS?G]Jc#MGSBI&UB(7^4-ZB8&8WY1><PZTN\R]46JKf#//KVIYO7
6FK[e)RL7OJKIQP/9EZOQ6f;PJ/^8RT+P0)5(INI6KGY6KN/5IQRb,OE\42KHU;2
29(?&ZM/WED(KfQ\C.SUd7J>(b=N(HZWX)b&B@G>(U:cfK8IR_7-#.<R)dZ^9(Y;
S3-]?6ZJ@C@ON0^7Q=N6[^XJZ\RT^2^^>,YZeG0f\&YgBP1;N;Q1EGd#]F.-+_b>
-/31:OdD=7Z(/&eJ_Ie-:ef+(89V6\]L5#4aM0Y?(3gPL0gXWDKc^VZ^Y]S4AOcY
4cf:V7DBRXKZF@NUf=26FAOP\D:?C@C\R\_G5U6;46DP?d9IXPEJY^?_[45J>K=&
/]6(1UZ2fUOWAS),:B:S#=5M7?DReaY@0&?a2-Z07W8BeBD#LVEOYEN++FC?C]97
1Y6?DeB](.XaKF4CO&.3]CD<\?T1>34LOK&]3J.<UNOQRT27JT?BD;JDLE)V6\>_
KDB[-4FL<.W_H8FW4KJTX]:,NYW=gR?FG.AV86-AG_?QW;SLODAf_BXD;;?VLfKR
3K9C<1GUX11BgO6\^KAF\HM/;V0Q:gf8V/<LLVJ-9aK@[Dg90U=B==+L<4AdH9U+
C,5,#+8f=Y=7f.K<.[b]2P&SeBR;cTM0a51B#+2A.,@TNe^I&4H6U@R9,7;U>NOD
?P4[dB:5312f/)K(Q<:#\3\AL331DL56AGbfY+]C6CNgUQ@DD:Q=D_J]A^\aOB[G
4(1Hg9<O3MX]A_F#D.I#<,7?/(.a5G@SRPP.KWPJ.ccW0A)_>WLYbKL]?\>P8&]O
&9[MUK&(;>?Mbb,\36,1,3_7<eH0/Ac.DCJ/+H^Fb@[P5+3aM3/@bNQO\e]>/Q96
>@L>?LBNNP#4c0<^T,2cf,52cZcXWF,4O&L.6&a43EfVFfW&GL+?-F\MFYNU^4-(
328e2+1A#\F)LT.IA-=&_Od>d&)-;3E@B:_C]b&AKB(If[D):JPTcC+0I)F;b1Ua
QT1M[1O]=S8b^/NZ<([+.-XUK&)<Z-\KHgE811Y6(.,(J<aMfT^GD2HSb9,+QI&Z
Qab=/,1bEKQYG[F.7M1MPKeNXCNHDH6SOX@)TO:cfc]Yc/W\4f2\1)[N;cN5[70M
<J)\/KWG#HB6Ff.<)#[4J<\QEd67>2B58.5O_788BU&WSU9If7&74,XN8N3Z\=UB
@gGCR3-FN)_\6HUc^,MWKI9ZcZV_JS>?6I(;=1bN:@QYX\G=gIaC#T4<Ga(;EE@]
MXLBACO9ZM?1+G<[KD,Gf7^eE<.6[,IUDbC-Md-U4Z?7b;VFgGB\61G+5JTA8+a0
T-);2BfD_0U--D^>I2]I-A[&0dM_eZII/>0F0aY38Uc[G+b<>H=_cU_@K5fMd:=(
J=TV@aLJ&<6cK@YHYMCJXIDH8DJKMf)^;8WeQ=+HC5=KBCf?/eJ>^7:./PMTVX.Q
WeQ+GaL#5LJJ]P2@Z6K\8cd&2bLQ\D+d)e/6d.U<H<,CM[+Ra8KZ[BB.7/d__A+@
T]C@8FA6&P-[HLR=9OK.I>.(D&OANF2Q0XM#QY770#AB>DZ2:I4A3,?e[7CM2Z>/
C7WMQ,FfS^(32RF4aL1^6NC#P@[)4_E7cO^NN#AJ..(Y3G^M.YQ-SFDKQc?ddL>7
8(e.F8K\VE9J>H6,3=-@0H^MW-aXA(?,CTc5;-)M9K]=0.5C:[/4LDRSJ[0^K^]J
?@(Aa[_d&GBaZ?\R(/3KA6(8;72N/d#O>KLSHfH2^B03+F)]9N-)E:Q2/J@>^A@G
fN6(R4<X=/e?Nbc^P>;=1bZ04a1cRO[0dV&IW;795)X-ME(DaPY[5T[TP[PAV:7g
d5;WG-eYN.Yc6DWV)E.:a\,A6^=#/3A<?cK1[AIT<5Pe1)SBdC[@88b\D<bM79)Y
CY_OGVH+2=2AYf>F1Z44UUD<Y(Z?[Rf7E4C>:\ZLW(f=@OW_4UR.273LSaBKd4PI
SVHbd/?gTIP#80DB9)\-3<6V^O3NAGF=<:8Z4J@50#TYeMY#/HOY(.5dL\C65HKP
a]NU1C9[?4gR^d@^MVTI-^6&Y<Y^YI)<O8^+2gNG\H/gN+=8W-H>8WH#AcE]1\\C
6@>VZ3,D-#e.;9ZcEN;IP,^f8+NcHS(OFeAT]_&NF.G>dSHXRIPBR(:9c,,M0#(Y
g_ZS/7HOcc9a3]GCJ<@7YBA(B3b=:4TC9J?e7TIK(DVZ&f.43[HJQg;9Q0S_OR^2
;B#Mb4+(/PY<9<[XF(F[_B_&Y)X@)66XI97Q.:DO&<V+OA9._Df-@02WNd5+gXc[
CL.5N53ROIZ,#;R34VZ:@LfPA<LO<EKY-EbSfJ1JM:U>HO@9TO0ELZ/40Q>INL+(
)JY:P,gTR?Z9C4dFLN+1=M-UdBcRaJQUaMVMe86=Z8HF01;5[Q3R3dJ#aVgb8HD+
W[:M/0YC2NYJQgUeM-ASLIU->RB0>7R\7VZM.7Z5(DS6D/G<LLX?4S8F1<_]-G4Y
++F4V)@M5\4QG?0NE&(5JH8G#B??(KTI8QebET0IGf7UUO[_9PS)FR_C+NF4XaGD
-)]VEVa0A9_ZGW,BBc;,XC5K9,3A0cZeJ3QQJN(OKMD=,g\M5):Za#Z]MUP^1.41
.QLXIdII:Wc?^-/X6E?47_]H,_,bJ^4IfJ;==X:VKAfWSKA/#45N;6&C+3G]66X4
DJ[+WM3VH5Rf-2)R1[2LD8@7f9QaKSRfV9<;X>S)#/6CKI/)[DZ\?@Q+XW#NKE]+
D3RBY_DVcQI?aZ>ESHFN]6AAQZb]N<GSD,K[>C;8TbfU+g/ST:NI10\W<;^ZK/EP
2EVXAI6^(=@IU=?fVE3<Cc0GHde_46_0#(aG#QF8.#D@2,AB]XbSC]SM6Eb#a4Y)
9If[\1>fBgXG\(WVe.\aM@V+#/gU,0aA[Q7K&<#.57:CI>_T3:4B)M;WL#cd[,OX
5?A3_2d8E+@O2W34ZU_U=[#,eWJFXR)Q#Z/E#F+dI(T6g9]X9?<@QP2<)(3_eKF>
T3]?WS_._6UEeU4I>Ud8VP\e]@=A+4H3JAd[6QHYOZ45XKZ3:g+TSID2#beK&9@0
V4/S+g&5PB5_4=gF\d8P6VB6QeWW-INT7;6;V6]W..AGc[f<\7S?=N.<Re-:;IJA
:PCIdJL,Z#;XJ:J#H.<U,>&0.M-T1O7V07E8#(=:L.0SfW=0Ob>9KD5;BcHZ;KO0
(8F\Wf::]QPA&X&9g=KcW+;Z_6_(?-JC6MP4YYUcDN/5M:SH_/E9ZaD=TV/4ZZPL
G+[]+#_<^;Y55R/^<TT@A4/Y>T4Y/U7RD@=b8:Pf3Z[SC7CAS1D_#^GV4P2,7e+O
b=9X6/8Y@XHPb2e(((@W:4Y2b_a-O8VbY>c#b/ec_CdQ,;RP[Q;(>M[e:/O/_YGL
DX0P8+63T6A@\eBd9<&TD)/E[Va0K.R2J9<.Y7?E[>.7,^c^MMZ,0-,?M@B+#6R=
PZ_\3?&H0-]WAFH(K01<;@b#1QF52=[RQ[P,]42A36XV+S_\CH^9fH7fF6=JPQ]Q
0EA5I<&CVY+)c>8Y/^0+YdX;O,,(Y)R@DTc)N9_&e8<CZ),/<(FBT,[-2G-DWU:7
-/BD&O:d&#6KR6#VZ?(E-ASfW,9AWVY>S&N[=2.b#<UDVDK>66eUY8[/JSJ0W._I
6Z8(6@O]eWdLW)^>61Z677#cb:Z\\^<A7]Lb3:Dc0#20Z+AC>?Z;CR9e>aLKgIV_
A[#IVEcL+cB^8D\M@NQZO3(?:>0OKOB3V4F^F#][26176EPQA?81.&CNZ-T4P9@H
WcFZ,Q<1L(]@86DLA4e^21cbcBJNWAg,@-IOO<=V>bD)425/.#\-3L)>HF<dBQEY
[@HEJQ8fGO^C^.KGBN0NbM1,Gb14SQO:.#H#;&NHG^L84GFJ0Z\Jc3LCNc#1LQWI
FYTRR5J[+Kf->L@_>IG]c?L/@_I\c+7IC9b,SW,d(=]JNC[=]I(ZT><-P2E)TA@X
4399[a,;@feNeBL=N_R:I(@3;(&;@BC4>Y@OS-24\1,KBV]AYd&BbEX;61.)OS[Y
-VT?+K<gC#BF..1G>@-S\P/D/4_CO))WT/&c?bW(@2SEC/_XYa\6JTTW-fF49H0L
R:<Y=#C3d\JC+Ia;1B=4;cBHTX9\KN(.KN-^Jc90KG.SI/F;/S4P4?aLf,b^X0.X
V/AfSM.:X1I4G0:d+&#+<6_D4#Ke4[TF<,UTg)>-eK-0=I5fI2<YIEF9,\e#XI&#
KeKdVbHaaED<AIL.+WgJa]72bZTL:#gdb/D-V)F+NGF/6G@2\LJDe-a>ANM6;QG+
Y(=LOJ(&Z+<QTXLA[:)G\9]5Z8&<K&J+5Hg8NWVYT41g41]L?OGA@O5:fW6WCb0D
?A#^S[f.b:g^)g^.G&gcg?>XL=)Ib]I(I)TVN5aFe=;@P]Xb0c;VL8N@V0XX>B+3
#BI0\7,GS)Q2Xba@_TeccH&Ld+NVb=C.Z.5@ZPSZPS]L6gaGN,V@9IQ495^YNNU;
Qe>)M?fabVSSD,MCS1OWgV(]O^3[UD/8@H_\OX0Y7?DU?gO,8W?UGM,63?c+EF/O
:.IF1TRFL[129M-N#=?3YdQRYCYXC1E+;AX6K,7&a&B)X-eX//2::BPPTaf]Q).(
^aWAM_D=f]X:0E-;)?AAXIg<O=W[DBTba;>#OPV=.X[Uac>@g3_JEW(B.VZN\8fM
fJ5NJ3fHWaK+;g_S+]_R/XBX(JN_Rf/Z@^Z<TGf#>BE9C4dX#;ff=F-4JM-8AWVM
5.O9C+2@<^-(>JYdE?If\,+48[<N#f<c\Z3V:KZY=9Va7AXX3L>DCC<Mc75_]0,E
Xd4=Nb?_X5;R&R3cZETM->;2N@<YdJ9]EDPSZK<_?OB#ac&I&X]DT484dP[X+FGM
V5O^>c_Qd[1cK^IEF@_bEN\CW16/C.04[AV7YH^=N)]A+?ND&Z,dZB7K;-_UL@/5
cIFY50T#T6de5YY->OMCJ4<^4O:<&#MC4=4=__OBRU)L/#G(d24cCFA&dTaK:G<2
..MW@-7DG9FYSUFW#Y^D7NK:S<8(IJY@,Vg(UD+=S0?B,[W:-K?8&c6JJb;N(dcI
]A9=,2#3#3-_(,KN+f3;?:4ZLSN>\eV#f)Q+aR0ePaEW1@#.V917B0,7&)5CS2Zd
UC7gK-A6EL;JWE7D5(VR:8KZT^)[.6/2.(U2T0XYKM@&F2#;cS24)f/JORUFa-d;
PQCDUL9C9U<I+A9bZb6T+RV,JO4G7ZY;YWP7,7:g]g:9TNC]a]&.FS=?,4=d<67S
0:C9DL&?AG<C073\V&RT44JOdNfUK0KOQ+C(7g(S7NVbCa4BO;F,LPK+9HYgHX5a
>eOYQM4GF(-1QB=@>=WKRE(BZ.[G&cA^/TBW,b]3G=U/;YJKG\Q:KOTd;1gM6b68
</Ab96AG>U8J(E)S9EE>(d]DX0Wc>FPf8)Td)^;GP+f,@R-RZ(]<9b.R?U>#dLLP
\LIAF\1Na<ggE<fWLB70R</\D6cD>51Q(QBIgSX=eFK]9^_NLEETMAQ\YL_]S4a?
bFNSa.c7NH]JcX>JYcP6/?R_HD<_&f&cX?(E95JLYS[)VC?96?FV1-:J->0\:]Ha
34.B5T9db+B]W._Jb7&1He\<=5@Lc83&V21E;OeWU0N+e@64J\UM_.Fc[5f(PcYA
PQMT19YC:N8D.UEF<2G?5GR);CXHIQd8N^+??DCAC&^(T+ceK9-AJ:,91TU,4?/D
.Y3=^5JY\-G:eNJTHVfR5E]&GOJSe;M@bK9G&^^HK)5Ua2Wa6gH)VVQL,\>J-:[?
aKIKe3\RNEV\5gHf)UM>eL;3+gC\K?4#GdT(9b#X1eCI>XY+44JG#cX8)#]8SbV^
]I/YN-eVTe2I9d_DX&c-gZYc,=&,Z/2JFN;7>H5b(.S2f\b3]@<YT#1S_TdO?]M\
C.^2@g>;#dV]6]O1T-@F/)EEN?Z=1QgO2H#ABLZUNX3L6K5,@+Ud>HPQ=U_VGQ)g
Md&W2bMb,Og/X\QJcKETA?V)X<D.,PIUQ(f)9W#e<+PaN>4&(IZPZHfe-S8C@8S+
G8=9S8J/JJ0GXW,WV(g:gV0egJW<K)KZa^2g;68XK9CMZAC)X(6e#7F6W=;^GNW4
E(GI.bOMOaZG:))7.]<dT)g^SHc:W78D6BF@VS)#O.JAb9\e4WB;/@-Jd/-]2R[=
VbHY?U?0U&bQ3Ib@YER(A3,N8YbV_Q#),IM38P0-f9NIBR]bQBLWAeA]=?UKGDKH
.NV)XCNUQg&J,MR/U[]4NB6<5C;#?e<3d0cNYY#0)+U+,PUM2Ba5PR1JLX8F<L\B
N9FZBKNQ&1EG4<XfU[122c6e&-/B/=^7f1G0a2/-4DJ_)O-+e1K+gZbPVE@K.fb5
_PLEgZ6N7QKND8Z6=N\.)98F1^YY:c=&.=?]2f).-ZVbGf?aa+bbKAS-]4ZW;P0A
+5:2SDU]A,;L]/TNgffbY8]IC(;>VOeUC(Z=;PU0&I\^;QW5-K@X2R@;Hf7]O5EZ
;19S?gY;CYV\XFX@@GeJZZg#YgW^)b3OY)5_6,8+WST&DMafRfDI5K[&L^L+_7+0
7YYN8YBT&:/PQVH+C[?Q1?1NNU[31>T8N=9UJ\Uba9BFSP6,R62:Jf,9X[#TdB>#
EfQ[1=0]AM&bK=6L:Y@^H=;2N_1[G(M:@fa@@Rd<ST>3:>>.@D@RW>N4&T9[<7-[
OQ:[#EeAH3^]HNF+K\Sg<.Y5D9]geO)OO+4Fd=I=.a@(^>B-=U(8A#Z@eU#BDJgB
H8,SE.?9b(HN&[FE;AU)3)U^6CeX7g_>/PQU:(H](TB5+E4X8]QAA8A7SNEHW]MS
1-ZDS+]GaZZJ-92#+0JeI4.6/S#ULN0g304dUL?&G0-ZR?JRa)ddFM0K=7W4/G^<
A_,58+0.RbCdR4\dd:-[V^]K@H^Y7TOO4RJfGD?0SF-&<H<4Ke2]D^(/UD1ZD9d9
XV[cLa&+F2?gY@<@B;L0?.MY)4X7=AMT&.FW8O9+b::a(N\;TeV^7c4IDWIL^_2@
DEg#CcKK\E</@LdPS0M6LV42N6UBV->e>6P)gSWFZ,JA^#;4=)Y]VYA,D3c#<0L=
)e1]6JHM+?VcK\-3[;[MR-7/05a]Ia,HCgab+ZLRJ[?:0,e]AB14I3,fMKgZAXYV
YbUY\)PbU>=a;II6K+0b-dQJZ(gE][;#_.3)42WS;),OL9-d.\TZ.TR,X\_U&;DI
[31F/84VV(#aNG/bG>RbN_0&+-R2>?,+I)5R-B,.>8K[f>R#BeT30E^5]U=H<d0R
?5F#J8ZbK3N@e+SM-QN[J06RfcNfdFPSde+)Sf)8,-b[bZL4B_dTQG(QWLU[KbbU
B_Y7:CEUT:F;Ce:IYLB6Q-^&V)G;OP1A(ITX_bBG<OJ#^5GVDF?/P>,;PL,_bMN:
>WP&4WM5TMV4?TW+;?JREOT8gL@H.(#b;43,MC_)F1YQFb-d.X43:LW2_OD\:X2(
T#JXC^K6QL+AKG/J^ag/SIF8GG.dH;V;BRI769RQ[bK9WVQ3X&bT@>_a[.d+c<-(
YaBe>O\(\:LL>C6USZ,GdW9NXXMG_T[3L5R1RA6,>(A8KO7Z0JdF-6NA?+C[A\2-
3>3+V?]EP<bQUSW-3CMgQd1Pc@@U[fcd6V</L&_W2=g2=.S(OBaO=X4?32G=EPaR
-_)_-QKW\JDVb0-5CRbgE3g=L&B;0BL91[QZ87[Zg4N_aN>Pb6ScLZ.(Nc@WSH.[
<S-JPFE.gc\g<JZc>N^T>.NIc54L0eCM:EHKc2U<00S4A[]eg7W-\262\0C4c65=
DG_BQXEN+Z>^@eYJYF>7YAWLd00bdSS^<I[+Y7:_)4RD;#7NM38<<dN>P673MJ:U
b->5Tg+M5]/KU[[G>JH@K#aD0-e\XQ;BLO?L2g+eF7#[ER/RDG.g2/\Te/MOGe0N
9JW]X5/25YH]\L3GX=-aS/BPH2ba..,6b5Q.a(dYD:SI^54N0f<^WYFa9Ke5.eSS
@#@/SZ@b=dd]JVN:]J1:VGC4RQB<Da4ffDYS/6>#\.5TU<U2-C1SOV[@fC/M6(_5
[]5@Gcd]RDN?BWQ(M8e5;BOVQ6B6c#D\,+@V,K]4AZ_=1BUXKQZI@&+Z8:dHY05_
[Kf30c6N2)5]e.Y0YKBK&RRY7O3.9&Z.(BPfYR7_&Z94V(SR:dDJ[Tf-/4b4DM7Q
GA3cLWEF7C0B^>)&##LNGUFe\)6YFI_a_JBFd,N//J5LOCTE7(=(.<M&E[F[O&_-
e[1>\e;bS#;/^OA.?86+6G,fM8.Zc6#NKD&R:P_IJ^/,26Qb?2&G4JSZSU\g@)e_
ZDS6EJFcZRd0H)9d3EU>E=9V.aB2(\<\:e6I>^5.U=eH9IAREU6bA4>XE03]49aK
56cd/LLaNGeL#aFf?90(UM.H6Y7LA+#DQRN;dee,4c0-bSZg5D_.0NV]gcBF+M@F
_?8/:_>5PMLYMYPBg5SegEY3f4KK,PQNAYeg7Je9H#ePX4b)J@dEYWG?BGT&N^HB
@A2Sfe7R9C2__<\7AZ990Ed5U-1C]E>M=)@bR7eF@T(g,0)HFY[,NI939SaB3/6.
YdS[CL&.F(^bF#Uc<0W-eIbE(=K8EWg47@NPOG?[@E18JE)<X4/a/)eId7.Ub-]<
^27)U:L6c,K([KJX&ADSRWB@:DL@K=J,9UR21EY2P/)/VW_98?62#.dS[ELCWHG5
,5?B]&cWSAVRLe4GPd=Z)\@([;Q?3??;e0@4cY6=bL/-W[9C\dDKAR190IRE/KNH
^\WESg5UTREbC)6Q5.+GV/[e-1918+A>UaeRF:[Ve7;)UD@3XWS=I@6-WNUEW<Pd
R,A<2/F+QfZbbQD6Y=M#9@bRC5&XX&bffYV<XJ2HGQJ\TG621Vf3-f+](4=ecdN)
8_S?R7a<eRL&Z,EL[Idg\=R3H\4SD2EKW3b@V8VNAe1Q=>P(O4QP3gaF+L[IQCR.
Eg)A;JYQT(5@#_.EafY]5dFI\f-:D0__1LLdc7@F)D)eOP:g+)Wf]f:DRH_)O]&X
=aG-)>(=THS^?9?W4X?\4ZM+3IKICQf7H=&4a(<5M5CXb>A#4>>C)\A&M[5_T[X-
-]DQ:BaUYR=OJPObb-0a77QV7H]XECd(4<(fJWH)bP0]D+DCA&]@TZ&-Z(XIR[]3
/ge-@cd:./_+e[];H:Z;0Z/K#.CB/@]F4]<9GgY^7N2-Z#=;\N.4eXV:&#0d31&5
P_/8)e.A5O#J@=<A@VI0JPbFEO]RALOeZ][d/)7618I7aCJUZTH3&5d[77TYafbH
Z86I7OTd2M1d\V96BHV<RTWg\La&;5e&0GP92F:]bK,7MX<_4&8QJ1^=aGWOJ1@g
ND_ab3VL-?N/U=RC8JG17Q<bX\fTd^U?:C_/#McP#QM<[U6H7e<=UCD-F[R-),Z2
_eSR:/TXF2,MPR_:^SRVPU\WML@(38-\UL[3eENUQ^KEEA,GHF1_TKf(=K?TNDY.
C759b0RY#&7IKSSGG\XC]Dg\PS,0)_SH#8P+.(a58M@fZ8V^g8c\DA6b6A#I@1,)
G>7).K4(XD2Ce?.:QUSPBF-9-Q;+A\9V2HD;H&BDJFAIV./R@A,LZ^_bP;dU64II
Ob0);C>QVaK0CHc?BFg6ZB6X(W7)?>aaF&&]Ra#QLZ4_KLZ<L0@.XV/]5-c,bIRT
DcPgCTT8PcVJB4Va)8Y0Kd/FL2/&/Cg5TM:\TW7>Q]]WdORL6E75FPMTAS>X)?;<
ID?RYI\-H4cPIeaXS+/a(b>O5D:M1DU)P7f[_S3eNSS&R6eYXTP&AZdcI<\MF4X9
EgLXB0B<8KAc=N^Nc<.9J/QK)93G3K[V+g<eRU\V,HOf96+:RW\Z1L&-a#GZUd<A
J=-3&1\VH3#?=T/I9YaY:<Q48UA>^V4EJ3-4@M0H4A[DHGP[9^-551XM=#=(d](=
=U6G[YJOYZ<DO(<II@D=fa:ab=<M+S=:7Q=3#b<M,>e3QL8Le+0N2R:ADC09/2]H
X_#Y-8_1K2E#R0e#5D7CcOGXCWT-6PX9]O3B\GFbFK)J+;4(>W9G=Gg3a^0:dUW^
C@P9<H5<4cc.D8D9G94EXZ9Agg+V3]cdReg0\QR7##28U^c>]7L5A<]FHJ^Z#gKg
8-LB684\XGd9(^U,QTM/H9025eQ@H85UYM\JV,U3FZW:0RH,EPMa#dDI/d+e_,9>
]5AZT7IUaFOW)[^]VS7>P<[X;XYQdL7E(9G;F>S>L,IeQ^/:KNN&fDI4_3\4&/JN
N@T1bH.T9eYb;#3GBETTH;==K?[dJ:L6IMe(+ETG[67LIKABMed7M=1HH=-/E1_f
[TNEZIL+9cE&cAQ[,e?XC#@RG[_fGW#J?+:XJ))-/5d+1IOe[1cC3]fS9D@MM^4]
;\&X,-0/@0IZ:(Z@dWe/-:F2/V3J72YfTW_Sb^N-dX2:;9KbCM6(b8CD&/GdS6MF
<V?@c>84]d05,gfLQ6?cXf6Zae(eA;MDSMJ0NA8D356V]@\)Oa^V3-=(_^N1FC/?
U^d^.+/+.L#Z,Qb0?H:KXS5TL?/&]]Z2MgA]@/e=5GBTTGZ]I;-b^5)CC;#BR4+V
OWM^fA<QXLd=OH>@eb4.GE.-\5fB4RJ@U]W>5+D4220-:He>)f5@MC-9L3gdHAf7
^KM56=E(P^)09AS2FVS7?d3=G_C&W;\^b7AfCIP#H(R363.L<W5#U?3F-d,KI3eR
,Sc\0&XZZX48O3feK8BIfI>IWec(])9G.(B95](47c2O>M#[[(G]Q13@A[UBdgJE
ARUT<X-,F7#;E&B)7.#eBI9<ObD_1KgIIGL@?&-M^2=cJNBX#Qf[LC=a^4fK8/1Y
&[#F(4O_HRE,-VBN9?aUWRb@1eN1^L9[.fLW0FeGGcSASfRNNQgDf4VF\ePX.0ga
HH#W<]OFgfO9WN45TU>C&#T&TE#W?M6dDNfS3C4M?P,TA:3fR<@=FSDFOdK@M/N8
:OIZ[^[N0S.O6+RG5?^[-STO^GS3Y5?S8)+OAfEPdPIG<?JDD9>#FBPJ/Z[HKd7+
^-W6H;(>/9[&E.1Fc,.)AVK[dC?ZHQE3K]1Bb3;M).H5<LVf=LH80.@EF-E@JLc_
XCgB6gc\-3F0+<0:2fB\-Db^VBK=Qb2=1de?R2.8H9Gc@edHZgQdHS@fG:TZK\Z(
?gWIJ)4VM-M49@aPX(O4)e9G-[JQLT:cWP=-CWKNHLX21:)[-F.dL-Ub7CAE#aa/
8W=Z,dLdFA>SL]5K8Z32JD?e@YDI,-FCJZ-4HW2F\?b+@c>RN/9S#g1d+VN/;N@P
T[]4;0O.D0FXN?]82^DC=,.DIeg0^d0OZZ6X\D#TL&/5.;KcXg_&D:Q5@bRG35B7
.gJ;e-YFJ<JH6B5R(-JM):dBPZQDCCf5AF7ZRZ5@3AK>ELdQ<b/,\G?-9HO#MI8L
#/S29DcOH1Vc+@+af9/YGQ<b0N67TA/e4U8O.3D1LB0TW[(?f0.aMPFUK<0=gBR<
c#eMVca71<AcXRDX.?@^:<A&g49W77;#T5DY8OVV6U2Z#b=0/a82G1D:Mc-[083V
c;M</ZWE?/YF3(SL[#OLO[]TBUb5O1;8Qa6@^X+e9:Lfb:#g6RD^33>>YW\R]-^^
B_,?\L+C2gV_Gf^7O:=>?EB)E^H;W[-M(bZVT6]Ba>1a\;d+=KXCQEPUWd8?e6b+
:&.e^OUE^XTWQ@IgQ1FcVZ?/@eM94CAK(<Z57W1Yed8<>fLX+d;M^XaUJ@:aHMOX
_^8,O<_3CY5Sf>X.3YB2/>^^2:W/G9gXP6;=<(LY.EbPE7Se&LQd09I=X&Gd8GAc
]DfV_]cOL[M1R;Rg5>ELbMJIWMMD/e#CL@6+?9P4S^UJa9_5JSgaY>N.c08bABc[
G.6#D#-agC/8N)/RH-ce)WcCG,96S^-(WU#(f&9fJ<,O9FNO1bR<0CAA</_:FW.K
f-6-Z_cbYUW.#=AE=EE(=UfV5XD28UEHfJ_1WeL.d48X[X(AI,SZ]&/2Y-5M#JbT
A_#Y+\K.a8eAXMeC+^DaF<6a2_P#B=KcKB7eA/FNgUa2E=cTF)A^Ma/-HF\X9f((
O(QI__4ZAW-JBQ&V@\:(\L:ObE.5)7,8?e5D,-]O1-#b^TeLU(d>.bW6B=_Sd)\B
U<15VL:Ta2?P+T]_B@-<P0;3\@70+_g.f,IYCC.>4.XJ++I(G:H>X.&#&(\0gVXO
BddFXB5#N4,]?dT5=Y0UNM;CI5#.5T2BAT/^I@,Z#ec4J78);^X/=A@&0&KZAf&<
cFZF^Db<JFa6;7_Ea3^;=WdT9BO52Z93Qa@FgPcS<>.)D3@&K;AU\?bL,<BV480.
0f,4K7b^?.ZII7a.[@gVQUSU6&f^V)(L?:VII0O0V49W/eC&:T_]9aP9>_\:IJb+
ZAV\6Pge<^MG7#fS9>fB40R<A->0fgS^C=<aWJ+WO/M^?@4/7Yd7)gX6G15&NAd#
.P@P;7D9/>;gc02RZL>+W;)gJc&CcR.X9NQ+8&Lb#K^2dJU6<_HY-Ld<G5>Oe<?B
EbM3.QY13+X#>;-G.=:>0ObO)X0;RBdU/V/CX\;FMLY/J)g>(G4_5Jf?g^N3eb_=
)_?-063H&H@XV:N+P&eA-b]VEcBYM&:X2E/F0(f.9X.NON>=\ROF@c3FF2?SZR-/
=]Y#dR,:0W&D5Z(;E4).82+&ZYDKQM1M74]:&+7[KBU#8M;:YC.ZQdFe>@K&cB@2
V+_5ISI3[XE-Wd@9BHeZY8YfI5fd>.E6>TVBQ&K_K_-2F/N;##MD#P8F<RX=ZO@Q
7;KYdW+2L&:U\f4)>AOS_OO6&\)bb]#.XDda98NgR06?6<8W<dRR#M,TR:7&2CK+
PU4&UK6>>>8EdQ7c;b5VW@RTTMN0T4JHe;bUKM7YRT8]IXa--(6Fg.bg;Mc6?H_e
O=G&3<Jc<f&CabaLRe=80a>;\7H][d:bN1;@W21c@-:G#&32/QXX1(\28VG=A0>3
@Z+e=D:+c_/9B#0c\I7fIS-TFf2MRB3=O=7F.DZEc#JGe0ZEU@ZXU)^XE#KR@,9-
HM,(DR[>RLOR2GF:@Hf;OE8CN[8D2;BARgJU6@X8CWAe(FC0HX=^a(0J7G;+TDZV
]-OB]3f/6>]QKP^2;A@a:N(^;]9d_B1Ce;A-<Z6+5RTN3Z1J@7,MdZL1P[RS+&H3
6a.<@_=5N-e_Ng<?5X7[c]CQEaX^?E0-[d)SJ&YY]Xe2We@C.f(eWB6XASABXV,C
K(>#e5bUO&YAUP^JM6NPM@>U<A?]Q=[P:L#](I4LKdD#Z?0]8TVd\W9-@J(]eQ_K
5YAESDJP;H,eQ.)>W&cR+D?[E=@ASd12:3[P4#feWaUX.8J.RBL7M0AH?9aGEJ.2
HfZg:Xc(&<+g4ED0HSg)f,<B>NdB\RZ0Z5_I96)K27/1&[T8e^F/YP]@QN_8c&ZL
6@8[2eMeRF0aD&g4KY2PdYgff;76PSL\FQYEYCX;[Q8#SO6H1Kg6Q2>5:4(C=K<V
7X#8NAXV(L8WQ1b:SfJ\_1:G9<,@ARaTVMgEP<OH5#:^8,3W97aE=FX@aNV:2bfe
K6XUcJE]8.?I-5JJLK.<6M?AFQ:N/KCG&J6(O+bP+[R,G(8Z4b5HY-NJ_/;b0]Z5
-&FNE4.29V^B=XOf=YA;3N:)(VJGf1@EV6-@LZ?,b+2XY1F0^N+UU#:,;9?R6:^_
,e;WTXIeHaC.eAUO+S?<&>Sd7Nbb#;e(.R:&a/;a<5XdQg6d6D\XI<WIG]3E1Z<=
>_R?NT6CX.ALI\ZIB9b<D:)^55,;)CLD=WKG@&5<E>D8QcDL_^Pb(7(<e\.I6^?U
9:KF>@KfIf=KA6-2C=(_^Hde@]9GcR&X(?9OA<1=<#_#QC/T7S&&aFcHCV#^<L:2
-b6.a&5>=6#gDJ^48_C9?VC(ZC,KFTY1g4,A6B3VKGQOQ<8H0EYU=4f.SGA^4Y8N
:fO2J8R[C&WXX1d7b2JLH(<b]QSS9^VMN\Rc;e#AdLNL#(.8;JY0.3#5-3dOM>NM
L^UEHA9IgSe=R&ID_O3UN2OWcF2.=5E=S5\S-eV,2\B8HFEU[BRJL#L0_Q,O/0M4
3FGPO6AMB-<9?R0);<I&1;A6;.cKW1Ed7fR[43;Q;Y9+=S56=USeBL?2Q684e6F#
#+_Jg5f&Y)2b/97;Z72>=(=1^aRLU:04<+^0W@5DV#NeCMd@2>#.>T1W.1[=[^>V
7GV8ZNdRLRLPVdX-VE^OG[^1G;W/BO-@GULV_3O@AU]Je.U.[.R1)W1CKd9594-d
?T,1LIUg09#Pa+#=1[RGQ-JfJUW#-@@4T_E?)3bVMX7XWdTO^LOQ_7099,?-O?\=
+J<I7d#CG0F^[bbIKZ4BL0Ce.0c)0J-YN?7GUbfGH=Cc3NU7&(L3Z>ADXXE/9C3Q
<2b.44e@GAg0OFIQ4_0HHA^4WEXBAdTL-:fW&]Y0V?NN90f97,3]DCH>;Q(cAX@;
N6@V@&CJ]U?BN8S>YZ;/(/STeCZb^47TK[UP:Xa[7SY:?C?#>HDIZVad(U]=\R4[
HgSbM[Z278_baQ^DQaCPQX?9CW-(>67M)[A?QfD1(SPb0<8EC6,LL<EB;eR-D=Y=
0-<6#1NdfD87G)Gd=T-_E_6,\].bb>He89N-PWU3)8,47#IL5XgbBbeN_C_<MP8@
:_30Ob80OL0HM^\0.fbfJ6FC#gW]:HDe[b8?T87g5dT+NId;a1Uga-HVG4JEaLca
d?:#N>+YC?F:K>1H5(I7]WQfP379B^-J\#X#-:^]P347#E84Ec?<III3ED8/].C+
W8-6N>I6E3.]P>7FE_L9T,BD_a_c\PaT6:dOI<Z-G>T_8cd-=MNT.,\;0E2[.<-(
19Pee?&a_Q(-,I4Meg(N+>FR.M1-5\;MW&HN2+:_4&bZ>)76D5/Y]e<YDb5?D]YD
QIN>YJ9b.&RSbP-<<?/R;Tf_eZ\;<a74GaIE((gT&R6g0RXVX[T90G=,<Kf4f#,e
;.75(\-_#eXG9AO\/W)/13eK?_B<XaEX@&0TN1cOdD_U>CISN9UGT9)MR2:;^CQW
>+c.\23LRLUP1/MVC#6;<L^H-S<T1?5PQKO:=<fJgP30R4>/_BM&b:4QI808Z>)O
^X0X?IKPOg7256#T5UbIV]?;\Q[Ha]VJ80e<&:b_?cgG4Ga+>&H7Y8(UOMcada31
&6?fCb7KB\[a3-N)0U/Zb>T3-RU+b83R<5HFeRA7\A0cWJ4\V@IE1X#\^/c>8N7^
C-NF[:9MgBgVK17?TfM/B+@)?LZ28H7@WbJYYP@:KL56MV;2,&6@eTfP+3VBSC6W
RBgbVE:c+cVX@L?.:3?L02XHG#Y6O6VK9[Z85E#^_QgTBC=AS=f)?F>ed>M4]B7F
^K&eD,]QgLP.FcL.XL^eMe[>U8a]d6]f?YCEgUL@Ecb-fLI77YD-S.8<>[dKBaT4
[<;:]FVKZVQ84UE9C(C/CEe\^87)MfM>\^70<e7=;D@HM&RINLBN9SVP1N)P[aBP
0)WN:^_6J3b^C]TW;YYN<Df5cV:S[PRQPPG-/3C&Db?4</AcgbQ1SR&/M-S?05+X
g(X3(/g1WV[dF)AN?a,-YZ(V<M/Q0SJ7)WDFTMO^GDCFM<D8R/;4^eId(PXVQKF0
CU:M8IgL]1,D/8D0a16K2/W:\Q^dS,KA@)E:R_P@<](NX_V-EaG],FUPDWePgY<3
E\.H<Zd>KJ2LOG6FQR]JVX-bHbb5f6NWAVR8.]G=>IV??Fb]7@4.?>6WPVV9+[_E
5LG_b\HTZd]A<cDY@Z9gQ+=QE^PDL8O1-\+aJX;7GQGOF.]&(JA@R3PJBJYH&244
2a=6T[d7;/&]4RAD(G]GMJL7LS#?HOZ[^,K,?F0+<9ID1CMK=cb2aV-Ueed@3IL4
;c,1@BeOTQG=)IaXJO=(C5PXKe01\]8KU+C#\ZEeFU;X4>9\/<&2]UX1EHVSR2;5
g/O?^RLJ\Uf]T=GDNK?QJ&969<PT=gIRcE;fJ3/)II\-D50+?VWc7^QCg__@^DE-
T/;#,169E#R,Pc#;,^FcZX8:_CTZVLV9MI7-?_dTL@f\LMP<8F@08_XC?;)Y,4)A
520EFL4Q&_c7,SR.S.Y\H5UTQXfQdR<Of55ZT-H8+1MaQ7H371I13_R1,Lf@RS[<
(CW?aW:>.05D6D,.N\?M3@,aEE8K/U>L)G-XfB4_H2Rf,c]7T]aXYXfA.c\4aC[g
TaN(&LP]:^/-TL_UF/bM.XEHdc<3[4dR;G(X<Y@fE#.VNIYS<\=ZK(]GW3VV]AB-
<A8&4U]a(cS0Q;1WS;6LU#g93:)V#2K-CeG#?VQW4]\U\YR;T]PE>4a]S]f?WYBW
,01af._KRJFT#.Y&;LAM)e.9M?YB^\I9I2^WS_\4#Gd(#=86>gI3;)WMU1e_Na&_
^CbN@Cf#Q]ddU97VD@FG86D<F)]gNeV0a3P1B>2e\2E5C&eJc):S31>6(,9AZ(B<
4.5BZ_c<28(M?A)V8Ke>fHT5PLMB5_Eg?[NJYKG,KCPHcF52<6:05,\B_:eN</&:
<.T,2LUL+MZG#10@EA-)+5?^=KV@;b18,Qd;<MOW/[W:#(L^G[1&c>3aQ8L+>#OW
+LDHK1(_:AMKa)]Vf@[UIgB0-P?3H_<Y9E==D_,H+4>L_d-f\^eEYIR.4(_LD>2N
7Bf;&Q7W:RTJD6BU8^OV1MT_;=6,,/00B2:edC#IIC-42)+081aMO][2.[NEXPRe
Y^Z.O]V\8:YU5RZ,GQ,?A@S.7Gc9QXC)EQAZ(gbf#:C@480S=^X1aRCH+SM73ebb
(?A7:0+4C:3H^bKJ-\P5#+:g9;S6.W,a@[[J<[_CbDfP(/f&.+@<Re]DV<eWb6@U
-+0@_VSU0DdDFO3MOTee<S\bN<[7\&HT>B,9[g21F@1UO6A^dK?.N5E,74-<IZTe
[a7D@D@HM=,7?W#?A8Q#XbOa+I-T-HeC)A:-M:N4QG=:8QT0V#-A^D6bFb47?43E
M+2B_g+=f._)IY17gIS+<UbTB5R[NZ]OFXOF?SGHK?0>G#aXTCb3=O,&e2\URc@d
DSGfPULRZJ@S78=:[4a54^])g?;Z/;4ZJbQNFFB4geO@.d3dTbeYVE[VL^g(J0JG
EKWR7.Z<Qf][-]<NT]-XU7+TS23-4DVE,&Sf,[Z&29Ta:<TP./T9cH=PN,PMdA.4
-(U)=PdL=gBaQa0[@:YB:4+?^Q&Z-9L,,D^JbXU/=Dc)T=TaU9@&ACMbCL0T<bUO
H2HL[@Jc@;>+DRK7#O;;bULOR?B\KH+cJ+T/Q,4-0PKB?BGIT\Se?5/0[B1[F\fR
.J:c.A3@S^.c6QUb_c\GAdO-LaGPGL6QWTZ:L7YbSK]Y>OfF[@)(@._(NO-adJ(2
aE579)gZ@I7WZC)/K6OYC-P1T@L-T^(]W?)+F[-\WHLD=^=e(/d9N,2AWdPK<#,_
-N^d^Za34FYcB+^FId/S5/>IG]^L)/A_#NZT[/N]^,T.YD4O.W+cc<]4PNYOLS&N
A;JF);dRABL8+73SW):21:#UW[.+OZ:85#(B9A04#a>&;Wfff8d.:)AXOf0a7;-D
<EI;R,P&GC#S/[HFL<SG,I<G(V>YI5IXd46?AG-&5-eBIGV^LJKKB9gc-\9_3X[+
=GaY9gbWUd^H[-Ia7]K:YB->J6JHb9?K(M@;[0QPRP<7)L9C?be8ESC6WEg\fW4d
(90=93d_I7SSW/_=c2+]:&FU-<Y22T6RNCXK)9QKCcM_@/;+_X#&U@.=Z[OY7OBH
[f\c1HSbdRF4?PH42cdH5VY)bcJ+Z]HBX.AP#c6GJXb]L.2<@^O>;/gMP#GbT>_9
(XF,MbG=/.T>0[U@dd4.<50g#)W:5QfZ1L&D+@@>4GS4X^DS(5V___-0/XCbP+PB
>Fd3DOIFU=B>?f,4S73AVUWHK8DR^UR5.Ua7WeL83O5-]VNV]5:,/ZXb&bPDF^)c
C#4\EQE]_10CBA_b:4Kc4<Xb1T>_c(K]K>M\A[S.Y+=<4IM,feB465)3/faPgVdX
MbR32?,KXf32+>0MYd1G=+F.]^3<>8GP,D)CMMge;RWQVeE:1Y\KP+I:^5PJQQBV
YR0240W>X?&G/,+NdaG@gU#Of#8,B9\IL@^0:Mf2#..?CMW&-1H]A9O;7WDRK-_M
H/R-8=^,MK)^-aYV5Z,T##(M,3gW=9&[]T_C4-05X-R/d2RC33Bb[>N7WNf;@4LI
Y7GP>;&I4@@O<c-^;F,b,E@&/6ZN])62=;=M;^PfFaX7TQ)EMK64b2]/A-g.)4Jg
5&PdS8PS2VCR\)GQGBQ#&\=SBQ_D9cc<PN:V^aS_cNH10QaJIHEIZWa1&2]FTa<>
>JAab/&IcFd@LGH@48[1&V4-7\6M-b^cU:Y.TPNA9cGHL<\:;B+>\cN:cI3(&L#e
]Ge?E^Q;^#2E2ZdP=CeW/-SS+,VJOC/M#+E?f53J^,cNZ1R:ANN9#EeBAJUAJCWV
I-IML#UIYJM2O:)ZZacR#=<.b(7FDef/S<(3GgHKB=daG9<BWNIB?WP0GSb+P/ee
BPIP\K&9JBgeM[6P[)OKV+ga;8X(K.UJIgA^[IMWV):d-aE_K=8T]3:-A=41e/>?
=9K4JL_Yb\PI??<U6NLeR7e4H;H2e7@:7bd9CT;VN^#\Uf9WSAJY)a0gPgd-S.c+
@=MT9Qd>7_L.N-Nbf\R?a:)C9B8HAUUOQZZf9;(BL;O>gM0M<VBLQ=_=,R#@KdHQ
e-:f&X[dU?cOM15VNH=e[M2&X<gD0QZAD60B.SaGg:WgW,O?H-ABeG7^^NZC5WJf
g39Qe;<EZ#CI>0@[22=@TRPMa3NG+CaY4K#S<O7#aX?K/-aEgFbO-UPcYZ;WSOM+
d79]PRT3Z5VaQD0487EbKL/H1HW&>1^I(ggT#M:?EMa)#C^5X]U9C,Wb:GJ6CW,C
LL;6YV7MT1XIJ3>?>-_:;2Sa/87a>1dg4C8b^@_\Y2=_d\6cW0DX?PDEcK,BWWOO
PK,]VBUY:4Q0=X425c3>QT5gTbD:X3a=fGNB3BFBQ/?5H0\:fC9F5EVS9gDAE>],
B[?19)a^[R:,5&/GRRJIU_>,@Z/ZU:[RQa-7JGIT0+3JF/3S8M-;G(_?e8Da.BS1
8fR;I8VZ&@FIJ\_GeD\3X?.K7N#+^5N=_,X_<\N+F:,5NF0B,_0ZWA<@VUc[B1Bc
42e^L.#H8G#=EG=.?R86EB[E,VD\:U\_JN>Pb+>A7=]-b-W=QcA?Mf-2LXUBf67?
-=]U_K=0X8CfF<IOF<\:8L+QZUQ#M,4:--#gQQ.TN?[e:A23=0B\QE2eU5@0?\S6
\)[EB>,Z/K1^8bG]8d]@NW1\a,Fd#>F@#f=Q1ZKCg@4C>O&d+04)Q_NI)I@6UUW<
46BfD=D=5T;KK;<LG>LX0Y2]987(L/J?aTMGCccGMIb^;bgC:E&>d&bY_]f3Mdc)
7+?Eb.;XKcMIJ_DA<;+VTX_QM>93:-^5FL>,CPVC.9FL5G?Za],.:0PQJ/:#ZM<L
/580O.QDb/[8cKNN1?<&5;3))53PR<Q0[-7ACKOb)Q?fOWfb^(->EbT1K?#gZ+J[
QOgg-+C:gDI@1YQ+:d&DMX(gAa.];G@Iddb^d3RIHBDWJWaL&+@\O>KRS2?QcH@1
L&O>6:Va]A+Y7D[@]\aRO@QP/SNA5VIcJZ3#^M_H1FQedO-T#8)<4d&6G-T9?C5a
g2EMEb?f-D)?++0^T6UTebM)3\H,2d=L)fb03H_()9?2#d^[BC/VZa8M[@0cMK:Y
8BIPKEXgYJ+/g,[<)MWI]J37(,/3eC]][CV)[AW&-<:b;-V8@5WW2[<G3</La&\3
#FVg2HIP1TZ.ULLJCbQF])cD#7aKJAQQfR;VUM4eYgX?8V4Z.FA034_YeP8T@K06
/Da8e^N1&(IeKE5G^Fb0L2GC6eAB:@>/1d2/]QQZQV<LHCAU41]Z+WA&f.O4d,91
:D-U5R8:)/a(#B2VWS^0Z0TC@[a-P+gFXMgEY<4,V960D5@5B=N_4(XM9O^J>g(R
]VR</cVb_e=YUD29<I2_d&R7=JEZ_4L>1b?@,,^fP)gN]@IaQWH7Q=8fR&H].MDb
Mf;b;Z_&A+Xf&c_;?]cb2gGS_5a5Y.9_:REP6S0W(;5.:P(9TD7/SIO3be8F#4M?
?4ab,Nd35Y\N>4@FUJ5#2Ycb1T0-3X?f^/S(@FLgQC]5ERS1aV8QgVa1B8eHC,/C
[2D1#1:V>8.BcFRZfV76BI/ENT/3\S7R-E1+,B-2Z^d+S/)U91NZYJ[:Ecf9K,\8
,g4.7[@=IG7MXE&AY/^>-2a,E#W?KZ/_PE_[T=^YCP5f+)Z3W#DdU6@;]PJ2V&_0
g?0JD=.DO)11b(aeTd<MPdaH<S;PJ+76I89g?PP4I.#]-4XIH3L+]7_aSPfJ8]K#
+C;E-B>)ec0V\TdC,cdQ1>.P&f1P#g\VU(L5b/8LDgg&F;\#O7U;VM1=RV^Gb2eS
JNg=87+N.4(b<?GI?2b5IKS,YV&:-YSG1Z7g4WFaL+_GIP\^VRVb)NVe+8aN9I))
R:,=Q<&;Z7ZgPQE9?U6EbJ7N+NGZU+NAXf;R#be?X3+Ac,gO[,2H6Z+68U5/)&eI
QW7U6cb5CdRU-0c#>]0-(#.DdED>GeH&;G_89VZ?0EX<M:8LDB5>:1)B61cR0:Tf
#eX-N.>YNL_@M#=LF;YMH-K5=7#N7:\09M,TW.U<D]2\0&BOGDQXIL1D0HJNTV/X
a(^Q.V:YDM]@@WC#=>cTTV5;X[IKFEag,&&@5IC#?U,#)_S&;b76:d5d);^BR:O2
JgQ0IQP+Z-.^Sg(C_2W6Db>]^aM9^GM>V]CaEbbdV\@b4I6))XPL-S:NSF5=4T_#
CBX.A(VWcDT>_CU,\P,.P>;E+U091:aeG(#DUf1ID#)^Y.J2TK_gHMN]cG0CR3dC
c(:/I(^Y^-ea<^AOb2..:IcZNbfeBH\ZMd81-M7Sc9ZP>eMc^R&KE1dLXWg--V9B
/LX))4>X.Q.H;CDd]630)IG3,#D):11]:#JFQ7MM9O<PCfed&6)Ec\UJG>=]8KKg
Df\;Oc3e;I]R]ZTJV@Jdd:=4&XeSe_)^cJ-a5]KNNPcfZ0V=N\&FTcBBZVg):\BQ
S8#>IN8R7fU.0FDL@AP;U.X;=RXV[I1a7?0@P5@fJSM.d.38-RF<YLVO&Zg,)><d
RNMAF];]OM=#[5?U/C:[S)U[3UKO\ZBW2A\\d;2M]TfR;=ZA=aW<HXFc@Z5SHL\R
@OUV[^Jg)5]YFU\N@+I67WH,64DB;,+/KE1@](Z@@&7Q\gP);R3K4?a6#dYZ]XX)
E#HR@1FS5]Ydf-P>Q>=eE62>:Yef,@53-AJJPaX)^fFI09PG6K6]0H@8@PfbE@8N
WNPU6FT&23e3O:)^:EIe@K=_D9IJ@b_;68f\ZWe:=IMVa];BN<72S3G<7LMPHbaZ
AbHJ.Zf,+gD+BRAD]X-+3SI>(^a2SH^1+\8aVfO7g6W@#SZ(>R.)WG,J9@]Xb6QM
gMJ]d;=B/@E9K7A.8C0>D+5X&^4>9;=,)b02#L?0+C4)c@LP1#X4dfRA<FE]0</D
gN8&065WdR2/cED1\;JMDTf/PP69/JGAHU)RfCB[&E2F(b#8J12N@bb7^2;52E@R
4gH7CNd24J\0+:d\cGC,#PZ^c>,_5f+CWeZ7C/]6U;,&()[.K&fT4@9-c7M,c(Zb
fHC^-MdC,7T)FE.6Td2#D.,-?6T)T?SU;;ND;7KHU,fd,C8S0E0KeG4-e/<U2BL2
-+V(=O/M=DQA1aA[E<6)K57d@:e>0A2(Q>(dgdV8,L8X2HJI:fb5fGIW^T-&/I65
Q2cT7<6/DN8^LeGGL,<6N<Rg(R8AVHX_]2Q[KC.X<21U/0:K?1cIE26(2>Wf-8U(
L,DE86AaSCD/XH,e-\P2b;)_ZOc0Q\_CE=@?e^V1<d&H].7>N9B81Q&\6&#HW\D.
(e#6bD-B\GZ0WI@d]V]9\,UPH9O6SN<[LASd&W,XDH2BX1-ad+HdJfM>X\^R6W?F
H6;K9A;2<]QG[M+d5-.+YV7RY;WA#RC&]bVCW;</WBa].A/:3:SV_2,W)A1(ZA,H
M-[=^0;&#AXH>/g<d)9MIX7VY\390]M?J(1^6XZQbED#3Q(HGLf;bI(=:#QNbHO:
1d&3-L[H_V;>FM]@VBGK43gX+;+Y;RMDD9]MMQ5)2fb),M,@OH-WPP[8S84YJRIW
f6?UKI1+K@2fZH6?\6eX>#;+MX=2e.gAJ/\(Q58YL>\_VfY;V_N^4ZQ::JM_\_4N
;d0>N,X+KbX0;269Sf.J#U+9<<;0b4[?XGY]A@UWP+3\^Z@8^JYJg1.c1^XHC/P0
BXF<8RJQ\Pd;]3DEIKc.,H,DN]WB8_Z1N.IE9afd@MS[T,>]>d;W:A7.@4Eef21L
NW2F:g7Y==I1M?HKE[@4]WAC+cR>2E-K2#^K@7]5B<\N]?-<VN\4G[OUe+97UHU>
I>CE_?.@9KeMR1+L2FW;^F9D\ED[-c9QDdaQ_Eb_KTFLV)WGa\YBF^3QD:f\5ME9
Q1.ZX<_)&3+4eDA_Uf[1HW<7;VA00/@^K>PPFOUVXW>aRYY+YR,C4VB\N^GKNbc>
.6I/+;07O7[-bU_#.54e>97DD8.TR,P9^<:T&I<(>0fTdQacI##eDeVR7J?CYP\=
..1F,#?bP85g4VGMgYdOXGNba9Z045N1_C.Q2<@QE?06.@=H,6-\0LW/GI\ONVZE
0.VTP=eaAEcO>185-:2L,80O&SCMN<1OZ4@Z3&NAA9V-G;W]#+3]bH8<___Z,M3^
M[BLWgV;]MC0DYW8S^6[LM+)cZ8,af/CJ=-=RSF.],LURZ&P:V5T?M4&EVM>5--U
3@fKcXG;Uf]:+.,G7R[\=@KK=WHMb^cZYAUE3SW5ID;cc-8B:OF:.DR,0:VSDg#(
YB]]4e(7S87UJ7#Z0LgA5c24VZ;M\D1\Vb&/+2+^&K;J\?aG^a^W_[P2e,<4#fV)
4XM>CMFPZO)cI9SMF6c74E2(/fG2L98[-^MM<5d?S&KU^<[579S+[Sg=_cLAM-#\
Pb:1>R:b7g/aQ+V6T87.IS1ZPAH_+?7EEBf,@BG-;A\NW7[Q2V&Y^U;eMRBfcHVR
VCcES.XL91KL02\&Sc))WS0,1>+bf?+d7c7,c9g+Z8H[f\fS425@541V@2D-LT8N
H#OD/TM0P=.<ED)5g(X44++-TH8ZQ__:8/S6Q5IP6^#M>]CU]c]MPDN#FK>OUUdf
f41&Ef5,a^ZN1Q#b@L2I3eKU59G9)T1(#?g2QH=_5fC@?+6KE(H0N]cc),af4ZLP
CXIIL63M,]1C?7&QL>N/Wg[CQNGbZ0_gKCZ_6@Uf)AR7#1\?1XUG8&C@H>af<E;3
5Z1b_P^S07:_?7aAcVK\LW<2BL2X@gAJeH5&D2EL3^e4Q>:De.M@BI]NVUGC\Z/O
fOKK>OT>K,2]G1A8dWd>/08T4Jd[^#=NcYIC-62M5d+,#.YB#JG?&C=5=WP(M[Y4
QWfMJKB^Z)_DdGGS[@WN7FZOG,XLdSMD8EV<dI9VeTcX=?&KgU0_75]>d6.B0YBI
6RaRB+W+3MUL,Z^b7]NG_2Y@ca?dc2+OB4CJX<c(ND2<b]PWV4G:?d_g9?e=PZWZ
1R)(+,RTP]c5.?#[_9HEU+L.TgC0\AJFcDb\d8aeM[K<df.0KcRD>M((/,D?\3eM
E2XS[-<Z^YHB.=MV]_bOG0EET0TYad9?\XB]0/eHOYQWMWc-dZ+P48\],;C7M(1S
HQ?T./+F(8O]RXY.2Se3_3\FOfT3E\Z1^UJ\GXZ2,L-R9g,K[3U7Zf:6/NgWMRB-
>N8g[-AVGX:COb3;3V;)D@.YeaIQ9-@bLaY8W+[>Vc4EI7Z>&O)A#eU9\Te^=FUC
18^?L#8@MCZI:2\6^>Y,.=U:=+&-)4.gP(1DOLCGAX?<PCSOJX^d+VWJVU@DgCKS
DP0P15L0O./Y5_?G]079BPR+/1fY@G@#?E;cS@IZgL[6ZJM#GSWdQN&;a5A(NfZ@
H]6,.6Q/RG2=eT8aI#733_Z@68GaP90,6/AR9Y>6L?RO#e9f(aU>_#V#3Ge?[I&6
6O7,/&>)XZ<)E2:Y,Y4]UV/DF?3X&e7\+B?GX9f=1@3d-d55Qb.55;d6MfNAAPHA
\^5I@8PNU)):7JR_B&,G.7\-Q/M1-XOg-eYZHG=R0ZTdc]Y?#L:-?1,Y0)^Qd-:U
gZaTSZ8W:TLKCI-9J>SUg-J[URE,dR;5[aeI<II:HDZK,M#0<>&N#J,EVIgTI_CS
RF.11,N<T6IgC6K47GYYT.<(g8be)PAVM1KL0D3DT@4^[]5NgdI944:,.&]I5RL]
TBM3B6&Y(]O+3SH(3CT_J-2e2b25VN+,9:<AN[4LA)FLb.eFdGfZQ4I\?LJ/QMM:
=D@I&><K2J]H77U6)NZZT]a,)_@ag6K:AT]@E,b0Af6&E?17dSZ2D\eS1/#JeJAG
3U4)bc=D+^?+G;V)gML,VI38#X4cTbM&9PL72If#E>D)UeKJ<J;^<,f\VDYS5[(L
^U)7=<(S4e9#/_M:eP3(XC;,)O>XNAN-)dJ9^VgU)ac1.+aScJ,SMgWMg.Z261MU
BE5(fcC6L)&3DO&3@2AUJA&]D2MgB>NbbHbI9EgNIY5ND]+[HD>&9F\X##LV;,g#
.\6Q\Qa=2+P:IWO62e9K)A5.CY4a>72I/>/_e9R7HcL-O\R9GE^@,,T1gGX;LQ]U
EcMe&bN=7NG(gNc?CfBA)LX1I+c./50]=8IIJM(B9;c=\U_W8V_>Ge14A2Mg10H,
5H7c=:-3#888@0d)V1D/LF/,0\Cb9SBaF-59&+/&IGU?K<K8&a<2C(-Rg4@Y=NVX
_#N+\W1\WM^MKIE\K_8CR2dMK;=ZQ4J+UNV>\L/1;][724DJM^F0IceNd[MFaSL6
I)W>)Q_\3CNLP::M&YdU9/<NJ7[O<eC7WV<bAG]46[J_OO3U0cFZXO]TMY62\,?d
OgKCH]XO=KDJL<Q-\>FPHE+MO>F6:IL^MT=I/]ba?0E.#/VNKV;5?5FUBd/[NRKL
1)9LB6W+&;Q2eccM656?Ia)C.49:c,R?KW3#@5-e?ea:a0CBQ-,d?Z3@J4FN2dOg
T:aQbeRX(3IGI]2<SaB7N)#.LGa)=HfY6WT#e1A<+4/:U#Q<T-?ad\TN:K0K-d>=
O-J+4B.&JWMWHgUSQEEa?c:-NXPcc&7K0:R#bTE/?Q>8BBeW)S8>]@CZf-7_b?:1
FgZ>D:\)D5W@Y4.c(LWF[^VHg+][#(+=E-fJ6e\<==[Bg:fS:30D]7N[V9.b/Hf/
e2I<1@1gMT+AbE;cO/BC7Tc02=B7.FcV8[O^\2;GT/],R>g#PfXPUO=]69L:aX0e
,9>fLK;/f)1+@a<<W#_)2>JLJZ6.RTRg/b1HgP6B.UTS:V51J1WAPI7IbW&)e-e_
A-0YFZ[+WZ[PV98:X_bXW>a\7Y-J9#Xg+V=ff9\/>-VD&K++-7DJ&OC54Q4UM>_S
Zd-:?f/)0S#QV?4aa?COL6MB@&P?,.B[.L\7?0=(?Y=X8^>I(3LWfeLEQPI8bZd+
AVK+M#F>D\-0Z@B55BDK8,]P243FE/15O&<_CH)cOC^Q:(=A>58a,(;edBMETCHH
&fX<(8gBf,0+;.]?/?,e)>WY26.5Q)ebe.,GN>+UQG))U.-?aJQYUOg,P7g3B5LY
LG1@J\(HP5.RdIYc].?\g5=#X5bAKZ1g)8Y(;T/(Y[(7/LbV\+9,aDM5R3+:\=g?
:7aI=.>Sd.OKEJF=]\48OB:gb4A7^XYWa8-4GFO0_M?[?G@_&g+5=E^#bMH?XQ^A
Qc:Z@:W0>=^I[7c1QV_;PF/\HX;E+2e].\]_:U:?9#>@Hd@SA^[7&&4&\#f-P;HT
B(a_TT),<B)&M,b#4VSFe?)D/DAUQG?<;WLaL^De5Z5S9)TcBJJ&SYEW^I^MNL.F
dL1,EJ0X7eNC<#4>20bQ8#5cOT9Q0:@b09CM;ALV0\>V]7E\_]OQ)\?OdYE0-b[5
CA,KTgD^.gHg1/\=B-PVODG1E4MP2U\_d[Z:S@4[)/<[3ULKWg3:Z0#<LW(STT?X
^IWO;>4T<L=6eCM=MJTD<CeIUFQUD5;8.?bdRX/1M>P]Nf&?(0d9VH85-CO1S:Y@
)Kf^<)79B4=OUP=>0L6VG-ZbZeJO1_IdLV(;OCQF?M1LK5Qe#2b7[:U(W;?W>M[Q
=(HKIT45Q.YSN^M]X>ZQ;Ia8Ic1Hf-LB&g<Z6a2?Ub&>P]=.Z6V&2EPb1E:;M+6,
]a8Y0OU:[ER6IaH[.W3<H(G6WO^])F&+M77A^Y0b/(-eSP,#FM91T^T>S^XNYY7;
4eLOeFKb5NR7VH>/S?)N=C?@JFMO]I8EUU8M:B?,,/RI-aY912]e4KL9^8C]IgUW
B&.E#8S+8@@PNPGSS_5+f4cf&#U2JL68Y\.1HGWC7)Da(aEb<FgO\=@/SKI0SD?1
N/[&EVe=@9d]3Y,FP(Ef/E,S;@_K@SKZT?5TB5L1:SB;Ab,^Uf2Zg#:K;Z52E2G-
W]^GROVBH3<S.;?L)G7(Z0aNV,3be)-YTW/5fOFU-=\[eGH\LA/<3H[<V:\SB5L<
>DYM<aL+4[gaA]T9G#63OOeV(N^\5&32ADE9(,):Z/BKK<5BgBAgY,\_H<HUbGYT
+;];#KHTZM7d/RL5]M0=Z35eWF&.59YMS,SU@^TCZEGO=F\JGg8Gag[HM-6/5>f6
bXFASNF@&_.)5>OFVSgH7K[;22P1,70F&EE?2Z>958L)O,dVg,2U7bLG?LgIb57_
49Ub7T37ZPEe+==]L?2d#HLQ+gSB6LSO_Cb8FX\F1GXdZ[]=2F=/S6B)W_)&^/VS
Q/G#c[TV^=,.AS0^&_f&^f7SX#CXZ+g,U4Oe[+&+[7f7/4GeBD(0QBL<H(=DQWbf
(-K7JX^1,Y3HS<UCJKCS<.?egU:_gEbD7EP?&SW+PW^NeUgMQYX-]N?aR22(L6Vf
#-N3G+(6Zd7FG/71.95+\1#<gKg@Z&@GCg_?.MA8:MYI8[?Dfc(DDA:Wec650R2^
SNIFM5ORQ+IU@I](2B?TB?BQ>@^#Qg8T][+<8Qf.5Y1IY?G.8:PWD0cXWYHZPO:-
c:,3Y9QX?&\/=NY//CP/5O[,gPP9M#M3H_HGBTXJ/3?5-J+<(=#T73(Rf:CYa4<@
PH1c7QK97TI,>]#,+[;_A.NgZ8gfc5^g8(NdMXV.HcUZQJ7Lb<GHaRD#aJY)Q0e)
:L\E-+I]2>SS>3SV4(5EDJWD_C.C?.58&0(#X>BU^,4^>VJ/ELc&+G]e)^ZB_C:g
a5QHPa?ZK0dN82gAJXHY58I179EE_G6gR48N8Zea@//Fg\?/2:5ONRJWgXRUR4;_
/#TM#1S8f>Y>MTDb?M6IV@/C7,H#/H@7;LVK6\YUf?10UC;V+GBfVU[IK71R=2.4
cHa)X[F..0_K_R]H+XMLP7:1)DKcN4=EI98)Ofb>8fQX_Y2._f>fPA6+cZ1dK<Wg
L6AL1\#O1b_LU>)Q#^2H8XH&ID2=/_T<Re=FG<;;V?#7+C4S4L.#L<<;?YDTHFZW
/6T2+,]W2ADG@RHHE)>?A#HMP9-eRR]L\/5dSB@V0BBEVMEH5-N#H).&RCU#gY7R
e7g>^fD6W>5c4FN6:Z#T<LJN:Z(O(@d@THS,-d)=VHSUM5I1\28[SZ]LQB3fGNbA
\g_-YfR-WL#:IE)b-DBY)186FL_;/W]=62MP.eDf#=gI)0.a@54c^C,F;9HYb-gD
R[8MeR9-V-_f(;^3&>Wc1)Q5+VX)DTZb#HadM#NeKX4^QE/98:6\)ggY.:RLF2M8
YgQDALYXc@^KD5)7I&W(;g:EY]6/H_&-17eU1(&<T7:):I3BeIb9DC7Xg,+C\43=
NGOH17>d4U=RU&T;Tb6K1f3TeAB;fXDR@O-N/499]F(RRL/86HD=46TW>c;U3G\0
;84NI.7eQ2]-aI]g;,^E#.62&TAAK]P]=C^EQV^L]Q,.Q3UQZQKeH9=FUI_+RgQ9
6,H/-e(P#-PC)=O(5&+3#aJ194SA,Q9FH(#LQReP5^(O?cZC&87+<^__PeRBZg=E
d976K)CfPD25Q4YUE&NO=2c3OT<8W)+5DP7dYYAN>F9^UA?(Z-3K.B?NR2,-MLDR
eNXbB8AaY>&<O]W#OA?<2L5,#]dM<[P2^C-YBYd01IZC?b]4_AV[XI[7>\1?(VLQ
4#AKAUJcEC,)+IBZI&XPb^#>=D2FIc<=.MfKZb0>+b.?R&-S9Q((?QQ7V)IdVY7M
F[P#XRWQ2Z>][)LIYg))#ZG/4<I_/U@:]FNX\W#018_G?P90(-U1I+B)09.14DNX
-98cb.21RHN\\)35-J)FV+8.ObXO:W(L>gdC3?))]VU1H/QT_eVYe]LGf]f+QI(K
;E_5>g[?0eI=OBWT[9]K>IMTFfXEGE8K_f[eL.-IN].U./3--<B\C=)d4\C0?8S1
LT\W1FX\LbQ6P.C;2DJ9?d,O#aWEW:^UXI5DgNEaR86HKMdXRbJAf:XWD6\F7UT3
8GVW13a^abJH..;N8I<(1[/T,eM3\[W<gJR7\]X,++g5);+=JLWU^0dCRbV5^&ff
Gc@3<_?2+-68,=NO?U[K[9eRS+2X(MIIV,U\.-I3^_f:@YJ@&4QaL\WVHPU;RLB@
=(G1]+2DU/LO=Z\+,E=eWD[)1<c46>fJ>2EJCF-1IMOC5,IQfN&-QL/7d\3\>N5#
CLSRV]K7;H:?Q1/O=LY4YfDCY9E(LK(\];6LKTT(_E<#O.P,,.ZW@V)+@^(GLUS/
/K3;)Cf[E#c;ITP.7F5b,,_S8J7)QV2ZBSJZ\0&HM6bL?_]U;MLZ^(0R3<P_[6:9
53Q>6QPT+g3+1J[aB/^1]eW3YY1V_RKM1bZTaMWd=-FIU5a-,5CIJ>.1eScVI^[<
VH60A4V#J&_+^6d(UEMHa;D9Y19)[.-<,\=b9g/bH<I<E:d4/G&QcH:#A?S>5IBL
I3G]9;8A<&fW)Ec:03YVSD4G1JJ>[7NYYAA(cYeJZcWC8FRR=S<+)V4@DAP3^a?+
TTaL]NT=,]Z/HGNFWH:d(R\@XWbAKbA#_A]:V^6B952&W,H/L6(?SgC6R)g&7<&:
8&89?bQc6J\7dP.TWANHDFP_gPfNL^950-b5(OPO&CU9g64MH/?/+M7gN?WEG;be
@Bfa:&P]dV-NB@RbMRUW7Vfb?9BJ9#>7g)S(L+Y<7eD5WGHK3X4M:c-gd=#Q\XR+
A,_7b^S&d>,/e)C&+3<:/MFdRSJ^T:f-YMH+<Tg12M^bSe.8Q7=bc[FKTbX>+7)c
;QbaE[1.A,5L[HKcV)cJ;PF8;GI?F3;e7K\Yc99?0Md8?+F[E=cGALaNKS?+A05P
XN0G[M[E#[2@2KaZ3??,ff@@Wc8)F>U9^RSfN_YY3)(T?PV.UEX7e5R9DB3_A+f[
IE:\Qbfa0cZ<:egW.g:G<Cg(#]M?9H26VNeKZSC@D6\]M9)KOd\-d7g4(45P388(
^8L<AM8+?Mfb6g^RfdbZ)ETO[#8H;Qc-639R[MO&YdDOSUU0&?FGZ#P06aT0b_2<
aA?.5H=AdMVe2GM8eRd#.F)f+7EbT(9MEF2fI2XcfFf&>@BFIS0aU?P-6OZ#f>SR
?T5&\P3ZY7L87I[KaE_&a#F2+W4Ha4=6Q+\I)4&fTOdEVSI2U>KU\?5S=D^B+#\_
UcUX@WC&YA-^9GA&+1@)@5H.#@X[).<NF[fdIAIZ),VEDZcHeIYFTb:Z_35[?OG:
eU\ScgSWIU\(/W@&&F_[2EM\[gJKEOD>FC(8EW:F1L3Y:dADN6D>@WN>.TcfK<,;
E/gS0<E[U&(==]&UA>67dVM?O_<OAC[Ud5H<^f+WPAR;A\#3H8JaC4e_EGS?4R2V
NaI2@0+Qa@6eeIL&6<><Y-R2g8NgRY01eL@C?g/DSHc,>c3P9Z_A]aI);4;NeHP3
H6DGO2&6:MKKNCg^5<,#V4d0\[.;J27#0]GMT0.a3I[dA+XV#.?E3SgVg.IKMMN-
U]CFO-[ITL8AbAH;_V>@-/ZS^UgH/_I-=X_I@-\bZ^W<)d^]9&R1>U9@/M@@]ZH\
;b(cLZ;E]K=0#0JK/B3fX&7ETQ&+K)BW/S:F2C1f+XK=8dUgF.M&4(<_07CHd58E
2db@3]I6<1@BA7:8SQ^;6JQcKVNZd1RUBC,;;#PQLHYR>KO&X;1AX<XSUcT5C,C3
PeK/QQ\5E[S,dd2/1BE5OY^g2-R^KP>]&Ng-#[cQTR5:6J9L,b\K_HVRTXe,R&[;
QaY4W,.cK;Ic>b\;069;NY57R:M]Z2]7\dI\eZeO869#+P^H&W1BE7KB7N3aMd#P
A=&:UG;A4^^;)\<1ZbcG20\QZAI[(A3cI87,PA2BV&=::93+8FC@g;1L[\XLYIMa
L?@;c?]f:d83dGO)X(7SK0/##fQ>?#1I.47D@B\g+8&CLJL[3B#<dWAS+/&5<JRf
3aMA@DDUPZ>L?QQW]6_9EU04]\(R.YP/=J<^E4dO9(5E9P6@^6_:QU[\\Te)8I=I
S@U3.HJ@2CG,EcZag@_?LNbec]gA@8A@OL;?e0_.&>G8;,>=^g<=g54@Ad7;4H_2
^QZ@K>+FQKTX:d>BS1O?\-YQ-<V6[>/\#/bJP]F#6)M3d;g6BWWP]<0=OZZOM<HS
:Vc5.]g)gbG]O3@aEM@BPQe\gVVG=BC0G=b@1U)#-M\M&1V]2fO34#KEaKg(4a:1
4EgJSYK]G_.B9EO]bOcP@g5K/UP6g.FWOKSC\3:cAZ^Vb[8e:4()cR:SDVT_1<?6
34PP&+_O1ZLQZ2d,).OMRgS9O#BI)KCI@+MZ2T07Wd@&LOPY=F;K)da+_=UK#8Bb
<U;8(@DMFbS85:-ZPf)#,#/7WA4)AAbY^)ffW;\?43\:SSL+<+WMLA8@=3c_3PM?
AA0]?IKa,#;?@.S3Lb94;3<ISd1d]D?N-A)2ZNaVIVCB>QG@UW<P5[f:YIR/?BVW
Y-RNc<CM@NZ&3@)XKX@Z;(D7\ESN=Q6:f&)#PEAKFa7W[P2T:Q4d70.XLY;VM(-;
4Se[<(Z1N+d+V&Ra1KPX?IOd6.<9IB(BP<cc9c0]W5KD+6J7Ib#69?\fX\5W&C^4
VW5M9&X>,FRL_K:)]TXG0H)?L(LUbV^BA<XUGPgQ4gPOS,:[8J7Ld_f66fP(<?Qa
+?eFTYNS&??H\2eRA,S()O7_ME?_C^Q:eVHXE-Wc2M[AY?=4TFBL0Rg&6S:IWK=+
B.&gV2YJ.SY5e7PQP8eJ</B-)@.AN/JBX[,Z?)D->N)7K0a9F/f8c2Y/<F[UU3Z9
3&-Y?dM4ZTJb,#<JIKWQX_M+\b<74(#\0;V=(^bQMe3HfC&[a83DcELL)VJ1E5QY
]AeM2;3=S/c2WTfLD6F,+Sg5W6[;C=:Z1R.cc,SPQ=&a2TA^6ES3fe7:(<L,\G1M
YbE;ZB_6208e)[#I,-;6aIBJ?;a?a[2[5aD>fE?1Z>@FM(M9AgXDD;fb#8eCVK/#
V?)g^9F,SeEf1\X+A:&A/>L;PY<K.4=6,Df+8CdUEDfMJAER83[PI4SSMVHF9U@C
#^YA]^251B\E&D7_P583HD5,<APP[RC,J\S]UdC+K5PZVN=+Z6ac^ES1EP#KT1@H
&F^Ef^G]/MW,J:ZY;0EOda>=>OWV3<^@>:L4B_;&HYM_f_MB41/Zb)I;NOOe#BME
CLA/a(.[SJMTY[-SCL^12YI.b;3A)AW^bORY@I=KOM([7N47VC:V>Jd\TJ/aC]?3
VXIdE09M>GK>00U#VQALQQa^6/MRG<F2#IWSN.V8T3&TI#dU;#\XGe2H<S3LJMGf
3Y3EH9EXA,CX./Mf:\e.^LQF#;5Y0/T:8QCER#3AM+dQ[5LgY5E8e.,f54ZLe>g1
b6>1f5:[HZGM_0BS^]XL\@Y;1aFAS(1A,KZ.]]8PN(If5\bC72O#gS@0PVfA9+TN
1<W@;P)L3H3\E7Wbbe\6Rd-8H\f]2TQI;,R-b+LfY[\-)2]QL)b^;eTMUZc]T>8[
:J#fQLWY9[dD(YZX:dOXK2cgIc=/3.=[L+fR&7VDb&L+21)d=@>3cVE=XEU]I57:
2^C1:<JL/b\>CUcA@^T5.NS?SF>K.Z+b#(d0?3..[?(E>-W8J3LRZDH9:&(\N7VR
4<IE=<cP#<\P&9V^-.&7<=_[1+Ab,2&D.3F]c&M7S5R]K1CT+XI&4dUfSD9FY><2
Y@NKKWOHI1V5RFc39JG[6&d:O;KJ>S_5U=W/J,1dHHFM&=6IdX6:+?g,?MYMA2G]
a/d1[@A@]f4A^K@c.gHH(YEf#7>F.cAHgE35cCd2Jc^GKMQJcdTY,aC0-AC4,gH)
1/PGB4bSR]N1&8e/C<-)5Ng.Z;C+C[AXG714L1KF5e5U\@\eJDM.7CgR_[X#QGPG
TXa.]K7.f,FZddN&SQNPW<EaeR-\d+baEe#@fdZIEaI^^9^ZDC&GJGXe^;b=TZOP
\-8SP-I<gaXMU-7X2@V?+g8HC4EY5O)^Vd:6(TF70beRZ#M+UbHH66&b3#SE0aY8
Ec)GL\HG\3SC]]f(2Q,WPIA6=LGEM1,WT\[-9J/L]7A-Z6\WRR/3,][93.JJ5c4R
I8V7S5E)KC]0)fHTZ1=V:V\DD;fQBcgB697+ULG/LJeC\TYT<5UEG@(GORE[,RC-
ZIe(D[fGYB7F@0WD4a+;:3K4G1P@eP+Z6E&Ad^:fBgYd:+9,@S/0PRgV;CIXZ8-e
+I]OS7)#dS&<JAg_9>_/3F:<LVfHQXHB=@T(;RM:)C\KD?H.RVTL5CHg8Ib67VCa
M(]MT5FE]9B)93JBP&34=[_[\&#;dLbU.3SfR+A5;V(_]DdFa:0&FRKVOFQ+7adK
[@<c[\3L(K<E9:\U[F#Gb<WF>8T2I-)C<,b_Ae6,#I04Nd1f_.1N;W-:,62M^4OX
?JZ7[I2BYc<8G[:5HNT=6BJEc<O:4Cc6JDS14J;:.(<<C-5^R<(XfP:L4M]0;+3?
L;?7D8O]OR2Z8NB99F_NK@()7CK2G7SRT<WCf;L[Ee/[[VTH2-?Z#RD,ATRW[THI
b@@0[-@^+LJ_;4eH3FV2.@g(aPES38?#24(_I@)fK+9afO1LX;?-=.)VG/cX)GaM
H/5O/TZGf_[Jf2=+\a7X.5dKX_BZ.TKd0:P#eW?GJ/b_SDbWO&P)7R=<T]MLI=4J
d&.b:2CD^^eUB[5Pg6P-+9cgK).<a4(fIc]6&a.SY=M1XVYc3&D(Gg,#(<.X4\/F
96Hb,TUEIb?S:b&SIaf9+&<MMN[b1M?-TV[Kf]&e5e05L)UATRGF\-EL0=N,2a7S
&g:cH>6W\Z\KK@<cKY2ND85WFC>?0^,0R7/0Q62G.^b(^=PbA_&#^7746.Y66C9Q
5#J?eX7SI9<OQK+ITK1=_.?<7/NPb.W>)A1F.]YRddf(GCf-BL5V@R2<\AJWICI.
S#\\Q5A_1.ZT].BY^b(db/\5VEDUXDK_U<gI;d(N/C7YF9\W;GH>MW1g]NO\Tc\M
))^/C@>9PU;VP0eE:6N>40=Yg/H4(UTYQJ;e1K[?#61-^TK[Xd[N9<f)BQU(eZae
cP&F&]B3ObS;)[@_PW7FULAe1ENZUb+ONS_e=-_S#C+>S7\6C@)4dE?BQdaTZP&^
\FJ4#U^@I:f?&N(Fb+W@;YDWMO;6?_8NL,@:ePf,Q@JfT4Id>Z>1?C^WH^Z\RgJH
7F4#S>NTT_/R\D4,0OSE_e85gfMH-T(>0f?8S1.MDE>G-8S<7O@(\0<7Fc/V^^T;
]fJ)(\>^a:639V0IQT12_UF30]WVG/;^abAGdIM2[4\SCe=PDE7Z.#J]Z+&YU7L+
+TZc9._/?6gZY\.^3IW^G3SbJ67\D;ff3NP+U[;UPD;@VESGF7I<LbVM.bg:=SAO
K9\<:JN1I:OZDBLdJa]bS^FDN,N.>^A]WQ7,02YbdcNOS3S12Lf+TG09T>W5b@VL
NW<gf2)2JQ1=V]Q-HNMVS:)Wba1VT4GZg1LMd[[0KYa[58V,V#B:I-F@1Y5+<WX&
5?9aHC6Z^-_51X[-12-RR>I:3d8H0?CR2J2E>Y<W0BRKGGFJbTF>@]93MWWO00Kd
#\E(H\&B8#A\<f1G#YL_W77JAd\IX1Z?O-:BJLE=fKeON^9NE#TGR4,6/MX=5PKG
_D8TCP0YV@SU+F_HRB8+M0,e_,PY[_^.S-,OUYf]Y1<3d]gF=WI3-I:^R/OF:c:6
6,YDN,K@7/N@6c7H1N<O^Y3Q2Ke3WL:@K??VageM2^3E#^09B;AUBgP=dCWOB9aC
OHZ9T8dQQ4g3Q(G^K0>H7L8d5P9N-YGb?LYG8B6#Bf_3#YC322^U[C7#cJ.:QTfG
X91Z,.:_OY0)^2XX/e0N^D,#@50)@2S99gI^4\AE2,_?LfK>XIeX/3]EHVBY6bEb
6F53TKE55H&5aQ:V0(I2aO/7_P?W)<44GL[U5>7UV&7.\6<4>?KM=;6A^9DDNN3]
Z,afgfeFJ?5e^Db7GC;S>CDT>AMWg,9A]1\9A@^8V:Sb>0c@b@2g67R3EEI47^LA
F,KaP3YY40IJg[[+C0:aL;e^\TJ=B(RK.+JCXYC^[GA.R\YQWJ:Uc9cT2b&[=,<6
cWabL3)(:9Aeb.?^P?=^1S53Mb81cK25fL)7g/?UQF:37fQ@7?;gF5c9T9GKaW51
W6.AL)O7-gZP6MaD/W=1>?AE>0c=9dDHB]).I5N0^Cg#L><T#8F:[Y27@.@F\U/V
@#EK13)HZ8d>TQ8Ac]7X<M0<dP)F/3SI[2f[VgX.O.:d&OV?U(B^XK&7HgVX]V+2
P-JS]^,AB@a(=EGSHE59=8RNb^JR.)-59.U4bd<\1aAN-W,QV;J#U>=2e=f\AfaE
+?SOFeM\f9fELF(F>-2,G77Z92EV+3BGG9&AOGYaA_OA+N+Y4YdFM@2=NO2+U-)[
7S^NISDSCfMS6/PTO\>17NQcIH&1Y#fN-Ubf@?.7:X5J:a>BRaS7&+N9H2B>@M,)
&6;HfHA8Se@^]G0>PP/TK8,,D(;fEGB(-b-VdBF_dAH&0IN67a,#,WZ(d=fge?,7
A[36.\9A)HMVa<dF8>,7R6XI/C9?7)9;?-:)[HK0d.Q?^_8J+dBI9PUDO94C3ESF
D+62?Z7_#08JCHgV7SM&89/M:.VY0V)J7PbR5=L75_&1G97/L+;A]22fHAO:Ae[7
&VK9+Q#E#.1+Bc&bFU0L53B6B+0;Ufac6QRCL@++NJT_-L4ZFH<;F\#/D1bJD+[b
=cJ[UY1TU1J0GIE:@];?PHOTX).#=UFY^COgPH>9HQ4?N#QT9T<F.DFEbIfE[P1g
5/^+L5EA?TR7/V_Xd67]#(G[g&:ZQI,Wc]dGZ6L;QcYF<DRL/YfK8P82(=&//d[6
IA>;>,P.(b>ZUb?B\QaDG1:fAHVVg_8&_->@DU=(S=R#YNF\/agCDJ34\)1V=2Xd
VH>LTT>5L+U3.=X\1(&0a\#>Ac.;WRYcF\E&_YG_9[+1+OI)5PHa(g>AK.;^I68J
M@fg1O^,DK.@OG\,b=0W<)7U>:f?G54\RJ3]K#Icg,Z;@gS45H+-6#)HG/ef4X(0
CK&AF(AS-7[&:eK&?,eOa)5.cdR/O3^V+eB8_MOJFSa7I(\H=A0()KMCM7H&7-AW
c?7.fTD(&4()3_RN?:B#A4a[1[KJ/=O:&J,:90Cg##D.W(S:Q8-b<?>D_\_ET>fZ
Ud3IM;7>,fge/LY:CT0BYKJCD.WS[QLfS(B9DC;g5H4dI-/d3?5]J>WHY[YPeOZ7
A:T##S5D[X([7Q1H;NV^cZ<@eJ(E7US2>3ZfPKRe5aB6Q@K+JXF)4<9Bc+-:HM=0
98H@3UE2Y8c\/>4(LRB/N_N+@NLe.=[4NBWH<H::/?IV9+=,df>A2V-9YEc.9=:U
FM[)5)I(90A+:-3@0ZM@9@f]TYUSXAMF[;4PGR1bY^XgF1SgWTca[fgKFfAA0ebZ
G[YI5Ef?R_6]M^O-.WZ^<J3,_d\-2D-28#=S]V@U52ZTg4dPO9/ObH@0P:1,ONYe
NOdTc?\Z?DP+>BTS/#BDec_?gEIcCF)Z3;J2<Y;&]:aXL.)+P1#IYS5de@_g/6d#
THTdG8-MA1#K69/9_4KJFcdV6K4.T=:Q85I;-_S2Y54<I<Y7[A0>=OH+_FPO/D1U
V1M(-55,_XY0IXF:^,IP_&Wd)VLOO,_ZC8_-Jg_bb/O0+CaeUI?eCD;N&+U<R:T)
AEBGW7dK;aMY[f7TIGTRX_4E<0&A6,F+,Q[2A;X7@.aZ=ERGF?fE4\?QdGT=^Z[B
T&b9fPA2M7<EAS^@DV[+g\T#])6X,NP<ISK[8GL-MN77FM6c;A^?XRU_,C/;X;2&
f\(O\W)fa8Zc7e4ZUK65a,ADC@?b]@DHY85J0C#]10de04DHOUU12g-_f-bB^fB7
U&D(8GNW(V]5eg)Bc16UQIMbT(1^:8R+<K32+7RfD2DN2P/fdC6ScDBPGGf@[CKW
3PRG1+4Gb-@dff<gT4OCQ)(;KIECd?AKJ&X5(Q-G7DCc-Wf.2D0I58gMgAcUefH-
+G-]/0Ba@?MO6D/ELNG;D+QU=d\Vd4)^OU?Z>ca:2UdVS,ZRe@(-Gdc7aH76\?8#
;dDJIXe&#N(2BeD6[/XE[K9Z[5,\4XENQKYd,c?1E#-;NHG_6\9]QPT&[dO2375Q
/F:/F4^MKJAPCFT]Z6Y&IM>gVO;)QT_2O:1QUON/.CKY[c?)/8)Q2dXPY_@MN0\B
?VTf.NUA:5f8XC5\C8RNML-]3\S+/2S^Pd->+/_[J&K(.CT5Wg#SRaW(TUK09BF0
>ECTH\X.RF;S;fP^@J93Cb2<c>34^JXNGCZa.a0K5B4-7QHgA39QJ7B:<\Y?TRaW
D\a1HJ<MA)c?gEQK@;)<^M3FP[Vd6JP>gP/?EY,7BQYD^_+[0.WDfQZJ9W./cHA#
XFKf_PbcPM7#Y]1c<P8H-aG#dBYW;.>M14:MAdEW12ZfB.=4L.EM:\YH]EP?)Y2]
GZg;dMfCCfRWGb[OWMgQM:OLH3a7;cZH6d\ZDbSbQ<bF[43-<P=V.?M5IAba<894
1Y-fX<^H4.,U;eKfc0>/@IQeOUXL.^Wa\b=@NGF6&dgU]N9.S\7W)[RH5LBF9bI&
J\)1VI1]_J&5b-f41bTWM,d,EXQB+<CYV_D#Q67J\b(F&O2e99)#.).@4ZfU9\ZG
dJZH@g+I#gP0NH.Z;WF.ON8@e1<QZ<P7?fDbBKeSdfR8@L4U4=H/4_L:<XSI#Q\A
2#d^CK/7Z6WULS/OCId+c.]PfS(XP@Ae=)F99>cdD+g#XFd5N[^6X=<&N7.M(\_S
d/fXRf&c[==UR[+4(]LSgeZ\(+@(3.SIaMZ/::Q1N>Jc&/]D+g?3g\SH0?XB]G5@
_(0(LGK_76Wc;aOH3+(5+fTQ0EcJ\141TZU(Y/E\I.LC.V\V/)b6O2+IVU@0?XB\
C(R@[KV(_d4D_JcX,^G3e;6(HLUG@#N]UD_3Q/BIC:0?RE2@.2c.^1BE3:7R0L86
(WNBU6X@dbf#^MFVS_Q01]A?LYY.bV/WOc5-1FV)ZL-;]CQ/]PKFR\E^Z+;#.9c0
aZW9dCdaYaN/?:_T@K6P7=:Ma-?\337G@N&MT1V@TaM<00b\Sf,cXJE0E&:\GWI9
-(,-DbIK7Tg7KS#M=)BVG4V.;ZF(1MM:S0](\KPg1EX)UTdO_X.1B\f0Q22Vg]YH
#;M[d<c^N]?D9.PDEJ8P43^1fZJ&5N(+5Pg-^46.?3C@]T^6;D4A+1?[SRHYHb),
3P&18:bJ0M>=61W6L1Y0V)dCH<Y/61KMA&-VK55BdIPM,5cD?IG,e9g+&a?E>R79
TREfU2DA)dFW&S>6^A5If4&D4I.;^RBJC44)=FRVg>U?8;f9FU?JVIUcA.7M9[XE
QW)a;FO@^<6.(a;54^(SYSeD1YA+N7=B1)-/5M@#Vb9NJKFCSZ08BeH;=96^:.PO
]fD=W3W[>0:V8X:24>V(=)]d1afE,G67=QT2GG]=4-6KFPHBJ73(>0-aSAdR/8K5
HI_6_IZ<)X9X[N47^+4bHKGb[Y)L\B5<Ra4PQ\UH4aMgH=?-3A1fKc>H;C]@76=8
#CRL6:DS>6N(G6EYZ5IK#cE(90K2)Tb:IKKZV0-D8R84W/KF8Z;#FP>aI+OE-K<Z
-9O=9C<.9#f1>UUDI?-be[YQDZSTea&gd[)JW?9]_S0,O@/ULFZO))^&+DJ3,b#A
7d>W]AeQC^EaP4.4^I0f.\@U/9UF:J^aE#D[cQ_TP;,^[@NT/U@:2F7CR+\1\NN1
2MdVQ.I>CL>R052PbDg23TaKVfSS/dAHTM(PW/PHfGBWQCO>6\2#R;#5cTN6aDA?
VAJQYV-[Lcf8>)a\X>48L<BRUHL9@-:B8?C#RY8@NQY5+=X[PCYFI\9gLWXE?K:6
N:X&3<@dPMg]?V1A:QbS)HcOcF;W3Vb/+g9>W=Z92ST80F>g(?&af=?K@A))?QQY
^D788M6P6YD#<NZXJNb&^]GLLFTGR]:8@C+,F/H2-7;eMB29g,\TM8fPPK<4L+(5
^-.>VX,N7P?T#FN4?./T-4&[S<fS^&7IK/5]W#1,P3b)W(7BbW<b+b9)@OD/^?/X
bMEYN.U8MTT9,H^>6^JL.UC6E2I9aXF7Y\/]A((a0RZL.84:#L@A]8\>J&[8A=(d
;BQe#RK<307aHH7cbMB_@:gEBMgQ2ISWg:KTW>\)._7L+&Uac+.G;AMZGa4&:FHM
J5SX;28;TMN_:05/cBaOdI).;_,3=CM+fXg@<6Z3(:BCbRLIVIQ6,I(M:VUT0D@.
0=QcN:[.ZS//.Vcf5+Gc]I-]6V6>J#e8RHbc(N;eEU\17ZbPLe7OOW4N.<LF;497
d^K^\WQ<da3YOC/_A1FdcM##5,AWeIS/Of9/IC#Z[C&,7[XSE&A4)X-Y+#&.+WA:
&?BIZ;U5J88NbZcT[GQO)Xg67QLW0^/C_NN-5?>\dBNL05c349LJ)9-7R\2ba?FY
Q</@J2e.A9)2CQ#QPOB2#fe#?R.?7@+bbE]K0@CM7O.<?GaN:bA5E+OYM<_8Za9(
?W^K3KAN>ePF8KY]>RHZKVL&B?)J&I4,eOUVY)C-IR?ca&I0ARSe46D3DDWQXfFH
>]4f&)DR.DLEcfJ0ea7[;XIbB7],9R3X+A\;^;ML;NDeR5<_8L:H)^-ONVS>DIb&
Y1);=Q8^.5W?(YfTGIY7.S@16BW)>f#<B#BB2<Xe?C_9_-.5CbL&c5d8XSg616[E
I31@>[<[[M:XD1,77c-XYH&_8N:,@&576S(]\<\+SA?DPfC5;9WBGFgMMd3-L1I1
HE>#+<@cf2Aa^3B?QSVG0b=HF<FaML7=>3F8D>4^1AP>^7e5:,a?d)aX[@-NE@=W
)J35/;=^)IFFF77)8/+;QABCK/YD-:[1A->PQ4_=(W&<OeUVdb=.)BCc:HO^DOWS
8A;BDN7\eWe_Q31].d2Xa\[6;?9]>Nbd.M6\W7LELPRUG&+V@&-?EQ4a;A.LN9S.
B8TIBYMYGdV\dFJ87_F:FQFKLMSSKQD6F#8\G7,M.4d4/>4QM<^WWB<WDG?S1FXQ
F>J0G;S?+4dcW:NAAaJQgcSOe=gg+S2B(1JVd[=d.a8AD;N>NBb3MWR7RD^I^W42
dE-Q+fP+MX)<@@b:V6P3MIAHSQNMHd>9cOM#+H/^8G?CG_REC(TY/A4P1WNFc/>g
PIW;P#V)dO[(G5?_OBaeX-6F^DQ^3F3C#]8EJYfbgNVdRaWNDS9eO\I^P<A^\9FM
]PFd=(6<(Vb_>-3DcF1)<d[;4X?4&=3O0VNJ)3^K_OB]Qc]d3>UcbA,8H@K6c<OY
VdUF9Q9@@#FfV0]N&Y@9Sb26eDIbAeEUT9M;2^\d=2O6a(F:=Z?7&,M5O3ATbbDX
W4;fb4BH&>3DWMg>693HGCBC[,NeN@3P,(L&I3WA4/c[ZIVI#VK?DOZ,CQSAAe9X
f@ZXG_[3ATdIC_9)D;HAK0[P8[NH.6Gb+gT@+MZ26G>D&#GZa7JEW?IP0V4D,.(C
O+T<d[(R4)D1]@=7&(\Me.OJ_a18+^Sd24YUR<--U-]CZ+_[E[GV._YW3@[2GNEM
d[<PaVgP8X7\^#/;e928@C>P?/_A1&:gK<068f4+/DHX1XJT:8\,:BRJ7ga7266b
:I05XS5MY74f@5NQb(=ZB)bFC./+,T_2W&H</S7JI/ZdF5:gQ=_@C.9S>?[7_0Cd
S81N_FS_.3@^_M]A6?cQ@;U]Fe9feHS818c3]NMLILBOYf84G0;KFX(J?0e\Q<d,
Bc?><]9+&:&J+XG7b7X[S8Y,+_c;0=E_e8ZT@JS#CW,_H-ML=&)4R5^T#6DaHAXU
P6QgVW@XNPJG@X)=]Se:?=Y@TV<F2MddbKWD]R,]S)NQC1f)\2.[9Z[VQS\a^+eC
c&C4_;2IRY5[[OT(9B#e-GLUE:G#,J]#(,JC_T4,K:X0V0HO(7^_7DRQ1:NaNH\X
J?KSA<MBDN<];?:f64(9U\T9aR2B4^c:PVEZaZPM[4Q@)B1JTee-)P0KS8a#?\b8
-MZbYHGPYZESc:.64ZR#W2cM^O6A1@&6GJ;705b5D.,UMAYB,6<X__g)\7\OCg-U
Td)GB(3c166RO@K5Keaa;@.1BIB5^9GPM2)2#<aH?<[1;KP7E:,#@E\YMS><+XeL
+TAM=\CS[-;SAgCFOaEQ5O(@.YICbS2_):9a[[O-H_=(^c]_FGeJKVQ[<6AX_Kc?
6UWaBQ)c,19OU?_b3URW,cgbP[>+\F7#00Y;ERGM>+=bA&6WJ+c[O/JUeZX4=0&)
5I5g^H1GNdaY;T/CP<@L6^TPU-=19,7A\7G#DaSZcEW5]IePeA]-e?edG.QGPFgL
1P9G/&?P;DZFDPT46&A0TJ?=O)&:W5=V8bSBUd,9JcbHgXP]QcbdZcR(CC#)C]Nd
H(e:XIc)E7ADa(?-\RgG?ZOfWDJ6FLY<AA>W:O3?V?0bQQ;0M_eM=OEO0bMc-2[g
K;VSO?LB^J[>>.QEMJEHC1;@V/LMB^)=,0W\N42<=/,]c0S&-aaT2a,@S5X6LM#3
S^Q_0R330Ze##-#SVFKY2&/,&W<:E-3#F[\F-,JHCbN^^(c0W:&;73#&8;.H?YO<
E1.f-S+SLcAO@M.B=Q=80/K2CFQ)a6Y3<]<IQ.Y?YB8Ab#eGOCB_?(<&bVN&SgT6
WeQ\01_0BOB^EeS+c,/=M[=SK_?D3BI6R:-I?@TGR:Z:NT1@#;fN(DJdV8gBZ6P1
QE=9]@_.MSb\/&WY0,b7W/TZ:E)R_<[:1:]1_DOZc<NU?/K5#IOcRO0/bYVA/3TM
F9X)]9BT/.>feV?@42>U:bXaIgQ;GC:fFcf@\.LJe,A.:M=Ee],3F@V3INf\#eaa
GO^M^C=@RW&NgD]WK>R.-QYT[[G2,&N&e[I6_gLD@I;P];X213VT/CG[bQ2@9EC@
4^VNA+CHQaA,MPV9WM3CR=,b,;/&f<_+O+12FO8Wc5GLI[:D;D8T@7N\@0.EJbM>
]X)7N]?<K&e-LI2cE1=2_V^FPB[\S\\_:76=O,-4c&3;QH92^bfFd1_0T8a.&bNV
Pa(BbN;cJ8=B.aX\3ZJJ.XBZ0J2c7,+gfK&&PZa4Bc2D5^_Y?965dE6]dJKCLSP.
K:C6=9^-)PP-=G19E7>A_9&8,GT(=eb2KaJA(H>O(-DIP)47OV]0C\da9a,0@9/3
M)gJSTeK=Q:cf=Z0+&,<?APd(^+DVggZ0,>;6XHDZGAP9/QW#Sd7RZWAKAQFCS6[
WAa0(\9-1\9(aEMOc&LGZMSa<g\]YND8.)T3R(feA3IVKE;NLHIOXDSD=CJN.V55
OLXf3gVR@>T?A4f&DRPC4/V,]H3BG7I4>E5[TC2G,Zd<deVCE6:02J/7bbBU<C7M
GOb@Z\Ob?4DZ7XUH<Jf6@(#6\YII45#C^L6L-[ZZ)<7feZeL6IR2DbB,a1.GU7C-
1b-fD6T^4DN?,5495VK.R^SZ.aVO:&.?#<61-#4f9gA53);&/8Z4.7H=&=>G&S:e
55LdK-:Z=@J9U\DA;3]cBMTY)L+3cbSOOEH.fU6V.3(\+J1./(g>1586U3/^=g9Q
0W=?MRKXD#4Z]:FB9Z>g,;EF;CD:bB>KC>U<YecGO4=DJ^8)6WfFXN.8MbDWD.3b
fW+(:)Rc:Pc#I2W7gF>\#f]3O5[A(T6JGAD\4/P0J9KeSb@_P(.EWXVAF#Z>&UOZ
BZa^RU0W+?5T1QcK<^IHgcU<L5(<])LI0@)5Y[7O;Z5IcW5[K59QXg37QJ1E_QHT
;+P(7,/L=@[TJeU89eHXCLK=#FMZ3GL6E>]8UQ203;5;IYbBE/cS(#HQL)6#QGKW
ZA:C61BdQ9ZGd60EFdK@<5_V5gSK;e&bU.<AAgMQ8MFDO)>5FR2KD^W5Q#UM[8.E
@DR?-+9Ff5_-&4Q273A=JY1T=5)a[8P87?(SXd=4[86<:.T-eYG8O]XTK<EV5J1K
39Rg(4VcAfBfUbH@/?@FX<+?I2UD3-Nf(,aQJgQWWD^-X:\cH^S:B4,8cJQ#O7&@
5;d9^S&#U[=P_^_L29P5(X+HI76]OJgCOBcAH,C#b161dacF&Id&8Y0:bQ^c+H9B
V722_SFB-5I@C]CXfXR<TPQ>Id[P@O(eT38-O;c6R[g]Q\:(;I8=05.TCQGN/P>d
_2X6+a9QM>87-.(:CK50QR6ReE-N]L>.8V\[I4c<4MCAbeRJFfR6F9PD50[B,A7T
@(+3E)_MDd17AP.S6LX]@@.6?GeRR1:3UV\1J>#9eN2969^YD9JDNO&(2#2G-SdP
;NB\6;5(/.+#A62</.\1ddKcafF49C-D-^=^H;G.<N=HF=1?ID50;8,:RX:HHaSd
6gQG]Z:XC48ZE.=P1UAKQ[F;JYa0M,e#2ZYNMa1&5(P[d,a0g9CEe5b69&^\1K.f
_U7TJ,;M+5c3]UBX9<EU#.E&0,ceUA/X4-J<LSZV3=UaYW.Vb^T8,S\7H\15.F+G
-+\;<dP_IIS;48:-MEA6F\]P,>6Y&\9W.@<XaXZc>^b]:UL?K.U:\USV)=>@FH)\
BX+(5d0AS3M>d&f+?#b07/,XB(I+LVPY1\@.,^gg)fK7<;WHMGF87(3#Q=S91FFN
-XI;A;DQK(CEI,)D)4f+KCMUe,.[HJU03TEP32EYOK5\>Ga67UCfS(V1I&IA5#VK
bg-1QXUMRb7Cd_0A#B)Y9g7T=(TaKOE&3>aHV#)<7F_FVXLWCTFa[A8RI#B5Na:0
+&AJe8L[?5U7\,4K]Ha,P@X:3Z<.Q?3#geX8RWV[4f74B,RgME4O8F3],=+HWT#C
Wfd[(e/PSa^M>P#(T?#.3cN7CH0f-]AFcHAXR.:6=&GdYYbPA/P7,Ta\[KG1^f4\
;:BefK\6;^U&>=6M[4Dg=(H+Q:<^V-_a/_8W(^Bd@AU1Y0)2T,g@WBB?ZGfAWfB2
b?H?PQB,gT-+2?g4LB6-S43<W-@/2]C&8VC&HNDg)&LNY:__CHVX5I&?+WT?M_aG
OL544cfI9,PO)XTHR55FG,MU43Wbe=-,(>FNFYgM=dCdZR7.[[U)2I<eff:YA?A1
?U>QU-L\.F>8\e@X_eT;4E^IM7O/33I>+PVY]dJ\T&-XM^WfV]L@6ME.FQc]R1,5
5N4IMHNIUQA4G8M_1[5=A9(TT_]3Ddd9PJW0XBV)O-V9W?cD:)4E2MA2=J,@1a50
Q?3U;&]5c+d(3Q>;-P_[+(a18da)eQ)I3)GVRX3P<@#VDBTN#\BEP]Of.^A.A37Z
M[_]AR?g=2M9+++[ega)4A0UWdFA1/(ON/C.,G2NO723HNI#a2E2]<JOL56VQ)<7
Le5Z5OLQ)=Nd9/QP-Q#1a)HB<)((EOKIQO]R3e#Q?@H\(YTHgc9K/(a?CgfM6CM,
H<VU/4JJ5,[ef^.c^KS^6?W6S(JGOVZNYLEH7QL1KC2A.8=ZTRY83CV1b;f6cG&5
4RFbVd&9aDA553DVOAJHRdf>=\>Ke1eQ^EE_@0JN/T>X_KK1<A@\KKSbOUZg+PM[
;5@]^Y28-L/S1H@11H?[0#N@OdSJ6Ra#7Xg2.;43NB/GA[#Cc67H.:C[42aMNYV_
;AUAXGf55O[A&Qc+T.)IH#)bZZIO)=L(D#(S1b(9KS=X9Kd4fbJ3@5e3^-cG#2PL
@HfaR?)5H,XU/f[>V^eeBS&4#C;\dNB;c.F1FRE\,H9V?MDL?1D:.]#_PDM^Hf2=
P/(2<-EdGT=QH3FW#=\::20aa1S5/F<&.8DUB?3+VVe74J-JM(R,gORIY=V]E(=B
,)5_)YPb2L#076PK(\3PQg8+6HH:[\C-@T#a:/;J7>KH?bD,=X(TC[cYIA]A5C<R
/ZEe4d)_GM\7CPR)Z8)0N_#6/9f;B9MdE0P]<df1KP=Tacd.8UL.6CNF_@WV:6)Q
fV[>@+,VWG9c)1=4Ef8&-L.B9FD,0^cD.=:.4GIB4gK=cV=B\&F#;c/a<Ug=T+CY
_G0M_@CZ(g>Kc3-R6IP/D(f[:.-QOD/YPQSGN>X<ULFJ+@]f_V&gE6)ZW_MUD(+&
E\_87@/=K>49OOd0bgfQ.]D2.F>5-RW51_AeX;:;FA:VFXO/7TWYL.AI(5]Se\(8
2Ff(R;K.V4Rg4FWYF12HVYV)]8[@(]&U?T@:UTN>RBLP=3TMD@WA0,/:JW<;5;6F
T8:.ZfVO[TVU;/N>cR=;fd=-VLUCRW/(LZ,VVS@R6+,^c8b8\<@aO1c+WY>OY4Z@
#F,FN[eH2.@9PKJS).Y_BS9dO]V3+0SD3R-RI86((G8[B5:E@+A40d_3XH:&C2C<
U\SZ+aXL,&c<B@>6M#U=e+JMNFg;<H]@U&77:gL/0L8C30dZXa5GU/[Z-JIbPK:T
4@&:W@KS\AZSNGe?IBKK;PK2Gf3b@Ud;DCbRNGfeF<PZ(d\BP]+/<cR>5V\VY]&F
X1.Z_]TYI.CIA1^=\GaKCFD8+)c9f(:8@c14LO3>AL\DT7-Z]3V[4O(;@SUb>K4(
OS?D)Y,6[Uf5H2T2dKNBc^C[T[9cVZ0@c.gC+5IR2<P#8f[gLF.V.c^YG^56=?-[
b(OYXWJFZ>OH]G#QKDA0__.G#TF_UOY=+R(KV7>TV#,&eK@CEW>],a81:XT2I7:c
?+=]71S)+5,#+-e;4E:55UOT9D.4,KW#O(Qd>7<0)DcH]7S5-@Bf?><6M,T.V/0N
KM^Z-L@)O_5=3)[JDW5HfJIJG2)5gSg#deM4N:22Y>CY]DfFS0e0TA1a/X_OZ3ef
E=++<@99=R4_GS2bN.HN,]Q49[Y@Y0R/U4@-gAHPPJW-OAegAeI[27+T@ea)NJIg
E;D)8]TfS0TCZ8I7M,T:6Y[@UZATQO[A:6WEbd#:/8M#d;GT.gb?fD57LB])bI9J
:#7KNAX=^,;.#L?UZ]40XM)I&XN1.B#f<_413-U9fe]b(M.Q8OF9/@Je=C1>DP+T
,6>Q8AcJXBEA_,\X9fEMVO65_8+,Cb8DEI+K^f5.#1D+UFeI\MQ>U+14L950NKK_
/8;d.GYPH[U2W^Pd<V4+P]61AYMNda&+YE)&EfK;.[dRU=4PC[TMC8bdg8V@MI6d
CQ?c9K^I@]JQJ&c146fW1A[(RB#6C=R@K:5QT>B-g>#+bZU>#?TFL\5gX31BS.>&
)Pd<egHY>1Y]UB6EIbX\,<32>c8gCF^,]ITC_Y_RUaPW>ZZ#ZXbSY/FS#:5?<LR&
2C+P]1=b?P@FAUXQ].XQR1?U^RN3/T7>YPKL1_Z>>?C7MXaOIZ;..(N17UIa/,W&
9ZIVY3YP(f-BHG^G<6@327_U]4<bCD]fPQS-U3dcB6KMbT@JFLA&WdIAB///FP.<
#dQF))H]GQfHFZc_E=NRGa(1XZ;0AMS?X/5#7f#:)2JUO,Rf0Xa_]_dfCOggdF\8
3R?2UUEI]Tg(1g6@)ecVL>=4b5,W@+#=F9Hc,:C_?U#>HOc)cFN67]=bb)=g&IfS
(f;:+3a:[8M>TY^4J23H>0CO(bZQK)PcMX,4?A#4aeP\K,f:Z@fU5K)Xb_VGb=I?
cdE(ASM939/e\e5X0SfR#dL:2K.:YV8RDLG29a\=)cJ<Q+LK3AU58N[RMO-(bD^1
LCO,-[CA7gS?:YCf=XN.+;.<XBO@COW681>W(fY):bCUN8]EB\HG0EH_@.LQWf8L
26=eK\C9YK9Q:5OK6bIf,/LKIX:K.IQWE4NW3,>,d#@0;\T,Qf:,G[VEFX1+C;=5
fAbQH>a/B_YJPSBD&F#O/074)R2;<+22<.=b0).][4C[1Jb?IC_YT1/egBVBWA<#
YEZ^D+/0IPS?&cNOIUT;>W@QgER6BdcfAfA(SaP(QPLg\1@&a&)\R4E.-G>/0JH+
0NXDL5/#9(9_4I_FSS@+<D0)?X97b1Y8TABL=&Y,2(=DV\MQ)<,TP;865-Aa1V#W
KH=ZeZ-TGRJ6bEaeSUNA0/d[8&E-?UFdL295K-@=;M2(egU7-9G)aA.]H(<4I0_9
5S?8NX6#XK@H^/KGQacP-0ReMe=(eJAQN?&6\(I.4X;N7.5F4VgOICEC?+T7?<Of
W7C:W=@/9&b1OW_STI(Yb90Ge&/^K&L^8]J6E(IDRLI.Q&)9-45FTK?MDCU(V2N1
K19:]RT;@2Sb1)ZV>F?-7Mgc@LWgC/T_A(+145VdJ(bX8Rc_^V8MXB[L<85OL4RL
4/PZUB_=Z9=IJaUf2N668@S9KUSc-JP@KO/FGCb)SX-=]X+.#M.BG&N#C28;>/Hb
)2+Q;Uc;S^ZM6e).>1b<V#7]YRTe:VTCV_>YCMTF[YSJ6R1-:6f[SgS2_MF.VTUU
/b=HIKJ4N<S6[:PJaGf\BbeG0H5L?S,PZ(DB.#\A5NFZZZUQ3JS/GLUZP6CLOI>T
X^VPd)9>e^1dY(8,e@gQ-d7PLD)778G3J_V]<^2GBQB,=B42RUa5)Q9@6c7,=SP)
WCV>-ED?78E;=7fX_>WfD,(2H0U:<+25C@6OG=6JeNQCOPO817CG0H7AW(fMIGg-
.5KD6AOR3S\geU[X4EBX-2O\dQ+R:S4g[d(.9+8DAV2V>0Aa9/Z7KJI)P,F@I^K/
V,dHUQ70.Fb(A&-#]N(+WGDa4WP6AM;7V(V8f8<.G[F=0bd8^aFS;3.b2S5KgN@#
.K<Ib8.Z2.Q(SU4S;&JT&I_O9XLEL\(?@(QUV66/SO54^:1?&]MRQbU4C9SG:e,9
VNND_N;^cQ12=EaUAg96QA#]gMW\?J8/Q#OWH[@)gABXK[\G@c@<\T5S>@&R#C_W
IU_F]\#9BF)+6N1G8:c/]7ZO,#GB=&(CI^CL-<9ZN1GEKSCQ,6Y@7D3&+NFd.4VY
G0]KCNOQ+6VEgTW#dI3Jg/Y.0BdbR-.0g?;c4XWfQFTL+fUQ^SO@S,&..#>,af@I
R?/PbCQCQd>V3\K[:J3W(5N7J+I2//c\ET[FN<(UfBWE.8E71/P_.TO6P,IX_JVO
N-72=6UZYD47\QVcA@?-d1g1ESHK.H?=>YPYfBG-a5eVK@QA\c@GSYg5A^\^2V(O
KCdf]<TMSQ?+.;\;d(eG+)@PV@T-V,B:=QCXfQ,G@6V70_>]3aOe.(?abN>XO[gF
O+K;)[<9LT\2f?IY/.@\[geKeA9g.\8>Ca9TXLeY+Y#RR5O[2\NfG?0/MTUZE>SH
#:94/X+dACUT[TXBP#P-J-Z[4.R&V_,T;GP85Wf/][R>1TReaH[daLF^?5AWf)Rb
,16QNW>H:0,eV.gRVe;c&Y\)5Rf;-VAbL0P?I?:LWS?2F?T>7^<Nf0d_X0K3YUa8
RaF9L0O&<SXeWE438(D/HXCU7,NON1\U#G-)PAO0MH_.aaQAA@,>FI61,X:(Y5c5
f7<X#O4>=NJWO]b8QIEUF:\cVe(Pb?[b0e]U#)>O&.;HV9CUa=(R,ecEd9=?CLHN
Y&TP;I5QLDZ[=(5RZ&]M3?L:@#SUBQJ@?G-UC8aWVXI3Z06\B/Y?_P(,>,--4eE[
ZA((ZI:Y)D(4efKeTU-U@=c_O8=]__<H&I?SaPfC57H2^/2b[L#/KGZ)^MG..&bZ
CP2]KP\FHYS8DcH1[e:CF;HRaX;M7N92=RS[BCf642VeE)LZM,T-_cGb_V5,,LI1
f1;Kc)^T1eJ#T;)7Q)6d\B6M>@NW3M5M+4+O9R1b5VUUHBfJCCKP)c,P6Hc=Bb,_
7T.1_U<MKg36f:E(DPMfQ_N,IJeacHK(/E4>/@LU(0)S38f:2H^c^I9UJAJQAET[
cIRe(:\^I)X=PU7DRS=\Ng1_S6#^FTOIPJH4C27,+/(fL];5/d6((Kc9@-_,M(Z5
Head7^FMdRLOa;cbGYP1Gd@U84/+8NI@@4A8&(E7=gZZJSfWD-^91Q3#CB3G#TF+
7+V<8BX3K@=7P_M\D9c\MXDBICY:SQH029<+cNHVD0U3P5?P<2GDV82Z7eQ_<+bU
]MX-[W^[D1afRBODc0bWUJZ:g&a[V<A>9@&^5gR]LJIV/(4+.TLcZ\7J<TYcM18&
]AU^P+0Y1c_RFCY.O+g@QSBba(aBKRCYYD73-0CT/bV;E1X08>L4_5VT7a12Z)-]
S/VZB4<e8_0MP(-BOf[#8PR/20AIQKN7N[;^1\PC-/NK8c:E.H]7UBG]#8=aA@9V
Y:46ad+M-P-ZE777D0XO/b#7HIcLdQ3@J?IGTH:_HON,QSK-?UN#ZBd8F>V]EN@)
2.JT]L)B4I?&Qa[aO77V6+dEg.:R]LVP3H4CLF:7NDS[1B:4:IE?IU2Y?TPgbZZ.
[6<V9fJIKGM1MU8\\M11U&gJS[=W4NeK?cPC.L8IL86&Ub4I&cg9A9IW@0?9)X:S
Y&/b0d51Cg+9-LfFSW0(JBbLQCV_F^5<+0>c.__BLdg6;@?&R7FQ1c1UU7I_?6:e
K>N=6>;HGX(P6M#Y&dBKD1,+^FE7@.Z^AA+TN1L(Z6#RLWG.JG9_5T2J8J/-ECRI
YMH7/<_5/2UY#@V^@72@EEGL_?K;VOcB^Ua>X;cVF0L>HM16:.TKS85Y[/BBg=J[
G:,O6,[:4\<.d:U4W\C3>?#W.f8;H-A41LKEEUW\f>7@S1]4,&4@O9/UI-55O1PQ
gA>;Q1V3WUYA[.Y1DX[W@KLK@;(]GD+\7AJ<P)fb6-3GVOTWU,7=@+?(a]dFY\gQ
[1)/8PH3OA:I]<+TIC?SD<+03O@df<O-Q]RQSQgCYO\7N0C4;9LQI(W2F6U7HIR-
KcB_e^>KL(d7RX\[/dO-^L94A,@B^2CNO0+DEBP.6=A)L4VCIe&VB&(4bT48KWB_
9I?R2df.HCCT=_8@aEZF:bVQC:5?HN#I@MA;@9D#O-/)JeN[X\9N2:cb]&6;b0TI
dT61IIG0)=-&GKT6.<2TFXB3Z,>_+RB6WR,<2&9@;2<2Q0LODF_U^:7KX5Z1(:c3
:d#>J,NWA?ZC=#SB]\<,[KSbRF8f8MXb5CJ?4b@JU?WO9.CZ]=LOVI):4@O;=D()
TOZ64S@6E@\<b_+OY@Y.(9H8IO5<F(Zc&0.QV?P>eU<3d,.LXG72]^KdATT2Ab5M
UCOC:H\>_<._RL-ETAX\8^UNM2Q[KX\BHU<2Da;.T7-ZQ;V?_\LB[[c5VW7Uce52
-3]cW)JA@0?/+LX4:]c#I^MAgH893B_d/T_RAO\(+f=bR,48,5O(5@L;-G8VG7:V
4O_6I]1]d,0:685EHTg8Z.^E61#bF6g\U+0aCbZ_O6T54C2>&EW1=U@TSPa#@V8T
ZCG_EDU(1TT@:R@>?N.<BG>;F/,9M[A-88B<OHX(?-6@_2KN.V,d)?<K6PI/,CF&
SA0P@[?+cdA2>6R/9W\)g4O/[:,[G\KACA[:+7B31MB)<8L(Q#?gK&A3WfdCb8:2
C/:.dWVG35[2CS4+[?Ya[KPeMV??XgI5-gS&W\SR4[/R4<Z1LRNdFW6)TG7B):9f
UQ,O,>TU80EI6K.4T(eF?7&EZ.\d\CLGWOFU@(gEfRaZI@&0?P3fA=0a43gJATER
U)2baRNA2&bS@YLV-P\W_P+R=7fMg6N^D#+Y14OZ<]_M-#R=PJP/_<I+C3Jd2G#S
/F_90M3#>1)^S:ad06,=E:+22K>5Ke1X8Sd2Y=:.,5^,MQgT@Z1GZ9#TLc\6;9GQ
J\(,-bdH_SBU7#.0Q:F+#[=/+7>_Z=5/CPdP:1fD&R-Y,>]Z>#R7M6a77L6;W1&5
05EOM\#^<24XQ^[G/Ac<2gaDd/E[M3TIPPQO&E&2;UH2>d:.UZ8a2Q.(7&(H0aD_
5,&Z]b)BIfX+D,>5e>8/G#e#+>e984_PdF,a]=fL&Q[b7OO[2gBL#-b>a#Gb,1a)
YFZ1[MH\PJ=b^#>Le4)NHS?2ELf.6fbH1J5B8VF89#U0\RX95JG3WI:&dg-:>TK9
W0?8GEH1@O:]@[CbZQ&(7d#G@E\^>-;c):T1W_Ib7=&1XMTeS\OS09\EOc@AN;gS
C\J4#E?TWP02-EOE\f&NCH?FbAKHSZbJFZ(S;C90;(I^[/I9AODDHa/b/(D_D8.^
I(AE?IdX.K@H=de]\)Ac0a-43Aa<XFB,Z[;P.N:34Q+F:-K^@fA4J#[Da)J]6W<g
7SK_A=UZI;d1=/F@R[JJ914GYP7ZZC6f4S4F?^.Cd1c@Q^Yc\N?ef1W5M=8<a,NX
D2R@Qc>E2PZNgZCYYa&\\6F&P;g_YLKCNZYM[QaL07\fD&+?7[;A]1BYV5TD9TCF
T\TfHW>7L(4DY1AgL2f-4=.@O:ea,-=<)Uf^HXTM2:bNL7eF>#/6Z2<&)2@SKR)S
@,dd?78JeD3d&CS(Z0Z+H_\7/ZY_WSPB_Q:IWEA1H0JPPN>;1+d=fUT/V+#(SW?+
SWb.5g)fgN+K(cLfX\=8Rb?;B]_8dBSg#5e?]<>\]#&Bfe48;_(b7LfN8@CbHH[+
IDOJB91..=G\aP<1P@T1?1])7@SgU+B\9J5#:6GV_E&XO6B.-1R]_Y3>9/Q(7?3:
^cA(ZZF@b:?0R..#2GKHK8+3=f>FMH95XHJ,C<1IP;Jf<<C/-/)b=SZ^fNP#HH?C
dVNFWQA61fe+.4RF?SI8GL#,QO1TM.342eAW\U6dF_2ZD5W]=[2MZ53a=^?a>=4H
L=9-U^JAcG/c&@H5?23acHK,/W34/@+U-I]Sbd:g5LfKYS[JNQ5FADD-LP_1N/AF
??,NJ_T0>[Y3)?23S6QOM28&UYEdC1e__IC0;F+JN8HC[47RJFc\I/A8a#;C8D(7
H-&7IPT^7NbK=-;Na=f[YD]g;26\)OgL+HTE\-DEa4;QFF4UWgE:;cgN\Qe/^47d
99P&;HG)dN,[CA38(8.D_+GU5M&HgP-SM[_.FRYASeTfT&^)IYH]W);5([2f/4NL
PeGETa+,;6WHV@@G=RV#=G56)ZYQ^C8aO<QWJ?d,X&8M;46YN+_HN;gKGC9OQgdX
]T+6W;RK&.(3D28S7.Y=8]BF#=^2UGa0@&bN2]Y,7@/KCM<>^#0PA]T1@?G;.0\P
Y@,>L=(cC:5+PTH#Se_M-_3#7FZH25RPgHZNT3JH<[@P_6DTF#<g7cX[[3A4dH64
)XRWIeIgS#8W\-N>WFJ]P2?f8^6]KHf@>OT\d8IE=?D^;a[(GD\e3dXS2ZWf^.PX
R\J&CA)TE(eXV=[]aR(=Y[CE8eB+38:c+0?;\U,,:2ZH&QK_R24U7#,ZTe+N7WVV
9c.E,ES4<aHZa@?;/C[]+]Z[>GSE-N=F)-N<V,)9U,.O-dDHZfbU6]Vb?SHV^dXQ
^?Lcc)Q89^4X6ZR1<74.0J]@_9O;Q?XICN[:ST]aA1RVf.Xa-;VP/EbdCB7S06?L
KcYUW?BLWQG79O^e4fd7CT<XF1f-GR_EA0;2=3WKf9aW>7FfCL#Q&)GaA/>RDE^;
7.>8-Z6e[6X&]IO/\W1&gLWP>3)T6?@W4YR;dS]L->fZ=3ZJZBIfA[8#gR5FZ1L0
8f.&NI>&E@BE=WS[U_,A0LcCBIg&3b(8a7Q)^S(5=;gY?IN,;Xc#aN8Hd.@d1KUd
(V\X&NR)))Cg9I#HX-3YGCa5aF:+:]CL.bE&#-@5gG?W[TII(3UT-QOIB&dGUDS0
L.Z#d\@6KBA9f77F1Q]?CP;W/?PPB0NV>&D[DT(3)Y<,D,=(_cRY<LY)?]OYZ@S]
P&>W;gZ9U7Y:+^eIG=+]@DL>Wad&bXIH<WC&c94-EN/Da.FH=;9V.0^9a.@bU;(/
)^>G#8:VL(Q5697VbASJ-?c\+g,c3aZO#]K6W2Hb^I<V&WH8<6KC0[2..D(;@_gF
\@=^0\LeWbLfWKU[,JQWcYJ1W3MH^GYXL9IEVLU+)BYSJIg7FP@7)66ESd@<-._^
_,Q8P<75fgDVBA-?A5D3:,<SOXf#J)^2K.,?FIT;3O/WNAA391-@,^U?6E[3@A0[
P1)^QC3-,BJP?,DI;Da2S7>WE9fU;,G-[6()K@TdDT1/C2@6FWb064WNgJ1#6E.b
B3A.gSU0/2_#Ud.+Z<2TCUbE5RUW-bGH3[S@b<_\;5(c0JWLI5?83^TNb3HF^b/N
2_8D9I^QDBCbOQ+0K=7b6MY>Fa1?-S=1><=I,:.a&bKg9URdH&]D1Z:UK-]T;>G<
<e.aLG8N49UfY-<Pb<[e5GO/5VV>WNe7UHaM5K/(S0LQ>f<W0T8Ge>G_=Se]b?9C
-.=?:)K@-@1?@ZcYNb_CV]M7UE@K8GPDCC6G)5QX3LEM5-UC>NU]8bfZK@+b7P5R
5;&)_[9+?PAdeGW0QV\d_E12Z&=Z8DAOR<Re5HgA&9aBb(JJ[KfK8\9\e)0W(d=\
\-(0<WJ9#gO-c0LB@9Q3,Lg)65,(BZKbB<9.MF][+04HBOY,B##d/<Vd+A@O7#G+
XFCW2FX&Y0]?CI#;IDCH4[EVcggTZL2EWA+VG@8X6E^<[&Pd9)IQ;UO+MTe.O;Yf
,99WB7RK89WAY]QY-BE1B?H0g(eA)^7X9Y;Y><G43<\FQ3b5aP/_H3[&)-U7N>+R
X1b[AULPD2^H>CD+e)/=>+D-G;3IR?-7R+(D.9-MU3\5PG_+N-S3QC3e>&Q9F/.)
+MT&T&@#TLQ_O@84eM/_2ZI=_d[&ND442=Re=B.aCQgW;9V^F-Ha_eV.a+;OGO+V
g)fO?MR?0(,6e)Zc:YI&PI.[UC0]U;O;D]4;O.A3S7AGVTO2@43)Ib+WEP(^g-Q:
9BfESS:^/AT@RfSc2:N;/BAaa-.BGPD@d>H4dNQZ,f@4d^+A\IH1WEdVNc76]_?4
,D]X0=9b=B1R-fA^CX/PB#.e?M]U_fZ0He9Ic&V2^c1AWB#3,_83[TK:,N\N>aCW
@MSfHf-aEE:RX7Zga=bKWVc_KP,7g4A24d+b5G?JRK6aNJW=?Oe[^I#dVBQ/2:]T
Yf]._]J,?e<\Y&:QVc:gg5EP[XH.I,&D+XN^UVJG>7MY(c_(5f(;I)B>a&(NH^,2
;JK&>+@M],GP3?EW.dV7S?Z;G)1_46;^:;?S9Pa8Y;f7\d5cc\;XdD;)bS=9P;0O
#&<Q-JaH-,_@T<.9SIfbCU]WQ7f84)5IgN4FJ;gVVcM=F#BCLTG[ccE/#RP/E8Qe
>B(5-)BAH4M-g/[17X[(4CD19#9_2Q--1)>deZCM4U931+4MA:TY.8[f]I7J^,LB
,R3f1+fBY:-/ZLYc^0IOD34(CA^\A&eR9d=fTNF?V6OF7+M-<PT2MDAVBMBbXf,e
3HO?M@G#>CI^76\AU916T?1?JUeK-B_/cY2XA)V?O=/274KO3-?D#<:URWGbY+5:
S1eL80/L]8?-TTf_2?c#G6Xb&+2)UfbJ9H10,G<Lg4Ebf;K/aD^=RabaNGS-#IJU
8c^43KaJHU_BW2NY\M?1RM/\QDJaf/3MUK?f]Q9PNZDJDDOTcDN1]7=,9Uf,\)YL
P)LOA/Y3F3QP,=^Ab92RfHAbPJM<7[J/6@6J=1)A=NAAP:TQWC2\[7GBQ@.<;P,7
gLC2cJ)0X6bGK]]@@_EQcS[(a+]Fdff<JPE]I&SN,e[NJ(?7KIJ1b/<Ld?AXR&S,
XYL#K.MZ1])G1BZM^(R39URLdgHbgb8EMTR6A:2S<85Ya&;_^B=R7O[:SN)+MG,_
DQfc^>6Ze,QYfCe=G5Ub3UbYD9:TX0aS/LR)7CdC2/cX.^Bg3DPAKK)EB(@G6e_\
2BPfDE>(@#IS]0Z)a#dC7?Q;/D[bX92Va+@;3bN7NT2DZH_FaIH+-C.QT^P+DMH5
::C2aK<e<?-#S;A+N.F9,Af]Ba-1W>3dUAfLYPNI?D^;SccfG+AMY5@Z>0NBM7dD
Wed[R=Dg977OYJ:T7YUHZC<AP++Yf0LR6]Nf@^aR(Y?>ZX>#]ENfHWe9QYLA+KM3
9RBR)_AB8X<<\DK3MPeZ^>F@V0fDdNIM,f3Bc(MG4J0J2eK#DgU-ZQ(eT76^RgG[
=a/21D,#H5[5#E4\(]g7[NQO-\BLRa@U7b_JN:ZT;F>,YE]_b_CaJg<>:A??LA[O
]3Mf0OdbXIEG7edbMDG.A]DRRZ<a+:_RgM=@+R8SJ<K)eS2b)[]b[<Z).Q_-6R7f
WgK;;Z>Ze\UB)gVbC0f^;IU^K68.d9dgD:G.9,S2<7\HeK^SaGffZ:T.M@38)O2b
WDaa>HHDUEe7>\aL27-+Q#Y9_GP4d\A?ASOOI8,<>@-8T4OaT-g7V2=IZd62.(Q+
3G=E/:@+^]9GcS,LSY#DfD=SZI>gg50e1HOe7,66TCJ&W?=PY.&=GP/C(3cQNL0+
gE=/XR332Q:4_b.7)9&#Z54Xg3ZAU_ASDg[<4UC+AH20;M#5M]QT631^ggL-bY52
A\.gfJOORDZ@48a>:ggU\D[^1cEOEJg]:G-Q^aZN<<B)[00]d5_P(D4a2K(+1YdS
eMD5(?b^0//Nc2;1gYC??/f;_<)TI1]<ZX_1eH/7HQO;:T.?\#(;SVP@VJ#PgIKa
Yc?2)AE>C)3?c\f9dLVVVdcDXEZZSbO\bRY\RL]d,,1fGH\N]<((1)AX1@>NKW,&
+\]c7:52KKF/+L:81F]U&_A5F:Q#MI1M/>Q/Q4(\\5^].JOL-(_2,E\UL\ST-4N-
cMdRKaGP3CT0_@:gS\)VSdB/a<8]aCAOXU4E_(:=Q#=aE62a3EU>IJ:1DPfbg_,L
T;-a62R\_-#[#b3+)-LGU^ZIQ:.W]A2fF(/<Pad8#BS/29?cQ]=3FIMc3<5e>:eE
F]dZB:g04f5CB0E2@8#M1/BW#-30.4R_N.BY8P6DeW2T0C^KG8A.]e.^L9K_O<_I
YU5W?D=^?1CD6K++A_FL37/([XQd<Y4Z(f/B]a>W2MMKaZ/I7;:YY^1@23GF&7A[
3=:XNcTABA64/W<Kd^dCT=Af9L[.8HgKaeIM:D7-R:WJ\Y98Y2U:4<+L5fQVVbU,
PVDLDa0K=g]\F(Y,6;C2@H=ERX>D/89XJP2OT#/<E#S#GVT+g0E<g=7IR,M@-D/3
FE,gP&f@^,:UPaP<bE(1GUYV9NNYF(KUaN.e^29(1&[:FPb86)P7bI3:a7:&@,0,
?,?4R46W\+:7c2NbU\3#<@EQ@eR2:<-90LHggOe6=b,\=-6P8WS>M9PBFZ4H<AA4
2=Ga)9,6T>9IcZU<1(0@0a3M]XP\5W\:3OM(cb[S41[]P92S^-8>O+8KZc<@DJ;T
E&H,bbF8g)RR[03:8He=YL<6N,(KMJ_WZ>>fC.CZ\<QAC/;BL<UT3C)JKcB_SNSD
<B5M9_==C>LQEM(K7\NEcM;_0-N(S6SSf.aP+I+bT<ObH^bcS-&980XVB3V;4_.V
#@\T&@b9\O]+UFA<6<O/NEFQgaf#DK)Z\@I=<1;/.T>7OI8LQZ@;#9ZCg/#X5)EL
.UU=];OT>;=M18A:P0(d<aB=f2S+W=@<Y=Sf1IfU/D2E&TFS]2X;H[BCVK,]g()R
F=:)NG-70X7WM7A@A0@\S&JR?,aY9]\bMS[WXQZ=_L3;#,KNUf3Qg3>MfT0Z26g;
\/a#PNaD;WBA-DB:6c8c.S/[8?I3Q_]OBYd-9dD#4TaF0:T)d:]WF@.6_Z&AS6C4
,_2Z/_\R<6;Y\7g_/UOCcd#.5(O]d36=&EM[g<77=U<[f7XIbX<4MI+f/IBRKX1T
X0K?=OT]aO2LMD&)14@M5g@6J--b6GYZbWWDV/Td0];a&8;O,2V<9EX>;^?;?:YE
[eQ_TbW/\UZDNL5-.KGM8<>S?-DcX<]aTWdB]40?bZ_3[8][U4ER_NO12g2F#@]F
WZ&YH(>+fUIR<?1_HSZ]F@Ad8\7_>C-A;7-bbJD[0Q0FcN4#eb9;OTcQ4f_FLe;c
:SZ9N5/HQ<?@+Za7,+WHG5:,)M5P9]B5?JL)f1aY5TE:_-(bV(:E&H+R7_.7:+d(
#2?(Qa3PfS6QB\(/OA(4=7=Ma#X/;)3VZG;]db5cIB(6&J_g22(<3P:D3U^LP1J-
X<Qb@X783D)X#W(54BIea4+0=I/+S<&;g;XEKZ?(\-b]EZ2?HeSQIFN=bVKFCB/K
2\/,=4&I24)<B>I]VIV:]OP_&1K;#9CeW17A5V?,8EL:R4>Me.D,EFeO>7K1I-JX
=>-12Q.F7ff;W(c5_5G9P=A643WDG^J<_I__^(J6=R_5^&U4Y0XfS/&1UK:e(?0Z
K&Vc>c,J=f52GBXA7efU[=QfFX;(3D>0gI.dWK9&P#WAYZY0,I7#+\LDR6<bTTQ6
J0PK^Z9RHA9IM54C(Q4.>7KK3]=&QYgK8X]QFF@a@G7W[KHUe9WUf07<)Q/@BX?R
)>@a[N;+0P8;d0<+dbCb&[N&4e_.;AVdVI])EJ=1:0f&9P0I94.Bg=f-?_:)XbB9
C<Z[F_&.<YJOZ-\Hdec:P:A\>1\G@(28Y^EfSKdR6.C5HfV\45TV-=)WDP]EZ+]-
>P?RVbNb5EAE_4]LX4LBC3Qd\/SBdON1D?.;VX/D8DO6/<f0/54UWK6?;8/IX-/;
NP]9U8KQTM.?GSWM@7FMX<3)adII7RYg-<<(e#1UadT#=3/HOcNKVPM,@UN=c0[<
J.&M@A\?38_>G[Ac-+E&,7-SAW#Z3N;9CD,PVCM4I83:F#<AF[BEgK?D7&d@0&(=
ZcUE>J8&>=2<+Q@5@4G7O1>gd4M.XZ(V33=IL[d>M^UW[TS96ESVWJ@A9-.c=7#0
?4?P#5eRK8Q6&(GR);78W]H1]KdFY1M38eQDYC(D\b@:VUKECYS?RLgc;^[[=Q^G
L.626)Y;fUTEcaDHcTXG5RKX6C>\NX_[O9;8a+:eH.#Ie,>MZaYJd/;]X_VF2.(9
GFf5XVJS7-,E<fUCQ/aJZ=L3+DE;WZf2(FD1L7NFQ4D8OZ[KQgMD[SOB&Vgg(P+c
(2.E6@Fce[IDJ>E6GB9OeGRb>-7I&)H7FJfI0]TUKM7:H?HUI?UHMUaMEHbI\gX8
(NKNe?&:fJR7(WRIC9;EeH\c&g#7f4NfOgD+,YWd)XQ?\PI3g.1)30DdFd&^2XYX
\X-E;9_O)dA=T/T)Y6HM>6Z]J@-/^Jc&C&6WMCcLEBa]cd.<QS[(CH8edZBRb;1K
M++c.LOT0=/-a1+b<4gYY9g^-V?.?g0VDcUC\;U;_M^NUOLN[VL3-_0N5_XF+0EI
KA2J?GHS[aC+I^6@71K/b-,HB<3V94JPAN?[H^]aS(IMICJ;g=1=L]@J+UJ=H/CB
9M_MQ1C_7\MS-=)f8RL?-d6eYf8-;HAJF_L8I,QD4LH8dIKH9)+_d::Sce;J6SY_
g>[T6^/(@T:S<WT1gVER6Q34Pe7-fg-9G42EGgH#D/.9C4)&+HTUTX@B5A-J-D2E
O[7=BZXNH@,8/2?X-N8=XTGSc2c\CO+b_>f<fX@F_M-_(,:O\gLf@F+_U09.QI(#
=1PSAgL9:7&..OCL33]d+K/A4_KDf]:8S5.CI:@GYHAO@=GZAO4H;JE9\)QaO-6?
/-^I1^<GN14Ja>3F;;[1,&BO5?</#J:L(6NBR3A=8-\AD@-0Z:G(0S)bHc(SVKeG
g-1@5+5K)I^[a#^7\NLD&3VWBb:R/+JX64HHI^Q>c-WG9DQ\/A;(@e<[5C>GfM7B
VT:#R3WB8SWJDWZD+E]gJ^(eBb4S6[Bb/.)N7((Q:Q07ceC0??2A#@CTH\BCSdWF
M]Ib8):)7KZBaY@JM<\Q61VX)?fO_BWH2Y0^O=6,e29-Yb/GUI=3MQ,X,KF=C#2A
d&=4AO.Cc>.?;g8.EDCBMLG\(U;^AIWfd^=?SQ/_L4e-R:J+XI<+(1[aONNI:>[4
.D(;)^F6_7gC+_7g2aJZ(U8>N/LX4bR7M4WO]]X^YXIf[dOVN[H9@)QCFX_W\Tc5
0^0_YR15YH<LP,0IS[CK4ed6/13d8\c&d__Y0Vf-O\WPdD4I2.SF6_RUCIL+dFF?
KFe=PVa=_IUAE(+e\C[UM9?P&Z<VgP1W2D^94:,,FZ9)65.b&30=E?S(X>93S\ZZ
]IV7BRGGW?<^R2F#4Pa^f:f>MbaN9RcZ>c):d-;?0)YYgGAF-&P5Z,af(ZfTe#HX
b3TMNHbH_SR_BQf,f;NIDD^C=EZI82[&gD-P^]UVIY.fZ4F?;GLW,L<[bf(\@@WC
+Df&\HEDHDHK[.IX4Q8:dPC?<[,]X4]Bb?W(W/+-b9C7:EY;ONLMB6QNa=FD9LS&
dWAPGNKE,>],&4\SD[=#83&T?XZa+f0=A?5U/6bC&ZD;PO3U/HUfd#0#OLg?E,_D
b@dge>=Ma94G7&7LN,g##bIH_[+7Ie\EXTg(U[+I#-9fVTTf[J(4X;N.O^VMRJJ=
f>BD<9I[[C-Eg\bWXF][E3<HKdC)LP&ZOMLc=8+C98^P_]JdG,9JJ^JB?LNDIVa2
FWQ+cfCA,;RLJU.0/3Dc)g[0V8RZ=AB6#,c0/;=++SSG)VFSQT&DNM_3d3Z^2g5N
HI/Z;5ZHK7bFVAV2a6?JGMR1B]UMJLG8eA1Y)I^02e?DA-/)3ZM>c1;QK3<JNA3c
K/&d@[)bZOJ;+71M4aSX).ZWc0;Z+>1M^]Geb+Wb/I17#86EFcd]2gQ?A[Le1\V]
02J\4]cc[/7R=HgcCU8@;(eU>QCS?;ORRL<aSTH2g0J-/R->[?:[#3QIZfY/;LRJ
ZLKCJ??:B-(<dG<5-)=NaM9gP)^EDaaf5M^3]89cKCgT5ZYYAG?00_888[G=SU2\
.9/^f394/P8g@B&0>RA<8&&PVD4_2fdLeLXF_<SVG##)N]+=@.[E?98H?>d4HM3?
F:7YS,;3e(>>_GCMTU0S0AGM;TdD_8Vc0@Ng-:Q8gOQE_NY&GE1S?T.a2g;6Z/Sd
bV7.2L5(PB=0=6Ea_^]4HT0feLQB6=KK&#(01LZB72a]4>:=,a:Y9b7_KJB7_TH:
Uc:\IeBAQQ6WcGPa_:?I<XN>IST,Z5)TdceVRO+C7e7&d7)g3@>&gTB6-H60.B,@
\9.I<\Q9a\2Rd^+C,D-KEH,WeBbIb^WIId_)9aDe]W&7b),.Fd#RF<^&I8UDHX[I
T4J/4Y1CDC3J4gC)N+dS<5O]JXCE=UIP:CCJOCdf[DOa;25E4[\Nd#Z.TWE-:](e
Tc/(6MNS,KP)HIINe[<6_,?\b)B,AW^?^16]VN=^;B<<5F;X94&=6;:=30+&+0Hf
?K4.-g;Gef_cQg5A,(1bg^B_G<QAT2;J?O-0d/X^7=<_YO;B<0.a8AD.:BD40\c]
d=\3=eBXabPEW(fB1FAR+@1MW7#M?=#NU2Ad(P=Fd@1OD//LG&?DL0;4I?5#b?NM
273@9UgWZLM8TCO635QGDW@aSY3DE#]9CG1US]G:D,3Y)SO<_G<PP4Qb4&GRS/D.
ba\FP_dT&Yb13M\fQ5JL^J5CR+K;0bd:67XR@H\ROL-1JabT5[c6;ge;#NF>d(04
4.Z&:FYdd)gQ\G))V^;>^YU+?,[a_/2OCF^__-UbTYKX>+67_+WO.AO32aa.F0D/
IP8B0(#BDP/T1<29gL5XEW>Md_,cc/#K\]S?&&f1YGHBY:eLe,;G<85feg+\P:/U
0_,NEXd+]VKKgf@SJC]VU)R7[-AM0b/f2GB)#bE7=F&XQ\-UB+X1,\&V+ZZT^_^O
#7.)H_g7F95:ON=BN445FeU&ac30bQGBMCg4@PV#e4OR8eA#VFBT<\HZJ06_1g:A
Jg&&a#_RUFRDDI\PX+2PD_21;8-HZR2)J#.VZ7[Ef-.MJ0BOdW1=P)b#AV;e/ERT
Ge/c6QB8U3/#>W(?-8QMN<RKS7QL7D]+XA6gS5d_UO@U2?>g#G39.B85Q:CW?,L-
2);DPL3#OdS&B62V6DFEKTGU<Q@a^U[3=)IW^&8=-.H&LM4&A,fd7&.F6?#WB/)A
0,Wf-]:N1V2[1]Z-AaN#a7efbb7Hc9VQBQK;O3S03LY\_cOeEgU8?YKPT;G6Q(2b
GI:aVNFaQ=<I9dG65(f5ZC)(e56b?5AQFa40K(&;FJWL#I0I[CO2e^+GW3)RGg7#
9W@4B?4UG7eG)_<R/FY:IE7.&3?6P2d:=^S0#9MFQUP]0H7a=+0eI<,+GK9<;KOG
/>,7<Zb7&g?@QCRH,/@>ING,fBDLAESJ3E6CR]>\C4NcEIWT3SV0d\9<0J8gNSF,
3<:Hg@(LSH4WT^2##V#eXbWaJb3?-cW,\ZQf/NBWL#_GB^BK^_>(/@F9B\Ue^=d/
e>W/=cBdSg)]f?HXLS#H&HaU]?[U7RK:Y;G)K50<,IT&a2g>.X@&W&ZGE>4b-3V^
,gBC_JRE9>[V3?A[TCZc[JO0WM0f2U[]HIbD38dV;GP?X0\NS;bWEb@/U]<Le8><
W6-FI6=I4/dB-[[F>Z@gT;gDB71PYdWVa5Zc?;.WacVa)N+>4BU^:dM)2<J]NG<Z
CV;13_EGf.)>XD0FJGe0Y/8GI9aXTA:FV@<+5GV+K)b?Y3GJB+;A^+&BDcK0Cd-E
RUAL8X^3B-#+3-2[G.P0MOC)KfZ=ABH]54bYg1@XUF1NR12F0<gXO1@<\PXK3Eb]
IEb77A=Tb2&\?11?LfR3K4)CXCFAL2MOF5SLFP?:AbU\R2(QEd;NJZ9=AA0OP&ZX
N=?,aGacZ_@c&2>:(L,1/Z5]I;_RXG^^-B3P:=^eY3@R)^?>[b5geg1,U9GEP/^&
WGc04<546ZGT(QD(HKAV>aBT&_-W8_CN-3YLC]016E]I+BcB6ET]O12K(Q-X[1V6
g&RU>0J+=J2ef2K9[69aZC-J.<+\82?6,OP^dLe]4X29+4(bVQ,Z<D\Y17L/I5L6
^I7&aU2,157Rf::P(:E.Aa79/7VVK5.9<?FWc](@XN:-;^T0:#AdZ8c(S]/2]?Ce
QFEOabFK/8\^1f/BcgW([I;&R.;[X[fC^<8?R^_N8,O8e?KgXYL&YSLfVEAJ(PCM
1S8G6cK<f]8Ge?H+O.\d#A<^#FD]b9TWC)HgX,+XQ8@/@-#PPFPE3_\:X1X@a>TM
F1\A#J2^9NT7.1]VdaZQ[GG1_4]#1WTfd;&b-WXLBZ68TUP)@bJ+KL#(\Hc\PZNd
2JGf;WWPLDWW+D;^@D57@HJQ=>O[B;O7ZfAdL39a^8fT-]gQ@TGd./BcJAN.>>W0
&?X:Pc/0(YHM1gP7c;f8(E31+HY,V-C[29B?VQ=H_\Q6YWeYbC[SA>]Q6T^c&^;f
Sed(:WNI@&E85/FFO/<=[_^EAeASC)I:Wb-8+M#eWEZH(DdK7E]d4Xg;b2HeXT+2
_&TS94=^7?=7&8:&\4[#^bW4HZ4P)=cUE;KbYTH0C0V9AMM.__^K6c2NK^[JZcQ(
MO5T)L[8[_:f?\H.V-RG),Ma65f&ac_MAI?#A2UaI#@f8Y]b+cER/?#^-;fbFeYV
@eB@EAO@eF35RcKGZM)cJ_Ob2d1G=1e#P#J]f4:=?ReV5VZ,923N[[LF4-#BI,)P
,V-@?<8O8^gU88N?aCeVCH4W,CQFOO:\a,8cNHS31Y)F(O>1J0)P5TS&gMT:TLSA
5f_:HQ1V,H7Z;1fCB^;deGe3;8V/Y[=.MS+.TTeTfI:=5<C[J9fARV4(Q<-AACXQ
;YU4TKYED3L;;40H:PC[Ac./UcfW_FK-<D39K[EIZT<M<;)eY3&\25RbOPfcaaWR
,.1-OTaGQ1H,>WT?I2dPf<T.R:>&SfE(VIUUUI6JSL7>4;ND47UEJJ_(&U<QM42M
fb(4ZQXF1;WXUPBcB2fG;T0)N]ZZDGNe^#cF7U[GT&);0O41LVg]4:@I)TNNMC<E
aTCB#^FK/-NWP<35ARJKAd0,/,@cFM<NVDW;2<97Ug3=b5M@=gFAgc5V75D)UEDJ
K/<KHCE0T.+eb-W)A:(g7@G@0/I\,(48XcBJ?9).Ig7=IK\@cSKN>7_=9V^DbWB5
(bT@&RU96fC;&dWT-J,,LWUbgKRbZQ7ES=;fQGYN?<,QRWYU3G\.[Z)Be(OL@7J/
a4>@APc:T)/JGR+P<J:_a(O3,Nd;>6>Z4d.7SF1\Y>4CITUC@UZd:GYJHY\F:fA]
#T^2\/7LAgeeR98E;B@P8?T+ddVXAfU^E?ZAP_4eD,N[:I&2#4X\^@<T8-:E].&.
K<=BW[_>Q3>JaWPb\U4_?)E-OG1TdgZ:[MT9]9@7R1>2N<@HISUadCW/A)2&BJQb
,-KR+O4P()5JP+\4Y00SGgJeR2-\F/GMKK6Cg_D&,XfM2<SW&AM8dYF2f_6@/X:C
:AgJSTD;YGDf=@f;PGQ7gBNGQ2U<Q[CDAVdJK+IgA3bI<^)Q)a<XM+OJN/eGZWeJ
=83HKKNMSY:RD?Dge74BMG&UcVQR)V,9;:4L#fU892>W5&O_c4G/9E_C+4>8^Y;)
?,+\IB/@YB5?d8Qa)ZFEV^a30[^42V(T(O,W&b)-?C?Db(AM+F=b4,8NX>](L\AQ
?+[Se_3T64DLO8(0;(;FVSK9B85<XA1RXEZH.>ZJ8^=3:WAB#C0Og5E8_S;E(>Y>
=DRWH\K(_QQZI&gRdM(RMS1;I,E.9gF#T4L5c?&[):O1c(G1L_NHNXY<Mc4?g:=)
]Z6=^IKVTBW&V0K5Q35Wb3OTT]g[^I=c\,8,g=.bDS2E[EcA4B#;-WG.5>f12AYH
#g<.,gVd-40g,-Z?MgG,RIQf.9[(FgGc,NJ41N2U@cF#d&KeI:eb=@P:=?92&>JB
\f^CBXTR^+F@5Z93ULXgV&0_B@/LFGf79R[OA:\;aR?Y6?AONTI4BA6J>aDPb=I[
;IVKdg5#YZNg\ZWO7.CbBg]Z0P0.AJ92/C]VUU=:=:ZR366J&Jg4.[W)W8OJ4Q(V
I+5C\>V]I:DZae#&O#NYL@fED;[1CYCPbd]0;KIH@HX9[4#4KgO:[.MI.RDbR>79
UP+Q,VT[c>Z9#^4/]-=Ge^2WXZdH7DQ?<A9b@ZBAbbM]Q.\)gLO=J0:AfZ2HD[&L
0X\YZ&FIQOQ]PfU7?+#Q(I.fN.4IWCA6a>:V;NQ)KC(Y^9DcgfH^E]B2g;Wa>K>R
fff7O_aJ#(DaYOU6UY,XLQIRc)8B:#ba(&LEDOXITF:T&aKbG#aUNfDL,60aB/D0
V.gX\]7^9(e//9cM<>U33V\V+OE/[Y0\GC#SKQ]9\cB-4W3SeRI29Z;&fO>OK/)M
&f/D\&^KQ=QfeJ2d1B\dg?VL8K/D-(Y(aFLfg2IF18M15;HTRF+X^1>^g74b2V+Q
F5Jd8ce_^&)^;<@E0+SA9Q,H7Y8;cN\9;gWA=e#<V]\WbE3:D?_O@S#G,M#c0,0W
]\>8<>bQ49H@fdH\SD\FP3+HUYH?1?Z,,=(BWZ(U3A-f0RL/M=T[SASb=;F-8F36
#,EZdcD&;0D]SJK\3#?G199/g52=:KdINPV:\O7AEF4g5VDA@45??-[)XVV_WC^(
48@G0R-J@-CC&V&4,agG^8[a[aJ2gFeU:JJ<OUNI&f0/YFf=7DW&UTb:9>S5RC;=
THR.KW7]eD]K]RT2+H-5F>H=4=B#BUSI>HZbB#O7&e=1f6a9]&_dHCJ#PE><E\EC
+YS1/S&efTYS?5-RRY&F^2OE02.G4N7aV?dAU4+B+4P+:@WL34e8-8UVH<Qcf&4:
7]BT^G_S&L,8+9BTL-(IPc^9==@W,9VLTG=,DEAV20N,CMOE^)JTRB,PB(\4@D?#
<]Lc;9<4.7Ad^FDUB;_\^6\I.F3Q-C,CH2SW>TJJ2C<WTNIaTPEY5RM.AF=0ZO4#
WD@..g_9Y+K.3Q62:1PLXI6Wc7(.aN9gbCdUV@X6KU-050JV>T@?+&UMc@5YYE+J
db)8D,QY(O0,[]?5#/SCX.:cH7N&#.T=cJ&Sb#_\)a9@?K]GTYe>5NVM?:YDZ0;\
]IB?4FP0JU@(:R,?Nd-f;V3\-;f86/:^0B+5N=#b,KK_FR[C2L:\@USKJ9=7.;Sa
.d&Y2.195ESH3KV/^9<AbaN2S+1\ZOE4M>dFJ&\P,&=d#UDU:/_RJaS+T/TR@B:P
4_-?W^PabZSC0\2J1C1@<5NUC_=Z][KS#VP4Q_4<WZ4EQ/Z@M3FY(M5[YGJO/K0-
T>dCQ9ObdNY.b/ZW[#N&4Y<W<?^B;K\28c3I.M2Z.ZPMMA9@8VM1B.RL0B.EWXMG
YHBQ])OE9NZVOZD(GW4=>./67TV3EL\4B:@G.L09.MKR1A6KI5bRHd]d)G/:\\U/
FPF5;NSMLa]PA.\ZB:EH&eU7&)Yb7VCffZaO36IJKH7=XCe\Q2,[G<(1-7\XWK.7
c8b8:-/ZL\>1VLBgIf@DBTOK^@:Mg:2.6_g_gWC;\=O<-HB=Qf0e8#WVKV_#7CEN
OM(-29TPNd;N9EIGN.#41)W#I7#,+-B^,Z+;YLdE&d25F()EYPP&:SeQ=?fGJES)
Sg7F23R_?N8=^+dCK8;Jf5/MX?KR6[7_+Y8T83G2J5@@)AFGS8=/+\>RIFdARc)C
^[<@4LUFVDL\N[__>K^/3V)R=DZF@>1OC-:]T\3Y8((-]/[++QAL1F[-0M+[^<\<
2eR(\B5S^A<PJZ?>Aa:.^M0<?+5PQC<CF[#]#Ub>Ub#2+&1AG(LHVP-f0?KE_ZS[
8GN1/GB&/(]Ma+-PH,A@(Gc5L1SI7@1926P.\Ae^bY;SW^g<?2^O3S[2F=fJ&F1L
f&IaJ3P:R5LRA4JCOg^;UF]4#b3g>BFY(:TIeUcFI>2F=f<8O#4=gE5YQf^GS\fb
X-=deN_d.Q;faRMV[9@0&04SN;LeMOfEY_5^@9,gW-)^:WD8N8ROB67K5gM;5Wd8
]f<4S-_51WTB<Oa5)HW&469OWZXS?@3/KRf9LHcDG3-87c.g]ZIQCB+e01I#8c1a
g,/MAP?\A5d,a<4=G4;:?7@a)Q]1-YNCb?NYU0YC+,f_be#]P:0.AOA>ga)S:.2,
dMA@^0-E]E5ZH8U@D4]30A1A?YA-Y#QM2f\dWBNS>O(Sa:.XX6S^1e]&X/cRQd7/
MbW386;<PLO-WM^.P>+e(S/<C&#_ZPE:)ZB.f6&B5:/@R2gZN1[_?&&B2B__@8R^
;+\-4^[;,2UQa]5BQ^HObfS<^]2Ob-1D(V;e\Q&#Bfg2C;^ZT7>42+4T^Td0_)8U
7aJ=Q6\f[F?NMaRY?-YHFG0#DABUK#e>P]:J_-F\fJbB^WaI<7bFWfHM:CH\8+(@
ad0gA:1EM&\AK]GQBW[CV)#7>gCJe);8:_=3CVcXB.V1YMVW+J-8+=Y.f)<U=._a
ZUS8L-+Fd09F;C92.T&:?17/78K[]MU#?]I?6:@BAOM)S:/#C>#O640U5(eI9T2G
FHf74eGR2K(F[&7OZVM,?M93Z7WA,>_K6bD07Q07eXC&I,2PID5c9U\3b_K:[#94
F,cT8-]3YB1(WPf;0=L;JSN=?H+\.fNd8T8#<C7X)80e@P<BK7#R(]2<-FR2A#7R
[aTCWTU:XATc3[L3V/^N[bVZbg9ZC&(Cg?9:N#^ZF&5fPWJ:U+[T[a7LT&2.]?+0
A@K&.)^c@4?-W,]fG.KM]=8)?a+S2Ga;L0R561a,FIPB]W5=32KFMLXgWFNJe-bG
BW3.UU0AT2_QdG\\^>HQfX7XcJTG.FTfAR,Z+Q>.[gR4\C8f;F+]V<]MbRU(&BV;
NID:.2L:GJAK09K13ARUbdFT:#b)P(\O8OaBREO^O=TC03=O+_.d5c5]L5AEUAe&
7HQ_L1]OJ&.O/@]N3>IJKUL9=a/UP>\M<e1N@7\.S/D1=Q0^Sa8L0G:1&VZ)aVEI
@f1:#Y#MUfVBTfZ/,ZSCSY2ScYc7MSR/AW-./BNS4P@^:P57HP(54MUHW_C9Yb#0
GQ,7-3T_#:G\8e:?8T+>@a1.VJ>[9de<FU\981dY]d>2M6QK1(4c.HVT#/_Y7@Ue
Xb?[7.bD25O\)CC;#=S8:#K9?88#cI^D9&T8>1ZYZ\>I,;Mf??MJ+W5_WM2^./F)
2=@=6W:-8aBYA8&Ke25VH\ebSYK06BJ4dLTS/aO]WGD4F[U/.>;g?IATe5/K0FLg
c0Oda+QGT6,Ge7CWKS)FU/VO^GOM()2?b,2RF;CQ]EAa43bR1?G?Y)F#3B_ALJE]
TR6MI2?#U(aeIE5#A6=V[g\>Q54Z2QAeHVA/N1Fg]Oc=eR_G>]Q9Sd:L]UH\YK[@
8:FN&cI\I6]_b2)\<ITNcFW/SbWc&B^#D0MX\IaU8gfWBdJQB?(T;5/;11_;#N,P
<@Kg^9aQ7ZX[B4eTZK^:F+J#DJgF>)a3f)\]@D3FPTfXB&BabTO9#.ULF@3Y2L\F
B\T9g^6H<g^=.\g,E.,/S5RD.P;]Wd+H][T]#;LJ-,<.HF2\CUT&..bdD)bfcD7L
X^@-_Ta#9TQ1XKSQ27d^\7_<TPAbec&HP]Hc)#g:d<&E&bR3C1/+?0I]e\P?CXYd
2JC<61L0M;VZYge.2gR,.CbC@9JbC3Q:X0Ma_Dd)S.D(:K[GGa<cD6J1)b.TV(1N
1RGXKdSS88]6bY\aD2SV35P&fX/JeVB5[^Q\Q?.2\=KQ)#EB=XFe4&U3WTLdWZHA
e+A&RgfBUA0,494FS=96FTK)RgA6eK55WREKN74D-X_OBP<aJ<8H8U[g8.fL(<E:
e2T@g9FBdJK7&bHAL15Me<J/;H#F>^3)g=UQ+He&(LX2=7E:ae7-Q)GeFGA4d5VV
53O6UM.(7=dd2F<?0&1KE)+X24HR?-e^F1<[??H;a]S/K7,54X76d\BB]Z9A/\eN
X/+^(_S1e<;;&Wg0g9\aSO0Rd3IS?17G6YafO0<(VCY8Wf\T>0&NDfR<N@67>,HV
7eH\:.Ucg6D:76@P(FNU;2K55K8DME21+@F]&,e1DF(?d,g3].-N7gdeT#aTCegU
BH3Ea.Vd8SdaKY=7Sd[bL4DYR=Lc5_)R?gG4)9XP5\H.3K;,HXe1L5]FZ6)<9TQQ
[46WdJ:JfG^HIB_D;CZ&4&AC10J5?.6.Jd<[E&&1IHU?P.E/IV^AM/_A2U#[X=KM
eD.LSG/(I2dM4]RX9YbXdc&9+)5/aN=\-_JEdREOP-9<30A)N0O(3KLFI^+OUVEC
QK#O1BGb+.^E8L/L5JeTB>[>:&.@0X(U70\2YZgZT)D[[c<_L3:N&2PdI[d)JZ15
M-3EF87P85)0GSJZ[D+eY=-T^W4E#6>-9HPR77,W&BJY96DOg;3ZNJWH0dVGDb6>
[C?#MY<2[8K^N50:Y3bM0<QR3?84:c9\Z(C<54##A:LBTP3(E)2A7)EV2I<?I7O3
Ra:V#;C>[^f\AUEbIV)Y?fWL:@UB(]DCTHF0)8IZ2+XO<[D\(OD66e1d:f^\P7&a
7HR/L1.EcN?Kg6<JL0QeeQY(,E?+,CAdbMdI;ccP4L4eQFIP6aDK<K7Ha,=,KNDY
GQI_<SObP\=]b^M]6J/E4<8]NLD&;27daJ@M>Q7?2#S^^=Of<9\;G4ePN_<24X40
QXa&ML7Od?7R:-IB]1/[\gLY_SZA-VELDFF@)e/J/77Y9C3WM8=6)f\BU:e?9/O<
>B7&KXGX2+LRI<S@b9SEP9=<)ZbVY=+FHV8YMHR]U6GccgV3I99>Qf4^ZY](OT)T
aC+H=I.K.Uf=QZe8d5=?RKU9b@(OW;&-f^??XBGORBQ)>OU5WM^,ZXUHJY344gef
_[WN8@UQRN78b[a:QO203QDNXc-Z)ee_N0N2)?Jf2F<-,I2e>\OZ_8.D@8^/TPBS
(QI;^M4eTb<]D\d^LY55+C4YRPfSV?QF?KWN3.0\5a:K[X9]DOe/_\OI84/84ZLO
<ONJTf>0NF,:YcM?UQ_Zd7P#>efGGc)6+1a58SSY>d?^D\AM=ec.aT=D3>+K_^=8
]-<;F&@^J)8NaOWDfII=E9>HN]48ST?N;^-e.Z94FIfJ->Qg_d+WJaaR&I9TLQ#A
H6C07+f<OIRV2,RHJ3EL=GM5Y.Pgb6WdUaI?U9,:09@[O,AMa/4UW.be@YfZaITO
E2,9-+c>C<XDC3;#)=U43VA]<18NDKLSCY&<HD^L_a-ZS]D@^[:b-J37NR6-OdGL
YZXb;Sa):QFOL-3D\83CL8Fb]2W<RY1=MMOS>.=6XZFJ=F^dNP7I><[CcX=.71<0
(959+X3b;E(FH=2LXQGZ[C8,g9FDX=]7[Ra574\Dc^OeZQN[WWVa_fO5JJ8YFIdK
fZB25E9/\&E0WU9^d\+2VW1J2,-(L.(6.20Nd[C/NWW2X0U7&WM@eI1Zc;K<Y;Tf
agVN5P1CE:C6M(/CgYV1c2gY[g3(PSXBWGK\UJRE6C:1,Q.#ZZY2#)4J?2?O_f=1
4=T5E<V:B0bF7O#XL?AgX[&RFZ@+[J?Q)R(UVK0?\]1H7I[d-B>^PE1JD9gEH7:X
MY)aN4_Jf(bYJ@2MUO)..W]a<:eFV.-00RRVAH4e08BVL-f28;#a4V5If(-D=J7T
W=Q-J]M2.?e(G<&2MP184PYB7:4bPTLW[D5]3XZgO_M2WU8/8EMY64\M0V/M)1Zf
+M7Q+CASfM(Ffa85UGd.OP]XDd>>@)f6:-FU4H):b:CC<U+TR6,+3_H_MK)_KRRE
Jf[;19^b</VaVS>a^d42g5UI?225N?BKK5GZ@JaY9\O\2+^]&YM2P<=[^A(LPJZ(
_Y0gI7U82b9?=KFU]0P[MaB:WOc,VJ65T[bg/W/7(QW5+,]P+Z^c<&AeBaD9E\ER
0.RZ6fC^XC@;>,/7:b(c#B0#DHEV[TG_>F;Q29QQaX.MYPQZL?d>F7bO)J\SeW.d
a8Pg4>:Ke4);_Q)TEcgH\RP,@RBbS<O3ag>5KALQ@bJL,O^C;5I5(3L(D&.6=I7.
g-8D;2\LN>W[1gCXTKX+F3N7^e>_<Z,^>+I&QU)@35O\87)M0,L&PYJK)>CZ+_E@
T._PTUPRJ>a>6R1Tfg-:YcTT&4+a<-R9aW#66S5H,7V+Wg@J7P=?[36VI6A/AW,2
6U_c,Y]O3>PNSP;#EZBL6?:05GLc/61+L5XDYTP/YDC<@:O>;baU)2FHc1O9^g36
,fGd/g8,?P.C?D1A_LgY&6I/VgG(e<)[dNORHGU1?0+DD=<XN@B+JRf;H9I]U9@[
=9\a;4YKJ,f&5[&7/_W[96L8^G4CbN4U,aT4@A/2]PA[A\-JN#b^86</[6Y3CC5b
UJ39BfZ2XL[RB=TgEdFe9Da+>L\(KSI_5,],#3?(U:/9M96dJ=OV.&(/eJ^:H-=E
P<2OXQ;0DJ_PR2(Z:]I2J[CT#:Y[RfVW:eWL[_WZME=L&TOR_fAN:^7TZ2_&g=:X
M.RS;:T=cJS0X@dL?NC-;5;Ua#S9Jd8MYR>1@+<YG+ZOebe4C6NAf;IWFJ]35Lf6
4=#&\DVb&3XP^;&RJa\XM:;GaSFIRNJS+V:WZ2PPI3#JMV]@=b9[:ZP)O,KXdfL[
#d6HMKF&W1J3#I)4T(ccd/PeCWJSJ?[YAXg)4-A;S,K0C?U+,.:HDNV9..NabCI-
782COFS3:2df3YGd,BKFHO4Hc+#RM[Q8-ENDUX,\<bVD-Y(R1P>8Lcb8AUWgYfSM
AVUVNF]_T;gEW[;M?/MV#5<1NfN3L[cKW];I,S:[1VV20(B^Jc:H_2Uf5I7G3MYP
&@/65+F/1?7^H^/@S]CQc/6>..@,(4FLg_Z:1N\Aa+19EV70_3;AZG[<<Hc;g3E]
eNN4aCN7X)cb2AFF4@gQ=-&#?U+1[=4]V-\?[^f_?)]Da+&#N8W]4<a98<)2:.Q)
FVZD@8KS9+F^UF\Q@C/S&&dRX>5_76AL1@8U(EQALS07^^2_ffS82:RC:/)@M,_?
]71H-e::eg3;/@SgG:K\:7#=1K/[0.;Ta\AWcX+:5H1b<H\R-NJJK(GdG;PL^22F
ZG\,5?dZ0dNVd6U8P#VR01FNYCJF3(H4TEUV1#H(VKUM/eZUgVQeTLI^-TaK]eG4
5.a=3#?VTeeCUJ8YdU=CeRHJ_(NE8Y+cHeC4;/FPTSYCJL?S:V,_R@OAQ+b5AOG8
Q:Q?V0?8+)F7-@cO9J/Ve?#DT+fCA=2FM4,2MWO@KS(I6FB(O5&GMIVM>M3,[J)L
fJ>^(/QBD6@dP8]U0=S,GAU=C\9dH7>X82X1EC\>RN91JR7\O\SVg]HNBV0Y&C00
cF>:V:2_A&=7W[gN-DcYWQ?4aPFA:.Ve_JSL-ZM6AXSCE@N0DOX^0E)Z;\fL&cIf
)9=,3eW&e4P1b3ZHTFY@Sc2Md6_CPEC-cPUCBYWVQ]3[64J)dO;<.-K(@^^^<W_Z
&948Z=1DYVK90BL,TV/U=)C8&Be16NA<OI&ZN/A^1FeL)cK?a)>W4VPJ[e[R[,S:
&e<a9+f,Q-DDNF[]3KEBDL6>6HN-F,cM4;Ya65Xb_XGS2:>80KK&UF_OYE,Xce,D
47;N(R@R2D(a?9-Eg-NdC0SFfDaTGB-VLO&_CMT]S.1D&>]RS#G<#=ceT.9#9BV#
O0U:_MAO-EbVY1@RQ,MQXDOR9^U#D-W)a<),T2e+Gc)L7-H@>ZTGF6^(_SE/GH:@
0[#bPLN]R(FO#e4#5(I3d8X3MDNa+0FcbBaD3dMH+Oc/<Z^7Y;WY(PJJb1_ZS+_X
U?_CE7L?d#<3aNQT_18C0:bTR3SQWQ[D82[TJ?:>KbBETO#VcSd22AcbOY;KZY5I
Y?H46?TEG@OQb8#))]I5.XFMJ/GTU(Q=A6PJVK,L]Bg6D:SRJ><YEeQ&0K?a_YE9
F+>)a_eBEccTBK6;,JT]8PAWZA&TLg6(Q<P@CgdYF>aLYSSK&H8EY1?B5a^a^a(.
Z[_F[BH+,#+0D3_f7QbO,@O-T-WCLbW-V6>_,f+?H],4#M]a+K#_/LO@[gNZU@L9
99BF\_--V+K4R2DS2Me1V<79B-WVc?][2ZccWfP:[027>Gg4AA1U\\F3g,+V>6+?
bDN>M89,;fB\[63-\NRRXg&a=^?R@+Vfa2\TN_Lcf+#XAK;@MFHTT^[IVTDYS^@E
e[LH<E=Q7YZ50FS5O;c\g0V>E=GdS+Hb8TMH(A=;3-Q(3]Q0dM4X9N4D[U7M2c,0
PO/JaKL[S1WD0Y26UZ<VZVF#QgHEVF3@A)NP/K2b_9e<UbV0N4g_^H[1K^[28e/]
&/HKfRS4EEJ.CISY_88.YP&A./=X=41=b<&Y#a&(JZRT,_4;QK22\T5Y9f=TGG>M
S,gD.P69;e4VH#dP[:K,.9PU50;H<[Od?XR)D]&SU\ICF:(adMM1fF)4EVd9UNTU
4\\egG:gG>bEG,gdFO23?dM<IP,U<?6\1)ZSK^LVdUF-MbYGdE=L3#13<//WEc5d
RMM\>/gJ^a:R6ZF3,QH19:d;Gf(C].D=D-VZIM/=?,KBKL8bXF/d\L?PZf5_;7U<
?2ZB,M<D<GY#S[[ZB]@)E]]ZYMC</9cf1BNWFG+QD6c^^8[bf)3S):BQ_NKZSJ(K
188KNI(A58FJ;8=WC^I@E9A@EW[JPFfLJW<FDSC[H9RCIR:]-&GT54()H/R+(,=A
V191+7C&@SO+]7TF+EE[5Q,>4OE-ZXJ1R)4/cd@CVBJCI6J4\V>+5.\R[F]0I8YJ
/:#3YCKG:JB8-6:]69X<9UW-Q^6A#8/B,_5)M;Fg1M?d>4=&c9>_VgU:]3IT<:ZW
0-0&>gDH2;Zg?K9F=e9X5WgR9H_fUgF_,gTQ&2UKH\21;^I6LN>Xg2372,WS<OWT
ZJ;L:@EaU^Lb9P#^UfF,4)(\=?>C3:(3edIc<MTON:H&,eVc+DBVI-:RWF8Oe/>;
UO<d2Ka,9#D,GNdNP_SFI2Ea@a6D#KE8c9Ab4S#F]T<O6=N1SSH6-@D_QbeN0W>O
DVfBG-g^7,54Y+P(3RddE(L<bJDeXYWD(KeBE@cECVIN675=-LYSM\6^5)bB_FM>
R)_<T+c]=+BDC-9.5N?d&+U_(M0R6]7C5RW0ZON#DgA_cY-_GHYK\1N@cL2YBE((
-M&QcaM#>;/&RVNG2F7B[cWZg;#V=?9fEgV3VKA3#.YV7d/N:==cIFE4?V_eN\4E
4?PVP_BJ(1bbRPIU@#L,Z[Edd/;>Y/-I[[EQL+0>JQTYXCBJQA3B4MZ7JOM@\2KY
>=G(MH1<bFN0Q9QZGS@V(M:TSN7DSX_;Y3<X+aR29BF<@J4D=4:7/IJ1SSG1-A,O
G:0N&e:b3GS.<[VBeDH>15,+bIN:Y0J)FTEFL8-Z\OO+5K(7R+QcSJXZ8:\e#X6A
F0PROg+HRTSeI+J48D=SYL1C2Xg)+N:B(/Ud-<[f+<Ld,J8N5^-KS>-MaEDfSSOQ
Zd?X#8CR[f5EW#WPE_W^JE^^YTdZ\eF??)Z,2\,d,/[P)E87Z+c>N9HAeXV^C#)+
e]0G=XbOf]LY_\S5^L)b=[&[]NM6Y/QB0X)4OWL.@O;gT[[^KEa=0<g=(_P\1.,G
-D??/Q4d[94+4VN1,M_J2;^OS&[9,/8Z:.;d1MGZNAW9c+]<-(O.[d@_X,>fVa&<
?^K_?5#IP(PUa&=SWLC:a;W94=Eg-:cT+1E)[SA:N8YA860fM<dbKAZ/+Ze(LgIL
G]64FWc4U)==(J.(\MIE.Q)DBC;.]X=UFCWc+S26PI0e71&EUDS:GCBGg6M?>a[V
BAS>ORQ31GD2HN<>@a-JZA](VF@EIbTd3b]Y);9_1H_W==JIPV+6WCVgXB>gS1BM
[\YB55_@5H\,TDX7/DZ??O]>Ne;XJIFg=D95;49TC&@+>9_(T(N4XZ.L5[2_?F[+
K=UZAF_0]9ee10aZ^UO@XN8</MLV3Y)[^d.[B+A&X13(6XG^N>,>TE/:,GJZ<=NT
S3EBJD1;V#2CM/3eT42fV7I^^Nb:RcOW:6/E<aU/B<G+_6-J\IP_,24GD0-;33OM
Y>)]1]AK<GeX[@<JVX8=]4>N&Q&M6GZ[Z2b48/N7:NS1_/DFcaa6L=B.Z?C3b84Y
W,Xd0<YR&UbGLTTUMN;R:g7NQ2cV<Q7ZGM?>_/TP;2(2SS2XSQccAe.V5X+ANa:L
+\Da@;&BLU<<H1bR=AKA<;?M6fKUV)I,NOZJ:(P_OFPgK6c0eKcEf:_f]QC3:Bf/
\72T6RC6BALaOAeZ)3Bc;_:V(&=Y-e03[g.K(gc^J=<LS[Dd-/Z,M1/b<5=>MKC5
26.[aZR?@N^(7c9E^HQNPC5+-daS0G1H<URcBU4f:8L4>)_B:=1,+eC8[dRX2SX;
;?4,=D8f8@7J8_PGZdHddEJARLE?)\G29(@GDUS51DP6b1QQ[MBGGMSE0@RJ]gOE
c4a-Y6@Y+K_(;=e=>QT#cX8NJ7eO+Z@c3G>g8E,),A=O4ACE=:8VGS08[M19d7a1
EY&7\3<=GeSDRRY:TPHJe73Q1XV9XMF3aNPB_\V#OSCQ6MLK?:+N?P?4dV8G51Q)
7>7N&JGJ.7PFR5RF,NZ8FCH1O4=aH<ea6f#KQ_E=/UPRLU]P231LM=&Gd?<-Z8;R
FO.YVI+O.Z_\D\=_&>UR\=]I@?I.6fM)/R@D1I8-/O^U^+3#=J#R)^C?Bc>39T(\
gSO8b&\D)/P:27AdW)Y6II:6gDMAX\KG?DB>d?4b5TYPX9a0WG9DMa?4FHFQTBT/
-cdR6=g]N9fU<<P=X\=_fKIS[,C<QDAAPEN<O\gS#>6>;5=<F,DUB@FGgN3NfL<B
]TYAa64[cHfB)V^UMYYFC<EJBZC4+;Z[49e?K6dgK0M+3+>51d[FQ1J]/SHg#[X\
AOf>.ZfXDEYR3IaN5TLV593[aF1.X_LO[Ke=\E[0P<FKWAFRA1(Pb@,848B,,@C8
CX2VCc<CG5O8?d-Y+TN?b@C6V6:;dEA#\AI+\0>8R3fdE+)DUJ>ZUPc[S>a.9#KT
R3PN#IGV388T^R#\>fC-D:>:JV6E]_+@Ac,O9491G7]TZSBca;M?5^]^L.OWdYd)
V+6B7L/5UX4(OZUAATH_2JfVESV.7,dcF\<0@V<^6#4IPS+[>LfQI7bF[,Y&7,UV
g3DW>6PLJ85Ne7f+IVXB,S#W0/ZETOV#KeKEORcd4U\#b/JOT;/DOWD]=N7^J7[Z
L_K/\98186KFb,L-(^Od0E9PV0^dYH)#<6C.Le[Ra08gQDZMKb79_H:R2(I8[L33
Cc^U&]KPVdeGg>C;EFT3^V+R=)L[Q8()B=dA3GdUbf0Z<:C>f/(;(Kc_7JM=H6X^
A<;-<ADeLA=;(Z]44VTI/)938eD\1Q,=RJ5^RC#^/T?BFZ[I-]GU8+/MBE#\YA.W
dY.4&Z.gZV#9PGI4=:NfbP\.:3+c^.D0,b1AQcDZ^fPge3X(@8(3,d-.ZfA#<Pd]
L:D)@AT14[=T@K)Z.>+ZbYW6c)2R<UHY[Bg@7aZ?7S:N3DL_T0S.HKJY)bJ2[d>X
Q_Q_TKXI1,=RNK>MPJ,b^0Y&[+2dF4.VB\HM)TgZ)CG.H,Q1#6T4^c9#gY@CCc/8
0,E(-AZc,6,-X_E9^OI;bd@f[HOZLWU.?WOICVFPB9.-T]N>H;MX)->A38:0g.fX
S<GC^W8LED1[5257BV)e#)2<44d7W,1d[VWY&;2-]0^,I:C.a;G#E(/123DV9:Hc
&fMR>a7QA1QH[g+dF9QJ<.[])AL._Z;X0@5>O#/8/][9,IH(8S0VZ&2-J2C@H8gD
KN@\Z8\[?ggL#[-3?CDOV9ZL?<?,M4]9GY?Q=KKcYb^6C#AU9T:+HQ:b#6Z8X=Ce
ggTC@W2#LT=XON6T#):>\Dc]D?(-N9WEcCTe<E(V&N4^9_BL^/(]V5+F><Y4YMM8
&1KUeH>I:PD?<&Y1.KIMP&L7f4?c<_S_b<Z&&0aa366NOXW@;-J7<VWFPg6fb7JW
fGaeMeOSC^Heb+@PEXH2@E<b&FWK[gP_JI:&A[>&TXNV5DZB;FOB#DZU843bd>+J
E>D(L@LY[RF@=1aa_/A\H[2+dLDOCUX9C05/d]J=[c=#3(52+d\I(6Z,VB,VLV\O
?9)BR:X]N:]K\aN(IX>@XADa9SJD^aU>IMHB/6)C7@dgU&.:]c(WO)]\Aa;c#];C
b[>A&3UU=-7LD\M\U@\[U,JEQN;9-=+^[Q,8]+NY?#L7gG[QfEfI3LYJ9SK&-)S5
UI3=0<bK3J\3JUTJ2.0M@?.b:e-IM-D,c41f>I60=KW9+f][0^QE&\O:K<2OPbe3
E/JF;.KaSF6bLS@(X,J\T(QU<U(?-1=g@DL@ZC04Z>@9Z6]@&1W/7F,I_&#c4/6b
<Fa=>ZdTF^bKXCRc8JH8X?#f2SQcTUIX7+/5#Z/a;_Ja_f(AYLUF\_;#LIVOAN@P
UXB[SKWPAJ(FgAd&L7b4;e(=4.a)Q9)e7dGS[;ae?MIc<99;9O02FG?Af4cZG&@f
8fKQ4=?SJ4>JKM)ODO5KIb7?G?FGPD3-fZB^UFI@6O,X73RfU[HD^a(KZ6H\>R56
C1<dD?BWdJ]WKDCH.G#bN\d&2OVZd(&;>AEK,,7-d><;dITFa]/R@JY^QGF^432P
SJ_2-aXQd[-aFYF^EZDG1HdWNIL5gA&:Ged?4I7BaJ0&e7<7GFW,6f(<60&bFL>?
7/\/Y=<HJ2I())6>T,T[\K6@d4.UX-^RK7182R4+G:VK>.A,d<C?f:>6Yf)2.]J(
87=E+F-E6.^U5g.G6^JMI#5_H>da),aT+BP=L/;ZLDHK01FWD4Z_-Y9CUc<SWS2N
GL(RRGR+(-]cLURf:E\]<@NZ+M3@M.E@V_D#5B01)9R60L=JU/?JWf<^cIb8bZ-&
4G=CdE^>VOUNN4eJ1>IFdTA]K>g4]a&J6=-VDgTX:/ETG-b9F/^(SKV2Uc92+C3:
H9-\TLV[<@9EcPF&@=2O3LadD6MUOPOb:TZc?.P?PZ+52afDUaEH=(U9e0:=JLcE
+3FA2M\\,&M#4b6JGL<YDI[IIH5MJN8HKV/gObcT;SXAXT.43DdHA8ODWYb?KTcO
EI=d82TG[RP>;.9/=DO1TQ@@@5W;X?6?1[DI4D/7e1d08XS7TYG]JA+X[d#EE..L
\dO2^KWFDd.d<.Yef@JfNKaMed>Nb_97,NKK?\T4M@^3J<dOe6a<>^VY<5Z\ebM7
/;Z2&gARMC[B0S)SOa-K?Q#CM?#66R<[AYVG#B,PY]W6c+N6H>^@+-Y?6)d-Q6.,
\DYYGV@KR&JGC+RYDf[WDGL&Jb@cQ=]EIJe+AMMZb/ZWc<=@J-8O2M3S3FQ/K<^;
T?gHeYD45(8D?aIWf(M\55EFM2?OIV1-12Q9ZIdS7Fda1O]UQ1RcF>)6S@-F^Ka?
7.<Db:Y,N.QdCU+?681[d[2W>46UVV>UMS)UBC:1+M<B^ObAUS=g6J(&<,])F@C&
X58UNf9D(&#DCTaT3:?_5c6DMZXaW_,0A6?+^9VRc&IN,KY>5\5C<<a>^<+Be;0>
=\E,BPCeCV7ELU(TZ>)J+T)4JW>Y-d1)1F^a\Q=KZ<a964Q?IP;Tf7Z_C^Ag:UN&
S<J_D-^bSPfB&E=\;XFbAcEJBITPFfd?cdd+_@YO]1TC2dV/R?9c(\L,.L-AKVS<
LZ6V7<bDSX=CI5&DM-HA1[\e@:X,71ZJGIR[E6ed,Y^6HdfTfF7?.g4L(09[RP+(
,.<TFC82bT]#=ZTF]XWXID-K82L\YX-[I+RD2dC=H5I82#O63W7HHD4&4<U2KaO_
6GK,\[JU)RKg92PcKU(X6GXNfV,Y5e]R[>ED]a@)OHRWK#\YU5I4R0Se2cXLO/Z+
aO6D^BSRg7b41=YZ\Z.N)a-L3\7Y)YV3NW[M,-=?A=M<aL0<F0.H\Jg4;HE]BA]1
Z)c_>3^,-OQZfb_TPGQ+3-6QTdO/N[O+QaO^>1Ce1f=BQGLE1HC#5\B[F6_DQ[Gf
^24@:W&>0Ca/\D5JKYI.,F>LU@e;STd(.8;46e4JOQ<HWXT>JEE>OQ0dH;#_3:Mg
^:[d4?SPAaON/J/#(<R3;Ca,]9G+;#&3?BcM4(Z.R5^Db7TOC-?50@+@(a9)WIYM
3FYS#/U\D4[0THS48F#5/dbFgJFRV].E5BL9;g,PYK27g:Ed#2\VE.=_RYIDG+&5
=Y<Zgb9K^,LFF2VC,Q^__3P??>D/gQ1D6:=/.YHEBb5VSN)1I9#C9LS@E3-+f8.>
9WFJTW_>M92KJBZZW76a#6RWE4,,A<R#F6XV+,LS>QEM/JNgDG]L.e:B:7Z.b^@R
fK.dWa81.RZ9]]D+4<QCW76BVabad<PVNWL)O.fUIbbTT75-@]fG)29KVNJOa./[
/L>QFeSb,Ye1+[NfZ0=DM(4@eCFN).LGI##CUA1KZJ-LA9@E:@P0M,3:gOe,ST#8
TU8Z(N@6GYc_)XcMIfD1cFG6G.51;H9Q&\WF;^5QbDgIdC?J\7>>_g;SPPVRI=Xd
MVBB;\TgG_[KHSdV3ED323HXOW^((9U#9I3DeC:QZOO/M87I3S.MDaNQ4#?H^)O7
.>QAC\))V5_OXVY4\@A]&2gGX<d0Ye\Vc:/1;0\,2+f.^)YZ96KNc?K\?+aPEZBX
^d(5KWISZd(</CK0LOFbbFA^G,EZE9[FEd5_DK[&T6d8^aa?g4g/HM.[E_21OR.\
@CWL3XZ4GA7T.C4GL81SAF\gFfIZYcV55X;PP#e;b,dU2cc):a&MA]^Jegg1MdcC
<#60@S9]HYAc5XgEN3B]RHg^N=.bJ(Z3gO=B,4TAC0<WP]cAB#V48KGS1UKXg&fe
bU#QOAE&)WAQG,NaDS\4P,FN^>Z?(J;&(D:_RB[a_X&gR^=Gd\06_812EJg.E:ON
-QA4EcG-P@P(\</,5Y-;E_D+gBEUML0UJEF]?7/S6?C?56W5;HD_:@&d=ZgH<..I
R5XFI8C[B5@XO)gF<6L/+)=4c&?.HX)Ya#bf<gZQE\K<_2B6gT>NLaO?Cg7#W&]<
TMX=?[6=Zaa/6FQKO55)31_QHee42^:7]]5(d^Eb/6YI@b94deCMP4/.dcSSJ#Fa
DU7@ZX5LSD/H6Yf)?S2Q4b2Y&0S.B\,<B6Jf-Xc1PGR6HFA@S3=OD_FDYS_5[X0>
:,,<CL:MF)DX]Z/JMIV[^,Q(?WNK)GcedW:Q(L&ac<ZV<g^S<;/d;gZ_g?]3A9@>
c9J/^P>g,(d4)FJX:Z:0]bG_BbSYMUG>6[>US7LO=c^H_<A2S@+05DS=+-[?X9#C
46U?J6A6A7BSMb@8[cJ23=.5T(EaJ4RSR,2278cD1>BY+AF^,LW:J#dZT2M#/4bF
IgC-a(f)>I6_gA57dQ#UEIFY@17XFJDRC,7CK;-)]NL-EN::Y47=f-d3E33>F)7B
FR9K5A3;CKLcM[2TLA5/CO8A)Y#^3P&9TgE]P\8T->>E8eA89OeDG@a?TKfQRFfa
@BUf&\?fIR,HR)NJbX_4BHBEdHTX3_:f6L;9?SgKT+)#E9Jf?W5;O5.]CEQcFSO0
RZ1cE]EFB>2aD\R#Y:0;(72=ad\C<AJN/H7ae_6H]XB3Vb\-B-:8aQH+fQfE+?2T
:Jd#U(<,8ZUU_?:7&G3U7(QRRfa0Ke[Y)0:7,XK;E:179[2W6#QcE.c2<3b>;S>X
[.L35-d>7.<\MS-5PeY\AS8(:(fg8YLMc-)H.&F?3O539K.,b>e\@X1XI@YS3?4e
F&c(]\Y&fdY-87X=:1V#/JHY/RJ3Y5]IT(3/<5#R,>b^YT799)Va1f@B=X7@(Z@N
ge2XN7[U>U,_JC)HTP):G-6c9Od^NT-QcZF>R1+18PSK,e/E;9EXWWN7b1/ZgFI5
@AHRH,LH^dD&<=:^c+MPVYSOA1#GP&R?;R5aRD:PZFF=aeM2Bg<65TOQ5(>JZQ;&
X/]@dV<2T<A6C&R8:RYc-C[<?U:R.ZUZ>a-^87T[A2^Sg5V,ON=U=4dLBJVcSUK7
?OCaE-L4^K#Y=Lc#]^\TQ(I,)5Y>F747\#2F9aK&(GL3d?Y9Hb>YCITCAU@RA33O
&5&DO?,)aBSN#D+=Z<FVXK24OA7:deeb:6^7.#@(B0R927T(GO#D?#[I7^e+W@Yg
X/=,GV)8)XOO\dZTNgMJf(.5PS/=H20/][[AOE==Y7M-SREFN;T_7\@)D<W1<(>G
&cX[9>PSCISdVO;R58)Ld;_0X_fgQC,-1eWEHSSZQVfZ,MF;f&eB:-F7_0ASSJ4e
T?NYE<>UHKB(&C_6F1MH3V2.A-+5-M1C_a:DGLU?09RZUS27Q1SGBd[UYU;XPf_N
D@J#8?GTCKWGPAKLU/Y([6???U3LI+H0]N)^SGZ6A-0:Gc\4W:O&:f4cDED._E6/
=DL0#MJ^97A]X-KbJVcM[6T/D0G#S>^IZXWYS?[EHTL+gdCTZ24a,Z==:GSA<9AO
D;[bZ?K?B\S-+)=7MKRHb?#<I+0@Q5:L5P7SG7P;RXL/HL\206d/ZA/+XTEe+_1B
V.Igc09M8CbJ:0PbC1#@40U\S7\_fLf(;)6HT[2d4Qg-^Q+Q]/DbX.b(+;HBIMM3
BFX16bS[=UcALT-0+I\A<0]F_PG/DCbQ0.TZS?9BBA4,a2NM,4a.=GJdPd^VULGI
ONR(372XVDYUM2G>S6?F?64FC:HF^(-#58Y<INX#XM7b2BIZH^F#bAbKU/62bW?]
+0.)M4d3Y04BB/A]8&Pg\Og)B9X.GSP(V^LULZ=N,=SAYP@CI50d1OKN34/U^LD9
V>N/04CE[Va@#<#0L1NXTLJ[I[ZYNNg+V#^ZD^SgM,eB93G+Z8J0QJJ7_4<NZDIC
Y+P^=:,AR@#JORUg0HO6?BR2RKU&6-:8_#4g5g6;^38d5L^73^6>U6R0@1N./E+K
g1KU-bJ,D-+71efZc)BB@8RHAMY9Fde-(d39QX>?:U3?043;U+^I]Ia-ABf^e,YT
4-g<g?BG8_5XgRc4Kd5;)J.18GOZ[HY.2<K=BZGV)<-7Y(We^CdWF==<7\K]KdVW
:JG\,JLc5_dc=H.O5g@eL_M>Vfa9[33+91>C#E9M_QLVfF/@_=@8AfbH+@@BEgP:
9C,IC60c61eK?)VNFD]@5ZPD8?_X7DZ?W\J>;H8Q)2#CXO0.OXC7.Kcf&NSF[a+Z
\)3.3.6B:Eb#Z>,C+7FMUO>4/(0f\GFC,Ce9\<K@M&?Y?+NFYC:5UHT._H?0TeTX
g1=a)7[IcNY+2(><V6UM8H@P70L3W5CK+A3>;GC:XQe9AU.Z\/Ee\(P\<]Ya_?_W
\;g@T\)_A5LGIY<8]C^c)E/-/ed@OZ)6DU7W-IEKVR[a.1B#<#5M5WTF>?[RK2]=
8=NIfOAE]aHYTPX+#PVgZIeK75f+-F0(<c&)?]2_0@WE-#OHUAQWUZ<c;T93)[BT
.a[dC(7VWFFcg_C#FH-]WbfLRT46#BV\GM;daUb6IJTM0K/@K<X6bB-LPgT<\LbQ
9Q+c8,WV7Af&YA^aIfF8:WaS>6:EY#:=e,H5DRJZb]B.:NR.7W6LV>Q(L>.6;F&]
8ACA=@bVI_gfN95Z2OB+2>Vc#<]Of0Y6C\=Ug5)#FYZ3N+2]Z+#[8L?BDN_Tc^ZT
><,066#[A#F8TA\S3Sd<HcDGLCC+C@Tac>R=9V0>68]V0Ke3VT76[EC5??2M(/Y6
I3F>SGG4a]?^C+_/A09E^)6fPE)-aJDCGD0VI-S8E\g:+>b>Y[(Q&T4N-C=(S:4\
\2&A7g@8VYL\3KG8G4WPe.MY&./I7dM,U?X(SW8BRE-cM)J(6_(<Cbd_e=3ZYS(:
N/KNYX,.d&^K&TU)OEC_J:Z>&R@0=ARAL+MJQ&(J4PN#F<:R)^DU73+7(NEA2P(?
WNEW+YK]f2->Bbc>Ma:LeYN=K#IA+Q;B6:8=70)]6SEgTY?+G3;_CE.5D;?\_JB2
I>D@8VXK>Eg9d[I_VQdRA2]^-\/NA4#H>QM,WC3Y,OZ3QUS@C)Zf2eVI_FQ9EGEF
1/V[c)K\A@NUW+/LbK]\Rc8NKdDHg1<UM7-/<0>&8aQ]?/g=<=:2Y6[>DDHM9Z]&
gQZXAJ7X&J?d@C&R?.@5Dc//SD;J.>+_6X[C5\B,JT7IgQ]CSC+HcVM@#P@PIe33
W&g-b_+K8&111/U,M3.?R)D:4DXb#;(YJf.1C:;/I)Z4]X5>?(1Ta,DVHfP=Z[II
Q^AXT/>^BL^>;SN2[#(HQePX)9@GON=.\<\:H@)+Dc7&_d2X:g<N&?N5dYM[ZeVN
G42>DR;10-<5b,YI5I;62De>;SMT7\[\QCIBY+?-66Z_GXT@H/E-1a46POED(>&+
#@Q;YL=4aEPMPE\+LP;K[cWWW5LQ;8@+V;QZ;KTJe;acNPbE#QXG\fc&69&[EV5M
N7SH#UYTMK4GO?Y_f=3Xc1[016_M3&cP=A2;e<I0c_5F7Tg3V_6Pc9JS6)L4M=U9
+Mb(^P-<fOW>9<GWdMU;DE?5fU?ffV0df=65a+].DVBAId]eTQG057+Tc?D(BeeE
<#+:@a6G<eO(1-e89e.QWQ40\^QgO/L.8TA/O)YgR4REB8,#PUP-3Kafe-=EUPEP
0g9V-8IR1CbY06<(:Q6LQF:WT/cI3MeC8cG&YG[9&UOTVJE0D/PUW-GTc\_WR)J,
7>Ya0eZac\+A7)\=5F1?0:[8c1IHRd6[.D+2F/97,Xd@75NS:+QI-:95ZE0EA8Wb
K)_F,OCV?(IDX0KE-NE0\6P7NDfT]XG.J3T0/<-Nc2?BGdT\.XS>4IgC&#>@J<OP
@J6_V(8cJF3-#SK8LKS#_<XA#cWM&_^@O\,[,c_&016VD^AW^1\8:+Jb;])dd_VP
VRD7M-cMJ>VI9I_ZK]#OSX63-WMd9J.2E.2FYWS<cgLVUHXRbZgEE<+S#HIZJZW?
W2<6:dPNYfHAf)2CTHaJg.\LCNL<&8KG&XC15&fS47gJQ3a.-LC@2P179D;>-&?Q
Za]8H1UQ#1V?V<FS[4.Y.?(X]PGO/-+I79#\]#\M@KM7^QOI9+-T]0[:6<8#)+#E
P+QO1W,U:(^EDX(>JO-C4&YFcLM?gKfSB9^5#I&FaH2JK=(1ZGdLP@6Y@Q_KP:5-
=F>[:cffS7[G,>H-O\7<=;XN_D6KMe;6F=AU.QWN?8[\3aGW73^GI/GUH_[R0DaH
J\CA>S\>K]4:E1A4;d9+;+^ZVEFgS9\dO&IJ,ff=.cVTbS@E,a]C=W,:&53P4#.G
:IQ133A=67:?>J(X5?^1VfB.<Bg#_[V4#QXg&X#0aUTgbGYG&:#CFSTgR&K.]2FR
LA-\^X^Y0I1EQbcLNMAY;(WP=THNO@dd/:1WL@]aO-UIE][c_M#dV29LAQOVa3X\
DI5O1G5XHJ:S.GBS7,##f0)Z80ZND-@^Y::6]Y,/Kgb@^[g0F?gU9P(a6O80M\A0
-WT1V3#,<H_(N[0]L>&1-QgNdRH>(@Mb3a3)Z0.581He0Q_FV1?47SR2V/#M&ZSd
N1><N_IIMEe<PC\K[4^H@1/Q10@E/(dN0(g[EEC&7:B^#R@=)UFF77cESF//GgC/
]5NaRHL9U98=L6@1aY5Af+\X0\B>V64fee/S[b?1@:C5]WY2,UdDa9@7?5UU=AU9
D(SAC[4bSO5>7?T+OKL_BU-^bFE[89X#=S8D^S(Z-,AJU.d>Z=G-C7-U+0:\E(0D
N0gIY;9_YG-Ja3B<=0P/Kbc?6SL-f)J-a].826^QYf,,8032d7@0MLGVUa3DZ,M\
2b+:F&0ga-2<>G-97AHSK]0][\52\L&[F/LP5](_.]#7KbO2=E95@22bbP9<Gfbg
2)//@(c:83c@NV;CbRMGg[GbCZ,S63[5NdK#&.;Z3c<1H\f04B7T2=MDVMW7FO7)
RDd#K,BYAGOJN>04<^^RJ1gYKY@5eb?f^D(db]K(PL:=QQS+c2OY5_=ZV-7E.U\?
aS7R)7J,ZW#ZK=Q?bE(>7eD^BI9.c_@JM73-2[9Y2KD+HF3Z-6[4Bc21N4MeI,NT
U2#C3UD]P#WQQMeGZI8BBc;A05,.Q1>F/[W)DB(PK<M[T^8Q9^J7+AQ=B=Q.@dD]
7A6ZRe@dAYb>HZNP;?aCO1;-2C^0E6N.>=MLM,<>O\&aYGf(-VbcURX^Z@?=F:S-
VP(?_WcVe(.\=,Q6a>1eS7ARZN#U9KBK.+,#7_5<SMXPXS-81<JaEFAcN^.2__-\
.f+FXg_^:f)LC;N;_=@CW47Na&^J)AH,W6Q<&@3@.(XT9#^//02HS0fHf5<HUEP[
Q_I-Pe?fKKWK0>VS/,63SA6K,:8HOEZ(QP@Y)8A#dLOgePEQ&CWE90K>P[_E@236
e8g>;Ue)B?&+?/T-12,eZU7g<DcK&B_CJ]/I0Jf)6\CV[B+1[B?]IV=88QaaV7[U
aS,2I@SFf2.E^ObT]7CgM^F^5gBR\,f.FfHb2J9[J9D+52Yd_:O)Y&R\@3]<Y6>@
GEeWZ4I@=GP8bY?3@#2M/[[[9\g5a10N+b\M?2B.];^fC2^4)d<]+U;J]6[:,9]D
bOaJOPM\fAGU7P[FXR6OB_BW_C>\,.^W,]../J@<VD4FeUZM+g,R?)0VNM1+S2>D
^2_#Fd8=/f:C1=G/^c0)>d,BP)).2e/AMRIVD)Ja2RR#6gH5,b[3EgCAM:_MUc=/
=8If?2-CL2/OH/E\\?R<W1cH#3:AcP3M+K2[KTQ^(NR1+41#\LY6Z0FW[,OX@bS@
GQ^ER2V/C7>E#YM3;aP?W(2^;45&V<V=<)2IWGI>TS#,:gXP<GA/&DUQLTXa9f=]
=bKb.G#^X(.C)5FS9961eHR+^H]\O4bCVe\dY_;&8I@81WPRT?P=HM[EW5UI</.G
?R<D->:J-R89=cF&4+5AS==H)68Q&9>cVSDS^F/1:K+4.WE43)0\NX<.D1a:9MX.
.B2SR(;;K\HD,AbfQLK(,F&7aI1UL\2aDT3BA1?L9BSM1^9JA6KM<F_F?G-)fCaK
48OZQ9c=[]0_^;(\VC</OEO7Fa/PI(fXE=JTUP-HSB)G+_;/]\2e,cA(Ng>EbXA<
+@W9Dd^g9-A8:?9RBf-H>O@K:38BZBD,Y0#BN\<_G;=XG#>&f?TKBA[)=<(^R,J(
2&dU[-BB;V0DRPXc6V\TS-CaO+a[c^8ZBQa<O])b>DJI-E\(D0^OWS?X#NO7EK=@
7d&EB4)XANGAV&fCUea2d/,XX+b181E9ABB@.D7P@_;4+(eO19HJ\Tg6VR4J?<ID
1N^(W/?P#HAEZ;Eg+f6];0e<_Q<@<6g72;X8^701KbM;f9XfZ]8Dg,+(\^e37-YB
T5GKQRdS;9EcZP<MfQNB1Y(GOOe]8ZgbSYA?H06T7^MRWN4dLX#2NTCE^;EUW-TP
DaaKe@I[2JHLba637c<RMJKUCP0K)&]L3YP7J\_[+PXQeW[Z+;S>e@O>4eB;N^P;
JaW/L7+Te/D_?<Ug;VWTQebb0P3BZZADU^WT.K[5,Y#OAJXH#BO]+PS#c7KEOB8S
&=>CL@V<c)1]_#TG\+eX\>SB;c65E>f5JXCY=-b2XX-V+Q@H.AMOV+0M0+E@Y+1E
NeT/@=#QJZ46(AP#_UEc1IYKF.1+ER.f#-.Kf?/]DHb:#Z;2?E\8CZB9(^#&(,,\
.+R[IU&F(P40-82K.6@DXe17)VE;_SL9-?N1:\b[AWSZC(I&>2W0d8&(>^gbae?N
=I)S?8;d5.>O+b/g[KT5<?U,LJ(#E,W=FHLf4O@9RK?)75MMM0Q[R>.0?e.]eSBY
Z,\dL@cK&>2)>;;.^R;6AXYcfNSO,XS^Fc-B0[YfX(_+2CJF7LLX#3fMf:UK(WLK
Y&?cX65Uef5X\a06WL5M95WP>SIF>GD;+T,+A1M?9@]dJO>Y?UAEB>L#S#ZL)[HR
gEaFDV_)6e,D&4g[(B&H4D]]f]+bN8L>#S4@cY=&AD7QHcEfH]c6=/.7G8X>PQ@-
);/Q#^+C>^K/[N@Ag_=YfaFK2J5WdX\5HH>L)\).ZR78HdP;7X<FVRTdMZ32R+T1
C6;d_U-IL=^69?UU\gIL>-O\QEGG>C]@EO?1?OCDM]WO8N#@d.<X6QgQ:N[.Z;0S
7Ed_DXg2e>QPZ+.HIQ0_HH//X.^d#(MJZ=;;#_W-0_<D=E[]P+DU_Y_S3UO[N\[@
>5#K.1VEe2fSJ/0dUF(MeJ-\:Q@]CdGP-Da6bC/b@;Y0Z@C_TFZb8aGZ[aM>):BS
8I2E\dObcc,QHcD+_N?OF5WbP/6>B^d>UZ2MR<Z@Uc;@WOE=P2#76dDb=Y=-c59)
-A=>C2+K\g0eFOR)M?3P/9JW)OYDa.>-9eT&]PE7G4f(f&/Fc<;G.2E(bM5Y9#Z4
PG850&5aADKb4+MP]8bF@P7g168_9a-IQ>I^@]#I_b[)^Z\\PN=BP;A0W-.acCR(
LJda9g0EZQLP?NNUY:6,,;]:?7-_;-/V&F-51HWe]5(f@XCQ<K@X<E?bC1XNH=VY
f?3I^8dZVXYI0cWB+8;9\>=&N8Mg#Sbc0dLD]NP4F0W.F1(/^1RJL,:@5g:LDMDC
H/2=>H\0OKXf]Nd51R^@YZL4_,+;?4ROB@@O2ZY>L+^HH@L\8&Gfd>55_b?:3ILa
/XBQY[3_A.Pe/F;/PfCH\OBX/;cO9;>U@3WB0>8)OeC8&7U73(JQIO-K3Cd]eU-C
>Aa^+45+R\.CB.c1AAYGH,Ue64dM5-a9Wd4G;B>4U;?,.4>SKf1<Ua]?V5Z>a^6P
BgYS\L,>;]A2W506].HAP<dPCMA6(G)M1U\8OA^4/9/YP6NZ-ggME89P7ODP4fO_
>,_OG<X.52f0S8.:(1XO@8+6[3KY]adHTZAZ)VQ0KCgBK?bFB1/XLS7BY)bA+08F
d3S36]CL.+57V^#7>dbKPV_ffUJc]DCM4Z&\>\R9/^Pg1(GHO=1_We&S=^WFG&LA
<=JaT:)O)AD^X3C6[N\Q<-R8PE?aZZgS-e4+UB)>de;\gC31AVP6^Jb+\HJCg6<(
WbCcW7N_FRN3cXXYV6,-Y;5?Wg=KBE)YU--V^0bL-6K:&3UWP7R6U5fV^1A.6c\J
Q5M;P<bVQNOg;1:d:O2:Y=LXV[#-L0AKH?56^fM>D9XaTX[PZ+fT)b:f.6)@g\>A
fDE\3I7DLb89/8@TAO9IGNH+P=>M[YVR@J<>JgO+d11]GEF_34->1OAEY?L;P&TF
H,O&Y[?g,SH-+:/04-D,J>b&F^/b+8UBXR;C\g9D3DD[U.QUc4)X&8-,07U[DUA-
-gNOC);^:413,GX#P:aU8=2;eU3NaMHe3LO4BL\b\8JXIV;0313?.TR.\\F0\](3
BZI&XaIcL\?F>CR)?UG9bBOQcPFg[3<@@=aO,V?4?T0:8Kc_a8NfNC>;99R:&OV4
6aZWD(JZ+f?b9dK(5Y7<&A,da#KMS<df;aL#(W)ZN14=fa9CP;QC^58U>6](CX2I
X?J6-81Oefe??C)[+]ZP73Z0J[:7TaBMD?c-O>LJB7T3B63Y0O<H2Ze=O4f#@?.T
#U825LEeU9e>_c.W3)>NUHaZ)\[&GTT]P&Y,/[O=?U]M2.cXSX1LbCT(IRfDFcCM
d]N8G7?\^A+N;+=W(:#D^_MV+<>A]c[d[+a;F^>-a8C@db5E4^8<0BWG4;<_\->2
e<X&]<d1U\TQKZM,#]]>;W&GJ(#14CDJ;0T4<3S9WR?ZY((MWRH>FcV0Uc?N@V1@
IDDP>egZ8SObK7g@@BfP8IF=Bg@B.-XDC:@2a-c960EFXK.Q1+-^FN,H1SESGE\U
Y?F/M0,H:?5e4C#?>aBHG:c2ZVU6YW;\V3-=YZOVIc_D0A6eYD&8890BFE=TH.=T
9;(]N&T:X[^3=0Q80NW4F77aH4D?N\N;0GR85[Z-1fE77AH/,I+S5E)YMf&dZgB/
?(O\[XYR0gcDd).\#M1@DX8.ML2:PKGX:^=?@YZ<g_?LNOC>G-C^VSKf,UTa@.6P
=aW.@0[1>-O<4U;98W\KDN(7#cV&MIB_\I&,>bF>>]G8HYP/K(2B3_WFIaS^ba&5
ZU>XYLWcGHP=/NR.@&??fL=MX@cf?9J5XM[?XdPK;+6YFf7P;#1;c:N.e,(JZcZA
ZWY(1#;Aa[I8-8SW#D7XJ7VN16XYBTaP..V1\B3-;fg;?LD9-S<:<1^>>5CAXEe7
c3dc<ETNANNF69@b2+D9AfU-PP)BO9dP#A1QG]I2K=7IggF1g01HLN[/21@e6[9I
41XAK/WaVV.]7UZ+-IL65C.0:]_XQEH#b73PB#J0]+b>GQ&XPR,7,)XH56M23JeO
U)6<X^g)AB_HFTHE9^KJ/.bS-M+:M3GM:gL99U_W3:YB=.K8?V#g-&[.WQ\6D>K+
DEePP)/:J_5.LTV^CK5U@V3I)C?\ZX\IV+]6?c(1S:_>+a^ceJbg9PVA_?-I=^_Y
GOYW2H<\[,YNF;V8JfA)+2O0P,///A+[H\:3_ac3dW+-;[R4X1Pg=fVV_#27W<d7
XWfMCC,KQf1@[<^CO)O0>BO5&JGLUIe^XXMP[&O0),CA3\Y:(fIHO5<\KNIaQ+E+
/WZ:R#C+aI,F<F^<I9H/2\KYQ7f?[OY.X-_#-Y+9#=M(P8efe=]U-#g<GL10[OEF
J:G\))0g6c]Og,+4GN=..EIX.FU8A=Z5bJ7]C;+3)I@6DV)QB4]0BR1CDg;;2>_:
7WT9XQUM-f,\;<#FTRW,6AK1a)#O:KgB0c4YUPYdDYaHV0b>2(_KE6-fE1NSfec.
eN1bG,J:./O_>/=PAE\XXF7\Xd.0K;PGS6cM[2:-X1JEcSf7\GQN\eHb^@/R=8:A
T)C_Z#AVTT=B#(=E4e\R@Oc/GfR+\X^J\bgJTHF>IBMfSe30b,.?c.^UZX51\c<Q
/GWaIVHDTd)QS3CGc:)BELZ>50UQ5^4(I0YF:g^cPdL2U6K=@K]C^Y4]2,_K5.:U
DAbeE+8eF_Z\K>X5Qf;<(^ZWZJc2+Ha-4;)STTf3]@87<I88GI.6J)PS0##CN4fP
O_CEU)=&HZ?JM@MV)&Q;-@HK-9W>./>6;WXY>4TDb#-#a<6:M@4XB3:-_]a88Z>:
MT2J3R[,K5W>2OWY87b[H<QF,eLO9#gTa\g5S6>SQ6T]Q8W(R=HZB6Ba98+eb,cV
^HfB(2Y-/9\^Pd-_ICF.W\V]T,VC].g4IV4</g;H+]H(=.39T:b8B@fPJbP8VLN:
R)N27(5C35-?<b0YYbIMKC+9)c6VN\_N8#.Wf]abSK16;R?X1G28HYD74\8U?M)1
>KWgGAPB,J<P[S8E+D,(g;.R&8bdC)I57(cJPK]H,0IBXZ^_K:F[UDaG+P2CWKWg
3F2R?S#7_)<>AG<F36?6A5+4JSW2Ib-CATC/A:3E12(+0([6P?ANb^CAcFZ<&SI6
E:1O@(-EKWY]UIf+d@\<B4FPeS5<RQ.1W[g_+B8(+LRCSLMU/fAcgM2AOg#H:a^K
YE<_DT>eBH-1P9c=aE@BV8)W[C)5Z/Bg7IZH0)-2SYc>,Y\Q-5d1F)7MZ-QDX<BW
=5&GT@?^<5_^PD3PZ(#1f_17:SSJBP>E@\0I&VCe7V]@^,?T0#dEAFE-PHbT07_^
aYH3]>EAKJSW^+g53^f?O>6df.0cfXWPVE01f=fU8<<TTWgGX_CH)?-\?0d7fI@(
CM&9=)R)FIRQ4^L-RM4](^f910da]&N(<:PgYS:<?ZMB1NS/0Y-LM-NA2A]Y.;-0
RH:3IZZME4E86LJFcg;?g^>.-@H-^HbOR><JYcFHY(GK^MW5Q7,)WSFfZag]]SV_
+X.7&B=>P>e16I_X7acZH\0ULU3+BM:;Nf?FLT;#;)MadCUIfP\fBd0XO#8FU5Z:
=-W^)?85]J(,)-FRPKGMg.,=Y+>a\#8GQCCO-R:-AD)ZM6)S6:fK4341f>PYOgO3
V5;EQ[N^H:a)eG>eQ&I9ga?F1ZJYE6EDXK1[0QXf/Z19XXaL5=@IW5L0JK5Z@F))
QP,/GF=;XC^L.4HH,BRcW=,X18-EGgJ[\(1U&E-BO#T#(gAE6a86Q[3771X47TgO
G__2DF5/]K-0D;7AMB(P1Q3G-#+:HYV(W(P2)>/[<g\@K0ba-E2\Uc_2)_<S[8B=
02[Z:KdL@N.&g_]SB##(=b;[2OWT>_D3)bZ(4IO]J5+PM.Z2Y-K\CLgR&=[a^BW4
+Q]BJIJCgPX0D?+LSB\Ke+5>^FXdSW>\&Y^UNNe^=>U,<3<LX5O#fK4DPK?ge2#d
B]IITN1AAE_;PCeLXH1T>@IV_YS=_DMK#71#>Q6KCKY>2EaD?TbaR,L.6]..)CA]
?7ORQ:Mba1VY8T_/1c[\(ZI@OS>UC=I/g,SSY>gO2g\N>3I<A-H0FgB[L<]G^:F@
0MPHaCWIOE&1&)]##64ET^YdK_NBXXb)[gYf1&6WBccJG]^,(B9W;E?[GK)UAGS6
If+I]H+&8W1K=B.R_\UaA=R@[2]DH+g=D=(C=5L6PY^0a9G\8K>H-9OQ+N))-QZ2
^S8^4S2SFKgcB;S&S<]g_0(Mb(V5D^84GG63L^I2fDRM_36Ld7VV\66Qf-+@f]TV
SV@_K-X7cARL(@^g7VH2#9gbF+?L(@bL2MUESG.H&d)#d-/11TSEX@^=5e4EC=^H
\(^3g98H<S\7Bd&\#(^-aP#)\T&d;Fe:gc5S@(<W+JO#feBZM&I);24\,e,?O&HJ
[A\<BbB(0.FAB,d_F?aO<TQ3G0C3g+T>.-:[7704?f+P>dVTe9Z&1T[:;@MX]7_M
?gI_YA&WX8V/2603gJ\F;._?>Kc7+f(;N95<\((QfBHM(U]GI>&<6J-QO.^I;C[J
?&9:^7c+S8G01#=IEb<16)G@NL,F@LKP67(A^.)a^.?=EgZ<YfM=6+bVJV3F=?7Z
Ue0(Ed4^^S\cZ)A4=B/#aCS(0T(5.\1-UR#Z@fdK?TF/#ZSMeX1M6/<OUG2WbB2.
@c+B\)95(_B^,@^R1IPVe=1@B+3U9gEgVFN-@9beXV<L,Zg6[E///M(0/08B)J?Z
M=B]PR_GM;J9/:HM.4caN9F5AY,XaFTH_]&[+/2AG6-7FI#T>:,bYa#HdGGCKI#T
aWe)^RBR/D#.C@99EPGdBGGLF@57T?(B<J^EO-b1-^&&\eO-ZWUCRKaTX+4V0[->
KUVB)e3gDbb1O0=MgBba&FHUV]DXI?&/?HLK#,VE.W,[WMGZO@_&5De#25Q69>.e
A+4N8/XgALKFGTZVR19CV[6J2eOHYWa8P=5F)cXLJNV31Fe:2_AOI#<T<Y;XXL_2
dLE^/B:Y(Xc-E@RO:11NP?.QCf6B\cc[-RLZBX(P#;P8CE,3U-5c4UO.FBa;aJIE
?XQ0[42c&1g@<6M+19T3ZG8f[&Ag_-g_[A=Nc8ba8N8RK9>2FU<2/:aX9^1WKgZe
N[abGZA2f_D.WVRF,1/d=B-fM^EBHFc-:+X[cPB(8N/_3STHEDVN\4b/ZQ<W<]e,
Y,\#LIe4RYgQUVB>GRAKZ-,8GXe:+9MX5^K9QdaUQ.QZD<E][^E@a#0aMYbA_HI)
P5DaWN^B(WI&d8Z3?;cI_:]e-1P2PSSP60_Cb[?5PZbQWY3gXW]X\^?fgHB4/R_>
U^@M3:D:PZC&VZ28(H4BMeS3@NA\0/eQRML(g.HR)IgXOE[A?+RZIY([5Q0]&b-X
5[K61DVP5A\?@->BY<a6A==gXg&NG?])XYa5FO=Q12U3:=(Ve9Y<C?8^;e9T_>d?
MQM-W=(X0Q?cgadgFPC6N:NAgA;b>.Q9T,3UQeW]71Cae>+-<;_U@+&fL8E\Wa\\
geS.UC5:Q+\]PKN.e^NX)UN1ED:4_A0JNE::XUfDQKM^PKZWgY&[)XVgAU)H>]IG
N#EY5E)1B.++HB12DD7b.@5FgV9LF:^DU\^f15E=[d[A;LCY[DVQ:NX9#R&OQgWJ
-ON2&#H>@-?2PC4H[;A):_?W8]<HcJc>VP>X2W=f)4HPc8L(edXXfe0SO;?+QMaQ
_8TPXRM[1F-2=6R]6[f0bR#N@Jg-[B(5>7JQU03TJ8:?QOAZ^aN,4E&cNWK8SE-5
KUU_JILF^3BdYC-Z6bYf9O&EedSI1P;E?_2/1<D=11<-39EAR@H1QI8RfD.BYgA@
V^@)TVI7?4ZcHEdI_e1aJ=-F=PDf8HO@/0:1_f,,gKf1E/U7WPZIDc\gK@2S>PS5
I5e,6OB_#+\FN5OHN?V3<.5MFA:27d#DS545/.VQDB48f4?PRLDH1#JGFa_0ULLd
29#UA4#51eGe.OWDT_U4,g@VK96_dU)a.Vf64Og:Q69ISNg+D:XA9X>?[:A7BI]X
aC=^Df<>_9_C4H7JE]<;EVCYdV2\>LA=:-;C)M#>W.^,&b6416Q3VW\dbcKeAJ3C
U9T)&?/B]2IfQ[Q)<&U,c>VBF1]01caNFeMPGfOC3;T/DZRRN^(5845N9[0;C/W)
g@5KDS&Kc:3]V_Bc7;eA8N@:QG:80\bSUQM-S\U?(>(5=g1d;R?LEM#Z<PS23<b&
ba;KQFW8Z9WLHN5aVRZ70@eO8_QLQ)=cWUBDQ(<R5a+&:-:2Oa&ec7\JL/MJ+4+e
DU1VaeX]^3P\72J\_\CfVBEF)+-20Xf&FeX?U=@[2P<5beE?<I;M4.[=Rb&5JI-S
(2IJEZ_0+<^6HFWOUdgOL3_E2ZB+g:4Dg^<W+MbHJ8>+,]H<(Bg/?]Se>)=YA[F\
Tg5YLIM>b<?\\?\;;H[C##T7J>[.^Y^7\>aIMIZMJP4>ZPTK/9&LTOTb5(TSXLC@
f=.Z_IbICUGa5#WSYR=1SJW^ON@?&D/Nf()BgLUI;93\S[5P3BR+MQ6BNFD4M,#@
I4FF[g.L&F6GGX6;93I6GJKIY:5H6P3[/;4,]BUMFQ//0N0FDgR)]B@03SEcDE^8
,H=eP,NS5G^-/DgM-@@;#G668J61SJQN>e+(SW2QJ7AeYA4S,B?H?O=S72[WSP8\
db52J=Kd/Y\7GG)F4)]5J;;d5@IHK383M2SF>^QY#ZPFe,,7TXMTc1_+If0;CXH-
[F0+^;2Q._R<;[1R+M]0+8fN8eARXO3K?J1YS,)=9V2+d[&gEKKZ(5aCJE,N9ZE1
O.=3aCa.BB[\eL71+X>.-d#KZ6_J5;V,FF4S)DQH[>HASX-QAc1?KD^3U4IZKO40
c[F8W4XJOSIC)3>I>/KW0U;e<AYIWa+>5JEKd\E2?Z2]Y3JddZO<8LSLCPE#.D#4
K6/8[&1E@W4O8ZBYcO-RVDaEAB4)B)JHSTd[EM-=;6-IO/8F#PS<LA+fe=)(,16X
H&6DIgSc\@_G\PQ(PCRF8M[VRVBd-LE\8g>C2Q3#Xe.8S-Ue=D84(S7(<c>\CJ?T
)0C4ag0^+Y&/)5CU,?MA9O:=]5WKET?DMb-^PMY+L-/@3Q?5N?>HY7C181HTb@0Q
HNa;DAB[.3]-.ZHHEN7F&QVGD96Q.@Ga]SLgN]\f,AbbWU)L9&U3D/^OX9PI1CYM
bA[=-A2D->bDbVf\@=M+E88-809H[(,YH.cCIOS4=<])#+&]^f\^Q<cRTfMY]Y\&
Z5]&>GSI)V^FT>X;TAB8_FLJIc62+30&&D,Y=1aW1C/Z0NI^KY.CZCA/e8([AOc3
P[P2KcdAMKZ.P]>L]=NLYBN5X]a/c^V9A4bRe)eXdOXMWCEc4][b2@N)II#HbXgD
dP>DP-4\_Q&@@Lb6?//d.#bB9)Fd_cYMD.]52>+bdfZ__1TVJ1=XC;E0/>5c/1LI
Vc+(76Dc1[&L,.BHRVJe5ffe=8<-)^9<<2#B9.S>T67=Z6220^5DEH+5B\@_d))g
gSH)a\WS:K-EfOBdHXAa-P?6]-7F2_b2.-J,65/gDL-F_AJ@a1LDBbCg8HBI<V,Q
HSZ1b.77g[\.FTNGe8L4UbZc>+C]<bBY3[7AMN+]\/W]SI<5998G&P-GHbY8PJ/2
Y?(NU(a9:P95bd.0V[_.:@1L.+BcXLQ^5YDCf4P:>G\&,Yf7(30ZZQ^\bI(5L1?1
)e#N7?a#KRc>I4MT1Ke(ed6PBI=C\R-c/+&c/GMK3?fY?EF?SKS4[X@VW?I,J0^K
g?=?)P@M0(5T7IaZ.f+AFD-BeMbIaNJJFg9eS5,X8/HX,[&2dA;DW5=+JJc@+B=F
U4;HAA3a.EY.+;f^(7TF.13=:>6@/^K-+DZeI5eM6?_5EfP<<?6.e+^TP+XR4[_(
A.IecZJT9.S(I+W)6FLI1_4:e>@3YR;:0S?6+]@I>V]<^:La&UYLQfLZU4#e0#X6
L^,GKA9bJ=L<(LTRHg_T2:J=dfK3C7V[5(bK8EWX>f:ED<[?7W;2UEZ8RcFe)aEV
(V/g3&b,>d5^b#4COA^+aS.3/Y(X+N0Z:@F;X<5@I?<9HB5FFGK:BR^Ve:d^(d[\
C&5HYX@fCfKB[/FcI&WU(EPX4UC4@UQ4R1#^E_Cb]SSQS/[&T>6UJdJH^AR4STSP
FYa_B+G1,\(3F5#cH:-:)V)<3=1EG_cCGK(a284.eYSbERXS:O(?aTUW&c]VDXE?
CLJXd(G>[#9V?4<@TPA=N6fK8MMg>SO5B[AW:eFIId906fABC<CTUg<5D9Z/GHD2
2Wd=0b?PHK\@V:O.e[:>ISL/FC64BZ^FQ^FC++BJ=g.\N(5)bVKcT,)fQ[+)#C@1
,^Q\/+<DD^,?68a(BUFeZ#+/7b,+)5bcVCU7:NY?/44WIIC1.9,E4O]\1-@4[&YW
9f_YcZ?<>+VK@e4SFgZW8.3)?LQ+_O&)MK@82K()R8=AcgN4(GMCPRKS>TB;QK3e
8.<Fe=8Hg;OB&-NSTd_>5U(<.YM?C4+GWaSDCdB]T9M1a8,14AW#1F4a_J55bfA+
)eJTF@=c\QgK^Wg,&ZPb1=+EF7PdSD48[\_1GR2_GCA\\UDG?DQMcKY4;g_\52)f
[2@NR/@(P#I((L/D(^MA_3K2>LF@S5^Yd7U;27HK<B;34e4I,SI/O74d9e_3(\L9
HD:^=.d4M\+0--=&(gV)d3E&b5ZTHFfSR,31\ZN8,Ia1N:][eVJ>-9TO5?e<NR(&
.F^dM4VSX1e1\0AWGY+de/abU#Xg8KB^5SD,MQHO5AAdY+W+)AgW>d[e9F,)8FD0
F1C.X[PG8S3RX)Vf24Cee<S[T.8W+.e/S.d/K&7/<C):dE2-FCY,b,e;2>T8\RV/
;\;M0_)\gE^J>MNWFD5(P,EW^/;3a9DaMbI:GNDY>^Q^@S2WSG@]X>1ZPXDOM>;E
XTN+<X5)JYg>,R/E:.C5W&1deZWCd^@1-=IN<d=^B@cXO+<d,e?UA7F,U2R26^^#
,34S/LIb+(T3\#SA.F<1PgFD+@J@I1DKKgf0A,gDV?2,;5I?JY86(]1KBSC&F.La
BMU^9\f:G>>XX#0OP.FMKEL1e&E6=H6cgY[3Z4YXc=F[3Rc/5O[922gKSR>H8U1a
fA(W]f4E^>c,8YU?G-^cU=V=P,1SfT;cGA^+N+,;_,)O5BK93YZgY/UHER#Ag-Oa
P=@1V]XXcZOH-=CfADd/e:RLT8,,:Kf7UEV+M^M9MR,>gMCHYU?P/^?9<G5L(f)b
FGIaP]a)KAI1E],b_,TJOCZI;](9\YMZ._^:Uea)AC0A^6<T;E\\T2,16&^,E[3+
0<6N#6bM+UKeA8H;JD-MPg#XEZdF]+(c-,)=]>NOTA9P(\@1;bfU?dY]:0Vg:(Rc
QE4A=T=eN[\bV8@>AN\GC)Xa+,D:S<BU=Nf(:/VSC-:7R#V4=+CH::F5d@Q(eNHX
,5#FD^TS,EZ^4QS-&HVF2(<.ec>_?==49<D@LO?TZ+_)5g4(3bLAM#8Yg6?\O&N3
4e\S_G[QMX.)#_4R50)8K\0B/UNM,[2,.4)933(d7QF>)7Z3X]_VY&MfR&YMCZ+U
K\,D8[dN\O8WSI<]0_V1Q>cSBfg;V19geEEGQNbaP#<IQ20ZacZ?+237e@g0:Y<Y
MdMd9OJ\gbbG^6c:2,d>/QTd]<QM2L0.We6J@Ff7T<T+)1Z)0cOR2SB7a,Uc8+Z(
UP^@2YV,P.E]K0WOcKJd5W/dLF7TEUb_6;K]G5N/D5gXH.0A(7gc@,[<Z#=MX8+F
a[UOe(UWge0YLY7>eQd:bPOV(,Q4R?N;)4@3P<L8FQX5cD;Z_23=](=8U]_3J_@U
>/b0OO9-5C62.HO)UF\13XM?-0]N_age;[aWfL#Y.=RM\a[EUE:M7bXB/]dAG&<f
H?26RD1;R^gOOCYI0UfBP0KND(c39?e2J]2:[34-.1@&4gYYYI:O/WeM=HbeA=96
HA]H\:R=+d-JV#B2M52#dBU^CSXc8>=K^0[>?@ZK4fTB82]8=9.:1PBF\(a36:)=
-bF#g8\McTELH<UD<@375ZC1LY13XC5W>[=caX\SG:FUXO+.b)Ig&O6J4?@)R5)7
OQ+4/9<GX+O)@K\VMK#\6C^L-Z(:,<:]Z0\/#gbB\_6Fe=&fT,CP3&2WP&JM,[C-
M-CXfMeBb2I@b4AeCG]D<85X]<7:(J#L?V9//O>I9C+==LcgV,K2gC(^JAU9U.MB
:\;&I]R66?L1Se)J:_T[<-?bcEB_]XWSg#.>XNZ=b><V]a=^3b33_#^?<#Rc#)>B
,JY4PN&4V^&6[5?Z\_8GN>/=I6f[T&aWT::MBDd3ZXe.LW2N\F[Q:=TTMU&-a&3c
ZSDPTcZ:0Q)8(V/dZe3[<FV/,,JL5Qf#?U?LKOW^LAJc[Be:E^8GMW?W-_BIUP@,
@0=@_:1@_(V8)H80PB)b4Y3AR-.LF5@DHO3^+<4?3d-f4SCaZgBT@Ye1W;7?_eFR
eAC0)F8Y3D<]U7d]:(?GYNc[7Q+Yc.GDg\N+C+FHG1M0Oc+;;e,DU/QUO^TUW+d1
WFDUc03.76T4&PB==a4B(aa@L1J699K-U;?@Edb2XLbB1/?(BTHd/O&,]_,ZcV50
cGK+#H3K(OKI[Z7MDGN6Zc63_OIK:OLA\_3Ie\I&bc,/_DM,@b?V(A<YR+3=4c#Y
N+#6;HQ>,0[CDe4^3Q.U:53NQFdLZAL)eJ/(5Q5f/Q/PSdMC=QYDa@#?0-DKJC=:
DY.FOJbC)SeO^J-UF9;\a#gA1<N#a]YPTe4;W&F<6455ZDRO[5J30g=UUW2O,#T8
&-0f)[7XfG6Zb6e40O>+#L>+;)B?Yf,-IQb9-]YA+=ULI7U[(=B_&ba_)9O(Q4G#
AH9<e&#V:>9OJ_A&EVTWOO;gVWZ#fQZ;SCRP+]b_H#&X5B2L[\7ZP=P@>9HU/LKP
/d).8[#R;PJX(?_BbQ/5BPSX3Vd[MJbMC0ed,YHfQf.#Z=1-Ed5R1-f>2[5T#[<P
-UICQN0NG;O.-3a)R=#ZAc7>-5-5beD1F+R,<eY^e_?W3C#;FGZ\9Fcf/W#gFF:B
/R?-3=76cZU?CaE9J4\.:J+@=(KT1gMOSUWRNdWX60BNRaFIJ2^D,V>ASFSa:MUN
N6VC:MAM)KGS]P&.XY:cB6;a&UTR6HZEW9&<KDd;0W+-IMR.Zd2(>P)6)O#CdgKT
>I?12.=d;6B\<]D@]8?F1AcV9c-R(3:a+,/,W=0H23@,CVcYdQEc72gNbO#(BMC?
2cSMPK,TAT+LOK(f^65>N^9#L;d,@(^KgT&CS?_TE3Tc@:PF3INNRN[<.;4WB[,R
0)QDTbScKa0\RT;9Y,&[>WR21GHTVcb>K05>XM;G8S8/OP#d^X/Y-8/OfXdFd?Nf
E)SHZ75LA(66JM(.a=^4TIg.X[Y6[)3;5U_+]Q+K:CEaa(0Y14g:]5(9[gO/?JBa
4b-g56Bf[Y4XY&XdeK[_.)@+fTO,[+0:^_\06?@PG9a[<&\XLa6Qb7[B/;2-B57\
5W/P4WX+Q\+M]K,?QI6dM_UXKC38V,2eCKb+5FS[\eBU?\^IAKP#87^KeV[&OYL5
Q2#55I_IHUA1#a=Gf9\^KOD8[PbG((c2?#\>@]@P?Aa.UDB^LBOXL1K09eU91-=2
GbLB]H.LHVgTUK/;/Q?,<2JYfZU[BJIIRS,NYN55U_O@BGFK<]Y?)INF]U]C3742
+PcUJN#,MIX>_\>KHAG_e>5LV,.WL3<9?eWN1c<+4&N?8G)eBU?EQb-=BeS2I.O/
E,)KEEGIDJ;)0W,M2U^AB&UUO+.\eMa<]PVY?WUKP7b()c6;B/>Hbc&MSV9PgKDS
.@MD@3Ag2\<(4cg&.LcX)V8Y&S?\->E@QK>Q)TC^X1]JI1g>::VZ0.8_RJAI/2R4
\?JMLT9YZ8.5<<)bT=PB#G_4XUJRCL5-g2KZ9A]D=G.>OfA7ZB&BV5V@CP,QBdGe
fC:RSHM:fSRUT0,b\b?)?E3D9Z\Va>dg^^S:KPKN[V8N/+EgH4\Ca1]S9LD-7]:#
Ug=Rg^D-&W[^D21N-JcOTD-RAB4X8OJ-#6YB/+9LS2f1:YW4(WGY[-_&He)SHP1D
ORBH<K0;Q&GM?YTN@dEdN,]R#e?]=,BCP\A;_BY/B8Q3C/Mcb\cb/HXQIab923?Q
LORF3Z273Z/fG0&e-<5=X&[^66>NB[+RWg#U97W?a<B3cMC/bWFCSe7<gML;S)_V
.K^IE69.2G4.]ROgL5>bgHB+&GGf\;g,</ObZ;efe6K_NT_BBT0fT:KTTTf>3K3X
YdGb.,Y2A4.7DPZEEaCHH77@9]<g#UfIFN+b\aZ\c3J9/&D[Y2(#&K08S+\0NH:Y
MMX6Z]Se@bIJVKTd4,M;.b?JUdFWeRU99cJ<U0@1ba(:59Ef+fc[V42L7D=Ia-d8
5g=1Z7Z+?28;dD)H0.U0;#:DC0]aUI]6d0c^SZZU]DYI(e;159U@EY<C]^Y3,(^&
&DMCH??JO<BYQV@Z-M&^/CZ.eOfK5&E?OefVJ_0T6eM2-f[5D7-H>0]^75KHB4fU
_Yf.VME-PY__Mg02U(&C)9Xg0=G;Je/d[KUb0^(KG1.NRWeCOZKacBNQ0;a2W5e1
S&d2L#>.db(ASHH)a19(AFT;I.HUb8I^GJRA^D&6+[5>QaKe4b:_3U39-#Y];09\
2LEQ-KQ+1)e8,.I2T\(,/<4WYSAAS;CXB0K>a+Q0a/V7#Y1T78cM:9&@7OB;.2c4
gg+;XKHH,HE#(T8[/Wd\c;FX6Cg/VD4a8(1>QG4)4<-Ac,+#LOW3gA__-\G2S3H_
T>/()ed;J_+EB>Zgc,^L+aL+,?Ca[MRA&YRRZ/V(2_>.XK+#=)D+I?^GOfFKSf;/
6X=W,YLRJc?QJ:P/CYI\>.XU//>7,:WUbe3AfN\EP@_UMJ^U#.14g;5TE-e_V58N
79SE##J9[+1LHBI?L7+cQ0F.,eg=FUK^f&dI9O6V(aN@-12#R/VYPU)9JP\/=U\>
,_Gb9F##_EbHB8d8I_A6Jb7?gPg8Wf19d.OZA]M[LeJbY7TF>8(P][]+dR<SC]23
NZPC(-b^L(dW\Wf@eQ>R7/eL(8CGC=]e)9XM<<#BTM1YAGb)f+Bc(d)QNYTYK;_(
gSbH<6_a)eNKcA[R_=-EaIbAKY4NXEN&B;_10915Q&E<4X?YV@Y>?3N3?\5@/((T
=.MV5X:8,gDS)6^dY@+:9<M)\c9;4Zd8Q9SKVHR9XZ3+?1JFFR@fB>GM;__c)@C_
S<QUY]F#d9N#45FU+Z3fD)g(?P=:C4CfH;AA,T_R4:1^LI^.bZ;5MNBYP?bfVNQ[
Xc>PKIHW0RDI?67Y]>e7fU>1acZ?C^=Xb.?PU]P(D[#L.Lfe?a;g4YbQg4VU=S6U
c1[T[Z-(Z1C=B9gE\Pg/SLL&Y-0_Xd7W6^PMQcD-,W6NEZ;QfL0D@WBd_D[_f#.6
BYSUJ.gW(0>X-76Z:2d.K^G@[F[)D]KdGWFCKPP#Of18&<3OI@Q?U=-B:([&aa_]
4J<)ZY(b(@cd?^K)T3cb#[#ZC\R;YF7TS>J0W:/_61c?d0K_[6G2=_;227]/2bTA
V;6CR</eF?>&00\XLD,47+0YCT^+fRO8ZdANR,6Jb4bJ^^M;e,Ua-b-K-^LaBF<J
[59Kc(<9gEVZ@R_#EdL><c-?[TBD<1?CS[7FHX;e7H=MI4O^C5FH:Q_f;FXA:(^#
7MC>^.T-c@WSaPB)=8@-/bcIfX9/a(=1F])c+7+]Ra3EW?A\+JMAg-WReeRKR;2+
J\NR/8b978W;;G@-V(5:HJ<9JPJg?]#P&N>7WU(WGW\Z6R.&/(6#SICYF.<e1+T^
)#TQB#0&0?(U/&?:6QP]Deb;c;)R9UbYQH1-5T-[#I340V.GSRI?+CN3-U[4:8:0
9<GUU<.Ub58M_TbMQD)@FQ7BDcM5ZIZMZIR-dH[BG12P54,28,5Zf1,F4geWdfM0
bc^K1;)eYK1QNF]KXdLJ^KSQ>B]RYb,,-fbd#;-ABV@Ad6f,0\BS3ZEPU27)Z&<;
YA>9X4/fG(G.NG6Sd&?62CS[QO5QFSCS1N,/-<cdFAD;DH),4c^ab1[b:AM4aS_g
P@(G59QOXBKI48,,<,(/#X4]BK0Q&D7P?Sf3Jg=F)>EM)NfF+e]HKPMN<#N92Y5G
)U:_\5O<H.bcHHI-GXb6c.T2ER949:_<Uf:-2/&f\#(4T=UFSS1187EYIaW7bJ?1
c=?1C71G,TJ1JLbKCI@Rg>>-XR2=2)GSB#N4ZGcNU/)PgSYHDEM@SgL\?#MgE(41
3LT8QQd0J^?:I?A[YZ=g);B9_YSNBLAT/UU/K&a#Z@L?aTXgaXK\+/&&<2^g.KR#
UW5[\PJ)bL#[0^<>0ccP2JJ2@2DQK)K+/DDT5S+9\WRHeg;0\Yf;\D^95R@F/:(V
dMEgMN7@JK;d,cQT,,,XI1@G3@c+;Z?04/CA7bV0/FF>.-e+X])F0YZ7KKAXIW/L
K6[bFbW&Ec7cQKLFT,<?)R2OFMa#(&;W_)U636e?^KRDA/F^W/4/2T/:Ae9.[XH0
ePS9:<5)&bIPIAcMA_c.F-P)W7YSa+d<>(+:6@T1A>RM2[-GDcM(I<LQ-TY2ObLE
7EUN2.;3e?\S/7.Q4e.V8a2I)1).8>dL\U^B_DOFfAJ<\fgWcHdAQ^]MR(a[Sg;R
;#NW\<CO-LeTD4MG<QD3f)5A44OLZ]Y?c)=bE6a4Z^0^UASAA#d07J(M1JD,]PWV
-J+H@C;D0\eE]:.#QDc59a2D-UCfGc4f<e(??/-aN&c@OL^ZT=fgBO?+.<+?_CNP
,(e[(gQV2M8(PaQ+e0b8O.O.6J>_+ICKHY6->4BNW;H]^fR_MJ.OAMTF?SgJ5M=:
R8Z2:-9,:JE37,AGZ?N#WLc:X<IH_5V)D_f9HT]7_6dDLe&KYgAB@([7CaH]/]g2
-G<ae119,S8:A/)c_:M[K#U?eL5Gb9/MGZ7]Vdb+F22_R<I<.be39?^>eS-X_N+4
_.<f=G.+-HB:1\:KERf(1IKC):9@NC0GV:Z#O0@L(P4f#]/RQ7-dHF?;&34F67>)
95>/F;;=/MIdf<5A]BG]:F?GOK;+]b6R-7&dgc.VK:/f7TgD+3@-9b_I^2PK]ESE
>@YGZ<;4PMF5K7;1WdP0<a+Ng0aQgN_Y)a-3dWag@VAg7@gWW9B>Q4K7c814+]0;
SH5/Xf.RZ_?LJG=@H)]UT\:DAe?P-I^+ABVU#?(R]cQIIe8<b#7<=CaA[U0/FHBR
/=,6>U-g1(\Y\@dJ](+H23>gEN\=59f,Hea(.5UV3c[=TL)5WPT4AQC2d1AcKSN?
-3Fg<7_@48]J5K-:FIGIa)<aMC&W9J4?F;_:]>A<]2R2f(MT9C[Z8X\Lb\(VYC=a
#[>[]BgK_:TXE(EX<CcOAE-c/Zc,@@Mca^=M.4e<&C6e_aT.;G3])66]^J+4FcfD
\V:DJ6H6P\LBA+<GFg)W>(EHff-5E.M^ZXOG46,>g(Xb\gV+LE:>QWcW^]F[Aa;T
eNJ)EV]TUIRTbId?)S:>0^M>=4.FHcM[]7C/?QSV4?>O8(9S0:c;3WCe2(]?TN:N
TSZIL?:^O]A,X>]^(eU/P0KSH09HGOTZ=/6[eX1=>6D@1K(/GXa,QNNXU7W0[fJC
?<_]FO4K91@Yg=b]bb@<05+5XLM/W(BD>?=bHI9LOXZ2@OWZL#[:N@\:1-#9&/0F
fXe#Q4ae=2IBKD55E-1H3Rg(gN>Z;KUF]T1T&KDVHIUC&[2(9Y\+(R,.fMJN(eC^
e6DXPI>N_c7+c:DeKD;aG59C]?9IdIU(:K+5G0#AgG:\W9QIQ=F(\Ef[LC(&+/ON
^P2^VO>P];f?63R2@KeDc_M.\>b1K&(MX4_EWSbZR;M@#3>H\=A?-\>V#N1JFWSK
KF4U&^XC^/g2:\e86CPYZ2<PFJ-73TBg4#+W(QSN/8.O2=.6N0D\7+9X[-fCgXf1
G8QX]NZ.XH,EV--R:PE)eR)XVQ?F^P5,HGV41.(7:e4EZNfG5gF59U(MD5P(cAU7
#IGFZE=26[?RAQJ0eN_.?Z-1Cb:EM4J3C95eaYUW^V?P:TNZ:4_I^d/@@@>aCgAI
gS<+7,Jb<GRORI;7Ob#NT]\\5Z9\-EGLE=e=T-X((H@<([DGZ@VO/[YR><BU91P3
8T?XZA;#8PSXO_TfML)P_.,38cA/bc1V#GDFdCE&gIHg9D.8+EgH_@YRP$
`endprotected


`endif










