
`ifndef GUARD_SVT_AHB_SLAVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_COMMON_SV

`ifndef DESIGNWARE_INCDIR
  `include "svt_event_util.svi"
`endif
`include "svt_ahb_defines.svi"

/** @cond PRIVATE */
typedef class svt_ahb_slave_monitor;
typedef class svt_ahb_slave;
`ifdef SVT_VMM_TECHNOLOGY
typedef class svt_ahb_slave_group;
`else
typedef class svt_ahb_slave_agent;
`endif

`define SVT_AHB_SLAVE_COMMON_SETUP_REBUILD_XACT(curr_xact,hmaster) \
  svt_ahb_slave_transaction new_xact = new(); \
  rebuild_tracking_xact[hmaster] = curr_xact; \
`ifdef SVT_VMM_TECHNOLOGY \
  curr_xact.copy(new_xact); \
`else \
  new_xact.copy(curr_xact); \
`endif \
  new_xact.cfg = curr_xact.cfg; \
  rebuild_tracking_xact[hmaster].is_trace_enabled = 1; \
  rebuild_tracking_xact[hmaster].store_trace(curr_xact); \
  curr_xact = new_xact;

class svt_ahb_slave_common#(type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                            type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_common;

  // ***************************************************************************
  // TYPE DEFINITIONS FOR THIS CLASS
  // ***************************************************************************

  // ****************************************************************************

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  svt_ahb_slave_monitor slave_monitor;

  /** Analysis port makes observed tranactions available to the user */
  // Shifted this from base common to slave common parameterized with slave monitor, slave transaction.
  // For UVM, it is available in the base class ahb_common.  
`ifdef SVT_VMM_TECHNOLOGY
  vmm_tlm_analysis_port#(svt_ahb_slave_monitor, svt_ahb_slave_transaction) item_observed_port;
`endif


  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Slave VIP modport */
  protected MONITOR_MP monitor_mp;
  protected DEBUG_MP debug_mp;

  /** Reference to the system configuration */
  protected svt_ahb_slave_configuration cfg;

  /** Reference to the active beat transaction */
  protected svt_ahb_slave_transaction active_xact;

  /** Reference to the current active transaction */
  protected svt_ahb_slave_transaction tracking_xact;

  /** Current beat number */
  protected int current_beat = 0;

  /** Array of current active split/retry/ebt transactions */
  protected svt_ahb_slave_transaction rebuild_tracking_xact[`SVT_AHB_MAX_NUM_MASTERS];

  /** Reference to the current master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] current_hmaster;

  /** Reference to the current retry master driving transaction */
  protected bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] retry_hmaster;

  /**
   * Current and previus value of HREADY driven by the slave.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected bit current_hready;
  protected bit previous_hready;

  /**
   * Current hready_in signal value
   */
  protected bit current_hready_in;

  /**
   * Used to track previous burst_type for error detection.  The extended active
   * and passive common files use this to take appropriate action.
   */
  protected svt_ahb_transaction::burst_type_enum previous_burst_type;

  /**
   * Flag indicating status of tracking transaction.
   */
  protected bit active_tracking_xact = 0;

  /**
   * Keep track of number of transactions since last reset.
   */
  protected int transaction_count = 0;
    
  /** To track if the hunalign value is changed in middle of a transfer */
  bit initial_hunalign_value;

  /**
   * Keep track of the addresses seen on the HADDR bus; Used for protocol checking.
   */
  protected bit [`SVT_AHB_MAX_ADDR_WIDTH-1:0] previous_addr;

  /**
   * Keep track of the HTRANS; Used for protocol checking.
   */
  protected svt_ahb_transaction::trans_type_enum previous_trans_type;

  /**
   * Flag indicating if we are just comming out of reset.
   */
  protected bit first_xact_after_reset = 1;

  /**
   * Event used to trigger passive monitor signaling that a new beat has
   * been detcted.
   */
  protected event new_active_xact;
  
  /**
   * Event used for handshaking between common and passive common to
   * inidicate common code that current_hready has been updated by the
   * passive common.
   */
  protected event sampled_current_hready;
  
  protected bit   wait_for_passive_common = 0;

  /**
   * Flag indicating if this is an active or passive component.
   */
  protected bit passive_mode = 0;

  /**
   * Indicate the last transaction start time.
   */
  protected time last_xact_start_time;

  /** 
   * Flag that indicates if hready is sampled for the first time.
   * This helps to figure out if sampled_current_hready is getting
   * unblocked multiple times in a given clock. <br>
   * Used in passive mode.
   */
  protected bit is_hready_first_sampling = 1;

  /**
   * Internal flag to know wait_state_timeout is in progress to avoid it be called for every clock 
   */
  protected bit wait_state_timeout_in_progress = 0;

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked previously. <br>
   * Used in passive mode.
   */
  protected realtime prev_hready_sample_time = 0; 

  /**
   * Variable that holds the time stamp when sampled_current_hready
   * event is unblocked currently. <br>
   * Used in passive mode.
   */
  protected realtime curr_hready_sample_time = 0;

  /** Indicates if beat_started_cb is called */
  protected bit beat_cb_flag;

  /** This flag is used to control the delay insertion in reset phase and main
   *  method for VMM while processing the initial reset. The value will be 0 in 
   *  reset_ph to bypass a clock cycle delay and in main method it will be 1 allowing 
   *  the delay insertion.
   */
  bit reset_delay_flag =0;
  
`ifdef SVT_VMM_TECHNOLOGY  
  /** This is required for VMM where monitor needs to know when the driver is
   *  ready to drive next transaction.
   *  This comes into picture only in active mode, however, the slave monitor
   *  has a handle to slave_common. So this member is added here.
   */
  event          beat_level_transaction_done;
`endif
  
  //vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
qnHFAP7zdZeR2a9/Jm5f4a+9f7VoK6+Rj1iicoRuR1ZVWd9XIjQHV96Twd7ewDaa
g+0hs7M1+BYyCJ2AriD/ryDiOsl698BrH/Qk5UaWLV4LY2IQq9kXKGm2Li5TvV8a
na877i6mYTPZ2Ww5KR2dzqOzGt707IqptLaeYPb5OlbztOpcKg3aGA==
//pragma protect end_key_block
//pragma protect digest_block
4nZUon6eaiapAYYH+HOkVh2fVA4=
//pragma protect end_digest_block
//pragma protect data_block
ABhH1TgRwTiKj1k/teHvvvPYPg7YNpIcqbV7BCSMMiDOmZDRnpP4FzdyEyXc3RXE
mt4oTpIB9X3uGfHPdjaPoNgGkg47XbpcpX4Mg3XQvYfy90SjXjjfJLqaldxu2AWS
VFgZZgk93j8vTmmScRW2NLGqynp7/lKwPVGYz5cicsF2mCDl3PptgdJZx1RSI6j1
G/ACdHibzbYIYET4u0iHVj6YK6e8ZMUUwiC5z0cRWcp7HRD58jknOS6m+THmZefY
+sdE4dez10rWMrVcTSfpoqlW8x9CCV1RlE9HA5iNyTN+9uhjXVkeewuvXUAXSWYx
bUuyA4AdFtyxvznKTM+kWWVXigbMJezzKmjavt6JUAOBhbJcUsAgM0m+9q6BSc14
FVbBJdf5cWINPFebS+EnJLXE38p/rJGC0ZBYzj1ksytGRNrqgTP4TSX2d/z01cCf
WXANV4ZXFMTYgfakvZnYGvRpnhoglzIO7hnm1mAygpxAa4SZIWzGMkehEx8R7cEt
Ii2bl/WzmCqnlzGnAk57xg7g4kP5/OLAvd55/XP/ZMT5QtsD1JMjptbGmyQ1ZgnY
cNNm6GuFFhqbmF67wunqRf0fCr+lb2Cc/JmsY3mKy/yI1BmfuENGMbRYW07/U7RE
Yxbe3PUHP/JjTvEzrv7wad3VMLIZSlIhCu7dWoBX6/GIXx8veP7xX+eM32PbBSiW
HH8MT70mba51OXB/zU8SEcT2mJ5H6pGbgg5gIXA6uWlxgLK7Djnewh0V85EeJiod
bIsiI3veuATUaY/7DH6u2E6wWpJTHbzNHasmFd9KQLpCFSzsqaS+EAOYIETwK4wO
HRMDlnYYG5NUTSjFDx0LzGzXqS1jq1BBlNW3pdpg8vrzTEPIz5QJH/gp1lkAG22E
O0b2fmiorN0AWyhUcN9tKrmQ6BcBqnETQIuq68CQh8MW5xoq70e25KA3BseloYSX
ckPknAfxmn0iE7tMyZXgBAuUXYHTwIKpVetC2V/wuR26mLfjSiL8/TzeeAbYD9bP
JjBvldSLgRSq5vCgAoyDgcJU6f2vjWjK6nTcnGHjCyTDbmrMa1LsZ95nMVHpbLop

//pragma protect end_data_block
//pragma protect digest_block
0Zu417GD9VhmKcOLw1Bpt6Itp20=
//pragma protect end_digest_block
//pragma protect end_protected
  // ****************************************************************************
  // TIMERS
  // ****************************************************************************

  /** Creates the wait state timer */
  extern virtual function svt_timer create_wait_state_timer();

  /** Tracks wait state */
  extern virtual task track_wait_state_timeout();

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************

`ifdef SVT_VMM_TECHNOLOGY
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   * 
   * @param xactor transactor instance
   */
  extern function new (svt_ahb_slave_configuration cfg, svt_xactor xactor);
`else
  /**
   * CONSTRUCTOR: Create a new transactor instance, passing the appropriate argument
   * values to the <b>svt_xactor</b> parent class.
   * 
   * @param cfg Required argument used to set (copy data into) cfg.
   *
   * @param reporter report object used for messaging
   */
  extern function new (svt_ahb_slave_configuration cfg, `SVT_XVM(report_object) reporter);
`endif

  /** Called when a new configuration is applied to the VIP */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** Samples signals and does signal level checks */
  extern virtual task sample();

  /** Monitor the reset signal */
  extern virtual task sample_reset_signal();

  /** Samples the reset signal */
  extern virtual task sample_reset();

  /**Performs checks related to reset and update variables*/
  extern virtual task process_initial_reset();

  /** Triggers an event when the clock edge is detected */
  extern virtual task synchronize_to_hclk();
  
  /** Monitor the signals which signify a new request */
  extern virtual task sample_common_phase_signals();

  /** Returns a partially completed transaction with request information */
  extern virtual task wait_for_request(output svt_ahb_slave_transaction xact);

  /** Check if a rebuilt transaction is complete */
  extern virtual function bit check_rebuild_complete(svt_ahb_slave_transaction xact);

  /** Monitor the end of transactions to drive the observed port */
  extern virtual task complete_transaction(bit[(`SVT_AHB_HMASTER_PORT_WIDTH-1):0] hmaster);

  /** Checks to see if a new address phase has been started. */
  extern task check_address_phase();

  /** Writes data into a slave memory */
  extern virtual task write_data_to_mem(svt_ahb_slave_transaction xact);

  /** Virtual task to drive hrdata when busy is seen */
  extern virtual task  drive_hrdata_during_busy();

  //***************************************************************

endclass
/** @endcond */

// -----------------------------------------------------------------------------
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ZiBaEFwVL5w14lY6FO4r2bstrlK1T/n68+PkpNoQ6eTqKIHSwJdYAKer5QXP64zP
RbwYB7b/Yk/hPrxmgW705q0oZHULK47S003/pCk8dgoQUWEzfnQMEAyi0uGrYyQc
OygTKCLEeut0s15p7bq3s2PXQSuxvW/0/RM2vbsiIZy2FNjh2r5DCA==
//pragma protect end_key_block
//pragma protect digest_block
wWLu48WzKzCZ16e0w7tnNjJn4Vo=
//pragma protect end_digest_block
//pragma protect data_block
Q7KKa2gEcHPCVq/ajxUegJmOniuCq13noE/mj/qyS9Hu3JaXC19GUMCJbCf5y9It
y8IdaAUhbVQ9r7XesArTfEYdO+a4tOjXi+d6ot/t8CsGqbDZzkgQ1sund19QuE2b
kRr2jUZZPG/VDhACPRJYmzBxp8GT5RYdn+BJKpST8V3A5xHKazz94HdUXvf9mERU
4ORcrJzukUK5S4G79b50sfjcJgOItSlbpmIE/DXw4EODUQllpLL2/2lqp1KfCpI2
2Y6xhKXYjESGwtMDq1K36wREMZYIbmbCbZsA4jfiEkSa5bhU2baMs44PENV/IF/Z
EjfbOXDkzfJttXrwqjqAHHxKEizP7HsD7WrwcnfbaPxRPOUBLhFgaeiId+6mAYBf
KIlmlTU6XuOe93D0Ok96xhEYwuGkAzBolMME+0/NNh5EiLpSs1ZTfbzMo82IMhba
C4QfWnRKrPNxHmNQohQ98XJzsWlIOGTjRPVvb/QxGloq2S3KOUeU5NVDweUVxjzb
v1KRwz662Pic2QipGNnnt4x6FlMsoh5w44bEKaV2iuub8caiPrA6NlAgOutR2VKe
jY4Wwj2cm5oo1rors5CgB/NaPTARvBnSIfK2gAtm3yY9MlU2ZKYPkDvDaVS/tFXI
HEmXQtdjIds8fD/piQ/ytDQkMYiFJCrXyLEX6wGq5Z/4hwgqgBfzsnqpSE6i5jUz
J5A1/dEbcg8XDcKkfHYVCLTG1lWFvg1BHufaz1Od+oS48LfYAvqUfIw0T/+xHB1n
HlEvAXDiPE8JX9bD5Hd3bVQIVS3+iLjuYX8f67xkqV0djEXAa7tMg5oyW0HFdWFn
Xc968H10Dt77mxG8pxqVtRy7m8ieB8BVtxMOiXUQUebO/ezJr7DQ0J54M9KbujWa
OurkoJYorVZfjf4SDyMMNBYZDgEMGe2z0I9yk86hpPuK1iZiwLVXu5Hgd12RI8tm
5mcvKF67VAwH3bJNurRKyfaSxhV65f8TcyPvDMVEFgiT5SZh4I+oFH3IOSyFfq+N
+UwNSGHxVMPZXEf3Yi+64BWfNZcQtjmrCyxHEkSnn2sdi6yipwzNs3Jks4wxoDhR
k4ts78hThKQZxI5/9VBabwvwDDBDA6D2GV6rxwlBwPpCvcVfHGzltnp1FjwycoY7
Zl28lfm4F7v4d6s/bCk2065DDKLu76i6rmKKNAFZyUK3n5bKbJ8DE3l9+9XopmEY
iNT2SCQ65TD563muWvWwyg7fVZq4wZVrRL7LFHWoU9pytjnW2edF6SCGYZE1mPBQ
tszeR5prpPNTz0S8ZTl4iA0FLNKVq3CXpGK8qaZkzngKtDTfMtvqpv7oFk+7467O
zhw35ykqzZVyfaGNHrF/XzfSbVBUBEv2ieoVlJ4zkXs8aT5e5DXkz6WzzRWywNAG
7hwuk6451ERtZPXRf9YfIrfHfNz6DIRNZBxbJbq+7DiUYZRouhrO1lsqcMQWHDRH
MW1XLzIk5Rhx4dhCxCQoS9d12M3jAYJmIWw4ZODK7eAEl4ev/TYyji2NXXhI6YhI
mZihtFRMImJDYrHY2GsCGWThqzhnmmERAzwdbeWh4raLgtpOJ/bePSO7ssyumAo6
usX+M3Mph3pR9ZrOvQtxsm5Ig2om7ULF9aL2cqjxtkfjgoneOpiO8Nn96uK8B6Tm
sMEiiOaXTOWyXZ8d8vDHD2xpkT9/5DEDY0Eegl3pL9Mri8Pu0wbRJe+riGLWgZG6
5MIsO/CTwzoA3OtBXRZNrP6wRPDyDYITALyhxpvUTH6KuKEyKJ2FEfLQ9QLPt4pT
IIiGv8wW2DsmNogIIkATMxD8AXpn8IemjbDGAwjGyNe+FEfREOHmRGivbnXH6TCb
9qyIYqVtcApsyO3bShoX+Nw1RkXfTXsBfigfjEw8Ei1QOkFySa7r2WtgWYrleoHc

//pragma protect end_data_block
//pragma protect digest_block
MX46AKKyFm5ndRkg2xF4vYjTXGU=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
DvVpzKdde65BfBB760RArAT3hMGFhZz3QzSnYBRJtUT8IUl94C8CJ8Dh/FyCBC+Y
UaMtGFWk2GG6PZaiDQy74+4Gc1tpz+a3bIohx0G4/Tp55TJ6PCLnqyZheNOMX1QP
YzmZ/LZAEsV7TtuJpSdM6MnhA4amG2tpwfUX/VD/JYmbXmWWa0bIog==
//pragma protect end_key_block
//pragma protect digest_block
YO4zOWcDgs9Pjnl0JcGZU6gyBa8=
//pragma protect end_digest_block
//pragma protect data_block
pv8HFD7y+t09OMK9K8dIF1zXT/lgRnlmkvW0TldbD3IgQuCOiwWxliU1L0BE2RVY
j7cq+pXheLI+RDnMGKXZUU1BV3Xz9EvqD6WSwdewO7AG9qKCWxcvqOYPAFjIjWhm
BvTZEdzYCK4xYe3ZrUTsNWZiyL6L7hCIeyLfWBGCXLNDjE/t5beGGt9buAQ97HMY
TQT0Sl/vdrJVHNLHdhoJMW78M9V8y3xqO2doPm95+e8R76l15UTGVkG978pbQ3EU
Znp5uGYZeE2+HPnfsAwhJrV48o2E8+pxF/CGxklxbVlJJL90XvkCP1aFVBQ4bI/9
Fb49QVzyd5HsQRCcs8NqqRPp3kwzOuMAvG++H72l6CwcYUjllBgm0ipGkp5NKpYP
S9FvMIAGsx5g8O+pjHYUnCEs51c9PcqGWT99vGtgYrOnvhUmbz15R/j4rUzkGAAF
/GX0XnHo7B4cnxAaWlTFaCjl/ILjG3rVosIaRO+4TjS2GVMeZrqR7lfY25sfQmV3
Xi8lEXkpHN34vE2OWnjujb5EqkcDqeiFoTlfhCb30zhlg+tvAXwfhOs67bsGz9EP
J1jlH5bi29sDociSvthuhiPy7Nu46QQ1o+aW7bE335T5jAVnNdmKQsu+7NdGSNMn
GVQ6Slo/wUvHVyYaDsyWlqyuYPxVPKdS/ObOhCt3bvpqCbYBxaPSapkZbZ0G7Bl8
KC1uLf2GYdQyVymX6nNzSTPN2AsqKQJXu77tQKMq0PNuDyZp+O2JZlizSm3TU4Ed
ubV22Ltigd3U9G+Psv4x6cMyFuqIBPyVc6cBkt5ezLPODuEA9qEkrut6MZyLN0am
A53t/hS2Aw7gjVtyXPkQXcRjyRL3KrTNHIn3wD2hopz2BNs4RWmy/zJ7kr8TC1lX
Z/A3MtC5BF8yuEd2m9PsD5Zxnzx/BYGFalPivcoFooFHN0Bg/t/s3K+AMOPT4RaZ
WNc6YTLBAaDuZpGLZaaCPFVKo7dpquOCulShOmC1cTbdlpSp3A/EIelb7gW21tpb
OnoFwkdUy5liye6EK7dmf5x/R/ZAdjCWT9G5IMn4epyUr47FTZ0gYZlkACJt6NqS
Eskazp6RpqgnU/GF3eH81lKs+UDRRGbfGp9tFTfHKur2TmhTqjoWeSrnHHvCDj9b
vguXE4J2hi24GtYdylPJxxeaUffrQ4p7g6xNCVm58Djmes4lB6Uldk7vilNH6MN3
fpfMU8olnIzYYCZ2AS6qmD9lOSF+6FZovfSsGOYrg/+Lde9FEYTtYU3g6dYEIG+N
DmKb/BBZ/L2zBDeTLGQPRbz85jB4mX0kkph1Qmbh0NSL0dnsJzVhKvuWXf7sZ4gm
AaZi9d28QYNm+XNluZkN9WxlhwkPCvQIrpqGvo+TPlpdw486twOip6ySPxz6+K0Z
EiQgjoK9L6aWRJlksUxahprzmtZgqw7kZ4pmm5abhDQy2AjXdqDw4H2b0jrdcVCF
3jrYl4PsM5wGwoThAjz0l6nO1q6mQHqK+uB+mFWORLEPav42GqNtRMkqChYPuVC2
2afgdGQR43GF5CXrALn5jHlFpSvMcOYzz0ODJl1rFrUmTag4cACfPPXjSMh/xc/E
74pn0BFoj1sMIDdtlbdbNAWsvHG5DW4xDvXAoLx3KtiBeALu1/p6sN8sneP9WUM4
rk028ur837iqCjv8m+guyAAvYQxPaq+WGfA4TclNkT2xN5Wfwfvi4rnezzFzKCOV
twLR1ElO9f9aEuO6zCWjr+t8ESnSeKtQOMM2YoC87ubo0VojqHqM/GGx575V2GCu
w2MHtX75wcCGeFmepI5Ac/D9QZl+20w6jUNe02JwFMRsILjmEj3PG3fRElIyy6Qv
5T4C4pREWojq3KluNSrJA/zGDlIrCT13bsOKUaBo7nFx645DGQkBOIti91zj6dW6
J2C22Tt1sccCHEC/ESrmxpORYdtrfRMuvKluKI/HCSWTQ7WDQfaWTxRtRhh8y7RO
EEgCDqrPxVHJYJs2tQkRyV90QOpTyQej1PHZ95HYaPp5B4FiAT0WJeikGEsX2vEd
79yWLKBpTXLUEKHQBomf8PknOUdhsYw8Rn6GNmaVzKXa532VMf8qCrboH+Cab+js
TD6pbeK6DFbkaNMDV6alCaMUFq/LOF0WUxTAnAaGHwl2VHTQkgHWf6naLar4JgSi
swauuFWROnCeGLR8GA7fEsjp5V9l+rqJrdBFxZnVBhzZArzSBzahFzVStATm10ye
Qiq/WwSk5hL9H8AFlmS7Foru+D+97a73M7mmw2sH3r05rfHQticux71r08zDjdkE
lbg7WlEu5fLAiQjbu6qvhd37o1gavyOmNGwmLBPvD6YLtp9zZt8Dt5aiaxCj91qn
X5m5WnSbG21GXHA59H/Qj5Vu/OGloXGgmAVn3hXKF3PU9AF0h20OUwu1MnQVwaXI
rQV9TPTEWFcisSHCQUbVTe+TFrqzUKnlsHvd7oXtNx7eZJHE8mxr2w37/4/AaRd+
uUqcnZ226iIJDcTT9U2EFGtLF5uEdjs43IxH5yA0b+vFjtKo04GVwCTX5tq2qRHG
1jN7aa+32f9Sbhnhg39GjLw2tdwpipPw7y5Wwzq/e4NQoTt5tkqQV1KCPMU2QIdM
K9Uh6Hn3LEoL7w9otB5WvTHrIrKTUR4bUOdlHwwMihJj4K3UZbY5OtlMCp9qgocY
EM9gQ/2ysDvTTlgqEUTbgEAN6kpjv9xlcZRPH9sG2jDIK4a7Ityf+lcfQGONN5kz
fPbVDOabpJoDwNb043GYVykRrRotwca0zRl7uhDpMKBapqFoV2+FAOd0NKc5xsQw
1621IlN7aXW+NMxgkQxjFwaL4qLv6Ob9Ovp72hQZsMNiFi8hM4gjSu7U5AA2wHNe
FwYiaHoG4JMyz6EJbwqdcEYoeRsZfleOvWFV9UiW0QRptHWimsjun5TwAOpvOiyZ
bJFlj7gN/8eGPVF/hpZO0P8Obj3e/rjS7DDsViiK5ASuGAI7NrNensg+UNJWxW5z
pYdOcJXuYWR9cqOe1cmCtkgIBFfBXz9GTkJUg11m+jus4vU0aHY7DsqtAvSTzdqn
seDVqeZk0OdQfwahDa2E8WIVZRK4O6trFuZRht7LQXVyYjUbsxkuErdkH4p+wkCL
0tsRH9/eay+1pD0MvlPh2Svgtp0NdXcCCdhEjkbUGGNdEQtosxpmYeoIYvoK9NfQ
+EWbQUEDSkowhhXQm/jfOqVraMGfZqjpgIkoTgpQg44kHhU3VKmiNmTZFYmmI/pY
UA0bZygUtXZCyuSRN+qFdkMHnjZom+C+iy1+HWNUh4WcMnhLHeDI9p8gXqx/72pI
eCtFJUKoWYc0n7dxnn5r562E4Xn5W3VEGWSLWLqfvArKuA2kBexa4h1qq3DimwYf
uUdwz6390acBnftCunjKAc7t3dv4w8C7r/hZAhbqhrRBrf+Ldl/riKJktVkutPxN
ykuIUEcUasaboSZZIWmFnFHHb0NqezcQ1ZsfnkBirOpDHWwOwAWbafxZQrsr7tx1
OL8oFIzL15JCgdCAEDR+6dqL4kRkrSukzwf+iUnsn46STJK0oniIIiQtk0E3uNJu
xqJ+0a268p/sjUhoJJ1ma/rTJCIJb97S6tYhS/o8HwXx8fkGHkPXsh+IPP8pgVPR
B8slH+yqeGRzzcXdke3BCP6na2NJl1hLSlCOBA5rhn/EBOeLaVFSEStrAuazQCNw
UwrE9audLSifShAogs4Gm9WpHVA1I4uO4RqMrljLwVj+WkSDFn3LqTmAy/FKnT94
hNIj+t8Rz8CTACpMqefOXF7SD9g5tE5g2yxI4Dofd2EBaZydj+xpTakNpjYX5COE
Gmth9sb1PuYQaasdP1rFE5/kQugBvlTsfj930z8TLAkLnWLsY/0kydQwyVZfov+i
t1AzBv3VZW93NZ6zZU9RqOUAZYcM2KGoGSJcT0GAqnPBG02JZz8WgtYSzRUHVQjn
XTdFeukj5JzJ7zcWJIdfWQPpIOLJyNP/qyrYSIAzKJVUXFZHaGhPWQR/83Pm9Bvu
8aSeU0qHCxKBTI/lTaDcSHBWj3GKo8Zi1cScBdvSTKrVvjacZGAqGU9AqUzRIaKg
va76wpWYZgn8ug8dPY7wFdbnSo5NYbPbvItVSLZXMCIBmp8ZcTDcAfTQdjiFV2yz
WUEMsCo453BmIu+iF2miwavfWQ1A0oERzZ6AM7YTcFX0uTeWCRNeymogswaSo5AD
i3EAJ8c3D4Md3kSVTT4a++pEr7L4CHonNHui4v+pTpUhknM40TxvoWTIc79gGa0i
PVAmvojtGnyGzH58Fx12ab468m+L1bjKwgR5M1U7NCqgOVlSYyIsLDOAjjnYCIjq
L81DXt7U1Z6luGAYXrle6gBEtaqm+NYuuKS2ceUfpaLKEs34eQIQrn7LP6Ey6H0s
VZdYJFafSNAEl4pzuXALRLuzKYABBIG0J0flUZrxSyBxkWLeOykDiv75W8qdF1Fi
RuXT6uknEYlfuACeYjn/B4rEIrNIk/zv0wMoMcG02WtHQnfeHcHjyqJQD9xhjunw
1y75BtnDahjD3PiLYFlxcmGL7Lj6zcpVr5x82C1SKC7RI31ds4xOzYKRav0ml/bO
26a6Y4hGNE0rLpk6rGlTykXA61GHAJX90/ilxlBLrmeJVM1LgLe+FE2tfX16kX2v
BoR6L1IbQ6KBhoxq7ALoBLMiRbEgNXVRaUJKxvSHO0/t98vB2y2zDFhyV9fgPnMA
z9+Ro89PJ27w7rs4YObsZrioFBYhUpvU1v2rz8sKX67EH1J4bSXZ9TIPwTsh5dcf
D+YKrL9J9YTkw+tMkbUy+gBXxK3bm1WYpP2lqFotrClERGvpcTjt/leo3sxIU7Kt
rTn2TRDDB07JFshBPdrIKNlgb8jzWpwQJmG8GW9DFbwN93oM1LzahGeMddD4vfKO
g6wHiyknDAHs0zui5fLkEEH461dV3T0qeyrBoOd6tKhoj0aCaDHGKK7v/XsLIUmO
YjSdOTcSiiTiOVU+q+sh68LQuW555BDCmWsEi7hv4+s+gDOczb0RPfDruRU59W2T
BIN57+RjZ63Qzxn0I7Nr/TcsiOyaqP7T0LO74iFCqn/GpDnSLzs2y8KceUSDjxhA
a4nct44YskcO0VhKa5gy/hyf8UsnWDprDxfrzjcmMyJCgHQrZFVShUbwOMqfp5Zh
7ufxjJFE6bn+P9eZv2XNHu/KHYj4NbAUNlKcmCs4V9XI66DC79iesuBf5JrebdX0
Hb/w8dLQN0mT6OeBM0aNMeLfNgZYM4Mk4O8/Cily0B63ZE+JYYiw06LnjitD6Chp
XG2YlPwaCmsEWaw/nSFf3Wqly4QfCg9bHuB6gwXFtK2rtVDpE5we3HyX1Uvbkt51
aGNn3NqY53LNXBV/+FKRuJvjdUQS8xvigNu6QKgtCXqHh7KP8LLCSzcKXpYLVkNd
zHU/3mbQzX94dOe6CxHqeOR1CEPhGiXE3rXZ7i/fSzVjWIxA76vxDxOLnojfh69w
AeJJnjueTNyIYKhljNEiIU6TRoiBK0wFlAmjQ//xQmfCtaA5ae/dsVO/CGWPyL+M
X1QarZExMqiNtUH22VW+SNfW4UjyCkc9mNOgAoTJ2nG1613PDaNH5TY/HhovN/D1
LqZI5pvSXmuIsb94qDWFAdOAHuUiG9bVrzE4oLavhp8YdcAn6xDGX96IEYycSJ54
GDet8Yrurs54Oen19Zne7BSpgccH4kCcxAToFD6x6CsttP5G5gqvZbiUpNEXZ7r4
tCBbWxfKQS8Jtb/gEu0siO25eZZDKoMuBzSmmuA5DZhlaIR4GifD4wfUG/NC9msZ
nOm19kC/pOD/e2KnMk52HTs8f+Hranl6QXuMgnkXjQD4hBsiLVNlfQeVV4CmWFpS
v/rdIx7HrqskRlPOW3Debzjusy7OKr1sXTMo9SWpHR5ycAD8Rn0uSVWf9VHF0x7n
wsbvQD81C3Uisw/n8Jx++SAxMHV2PYUUu+GgqDQjbZ8cYOeyMYUpCLOl6fBDkJJc
tvvCqYbFjFIJjK5P6Nv9SqBYnJ29fjDiF8je62ipAZ+vtWcYvXRMhQQSa/79RlgQ
wPmnB1CoTYaJWPNt4DbiCrpUAluYMehL6/KL/mv+Gv1hTbSo+qbOtLlVxfab6uZg
hQZ2b34Bs6X6fCL9hz77q+2sVR22jVq39H+ChK/rS85kcLOFFLMLtjXCbzPyWRqK
mnYX+mjBd5sncEW63dSjJksjG5HHvyIdAkug60O0PWchoI5zEhQ1hsabf4WkZJtH
RVC/CE5CGHq3uokncz0NcaAooozaB14d9+VvIXqWd9LjGblmcXcWEg5crq1pY9MJ
HcSa7CXxWGWfFu3IbanZp+nXhwA+UY7Sx6neh6PDH55LnntlzPmV7aOML3m6y7xX
eq+AUQt+yEDZTCgFjAAk23EB/5+2bVATjxIZAoV9LQ6yVk8b1KgwUDvi9meyFBXf
uIK2cCy6Aq8jw6xQgkUPMBMhaEPmF11TSKNfQuEcjsCBz/FtyhG8IprMO/Q3km+N
T4U0BWP8pMW7fdGwgl62X/25M7Hw2tlSRiPcfBNyV0ALkvzH+L0gbTgDd2PaatyU
8GP0yzjklnJXgax1XgvH86NtgXvSsCahYo4+Eind2GuPbf9/necjyTS6M+7JGH2v
ZG+1t61F4xzu04B9Laz/Y/vI/FehT+qc794kZbrlVG2zOG6OcnCNa2L8HkJ7M8Vj
oT33cdQuP62gzsv0zaDc4F+DrdiNvztSIAGb2fCiy6XJFdm4dX44is746+bn57WQ
uw2LRyyxrlm3S7O/VruRYISkG9t60BwvXnI4cVvk22eCNW8YQS4BlrQ85Ku09DdN
0zGrq2iAZuZf6IA7WwHpbAzhGralVdTCFtMGr6msV73oFDizLrC5Rk4UydCoasv8
uYU8JLZ+bCSfDCFR+HpL5TlWVXIH73JqdQ5MhU41Yik/9jvosN/t9wu8tcUTG+GK
8EZuBceoJQhOLpRAdKvHRqqM+9dn7IBixQ0xjCxcdxxuK4/UR+25caBfl1+6pSGq
iW3yC8/MlHzKa+AMbHKB+FZZzB2sGgeOLdue+1fbEj3xx2wy4V36dawarGtpxJ+N
hRzqdmblIHVvGzN40iPyXcqQvRoqLz+D93BFNqHpAB4IrjofoeNHyVO7eJ7frXgR
ylM84NTqhbkdoRylQCvBZ1Go0dAJadjI0GpySQyLG2EHtdnh+rMOhgYLNQ14oIC0
yloYsZllplhqHnkLB0al8KxD81KUZCRfgLKZ3YqRcc1bq2qJlPRJO1U1ZwLQR6BO
f+tbIWd1KtER5FucdbLZKeW+osoTL+trkFbkDiYx5iTdtCB98+vdZZvx9rh95vb5
g9kcuO2ahdOJOozVmKut9wj3fAxH0i84qUn3uyEIPNrV2GE3jog3YJ39bZqUuY4p
USYRV6P6MT8nYtLnqUwvLFVdIuGp5tE/g/0PpRQEhQBlQbpb4RULta+TJsctpHtS
+Wwb+g7cNftq+bMiLdFAtwPBZCNF8Ed1qsXJySG8vYAN/P+2r97CW3EPSsZGrKxC
Q20u7IANnyBSoCrrYlTbQEoTArwEn13xuXXtNM30vrsVfed5LLDTnDGS+1E8yqIC
i7+/LzxVMgJjcDKwH49iRXUAUOX5y4yKV23Z+u2EGVhziReD1YSoaznNeZ4RgYcY
Fd9esrDcNvmghzukgSHAC6AmE/OBYC3YtaDvRPqfijiGN0ac5a3BguWlu6BVkDuI
xsNxcsrQZPrsZBqZmp/8eATmaTIkCbCRdX2T7i5EFJCRAQcHEmdP4Zzx1sGG7BZU
eCXwr+8pdadIWzTdAOpEt5D5qxLF1IITjTzfK3mJArnZkA2MG063Lnecr8Z9yMvy
7Od8o+YuJOmK1nIP9ev89g2vAdoXMkfugxYoSfAjFh2IMvEouvaP28h7b5rQQUuB
kx2lio4+EdBSy2zWybmqow7hVKRtGSuLWVWr66NOX+bwYClCBt1Xw2rNTHqG7+Sh
Xr3Wx5Rue4oHesppVgHvxCI98+1PDLZlfOCYKC09366vUm6FcLOp4+VHdKqIJzUS
IXlJ5FqPDmu9YM2fXmkAOUkmbnG/zwBJ+JMm06sIOeIRrtePcg3y/+dRxBmtGENr
JwriFfEmWG4pipG51ydRpIPe9600D+I0b9eFhVKQqErUlJZKgV6VeGo5pTGtOn1F
X7cVOnYUgNdVD7/qp6WwJOdVwwEAqVQbQzdaFq7ztEL+4ZFhLy22oJ7FmhqIpxes
U///gEcuHlP2SWvMLwachr0uzlB2+/ciq2slY3lET7BJwsf8UNL+OyViqNXyt0rr
AyCjcoXJKu9CsWrjpCOqqfYLvj3D9+hPjbnJick+I+0X/7i16QrIjTNhiuAS85cv
MnfDBu9UxZ0nEMZicunEUrzak1EmQsyAENLcU6YrpvicNK4izrzrZ+iAv2OaKjqP
pHogz9l2KGrkM+O4zQQk46KaXXBsm5EYw7wlf+dd4A78UJsAVUHLs1FCBS4F6IyF
9o8wcQSsU8R1PYpN/fbr/7nuntVgUv6mUMY/x8jrL5qIPWIKJrB/bMufnQSJ411A
7sDGyGt6MQ7h9ZXGFA0yAZXJdYcFaQx3UWkqqfvBjtPt+19oRw3Ulvyv70777TpN
+b9DZpEr0hxlb62IAKXxn9Bb8wfoCSO538LlUwiEE3a6DE0xyrtWfulUMkdLqOfp
iBOlGhyvKn+z4WnkDhX2lG7RV7OyEF6HnMUBiuO0cLBEwohdg/st0wyosD2P0jHV
ayi3MdCpPEgC+FPxAOUWY3Oi5U59mZUuv2IR80LxNedhgVIwO5WIUQ+TG5NIs+7Z
QVXvll0qyflZfjRfeNrXcOgq1ZXxGbsbth0fHN9+IefbKqhZiGya/tL43zqhDww8
EmL+HE84O8lqyKqHaU7dTASFM9/Np2sCMeSVEZLbYj3Hh9tqPHTKidYP3YoPjpzU
zAnzUhjt1d6Pj2t3r8g7ykSbA4+uL9dxc0dl46QyyL/dM/+5qrRxK0VY1oe6+a8r
U652thCW5H0toOf3aCEMzN2FT6rQ6LF25ken4PGQZm882tFC2KqZPNBTetO6gt1H
OQ0k3XmhvICIaMtaUqt4uAcQL1QD9nki1KbV+XvAmxyJZ7HQdyAH2VD2vSyE/b3O
G40Uh8ujm8ZeXQocFHFhSNOYuGLC1P2VSSw5wtV4FTTR7GilgGidFKs/JQnadp28
Z4i6vVYgmEp5GfSsAqtGnt8POz+rEmgMt9/J1waNcvwEOoRwG75JeQacIscQadZr
htCsw4nkGigfk0xQKOw6EmronwQbu4iQ17b8hqwLeWbzabNhDNvc4I5VirQD5onm
VwByS3oqxPEH+ktbMcMf/wegHZs9kzOH1OYnW9WYI3bNLNgXhf9W35PMBFSwWKcF
htD3yO5uiw7tzWZL5c14s9lO8L+jVIQw16536E62R5v3T78ksiDjR+E18sUcmZ4t
n7EZJz5rIoC4JF/L5rDGGoOVkp4CNoEftbp1FwbR/KWI2sqM+P2LCeEBfrUVh76f
eyj6gOZR5Cq7TF1pxabHpDH59Bh4lWtSUaaSTXE9WqgkFN6f5lOzzsGxAb45d7ic
5W6MWRZj8swExp89qSv03zdnd/ikRAGuWvz7OeABIoNJeAQ12z4HVB5/5rmlfoXz
EteFRc9JylYHEE+9QWuPvnrG1cZO7rHUCCXE/Gxpxd8jJXGS42h7rZ789Lv9oSQA
9J7qcKyMKkIwa0ERPRmOcHZAKEelQZCOsmzAbd7VIiLkC8mhB4e/Iq1qk41rikOV
tLStS9lBdGwBxBFmZR860hQOfSCHQrynisVyDMmpuLk=
//pragma protect end_data_block
//pragma protect digest_block
wz0mYY8keo0FzVOS4FwZ3NMEr7k=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GiaZ0z6M+zDvgCZCWjv7YIKbEbjZwdsvtC2jTxkvDIwG9uwEghehjUpAqsfeLPaD
Q6S/9P/Oiz8X4JvO27UFCr7pwu0VLn1HBdv/iYgB7xUuT2hj0qtobF0rL614lHFP
ULlq8kZlHoBbXEyKpUzq4K6eFgnAH7EOmKb0lV8Rouw+dxd+r1aXpw==
//pragma protect end_key_block
//pragma protect digest_block
Dbui1ASk2mqUsQei3dFa+gBrwe0=
//pragma protect end_digest_block
//pragma protect data_block
W6rneWfAm20k/VmPv4faYcLVF3ahV11C/F96+eCgu7C0dnrq78Ojtr/yn8t28TWN
Zj5assO+b/u2iGo7DaRpA8sU32OnZWKexCqXDikl5jAU4Z9d83IicYiJJu/eJI6H
efA6zjYcKkjo4ECan5VVn7NsB5h5l+hr6jCjFv1X2P4dGgvQ4rUX3Ec4xpaptKby
Ktx1JmtphpMh0dZFuBzg16mfNwtKiwxpr0/ageHt5hmLNMTmEQOIX6G90luPT5/Q
uK4iZG5sATyVO1zIGmVMysBARSNsZV+4hJ5kXvTQLJfXfoarD/FN5bTHQCBj0CG8
ZBTv5C1jfUOyfc/d6drhN3o1G9AMQrHbnFxgDH9JjCuZEDIm9P3G48kjS3HwuqPK
3oI18Hzd1BKytOK5KLqR2MFwYziZyf2IzIMOu4a2BjDpJdIkbvxPNhM4CXFwUz2C
nPY1+lf+CkNj2W2v2fJF4txju7W8+a5YBMfthLk1Jz0=
//pragma protect end_data_block
//pragma protect digest_block
IPLJ937FIsLg/J25AgBPk0wQOLQ=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tJs+4KFJkEAyW2tc1cRrCT6nH9gYpr7hIRN/kVj+fHwILvUW/mxw6nQO4aR9aKov
GrS7yt2Cj1Js0l6SYfziA6Z9dYkF3elVcUx6p8CURLdO+wvLghFwe01FV5b+35Pf
tKVTLPtuuSoQLaEWmZw5Ap5IaFCmlXHvj2OgMdh3/mxyi1fV064bAg==
//pragma protect end_key_block
//pragma protect digest_block
ZdwATxFZH/0jlUh0XagE7zyZcBg=
//pragma protect end_digest_block
//pragma protect data_block
4OqQDvmPhNEJL4mNccrxAbbI4K7QH/aQpoHEXzUXdjUR7vmcJMaXN+qXVbC05kPf
UlCgWRXI4IXUheW3fVv1XSjVgOHEAkKUPyJtQXDmz1qChEvtMIzQDuSqxORbJbry
X7PZglbvnVQtvh/vvUSzkVNCcCGf0Szn95mR4ceceiv4SbvrVGGZvo5bir2tQtDJ
e15dMkSzb1QvUONJ06/68hgrOw6pyYIqZ3SEX39i4D95yMD3mE5fbd6sbo4zlyp7
wrSdIDbNc5jFlj2jDGZw821dZHeI1THHG0UU80ySj9WjanQQotLmAASJOFiZz2le
+b41SzM4hsrYqc25iOlvkIiMfXFpY088v7e+1mdpB1tdr6/h+QNKZhUxJBRD4Ltj
WS+kRHjiIR3n+1GgRpoWlvUnnxWV2tKVseHiLvnOVHtQoBd4kZTcunMFKHpzXdrp
sRwytOSnQ1AZ2yBhbocm8Uzj4Y0lnKJYu3dn2GZrk/3i2Js7iGHEwT4O3a0Bznr8
bg6H3pCZK/kyaRbud9nrkE2gfBiqGW3rAOFlsfwxgQ0HWt99AtdLMq6O3qhbt59Q
Q3jEiYgBEE4KNMclhWeViedjjLW6ZNM5350DDEMMOCF5QUeA+ev6UBOEe3MlPnRv
qZFXvxpK847Br9oD4Q4wRamRRtDAgZHfzHO7VSPpjDgR1S1oaujL91/dvaC2HDeu
yNu+tex0u0nG/CJ/wHWDsSoBHtHuTPrXVz7SK1jTJyCXq6Os5acVQtwo2rSuuJzA
/p+2vSiXF1rQWiM8rcwZyVjljBLBD61zq0OCnDVB/nCx8lBTUXt0Wk9kPxH0uf/5
xmLO1lk/EXsrC0xBuWOF0YGvYM8MxmVVoj/4dtJjQSqejSLKIFTt9ovPywcfOIq9
zbwOWMPQbk6m+q5hAklgjjjsc5tD3r/JC8ZFsmVw3IyswAV8adkHK/b7dhCIAVZN
WgLuBN52dvqYkROrDS0GRFw/Kt6ms5RBrfoENv3CIQtpH8+GaVeVAD5LFJ0y6EJY
m7JNQEKFafv8fQOQIoFTzwiFex9+m64dzBaMFLKT96cU+6XoQdmc7WI3fX9sWm5A
tTnKxosHeWz7Aat+7sWJDhjZwtM8kXF7wzOYIY8/qLLmDFVd9QwSkwX+xrvAtkJl
k7q12cV5m530D2LllqBnLrdkFp5YwfMx+sBrLNv/BKCDul0wmSL9rMGL1WJ5yQT5
5vrwPn9XrXagJe3wdO4vBxatenynk+OlNLFC6Xvy6znowhyLTPb2M5Z9eSttYljt
lVgApfYa/wU2c291iuVySqi6YGWndEUCdloZc2kvFPhCBKgMJY+aqZ1zHEpT9r4J
HTl7y/BoFrYCJGSmalfP8C7a/bMBU50dE6AFTeJr4PU+7pcwy2Mm3DIYN/vqYcFF
flfW+Wc0GMY9CvrW7cg19nu4GN9AnkE/gFdtw/y+gXUZ9BPknYkryfbQEj/wDXwe
f1lpnVL2ZCKExD9PoCL7QOPrL2zIJp84ILjWMylPbZqM1gtEjRNGlsK4FtMOjiz1
1aAbigx2I55NXowKL/vs3aZnUTJHQBdKS2JBrDzBav0CMv1cOe6lsUG+IL4iS5s0
PToBM8Y97BBojZM0JQnRXB+iEnpt2+NIcyNJ4CvR2uC52lpB7f5k0NFzzB9loGTb
xRmbNgr979YV8vnYG6Ikww5lWf8Hxk4nubZOlAiWeD0sc59iF8f+sxlyGLgDy7x3
Gv1a9r2AO+1xR1NTl18fwFd4A31DLQlTR52T2HgkM4EEc8UUgJrb/kOgXB3ek+3b
jzEWfNakAXij9HpOZ2OSLEf+ZiYxWO5xgM2ZNLD1oBZk4ehsHNJNp8SWOBi/gzom
PVAZ4xT58f7LOjLNTVhWdwFKO9u61kyap3qIZqkPZ7nVit/MIb5IlUhu9BhZEbz0
anZTKHueSYieYF2vZJggxhMo+3d0LvlH7Vv3VqKESClHE6BozNoS8y/92sfN3NwD
0+24CCwg2GDthkqCfjxOyMwxVGfZ1VPLwmtvq4fvMLJwZoHmcjjXve966JKUV3Jv
f2FEZ67rpRSyau3kVV7mJCRgAYSu4LLJxBVuB2tdzGrVMVPCHJ7mSdSQLQWzhOEv
Kb0g7DLaG9/nA3gSu6/4TP1K3gQPaSdRtALhx/b1/BQqHa7wAke4xpGiet+MF3Yk
ae05jFryhX244YvKn3n6sWgJI1fX5bQd6SVeiBXcM8z5S9nO2Pw6Bcc/P1/5l7WV
0yVUVTThK32/rsmdVIptT0dpYFZCc2VqzZduuPErAsKcsNmF/bcfes3RJb55Dvdr
vTh2U9qssMMDrqq7Ylag617zhw4UFeqqKgkCf18LiEErSGfpCsAC5tjOHOPGSKWm
QgdSMrqZkVak3B46Q8jYmJ80VeaSCrrP21pVSBLppmAwCI7tqhlUlzyEzpUa81VB
g826+zWVY0AszI0VE9HlQGbuDGiSMVigWEmVxE/oTYhNfKIA2BN7wgrIMo0Dx6E3
2qMj10cUmrD1G37Ppf13olZpDDLGpQzX2+iu9JVCECJafc5D3ISr+jIy3xpwqsvp
ftSMeFz6YoKrgcsoC07M+lgMP+irL27O6yqx94EzvSEDLB4Aw+asNEYSObIkMyrA
qr8C6c/Axb5OSuH5MXDkZDooDoR/cGUyxtIcU0TC4ys3xEne2rr54CtvQ0R8a3C3
kCJm1NubfH9muVLDoXOmQ/FXLn1kEteYZFS8cZ/+9UjE9wDyvKQZLDpBatAp4sD8
Wqx/oAZEASSSq5xDSUeJkaDWHWHi1sfP9ZCLRwzQahIcLg/Oy0Yi00Ia+IYGJuMw
KiMhjabHitobuagrlVhDORNdgOQx5kB/YugvoZo8MQMLAwC3V3RtPFmTneLDzySD
4v8wDrNboRx9sUWNdGdFu6dwYiq8cm7n5e3okh99jHMunmvLoSbD1tbku4FRjYV2
rDkuHyFmSR9nbMzH9PGu849Eez6qMxMun03IyMjR05M9P9zGxctRTpRlwHRiLOMy
1KGsHTlrveT3QZKGNEayz++48ZTb59O6p8c/zy4WullursOZooIECZG8wHAsrj43
Vi+lSPvqnrGJQ25ysMUgsrbQXafNhXfrpO2w7DwE33zFBdUylBuyNNwFbAS+6Pdl
TmJxeLm4WPAjbIrtCqs/fubOG7biBVo9XXuJ9lP1SeDbMXRPxftzsvxsxJ0hUuil
LN0gK723VeDv7nU4XD4dIAQEaCncAVt1uFQsSWCtgaGNewPKtmG4w0ttsZraafgs
xAoSiAY1o926R4tzktlwVvG41T+wLWIey7znMW2ImOb1OzmQ1EfKrJwLaP4gcnQd
AtXf1nupB2jAHlOVYXTAic0Ad/POJeSiNpPdvSEmKTL6clFIbazjmrd5bOGF2QDW
L6xGbvs+7c46H/BfEBBlcM9N+OqSsF/NGuftMsHv5cjZXlx712v8KvF42N1zJTMk
Uo7OArOHwZXUy95IJBls+38YpEoeORSquEYpMhVouewHQwOBk+m+t0JWfzZytYMQ
fd1AkZa+M/wKR5wDftKORNaJkvCYzBnsnUpm65iMRf8bCoAqTdA8fDfscTdFxTSd
XEBWL3iOwXilapxTlpE+M4ey7zEQMLGsky2uyee/ayLBn5hc/uwO7mMCIn0Ui1b9
xa6oLJMZo64chYpZDg8PYHtKtof/1cTY2Co0GEicSumhbWZeeZXZWVfBDyMi3jBn
muVng1HlE/xqNnhzvYKzSaxjIHA2Q5li8N6PZEHNWh1bTdCOKetejOb8zb0lKSpO
gRIpZGm2RMmcaYyVMOBhKZtSwKy8NyAi6mQjDz9ZcwpYurjZXWizts7J9gIWMfRG
6GzJ/MiocpQULBbjZPyI16VsAM6HKAchJbqLACFt5CZmIw7w2CcQFnR6Y2jadX1Y
jW6lC12v2bTtAwIbFQaCXscQulbW4z5iMN/q8cuTc9GoYS426z9/euuT4CYiAlFw
EOm9kbESX8xs2v3Vr0P439fl20dNTXigJv6CcmtdSCw5ZyAV4J7MtJmF/vwHHb5p
YxIRUaztBEKCAHj7WciBWsS6Zn+1AsRglnUUhvuFwUbiU12RzwGiwiSgVaaAZJrq
ttjjkKqBLZuM4HgTaGy54j4pqK6iQ6h6VR0QP0gH9qaVBqwG6DgY1c+fm9O24159
vpxeIZKGqz/qs5mG3KWhx/APg+xo7iELCFJlEVjRfSKu/b0xCa60r5hDHusf9iux
mIP8F5TvfQATQ9bl4GAvRPFW6ehHj4HgimJF1K9kbL945oIiykFR7okh8IKYgnhQ
K4aY1IADDsmOI1XzYdP7fhXVPbgfG/x25E6lIWUo7/ifsLm1dQSS0igi6AKhrqbv
dryJ1rTohhw1GwCoZAcJHxOi3PcCoj/Z5aQZn0y1GkrUrY6+uATHsycY8Q/EVt+W
B5HAw3gGJHzgmWVWz0fByRwZyMPuIAKgwo3TLcUL6aE0gd+b4VzAEH0aXKbtFV+2
+pcHoXTYOV4OMLadtIo7YsKqVecuQ7JKi5BkNE4j/hHrijHQb4QrBGvtqVPu4I3Q
8f+CMJ93mao3ZbjDarXxaoBdpapXCLd7R8dOtxl/ESHXUs9QbyX6CIjH4qPwSuVW
ApyVljOV3NrEv0Dr56FXCfHGD5ZK36PUM2ACnXXmD5OdSk8YXFN5mqWeoeuQsbj7
u6kKMXz0VYGOuYTqu0HsQpChEQGMkXTrIPS5W9JV1j74UrJUfw0eLbRyXdHLQSMh
ZVlsNtGaHypQ28/LHlzcwhvNX+cKOjR96x/a3yJ9NHjgAupOygPs1cfOdO7/KMmP
5WNyg11DxB9h3k+jlpT0Tnv852DIdVveBsPY7nqwbTBlOzR+wt8dRMbmn5HIlxvU
aUN96DJvKliaHTMhwnCuaPUzKabJ8GNMIDxIdBQ1D1TBbHjGxIW8YNIQAO0OojiI
FmdzfFu3GpbYEq/SkgXeshZERTwlxpemWVHjO8uEYvqTPTS+sM5+Hg6LR8XnkZwy
I2vhagNuBJGpqVVFvnR1VTPdGZpcmJ0+p3+HW5x8nRuE4P4A4fO4UZkQv96roR0b
eYCG1O3uEfsKo3+t6UaR8cjb2iQXben1VAytkcvcAlb/MYjgNx78nHc4PgaTq9sI
n5dDQMGC9U3zo2Dla5+Wd7GpnirfXofbLmNerFDaKGYDJTqASVhbUfbDe06VvEWz
VjgVxykimE0HPY9tXE1N+oinRhJH2Pb+42KBYWOwCq8txNWbGofPTEHtrFA/MutH
A728NwkX+l+PsNvoELrA3xVLBpT4sr4qjIIq65QfLB8Q9DqXJhODT/kmcr7KIqKm
YjA8z/CBzBr9vr+aepHQzMSXP1JjhT7/++9gCPybIX04BCAA6VEfs3E3YwmF2oed
XLl+hsrid9/X1wo/oiSlNnX1wzJ+LrMXHVi3I1wQzVREfXEO8ja/AyJDqbR6GEr3
dcRcya7euqu1AVPYgDbzi7ez3YcoCS3asmDOY0l+tCPH7ow8+ec9d4c3fiWLQCrR
n+t/UZlXZL38tgUzY4d7gRhDj4/Zjp2XIHgNSDAwgTf0gMH4VXu4jRPyUE3rGpmp
TucNBg1MayMnumLLgnsqZIqTw/0VrkFZyK+Ac3PL0geGeVIz1sCD107vIK8NTSD/
ztfKCu8II3ry+lMEdkSSvWN2zPhWxlhd+WckN2WYSW7uSU/xvCuAVLA1ta578WSl
t8jeUDR9Kup5jhCQbKY8oR1phveRWkZe91KZ/28IhDaZTSiQJiaPz/fz4OZN/Eiy
0QxbuZ9/+WlyIg94b0sV3l7D7EUYDapnlxAa9pIRFcRnm8FuhWxgc8m08RBKwe85
EKy7xvy8LbhHGrAhEp1lY/0yrdh20AXbad0zNcDpk/bTchcMEcCxihQydYVWYumd
/s7qtATz3RJX5vQzpDe/IzqSAtyRmkeXX9bkTvSehI65EiwP6AbvSJ8POFLcSv62
b1VdNkmHaJQ1Agl60mZsNH202gVjen7Vp0J2LDTApfP7AifZdTUoo4lNvwBYcBnG
yhBE8yVQlCHrMSb2HJH3G7zRqxhw2FQVHXUf3te8i7YjsWpHR/ZFNUMlFsNpTP4i
T7inWpSA73heSzG1Xijdd/yoTVeY4WaXlwn4AGE/CKr+W3ubmgFQ6LLfirrBpzPM
snM2qPiW9IZQJoDDUE4HAkreOOMmktzbczKYARkP9bnfGp1695pbr1pc2eLCnYGP
ohKFc/bPai61PHrH7KLOnLdCQBB0lp0Sq9T1hwCKXImOtG+XTR3pIp9T2FjV9Iqq
o18vZW2bePz8ZYGwI8hnWREwN7+XnE4KtsbxKU+mj7gtLyhY2BCskF3/2aS2+0mD
B3yvmR6uXwSUyPq5XKAslqTV2QhgIkI2ySChsuse7ABRaGXvPDKqVdhTDwfGGIDJ
ZHoWBg5S3On0wiQHDm9JUbUphBC5z4RoHjO6X8kjqz+o4jv26pX7UMfv9+pLxUG8
io6NfNXh5ai3STE041uAATuXFTM9qVHsXb/KhsRWAL6s9iayt11mPRt/SwM+M1TN
AqnHwRiW7TdKwgpAOTQMeRWi+Qs2HWprzHTWpswjIP+HrRa4DgWRX7dUW1AIX2rW
Sr7rLYGiCr7EC+j89bDQtOaoLS6thfS4kpsuxiuC1g+YzCdHCrdeUXP5crXWCrcq
ayG/Mw47oJhImttiGPZtxnUOM35JPughsDVd4I468NP6TeC09mI0fAz2xSEN/+jk
bLl9txB0IyKlEHTKRjib7t4paX07YL61wzyT7B9KPslWASq/8cb++iOgaGdOYhn4
JNewXuARCkxwObxZHcCQe6316n/Z+tH/uXE6LRzL0xgh4mY+1JkAnjXpaSw/z7YC
NPtjAoc1rCg4Wy3L5H/6v0LaIR9urjhbZkfRRrPiCArbE6nn108EfhjJzHlp0JIE
xhobp08SCngWzUaG/T9QmkzU5f4fTwbZwVB+qledbEdvz8PFUib4EyK0GkrAFY1A
thjsyDe/p7epRPdAH3Lq5b7rYU8y7j2C8LNCoZBH3P/ZD1CvkLV8efDNAPpYDctL
9f302dCUYk0hmC+FunKxCrPQOy8HFJsEEvQgvN4crpAHj+HIqgGZX4BWHMjffJnB
Uo251sLnnzO0RqjC0B7plFjOhhYPl2tfPLoQ3djKl2qr78dz8OAFFByd+NGHydYc
KopLy5VWsmO7LkDjs7cHtHW5mXNm6ZMx/mgew42+kb6hcYR0JdgWsJUgx4XFtKhr
gd27a+X1Sc/2mv5khOi6Dv8g63hNpnwgl/kB/sOT16QvoGb+7O3vIx8iDvQg41++
6JAUdGe7cN11OZn5hqaCwKpnFT3TXIZ8O4Q9PHbDcMDeTQ5vLxnWRkHlHnm4uoyy
INlOXUJEsXKPijtIwNc+HZmWBuDS0sRQcU1qLJEsGkeULe4ienwjol4i5cK9wEMB
0Jut7lB15KbCPyqbApStjswlFfqt8+bF8zY3KWuZtwgDZjI1k5yN+uIxuBLMlAZy
qKQUdATRwrEFyYhnhNWcDqUkcKEEa9XnzlN/0X2bC6L/7pyW5B71bHdiO9VoV/rE
oISWCeskwXcwQWqdBBpm1az0Ncq5ugIP662FKAALQjsoXxCUERM8WQbXxJwPXezn
CIASE910LGHiNxc7z5YWPJfU0ckhJXjNuQ2Q418U6352S/PzLtFcQFEryNMga0Wp
lfWB5I3/kOBSxexYsoZOvDqqnKaLfpfbeBl2Cmf59wdUT2C65nK/XP0CV39l15L5
lyNfU9uES++uo30joJJdOOAFjzneGq1pXTUfQdNGPY7+pqVPLtEo8Eir4EjOkSQR
GabYOyjmFiHr9Ntv2oATu9pUNDHzHmHK3P1bI4yKqp/bKFwjkCrDMTq/gWuIskIC
vk4X2p+DOL+eyTCUdaXOis3tsJTKxqLOUM0YoKDXZ9powDqQUD8056GU+65Pq1R8
EJQhVLx7lqC/Mt63AXJqo/QqadJTSAUjhBiBsvRZ5LZIPpPglC0w3mxgk3e0WF/C
bFi9heLcYmC9bJVDcSC5y4yBDYkTLfepaWxXi8vKXJT6jYoQJRKHfhWRJbyxy/Ip
nLspkH4WYEQcLPKf82TtwwHtN93CV4kk6EUOzOoofHUMIubwaRb3JZ5p+w+NbCVo
tp8B5QhDHDWm4zvfBJ+2KW920SgU01G9yGTnHAgnvmytH5GXWEPphXmIGw+JCaKt
0wD2gN4Z6yefhn76sgPdHZ+8U3N37HtQfj2rQDMW6MjKJqt9Rg6r49TRLXFMCI2c
UcR2om3DltUy0GKDTUUkc69DG56z7c/Uh+3xTM8AtLo7dGOZqLhWF0G63HgBKxoU
ACGUaqvAmH3aaDjzc+VSmOf5foYlbOizNkeUpnIVNFxuMVGSAm2HbiAB7NsLCYyQ
sUI1hJ7pSOgqS40QjfaRU/F18VIH6K5RjGmNUgZVy4jbapNEnGJpI3w4lqVJwiD+
LHwAd3fJQz3l6/C5q3v1sxzQjT0PfdYS05K4vEsdKXS/uKfpHPdDePWz46w22mV6
hUeKuLtIyMcClQ7/ApZfBBUQARpZ+ePs25++8kCy1lTNdxsvp7pgxP3SHLEi3UC4
9MsgeUDoD2GPVe+x2a5Mvj5ZztPQTALKzQV71/juL0m/Cpgf2HtEiyPKg3kjZyx3
8/uGQg+3rlttw8HoQltMHIUuMbLUUSWgUDFLwZhQS1FTkpcrZdcGS6L5TiMuoyML
VajyHrZNigCRt19QwGE099UhQ2L3du9ZluzitzBq6sCe7bC4nJ4Qyf7h3m5UE+Mg
HnbUnFGE991ocqkPmcs+3nCc5pYiwtRNyObcxghL9xoXYeHOMAFnAb6QiS9z9WYO
1OoFSSMzaKQq+mO3zTkgavg6dWRYS7/Dv0QUrniGdF6nOlxsLN8MwVFHWDLx5zmT
iap7+bEYUUNk8qe37tGcrAyULkqBx0zY7JlspZs7+f6WB+gR0pfbp6owj29czqiO
NpCGXHfr7zEiyZFT7j52QCDfTjU8NhPDKrxHXbGEbOYf47W6au0qFg/S3b9377Nv
HpHaCNf5HE2AkMrkBHxNxXJAZoVbv2CYorDdsnfu38tniOvSi4RH8rZVNv5znOTd
S/Mfi32pTx+E2liZvwq3dsmt3X8K0rY/I6r2t7MLiwcvlgsW5/kEAn8fNDjlpXKB
x+vO+3aB07/GWozuEaGD9WAYg7GuMXWZTmcbdFKplcRi631TtgWI7sG9rAuv9JZD
n/ghUYGG5Lgig2HLhxCbLaCpwoH4ktg0i5I/zO8HMp4D0CceSXTaOht75kz70oMX
rrPigqlKYHfWJR/e57x5wODEcWrR9Ubgcu/332bZjflP0/k7htQTvFH+g0pDyul1
0LDGkEAY/SxhA34DKHDSFBTcSYatafbbfbq12DItYN7U/+f6B9xSBXIY23xtXNnb
q+VOS80zXgQIk2tPMb+yPvX6n/kC2yyHNwpJiJ7a2KD7ojNS8XEs9jj/Sr8dIp+g
pUGZOIz2V+v9ZLSC0Pnl0hpBdCwEsoGko1pxJKUhQAfg+ZSB3IRM6SA3H87OhKz4
sfwnpljtKkOpQeO1CCwqY7YclEgFdxN89+cJOlkBiANDoj6NubW/0YEDvJ/yDtfN
W7Y5K9aYHrRib3PDgkFM97cpzdegnNtT7fKhy2CDrWwsFm99HUVYZ4nsuIoJQhIJ
b4YpZAiGBn5oVkosa7A3GSqs9ap59xN0PceaQrHwF06W8OiUhV6CmTp8olvBKNXS
JE6aaePgKXtxn5DEQ5m8VRq7SYk69SpI08xxWzt85pHIYjd1VzOq45pTVrXX+nTp
kFxHNGmCU4XQbnkgaEhMgYXvg6hb6/mt7FDjWHDUNaIMfNU0XEizoT8Dzw66WgrF
UxxvDYxHNNV18/arCcFj5nvEgTrHxYXmZRu3bjWFYip1xrkeKrJ7nP3fbn1mpmul
VLrHSAv44nRlFSKWjn0anH3ovI+VCtXXWy6Eegh3AYrAz1MWopzY/Xyr7XVuqL1p
K3QAj/KQv+hgH/XmtNXMlnuoOYPl5uiHQtxA66ddfBsjv12xzK0K/6iKOhPwZ97z
4LBW5B6cAqPG4aP5MgET7QR2c3qYx7CqyapAe/PukdTgkzWlCJAIGENoW/DezqnC
QmNDzLfh25DNHjsydOFSAEUSAp14B6uslqabkWvrOEaM9x0SF9BH/kDNvV624txY
AUhdEWuQL14K5/p96AW+G0otKw7+qBPFrlkrPTvldU5yI+8uckCZx3cowDhFwqf7
46BNm4nwk1moq/sI4l/Pw9b0qg1LOoKmrNMtkXPOLul441kvU/R+qKuxaL93DgYx
DbC0P654CRDJwNGNB7qJ/v8FEs/JyHoqJcY8orYtyzUOe3mKJjleEBsUa2R6DbIA
zvq2GJrCfwce4iEc97v+jkFjvprPXG9OjOl+KPdjcCO4tpgFQhNlnOnYB1+3gUTH
VcGkF6GROONjFMBaOidgVxKnQlZQfRVkcrfPAOoLXGbJPRmJr+aEI/hcSd2CMzNB
IzTUDNP2qThyFqZrrHDzyfnTJPgmKuxtSm6MLrZ9lexVbbEVrPsrDIJGhwd4kRCm
Qm/ng/Vr6/GagB1xUiBOyJqt9gAEJqSQwND3/qT6J/3A2JyFR5xTDUcP5JizNuAp
NtkvGnybYGSpf6kx8m2FUZrJAVMU1qrlOCZuUfHYTPICmK0VP2v4a5qrJ2L8td5P
j92DRYw4NTXU2FLVcfaL3Ik8LL8RZSR0Jq8mjLs1/yit0gGONgfXpfk3xZDeR/3t
Sv0t+WiYB20oay6u1jAgwheUIoay7ebNlLUcTeVRUpvAFPRKMT3L2WNC3Oko/xFL
bQNNIKLNN4Dbzt1/lFNfcu3izTHZPwWKP4pq38md2VhXN/GKIrcJhV+vM8bytP+F
HoVaN8mX/ktPQPOinbuvEBph+fzGs+I4TV+LVRZGWojYBcY0A+yO0+GsbtnB1Kpm
meeF9hxpwFdfGagISATEipi5emoZdXzhDZsrMvDRw/+jo8PxG/0wyBXA/rcjr0Fs
2pP3JLYA/RN2suZKJuKEcslJqCmNNicVPgUNnLdWrP7nzCFLCcd+hkvzDxL93MyE
kNkegQM+kxec0iBo4WWabb5AgkqcBVZc/Chuub9/aUqou7PkSGvzv35J5t+BV9+z
5JxqaJZt3Nxt/LSlgK6HGA8CtnPOtYhP/Kr7glOEleC80v4GG7Z5mSEf0l5BRRTU
jhzek1kBcTuanSVFtpbFdc9slF/C2klqjpkxvOvEJ1r7+MNSDo4uOq0MqAkfN7f2
zVYFu9rd/WHwlQj/SnckL6d3ci+d+dhZXXKWLWwldhkb6mGJM7bkbPAgflszTXHS
WdVv6ABW1+5Sbs8nSTth2BeiVxxIjXAM5VF7a8wUzeS33I2uQV4IN7iHC2KqJhrF
nQWepACW6NbaZC4+9Gc7l9hip9BHkBMH7cPw0NafscRbi0aAj0CcKPedd3SIcl9a
5+kvTEDXJk28yJDb090O5YA0FhIzNbk+zhsq+3ZFnDs6D1ZEy70LIc+zj2RV7AWT
Vh2vBENzD1cbkjbP/ZizDGmp92r5NxLsdg4JYV1wg/phHKgIw60Cv9xmiHM9/6YX
zwRhLrfYUMAjV90aVS1bjXtRWqcHmSRXqkwsbVrUyARUs60r+MA3bVXYHLzV0vKG
+JrBJ4I18Gr48Ox9/AdnGavusLLPEL6giPEMvhvjNMaVQtQKZwcicgIiPoSF6xP3
9UkuLTiDViQRJqn1YG2SkXQULNTA5LiM5TTAl5GmwGNg8C5uVpWlqtkC0XS7nyG5
D5dTxle7OxcWqdvEO8NQVOaFPZVfYMOPgdOvX5laMe54nqFEir2TKCNtdxW8TQqH
iSGVHhX3w4GX/h0kLhu7fTOz0kJnGgNBejFiG0aV0kjXTtKoGsJLE3EAMGfe/egj
VD8ae7YAZhb+K5/uo6MAr9IncqU1l6rLPq/tTq0qYAQLUgZJAph8L/ByBcsIkQkg
m6OTLxdhVIGX7Tg8GbuNpvn+OsvIDJ8a26eGP97vZXcqBovin6+Vb5rqsaiGxcXQ
2etuAgjaVrMhYYaAzatOHZ8ATWjqLmhup4/c51g6xHv1oc4KDFqrnFIKXsaWxDrC
D44/vatDbVK8QyKnnirWnEVzpJ4IrniExzSn314MAl2rWCuPEMJ7K51rP+pPsR1i
iA2troqAzoDZhkwmVbOBQd2zg6zlnZzXCs9+7lDIfHyyJjEi5BGr499DsG86e27C
H18SjyzyphkB79REos2NP8j2Jj3zidluQCcnWfyglNETiDgIv/OzbrJvAdg6ARe0
jrGpJw6qtiilceKdOmqAD5ybFKpqr6m8BEfxPw9W+nnxNThqc/e/RsqmpdC25qTX
EpuJbOQiiPvUw84SFnMV2l8RVDhSp6U+qRb1kZFDJ3JbZ1ZXHid49kZnHt3E+yO/
acI/yZDxJvsAVe31NPLqb3s/MJWVzVQvFFT5/kumrqg9Fbdb9NCSebC3fUrHHCyE
VFazDeDC5Qq8nMbq0bmkb7hMQdvdEfYgV4jcVYj0nED/CL2X4OTuZF1vdNe9BRGR
yEgrkoRZw1gZFNR0OEqc8oEicLF0G3FovEy5bYa6aDJaoImqXKJFV1JSpg5MHG6u
zE2ZPRELzzAMCDe+tBojsbLOHfqKjMjqYKK8kqRdM+z4enAGxwpgDOHM4TYizWsq
gqq5pRFQD75RtwoxrF2GdoItz44IxGbgsrwfWCbi2XW3GCuXhc/3FycZOUr2hAVx
46H0F0TRP3KVejQgpnHFxlEuY8eCvjbprbzJUDTNz5FYigY9H6EgJ2wVqP84LNQI
UJ6Ai9QvNqLHvfbAvpEdSlNNgoOGKsvVhEyuTTyZ0rfbzJ76K4vFJjMYRp3ftd/M
cKHGMSRQdQ6AtQv+GT0D4oDfvgBeq0Jpbe3tYtxPVOkpBiFmUQsWJ08lP42jron8
nt0qwcqdB1m2hqk0Vj3KK4pXdTUZL1OosG6nd5+9H/PL4XJo41QfGdxdQkQDP/i0
u0vOA8kQ30neFBZGaAQMejrvugPkN6TJGslMfzFFv9wOzzt3gRvosl1Be0deyqWc
BCZF3exI4FOjpJt1q3oBZrkqy9s81dwtZL0jObPOEWY=
//pragma protect end_data_block
//pragma protect digest_block
VUfcHVGwWmsLUwOfmngTFtoIg0I=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
JtF53LnRg8XtKr7lkd3f5l01y+QEs20y1FiBW6ESondmwMCmLb8An4gUgc+la/QJ
IIRT1LOlMxMZlvUGXCXKgxoib4un81IExP9W8O3ClYSIujNjtOr4nnQ9Ssu9HQ+7
PzoqBx3aXzIkB0i4060ynrUmh6/bgQ/QBuCMOUd9QWHbF05jY+qFwg==
//pragma protect end_key_block
//pragma protect digest_block
NNxYt+CE/9J6I+Y4kSyKaen2GFE=
//pragma protect end_digest_block
//pragma protect data_block
p6kYRmMEUNFGjCyWlgprRye6KmPxIDzuk6HQa3hKKniD1VfyrdLT+d59R5DHvrfK
G9J8QcqMRaEAVojy6CmK18Ptn12kMJQ6ElIgHp80txGOl9Y+QrqrpdkBpvStQsn8
aqfHVGcBYXQ/j73Lbbfq9jNUNRpqhMW+E+kAQXAat6aPNmvuFGUBLHZBW29oitn7
IxqK22/nHL5/4m3+PJoWziR8V7etRpcYPc+BW1Z+VlbdTzEIOalpasumg7EpFWOr
ItPpe+NyjaN2lBt6U5tFXr9Jh4T4iiP05tg4MjHJ2//QbooE0cTndd+BMsDqHu3i
n0dY4XMMAXtY1FU7LL4+Or3bqIHNGncLXlQijFQ8X0tUt8spT3fmo6ySelF5fqhd
+Wwgnkekenw9/PXJw4Pk6WOm8n4Iml85GdIA9xiGN500cduxB7BiQ2gDPDvC4aOx

//pragma protect end_data_block
//pragma protect digest_block
3zijji7AsCpuHXop582lAD1L29s=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
fPfVOABdYTzbYWuno1jYMHpc0LBhUtGSLM3/BG3+S9qDrVXHliTbHcVUx1/l0TiP
8U9NuA/L1p36JpDU+nYWoTiwir/WGQyHtNdR0QaigBrUa9L2Ymd10SgQ7ahBTH11
xBKROIiQx9PI3uswJIYLk4RXQxI7+c0jw4nRxxQGSXKGcOCP+/ev1g==
//pragma protect end_key_block
//pragma protect digest_block
lg7TTDzbMm5FAw35iQ5tUdDa9QA=
//pragma protect end_digest_block
//pragma protect data_block
AKdmk3LIq59T/PhwMbnEgWj9cpMKQd6LTIkeQpBM3mEg8oCBYYey1cL4bt1k4hdX
O6laHl8qNXCDowJtw0qpHV+lzUMYR3RAPupVdTF+WRAWPtxRcBdYRiqRE+UDQ+oV
gtgqwS5Azq3wFpvBcP6qMZyrzuvi4ZQC92RmzN0VqML6xdmQPaYBIadvWGMzIZiQ
E8G9wK8nc0uqw9qgl2yAOHzcvrHhdKkvt1uJLZfwcz2eEgkjtc0HnkPhsJ1PgADv
RK5ugl7FPhx1dncaDakj+xmFeafyLGulmE2cAS7jkAayn94Orn/R4cHydDu5M3RL
SMFe76nBrFI2/Lx0sayAcK/QRLWAdFk/Zl3kyhbtT44SLCecRC0N12sRGsid176p
r81gdx5Pdlt/0SBt3remcMaYLC5fmJ3DnUrx0HlL7QrB5i59ClHE/Bl3LxgxVFEt
2PGMcGNnAgZqNOjvwXM8lcqFGMIju1deJDNkw14jf06AadSfApTlFIn8B72eVWLQ
th9aeZNytaQx4231ydbxU59yS6flN6g3kMHw3YE7uQdYfD7k34DdMm8vdPhxAXDw
/9YugNJNvkqiGl6LqM1j3n03gzMCpd2ubKVFEvc26vFozXBmwrm5QTNgAAdktkxF
MeyIhaA9ygFHFzOKFp8HjoLFhOLkUjw6eDh7gVf3bQ764qi4av/O8qolX9CZyzZr
F0PAba/l8OIP8gUqOEyOU1tz7Y/t6NuGjJTZ1Aws8T7WeWNFMjVsM52QqjmhiWLs
B9VRBvU+F8d1ALN+HFPt+nRf8ugkX/B2BDQgvJyI6egSzYrBsyH600TAbTKmsIp2
NmJ4n9f894dGofUZDrwVCN3iH1g253cgJws4F7OWINtEyg3FZf4b/Ht5brqivUo3
QlXbYd1Ioie8d98nyeU/czjLDTVj1juKua6tdS2cRjMcVEwZGZuEYOf16kEE6Ot1
l/V3xdqs5XmSuqg1sgIoBrBqdKGfeuBYV9B9jCeh52FTsL+uiTrsMZQRueSny1g3
swLbDHpH+3xVfDpukbtv74U4QWHX/yfCdroVtt+QZoXcDKnm9irP/GNL7rhBCHA6
4Hk7yNAL4yb6X18qykW5Yk4B9Y0fXHDHcvNWARZlAxpN9YvwwpuC0nLCH4R+PvUa
GEA+T2Q80nXxchCzXYJd1IPGHvBtjKqtqCWMy2uFPlQIjwllZ2GgwXBoI/jabKiQ
lX6NrtXJC5cuIQ1IOVns+OQ8lsIU4ct4M/ohXSwhDAgbiCNq+5kYZA8tUXiLmAXI
wc5bIfCnUp7bndiL9mJR8ciLzBN+BRC071VXM5syIASi50uxyysiY2Rq5dsv5llX
YfT2kfE3f22KDsesXkKbRtFhEonMMuXzR6OR/75+6t5WKR7xpWv65/9fdcgqwSaI
44xDa/vf//REWGF88IIE+ks4giGOh8y8+5sKJ2gBMQd92iwJztGWyDNC0JF5eIj0
KWqCqGd2YLNHkQu1HHnEkdQjPFDdzIsXqE6wRYvxcSL2N1G7S7I9/44UQB8POHYj
piNT0AVAWjgJsssCNcGBDOo0sshKbh8RYw+KKtfB/CuqW0n9T7kJU9gQVu7+u1KU
3fyLzv3BE4d26CGN38hhTzXwD7vMDGEd+trnjnoVnMYJlyvKLe8pXr5wp5UKUBnS
XuCMvxdBuAqM46BOz9Mz2ZuwGdloG/QB7aEukofbNKZbsoPah7WMq2yQxqKR0mjt
KJR3WTNMhCTGUmL6sCr9LFInG9o94BWRTIVGU6UFoXRIc73epd3OErvPWZAZ7u6o
cff25YM58bHR9Ly78Za/Oy5KApb8/aOS5sRiuhHJn9L+0K/fpqnPdqmhUPwtHJEr
G5ekopdPL2RnoETCZLij+kJRSMCJ771lWxljfHBXyyVd6Sklc2vQtUsnKYFaK23j
8cLaFsilKbRdbGGBKNgdISCQ3Tmv8/qRnnJSS/R57a+gZSSl//dNNXh3NHt8AdLp
x1jQ2m3b36yvRP+3LO9jMrcjPx/QAigD8NGH6CuxF5r6kd/Dxc6NVUoNRNYkJtrU
cKJpUxK7VqJ79xC3UgS98vnqRJVMGuqEbwm5XbqsQ0qMk8RSZ6BIqNdGRhI4+eK8
UIB5dC6iOVgXNdwWruWi17GdCz/vQtDhXOqBJwHn6W5Usau0pFUH5yEh3dsTvona
7Ezzvxal0vr8vPWjk80wq+NuE84tYgh9rK18/dI1OMJbHnQfXJeV9v1/dKwcl5aH
4PjHEMvW4GcvjYSZ2mlub+o/4pRUV5Fib2coOxQR8cWCzP5YHxp+wTgQDLKlXgv5
qIkZBXhTtOBLmv7iYCRxOPwmeJxGJOKjo5c4nrBj5uYoHmNoaZVrU/u3CsfVRxF1
LWtyPSg0pksha0YJslEenzGBfsy8nQDugURxAXG4bexcFulFZY+BpBZ/2jsyGi/L
dWpOVsm5SWMzMBWd/vbQz6+H4CqlMz0FzNOCJPBuArp+lKHqB0pO0O4iH9+YRGcs
xj7abI4MVeTLFTyasQSSzCh2z0XViiNG4y6pvXc4VV4V++GeUyYWnZ1OXQs2//dZ
oJ85q88nMWOx1ZUyF2I/43wlbNS/5zUVh2q+1ZRbas6kgSTReXLWy2W+WEb4hj4g
6JC2GNSdOzfXHIJobg8HjzZAs0k13wyrBxr4aJk4jR1cPamg5dTlyVaEVdqOdAhX
/JNfv1yi/YQ6s9QNc2hEsgD3zuUdbTXzzTsKbor/tAAt213VMQSp/RpjuSsyrl4q
bB0FJqaesHT3qw/Vn/giVULSuvjyk8yYCzsnFhYIPU9Wf0XhlVbUpcqzm1+YkR+u
lMOYBC/h982jhmhDQT15gMJHwbsN5JIfezgGijRjcnugJwN167a/9xv7aTEMBnel
trimeH9yJ2R3v3ACXbRsEzqjariPpTO2+VSZBm1h7g5GctYslpcEfqlgWXgruSvJ
62cPI8blE+DOo9JZHwxwQFUNMRpBgmy2lwu/iaLJYPglyla/PCK97qACzvu5fFbp
QvT0CAU4twC8URKwNJcPgX867ZWMYT2eHJVrKWewlqL+aCgeuBbBTSs/aVSV9AcT
TaWLadEYqIESs7IUsuhuombHNiwtvZkAGrNVm+/d6UHMlGYtUkHaDO/x0+lq3IqL
QhhMwD7mCT5PX/L8uBzwSCuCNn4UmwUq3McKZ4koTseO37Y0eoOar/56DSmunTJg
wdxGoJAhRo4rcVfYFQCHuRuMeC+DLYQSMqCkQcQzRnRQdGwx7z2b2RBei9yzckwt
Pi2WfNs4jU2SLidzjBv/3h7toXIM89uT4WsckpQkB+OScAs2VM+FMZcdIGy/HvTA
rvoVTV2s/DWUrIDNGtBTzLAv5hZ4QmKp8FAtnoJqECDFARuZlhVPiLqVs+A38j9+
fEvU2OKqEf4ZjwMzttSghZdumjTFUcSuQJqMspaVNwyb/WEk7W73viq9zATybaAJ
pb2b3qgtaZ16iqlKd1Sv719m3fV8bwoeRrdTZIjebr2O0iXxoUYjtpTuj0k1t7jk
iSy4dkpYjw6YdegHd9PNhfXDqc8W0QnTSzdYEdQGwXW5aDS47QBw5/jjykCCahHY
Csz4bGQBCwOklM8/CZk+ZBBI+UWroLFJLkksN/BFEbVJtHVDPze3CkcbFvUPW82j
BWy+9evJ5Dmv6OA3W5ZTKdfRCmYycfKBmjucgeYcjp4L7eRA436HBm8DnwSeewol
5eC5rA5sx/7LNWrMdZbFPrOpoymh9AxxDTzOWwRzcCkOE0mKgguFCPJtgLzqJn1h
VoxpjAVV8swZMy4A7l9lPuGvRzuH36uFFGhEya3QW9ljZ+J4t6Ns/rPC2pMwwLvj
cBEX2ceE/2DmOcICwbcMJKsmHn/chUJdPdE9CLMB0RrbVHAjf1scHD/kIY+vcMPN
nuM/hORgy851S99wdJGSq5X4mJ/r+hOGU1dlHGNY/5pHYwKwQt50JJ/5i8BCWU+v
j5fSLLb3O79pB+KdFOo6pPaqk7SXSftLiNvIv+lqFXkYEzflrzI83fou6/TqpjRT
HBsklfrczY6enUwvmxiH0rr8S5Eb14UgYdhjL2IgzmPqNue7ZZMxRKMuGR0QE+Em
1hs/s2L+16rEw/qXgzj8X+b7UK0alkA/SxDrxRj67gyffx6H2q03+wqEFXB2Rvoz
9wNDYhbThJwe77lXhyshJElr5ycGm4do1J07NBs9xOU8w9/Im6jq1JEhq5b8g6y7
RE17hgbLpG1phB/HmCdQMOUR9f3AeaRI8CDVSjW/9N7WYn3poMfFzYl3IK1m1rNB
rO21vxB2PnxL9XPY3mNxnnPSPrsvC9Gyd+i8jqse1zvEFIAi89KdtAAQWcsd0sAh
SfmjKdLN/g68swGAC0ig87lrMrhDod2htDGQ2Un0SSmzP6MfkhBy2eRvfeBlZ6JO
DX6NAZAmWc2SLpQcNB/vgUF9L5fJwJI9kgQMCTwDQVuPrU0CnzU0g1vA/2P2N5Fc
spA4NCG7L7k/I5mgYxgnWd6nngSEOmjwR6SwyXdlhvWRE0T0eAPfb26Vxj8T6g/K
NMsGkLDURqsAJ6UsOunAFdk6yeUOjhBnh6CaxhvwYZhglM3BqAbfjQBYDRXF6Rrm
Bhwy+2KZCcO/q5S+KXRthk7qTA+P5geOe9q7FT8JtJC9tUPH/PqCDB2mpjWH2fND
+sZg7hAVM/ZhzkfpoUh7JAKbOyoXL0JiQGBYKMm4xOekTfi5qC8C7xLD8ww3cuVQ
xx/xxThDYjQy1BxwSSpIZkG1iP3HuvDPAI7JUc8pZIypIdVwyGnMm1N5gPalOPfS
PaRBmFuzY8+0BotGspUBGzAuVSj79QSDXd1LY2uzvJ0xAS+RQXiFsSSTTYiByNIc
3DD1qud3qvDSzvPtzWocYckcmmvGI+94uZPMieUfGmCYCFZJzcivzoJF2h9Vc46E
cTrjRfhooTbOnwEOCVaLPPNFtJwLhKOa2xkIqNFTM+jGtwpoFTj4CYMDYTWHvYH1
4ItYBr7FsQSkxyAE2dHSKMNUDedf3YdEhgQdbnYE8zY+y6tjUT7BxChWnS8NztH+
Cfvrwma4fTECfIHpdII/W2E8kxByoZKl+2GTHd5YFh6dxur+5dj7HPhPPJh3Aehy
cf7gP9eR0m3oRvwItaxj0ND5FfIrSlENal1ylBezZ9LAVtB3oVxObu/QRaM6pCTc
0HlVjOQurqfiPBrTOyGovxltlzgWSGZjnVYP6zk0/4OfRd+Pnfr1JkflAltRc/xi
ISqW3O9n3LztIna2yQYIKx7bU/PYHOPPXwAXYEBC2wJ5wFQrsszHqgKJtbCODygI
JabtogAk7vvmVekO9aL+tGXKQFw6B6gPeM0rkdlPtz97oQv4uCSD1jh0zzbsv4Uz
OxzFVv4gxqKGVggZDfuFWX93TWCyZzAkGsNFXqVRyN+i5lAtpFxsYVHxQY29OpMT
TOBTFjrsWl6ZwpwparSijUBKYsMB8ZyiMiwWa1ZINSLzAdAWqNJxTldQZGWDGn0p
Qh1dW77PCNot4czXIvRJBsUWhLqQbkeyQiEVYCt1XBolSP/4nDGKCZeBUT7oEhGZ
aimXDB1nTAl3q+NJwRKgUmnCNQy6m9WD2I9y/rJ2r1WKRr5Yibrykyy8elq58awP
qxA5ZL1edwDoQ5yd4IqhYb3r4/7I+F4MD9NeLYcpPJm9rEanXHMd6mqj5jlzi1Yl
1I5tehvLo9pSFE/wMWyo9XG5J3XgOQ9iyewpPvoGai1M3pSF91E2m39KRm9zBW3X
4X3zdFHMd0bf61+fdQ/YA139Yuiydmbwcv+XNy4njZeCxA+dtyMMHXYXHpisKvpc
HhKikMYcWaWMJbAagR7cC/BgEHqdHfEySt6PegYc0C3hc92HRWpFZM54xdRIU12e
s67W2UPZ6OFURnG0gim3pCjdmMsHRPdDvBY4wXqqularulQg02k5CSr21zOwypEa
y6NowT3WV4S3WL1R/dnIt6dqhwbcriAnBGhl3JKTURt4nYgCrYyqIOx4hhfk9IjH
/puVqbIKWl3niXFH6iTFAxChYCpqTUHsPWfZR7d3psmoEPNkvCAgGd4/xcPz93iF
YaCJHkczqm+QufFmUanImvNNr5ktK2/clr8xHSnJbhynNB6ZDWiYHNfqUdpx9tbD
Pnc/tigRwit4VxY0sWs1sWCZZir8A9HBbmBcWqBLPk0HX6+39ZUHuAULkv9q5H8M
svJWBti+4q+RP6/13XsV2rfjFV+0UTixqAGGxtxmLTKfKzI3O2j3NIpC7S0kTLhd
S+m+mS4sz3Eq4/7YkFmZRirFeE/mRb9hlYFGhZkOzic+FFpn7j5gG1m914CtGcuW
grKbY5/4tFlV7jwD7bqLtax6ElxAmqYfIp6STybowB4feEPwJDbZzQpyZeTVcenV
0dREE0O3R3jwIF8kbeFIWf3Nk1F0MuSizNsfz1ZuaKCMbkwXZwTuBCE8trvlq+YI
Oo3sM73s6/fffkqVFfr/PhHKcV8Q48aDVKHxXLen6/p4FtDMavRyGs7sdOEOqINT
+6noiC019hM+LTxSkTts/0ccQn7ANucDmw3wOKQHMdQnAQVdnoQHcJxiXUxWPDXM
PtqPdjF4oV8rqTFFs8nzG8yS6OlB07B45/k2F9OZ/7Vq5joqGkjg9CspRZwmqsFu
ahQD0+3GXW7a+VyN8fJAsKipNIN+OIoxXM0SGcVHIqR/TraNJ7UGxUDmhAtfoRFA
rGjh8XJbFXCPvHCKPAQkCoEfZAE2raUqP4crJWn6m4fEIrFNYAuVTrdvaevhHvnk
pdUo4oYPLlOvREeVYpwkZ9Qrf5/+AVsZgDCmBtqOKUBVacEy2HRHof/VUSC7kn7Z
6HsDua2q7Tix4jHssrqa58i1+1yOMK22/TXGnXDmsYfkQyiCW7JFtN5xtyUcY81i
hVf2DkSbIWciyJhER31VuFjNy6xD3Da2iHni77zaqQKaGbBnYusgApEazjxve+ue
cUAKGg2i7GHJ/JikmZrG1wZ5ewXbrUNgppnbeG8l2BLUjL5HE5ns8b8ROhgXt9eS
Aqj/v8z6J5S7ct4x811JQmHze0HJh6x6TmaHqMlolH1L+wuoDjTtehpOFwgyDagx
9P0VIB9dgb3mMLcKPs87TGzvSQEk89kLxACDF+/U8JUZCkxfbD8CMZBfxlLXgMI1
ZJcvfcs4xUbh3l3KAYleQGkppNRvRbjPIxalk8ZbmtoaJUqf1ZTT2nEmmBxgj7gO
K2vzRRear20UFSF0QxCJH2h48Q2AQuhxRaNANzS7zU0LRhwWWdgNe2v37sY1tchL
2sbdH0ev/YrCrQbxCrgQxGR0/nuvOcEZ9z/F346w3KLAdczf7x3DBPP7eZOZ52EX
HTeosXVUNi4R5y/5Jqw5ADRKO5gB8Odxbx3CNoyjKoEkePlC8FGlmpuE5gQ7EfUj
rGDMm4VC/F7lbtM6dVuBL4x8BVoYF/fvEmITUAGmhInC4qiWtlhavXylHlD7YVEN
rn3dYTn8fqWMv1UMEWNtA9S2vvjzf41hbsdp9qQkUuW+d5NGudYEl0p0IVgr1hA5
Ui2ypDyxvdGrhDKJiaLQXTMvu9T9O9tCC4xfTknlN1YHi8oaP7d9tCrpm99SrV2p
zoP48x+o9VmUrlWUdEd7elaR+r6Tsh279OzZ1Mg02vo/Pb/N1mxxNh8pHrI6DAP1
LmmbV3noYVxuhg1Qrg9B2qeUA7+dvj0qWYD9VP+AYW5zGeyb4d9vBKyfZCs5iLo2
QNOZ5IBYe3Lo2JJmbemaKOC2lWlbiZyjp5gPlYTs5/qoHEtviyir8PVjlzXGWnkq
ed+M+ipunrxGA2YkZijNPGd0hdBd2sLERa416UVDgqUSAJLdLC5ZmnTcIvhqbvxP
SwqV7xH2sSUi/qAFop5HEa+PkLF59G6M8MA/XR4YtZH0egTbESk58AnMMwBgmlMT
vGdXAfr381shVoGgF5EyogZqV4fasP916WO7bA+0qmALmm6MAKfpg97Bc79JPjeK
Xcg7Lr6uSH3yBiuq5qKYE4NYZ1o+PCjXnBcWFRXPJ0MdMHOEE7ZwVlYsoSYM+ZaZ
eXurFVrfmNpNg6A1d6s+blLSUyt+KT6Okxts5yM8hQEEGPCXNFOXi9Y2d3nvgy3Z
e91nt38aWfmqjzDkXOF41NgfNQVPuNEi14I8Oi9Il9yokEzoSD5VivMRsEtE37EI
ayVrZwpxlrHSvo+qBxFbVNlv/qvQjK/Xon2KRRGtUgWuWQJ9qZ0W2F+7/cBYk15i
OiyaKMbDrT0CwMijyLxZjxIR8RBIUndGycjvN2KFGBPC43rD2XC9kYzkYGIDsT6J
LHyHw8OP5I25GMuxmOG0YwjqOK6ia1v3cI/XRyqWMh6C7TMSY+8KPXTweSpYjYDz
5JIYZPw5yaz1ppf92GXHA7XvHlQiu2+C6d5CObKrxbElS8KKHzfKjXcc8KhzrQuU
JgjVR0FTwxQESkABCS/V27g2cDmfB5p4Hmffgx1iR1e5X1zkx+ntEAfFLT3N2f+z
PSESbGhzFyp81fP8qr1cikPJDYW+1XRV/qRMX4yseZNsYKNn8oKkH9af/Mfflov9
Crf5P1NeVs0iwJdTzMuJn4KrAgAUFXKCinLXLUMY3I8PUDArsQ8iTrzDLiIq81MN
Ns+wqUdQSpEmo9IHe68tynKbL2Nq+Vc6D3LZepc3TN7Cl6Hl+9rGsdi80pIx7W8g
UxvHZz6E83oGxldlUfYISjYtLBPm21rN14B2uIphsoNF0rhTHONJD5WMhM5AETKu
0uc18AotTHqtC/gvRS/+uf5U7l44qTopzQ6as5l9gvGbnpLw4LtoiCscguUQpMM1
WK1o/OgQMjRhx+p1mxXBITTGxm3+SIe5sP8tqEiQ/UOd0OUKQWtbAWYnwVkEKGDB
VGrzWPtF6DcjHuLyOpBO2FhQaqVgCtayJkNnMFV7oBBN6KzmZHSOZoNIzGpY5FWc
aZ/yP5KCx6XjASLWRIa4MZer0LiXr8My4k3O8pNVOjLNGEb4P5d4r8eNzICnxdug
F5+MS+XDUNwBcrGVsbq/PrdcRpGErPm/Cavfuz4jkUZAkrkYq8fDJ0gX7ekf65B5
8EgzBYW1ytH5HDyjRhHGL+jdjxZLfFjwhFgZRl77xCpPGaiV4LyBlSHy/o8uD2rQ
nCvvA4ZBdh3/D0W4OydBfiHKBgAU5rJm6OT0ZA5AB8FWy4WGP9MXiJlCvoBOD375
9qjGdRbozlDlw/+WIzrThEHXgbZNBwRCgk43M6eLtCeEzqTDzQg2Zywwx2zWHQVD
PRQ2W88q7DwA7TebzpZ+yy8HT2fd+7+kE1Xkl8lAU8FkODg50r54idopqmdQQr+6
iLINeWH0S+a2RFqsJh3ANQzHwmD1WermSMI3jn6JedgX8wqMxfITylMiWTPFBnWG
utQHPDAsAof4Ymgw0/4ZGK23TtKySx+E3IYmgpPCBVCWgt9lSECK4UPk4dDDdgBt
gg8/CaOcjdECSdH4dZJB3+USeR/asGb1XBovEezaky3+C2zg4S1+Xw7tWNGHyPmf
4hJHGq42YbYt0x0JR0RB8Hrj/DDVXvQM8UKdBVqP6n35qQAFWrBNVcSRA5K6w8xx
4sjwsHoO+xDThvDf6PbuUyv1l0tlf2cgW7lA1ZbIqgCJnH9RN3hPyazZAsNvO9th
1NLPx5087Npvtvvw8X8BWqTJ3lYOfV/AxBYvB6hPgNaSkCqXdNv+Xx61otwgfANS
WFMqQBB7YnA2M/hP/2esF7pWO9UxVeGj61ysJOblJICVZQYuvuXDnxHVSsSivVta
1lk4/vTwBfcMLEDq+HP2WYZ8VelONbwLvznWSKX0fDALwYrdHU4xCkLZdAg4s+F1
FVXVWzQcPKoVjbLzp0rEel6OiBc505DvegkjjIj5bOu5jjiZTNP85FHN7g2gEvtd
wDLsFxDniFb7LIGfa2vPWBB92g0qOazQe17ICSS7+CS+fz1+9ubR8Jy7J4esPPpx
t4WTLKD7R8tQUCXJTj42bmwrusCuk571FCo2hhJCd7ARHKFpw/w740Cz3QCYkZeF
xFWo2TkrlGXYUBo0FtuX9IJLsrApTODTbUSw+CjTkQb/Y9DuFsIRLFu5CI5cAQM5
uXDGxXhvyeRt7zkxN474+1d/5fiSWDBD4YfGQTY6AzUgotvBrxiLGcOzG8MKjJRP
Is6dE8VJdzxlkUT4KUXyxdhfJA8LLbzd1cl+hZlMiLIW44dxKcDxto96ZsIOhzKB
IdR/efytuNXLprFNl6iIc0E/9tQQpW2z6nPE9qQN3XunlS8PIMRC85+q59OzKmSr
qKFq+UU5g82ZlIMZeOGDS+N5dDkhItPBOfDGXm4+TNN8bkvc/xHn7/8QWriDK/Dk
wzdk9chYMmcwjHSHXEdyxh/jFGgoP3X+FdN/LB1eTcbDpksg8nxQ/rZf+4SIXeDf
SIGN8cIZ2ilIL27bv7H862iPAMJtFKu5dmaPhFhokDCzq4k6eCClsol90YSQ9eiV
stbjDk14lmvyH9gcQzBOYM7JGdcteHlPyBIzSW4cPe02vqbgzlfN3NdxaOYqezL4
L086qsRhdO004FPh7mYRNCkkj7lJ04lfSES4w9J7/sL6BLzdV3ZPjPew2RLvUs3g
U3smbn9V+7WbPv7cZmQ3vFFMKtKqb5tvdHx2ooudAQI7m6NKfWAUWs9wMG21Es/G
/48xqG+NhrZ9W8J6Yc78ILXu+gAASf2nA/MZj7XEK13tmKpVw09n55KH3cwjvFDG
0gmoSSRrYK+qewDu74mvzYz/Le8OVqFOaJd7K0wAf6nlClx1WiQpsp/OVZ7AA3Lv
hBmRfeglJD7dpyRNcEmFcDbUf/6RrNEbM1MWsrkebq2/pITUZN7RSsTwTGgxw8ts
CIkccGPYQBqc5AcqzFLPPhtB9YE7iJhTGHoz76wdjVrTdjLP3UdIkW5hsTNHVEP9
3L1TpoCdDNgTKJnlou1S/jaGHkBAW7VYJukpZQftRc3ap3qlZhy958rsJUixepZm
BNiKfssqOTTBY0DjR/omrb+1qr2kyIfCdcxiOcaEXnPyidUBCdfHTnaUIKEtHoYy
XppxbdQJ7tnwhD3O3MoiFWd0PjjC4WI0j3ePD4R6whUJxNzxmmjg9A2FK1yFnpFQ
A37jLZCmisEdSDDu4AHjeQDtaoJkfUr382YHG4o8UZQDk+ScuO37KCoKh6vxF66r
mapzQTG7WzjciswMb7ELkH6mI6tu25+YJUlwU2Cg3ueeK/gUg1DR9CiEhCsZHerF
Jvka09cO1iQSJ48wgIsqIK4HJezTiJFj7kd+2GyrRNxLgxDBp1Z5Q6xI3ykWSlnK
VqLCL1YSPZiIVqa9RVEG98La+s+v+447Tf63qHIAF1BU1wvoW/6lI1XWwQ6sdxry
ZhyTZlnbn4ViK6ncNxhNuYGvXsCQn4wOYioIPyZ1vNeDl1dZJGvNB/2R6IcvIGwn
TEtBID+kxyU2NwqL1rl+LU82lE/9pxJaycPLlZIyPM2IsMFjlnieZLSAvvXMnI8v
FkIiBa7NipL5Ml5sBtPIeL8J4PnGYpDnHCmDFo/69UeV3bLw9VpeAEMLKoZiMcgQ
uboDYGNcH/hDyNBMBfHrV6hAu0SRfrWUk43Mrm0N5Lh306II0udyehE8g7sCXy8j
3uteVkJcg6mluFWp0k21pu8Q3wwbes09U95uqOmMRIVyCEZ6GNS91is4OMJdRoER
la7vSPax2975yTF8C6L8/GRFeLp62Mk8PVE7GKxEbnlAWwkTXfWH9A/wieTRm3Fk
1io1vU7e4VlhduLwsyPMx9PS0DIad9hjz8c2z0TW1Mr5IOrCgPPWoLTB6t/pN4fQ
P5ym+kYaszylJ2y6IKgPyJsVf72DrRv7Fa2S45D8Q5kvOAGSr/+pmkVr2jms0sny
mxOEDLDl+2dOTQr0ouZRD1Ddq3rIbvhmSyStuDpBoWDmKO/uAuoH5/CGMJbFAc1o
mF39DEjSSQ1NEPZnN9MhgCOihouWV5mrJ6ICDpeirGi/2+EM/AwHH2UCdcmaPmzT
ys0gSKtU2o+Url12MQb8yXR61SiZdpW5Sg8BSMkuDCjxpTAgsqFSq+bDcJRtcYQh
Fa8Ac1TXEOCFxgUsEEg3EZ/5lNkfoGw1mCj1l++szxWjaFbDcmvt6BQi7B1qKOIe
VhOZXedSjnXc5B/JiatKwMGt8BUQxebyqM+bXM6amrdMGWVWVltt4vsbWOp4kLsr
Ihcyb1oOJABz+HxJpQM0Dxe2TlJiz8lV118FMAc1G7Y8BQLcuqQ+DA1NhEWT+52I
2fm5fjoCU71lyjTs+ATV6QwofEFX58CHMVcmkUEadRD8i/3mm1Ullz5fPv0ydbhO
J0FhwYx8DkInL0jHZhKllvroGFAqPXJFvLU5hdiBJyaXlCk7thnGoJyaGeqBPqhl
69MBrUkP7mqtrKz8s7vgE8RO2Eb1etRmPMSDPRoedZc0Fa3R1iFRRttm1eUkM6Wu
LsJI+iBIymNiBHbGbdOr/KuOdFRVFstQnJBF4i1aUSTOZsvePBa9viX+CHXE6gin
vnQdOHA1EewVUCm2Yb85jHsoin/JVtLn6BHAA+eOARKzIunvbUE6Jxy870T88bGx
XU//N9RDKC+QKNat3jTp5SSouFpjdpmR1lSxHkphex43syTNQDU2MXfF5Z9bRbqv
EN2+P8NScvG5FURZpklcSlL0CN5FBU90rMePSOmCM2EaZ9rqBt9pf4Ct4H23aukM
4k0/4Hz6N+Bsa1qVkTqo6kjpkMJgDmysQ9WiDYDZtQXBLNqyuPWQ21EXUomYvEzg
GegKiRZAA0s/qKZIqY4tsriSpjdXysFRwqq3BCTmnYNOuJgorbP/p+kl2Nq7aQ0D
wQviPjQcCl5XFPJ15Pm/b8ahYVw8ZtjaR+HXpIa9lGvNidHAvu7+Vz854Ov6jwVn
5NwHBuhUy+T0e0cSG9XAE5gzJUzrViFmmBpUPL5PY/JobsEuOYWVUcVeYmLwBdCQ
qCxpogWJZ+sOx0yPESOpz9zNekSBoL9W776T4yEj06PRUPgkqowViH3ws8YRcLDk
IWV9vnlFQbjOrXL9EVhJmMU2NHKGG2RbKxGnOrVO8y13kDhCBK8if4v533lXQzH3
f9dfcz/L0au65BbHvw5Bx4m27m72omRRG/s/cZ3iNrKIOPp1BC0fEae2BdzlgumI
YdgqCOpIAi15MfW/rEnLZOZjBf8q2TTGN9C4xX4m7ijd2ts3ILWK5mTudFmbcp45
YuXWeL70tg3fKOZWaaEWqoSAxzYObK1fujEvvo8TY/AL5romBTm2cAipCWbrHQaq
JkXbnP6WXfkbR3VLfRajk5CdcMCZiinlbZFes165cFiWCbGWcWAnFLhWxe6zSofP
0RzMTHvWHR4NJjZ2MA7/4z48zILFITmRS0NKPZIsTMIL7RaCN56v/gUlYVybhIsg
QZRfEbmRw6ghVI75pEmz6e/T89yJdJJRtbQ3uLT0jcd/ZAiIa0k3QHTbOIAdvC2v
92vUh9fnKPBowjhOx0sH1LNtkrqnTjz34+2l4zmnqqatDxnqyRL6vm+TcvKrDoB0
T5jVCF5HxTH4aev/C2xm5rzwn8FTzI6j6IDPSkC0k4k1ziduIMZoRs81kog6+/AU
yIHgIwyjTy9O4uQXGIWA0jkVGB8wV6gdL6m43RU3CxkYWK7ikIHkT887IJP6tRt/
oUrHWON3BuKnuDPUuYw57q3b5vYnedOmhpoJ97u4rx9g+4yNPAiUyPJ9Gfdv0xXH
lcvQwdX2GXMZ2huHQxDEfBlj6biVNJQcb9UlubL5m/pCFoKeqE4wHLaDSr3oc6Mb
Qr1J9Ixuhbz15gvPOZwcQhhKBhSB6DZFuGMLr1VJDtzNWFTt3MynAvzneehl4MWW
C69NvC9aUlTMIUiyZ02wHc53F/UM9PM61qba6btrEtACKfrU1YTUo0TK35+W8avV
jjKT9QdK5zKTDlrwZ9mO4PEpPCs3KFyYD7MDxoBibVITlkZ1bcVIvpKzIpOxoCKj
0edCcnaQgIYAuhYDcpgha/T8QmfilKbGkX2rkoR9eCStP+I/Dggi3bpQsrdsBrJU
usPKabPas9vuXVa/PhpXot2wIj3PU0EUY48YIZ1EKmRj0fuEBBCeisfAKi9qu98f
Tl6QJxxLNOWQDKhjNe9WLiJGtYtelG/RmxwzNPp+lMlUa2nFSj7HnwBB37PPbUOF
zahKu5N1JMO7FMFCLg6cK3BxnPv4ZZHPy5cD5JUkOLBLALSk9YZpjGeYCFJkw1X+
+0xKCBS+BpUT37dn3O407/PTV7KNix9VsUcWp3+G4rOkJ3pPoObuseZSubGGygwc
RaWwkR7AA0axfhD4efFsM2mlIUrH5PzBiTyZpa/1Rju/SeziUblvM592AemV3kg+
BAssKgkgf6qTha5b1PhPnZnxx11ZUJI2E1/Yonw211/7YaGTNb3A5pNGaL3qU79o
WYy4wdLDMmghWt4SWmGiStR+V4AEDAc9SXwVkffjou3qQ+Yd9OCFnjANv3vxaWle
kBIB367MeXoP/oxsc6yOLB78D5t2qOUgDC4yU4NL7u3EDlAMhhbzu0QMy1WwG14p
y7bhDW/AbG5NLk3eIhK8URmjOmPLL/hWWqElm+7mac/Bs4v2qyNbcIPa6QBVYuX/
PiikfgJ+O82zyHFplaSZ0IW77iHn9FAno6uiVAjV6QTneUFhjeNbfDu5d2drFre5
KBvFAPzgGyDn83VRsn3BOsGnkQ8szx42gWrOq9R3uTK92ZhRnTnVAJm5wZIqoHrv
39/NKQ7smsW3jTmz3Z8sYqHFS0BVATeRWEhC5wSD6Jy8Kxbh6/ySxSr/YsESIZau
Jq9jLFGJZQO/u6vI4wJAMx/SEw5m3pUkFihmhebnLIy88Z9AykBNQ1w/Y9u9rsTB
LIf5hLuGf7y4iFnL/1zUsxOUt+ICk33/79Crmey9dRexmYk4RzHYPd97zRmd03cn
AicBAqf88v0EC7/j7OrlGhOqSG8oeW2kA/TztajH9g1NCaHCjXSPuKtqBydyYaeG
8Evy1CyxX3XGybgLuSmp0nl8qU9PkgQkQj/1cZelRt9OD+5jzFLw2fkBp2MrCbbJ
bj2mrVc64IfFNIdsDoAo30eDW08+hectmoEP7DNRtzAJf6fF+/2zSX6hOowFUS/R
c2+oXMtOcV97g9APeMlMnpXsg9xy8kMET766ZijadjrRw5I6+4Rpn4wJ4le8QYFM
yjfthsvnoX8zr5xQbyQkPwsZMbRxPU/UfJhIXXSX9pIAqdKp2qGv2R2AyZte8Wn7
/ujwXBnAAkim4CerhSz+zp6vZMZSvtRGanvzKZ9EVqb8W+66nn/BIkAJBg56L9AX
SknPmeQFfzUg77V+drCNlgcNKo8np3ht+5XZTKpx3sIXRdsshA6wCWcd7nVES3HP
a48xT0+AIrqnLM+lqx3/zmuijIUsPuFzwLagt6nl6SpxHpGNT9BcP1eeqz0Od+Ns
eWNmEkfnMkdjlBU/DlaWDe7yXwyweHoqoLaLclh9EZHJzoaU6rYwhfqG1gaCorfc
A1PcSzkU1bnRd8oFJ+VJZi7hhwZHEVpEIyzRiBSoJQgu8+Ehkx56YM68INjE0Ddh
wAJC+if+CDiffOCdWglBkcHlKWv0to6hMu9BMKrl7F9tHE77hxYIZyumRlUjyGM2
6Vpz6OiZpTvWWXgrmvdZDUdusl/vkpBNDTE2VWAQm71ecTLWbw83WMH/Z+KE3rFT
RwOtEbl9fLjPx1mRDSxkYYTLMwtNO0CzSjPzFA9YWIESbSuGOQp84nCMwCL5fb7N
OtTRy1e7bIQAhRTFNG00RNQP/IkzoGm79c+0tRh+I50mF/zylY76v3F91aqbsDou
l1/LLUlHAoXTeIlZxCwHP2rgiCNMdgmzL2dSxQ/46HtFIN5wT6SAC0qQio4K4Qhi
W5WRqMjwZFmA7amNwnIUBPNG1xoAkxyIcNrPu+VIDnoQNUDkD7WZjCOK8ztt6984
P0E0zI1ei7rqijBF1LU4U1RTKNt/TKzJB1CnS8/PuU/Mc/mT3iSPYMlqY5XhBjUn
sg2nWtqP6iYVlDCcpt8ndBleuydY8d9bd9XJ4bwAvKZSiG4hwWEvYJU2iAKRMuYp
LFV03tS49Y3oef2yw0v3SYHKW7ObbTFbZ2qE5vJnLvctwc5neRI7VpHKswbLSspw
l8y3Yhp3690aiGYZd5JxLn1PkLSfZS9aDhijwGn0qeS9feYfp+gpMjgRRaANou57
eWvWl6LJvWDvinOQd7fnyalrUrpWiL+LWR+xxIhEdWA8EhDetVUzPfBcvuy9ogRi
qP0v4CGew6Jqh23BolV43QHBcB4YlteTv/EdY09WYD1M4g9C/w951fIJu2987YCi
Zv5BIZmVGSuxCSYubw2ARevL9vr5aD6Hs9GEREiL4t5n9pFKlkqUNRv0WeoobOWZ
Ff+Q8djghjlb2pOsCphgVKVnu8LsI6F4chfIluM0FLO8wtCMYRMnEiYK3uYai8rO
AoHURSkWO2+1FKl/oHkq9Gvx7DaTT6TIGqU2GVljMeuajyfQ7GqDUvv1oIceITTj
U/o6+XrgiJ7ZM2QXGKMxms5s3vpb5fDLZaXK6CqxzJ7QDM6qReOpII6Vt+BkjhWj
cPtFuOFjokuihqPL7FRlLvVfo7C9o73yUnDtwvHWgf2ndETBduzbOhAmulFHEFwY
+QQSWwN65cOqDgKTeyC3Bl2sEd5RDsmkzTlfK0t8VniOqcph5FeIaS+T2W1vTp6V
fubKf6JcK5NQGiqfRy7eWv42CUemgUDvqREsij/qqxSZpVNRSmk9fTZd3tRjpb7f
lXAqbuyc6VnSy/NJqHZE/L8OwE/lp6iZNQ5dZB5NZPNuF2TscOX1fOGpde8aTJeZ
CV0DeX8zs3MBo7B1u1v0KRkctm9JDVWiNKgQpGn3BzTDQzoNSWvwuhExw+80w2md
MqZqoJUSU9yAxlaO8vF1ZeQvqC7fkWFqKParVs5xeGqsmtNKQmz/Jomk0gwsihrw
Ttl6VOiKf9dY0jfzijXpkW7yanehSFmfTttq1Eg0yWhRQb8DjlOZLqCbQCLhke/x
m9FIWR5n7A/PdXTa2w3B3AM+eMGTsyQMwS0mWSqnsME9GCiRIBLsQ3kVrohsp98J
PhS8cwhsEmJ5F7NvU5CG6ODsrtvJXzLFip3xCCq5CF7sIe82MS4YvW2UzwqSxAJT
kKsw4BBWJUvJsWCPMJ1WvzBBukXvNMHsPPQjw2G3xErt+2JfcnlswdOAPqOq03XD
ebmk++e8/M4S/7dwp9xDQjlQJAaOGsAtOXisOG3EUwf9YSv0YRSygd1a0gKYtFzy
ri2tsSyS/Z4iPH//GfrW7j5JNs7HCi6hqPfTXdcPVHz/XeEyXu3BLNNrr+v4n9mn
GITjgWjeZXM5sD/++6HyycH3wqIZkrSNePsJ0goprOMOLLrFHtNFzRccySN+Fr3g
Wq0sM6JXZFh37Bm+awiC+jIYvUKwHMNaWmGnTjYSqPbuZjvDnW/9gF0IqFUviZ9K
xYoJuOPJc6qEMC0pMsAsJ7NAu1ojcNesZTjCndvBvGUiiTkQvo8oERp8nZCGhKh4
N3TW8zpNTWJVcnBDNf60b3FzB54Czti0NyiezUNpp0iN5HN+TQSKFMwJg0IzJhXh
YpEfouBrc+JG3AlX7x5H5Ho6U1v4kfG8V2YB7JTtCPDrAUmMf2hHrhmk2voMcaDk
jEC5eB/5NMzPedueGx0/HjXVsKSdMjHnlcY54B93egP0irYdW8rzRe06f94LTwi8
s7S/v3icDPhSqm5OC0mTvOdmOE8unYklaBYx6EIKKpqhNTy7aD+81H39jgtbLuV0
9mo1fDz/2AtoPYV/uMnj3yd/HMA23FV9iENAsxwsyZ02oWLSOovabb1kQcpiZb1v
JuQmNT93alP+ntFJAA9d5wsBkNbbcbryPUpn39eG5ehITuHGFQvCzzWawEeojter
ynB43LTNLKg+BTuCjqhMnMm2t7k7JUgOFZXYIEGtRQyvsJTmK0iTlcvq/2+YBL+j
1KCY/HnqUb3Feu/xbZZkeVUPaf1al6FijH6h83qjxj5SVzWXu4zjLB1IRQFE7zek
CjNRxbxqj9eMOaD8fSTyVxBtiO4zlGjKQ4Bq2Pv8VYYwSgRpOvZIuNm3rpSr1tbp
C4AW3gv/zMXBO9wktBxLCB/h79pQJpUhbpgPL7BAKKpHqySmJv999RDVA7BEvZKJ
tXBzZc9u1RA6eZ57idnwolATO91FD2s7PfGJmPzt4GWczAuVCWXnVBpOXqmQr9Hp
Zdixqijp36UVZ/OEEl3ObWkVgtGvcbBkrXXn/9bFvvv+nUyYyagSqEUDXZAwxKzg
0OzqWNJpZ7EUXgflvR1cm/8TdcwqOMUz3UA3fK7wYlum/Cp2yZAanNFuHmiZpM/Y
jgV2AJonwlm4sYsOhRmaDCzIuNdC8Rx2Qi4WofnNTA49O9UTiPyA0uO+hBVYpG61
X+/x444bfpPOr1iRhq8mvxRqafv+KIqkyW2oLFmDp9nDiorCoU7gNTqYglge3kHP
lvW4VqVOxUiiYLL4dhIi/iyanbVOplNM/6yAiPw4zoJBUtVIPHjp3ZUfIQkX6CvP
VJCiEfJz2KUWHvLjx3zT7YhfVLwvhbe44EsP8Lcf0w1OwqCR8qMc03D5PGsMade4
CuBf2DxP0dbqsO2001eIJF03Lq5iQ8U6OW3H/fZFZ+U14wLJYF81BxUDsVbT0oZj
x7uVcQiEPSnF6u/EO7UhoAci/iZFQkiEey9RBmihKLOLCWJr/c1Kj4tnrbI2JGF8
SLcrYd+a0fjXuQhfqTeytr136CRdvYuTN1ly9/kW8kIEccpzuorBct+FdORx9Fga
ZZXo7WO1p/XxfM7uPv0AgowKewXJpz86umXS9j6QS4YjQpU8J96POnyAdDUEpuxK
bIP7DuXgymkN5pLSdr/ZnBb5CFUbUGrfYeU6HcS1aFXwyODs8eYfYWdx+llviMVZ
P7lb4tm9f83Ha1VT1WVC4Ku1ZZfTRtJIPiKWbs8EsvspOrU7gmnBs/PnhlA4NAok
NBk8DIdHuoVwaoSP3SPoc0vmM2VojlyrYPCc5L48xcTjNXSmPfcLqWVpjxspTD5v
tYnmlLx46Itwo8k0TvZP9FhMcbe1a6fuCDXcM3BeQ7pkGE6dW6OqIyHP6kZsEJEd
zTKD/l2uAvJ1Gt+CMye2e+MRQf3O5c4hGRQCfu3B6a2NGjr+vP3OfMAknFEIdq3T
pYZfVRznnyreVroOyQ7vOtoN8k8B8MIE1gQibZdGxIbC+lnvNtyqks2rw/lKGRD+
5MG6UO3cmt97GYJihMXt3vjR2ZKSal4HS+r0bew61pFbvBIUyucxrjtphI+8mTDk
29DgLcK6zxm3W/R4CrckL/SUrsdULPIk/HUd52eDblbSpmYWo4vgZ4WD3/DN7PPx
+3QPNOt58qxxDuvBs0vmGMyY1sLQMkJzSdOsKYdtZYkKp+U/cidb0TVZGtJnzHqc
9lhWQAJTvA61xvBjCczyghaWuWnHCC4K4B14aMmM7HGg1zCauWFR+j7FjBrjmBB1
LZ5nHiO/jDNHGF1EYKuW1BL1vIy0beWRX5n2rE56y8Ii3YBeGwnNMhmBFDhv98on
QBpnF6RowDEFe1HZPjA0maBvsYUv6WqUvxWf8U9x8VFWTXJ/u021leGQPqZjN64W
q0nRSLl21r+JQQ6/Lv10orjvbQv2NoKDxQNylcAW7orVi6GnxzIWwti0rbjPFm8f
Hriu7b/yBlqimmBGviVssQeJ+iu9b1OPu9gxUEzkm/kwozbfyMoIxmBuMQVyHXDv
AwNKFrKJfdPXpcNS0+gbHueuXHKRQptYwm0+HmNsyr6+pj+WPW6i6s3Zj0ALU/LT
PGFuHE0TMuMz647hJyGyLYA1v6V6+RfRNmnQ8ZTdl0jekxaLBisUhD2dB19evwee
kI+uRsuYeBxrbdlbU1rDhXjRJfHArOh6jsLswU7wPnUm2omrBvsRkNtgMEK/T5K2
u8IHm+bBt3mXuCXrGM5LMQ/4EnLFw1VNC1Z7Is8uN7791CMDtr8wMQCN8jnFelTq
ZDLG7UsY4mT3v0Hred3spU/Tf4d9Ri9YIelDuE1QYGAPgOIm4OQ52lI9/UBwedAL
10PP4ZPyrPyvB6yzmQ5jxx90wLmxlFJ0bw4Tfz2porQcGYIYNrhEI1cXadTPyJ9R
V7wW+CDa9d7tzJF+AvdX9vpCSTVxNqicRq0HJkzliCUIPWzJB40AZqOJhMHbyY+U
/pn/XWaY0rfvqZUYz233ULmgj1xhiwicWJedpzT5YMLsYYUvKy1CTkVWLEG1zweS
9lnYuo1bLICT5xowtL3K1dOtVuFU3b8PaY6BMmL/p9MqO/ZWToyvR+3fHSq+1zpw
GSzt3vafEv5gLRiPWgZ/dubC3xFhrWCpAg1kxHJ1lFFwPL6mAOIQX2iqN/SPlW45
pukpk55V9uFSp7UAaHgLS/jLU7DBE3QEojmvsncU2/l9LRqaIV/ugLZv6hHjPB72
h1xCfmcmIoCn/fEnvvdjcWWmzmahnFuFgW2y8hH9PHKlQ1EX27A0HtNRrCGvUaEF
aNablPtSf+3cu3Xz+CSBQ1tG/jBx7W2oaL9L9H50JUk8ODdQlLkU9XAu7ruSPZbk
zRNI4qy5n3J2lp3J5xdDyqqi/B5ooJRy6+2UI6C9e/cx3sm6Td+MhQeGjUS0aHzx
/FTtVsX+e7LcPo1qLIDEOOryQH8KkHYyAfNCDuuBhWEYyW2PfUsgC7kzgdlzfCsu
8LEd7/SxB5FCFQALG0kf4Hbhk1g9cLH0WAtuZju0b/h9RWFP1OVkDeHmT08/l9eI
GXs7DAo6yLk4bwAT5ovGxljmqROJrZqx6Sv3oQPqvArqDIhzAzFyxhb5Ehn40B/j
fc7xRjKLOV0ufkuayB/w4QAIN6AiH7RgknFnvFrY8G3W/hz8MrbjGeE0HodgS/1q
ym7vsdx7Q3JXAHNl51NOSIG47AGs42NsvXoKe4yNUyBMclMY+PgOnYmU1766kpBD
7jKMDLTxsQOdwduobPboO84SyzSdCPcvx2lCWf+hJ6CxRGcxKfE+OP94vnNhUgKB
kH4czv7yhrjrJCUqMNp8MdtchU+wYt9wASoc4TNRh6dkuX/u/QMIEdjEFez4ivMG
VaVoMqJGGVpcY4J678ele/GBhVdWvn/yFhNcL9rxXqOx5QQbUVBqitCIU7T3hnRe
CW9HdGYjDlYLAHMoK8eK4icx3R7ZW9kcwF1g4y/FnvZ1bBfII1ru+rfxDaqJ+OuK
ErbZZMERJGT+3NZuYssdXf+veYRJFN0KTBggq/tIE+qJBbW+fCZsKmzgRHBGM2id
ii4TryWGRQK/3JPedvjvshJ/qAPPU/SLxwv7DHBhv9pcFFw60haqfLH02Hv/XKkG
Dzi5Nwhv4t6XvE+yVvMdvzBptkYfGQEyM/SKhp0IHvyzHQvVZo4Hck1EWnClyAqg
0vC34FefdGvK4Uko5oQu76315/I70AmLSG/EEPmBnon4QgxyDO04r3eXqi0naHeu
bJaRsFXyqCnkXp5Xy3qKv7pLWjl49/1HFs2w/Qu709YFdfIJjj7hHcENUbkabdeM
JUM8XlJBf6uZNBgoto50DDh0Q4i+sHj2aTHhWEwDg/OqNjEvPoAHYAtiUrfiBxI4
k+xCRYdg4G6isGRjVJV7409pnmVJkVCAB8xxJoXksQlwpMMZTXp6qDFm1uCcldjw
3INBdlRBrc/corY9mLJQDQo9uu8ihVivjFH1EqRb/OQyqeJ3w4x7UhoPHNCfjpq5
UbWt1LdzWl9ud7eOhz34EceqdOEhRNjKKPFb9UyxhGQl6QsEqbNgTyz4jCWNLaN7
bVqguTNmYxyfa/oHFpRhCzOU9ms/dsdH9NTddidGZAyxpbtp0wG3/srm9u408gUf
F3JEw0Dm/T1Lx9s/GkJNGqhL8KiJIH3nC40pU6SJP6Ia/iCWiwE8GiDswM5seWy+
7kZ+zy6RtOIZCPeq8MXFYDjcPyBppdJcRjMkjB34+vrs/VDBxih0NNrJ8TC4CZ39
6caxNSrxyKP36hIz1L5sq2SWdoT3XdcKAyxh4gDDfJ3XZVjJSQFpmRomyf4NllLc
IFvDh93q01L5en8SzO/TISFHZBrjraqndOCR9yRW5h2uwdqqiiAlXCgJDxz6Bw6P
ZdAhuoX9bpL0TEpm3ybrmcvEBSnZ89TIutPhRpXAtDOAZErS8nt29H4Gt5kszvC9
EOxbSkoOmq37RgVyERcR7t1rrtOYpG0c30iEdvJyAhDfGe+KdJQsKJv9fj5RaZ/q
DbeaV9x72lCIqlTkgkOxNP1uy4aYlnPiEardxssCNlHMlV25q7xfKEkduURlmYTh
UrgAMMLrVyFUcWCnwvo4xgTiDb5qRx1F09KVRc/OKebyfZcsG9ybcnqr7Mm+F6fC
LWsr7ifTGSzt5EyModisXf5IbuxfKgR+a/FgyDQugkLBQIWvN2ZLXnxw9LpBusS9
7qz4HbyWj8o28VpcuqmBITwNn/e6hycgiMh9Gwv+37dwu8uIJUFi5Y7RcOUnVsyQ
J0k9O9LufPNNJeXeC6oZkKGtXvCGLF6c6EWGUJy0xVI2xHfRxCEitYSD89RWAt3k
jf5sZvwBVeCGXLO3659cpdPY4OfLRbYaMijB+ilBilFAf2hEV46DWotTJb8J0sEo
NsCoECwJ8k2AwQp1uQyktO9g2T8mLCtwRGOZBk9/seiyeZ5AHjD0xhGKwkJsOoMZ
b1eeaVLokG66ISW43QN5mFQ76bE/AksTg8vgwftQH8KB4x2aJXBM9Zj/4GI8RTtG
p+oax0SS27xRhxIzGZgc0VrryQ84yZbdb8nztZZgUSBy35KS1udmbmdNGujV8wVQ
yUBd9q29bh/woDL8cyiH1p5dQiHXx9gFSyI7IrlOxVWfoubS7lHZvcYfrdWfFS5t
AjK55T5q7R4kMxRGZfaDZimMMh6m0oXwoWPjQNIuZCiWc5Bp/albXoeaumlJOMFe
kcYpwIJJy01zjmFz24Zu0V8Bw5iOVBYKrKq0LSQ0aemLrZ3xHNRlMnR3HmpBnhpm
KS9LimPOKnQOQFUsnH8JGBxmB84ox/YfhOJf2PC9NBEj+MdRwAMVibLzXe8jbokA
MfQf0RAS7xPnz+8SILxAdhCLE+0UICuSU74XH854/6F7lZurpHUykQSu9si1ZjEj
hQGtMxf6e/Uw312FLkCof+y8ICVOqGQlbZkRkX8gFDna0yWChn1IowvgSLaPcfNv
CFTv/+fBpV9Z9BDkZulSumlyX9rWMjBDMVH3XU5tf8tkWzuusvbTtLvvpzXaz9+p
S0L4627Kb6ZX28i0QMmDRN+veF199ou1wjYhO0ylF53IlDDi25V/Dm94HBifAXBD
Lzt9/fndjD6jx7Wde6yKDWABcwHYCJev5I5YIjjYIO5WbAnk6oeSW5wHARuIwTmo
aQQi2TeCFpUaRSaUA7ciQnsTCVcCBp+OPxAqHPuYGLxqmSL0TSYzXOFXB33wKLzN
rzRUlC1YGhfa/q9PW9b+F35mWvwYzE2Z51d8N4kPaUY/LwAUb6xf3HgwqCwpcBvD
1fv7pLTfPUiavQCbEzIIoKWuLEwo+PmQQmyALDlfTKXvYAF4znVqVfx7TxhadtPX
jvpdKKWG0RxswItKiOElpr4PRGEQ/5ef20NSJmRp27YT6ZEKvKdHt8O8MgTMdm29
HWARQYkmx44HHSHLw+HnA+1R4Ua7saC31CzuQwyi7lKd7qA+mKOahzygxXk5WfFW
DHVshS31AvJvFOSAqjABNsA90cT3bozV+G1PjvXSlZRaBHHQRNgTX8d0rZdXCSfm
JJatNZv/iY+K13tXDtzRbzYZFjr4Nxb/cL3DgfGgfVfhFv8O8KlxVcDVtaNONEix
CLk4Iln2CvsTDHZ9Wf9NQQd2LZCAVylwj5J2OsjqRvM9yz1UDjtawBfgWxX9HRTB
f+79CGok01azPRYIxn5mWXH8RDpUC1T95eEnfycqTugNWMwKiQXa4E9K+GHhyYWb
1fboSAOZA4C5Fym9r8eRmbAqQqx3u4Hon9S8ce9IXKOUULapZQsBfCZefkKREmEX
uUQQZA33X1ebEEvMLH376ewdL2GbaTMBcyVsPPF7R5PDysW80MMr0yVGUzRszWp/
F0AUlr+6Buwv3k2xUkaOYUsLY/Sd26BdNT4UHxm4GTjLya6xZMJ3BIdPNOlkLguu
oUMDKDbqnZ8s6tX7eQsawY2+zbKAmdvfXEHeBEhRdeXM6vSgerBLtVbRELS4kxH+
xr2N+mhewNgbRAjwFo74FT+NSZ+rotFGbFzYofEyC5Y/mKYnrJKsaxC0POaKemeR
KScMD3kYZwOF/oXQXWT40TgoU0feZLBl6nowSWP668k2xiuFDLZW3e4z52UmIlX1
DgVFsSuEX/T5Lv428qPP7LhoXiHzj6hPocZVkalbCk7sB7RACeCFw4pY1ObCO1wo
Es6iHBwVcPV/Qt8NoxWPt5ZqMzjr4WmKmIgdB+/LCI81DTWn2fCtBCTdNr1QATtS
L1oEU0TxNTADAC4R03xqwA2P3bFg8C5C4BENAzWnRZBbhIUHHEe3IzkCyKAtxUAO
6ham8H3LgeoC+/2g7BOA/pCtifIriJCCxl9UmSmxPvQwgIzb915JkUYIbBzjRe62
81TZnGrIO59ZNmZZx1sgUWh71t5lraS/Cz7QFEvGPdZ3bxCZHbTMXHb55NzPQs+1
RondFaJ14gkCeKREvjc0yPWlcPpBjGMXxUkMA2SO0y8tLGFwGhIAG56ZrLQSHuYz
oNuU6UiYgwkuFDaySKf9Sq44ZKFWbjByLXKViXpII+pexl+K9VTpGmsyTvCWNnOl
mEuDPMtQKAGxvEdbr2SSgdRf2jQlUbGh2Q1yXadj6bWpcVx4wXkXrKqTm8bMWNDp
4SxSUbRZEmJsHW5O0fplW0cpVerPlaKsTLUtOJSIPMckL01SzS7uXAk60I/RbzRs
jKpmw0+6SEtkQwvEAE2Q0nZstJrUKYwtJ641tojvXbmlcdNgjeaUCkMCNGJ3loDs
0B0e426P7cJJ1jIMQNMfXrW/7xIxDSsZP9qKqZBYhFd+ThKan8aL5jBWI73TwL0S
Q1PBD+tMK3geFzoezD1DmfOioO9BtSNGR1yun/3W0iFa5VyluVdtyyHuFXHiEyQf
5sSc7fyw+kDF1B9W7FL2QKs2Asf1ZnQq8o1six49k6es3t7bUbRxWq42GRyzIHXA
n4S2EO+C1ezdg4m0tEpUjv9/L/L+CLofsH/TR4bc1Iv4BO4cn0Ecrc15IJCKhH0t
ssK0/2BgvpdS92dxJHlJbmDsOnI359gIw7KNAf6Gh2Ze3MfMHBzBwrHXsvrSWWSj
BhsNHoYYwA4NYbADusiTNov0TM9k3h54ej1IDUdRxyOwNUNEgMglsj1tAGglU7c1
QhLcA2IJ5N+upmniRP7+kM5ks1YqsJ/tdTit0haclOYSbWZN9tUv+ufV92ICUAax
iuI39I/jKVENK/vvpmlUltApxhul+bzVB0nEhiXj/jOS1H4SU/kxX/pEsNmVdy95
fk7lVLHDWAmdVKhcqFp784vzVlubiYtWR8JtDrNmWOTrPcBfrqb6hOoHiYaAwqTp
rdMX0ObE08iZbVoBOA/RDgWfokcgFMQKhoWo+Qeh3A7h9SFfEsSiNnYO6HGfl/qK
XljlkgdRCemcFOIxhcT1YcKziQ+n8grdqAQvvIVL5ogBQco0O7FDIwoL+O64Jv9m
96Y+BgUHvQvl8OQKWKyZdXbPSKW/mKtImc9DaQrglVjUKme7bwf5zgJppClPzaLY
+Cvj99CCbVhC9PNz+ZUiZzpx5DhxrihM5EpyKtbUzVhm0vI0vnXdLtF/Lwu25on7
aLlOmK1jG68O+92HAOTSvIe8LuyfcKJuddgBNYkGPtefxQ1MZMlrn6yMw060yOGf
nMZyqo87cRGueK50xmizIQDgPF4fBCzMXwbFOyYyvX/Lx4/cfBvpE8rBVa7gpvLA
QM/VRKiScU5z+uv0lPvFEuJhOVFhMoT+pF8+R6Cz29a9dd2EIrqNE77oYnyfIwav
7YXWL4DTHxip4rWHYKpekf946nn/FOfxUx/U6nHa2aHfG9f98ytcUVUZoqYhgNBv
D1KhOfoKc3pV/Dtxt68xAFutZ3Ow+tsP3as2LcBacXA3F9PYtynzNqFl4amI3t4Z
K/y6sBd1cJRVKHjPhDIOKGz0/WPyjUgUUMMm4adJ+mFSYgTkQKn4PfzXObkhXvl1
YD38H/+iZNSEw7JGekQ5KKLOOLoc42sotat8tx6zwPw7uZzJgSdQyqeFHTQh0aDH
Ee2TKCuTMa00G6C9KY0TPmsZQ80Xf8e2iZPUf/NvKXvcE9CC3obeciReTza5MdVP
1CX45lsaNsrADZ2wNQggjfiYA019ko6BDSfo8XC8Mbutfe9oKs4xJ6KFxfjwKG8K
yg2HkRAOsjQiHoBZxA9X0w52+7Op0dyFlhqLLYJNTHLle1/AMdDlyao/cdHMHMii
/U62EgDaNf1fmQE1vwySaQ6p5IMl2e9GXG56BCKwGi+HdzotOFZO8bCEj3dPosRO
+ybOo2FL+NbvWIsj6rIUFSHdsef24Y9cI7oNg0iYK9uYM/jhRbtgODdcREbK/1K4
45zY7Tv5DCiiTce4hXcm+2E9+GYa1GIf0/ziLVDgdyOE1wih1I/tgVekjDzZoziC
jS0m41EUnp4trfk8hqfuKG3lOJF/yb3NJS1aSl85QlbqoiZnrrXhHcITfr4VGCwB
+FjOwWlTwQjK638xbpmmxgX4MU58z7EP6eh8zqupWVkljcbxsvNrFpwKZHe6MSf/
QoYXd80rKveBcIwLAqr5pg7RDMt3IRWLL+mRJswlwxPVeWJPL1RAkvWntwaRCwVZ
zkpasRw6+HlYrD20aMOB20qSPGlNx1u28YzxXJP8t2hCCSIH7b3VAi6eB7dX4/Gv
QyuiPOdUtA9/hddsGML0rFR2/8ynN2/cIxt657yNR9DRNb8trr+ebYxCGCHgoTKt
i7kQxK+54KJ+LdAuytDVj/MIlqrd0ud9QHZkb9ERWtceaoJ3t+S0oZ3HSEYafijO
EqGl9hNahOfqxlec8RREIqg7NTm8yi0QWZJR3b8Uet6eaAEfPqBvhm3jQatb1Y72
Lp1kHW/bRRwuhFpo8MAsQi/58Hn5J1xXOaGGUAY23f/nqGes9/HVuv0Et6OUuHsJ
SVuojTrpuGJTQLd+iAI1AzNSSt5Cj8HHs3bv6kiyhuc+ERUW/FQurR8L/mHWqZ8A
vxRRl4tWc2cWe0fDEmy/9Lh1C9AgV8zalwrXUOxptDOy9k17pu/6UgMJ4ZY30MGP
pPk0caEraWFxF5AHbOQsYiIVUfCRbIkJk5ClTSozkJhsCcGWPzo/rxtNMf2gyNbx
Nh6PHUFg9bIZxM5TAwgQun7rUmkR7xCCSt6vg1Zp89JmA+uRWtTukl2tgRFixtCv
yljoU4oPDoVnEhNNHUxKg18Wlfl+m55cajYn1DI4GF9RecgCvvhEwxTJIuh3OHV8
6OS0IaJmqGpZGhqUaonoY8aldEsBU20B5QQaO8T5sAMBhc8RuMVYBhqPVVtlHwo2
VwI26ciAcr0wwtx9OTSrl3fLupPZt6238ozUYXSeNIV0FWsvi2XtflNgARtMfXa3
hiQOPkfhU/6nZ7+9JfaC8I/YkpyX0mvM/SZdDGkS1NLDeR8YrHtnjzpdhQaZ4bsK
sYIWdv2cPQGGuxzDh86fuCbcDi8maBd4ioHykvBwyDPCyo/rNSnnnwEClQpRDlPZ
slgAlvDcn+gyHtCeeB5c6gUlnw+XVcvvCMhIv3juDO8x3GtOUYkzo4T1E+FZvoPD
eadV6XsQCCh/jlnjXMonyvPgu3nKg3x+UlSsCVOvxYB0JS31CFljlDEaL6SNLbx2
V5U6j7y4/+hHICZM1pzdJty4e8ZWl3Vt1GFdbQgSDBQZyjv+Xh1m0JC0zDZJ7hT9
3iAO2sneXtHwkeOgkFY1LORSGEx0+kU0jFy2G6jCdwGBH6aq0sL/gMgNAJK1UAHK
Yat6SU/9B08Vr1yh7dn3k1/eoDlMKIbfA/n5tS5sl2lXteC7x5jZTDgJFOpJ5RTs
mmo5SOmgLrTiLQGZGEb/4E8XrF1CbtV3BLTM9jMW5nnQT+dk6S7owXjXw+DEgxpR
mK4UgXGYa27xAXtUNmkpuVCvFUNZ4v8ZstM8UcL1PT2k9qBs2Bieb4ReYj+HmUvP
13QrNhGT+/LQ2dyhimmQ8iqwyFGTl4hps3Cu7jixuueopOiCYyesFnT8l9r0wK2x
UeqKzildKcoZo3DUkFFiNn12HM6jWh7ybSTnz2U66VvSN9vyY1B5OqHtAf+x7Nb5
3NqweZIBPLvQOjo5Xcd5VTouSZBd7ZeYaBeUizyfaMkgDgWdZgh0WgqqO0qYgcoa
C62RPdRBtbVhc7S/og7vBxdcSlHe824LtNAyNLvrO15wmDPpkxPE2EkeiANg5Jqc
dPUI4hNuFH8li+Ij0jsNNxUHj6Owk3HG7DHUHcVr/HB6IuEeEDDvCFO0H99G5RNQ
2VqaA3oiFWqENTcYIK9kCvsqeAKeLqOHXpwAdXaNqTC1X09R6EK5rOYDgAL5qcSI
yO+LJfoIJrTW9aJyCCLGgFdpjC7DoxCmkzynJbvyOywxrWvjBgisOTfqL+KibVp5
m8G6LerRylEJjfiGYPg3TUzTY5xFNsl01lTwsUWIOxW9MU+vxM+wqgBso5l15JrQ
v/EGgjq8CP4PQEN1p6LIFNs2J0BP6daLLtrCmXpEdbXClUmDRlRukMB2HRgR7n5x
SpumKWTiZRCr99oPse+PxEckRtqmdHOIAxyFm3GkSHur0rV85BwidruMA7OkXu0s
h8/k1NrdAaffqrlkIBLAJJQdeBTONimJ/8KsOwBTeoubYmJGcmgZR//GizRftvbD
lS8mQsk2pxrieUBnZShNcyhf8Hu8seQonHj5FrUb5wiumJR0ZAcqhtrWj9/aiOT1
YP6VkUs4YIrgYDqtY3zgHitvZQgu1jVDcqz04aB47w/F8U6CwxKv59AQoTeptb+V
j7el5qzfaKuEbyFIsKsxGAza4uVrJ+YXNUMxu1tGtksE+vX4Jjz1+q1+3anEKVKR
qkSpBDX80mmxZEC/3qep4AwszW8E3s7IyBYVqbC41vhIvpGOcJUoAa6Ww7BFS7MT
EB+DCbnhxZRc3Wdnrv2SoSpZdvYhErm9XJh7jLWAuRuKQCsK+AU0b5swtLwQKTEn
C2Y7M1sQXUJuDGX5kVu4GxfzUutaXQ4HnpctziN9g7TQ8PUiGTkrKwb4BrY+KpU9
LxKJaeHktMaYpOhyklEQlP0bZRY9Ojs+hCFEUPtNZ0UZv60xdpDRlbip6Bc0xYa7
pUdeaEcM/2W4nvzyEgxzXC5ET392tKnAmWRcOViydgG8uRVS44pUPNcC6TsfX0sn
1TTSmFPr7g0MTzNc8qNmjaC51iSss+OyZgYAv9KZiiehHvR1+MxPotWLbAw9ZdQk
VC3Xe2zRHcog1QVcKEyhO3nk0K9aDa/kK5sjgduSpDNaCOSBX1CLs6YzTRSqIOCa
fD4SkMfSWi5qyXhv+q69k0+iyRivevaDf4nWjEgeIHVQYSqhUXvP2PmRIrf9BPDt
IlLjjhTJp2csfbCV5r12snmNM2H5Y6Q/3H9kBciF+rhke2JqBo0WVFWCHqiMq1nj
a+MAYBvR8meY4b2XxSqGwbFzdx4Ob4QpGfxfLBK0bXOI2SAMn4Ug7iOHFhmCp4tL
u+EQZ8d3bOmqEVRQWa9e9Tpn7GkFBsCGtGWF4+60ram/vniZdNKoSIu9DCKJdOHk
eBrWDemwUlJh8rAY54NUq6jgRhZza8fKQrUDYH2AEzYXjr9MN//AeUwZD/iQSoGf
GOmndt6K32NzyDrHQ2AN/iASFx3wtzgJSB+7l0Bcseu1ZahYqMAE1tAqxiq3LeqQ
tze9Nmjn+mLpQ1cme+wyBEdyHle34ru0GKfmmsmDzgoUXRK4UnfnUkJwHEula2EL
hnYkKlTNOsQsI6gezMtPdQqc/XUAFVfg2EbpRx5aKILYV+tNcPNprFDh74pfNQXG
b1vvCN/oY1HU1WG5nLUVfNsEZRrP5a9qA2sLm92yDz9PwdGfePBcRgH2cYspRQuR
OJkwkJzV7qSskdTBIgOoX2mZLYHPyk0Bk1T+bGvH/eQVKdh6HBiCxfa050zUbcL8
M8sYctjyn8Z464RFO3HFZ9GWE55ZKunRojD8yOEhMOfdgLBMNQagialoIPGxkhXZ
7j/J7ivKa8I3/LOC8Ha2rRNAjx2/ux90Z/om87PumH4RkLsXWPFCR7jaUKTwjlQw
KWyXuIzrHfH7mVSR6R5Ql1WPWL8sFnVWLZqZrjwhhB3/lvq3SgYskaPJY1eRWqij
/kosRgw+gNG3vUKjWywhLP4NF5dQIwsyLqmS3uwcuHsv+uBhe7fkIIO5Zww++6ZO
tN5KJz13LZCeshZ6NnFfi97jx/Xqeha8QEDeRg4nWo64oD4CqOAOyL0BTsqyWCLP
7WUI+m8mQY05aP2EjeAdXHgJ2Sibl5tebdi6QjZ+dZtTD46VNcd0h/fFug2xoMKN
b2nad9mXt4AjtS4NpG4DiTxStsC6jpwMYCUOcFF6sCRAIN3CONqCLOQv08afEuDK
Ef5TJxFrhFZxD2U9gVZ8ZurwfO0joGRkeQrbUMP/06+q1BttlZqp4jIbJQpYZxuF
V4mR1cs4pYcZ3teeJbjbTI168j/gEXaJLpfHegL0koHU4O2/C9Cwkm7vilP9phKZ
WP5iw4Xih3ftvciPwAkxRebasLWaN1/mUrhETjtkJ8I/oZAC1x4cdi3/sUY/qsJo
Y5TXU4n97xW7fo725lXgFhTxPnHV3sC3Bkg5A7qJepgO/uPs9nI+Xey2XFc+YGcl
O76RLph46kTw2eDQGqmoEqiVF2AXYezqa5M06uvuMqw7xglCH8q6qPUMP3DIm2QY
kvmLGhBhme+JwVD269oXIsMMJBAJSyB4Xbr79sGXGl+zMTw0Vw56fqoLySvkFk0c
y9hWS877iAMMvGBKCaM6k53y2cG9itXG+aW0qQ6mxRgloPis7+ZEVxjEnVNSm585
4l1jlmGG819WaFu30WLGhHihXY/mDmYC8pZRlm7VM8SKeOpfsR1VrtmC4tHpRZBt
T4Vl5HuXmbWRUwh/LGUrcMPQ5ySUHYokGORPqIgYJrXZfGGlsPr0QL3LGjc4xhwl
qtb1h2EDP5p6HO1SW/VNMonnxex6XsstexUJSvJccRF+Hknw+EdoJ+G919oUE5sn
qSeGlYSE/M9aX5wrwF42n+3iMn4k//vqKLWtEoIQCoM/N/toZw4823VpvN0Xy8ZX
tSdlhmchQyUZI7035kUUz7bAS5HS4DLBtXiYU/5tk4qqyO4S9nd6ZKvNr6m46pyk
ukYZMUq9Yu02rJhuyPbB06wW1FLjJXLpafkTK376shE8eomxYNsaUmGnUOVG0FUA
ghRYPN3s23L10EG3aOAUZ30Wt1U7a6u6QDWqOw5qSuS0bBcmWb0YzWuoR3m8b61H
QvaMfxe/44vMf7kl3UYSU6TgkD6yZKxpD9iahRSCAq/S0ccjlwnf2w9Z6qUV1f4u
RW3xI1dbehrcsDUBrdadX1LvICoactnTOPPtqYvsYDm0KovDwZ66e6E1PRnMZF7M
3MzjiP4Knuk9aXoNcJKNVezUyslftdt5EGgUJEg7y3bE56SOTGBDLWWu3jn3bp/e
HcX8om8zXn3TWUz8ulDUVO3Qfj5FByHL726jzAJUW7vsJaGqoijehf5O3MfRRkXg
UiDvOJr5R1nrKH0kdhowa6LvszWNSJgEPZer1eKNORxQZevkiUWpRJd66GmAFUEI
9ghkwkMreGwI7p4ZSv5YNDWBbAVI5Sy0tGR6gb9AY9OjDQ7SIztM1IiFZEeIO0OU
85p49ZC+gdDokSZ3KdPT/dfF19gE3pLbVxISS0DEP3FeunzMUiE4i8Nc3+PsyvHv
4NMkthXDh1YBEzYikfDAVzVzj3aPteNmv4cH6eE+YiAA9zaQx+FyoLU1I1zLrjPZ
9qjh3JFw1KlCehLvJAyMZjGl2tfu6WC1HNTvEKpOFofb4/tqWPp1Xg8Sugrcfljy
q8J/4Ig+kqHMhuVSuocvfhQnSEhNQroBJZmCHchdy9ino4WpUuJXejXjeXPZy24Y
m6YEnbYJ3deKAPSjDjZqOuuSLR8xvMTv8GU9wvx85rwHm+T7DqmDYgU1PcxHD2gF
IJ1pshyQujpScOhb8bU+MDIMojxlTpQO3TcNMEymdrMEccgwt0xEFLczMsKHVTWA
GeEmnVSQtQ1/wTw46h0flo5pdCPzaMGxrIm+RBV9VHgqIu2Tl8SHL5C1PvtWtXjU
HiFY6Kmtp5iNWTNpu98IUEa6zCtPRGK5z34+s/VSmzmIgwyt3iRFd6a9QKtrwozx
GrUnSDAgizuEfx/hRLorVCN3+nNUrKv8Le0SE7mSLCMoMIhLiU/+1zUfe47+eXyh
JoB3e8mPU3c8DKXVqsltXDpYRPrcAkPCkvRjQjTgR9cn3+DSp8eJjipvtdorS5XX
GeZvfl8yEV+IdkwtWFxHGva8OFIhWeRYncu9eB7JAoroSd5/4OuQhZS0LyO3O1/d
HeQ5y8IpnscVPx7HtRePwEWZkPaYoikf+Ff29gXzNSZVsCQLYEQxtPNfW01F1OLI
Jm5bUPWO09PXRQ1M+d8bk7jV6bhalffZlzytLqbu/1hXyjEPWstF6fwjiWrhLVxC
KwOgQgSxdBf1agtYRKFjVjthSSQkr9ObmzZlFpJ5vQ0UARRK4OhWN7iPH1TfHXUh
/8B+SOycxveAGUKkd/HSAmGX3gmyr7tSSUSburHJeehi0lZdsLKL7w2DXMBL0KEZ
N2bH58OyTMIhovoyeh6ZhLwLcR11QmgbTkDOBIg17VhUgCZDC587obV/DV95B+oI
/niu6sTSUogrsSYvaXGdB0ITY3La+5ep0VhQ4ZdGKZFWo0jUD7kjyvjQLkfwMoMe
DyoXs5SOZRr+Jos1elHUxhOwhImRq7idkl/6wgZ/bt6Ec2GlM1EuILjsxFWPNuxe
PSanjoS/HgVYT2bb7M42dc1VPXlRha1CJ4zhx4PFIghC9gjlpnEC7pSMt7CLWGhW
gVPrEQlS6+1I3+8kYojkVeZ0d3Ygc1qWBT09fj61doyMDVwZUHGSw05o3IVYf5nl
cJ+0AuqhYa8vdusddETaNPstY2Trl4xzAg6M543jt7G2q9B8K398C6o6lZKiLNaT
WiU6I9FY/90xlRhCza1IPBUIN73iV6aMrD6D0sBJ/Y9Me6ldhqSLCB22rmfUfpDx
edn8Xlos12rFxhy8rD0O99yNT3+zo24dYvkyhEZyx0y81N3Bmkp4B5vJZQT89LcN
OaJWRjMmRT+PC/DdfZFH0HKRG7vOxkJ4KwKkpXkfZFnTs08XYyhqRNFIQ0UYRzsC
+69TIbMASJ/shpXmnzVRbnYi+A+7IVfG4GjkxpJYFcmQuvVxM6yLoCXIYF3sN143
ifqodJWLOCm1hj0aKbVE6vUNqQSV/JRxirxpTBkqB9U9j5qII82IYfkeqzLk2Gve
tpeQ08USD08y71XsQpC3cBUOuZBfz8en7NF/yt4QLvKz8fkFwKlxtZAQHgKcURJV
dJYHAJfEX1TonaVG9/xvoKxprT2FlQhmHyPEdFTsMnt48XfGcH1r7Cnv39WdI6RG
YgGGjkpXKn5GHyBL9hLdVEpxFClvVDFbYKsrfJf1upBbOec2Jh014jgCi9XnbhBH
4+8CuKlTC5nnzGwOdICalcqxGGydyhFlnMbEiUFftHiiBi3rbAG6MUQD5BRW2IfC
svXm+6vUR+mJPQwXXSCvWpnWV2s8EQalSVb+3JQNxWszTGKeJsR3dyZlQ5HJQ2km
SgjvE5Kg5EgRcY4QPo2h8aSoitrDkbl0cKuP5OWnzKtUv88kpGGHea/jd4IG8ziA
T10von89BOnKa/DkivnV0HyVI++y4DCgiAc8Feg0kefFHcDuUr9FYhl2LgkpNjSG
CeT3nWwMiysDGu04ZNQsneFjAbztqAYu2E44zb+EfgOVWWHW3zEeqeSyV+F+dpsc
1dbSptYNOYj3fs/ILkp1LnGqOcG4JqE9hx3HAFX7SYq9iPokaevBH56iNKOAovUq
qJ+8gRFS/HrEZvXw8s2ldV8iJFZqTcduSaf/DEfxI8OfneHMssyhAS9mlOdwCB9y
uG4JE8coGr7P4FDJtulAoxtGuutz6p8ycRvWDUjNKjJu0i9bd9JjCHCxNSNYpT/J
5dVxRHPTqXf/M+AmTsK/leYhXYDPQGVnV2/ALwpYxyPJpQWOrbj+gLMFIzUPVX3R
wehz8IHo47AwwlfX1/0phc3ioV9WttsJMO8IPWumccY/UNSSBlx/mIynvyymJkzF
8bHd7ib1GzdinnMydKlIxOFBPJDQ0fZXwx79f7LxLSZVIEeIfsKVaJjv7QFOFMpv
rWsksH4E1CiUTcg0qZreAQfLp2DF+F+Qg3x1W2pPA2f6x3K0f+9rgiHEQljBjUoH
iwFu6CbdWHpLHO7/ocPftVxx1lzlBClLlH0e9SyusuF/CSHis8IWGyCiEiCtOrcg
AdUNfQPS462KIogoJfnqqMdigTvbXMyMC1me/tzupLFL/h8BGzhPyB+n7DMJ5a6o
zMUQhRu7rJ9PIomg8usbXeP8A9urcsO49/7NLNR/psEG7HorMuLrUqfPeooN2Px4
yKa5a6Xyj5WwEDV2PsUdCeF0VInFReCdDz8VBooECqnE3qmpLE0dJqrbQTBYenmJ
xASeJeQlfaZ8P8JB23qzkecpMTQByI6Z7rJhTBE7VKofUYiHd+WgUPNA8r/2laov
c7yDaOB52mhruiQ7qgh5Mz0TLIDP9YW8n4zKpiVveIwQzMo21F+MYPfWGTo2CrRC
NiUf50zg5urESuACcOIVux/74xwV6cEt9Jw/94lPvHZ3GovF8lTrXYD8shYfBAGi
fkOJjHdxXNPL4C68RlivROAjAgNK+XFCIIDOeY7JUlDahP8h01xQBV9/a3pjvSXY
XJBC5Ve9hcZX9AcKUUrjhFk8vjcvi+jUjSzTmcJ71OWhYAk7QDqRi+JOxBfUEBiR
sKmkh3FAk33GzcFy+b68HAtIYzjN9rfBwReTyKx2D4iiG2/chImSsB+cWjMJC38h
BzZ9muMpmcf4mPLWnp3ZPUwAn+2tycUcmVy3+o3cRfldp9s7YfzqeuYad3ewLlIl
WGsloWWLhTMARLTzRy6kc7egYsZcHSv/avOrjEtKVTHShBwCw5lnuavxgFIG/ja2
/FjYsWjD9aA2fdz6QbwP9N44Y+T4XG9Ia0K3HK3osrKqCYW0cErZpBxABsXDeXcz
nMWXFZUNJcoBd5EOsCFE28040sYKfTpFVxhfG2gtAjkS+3tGJ162Y9mYoSS3SViR
2TzZxJYuhyDDQapPfAsZW+CeeF9CpQsBquntY4MIBOYArIN6SiwsAtXJf73Wmahb
vPBkB63qtHd27u/N+5VREvJ80DJb32V+ogysKfWaAD2qu7rEw0LD/IVUkSIj5T/x
3LhAbCkg6iATaJxy28tNKSp1INgFth2tVDMSsKHqy56HHQ562/HWiFEqdVVgRpIK
+d8FAz9QFhAj7dUbRT4HWOpw6upV1lnoQHaLtyiVXcidUpWNTjVFqKNloJIjcaTV
PdlmBk9JcUQBIuNEPseMpa8HMivtvGo08KuMRKIuw9bRgv/I37OOGbRX/C4kZiJl
Eb13w6XkJO3b6EZId0CFchC/b6Q24QgUQVBhB5SQUSAWPicqPMjGYqPDT33VYYfX
rlK7++nd4G5dMnveym7heEwR0rXdodayN5XUxffoqW3pFJz5dmWe6mBAamRbNccC
hyQUu7/Ya77lV1VyoMHFp3OPyXLHqiGPPZVyZY+yoRnaCa4OpqwYPSWDmNvwREu9
uBRlaw2Qu3zPkrppp6QZHK3c0kNIhhlsLB8u6YGS/8HD4L1268vwe/7CLnNOxisa
2elFBsH88IZGIIt8nWdtGmjjU6jMncTtT4994JggWyJnQzUg4OczMpEbmHEn7odK
JfHu/L13g50hHYdLsldSF0tHMc2YjL4wVkQZZafvKm1hEa0lPQQdcKbmJ3JfC4H8
j/wVPlfviqWKMHaRYEGiqZTFKWF9EUL1oBViUgQR1yZKYYSYsB9FnhoFlZxo/Fve
vI7cV9Vqbvxi3X4FYo47T04i8gKbYrQ43+dm4O9ksQZMvkxBVH0Ud79F9x4Hukut
YpuZ3IR/y1yD3aOSSahlcFzvJEZgoMHjVlDV0d3xXlOnTlWzgoiAWlpBlbZ7vxON
8IdjHzsQCkJNVc24QfAFz4g4Xl8i7lBONJsePVD8grOD2Oeo6Ng+RZBCDGJDOpGC
BCxVfKfG+HvUL5z9McPACzHotXTo66cw9pAziTaq25qBbr2V1lMAlRD4JkS+UIzP
sr0czPiOStT/UdwD+3szNpdW/SYgc8F+cb5kHfqLOsp/o5FewHT88IDZRflcdWYq
xdYua6B70Uq7ZMcDOFTNqSIB+i0gGJUrsIjlHRgKVUqA8s1carb67Ba+r/bLJG4o
VhobjsF1qRLsnygRyeLU3ILHm0W1u4Fk8l7+LGVQUJmYnT95hjPHo+aiNPm0azba
Q5U92SaOnFW389Ry7TJE4oQ7FkZvBZpZSt8TKBQUbkrxNiaPboZxwCjVTFsipmzz
57aFfv2i+EpgsRvHILDIlm+aoqGnu7HqCsMU0w+0u+yYdGVbXjrZgpdsRwt7D62l
TVVwtKGnNG7PCOwJFpthwmyjulFu2Bz/wVJdvxxFpcR+yE8G7/cVqb95Y8UJxocq
4e5if4IF/tJ9ozpIjQe+6i9DN92ryuihvLO5B/WbfF9zWMJ5x2q9LVw91PW7zkrp
KKoxOuv1O65CTaTEYLn6ghCj4jvNnfxWoGntmllagN3bu6ERKHZkJXSCjgb4w2v/
U2GdbkkQjbTDVelMuzEt2mpz0vSLm1heiz2L54BODMZazZcXIbFY1ns2ty/AUQFc
8la5VOiwSsADIpuR/XBdAWHLEcIan+rKIScikUmyBDGK7+WGc5ohQz6nbOkvNDks
IzyxkmI3TaDuG+T+EEgFF0CbQBhYYq+oV4R/6sNOpvexY2aFm7dAM9j6CUPyIP/7
MFzASehrVFy2IVwQD/WjjAt6MmRvYl9z3F/2YdF3NccWH2pfyU7x0m1oxEDo4mFR
fUlDs35qdvgO8cIdZROhgWI64/UXszIqF4f+0DfeUgnbUGt/8nCtP7B7xs5zLYcN
2mzjYSQRqnW3vVSHsbMX0jNaICtrkey0kDbXQAZdm1cJySYQgVez22opLa5h9duJ
oNRO2Dv69jDelu5nQfLlfgcxz2M6Bco0YYkM7hycv0LV5bPNGGTqq2XEMWGhx0v3
hgSeS2CNX4R+iejL/CYs3X0oPA5yu6h2BVwI26WqUnoQo3YeR7Q228VqzA1zjo92
4pjy74E07HrQpEVLXlWlMPpmSD1gHrG9mdT8mvJmk0w5AIKnpLfxGtcIol83aVwl
rfFWn35khE3s1EnaNgRuO2V/4Tty4UsmHFEn/sk/xayvSapIGaEifeN24AVNKUPz
P7RAeJ2d6jO2SP9+0z4agE6n40QfpDIYGQb7d6ytEvmHkHsRArr1aw5XPVloJM10
flE+AxrFlpbaCroGnkG8ctQoWwzPRNTDJZRNqsWPKFa4GNlw8PyPTJ2djRg2Ztkd
vGO5o+RpvTh7qJPuT2pi2kl8mgQ2QxElG07rglyCsvosHTXXvZJ+YNfJ9S2GbaLk
TaafIzBIgz6UTSvaeWS/P64pH/LR8mM5VNv07ST4rlRTMl7TLIJYs04o7o+OjFx5
fOvLsoaP0wB5rI6PM5F04hxdPF2PMiouNFEn2PnK/YVmftE1p+z3XG5VWC6q/FnL
N+6IrSix6wCJOU1UOEWIM5BbDHTB85GUfJ+aD+5wc/zlMOV+txbVCIOh31QrRipt
5Y5nikeW5xKHPQC69pkv9byLOzhnEAG88SY/di2hhg8S9WV7/fG4Zp+uNFxkhAsE
gNsVFe5GB1Su2XcJVKegI8w210KhpB09+wwDARcd1sBDuSgcegBshoDWlJ++YVtl
ZBZDcl7C7lfPMVvcDTJc+zalkXrYB81i1I8sGaXyJXOZOzXhpyEL6O3SqWALcwev
RXPQ7RvFHuR7//BAx9Fi2keD22GZKwqkUl5s101eFGMq1qNoUmzaNOf2KjeCBBM5
7jSVw6mlWevpxXv48FoYTqRSsq7aLJpd7CQe8Y8+m9BC+tU9bFm2vgRhJ0MdBTIs
eKpFyNYhc2j/bEMYGkidleWDA348P/GUpaoxx+oWyXmoOOB1+flRAFQeDtGclHzD
PTzSupSDAO6MAtnHVtBthSGVt0be4/HsPHnpZXg/qfVnKXvpDZakmnTTrUwwoCYo
wAyxcSFodC4d+UV/eTAvstjTBAUfd6Yku3GHRhWiiqH69/TWa3MM7irBISIh1B+h
YVso2Bp1+JllCRQO8uhGosS8UMnp7RMtZVBA/aAYVtRhInA/0cXaNYqqD9W9RctC
b7zO9oxrBXPPuQuDNdQDFhJnPM4kvaSN0phAJDwE84iTtnDn0o73X2MMPQp7QH0e
BAjI5ltM6GyVGb2T1WC7aiz6oG+uD5sFuvba3Kn+jtj7IohLuoLG6hpu9pf79xFi
0zgCiILODPTFdOU+33Y/iSjG5EcPOJGkqjyEp479ryEc5fOmEYv74h6ryQkdHL6+
H1YO8GAptMttp63nl+mngp57gJz2yUDZJbNDl7FNR6ktEzZzgs5oZKETjn3L/J5x
GIxrMcy8C4svXB4cvmnz8M5qQcCiVuefC+0PkpO3+zJ2goLkkBn00agGHsTxAPKI
ZsPVesYyXzrbbHH5jOp+45e+290GGUpnrTavzaa9oTdR5KNmW00ClVtWBowMionl
I+9OBCX5Bq6pAZ7zP99/WMUfkOHxojX4XgfdcbYTIff98wDiHEZJ+zy90/l6StAV
6/NFSNHRhmYUDPKLa278h7Y0JqhIVk6QokObmjQTrO6kRTdXb3AQPHhxHwOndRyK
2tReFberJTQS585RbmQHrACPGA8NUSgSGmPw5FG1wv5h4Ei50W4c1E5UWDeK1VSI
gVM8tqXv/FBnAONNz1hvtHPeK6NkUzuXqcDnCBD+0e2EYBGZLbi7fMQxjAXQtbdV
/n3DR4iwzOg0LoRs0cNkzwioy77jqZKYDm8kheaCXl2+EY/+ThDU4NqFP42zLaBl
z9yWIwFzR7uqO0J8V9PRAEKZ5Gc2ULuKGiO4HnWnUCOqlu6EPtdjcOHQs2tj1F/E
g2rwlHVo4JjGfKMg1ir7tdBuR63cmrpXI76SBRESIobtd8R5GGjI1xvOVczZmylq
oYdK0ZkMDgO40PkFCWH91UwNkyRIzoND47LltYRk22pWDZ7UDf1uMRN34fPbj9sx
fOQySzQ+gNrhE+gnvudZbC38skhG2IJAILi1nhVR2pXrvHSGBF6rioSMRudl0FmA
AWLsRXAy/L9hKz0lp+2yfaSaSscUPQ/nFC2EJZEjIcr4nHIoP+kG5ljXU7Fh07oJ
09qpkL2IYm+nexsvd69yquEuJEDeUP5TskABcleffD4e3SNyc6Nww1bbo5CwL2Kf
nW8H6dSsHQcq67BOCHIc01e9uyi/J+uTFcKBlzdqT1w15oBg0IW5Ecjc4F+82oWp
eczjiVWlwUfUi6Qoc6ILxWYOUM3UQq17K9ahKRhR4BkX1oIxtEyctVsmF9o1Uo5A
bu6STxBgzHIKWwDC256d+Nr87lKgMTs+H8NZbbWnZfboD8JbULczUdjPZ5F1UY6F
Diz26ziBYwc3Vj/Pxr312WVlP4QTWwD5GQXyF+T9840uFPrfQgPJZsRyCWZTcV3L
/j3FTxAMWNTvM8FEl0a4KRR2HrUCEcaQb63SOeYg6gseAgSKgSURamANrv4on3bZ
8a0PsaH/X/avFSEc1rcBMc5kkv9QRToGeBXGQXXceHNteW6A69RVe2q/w5Vn3Bib
9moxTNg9oPPl2nM+kDjSW2ilVrPvU0y2HhcimwH2sJnOWiqnJTc3ypEjBA2ZR6Kw
AG8Qs7ynbbS6cJ1oYHA+RjoQ/ci2ouwRnrgAv5b+3E0MOPe2vbup8xIJzjcLmLJv
TRP26sYayoCypcaXlSAKZAmwpewbMdpI5wTdx4mDl6pWhwZ7oWTCOz6UMMi96nVo
dIYeqC1973N4pCEfJXmgcW3mSYcDfrvlHbiKHIyTWEW0M2gYLj5dZ/hoHWW1PTUh
DMNVkgs7D5zUimHb/6vc5Zv/+62NZ0JQno0K9mYDUGi0rRY990uiws/1p8eJnNJN
+eweH38Qk8oRx+W2qNfNfiXKmoucgbWIhVXs/dZPFsRd0VTBpDMy9KGiL57leksJ
I8yj+LuDpBUnqNFDYS/ZwEldDwKnWmzHMM3wHBDTRYgMRbMEVkdumzUPHnPhbdiH
7gHBtdcxKZO7A5ufjYWA81e4ke9dqwma/yU2J5v4JmduxrDr4vB6sVZ/vt/qOWQi
5F0lIr+YtvgQ5J/BvrdKe8hEPWRmH9DhLP3+7+iC3EUKFK+Ia/z5rnF6xRyXRxX+
vrzR748r0qElX7LnJ2gNyAZfBvnvOr2LENUQ8chXzPsW8BZgbzB/cKcRfQW6Er0e
Iff2SxE9ZS+vLxnsK720yiG8JpMn2SMInOqyz3sPde0G+1/WbWx4HNhK91x6T9EL
z+AJdDJQSWmkGw0vzhTM+MRVbCU5D6HeogqdBBLmLTDOXHKl8cskHsevY/pVz50O
TUpEkE0yPw1yL3DqW5gAWebxpqcXzhOMIa9Z2KVrIHtWdyGjIzhqIo1dmqacmK1u
FVHj473i5Kxs/f2CLyCZKCzYCC69sjBsHvHZpOVxVlkOscy8RVvjaz3K9QEkimue
k5zJYCSuHNJho0V9pdcCWVLvaPD9KFJYELgI+wwxJ1HdeVgj6PDXd2BkOlJybUCK
xnFbJEy1RyOc/P0VfX/PWBJh1SQkTiYF8Gs0/CDEBC7hgfeyYIVlfLaveUag8pnm
AvsDVUsmB1OYZl95J8pswjv2E/EzmCop3CPiglMkpLIVg5JVzzT0iUeT3izavzH6
h+H/vw08wgb3On649b9xuwtmdAmDdaPZIRmxKKztfJwXcmiC97ngtlTPNHKtNLRG
oMVirxSyVttcs7esfyUj/yEzPPQgv6s+AG5/p/CGRNCz+dmdrWtnNzjqgEFRy2Ye
d1oxLdR2QlsYpSaYW7gbps7HaEPk+1h3P5I2jQEc0uD/JVHctLm29zqV3zB7uTfq
D8fp8czpNWfyM2/6EpWkzJBzUMk5q7DJJi/FgC07d0lUI6eOkBd02Z/qQg2ZOTwo
PVovkdnG/5IS6gJ62/SwmfPAGEndvDYv9ME4x6MolcfjmZwgLmOWE78LAK6lrEZO
lB4nRsfRuGt9wPp7r691TTb+z8d+/bUW0VeEKrbhu0Mf4mC4KbGfD2E75mme+PoQ
VZ1B8g4jXyAX5GKpLyEwPSl2scMagHcSlTbnKuKKwhQsF+OdU/Lajg8mamMs7Gu1
SeNHFHzcsWpo9Affg7hKhl5srBrhaOO6uP0awCxmZushQUe8dAtbv0zHQoLSYICw
RcfitwePuxz5W2977nlc19N4Nq7IQzB5rAzJM0182qzdjm6ww2j3wlYFctP+BpR1
fyJD8/O24aWOfya25DOwD951Vk4Ho7IyU1QJKR3HPQlbh8CjLKVTFvd9PywXbyUB
rLObq8IOD3J2e91Gx8PBdcElF4ZYh3q9jE/u3cFB3zXpqd3+pDwDSqsrrGBFv4RK
iKUFkHxK2KCemg8nMOfwTy/2QCwnjL+3jC1UW5ojBHC2oA/AJvhiDYS8G53aBJ97
JAtxCo5X78dq76bL5nWrEoPu8sgrfg7aQp8lWIbH1KDDhhbv+gj4xUSj0oa6ZKPF
+sbLe6vNrb4rweQCR9TRdpjoXnjF4vM4Yf4tEbWZhsFwnjQ9oR2e9NTVtqDfFMzl
ACoBrYz0690v99x0eRazEIEgveiwmhEkOp7JvLEEch8SaDo89JIkFXhFNGIVpS6I
0GsDcxmzV9y243Wyss5z6ftihLWVMmUAam3YK1NB9kyz1Hued1YdHSdROWhNW+KK
P58CrfGDFsXSB7WxE54YKY0yF92vNUjJ2/d7fNmm+v4nt9jJrP1aWlshY2YjlfJT
4qaMkuP3aRhG2SKurpRIcEd7oVWG64L8H8AemGRtujEaxmJ588DZ6G3ra3UMHUbA
igxU2OWeRGBiAV6thCbkdh8O51X8IZpHb/r7mIgrrtrhIkHu9lbhaFheWLeVKMjh
SBYR/U/nS58v+C9aLHfhPuCDb/4sxO4ReyZs27puMRkhb/OWUYD3xN0XzJOotaB0
AZ2IapGHlAAXrrIBa+8BrJVLWLVAUnPtFHk1hpH1c/evCCE3IWblAwcL/pk132+R
//ZVNa5VoWRhEOJ6WHB7046quuNcXGR6Wff6bk7++abe0jEMYv1o2XntqczC6idr
DIAi+y1lIWkwClt4DZ3l+rsD2D9YEk80Uohj48xHuzvR91epw75tNbHCkZO7uh4N
RoabEXh7DFKJ5UVu+EWmCtvf1hNdmpIk1jLBgGuilBAU0RIeoGs5B7c2/Us/9i/M
0Ausp0W5nmv71jj2sUExicjt6pe8MNeP+gkoKWMNRqo5M2LcKGiVp3Ki+pLh++yn
SsTFBeeeCQVUjgSO1H1IRYKYzFjsuKpORoXu8aFvcOuwKRiBsdm03zWVIXQ3q0f3
DuqFeXFLzd7mUaFSp+G7nFLqLC86m9AttfW0HPu5IvnmLdctoPu3s0QKq+s4pqJw
XWh4wGa2pzvV/VGKtMC2+n9UmgHbqKZwGhmHX1UVFmG7v/C6vo7GzPrdFHRDfYd3
2teIrLsHvJAVQbgluSeFsL6f6uPdUjnfzQzsgo5E8AySIgmGq0XbQ8TyqMMaqNYv
QEWepiA6H6hvm24Ip1CaluszxJyhKV+g7cDkARiBX469rNx5S2lbMlXpgTO/REs7
ZqwVBkW4z/uPlrqWETwLMpB1+bgEjiYzKrWSO44uTOVC7LdmTld1wiSyedJTvF18
eShP0ImJ+aK8Vj3m9qBpqclG6angJ5Wos9lndtkJXxOBv26/9RAUZCM21MlHRtkl
/6yNuYCjhvyA/NF9CosX6eTKGbxx0tmaENpjrjapITVxtwow5qWM/J1OOu3ulrDk
0AfJ/WhbUe2Eij3mamQDB69NQOYsxxs5H3SY4wGjQikQnGrMVpfOERKIHOPCYGm1
ZqSXQVxgt+N8o54WivSTBWZWy/e5SMKzQqIPtU7ntlX65KbhWmFdIb9JV9+NdlYO
8LnjcXpOkI/IzU3v/wTVkvOCqZj+4ciZakVOK6EPBEe5GlCBcjxiimT6iV/5/mPb
4mAjQcsfEEbMrrBXN6Ct9zEhL/1YIwXGnkJoIcdYRGbxcFtcDMar/J8ii58w9ZPo
qei0CAY0YpDAT3ArpNTxW7kAxIQN7YypAMHZhlX3Vq5wErM78LX2xIahkkwvpw36
utApPXyj37tA4A4O0KfhC8ZH/HDu69cdk9e9NyqZMytZLTg/do6FwOIsW14pzbKe
v/W4ywcxsHCuh+lP+R+wF06zKJ6F/8c9tW7pWThE4vkBMLXYq+BgBgp25rpsDRS3
meSkalWqgMhgI/h2mWwMZWkCfx3jqVw5WXBHJCOJwX1IUNmv1mRlFRpAeN3VB0d6
ZT5tqFLf4BszYQvjW0+WohKYQrF8ZwYI+bA2QvwEm4l1MQizfj6Hh46i/cJ+S6Rt
4cWkYNAW9aoMZFu4j8135IBNDg+/iJ5RY6ej6+HqCwAdZS1DjDNP9jdwn8AHfLi8
whyJam8kmscPZ4hsS6YrtQ41fEORdiOe3SX1oo7NueHIyF+gmZ2pW/z48hsYzX1F
1crcLH8tjceGAmSUu4LcIBG6egA74beeWyZf5fhRpr0pcI6flDAPB+ItZ1zXSh4a
lils6tjlhsPPrH4xiYwLUp7O/1VemA5oEtHX7qeuWx5H/dvpAFzPxiEALS9B669y
1YSrulAdIS93tMIXashvS1FwJbKEGx/LlwTbywq60eo0DGVZOFlSNqY/C25XdAcw
NiJ4GtRmYloDMXakPktiTQdLDdDJTDkmxsb+i40CKthvGotsrcu4mbQw6dx61RBw
wL5AfSqtm6WN1KmkBNEGZEjT1CSA3m+qg1idtcokMN1a85kqyTiG6X/CtysPyVGE
QnAwLzllzKnETqpgSdDAVljiGbzdzvuzgPm0ReEAJPn8J4+Q3FiTddXp2EF/kdRP
fE7PTbuwrURbKNU3d+WO1svGRUi9/9CWFfy+vOzDxAPsK1Y+sty76v6DZPvMB8Lp
QYuEICP0KsAW9qN8zaS3oik6sKZ6FpwqU66bcYc6SKpwlTGenMx0nFR43H7LmEJE
m8gIgrSdItfb2Q8cGpspOBkRLg47/E/J9xbg54lwNsI2cwK1qVEncg+FhHzqhoDX
L2VFV/+bSC8YXiL5K1HZ+bfx4+8yz9kI0OmEQIIqCExfOjePePlqjX0do1K2bKvb
Rw29496p35ol9bc6FpSLC16CU1tjorGp1JC/zVvexhxv6l4yRdhptonxQn/UjCar
5yKhacTVEpvgfPCzrq08734dOIfVCRklTc/X5A8JjKuGaGnqn3iQs4IaGnjIAC3f
u8kQcDzrFlOFkVuJn876Uu4YSj2lXgJOuOPuhQYv6jtNDkjQej+YE0WxmRWsMGuX
8LULioE+vE9SP7whvxrIQ1prmIPlXprxbOonWzPyW/HBf6o8dg1o4bjRIB5tn0J1
whaTMj59Mf/xuBnlb+g0+i7O6o2TMV3O7Q/duT43bEpWcT1H8O731yd4WdP9Sejt
ovllZvaWsOvkda37hnuQrzm8y/kJuZpZkE0L0A8oI8MSV1TK6uV+kMz5DqiVii9H
ctm6fF1KI6tJcf82R1F/L6d8zn/cgyf2Es4K7EBWArT6/atF3l2Y/UQPpYvhZZFr
lAaVWLyOQ6t4se0XoSce3G4QhL3dyyCYaMZNF2hiYIRn37AiNd4l9er74E5KpYkI
hZXybfYOQSxL82gOPif4kPp1jifjUvLPsKk1x0E9bTQFtCA7VwmjBHo/cx9VIloh
9kaGgVgVyZkgE5hxuJBnEAYsMF1ybapGMPSfsLhhLL0fm/uohA9hUB1ugQJPUFop
1uKiAeWd+11nHuvoZKdG9D51ybAm/n6H0JKy2H2bKcZXOlRbBEeVuT2CjWRDPW7l
ns5Wb/ZvcGzjBGHwRkbnFlWjguNJudbzMqKjkEkG12GqZxce8VGSua9b4CUqEn47
mm9gyITukBomOcvHwj/uYXgHIG1RPu0xoP0XG1ePPDur2CgjPcjrabKNhJnys62K
izdgiXbgPnfV4s1gI+YbImX8GNiL1urF4K2HZ5rCjAR/AoAQHVd/aQIC1hSnHX3C
Ye1nun+SNeN1/447Ojpb9Z0/23xajXk4Jc2c9x+hshFcrzNJRqi7oIL2XncxRjSE
D+ZBiucVKdlpLhcs/54Q5WfuHvDv8iyaOl+oAtCPTA9+l+Z0qwvgUgrKBtjsrt7q
yitER0+yVq0FRhd/ssPuueJl08cv8Bhotvb+kA0VDutZ34Ug/LFVuPqqTmD4TPD6
c3fR4bsqvb1zspeMrjKVcQHrgQd/NPAfUf+lVaAU2a4HiWif/UUGmbinqiVPdN9f
3DrfUekOmRGQbdHMLvI6OC9M6p0B1Xn5yZ6/IYMEL9XrTAnSiz9D4+cr1vOhBxsu
02O2NDgX5QrznO/oqVKg77jDLETrLmx3u88wAWInazkKISTybr/kN8zcFnxkzb6I
Vn7BckNzfPhJ19HhtxH4QFQK+/6ljo+LVcQxiaqsCH+wDrBYbgSdH5fnNj83r05T
TPTBjyCEw/4e/lTdBtF2HtVA5VlcVIKbPRIl+FWqqShkL+/v+coP9D1gkl2poad+
Cds/V3JyG/MPsTr1+lsF1mqr84lJMMHponmBc9s1J7gUkDknQbHV9N+rekV6BxFd
2qh5W9d2NEkR031avuWY94JmfvSkcfBgjX9w9E3QFf6HqqKzaS3K7HWdzzfmqxyk
7pt2WeXyAKJgAWZiRk1YUIU1ziyUL/iD0dG7pYF/q4IlUn6w8UuXcJtIiJPzJG4S
trym5VRCjaO8V41G59qk50VcJnkvSTerAZChZLkyNaS0/w9ngLv8y8KOUyKejf7U
Y0gFC2zv9DESw5MEwtm3QeAuLwDmaMs5p9Jkot6KiDCvT7TPNv55UjBw4EAvT2sq
smdJlgVhZ/aX2hQXQCOlCYkDB+i+qdxaJE0PkDDUK5mfvb8I3Yywnw3G4DTbYezC
TO1qbyowPt9MR5ezm/iMBDMGd7whY/LCjpwB2D7znzcAH+HYQ6pB/YLEh6qIBFHc
mnZOIIqTmYlJt3vKi56RZAoWKSJGV1W2tU3H0LxF7mdpSP1MdqFXxNW/ZIv2vZLd
ATHWY890VjRFt7p+hhBjDweTu+4zUnpKuAsvBF4VFYbtWhAeWRrfidpnFhFWLyG3
8vWywiaINRoawsv0O1Z+h/4Gag6lUE6Ox01Bi0ZBQud2jlTNen8hV4KpvOqPO48r
nj4YxFxhPgjsaK8Dy1BiRCKBS+83ryoMp440ybyeiW3j0f4eqpXFzOzpSlScLCJS
c/nsAq9pNAiGXxmd9QBJufAJqDfVaYIbTBhcr+JWUTNayJMDBRPAsNO4zEXsja4c
njM73fAegxS+tulKrNH+OJwSphsCBNMXBy1oROhBoNWf8TYAdst6mx4YbSlJPzx5
QrjJ77DzBgRGWUc2X9IqoJ41Jqjbk8MMC+xzXZ61KcDbe2frb/lhx29HoW+CMMg1
IF1RqMFvoFLgEclS2+tzMtaFga2GSPOGyfniYTVgACehvPV/EFj12m7vp4DWfIhu
BZwZLWzP45QzrglnSL2C9H3s2sGzS37yBiG6h3sZ7D/S7fo51YCY3ID/8T7NI28C
JL3V1Md40ADwZJWiDoQ+OhYwk1cKUyE/WA3LA66/WbaAcYXwpUdQVqRGHP+lGpbW
yZBH00mW4DwyB8W1/JfblPPWQ4V9mvyLoTP/5JRL7FhM8+gbcvt+u4KHkoprxk67
AyzrNDTlk1hr95AWtsan0eSEgBLYUd+WhFi6PN/Wz+RLkXJMHRESEp4vDhEiqqds
HVKDdyNYhH+V4yAO5qq1YcPec+GwEDwv+9tMaE9f0MIXUnRaw1Pzw0FEBdluNuMt
R7z+OX72YoBUTXpzVGAFYDObTU4QNDiOg9nJNWU0jYkWkEy4/utzb6ayN77tNa5V
1lEDLp9Webz+kIuZG1kUjIgcS1j3PrO9xrxHtZfOStfiIPOc3d+qJuuuavuZlMAh
wqfMiblZ1yRb57RrtrBggVoeHgpsnJ5CSJrWYAUxUDCY8X2b9m+BS4Lw8D2iJUvO
gKR9Gu2WT4gjIYsrBdu1hF7UzcMjioPCDbAvpCoiBRpejVaqItgd9p9Idn5If+VD
iXP57ycpGzNVRZdrKmHVbMGtrO9sQtrGWrola0mJM2zRvWJOMunbVdn+CTiTHYB3
ao+shmX+v4YfdIhTOR9YMbxKGiIjFAKS4s6C+XM4tx6ZCHUo9IkN4QJB4rH7Br/a
h7O3keDUySCntk56IJqAJzgGwIv9r/UUxJRkTZ1kbaLy8WrpsgWz7FxA/3+WBivv
3sUbIxt1RbAR4rkcwJJTaYODeNmMemSK6GgdapanzOtPzKbDYfB8TzVjrWEp1moh
jHuzmxk5yfCeq2he8SFwRXaatz/OhslwNRr3wbflRQq5029C2goizpHItxTvy1t5
OYNsa/Vy7qZ1IyM5MNpBJnDehun2TU8xB+H3NaMUes5MNLl21YmQjMNkZjAcqor+
YzLvFLz4IsNErfuWW+U3oynwfPkl4SIu3cpGLGPTSTYBkB/pbXtKVBnwu8YQp1j4
nFns3dRBs3M9n8sEkjcp/VzsKr5owKfGWyV2V2luW6TjtBcI67TiZ3fF95FqGY2J
VkZwtL1HV2cyToRaRgvryz84/QuzYa8nyRLocbm4fOYzt8GhCWnO+fqqwwnb44pt
xB1b68RVdTx7qHyggybhv/m4t/xo//8AGg+At6LHkrtOnNHMlPLePIKcvAHY135j
sIJJk/bQbFLtDh/HyFuKkts4qkc95lGdb4Ps+NXSD68TWsS4wZQ0WyGVWXpCAyUz
oIC78xoqmPF9Ot/xn4zrCtQyjFpdN2rDiSYdfN/CiUKxXzcVkzyyo5Bz6G/C+VtL
UMRqm6yVARHYJatqe34cx6eyO06xKU5SPc0Whcbwmko/4kjH7AtrXfG6Yk6eSTh8
l0ZjTG5fQu9cdSOt0+Ovb+ZTPA4k/uUmLUDS7slaLK1KbBTjdJF/AVwkHKR+eals
rtQ1alyQ+QxcOR+KAEfpzsTv8l6WypKKpmrdQvzSFpKXivFXFj39M4wYS4P1Uubl
sT4D/3ge7Ania6fcaNNkM+y+1cr/VnaNHTMIstRGb25gBO8e/QpUjgsmJTFN94oP
6QAgbeQ2DJNTowVJw1GKsCNcLQs7U2DBXy8aShPVO062c4gVgmlxFwtem2m+cgoa
H1PRmas5Gzjb6oR45eDVQNzTYiaNqr+jb7zu1ctaNohe7vroP1/XLLFgk/fJpNX+
7w+TnF60dbE1Sh2HkDQy3Z+gMYhtMUI4dRUBbL+XAO+7/PKrsbBw4UX59R864Xx6
3xEdt+xe5eajDxKj9H0Y8Gnm2nEYqQyloHFb9RIZRL7DurSuEHzj+Xb9w03/U5RP
qEYMImivqycq5Uzssrlf9c2IeZI6NRxSyQPZEFUJq46HepiGHtTw+nYKSkfS6F9Y
vsLhCjXiYp5D9LUVHJve77qeGnzBalpn0Mj8VOqGhTndNDTrkZIRZaViiyLUjw0R
gg03cv1aqWfx8v5MptftELjp87VkUrvyQYAC0+KlHT2fkabK/BQc5L5Vn0hg0r41
YzKfKuuaY6q4sbKy94rEDp/+2h2ek+wZ4WrzPxkebe6NN9ng9sKGQ6Bzkt6eMMwP
LYFO4HTomI+glLypujvZsrx3KADN8cYC2GXNMOuUVM46ux3LIrq7h70i62cmhXGp
uwgxf4ujq594o/8y06JHXQoHYU+rnr064EXd+LLX6iabh1VXVjREpVMkImT8ATsq
YgEcR9qYtOMNrU2tuKRGAYjvwH8nfH0y1fEFa0pF8PZ+usR388wJFl5hwWqcr5jJ
XrQxiqRihYktUXGvzVMZBMH0+5AbroQLHqTOkv4zEOWuCF+bNVEXiIPUsdzFic3B
bZ3VsIb9Mi2d8XVv6YmQHcNqrls+Q8+95okN4Kn2Cfi6k9VYNzVCvJHlMYAHLLsb
jXD25SzoptpmLcILNPAiRaKYVsYEgE9XE5ux9FQjttxW4Epyk7AUx1ZnzfeJ+oub
TH2C7DsI4SztV3L6y2bfHQkrj6AXMQbxjg74/U3TVVgL8F/THeP8NpmxqJIy0bTg
wLvUL1FzQvhN3yAfreMh+ijzfk2rKjL/+OsYUWufsbWyiM8L3wex95p55I98At38
S3FSTXTNPgmosaA8Rj6ndP7QHVTphn3GAmoy942w3N9CBwe0iyTxO74nph9xZsUN
t+2R7K3DhqKKs1AQV58eYWvnTWMZJ4vgWF/+z2rK6BMIgYN+G2aK6ZNA8//YRdXP
LZcSzmVOyCFdwxRoWa6UiqMGBGzikciJCx38peDrzgwB688fNVmNW8Etp5BUmFx1
f4A6q4/x6DahSwUzv12bxoNCnIghzYpIgjiArazvYB761n8YwbPJkkXxO2SYsQYQ
Tbt1DZcpJXgod1AGhwVZngBgsgTTaRcOVA1RVzQ4Nk7omrCbM0U+9B8u18D9XX6e
/EWBKgNfx+lFEKZ5VSL34Lv2NqNffGjysUiIgsRS8qGKL7MGBbvkuiTWorT1umGj
fFwa4WqiyuHdWJsn2BJMsYog1KRqCJ/pIMQgOXAtzOl+UM6NidwqW+W674u0lm0a
o90Y+9KfCYCJBvxKHGdopo24ISR10CkKLxeaLbhglou85AaupENyPBXzy/VF5qa/
caKEMrIKjyR0ExDkI8ZoGZEU8I4HbczEm3Vo9SY/3vZqbWAzYwSTQQKn21q+OX/V
c/WAtE8BIIaaDtR/C3NMaDL0AF48Dz3iCqQp9Yf1/fetZjAfic+brO9CRN9xQFKL
lWHg0+Es/95EIDvT/RRu/KEYrTfI+wpx38ss6v2Z9XKTH+Z440Jb6DkrFpgllr5i
eXGpe/A7+BWNdNMWx4vPt4G453pocrX15a6H8rwSQgo3vZ5IISmwcGlvyZ7wkuC6
FbWl8AgsD4T+vLruuNW9xpWQlANOTkxOnTMRkHqNQIdn3ElIubYHYUg6+25JVmZp
JCfCzwwd8vEU6IJ0lVcUn69SP+8JzRHXzRpRW378qILlIyr5qj94nGj2rFAZx4Og
MiiXAV1BKrOtXZzslAX4KP/gCJXV/7pHMW7k5QgOGMvQ1DJLfbLr3l0TqIOp0xox
rFFenV6N5iyOw6Fjx+rkfqu6ysgdxZLFX7QjYI0k7AgyTHris9KR+PzbA0ikuJK1
nWVhGgA3tHbfse4cxmw9aKjjw5xU74++sz1gS/ZFbtupRdJvvHPJeR5S1MwceUfV
JN0H2TVfmNAA7/2VK+QWVpSlHH9BWzKVJuAH+vpH5RxFwMub/OpXNzWYeAW60bv8
czzFjsRq5/2+jctuY/vp9BH0ZZRVnWxOiIyK1tvvZTxhJn2C7AfM8a6uIqjjVm/z
V1HwFykNFD5jDj0d4exs/n7TUpaq7uhN9de54N2bQqjpnFipAyAidcPxRCiior1z
42KxXPAP7Ae8PDqx9+z8C0EpOLYiY9D9E6ozUASWDvJVjUcSJlkMKPn3TsQAMytr
UQzODCQViJlh1jl4vIAuwWWv6k3tQT9ifoqqhwUvSArRd6+Mu8VQyp2uEHtbNwc2
tDUyD+7sb+/3uL2B9UKmQMA+uj8ceR6BA592icA36VQXt3/Arb/8G9IGRuWdo51X
l9ZoRXIdypHnRTnh7WI7UnzI/JhHs1VQXzcpI9s6pyfBu7GZ2guUSddor8xVFLb0
HDP1eTnl1t3lhh3kUu3JlaxcOPUu7RQ46ipqkx+UeARmZXlX7m+I+Aiu0O1bA8VP
gfUijYo+To8vRq0HZDo85ercRSVOKKV1Un4Ma+Q46EBzrx+/DpMHCAewsvg22nev
jXFf8TvM8OR5UAjq4SrXixxBv58e/CwuKH92OBKq3zKF0nfMlyqn4tkugsKbnumC
0LYIkt/CwMNaLkJkU0ddpY+KlFI+l6bXM+yAqAkaEGWhpV0vtl1Pouc6xW9YBFOp
bHfObxcy9N8m7bWitBshA648Lb6mEQiKYWX9gLWLqm8xJktwqLzPc0epTpoQ9UT6
Z+4LY0wPgnuntsSLFKChNDrpxH9kpyaBvdI7zlRGrPUS6O84yZNWwu3bBE1e5ZAG
bcEHNXkZzE1MZvW0hW/h46PdQJxwjcU7//ec1DOrgyubAVvVN8dKJqSDl3Tr4F6S
0bbNpt60P1UlrWxIPJd5QI9mblSD1xPAx3QHZpLfgr/EshV2XeNOM0gMWzQ/greC
pKNJ/tqGWy39FkBDPdWo1qBKmStZ+NedAK3nHSVohjzAhn57bZXB18nARZIwEWgl
7d2AaM0jFjELD4khVaLD8cP0jRpf1gjx+Z44Jqrpa0xAliF4aGbNQjeqgG/DrwOW
sNdbCm7BThMTvw9rZUUTSJOZKLdCaAiG89haz2xFB5r6FpjB3riZDVgilBKYEBFH
YdMd66lEQ4e8yoX9SubdZ15/+AOf770FB31kCRxHaKoe5h3gYb6jGFRLB9iWw94Q
Tnjs4mRvRZecU0xA7khknlc2icYy4arxAVYcDYx7rIGG2/hIkAK15AAA2b5bPUCY
2QlU1qAaoe+FfV36xMSpqPVeRmXb6ixqqSEZBaCbAjBnH7GQXJ7zaGFND8lTREjt
M3KqJGzXyKvrVcKSVPWTX9qZx63Rk0POyMtAXT67ezJ3+MwSijXkPHrAK11NPX2Q
eTqDoyEf3spPG53rGxQGzIH3Sr49E77QgFW557S/HN0z+6qMHiu2vhhHyJWb/3/T
wEI4+LLnBugV5ZkHWkv7YR/3ohtabPOlIgCbcFkbKZg1CFXECAl+copQStTVGpP/
lVXpFv38JeHrGtnUjoWtz6CL+H0AAysKJwxl/uv98gwSfB2lBBbAmZ/5PXifEL7v
yZJWN7Z4F1eeLF+PPZc9RTgPaYvKpQRPuOESu/rskUD+6L8MzAqvgHZkRnyE68UR
yiGemFU02HGvoKeKErJ7rr7p8o/FKbC6+ndOzo0yPPoFoTy9Qe61FTsqgzANR7l6
kcpjysZfIkiT/JCEplnvIiN9XJZIl2pKvj2CHjM9zDICII66qHkwwmIh7+hDc9/s
jUc56PnFk+lUxXXHeYPXO7hlAJZ94WpTQHo68Y4mZPaLaazwSgxJUp6cGhyA5QH3
ZpyJNvUflhwApIWu5IBMgbABM1KxGpbjZz3R0gA7O/GA1GsiMPgHgMk7zD2pc/3t
YUgs/V0PYPbsdTBIeLdaC7FjXulgVdtv1Cqw3C6RLs0DcQDfjHB3phcQIjqRkr/c
0H33jZO1MgQT4x1v+cYuAcW7mxD7oyHCJZNxIimc4dVDOC4I/P9binmLqecsQNC8
dzOv8JWvIFxEFs2Oj5NtvC1tq+6Eqg6hQaMY88F3LGkOiftZViyB8C7JtzaqJztV
GFXPQKtx/cwQQkr60CI8wGFYKlPhgOVYfXfJ1N3TVGLCevpdEM3apAbD8kV2ZvRv
YxwgyzH3tIyKTJMmjuy0YEGR/SSnQOYSFcIN6nE5ep9HbNPhO/AoRdKZAGLjU4GE
muA/RdJWqpWuVARm2YpF8bT2VSR7ChbqH2QHj37/JqsxUNwZiJBZATw6ZvluDeL7
nQYec8Nz3vQypm4eUIWVJkAidzkipgfIw5dyysXg534Nmt+6sC3eybh5xnHjkJ3f
0OfAB0fJmUKTBxP6/wvkmGHX3E22Q8dUvVNqTcjg64IPaUjNfJXFrmgWYDtAdn3i
Gt7Naj4Sn16ehsilkflDppE51be1dkqK/6xfmlDhktaBAKXfrpj1EJ6pHFYhY3/+
lmPYDbgGhdfvpCFJ9tQHyP7dDNxYgY3rLR6eKHhBhRAraxrLNMrbYq0EybB0dgZY
x5WBH2d801OYJPO5if0LAkfbft1IZhoqH0ET68V2FvDwWVorooIgsitgXwHSjw9G
1uL4SRzC9TDFg6bF/O8mqLz6tJ43yWxKuEjzDpcDD3ljng1kn3jKNPNKMrie30Jx
Y45UTIs853pjwHYnzp6Yx4E+GG7jebpPx18+RphGwMz+NaJZc0ydf4FgF3XOPZBc
yPAOCFtuok9HtWRLLfAPtrR+RnibvBL41zjcLQp6Ttf1JFcHF2tjWGsXjlKZNupL
9XWejYggRwanXXt74dGfG0FHLnFW1u3IiccMeBvCH7yZzGyQhWKPB1vQfCGwvQ5w
55qpTs/fJ7ImtPl5rCf7XkeUCe9ppL6a1yt6ULycBvSu2zDRpdsXud6eRMamIFZA
6aRjq0voeOZy/yTv0eeIC2GvmCt9KrGCcPqwRi81PIG9rJvQPLitRFzyKZm/frjv
7qw61hyEE3nydBYBIbH7UjuomR/GwjpHAjfujzW8yFH4YcRLPwoVNcBI/x/7uqtK
iQHbdM4xZyKLKBzwMSQqx0eA950gjeVV62Ti30CEXDqeNFtmyl9r+z+ATFSysgr8
XgmHuOzyyS+rZ82lkvCvIqqA0kL6dXDEIyQnFcJyvPUWJcK8W4QeabQh/H2nmsjq
EZ0DpgLlhRoeEMHQ+cCgc/wbesfkPBCLqIkQHiWqULR1zrqIg4L035daymZvzkev
4lot7aKZhMvscrDXsqZAT3kFEUqhvh7jpJGo2S6jF4sAYV5Whh1+qMXYCONazVSi
ZAvX2X/EBlyBCDzEIHucam7OE3Prqv1SXNnchTjBg/1CMCw9Its8sgIAoKadjI/5
Uej1sb0usQoZLu9G5utwwarWwgyFzOL0rDl4QSGNmiRcTWEFsT7lHWedPfWxrOQQ
xcvjAIpY3mH/INFNQNzmVWoNzjOsfO3mFl+IZls5abj8sVhG5grJ1DTJyH3Nc3l3
1ro8k/onmRQqe6v6hALOsJ/K6JzUxSx9/+zLYxfIGpzUTUGL1we4OfTIk2p17iCl
6UEIFAy9NVKFNCP8dsbJ2qoa5h+pKZcqHtKsp+LRmIQYtiUGnl7Bz4qjyHRNwZct
kGYzlGxSAX/zURtH9NVa0F6CuQSCecMZvjw5vtlbSh4PwwiDP5VK9nhApqYC5cjn
fc6jd5YJHTpaAovPYo8YGSfZ/I1z91ejJd+aEzzQ71xSI2L+4OkGIdt7r8hyICI0
dNAcKlsexnS1pOiYgetEQMl44oyFzJfVxg/h+xTYw8s4GtiC3XZWbRQD/i3Hau96
+rWDxoM6RsxL1eWcI5MS45d+gpRVeFvzwL4BsaMzDuKhQU1PmzY18UJDyMA5BGhj
DXfRNd3R93Gl0VDMcVxfTSq4/c1twYUbBiMBKsXKus5bYG+tlFiKuA3zs3xVU9sa
t4vKV1xI6l+lweGgJrxamHEN5RVrtigwfTTGeOUA0E8Jo8VnGQQxTO+YUzkyb08j
X76rcN1FhAxnBvfrDuRFU1iTNwmiuZ5AJu5QLdJBCHFPwBoNo4kVPVmEOFywGh9u
v440OAwCSr0tP/e8iTfXZkcHfS3znP+pro4zvPsTJsoeMgLDquUlzPB1pkQruDcP
t4tGjDaNqu3iJPUEj2dpgG2o4K2in/dND3ybR0IdsCFFWqpnXd/lDflhWuhnPg/z
2l0fg+INFX2YoBT0B76zP6dfDxDlRmx/1bxWpcC2sZxGIm+sxHUz6AtNrDNkKpfV
pX+c0mEccf7kK+UGDFj9URFbBBMwL6gUl/knnG2wQBtLNG8sT2H9wrI1EBNhNOAn
jtZP2iNWNG+5DtEfL1ZQajTRyEFOHN7RaRnXk7TUADB8427ZCduw8qxcbXxFxzO3
9p+MVxz7wDXk5sxwUv/Ood+5IVVjBP3MXE/+mXCPvU7so39kNJ+WMpOaFmLZ4f9T
iALvCotFLPnPtg0T356c3lvWNvfmjZh5jx0+yY53ILOBzjtY+9LuMW3Flv4Hif37
UFrW41MBdWfBpmAoD5jIyQu/sYYyzcFqVCO49gLzUsfdrl248U91bwFZeV48Wyls
z4aV2ldvMLeZFqovahrIsB6Lc7SAMZqN8ebggVdUXgeYPbRd81jx7O+BK/CQaWzi
6fX4++o+sQIeHHR6JEqm/hZnfGRnWKCSwavli7d1fTHwwpolbagik5scJQSuMfN5
Zz6QMOyLva6MrYx97Bih/vg508x5xbjyBHxdmJH1K6bgN+4i6FMPXoYCxS5Ibhxr
p5LO6djic2npVjZOXuTlfAh4ZG+4oXigfa6IaVmaGQpTV0G7eAYJBEKbH9Rp1+w0
iThlZi800GL9CeUOe/LE537EXWjnlH5ftdAg6k29Yh2kp98EmENNp8ztKj7FLX6l
IK0fca+jAtayM9RzveM7T/I6QVpU8b9NRIgWswhtXPNOX3fyTFSg7EJ9kKuFSQ7o
iqGbPznCDyaQ1E0QLWzLsZstvepyfqI9FNSTnUiOsUYKimBLr0tRwo2O2dpPFDpD
iO+6gxuue7AjhuUoJ8l5ejbuCo4odFiVk1C0gSHa/vTlrHuetZxXghZdWF7VVXPO
sS3fVB9+rO1Z81MtOdXeXQdehuuKc1+uQVoCQiWYjzcB9wLD5AXJ6xHFoZhW316U
H6offUDWkinGnDgkggIiNoVnqnXmESeUQQ9XSx3oni3vreyh5E+sTAFej9aMLFfn
PP/Vx6m4eNmFEAWfsPg54T+DJpruxCI6/n+ya5h8iyOYvs2SLgemLWe2h5ircYqN
4EH71Pf8f+gXH7ed25wGpOYNsFHFriFXlun+rViTZFIRgD+yoDuWsKoR6csSGn4L
OM91KL4k1TjTkjQyPJSJyQwhtOiFTStLH9HSSJZMWH+MbJ5bMPpQEOE1pUWr9RPS
ACLljuHxhFNwnDUXHdoXRtG/A2oKwDjBG/RrkDdct51jh70Y3kxTH9ivqQRn3pOp
cT+WWaGiS0TtGF+AzQtx0ubhR0YdcBnXQ5GFr78a+jqglLgv05VPw0Oy8sKay1Xs
2On9245wFzPKjpWiIYnUBRl24W3yA4YlvDt6O0SNY0ZuXsZErc5KJNtoi5YAgXB5
9jTXF3bOeKXewxx0RCWDYgX748tt3ENphXkmnqLlxDUB3idKMza4Kgy960c3259f
24JFTZrA9WREwjjr8sXsN7qUl/RFDNbQZLR9hEjpn1u8lf0UBpKKdGKrlr+ShXHO
FG5yqKBacbYJoN6zKbnKro6QoczwY3KJB12b+TdHQQZfGax24AN08f8qlepag3ur
CjXi2wur4S6JHwRwxzdYoPisVZKHlj9QmtjNUC3dMxkj0fK7ZICGnko2h1hxNT2h
YUrmFZPus4uQs279IU2nI3U5HrHhZSSHUfWQ0gPTo5acexKj0x2rBuUNThVWmeqG
o1WPIVLwRfCRhNVcWVufzZkTTqa/SUtiM53w896opJTKcCi7OFHJFE1skiqCqiTg
XDLG0pzyT0kxSyzJ1au4Fu8GOylJ3kuySuBBJkTVSVarXHMFrbjgprhGsuBGobWX
xN4SGWrzkZurvDlT0MtvsF7S33fXVYhL/GaoGnCoQdRM8ZDOeWo4Kn4stMantX+m
LMpMh28/+8d1jZJHJCIDmbAnPlZqT+mcDEupadKdfW2bqF8ksEjn30/wBHAZtiNe
X6TJCaTrxLZlcRTId+I3iYlhCjvlDu9IYzT9/ENwlsNmYa/07sdz5Zfm7NPJm+nq
5ao6sD4UZOvan8AYjb2o3Mujp8YBYKwGo2lONTyz3X1p6VhfNbnq6xMzvzInudQi
ums81EJgp33hqJvwlFvoGO7As9BGPsiBaLD1+Y9A/wfT6VYgBJu36PElcjT7+R7y
6sed3OZIQsEs2iv92kilgsamTeYBXRmCmumM9TiZGQKR80cCNQLAfqZCGhF9HgZS
FeqKsSpRejGOqQUjdhYckQtfxJxZ60Bx/Ts3wFUOWxnxDKSQmSWRM94l8YU2SMhb
JtGI9opiCMwlaLuxqNKcBTinUMWmP+LhpoKD0JlgyHQ9ZnSsjGC8Rt56iIBnTkF9
v53WWW9rB2GAO7APvfUPNPv231opQyq5Ia2esBxzNIX0iFR6C5NG/z0JwMHzeh73
Z+M8iWtCRBroM/VpgLkLUQB5+fLuAcokDvoQCHE6EFGHf4+WUQW7tYTiZqPAUvby
NsY2CsiF0Q21iOfNdeEIkmBfXZsGEv444uxh7nSujebPbCP9qcV1lJpImnzod6v1
DcFxqkBdyzagI+0XANPRzCrgUuID1o3lIRxw++wsq/wg9VYpjKK5BvCPjTZLXbDj
bsLftn7YGXDYg5TRsdiPj9n1+cXfPKc0K4AX5ktfKSVVavj2JADJqUEYOavg5H8a
4Wic5mUVGBlUSSn7ovFcCFY0t8DvjEQdq/6CF/4WQkz6BRFhyr4dc8rxWbEc8jhL
eQ9QUE34LD2kRN9VAOO2NjLgkGWhtNIV1U1wvTa53w7fBLojuDmpTHUQ9qpeHqSP
unmDXTmoU0g+t0c0LEjdF2a131aykKBK2JQrLQRD0axgs7v6RXJLXZcv44zu9nFP
Sf7qdAgMSt7FNyrIR0E1Wl1eie9CpcnMZdaDE0J5gEEA4RVPILeR75CCUwn5J/gc
AdxRzq7NyycoLldwlMmx+0HsYnHzr0S+D08uWKGKM7lFkQ4qzbjc0rV7KKotAuyj
69SHhjTEuFUKrT2N0xjVQZpy3Y6REOq78NaRbaDkJrD1v8tYEsybQyaK83fJhf33
9qngSc5M3o8O9H3Gkt9CIgh+E7ZJsEIpBXHgXOaNUit23il2CNnjV1ZOO6DeKD2l
nlADP74GVQMKyRQ5e9S+ssvWvPDb0O8SqYlnCEPVuHlo0yiBDrGWSD+nTZjjA/s0
ZqWcejz7F0X3nsOjmX//pTChZEZ9LVie2FOqGqFMjlCzJdzvSsz7aqI5p6oCObfB
uvI24E+koK4YRUW6ixeiNeYEw7q0Lvh5/CDoYuASX3NGeZw0iiknVNLxPSiGb+VI
Cq7t4w/lAsGK0huI4XXidH6ODhBD7gyHQ429ewEbKj57ihGhLkFc0d7tEa30LbEk
CJJol7ZXuRhOa8+a2ls1sZPRtMC0emhDNu7jFahGqcpq2GgJ5sf8/gk5YHBOOybc
8IOP+F2D0IZ+jyJ4DXQhg8Epxifb+5xN6gA5e4fk9Sr+tqPjvUrbATOqoHqk+OXf
7OhCmFWR0Mxc89K3uerqStev+VU8pu7Zi2fje5WCw97lmqhatWbd6d9ls9H8vMi7
U47mCK4fX00tNPyQyOrpsnTsgESNney2BkM5mtSdU+RMP64uC1VkUwc1dUQTek58
mu0CjFDQFNO3l5u+zgwQoBgmkkLUKtbg4F6bJ39budP0LnLi3zGkieBci9WZSYq3
Xp3e4yQhEYUChfO0F+Q7ALbbhv14LId8L93TnTwJBKsAh6B7XcmYRVEUzZ+lNwoB
27lxJlGjK3rpgVv0sh2PKY/MZMIs2m06csm0J9xpfxPuUojpUUamCsA4jiuIKjAT
l1q4hC+P5XhxQLhTa1p7H2oKI9lP22a1XOOKKPg0QZv0HQhKRI278uxKu3q4vg0w
b+5tx+obPiULbI+AxyH2FehcRizCPXixhrOW1UV3Qhwezk+Tgygj/s/kyn0EoRqi
iDT/m8wK4eLzzB0hq6+0Zc3GU11THUZp3ZDqV3s8fgkh4snuX1jzUx4dDoe3aYet
BO0+T9y0G1xgqtZgovAneI0IxgN8JUJpFt7shh0fhhqQ1Z4IUiSVYtt9qv0TSg12
bwJNCaZ+VzPh1fDOlZJa4MGxWZTsONA649CZ9Pi7emIFzbrPWuRkaVGgK2PgjMTd
8taHtsdKNdnWh2omDnmrMT53aQQh07Ityq1IlHVQXWGcsK82xnmzGQiyFhs4FA/B
1y3pkj6MdVnDQSpiQ0kGwPFChuipS6DFQua33AKtSRM84ESAvO7c876dla+wELyp
gnIjvzsL13woov/l4OQ8L064/wNXh3nPCd9wvSs0Rl7xxQxU43YIvBfYCjZbF1hJ
4ZNUm7lfyedODmgYZqFtSaJzFkG5IaN1blxCLMEEfj05YwXkmUJ/7jDtd/JLXFOs
CSzM1V7wGsFLzaKrwZWc31xj3KFx3OwyhlL992ihveBnXwQyW07lLCKCPWYRemfZ
+8EljoDRAZ83cwRYKBTKLP+LITDoJtuS0G4sypG0VY4p5iDG5xw4PASqB18bPA+G
Gckkz6oe0dFVJ7x547cEmhQw0f+Bn6D8tpKBsN99Neq+/Py/HUmg7PsKk88jTJIl
8VGsxOBDa55H2QcMkHJMd1XM4PX0oQsFL+wRsrhL9Th8hEARnRVnbKQR5n8eXwhd
52CgBeEClJ0VW7RuOQs6NHf0Mu4k7nYKEYJ2IPhAq9gwgtUCTq8sVveWLUuVKL3X
3+5ToABnZmDAHqzD+bd5xFoj4+H9W70EPbZQAZ8IV6UhgHHjJE3TIqJijwxF+ENg
EyPBNaymL0ptewHj4o6aNs/w5v5V2ReVStzgn6l3wJtJdVChOERULHiHmOtbK204
oMWLnssnvTTV5pVlyzkLqknG4ebJ8c2JaO0xzC7zBc7FzdenUqajrSjBpZPp2/pB
FreYFfgGK08Wd9equ2y8Rgo/ziwwItyylJVaqwCxvPCqr38mPZE1IdKnJsuFHFVb
vW5hj5frvyHd3102iDJjdY/0DUjp6XY22tllDY4p2Qh7IbK7K49/orF1SpswAzzM
rTthhqh4phAPMQaBi57CPtZ1H502hhWGQ5nUmandemVht+rpXyx5Rpk/jjjcZVMG
QxVfaHLfJ+OcviN/OZ2qLO9sywu3bWny15QUuyr9o9Jb6vK4hD0nugUSHsmFseIz
Eu2Ov5/tPpj2egnpErfN0FWlhVBGYRjxz74So7bN5nDq3BSlSzbKDN/MUS9pT15E
f0UgCJ9xG5CywMOATifVnGwofN2YwypL5TnYXaVKW+/v283EFlEHoz2LypF8oMqE
9amoDat9W/0XFYlyr6i5WqQ3XmuuIa3Y0Ivp2ML9gwFtj43vr3MC4xeOf/oi8vg+
XHVqYB0/lXJDVaDnQue4pN5lyqDm4N9PLjE+huHkrH/CQaEMtHBf3p7N86A/+rgM
s//yfy1Rt3vkUyPkF0GkAHiBSbvyEDjhDw3H2pPMfO+DOieQePp7jEASrSLE/2/c
E19FBJXuYWVQd46q//31MrOsU4qCkfvPTGKzu926wBDlKEYtODO+NuucGHZ7+RwT
uf3quuLSfv3bCAT/xBxfVEz1lW5UsQwn/P+o00TYBAOwXieu/+v6ibF766f2eaPt
P/4qUPLrVp8cVVqEkoqKsdQDsREXM5nwqjpLCZ9gPj/RCEuHaNgEJA7pQcBfM6je
uTtsFFDNbAgtJNJajCEqWA2o2qzhxxtGQkAEAvztewuv/7cbExpskW5pNKU5jy6r
8tRzRP5rj4vpNpqt06wJXkGlNu0Z2s1juptgoFvLfw5pUP8rvYUoifoz6Sir3+fW
X1Eeg6OQFuCY5kOl9Bnrn7zP6jHULZT2DMIhdL3udVdBSqsHSV/bYHS/T0Qeu9OI
ITzQs1sIZQEKFCtGwP920PQUzq52xtIzYg8eSYl0Q/ZJ/nBHrVql7gvVNQ1hFBv9
Jx5wn8tlHZXC3YP4qTNwst60wGMh2tDcxgM6r3GjWBbROhU6mfxEOy2zkoJ7TrJA
dWErL6oghzLnr5HdkIlRAjm1YCxT/ysItWdISkPH/MGXmeP5knIYJBcN5Ae/3OPr
SVO7DKwDaiPIwxegAlTp3HfOiTRfdOMU1TXyiFs7FVY9+dYCWpw6NSjsdJAT7Qi4
grUwkwuHSm7DIm8bSvT6hWaN1DdbSxNYRwh2JJNG1ghW2GrRylp4WUK6mJ+BpgaM
w8vvHoRrZqT+XHgPJ32m391QGKzPzNNu24CTbdfn2fNsdO16PcJ3WqWIsBwnL8X3
Zuds5JrODB8gXyBoe1QpqFk7WnLwMIPbhnmkKE0MDNCYYTtvx5LPTRrvEcxoHU0m
oYY+vnhmRNs3SN1yQweV5ZnHSWnFbOS/6P5xwAv6EzOFxMmEndnroS9CNXVTdirk
efHcsbeHEukXUs5UYX74FaNVejC9SG9tvc+0FNF/pnnqaslTTrZnCyezo5fGTTyS
kLnCgQx/EphiF3xoq30DG3RWEaZzpZbFXiRsrt2R5EZlm8c+o9ciVRVWVM0oN7NO
oV1mPe6Ihl5PAE4dWY/ednqTwRsO3EDZtFCm13yfbhfoP+4hmxREo6faqsJjsVtG
nO+Yo09HiaD6eIYTovetY38f4LNJ3nMBTNqDLYN9dM+UAJXZWdO4i+fqh7BUInJh
nIt+DgOC7NaZ6pxX/SphZJNFi0zzgPuYnQhXg7o6NFcfV/+mBrOnSBN+ubZZ7YF2
U8wpqs55Apz12UgnallrBizL0tahpGsQ1NS9+cgOxq77Iyi/xYLraDtxqOdy+Ta/
tpUnv3q41Yfvbeqog5I1qKWPtLcrxi5qsiLW+AEqs5TweTyioVKPg9MwbhwXB76S
ZGHK8EGJxDvC8cJBg36Zm5JqM2yKOA40s887lSCKnSeKZstPkLS8YYMT2Rq+MImk
kR2bydjmIPO7m2ZeA5TIla1K80Ha7+QJMDrK4WHLTQeJt6SP4yOvJmZmZ0zlgRsE
6EjN/FR10BlBcoJrlpTJNNk3EBI7wMSpyMGkKksahbJsr7PkHlLD8ERFZjk58lm9
9WdS/1Oj53UqimL7e/i5CCc72aORo8OPqQJhMv2ojXsIcD5yfFh9oYZIk29SsKmn
I4CEQPVn7ol+O2U5364pRIhp+vVcjNWPa6IqPIbWx9bD+UD00MqQEA0JqqX22Gnn
0I+2pACrGLk/w0SAK4oR1aLigarjYi2+6Yo4omktQ0ydVU4dVxjcqLFAbkUUfGZk
SXEdZmUhLqHPZ+8CItJX8F6++D7IQ7dIUXpFyYkSgqmt7RHAPP09RlsMWY9K/8KJ
v4KRy+yppkLuCOVEnMpC2Or6qzcKxv7DiQXk1N3uMgyN1gr5RWdFqCLOYPnH5UqJ
5FqAkz/uBe/U8AomyQHkiNsJH1/NHvneFAIiHFxecNGvE2Ck6vv+a2akbOkZVW0+
sA1XE0H/kpPvbPIFpx0TfJHo/Nxp2Q1PhIBhE+s/1LEomAE7zo5vQeZ6N/XnRhYd
UhEz1aiWH/TImsiNdKxzK3I/0EnV3VbPTOIgL/3j/I3PxMwl2Gfz943z6+3mT9YD
buOAcPmOSMzi5Xr3A3ekiupPvT7qllwsADSkXd06rExs6BMOU5cQyjMXcXBaYs4N
9YYnioVeyA4QHfmU2koQ/l9jRB/SAxsJM+CXHpGAhou0QHjOZ0eb+l9/9gl/az1s
ep5By9TTgfEi6fhmr3a0Q6x4s3behTLV5kp34XlW/5L7NpBOKcVf5OAgE1NI6eJb
kTYH3pUJ2atWb4N8ESchiR7Fhvo3t9qJ9VgPR7nkEEhmvtFVq53NWzDohFvzEUrL
g9qSJlzdT60pQ4xM4gZ/I1zOR8X0ZzHAIebtSZqgjJi0TFD9ZD0fN+4KIikFSzyY
cfMUfvgHe/HH2tq0BdcgjIbYC+5oN/9GIQ201c+ViiTOYs3g6oo8sLzGDbD7E/kJ
i3d4rk0P87WUh0cvx5fwrOlhxFNY+O6KAkLv5iVfBoJ9nTizCEKxwZ77hBlp39/k
P1Ovyc+7rjeQsFTPUzyX9hsQZCnw9EC6UHq1ZtzmQKNW3+EZBRoJxnasUJJAtfWr
gOdMg09yQHmE6Bzq8eYNKZNWwgOAw6RFjmeMcLHMao2G7AKFU2udPmO3HdU+SzMs
kQ5pqe9rUwXg8X3Y37nraeKHHNVbW9sZkJuvRmahxoI/9Iqxj85XOq0FiB1U2eye
U17kTQC9UVayhZg2sYgBM45/+PldqAYuLi8BwHRMwp8z0hjAGOK1OU+3IcMQPk2s
SriGD0X5HA0/Uq7mnjaDqbe9o3+0It4lpthH+eDfYMzNPFUFZQl4iu2PGfbrfQkN
T1GoI8plv0FV0gWdRfXvSVXZnV/1VGGqWJEQcowaNQNVjY11Ns1vnqmmH3vc7sWM
PGkp7+b9PrMwLFzaaNXVMUoWP/u+e1y+HQptjrmLiMPMgjvDn09VNUgHWfvT6qyC
7IqejxWdrj+G/jzAR6COxrWcE9cQZz7tB6qc/ZOyuXdiNgtB5iQAuIlcTho53YHm
tRsir844stH/TqsjzF6EpDsiqj32jNvobcmbQohfPnkKvNDvTHtzLTn7g9utt4Cp
VFHc0QCQcJROiCPK858k9rD4GABIp6V3jr+Sth0Zb0FlqGWMhdrX1cUvBi4xbAor
2bG65nBGfJR+bkLzFdsaRi0BK+toA8HvId32WjTMi17UQzEwlcytldmdKyq83hcB
MP+HyhxN8RGV8D7oFtmQukYNbEVNIUMinumjv+5XHTa/RbvwyrPqYsChzG+nsg9b
y9gk6qr3cVYA/exUXBDG+sihZPRtuFd0TMN/LKT97tXpJHRzIMZIs1f6QOMi2VTW
os48H+XBg6Q6LFqGIYRo3otP8U5XZXPkN64rOnv4Al6s9F7TgRCAU/8BFLXrNztw
PctJdiH34rZqhBpgMtkY+lgbzZrem5NieX7AYWvaB3Hb4ZM9KUwyYtItQ9Byxg11
434uZYov9/ccZSzshD8rBShkWPqNNTanZxUqWwI6mcQsZXiXd4BsdfivpY0KwfWT
l7OQFKeabAtxjm0dsYLCnBBH1d8MmVLFcHrd8DZnf4rIZZlFJiqU1XzucLSSrjbY
jt+X2KTqrOgxlVTc3g9bWORsGXSwVYNsNUkSFtsWFJ7yjsIYMGtKCycFg0/y9Auo
VJ6qDSYenJnJ0QyXH449STAK/mitcV0NUpMb7VkJT3kcb8Qnx0Clo3BQpnCeT3hc
RngsI3W8vxoh0pepwdstlX3fnxMPvXx+Hm35jEzwf1Byz8sB+lVYgbAfmI3IrjgQ
N1F5K4PIv4ozVWdQIBLXX+ez9aJGcEcOpEzQcMtu780/uSY6cTpMZGnEbZIt6rGT
R2cOh7ByA/Fvejb4E1W70tdfNMn9Lzl5Pi42/Gkr71JA5eCoRPmev+PnL9uPIoCC
sEWL4tcQ1wprgKIjlx6jhozRJjk+LNyJ15ABE0XkCnPysnVud9GzOu+09a4AJphW
pNw1/GlFUV87nFEYffGwydkIweo/xi5RmO7mOOrMi88T12AsPL8myTXm4HxkKbUN
WyPjhu2Fiv3YFNG1qyoAOoSH9TcWmLcmJztS0lGfjIpoPG0jondeB1G4egeF1bXq
5KfJPHfgzDvPhGA5qtj3rj9tXqFM/qhdjfEKvv3h3U00CY/ek6EWdQXTi9mD7WzP
qDX44PmXtc3klBC95J95zPCY+QExobF/mUOW23cObunEer17/M22ILEh6BR0yZXr
YX6dvQY5DB54yqIrQu9q55JqNnwfgMXI9FzbX+wFjEI9mmhOTNyCvfhopPosAXqF
j0W2li1aGEZ4d/W++EHe6Ea0YeIFOFwk7m10InqIDSqOsMiXPHWmsUfnvwgCkAnh
60qSghXjRuP3sdSkIjXUTUxamJYC/1RvQ2aQP7UBXGqasYzX9odvPbK3F1G1VoEL
T204tzgUT1K7oYJaMW2ASnURR+yfAugmsHTjoxDdC9s90MSCgUZ/+8YZqMUS2tTl
C1YxOFkFICfY2NCU7P9asnZSxk1N5IueEs20g01BvtXsKITyO0oklaeJ9hvT811H
ku+y81bVPBw5dB6MW9fjqb/p8moTY7WnTWPKATOAw0QtKTG1a6OeiuhZvToRIyvF
ROR6PnXHPG5n3vzzGulR6LEGwk8mJQC1mgpmiuUg5ASEZyfkateoOaiGtjpNLVNb
vj/OfwbUJfSFp7jDfBl8MgUUBg/jzKespDKJCyFhblDSRa8n1svjdROEQLaw6FAh
JhESCM8gsQbQlx53tJH5ku90pkP3sMNFsb4IOT8GWlAXblEqKbU5oKn5odDzSqa0
EknSoGvdp4YWw9v6nhZrl/mofjQYZZLlfb3v7jVgaowHitRWqygNANAFM/4jpvfs
6ZjClpIAItaffzyqha28zRQe/gpuWw7PQM7fMFXyD5MjHZtj2Xi1/sP3de6LYd0j
eDmwI/x8hdPbNaDzukv3Xkiuk2hhbrxDwRy/qFnHqVL8rZ0+hDrFj017lAe+87OX
RSWa3FqNx3paTn8/e72+gA572iHn9rafRibEWsF+BzjvKYx70IxXkOu5Ur55RgYJ
aBQli/9PZQnkuXKaLaCk0g5necVdPT6S4AgL7EHS198knqHFjbW4sNGQfElQG6cA
UhTmWJWIxb/wIQ1SxMlDdQ6S5IE63pmXZ/nX89L7ES/FAzvmmupMThRNPzgpThS1
1m3dtkCiIzprTvEX4jEmpnlwtmZxF6/tL/Tu1fYyUbcBXb1/AS8r8CSBgGI/5Qb3
407QkRzqy0SwIbp7MN1IerQ8Ag/gfqFi7lFmkMGyK4/2SMF/5Uk2zXBcfWrDLj//
hUA0d1XZrjzKqB/SYxmOHJjlToqX1gFhADXEfYgvJCQkm5DI/O9lkQD3ye4EipdR
fUsdE7JDo8QdoAiOE0Soy4gz/HlGanrHFe4mV97jY3RAB9G5i46Cn/pZJ+jlQS91
n2MiysUX3Y/5sSXddoA7pz0i7FS7FPzpwWatOpwxDzKbf/EXtMoW99DsPN4OLdQO
rWsimuEo0EFBELoR5o/HNsI58FWgS74FToZ4B8WzxOOo5bEzFCLgqnBlfadUf8CZ
L00O9eLPfBvrmVjb5fMR56oC9ET5QXkkXbRPOgaTvsKducI0HihCeifosYjJN+jW
w0+LWT8q19QC57k2BWrB1Lj/2ReNN/mPjpYMGT5sdOVH11yQs7mOt6IJb08h0XEN
8Y76NfOrXfH5TIlwNc4twAaGl1M/s7yG6/r/AdPQoJtsilC/bV8StPV7PIQIeDDf
ftvN2xTe1Gjr78pqVEOww9ivDFDT16Xni8FsH7fvSecjsAhhQ9llVeeQ2tlq1L3R
DPq0E+cseEXs2Jh265ZIOXWoTWNPwIYGvsusKINTy1Oy2lUfpEl90BmAk3sD+ETV
8cp4hgQlE/XJQyupELrPKksvUasctTvF979+GFlq5xtrpstkmu3wEPopo+OyyeOh
gZVA8cGUCxNDdPynPFPhnrl1v/RrMI2p3ESrLYgHtFI6+Ndfpy6eMAOMvnMoYPBV
NNx308rWry3+4SpahSDVZi/xvpK+sMpcdQfA4y06yehB1Sk0vf8YMbByB2Ta3cbl
sPWZzgD0qqa7Hc547hmg4ni5Z0RvkfdGkOBX3Bx5D8M1/KdTKqRz5uLOcfJLZGQ3
amhB71lLjTTCznqMM6qu3f+ua8NDw2gtfefRo2mG/Xlm5qSyAR0EJQFeOX92eVGD
MCKVgWc02oXAltOjf0s34T1TqnUYXDjVb4SEQ5WBMVSdunuB8crlH6LVuVKlPRKz
t8N+ujEOrHGYMykV1NLKhdj1eZYNig++vZ2HM7+VDKXak0umLg4Y15Pf2OjS9dOY
UO0kLCzBjvrP4HJ+O13xphaHqYArSvj6WTdLo15ALorKElZdAsT1RXcajaKCPZAZ
uJx2Em1FAKmkgtfCPJFxs8SbO7dlWbY3edW7G7dHEUw5Z+6Q3QyOYdR+jsiNpF/6
DZBdY69SRB74OFp8M1njt2gfm3tWHVEWDZN4XlpgG06dF8gJYJtYeoljH4YGfw85
tahKMAdyMRbJMTZlRwUPwOBNnrEn+BNMg4pa7d7njQ5uvKoehI3CP+Rmo6xmQBuf
YYqIPDiANgq61nOfkyWtn020V88+fX54Wd4CJHzNfWTc4+r+On2mmYRa2OO4jGUf
o2+Kb+jNiQGoSfKDrkfI5daMQ+Graj/5wjapwuG3/Ucg/+6ToCyRor/M8xhO302f
DHhiUWa15xmGC106ferQ5n9MS3UlhdFDIqr1PflusrwKo7aru2QtmyHBYm/vVOK3
Cf8ambE4WjWzkNIKuiKiVRnvV5zsvyTC+M0v89HJjxiQkj1uqFDsUw7aOyulJdT6
E/vaQjy9s2WCfE0pUMDUZN6pO4zzlBT/GX6YZdj0HnTyFrlu1AHWR8oqY7QawZTT
MOBrW+KMdlWQWCkpuw19QiHBudxEHsHnjCg/NcCWtIJTvASLmcoTxxC4LfeE56ye
ZBI7SJi8iTLkCyMpghAnQ9PinQiAr/UsvR1xheWFBS/h4FxByBkP1CrS0xZsOzIy
uhQ1EU0uiaG0Gd66lcLC26caqYLdkU+6WROqLPFIcLxYdH7oYj8pQAiEq26VXo0U
LTM2ZRGR+cN8uwiByiPcazZpTRNZP9kN5y6Lg+ehZv2me5uWqhI0R6KxzZYy6IRW
wBsrIg9q5pu5krUF3nc8QtTqZvvFqwZKxyyf3SK5unDSfJGgZjlm6cygPrs6tea0
xg3Q3Asdx/2C3z1hFtwO206ocssxVGHs1L5PWiX/IjWAF4hlKMrOnTRLoPBILriv
GuZ09s4IyCReRjXNLXJb7/bmK5ZoX38IuIpq4+v+5hDS5O/xaGFA+zpHcn/c0/4G
uvSQ6F613r0e3FLXwvUdjqDf7GLOOjdNQnXSraQd0s3Gr1Sd/t/Vk0OSG87/MkEa
VdAWduqdOkrq9iNup14TUeJWqT1xp1PF8JuUHFWSX1Umb3I6hpAvGsGFdCrJRMB1
4+Cznh36H1LGXGjWMwOjV/Q2louOItNin5tDd/CNsC42Wf6h+moglJJWlDog7DOP
y4LBCXAPFZAso7Bo3GVbJrW+swnXF/EPFrVqhaMopYPdcwwbDL2yP061E4xuK9Cr
GGwlaQwxkoDda5K193/wM7MSft9DeQOIcGSw2MBrK2RJ9Co6wc2sGYAZUY01MVMl
xkOPABhmhW0BaK5by+xZb1ub16X1IagOhUPwNhAQz6l4Xzf29gjWObLvzArm3pL5
SNLnA5TEQj0XIBd5l064iVMvN7Z4LU7zGNSlJjTC499bBuPxNyfO+IF0J1Vi1Rq0
SltjPPl/aeSUsdmyf97F05mBecao/hCaOIWcbtrvPly9DQTjAXDCkMOavpCt47Hc
H3eC/HVyuq479b3n72ERAt18jYzkotlXCbwR4Ju/VKbsAMiZ73Bj8baLYim3G8m8
3dP6FUhKN+4hAarRSvCw9h/JEvD+sP9nulxOVPoGhFs2AW7BgyczY1/7aTKWopiO
Iwszm7Vn+Crouqbz9FxqavjIF16U6qNWNB59Jar9owEzvm7CLbLnHTYkjrDu6laX
k0qS7IwFF+AcsjywccZAOEu7ArVLTmfDtMke8rHw3629Xnpd8DKAIdZYGVXXGOVw
P0bj2yx0lc51czZ9TIKGO6FZ7tHf3U1MbhMxnjs/0uennXjox666ParDmMBJAiq4
NTeFxtXaJUBoCvyNIIgnhzTKwIpPzPyftKM7LaTXHkLxQV6HUlcrHFkk3tDTMjbl
cXid0W4KKnRTdJk3Kng8gj7tpPqYKP6LufIdYKiCYgK+mmWx/yORjzatEniR1Jgy
kcTcW75fL0pZ5j0sdquGWMfZx9Ky0tLPltAESeljfxYYs5hX+KHhHMd8xXYv9qpD
cK3aD4tb8d8loRseY2Ixir0c6EgLdMtH3KSmoh0VHzygx4EIstBoJuji8hKEDLqQ
j/6q+VMCUfbuF5rJLRFJps5Zcr36mGSejmfJaqX6Pzy5pdWmMwvcfS2Vc9C6Q64z
2efeHMPv8CFD56oaSPVQ5F1XDl8a367N1dga5OVNbgKYw4m1lqvclL8+k6cTwyTn
k1zCS4Lq5TnzuEzrtUpeVE6eXuZowRTy0xAT9/udCSDw+zVm1e19hnqxZVspX/1m
BIm5VpYBaozbBjV3B6xA6f/5rMSRNfOh3E9+s2KS9hHiOQmi/d5AcIzKi5cBjj8j
+mkTjtefh9et5tItBmvv9lj1jslrs3IU3vPB7pzJd93RyRcWcgvxrJTqC9Vh1Ptr
IK0UBZj6d7dtQYHDUWyLzF4HqSGfkqcfg53lJcE0ZuLeN/70mG9QGRccz2Lg1Dfx
JL5bTHHQsrP3z9OXS0aJ4i6oSYhytVDGELwmHdnpDJZNbipaYCh11/aKObGCReTE
xRYKYKFRmOwehqEUZvoP/eRDlv6fJvWKSzPoxwvpzTcxnMyk8ZLVM6har5kQnGm/
zCUTX4uSlzRhIRm1rIis1JPGoMtPC29zhYB5yduTDLuMJnRz9tPD3qsHpTbU7ybr
oywogYyeLrtz+37Zf2MHO1YoZ8lAZuoOcb1jHYz14Kf2nvcby6O5Qxo/87LgbBDJ
/ujQCWZAgy2nS+B0MbORDKf4d3owW46S0oHq6+cKqe66AmD11aJ7pJC7uuJ7LmYD
L5RhZ84VBLK88rDoMcIoFmowyXpAqMo2dRsLlhCZ3TrYCOdGsUFvuKMTZA5xgwmc
BI0THO8Gt3zHKZPhlm4tXvIqQna3AIlznux9uZAr9XoIiA/5ktU2HdC/k9DIhNl2
WGDFg5YLNQKLiOh5oNCz+7u+lMVUpkBagMapCSUcZ4WVVfELR2orjFcuV2731WyP
dLaUl1MeSXjtj38DyxPjb2FdH5e2J8PbQ5dQdgfSsYzIF9s/Ea7RiO7IJaoea2HN
GILrfERyyRu+VCQ8+bbqj0tg1tCuboRAgHmBXHV5LrjU4NUqumnlJe7Ca9WY0Rkt
wyIJrXb7zpx7YSUdoW4fiIofQxqo8JNSTkrPV8g81ciCXrsGNez71coLGkMIefXb
1IlyJshtqWumMMl2tCQVbXk9sEcgZdihXZwoV9oSVutM9MyirPJ6jSoEqvkHfAxg
zz+rSU2x7hu8xNvqnihXNPM+b56b3JS0zqSOJ0QcLpzE4zN2YQn6ieFZFMGWKfo1
e0EzmgogNtD+myKqg67o5/DqAS18NKpApyWDVp1wH5gw0yeL9xG+LxGRApb9+wc6
dWA1+xMcHDGGIc1Bzsyl4NAbfsIrz51pZG8JAB9F6RtDrpte6c7Wyv1LTL+mlwW1
gstlgO6PBzuvtegC0ThFra+aub6pAR0paovdFL+UdRNg4CCmX6Txg7IIKyV27+ss
VGHr+JdW4WMzgIiFv3FGpdgnOW1KwyRh8LvyEHhbTG70CoyUydNnihmo5XboQOR3
3DehHsdhWt75dxr10B8nbO7I00P+Lxvfrk53sUEDotRe+/48yKaXA2AXtYP6XBzF
ChcSA4RsQa7Qttt1JqiJ/VZ9nWK8+ppkcu0atg/E5YScocUStGhHIWAvoy7MZilI
IIyCNUrkqwBCDpWlkuP5xkrfkmd2aoauyvz5xQ+EB/Ji7iCKVCNPjVkBOMHTLqq1
NQL7esBZnYPMsSIXwjTgbNayE0IpDiwLz1QI7CpPU/wC3ITITbkJexn3mlOzPdZz
gMXtQV8X3Q4nw+6/22Cje/jluKCjPGYMJm1duE4Sg/IVaBukh42Rn1g9dMDFW2PK
nOeaB8YJMi+0g8F43TRHUa+scUdj5o4YESpDoJ0c+RBfEtiw+iAfNOmWVn7yefGi
vB5bf3pItMLrQeXNn81/l6rLaBND1JeDI1glpkYdMe0JG6DgPSyYXRxSYe8O++SM
dVtP4Tj7IOFn0c7tN1pnOahK6OKKwqM57Z/ZH+Bftfr07NhOUi8T8dI8BYFBt/h/
KGgCkbwAzOnXsAKVVLQFAmDUOEnhYEBQ2Djh5XGPl9h6GGGHtaqRjPYdfQ0kdA8d
Wc4OnEyYJeAq3FsaWedjsSnaQGI2GCXlH+S33fjV7MlXIhL3/yKuZBjta9F3RJ+m
rs2TfVernHDiY16IRJnQ++1cHTqQyLIW1j6SIOV6N2unnSXi6US3Z8Wba0DfjhVU
HqGGpvNQGxWojzRjPqUy9MPFIj0dXzHdolHm0oXlhPx9O7+hiJueF3D11cSPMimF
OsH4tiDbypBV07mZT/SDyOVIeLvLT606jB5xggubG441lkjXhcL+yv4XHO1i60iw
dCV8B8ti4oGwjrf3rXzAg4lqjARJTkFvZ9OBOf3Mhhpp/Chho7e+xdui4ZNcyTdp
TuBLHvjIER5BYslYRXsn8So3kAtuyPv5gLjKry7yDRMMH02MxDStWbLBXaCN36W0
cd3rX/0g1E6TmyDMX7Rj3TKPoeyrXdL4h3xBKwnt26xIfpFOfbY7zUqAay+dZtCW
3HWP7lnEZQI1iCYTJVBc6lYlsOZ3ylKstYNjsIveJKQkHYwfr7hms9TuYmYorthB
DSH+R+Yaso+CRGJkOJd+y4Dsgx6dfsT0HHnGnOx84q/2r6nTDyCC06qpmm1ZcYn4
R1cpuLh7SizGkPH5KP0ZdzWlBGhLS/JtAfm4kRfYa/Ofgg6qNFf3mfqsd0sUbgP5
gTusCH2JpdG/gZ63qcbc/Ymqa4GbJXau7U5UZZh0Yb6gEjjIMRpsGnS1S0AsW7JM
Q4kcQoqdvyqaItJYrk7Bw5DSPu/shJMJKuMeKltVRMTWSNsc9NvBhp+xgqAN0OkY
pL4JKLtE216R72uNwcWWLLZKQ6bdQcEgiFBHkopVy1JZGHvBySnIK7Kj9n4p54FK
lQv/YrvC/8gLBUABMJWeXMfX5GNE83hD4YEKtEqN+pjptHUL5xM085O9CUD4GGqm
KjJpETkGdvePCM2c9tt0wttxGggw4/LkE3HZg760aY7dqJ4Rd7r2YKB1uiuga4uB
xnParhb8Xkb4Raop39QdsYZEqBYHHwKQ+i7nkJY2fB4xXdQy3MzSDNE36tlSMOv+
DXOHfNrdLBT5mSZVsB9H2BjYHmgiCHT53uYMY58TYc3gqcbP05lttN/FPPtlLR3j
OElTwHA3SeypYspZ//87tDqY1hiiUoslya7yv80mcTAKlq4MmlaOWQzppjx6sgG5
BIm1fbY19TuuiMs3nSlhjQh1ggY5c1+OJmM9GlUlmr9v73VPhd3eCaaTK9OopnkY
jyMpAfHgFV0h34lDlh8nimO32J6H4tREB6y+lz2yTlQx6gmJNoNUbtSJidJe+egI
u2qjyS6HtV9LTQ8V2acW3OH/eAxHOLu8zwMujAlqD5LQn6jwXbMUe1H17d/+0VXw
NV8yqeQDa9dh7+xaX/vLMONylAKmgZMdfFm2WLWtrNcktLcZ+YaP6Qw874ZWSyvy
gBu1IX30jUSw8Wg5GrDlAc8wSUaFUtGLSu/EujTasF/FUdJM5wExxyEzyY/rY+B1
2rVx1JWblizLQgNcy84t8kJ7a+DtwxJmVS8AP4ce5Ka2nxoa0p5Vw1/KePurBXXM
+w3Yp7y0314me+/eF96U3l86YwhkOxeUCWu4YPpZwAOtpGSRhEl/ARxH7QuWpPj9
snqdAAdTgZ/56D/1CsKjdrChYHCd2pj2bHEb/OhQdLtgUrLOFhFvO9o19IowjamI
tQRD6uV868YFkqJAc9qORI7b5QkUpFywtxUpCD7BTk9HrVG0GpK1wqZ8w9sQdGOA
dPghwVrMQF1DBQtDBolIt2vjRw+GZr4Ine1/6nq+K2C+q/yhpo9km5sjbZulU9zR
rZzS2hsk2gtjlf4woeVCM0kZnKeklSDKooYwCfpBrTepypJ4iUwxGVzN20sN6uyA
z7Xhu2O1mtPzL5gUNOlybEhg68dJKf5MrH6WFBaI1Zp7L4w8rMa/Ge/4NA/pZJBS
FsNazfhTIAUHJUfIJdzomsw+UPng46wuzrqh0vTKLmV0qLB5yhS3h1una5MuwiAj
z4WutvpWBbjgsbmyYvV235GTLU43RGclNp2IdJk4qzpaX0ugck1WQbh8jisKmR7F
EiFSXYve+Uog1rrbZtx5dKavvSX+/IEuhW1jGEL+5VFKq9cOpJlr643dky9OomRq
tacrTml2D2w06gKxr5kKH4zly9TOC1SrLyPZsecZQBEH5Wua+pnwLxgKN0Lw8opc
vuCbTXxDQpVXDy3oB3Qjo/oRk05WY7UovycwCAvCDLgkm+wIO7gSYGc41023xko+
u/5zqGQmVt94wxDGXGO4GfGUmcx8eimwnrZDUa45Qa3m8U0kjurOOvPmRhWOmn1V
F6u6Lzxk1hN3b3ruXMFxTWUSAhxYZNZc5TBACLsOsGihx8ql9DVDp03X85RRPRxl
8qhmUdT/ZeeTxm5ghfenH023p5LYtXgxUk1rtngMIPzqeIcFdncaSP8glmljmCEJ
DjgbwPtkqzdL8aSvMbqbhMFiz5+zB/GVuIIxRlCVqnHByzTZSSBRX9uoQBh0mUCv
XubNOpLbR5IaiJDm3raYsPp2SJE5YjmvlsldfhkIxyn31vxEGMBmImpehMwgcKek
atsBrZYkxRagqR8ZFv+n8SZLFoU8uuHZXfY6elr/eIW1wobE+VmKAkgK/jST6GLC
eE4HcD/hJMlm8b+kULsOr75Ycb+rN1LjjrcLFJU3F/NkNvKVr9XJ4VyAfUw4D6Nv
HbHwjFgnJv0Xo/COtMoB9X7fQJtKhUOGpi4sc6O0j9XAaOAQHRtkf0cjl1f15wdJ
ljgGcjVUHyxxBkqA6vg/I1ayOWLYKPrvQImjrhh2Mdzu5voXZzDmFmNYbyovQY5q
Zpp7TuVLaNlzITYuO0PxbuqoU8ZbYvU1S4OxdyLRLuSWav4bFRtvrbDdLTLTMlo6
I+a+5Fw9JyTyzIQvZimHbCZgfu/mzydAcLb+ja1yaY5ltM4PSV0uvkHCIS461IgT
oGbARwhNm02QuQ61EmkzWAro9q3Dl4Qm4F3NvymHxyatZuWLcGZ0PMzw5ijOGKJC
J5mwsV8SdwNXUiA4f5Bm7KN6V4r84LD4WRqH1TnYYp7aCnoAZtI7yZ+XfYO1EY8V
nL4UH/3CKbGH6Ri9uU01rRhMbZcO0FPF8p2mccq6fPXZAj/8N22IQ78K8fm8vhk2
/xLEivGbt1ovjFB8Ip6O+JQg/Scmj+C+pVa6moQ6ebCtDrd9u57Ox5Q4KXGvY809
6MY6HvnxqszAKgoSaSXscAgQIrXqPI/3YXHTCTpp76pRUnIKjTNJUGtFQH1/GF0Q
uQWM6qbZKaNJMt9VppXDkdeWbiJ502o1alZg2jkB4QQaEL3voQyiHbwgn91jaMws
mlIjVFhJ33bjBD8u3gpS7XZsSCVB+yzU+QYD6vKzwF3RkQ88S71p8nUoZsPuJ2k1
4u5P4gyaSBaFFY3k6OyFXGGCo0/eb9jiTIb7KaPDlvAvW/1QIdHBCEEW0HbIQzR3
d7Nz7iJt89bfSgwm+o5uzV7GPOqrGwHsZSd6CMQw0UgVbs7q9FNspe9hrb/vtKWs
HeNE3EYYTRQYbJjbq9AS2AHn0PaZYidXD8I1FCDMPYzl8n0HAQd/gDFy7J1tl+2X
VPykLKRTmjYksJeyxZV2+V8QKW+ERNZrmcJIyZ08fJ67tLy+2ru8fyeutVXAuggZ
QHQiK1nMsf348/ezWwjiceD0KbDQMS+NV6KoEj6NzpeLXu4TJP19a9z/lcvcbBbY
WhCVFLRQN+JLgRCvx3gUPCtSiTbeT61lOgtd3ndvc3+fIYUNk4RwmI31Sfzc3a64
VIGMqBP2J6T1GIk88T4DxTwyNyP2qhwLJwxU5o0NV8p47mDtnt/JdPTUGKzuroz8
5lOFY2JMFNfOYjazMVfxaXK/DfsNVA3W4bdGKBRKkJenheQRtQZ04hBXh1vOStzk
BR1gjgd6KIAsp0vDh3oCd2l2Qq6Sxan4EwfL5iFZVEqWsuwWC/tzHiHZ6YfBn/bc
+1rxAzLPjAThVCLJKYXxSn6Azc50v3S5rRxw7KmDI76OGEWolBSqpSznEAojtuka
+bUDVN80YK9N80w3VLO1VOLklTzKrJBjhJIPSZXeBlKYLXCWQ9njf73oYULsTkRB
lzZrOlSqvE7Z/TXfP6AOc6/m8djwRNojzk4MPGIRBMnFFoYLdJouhvu/xJTo50KJ
NxskbSkG5cCqhAoB/yCJdLkOJJ+0iJCUg9BOALn1wrJEqEheORsxcNxVDGdpQXej
WSTQJdeT3Xs9qynjxYbPAro7FWN/sQOFQFjSqb2fUXYDhNwyyaLECaNK9Eq5Re4g
6kkOml6q4+YdO18u9mYld2WH0PydAWHanfgv2opzrA5LckFRebvfIEmDW/83KB/2
yyGXQUQ3coV9OupEnx9/Maenhd82Sq8jtbv8qUFL2wGNoYe4cwMmOsllxOQf4QQb
ZuYjxFm/z4yOrku0MagOOsP7XO5gkC1RSPWNbv/J3f+oUjYhUK3YTzbfM/cRdgKw
jhVe+DOY/OCRN+4hHA0uHKbMGRdXB13nVttOik3xYVx1QkxGkDt5rwQusxxADnBL
5+8RBye2+4JMO4JN9lPh/nlxl+pr3hvG43s+ppxoqHAKznGIdOyMkiRrTIKg5T56
aRRs9DSosgcRoe3W+zCaB2spYHAXXtmGw8XVZY6Sck83CHtbh3Jq1NSi/byFxpRE
5ri9sBHE1szBwv+vw1EJr0/ivKVZMHUB67zVdnGHLpj60exrvTU+2js+Hy2CvSIB
cMgy+65z60YVa92Btxz3tF8R0Ns/ZZdmktGtua9DaQc1vYOfKfzKrUjRTt5T+e5x
gz6Ixl1Dv52LgWWBUWYDraxOFxvS3le/JiCzB+ouMza4DWBrJkkxZ93sAAw59avx
o6t7v5RG2CTawbG9+0x/GMZfF1QQht5cNgMFVelg+nUl6YpoKcDM/7/MGvgmqFPt
wRTct9ZudDa3r8L3MRp3lH2u2y8U2n5e0w2pKqLExZik/a/N8dJkiDoxPvGyComd
ofb4bNTc8zxRo7vKJWUxizmTu+vVrgcrnv8GZLURpGg/3aHQ5KsgtE4ULxSi+2J+
eSJpMHARaG2gZaGVYWThZm4aQRH3SV2COPc6S53t6lELJP8aS8EkpfRdiUpLjXk0
6F0RL1yJquKm3htCvqJv2SU8H/HWk6LWeXCMPUmxeQYzsb5kYsr5Y4l9fyWpKsXt
WhdOMfpUUyloGUByuRKl/vmiCzzZQrPBxUzj+ZqBwp0j2rqlPQPV7HyRcSGGd9Mz
nQe5Ui+zIp6GHsn+KhKLo/zHfCG/JJf1GL+PrmUAGJi2y5p6gXeeyIzBrHoDJBbI
v+t29rZSWHKc5PmUHg6uW7NHFpPKWOmM/CmYcGgda51REtKfJyjNjhX1Oi7h0FO+
IP94INfL/Q1+JLos5U5FwageI9ylv5lySOc7q41A3RDhG5WjR+pub6foVK6f/cgn
z8xfHDG85T0aq7i9NU1Lemh84QgiQgpOJQAYm6oxWWlodYPQZSlLtS3apWmBQyr2
jrNhCFaVtXk3Wqt7PoSVEdmEZW11/2+ZF6NqARijn6Qu+QHoHQTWc5rJaFzDGvs/
5zupvX4nlYVWZGrp5gnyNhCResRAjOITejEdSFwk4KQWpSwE3FVs16Zo97DbQI3W
Le94rlMdl52BJjaMCoeNiQvkkITtiVXdscqJ/s6LXvp03ZKK1xPLVxH/EI4XNIW8
xqU2cKa4t09aOKOOO+ex8OZzZ8T3QlXQqcn3xl3kgvYI9MreHfd+Ke8yoqcP4pL7
5mscaKNm+nETNk4xL0LVCBMpkZy8arVgOkU/6bcBLv1eVHc+6YY1qGTd+/VM3G3D
otpgjCToieeaF8upChosnctmZ7BY5zh05FYe1QtduXfJN99bkyUX6f+LbBBBx4xo
IDXuNTmwfspQZd6sFnp4Se3RiDO38aT6LXGUT3rVpQmy7nW1ck3/X++SYfBpnpu6
4IaPE1DZokmWf+H4uX1uJTW3kbFMpTDOnJzwqeleIe6qctyUYorQoD0DIpsudJAC
DUX374luE3pc12Z8MSQ51nzJS5McNN34ySNdHoLXkt8NwdXi5GQHVfKLnOwysyWM
kYTSMII7x9eTnEYK5F6S+ofKx6kw7kRn1A1yrwxMm1KXd1HGs2hr2E0cMNOyH0ZR
+Lciv9pIhpQM/hX4H1sD5+iSlgI5tW1aFrGzN8oAQbsa2xeq5wAQIJuTNPa2K0p1
otNrDmBcpoEgmt1TqPpmtcrR51JCt7pCryV6z2LJ/PT2gl7puQ1RFxJHiybQrM/J
+gYUVBhKxLhzPQteqPet0spqOoSWnB76jzZ1R/AtZSipghcu3a4IPxxnsIADRs84
TwyZHtFlLZzEqEB7Y5lWgK/ye1OBQneK9M0DxG4D5uwelNdBXa58f6RV7laFZ7Pk
JXN793Z2fi05mr4So74Sq4lKTiTygIJ+8jpjdjr717OXsfoPiKTZJzWp20ESn2Md
p1Vox4JW/4v3VUtzB0HwA3NGjnD9mFj6oWiPPMkp2C3vb7PBz1joZxecb7X7jdns
f5uq4Djg515IAgnGvWqmttVXqVD21Vc9g3FxYE74QLBMA06vmNxI+IK18v0YTDLl
zhx2ZohxNaAbngQQKsByeFqe4eAwHnZIcKqSfgTCYVsFQecJDqDOREyhGO/92wSK
qr6WA5TcXhLs9s9C752WZX9a6GwM0mG3OipB9P6yig23dpV3QENYvON6rRAcA/BO
Nxf5dlLLUr/GNdof8/4Wc7/qEJqKUCS3Qth+0w6aKR4pStNnQImTo1qDyj/yNyqS
228YedWj6DXRWopsYk+HmRRmi8i+MAMGOuSX+C0Kk/kdLIVC4P9mvFEFAjimrJ8d
ZrcIel+rAr+un8kzVs2W28QzRnUyoSzlbwggf4qTYOKaHQIA/+i4qQ68K1qrycg+
FD3XGCVjtG90qqevwGiWV7zLXAGFUoNFrFWFIXf3MqBDuu1Ue13sN45Kp01x0x1E
N4wjm70pWFd3BP5Wzu8OWirj7xA7YW6yaSY0gZE4Oaw8ZuH/nx9F5Kc5pAMiHkXb
ay/oX14v1vu9mwZDmEgg8eWbhsgDzUKV7hBx626NuraGmt4LnkhUFXkOvnmpasTm
7aoojgdLWaRarqLIli5wExrRENx44L8djZmU/8kQLlY3sW5EqjDb+PtdVlH945kp
wjZW3G+1httnjaYYxI6lWoNm3Hd/IcBo8rrpaZLK/MwTcS2oy8KkahE89WVH7p4s
vV4gLpyoyTzVVMZZzH+UHFW605NdmLSZ83m+9ywd6v2DlkazBoEaHSJsIOsNELYQ
w7W9/3CNpUo89v4kQ1gi8iNYRz6ApwiS5CvgRL0ujLJtAec4EU1ESGLpUAwNih9V
yg5h4QWI26e9iIAMN7inUv0eEFxZd3vHExYt3y/LUHaDx7opEpShEn5LFMw1V2Ov
jYTn2AlSIMO9LOWn73Yoo/ubT/vEU9lrNLxoyjlvu0rhyQj1VNFoQAUM/WZg17lg
4u38GNftYrOw9xi1rLYUKlvS3TlbQrikxVlhe6MqgS3d7+N+VdS0zbP8EbxClG2Z
+wgczToW63p4AhQTDjZakSUC2dL9bwBGWTnVwPsw4uv/OVkkK2FJvFq0AxAxYTZ4
EFWSPjCd7pSxEBgAHCqCxor4Df20ZMyZ9Z4xHzXrxdVw5zcZR5HAMbpiL8dE7Iji
UL/3pkfdHFJpjuRaYjnY75wbUcb7JDD6GOE0I1NIw2HG8fuhSw3wecjOE2knnK+j
TVBvVzRRJ0qnUAJ8FKSZQ0Ih7J0CDvgVYMwf7LUmNohnTec4DvKx6RYpvLGt0ze6
CchNQZblReHQvm4DaeW0WiQ0HUAQj8J8CyDbf/qnMWZzzDzO/J5+BVqXFOtSYBlP
gHijNCW0RbPGHKlLwHlHVoUbjrzf/l3uEjSfznIQx0XDACAvpwPfNVO15VgdqyZT
UK/7JUb6NVpvlYiqWBGKYwpJpUpJ5Pm4x26fvnjh3Vj5w+saPjJ/y2HFuBFhLtC1
CgbpFytYj7kPW7qC4wpZ2IdIlMxhIfezWztXgZ/dRhQRKPu/WLLEeRYuxPf0TBSH
jxidCSMRRb7xcN9g3oOABY3XfLiys3WXT/PTS/HGC0Zmk9xcWR3BKcu6vD4Ljiyl
9qoD2gV6wlbNjIbgv1XwmHDsw4Yena5QrEhXhiGe14c3pAXqA+IiMkmndCbhKOKU
0vMLb3nv8tXPv2uN8sqWTEQ0j8JuEDs4i47QKwiE5nybpduZtPxNbD5sa9bOheWi
Dz7VyxnndzBJCfSnzv5NGnB11W7TKRTsFT8bpQv86nFM78EX+5PW7adeaPS+1beR
2GUi6mzQtu65nZoCJR5a7Qb+pBc5lbDbPFABqrThz4HTVJ6UDL80aZQSH1dvCrNn
6NUQSWGlJZME6AsC4Ax5TzJmohvn19mH989uCK0yXreJdn7kzbaOH/k7q/z7tBQ2
wXvB8bKQ2D+8EzlpnbfPMXLhZjnM46mYwc5sOg/4uB8aODyRWjD/BjGTk4Jwzm5K
uh9kNNexz1TXwkNh9V481zUum8OOjMy6v8d97hjnH6UMHh0/I92XV2LJ6kgdhl6i
spWPeO9MYwivhqPaepWCRGuE4m6rIr71mjnrfyVW3ebv6VSKHSqKOf555DNq6ezv
m47Vavmr/5cZ+gYKgo+oYPA9HGo7UQjflMaSutjcpAlTTpUGbmZ6vm2mZP0va9Zw
WnvT7a6MB7JDGFhQvc262ZU1TItKdtXiktFIntVVsd0UFoBqeiURh2o1X6VpT+wW
LPdvAt6itpbQhcybrKiCVpElvJqW8o8r50eZ4w4OiXdhaL1GkwUYUGuxhC2jcvnQ
KipNqUhigpNo7sIJlsuiKeOiLpXWj5uxlEFEmvJuV2u7+S4eFUnG4Ho93CEhDCHD
swXRM1g2vUhNR6dzBPn5yXQSHvkEKiuqvPCQ+Qz4FzyHD2/Yv+WiEpUvBNSEePIr
DTJodXApZ79qmxLa4H5xHluLBQlpI5LVrJoLY/7SQLWVYzQ2/MMoKQudcwnKxCLc
FbADFBpaqRzYyIuQPJdryMFR/OCG2k6AgMJClfFLVT2gllatd2JfoYojV1Eh4SUO
7QMAalYIuhxaR3ny1l2oOXVPbyr6ZhDq3Z2h6c6Zlnbotif7DHh6dziTw4q3SkqA
Jii0puppWlpn6AA2b87NpDEggk1xZboM/lF9wQ1cDtVv48IFAW+bBTIk4eX5mQ36
a5cmY6s7ROwyVJNepDQs17ANBwVZwa1h49Ugf79Yha4IUx8tmD512NPI5Yf24ic3
z8OX1z9v3NZs1mGQCgAFKdKN3w4c2mDIAaSQOgxDADUfDxp2GCRpVNqRAvOn+pnI
btOh70bq5FGlw7jq6PGcQHb7irwRD8ckS+tml0YjWX5U/CEwWzhD3pkqQSwUS7j7
r6Hm00dRZhmYbWvr3szuVYCK81dW3x2SNBBWULCdSC+oQ6BhppSN1HYSrRrFr38G
3lLMeyHMuoEgSj7FQe1fb9FeFAYBUWt67e8OJ6IvXq7bEOryR6h5nnyPEKxQRxV0
XiR8dSfY76W5K3olfnNbt/NTlxaVt83OTlsPm0q+f2LaXpMuxuNocfVXnlwOBXeH
h9xCwofrmn4vZ/c5sTmy3MvKbehWqHTDfToiysRCDx3KOxaSHO79PCqCNkD4AZgJ
bkFTbPg61aRM3LFWPsIseJDn1RuNlm8KSzlMP1DLgUI4zqFfR+cXZMSqIMdTT5I+
aKzLQtchDZ4kN8VHDWGDnDOQUbZjQ14R3fdoHCNHH5yD2zdpd6jPAwOyofzcS1pX
3/CP5MfEOqy0/hIG7NJGY6Rbm44reHzaDirGJakxxPXQjS3h+2vFNahwwSnMsGbO
aDhgyFF8WTH1XLps2OPUZ54BKWzhONRUqvTPBHHvV0NT3/S7Mm0rgqU7hwA9LGeI
hSPt5MxZl/y57sJyFPCLJr/suDxplvQ0OFhB3ISZbfO1434UIGDBNVCOCX8y59lU
/eM/71F4lh0VPEVbdCfg9g2f9odlstBgGwc/cxKlsLT/MrnCAz/0w+HEvmv9sOQP
CPY8uN3d6ZCKsaBWmQesWsQAYw8hrcCltnexHPW6ipAYRRJwj5Wbp9yxwSPUsW69
jZecMKaZ1oYpv8pvEvOvmJrTJipXm1bqUCclVRwQbS02xP8cDAVkd2CTe4/ji1Rc
/j8lhFz2D5ruT31Y9+bAdWvOWYPd2+ibO6WY+ONs71kWvVEsO8fghvC8VDUxr+EZ
uLDG9CvNlUwfKjZ8powUdXrwyo/04wf25MSCYP+jtBU3zfHpKnQ/EJq5QSl6YD9v
ymJKzY+GgFe8/MmbB6BDygUlPmBnXfdKk89RxCXy4RvjyuTVQgyGhwWuqvvG6LwF
GeGB51fjjseQpjPkLGoLFeRX83BO54giaEkinbDvDjOgxQ18RK9eURgHU9ro0yld
G536bsTiVBS8kN/vmWEhDV0QXMCBHohtKSBziOO95xX49EFasCFMxYSU636XssGF
vfMa09kDxdpEewTc8pPiNHNoKMsh3hFWNjmhF+u1zWGg2YS0DNrdWBc4tSi5FP0/
CLB2cGJcXWOJe7V0l50lGujD4xc3OMsYA05f6vGLJ2ohsm5D0VNgw4pyZ8+A5Cnz
9DN4h0/AlTlfVxPB0ZUXgkBA26MCgxMpjHDtEuxtq/Q4KyP9LC9GTbqMPbLjx1TE
7yo5swsmwxUjIeybHy2ksceDtogwmP1+RYjcDXHDREC3QJ30s3xKeAgeFL7fCLFx
mo0+42RKxPce1da3m1CWvkof0X9LkpFbe4m+Pk9YcFnz9xgFD8oigS4Jf25siT4w
X2hWvtr6aBZhiKiNLpVsXou9rQnc1Fi/FJ6haei5CDzrB/Ka3wLwNyu8RPqUd+Oo
1l7zv2jEeL0cmGjJvjUSasRWPWWlJZLIReKCXsr2qGS6/ma533+DDgiF5617E5xT
sXFTxSGyW7DoysWEqO0aKfM0n8yaBU2bKKX3cze/hIJOkh5JRnR6G73HQL+fZDtH
uVXx0LG2L9hxFDLdzkyo202fL7eZRn3xcLLJrkX0YUljK5g1UtepSm9JFB60aRP5
i+5kOYVXXtL2RpFG08ICaPClQD/0SZJSs385iCadKkp3wDXwKQ1Bg5M1tetpmVvK
3yBDBAoVyH9loyNXKyn74VM+bEVI2Uf3f+5dIoDP7JxxZDM/eHFzY+KNTtgkyMrR
cZ0/I8KlSo+fVEeaPG81ema3vForWCqVMrzG18P4UOB1Ftn8x3asCprui82As7Dp
+DRNgMBY5tNYDCgq+AutF5F8xRxUBCtkvd6Az+z+9/BzzqPiAN8F9pZKk5sr93Q9
OwDm46XAhbGgcsULeWaweqbg1Ii0pWVBze0vusQdcG3b0x4RPvZ1xVYuki38Bgsg
cyyiBh5puKgeaIYf+BLI4eZwKKUOpQZ2nUFmkT0X9u+VIzlDqNTAKS8twWf2ptcN
Wwl8BLQLujDenvg3OiECpjIpQIxsT6eIVI0UHpgNkBcDURl9glmwzVquSXGuFJpW
RCKkNW1DBF58VOacneemp7PWSb+5EcV1vD8fgs40zbB4eb2gbPTYIGwCWmszVvJb
Agsplec9GBL760EbexsUgi8Yg2TKx/FElGTNKX76nbznHy3B4N/9MxI5QzgHmUPl
7zcEgpw1Z9TUtpjCT3hAweY6/2IYfQZjhf5kj8SXHDALcoG3DlKvw9EQioMvpfFt
e0pikwV3NByJex+yuCAJ2nlTCZjdAXJPTBPdJom49+BiACPL2Hzgtsban/ziN3CK
QFpkMqLxFrZ9cPxcxeYQeS/xr8PaRUgJPRvrnCAR/K5lhDcjuqMpSqH6EhRv23Uf
xOLPeudluh2+sPafo2BtCfloprpqk4VnTJ7wFOpVWpF1gsliLIar92Rw5UcctKY7
5912aybVYGpNV4BfjYIigyL2UVcM/1Li9lPHfmc20y7FNiXU6m+nnMeeusUypPt7
VGp+mj0pltQm9Ryl3DQ89Ba4LXViwgptdKgId9Q4vH0kONrP3IG9LkSR9SNxzD2J
ed5fH1Tb0IQqDrbr6UMSpHySvqQIZayi2IdYAY5/d2Zf4jHqVfUqHjmnAe7vs5gV
a9NgmK4jkE0+V/ykgC36pkWA5trSix3xhtqEZwVje8VkXqWyt/d0HxMqKb2c7vQe
ZF8Gsy8bmjmvVesRVCnp/0rbu+u1JuLcKL47C/g73OOxRqGncUuTprqslxyPKpyf
rkd9PNM4hG9FWnJXDLILjeDOARXspAldvzgm+dKjjzL+Ti2YGo7LCStmHgePscO+
wQNQs1evx0w7RWnXp6aKwIKuz5luR1gXKoqY0yOw5EUy5TbKECk3szOBQBqTdHJH
sVd6SVbMOaaSvxShTdA1U8l0/M7N31GALe6Hp8of5FzpPdd5W9hdBL+gr16DyC+/
ys1wzPXSnEyY9EcGZzU49iv06TmD08v3GPejHJCd+8MKirSIoFg2HxMeEartmbny
0navQbiF03xuKpd3sR1kaPd6ZSxC8CX+BD9mYGf1ShartjlCP7L7bUs/OV5MOhEd
DkK9N68pJ7gAq6DvcIiZ+Pzko2Eg2S8AseQPEgczFyB+gFdaAoZt0qbfZ79T8p5/
zI9jvKhOP+uM1zM0z+nDdvN06t+VYsL0/U9hQ2qYjOAi/yR+O2tQQKsAc3TQTux6
V22DEXJozVWxL51lcCg2KiVPx7eFyBYS9nq7x+OG4P5L/jf8q1u59R8jPchu901Z
OccCHocBrSiQ8lQ/gPapPRfxtFC3V36vQtwYyKkiMrqGFNfefDzTMP/nCiikLQC7
FMC/nv8vc/m2Zc3CBKXrkn3e+dW3FHSN8TBUjL7FutQLVE37XEskQHBEe1PjR+7G
et+8nv8u9CxU8Wsk1Zxx9fG7+W9u8YI4qtoKe3OVYbZFTgqmH74fmH8TYaq+K20M
Q/5Z88sCDTHB6Q3+2UD3I8dnATA673VDsC1roCd3FoDG/f1Ze1ffyykuM5CC7Svh
/Fn6ggUeuSPpzsfzej4S4tbys3rD7zvFBkqT5An63gP6BrEMn0MWLBiuQjzmjcZr
CcUn47qQ9cRWzyF7y+i60A79k97epPVXjIlJeyn0+TU0I/naqILxsZGwbEML2zhZ
79TkzPmjCOQguMGhYg2I4eShlDdDen9FQYXJII8d2xhT2QGYQeZ4wFXdAKqF7C5p
YA1CsvMuivoGXJYASiBGI+NBMMdCtr9Ssk4DHbHto4N/Jpm+5tdJxxZaFbVPvFRx
/XZz5zqkvJX6IsNp1PDFV25y8qZrAqnifAIUnUIHAaxyA7k0ssdohCcyjJLU1agd
fAG/L0W4XuCOJepRqw0ntuTdihTmP4iaOXeW4jrpgrR/H0bN9ePIpsWNf5n3MZX6
K0z3FLcPhBQtcbKWGKmphnD1GVAMCvXNJT93/MX1kQmVAmS8zLwSYEjI2WL5vuL3
x8k59iN1upxPCu8Dtig0d925tuzlS5hDTGir1oPnsrRzJzTVb8+NIkk4eFLHKCPV
K7fTRQ7PKWzjpL8jmtTFIfq0GwNebBdRRBYcyiocwcACR3ni0DiXNjHyFSuZGb4e
HYt0DCWLinJhhjrk67TOGWNcYvOGzpJPL7ZAoQwcVTjwL0jkLtSs+yQjaebRzBDQ
1710NxNWEAyK5/4SaeDIsvd3uxQ4aAWVKcDTMQOeiA5ZrqXAxKWo/s1MEsT2lQ5r
I1pak3JieIn8aKJGKMRx/oJRo1oRlAau5sA0PNulmq9amJ63p1Ox+tpawSwXE1+3
uSh14x4k3PBomWDstPYjBteehuGMEtcnFamZFbhw3g7kjrbjiwP8NlXlqXaaeK/4
kBmO0oA21X8uc5IExauZV4L2OUEqPsOxRJHf5UBKrfOv2Dynq3mZsi9vgaaD5UWI
ioi0k34LBVe503Bz3IIbw+iY0ocdduSXCnPBWK0cCSUknVs3waE1UUucw3GiJz4C
wUDNN0tPE3uAT0R1cPU2kzTvpt43pABBSgHCEFYeduMj2lR5u/cVOydhWH1Jus/q
wCgMZTx3HlBvLYBIU37WEO5pei/3ymPbwMEqA768sC2tvFwgMhQIAnl+nlryRAG4
cRMcoCrUo+gmUJRw/I3y4nz+GnAmhmb51xISYRlOfw/XP9+jWypabvkeeiM69oRn
ahBEcSTPXRhILv7kCMw8oh8n/sN2NdcyXH3YrmusekMt5oyghU/QRARWdz0Wxj8b
0hdgagjZRoXnc+68CbzYfdKrpTkL/UTs3AGBgfEEGPeRSnnyT/FB2pR01cXXOxQd
htktc+RwddIL2Q5Tln0KDUPfKsYfof6Y7tXbIccmtFdbRASLwgzBq7AT/WHbaYrX
4MiuytEvRyHoyY2sv2O0yHUS+mFpJqIrrh5izYR/HmPOf6bRTeaqfe/q3auTEhj1
UpgZxb5tfpH1Jd5Pn4LG/uCXJ+5Y9/0ZEUSGKO9GcinyXmp1Desk5NG4D2vLKsm+
z7fOZu8XFBFwdGlER47mUNZCl+7gWcq/1qxsBSREwYzmUbK/FojOWV/Yl2XKBvfm
Z1N0Qn7xx3jKgGpTfroJ79Xjo4meq1WPQGDE2+DognBFB17cUzpbqWJfBvHr1Ei7
E6Vb/4ucPeLqbV0CjUVq+bZNGwKJa5V0/dT1rZb8gJrL5kRfTVgj72ZcdmY8g9Q+
4Tn/gDINKPVela2Ov3wE48oVP8mFo1W63hgouCxoBbTy+8c7Nm9i2i/Riyud0F9I
bKiwMJ6F8CqkKDlfhZGLesMd+W1GLodbNftLn3zMfxesyuu/C10JTiiH+HybY9Xo
nFsHWk1C3uzAtan0acZ+75US5PeOFMmhKBfD5MHEaXLKh8GulfX5xYXNQD/WZui9
VwfJJHoBd+4cONt9n1qmL4kGevQ34JaUvM2OWJSFtU33HgoYHZYDqbQ8GtWPcgaQ
lkqhmU9+Uwm+VG3SJNGqFRts8lru66nxHk8YcnfUPZM3dHy+iZU+uGY3tqcBOxA6
10s5PFXShZoKV6kNNhN8A73Y1tXwOk+7ghgxkWA6yP+uVNIRH4NcvmcXXtJJvwdn
EYLZP8aj7UtETgu/vcSt1r7NwXX7j0QtPN+QYuPLR2EnicjsDZG/Mv9+YlLTUeuq
MUVgmIJoMsTI1exL3768iDeTV/5mKLCdromq9yAHyFQnx3Ci3iJg92uSHPxDgeAv
T0e6nJyN9+gJOwNIsUZ6q0v90ZBZPyre87XW94FKcrA5cVS7ElfID2U9JV+hZ1/b
Ckj8Oyz5BlJ+qgYqlDSIzX2D50o0jT7mAY10MqOlEB0EVNqtFXdVvK5xY/3d8mxR
pW4B1MrFrJXT0oatqqUXvNEZS14ROgNI60k18yKC8XBH1kxzIYe7rUC/xDRaxD4P
3b8Uh28VpfoItwX9JuHJsyUGCdUU8BUFJyk0nHHPlad+qFvLHMqFA9jIik/9/FZn
2phrOgY6boEGLzCVB14aviKNX/8l7o4plxng1f0b33qVkHwz5+NlneOO1jGS+xXN
ZlY5G09LGNAyiNuZzw/u0jcYFAnBxCMdwcmCWC/XqqkYY/TA9fea8uXcQTSbnE6S
mhqRbERsumfPKjVQ5OOlf45a9PcedgF9YMJ1RNhNsSsNB+XLKFl0aTPWkcUCEXQ/
QHryA5aLIWJKQEMqpf15hq3ipthxoX86wWpKP5RcIvb8qaVtGLWOQnC53sfJiap/
TIUt+vVFg9iWMjpDvBK3LwCdjK0dBCa82N0q8RgplBLpn0DiEH/UTZfkW4r7TR9S
kReYCgsNIfOId7zuHN+cv8nJNB+mpU9rXtizfGOfkrwu4cV+HKCpoAEqYQcjjgH1
fPbd79Ntd6SkBQbKSYGs0F7qjvxD3rFJS5QjwC2o6NTjZuxO99dlOKroRFUHFSRy
4A1jnH2z2Kex9Hj9y1vrCc9wW5YPjhJ9ggWaPIwHKG0HhImzYakA73h2tFd6NJzg
fwppfZCAo9xG74ktzh03EYCHifU5xRwIkhpVbrultbB3JbhzBsohs4GBB2gN/hby
AyR7dkXTvhfhLfcIVzMupgoioeOexG4b1N9oPWUZzKHgT5N55qhZ6k5PIllVEU96
8Mj/jYKPZEMmZPomtKd1X00SXiP0QgwfBiWctINlS6OOv4ER4GBfC+HSmBdelZu1
UnzyFcHU2HFCgPZjqjqynca7VRweW5ddC0Nz3NETXThZrViMo3x1OcPs9p+SDYn7
FtlEWpfYsBXaedl/f3XS6z7Kbu0IGDPYKs/SJD8DmgB5dsnlwsHj4RBm21vHkQ7b
xijPajsMsemSEAsCXenQdT3uSyqZJhCY+/U69H/b+Az/6G8fgYRe1qkZrgzt3KED
RSZy3GQgseUKgTfUCz22+U8TJAvmCrkxCN94T++qEWHMHrb9Ffs+LdybHYKRRuTn
FLpph9BWeKS6U2Tl12Wae6GAryJd4QtjlkFRDvGHMF0S2eIs6Pd34btONuh2//Tc
Uy9WI0pAQ5KFzf50xWG9LFZqi96Usn7vAF7vmYSH154kijX1r6eTdapkkiI8Syr2
IvRqcoCbHrVTVypZP5PwEkAAyo7DWnS8/1ppzQus52szjGjIzGn8Kmy/w9hjPqxM
ACXAroW7SLMD3cm1TQVlxS5xYGNxIrsszOdHnae7PMOIBJo4+Z5Zr6dT1KRzs1D0
tXOGk1qydg1b3q7O5/ud1EdqcpJ3aZErJyEE5QgJLE2PucPmfIq9GIyCmTlv4B6l
0V4A7KUNoP3REsWDYv/Qq039REp1xs6IjluBjP0Ksgpy668wDsrkSQSPdJbQqd1g
d020oeflp7FRRtd7l7YO7NnefaNKTtDzJNTfWvu9VBoi1mHkRskpoL3h/tx3L9we
WYP1WahKLaD8KmqUnqRFLb9o5pOxgrMlNgxcuMtXIVV4Ec8teSPqhdMZ5cw1X3Y4
Gc28gjqaisiRsJ/D5zjSKY57PpQMsJvJ7fUYl96htV0ATjxISovuGkpdBUONNce+
a4uDg7F6DZU2jfthR5CqZbYBIKqJ0o0wEnQZfigRtHUwb13C7uazXniqaBY8pxRa
ffWEwLHB41iidvuOetZ7b6MNsxukFHxQgAuJzra9zVZID/C0hmOZK1Ot/XFzYoMV
HiB5Md/pV45SE2g+cL8Iv5NTZNUMkhQ24KlZc74ui6Cygnfn+RGkQoKYA5xkdxrb
k9gTOAABXouquy34dPpxVyPZ57WCf/wDsAMn7BpUSaECkJQSTCEDbjC/MHoqCwMA
G6yZqYOZkXPmg3ek/LbGSno4z1n8LwaYkfb0lcWQyD0sdjFVrn82NiV6jg5OnJgK
2E3+u69xb6w0Nl/sJDeoLwvMMCdZJQCOrhKpKBP2IN2lz6SRallxlpVtRNhEkn1R
QitA7uLMAIjclWI/u0O4ZV4tY3Lfcsahc+AmdKciZRvyL8BS9jqBy9bsjmrbz7Ko
4Idg44hriSm2/x71MPI/CmEaZDJanusEYFSICaqkAVvU5mzs8EPpQ/R727OXcjFU
tUMrKKP4KVPq4Uq3crp5rpI8bSdKEyhwDqbeJdYtZmo7OB7XXmmEp58GWM99R3Qz
TROVlxa4jKbD/BW9nMVE+YNWc73Wbfo5lopGndOKoxrXJ4HfLDAkN0YQo4NRVqrU
FADBxr9NGyuFZGhUqous7E5LiGMLnE5ZDSEZiGrECIRVBboOW2BEyr96gDVxy58C
Ons4dQ186N1WCzSvYp/Ecwu1rE2n4IRQPBfeIMxZHKkXPHLKybg3KyAJpHl+kKcR
YDVqaInnU9lFai3BC1DRDl/DzD7/BoVAmQ7OhPC2dVdTL9Q8uROzDYMvDsX4yVrn
8wIoLfln8KwAD7QvThjja6v49QZZqp0q72QmwMCfh6lnTz4BILfKmbzLQjY4FadC
EBLHCTFkXx42ZDuS/LFCpvlw+/6JG5fn992SKbESe1OoJWlNlMPacmI8e1A9WpPY
G4qQsbH7y080mXeE7iFjRb1lcL90FkBbJrc/hgh+QKGg30Xna3rj1JTI18n9Qkra
/DUnSHNauJvyeeXavtN2Lkkd/75AtQeQ7nOkgdcA1vbsm9KVzKJAJIgjOd/wI+IR
eHV87kdst9tIFS6I0K22Txl5XaDKu7EAvOQdbTuta69qB1Hku9AON4a7SSdEdlzc
eFTM185kMP1Wrd68AdEKrlr+bKhxqV/pBUF/97+n/m0K46/s+vPD8Vsi8hElgu5X
/QTccxNnPhxVS/4XNuNGPS2r4//lGe0DOxoJjmULUqXUiXTeJANaRZexeLrtYs8t
LRwkfHQL+1zzIMZZM4AhZ4RYgXg95M5jkjVKKsuq0/kBMnQUhiFohkjd2EoxJJs+
E0WehOOh9cLFDFCVKZ4zvHnEolkNmsY4RMXnafUU7TwBSqaJFBrou2IbSq2KZ2lj
iVM6D2i6B1FCgcdCqRCMVCGmbob3dzYG9+2nyKfs3xGYNoo/t2R3s+EROhv4xiGL
YEJPjNlBRgyeXaSu5UWPSG84ckVum4zdDB94xLzdA81h4xDxepQrlTKP4y67vBA4
9F9QjAeZiFZ2wUeg3c7EEgZZJ6hN5GjW0xAa3PqsXXiFPhh2FcCwWWi0X4FXtqOI
5zA8NVCrLINlSxr1Myz+lI3D/fYhxNDk2090btD5K37AF9ASz/j5ba6vB/m5un+b
AzbVnsTh2DAvjloiw4quvEYc1MZZF/SYFjV/DhRL4HxM3WpIX83dcw4wFPQbrfcW
1XpZJvlGYsrMLfa7+Y34i1RHe2tIbKSijI61ze/l3uwnbSSD1F0IvGM15zDVlQNY
6w8cr8E21K9R/ZoakMTS7G/qbcWDuwFRNv8awR9Ycu8+MOOfZoeqBURBHQc8wIFn
qTpYLC0+4tnyBd7SrpS8IiQJDoToXB+yOZcON8cbsfki3sSIKKEJU7Tm7a8N1TdI
liSO2QIh0xqNLhkMdAO5JygSVu9G7vp4gIK0HshzShRQMAhrjWNfPCSIcvlc4Qhs
KUYXDmYJWqCGSDpYHI9Y54SPhuPZdtnQpj+PE4X5sYnP//cIOjJHJpw1Lf4aFyEh
GBJD7bdrnEu25ckTcM2WO52bJvbqzKj8XoQoRrJcbo/IclPgIeYTYM4lFGpvXVhr
63+AxkdmSUGjIIxe6mtOCBqIEFlSkHqU3vfu9hr8jcBWnzcP7X/H03XMRMB2UH9U
h6UE+rpp6TbPwXH2cLDE5f2UEIOJVuPYoZiEhPApCr+jCvRF4sotvCrCt9TOywjo
KfXoRpw1OsvhElDYDBULn5JPnzgWHJhbRyv/s+uwrDKutfZDUxZyp61/x8jbPmuB
ViQ6WZOsBlgCKfCUNEL+6YDAGBoW26NZsI0EVb4SYelo5SZ+jVIwBaEID15vSN15
yiRt4/9kkFQgfUBjIwYfsNoffgsJYCqpYG6eGI+j9G6G4U+cEiPl9voI1IuIDC9t
7xgVcyk/n6VskKpbKAcafB7e7fr5aKgPgS2koTJ+eDT5YldGFEQ7r+J8DhRGRl88
qcNhGsmRz6q2tGfhcBaaSGTzE+oyGIM7ZO9zJD8izmVWSkRl1RKwOGEkBSJFg6yw
pzXpeyTi9i5qOAPBSxJsf7l+PY+fCF1hzB7+H+Ox4sd4PXm1FfWJEEnnmvqkgxwA
jrZMB3e9pC4PZpNa7As9YgVhX0FOzsfLXVzPLhpCX19wvexAOdQXqpd80zBk57dt
YgWT9fikgThpsP4HUyyQffrptZxqxAFSf7f7oieQffzCUQHupAlAIaka8O1u4HrA
w2voVfRqz9N5HyJU7z+W8B4MwzDDFbIWc/W5t2RCWQXCuZKgwKxBMVx/zsUemHD4
E71uH8LtB+g4IVxxE7Da9HXBskekLmP/xUddOMPoymkS78ooDcC6aWKXTlGvsHCK
SByG4eiwCN0CXiCB30raaoA/UO6dGvDH78FFMUu2UYsU/+qKpxuJzhUZBhaZGmmQ
kxHLP4mbhNDap6Zmg0yuL2bsKGM9sJxxfbGnsXLaS1t08ljvXsLPJqF49kxpWzXF
8+3e3oKGmqh3MK2w74HOoJphoHY9XUM5XzwR2pIae57A9PebIbTPAY0GoYPBcpJF
qjPK3XrNxsrR1kcXO8QATFu24mJJNp33w4pD1LrxJIphqpj070/Vej72jjaAAdLQ
ZEJcNJoafDxD0wNWwXIZOyBASqQSKG+fM31qBYoYaaxrk4F+vqRCuKkXnI3XJIsD
9UVuyK034RjdIatxVcmxQBkwVC0m0unDMnVonAn9XoFppDdyd31oUCx2gtfiBfCv
zA/Q7yI3WZXiXhcy5L6RwSBjzFd7fJICprJm1o8v13vETV3A5ZcWSKC1XP4LK6LT
AmKHzMcezZnUVWhMjde8nYJkBHtKCclHdU55B60kJT6a0K4jU0ERvWb9Y1Zs3Dk5
dD3Zg66nAGYZ4lYCsdHyYth46h6bWQttW7BCpP6O/QBBj+yVGQ0nnaFc44Yr4RQ2
h0YuZrBCkFRCVg8KZpXHyvV5mfXlCUCZqCYepy5KHesT9mt5J9dwZMqvFTj15Fem
hjW25NRTvZAkC0enciC7+0v8sC9bbJZayfdxK9vh8505oiVsHQvT9RYm20hAWu6C
xQuPr7ZDgu1bHdku7XKs1h6XbGg6oEMcwE+YBTttj3EVLGcEETqM2TarDyeFOMZu
oxqO+Qh8lmSKwcVk2VIWmEim7+GiQWB3SntrhZ42UmIQt2VvvVYRmUEnbFIaPsOH
V/TDKmeiYO3C8WwasDU6RYySZBynb5qramEMlYh0ELLTAp1Cf0Uk7G9y+AbilfdE
bNCMZb56V4tuYsuoZOfoM3+hUXdW6Qk0d3aZ+oUbpLuOE67QcwEfoOyWCcYJLXYs
xg3M7AzSE/KbNpwB8U2Gk/kALfEjn+aJGWLbLznNANqgxVYmMQtY1AB0t2Dub5KH
F+qBktWNFi3DSKF78K6LI3kQPFzvlptMDOs5DC4qeYmWUPjeoL9Pf227L0ZGDHWV
sWcSgcSqZ4ZXnFISqal+WPAFSQq+Z4aFE599UapynpkUeGfKUHZ7RIBuhDTMDnt1
nAQhMhAgpqys8WvYX/wZC/G8n+3U7YR1g3EPL6NE7nBGZoWrQmwNB2Xvhzi+z/SK
2Tx9Lw4e5SYCpHu/wjAaH5g6qVfDkuuhHhr999ZV5TJTltU31LlY5d6BDh6l5Cj9
Cvdh/u7SWP41EzSu5AhTLELLhjpkME3P2bxynh8KAzLBktWDGxBeOxMzTWvrsQI8
CWOQPFnTe5qheak5igpdcKTICzd6X/Ll/2Ef1FMJDPKx9x+8uOvwb4AaoFzABg8+
8jT7qihKu0YEzbu8P1JIHha0F/m7FO0dBtlYGlBrSoZpV+tVSVUY6JQs9FM/3Qcu
m/gsQP/2O/0yMEIJcL0Sp5d+6NhKqqc43qP8Bv219pP4+DoTjlPiMc3mdLlHD/gT
W92wyoA9pM6Xe3sA7tPzkiuvm+yYTVfGYRwT2kgvCRn4gWiXvOFJYqD3HlkhoVTv
4I4Tuc+m3s5pFiKUN2j/HuTsK2jmnZfDTS9tDag03ry3346OE/W26NWBzwqpDPDO
2ph5BvHo9bpX/TY3ryq6Q8XVEqxinA7y4JVLCW2/SEdcqcOVOFJcMGAtmxb8hH7A
88+Se/ZBTqPLcY5hoDjSRc+gagILGlPmWsH9+5XUGzxUs8yldVqaoNMT9YXJm3EB
NdDGEywSqM6Mjv1F3NRdz3e5qowy79DznmgGNle17y/CE8bqVe+aR3VBF8p4X3/S
8kAQja4/fWtMyGcpe/uaIQfchNuVmyVii2f8yV5fsNHwMn3pWNuNVNPDXcfECXeP
13CwIfHlO7slNk2S9OLFmv2KPzcQ9ojtjvI29d9uPE8CiTMHp9rlOJ6CeNEs5MPe
RUB5xLVB7Tpj5+ENRl6qcIxy3CSrFYJKqj6+gvZikMTeenyDyI261VH8wCLH9fxI
0WiniRrH4Jp7HlYca2GbO1dgXP9gwQ7sbKA3B0l22QRHQ793UrH8ky1w10LSItZA
S/F93crrOoZrERqoj2Lrz3jpTfhxBkk1//x0TIHetMHc7f9eBRVyl+MTZKs+Y0VN
UH5he0S+0WeVjWj+iUfhE7ZlNPjJsZYOx+aC5xzv15wQopHDbVSokNWpdBPRr2Wv
isfN6IfWZfIlfkMHX6Y/a6T7VopKENNqZmTj1SM3oBe8nB/JniuxfUa9G6vVw+8o
IY91b3Bf8WQ25jWdbfXWM9dpT/EPRjMOMD27by6LS8EqUMJGafVD1xEzNIM5001E
eJ4mJYRZQGDe1GMvwI+PtBJ5eT78XI9KJIHtPFCtMM2DqANdNC+BT4WKF6nCRREU
jiR7MmipEG61SZwQ3TAkprnW83t5cs4tW+CST++5YGFLVB7rU5NFyd3JZX9xipHU
vRHhbi78n8kuaC43ZAe8OVCSf67KadtuK7WbkryLodCaabUMbhjS/bw/FsDtFFpQ
RdIuWYtYMIYl33KHOY4CAoBLxE4yk6qqjWjNhWvcgi7mvZKXhkYAovtBD3STPEpo
9O1TCQPXMHD93mkElThqlWwoblbhLQ9Ya5s3+wBtX3lHJwcd3arXyYS/2BIiRgPS
m6ihAjc5O9qNhCeaTKt8xpvp73+lw9YpqgxLrurzVhwRvkXqMCAK7fVOMLW4JxVE
3FukIxl23SbwIfqPekvTgz11lYPuxrBh6X1vsmELO9Nm7ZSj2IrREdvHVQlFIvhf
tBA3vbtlIpQ4fm3clGr3e351SU8/ohg/H1sqxG5vtVCuLUxSdbk5QjseohMfKA+y
kpgaXOUmlA6t0mwqOKnLPFWJGtzSy4yor6gEONXwjMtfXo02eGRO3Ki/CrRogxqs
MZ2xm8E4zcdiBW4IqfHFPnuRCAqtbtW0eaTpwBMTY7uHBC4Z/IuQRYAfsMTK+pYq
3S7gXtq4eViEgzgXXAj79PCls4ygmAZKsxsRNePd3SKrkeiz6FL8RRNrkFI4pLQW
iWw4FdQ1qWp4eepAIB35MbSJ0t84juyitlnSJ66FD37O/EzKx9avaUJsu+wtrUGw
j3VjnolfLOuUEvVqFHLNuF0f6hHhpcGsI/wTLh6OoYGKVucm7M4rlGAYDTNuXpeN
7omp66W4/SjeN/FgBAgX5/4zf0tKE8Mchjm/WI2nvFYjDRVQkcCEIisuVXWco1eq
Ff3aXH/iAqzVFGqPXZQ1TZrScEPaJaU/SCKQ5GtlwU9rCYRIdCxsQippAmYysDXa
rPufwcc0pRQs6XRL0ejOxSXjW0jpsZw/9p2Jv/wDcOISfHc2lHB22w+BiOjlc2En
lrflqqkYWv5GcM6cDPNnuqFXOxaXviH6dnoRs1KNKVG753MrHaWDJYjVs/OJrxq6
MASV1+VPQFzWvRF7Au7kpMGwYGe0UzaX27vE94vXUuzrE6hCByhB2Ylbt2bBQEfD
5rrUmQbNWWtZ3382Pc17tE3Pk+4ys+AEwOsUxfT/0pXUxx5IY63i4MOBX2Ir9HZw
TF5vi3wu//Cv/hHBvSL9Rhd4aa30V4jxeuO0spqHkoq2GOwFIzrNnz8meNz357UG
Me7idhaDj7Z/auCziI8oINDjecHdRZCFNzLwvkAfPowuzyxDNK2+9OBsGPtSvL5g
5+voeuDq4rGJaEdOO889iBdu8iGKCCltH2hpFm1SgxGUw+agIvUzc8gjREd60YBv
GSkmGJorCxEC5xFTAGXGK1iWHd8jWXHZuQYH/zB31hItVLIOBjMcJyC4Vce5xXa+
vnuUS+X+A/YigMv/a0z43e+HHvbkkW1SlBvdpAuCFa3FEvC/HMcsYq+Vk+bwwtO2
oo2XbWwCr7tuT10YyL4ML58URHfg8KCiTUv2C98a6TXhtSKjmjvOzaMsanKWnxn8
Kdc35jDDLZWPE8laKmiwOQpXPyI+Geb2vfmaS/skkijvUBFaPcXBzVPgCdmDQ628
0U5jkUOukOqgk/gdCDTfOycxiHcnNgWXVQGVO9y2LefVGYBW77tOJTY61wGWhOF2
jK3fjW+fWXYHUFhG/Kchh2p51WMC+A9DAVVFS+8kh7tl+OGiFh3cJADu5iO4Syq5
SYNMZZevf3oNGM8mtQlQHpuMVIeiSzLwYVhURFMwvwDvXFZ6snapS19DidLamzpu
ElsFUybv3pz5uHYN0rl06YAPMpRTzHvu2EvACC0k9D82XENGKl9KdBNnSA0auaGm
cdUDfH5Qz+Dszz1TFFOYx6kkMmMwsdNQtcKhHy7vsdR0kXDMNrlXi4/pTR2pqnsZ
Z9+N5nj65/EzX3haIqSvw3P6IrltkjIDfmMUrEI6wRs/EMQsrKalm28WlAz2wmui
k1n48z/+zGtaC2Aftas+e1zI3CVFTpBAjW8AEAZ7GgSLO6N5shaECt9W3jyHOyyZ
j8/FPJsKmIsSiSVeX0MIBt8s13coWkIIwigjRY55p6OOsNF4Hl+7bUTzpr419ZpM
lpArM6Zx9hRxQcjlY8O85PeTacxa/Ylk/5Ep7t2lwuOFvMozhsn3tqZFPUGGGhfM
5K5mWjj0gst9v2fgBnMC3cN9yHnZiMJOxeysA/fJkFac65ILpjHeEyMUixD/3n6U
O5iDeuUNbL80WhkFJzm6KjRtQ1o6EQtEKlfMA0AB8lBXNmgC0TAz72yycQ8kc2uw
SgBm4NxWr5pwaOY/eKdovxoOnTjQISeUkjoj25hDbN7hNqJx30T2vwDElhMU0GGn
I2VkObk+Lg0BHpvN4EDLbf7KcaVsfraSR6YpACDoEKQz7GbHDzTOKjBtSRH4hEzP
Jd043fRn1cUVN+PyZo+B+CDOl6Fwo3+Yr8gI1PwOxSOEYlqxnxpgWEWsI91LsUSD
8dMY54vKMPlHhWaBNx2QTHjOUewhSwyu2ukCH8tNSXowVjGJ5u/Ay2kOhaArAs24
8s2UlHwj5biGn9Wa256NadLd/t0I8mrqRO2NMB/MoMdVLU9IjqZ+Iwg5+Fd8RjRf
BbpaFYQ65p9q9YF9m4lJkRzO4PhDgxfpTejET81o9CGmibO8sOOnrHYQf9FsNDPw
xXqw+w0ghdOxm+6qcye4CnxaR2O8lQBqKdmAarihjOHi60snn3amflEZtlLcyAWL
yLVLeiFiPOGsNisYr/nI0dyplCYuO6H3HVwuJtCIdXWsNrt89lDL6LLi6MY+DGui
dWGRxQ3g5GnDx3A14f7GC4ZmfYTaWXac/z1gxO1p7hh7iPMU+BQrwJxbJUJxKWJn
g1ot2ZU7suHpl/m5ftUYv1hCw9F+khvSzW2xFIvY5OM31GGJdTnyICU4jNqzaEZr
zX+b/4Po9TEoiAlhOqLkxn3XasGIvisy7AXk2ookC1RYlWTT+7+CRQ85sMQOycUf
2nqNT7iiXJ73k9/JOjzsc5x9NxrZ8OzQQ4bX1LlPopmFi1WCTcBblxSH48Melc+Y
3h38gOZIuQc4lsFGOY/CLyhUuNe6Wzjd+iVIruubqdVRw5u4Zm3igRClgL4dBpcx
uA+8+nFwHFH+ark3ajTq6MqiKcIsxTWhr9TmQo7f+LwbhZ4Jm5EEWTr7ujLuXXzh
hL2EC4NxsieU/H3JAHeGdVeosYwdB+ksAwRMBA+8NMe3Dkx4FuVOe8afTEWOvren
gIFdiCAP8zUpQhjNym7F3D1oEC1bDiJQyLV8/tsGHvuM0USmBkwBjP8amb+V3dG1
HwMeDSrNsv6j4SziXRpndQuWUHp/jwWWDjRfrp4UVaTlvSv+Pvv10fSJG/qzWZS3
DBUbueaVsr9OW5dWrzljM9DLz4BegJ4qvGhVJikMQLQolLpCGIJX2e9qiOhKu/ld
TYqFyuneOBeBDf01aSJBcEiQJleNCR2v03WYmPVE3cusYJtJP1G50GCw8k8ZfFjq
E2/z4XmwU39/Ba5bxSW3t1KH9iwhOwHe8Xrc4iNLpfcrdYO4fOsyO//cfdNhQ3gJ
Umm4suh2ydPEqtzVvr6X+jaAJSMhN53vBDL0/4pqUKIVPDlR2ZZujO6wUbQHc/g1
Cwzgfe9qoYbygrDpXZB8hRvoO2HW7jPgdbxOdK7kTs42eB/DnZuczlEA+j8YxAnu
SG87rrOm4T4AwxO9rmrRtsGS79kdLp9mH5Km8/UvMkJ/ko+ViMkxx2Hq4N2CtLk1
O8HvuwjsyI2rYJSRDMGovEd2JmCleKzH/I4eeg/mrXW4BKHfseiL+6fNF8VsaqVE
GP6I05zm+9WLgdvYuU3kTnV69CzrubeH5vm3LB4CuK/Ei55icsrpbgFfQNzP2MgQ
ZIXni7r99OS1q3MBxpK9QMu2ac9TpMQRJNNj8hrHxsqBJiDaI5O5qPltsPz3Gtp1
SbazSR9DZbdlPJGx15/bLtvXDN5DbOe25mVrLwMi+fqQuFkYvDKLQW3/MiVdnKvG
JcIuIOAjkhpr/NmecZbG9VAhLAH7n3dwppKCPD521Cnr4HKseopnjBbVSfgWDnQk
/y9wnqanQ3MVoPciscwRbq3A+td+GaFThol3lD12RyzFcS2CG0Z42nwpbp/BTwC3
xgnpylxEH1nBLoZBikGbbSwCZTSuJGnzP2LXbLQc3vjaP5jeaQGvo5MwaMxyT1J3
MZSyJpksnw+y87WnTotaDt43hYFHdV9nvZwHiO1tZHDa8fZOhWSajKIM1QXi9Y1M
eupB8B7C9QytZPSE8xN5B4PvxQ+lJx2Fu2mWZp1CFHV7Plh5W+J4DjOwcbtU5AsO
CAKQqV/hVwibwm7yXzD1S2JbnW60n5RKuFMQXwV+Wqm81Rjx+h4A5tiEmgG7S8MV
nRxBAeqyQ0//wgtl0VJJBqBU/Eqo/vve1Yklq3lBZxMvZq7FjQDVlnCJqb7dwZfH
/nGtlt1GQQaK0e7IqeLy/tdD1f6RXuXXqn6zzmVt62rQzf/OMsjCMS9Mf3PW6cun
M+7fwXNcoYTR/9hCPVT9wxhwe9xzjXsdxSthcAEyLwvPsTGtcLordWerxAr+X9XF
WZSVgft26sO76ux+H4ZwW3xfaZ0jm4t740X/x36YhgQqDsAveiwRaKrjAJef5ZG1
UhdKgPrZNDjfvNDVV27YLPAzHd20EgQlvKHlZsJOBEe+vMETJM9dQKN43KzHPVTW
YXLzBvhmJcXiQEgYIf47iFKgP4lLZumKewXchoOZko2H8xoPjpbk4VHcadBVHXRM
QyIYb2d0J+3Iz0DbdQoA+ksWdXssX+Ml2gUROCN8fqZhHegCuIL4DkDZshc6aM1D
i3hQ8sU/t4/pGxIYRrE8nyCbXjBqQMWSLkmXxC9/ZzYA2tuJQhiy7zTS4CxeuQr4
TfLwuZjjCblPgfKva9uUGKK5WV3528sGwCBC1ft1WDVK0JV6Z5y474rlL81eKq2x
3+sCtY9Y4m1XWT7aUp52+E6+3yY5TY0yN8QD/CjJjg7t0zrhkLOU5vWNWRILDMy+
CAnm9WRQn/R5KGatnvUWLZt0Du5Iog/uYeVZk74El1jjANaauT1OzBsQ4/gZCFWp
g1hMH96bda+UoiS1CcNFOmtQsR/Gh2MUHnJH0aGhTX5tDrPt7TMAt0N0pMCAIoBx
JruBKeWM/pmJ4bw5BMtN6KNSR1xPTfoYoAuGcKkTC/PpGTwGm3ydoKKLdU5CXR4c
SkOj9YhPH8sdw1Tpe7ure0xcKXWQ70gEuOSebWNifyCWwwtaJGQchI7tDVeHESTM
v1pCpE56nVshbHfjjfC+G1FrgWWf4Jt9Ynlhwu4f43sMfjLK24qLtGhP4LYuZXzE
n00iJMlmDrddVXkuqJmRhZ6kJwTgUEJwbn5DiHFUcCQPwOZ9LtsuAWc9wAFK3F3g
dTkgP8K5/CkozlGg5OQ1HZACyDJ1CtVJtRXQENjCmCx6xveIotmqK29OkuoOkwnK
0wVjavEyxRN6QLfEeQmaUsXRnR3/N0j/mOVnX1g4XW2OCtzQIoMBH+4S1r3CS71H
Y5CmoygfGvkicJGEI8veG6CYrj8z1AN0SRVT8nenASyIPwTa5cEN0GdnnMkEG98i
XQ9eEA0tLcDshjuIfGyJRrb21l+LJP+klmRn4bNOn/3O4Z4jLNIY/Av1N70CXbLW
X9AvNcZL45YR/qRwBjrrAt0HUw14kbqJsmWZtL3sTccB3/dWAcWp5d97uE7qICx0
/qqCPmvPw9wPrYENWz1qsNia5iSKnDRRB8F6C6YwSd6YB0wGWK2U2tsUVXSDNhY3
AWQGcyT9ON2v6+L6nrg8DZerbGbQ1bRj45fFGehtWK/7M3klHkRUnWNLlSwf1hsl
+gv5BZyI1hY1e9C5esZfy4YAJpT3ngkiGQ9K5UvvgGKYJzcQFnmmo1eLlUb9ZjTy
6mMjTdTlJty+IZKm+cl4f2LRW1F0AfIt/8bRTx/wZEFIBVW2bat4+w4dPgQgtWzN
DcRRNIt98THguPR9AzPr8alAXHbq7gjoyICYniaMjWyiE/89DpPew3st4xlh7wow
cUdSaYYsXQvevGb+bLRdHHtGQhY4cH6B7kgHYvWY4Wu19jimKk7Uw0Slx13BEOZZ
5s2xDDYVz89AQHRScNvv1xDBjWLlk1j3lhC22KRWtqlofs1D+DoFY99hDyBgaXCn
7VU5egVrZC0rR1IbjSNwJKtclYArlBd8YasmV9E6BLXaJjMF1Ma86fWc+oUd5Y0l
977SWr2DjfNUjkO6tm0EtGOU+36POqomeK0IpZ3IpUDWcz+GxMdpN5s61TCz/NMr
mEOFeReO+eCWRh+gGIMEhATjACDhECvsSOOre39YKcTMGh1rw39XaZvTDuV5cxhQ
waoMrK3zFVnl83dI1JJBByHbI3jx5fnlyTkbw0V72zolgWJVnINlfYNJnrtfRs58
j+wZcwLDbtqNdAYV08aLniclixW7igFa/7GHKCiOi62MOiTEmXWltHrnPXqtIvAQ
91NSpKPAWprcVgTqo6OW/+P5OjsZLBywc0lQvaR+V94daCwNSFOpiV1GHaXukWMc
GhEsqh2yZdON3uO9BJ8y7xvqyn9Hv5MF9xLRzeKGRin6qXa9AYwiji3Rz92XrY4E
4mmz/SxrYNRKbpjeudy4vBMNdEoQse1of/HsipDt9WRzUCSKe4dhnOBPWhbVmCkp
NXbry/96wdM1CIihq1xVWXKByaZufiNYvI/JRv1ouSeYbpvPibW0zg7S64a8vsFv
c7PNcO90E53UB8tUQa1j7TUMZVZVIGxb/Id7chgcX2tFtC8yIbiRXrfkaJAaITrF
0sY6ttCnOcPk6tyZ8MZJFc+L34+18/7QEdePQ7ik7hn7IOOiCkMmTsGOS1IpGzFw
8ouc+GMHooXTP89Y/GmHN2kPlBsR1Ef/ABgtjlhyubB0MfBGpZ+sRHObEwnhXK4X
fxIxdyl0gRZl2BelxLDYq5PEIqv1IfWmz6HLG9tVa3ks+g0HFts8zPCKUnOCApKy
LXlLbNrQCH5Dnjh1oHVF7dITqF2l0IeZPpfDdJHLpqPi6k+/FqZ9GaiUc4JDPwmS
8b29QQwh3hs1e30S7MfKj+52JbBUVLEIZpVNik6+PVF2TujbrDfM1nDpqIG6nXkR
45yqbBsTRDmjIjpF6jhdnvDBCltVeeSWjp18mnLeZHLNkG4bErUvAUDfin5AsikK
mcwYDIIx3KlNHfuimrYZIM7SBKpbInhW2re74R3OsqbK+S0iKfGFjFTGJLlz1UFO
1s1hEMq+Esx+W8KtmZ4IFNSy8jZHzrY+JpJtYjQ0tPeBBA8TGKFZ/BaTLOqDUNPn
Vf5lI9rL8wAfM9ow88dU+k9Hq513F8qiSnO/VXl4lbuk0epJ5TmI86Q+8CPLaME+
T7UmFJ0h6eH+3DaGQf8E9y3ORSPqaO3yIjU4WEHK9L86Yiyudn0ZbtWnJmymX5ks
X3FdZWyYxLVwH4qJWhdUPSL9YMjveT62jlXCh0FG6Ts6AZSRJSRpZReZ1/xYKLff
Rsy+Jr6Tjeu2W2n1xIeS+mEhUa2J+XT/JS1VDiXqezx3mld6fQtT1qbFdga6RLrk
sJk83zI7lhjEHFHPljYOUQml4XsRJlBh3b4GKJNOqJ8wRBqhXBmQqP8fJFhyOjy4
7G0SUtMK0GRvJOs6WvGxEU6xIro/U/lSWzJgUshQOCqg7elZwe+Joi9OYscoVfK2
NBnCUC639htyCPAWaS6vB0+0YPWYoXCxkGsRqxWmWgB/UiL7WWNfH8t+Ieo1iG0V
L1mzYwex7SSX62xHsR2tzqSsFEmZ33t6Dhg1SB/8kylJHBQmqI5EP7NW0LSdmom9
xZk8YXSPe6/GiJ0b+NfeK3AYsJE8XjmFHugBW5TrQ7JrmfOLsJlJZurt2k3dp7u+
F9UaJbHw9ZezAv2Z4DkiszzFpRB9T72GLjTsex1qP1Uo4bFk1jV8sfrqo7dgpuDD
YPjVnnp9csalfPtzMX2enVaBR4Ln87gbV9RaHYPdzfBwdFsl1B2bf9f6fJQQ2wqh
Fmnrc4eHioki3gv+nTXFocbUevFbrgnYGsHGlAkpMeC6IeN2RTl1QJChomBMsYXe
QxP/NQg7FDpcsEKZKvN70iaiq9y+tazsYJiRNQZgHbGNc5rUubacFne2vwiWp66G
4ROewECPofk+aQmbRaG0rDMh470QoaG52L0jdZWw5lN9s80DQvFyzqZQFWZ9zzJZ
Ve1XfPq+OCDa9lLXawxchI9dWxIzjohTCtTng4BTHtOxOoGRho0IVHWUv/AeARwn
lPJIUJ67iulUEanNpQmHWpze7jslL/LSnwvizddZsJUPEnQ+DL4G0CXZfWOjngZS
NPhVM/ylPbi7Cwy2lOmPzViGHuXrDtJcK57/zwwedkDSz+TadGAJ5fkr5LpCVOtq
LyJQiiNdrFXM5mL03JlIMB9Lm7oG5/9CmKAUOMRew/QqjeR4PGGHI7B9974RfbM4
0DISOZWkBknnCve6JRH5Fyn/9yews1xglKKRYnR+sbO1Pvbc4gQ1sq/6TxKYAkj5
GUzHD2vfq2s79DvEXgfJU11DgrZBrbIldsRFOLaAl42hSBRjhPiSh+rs2evCImrV
w+umcs1uylHTnHhY3JIhyH5zm+Y5/ZJcKiq4zGMzbONcKh9iIas6AM4IIvSv4dPR
RMWp7kkWXfIctAnJzqKAPwH6YoTA4cRTpjbmCyUlP5XxlDx0GihAh3hP8D5ZOKNV
yBQQ0+ECAg3nYFKAwxcf/3JEn2gSQPM3BcBpGKmQMBNnnDg7rYb7+C/BpCWBTq6S
Ecal6hxuEr5W7yOKWJ5Urlcrqw8i4otFUecD7pZ05+ba2KmaX+Bfwk3aL2odRAue
J6m8dEghYVUnwOGz2/sFE2FdnWlSPho4b8A9gcvvQR30ZTwYQ1oxOUMlZt7blqZ2
jL34L1x9ftJxUOgP+C6/i42CYiaPzTW59dzzRVfVyI4RXL4IrhgXnQDWBi+IE6S7
F9YWAQUf80L01dYc28JpDkI7EvxYMoOA4g9+4DDA2C5OBYZqHAkKu/VOdklImvTd
QUTqWdXNHp261K4UPofJorhXwcXFrA5S7hSz14LyVGfs8insQla+9PJoSn/Bb3qT
eLY0d+XpR5XrIcnM1Fc12OY40J79VEdSK5fBKLksW8gz3HZ4wKMrF+VCyquuFWSU
khuM3WvXCaCDR6UGmncJN82/bDFkZo8X6NOSUO2X/+K8WTVCLGhPooO5w3fAIva5
L2e+TRhnlfAk/18RNa41NOapBP6IVCcvoF7F+UXumui36kSE4N0mkAr4Fdflie1H
inukQzpdUeB4pNxGAO1EF8nUVhktKiVDzVUvkjQCMtpmJT7GKH0kgTOTSLdVuSyZ
bYdriifkcf24rJAuEy8/BTEm96GxdFrmVPXwHD8fBZCxETsf+k+71djoCV5Pnm5q
XWedJiWFyj1AUWZUEwKDUKT55XErynA+blOFhC32cbCH0Y8BobWM+LIjC8OtOTsP
Jx5eD/1JCmwrumVvBYrGVwwjRiCZ0LFoBB3AvDs5ltD/qyPQDfDX/YLexyKp2cRB
GMG5Ao+M6JlH7FNL2uECIHifhguW9B/zzem89GyCFHGdtRNiAiaAvnxcchyVNjPD
jBVESRqt+MAfPq8xwoA7+WLkzbYWF1mUk5vP/nV7rzh9VBIsGcEr0Wel7fLgg9DY
AW00kQpoMwww7IUAJbSEFDsd0Rjv0bXrcR/FHJKlPh3fQJRJtWvvPDCHs83pF1ns
duFCKtuPTOglucEzGxmXgOURyC+YbLrAOT2/nwxlqtMjaWPV07G16iQsGccOlJ/3
r2A2VDDzwnWewgpJTeXvlmXiJYOGKkJLqTr0L8ivaEZb+Ns4MlMc399Ui/haweUo
z59DaiA3fSMs8S2/8IehvKYMP+SZOKNZEfHtVFfX7IFt7R1desQ5rCh3Dm8UZkxm
2l5NyGRfLo4Aes5DnarP3tCYMvbrtHHrdEyGUutbDkmYjnVBznSft9rd/bI2gfHt
P9rse/58U5fW4qMUU67nE9pq/l3pdBbcU2b3ASrZN8DPRq9qgGuPT8Rw86+DCeT8
636natadf2eyWR+jnSTCpHiG57i9D0jVD1fMWSslMdR39RJ8YwP9qTaPTbWppsJ3
XH/SxRDrBH3SLoOC+zUnaxATU3z72m1Az/sIqdM/JpYEeS0hM1OPYpAx5aKBBGV8
ZF2zJLrYwS83THKvUt0zycbGhpQUoIzw0fs+iIdXswBxvfv5NL79Y+/lm+En/lQs
YLj2mlys1JtUxJrifeQckYpFZgMIEb26hRAk3XeIk7Pu9KkBJIwMpm/eMqrVRRu+
Dqec9YxRILX5nQtmhoV6Th190HdM7DS2lBNMlQ/z/npHjUL2kyKG1noOwwP5EsIp
P1XT2g/YpyUN9ciLLqmA+7S2zpYbb0BYy+egdPEFcXpxFxivQlRtqjXSHUb5ogns
MRIIsyCg5zvJu9lsGbI8BnE0klI+ceTcKXsr/+sI12IaXbBTCmJLLMwoDMgqRseo
Tpy1eUje6fZpTK3mpLYIRyGGp0QaCY5cNuYUJ/kJ9QDDLFHJ0xctVQ5Q+RZMAxO9
4uEH7i0FKTftCq/RZEwXl9gHtmDJ8X8RAirRwx+0PaHB73XDrzCBCCqYcs2zoZLA
nUb3oROP1HViZUM7YV3JAfMGpy4OEWfgjyqOFOUBZSC1yUFrbb/VRdLX39ZA76bL
HlAdl6ICYfcksymz1H1UhPWBUdKKGihvenVbx3Sb3DjUEWncZ1DielPvebTFVawz
UAoJlJTP/Sl7iqiA9v/Tqs/MWKn02rwc+3rCMLPgyBNlRYzCZpwDjuArgClwCPkw
YQmSfy0Ph9ru6I+fKEHP/H7mbVlCFcC1ThCLAS/8iDYofDAMYYgOFlC+reqgrMBL
EERm32ykzqCuwG0SrZNa8ECpKlldXBJ+xq/YFbF7/yYB/LGdOegBfFagsSVoKtuv
y/14Brfab0oapbKYUkM0tq2MWAOrBvlq2swyDHocp4dVrRqwlKErpHH8ccTaKPMS
1x4cscE6wut7ARw4YoQGMzEwLqQuPbgq7yhsyAcZjZTbikqEGRtjHpOw8VNNZfsZ
wrIJk9vnzIAOvoeoST81UFrRelj2eFqrkL/IJx1MeECauPwANDderDIgOFizkshm
IUx5bTW7LrK5uEM7xMKkO4YALzuS6JDPVKWB1LKO2pBfu++NFyF5LkA7BAASzfxz
dlTbKfEs4AiTfQlRMRZSfIxfT4Bem2vDlqiniGdBNl0JTDXg1fDUfyGSB14r3QRy
n/KTbmwJX+sbNhq80zW6EN1i7uVcLivGyQytOzlFeIp3R1fSIJrYWWHFzbQODRiX
0Pwr0+mRbhVph1/UCbM7uJOhbdeqYt4jztNqHPHBppbpP0K2MT5Fd7agFmAq1Wdj
wVa8qqFh22zLpD4JhbFKzC+br7vbVmF3p+BLONfxCzLw8d6aiOVXpYdtXHHzvwXC
dwTqshQU0np8zX5UY/z2FsFWL/UZYq6Yh+4cTFbEHZheBCgNO5c1gSVnys7H4uq8
SnUVxqMQhsHkqBV5pKC7YCsvfvwe83rNEyEO592UprrNBmFgtCHs1OpxyKQzQkmX
P/8pdDFzMVa1tiaxa1tuxbSZVRx1Xeu/bNTkQg1zuLqCorssrrmZqv7TKdDWci/u
FbHnDQWP+eIH1dKFsje7NdoNlSeYZCX6NLpuKUHHKzGwLnCTZz2j3v3Qh0jbv9qJ
f3VaJ92r0ecpDWnwxcMQGZLdkzTYX5ScDy52JnpzR/pIV1SSPAXXIaVCVgbyF47N
6AswxhaZe8sWoKL7aPKGkkl0TJjNMPqzPAh5yRafppy1C/Ctk2RFeNFRLWH48yU3
0nzIEuVd4i6HvyfMOVudgm/gozdOHbduo/L65O5mFGHz85+ZCAyqCZ/uJRUSvkqe
zFKmdWUQClcu+rfkFepVMakOPoQWTbjCcklF3uUB0dFwLbPD05QKmk/WK4YawBQw
sIVi8v/a99gepjre4KpgTwmjQh8HI5WhCcXDYfIFd8u4+CppHsvdHXO+uy/KBQ2g
Xu9zdoftC83OWqa711PJKWVWYeN6BQBA7v83LynaLxausDS1NVVJEg2S4S3u4He6
alSaYSFPbCwmHosgXgXnfUYaAGy4rHM6rRo1Oh3Uwr0vhoSlJHDhappOvPyaz4XS
M32JpKx2L/OUNhMwpNaLHsbyfiw5HQ7QHVNIVstGsFE7g9M8X1cTtEbUzOyby9V7
z6L6oUjMT13saH/UpyF4jAortAfsw0/6Hwbp5y6gSABQ2MMaMFVFxhynuxn7i6Ns
a20DCSf0GBO5BJTtztGE4uAKJu7OEkrZKzVVkdc8R/9fivUjAwCPgqW7oSNCvhqD
nq150c/i1lymCloPdKYflasWDjitEM7Em016OSQLhM7nMat8KQT8ZKcgllERrc7g
tXt0iQsCDsAX36oq99LsDFns/GXgqfBMraabWZ3Ah7vbDw2PDnn5EdT72WoIkJ6w
sTgenH9I9ToDVKMiZZ858qMd1ZfY2RC7a0WI+dE49l8dEp7iAy4tmoh5ucx3NzdN
T50PpPp0213EPNc+dKJZBd68GwiFVQrqBEv076tbCQ6la3Ac8Cwa74GphouHTCXL
kvYzs46hX8YxJcsiJO6iPsnXLd5rNSsGhYLs0LSPyPXR2c9ocQBZ8lBFkYLip/py
SUzFcbB3zpWYrdgYfBWKPhZEYqPVUA07QWkfGxSZuyDPRfYwFIuLFFsUS3sV3OvI
HbcvJ4Mex3VsJXOVzDKVmqj6piO3xXbcpXF8+anGYN+aJN4esfSmetVTHUJd1gDZ
c4P4xY+9E/aPL2pv+O7O4lPk0CGAcf3d63NOk8pw3nDAhX97G7yJmSzTXQO0W//c
9lbLa/7bgmMjpakwsFbD2hKGZX4fbS8Sj1UyNXAsfl/3AZW5JlvunSpY+80wVs4x
spBZyEVqiWcaBeVP14ePy6I66Y2mV2JQtAdYt6n28pFftTTpRmXldf1L4/x8nDBK
48sINU9wFf6hwFk1VaifWWUo2HYdtCQQ9jFFNlfnMQ4s+294DW2jCWXbfuaTxWqQ
zlqgXw0OJyKM7D1SuXFjPvBhzXl3dVdXifcVymTbtZpyHv+DG9CICTYCQ7a6oejj
Xo7T8uHKuhcQA0v+oiTXqfVMsykSlPz87LcWafE95H4uDEvG7GvvtxQ6AqyHMYpB
pJb2S8DF/rxPqxigmUBMfwWStlsXruN2+eFulpD8Vb3B5rkLM4wJymhiTZiZjm/O
J5zMFCGSKKc8KfJfis8EZNnJbRccE96RQBq+msN3b9Pe30vSrTKMOkJ2JL1Nbeuc
6n2Q/ioWmAPaf8QkYeo9CeowcXEu5Ve4sURjJRZwgT9+TknqaHq9z4BiYMpU8FS9
YRcYTiuZakym5cyj+258LDwGEJMvZgFr5QMny5x/fatXy/6nkUNVs5J3iZCjUUvM
RL3AcrAhoZYr4A2KUAqnmxRxAlvLzXPYuxEaIO1P4CN2KR/bp8WsI2PEXV5mFuJE
ZXj3eGqsfzRjGUfxhTfSUiUJcqEovxJZa18x8K14sdLquMfeZ0RCWNBy0qnGvPhn
ml+xHHC75SvImmtAavQLQPR0iLI+vj6+3I91YH+UARfh1op9kBtZTUXDHOMKktFJ
eAI0XiEWWzfB8k8KXVv5pxs0JvkpBFsycEhWNZSYJLcOyxSwvUTeru00LgHyOOwT
KFv7WpbN0k/pfrQMflCrCixGY8u9UNIKzk07Tgnt12Su+TXF+iOzjD7fuTdBgmRH
9j14aGni6w3xxcg+vqnNDx2KopD0pkofgU3x672nYtlBLasHUUN0XEmp8+8zcU2W
uWpiXgr5MaSgX3zxYH0qPCQVq1mSlKfQ87RQ8EAMZ3bB4wrotJCTFMOvw9/cUjs/
6DSkpWvvoVqY5YltDJGwcRe3HQxtdqM5DLMbCOYjwZ23OE6g4vasRVnG8xHIEI4C
HHV3s3ZSslN9mQ8CqoCxzQZPU42f6W0GUPrUdXXI2WZ0PT/VsxGGTn01MBbZ7d+5
+0SqwTJGCIYzXrj3F5nAwhJb7R37RP8qnm057iXFq6YT0CdG17vhNCiGrurhxbIw
+3Lc0Fb8cWQ9W2fB9H4t4wsc6zH9wWzrAf8k2nk+1yg+68NqUrZLSgCS+hqembK7
nNyO+czhxRWaIIEO3gmaCpLLx8tXU+nkGHFsHgLdPLm5Gn0eNZThcdTCajqU0APo
hC82Gy89m1pjLkxIDkTphMEp8F+t2bWwToWlNM7Cv3wxrs3KKPMnY17/Y/XGrA55
AbcK/Gr/K4r0lP/+pAwWsTLpTeHdGviY+SizyNEELwYO75YkBDbrem+dUarlOz5G
rkIlAc8iz5kvtM9lTCZZVDkph8LTsqHXGVCRF/mXPstXStoAh3zqQqhV1i4u9qE9
13s0vgVg2jN4fes2E+V/AweHxYDNUTK32yB7lx3PUT/uZb2DmuFA5HDToFEPmFKd
lZVayVJa5zWL9hXVFZWZDuGxOEBeDDI80fCyfsGraUQFLvOA1rRKlSmh0EoXb1Uo
gl67UdaYAoiZ/23fvreKJbxoLbp/2TlP4fVNnfoVDSqwWimO7p30/SbNaPOJ6tGv
7GxbUtSsN9X/3Omya2m3WNOoso58RjxQwPtgpWziv5tUhT4tPb0Rk6r3cUzpw12L
Ugic3OzP8FGRQZhCvHsI/94sh/xpVqT9n1bz5aLEPo4/p1ZTwepe3SBt4imoydOR
edp5utXg8UyRLeIB59E+l8EbwiOQMQsBv/J3Y9TT27ykpsJ/NS5E98gvKcwaiV8F
0l69xy9Zvvv0lvdOyb6PMaV36cT3Q8IXmZmlHClCJYvriCdlsioTgrpXPWwwrtkk
/CRCmQamJDCEv9e9MdULqENlh1DNwCXC1xWTlREoAyg9Uxah/yMkIi+/yEtPvydV
LO9piEw7aSrshhHxcnB4EIfv9HX7QeEBuRUGZPYo5hQ/mSyC+JRYGi/1U1y9iYk9
aruQePnfS4WVbVpsKaact1CpksPI7pPKrYjQI0DEX+6t7jp9mzDpoXwsnQRGZrS1
t8Hp/3Q+R+UB6wTz3yHBpdSOjIkp54jF973dj2+XkNO52M1+tcUePzf/qgXUyLvf
Br+qcXrtEDdfLDgrI4da+MJRnwRQCtQYQGqsbPs1RpRTSyh7OHh4HB8Vjl4osoRS
KmG1iWTaXODqlZNhvMAyJfBICq1dYCs0hmnEWeWXXhWNYDvrVfe98X/92TEmOeLL
y+4yph20NpE12+0uQdaFGLVA0tiqOFkpmr7/opfGMs3aIEmz4T+NylhyMoi1Jv0d
WUnFMcCXsJUa2FsLHpoeRtFl1g8KdidUXFYR2eQ6JcWOf9ez4FyQ/gLnzvpUxJSA
EaG1xd2pCpTmnMiDge5vGVQPBVju7YB7MpGTKwsKgIYlTCqZR4adrt/fPHJr7+Xd
eNvxHl7Llfc9QCoinqfcjzcJACAsiKLlyEHphSZ8t/FtzlxfrVevtSdfH1Oy4YHe
5vkiaoIprb2IgS91JtyHMMUVd4+v9l+BBNfHxqLUWbfuwkMEeaXNli4EIxtBh2x4
+8e8D3nmtYMwZOk1wUIwyNPU3VKA9A9j+NT3TZx5tYKk2c6IeffdSxVkf6tAyMLp
zRhwAYRSWD1d3p8pT9AKPLkBvoacEVwh3Tm7Z6E49uBRv0DEBk45nufwJXv0rgQi
9XnQdzaewX+dbsh0lcEuefidk4Ij2QF1LGN5hB9EpJV62i05Ap2vhSDviNplIx2R
oKf5kZnNZI4iR763r+eVTVzsxuEyhtdJVAiKI8nSYRqkhCplnMU0NR6LxM/39e6j
OghmWYLJJ2qzWoU8X+NJoCWpRE+8fyHhXULy2RrC/cx8HP3PqjRsTk6y4D5QqDI/
mvYRX4ccjPOTH/n9CNkVse9b/ay082tGbsghCRtXv7Oufg3O3jPy0oVpZy6df34J
F/dsVLwi35dDHak8eMTS/cOBVHz8GYDjEYzCAsTLPzxXY2fBJiYqXHB+uwQdaaHQ
LZmulebiNctnF3nt5yjXLMDbWRN3AWTzXKdur08JX0GD2lxJcQeQyYw7Yu9wA4Ib
dytaz5FMP7dOtaaXVreVhZ00AcU1uO+T3J4CBopCUwhDWMYEn8iAMgRcYUfWl4BP
TktrCTRW445RPT3rbelRv0wbTGu0qKmKMzJt3xUZRG16lrI+bhMxJMBrQFxImLv5
MK1HYtRF6HdJX2Q1SlBWqTSNfnXqh/fLlB4gnKmQOfkBFuXPxqSCnayU0+Mplstm
aJHYNzmZF02E+hgJtZyofOFpcJWx7vDrUXx4RDXiw2NZT7iz+SEn7lqggSUr+uI0
9yQ7gfdC5rweZAjstQ+wrZyJBouC99Vu8HTBqZdIY7pIIgDKGqf4G6FIpyK0nh5Q
c7IDEJOK/lZQbPLd0gGtfQu0lRARx5t9JRgbu3OPt5mtQk+F8jrBcqbPDRH0zHyB
Aa2lE71oGk89CTSCh3/rW+jIOvjcgyint7eAsMmsd76nqJ60NHqjVxlJkWOSotHQ
8KGiJdSKxnfam0UWdq80pLzsrgNXbxPEpvUZ9xr1Y4nBFl1VZWET2H1Ta9AXehfA
ZeDsnrKDjGxvhSinPJuCEwIED/t44+CVXIsoQu89hrEQzT8Gn9F0g3SVmXMPfJmo
t3rvX9dK3nYxU1NLPde4uoOBGrTZo0vS6KSkTs6mrzmpRi66Uq+67BgcsZzFLok7
zxAoe68HdMbwgJ8evuLPypFpyKKig2hRteXzFZjGvE/PMkxYsP6M02KWBdQLx/wU
eAEhgnm0N8kOnSMgy8gcXJ3ynr7OEfNzcNRuNTWfh9PRh2+ZhvXVSg+e+ipTAJbu
+8+BmYEprPqBrShvUdULuCHiT0elJU7hvQaA1wABWIJK9sfLSp39ZBfXvh6RYZce
UdWuhb0Roq2UH7WkqLIeP//L6QrRD6j8fGnUHjq9AknHmEwTHBjdvip8ckkZm/i4
cHv345+KFwwSQa5vgFsIW/Kr4GJBf8JmKvw4uBxAHlSBkpOD7Pt0qSq9+NN+cNJz
Hs44CpEdEB0xdTSY4FnYhtXvJtMRcVJdfXxIcBc+yGyJAEcGwdNpjz7s+hNE8+FY
3qIAsFovAU4B2fVdM3wFUXA4GXucZpj27K3+YNitorMTS1TevHd5CbTm1Q08M0OG
gUw2oaIcin9DliE/Y4dn8mQ4Fvbssi9zNGonBaslmx9Tk2KRRGeZrs/8HolFpx8W
pfPIkZDxknFcImeLV0EzFDsx/hKAu9M4KQoetpTFYTJ5T8XBgIYXL3Gh+gKyUGCh
SFsuOl8YzPWhNdY6VmbtP2NkfAsxiO+O0FPTng25RgNMJZ7MrUUfWr2/IbfstLWU
8lPA/BCcKFmaIR6DVXjMF+el6KgiYBrZ4ddTPIjPjN3LQFkfgeHujod3a+XqzlHt
uOrNOArkowI9VZxiOdNx7HnzFxbi3zrXp44ABaCTOL6ngs9sd2FNzjHAK6L2hcYg
YMKAtdDZNfdd/KCjxuENbXRNV777o1FRLjdlhcsm61jDCyH+jzDSpq4TGerkw41+
M6AdRV490kzPOmRWlLTuhMWZGdSya55dnJHj46dyYo9k5Nz0cyvkty0vWT62TUe0
uD4LUJGJu7BnvQSVQBC6A0sxKpMNqbQF1pvuMljRL3bg8YVuH3/2HN5+gWf2qrnL
jAGYlcRUhj2wdO6BZ/v7eHL3D94P3bFdqEt/zixDvI1Xz5ltmEs52DucqNE9B+y7
0mw7APOkI3z3AZxecD3Y23QgiUog4FTTcAbl96waZRTqWgjCOI882yT6IMa4PiJO
2big9Zm7IMYjbkL+KrE3+ykz7MYmkg2hMvfKPf30GCUDFehTWzdbxhU97D3sWQvW
F2E9ffMNCwJ2L8xowm+6tCI6fSI1nLCcKZCQe9MRnWYNjyeMqyw5B2V95LBmZ0Z8
QQhqvO7Z2icb6J7KJlHmWHcoqU0MlIV/RuK0lzqVhO7iEuD68kmzlp4MGfWm/NHq
fQLuzKw/HLis0FM1xImTeOh/BG7jc44ck7upeRkWgZGF4PbnJI79d+1qYLSa5AxS
SS1+ioQbdOy1/nDuO++XTALI+qkUxU+KoXJbgHH4L7lyytzOP8DONJ4MKuhQK4xR
gnknJu7jNMmXAm8tsa2VRKXzPsZ+1nbpZvRdgDfGq5/UQxDHH3BTwj7WPO3PqLTs
KP/ijXu8AwmQfAnz50FTD9PDtwvfUHe7/mROMccdkZE13LDGroqteb+ggExowglk
6Ntt2LCFUR4xXwPUB6iyuTfp6+cdVBsfkJbgb7iKWn+gTV6fnVk+i6t4kEABtEHZ
x7ReLzEKQgd7yAL/HTXVR0SNNuskmkA2W8yMPflZcijCBnYeLkQ92yXqiHTY4FYh
7XCyD2cCkFfeMIs4R/KSLwV8bJsJhv9VKp1TCGbWuhLD/RAR0qXVvDYQg2hInAUC
ZwY6o7xtZ3GspWjobnHdwKbjLXOa2OtDtu2jrDKo5xwgHyGuR9m1Mj7xNsF5oWMw
a+F91Py2QWo40arZcJeGXgZ68V7LaNTZGQENIgdcDW3trs7PrcYq2vWxXUPozM60
FRQ4AZd6HHl9HafMHv2SOAQOw6UGSsmiZhRZhr8IN7jW4rwlVP2zF7tpHANwByZj
iS4p/rhA6l3aEX+zEgxJj0/OMU2OVibSGi8QXxOll4ull+vaHh7X9qo1L91p8rRH
PQQkHInDjdf3n4Q7gsDtnA/A4FRBnugD9Eh0R8aXARtT87z2sC6ECTYsKyDE0YgW
mybD3+v11lTYwDuYEDMKKHW64DY7FrfG9X9IwyslXsb63N9/e76DP+pP0+ULbPml
0fPRT7K8AUBU4msOVTL59WycZ7dchPBFPO24dfsHnGrXMChgiIbHgdifE8PPutzk
aTwwAdVTgIla8XcCdsi/4QOr5nRlqGEDch96HWqwdN4MHu0cFAtJvC2BSFetvHPg
fHuq4PBpa69hV0ZYOFUMIjPoIU7NyJUpSyVZ9vjHXn9mbyi000Xgw4cNZaAQr83i
rWj8UW42B1+hxg0rS7SALWuxA10S1Mvs0Jq6li2b4vfnMrn0kCzVV3WzL317AXs9
7qSisfWI9gp61Fq3BUwkQk8mh5IMJgfQN2g+a6/MqrUHC8S0jML+6C92oCjJaJol
+uMUA7h1C//GUWJuFDFyMaDrpoF4Brvah2Ql43NK/GH5UU4S+GUTa6EVcD+0eTa5
FelR161F4ytgfGAhT0GbEwU4GwFr0iPOvbTfueMpTVDXUJIXUGVGmU88JYFy33zF
4v/zwVTy28A0jv+Wb/6RsYqcPiOQQ8HjFoscwC84U/IYKWGdAza7eMaZRu3O5q3T
5G78W001JnrLE/IZevssQArLIbE3iADMsVQ+OWq4tmxwvsptNzJUMWlSDWKzi9AZ
Jww+KzZVWy0cuH6c4afPaP+OviJX7XZnP92aMlWKQ+er5L0cH3ALUr9tSMN1QqLw
O8UVp4a6HrhX8Y90N33PvdY59d5JHahXgzyH0Hs6ezyB88lNrWb7WZvR1SQTU9Wi
VYfSrG1RQYtBERMinPK+len/z1Ts6N8lYrdmb2ruzZT7745wplj9dEnhErIm/yTU
U/1rKnJtZxrQSeafXzLg083mtL1GtOciftgg7SxcZGe/s14o7ouhdO6LOvzL8hTH
WeKHoEABKodMSieefvvEEG4hDcpx+v0ATBZk7nYsvz/QQ8zm5FoSk+xkoIwMRUBS
88y8yofhoIQZzq00d7bh8eYlZA8l/59BlGZBT3k1jRcsT/N6GXgL6jCoBXqJwwwy
QBIKAI0FzcF6d8Bto3ndpJont1x1zc0Wo6IoPB25zn13yWoGIljXFc6w8BeBjLrS
vi9OhjmycT23XD6CY9umrgdZGzBWikrSlqhuhAD+L5Esa4OGEHXQZsx/aZe8IiAD
rm/Mh8IcTFOoGIi2iexAvYSDcecEUUgJ49uV2a7v59Ve6wlWoEaBpHqgv535WaH7
0/QwQWkISQj4g243VW9two0AxB9AbiX6lp09PVdQdgnFWRWEonVgSHhesyPo54zn
k2jzqzPlzihMkGQlvmz/HOPXf9C7LPDpOT61BM2y7yw2+/GCTMIFF9tOuImRY7Ub
CR2cAI18/tVyxzgH5dwcIsluRg7o3NLLDUzWbKl1UYe+PZixUgh5JV/vFwsRB8hh
KEi4TK32Nye+mg+0Hj1JgyktqVdD+NplXHHNopOiP/+HwJL/+qY8e9VAjOLKQQKd
2pDwbRpT+2KxRoXnzkqpmi69O8obU6XO3UjWToCM+ErwQkXMi2qXBPq+96Sv7/jl
9knCEXylZTms2qLKnlThL461C9uiI66XFD4+U4zAsYD24ouAPQ4NAQ52j87bxLFS
1iFCz6DJ5uZI/A3QyxrKTrRw+qq2+wmg/S7ja6zxHzv+SNOjOClXoHNZO5qg7Srp
FQrS/d+BRXHWcBv8Gra+p5trk/BSCU6Em6jyvui2/3mP/GpZX7EnUxLNDVY4ZFz9
7Oo/qswrZKcaVxlsodIBQdd22JcwdyTkB5TTzcpfZc6ToAcvoSblNzzuscS9aITb
vR8OtQmMYFisMO/Vww9vH9eayur7Y1FEaP+02d9dSXUySxlPc7AQW3PoggPKmVfn
oVmSn7VUFrejfjFbZ0AfDJdcnt+QRBIvtxlavS1MPyvwbd/1nLgK4Q9ZUKp3bpcV
cTnr2AHNORc1h4pn15Abp++FsuG2KP0pU0hyj/MRxGvZDwLdaUjL+EfJBM3c5gSk
tkR82qt3fRKHocZD9gBCRrJeA7+Z+6F0ahHiQa6ABUPjODl4+lQD38hrV09QJLHG
kTxMXuXaMyUfg15s4qw1Zc/tTOeOkUP8lDS2vzXQk2owP8dGzJrfZajCo8wHfo2O
re+D8mn2bje7Gp3/ZfZuf89FUkIAGE9cfEseZ7kr+QEsHiQaH4fQkIDdBt19+I14
FiSclPYw2QoFm3QPmdXVxAtIRotTtkqF00vTy9BtllWCNM8+myxxQ5lkEkVumjmv
MYmIb6CJE/PLUrFmcN2T5dbuvTvY+bWAvQ5unmM+HdHMsQ4VagXj133U4jFkUAJd
c2vPLy5VN2UxZ4pWdcX6vUzxeK0Es3AIgYftHdBG3B7IcnI2kfdjcX3jW2vV1Dcz
nswn0SjJ3/Tdyz9WKv0pwcHt+IcVgKqv5Ph9wdnceJjNTxZbGZbZxtoDlLPgUREb
MxojlX9SwQcMUiZ9W2iInPY4OC8LyKkrEAikAl72B7p/DKE/aarFY+G12sLqwKf5
hm0LT+21zJlL3fjqJ3+XgfDX2xJgxDUTQ/sySqLbY+hpxmGNla7g7wCMKokHeNhp
ZnNFQ837dsGh/pyUZMZZRQLbv/JkFzIpBhoV850rI88gzXNRjzMPL1U7BCVrEHH0
xn1OnQ4/kXsHd3j5AvOQFLVn59A6rS7bJigx2twwv4O9B0KdsJCI9CIRo//m00RY
yCYa3K8E4dB1xiLqEvAb9/U3yuOlHvFBjUO09rFZLo7KoDWP6VvNMBa1FeRvRFCp
Slz5V2LMjwolAvvGQ+dyxCPYRyrGG4lmKx5jisR2/3SwzQteaAKzuRe49vY2Aw0H
/+BXipj2LFN1uZYkxrKmaWbpQHcgsD9lAGCX9e4Kx2Jaiz51p5Gt2syeu7bIg5qi
or85yxWdCIbXBVoTUMAf9Z1Admar5FUNHQ2ozwi9E8XZHSI/uaun1IJZYnyaKi+6
0fZPec+ufUcSoHCGwaARpUgffS49yvna9ajWg8RHrh6WIb5VVyc2VihsYmlInHvj
yTP4V7Oq/pptUyvZWM8GegTF5g/x6YQYSXJoS8r5RhfhS6QxEtTBOi/v731hPy5T
46/yKlnGAbA/DMNAkGyc8L9/LM67mTJW4QwD4AISxiYMWXy6lka5GP4jm5OH5I3t
xDJdks1yhBuU8ktfiO6bPUlF2da0z87evTDHTL171PA3Mv0je1koh+njaskBGbIa
F1/j7NfjK7oL4IZPdBLh5ya3sndpPxmdDOIrfh99BYCh6cqSpQTFdal4Ut4Jut1x
MKFaPzmIh/zzRQfSGXH/o2ZTPSAts4ETX21a0FxSAFUO3s1pZ+4vD6c2fbVD3Hzb
/OxH5gX/rvwvuarF8yLuOsUtrb9agkczGL/89DPiafMlr+41ItlYGOOymG5oMo8m
q5Q9G/JCMGnc2/5+3dk69NWMDIbI06FiRIHME6tVe08/aA6A5EAyibbixn9/5E3s
osOeY3i3SqBww97EK2cvrR9ldW+kcWJytL78j/+Mzgbu/J2B/n33L5lfcMT7HUJ1
vFSkkMM4f1WAzXBxFRYZaxUxyXSyJbT4Xza0f63IPYkdzw2qkq9KYM+cFyvyIhIU
PuRRERRhjOrTgW8KvovXaB79OoH0+dntRhPAc4QaAN79FwG9VLN0/KuMtpJrhs41
0+pT4+g/lRLAEEQN+rVhIQPK65PoMvxkzPPqGhsRlcIBxHfiBMLlDwG+pIvsr29F
YLTe2TcVL7giNeAqM1X6V+aORcOUwNz5AawfvJL7I2KM+0megA0lgvJok4EDRe57
2T0mYfxgL6rBRnoRhe3DQ0OWkYnlifCA3HrgqVn/yMSKHz3Pn6CnBGMWQuzDB1Eh
HiCZ9rZKsNBDm49XDrVZkXHmtFXgWX0rOmzVGKYT+ICJM2l6btij7YFimkdXiO3q
OVxFtMGJajNGn4K6ogjZW3szUTUieohjUB8L53lqAJ2sXAbSY/g5Rzw0gPV1GFgZ
UarE0fJLJYfNf4x+TnArw1+Z1rjLuCKWhuDLlNpif5MqTUwTATePUofkL6EEs4MP
BIAO0Dth76KW5060NLKYtG5e6SE3fdEUVIViv/w9mh1S+gghz3zFGQ3Y0k2WIYVe
X+QrX0kkZP8/OsAO/NMtkAlJuC0Td8WLrM2vaTaNAsYtDsneSSjdzPKwPyKPrmTc
v6duJzs4DNy/pYpHMhe2CvDBQnlEaKSixTDe39kPWj4wvY1eZE/QYTnzsTxm0M3K
ZqpsKqInzli19/PwZSGbi83uStBGnDCH3L82eQmSsOoU7qJfN17X7SyaakMzN11J
ol0oFFJe4T5A0AvSx0QjF1wwbn1TEfcPa0V2dpEiYfO4TjGyBVSkBxQZF1ZYlDQE
iubKTwxF/xSTUF15mg2MUZBqCO/v+MfbwQTeTcgUfo5xllXel3KYXAq8g/DXK6I0
WS0D/mbh67IxKyt9Y53WxMy/CI3fosliSEg0ax0rjr3WK4aYZChtmJrLRsEIqF7t
pdTL6xigVpIktF9Nh7UEYljaWFqve8fHQwPM3n90vc6sfTQoy6/tnQR3G7S8+Rsv
GgtY1Wg6WXk+ws1dfz940p+/4z0Srd+B2w1N0829gMNKBVWXBt/w2y3ks1m1epXu
HcByNNPUqciAwifnY0bOT7TQ9qB05UygWxSdgqlvKIXZqcJfklam+S4Qqr3qlurz
vXI3V2uVAvokEm+tSbH+j1PcoEz4n/Bz6EeCQ0EC57IMUXMLk4v0mjEd3clMZ8ld
IQoYLZMZp81mBd1+g1FpJOPoEKZeFzNgQ6VzrlbKmSwq6JIdk9rC2JROX19wssKb
D27HkU2wxwCDC8LgRj7ShmFfMdTZ7SdSVOixrlenSMQdSElpOCFMpU1mbNEOPvL0
uigVW27vKSsS/csCR/0gf/BPUTloIIAhbAZ82tiXeONsB5aypd3az2HTypjWxYA+
WyIjiMu7VlM3Z62AELYDSa+zBBy4AH7ozjM5o9lHALLHdY1myy1qQisaXgLXyMRq
p4dmfq8i3rcrTKNzVFO4Opg+qMVx1wCxhtEdcvlefFuuuxgM5uzCEMNH4gpxEaFi
J9Qkfbp/qD71T/sKF2sDMPeKkMB/6XaMxWPpa4EMt9VMkl/Wi8z2xIHvGNaLQQlB
3P4XhHZFJ744jEUggmDPJvtKYnahM3DC0YelsMDlQW+BKwMWpSmcQxWa/p5rJnRh
y3OXQYgXogOom8NSdG/oAhcwDwnqJQ41A8mP7yJjzBTuJ7PfsF4eWz+Ku+VJT/q3
UK+fBULfYzTJH7VtTt35HNBy76HUeONRbKY9rjNP3ydfK0soy9fhDGVU+EVXoynd
FqlgIQJGqJxfEjQsTW9V58I9TzBX9py/goT2buGuxGfytCuzo2H7CZ7ozd1Moup1
N4xFaRR/WpjONBbnL3tiOwOGBkCbeklAlccEEOZDISpvX4+sxRnl9pKLUx9mPNS3
+L5Mb3d6WPc1kKz7t0wctKgtMz4Hjra8qcyNbQP62hB428A4bbQYkoHK+de6gc+N
ZpMLVsqlcd1ZatFKpqwXsICjmOgkHXdjdvOVE6ri4ojra6E9FUOhAn04gp0fW8ho
Yt03WHYPLI7NzjJploFpRiVhjhBLmQbKe2dyUBmH6c/JfJtfF/pgqBUqOEnGAPMO
AA1Wf9lqp5nx6OOUANYbTQ38JiQZDZsSAJDuHBvdGAMwZ2/H+26f5WXiyyrnrBOa
tn+4WAUmCnzYnkZR0pyUeCZi+Q/byIXJ/VTStv1UTCvbCFGrYfGDGNwwD/TJPkFC
vyWR6qPiF1rYI++9oqXz0IMUfEer5M63RfN2FSRlU8e6E0GXzN8SX8yUN5P+jrjD
oLD2LJYpHljXg656IzYpVmRWQlA6uz0c/EAMGTACzvXBN7wejYceVX7hvlS7BA3F
Gzz/gNgGS2G8VD/kxcjRAe7K94n7L/OaymGQJAqXi6KSNd6dsZy89TWwDM+HRc/q
5ac5LNDLZMv7uBiUeZw2nTuDQMbecYnYoo+xx64au9AU1eBlgEHkt43y+2T7sC9N
VVTMWa6v9paFjiaBlnv7bykjGALT+3ekOCkucPMkS//Lqm5WhDpDo2QWb8w679GW
9Qjwh7T7HSTnNDozrlN5PsZMsLQy+F4frTirB4NyLOz+KqIW9CYLCwbEkny8sp6o
wVH40jQ1TWTfxW2rTC+5lERW5odqC32Gi23FgK/kyLwaLitYsMZDG3glkfPLOgvv
2j+KWi//gCFXrWWEHUDTB6zFWFDcdV9ithE1iKF+Ob1AtwPMgR78cPhIxABQIgMT
WUyVjQijW2z7JZ3l02p5I16SsMHLw5EaxPBZwmEASjjEw/zX37zA977rl7LaYTSk
rBYXtTibAP/cFs4lupNhqvmiNjx58Le1NpqMwkqQzjhcddIYcEvsutLbgGgjt8jN
tuGwaOFD7YJIUk9kAvJzz/I9V7oaMcqjdk9PQSxpMPWa3qJuIgEuNnbASX5qDF43
ljKVIrwqfDVDiA4YkebOLEcSJgedeVWlFT2r2LtDT7l+0VRSCDt3Hhm9C3kQqW7M
4kMpQDVgJI/uZRNGGcwqb07CQNpORnGGJMQ7tk017Pn7Z2gK1Th9+NvmRm6mLaPr
vVxTEkm5RXvJwWXHDJ0qn5vZOICHIvXsvRxSuqVMYchRRNhmTOIJITVCdQnthtmT
6/XcuVcZOnJklMF5oi4YnXRUAGkyMJun0GiRX06y8/sELKJoRFo7wkWq832odJ6k
RHBhBPFGltItghVQ7VXVfbeNbQTY5mKn1PCMv+Uw6+71OJ9XW7hY6yKZxPboKEYZ
WpKjn2cG7El32WsBd7sNYI+hcFQ1zKvbTxPMu9JuMkQhanOBJb4OSlRc0kcFmjDM
RO/VHJnOi6LUgYkphufkSSlcddmKrCE3jfNwFZr536el86beCsLknqwh1ip/lcel
L4TBQqSwogJXNi9Za7eOCUivXr8C7DJHlSKMxSEgFS+hep0hDArKB4gupXto3MLG
4ULo+QyswxU2xRHBs69+xdMq7mpqQur8DRBHjtE7c6nFVItj88jOoJdq9F2hNuVw
+iJZASe1O3MztM0L2CSbiklPiFORWuYJuvLw4Wp8HB0eTNYUDqvfEWTCVDzGws2Y
ogup0v6hGDlBQCc2G/+65Lgisb+3Uqw17MhogQVVduPxg4zF50j2vNMFtFy6Tw/r
5UdINyd1B1g7qKwHKJqJnhNrqzzQteD/DSgMLUEJdQZn1XNTNYRlRcFQL9yUiS6a
Wz2dUhYdg/9sU0kx8vT3Xr8x/Bj1t2wtP9FtwqoVA3JP2rDArh9we6CVXeFw13oG
p+is83bBQFUUx6vaDc/zwX8D5fs5bNA1HzFwkNs+RqpV3dhYQmdoK3l1dhpk+Dek
ei4G5NPGiTd68AExSv9oKVXN6vi/YfAoYcenPVgIYWrPo1yq631bXdIIQBLO99Oi
XceQ0Y25VSb9SmLMtlBTyEPV4lVMhYdUgR4IrIksMfa3YEWkfXwdh5q5Z/6G2Mgy
jUgbZGiKW23VTvAAUbDjEwfa0qx7QnqJ3IJ6gnoQOMQb0p6k4CzCIuuTSAuk6N5p
MLP39xrmvwCH7ghN0g2YZMm421xNDU2JCKvkHvU5FiiDYLtD5WiS+DdDqwIOh7kU
be17fYYdc/hpMcX5ShYHyXjqyh3AjKHx5a7PDmIYeE6syUrUXOwxLdhRjBbrfbeU
+IHQpS8PreHvx5TauVOUfEgXU3nbovEo62l7ScN5/xxb3S+z83Pb8NAX0WMHbHu8
UqvN7QzBtB2IPFsyDFE3lWc6gFN9U3Xj6QZtW/z/QMNqarILNzibt4gdneyuSJeO
W9YHSyPHv/+8SphB1je1hGu8lwGmGmDVDeqdZbW/77LuE+8NUByXjFEjva2wjeD4
7Yi8rdwGO6XQAVDrpnbIwd+/PpirVA3OUUJ5T76ghSy17lESQ7mWEH+QXcPJxEu1
EOePOd7yiyJKlZZi/KN4bdABpFT3Wcd8PAZaYwtzokq5bD3f7RLcDqF/0Ht4SJqC
WNOCD2ehSNBkHmYWdfwMBO4zh4fRbCa3mc1Ad7DUphM1qlRCiRnOMyu8h4g3qnQJ
RugPsA7YlyGTCeVJGS+QZvyYLD5ZwZblKbgHJWB9wI2P6b8kA6SBoDd+8YONXMaH
Ud+72GhdA7ReIDLIYd0/sIIPU2BZRPEhtlZVRI8DZEE0DkzUlWbxcsbPJcCxnYe0
wix76aUmTVuCfTxDQrtKmFDBgXA81a5j0jJIK+3qi+CwCJYCEPHD0TdluMjxF3xL
eC9yUhoPJ2Kw2bHPfK+a30VxvFjpZi83ISyrCm41vYiCHrIMC/cjUSI3A2qcYgc7
baXL8sXc6V8UJFEzR5Mwnf2JOZgmUtcCmotcsXtgYUGDylOZ483TvCRc3/u7NfjU
bT6dSptnMDhUiaH5PAiLacxqFZpPGMflnejbQQCxQAxSLfXJlW8pddg1eCetoF8l
E0Lf1cJsOLDv3/RkxSiWLK7OA53SGkMoRE7kh2GfTLPNs/3LqtwOgeliQ8eQLsy2
zfbj/0SI2wId9B99RAH6uQrsQ/dNk97VKACOCYtntgGd5D9fWoaztiYEHdPh5zuN
BMXljdgArTyhInOi2+uGWf0nVveYu2qrmt5qLW1wM4P3DfCc24BlcMRtmngiUEvF
ZvVqGJcsLmqXi+/iHfioptiHvwiRRsdx6dxP1e5mRCfVcu9W87wNpP3WpYCcyKbh
URZa+dlcd+g3vOhqrWoCPOSWoFsapd2W5Y1767Ufzp8jGEzh2AP+u+WYUFVt8OD4
EWyI01QIugMNxaZA7XBA2fg2uITpJENF1Yto8MQs2ujPctDgERQHVjZJodYNAeYg
5l+gDk8e1G9njmuvCXAJHxbyCw8xXJNl6svc2TdP3jeU5Kox5hbfLZLYNG/kRuxS
TRHj4s8/OqHw4MyzHfmuOp4tNOlxZl6q3QIRZIl+VvJrNbthVfeOcFKJdXMzHgKc
njzwRgvrMUbMjLgqWoCBBET4FFhu1DMdN1g9e4qbSFszZgt2SdGbUxkEgyK1NmPa
Sbz+mt2/uHP9FFaSz3Nvkn8R9bsmWH3IcuOtU3TCyb+FWy6DRsKpqXoZJC5ivDDQ
qOQG8iWQ9/QFPdJlh9OuZQBcE1fuoK4O1LYuyjx0TFY00GI5AkJfWqgneNVuaU4s
pwFNhDY8ZKdGsx0W2Gpb42aAgR4ofm0CSSkzi9wA1SxJEJjB0ekYiyBRGrkNm/Xg
5vwndqCxd3MSDWnep/NoCnfnpMjdfCaImqAGJnoL4JuVcHMydyhXtIRME8dpCc8n
gGAowaHgQP5eloOnTQYlQejrLYrft7R4g0Yp1Gu1LhrgQd+lNDixxfExOil9dLDU
1usvy9mWYy78+SPmABmDp1x2dJ5E0XaEqqfRLxIMLFoOx84UN2EGkqZH2PlrsuWn
irnxo1ICKLhPLVobh0/A9xsFpdCBzH0vvX8j/8TU4xzCkkKt1XJdPPMCb5QSmntE
s0JuD5b3rh5xs+WqA+urATmbK/1uwrs6mJN9+kOskU+FPibdV5p7q18AXen0IekH
02DHmuC6S69k80JJBenG0GeOglWJQAZYgLCzTFRhyYiDJ3rmB/MyzsI57lrj6UBA
xctmuaYRFLvaQx8fr80E1tuNT0NLYaheX68nit5XBxbcCLPzBvv6FeDPrJvNuRe+
WUOgWq9V8XNm4Mnt/51fzA+970Z65w90DQ6u7WSqhd8CfdIhe7hqAAcTnb+gRggj
DndxDBntSkf8o+FYM0Qo9fdiUzQbz5XDyL0JNZnHIeQ1x9mTqm9nFDS2aSjV5uq7
LVhp9odYbjQQNS9DcktaXZmnoXIyp8zhepvvVpBVd3a/G4xdBWC7GYF80MDgqCft
201xrPF0jfdq0KLmOEjlsyF8UrB7/BK/Bk98cBMg+qq5YGnHJKyjhwxNrSJrHIpu
NTjobxxSQDMBbi9021HMKyW3kvKFgyACVquMqVrdtAFmW6Ak3BW4cJ21nRSOYv/x
Mm/BwMUcYQZ1hK3R/fB9bfU0TTzaf1vEjKKPew4QK1q+bCUPJaYYNLWm8OzsB6+4
Un4wktRJZyszMUzBvGXzlIYe07ssJ3xgsD93fllrDoFvvRl7rB6IcyRmMg0Vjm+4
FnONVNSRDj0BPBsjXSsI4dUKWnwDAJ5Tcl2kSyUIZmwkj/b4KzJvPBDj9nftWE1+
bPHN3F+i9TERfM+8Y+9oGbiqUVv4CH+MxSnfkohoMeFDUapbmuCn6NRBdTTgtHr0
NB+ghWnkrky+J7zild9kDu4Xs6LYF4JHuKkhU/idt6/YK+YF7DbxjFnvLvG73uYO
CRVCfx89UvxXpQ+mHLrIpiMPxmAgWu4DcRV09jCwwgLmlTIRz6TcFm93wlw2PFtA
d2lyTf0IUemjVFcZfbNJ6BFxgoAjNE5mZYhg4LUNZACLsigkWaA7CyNjMlxKW2CN
M6dhXpfd1cDugUlecxq1TU+aqF7c4pSwuhN5B2SF6naHF7cqjyq0tIz/7Zpl7NCq
zwkuyz51y8pSyMdMUKRnh8SHDu7mVpUcUobKtR9lzLtHVaIbjado9pkrR1DLogIr
auoBpz7aRqT/zopCVYjmQlZz3w12F1DA8nYhNASYHi12v+aui5d1JHynn1u2F4Fp
nuhQNNjMrsJBWamxmxALvVQuiS8/TyWZVasXisW6kQhp0/pnloXMx2hN9ma6nqGb
3T+NqO/fpfehJukQLy+XeE5y1JRGreA05V1XpJQNVbh32ZOAYTPCg0O0MciAspsA
+y9BsL3un9SsUHNz0ga5ZjH43VcyMIj4M1IuMyLLErA/SA5UHZEikGCcDABRKnaG
cRpmtzSNtODZVpR201Y8WsSuD1ZvXDPPSbyNKz7DUmKW4JW94epP1Ok66O9BDVH9
pblmwdm2AQqaVrabxEMgxLAnuQfMcVWfghTFDqPvJjsV0GZ8OVWWfZ9W3kSztl7T
PBhLWhLZfUtWlCNF7vvZY/hxml7waq/UmbautThEFYsIMV5+Dtfj7I4xIRBJzFBq
tNT+Pfb6uBsl2Fj9AwrGt9tS52qGqe9L6Yla3htePOuLId37719PJ4t1ZCSGNHxp
7Qc49UikcGSx6xT4vHypBbFBDHxc06/r6Sh56mRg7MhGAPDwWfh4Vujf2Ai7amR8
BkFX27Hp8iiMGX+63OjcVwLekSjMvmaIPFTwwIJFJscX+KhlVzl8L98PhMKgGozA
jXvjTzoetv2+WcB5fFn13+o8LA+BnoehEqEgKoZzPknDubhmRAY96NGgSXV8BqoY
raqonx3LjAiVGY2i2yS/j6WzsvMe+4WZqPeOWONIHIz2suqDaYt9FM6loTuXM6pN
dgC1MmS6oDP+w85b1vQmgFrCb7Ir6cpcwj+XcFog86abnXMPZc1Wk+5Gs7jAXyDY
Jr3Nchf0hun9REJORs4LgKXI3S1vk5kqJs9ITznQy56ib+U4o4Todo2yEiHPclzo
JKoJj9ktLVNO1PCNak6w3omS9saVX7NBxZVwbxvJ72kak0PTZVOjj7DCS6q/O9Ip
wGx1Jm2Q3BbiPH3LjiuBTzEWkKag4rOnwatNnlJGBWUei61CkSiQUaTf51syIk2T
pLcJKXHCR6AC1srJqqqh7q8SBrIDl5K3tapI5BKeEPUw7BBjHVz9K3sUDLtNf14l
hHWN4RdYryN+cphTh0A9Vmq7rEBCywfaJf+n+P8yLwIBhJYfneziMgFk9/QET7Hk
vsaYEX/8egMOy/ddjLwXHIwSuITwOsLnDOtpia1J6GpjpOVdLhspIUHOQuQEgVsB
uqpEP5Z7DtQSTZxGl7IAKSJuyAMkfEXX9GspeWpv8N2uss+S1dCIgQU0yBaEtFL+
FQc5dBuKjqhULV0uzbqAi9+Z52apZjnRSosd2izmEQuLzdZ+1OrPViE9vlfFSwc4
QCwILS9o43lrYy++cX1o0s+ITHcCBMC+ml/nPDWYH6BxXQFF/NuM3RTeGuyYTZfV
mHr4ITYjBH6Dm2oHOO0PCUjlLfTYDK+s4XZrdrKM4gb0Sh7JN3Wn424PvhQhVOPa
5E9Ua9JLoDq/uEZXuNw33Ra2t8yUmNJyFYHOLxH13mTyew2xAHsc738ETwtYb/UQ
BH10aGfgzrAy//tzBohzRzVMiJ8CK22U1RelXpGrv0xnHHZDoacZO24AIWtlYwF2
70//sCIwq5RVwynZo1N2d6JpBeyU/zxl8vF+BhslgZje+LBW2lWt+biJYsEZ86PL
WqpnM/Rrde6OsGs8c6N5ll1BtIFcJFZSQBcZAFk6atOcReQ51P9Xyx+dItVigqRq
8tVfmJXThXRFWTKsa4bLHvTwybwA1zC3JA/WS2bu1p0fpY/bUZUxSy6uYFDItswP
PZPg5gKWcZsh6GZzIxG0+xgicKmvL71308EDn1bRXbC5V5mkHz2exDpROnGL0CEv
OPlNq3Pbk4jV6179DbSQ90R/zrZ4oE0Dx/Z8QV+Mh7mSM97N997HZ4lJUE7rA8jT
4u1EsxK+qnPiZQGus00jM1yQltae5oYuS2b42x0GRi88yjoQjKfTJXlOE+UNiuAS
xtmRxo1LUNLuuIK/CNR2c81J4faJv+c96ya4eStHpW8ru4JQuV1SkNsBQ5ryawsj
FvzOTOXoRrMGGx8mmrqr+sjjF9SEFlerRnr/9DWvuf+XiGX/xi43c1oQJkZoESHw
NEV6e3QvqNyVsyBAZXtIyC+JApWAFpLr3k/5SsBrU5+wBeGSXMbGJNRyUkF8ebqd
JJ1Qt1YSeQ02oNPlArcBuQ9MHeFM2uUX8/wdENWuAL70KgIf+Lks/e0EXQjuLdTC
eWpoOP8rqSCN0+5HfZOhskjVkujbcQKalhtKv9CSvdekOh8G4n+64h5WzFibMt8H
J7ZaKGVjjzNHYr3OjVGPpCiOjHN5GIX48My8HEffIllKry8jDGwCRlsNF1LLIlKf
cEER0GCteH7TlX/uk0swNu8a8myB+Tdczq4lms8wI4nE31aqKs57vFkoJv6v3CaN
5XfTpo5Vu+oJW4PdidCqu2qV0wplnzA7L20xSH5x6oFMkEwU2aQrYgTEhhEp3rTB
WpRgTgRa4Dsd5e0tJDhQzzQK30hUBkB5EuYN+Xep5vPcyEZu4EJ82bXqXDGaTwfG
X3eXQghbH8Of7oDjzDI3fXWVUQh1LXKh9qQhfLSHov1LwQVIzxAc1b2+ogikBBMw
XNBjsujVnAAth4GihJippc73G/XU0BtI47OTgt3Sxy2EoyO4D0IMHSRx5LxhA8tE
PIwBbKQEXDbCTZq0fWR0xd7AAuRgQBtQ7ha5I9LjbtKvWkHEIk+EI2i4irQsny9j
Jj+MsTLAwaUgRt1Jce9th9yFW5kaAp3zyfhSM8+QveCedOhK11dqhZVzRU8aUUfU
2Fh3zLu1jlbOftYVXDtUkDa12R2iEeWpvGvvX/kHyst9eFwP9CXvvwCXTc6kZdm5
Zpy3OsPU8acX9FUA/Jz7G7rv9Tdri2F1mjDd1ds/smdF6p6Ml52aenFQIo1wc7tU
siW4l7qbKK6J2qAYESnywuNvhyZcX5TLjD95Z/kSlAJw4lV9adq1htSL2WCG9cCs
X+hp0QlO2ZNRdtoUfrBk6sJU0pZJMFrM2qBnkJ3SfZRgGHinpY7LTX2Pz1GARmlw
jyakpG2UwnLboNMTXInwk6PvWcs7Hd5s7RzH6zCjW07txyrbCZnB8PPac/qyKhm2
Wpa+Hu1/3/U/a7SH+hJQZuPJkoJJJg4p7QsxuEQVDji95HeBsgeG1/Eir8q35ghu
cJnon/Ylkdt+ED9I3mXoeuvb/LYz50d1HSb2HaXcHqMADHkUwu9enBaYDD2muXXQ
RYZt4Uo7zbL+uqzTqpOBq40JGLAwTDPBP/U8y9UKJBsR+r2O/wQURua5nFOFBvi1
+6IrAPywW5Ik1w2+YFUEjVpISE4yv8GMcQWSpJi55ahli4VKBvnYHyoTACnFsna1
dz9yVGNKCvwLQVTNyGYVBkk6t0XSGGm18J3QqSoQeidPJqTeUYTD6Af0X6wOGxsj
h7m2l4MDWguXkQf3LA9/yKueMUqkNmK4IX7HzX5rZgtAkfgjFSbCZhrKlfoSttah
lnTBHt4GCzHLfbXvj0OaOnyn/P4ty5aA80B93tUlguKo1mxpGQ+mME616y1+xnDF
M5aBiapYPCpN5UuxQbrF4GEz8jtQtyVgfkBXt/0AqqRFjB6l3ClNW5UFoTwKJXl6
VCFn2xcOIfU5EVQ8p3b5CqOQjXsVorP574Qla5bsQZW5IKVwmL6VvdRTru2VZQL9
YrvXcf17i8syVvrDwr4YPYjBtnzWVGZPHqKKhQyYPsvPZLe4sYs4MAu2iRxxs/SP
1WLPMjMxN9+GJ6Q08fCSLgS8tO9ZWYmwWVUNNWOG2tIil95zmc3n5kJjep5M18dE
2FsaLW4uJix34kjM2A6+oeRuwzc1mWVs0knmHx4CVI+e4Vj7LNjnyJgVv4Z/i64B
uA71+PbQcYqwnMTlfycfOUpZty/qXqhR8+lkkukLfwcYhViOYh71g4ZpssDaCVeG
jhkG404LGA9QQGFEZjctz7eJME9TPQnRFAM8egsRYwKiHaGlg4GJuHiSm3Rnr9Az
LUGR4i1CZdwXNcihIv/PPlOv9gT1Cx7ZqfMCHeqVi06Q6U6BfTcZ2kxY9IOYaATm
QlvVR71LtskPa1UsxCJm3QFx6CeR0ss58BwJlC0So6VQI50n367kBsAXbCiwpt1L
dVfs5ZPHpH8AcwnHm0QVQjxoseAKQV/sJJ8+Amm7vlGGkszZQyk0FSv4JZ6Yl7Cd
aB52Jls+sFEDVuq92jrykpSchqfi/lSt4pmAcd6huaLcGf4kFI2D1u6GmRQCJc8c
ORtO8ZLtRvmM8iTOrmZBAZpi62n6sbTxao8XhdH0MY2ibSM/QrUsnC0Xf9XSATch
T8W4rLHDqD+qPliAiOMrKqyL5swO9F6F4xofu3MX8E6lO8JTSTaDoq4ee3p/kZN2
A5a7NrKYWKX3F7o61J0PPQRAIX4B6uxz/0dgszp8ODyFofFPGrzM/jOEMg5g0TSZ
U+8hu2godRwno3xxRpHcwNVaDwz3MfC/d/WYNhAagBPWEnI2pMEgUY+5tSXJgYwg
/P8A4EYkCkol8s1n4mPnzNuZNHZ2Rf4illQWG9QXxUBJfOR6yAdUIAsbon1qyTvz
i2HNFt/fCF9Yg9wUbLN3AqvzDtNRwp9Wh/nnekoZpS2HP8RKMV9HDW9doeJUCesJ
q6SBkisFWWfQX3BdLEMt390vUtsSNeW2EGLJVONMQsxjForF3qAB0XLCCGBPlghn
Lq/n5WW0nW3uqrt6oHivUJbDDA2hD7bdvRBhqnwA9qHogSi5AOKP/qfbXzz27Nqi
VmTGSGDJxpFY6ee1Tl1myW0FR5B1Lqs5qEKozLvrX3NTEuJ57n8IWgLdj7ifJjl1
WN5JVYsMfpD666aG76UCJD9FInhH9LOvQ24h3Vd6XuXI0wOV+d2QQdVJBcGJWvap
Litk15VH20SdzUWyAVpjjVFNRJS/L9M3ZDluZCrUVaVEmPNtnMIqOnoZuuLXlpQB
GNj7BqkeoSzz8SEmA2V5GnclH+7Jbym1vfbqw8v7OFb8JsQiwHpAdYWbAtTywOIi
JgP4gTtY35dpVUB2BmJvhPkk6vV6cXtIvl9eWxfCk6IOJ6Hl7Y64JyUQBSH8H6KF
PlegwI/MNrBTkXUQNBlAI1dOb1aNZUFZIT/FPU160iyJUoarUdGVxXZQrfrxIPAr
xHrF1gQGHqwj5j15y0a8Bu8AiDbmRAAa0G73Y2O+pnYqeMr0tHHsmZUu4Ybe3iMa
7jcugNCLHfiGYgwx00ZgBK8+PEl8yiDr6lLPKKmo+EN2iQd/8jKDuta2qZ0utzO1
FPuAByR/hDYmple6gIZUSp3q7W11JVMnz4edzrJx1UT7FQqyA3BwOCQ6YhCA+UkC
LGREjOL5TP6IqdMAoEffu6A40oxeI4Hs+nuBwTmXw+5HZjbZlAK3I6SxiKq+sUe/
qk1mTTrz75/ynT/sPLDQMmc3bLcl6g8YwqWlzk0N33aHVdBMafTLGBbDJCHCc+V9
RXSjzyXIhnhvhEnDjXORkSmqwIkgDPp6UE/w6cVi6fmuH86IifaZQxmMvHOr1AZg
DP9hMtFPomV1iLsTB/GN0NXtGhZA/KuaibljtICHOXpSY65oX7BTGpRq7A+ePocP
B9qLbdUTh/PD9ull49HPTR5CTOzITtDL6MubGAx4Ih6xumoyTJRP8WrChygtUGGz
tyLEX7pfDwiG8dXF36bR/V80nxM6HgqCzEclIiVHew0vhkE2EdOkl+MrTrE5QDM8
HLZSpP3M2vseuqRP8eQuQaX4vmG+CUiVg21XsNc7ObhjAzynnQNDnjnxhm7ugkue
VP+B9kGiYpLiS7GHaq0AhYZx059wjR2SEWeleTQBW3qokLcKi9PznnK3GejtJYyQ
k+6hnxRFhQyRts91+J0I7MNlaGy0+iO1TgzFHM4FimWTBeTXAv9xemJ10ZOFhFwk
74rH8dIHpHqsXAJ9J2Rb4ZPkKTgZ6tL9aMLOCdte2YhSGfQNieo7f2zhYfz5STT/
TxExkXGjkn+KUDfbe0oNidj/l5qX+abQ/YMVZppfaYUSIBqGQevipvnzPH0sF9vE
hcI+SXApxoG6/CWuqCa9WR5FgE2LgKVIbJnSSa4VozcTNNXMYXuVkLVklaYggSP6
J4k9YBVXiqejrSFM+iXH03P/XwkDjx7AyCrjkAfVF+tTKLmjeV66mDTOktYXm/VY
OLMRIApImt+cwIBAUMwH7JzXXEuMWsxzjmoZHzplgO+8e6mtDxx04KawbyLf6jor
7jL6St4+8hxYpE8mLbtH/f9377MBGmv9mTbaw/2Gna1WD0chtTWJzROpcDcqmH5C
94FQ1EJhRYugEBDl2dDjL/xWhTm8jHhvIH+qEkCJ7NlrG/iH1jkWOlwB2w00BpfL
84kVpdEI8QQFScc/k//TwtjA5HUF42Ux+0UG3iHkzzfXzWKqyuCXTt4ssRMvl3qv
kxGNc7nNNjYcKZ6IgFEGNrlx3WMlu50U8np/KGm/hnifd8zNSgh5/0yFfvbjlGjE
p43isXYEHr2EAC91p5UMWagq2jqCiPKv8+jX6zKUXP1Loh4Wtg/m7l8SO+iIf8eb
NNEIvb/2zm6/jVSBSJPjDMMHxLrSObc4Csq0dWY1xJ98PMrssf+BbQYqMvsazIs8
yq8mJQlQ1dnXIoA3LCqDtexO978jn5RjpG71al6OCMrUlDo76fE9TbFhaOGAwzCs
T+k5l0qBRZpI7UwbB+387hNk50OT5jZFzmiRHZg13QZ5AkhwurjE+7NtUs/pdgod
lVzsqg3HTNQ2FA1qzlvr9CrWIJ9rawDailPN3mgZ5re0H3g/lbNyD7ji9sMuJNp4
rPa/HCnbeHyFw/v//aCC5HHXXDMFrxHvFy6HpWaMjJq8hGYk+COLuwa9gnydpmvQ
P3EMMV+9+24hw9yrYeG2hlW+jfmWVSdoNxs78ZWodfWjJvmT9Cn8HPcJqzC31OsM
ciVdsFHAQZDKqlGWnD90N6djDbQejGcTpjl4Eeulb1nRkkVldTOqekkpaoefTVVo
0GNHUItyfoNn0I5rP96JmM+1ZMDZ8Da2A+oKlpjZX7VSYKbVi9KPhgQVhlApIKRH
+cHWmON6zW1wHsQLJX5mGscMc4guorQlYHkmte1+KqkUTa0ixlnBrvkYt/f/TJUh
fZ1h3TSRRmPc2G00+wz19tcY0FhirWNgw61n2twv7tdfP/xD9H2UD7o9dnmBCIKG
oKXbg2vOqGvVosi/URIL9Sm3W9XtHXRcn9ECfwjQ5/0uCxVVgVtGY9jrB6XbbaRX
Ww5DOru926hTPkvv8x2B8f8jusJzkqn47UoMW62lKXqalUwoimvzO/cBUfnQKwCn
ssG2Sc9KonmxIUzdc+2PI2sCb/9+EU4xsO92bny95bqwD1Y0/Ih/+elaABZjoPGg
try9fyfy/b+MfYiNT8G3/baoxUiwDBkMo2qSzJDMSx4vk4A0jS7D+jFoRsd0URo1
g5Y4X26GfjjPFt/eOgD19xBSJQj1/V2DNjcx054NhUbqNiycNILxrCJ1hqMU279E
tOny7+5qhrZ+rD/+dI4OAz1pYHGo2/mfZog7eyI8Rf3NGgKtEOpXo40yLmsAGaJS
zFPtlDasBgIuctlYB0AnUEuVk7BTMJW68PDcnCjQa6mvrov+kdgAPzXu2vthV5TS
cHJlAi927PF7oM6ws7lDi9BgWR8tV11zrrgdRw6nHR0hwuX7ct7A1ZjLNRWFJVP3
ugnUpzTwOjYHcR/INgpdGtLqHJgp3C6q6Zs6sa9DkeFImleqZhBFb/pEk91lnL2d
bUht48b9CBmQOc4N//HMc+na54CpaQHpyUKSnpN/0KiozlGjRoaOBkQt+yjMu+O2
IfIzsRzeYgkIrB3Si2b/Jzsl4iKYZ0wlPCRT9bnYtSiaykRyQYcCQmh4HjLx28Zx
vNnozQF0Z1opKt1kjYDgfsP66Zkp8qod7QNTjJfy8hZqiJhorgOV4sVhtIsYq1YK
vlQXn8s/J99fHoGuHS7vNEiH4yCDgLlIlaghR171Ic35n3yVgZDzhHkvdntvf8Zr
sJkpeMgR24ecdCy/HIaW6c5oXZzMPZ9p1EMrsv8W4JQEz+cuk76VMq9HErUAT0lS
aTkBX91u/gW/kevyEuky5umMHld2gDJKFuuRrqQtaRvGN9zbv5Qx0REgD5uwO9Pq
6N5PTPgaue+tKLMy+keS/F9cbrVWes69ohqNSYgwREY2nvfQXzdr6rUFdBraZFUf
r2YgPSQUBP8t97uEmVdZ2m6sjJA7qAiWibjzcscuCjS+ZcwdhGJK9gP78XI1Tkwn
w2dXqATfyTkLXnCgBJIYx7Uu9bSaPNvh+djS75SyBt1cDYoHri8GDXnUFVn3rvt1
9kgWo9kQqVYHeR8NpjUfQ1Hnc/bYpGu398G3BFtDnpQGuaoPMRLJ91THrUgcqeTI
nzQUYn3e3boaYMzotw7r/SNunp0ythHY1X2LG/pHTgbDa0yxzYXQPD8xw4YzvumK
EI9tc6f54JkbabMqCj2w/fkiEF0VRQgcfeoMawfAASnrzyuBti5aeioyM7LRO9Zb
H6rQD2JTwDEqq+GXLE+Db8Fn546FWUEHPGbo/U2q+ci2QK/r6Z9EQNpIxPBnenfb
0SNTavhhXDzcKyxX0Xk7CDcpoOlYRbHugyjDaCcaYxcYDG4kQWUBCVD9a8a3X+RP
WqPCDBA4S5rf3nvYUljYLHi8xA9KmVcSRnOHJ1ihThFEgQ/OWbiXVjuJM6m6papp
eoZad0nYV1AQPTcyQRdl2LXMIyQV2mQmiU1NqheaoIhRmvZB0VEUOnR1tanJC1HW
TIbb/6gp/SqaEUxJtYBZMDeXQpoIzR2rn09V7sqdngUOXKB4vk4xWAPHdvW/o7OW
Vce9PPL9o+g6YKVFEGXvuj5T7uISvERkQLTgnHKmWjdURd3ZKq89b4AcjvnLoDl0
yjaarCQmODs2p3WMTCG0EgC21QaoH8kRmVWGuyn+Kq1xCifraQ9m08s2RQhN5V+p
vpnf+ksdordwGRjafIjXJpQwyse1KeR4n4S6YypqUIA8tqs0b3WM6gJxKgZJnyG6
2pcWR1WYs7Mo95Oj4YxIkibI4QG1czYF/okE+sA56Cs8ZV3at8DhcCzSHoxNUIfM
xoVnCfvRCg85TwgVUU8xznJ6kWusTv/Iz7jYpHFwhFHlvWg69LKeCbiDBOr/TOTT
kvoH0zBAVAf04D1ZKrvM5Ffkyxt2djt5qwGh5KN9bqSDw3RWCL6G2fI7DTda2oic
qb8as+EQ/lMNYm5aDqq0soHQjw9YK3Fv78rkKOxIrmACJaKUWv9r3/+yw8YPScNf
2RRpgToPN8GzjRf4oBSwMYLNWh/gFt9+1Bu+8sSi7xG2NpU5krzNCCAPTImNpuzH
SIYug7RtEvil0Uwe8UYdHo332Y2y8sU188WUrbDyxxRIEBSZksaak5w/AbhQLHgf
m7Axt7YFB8QBKsHQOJ6h3heqOsOsemGeTYRlfeOhtyNTSEFV9XCsMcy28QL9k9iO
b9EwiWBsBxSD8CXZqUYKk8UHooAEqvvd8OLnumzN3S/ep9tsSxqi9p997zn3gH+2
GKcFGynzsF7GKsvzLddegxmkNd8QyUnPF87JN4FLX4KkzzASxQKLy0JNl/FIjrq9
iL6BHvvyutJ5C7F5NqObqsmtHCriQtOAc1Y+O0PWgsLkmmEbiJ8XcadVHSGO8E6h
pyrny9sHqVoz1pvVKOKfsgBizi2UGqA4dlD1Ez/soA+ChrSaAyDpV7OnrPePl86L
Cy03PQZC3TGmfrTDBS+5hikqdq1+sdCpSI/7LfXxFrACU9zOTAOpN5/KV6+AzG1p
lcI9Ho9HgJ0mOzQ/ao8yRdoECPPUu3wSZ7Skm/E/CvuMHqiDibT6ug6sGTUabPiM
fMaZHKm1QDz6sw0KznznBjz/4WrZMOzD8i0DG0VdwTuOs502JkGp+HRNgCrXIqq4
VniD4czNo4JaZ83xdYEKf5bsv3KcDtP7JYblFZ/cGMSJWPWkuPoiQCcqWCO4DN4K
dvueBJeenAem1vgFmbq+W9BtfiLRPuZ0t4NCrrBAZlZa4V3H+ofK1SL0kdXDrl0U
vGMYkYj8YTan55Ldrj//2H/7ZgmPhWp4FyvVfqgSmpWOHBxSKxPCFQ+5sBlsZKnM
6UzRfwF3UJzwpsm7MQdCDtJhE9OG8uB7qA4tH/losLwLBe1+i2k7maNLDoBo6HoH
5FEHyQ2jboQJJ/l/OIsbDLLpLi3RVqLca9ci7HZy807Lzl7+PdmuP7Mdx5z8SlG1
nbkkvxScNN3NY2uSZcTiVUz50P7je+/7YIK/PukXtkWfVbGDD2wmYHvhK8kj9peo
xWd546iyjJbTRpYwVg+/p4JMtTOrD4LEnqQcZP/z5cAXH1ocDupKZ1i1w1qB0OVx
1BjeMjv+bGfmoCvp4qqvii+Ww9jYxuBRUer+Vxr2itYEk5OFsiB0+6fBF2tTgsvn
zjVwW6xcPB7ZtpkiokQK+Q45FxaZ8NjfJF2sOXZAmvZsf9cluO+lED71cIzQlNys
4UprCcn/xZ5veO98zDOr32ggPQIpvrCbMq7neEdgEsjsTl/yo72WN7j+P/uxG9QW
emQ58dLFoLmoHLGPBe/QB4KIMiJqdZp0gay0GkI7k24TkoVKXNU3Zyq8wv6NKr3m
LO+qfVwaLZJrFFsQCMcQLtzxuyObvXDhZ12yrr6wEQ6tjz4PNVBrmdHGBBwoAJnE
KaorYp2xRFLn6D9Yo+UUoeijObuIyS+W0QqSp7D3cFXUJrG9nYMlax3MiTVN4O9P
lZL2h2WxHLM6KqN4mML4iG3GZaPoA+4qA5J+QRsuo3o1Gv3EyaQrAqCXRm3aaBlu
GfiIjFlneLVcrTCln37zAetvkrX4k4GhMhamxD5PZwSutaBgPcdYql9B6VREPZIA
zAK5AE28sfq7Sm/LnNk0WfMCCfDDyy4qxXynaKW1SDX/3Uv9R261pzrin7LHqXuw
xdEhvTYH2hiRoFM0CiodvEga2MFBKo1SYcWMVPzh/J/dhciqF64hcaXpZ/J3jIJw
2Rz1VDG5lyZMv99tMdYHIbhkH0vuUUQGMykpCYhAF9+SkZvsi9oah/fI+Cq2V6VV
HRYexeX8/mia3xTDM0eREek10cBEWLQ2lc2VMePf68RbpHF9S0HNvAkH2djmn0hL
5HCp5I1+EoOI5ose6faFCYmRaCjaAe07EQ69a/owG4mDyBHRi3fgv3yDnSLSrK4x
Z2LEqQL6iq0CJpbUdYr0BwmXdzgyM2H4WAsrSlUbYNZdOIo6g1SYb1iuWB5HexRm
RSMG0UOrB2tR0SoslpB+SlHukogc6OR+l0dTEF974XFB96HQtA4jmfIx4h20t/I1
jn3S6g9xehvRkdnK0zYuXUJ2nkpUM47ShvibLCvKSOgEFS6RN2jxdIvGjXng5CrK
efiN/RfKZ6TmqzlVGs2wvszU46msdw9poqrqX7yw+4o6Sb1ihWK/iUouOjkc01cM
0jTscwhze/ahBRTXVnarkrLCPG64C4i7/+k6NXLQjKRgb/+dv7eNse6gX8jZ/rpg
tJvgzrVrsCcuGpVSpK6klwqOd397TmNn6kq9LBRAf4sF63V4l0G1fWbfWaGKkytm
SEWpkwl95NCm1KXQAl+vAUcM0jsi5knxu4kvwesSM64VYp9qMmSBNQBOMvy7r8UJ
0REbfcmDedt17EBhtfI5wgin+YUcxL9t8fMg/Yrlt6AZntoz0SZA1eGSZiKA6rfU
1lHLJ0q+pWRSfNwwGo4/G0D7t+GEoEiYL96032ziAS/yZ+uWNCXdfkwWoPZ1+ouC
s1FZvZMU+X+rT8/Krh04ilJJsMltpaS4ex+3XBr03opO/n5TNFca72RtpN8Kr3Y9
7Xy2ZSLmfP4ezTMAAyKb2DUgJezgNOiGT8aW5rl7qWQ5SdBRYkZtICPrtN5mdCkL
1wdq9XJGip+y8TkOZ+3ow8RNzE1nE25APlDBd3X+Zp97MttRMAoAOvjQMIoBjm4i
wbC0QKtV1CmBCImS1Awkfhv63tmcXfj8pXwO4Pl2rnDpceSuuUa3TnI2r5KUt5Pk
rYnaZfXzI5k70LICYBhW8uYCOSpI18Qv3tcJcmcHM5yCgNiaj0wJs6NSVIcJLtI6
UTziM476j6H7EVS1lxpY4sGBYFRmSSljimXomZiyTzJi3UgzZhmmmECPOJARVb35
+G4eSTY6Eg3+HVrC9DGtnBsN+BIJidYZiEQvwdIxstTFlwQMj3/5eZHjCsvBeEPF
fHtsuMM183xKDC/jyrgORklUUOFFtxd7KBigd4xSRfRsI1ioxgXmpRzRzwyZ9hWZ
EjsNDLbxxqPiR6fHaElGa7MGKvEWvIrNj31/lwhFFVQv5Xry4TiqMpc7UQAhkrlW
hZaOpn7A3RraXdjPp6CSftvmXchCizZ87HBW//QkmtW1OTzz+3UiTtAvvzAlkhKm
AKsPm9elmPJg17mVpOXBsUiJQ5nrzZ0Nkvfrr67rHMlwizaWM8HJwzFusy1Hm4fF
Hhr/QN/XEyJW2CCzI72m7m1K2/wXcy1zh8bIndw8maiHq0qBaxsSherY6sgCLxa3
N/UYN9CG21V68hnJHK8bFeZK0IjIC7ElXWk/lc2eP17NxMaJBeoIHbGkpNxXLVg5
ZD77qHbnjnO8KyrPP0BZ6O5psseZ38tMun4ZkDGe0fBlA2l8Q4pBzvtoK2Ntwuog
MEhLFD5J6q9ab42K62p04vUcv9WmggDwqb30Q1kLQGPJbeA2tuTs3pU9R+OH3f7+
OIC+AKTqmUtM013aD4q9pyPzdkPyy1x/HwLYLRuptkcFrLJP9H//zOKwnJTHjPUc
gx3DmUaraRJuAQTGypNwWm5dVkZqbfBjaX0w2EUZQLtY3Oywda2d0zD/i3SMZCER
oX3AZrl6fjpw6CaT4e8RHpDadCcv2FiJqmow/FAhc2rGeiSmMhrfvWOC1da0DTzG
uvqSx8uNWCFxIcMQYDEzLgfAJ/nvuWjyO5y5zkwF6GNV/4SrcPyN9/zHjX4qEk4B
6MbWWVi6WmGKgpSGq0k9TIP8L8TYKYE6/8QiStAQElW+QeHBTkYzMuAEYlsrXBqc
gjtoOMOAOk9pRWuEIPBRHRLq7q13HYIsKLgfjYY1dr31z1F528laeGVuqWOsfojw
cUjL7B3F8s7aBnlM9z08TLf1rlyJCtnGBiADOov2hbr1CzYWg24PX7NvRCypF0Zg
oVErWiSbASQ2JZ2ac5RejmQex3mE/RPsBQOilzvbu8VoR9EqKXS6VhoWbQ4QIxAz
HuQ0nOan/y6oSNeEw5OqVsRJmWiZg4gwM5Mu1MzfYvWyS/orGR9Pr9Iy5+lshRIx
dN36DmleVmvKXwdsVHqpERnly7rKfhOx/cJ4TKWseBnjev27EjTtUhYtFrGi13Pe
X78rvtDGNDOKFf5FRmj8mmdFRsqCLAik/pgAbwaObLtxRcJr10VdYsC8Morl/ySh
OEjThEFCi0uWDc9zQG1iNcHJMFHJ6ykGLJ7qey5cf31sYIY891vIDoLCEvkyyFhG
Jfc5i1p4y9nnh6pdxxYWzDbKLY1lPvQCkYkFdxq1/lI6msNTPRdeHo40hsHpPhPA
S95SkOUctvFHehV1Irliq2IGTkOrCHHsSOyVjlOu96725Xxx0COAO2vTEdsgQ/qt
Bqbb+4yymM+wJGoAjx7HFFBl3nUvxnOEHFyj5VTxMKdt6Q6/utP2M5kT7vEeWkO0
H0kGFZ9LgjvTvREGjDona7f96b7XYPpTIN2C0JBPAj19X35A4yc54F8OJeOjTjg/
bu0GPxMZHT5q0bZ+4n0Gnbvj0y8qW+qYNpZLmzn5cGTFgzR6SC0eS2gzR7YegJL0
kq87Aq7qQ2sIiC/5AVwx+mMGhkzyHp6GLFjW7EP7ioWSJH+XfelkpopBQtjzYbuB
TEXnLincPKVTzdO/xOwOyE7HqbneWA2pv46fEHTRUvrL247dhRu0ZqZfyZ6hwtz0
/S4E6Lya/dTb4Lj3ijUQGLCnPD7yGQ8bXIy6gZ3uPyQ0MDHes/ReEjNVoRXOLnBD
k8D7hiA9qJtVwaK9jA13lvUp6+caQwk7D/1wDpkow5syMz5/wpKM14mXc+cBrPKP
Ebm6Wku/wLNo5odMX9Bu3MhWsfHLUaRZcTillF8UjT/CWocP4/78WdMFyUICrWui
BGCFqIKL+shR2oMGNtelDEDaLidg72Gjx0rw+I2Vw6t/cuKhhzLhzrD3t/sdz6HH
ebQejd1Bm0Z/HGYKrJy9z7oZqgamxq+naOfe1Jv66k4gbUx4jdWaFfPJMwCRjbEW
NCR1ag7hOHt0fVSrlfCpNOUQglkhMeDfqskVDxAetmUfsuB4N9O6VMvb/7oxarXB
8+BQFptea3Uvj9kU066mv/U1RzjbGBpqjIBbzbh7T1ENbU84FyMI4GXJp4ygSODR
+sS3A0YTekL04FZjRuc8FkrAEpEf3yHRMT4t6iXQedpPo6CpbsjlRvORgxTHISxe
WSrowc+gz4VioPD2rpowAdD851R6itxVYUxMTY6GZCtI86hLcpWN8tR2g+w/XkZ0
Rrw+I3zF/hs8lR/N1eOoIe73pn4r7J28ya3d6a3FqQ5CnoV8bOrevzwdtv7gQZfN
WKr2vmd4pnFg8zbNSj1y7l+YffGjf4bG22P45/AVRQw9hlf+zTCa3H/uXFR5+hUQ
dpQ5SzFobxyGKo4XXnhqHHhtJdpXnGHTfQ73Aijih/0AKXdRjjY1EAmCldQnQ0Qa
0x3Ajie1zIhzjHMHRZQ3FUX9VhwfA5luBQ/Au+PGAN1k1F/xK/MOtQ4cPK8/5Dyh
oyZgeyLV+O8h7KYt65ZfSdTGbwCreq7FMPvj7DCYxF6Kvo40y2IKRXAur5pdug38
/DSZ6LIWf4xth+6A6RQf0oCGvMjjf30WLywALI1BA+/J+J2UN4X6Yd0o+AUvUN/O
O/IVBSZaHXqenjjU7Cjx8daWUnCPdU80DYy5RdCWE306da6Tgy2mnRQtrrScbOv6
IUczsXwBfG9ohd/wUuMsSEirLy65sd4tzWzlsRqdjbjEbZKst2y7WQh+c8HitKku
bNfjJ+aTrNldbroSF8CzFCCVHekWu32ljGUzZ8ZwW08ztze/PDXzyMlNeVRVugLc
QLcFgJQhM7P3ZKynXH7XxFHP1RIVx9wHKDc4vfrOWW27xHU5e4Y+bOfgXB62taP5
ciB2zs/lH+xKQda9QRAoc2GJG6kYh1P9IZwTRwBwCGiPY8wl81oWHYu3KRW6W2x+
0p3kcDg8vwG1bPlkrRd++Iyxv8TSFijF8XdtVYGt1+B+8JOCRDOFMwNeOOdDkHz8
x5gSiFyAL8TwX3TnxNXbldoGVmjkykkcqQ/VbWUKuIAD2ih0mo3RIDz4Y7utPPkv
iDY6BWqj6qphKDycuYz8vC6lApPhh9siudR+BuKPI8mMv4KiP46gwXbk0OLNxckv
zcjja5TDcdWkMZYCtJX7EkUk64K2Le5EAVKWdMbG7oQMn7MBxiJdatLOW/I020rx
v0+R5BbMlvg26ss2ttSDO9FL/9bY953WmF4RqFPqH6t5G7EoyEFkuv61xRLSlfdH
50gbwOWNls3jhiiOnRbdez0lSXi+B+4fD929ceePpPGMU05rOeLvp74kJ80NsiFT
VAemI9mOZXzLzG9XHtA/u8WiSsjfz8OgcwzNf+7/XSjpsT6L/Pef2tnuDDneD/yI
k8LzF542Yqt/svc0nwSAIsaG7kbpPhCwz/I7UQRv1Bcz/FRubAM0ylh1LeqaDh5J
akZEOK9jNvSNxMFwfzX/A9o9ZKJA+IH0i4l5k+zsrjUrIoUiJu4DuBfAuFBIW3ey
3l62Q387Ukn7Iwa5MVbv3Wm+J84EBuMw8A5iJcipXmLBeAjImx/p2+pwU5oMG9dM
7Y1fnexHPz5RqBxsO4XWIz8XQPoO8orBLg/AIRmGw0F3Nm2KpIOFQ7GS8cWmhF5j
jdYxB8CZdzp6JQ/ehfQ8OSPWZuxC2uCjOI54yl42hSvHfSZdkQqqFooL+q5+zrgh
i4Wh+Onkrav2lyk7gWdvJu0tC9Yc/bFEQS711V8Ohte9w5IVz6i55113VksmMTe6
ialQ2rlpYn3q8sJMEooPhUA9sZY9k96SN8aVy3C9ijwOt/6QjcjOXmfv80xHHxo7
Cv50Jf92HkTB2XNeAT6+nkS/jOZekVI+orgNia+nvvaJLh4Ny8lrAxMw8cDSiVVr
ifcTlBKKWi8RORYXsvFoyvkSN8RHzM5gZUhOBJex2jsn1wUlh6cv+AnyDN70rOZE
dwwhMOrFwwesjZua81qZV4Avkcn+aOyKE3DFZxB/Q4gfP2ij4ww4n0EhIJbDRwcG
MUFJxV9ekmju4BaiRNk2JToKv80Q8tTAmbY69U85FGEk9bKt6ZqFCK2CwPwvWrJK
b5Te/UWwUzBxQmVvKMnYPXJjad3O2ptCmw4gcrte4tRFnyYLOsEmtSFuqDGlCeDm
a3UsRLDp7KH0Y96tUtCG8pgT2/HSivP0RcYLV3RL6F0oRAgnQJnLbiGAgZJcaRHn
A0HI2gwvBDCbAD8W3PJFObj4npAG50Y6Oyr+4vFZ0UxXxzKhsGeu2MW1QmYNCh56
SOKCSZsLr+nvDtlpC/AGNOl38em2Ihr68tRdFrjJL/nD92DWXt7vIpSq31XKriah
aGfkyTCMbfjoGb130/G+6nSPhm6V4hhRX8qKLU0hHRVPVMyz1sJCJwwjj0D+ZhvG
cEBQvuf04asXW8VRUOWeFV5zE/09zM+XY1gRxBFGsOd2xhzICTqThlQuZC40ZGy9
Kg3V1gKldCDN17sPp+0xtQOl8QexLWCiiookhxlVz47PF9EuENpQq4id/ZjR/Vor
ovOHSDYnyI6ILRUdlfY4fIl7EKaoo1kovr/1f/NltkCYYiHxvTArzQBnBh0z3CpE
FFNfBN9yVL5B749QoMXT0AAaZYXXLkWB9TKYMVki/n3HuMAlfuhMC2qaFhVxi3zN
wvXCr0m5Riyu26keeEygadTj5P7NjuBS9WnG0b++4Mfulr4gt0ajHCOdnoEIu9iv
/7mvIgqBet0XN61D4DHENSJ0NGIhgkYq4CbXLl9Uekjeng+1HUEkdvGGxsRARnS4
cWkBzxs+iJVFAJm5S2w9+zwYxO5aM7meFfaZGHxGjO55DirK6+bLRJLJG0gOKuGf
sc0JxM8dQQlkJVJm+eLY4LUvh9L3usq2r6Jhoea91yibkZBEjH0IGmocfbHHr2nM
kn10bJFX6LHqCJ+LrAwxJ1ISsxyizKdbF7ZDBkzn97U7hVOpbOl22QdKjYp6FY1q
O2CebwAlmkIh0sjDVb5D02U10BAXl0e9W/cugCOkaPgr7ll/dMDCFR577y3GbM0/
sde4hzrbv3fvYf8GN544Po7FF1MJZbhDaCfGaaRrz14NTauoDI8D5nPynJpnceGr
uUMBwG+PQ97sGWPaLCtntH6VctrWl5odaD8tRx3FVaGwKvtfALNHAjo7jCKU64o7
ERM2hODBizJYrWhSsulyPoFRqovYY85Ch/56JyQE64RLBeCvnfhfdWRPyK/CH/j9
6v8AfDAnCFavyOM0X/j7Fk9WjeqbP1/X8F3DeG85NLAUi35INDM/sPTuEqBYpP23
aPOzeNG/4N9yt5Zv3LVzs4MoqhOLr3H2w/OJNxJycQ68OW1Hu9ZSkBFQV/lYKiIx
vSsHUEnT+dBF5TS18b1BKo2Vn0hVqnOdzjtLX9nhFyWTcMrlL5EdAzaxIeru+B7e
wMBwIwOdtv937DncOpIjwJrwNpA5cOPWUk2q+2c8f93dFTzfhBmzxM0+xl4PYht3
SOKgI8nRblj/y/Gia4ILZzajK2nKPpATVSCRIvaieeTqkRI0L5cL/C561XfWpZuW
/6l6tULe6D28w/gGoqsEkY/Jk1PKfO61xUiTTHBV3/2vJnJvR+9gvG9bUGK1R/HA
k9VBnWGCar+6aeJovOUoJ8MuOUQIst2bw8wGEU2Q1v0XhdaV7Ee6wmt1uUIPcuHm
PA4Y/oyk//Y67+b2JkwJsK87OCoZzeWfZ5b1//r7z6i1D5l9Q8QsIdUvNrnxN553
fH6cozh00EkvNTWZtSYmqTw4yYxOGls89K4EOIcgdG+AAjAvIZXtgNZ+/7GdAEkW
n3IVzx14Cna+ikvYEpTMagwHFMKMa3IsNldFI0+DBu12JFN8RZWS/9YdgQGtULPk
ksyI7SuIBTuL0Qfu3h33NokU/bOUzwSLGQXzPNBlYsLqYNRmE38m68CeckeRO7xO
sfF770NDJGTw/yyRIPkGreZYtGHVbUsaAKSnDbYoklrB4w41N+pPKTpUktRyHqnH
RzOLIMXU/I9tmMlK5WBMUGk07zFeK+2h8mD2yMJPFpENa1pei3Oy+AVBc3Yo1JVZ
pltPkJf8eESnD5vS2pYWHNZHk/fVS//l5XzDSqDq31jaxUC0TWSvnOnmYGCTHICE
SMoYd4F0DUO3hBB9/RT53R4lALPi1mRB6GL57FJR2AS5+TBRT9apknjEyO/bg5oq
qklYyxqMLdM99MsxTqBuvzE98VmjihQ2tskzu7b2vkgqwZZqYU9QNy6y5QCsepw7
13ks5XoV+NpdRTL5w07W3WVWzUUILMiqNaG55x72qOytN7nDh5SVOXQTeMNFb7jy
yxKYRtKu7MIlaytLxqytSMErNcjNsfQ7Y3c6pEUfWrixNtMXaCeD3+3WHX93Q6G/
WRFp+EpGSQg0VltONn8iXpN0VJxvDP5uSV2bPefLC2UmBi7dN7Vx8ht+o1lGPmFO
Z0+rofdmx0kyFh8tU1PhWBseQ2SKzBUNFhoX5Oac8Ltzwp/arXNg27jcQ2zZxkQG
1IP6xjm/WXtsW6YKVIQAQXPphEY4P39RDy4hHBmQfQ9WhZCCrztPwoYKN6IHzGCo
GQeKq78b3deM+/dZT0RXmpaSKwAi0OSdUnOGrfNrtK39ONq83cRBioavvfMXGCHl
F/O3CMycyeCt2kC02RIIAOJQeTZkE6biQ2BSderxi9p0cEfXC9/L1Wwm4vUFAUxg
almknj4O4oQEmZXKL/hCnTMGiLBTd9NdTHPF3Apnac7G1QweUU/YSRn0fEPLsKDq
2W4VtKYDJVWi8zze+xSmMfLQ9oThAyW7O9jTMXLZ8ysGQSdJO5Ga7TckIv7m/5fQ
UQW8kyMarpYesJs460hBCBy0y0F950eOmarrkA0LXsdQXNG59fXaQkDh3khqgGdE
pJ/6l/rtYNevBzw+au1lf1b5LiwPNEmQw+cA/7YKj2TNwH90ARqvoVOH80XjcIdn
4/SJf/qs6vOXc7DdaCpm3rEbN9HLF7b1gSPQKKIj+3bler5gpW3WaGatv8bBR5d0
KS+UxNrOwO1Jy9mXM/iFdIunT9RpComFuEsjdsrAs+a/P8z7lF8yVtcjxsY9uOeP
B1S0PaMCJ8eyxkej58acsLlOjcwIbbSr1O1XUsxlEprfcpOq2ksKlX/tFDTf+jhX
7qdD1nouicV5lttkzTFLiSsHOCnPDOJfQ9x1f8lGeQiEXxdVdp0if8Is1DemZ7PS
0pXWaCeLzwt7FnRgodw5ymMPO/nxewORxFXy11nYT7/49+3d66POTBDDu/r7lKID
gmpAEM2tva/R+fWv1hlNY4UQnimfRPYFnEaWVGVPU6yCLkF6VstLSuotBKrDu+Ps
jRH/odDwzRgcrxyv/Gxo/Q1dfMxwWp7wtFx6+dlD3pm+/rokd7hcVCTINH/mwgGO
c+jX/8Ec7aa/kmse+ENhenAQD0WttX9tRqImhLvHG5s=
//pragma protect end_data_block
//pragma protect digest_block
0mMMaj8RtdMQml2MY07zFb39ViQ=
//pragma protect end_digest_block
//pragma protect end_protected

`endif

