
`ifndef GUARD_SVT_AHB_MASTER_AGENT_SV
`define GUARD_SVT_AHB_MASTER_AGENT_SV

// =============================================================================
/** The svt_ahb_master_agent encapsulates the sequencer, driver and master
 * monitor. The svt_ahb_master_agent can be configured to operate in active
 * mode and passive mode. The user can provide AHB sequences to the sequencer.
 * The svt_ahb_master_agent is configured using the
 * #svt_ahb_master_configuration object.  The master configuration should be
 * provided to the agent in the build phase of the test.  Within the agent, the
 * driver gets sequence items from the sequencer. The driver then drives the
 * AHB transactions on the AHB bus. The driver and monitor components within
 * the agent call callback methods at various phases of execution of the AHB
 * transaction. After the AHB transaction on the bus is complete, the completed
 * sequence item is provided to the analysis port of the monitor in both active
 * and passive mode, which can be used by the testbench.
 */

class svt_ahb_master_agent extends svt_agent;

  // ***************************************************************************
  // Type Definitions
  // ***************************************************************************
  typedef virtual svt_ahb_master_if svt_ahb_master_vif;

  // ****************************************************************************
  // Public Data Properties
  // ****************************************************************************
  /** AHB Master virtual interface */
  svt_ahb_master_vif vif;

  /** AHB svt_ahb_master Driver */
  svt_ahb_master driver;

  /** AHB System Monitor */
  svt_ahb_master_monitor monitor; 

  /** AHB svt_ahb_master Sequencer */
  svt_ahb_master_transaction_sequencer sequencer;

`ifdef SVT_UVM_TECHNOLOGY
  /** TLM Generic Payload Sequencer */
  svt_ahb_tlm_generic_payload_sequencer tlm_generic_payload_sequencer;

  /** AMBA-PV blocking AXI transaction socket interface */
  uvm_tlm_b_target_socket#(svt_ahb_master_agent, uvm_tlm_generic_payload) b_fwd;


  /** Handle for uvm_reg_block, which will created and passed by the user from the env or test during the build_phase, when the uvm_reg_enable is set to 1.
 */
  uvm_reg_block    ahb_regmodel;

 /** Handle for svt_ahb_reg_adapter, which will get created if the uvm_reg_enable is set to 1 during the build_phase */
  svt_ahb_reg_adapter reg2ahb_adapter ;
`endif
 
  /** AHB External Master Index */
  int ahb_external_port_id = -1;

  /** AHB External Master Agent Configuration */ 
  svt_ahb_master_configuration ahb_external_port_cfg;

  /** AHB svt_ahb_master coverage callback handle*/

  /** Callback which implements transaction reporting and tracing */
  svt_ahb_master_monitor_transaction_report_callback xact_report_cb;

  /** Reference to the system wide sequence item report. */
  svt_sequence_item_report sys_seq_item_report;

/** @cond PRIVATE */
  /** AHB master transaction coverage callback handle*/
  svt_ahb_master_monitor_def_cov_callback svt_ahb_master_trans_cov_cb;
  
  /** AHB master Signal coverage callbacks */
  svt_ahb_master_monitor_def_toggle_cov_callback#(virtual svt_ahb_master_if.svt_ahb_monitor_modport) svt_ahb_master_toggle_cov_cb;
  svt_ahb_master_monitor_def_state_cov_callback#(virtual svt_ahb_master_if.svt_ahb_monitor_modport)  svt_ahb_master_state_cov_cb;

  /** Callback which implements xml generation for Protocol Analyzer */
  svt_ahb_master_monitor_pa_writer_callback master_xml_writer_cb;
  
  /** Writer used in callbacks to generate XML/FSDB output for pa */
  protected svt_xml_writer xml_writer = null;

  /** System Memory Manager backdoor */
  protected svt_ahb_mem_system_backdoor mem_system_backdoor;

  // TO DO

  // ****************************************************************************
  // Protected Data Properties
  // ****************************************************************************
  /** Configuration object copy to be used in set/get operations. */
   protected svt_ahb_master_configuration cfg_snapshot;
  
  /** AHB Master Monitor Callback Instance for System Checker */
  svt_ahb_master_monitor_system_checker_callback system_checker_cb;
  
  // ****************************************************************************
  // Local Data Properties
  // ****************************************************************************
  /** Configuration object for this transactor. */
  local svt_ahb_master_configuration cfg; 

  /** Address mapper for this master component */
  local svt_ahb_mem_address_mapper mem_addr_mapper;
/** @endcond */

  // ****************************************************************************
  // Field Macros
  // ****************************************************************************
  `svt_xvm_component_utils_begin(svt_ahb_master_agent)
    `svt_xvm_field_object(cfg, `SVT_XVM_ALL_ON|`SVT_XVM_REFERENCE);
  `svt_xvm_component_utils_end

  // ****************************************************************************
  // Public Methods
  // ****************************************************************************
  /**
   * CONSTRUCTOR: Create a new agent instance
   * 
   * @param name The name of this instance.  Used to construct the hierarchy.
   * 
   * @param parent The component that contains this intance.  Used to construct
   * the hierarchy.
   */
  extern function new (string name, `SVT_XVM(component) parent);

  // ---------------------------------------------------------------------------
  /**
   * Build Phase
   * Constructs the #driver and #sequencer components if configured as an
   * active component.
   * Costructs the #monitor component if configured as active or passive component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void build_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void build();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Connect Phase
   * Connects the #driver and #sequencer TLM ports if configured as a UVM_ACTIVE
   * component.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void connect_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void connect();
`endif

  // ---------------------------------------------------------------------------
  /**
   * Run phase used here to set is_active parameter (ACTIVE or PASSIVE) for master_if
   * Start the TLM GP layering sequence if TLM GP sequencer is used.
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern virtual task run_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern virtual task run();
`endif  

`ifdef SVT_UVM_TECHNOLOGY
  /** @cond PRIVATE */

  // ---------------------------------------------------------------------------
  /**
   * Forward TLM 2 implementation
   */
  extern virtual task b_transport(uvm_tlm_generic_payload gp,
                                  uvm_tlm_time            delay);

  /** @endcond */
`endif

  // ---------------------------------------------------------------------------
  /**
   * Extract Phase
   * Close out the XML file if it is enabled
   */
`ifdef SVT_UVM_TECHNOLOGY
  extern function void extract_phase(uvm_phase phase);
`elsif SVT_OVM_TECHNOLOGY
  extern function void extract();
`endif

  // ---------------------------------------------------------------------------
  /** INHERITED METHODS Implemented in this class. */
  // ---------------------------------------------------------------------------
  /**
   * Updates the agent configuration with data from the supplied object.
   * This method always results in a call to reconfigure() for contained components.
   */
  extern virtual function void reconfigure(svt_configuration cfg);

  /** @cond PRIVATE */
  extern virtual protected function void change_static_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void change_dynamic_cfg(svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_static_cfg(ref svt_configuration cfg);
  // ---------------------------------------------------------------------------
  extern virtual protected function void  get_dynamic_cfg(ref svt_configuration cfg);

  /** 
    * Retruns the report on performance metrics as a string
    * @return A string with the performance report
    */
  extern function string get_performance_report();

  /** @endcond */

/** @cond PRIVATE */
  /**
   * Obtain the address mapper for this slave
   */
  extern function svt_ahb_mem_address_mapper get_mem_address_mapper();
/** @endcond */

  extern function svt_ahb_mem_system_backdoor get_mem_system_backdoor();
  /**
   * Set the external port id and port configuration
   */
  extern function set_external_agents_props(input int port_idx= -1, input svt_ahb_master_configuration port_cfg);

  /** 
   * Gets the name of this agent
   */
  extern function string get_requester_name();
  
  //----------------------------------------------------------------------------
  /**
   * Function to get the configuration that should be stored for this component
   * when debug_opts have been enabled.
   *
   * @param cfg The configuration that has been supplied to reconfigure.
   * @return The configuration that is to be stored.
   */
  extern virtual function svt_configuration get_debug_opts_cfg(svt_configuration cfg);
endclass

`protected
eILDB>]2IR<=7=],.JcF5e\X(=^/8bG/E-81(P9=C4_4PE>=Y_HF4)83^UY-Q4Va
@0^)KKP-D^:2ZSd)1#(N571Q1dVNDPRS.e+YXI6-TU(_;a]_aRJ&>(^7BIB/6a+g
])8GU<T/F5\MCcF0N7=[Q0A;J./-YgZYB(WKFgaR+#O<F.>>]b0SZbD\0b7K.4L5
N34@d]@G8bZ<?.AQZ18:T>93HQ+Lb^K,:fCc88D;d/0_R]b4<WC03<7#-1.\7g#c
GEB]89+H\JL=I/ce1@QfCTC9^^2VHC+@[<H&IO(<\);_C$
`endprotected


// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
  `protected
#a0gE]3/4,]FB8PVGL[b>B\:=F15f[XD\eF6.+QdCd9[B02>0PTa+(dLC&H@Odb4
+&f5P<(N4<Bf@Qb4N2Z_SF9<WMg5d1KdeBX=H)IW0+S5ZMANC[g&[O]9J./()30J
+Bbg1YgLYDYT=&d&MFfLJ1ef6/-E,&4&a<b0S43fYXSB,1#23.KKBUfd+:gdgO4+
Z4UFSH+(X<?PB9]I9I;9U.K<[_L?EZ;@48B)=gK/AXYNLd[8JCTaZ=MDX_Ff.J<4
FRM98_?/ab30c=K:#XaM=4LJ;?O)8fR1>7f-,F\#V#F(N4[:C989V5RAO4+-0FWA
TXG9.)R2T0fP&FG\<GLaMA9P?.<dYQMAK]0ROA(deKUa3,M#E=AUTW<IEX<^7(-P
8Kde[]_fTZFC\U,P+N]F>AZd@KHaX#GV[FJI4aTfRZ4<7W7&+gf@d>Ib\a&GI4eL
bN<LQ/T,QAcC(FagMQ+aB;TWc2E7P7ZTKI-QPJU8&F)D(9cSI/4W&Ae>&VB>Y=_>
A?FMWgTKUMIF7Md&De9M\-N9]QPU<S;U>:MF:)IXY7X4MQU@=bF2,4AXF-(90QFW
e7A-HQH><>SN;[.JG+^(0,2/U;PPTJ^R5gS/[7;gLdLC=0LZ^Ib\HL=@#2&)AG9b
VFS?c#Kf6[9O;BY?FK&?>D&7FI/654Z1Gc/V_Ne&:4d5B;6L45#HW5SVHWLB2<Q,
.LVcOY2FSeI&,+\BdYd+NY,?3K&(TFG>P+X[7PJ_1Q9Z1[Qa\J(Z/ZNYJK_eHDFJ
=;YON:ZMK^,J=Kd9Z9eG,&_.d:UZ?3/UWf8RcVST,b?g^1AE2b+G>ZFVHfC5CPD)
PI7H7O>G54,/A,Ubc8@_Y3UWIa&d6Q;],>ccRC71f]_c1_=Hf@Z==?J2W>I[[#Ua
/T)#]c[>K6Gd;E2bXKY/5)P#\3EB+aX,>G6F]S:#eEc+61>)aX&9R8]U\STQF>K3
1=/Lg+g^N<I@ZF@Ec?VKB1+Z^7Pa<#Z+a:)Lb[g[N_:-Gf4_P?J,9_4DZK?QDX)7
FCIQO?Vb&@5+@OO--5I3M=->1A.,K)WH+Uf3VMM<QdE]/b?YRe99QcQMAR<c:N?F
0H;Ba]>XdbD6He=Y#5&^OLC,Fb+A-b66D0B6KPK=a4KC@1(0AYL2+B3DXA\b92g@
T2?S?TGDA\[@//I(OMRUE1GQ#G#1b2M^HN:e0U^Y4+)V_?8XSEAJaQI_PLQ08FZc
@O#)4e,-?cS&>VZOU#a4fA@VN_>7]e-.Cf?&T47KS9#1J9WQ@cbNN=5a&35WGU=O
+5K>1ABWeM#=^5YD#Q7G]G@++--Y4b\XC(a/8^5#D#8Me_J<S:5C,<7C^(]0,E=G
I1]G^O8<+B>JT-[)S(<_3+[[gH_1@L40a=]_=4@U2@M4]#WT_D:HUPHg)KSRL97L
d40JW=)BJG?Ig47dLQCVF1956H]@Bd>MB[VT]TgKCPJ.UB4)Me1F7c@3Lg,^_)SF
c#];Y33,N#c)#N@\;=D;/(fI8,gVH.N.[AB))K;6Nd:W80cAVe.7.Tc8#7AW)MQJ
,dXO_JBdH,f9+]f]J8Q:F=;CI+9KC5CC>(;@\6@WXDd1NT\JV4_OYg4Q/SC=LPPN
Cg(bcCW=5,cA7Tfd(Dd)cDfTaMJQEYBfL6[YL&6\a&:-9FBT+5#?BP+A(T8R\UAB
?10BU-NWX>5c0@9-2_:aJ1_gHM3?=O>5UMJ<4aY5PD5R)?-=d^2A^+RE4+_J18W)
D+M_)BH7aEDQ?INVX?>0T[]V[:C21eC6>?^.U=G@YP_H,fK2@9L?<ORH&Y@,K<b#
>b#.B>\Ade0Z^1>DD.P.KY59ZZ:WO15_3O5FAfWZC-M@3R0,Q\OF_eBJ1_2Ib9/F
#JZ>40VPXP.HE0/>0]X-HW(1e\eI4@NWWEE)Zf:FK5a_&U1VfKIbU#F]@93=,PN\
@?T@UJ[#9//.D@C-ccOZ9YfB]6AS/^Z24]&3Y\-HR7;<b2)fR:::eLY&W:DCF/Y;
USETcg]SZ>_C=U,/K_QUR@eE#4&6DQOU[-gN2T[c31fU;+8E<O[2A0AG^YP>GR49
5\b+d8Z+T^B==^7BT(UZFHER:1f7a5=TB3O,#cS1>9HE[Re#WcN]&5f:b=4B6B)J
]C=5U6eN.=&]7a?Q5U],O6YSS+LH2++NcE:Q)<;A5bLSI\dR@:^ZEIGWJ5,N[2EX
/:Qe>\c<5d[g@C7dMA01PZ@:b8RK0-BPG#?:?4.d\SQ]-;\8g9BF;/PL=(bfHVcV
b1^0faOLJ9F&6R[DgT]e)aUBc(5?W\Z&S&Je-83;?Ag&RL>eZ\cbbM>OQ7:XX1I]
E0D8WX+MDgD]4,VI/Xb=R3GN;.RF8>]D?S_gUN]bBRSZRI1/EV(Z+c6ME?]_E&3L
ga-:2O?</5JF5G/I_:2.F>GTdFU^bGaGeRE1gc71bKFd<27c+)gQ<ARR&:W2WHf2
<DF+A92P6-V;J^#&DR5Y@4KEC+\A&QA/_:Ff@C9^J+NePE&A<#6&6Y-HZ4/7KWU6
a=R#IG^fN+KA:g_D37ZD?U42:RgHM/S4P=,82F215#1[99_0B/P9FA^AU+b(EO-,
agA@R;NXc1HTC7(2LTPAA^@DPZI1G5/e9Ug0^CE3Kd]B7&VP7VeDP?;eMP?HRE,^
C-F&?Ca=Q#,B28&fAPUCc:;S;9KE+OH,&6]BBd5E>C5OAZ;dZI7JKfJd-a[WSE,/
F\TCR)1fcM+#:Z:N8e4#T\;P3UAfHdgV4<[/L9KTMZF)392:;<aVGa1V[U]\PXFb
IdFd-BKWGN3MPdfPZEUH1CefcRC0fZg6D1]GbMF\caAOK/U(<=HWZ&<ZXdF^CB<W
S+6(]EX&0W?<ZDRV9SA1CL(1L,&:.E#T;#DLZL_Pd2QSfWP<bg;5SEUN>fg61A<S
(Z709Z(F^,4+7=^8)2TT91Z_=BX&?//26,^EW6dUW=UGESE-:=EdR_4W+ZY_f/I,
P@)R4/H_F9KEF62M.\fS0RWbFMP/>.6TZDAg5_Q^Z=EBDEY=?F^b,Q&3@&O2Vf)0
D8V6-EIc@4;<=IC80ER)5CAKUb/d8NN39]<;-a_Z]V7P=;W+J:aE>,/FRb=XWWQR
703]B#Re\T_FT&3&ZJXJZ,W+IHW,^e9S<GPa_9c(QJQ6D8O#2aI;]V6>.1;F/-bI
+22C(+NJGbKd<EEW&Ef6//P=5:R>P(,2VF\KYQT^0SC(\)[#T[YVDEVYE:dBDT2,
R/]99Q+f)059D=JL7@>V]=.-[46<F>^gFZZ0Na6bGW:;EI\Tg1Tg0G#[BHYCJVFd
K[UNE8^Zdd]b,S.aB6.UKQ>KR=_YAbHK_2B009^d7N+VP&Z/P_TM1N.\7VCK;>If
0-9OG(X[<:(MK7:W[.?NeZ.2SGBUDJD2-B]L>HCE4YEJa-VRT9\I<daW25a/&J?T
0^>JN>/G9.7S3<R-JAaM7326G^^+5U&,0KU\-^E5EFSE2&04&>e8EM]5I_B:1f1)
BUJOJ>(59)Z#;LMT1O_XfLC(C3>Y[1+H?].L=O_+gd3HdaM/\aG4\L7P[ZN\;Z+b
#GVMeL[A]gGKTf/>E5X^,69T\1PgH86f\<)NGEdXdFX@),&.U;F)4Oge44#>;8RK
A3ZBaF2OB-eA(]HP#&(/)AI1f[X2TZ4+=eP[<_/8Y/^bOb9.<[K&#1+I]@Y?VSa0
HF2a@YMKd1YC?5.1-NQVb2E7,^TCA),e?=(<OI+-dg[U_J.I.K&>N#WE#+<H14fb
cFL@(@#.fSIDG(/&gQ(WGYK^1H<[L[LZE\:37IGT4.)53+-\:C+4SO#PdVa_EG6b
2G6e(V?6SMMS.FJ4SQ/75Y&<62X2@X>[O&3Ga7L5IV4LI3Fc^AXeN?OA3g9bU_Sf
,^58?8TXga\6]/=d)A<?1TI[F-AgN)UHG6c_G2GL8OQMLTX/8+0UfII7D&9J[PgJ
&YYb=>(<_EG44S[GKS3PPE_RY3c^LNVe3b>N3eB.g<b.QL+ZOC&.0-2;BN,f.+3^
gYHeXU.>2(bb9)352+g@4\PXH41#6HUN0DMJC)QGC(=1R<+&I<6F_E2\eSL9f&F#
:0b?/bQK:@4\ZKP()A7DCR7VaCJ7MU/ABZf9ISFDSbfR6N<a<bUAc,Jd:8_fP.;7
L8UHE\AW4/P0HPEb<<^<<cX;H(PECC0AO37LM:@HfBGY=8+3S[L=[HY3U6fE5Lf\
Ia)eW8Bg+),4U>4fK6S23-KKF>3HQHXLJ_:2+P@@.([22SO)K9-G8T#/P@M/T>>S
Y\T^AA,_)g/=JA24gE01Y#?=@fABTI4WF0>H\C+9BG7#^J[(RTAIc(B8CB9G3LKQ
3V;A;J#69L@7MX-Q/B8A5A+RUV@7ccK-_#+6M</S;W,#d&?K&:Y9E>+9<1aGcX8&
]8cY(L5Q.-[I+_ccX-B:5TR128:PPZ;O#P8H[XH9aZB^.?.7HAOZbK2VB/Q0_gDL
C&KI,<ME=;:I-JRddb_J(#eDJ?f&#Gf#624IYDH^Fa_\#-eQCF8DA?EAY#R2b\K5
:.XE=USS6]=Y\=_eVVE[?)e&P\U=DF&,KWZ&D?.&H>0=(S.VH/N?cb)bAEV]MU91
3a(_@e2;7T&A8R5ITTS9SIRA85&F.4=,@CMC<fV#;]B>HVUG<:MdZJB7_#f_e?QN
\S[<(f\I2EV>B05Q#7NNI]6\1?M)0+_Z9Md,RYaN3DST-OeAH+/cK7f#Ba[G3.R>
AMeE&#,/V_CC?DAe==geCdA3FTNgFB;7-U7H4KYR.J0XVYD)L;8b+cE83F-+Z<3Z
)8>9>>((P\^=O?:(_aBDTd\WN@gUKa=4V9U2V<I3PEW\T;2<<669G,eO&\\PV,;#
Z\I)J5LcDXP@F_XDY(-?RYbJG[=KbVHI8E)P?A;&B6e1b=QbGT=B4a9fNF>4b4M3
Z[_2#EC70LXL.Wa9XbLMDYaE@E1)#_f,S@_<_1Pc(&PRR,LH.ART6e?e8A0313HU
ML#AR<Qd+X#R=KDa\K[,H2I<R+d^S;ATG_,2]M_a/GMV,2_HYH?G(7/T^R>=1ZPF
<8DD20_VDe1<JdfR15Z2UA/f2Pc4/P1<bXOS,4QfJKWJgC=bfE)E^RN]DA.A@_[,
C@2g/Q2gU9HFB^RE:\\;[4PBLAI.(@;b3VF;D1AJ.0\A&Q.)f:,>@eN^WR--O+fH
c)YaC5#+5U7=-^8D[(6@]=YTC2S#2FO;)WGa.ZJ[Qca:5RTH6&26_@]7VPfTd.E_
5]5f&]A3BV[0?/:9?/CE.Y9_TGB,V:+?YP1F8UQRdKR=E\-M0Q3TLMC(H3/[A-6-
P0ON3>.O\)1e_D:0_PK]JNH9XB3VNPfP=/MJ1GX^1+&1Y#2QE9F<f^<\CUa2DS]0
_PS;^5)[WJ@O([cT0gO9H&f5]_BS1L5EfC^[9Gb901LU-JBO,gPPGW<(L;^e#5WD
/0FFHE8FW<.ZK/Y6gf@7<L-)a1f9,RXXDXPF43:>#ATRHaCFGBbFKcgKHKN7D+#Y
&;g=32T?CgC7=9T[:Td(Q[2@.NX-DO]M72Gd6eY6XRZEZfR/Vb7PAX8bU]Z5PeWJ
M58,a:f?6d[53,Nfd>/E/R7[,MF?e3]bd-E:\M(VXV@FG(b:B_H(ON+&+eaP.CNX
dK_-@3L;(87X.3Z=RL(9Af/;E;fAM8F7@fLJVMaK2CG=0P6N3#TAIS@\0@Y\-+/a
,9gRNKe5gC\;,-BeN2RgH-8CF>3B6O:M@Mb]MUW2f[TFUU#EBCRf^]I@1f1/d._e
MN5-1<E=/NPL:(VD3eIOXD^EQLTY--+1-IW&YWG>,+(:=.d8S300gYf+8c1@X_XO
,\bIYaES/XUDBgd)^aeRII[b8CIQ,C+@1dV=f5NB[Pa3N+CJ@CR@L_1UaX]#<C[M
22F\B(O5:N84JEEVV[HfZ6;5]S6fH_H,8XBC)91LQea:XCV(a8[SKCa4W3OP1YV;
4.fGTcW5,3<3XCfF=#NEbD2YMWOf?d4S2Df&H@2.;;[S<LB3&W>gG+D>KSaII;[G
58B-b3-/B5[87/NK>&ZV\??C/-R8Hc88&H&RCfcJL8W?,TS0&+).&3([Y)+7gaR9
-db2:CF.BW)=M\#@^E7JC[(M5M[eab0,aKE/HO>/D9-#HgCOOZNfQ\Z.QT1W[g4A
Q@+W/:-6B-DH9FdKe_UXH;[NU.NIR46N8WOBPU_4XC_GBaa6EeO#KGZ4^LbY9T@F
(_BNF=2&?3,P]>+/\)_/6O91Cd00]R9a(&g\5K55-NYNcLXJ=QI>X59;1./_G+)Z
PVZ+e_0-B8D>JN#^a6XLMDeOe2,OAC<eXI/05V9gf@,=K#SgRO[.Z6M0dX&f=Sd7
I:Y(LF[<TfaVc)G7K53fM0.a4D8a2HI:X\XNKH/E0JOMOP.X@ADSOf)?a&#B9[OV
7/B07aN@ED]R==_U#(E[fEfN^@2@73\[@gQcg,+D:UF&?cC+D20YH55XR2\J<1,9
a5UeXa;ERa:8b+:?S.P-[;6XacUW)OPX;7g)38:dEfBX(c,FA?fP3FN@IV,2b-Ib
<HP:A>.E>b]0>bU+H95OD;N1D2Y:MGJ>S<><M@a#Sd)>d-Y5(VL;S(TVJYU+\]=W
/M+/XN8P00N7<U-)F6529d,A0_&VgP=#TK[G][W0W5]N[;5<83bbGdU;045^@VMG
A&-H:cWTcK\M^<MXMD[Z8XNL#>9REOeG_gYU468G9SH.[^[HX3QZ49gb=6CY;#9C
KcHAb13Bc96B5ZY7&^X:)aW23d[,WJL0K,[8@):c_d>\KLZ4E..BU?0_2UAfBAaG
8Sf0TC;Yf?G\+[<[+,.L,O;.SALeY5)6DK^dO]R\+[VRA<^\?UW@C)>VD&1IH5B5
,);+50_(@7FTO9)aHQ6A?4b?GC[-Q+A(]JD9Ba2Pb\4=U;\^L]08Qg7dY/d\3aTB
@^f0.24FD29EITG>2Q&Q]/90,d(>LS<7MUL&2DI;Ba,^(2N0T>L^EJI#POU\26D/
S]aE+]T==V]aKa:IS<@O9;;5A84A&7fU8>VQA::,=52SX:S/#;f0[aYccBeMTREX
+47#X,=JWMNZ/XOU@UZ#?e-C+A[=&0G(&T-5N-Bf2:dC8,>=4__L_WR>?gc9-EJ=
g3#J_[\;:><GFT<4>K<Bb1[IBJV04(T;J?dPKW5e2cUO9YK-H0FOdb7NK2c.a/eZ
c]504ND<b\I->THW>L7BBWc4+8Qd:V2\Sc:&,K[?eHI+-cXF=A+#;DIgg]6?^=\7
UbQYTI(J6ATR/T6a<<b7CJ3LMbdePH4>:0;g&Z]5c6NYBGEBegJ3+Z+TX8Pd],B9
SN^F@KW:5[eHY)fEAb/NF\8&C(=E/S0^5I9U0(])2W)8b8#SY<2:TD3c8W3WQ@QR
@2O1FHgc<2=D3Y2TGbdIK@W([:\J,a6?ERM=SFHH1-1S9V4c:OSLF+K)?RQ=^F;T
T>J\R0Rg931Q),92O5;g#LC).-Q?X?\EWaE91Q1gH(3QUY+<&X(9W)<Z\[40(P:(
14>QF<O>)(V\IUY1&(=Gc\[6.Q&@9L3<dZHOfQ5ab@MUX1N?182_N[8@ZcW0RA&J
N8,H:5P>Z#cXBP:_46KXedK5DefRH;^aHHE#Q;T+^1^JDIOGQ)9eE_?cd>C5Y)[b
OKFM2+<eL.+=S\Y37F;K5_7A&P)?+6OWc5D,D=1C)V[fFfJZ-2:N^M<CBJC28gMQ
S9g5KV]9@]#7b1#_HaH;U7fd:#W]G[_6ge9YVMO]d[#KE>:0[_(<@YU(,d(J\.3U
>I4?#/:a:#NA(D6F]IZ0Fb#Nbga<?,@N71Fd,].J[DMBFB24BX#&7,/M7W:7CV5b
07ZE9ER7U.9fdJ8P[F:a95.7@F\:T(WEg81EJ\=N89+#35Q1>-\J0+Pffa??I3@K
N+NYNAaI][=NWWP^YW)DD&>9)(9C-+Za=H(Z>,;d[EZ::7#.[JU?W.MN]S47^/XS
#/=,AI@0EEcWR.B@-S:)H&7NfA-c..Pa[4a&X(DNLVC2,S@GA>2LIeA:(<5B#+&=
6T&],0A328TbN2OU:N>8E059J^(T.T:FRbT[,MH>@YQLaTfcfCc)^(6>S(WgZ)Pb
e.Q/)R>bNaN6Pd&ZQ2a#E_0b_U\:WM_5H0U7VY&:fe65CVF<OXfaX6L;Q42B6c#<
P[dKg2@5dRIL\ENM@\,:IB3M\MM0a>G^_)/O&<(]SJ8GI<[:1e6(7J:,bZ6)e4(4
dR2]DI@cF0.W#(_dFX#;[A:>H4JIP2=SS_(P]<a?RbeOD9T>;O8RA=F>U6>[=>_H
QCZEGbWYCHdX#[gM-BIYN0bW@0=?(+cKdf#]PWHW9S\1B]/M3)3ee#-&Q7A715V]
68Y&&E@JD[AF+EbeNVFc[I.?fXN;T1+<A?R.OCZ3a])V@O..A;1>I;4eQ=M[DSW=
/SgbSN#.S=gA.ae+a2c^=76/SVE@O]-P&#Ne,dXME.cU?IBV9g5B?bGP=2f&>Yf5
?V:-&TX&d:K5+TDAS1X_d+;BI36>g)::H:[LJWR3g)[bVW#\eO=e4&_YE^Ka=GfT
>^(^gK1aba>C_9Y7A+Z2dA@IefEFfP&_^]cYQ^O:AeRaNV.&6R9X&[)_[AQ5UF0Z
8_D=YgU&)YQ#]3&V3#>;eAU&P.4K=d\-XZIAB7((YY3J[ZRd.-g@#X;M#YKLDWJY
a>ac+AfU+T5eCJ3?1&[M6W:K\H:L^+IG?2>QF3+UR>4?P>D_a\(?[3?MJ36b?JR=
V_3bWT1XLSdIRC<=aV2]Y=6I(JY/ASK(H>6NbYN&MTLZ,5:9^;R+GCA8T>fMdXZQ
e0@;/Jb7B8]JK#^GZ:H=D=P_&^WKa(\N\a&;];H/@JdUFe<EGb\\TRZ]GCEa&?./
XcWF/Y78[]J/VJ#Pa5XK7+#>a>A)IZ4Y=^=APAO.Ob)fA]9.VR1T)/EQC7)PCX;L
;DPO0gOZC0<1EPa91<S:G8+W:@29-.?dBE]ObI2f0bGfL>IO4\ZN+D,>;?b?9&4>
TNPBUZXW?=QQWCc4<6.GX5[=:7)MF.e[]@5g)G()ac>\HDD6O2@BE(E]R129d/7(
@=(_c=(/.Z@BV<752K^TP@V[fQfZT,,/?=DMV+(<P@@7[BL0Z1NR;ReQ1@R2H9C[
AM_:[8Q@@#1D,#D^gK+ae6PW&A8>Z^CaO5ZV,E(96.9G_-HbZP710SFC\Sb47=ZX
SM=,7I5;0)bLcd3Be#\LeYWB7E)C80L<8bQH?ZT:),)AZXP/@b(J)C=YJ@aH8ER3
J5T(^-B&7c/01>,4\a)1(3\:g4\EKI65476GM+\eK1_SQN6I1eTaZ\g[)Y>aG@..
-P@ZA\Jf,=^1E>dOS[+Ce7J?S8]eBQb.S;EaIAVY0f,L+2T=Rc50(T8335C:(=cc
P29Z1,&(eMT0LLaJ=LDRdYe?GD[NZE)YG:fV([2_.-[G;MJ/NabS6X;G.\8<41S>
SWA-@Y.4@G]HYV#VJEIE&]&b)b;]CMgL-XM1KDG<HE,:0;V.LZJ>\=]JM[0=]]XX
(-6:(ZDJ#JE7)c(W#H(4dfOK?[8M]<>E.E62;gaYgG#QLYP5NWIF2EGY1>FeJ6O1
APAM^1bU;=]^/#>7R=OH?7agQda4O=:1]PeP,(O6?KB<(TB@[;d(aA<IN?Y?\Z/2
E\][@dFeH(Rg70f8P.TC]^;CZBLVEV<Ob]]YP7_ET-A?+T)0bd5&TZV,W;L\YGag
26EeSN)]#:7cR&@bZ,/SH6WUBVS#=5[/&Fb>&BN\Cf?82\?>6D#G/,Q]&TcPJ5+U
fR.)bU/B-M3Z(RNf3#[<_A;c..L66CE<J,EIACe9R=OZ?G7YJBF)\+DSZ:3bTK5b
TI<4Vg(ZEO=V3gOYJe1F;?:S+J=c=]0TfUXJZY:)/EE^+GQ8Ff#7[K^W;.N;]2g>
W9VU8HN3,#F-(Y0ZX=Q(N1.E1MHeH&/YEXZI[#^8AK#]0/XU_<R,e:#L^NI9_a81
QM,ZJ78+VQd>7G,aDd\,/Q0;A+<XTA_Q#?g<A3[^/\250D8G<A2M/-646C;4Zagd
7[da+\&)g[#4Hef>TdZWL2Ud@cZI3_BTSP(.<:R@Y5YdN;14]DD#;Ub2/fUP3NT9
XfUPgZ&HC#7aBYFDNHZDCaV]>,)+,IFb+_1\S;5+L,K]@S1D+0(C/&(.=[eK-Xd[
.PNBB[g5;G.LV+&,;aJ?JbO/M</Ifc:F6/T#KJ?)M,K4Z<_1b(Q4=+0]]d<;<c.H
H&_TI>^HE<>9T++a((N]5-M-<9W;9I.G-HE?;adE8[6L+RGL1\aN6#95/\28e4XS
dDA][(fD]KLGYU;T.@eKDcHAF&,UCBH?dFa7d-D@6?+07D#;gW[7M@3<0R<.E2d&
Te3_Mf0_OCf?-4DRBHFfXRD0gbWg?OXN8c?AX-b,M-?&6A,7PA3L8a#d]Q0Z?De4
CcJU-,9:EMXMDI68e5>F96L(V:FCZ60WbX,ZR7HWc\8:g,Q5J5McWLe+=ETcA+;L
02SB6e^A?S(a)B^I]E2^F@FaVC0,43VW?R90/9Rf7OX9O6,\+I7TYgcS<eY]A)3/
9GfVF#4@&G@[FgGW13fc&d+Cb3FSR>(dJZ9R#8#Jg,=;TV9O1^)eMVXE;C>\-a[-
IJGI\CXWc#C>3D7+A28Hf+0gB]g;>#YLHIJf=IJbGZeSeIcPK:13R/O,Tf>>S<Z5
C0:/YI7A,,U;O05\C3_I+N)=547AD0cXa]9LQ[C3&d);33+;Q0e(U.BI;L3T]I=Q
.gKJYKL6\X6Tb6OeO\57#REDB-8/\FG4SY?0\BU400HDUJT[;47BbB]FTL;WUF8U
D/#W[U@4=Ad59^>)a3ca/+9IKNE,Qe3@XY#42H&<6L^>5)A9:1b^+\:FAd&B>Ea?
X)4V8JWIY]\+6-KYM0)Q1d8g#8Md6HU\dFM&7#UD8)aP?G\=9@B_b\/O3_RT#8M>
;?F6S43>bHCPGdNFK,JG@b#@fQ,0V-I-Q:[Yf:e_K_[=d<d^A,+c#SL;4HO7KM)F
Ng?#KQ74F5g(K0>a8H+BM6c87SUeWW(_LD#:=0KAg9IgR(DU9QH0G,T1BH43L_:T
L)3+QII.eQPOR4Vc\FG-44G]dQ]RM/<W,UJWH^9TM9=C1U&E8?c.3W=2TeS=g&2G
g[AeUSa;cP2S_C[R>#3=DGQd4GY8b;=85>6.JW@_GK2,DK1g4EE&CIGY_b-;6Fga
+PcC#Y3\)De0N67OP4YJb/9cRe,T/:-N6c;_[(PeF5,S.-/=(7VFY8NEJ)@F)Gb,
C(6DU&cQ]_&F<;S-cFS>5gLD&aP6ES0>5:2^#1AFL;2D&&([c:OOI&J=A[)^88g1
T]>.KZ?]N&A&.8HK7K<BXdLaN</@N79(CLK+6-Bd[48[)_23>-Q.KC>/;6fJ[Qb5
#7>Ng5>>0(Z)V@Y_^69Qa_\8-1[bdD1Qa\:I^OeU+BU^K>L):J2f?\VIb7NaFV@/
BD7C(/,0)>fLANBEJWJ]Od;(DY3UNaR@9N/<[;..Jf6gDX4e3dL4(eP1&LA4c/WX
+G9CJf3@H:^&@5:2;@;RI)@.B6a=H+d)?eKBa<:^GO8/N_?E1=0G)Nb^-8\A1\8C
\G)<0=J0F\;G.da>Z]:+]Z]@__:<0CWO<L[/M0YRW#K<O#fN2Qf_LgM/T6DY7YFG
)E;0I^V0PIB65aTR>PP:J<-FTd7[36_IaBZe^OI9IZf(H_8=ea>M7(6SJ>L,V#ce
>I]N4^JE89#>@:S\E[FK7.gE>,cf?@1Y);c/SACL19BZ^2c^0aT10/A_K^F6+^eM
Dd3RLL&A9OVNd=b3>=+b^T8>E1HHD][9bYPVX-]4B5aD<3=[^D;IYJF]BPG;DL@C
Y[R-609_L3cZa<d]MV@:;=?>g/dVS]P0(=@f,S^BfFQ[79eF<]H;/bS;[2&c<J7+
G2MVU9M6KG]R#d/b1>?\-G,&9Q/4VK3K;;XG[#T^K2(O#6fMUESA.W?Aff_g>ZR4
QM47(8[8cZ;463U^MHL^XLIWadT5MK)VTJ&?&(eH@]GM<(UFZB_TM^4B=beX];7^
;:?CWfAc7WFGHb=>YRf]BHbHC8A,W+]5(\ZUX7]1W\YGIRcUWYO_^CO<Zb8G&eg&
S3aDUA-+_?90([fK+d,_B#3@(Jf4c\Zc]N:eXF=.fRfVC;=Gf<L>:GdMK[3cbC#Q
8Z183\9#495L#VBO5_/2KJcYC@^Y40RG0I[T#Y<W(R(-Wc<Ha+O&P<]&e9FX4.Vf
6b#EJf@B>>\SDY7:]YB)S=?83.0#?O5FVRZ&&<8e3:CQ^(Fg:H086/=g9;O(-C@O
M(a&P]/@)LZ(G/C&4#bNWV-52D/NV?9QLV=e(<Sf)_X#N78#<b-TREY9;DBe,]LK
K.ST8.Dgc;?PEZ<LH[W71A/8YTe9DQY#d_WMb=SV/HC1LbO>MHfEWV0VNI@5.QF<
7?^BX)829#+P,D.>N-H<:Y12#S)TA#MU&;,IY^E?KO;6A@[gJZX2/]Yc^#Gg2d,G
#O4a(V[,3ZPCGN;@:GG7f8,.P<#cLR5e\S&f[CY94W6RIIYbMW#e..O>Jg)GX<\0
HWUT&Z54eJ0Fd3;:U]973[B7SH^f8:&(Z/58[MAN+[#-37a[/_2#d6XeM>E&Td3F
FU,fO]0\\SNSNXWbXBd.RV@M+fT1+8>R/#eQIbP3@MM5TT>-@U_f(4gb<]6^L>\[
B=2H8T6+d8;UNcL56B=d]#EUQL)fIY[OJ9\C_>S##NEeUEfMeD;<g11<Z:F3.?dF
dLQ5KbFWUI/8E\5Q(B5eUSe8B,c&[X9Y9HZMXU>V_PMZF-IKWL.#X2=2GM?7O=f2
JSB[C\ZeSP0<O-5WfATFYK)S[\A(D=N?:Hd-R8]ZBfV;^FR]]NTgVYP)g];:80GE
MBQce:?aN-:V7&>E9PI/B4G2CD/8+Qaf7-9SW5=f2>.JE_HJ^>2XaK4_8SIgKc[^
]H;.4J[//YNc\aVfbI63?4-9=Ig@TY=@21A3P[-+S>Wd#@83MeA2U_+a0?-A@dZ5
+5@)MRKOG#A3d&L.0R.-EXHJHLOAe^L=U7CG[eT<6)H>H)?U.6M5@5<7\a.;]Xd-
c:WP<g=&ZWJ(7A)3DV]I>[Z\7+VEEb?RePIH0gFceF?QDLT#8?H70OedAU)X50ZF
.;QWH..93T;IFD99b.BU?QeSWL^L[,2&?,,F]5cN&EH4gb?<c+[.=\=O-?<,Tb&>
L)X2DB(MP\DeO4-T[,Ucd8HXJD@Ea;(LYJG/4gPW1S#JC<K34C.3[AaAN3?FM]?J
dLa_;J-BDSdD+G=,_0L?UV):-1bFU+BXSO6]3EK,C+&?[Vg@6.EH?(_8KT6P1e^M
W@0McZ4\RfOcE/NR5W.6=?^Zg=c1CWAc7N;83^P6cY+?0[0eb1J/\cT<ReeeG=I9
J4-6QN+.HVdM6H=I<X5K&L+5:Z[PC+II3Z[^W>^;d1c/CNH?E@X,-1cc?95_6OI.
K&eL(FJ+]HF@Lb02+X+9\1Id&XLEWf;-#:JF)9d3ADXNPMN[HO>X&Y4,BReIKJBK
9I[;84RRM<U=+VWHR38Y[>=Z6S\4B5CT1a6c5UN;J^)bSEfQ=WL<.DDJFX0/JM?:
2@e^4I?dg.=6ZO2)A2_(^2g0[2<7fdU&G^9/J^5\PD@BLKU==NFe<;7D;dEH2.LY
+@-@VGG/Q_]UJEEWX?NC\0YX2GUB)OW0E93<1P942;&64]QS+:,,\PO1<UO()-Qg
#FRJfDfFW1JU;.W5641+JCW75O,DgW3@AA5VLg;[8;#b>57<<29.Yg:#-=3F][:L
+A)T#RE:6KcC(c1DL?&(ZA>IXVIgPCSP=SFUDY,&=Qc0T]b1X(d&1=PJbNA?f2fX
\+8_HZB.4K&MeGK>APQc(#WC,d2K(O8=NY)\#K^6Hd5#W6HI._1ZETD8+C;1V\+[
8#1?X_2)C5RCXYTEN>@Q=GQ_Pf.[Fc3bb5?caCO5[<T(/+)(^7)BfS=GW;XLSVKZ
060SP^G/;MfRL\W0;SG:[L/-2BE9>KL6Y6aeD90J[DcNH93EIbPeFSU;92MM[5bf
[Y3S8-EYb9Q\(_QX?O7EMPZ=NI6[TM^]ESDb^FS#fCW+-AJW_V;d[eME59]H=.7?
YX7bJ(4RM)f?;@)KNXSECd;97JHAJa[gM\7&S:3Fc5K3SPD9XK>\UQ;2:OFYga4P
JZKYbTL>[gD)A&BT93Q;]+10DSfTY+&2bCF3Yb_3c)bDQagKR69&=.AIB3?I5JgI
F>]@1Q9T+d>\ANJfEKK6HaCI4GRId7bV,AB+U-?,,I^XdWfB1\TE>d6RJZG,#O85
9IH#-/WO#@12AOKJUJ2P\d?10eHIbVZ:;MU9CLB_LRH)N=[&9@VeCZB?Q?<3Z-WX
I)aO28L3?DUB/8V#PWQ(WaI-_cX(G3,7H_:f3_L87.F<7,be2=1PN71c6VM:1QJb
WM3b<a0.\^YC&Jb[BH-4AU>ALaPY31AUU10XIE(+X9>:E<cGTN(c.FZN:&GO_D(?
>Kf_RGQ-f6f0QT@+^L=H68+&G3>B=P-O2\KFN@,M5@BX^fRF#U?EH1eD.IUZSE9H
PM(5dQeOV2gDWc/;];EM;074:AJAWf3\U.#AP:M\2(9;Ab]GQY@/,#5c]HJ1WG;,
5K)+4E04(2:T04X1Jbe<=4)R3)EC>L+^>_=gHSe)(<5>O8HOWJYcCB96Oc(FC_M,
L<0efUF>b87\L]MU9E(&/a:JC+Wb2E?/5YdH@PJEV:29a7K/FCWZGW&a7+,,Q0/X
?-CYWUBZ+8XfYV7&<C:YJU.4K_0=M\Og7A\PGK=H4@Bd;+IBKS5,756XZH@R>ZHG
56?Ig9#;BU/,f&@ZPX#b^<[3/eABY/:C)6:,XA<>_c\gD]?MW)Eg,>[O3_[W^[K&
R[FZ1LKB=UD3.B4NJYCK[3REe=]Y;AJC8YC36(,JcN+,Z<fBT67.K2@AS:DP,?U;
V+0>B^6UcU9-U<)UL9R)FR^M+P(SG4G&0^-1]C8QULE1<@Qd^N5f?H/fAfTFP=81
(:eBBNc[#64LgQ:W;.T#eE]I4R:bWb6b3;J-]d]2d?W@,@.-IQZ_7T-)?]1394,5
3S@VF=+22XHL0NQ7GLEO-BAH38KJJ5UGC<;E4Y&1ILLYH&(P2X3GAI-Q_g97.,N[
-QPXTPT[C8AU5BFCX=(VCZ>O)\JFc-BLK7^OVG5G47OL(N@f4,HP9b@A[,Y>c996
UX=<2?cfFX_CG)cQ.<K[YD9.A#):b(g)(\T<ac[,RIVNbKJDLJ>C5QM,g9UZZP+R
AO-@&.RZH@G=#?B\QCH-:cLHO(#QddHBR=2>2UQ)R@)>+?:.E>-]O-U->,J1,=HW
8V.3F^ML+dGG.JURMQ5:VT/T81W8YH:)I;F\/QC#c,LU2WYdE;P,TW/6<fDg_IQP
O/^eM7eT\80Q4e\S4d<WcY9bf..XJ@8K#Xb;PFMd<d&Q[f235AEX3eG2-VAbV?#b
5&6EbgfYP-7Y?ZgJ1B>MdIg4[eT5BbL+;bHHX>TfRI(PB0#<&#;6U_a=1,F;NT?4
<Q#A=,eEQF76.Y/6Te5#38ZIX._Ka0gH;S?0L9L.gLSQ[8-P39WXZeb]#gO;T#4Z
4-(KO1fL<,UeOTWHF@QX9U<H570e5(bB<35+G2VA9+d#1GBe5bCS@cb#(79?_P95
U/N,TAf-TEZg?3<&0e^Q,P@Ac;:1OCEdEB\0(M5):H4D4NF]\:#KZPOFLE.OKL0^
((&1F:7\bP;M#:PXAf>@GcI=_&,MW4?7<Ef[_F0:9LF6/a89>=Z_f&Zc+D]gRYUS
gcd1cR-+_TGcfAf36;>+_W<G#U^;MIY;9]O30>1.DNb1]PW2Y?V][UW&6ARY(SJf
DF<F[H;H9@,QM2:dR\fef_-VXe+EUVG7C.\SbA9U&E]a=4K0Ye#(8UcbNf>-2S2V
@\33))]-]U@[3d?CU&2.E#AUQI>g99ITUYb2]SbLE-&_[K1CSN3-55Zg[H\-CCRE
UK6WYAMXMM=[_G[/^O(PT#AMdb,+ADEZgO;&TN+OR]O>94Y>A/;6b+^YU[DeIW.P
VcPECd<EfYfgSS\d/fb[@(F[<eWS3Y6YDdJU-e[W6ZEb(7?-0K<9@;@1fZ;3VOBZ
=PVG+SV.8SKg;SN7D6Q)?fQ)K1g_T8\HAa).T[\f&5HE/D=J7_-@E_+MW+Ze9RUO
87IeP+#30D03\^[_5^3.d:K>:GKDK6>_,EXP>^d9Vag?_#(\5DQW;I=E_:XM]<I=
PH-Z+9f9GF+C0(aOOGU.,^<Ka=LT;Y?O>RM/G&)&BMa;[dI@G&gK0:[1ed(QOBJD
IgIXA\T#^0C9cV];Wa4^E#R>XUa(1AP-FSK4@^@H]U]9fR1^KAVC5NXHA)FX&eFL
XQ/-6&JB&-4:_)2QJaL(;a9:((a\M[).W:+Q\g-+0<\?Ad,2[_71JUBI#HW;@<6H
^8[aL671W(JB0K1:I3;)N^FeGDJBR@PQ&0KB&eRZO@5@A7g#J3ORU,d/D_>feM=9
I\D3N7TC9#\KN6)\/VHOR(S]5+A#VdKLB4V#;R1D_5F5fKe^aUd5XT];#a36\@NQ
bH8B2_L(d@,_b4/0]J)Q64eP(Y+8;#S=OYV)XWRVfE=I2Z9N,LO0aI2&&]aBT#6c
(NK^Cd>]A6a]OI#T-+d>;DX_+FQ/RS\f.Laaa[DMQ]fe(1KO.Jc&;@)WHNF]:B[E
B;TWXV9-gS+HO+g(e(?C#+1+MI#fS?>?G\-Re+:<S/-\>Q]__U\RX#1LJWIE,EQB
eK7&X][aX6;c+KWBA-.cOfKg=A-@VKGBGJJ#S:U;<:^L(M5H,ROe-C;ZCY#@f0e7
WL8;faD)Z5M6b<:]>30#HT3A1O#UQd#:U/+AW(:#5dJg]a.4YEXQc(@&JQ^a4W5R
e&=gZ3)G>Vc_5L&(LF[e&T(1\d9]Lb?>AcZ5_Y)?S6f[e)eJ1?65NH?/;=K.T;BR
,BJHN;RQ>8_c>LN<P9/U=4)CF&bG)DaX+c3dC\Lc<:4c?ee<&Q7fA@P)Ee)<0aJ_
7-3dTI-a4D6@ZXZ_XG^3O&(\/:NTf^E_4b8E7aO[Ub7+V4S)6HR=8,g./+)7c4f&
L;+FG4[].8V](.;g.:T]KD;@c[2QFQ,[P-6R+:<KJf4EY,Q12^.K10E(aW4&=<dM
>8C_PCV3Yb/7@Efe6K=B=eCf4)a+KO&R1F&_G9#1b<3YD);)b:++&=+AagG4?IL@
c?&B@V<S9_f^aIX/0bL8]SLFN?Uf?Z/+9g88EEF=8bY=#eH=cT_f894V_3Y[(5@:
,<2O#X?SfLU;T]:M@6J4M52c+P2^:a7/OB,Sg-=?9B:>@4,ZVKOX>QO^)&5SMD(#
M?#a.Eb(]:/SVF0aJffXM?\O=HIIG;:#W(4bM4YAT=/GTD/07aE3QFNMWF:SML#W
DLeN;_aT?9Z8geT6RFACY&RGGd4<PQ<2BL03?#D;cMV/=U[;2D7RH.FB,0XW;X3]
IV\EJeK[>Vg^E@g<TZ.JS1IY93X],\V;WN&c/fTX>>C=JKXYffBA>8KUg(KQ8YW)
;5eb01N9CH+3:/8aRA;#RG.30;/^FCbU5HUYd+2Fd#NW@/:MAP9bOQ0N[UI2F+cX
-<-+f[a_ZU@QC+NEcC]82WXPVc2+R,Zf\H-T0OUDL;]>B<_ER3Q?.>T/.&#5-R.U
II:I#&;6>/+/JR9bNUQ<N83A-Y?g.>eA9#.L=[/?NXJ>.;_53AaWfd+HO@[9d&c#
EU?@^/#+^D+PMTBa0/3]T8P@L.3-H@.^HD13(Y,;#BfO_g^#5C,_&HKWQHfeSD-V
0c-EMb6?Q]V,c=_Df3^8,(&479M3F#fE.6K[5Ff2+\1UH.[Bg6@C<YY7BM_2@YE=
U_\=K2:QN^?2Z2G)V?LG3H&MSWf1dc\YY,C-SY;G?/I#.PY938F_f+BUOW52JU:M
-_XS(fJ;UZ(:O;d=5@@K@CgD>V#TVDJ6<H:QH#R^c@d2g-A^)MDCB1[9EH9&4EfL
(1MJ+6)gPY&.JAL@.adO[8Qd[)]K6eW1D_[&-Aa&L/b>>\?;GBXCd(0e+6eO=:Md
e0J6U0<A>X_34SU62OC+g5[0)<+PQ#A=5@M:bH7G+G8TaLYGDVR69PaHTYU^1Fe=
N\b,S_4F://Ld&;-BH[dSF<aaK0:LR^JT9#Q,(H4fG.]E[T[O\,=U>V&aWf84+95
V)094CeAC[A#b(T89YbZKaXE?Rc-L:M)e#?[XP\[&Q./#/@Y]W_;2MeW167cPT+I
?#>BLSOMJ(e<f5\DMf31\??Yad@X6+.W1>.)85T.11L&=Mf2>O&;@0FN_5_3Lae&
HOUDN)/RS>7Pd2P73Dca]B&fEPVD^80^6\:^9);+CbRda_QU3,/SW#]XF-04\)JK
HQ900C90d8-BPf2YYLLJG+J8bW0B]YW9U;CI4PW@=50ZP?,PG8<1U,2Y4ca2K_,8
9QV=C^11+GNa<G=F79#9)DXW=WT<<:a^?d#c..Seb;\DET@5VJS;BRQKW^Df=ZC=
M2&[dECVGQbQ(YNIHOO=(dMTgd50V[/&YPd0=MfQK+PQf\L&^9KTEgYU6Se:^PD6
[9(\<#P>BYD_:=FQ)=8e;5e1BS>,A3_7U)X[^F;G78.#b^@)2S;\0Y58=^3YHUb5
cV4WeSB_d&b?UK#M3db+@.D3?)-,)RH]NUCY>(&VN6IWe9fIce]H(V#d8EfVH/+1
P8\LdGBa/#6T[a:4gJN?S<D9+af1[I1-J>PR926Qc@7OIBfL8Y,0gHJ-dC@C[DdL
K,K4V=DNF&NM64D8Nc)6USE/F]R6fFf)3?B]7@:dOH+4gdg:)(7B+=A^O+@dZ.T(
1FXfL?Q4KTeJ;[eIO<E)8?AGYY^9Df<)@G3(ZC/K0]:&=(G(<-V5&=SCQG66MO6,
TD1R1O3;_IaLCKBQM>ge-]/SAV=+]bVed@cb6g?FYI/B.^3Y8gCb3?4U8Va>d-YC
9Rd387c)fbYH59dEB#)OWMeCDLgEVQeA=[2@NLIOeI1Q]+O4X@)faCN0_^.NN3_e
2)YX^ABd^#IdOO,N<bCC>dK(7##0)CPS.KWXHdSC-f//QTY4PZ.HTV>Ne#V74EPd
=C[9Bc&RZB2VKBQd.fW_4[If.]FHF([VZ0^,1gJO^N6<_Tg.f.N31V&0LJ/,5GF-
?gM5]V8Hc)/gd\Q\^M[Y4)F@O.1;RI[9CF\Jf]CObRcQ22/OUa9)]S.I6ePY.gZ+
_0GV-O&+HG)bKCcTG.YbQ\X27R#=STCL^E)e/6L;>cY)0CSG;GDS,OV,H\Kca58U
TE)NgNLB6&Y2L,+J#[4&5)U65J?5&B,;0Ve@cIaXH>:7+6YBW,<5.H7(RJ.]SfS^
[d3cX)8\(/YcCU.V[?C(J5O1R.LHGQQR_+@:?f@ZN)Y1RD<UOG.#e,M87cPMSO<K
V(.9>0AHXSZ./WY5HL8d^aG2Y;TaO0?7>ZN@@@6]Sd>/E#<3,S9_18fdHKc,<X7F
135SF,TN\X3UK:3ZAAEb=4122\:3>LH/?/B9XB>gP[51P:>9:3VI7,gHeXd(HT72
b/3:9-]bb];U<F:/&+VEVTXHIBcS2-JaUe.R<RMW1UE8CW-eTbD+-W9TASf[B(e9
8O#b-MA02GcC7:<QV84fN@Q44?@^571K-7/,MX(76#3T?@,C,J265d]U7+U=9K7[
+/W]0Pf\GLK7gg2H;Q\gD7\0X]-W5_U:EcGa?2RO(#3.1_:@X3-/F9aJN#.fX:ZI
<(NTSTIRC3^#N^,4-:>MJN^R2T==&?8H9?MT273-=TQ;L:HfK/[S/MB=5&1XKV^\
G]P+&U[)-8.Pb:F/)X_a0S/#?.TC<a>-M+/EYO^L[\bZAQ<OA,#<WgQDV,@,AGL/
;HHKX+F.[M[gFg0[RY++aEb.X8.2O[dPbS3/I2dX#&3bI1N?,;6T:^_L\KO#V[d@
:)5DJG]9F@\[4NPbOc_JL.JSe#9L0Zc.VO+7bZf0NF?]5&FQ;OS-UJ,W>J(XG;HC
[)a@eM)YF#F3,M60bEfT[U&L+gOcQWWJ42Fc#LC5/fZcWPUF[C\?][Ng]O(O[a82
=NK(,N?RT_JGH0#0_4.gC2QXXZ+bOC:[W#a:1.-6)QCJa;gD.;)Pd[0@XMBf<AV6
U;_6VfdF59)]?62G7_NgEG-IKT18<4HeIE;7@#Y_cPdDQ\/XV]#bQ/eDTBSMMKWP
B.bKQA.:^>^S0Q<JB,,=ebc=A-P6\BBDTYgX&9:(P<M@3g70f=XU:;aZ?-,UTAdS
TQR6+d2B+Hc=24)D?fcE2A,a?Lf?4OP6XIQT9Z1TD#c,\BN]:^1UM.&+AAX>:-XW
7694VKV:PNdF3H6)21?B&R=FZIMY?ON8:BY/S<3-#?[b\7WJ((&&;?_+IR7g,B3+
XB1#9L7=O.DE/3?,HN)SF[EA#D+UfS<9TFdKU37Z+?EI+TcAV&4JE7UTE3;]2(cL
6.4CK/=Z86P&V=76-+Oag-&37V8#+@QI&RDYg3QHKL_,\L=3BY(IA/4#XOM0Tg.,
MWPT<g:,RSeRKcUL?a,+-<JYc2)U/)eQX6B4;PObBMIa1E?<IBUfPCI>+MXE3Le[
:TZ;K2[7GcQ/O4O>1Ic7A>6e]DP1dS@dK:)0:++?N?9GCP9ZX/;>:e]DaMIWfNXU
XYE(O1XC_(K-bP],7^5JKDH5V+/Yb+F3\D;dB7S@<,gN#^cOgU72Q>KQ[/4]G]T]
UJ]:6U7fZ]>67_+ZaAC;#-;cD9W/a<fa^X@0@C,6?\>1cK^M.JdB5bPNdF:PC4]T
Fe+2A0&,31+:N0/ag3EOO207R.B+5bWJ1eF[BR.^N#;Sd)UL_QMW76Bg[bIH1SRS
AKETad>2\46GDGa:9\:66ILZV4VQ:K41cHa7EGQc4d_aEC?9^0fTP+P@5U#e\=-[
/GZ(K3\4A@YI#a]>4V=IK9V1>c(N3R1EF6(-IH[gU7/,/D_(#7K?PX1TCEAZVBU\
\gX+eQg/Q8RQK#b]1-.c@QBCeQV7C)OUXEEOB9(3aINGX@bUA/Og]CaIGF+^FXRI
g@8-GRXBM/?]Q#deb/NL7N79<EB==fAE-.R&FTcRgG.LLEH.;F4H4aU+?0I7J8LO
/)N^4FCV^0VUaD.8;Ya2.9E:;^_FRBdXMLBad&L5e,)I:47RYN<D^L)O)9C0EK\6
<KYHNU9;H1,C3ZZH?G48Gf</9(7@P>([BVEMS(ZcU1JJODF)^GVeDSBL#Z<a&PFC
=@^6OA]\Z)d2)51?8-4</f#?4H1GJ]/K27;)-#\XB\>X@b?^/\c#.F_B5#4/\(4C
fK0Z8M/XC-M7FUeOaSNN5^AI3c;O>62Q9g@^=gE/A]BcASVUU(?&+ZQ.3;),B7.+
_6-@EWOQ7W&@K.I#LEcB[1e.1Rd]M.E^#=U2aSVS^:CLaK#2>.gJVF.g@VHXT79;
27/07FZ>K20@307ELd48+JDTf8_@Vg#L.O3G)5/TIIQ?PY5YM\;,S)K;=7A\T/):
]ZPSO9BY+ccGTJY)JS&P2V^KHN]I9>#;QU0=0:+,e2K^5.U):>;N>BS?d9AQZ#UW
A3(E6HX;(A=V(2eP.<[IQ^M+00&SHC6-4-5THCKL&^HLVcZ^B,W62S#,9H0WS=VL
UD_(-[--3?g9b_b(5@.3GMb-E_^)F9BJW\+;b?-X3OJ^f3#J0Kbc_R\RVMO/NS@;
Qa[57<7=)[+</NQ>W0?7>+YD^TLfJK61a0)QX6):QLL47(@g:D1]XNf?224Y,5JT
a=ZQLSY6&B4XZGU_g3>M/gZKJ9[BDA<_;WHNV0<e@:6:D?c9X;DOPb#&dXRH8JaQ
,HMY@aNY6E1?72D(SgKgL<f8GR4#QU9]A_4G.@3Ja03&_CYEbLSH/Q8:-QBR#R/g
,2YcYeb3TTQ(D[M+X=WWaW@AFX=QE\ED)&HNDF);KJ]I2d[1Ub-I=]Z..>/^SWY4
D6dQ,N^.CI?dL#KQE/LM&[YP_b-PKI0^cM_Ta#/ce^NcDM3MOA?K+6g;.4P:53:#
\:MJO=QFC@Q3IHNP3-PCeX/1DJ9dNMZ(B6?;8JFMe-KD5IJKbPG/a\BF(5/5cHgG
gYLBeW>X>M@F7VF&aRRc^=NI--#QgQ1EF_(8=(F<THcbX_RJNY&<<^0^7_,3Ra9<
dMLTQbbZcT\Rc/->,15V^JdV4Le4.A]LD\F[B-]7aQe=_3[e5J\:?Ag7c;.3UHU8
A<([Y:)^U2EffP7.bO9We6SGO].UPO.>Q,NWA<(1<Ob<=E?JTJ=,B4Z/Lad2[Z&A
6^1\U?]2:bdMAAL(6T27;-NbQGeZT2?6^RX)9\=<Y[6\=]BN0eKe/+Q7@ZU4>/[g
>F2Ba@@U^\Q5Z)OacD,]L8N[HOQe81PI47_9+8dB8E0R0R/0<(YUYUX\D41;64P=
N5K9Ca5fYYF=KX+7,X2[32/2IQE/;C>R8(c0B^:1#B._ZYP(-c8eAVNJ_XK>_274
g>>VB<fe4g_&&=KPLJ3[a@>^+-g)F05c++.^M-/aU/ED^4=gQAWN.L^N24BT.J)[
+KXKBO[bMVeTU&,#GDb=N80O)g6D</?V>SDg+gb->4KSVY(5#&V)eV3?Z#08f/5]
_D8=72gDC&\Gg,MaHI@IW,5,HWM;WKFdVC(aQ/\OB38[0W(OU8-N6@<.><.Y):5/
]6^6/b@a^9HV6?_AdBY9;R[/L@P^b0L,1>5IS_?;bFH1gA\+/T63;b?(,1OY4bg:
Z<#=#Q\JObaJA0)&=BQ#O\RS3Q+D,B7EFXcE1P,6.6S2Y;;7[eU>RGU^67AR]#+W
J7b+(:^T3KA3R?^LHGN@H#MPdD5:S20A@<G1#\Z..e;-XP_25FG)SNd,OZ-,eE>I
SLR/0H88c[VIf[YVN]3Wfe>5&SF5aAMRKURd-Q;;]&_f,c)W11e6@(cg_H3f6@NV
,^=N.;8GE1d5TK^:ON<E:XWGTE;+\ET.F)2GX99W99/UBI5?E>bAO.U4-OD;MJ;P
9./M@fF8DTZOVP1\+X5eE4>,?:1W+]3Y)KBfNG_&TaY2SJcNdO)LW+dK038=Hb:2
T\8A/AI]AMNH2J[KUU._4Me>-CY9d.20>/S_8IHY1F3eGg486P6/SETF46.J<6\C
^+gC,LI3)4d>^@MDTbY-45AWFCJ_56^2RN)XEce>7?_8(PTTL)W^+&8<2M6Y2S]D
PMI0DR>&:^0C=/S>B_N-XgC)LY:aQa;,<+0:^A.TBFRGYORU1.J\BGHR_<GS#YTG
gUU9&eWMS9G?d[M\-G]O+.-XIbX\gfJ;653d[-SC4\I&8(]DNI^:<I=LS#TcNB_U
V&>SBd\O#YcI@gGYAQ3#L:CP+ddN+X_T]Q+A^9<cf=\MY4C1f[@73/,TQ>@Za&XA
=X?=N[##69M-TNEE&5;V]2UP]N;(+(7),YWCRdXTN<XdLIEe]-gLcXYFO(8b=[FD
U47CbR1@WaFAE.JGQ^U#44eFeHTXbXVQB)7YO7=;V-+)VX704=<R?WWC7WSg.OCF
bC>.\28C\0=MRYV3;V>#XV3C@+Q31VH+2cQ\F<C.5Xbb.ZX^<fb#6N5U;f5V.\[A
SF]cG4GFA8@AcKYfIR1:EW[c/K1F6K_[O((&4&T1=6\1W5D^030cPOSREY:dQcM&
RV;Be(>E4-24J_bF\DXDY@&V3,EeA&eTDI0]3#@<^N-68M<#C45A&a.@P(FM65+>
:81U4Q<8>V_/KK&aJdLK7.DUAD(cWY\A[K5]NYYO7D/PTDZ\_gT0+R[HVQ<1V/gS
cQJ9TSTE[fHY]<FL9H#0YGc03)P&B40d]P>J8@<Z66=fTQ-d8LVeRD2(]Wb17@[B
&a:@5V=2DZC:OWMB98&DOd^,W7T??XQG._CaWJH<cKfYIZ)OY1D.E2N#)CdL1X)/
6?N1/;8EX2>XYC,OO]/DNH>_Z9;eZL\N6NbOBM\3_LeE(K2Y&6adF6b,3-R\,Zg9
(S1\[#.5.f6R-C+.c9\g=_R>>Q.,E?QW[Ge7SJUe@/19f3)H+Q5[L4Z[[dS45;d4
/#+_]285>6,JI=Z-=;]CA>9XdG,HIKRGAcRAFO7Z>feI8c/05KIfDY;ZB7WB9C3+
QQ),)=D?<X@21]/[\&EX[:\IK\f+Y]A@5PFL])MO@G6_SgCOCX?<=I2ECW&3=BOB
./W8_Q&78L]L_C5OI;1^,^HeS-9<ZJ=He05,\Y9-8]TL=9:E[[Te#W<\+g4(FH[R
^0^BHB4)E)Y>bda?\1=T+_DTC[U?(^-FUHa\I<92a=07/dO.^eO,P/W+MT-.F3.P
2QVN?QA>_bG\Sf0X-ZWBGDXHSY#[d<EPFM@a^Tb1VEf,+/2T:=aVHXD^caK#-UR7
?EU]e(Z_4,:SN>.YPf#/FJCHQL]]8L#AQBU;/\e^-8d1#/NPa\@&\d62f:(2+d1#
@B^3TGg\OR^@_Fc,P5d)XD&fdb;=,?cB^-M_Y0b7]1F<55,E&XYQ@]WB22SJ#IRW
\Q+W+X2>I\]U6.6&;?4NUHZ+A9MPM;D5e,X_aQYMdUQeSfB>=X0JTCaSY+G1.bW<
SMBb)A.;<<A6P6],_DaI4#B.S._8)fN?eVS6L)4e==GNIG?f^F(T-URacgU#c]+,
Lb5/AfQIcCE,DL5:)+eG+3YBJ35P++gJIVDeGA__.71N1KM+.5-E+\X6DIC9^9@a
MZSCYc0@H&7)e_B+T]>>R^d]a.E4a^/X;e.6/Cc_MOMgVf>4Z]gXK-+KL)>I58d4
BUB33+^M<b]/NLOeH5<^94eL@34Y7Agcc?;8TfT+CTCPa97(g<E,<Y#_KTD0M3=d
M2I)T\a&;b.ZA+E=(N:Q6ZL-UH\QH(eK)-#?X(\_6#T2GI&TV<=ePQ?L:fQ7bVSJ
7I[Ad#5#&XX]2+>X8,0<K1c7aegM@b9R+,1=d-6EB21=Y/CKPYA]V0g.P0UY[a?4
gc_LV@\:=>Ic19;7-9,[(N.>cF0=3XS.UaAF;I[OK@cgPY_RDQU7T4C+^\3/PWA]
ZFRb?@5SF&JbHFF+eeMI\6#a\GcTDNM4IbPa-YS@9,2eN5)/:/X,&+<Sb.]>S##c
2BAdGEKdAeX-,e=?NTBI_]fDP2-;]^d]9\bdR_,TS/@_=f6CKI8P(VK--IM^@?03
Y>)/3TedBA7MI4_W../N7_3d3W()Z2<#=7U6^MFf(&N3/J@H<>&(0M#PIC2Z\9>1
CXg\KB1V8<1a[][Oe1UF6-6f_DXB1D7L_5K[cE\dD^[E43I_bQJC4[(V9_]+4(aC
)M:+X(FPCE>56;#(NP-M4CM<^38[d>O6f37X@^eHK(?I1(FE7<:BW3BA45IA>3U9
9,eV:GH8;H.CP,A5_LWGAcFZH(AO;[]ZKFMY^+U9M[F@&NOaa[N,VWN/.]D4UJ2M
J2MC.@P.cbG+:H1><-+AKD7WK?CNDDU6)Hd;F[g>gTDA^b6YJXXY0L+.6/dO&U-Y
F^ABeG=^ULbC>94aY.P&6XHbf[K[OSLUe<TQ5<8T\F]XSU)gU2STN(S#U0K9b8<c
QVacYQ1C,0>E_)]-2)V,.Kf38C^eE<);(V+@-TdX<cV5_6g,E_N),<7AM5_UbRV9
Q+aXXP2,^Fe\8P+0\=D50^8EPG&Df;N(^]=V:7K,FJSeZ81L:.d3;0/=b[C1XXgc
CL)9_TBf-H]b8)dSECV=WPTAOe/MCK:#cY07gNQ>LYK+6COWHIgVg\)MNGDW7Z@P
#<L60QAfWb]-3:>1UQ.aLHJA]dPAd9Ma66ER]9Ca,c/IUM7.#P5-J3>PDVF;IDF3
6.eUXP>@8a/MG:-:T]Q7/[?5_,Y&RIN1aHOEIM@Z9HA9MX09PISUX]/8QA11;=E)
g;WP.G96VY5LcKDWH4W(0?ceTE.>Z,R<9Ucc<9#R3J?.A[(5gR7<afKYO\^Gf;Ea
:X9D9V=@QAaZc6/T?,b0M.fY9W^H]XWGgVM\/1456W\bZF7=J6?RAfPREZX]Y7OJ
,US=P/_PEUJbO90\Q,C[P,R(,_H7?J/U0bg+PSUJ.?RD4PQ<@2Kg2@0gOfgET@GB
@YT.fcZCB9SPEYW4I>C/[9]DNM22QJ>-AG)\9OFaMD^4J?7NCAV5CSP6M+-e=Z.2
Z[^F7RDd9L+g?&:H2\RUIJ6ZU=W_#dGg:fM8f=PTYNVY4EZ</L=f,SPbIQ+DR7B4
4N.NIK9Paa/)ZAM1_8-=BKM&S_C@Z714W8D;#VOEg+e+GP@U9DD-N5J[]Q)+f9CF
Ddc6cX,UR20TDB]+L@8T0RE:..9J:&)UI3<JFWQ6@+]]3fZeGIDbfg_#b@c8HL?[
2TJB]4b+L_g2:bEBPJa\[cgB8S_2\+=c:43aU)FR)7\a+Z]H+d2AYbFUFT99S.4,
KF].f^98>5OZA<:1F=>UQEM+I-9=7]JT;E>D[W;C^A-25\E1YRT.A)#T.@4M)<f.
I6N8JMNDQLXJL&69\;)4=#M?:8]UQLM\K3IKCb[CKLe]g@91RH:@>2@eG#JfgJ<D
)7X?[ZFbQ-\fMU[d7eBLcfW-<9-0IRD\JeIJBf\VdC,BgU/5P^_70F:^(?YF^LNF
#Y-@40BW==-)JbG?Pfc:WW^X8C9@8M?]0c=2JF0:GFP3[?[P(fcV434IfRQ9]Q9U
-\N+=7VZ)+&O1GFbMFY&QR<Z0<[-Uf93KgEYEXXYBJNM7]a[Ka\?DS\D5.:d?NT_
.g6Y/-ME(N<Rg(HGXR^9H@aPXfF7E.\S#&C14FBe<b=1<aa?.3-E>D9>fe)^CPFK
YUg0+1F7VELNTb::TeEcZ5E@_MNW/L4?;=77R>:.WEfWR8?7)<._[9V3Ic^&gB14
\PcgbY1b--B;ZbI35:/;+DNL=K7B_VOSF\/MW8T,O3SQ.Ob<BXb5cbI@Y+56D8)c
ZE+FE&S=,/7YT1fYbaY.?QP:3EJTc8YO?R8;F(7#?>Y:8I&BAVH^FKPHT<Ca>.=2
ZW[[c_;Q]HNBGF3WAN.df.-OLbUM=.7:aZDZ&PA:1>QXWcGS;R^T&WX5VNK,GW(^
5OJ431/R-US\.\/2O_AVb#1ZR:(V)A6G;J_PUJ]P#b/38326[WY]8=HN;BCZM3-W
K^^52K+Ee7V+\SL&YNH+#V>HQI[eJ7PIKT[R/_c7VCPa)=9&BILH([ZO6,NM#J@M
S<6^Q)2P=&+[A,GL=DHCV@TQ;DX1F(O=+R\J[,&e(d\e#^XT4MbUIMOO^PV2R1@b
(?c3A#2///4bCWILS]:7UILT5]L3)RD/EAO/]?6WFbL^4Nb)HE>/^&X=e8O-BG]H
7ROc-OWM,.5@Ke>.A]ZdV^.AT=cgDcKI^W0_<:VBdBcb4T[FHS>:bCQeT\#QG]B\
Rc84_@@K[&4aCWU?E7[;>#,c)HB1(=@6X_cd0]?_Ma5VR3a,5O[([d[JK2A5(M:G
?)K,dWa:+1dLa(>G-1X_7+6<JH)MFULHU2MI:(O8g/:R5>;,L9gJUd=2E;;/F?.R
KPZ^Cf&,.0R1ZCCTfbL:A(Z>\O4cf01E/UdNE&2gAP#0<AEK,-UC^MMCe66]X)Lf
I;(0NLFI=A/S^7=E39RQ/2U^]E8=MUKb#Z2A.Z3+>;d(MVffT.=^YZd3+K?0Xf#:
JNOHPN<0)WEJeb,C,)c\5-FX+4A4;CVL&\?#dBC+K>:UU-,)?7(QOTa/GW+?9]VU
f7KCR.-J5/Q[\6Y9TZeR66S<]1[)b<I9>@>+-b0731BVRA&KFOSUU^d-A#?c=\bQ
TRR>b78Te,=:+4IWC#-\fPKHX^U[J4-2(>.MNJ>M5Ug+EB#J<((M_#AE8U6E<OBB
4-/Y._;&WRf)(6aY1)CQ].PVeU;BPb)c>FC?+DT\cFc:fWb^8V]B)OR:@L-Z031Q
NV3F7]G6;gTf@/L95\OANJD4e&cVBF;6&.dCERPY>83S[JAgXMGKEdC<S(QJJ(Nb
3YS(&-0([MTL62YgUgQ7U<MX\[B5<fWe;&_cO;3WI31E\1_K,6MU0cW0SU\HM5T#
UHG:1VR;g\(FN;:\Z,&VXP6O-LS-[>_/ZMET++F5\E0PdU=Fd4JR45D0[))XJ-;b
3B]g3#DUA:dQ;/#F4>RK2P347fcd@F7T/XLV6<2XCDED7TD4Wec)@P5W8C\/d07(
g)XPI]fe8H@JX,>S(K>NXHUE#G5AFC+E6cHTb&^B<gHQ[-9e5,_Id_ONY;#C]-XA
[+Ac<Vg_/c5<M6L+=f<=G4eP\S7M)f[@bNb;EgU7,;IF?\8HS:A1e7gTTeYK<+VL
2-aMS^GA<6HANX&c^?P>D#bHKB6fY#bCX<V#393))O&]YVJ;[5#HQf6_3g2G#C4E
f>2H<,_V/G&-C_5QYYPb#^<Id,6G2d[S^X<c<.=\;9O^f;1:)fa6_;Vgb8II-F)&
B6:[-59<<(aIZeM<dWO=<UVa>E.,AdFAY<06YBTNeC7UcSb7:NOVT]N?]OCY[aQX
E6bR1>EWSV(_eYOX4eRF(+A8,>LJL2Y#B/U[=-DJ531Z>B0^KAOIJ2JV-/d)Z\F?
^T7M0F+@T[T-.#T5T))@A383QQg3#fgE@3a<3UXWM[_)N3X9E/N(X[<4b3/_FWAW
(;,8@2>Q?G2&2:.NI]+GDAMR38ad,V/eTG,R3QT3:8A=VBTV&e1ZL0)>DU.;9)]0
UE6-9eX>I3ZA^M=3_GGF08V7NNaBBa),_=5\LBY<PR-Q930:_KYeJ)IQW13(#CG/
g-ZD#7V,B&#e3)dO7.H4\D#C3K]U[YN\B@A#FSU8>G;\=&0WL>L^G1@L+Q:gQgW^
^#QR]c]DJ&eZMLfB)WcG08CW+[d<4A<\T<A>0cQ32-H#6T>bYJL1;g&6,ZFWN=]4
D(>(/7^(eb7<JcTXXbWeO<+-<;FeA:1BN&M02fbEd\#eLM/NH:A)G-\FSZ.[_7+8
EZ>_ZgARGbY4Rg8ZM/<N+>FbJ;b]NR1e\\4DfaaTIHcBJZ_dH(Mb2a:>DX2;DBY=
_=ZFd.BJ15WB4g^6@9Q<5&?9S=WFZ\VDO8Ud?eBcegELSPA.IX<d)<U5=ad.1;CA
SH&MX;UAPJK;1:+YLXJ+X)e8]1dS]#1@.KFCe78b?9#9c8b4g=:T)X2=K)98bQF2
^):D5bXC>UQ-M&4@UA>NCdeeD3#QJb+5D47GCOIWbdO)/R0A=>(Oa;T7X:[dZ=SZ
WePPHR=(P@SRO3]dWA\Q/+g\[83M<)E-ae,KeS=1H@GG&XDUK:B3H(TfX\]DJ@;c
W12,1XP&,_@d0F_95/^DBE4Z0_+1J1cHH21b/)M[1NHP?P\9/g(>DcYdQa;dL?_2
+0]FeQ?=T#+/10Tg7X:^:2;B9UXYDV4VT:)H/(+SP^b]4X07PC@<&/?W\6@&CHg]
B,WRbM?55/AF6GUPM(...>dUTGQf)4T.E8@;A5J8bXP<+YB_N#5G5J7Q,L^81P[;
G@)&OI@WVKQJc<7U/&#LQM1(+THZZgD&Q.=?FL@A_\cIRGSU\ZQUGT\:c;(4XASd
,8>MPH?2R2ENE^/<>6Rg(JYKHDC&I1\>RJc2(IGbFgg@(\BMbGQRH-CD8PWB5JG#
N14](9[bHH^fbTG1ZJ1eaLIbL-#EDK[_Lc11RW0QU_fTHM<N2K?J9>eX;KK2D4Jf
:_8\^6>NVdcLKZA#J3=E5f_cPVcCCPaFfI<1]DI?a#f1HH^X=FW42=_4G38RACfG
F:H[\[D7.ca.Jb0E7dN[?(0W>6g(NdVMd=SgOCW7cD@e3W0YWU?Y)?_?C#>P=58e
PV34.?[F5gOZ,[E)(#Lc(&dU_5RYJ1dF@DYOdIQWB,^MJ3,HRL]Rg33(Jfg\RagD
]_:/Ub2QJc\&<fLKIBV[NU]S9TgJ7g6TA-5SL-I+c@TB35J&^;<7#Fb^Cda_B\:N
b^7C[+IBH_JPJJQc\cC/TYRe#]d2_5VPP;6Z/&I#[c<04gB01_=M[>I<]E9E[a(C
#P]/W5U11[OP_WX#(,&;QS=/S<I\dA/>e:RDKQTfGC=7LW-.(-eM;/QW2VUV80(M
Wf8ZaJ\6,NT>CGE2.1IZ-<4@8aI9D+U-U9ZbOXOYg[+5;ESR&Cg]P>B96H5O=_WM
cNe.FcdFCY_>XU/HUX1H;G^SVC#9Y4CK+@Ne(&_9<ZRJT:RINJEOMC.,RZYBF::g
3HJRW;)0)S=DGE3#BSfQX,T[P]Hc5D]R?)RaSg\#(?>71QDYJCA-BFe=Z<cEf^>=
gGfFYF9S_;eK[=>0>>gf=5<]&B1SC#a0JP6AO1:3U#7:^Z-0aIEX;<9<YaPL-Y2D
A8>2dUIQZAJ;K(_^_&;Z1:;HYUNC#=B2.L.6<3V#XaOV]0@RX+a=D;E.\B#(e(Pb
\5R>XL9)W4Bf.,PSe7Q#aJW\70eJbXYAT/^7^G3UW;,ZD5-JJ]6-XD/Cc#>dZ6Ta
_6_6R>bFbBWIIQ<Y2->G3GI(DW;Kd:-[/0GE:]&2B05L-28.6SKc>_@\[LE)^QOA
FfL-8K_-+UOQ,8#-/TE4)d:ffW#?2PZ7Vc1BGWVE)[9<0\bdBf),#2MS-IDadJ89
P&=:f<e&TGd\dZg?KE=@a35d=,QLV:ELP@2B,UUef]FXOfOQe<(1Qg[._IC-\>=-
fOYG)50C1#,C3SB.62cAa90SDO7aK?9YC.CX28)<]&XgS:OGW=][<?c\G?L24L+@
Se)SeA,>0O8L=RFGefJbIQ(=V;g:EbI>:Z0J.40b+P(7QTB8[D058adT32\P01,Y
.XTCG&G/F1QU@X1:0WQ/@ae##(^b]C?5[OLK6J<UQYZ/S16cKbHW9X?(dDE<+L6\
ePcH;G61cUT^)A/Y@G8SfOV6KCfCR+:RL[)4^eH4BdQ3=\_[I8&QUHZS\SUCJE.F
<3Z@R4A#^c7YJbc1(fa9Oa2(L1g6HRP>.H)G(RO#4Q=GSF=d+@HNCC/-B7f(YYe3
ZQOT\OTW.O7F7,:IG9(>+3?MF=(L=b>&J[0^VC3V[gZV(#>31M&FQ1;2=@+;P[+@
TX@L][?[.),X0MSLS/F,1<78)E-G=16__T67)7c7H856VYT8YA?_\aC/GL_.Hd:?
c];3F.9WXK4\cS.(MPCG<8#?,7Q?]TPGT]1_YOLb<.3[fDAc6M#^(8d161LK(6eO
&S\B6ZH?1E<ZKWV6Fd^d7DPWCRefC:I^IeK<LO?<9K\D)&>Y/.dFKY\NRSM4)cc?
F_g#>XG@MM>TDQ>+f6)M4N:<<;3fZ+K-^VC11JTAVIgB1=MdYK#H6dR_:&[DPJ0#
(R)g5FBOE-9T*$
`endprotected


`endif // GUARD_SVT_AHB_MASTER_AGENT_SV

