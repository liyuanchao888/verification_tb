
`ifndef GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV
`define GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV

typedef class svt_ahb_slave;

/** @cond PRIVATE */
// Note:
// This macro makes sure that hrdata is not driven beyond cfg.data_width.
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Sf1Mlmh0sLHfEiaQRHU4ddym6Sd86Wg9o9XYNaKHj7OlxfMnhRDEGDO3ffd48f/B
0HzfC742s87NVlxTkHNtPNuoOb+0ZGA3cOWPsJPk9oAMFs5uyqTpv9oFQ/e5jFMu
m2r5/hv6kpjYl+FS67xyvSQWhvVZNkeJ4QTkLlq7rBHsWng1cmmbGA==
//pragma protect end_key_block
//pragma protect digest_block
ZdHwrVL/b3iXOYI+xIjB97vBAeQ=
//pragma protect end_digest_block
//pragma protect data_block
ahlX60uABYvwus/nLZtt39XmDsull4/aWuFSwSzRWOHR5OEOCkuxfr142TYtXnaA
yhDpjMDEXipSgMkBZCdbAmLOuMCHajOeV/6BA2865k4+WQZJWqTtMho1aq2Fum1/
DjeDy17dXe609hwXwlOABpehroM9ZKiuqeyjaZ83pULwZ6JI3UhzwpsKFUD+sngG
GruImiZDomtt9hNQBhF/nTNVr663mtvSx3UI5P0iBxFQVjgsRHIS3LLGx9/wztNW
jBerabRnL9zGQoQyZTOI5F8M9tE3XAvDE15NRhU1zJ4F0g+3NEA5hy1ir2sQGmnL
e6ikkLu47RQeJYC0GYEEsJ9lnsoafV//iO30yqvvMby0EK5IWqsDV0g4S+IM2L9J
PojJ0KyZ734gesvu5JHC02/WbfhLyjsChOWmv5XHM18oItDdR8+gnahNaY4abuUb
WSbjxAtklzCUf8hBXxic22v9FO6WolxSRAzsbQHjiXI13uBc/kX0e73FkPjeRoAo
5R3cgMF+I8rUPeqDzLGDyMCaipq0Cr0/uwt/GEwvYlrkVWy5Sv35KzgH0PHF/tNY
E5jVOnqPBypvvrHwMgrIsRNFFFfcgq60/eJ/M+j3z8RBZK29+4uh5LvYYhmh8Zl0
PPBeNvdYDME2sQKfOa41FIbWpSmCpCrzhL8Cl6khc+X+ri/asGJADEiCi1OT1C1R
b1ttvWF6hs0C9s6xl5p1lg==
//pragma protect end_data_block
//pragma protect digest_block
qilQPsv252FWjbW3wCUrgnpXUDE=
//pragma protect end_digest_block
//pragma protect end_protected
 
/**
 * Defines the AHB slave active common code, implemented as a shell assistant
 * which basically just converts requests into VIP Model requests.
 */
class svt_ahb_slave_active_common#(type DRIVER_MP = virtual svt_ahb_slave_if.svt_ahb_slave_modport,
                                   type MONITOR_MP = virtual svt_ahb_slave_if.svt_ahb_monitor_modport,
                                   type DEBUG_MP = virtual svt_ahb_slave_if.svt_ahb_debug_modport)
  extends svt_ahb_slave_common#(MONITOR_MP, DEBUG_MP);


//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
yFP8wFwl8rIOqiw64P9vRRiGjw3NQRtm+IMTXuzhLC73MzkE4wdyYzd5RhrtzU6t
YgTWFGHOd1xLVGGJy2JXXQPtDmH+37Z/C871sb0/AXMNayAWwqOqxjEpy+BJIdWt
VlxHk16qeMbqPBI3J4nlauNOZUCLAgqNW4QuC3dn/FmtBeQQG6Aupw==
//pragma protect end_key_block
//pragma protect digest_block
LQT4ZX/MMmI78oucZz1IpYSac9Y=
//pragma protect end_digest_block
//pragma protect data_block
WZVaMxCk3HI6PuKYW7luoI3NFQy3Y23RTw+WHsq5YvBEy6D5yAWWejMEHQxtEqkR
DWPT8pgTMe19pOuXWzWr3pBW0n0mTJ2SoKO4MMIoNbWFij4Z2mNDudC/aYIEZsvv
iRlsHSq/ofQTu1/4HmDrGvIm7SDBx3yIWCbcdv1KHjRTs2Rnf0WzvzJVHz5O1oi/
BLSBkifIKdxMUYUQEHIY+wGnJpV4qroPoLw9exhmSaIxms/CypntOqtwRo7ejU94
Yscvvrli6irAsA1w0y6GK4dqiGHbWg57CWPAZtXlkQ81m367OJHkl8Eg/iHNjdCp
0inu6KrA/wKSnoaZjmGUEt0CgSGiEENOR6bYmbI2zHtx11JtE3lxdHJjML13edP6
n2qkZHO/w0UkSm9ti/rsdxbC4XW5iCwzD5Dib8FvJVZt65udHkDGgT11h7SZXGjX
lrX4xjrjxjv8NXmGYgUIo0Yw+THAgQOC/0z69+kbfJa4bNKeodZoUM3olcdqdlFI
9c21BVBOLe/xRCZMNLspUl6Od4vXT2+PeLTynw+EwZzp9fh6hSkWT7YyItBSZ7xT
4PmadI+AYEE2TDbDUDYytElP9gUujDQ6kqO8Plr3KTfZ8yjcbVu0uY5oD6VTBqpe
3vRwkXUC2mZo4Tkqwt+thScYG8w2560wYtbeswfG6gPTaTc7FxeA28bNo/95iWth
0geXh0cq+HBUz5XosHvACqBKU2xzqKOYgkLC6yf+zytJY/bLJ4Y5lIKBSPrfeqA7
n/zdS+oEHOIM7qLJxEZF46J8Q8eZzgtx68GS/p20lcArvRZRZptDt8iReSy9NrLm
uuDUmexXr/Hb2pdiCC6DxIKU5CRPZI6lBz4rFm9ZzZzwas9xfNuxWqYTLng5/vNC
5gENXmF4KzSO4ceaggxcK2yCM7OMICcxvLu0REMsJuL+z3Pqib6myiuuw98PUZDa
jjdL+YA4cGWLIG/zK5304tjVHA8Z0vaKkq3UKoXNZkYFcPXpkcB6YWx5PVceVs9n
XKPNAxxI5DkuXgCMb+Kj6ROChXLjGx6Z9wIrXY7Hhork+FLDyRLtMgcrlrGAJtXi
WGSuhHMB+0qcnJVBXehDliqDnlzHEdzWq9CtReDhZvmTmGYMHjFC5MA/2MH+YAR6
beRA7R88P0BXkeSodRpasq0aJ37tiyML3BAe3LZUdg77/Qk/RmjDrE/gUj8NzAQX
PEAP1DRVcLMFDUyNf4fOU6BRY1thJ7aF/QdcCCHE4I6C2C214x4eTaTN8nmL7PeH
Bz3WjaFFB39JEO78LKrYi1VjUkzR2dAlFgSr16IqUw8Y3I6xk6LmcUSbAws2o87v
YNCdvfTIXnL/+rOw16JkOHKDBWJK2RelSBXwVU18jO4VlF6nscFMyWLbiuKLlmxn
lzpHmY6m17zqWe7x508pLqRt776wGuN8x7KoeofxfxjEGzyiwm9DO5PmMfjUVIw6
SBY7hethn+Er8ux1gJJhZKLFMOEr/yX+GeL+tuVwYjyX1AuFU2mlW9sxUpDcHiPE
Tae/hpNLzlJcqmp0DMg87a6FEWkOu62+f1M603gnrdnYT9BwgpdrZJyOQOxN3qIi
ifaPaLA3gnUEdqgMk8IQw0crJjmHtaPe5RqjAnIRypqGtpf3xlz/MYAqGaPJSHr4
RqXIJ5+tWhvu5MqlRhZic20RUnGr5fNXsyHV/Nu+Z6S+yqBgUMhOnaGzlaYGI1t9
75ETzemPIFT4c5ASpnRYVvA/+ZJTEWebIcUXYqXZFky5df16jFyH9gVxbv/U6q4t
iiq1WO2EYDpYFTm2Ynlha2rNrCCjSK95Bwecs/wpNzJF1DeiZftWwhKjlep/h3J1
mSev8WwS+Uy2TVXmLt0NjIxnTAhtuSx5krlEU+SuT+Wt6ceEI1pmdgDGuiGldmx1
LxEntS7P44ow68k/MT5ML+UkpCr0dFP+fV+X8/KDwJ2LytWbtIL02lSsWjXJU2fQ
ahrSf/swcqEBR4ItAImVmBxfmvA9Y+KZECHcFdvM9jRAbH/NM77Kse6n1dDi+t51
KzXkylxGm7Fe8J2C/MDDIGp9o3GNuH8b6wZYV46/7oGWgoPI6DV1SSjh3Xg3jRBF
R0VkH1QhhaPFz/lnvp4glHFHruAR85KYg3b6G9teouFtGdQsrYKiBKgUy5r5wHme
3C6LIskv630+VnGmOF7pQe2n5HjidbM/vstLNY53h9CKOid83S3Yyras8uZl2hAt
Ox4mBiBOJeke2snxXeHpwEEfOaMbwkN6JigOaU9XEuLT/PBqGFaR17CV03M69vR9
qLc7AIR0ACRFnHP9cC5ryqt1edunw5TkmId18b+rGSdu9NGbZ75erwF7pNzxgB2D
87gCzlxiz2nAR0adbjBwdJuv+6BOxIKDSXNY0OsTbwmzhxuQedBzfEilZ/9U98gm
DNDF7u6NLkcu4X3vyLQYvX1UgKJ1nIbCl6gSbYMCrg+wUREKxgj1cPpjtEiuCa5d
SmSgXrGrCcR9fDVvebq49b2rJH79CwtChNzqLHvTgTNQ2FnxOl3lJv4/eAymbrkO
9k8oMHmfM1nsF3ZfIeM5Keaz/ykiHzJTogzevp2TP25yGgvkwW/xrXfxkc979Qmu
uG0t1V0wAPpe2atirI65EcldwS0Vd8VRfQ1fP7dnJ6Det7/5Gd9Uf/NFIDt8Qqqa
DUj1G1suB/IxngmI7vqttFnZINRgYlm7SLavZXTyT7+X7fNtD+ZEsnNM3aw71y6q
nkA3uU7WMo54tOkVFCGmYm7bnMq9hEZAVgX7E+zz3Z3Dufk7CMh/9gyqwVvozJq0
hW2dNY0fWI5VK2YVbff+2R4vE+AnaqfLP51aNWgEvmviasCEhFzR2TOMUr0UOS6T
ZO77zKdjfbN0oZTOMBir1EoqDbqDGiIL38EO2rsKMt1fCO9wyyeWSz3YeQTFJoDk
jBGNM5ndc3CmFuVI5ZbxLY9A3Spq7Lj18FXvqtLBUuctnIU6Ko+M/5z5SFOZ1t5a
8wjYjGGvfSCW9bONJFFtzU2yDUA7fvjYITw8Z0Aq0VoJtJ17d/fXNUEDqmW6XJJL
XG7Mwbeb2iL7ZVZcX+W3Xh1awCS7rSivLr8zMydmV+aKhJ+3/gNAA6mcnJU3GesK
Eyx2GL21ZSBZrrEkUZk8zBzskyHGlaH5o+kP/xvZwRIflYOczN98bmFW0QY1xW0y
8s7Wo1hzuIM55VWrU64lONh3e+2zJQvUh1pXZGPJ4S19uhcz2iURuBGpgC84Th6F
IakhlndZaHlb9sfa7BJxXTfdO7mLqI4IbJ4z2sLB/9TRlvEptIWkBQVVPTAKH0z0
ORvVBDJGGgSVoyx5mMlb3mA/YlrC0gf8q3Iw57CLUz+Gi7UtAHnINfF5l9Ayh6B4
jZzZlKi8rRWq1boPU2KOS3PDZZmWeyUlTk1XocSVmmw9Z1+q61h4JTjykxyuN8IO
GXKqlkNYoQkIxk4f8X0nGnPVoJVlimVg8iZ+wjsAeSUyiL3eftQCjVktK6RKyNzg
iAiinrrmktEPKoVM3pK17AAlxMIS6aNVjclxmuDMIFGDpmX8hItfWxGilcM842tG
Amjz1QaEJAukucdwNAmtdfkCjTe80U7Y27flQ6X8fu1gx8e6tda4x3pDUKcekA7v
yWAcA4wUkX03Loso+gpe164fe+2xU3USGgctoB5TQI7GtgrCbKYkdFxIKTVu8Rjj
8CE4oyCn5OU2YpEBTiiLzKX7A9N/NDQP3FPJdk740eB6yNeMJQ/C2JjuZ7Onl1q6
qRJTuXVMk/i+qkeqD95dkzVB6I9ogybvG/I/Q0OUfH/ngaMlCJ4y5b0cpGH/aO8N
ufTIkzPgnpkY4lNfU9DKeURtTpkdaG1vOkxilq1CLSXOj1JUqmWIKEJifsbblUN0
qiqpTb57py0ic3imrfTTK0ppQ2k0CKpajXuxu/uXw+fEOvfwDHALprcIbd1HRBO4
VYsKXDymbWUHJ5JNdbgE3tP+ZxeHPXu1mqlGEKHlypXTNReM+nTbTYpzBdLjSxmO
Ylj8y4keUoadPJDFyx1E9LKl/Ab5C0E+EOED3Fr8krS0a2ZItHAnzvjv4N63zugb
GqCzw4P1CaXjmqvgY5kVrfVvLdNhqOV2F6litOGpCchmpCI4Vgntt3GphPaKJbbP
0/s5dc2NjQz8pbLMCUuvICzVHA/YCTmJwZ9IJp62tENJEPLa/p8fCiHA4NL1uY24
unVFwbLgNRLq52vJf9zab2npMPoLStCjH1wB/jNY84G0fGjGOyk6AySi4tskPwMR
kkmRqToyVGB21x9c59BV/CiPmd+gaQGDpD2unVsNQDtPkLThYDGvK98AhHCo57uP
FTxRPXbQplSg49Hb+YxwMhsFcDA3SJ0y05fDRO/Erj6THaVvzxl3zrofi63EJ5kw
wjV5YC0n2cmZTodHCnqvFM9TZYhqR5LYdLP5d2DreR531lSjzFe+4w6mRYn1uxqq
CzCFI2Aw6CSy9LvCFpYOi2iH++Nn+2xKyOMvfIcQMLZ/GljuGFPWjveoR9Ei/C0H
RdAkm3BQapiSGmfe3Mc/VzQxUOsf3N11s/9BYqFI+0cV4eBzZkIvPadKAMlPKhMh
1/UElG0ir7NZrdpbrThYyOiWmW7TOj2z1v9kzqpaTZbXRl9WIodIaEkZ/1kDEPRD
fsJHgbqm4cUurB3ymVgPm1/QxREHQJ3oHsLadGs6aKofaqBcSeaAe3CpGZ5CIxXO
fExwoYI9Ylfnncg9c9DwN5fSW0jY786w+trFOXbJf918aVPdXlJOwWBXXzzBtDoF
0QtTlnQfunh6W3sry+grH7w8Iym0tCIlkFxaVX4y67q1BdHvrMCFwQG1KIL4N9dq
uQ0NA5YUUCLmquxfywrl5P31YBJrinie0BEQZATfieK9uJ62cPNqSTpl/KThzuT3
l6csypU02l5KjUwLDQnfrv+Z+OLgrYwvfUpZk6l7CFBAtcG2lkeiJ5TgJzbXREQO

//pragma protect end_data_block
//pragma protect digest_block
3JPOV1X4vy68V1WRmWreOgr5wIU=
//pragma protect end_digest_block
//pragma protect end_protected
endclass : svt_ahb_slave_active_common
/** @endcond */

//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Ivs1bNhYeywDMVRjjRwkbTkSsO+qtSqYlkStzxrNx8Z2pfls2DmrxA+FMrOcJLTj
FbTnYNy1s6bec9R4tKk1z7HP7HDs/IxJ80r1D6glD+g8lD1GdnQYrk//opKCmY5w
D/uWzG4xH3q6spphfdH3Ky5N4TSyR9Qdpvc28ZEuuDgT/C63b1CujQ==
//pragma protect end_key_block
//pragma protect digest_block
kfLukPC3GpQx9z8GbXtfZu7jpuI=
//pragma protect end_digest_block
//pragma protect data_block
si80c0Ec8376Wiu1iozgIDxTZFRl89N2kuBFT1BgiShxTMTic9inkctMyydHBAaF
uncCSSOXZxHl6FUHYf3/dlWETx0ntWJxWsF5e8cQmrDUkRjEId2rwS+Yf7cKQolE
ifGLRviR8HlnEZVZM5rWGD1ITjFG+l5wI1Pr5SV41VBjvcoc9SdToLNYjeQVndbd
cAqxfZ1SZf/0tfNS1A8TgTgkeS3TuUvwI5ACOi46t3nuYW887Fuu7z1IUgRYaeOo
Drouj+S27UAY7EboNrF+brGn71ZVUM/cU90uBBXctJbQHn8PBOc8Rttr7ZBvVzHU
pZMw/AL0civu2AQyjyvjjPCvz1cBTuTYMgJClAaGNB6CKgjPG/SH2t3CFGX2hXGX
1+Ebp7HEbGBD9m5Q6j9O+tR57iPumMu6mkzYgtPk9VTz8hcJg9Dn+bqhVggEoYMK
V4wPxt/a6BkWHieH+01SgMgjZ5QIYMIwlc9nYWYvCR2ilLLMZR+V5TqlZ5E5m1SA
5Cbv53kZahIV1JODTHBeeRqrzQ0t162OoIPMwZMhjFCFA7YdH8fjnFxzOvCPjVgu
8XxSFnjVQY5Bj6sIFbiQJJQEt+6Gy715TvxYghSRN9RqRwO9PP8bnUptZBtdOSAG
IsrjTCG4GI60DWooSRnL3RtcAyK0xeT8ZcG2hrmukcdHTSpoFizb8UarnUHhIt4q
KbZ+44zByDRT3WLbaixxOOaa5tTPaDzwrpW+7R4aa23IRRYOQ2QNCFkzsiy1toG6
ko9a1c+VvDtc1QlOayj0jgOrP8gHt9BS7IlZDTVDjFrWlXFTYV8Tnbr9oxaJwjZ6
y7lU1yDzxYjY9xtXpjU9XC0RCuGqcu+VjM8JxlNunAnk3TQrPgEQ38mWjvIMQgEI
d558l6BuayOK8wViT6m7Du0PV3YeUiIdwLW0BwhUL2mQJL0pTxmwO5fvSh/6kElW

//pragma protect end_data_block
//pragma protect digest_block
wGvY/BZsl2g+cq0uLLh5WuS4Htc=
//pragma protect end_digest_block
//pragma protect end_protected

// -----------------------------------------------------------------------------
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
tQ6TwRmu5DckiNmDqScuwkb9+/6qQnYw/UNvpD3fYlkX3fgv4cAZJat9tnJqt3IM
HNNItONS1DgVzWBCP7M/QrMuy93ro1+Ff8zWrxDgSxdNIIIjAPb2g5UxWxkbJrQT
lfGe0GNJpWVLnTokxUk7fNC+LJB8BSqZF8xmDxqIoFhS13TCDg5MTg==
//pragma protect end_key_block
//pragma protect digest_block
6XM1Pqo/CREpkKBD0PnJ+yqLJ2Y=
//pragma protect end_digest_block
//pragma protect data_block
VoWDsgJM+YQraQ/zdH8NjWMv7VHTeURlCJ0bbOoHjUgJI7OdoIvd6avjyVFGpZj0
kKgUQ9vurzb0tLyvb4a0C00WwpEJWp365lhReyCl7g9E68JIBEgW5rrvzkPi2XUr
J/3ZgcWbKlC97rWj6jJzzAmhvYS5X2ffLuZVKjpWDjzfs519si4tMoBHML7CtpfN
UPguyWZL2ZrdGTw+7hYsjkcwLvOJR1N8HhLWyE4fQTk3SffiuceZ2sXR3ZVrJFlc
047qoSdz8YR49c3BOHhH9GIHOGEt0XJNN35JS2+peLjBm8BWRZtOsEyhYRTtcEb8
qA7un9vGB0Hq9GkbfBygQo6xuXaHn7bBUwUoWuiYlctVr+FL/rLUBDA5XZKcEuXN
KUSPLcux8b/cb4whK/BeEObJaBfmmx1hvxlhb8NjGFjEp+oCF+BQOqpXcLpbFMxY
I1ED9LKUqJv5ffTehNpLMyTuLUUaIZ28cR3nYY9QU2okDQigyu4zmoJ9+DTRVfT8
4cUwIIJUhgkBAGVwPBItLCybnYqVxE+wB8KT419PkNpTmV5EZ0WzvEibozC+jnDd
hkTFx/FL7rcdXsvvMGFDDCGS8WJ1QiC218sV3IjE1QLolk3MA3vnUHPpQUOPqshb
i8CSSFHewtE3WmF43cPvTS74Wewm+bN2IRcXwp98xjGY0J+676fdVgLSkwXaRUbQ
JH2SqfCpur14IP3d4wPtX+bcN642BovQ8rIktL+WmyO3efYJ3L99+t2ETnXiuvbm
GkwUcL+RZxI1b3JixzEGA5dwlgez4kAezqtNaO2Jfmw4NqmqtJf+3/XeCn0KS/7w
gC+UFbfpgBz4rcTM8Q4kF+xtuPoVJAwNCydowWuzAzoyzkf6OAp1W/fHRYvNLKds
QBoGzl4qjVu6wQSMuWV72EZTCr3QKEhjnycBKMdOmjtBs5vuUkEwBPtBixXjszUB
IQV1K+jVeixDnpR9OCk8CceQtMmRxwfEy6yORHnq5b0jf7AQkg0D54dteJkWKuZt
orcRcUeE34O4CtAPV0m2QpqHUpeP7tUoF3ssuzBaS7nmvJWDXKKnij5pZUwAuKuI
TGsQ99EvpXFYNBlJoLeW+ZlWo+eCjqWDQNgjczYOJCQiiKn7nY1ue8XTJIsL/Aix
ioKhyOnjaJ9MoqQxZHrbaTL4JPSyEwmO8s804RF6MfCNBYWZXVIoZV2hmLoTGyhU
0BzPXQ+sBr18qSQlUjed00ydQ1bvHdyRTm3+hL1Ql6RaQvcUE6wd3XkWHiXT7s6l
YUkLiqMCiY2hiphn6nQnPpGio19LGy1aOKhb1k9BGJNu4XYR9aRjrycjoUe20rtm
EJtrwDglWIHsc7OmgIgRBUIxMrFSPQSMVX3Fv1vOxpe9eWZPWn68pDFN7t/Ujyeu
d7uaIwyIBlx4fi2Lc4LuztOxdynbnsv/xayR6GWf35wfQUJ/Dxyhp6K9PNVqf8Zl
mCx70sUy/rENlJWquLxdlr81PsPMZRFde9D+qTJO0nNkyigM2HBa9y+c5sBRZvHd
qyxjC4CkWRKotK5+2eXRiMXOHNVpENXjYK2cRugh8+GwRIgpfKdAcWRW5U/TSgpl
kBNfvEwVlMpNpHt70iGUovdcZg8St0urm3PdoYuV5/kohTxiy3MogInUaqwpyaqZ
4ibhNqO0FVax51F++Fxe3a7SWdPz0tozLoUVx0gTP7GNMT4DtFCCZw64oVsUfHJK
nvm1MFO1zWarXq33jgHu4Q5u6zw2VP1KjEtKJ0ZzvJbrt+Lg1mhqc3BAC3n8XBey
OP2FJhBorZilLW4ouOdzSMcLp/Cod0PrgAfWCq7R0ce+Q24ImN6bRlRWzingDb/N
N31Ab01IRiYSBViE/OGzlJ3QKm0iQQXM1Kf3wN/9FyFDEWXVRmFXGBdJWYOMlAu4
y6Phx8gBDfMLu7Y+U31iK+4UBkEdCyEd0OiW24c4sj9MewJsWGtHriuIjkBFhFgP
zjqpKOBTwXNMy5+6YWt2WU8Rt3UYL2PeL5kTLAnPZob+MOpbzy52/iDleJslhRbV
DXaF71QnOQLCAAxkxuy8912Pa3L2tPhJgD7LRpmEaeNP+fG9u94xT9yDoeQeeXRj
1QERVT0BO02wg2hhqgO19I7Sh0WteVL/lI3DxE5Y5FYcmsaviXCOZi5uEZCi0jmx

//pragma protect end_data_block
//pragma protect digest_block
J7QDckyt4elWrkuM2jubBNyKUuk=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
XHFQr6469f6LoqKiU+Hy84e+YqQaIZS7zgIks0gMmh+y/8NOVdGBV1Ihi4tlbOYc
DdVDjOd/HuuBYaNH+UZc500Xo5OZv/4bVmnxUxGJNJYU1k+ZBc+RtoIieSibOECj
/aig+uAn9aPLGHJUBmcVEBLuF2QtcikyhDM5RgEpo4uDBV6CtJkfKg==
//pragma protect end_key_block
//pragma protect digest_block
isMPOqGvp4/5uT9AXaToQmSlOmU=
//pragma protect end_digest_block
//pragma protect data_block
B2JR9YpJ9Puj2xrRwtDUmC7hVR+tN6/5GffsdOiITsf0/vnVA7YtpmqvS312Eceu
/m4NFxMp9Hm7NIhHfzTF2Tuo7rqthV9+xTOrQJevpCz80zYWwH4c3vuXeXYpa/cp
qg2be+wM0IA2Pllxc93Wx2TaTal0/YXSkdXADRzORhsNkFRu8Hn4uHp4wByWikd+
6u6QfHmjraVTl1PCV2PlcQC7VyTNVKZMuchf9jX7k/uGWVq5p2lJaXcLTERZah7V
9EJ+ySgYVMqa9KPErC5/mUAHkp/emwyQHYD3B2sthKFG2PTMGOrpNGNzucbS1yDd
1zxr6POZfrYYYLeIYtlpCwAFTTWs+RGMMMFA9J6k++uCBZ0VA2YdT0gEy1WTrWKU

//pragma protect end_data_block
//pragma protect digest_block
Pk7eHWC3V7tWSAQANwx75M8H/PE=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
EvqT677fw8zXZboFFh8ITXWE9vU/Dd7QvLOOk2goN53yFj/InoSukZ3ymhzEIqna
WIxg31j3j51SXTz+RMYTHU5QQT5FV5oL01Rxisec5CNNzwBPXmfMNXscmyBUXgZ5
EcH75w/uQclaCh0jYXqigM8ASDrULjESiRBUtJACBdJDjoLFYoTGPA==
//pragma protect end_key_block
//pragma protect digest_block
73q+zpi05gn5X632AXVNpSYCosk=
//pragma protect end_digest_block
//pragma protect data_block
SEq26d8F3nuzkmN4qYgcOXmFu8qy1RbfKjxkKwdguiA6/+9Rpw5+KA2jkkzK1JeB
OZk0nHId4ycdBoMzQsqYVff/PCsEkxbh/dDSw/SYitYccgO7EjwT/By9N9KK8xyH
fak6EPxVd+ZNHrSOO7O5j/7ab6LoTcAszXHwrmyze0TAtae7yMEeM4FYCTiRTX7p
l/SEMyYMB0j8kzWiAMudnL9haFezKLzfXmduLcUZXQo8t1LUdw9gkNpfRuwPWI6g
QsVG/UV9pEdtvKljea1uX9iDB+6zRUyutSzhzac35fRKbi1Mbq95fp1GKdw1vVhx
NwuCk+ECND5qxwslZhXn9dfS0zbXTXydlbrGPfNnsXYgfHqkmDBVW8+/jjhA/Rug
prEalMdc1EevLRUDb4IyKYWUqc8AdFIcmsohS3x+JQXu/DQc6WDwEo/iWmtwngO5
7dkc2O9+jqowSCZfJFIELtF0xToOXvoeshcXHH96UXhRzrI7U0ZPddUE+mAZGYPm
7f1Qse9/mVmgiNqrQhFenzeWER++ou8ZdYJh+t5EHKzySrwbKRV4tlifdDpqfNEW
vPC8aIaofothdLDQagDTW+/1KAQ1MTxCraH6xxnFdUBI+WmFxCy8/BKEwufGdumf
V0ApDYz5+ZWXN0B1vaGFIOf0jkwX/Npzl09O11gJFez2RtpZOQfZTXMODkkrvS7P
gxzyPj397zDrnYEW0k1cqWiXS5X7QJyffcz7hR7KmBTWA9L0c9hlVDo5rRyOn2nC
R9OPNuRlx+iZc5YW/7aJpXPadaoef/Ye2ONBw95DT6bS29F7ZJkpEcx26R+C8MYk
UV8s2nIh2g30FFky4HaSU1dSBSr30vTR+t4quejdnH51+9CfT+hrdtrlrk9x41ad
owYl15F1bY0HbpUas8PB+/th0Kav5RHeVX+/+B3POMrDjUNI5TCHv8FPryVvBTrh
1+RCfe7EemYoRxcYFWVWT0xKUYZFKUJa9eH7jufu5x0g5J5v3xwSWg9Qsd8/7Z/P
J4zQ9hLJ1RbVvDdhLs6jyp53KxNo5VZKw0ptGqNsDiJdllyi5s4vSnM8J5DNBY+V
wtjsXyPLLYaWiK+lExHGPqhgRdnPpAyCgta/rBt7WK3+dDsybrw8HA00utuctc+e
8oELaIXqPh8HopfHrSApWBBR3b1UNqRU5UHOHv2tkLKmpwYMfN90132dGGu2YgZx
Zgkq5mOUIz6tUXlMkJzZabKtzwZD38A1sJImGny5/EmXm7j3XXo82emLEyBTSodz
ip4seI3n/581XxkKkmzjWF09X3nhhPXiwD3+9RrU5T3XMvWcUufLwhbqpcDhZAkG
aN0XEsFxss9NuIm6vFur1vH3kA5xNEwNKEhL0h8HY2llGiPlHyML0GE6iitdnTCe
Lx4yAD8lyFLUF55l3wPJ8C7yW8Q6BwWlNXWwpsJ87qYDaWqlHJHZgagADrmo2AXC
vMH2PDL5b6XQGuEDLm879naUjiRyUZtYP8I/pyEoN39QHeUdILVcUmVD+Djm59Dm
le0dYXqDM1Sdm1z0HYXMhu2G5yashtqh7DW4hVq/+3DYtG1OM81xVTXrimgpJNIo
QptvBAM/JTIHEGXadkfyqetPKCNTRXLAqcqpLo9Lp9M1+3LndaSKql9gn6k/OboT
ODez1cEfZcLx8BXyOL/q5iNE5QfH5uYGYpyQ9WBN5yYs7iPiGqrdvNIvAkrEVCqZ
iIuVyw8fgRJHlqxPWghMKGSLyW7OY25zu5M8tJsm11aeAv/zyI7XbH98VyWm1k4v
kqbNXb6G/U3/0HdIxQSkc1tlhxqx6xCrRQull8+qcxT4bePIkWg4NymfDLH2/Id2
Z12FRpsrmZ/oRQFtGyNjfbG3XPn0uQtjEGyDG+ZqfQhzFDQ/Q+B9qXsqbM9iFsUG
zaiWWmh9EZZz8K4c1Y0/UdhnRYyeGuWa5tL4xBB06+7jSdYKAILkbOZ8wrTP68BW
0QTbmh7hq4O4t/m4eiVubMY71m05oPQNMMmuFwWILOzKWhZILa/5H0y8NPh5KKA6
CazQnmlc/Apga5hjPQ78XTM6wok3+rTDtJl0SbnlRBxWZ2ysj7wopYwr8EbOuj/S
IggyO9q1zL24wz7Ii+1uO+SHKiKun7LWT50i297csZD+DhHu4960mNVs37Gs3aNd
QswoGThb9Q5rJGfWv5vW/D6DpOkMlErpvzv+KOEuwEFOUWWCJ4VRWgIYv9AdG3eA
xNEeU76SycyrIDq6PH1xWkdGlDRak27yaVKkzHiOOENb0OcVorr2MnXlXeJlHXl5
gVljonSPi48EiirLGE8NH505Ygoe6RRZYziFLjdW0tgtBcZfUIv94vEXq8wQAOH4
uVlwcBGT86pSt02UbyhXhLoyqn3Rct4UTSYn3hiLts7SMOh8LF28CqoSIXDQijDn
f9MWxt8kwAHu0DhWKxIAUEow4p+cm57YrD+DKXJesxi/z5PCUdF3KDwEVZKjykzk
IZmSMBsuB4CTeUh0E9FYehpewPPXv1FhfTEqonbl+xOTo7d0nRoVW6nRkgOihcKy
3FfPxqVfrAmHZKjWRR9Dz3sxQd+7T8xn783Dij0S3o654Xtstc1h9aKNzVyODxP+
Oa5gW7Ep5q7xRC9dRSXiTG8kBe06LhaQvZ903JDS3PmjgM3RA7n6WWLUi7jVt3qr
kqccZvytm8xcREqD+3XVrIbByUfwz20dmEVLgUGD3qU9aCeIQHy+qjJ0rpDpySkP
BkqoUmxotXE9sEu9+AyyYhaY5c9wXpRFaXaX80sVTrQy/yaV+DdysA7gYWabO/NL
Mq+Pat0UGfxx/O8IgujZVohZgvZJkCY+afQdVMNdCsuB3ynScyyBiZ4gEKZFUIDd
E42Xd1O//OIJtglzBzYMRIclSxZQm1B946FJmUs8DEZFm9NQfWkT2ntG7rHuJuvm
+/Qxh2psmqaA2RD9u5ywxVbLCpyUlZ6kyMwKYZf8FUGV3+ITSjJpHUc/qL5lwESk
1iZy1/TKNlkVbTYkuZKDC5mhLsURrlyKFKiBj4Jg6lx5dO1Q+L560mo2fd/yLvuL
z45tueAAW39PzRHXeR0NEqYkXNoa1P/A00maKdf+3QJDJRb5ax3E2vq2lQjeTdBe
PY8VsHCVMNc4ouC3JHDBp+MsLjyA2WNpPMNYIjRy8PySd8LAGLIcIqXXIiLFaA/l
4BHilymqt53wtrwG6Vr4rhHiGPBfOYDLNf3RFjqpWjNM38kpuyqQeFSUdRaEtifK
L0iBrAyXjvZvubt6TxMRqFB7E/b/389LBYor9Jz+ofbsSkuq+wANtKO3QEEPkKM9
5CHdeLtEyhASI0hv7Gey8RnwUCiez5ZTjxhelwVw3Wk8DIdisliG6TXFCymvWwxJ
nq3hxDMyfhqeXWeXWtFw56Qy/j/bJHPhZDXVrZd2nlzHITg2luyFwArh94Ed0hje
qdPRGjH8WEKgrFrhlpntNRi7+SiSt9zKSyKzfg2EpPD0hvv058Mml4xAXKOKF+jt
aJK67MexBF4ydWI7ejgFXkK0DaMgT+NLpzZn5LhhgOQODCsEk2tr5JIQH18eqbXN
tgggnArXpTrPNWY1XuP901GMPMJpaKdeYU5flsGg0//825siyxW6YRZaqGW7SO5a
uD2VHFl41oSTMkmfD/0iHcB9pTEU0N/NT6hwB5ExDMLjT6vGeQ9lOXgFfWI9Yfhl
lsk71iCseQWDpgz1MlDiKM++GfoCANALTC7blf+DRwS6NJDbly45odvDXipxS0OZ
+fkmXk3LCe2dxmO15Kf2pzYVm9wcXw7LVNpbX+1KYIJYDJ/HfPZgzPZoqti9Wuec
4akMdOQW3/lMUoTabCIYeC553yKc6OlgN3BYpR5LKnIzE7kunAyDooc3XefH8JGJ
2hbeQstXSwrNoxgHOsmKfmQ+ZcDafHwRiYaf9DKv+PXV5Rx2u4eNFo2HOcyP2aMq
6avnaib7uaNiaPvYbSJOKipQDmlX1dxNpccrmGiJZTi7Li5aLGNTYdkn6QoZ+7cJ
ceGKqopoca3yB/KfFX98cwPkzR38PeC/kyu0hEW4oEwICzYAJlLuEEsfhmo96Mqv
bZbBpy8KO/3Q1e/H5e6l525k7Isz5E8Ub5+YZ4x4slzDfBP6Zd4w2LrORWVDEWDg
arWon1FNgN329yfo0PsOBCM3EVyyEqlZP2woe3uJd1L9GVCJ1w7s8B+pnvCuYLHY
RFu7HHrMYXJ8cRDIutMnBucnJ/FbU2aZpdxCIJ9auD72zYYFqjvhgzprcY9lpr9F
lFJjKUpAgrWZzFoIOb/12jEwSDF89iJV3XkWkz0PaaWv9e40HUqtlvlzdCElCWEe
ohykD+94xVwISx1nvhJiuOLKUGDFn+5HXqDstwhEgI94xGetCLrUCll8wiuSkj6F
h8jYHeWQ5SWelBCt5LIQYRWF7VdG2WoGT/iVIwp4guS7YEQZHrRe2WnoY2VT9Ksy
4ZFj/rQhWfh0Z8ORJXXS9Qoljk8dqtdyaZi/MOnlOSUDRQ2KoKyqkR7HkpxDKqtd
E2kJHbQfYEbnnyR5j3fDyZyVZTdef+tcmQQWTWoGFgDlbu5E2frQ1JjMWBmrF2Qz
qzoKwfNdig4tVQnBMVYqo0c9iGajchCs++iSU4TpaNprYfh1IF8LCT4+MlrCWo+R
9mFrxkrL/8wwQCbTQhXQF4nCTxGtd8oJXIxa7GqSz9XXz2Lpqvgm3QMrf5jQWWYE
Lm/a8e3yOl7gX3OmHc4ZjipKdIc/VwYVTQvlGhU2tQGSCL7XxhE8il28fORRBnuJ
PTAsNnLgQAsaF6aAFZbeO6CWumlDgPwVLKqVF0OrPao8JYPWRWLnpeJDZ48B73pC
H0dOueosGPkYRhRDFks+M1Ch8dKqjp1WVla2nZi14FbhYXKZgZqAxy/5vhprcNNd
fYrsH9clPcmFH0pUYfU88YzKz7ZS2sxobXXwsC+PQczFpQWYQtQzQEGscACILmfA
Em+nGuuvbRrBNLlmPaVjqsZeRQujWH3ikWgtb2hhAg94mFfOCoX6k8whxJ5+fG2O
HFCJ9z0n6dtw7hiMpRMhFZ24X24+z5FRViJN9zNUo2rLreDNiJyhssRMDd0i928O
tG2vJeUGa6MR0quCmbUWNOXVnF9WmWtqo7sdgmWcBoFeT/NhtbF28jtXpV64j3n3
nDo0uVcws1cE5nS2zv4vEeDlavZ3DTG1cCB+YeNmnCaxXFTaif9OnZHG7pDrXgBF
sRIYXkQz5Xfjlk7z6U1zcWyXhu8pzIvPVKlKRdEXKfAOrhGa0lEZBANqb0pe/4/Z
ZZ2cXVqIFRsbEEt/Ny3irry/zI97UF9QnpIvxbT26Plf5dUPCKTvwwYYya3xo4hQ
tbTHH1q7OV2lfe+kEtTSfTAdh5CRKJK5fN/xWP7pO1W0oioTlEz8aPuWdboiEizj
i7+CJYhF5vqOkGXYTTZPTznBHaTJ9wsHU7DTs41xHpl6CGsDePclmJCtN5W//qFa
nQiYml0OptcufPl/C60JOreoDYAE94hvYkPtdfxM0qcYiQAqCtUedc52MNfFJxxF
atxYX5r5elhSBMujGRmRgZjjrEO0VaZK96x90oB+WTniXWGpnFZZRoki1zeZ8n0U
ybPCquEUQBfT9pzgMbIGGjWdEAnn5vInaQXe0ICNUPsI0gNBIsWd3kKj0BaF49M9
cdbZcJNozaTPkFbce1PbIlREdHFe147NP5n9X325lP/EzcojsiaanZp37XPbwV57
D/I8rLOC4Ra6c9wlEFPB0eUBzimZPevcomL/0CHJG41VNVAuqbgByFwkoqQrOwqm
WgJaw5K6195UZgptQW0w7hoKhZT6H/+6EQCz6avf/IfOrURCbq1s3SlZbcB7H67n
v7eN6MZsJJ4ZE88E96qqI6X+rCkAy8i0xCDwC6IayxpBWbWwmwj5alU/b1VmYc73
zh+Z/mumxiQHVADgNn0yB8LSA61eqGn6dS2uJUd36ipdzFJWIQMnY+pL1lkBVYP4
fVGYdWYdZq6ypYBpvBDw1efFPRL+SrlbvDv7U2MkGx6J28J/exB8NYRN8OrJii15
PX4qcFxaCt5NiPMMrVIH8QOKmKlNj6lWVfqVdicm6OpC1c2NzZ7kNNAg+4XC/njQ
o/aQq8vc/9sm98c+AEVmFZmK9wD9zl4Ha5dVcoE2d/o4i9O7NN9wwnfnmAlcatYy
sPMrf27urcgNuE8TA5Xe5sr4zZFdslSA2AG9GUCMiVRlj2ujlwLygcJ+8dSQhvEY
Y3ZXOOR8d0/rq3STtcO2T+4TM8FU4CwariLdSbr0YVkCjZdQXSFxzsTBjwceND9k
xfovfzWUxOnAbI8grlV6v3gITba397hDvEfLrasWx9ZkPmhMv2EI8tcAklA93uvT
53xwLEyyQMMCxmdoEIUHVjidPmGhFxX9t6LOHamN0UOu/+C5WXhL3UlOi7QNeQrK
ba5THg0y0woaCKv7RqPRosn90achUjdiChUsIwTJW1+QfBjQbNRIP1YeGIBiY1TI
uboZ7N4M32uNQ+OEBpqSoAOnS80rpvutU52rPDXTOiyBjhkSP2nJq0cEmvQEatFc
vz4p6IssYyaDdlADR5y9NobnW4hWLPwPHI2RAWU7oPfMmxBx+gMlivvqTgRuugDj
59eRK37+lwDnHB0WzTpkpASrFAz2HkIzog+3XJY+CT+sORgYvbH1LhsRs9dtJB3z
8n2bhN9AtMd18gcFbr3J/9iUeOtsVlGVAMxrAyrQx/MmmTQ6nxtHklOOeJ9N2OxI
RrbrL6r6etzvGq4CJ3dcp/9Mk6vUSmBBtL90Y2Yxd0Vr6ifEW3Jv18fi6/RaIvoZ
N8Tdgx84BbDtypfbeLruCszkzRtcR8YdPn33F8ViWy8du+5UU7q3UDwDbaGm7cV1
izbz3c12OeBtS/WOpPdBgrMU3U0kdLDcjUaFvzPgSXr51YE4oQuGyxMt9Oai2EXf
ZPu2nK6l5mPdkgb0KaRyew1OO3PPDcMZNl0XlU5pYldNqqL2yU8z8FYFWwxvgmAO
Zpch6EAWhUvTUMgvf72RuFBfqDTPdVSufsmIfIJ6npqilqwyMpEWHOziGiiJMp92
K4z6oSmsoUQrSOE+841UBatFS3pRX3MBza9QreRDvDhdbXS01fLUnsVCwe7m4ktn
rf81548klHQsqjeJwJfLyU5cOfrOfEuk944i80Ua08ACJWU3DiAr3D+XP/KYo9KP
EZXQLqiRzYP+tA3yKDb0N506cQ64G2u8UDETANV3pLHCdnrEl0Vj0LIfJ7a+Oj7S
wgl99cxujqkM1xIBBfGWFBZnSTwWp4AVBf0nbshR5OMUITIVmj3fGt2IcOF6+0ZI
AIFIvhQuVzEzVAABh1fzoasamfmFFDFneTSX3T8O2F2l/U24awPJECoA4lcSL38M
6+uMCLGhpjfvGBS0BXl8ghfvwuHnPy74HqHiztFeNZ0QIPxiyz9+iZQLsMl3betV
yBhgLuQPqkUoQ3zJh8zWWHDbw2qv7zgWZZosYMFtDtr7oIAcv12MOWX9zgs8TLw+
FOzvoNpN+1NZEYRUtt5SE87pn2NFjZaI4ndEUsaepxghhBbf/fwiYBpm+AO9ocUE
wiKkrbFhaIK5dbalx8igjS919a/mAirS6ecuIOQJZ1lai5AXQI8KxoR3ME04ONgm
jts4elol43Oyy6crgSCzx96m2KIe9qEvfogi4z4BL1xl3N03zb5SLOsfrFKJOPYS
Jk3FACujBCmk/pp8RVgNBSCYy9LrkM2lq1POX4ZVQk22IycS9wcyuvKLroKGxVD9
vZeNkv+SaW98Myc+WjLEXFpr2G3MoDhBe+gJs/UZuhFSTvhxK20uWKg6P2/sd4PG
/jO5g3Kf4SovzToq+INwGLt43MQTcqu0g+UBc6lbv1ONpPzFX34kobJeabppwTaI
OrV1jTJRm6sGjKWa4aRIamrbiQYwPfTj+FfzFg2mU6bE2x/BEYXbXCFCLtGOI+Pj
Zjt8ZKxtDWunxSBV/IokcnKAmuc5tRMxglLYuMPD+ihthSj5Jb59PNrvmShZxUWg
rXa2oxtfNTwfQ8KL6adu6i3k+cIzRDzZIa/pj7S4ZN5UuyTMVS8UUJTy26xK7i1O
qLO6qiZqvZ0VmLk7471XKsDoaCXoa0GmYf30GJ8EuKBkIydLYwhiy7JW8PAF3Gay
FE7d6A79/vwRfHbvt3vpEm6pbMCVsTsJwVQ2Y++Gqh4gKyZXwP06CoPCnBd8IQCh
4ANn73v7P7XDCc88WYVQ7fP2rx6rjdTDd7m+uLL1RVjhw56zrDOIeXLxLuDv2Psi
2o8BBry3ttlpO81TZMip8Bmgq0H326vwB0Np/OFMU5Q88NXC+lQ7j0MZgi9EeIfQ
nuiWjv5N6h61TOC0QOe8ZkePcC5PSLq2XpNqFxR34gFBp0Mjxi2Bt9ICohO4QiNY
rGdgTj8vZLz9Qq+LVQA0SZT/2JM3ICwcvfvtpVAxq8/a37CTPqS01J4/+xc+3VUh
GFwT3llFJDc6Ug+O6R+lCec7dwJyza1t2Corw0z07v8SD17zz2hCppzoRhspvoj7
HE30K2ezpBukIxaqTIe4jSSUA2SQsxKqvCL5egHI5WBeIHXV0m7R59mzt0JM60xl
jXTuoCW4ptJRF3I4qv/VjqULK2voe9jcrz8CzGp07UG9KiytaP6vG1jwLmrOSND2
xY52GC4tpSwr10F0fmQ9fLcZSYSqMcGL84tgXyo81UqH+O8wsaBtSzMSkJq5/tFP
eGLDHxMhzseHi7OE1kqkWwBoExGNXtFzoqHlAh/+aPG+IVOu9QwKs6UsFiac9zf2
5+PSLl0VBP5TJpxHJhTsdnFJrYyGvJaS62SGsgB9G52fcc/bZBptlci/FEIMfyaY
w2A9G+VgLbUR0mMZn7VKTtTegUjsxXSg7impu1HMnzSQjubu+wwfjAiTIZQe9IU+
+9Te55cqJ6lsI0YhWI+tGTMEpGNvVIzmJwCTw1tKKlF2FT50VE5GP6sbfCXm2I5u
33viDftN1bmnqNSwWcMV1Q8Uz/6RO1wBcR2Lg0mNdOEb0MLuWy9EmptuJ7Z7NjJL
OlYGPPPPNkjbUOm7mc42wSkK3EMDs3C+Y15XYHX4XNR81Zh5gCjTDhef59/gWvUt
S87rLCnI5XuT7pvW5RscPSHmuCmIacAUwvhQZyOKE3SZgyMPyYPPlmU+yXa4U1Yi
NuXbrgyU32JP12qBvNPeYMiFQ33/yXtOBLGzDFZIdHL6/KWe1G+4P48QNSBI+j5M
+nKWJKQ/AFPutq2ahe23cKL3+ou3S5LyvbOirDOESbG4+gfoJZGijuBTmNc3OEUa
CZw5MontLhpvia8ct5OUBHksJ1Fz5XQ4C8MVkPg7oP6AyVHtP2GaG1dHyOmhvFU/
vyQqi7Or8gVmfSH3ecG1Abn1itxZTYSycTYelirrQ5jfvzlpy7teG9HmLkCFBOTt
ntTKESukv9OkDQP0wwSLLyzzK/gxSFrw5dgMLSdKh2Hh8WxAPpQKmfXYL6hmp993
9OLwsxyKA8bhR+JX5uJNP/ZY4Sqlp+Ku73ZQGFjVpokIq0SHphBev/fYPDqUgryn
Stb4YuNqSj2asV2U+EPzUZQfa97J2C2wXxPNWQG8wKmD6rxuN89aSuU7IamFm9cW
nHdCt23gSpa4jSVpfJ9KrEUCwsVLKwFQ5IQwK22UoKhy8C2PCF1glfHkl0jXOiGm
HWOr9YsmP0jD8i4KpoMmI4DrwAIJeJXMzsKRuWZSgZxrqQH932IUT5O4Cb5l70gi
pcojrKKw1ehH7VPK7J32OKrPTfqa9oalC6S7WU6Kzeg5MsWR4Ef/yamV5lJDIpHT
ZF7vGu9yOP/Qw5hGl344uD9RroTa84Jt2GNOG/EAYTvibi7Ldoxbbhk9997Qnl2A
PhhE4rLYmtlV0UfFq3XzBE9uETTB0KO5fYBHqYTpenDcgHLxVGupJp6/hFnSvD5v
QS2/ZCD4tzrFa0kI1AXxcV8275KudQfIJWqFpZp8n6ohGaoUBDNCJc8yrQ9D5Yz/
t+og2rQZ3Cw9ntBd77jzVmYSh7VtWOSxRH5W+mBdrR1AiXDPeuMQI/ZeFUc+rTjL
+w+o0CdFX6B1ie5BQK/VOcZz5eW3Y5+TY2M6RXt4KsF3rZhAb4CJyTkUBPPUqv9m
eGYcH7NBAKkUNGdC7ZEioCUMmg56wCsXmCGguJRioxrccbTdpOhHkNnwdfM2PGTv
MmUOUo7dMV2FDufrAFRDeFz9Qx4/FVCG4JdxwbJTIfqrudHf8iiE5+cksaeznhIR
tdX864lxUVDCbBydSRnK8A/rZu7AQ3JczPq5QibfJ1kCCZOKnm5T0b1WkHAhn5bm
Zvm/orUyuUeQnkQJXVWXm3MnGGKbWmiD1sqA0/UbV66DGHvWocP8YF3BMGgWI65+
Skem3d4zSXG2XMFqHO8cDOD+ptQQCVOtZvMH7bd2AB5YuJ0BJ5+5miag4LsfYQog
Oe6KCoB78jJ47cZEbUO9EUtabmYy47aAWiT3ARyxYMTIiZIAogPEBpWoMenFSxsa
iM98/eDFjH3yWXAk9NyCLhVK9vgfJ3PU9Jk1B6SC8fSj8jxQeUlw9JKfh0571c7B
DhV3vpbfeNT0VvY1z+4jOjgPkR/5TScn95UfNJBEQSVeECDtRlOb+N3BGdHxZ4Ph
a3pMgxIqQIxMRkAI7L/hcyFOWTCw+4F1dpNTXfhbeOWQk5Dwj5rcuL1ijzNtqm1U
So7nCVhB0sCSQmQiypM1T0A9+1SgUIQJaZk32vEXcdfZensTtS5SmbbiDoXeyfgS
EVET7lO+YxO6Ve/ZQXbDItwnWvAWEoTJn90FY0Rt6OfOy53jLBCY7uHrPLdGKDbP
EsOfZafsY5syG4F5SWOEGHz8uWXrF+rf9iCUy/UaR/c6uJ9CLTZF6lwJBJihJj35
yCxyDs0Af55y9o1WQ1Fmjd8zXfN0dQtwLtttfxEsIFs+6tvAft4cY0/4Rp3Tj5Fm
SWrpkm+sxo8f9wRL/In7VQAZNsn1hgIMRupZ0hGYmW55ht/XpKmTNr0VLBuyyvmI
C699Y3AXcGobod/V3BwC3H/2SEqFkyCnStDkVC0qRzGsd1UubaBN16ItXfEZboja
FIK5p3udKrXBsVWJyIvKP4YmDo11jXCox8tSRl1UqMAVj8MZKAuyohT0Uz9kAdOL
Esb15yjmVwdJ7Z6F+5H886ZZhj/TrjuNvrtM9NYzb+z/jCjimjDPqiEnGtjtexLN
/0eRTPBKoXWadblpTPwM/TQGCxnZ792xAc+BsVNgOosAFTRQoamXYQeuQvNZIJjS
rhXMDAiRI9BqCNDZPKcXUgE0IB7vl0bDsHPoalanXpguhOX52qn4WG9GGTx+J+TM
EbxIfnZyDii0k/RjITy8VecgbVhh4e2cYFG2+zxJBkGE96u7AzCkZWy+/MxzZ73p
iLCgo5CAJxq0+47BBRn+9bktemGbaJ9V/OTiyJSLD30EctE9rYaceAfwOwm/vVqD
TB2/65HYdmuhk03naQl1zfrA1JNN1ZonxsWvwdogQM2vifjM1G30f037bj7dS9Rq
RqxqTbZaXpk/xabWSvzfqiIqd3buLR0raib6iVMnqJlaFUDKNCquvKRd9vlvJLEl
NDuVw5DapB7SSnWfRur0mAMPlU18mSwGtW7t4Ngmsx/bNOybzarQpupIiYmiayOR
cLVc1HOHoZhFVAQev7ttntFBMiYgx2eh4VZwcbbwxezVrEiOTh387TxE1QrfrnJ6
MbQV0JlhKieocnGTZ7YwovmNOGojEQO8rBtRUhsiIK1o+RkYN/VraQ1yyohhDkjL
Maq4sHs8+WjR7VXMgen3eTSgntBzzxeK09xe5J6E8TYBu2ZwzFfofDtMHcezOPmy
z372yLSEOs/SBltvJPaKLECCGlR3OC6Sh/UCnpxgAmEmbC8GmE6Tdsv978JYliEp
4mfsFW4+BXTgVJSD8XhGFf+rM9UfEq6uPWZPuOEEh7/xaNJxAMFopJLdUv3VCv9X
MtVGaphOQSrw/utdL9xYXTYHKvcQ1KWv9MJ1Zk6ZlH3/0xgpl/bs/5CLEHpGwHxf
NXWsSnP+lrVI++o3NqO25PNxEBPDFAoKfVNTQCJpIk47FIzTQ9jevpsgsTS55NlQ
jPnZdIfvza9Agoi2pNk4sJgB6QsWHPmj30BVvLu8mW+K5gTLrd+HIQQtZisMRzZM
Lu5dNuHaAeoBf5iVJZHYO3DgL+YZzhi6YsMmHPLytsEVUiYUgoi6zogdV1sMnkw4
3OZu3FjTAHNeevx5uMh3rf4T/cAH8OWmGcjHQPYAkIpU8IwmFJExEP28AAuB55QV
8O2HSskXBJIMyqebaBYGsWI7ItEuOg/XGt5SIJyvTjqOUy95n692+nsW0I69MYmx
XbqWjQGN1VAik0t9803qv6O/+ZQXyfH1NLErDa4UHb58WTU2szTAI2lUpM4DOVHe
D4vYSsxqZfwdrkT1dO2SAFhYQHuDnTdmSIZsBK8Dl7Yef1V2IGuNqatU85hrY7ee
Tbs61BpVZ5uAWsDhDk0iay2GHRoXzUFyrHNVtNNkYkCi0ImYZNsPYkOpb3NbtS7O
9XC5gJAM8kLbXKwx/KMtUVkd87S7jmNSrpiiDxbULdqMAzyCMRrW0txtumWxLlo8
JaohWLeIvXDJlEDNudPNj/enWFmYTkr85ypudgN0gQMzEVEHSwqBIlo+5Cha/zE4
TCSO1S5LXmVkAVZFnYLgX/9nXBv14ZTcqClPn3vSlvoD5OI2YyQzzaHD82J9bdq9
VfDUfD1Ue/sOmLkjl7nsmdsy31A3gpABRzKaA8davf891KFNYslsnHe4dkc8A/bi
a+lLZ56xJETQjktFYDCRbn4jCRGgiFTdlH3k44L5TMqsF9/+nqOPk7PxiG7nsaho
+IXqfDgGzXB9YlYtUIsUUpyktTuazPGFvEQzL1AScm7IK7KvwOVv7d74pZBVkScV
S5u8J7qZpjFxxqGNqI4WVDNc3ZGyAv5O10J9R55wdLgWfOKD+sS/DopTTwGwPEi9
HDPd/V2mR1f5WfeHGvGdMxIiLsAHQJ292QHErxGnLxWEeWvmAK1LgiT+sY0VuFT2
23E9WurTYmdJT4LN4lZBdW87mbH+MVpI6rYle5OVUtPzBCUi+OJWhP41FCAmUwEy
WUJ+qkUuqKv0YeJTyw6GAEke/rT0Tt0TA9cpVLEEfdq7Y/TdAhNWSq9GIreYAzQ7
REmFzhp43gNVGOzvZsjIuIAWYKAiGlrwJwut9M+TyM5yPh3ld35kJ/ClvuEjwTV2
i5SdiX+k9HQeIAATMLFDigPiSTcUePGJr7YjpFSpakANMz/QagaxvrL90FqB2xq+
V0/uCM5kaovPjTcm4QCdJR17bLtcmXaC0RDQt2OgYzWZrdjVOkdvbCvVFaDfAqq6
LLbcm0oBO2T+m9amMSIslkfNC5R67wl3EdflHQD/1vifaJBbucagrzSw82kbpfYb
DIu3UDNyifdIochLq/LyedtkYSvghPQaLEgCOhUj29wQidu/hCGdcOW/hQM8fAnT
N6BUOWLiYFsBzdUV3KWnNe/5xBZBYVw0ty3M+UtQPweIm+MdILOW2nXMZGEppWmI
eHkE5xcD9NdqADHahlTv5+Xa2nzM5O2d9DGWa9E5a3CaYLvMUrpEQKnGE7+ao0J6
4wTzaNkuM/N3ji54fjLVheMv5pBNIIXHV4Lf6Y+/Va++cu4o/HKJzy3HdTdUMnNU
0+giTkZ5+mD3fB/U+DiVR+4j1yl5H0lRoVnjDp4AyQPKDohMurYB9O5ksQuw4DU4
FkAQF/6219+q0pHuU9OvSbaisQGs/vMPuCrfIlGR7jAX8LZqQ0yFCm8wzMC+s+mm
SV/9e3bLCipRCVwi7+//a2xBWp7Fw63wGxAmy+/YOS5R14pRMa2M3OFvMH/ASazl
oeO86GVFqke4eoX4JHyzO2+LcEiPcxUFYXoEHRumOGT2eOLH6gee8I6E9/mD2hSN
NHX1HcZI0jLhjtneuiW1saSMDoi4SiHB/GnfjI4I3rJO0AhjzhhYDy6UU79ZRuf2
UfG7PPnmSj0xTMB+CLJgRw8lG3AwuGTkQ3EDLkiGqzXQgdxybOKiwKO2Aj7ir8Tb
DSan3TVhlgD+CjBqWqz6MFTYxLDmsqBPExbhnwpZ/5u8/VNGWKxpO8YtVYCuWzpi
mj0V2EzxpLzXgDiAZ2lMZGC9OlBqaC6TsCQNN4pSQ9/YX3FL3l4u7xIhjoC81NCh
ln3LHiioC5DbkTFZmpXlN3ZsTJU/sgnpY1Ce03lwDNuxL2kYw3c/5koxRZPtTn0x
XOV8+FvXezubDRpBlsGBrZZMh2KZ5C9dXQrCJlZzd+4E9HHSOr1Zlp+zXwaTZz71
e9riLHO/kVMMOmY1gRB0iC82xgq8QPWoY+FefztFEHJCBTa4SOgNmXHFGWk/up4/
HpFNQDvwZFg6gm2qCiXiLoLwJn5PUzRFeGuLJeWY5VoWTeWydar4yS9vYZcq4mWN
6KD6Oosm0IBJN4GdosfX6/t9r5dzx9d3PND9w/+3YVLPJdQLMNcA+hUIcOF+Gwh8
k21pDuoq6ucVCshjXAdGW6YOtpe9STxVZdxCJUBZnKPBXHTBFBM5uBjY8Qvv+Ruy
gjaNC4emfFU9UcDwokdPvKDJiZIRTJpVg87LdonGFgDvr6LzVzmilxOto8raNh0w
I4xCPZ96dlGM7Hhiw+6HpYEENqLe7gqIKTAsPkw2Gnxm2HIGhzoONrLRnTP1sYY9
zpPglLdkKmvaKBjMlbRZyT5hlVW17vdy4mK7ZBtMS/lggStlsKcNnU4Fslzfs/Om
ux5Igd3sqXpk3eNRKEBlBDcnX8bECGfbnxkwPbte6f4R3Wp0z68htuK8gYKJnrIz
ZpBBVI3R4L3h4+HkXyKwfD47RlmOYK00F5nUMBs6E4TVCqpZE6es0z6cDnp7Q7xj
fmXHDHPj7WFQa8traeKq5qzlDXUMWjQFocioOi0TyyJ1PZvDJ0NL92bZW6JOKJBM
OhPn4/Pz/eN/wr+tv0r8EB7qjahiD7XOQHjPRYjgILWYQRkWrr+fgi/g/h3qV3Bb
oIaGT7OoXxC2eaDBlDm8swoGsIhb5/Wy7qNtqBGGrr2zby+3RuVCzYsVGYEBoFnX
KsGq+RseQqfldIlwkWUudNbg+5aKQJQT9kTEkYwtuzPA5PmPX2dGHXGpt/P7570Q
SB8aKT0Aj7H7LmafUmTGMcY+BRYERAFNKoanXXH7XKX/re/dYv7Guw0VRuRm5SBw
Zvj2i3ouxDpuSnk6dTVm5i/v8iqXSsq0MfWXaRRvcnwmwZCRCqlgo32zjyhc8Exx
10O2y6c94HFrmKJIgdOaGq/HtiEAvHm5/NxvjNYcl96UyB9GCfiQRGtqq7rZGWcB
//qoaCqR9Lv262NVvABP825+A+yKgcfqAjeLqu6yVg/LSPz1/cp7/lnKsi1VzHZ2
ejO0YbUxD6NERkp85Oyhx/5hjhZA6gCQN6xFlzTEMGeiIulQj/T1Iw0oeEARLpQ3
RlOjqM5Pzz1D+2ERw9j/1IV6T7FFr5AjM7j9YbwjOcTcStHWNVfJOPqQnMjegyHz
VJ1SnFon0Z8F7l7qn81PlAemDb1RiZiR2utzw3NRDR1l4A1MjA2mQK7qNC+Jaif6
kx/GSv165TolR/hh6ain1CVnelzJ1atCCiRTYdsgLuCnqVjkBAZNPC8w5A4EMaZs
F0lfegeLsQEtCTo16Jq815LsQAESup+D/IaX+jE8r9IMCfM9iZ1Y/oOiQkxFjsjQ
ZDP6hPmuP25ySWqEnjYrt9emhyYHYc51+at4PPYCOPQL+PeA7EU2/uDK6klmDnJA
qoklIFvJ376P6PF88mVOSSy4MhBeenmYt+xwsoeU5AwnkhNKw3dPbPKbSGb/5NoK
PURJVriKe7GlpqFkLr8JQeRkSyAHZ2VsCqi+MYmYwfVx1IGb6KZrWALT2nUJpamZ
3G1cKV/Twwr3XFW2X/oCN2IhdI7Zs2KUCrTJKmV64rZRDPR8zcj9tpgUxdWBGjaI
XmlU7iqcmjTnSZ3TzBqg17WYJTLo1W8MLguhwDTN79F1wE6nXufYE5d8ZXFeXUL9
WNU4tnQThDZvCnDKhLm58ntR6AdqhWmLMcQvfK6ixb+VPk7GlEwQeJCFX13wqbiG
gbqtojEwZMha+JU/Usd+4IK1M8dowIB7Gq4/G6M2yEfSUMOpJAObzSdaF+YO+ZC2
XpCxQ4BYqxGTOfZ0/+HGOmn9gD5A7jQ+NpuVB+q/VIXQYkrA/q3Gc59BB/qOZATG
mlp8EV7TPnhXoKevTIbol6v7XNpTkbNliXzr//ALqyu2qt/KUvAFvBapgVErnfXf
PAJisN9BjNsrmRc0OkIeWer8qSQX5JxiVEjMblKWwEwspOgGwenT+bstpJ5S3F1n
V8tBoOC2XkuZNiCIQVioOVuKReAE6gkR7S0ZGEQ8avBc2vHE/EQJ7hJ2Wht+4O5+
LZKHp2VSJI0q9FKhaLKX6nv78kKdJGrjN4H1hfXizdhMYSXWVW/jA/UO6/ycj2mm
uB2iy3XtCJLLYuAbklzcOwndtQn1uual5AVgg+QXbJN0kWJUtcKB8/wdLICVs0Mp
JYBK6psOJd7Z0JU1Mdf+hUxq4xBOOogMm/CPZAjkTgMOrUFHFw1Uzg6T5auhnS5j
aciocqsvDXaSmisxvuIiOjAgp2015TrrpP2wXlkZjatrQ0G7Ng+O4VWv8qqYmZYg
cJ3Cz7OPsWrBfPpRoP1F5bwyhl1aWI/aSVnaMyp+0qUip3Nv8/cWr7/7Bny6nA4X
gcPAR+Nd3FlB4dQlaWJT9pjjhVaYlGYN6AaIvLFKoWBZSrtsygmoupv4MYwr2zeg
O+o+f0G0v6LukC/AyDpjPhFhegaSM09XZKzbM4fddUT9wudAykml5umat1huPLtr
wi9B97sgSya2NwO1oCDTnuXpw+zojQSdnadOY6ivn5KrJ9l9gAGTnnTUxspqTXhf
ZEjFOLawdfR6t0rKlxtPAkwegXniiUHu5CFKRwganUiCEsuOM9knU2aWnehuU8gt
Pg+3DBMyfRqK2X3QlApZTh+t8ZjBXNAZ3KgXypLZlzgfTtw3THu8Wrr4Wjtn/FzI
b9xAiCuRtBbiF0lOWAVYvBDsLOpc6eRp36pYwov/bCaQCSWgWYPIv8C8sXXH1AFo
JOCVeNxAHF+YhIGAUotCzNvj94aYAemzhs9UNCekzN5dxlowm60wc9YKpS0J2NYM
64DLj+SoF4J0joKbTFZgciUsqWAT8hr/ksl23UO9kdl8W3ALHCYdas365EwFla6M
+FeRVBdaqbj5hl1wOz2rStLxoj4jzJC8Uk/p0NWguYB86NKxrH1VFLeXY8KeTdTZ
ADkcOXjZAd09iLvH/gZsckTRPKUcZ2mbQKKfDwlPu48woRpmy/F6gvnaONjrh1pQ
A0iCk5zEuI11L8xFd/OUEprJTE4YZzkRcW5bNtwrRVAfOt9Yal6v5yyOep9kffLC
bbnUin40sr2LiZbhvq2WPPrrJcYT8qSFr0cGjo7FEDoP3XXbzV3AFLXllyWltgJ8
BwVyBgIAzc0dw/ldqZLaep1EWZZcyym/YBpsjQqMv87jd2eWrXcPYmWxEvQF6lGt
waf3lV3007FE0RBcM8b+6YlVXvj2iEdUKl9KUH25IM3mzNGAwJ/3eLrqCKOCd51X
7qHRpC1Ry0GhgkbiR1tc7X5iSsAxplCNv0RwUesT4Ybrc1lfcqRcicTvxBFLTBH/
p6f/dksu3vtcMP61IAloIQnE9E41BU9C1Kgm4rfsb6tFUedgPR5/bC8SbJRWOCyG
Thdh6UTIACQ2DOKcztjcN2QuUZwcGo97/SE5kMF2Hy8LD2BzH5f2ez/6TbJuIlW2
yqmZ4roAssDXXyMmqTffmtBhQfkzoDNqQcJ5kZcsHqssz3Ko70/hSMDGIVCZapNS
/5iJlXFb6CSYtZ+CoaCHHpbI84Jv+0cpE4tKqKx4ECTYKzqk9vaGPQqG38o2LtEx
eqCNWa6KFA96S5HaPoqbOZQxew4ukNutuyIfJNNAbiIB/qsTW/+I/EcE2zZ7dbQ+
lo3Dvm4ez5cuSCnTnH77k7ra+EkFAix+/QNm1GsaZWTz5/FkcyCSH/kXbPACW92P
5+o33Nef0s8KtRGrgu54nZo/I2EYL++IUTZAr0Pdqkmr0LssUIVIvPnd61ybF9aF
lzeImG+ytoOAuDnSJBiz+mu67+tqBfUhXV7yfnZfVqIq7l5T4O7utwq2bcALu0c2
w9Vzf720N+YEnOV76un+Whni5/UFTFvXd/kCYACrMo9+h1REyNEQmtGtOjahJDBP
yWnaFF+wAakRwSLjqsURpUQLNpCDWhamCWkgQ+GOQ7m8Oe/frE7jHWzjYSJTwNXc
/+VV/mkszP3Sg6ZZnfQyU5FVvpzFJ9zoraGjFgLQSL40QDQSSpZjzwWdZtHgy5Yl
us9GVqEf1FDwM1PLwna4mEVchYDBHffiklfADCt1Yo1FZJIdiwXdBS8eaU6p9i9Z
cb7MYEQ0HjySc5wq7p/pNazwc+keCtgnAbGh6QHM2WWxcyO/XQgQx92r1GgGwuWn
iqgREgeBi9/RE/WgNA0FZZgyTMltTFC+gzIlcHz/77GoAxB46wFvYngqgNtniF0J
j0Ftj6kH+Tmm7bRcXY3dZkaueCQbevewaHa2qEUL/rTERRBQFnGBhHUPXM6J+fug
6PhVtiGCpHrZAk7mgGDAwAQwwnZ+1CqlorQMF+rZiyNlHvtjSN+Nz5XgHw8j1q98
CyED5BGd1AYTLHIpcSrswh/l9amh5E4S+/9sngaHpzbXMh5XxmpNEhs6FXTtMkwO
1zOH10XCy6bloWLt+Beb8hKSzxn09n3AgHPWXqS8y5mN7VuGT3BA8tmdulLIu4I2
efP7DKFv1KZ0KEDUIaNyTXx4p4ljt0+wXhxtMFsHfxHJzqsvQzpef+cRnePVKLvS
zdEcSVlnmhYAOuwq1MjCQzbMFQR/fkia/bul5YLxkp1QcaPj1t1bbofqSQd6pgpu
5y5aTLpsCBfKVMG/9QwFpmRezueNACMq/SuhlvWrh63FGWD+9jv4dMceIeCFqGTx
BSXdP1JKOtk7/Ut78lDKqioO6R2e3zPCdxPXHGZlgcJYtZWOo3wrmes0XNATzNX6
HreMwDY/JIFi+6vGV09kJT+NHK8ccfjk73h342LlC9y12C/WHdt92pfIIMpOGal1
j2lFaBppZ67g/+bYUEVmgJDSU8m66GQJpl6OQq0lA7qn+lGW6lHAb11OvsI8JViQ
ek0acKzISSxOcOOCHYxJL+2ubzQyzEMMnvoLdkGP/MmRf6TY529E48YsIFkzHxz0
fu48YDutny4EztWtSzU7DzcM/WkA2dZHkq+iHqtJltt8IFTth3Tfe3vbfgRjMWn0
Dt7pMd55tUuJLJn0DyT3N0n+XQvfjb9zlTQCEP9C0r4WCdQqzll5nAkH9NwLp5vR
3dIcimNVWZEV1ffvSPujkeB4cGT7d3oz7suLeR80Ho3D0SU0wSStyH/2r+BEENg+
cwzT56cqBi7WbOG6Pt4if8GKADO97jAjhWnElOTFgUwopmu8lLLblawHa7O5Pcm1
j/UTEQWGaygrXP57Sp0h7o+tG6eOfH9ZCy1v7uUlpyrnA7XOvpP2OucOk5IhuDTd
i8DXqsqjRely8E3leJgkBGf267sR/zSUaSRaqLYRAdmCIo/NIxtwmCoYGnVdjv0h
fQXHQZbdr4iDaYuSVPGc8DVxGbqna+D3UtlAh+Di0HjX4xPtaTD68IPbQfWHD1PY
QRZyPWRM1ZnCtqTGub4G+W4i0lA27YjhcL+BjzHxAipT3hSUmeSxxOXzbgA+2ysT
NrrnzgGj+i15mtRL0dzeMobQGHt/j9rOIbHFCUrgyLF9uVMalK1YgkTeh1Jp/jjW
umPEjg6XFwbz8GGjRurRATNi1QLMh2YeLDN8cxV6+mvQIScqmCCgmx6hkwbKux4f
FXn64/jSrF+GwNSSZjNsTkZ161bjRtGrPWkUnCLC/LiKmqMIYGwBwNW9YWnfMSEm
9Wv6AoiboJ6lIMqOmxfI0YzlFOQtylpJQwqpiWvmCGM9cYesXgDQtEhx0A7poSzX
jyyqIFeanx/m6M5EiiA3eqV7VS78q5JXpszINdOf42mjbC/f9L9IiIoijjeTSOIm
3o8+9kXkm7cFU6kFmDvjC4Z5udk+jgFLRf+ROs37cXyYE/YeqKChBcYxDEFoW4NK
8LyB5MrLpMhnB3lMYWDCq+GGt+AlgaidBj3rpvAh6GiEhnOpEmciBRmbQmAzDqVJ
y0dXStZNIiTEOhnWFjPqacuMOOY94bmtnkAGO7AUD2PlpY2ZgjuXEdM2kqn1UhRY
L+9Sa++datHcrWYCPPLwWkbrts9N6050TDsrKOpktXlKxsqiFeZmHK6Sd3HkCbdq
/RUQ/05WprBkpOHp+qHHdVRdc+TQ1XYXRBvrc5bcKmd2cGgeSrpO7mFBfLmn5o9b
0yd+3CrMwAgP5F6XB2igZuIoBCNaynCzYdmnjxLcfP8ctOP10FM/UVtaL+FgH5/k
xbmORnyTL1q5HzxPlMck9n4r9C+xX+FO+8aZaxabNe/8y0P/1qiPkzY0ESvModKD
JCU2/dtR51SzRV+Eq+xR23qr7vmnlJQik9mVHPjzxTevQKO6YKjzEc+hZbNZGwWE
7J5ezVoz0j6H8AVSz1J14lAzlEizE3zn5nIGZjwSbe1Ihf83yTJGgvYGCkOvZUFW
SynxzXI0fqLzfM+A1g2xL4zg97f1K3waADQPHl+HORYqC9IwbTeSXss1IzW31GeI
F51tkbBryKBzENcf4KUZhR7Lg4buQ45yksX+wK9efPP6/lyMIbG0MVx/NXBWAaJm
k/rrgUmcv2mhPWGYRWEDtmsWeGcgwt/xd5QwGcwyGC8hjsSkY7xIgtHsgK7u5FQQ
NVyvSKzv33dVDMqf2lGLzlu4PNGlJUfmh9Uhqv3YWU7cCRiLlkEjtz3G5gPYPpzU
+oe1cEyFqIUHEOGmSmMSJ6BBk3YKn9wbj9ZwMYSOOMfNwneb5oHi/dJfzRhxnnMm
qNY3LBptNg8f5ZUeQYuYYAIAnepdT8rNUcRC0XAJZNFWG8nKHsTagzPM8IxF2WmL
cMREy5A4beFcEImfEHIttwKiMcQqdXbHmYD2QXq16bsmttvxJaHD8sYnoq8xKDIX
ikKKS1fTlLPsEYnPxZN9rVzQCHdyRs0BX7S1wFsOSCHu9CaVt9A+G8w3qHRVJ8Tq
bC0gj4ZdAvZnp54/jLwl7lj6mjwfAWrU+9h4VFrMeV8NMusfCQZucBg/KMaXJ0gi
wISZWp2Cv1kRiN7J8YLf4f4f397lbIrISJ+i+aZL7NNSZpM5+4AQr7zp7cxmVE9y
AFqMAPlbsbEv+0lEdC28usJ4hGAnZx9dIu+61UlLrs4B5Sfk3sWne/4eCHSZxhyv
Jy0ae6V3HDnQQYcIeZhIjN5JbbiucfaZJgq3/kTAVwi80LtM2+ai361LbcDl8zR2
9kWwLrBQQS4iTLd6YE3NbXiwXX06aH2SgnaKuWEZdDpZsn2pRB6tNxfVNhjkYrjM
XZREFQoBAk9kOUMgZE8pDigzHAE89lqwQEpiw6PIhW2qOvAvzkIiKVreHPb+dkbi
Y5jr6e7N23I/j1QH0b+MnqHfzu3yG+wBWqTOTR4Ryd4z6M9sGXV/c83Rgu8nRgJr
1gQdHE/xFZbzYdkOZdYcK2ORDYILxYZKdIKZunrGFKxLm0bvIOqdGdQrbxmex0pf
ql3sqNzdvGZ/oZevWANUBnsnlRTrtbVq2YL5KsJyhwIZRHosG2i0rzagLSeJvpuc
4r9Ie72WWOe2kDvkaqswdjQOEocrrEbLkH50UfYWZSB1HmZ1DAT62xhnRZh1DKCP
+Hfa92xk9V52A+MSniN9Jd/VdPQmroiYlgTwxIU7stVmgLjBE/EymguUEsUefgS1
0Qvj4LUMvfTUtyiMLSJjrXVr73sloXkDVHm0H5FOSCzUe+A+IxBhzNmGY6h+O3Au
2ML9s/Ki34HFE4S59Y6R7CBol0HEj9m/yqF8oXuPQR86GqK+WWf/Lk4O16z0lR2n
xs7gkUsDkK3a795BiK9M9GNCtOlmf1zpD47vdsWi3YWZ2fkbGAf8f0OiQ6ExIv66
++FRVFIrVUivTH3ETD52V6bChPRkUO+Crik5bGtOWJV2PNc9IDziyuyOi00Z7gLY
Z1S/LjYyQZCpA4czWSsGJdPfY5lH37mPIxFLV/mNt5J0j4pw5u6OM2NnZe2Ty7qy
iqmcnsT15ACV97s57SDdTDL3iWo40lckfTjo6a789aqk4jrdMb+ztGiEGZzV6boW
lTu1ZSbqa2qkitTb0hK9q0n2+s6rFD4aMiD7gAS15ED99x1eruU4be3XwyiORK+F
is8y7q3JiZTX9Q6WKe+ML1Y2CsW5hLPsiyB0j+Zhv1MkEs9P30WjmQH7T47cRaAt
7er4hGivkerDHgW+hmk54X2BFzmv446MjuZ0CHo4G5/kS7u+7D1mGDRBRxnQpygu
A3IqiH6Nc95MDIrefNGurWdtollZX8bZIJZpowKMBRpIG67d4sQ8c/ifOYaug/k5
l9M5MPYfnz50BQAmp7IOTdAaXSkeQ3G35BkamSDVXTG5vuDtbviqd+8h6gNmXrwm
BRSglVEIdfxyEHulpRiBmQwR4OiuhzFe+5vh4tvBwBLYkLIN3DeOsqkb4zgAyIka
Bszf/NT/2tkhmxPeFFiENIkoit2PwaKOjNntbEOYuWmu6JEph1YLeic0AqeqWN/o
3Clv8rcj2/0YZmDymwTccshC9Fp3Ka1s1/448khal+kBaXHcVVAHgA3N6xacxUuU
YdHcitxYIAP0qQ9TcsAYc3MOrwgqBG3ituBwxLBRHJYeoCg8l06FjtAXUGF3Lb+z
nlC0CLgG8d9p6boIiEtbJno25tFqWQBazEQ+TZp9FloSPAS9qlAWdqX9t37IgXvZ
Kw3Z9v/44VPqOdO8oghHgCVAMNOlZbnRf6u7Q+MorDUT/dk+x7KFINMtpjH/UJiG
t7oI0jTlsvYvv45eg2imYqXggV/dNM7QZjjWHLJQWyWaqgePs6l1ZtFtEi5uaKq1
X1pAOOaghUzo5xB5hLr9iDWRM4qhpXkSgScZwyOa6OiJOG4H08Led+zV4PLHcz+D
uh+tBC/9L/MWLEEcrS5gM+DldphEjmIj/L2LQKu6/R+U8RwWyfPZo/5+bdUWU4X9
wA/v+UaMgsRr7spl17Lsyts9SdXKz+ywJnPJVh0O5qwY3yebjQ2eLHxnOlMjGfHr
z5JqZB6fQ5+axNsWLaaNRlq1nfE2kn1oP7SQeCvQj01mFEycryNAl3e7NC3TZpdB
XWZIT6IinPhRBWmyUGQySHtxiyE1DRvhOJkFi2HExpxsfHRn4BBABzS6f6kkrD4L
NtoTqIkpuUzv2SYvJZHNDeq2xWclGhWH+X+DX+dhpdD/pvsOPxte8pz4ssBYAufK
GTZAaa04E688c2S9Kuovf+Hsdo5VfA+dL5mfKkn92hwUY1F0KfZwBPQco8e2ly0+
MVSaK/XvyToAf5O1CB8kebcMAXi5m3F+Pnn3rao4KoP020KFryy5cv8R0BMuvftw
BKQ9UhEhTNsTCZ2dqH+i0o5pngcdFWnwcUxYRqi8TrijtzcMipLILHabguma9w8l
fOuz/KWDOeMfIftCyr8/H3XZlJEFsdr5TTRs8GzzDtp4IpFPO4BANVmzy0hIbSVG
n3HsHnP6obYe5MdDPswxRZVICIdixR0IKfA+y4HoeSylHYPulrEn6VW6a4TNEqkh
Gh4QXrzGat5cO7nfQhMjiZa3uvrqWXQGR9Bllu+PkvzCvpGr057M65Yi4utzLn6/
0nfUWpt/tnYT6Y0drbocr8KXR65WDF+85Ozqbdz6Iw3htxRuJPAz8dHCRXTdKNP8
6StsRxr3uKGuO/RQ8TVf2iu//A2yuv1tSoRk+2B8UgEuclVYxf39bqhVZpcEpKju
sKgUXwln/6Y9zfnqYTx6TdGfsghLdy8r1FVDE7oeh6lHaTrHE6O0zfz0GlNjD9FO
M1ifsAWaIgge/qmPLDZdUZorB94GkDmd7oNK24nPipqwB0lgWr+hIF1ona04kIqc
0+XRyG0Og9ysOwStVKigBuo2WCKrLKUZ06d2a2SYM3JsJyKCAIpr3ByiIhcW+Yyv
XcC+Zd4cUiaca7aPUiMI3Zbc1d+gtNSviPzbJ/MjqvrNXHd+omvXgge6VaR9FGKQ
TyKpPHoTGOkAOGINMdPUjoxDTNFthXlOTpEL1ul+GMkbFrG9TfwZSEf3v4mHwYNh
LGxnWpRHQUdy7hj5dZyWxWTuggH25R2iN2M9EaiAZ4zxNce7wKrAbU4+5WzPGojI
7yMNAyg0oY2pbqem264AH4zij2J3SjFL4LWSA6R6wKv7JqqO5DcH5ioYv8zbIAX7
FBe8FDShaN+r7UsLqubiFQIAaD/lYrdbGv8NTPECddqPXBa1O511p2RVqL/7KWHb
8tVGaAnE2S0wso3b86VafupyUSQXac+UkVHdd+yJz/6fQNc0ucgNW5L81SfuLMCc
thYM1XaPZyHBIDwYh6UCagbby4x/0BrzcLbsPFC/HDM7xpJ2nEkUijcLmCu9uwpA
UZfBa/ySu/SJeb08xm81pzZw5i2z5Wf9g9dAOzDlbGOuIAy/xBoE+FSAWP16DDJa
qFsm5Yt2NThlis6CJ2jv2JMjdTDIE1vnLj+AL8wrH5tqDf+E9wdGHgCa9kmo1fWh
jH3iLXEOSzXvhH1+wkXfx5zk7hWTlh/6NH8PIQbhQgM6jl14H952ggl/juXJhgcI
VS9k4fbdf0qZSsieSqgGj5U7vo97Y0O+3OAqhgJ4hmNM61Q2YQNec+UjPICBeEqq
SnSy8n4TnmIZfYSPt6V0q3JY2+tZvGMP9Gk5WqxfTAO89Jch/gbbWydWcNvye309
MGmo44v/Y3QPOj7sOA15Knr3rYSIAXClvc60JI0Qwf1oHjHNkChITPElEUOhWavE
G8y89+Uhmc0M5X4cV6ndlsJc3YDvzIHZKnr/WdLgK9v2MHyTQb24JD9EhPmTm+Sd
4Gn5PSM7BmqC0piDEDftZhbPUawgUH4GzstaLT8Ym7X5EW5jrNhFgA1uFpt09Q8O
KoLRAhwtqoQMFpP/JmXFj3LFWmH288VWIz+dzLtPpEMQ8nL5bvxlkVPI/8hZFJzD
11qj+Aw15n9DJN9+9YnWwAaI9j3Crmf4LHBMJOMG4Odiv9jbpCZKsNtdTZe7uhXo
s0eeJISHmTGy3QkzVTP4r8AXIV2DotFz8HlNP37zMPVgQNJDyvcasALLq3ytkTMP
DmvNPuBPmhR+luykIx0jIWIjwh9qmgazP6QuRFbAaMhA0l76nkwbssLuhMkAmHKy
izVZycSNqdXLeOfSWBTHvqnuxtKC/4Mh+92FJyHqviXu3eOgWThkBiNZTFfFR60Q
+dBKEnJdtMzX+XyK3g5v9IlDMndr8rZpUtBrAldLC5nLtfY4RbVk6BwJDpFW/JrE
odCqU8VYxG6TlRXlNw0uG+YQLU8aTMiTlXZGOcnIZ0cph1kzuRxGJJHmI9t91vmJ
dJNcjZCjnyoaR+ynqhNCg8tCMEl1kcajDCYip84g7rjNOGNOJFNV4Nvx5A4rsQ3n
4qNKU1aEBgBpp5+iRH1gpeiLWeaenawggwO3JWeLrBb/hpaMdAfGZ0VqalFEyAFY
ohNoFN+QBK0nWp+Oxu9Ddqq5TrGuXa667yp2j9pdZGJpVapRDuoN/Nt7OnOIElXQ
XvhwLRcMIkoURMp3OSiFzHQxyEzN2ajcD3UlqiYJY3n4qw83j7sH8wfEefo+S4ai
hT7uX0/LEwUhj+pCttSQCgrXy2NYme4bukpO+LM83cvjZSISRvfLRHhnJflqGdxW
B+S26UIHUyftxrMMUXY+l4IYmoadqX6fcy1owI2llf4R3E3GlQbEUckdtmEoh80S
ILYr245AuMrbQx/gKaL2WFqKRwCvptftylGZ3NmfLwCL5egEAdD+Fp112d0m0Q8n
aZPgVizXdcTJH3kFCx5ita0Sgjsu2U5lOtUOYT3CkEfInXfL0VlH6KQT/S3XDy8g
zWdofQaGqHcbGIwpf2U3JVbnSP5Qe0k0Q7awhcd2gap4SSMkb7IsVaUsSfi68NHr
fqWgeFvNxREJD5ZCaxncGZpQKXWlRRcEJ6sJV3LZxA17HurE++yee/v6D38F4U0m
A6Nh9GJ/sF4NH8W5VODkRLtUTycZ7/xVGMV5yfx0OKnpd6XhyfFtblLwJEZowul/
MK0lj8uAJx9V3cd3h/Kf+Uh7bZokskYgrNNisPf1rEJJGcEs7o4moAsCL7u7xZcJ
10QRWL59vZW9rLNA7eqICdH/CsPaehHbFqS0aRi5a6rbzc0mRnHfRIuNFRBr0H+r
cnutdQp6dykrHZzrEVTeqM7iquYhP/nWxGO1NMjXXbUw9Y5Jp21CayWPCJcXsQAN
dkAD6vp/c662WQuqhVLOrdVJ8jEv2rBkpscecC17vIcdNOX7Sj9SDnmdCtIFxo6f
0LFdjMY3jFqYuncHg5EHrZmhjeExPXgvLQlA/fZoW0V0O9dCc8QrwlOOyDoIn0Wr
8DB/3mT09irDPVxC6OgaLX1lDdPG3+0O3hq9m26XMBqJurAQPSOM3hjwnd2fJMmz
DInbuSNpO7Iy6Y27s0uGEWJVXwS6/U1rOEv3MUKexB7vWyT6nKMWzN+5F8TiKLop
zW3mvK4duC2Yh/oU3gWU78kSbUIEG/xbkQG6wa7r16H4EO4z2xbv0Z/QSsANb23h
GMdAmKqAI8WfbZQcpj/HV2xb12+0HFO/js0LS+jy5gBozi1DwplRhTiIX3DxPpCF
e23FVuq5hfbPKsHK6yICJ3UHYImLF526Dcou4MVgrzTQyRUDmdZ7en6jwb+iZui7
b68aS7ByQV8Q29WwKmGd+MY5hB2Qdu71HUhJAIrh/33ybSRPlsprscBX4PlfSpdS
pUysS6JHqZwAqVB10VnXNHCI6tdcTlOwJNK1iLnz4Pu3bWYS7L2wVx22r/UF0ME1
Xlub2hu1h5UDlZGqD/g4iSCnrM+5NePRMmGIc3aAf2DaGfDFjfceg1kgJ00zHqNj
ZhNrTR7iYgmjKJfJCNLVhsIZt8iLWa+3bP1tUZ/qOYvW+SdP32hfMPYROhcGUyVQ
blNXF+Z63m0cTpLUQqxXNCZlbBeuhSu91o9WEjha+8vAukoq17KAsVwZZWVLemKQ
zck2z+ci7uBKoX+hfS1KlssS+a78W+jvWAD2tlJgeSXU92+u9gK9zBDC0aSQSqhB
V1SgtVJ6DaJ7WpS3/4xp1qWSbK5fezXDWBUzT6z8cy8MfKVzlVKqo61fu86eTUUF
z0JoFxrD5ksMHvEzMrFFMW0tjaWxtbu/SYQQeOD1sqVXvr4Jt8JvInnp9F/sGl/y
E5Ljo1XIrb+jiBlhyeVR5pU96YWef8K1xaSvg6WKpK5xWAA8TA0VGTQYVh3cVXcV
1AnnO5NeqHCxlMXShDtqodYe5fODiAGPcMX8/ShHcODVOPG7ChWNbgc/LIq8C2sD
EJA2dYNYnGjlKfFVhABpYVv9Ee6TXIhqdn5rUpoOrfoGmTHOD/IWuIy8batyQGHj
+CE9fEL+aSq36r5bZ/Rfpfae43LED/4VmxAH6xQuoo2nmj60f3pCXXQ2vtQi1bLq
yJIqqhiqWGzpzLMQ6X/+QbLkbn0QXaL0Ax6miKkbuI7PuACxa2KkemW1cGLPzuVW
9fX6aK52Le1dSZaV8qxLRmi+u57ZoFN1RI7AxOQ6kNnQpBuQCfuluiK0oo2Sa1v4
ipRK0rLAlLY8q45kcsFPDFN60+P/lZjNjnkl3u3LNqnKFctNqW5NWRC1u51RjqvI
nPLqXfjtn8VxspW7tUG8d/V7KX4pvlEoIBexP4EYnoK2dsZy+FG7T8OmFwYSbBix
LHJZPmQrv7TF6pQfOysbnvXBQs/0+XqouKOaJ+9ba793AkP6akXpaFqvt4V2dL1y
IFrbleXJ7bFq9/uwsEqmgAYLg8y2yliEI2QRcglO8XnqRVMYOhl96aQ6aIg2j0At
Mw+wl+JCs6FinH8Mei9Dydy4FIk6uKxshYQ+SIBKS8Ld0RWDj+LM33OeQqMRqu1M
aRzBmZuysvuw/P5+F6RbDQdPPb729cicRRGBHENOZ134sKT6NoUFrgJVK4xgSMIh
2Ek5FjnuK73puuhVqvUUjmIK2K9nPYMRofh2oRkVnVddj9ZBIS1AWshChuOY4hg4
slvFJt8B9V/RZuQhuFH3SjXRpkJN7g+DliFweGYBKHb7j0CLwpcvhzvazgK0pq4q
Y6SRWnNuSdqEgV0K1Qrpx+qBBS7JGC5VCSdEAxLlUnsS2xJCQQsd+VE2z0ej6oLp
5ekrt0mGVmCX+jdlxnwZHiKqZvGcwLUcmwmOC7a3Y7XSLVh3IUj2qaVZwSW68xHX
q5YGOMkamkPaWt6Sch7lyt2SDsVp0ZAdpt5ppM9a8W+KtYACqPb0nnxGBLQqc+uT
givQAf+VB97FF9gUKGoaBT3QAMXUINPzpnFcyCynlnod4fA2ZGCkkXthzYcLUpSO
8IxGCpruRGq2AQJ0VCjEL2rG9/1IBl0FC05H3uZJotM1k6ILzUx+2saworpM8j0D
l84gHUfsPMhUZSKFN0WfKd/+enenniW6vsc3DK7drSqZZsBtD+END2eyL1De/JuJ
aXKI51LtoDcpAmNv4md2LHkG7sAPi+PfssFlyvT8g1I5wDMNXai7S/pj+Iv+LOlR
5jMWaC2+b/Lt3yKTptikc/HTa8+Ews8avcyGk/HovzluSfQYXZxMkIIeG8KrJtjn
GNpkQXttiP/5Wja2M0YNFy6rAHWVzsIhZsQ8NyZjF4hLeDk5bwxnQ2f3cD+pyPyB
pgq9MeBoP229IEWqVZG5uZ6AcZQA4Mh6grKrwu3NKrCAo7c+ZZmfIpyxrx9jXF7s
od59utewFgchYdlRdTAKG8miI/kL1iy0TcXrCEujU9a7/k+vGXRRhNgYrYmDnwUF
AaklrfZ0Md4WEQThj+jOmdeoiig8o3G4ApP9BBrhy7phH4t0ZqQ6MawdpX6BOtGb
J+bCujcKWH7V6XGjlmq5GvwJ9ozuqx/n9hfLZBGCN1yaUXKrxp/LS5uAx6EusRB/
o+FjmzkS4W+I80EUp4m8/ZyMNy8hCgWRbAUhuLoBx7KqySxNMw9xXNMnoPdmmk+x
uKMvFZ1MaRJx9WXKn3ftQMjjyj2AJh8XhctTBNY8Fz0MFPs7H/qe78ynA/urb+1j
c2w00tIUNx8fEElTE0ByFJ/j4l3r3ah32WVJsZle5+Mc/T51ZdGskZeQ1I0eGWQg
vcU7cxlb0cYKrDHXPyNr+Xrrpnn8A7BCZe08db7Z9ed5Nqh90S4AkjE2CMO4Ii4B
TOE47+1J0XR7oGLkie6OFYxmw7Bibg9dqY9ph7ya+7LZ7RzcG8mLH9/t2kgK3sas
iiiEJTDjJBhLA4LEuWJBUdBtgZm+FsTh6Cba18lQApvZ7A1FAA4RgvgDx823mcnn
iq527oZoVLHGJnZfZ/2u90tI05a6VvoXYln5X+7JY9N9/kSuwFImEt0C94KmoEn1
K5/5E4A1ai+gXjcc2UCxUbXinCrnG1IaIJDrHSFRYenCZknPpYe7mwWtZIeMsvDP
6Ul965huTuw52gKUOxk2C+FUueJDr9Ks842FZ2fU1WR7dkg4onEy5zaRElv3olhM
4J/dRlxhcp5vCJcnM3IAWk351rellDBYlcE9wA50d2U2nF8fTac7UYP064HgnS4q
mknjlMRs9+1mihjMlEyAbOV2GUqoSSqjs7FU+UTAuorSj+DUlHYHUtmZ958qVA4+
BuVzERSvEm/1y6OFdAfw50A4iB56k9uF9sAqPWF7kgwLc5zIRFirfeJToX5uWgVi
QaWlsnb22Yn15Tk6UTiSdxey/4eXsRPuIFq9xYP5OhddE0N+AWdyCktUAY/Xw7qr
o2pDS93ZTSctMrBZNIB/DTjyjkw22hrL1Fg5eTsHP2Rb1ICnCCmhHxgyGdf94rSS
xnKBsrMIm5j998JWAg0J2c0f6Eo1CfL1s7ljEWALBf0rNrH33jTAwojX5a1OnNW+
FjO4CF2k89Uf7fROxLFZKiWEfyIaOf4Gi7+KXGaGsOdeMyrCAnartc9pTSw6XaLv
hePS/K8cUEuWpehxk1c2oNyuArXttU1JbmrsFsySyjwshQmxoErnUePI4g2db8XY
MaJaYwO8b5TrahGTYY7c4VnU4S0eQXs2Fgudd/5FX67cM25WnNHgOFNSATkHonua
9KZYaIPpAFnFhxJTg3S5Vh33g4bQu9/gUOkJ55chnfDoxK4PwRE82ofva/m2GYeG
W+pCNYk1vWEgp0CgO7BoJKh4DoJ0TTAUXU2QoRsZz1jXOl0pY+395HsjhXtBNYSa
VpxzhIvBb190te4eY37+WJ6BGv4po/jlvFZDFksnrcZZ8ZLXnGhRzkTD5cJbSyOU
4aCGjv0Af9o4yUikZuD0zRJ9/ccqSzfyog1Y2GVM/d66YyI3gIrsyGMqrPvclyhs
A07+hlnTL56/W5AQqAzXxgxwNgZ5uFZVY7Zn5vwSGDKNAmlD8bWk2emTGHqhsbfj
8HWunMO3XSpvf74/nEKKFKhCr973aAfvG4JaMxQzhSIAsWsZG2LZL+pvYvCx5Fv/
RnhGq9GvyCxxzy8FBqeEEqetzEIPgdldK33H0XaXazKg6XxH4nLOje8jl5S1ysev
DL6dYD+V9V7GEukje4tKSDU83T/RudOeioLhIHzfF92f2yugbvmHHCFoR+vVRi69
WS6jIEVoBux4fw0PiRDSmpaP3RLr5EgP15mEEOL0cX7IoHbfolLgn/sqMqJ/Hz/3
HTNGQCr1LwAr03pl/XJ6k/PztpqqC5lcr8A8svQaHHv5k3hVXkU55AGWkQaFPr9J
Iy938015ShB6j6RsX+VA7NJYSiALLSuvqmz7A7Zlm2ChLNzVdlid6s+ntElR37Sq
Z1teJyMXVI85o4Og0gViZ5vsm1Q7TROn7g8kvDFywm/QrFRKTagcvvcPkYwvQz+2
vtTzNOG2Qxn5uULAmmQ5oiM1zbjBAqNtTcjPJUPQUOdUlREc+YFLV+YPqRlRjHtb
DzPOAQ7PyVIkCEOFt4GyOl6A54FQ3uWjGmXXsxXIkZGfQ5gu578P061ICt2FgMeT
8f+PHM6bqjXnwSGr6u09BdMyS/dLvXn3kFlS8rcqfpSzNbhUYItQDxF6azOreDXK
ZQk/Kr87jtSG03HDf6MC+VmlndB3evOBGO4V6oo4jCPWBmDHX4sM6Ciaa3OwG/gc
pn6uyZoHCzdhd4Jv+hq+Oqyb4UZvZxlDYm1qSVZim6RE/r1m9SwDyog1zVfeBfVn
To8loynvWHatsIApiQfTQNpNSsK+Dq4SjxtxQrwEqTF1Pj/9yY0nGZyFUH6+wDdO
Fl/Qr9zmnTQkcbOzF7owgWwCmk8Gl1ALA/SwR4jVCt4=
//pragma protect end_data_block
//pragma protect digest_block
KfVhYjMovblkx1czb4koL74W86g=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
i2sIZAx433WzzUCRy2rzi5fW38aZfNs6PTdUcxhqmj1JcQPRwugLhD8CsrCr1mhX
aMUMmLQnJrnLWUsAhBl89uunYXw7XNHMJ2/C+oss1kuqI97GhR8YEl+9GAqs1vsG
xCmDJ5CuminVe8oKQi6RR72UBxJPemxtKysfBz0Vlo4CgSEqKOWkVQ==
//pragma protect end_key_block
//pragma protect digest_block
BBZpQ4lkmANUli4RgSgzpk6qIF0=
//pragma protect end_digest_block
//pragma protect data_block
1g9n2c1tvG27hkRHzsENJpV2BVBZipSynT4AM8qrf3vVKn10mwAn8apg8r4Hc18u
Y7b5JrTpfHxmBpBNZ2juN46SElJ9WRTqZqrd6sDaSHhWkI6BSkRwuMTu+X+dnqkD
la8r7Cefn2+Hzxnq6BnoGtHaTa+BDFM7SaAgY/2GZmmyiGROs6LRm1ynOmn5AH/z
3FlK4uwkCEcvagcL1LDpf/RA+AkHU/M+Huy5N6KVNZZTEwW/DLzp69eejAqaX/Hh
O4ymcZnqNIX3zIZORhJU/227L29vdssr9zzpKYJQUUC2jbqGmaHMRmQHbiIqiHxv
Uf3Hx9l1uyNt1KSPspuONkgv+AQz9I7VUWure2oUOxmlsXrc9BY82uBfYvDHy6yq
jR0+qYMjVjjBhB2EU5IcNnFlnynkY04HoZChWTd0WvT/Q6gaJ/4CdLYEdLVFDyFN
YAc8M8YNWgJJd+RVQOnTG/xUhKqUqwnRC3C9Te+69GdUVB4Du8ksbHsUdznTTi+l
WP0KFIx6vVjsG678rZiQP1hetHk9oYUNuUsVIdtUcSFYVHuKKQZAPG/0iBlNkdIY
pgOvqpgWIgJ1OIR/exHjxhY73nQPZnievghBl+Qa1UQjDRfWsJvj8EHrjLo0hwj2
s9lTwwb3fVBV9pQuaN6D0FlAVC9ZibFmBLATzlvTvHBoH/skfAhiEbThuxHMJw+W
DPfUnjpkkdNmhbyNC/Xj4bcHYRmFCkiY+yim4H8yUYpTcqdJGy+t4XFw10mhx6MB
lBzyNoFbajoo+U7M188xmYglyi4iwQsa9yzFs7jOPW4jL6DvifQe9BkgMpUDudVO
Po0ULrpDSMx1xhZCP89wM/im/fNg7LukpRnbMY/kexPSzCL3vzIzdfpA45kFidGO
egjEXn8LAVSPURAtVSl866Qi0yZK5u4+OVP7tLxUVP4h8meqIPip2BpUKZdxujMS
ZPeNw0g6c6F45uBLaiGqmw==
//pragma protect end_data_block
//pragma protect digest_block
iU6+f7WewKV+Ek37NEL81jMF9I4=
//pragma protect end_digest_block
//pragma protect end_protected

//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2r6dKdxDY7I1pvXsfeaYOoFfTstxolmBTX9p36RW4MVbfJVxKQtkO2MTj+wIBC7T
ujI2TlaOIm9p4ehAhdBsmWQ20tCf6hlc3F1fpKnwLl/0RPCCzqyH/myr4l/vS6lS
/VGhfpVYdLKAQBrTjYRQdt7yY4HRtuYDArP0w3lxxFPSKRaY7nmpiA==
//pragma protect end_key_block
//pragma protect digest_block
p304yLmP69PhZByiKPL7EEmJR8M=
//pragma protect end_digest_block
//pragma protect data_block
9pTze9CDFHLRN6EwmLPLLCiHU1T11XEi4t48pe+LNf3w7pFeaK0XBq8iJ9jvdYVu
eBwSl+6enr52mNrss4g2YiN5fwMQR9ShUgwgNgyyrviro15kJ5fbpxHECwuSemCE
oIHwkuqjoiFTkVDs1QI9D0R7V9nab8P0uiRIM7yAkLXtVIuo2ePZreyuUjsCqWkn
p3IKqJ1+a5dGy72QmrGy/YgEylqIxpX+i9bIVGDCO05rUGGAX6Vg/s+RxLoVp0Ih
npNu1yhaXVTNwkzY0y3VProJePOwRts3JIgDs3zkQL0tMqVnquSqVvHDnO77pvzT
tPHhcA2I811b50u31GvKH169dWvM8ifUPph+sJu3W3UyZrsuMzanb4w1DOF2WwX0
whA+c5ta7kPTQGK+xhNLqO/ahgLAQqlKT0P/J2xAkrKCi526KoE98gxQ1UGxIMRE
69d1w4MGquUd2v9zxw4n/V/wxy47DghFdiHIr2E/liHelGKs9aHw+POAUHVwsiI+
6KuyEeJPdBGt+XBMDteOnd0WBS7mrKz/WzwsyQdLTin9RyRexFmF1t+vXvhxMiWS
MMSD2mjIoQG0jBX4tDIvDNTs9uO9LGoZYtwitN3Kzfrwvm1SiuzZk4WYOWM5SbRS
U1Z+oGtlvi6kzLEe0swZangu0od3VRxSP4tcDjToy/qjSq12qlSTcPUoxw13kjjS
2QJzbLWXsYv+SgRuM6/4wp7hDa7qK0mnpSClyWNSRdbrRlsINyWZkSJNDy2bcXyC
umEPcK9KdZBoIl4InRkDWOZlagttYgtlkzYvtEwG9uaMwfntsvjTJnozxxhHcJgM
nFcZBVJeB1FcwcJucFOB6wdihb+fOPezZewSvviVdlaqfJcAbRT+pZwTbstu7+ut
XFVZC6lPEAURwETJa7hz9eeuSvuTAvzQdkLTSj6+xjExE3/UG6hPS0xaXZKpZW8+
zj5ce9kjUL0cMxzvX3ksmVBUooTCL1+O+it1hMblnIQET7kmYbmVLm9fKHvaaii5
7iDANZcYOrSQE3k3wYKgc/4zV+wsFHMmUpvxO3ZTUB13VLq+xyKauEPKRfhuz3e/
2rzlivQwKGDDO5zZ34jB2U/vQ2Ph/g7+uHCd5o1sFdLwAlyvcFgwhkMhNrZhC6Xg
ROzKG3FUfGBWsfzW0iWIw8Y2TtKPzAtKCNa9BIXKO/ftWa6Xj305WPy/LpLfEYPP
NxEwv8TzKhHywcXrGfsVtuiYnNA6JUQtIJl5c1MrVe6tbK3FZT9sjrEo/pPolT7U
KCeRIokIhMFgcVWtLzkMVSBx4y/+VyJDSfUqAz4juDdsPa/e3D7FPFUcxJ+hCufa
+Orp80o3wn3ikBuxLtjDPHYC04kFECDsbqUenasf8xG1jTtaeHmvIO2eZkMhLigO
kmvkkXSkm10khCD3s4/wgFf5k6CjD+4ZHgLgiEg6BBKmN8ahwqhZsN3iJkZ3BMes
RCyQjr5Ss73l+aYc3NUlSZUD0lDUbklPWdUDClBOId5zIIf9XmpE5syHWp1EjV//
GKIyP5hZnImdrkLHY964/lI0j+WWl9S1kbWkylArO7BUwInpdLjZ7/GnUTRvQ9dy
IROgNZU/LxYbg9/t3uKEaRx9QrTpx9PmQgK4Ti2R6S5IreF97jPih9U+Q2+5YLGq
LenkmN9OWNocKonvxMsuMA48Qn12gYkanciB7vziOMPOpilFIn2DYTvAWVUjpkQu
LCBTouj7Cz6CADM4LAb82d74lmB8nxCk5MEtfVmTqeX/etiNnwoFQKoSIouzL2g3
q5VBbC1szJhXoGjLcGkj5MKqkW/RgTP00K/+q2YsRJm6q1Y+2YeTfP2+yVgWdAYW
RKnvm7rIU6RT5pfPBkVp7bJu0fJpVh0lIz/Va71DI5M0vaFNnZDQhOUd9qBSMKnA
jDF2D1dQ+qI53jvsvP+Jvs1FWV5XY7uz0lqjNl9NNsmKC7ti7L4kqNi71c4RJkZG
ykzqzJ447GGTWwbZ11uweIWkGyYcKu6vt7S7sgorP9Y2sqjwloEVQ5H3Hvd2ByX/
6OGkrB9pPhhqNC8/KhDv7NaI/7MXTBiZLr9g08C6tU7p0B3r+6Kxep01nY/XwOWr
ExLoefJlLkW/H6aFJe3tdsIcLb/4uWBadrcw5JFvrw2wtAGiDzb1JTFhfpZS2Jn6
l4gp8qI4rkjiA8pfIlbVbH2CyXcnIgGbl2scZq2zoaa8P7HB3O6ZkMITH9PGkfL/
B1Ny4VBg1bst46toI5aU0AA/MM+ylilku4KgmBmogswZhqGJv4d7K9oM4a91hsKw
FJerhdA9gKCj+DTLbVeB6bmX5x8AYcwEWrl3g+qgtdo+/CDpqhtgjL9HcxqNePxW
7ZWChZXs6Jtnc5fv7VjGjpFkGX9IFVNkDaCu9bauKC8iJp/adt6v1GXV7Yu5o7uV
HlVfx6mEBNl/NPtyPmiK3UrwH94xp4X1sQhynEsG/ohOEOA7WeiCoo7XyvaDkrQN
smb8+/OhNfM7WB4eV7bly+eOla8mwV4P3urMrEHCrLu/a52FMc4Kw+mDBk9UgrF4
eGaKmCduMZqpXvUFIUYe0WNcv6wL6Sdy3KHsJE0Ajg55hVxT1ge/H1vkQ9FAUM9r
Ik1ztDWtd+Ix9ayU070TCk3Qg5sWYmvqHibXSIsXSwJ7cKMBYYqrKcEuhP81a+oi
f3XOk9nCQ0Qd2bgKuhvntCODnLcS92kVt5DrhCxLoYEpwTzNs9dwoWJzUukGN6nh
cdSHKpdXaaD1NwLl1hGjWD+RVSGagNUsYR8dZW469o6OUIalvMcdh5v7FmWy/TXR
g0/MP0+RCK6uRizGPTFyve9glD+JdQtuGQjOuPY+z8KAgNcPB6V5tTL2yRehZe8G
4jCwyMcOBNUZbItZ+CQ1kSUCA2jBB3s4vZK92EoJRi0xLodh0n+G+Cd1A6zUBLgo
B7vxjThHJs1LZrRU55SUKua2sY6dZYRCfjCI4MIby9AEeuBUVpky0fC2cVFLwVU/
+aZc7YNEXnPt+Eun24OgWtux35BgRQixO/dIlrqDfOqPMKUqUUEaGO3TQpvbdIyc
VBafh74D5Mo5t7VsMIYOF3229+LxorKi8Rr+DHIaPlfsKsCmuGhPuM2haIlN83y0
8ruqFteEIhgeVK2mlGIxByDVbwRXx4zxmbO2lZJZZf65mnU8NGDfCRTAQHf3Jr6J
mziukogsxOC7XGSnjKQU6Zi4kkEpy9jh33jRSUHbXygowQPi/yCojOlX00FZ6E0+
Vtda+jSEhmooaAuPS27YK0W+rVXBXf6xwnjc/6gHcefi58E6baPbLX0OWAu6FpPD
0gEXDe/ajRo542v08uG9dPwd6q4G1ujzh0ZcwYO/5pc7058KrE/Cw49Cq3QB4RFi
OWUq+hz+W1sFER+hZD+ZLf7Yt1h8BstvIcF2KIrnpA+2RcVzGfU3kHKiIUyeg8NZ
lTpE7pjzkEzuhlI4LHa9iaAPYAmuyg6dOP9yjhhNOXLLvw+tRNIwtkfO17LmmDjn
MGWewix9J/its8BpWz8P8iwgIi2OM9XHI7U7ZdEDr8+nKNdIqnQZ3S0E4bLrPtow
+IypGwpCLicCkJwmjSmVy2vuy3GmOli0gFwQSDnsKzi9hxK33nNMbFIsyNPRwBNK
+D0+GigzalQMjPCIDS2B86i8MgEkGgIf4z+U5OPZvfn5z0bjoUaQi7VLWkSfJB3N
bnX487IH0RoSZGpHtBLnBgOA26A0JVR7y3l9PKUSR8Vn2b3dvGr4a89a/3lRAOrb
Wb/ChdLmqxxJWizK5s870pqiZ7AfiNg/NzLqLXgqgnhM2ibO5/8yXuXzC+kIzgD/
HMEkPIFMvNg0Q8UK0KeDii7ECNXEidL9rmI1rGnw6pKcHnXy/W2rLsMm9SSkPfRN
zROiOb2mCN1bhKZuOwua6rJlvBMnnnaTBxlBbnG2zguDVv5zW7su2eCfBSNmuR7q
ti09eaQuZ7ldHgHsJAbwmMcAuI6uBd+UtBHVfwLZrgllzR5t9lZkpEeZr8u10XDH
xMds6lhm95PZWiuS/7m1kheIuOLZYe7LQbUXnS9OP7CRYhfXi/J4VYM9yQpb74dC
cBXw3x7nUPg1RTOf5/BBCRdQhOHWnpshlVZQpca2sfVXDO/wC2pqnjvgBfLWej8t
ft6eE1FF8wPydtD5XXMVwfva8PRTkE5gTInf/3x71LwKXXTe4hlAs5v/ZXZSbts7
i/Rw2BCoruRE+QVGkiMqoC1jjOPOoQi1pchHqjvwj6FYxidf9tmexQxHBb0cKU9J
f8QjgyspJH/pwnr1XxYKU/opIM2NOleRopTaTTjVIeB9oSf37j99Hx8+b4p6GnZo
I9bm7G50M36GtKdhNpp0GTV5sNS2LVV+d5uJ4B28BYWBjrjH9ku7mXfp9mkfZSCt
WA+FSiwHtNpczIutamX3ZT/GsXGb0SxPxMFvqxziuS5nuFPTOduPPMugknHDlOgX
/+gX8dcEAwrPpK1+cJiDhqj8OQjiVp64gMCn5XGHtjXq7ig2FEhzX71AxrYJcvIW
VZ6OF+9Xwq05NGhaT/QnHTJEKYsWuXLYCaoYRYdvJU8q0DOkM3OwiN0UbLq5XjMl
LK8gHNToMXZDZVHz3kRbeuxTGEBqIw/sSSCm/+U9xQLNhK7RiCy2VH+CnyS3S9vF
oCU27E/tiYF+utnM53mDaozdYlGhxRv4AjDuvjorqNywMS3ZvuhrYyQDi8hnqbHG
yRy5WMBGAjORDHVvxoAfwfryTjk8QNcLo5vQecf0UsV64ruKHSyDUzdacjYHjaas
JZg8fAZgz69JgHzpU758FOBoGE7WuxRELglAt4VqJMv/5sZ4gIAu5EuQVzKy1L+E
EN4GZdq+KpptKxAQmEmxeLr6gCK7IboKM7pGlLoej0TlBCFMFH0LzbJQDNJDREx8
4vz/aVBoS2VeOegPYReUemGCyB3z+FSAb1CQAXn298UChp3CFDl3ndjO8jmuVldE
a3MFl9OPGBhyDIqe5GTzfhbJVnMmJfAgpxwAh0Fx1SpekURipHHduPxWF1bbKwcF
+DFrhxBVKZgAcyYypW/aceWfK1dMZyZR3xKmR4z98LARwW4ZxdZiOdCz9mUY4jKH
KJtwCIKfA05TtwVP9O8C05I1oGSvf7TGHE953hR0dBasrcHdBKWD2gGqe0KHCHFO
9ed0+dHdcDe2baVJq63GG4j65rECmr+2rsRptu8kXrWutJMHIQRTErgBR6PQ8rIc
0w8wxqcsbb8vcoQ7+QzZz2i1g5sA/liUgGcQ6RcLd/01xpm42Fi1fBBeMvz7cGWy
cwf0XVaQ+dMAF80ENvzUed53u9lIv0fTFXOwVlcb2CWD60OzNxEOpHU6oyLTqJl0
gwXP0VoerXxL5JZeA+fBkwkeVVZMLWhoVzH3dmIRrAtP5RH4xSNqcVWQgj47E2t6
/L9BxcCn0LVDzTn7J5xRDlHWw9xMUt9qh+RccyxotqA+PlUXncdptlr5X/xGy5di
0DOwGs+2DXHslK+FYKrvfZTPDR8J7s4yvrvA9GNcs1TqNnM4QZ6DTEgIu9uRHYQo
wQhQGBhgqGmtgptKd3Uj8dhEIoaDWhBih3U6Bb6Z3vPGm6I95KBUuuVM4TnhoAtr
UFp/WpJpnFl38GiK+Cn1OSW8uAz2Kcz8+l4ZzGzLYDordx4zST99oZ8Iv7S3Io6p
jQn6+I3NzLRGZ3/9eQ7XA7Vqt4N6VEtPdF31B138CmFsca3rD6LShXWKEaZwPtBC
IQY3+CJb+kZx4uzIsZTwWYkFdK9MbrR6tL3NBEPKu3j+ijklKDJQoOJPBvLs1AZN
XstfiJuM79lCUlam6ttJVIedKbLS5E7Crgr09tdGJ3aL/XjHVygjp+ut/evSNABg
2VLDufvutqPMBh0rsUPSbfz+s1M8w8lgFGgC7j35truHPG/MAvVzJKReBbQSTSu1
7GGKDN4yxQ0+xFsj9ncV78XYOFppniXhbsxRx3aRSGtfa8Gukr40NM1j8wZS4dxv
tHsz0xrrvaMd+tHAV0EZSIUmAA6Z2jvfyrVDkYrVC7osKSidgxHTmQJloKCaXmGp
XU8Sqly/r9/sHiTW5VajrOtm0GwG7z/CyRmivAQq92s/nq9G61T+o0rPlMR+T+GG
EdbhoiPv3M3/tfJQXVsVoSQqmH/ITZbWipG3Uxrv1Ly+N8NbTxMes8mO+D4EuSc9
RycvXzTPlgfFEd0iCsyXe2BNyWvYQXsiBsMuJDY7qEQvfxEtNrQ2wrJxjYYpB7hR
imGZkqTlWd9Fy8o+df29u3TZERcOG8iRdELOYVroy1LmJAmpRddo8Eq+202Ke+FA
z4+kSALglLz4wlmAcvezZvYlDABsq5UYlIsy4sL4+KOcvwZu93mwMGC//fYcyk6X
iZ26vXqP1lKgQezoLRbU5WXt25AdAvYaFMOFdbOb8ReIJyuD7WsUifa5rpnPTrpt
FyKO1mPpg/3ccMI/GPyM+DBx+tM9aVMoATVYA44+8jRL/bitDwowyGbWKgYKPoLp
QxtEOV02+cG60kcRzwSwMLZLe/7xuG0f+4FsBmvK2vUU7psR2fTpLek/OfwRpxMy
SHOdfwvriKaXitkW00CgAdfWwQYcIJ5a5qInkqERfHoRK/YwOIuMhjeA+ZZn30pK
vFKBuX2FybV6T+NuhOTvCQiu9rNrGENFQ/+Bvx7fXLpdNsmgp7IGoIow9/3GrRGI
NuKLSsUw2pk6SFGYk2OyXWuVWqAfxnSpqR8EskcyucQauP7TZLNntYqC43AQtv1E
Q5hSY3uM8by1L4Bepi0DPos+xaqw1DqhrCa3IeBQI8eNjoPzHP2mQ9W9k9bv1BuL
AG2SAZ3ya/MRv7N8BMdItg4joS/nuf4gcHv/x2c+IyZQBNuYZwOkVKnb2PzyJKCh
y2/HmjFJH9hY9Lp8VLbZ2GGZ4FJB83hB/HcHoa4n5PGZlVxe8Pn6TYWnYGATowVc
Wi0cXMqcddLMW7AfZZKGiWdmJnd8au1old3v2EiFglcOlLcM5JoaxDEM7iy/V8um
P2HzrkLFYxlQBh07uWO8OChrYu8PiegrxbVAONd17kjJDxYmjcDXYbMUooIBvwQY
rML8OJ68CuDsvDGt/5eU+2/7FcydAF231ph89gUGHbep3pyVO2AD+FZ9utOBSu2I
bKZj1wOJk6eD9suaUBMN+U7N/a1Sj60tIgOhQG4GHM7xRviyxxZ9uE9+mEUrgG8g
V6EXs+Nw/s2YwNP3xbmk2ssqtvpdlNZ5C/yDw1Ni9dOMadSgpyailNG7Hi2MyrVS
hvn4375D6IlkNUwz51BHWMYl86HRwmF1ncD7/Pyp/X2WypwUwX+3Hnez8ZeSr2W/
5t3xdJP2a4fZSX5i/on3xE8IJICHhk5Q4fYv7tGD5oLC2a5t+mHNtbBP9fef12BF
fJhXOTPYsHVvXYV+LrXxYL7CnY/TYuDMnbB7nrKDg1xJRomx3SBRFq0CTAms/qqc
+6QI45WfH9h6yJYtd+Da/QwzO+wcyczpA8+n4Yqv6fZmidUq+wwfGtVcxtmGQnvK
1ln4w4PUVmeK2wEx6JYPHmKiUG7t42EdfJ5vF213t0zvYWvMQrH7a5e4hzrKbIYE
ArXISMWbvm8ArZW2gddl9HUtBeplnz90oGhgBbHHQbwx7NiN1wJdt+rQEYZPAX8Y
T0YWQ6E/m7Wly1XlfXO3Ts8FXkeHPKcyl2RntprhwFN5vHIjAcVHWu4gc+YoaEg5
PJO22tMRUQKj6C0XLh6epvfPxPwdOLFE/EvPqb8SEEbMe/rV16Dt3VeqAw8+kznt
7R95EWPqdcA3X8xS6B3yII6kkNwbmu1GohoHJmpP28aJmM4jwVEs8rB80hIqjIK2
3v4+K3mMn7+KML+wIDheovcrDIIW1sWv1UTyb24jK/q/zsbD4GS0iWfMJS/m/2gl
rcekPBg7i1kinCRgO0fk5fC94ec4YeI7/am7hd24KTzbGkoExKa6KJnyejXGTJ3Z
zNl/9DoHyOruG4wgupw5OtwTPZsA862AIFKvvByhSLHHgtcw2p+OMcZVubfW6gDZ
A/x9od5HPOmQ0NJB9SMUju9wgX2zg7gBCm47Fl/0hwe/WO1JFoZjom9JdoW6FXJO
rvu0soNgSU2lFRj4jGv8cXET+4Tmpeg7O8x3qxC3B27L79IELBWq2gadUhniOWlB
nD4/t7XqoehVCzey5tkXcg9TaSx1tvgyJbZr2kmI1/BkjIwjoOkOZedCOBvN3ZSO
peBsISL6mqKDC5OBfSURmLANHawtHarEGOxJHlmhMMM+DJ8k/922OsA2ah6FMg0q
DDACVViKmJbuYpOyxxNVL10R4jDcNVE9axP8N+oR+F82ROHad74oPoIATp0RtLog
t4Lnk2BQI2knHDeDEPhkMPeK2oq0majzyQfNxMOd0Elp4Q6tj5thSrvUopFypMYA
7LIFwuPxdcQ4vPhuD8Q7VVvR6shlCk31qaEYPqds79UxNf8ktShGvoAPnlWIPWBS
Qmix8lXtDPzts/b1I3wqVHMQPRbPBSsAI45bhcKuShN6zDbh2ASq4gl1tf+kwdXF
07mtQ4QF4wOMYikJmqE6aisUzLr+7hPyw7l2Nic53cCqOFMBJ58nWJd+iuJZgljA
x4jamRenJfG0k9j6Bib4WtVf+bKbbaLAoCXKjWWNvzDMrTdIvLE0oZqRU5MFLY68
BY1uAwtMIGaz/ZAAgs7WpFxxfKwmgPeIyKjdyg5ldiWET59qcds2D942X+9HCI2a
VzBtUmD0os8NKekqn40RrPO+tDLbuThsN7Vn9UMEj27wcduOV8xR+uQ1XM8q2m3W
aqWNGUy5MhB976akqA0xQZJBod04Z8cHFpOUGXI7QqrgNvaO3/iT7q1ew2x2p6qH
Jl4cxYK8DPuLBxWgv5aihm8Mz/QLOx5P8F4ybn+tD6qpvtKuHIys7j4qszgDvyIW
6oLxKWe1OdcvILYY/U+UxKVgRdagNJVKn3xxbNQse6pdzg7yP73Uy1wRv2QA895h
A+BX/iv5O76uxhy/aTLihZDGBoFdVbnNfN+7+W1rwdL3LFO9FXdjmm5LEECFbmd1
lgmV5xwi4A/14qERP8PHJXIv5uvVELXPJ9DFjMwFz0u/HsZtUVP4pRp/yM03CQNy
dg5l7IUFVlci022V1pld6Rjem2m8h5grXHI5HMdKrNo/P94ZCI+XhYw7s3P9VftE
deaAu3Ruzpjv1LmIkaBjLVgZhvPr3aolvsQOv95CHC7MoBcAs5uGYmZEmAjFeFuG
z/S3g04UEounmGQBy8laJ47HhNjY1qAsVi45CyZ0yLtS2627JUlDrb89aUo+sX9P
cY4GNjXDXG9ei+wSYwVrdmB7HiWju3zejJcQb3JhsISM6GbTgQ/W+K8yYKUO94Vh
DEd8WRGqB5KOrHtGfpX1fVUejtAbJaVyELS6AuN0ZnmrNq64j9rF3qH7b397a5kj
lI7Fv68PbYZlD9IqxioaFns0mB4UZ5E08Fq6X2JKy9Ff9jcdL92iD1yoZbcPXnEB
1wY/4kCWDbw/3JY4H+7oMqVUoVfH7nXllVMKMoj17jUV04xLPKDIfHN3pMDWU1A/
ukGI1JfBGKKYJ5Ldvjl0nZYZTDesEuK04juTdSdi68kH0PdZU2IRcndEVp2XBtMk
DEKt1ZUHZk1TAeaqVz/tCg45DFvkw4U51Gei9cvzELtbvXl69bx6mBqvEw0RqEHh
CnX3XAsliiIk98YcyDegp6ijj0KAwoeqy0oZmTx9X7W3acTagzMNxPLF96JHhQFo
7Pq/DdhpmERG439FTORg27/s7tmQagSd0An1o5zgQy7hyiZvgF6FHLeSU6I6f5jK
UZ/TGGb5082yYMmJcQSDU5yc14X+RGrdkgErvDcBUnbvoOia8SZeFNvyLOh4yhMD
2iXkwzRJiNc9k/e1ORmg5B6UOEtcYsHgjIcMb1RWF/K+mXLrNoBsQ0oOJbS+vs4j
I21F7QWwrCRs0CqxMk3900Ned9tqikmNi877d6ON94opZmxFKj0N18XF0UsTCOrH
m0kJvhur93lSxjK/GTaS5j4HRNiFByLeevHoW6oWvGPGtHHG1rvSYGMgOHOkPzLT
FcMS75F6HWz7vWoK9exMGrsfmrOdzplHHarW/ocPBaOsdzlHJR+wzCBnXJVnnIfk
LveOpKTFUg4/14SbLlhkNTmM5jmygO9/2lDQ/Mk4kVuMbOd3Hs7SFPqZP+w3JJeP
NhHPnw6+gnGqPpEglTzIeY6GWEITnp4P2CBd/LwxRRmLiH3MP3UU9zineEBujlyL
LzhqvowPxW73iRnPmHnn6Kyda9TuQuL+0L/YGeXmSKIQZsHbku267C/hymoRsr30
9+sLJYzyPeagHBQ8JgjuCIMMXbz/ML16u3Uf9FAbf+88coQ5q7pLO5V/XzYSSuNu
hea4SY7yVJnoUikHWAOoiDA/lfugqT70m1pcT1lCDdC0o41mgPyK7Xxmu6Bns3xc
mNDmCxRdApp0Tqsdu2dzUwCdlBjbpOB3dZx1gCK+z5kRwh8xDptfBE8l3Vf/Zyyt
TgsCNrWq5g/+fiJxT5ed8CdhlzqD7yHe90/E2AAxBD29JL3kBKDUNOE+RQC1z+f+
T3u/rHFxhuuyUvJRsbJAgl25pRkX2d3/YGWHg7qloB5hAmZNb8nRlByCkpoYnpKu
w812oWfQEqNxbEzKM83XsOxcQ0YxMWJm96SmgxW1LpOde6gkqqvlonAN0pMjG51C
r9fLuDpwhcjghPBKiEqUYUGizaet/aiyFYWhFrnmwW0ldMleI/tl0i/gABBwh0n7
DGy6du2F9uBNsWtjJxM4y/rPbdet8HMDk0FnyAh/dT/Nz0vxegqRu5YpZrFT6LU0
cXuASQ8DvFIAC7OjNxI2fYv0dEAjtPMDILF5hcOscFfWmDg6aGHFWRF6u/pvpIqg
Iprga1lmdqaqbqrmK3dAMCBsiPYO8NQLyY2I5VmsUY4rC+WFlIRRPPeL7f6rGHhh
5Gg2EPl/VMDb50mMr1skO997jGU956iAVKCc20os5Vk9M6drsLARpSPbLcecuIC7
TUQASu/jUIMPr4U53L0IL50tuKHEIAE0CGodtppo9pkemr2jG1yc+L8BJqF9Kmvv
pnW74vticollx+TUZMm5WHNQTNc62REKIY2PXc17O8vp/Skhdmhu5qgAM2PuN0bt
KJFvb9NFHqNonFSENJlniMmA/LCyfUbBhw4DlWMdb6zleq+rMh15HIBU1dPqID6a
QJ1BElcjP/7v2wBx6kRr/dws48Ego2F0kkemltqlNjm8oSyWslv+zzWObeD1Q8fY
GObYy3OrJiO4FDeGamJIrQmdXxx8sZCsthWXTGtE5bg9xv9x7ke0iUb9jGS31VfT
G+LnC6wYNh5Hcdb0QGXcF3sVRGmy8qWwSo7SLauU0nvFFBY3WyemwBphBOwRxjlE
o+ozfmgw7jq0yi4YshqbNU23beP4+CB3jws63hrCkPX7NvJGe5AnvV/jZDiEPeF0
8TQsrFnmVdatZBAln2II005jImNhbqq8or3znzIE//qcXVXPVMIb8OC8k7JiwO6A
PJcYReo9ydCIE8MiRRyMD28a7Tp+4LO+ZXGAzeq7VK6rkyhkl3zmspDFpikdrvNd
8iJYIS11fg9dOmfD2fZs2RP4JsioPconehB2Vglkxl40SApvfpSyzbUVQoTIwewj
m2uH4rtgfbmPoRKGv6pGLOaXu81ow8HjbnMjlxgjiv3AGdSkSWrW2itusdp6+SPl
4qQP1FYtiQSP0ItrI+CeCyD6FMYE31Im1raQK/lIpj0tIFdi2O9NjkgB03g4rPbK
4QDJS30VvphM2HOTLwT7GxNHzuJmo28LnMLw0nwvsUiNp8+2+FPAUArpPtht6RsB
nH71KTPCTYq1ufF2YLP/pehEG5+lqxr3cbjHayRpmiTFiZ8qhChK1T8nWyUGAzl/
VarNSxNLmSVbfCyS7UZOLaIUsYohWakLDEBWNaXIpDmiBxb/YfH1EGXdLdEpFNkf
KAaEPDtKTxugIhYY5PdJ1CucaNAzhCWp+SfObTfkY/2fWPKNn05nYkbfdwcHeZQU
h2IK/HawgvZrxDQxxEcbKSpvJYdZdbIVO4m9NY02QsdSZoBKpPmx9vx0gK/DLZ7K
fdiO2BDdOQz6SrEU6GZVCGjzccWTp6Jksf5JGflC4dD96TigfDLeOelmgvod0PVb
pHYHNBtdkpmuYcekpPUO3/He4s9wl4EmyUwmAHYRhE3SSMK1E9Dz8rafw70CaSgr
eoMPNI+if3HPTJ/hs0r6C6kkNBSsG2HrLm1ys2OS4sTr+Em2W1B2mQ5aEPpx3zej
418fjukWsma/L9nvreZWmexRV5n/Hsq78e4Fd2P8XXyyyNaKUcLOgbgp9WG19+bf
CU+GqfZCt6X1OhI6FJ6wpjCZjatNU+gvoSxl2vQbAJRZTduEve4TPXiDxkUsUWgY
k3sKwxnKz6Y1gTdOA9iC976NdxRfPExwn/+Gck/C19QVCXen9UC/RTptoVDTs4K8
XEJEXHDbuhcfqXFcZMksycRi/yJA7iwJqkxT020pDxFqEeYla2Wnrtmn+JYLaIVI
rwT2c8mI9YcARhNoebTW/WnT2+pw9gDp/18SCJxeOF70IK1age873TqWIub/Oy9o
7t/M8m1wdrIEVvRxA7KflS8h6XwjOES0dw3ZnVHABBdobP5ZHHWm5zIEODBTHdQQ
mTqdbnnDsNIWrsxnkyqJFZ6MQQEDjG5DjVra/b76vkkxI6b8duCk0zmqq1vD7wxB
m2Xw4jecYkH9RylUQZMoIdJJllBIY6Dx4JknFURuR4Ti/l9y+jMbbcxVvwcpGOVh
j4EYahhEIFDkCW1P5j6TfHpYNtjLrW/rx1E08pFUZosCIva9O9nx4SeDj2zwEMfQ

//pragma protect end_data_block
//pragma protect digest_block
1r9gcj7zJel+UhdggRQprh9xYbI=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oDS2gXh5MQvhkGBGyonUWxLpwsN4zLVc3aTwktM0FyMJiWc8pHa7w6ZHnKyyOm7m
lht+uWnqYyr/geCwSnbE3e8SMFKXIxDbf6RekWsz6sUYSrcsw254up9xb7PEyQAZ
V4IM/NLCi8qd+t87qdrdWQGEY0fLeGoWQN2SSwcFGCmoFyCNvRXFNw==
//pragma protect end_key_block
//pragma protect digest_block
y6E3sDf3gXgFU6xjkf/Xp7U/GQM=
//pragma protect end_digest_block
//pragma protect data_block
Rll45f9N9j9T4/p0P+DmFYoqKooa6NCWuCWXD4HiUpsHT28+Xuh9rjy0zxwWlG68
v8PIFeHNPBTZKWDhvlLcgSjuwemArlG8i0sdAfLH3bRfRv+ipRxPeC89HeB+pH4J
09KNgP+niavzrYXcO+Lq8fvAxZRcWTxJe+PvBLAfuiyrxo6Ar58I0TtKBRk1rc2j
veADP5fBCn3vkptP3+1kjMLhJblffkF7pyzO6IqM+b35Lqjcsi+bbsh8a2ePKTuP
GcLH/CS1Y5po27pB6LHDu+JTgspfahjvasWUj+bGGEYuGNsE4zqdxQSqdJ0mwkDz
KjfIx7Q1Wh1h3MGtSmy8gTd8ec1tuaGuqLM2Y5TRYxDYG7fffIGNSddUnUw43CWt

//pragma protect end_data_block
//pragma protect digest_block
Zcj2IAGKSoFnvGIervTaVZafEaU=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
PYwrtYC9UPK0Ttj8w4uoUfWtgKY1h6e+WzWAKb+4Fxs8TMTCgSq7hF7XZ7KmSLsA
zIZmHHZgZxRedlYIw9qp7c+4bZcilyYo0510L2HPDcn23FIhAi0/d04Fl8yU8b2H
7QjwLznuvCUt1UQKb5JOV06K6mwf17QWFJXIVmC9gwAU2l5UMSfjEQ==
//pragma protect end_key_block
//pragma protect digest_block
4jLwsoG6SujRcc2tyW6yel6Hk+0=
//pragma protect end_digest_block
//pragma protect data_block
02Gi8GaW/KGm7zI22cnHDi9u+POz8QOHUS7T9MnowPx2LUL5MmHdEvBlKC14kYjI
NHTr7/63WsRvKJAsWXqOA7ZF1lr9HQcYsaW6et9Qw4LesNBQtVu1RFj17wbM1ti5
/21EJY5B0e/FxhqHaYUKJA06EXxqbdXVFfIoMBEinJ6Ud+pLegbSINHuk7VWg8EL
GxKsP2WEuwYRnZCjjxk7qodU/TlItZKwyTxUhCoQqgwxz0EMJRxLuoTnphm71+Tl
vqZMj4K/EdhXddor452/qD3w0PHECGPSq4CbehSdXG1hRM5NLWmfmTt8Oip99bjl
dk+o46rPo1VNprw4KDA7p0ngCyh6xRo+U3TBZo+1zJJ/rPN+7w5VMkhwzHKM+aUT
8AVco872aFc1rfo6TbwtyWLTxUfiTPyXc44ec/T2LsrIHXCxPRKWpXSqxn+bBeGQ
4mMekPfonUcQpegcfUFGMsBcRFzXYGF8auPiYb8a44JFywaLgJRRb5s+sVEDmiI8
qQ4hXQVUWTXwdgHgrkmtMIf0x9B98+4Tu773TZDuxBPPbo3EWXh5GnflDnxoDVxq
+sNuUjmwTdixWl4lZQPvlqK9Xc3fP+B65cmyDci2OJaeZSvu9ezZkLzQ3TuzKX20

//pragma protect end_data_block
//pragma protect digest_block
zyRJsGXPhpuafuhkEzKHxaHzpjw=
//pragma protect end_digest_block
//pragma protect end_protected
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dexvbN2YxYAL1Q6qwonu7H6et5LLQg21e4+udn4A6kdoCHUjCtdy2AtjROUh+C5n
pnS6cqQGKrzISlC1x2q+D7dKWCC8s370o3SuXhl8TaxtUz2tWhXp/YaNinqjfHmf
oT3wVB2AOlRu4jZkLyO5TRLFQYf4T/yvkpeJqk1JWic36i7rcAoHOw==
//pragma protect end_key_block
//pragma protect digest_block
1y/d37aMWPtVp/9jMKe0i6KCRwk=
//pragma protect end_digest_block
//pragma protect data_block
pMj7PrcEeggTo9XfS24ouybPv/OXoedE7tprGVggka0F68H9X2K8ek0kmtlNsaho
mZiRY/1jQMQPEu/tm0ZEPhGagkzQmlBiKPXLeszgqHtS3swK+gDn6IN1Wdmq+Lkl
LZBa1L56j4BH0q0ExigyGtgaRNJCcJrM8/S/AvTsfUVwqfmg42OYeFjt5/JXV7tm
TCuM72+BW2tW3lh/L0Tl/m9UHA3qqzfSygXmaBNw50zY7ssH/KW+ZTdr/HA8mLc9
h6/5bzLDL9EoXygDIDyCco2Q/PoZWMXlbSTZlxrfWL85bFuWMYAGBdBsndB7cpdl
rEoY1kaagnQpb+wxdwjfVCl8J+TSA6snVe/c1LTz4U00n5pbFyfl2kEDftGWBCI4

//pragma protect end_data_block
//pragma protect digest_block
+kfvA5a6hygjS9QkMKw/5YM+5Rw=
//pragma protect end_digest_block
//pragma protect end_protected
//vcs_lic_vip_protect
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AS4IJscnZDTjd9PS954MzXDT99TMKrlRSmaXTJ6G1wuAHP5e+HHBb8y1khBXPTZN
KFOcHc7Ch04w8rQIeEAxuKuyBhPwNj7TZ49qlYqGid61T50LtTio1yHANRjmF/MT
1Ujnlzvyzq0zHGH+WlWLyJIQVXJEPdV/5hbIqg6DZAXQG4jd+BhQsg==
//pragma protect end_key_block
//pragma protect digest_block
uE40atvxHeBahuTRe5R1Y+C3hg8=
//pragma protect end_digest_block
//pragma protect data_block
jlpREOX401r6Y3xLUpwin5X3T4Qrcf1ClVrSOQ4SVI6W2Mybc0aSkeP0WD0HLo9A
nfcRTDORyiTImRcKKKa65RsmF6cplFwPx9CuM68UjcpG4nRhK/calFKQTPlFgXwI
97A3+BbbJY7c9VwbBUrO0pdYXlICt08rofM2O4mWH5i00mFdQQMYBx0dzc65PvcY
QARI5b9SnIKtEqVt/JmxCr4um7kGCdTE1UTqLJNv6ocdUVbmCsG7gYut/iPdxolo
sgOAvfBp2ko1E4eazGFY9wtDwQnEZ8VvsX7X7inGMZ9v/0OhS7AJ8HgI5EsS56n1
sRhfvSvNWmJXjs/iF0r7Vlv0h24TsNl/dA7ICz8dWslXU9UA0tnNtNPnQYpcIzdO
6ckXLevY0q3IGuHZsSIBBDwyqmOyEUoeYJLj6/SlLTk=
//pragma protect end_data_block
//pragma protect digest_block
EFdoahSfJpz8iIVy0mPXrjeYy4g=
//pragma protect end_digest_block
//pragma protect end_protected

// =============================================================================

`endif // GUARD_SVT_AHB_SLAVE_ACTIVE_COMMON_SV


